�	  �   ]��?Eb>5���r޾�ln�J���羫�K=�v�K}U=�F־��~�m^�=}�	>����'� ����ͪ��/J?H-l=sA��pbU�u���3|>d��>Dծ>�d:���x�u@��Ȭ��\�='�>��9>����1��yG�Y�ԇ�>�C?/�^?��?QI|��o�d:����>����|�:�J?��>�P?|iZ>���=j��I���Tc�6�K����>�?�>�u��EH�KL����$%�?�>?z >��?2OU?|g?��b?��)?��?`��>���_ծ�9�%?�E�?=Y�=%9Ƚ��S�L<8�C|D��,�>*?�FC�sm�>N�?�?#�(?�~R?~?)�>: ���@��͔>�<�>��V��>��?�a>c�I?5r�>axX?6p�?8�:>x�4��C���G�����=��">C�2?�g"?t?D��>Z��>�H����=�B�>/.g?�4�?��q?��=�?�1>���>P�=�ި>xd�>'?�GM?Ֆs?�K?���>1x<[ٵ������1a��+��:R�<8�v=;���n:���|��<]Tp�%�輱�Լ_5�'�C�a^���`t<�_�>#�s>(	����0>��ľ�P����@>�{���N���ڊ��:�^�=1��>o�?���>�U#���=殼>�G�>����5(?��??|�";��b�8�ھZ�K�b�>�B?8��=��l������u�h=/�m?��^?>�W�%����b?� ^?_��=���þ�b���@�O?n�
?��G��߳>�~?�q?���>��e��?n���yIb�t�j�O̶=�q�>{Q�'�d��6�><�7?yB�>�b>��=�p۾��w�o���?3�?! �?>��?(,*>K�n��5࿠��)��J�O?$��>�6s�LS1?V�7�C款����Jо�q̾�灾Bbξ<೾v���	��s<]�d���md==�� ?Ay?(5n?Ck?1�ʾ�b��UV��$���\T�����20�-�_����=�?�<�n��&�y�����]��=��~�n�A�kv�?[�'?}�/��%�>մ��"b�u�̾7}A>,I��;��қ= 獽n�>=\=�h��.��*����?�Y�>d�>��<?�i[�>�cw1�K�7�1$��C�2>P�>G��>��>��:��-���B�ɾ�A����ҽ]y>00z?׊@?<Vd?������-�����U�,�+�g����`�=��0�S�>�_$�J�+��;8�&mY�o���x'�W[��<���u=p`j?���>g^>�g�?`�>�|
�{G5���@<��3�=7?ӵ_?�F?���>�7�=g�I�t��>h3n?�O�>���>�c��U!���{���ս1q�>��>!��>��^>ψ#���Z��썿�[��?�<��g�=Ul?��VW���>�FK?��2�m���۝>�$r�y�!�`A�!�	>u?4u�=x�I>>�ƾ΅�V{|� `��� )?�F? �����)�>?"?���>~�>ND�?۾�>�"þ�1;\�?��^?�J?�A?���>R=^g��'ɽ9[&�Ŏ+=��>�p\>ݒt=j7�=i<��f\����K*@=��=WnԼ�i��=?	<�����O<0��<�#5>e�ؿ��@��>ξ �
�WXɾ^H�W����𖊾.��a��o����S��F��a����f�8�v��+��g���x��?�r�?�Hk�e���퀑����� �sd�>۬b��e�Q��I�>��7��fJ
�V߾"V'���[�2�h�x5N�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<
-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾t1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@[{@?�+����:z>=��>��?��<>��#�F������X7�>/�?̀�?Ҭ=epV�O�Ӽ��d?�!n<~�D�k6��k�=���=��7=h��sQ>R�>X}&��7O��p�}�)>S��>��漧$�(]�4<ȸV>�J߽|��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�����%��18����#�=��=�w��#�6�
B������NѠ��(U��y	;�D>��)>�A>�R|>�?>j�=�S?�t?���>�;F>Ja���1޾&�c��*���D|�WѦ��x��Ǿ�j�������tA�=�$�����"=��=�3R�4���޿ �6�b�n�F���.?�q$>��ʾ��M�H&-<�mʾؿ�����륽40̾Q�1�!n�S̟?��A?�����V�]���s�������W?�J����鬾i��=

���9=��>�q�=\�⾐ 3��xS�6t0?�N?�|���b��R*>�� ��=�+?��?\X<I+�>�O%?<+��o��Q[>޲3>qۣ>+��>�;	>����`۽܈?��T?׼�윾!ߐ>�j��	�z�A�`=">�B5��F�(�[>�u�<������V�`e����<��O?�*>Y��]�������O=�=��|?hG?+�X>i�g?F�J?"s��Ц��K�_�|��=0�U?��[?+�==m����ɾ,����.;?�Qj?u�t>��v#���1�W$�UO�>��p?��?r1����x��Q�����	#?y/�?��]�v@�� ,�H
��Cޞ>���>%[%?!{v����>��?[Ύ�v:�����v�W��F�?$1@P1�?,5>is%��� >~�>zI*?�=���!ܚ���k��k�=���>����!F�P�$�fξ*�C?��Z?�\�>�,�@����8�=Ҕ�����?0 �?e��c�=xx�l�`��c��C�'���;�͵��?ý-��h�4��Lƾ�	��ĭ��2�<�]m>^�@Si�����>�i�a�ؿ��ǿ�3���꫾,c;�P��>]�>��'>�둾-.h�����K��Y�����v�>��>l���V���u'|��_;�JF���|�>���H��>�IR�����ǟ�f�*<��>4d�>ц�>�/��w���֙?h���IZο������OY?��?⎅?��?<E<e{s��{�z���`G?�Ms?5:Z?L��EZ���:�%�j?�_��sU`��4�oHE��U>�"3?C�>V�-���|=�>~��>�f>�#/�w�Ŀ�ٶ�(���X��?߉�?�o���>u��?js+?�i�
8���[����*���+��<A?�2>���L�!�<0=�OҒ���
?E~0?5{�b.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�˶>��?��=Z�>�W�=����f��:>r��=�$[����>C�J?��>ε�=�7���1�j*H�TU�"Q�m�A�`z�>#!a?-N?��]>F��S�E��`$�2�Ͻ �)��ļkD���A��T�+K<>�H>M|>�BF���ݾ�4?&y� �ؿh���t-,��a4?�҄>Zn?]��t�S�����^?��>���3�������U��
��?��?�	?�Vؾ3�ԼNS>�0�>G�>{	ҽ]c��+��W�7>�B?���5����o�S��>��?F�@�~�?P�h�j�?Q1���:���BO�{�I�]��>4R?����6>��7?���<�h��ޓ�2��Ŷ>	u�?�Q�?П�>�bo?��v�G\K��E�<��>nz?V$?]�=$-4��Y>�#?�-ܾ�#��^�ľ=,?��@��@�lR?���JԿ�������������=�<	>[jg>�����=�w�;����"?��>�}�>�9�>�q�>��E>W1>{�R>'Æ��� �ם����^<�"��8K��� 0����[����C"�l?���oо ��y�/^l���H�4�#��gJ�A��=� H?�8??K��?��?N>n�is�>�����=k('>�fa��8�>7�T?�t?��R?�	�=If��"�R�5��Ȍv���U���> ��<�Qp>[��>ND�>��@=V}�>�>�S�=���>�<>�=�=ۇk>���>P��>?e�>!��>�C<>��>Fϴ��1��k�h��
w�s̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?%���z)��+���>}�0?�cW?�>!��{�T�4:>:����j�2`>�+ �l���)��%Q>wl?�f>zu>�3�Ye8���P�}���d|>�26?鶾�E9���u�v�H�fbݾHFM>�þ>�ED�ul�����#�Hti�B�{=Sx:?τ?L:��Jⰾ�u�TD��mPR>O8\>�V=Ye�=�UM>�pc��ƽfH�l^.=���=��^>�)?���=7��=��>�e��D�O�'��>�$}>��Z>��+?��#?/��;�S7�����;H���>�<�>~�>�f>Z,\���-=��>SX>��[����<O�ѽu�T�TJo>˶��Z�O�qvr���W=�͞�x�%>K��=��ս�/���=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ	��>�e����m��Aw��M=�q�>\�H?:b��� X���7�0~	?��?7l�M���o&ȿqu�B��>���?v�?e0n���QA�J��>��?9�Z?:s>לݾ2aU�1�>��??��P?'V�>Br�����?���?ڗ�?[Zc>xK�?KU??��=u.��\��K����q��z�<-d��dO��Z����=3�n|s�����xs����:�I|?i<(��>��)�>Vо���<V�8�y����G���E>E�>��%>;�|>d5�>ˉ�>��>E���I��������n�K?�?����(n���<l��=L�^��?�L4?�Z���Ͼ
�>Q�\?�À?�	[?�h�>����:��u濿�{����<T�K>	&�>�S�>��qFK>
�Ծi%D�끊>�ϗ>����Jھ�9��_���xA�>�`!?��>�ͮ=K� ?#�#?j�j>��>lUE��+��2�E���>���>�.?�~?9�?����+\3�h���衿�[���M>6y?�J?��>����Æ���JC��J�풽��?�hg?�Q�:�?0(�?7�??��A?�)f>����ؾ�Q���>I�!?aC�(�A��L&����~?^G?���>����ֽc�ռ���z���Q�?�\?dC&?���z a�Z�¾���<�l#�<RX��^�;�D���>L�>ŧ��]�=��>'Ȱ=�=m�E.6��Mf<���=�w�>n�=�&7�ņ��y�<?���IPԾ��=��Z���v�RO�=U� ?����g5?�^d=�Gh�t��9���I���?�?�S�?/Й?�L1=O�^��?B�?o��>�?�����꾼#����ҽ`Y���,����<@z|>���;�:�O̞��3������N�����>���><�?�= ?��M>��>������&�k��FI��f^�
��7�8���.�b4��`����!�����U¾�}��V�>�ˎ��z�>n�
?Zg>A�y>�P�>�
ٻ�ȋ>nzS>�}>-P�>�@X>-j5>���=Ⱥ
<A�н�KR?�����'�g�辸���[3B?�qd?,1�>�i�7��������?���?Ts�?U=v>�~h��,+�wn?�>�>B��Uq
?XT:=�;��<�<V�����	3����"��>E׽� :��M�Ynf�xj
?�/?B����̾�;׽�o��_�=ҥu?��
? y��D��n�S���6���]��q�����R���o�4͉�YF������R�6�n#�=�f-?��?��:����~�0[\�< ����>���>y�c><ן>�D�=܀��B7�	�~�?/�����z��>� �?��>K�Q?�;?�I?z~Q?�g�>>��>:����~?��+>��~>��?uD??�=?.M?��?y�?UK?>Ef����5=��C>
?�D?o�"?HH?�s
?e�����v=�=���������&<�n);��.��Y���=�'>�Q?�%���8�������j>ie7?0@�>��>�
��!���.�<���>`�
?��>���˒r�w�(�>A��?�/���=�)>{>�=�����j���0�=���iD�=Gт�:;��M <Q�=�<�=�9[�{����:�-v;Y�<g��>پ?.{�>H�>���	� �������=�\X>�lR>EZ>�BپZ���$#����g��iy>�i�?�m�?��f=[R�=~U�=���,���{��D~��1��<tn?��#?�*T?�q�?2�=?(#?�>��..���h��cM����?v!,?��>�����ʾ��։3�ҝ?d[?�<a����;)�ސ¾��Խɱ>�[/�k/~����AD��셻���V��4��?�?WA�S�6��x�ܿ���[��y�C?"�>Y�>��>S�)�w�g�m%��1;>��>`R?�u�>l�M?+&w?��^?��F>��2��i���˙��B�<��>��3?�p�?8&�?r�?Ol�>">&{��۾���#
�m��m���q�9e|U>l�>���>�:�>C��=7s
�&/��e�=�=7�Z>#c�>Qƨ>۞�>�R�>��d=L�A?S��>_���4��/����V����|�x?�_�?ƣ?	�=b��d[^��� E�>�q�?�8�?�m(?�\"�e�=�|\��ľ�]Z�4d�>���>D��>Lqk=��ƻ���={��>8��>$���M��ޓR���?Z�=?��c=rʿ��t��Z]�?u��wٛ<��t���2��j��@�W�'�=[ ��Z@K�4����9M��a�������C��ox���g� ]�>��Q=4�=/��=�k<�Щ�0�K<��2=�,�<���=�(���L<<��!��B0=n�h�+�u��b�<WE<=��,�˾��}?�;I?ݕ+?��C?*�y>1;>��3�[��>�����@?V>.�P�����i�;�F���� ��O�ؾx׾	�c�ʟ��H>�`I�$�>�83>�G�=L�</�=�s=�=��Q��=$�=�O�=eg�=��=��>RU>�6w?X���
����4Q��Z罢�:?�8�>�{�=��ƾm@?��>>�2������zb��-?���?�T�?>�?<ti��d�>R��`㎽�q�=I����=2>d��=�2�[��>��J>���K��S����4�?��@��??�ዿϢϿ3a/>�a9>	��=:cP�?f1��<_��X��W[���"?h�8��{Ͼ�"�>���=R��ɾau$=o;>y�u=c~�&jZ��6�=�^��:�-=_�v=m/�>�5N>���=�
���:�=Ob-=��=��L>V�;��>��#���!=���=�x`>mb >Y�>P?-L0?�Jd?��>��m��ξ����z�>��=���>���=�D><Ź>`[8?�D?�K?K�>���=��>�S�>DQ,�
�m�-侦6�����<�?i��?�*�>;tT<WB�����>��V½sq?��0?xM?O�>@����Կp*�ߩ.��%;=�1�>E��>T�9�=-'>��x>K�:���2��=9>H��>x
�>s�>RA>��f>ԂU=&�>%��=�0��t�����$��=rʻ��T����߼+�ӣ=_-?>��L>dL�;�>*�=��<D���t�O�-��=���>4�>tC�>���=�C��W�*>����]�L�w[�=���P�@�>e��}~��:/��!2�MF>%�\>�0������C ?Ke>�:>m��?Xu?�>�����Ѿ�Н�r�j�?�Q��
�=mD	>&\?�6�:���a��|N�K^Ҿ��>�ӎ>���>��l>�,��&?�}�v=��ᾮb5����>Rm��e
��^�:q��=���i��˺��D?@B��U �=�0~?�I?ڏ?��>qa��p�ؾ@�0>�E���|=e���Zq��L����?�'?gk�>A$���D�<ޫ�v����4>hա�hna���|�.���7=����b>>x�}�ξBI&�L�#���YH?��ܓ���>��^?$q�?�����O��Zli��[���=�%?9��?��l>3{?��M?�I<����,5�%ؚ=��y?�W�?>C�?$�'>�׽=�ҵ�?K�> 	?��?Ѷ�?(ns?�?�/��>��;B� >�ϗ����=j�>s��=ס�=4s?ϓ
?{�
?����S�	�%��|���]��c�<�A�=�j�>�<�>qTr>O��=8pg=��=m�[>�Ǟ>7ď>>�d>���>�H�>�eB��=�~$?L
�<AUf>�9�>�E�=��t>�;$���(�O�|<e�(��(þ7�V��5c����=ƪ\<:�=b�t<�͢>��ÿ���?�H>����*?Ç����>��)>��� �?��=Or>��>�%�>:4=�/>�%>�8߾�>*��.�3�9���R�I�ھJ�S>�ᙾ�G��
	�)��|�?��ν�c����j����?�r�<�ŏ?,н/�e�X�%��R3���>VZ�>��5?贀����U>Wn�>?�k>��}��b���=޾*��?���?�;c>��>R�W?�?�1��3�vZ��u�E(A�Ie�L�`��፿����#�
������_?��x?�xA?Y�<�9z>m��?��%��ӏ��)�>�/�';�Y><=�+�>x)����`�|�Ӿv�þ'7�LHF>�o?%�?JY?SV��n7�\��>^N<?%;;?��?�<?�y_?�:�ȘS?6A�>���>�*?q�C?W�T?�!9?
>�P�=+i:=>=���4?̾/4���Py���*�׻=�-�=���<6�Z<#��=�>n\�<����ļ@tV��]��fcE��v�=�'�>���>��]?JO�>M��>z�7?!��du8�I���y./?U�9=q��������բ�`�{�>
�j?���?�aZ?�Yd>a�A�uC� >V�>�y&>�3\>l�>,wｋ�E��ԇ=aD>�W>ɥ=��M��Ł���	�6���J�<�>���>"|>���q�'>q{��P#z���d>j�Q�[˺���S���G���1�/�v��S�>��K?��?|��=�Z龵+��zHf�r.)?�]<?8OM?��?��=-�۾��9���J��C���>��<���˿���"����:���:��s>�1��J�žn�s>�Ѿ&ž�iO���b�������7����y��!�HΚ�Sr*�lI�=�?�=Ƭ;�(�<�����kSD?��=�_���a�5���%s��B>j��> �K���t�A�2�Pd���f=̇�>�U�=�;��ܾvK����$�>��D?�_?Y�?2S���[s� C�� �������ܼ�?8�>%`?�TB>�8�= 6��8<��+e��H��o�>?�>���u�G������6��cW%����>]�?�->�?ڪR?��
?8c`?�s)?v!?z�>��������A&?(��?��=!�Խ}�T�) 9��F���>��)?x�B�k��>W�?�?�&?�Q?��?=�>ح ��C@����>bY�>d�W�eb���_>k�J?���>O=Y?�ԃ?0�=>�5��ꢾ�թ�"V�=�>j�2?�5#?/�?���>П�>���j��=�(�>c?�2�?A(p?Yi�=oH?�2>h��>�ۘ=��> 6�>�3?$O?gs?�|J?F��>w��<�S��8��;�u�$�o���;`?Q<��x=���=�s�O�����<��;�������ѵ��B��n����;#`�>K�s>����0>��ľ D��Y�@>�>���O���؊��:�$̷=e�>��?���>�N#��ɒ=y��>�E�>���5(?'�?�?y�;��b�|�ھ"�K�?�>g	B?۴�=��l�⁔���u�A�g=�m?�^?9�W�F ����b?� ^?\�I=���þ	�b�����O?��
?��G��>:�~?��q?���>� f�g=n�����Gb���j�|Ͷ=%f�>�T�>�d�+'�>
�7?9M�>��b>��=@�۾9�w��`���?��?��?
��?� *>O�n��5����)����[?��>'־�??Ƒ�̾6La�:J�e�Ӿ#�޾��۾OPž���`��JB���C���=�f?��~?;�^?�Fb?�c
���q�K�M���z9�p:���8� eI�}���D7�ܙo�<����unž�Z�=��{�:��2�?�=#?�����>獵�p�3�ξ�h>O�����W|�=QⒽV^=�W�<h�y��m@��{Ǿ� ?F��>{��>�1?U[Z��7G���8��;�vh�S�+>|Z�>�=�>�q�>i��<�	8������ȾES+6�eރ>�v?q:?�^f?S���ݣ>�P<��r�}�P<T����	>d�>h��>9�U����I$;��uZ�ׁ��y��}s���$��Q�<��?���=&�w>��?��>~���о���n�����?W�v?���>$\>��=��J���>��w?$Z�>L��>�����L!�^�������>e�>���>Ӆ> �RbW�e��J���D^>���=>�n?2w��j�];t>w�Y?���(�J�&~�>�kW����g��;�7���Q>7D�>�_�=��>A���Xz���q�����tp(?��?������(�̯�>y$?���>(ң>��?V۝>��ƾO�;�8?�4`?�K?�??u��>�=���FW���"��S2=�)�>=P>Jv=�C�=u��lI]��#�O =} �=�ܼ����Q� <�9j�B9I<�?�<�)>%I׿��A��@þ���<!Ծ�1��\���6����y�?��Uɾ^"��Kz�4^���O�аw��c�����9Վ�%(�?/��? �R�ȃ�rғ�2���"�dr>���I��Wk��X��:[c������`���"���J���r�0 |�L�'?�����ǿ񰡿�:ܾ(! ?�A ?3�y?��8�"���8�� >�B�<?-����뾮����ο?�����^?���>���/��h��>ͥ�>�X>�Hq>����螾�1�<��?,�-?��>��r�-�ɿa����¤<���?0�@�rA?��(�OL쾝�S=l��>��	?�?>`0�2P�����|�>��?���?��J=Y�W����<�e?Ԋ<��F����,��=>�=�:=���״J>?�>_���?���۽��3>0҅>��!�B�)e^��(�<�]>��ս3d��zۄ?�t\��.f�υ/�]��C:>��T?^O�>��=V�,?rH��sϿ!�\��`?4�?I��?E)?�d��6�>��ܾ��M?�S6?�>C\&���t�(3�=�༦;����㾐V����=\x�>M~>,�C��kOO��r���=�9�ƿ��$���=̺�#Z�)"��O���,T� ����n�,���i=3C�=&�Q>�`�>�W>�HZ>�RW?�k?xK�>��>c佶|��^ξ�/r��ܧ��i��E���ߣ���Y�߾5o	��������ɾ�&=�H%�=R�r���� ��b�B�F���.?`9$>O�ʾ\�M��&/<DVʾ2����l��FT���C̾�1��8n�Gȟ?3B?煿g�V�: �c���m��ٖW?�g�L��Q���g9�=2Q����=}�>���=����.3��S��u0?
U?�~���`��*#*>w� � �=�+?��?�/Z<�*�>,H%?��*��D�O^[>]�3>qܣ>m��>g1	>J��_O۽��?�T?���k����ِ>fm��ܗz��3a=�$> 95�J��X�[>U�<� �U�]N����<(W?V��>V�)�	�A`��J_��I==w�x?�?"0�>�|k?��B?��<)o����S����jw=a�W?�#i? �>
�����ϾW�����5?�e?��N>�gh���龮�.�XU�%?v�n?�[?�H���p}�'�����Mi6?*`�?�=e�T�ÿ��J��U�>Z�?y9(?�$p�RJ�>��f?�*��P̞��¿�᥾���?d�@���?�a�={�*=�e>È�>���>�&����i��X���D>�?X(���3S��v�g���؄?��f?���>|�4��ž�	'>ވ�"I�?Y�?8I�4�=/!��i�S4�����xV���j��1ν��F�B�s������t3��Y'=[�T>m!@��U��г>t�����ٿ�˿q\{�V ־����>��>�x�=m]���i��H���J�LN_��S���M�>��>ɔ� ����{�'s;�.���>J2�P�>��S�.��D���Lc5<%ޒ>��>���>���B޽�}ƙ?�i���BοJ���
��H�X?j�?q�?,e?Km9<�v��{����(G?=�s?�Z?��$��]�$�7�!�j?�_��mU`��4�sHE��U>�"3?�B�>O�-�o�|=�>q��>�f>�#/�v�Ŀ�ٶ�4���T��?��?�o���>o��?ps+?�i�8���[����*�՞+��<A?�2>	���D�!�E0=�[Ғ���
?H~0?*{�].�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?Q�>�$�?o��=F�>�U�=?�� \=��!>�@�=�)A��|?��M?2R�>Ę�=��8�DO/��cF�RbR������C����>��a?ȔL?y�`>!��� E0�Ե ���̽��2���7
?��Q.�֧ݽA[6> >>O>�{D��Ӿ�?Rp�F�ؿ�i���p'��54?���>J�?I����t�!���;_?Fz�>7��+���%���A�h��?�G�?Y�?׻׾�W̼�>��>J�>��Խ���������7>2�B?���D����o���>���?�@�ծ?Qi�u�?H���מ��q{�M&��F�zp�> ]m?�-'����=�?��d�>,H�����]�v���>��?)��?��>g��?i��!s��P>�H�=��? �$?���=�cL��&(>b�?S���Mw�B&X�I h?�@/?@��k?4䓿J|ӿ3̖�G����ﾊ��=M��=!��=f�߽��>�x��ٖ��>q�o>£�>]Jr>��I>��\>�g;>7�>H-��h��5И�i(��ۺS��
�)� �SUS�����^��k6���%y��f���nI���ͽ�t���	�̱�����T*>�"P?�kC?>?]D�>��Խ�:j>q���p>e���5>�\�>[�,?��A?k�,?෎��H���oM�k�m��s����p�>
�>	��=��?zG�>���>���l�>��>Ժ�>�&�=1��=�E�=M�<14r>�l�>ߔ�>���>�C<>��>Fϴ��1��k�h��
w�s̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�4`>�+ �~l���)��%Q>wl?QQf>�%u>4s3��S8���P��Ͱ�]�{>:�5?2��9���u���H�+?ݾ�KM>b��>��F��q������=�6+i�H{=n:?"y?������}�u�����8R>�\>0&=hs�=�L>RFd���ǽ�H�,�-=o�=��^>G�	?W���>
0&>�\���`�=H�d>�C�>�� =E�-?&@5?fm=���~��S����=�W#�>���>>2M�=��d���4=���>d��>���(��m=�3n��g�>&����7����Д<J�ý�l�<��=�f���I��Fq=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾM��>�N�����.a���xo����K��>��J?�����L�q8� ��>��>]��g����zɿ�v��:�>Sw�?���?�s�4���HA8��P�>�?��n?J��>"��X�P����>FR7?J�`?#;�>7��즎��j4?��?aw?�s>㹜?gsK?�F=9��H��}{���c�����=bԳ�z�߽k��/�B��Ĥ�ŵ��1�r�o�>���=?V�ȟ�>���Q$ž�T>!��훾�i��Œ>'O�>���>�v?���>�N�>�K�>�5�LE�����,���{�K?���?���2n�xO�<���=��^��&?�I4?Fe[�h�Ͼ�ը>�\?n?�[?�c�>1��E>��:迿!~����<~�K>4�>�H�>�$���FK>��Ծ�4D�gp�>�ϗ>#����?ھ�,���R��OB�>�e!?���>wҮ=�� ?�#?��j>�#�>C_E�#7���E���>��>,>?O�~?��?�ӹ�eY3�t	���塿9�[��,N>P�x?�S?3Օ>8��������D��OI������?�og?J归 ?l/�?Y�??�A?gf>����ؾ=������>��!?h��^A��J&���n�?Z
?G�>�a���zֽ�Dмg������8�?��[?0J&?|B���`��þ"�<B�#�Y��<�R���>�>.��a��=A�>g%�=6�l��5�X4l<��=0J�>ɪ�=�7�Zč���O?ٱ�K�ؾϖ�=~3�������>��?�,����?&�>$���1���"���&�6>!�?l��?�?3;�&_��j�>O��?4�?>O*#?w��<�ľs�v����N�j��
���f�?���=�.J�����js��b����OO����+��>@8�>o�
?�  ?RWS>8�>��o'���������^�����8��.����=ٟ��L!��[
��y¾�$|�B�>U��D��>��
?d�c>#'y>LS�>���_Ȋ>VT>JK~>Qԧ>��W>FB4>ұ>��<�Iѽ�KR?2���;'�1������3B?rd?1�>qi�������t�?���?Is�?�=v>�~h��,+�Hn?�>�>��Hq
?�S:=�L�f/�<�U��μ��2���ת�>�G׽� :�rM��mf�Uj
?{/?���̋̾�;׽[g��i>iPn?���>*��i���1	z�Rl�� 8��ث�(���V�Jp&�] F�\����Zx�X���6@�u2P�G�?�M\?��徦���|���7�ۨݾ`X�>O��>VD>���>����S(��M1��(]�z.�#���G:�>�Ȑ?��>�I?�<?�R?��K?���>�h�>�7��OR�>�<٧�>��>B�9?�+.?�0?�? �)?��^>qL ��h��ԥ־}�?�n?>�?��?~l?2��YF��z����C+���{�w��2�=�ȼ<Rͽ�b���\=�uQ>�X?����8�4����k>=�7?���>N��>����(��:��<��>ζ
?�I�>�����|r��a��T�>���?���6�=�)>v��=�����Ӻ�X�=f�����=�"��1v;�%=<d��=v��=j�t�*�z�Ñ�:O��;@e�<�u�>#�?��>�0�>�C���� �����۰=x�X>,S>�5>(Pپj~�����J�g��y>-v�?t�?�If=���=1��=o���$�����5콾1��<)x?�g#?XT?��?��=?b#??�>9+��D��X�����b�?q!,? ��>�����ʾ��ŉ3���?S[?�<a�4���;)��¾��Խ��>�[/�e/~����CD�2ޅ�����~��-��?ܿ�?A�X�6��x�ѿ���[����C?"�>3Y�>y�>W�)�s�g�u%�h1;>֊�>hR?<��>�O?},{?&(\?k�T>�8�(���ꏙ��1��!>�p@? ʁ?�׎?�y?���>��>��)�j�߾���7b�y������U=�r\>�Z�>b�>.�>Q��=5�ɽ"�����C��#�=طa>gP�>x�>`��>F�w>�<�9G?Ֆ�>&���Μ������k�[�`�x}v?<��?�<(?��9=x��%xG�����"��>%��?�5�?�9*?�X�[��=�ռ�v��,�_�S��><T�>�U�>�9M=Yy�=�>���>ڧ�>U�����6��rQ���?%1C?���=�)ſ�n�I�h����Y]<�D���p��Ы�mt]��̒=ѝ�i��Ȧ��W�aϟ�>N��1T��l�������>b%�=��=���=���<�-�f�<P[=��<�w=E�p���<#�`�Zn"�ƺ��W����/<��:=�"$���ʾ�p}?�7I?),?�oC?%�x>)�>8�<�!�>��|��3?'�Y>�OH������9�$#���֔���ؾXm׾�d�n#����	>�)T��J>b�3>���=��<G��=bEt=��=�*i��p=���=�)�=î=lq�=��>�>H�w?V����3��XYP�f�]�9?��>K�=�QȾ�D@?�oB>r$��I׹��%��?@�?��?�C	?@{g�o̟>�s��9҈��є=H	��<�/>7��=�2�3�>�HK>�`��Ӝ�\�����?t�@�>?aJ��b&Ͽ��/>E>�o�=I9G���1�SiW�GY$�#�k���'?�=�`?о䭏>�n�=����˾��=�(K>F+�=8���+�[�f�p=ͼ���@=XB�=
zu>M>'��=
5����>F=���=��Y>�:�頼���'=���=�._>��&>>��>L�?�a0?�Xd?i8�>�n��Ͼ�=���N�>��=�F�>#�=!zB>���>l�7?b�D?>�K?
��>c��=�>��>T�,� �m��i徒ɧ��z�<��?:͆?Ѹ>�\R<X�A�i���e>��-Ž�v?R1?j?T�>�<��ӿ��+��T5�9��<�ם�b� >%E���=��s�����>h��>\  ?�9�>B6�>��>qE�=��>�-�>6�=d�L��- >2�#=&
�>z>7�=49ν{��=c����k�5ͽ��*'=���<��W��#��b�*=u��=�^�>�>0��>y7�=j����1>�����N�p��=�N��,�D��md��\~�56.�\�-��	D>Ο[>yt��*����T�>�)h>O�1>���?A�v?>>�@���о���f�a��qM���=�8>R&J��o9��#b�zmN���Ҿo��>���>�>��l>�,�["?��w=��a5���>�~�� ��.(��9q�2@������Oi�� ԺءD?FF����=�!~?�I?1�?"��>5����ؾ;0>�G����=��)q�j��a�?'?��> ���D����]��L�>u@���9�g⛿�W,��=<ʳ�[D�>-������W(9�A({��3����X��]��,��>ʿX?�
�?����Tw���lE�f�0�ZT�=!�?3w�?w%>&?t?<<��f��� R���=|�_?^�?�%�?�&C>��=)!�����>!	?iɖ?��?�t?u�=�A��>%�;�c>#t��p\�=��>&m�=Y^�=�!?�$
?kZ
?����|	�Vt�S9�ʷ`�� =mɢ=��>4ˈ>�p>,��=�ac=$-�=�[>MÞ>~��>Iod>�)�> ��>��\�����'?#��&g}>,�K?�WA>��W>׾H��=�C�=�a������̤?��w�7��=6�5==W�=�٥��H�>�p��{i�?_|z>�r��}�?�s�%r�V�>V6=$1>��T�>#�>�>�x�>~��>s�5>�}>�b�=2Ѿ��(>5aﾢ]#�f�$��?i���޾��E>g���_���
�{L'� ���ߪ��~���7r��I����7�<��<���?z&�%o�ڬ$���7��0?~,�>�M?C���Orv�� p>Rޞ>�e�>�ݾ=D���抿@վ�?~��?�dc>�>��W?ΐ?Y�1��v2�w{Z���u�nA�He�:�`��荿3�����
�ZG����_?��x?`RA?��<W�y>���?�%�
�J�>N/��7;�S*;=)�>�B��c�a�_�ӾXDþ���1�E>�Do?��?�?GU�Ҕ=�v�>��;?�;?tF�?�?�d?��U�~?�(	?���>�X.?��g?C�g?�?n��=B�q=O�нPb��E��a�������;�i�I*3=,��=��=��{<�l��k:N=��!���t�e�<=��<���;��8=>�,;(��<�޻=�¦>�]?AN�>>7�7?���x8�����R /?y�9=)�������آ�����>`�j?���?_cZ?�Fd>2�A��C��>xg�>�J&>u\>_�>���c=E�i�=4>\T>�˥=�GM�;΁��	�\������<5>4��>3&|>T���z�'>G}���z�2�d>��Q��κ���S�-�G���1���v�zQ�>�K?�?۟�=�Z龢"���Gf��.)?�\<?]JM?��?�=��۾��9�r�J�E�A�>�u�<���꾢�\#����:����:��s>�,���.��h�a>H�
�<�ݾ"�m���I�?	龡v>=iU���H=S<�wԾ�Z{�`��=��>h����*!��*���l���J?O�{=M����U�н�Rc> �>U@�>;�F�H]w�a�?�><��G��=X�>�9>���%I�ˤG�����G�>�E?/�a?�B�?CL$��wi���Y� �s����8���?�@�>��?�
�>��>橤�����\n���5��V�>�>����4H�����:񾺟$�J"d>i�?
5;>6�?�_?�J?##\?z�.?x��>���>�����ž��%?y��?�V�=�_̽��N��q8��D�"t�>��)?|(C���>��?��?��'?R?E�?��	>ɚ�n�?�g@�>�-�>��V�Z3���a>�SK?ܻ�>+�W?�Ѓ?��=>��5�q#���į����=�5">g�2?Ӷ"?�S?�
�>��>������=Ҕ�>"c?�0�?��o?׋�=�?62>��>#�=���>t��>�?fXO?��s?��J?���>���<I?��wC���s�~P�z]�;�
I<
�y=>u��s��8�j�<mf�;�ķ�,�����D�א����;�d�>^�s>����j�0>�ľ{G����@>�)���N��Smz:��v�=�j�>�?	��>=B#���=��>�9�>���,7(?��?;?�;i�b���ھU�K��"�>?
B?�Y�=L�l�y��j�u��g=��m?�^?��W����b?4�]?�f��=���þ��b������O?:�
?Y�G��>p�~?�q?'��>K�e�e:n�0��Db��j�[ж=�q�>X���d�@�>M�7?�N�>�b>�&�=4u۾s�w�q���?c�?�?���?K+*>!�n�$4�y_��4t��t=X?���>����!?�_ͻV�Ѿ2솾󾎾Ɠ澸ѫ�c���.������W�/�$.��_�]�=Ϟ?�Gv?�|s?	^?g<��Wb��m`���}��6U�sc����5B�%A��'B�qm�������i&��g@<?���UG1�)Ʀ?r�?sM�����>�¾#E	� sþ�֗=����ý!�>;�;;Bk~;A�������24������ ?6��>kk�>��!?����Y]V�Q>���,���G}�=���>lj�>�H�>Η��SN'�<���IAھ�j��}ny�
��>�Xp?�s[?&;Z?���  �{�~�]�)��=�Ǹ��{-=�">�C�>(���M �P4*�QTK�Hpr�����䎾{T�1��<o6[?�-�>dd�>�?�?���>���S��Έ>�@I#��k>>��>��U?!h?���>��N�������>V�i?���>Fۭ>���V"��)x��ǫ��	�>�ߧ>e�>�S>-x@�nW^��J�����5��s�=�c?���2�A�~L�>\�Q?4��;,4N���>V\�����	���l�?�� �=t	?� �=�u7> �¾����l{������/)?jq?�ґ��`*��S>)l"?#s�>I<�>R1�?��>~þ�_1:��?3�^?WuJ?NA?���>�=qв���ǽ�]&��"-=�8�>K�Z>X�t=���=X���K\��2�#�D=ڦ�=��м/c����<��^�I<�^=q�3>�տ�H��Ѿ	����ƾv���W���3 ��|����*�ƾJњ��_`���ҽ�#���y��|�d��ꀍ����?��?�5F��u��ꠘ�")~�����>췅����뢾����̎k�5߾�Щ�.d�[�O��t�JSv�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@}A?��(�
��V=���>ΐ	?I�?>�N1��I�����aU�>�;�?��?�nM=$�W�S�	��e?m�<��F�5�ݻ��=�<�=@E=����J>�T�>}��LOA�(<ܽN�4>}م>To"����c�^����<�]>?�ս�8��ׄ?�p\��f�/��V���>��T?�8�>��=�,?/H�wϿd�\�qa?�.�?t��?b�(?;�����>I�ܾ��M?uI6?��>Q`&���t�A1�=�߼Z���a��3V�+�=���>GR>L`,�4���sO��������=���۱���V'����L>	>A?n=ݭ�<EsA��,����p=�m���G�a���*M3>���=]g�=��;>�{>N�>)�M?�j?%��>��>:��=���1;��(<`+��]����@��՝��>����g����
���
�����Y*��=���=5 R�Ԍ��	� �w�b�x�F�F�.?<V$>��ʾ��M�;�/<F?ʾ��������v.���A̾��1��?n��ǟ?vB?xⅿ�V��"�li��%��ęW?p�����ά�a	�=Ŀ��hw=n�>ث�=3�⾐,3��S�z/?ź?���S%��1��=�ṽ���<�/?���>_��;Y��>Ļ?�]o��/4���A>�W:>��>(��>���=�/����ڽ��?�=[?s ��۟��8�>�+��f�C�.y�=5�=>�#���Ӽz>>�3L;}�����8��O�����<�'W?i��>�)�7��j��� ��;<=�x?l?L̟>��k?7�B?�	�<x�����S�����x=a�W?4�h?��>�7��<�Ͼň��&�5?E�e?e�N>b�h��n龧�.�.X��?��n?9h?�;��k`}�������7W6?�V�?�?�ү��C����޾z�>�3?	?��c��I9?�qu?�����M����
��7�?4w@B��?��:>t�����+>up�>��>��������������>�W?X[�Bɞ��]��#�����?���?|(?e�ۻb����F�=5쓾�c�?�?]c����<V��J=j�����ry<�=�5/���.�|
�Tg7�cȾ�e
�e[���]��&��>��@ !ֽo>�>�<������ο����Ͼ�&v�?�Ϩ>�+��	���h���r��H���I��C��?N�>��>ί��G���!�{�_q;�D0����>i���>U�S��'�� ���k5<��>���>긆>r&���罾�ę?Ib���?ο������P�X?�g�?n�?Vq?S�9<��v�̐{��d��-G?��s?HZ?�k%�N>]�C�7�%�j?�_��wU`���4�uHE��U>�"3?�B�>T�-�S�|=�>���>g>�#/�y�Ŀ�ٶ�<���Z��?��?�o���>q��?ts+?�i�8���[����*���+��<A?�2>���H�!�B0=�TҒ�¼
?U~0?{�e.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�%�>��?l�=��>��=<���G>;���"> ��=@�"b?��M?q?�>V��=�9��9/��uF��WR�x�e�C�r��>��a?p�L?�b>j���-�.�e� �R̽�n1�!��@��)��\޽'�5>��>>�r>Q�D�Ӿs�)?�~�d^ؿ�'��m𤾈%?�R�>�z?$�0��p���N>5;f?�	�>���o+�������w����?o��?��? ����+��5>)ǿ>Q�>�Ч�v�-�\�۾�X>huE?��p�������y����>J��?�_
@�1�?�0u��Y?jb�H6��5�t�N�����v��>�E?s%#��UF>B�?�'>�)e����燁�OR�><޳?���?|1�>B�j?u���@�xI>�u�>�-a??�>��k��T���>I��>$��_Q�����\v?J|@��	@�m?���5]п�c����P2���V >A/�> 3>�q��Nx>���=߸;���=hZ>�Ѳ>ܘ�>.�Q>#>4d >�~�=�����M%��h��pލ�qI!�������
�=TʾV_�^k�񈳾�ޫ�3���ٽ�4�r�	����R����>�^?�zV?���?�c-?�ǝ�ja�>Ux
�d�4>}�y�$�
<��>�M?Vh?V�1?���=�ɾ�qn��nK�吀��M>��]�>���=�A�>�>�ĭ>9�=�A>�O*>�N">�(>+�»���;j33>e�>�0�>���>�e�>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?m�f>�u>��3��f8���P�]w���O|>^56?�趾�c9���u�'�H��jݾ�.M>ߺ�>S�C�d��������vi���{=�t:?L�?�`��ڰ�W�u��S���bR>�G\>L�=]Z�=�mM>Sec�V�ƽ��G��}.=��=}�^>]�?��'>vf>��>�촾0&3�.D�>��>�8>��?ע?���~�s���ɾ�yK���?>W��>��>r4�=�pU��c>v��>d�>���}�o�e[��Kq�>�pf�la����ǽ n	>�a��`�=Rn�;�YH� ���~Ӂ=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�5�>��^�[ԑ�:؁��Ї��;)��a?��N?�����»�?n�	?�^��0��V�Ϳ��f�gP�>6��?LG�?\%t�������J��n>���?��?R  ?ǭ"�`ݚ����>�S?սO?V��>E*�8���]?�ò?�Y{?�1�>�?y��?r>������!���Ah�ubS>�8���ah�.�"������$�#��J���j���Q��=ė�:΅�>K�;�𾡽�>�=UZ��ݼd��Dm>��.>�~�=0��>
?GM?��6>��߽�-z��j�w�F���K?ǳ�?Y���+n�"��<T��=��^��?YK4?��[��Ͼ��>�\?l?�[?�b�>g���=���俿�y��fҖ<9�K>E,�>�L�>�㈽�HK>�Ծ�'D��n�>Ǘ>����>ھ�/��à���F�>wc!?*��>�Ȯ=�w ?#�#?�j>�>@uE��l��J�E�u�>lJ�>u3?��~?��?����
B3��#��F����[��N>�!y?��?ĕ>>����v����j���E�>h��Ղ?7g?!�hY?��?��??jfA?��d>�O�<׾𨽿E�>��!?����A�od&�Fl�Uu?6??�>q���b׽~bԼF�~����?s�[?�@&?�]���`���¾"�<K��=^��<ãK�@>��>�r��h�=׷>"B�=3m���5�Q�b<�4�=癒>�.�=�B7����a\F?�Ӵ<�P��0��=�3���S���>#?^W�Xq1?�BK������T��/U��!Yh=}�?��?&��?�|�c�V��{�>�y�?`M>-��>���v��ƺ˽:�C����ՙ��>0��>�q=���p���禿�qr���R����>:�><�?Q��>�zK>�k�>;햾]�%�k��f�z$_�G����8�h@.����'ݟ���$������i�s����>g�����>Ɣ
?�8c>6�q>��>��
�I�>B�P>�{�>�Y�>2�S>��4>���=�]�;/�ͽ�KR?����!�'��������f3B?�qd?T1�>ui�<��������?���?Ss�?=v>	h��,+��n?�>�>H��Wq
?}T:=
9��:�<V��x��03�� �2��>E׽� :��M�Cnf�vj
?�/?�����̾�;׽蝢�R˱=)�~?�.?� ��6x��6}���Z�Z�Q�:�S1��D�r������P��Z��}�{�]ц��;�4}�� .?=m�?��߾��̾����/����U�>ƥ�>���>"��>���=r��!FM���v�v�3��(���Z?߭�?E΍>�(L?��=?;�Q?-;Q?ص�>g�>�������>�㛻4�>�4�>��:?C�0?h\2?��?H�!?�G>p ���Y��_KӾ��?��?��?��?ִ?��#�߽��y�HG����z������=5��<2�Ƚ*�i�-͒=�T>�X?L��4�8�A���{k>L�7?�>���>���r-��i	�<�>V�
?�E�> �Z}r�Rb�
W�>Q��?~ ��=,�)>s��=������Һ�Z�=P���-�=h&��7�;��a<���=���=LWt�Ye���+�:L��;�o�<I?y?�e�>q`b>�W���=ݾe��=@>�p`>y�N>8*>�R���/����R]�I��>@��?3@�?��<��=$�=?���섾�Q���¿���f=�4�>#m%?LR?u�?��8?�3?�ճ=	��8���On������TW?l!,?��>�����ʾ��܉3�ŝ?\[?�<a�3���;)�Ґ¾��Խű>�[/�`/~����@D���������~��/��?濝?�A�e�6��x�ӿ���[��t�C?�!�>Y�>v�>Z�)��g�q%��1;>��>jR?�ջ>*P?�{?��[?Y>��7��ڬ��j���8ڻ��>~8??:�?e�?�y?���>��>b-�x�⾀���:��
q��Ă�IH=f[>�>���>E�>��=<�Ž"~���9�,��=�)_>���>�Ӧ>O��>Vy>�@�<�F?���>()��b;��V���Ec�����<t?ީ�?7?r-=�T�˸I�����V�>ޭ�?!��?��,?� X�(��=�&ü�t��d�M��a�>_�>��>!2=a��=�S>3޸>~{�>�H��O��Z/���/�1�?��<?���=��ſ@r�ekt�m#���<�g����c�ƙ�?KV���=����z�?��φW�1ើLᒾ* ���͜��,v��1�> ��=N�=L�=�4�</,��w��<��C=��< �=��q���i<��0������l_���K</
R=6�ɻ9x˾��}?�?I?��+?��C?9�y>%@>��3�I��>�ւ�$4?�V>GP��j��ρ;�����>4����ؾi׾ �c��ϟ�0=>��H�M�>� 3>9��=��<���=h)s=�;�=:�L���=���=���=��=���=w�>Y>�6w?N�������4Q�c[�z�:?�8�>|�=��ƾ�@?��>>�2�������b��-?���?�T�?]�?�si��d�>��㎽�q�=t����=2>��=B�2�`��>L�J>���K��}���k4�?��@��??�ዿ��Ͽ(a/>�,o>	��=~�2�J>�߶z���@��Ā�j8?7�����&�>�P���
�S�Y�<d@>L@�=��%�V���=�鑼��=�0=p�s>��k>���=��g�×O>h�w=	gw<��=>��c=�-���ߥ�$.x=���=&�>�">p��>��?�a0?�Vd?N9�>�n�cϾ�>���L�>f�=3D�>W�=�B>��>��7?��D?��K?z�>ⲉ=)�>U�>�,��m��g德���]�<K��?�Ά?Ӹ>I�P<�A�G���g>��Ž�v?�P1?kl?!�>����Կ�W@��n#���>��>|
r<;���W�w>?ְ>��B��xj>��>��>��?,4�>�i>H��b׀>��>�=][	��F=��ɽq9�\&B;>���г�3��=b����U���=gG�=���<���ڨ�d�;(P>�J >V��>��(>>��>a�R=�@���E>$և��zC��ơ=����Q�E�#Hf�٠�e�,���@��V<>�u_>Ia���쎿�m? Of>�:>��?Omi?��=��6�@�˾����Y�y��W�V�=�g1>[^9�%�5�1a��N���о���>:�>3"�>@�m>�,��*?��w=����'5����>������y��WKq�Z/���ꟿ��h�賺�|D?5���_�=�~?��I?�Ϗ?���>^���-�ؾ�70>������
=��LXp��G��<�?��&?��>B�=�D��þ�.��P�>�p:�~R�=휿��+�_�X�@m��W��>�O�ξճ+�)��*��aeL�q@���:�>#�V?�4�?��Q�I���KfO��F!����L�?a�x?�)�>�?��?���^ھ�|��{�(=A�]?z6�?���?c8r>�P�=MD��`�>��
?�Ɩ?�,�?O�s?�@���>^&
:� >S����~�=Y�>"�=��=/?�	?1�
?�~���	���Xn�-�_�ڃ�<s'�=gd�>S|�>&t>���=u�q=T��=Ya>՟>=;�>��d>|�>pr�>b������&?,�=���>;2?�o�>�Y=R:��Sk�<M�I��M?��L+�7���%Ὗ�<����
�P=��̼�%�>��ǿ|3�?��S>����	?HR���A1���S>�WU>��޽��>0�E>$D}>Ol�>"�>�F>�j�>�$(>��Ⱦw�/>B��{8��C��%s�&߾ݬJ>.��5��7���l:���o4���q���t���*'7�:�=�?����T�v�V�$� j��Q�>���>�EO?�s�/#��q>�u�>��{>���j$�����H���<`�?]� @��d>0q�>5�W?Eo?.�3�5�4��AZ���s�F@���d��)`����-������^½�^?�+x?�9A?Ei�<�w>���?��$��z��.�>`2.���:�,�=���>1���\�d��EӾ���1��7zE>�*o?�T�?�
?H�U��� <���>��J?)=?S��?o�<?�I?����f%?��=\_�>@�?/�A?��M?�e$?��S>iQ��}�!��<��c�9��Ʒ��nv�o�=���=8;�=´,�xG����=�I/>�_�=2KU=��=�s=f�1<&u{=���=Ւ�=>�>X? ��>=�\>g�(?|��"�5�@���j)?JI =��t����K�e �@��=HCj?��?�/[?��M>��F��D�|N>��>)>;�]>-E�>u��H^�l`�=">��">���=�����hw�;���⑾^�<[�>L��>a1|>����'>�}���1z�1�d>��Q�ʺ�:�S���G���1���v�4T�>�K?e�?᠙=�[�60��THf��0)?�\<? NM?��?4	�=��۾�9���J��>�z�>�K�<���J����"����:���:1�s>1������vb>y�'\޾�in��I����h4M=e+��	U=q��־����1�=��>������ �����������I?�Bo=1��W�T�5��2�>k՘>���>�;��xt�$m@��A��`]�=���>{�:>Ҟ��,��G�����%�>QOE?�N_?�e�?������r���B�����B��:�ɼ��?7��>q?\B>\m�=�������d�S#G�P)�>���>���0�G�<��=����$�뎊>6?�>W�?�R?��
?��`?�*?1=?�%�>K����ɸ��k%?�:�?�E�=$�νwcP�T%7��F��Y�>i�)?a�D�~$�>�W?.?Hx'?<�Q?]j?h�	>�� ��@@����>9��>�V�f��]>��K?�z�>s�X?���?J^9>M6��¡��x��b��=�� >@2?�$"?��?�u�>�3�>�ޢ�Y�|=��>=�b?؂�?�Ko?|��=à?��/>A�>���=�N�>��>Jk?N?b%r?�SJ?#�>I+�<;��n���ta�3q0����;��;<+�z=�����l�:�1�<'ͧ;�ż������cv<��\���<!h�>��s>ᕾ��1>�ľjP���A>i���P;���̊�!�:���=k��>�?���>�g#�~�=k��>�,�>���(?��?�?l��:Ưb�j�ھ|�K��ٰ>\B?�O�=��l��z����u��Ye=s�m?Yx^?�W�����O�b?��]??h��=��þv�b����f�O?=�
?5�G���>��~?f�q?V��>�e�+:n�*��Db���j�&Ѷ=\r�>KX�S�d��?�>o�7?�N�>.�b>(%�=iu۾�w��q��h?��?�?���?+*>��n�Y4�߯������X?,Q�>�d��N?k�:�M�̾��u��1�����#겾�������e���"+�os�; ��	�=��>�Z?��W?FQ?Ps�6Sk��B��Xq�P�_���ɾ�����G�Ӿ+�DI�xJx��V�p���T��G
> E��;$8�?+�?[, ?�1���>1���S�=���)>Gp���)�Nj=ն���7<FI^=xiY�e�7�_���4?�~�>?_�>68?��P�SG7�n(�w,;�:�����7>f��>Ҟ�>x��>d�<�%�i����ݾNt��ѾV����=vB~?�O?M6?[_ݼ���2ދ�	sJ�ϗ���뾢��>��m>���><�"����C1�jT��A��CN��炾�8�]n�="�S?���>��p>��?}�>/���>3콙���	�>�?��>?�?O�><�=�����>�l?q��>EӠ>�����!�E�{�h˽�E�>@q�>���>��n>��,�
	\�{b��La����8��{�=�h?Ie���^�Mą>��Q?���:�|F<��>�cz�{�!��]�<(���>�?\߫=�;>��žie�s�{�bf���q)?m�?�P��h'��n�>�"?�>4��>�-�?���>p%ž2�<_�?߱_?�J?��??�9�>cP=��Y�����'��<+=m%�>J[>��u=�;�=��FqW��*��D=�]�=��ļ�Ƿ����;F�����n<���<e�2> ۿ� J��Iؾ������:Q	�|x��H���ԑ��
��˵��͚���x������4�-IU��Qb�fC���*i����?8(�?}瓾~������/&��*<��H�>�r�r�y��¬��P�8����޾�ƫ�v�!��P�L�i�s�c�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@0�A?	�(���쾌�X=���>D�	?�!@>f[1��"�J��D�>�>�?� �?�bO=�W�+
�&ae?��<��F�lԻ/[�=��=(,=����~J>A�>�s���@��۽J�4>Յ>0�"���1�^�VL�<�]>jս}���ڄ?�\�91f�S�/��P���^>�T?��>N�=��,?�9H��~Ͽ�\�%�`?��? ��?�)?����!�>�ܾ��M?Y6?���>�M&���t���=w޼�e��+��@V����=v�>��>ׄ,�w��O�
����=�� ��iÿ�� ����Qa�<̾�;.6��a�սpሽ&�y�g���mAw��- ��>=@��=�R>��>z�P>D�X>�S?��m?�޽>I�>�˽0����ʾ蘰�W�T;������� ���a�޾u$�������"��[ =��"�=�#R�����I� ���b�{�F���.?��$>�ʾ�M��f*<[wʾCȪ�ֆ�̥�̾r�1��n����?=B?���V�����Q�:W���W?@S�Y��מּy��=���b?=\�>���=3��d/3�6_S��b0? M?�p��#`���*>�� �<�=d�+?Ώ?OY<��>�7%?5&+�=s�[>��3>2�>j��>�	>���l�ڽ��?P�T?ٷ���
Ӑ>�m��!�z���`=t'>*5���漬�[>��<	���Y��Ӑ����<�W?���>�)�h ��`���t�͠<=��x?��?��>hok?��B?,*�<Nj����S���
x=�W?�i?Ч>
ŀ���Ͼ$h���5?�e?��N>ֈh������.�T��?t�n?�X?+��By}�g��"���t6?>�?ӥ������� �\�վjt[���$?���>��h��H?��e?����e���	����tШ?<N�?���?j2>�V�=~�#>�`�>t<�>O�=���N��"cҾt�>��	?�j�I�؛�T���-�S?�>�?a�>kf��\ٽ1�=����y?�?��?�s����m<�����k�����9��<��=""�T#�"��{8��ƾ��
��������>�R@���>��7��	�U"Ͽ����bо��p���?�[�>�ƽ�@���j�	Zu���G�{I�l����K�>k�>���������{��p;��:��R�>��A
�>��S��'�������e5<1�>@��>���>'(���罾\ę?�`��?οz��������X?�g�?gm�?/p?/�9<��v���{��� .G?�s?EZ?`%��@]�Z�7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?���>¶�?�- >���>���=�����Wu��Z�={�=*�m�Ő?UM?%�>��=�m*���3�0[K���X����)?�~�>2�_?!�O?�qg>�&���R/�} #������?��S��D'�s	��0�-'>9�G>�h>��*�/���?Qp�9�ؿ�i��Op'��54?F��>�?%��u�t�t���;_?Az�>�6� ,���%��oB�`��?�G�?D�?��׾�S̼�>H�>�I�>,�Խ����b�����7>:�B?X��D��r�o���>���?	�@�ծ?fi�$^�>6��XF����~���.�6�I�ɢ>M�b?y�-����>g?9��=�ep����D���9�>�^�?���?ܚ�>'�?��w�_N_�~�a����>��i?�??���V��
|p>3@9?�u9������wg?b@b
@��|?oZ��pӬ�t��Z��M�a�Ȋ�=d�=#�S>����	�=�H]=pػlۀ�W�>a]�>� m>�P>}9>bb/>6�>�%���M�u���~�w�_�|4�����fL��o���n�������¾\�`��z��K�6�M��7�CƋ��g�<=�F?�L=?�]?�?$>�<Rf�<���s�>�D���&u>PI�>��G?d"^?N6?M����XxX������ �c�c����>g>���>0��>=�>��<nj>��%>U\�=$�=�Nu��7k��6�=��?>P��>x��>��>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?�e>C�s>�3�*8���P�,����y>[[6?_ݵ���8��Ru���H��#޾sUK>��>�i9����V�����~�Ai��t�=�1:?ǃ?=���?���t�:P����R>B�\>�6=��=�O>F[���ƽ7�G�'�+=z!�=�_>(��>�l>�6�=G��>�"��&AC���>�.T>D�<>�,9?9j?�t���ڽ����_G���~>��>al}>�"�=z�G��=N��>f>���y�f��� ���U��LZ>Kw���[�Bv[���=��o��K�=͓o=���X�\r�=��~? x���׈����>?���VD?+5?z��=aN<�"�����N긾� �?D�@�o�?�{	�w�V���?�*�?KJ��6��=C<�>	�>��;5L���?��Žp����t	��#��B�?���?�}0�X����l��8>�V%?�Ӿh�>�x��Z�������u�'�#=n��>�8H?�V����O�v>��v
?�?�^�橤���ȿ |v����>M�?���?p�m��A���@�_��>9��?�gY?�oi>�g۾R`Z�⋌>ػ@?�R?��>�9�4�'���?߶?į�?jX �f@�?ӯS?�ږ��B�;E迾�樿5F����>94���'>,k�=�����V�����{�4�_����>�;F=`	?%l=٬پ�AG>|#ս�*���&�G�M>/�G>~��>ȣ?�ɿ>�C�>��>�:�� 쁾P��!����K?ű�?�� /n�%��<��=^�^��!?�J4?�J]���Ͼaި>l�\?À?�[?�a�>{���<���忿�|�����<#�K>B1�> G�>�
���HK>[�Ծ�0D��t�> Η>�S��8ھ7'��Gɤ��C�>�e!?^��>��=ڙ ?��#?��j>�(�>BaE��9��X�E����>٢�>�H?�~?��?�Թ��Z3�����桿��[�o;N>��x?V?uʕ>a���񃝿YkE�9BI�@���^��?�tg?pS�0?<2�?�??`�A?})f>܇�*ؾu�����>��!?l0��A�s<&��`�av?f)?���>M����Iս�aټ��������?��[?*O&?	j�a�$�¾���<&$���W�=C�;�A��>۹>_�����=n�>f�=�m���6�Pg<���=L��>l�=mG7�������?�h���?��+5�1b�*�B�k�>q��>dҾn#X?�Ⱦ�����1��谝�qN���?�/�?��?{�0c�05?O�?��>"��>����_/����=��]��f����T>c�>J>������A��ak�������Q��r�>E�>Ú�>��>�Y>���>݄�������t"	�ІZ�����1�}T2�|4������I�},=�����>Y����n�>n� ?Pp>�&>���>��<y�|>�`>���>l^�>�$n>���=F�`=�)ѽ�q�<S?:¾�l&�޾�7��uY@?r�d?���>��>����M���b!?���?��?ǂ�>�g�&�*���?�A�>�ev��!?��={Q;C8�<�䵾���J�����΁�>��ҽ~98�~K�0�g��`??]���ɾI~нN��,t=��?`�(?ܩ)�RKQ�v�o�S�W��oR�2�c�i�j¡�:�$�O\p�fڏ��-���� �(���2=-**?�3�?�J��}�����j��>���d>���> L�>q �>�zI>�9	�k1��g]��'�����k�>Fl{?���>t�H?��;?��O?ʢL??H�>���> ���	i�>[�Z:u�>G��>M:?=�.?{�0?�?��)?�a>y������yO׾�?/[?��?�+?ss?C���y[��[��.^m�]z��b~�G��=��<m'Խ��m��-U=�HR>�J?M�[�8�����yk>��7?�G�>���>����,����<
]�>��
?ؖ�>m���[r��p���>���?����=*>��=N]��D�����=�(ż�ڐ=�=���'<��&<d��=u��=�ꆻb!�8�p�:�;J�<�o�>��?^�>���>ף�������5��=`�X>zAL>�S>�߾b���5�����h��}y>�܎?=j�?�%=���=D&�=,o��;���,���ݺ�Ƭ�<�� ?dD&?��Q?M�?>?�#?��>j�Oϒ��M���H���)?h!,?�>�����ʾ��щ3�ĝ?y[?�<a����;)��¾��Խ��>�[/�Z/~����,D��􅻻��O��/��?꿝?|A�L�6��x�ڿ���[��v�C?�!�>&Y�>��>;�)�}�g�o%��1;>�>bR?���>2�P?$�z?��Y?Y�V>1�6��������|�0�~�>0@?���?K��?7Wx?�r�>�A>��/�E�᾽����3�́��hʁ�{�m=��Y>'~�>J&�>�~�>���=	�ѽ%֭���=����=)�g>�"�>E��>���>��{>�ڻ<8�G?���>0V�����������1=��u?o��?�+?�#=f��]�E��H���;�>Xn�?J��?V0*?J�S����=�jּ�ܶ�Y�q��&�>�ڹ>�-�>h��=$�F=�K>��>���>*'��]��k8�oM���?�F?a��=<W����_��j+���������xu��
���f<���=�B��mn��>ݾ��.ʾ��(���~�np���uz�&G�>^>?�=�?�=�\�<��(=�t�=Sם�}��<�=��j��}Y=����8^=E��˕E=�ѳ=��I��=Ŝ˾Pc}?#I?�s+?G�C?5�y>��>�Z3����>+J���)?��U>�R�nn���;��W���ܔ�3�ؾ�t׾|�c�����_5>��I�'�>#b3>��=2+�<���=��q=� �=\=L���=1��=ʥ�=��=���=��>�d>�>w?5�������G/Q�5��[�:?�K�>Rc�=Q�ƾx8@?�D?> 1��鎹�5q�a?��?CP�?��?=i��k�>-�J����o�==I����1>^�=��2�?޹>��J>��V�������?"�@��??=؋�%�Ͽ��/>��j=�?�<��#��.%��񓾁��Ľ��h�,?y��Kn���7<>��������2��߰�>��->������I���;=�4�;/�=6�=ӳ�>��M>��=F'���F>��z���&>:�c>;��='��<.�����ζ�=�=�8>���>e�?�%0?�d?��>ehm��'ξ�+��N�>�O�=�|�>�ˊ=�SD>�{�>�K8?L9D?IK?���>���=z�>�
�>s�,���l�!���E��t�<a`�?�Æ?�ɸ>�iH<�@�A���/>��SŽS?S1?.y?M�>�M����I&��.��왽jw8A�*=sKr�*�T�������^��=�O�>���>�>�y>.�9>�N>;�>t�>r��</�=�i����<{����=�ܐ�n��<)ļv܃��$4��,��b���z�;<�;��\<?s�;��=�[�>��>�s�>�E�=-窾'�>R&����C��h�=$Z��k�A�c���{��L0���-���I> O>�n�r��^ ?`�Y>�C>���?��o?E>��۳Ѿ,D��K2k�oQ�1)>�>eQ>�e�=�	d�^/Q��������>#ߎ>)�> �l>�,�#?��w="��a5� �>�|������)��9q�@������!i���Һ��D?uF��՟�=&"~?ذI?+�?���>e��g�ؾ�:0>=H��N�=��(q�of����?�'?O��>s��D�������g��>;]���p��[��/�5$�=�����>�J˾�W־W������y4����G�jrR�޷�>a;I?���?�]Ͼ̗������*I�J<b�ף?�l�?��=yU�>��?Ht�9b��v���q�a]?���?9��?��'=�� >ybؽi�>σ?!Q�?�%�?'�s?A��f�>��]����=�2�=>�f3> ��=�Q�=�%?��
?7�?.�J�b�����8cվ8]Q���<��=@��>���>�>��=��t=���=��K>]>���>*�b>��>n�>M�������&?AN�=�]�>��1?�Ё>��`=�ऽv�<ԩP���>�1�+�O����zὊW�<ꅻ�xU=�ݼ���>L�ƿ���?�V>47�ĵ?���x;�U>m�V>X�޽���>W�E>9~>꾭>�ʣ>ĥ>>�>&)>"vﾴ�>��������D���X������b>�&������[������&6�����1��Pi���}��88���@=��y?��P��Mp�|/��0���!�>���>z*<?����_��j�=k��>�s>D��Le���ZUѾH��?�s�?�b>{��>ؓW?/R?Rj2�&�2�oIZ��Au���@��d��`�Ӎ�ŧ��o�
������_?A�x?�?A?�͑<��y>я�?p�%��܏��>�.���:�`�8=���>�����X`�u:Ӿlľ�����F>upo?�'�?�?�fU�zQ>i�=O�%?�P;?\'�?^�D?�'?Oh���@.?�xZ�S>(#J?q�j?�bp?��T?��¼e�L����ޯ�=��=ޱ����B��aw=_T<m� <��V>�='���;�o��W޽(ă='5U<to�=ͳ�<�9�=e��<h�8>lC�;(�>\�Z?�"�>�X�>?�4?����8������9/?��.=�;���:��7����򾟆�=�<j?�}�?:PX?w`>�@�?Z9���>B��>++>�Z>�>�N6?�F�o=d^>Dd>��=}K����)�
�F
�����<�">���>�}>!�����->�����z�>�e>��R�p⺾3,R�|�G�U�1�a�t���>XK?3?4~�=���9����h�W&'?w�;?eM?�|?�c�=�vھ�*9���K������> |<����9��n����;���$:�Dr>9r���.��h�a>H�
�<�ݾ"�m���I�?	龡v>=iU���H=S<�wԾ�Z{�`��=��>h����*!��*���l���J?O�{=M����U�н�Rc> �>U@�>;�F�H]w�a�?�><��G��=X�>�9>���%I�ˤG�����G�>�E?/�a?�B�?CL$��wi���Y� �s����8���?�@�>��?�
�>��>橤�����\n���5��V�>�>����4H�����:񾺟$�J"d>i�?
5;>6�?�_?�J?##\?z�.?x��>���>�����ž��%?y��?�V�=�_̽��N��q8��D�"t�>��)?|(C���>��?��?��'?R?E�?��	>ɚ�n�?�g@�>�-�>��V�Z3���a>�SK?ܻ�>+�W?�Ѓ?��=>��5�q#���į����=�5">g�2?Ӷ"?�S?�
�>��>������=Ҕ�>"c?�0�?��o?׋�=�?62>��>#�=���>t��>�?fXO?��s?��J?���>���<I?��wC���s�~P�z]�;�
I<
�y=>u��s��8�j�<mf�;�ķ�,�����D�א����;�d�>^�s>����j�0>�ľ{G����@>�)���N��Smz:��v�=�j�>�?	��>=B#���=��>�9�>���,7(?��?;?�;i�b���ھU�K��"�>?
B?�Y�=L�l�y��j�u��g=��m?�^?��W����b?4�]?�f��=���þ��b������O?:�
?Y�G��>p�~?�q?'��>K�e�e:n�0��Db��j�[ж=�q�>X���d�@�>M�7?�N�>�b>�&�=4u۾s�w�q���?c�?�?���?K+*>!�n�$4�y_��4t��t=X?���>����!?�_ͻV�Ѿ2솾󾎾Ɠ澸ѫ�c���.������W�/�$.��_�]�=Ϟ?�Gv?�|s?	^?g<��Wb��m`���}��6U�sc����5B�%A��'B�qm�������i&��g@<?���UG1�)Ʀ?r�?sM�����>�¾#E	� sþ�֗=����ý!�>;�;;Bk~;A�������24������ ?6��>kk�>��!?����Y]V�Q>���,���G}�=���>lj�>�H�>Η��SN'�<���IAھ�j��}ny�
��>�Xp?�s[?&;Z?���  �{�~�]�)��=�Ǹ��{-=�">�C�>(���M �P4*�QTK�Hpr�����䎾{T�1��<o6[?�-�>dd�>�?�?���>���S��Έ>�@I#��k>>��>��U?!h?���>��N�������>V�i?���>Fۭ>���V"��)x��ǫ��	�>�ߧ>e�>�S>-x@�nW^��J�����5��s�=�c?���2�A�~L�>\�Q?4��;,4N���>V\�����	���l�?�� �=t	?� �=�u7> �¾����l{������/)?jq?�ґ��`*��S>)l"?#s�>I<�>R1�?��>~þ�_1:��?3�^?WuJ?NA?���>�=qв���ǽ�]&��"-=�8�>K�Z>X�t=���=X���K\��2�#�D=ڦ�=��м/c����<��^�I<�^=q�3>�տ�H��Ѿ	����ƾv���W���3 ��|����*�ƾJњ��_`���ҽ�#���y��|�d��ꀍ����?��?�5F��u��ꠘ�")~�����>췅����뢾����̎k�5߾�Щ�.d�[�O��t�JSv�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@}A?��(�
��V=���>ΐ	?I�?>�N1��I�����aU�>�;�?��?�nM=$�W�S�	��e?m�<��F�5�ݻ��=�<�=@E=����J>�T�>}��LOA�(<ܽN�4>}م>To"����c�^����<�]>?�ս�8��ׄ?�p\��f�/��V���>��T?�8�>��=�,?/H�wϿd�\�qa?�.�?t��?b�(?;�����>I�ܾ��M?uI6?��>Q`&���t�A1�=�߼Z���a��3V�+�=���>GR>L`,�4���sO��������=���۱���V'����L>	>A?n=ݭ�<EsA��,����p=�m���G�a���*M3>���=]g�=��;>�{>N�>)�M?�j?%��>��>:��=���1;��(<`+��]����@��՝��>����g����
���
�����Y*��=���=5 R�Ԍ��	� �w�b�x�F�F�.?<V$>��ʾ��M�;�/<F?ʾ��������v.���A̾��1��?n��ǟ?vB?xⅿ�V��"�li��%��ęW?p�����ά�a	�=Ŀ��hw=n�>ث�=3�⾐,3��S�z/?ź?���S%��1��=�ṽ���<�/?���>_��;Y��>Ļ?�]o��/4���A>�W:>��>(��>���=�/����ڽ��?�=[?s ��۟��8�>�+��f�C�.y�=5�=>�#���Ӽz>>�3L;}�����8��O�����<�'W?i��>�)�7��j��� ��;<=�x?l?L̟>��k?7�B?�	�<x�����S�����x=a�W?4�h?��>�7��<�Ͼň��&�5?E�e?e�N>b�h��n龧�.�.X��?��n?9h?�;��k`}�������7W6?�V�?�?�ү��C����޾z�>�3?	?��c��I9?�qu?�����M����
��7�?4w@B��?��:>t�����+>up�>��>��������������>�W?X[�Bɞ��]��#�����?���?|(?e�ۻb����F�=5쓾�c�?�?]c����<V��J=j�����ry<�=�5/���.�|
�Tg7�cȾ�e
�e[���]��&��>��@ !ֽo>�>�<������ο����Ͼ�&v�?�Ϩ>�+��	���h���r��H���I��C��?N�>��>ί��G���!�{�_q;�D0����>i���>U�S��'�� ���k5<��>���>긆>r&���罾�ę?Ib���?ο������P�X?�g�?n�?Vq?S�9<��v�̐{��d��-G?��s?HZ?�k%�N>]�C�7�%�j?�_��wU`���4�uHE��U>�"3?�B�>T�-�S�|=�>���>g>�#/�y�Ŀ�ٶ�<���Z��?��?�o���>q��?ts+?�i�8���[����*���+��<A?�2>���H�!�B0=�TҒ�¼
?U~0?{�e.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�%�>��?l�=��>��=<���G>;���"> ��=@�"b?��M?q?�>V��=�9��9/��uF��WR�x�e�C�r��>��a?p�L?�b>j���-�.�e� �R̽�n1�!��@��)��\޽'�5>��>>�r>Q�D�Ӿs�)?�~�d^ؿ�'��m𤾈%?�R�>�z?$�0��p���N>5;f?�	�>���o+�������w����?o��?��? ����+��5>)ǿ>Q�>�Ч�v�-�\�۾�X>huE?��p�������y����>J��?�_
@�1�?�0u��Y?jb�H6��5�t�N�����v��>�E?s%#��UF>B�?�'>�)e����燁�OR�><޳?���?|1�>B�j?u���@�xI>�u�>�-a??�>��k��T���>I��>$��_Q�����\v?J|@��	@�m?���5]п�c����P2���V >A/�> 3>�q��Nx>���=߸;���=hZ>�Ѳ>ܘ�>.�Q>#>4d >�~�=�����M%��h��pލ�qI!�������
�=TʾV_�^k�񈳾�ޫ�3���ٽ�4�r�	����R����>�^?�zV?���?�c-?�ǝ�ja�>Ux
�d�4>}�y�$�
<��>�M?Vh?V�1?���=�ɾ�qn��nK�吀��M>��]�>���=�A�>�>�ĭ>9�=�A>�O*>�N">�(>+�»���;j33>e�>�0�>���>�e�>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?m�f>�u>��3��f8���P�]w���O|>^56?�趾�c9���u�'�H��jݾ�.M>ߺ�>S�C�d��������vi���{=�t:?L�?�`��ڰ�W�u��S���bR>�G\>L�=]Z�=�mM>Sec�V�ƽ��G��}.=��=}�^>]�?��'>vf>��>�촾0&3�.D�>��>�8>��?ע?���~�s���ɾ�yK���?>W��>��>r4�=�pU��c>v��>d�>���}�o�e[��Kq�>�pf�la����ǽ n	>�a��`�=Rn�;�YH� ���~Ӂ=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�5�>��^�[ԑ�:؁��Ї��;)��a?��N?�����»�?n�	?�^��0��V�Ϳ��f�gP�>6��?LG�?\%t�������J��n>���?��?R  ?ǭ"�`ݚ����>�S?սO?V��>E*�8���]?�ò?�Y{?�1�>�?y��?r>������!���Ah�ubS>�8���ah�.�"������$�#��J���j���Q��=ė�:΅�>K�;�𾡽�>�=UZ��ݼd��Dm>��.>�~�=0��>
?GM?��6>��߽�-z��j�w�F���K?ǳ�?Y���+n�"��<T��=��^��?YK4?��[��Ͼ��>�\?l?�[?�b�>g���=���俿�y��fҖ<9�K>E,�>�L�>�㈽�HK>�Ծ�'D��n�>Ǘ>����>ھ�/��à���F�>wc!?*��>�Ȯ=�w ?#�#?�j>�>@uE��l��J�E�u�>lJ�>u3?��~?��?����
B3��#��F����[��N>�!y?��?ĕ>>����v����j���E�>h��Ղ?7g?!�hY?��?��??jfA?��d>�O�<׾𨽿E�>��!?����A�od&�Fl�Uu?6??�>q���b׽~bԼF�~����?s�[?�@&?�]���`���¾"�<K��=^��<ãK�@>��>�r��h�=׷>"B�=3m���5�Q�b<�4�=癒>�.�=�B7����a\F?�Ӵ<�P��0��=�3���S���>#?^W�Xq1?�BK������T��/U��!Yh=}�?��?&��?�|�c�V��{�>�y�?`M>-��>���v��ƺ˽:�C����ՙ��>0��>�q=���p���禿�qr���R����>:�><�?Q��>�zK>�k�>;햾]�%�k��f�z$_�G����8�h@.����'ݟ���$������i�s����>g�����>Ɣ
?�8c>6�q>��>��
�I�>B�P>�{�>�Y�>2�S>��4>���=�]�;/�ͽ�KR?����!�'��������f3B?�qd?T1�>ui�<��������?���?Ss�?=v>	h��,+��n?�>�>H��Wq
?}T:=
9��:�<V��x��03�� �2��>E׽� :��M�Cnf�vj
?�/?�����̾�;׽蝢�R˱=)�~?�.?� ��6x��6}���Z�Z�Q�:�S1��D�r������P��Z��}�{�]ц��;�4}�� .?=m�?��߾��̾����/����U�>ƥ�>���>"��>���=r��!FM���v�v�3��(���Z?߭�?E΍>�(L?��=?;�Q?-;Q?ص�>g�>�������>�㛻4�>�4�>��:?C�0?h\2?��?H�!?�G>p ���Y��_KӾ��?��?��?��?ִ?��#�߽��y�HG����z������=5��<2�Ƚ*�i�-͒=�T>�X?L��4�8�A���{k>L�7?�>���>���r-��i	�<�>V�
?�E�> �Z}r�Rb�
W�>Q��?~ ��=,�)>s��=������Һ�Z�=P���-�=h&��7�;��a<���=���=LWt�Ye���+�:L��;�o�<I?y?�e�>q`b>�W���=ݾe��=@>�p`>y�N>8*>�R���/����R]�I��>@��?3@�?��<��=$�=?���섾�Q���¿���f=�4�>#m%?LR?u�?��8?�3?�ճ=	��8���On������TW?l!,?��>�����ʾ��܉3�ŝ?\[?�<a�3���;)�Ґ¾��Խű>�[/�`/~����@D���������~��/��?濝?�A�e�6��x�ӿ���[��t�C?�!�>Y�>v�>Z�)��g�q%��1;>��>jR?�ջ>*P?�{?��[?Y>��7��ڬ��j���8ڻ��>~8??:�?e�?�y?���>��>b-�x�⾀���:��
q��Ă�IH=f[>�>���>E�>��=<�Ž"~���9�,��=�)_>���>�Ӧ>O��>Vy>�@�<�F?���>()��b;��V���Ec�����<t?ީ�?7?r-=�T�˸I�����V�>ޭ�?!��?��,?� X�(��=�&ü�t��d�M��a�>_�>��>!2=a��=�S>3޸>~{�>�H��O��Z/���/�1�?��<?���=��ſ@r�ekt�m#���<�g����c�ƙ�?KV���=����z�?��φW�1ើLᒾ* ���͜��,v��1�> ��=N�=L�=�4�</,��w��<��C=��< �=��q���i<��0������l_���K</
R=6�ɻ9x˾��}?�?I?��+?��C?9�y>%@>��3�I��>�ւ�$4?�V>GP��j��ρ;�����>4����ؾi׾ �c��ϟ�0=>��H�M�>� 3>9��=��<���=h)s=�;�=:�L���=���=���=��=���=w�>Y>�6w?N�������4Q�c[�z�:?�8�>|�=��ƾ�@?��>>�2�������b��-?���?�T�?]�?�si��d�>��㎽�q�=t����=2>��=B�2�`��>L�J>���K��}���k4�?��@��??�ዿ��Ͽ(a/>�,o>	��=~�2�J>�߶z���@��Ā�j8?7�����&�>�P���
�S�Y�<d@>L@�=��%�V���=�鑼��=�0=p�s>��k>���=��g�×O>h�w=	gw<��=>��c=�-���ߥ�$.x=���=&�>�">p��>��?�a0?�Vd?N9�>�n�cϾ�>���L�>f�=3D�>W�=�B>��>��7?��D?��K?z�>ⲉ=)�>U�>�,��m��g德���]�<K��?�Ά?Ӹ>I�P<�A�G���g>��Ž�v?�P1?kl?!�>����Կ�W@��n#���>��>|
r<;���W�w>?ְ>��B��xj>��>��>��?,4�>�i>H��b׀>��>�=][	��F=��ɽq9�\&B;>���г�3��=b����U���=gG�=���<���ڨ�d�;(P>�J >V��>��(>>��>a�R=�@���E>$և��zC��ơ=����Q�E�#Hf�٠�e�,���@��V<>�u_>Ia���쎿�m? Of>�:>��?Omi?��=��6�@�˾����Y�y��W�V�=�g1>[^9�%�5�1a��N���о���>:�>3"�>@�m>�,��*?��w=����'5����>������y��WKq�Z/���ꟿ��h�賺�|D?5���_�=�~?��I?�Ϗ?���>^���-�ؾ�70>������
=��LXp��G��<�?��&?��>B�=�D��þ�.��P�>�p:�~R�=휿��+�_�X�@m��W��>�O�ξճ+�)��*��aeL�q@���:�>#�V?�4�?��Q�I���KfO��F!����L�?a�x?�)�>�?��?���^ھ�|��{�(=A�]?z6�?���?c8r>�P�=MD��`�>��
?�Ɩ?�,�?O�s?�@���>^&
:� >S����~�=Y�>"�=��=/?�	?1�
?�~���	���Xn�-�_�ڃ�<s'�=gd�>S|�>&t>���=u�q=T��=Ya>՟>=;�>��d>|�>pr�>b������&?,�=���>;2?�o�>�Y=R:��Sk�<M�I��M?��L+�7���%Ὗ�<����
�P=��̼�%�>��ǿ|3�?��S>����	?HR���A1���S>�WU>��޽��>0�E>$D}>Ol�>"�>�F>�j�>�$(>��Ⱦw�/>B��{8��C��%s�&߾ݬJ>.��5��7���l:���o4���q���t���*'7�:�=�?����T�v�V�$� j��Q�>���>�EO?�s�/#��q>�u�>��{>���j$�����H���<`�?]� @��d>0q�>5�W?Eo?.�3�5�4��AZ���s�F@���d��)`����-������^½�^?�+x?�9A?Ei�<�w>���?��$��z��.�>`2.���:�,�=���>1���\�d��EӾ���1��7zE>�*o?�T�?�
?H�U��� <���>��J?)=?S��?o�<?�I?����f%?��=\_�>@�?/�A?��M?�e$?��S>iQ��}�!��<��c�9��Ʒ��nv�o�=���=8;�=´,�xG����=�I/>�_�=2KU=��=�s=f�1<&u{=���=Ւ�=>�>X? ��>=�\>g�(?|��"�5�@���j)?JI =��t����K�e �@��=HCj?��?�/[?��M>��F��D�|N>��>)>;�]>-E�>u��H^�l`�=">��">���=�����hw�;���⑾^�<[�>L��>a1|>����'>�}���1z�1�d>��Q�ʺ�:�S���G���1���v�4T�>�K?e�?᠙=�[�60��THf��0)?�\<? NM?��?4	�=��۾�9���J��>�z�>�K�<���J����"����:���:1�s>1��) ����c>���!�޾H7n�ۍI��I��N=Le��MS=k�S�־BD����=��
>o0��t� ��K����l�I?gg=XG����U������>�1�>��>�S5��Oy���@�����p��=�:�>3<>��E�G����=�>XTE?MW_?�h�?H���s�n�B����+W���Ǽb�?8}�>�h?�B>�ɭ=˥���	�@�d�HG�w�>#��>���z�G��0�� &����$�9��>�-?֧>|�?��R?5�
??�`?%*?B?�*�> !��I����A&?6��?,�=��Խ��T�v 9�@F����>u�)?�B�㹗>U�?�?��&?��Q?ܵ?��>� ��C@����>wY�>��W��b��c�_>��J?ޚ�>v=Y?�ԃ?n�=>`�5��颾�֩��U�=�>��2?6#?V�?��>ab�>�%��Φx=���>�c?��?d�p?Ð>�.?U&>%��>��=;K�>(��>�L?��K?�p?�*K?<��>��<𿭽���o���Di��3η;�y<�b=�)���E�:��<�<!��;�M��<h���/Ӽ2�:����Q�<#`�>��s>j����0>�ľ�M��n�@>����MN���؊��:�L�=��>��?���>�Y#���=Y��>�K�>���7(?�?�?��$;>�b���ھ��K���>�B?���=��l�����U�u���g=?�m?��^?͏W��'��;�b?�]?�g��=���þ��b���F�O?G�
?��G���>��~?U�q?��>e�e�0:n�%�� Db��j��ж=Qr�>@X�;�d��?�>_�7?�N�>��b>#�=Gu۾��w��q��s?u�?�?���?A+*>��n�N4�.����քP?f��>Y�žR� ?t�Z������7��z<���z�?@��(���s��:���3��G�����)�=^,?�l?�b�?�]?����[���f�����oG������o=/�a"a��J�cl���%�*n���t��Y>�)^�$$J��?�?�On�ch�>m%���M�q�;�Y,>����RS=�b	=v�r�Ķl=A�=�po�ف������&!?u�>k��>�,I?�E_��?�+u1�^N�5���>>)f�>`U�>���>���܇��-��쵺��g�[}=Zs>;as?)N?hJV?U���h!��Qx�#�#����cn��u�>�bO>	]�>7t� �d�P86��@�*|����Q���S��Q
�<�?"B�>ا�>;؛?p�>��:��͐����m��gl>|�>��b?���>@�>��潵�����>��{?l"?�r�>\[��K?��s���h0�=�2?"+�>���>��>=�I��\�Mې��l�����> �e?�풾���{�\>QB?<��>�̻�-�^>c/Y��b˾��I����>���>%�>�Q�=�������?.i�����M)?j/?2䒾�*�Il~>�-"?-��>�N�>�/�?H�>�+þ1��,�?1�^?�:J?�;A?B(�>��=ӥ���/Ƚ��&��,=?q�>N�Z>8Mm=
��=���0�\�ݛ�7D=$h�=�0μ�9��cu<�����tK<��< �3>��ۿtTL�V۾T��>:���������ԻŽ<J�����ѵ�ؓ��N�w�����#��^W���d��ߓk�8u�?��?�����4z��2�� �"��>�7r��ʆ���)�������n�5���7s$��P��
h�=�b�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >ZC�<-����뾭����οA�����^?���>��/��p��>ݥ�>�X>�Hq>����螾z1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@{A?��(�ָ�PkV=���>��	?��?>xG1��;�-��,Y�>u:�?��?(oM=��W���	�|e?��<a�F�@U޻O*�=�,�=��=h����J>�T�>�v�:EA�8jܽ��4>}ԅ>^c"����~^�u��<��]>s�ս�4�����?��=�5͑�	�c��\}�^�U>��J?��>Ʉ��n�d?Ŧz����KM��Ȳ?+�?.��? �$?S��=Q>qꪾiJ?L�?S��>/��. ���n�>i]�< Bl>�� ��q��eΛ;��5?`�F>�-����&�6�oߊ���=�E�kPȿ|�0�v�R�?�:s8���s�1K��ʽU�3��&����C��"ͽ�p�=P>�:E>ih>b�e>��@>�lW?��u?y �>x�[>�q	������7���⟽�^����S������>��̾a��������%�cL%�8��4d��� =���=7R�;����� ���b�ӕF�u�.?�t$>e�ʾ��M�{V-<rpʾ����҄��ޥ��.̾I�1��"n��̟?�A?D����V����J�<���ޮW?�L����鬾i��=v���r�=O$�>?��=���z 3�O~S��s0?�]?�p���P���&*>�� �{5=��+?��?B[<e-�>DO%?M�*�*i��A[>�3>Iգ>f��>�R	>����G۽�?ɅT?*��w����֐> R��Z�z�sa=�>�05��(�+�[>i��<i��V��A���%�<�(W?���>v�)�:�Qs��p����<=��x?#�?p&�>_vk?��B?�<ip��7�S�����w=U�W?g5i?6�>������Ͼ�h����5?`�e?ϜN>t<h���龘�.��N�-(?��n?kX?����ow}���9��8q6?ôt?�>`�0������F\�
^�>��>�>%�@�3 �>��:?��(�hp���/��N75�!��?!2@��?}B�<+�� �L=���>���><[A�3i��e��v���P=G?罙�Y�q�Z� ��r��??x�?��>y惾,��O��=����i[�?��?������h<%��f,l��i���<�~�=�����#����7��ƾ��
�nŜ��������>�R@tz轙#�>�H8��,��@Ͽ���X'о0tq�1�?�Ū>�ʽ����p�j�/u��G�2�H��\���K�>��>����v�����{��r;�.����>�!�4
�>�S�(��I���c?5<��>/��>麆>���T佾hř?
f��Aο����"��9�X?i�?�n�?fm?8a:<��v���{����<-G?��s?/Z?�0%��3]�;�7�$�j?_��iU`��4�tHE��U>�"3?�B�>K�-���|=�>���>g>�#/�w�Ŀ�ٶ�3���W��?��?�o���>n��?qs+?�i�8���[����*�ʷ+��<A?�2>	���J�!�:0=�VҒ���
?J~0?{�t.�g�_?ǣa��mq��.�5Nɽ���>f0���[�Ĳ���e��/�� .|��%�?�n�?hH�?\��ޚ"���$?�ί>�B���Ǿ�9�<J��>��>��L>��T�\ v>[.���;���>Ch�?]��?�\?:���k���1>�}?��>�L�?;��=���>J �=X{���
���">8m�=�$���?X�M?�N�>���=0f?�?�/��D�7Q�Q��o�B��>%�`?
LK?�,t>��V��t-�AZȽ�/���
�U@<��0,�>�۽�6>6�?>i>5?� Ծ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji����>9 	�����3ɖ���.І� ]>�W?�#��>.̲>���ʟ}�A%���r|��;�>���?\��?*��>AZ{?�^����u������>��?��@?w����_4�
��>++?uҾj
��Q?ɾD�w?��@@�m`?�����ؿo��Ɖ��ٺ���>�0=��=�J5�[��=F��q/=7�ټnj�=(�z>!{p>���>�">~0Y>f+w>���T&�&)���ʐ�(A�y&��,�\¾��dOG�I��޾Kn��Y����:��rH�c��"��>�G=.��=~b?RS?��]?��?C�Ҽ-k	>B!��	��n��N�)>���>=�>?1T#?��?XQ�&䐾�@b�l�x������Z���f�>�ۆ>�Q?��>Ǳ�>��>Xhf>e�'>dn!>�BT>��==�T����=�ҕ>T��>�k?�s�>�
<>O�>Rƴ�-*����h���v�M˽���?����ɶJ��,��s�������?�=�`.?Ǘ>����Fп�����H?���� ���+� �>��0?}>W?^�>w۰��;U�>�a���j�e�>� �$Xl��s)�0*Q>b?��>��>��4�9�5���,��w����>��$?�_��aa�ji��
c���Ӿ�0>_��>K{=��$��e������XRn��34;�$C?*%�>��"�`�&��}�h����>��>�M+= BH>�*D>��<�(I����*��=b��=��#>�N?s�,>(�=��>n�5�O��Ĩ> �B>��,>��??��$?V�� ���냾(�.�	�u>�I�>y,�>h�>T�J��t�=�W�>=�a>�P��^o���1���>�/�X> $~�g�`�~=v���u=�$�����=�\�=�� ��z<�m� =�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�w�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?uI>=��?:�x?w��>�w�<�.1�_r��)�X����>Ub�=SL�>�F>�2��a�<��������)�{�j$�ف:>b1�:1k�>����|��/<gA��#��0r�M�>^$a>̣�>6�>��#?p�>#Ô>j=���=�������\�K?���?����2n��S�<H��=�^�v&?KI4?!c[���Ͼ�ը>�\?@?~[?pc�>;��S>��5迿5~��ը�<c�K>4�>TI�>|#��]GK>I�Ծ�5D�Ap�> З>I���;?ھ�,���B��^B�>�e!?ʓ�>�Ү=�� ?��#?%�j>U%�>�]E�G5���E�L��>c��>JF?S�~?u�?/׹�J\3� 	���䡿މ[�jHN>��x?*M?_ȕ>͈��j}��'�A�9�I�&��*��?sg?_"彺�?y.�?0�??��A?�f>l��/ؾ4ۭ�-ـ>+�!?��A��G&�J���z??5��>���WJֽ�ؼ��p����?\?I)&?���({a��þ��<u$�g����;k%P�ut>l�>�燽2=�=�>a,�=l�=�5�|�t<���=���>]#�=��6����=,?j�G��ڃ�v�=��r��wD�0�>bGL>���w�^?l=�N�{�����x���
U�� �?!��?ck�?�����h��$=?��?�?!�> K��4~޾���iPw��|x��v���>,��>��l���1�������KF����Žz�,���?r�>�8�>�V�>�$R>JP�>�y���\&����V��Ymi�����{7��"��������		��[����ʾ��h��}�>��7�>��?�!w>��p>���>�ʼ�ߝ>��k>\~g>�ۦ>��I>�\->+D>S�����KR?����'�Ω�����3B?Hqd?6�>;�h�8���M����?��?�q�?Bv>�}h��,+��o?4�>����n
?�[:=y��1�<�O�����7 ��!��+��>Q׽�:�>M��of�ig
?D.?�獼߈̾ZA׽���8�D=��z?��#?�N0�fUw��@���q��s�G�\�Q�\�,��=�/�vu��荿q���X�����,�U>�x&?�ό?V^$�@~�������
N�E @���t>�П>Q�>���>(RA>�\"��A5�B|�!��J�:���>��~?t`�>��L?�C?�,O?��U?rZ�>۠�>bA��zx�>�N�<wZ�>�}�>o�<?��?]'?�?�q'?{vL>g�罯���h�ھ(�?6�?��?r|�>I'?��i�8J���g;��ֽX�s��â���={�{=�`N�D�*�$��=��>�T?�D�Z58�o���4�p>yD7?6X�>�c�>�:��su���#=��>�r?�ː>}���X�q�0���>��?e-�T�<��'>�W�=�_�>c�o�=���%[�=�i��H���;���=�ݏ=�=���$8gid;x�<�:�<�H?��3?J��>,6�=�����t���u�L�����>Eh���>�+���舿�����g�r	i>���?�Ű?&��>�6>�:>6B
����2B�7�˾��g���&?h4�>h�d?c��?�	?]?N�;������6�������U?(!,?���>�����ʾ�񨿜�3��?Q[?�<a�W���;)�ؑ¾��Խ��>�[/��.~�����D��$������~����?ǿ�?A���6�lx辮����Z���C?2#�>�X�>}�>s�)���g�j%��0;>��>�R?�ܻ>8P?y){?9D[?�V>�8��ӭ�����S`8��">"2@?���?0�?7(x?�R�>f�>�)*����?��� !����bI��X�[=�]>.��>���>m|�>���=#Fǽ�ʰ�~h=�sT�=/Ta>u��>-�>���>��x>b�<>�G?��>9����Q�以�� ���=�޸r?.��?�|)?3|=��$G�����>36�?�z�?�*?Q�L����=!���.����t��\�>ޠ�>���>@��= �X=�>���>��>X�����r�7���T��h?SZF?��=6Sƿ&6r�{�r��C����L<����`�e�aؘ�M$[�Շ�=�Ę�6��z5����Z�O۟�w����;��������z��a�>7�=^��=C��=<�<bּ�	�<�CI=DP�<�
=�<p�K}l<��?��x컷g������ƒB<��I=���l�����s?�DC?�Z,?�R?�m>&^(>7�%K�>�|O�!=?���>+�B=�¾љ4�S���gF���Ǿ��о0�Y�3��V~>�:��� >39>�.�=<�=���=7-�<�}=�Y�<�$=��=��>�"�=jA�=�>>K�'>p�n?(������s凿��]�6�g?9z�>g�=e�@���??OI>���<$���X��b�y?�W@��?��?-�׽�r�>IRc��=t�h��=�L�����>�K��Y�����>�e_>E.	�d����5н���?/�@��?V���h�п\�y=�2>�>��R�01�l�W�ȧ]���L��p ?��:��˾1B�>�'�=�߾QYǾf�6=}6>�6@=>�+��;^��Z�=x�JT=�Y=��>ӚK>���=u���V�=@M:=Ѕ�=d�U>�Sx� ������8=�>�=�_>�>���>�?�0?� _?+d�>��_�2̾^EϾ��>�l�=V��>��=��>��>V�1?KE?��Q?y{�>w�=
��>�6�>/��m�]�ݾ�ء��ʰ<\�?z�?�,�>�d�<��:���V�=���ǽ��?;S4?�n?s�>����
�6�+�j��MP��Sm� ���/��_�g��tE��<���Hc
>Ϊ>B��>�,�>���>6�K>>�(>��>*h>�m��`>[��^<G��g��=��=��ҽ	��C�n���<�֊�Y�����;����W1��֠��x�</��=�U�>�>3�>�6�=a
����2>hӓ�&�L��O�=_>����C��c���}�@Y-���3��8>(�E>'���C8��be?�Y>�?>�X�?,_u?� >����"Ͼ�V���S��Q��d�=s��=�;G� �:���_��.N��z־���>���>ҥ>Y�n>�6+��0=�-==��ݾ�3��8�>ʊ�`������wq�K=��Ц����f��V;�
E?����=�b}?��G?x��?E��>�F���1־&~7>�3�����<+�w��솽��?.%?!C�>j��>�H��t��=�{�>�-T�žb�������K��`��0�ɾ�YF>���Ӵ�ܞ8�Y�����{�L�Z;�����>��^?��?���M���៿ ��<=,P0?6�?�$9>�A?
��>Q犾0'��3��c<�=�.�?�w�?�D�?�==r�=+۞�uq�>*�
?XL�?�Ӑ?r?1�Pm�>�.<M�>�z�t��=��>��=���=d�?F�?��	?�g��m
����꾍0Y�ŏ=��=,�>�Z�>vw>ب=��?=$��=��a>���>�f�>�a>��>,�>����Q��,=?(u<1t>>��8? O�>tO>Og����S�|�=�Kю����Ņ�J1�;�ߣ=pU���-���(��i�>P�ԿL�?�s�>�%'�.�?�F+���ս]�%>�x>����>w��=�3q>�Ā>���>��'>�-�>a�>GӾ�~>A��{d!��,C�2�R���Ѿ{z>ݜ���
&���4y��%CI��n��]g�cj�:.��s<=�wн<H�?O�����k�o�)������?<Z�>:6?�ڌ������>���>mƍ>�J��y���)ȍ�|gᾄ�?6��?G��>3MU>�^[?v��>mȧ�4p����;������N�#�^��AP�:tW��X������}:��`[?y�?"W3?�-�>l�L>�*�?��6���ľꞥ>Z����!9�<�m?�q�y0���+����*@��2�=��Y?;J�?��\?@*��T(>W�߽)Ь>��k?ȷ�?]H?��/?<Kt>�i7?'�d3;?��8?蜀?Y��>���>�aB�q&h�b�}>p�����$��L����6�[�}��H�(w6=�8�=#��%<j%�H�y=T�u����<���=C��<(Ǯ<����h�=��m�d�>��[?��>P\�>��1?bn���5�tS��)�0?�<y��/?��g��8���=�~j?��?�\?�Cx>n.B��N*�s�>�Y�>�>�[>P�>�Ͻ��3���W=Q3>�>���=w�|�߁�[7
�oO��)N=>���>�&�>�K�+�<����tD�����>w��QH�S����o�S���=�Ti�>Ʋf?A�!?ƺ<�"�]P*��~��-c<?U_+?�A?�.�?1>7k۾�#��*�Y��W�>J�#=No�>�ſ�E����B��s^���<���꠾׺a>�����޾\@n���I���,5L=jZ��cO=T=��c־�9�2b�=�
>�r��d� �����䪿6�I?G�g==$��f9V�}���Ș>�ۘ>�/�>��9���s��+@����=��>��;>����&�,G��#�Ň�>�H?��`?ݬ�?_ ���\q���>��뾄(���}�dy?]G�>B ?_�B>�>�=&���*���g�tH�G��>�s�>���GE�������m��+�>[��>.�>03?z2N?5�?4$`?�T,?��?���>�U���Ǿ�A&?D��?��=��ԽI�T�2 9�CF�Z��>��)?~�B�Ϻ�> �?G�?��&?�Q?:�?��>�� �TD@����>�X�>^�W��a��h�_>8�J?i��>�;Y?.ԃ?��=>d�5�i뢾�ʩ�W�=H>��2?X6#?�?���>�<�>�����w�=��>�c?A�?ԇo?C��=�u?-�3>\��>��=���>£�>S*?XN?��s?b�J?�j�>�\�<��������6Wu�;^c��GP;�Wa<y�n=����?�����.�<�@�;�1��ሼ�켚�G��t��/<MN�>ws>�ɕ�9�0>-�ľm[���@>r|���^��D��E�:����=!@�>�?�}�>�#��m�=���>�1�>Y���^(?�?9?-� ;x�b��۾�SK���>l�A?���=��l����u�u��He=;�m?H�^?@~W�t���"�a?t�^?;b�:�X�þX�f�13�gP?��
?��I�H��>��?4�p?���>1	f�Z�n��]��"�b�Żp�6�=g@�>u�`d�}��>��6?_�>%r^>o��=�ܾjv�Ǳ����?ر�?���?�;�?�&*>��n�,�߿������#E?D��>�h�1�? 9��h� �G���A���K��ٰ���AM��(��T������o�p����h����>xWu?x�r?��s?�����x�Óo���a�ǎF�y{�!�о��R��/m�5�Z�"��r�������,�<=6>V�~��B�|��?�<&? E-����>�^��H�D�̾XB>襡����O�=�I��K=�_=i#g��.�绮�
�?rg�>e�>I{=?�j[�d�>�u�1��7����:�0>Oޢ>�Z�>���>6���:1�W�IIȾ����-�˽�Iy>4�g?kJO?�5l?��i�0���u�w��erJ����e>�@]>�=�>�;6�G#���,���J��mx����C��`����<�#?M�p>H�>X��?��>r��dR����k��(����=���> mh?���>x}�>"�
�h))�F��>�b? �>��>�־��8���V�?��=y
�>��? N#?�F�>������q�d͏�:����M�I�=�nz?�W��E��Д>��??�(�=�>ºQ>�&���ؾ��)����u~=�>�9>�ͼ�������`$~���ܾ��&?�v?_Ȓ�oR-�L��>�"?i��>錡>bՂ?a��>j�Ⱦq�3:ˍ?�(`?�RK?�	A?qD�><X ='�ý������0�u�p=Y�>�[>��I=#��=��!�p�]�h��~=�=<����k��0�l;1zż9%X<�=d�?>�xۿ�CK��vپ���A�PD
�\,��}����c���	�
`��_�7x������'�'^V��]c�M��� m�px�?�:�?BW�����%�����������饽>urq���~�����2��m��R��C�S]!�G�O�ki��e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?7�y?��7�"���8�� >eC�<�,����뾬����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾y1�<��?7�-?��>Ďr�1�ɿc���|¤<���?0�@}A?-�(���쾑V=?��>'�	?$�?>�S1��I�����pT�>j<�?���?H}M=g�W��	��e?�|<��F��ݻ��=><�=�F=�����J>fU�>"���SA�l?ܽ�4>1څ>�~"�j���^�g��<��]>��ս�:���e�?.mf�Q〿1����7�����=�wj?w�w>�f7�1Y?a�[�EϿz�&�ӑ?c��?��?A�H?�)ݾ~%d>5¾N�[?�i@?�n�>41�,R�0K>3̾q�>�~"�m�h��ב=��?3�>�.����0��Bo�&���t�<�� ���ǿ�"��!�܎&=#v�;/�:���x��T�I�M茶�?l�w�ս�؎=$��=�.T>�>>�O>0�O>|�U?�4i?��>�[&>=��]�� �Ͼ�q��u����!�@%���?$�~ͤ���>���d	�������Q����=�g�=.8R�{���=� ���b�}�F�~�.?�m$>��ʾ��M�|x*<�nʾRǪ��}��8ϥ�C,̾�1�)n��Ɵ?��A?����V�!���N��m��"�W?�D�x��nӬ���=���=�(�>���=t���3�{S� j0?=\?X���P����)>�O���=7�+?2�?�[<�!�>R%?�+�t�k�Z>D�3>��>��>��	>���<zڽ\v?�oT?!"�2���ː>�A���Qz� Ib=�{>Y5�,���y[>��<�
��(h^�������<�V?/0�>�'�ބ�J��I���4=R�y?A?���>P�l?oFC?�.\<Fy���S�9�r�X=dX?�k?�	>���RBϾ@�����4?D[d?a�M>�t`��f�(�+�7��O?6�n?�4?�XƼ�}�
���o0�R�5?�v?b�^�{����&��'V��b�>~��>
�>�<:��Ƴ>�s>?�\#��4��V���1@4��מ?��@Y��?��J<���ċ=�?�>E�N��RžN߳������l=���>{����Mv�p��Q+��8?w��?N&�>�ւ����D��=#4���E�?���?Oj����c<;��Ul�m��^�<�٩=��"����7���ƾڌ
��_������ˬ�>	U@U罗u�>�9�;"��CϿ�셿�XоG�q�M!?7�>D�̽�룾��j��u��JG��H��(���J�>�>4�������x�{��q;�2��.�>���	�>B�S��&��+��� T5<-�>Ԯ�>丆>("��:潾@ř?�d���?ο�������c�X?�h�?o�?�n?t�9<��v�
�{�if�U.G?y�s?Z?J%�t6]�$�7�#�j?�_��qU`��4�wHE��U>�"3?�B�>O�-��|=�>���>g>�#/�w�Ŀ�ٶ�E���X��?��?�o���>p��?us+?�i�8���[����*���+��<A?�2>���D�!�=0=�`Ғ���
?R~0?6{�h.�9�_?�a���p���-��ƽ�ۡ>߲0�WX\��Q��"���Xe�0��L@y����?t]�?a�?_��
�"�3%?
�>c����+Ǿ;w�<9o�>8�>�2N>��_���u>�
���:��Y	>׮�?�}�?bj?ڕ�������6>��}?�f�>�o�?eP>s��>_��=E��h�7�-0>g�>�x�Ĥ?�kQ?V�>�l�=C�;�*u1��K�t�U�2P��	?��Y�>��X?�E?�`>K��� 鼸 ����c7�tt�U2A�Bp�����E�C>��C>��>��K�R�ھ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji���>)��@��:��O����Y��@L>��L?���V��>���>.�= /q��e���Nn�<j�>. �?4�?o�?��?�%���e��3p�=��>�^�?m/?�0Z=�*�{�B>4�?��NCi�E�����f?=�@�@�V?2�����ѿ䲖��������d��=Y��=���=sz(��q�=>Gb�4gl=�R�=I�a>��>`�q>U>�>[�\>�=�ǂ�;l�t���i����F���.�|t6��-��u��񚣾�H1��Щ�7UԾ�����"��V)�vs��~�F�(aU��9>�*\?ibO?��k?K� ?�x�;E(D>�dʾ���=��P���=>�Ӭ>��G?i�@?�?���þ�d�ұ�������Ir�:k�>��t>�?ܘ?���>����,�>gt>̹�>�7��/">jH׼~d�=�)�>�>��?m��>��;>��>F���&.���Xh��u��8˽��?�R��E�J��+���������8�=�p.?��>����:%п��K
H?�`�����+�,��d>�|0?�XW?M>�հ�j�N�N4>����i���>w��2�k�MN)�~uQ>�a?��L>VW>��5��;�O�D�u2���y>0.?�$��x�m�)w���K�>ؾ-69>Ո�>�����M�,����^��I�^��<k�7?���>��ӽ4ɮ��V�寇��O>"Cz>��\=%��=��[>����HYs��r-�ԨS=�!>�W>�?��3>���=�M�>>���[>^� ��>�}?>">,>ĥ9?'� ?~����<��>�Ddv><^�>σz>f�>�1C��\�=��>�Z>x�\�����m
�r95�&zj>�5/���B��^�`G=���{��=�*n=�g�`�5��|0=�~?���%䈿���d���lD?T+?H �=�F<��"�E ���H��C�?q�@m�?��	�ڢV�8�?�@�?��%��=}�>׫>�ξ#�L�ޱ?�Ž6Ǣ�Ɣ	�<)#�fS�?��?��/�Xʋ�9l�}6>�^%?�ӾPh�>yx��Z�������u�m�#=Q��>�8H?�V����O�c>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?toi>�g۾:`Z����>һ@?�R?�>�9���'���?�޶?֯�?��]>p��?=F|?w.�>0#���"�誠��1W��H�>���~;>�u�>����v�1��ۛ�����4|��<�R�|><��;�U�>�E����V�!>��S�)��q=���>�$>ߔ4>؝�>��?�5�>w�>��C<"Q���~�0�Ǿc�K?���?5���/n�2?�<���=ү^�D&?aH4?��[�^�Ͼ�٨>R�\??�[?�^�>����>��迿}����<��K>�2�>�K�>�	��/JK>X�ԾY4D��o�>�ϗ>^J���8ھ'+��9آ�7D�>�f!?O��>�Ю=��?e*+?�z>H�>��M�����>��1�>!��>�|?���?��?�Ѿ[�;�"����B��;�Z�l}�>0��?!�?^��>|���Ǘ�����4�aQX�y�?U?�`��}�?���?��@?w	*?�T>�tG�N�xF��O=�>t�?(���iB���(�*���	?�Z?{�>|w���-
��%P����0���?
?�
[?�#?��,da�.VӾn�<J ����<'.c�eüI�>�#>��E�$~�=6.>vP�=^bM�u�#�I0=2y�=K��>]�=h�&�����<,?ЧG��ڃ�5�=k�r�:xD���>}IL>:��ӫ^?�k=�7�{����Px���
U�� �?Π�?�j�?�����h�%=?��?�?d �>�K��G}޾A��<Mw�9{x�pv���>���>l�l�����������F����Ž��1�y^�>��>�Y�>4�?;'�>�N�>Lm���Q�u�l���j�a���-<�������T��El��`�;�7���TՈ�!��>+�*�ī�>XC?^�?>XN�>]-�>������>�*>�G>��>"�A>��>"��=�x:=
n*��KR?�����'���辪���g3B?�qd?81�>^i�4������~�?���?Ts�?R=v>�~h��,+�qn?�>�>;��Jq
?�U:=�5�;;�<!V�����w3��Y�$��>5E׽� :��M�Onf�ej
?�/?�����̾G;׽�Y�(�<�6?�$?����mZ���{tk�
??����0�q���h����1|j�#��@u�������t��я�2�/?�˓?��Ǿk�߾Ix��]Q{��QC�k��>S��>��>��>�|=��6�mJ�(�m�|��:`����>=d�?(^�>#aJ?Z<?��R?�O?"��>˃�>맾���>���;sV�>[K�>�^=?"�+?2-?/v?�
'?�Z>Y�p����Ҿ m?�v?&i?�c?��??�z�۬���֒8�S��M��r[���f=X�=��ŽN[�|z�=-�i>tX?Q���8�����"�j>P7?}�>���>)��)���:�<��>�
?oC�>�  �;}r��b��V�>���?���x=��)>R��=������ҺX�=���q�=k(���x;��T<h��=��=�Wu�,􊹸7�:^\�;Do�<��>"�-?�j�>E�k>y�"�$�w���=?t}>GJW>V>�����㓿9���4�]��F>� r?�ɛ?�L>Z>�,`>�z�sK���A
�6Y߾�ـ=#5 ? S?J[?��?�[[?%�?z.�Ğ־ ��f���	w��m?w!,?��>�����ʾ��։3�ڝ?i[?�<a����;)�ݐ¾��Խα>�[/�h/~����=D�u텻���Y��5��?�?GA�V�6��x�ڿ���[��z�C?"�>Y�>��>U�)�~�g�s%��1;>���>kR?��>�7P?=/{?\{[?�FR>�8����T��=�"�۵>�@?���?*ώ?5�x?O��>r�>�.���������򽽄���S=�R[>�>�k�>q-�>���=�Ƚ�����@�S��=�cc>���>�>!��>��v>��<��G?���>�O��V��G򤾪̃�9q=�Y�u?���?,�+?qN=�����E��A���5�>�j�?���?�-*?��S����=�uռ�඾`�q���>JŹ>+�>5ؓ=0G=�v>��>��>6<��Z�fo8�n�M���?�F?B��=��ÿ��q�`w��f��z�<4刾�3`�{���͞X���=A��!!�خ���hZ������t�������a��������>��i=�Q>��=?b�<��޼��<��d=`�<�v=�S��}<�7�8���\��!uV���j<�8`=�|�K ʾ�g}?%9I?�+?�D?-�|>�>��*��_�>Mt���f?�UV>��=�曻��W<�w=������Oؾb�־c�����?�>^�@���>��6>���=��<���=��}=jʑ=�'���#=���=q��=�f�=���=RU>�>[ox?�֌�B?����P�{���:�B?:�>L4�>�G���Y?F��=ZHy�)��}>Ӿ�m?� @(��?��8?ӕ�MF�>�uľ�ý�>�gR��n6>kK�<�1\��KQ>�E>��7�O��J��)��?#��?}�2?�6��	�̿��b#>��=�}S�LV3���E�C�3�m�P�??��4��ᾦ.]>��<=��ܾXZȾ��k=Ⱦ6>1�8=��5�"�c��͒=�Ĩ��b=�!�<� u>��7>�@�=vP�3��=ٕ=��>�g>d�<	�»�':��Db=�-�=l�k>Vz>WS�>��?�F0?��c?&:�>��n�uyϾ@*��7��>��=׹�>٘�=
�>>f��>�.7?�zD?tL?�<�>(ԋ=���>fS�>ek,�+Gm�l���&��w^�<ol�?��?f�>S΀<��A�����=�`"Ƚ�?B1?��?�2�>
F�|���F&���.�<̘��ʤ987,=r�I4U����M�H��j��=���>��>p�>g=y>��9>MTN>K�>�i>��<���=X׍�a"�<����΃=�y��)�<*ǼV����)�E�,�4���k��;��;��b<ԡ�;%}�=E�>��>J��>J��=$3��D/>w���XL��S�==X��_ZB��c��~�*B.��
5��&A>�T>&a������?D�Y>��;>�z�?�t? �>_&�X�վ#&��\qa�lT��t�=��>m�A�5�;��t`�e�L�V�Ӿ���>2�>R�>��l>�,�t%?�n5w=��ᾄL5� �>O������W��<q��B�����&i���ݺ��D?(>����=~?��I?�܏?V��>@����ؾv0>c�����=��q�����b�?f'?���>�*쾼�D�?�/N=Ef�>?����$6�]5���_�^ۯ�&"��㚺>׀��{����C�S�������+L4��oW��8�>H�b?�o�?���Ȋ�0싿��,:�;��E?�`�?���=@x)?�
?�
*�ޫ����T����=_ؖ?���?l��?�O�>X��=����m3�>D	?!ϖ?���?�as?��>���>�ۚ;�-!>`�����=7>[�=���=V?JY
?\�
?�H����	�������c�]���<���=*�>�l�>�sr>n��=�i=�=\>�Ǟ>�Ə>�ce>1S�>Gk�>�̣��I$���>�d��|��>nv9?F�>���=bӂ��+���6�2F�� ݽ�U�<�\,=nq�=tGQ�]���G����>�#Ŀ�͗?��">�?����>�ľ����k'>k�>)���?`��>9�>Oè>?C�>�\ >P	�>>�>iGӾ�>~���d!��,C�~�R�j�Ѿ�{z>Q����	&����Dv��-CI��n���g�rj�>.���;=�н<H�?+�����k��)�y�����?[�>�6?Bڌ������>���>�ƍ>�K��P���0ȍ�"h�y�?1��?"ud>}R�>�GP?gE?�O���T���S�+*e�]C8�� a�{ P��������e�=���P?�x?u�3?|�L=�Ro>n/�?�]�6p��C{>�).���6�3�=�\�>�m���S��Iپ�}�;��RK�=W�U?��?��>�eڽ倾<}Cu>u�5?�\?���?�g?=tI?̧="K?�>�i)?��;?
��?�%?9�?��9�^�=�P<@�=#DQ�#X���4)�Wb�@~/�EY�<jd�;T������=��7=����A?2>>��<��=&�^=��%�>U\>o<B>���>�Y]?a+�>�6�>��6?=�q{8��G����.?Z�6=�Z���F��Ql��C��� >��j?��?o�Y?#8e>�:A�i�?�e >�ى>�#>#QY>��>����B�T.�=i>� >ߛ�=L� 	����	��'��Y��<Q>?M�>�`>��r�C2F>�G������Dլ>+��t�o���[w�b�<�84��5�>`?Y ?U�=~&�7�0�w�k���?��(?��?>��?OG8>(�����.a,���t�콍>�%J=� �ʹ��ӧ��8M���<u>>o޾�Ԡ�Iqb>����m޾��n�pJ����VOM=	w�nV=��b�վ 
����=L9
>������ �"��7۪�D+J?��j=�v�� U�8t���>8��>�ۮ>y�:�r�v�h}@�4���:~�=��>�;>�9�� ��yG��3��|>C�A?md?po? �1��@j�g(�k�۾@pG�<�뽱�?$�?\�?6�>���=�ξn�*����#i� t�>���>(>�"�J������Ҽ�P��r�>��>?�H>0�?�{;?�?�@S?Q,?���>!��>S�&��J!?	�?O��=�M�o�T���,�W6�޿�>��#?C�?��.�>��?��#?�$.?�qO?D��>9e�=�f�E�V��`�>�Y�>�TS����'�<>��X?� �>MZM?@+|?��C>�+��վ�砼m��=�N>l.?�&?�m?���>i�>����D~=���>�%c?�??�p?�^�=�6?A�0>���>,�=�|�>���>j�?�M?iur?@J?+��>us�<�3��K����o��i���:�!E<��p=`���xu��6 ��;�<8�;�˶�Қ~����CG�E@�����;:q�>�r>zڔ�G2>��žie����>>�{���㛾Pr��c�:��{�=�_~>�?���>�R"����=;�>H��>���Ӑ(?߀?4h?��;ջb���ھ'hJ����>�WB?I��=��l�/�����u� �a=��m?(�^?H+V�9����a?&B]?�X�F:�h�ľ7hd����}�N?iJ
?�}C���>3V~?\q? =�>��i���n�(D���Nb���h����=깛>���+c�6J�>��7?e��>�I\>)#�=�z�o8���?���?��?��?��(>�Hn��߿�AҾ�(��#�d?
:�>����Q�?�������]싾r���at��D����W�D�w#���y�}��rwν'8>rc?�l?^q?�<e?/G���r��+b��S}�Hf�?��6��'D��[��/-����0%�R��U����+>by�ͳC�l�?�'?d/����>I	���ﾤ"ξ��6>H؝�ԙ�v��=�hz�!�F=�^=ej���0����� ?&�>���>�<>?+Z]�?���2���8�%��2>:~�>j��>A��>��;��>�zܽ�5ľv�z�:w��?�>� Z?J?d�i?xU'��)�`r��3��&�<�ʚ�}�=�Z^>Xu�>$�ͲA�QE7��XQ�̴u����̶��`�辨W=@�?<��>\��>^�?c0�>I�˾%���.=�����[�;���>y\p?��>o:|>��<���%����>�jt?�?p>J��0�R�k�O����>	Z?mR,?�/�>+��L����"����;�ȿ�=�+|?0�D�Zf�V�'>�G?�i�==�9<���=�X�����]�xw���)�<_:?c�N=��1>���#%�qaq��ݭ�K")?/�?�摾�*���>��"?�d�>�p�>DF�?��>Eb¾�S﹭,?'�^?S-J?��@?V`�>��=��� Ƚ�'�Bi+=���>��]>�yp=�K�= _�	[����'�?=�=�ZƼ��>Y<e�����h<=I85>�:�\K��Ӿ��w{۾A�	�θ�5R?�Љ���@��G;���Fxx�?�7�>i��X`��-e�����%�&��x�?���?2.C�/�i�踙�������E��>�4���¼�ն���^�t̾�����OX)�eH�,eS� �U�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >ZC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾k1�<��?7�-?��>Ǝr�1�ɿc���s¤<���?0�@�zA?�(�����`V=���>�	?$�?>�Y1��B���UZ�>�;�?^��?�nM=�W�J�	��{e?G<(�F�z�ݻL�=0�=%L=��(�J>aI�>��TMA��@ܽ0�4>KЅ>�"�á�%�^�d�<q{]>��սY���A�?�Q���w�/{��ˀ��;پf?��>�Ր�aA?�%g��.ѿUgZ����?.��?�m�?J>?��k���>,fԾ:T\?QTI?��>g���`�e�=�L���I�>B����^��
�=��?(�>�԰���?��p���ͽV,�����(�ƿ�R$�w=��je=�Z�:�佗�<�7�ܽ���o歾}�н*X=n5�=q_D>��{>uU4>�9m>z<Y?�p~?V��>�u&>���}���N�n�ռ\�T����/���2m� �վ����g��������F��� =���=�6R�����l� ���b��F���.?4w$>U�ʾ�M��n-<*qʾ���%焼Cޥ�;,̾��1��!n�P͟?��A?���S�V�+��3J����3�W?�Q����ꬾY��=���4�=�$�>���=���N 3� ~S�`0?e`?a����;���M*> � ��o=��+?1�?G9Z<��>�+%?)�*�a��H[>n�3>���>ė�>�
	>����:۽gz?�zT?���ޜ��Ґ>�r��N�z��_=.�>V�4�:i缂I[>i��<��BD[�v����<��V?�_�>��(�x2�������(�!�:=�Bx?��?⿢>y�k?K�B?�H�<B����TT����Pv=�aW?��i?�m>j
z���ϾO����4?�ud?w�M>xIh�l1羪a.�t�_�?j�o?TU?0���u~�����\�Sq6?l�u?|g�������.��,�>d��>�H?�R��h�>YK-?@5��B��s��ݳ5��4�?�@���?,����q�]H�<8��>�`?�N1���������ľ��
���>������j�1k#�����H?�3�?��>���,���!�=�(�� Z�?��?~���i<A �9#l�eD��!�<3�=E���w$�Ʌ��7�\�ƾ�
��~��Wh�����>�N@���(�>��8��/⿘CϿ����Ͼ�
q��?��>��ʽ�{����j��u��SG��H��a��G�>��>�ė��\���~��!A�!�(e�>�*ͼ�E�>=r�]^¾,��t�
�`o�>���>H$�>`G6�����5��?w��I�п�t������8x]?��?�K�?��?�V!=D����d�c��8UI?�q?��b?�4#<��J���<�$�j?�_��qU`��4�xHE��U>�"3?�B�>O�-���|=�>���>g>�#/�x�Ŀ�ٶ�<���X��?��?�o���>p��?rs+?�i�8���[����*�%�+��<A?�2>���C�!�B0=�VҒ���
?Q~0?{�c.�l�_?5�a�{�p���-���ƽCۡ>��0�e\�\\������Xe����Ay����?7^�?��?���� #�W6%?��>��8Ǿ��<��>!(�>9+N>DJ_�ݴu>����:�Mh	>���?�~�?kj?핏������T>��}?�{�>n��?R�>]�>b@�=�ٵ�(_�����=>�M����>n�R?��>]_�=��3���2��BM��*Z����b;����>��X?-�9?��>�rĽ�^L�!�d]���'W�d.
=�޽h��Mت��<W>@�\>WH>Fi�����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>D�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji����>c��H��|��T��f�1��W�=�m?��ap�>�fd>>ٵ���k� ]���z���?>2�?���?u�>�w?�3k�0V����=	?�f�?���>�A�>�C��B�>�2?QҤ���Q��ھ�fN?~�@�@X[?����+U俊묿:^���玾��>F�=;��=�J���,r=q��<� 6=/]��-��>�>��>��N>���=4�>��M>����.���睿�����<����.�����*�o�վ�}	�?;���~Ǡ��� ���¼�W;�����AЌ<u>1�j?��L?ƸE?8m�>hA�=�b>+)Ⱦh�%>��0��>\��>w�C?��E?jH"?F��Lo���y�[hu��X���
Q�@[�>�f~>���>�?���>&V�=WR�>��^>ZB9>�?�3�=�Т�S�Y=eV>���>���>G] ?pC<>�>Aϴ��1��@�h��
w��̽.�?i���M�J��1���9��̦��h�=Bb.?|>����>пh����2H?���k)���+���>|�0?�cW?�>��#�T��:>���h�j��_>, ��l���)�d%Q>�l?� c>�ty>�a4���5�U�L�m<���4v>]�6?�u��\�<��iv���I�][ܾ�b@>�Ծ>����Wߕ�Y��qm�՚}=��8?\�?���)���x
u��᝾x�O>"�T>��E=/b�=��O>���ģֽ��M���=�P�=�f>?�@->��=��>-W��� O�6w�>1@>A/>��@?\&?@����[��{H���[/��s>��>�>�@>�QI�8c�=���>[�_>9��&����c���B�w�X>n+{�(\�^�|�r�=(g��-��=y�=����:���?=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�w�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?�jN>���?z�r?T%�>�㞽��0�*���@��55�=��<<}�>F>9���ٔ@��l������~�k�����c>^^=��>;-ؽ�����J�=7n�_��)?;����>��V>A�:>�,�>)�?�>�>���<��pW�������I?ܐ?�Q��=k��Έ<��=�L�fM?F�2?�E��޾�%�>�_?˸�?0Y?r��>9�������������`M=8;>���>�P�>����٧Y>�r˾��&�3�>�Ï>�����?˾�����SO�>]v"?]��>�>=�?/�%?�w>-�>�H�vi��^:C���>g��>�s?��?�?�����{0��o�����YiW���O>��{?��?�<�>Q1���q��j��gT��U��C\�?*�g?��ٽ�?�s�?tD?�;?��^>b�/�G1߾#��廆>��!?���'�A��,&�q���?aZ?&��>�3���@׽��Ӽ��{@���?�&\?* &?s���a��5þ�>�<��%��DH���;��C�N�>�m>[m���=V�>=��=a�l�YJ6��bj<b��=%o�>�@�=�,7����=,?̈G��߃�U�=��r��vD�X�>"LL>� ���^?ȃ=��{�D���u����T�� �?���?j�?F*��Y�h�U%=?��?.?�(�>�A��؄޾��ྷEw�.}x�pu��>���>=n��循���#���*F���ƽ�NB�r-�>��->Vf	?Q�?K��>� �>{�`��_�#�#�����T�������Q�M����:��k/�����Y���p���Z����>��,y�>j^?�5�>���=�G>(i�[��>/��>w^v>Ᏹ>��d>��=��=!'<�Y�cKR?x���g�'����{���c3B?zrd?�/�>�i�򉅿N��>�?s��?}s�?�Av>�~h��,+��m?4<�>d���p
?hM:=�G�RB�<U��l��|6���%��>�>׽ :��M�of�-j
?|/?5퍼.�̾�6׽��۾��=�}?�"?�3%�:�X�x@��^	k���I�����f㉾�þ�=$�4�Tݐ�q(��1|���Q"�_�=1p6?���?�{Ծ`�gھcw��+:��\>@�>d<�>G�>f>Z��q<A�I�r�C�#��b�WD?|�f?8ݑ>�S?#V:?]JL?bxS?K��>��>�����c?[�)=���>�]�>�H?\"?@$0?�A�>?,>։��A��v��zH?'?�E/?��>cw?��G������=C&��?f@�>��Td<l��=U�߽L��<�G�=<M>�Q?S��p�8����~ k>	�7?���>0��>���t4�����< 	�>8�
?�@�>�����vr�
`��N�>Q��?����Q=��)>%��=/����1к�f�=��¼k��=�킼F;�Z? <�d�=O�=0�p��R��a~�:Z?�;b��<��>� ?h�>�Y4>�ž-B������=�'4>QT�>U>p`��y��y�z��t���r>�?�R�?Q�&>1�=�ԉ>E���N��8���(��63
>�d??yZ{?y_�?�H<?�;$?�<����>��x�������W�?p!,?��>�����ʾ��ˉ3�ҝ?m[?�<a����;)��¾�Խ��>�[/�]/~����8D�)����B��/��?뿝?�A�K�6��x�տ���[��p�C?"�>Y�>��>[�)���g�v%�}1;>��>mR?��>+HP?��z?�tW?��Q>57�b쪿i���D�M���>V0@?��?�W�?K�x?���>�v>}i;�q뾨��?�� /ٽ���M�=(�N>G�>O��>0�>�R�=�`��Up���N���=�d>_�>��>R�>�uq>���<��G?���>&<��,������nу���=�]�u?K��?x�+?�=lz�: F�-���!�>j�?x��?,4*?ϗS�E��=͆Լh涾r���>�ù>�9�>5%�=�BF=|�>s,�>���>�@��`�l8�
�M�,�?�F?��=��ſ��q��q����w;h<�ђ���d�vǔ��[�Բ�=Ʃ��خ�����$
\�/����~������Ꞝ�=�{�a��>��=w�=��=�3�<�ȼ��<�K=���<�=��n���q<T9�p4Ȼ����s��>\<�H=�.���ɾ�B{?��B?��*?ǚC?Κ>.6>T�4����>�Ʒ���?l9P>Y-D��5��5�1��b�������Zؾ`�ؾ�b������v>;�d�"=>��6>���=�#<�*�=a;4=J��=�b�<�E=�$�=���=œ�=�=+C
>.T>V�y?�����沿�s[�(�����0?VM>y��>��F���T?e�A<�儿D%��+��}�i?�!@�a�?�T,?�㈾ɫ�>ҟ[���=lqh>l���M����>���T�>�F< s�奡��KM��q�?أ@�E6?�2���ٿ��h>�� >4�>��T���#�?q��2��nW��N"?U>2�[#پ�Z>�!=F<׾G�ھ�m=��3>��<G��_��U=2}���k=��=���>@R>���=�ҽ�^�=�Z�<��->Vx>��7<�]��7q�>��<�@�=�M>��E>�\�>6�?I�3?��b?�X�>^�z�VaھƤþy��>A�=��>W�=w	>�V�>u�(?D�B?�M?ȃ�>6��=��>�U�>��+��t���ܾ����
��<gM�?��?|V�>�ep=�eM�#�$�b�;���ܽQ?�2?J�?k�>�U����9Y&���.�$����z4��+=�mr��QU�N���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=$�����<�vż�����u&�:�+�1�����;r��;B�]<]��;�c�=Q�>ץ>��>,5�=v0��g&>b����H�?�=�����oE���a�`�}�G()�}�+�c�<>	fS>�ýS����(?��T>�	I>�0�?��t?�:>^��q6о.�� tN�-K�u��=���=��Q��t=�ܒc�@�M�)9ʾ���>��>O�>��l>],�a!?���w=�
�[5�F�>�����t����2q�>��1����i�H�޺ΜD?�C��c��=~~?��I?1��?t��>\ژ�܉ؾ\M0>�\��=��1q��9���?0'?n��>���D�����6X����>����q�3��2�S���\�����}">��Ǿ���>�BW�� ��%d)�ό�2?�61?��?^Va��Hq��,�� ���dU/?p�?㠎>G>?���>��p�3s��w���P*�=5܅?Y{�?g��?�,4<�)�=�k�����>|�?l��?��?-�x?QP9��:�>�7�=m�_>dл��Z>r��=%�=�$�=�u ?��>_V?����,�
��e辈�վ怾��s�	?<U'>g�x>o^a>�n">f=��=��c>z�>g{>r1>���>ͥ>Vu��̖��G
?���=�>\�I?��>�?�=�9e�iK����=A�����:���]��}=:'�<�!����-���'�ݩ�>K¿~)�?(U>C�����>����>X���>>�)�>�7H�s�?�5;<)��>`�/>02�>R�=@�>��>�FӾ��>��Od!��+C���R��Ѿ~z>(���C
&���|���BI��o��5g�j�&.��<=�P��<�G�?����k�k�}�)�����?�[�>6??ڌ����B�>��>�Ǎ>rK��Q���>ȍ�Rh�e�?���?�~>��q>�_?� !?�=�C��_�cs��+���h��U��}� ��S޾t@8�88W?_�r?��??���=j�c>6��?]� ������Ag>��9��H0��S�=[��>D�C�+�U���af�����ۿ=�^?祇?�?�/]��ck=�+�=��?|V?o!�?�.G?�Rz?�*��9I?�H�>N_#?E� ?�r?�++?Bo9?��ý��<\j���K>�dP�����������w�Uߗ���o �M���ʼ嗖=���_X5������=�7�=b57=��7>���<�>)�]?���>��>��7?��6l8��y��B/?מ8=!ς��A��hҢ�g:��>��j?��?�BZ?��c>:B���B�t
>6L�>��&>�$\>i�>C��ΠE�d��=F�>��>P&�=D�N��߁��	������Y�<��>W�>4��>�FJ���>�쏾\�Z��0[>�'Ƚ5D������-s�;�J�9���K�>�,V?y� ?nm�=�pY���i�'+?�x#?.!>?��?2Zg>���q��� ����m�>�,=�Jʾt����N��u,c�"�x��"�=X�ž�꠾׺a>�����޾\@n���I���,5L=jZ��cO=T=��c־�9�2b�=�
>�r��d� �����䪿6�I?G�g==$��f9V�}���Ș>�ۘ>�/�>��9���s��+@����=��>��;>����&�,G��#�Ň�>�H?��`?ݬ�?_ ���\q���>��뾄(���}�dy?]G�>B ?_�B>�>�=&���*���g�tH�G��>�s�>���GE�������m��+�>[��>.�>03?z2N?5�?4$`?�T,?��?���>�U���Ǿ�A&?D��?��=��ԽI�T�2 9�CF�Z��>��)?~�B�Ϻ�> �?G�?��&?�Q?:�?��>�� �TD@����>�X�>^�W��a��h�_>8�J?i��>�;Y?.ԃ?��=>d�5�i뢾�ʩ�W�=H>��2?X6#?�?���>�<�>�����w�=��>�c?A�?ԇo?C��=�u?-�3>\��>��=���>£�>S*?XN?��s?b�J?�j�>�\�<��������6Wu�;^c��GP;�Wa<y�n=����?�����.�<�@�;�1��ሼ�켚�G��t��/<MN�>ws>�ɕ�9�0>-�ľm[���@>r|���^��D��E�:����=!@�>�?�}�>�#��m�=���>�1�>Y���^(?�?9?-� ;x�b��۾�SK���>l�A?���=��l����u�u��He=;�m?H�^?@~W�t���"�a?t�^?;b�:�X�þX�f�13�gP?��
?��I�H��>��?4�p?���>1	f�Z�n��]��"�b�Żp�6�=g@�>u�`d�}��>��6?_�>%r^>o��=�ܾjv�Ǳ����?ر�?���?�;�?�&*>��n�,�߿������#E?D��>�h�1�? 9��h� �G���A���K��ٰ���AM��(��T������o�p����h����>xWu?x�r?��s?�����x�Óo���a�ǎF�y{�!�о��R��/m�5�Z�"��r�������,�<=6>V�~��B�|��?�<&? E-����>�^��H�D�̾XB>襡����O�=�I��K=�_=i#g��.�绮�
�?rg�>e�>I{=?�j[�d�>�u�1��7����:�0>Oޢ>�Z�>���>6���:1�W�IIȾ����-�˽�Iy>4�g?kJO?�5l?��i�0���u�w��erJ����e>�@]>�=�>�;6�G#���,���J��mx����C��`����<�#?M�p>H�>X��?��>r��dR����k��(����=���> mh?���>x}�>"�
�h))�F��>�b? �>��>�־��8���V�?��=y
�>��? N#?�F�>������q�d͏�:����M�I�=�nz?�W��E��Д>��??�(�=�>ºQ>�&���ؾ��)����u~=�>�9>�ͼ�������`$~���ܾ��&?�v?_Ȓ�oR-�L��>�"?i��>錡>bՂ?a��>j�Ⱦq�3:ˍ?�(`?�RK?�	A?qD�><X ='�ý������0�u�p=Y�>�[>��I=#��=��!�p�]�h��~=�=<����k��0�l;1zż9%X<�=d�?>�xۿ�CK��vپ���A�PD
�\,��}����c���	�
`��_�7x������'�'^V��]c�M��� m�px�?�:�?BW�����%�����������饽>urq���~�����2��m��R��C�S]!�G�O�ki��e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?7�y?��7�"���8�� >eC�<�,����뾬����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾y1�<��?7�-?��>Ďr�1�ɿc���|¤<���?0�@}A?-�(���쾑V=?��>'�	?$�?>�S1��I�����pT�>j<�?���?H}M=g�W��	��e?�|<��F��ݻ��=><�=�F=�����J>fU�>"���SA�l?ܽ�4>1څ>�~"�j���^�g��<��]>��ս�:���e�?.mf�Q〿1����7�����=�wj?w�w>�f7�1Y?a�[�EϿz�&�ӑ?c��?��?A�H?�)ݾ~%d>5¾N�[?�i@?�n�>41�,R�0K>3̾q�>�~"�m�h��ב=��?3�>�.����0��Bo�&���t�<�� ���ǿ�"��!�܎&=#v�;/�:���x��T�I�M茶�?l�w�ս�؎=$��=�.T>�>>�O>0�O>|�U?�4i?��>�[&>=��]�� �Ͼ�q��u����!�@%���?$�~ͤ���>���d	�������Q����=�g�=.8R�{���=� ���b�}�F�~�.?�m$>��ʾ��M�|x*<�nʾRǪ��}��8ϥ�C,̾�1�)n��Ɵ?��A?����V�!���N��m��"�W?�D�x��nӬ���=���=�(�>���=t���3�{S� j0?=\?X���P����)>�O���=7�+?2�?�[<�!�>R%?�+�t�k�Z>D�3>��>��>��	>���<zڽ\v?�oT?!"�2���ː>�A���Qz� Ib=�{>Y5�,���y[>��<�
��(h^�������<�V?/0�>�'�ބ�J��I���4=R�y?A?���>P�l?oFC?�.\<Fy���S�9�r�X=dX?�k?�	>���RBϾ@�����4?D[d?a�M>�t`��f�(�+�7��O?6�n?�4?�XƼ�}�
���o0�R�5?�v?b�^�{����&��'V��b�>~��>
�>�<:��Ƴ>�s>?�\#��4��V���1@4��מ?��@Y��?��J<���ċ=�?�>E�N��RžN߳������l=���>{����Mv�p��Q+��8?w��?N&�>�ւ����D��=#4���E�?���?Oj����c<;��Ul�m��^�<�٩=��"����7���ƾڌ
��_������ˬ�>	U@U罗u�>�9�;"��CϿ�셿�XоG�q�M!?7�>D�̽�룾��j��u��JG��H��(���J�>�>4�������x�{��q;�2��.�>���	�>B�S��&��+��� T5<-�>Ԯ�>丆>("��:潾@ř?�d���?ο�������c�X?�h�?o�?�n?t�9<��v�
�{�if�U.G?y�s?Z?J%�t6]�$�7�#�j?�_��qU`��4�wHE��U>�"3?�B�>O�-��|=�>���>g>�#/�w�Ŀ�ٶ�E���X��?��?�o���>p��?us+?�i�8���[����*���+��<A?�2>���D�!�=0=�`Ғ���
?R~0?6{�h.�9�_?�a���p���-��ƽ�ۡ>߲0�WX\��Q��"���Xe�0��L@y����?t]�?a�?_��
�"�3%?
�>c����+Ǿ;w�<9o�>8�>�2N>��_���u>�
���:��Y	>׮�?�}�?bj?ڕ�������6>��}?�f�>�o�?eP>s��>_��=E��h�7�-0>g�>�x�Ĥ?�kQ?V�>�l�=C�;�*u1��K�t�U�2P��	?��Y�>��X?�E?�`>K��� 鼸 ����c7�tt�U2A�Bp�����E�C>��C>��>��K�R�ھ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji���>)��@��:��O����Y��@L>��L?���V��>���>.�= /q��e���Nn�<j�>. �?4�?o�?��?�%���e��3p�=��>�^�?m/?�0Z=�*�{�B>4�?��NCi�E�����f?=�@�@�V?2�����ѿ䲖��������d��=Y��=���=sz(��q�=>Gb�4gl=�R�=I�a>��>`�q>U>�>[�\>�=�ǂ�;l�t���i����F���.�|t6��-��u��񚣾�H1��Щ�7UԾ�����"��V)�vs��~�F�(aU��9>�*\?ibO?��k?K� ?�x�;E(D>�dʾ���=��P���=>�Ӭ>��G?i�@?�?���þ�d�ұ�������Ir�:k�>��t>�?ܘ?���>����,�>gt>̹�>�7��/">jH׼~d�=�)�>�>��?m��>��;>��>F���&.���Xh��u��8˽��?�R��E�J��+���������8�=�p.?��>����:%п��K
H?�`�����+�,��d>�|0?�XW?M>�հ�j�N�N4>����i���>w��2�k�MN)�~uQ>�a?��L>VW>��5��;�O�D�u2���y>0.?�$��x�m�)w���K�>ؾ-69>Ո�>�����M�,����^��I�^��<k�7?���>��ӽ4ɮ��V�寇��O>"Cz>��\=%��=��[>����HYs��r-�ԨS=�!>�W>�?��3>���=�M�>>���[>^� ��>�}?>">,>ĥ9?'� ?~����<��>�Ddv><^�>σz>f�>�1C��\�=��>�Z>x�\�����m
�r95�&zj>�5/���B��^�`G=���{��=�*n=�g�`�5��|0=�~?���%䈿���d���lD?T+?H �=�F<��"�E ���H��C�?q�@m�?��	�ڢV�8�?�@�?��%��=}�>׫>�ξ#�L�ޱ?�Ž6Ǣ�Ɣ	�<)#�fS�?��?��/�Xʋ�9l�}6>�^%?�ӾPh�>yx��Z�������u�m�#=Q��>�8H?�V����O�c>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?toi>�g۾:`Z����>һ@?�R?�>�9���'���?�޶?֯�?��]>p��?=F|?w.�>0#���"�誠��1W��H�>���~;>�u�>����v�1��ۛ�����4|��<�R�|><��;�U�>�E����V�!>��S�)��q=���>�$>ߔ4>؝�>��?�5�>w�>��C<"Q���~�0�Ǿc�K?���?5���/n�2?�<���=ү^�D&?aH4?��[�^�Ͼ�٨>R�\??�[?�^�>����>��迿}����<��K>�2�>�K�>�	��/JK>X�ԾY4D��o�>�ϗ>^J���8ھ'+��9آ�7D�>�f!?O��>�Ю=��?e*+?�z>H�>��M�����>��1�>!��>�|?���?��?�Ѿ[�;�"����B��;�Z�l}�>0��?!�?^��>|���Ǘ�����4�aQX�y�?U?�`��}�?���?��@?w	*?�T>�tG�N�xF��O=�>t�?(���iB���(�*���	?�Z?{�>|w���-
��%P����0���?
?�
[?�#?��,da�.VӾn�<J ����<'.c�eüI�>�#>��E�$~�=6.>vP�=^bM�u�#�I0=2y�=K��>]�=h�&�����<,?ЧG��ڃ�5�=k�r�:xD���>}IL>:��ӫ^?�k=�7�{����Px���
U�� �?Π�?�j�?�����h�%=?��?�?d �>�K��G}޾A��<Mw�9{x�pv���>���>l�l�����������F����Ž��1�y^�>��>�Y�>4�?;'�>�N�>Lm���Q�u�l���j�a���-<�������T��El��`�;�7���TՈ�!��>+�*�ī�>XC?^�?>XN�>]-�>������>�*>�G>��>"�A>��>"��=�x:=
n*��KR?�����'���辪���g3B?�qd?81�>^i�4������~�?���?Ts�?R=v>�~h��,+�qn?�>�>;��Jq
?�U:=�5�;;�<!V�����w3��Y�$��>5E׽� :��M�Onf�ej
?�/?�����̾G;׽�Y�(�<�6?�$?����mZ���{tk�
??����0�q���h����1|j�#��@u�������t��я�2�/?�˓?��Ǿk�߾Ix��]Q{��QC�k��>S��>��>��>�|=��6�mJ�(�m�|��:`����>=d�?(^�>#aJ?Z<?��R?�O?"��>˃�>맾���>���;sV�>[K�>�^=?"�+?2-?/v?�
'?�Z>Y�p����Ҿ m?�v?&i?�c?��??�z�۬���֒8�S��M��r[���f=X�=��ŽN[�|z�=-�i>tX?Q���8�����"�j>P7?}�>���>)��)���:�<��>�
?oC�>�  �;}r��b��V�>���?���x=��)>R��=������ҺX�=���q�=k(���x;��T<h��=��=�Wu�,􊹸7�:^\�;Do�<��>"�-?�j�>E�k>y�"�$�w���=?t}>GJW>V>�����㓿9���4�]��F>� r?�ɛ?�L>Z>�,`>�z�sK���A
�6Y߾�ـ=#5 ? S?J[?��?�[[?%�?z.�Ğ־ ��f���	w��m?w!,?��>�����ʾ��։3�ڝ?i[?�<a����;)�ݐ¾��Խα>�[/�h/~����=D�u텻���Y��5��?�?GA�V�6��x�ڿ���[��z�C?"�>Y�>��>U�)�~�g�s%��1;>���>kR?��>�7P?=/{?\{[?�FR>�8����T��=�"�۵>�@?���?*ώ?5�x?O��>r�>�.���������򽽄���S=�R[>�>�k�>q-�>���=�Ƚ�����@�S��=�cc>���>�>!��>��v>��<��G?���>�O��V��G򤾪̃�9q=�Y�u?���?,�+?qN=�����E��A���5�>�j�?���?�-*?��S����=�uռ�඾`�q���>JŹ>+�>5ؓ=0G=�v>��>��>6<��Z�fo8�n�M���?�F?B��=��ÿ��q�`w��f��z�<4刾�3`�{���͞X���=A��!!�خ���hZ������t�������a��������>��i=�Q>��=?b�<��޼��<��d=`�<�v=�S��}<�7�8���\��!uV���j<�8`=�|�K ʾ�g}?%9I?�+?�D?-�|>�>��*��_�>Mt���f?�UV>��=�曻��W<�w=������Oؾb�־c�����?�>^�@���>��6>���=��<���=��}=jʑ=�'���#=���=q��=�f�=���=RU>�>[ox?�֌�B?����P�{���:�B?:�>L4�>�G���Y?F��=ZHy�)��}>Ӿ�m?� @(��?��8?ӕ�MF�>�uľ�ý�>�gR��n6>kK�<�1\��KQ>�E>��7�O��J��)��?#��?}�2?�6��	�̿��b#>��=�}S�LV3���E�C�3�m�P�??��4��ᾦ.]>��<=��ܾXZȾ��k=Ⱦ6>1�8=��5�"�c��͒=�Ĩ��b=�!�<� u>��7>�@�=vP�3��=ٕ=��>�g>d�<	�»�':��Db=�-�=l�k>Vz>WS�>��?�F0?��c?&:�>��n�uyϾ@*��7��>��=׹�>٘�=
�>>f��>�.7?�zD?tL?�<�>(ԋ=���>fS�>ek,�+Gm�l���&��w^�<ol�?��?f�>S΀<��A�����=�`"Ƚ�?B1?��?�2�>
F�|���F&���.�<̘��ʤ987,=r�I4U����M�H��j��=���>��>p�>g=y>��9>MTN>K�>�i>��<���=X׍�a"�<����΃=�y��)�<*ǼV����)�E�,�4���k��;��;��b<ԡ�;%}�=E�>��>J��>J��=$3��D/>w���XL��S�==X��_ZB��c��~�*B.��
5��&A>�T>&a������?D�Y>��;>�z�?�t? �>_&�X�վ#&��\qa�lT��t�=��>m�A�5�;��t`�e�L�V�Ӿ���>2�>R�>��l>�,�t%?�n5w=��ᾄL5� �>O������W��<q��B�����&i���ݺ��D?(>����=~?��I?�܏?V��>@����ؾv0>c�����=��q�����b�?f'?���>�*쾼�D�?�/N=Ef�>?����$6�]5���_�^ۯ�&"��㚺>׀��{����C�S�������+L4��oW��8�>H�b?�o�?���Ȋ�0싿��,:�;��E?�`�?���=@x)?�
?�
*�ޫ����T����=_ؖ?���?l��?�O�>X��=����m3�>D	?!ϖ?���?�as?��>���>�ۚ;�-!>`�����=7>[�=���=V?JY
?\�
?�H����	�������c�]���<���=*�>�l�>�sr>n��=�i=�=\>�Ǟ>�Ə>�ce>1S�>Gk�>�̣��I$���>�d��|��>nv9?F�>���=bӂ��+���6�2F�� ݽ�U�<�\,=nq�=tGQ�]���G����>�#Ŀ�͗?��">�?����>�ľ����k'>k�>)���?`��>9�>Oè>?C�>�\ >P	�>>�>iGӾ�>~���d!��,C�~�R�j�Ѿ�{z>Q����	&����Dv��-CI��n���g�rj�>.���;=�н<H�?+�����k��)�y�����?[�>�6?Bڌ������>���>�ƍ>�K��P���0ȍ�"h�y�?1��?"ud>}R�>�GP?gE?�O���T���S�+*e�]C8�� a�{ P��������e�=���P?�x?u�3?|�L=�Ro>n/�?�]�6p��C{>�).���6�3�=�\�>�m���S��Iپ�}�;��RK�=W�U?��?��>�eڽ倾<}Cu>u�5?�\?���?�g?=tI?̧="K?�>�i)?��;?
��?�%?9�?��9�^�=�P<@�=#DQ�#X���4)�Wb�@~/�EY�<jd�;T������=��7=����A?2>>��<��=&�^=��%�>U\>o<B>���>�Y]?a+�>�6�>��6?=�q{8��G����.?Z�6=�Z���F��Ql��C��� >��j?��?o�Y?#8e>�:A�i�?�e >�ى>�#>#QY>��>����B�T.�=i>� >ߛ�=L� 	����	��'��Y��<Q>?M�>�`>��r�C2F>�G������Dլ>+��t�o���[w�b�<�84��5�>`?Y ?U�=~&�7�0�w�k���?��(?��?>��?OG8>(�����.a,���t�콍>�%J=� �ʹ��ӧ��8M���<u>>o޾�Ԡ�Iqb>����m޾��n�pJ����VOM=	w�nV=��b�վ 
����=L9
>������ �"��7۪�D+J?��j=�v�� U�8t���>8��>�ۮ>y�:�r�v�h}@�4���:~�=��>�;>�9�� ��yG��3��|>C�A?md?po? �1��@j�g(�k�۾@pG�<�뽱�?$�?\�?6�>���=�ξn�*����#i� t�>���>(>�"�J������Ҽ�P��r�>��>?�H>0�?�{;?�?�@S?Q,?���>!��>S�&��J!?	�?O��=�M�o�T���,�W6�޿�>��#?C�?��.�>��?��#?�$.?�qO?D��>9e�=�f�E�V��`�>�Y�>�TS����'�<>��X?� �>MZM?@+|?��C>�+��վ�砼m��=�N>l.?�&?�m?���>i�>����D~=���>�%c?�??�p?�^�=�6?A�0>���>,�=�|�>���>j�?�M?iur?@J?+��>us�<�3��K����o��i���:�!E<��p=`���xu��6 ��;�<8�;�˶�Қ~����CG�E@�����;:q�>�r>zڔ�G2>��žie����>>�{���㛾Pr��c�:��{�=�_~>�?���>�R"����=;�>H��>���Ӑ(?߀?4h?��;ջb���ھ'hJ����>�WB?I��=��l�/�����u� �a=��m?(�^?H+V�9����a?&B]?�X�F:�h�ľ7hd����}�N?iJ
?�}C���>3V~?\q? =�>��i���n�(D���Nb���h����=깛>���+c�6J�>��7?e��>�I\>)#�=�z�o8���?���?��?��?��(>�Hn��߿�AҾ�(��#�d?
:�>����Q�?�������]싾r���at��D����W�D�w#���y�}��rwν'8>rc?�l?^q?�<e?/G���r��+b��S}�Hf�?��6��'D��[��/-����0%�R��U����+>by�ͳC�l�?�'?d/����>I	���ﾤ"ξ��6>H؝�ԙ�v��=�hz�!�F=�^=ej���0����� ?&�>���>�<>?+Z]�?���2���8�%��2>:~�>j��>A��>��;��>�zܽ�5ľv�z�:w��?�>� Z?J?d�i?xU'��)�`r��3��&�<�ʚ�}�=�Z^>Xu�>$�ͲA�QE7��XQ�̴u����̶��`�辨W=@�?<��>\��>^�?c0�>I�˾%���.=�����[�;���>y\p?��>o:|>��<���%����>�jt?�?p>J��0�R�k�O����>	Z?mR,?�/�>+��L����"����;�ȿ�=�+|?0�D�Zf�V�'>�G?�i�==�9<���=�X�����]�xw���)�<_:?c�N=��1>���#%�qaq��ݭ�K")?/�?�摾�*���>��"?�d�>�p�>DF�?��>Eb¾�S﹭,?'�^?S-J?��@?V`�>��=��� Ƚ�'�Bi+=���>��]>�yp=�K�= _�	[����'�?=�=�ZƼ��>Y<e�����h<=I85>�:�\K��Ӿ��w{۾A�	�θ�5R?�Љ���@��G;���Fxx�?�7�>i��X`��-e�����%�&��x�?���?2.C�/�i�踙�������E��>�4���¼�ն���^�t̾�����OX)�eH�,eS� �U�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >ZC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾k1�<��?7�-?��>Ǝr�1�ɿc���s¤<���?0�@�zA?�(�����`V=���>�	?$�?>�Y1��B���UZ�>�;�?^��?�nM=�W�J�	��{e?G<(�F�z�ݻL�=0�=%L=��(�J>aI�>��TMA��@ܽ0�4>KЅ>�"�á�%�^�d�<q{]>��սY���A�?�Q���w�/{��ˀ��;پf?��>�Ր�aA?�%g��.ѿUgZ����?.��?�m�?J>?��k���>,fԾ:T\?QTI?��>g���`�e�=�L���I�>B����^��
�=��?(�>�԰���?��p���ͽV,�����(�ƿ�R$�w=��je=�Z�:�佗�<�7�ܽ���o歾}�н*X=n5�=q_D>��{>uU4>�9m>z<Y?�p~?V��>�u&>���}���N�n�ռ\�T����/���2m� �վ����g��������F��� =���=�6R�����l� ���b��F���.?4w$>U�ʾ�M��n-<*qʾ���%焼Cޥ�;,̾��1��!n�P͟?��A?���S�V�+��3J����3�W?�Q����ꬾY��=���4�=�$�>���=���N 3� ~S�`0?e`?a����;���M*> � ��o=��+?1�?G9Z<��>�+%?)�*�a��H[>n�3>���>ė�>�
	>����:۽gz?�zT?���ޜ��Ґ>�r��N�z��_=.�>V�4�:i缂I[>i��<��BD[�v����<��V?�_�>��(�x2�������(�!�:=�Bx?��?⿢>y�k?K�B?�H�<B����TT����Pv=�aW?��i?�m>j
z���ϾO����4?�ud?w�M>xIh�l1羪a.�t�_�?j�o?TU?0���u~�����\�Sq6?l�u?|g�������.��,�>d��>�H?�R��h�>YK-?@5��B��s��ݳ5��4�?�@���?,����q�]H�<8��>�`?�N1���������ľ��
���>������j�1k#�����H?�3�?��>���,���!�=�(�� Z�?��?~���i<A �9#l�eD��!�<3�=E���w$�Ʌ��7�\�ƾ�
��~��Wh�����>�N@���(�>��8��/⿘CϿ����Ͼ�
q��?��>��ʽ�{����j��u��SG��H��a��G�>��>�ė��\���~��!A�!�(e�>�*ͼ�E�>=r�]^¾,��t�
�`o�>���>H$�>`G6�����5��?w��I�п�t������8x]?��?�K�?��?�V!=D����d�c��8UI?�q?��b?�4#<��J���<�$�j?�_��qU`��4�xHE��U>�"3?�B�>O�-���|=�>���>g>�#/�x�Ŀ�ٶ�<���X��?��?�o���>p��?rs+?�i�8���[����*�%�+��<A?�2>���C�!�B0=�VҒ���
?Q~0?{�c.�l�_?5�a�{�p���-���ƽCۡ>��0�e\�\\������Xe����Ay����?7^�?��?���� #�W6%?��>��8Ǿ��<��>!(�>9+N>DJ_�ݴu>����:�Mh	>���?�~�?kj?핏������T>��}?�{�>n��?R�>]�>b@�=�ٵ�(_�����=>�M����>n�R?��>]_�=��3���2��BM��*Z����b;����>��X?-�9?��>�rĽ�^L�!�d]���'W�d.
=�޽h��Mت��<W>@�\>WH>Fi�����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>D�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji����>c��H��|��T��f�1��W�=�m?��ap�>�fd>>ٵ���k� ]���z���?>2�?���?u�>�w?�3k�0V����=	?�f�?���>�A�>�C��B�>�2?QҤ���Q��ھ�fN?~�@�@X[?����+U俊묿:^���玾��>F�=;��=�J���,r=q��<� 6=/]��-��>�>��>��N>���=4�>��M>����.���睿�����<����.�����*�o�վ�}	�?;���~Ǡ��� ���¼�W;�����AЌ<u>1�j?��L?ƸE?8m�>hA�=�b>+)Ⱦh�%>��0��>\��>w�C?��E?jH"?F��Lo���y�[hu��X���
Q�@[�>�f~>���>�?���>&V�=WR�>��^>ZB9>�?�3�=�Т�S�Y=eV>���>���>G] ?pC<>�>Aϴ��1��@�h��
w��̽.�?i���M�J��1���9��̦��h�=Bb.?|>����>пh����2H?���k)���+���>|�0?�cW?�>��#�T��:>���h�j��_>, ��l���)�d%Q>�l?� c>�ty>�a4���5�U�L�m<���4v>]�6?�u��\�<��iv���I�][ܾ�b@>�Ծ>����Wߕ�Y��qm�՚}=��8?\�?���)���x
u��᝾x�O>"�T>��E=/b�=��O>���ģֽ��M���=�P�=�f>?�@->��=��>-W��� O�6w�>1@>A/>��@?\&?@����[��{H���[/��s>��>�>�@>�QI�8c�=���>[�_>9��&����c���B�w�X>n+{�(\�^�|�r�=(g��-��=y�=����:���?=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�w�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?�jN>���?z�r?T%�>�㞽��0�*���@��55�=��<<}�>F>9���ٔ@��l������~�k�����c>^^=��>;-ؽ�����J�=7n�_��)?;����>��V>A�:>�,�>)�?�>�>���<��pW�������I?ܐ?�Q��=k��Έ<��=�L�fM?F�2?�E��޾�%�>�_?˸�?0Y?r��>9�������������`M=8;>���>�P�>����٧Y>�r˾��&�3�>�Ï>�����?˾�����SO�>]v"?]��>�>=�?/�%?�w>-�>�H�vi��^:C���>g��>�s?��?�?�����{0��o�����YiW���O>��{?��?�<�>Q1���q��j��gT��U��C\�?*�g?��ٽ�?�s�?tD?�;?��^>b�/�G1߾#��廆>��!?���'�A��,&�q���?aZ?&��>�3���@׽��Ӽ��{@���?�&\?* &?s���a��5þ�>�<��%��DH���;��C�N�>�m>[m���=V�>=��=a�l�YJ6��bj<b��=%o�>�@�=�,7����=,?̈G��߃�U�=��r��vD�X�>"LL>� ���^?ȃ=��{�D���u����T�� �?���?j�?F*��Y�h�U%=?��?.?�(�>�A��؄޾��ྷEw�.}x�pu��>���>=n��循���#���*F���ƽ�NB�r-�>��->Vf	?Q�?K��>� �>{�`��_�#�#�����T�������Q�M����:��k/�����Y���p���Z����>��,y�>j^?�5�>���=�G>(i�[��>/��>w^v>Ᏹ>��d>��=��=!'<�Y�cKR?x���g�'����{���c3B?zrd?�/�>�i�򉅿N��>�?s��?}s�?�Av>�~h��,+��m?4<�>d���p
?hM:=�G�RB�<U��l��|6���%��>�>׽ :��M�of�-j
?|/?5퍼.�̾�6׽��۾��=�}?�"?�3%�:�X�x@��^	k���I�����f㉾�þ�=$�4�Tݐ�q(��1|���Q"�_�=1p6?���?�{Ծ`�gھcw��+:��\>@�>d<�>G�>f>Z��q<A�I�r�C�#��b�WD?|�f?8ݑ>�S?#V:?]JL?bxS?K��>��>�����c?[�)=���>�]�>�H?\"?@$0?�A�>?,>։��A��v��zH?'?�E/?��>cw?��G������=C&��?f@�>��Td<l��=U�߽L��<�G�=<M>�Q?S��p�8����~ k>	�7?���>0��>���t4�����< 	�>8�
?�@�>�����vr�
`��N�>Q��?����Q=��)>%��=/����1к�f�=��¼k��=�킼F;�Z? <�d�=O�=0�p��R��a~�:Z?�;b��<��>� ?h�>�Y4>�ž-B������=�'4>QT�>U>p`��y��y�z��t���r>�?�R�?Q�&>1�=�ԉ>E���N��8���(��63
>�d??yZ{?y_�?�H<?�;$?�<����>��x�������W�?p!,?��>�����ʾ��ˉ3�ҝ?m[?�<a����;)��¾�Խ��>�[/�]/~����8D�)����B��/��?뿝?�A�K�6��x�տ���[��p�C?"�>Y�>��>[�)���g�v%�}1;>��>mR?��>+HP?��z?�tW?��Q>57�b쪿i���D�M���>V0@?��?�W�?K�x?���>�v>}i;�q뾨��?�� /ٽ���M�=(�N>G�>O��>0�>�R�=�`��Up���N���=�d>_�>��>R�>�uq>���<��G?���>&<��,������nу���=�]�u?K��?x�+?�=lz�: F�-���!�>j�?x��?,4*?ϗS�E��=͆Լh涾r���>�ù>�9�>5%�=�BF=|�>s,�>���>�@��`�l8�
�M�,�?�F?��=��ſ��q��q����w;h<�ђ���d�vǔ��[�Բ�=Ʃ��خ�����$
\�/����~������Ꞝ�=�{�a��>��=w�=��=�3�<�ȼ��<�K=���<�=��n���q<T9�p4Ȼ����s��>\<�H=�.���ɾ�B{?��B?��*?ǚC?Κ>.6>T�4����>�Ʒ���?l9P>Y-D��5��5�1��b�������Zؾ`�ؾ�b������v>;�d�"=>��6>���=�#<�*�=a;4=J��=�b�<�E=�$�=���=œ�=�=+C
>.T>V�y?�����沿�s[�(�����0?VM>y��>��F���T?e�A<�儿D%��+��}�i?�!@�a�?�T,?�㈾ɫ�>ҟ[���=lqh>l���M����>���T�>�F< s�奡��KM��q�?أ@�E6?�2���ٿ��h>�� >4�>��T���#�?q��2��nW��N"?U>2�[#پ�Z>�!=F<׾G�ھ�m=��3>��<G��_��U=2}���k=��=���>@R>���=�ҽ�^�=�Z�<��->Vx>��7<�]��7q�>��<�@�=�M>��E>�\�>6�?I�3?��b?�X�>^�z�VaھƤþy��>A�=��>W�=w	>�V�>u�(?D�B?�M?ȃ�>6��=��>�U�>��+��t���ܾ����
��<gM�?��?|V�>�ep=�eM�#�$�b�;���ܽQ?�2?J�?k�>�U����9Y&���.�$����z4��+=�mr��QU�N���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=$�����<�vż�����u&�:�+�1�����;r��;B�]<]��;�c�=Q�>ץ>��>,5�=v0��g&>b����H�?�=�����oE���a�`�}�G()�}�+�c�<>	fS>�ýS����(?��T>�	I>�0�?��t?�:>^��q6о.�� tN�-K�u��=���=��Q��t=�ܒc�@�M�)9ʾ���>��>O�>��l>],�a!?���w=�
�[5�F�>�����t����2q�>��1����i�H�޺ΜD?�C��c��=~~?��I?1��?t��>\ژ�܉ؾ\M0>�\��=��1q��9���?0'?n��>���D�����6X����>����q�3��2�S���\�����}">��Ǿ���>�BW�� ��%d)�ό�2?�61?��?^Va��Hq��,�� ���dU/?p�?㠎>G>?���>��p�3s��w���P*�=5܅?Y{�?g��?�,4<�)�=�k�����>|�?l��?��?-�x?QP9��:�>�7�=m�_>dл��Z>r��=%�=�$�=�u ?��>_V?����,�
��e辈�վ怾��s�	?<U'>g�x>o^a>�n">f=��=��c>z�>g{>r1>���>ͥ>Vu��̖��G
?���=�>\�I?��>�?�=�9e�iK����=A�����:���]��}=:'�<�!����-���'�ݩ�>K¿~)�?(U>C�����>����>X���>>�)�>�7H�s�?�5;<)��>`�/>02�>R�=@�>��>�FӾ��>��Od!��+C���R��Ѿ~z>(���C
&���|���BI��o��5g�j�&.��<=�P��<�G�?����k�k�}�)�����?�[�>6??ڌ����B�>��>�Ǎ>rK��Q���>ȍ�Rh�e�?���?�~>��q>�_?� !?�=�C��_�cs��+���h��U��}� ��S޾t@8�88W?_�r?��??���=j�c>6��?]� ������Ag>��9��H0��S�=[��>D�C�+�U���af�����ۿ=�^?祇?�?�/]��ck=�+�=��?|V?o!�?�.G?�Rz?�*��9I?�H�>N_#?E� ?�r?�++?Bo9?��ý��<\j���K>�dP�����������w�Uߗ���o �M���ʼ嗖=���_X5������=�7�=b57=��7>���<�>)�]?���>��>��7?��6l8��y��B/?מ8=!ς��A��hҢ�g:��>��j?��?�BZ?��c>:B���B�t
>6L�>��&>�$\>i�>C��ΠE�d��=F�>��>P&�=D�N��߁��	������Y�<��>W�>4��>�FJ���>�쏾\�Z��0[>�'Ƚ5D������-s�;�J�9���K�>�,V?y� ?nm�=�pY���i�'+?�x#?.!>?��?2Zg>���q��� ����m�>�,=�Jʾt����N��u,c�"�x��"�=X�žfޟ��b>�����߾�;n�_eJ� V��R=�#�8FK=z���	վF������=*�	>�]��n� �t>���ު��bJ?K5j=����IV������>�>)S�>��?���x��Y@����=��=Ɨ�>�<>Bs��TﾆkG��1��>��F? Wd?G�?����	�s�woL����u����f���?��>r�?��B>]�X=B���h\�Z�e��'D�u��>���>����KH��Þ�6��~'�3�u>:o�> �<>=�?2N?`�?
�a?RW'?#(�>��>ҥ½u�ľy4&?��?�=�KԽ~KT���8�@(F����>b)?�B�ԗ>(�?,�? '?e�Q?�?"T>?� ��\@�~m�>U�>@�W�VK��5�`>�J?w�>�ZY?�؃?vd>>��5����𺪽��=	�>��2?sB#?H�?Tθ>�>�������>�!�?��?��?6��>l�
?�K�>�i�>��4<�~?y?�>3G?u�T?b^\?"K?�: >�w�����/�X��F���뽰b�=s�*>��^�c�ڽ��N�'=4⟽��-���S<�=��߽�*s��n=�_�>��s>4
��?�0>v�ľP��G�@>M����O���ي��:��ٷ=���>:�?���>gZ#�ȴ�=@��>I�>����6(?�?�?��!;�b�e�ھ��K�4�>�B?	��=��l�l���K�u�uh=��m?=�^?��W�'��T�b?��]?Kh�=���þҶb�щ�j�O?�
?��G�	�>��~?C�q?��>�e�:n�'��Db�A�j��Ѷ=Rr�>iX�T�d��?�>{�7?�N�>`�b>�$�=eu۾�w��q��c?}�?�?���?�**>~�n�R4�t_�������rK?%�?=�¾ӥ?�TN=>���a,w��m��f���ӾW����|m�
���Y��ML�c�����=!?�Jv?���?��J?!�#^���d�!Vs�Ӡd�J���� �վ$���R���/��e�h�	�,���_�D�\�����;B��ڴ?+i(?&4�?��>����[���˾�K@>����A��+�=p��ar<=��\=��h�Es/�I��V�?�;�>���>tD<?�Z�a>�F2�ֱ7������+>���>t��>�(�>�,�:OE/�����Cʾ�����ֽH�v>�c?�_L?�zn?Y����0��ނ��@"���5�"�����F>8�>M>�Q����?%��W=�� s��r�%㐾�	��|=B�1?�ւ>���>�?a~?~�	�լ����t���1��y�<wB�>xj?�U�>0��>�,н'!�f��>��l?x��>< �>M���;K!��{��ʽ#<�>�߭>���>��o>޷,��'\�bg��;���d9���=2�h?Er���*a����>�R?��b:�	H<υ�><�v���!����!�'�g!>4�?�Ū=e�;>�sž�"�B�{����0�!?�?�>瓜�T��f֗>��?�n�>�<�>��?�o}>�[;<��<I8?�^?X'H?r�D? &�>��v=�O��N�۽���(�N=:Z�>�B>[X<��>ˡ���4��ZQ����=O'>����Hp�@"+<"������<�Q=��>��ڿ��J�� ־� �u��b�	�)�����ý�F���b	�㸾����h*w����$5��VW�]qa������p��m�?O�?�����D��<ޙ�+C���������>YG}��ŉ������2��R���ྫྷ﮾Q�"�S���i��Pe�]?�����տ�ι�u�a�h�>d{�>�_�?)�&�P��քK��>�oR�Ľ�H��姚��:Ͽ����u?��>"�Ӿ���J�>��#>&>���>�k� ,=� >g/�>s0�>U�,?@*�< ƿ:t׿�>!S�?p 	@e|A?r�(�i��SCV=p��>%�	?��?>�V1��E�E����P�>;�?)��?3�M=��W�|�	�I~e?z�<=�F�o�ݻ��=�M�=�m=���7�J>`Q�>���iSA�LJܽ��4>�م>m�"�����~^��˾<��]>W�ս^=��3Մ?1{\��f���/��T��U>��T?�*�>y:�=��,?Y7H�^}Ͽ	�\��*a?�0�?���?"�(?3ۿ��ؚ>��ܾ��M?bD6?���>�d&��t����=�6�㉤�����&V����=R��>g�>��,�ً���O�eJ��I��=�{�����.쾀��G�A�[�ɽo���o���>�9���\>����RC�� p�<���j�=oi�>e�>h��>o�m>>nM?��W?�;�>3q�=�������y�ƾ�h+�;�쾭�= Σ�rF��B�%����	��`�R��߾�í����)�>��C�\��ԑ�����;�W�2?�(2�����k��=}	����<�a�o��;��=O���q�\L�?�-?`��,'o�KTʾo]=P&|���l?e���-�]ę���o>u�	��9���>�k>�	̾�'4�xT�$l0?�I?m���EJ���_*>$� ��-=��+?�?��X<*�>}L%?��*�O��ā[>��3>�ݣ>��>N%	>i���=۽�?�|T?;�������>@T���z�JK`=WO>%5��A꼾�[>Ӎ�<J����U����+/�<RW?��>��)����e�����==�x?�?�-�>�zk?&�B?v�<gr����S�� �2|w=<�W?L%i?$�>Y큽
оEs����5?��e?��N>-ah�=�龮�.�0Q�&(?��n?�^?gm���n}�������u6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>��������%>�V��D�?��?Qlھ�̤�"���j�`�̾I>���R��u9>�e��O�Ⱦ%<1��7���kþ�A�=Y��>�}@�ל=�\>��2��.鿆Ry����|嗾��?��?���<]���6�|��^���6��J�A径O�>��>�a���䘾r�z��?�[��l�>h�E����>f�C��n��[������>� �>��}>sҽ�r��q�?8�����Ͽ�̠������U?ZA�?�1�?�i?h͟;��l��%a��4%���A?�]r?R%\?J��f�a�i�Y��Ȃ?�U�$
t�R�F�/:0��:��4?,�?p��`�=b�>s7�>���=3t�d�˿�Oп�t���?�`�?���S�>>�?Q�[?ߘE�ޮ�����HY��;�:#."?v��>��	�M�6�G������(?\?����:�[�_?/�a�M�p���-���ƽ�ۡ>��0��e\��M�����Xe����@y����?L^�?h�?Ե�� #�i6%?�>g����8Ǿ�<���>�(�>�)N>�H_���u>����:�i	>���?�~�?Pj?���������U>�}?U$�>��?2o�=�a�>�c�=H񰾸-��k#>�"�=��>��?��M?�K�>W�=��8��/�>[F��GR�Z$�=�C��>�a?�L?lKb>���2��!��uͽ�c1��O鼄W@�Ԛ,���߽7(5>��=>�>I�D��ӾW�?�o�A�ؿj���o'�54?��>��?���"�t�)���;_?�y�>�6�	,��#&���C�`��?�G�?��?>�׾QE̼.>��>�H�>r�Խ& �������7>f�B?- �FD���o�g�>t��?�@�ծ? i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?pQo���i�B>��?"������L��f?�
@u@a�^?*Hfѿ���IP��]y���P�=ᄦ=7>�A��d �=�w=p�Č��>}�>	{>��y>|6z>�bX>\�;>J���H"��B��$֓�W�?���-f�
�n�\g���b��		������&ʾ�����e۽Z����z%���ག<��6#�=��U?�R?�(o?� ?�i��>�����g=J�!�^̓=��>ʬ1??M?w�*?o�="M���~d�Po��ˏ���1���.�>��G>���>���>=A�>�\�;�EP>��C>��>$&>6f=9p���=�M>n��>���>fI�>*R�>�0d>�`��(z��i�>�I�����j�Ģ?�y��,l�L&d�!¤�u��A ��_?-�@>�񖿓Gڿ.����9F?�����8�	�0��L>��U?�R?�FO>'�p�n�>��Ӽdq���-�gW>��n�h�7�&)3�<N{>ʊ%?e�f>��u>{3��U8�x�P�%^��ע|>N&6?s����'9�T�u���H�>�ݾnM>���>��E�%e�� �4�i�\
|=�q:?�e?&ɲ�k���{�u������R>߇\>��=<H�=�=M>�[d��iƽ��G�!�0=8G�=�^>�?��+>���=!ɣ>b���N�E�>��B>H�->�??4�$?����L������Kx-��3w>&9�>d�>Z�>�J�'l�=J��>G�a>Nv
�Z���h���w?� W>���6_�r�n���|=�@���G�=�F�=O� ��s<� *=�~?���#䈿���e���lD?`+? �=N�F<��"�@ ���H��;�?l�@m�?��	�բV�;�?�@�?����=*}�>)׫>�ξ��L�ͱ?N�Ž1Ǣ�Δ	�y)#�aS�?��?j�/�Pʋ�l�z6>�^%?��Ӿtg�>�t��Y����j�u�ּ#=���>I8H?�S����O�s>��v
?b?�^򾂩��1�ȿA{v�3��>	�?v��?!�m��A��g@�)�>s��?>gY?mi>ng۾"aZ�1��>�@?�R?��>q8�*�'�t�?y޶?��?�[>�l�?��y?���>_o��u�3�?B��F������=�9�W��>�d>�b��b�;�I���Z���}f�ȭ���H>{V=�R�>����ƾ��=+���iܶ���½sݪ>�&�>�P�>l�>̅?N��>hO�>Ǽ�<���s‾���v�K?���?	���2n�+Q�<�=u�^��&?rI4?�j[�P�Ͼ�ը>�\?y?�[?d�>��M>��H迿9~�����<	�K> 4�>�H�>=$��GK>v�Ծc4D��p�>�ϗ>�����?ھ&-���G��9B�>�e!?ғ�>6Ӯ=�}?{+$?�Ay>�W�>2�D�N{����H���>3��>&�?ڋ?�"?i�ƾ��6�]����5����\���2>`?s?�P#?P��>~ّ�L��@��;��g�� ��pm�?f0^?�q�=#?2��?s�;?kE9?z�i>����Ͼd༽�Dr>��!?DR�k�A�~<&�h��w?�N?$��>�����ֽZ�׼M���Z���?�$\?�H&?��ca�/�¾3��<�#���Q����;qF�[z>ʋ>�v����=�>{ٰ=��l�G=6�5�h<Dp�=�h�>�=�7����0=,?ÿG�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>$�l���K���ڙ���F��_�Ž�\,�+(?T+�>=��>_,�>�2>�~�>�l��#H��Ӿo})�=�w�ݱ$�,�!�a��������2�Z�s!�x��4�ҽ$q�>Ǒ���>� ?d�E>w��>��?�ie=�b�>M�g> l>�"�>ʦ�>��a>i4�>� <c�ýAR?J^����'�<�:��[>B?�d?���>2|f��u��d��{e?dx�?Tk�?�^v>�Qh�3+�Qh?c��>o��XI
?�<=e��uɇ<�%��>�����\��m�>�xؽQ	:��M�H@f��d
?�G?Dݍ���̾vR׽]�����>�(�?�g?�(���d�B�k���j�Lb�^�_���9�Xb�H�J�ͥW��#��O��!A��j�M�"Ω�r<O?:}?[����-��}׾�=��\kO���>��>B�&>�<?r��>S�2��>�EP.�����ԡ�� �>1�Z?f��>:G?��;?X^N?�L?w��>��>�l����>�.�<�u�>Q_�>9�;?<�.?��4?S�?^�-?n�`>���v��u,׾B�?-�?Z?�D?'�?����\M���B���gP�	!��3���ˏW=���<g�޽��p����=��X>�K?^���8�����9dk>�e7?Q��>���>�����R�����<��>�
?�g�>G���=Pr��L��]�>U��?	_���=��)>S�=8҅��:��"�=�7��
�=~넼�K:�o#<�=J�=�Eu��g�)�:��;خ<�i�>��?���>�<�>�C��� �����c�=,Y>�!S>�#>�@پ|��}$���g�zGy>	u�?w�?��f=�"�=�K�=����K�����{�S]�<f�?-A#?4PT?ݓ�?z�=?�n#?S�>O(��I���[��T���?-?�ˑ>�(���̾18��܊3��%?��?�d`����)�:-���&ֽ��>�;0�����ޯ��B�
�;���^��E^�?���?�.Y�H\7����͘����גB?P��>7b�>"*�>�)��,h��#�r�<>h��>�&Q?�u�>��_?	O�?D�N?�e=���Ǹ�����S��5�<�=^?���?��?���?Zr�>`�g>濿��!�t(�]����+����G�G����>v�?Ⱥ�>?)?Y⽻]۸=k$�<$�ƾ�l>�<�>C�>?]�t>bX?�:[>,����G?_��>�Z�����餾=Ã���<�Y�u?��?;�+?�P=&��s�E�XF��0J�>Jn�?��?�2*?��S�b��=��ּSᶾ��q�s#�>�ٹ>O2�>�ʓ=~�F=�c>��>0��>t&��a��p8�=WM���?�F?B��=0ſsKr�|�&�9ƃ�
[������ǅ�t���~z��j��=Rɸ��Ԓ��¾���w��{��+���ʴ��;M���>�,�<��o=�%8>�D=��"=�+#<��R��T5>-�t������M��K.>I_Y���ý���>�y:�,�r+Ⱦj�?��E?��?u "?�>ֶ^>.=��t5�>��<Qh?=�=���ྯ�N�x���Bf�XJ��_EԾv:Y�:����=`l��v=��C>e�>Q
�;*�=�ӧ=��Z>W
2>$ >�H^<ܲ�<��=�	4>r^>}6j>�6w?X�������4Q��Z罥�:?�8�>c{�=��ƾq@?~�>>�2������yb��-?���?�T�?>�?=ti��d�>M���㎽�q�=L����=2>o��=x�2�T��>��J>���K��E����4�?��@��??�ዿТϿ6a/>�t7>=�>N�R��z1��|\�ɜb�_iZ�a�!?X/;��P̾k�>̺�=�#߾�oƾщ.=J�6>��b=�=��J\�0ʙ=�{��;=�3l=tǉ>��C>Q��=�+���n�=��H=��=��O>����p7��?,��!3=��=N�b><&>'4�>4?�*5?H�^?Iq�>��ٽR��G䙾�o>�v>	��>���=
��>'��>�L?��=?��[?��>��a��3�>��a>�W;��S��]��䴃�a�2>+[�?pr�?���>��ҽ�KS��.#�&�X�U-0���?:6?��?=��>����ٿ���tc�-���Ґ;��u�}X����|k��94���_���<�?�>���>�v�>b��>H�]>�T>�q�>ؽ�=��A<6@�=a�O=��*=aN���=���sS�=�����x9<���=P����)<jnX=�=aM��]��<��=�Y�>3?>4��>�ݏ=⳾\�1>����E#L�풽=����U�B�d�A~��+/���7�c>>�)U>�6���^���p?�lZ>�7=>m�?�u?HI!>�q
��Ҿ�Ν� �e�d�S��h�=߫>�25���9�l�^��)N��sҾq�>�F�>�A�>�I_>t�C��L�g�=�W��,� ��>4잾�Hc�҉,��p��i]��0Q��A�z����=�$?����$DQ>4{y?�9R?ˁd?�?�qV=����'>��w�<!A�h$/�_n���6����7?�JP?Lξ>-9�v`�� ¾�ˍ�3��>bhh��N���9t6�۟C��ľf��>	Е�9�ɾ,�<�&_���+���C�%���_��>�`F?8��?a*[��؅�:_��a�T�����>ڍr?�ņ>��>�?M����ސ�[!�=��r?Wo�?Fػ?�.�=)<�=�{�����>��?.Ζ?���?��o?g��'y�>���<U�>Kc��Q�=�>(��=�>u�?�		??i+���?�=T뾪�뾲/r��ż�l=-��>�3�>��9>���=햗=N�=Il>Vݐ>��>��T>k�>Q��>;�p�Cn�ݠ�>�j>b�"�s+?���>�O�;M�=>��9=��<�i�֢��ٽ�`�W/��'a���>;�>�f�>eݿ�GT?J?��%�	?-���l�C���>�^�=�7��1��>��u>�9�>���>�q�>�{R=��0>�ݫ>��Ҿ�>���[�!�(C�NpR���Ѿ1�z>�&�������:�I�2���6\���i�>5���G=�H�</>�?����k���)�x��J�?�e�>�6?㜌�����z>���>Z�>w�������΍�
Z���?���?�2c>C�>^�W?n�?ڔ1��3�{uZ�Ưu��'A�me�.�`��፿����l�
�"
��p�_?I�x?yA?
H�<�9z>o��?��%�=я�q(�>U/�9&;��0<=�.�>p,��@�`�ȯӾ��þ�0�3GF>��o?R&�?cX?�SV�i�6�U;�=N�?�f?P�i?�B?�i ?�Կ=��7?(�4>� ?�?�N?�k*?�}@?<݌>�ܿ>-W>y�p����|�4��8c�f�˽5���]��=Z[>	:ʽ�pA=>�e��:>����&��=<��=�g��|���W>��=���>�]?�[�>~�>�7?o���;8�5����S/?PX;=Dv���0��"��,�@�>I�j?��?c=Z?Q�c>5�A�&+C�� >�.�>��%>C\>]�>\aｭZE�[J�=f>�.>6��=yO��݁�5�	�7���(�<�>,��>R|>������'>툣�/z�U�d>a�Q�������S�T�G�k�1�,�v�FY�><�K?�?���=�\���Ef�N4)?c<?�JM?�?��=�۾��9�L�J�_�w�>GE�<���ﾢ�6#����:�T�:��s>�7��fޟ��b>�����߾�;n�_eJ� V��R=�#�8FK=z���	վF������=*�	>�]��n� �t>���ު��bJ?K5j=����IV������>�>)S�>��?���x��Y@����=��=Ɨ�>�<>Bs��TﾆkG��1��>��F? Wd?G�?����	�s�woL����u����f���?��>r�?��B>]�X=B���h\�Z�e��'D�u��>���>����KH��Þ�6��~'�3�u>:o�> �<>=�?2N?`�?
�a?RW'?#(�>��>ҥ½u�ľy4&?��?�=�KԽ~KT���8�@(F����>b)?�B�ԗ>(�?,�? '?e�Q?�?"T>?� ��\@�~m�>U�>@�W�VK��5�`>�J?w�>�ZY?�؃?vd>>��5����𺪽��=	�>��2?sB#?H�?Tθ>�>�������>�!�?��?��?6��>l�
?�K�>�i�>��4<�~?y?�>3G?u�T?b^\?"K?�: >�w�����/�X��F���뽰b�=s�*>��^�c�ڽ��N�'=4⟽��-���S<�=��߽�*s��n=�_�>��s>4
��?�0>v�ľP��G�@>M����O���ي��:��ٷ=���>:�?���>gZ#�ȴ�=@��>I�>����6(?�?�?��!;�b�e�ھ��K�4�>�B?	��=��l�l���K�u�uh=��m?=�^?��W�'��T�b?��]?Kh�=���þҶb�щ�j�O?�
?��G�	�>��~?C�q?��>�e�:n�'��Db�A�j��Ѷ=Rr�>iX�T�d��?�>{�7?�N�>`�b>�$�=eu۾�w��q��c?}�?�?���?�**>~�n�R4�t_�������rK?%�?=�¾ӥ?�TN=>���a,w��m��f���ӾW����|m�
���Y��ML�c�����=!?�Jv?���?��J?!�#^���d�!Vs�Ӡd�J���� �վ$���R���/��e�h�	�,���_�D�\�����;B��ڴ?+i(?&4�?��>����[���˾�K@>����A��+�=p��ar<=��\=��h�Es/�I��V�?�;�>���>tD<?�Z�a>�F2�ֱ7������+>���>t��>�(�>�,�:OE/�����Cʾ�����ֽH�v>�c?�_L?�zn?Y����0��ނ��@"���5�"�����F>8�>M>�Q����?%��W=�� s��r�%㐾�	��|=B�1?�ւ>���>�?a~?~�	�լ����t���1��y�<wB�>xj?�U�>0��>�,н'!�f��>��l?x��>< �>M���;K!��{��ʽ#<�>�߭>���>��o>޷,��'\�bg��;���d9���=2�h?Er���*a����>�R?��b:�	H<υ�><�v���!����!�'�g!>4�?�Ū=e�;>�sž�"�B�{����0�!?�?�>瓜�T��f֗>��?�n�>�<�>��?�o}>�[;<��<I8?�^?X'H?r�D? &�>��v=�O��N�۽���(�N=:Z�>�B>[X<��>ˡ���4��ZQ����=O'>����Hp�@"+<"������<�Q=��>��ڿ��J�� ־� �u��b�	�)�����ý�F���b	�㸾����h*w����$5��VW�]qa������p��m�?O�?�����D��<ޙ�+C���������>YG}��ŉ������2��R���ྫྷ﮾Q�"�S���i��Pe�]?�����տ�ι�u�a�h�>d{�>�_�?)�&�P��քK��>�oR�Ľ�H��姚��:Ͽ����u?��>"�Ӿ���J�>��#>&>���>�k� ,=� >g/�>s0�>U�,?@*�< ƿ:t׿�>!S�?p 	@e|A?r�(�i��SCV=p��>%�	?��?>�V1��E�E����P�>;�?)��?3�M=��W�|�	�I~e?z�<=�F�o�ݻ��=�M�=�m=���7�J>`Q�>���iSA�LJܽ��4>�م>m�"�����~^��˾<��]>W�ս^=��3Մ?1{\��f���/��T��U>��T?�*�>y:�=��,?Y7H�^}Ͽ	�\��*a?�0�?���?"�(?3ۿ��ؚ>��ܾ��M?bD6?���>�d&��t����=�6�㉤�����&V����=R��>g�>��,�ً���O�eJ��I��=�{�����.쾀��G�A�[�ɽo���o���>�9���\>����RC�� p�<���j�=oi�>e�>h��>o�m>>nM?��W?�;�>3q�=�������y�ƾ�h+�;�쾭�= Σ�rF��B�%����	��`�R��߾�í����)�>��C�\��ԑ�����;�W�2?�(2�����k��=}	����<�a�o��;��=O���q�\L�?�-?`��,'o�KTʾo]=P&|���l?e���-�]ę���o>u�	��9���>�k>�	̾�'4�xT�$l0?�I?m���EJ���_*>$� ��-=��+?�?��X<*�>}L%?��*�O��ā[>��3>�ݣ>��>N%	>i���=۽�?�|T?;�������>@T���z�JK`=WO>%5��A꼾�[>Ӎ�<J����U����+/�<RW?��>��)����e�����==�x?�?�-�>�zk?&�B?v�<gr����S�� �2|w=<�W?L%i?$�>Y큽
оEs����5?��e?��N>-ah�=�龮�.�0Q�&(?��n?�^?gm���n}�������u6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>��������%>�V��D�?��?Qlھ�̤�"���j�`�̾I>���R��u9>�e��O�Ⱦ%<1��7���kþ�A�=Y��>�}@�ל=�\>��2��.鿆Ry����|嗾��?��?���<]���6�|��^���6��J�A径O�>��>�a���䘾r�z��?�[��l�>h�E����>f�C��n��[������>� �>��}>sҽ�r��q�?8�����Ͽ�̠������U?ZA�?�1�?�i?h͟;��l��%a��4%���A?�]r?R%\?J��f�a�i�Y��Ȃ?�U�$
t�R�F�/:0��:��4?,�?p��`�=b�>s7�>���=3t�d�˿�Oп�t���?�`�?���S�>>�?Q�[?ߘE�ޮ�����HY��;�:#."?v��>��	�M�6�G������(?\?����:�[�_?/�a�M�p���-���ƽ�ۡ>��0��e\��M�����Xe����@y����?L^�?h�?Ե�� #�i6%?�>g����8Ǿ�<���>�(�>�)N>�H_���u>����:�i	>���?�~�?Pj?���������U>�}?U$�>��?2o�=�a�>�c�=H񰾸-��k#>�"�=��>��?��M?�K�>W�=��8��/�>[F��GR�Z$�=�C��>�a?�L?lKb>���2��!��uͽ�c1��O鼄W@�Ԛ,���߽7(5>��=>�>I�D��ӾW�?�o�A�ؿj���o'�54?��>��?���"�t�)���;_?�y�>�6�	,��#&���C�`��?�G�?��?>�׾QE̼.>��>�H�>r�Խ& �������7>f�B?- �FD���o�g�>t��?�@�ծ? i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?pQo���i�B>��?"������L��f?�
@u@a�^?*Hfѿ���IP��]y���P�=ᄦ=7>�A��d �=�w=p�Č��>}�>	{>��y>|6z>�bX>\�;>J���H"��B��$֓�W�?���-f�
�n�\g���b��		������&ʾ�����e۽Z����z%���ག<��6#�=��U?�R?�(o?� ?�i��>�����g=J�!�^̓=��>ʬ1??M?w�*?o�="M���~d�Po��ˏ���1���.�>��G>���>���>=A�>�\�;�EP>��C>��>$&>6f=9p���=�M>n��>���>fI�>*R�>�0d>�`��(z��i�>�I�����j�Ģ?�y��,l�L&d�!¤�u��A ��_?-�@>�񖿓Gڿ.����9F?�����8�	�0��L>��U?�R?�FO>'�p�n�>��Ӽdq���-�gW>��n�h�7�&)3�<N{>ʊ%?e�f>��u>{3��U8�x�P�%^��ע|>N&6?s����'9�T�u���H�>�ݾnM>���>��E�%e�� �4�i�\
|=�q:?�e?&ɲ�k���{�u������R>߇\>��=<H�=�=M>�[d��iƽ��G�!�0=8G�=�^>�?��+>���=!ɣ>b���N�E�>��B>H�->�??4�$?����L������Kx-��3w>&9�>d�>Z�>�J�'l�=J��>G�a>Nv
�Z���h���w?� W>���6_�r�n���|=�@���G�=�F�=O� ��s<� *=�~?���#䈿���e���lD?`+? �=N�F<��"�@ ���H��;�?l�@m�?��	�բV�;�?�@�?����=*}�>)׫>�ξ��L�ͱ?N�Ž1Ǣ�Δ	�y)#�aS�?��?j�/�Pʋ�l�z6>�^%?��Ӿtg�>�t��Y����j�u�ּ#=���>I8H?�S����O�s>��v
?b?�^򾂩��1�ȿA{v�3��>	�?v��?!�m��A��g@�)�>s��?>gY?mi>ng۾"aZ�1��>�@?�R?��>q8�*�'�t�?y޶?��?�[>�l�?��y?���>_o��u�3�?B��F������=�9�W��>�d>�b��b�;�I���Z���}f�ȭ���H>{V=�R�>����ƾ��=+���iܶ���½sݪ>�&�>�P�>l�>̅?N��>hO�>Ǽ�<���s‾���v�K?���?	���2n�+Q�<�=u�^��&?rI4?�j[�P�Ͼ�ը>�\?y?�[?d�>��M>��H迿9~�����<	�K> 4�>�H�>=$��GK>v�Ծc4D��p�>�ϗ>�����?ھ&-���G��9B�>�e!?ғ�>6Ӯ=�}?{+$?�Ay>�W�>2�D�N{����H���>3��>&�?ڋ?�"?i�ƾ��6�]����5����\���2>`?s?�P#?P��>~ّ�L��@��;��g�� ��pm�?f0^?�q�=#?2��?s�;?kE9?z�i>����Ͼd༽�Dr>��!?DR�k�A�~<&�h��w?�N?$��>�����ֽZ�׼M���Z���?�$\?�H&?��ca�/�¾3��<�#���Q����;qF�[z>ʋ>�v����=�>{ٰ=��l�G=6�5�h<Dp�=�h�>�=�7����0=,?ÿG�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>$�l���K���ڙ���F��_�Ž�\,�+(?T+�>=��>_,�>�2>�~�>�l��#H��Ӿo})�=�w�ݱ$�,�!�a��������2�Z�s!�x��4�ҽ$q�>Ǒ���>� ?d�E>w��>��?�ie=�b�>M�g> l>�"�>ʦ�>��a>i4�>� <c�ýAR?J^����'�<�:��[>B?�d?���>2|f��u��d��{e?dx�?Tk�?�^v>�Qh�3+�Qh?c��>o��XI
?�<=e��uɇ<�%��>�����\��m�>�xؽQ	:��M�H@f��d
?�G?Dݍ���̾vR׽]�����>�(�?�g?�(���d�B�k���j�Lb�^�_���9�Xb�H�J�ͥW��#��O��!A��j�M�"Ω�r<O?:}?[����-��}׾�=��\kO���>��>B�&>�<?r��>S�2��>�EP.�����ԡ�� �>1�Z?f��>:G?��;?X^N?�L?w��>��>�l����>�.�<�u�>Q_�>9�;?<�.?��4?S�?^�-?n�`>���v��u,׾B�?-�?Z?�D?'�?����\M���B���gP�	!��3���ˏW=���<g�޽��p����=��X>�K?^���8�����9dk>�e7?Q��>���>�����R�����<��>�
?�g�>G���=Pr��L��]�>U��?	_���=��)>S�=8҅��:��"�=�7��
�=~넼�K:�o#<�=J�=�Eu��g�)�:��;خ<�i�>��?���>�<�>�C��� �����c�=,Y>�!S>�#>�@پ|��}$���g�zGy>	u�?w�?��f=�"�=�K�=����K�����{�S]�<f�?-A#?4PT?ݓ�?z�=?�n#?S�>O(��I���[��T���?-?�ˑ>�(���̾18��܊3��%?��?�d`����)�:-���&ֽ��>�;0�����ޯ��B�
�;���^��E^�?���?�.Y�H\7����͘����גB?P��>7b�>"*�>�)��,h��#�r�<>h��>�&Q?�u�>��_?	O�?D�N?�e=���Ǹ�����S��5�<�=^?���?��?���?Zr�>`�g>濿��!�t(�]����+����G�G����>v�?Ⱥ�>?)?Y⽻]۸=k$�<$�ƾ�l>�<�>C�>?]�t>bX?�:[>,����G?_��>�Z�����餾=Ã���<�Y�u?��?;�+?�P=&��s�E�XF��0J�>Jn�?��?�2*?��S�b��=��ּSᶾ��q�s#�>�ٹ>O2�>�ʓ=~�F=�c>��>0��>t&��a��p8�=WM���?�F?B��=0ſsKr�|�&�9ƃ�
[������ǅ�t���~z��j��=Rɸ��Ԓ��¾���w��{��+���ʴ��;M���>�,�<��o=�%8>�D=��"=�+#<��R��T5>-�t������M��K.>I_Y���ý���>�y:�,�r+Ⱦj�?��E?��?u "?�>ֶ^>.=��t5�>��<Qh?=�=���ྯ�N�x���Bf�XJ��_EԾv:Y�:����=`l��v=��C>e�>Q
�;*�=�ӧ=��Z>W
2>$ >�H^<ܲ�<��=�	4>r^>}6j>�6w?X�������4Q��Z罥�:?�8�>c{�=��ƾq@?~�>>�2������yb��-?���?�T�?>�?=ti��d�>M���㎽�q�=L����=2>o��=x�2�T��>��J>���K��E����4�?��@��??�ዿТϿ6a/>�t7>=�>N�R��z1��|\�ɜb�_iZ�a�!?X/;��P̾k�>̺�=�#߾�oƾщ.=J�6>��b=�=��J\�0ʙ=�{��;=�3l=tǉ>��C>Q��=�+���n�=��H=��=��O>����p7��?,��!3=��=N�b><&>'4�>4?�*5?H�^?Iq�>��ٽR��G䙾�o>�v>	��>���=
��>'��>�L?��=?��[?��>��a��3�>��a>�W;��S��]��䴃�a�2>+[�?pr�?���>��ҽ�KS��.#�&�X�U-0���?:6?��?=��>����ٿ���tc�-���Ґ;��u�}X����|k��94���_���<�?�>���>�v�>b��>H�]>�T>�q�>ؽ�=��A<6@�=a�O=��*=aN���=���sS�=�����x9<���=P����)<jnX=�=aM��]��<��=�Y�>3?>4��>�ݏ=⳾\�1>����E#L�풽=����U�B�d�A~��+/���7�c>>�)U>�6���^���p?�lZ>�7=>m�?�u?HI!>�q
��Ҿ�Ν� �e�d�S��h�=߫>�25���9�l�^��)N��sҾq�>�F�>�A�>�I_>t�C��L�g�=�W��,� ��>4잾�Hc�҉,��p��i]��0Q��A�z����=�$?����$DQ>4{y?�9R?ˁd?�?�qV=����'>��w�<!A�h$/�_n���6����7?�JP?Lξ>-9�v`�� ¾�ˍ�3��>bhh��N���9t6�۟C��ľf��>	Е�9�ɾ,�<�&_���+���C�%���_��>�`F?8��?a*[��؅�:_��a�T�����>ڍr?�ņ>��>�?M����ސ�[!�=��r?Wo�?Fػ?�.�=)<�=�{�����>��?.Ζ?���?��o?g��'y�>���<U�>Kc��Q�=�>(��=�>u�?�		??i+���?�=T뾪�뾲/r��ż�l=-��>�3�>��9>���=햗=N�=Il>Vݐ>��>��T>k�>Q��>;�p�Cn�ݠ�>�j>b�"�s+?���>�O�;M�=>��9=��<�i�֢��ٽ�`�W/��'a���>;�>�f�>eݿ�GT?J?��%�	?-���l�C���>�^�=�7��1��>��u>�9�>���>�q�>�{R=��0>�ݫ>��Ҿ�>���[�!�(C�NpR���Ѿ1�z>�&�������:�I�2���6\���i�>5���G=�H�</>�?����k���)�x��J�?�e�>�6?㜌�����z>���>Z�>w�������΍�
Z���?���?�2c>C�>^�W?n�?ڔ1��3�{uZ�Ưu��'A�me�.�`��፿����l�
�"
��p�_?I�x?yA?
H�<�9z>o��?��%�=я�q(�>U/�9&;��0<=�.�>p,��@�`�ȯӾ��þ�0�3GF>��o?R&�?cX?�SV�i�6�U;�=N�?�f?P�i?�B?�i ?�Կ=��7?(�4>� ?�?�N?�k*?�}@?<݌>�ܿ>-W>y�p����|�4��8c�f�˽5���]��=Z[>	:ʽ�pA=>�e��:>����&��=<��=�g��|���W>��=���>�]?�[�>~�>�7?o���;8�5����S/?PX;=Dv���0��"��,�@�>I�j?��?c=Z?Q�c>5�A�&+C�� >�.�>��%>C\>]�>\aｭZE�[J�=f>�.>6��=yO��݁�5�	�7���(�<�>,��>R|>������'>툣�/z�U�d>a�Q�������S�T�G�k�1�,�v�FY�><�K?�?���=�\���Ef�N4)?c<?�JM?�?��=�۾��9�L�J�_�w�>GE�<���ﾢ�6#����:�T�:��s>�7��W-���g>��
���۾�=n�nGJ�<)뾟�,=����;=�
���Ծ�|�d:�=Q>OQ��T!�햿G�����H?���= E��=�_�N���D>48�>��>�P"��{u��6?��D��	�=h��>[�8>�WT��v𾠔H����6��>��??��Y?S��?��y�� ��4���@��M�;=f�>�?�5?��>�C>�݄�Tk��Pn��o�]��>�?�g�R�J��+x�%��0{`���_>a�>��	�	?fsA?G�@?��a?��)?J��>x�;>�*��o����?�k�?��=�m��!���5)�'�H�{��>j��>�`����>��9?|�B?-uS?�kb?��?�C>
���-�Q�a>c��>��@��q���+ >J�q?���>u�?c��?uہ>��Љؾ�-��J�>�"q>��.?��g?�y??��?GG�>b���>�H�"��>_?��?�l�?�+�=��?��/>��>�O�>t;�>��>7)?��D?�v?��K?���>��Ỻ�2�w���Q����ׄ�O;�X=>d��Y8�<��>z�ν7B�E�8���A;,�ͽe �m�d= �?��u�=��>Yt>!��g�0>
�ľ�È�	B>Ӡ�ٕ��.w���:��L�=�^�>��?a��>��"��P�=��>3Y�>�v��$(?�,?�?(�:�Eb��ھ9�L��а>>gA?���=Ûl�b���4�u�2�h=P�m?�'^?��U�^���#Yc?��^?�󾋸;��V˾�j�@��n�I?�/?mH��3�>�V{?Sq?t:�>�Ml�_ui�U����b��H|�WԳ=��>.���ag���>ٜ5?c]�>nZW>!�=\ վ�u�-��� i?���?�&�?cz�?u�>� q��ݿY,�~R����Q?.��>��ʾ�=?���\��Hɛ��jԾ�L�Q��Hzƾ��ټ��5xD�����3o��5�=�?&Z�?r�?Y_i?����Q�G�@�=Ä�E~�(��?�	��y��W@���$��u��3�6����_@Ҿ����W���J"���?y�R?��ƽ���>��?�yH)��+�<�,=_�t�Ʈ�|~�<N��=�ӷ��¶��c��맾��侭�%?s�>qi?ӻI?�E�9Z$�>�6���-�*���=�i�>�f�>�_?z��>�E��q����	1̾��Ǿv�>��e?�B?S�X?��A���'������5]����">	e�=�e�>�?���J,����2���u�������'��c�>��M?P@�>*��>�ʩ??�(?},��>w��+f�H!��Χ��؋>A^}?��>�Q�>�FR=|d�8v�>��t?-��>qӀ>�q]��t'�X�f�9:;\�>��>�k?pH>����\X��%��?����3���>b�y?�j��	���>x�>?@&��=,��K>E_�����ξuмW<>ö�>52(�/U}>�������I�k��;��%?�,?F��O
�#��=�Y:?[%?P>@b}?���=�޾��M����>�\l?ߌB?@cQ?�*?�8z>$ ��ȧ�R���zN=��|>B��>�x�=�J=)'��)��H ���@>П=>bQ�=�;�=尲=y�v��l�=�K=|r>�@ۿ�K��vپ��dF�T
��a����������c	�Q����K��?Ax�����&��YU���b�2c���?l��d�?g+�??w���������xv��:����>��r��ς��@��L��y��
q�Z��W!��O���h��e�AiN?k����п�������?xo�>*Z?=6�#!W��\�[>qS� �ƾo#�Tŧ��wԿ�2���	f?�F�>U�ԾX��<�>
�5��k^>�dv>
!Ǿ(�=��z���>�R�>y��>�Z��߁ƿ>Wÿb}ʽ�Y�?�j�?SuA?�(�z���sW=���>�	?@>991� T�DӰ��+�>�7�?���?qgM=��W��$	��pe?j�<��F��^߻%�=�b�=��=ߛ�('J>�G�>�}�JqA���ܽ�~4>0�>>j"�����D^��w�<jO]>t�ս���3Մ?!{\��f���/��T��&U>��T?�*�>g:�=��,?_7H�]}Ͽ�\��*a?�0�?���?'�(?ۿ��ؚ>��ܾ��M?TD6?���>�d&��t�ޅ�=<6�%�������&V�l��=O��>m�>Ƃ,�ً���O�I��"��=�� �V�Ŀ���h"��Y9��J�V�7��ٌ�s���ò��J����|���ֽ2T=<p�=�X>f�f>ߞK>�u>EV?I
t?���>�	7>xm��P����ž@�\a��4$y�~𫾑q��_=����Ͼ�<��4��&q�2t�pa���g#�rv�=�zN�{��H�shg�;0L�� 0?���=��վ;�8�	9�=C���@�����g�ѥϽ�zھb(6��tj��0�?��4?�᏿?:X��E��*ϼ�-��۟d?�M9��������P�>\��,�`=\��>Ք�=ُ���"��@��@0?"U?���Z���{�*>� �:$=��+?�E?q&q<$(�>�$%?*�]s��R[>��3>sף>���>�G	>����ܽPV?�vT?t �.U����>PC��_�z���_=w�>��3�p�/�Z>dS�<��8^��ʏ�s2�<�X?��>�z-�I�M���X�A��=��{?W�?�ו>*ih?mD?iK��{�����R�N%���/=�
S?��e?�X>����34վb,���03?�qh?��P>^�g�:�۾�-�]���	?��n?��?�ܼ�}��Β�P�ݑ6?��v?�r^�vs�����L�V�v=�>\�>���>��9��k�>�>?�#��G������pY4�$Þ?��@���?A�;<��K��=�;?g\�>�O��>ƾ�z������B�q=�"�>���xev�����Q,�`�8?۠�?���>������[�Z>w"��zX�?Q�?}��Z_h�n���?�d�;�;{�<�=y��C���)�����4�WΔ���cE��)��Qs�>��@cT��p>�#�_ӿIWԿ���U򌾓9���>���>WF�:����x�4f�G�6�He��`�bͨ>b�>G泽}i���v�+(8��X�����>��1�Z�y>�'K�+�������x���ԋ>]:�>�΀>�h�����?���|п�3��?Z��RR?���?p�?��?�'߼�}���i����@?�q?�V?��t��!;�a//�>�y?������_���C��0Q�M�=� �>�>����1�:�r>��>�T��]\\�?I˿޲ҿ�R)��O�?��?���R��>� �?"5?�4�]q��tǱ�0��|�[�>vn?�ނ>��վA��������,ž�?'�L?E6*�s�-�]�_?*�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?ӵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�
i	>���?�~�?Qj?���� ����U>
�}?K��>B̄?�+�=���>�(�=������%>zo�=��/�ӯ?ՋM?@�>��=*P8�&�.���E���Q�����|C���>QLa?��K?�Jd>����L�9��� ��eν�$3�Ҳڼj<�"�+�FX�t�7>�:>O/>�E�N.Ҿ��?5p�*�ؿ�i��>p'�z54?	��>�?�����t�����;_?z�>7��+���%��C�R��?�G�?3�?��׾rR̼(>�>�I�>��Խ;���������7>7�B?]��D��f�o�v�>���?��@�ծ?Oi�<	?L��P��}`~�����7����=R�7?X/��z>���>w�=�nv�仪�>�s����>�A�?{�?4��>g�l?��o���B�k�1==K�>s�k?�s?��o���o�B>��?��������K�t f?�
@u@�^?��X�׿`���ƾ�6ʾ9�=��=��A>����Pa�=��7=�~�<�y�ɒX�><�>Z�>?�>��z>?">JV&>�}����c����2����C��&��;x�����YY���9���꿾'k�d ���H=�_G�

���F�#���w��=�R?C=Q?�r?�?���U%>����D�9J	�}�R=��>�1?�I?O(*?:��=���Bc��р��ѧ�������>��R>���>o��>r��>��}:��5>.r+>�:v>��>o.=$3�C%I=չ6>��> ~�>�8�>�p�>ެ�=�,��_��J�E�����5�@ͨ?z`����S��)�����Ε��u�K<��?WW�=s���ɿF"����G?~��v�+�6�:���A>��;?�M?�eR>ljD��ѹ���/=�?�i�0��*>>�Ͻ���;5/�u�y>< ?L�f>�tu>6�3��_8���P����� �{>c�5?¶�H09��u��H�\ݾXaM>Ћ�>�o>��o�����;�8ji�H|=�h:?d?R����İ��v�<V��3R>��\>p=x��=&�M>��b�C]ƽR�G�ݧ-=��=��^>&��>�(%>��=f=�>p!f��D�:�>�GV>�a�=j�C?��?`��:e;��������t�>���>���>��=*yN�Ry=m��>v}r>�����	�����֬)���2>�����|�����8{s=�љ�O*>��==�'���P����;�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�m�>!z�L[����_�u�\�#=D��>_;H?�P����O��>��w
?C?�a�����ȿf}v�%��>��?q��?A�m�8A���@��|�>
��?�eY?!gi>�[۾[bZ�U��>��@?�R?!�><:�̙'���?�ݶ?���?>"O>���?ҙo?���>�(����/�����'�����=�˾;�_�>��=&e���7C��d�����0j�v����U>�S=.}�>D8���Z�=x������<e��D�>F�x>;�K>[֝>�L?`��>�>7U=*������Ś��O�Q?9��?����-i��Z����}��R>?g2?ɱ=oʾw;�>Ղ{?x?��'?K��>��N��Ǌ���S��sC��S�>���>U�>��?;0/^>�/���փ� ��>av�>��O;������W�M�3>
-�>��?���>kt>*�!?�� ?;Oa>�c�>��C�����2H��j�>���>|�?4~?��?bpȾ��6��^���a��>�[�U7>��q?ޢ!?8d�>������,MB<��Q�`ʆ��4�?�+i?�V���?�ֈ?;9?�??D�v>M"��ݾ�V���u�>��!?���D�a�%����Q
?��	?��>�C��1���ql3��	�vr���~?��Z?��'?Dg���Z���ž(�=��ӻa(����;av�#>ߩ>U���C�=c+>���=�#j��5���<��=m@�>�N�=2�-�[ؗ�#=,?e�G�Bۃ�Y�=?�r�9xD���>�IL>`����^?�l=���{�����x���U�� �?��?Ck�?���-�h��$=?�?Q	?�"�>QK���}޾���Pw��~x��w���>���>]�l�\�H���Й���F����Žn�3��h?��>�{?m>?#{�=0�>~�.�f��r���r��$�[��:�a'�X-A�R�%������	�æ�;�����_u9>�}��?��>��?��a>{�>N�>͢�V�>�Î>N�`>�f~>�~�>S�=R��=��>�֫=JR?F�����'����<����3B?�sd?�*�>"�h����O��8}?0��?�q�?EBv>�wh�'+��o?�9�>f���r
?�:=z��=<S����#9��_�朎>�Y׽�:�PM�iqf�h
?h/?+����̾	Q׽0*���e=��?�5'?�����T�g5��H�^������n�������f=��N�Ef��߃���}��
Y��S����d?�U?��7��W>��F��*a��=�ǋ�>�} ?��>�D�>���>�rD���r��H�<O���a����> bv?�ߑ>��;?i`5?fNS?1�D?r>�@�>�pr�*<�>�h8>��>���>�b3?�#?��.?�i?�Y$?�)=>����)���(�Q�?��&?��4?<�>uY?�	D��]�ҁ�ׂ_�6d
���ض���ܩ=��7������=qSA>DU?����8�������j>Y�7?p��>���>�
��5-����<w�>!�
?�D�>O����ur�]��Z�>��?*
�ki=p�)>`��=�����2ۺ�b�=T¼D��=ḁ��S;�ĝ<?f�=�=�w�T���9�:�W�;s��<or�>?�?b��><C�>>��.� �G��!z�=Y>SS>>�Eپ�|��$����g��Vy>�v�?Pz�?��f==�=��=�~���U��������S��<u�?�J#?YWT?��?��=?�h#?��>J)��L���^��Q��#�?�R,?�
�>�/�&c˾�쨿�G3�MI?0?�`���U)��>¾ǥֽ&$>k�/�%�~�����C���e��������?j��?$�A��7�MV�A��������]C?���>O:�>$s�>N~)�*�g�����;>d��>�R?���>��P?.z?�9\?�3[>�9��������Wּ�? >G >?���?|̐?�{z?�>�>�>)l)��q��������Q�ڽ�酾�=RR>C��>6��>E�>a��=w̽y����;�VC�=/�j>��>�"�>�c�>�}>��	=�!C?	�>�rվf����e�7� X=4�]?
��?=S?��Jq�L�B�;V㾯��>_��?0��?��1?�fY�њ> ��;�!ɾ��{����>S��>���>Y�=b)>=|��=�>B�>�S2��I��4�ƍ�l?a�K?��!=��ſ��q��{p�.K��@Ce<������c��M��nZ����=&�0�����2\�&�����A����P���{��~�>]��=�U�=	�=*��<�>Ӽ'.�<V�E=���<J =��o�Y�t<�9����b��~�:�hwe<�SG=�B𻓋˾�}?W8I?"�+?w�C?��y>F>q�1����>�;��B8?'V>�P�T���z�;�K���� ���ؾ�S׾d�����>ҹI��>�3>K �=3�<�m�=�4s=���=}kG�E�=��=u��=�>�=?��=A�>�>�6w?V�������4Q��Z罦�:?�8�>V{�=��ƾk@?k�>>�2������vb��-?���?�T�?@�?Fti��d�>I���㎽�q�=R����=2>o��=s�2�S��>��J>���K��E����4�?��@��??�ዿ̢Ͽ.a/>9�<>Oa>�eT��=1���`��yX���L���?�8�l#Ѿ)N}>�ֲ=���ľ��:=�=>�Xu=E=��[��G�=]@n���=�Na=�8�>�E>�d�=/���L�=�"=���=�pK>�����m�¶3���6=;]�=�g>V| >h�>aE?�?B�F?=6�>�%�(����p���ǚ>(D>�>F�j=�n2>�=�>�@?!�C?�W?-y�>!�=̍�>9��>	�4��*g����i��,�\Me?q�r?��>�¼�hw��.���A��j��`�?L�/?�!?�>��K���4���L��ì�-�<�mZ=D�ؽQњ;�5���ɽ����潵O6>}G�><�>Cq>!��=�=D><U�>:��=�P<<K=�΋��p�7a_�
�>���=���<z������=n��='��2b'��;<RW�U��M�\�XV�=��>��>�u�>{o�=��Φ/>�d���L����=�~��5JB�W1b�݇|�{�/�y�8���?>�R>����X����?_�[>^pB>�P�?�jt?k�$>
��F�Ҿ|e���c�nO�#]�=��>K3��H:� �^���K��Ѿq��>��>���>��-> �)�V>[��*�^s���'�!q�>�p��^�:�eL
���a�p泿;�����Y�S���j7#?�F��j��>kh�?��L?��?a��>z>����_->>4�u��8��X��zc	>�:,?�X??(�ھ_WQ��]ɾ�������>LFF�6*M��\��&�0��!e�-+��p �>l[��w@ξ�G5��T��ꁏ���A�@W|�)�>��N?b]�?�����À�t{I����Rh��T�?5�c?�Z�>R�?@+?w���eT�󲁾&��=;)r?9��?j��?�a
>frh=u˦�m��>�?�q�?pm�?� d?a�����>��=ߵ>���ݣ]>�=��7>��[>a�?��(?��??�Ľn�!�7�Ծ7ࡾb��-n�l8>2��>�_W>��*�ǭ(�&�>���=�4F>�>��>��<0\+>�t�=Nx��n����?Һ\>E&M>}=�>�N>P�~=^�μ >>\�=xUA���������f��@S<H��b �=q$,>��?s?Կ=��?x��>��0�Z?Aǌ��,���`���N>�5�h+�>���=1A�>��
?�]?��= G�>�޻=ʗ���=���+��-�3N�s㾶E�>�:��"�]�*�S�����ľ�<��rk�]}��@O;���<�Њ?�� ��{l���(�c���;?k�>�f$?U�0�+@��eR=���>_�>|[ ��$��d���3���\�?���?�4e>a�>��Q?�?Ci5�l#�?|R�~�t��t=��c�{<a�R���/p���?�����`?ƴx?�B?�(�<��><��?��(�Ж��&N�>�,��09�4�/=�ݣ>�ݼ���j���ӾŁɾa[��A>�:n?q��?�S?0�a� �׽
�9��g,?��;??pX?dY2?��]?év���$?5>�G�>�	?�>4?}0?�-?�=m>��]>�Z�=�;�<o2��.>�L>Ž��e���<D=a�=-mȽH�<2e�=�ҧ������6�Y�	>ʮܽ��<�0�=;U�<��=�~�>/�r?u��>�ӑ=~�a?��>
!�"�;c�	?���>���>��1�w]#�L-��]�>�fY?[I�?�B�?���>�FF�Y%��/P>�z�>�@>%�>Qc�>�X��a���> ~�>���=�	>����J�߾�~��v���?w >�>���>�z>���� 1>�����{�|af>V�J�(q��"F�SZG�b�/��p�L[�>;<K?��?��=(6龠0��G_e�q&?B�;?K*N?���?�~=�CԾs�7�I	L�E� �?��>s��<��	�|䡿U��x�;�� :ibt>N(��W-���g>��
���۾�=n�nGJ�<)뾟�,=����;=�
���Ծ�|�d:�=Q>OQ��T!�햿G�����H?���= E��=�_�N���D>48�>��>�P"��{u��6?��D��	�=h��>[�8>�WT��v𾠔H����6��>��??��Y?S��?��y�� ��4���@��M�;=f�>�?�5?��>�C>�݄�Tk��Pn��o�]��>�?�g�R�J��+x�%��0{`���_>a�>��	�	?fsA?G�@?��a?��)?J��>x�;>�*��o����?�k�?��=�m��!���5)�'�H�{��>j��>�`����>��9?|�B?-uS?�kb?��?�C>
���-�Q�a>c��>��@��q���+ >J�q?���>u�?c��?uہ>��Љؾ�-��J�>�"q>��.?��g?�y??��?GG�>b���>�H�"��>_?��?�l�?�+�=��?��/>��>�O�>t;�>��>7)?��D?�v?��K?���>��Ỻ�2�w���Q����ׄ�O;�X=>d��Y8�<��>z�ν7B�E�8���A;,�ͽe �m�d= �?��u�=��>Yt>!��g�0>
�ľ�È�	B>Ӡ�ٕ��.w���:��L�=�^�>��?a��>��"��P�=��>3Y�>�v��$(?�,?�?(�:�Eb��ھ9�L��а>>gA?���=Ûl�b���4�u�2�h=P�m?�'^?��U�^���#Yc?��^?�󾋸;��V˾�j�@��n�I?�/?mH��3�>�V{?Sq?t:�>�Ml�_ui�U����b��H|�WԳ=��>.���ag���>ٜ5?c]�>nZW>!�=\ վ�u�-��� i?���?�&�?cz�?u�>� q��ݿY,�~R����Q?.��>��ʾ�=?���\��Hɛ��jԾ�L�Q��Hzƾ��ټ��5xD�����3o��5�=�?&Z�?r�?Y_i?����Q�G�@�=Ä�E~�(��?�	��y��W@���$��u��3�6����_@Ҿ����W���J"���?y�R?��ƽ���>��?�yH)��+�<�,=_�t�Ʈ�|~�<N��=�ӷ��¶��c��맾��侭�%?s�>qi?ӻI?�E�9Z$�>�6���-�*���=�i�>�f�>�_?z��>�E��q����	1̾��Ǿv�>��e?�B?S�X?��A���'������5]����">	e�=�e�>�?���J,����2���u�������'��c�>��M?P@�>*��>�ʩ??�(?},��>w��+f�H!��Χ��؋>A^}?��>�Q�>�FR=|d�8v�>��t?-��>qӀ>�q]��t'�X�f�9:;\�>��>�k?pH>����\X��%��?����3���>b�y?�j��	���>x�>?@&��=,��K>E_�����ξuмW<>ö�>52(�/U}>�������I�k��;��%?�,?F��O
�#��=�Y:?[%?P>@b}?���=�޾��M����>�\l?ߌB?@cQ?�*?�8z>$ ��ȧ�R���zN=��|>B��>�x�=�J=)'��)��H ���@>П=>bQ�=�;�=尲=y�v��l�=�K=|r>�@ۿ�K��vپ��dF�T
��a����������c	�Q����K��?Ax�����&��YU���b�2c���?l��d�?g+�??w���������xv��:����>��r��ς��@��L��y��
q�Z��W!��O���h��e�AiN?k����п�������?xo�>*Z?=6�#!W��\�[>qS� �ƾo#�Tŧ��wԿ�2���	f?�F�>U�ԾX��<�>
�5��k^>�dv>
!Ǿ(�=��z���>�R�>y��>�Z��߁ƿ>Wÿb}ʽ�Y�?�j�?SuA?�(�z���sW=���>�	?@>991� T�DӰ��+�>�7�?���?qgM=��W��$	��pe?j�<��F��^߻%�=�b�=��=ߛ�('J>�G�>�}�JqA���ܽ�~4>0�>>j"�����D^��w�<jO]>t�ս���3Մ?!{\��f���/��T��&U>��T?�*�>g:�=��,?_7H�]}Ͽ�\��*a?�0�?���?'�(?ۿ��ؚ>��ܾ��M?TD6?���>�d&��t�ޅ�=<6�%�������&V�l��=O��>m�>Ƃ,�ً���O�I��"��=�� �V�Ŀ���h"��Y9��J�V�7��ٌ�s���ò��J����|���ֽ2T=<p�=�X>f�f>ߞK>�u>EV?I
t?���>�	7>xm��P����ž@�\a��4$y�~𫾑q��_=����Ͼ�<��4��&q�2t�pa���g#�rv�=�zN�{��H�shg�;0L�� 0?���=��վ;�8�	9�=C���@�����g�ѥϽ�zھb(6��tj��0�?��4?�᏿?:X��E��*ϼ�-��۟d?�M9��������P�>\��,�`=\��>Ք�=ُ���"��@��@0?"U?���Z���{�*>� �:$=��+?�E?q&q<$(�>�$%?*�]s��R[>��3>sף>���>�G	>����ܽPV?�vT?t �.U����>PC��_�z���_=w�>��3�p�/�Z>dS�<��8^��ʏ�s2�<�X?��>�z-�I�M���X�A��=��{?W�?�ו>*ih?mD?iK��{�����R�N%���/=�
S?��e?�X>����34վb,���03?�qh?��P>^�g�:�۾�-�]���	?��n?��?�ܼ�}��Β�P�ݑ6?��v?�r^�vs�����L�V�v=�>\�>���>��9��k�>�>?�#��G������pY4�$Þ?��@���?A�;<��K��=�;?g\�>�O��>ƾ�z������B�q=�"�>���xev�����Q,�`�8?۠�?���>������[�Z>w"��zX�?Q�?}��Z_h�n���?�d�;�;{�<�=y��C���)�����4�WΔ���cE��)��Qs�>��@cT��p>�#�_ӿIWԿ���U򌾓9���>���>WF�:����x�4f�G�6�He��`�bͨ>b�>G泽}i���v�+(8��X�����>��1�Z�y>�'K�+�������x���ԋ>]:�>�΀>�h�����?���|п�3��?Z��RR?���?p�?��?�'߼�}���i����@?�q?�V?��t��!;�a//�>�y?������_���C��0Q�M�=� �>�>����1�:�r>��>�T��]\\�?I˿޲ҿ�R)��O�?��?���R��>� �?"5?�4�]q��tǱ�0��|�[�>vn?�ނ>��վA��������,ž�?'�L?E6*�s�-�]�_?*�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?ӵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�
i	>���?�~�?Qj?���� ����U>
�}?K��>B̄?�+�=���>�(�=������%>zo�=��/�ӯ?ՋM?@�>��=*P8�&�.���E���Q�����|C���>QLa?��K?�Jd>����L�9��� ��eν�$3�Ҳڼj<�"�+�FX�t�7>�:>O/>�E�N.Ҿ��?5p�*�ؿ�i��>p'�z54?	��>�?�����t�����;_?z�>7��+���%��C�R��?�G�?3�?��׾rR̼(>�>�I�>��Խ;���������7>7�B?]��D��f�o�v�>���?��@�ծ?Oi�<	?L��P��}`~�����7����=R�7?X/��z>���>w�=�nv�仪�>�s����>�A�?{�?4��>g�l?��o���B�k�1==K�>s�k?�s?��o���o�B>��?��������K�t f?�
@u@�^?��X�׿`���ƾ�6ʾ9�=��=��A>����Pa�=��7=�~�<�y�ɒX�><�>Z�>?�>��z>?">JV&>�}����c����2����C��&��;x�����YY���9���꿾'k�d ���H=�_G�

���F�#���w��=�R?C=Q?�r?�?���U%>����D�9J	�}�R=��>�1?�I?O(*?:��=���Bc��р��ѧ�������>��R>���>o��>r��>��}:��5>.r+>�:v>��>o.=$3�C%I=չ6>��> ~�>�8�>�p�>ެ�=�,��_��J�E�����5�@ͨ?z`����S��)�����Ε��u�K<��?WW�=s���ɿF"����G?~��v�+�6�:���A>��;?�M?�eR>ljD��ѹ���/=�?�i�0��*>>�Ͻ���;5/�u�y>< ?L�f>�tu>6�3��_8���P����� �{>c�5?¶�H09��u��H�\ݾXaM>Ћ�>�o>��o�����;�8ji�H|=�h:?d?R����İ��v�<V��3R>��\>p=x��=&�M>��b�C]ƽR�G�ݧ-=��=��^>&��>�(%>��=f=�>p!f��D�:�>�GV>�a�=j�C?��?`��:e;��������t�>���>���>��=*yN�Ry=m��>v}r>�����	�����֬)���2>�����|�����8{s=�љ�O*>��==�'���P����;�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�m�>!z�L[����_�u�\�#=D��>_;H?�P����O��>��w
?C?�a�����ȿf}v�%��>��?q��?A�m�8A���@��|�>
��?�eY?!gi>�[۾[bZ�U��>��@?�R?!�><:�̙'���?�ݶ?���?>"O>���?ҙo?���>�(����/�����'�����=�˾;�_�>��=&e���7C��d�����0j�v����U>�S=.}�>D8���Z�=x������<e��D�>F�x>;�K>[֝>�L?`��>�>7U=*������Ś��O�Q?9��?����-i��Z����}��R>?g2?ɱ=oʾw;�>Ղ{?x?��'?K��>��N��Ǌ���S��sC��S�>���>U�>��?;0/^>�/���փ� ��>av�>��O;������W�M�3>
-�>��?���>kt>*�!?�� ?;Oa>�c�>��C�����2H��j�>���>|�?4~?��?bpȾ��6��^���a��>�[�U7>��q?ޢ!?8d�>������,MB<��Q�`ʆ��4�?�+i?�V���?�ֈ?;9?�??D�v>M"��ݾ�V���u�>��!?���D�a�%����Q
?��	?��>�C��1���ql3��	�vr���~?��Z?��'?Dg���Z���ž(�=��ӻa(����;av�#>ߩ>U���C�=c+>���=�#j��5���<��=m@�>�N�=2�-�[ؗ�#=,?e�G�Bۃ�Y�=?�r�9xD���>�IL>`����^?�l=���{�����x���U�� �?��?Ck�?���-�h��$=?�?Q	?�"�>QK���}޾���Pw��~x��w���>���>]�l�\�H���Й���F����Žn�3��h?��>�{?m>?#{�=0�>~�.�f��r���r��$�[��:�a'�X-A�R�%������	�æ�;�����_u9>�}��?��>��?��a>{�>N�>͢�V�>�Î>N�`>�f~>�~�>S�=R��=��>�֫=JR?F�����'����<����3B?�sd?�*�>"�h����O��8}?0��?�q�?EBv>�wh�'+��o?�9�>f���r
?�:=z��=<S����#9��_�朎>�Y׽�:�PM�iqf�h
?h/?+����̾	Q׽0*���e=��?�5'?�����T�g5��H�^������n�������f=��N�Ef��߃���}��
Y��S����d?�U?��7��W>��F��*a��=�ǋ�>�} ?��>�D�>���>�rD���r��H�<O���a����> bv?�ߑ>��;?i`5?fNS?1�D?r>�@�>�pr�*<�>�h8>��>���>�b3?�#?��.?�i?�Y$?�)=>����)���(�Q�?��&?��4?<�>uY?�	D��]�ҁ�ׂ_�6d
���ض���ܩ=��7������=qSA>DU?����8�������j>Y�7?p��>���>�
��5-����<w�>!�
?�D�>O����ur�]��Z�>��?*
�ki=p�)>`��=�����2ۺ�b�=T¼D��=ḁ��S;�ĝ<?f�=�=�w�T���9�:�W�;s��<or�>?�?b��><C�>>��.� �G��!z�=Y>SS>>�Eپ�|��$����g��Vy>�v�?Pz�?��f==�=��=�~���U��������S��<u�?�J#?YWT?��?��=?�h#?��>J)��L���^��Q��#�?�R,?�
�>�/�&c˾�쨿�G3�MI?0?�`���U)��>¾ǥֽ&$>k�/�%�~�����C���e��������?j��?$�A��7�MV�A��������]C?���>O:�>$s�>N~)�*�g�����;>d��>�R?���>��P?.z?�9\?�3[>�9��������Wּ�? >G >?���?|̐?�{z?�>�>�>)l)��q��������Q�ڽ�酾�=RR>C��>6��>E�>a��=w̽y����;�VC�=/�j>��>�"�>�c�>�}>��	=�!C?	�>�rվf����e�7� X=4�]?
��?=S?��Jq�L�B�;V㾯��>_��?0��?��1?�fY�њ> ��;�!ɾ��{����>S��>���>Y�=b)>=|��=�>B�>�S2��I��4�ƍ�l?a�K?��!=��ſ��q��{p�.K��@Ce<������c��M��nZ����=&�0�����2\�&�����A����P���{��~�>]��=�U�=	�=*��<�>Ӽ'.�<V�E=���<J =��o�Y�t<�9����b��~�:�hwe<�SG=�B𻓋˾�}?W8I?"�+?w�C?��y>F>q�1����>�;��B8?'V>�P�T���z�;�K���� ���ؾ�S׾d�����>ҹI��>�3>K �=3�<�m�=�4s=���=}kG�E�=��=u��=�>�=?��=A�>�>�6w?V�������4Q��Z罦�:?�8�>V{�=��ƾk@?k�>>�2������vb��-?���?�T�?@�?Fti��d�>I���㎽�q�=R����=2>o��=s�2�S��>��J>���K��E����4�?��@��??�ዿ̢Ͽ.a/>9�<>Oa>�eT��=1���`��yX���L���?�8�l#Ѿ)N}>�ֲ=���ľ��:=�=>�Xu=E=��[��G�=]@n���=�Na=�8�>�E>�d�=/���L�=�"=���=�pK>�����m�¶3���6=;]�=�g>V| >h�>aE?�?B�F?=6�>�%�(����p���ǚ>(D>�>F�j=�n2>�=�>�@?!�C?�W?-y�>!�=̍�>9��>	�4��*g����i��,�\Me?q�r?��>�¼�hw��.���A��j��`�?L�/?�!?�>��K���4���L��ì�-�<�mZ=D�ؽQњ;�5���ɽ����潵O6>}G�><�>Cq>!��=�=D><U�>:��=�P<<K=�΋��p�7a_�
�>���=���<z������=n��='��2b'��;<RW�U��M�\�XV�=��>��>�u�>{o�=��Φ/>�d���L����=�~��5JB�W1b�݇|�{�/�y�8���?>�R>����X����?_�[>^pB>�P�?�jt?k�$>
��F�Ҿ|e���c�nO�#]�=��>K3��H:� �^���K��Ѿq��>��>���>��-> �)�V>[��*�^s���'�!q�>�p��^�:�eL
���a�p泿;�����Y�S���j7#?�F��j��>kh�?��L?��?a��>z>����_->>4�u��8��X��zc	>�:,?�X??(�ھ_WQ��]ɾ�������>LFF�6*M��\��&�0��!e�-+��p �>l[��w@ξ�G5��T��ꁏ���A�@W|�)�>��N?b]�?�����À�t{I����Rh��T�?5�c?�Z�>R�?@+?w���eT�󲁾&��=;)r?9��?j��?�a
>frh=u˦�m��>�?�q�?pm�?� d?a�����>��=ߵ>���ݣ]>�=��7>��[>a�?��(?��??�Ľn�!�7�Ծ7ࡾb��-n�l8>2��>�_W>��*�ǭ(�&�>���=�4F>�>��>��<0\+>�t�=Nx��n����?Һ\>E&M>}=�>�N>P�~=^�μ >>\�=xUA���������f��@S<H��b �=q$,>��?s?Կ=��?x��>��0�Z?Aǌ��,���`���N>�5�h+�>���=1A�>��
?�]?��= G�>�޻=ʗ���=���+��-�3N�s㾶E�>�:��"�]�*�S�����ľ�<��rk�]}��@O;���<�Њ?�� ��{l���(�c���;?k�>�f$?U�0�+@��eR=���>_�>|[ ��$��d���3���\�?���?�4e>a�>��Q?�?Ci5�l#�?|R�~�t��t=��c�{<a�R���/p���?�����`?ƴx?�B?�(�<��><��?��(�Ж��&N�>�,��09�4�/=�ݣ>�ݼ���j���ӾŁɾa[��A>�:n?q��?�S?0�a� �׽
�9��g,?��;??pX?dY2?��]?év���$?5>�G�>�	?�>4?}0?�-?�=m>��]>�Z�=�;�<o2��.>�L>Ž��e���<D=a�=-mȽH�<2e�=�ҧ������6�Y�	>ʮܽ��<�0�=;U�<��=�~�>/�r?u��>�ӑ=~�a?��>
!�"�;c�	?���>���>��1�w]#�L-��]�>�fY?[I�?�B�?���>�FF�Y%��/P>�z�>�@>%�>Qc�>�X��a���> ~�>���=�	>����J�߾�~��v���?w >�>���>�z>���� 1>�����{�|af>V�J�(q��"F�SZG�b�/��p�L[�>;<K?��?��=(6龠0��G_e�q&?B�;?K*N?���?�~=�CԾs�7�I	L�E� �?��>s��<��	�|䡿U��x�;�� :ibt>N(��,���2�a>Pc�
�ݾM�m��J�A����S=-B�M� =�g
�m�־pǃ����=���=o¾�t �B���A�y3J?e�=�Ъ��5^�$q����>�ܒ>.H�>��*��<��p?��s��Ӭ�=���>�4>@9u�j@�F�K��7�>�-K?��Z?<q�?m䚾_5v�a G��������	׾�l�?�f�>(w�>7��>Yk<����=���`��tN�l��>�;?4$�9�H�Yr��k�U5��N>��?��>]�
?�T?M?1�X?a�?#��>x��>�]ܽ�+ؾY�?g�?0>�=�~I=�Z���+��F�� �>�1?U�����>k>?Nt1?$�?�a?�d:?C�>l�+�F����>��g>��Y�Ǵ�� >��V?��>�C?��?y<>|#�5����6�H�]<�V�=��??T|Q?�3?���>TD�>��콋�0�Ω�>��c?>��?���?
�>��D?��C>�F�>�6�=��>�ؽ>9�?z0?rq?�n?5�?�V��Y�K'��Y��ĽnqI�V_=�>Q�S˧��"����9�f�3:���=A���Ѵ������=�[�>��s>)��&�0>��ľ�L��j�@>�x���O���؊���:��ڷ=Z��>��?X��>�[#�Y��=ͬ�>�H�>����4(?'�?w?^�";��b�&�ھ�K��>B?���=��l�?�����u�zh=�m?��^?�W�$����b?�]?�e�4=�a�þ��b���W�O?s�
?L�G�Y�>S�~?��q?v��>�f��8n����Bb�`�j��Ѷ=�q�>�V���d��C�>К7?�E�>��b>,-�=+h۾��w�j���?�?�?D��?,*>��n�D1�zx��l4���lZ?)<
?��)�?�F>p4þ}���,��ݪ�፨�����`뇾oɓ�Z���d�<`���hy><J'?��c?��x?93j?��(�2m�!sN��}p��2a�2�/�YA�NjR�AsX��I��[v��9�ͣ��]���.*��}���Y=�B��?�?s]U���>P�g�7H�[U�5<>�
���恾1��=�4�<�!]>#:��Q��y�l��Ӿ�q=?���>ᗎ>A��>s][���Y�n:G��� �j,���.>gt?f.�>:Fh>�#̽:8���n��s���6����b5��8�>�$i?8?)�K?��R�4�r؎���-�tv4�s��W��$>�L�><�*����<�255�&�Z���#�'i��R�
���<>�A?OG�>E.�>��?/�E?��1��*R�d��O��}�=���>d��?���>#�>�uD<)ᴾ��>L�l?���>��>����bo!��{�+*̽�>��>gc�>z�o>��,�!\�$m���}���9�m��=#th?b�����`�)�>sR?�z�:�L<���>>�s�Q�!�hs�E�'��->[�?�%�=� <>�TžB �|{�����k))?`�?�J���)�3K�>��%?pH?�m�>6�?�Ԡ>����[�ϐ?�G^?rKH?��B?���>�N�=7�t��3���Q*�T�=�5�>��_>��&=�
�=��%��\�;@���ݙ=���=���)֝�C���[�޼�/<�i�<e�&>��ٿ�J���Ҿ:d����z�
�8M��ꣽ�0�����0s��_*���y�J��Ҙ�Ga���`�v0����r��}�?��?�@���'��i�������� �W��>Ip�雋�����������1�޾^t��� ��qP�2i�i�d�`�7?�.��3Lʿq���D����?�5�>�f?����Z"� �%���>-�[�D�M{��&���zҿz̾?Z_?�k�>6:ľvB�3ݦ>��>��	>��>�e����U�� �=��>K��>���>���%:Ŀw����ཽ#��?�_@ҁA?��(���쾆�U=w��>�	?/�?>�L1�]A�����l�>�9�?(�?W�J=̷W�r��le?�<�;��F�͔ܻ-�=�^�=,5=���ȼJ>#W�>.���%A��;۽m�4>⢅>� #�����^�3<�<Vo]>��Խ�/��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��=�����M������t�)D�<��R�PM���n��MI��x�*�ž}ª�zX���� =�e�=eJ>��>���>�<X>
�K?�Em?��>z=z>�ճ��C���޾�'e�����X�����6�mo�9��@Yھ�z��e���2�#�ܾba�1�;�O�����:���#k�Z�M�;�H?Gɺ�����#��x��V���U����U�x�V�!���l>��v��ߦ?k�.?A��N.f���о�\Y�������`?w��KR!��>޾B�>��8�o��f>��u>�����:���K�@j0?�T?AC��T��*Z*>� �G=3�+?��?F�c<ͪ>?%?xm*����(d[>|�3>f̣>B��>+4	>3����۽�?�T?@Q���g�>��S{�Na=�H>7�4���鼞�[>���<E���U�Dӏ�,ҿ<+W?{��>R�)��
��M��l��&==�x?9�?B)�>�|k?��B?�	�<*�����S�8��v=��W?O$i?��>dy��0�Ͼ����4�5?��e?8�N>RUh�L�龺�.�[��?��n?�_?li��U|}�!��[��3x6?��v?s^�xs�����K�V�g=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?}�;<��S��=�;?k\�>�O��>ƾ�z������.�q=�"�>����ev����R,�e�8?ݠ�?���>������C$b>n�����?��?��q��T��
d�v��T�v�(]w�%�T��P>��~���U�ƭ�#z��柾VWE����>R�@jrO�%uG>⒀�:�ڿ���p���!d����Cm?)nh>{g��
C׼����މ���K���_���#���><C�=��`� ��,u��6=��<�Uy�>(����]�>0�����nQ�����<稑>L��>�8�>��ֽƦž/e�?��[ӿ�~������M?U�?M�?��?Hܘ��1l�]G{�dM�֬@?0*d?(�W?����X�i��lU�C<l?�X��a���:��NA���:>%.?1L�>۟-�L=�o>.��> ��=��1���ÿ-2���Y�=Z�?6��?��G�>��?u�,?������w.����/��⻴�B?`�8>�$ƾU+�3�3�z���,�?��,?O�MX�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?`��>���?��>�?��(>����5�i���=*́=�>,=;I�>ݢd?���>@�>oR��/�/��=�x�;��龡G���>hXV?�Z\?S�>i@��J�g���$�vp2��<���3=��U��<�]��y�>�[I>��>ç`��ힾ��?;p�/�ؿ�i��/p'��54?.��>�?���1�t�����;_?Kz�>�6��+���%���B�R��?�G�??�?л׾gT̼	>,�>�I�>�Խ����e�����7>,�B?R��D��c�o�o�>���?�@�ծ?Ri��	?���P��%a~���#7�+��=��7?L0���z>Y��>��=�nv�ͻ��8�s����>�B�?{�?b��>4�l?�o��B��1=�L�>��k?�s?�bo����B>8�?"�������K��f?�
@su@y�^?�9ҿ����s6Ծ��⾌I�;��F=�w>��<�^�=�M2>�ｭS\�%ϭ=��>\�W>�r>���>���>��E>�~���!Ɠ�嫖�W�:��"���X���F������v���������٫�vV�<y�ý���8��Jj�=k&P?�[R?��k?�?��g���>���s�غP�(� ��<ɕ�>i�1?&�L?~J-?�1�=�l��;^��&y�Ws���+}��.�>�wV>a�>R1�>N��>�QU<�k:>u7%>��x>��=W E=��<KG�=`f@>@�>�%�>&�>e��>T{=3rĿ�f��{-��=���M��}�?����n���u�	�-�Υ����+?���=짌��HҿK��l�F?���z�e�"���->Qn+?��7?<N�q�����z:^4<>��Q=����W5����pR��!�?��6�=�/?�f>9�t>��3��f8�:�P�tn��k�{>6?K���g9�*�u��H�m�ݾ�L>���>تG��m�����x�~�%@i�T�{=En:?*\?��������nu�� ���gR>�b\>�=�T�=�EM>��b�A�ƽ8{H��-=) �=�>_>�9?�U,>��=�գ>D��5O�֋�>�|B>ҭ,>�@?�@%?BF�S������F�-��v>��> �>u�>*fJ��y�=N	�>6�a>���1��!?�M�?��VW>2n}���^��Ws��y=ꓗ�&u�=��=\C ��w<���'=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿla�>�k��X�����-�u�S�#=���>l6H?�H��vO���=��v
??
a�G���)�ȿ�zv�N��>��?Y��?>�m�A��u
@��}�>R��?qeY?ai>ph۾7PZ�Ս�>��@?UR?��>�7�@x'���?�޶?��?��>�В?i�@?2��>�-Ͼ��C�����H۠��`>�n5���{=ؐM=�ľ�������[Yy�~gW����hg��[=2.�>Ss��8�>�ռZ��*����>�$�>cd= )�>��;?+�	>�8�>�A�=e����z<���Q��6L?ỏ?_����m��V�<��=h�d�R ?�{4?�@�f�ѾxS�>�J\?X��?*Y?���>9��v��s��n���j�<)HL>Xh�>�2�>����K>�nҾG�
��>��>إ����׾4у�m�ݹ�0�>�� ?� �>2�=�� ?2�#?Ŗj>�'�>{aE��9��z�E����>���>)G?3�~?8�?�ֹ�^X3�����桿;�[�6N>2�x?�V?�˕>叏�2����lE�,PI�9�����?gtg?�V��?�1�?�??��A?�!f><��hؾޫ��_�>��!?<U���A��h&�o~��[?@?���>��0ֽEdϼD����؍?=\?�(&?Ļ�^La�y%þ���<�� ���F�A��;��G��>�_>"���g�=�>0X�=Οm�Ms6��f<�˻=��>��=��6�!��0=,?��G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>�l���K���ڙ���F��_�Žw1��� ?[��>�o?^��>_z�>*ɽ>�6������־���bVN�'C��$/�0��@����]�L���2�`8;��'=>b�Ž�-�>>�?�.x>YȦ>O�?f�X�!ʲ>ո�>�`>W�>J��>��=Q:>.�i=�5� LR?1���	�'�F��L���
3B?Xqd?c0�>Gi�3������W�?|��?Us�?W;v>�~h��,+�Ln?�=�>+��Pq
?�S:=B��A�<�U��#��^3��R����>�E׽� :�AM��nf�zj
?�/?y����̾y;׽_g���wG=�B�?-A&?B'��Q���n�.�P�n�U���� �M����#�a�j�H���px����)���<![/?m��?���eg���P���m��IB���Z>���>{�>SV�>lJ>&��π.�5E`�q'�AȊ����>�u?UL�>~�I?7�<?D�P?�eG?�>QF�>2m�����>��m=]�>���>_j<?''?��(?��?v�)?�)�>v�Խ�h�p�Ӿ�C?�x?~#?^y�>vM
?�ol�T\���7S��@�;g�2��ZT����=�ё=�a��̽dp'=j�f>�W?|{��8������j>��7?�>\��>�폾 ����<� �>:�
?�b�>�����jr��D�Vw�>Ꞃ?e��\]=��)>���=����$ںb�=Aq��x��=�ၼy�;��<X�=�Ӕ=
s���s�#��:�d�;�0�<�t�>p�?���>/D�>@���� �+���c�=�Y> S>�>�Eپ�}���$��1�g�8`y>�w�?�z�?��f=��=���=k|���U�����D������<��?�I#?VXT?i��?��=?Hj#?<�>/+�|M���^��]��ٮ?�)??
�x>�T��]����kS����>� �>$_�"�޽�	���J ����3`@�K�H������d����F���5>����M����?���?�g��|�F��������~ƹ���`?U�>�8?>�$?$;b�֯����>Rl�>�^ ?U��>��t?m~?c�?��>'�7�M������?r=䭿<4#?�^�?P��?�M?�?Cv>9�G�
���G���ϡ��E���1��#�=�*I>{��>���>@��>��>�-��A��������M>�&;H��>'q!?���>���=�����E?�B�>Jy���#����Fk��(I��9m?�@�?�T'?��4= ^��N=�� �%��>q��?��?�8-?�I�`7�=)���4��W�����>f��>ѡ>��=�I=VMG>�k�>�B�>V�������=��t����?WQ?���=n̾��bO��ܴ��h[�KXz=������B�P�t��Ҟ�V�<�X�+y��/�V�[�� �E�x�;�|��t���釾o��>�i�=fK>�/�=
� >"��=!/�=E�=���8����d���e�= yf��9>U�>��<�	�=�v��U��S;�}?�z@?��?�4?У>PO0>G�v�)ݱ>�eҼW-"?nQ^>"끽�����.�B澾�ۢ��۾\��#�p����[O8=敌��1>T}>A�=���<~2>aϪ=h�>}8�<'\=Cv�=R�=�Q�=�%>H�6>hX>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>:˕>��{=!Jr��A@����"�z�_���?%R���پ��>!�7>���Yc���=�].>����L(��cPd��u�=�+��F�=;�d�\>`�V>d�=�k~���>�>٭�=d�>�y��驽��V��\*�/"r��k>(��>���>j�"?� ?�(n?_ �>��0���Ӿ(sɾs�>8U��z�>ʡY>���>P�e><>?z!k?$V?��>�
�<<��>7@�>'�(�q�Ţ�q=@�μ=�)v?�ׅ?���>��a=������'�S�2��d�#H?.\?�9?���>d��p޿��1�d.U��cz�㔽�R�=%A������ch=`�L������=�K�>��>T�>��>@�>Լ�>�=�>�8�>���<5�(>���=?A��'Z��v���W����X�X�L���S���9��qJ�
�[�`� ���=�	�e��=� �>�$>�^�>9�m=�M���2>[w���0J�M�=������@��{a�'H}�f{.��f6���/>|PI>�̉�����?I�J><>-��?��z?�v,>n�罇'�������V�	 B����=R5>);"���8�!�[���I��[̾���>��>fV�>Y�'>tPB���D��<5:�-�>��7+?(��&H�>+7���^����}!����x�`"��3,?�����F=>;]?%6Z?�\?��L?�=<pڽ�F�>���J�.���!O=�����,?�uB?��?3�ɾ
@<��A̾㎾����>/I�i�O�`����0�='�ZK��z�>���ћо��2�J^��揿v�B��~r����>��O?)�?n�c��J���N����έ����?�7g?���>�=??c�����=���g�=R�n?��?�:�?�=>�6=/mǼ���>E�	?�0�?�٘?ɑs?�"�K�?��3��_>��9� @>tB>��
>��>�?C?+�
?r����9�I��Òо��뽥4t����=�E�>֠u>�>+>O�9!��=�0��0nB>��>��?>�7�=ӛF>��V>$5��8���c� ?r*�=�jX>S5?���>�`�=`�(�>���=Se^����%0����<�B�j�M<�\=��$><�
?��Ϳ��?�7�>r
�ʧ>Bd9��ՠ9�Xм�;>pS�q�l>0�@>���>a7�>%��>�V�>���>E�>�B��@b�={3 ���0�} /��yK�'���Xi>����� �������wZ������Jeg����H���<�?Z���!W�4�.�AD�/�>v��>t*?&?��e���=\=#=�>��>�>Ӿ[��O��G�� �?3��?v>c>R�>7�W?#�?��1�!3�vZ��u�1'A��	e���`��፿a�����
�Q��3�_?��x?wA?�
�<�:z>֣�?'�%�׏�J)�>_/�s);�'+<=�.�>M)���`�ԬӾ|�þ�/�SAF>�o?�$�?)X?L`V�����
�=x�4?�$?��a?h�5?��G?r����?0.X>.�>��?\88?U84?'?A>K@>�1�=E�;=ĳT��Gw��X@��B8�u�7��=�'V=2;+;7��?>��[�����ޤ=n	�<�D'��=f��=�۱=5�=iâ>/k?��>S��>|3/? ō=y���о��K?q�)><-�C/t�D���k� ���=�[�?[q�?�2}?�u�>	KM�:pd��<>7�>�>x�>�+�>7���9]���:>�n�>gy��vM�=Q�=lf��co/��f��P�X>�qu>���>�0|>2��%�'>�|���0z�Ĥd>��Q��̺�l�S���G���1���v�Z�>�K?k�?E��=C_�.��QIf�0)?�]<?�NM?��?�=X�۾0�9���J�/>���>z^�<��������#����:��N�:[�s>�1���*����c>�-	�Hپʄk��YG�����Q=��1�?=�)�2lӾ��u���=;�>Bʾ�c���|������I?!-�=����
�Y�~���$�>H��>��>#������H@��嬾mܓ=���>fO3>,�ؼ��@�E�l���>8�D?= _?�-�?ှO|q�n�A� j���t���ռ�U?o�>%3	?#)H>LV�=_̰�]F�z/d���F���>��>���H�����;��!f"��p�>�#?W�>)�?VP?��
?pi`?�(?��?*��>�a�������#?���?�z�=(iȽV Q�r6���@����>o*?��N�R�>�?��?u,?1�Q?��?�>� ��*A�c��>�F�>��V�zj��3�U>��G?��>v�Y?��?�R,>U�5�9ݩ��շ��+�=S�>��.?� ?l�?�>���>Џ��R�=��>��b?=*�?��o?Ý�=m ?��1>���>��=��>Q��>�?�IO?��s?>�J?�[�>��<Rì��u���t���R��b�;��M<v�z=f���Au�����(�<SѰ;+���J���@��J�D�nv���O�;��>��u>�Ď�L�3>q�¾u	���B>�$�=��kӆ��>�e��=+�>$� ?�>��5�|�q=�^�>[�>�2��0)?�"?qf?�w.���b��2žU^[��Ա>�>?�o�=!2j��A��2bp���c=��i?�)\?R2k�#[��Q�b?��]?9h��=��þ��b�Ɖ�n�O?2�
?�G���>��~?h�q?E��>�e�*:n�(���Cb���j�AѶ=Xr�>PX�L�d��?�>n�7?�N�>�b>v%�=ju۾�w��q��c?��?�?���?+*>w�n�Q4࿴���G���I	[?���>C�����!?�Fu�/�˾���j#��;V��J��F���.���䰦�R~ �M�}��*��b�=$�?�	s?1�l?��\?����V9a�]L_��Ҁ�خR�5���!��)=��3B�=]B�8Wp��S�`P���	���=����fg/�h��?�/?�Cý��>�e��{lվ^UƾZQz>
��z>��!�<�?.�nnV=��M=�(��,��ξ��?߳>��>u)?�jQ�e!/��Y-��K=��P��E��=1��>u�>��>��=�b{���R��{���o�=��1t>=lc?��K?��n?�W���1��y���r!��:�������A>��>嚉>E�X�Ү�yN&�^8>��r��s�ن����	���z=�3?���>�Ü>�ۗ?2N?w�����h�w��y1�0�x<��>�Ai?���>�ɇ>�ѽ2!��Q�>�Id?��>��=�'�����\�����;x�6=|�?��?�(�>?Ԏ���X�����uS���p�p��=Ʒ�?/������>k�?�C>��	��m�>a(�=�bo�p��,���T�=O��>�\�u6>�料���R9��Y��)(?/C?& ��]�)�c}>kJ"?�$�>��>D0�?*�>#=¾�z���?�_?T�J?��@?\ �>�N=Ϟ��bŽ��$�s4-=���>�JY>�u=�>�=�r�[��d�!I= ��=�ټ򣼽B�<i��G/<8*�<q*1>�cۿ
5K� �پ��� �.
�����󕲽�N���n�䄵�����x����X�'��	V��c��ό��6m��q�?�4�?���t'��X������������p�>)\q���������V�V�����W�u!��P��i��e�I�'?�����ǿ밡��:ܾ!! ?�A ?)�y?���"���8�W� >�D�<-����뾫����ο)�����^?���>��/��J��>ץ�>�X>�Hq>����螾�2�<��?&�-?��>юr�%�ɿY������<���?+�@�A?n�(�Z���V=���>��	?)�?>�71��J�����/N�>�:�?���?qaM=t�W��
�vxe?2�<��F��kݻW#�=%@�=�_=e����J> [�>����HA��Jܽ
�4>4؅>Ϣ"�����^�C�<��]>;�սN*�����?����Fʒ��vF�,���	>?��h>�Ʀ>�,?Ao���YӿHƏ��O?�%�?Ժ�?�O?�E���x>Z����E?˷?e�?s��O3��݆=xN�=��F�Ok��hW�O��>��>�:��E��6(�P�!��S2��&<>��ѱƿ��$�^f�"�=�aӺt�[�?=罬���d5S�6��o�o�u��Ug=���=0�Q>$x�>��V>Z�Y>#VW?�k?f;�>�z>�9�v��ξ��NG���/�����f|�B룾�W��߾r�	�V��b��D�ɾ�#=�<7�=
�Q�6 ��/ ��b�Q�F�ח.?�$>�ɾ=8N�l}<x�ʾ�૾�������<˾�2���n��@�?�B?�����V����~����ޤV?�^���G���|��=g�����=^:�>�%�=���w�2�#!S��G?y�?0��c�t�¾F>?1�Uϓ���1?`��> �<�8g>�g?P�F���8s$>�Z�<��B>�=?KJ>��������4?�Q?��,���Ѿ��?��ھ㹊�|h�<aT�=@>J��'�9Љ>�>�&�������9�V6=�_?ޫ�>�b��a��[����h��e��a�?�[�>���>�l[?5�B?�	�=���BF��`�_�;�#p?mN`?,�(>-�\������|�6?�`?=k�=��p�W��?�.�޼��y?MW[?)@!?� ���i��ه�4���4?�u?6h�S����[�R��̵>��>�V�>�3�e"�>�K?��)�𮗿�m��ۀ5��h�?�~@*��?��8b	���K =��>Aq�>9,�S�������zm���:�=���>q\��Pcv�a]%�/�wF?k��?�V�>Mڌ�q����=靕��?���?!奄	�q<w��zk��c���Ǯ<P��=��Q�*�J�#�7��_ƾZ.
�5��҃��ۅ>G"@���c~�>�=8�����7Ͽ`-���;Ͼ�	v��?�q�>�Lƽ�)��Ck�ʧu��#H��|H��Ō��O�>z�>������ �{���;��0��c��>���#�>��S��Ƶ�9���.�<Ϩ�>���>E�>�Ҭ�I���D?����F ο��������_X?/2�?���?�m?H\<$�u�]�z�8��~"G?+s?��Y?�1(���Y���6�l?R��4�[�Ɓ1�CC�BTB>�Y1?�_�>��.��܃=l�>A�>�> v,���¿Ķ�*���d�?�?�?�P�)�>�ݝ?�,,?'
�tJ���h��(1,���;$�>?��7>Ow���'#��9�oN��2�?Y�.?{��+�ɸ_?2�a��p�F�-��ƽ�ݡ><�0��g\�Y&����+We����\Fy����??^�?��?ɱ�� #�H5%?!�>ʞ���8Ǿ��<L~�>j&�>M,N>�G_�Ѳu>���:�ug	>Ю�?�}�?tj?���������Q>�}?�X�>;Y�?�:W>�,?��=�.��%1�=F_�=.O=�镽��>�;?�F�>7�=��B��<���B���(�:;ž�N�AX�>��a?��J?�>R>�~�<X)O=��?�?Γ=�����;�Z�������c>쥠>8>�u�������?Mp�8�ؿ j��%p'��54?.��>�?����t�����;_?Oz�>�6� ,���%���B�`��?�G�??�?��׾�R̼�><�>�I�>?�Խ����\�����7>1�B?X��D��u�o�x�>���?
�@�ծ?ji���>��%�����\��q��x9��}L>hf ?�����E>�;2?Y��a�z������2��>Y �?�R�?�o�>��?�q��~l�,�;2C�>VI�?��?ˉ<����b�<Q�?��Ⱦ�D��xW���P?��@�"@��`?E���2s���{��5`�J�����=*��=�?�>x�0�w�=���=u�+=�2<w�Q>]��>�R7>s�g>��$>�R<>��>�1}�Q��dj��ֻ����T�x8�a+"�{5����E�jjԾ˫	�����Ͻ�	��[;9����,	<:�hS=�=��Q?Z�J?�c?l�?p�">��>Ɠ˾<>n9��
>�Ց>��@?�h?��??{�=:�����a�G���M�w���\�T��>�y>&O�>�>D-�>r䙼��)>�J�>Rr>��M=���=�t��?qĻa�Q>�N�>w��>[��>�C<>��>Eϴ��1��i�h��
w�q̽1�?}���R�J��1���9��Ԧ���h�=Gb.?|>���?пf����2H?$���x)��+���>}�0?�cW? �>��v�T�2:>:����j�1`>�+ ��l���)��%Q>vl?1��=��	>o# ���^�%d��|e
>vp?45����v�����d����K.=bf�>�n>eL��?���f���~�oV=إY?�M�>�R�T�S��ӛ�il����>�{�>�M�=Y3=�>�Z��Zּ�ߴ�~�_=gE�=+U>>?��*>;�=��>^
���*R���>��F>�x(>hh@?.#?M=��8������J-�s�r>��>�N�>�>��J��=K�>�b>V��T��4�	���E���W>󂽺�[�xj�ki=�K��>h�=)"�=~��̋?���#=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾA/�>9w�9�������u�!=���>��G?
2���G�I�<���
?�?�#�ᦤ�d�ȿއv�ˬ�>��?��?L�m�����@�?�>o}�?/Y?|�j>�۾+yY���>?a@?R?�i�>��ɋ'��?�ܶ?���?��G>�w�?��r?��>|��3/�u���P��
�z=�<�8�>�s>����E��ޓ�}a����j��e���e>5�)=���>�Ὣ༾�C�=�`��9����W�7i�>�*q>NJ>c�>�?J��>"�>Ν=����z�}�����}�K?"��?����-n��~�<�͜=b�^�{&?VJ4?��[��Ͼ�֨>��\?�À?O[?d�>n���=��S鿿�y��θ�<��K>8�>'N�>���)RK>>�ԾC6D�Zy�>"ɗ>%&���9ھ�5���"��wB�>Ib!?��>9ܮ=��"?��?��>4��>��;��挿BN��(?�]0>7x%?n�_?�J?'�-�^?��^�������jX�M��>J�c?�L(?�K>�4��A���=O�u�Y<���ki�?��l?�u�=g�?D�{?�??��F?��0>����eӾ'JH>�Έ>+�!?j���kA�X&�@���? [?���>��1׽ӕռ��������@?�6\?� &?�p�`'a��sþ���<���I�Q����;��F�$ >׭>JȈ�Eu�=��>6)�=��l��j6��S_<D�=�<�>:��=�E7�$2��i�:?����5���]><p��Ac�~�>��\>�3����Y?~M�A�o�o���A���p
���?pQ�?,��?�R���i���`?k�?�*?iF?x�������ݻžUʥ���3�	�+�%�>P]?Yۖ�F��q럿3¨��o��#+L��h��?���>�?E�?ҟ%>�K�>+f����%���,���@�1��.f3�B���#��]��|w6�����nþ�;?��|>���<ӕ�>,X?�ƾ=���=0�>�Խ��p>q(>T>-,n>��x>n-�>'(:>��+�3lR?�����'�.h�B�����A?�4d?GT�>˦l�Oe������t?�y�?.S�?��u>3�h��2+�A�?�Z�>=2��O~
?�n?=U��g�<�����!��戽����|�>vCֽc:�. M�תe�F
?Q�?P׌���̾e�ֽK�Ծ~_�=,d?��,?����)8������N[���*��k�jfľ��ɽ>p���h�V���_�t��g���=��~��u?�w?'�ԾL��Ng往�Y���&�)��=��>0=�>��>bt�>���0$����U��:���ɾ�h ?5��?��>�I?��;?�P?��L?���>
U�>	���{��>Z�;�Ϡ>���>�9?{'.?�{0?$�?��)?s�^>L��g����;ؾO�?5�?��?��?s�?�~������N��,|�K}y�y�x�B�t=�$�<{�нzw���N=��V>��,?j����	/��T�c��>��&?A��>73�>�e��KzK�a���kn�>y?�b>9x��o��c��?P|?����tV=pC+>�h>ǎ�<t�-��%>L���т=����ܽ�m���=6�=�c��f�*��/��z���b=�q�>1�?$��>�F�><��ì �����=��X>kS>�>~@پ�x���%���g��Hy>Ms�?ux�?��f=~J�=�m�=����#b���������
�<��?"H#?&]T?5��?��=?-m#?��>%+�kK���]��n���I�?�/,?ƌ�>�����ʾ�㨿�3�9�?�`?Ca�(���6)�:i¾0qԽ�>XT/��7~�l��	�C��{x����1㘽*��?軝?��A���6��������mH��sC?�&�>@?�>���>!�)�=�g�� �*8;>�5�>��Q?��>��O?�1{?��[?��T>4w8���RÙ�1.��!>@?���?��?=y?���>��>z�)��`�����i��)[U=oY>,`�>_�>*7�>?c�=��Ƚ&����r?�s\�=��b>
h�>!s�>q��>#\w>���<�G?���>�Y��߃�|Ƥ�޸��BL=�^�u?9��?Ԗ+?�=���k�E�BM��n>�>k�?_��?*?�S����=ּ<���Լq���>7�>��>ߣ�=�8F=��>c�>��>[0�sb��a8��jN�N�?�F?5��=��ÿ��i�}g[��冾�6=����w�ѯ���p�SՇ=`ޛ�#���ȥ��.t���������4��?���|z�>i ?dAZ=�}�=P��=��e;j��^�<-�k=:m�:H�=R~�!]�<������Gާ���$��c;e�t=��Ի��L�?�rU?F=?f>?^4�>�B>�����Y:>l¾���>y�0>�Ӄ�5ɾ|:&�����k������l4��8T��I����T�U�A���n>B4�>Z\̼��� [>^#�i!�;^=q�=G�<CF!>C�L>�_>t;�=+��=�?to������v΃��"��r?+��>��y����A� ?���>�a���ƿ�о�~|q?H��? ��?F�?����߽�>����=���X�=�B��fF>��>�7��?��l>)*��ʥ�w_>�3��?��@kBN?aʍ��ӿ1o�=:+:>�C>�Q��W0�39Z�ߋa�'`��"#?��:���ƾf��>U^�=�+ܾ�OǾ�.=�~3>��_=����1[�E,�=8pu�)0=�`o=��>�HE>�q�=������=k>>=F��=�pR>�;Ȼ�V/�(&1�Y�#=��=�b>��&>�\�>�Q?e�/?�Mb?�>[�c�E8ž�̺���>���=���>r�=}�W>s��>�69?��@?D]H?"��>^C=��>��>?	,�0Cm�&龼����==�/�?F4�?�N�>�u㺿�W����R�8�\3ʽ?u�-?5�?�Q�>�U����9Y&���.�$���[z4��+=�mr��QU�H���Hm�3�㽰�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�= ጻ���<� �����=&�����<�vż�����u&�;�+�3�����;f��;@�]<Y��;�$�=_��>�ٛ=��>{�	>A�����>;z�t�2�#,->.�ؾ=�;��_�7gu���&���ν^(d>-ph=U�E�����&?nXw>8>>�i�?I\o?��F�����㮾\ݞ�p[��W�����=���=L꓾�>�g�b��G�ƹҾ*��>�§>f�>�?>�����F�t��:TY��_�i����>3Ο�,�=�gH��qk���������Lm��`�;��V?�����W>�o?�g?*�?C��>� ��T ��g>�1���Ĺ�p!�zJ���n���@?�� ?��%?�L뾆E���꽸��>�'����O�.��
�$�H���i����/�>�E���-羉"��t�eB��#:8�:G���>>}U?���?�Ǿ�,����g�t�� ƽ0z�>��h?P@�>C0 ?�?&�̽���6����k �l�`?.��?�u�?�
g=�dW=�f��U�>I#?v �?��?�i?\Uv�/q�>\�:�Q�>I(#�[�>��>�5�=+�=�?
�?�?ޚ��vp��3�ua��:B�g=�( =ĉ>��>��>�>���=�d�=p��>F�>��>6
b>��>�u>`4���i���#?aT>�>.�1?n�v>-6=�5��`��:j��X,;�(K#�sYƽ�ƽ���<�B��=�ݼJ��>"�ÿ�!�?m�K>E��`?��rY�6XU>�<k>�ĽW�> 5U>�~>�ճ>Lɠ>ʺ>sԁ>D�>�|۾��t>v�ھ؇��gH�@N�&�	�J�<�䄾�"%��gӾ>�>����ƞ��G�BUi�LDw�@8�Z?'>�|�?�����L��L@��������>x��>'�D?;";1n>K �>���>���>��ƾ�S}�k�~����%ȕ?��?�-c>��>��W? �?�|1��3�vZ��u��)A�?e��`��ߍ�����D�
�%�����_?��x?muA?fa�<,5z>	��?/�%�kˏ�G,�>�/�(;�X<=�-�>:-��4�`�&�Ӿ��þI=��NF>�o?�$�?�V?�]V�D�C�,Օ>�,?qd?�Q?�G?��"?+.���9?(S1����>���>}kH?��z?"�A?�>h���i���[�M>F<97Z�v������`N�r��=�Y�=��>�4�=~��=�$>:�<��W=/�Q>1��=Z��=�|�=��n��Y�갠>WY?���>	�>R'6?j���
7�Ȣ�x.?�2�=͊��쒾�4������>�i?�t�?�S?`Q>��@��?��� >6��>�~>l}Z>%��>��L�N�Ƿ�=�v>�`">H�=�g�9��J��C�����<T(>P�>�u9>��"���e>�V� 2���z�>�k&�a���7�	��R��0�很����>�O9?c(?�@>������cSk��I>?;xH?��7?3��?q�F>�~���-|:�B{'�9B>ɼ���0A���c��X�1�3�,��B>L͞�v����Fa>:��oݾwtm�"�H�n��`FD=���_yP=O��B$ؾVK����=_�>��	� �Ȗ�����.SJ?ENn=3���\S�퍺���>퉘>�T�>��C�����@��̬�:�=���>]U8>B"�����F�����7>��G?�/G?s�?�G��m�h�,�2��0�z�o�%�ɼ>u?2#�>B��>�_>j�=Z#��q��U�o���?�pD�>�?�p�{_K��R��3���7���>5|?�{�>�?��I?3��>b�e?d�?x�>2��>��ｘܰ�<&?���?纄=��Խ.�T�	�8�F����>��)?߅B�T��>��?K�?��&?{Q?�?*�>.� �/@@�_��>4c�>��W��`���_>˥J?4x�>
&Y?�Ճ?D>>�x5�̢�b
���~�=N�>��2?�0#?��?���>���>F�����=]��>�c?�/�?��o?4��=��?9B2>.��>���=*��>���>�?LYO?��s?+�J?��>���<�B��b���Ps�NpP�#��;	rH<��y=z���+t��0�	��<!�;W)��gj�������D��
�����;=��>��t>>���J3>k�ľ6n��� @>��#���m��Ϙ;��ܷ=���>��?�ޔ>��$��=�p�>���>O���(?ɴ?4d?�i;�b�xx۾P�N��k�>�B?�_�=T�l�������t�@�f=m?�]?O�W�������b?:�]?�L�t =�v�þ��b�k��{�O?��
?E�G�-��>�?��q?���>�5f��En����s+b�Y�i����=�L�><���d�K�>��7?�W�>F
c>͙�=#c۾
�w������!?g�?���?��?p)*>��n��5��*��o��v�P?T��>�W��ʬ(?m����^þ�����푾��
���׾�����5������M<���F�����<6t?�qn?�Y?��a?.�龎_X��^Q� �� �S�@�����nI�M�:��6.��j� ���O �����0�;(󕾓;�5E�?f�%?7��*;�>>7���z�����R>���>U��ߒ=��ν��<���<��x��'�XA����'?:s�>���>�;?�^�@�D�3%�7/� ��W�=�i�>/��>��>�
�<�QD��i���s����f��2Žc�u>�cc?	L?cn?�N��)@1��^����!�h�1�
��B>4�>_��>�V����P&�n]>��>r�r��	����	���~=ۮ2?d}�>���>�.�?�!?�	�Y����w��[1��x�<��>W�h?���>	�>D νF� �d�>��R?gQ�>�E>��s�E��{؋������(?6��>
�>$� ? ����#�����D����J�6\>|�?�A��-��0��>y_B?�>yD�|y�>��4>��9�Ht����<>{?�P�<�YL>�u����־@7�2�7�R�$?�5?�ޗ��E*�::U>ju#?�?d޾>L��?E��>�ƾ�ݝ�f�
?5s^?�JK?��>?r��>�p<ǛǽW溽��:��r�=͉>��G>��<N
�=G7�9[���4����<�k>K\=�{�����<�jɼ�+�;�<=�-7>Ahۿ�K�f6پ������g 
�`���²�6͇�"�	�����晾��w����<(�eV�Ozc��Ռ�d�l�-G�?$�?�/��6*�����򃀿����Q�>\zp��ku�jy��%����6��>��(]!�p�O���h�X�e�|o'?8ᐾ�ǿ����i�ܾ��?ٵ?��x?�g���!�VN8���!>/��<Cp��6��a�����οP嚾�_?&��>	L�+7��U��>h��>5X>Fo>��,�����<��?��-?��>4Fs���ɿXu��J�<���?�@��A?��'����%S9=���>�?�A>�2������ev�>�͞?�r�?==��X�$׼u�g?Co<S$F��j�8�=�u�=C`'=d�~/E><��>v]���B�6�9�;>Å>�&�����_��R�<�V>�ٽ�5��Vd�?R{������ �φi�۔�<�|?f�?�l�>�R?@O
� H��Fs��]�?^�?�<�?y�?�j��/J>-羀`^?��D?+��>��^�M�x��-�=�j=���p��p�8���7���>���=�Q��  �I��I��:8��;2��Lſ&!�����=�V�;㉽�p�/>Խ��e�;~����l��!ܽ5=�,�=�F>ES�>[�Q>Q>suU?��h?�d�>�)>�E����1׾�s�L�}���4����� ��<�����=��An��@�)���^ɾ=�*�=�0R�����K� �Y�b� �F���.?Fk$>�ʾH�M��[+<�mʾ����?��( ��;6̾T�1��n��ɟ?��A?������V������ ˹���W?_5�ʭ��ج�ڝ�=����5=T�>z_�=8���3��wS��?2?�1?����嘾�D(>���K,=�'?�� ?>��<`��>>V%?�w#�W~��rx7>�G>�>�.�>��>_������/!?�zW?�Z��e��sU�>�ʳ�4M��8�)=d�&>BK1�5f
�v_a>5Q~<�i���s/�І����<��V?eۍ>8�)�s��􃐾�� ��3=�x?@�?_��>�4k?I.C?��<���T�G�,p=�W?��i?c	>8���6�Ͼp@����5?n2e?��M>�Rf�t���/���;B?��n?�?�8��D7}������`���6?�v?�]�g���'c�HP�Ve�>��>mG�>�8�J�>�<?�6 ��>�����y4��M�?-�@��?4�;,l	�|�}=j5�>[�>6b>������_��+x��&��=�_�>���ݶr�6��z���4?Nz�?��>A?������=������?�(�?Hg����;���ec�}1��"���7h=���f����0�3��{ľ���X������Q�>]�@̆ ���>��6��Xݿ�mп����5����I��?	��>9%�b�����l�Iw��$G�6I�汍�ٻ�>�F>�p��F��WOx���;�����a�>��1����>caI�Gٱ��|��5
�;���>��>�6�>6�����?44��=Cп)����	�ͧW?���?�I�?ro?uC�;�Gy�1�|������>?V�o?_?m�˻S�R�6y*���j?�^���S`���4�(GE�]U>9 3?�C�>�-���|=�>��>�l>�"/��Ŀmٶ��������?���?�o�r��>;��?�s+?�g��7��*Y���*�/1��;A?�2>������!��/=��ϒ���
?M}0?�y��0���a?�j��_z�
�1��c�I�>�����7�hF<b^	�F0Y��s���^���L�?]*�?l��?���)�J$?�W�>[����ž���=S��>8�>�p>)���YU�>���S{9�l>���?ߛ�?"?"������`З=`?p=�>da?���>Ld�>g�>�]��C�A��%�=D�
>z�Y;ܾ?OOZ?�?W��=�����E�!�T��@���G�i2F��j�>J��?p�?�N�>|���N,>C
C��I��:���L[��k������a�n�`>/Co>��="�/���N���?Lp�8�ؿ�i��p'��54?*��>�?����t�����;_?Rz�>�6� ,���%���B�_��?�G�?=�?��׾�R̼�>=�>�I�>;�Խ����\�����7>0�B?X��D��t�o�z�>���?	�@�ծ?ji�Ӊ?��u���~��d%��喾K;/>WhG?�T��W=Y#?=+�|������;]���>���?U�?���>X��?;ʂ�:�e�׉�o)�>*x?3�.?󰯻�(̾��h>�k?,�޾�疿,�����c?Z�@�$	@�`?���6�޿���P�������M�=� >��!>�g
������Ot�j%m�����S�=P��>�1u>�N>�5:>�_#> �
>����p��/���!�� �?�D}�^Q��F�����ZS�����5������C �P�4��ý�XB�_h��w��SO�=�;U?K�O?,�l?�g�>d��y�)>SU��=�6#�Z�= ��>��D?,%Q?a�1?�Mg=������a��z�Ë��1���8t�>*�6>��>�I�>m��>n�;��->{|>>�{o>Z5>d�=��A<K�3=�fE>x�>J��>O��>C<>t�>
ϴ�S1���h�0w��
̽f�?����J�,1���;��>����t�=�a.?>~>���>п�����1H?I���;(� �+���>q�0?mcW?O�>��h�T��6>ڼ��j��_>:% ��}l�P�)�'Q>�k?�O>�L`>	
.��y%�0WX�,�S����>�4N?�'P�w���6�d�"g8���־��>Y��>�J�<��D��!�b�|�@����<�.3?v��>c:���̾�ъ�ܾ��W>B� >6��Z�>���>8��U��G_n�C�s��=x�y>$�?�
/>���=�-�>�y��W�Q���>Ό9>��3>��@?�"?��}_�������;�F�{>�}�>b9�>��>v7I��|�=���>S�g>�'��f��X��ݓ>�"O>>v�7�K�WU��o=ַ���6�=��_=.N�H;��?=�~?���(䈿��e���lD?S+?b �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��I��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l�6>�^%?��Ӿ^]�>�����C����u�S� =F�>��G?���>H�=k=�B�
?��?���f���w�ȿ�v���>D6�?�˔?)�m�����M�?�{��>�?�?�X?"�j>�۾-\��l�>��@?�R?捶>Z:��'(�F�?;̶?��?I(E>O��?I�W?|B�>�k�y�&��骿U���R�9>I><��>�,>q)ƾ/#�Ό�����.�i��$�[v>
D==�e�>�U������i�=�|��fξ 罧C�>V:�>%S\>�[�>ҫ�>�a�>��q>�ӼI���.�c �{�K?�?0���n�N2�<V�=/�^�c�?z4?V�E���Ͼ�Ш>rd\?�Ā?��Z?��>7���J���ɿ��S����<�K>'��>!�>�ˈ�)J>�Zվ�\C���>��>�>��z5ھ�����"ќ>=A!?���>���=��?q)$?��g>@˨>�;E��2��f�J�^��>��>v�?�3z?\?d²���-���������3?]�=QI>H΀?��?'�>���������;�A]�����9V�?1^?�h���?�X�?�eA?�3;?��P>]��G�Ӿ��i�p9�>�?$h�ߋH�Q�R�0�6??��
?F�߼v��Ϲּm'�)q�V6?/|M?��"?�$�e�]AǾ-ފ<P�����<��]�FM����>F>ӄ	=J��=�Q*>��=r4�ћ<F��<��9>΄�>~>��ӽ�Ԉ�}:;?����D�=��b��2]�5m>��_>��;F�A?��&=��D�&䐿�{��`@;��?ך�?�J�?��˽�J[�� ?�(�?ȨG?r��>
�龚�ھ�;�������4��L���μ��>1�=�N��P����ᶿ*�|��)�>���?��>@%:?8A�>J�>
@q>o$��������5�N.U�����G�"�'�������q�8�x�B��誽��i>�)�U�>A�?)�P>W"_>.��>|���X>}5Z>�{>%�>}˒>$>�O�=}����(��BR?Q���W�'�_��,���j"B?�ed?Y2�>Sxh����G���~?���?uk�?}v>�zh�M0+��Z?�F�>����z
?b1:=A���y�<�S��(������t��v��>J�ֽ�:��M��>f��[
?�?k�����̾��׽P��c�K= �?:�(?^��KxE�޸r�̍Z�-�[�����1��6������gq�F���u肿
����$��p�;�:3?Z��?34���;��Ƽ�n�s���3�	f>{��>�u>Y��>�U>*��:Q'��[_�t�KR}�c��>�v?�_�> �I?�<?4pP?�OL?4Ҏ>�Q�>�n��/R�>�T�;��>F�>��9?��-?&?0?H?�9+?6�b>,^������kؾ�?Ou?�'?�?��?�̅�n�ý>��V�f��Ny�;������=Y}�<x׽Yu���T=��S>�?���)p6�%}��z�j>��3?+K�>+X�>�[����}��� =}��>�=?^��>��t�������>]�?�a����<�'+>Л�=�/�Ӓ��Ns�=3����=V����%�"�B<#�=y��=���;��i;ul�;��;ޡd<[�?)�?��>�y>�	�������	�
E�=<Y[>��Z>�>DdϾĉ��Iɖ��ek����>$��?��?F�Z=���=6��=%ϐ�~����
���ž�"p<�?H�?�RM?M�?~C:?��?�>���'���E�������>?�,?Ѿ�>�����ʾ���x3��~?g%?&�`�q��b*)��C¾5�ս~>�N/�*~�&���)D�?��I������d��?5��?_�@�Դ6���E���E���C?X�>���>��>A�)�D�g�<.���:>���>5R?H��>D�K?�V�?�N?�_B>/L'��t������ּ�#>N$J?P��?W$�?�H~?XH�>��=��O�t�˾6��ﬂ�SD���r��6�=K�=\~�>���>��>��=j���]sŽf+�o4>i+I>I�>!F�>�k�>�qf>��&�#�N?!�>\������.�w����"=��X?��r?a� ?���S���+/�pQ���|>���?&��?=�N?ߜM�g~>������ྦྷ:�1��>N��>�p�>n�%���5>��`>P^>�.�>���2�`�]�#I=�x5?�!?b/�=��߿tV�V�,������Y�=.�����~ν����,�>�Ͼ�Ƒ���F��C�Ø��Tg��zǕ�u�z%���X?4Ƭ=��>{��=��=���P�M�<Y+=&z(>�1�o���� �K2A�y�ai����k=�<��}��{Y�?��T?�;?�SP?p >;��=��i��>r�1���>p7>��
==Q��!.��9վ6���]��諳����
���_ԑ=�-ٽ�$5>(@S>�e>��\< fM=��>�{>���=���=c�4>P�D>=�>��=<e>{ �=3{?��������ˋ�;.>��5?FT�>v^2>�����!?���>�
h�%R��n����-�?gA�?�?�?�?Ǿţ>
̾=������=0?`>s�>2*>���[y,?+5�>w���`����5��?'��?(c0?�����,�iI >�6>�>IS�u0�	�[�ZV��N�:�"?�9��˾G�>]F�=I������$=��8>\�a=?�!�B;[�C��=�}�<G@=t�J=}ن>�IO>�=�I�����=>�E=���=�O>t�j;i�(�$��.=>P�=pf>�$>��>�V?��E?^�b?Fd�>(\����pݡ�c|>�=��>-�=��]>P_�>��&?��7?v�A?9z�>}��;-}�>��8>��j���I������h���=�a�?��n?�݉>�y���R�|���^��i��N?Mtl?�?���>����߿޻#���-�ki���&�;c�=\t��Ԏ�J-�� �l4޽7�=[��>���>JV�>��t>��5>2�H>0=�>.�>�$
=�5|=�',���'<�q �VɌ=�ѐ��==�坼�p8�x;Y�K����o�4:֚�;�(�<Nf;�3>���>�c�>�!?����K߾_�>�I����e��ܯ�~hp���4�����#^��)?��|��`9>8�l>��������S2?��W>�ګ> v�?@Z�?�&���bM����������(&>`��=U�;��C�;pc�JJ��D����>~Z�>���>�Q�>Iz"��r?��)&=}u�D~2��)�> ���K@ּ�g��j����ܞ�(�g��M�;U2B?���	>;�?n�B?��?M�> 1���m�{~+>�7��K@;���s{��Ӧ����?�#?d&�>�����H�7 ھ���Ķ>y���^F�����&3�����	���	=�p¾c���rY�������_#�z�x�*��>��?���?�ƾ)s����Z��@�HU��`�:?'D�?)^�>�R�>�JM?P"Z>����K¾:k�=V݊?֕�?�L�?H u>��=�?��`��>[�?1��?\��?�|s?�>��N�>m��;5� >k����=�=>B8�=3�=�)? 
?	l
?a˝��	�7`����^��=�e�=
�>�,�>�r>�I�=	�h=�4�=@P\>�F�>1�>�ee>CL�>���>�Ģ�V���.?���=p�>A)?N~�>�=�����=��'�@s5��")����?�����;�噼��=�o��9�>0ſ���?��i>O�
�k�?�-���m�K4=>aoQ>��Խl��>H_>�d>��>���>��7>0{�>>X���@��>5 ��X��L��a?�������=̛��yI�=���F.�<�V^�=8p����
�q�7���@>�|�8>[��?��V���6��8�E鋽j��>G��=�!?��������>�?���>o�������⊿jlھ��?t��?�ac>��>�W?�?��1�x*3��^Z�B�u��#A���d�@�`�@Ս�\����
�^��)�_?��x?y�A?�֑<�Tz>ї�?j&���� �>�/��;��<=�E�>����;a�B�Ӿ4�þ�z�U�E>U�o?<0�?lP?�.V�h!!�s�>�?;�?��i?Qx?
?K&ƾv�(?u�*<W��>@I?�~a?	<7?�:?��<~��`޼X>�1�Wˠ�9����������N�=��=�\=��;�m<u�c<X��=#o�=�2>{��=��=���=��=�`>���>M?���>���=E#8?���Si�5���-)?V��=����AY��ˉ�Y���8���+w?Yi�?o�d?"@>^�/��LE��ic>��>�^�=�.>�.�>g�p�*� �X=ͭN>Z#,>���=���;�i��/L
�1_�������>��>7�>yb�m�z>�T��ء����>���=5�q��+�S�0�\f=�B+��>��>��D?A�??��<Qs!���$�r�v�̳o?��'?5�1?ls?��P>MC���C�%�5��7>�9RH>lp��'��|��:\����J��T �{E
>i�d�l/��D�b>b��{�ݾ~n��I�!I���H=����U=yW�:�վ�����=e�	>����\� �#��Q���o
J?��j=�T��?U�3.���<>e.�>|��>G<�9u�1.@�8%�����=)��>6;>G���XG�e%��͆>9E?l�^?�o�?����@r��MB�t���I��A���?�Ϫ>?�?<�@>�ί=8����`��Ld�F�^��>���>��,�H�w��IT�n$����>�?-� >Y�?u�R?A??�_?�<)?�?�ˑ>𩸽���?&?ۉ�?9܄=��Խ'�T���8��F����>�})?�B�i��>�?o�?;�&?��Q?��?��>�� ��@@�>��>a[�>��W��a��g�_>�J?���>�:Y?�ԃ?*�=>Ԁ5�X墾ĩ�)X�=>>��2?�5#?K�?���>�a?�¾��=���>�,C?>^?Sb\?�D{>�
?ޜ�=�? ��=�3@=V�	?;�	?�]?��r?��U?�b?�3==�8网�_��\���>9=K�S�d!B��i�=LH����ʽ�e(=�{	>�h����l���}�s.���G����}���Q��>�e>�E��/�->��þ8
���dB>ͧ�!�������N�+��=?�>)�?�8�>�`�=���>���>	����%?:?<	?�*7�{_���ѾY�E�7P�>��D?UY�=.�k�'啿�Vm�I�z=#l?/�\?,�Y������b?W�]?�h��=��þI�b������O?�
?��G���>_�~?��q?���>J�e�/:n�^��pCb���j�sӶ=9t�>�Y�)�d�_?�>��7?xP�>��b>11�=q۾�w�%n��?��?� �?G��?�,*>C�n��2�>K��EՑ���]?�w�>���!?�o��Ͼ%c���Ԍ�� �nI��O��p����"��n%�<⁾6�ٽ��=�?s?UMo?�a?z: ��c�	\��~�VV����[�گF���C���B���l�.b�/��������@=����y�B�a��?�&?��Y��N�>����$��/���f>�Ǿ/}��3��o��6�3�x��<���
M��!���/?��>�W�>G�`?#�X���F�~�?������$>�2�>�:>��>a��މʽ�d>�{J���W�|���J>��T?��Y?Y$j?J���
�)�<.��[���F����&�i>�A!��{>�/����9�N����K��v`�/��������i�=��+?/��>���>ҿ�?��>���,���K6���[=��>bd?�+�>L>e����)����>h'??�y?���>_���OH��%��=Ӣ?Qd�>��%?���>� ���_�m���-���?�b"��?�'[��Wc�t��>d�;?��`=��<=8�>�Sǽk�%�@���F�@���@�>#w�=z;
>�碾�,��h;�"���j.?��?D ���Y$�.��>�z?���>hS�>Zw?���>귤��u�<6��>>`?�.I?��??C�>�p=;����ѳ���1�Y΃=�t>�Yh>6�=>є=�� �F�g���/���=�F&>�]��3��e=�B�;�I(=v@`=�
>7kۿBK�4�پ[���m=
�Ո�߲�mt�����Id��{���ax�z��08'�� V��(c�����
�l����?�:�?����q��б��!���Q���c��>�q�,���૾}��*����a����e!���O��!i���e�|�'?ȵ���ǿج��}-ܾR! ?k@ ?��y?��ͯ"���8�ř >���<���_������M�ο\���u�^?#��>�x�����>���>��X>~Uq>:���؞����<��?��-?]��>
kr���ɿň��a��<��?��@��A?}�(����{�U=���>`�	?'�?>t1��B�x����d�>�:�?���?�M=��W���	�~e?3<z�F�)Pݻ�+�=3>�=��=����zJ>)Q�>:z��_A��ܽ��4>/΅>R�!�8���^��˽<o]>�ս�W���΄?Ў\�!f�j�/�Q��.H>"�T?NA�>7^�=`�,?�8H��Ͽl�\�>a?�!�?���?�)?����O��>��ܾk�M?1E6?v/�>�x&�?�t�N��=�ἷٚ�����V���=Ɠ�>��>�x,� ����O�j���._�=N��ƿ�$��|��_=*�ݺ �[��}�h���S�T��#��/fo�ŉ�Y�h=g��=�Q>Ml�>u$W>-3Z>�fW?J�k?O�>��>}5�Y���ξ�-H��H�����]���죾�R��߾x�	���������ɾ�.=�t��=w�Q�ڔ��� ��b�&�F�k�.?%>Եʾ�M�<�)<&Eʾ�^���<����0m̾G1��n�W��?�6A?���:W�V?���	��5����W?��������b��=�Ϸ�f�=�ś>��=-��:�2�QBS���3?�A?�������&>� 	��=*R.?q��>�0<�Ͱ>��$?m�1��սzV>hp:>S��>^��>�l>JD��DPͽ�~?�}T?|���'ޞ�@��>U���Y���{=��	>,><�F&�,X>F^L< �����
����a<��j?}H>�d�V)��y�� ���=h��?�4�>�8�>Es?��B?�S6�`�Ҿ�H�C���=z�S?!�n?|	>�S˼a���{�6�,?Y�H?f9>�QU��F�����A�辊Y�>��?a�?�-��|����� �	�֝?�\k?E�n�����K�"�I�`�s�>	��>%��>�a6�`��>eo.?J�H�����h广cz:��e�?��@�$�?"���{�;	?�<���>��>_|��X���4�)���]�=��?��Ӿ���h>��T?��?n?�t�I4
����=�ٕ��Z�?��?���5g<��l��p�����<�ͫ=G�oN"�!����7��ƾ-�
���� ��T��>Z@WZ�,�>hE8�T6�TϿW��$[о�Rq�)�?��>��ȽԜ��D�j��Pu���G�_�H�����2��>L�=vaZ�����T�����z<���>�G=����#M���ݸ��k�_gZ=�Q>�م>֕ >� >֪L�l��?�8�����Ώ��&��5?� �?��? �E?VX�>���<{�/�����/�J?�Z?�s?P�|>Z��p��>��j?%f���H`���4��AE���T>�3?,W�>��-��|=Q>_��>Tk> /�L�Ŀ�Ѷ�;���	��?��?vu����>�}�?�w+?�a��3��1K����*�<�6��>A?�2>I���8�!�)&=�ϒ���
?kq0?�w�3�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�#N�����Xe����@y����?N^�?i�?ֵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�ض>@ �?~��=MH�>7��=�I���d���">e��=ߒ>�4z?�M?�k�>���=�7�/�	MF�IR�?��C����>H�a?�iL?3gb># ��*2��!�X(ͽ�z1��3���?��S+��޽Ӂ5>0�=>�>��D�QӾ��?�q�H�ؿi����'��-4?{��>2 ?N��a�t�6��3_?<p�>�3�j)��z ���7���?�E�?��?D�׾\M̼��>8�>DG�>`�Խmޟ�r�����7>G�B?�NH����o���>h��?׵@Ү?X�h��>(�1����������tT����w65?&��:�[>C��>���=�k����*r�����>\�?�b�?rr�>��t?lg��I�f®����>ɹw?�?�'ǽ��׾ɞ�>�x�>���3���6����2Y?m�
@4@�AH??���԰��s.���<D�����P��=H�R=zS>?���|@>l
X=b�J���@=bT1>�>#�p>��l>�>>��O>���=|��<�Bk��Ѩ���^P�J:��T5��Z���+����g�s� �Q3Ծe�׾́��?��RؽE)����u<�Ľ�͜;cj?ZI?��`?G�?�r'>ݖ>���vH���8�U�=��>��=?<�]?lM?���<#w���_f�,�a� ,���/{����>(�Q>���>�h�>Rڑ>�V��4>�7>��>)�B>�դ=��V=��=WzR>��>Jf�>gb~>�C<>��>Fϴ��1��i�h��
w�k̽0�?����R�J��1���9��Ӧ���h�=Hb.?|>���?пe����2H?%���z)���+���>}�0?�cW?�>��q�T�6:>7����j�5`>�+ �{l���)��%Q>vl?ٯF>�y>��3��7�-eK�樾K-j>/�0?����=u<�%�x��H�\��K>�L�>��W�����*��L���s�/o=�]??�U?ލ����3�o�i����QF>W�_>Ѕ=���=��U>� ~���@CI�i =W�=�`R>��%?w=�1:>��>5iľP���YlY>�<�>���>��<?:'R?4�=O6C�`p�k���8>9��>�B>I��>�mL��i>��>н�>��\�����϶�D��5>�c$<{N���A�̣+>�yI�+`='Lp�w�W���V����~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>J������ݲ���t�Oo)=�r�>yG? ���u��>B�ڛ	?s?-��g��-�ȿ��v�3��>}O�?[2�?��m��o���1@����>���?(NY?�<j>cbپ��W�b݋>�FA? �Q?+I�>���P(��g?�?U?II>�t�?=�s?��>�Uy��l/� -���t��X�=H!y;���>�I>����eF��Ó�q��h�j����b>�5%=��>���>���@,�=����L���c���>Yq>t(J>�~�>�� ?�O�>G�>z=�艽‾�(����K?X��?��|n�#�<�y�=1^���?x4?�Z�i�Ͼ�٨>ԭ\?���?[?<�>F��!6���п�'g���ޖ<D0K>���>�;�>����K>u�Ծg�C�`;�>@�>�8��@ھ�2��:E��g�>�n!?��>J�=��?���>A}�>:�>�JQ�������V�Ͼ�>v|?Q(?��?W�?���A����F�����v@�=�z?�~? �>��X���������\�	␽��?�d�?�{<>?�_�?"�1?8$?�=����ǚ� �9���>{?����B��X�Bw���V?�n
?=��>	���
>��T7������N�?r�]?rN?n��d�^�����Jq=��vB��K�������l$>�>3��� �=B>���=�K��5�N�<�4�=WD�>P�
>Z1-�z䶽��?p�Z�����F���Oy��01�b�->Bb�>߄^���g?#�����V���*4��Y�&�׼�?��?�G�?�	���o�#+l?�|�?&�D?Zx�>�A��.cʾ����7
�͉��:(��<>�է>D��=7���<���㩿ڢ����Ľ#k@�3�?S�>H�?��?�P�>�{{>ܪ���A� ��h��YY����"�2���_2���	���.���W�,ד�`&ҽ�x=8�*��<�>v�3?�O�>��>9�>�����=W�>�a�>���>uw>��=E�$=C8G�K��.|R?I���n�'����I�����A?fAd?tU�>;�e�iu�����/?Bh�?h[�?Z�u>�:h���*�Ry?8��>�~�u(
?��9=��)#�<�|��H4�7��3p�擏>sԽ}:��uM��3e��S
?�q?r���̾Խis���AD���k?��k?;�ϝX��7�N�D�>�f���=ߊ�:{����&��o��6y��솿~&g�V�(��.Ž��@?ovu?3�վ��ξ-{��ԁ�>M�����>��'?�c�>��?`�>ݤ��~/5��5'���.����<?Q�?��>��J?n�8?�7O?��L?,d�>�ح>}���Zo�>~]�;S>�>O��>�B:?�/?N2?S�?�o)?h	Y>����/	���׾C?h�?�S?Eo?-0?�ˊ�L�ǽ�����)��q��`p�$�=lh�<4�ܽ3�|�ϾM=%�N>��?k�=9��K��u>�9?^��>=��>��\�~�ͮ<�<�>g�
?d=�>����q�)q����>���?����y=� >T˿=]mv�n�T;���=�vμ���=Dp��h�R�f<1�=�G�=!s�:~��;
�<c%�:��y<jm�>��?Ǥ�>}F�>�V���� ���L��=�OY>�KS>�U>b,پ�t��%#����g�by>Vr�?�n�?k�g=�5�=��=�h��$t�����R�:��<�?�V#?�ST?擒?V�=?h#?��>
/��@��O�����|�?�%,?��>����ʾ�憎��3���?�^?�;a����_4)���¾��Խ��>�Z/��+~�}���D�,ڄ�����X��R��?保?�A���6��q辡���,[����C?u�>[J�>H �>ؾ)���g��(��%;>���>R?g�>`�O?�0{?ͣ[?�wT>B�8�z)��HΙ��i4���!>�@?���?J�?#y?w�>-�>e�)���S?�������(삾�V=wZ>8��>)�>�>���=�ǽ�+��;�>�ュ=��b>���>㦥>� �>�cw>�ݮ<�F_?0�>�=��T���3��0���P���y?9!�?/?ʴ=���
R��e����>Q�?v
�?�-?��z�>�����⊾'bp���>�O�>:w�>�|>	�<�4>�w�>:��>������nd&�Rm=5)?�9?��=-Pǿ�S[�äa��A��U=�.e���y�~Q���I��e�=$Ͼ2<!��{����K���˾�㌾�4���ľ'��K��>ѫ4��L�><�>љ�<*�!�/>�=צ���U��C�=�C��P�=�D<��V�����1X�Yp�;p7>=�n"�� ˾1~?�lG?�"+?�^D?W�}>�*>�J>���>9��tT?�X>e�E�F���1�5��G�������Dپ׾>�c�kR��b�>߽O�L>�92>U��=�(�<I��=�Dq=�=^V���=��=���=���=?��=�u>�=>Q�e?vʐ�џ��փ��PZܽ��'?��1>�],>X���NqO?}�)=����N����q�t�]?ϧ@R>�?�/?���@��>ഌ�iS��R�=/��9�=��=�ԃ����>�&w>�_�P���@{	�WԹ?
��?]/ ?I5o���̿AQ]>As:>m>LR�d1�Z"Z�zPa���X�B�!?��:��.̾��>{f�=P|߾��ľ'5=��7>�'d=4Z�.*[�(�=�Ky�Ue:=. n=Hȉ>��A>��=b������=�J=� �=��O>03z�Lk<���.���0=#��=�
a>w�#>���>*�?�90?�c?U��>�zn�oϾ������>��=���>xO�=�?C>f&�>��7?�D?]�K?Ų>�f�=?��>fa�>Mx,���m�������3�<$��?{��?��>�p<�q@�l����=��Ž �?�1?�?��>�U����9Y&���.�$���z{4��+=�mr��QU�M���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=$�����<�vż�����u&�:�+�1�����;r��;B�]<^��;���=.��>�Q>Y��>���=�9�����=^Ul��U)��K0=I���X�vI�%$��������ک�=�>{e�����$KT?�P+>�܅>7.�?���?�$\=P� ��6������l����e����6<���K�>��q�1�Q��־�L�>��W>���>�L~>W�0��_G�6���J���h���>"��}��d{����j�I��角��h��?���f=?�<��$U>#�o?-_??��?�A?/R��B�����e��9-����?�KN^��B2��3%?��"?��>񮑾Yw�X�z�J�p��>G���_W�����~XQ�~B�=혾{?�>�[��M��=h!��˓�ޛ��i0��F����?u�$?Dm�?H�œ�J�c�Ԇ%��?M��a�>�Rf?���=mT�>��	?_��| �􌹾>��Ub?���?�?	3>�T�=0���Uv�>Q�?}�?<�?��r?�T��*�>V�<���=�r� >�$>.r>���=���>���>At?.O��$� �,���<���jfM�4RD=��=�>��>�wj>�5>h~�=0��=� P>^=�>�Z�>;	}>���>ggl>�޾�S�aP$?�	�=#��>b1*?l�]>�{����\=�4�ĵ$���E�!;��`qG�5�n<N�:;�VU�t��x��>R�ǿϡ�?���>a�����>=Xz���ƽ�=�>Ȃ�Z�>U;[>�G>��>�Г>��>>WΒ>8��=Ɍ;��=bm��-;�D���q6��ξ�O>l���[޾G���G`�)���¾w��\d�6��}\���UB�z9�?7�b��Z��§<�\�x���>�ר>	2?����<��8(=,	?%L�>}$ƾ(��O��֪��c(�?��?d;c>��>Z�W?)�?7�1�3�vZ�
�u�l(A�Ze�@�`��፿�����
�����_?��x?yA?;P�<:z>B��?��%�]ӏ�*�>�/��&;�p><=+�>p*��Q�`�;�Ӿ�þ�6� IF>L�o?%�?�Y?	TV���־�'?�\%>%��>.$�?4�z?c�r?����p�>n	>6�T>|�K?9Af?��`?��s?���=ZO��nþ3�fŽ�ှ��>s%۽�o,��Ƚ	�=R�;Ӧ >]==Ek����b%=1�$�#��(=5=�OO=P��=�!�>�h]?nU�>il�>��7?	,�g`8��K���#/?��8=(I���Պ��'�����%�>��j?���?�dZ?e>ۚA�2�B�Y+>�r�>�{&>��[>/�>����F�+ɇ=�w>�u>��=s�N��⁾�	�Ɛ���;�<d�>4��>��y>�݀��,)>d����}�eb>�WL� ᷾�YO�iE�V�1��q�[�>��I?_3?���=�V�Ȋ���-i���(?�I:?N�K?�d}?g,�=ȾܾGl9�1gI����Қ>F}H<t�����������;���ĻDKu>�Ӡ�����"�a>u��W߾�Zn�J�I�r���TL=��IW=�H��k־&��
�=-�
>s���� �5��ت�R�I?ļg=A5���2U�p��U�>�q�>���>�;���v�|@�̼���=*<�>;>Q������;\G�^�B�>�F?Q`?f��?��|�X{p��D��������0����?���>�h?s�C>���=����>j��Ub��E���>���>����E�Ҥ���򾔴"�g�>B?��%>t�?7wP? �
?��^?X�)?ݎ?�	�>%��A䷾f@&?��?�=<�Խ�T���8�VF�F��>��)?{�B�&��>��?��?��&?��Q?��?��>?� ��A@����>�X�>�W��a����_>�J?���>j;Y?Dԃ?@�=>��5�颾����e�=�>��2?X4#?n�?ܱ�>x[�>+W��ܽ�=���>�c?�A�?�o?�+�=��?�2>~z�>Ft�=&�>[�>G?�EO?��s?(�J?�U�>���<5l�������Bs�t�W���h;y[G<�ux=h���p����_
�<���;����<�~���V'E�ٻ���X�;�V�>��s>)핾�1>��ľ�2���;A>eA��=g��Q���H�:��÷=>�?��>�d#��f�=���>� �>����6(?��? ?TM;��b��#۾��K��G�>��A?~�=+�l�r��2�u��h=@�m?#X^?��W������b?�\?O�쾪w<��¾�-g��d��M?9]
?�^9���>�~?�r?#Y�>)�m��m�����}c��c��^�=Kț>�t���d��ɤ>��6?��>9]>�z�=�۾Syw����/�?�?�^�?�ډ?�	 >.>m�%^߿o���x�K�"?�a�>���A�?^�N����-`�G#��cl
���ɾGIL�� ��Z�ӾE�L�R�F���������?Bs?[q?Y~?kپa.p���v���~�5CX�$�!6���j���p��Y�t�� �����*+��Ȇ�=a?X��
C�J��?-�9?s�����>���.�r���.v�>�k���)"�� z=���=Y��=�S=��=�	rm�C;�A?���>�e�>ZI?��P�RHT��?��)�㬦��l>B��>W�L><�>!�!�n����[C�,���׾���L��fd>�Zf?D�T?C�b?5�����*�I���le%�s���yﱾku4>\�=��t>r:3�����,���C��ii�p������x����=<�*?Ρ�>aģ>^ӑ?�}�>+3
����DF��Sf+�K��Ļ>�0c?$a�>秙>�]��.����>�\?!�?���>)�쾗�!������#��|?��?�} ?b:�>g��?�J�ާ���h�<��[���~�?q�;�̿����l>�� ?���=��a�,�}>��C���3�cxϾ+Z��� >-,?�=E��=Ҷ�����og�/-Ծ�?��?'�� z"�.h�>�-?���>�w�>;a�?ٛ>�Ӭ����=��!?N�r?��`?˻F?2d�>�H��'������Hg$�͊�<��}>��Y>���=[ƽ=2���eS�����$f<S�=��e=�A�]u�;�e��{��W�<� N>�jۿ":K���پ��`��H6
�\�B���/^�����#q��� ��Cx�{��݁'��(V��,c�������l�q��?9�?�k�����箚�*�������~��>x�q�B��{﫾��d@��)��3Ǭ�Cf!�;�O��i�F�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@��D?�(������E=a�>vx�>crW>vB��&�9��&��>_�?��?k2�<K�T�l�$9�:h?]�:�a�C���;�i�=��=��=��&H<>ˤ�>�	��7����4>>�B�>ջ�����o���=��W>~O��#F��5Մ?-{\��f���/��T��U>��T? +�>P:�=��,?W7H�`}Ͽ�\��*a?�0�?���?&�(?5ۿ��ؚ>��ܾ��M?_D6?���>�d&��t���=�6�����y���&V�}��=[��>b�>��,�����O�J��M��=����?����+�cD&�閴=4�=z� �������"�R�k� î��E�wnP��d�=�g�=WsN>��>.�;>�;�=�S?�g?I��>��L>ː��J��G�3���ܓ�S�,�o�����C�oy���F�����W|�ڗ�����g���E��n=1CZ��I�������^���D�w�*?�.C>�����P�]�\Ⱦ;����|�:Ʈ��ҎȾ�2�t��<�?/�3?�胿��W����]��ܽ��P?���e��̷�N��=�oX��q�;ɜ>��=]�P3�wlR�Ĕ0?��?���~&��[�(>'��� =�C,?��?OoV<ū>��%?�m*���何,Z>�65>�j�>�P�>,�>)Ү�/�ܽrk?�XT?3�����=B�>s���+Sz�i�f=ٕ>��5��-⼂�\>v�<����\��R��2��<�#]?b�R>��о�������t=(}?�?���>�si?�[:?Y=u2Ͼ6�S�S�ﾑF�=v�K?�tb?Q��=�i8���Ծ�����2?��a?ɵ*>����1T � �.�-$����>j�_?j�?1���9g���{���z���`(?��?ar���`�����������>��?G1?�8T�:1����?��=U5��Å��oxE���?�N@wN�?�-�>җ=���=��>��?Z�������p�O<����2�p>P?'�z�}�,���>��| >�if?*kk?� ?��˽��5���>��u���?���?���_�����p��G�a�:> �%=�
����'��慨���8�۾kA���F�];�؅�>1 @ś����>�w�7�ڿ�ӿ2i����9~���8?�$�>���*#�z�E�t�z��>]���T����<���>BzS>�B���a�#%z�tE;���M��<?\J
=��>ѱĽx���x���=qH�>5�>���>]�<�Hž�y�?7o�[������P,�SY ?|��?�5�?G*1?2�=�^=�C�=�I�=tM?A-#?fhk?$6�=H����T|<&�j?�_��wU`��4�uHE��U>�"3?�B�>S�-�_�|=�>���>g>�#/�v�Ŀ�ٶ�2���[��?��?�o���>p��?ws+?�i�8���[����*���+��<A?�2>���F�!�A0=�NҒ���
?P~0?&{�g.��_?�Ma�_�p���-�/ZĽ5h�>!�0��C]�%G�&'�Ye��қ���w�G�?=u�?��?s���#�h%?��>�}��ugǾ0c�<̋�>�<�>YN>[F`��u>2����:�iF	>G��?Rs�?�[?@z���릿>>��}?uo�>��v?>AM�>˱>b�ƾc;���1)���ɻt3��>�>�'?���>o��=�7&�Η?��v���K�������M�;ڪ>�W?��9?��J>BaռD<R<�����(8��L�<�g���D�X�r��x|>�h�=9~h>�=FWԾ�$#?_=+���ӿ�`����Y���?G�>1�	?��C����==�	N?�|>Z�
��6���1���r���?1��?�?�|����i���=I��>U�>�+���=��Q���O�=JJ?L|�f����w�\&H>&��?N@@���?�k��{?R(�?ӆ�@����މ|��n8>�*B?�����=��?pQ�=Pk�v����儿���>�e�?��?x��>+b?��n��2��+�<X��>{�k?r�?&p =��̾��=��?�M;�˒�mc&���R?��@A�@��8?Rٓ�Eg¿%�m��x��d��U�=���=5&>����>k[�=|;�y���k->���>���>y�>9�->1v�=�'��w�p������hY����:�� �S���')��m���A��O+�����$�R������-�ɽcrY�~���{���L�=Irc?R�f?��s?��#?��>��>Y��d>�=d��/����>k�$?��:?��K?�Ym�����2�f��LM��ӯ�q?:�c��>լ�=s��>g��>)S�>}�T>6@>���>�~�>��v>$��=�� >�Q>��j>��>.?�ر>�<>�|>�ϴ�4���h��w��/̽/��?�n���J��2��oK��0���Q�=6d.?À>U��=пY���,H?� ��+!�h�+�F�>��0?�`W?�>e��G�T��,>|���j�D>_( ��zl�,�)��$Q>`j?�)a>
�r>U4��69��LP��篾
�z>o�5?\���Ƚ7�3v��7I��Rݾ��K>NM�>3�6��2�l얿�h�d�i��t=�j:?*S?�&���⯾pu�p$��)Q>\�[>}j=}v�={�K>�Rj��~ƽ�G�%�*=�@�=�_>8�/?ԧ��~�J>��>���J�⾐��>�z?�
�>�C??��??D۹>�/�<�a��L|��?�G?�8>���=���v�\<�j�>$�>�޿=�Խ�®��@���@>�+>����ο���W<#w>}5=�s���=�������i >�~?���$䈿���d���lD?T+?> �=��F<��"�D ���H��H�?r�@m�?��	�ޢV�:�?�@�?��7��=}�>׫>�ξ�L��?��Ž;Ǣ�Ɣ	�5)#�gS�?��?�/�Zʋ�:l��6>�^%? �ӾI�>g'A�跔����)?q�{�z+�>�J?�4������u��>�<�>I�ؾ�>��?ʿ�u��Z?�*�?�\�?�ڂ��ggV���>f��?�c?[ؠ>0����I��S0�>�\H?�:D?t�>!�)����=�?7�?�Jt?���>�Z{?>F�?�u�>�0]�'�$���z{�+u>�N�>�/�>�bR>���Bv��狿��x�8�u���H��>?E�=l�N>�kܽ��پ��a>�r�3k��ײ��-!�=o6>�6Y=�>>���>�'�>*n>�@�<h.�	���z���x�K?V��?Z���2n��Z�<I��=�^��%?�H4?�D[��Ͼ}ը>��\?1?[?}b�>1��\>���翿E~����<��K>�4�>�G�>�$��/FK>�Ծ�5D��n�>�З>k���9?ھ�,����pA�>e!?E��>�Ю=l�?��2?(�|>C?dCK�.��Z>��0z>���>��?q�r?c2?����k�/��]x�Cɝ��Tb��>T��?��?E��>Y�K�A�������O���f�q?1,�?l���?�}?�,?�D? �t����������혾]��>?�!?���A�	K&����J?�N?���>���y�ս��ռ���zj��E?,\?C&?���*a�U�¾�\�<�#�;X��S�;�C�%�>Ӊ>����7��=k>fİ=Im�`!6�g�h<p�=H~�>��=+7��V���n9?�mg����^�C>�����V��Q�>nS�>p��<?��;=u6�0���7T��-�Ƚ���?�A�?2�?��U=�c���T?Ǵ]?8?��>�U��b�޾���6,���V����2ܩ�_�>��;�"�Ͼ�����8��*���￱�;�� ?�
�>=?��?�Ө>D}V>n����D!�Q�1�����:��<�"7"�����[Q'������VK�M`��YRɾ��5Γ>~����>k?Oׄ>��B>���> ˛=��<���>Ů�>���>n��>�p>�>���;^W���JR?9���`�'���辀����1B?�qd?�)�>�Ci�������|?��?s�?�:v>G}h�Z++�:n?W7�>?���q
?�s:=�x��D�<	R��}��zH�� ��-��>ea׽� :�|M��mf��k
?+?�p���̾�8׽������= �m?�o1?lt
���D�Ht���a��A���t���'�۾�J�[t�ّ��p����+w����O�I��8?�X�?ܞվ�Kɾ �׾�m� i,��B�>Xa�>��>�e�>ļ,>AE	�%�G�(�=�O��>�х?!9t>�K?��;?��C?�YQ?���>�x�>�ʽ�/ ?���;��y>�3�>�M?�A?��E?�?C-?W�+>���"�ƒپ�R,?�?�?	��>Ȏ?��X�r��e�2<���i�	ٽߙ��K����c住y뼉_�=u�>�T?�f�i�8�)����k>�w7?�_�>���>"���!���E�<N�>��
?�4�>[ �iwr��j�}4�>J��?�I�w\=Դ)>��=����eź߅�=��¼_��=�+��X;��W <�=�O�=��d���z�/�:cՌ;
��<Mu�>�?���>�C�>A��R� ����.j�=�Y>�S>�>�Dپ�}���$��9�g��^y>�w�?�z�?F�f=�=��=s|���U�����5������<�?1J#?�WT?L��?��=?Rj#?��>E+�M���^��k����?v!,?���>�����ʾ��Љ3�ٝ?a[?�<a����;)�͐¾��Խ�>�[/�]/~����5D�:���6��1��?꿝?,A�R�6��x�ֿ���[��x�C?�!�> Y�>|�>K�)�p�g�p%��1;>��>hR?mZ�>�4N?�w?úR?9k>��1�#l���Z���e���1><�9?l�~?�
�?��y?���>N�>�,H�������a���h�0�����v=͢]>fo�>���>M��>x@�=���y⯽K�=���=lXo>���>���>���>��z>��<?P?h��>�ާ���U�Ǿv���T�<�(�?��?qp?NM�=w�Ծ|D3�p| ��կ>1!�?��?� ?L�V�*>fD�<Ö��)f����>_ǜ>5W�>��>W�v=S[�=2�>�C�>h��Y�B�?�
�;?��&?��=+�ӿ�XF�����K�uʉ>��=8� ����L�>,�=)-3��ᾚ�I��<���c�-�:�����J����>��t<H��=ALL>p�1>+��=��=�����н��w���<#�G>��R>�k=w�\�t᛼�m�=��= 3�<�,ʾ�?N?��'?;G?D�r><��=,5��Օ�>񣺽�z?��I>�都�n��*�4�ZͲ�)ʛ��ԾŁӾ:e������>rv%��:">t ?>�K�=��<���=�,=TZ=�� ���<v��=�=P�=�>5�>���=��w?枂����&gO��A��I7?)�>�,�=�HǾ�_=?�pL>Y�˺���	�-}?�>�?Y+�?^&?ΥV��a�>�����)����=�]����#>��=�H5��H�>��O>$y�EE���������?o]@�];?�%��r�οh�%>?�I>a�=xM���,��(j��?e�
D)��*?��4� վs��>_� > �پ�^Ͼ��<�L>:Ͱ=�q�4�W�[��=�	���]=|0a=���>�QH>-�=���X��=;�s=?��=%�b>�:=�+�!y#�5t|=��=��Z>u�>�	�>>�?��:?j
^?���>);K���'þ|�M>�WL<9�>;�Y�>л�>r;?$s+?�Z@?ǋ�>��8;���>t>3�G�#�Y�
��"¾^>K[�?<ڍ?��>J9>�6�������,��
<���$?�EG?u?��>��̑ٿz�-�>�5��"꼶@=U_B=z�j���J�S���4��t���R%>���>�5�>�=�>Pf|>v�#>�->�r�>]2>3�=8��=�}��JV�<����^`_=�Ƽy��<�����z;-$<d����ȼ<����)<dˢ<}�{�*�r>�Λ>��	=�
?�-�qG����R>*�j�8pV�����3�G�@�s'[���T����Tؑ�0BI=�0b>�x�����W?׳=qB�=y�?qʣ?)��=癿�%���x������w�Ļ >����#|��[��`]��*L���;��>��>�*�>T�>܏(���1��e=؏��1��?�>�7��u䭽�����wh������j����hF:?�t��!�">.mz?�H?�Ԏ?}��>$䦽rw�R�=>к��Yc.�}4��e�m5۽f$?��?X9�>��E�=��#��������>5��bsD������	-��=��7ɾ/�>x:���^�+�+�G��K���KP�C^��R��>�H?��?����K�#�[�F"�UK��r?{�|?��<>��>�r!?��߻�پ�| ��?=D-V?&1�?���?�^>?�=���=c{?��?�
�?%�?T�s?8��Mb�>�3=�	�=C=��>�>w�>tZ=b��>74�>�!?Go��E���n��|	�
|���=��>�̆>�X�>XZ>qG>�>U�C>PJd>�q�>>s�>gNo>��>]�f>c��o����>��/>B�>T�I?���>����9췼�:�?�y�����Ľ��6=\��=Q�0>�����>��ʿ�k�?�ɺ>bc���>M���H��HZ=���>��5�:�><�>`u�>Ϙ�>��>c�>9�>�L=#sѾE�(>?�'m���3��X��%޾��D>st�����1���g[�O�Q�cCʾ�s	���p��z��#%�e��<{��?�K�I�e��}0��Vg�0�>���>0�M?�W��n�!��f�>�v ?U��>�Ǿ#���\��)����?P��?��^>k�>�Y?�H?�!�[�.���[�B%u�e�A�T�f�i�`��!���򀿡��A�����[?�v?�4@?�G<95�>?&~?�'�9ɋ�S��>�`-��F8�+^]=���>�H���_��<Ӿ�ڿ�3��FO>�#p?g�?!?kZ�G�ҽWϰ>hTA?��?�{?)]?��F?I|��.M)?a�+>'�>K�?�N?��:?F�<?��>O��=���<��=:����l���p�����<��,����<���"\j=L��=�V*=;�~���:�✽?V�����=�Cu=CmF>�=H��>��]?tK�>ᘆ>2�7?����s8��Ů�;+/?9�9=������q���>�
>��j?���?�_Z?�bd>G�A�o
C��>5V�>�n&>�\>Sc�>у�%�E����=�?>�O>�ԥ=�JM��́���	�Ƈ�����<W#>ɧ�>�Hy>�l����(>v���q|�5�c> =P������eQ�SG�v�1��Du���>:�J?Ad?í�=���㔽Mf��)?gn;?��L?�P?A��=�۾:�:��K��!���>�I�<2���d��l���0�;�V�F���r>�ן�V�:b>���w޾\�n��J����d1M=z�֎V=����վ�+�!��=.
>���\� ����%ժ�!-J?�j=󁥾v_U�b��w�>�Θ>�߮>��:��w�΅@�/���e<�=��>W;>���X��xG�:0�䥆>xcD?.Jd?!��?r�T���q�cK�i����9��N�<�ͤ?��>�z?	6>�*�=�i��ނ���\�^�D��=�>�Y�>o"��XJ��X�������#�؜>�,?�[>�?Y�S?-?�Z?W�&?VH?�E�>Z��⯾*A&?���?��="�Խ�T�8 9��F�>��>ҁ)?��B���>��?`�?��&?�Q?��?��>&� �5C@�ϖ�>mV�>J�W�Wb��F�_>�J?-��>B?Y?XՃ?��=>�5�l墾D����Q�=>�2?P8#?[�?b��>}�>d����=�k�>=`?��?Hfq?�N-=
|
?���>���>t�=Nn�>�*?s�?1?E?6�g?c�;?��>(��<�W���,������b���������<�6P=��Ƽ�˼�d<1/u=[���P�^�=�ʻq��\-ܼ5�����>(Yt>`��?/>Ŭþ����A>��������ډ��8�'��=죀>�,?��>g�$���=J�>���>���P(?�	?SF?�Ms;VKb��uھ�N�xڰ>��A?�}�=!�l�~c���Vu��sh=pm?�R^?��W�W
��N�b?��]?1h��=��þ��b����g�O?:�
??�G���>��~?d�q?O��>�e�,:n�+�� Db���j�Ѷ=Yr�>EX�N�d��?�>n�7?�N�>2�b>�$�=mu۾�w��q��g?��?�?���?�**>x�n�Y4���������4?��>A��1
�>�˭���Ͼ;���g���ܔ��T���N���Ϣ�,|���-$��̙�@.����="h)?���?Z��?	�h?����X�S��l�A�[�̚\�Q��~� �C!Q��d��_�~K{�+���3����c�>~�<�$W���7��g�?�j1?�������>�;J���پv�;3>퐡���U�L2k�"���#�=(�=�1��.L����<�?�g�>G�>q
M?$�Y�D�O��H���N��A��g�=H�>e�>��>����Y+�Lyj�SJE��Mo7��'>1�`?�N?�7m?�0	�Q&4�i-�����,�����
 [>��>�3�>�YX���2��E(���B��wp�T	���������ܥ=��1?�>#�>yX�?]�?���.���Zfo�/��I�<Y��> �g?�Q�>�}>�}��"��[�>p/`?n ?ʱ>��ݾ�V��E����'�u�!?���>��<?2B7>�u�v�4�Er��;֐��Hg���X��m�?�%�M�Ǿ?�>4A<?�=s[�|��>��>��N�	z7����<�׆=�l'?�E<�܇=ۧ^�>]���������;%?S�	?b��E3!����>n�'?&��>K��>�M�?���>�������;|�?0�a?��M?�~??��>04�<�B���廽���~m
=_�>�s>Xz=�0�=T.'���o�Y
�X�.=�í= !��ѽqu.<1q��:]���(�<{�C>�ڿ0�J�M(۾&��SV�y�
�{u������^����
�NȺ���v��,�"`5���U��ff�7���=i�3/�?�3�?@p��f��K ��(����aԽ>c_v�٪���Ʈ��2�0��`(�C����!�1�O�g���d�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@ӗH?R�#��پ�H�DP�>���>�@>;�� �~�оT7�>���?���?�+n�Ig[��w=��^?�3=�<��S7<��=��c=��'=C'P�JY)>��>py��(�ٵ��>ȿ>dՕ��_�D?T�O�K=c=d>��!Jʽ�ϊ?�҄�nl�'u
��B`�g	>S�E?qM�>�s�+?�������-
���E?�K�?���?,:[?k�Խ��M>��;��Q?�-?�ț>�2��o|���ؼ�҆�s�K>�Ӿ�3G�4�"=T��>�q�=�(��8#�ӑS�b��s'�=�3���ڿ�^�;����?���_ɽ���v5��n��;@*�4����.��?*�	��=���=.�;>�T>�>�
t>h�W?pl?��>��>�e<v%k�^��?��������*~���ž	8R�YW�^��^Q�+���N� �� �%}��;=�X�=�(R�����T� �\�b��F���.?	p$>��ʾ��M��*0<�Xʾ�ժ��p���f���̾J�1��n��ʟ?�A?u�����V�������˸�<�W?wH�h���Ь�|s�=b��$5=�>3�=!��b3�wS��f=?v�?&\��o��"ʟ>��4�6��=��>?�)�>�]Y>+��>HT?���H�=�<�=��1=���>I ?ӑ�=ͦо�;=��2?�Y?HZ�;G�{�MU�>����F��7|>U�>��꾔#���W�>�,�<ݢھ��b==n��(���0k?�~?>}��>�\�]��_�e�>�͛?3d�>�Y�=\�N?S֑? ��=�p#��~J�f���&>�S7?XG?+��=վ�=84־4���RR?i�Q?<X>�7���e���;�ʑ��r� >��V?��u?ec�;�����f`������?ش{?tjo����n���g��h�>=u?u��>��O��3�>#�I?9�X������ܻ����6�?��@���?�^�5Gx������m�>��>,���Υ��V���P���c >���>�����"]�b0� ���y�@?"�?U�?�}�$�ܾϯ>�o��oE�?"��?�A��X�/P��&Af��J�� 7�z�.=�ƽ�������_%�����4����F��($�W&�>�'@�&�=�>F���Jܿ"@ο�����x��dl��xf?2 �>E�X<��u?i���Ǣ_��F�ur���:�>~�>���L��%`R�=��ʽ�o?!ꖼ:�)>�<������v�qI:�X>�g�>\�x>��=�4��K��?@s�ެ̿���`}&��B:?��?X�?��?	��D𩽼�x�D��<7�?s.R?�i?ܮ�=%�[�ˊ��j?�?��0G`�>�4�4E�o�T>+3?��>��-���~=Z�>{�>��>�.���Ŀ϶�O������?�u�?\x���>�?af+?@��#���?����*�����5WA?qG2>�%����!���<��ɒ��}
?�~0?E�J:�\�_?+�a�N�p���-��ƽ�ۡ>��0�f\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>c����8Ǿ��<���>�(�>*N>jH_���u>����:�i	>���?�~�?Pj?���� ����U>
�}?�w�>� �?i4�=���>o�=E��Q����#>���=��=���?K�L?TN�>��=�5:��x/���E��bQ������C���>��a?;�L?x�b>hس�A,,�2[!�o�ν��4�i`���~@���/��3���5>�N=>�s>�D��MҾ��?�o���ؿ�i��Gq'�q44?㸃>X�?"���t�m��k:_?�y�>N7��+���%��HA�{��?�F�?��?ʼ׾k̼>�>RJ�>��Խ����?�����7>�B?��D��4�o���>���?,�@֮?�i�� ?�����^������X!K>p5?=��SE>2�?����Zl��访��q���>��?Ah�?,�M>�By?K���3�e���N>d�s?7;7?��D�%�̾�5Z>k�5?g�ؾ�i����
�H^�?��@�@�.p?�w���ؿ#���7��W��d�9p�=�]>^�"����=��:�^�<�S>�{>g��>A6�>Zk]>t��=���=pla=������5���ϭ��o�ݻ��R���N���t5�۾��a���F�f|H�H��o��V@��^����]�즴=)�L?�H?�Pn?��>�ʹ<z:>�'��O�=_qƽ��
=/O>�w4?�;Y?Br#?� �=/x�V�d��;w�L���ĕ���>k��><b�>#�>���>�G˼�)>dV�>8i\>�o�=!֥=D�="Q"�y�.>I��>���>���>�C<>��>Eϴ��1��j�h��
w�p̽0�?���Q�J��1���9��Ԧ���h�=Fb.?|>���?пf����2H?'���z)��+���>{�0?�cW?�>��o�T�5:>7����j�3`>�+ �{l���)��%Q>vl?[f>�u>[3�=�7�
P��g���[|>�36?���N�8���u� �H�lQ޾@�K>.��>��&�Y��ɖ����Nh���q=P9:?��?R)������`r�������Q>B�[>��=>*�=��M>VOe� ���7#H�<�1=/��=��^>N?^�D>-�=�h�>=9O��`��߶>RnK>Ӣ>�G?'�'?_��(C`�X�6���=��]2>���>�>�>���=��z��,
>�>��>��/���J�����_����P>��-���陽}�&=W������=�M9=ܹ�v3T�eD�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ3h�>/x�nZ��n��v�u�{�#=ݨ�>�8H?:W��/�O��>��v
?�?"_�⩤���ȿ|v�<��> �?���?k�m��A���@����>��?�gY?pi>lh۾�_Z����>��@?�R?��>�9���'���?߶?���?�!~>�h�?��?Ж�>T��C��@�ƿ�m���l>>o�S=�%>��>��оت��e��e��5Pp�`,��?�=���>)���j���`=�&��LžI�{���&?_��>!��>87C>�?�޺>�K>��w=�D<3�r���ֽ��K?���?)���2n��O�<P��=�^��&?�I4?�h[�o�Ͼ�ը>�\?k?�[?d�>4��K>��E迿;~�����<��K>34�>�H�>�$���FK>��Ծ�4D�ap�>�ϗ>�����?ھ�,��/R��:B�>�e!?���>�Ү=�N ?��%?�{>
��>$cC��͏���M��>,��>]�?�s?П?� ����0���z����\�$e>�}?v�?
4�>t��������Ʌ�aڼ�� �xm�?�h?$	Ƚj
?P��?;�>?;RD?�lB>[)���־KZ��ʠ�>�I!?,��	�@�g%�^���?�?W��>���żҽ{��h�� w���n?[?�q&?�����`�[,ž���<�T���s�c&<�B���>ۉ>����?8�=��>�A�=V9l�l�4�P�Y<}��=5�>92�=$4�
ʌ��,;?�8��͗�A->Ҏy��C���=>��>�ɿ�<?�ʽ!J������b��i!��I�?�t�?e��?�V�`|���|?���?�&?EC�>U$���'�W�㾗�]����|8�3;l=͂�>,HW�'%K�g��e}��©��i����#��c?2?�g�>ok�>qG"?���>/��>@������#��7*�cPK����`�	��1��K��i��I�D�HIw��̾ ���߽>6��%�p>	-?m�>#">��?��q=�=�l�>�:>�=j�>&�>�k%=���=tl�{DR?�����'�X�辻p���&B?=vd?��>�ui�Ã�����1j?���?'q�?�v>o�h��+�Om?�>�>�4���y
?��9=a�
��>�<	��N�����KN�}c�>@�׽�:�hM��f�]
?!#?uӐ��̾��ֽ�L}��%>�nk?��D?����oH�T1n�?WL���F�8C&�)w��i瑾hl%��dq���H΁���{��).�e��=��2?(9�?DwѾF�]���O�M�f���>|��>�wn>q��>��>}n�q���Lc��fG�-������>$�?O�>	�D?7?��P?!I?\�>{\�>,'�����>k�/=���>�k�>�';?��7?D+?l�?fF,?U9>A+��u���۾ʒ	? �?]u ?AW
?�Q?���a�нZ��<�i޼�5��͵�}�=�?�;���m�0��=ɮf>�V?�����8������k>�7?���>���>���#��'�<4�>��
?�G�>�����vr�>b��L�>���?.����=��)>���= ���O�ͺDf�=/�����=󅂼�;���<}�=�=]�s��Ⴙmg�:�S�;�R�<&u�>��?֓�>7C�>%@��'� ����i�=XY>�S>�>OEپ�}���$��F�g�_y>�w�?�z�?��f=��=���=�|��U�����������<��?�I#?�WT?9��?��=?"j#?�>�*�.M���^�������?�!,?��>����ʾ
�҉3���?�[?N<a�߶�O:)�]�¾:�Խ�>�[/�P/~�=��)D�`녻����z����?���?BA���6��w�󿘿$]��z�C?�!�>jU�>�>��)���g��%�2;>���>(R?�!�>�O?�<{?Ԥ[?�nT>#�8�30��qҙ���2���!>�@?���?���?Sy?�m�>/�>T�)�`྽N������4Ⴞ,�V=FZ>]��>�"�>P�>���={ȽVi��'�>��m�=P�b>ό�>���>�>^�w>�D�<)N?���>>��~��:���И��$��1�?���?��?�Z�=�4����6�ˌ���>h�?5�?7�)?��I��>�҄�S��7o�99}>W��>���>���=/�=(k�=rR�> K ?O�#��S%��	3��<.�?ʣ1?Laf=x�ӿb�|�;�������Ѿn��A�V��_�t'۽ƅ>�#���*�T����`����蘝�Dt��|����돾ow�>��E=�>��d>��S=�ET�Xi�ri�:>!
����=B���������G�8���B-q=y?�=d�<�mǾg�?��Z?��?��C?���>��4>����H�>��u�fl�>�_>l���f���Q#��v���ë��󳾃���6�v�y����=��f��x>��=F��<���=&A:>�=��=��i=��=���=OV>D�>oY>�V�=�wz>�E�?�U�� -��E�&�>+�" ?�?ҷ�>\B?�9'?� ?�́�|�Ͽ.��$�?�r�?���?��m?2u�����>ܝ����m�>a��=�)�>�߼dy��M�>�N>���q�\�) ��	��?���?�h*?��c�@��p>>��>��=t�=��=:���u��:��_���C?�%%��a�_��>╛>r�ɾ9_�Pм7m�>޼=�����R����=���gr<Q��=3Bw>D'>�>�"�����=�'K=�=Ԛ>�3��O��tq<�<���=k0->]�/>�*�>l_?�1?P�`?5�>�r��GӾ����.�>�ٿ=K��>*E�=U�B>���>r)5?�D?�QI?���>�=��>E�>'�.��Dn�+z辝��Rm�<q��?)l�?Ft�>ֶ�<b-3�D����>��ǽ>?�3?�&?0��>����ǿL�h��Io�����y��(�t=���T�-<�0>T��8��Z��>{��>��>%>�6�=�$*���(=T	�>�!>Z����>�R/=�����Ю=sH>-�7�l�л��,��Xz��\�����	�Ȼ@=��m<(��=�R >Ғ ?��j>���>��>�4����7> F�t�?�ݗ�=Ϭ���L���N���:��36��u���n�>� >m��4��'H5?x_y>�=�>�׫?��?�%�=�F�������|���"��=bٽE*J=%�v=�����!�`6x��Zr�0\�����>�T�>��?"1�>��A�B����V�[J��:�=W��k��d����W�ɘ�W��M��_=>��,?)-��\*0>��?v�?9�?�?�;��WM�ZL�G�H�_�@�o�*��þq�5���%?��?��>UR=�3?R�r�����q��>!�=�����ț��_�N�~D>�������=�Gܾ�"�\�{���o���gBF�����|��>�\?q��?�>������G�Z��O7�����G>9? V�?`ӱ=F��>E}L?j��;�E���5ؙ=#TN?а�?%��?{��l�k=�탽;�>o9?�M�?~�?{l?䟍��r�>�]>��=0��1�[>dΠ>��=���=Y�?�r�>�?O
A�a`	����9߾�N�s��=5 >�6�>X��>��>
�">�0>"Z�=�O@>�Q�>��>|k�=��>I��>���	"����"?ۣ>���>��3?DԆ>�W�=�Q���8�<�����*^��?o����^z���v�=�6=�F�<�Q�):�> QĿS�?4��>.���$��>�������z@>�O>Sf����>�RO>��N>�>A��>N>��>_H'>3yӾ�k>�w��X ��VB�ՑR�Ӿ�`y>dG���$(�C�	�ٽ����I�ܐ������i����2�<����<΄�?�d���gj���)������?�X�>\�6?mˎ�I��pF>ԭ�>���>՗���z�������	�背?(�?�b>�:�>�W]?x#?����:���_�*s�G$@��ve���_�Eꍿ'�_V	�\�ҽ�Z?�@m?�A?�&(<`�}>SD{?m�*��똾b�>�8.���;��s=�i�>�*��ٰm�X�˾	5�������B>��o?!��?G�?`�O���*�0��>!��>�<7?wi6?S�y?�%?/�D�P?�-w>E?0;��?�p@?�3:?�>?��+>2e��	s���Z�>�� p��-�V�vFT���D�>x<��~=�մ�Bސ�O�;���=t{�m��<���=k�?=�#*=��=�o��tT-�A�>��[?D��>NՇ>H�7?i����5��s���z-?X8<=,Ƅ��s�����(�{U>m�j?K^�?mBW?��M>OT<�^>M�gW>>p�>J�#>��O>��>mU����D�3��=�>�>b�=�W���s�!	����N=�<
�>3��>ǔ}>�0����'>�0��y�y�Ϻf>�rQ�0̺�\S��ZG���1��v�P��>�6K?�?]`�=�c�!��5f��6)?O�;?6�M?.�~?�ۗ=�ھ�i:�!rJ�y ��p�>ˢ�<n��ⓢ�����j�:���jq>c����͛���>���� ��Q�o��VI�#"�����=S7�P|�=�Y��������=Q�=����`��a簿0dT?|��<J�־�C��1���MU�=뗾>�>-JŽX�����W��J�X�=���>�h>?[�<W��b�`�F�����~>�_C?��_?+X�?��z�d-k��<2�[M�˕��E�<�?ޕ�>d�?���>u(�=o�����?[��ZH�"�>O��>����,C�u�������&�6Y�>:��>Q�_>:?��B?!�?��_?N(+?P�?�q�>g4������"?�o�?ħ=on��b32��=�8�C�cu�>(�-?�
�}!�>�I?��?��&?P N?��?zq/>�.뾑!D���>2��>KaS�����R�c>��M?�{�>��[?/Ĉ?I�9>;�����X�ؽ��A=��>bY0?q#?;?=��>��@?򸿾�B��|��>p8>?���?b@?BN�=��?�Q'<�İ>��>�H�>Z�B>��Q??t[?�G>?`\?�m�>��b;խ�5#���P��aE��6<m;T�䙽\9���(��`��P�	<L�$�X)>�"�<��=��2���Ž� �����>Is>�-���1>O�ľ�����A>{����ƛ�������9�]�=0��>}S?�ו>1"��M�=��>W�>��(?��?$�?�B;��b�5۾*�J�R��>�&B?N��=��l��]��Iru���i=�m?�^?�W�wu��O�b?��]??h��=��þx�b����g�O?=�
?1�G���>��~?f�q?T��>�e�*:n�*��Db���j�&Ѷ=\r�>LX�R�d��?�>o�7?�N�>/�b>%%�=iu۾�w��q��h?��?�?���?+*>��n�Z4��"/�zh��L�c?���>n��H��>1\>�K+˾�i�������ݾA-ɾtʰ�B+��(4þ��q�s���!���w>�7?���?�h?��?g=ξB@��VI�׾��M�V�u'�	V�V�<�{e��T�<��1�L��1��=���J�<F���6B�%<�?�#&?��3����>�j��<��o˾<�C>È������=Iև��E=�T=��g��m/�;���F�?gж>j �>�W=?�\��2=��1���7�\$����0>ǡ�>�W�>!L�>Q=\9��/�v���ɾ����Eͽ	�Q>�sq?��I?��m?�_9��+���|� X@�*�	���̾V~_>��>P�>j!ҽl*��;��'��=p�q��zڊ�*�^b�<�|>?�>���>^��?i�?b���ϾP}c��z�HE�=��>K�?G�>.�>�C�_��`��>	�l?���>��>-���aZ!��{���ʽ�%�>�߭>��>-�o>b�,��#\�k��?����9�Tt�=שh?򃄾f�`��>uR?'�:��G<�|�>��v���!����e�'�v�>�|?J��=Z�;>�ž�$�[�{��7��w%+?7?<��I�&�(��>�c#?��>�`�>Ja�?~�>N/ľ
c�;x?B�]?RGK?�~C?��>TX=�޲���ν�"��{G=��>�D]>f=��=5l��zZ�.V��(=_��=,�Լ+&���<zC�����<���<_*>jUܿ��K�RkԾ���_�h�
�M�����Hϊ�m������G$���Ȁ�-���ON�da�g�d�O/����o���?u��?����)��������| ��p�>4Ms�o߂�x������4޾uꪾ_&�(XO��9j�re���&?ۙ��ʿ�礿|$ݾKn
?X\?�nz?����K��B�E�=jA���q<e���Ě�oiϿa�¾�W?QY�>7yӾ>4�>$<>�>S��>�2�������#�<.4?�T5?:�>��b�>�ǿ1뱿�ֈ�2��?md
@�IA?��(��t�)t=�z�>��?�?>Iz.�������	�>)�?ɹ�?�2@=_�T� �ļ��c?O�6<8&G��л�=s|�=�.C=�����Q>#��>A���G�r����)>@^�>Ű��
-��c��y�<��Q>:��4蝽5Մ?,{\��f���/��T��U>��T?�*�>d:�=��,?Y7H�_}Ͽ	�\��*a?�0�?���?&�(?0ۿ��ؚ>��ܾ��M?_D6?���>�d&��t�܅�=�6���s���&V�k��=U��>_�>��,�܋���O��I��B��=)�1�ƿ.�$�Jv�t�=�p	��_�W������`�T�0៾P�o�/꽊�c=��=�Q>4b�>�!W>��Y>�hW?�k?걿>�v>=��$z��8�ξI���w��T���B��f��'���w�\"�Z"
�������ɾ�G��1=��F��M��|�&��b���_���'?6T�=��Ǿmu/�� <���3����u���P������/�|�r�r}�?5?����4f����/I�I��;,m?�r'���Ⱦ�.ԾJ/;=�3���=��>q=������C�ˍX�� 0?�R?v���͐��Y,>{����=8+?��?.D�<� �>�$?E�(������^>��5>Cʤ>��>C

>�S��+�߽�?�kT?ô���������>�����}� 9Z=��>mz-��t���]>;��<i�����SК�N�<��U?�0�>�d'����42���g߼?�O=iv?.?㧦>�j?�IB?�I�<R'��+O����>�=�}W?2�f?�[>��5Yʾ~S��ޘ6?=h?��L>�yi����a�-��"���?h�q?HB?��㼥Dy�/���w=
��+1?��v?s^�xs�����K�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�%Þ?��@���?��;<��Q��=�;?l\�>��O��>ƾ�z������'�q=�"�>���}ev����R,�e�8?ݠ�?���>�������;�=��>��˧?D7�?�c��1�/-���~�D��ِڽ7�����Q������9Q�֗־L-*�.޳�dB=��m>��@,T˽v:�>_*o�`�ҿ��˿�Ȝ�e����ƽ��&?o��>�zL�~վ����T9h�s'��=�~�˾eO{>D��=����骾����2;�
��>�>��s��>�6�Ǽ���Ⱦ����>�(�>/��>E������o�?����Oٿ�٣������K?���?8�?�� ?UT�=.Yξ�~ž?�����O? i?�ZR?�]ǻ�¾qP⽜�j?~^���U`�4��IE�U>�"3?D�>7�-��|=#>���>�]>�!/�w�Ŀ�ٶ�2������?V��?�p�A��>���?hs+?�i��7���U����*��*��9A?"2>�����!��/=��ђ�{�
?�}0?[w�7,���_?�a�L�p�+�-�M�ƽܡ>��0�+e\��C����#Xe�����?y����?*^�?H�?>��J #�.6%?��>����?:Ǿ�<#�>^)�>A+N>�F_�,�u><���:�#i	>t��?7~�?�i?ƕ������SV>��}?�#�>��?o�=!a�>d�=񰾈�,��l#>"�=�>���?Y�M?�K�>�W�=��8�v/�_[F��GR�-$�5�C���>n�a?��L?Kb>{��($2�u!��sͽb1��G�MW@�Z�,��߽�(5>
�=>�>T�D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*��п�/��dX������C�=#qm=N5>9⽜��=U͖<�*�}M��S>f�>Z%�>KG�>τE>�oH>ǉG>g ����%�ӏ��i����@�i�wj���r����ǘ�����Ͼ� Ӿ�������ձ��/V�r�'��+�=y�S?k�M?H�?c��>����I>�P��2���=>���>l�.?�^]?ٴ?�q�=UU�`V�IO~��
���[���'�>h��>�?�>��>
��=j�>�o>i*�>��=ud�=r�ͼD�=��:>�2�>�T?�ɻ>�O>G0�<𡾿�w����W�]�������??4���"���������&>
H?':a�{䉿��ؿL~��
F?��u����\��"6>��?��O?AO>7��fў���=�2'���~�{P>��s���Ƚ�Y���=�)>?���=��>kI$��gH��F�M�����>@?�q��sq\�0ts���G��ѳ��+a>A�>	]��a,�I}��B�f�<r�0��(.7?3��>%?(��ѧ��[��㗧�eBk>״�>�r�=Ls=�T�>f!s�P���� ����=�f�=��G>�6?��>ؚ=��>�����r�-R�>��C>fM>�I?�o&?�����B��j������3�>���>�;�>�>��&�u	T=�9�>��> �<uj�<�}���J��>f����tP���<�>[4޼!S�=��=-h9��z� .\�!�~?���,䈿���d���lD?V+?Z �=W�F<��"�= ��yH��@�?n�@m�?��	�բV�H�?�@�?S��8��=}�>�֫>�ξR�L�ٱ?��Ž.Ǣ���	�;)#�YS�?��?��/�Rʋ�*l��6>�^%?�ӾOh�>xx��Z�������u�_�#=T��>�8H?�V����O�j>��v
?�?�^�੤���ȿ6|v����>X�?���?g�m��A���@����>;��?�gY?soi>�g۾A`Z����>һ@?�R?�>�9�}�'���?�޶?կ�?�>� �?�2x?�W�>�<!�1'�貵��l���)���,�9��>�H>q,߾َW�:*�����n�P��t���>��!=��>E��e���B>��Z�I���B���cv`>��O>���>�7?ox?�H
?_U�>{�=��>avr���Ⱦ��K?���?,���2n��N�<[��=(�^��&?�I4?k[�|�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��M��<��K>)4�>�H�>�$���FK>��Ծ�4D�dp�>�ϗ>�����?ھ�,��8S��GB�>�e!?���>�Ү=ۙ ?��#?��j>�(�>CaE��9��X�E����>ע�>�H?�~?��?�Թ��Z3�����桿��[�r;N>��x?V?rʕ>b�������vkE�9BI�6���^��?�tg?wS�0?<2�?�??a�A?~)f>և�(ؾo�����>$�!?gm���A�V3&����:~?<Z?���>�]��^{ֽ�ټ&���2���?_5\?LZ&?�q���`�X�¾�w�< �!�ӊA����;N�C�Λ>o>����
��=�]>�@�=.�m�xh6�h�f<��=i��>���=K7��I��=,?~�G�*ۃ���=�r��wD�s�>JL>.��٬^?<k=���{�j���x���U�� �?��?Qk�?�
��˝h�E$=?��?]	?S"�>�I��v}޾N���Qw�~x�/w�K�>h��>�l�S����ә���F����ŽDx�k�?���>���>��>2�'>!b�>h��������7�yV�Uv��Q'�~@�-��پP�M�p�S<�T�Zb����>�ʽ}��>i?�a�=�-U>�-?=�p=Ȼ�>چ�>Gt�>���>l(�>��>qe�=m\	>�&H���R?�����(���o\��6B?.[d?�I�>�k[�����eV�%�?�F�?bJ�?&�y>�sf�[*��-?�c�>�瀾C�	?��I=�-�j�<�j����r�������>݆ڽ-�:��%L�g�a�*
?C?cHb�>h̾Z�߽�I��B��ۃ?��?����@P�@z���;`�Z�W�3��$�+ԫ�30�RՁ�F�/����Ȁ�L�!��<���08?;��?���O̾�s��h^�PCI�So�>��>��|>� �>��>Ǎ�M���C�T|U�������>��V?��>:�D?2�:?lT?�L? h�>fx�>�
��~��>�����E�>�M�>�;?�Q,?�c+?�?��)?�}]>���W���!׾�U?��?�?,?�n?ebw��ᓽ�{��?�~���j�_������=S��<7/ý>�����\=��K>�v?z��L�8������k>�7?��>y��>B͏�Xh��Vw�<a.�>2�
?�^�>ٓ��:r��M�P��>颂?�E��X=�*>4k�=7���$����=Y����ʐ=v���Y,<���<�b�=ݕ=�)m��i���;O��;٠�<hm�>��?��>�:�>_2��� �������=55Y>GS>�>�Iپsy��/%����g�nny>�y�?nz�?� g=/�=�C�=���fX�����x꽾-��<�?!6#?ZNT?v��?J�=?�f#?O�>��,K���]����9�?s�&?kr>(`)�7E��/��9]�og?�?A����e�A,(�� ��ϱ���o>�F�k���z
��Oh��_}>��`3�==\�?4�?�GF�[�=�ņ��R������z?�>'�>E3�>���R�̃����="?��t?�׳>ouU?&�y?��[?ݦ6>�6�g����+���H'��F >�>?f��?�1�?07w?�Z�>�>9����%����'�t��ڄ��<��=W�h> �>�c�>�ź>���=����)����D�s^�=��>M�>y]�>���>!.|>0$<�/E?��>V����y
�y)���.��?=��+u? �?5�0?L-=q��B��D���S�>m��?�?��-?�<Q� �=S���ݴ������w�>i�>�y�>k:�=�%l=/�>ݿ>h��>�^����6��pW���?��D?���=�ſj�p��!n��횾c�<�Ғ��Rd�Ɋ��8X����=�䙾ø�Vt����W�����Go��궾�)���x���>^�i=Cb >�q�=��<��ǼV��<L�7=w�<��=T�e���<��/�y�λ�ċ���D��}�<�aE= ����˾��}?�3I?^�+?��C?'�y>Ɩ>�Z4�ř�>�����8?xxV>*O��8���e;�������
�ؾ�v׾��c�
ן�=m>�FI�0�>�[3>�U�=���<N�=�v=LJ�=�^��=z��=�J�=�ˬ=U��=|*>N>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�i6>M�>�R�]�1��U\�n_b���Y�ҷ!?:�:��U̾I̅>�=&�޾ehƾ��1=� 6>?�]=�U�a\�ט=UR~���==�j=j�>�'D>%��=Ѱ��ŷ=<BN=�y�=�O>A�:��5���*�U�7=մ�=Q|b>�]%>#h�>J3/?2C8?��s?�s�>�վy�����;��>]�>�a?V>��x>�
?�?MA?�1Y?Z��>[_<�0d�>��>���,�w��Y��v����6c�?L�?���>�^�������W6�%W�N�P�?�55?\�2?�?�>�U����7Y&���.�/�����4��+=�mr��QU�J���Lm�;�㽾�=�p�>���>��>2Ty>�9>��N>�>��>�6�<~p�=�⌻���<� ��x��=�����<�vżT���$u&�:�+�H���l�;��;-�]<͡�;
��=���>	:>L��>ɏ�=���L/>г��-�L�=��=�I��|+B��2d�}H~��/��V6���B>{7X>�p��r3��6�?��Y>�q?>���?�Cu?��>t �޼վ�P��4Be��ES�s�=��>��<�w;��Y`���M�2�Ҿ��>jL�>S�H>]M�<5<���\��u�>��Y��HN��3z>q����������!�E��ݛ�ۡ�����E�ьj?N����;/>�j�?A�5? ��?��?~�q�˖����>��ؾ�����vھ,�[�}�6���=?'�*?�?�[C���V�ɵ���ݽ�K�>�>�\�K�k���HH�`��=�þ�m�>�����þ4�5�����v�� mQ��)��>"%A?��?��A�SU��R�T�j��!���?�\u?��>�?���>ߔs���CVL���>�)Y?n��?j��?�D�=7�>�Fm��>Hk?7�?C��?�g?��+��>�EM=��>�҃�lB>&��=�|�=��1>.?]B?��?�\��������n��W�����A7�=Rϑ>Kۆ>y�j>��D>���<<)�j	>�ߤ>YF>'��>Z\�>�E�>�ݾ�=�V�?Ԝ���=`�?G?8>�4>>���Kl>=k��������,<�ƒ��;��˭A�BG����ʼ.L�<��>�˿VK�?�	�>��*�=�?A��,�/�GQ>T�g>��2w�>�k=>ۡI>�?`>��\>+�R>��J>tWZ>ebҾ�">�r���!��C��R�z�Ѿ��{>���3/$�(	�[*��NoL�Ws��t���/j�nV����=��g�<^�?�~��c�j��w)��!���? ��>|�5?:��Y�����>,��>�m�>��������/��F��Y��?+�?1;c>;�>U�W?+�?֓1��3�vZ�m�u�e(A�,e�m�`��፿���1�
��
����_?��x?�xA?T�<�9z>m��?��%�ӏ�J*�>�/�[';��6<=�*�>Q)���`���Ӿ��þ�8�GF>J�o?Z%�?CY?lUV��3�%*>X�:?'�R?Yd�?oZC?��)?�'H���?/55>��>�-?��W?LW"?C��>� ~>V
>�%<���6;��2�)�.�i5�(���x=b==�=]�=:+v>Z>=jt�{G���{�<�����=c�;�|<>_o>��>�y`?r��>��R>Mb4?�����H�WZ?nq�>�;@��Ѯ�߳���@���>�If?;B�?p?�Յ>Id>�&���di=[��=��w=��>�K�>��"�Q]����\<�[�=D�>'�=Dp�	b�$�������<?��x>��>�/|>#
����'>B}��u0z�٤d>[�Q�O̺���S���G���1��v��X�>��K?Q�?ژ�=K_��)��If��0)?�]<?OM?��?:�=�۾>�9��J��=���>]�<�������$����:�6v�:8�s>�2���͛���>���� ��Q�o��VI�#"�����=S7�P|�=�Y��������=Q�=����`��a簿0dT?|��<J�־�C��1���MU�=뗾>�>-JŽX�����W��J�X�=���>�h>?[�<W��b�`�F�����~>�_C?��_?+X�?��z�d-k��<2�[M�˕��E�<�?ޕ�>d�?���>u(�=o�����?[��ZH�"�>O��>����,C�u�������&�6Y�>:��>Q�_>:?��B?!�?��_?N(+?P�?�q�>g4������"?�o�?ħ=on��b32��=�8�C�cu�>(�-?�
�}!�>�I?��?��&?P N?��?zq/>�.뾑!D���>2��>KaS�����R�c>��M?�{�>��[?/Ĉ?I�9>;�����X�ؽ��A=��>bY0?q#?;?=��>��@?򸿾�B��|��>p8>?���?b@?BN�=��?�Q'<�İ>��>�H�>Z�B>��Q??t[?�G>?`\?�m�>��b;խ�5#���P��aE��6<m;T�䙽\9���(��`��P�	<L�$�X)>�"�<��=��2���Ž� �����>Is>�-���1>O�ľ�����A>{����ƛ�������9�]�=0��>}S?�ו>1"��M�=��>W�>��(?��?$�?�B;��b�5۾*�J�R��>�&B?N��=��l��]��Iru���i=�m?�^?�W�wu��O�b?��]??h��=��þx�b����g�O?=�
?1�G���>��~?f�q?T��>�e�*:n�*��Db���j�&Ѷ=\r�>LX�R�d��?�>o�7?�N�>/�b>%%�=iu۾�w��q��h?��?�?���?+*>��n�Z4��"/�zh��L�c?���>n��H��>1\>�K+˾�i�������ݾA-ɾtʰ�B+��(4þ��q�s���!���w>�7?���?�h?��?g=ξB@��VI�׾��M�V�u'�	V�V�<�{e��T�<��1�L��1��=���J�<F���6B�%<�?�#&?��3����>�j��<��o˾<�C>È������=Iև��E=�T=��g��m/�;���F�?gж>j �>�W=?�\��2=��1���7�\$����0>ǡ�>�W�>!L�>Q=\9��/�v���ɾ����Eͽ	�Q>�sq?��I?��m?�_9��+���|� X@�*�	���̾V~_>��>P�>j!ҽl*��;��'��=p�q��zڊ�*�^b�<�|>?�>���>^��?i�?b���ϾP}c��z�HE�=��>K�?G�>.�>�C�_��`��>	�l?���>��>-���aZ!��{���ʽ�%�>�߭>��>-�o>b�,��#\�k��?����9�Tt�=שh?򃄾f�`��>uR?'�:��G<�|�>��v���!����e�'�v�>�|?J��=Z�;>�ž�$�[�{��7��w%+?7?<��I�&�(��>�c#?��>�`�>Ja�?~�>N/ľ
c�;x?B�]?RGK?�~C?��>TX=�޲���ν�"��{G=��>�D]>f=��=5l��zZ�.V��(=_��=,�Լ+&���<zC�����<���<_*>jUܿ��K�RkԾ���_�h�
�M�����Hϊ�m������G$���Ȁ�-���ON�da�g�d�O/����o���?u��?����)��������| ��p�>4Ms�o߂�x������4޾uꪾ_&�(XO��9j�re���&?ۙ��ʿ�礿|$ݾKn
?X\?�nz?����K��B�E�=jA���q<e���Ě�oiϿa�¾�W?QY�>7yӾ>4�>$<>�>S��>�2�������#�<.4?�T5?:�>��b�>�ǿ1뱿�ֈ�2��?md
@�IA?��(��t�)t=�z�>��?�?>Iz.�������	�>)�?ɹ�?�2@=_�T� �ļ��c?O�6<8&G��л�=s|�=�.C=�����Q>#��>A���G�r����)>@^�>Ű��
-��c��y�<��Q>:��4蝽5Մ?,{\��f���/��T��U>��T?�*�>d:�=��,?Y7H�_}Ͽ	�\��*a?�0�?���?&�(?0ۿ��ؚ>��ܾ��M?_D6?���>�d&��t�܅�=�6���s���&V�k��=U��>_�>��,�܋���O��I��B��=)�1�ƿ.�$�Jv�t�=�p	��_�W������`�T�0៾P�o�/꽊�c=��=�Q>4b�>�!W>��Y>�hW?�k?걿>�v>=��$z��8�ξI���w��T���B��f��'���w�\"�Z"
�������ɾ�G��1=��F��M��|�&��b���_���'?6T�=��Ǿmu/�� <���3����u���P������/�|�r�r}�?5?����4f����/I�I��;,m?�r'���Ⱦ�.ԾJ/;=�3���=��>q=������C�ˍX�� 0?�R?v���͐��Y,>{����=8+?��?.D�<� �>�$?E�(������^>��5>Cʤ>��>C

>�S��+�߽�?�kT?ô���������>�����}� 9Z=��>mz-��t���]>;��<i�����SК�N�<��U?�0�>�d'����42���g߼?�O=iv?.?㧦>�j?�IB?�I�<R'��+O����>�=�}W?2�f?�[>��5Yʾ~S��ޘ6?=h?��L>�yi����a�-��"���?h�q?HB?��㼥Dy�/���w=
��+1?��v?s^�xs�����K�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�%Þ?��@���?��;<��Q��=�;?l\�>��O��>ƾ�z������'�q=�"�>���}ev����R,�e�8?ݠ�?���>�������;�=��>��˧?D7�?�c��1�/-���~�D��ِڽ7�����Q������9Q�֗־L-*�.޳�dB=��m>��@,T˽v:�>_*o�`�ҿ��˿�Ȝ�e����ƽ��&?o��>�zL�~վ����T9h�s'��=�~�˾eO{>D��=����骾����2;�
��>�>��s��>�6�Ǽ���Ⱦ����>�(�>/��>E������o�?����Oٿ�٣������K?���?8�?�� ?UT�=.Yξ�~ž?�����O? i?�ZR?�]ǻ�¾qP⽜�j?~^���U`�4��IE�U>�"3?D�>7�-��|=#>���>�]>�!/�w�Ŀ�ٶ�2������?V��?�p�A��>���?hs+?�i��7���U����*��*��9A?"2>�����!��/=��ђ�{�
?�}0?[w�7,���_?�a�L�p�+�-�M�ƽܡ>��0�+e\��C����#Xe�����?y����?*^�?H�?>��J #�.6%?��>����?:Ǿ�<#�>^)�>A+N>�F_�,�u><���:�#i	>t��?7~�?�i?ƕ������SV>��}?�#�>��?o�=!a�>d�=񰾈�,��l#>"�=�>���?Y�M?�K�>�W�=��8�v/�_[F��GR�-$�5�C���>n�a?��L?Kb>{��($2�u!��sͽb1��G�MW@�Z�,��߽�(5>
�=>�>T�D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*��п�/��dX������C�=#qm=N5>9⽜��=U͖<�*�}M��S>f�>Z%�>KG�>τE>�oH>ǉG>g ����%�ӏ��i����@�i�wj���r����ǘ�����Ͼ� Ӿ�������ձ��/V�r�'��+�=y�S?k�M?H�?c��>����I>�P��2���=>���>l�.?�^]?ٴ?�q�=UU�`V�IO~��
���[���'�>h��>�?�>��>
��=j�>�o>i*�>��=ud�=r�ͼD�=��:>�2�>�T?�ɻ>�O>G0�<𡾿�w����W�]�������??4���"���������&>
H?':a�{䉿��ؿL~��
F?��u����\��"6>��?��O?AO>7��fў���=�2'���~�{P>��s���Ƚ�Y���=�)>?���=��>kI$��gH��F�M�����>@?�q��sq\�0ts���G��ѳ��+a>A�>	]��a,�I}��B�f�<r�0��(.7?3��>%?(��ѧ��[��㗧�eBk>״�>�r�=Ls=�T�>f!s�P���� ����=�f�=��G>�6?��>ؚ=��>�����r�-R�>��C>fM>�I?�o&?�����B��j������3�>���>�;�>�>��&�u	T=�9�>��> �<uj�<�}���J��>f����tP���<�>[4޼!S�=��=-h9��z� .\�!�~?���,䈿���d���lD?V+?Z �=W�F<��"�= ��yH��@�?n�@m�?��	�բV�H�?�@�?S��8��=}�>�֫>�ξR�L�ٱ?��Ž.Ǣ���	�;)#�YS�?��?��/�Rʋ�*l��6>�^%?�ӾOh�>xx��Z�������u�_�#=T��>�8H?�V����O�j>��v
?�?�^�੤���ȿ6|v����>X�?���?g�m��A���@����>;��?�gY?soi>�g۾A`Z����>һ@?�R?�>�9�}�'���?�޶?կ�?�>� �?�2x?�W�>�<!�1'�貵��l���)���,�9��>�H>q,߾َW�:*�����n�P��t���>��!=��>E��e���B>��Z�I���B���cv`>��O>���>�7?ox?�H
?_U�>{�=��>avr���Ⱦ��K?���?,���2n��N�<[��=(�^��&?�I4?k[�|�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��M��<��K>)4�>�H�>�$���FK>��Ծ�4D�dp�>�ϗ>�����?ھ�,��8S��GB�>�e!?���>�Ү=ۙ ?��#?��j>�(�>CaE��9��X�E����>ע�>�H?�~?��?�Թ��Z3�����桿��[�r;N>��x?V?rʕ>b�������vkE�9BI�6���^��?�tg?wS�0?<2�?�??a�A?~)f>և�(ؾo�����>$�!?gm���A�V3&����:~?<Z?���>�]��^{ֽ�ټ&���2���?_5\?LZ&?�q���`�X�¾�w�< �!�ӊA����;N�C�Λ>o>����
��=�]>�@�=.�m�xh6�h�f<��=i��>���=K7��I��=,?~�G�*ۃ���=�r��wD�s�>JL>.��٬^?<k=���{�j���x���U�� �?��?Qk�?�
��˝h�E$=?��?]	?S"�>�I��v}޾N���Qw�~x�/w�K�>h��>�l�S����ә���F����ŽDx�k�?���>���>��>2�'>!b�>h��������7�yV�Uv��Q'�~@�-��پP�M�p�S<�T�Zb����>�ʽ}��>i?�a�=�-U>�-?=�p=Ȼ�>چ�>Gt�>���>l(�>��>qe�=m\	>�&H���R?�����(���o\��6B?.[d?�I�>�k[�����eV�%�?�F�?bJ�?&�y>�sf�[*��-?�c�>�瀾C�	?��I=�-�j�<�j����r�������>݆ڽ-�:��%L�g�a�*
?C?cHb�>h̾Z�߽�I��B��ۃ?��?����@P�@z���;`�Z�W�3��$�+ԫ�30�RՁ�F�/����Ȁ�L�!��<���08?;��?���O̾�s��h^�PCI�So�>��>��|>� �>��>Ǎ�M���C�T|U�������>��V?��>:�D?2�:?lT?�L? h�>fx�>�
��~��>�����E�>�M�>�;?�Q,?�c+?�?��)?�}]>���W���!׾�U?��?�?,?�n?ebw��ᓽ�{��?�~���j�_������=S��<7/ý>�����\=��K>�v?z��L�8������k>�7?��>y��>B͏�Xh��Vw�<a.�>2�
?�^�>ٓ��:r��M�P��>颂?�E��X=�*>4k�=7���$����=Y����ʐ=v���Y,<���<�b�=ݕ=�)m��i���;O��;٠�<hm�>��?��>�:�>_2��� �������=55Y>GS>�>�Iپsy��/%����g�nny>�y�?nz�?� g=/�=�C�=���fX�����x꽾-��<�?!6#?ZNT?v��?J�=?�f#?O�>��,K���]����9�?s�&?kr>(`)�7E��/��9]�og?�?A����e�A,(�� ��ϱ���o>�F�k���z
��Oh��_}>��`3�==\�?4�?�GF�[�=�ņ��R������z?�>'�>E3�>���R�̃����="?��t?�׳>ouU?&�y?��[?ݦ6>�6�g����+���H'��F >�>?f��?�1�?07w?�Z�>�>9����%����'�t��ڄ��<��=W�h> �>�c�>�ź>���=����)����D�s^�=��>M�>y]�>���>!.|>0$<�/E?��>V����y
�y)���.��?=��+u? �?5�0?L-=q��B��D���S�>m��?�?��-?�<Q� �=S���ݴ������w�>i�>�y�>k:�=�%l=/�>ݿ>h��>�^����6��pW���?��D?���=�ſj�p��!n��횾c�<�Ғ��Rd�Ɋ��8X����=�䙾ø�Vt����W�����Go��궾�)���x���>^�i=Cb >�q�=��<��ǼV��<L�7=w�<��=T�e���<��/�y�λ�ċ���D��}�<�aE= ����˾��}?�3I?^�+?��C?'�y>Ɩ>�Z4�ř�>�����8?xxV>*O��8���e;�������
�ؾ�v׾��c�
ן�=m>�FI�0�>�[3>�U�=���<N�=�v=LJ�=�^��=z��=�J�=�ˬ=U��=|*>N>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�i6>M�>�R�]�1��U\�n_b���Y�ҷ!?:�:��U̾I̅>�=&�޾ehƾ��1=� 6>?�]=�U�a\�ט=UR~���==�j=j�>�'D>%��=Ѱ��ŷ=<BN=�y�=�O>A�:��5���*�U�7=մ�=Q|b>�]%>#h�>J3/?2C8?��s?�s�>�վy�����;��>]�>�a?V>��x>�
?�?MA?�1Y?Z��>[_<�0d�>��>���,�w��Y��v����6c�?L�?���>�^�������W6�%W�N�P�?�55?\�2?�?�>�U����7Y&���.�/�����4��+=�mr��QU�J���Lm�;�㽾�=�p�>���>��>2Ty>�9>��N>�>��>�6�<~p�=�⌻���<� ��x��=�����<�vżT���$u&�:�+�H���l�;��;-�]<͡�;
��=���>	:>L��>ɏ�=���L/>г��-�L�=��=�I��|+B��2d�}H~��/��V6���B>{7X>�p��r3��6�?��Y>�q?>���?�Cu?��>t �޼վ�P��4Be��ES�s�=��>��<�w;��Y`���M�2�Ҿ��>jL�>S�H>]M�<5<���\��u�>��Y��HN��3z>q����������!�E��ݛ�ۡ�����E�ьj?N����;/>�j�?A�5? ��?��?~�q�˖����>��ؾ�����vھ,�[�}�6���=?'�*?�?�[C���V�ɵ���ݽ�K�>�>�\�K�k���HH�`��=�þ�m�>�����þ4�5�����v�� mQ��)��>"%A?��?��A�SU��R�T�j��!���?�\u?��>�?���>ߔs���CVL���>�)Y?n��?j��?�D�=7�>�Fm��>Hk?7�?C��?�g?��+��>�EM=��>�҃�lB>&��=�|�=��1>.?]B?��?�\��������n��W�����A7�=Rϑ>Kۆ>y�j>��D>���<<)�j	>�ߤ>YF>'��>Z\�>�E�>�ݾ�=�V�?Ԝ���=`�?G?8>�4>>���Kl>=k��������,<�ƒ��;��˭A�BG����ʼ.L�<��>�˿VK�?�	�>��*�=�?A��,�/�GQ>T�g>��2w�>�k=>ۡI>�?`>��\>+�R>��J>tWZ>ebҾ�">�r���!��C��R�z�Ѿ��{>���3/$�(	�[*��NoL�Ws��t���/j�nV����=��g�<^�?�~��c�j��w)��!���? ��>|�5?:��Y�����>,��>�m�>��������/��F��Y��?+�?1;c>;�>U�W?+�?֓1��3�vZ�m�u�e(A�,e�m�`��፿���1�
��
����_?��x?�xA?T�<�9z>m��?��%�ӏ�J*�>�/�[';��6<=�*�>Q)���`���Ӿ��þ�8�GF>J�o?Z%�?CY?lUV��3�%*>X�:?'�R?Yd�?oZC?��)?�'H���?/55>��>�-?��W?LW"?C��>� ~>V
>�%<���6;��2�)�.�i5�(���x=b==�=]�=:+v>Z>=jt�{G���{�<�����=c�;�|<>_o>��>�y`?r��>��R>Mb4?�����H�WZ?nq�>�;@��Ѯ�߳���@���>�If?;B�?p?�Յ>Id>�&���di=[��=��w=��>�K�>��"�Q]����\<�[�=D�>'�=Dp�	b�$�������<?��x>��>�/|>#
����'>B}��u0z�٤d>[�Q�O̺���S���G���1��v��X�>��K?Q�?ژ�=K_��)��If��0)?�]<?OM?��?:�=�۾>�9��J��=���>]�<�������$����:�6v�:8�s>�2��iJ���9>qN.�ϳ3�K���}4O�"��ǳ<�~H�vm>�cվo�*�4j �<�ؼ����u���4.�����]�I?��=�������ެ�^W�=O��>�5'=��Ͻ6{� �B�N^�j1e=c��>�㔾,Mu=��̾�a�&�ξ�+u>U?�.Q?L��?^OQ���y��M�����)Ⱦ)�^�?�H�>�/�>p�p>��=c[ž!����X�ɇG���>�&�>dq�>pM��8p�م�ۗ�[v�>���>
�=�?��W?�u?l?u?��A?��?��Y>�̽��߾�9&?O��?#�=��Խ*�T�}�8�'F��><x)?.�B��՗>��?�?��&?r�Q?�?0�><� �;@�ȋ�>�G�>\�W�:\����_>x�J?ׇ�>a-Y?�Ճ?9>>_q5�fϢ����u\�=�>��2?�(#?C�?'��>q6?m�#��͑��?�Ȉ?�AC?�).���,?>��=�2F<��{>�d�>W�>`�7?��w?�=�?d�i?��
?d>1�+�1�.��zӽ�<:����=���^I>[�f��5�Z@��n<�=Ej/��rp�h�=��/=>��=v��<_W�>�s>���z�0>��ľ	K����@>�S��IF���Ί�(k:�� �=Ռ�>�?���>uK#�2В=4��>wJ�>����0(?��?P?�;��b��	۾*�K�Z�>B?w��=O�l��~��w�u���g=��m?�^?L�W�g����b?�]?we��=�c�þ�b����^�O?[�
?O�G���>x�~?��q?���>h�e��8n�	��Cb�G�j�#Ͷ=�o�>FW�'�d�!@�>�7?IQ�>7�b>23�=pu۾��w�l��?���?c�?	��?#*>��n�L3�DK������ ^?\�>[�w�R�?�d��������4��l�������[��(����¾��;��Wa��Ž��
=�?���?�?�̏?�r���e��fO�nr|�Q�y�S'�Yr��@��R��$�	�7�"�+��=��о��_��QҾr�D��y�?@2?-�ݼ���>0-־�R�j�V�=O���i�`��&'�J�ٽ#��=U1Լ��������߾��(?u�>2�>M�S?�_X��I��38�N������J�>J��>6?�>�{N>�=Z=��}�����v��H��J�<��q>?Ff?�G?Prm?���}4����M��1���C���O>v�>�o�>�3��d���$�u�@�_p���������^�k=�)?��>n@�>�h�?�?�� �AH���Kn�hF'����<���>Fm?y �>B�v>��н2,!��_�>��m?�`�>���>�%���� ��{��нZ��>l��>gD?It>sE'��6[�Û��K��>=8�L�=�/i?����I�\���>L�P?��T�rqa<;��>��������G���+�ݮ>3�?f��=k,:>�|ľ#9�^ |�s����j?�3�>�����p�+�>��a?w�?{� ?֒�?3$G=���̙>�Y'?̹?�>?�Fb?�c?˥O>��'>���������X;�xk>��>J�=Y�9>�I���1�V]½*�˽P���N��ν���=��Ž�-����:��=޽ۿ�K�,�־`����m�	��Ȋ��ٹ�TP�����;��ܹ��a�y�lp��U$�R�V���d�k��Xno��?x��?������Mՙ�ꦀ��< ��>�az� yr�~:��"���^���}߾j쩾+#��5Q�~2j�84f�N�'?�����ǿ񰡿�:ܾ4! ?�A ?8�y?��7�"���8�� >)C�<x-����뾬����οC�����^?���>��/��l��>ू>�X>�Hq>����螾v1�<��?9�-?��>��r�/�ɿ`����¤<���?/�@E�A?`)���vN=�r�> �	?�:?>�0�J��`�����>e5�?��?�N=�YW���ye?�#<uF���ǻ�V�=��=�=,I�v�J>=o�>Y���@��ݽ�-4>#C�>AW"�s���_����<��\>hoؽS���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��=�����ȿ�1�p��#��=��w<d���x/�q�)m���]ʾ/����]�Fi�<���=PST>,i�>�H>�B>��T?��n?9P�>�y>]=P�d���!�W������}7��4j�;&'����%*��]�־sQ�}�(�����<ҾU=�	��== R�Fx�� � �C�b� �F��.?o�#>-�ʾ
�M�ƫ%<��ʾ�䪾ƅ������%̾�1��;n�ϟ?�A?-����V�J.�^��-���kuW?���[��U���=x@����=GR�>"!�=(S�\3���S��g/?U�?5���M��è->ި �O�=/�+?F_?���<P��>)�%?��#��|��Y>�5>[��>��>�>R歾�kֽIQ?L�R?���wI��L��>������q���=7>�2�DP伟�X>��h<Z����|�7���j0�<��W?`S�>�*�6����������)6=
x?��?�.�>��j?"+C?\(�<�1���R�c�	�ʚ�=20X?ci?p
> ��W�оK,��#^5?�	e?E�N>�hd�H��%~.������?��m?��?�V���k|��ϒ�.U��5?��v?s^�{s�����8�V��=�>\�>���>��9��k�>�>?�#��G������mY4�&Þ?��@~��?��;< ����=�;?f\�>ЫO��>ƾ�z������"�q=�"�>���zev����R,�c�8?ՠ�?���>������As�=ĤS���?�S�?���mѼ�A�ʪp�ض��\��#��=$ϐ�?R��Ѿ��:��ξ�����������t>u�@a	����>���	ܿ����^���Mm�������>�y�>Rӽ_;��	�R��oy�~T���G�ٯ�����>X�>��F���KDy���8��B=�&�>y�N��܁>�ms����󰥾z�x�6�>��>��a>q߽����P�?/����ο%a��#�価�m?�;�?]��?23(?	�5����W�/�L�=/a8?�3t?��a?��G����ǽ!�j?�_��xU`���4�rHE��U>�"3?�B�>R�-�S�|=�>���>g>�#/�x�Ŀ�ٶ�=���Y��?��?�o���>r��?ss+?�i�8���[����*���+��<A?�2>���E�!�>0=�RҒ�¼
?W~0?{�e.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>�(�?4��=�>�M�=�ڰ��.��">���=�]8���?�M?&o�>��=��8�9�.�@F���Q�����C����>��a?yVL?èa>N[��/��!���̽�(2�d�켡R@�1�*�|
߽`5>۸=>v�>%�E�BӾ��?kH���ؿqc��Nf&�dA4?���>D?A���`u�2��SP_?�M�>8����~���k�%p�?��?��?��׾��ͼ2�>v�>�{�>r�׽j��,+����7>��B?�Q�L�_o���>�	�?�@�Ѯ?��h�	?(�Q��#a~���]�6����='�7?�-��z>���>X(�=�lv������s�㵶>4@�?%y�?A��>A�l?�o���B���1=TQ�>�k?�o?{�m�)���B>�?5��Y����H��f?��
@�t@%�^?����ؿ�3��kș��-վl��=�~�=�*O> �^��-�=	�=�Ss�(�y����=9�]>�ō>�G�>iPz>���>�>7|����(�۴��t����<��6�Y��T�����Z��_B*��(�;���ָ�Y����i���똽x��-�(��C�=��`?{XE?��c?Of
?��F�(�>�f���m";�}��y6
>'��>�1?�?J�:?�o=	�����S�I�}�u<��>l��߆�>`�B>>��>K��>y+�>�,�=-��>%��>��+>�Q�=�=�{�= ��=���>(��>���>;1�>�B<>ʑ>6ϴ��1���h�0
w�y̽6�?h���K�J��1��{9��妷��c�=�a.?{>����>п:���[2H?{����)�	�+�!�>��0?�cW?�>S��5�T��:>}��Ӥj�/`>�+ ��|l��)�['Q>�k?�f>a�t>��3�&,8�2�P�Dq��{|>�36?"��q�8���u���H��xݾ�L>Mǽ>�M�N��얿b�~��9i���y=E�:?�p?jC���U��މv��~���DR>��\>��=��=:�M>+�]��,ǽr�G���.=���=��_>���>U�>��>t��>��~�M�4��>l
>��>��e?��C?��G=���;"ヾ�����>��>��>�r>N�;� `�=u��>w�C>�Ž��`���)F���8�>������k�TqY�G�e=����=(��=�.��Pz�q[F��~?���(䈿��e���lD?S+?_ �='�F<��"�E ���H��G�?r�@m�?��	�ߢV�@�?�@�?��K��=}�>׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�<l�6>�^%?��Ӿ���>��@����G��V�d���`=��>3�P?�*�Y��������?���>���C���!\ÿ��u��l�>k��?N�?�/n���OI�_�?�!�?W�U?�|�>-�������L�>�@\?d�]?n�>N��j� �ۼ?�y�?2Zg?�$>���?�"x?�?�XJ��9�x�������f@K�W���F>�/j=����G'��Y��]��4�q����V)>�e0=:��>�R�rf��X��='	'��s¾qr*��=>�;�=�r>)��>%�>S�>��>�U���ͼլ��\0��i�K?���?���2n�Q�<��=7�^��&?aI4?yw[�5�Ͼ�ը>Ѻ\?}?�[?�c�>]��C>��B迿1~�����<��K>4�>�H�>0$��?GK>��Ծ�3D�wp�>�ϗ>>����?ھ,��QB��uB�>�e!?���>Ӯ=�� ?\�#?��j>�7�>�~E��C���E����>�I�><P?��~?��?����Vc3�����꡿/�[���M>zy?|7?���><|��>����=�AF�������?��g?y@��?O:�?��??!RA?_�f>�a�d�׾W6�� �>!�!?���9�A��&�����?YR?���>3�����ֽ��ڼ������T�?�\?%b&?�R���`���¾��<>���m�G�;7�>�_ >:>/���F��=	�>6�=�,m�m6��fb<vP�=���>��=i�7�^Z��/=,?ϿG�|ۃ���=��r�>xD���>�IL>����^?`l=��{�����x��	U�� �?���?Zk�?[��?�h��$=?�?T	?l"�>�J���}޾9�྾Pw�~x��w�V�>���>%�l���J���ڙ���F��\�Ž�,��^�>^��>\��>��?�g> >�>��`�7���,��E���L��Y�QI�?j/�(������� �9e	�"žl���I��>n
��K?�> 3?J8>c��>���>-�����>��>�Ҝ>�Į>�Y>���>Ø:>T}�=����RR?:���@�'����G����8B?<kd?w4�>D~h�^������}�?g��?�n�?�Dv>�kh��+��r?�B�>Y��p
?�9=�*�0��<@I��)��M������K��>�f׽:��M�sf�Mb
?0?5�����̾R=׽�R�/�<哆?�5??>���>W��;��y�.�i*f�'PX��/��Hľ�pJ��4\��ig�i=��5���B[@�bc��aB?f�?-���ᾕJ+�	Gg��J!����>8��>���>�e�>z�%>�I4���'�yyc�c<�iǽ��>3O?Oc�>�sL?vY=??]M?�J?�V�>x�>����m�>g��<&�>�z�>9:?#�,?u/?h?x�(?(�h>^�߽����B3׾B�?��?I�?b�?K?����tK����f*��Kx�4^�.=��<dҽ(i��3)=�?I>��?)Y�k�8����sk>��7?���>5��>�,��kl�����<u��>��
?߯�>5P��c�q�������>���?����=!�)>k�=4>��E~��Y�=/���=��=uo|�V�<�q$<iT�=UЕ=�n�	So8x;�b;��<Do�>r�?n��><�>7"���� ������=�?Y>y�S>v�>�(پ
p������g�ny>t�?Dz�?Mh=��=���=p���S�����v�[�<܃?�U#?�eT?���?��=?]#?r>1��F��;]������?�z?�\�>z2��uP��l����U�D�>��>�q~�`����C��'�:����>�m� C��N骿E8v��J8�О����;4Q�?�y�?,�3��UK��&���R���u�,7?��>Dm�>�4?(�'��|M�= 
�T`�=�|�>2��?�޸>��S?bLw?b�X?(V>�:��������z�^��>#�A?/g�?]q�?�.z?3��>�s>�5@�+ܾ�m��m�.��C��rx��=�'Z>LD�>��>�P�>��=�wֽ]ⶽ�w*�]Я=��> ��>�ԭ>?�>�e>l��;_�G?ڵ�>so��4u����qӓ@�qu?s��?�,?��$=�Q��VD��&���_�>H+�?��?��*?�{N�<��=�R̼����<s�-��>��>�&�>�3�=GTU=I!>��>;�>D>�m��I�8�23K��	?��E?��=�Y����s�pe�.���U@û>��XPa�.Ǐ�/�G�<M�=RK��ߝ�����LO��ӧ�b����Q��Jf���u���>�]I=n�>`�>��<�{��<F�ֹKd�;�=k�x����l�=����fL��I<��_=DP���ʾc�}?6cI?8+?,qC?	y>��>�Q8�˗>�w��?��V> �J�>��V;�5���L�׾�?־G�c�V���N	>��I��>��3>���=�ׂ<�5�=�kj=�=�c���=���=��=F�=M;�=�I>�d>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>}�>�Z�=��U�a3���?���C��%��;*?34���Ͼ���>9^>&gվ�޾Y��<�.>(�N=u�a�U��C|=�����bf=$�w=Oȅ>�<>�=@ڮ�>�=�e�=6>b�c>�=�ࡻ[g�U�=.>��r>ŭ>Ұ�>(?>|1??M?F�>F�l��,��>�;�_j�>P�]>���>�B�=��>a��>%�7?��A?�eK?+"�>Ԅ$>Fi�>�Z�>z�"���]�[
����'9���_?��?Gz?۳�=|���O���V�XT���?K?b?��>�P�4��xP&���.�1�����ն��*=kjr���T����Z3�j��d�=�p�>���>�ڟ>�jy>��9>e�N>��>5�>qy�<D߅=8R���`�<ɷ���'�=�����<��ü�0����1���*�eV��@�;�?�;`^<���; ��=V��>0P>���>"��=7	���>/>���>�L����=�G��A+B�(2d�6E~�/�i]6� �B>�5X>�x��-2����?��Y>+y?>K��?�9u?8�>�(�b�վ~R���Ze�RWS�&Ǹ=Ү>.�<��|;�\`���M��{Ҿ� �>K<�>[N�>+~�>�"K���Z�~�==�ξ-C�=F�>@.���!7������F��q��O���t���2���Y?	�����$=�Y?�?���?f�.?��j>$��ݝ�>cHؾD.J����g	=�,��,HD?�H(?�C�> a.�jd;�ā;�����>WC�	�P�Y�����1��k������>�d��G�Ѿ��4�o7�����;�C�Mu��>u�L?:�?f_��Q���RO�z��c��
�?�f?ݝ>��?�	?�n��K�ﾍq����=��l?���?�y�?��>k�=A�o�;��> ��>8��?�!�?��w?�E��!�> �p;;�2>g"���>�=�@�=�`�=`�	?(`	?�c?����a�����1�f�O�e�=A�<�Տ>�9�>gp�>�>�E�=���=��C>��>Ț�>}�>�O�>�`�>8���x��j��>����^>y�?�"o>��>���<�[ϼ¢�<6�+�������T���h�Õl=��a=^9�����>B��$N�?��>Q��>����/��mQ>-�>�I�=��:>��,>��?oH�>�X>���>�c>.9�=�(Ӿ@�>S��%!�U]C�F�R���Ѿm�y>����^%�pe�̱��mJ��]�����#j�F0���l=���<r.�?i��sk���)������`?q��>96?����`��
�>-�>��>)���v��ṍ�{7��?���?�;c>��>Q�W?,�?Ӓ1�O3��uZ�1�u�j(A�*e�Q�`��፿
����
�����_?��x?%yA?�R�< :z>T��?��%�Fӏ��)�>�/�$';��?<=Q+�>>*��U�`�{�Ӿ~�þ�7��HF>w�o?1%�?fY?LTV�-dH�{*�>�J?/�(?{\�?p�?HNK?Q��h�?�ɉ>C�?J^?�	9?`PG?��?M�A>�>��=�<��#�;ߚ����$E����� �=#%=�5=��ԼFK=���=�ď�bǴ=ǽŽ�b'<l��=��q>Y�~>�D>�u�>,{j?���><~h>�5?ջ'��J7�>$��( @?<��>J4���p+���R�8��2��=#Cb?I��?�Cc?��>�.�'4뽗�3>Lo]>ݐ�=��Y>&�>�V���f�ݨ>c�=g[2>�gd=�载jl���g���᩾�/8�C>���>	0|>Y����'>�|���0z�C�d>L�Q�x̺���S�j�G���1�؄v��Y�>�K?��?֝�=;_龻,��[If�I0)?�]<?�NM?��?9�=��۾��9���J��>���>�U�<��������#����:�y�:}�s>�1���ՠ��[b>���n޾{�n�J������L=�z�ʦV=��`�վ�$����=�*
>ܱ��/� �O���Ԫ��0J?�rj=zz���LU��`��Q�>�Ø>�ۮ>S6;��1w���@�Ը��;�=���>�;>����m��ʁG�~9�z�>��U?tlX?�r?��i�ŮS��;�Qp���a��Po�?�@�>!��>mU9>ٰ=뀝�����"�e���7�%p�>x��>�����?�����H� ^�qP�=�Q?X*E>��? q?��?��d?{6?�V?��8>���bs���&?�i�?�H�=k[ֽ��U�5�8�׮E��a�>��)?�G>�+J�>u??�?�a'?�Q?a?F>ū����?��u�>���>+X�����Ha>K?G��>2-X?�3�?� =>\85��-�� Y��N�=,r">;�3?��#?��?���>���>O瞾�I>k�|>�c?�?_�\?0��;�w�>?D߻nq�>�S�>���>z}�>��
?p�R?.c?_�d?�Ժ>�[V<��������2�8�>"(���<��b��z��;�<�r�c�p����<���1x,=�����>�V�'=C�(=��<�L�>g}r>|¤�L8>|Է�Q7s���T>��-����D����C0���=)V>ґ?�A�>d�	��r�=x#�>�W�>==��'?��>��?_2=�o_�3?̾�-�-�>�o2?x)�=MO{��=���Zx�H�>=��h?s�\?�=q����2nZ?=QZ?5���7�saɾ�S���ݾ��4?�#?wV��u�>ш?əo?�1?|�I�7�]�$��]�D�4{a�˳>`�>��A]D��I�>#HD?��>%>G��<�Ҿ#l�����J��>b��?aF�?v��?�Nt>L\i���ۿuw��p���	T?��>�������>9?��I���F�ƾ��վ�־�׿��d�����Ⴞ�%0��`�`d��d��<�� ?��p?gVy?�Q�?͇�UG���q�\[��;���M��侜C��Y���F�_�s�3uK������Ⱦɍ�с��.>��p�?u,?��-�w��>�뤾�@�0�ھx�>4ٜ��<$���f=15���*E=��=dm��B7����U{!?;��>X��>�??�J]��=C�Gk5�+5�����2>C��>�i�>wB�>?�+�6{<����4־ @�����gfv>ۍc?c�K?��n?�P�n1��}��B�!���-� i����B>�>��>�W��-��&��7>��s�C��-u���	��}=a�2?m3�>ʛ�>?F�?��?@k	��G���x�bO1�~L�<&e�>�i?�\�>���>�[н�� �E��>��l?&��>��>F���sX!���{���ʽm&�>�ܭ>��>Y�o>3�,�o"\��i��\����9�Yg�=;�h?������`���>�R?R��:ƛG</y�>a�v�?�!�k��¼'���>}?瞪=Ӣ;>`{ž]&�ߦ{��6���U)?/�?@֘�ZJ�儁>�.&?��>�h�>��?���>�@���=lB?�&g?F?��>?
N�>�&�<}Y׽{F��^�.�rf�<װ�>��>��=�p>�
��兾R�B��/:���;8"��@�ӽ��<�V!<f�=�����>��ڿfK��־y&�X���
��2���w������`�#s������y��a�"3�FtT�\5_��I��D�l�O��?f��?ɜ���Ӂ�������� �>��>�܀��1��pΨ�����6��(��R��s�$�0YP��ui���f�5�(?�U���ƿ�ҡ�
�߾��?q)?g}?-��`���&0�9%>�Gb<&�a��I����|�Ͽ{�~b?� �>��o���^_�>��}>_-Y>1�w>a���������Z<eo?r+?G� ?��c��ɿh���\�<�o�?
4@��@?"u�a����W=���>$�?+!@>Gd���sʈ��P�>��?�0�?O>��F��@���a?�r<��A�?��<͈�=^+4=pt�=y�q��y>>�>���P؆�������=�";>�С��0��7����=gw>K0�i�ݽ�Ԅ?�x\�=f�q�/��S���V>9�T?-)�>44�=��,?�6H�.}Ͽj�\��*a?�/�?0��?q�(?�ݿ�՚>��ܾ��M?�C6?���>@c&���t�[��=h������*'V�3��=���>�z>��,�#���O�N�����=���Ϛƿ�$��/�,� =�C�0�\���潲c��o!\�,4��p�L��P�d=���=ܝQ>��>ҚW>��Y>�XW?��k?��>�>d������ξ��n���7���ڊ�~ ��y����#/��0
�~��,��Y�ʾ =��3�=�3R����$� �x�b�V�F���.?�$>��ʾܲM��~1<�[ʾ4��� ����5'̾�1��n�w̟?B�A?������V�������X�����W?]O�����٬����=����m_=�B�>$)�=���:3���S�zm0?�r?��������*>*��N=� +?��?gRf<-�>dh%?��)� �޽��[>@4>�*�>o�>P�>�]���p۽�i?-T? ��7��g�>z��{�N�\=7�>
�5���yZ>���<�ዾ�PK��;��@�<��Y?�Av>�+��#�䚣��놽�=�x�?��>� �>\�~?};?�>�)ྮgS�n����$��f?��w?��>�逽v�Bʾ#�)?mv_?��m>�S_��'ݾ��,��j���?3|t?��#?�[��R���:����Ӿj�7?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������[G�=m����T�?~&�?[s��[eV<*���k�� �Rܓ<-ͫ=���i=%�I
���7��Ǿ��
������Ƽ���>�>@�i�;��>o	9��=�;SϿ9�ڨо�+q�W�?�N�>I�˽Cͣ���j���u���G���H��,����>��>�ȹ�����T8z���9��
�:j�>�hC<�ǧ> s�'V��2���5=�_�>�w�>!/>��[��w���F�?�e��ο+���M���W?D��?��w?�<?�+=M�Q�L�H�dÖ��L?�'|?��e?��<�|J�������v?�-��1O]��X��}r�����?�?�#?�uN����>�`[>�a>���Ȳ��ʿ��˿`�0��?]��?=1Ӿyj?���?�?��<�ó��s�&`d�C��<,�?�]�����¾z�_��	����>�(?�p��i`
�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�)�>�?d��=�r�>���=)ٰ�m�1��d#>��=8N?��?��M?�E�>O�=�8�g/��LF��3R�D*�y�C�	�>N�a?�kL?�6b>*6����3�6� ��ͽ� 1�B�缙G@���,�~�߽p;5>��=>"J>��D�'�Ҿ��?H[�h�ؿ4g��f�'�� 4?.��>g�?(���&t����%J_?���>��^"��p��3@� ��?s9�?}�?�׾bм�=>Iح>�Q�>�ս����eu��U8>2�B?���k=����o�AQ�>�?��@(ͮ?�i�	?���M���_~�;��
7����=n�7?\�{>��>]��=�^v�±����s����>�;�?@x�?5��>4�l?&xo��B��f2={B�>��k?.m?�<y�J��	�B>�?������
:��*f?t�
@tt@b�^? 𢿳п�A���I���_ݾ>��=��;=��m>�Eڼ-~�=�X߼��(�%��*�=�a�>�W�>�y�>$�>]s;>�[D>�/��_G$�]Ң����S���7�8Y�\OF�+"��>\��Y�������پ��ɽ:Ľ@ʊ�i�����#��Y���*>.(d?g=?��k?$?�I=i�*>v�����=��b��]�;�`�>�(3?�{X?%2?V#>�Y���=[�a�������𐫾���>e�U>��>��>�ie>�t>�EG>U=>>'|2>�T~���<�����<"M�=�w>��?�>�C<>��>Fϴ��1��k�h��
w�r̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)���+���>}�0?�cW?�>!��t�T�4:>9����j�5`>�+ �~l���)��%Q>wl?1�h>,�y>f3���6�_oO�7����~{>bs5?읶�f�;�®u��iI��޾	L>X�>�+A�:��ɖ�O�~���h��e�=�;?v�?�ʸ��毾̶x��I��@V>mZ>�=�F�=^O>�g��Ž�VI��"=y�=�!`>�v?�Q>�Tz={ɧ>�����5����>��+>z->�K7?��?�f��Т��`o�o� ��4r>l��>��i>���=�4=�;S�=���>�GS>��#�I�C�)D�[q\�~�d>Ը��2V���:��(�=���Co>ၧ=��ǶD��y2=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ� �>��1�屘�pE��K1z�r9Ǽ�x�>E�a?ȏ����=�W9<R�>p��>{R�����ʿڹ���-�>���?�v�?��Z�ȍ��Rc��g�>Ɂ�?v�e?��>�4Ҿ��M��m�>��:?��c?$��>�U��������>[��?��?*`K>-ޑ?p2s?��>n�t���-����ʽ��h�=M�����>�+>֊���E��ʒ�p����h�����|_>Ջ=pL�>���ʧ��uX�=�����4���'��A��>�s>�%O>��>ƕ?A��>�N�>�/=v����/��������K?g��?����m����<O-�=��\���?'4?y�Z���ξ�3�>u\?n��?`�Z?��>� �`6������s��<�YJ>^�>v�>����vL> �ҾBF�?L�>�W�>�¼�+ھYm��A��R�><� ?��>�Ԫ=2?�{?���=|�>D�K��Q����D�k��>m��>�}=?p��?�J ?��ʾ��'�^)���2���bb���=3�v?��#?}*�>g1�� G���sؼ!� =:��^eh?T�b?��)>��@?Z�?�4?��]?�Q�>=�du��t):>li�>�"?�J���B�~$�]�
��	?/�?�J�>�?���̽gAǼԅ�AZ��.�?�0[?�M&?+���a�ľ�G�<�gĻ��HX_<�0��v�>5�>s�\�=Ԏ>y�=�ѿD��fZ;��=J��>���=��?��b��2=,?K�E��݃��=��r�VqD���>QHL>l����^?+}=���{�=���u��iU���?���?�e�?�$����h��*=?u�?�?��>@E����޾V��$7w���x��t�F�>3��>�@m�P	����
���*C����Ž,h��/�?5�>��?��>�r]>t`�>�U���w�o����Z�;e���2�yi/�eH�~��*I<���l����l�E��:�>:-彁��>�6?,�>}�U>5 ?���<Bͪ>i�>/�>K��>��>.�F>��=���< Cɽ�3R?�`���4(�iI�c����KB?%d?L��>b��p�����U ?O8�?e��?wMw>��f��)��h?�'�>�v}�{\	?�Q1=$)��TǺ<1���~9�>���o-,����>��L�;�d�M���g���	?,�?Rr���ξ[]ܽ!����5ƽ�,v?�5y?�9��7��®��T��뀿\"I�ug����p��?�����0 ��-*~�8��?|��Y?�?^?�1�𳷾n����e�]/8���s>���>�n.?O	�>�y�=��H���-��wg���$�������v>�~k?S��>'�_?J
U?�>?�Z?��>>�&��:0?�������>*��>7k?�V4?~7'?V�?�1)?-<,>c��Kɾe��G� ?G�>���>3K�>���>�K��n����o��dJ�A���F��=�\�<"Ы�������.�H>�X?%���}8�����̷k>R�7?e�>t�>�я�ȋ����<��>��
?�ߎ>H����r���M��>H��?��S�<�S*>:��=�Є��uغ+��=�����=#و��{>�Ά<BV�=�Ŗ= 4�����7\;�n�;�<N��>�?ꇊ>;m�>��� �.����=>�X>�yR>=|>gپZu��R��A�g��3y>|�?8P�?�e=���=,��=�ٟ��n�����Vؽ�Q��<�`?Fh#?�7T?E��?�>?�y#?P�>G�7���b������ĭ?�$,?���>�����ʾ}���N�3�-�?�[?@a�����9)���¾�ս��>�d/��7~�����	D���~�����>��Ι�?���?|A���6��i辺Ø��W���C?���>�O�>�!�>5�)�J�g�;�'.;>�o�>6R?�u�>�<e?)(i?IJ?�cI>cW�l���iϬ�Rq�=?��=�2?t �?��?�Z�?�
�>��[>�m彈��������1>��ʞ�=�=耔>b-�>MR?�y�>�6=�����e��>��`=:>"�>�a�>���>�,�>��T>Ö��R�G?���>;U��T���ݤ������=���u?K��?m�+?�"=�~�:�E�S7���F�>�j�? ��?W,*?-�S����=�xռmͶ�N�q��>�۹>�!�>q�=�F=[U>��>ī�>G$�\Z�i8�dM���?�F?��=�*ƿ,�q��4s��Ϙ��nT<�Y���d�����
CZ�c�=g����K��q��B:\�����F���ڊ��ib���{��j�>޺�=��=�=�>�<�GƼ3�<�J=���<��=PBo���m<��5�n�ܻ䍈�h� ���j<;WI=E~��YOþ2~?�
N?$�*?�!F?�~>ě�=�4�B��>+v�a$?цT>G8-�ø�/'$����d΋��־�ھ+~d��㢾һ>}A{���
>�7>#>	��<�l�=LF�=�(~=��L�+�=�)�=+}�=��=��>�k>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>ٽ7>=>k�R��1�\�H�b�rZ���!?6A;�FB̾K3�>=�=�$߾	�ƾ�.=��6>��b=�m��R\�U�=|�z�@%<=$l=i։>2�C>�g�=bS����=�cI=���=��O>�����7�,�+�K�3=)��=��b>0&>.��><�?�M0?uBd?��>�j��о����r
�>S��=�:�>�N�=�aC>*�>�7?�;D?��J?�	�>X=q�>�=�>\�)���l�E�㾣L��tsZ<��?(y�?c��>y+w<
�A��z��O>�����f�?n�1?�?��>=A���ҿi�g��Z�O�=�u��g=Va��P=� ��O�YS\�)��=_d<!��>3��>�V�>�r=ݝ>�P�>Oc<������=���<�:>O =-B=&	G���������=�޺=*hd��($�S�(�/V�=��}=��ź� �=!��>�'>P��>��=:���"C/>ٲ��=�L�1��=HR���4B��3d��@~�l�.��L6�%�B>KX>~���c/����?,Z>�\?>�{�?m9u?��>}/�n�վ�M���=e��#S��޸=<�>e�<�Pz;�V`���M�UkҾZ��>�G�>� �>���=��_��Z�%Ē>����T�4�>)-���s���i9�'��B̿�w���q��s�'�a�?���>E.p?��)?��?FA"?��>�餾���>�ִ���==�6���B�=�����S?�'A?��>������5��˾�!���׷>��I�G�O�"���Rc0����ⶾ! �> $���9о�2�o2��O�����B�ҕs�&f�>0�O?���?m@b�%m���%O�d��!-��Ǐ?g?=��>)?{.?=����\��}����=o?��?��?�)	>���=���\�>"p?���?ݺ�?�Xs?��A��L�>�:�1!>o�����=�X>��=<��=� ?�L?ԃ	?������	���ﾝg�1�\��=�̭=�Q�>���>�)r>2�=@�=�S�=��X>�h�>9�>޾g>��>�f�>�ǥ����n�&?��=�č>�%2?�*�>~W=BӨ��J�<15L��?�(+�^���W���C�<˰Y��BM=�"μB��>�2ǿ�%�?��R>�����?ߘ����6�TdU>q�U>ܽ���>�/F>��}>^ݮ>�g�>.)> �>��'>#��,��=���6d� �L�\�>���>���D�ý}q쾾�!�H����ɾ[	�M�k��e���F�[��<�m�?�ս"�s�!?;�X-����?F{�>�;?���!�<!�9>�3�>y��>��c�������>��	W�?8�?��d>�ޠ>�V?��?�'/���0��Y��t���@�H�d�O�`�X/��j����*
����_?(jy?�@?~K<�y>���?ʸ#�v������>�d.��d;��`4=|$�>\����`��о%u¾�Z�.mE>�n?���?� ?N�S�9�=�Z>F7c?�L?Lt?l5L?�91?뺽<7?b�5=%{ >��>Q0??�	?�j�>�l>g��<9 ����Ⱦ�ཝ��Ms�D#=k玻�$���������¼�m��|ս+��|<�U�=՞
�s��=�>6�>h�`?&�?{�>I9?m���`6�����I�1?��9=�u�B#_�z��%�վ�_>G.g?��?>RS?��=>^�1�mY��>4v�>HM(>j�g>)�>��3��B���=��#>/�/>�4�=�Ե�L�}� ��iĂ��ϻb�>Xs?�M�>��p�J�>� ��Q��.�>*D@� |����b���>���Y���L�>oQ2?/�?X�>&��H�J��UE�c?�,H?;|9?g�U?G��;V�m��Se/�l����>m�,�+��j�����U�?��E�=��K>�/y�iJ���9>qN.�ϳ3�K���}4O�"��ǳ<�~H�vm>�cվo�*�4j �<�ؼ����u���4.�����]�I?��=�������ެ�^W�=O��>�5'=��Ͻ6{� �B�N^�j1e=c��>�㔾,Mu=��̾�a�&�ξ�+u>U?�.Q?L��?^OQ���y��M�����)Ⱦ)�^�?�H�>�/�>p�p>��=c[ž!����X�ɇG���>�&�>dq�>pM��8p�م�ۗ�[v�>���>
�=�?��W?�u?l?u?��A?��?��Y>�̽��߾�9&?O��?#�=��Խ*�T�}�8�'F��><x)?.�B��՗>��?�?��&?r�Q?�?0�><� �;@�ȋ�>�G�>\�W�:\����_>x�J?ׇ�>a-Y?�Ճ?9>>_q5�fϢ����u\�=�>��2?�(#?C�?'��>q6?m�#��͑��?�Ȉ?�AC?�).���,?>��=�2F<��{>�d�>W�>`�7?��w?�=�?d�i?��
?d>1�+�1�.��zӽ�<:����=���^I>[�f��5�Z@��n<�=Ej/��rp�h�=��/=>��=v��<_W�>�s>���z�0>��ľ	K����@>�S��IF���Ί�(k:�� �=Ռ�>�?���>uK#�2В=4��>wJ�>����0(?��?P?�;��b��	۾*�K�Z�>B?w��=O�l��~��w�u���g=��m?�^?L�W�g����b?�]?we��=�c�þ�b����^�O?[�
?O�G���>x�~?��q?���>h�e��8n�	��Cb�G�j�#Ͷ=�o�>FW�'�d�!@�>�7?IQ�>7�b>23�=pu۾��w�l��?���?c�?	��?#*>��n�L3�DK������ ^?\�>[�w�R�?�d��������4��l�������[��(����¾��;��Wa��Ž��
=�?���?�?�̏?�r���e��fO�nr|�Q�y�S'�Yr��@��R��$�	�7�"�+��=��о��_��QҾr�D��y�?@2?-�ݼ���>0-־�R�j�V�=O���i�`��&'�J�ٽ#��=U1Լ��������߾��(?u�>2�>M�S?�_X��I��38�N������J�>J��>6?�>�{N>�=Z=��}�����v��H��J�<��q>?Ff?�G?Prm?���}4����M��1���C���O>v�>�o�>�3��d���$�u�@�_p���������^�k=�)?��>n@�>�h�?�?�� �AH���Kn�hF'����<���>Fm?y �>B�v>��н2,!��_�>��m?�`�>���>�%���� ��{��нZ��>l��>gD?It>sE'��6[�Û��K��>=8�L�=�/i?����I�\���>L�P?��T�rqa<;��>��������G���+�ݮ>3�?f��=k,:>�|ľ#9�^ |�s����j?�3�>�����p�+�>��a?w�?{� ?֒�?3$G=���̙>�Y'?̹?�>?�Fb?�c?˥O>��'>���������X;�xk>��>J�=Y�9>�I���1�V]½*�˽P���N��ν���=��Ž�-����:��=޽ۿ�K�,�־`����m�	��Ȋ��ٹ�TP�����;��ܹ��a�y�lp��U$�R�V���d�k��Xno��?x��?������Mՙ�ꦀ��< ��>�az� yr�~:��"���^���}߾j쩾+#��5Q�~2j�84f�N�'?�����ǿ񰡿�:ܾ4! ?�A ?8�y?��7�"���8�� >)C�<x-����뾬����οC�����^?���>��/��l��>ू>�X>�Hq>����螾v1�<��?9�-?��>��r�/�ɿ`����¤<���?/�@E�A?`)���vN=�r�> �	?�:?>�0�J��`�����>e5�?��?�N=�YW���ye?�#<uF���ǻ�V�=��=�=,I�v�J>=o�>Y���@��ݽ�-4>#C�>AW"�s���_����<��\>hoؽS���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��=�����ȿ�1�p��#��=��w<d���x/�q�)m���]ʾ/����]�Fi�<���=PST>,i�>�H>�B>��T?��n?9P�>�y>]=P�d���!�W������}7��4j�;&'����%*��]�־sQ�}�(�����<ҾU=�	��== R�Fx�� � �C�b� �F��.?o�#>-�ʾ
�M�ƫ%<��ʾ�䪾ƅ������%̾�1��;n�ϟ?�A?-����V�J.�^��-���kuW?���[��U���=x@����=GR�>"!�=(S�\3���S��g/?U�?5���M��è->ި �O�=/�+?F_?���<P��>)�%?��#��|��Y>�5>[��>��>�>R歾�kֽIQ?L�R?���wI��L��>������q���=7>�2�DP伟�X>��h<Z����|�7���j0�<��W?`S�>�*�6����������)6=
x?��?�.�>��j?"+C?\(�<�1���R�c�	�ʚ�=20X?ci?p
> ��W�оK,��#^5?�	e?E�N>�hd�H��%~.������?��m?��?�V���k|��ϒ�.U��5?��v?s^�{s�����8�V��=�>\�>���>��9��k�>�>?�#��G������mY4�&Þ?��@~��?��;< ����=�;?f\�>ЫO��>ƾ�z������"�q=�"�>���zev����R,�c�8?ՠ�?���>������As�=ĤS���?�S�?���mѼ�A�ʪp�ض��\��#��=$ϐ�?R��Ѿ��:��ξ�����������t>u�@a	����>���	ܿ����^���Mm�������>�y�>Rӽ_;��	�R��oy�~T���G�ٯ�����>X�>��F���KDy���8��B=�&�>y�N��܁>�ms����󰥾z�x�6�>��>��a>q߽����P�?/����ο%a��#�価�m?�;�?]��?23(?	�5����W�/�L�=/a8?�3t?��a?��G����ǽ!�j?�_��xU`���4�rHE��U>�"3?�B�>R�-�S�|=�>���>g>�#/�x�Ŀ�ٶ�=���Y��?��?�o���>r��?ss+?�i�8���[����*���+��<A?�2>���E�!�>0=�RҒ�¼
?W~0?{�e.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>�(�?4��=�>�M�=�ڰ��.��">���=�]8���?�M?&o�>��=��8�9�.�@F���Q�����C����>��a?yVL?èa>N[��/��!���̽�(2�d�켡R@�1�*�|
߽`5>۸=>v�>%�E�BӾ��?kH���ؿqc��Nf&�dA4?���>D?A���`u�2��SP_?�M�>8����~���k�%p�?��?��?��׾��ͼ2�>v�>�{�>r�׽j��,+����7>��B?�Q�L�_o���>�	�?�@�Ѯ?��h�	?(�Q��#a~���]�6����='�7?�-��z>���>X(�=�lv������s�㵶>4@�?%y�?A��>A�l?�o���B���1=TQ�>�k?�o?{�m�)���B>�?5��Y����H��f?��
@�t@%�^?����ؿ�3��kș��-վl��=�~�=�*O> �^��-�=	�=�Ss�(�y����=9�]>�ō>�G�>iPz>���>�>7|����(�۴��t����<��6�Y��T�����Z��_B*��(�;���ָ�Y����i���똽x��-�(��C�=��`?{XE?��c?Of
?��F�(�>�f���m";�}��y6
>'��>�1?�?J�:?�o=	�����S�I�}�u<��>l��߆�>`�B>>��>K��>y+�>�,�=-��>%��>��+>�Q�=�=�{�= ��=���>(��>���>;1�>�B<>ʑ>6ϴ��1���h�0
w�y̽6�?h���K�J��1��{9��妷��c�=�a.?{>����>п:���[2H?{����)�	�+�!�>��0?�cW?�>S��5�T��:>}��Ӥj�/`>�+ ��|l��)�['Q>�k?�f>a�t>��3�&,8�2�P�Dq��{|>�36?"��q�8���u���H��xݾ�L>Mǽ>�M�N��얿b�~��9i���y=E�:?�p?jC���U��މv��~���DR>��\>��=��=:�M>+�]��,ǽr�G���.=���=��_>���>U�>��>t��>��~�M�4��>l
>��>��e?��C?��G=���;"ヾ�����>��>��>�r>N�;� `�=u��>w�C>�Ž��`���)F���8�>������k�TqY�G�e=����=(��=�.��Pz�q[F��~?���(䈿��e���lD?S+?_ �='�F<��"�E ���H��G�?r�@m�?��	�ߢV�@�?�@�?��K��=}�>׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�<l�6>�^%?��Ӿ���>��@����G��V�d���`=��>3�P?�*�Y��������?���>���C���!\ÿ��u��l�>k��?N�?�/n���OI�_�?�!�?W�U?�|�>-�������L�>�@\?d�]?n�>N��j� �ۼ?�y�?2Zg?�$>���?�"x?�?�XJ��9�x�������f@K�W���F>�/j=����G'��Y��]��4�q����V)>�e0=:��>�R�rf��X��='	'��s¾qr*��=>�;�=�r>)��>%�>S�>��>�U���ͼլ��\0��i�K?���?���2n�Q�<��=7�^��&?aI4?yw[�5�Ͼ�ը>Ѻ\?}?�[?�c�>]��C>��B迿1~�����<��K>4�>�H�>0$��?GK>��Ծ�3D�wp�>�ϗ>>����?ھ,��QB��uB�>�e!?���>Ӯ=�� ?\�#?��j>�7�>�~E��C���E����>�I�><P?��~?��?����Vc3�����꡿/�[���M>zy?|7?���><|��>����=�AF�������?��g?y@��?O:�?��??!RA?_�f>�a�d�׾W6�� �>!�!?���9�A��&�����?YR?���>3�����ֽ��ڼ������T�?�\?%b&?�R���`���¾��<>���m�G�;7�>�_ >:>/���F��=	�>6�=�,m�m6��fb<vP�=���>��=i�7�^Z��/=,?ϿG�|ۃ���=��r�>xD���>�IL>����^?`l=��{�����x��	U�� �?���?Zk�?[��?�h��$=?�?T	?l"�>�J���}޾9�྾Pw�~x��w�V�>���>%�l���J���ڙ���F��\�Ž�,��^�>^��>\��>��?�g> >�>��`�7���,��E���L��Y�QI�?j/�(������� �9e	�"žl���I��>n
��K?�> 3?J8>c��>���>-�����>��>�Ҝ>�Į>�Y>���>Ø:>T}�=����RR?:���@�'����G����8B?<kd?w4�>D~h�^������}�?g��?�n�?�Dv>�kh��+��r?�B�>Y��p
?�9=�*�0��<@I��)��M������K��>�f׽:��M�sf�Mb
?0?5�����̾R=׽�R�/�<哆?�5??>���>W��;��y�.�i*f�'PX��/��Hľ�pJ��4\��ig�i=��5���B[@�bc��aB?f�?-���ᾕJ+�	Gg��J!����>8��>���>�e�>z�%>�I4���'�yyc�c<�iǽ��>3O?Oc�>�sL?vY=??]M?�J?�V�>x�>����m�>g��<&�>�z�>9:?#�,?u/?h?x�(?(�h>^�߽����B3׾B�?��?I�?b�?K?����tK����f*��Kx�4^�.=��<dҽ(i��3)=�?I>��?)Y�k�8����sk>��7?���>5��>�,��kl�����<u��>��
?߯�>5P��c�q�������>���?����=!�)>k�=4>��E~��Y�=/���=��=uo|�V�<�q$<iT�=UЕ=�n�	So8x;�b;��<Do�>r�?n��><�>7"���� ������=�?Y>y�S>v�>�(پ
p������g�ny>t�?Dz�?Mh=��=���=p���S�����v�[�<܃?�U#?�eT?���?��=?]#?r>1��F��;]������?�z?�\�>z2��uP��l����U�D�>��>�q~�`����C��'�:����>�m� C��N骿E8v��J8�О����;4Q�?�y�?,�3��UK��&���R���u�,7?��>Dm�>�4?(�'��|M�= 
�T`�=�|�>2��?�޸>��S?bLw?b�X?(V>�:��������z�^��>#�A?/g�?]q�?�.z?3��>�s>�5@�+ܾ�m��m�.��C��rx��=�'Z>LD�>��>�P�>��=�wֽ]ⶽ�w*�]Я=��> ��>�ԭ>?�>�e>l��;_�G?ڵ�>so��4u����qӓ@�qu?s��?�,?��$=�Q��VD��&���_�>H+�?��?��*?�{N�<��=�R̼����<s�-��>��>�&�>�3�=GTU=I!>��>;�>D>�m��I�8�23K��	?��E?��=�Y����s�pe�.���U@û>��XPa�.Ǐ�/�G�<M�=RK��ߝ�����LO��ӧ�b����Q��Jf���u���>�]I=n�>`�>��<�{��<F�ֹKd�;�=k�x����l�=����fL��I<��_=DP���ʾc�}?6cI?8+?,qC?	y>��>�Q8�˗>�w��?��V> �J�>��V;�5���L�׾�?־G�c�V���N	>��I��>��3>���=�ׂ<�5�=�kj=�=�c���=���=��=F�=M;�=�I>�d>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>}�>�Z�=��U�a3���?���C��%��;*?34���Ͼ���>9^>&gվ�޾Y��<�.>(�N=u�a�U��C|=�����bf=$�w=Oȅ>�<>�=@ڮ�>�=�e�=6>b�c>�=�ࡻ[g�U�=.>��r>ŭ>Ұ�>(?>|1??M?F�>F�l��,��>�;�_j�>P�]>���>�B�=��>a��>%�7?��A?�eK?+"�>Ԅ$>Fi�>�Z�>z�"���]�[
����'9���_?��?Gz?۳�=|���O���V�XT���?K?b?��>�P�4��xP&���.�1�����ն��*=kjr���T����Z3�j��d�=�p�>���>�ڟ>�jy>��9>e�N>��>5�>qy�<D߅=8R���`�<ɷ���'�=�����<��ü�0����1���*�eV��@�;�?�;`^<���; ��=V��>0P>���>"��=7	���>/>���>�L����=�G��A+B�(2d�6E~�/�i]6� �B>�5X>�x��-2����?��Y>+y?>K��?�9u?8�>�(�b�վ~R���Ze�RWS�&Ǹ=Ү>.�<��|;�\`���M��{Ҿ� �>K<�>[N�>+~�>�"K���Z�~�==�ξ-C�=F�>@.���!7������F��q��O���t���2���Y?	�����$=�Y?�?���?f�.?��j>$��ݝ�>cHؾD.J����g	=�,��,HD?�H(?�C�> a.�jd;�ā;�����>WC�	�P�Y�����1��k������>�d��G�Ѿ��4�o7�����;�C�Mu��>u�L?:�?f_��Q���RO�z��c��
�?�f?ݝ>��?�	?�n��K�ﾍq����=��l?���?�y�?��>k�=A�o�;��> ��>8��?�!�?��w?�E��!�> �p;;�2>g"���>�=�@�=�`�=`�	?(`	?�c?����a�����1�f�O�e�=A�<�Տ>�9�>gp�>�>�E�=���=��C>��>Ț�>}�>�O�>�`�>8���x��j��>����^>y�?�"o>��>���<�[ϼ¢�<6�+�������T���h�Õl=��a=^9�����>B��$N�?��>Q��>����/��mQ>-�>�I�=��:>��,>��?oH�>�X>���>�c>.9�=�(Ӿ@�>S��%!�U]C�F�R���Ѿm�y>����^%�pe�̱��mJ��]�����#j�F0���l=���<r.�?i��sk���)������`?q��>96?����`��
�>-�>��>)���v��ṍ�{7��?���?�;c>��>Q�W?,�?Ӓ1�O3��uZ�1�u�j(A�*e�Q�`��፿
����
�����_?��x?%yA?�R�< :z>T��?��%�Fӏ��)�>�/�$';��?<=Q+�>>*��U�`�{�Ӿ~�þ�7��HF>w�o?1%�?fY?LTV�-dH�{*�>�J?/�(?{\�?p�?HNK?Q��h�?�ɉ>C�?J^?�	9?`PG?��?M�A>�>��=�<��#�;ߚ����$E����� �=#%=�5=��ԼFK=���=�ď�bǴ=ǽŽ�b'<l��=��q>Y�~>�D>�u�>,{j?���><~h>�5?ջ'��J7�>$��( @?<��>J4���p+���R�8��2��=#Cb?I��?�Cc?��>�.�'4뽗�3>Lo]>ݐ�=��Y>&�>�V���f�ݨ>c�=g[2>�gd=�载jl���g���᩾�/8�C>���>	0|>Y����'>�|���0z�C�d>L�Q�x̺���S�j�G���1�؄v��Y�>�K?��?֝�=;_龻,��[If�I0)?�]<?�NM?��?9�=��۾��9���J��>���>�U�<��������#����:�y�:}�s>�1��Oߠ��Vb>���s޾��n��J�&���EM=��UV=����վ�6����=Y$
>������ ����֪�B1J?�j=fw���aU��o��\�>ܾ�>�߮>��:�V�v�)�@�h����4�=|��>��:>�`����~G�8����>��H?#%d?���?�\��'h���8��W�ߐ�ܼA:ߑ?�c�>�?�4>-f�(Wپ��!�St_���)���>L��>p���ڸh��;;��|�d�*�ͤ�>h?�?����?U/?���>^�n?��+?�b�>E�>���gʾ9C&??��?��=e�ԽU�T���8�"F���>^�)?b�B����>?��?J�&?�Q?�?`�>� �M@@����>WX�>��W��c��_�_>\�J?���>P>Y?iԃ?3�=>�5���fϩ����=I">��2?L3#?٬?���>ԩ�>�����=Ϝ�>c?�0�?��o?x��=T�?�92>���>V��=&��>M��>�?�WO?K�s?C�J?��>\��<�9��5���=s�}�O����;H<��y=ʠ�]7t�iK�T��<~�;f��F��u����D�Q���x��;;W�>��s>�����0>��ľ�P��X�@>$���JO��Dߊ�4�:��Է==��>w�?���>�X#�kÒ=˰�>G�>n���5(?U�?y?�5#;Ɵb�>�ھ<�K���>B?��=��l�������u���g=M�m?��^?��W�\%���jf?]�e?�����9���꾁�\���HGa?�G?�
���Ȩ>�-v?���?�?C�f�n�n�D؞���h��W��$S>Hl�>��6�
���S �>�yS?���>5D�>��z>
��\Y��
��^L?ާ�?��?��?ӿ%>~~M��ܿ����񑿕�e?%2�>,J��r_?�켬q㾞E�������������%n��矾!�%��@�����c=��?�w?�j?�AU?f����g���Q���|�LJ��9�f���?�Q�D�QAL�8�m��Q��i����4��8�=YKf���L����?��2?O/�@�?���cN���Ӿm�>�	���F��82=I�g���C=��=̈��u����̾U�!?y�>F��>ff4?1p��>��"�,�E���վ��{>��>���>"��>#��P'e�pн����d�Q���x>��b?L�I?-x?&�Ͻ"j7�T~|���'�������V1>�2>���>dc�~:�g�'��D�	�r�(C�賏�	���r�=.�.?��>�H�>[ؔ?���>݄� _��,|l���-��Ӻ�$�>�e?m��>�و>HŽ��*��y�>_��?~B�>?�R>��ɾ�-R��+��o�p	:?w'?.�?pH?
��=S�I������I��+G�(s�=��?0Bj�����3d>��?�=����&?C
��k#�PY��V�D����>Z?� �����>������0�Ẃ��_b��R-?�d?<~��2_=�M-�>��=?M|�>%�>,�?�G�>�ȍ��= H'?��h?�1?^j*?�J�>�h<� �`U��8�dP�=�y�>�)b>eɎ;k�">�޽l���'�3�{��=��->9�<�ٽ�%��mɼϦ�<�;=3qz>Giۿ�DK�	�پ��(�@
�D
���(���b��U	�w�����&ex���G�&�4V��c�����l��y�?*+�?pn��c.������b������ĵ�>��q�ҏ�����J�Vx������Ҭ�VY!���O�Q�h��e�M�'?�����ǿﰡ��:ܾ,! ?�A ?A�y?��4�"���8�� >�B�<-.����뾦�����ο�����^?���>��0��w��>쥂>&�X>�Hq>����螾p1�<��?;�-?��>�r�.�ɿ]������<���?-�@zA?��(�t��OtU=:��>��	?�@>1�N������p�>�6�?H��?��L=�W�A�	��ye?2�<<�F���ܻ��=@�=E�=k��!�J>OI�>�����A�*ܽ��4>�ޅ>R"�~��R�^�O5�<�}]>��ս�������?�W���t�n2���h��C0>��f?T��>~��;��l?� <��|ο3vU���J?��@n��?`� ?� �!�)>/@Ҿ��@?oV?d��>mX,�Z����̉>l����>>jܾr���]N>�z�>Q�>�>D��!�,bI��e�;Q
>nC �M(ÿw��DN�d荻�ؼ	iý&��;p����ϽX]��9�u�p�ի\=l��=OJF>�Ƈ>z�c>��Q>ݿS?�/d?���>l4>g���o�������R=�;������#S��u�E�~wȾj��$/�����z����0���<=��o�=ΚQ�����I� ���b���F��X.?��#>��ʾ�MN�X�<d0˾����3��c���2ɾ=�0�_�m��ȟ?UB?�˅�2W�S��:��i����2X?e���<[�����=ah��|)=ZL�>�o�=?��S�2�9�R�a�/?� ?Jg���L��nKG>1�˽}�<=[/*?<?O�W;>��>a�'?۸	��6���7V>H�(>�>sJ�>��>0���a����K?
V?����ߤ����>oC��96����>=ö�=��#�:�#xX>�9�<��|-��G�}�Ͳ�;n�U?��>h�+�A���4��gJ6�~=��{?� ?�>rl?<�A?��0<����P�Ռ	�DM�=uZ?�#i?>c���׾m���t6?�(f?�O>v�l��f�}'-�ئ��		?�n?��?T��L�{��`���&�] 6?ىh?X�U�m��R����4$���>��?�Y?�=m�ԗ�>��l?�V�9��9'ÿ�N��Ҕ?N��?�H�?QG>׎=,7=b��>K��>���O�Ͻ�)6��$��<��? Y�.�s��V�V*Խ��)?g1�?���>�d��,�����=Z��Gi�?��?u����l<>���2l�<s��P7�<Lժ=���� #����z�7�?�ƾ��
�tӜ�eļ���>X@����>W�8�s5�u2Ͽ���-оr�p�X�?j�>b�Ƚ�磾��j�u��7G�a?H�.1��H�X>W$�=�w��u�ؾ.Pu�W�;�^�5=�{?ep��opR>�W����ھ;uؾ_��ƨ�>g-�>:�?�=�}��*�?�(Ǿj�Ϳm����y(3?B �?���?��>�5�=��<%���}Ҽ�� ? }?�8?z��3��!�=%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.���_?)�a��p���-�o�ƽKݡ>׾0��a\�8d��ך�We�a��XCy���?~^�?��?��#� 5%?��>񝕾�5Ǿ{!�<��>$�>�+N>9_�}�u>��N�:�"h	>#��??~�?�j?ŕ�������S>��}?o��>���?��>���>�C�>�qi���)=�>T$>p��><&[?�?g�^>58��9*��C���<��N�2A�$C>�e?ÞX?��+>%�1�g�L�RW�L�0���=�q�{��wҽ�D�"ĭ���+>��>lW:>b��h*����?Op�P�ؿ�i���o'��44?"��>��?A���t�}n�i;_?�x�>�7�m+��V%���>����?QG�?G�?|�׾�p̼P>B�>L�>�ս��-�����7>��B?�(D���o��>���?��@Oծ?�i�vI?d��Fŉ��fz�x��7��7>Y�:?!���B�k>7?�Y�=P�u�����>`n�pM�>G�?p��?V��><,k?�k���D��z8=;>�>iWn?A"?���m���O>�?DG�2֋��<��^?�D	@��
@$�Y?����ֿ�o��󒾳�j�K6�=��==v,%>ṗ���=KYӼIZ�,��=@Z7>^��>�>>��f>UMj>��?>��[>>��Y[���������F�p��.���|f�����G��F��Q��f��Ǻ˽��X����<�=i�~�%�"�����=�U?�R?b�n?-�?W�m��W >�����==�%����=ξ�>J3?BWM?
�)?K��=�ǝ�[�c��%��+���=��^�>f\O>���>��>X��>��8�8G>�<>>�s~>!n>��'=��N��=):M>σ�>��>p��>D<>)�>2ϴ��1��T�h�
w�/̽2�?���Y�J��1��v9��X���k�=Bb.?�{>���?пi����2H?����)�#�+�L�>}�0?�cW?��>���j�T��9>r��<�j�v`>h+ �l�~�)��%Q>Al?ԡf>0u>Ù3��N8�f�P��v����|>�-6?��?n9�P�u�ùH� wݾ��L>���>"ED��o�O�����b�i��'{=�y:?��?����ΰ���u�Y)���[R>(�[>vU=�ū=�]M>R]c�X�ƽ��G��(.=E��=v�^>�W?��+>[��=_أ>o]��|<P�ڇ�>Y�B>5,>�@?�*%?�d��˗�Ƅ����-�iw>�Q�>
�>!a>vYJ�F�=wj�>c�a>�>������z�?��gW>��}��x_��Ru�P�x=3�����=i"�=� ��=��%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿhg�>���S[��+����u�u#=��>AH?�a��%�O� �=��t
?�	?_i�ڤ���ȿ�pv����>.�?���?E�m��C��@���>���?'eY?[]i>,z۾\Z���>T�@?�R?S�>�;���'�k�??ݶ?���?*\N>�8�?��o?Y��>S7��4��䭿AH���Қ=(+�=޻�>��->�ם�V&A��H��BC��n�k����xz>�$%=�J�>�������8�n=߳��` ����2�ɤ>��F>,f>3��>���>n%�>�y�>2�<:�{�_�u��6�� �[?��?<��l���U�>B`�>�.��?�K?C���'�߾B�>�yr?�Ö?��=?�!>�@�Ḉ��й�1d����A=E�=q�>�B?l��<mV>Yy�w(��ļ>T�>�ц:f�cr��=~�����> �?o��>�[c>} ?lB'?�u>ͩ>d�C��$��4$I�m�>O�>�?5�}?�?�⭾�%.�)���Ԣ��;Y�"�P>jw?ej?�ݒ>����^����S4�L�� ʙ��|�?�e?S?��?�?1�?C6>?3??g�k>����.ݾ3	˽���>u�!?v�-�A�lN&�/���?�P?���>5���ս��ռi���z��� ?E+\?{C&?f���*a�#þ�5�<~#�r�S�O��; �C�ί>T�>�v��ؔ�=�>�=Qm�`<6���g<y��=�z�>���=�/7����*=,?	�G��ۃ�7�=��r�QxD���>aJL>�����^?zn=���{�����x��U�� �?���?k�?��G�h��$=?��?7	?X"�>�J��L}޾�ྈRw�k�x�w���>���>A�l���a�������QF����Žk�7�3��>�\�>q?��(?bo'>��>�k��U<��g�
����j�[+*��qF���R
�9ľ!���-���Oþ��j��>.����>:S?���<�>�7�>�ڽu�>�e�>�<�>���>\�~>�HV>u�=�!�����LR?����m�'�z��Ln��5CB?�hd?)8�>��g�񄅿�����?8��?1x�?�0v>sh�f0+��Z?E�>#���Y
?��:=V	��!�<�]��٨��J��e��)��>�g׽�:��M�~Cf�qc
?�?T����^̾�׽]���6g=m��?�T)?L�)�@Q��Yo�	X�k�R�����h�����9�$�Qp�����A �������(��v$=�a*?�e�?M9��V��אk��>�Gd>~��>�)�>���>�3I>u�	�k�1��^�x�&��q����> X{?�u�>�qI?�A;?<nC?�R?�(�>q&�>����6�>��5�>�� ?jC?b=6?h�'?�?�B?g�a>�x�#k�$����?%�!?A�?#��>>>�>�)}�4�@z���4��M�l�c���D=�Gq<R��S��,E=k�7>�?�B���!6��T���>hU;?^7�>)��>�Ǉ�w׀�g^=���>�?]�>j����to�A�� D�>�΁?8^&��I�<$1>���=Ssf��8����=�鍼�i="n��u�6��y�<v�=VZ�=`o���H�jg;ܪ�;��<
'�>�Z<?X�>v:�=�������8�xk�Ѩ�>ս&>��=U���Lk��ڀ�%��.=P��?K��?�=ƥ>.�q>׉侉���������:���>�(O?Ay?J�?T�)?r�&?�'�>��%�Qh��� ���\��1#?w!,?��>�����ʾ��Չ3�ܝ?i[?�<a����;)�ސ¾��Խӱ>�[/�g/~����=D��텻���S��5��?�?IA�W�6��x�ۿ���[��x�C?"�>Y�>��>U�)��g�s%��1;>���>jR?���>=�O?��z?�d^?[Y>ַ9�2����D���#*�#},>��=?�%�?w]�?<v?&G�>q>w4��7⾆��Dc�K�3;~�W�@=6U>Á�>)��>d��>K��=T;۽�s��u�<��1�=�k>��>!��>.?�>}w>"N�;1�:?�>��龻���B���*�����=�Ջ?n^i?��?���=�0��M�w���;�>?��?�z�?�B?�罌�J>ɱ��X�����j��>Z��>ҵ>H�==� �i>[C?l�>�1�������9��$н��>3I?��>g�ſ*_q���j��7�������t����w��鸽;"Z� e\=G����������yCO���>�����H��,�v����>���=Uf�=U�=s��<�Լ���<�JQ=��B<���<B�������4(�.���MT���=�e�=�!��˾}�}?�5I?ѓ+?F�C?߻y>^G>Um3���>´��-9?�V>�P�D���V~;������'��,�ؾ̓׾zd�bП��d>I�g�>703>�=��<:�=�r=���=�jJ��2=�"�=�`�=7p�=��=D�>�Q>��q?�Mq�����<:A�G�W�o?�c�>��=7��͜d?M�>/���"���h���?��?	)�?@�>��ýo�>HŬ��C�<�N�=0	�k�8>�î�G�B?��>P*��t���އ�c��?��?��D?+֏�\�ӿ�w���E7>{>��R�b1��~\��b�|�Y���!?�n;�bw̾jW�>Jh�=�Y߾��ƾA�.=�l6>�d=�R�&\�)��=��{�[Q9=��l=�(�>��D>��=�İ���= J=:��=t�O>��1L;��.�v5=O��=��b>�&>���>�?�a0?RUd?24�>�n��Ͼ�A��~G�>s�==�>̅=�fB>Q��>��7?��D?��K?���>2��=r�>|�>��,��m�hj徹˧�,Ĭ<���?*Ά?�Ӹ>��Q<��A����%e>��)Ž�u?(T1?Yl?E�>�����ѿ��uھ�d������9X��B���=/�1��hY�l64���<���>� �>L��>@]�>��>Jֱ=6(�>�}>�J'=T`O�l���~�Q��1�OF��^S�%���ԥ��~3��rN����G���XQ/�ɀ��sn=P����պ=���>.��=;A�>0�=���ܐ>����b�[��]=������P��vl�� y����1�4���=�=�	T�Cё� ��>� >��M>���?�/q?�w�;ӱ��� ��}�%���p���<�Z<"���TZA�Û_���L�%����>�ŏ>W_�>#_r>�+���?��Fv= ���g4�^��>�|����	�h!�fq�2��Tԟ�i�i����ˆE?k��Y��=}�}?�I?9��?z	�>�Z��L�ھ��*>T���"�=O�z�o��5��E�?�'?6�>��0�E��T����+�c\�>��s��@�P ��1�7����������H>#8�oe�lo;�;���PЃ�mS%�%3����>��2?��?�/���
d�AiN������� w?lFj?2�>8?�>i�"�N��5��Ú�=U�s?ݢ�?E��?v0�=��=+L���*�>Z	?|Ŗ?���?�|s?]?���><��;�� >���3/�=O>�c�=[��=[?2�
?��
?ʾ����	������ ^���< �=�>�A�>pcr>
��=�h=Ր�=�\>�ў>?ӏ>��d>5�>�G�>>{��R�"$?�؆>?�,?2�D>��=�a��[>���,Bp�������!��^�=�k�JT�fSx����>�ϿU�?��M>= (��r(?fo�42����>�|b>�B4��i�>��>���>bo�>O�t>�>�=^>��{>,FӾ~>1��e!�-C�d�R���Ѿ�z>t����	&�Y��~x���DI�vo���f��
j��-���:=�ڽ<1H�?�����k��)�-���A�?H]�>�6?�܌������>���>�Ǎ>uK��5���Kȍ��hᾥ�?���?$GN>��>��v?9�(?(�R�l>q���H�mw��%�5��BW�K�Q�Ǜ��U�o����W�,���D?�gq?�0C?<���Ji>U��?͐+�Qs���Ц>�:@�1l6�B	'=�%�>���m��Tr��2�Ⱦ3/g�4��9��R?���?Yrf?�+��O���w�3>�OF?0�2?���?��1?NP:??$	�F#?-��=�?�|?��9?��??��?���=Y{�=~����;�|���葾&���z?P��r?��ዻ]j�=��-���=�o~<'����������H�/<��%=��U=���=TH�=���>r�]?�L�>��>��7?����~8��ծ�0/?g:=h���4��#Ǣ�����>�j? ��?0iZ?Wfd>1�A�9�B�>SI�><U&>;\>�W�>S\�WsE��@�=�Z>Gj>��=�3M��ҁ���	�����T�<C>��>��J>l<Ƚ�.e>t{�����|��>��T�T�����x���`��A;��}��O��>*U?�w"?
eA=�
�#|��)w���0?�E,?�=:?�Ā?�3p=e�Ҿ<:@�׃a������?�>E;v;�������[�� c�[`)�F$>@�׾L࠾Sb>A���s޾��n��J�B��|5M=z���MV=����վ�7�ܟ�=�"
>K����� �"��dժ��0J?��j=s��[U��r����>���>�خ>��:�V�v��@�����.�=A��>$�:>�}��� �^~G��6�|�>�qE?��^?"�?BR��x�r��ZB������v������$?���>,�?(�@>V��=Y��O�r�d�܃F���>K��>���ĐH�I֞�����$���>o�?�T>\�?R�S?�?J�`?:�*?�!?Qܐ>�N��]G��VB&?o��?G�=M�Խ��T�k�8�[F�6�>��)?2�B�Ҹ�>m�?Y�?��&?�Q?v�?��>¯ �MD@�f��>HY�>��W�Ya����_>��J?���>#<Y?�ԃ?.�=>��5��颾�٩��X�=	>�2?S6#?��?���>v��>����Y�=��>�c?$)�?>�o?��=U�?��1>[��>�ٗ=7��>Ԇ�>��?�2O?v�s?�J?�W�>̧�<f2����s���P�P}�;߆L<�^z=,����s�P����<Jl�;Ly��0f��J��D�1������;_�>��s>]����0>��ľ�O��C�@>����PR���ۊ�'�:��ҷ=��>O�?���>8V#�I��=��>OI�>����6(?��?�?�\#;��b���ھ�K���>YB?���=e�l������u�4�g=��m?[�^?��W�
'���b[?M*l?4TѾ��D�@kݾa�	�� ���HJ?��?gѤ�zd�>�V�?|�y?�c�>�p�]Iw�m��Ǩn�:�'?>㻛>,��C�d�%��>��8?>H�>H��>p��>`G�]i�݄��a��>iއ?�)�?�N�?�>��a�n�ֿ6D�4����`?z��>(�����!?�2���پ@đ��ǉ���߾􈶾�l������R����$�6!�����h�=��?�o?�v?-�[?	�*�d���[��ƀ�_@X��m��z�?F�	�?�gA��1i�sU���徽.���'�=�$h��CD���?��?T�1�� �>�*�����aҾ�wE>�J���-K�"�<$���1�=��4=�/y��3�+]��:�?���>��>��7?i3f�[�A��5-�j=�ū�"�s>��> y>(h�>����)���r��
���-Y��r�q=v>�wc?��K?ѷn?'X�:%1�C���M�!�d�/�f����B>h>�ʉ>,�W����X:&��T>���r����:z����	��7=ɱ2?0(�>˰�>�M�??�|	�uh���kx�I�1�~o�<4�>i?�:�>��>��Ͻ� ����>&r?7i?6�>�ݾ�`��ZO�x����9�>w;3?�v�>��>>g=$�#�w��՗��/����B��l.>mXh?�<s����%D`>��a?A�Ƚg@>�?K�ھF�`Ͼ�G���F��WnL?YE&>l������6�4�y�����ʽ_=)?NU?���=�*�s�~>M"?Zj�>�	�>W&�?,ݛ>7vþ;Yn�C�?W�^?0-J?]KA?	�>a�=����=Ƚi)'��1.=J��>��Z>*�m=ܫ�=�T���[��k��E=��=U�μ����%*<n�G�K<~��<�3>�qҿ$ P�l˾���a���M�� ���ڨ�}�ξ���`���)��ELa����5�/�Z�h������`�W����?A��?ô5���8����� }�����r>��>�+aZ��{�V"Z������ؾ����i�$U��q��KY�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�|A?,�(����DV=���>:�	?��?>GX1�nF�p����U�>�<�?L��?��M=o�W��	��~e?�?<p�F��8޻k�=0K�=l=��1�J>�S�>A��EXA�6ܽ��4>م>`k"�N���^��_�<��]>��ս�4���ȋ?WG]�c'u�Е,��^��/?J>�/Z?|��>�B���?�u�u�ѿ�h ��Z�?y[@~V�?�-?3��?�����G?�@?��>��W�鐿F�>S|���5��$�˾�t]�7eF>�f�>)%�;ב��L��U��� �=�F�=8����ſ�,!�z%�:��Z3��Q0^��h��ƂB�?�Af���UC���нr=�=�?(>�j>�;M>��b>ff]?�m?�.�>k>�!��������������ZG��^v�X#8��������(�Ⱦz���!x���"�Ⱦ?!=��	�=�6R�T���Y� ��b�D�F�g�.?�q$>E�ʾP�M���-<pʾۿ��T݄� ⥽4.̾�1�i!n�V͟?�A??����V����o^�,����W?vO����X鬾���=����t�=�$�>͊�=D��!3�8~S�9w0?;�?[��������,>�H��$S
=b�*??Q?F&;<��>a�%?uZ%��߽p�Y>cE1>�a�>��>ٛ>�Z��3߽6�?JU?�������	v�>q���[�|�w�k=�>�4��$Ѽ�\>���<�ɍ���0�����)�<'(W?U��>(�)�)�b��3!��9==7�x?>�?�1�>S|k?o�B?���<k����S����fw=<�W?"*i?n�>����о�{����5?��e?��N>�eh����-�.��U��$?�n?�^?����zw}����7��n6?C�v?Qk^�������V�2��>a�>]��> �9�1K�>�>?�#�!P������NL4��ʞ?�@w��?�<<���8�=�?�Z�>/O��ž�A��߀���[r=En�>Cr���rv����9�+���8?:��?�~�>Oꂾ���}�=#ە�%X�?v�?F���f<V��fl��y�����<@ҫ=���\"�5��r�7��ƾz�
�=���F��J��>�Y@c:轙-�>�U8��4�XQϿ��Oо�5q���?�v�>c�ȽT�����j��Mu�βG�4�H�昌��M�>\�>봔�.���u�{��q;�7)����>��	�>�S�:&��Q���ba5<��>���>��>4(��潾Vř?mc��5@οr���p���X?Th�?�n�?q?�]9<w�v�_�{�g���-G?߉s?�Z?D^%�K:]���7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�pq?��e�8��h+�rQ���y?(���@�4=W��=%$@;�JV�����������?�@$��?iRG�o�A�]o*?7�>��_�9'd��>SY
>�~>�،>�zy���=��,��t����'��?.�@��"?M4��d������=U�?��>[�?Hr�=�|�>��2>����q�Rȭ=Z�;>�����?��V?.M?�>��<��Z.��7�OL�C,��?��R>��j?qV?��>|"Խ�=�f�+����2���>�5�B�r�C�"���[�/>��>��%>���c�����?7p�0�ؿj��~p'�x54?��>�?���t����;_? z�>7��+���%���B�\��?�G�?W�?��׾�X̼Y>I�>3J�>��Խ����C���8�7>>�B?V��D��q�o���>���?�@�ծ?hi��?uZѾV���[�
�Q]��T#>А=?�	��f�=)Z?YB�=�僿] ��3�h�GJ�>
��?���?��?ʬ�?<�w�qty�P�ὦq�>8��?�8 ?��<��˾���=��5?Y��j��JoѾ0�y?�b@<�@�3c?) ����ڿ����`��_뷾,���	T=�~�>S������G��7�M;je<�">lF�>��>;�7>P�V>�f�=r�s=�M���\ ��������0�W �,a�]A�%r���������ҿ��S���)ʽ��i���Yx��$��*����>#�Q?�R?A�n?/�?�0¼c>>�P�=117�p�=�[�>�I:?H�P?�!?�s�<�����X�|x���;��Ii���4�>�p>"�>���>Td�>r�<��A>s�:>�n>���=�a�<�8<��N=L(>��>}'�>��>'E<>��>�δ��1���h��w�W̽H�?���n�J��1���7��d���@k�=�a.?*{>��?пM���B2H?�����)��+�;�>��0?KcW?l�>����T��9>o���j��`>�* ��zl���)�$Q>?k? �V>׉�>�7���+�I�5�����Cz�>|1?�����]�Y�v�E�M�J���*<>�{�>|��<���_w��[s�y+g�\q�<�B5?�5�>8����S���~������4o�>: J>d�]=�>�,+>VG��>��ۏ=���<��=�5>PV?k�+>���=�ݣ>A[���>P����>�|B>A",>�@?%%?���|�����-�w>|L�>
�>�X>�XJ�sݯ=�n�>�a>LB�O���L��J�?�,�W>
~��z_�Pu��x=�+����=�=�� ���<���%=��~?!T��� ���Q�}���SfD?C? ��=`�4<�;"�j3��㻾��?�
@}�?#;��V���?F��?���=I��>C�>�`Ѿ�pS��\?
�ǽʡ��R	���&�I�?��?S�2�ʠ��\l�>�G%?�Ҿh�>�w�mZ�������u�<�#=���>�8H?)V����O��>��v
?�?�_�㩤�u�ȿ|v����>k�?���?(�m��A��@����>I��?�gY?�pi>Ag۾�aZ�'��>��@?R?G�>e9���'� �?߶?���?��Q>�/�?	q?
�>j[ҽ�K3��˧�z��O��;���=1�>���=pO����I��)��'����r�����ϒ>�wC= �>w�r�۾�g�=s]������6���ϯ>q,W>D7p>D�>���>t��>�?�>�ב��j_��u��(ř��<L?"��?���`�7�3=NC>#�%�X] ?<�V?}:u����0�>%9e?��k?�\2?F�h>���+2��/5ſ��7(�\�>չ?Nr?��o��E�=>����>�!4�>�t�>����v����W��M���n>�:?���>�͆<�?L
.?{+i>8��>-�<�#��E"��wN=�W�>�{3?�}?F�? k�/7�W���'����j�c	{=�v?�s?k�>���y(���+�=Ѝ>G-3�6,�?~3k?^��=?9:�?[??EoE?��>?|G��̤�6Q�����;�?�?�ΈB���#�/��vm?ּ?^��>�A��f�罯��>R��'����?�#Z?|�&?�>��Tc�³��t��<�E��V�:׵ <hi(�C!>#� >4!���h�=��>"��=��^���8�սu<Զ�=ζ�>��=+�3��/��=,?�G�*ۃ�z�=I�r�pxD���>�IL>�����^?Kl=�	�{�����x���	U�� �? ��?xk�?����h��$=?��?5	?�!�>�J���}޾Ӕ�[Pw�@}x�2w�7�>���>��l���L�������zF����Žzd���?6x�>>A?�?1D>
�>��m�:b+�ؤ�p��?i�k'#�^-+��������p���z��� �����l�}��.�>>�B�k��>?�?|�E=��;>�$�>#���瀏>o��>&�7>�N�>k�U>�)>���=�����KR?|����'��������a3B?�qd?{1�>�i�L��������?���?Ks�?=v>�~h��,+�Nn?\>�><��Lq
?�S:=�6��=�<�U��V��*3������>E׽� :��M�nf�jj
?�/?�����̾�<׽������2=~�l?.7?��Q�C�b�;t��b^�s^�:!o=���g҉����[�Z��W��(�|�$����8�P<�=��/?��?�!���.޾����q�k��e��l.>��?l�>���>�e.>���[JM�.Pq��"���s����>��?�&�>jC?&�7?�
L? �X?L�>���>�����@�>_꿽Mذ>�p?�,V?��:?I�?���>s�?bA>y������s���;?v�?�d
?���>��>��3�`����;����h�������v>�6�=����>���=��=w�=�X?V���8�����k>:�7?M��>���>����-�����<o�>��
?�F�> ��}r�c�LU�>g��?Z��p�=��)>���=�����{Һ�T�=\�����=�6��5x;��z<��=I��=�-t��怹{�:☇; h�<)��>�f\?��>b��̠��v�G�����=H>�m>u��><��>B��w���l���_m�٥�>�p�?'�?���=R��=�w�=���M��ʙ�^h���mͽ�?�?T�h?)��?6{�?Δ�>h�);}m��R��[ ��gR��c'?u!,?��>�����ʾ��щ3�ڝ?`[?�<a�	���;)��¾�Խϱ>�[/�a/~����>D�텻���J��1��?鿝?_A�R�6��x�ڿ���[��x�C?�!�>Y�>��>S�)�z�g�n%��1;>��>gR?�>Y�O? C{?�[?��T>Yy8����Cə���,��!>@?4��?d�?Gy?�j�>\e>l|)�����o���[����X=�Z>ց�>,�>��>A/�=D�ǽ�:��J�>���=/sb>���>�l�>I��>Uhw>_��<��F?'��>����k|��z��p!���MZ�J&p?U��?��(?�^�<�`��XG�*V�����>%d�?6��?��-?�Y�Q��=�>��4����h��u��>
8�>9��>���=�Y=�>/a�>"�>���&��9�8��s��?��F?�t�=Yƿ�t��t�=b��O�;������`�B�~��h�5��=�������𤾷�T�a�ԕ��p�������l���?�B�=���=�=��<��鼑4|<N�7=���5�<̪a�X�8<j\C�����L{��$���;%�%=r�P��Vʾ��|?��G?~�+?G�D?ҝz>)S>��2�Ö>�=����?�T><�W�i�����8�9I���Z��_ھ�׾.c�!̠�41
>�G���>74>M�=W_<�K�=Z�j=b�=L{����=4�=4B�=�N�=Q��=��>�X>"�~?D�~�]���hq�kL���U�?��>>�� >|�=��8C?J� ?��p�yK��4���u?TC�?���?�|�>�D9����>����No>��>��}>��������>e��>:U?�����i@=���?�[
@G5?�{��IU��A�=�d5>��	>_9S��k/���O�Q�_�W Q�D:!?��:��,ξ�7�>��=c�ᾗsž(@1=�1;>�GF=͂%���Z�a��=H:���B=��m=�߉>@�G>�n�=�+��ե�=�,D=��=n�W>�`�6r4�����p4=c��=̍_>׸>e��>Y�?R^0?�Pd?'7�>P-n��!Ͼ�I���?�>��=*�>S��=MB>B��> �7?��D?k�K?���>C��=��>��>��,���m�[徣̧���<m��?}͆?hŸ>=�R<��A�I���i>��JŽ!o?7U1?
p?�̞>�����ڿ$�n�-�rnt�5�<%�=Gǀ=���=t6�>hRS���E=�:*>,܆>�EH>�5=�=V�V>3��>��>+�>΃Q<����l)*� z.��Jѽg��=�d����<��E���=����aU�������K���%��G�<<�=�p�=^�>���=���>ez�=+G���Tr>-挾�T��k.=B�J��ld���u�R�)��`��+>��4>6];��>����?V>�OE>mC�?�s?��=A`����|���E�O�b���A=p8�=�B]���6�Or_�[Q�ێܾ1��>���>+�>}Xm> ,��6?�8�y=�a�ms5��b�>�\��c�����?q��K��%���H,i��R�ҽD?3���o�=��}?#tI?;ُ? ��>`����ؾ5�/>�Z���i=���'�p��钽��?X�&?(l�>53�<�D�E�ľ��H�9��>#[����]�����8���
������>j쌾޵��32������-�:��ŗ�<ò>�n?a��?�6������Gb�;���=��?�Zt?=�>�w�>_
?0E@�K�%$��G�=�w�?���?҄�?!�9>V��=(*���A�>�A	?Q��?���?Bs?�]?�@k�>j�;ܤ >�h���x�=�>���=���=�a?�|
?�
?
(��	�	� ��'���^�Gq�<���=K��>��>�yr>\��=�2g=�<�=�#\>�Ǟ>�܏>h�d>���>� �>�"�����#?��=�d�>@�.?̌�=����9t����2����Ϯ��c������s���Z�=���h��s�ཌྷA�>J�˿��?c
�<��$�gS?Ϻ�=�H����=Z�>t(�r�>�>S:>�<X>��>~/>=o�>�u�=�]Ӿ��>̑�LR!��~C���R���Ҿ��x>�朾J�$��F�����DI�W���H��bj�1H���J=�-}�<�@�?@��N�k���)�#2��`1?Щ�>�6?﬋�k�����>O��>���>�7��ޘ���������� �?���?���>wҳ>A�T?-��>j^�������o��듿�ZQ�W���̓�პ�1����M��m����?�p?�qJ?H��=1QE>�B�?��B��灾�C�>r�R����"��=�4�>[O��u���N;Ⱦ@ݞ��SF�>#>���?hM�?iG?GsC���?=���c�g?s��?��?�n?�?�6D=?,�b���>�hG?	GH?܁ ?���>a"V����=Wo�=�z���k(���e�>.������5������m��=B��=	~<8��<�=�� �D���-b2�)C9���=��<g!}=UJ>9�>	�d?>��>Y�E>�P5?�t��8���ɾv?H�+<
|��n*��R�þ'�����=��y?���?�r?�>� :�9��t>~>� >�cP>�u�>Q�����/��L=�^>�3>�\�=����������7
f�|=�B�=t�?�y>^!~�~7�=�SӾ���*�)?\a�\�%���z��w���E��_�F��>x{W?��#?�М=�����=շ����U?[�?��E?���?�K�=\a��dQ.�aI/�"��0��>�;��4UG�R���N���|�����'>]~־N۠�^b>|��q޾��n��J���羥M=�z��V=U�^�վ1��m�=�
>����� �E���Ӫ��1J?��j=ł��|�U�ej����>�Ș>�֮>��:���v��@�����Tm�=O��>w�:>S������Q|G��5�A#�>FE?�Y_?}D�?j�����r��OC�;�������sѼ��?�«>��?y@>��=�=��W:�N�d�I�F��[�><�>I��8H�6���[���N$��>?N!>�1?XmR?�'?�`?"�)?��?.��>^��������A&?%��?q�=2�Խ��T�z 9��F����>��)?��B�m��>`�?�?e�&?k�Q?=�?��>� �oC@�3��>=Y�>�W��b��6�_>��J?���>�<Y?�ԃ?�=>��5�	ꢾ[ҩ��Z�=�>(�2?�5#?�?ǯ�>x��>D�����=Ξ�>�c?�0�? �o?���=>�?�:2>K��>Q��=���>j��>�?MXO?:�s?��J?��>1��<�7���8��Ds��O�`Ȃ;�uH<��y=��3t�K�]��<"�;Dg��I������D�g���e��;tZ�>t�s>ͳ��)F1>��ľ�O���4A>x��̍�������:�R��=	��>�?���>l#���=़>�K�>��~K(?��?�
?��;��b��۾��K�=R�>�A?=��=J�l������u�h=&�m?ߚ^?(�V�g����td?~2V?�ܾC�{��)/���+��lӾ	S?��?�����;=��q?�Ȍ?�<�>��o��y��W��@Vd�gm���[>h�>e�'���ռ}>3�M?�p9?6�;>u�=���<1g��҄�6�>�<�?�?D`�?UB�=�9]�1Vƿ����<��V]?���>\R��@!?��G��yӾ�܍�ݍ���ྑ���Jb���T��l���$����&ܽ���=bD?��t?:q?�Y]?x��kbe��7^�hV����R�#U����;F��wD��fB�EEo����t��S����q=S]�ʕK��w�?�/?��̽�L�>1[2�u �͡���>*�����2�<l�=�ƛ���8<���=��q�]�S���̾�%?��>���>%�.?��j��u>����7�>��ξ�d>'%>z��>���>�N�<!I�Ax����d1����>�v>;sc?H�K?��n?�0�(71�[����2!�o.��٨��RC>��>��>��X�1��J&��p>�2�r���������	�xd=�v2?���>�̜>)�?k�?w]	������y�'n1�Zق<��>i?j*�>1ˆ>��н�!�*��>��e?a	 ?�1�>�R���v@�1菿ʥ�>���>��y>:�.?7��>��<$7o�����ʓ�A�H��6�=�r?����$�=��4�>#k"?��>8�=��ؼ�)�y7 �w/�E���@X�=h�?��&�o�>�Ԉ��q$���{�
m��~�)?"�?����T*���>�u"?5��>dТ>i��?ܚ>�ƾ�.&<Y?U�_?Q�H?��>?���>M�<"پ��Ͻu�)�s}C=� �>CT>m�?=lm�=P��~+Z��V�R_=S�={�ü۩ǽ;�7˼���<�=�n;>�޿��P�8z;h$����i��?Y���x%�=��.+�{⫾9~��g��$���)���#`���V��f����L��}�?�v�?f�U�\��������k���>��0��\�WУ�tL�M���m�ܾ��Ӿ��#�U�N�0zV��K�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�|A?1�(�&�쾄V=���>��	?��?>zV1��J������S�>�;�?���?�yM=�W��	��e?:�<F�F�V�ݻ��='=�=�I=���J>ZT�>C���NA��?ܽв4>�م>��"�ݩ�i�^�J��<o�]>��ս|+����?��Q��|�m(��mt�];�=��Q?x��>�.B�ق^?��*�[�׿�oJ�IY?�@ =�?ߪ!?��g�0%>��ɾ��;?�9?dI�>/I8�/��n>�R�=g�����bR���;mC�>ڛk>����(�����'�dr��F�Icɿ��!�}��o�<���<��ѽ���Չ� @�¨���k!�#�ý�Ĳ=�\>¯1>A|>�!>*f>��S?߀|?D��>�k�=�2�$Qž������2G��RK�O��8*�B+���Ӿk�߾>�������	�Xw��p =�-�=Y6R�Q���v� �;�b���F���.?<x$>'�ʾ��M� �-<Snʾ���0�w襽,/̾(�1��!n�f͟?5�A?,����V�����Q�Rz����W?P�ú��묾���=������=g%�>ډ�=��⾄ 3�"~S�u�0?;� ?������&�>>-��O@-=�O(?��?�<P<LĜ>��'?Z���U����Y>�v&>N��>,��>܋�=����*E콷�?��Z?����ܤ��>Ʈ��*pm�,W=;[>��4�����I>�э<�����`���fh�a7==�]X?���>z��d����۾%.�mb�<2e�?��??�>+ف?�nD?M��<Ė�d�a��kmh=U?��m?5��=�ٍ��oо+1���<?�sV?U�=�Ė�5+��e���?�+�?jH?LB��X�������S�>?޶s?��_�rs���.���e���>#��>���>��8����>W�G?����c����F(�xΞ?/�@��?�р=O\M:?g'=1��>�n�>C�m7��1vѽ}�ؾ���=N�>��4�i��G��R��a�3?Lq�?ڽ�>�,���a��x��=W����c�?��?�m����d<[���-l�����{Q�<��=7����!����F�7���ƾ��
�~���?㽼���>U@�)��>��8�/,��IϿ\��.�Ͼ[�q�r�?�R�>�:ʽs��٠j�u�xcG�pyH�z拾>S�>�>�H��s���{��j;��"���(�>����>� T��浾/&���v.<<��>�(�>KJ�>}ׯ�'����ę?cH��CEοÞ�[��M�X?w�?pZ�?2S?�C<opw��{��&��_G?L�s?� Z?+�&��.]��8�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�d�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�@�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�`�_?'�a�m�p���-���ƽ�ۡ>��0��e\��Q����mXe���5Ay����?U^�?z�?G��� #�D6%?�>H���n8Ǿ��</��>((�>g*N>�C_��u>j���:��g	>���?�~�?{j?���������U>��}?��>`��?���=>��>��&>�(���nw<\�3>1FB>kGV����>��P?�5?|�>f��@Y*��?A�KL�r����@��Z>�Tf?�5^?T^9>��ٽ�P�����|��%��zC=�~C�Z��⽳�1>(>��*>l>�������?Mp�9�ؿ j��$p'��54?.��>�?����t�����;_?Nz�>�6� ,���%���B�`��?�G�??�?��׾�R̼�><�>�I�><�Խ����\�����7>1�B?Y��D��t�o�z�>���?
�@�ծ?ii�}L�>��Sׇ�K��^s#��/ýp�&>��0?t�
��)>��?�a���s�����9�S�T�>�+�?R��?�?
��?�#v��l�y9�g��>SN�?��?��>����w=�!?ja���Y��wAϾ/�?4�@��
@pw<?+��mpÿ�N�����D���>R�M>i5'>U�y^>�<��;�v=O�>t�>6�F>!�=V#,>�.*>ԉ>�v�O������ε���8�0�Ծ�_���̽t�оSbb��M���R����Lh����*-���Z��HQ�P|p<)�=�lU?��K?am?�h?�gQ���(>���S�=��"�j�S=�t�>A�6?�M?�Q&?W=\���ra��z��{������EG�>-*z>�	�>٤�>8��>�x���{K>�:>�Ҍ>�� >e�3=� d�g�=1*B>ey�>���>ӊ�>�C<>��>:ϴ�2��C�h��
w��̽.�?Q���E�J��1��p9��}����i�=Jb.?�{>���?п]����2H?����m)���+���>��0?�cW?�>���%�T�:>1���j��`>+ ��~l���)�1%Q>Vl?�rc>�u>�e3��6�aO��2����>G�5?4���>��u�ǽI��`޾F�J>8F�>�j����u���.���*j�?�v=�:?�;?�x�������ey����c�Q>{~X>�\'=�ȳ=$�O>8�_�9ɽ_I�(1=l��=TB[>�W?H�+>1ڎ=�>�[��V?P�H��>/mB>4,>y@?"%?et�8���e~��v�-��w>�J�>1�>�Z>#WJ���=�o�>��a>5������o�?�j�W>�$~���_�U�u��}x=-��X��=�5�=/q ���<���&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>Yn��W��F��-�u��#=~��>�8H?dN����O��>�sw
??a򾞩�� �ȿz~v�;��>��?���?��m��B���@��~�>~��?mY?�hi>�f۾�IZ���>��@?/R?�*�>4���'�>�?*ܶ?���?��'>��?�|?�#�>��j;s�2���ſ�S�wO>�8Z�A�>�[W>ڵ���/h��m�������s���T�9>�si=�Ȕ>��#�;���$>r)�i2��J%����>���>�<t�>�7?#��>�+�>��ּ)����⏾�����Y?΂�?k��<����8�>��>�R����>ŘB?g�{�I��i��>�,m?R	�?.�K?��)>8^.��圿~���
�����&>��5?[��>������=RӾ�n�Ol>=͡>� �<#ſ�o����fϽ�J�>�3?��>ޚ�=�?��"?�i�>�a�>��5������\�|%�>��>*C?�:m?Я?�v��%;�^���*񤿱�]�'�>usj?n"?w~}>hɔ��x���w�<	�#�a' =a�g?XqK?w(.;�p�>J�s?EbY?�S?��^>�DS�����<���[��>]�!?P��a�A�l[&�t��l�?�U?7��>O���	 ֽ��׼����_��8
?�*\?�8&?����2a�Jþ�0�<�!���T�
�<��C���>R�>1���)��=��>[Ӱ=	Nm�c6�Yih<G��=5��>�G�=�;7�1����<,?H�5惾6��=��r��yD���>�NL>	��P�^?5�=���{����Zp��\�T�Y�?���?�f�?����h�(=?��?'?�%�>'I��o޾[���.w�a�x�H{���>���>rNp��$�����q����G���ƽ��o����>�w�>ǡ?@e
?��>�o�>8�z��E���"���澛,~�S�$�c�,�JT�����K��P���j��B7�� ���q�>q�
�i��>~�?��N<�
O>}s�>�Iv����>-�>PǬ>�)�>��>8:	>���=�:�<�B�uLR?"�����'���込���Z3B?�qd?�2�>  i�{���k���?膒?xs�?g@v>P~h��.+�{k?�:�>���Yq
?!U:=����:�<`Q�����3�������>�C׽�:�5M��df�l
?�0?%��̾�B׽��i�C<J�u?�p?Z�.�M�X�D�}�ex�h:�����S�틾�����Q��������b}��$�M:(>d�4?�Ď?&���:���Ԭ���e��/$�Y>���>C��>R�>%�R�s=���I�jf}��,��ǐ���?3M�?r �>��H?�'7?w"U?��L?Q��>�_�>�Ҳ���
?��=<eϗ>#&�>"E?>a4?�)(?H� ?��?�3>�zŽ�� ���־�?�T$?)?��?���>ϔ�����UR�c�G=VeS�w=����=�b=o8ҽ^���Q�=B�U>Z?Հ�̪8������k>�7?W~�>���>����)���c�<�>|�
?O�>b���yzr�%c�K�>E��?�"��\=��)>N;�=<ㅼR޺�S�=������=�5���:;�mt<��=;Ք=�Ru�f��9�:V�;X�<b�>R6?��>�`>�
���5�$��
8>E�>y>�=Ž�>��B��ᔿV���o���~>��?!�?㤼��Q>3
�=�ӥ��ヾw�F��x����Z=Ǒ?��6?X�c?ʆ�?,9C?8�=?�=o=�'���m�ں��?o!,?��>�����ʾ��Љ3�ޝ?f[?�<a�,���;)��¾	�Խ˱>�[/�d/~����@D�������c��2��?꿝?�A�Q�6��x�տ���[��n�C?"�>Y�>��>Q�)�y�g�r%��1;>��>bR?�#�>t�O?�<{?��[?hT>Q�8��1���ә�73��!> @?��?��?�y? t�>i�>ܺ)���RT��<��Q�4Ⴞ		W=�	Z>s��>�(�>��>q��=� Ƚ�\����>�aa�=b�b>��>+��>��>��w>+K�<�G?"�>n\���=�W������1}@�Lu?�i�?-�*?�c=ZV��WF�E:����>\�?7�?F�*?)fS���=pͼ4���g�s�h/�>nf�>��>�(�=ʱK=�>R�>���>  ���a�8�0R���?�F?�Ѷ=eƿ��q�J0q����^�f<噒�� e�%۔�4[�5�=�����#�ɱ����[��v��P����ߵ�񻜾�z{����>i�=i|�=��=S��<�aϼ8�<1�G=��<q`=��o��q<p�7�ߴ˻�:��Y��p�_<�;I=y���d˾{�}?�"I?r�+?-�C?��y>W]>+H3����>V��1$?� V>:�N�aD���O;�ľ��" ����ؾы׾.d��؟���>��F�B�>�B3>ҩ�=���<�?�=�s=���=S+7�v�=�<�=�G�=�D�={�=��>n>p\r?H|�����D�T�����y?���>�\�;����v5?�l�>a�t��������r?��?���?�=?.�o����>�9��u5�U�>��|<#�>�
vV=_��N�>���>��,��뫿�C<�?�?='�?q�E?eˉ����������6>sb>��R��)1�ǵ[�2�b��^Y��|!?dw;�:�̾��>���=Rd߾a�ƾl�.=��5>@ub=d~��\��<�=�P|�ϧ?=�_l=�>�D>���=�=��X�=��G=J�=�3Q>M6w���6��-�%O3=M��=�b>��%>|e�>�$?'7?��e?���>�Tr�L꽾�"̾x�i>#>E �>Sb=��:>pP�>d�0?�bE?3	H?��>j̚=r��>E��>�O(��i����ذ�@q�����?y�?�Q�>�,s�=�=��V$�++9�GB��C�?��5?��?�>�����_V'�
����?�3t>ų"=�1��.|��tս�u޽_~���=46�>|@�>;�k>iY/>y��=M~>�Y�>6cR>,E=��=�E��17���ڽ�H�������������=�$�<�y�q�A= ��<b��<�����W�-P�=�X�>4i�=���>#g�=�s��a�>�:��Z�F��=�,����Z���m�"u�6y�h2+���>�8�=k?��������>��_>Y>`L�?v�l?M1>�6�c���ꄟ�w��(���Y��=�"l=涐�w�T�q?O�w�V�,f
����>��>���>�xp>K�+�vF@�@[5=��׾�3�|��>Ŝ������5��Cr�_<��M����i�%(*��E?6+�����=�9~?��G?��?DC�>b��Y�־�)>�ԉ�V��<����m�={���U?�'?ѻ�>N�E��>�������[�>���ZlN��ے�{�2��f��Ӛ����>�W���&�+"�\
������&R7��3|�UY�>��i?7�?A.�5���5S��N�3u�<��?n��?Z>*��>�w?2�m�K��/�׾��>1�?��?���?�Wy= ��=q���;�>�+	?Z��?ָ�?(�s?�{?��z�>'}�;�� >����ZK�=��>���=�)�=s?+�
?=�
?�i����	�$��U��$^�Ҏ�<�Ρ=���>�l�>K�r> ��=�g=5w�=r/\>�ٞ>��>W�d>��>�P�>�E����	��$?05>ӷ�>��?�t>�o�<�"���b�-@=-���<���گ��9Y�<��������!��7��>�ȿ��?�N?>�� �	?�����?�2�#=���>!=ֽ�)?ć�>-�e>��o>�	�>���=k,�>Z��>ߠӾ6C>����T!�^!C��R�p9Ҿty>�_��]�%��������H�<[������j��(���&=��h�<(F�?����?�k���)�9����c?2w�>��5?�{���↽MZ>���>;��>�}��\�������Ufι�?���?��b>�@�>�fr? )?T�����f,3���t�NB���9�Iw�6���s~�u���"�l?m�v?d�Q?:7$>I>iJ�?zw.�nM��0�*>$�8���R�B�<>�n ?���tW��㕾3�/�58�C�(>��M?dL�?�!T?����o[���>��K?�Y?ty�?�0:?ۼ8?aҮ��8?�[�=i��>��0?�7L?�W?��?��=�-�=��~��9A=�νK�]����<�t�?:�=��=��>���=?�=���߼��X�,ʜ=4#���
�=A�;D����=�#9<�x�=���>P�]?���>���>�@7?���Td8���;�.?�]%=\���芾D¤�H���>L�j?��?�'[?��c>=VA�"@��>��>��#>��Z>K�>�Q��B�Yk�=Pg>�>�D�=�
Y�֪����	�|̐�
�<��>l$�>�+m>|h�'{H>�gȾ���Sf�>t�6�a�ξ9��M]�!�H�\u����>�Y?�$?w�=&]߾��꽻mo�r0?�31?PYS?I�?��=�\���7�ʎ;��#6�>n��< L��k��wӧ�naS�h룽�D=�Xɾ�堾�Wb>���u޾0�n��J����~FM=A~��AV=1�t�վ4���=(!
>R����� ����ժ�x1J?��j=3v��$dU�Kq����>��>ޮ>�:���v�l�@�����8�=u��>��:>ı��� �%}G��5�<>�>KQE?uV_?�k�?�"���s�|�B�����oc���ȼ�?v�>g?5B>��=�������d�aG���>q��>���'�G��9��a.��@�$����>�;?��>��?8�R?��
?��`?*?�C?*#�>���Z����A&?4��?��=/�Խ��T�� 9�8F���>d�)?��B����>�?��?��&?�Q?�?L�>í ��C@����>�Y�>��W��b���_>��J?���>O=Y?�ԃ?��=>I�5��颾�թ�[U�=*>o�2?�5#?6�?ʯ�>4��>������=r��>�c?�0�?�o?��=�?�=2>k��>)��=���>��>�?1WO?G�s?��J?���>*��<]7��+9���Ds��O�Yӂ;<iH<d�y=����1t��G����<�;mm��DE��<�񼮿D����u��;B`�>��s>�
��[�0>K�ľ�N����@>����N��ۊ�J�:���=V��>�?l��>EY#����=ѭ�>�G�>j��f7(?��?�?|";(�b��ھ�K�K�>�B?���=��l�������u��h=��m?4�^?��W��%��/Gv?�#I?�T�D�E�c��;.��~j�֊V?d�=?�X��u>�>2��?�!�?�O?_���뇿:��o�E��fA�)T>>�>j�r�u� �O>�h?�?���0>�(��������%�>`X�?�ư?�?�V>+Q�dD��~w�5͖���l?\%�>�����C?Q���fپԂ������|X̾�����ѹ�@����7��1N���>���lڽ�~�=�F?ZCq?:�q?��]?�0���e���[�Ⓛ�J"V�!,���]���I�vk?���+�*Ra�D���Ѿ��M�e;�=��u��P��\�?LE?���;�>b�����g^ᾌ�6>\C���"�-=1ͽ//�<���=�D���1����� � ?���>6+�>o+;?�[f�7=��4��r@��4�.o">���>xz>�>�0=s�*�����4���k4�bLB�<v>u{c?9xK?N�n? =��0�ف��P�!��.��p����B>��>��>>WW��e��?&�0P>���r�5��������	��n�=�2?m�>"��>�F�?��?�}	��?���x�\�1��'�<�5�>4i?%��>��>�oϽW� �m��>%�j?��> �>1#���^1��v�H ӽ࣡>�M�>�?��2>N�P��:W��������~�%�
7>>�T?�׆��W�&�k>ҕU?،=x�<��r>W��}������+��Q�=�?x�=��>L�־�<���}���/��O)?�O?74�*��8~>x$"?ew�>'(�>	2�?X �>�rþ�'2�R�?n�^?�@J?�PA?z@�>N�=���,MȽX�&�!�,=Ċ�>��Z>�m=b^�=E���z\��k��
E=\b�=Mjμ�c���3<������K<�<��3> ��#?�����J���ྒW
�E�־�F��'�*�9�*��%p�;�f�KL��� �.�eD�Z2��Q"���T��*�??�?T�Q���¾�g��-�����TS�>����i�����O9��*�Y���<Ͼ	�'�%'U�X�b�W�K�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >_C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾y1�<��?7�-?��>Ŏr�1�ɿc���¤<���?0�@}A?��(�����V=(��>(�	?x�?>+T1�rI�����}T�>r<�?���?�|M=i�W�~�	��e?|y<��F�$�ݻ�=�=�=>G=�����J>fU�>��TA��>ܽ��4>څ>}}"�F���^��}�<�]>S�ս�;��@C�?n�����~�����������=�y*?F�?]ػ�x?(�{�
ѿ�jJ�9n?��@�d�?jN?C<�X��>���K�N?n^E?��>i#��΀�#�>'鯽Y	)���G��6>�03�;?H>>�?���\*���f�Vut=��:<[���rſ�S"�U\���=#$��#��v��Z��l����4�h�ed��(g=7��=Q�M>��>�OJ>0�Z>T�X?��m?ݠ�>~�=���!�����վt�u<�2g��F!��͋���b�������۾�)	��B��1�zs˾_,=�:�=S/R�֖��t� �}�b��F�Q�.?K�$>`�ʾ �M��.<niʾ���/����襽�5̾��1��n�b̟?�A?�r�V������մ���W?�C�P���쬾��=�_���b=$�>�@�=m��3��uS�!H0?� ?[���y���V*>���?��<XN*?�
?3�0<F�>R�%?�M'�(὜[>R�0>Oɡ>�S�>��>�˯�0��8?��T?F6����c5�>�j��}}�[�i=fM
>� 8��]Ҽ��Z>y��<�b��S��=x�����<\�Z?(S�>C%����^К���!�G�6=SV�?B�?��>y�m?�HN?@$>D��,m_����Rϼq�I?@(~?��%>�֝���A�۾e�;?�>q?́�>�|���ӾˤC����b}?��{?�W*?`c���|�G�����pv"?�Hq?t�W��٢�����-�����>!�>9��>:A�*�>'�G?���Y���D¿)c,��Ν?Q@Iv�?��%<~��;�˼>Q�>���>bO�W��s����ھ�>>��>�G���1y���$�@b����D?���?r}?���������=�ᕾ�[�??�?���[g<����l��r��<e�<*ӫ=���k"����&�7��ƾ�
�����u̿�v��>zY@"G�r,�>T8��5⿖RϿ@���]о@Rq���?�w�>��Ƚ����&�j�5Ku��G�Y�H�]���M�>��>���]���k�{��q;��.����>��m	�>�S��&��+���	W5<��>��>���>�%���潾Nř?Kc��@ο\�����ϼX?hh�?�n�?)p?��9<��v���{�����-G?�s?�Z?�b%��:]�}�7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.��*l?M�{������1�h�.��>�ހ��.��<�ԼW�j���n�K���`����D�?�@ԩ�?h�����(�n7?���>�⏾Ϋ���>V��>��>]]/>#��=�n >8���;�^�4=���?�'�?n�?�L���ީ��dd<���?M̵>[1�?g*�=�J�>{�>9�V���߽��j=S�b>���5�>o'R?�P?�+>L���M1��>�^�L�<�<aC�E~>��?�H?�4>Ź��;��;�����=��㵽�S=�R���\W=>h���>Q�=/�m>*��*fؾ��?:p�1�ؿj��Xp'��54?��>�?����t�����;_?=z�>7��+���%���B�`��?�G�?L�?��׾�T̼�> �>�I�>V�ԽO���������7>4�B?b��D��u�o���>���?
�@�ծ?li���>�ӝ�2,���ܕ��)�V�A�6:�=)7?cD�]l�=��?��3=I�t���¿y�]�r��>W��?�n�?YV ?���?�Ok�~^���Խ�Lk>�'�?�f:?�=������>]?�j˾9��D����}k?ц@@@`�[?絞��߿|���
���p����2>x��=�1�=�K���;�<< ;=߶�<�,�=3��>�O>�>:>�;B>:�R>��7>�b�����IL��H���{�����O��4o��h�~(�3f�����*�ƾ$~ٽj�ν�Z�b�J��0��n��Q�h=�J?�rT?l�O?r�?I	(=w-=��A��=��6���=P�>}�K?�PG?Q?p$���t���Y�A'��ծ�����'d�>8�}>ޡ�>8/�>E�>J��;b�=��c>�j%>e�>�t=�~���#:��D>��>EK�>��>\C<>��>Eϴ��1��F�h��
w�̽-�?����]�J��1���9��妷��h�=>b.?&|>���?п^����2H?8���d)��+���>t�0?�cW?I�>�����T�}:>=����j�@`>�+ ��l���)��%Q>ml?&�d>gpu>�3�{�7��O�֚���Q}>X=6?p����;���u���H�;�ݾϥK>l�>3��W�����~�z&i�p�r=��:?��?8���N���hv��!����T>��^>��#=�(�=�M>�`��bƽ��H��!-=���=M	^>�1?�8.>���=��>~���u�T��>$�A>M(>��??��%?�������;��h`1���t>��>؉�>$�>s�J���=�;�>�'e>����`��v���B��E[>\m��hA_�*���x�= 3��o8�=�=Տ��@�{b1=$�~?���)䈿��Jf���lD?Q+? �=i�F<��"�L ���H��4�?n�@m�?z�	�͢V�'�?�@�?���"��= }�>:׫>�ξD�L���?n�Ž]Ǣ���	� )#�\S�?��?��/�aʋ�?l�l6>�^%?
�Ӿq	�>����+��톿P�u��y#=$k�>��H?����]�J���;���
?��?���¤��ɿW�v��K�>�2�?۔?զm��;��@�@���>'��?��Y?��g>�ھ^�$�>�
A?%tR?E�>%���(�LO?���?tC�?~9I>���?��o?��>(���@3���4h��@sW=��;�~�>\�=�4¾�D��v���G��6�e��c�)�`>�3=�δ>j��d������=�x�����z�d�Xr�>�g>|@E>~��>��?<!�>>�>�:�<C���	��OĂ�
"M?��?��*��se��Ő=l�U>bVX�u<�>/�Z?e��2ᾙD ?�!O?zx?�T?w�_>U*�֣���Ჿ�Qؾue�=��O>y?�<?�Pb�c�ؽl����z�+��>��>���ˤ��7zϾ�N��Ĭ�>Ev?�j�>s`>��?&�*?l�T>�>8�I��ތ�1<M�{�?a�?�T%?+��?�,?t��T�$����ٝ��GS�Ġa>kg�?{�"?qs>v4������&<�.`?>:�=�M�?@i�?�NԼ��>&\�?J&�?q2?��>����v�!��Qc� ��>A�!?��[�A��M&���=~?�P?T��>:����ս�Pּ�������?�(\?{A&?���e,a���¾�7�<��"�ОU����;!zD���>��>�������=/>�ٰ=�Om��F6���f<�j�=\�>��=:.7��u��N*?11�= >S�ȶ>�1~�)�P���W>m֐>�u�`�l?��Ѽ=d�{7��,/��煄���?ˀ�?��?��н�>`��-?0Qr?c�3?��>�﻾L�ݾ��� 샾�&ž[��:��>��
=8{쾜�������r��+����`����>dCN>GF?R?ut�=�x�>��H�,�8�,|�j��D�e�i�$��e9�9�����S���������\ͻ��H���	�>��e��>���>ʕ
>uܤ>o�?Ny�= �>�0>{SD>!��>(=6>	Ǥ=�b�=�s��h��'/m?����F�.����ܾ�tr?��z?�i�>��> ���cO$�%A?�D�?�j�?��>|�g�k�>���>���=�x��I�*?;-C����<5�=�O���w�z�H��6��>hf>�+νS5�C�}��g��[1?�%G?�4[�|�
�;Da�����'�=�w?��?n�(� a�2񂿯/O�h4��8����V��֍��f��i��r���D��r���D'����=
,?��?� �E4꾴㫾�go���8��=Y>ފ�>�ly>��>�z >�J�5/I��Yl��~�3�Z���?�"�?���>C�I??�;?Z5O?��K?��>���>4���&��>��a;�U�>���>�W:?\�-?z�/?��?6�)?�R]>�������:�ؾZ|?�;?s�?�?F�?� ����ǽ2I����h��y�d�q�";�=��<�۽�Qf�3�T=��P>�X?���Ȭ8�����Vk>m�7?	��>v��>���(-��E�<|�>�
?	G�>E �#~r�c��V�>���?���!�=��)>���=w����Һ#Z�=������=�5��z;�$e<���=L��=dMt�0���6�:ϟ�;en�<�P	?jg8?ֈ>�aW=Q����.�&��y�=�)>M?�k��d߾qI|��Y����c��h�>���?�?������=���=�S��ϩ���!�o��x�0��?�9�>m}<?O��?�YS?��>��<TI�Γ�·j�})���>r!,?b��>�����ʾ�񨿖�3���?-[?5<a�����;)�O�¾��Խ��>�[/�O/~����BD�����������?��?⿝?uA�:�6��x�˿��\��y�C?*"�>�X�>��><�)�f�g��%�@2;>(��>8R?��>X�O?�={?�[?=�T>B�8�/�� љ��13���!>$@?ు?q�?y?n�>��>(�)�L��]��������KЂ�o9W=2Z>;��>3�>���>���=jȽ������>�EW�=J�b>e��>ϓ�>���>dvw>9z�<��F?�z�>�﷾����r����`��h?�
�?4/?�yP����bC�ne��í�>h��?wB�?��-?}_a��A�=:k��(���n�#��> ��>�(�>ϝ�=#h=��7>��>��>��]��<6�*:��R�?�%C?���=�ƿsq�"�p�������i<h!��'ie��/��N�Z���=Z�����ϩ���[�����q`��"���	��/�{����>�#�=��=Y��=�y�<Mͼ�V�<T�K=���<>r=�o���k<N8��ӻ�%��W�F�\U<�I=��"XȾ�t?aoN?�!)?�CM?�K�>�b�=dҺ�Z1�>M�=��?߇�>�=�K���� �����&���0�2|��a�s�� �(>*O��z�*>�f,>�	>��=���=�se=3=��=WH�<��=6�=%&�=��=d�>��8>=0x?�Ɉ�l?��#q��֚�v�_?25S>ܰ������v?sU�>!�{��������?���?7�?t�?��>�n��>m����l'�{�{>���x��=i����=03�>=��=ݭN�=Q��_O�/Y�?�@�!J?zt���%⿺ޏ>f;6>K�>��R��1�#�Y�Lc���X�\�!?vv;�Z\;�Q�>��=��߾0�ƾ�".=k97>�:_=c��[\���=���'?=�"g=��>��C>,U�=a��L�=5eQ=�e�=:�N>����g�4�,�;/=_��=�4b>_v%>���>��?�X0?{=d?�/�>�gn�=Ͼ(]���)�> ��=��>1Ԅ=�B>�o�>��7?>�D?I�K?㬲>G��=a�>�>`�,�ػm�dR從���T��<ˇ�?�ц?��>}�Q<�OA�͂��d>�D�Ž�h?NT1?�\?�Ş>�U�Q�࿫X&��.�����F�+=Ror�NU������j�R����=p�>;��>C�>�Qy>��9>2�N>��>�>�:�<�f�=���{��<&��Ҿ�=�p��!�<�~żLj��%O&���+�������;A�;�b]<�W�;u��=���>��=4��>7��=�ľ{p>:���1j�?�5���gE�^��K{�^�!�􁩽�w3>N%>��j��_���_
?e�>P[0>v�?~MW?@ݘ=_���#���6��k�lI$�H�;k��<�M����4�c]��i^���׾6��>���>��>J�l>b,�p$?�l�w=Y�c5���>-x��8���,�s9q�@�������i�9WϺQ�D?1F��V��=� ~?бI?e�?+��>L"��+�ؾ�A0>�L����=C�?"q�F_���?�'?��>��k�D����o��<��>���WR�Ϫ��@�^���_<��s���Q>�B���p��������X&��#Y6��L��Ǆ�>��w?��?�7����8^�C����<@?��g?s�>��?��?��U�	��Θc>9΅?���?e�?�N�=�b�=f���N�>49	?m��?��?�s?�?�md�>���;Է >�z��8��=v�>���=���=ac?�
?P�
?�Q��W�	�Z��I��^��:�<�(�=��>�Z�>�vr>-��=yg=?Y�=� \>�Ӟ>'ޏ>��d>I��>�;�>�[��:�7?�9�=��>�?�&k>#R>>0�'��_���|+<U�����K
Q�	a߽y#�=���5<ν`)̽b��>��ʿ,x�?fx=�#��G?���xc���>�+�>�=�w?!HD>��;>�`i>@ߐ>Yl�=s��>O	>t��E|8>(t��]W#��A�,fZ�Z��۲H>��}�Ie_�9���*ǽ��&�@�����j�e�J��-@�].=,a�?r��P>^�� �c��wT�>(G�>��"?��n�a򽂥�=�*�>3�>��
��~��ܙ����۾W�?5��?�l>/��>��`?���>�)�ʾ��:��8r���^��8�ǐi�	����(��1.��q�s��?�z?^�Y?x�=:�|>Vu�?FV�M¾�n>�}>�I�־w�	<��>T��������J����
�"'>��p?�?��?�z`��8���w���QX?~)a?��?�Z:?ׄh?��V��J�>�P�>h0�>�?��?��O?4��>7b�����Y-X��(��k&�)a���� ���=��#���=���=;�v������>m��="�)��F��6��
��9:�=��<WT�=7��=�!�>�Ic?�P�>S/>p�(?}ʀ��/�E���e'?�]>�ε�;���b������Ac=��x?vԳ?��`?�>�Q��s�Hv
>�NF>���=��R>mЎ>�.[�6-ý`LR>&/�=��{>:��=��ý�ɓ����_v��t�<���=�J�>�M>v	<�l�q>�YǾ����O�>����4��@��`a`�_~K���^�i�>�V?,N%?ȗ=��+�<;A����V? �+?�pK?F�?�ȸ=�q���<E���V�������>�6#>x�	������-��u�(�{+��;PC>-ع��ޠ��Zb>���m޾P�n��J���	&M=����lV=T� ־�:�o��=
>"���h� �N��Cժ�;1J? �j=cw���dU�xq��J�>��>g߮>�:�g�v���@������8�=ų�>��:>|b��:���|G��7�a��>>[E?e/_?�܄?) �� �s��/A��c ��7������r?d1�>��?��>>zF�=�α����[d�F�}0�>�g�>����7H��5������#����>��?�!>��?"S?�?�^_?��(?�?�Ð>����:ø��A&?G��?a�=��Խ-�T�� 9��F����>E�)?�B�;��>��?,�?��&?˅Q?ƶ?��>^� ��C@����>�Y�>��W�jb����_>�J?��>"=Y?Ճ?�=>�5�t颾
ש�MR�=K>j�2?�5#?�?���>��>����^�=��>�c?,�?�o?��=��?2I2>���>V_�=ђ�>A��>n?�QO?f�s?\�J?J�>t��<}-��	X��oss�.�P�闁;�JI<�y=M���It�>=�z��<纱;$D���\�]G��XD�����I�;�o�>��T>�ʋ�<W)>��¾Ա���O>���ՠ�b���N�=�o��=�4w>��?"A�>xX�j�G=�O�>� �>���Q�-?v�?s�?oPr���a��r�pr���>Yq4?�~�=.�i�w���O�w�I�=�}s?�c?�tS����r?�A?�A�Z`�B�r���>�Q���R*?��E?������>��?�a�?��>*����Z���z��=�ȿ;��>�ƾ��I��j>{?���>G[j>V�=�rf���g�-M�O��>V<m?4\�?���?�`i>�!o�������澩@��h�Y?P��>�����?� �<	����T��u���2_پ.���-#���T��y�}d��͖��p�3��=��?P�~?��}?>�W?�O���b�ېk�����~K�{<�H##�4S@�k�I�MXM��Y���ǾЅ��0c��T�=��}�[B��д?�&?0.�cu�>�����C�;��=>�d��+L���=GQ|���P=+�U=Sam�O�&�gƭ���?��>m��>��<?@G\�/�=���1�+?9�݆���"+>;�>
A�>R��>p�i�M(��ս|�ľ���ν� v>'xc?��K?�n?�h�?01��}���!�?�0�8Q����B>�:>(��>��W�V���5&��I>�H�r����v����	��8=*�2?�(�>ᯜ>�J�?��?Q�	��o���cx�o�1�艃<�4�>�i?�*�>�ц>5нd� ����>�Rp?#t�>���>ȴ����3�S�f��y۽_��>��>���>�>)�e��W[�����N兿��ؕ�=� X?�x��mzg��ڎ>��e?��E<���<Z��>O�H���0�N��<�4�=iU?�.>��:>	PϾ���d���8�pO)?�K?�钾��*�<9~>�#"?���>�/�>{0�?�'�>6qþ|�F���?�^?�AJ?�SA?-G�>�=����@Ƚ�&��,=���>�Z>�m=�z�=����r\��s��D=r�=l�μ�R��m�<s��B�J<��<��3>J�ۿ�.K�p/پ������	�2ψ�8J������
�i[���Z����v��E���$�uV���c��O����j��K�?�*�?WQ���N����q��j/����>ڹp��bt�����e���;��R��G���N!�r�O�c�h�ie�J�'?�����ǿ찡��:ܾ0! ?�A ?9�y?��6�"���8�/� >�C�<�,����뾪����ο0�����^?���>��n/��W��>٥�>9�X>�Hq>����螾1�<��?1�-?��>��r�$�ɿ]���p��<���?)�@X}A?d�(�d��MV=
��>ܑ	?8�?>QR1�]H������T�>�<�?��?�yM=��W���	��~e?�V<��F���ݻ��=�;�=�@=���u�J>�S�>҄�oRA�lAܽ{�4>م>.�"���.^��r�<;�]>3�ս\>��1Մ?�z\�Gf�u�/�HU��U>��T?A+�>"6�=%�,?�7H�}ϿX�\�F+a?�0�?s��?��(?8ۿ�ٚ>��ܾ&�M?�C6?X��>�b&�%�t�|�=�"�m������&V����=!��>O�>��,������O��B�����=��]������I�r^�eS=��l���Rʞ�'�-�RNϾ�8��+\���=��=Zx>b`@>�&<>�T�>�[?�?.��>5H�>��<Lה���Gv>߄_�][�0@���8�<堾��߾.3�9���F�x[��g��� =�v�=�6R����p� �B�b���F��.?iu$>T�ʾ1�M��-<dqʾÿ��$ք��㥽Q.̾}�1�d!n��̟?L�A?������V����3[����C�W?P�����謾��=������=#�>z��=����3��}S��t/?'S?�ع�D_���K%>����%=�.?h�?u�<ȍ�>ܿ"?\�!��q꽑![>+�7>lJ�>���>��=�%���;�j�"?VuS?����ߜ�%��>,¾/�x�}n@=�>�00�L�+��.W>c��:���f��;)�9�7��<�f?�2�>�(3�_��f�[����=W�H>M�?�'?��r>�e?���?�j�>w��0���#�6�K�&�!?O��?�2>��������Ѿ�<?�J�?}�=봪��y�Dl����v�=?ԑi?�H.?�Ir<j*��0P���-!��SP?��v?s^�xs�����P�V�e=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�%Þ?��@���?K�;<��<��=�;?j\�>��O��>ƾ�z�������q=�"�>����ev�����Q,�f�8?ݠ�?���>��������=�ڕ�tZ�?��?N����Og<3���l�0o���D�<-ʫ=��7M"������7���ƾ��
�����ۿ���>@Z@�H��)�>�F8��5�\TϿ����[о�Xq���?�~�>2�Ƚ�����j�wLu�S�G���H�ߣ��G�>�>�:�������{���;�V���K��>�M	�YK�>�S�w<�������K.<���>,�>�Ά>宽�½��Ǚ?&M��<οF���8���X?�T�?^��?��?�<@<L�v�9�z�j��DG?�Ys?�Z?�(&���\�b7�3�j?X_��U`���4�=HE��U>�"3?�B�>�-�خ|=>[��>h>�#/�x�Ŀ�ٶ�����&��?��?�o����>S��?4s+?�i��7��\����*��q+��<A?+2>B���<�!��/=��ђ�y�
?=~0?�{�v.�U�i?T�������4�n��=p��>�Ș�1�O��;n��,�=)f[��������๮?��@�æ?�Z�13�$t?���>�+������r=>�Nx>_G�=���>A'W=l�>I[=����p�=@}�?de@�{*?"L��㼨�3�O>���?���>�-�?�\&>���>e��=�ʯ����<��M>�+%>;zu����>	�A? ^�>���=��/�۔ �_68��V��V�T�G���K>E�v?*	I?��{>Ӑ���1[�b�$�����o�79�;���i�=(}��R	>71�=�B=>MŽ�`����?Lp�9�ؿ j�� p'��54?.��>�?����t�����;_?Qz�>�6� ,���%���B�_��?�G�?>�?��׾�R̼�>;�>�I�>J�Խ����[�����7>0�B?]��D��s�o�{�>���?
�@�ծ?ji�+q�>9Hվ�����恿�10���w���Y=�}O?������>p�"?k> ��m����g��2�>L�?m��?���> i�?@�����p��fǽ7��>ۚ?�9?��HE:���x><�?$*3��׈����R��?�$@�J@��\?5�����ڿw�������v��Fa�;4{>�KW>�D�ώx=���ぽä��.L{=�Ȇ>�aY>�φ>&+�>8HN>?>�<���i"��y���\���JZ����z��#a���}���թ�+6ȾrU¾%琽��b�11�X��_���A���#�=/�M?�\?��a?4Y?#㎽b�!>�Mپs�?=�W�wU�='݆> W9?S1<?�n!?�(M=<�����c��F��Q������|�>���>`�>���>�ύ>f�ּix>}�>. �>���=�\J=�g=@�~=�A>��> '�>C�>�C<>Α>Cϴ��1��[�h��
w�̽/�?h���N�J��1���9�������h�=Eb.?|>���?пe����2H?���n)�ܹ+���>g�0?�cW?5�>)��V�T�6:>M��Ŧj�$`>�+ �?l���)��%Q>fl?��q>���>T�,��4��4I�Y�����}>�>?o٣�S�0���l�5�A�60Ӿ.�<>в�>�$&<��� ����r��GՀ��<=-C?� ?rdƽD���'�v�G�����K>q"X>{n=�=�qc>��6
��CV���=N�%>��i>��?�].>!�=	[�>C>��F�S�4Щ>y<@>�X&>H�??(�$?l!�́���Ճ�t/��u>���>ƽ>��>�6J�S׬=W��>�d>~���⃽�"E�p�S>�A���U_��Jy��Uz=�n��jD�=uc�=˲ �y�<���.=�'�?�0���N��Ce�O�(���$?�L?�+�<>\t��'�ô�������?��@�X�?O��K�~�B?]��?/���>k>���>[|>��7�虓�dd%?�;ɽ&_���>��EL��"�?4	�?�~̼D0����X�)�A>dB?�����x�>'`�?Y�������u�p$=:��>9H?j6��d2P�s�=���
?|?b�>�����ȿB�v�b��>a�?��?��m��=��v@����>M��?TTY?r<i>S۾b�Z���>�@?�R?s-�>-�[�'���?&Ӷ?߬�?EzH>܂�?�s?��>рz���/�8Գ�����=s=%��;=X�>4J>LR���[F�aϓ�H��l?j�d���~b>�&=5��>�z�(��'r�=c���Nx���_j�W�>Q�p>qvI>�Q�>�� ?���>��>k}=5���N���~s���L?�d�?�/	�|8v����=�d)>�o�;��)?Z>?=�|��Q����>�jC?'-L?M�L?p_�>#)(�퐻�g¿��ʾa'=�i�>`�?�-�>}��;Y=46]�	d��p�{>]��>�b*��������=Pt�>ʕ?�o�>�S�7 ?��'?#M>��>$�W�������l8�>5�>�}<?X�o?�?`���C�qJ��ʙ����1�1�{>�n?,�7?�"�>�-��������=��$>�5�G�?P�?�NսQ?�k�?��m?|�?���=��G%�P6A����>ä!?ʔ�v�A�V1&�T���U?�H?+G�>�@���!ؽfOؼn��/�����?7\?��%?���E�`��	þ���<�o'�}�^���;نD�n�>C>ܸ��0'�=��>DR�=��l��z5��d<�?�=�p�>���=��6��ʎ��$$?�E#=�n��J�=X�o��M�Uhn>�k>��˾ܻc?8>��[v�D��ب���;y� ^�?�:�?���?�ỽ4d�#1?&��?�0)?�s�>�t���^¾s.�!����n_�v��OM�=��>61�<�o̾O���y��,����m�!_"�D?�9�>k�)?3��>��	=��>�G��/�N��D־/M�Gk�(���$�|�!�����ˊ��)��<�i����{��I�>Ed���z�>8�>��v>?">�0�>�*M<,�>�%c>��e>��~>g�=J>�#�=�wY<ˏ½n�c?	����+�����J(��*7?�/�?�L�>QOX��~�B�0�WU�>+]�?�=�?Յ�>Q�P��`�i�>�?뛾٩0?��S>��<"�W�l����i=�cf=b�=h��>>0t�gi4�"�y�
���$
�>�h?ʙ�<	y�=�c���{G�=,�?* ,?��>�`?T�V�g�G�I�g"�<�=���h�f�7�/�k�ؿ���pm� �s�(�/�=&i7?�}?�4 ����Q�ؾ�{�R�T�ݪ>��?�`�>��>�Q�>f� �Ua5���c�s)�ą��b�>]߆?aH�>��G?��??��H?�I?}��>�>�����Q�>]��ö�>�P�>��<?�&?y�)?��?�&?JB>"��� �޾x�?��?�j?� ?���>Fg�����s�S��nt���j��v$�5��=#�<X���~J���=i�W>�?w��Z�:�e���zMr>�G;?���>��>�r���؊���%=3:�>�?�{�>uf�ָv�����v�>ix�?����[�<'$>���=߼p����<+�=��6�ܥ=��üܤW���<�W;�=���=\�<<��L':�LF�{�d<���>�+9?S=�>;
z>����A'�0��]5>�-J>6��>��>Fc޾����w]���y�� >�1�?���?#����j�=�	T=�݁�Ҟ̽������:�.>=n?�y�>��W?�0�?��0?�k?�>��㾐{��`䍿�Uľ,t'?�,?�>-��|�ʾਿ�3�ߕ?�x?�	a�����$)��z¾!�Խ~></���}����R4D�𤚻���[ϙ����?G��?نA�l�6�Kh辦���RE��{C?�,�>C�>�4�>X�)��g��(���;>���>�R?v	�>��O?pB{?-�[?�qT>n�8��.���Ι��4�">w@?���?��?�y?0[�>��><�)����P��/��W��?Ⴞ>�U=�Y>���>�+�>{̩>&��=5EȽXv���>��A�=��b>�l�>��>���>�nw>�Q�<x0??��>�޸�7��n
��4N��<��65^?懑?�?�ļa��HpJ�g����>4ܮ?��?�/?�煾��=K�7�o��!Y��ܬ>��>v��>�$�==�=��&>p-�>���>�����J�W�C�)Ħ��1 ?�FC?��f=+Fп_^J�����P�վ����E�e�P�0F�*V��ʓ=W����T������g+��Ƙ�������x���H��'p�>�Wv=pg*>&h0>>�f=���;ָ�=����#�=�2u>Ebf=�ט�������s9�#��=8G�=�"E<Ϭ½9!��g79?��k?�(E?y5?0�7>�`K��Q���*>���;�3%?�/^>�`>^C��q�	��NȾ~�{�(�վ N���A��5��%��=�i��Ĥ=�<>���=8'���8=H"=|~'=�/\=�;���=�O=^3d=� H=���=�N:>O�o?�鏿�����|l��u���zi?�h�=������n?&��>�v���s�����I�v?A��?sW�?�U�>@������>����
�:�=}�a>᩠>�۽O�����>��>m�H��թ��}>f��?�K	@;G?��m߿~C�=K��=B>�|g�Z`���F=�<s�Ȋ�<?J#W�Vs���lB>��X�D��]�f����="�=Y���٥��E�p� 8� ��<�P��Ao>��F>��Z=�������=y�z>�s>	ʁ>�7
>ƛ���Z�<��<XRU=�j>�>E*�>�!?GI0?uzd?e��>U`p��Wξ`c¾#܊>7��=鮰>�=�#@>��>�>7?J�D?��K?�R�>۸�=�t�>���>�,�4�m�{�徨ȧ�7�<Ñ�?�?=�>KPX<F�?��!�~b>��ǽ�??�1?[x?)>�>�j�&	�k" ��#�8�D�gş=v��=ɕ[�PI���rL��`l�2�1�dy�=8��>���>��>��>5y8>�%>5��>�7>b��=���<�.���H=�@�<.�=��&=�s<��̗���{=�}�=�f�kE=X$��vP�P� �<y	�=�@�>�I>{>�>��v=T�ƾf�+>̼��	&R�	��=�Y����D��c�hG|�;�/�5>:� U>�wU>��q�N׎����>q�a>1�p>4�?rIn?,M1><�?�0J侽ؚ�V�i�0'm����=G�>ou3�OD:�Q�d��hP��ɾ�n��>}��>B�>8�l>�,��#?��w=��c5�G�>|�����+��9q��?������9i��pҺ��D?CF�����="~?j�I?��?k��>r����ؾ)70>HI����=��Y)q��d��^�?F'?}��>��i�D�Ŀݾ���:�`�>��l��I���8��;>�^dt�|L�>Y�.�����]�=�����y��|�8�4c�
��>loQ?���?�-S��j����f�i�*��b��>��{?�#�>5'�>��>o�����߾�tþ�yV=�oa?C�?}��?:�;>�r�=���>��>�	?�?ޫ�?�ts?�+?��=�>y�;;� >&�����=�>3��=���=�[?�
?�
?�b����	�b�����^�k��<��=��>As�>��r>�=��g=�Ϣ=O\>�ƞ>�ۏ>|�d>�	�>�P�>]����l���>	}�<*��>z/%?�@�>�Ht>�26��7x������v�/�lf�=M{^�*sW����?8>����&�>�Ⱦ�3N�?9�n>�"���?��ƾ�Ю�ڊ�>*r�=5�����>!�6>�T�>�{�>)��>+$�=�'�>($&>dվw�>M'��� ���D��sS�4վGQz>������������!�M��z��ޱ��i��み�X=���<�x�?����pl�;�+��U�B;?'��>�[7?X?��"t����>u�>*ˋ>K=��HD��{����Q޾�E�?���?G15>��>��B?��>.~ͽ�%��Z3z������9��h�ٻt�T$�������(��<��?Nr?;�K?�B<PGH>ww�?�0�־���>�?�%�L�H)����>�3����.�վ���
䵾D8�<~�?+7�?k��>�ԗ�Z�ʽ�&��
�?�TM?�5?���>��>�����>6p�>GC*?+-?6?��>��>>B��H�����+�����}�� @����j�:�7��6�<r��=���ǈ=��>95H=���=��	��D!<�k`<�]p=�K=��>�^�=���>	�?Et�>�E7�N^??��־�b�Z�農R?<;������ ���
h�fW�?���?�q?j���`	��K⽉}>i�>��=���=�>h
�= qʼ�>J>�Å>��>>1�=$cD��Gﾥ+��hx<�j�=�,�=��>�X>��@�"X�=������s���>�)��_P�J�����[���?�;����>�Qd?K�>o�9�"��������Y�E?W�>t�F?[a�?�PD��.������<��\��X�>�QݽZ�>�-�����./��н1i�>Yܮ�!+���q[>
�#H۾�o��M�.��>=,=ϳ���Q=�'��IѾVt~��m�=�w>[7¾P� ���NJ���I?�n�=�}���&W��$���`>\��>ب>Y;��Pd��.@�����V�=�,�>
�.>�^�o[��F��1�Ɇ>��G?�-^?車?����Yo�)�D����¡�� ���`?ъ�>��	?aB>���=LU�����?�f���G��n�>b��>�t�aED�mo�������!�g��>��?�45>��	?b
Q?O�?�\a?��.?�D?Mڍ>,s���y���%?�i�?��=����!R�7��6�A=�>�F#?�"��E�>H?��?
�'?��R?2:?<��=�� ���;�~#�>lՈ>�Q�߭�aqR>�lE?� �>p ]?_}�?��I>�2�����5=ͽ�{^=�|>z4?#"?�}?��>���>F��g�=]�>�Gc?��?S�o?�q�=�P?oG1>���>Ɍ�=У�>V<�>�C?�O?�es?��J?��>�\�<l��fR����s���Q�w)~;�[F<�%v=O+�D�n����`��<��;qP���{�:����A�"�����;�b�>�t>�����1>��ľhT��pA>�u��YR���Ŋ�"n:�w��=��>?���>U#��=��>"?�>����0(?!�?n?m�;h�b���ھ:lK�A)�>�B?J��=��l�䀔���u� �g=��m?��^?SkW�����b?/�]?�g��=���þ�b�K�龎�O? �
?a�G�5�>}�~?|�q?��>��e�!:n���1Db��j��ж=)r�>1X���d�h?�>�7?�N�>2�b>c%�=�s۾��w�kq���?��?H�?���?�**>I�n�4࿀�ʾGꖿ�l?yn�>�$�= Z?���=��*$��A ھN�J�H|ܾR����=/���<��6���
���>��?.�/?Y\Z?����?S��<��L��>�W���!��~4�M�S��F�QD���W�d%*��!�Tbþ$�"�nqb�}�V�j��?+$?�7v��K?�Ƌ�_vɾ􌾑�>�JB�� %���<M�<B��<���=Ϗ,���r���/?�ʶ>,�>�H?'�j��<A�C~D��ʾ�>2��>Y$a>/��>�@==��W��/�5�о�7��l���1t>�Yi?Z4H?+�e?</�^*�.���W.�)�8�&�����T>��>���>�<8��`���r'���>���w�ǹ�����F����7=�p2?O��>���>zR�?6?�� ��o������x*�A�*=56�>� w?� �>�vs>������d��>��l?���>~�>0���8Z!�0�{�m�ʽ &�> ߭>*��>B�o>˫,��#\��j��P����9�lr�=t�h?΃��a�`�>�>�R?�`�:.�G<�|�>��v��!�p���'�3�>�|?���=̞;>�ž�$�W�{��7��'T)?k�?Db���)�Ŗ}>�n!?ji�>���>I�?u��>ݐ��r�8�b?o}^?��J?��@?S��>3T=�-����ƽD�%�q.=ؑ�>�rZ>c"l=�=�W���W��m!��B=��=jcԼ���<&��;�f<�=+�3>�㿓�U�xվ.���̻���-�*�l�p<׽S*��i����߾��a������岩�$=���@�m���!ڕ�G��?zx�?q�����L��G��'xv�X��B5>U��eՌ��ľ���t���⾋b�@m-���a�; ��|�{�L�'?�����ǿ�����:ܾ6! ?�A ?=�y?��'�"���8�Q� >�D�<90��Ν뾧����ο����^?���>��#0��B��>㥂>H�X>�Hq>����螾�0�<��??�-?��>��r�'�ɿX���FĤ<���?(�@�zA?V�(�����-V=���>ԗ	?��?>�C1��?����i_�>�8�?���?B�M=I�W�x�	�Pe?��<��F�l�ܻ� �=)�=��=[��N�J>�^�>����?A��Fܽ��4>�Ѕ>��"�ל���^�^�<�x]>m�ս�H��5Մ?,{\��f���/��T��U>��T?�*�>N:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�ޅ�=m6���{���&V�{��=Z��>c�>��,������O��I��U��=���8uǿ�=+�����K7�����ʼbE��߽Q�N��괾��>����Mא=��>F�[>���>H�n>��`>�U?g�n?m�>>���;�����۾����w�ɐ7�\A����1��ξ\��X���@H���)���ﾴ!=���=N6R�	���� ���b�>�F���.?�t$>��ʾ�M�ڰ-<�pʾ]����愼�㥽r-̾�1��"n�͟?��A?6�����V�����V�h���D�W?�O�����ꬾ}��=Z�����=�#�>ņ�=���v 3�~S��u0?b_?�t��FO���%*>!� ��=��+?9�?B�[<C/�>�I%?��*���g�[>S�3>�ˣ>V��>�6	>c��N۽Ԇ?9T?p������tސ>�N����z�ͧ`=_+>�45��,�݄[>q�<N쌾��T�����}�<�(W?q��>��)��qa�����Y==��x?��?%.�>k{k?��B?դ<'h���S����aw=�W?/*i?��>����	о^���G�5?�e?��N>�bh���>�.�[U��$?�n?4_?[~��'w}����n���n6?��u?�K����`�!���<���>璋>���>t���?w��>��̾�|��"zȿTqS��ļ?`@i;�?�4�=�J����:>YI?�p?w*;;0�\=/��c.��g ?0�O���`�c���XD?Q:�?I�"?S}�5��m�=�6y�uy�?t;�?Į׾�'>e��k�i��B¾�%��a��<� v�@c^�3����1�%��_������&l���W>#�@�iJ���>Y��<0�Οտ��r���������>���>;D�<����d��j�	�O��P��M_��M�>�>���0���-�{�|q;��!����>M��	�>��S��&��������5<��>���>p��>�*���罾(ř?�c���?ο.������n�X?;h�?�n�?-q?�9<��v��{�z��.G?��s?GZ?wp%��=]�c�7��j?`��V`�h�4�<GE��U>="3?�C�>��-���|=K>*��>=e>�#/�m�Ŀٶ��������?Չ�?�n����>D��?t+?�h��7��\����*��h-�=A?�2>������!�0=�dҒ���
?�0?�z��.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?X#�>l�?1��=tt�>���=�۰�0�*���">�J�=�=�M�?Y�M?X�>�p�=O�7�F!/��`F�rGR�i���C�R��>�a?�yL?�&b>!Z����0�� �6�ͽP�1��A�%@���.��޽��4>=�=>.�>p�D���ҾI?�;'��`��-���۩���H?ȕ>-G ?��B
�Q&?��i?�*`>Ll.��ɵ���f�.�P���?�� @��?�Ⱦ쐽jc�>g�?�͎>#�0�+_ؽ����>��=�-%?�}�X���y���^{>��?7S@J�?xn���?7q���{���پ����e�=�<;?{s�����>���>X��=�qt��I���)x����>�ݭ?&��?�+?��g?� a�J�4�M��=��>�Y?���>a��w���38l>
��>d!�3�H�
�WWX?��
@zg@�@T?;u��+ÿ�I��f���lGW��b����%��>!��<�؝=���=e�=M�=��m>Tt�>sI�>g�/>�->	?e>m�:>��}����c��������h:���1��	�<�P��X,�{����<YS��햾(���V}I� ������P���U�<�L>�_j?�0?�]?���>{�8kW>������|k�=���>�ƥ>Ni5?�~l?e_?����ѹ��c�mmI�i#�`�y�>�Z6>l��>�̅>��?_��>$�>�D�=#c<>p�k=�9��g���4���.b>�Z�>�w�>���>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?!�f>u>H�3��d8�K�P�x|���h|>I36?;鶾�F9���u���H��cݾ�HM>1ľ>�'D�l�u�����kui���{=x:?h�?�3��t㰾]�u�aC���PR>l:\>�T=�k�=FYM>hc���ƽ�H��d.=̻�=��^>!�?2^/>3�=!;�>�;����P�{�>�nC>C�,>�,@?aK%?a$�D����X��p�(��Yw>���>8�>p�>9�H�Nΰ=J��>�l_>�p��Ƃ��

�u1:�)=]>����?�_�Ӌx�&,p=a�����=�W�=n��_9���&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>��3������痿0�e�Dmu=;#�>�O?2���`�<��v���?�
?qp�e���쵿),��/�?B�?z �?�i`��)����x�w�>��?��;?*E�>��۾� ;�D��>Ƶ[?��V?�C>�d(�в��?���?s��?�D0>er�?�8Q?R߶>��H�����������=c�оZ��>!Ӈ=v��zN ��⋿\����_�xK@�`)��Ґ�=F��>_^ƽ*i���ܽ�d�Ԕ����w�AD[>��?`i�>�Y�>�zK??|~>�>�K�=�b��s~�̱��
�K?޳�?����n�#�<8z�=e�^��?�>4?�eW���Ͼ9֨>Ҿ\?/À?�
[?�Q�>���<��⿿�p���@�<j�K>+�>�N�>��{�K>�Ծ�)D��m�>iҗ>�R���Fھ+2������B�>�^!?I��>��=ڙ ?��#?��j>�(�>CaE��9��X�E����>آ�>�H?�~?��?�Թ��Z3�����桿��[�o;N>��x?V?tʕ>b���񃝿UkE�KBI�F���]��?�tg?lS�0?<2�?�??^�A?x)f>؇�(ؾp�����>��!?�l�'�A��"&���_?�u?���>bޒ���ԽC�Ҽ���[��a�?�2\?�3&?���la��¾���<�!�n4P��"�;{xD�X�>��>o��^N�=r�>;s�=�]m��z6��Z<IJ�= ��>qk�=0�6��I���S%?�����N�����7�W��;��z�=e�\>P��[�}?���}���ԯ��g��J���Ԥ?��?��?�=�\�k�!?�?�?��?3��>���i.��9�� z>�᪾0���Lq>�RE>:�>��z���C���ns���?���5����>��>�K�>uw)?[2V>�#1>@�E��
�{a�����)>Z���4�]i<�}&;��_���!�6�ɽ�>��<þ�����>�����C�>��?z��>R�>SO�>�o�T��>��>���>�Ţ>(��>/�C>cy�=�3;ҹ׽�KR?�����'�W�辨���a3B?�qd?J1�>�i�4��������?���?Ts�?G=v>�~h��,+�qn?�>�><��Qq
?�T:=�9��9�<V��4��3��;�@��>�D׽� :��M�Onf�jj
?�/?2����̾�;׽�����s=�&�?�f'?�D*�||T�2k���Y�S�O��'ͽ���=̢��%�4�a�ʌ���������,�>�ﻄn'?�e�?�J���r���ˑ�w�f�(tB��[>���>!֜>��>�BE>L�����3��a�Q�#����>��y?3�>|bI?��;?�hP?�IL?�+�>�˪>1��s`�>nX�;��>�^�>��9?�1.?�0?��?�o*?��`>���5��� �׾x�?s?��?�?�?T̈́�oĽ	�����`���y�%i��R�=Z��<u�ֽn[q��Y=dT>�X?����8�����k>_�7?o��>���>[���+��P8�<��>.�
?LI�>]����}r�ec�cS�>١�?����=��)>3��=����WwӺ,]�=��� �=�Q��l~;��<�}�=��=0�t��������:۴�;or�<�n�>�?>�5�>�7��O� ����y��=�Y>�BS>��>�]پ����&%����g�ay>�x�?�v�?مf=@��=�y�=l��tQ�����彾���<ţ?NV#?�JT?Δ�?��=?�a#?Y�>�0��S���^�������?w!,?��>�����ʾ��։3�۝?i[?�<a����;)�ߐ¾��Խұ>�[/�i/~����>D��텻���V��6��?�?KA�W�6��x�ۿ���[��{�C?"�>Y�>��>U�)�~�g�s%��1;>���>lR?n��>�1d?�ke?t�F?8a�=�F%��ɧ�qL��̼ۜ�`> $<?i�m?a��?d$z?ml�>Z�<����E�8	�<q׼������)>X��>�ED>�?��>q��=v�=�<̽�#�6Ź=�o�>^6?vt�>�>�m�>�0r=�G?���>QX������ꤾ�Ń�.�<��u?㚐?K�+?�j=����E�=D���L�>�m�?���?�1*?I�S�k��=��ּR߶�r�q�1%�>[ڹ>�3�>�ޓ=��F=ZV>�
�>ٞ�>4,��b��o8��QM���?DF?饻=#Pɿԑm��{W�#0��"�(��;þ!�n���꽜���=�=����\׽䚥��wU�`�������3���&�������B  ?C>R�->z�=8�5=������A�?b�F�X<�9k=ˬ�H얼wsD��{����g_���z�A.1=�K���ʾ�}?H-I?f�+?�sC?ܐx>T�>�=,�xd�>�[��p"?;V>GN� :��?n9�HZ��> ���iؾ�׾��c�2���z�>�&H�u>�42>�S�=F<�{�={|n=���=�]'�_f=��=c�=��=��=82>��>]"w?�8��꧝��QQ���彠�:?_�>=��=�ʾ�lA?�
6>�ф��n��,��BX}?���?���?L�?k�e��)�>ᠾԄ���=]q����,>u��=��2��p�>4�J>9{�����<A��r�?�t@vB??㌋�_�Ͽ,�1>�<7>m�>F�R��1�b�Z�s/b�+H[���!?�;���˾�ͅ>ع='�߾a�ƾ��*=�*6>��e=����a\��B�= m}��]==k=n͉>PcD>�O�=�x��Mض=�E=��=�tP>�Dw�07�l�'��5=���=;~b>�%>$�>�Z?kQ/?Fc?j~�>�u��}���ʸ����>�>�m�>#U�=gyG>��>�<:?Y??g"A?W��>W�{=C�>	h�>�X&�r�k��H⾽���&Uz=��?��?��>�&;SU�ck���E�Lý��?��/?>�
?���>g��A�[�2��u$�U|�����<D�=��Y��ʽJy�ِ5�:nn��>�ܬ>�>�>��>ꥅ>�[>P�n>.+�>�> �=K(=?�1�94Ҽ��<��=�(��щB�%����޼�o��6cV�3�����<���<�e�����y��=_#�>= #>�3�>5�>xh����8=��o�S8��z>tþi�K�?�q��&��g8�4�<��6�>@�^>�eZ��E��>Ne>go>��?��z?y�
>��F���̜��w+�����X�=\�,>2rb�=�J�տ\�v9D�m��`��>Rߎ> �>|�l>�,�L#?�,�w=��Zb5�}�>�|����D)��9q�&@�� ���ni��`Һ�D?�F��p��=o"~?��I?b�?��>;��Ԇؾ=;0>�H����=f�|*q��h����?'? ��>�쾪�D�P�̾�N��t��>��I���O�x��� �0�!%��������>eI��;�о3�!d��������B�;s�%��>�O?���?�%b��|���O����㈂�#Z?��g?�@�>nR?\?Tu����쾨���&�=��n?��?�X�?Dy>�F�=w+���6�>z�?O̖?��?QCs?,�>�>t�>�Α;�K >�����=�C>I��=���=h�?�
?ו
?`���,�	�h��o��:0^���<��=��>a�>@�q>}��=�h=���=�\>�1�>�>��d>��>pQ�>����2��=F?.��
�>�)3?���=j_�>xǞ=joн�f��f�~ԉ�*����Խ��>_]>m��=;�ͽ)}�>�ſɱ�?��>qfQ�w�.?���7���1�>zL��Ҋl>7��>|`�>�I?C;�>�]�>��G<y�>���>���f��=�t߾	z�%7?�(ap��{�����=�j����ν��*�v�\][�-Ը����=/f��܂�qR%�]�;��?��������\q�����6?�f�>)�`?����=��d>��>�ٸ>!'�;��u�g�iS��F,�?T�@):c>�>��W?^�?��1��3��uZ�Ѯu�Z'A�)
e��`��፿*�����
�i��j�_?��x?�vA?Y8�<E9z>��?��%��ӏ��+�>< /��(;�=<=�)�>
)��<�`�`�Ӿ
�þK;�[CF>��o?Y$�?�W?�RV��0�>���>0\?
^A?�2i?��>^U�?b.�>>�V?c��<'�?<o,?N?��+? A?!,'>a�������/=�뼩����w��ꪺ�Z�=���=۱*���ܼjj:����ƚ�<��S=AZ�=� >��ü����ѥ=�H�=�2�=�g�>�\?���>���>=�8?����)9�~�����.?,�B=�샾������U���c�=��i?��?��Y?�)_>��B�2E��
>��>�()>{L_>�²>�B�D�y�x=�>�J>9�=p�G� ���:	�C+����<g<>���>�0|>^��-�'>�|���0z���d>�Q�'̺�B�S�v�G��1��v��Y�>��K?W�?@��=b_��-��6If�?0)?�]<?wNM?��?G�=�۾H�9�n�J��>���>�a�<��������#����:����:��s>&2���0;��p> ������K�g���Y��b��O��h��^���F��L����o��>���=�����!8�͵��ϰ��HQ?�(�=�K���j��_��G4�=�No>���>�?`��l���@��N����v�hU�>��=�3�d{��5�w��x=�>�WM?_<\?�:�?�銾Q�|���>��^�֫�����q�
?�`�>�{?��P>5@�=��;}��Lo�%}O����>���>}?�n�N��f���cȾb��Dx�>
�?UG�=��?t\P?j�?�S?�%?%�?0i�>�bx�����?9��?2>{	μ��+��5&�V�����>�?زY�I>��?�?��?�fK?�8	?��~=N��L�)���>��Z>p][�&"��c�>��Q?�t�>��Y?Z�W?�n�B�P��ӆ�eeF�	��=����k�>DX?ճH?�7�>��?�ֆ���=;�>�!?��?3�w?�ƃ>q3?�<�>]�?g�>�>�+?��8?"DO?F1?�B?��>Q�=�Z�<VV�[-�,����<�>��	=R�o�!��Uc<��(<�`�P�<~x�=�8���Z��<WS�<�g�>-W>�l��4Bh>�Iھ%ʖ��;d>�<s�������e½V��=�^�>@�?q�>e��+��=��>�>�u���?�u�>�?k=��� W�J�Ѿ�.T�`2�>�'V?��=ZZv�q����f�7{�=:Ct?��P?}�y����O�b?��]?=h��=��þz�b����e�O?;�
?;�G���>��~?e�q?U��>��e�(:n�(���Cb���j�'Ѷ=Yr�>JX�P�d��?�>m�7?�N�>-�b>%�=ku۾�w��q��g?��?�?���?+*>��n�X4����aߚ��{o?���>j��jD?��;�1��K��}:��;[��Ⱦ�����i_�퀼��Y����Xɫ��P>k	?�)�?�V?��q?v���p�R�N�Y.t��,L�p����"�\[�^�C�MS�XHc��,3�����˾�r@<Ҕ���O���?��?3b�E��>�~���B�s�����=�����ӽ��x=��<	�o�=�|"�����ݗ�� ?㭿>Z0�>�UD?ank�[�I���!��,�
��9[>�t>Y�>N~�>�>f<��J�n�J�F�;�ت�$2���E>�.�?)'7?g�n?�*�rs]��r���_��N�
=]��.V	>�򱽋��>�ZʾkJ�3?�o�?�6q��8�+�������.~
>�,"?�;Ro��"�?�'�>�xJ����������(��$>;7?���?��>[{=�C�s�.�ĕ�>��n?�U�>�#�>��u��"#�����B�3�9�>-��>yr??/W>Z����b�����z]��"I3�^v=9�]?F����.C��>U{N?�3�Y��;-�>�^ν�f.�����������=^?���=�>�$;�
���w��ء���'?5D�>K(�V�˾��<tf)?�?�9�>�=|?�H�>���~p=�� ?U�R?6�D?H�6?���>"%l=���wϽ��T��}�<�P/=��>i�*<��7��l��A�V�Zj��sc=���=[Nj=�h�纖�1{:m�d=^��<���=7�ݿ��=���������̾�;�\%�E�:�{V�z)��	A���D�����4oz���$�����WF��c���]��?Я�?V������[����ꁿ����E�=@�e8����������r�B�پ% о����yS�4N_�I�s��S"?F(��hҿT,���,����$?�v	?��?g���#�L�M��t%>�˯=X{�8w�'┿�ֿEZ��I�?�P?����&�"�>�>��^>7T^>l?��͟����<�T?�jN?���>���OsĿ	`���A<[��?��
@�lA?��(��-��W=f��>͂	?: @>f�0�{>�})��l`�>� �?��?��O={�W�O����e?�V<�F��ػ���=o�=�=^���I>�Y�>���KA��ڽ}w4>�]�>�#��a�h^���<C`]>}�ֽ�ڔ�(Մ?�z\��f��/�%U���T>��T?�*�>�7�=T�,?�5H�=}Ͽ��\��*a?q0�?���?��(?oڿ�.ؚ>;�ܾՉM?#D6?���>�d&���t���=�#� E��u�㾝&V����=���>J�>W�,�@��ևO��a�����=���mƿ�L$����<��^���_��X꽦e��ƨT��X���o�U���j=8��=O�N>�+�>�ET>��W>�W?l?h��>58>�]��w��X�ξVYs�����q�;���f
�.���+9�!=߾����%�2
˾=����=KR�ʂ���!�%�b��oF�y�.?�$>5gʾ_�M���<��ʾ���� �������I̾Q�1��	n�g��?��A?�܅���V�����4��ѹ�}oW?ݳ����Nج�(�=���4=-A�>oʢ=���(3�8qS�71?,�?�����hz���,>�ýr��=��$?j��>����{Ũ>LU?4�����ڻ}>2� >>��>c��>@0>�Ҩ�&�Խ�?eL?���S���6��>�K������x�˻sO>�Y8�p���?�>�E�<C?|������*��y�<,W?�F�>}�)���M����h#�ޮB=�Nx?��?��>Īk?~B?���<������R�p���x=��W?�Ui?~	>����0Ͼ�b��Y�4?We?�O>�i�����Q0�B���?s�n?P?嚼�|�݊��5��zr6?wq?��;��n����/�o��<�a>��y>ԫ/?{�{��^R>��(?T�U��r��U6���0S��q�?ݙ@�� @�}�=������]>��#?�y�>�_��h�G��=�=��??S�S<�>�^�z�c�@BS��<���f&?�'r?�?�˒��r����= H��k�?̴�?X���4
۽xR�7L;�G��%4ɼ���ܫ�KL)�s  ��fJ����6u���{��Tn�=�Q>	@|`���	�>��>��)ѿ@ؿkY��3�$����d�>�0�>ug1��23�-����́�,~��8a�ᕉ�:��>�	>�����>��f�{��;�u������>9��ʻ�>>�S��	������|4<˴�>�z�>//�>1���!4���̙?zK��ISο����e���X?]�?���?]h?ʚ9<��w��b|��4���F?&0s?�Z?-.%�m0]�§3�"�j?�_���U`�;�4��GE��U>�"3?�C�>��-���|=�>V��>�e>�#/�s�ĿSٶ�o���y��?���?�o�*��>`��?�s+?di�
8���[����*�D,��<A?f2>������!�0=�Ғ��
?�~0?�z��.�]�_?*�a�M�p���-���ƽ�ۡ>��0��e\��M�����Xe����@y����?M^�?i�?ֵ�� #�f6%?�>d����8Ǿ��<���>�(�>�)N>iH_���u>����:�i	>���?�~�?Qj?���� ����U>	�}?k(�>��?�p�=yc�>�M�=Y�|,�Rb#>u$�=I
?�?֡M?�R�>�b�=K�8��/�_SF��@R�f��C��>��a?�L?�Cb>����1��!���ͽY�1����?U@��,�Uw߽�%5>�=>�>a�D�O�Ҿ��$?��w8����G�|=<??��j=�VF?��7��u�2�S�~˂?�0>��/��5�� 5X��]��#'�?��@�?5���gy�<��>�F�>%�d> Խ�<�l��} c>��W?!"-��%���^�P�>nw�?��@\c�?�p�|�?.��>鐿Q݅��׾����-�=��D?�7�Blx>ڬ�>���=��|��3����x���>�$�?�{�?4?@c?b]��3�5��=�2�>��V?A��>,���󾓶)>��?���i��W��^?i�@NQ@�Z?7���G�ſNG����ؾ=�R��0���=/>�UƽAW=���=ҟ-������a�=B��>�D&>�ս�:)>i�=]:>03��#��ۼ��U�vp�����4��=��"��f{���6��m
�Q�����9��6��}ξL���Tx�����=L�?�wB?7�K?��)>�т���='�>���(>�����@��"�>�kk?<?!�-?��>�w���L��<.��.��!� ��j�>���=3��>�<�>*_�>L�,>\P�>5'3>εM>V�Y>b�������>h��>�%�>8�	?7�>�C<>��>Fϴ��1��l�h��
w�q̽0�?����S�J��1���9��Ԧ���h�=Gb.?|>���?пf����2H?%���y)���+���>|�0?�cW?�> ����T�2:>6����j�5`>�+ �}l���)��%Q>vl?)�f>�u>�3�w`8���P�ev��o|>26?ᶾs>9��u�'�H�b^ݾKM>Iƾ>|D��i�G������ri���{=+u:?�?[/���᰾R�u�	@���LR>�5\>Wt=�z�=$YM>$Xc�3�ƽ-H��L.=��=��^>��#?Α�:�F�=7�?7w�Xv<��!�>���>K�=*7,?�.a?�f�gH>ITe=#��=�Ų>U�>�@e>��
>�j� �= ��>��	>e��6���F�#�r_8����=����)C�����>��	�A��=cS2=����8����<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�Ž>4���{��ߑ���a��&�=Մ�>�=J?v �C���Ǆ�=I�>É?�*���|H¿�������>һ�?Pę?g<r�{٢�S�4�(�>���?��Q?�>nB޾�M��9~>�L?G�Y?�]�>-u%��2�{�?o��?5�?��3>�ԍ?yu=?+�>M�=��;���ѿ�l��>��>�>�>�{�>;�=Jw��󵀿�㱿�t�L�u�7��q�>+�:=�=�>}�y���~X���:��zپ���{7�>���>��>��V>�U�>���>Њ�>?�T=��u�+�Ͼw־�K?h��?2��*n�;
�<��=�^�A?�H4?�H[���Ͼ�Ԩ>%�\?ѿ�?�[?xb�>���_=��i忿v��?��<��K>S0�>xN�>&��HK>{�Ծ
/D��r�>�ɗ>壼!Jھ�*�� ����C�>�`!?T��>!��=�$?G $?(g>�G�>Ý;�Mʑ�y�K����>L�>�=?[�u?@@?j̴�B0=��h��{��ZY��b8>�x??)��>z����ڛ��t��J�y �c�w?�v?$�r�B�?�?�A?�.8?b�4>2~ѽd�̾z׽���>1�!?;6���<��/ ����ٴ?j5?<��>�Sp�1ǽ(O#��O�7R�v�?�r[?�&?p���_\�H}��.�<s<h��ߝ��;,hr���>4`>+����b�=��#>���=��e�=O+�i9�<)��=oُ>ư�=�9�V��'?�kv=𱦾DB��B�A�|� !>s}>>���;?�}޽�c�V�Ϳ_��3h���n�?���? ��?�J���v�`�C?���?Z�>���>ӈ����˾����U�2uv�w��W=z>��>0�>���ү�GD��<����~���(��p�>9!�>\+�>�?��h>�O�>����,�(�� ������WK�����D�E�2��;�1��+ҽ�<�*�Ǿ����X�>����]ߵ>�?�{>�[>S��>�~����t>��\>�{�>�N�>�_D> 2>,��=}��C��L\R?����uq'��6�5H��W�A?�\d?�M�>>�l��ʅ����IE?Wo�?PJ�?�w>Yh��m*� y?j��>dF��	?�9=�d�q�<H��� ��ņ�����9�>�(ֽ�8:��M��e��9
?�?PC����̾�lٽ ����`�=�Ё?/� ?�"��]��/}���^�(QE��;u�6d��<������x{��є�����l��+,)���<�R(?�W�?���c'��Y�-WQ�<�g��L�=�U(?q��>��>]�>"{ξ�uK��{��Ռ�1$l��_�>�cd?0��>�=?w3?��@?}[?���>�?�3s��}�>�/�="�>��!?bh0?��@?�ED?�� ?�?i�Z>�����Ӿ�#?eC?O�?�W?RU?��]�Q=��=>�q>�YԽ�DW�� �=�����	�^I���,�=ճ�=
t%?��q�$��m��<��=��?�n�>�j�>�󂾾����L>w��>�?�ޝ>���2a��¾�y�>�3�?^��a;��>���=dx���9��\�=*���S<�϶�섗=�w�fH�=m�=5��i3�=�3=ɥ�<��<�t�>3�?���>�C�>�@��4� �b��f�=�Y>6S>|>�Eپ�}���$��u�g��]y>�w�?�z�?�f=}�=���=�|���U�����8�����<�?FJ#?"XT?\��?|�=?bj#?µ>	+�hM���^�������?w!,?��>�����ʾ��Չ3�۝?i[?�<a����;)�ݐ¾��Խӱ>�[/�h/~����=D��텻���U��5��?쿝?HA�W�6��x�ۿ���[��z�C?"�>Y�>��>U�)�~�g�s%��1;>���>kR?ᦷ>#}T?��x?[?��A>�=�@w��Ü���v	��i>qs8?�Tx?���?8�u?���>��>s4�9���'�����O��~�D��<ZN> Ԝ>�c�>���>$��=���_���w.�k�=|�Y>ل�>"%�>[(�>@X�>��<��G?���>!��[d�������Z�:���u?q��?3�+?��=U�h�E������d�>�_�?m�?�*??�S�b��=��ּ#¶��r�=+�>c��>��>���=i�E=�k>N��>��>e&��X�1_8��O�B�?$	F?R�=������.ؾ5�,v�Iח��>�� ���򣆾0Y)�C����ھ�辯tҽt�+���R�ZF��d��X��T݉>�o>2n>nMn='�
>��˽$9^�l�z;���<���`�=v�j>:�ƻm�=oe$�<�M>���M��Y���bʾ��}?L�H?qX+?9bC?��y>�>��6���>������?�-V>�qP�Y໾�z8�(N��Xה��Qؾ0�־]?c��s��Ä>]�J�	a>��2>Z��=/�<e�=�.n=��=,N]�U�=(?�=]��=�۫=���=�s>!�>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?��>>�2������yb��-?���?�T�?>�??ti��d�>M���㎽�q�=M����=2>q��=x�2�T��>��J>���K��C����4�?��@��??�ዿТϿ5a/>��8>�>svR�#�0��]���a�Y��!?��:���˾�C�>��=�I޾Y�žT�2=�F6>�d=�����[�љ=�{��;=�i=8��>@�C>L��=�|���Ͷ=dLJ=zP�=�"P>���+z7���+�`�2=���=V�b>�#&>n��>��?U20?��c?*	�> n���̾�p����>R�=���> &�=v�B>�L�>�8?]�D?<�J?4�>>��=�P�>jV�>�,��\m��]�h�G%�<&��?
'�?TU�>��)<��@����X=��Bɽ�	?o�0?z	?�:�>���]�׿������O���0����<��c��8��6)j��z�H��} �<�Ӝ>K��>��>�W4>{��=���=`(�>mɶ=�=�4_=�#�=�u�=�7�=��>�c;�/�1d��?�;|'B=�1¼i=��6>�P�=f{=����,c�=?/�>]f�<�#>��>�W����=Ƿ����T�csE�P�w�4��ʾ��oo����5���i��>��>@8��KЗ����>��U>��>���?C/�?�~%>:an���X��皿zl�@1m�c-�>߯">K�N���U�H^i��\H�����>��>s��>��l>��+�Y ?��`w=&�_^5�'�>2|�����.��Aq��A��O���)i��кi�D?�C�����=~?S�I?���?��>N��T�ؾ<i0>�7��I�=��q�:e��8�?�'?ݕ�>��-�D��N̾���V�>JVI���O�jÕ�n�0�_�\ѷ����>c�����о�#3�f�����e�B��nr�g�>ݩO?(�?�3b�l\��}]O����v녽%p?`�g?
#�>�I?j6?�i���w�(}����=��n?���?68�?(>���=��?�3��>L>?,ώ?�+�?C�q?�����>�¸�Pl�=H�?�W��=pT>G�=%�=��?�?�|?��d����x������{�&��=���<=�}>��w>g6}>�4>G2=��)=G[i>|$�>��>
l>�Ƣ>zǓ>�S����"���2?�$���???h>��<c�i����O����q>l*���`�|���*Ȑ<دn>yh�>m�="M�>�k㿗��?�?�7�?�>�r��z�;>��*>`��=��.��>Ĩ�>]�8?rؕ>��?ժ�> �+��|�>��龕�?>-=���+a�
� ��DF������">w׾���kv)��Of��Bz��µ�8b�I;J�i���8��l���!�?<�j�����%�X��\>��D?n��>g��?�vy�HTI�H	�i�z>�Z�>G���M���g�+�о1y?� @�;c>��>-�W?+�?<�1�v3��uZ��u�'(A��e�I�`�l፿��
�C	����_?��x?�xA?[W�<R:z>G��?�%��ӏ��)�>�/�i';��<<=,�>W)���`��Ӿ"�þ8��GF>��o?.%�?(Y?�SV��R%>�S�=�L?w�
?�;?�7?��Q?%�j=p�7?��3>�f�>=?��?H 1?K�#?�D�>횽=�2�=F�<,��0.���/��`Ii=łr=����ڼ�Z-�Ei<bZ�=��Z>t�z<A6F���=ۨ��OB��o�=��=�|�= ߦ>��]?��>�_�>�7?���68����/?K�8=�ނ��݊�跢�0����> �j?kݫ?QZ?B�d>AB�6C��F>�4�>b:&>�6\>�\�>�A�|YE�ȇ=��>��> �=��I�ދ��ȗ	�z}����<��>���>�|>�덽��'>Q���^z���d>��Q�������S�2�G��1��`v�ka�>��K?h�?��=�W�X��Bf�U()?,X<?�=M?X�?D��=�۾J�9���J�M&���>ۋ�<���4���� ��g�:�r�:ȹs>�+��lQ��Ũb>���޾��n��GJ�N�羦2E=[=�y�P=-)���Ծ �~�x�=�`	>�R���� �6���ͪ��aJ?߃m=�&��P`W�����>JK�>6��>�9�Z�x��m@�����Ck�=��>�:>{���S��~jG��/�c��>YlM?k�Q?JRz?�Ҿ��y���=�mv�  ����� ?��?4_�>��>�w
=�Ⱦ������v��@e�6Ⱦ>���>�C���H=���E�-оk' ��J�>��>��
>�h�>��L?�}?(�r?|�+?%+?st�>�_#�;BԾ�>$?��?t�=�A���xr�>>��@�La�>H�?H�A�8x�>�*?R�!?``&?`|L?��?�K
>� ���S��_�>��l>�R� ⪿S�[>6�I?㜶>�\X?�-�?a�q>�=C��3�����T�/>��i>��!?�k?o�?T��>���>����	>�a�>�c.?��?�Ђ?��@>UV?���>P%�>EG���}�>)?w�C?��K?�2?�^?썉>G3(���<p#B=dN�l�=e�= ^�=+�=/�:��U�ٰ����^=�$-���[<�Yu=X<	���4�=�n�z��>R�t>ƶ���0>�9žd:���A>�i���ͯ��<[:��C�=㒀>� ?G��>�#�J��=g��>��>���W(?��?_�?f��:�b��۾�VL����>��A?I��=��l��h����u��af=��m?lq^?�W�x�����b?>�]?kd�=�4�þ��b�ǉ���O?�
?��G���>��~?�q?��>?�e�"9n����@Db��j�2ж=p�>�W���d��?�>�7?O�>x�b>�8�=�p۾��w��o���?��?�?���?�**>U�n��2�e�#����f?���>܇���#?nW��Y�;5�~������ؾZȾ�@���4y�&���(����o�,�ʽ���=Ԟ?[xq?:�g?��c?��x`�t�R�Zx���H����"�	�ȲA��D���E�Ęv�c��7����D����N=`1�,��?@�	?𴎾���>_i�MZ�@�����=D��Lۏ��J�=$z�=��=�}�=��ʽ�ۦ�*�p��*?&�>�3�>��?�V�ɃB�S(5�Vp@��¾�_E>{q�>)WN>Tլ>��V=�����[_������f���1���|>(�i?��+?�a_?�9���MO����gFO�\��%bw�~��>B�X>�C=�uо�����q�o�C�`���7��{�����_��=�?�9<�<�>��?�?9?��$�8��&ܾ��'>zb�>�|G?,I?JI�>���0���>�p?�+�>��>fR�+�.��j������� �>��>O?��h>������p��K���2��?OD�	�;��Y?��q�zt�
݀>?;?�NȽ8"<���>���;�H����-$�+H>!��>PB0>£�>0ؾ������}�������)?|1	?F�����)�?>�H?�`�>x�>d�?]�>G��Q�Լ<?t�^?a�M?w	C?���>��=�,Z�����j8=�_V><[k>җ=x��=��@Q<�D��5��<b$1=ۑ�g��@�<�^�k�	:�4(=��8>�0޿�i=�({~�C�'"����8���ċF���m�vi���־i���m����	��c������u�C�������D�?jC�?<$��RӾT���"����'��*�>�����<�ాK?9;����P¾����O��RSN�Ժl�aUh��?̎�����
d���즽��?���>'+�?4��8i�;K���ɀ>u$(=@]i�l�'�������׿���d�?�S?`{�Z�K�"��>ՉA>���>�<_;��ao۾x��>f�*?oF?�t?�1b�P�ӿ����o�&=�3�?��@�|A?;�(����\V==��>�	?��?>�Q1�wF�/����O�><�?���?r�M=�W�*�	�1ze?L-<��F��ݻ6�=�2�=\�=���t�J>�W�>X��EA�u5ܽ��4>Ʌ>�t"�����^���<#�]>��ս1��7Մ?�z\�mf���/��T���T>��T?�*�>�:�=��,?P7H�X}Ͽ�\��*a?�0�?��?+�(?ۿ��ؚ>Y�ܾ��M?TD6?���>�d&��t�\��=-8�A�������&V����=O��>[�>�,�����O�~I�����=�$�l�ƿ,�$��T��=1��d�Z�Eg�N�����R��`���o����)�f=t��=�Q>ҍ�>��V>�)Z> FW?L�k?�r�>>佔ʉ�Nξ�s�e���������r
�k�����%�U	����l���qʾ(�B��=�=��啿�)�2L��NQ?�q{?�J>������g���=|߾<"�������O��N��,�?���z���?F�3?����ᇿ�B��kżFEO��t�?��	��k�{	��D�=!����:xh�>a3>8��38��S0��w0?�W?�o��L2����)>�� ��=��+?K}?�Z<�>AT%?�?*��$㽈�[>�d3>�ʣ>A��>(�>����r�۽N}?��T?ͽ��ɜ�d�>qU���wz�8a=G�>m�5��2꼜�[>��<�Ì���U�5��MZ�<39W?�>B�)�1�����R�ȑ==�x?��?+�>f\k?��B?k�<f!��5�S�l��y=��W?*i?V�>������Ͼ�����5?��e?כN>��h�(�龞�.��K�1?��n?ZH? s���n}�3�����qg6?�mv?!E�� �����,u�58c>\��>�"?yZr�h>�]%?��Z��c���S����Q�ሦ?��@�L @w�=�
i�Ž/>�-??4؋�v3��q�=�Q��񀏼KX�>Hƣ�Sdl����|��dnD?I�?$?�*��h��K�=�ߡ�]߫?o�}?�_����W=����W���X?2�{)>S*��g���B׾sB���P���3���&s�==GV>�j@yU��A�>���=��п�����y���������?9��>)��2�!��f��~���Q�E�E��_��E�>}�>�Ŕ�a��A�{���;��[�>�����>�`V�+쵾Zϟ�>H<���>��>F�>߯�໽���?(���5MοLҞ�X��3X?��?���?y�?RC<k�y��2{����F?H�r?i�Y?�+��H]��K.�+�j?�_���U`�V�4�<HE��U>+"3?�C�>Ô-���|=�>'��>d>�#/���Ŀ*ٶ�������?ى�?po� ��>|��?�s+?�i�8���[��B�*���-�<<A?g2>�����!�/0=��ђ�E�
?00?�y��.�~�_?��a�d�p���-��ƽ�ڡ>��0�g\��<�����!Xe�����@y����?^�?�?޲���"�l6%?j�>����o8Ǿ9��<�~�>'�>�&N>GR_��u>����:� i	>��?+~�?�i?ܕ������EV>��}?�-�>%�?�z�=�g�>:��=������-�NP#>���=�9?�h�?��M?B]�>���=��8��/�yQF�)IR�7.��C���>!�a?V�L?�Pb>#㸽��1� !��Uͽ�\1�$��5}@��w,�t߽]5>}>>x>&�D���Ҿb�%?]X���翕/��
���j4)?f&�={�?����'��k��g?܏3>���S��Yz���t���?��@�?�L���ǃ=9D>��M>#\v>����[��{پY�=ɑt?r��c���d�5q\>A��?�G@��?��t���?���n������G��Q��0�Y=N?K����_>0�>`ʈ=�o��e��u�����>b��?��?P=?�X?�R������*>��u>s4D?h��>�Q=U��'�=J?4 ��(��oQ��G`?�@��@�R^?�(�������˪�%��o��H��>E��<�D>ސ�����=is'=�S���ԍ���o=9گ>f�3>kh�>v�7>p�B>�+>+_����!�i��Φ����)�*�(����!9�5j��2\.�G+�Yվ�vξ��"�
�+��$	� <)�� !���G=�>d7?�"?=pp?A��=�F\��Y�=a�¾�"=�8��a�=���>�1h?�i?��%?���<R{A��*S�SF����Z��׎��k�>�m�>U,�>��?��>5�V=�>�2�=� �>y�F���O�L+ �њo���>�8i>w��>���>��>%�>A������(M��h���ɽ�?�����PX����y��ڡƾV=��?<>�v��>�Ϳ�-���P?M�����9�ftb����>0�C?�X?��>T-���ė�u�<����2�� >�B3���D���,�C�W>�.?��f>�u>n�3�6c8���P�{���i|>r26?�涾B9�/�u�l�H�y[ݾXRM>yǾ>>ED�j�������oi���{=hv:?��?�<���ް��u�C���QR>�7\>�h=�N�=�WM>Qc�U�ƽ	H��h.=���=ʲ^>��?`b:>��=5/�>
��Z�B����>-�4>�DA>
�=?v ?�<�)�{�ߝ`�~���\�>�&�>/݁>?�	>�7�˶�=���>3�F>&'�$b��-�h>���^>AQ�� �n�����e=��=	�=#����6��]=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾHr�>���5q��|(��A�u�3$=Vu�>�JH?3f���]N�4�>���
?K?�L������ȿ��v�b��>��?1�?�m��0��u@�U.�>v��?9Y?�h>.�۾@Z�+�>D�@?g�Q?�ֶ>iO�ue'���?���?���?��>d��?U�2?d��>m�3>r=��۽�Sq��g��>��z>�>�>T�ͽ�3Ͼ爿����_V��lUv�p��rf�>o3=���>Za.���Q���=:�L�U
�o飾��o>�0�>\U�>2C�>r�p>2��=;[r>�*���*�_ܴ�b���3�K?�'�?���T�k���t<���=�t^�ZD?A�2?dQh���ξ�>�+^?�!�?��Z?<�>N���ښ�˿�oF��BS~<q�J>sd�>���>'t|��RM>d:Ծ�@�'ى>��>
6 ��;پ�\��Y	�ӳ�>h ?��>�K�=2� ?��#?]�j>U)�>a]E�M9���E���>���>�I?z�~?��?-ֹ�7\3�e��a硿��[��0N>��x?�T?�̕>Ҏ��炝���E�JRI�������?Mqg?�T录?�1�?�??|�A?U-f>���ؾq���&�>y�!?C����@�bD$�vc�M	?�?�w�>�����]սy�ż���$"��S;?GN\?/�&?�	�=�`�ֻ��q!�<�=�F�����;�����>)�>|q���_�=��>@�=/�n��5���r<���=�p�>��=��4��ǈ�Y�/?'�>$�n�uϠ��d���as�y:%>���>��(�S]?rB�g�i�#Ӽ�Z���#��{?�?�L�?mt�?�o�O�b���E?���?��)?(�>[����ս9$�[R;4j��U�ߨ�>x11?�F�]��r���ᬿm��������K-���?,��>��	?��?�}�>�=�>����&��j�h��8�H����|E�A.&��� ��>Z��7�ۼ]=;4r��+ٞ>Hf����>�?E�@>be>�R�>A=x��7�>�s
>���>��>˒�>dZI>���=bu@��?��mMR?g����'�G��°��+B?)ld?x'�>�h��������2�??��?�s�?�Kv>�{h��%+�Mj?�2�>����o
?�T:=y�����<�O�����qA�����X��>6׽u":��M��if�_c
?Y-?�����̾�׽}���[m�=j��?_:(?Ӫ#��TO�mo�"W�DXM�Y��n]�_l����#��p�^Ϗ�d��x3��K�'���V=�(?�?V��������k���B�b�U>p��>�\�>�J�>1�R>���6���[�l�'�k���>x?F?�>��@?�1?L�Z?�8?�.�>B�>G���!�>�9�%k�>�z�> XA?��1?�^.?�?�E"?�)>���Q�����Ӿ�?��?��?�o
?�w?�a��o���5����~4���֔�"=W��=��d��Z����=ί�>zX?���r�8�0�����j>Ձ7?���>1��>����&��� �<��>�
?�I�>.����xr��`�bR�>��?�
�s=k�)>i��=�u��s�Ѻ5S�=������=���w�;��<��= �=Ws�]�}��m�:g؇;e��<�v�>��?̑�>�9�>K��/� �������='�X>�S>�>yDپ���W%����g�-my>�z�?�{�?L�f=���=׮�=vv��G�����*����<՘?bN#?�ST?\��?s�=?t#?�>$�P���`��?��2�?x!,?
��>�����ʾ��ԉ3�ם?f[?�<a����;)�ϐ¾��Խ�>�[/�h/~����>D�l񅻺��c��2��?￝?6A�O�6��x�ٿ���[��x�C?"�>Y�>��>R�)�}�g�j%��1;>���>kR?���>��R?�Gm?~�O?/�=��?��Ԣ����ᵽ���=�e0?�$�?;��?yp?���>��=��7��� �@��]��9��n�A<SX>��>4p�>�>�P>`ؿ�#9���)��!2>Xf�>��?z��>b��>rb�>�T�<K'L?���>ٴ���
ⷾbቾ5�)�]�k?&�?s�%?@��<�~�>3B��x�Z��>^�?��??"+?_j:��?	>o>Źn�����x��>�6�>�F�>?Hw=�D=�	>��><��>�:�_���8�(hw���?�[A?�v�=0�̿�Um�EN�X얾F�.=(��S#X�g��фa�����ͷ�B�_����N5b�#��|	��6ɸ�K��|���z?���=�b>�{�=�bͼ�o
�a�����<|��=}�<Y���	��=pn���=�Ž��5=C�O�����/m���˾��}?�:I?h�+?��C?��y>#Z>&O3����>�?��6?��U>��P�P����j;��������[�ؾ�m׾>�c��ǟ�}K>�I�!�>{M3>�A�=�p�<( �=��r=���=d�U��.=_2�==K�=�g�=X��=��>pb>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>s��=w�2�T��>��J>���K��B����4�?��@��??�ዿТϿ6a/>�7>c>�R��o1�]��b��|Z�>�!?c<;�i4̾��>ڍ�=Q�޾%@ƾ�/=�$6>�ab=ò��i\���=͞{�d;=��l=a��>�/D>f��=�ԯ�3�=&TI=���=�VO>����6���+��3=н�=џb>�F&>�I�>��$?��.?�E?ҿv>b�y���(ž8�>���=�˞>ؚ`<^�(>r��>��B?��=?2.P?Z��>�'�=t��>�>�����s�Pg��aо�0˽�y]?P u?	�>De��?�*�����&�< �;��>�,?ʰ?��>���꿙��V!�Zqͼۄd�"��=nh:�p�E��z=��?��H�@�>���>	�>:�>��>a�;>LT�>��>��>5�=$>!�_=>�V��c��Yd�<����v�=��x=�+<)�<����9�FO��_x�<��=����1�=��?�%�=�$�>4O=������2>T��f�X�@��̪��(H��Q��w��n�/�b�L��8�>>R�>�m�S쓿��>9�>�P�>���?���?�#d>�di�>�K��������L���C�>x��=8CG�A�R�w����[��_����>��>Y��>:�l>�,��?���w==�d5�*��>'w��u�� ��>q��=��<���Ni���ƺ=�D?�F��gv�=7~?��I??�?7��>���Q�ؾ�Y0>�M��-=���p��N��5?�'?�z�>���D��H̾L���޷>�@I�5�O���T�0�V��+ͷ�(��>������оm$3��g��������B��Lr�P��>�O?��?F:b��W��RUO�����(���q?�|g?.�>�J?�@?�%��z�r���v�=�n?ų�?M=�?d>\�=���x�>��	?��?CP�?qJp?#D3�E �>����څ&>ל�ɂ�=�U�=bo�=�<�=��?��?�??l��Bn�O-ݾ�����Y�k =�wm=a@�>���>�&X>wջ=��	=L@�=U�x>�D�>e�>u�b>���>⁋>����:����(?�b�=i>�>P2=?	�>�<����@���ه�������+���|������=DH�=T>g�=c��>�ѿ�̩?c�=P2���>���?����>�1
>�����=���=�y ?�>>Z��>>oG>�t�=��Y> �оZ|>C���&���;���R�ڻξ�u�>顛�"7�3�>����O��,�����`f�q⃿��>���<{"�?HD��Fo���(���ν�?�_�>��8?�莾637��i>��>��>O��C֖��� �C�?�w�?�0d>(�>@�W?4?�&3��2���Y��hu�^`@�pvd��V`������e��*�	��ߺ�?�_?�x?�A?!g�<K�|>��?"�%�ɐ����>	o/���;���/=���>ˑ��)a�58Ӿ�Uþ���q9E>��n?��?�Y?��S�+=�M�
�?��(?�4?0T?�yn?�n�<��?�K�>���>��>6=$?��)?Y�<?��>�`�=�y=�x�����`d���F;�Y㊼f����0�=p!��9���a>�H�<�'��<!�ñɽd}���Z=E!"<2�=�g=cæ>��]?L�>���>!�7?Y���t8�Ʈ��+/?��9=+������;Ţ�t�y >e�j?T��?�bZ?�ed>��A��C��>SU�>�n&>�\>Pb�>�|�J�E��ه=7H>�U>W¥=ugM��́� �	�n���B��<,>���>�|>�L���n'>D����-z�~�d>mR�������S���G��1��nv�,��>%�K?;�?HL�=�"�䅕�uf�L)?<F<?@,M?��?�-�=z�۾T�9�J�J�-[�L�>��<t��᳢����`�:�v-�:קs>D���~���u>;޾60ھ�Hn�]�S�}������~���>���������x�7�
>�>&�ξ�2(�#������WH?my�=����!�� ���[Ί= ߝ>���>������	��0C�ڳ��|8=iw�>�i�=�̅<���@�����l�>q A?(HT?X	l?�����N��Ky�R�)������߇��s�>�p>��?�>>G>ԣ۾�e&��a�۹J����>�V?Z>���S���	6�E!;�v�5>�;?��m>,��>�2?�?�2?��;?�U�>�k>u�������$?�?�?��=������r�0�!�H�6��>^�)?�*۽^��>[0?�]?�?��S?C ?5*�=� �E�@��I�>�_�>!eN������L>��=? ��>X?B��?�u>�3<�͙���_�=��=�>u4?7!?�?�<�>9c�>�ۮ��U�=���>��e?�T�?�Vl?f��=G,�>s>�: ?<>�=%�><��>��?�.E?�o?�F?��>U��</��b0���!9��˼%b���<׌=�fL��"W�=�C���<� <�%�M=�;:?��p��Lk��<���h�>�5t>x���0>�qž�C���?@>�������W���:��=�=&��>��?�ו>f$��}�=�Y�>���>=��|+(?7�?�?�v";�~b�`�ھ�K��2�>pMB?��=s�l������u�y^j=��m?�f^?$mW������b?��]?�d�=�f�þ��b� �龴�O?H�
?L�G�L�>9�~?W�q?���>5�e�F:n�����Cb���j��Ҷ=r�>OW���d��8�>�7?�Q�>��b>�:�=,p۾�w�r��"?�?��?o��?P,*>��n��2�	h�)M��kX_?�>����-)?��<i;ي�Qʡ�mu��w���d���yNx�����Ƽ"��w��нH��=�e?��}?_�d?c_?V��Z�c�iS�,���b�r4򾊮���9���4�-�<���^��f��������{x��8J�es�?��%?��
��Y�>����m��Dʾ�2>8J���8����=J�&�ܜ�<Y~I=��\�k�*�]����?�V�>'+�>S<?�X�B�>��Q*���:��4�`5>�:�>���>�#�>��� .��P	���ܾ]����>��b?��>?�'E?h+ξ7�1��+����2�h�=�+��(�0�`���>�b���ע;�=���=�"�p�����)]�/�־j��=Xm?�=��E>k8�?�l�>�F���1<��2�d���ʰ��+0>��Y?E��>dk>уe�ơ���>G�l?z��>�-�>2���fi!���{�7l˽�`�>��>��>4o>��,�c,\�RB���z���9����= Uh?xh����`�oŅ><R?*��:@:<�R�>T�u�2�!�@���o'���>�p?�S�=�;>/bž�e�{�g����6(?6?�^��^7(�G]>j�?�A�>��>ꌄ?�v�>�ξa�Ӽu�
?i�X?y$J?��=?&��>W$�<�	ͽX�Ͻ3�&�7�&=��>h�a>#�c=���=%���`W��5�%�)=p��=V�����qn�����IM�<}��<��*>3�ֿ/xJ����j��sҾ���� ��-�T�䥾k��<����q�y�_��<s���T��O��*t���G��MRP�`T�?e�?��D�F����f���������U�K>T���սQ���˽46�� B����ɾJy���^��d������&?�百A�Ͽq������^�?�(?]��?n�����O� [�>2R>ڜ =<�	������WԿ|���q�x?��?i���M�$֔>��>;��>�d>,���kX��2=�.?��T?��?&.h�JPҿ.���*�U=G�?�{@�xA?��(�}�쾠EV=���>R�	?��?>mS1��E�E��Od�>t6�?��?/�M=��W���	��|e?�< �F�̡ܻ��=Ja�=U�=����J>�Y�>u���iA�sܽ\�4>�Յ>Ln"�`����^���<g[]>ֽ�p��4Մ?'{\��f���/��T��U>��T?�*�>h:�=��,?[7H�a}Ͽ�\��*a?�0�?���?"�(?<ۿ��ؚ>��ܾ��M?^D6?���>�d&��t���=<6�d���~���&V�]��=Z��>f�>ʂ,�ދ���O��I��O��=�� � ƿ�)�%�M�=#Z��LI�65��K��Q0=I������wIX����=Y��=O�>x�>ego>ܺ�>V�S?�k?�N ?�Y>��޽l���!��<� ��}Ӿ�8��򊾙�"�)5����Ѿ78�{���,)��k&�z�о�<�쵂=��D�ⳏ�.T��t�n�K���?$��=n����A���I=N	ʾ����G��5ٽ���ˑ8��o�uޡ?�y=?Zd��,�m�P+��X���А�J�k?%�'����v�ľ���=��
�?m?�1)}>TF�=��ﾖ+���F��n0?�g?!f��S���)>*� ��D=1�+?+�?PL`<��>�*%?+�+��O�[>�w3>��>���>f�>����Q۽^?��T?=��
����א>uD����z��4`=�>�I5��<���[>b�<�㌾�kT�
L��w|�<�(W?t��>��)��ia����NY==��x?��?.�>j{k?��B?HԤ<3h����S����aw=�W?.*i?��>����	оX���E�5?�e?~�N>�bh���@�.�VU��$?�n?<_?�}��'w}���l���n6?m�?hZ��{��e��KV���>�ȏ><?��p��Ma>�?+�v�&¬��κ��h�2�?:@2��?�D>3�޽f/�=��%?.?M�辞�Y�=��Żg�?���dۖ�$����H"?���??�n�����qS�=�B���J�?Rd�?,�g�@#�=�`��j�_�
�% ��Z%>打��Y.��\̾P�/��о���XF�����(��>{q@�� ���>q��8�׿܂�~p��K�������Os�>�ڞ>]�b=�G����+�WCi��?W�2^K�ߕ��ݢ>Z�>�[���o���{�v�;�
]��B0�>�q�xԈ>V�S�ٗ��@���ċ<<�>��>���>�籽jE���Ǚ?Z���lο�Ξ��P���X?uN�?��?�0?�<�x�#�{�=����F? �r?]	Z?S�(�Q�\���4�1�j?�_���U`��4�IHE�9U>�"3?7C�>m�-���|=H>�>Zf>�#/�~�Ŀlٶ�����m��?���?�o����>k��?�s+?�i��7���[����*�k,��<A?�2>������!�Z0=�OҒ��
?�~0?�z��.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�(�>_�?�(�==}�>o��=�`��R7�+�">a�=u<�MZ?�uM?!�>�o�=B8�P/��QF�TR��4���C����>Ⱥa?�_L?�bb>Ӹ�c).�T� �6�ͽ(�0�\���^?�"�*�߽��4>OP>>�?>tD���Ҿ1�4?B, ��忰���1B�<�2?Ź�=�-?]��k��xT�;3��?A&�>���x���^m��|����?�@��?0ϾC(���6&>O�w>a_�>Ʌ�������9��(�=��q?5�5����tn��_�=��?��@��?�e�=�?������Z������8|ӽ�6s=��F?�����7>��?�&>5�~�Ո������a��>��?	��?��?B�_?�d�--���>Y�t>U!`?���>�A�p����C>���>,�2��♿S��}V?�F@xe@�\?i���p�ܿ2Ҡ�Sٴ���ľZ����I=���>��=2�	>F�+=-k%�~�z��h>��>6۲>�4�>h�@>�r6>�)R>�����9��������vZ�5�����=]IݾښQ�['��B޾|��^�7�.{�=QM�4A�����(R��|>!]?�D?�Hu?s�>=A���H0>�?��r>vQ�<���9C��>��=?ˎ?�.!?�=#={I���W��f���j���ゾЬ>��>%��>�8�>�>�>;L�z�L>a0>^d�>uy>�	>v��>ч�=��>Sж>>9?��|>�B<>v�>Iϴ�32��1�h��w��̽� �?ك��s�J�2���8������Wi�=�`.?${>6���>п�����3H?�����+���+�K�>��0?jcW?k�>N��`�T�
4>ֽ�C�j��^>�2 �#~l���)��(Q>�n?4�x>�>r��O"��lh�ǒ��;�M>
�?��4�g>��ꄿ�_�{���H�=��>��lb��@��2n��o��=�3"?��?���<������z�Lfv��/>���<!g�<4�f<��`>L�f���U��M� Ћ=�y�=H�*>�A?Pt3><�=�>�*��9#P��^�>@:>Y�1>#�A?�A"?�m!�����cƅ�&��r>+!�>�/z>��=PUJ��2�=�o�>�[`>�\��ଆ���Ԧ9���Z>��t�0Yd��s��	>p=�������=rG�=)���ʦ=��p*=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>���T#���㈿ݳn�Ȁ!=�5�>�HJ?����mm���T�?��?�?뾈|����ƿf�z���>S��?��?P~l�᛿z�@�C��>���?O�V?�9w>{�Ҿ�S����>��E?�YT?��>��!���'���?���?0�?gzr>�}�?��Y?���>:y�q�'���^⇿�P\>���=��=������]yO�CH�Ů��I_���$�#2q��1=���>���I�c�3e:>]b^��O��U�ܺ՘�>�p�>�pB>YP�>��>A�>>��=�M��Ăv�E����K?���?�X��m�`;�<�ě=��_��V?MR4?6vA�Wоr��>0\?�M�?z[?KP�>u���#���ɿ��C��鏚<�K>���>q:�>�L��A�K>RԾ�B� 3�>���>�U����ھ#\��	I���V�>�!?�'�>G��=ٙ ?��#?��j>�(�>PaE��9��e�E�~��>ע�>�H?��~?��?�Թ��Z3�����桿��[�(;N>��x?
V?yʕ>X���ꃝ��mE�uBI�����W��?�tg?cR�?12�?ω??H�A?�)f>���ؾl�����>�B!?ʉ�7�<�x%�s�)��?�4?��>�`�g���N7���V���A�	?#r\?�6#?�=�HPa�H�ž��<��޻(U���&<��,��->�X%>}O\�|s�=٩>��=c���4����<�d�=���>p��=��9�=A���0?��ؼ	��:y�<�o��/_��ς>y�K>��4�R?2`��W#��`{�����۾9Y�?E�?���?�S�=��i�;:L?%3k?�?"�?gލ����5����R=�G:���x��=u��>&������������[�����!�Jk�>hX�>K��>�N?>��>��>>C\����E�|	۾>�c�A;���M��=���&�i�b���e�4D��Jƾ.7��?�>��+��S�>͖?
[>2�C>d��>�!��#�>G��>���>�?1�>��>��=ClX=ɒ���JR?����6�'���辦°��.B?ed?��>��h��������y?솒?So�?uBv>��h��-+��g?�/�>����n
?�P:=�K�kL�<�S����X'�������>&F׽�:��M�Y�f�Qn
?:+?�	���̾/B׽������m=zC�?��(?�)�4TR��o�tX�KS����Lg�\����$���o�7���MY��l(����(��#=��*?��?���������:k���>�+g>�J�>f��>�=�>u�I>��	���1���]���&��E��x�>5�z?x��>��J?�v=?'lQ?�FJ?�ւ>�e�>J밾�?V�	=�Z�>�s�>y=?�0,?B�2?�?�G'?�N>�#�yL��(̾�w?(�?�?���>>�?�T���^�e��_}:�v\�I�e�,�=��M={n�SA���K=�X>CX?b���8�����ek>�7?��>���>����1��7��<��>�
?ZO�>�����|r��^�yW�><��?���`=��)>���=k���{�ֺ�T�={�����=b��Cu;�؍<ꂿ==�=ͭn��[z��:��;�M�<u�>0�?���>�C�>�@��<� �Z���e�=mY>TS>>#Fپ�}���$��r�g�8^y>�w�?�z�?�f=A�=V��=�|��TU�����Z������<�?AJ#?XT?]��?x�=?Xj#?��>�*�lM���^�������?E!,?��>���޲ʾ��l�3���?PZ?L;a����%<)��¾a�Խ_�>�Z/�P/~�}��ND�b��f���~�����?���?�A���6�?x�n���#[��T�C?�"�>�Y�>��>l�)���g�%�1;>���>�R?L��>{EP?$z?��Y?�E>�7�ǒ��=˙��K���'>'<=?�`�?t��?��t?���>�>�/�\����������:�X���>�B=�?X>o�>���>�˩>"t�=�4���ɱ��0<�G��=.�_>c��>�l�>|l�>=�u>�2�<�G?���>�U���������,Ń��=�`�u?ߛ�?�+?9�=v����E��J���N�>"l�?G��?�,*?��S����=X�ּ�߶�V�q�*%�>Kֹ>'4�>+ܓ=*�F=�R>��>��>�$�j]��r8�<>M���?%F?u��=:�ſ��q��Np�����/Tj<����=�d�J�����Z��R�=�V���������x[������f���ĵ�����/�{�k��>��=�C�=��=���<f˼�]�<�
I=m4�<@�=��p�#Fm<��8�!ѻK戽`�.�/VR<�(G=�V��ž�~?��G?}L+?OT>?�ni>��>��[���>܏h�D?FiF>0oV�߫����1�����#���Nܾ�-۾�A`� ����4>/����>	�!>b	�=+7�<P��=��o=k��=!�j<��&=)K�=`
�=��=��=�c>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?~�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>s��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>4�7>�>��R��m1��\�lb���Z�y!?u;��%̾���>aŹ=A:߾кƾ��.=�6>��a=����U\�~��=�R{�T<=aWm=���>}�C>ӽ�=1��8��=�<H=_�=|P>�r��OL7��+�%C3= ��=��b>>"&>���>X9?YJ0?3�c?rF�>%�m��Ͼ�'¾A��>�u�=zs�>lF�=z�A>�l�>�8?�D?�K?�v�>�&�=4��>hQ�> P,�z�m��>徨���塚<�~�?B׆?&�>��+<R�B�����>�SJŽO�?�21?
?��>�����忒�&��\,�$3�:�:�D>�:>L��=��<<9�z�F�T>dW�>5$??��>�To>�=4>�F>k'�>fn�=�a{=�>��/>q�0=�a����I���G�d�$=��w�:�׼�i�ک�{Խ��q��w�;t�X��:��=���>B�=v��>�P
>�ߖ�@9>7<`���G�į=�G���\R��s��ʍ�H�C��p0�j�>���>����e�����>��l>�o>_h�?�w�?Nh>~��K�f������)c'���=2�X>��1�m��zq�T~X�M����>�>v	�>w�l>�,��?���w=!⾷[5�#�>���~���!�j8q�q:�����si�nFں�D?�C�����=1~?L�I?�ߏ?e��>M�����ؾ�D0>-���(=P��Dq����?�'?Y��>���D��H̾6���޷>�@I�0�O���[�0���Gͷ�,��>������оh$3��g�������B�Mr�7��>�O?��?E:b��W��[UO����?(���q?�|g? �>�J?�@?&��z�r���v�=�n?���?K=�?�>���=q����p�>DX?���?)ɑ?��r?ф;����>W�Ż�+>����9�=�
>��=��=��?�#?$�	?�4����v�쾵4_�Q�<�`�=T�>j��>��h>���=.��=Z�=�/k>��>c��>�uf>t�>~��>K���9��S?i��=�z�>�K?rx>3V�=��ٽ�����7>��K���g�f��5F����<A�=�yA>��=n�>��׿o�?�!�>�}���=�>%*߾��&Ct>�*>���<(��>�G�>��?��>���>�{�=��=��*>A�¾��=k���B���#�ەj�G�:�}>�@�g>p�d��9wT�q�Y��ې��1��	S�������I��7�o�?�n�ʽ��1zN���'=[L-?=s�>{fx?��J���%��4��;��>�C�>�d������l�w���?���?	<c>�>�W?њ?�1�[3��uZ���u�'A�e���`��፿Μ��5�
����-�_?��x?�wA?L7�<�8z>뢀?��%��я��*�>�/�3';�f?<=�*�>�*��b�`��ӾĹþ9��FF>��o?�$�?Y?�RV��R>s��>C�L?{�e?2b^?��+?��r?�~�=�Q@?N:�>�1G?IV?�S?5dO?5�?3)=���>�����=SnE���{�J�������`<G�M>0L�;ޚm<d��:+|�<@/�<ˏ���ϼ�?>�m����2��=Hߤ=�>���>گ]?�L�>���>�7?���n8�ٮ��8/?F<;=����le���ˢ�,��.>x�j?߫?�#Z?Ġc>w�A��C���>p��>��&>��[>a�>�Y�0�E�m��=�w>Ȇ>.�=N�큾m�	��j��jr�<P#>/v�>B@�>k�J�j)>�E��Yw�R�O>�?_����yF4���N��E;��dz�Y�>�$I?�s?yO^=���!��C�_��!?�4?��M?k�?�i=�]�!<4�T�G��:K�^'�>��=�5 �Y���ܠ��9�g	<N�w>�[�����w_`>�
�[�ܾ,�l��QJ��辰�,=���rx\=�/�rZԾ��}��}�=[\
>�꿾�R!�v���Mڪ�]J?2�w=�;��x�V�.f����>˗>$�>�@�#�g�V�@��Ϫ��}�=W��>�54>Ju���k�{E��r�#W�>c|F?#�f?J{?Y����l�S�5�,s��Fg���;c�<|	?ʠZ>�:?8��=�>�3߾J
�R�h�!�J�6y�>�;?X���yM�u�]��Ⱦ������>��'?T�=���>�<?���>~Fx?��=?��?�!�>�X�~,���f!?���?��=�^���/�����Qx�3��>l�$?�H���`>���>iB-?a�?�N?0"?��=���7��y�>�П>I�(�����=�D?	K�>f�f?B�u?SE�>Υ'������?���>\�T>e�@?��?
=?���>s�?��¾����J?iU?���?`�{?e<>b?���=�?�GD>f��>ǖ?l�!?��-?�Mo?��@?R��>t �;� <|\P�> ��rd>$B�<�r9�;.�BνcC�N�I<��=%�)=��A=X�i=z��<0����>��3�=`�>Su>ꕾ�h/>�ž�F���A>].��V���1z���O9�p��=��>�3?Y�>rO"�zA�=�V�>�e�>�����'?h�?��?F
W;��b��۾�/K���>³A?�h�=��l�f����u�l�b=?�m?X0^?�6X�/m����b?1�]?�F�=���þ��b������O?��
?+�G����>��~?C�q?j��>��e�9n����oDb���j��϶=�i�>R<��d�N�>��7?pg�>��b>Ot�=�۾��w�󇠾_?���??�?6��?y *>
�n��&��a��˙���e?�Y�>�ڝ���*?�Ż��ؾ$ ��:㟾o�پ
��v�����VV���;���u�IzܽR>��?ӌg?i"m?��^?�����i���S�bar���W���go
��dC�̺8��&=��s�4I�0���趾�]�<�g��0K0�W�?qk"?�J��/�>0��hD�MS߾�&S>|p��pb[;4��=V��s�n=�~ջM����F)�Nɾ{?�#�>%�> �S?IdG���3���$���4��3뾢�8=��>���>O��>o��<�����&:��~Ҿ�Ԃ�Q�����>4�B?��U?�11?$�B�|�4��^���>��LI>��i>��v>$?fnZ�V!���4�"lC�K�y�A��h�Y� @̾�}�>.+?��t<�m�>�0�?IX�>�R�t�������H�P��=�F�>�n?���>�=NA6��� ���>Uyl?�$�>e�>ϓ����!�>�|�.-ҽ�!�>�'�> (�>��s>�")��
\��3��i���8�X��=��g?�E���`�U`�>H�P?bq���o<��>�t�;&"�0��s$��7>��?�\�=.y?>�ľ�-�D�{��m��{�!?�Ue?��@��O���+־S�4?��S?�h?>K~?�?J�=�����R>?��?bU�?1�?��>�l&=wa[�Kh�eK�T��<�y�=\�>1v��tD����
`)����"2>C�:r���X�=Q��2 ǽ>}q�r�R=��>�rۿ�K��!پ����#�*C
��?��������ſ��ش�vh��6x��q�F$$�*�U���c�:��<�n�kY�?��?����#��4���H������'C�>�Rr�4�~�(��ֲ�����J��;9��	!���O���h���e��	'?
���&ɿ�=����վ� ???��z?����5"�k'=���&>:z"=L.ݼ
��_噿�ο8����c?ϓ�>���|ƽ�.�>�ą>�M^>V�i>��x��n��[�;�?*�.?2��>�w�3�ȿ-�-��<�3�?��@�D?�10�k������=W��>�?u�e>P��H�	������>�?ʸ�?���=�GM�fr��B8c?oZ~<�@���5<���=�4�=��l=p�н�^L>L��>��+��*�Xk�<�.>�J�>���;���]�.���<�Kb>�מ�.�W�Մ?�y\�f�9�/�U���T>��T?�+�>Y>�=y�,?G6H�%}Ͽ��\�-+a?�0�?���?��(?�ڿ��ؚ>8�ܾ��M?8D6?��>bd&���t����=#��������&V����=Ѫ�>q�>�,�5��N�O��V��7��=����ſ����#����=}a5<l�m�j���������6���z��?z���=]�>�EF>��u>]&2>Z^3>IU?u�j?��>��=�b�����u�ھ��:�@�z���C��2k�F�½����|���ξJ�����7t��rӾ{=���=:(R������� �$�b���F�w�.?x^$>x�ʾ�M��0<ʾ8���d��5��u>̾
�1�1n�:͟?��A?/���W�X��+���F����W?k#�����!��!�=2����=�՜>몢=����3�:\S�T�+?3~#?�m��#���ت=����=�/?��?�3=iU�>34?XJ����J�>�0M>$�>���>�N1>��.:&�]/?��k?��[�r��)Q>�ž�*���,=��=Q�,�J����">�s�B���`���s۽��=D�W?'��>q�*�͟��f����ڼ�Lm=��x?q^?���>�!l?I�A?�j�<���zQ�X[�%a�=guV?��f?c>�z�:о�n���l6?<�c?I�R>
�k��a侙e.��o�:?پl?\(?��ӻ��{�[�����*6?�{v?�l����Q�羓m����>�8>-6?g�]�N@e=�Ǵ>�s����09��L+j��/�?2�@f@�+=�洽���=��6?N�?���r��i=�}ɾ (5���?��� ����	��"�� 4'?��|?o�?���"Z�+�=Q!оȩ�?ke�?��?�*�������c�N�1D��X>6UN=�=�<%%��T@�MG��Z� 햾zG�=��>�@�s����>�o==S�wٿ�\g�6�!��A���>C��>��4��� �׷}������B�`?�~fѾ\I�>�>铽�͑��~{�i;�*�����>f��eJ�>�eW� ���
��-8<v��>t�>B��>䌯�0H����?=���l�ο?����:�X?�
�?\�?�?�M<�|�3�1�����D?0�p?[nY?���}]���&�%�j?�_��yU`���4�tHE��U>�"3?�B�>T�-�Z�|=�>���>g>�#/�y�Ŀ�ٶ�=���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�ü
?W~0?{�g.�]�_?%�a�L�p���-���ƽ�ۡ>��0��e\��M�����Xe����@y����?M^�?h�?ε�� #�e6%?�>d����8Ǿu�<���>�(�>�)N>jH_���u>����:�	i	>���?�~�?Rj?���������U>�}?���>���?^��=�^�>��=�X��{-@�p�> ��=0�=��?�:L?���>
v�=3N7�,�/�nkF���R����T4C�Vو>-�`?�NL?��_>�`���|(�
���(ֽ��0��ʼ��A��>�M�߽ 	0>ڵ:>�k>�4B���о�^&?�~/�A￪������<9:?���=4?tc!��E��(�^��5r?��>� �n���aFa���R��T�?��@t:?�%ʾ���<V�^>>Э>8T>S�4�a�<���1-_<�Pf?Y���d���F�w�w>���?�@�h�?��l�"�?��+'��<�}��	վ	�	�vP=uoH?���>]K�>�7�=  ������s����>mw�?�6�?]?�_a?�$b�
'� ��=��>�Y?��>��λ���U�!>� ?q� �c.��iu��X?� @�A@f�c?Ty��tM޿�Ȓ��Wp�;o^�2��>1:=v��=B�M��������b̙=l%�����c�`>�3F>�d1>���=ޕ�= �>X���O��+K������$������CDK�?n�v�ڽ��$�&2��c����s��Z�T����;:�9$��ܠ8>΄R?�5N?'xY?b�>�ϴ�y�>bM�#@L=�eY�#���,��>�
j?��"? �?�
�<�ף�ѹv�
/p�z�{�D�н���>��> ��>�Ʋ>�X?�`�<�����4>�z!>� �=ƒ�=�^��Q���U>B�>�>���>�C<>^�>3ϴ��1��\�h��
w�̽,�?b���/�J��1��S9�������i�=Cb.?J|>����>пO����2H?����y)���+��>��0?�cW?D�>���>�T�j:>I��r�j��_>a, ��l���)��%Q>Yl?�1g>)w>�3��K8�RQ�ύ���)~>-r6?�l��M�7�3�t�?I�ߒݾ��O>�+�>}�&��
�����}��zi�B�p=�k:?,�?(���l���w�&v���P>��[>PH=�m�=�K>RPk��'ʽ�YG��,=�/�=qv_>��?��>i76=逷>����VvW��'�>��r>�Y>��5?M:(?,J���ƽ�����Q�s>�S�>��9>�&%>s�,���켯R�>��>C�<p�>��8 �\�>�ա>߀��o'��8=�v�=�A����=�:&=ڶ���C�{�i��~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>��B�맿Î��tJ�El�=���>0JP?sr��� ���޾��
?��?�� ��˫�Kռ��{�Xʻ>�|�?��?~l�������<���
?A@�?��9?��>�������_�>%�@?��f?��d>�4��Ľ�h�>lo�?{�?��g>Nk�?�J?D{�>CZ�=��]�4ÿ^�����>Ҏ'>k�H>Ē�>�L��_�&��#��NWT���	�vk=W =���>,����z׾c� ��n���~����-�%%?s��>�&�>G��>ק?X0"?AU�>��=�5���t������6�K?8��?����m�l��<�Ɯ=��]�1�?�=4?%=^�S�Ͼ��>��\?ׯ�?��Z?�v�>���=1�������9���_�<�fK>R��>���>GU���L>��ԾaeD�la�>5T�>_v���ھ*��$���R�>YJ!?�p�>1��=;H ?�.#?>�j>�p�>�>C��}����F��n�>�8�>�?��}?��?���ɐ4����=$��+^[��N>$�w?�?�ט>�����/�� �*��Ua�\駽rʁ?Zti?l�׽�}?'��?[\??�A?5�c>�����־�����O{>�� ?U���):���(��?���?r�?�g�>�4�[gu�~�9���pr��?�_?�'?*���yX�7'��m��<*�K�񂋼hм$��Om>C�>G���S�=x>;̋=��o�)�?����<m��=�b�>z�=)�=��?��&�+?�垽ʯ�����=R�o�.^j���o>7d�>zN�dR5?�ս~nu�֕��R����ؾ�V�?���?�?�Ce<zIx���c?5 }?F��>"?)9�4��_��n�q�S2U������>�8�>�h=}�ɾd湿n?�������i<�cS�>pʱ>Y?ޯ5?��>��>�܍��}:�z�=��5�+O�����K���2��! �&z�c߳�����]ľҁ�m��>�گ���>�,?p;>ɟ>�D�>Bb�����>�>�e�>D)�>\�>{�+>���=d�=H��Y?P�羳q0������Ѹ�f�J?��n?��>X��=J넿��Ӿ��"?ۈ?���?��><9i�7W�	.?���>�z[���?��"=�0=2��=/���il��罪0�Iz>$氽���[;�"��?5�?_�;���G�=��k���g�;Q��?�3&?Oc�yYZ�Z�n�p�o��uG��Ǯ=u8��'ʏ�A� �S^O��Ǆ�xM��Ϊ���Z�7�i�d�,?5>y?<.�8_ �'���=F���6��}�>r?���>���=�rR=u�øM�f�����h)����>�W?:�>"�H?�c:?�&P?�qI?�>}թ>V*��u��>:�B<,Q�>)U�>��6?��.?kC0?i?4z)?�J[>�3��;����۾�?�w?��?�h ?�� ?�2���ҽ�x����'��Lk��j�^t=���<v�׽O�c���;=�K>��?�c�(�8��%���h>��7?���>�2�>����q}��X�=DF�>YG
?�b�>�����\r��r�vX�>�?�?C����=7�(>���=mR�\����=Zkм��=�����;���K<�=���=Z7m��":��;@��;o�<�t�>-�?���>�C�>�@��,� �`��f�=�Y>S>o>�Eپ�}���$��x�g��]y>�w�?�z�?޻f=��=��=�|���U�����Y������<�?=J#?+XT?b��?z�=?Yj#?ε>+�gM���^�������?� ,?ď�>���m�ʾ��3���?P]?u7a�d���7)���¾ս&�>�W/�-*~����oD��̈́�����������?;?��@���6��{辚���\��[�C?��>OT�>��>��)�G�g�&#��,;>Q��>�R?��>�kN?��w?�Y?-S>O;�H&��U���9��<��9>~>?�ށ?HN�?Sq?�u�>0�>r51�N5徐����� �j���~l�4�'=��C>��>� �>��>�P�=��ӽ������B�^P�=��>�A�>*~�>n�>��d>�i�<q�G?�@�>J���O��ƥ� 䂾�.���u?-h�?�]+?�I=;�BE�ڷ�����>EK�?֟�?�)?��S����=ӝ�)޶��r���>5s�>�D�>�H�=��J=T4>P��>���>��������7�<�N�x�?�E?=��ӿt�A�0�=�-��k>���8*��պƾ�˾	��>\�s�Y5��k|�����=�	X�Uǅ����A٬��� ��q�>ϫ�=O+>..ѻH����B�&���Oa�*T<�\5>��(�P�a>Z7���	��Ký�������i�=H�v���Ǿ��{?��J?�V-?��??p>fa>��]���>�U��S?*WR>)}��h����9��֭��^��gE۾�پDYe�G��:C>��:�T�>�p)>���=i��<���=�Qh=��=}`'�B��<���=�а=͢�=�J�=�M>�5>�6w?X�������4Q��Z罢�:?�8�>�{�=��ƾk@?b�>>�2������~b��-?���?�T�?H�?;ti��d�>B��O㎽�q�=�����=2>���=��2�I��>��J>���K��Y����4�?��@��??�ዿϢϿ<a/>"�8>F�>�R�*N/�\�]�"c��oT��"?%:���ʾ���>�ƿ=�ݾ��¾�>=V�7>*:i=����@[�M��=��q-=�_k=��>$�I>�G�=(��M;�=�&9=���=��S>5���I�;��=��+=���=C�b>��!>�X�>�x?nW.?��_?h�>t�^��߱��Ӻ�h��>�ή=�>��=�p>�G�>�+6?p�E?E=D?�o�>�~=;�>��>I�(��ml�׊��W��tв=���?���?O��>�X�<U8q��O"�J=����*?�*?m?s��>�<��xݿz���Z%�z��;ov׺��<�ˀ���X��U�<Z�4���E���5=���>�G�>�H�>�-I>/� >�XS>�}�>~�=��kI;=Pi<]=ѣ��z�W=�X�<�5=��;�q�*�;�<�<4��������>~���=�"+=l��=���>Q��=��>~�Y>5=��FpI>[f����`���r���Y[A��`g�у��oE�#@�t��>��i>v�ۻ�[���r�>�K�>���>���?b��?��>�n��B��c��~\վB+�ϗ�>�'>BѼ�f��6��m�W�u�پ7��>pߎ>��>~�l>�,�<#?���w=�1b5���>�|�����|&��9q��?������Ii�4Ӻ-�D?cF����=�!~?İI?�? ��>��ŅؾU:0>�H����=:��*q��g����?�'?,��>D�1�D�+[̾�k����>u$I��O�պ�� �0�q,��Է� ޱ>G>��3aо'13��O���ÑB���r��׺>�vO?�?�a�Bv����O�������[k?�g?tK�>�5?��?Xࣽ�_�����=P�n?n��?C�?8t>z5�=�>��vB�>�?_W�?��?up?9A��A�>״Z��#>�[�]�=b��=�ʁ=׃�=�a?O�?2�?ת��Q;����m��6��X�=��o=��>s��>ʈ>�>A�=#j�=]�V>�˫>!G�>��Y>kۨ>�b�>�K9�,�'�޷�>�t�>3_>�4^?��>w�=�>ɻL���ƋA>i.2=�V��o5��i��p=:�Qk�=�Q�=+�=��?}�ѿї{?|*I>_q.�-�?2����:�!�?��U>��.�8�H>�.S>�Ef>ci>��A>��~=̯T>��m>̐̾A��=�� Z(�6�3�LF��ؾ=_>�͎�q�D��f;�6�;�{U~��z���z�C{d�B~���,�/���A�?:	�:��[�R���<?�M�>�?��o��Q��옽�!�>���>uQ)�؄����q���¾ԝj?0C�?�;c>��>H�W?�?Ւ1�23�vZ�*�u�m(A�,e�U�`��፿�����
����,�_?�x?0yA?�R�<+:z>Q��?��%�Xӏ��)�>�/�'';��?<=u+�>*��*�`�~�Ӿ��þ�7��HF>��o?;%�?vY?ATV�_� �E�>h4+?�?6?�l_?s?a:?0K���"?��:>�?��?F!)?lO2?8�? �E>�9�=��n���=�c�$e��,7	�X���"�)��&�=W4�=(h0=�~�o��N��=<�=�)�<u�-�Y�F�<N��= �=�D=}¦>��]?�,�>p��>��7?�/�G8�����'/?�V;=�r���O��ߢ�Ϝ�2]>��j?��?�/Z?�d>~�A�ѢC�b�>i��>��&>þ[>s"�>�d F����=�s>��>0T�=�N�����>�	�[��c��<Z�>���>��>�����>����Љ��D�x>��#��l����8��;���8������<�>c�I?3�?���=q��T�R,_���?��8?33_?��?K�)=�����:��H�L	�Ð>b�<�����A���vy4���	��I>���zݠ��Tb>ܽ��p޾�n��J���羱9M=��VV=A� ־�3����=R$
>����� �i��y֪��/J?֗j=5u���aU�om��U�>`��>߮>��:���v���@�ﮬ��4�=*��>��:>Bn��V���}G��8��U�>�3E?�E_?�n�?�ڂ��r���B�?��Y���
�μ��?Q'�>�Y?��B>Z��=�H�������d�@�F���>{��>����G��垾0��T+%�+��>��?̫>��?v�R?��
?�`?�E*?�C?��>ؚ��j���RB&?��?q�=��Խ6�T��8��F�B��>ǁ)?H�B����>i�?0�?��&?��Q?�?2�>-� ��?@����>�Y�>@�W��b���_>��J?
��>-AY?3Ճ?��=>��5�ꢾ�����:�=g>��2?�7#?g�?Ч�>K��>�С�3,�=��>x�b?�*�?��o?�2�=��?�0>�>��=���>ʲ�>��?�3O?O�s?�J?��>�O�<�����붽��q�6}b��o�;/�9<=�v=��Nx�O[����<ꀛ;6���G�����u=�����]<Hk�>�s>5񕾔�0>��ľ9,��A>�դ�b�� ���G�:��%�=��>
?��>�#��y�=��>X�>����<(?�??� &;D�b���ھS�K���>\�A?�=�=s�l�t���$�u���f=��m?܄^?�}W��-��~]?��b?މ�1u=��������L�͏[?��?�Ԅ����>u�?8�p?տ�>˟��Ⴟ�\����b�M�e�N�R<�v�> �Ҿ�"^�/�>��?ˁ�>��>�'��.����n��B��� ?��?r��?/�?���=�`l��濒���߇���b?�D�>�־Ua?�a��f��ʛ���r�0۾'��9܇�~�.����jL������Y����=;4?\8�?��?��?3D9��~��O�.����vj�-n��&YJ�� ��_:�JbS�0'{���(�-~�,�m��?3>m�8���8����?H?+?b𽭩�>�����/�Ҿ��=
Ʈ��`�	gZ=��u�oƌ=�=��:���/��Ã��;?��> �w>m�??�PN���(�{kY��^�6h	�>V>�'�>b�>9��>��0=�_���*�S���i^�H򭻝�u>�c?��K?!pn?����"A1����M6!���*�����+�B>�>�}�>^5W���O5&�$y>��r��'�V�����	�-�}=�~2?#��>��>@(�?��?:a	��z��Bw�F!1���<�>c�h?z��>6��>��̽L� �b��>��o?�c�>[�>En�LB �̖u��壼m��>_��>��?d4�>o¿��V�B��'@��q�@�u��=Wsz?�ȑ���"���>��*?�vw=Ao˽�#9>�<�<��2���'������k'>��?�G�=��>>:	ϾO���ڎ��Iž+Z)?r9?������*��y}>�*"?ւ�>#B�>o!�?���>�$þ�d���.?w�^?�OJ?�vA?���>Z=�泽:FȽ��&���,=C��>�Z>
�l=		�=�
��G]���D=l1�=N�˼0���QR�;�d��|H</��<��3>�ۿ+�K�5Lؾ(��05򾱬�����º�:��,�)�������r�E^����T�J_b��{��So����?j��?��G�y��=���e��]���K̶>9�y��t��U��c,��1��߿��3	!�F�P� 0f�b�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >^C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾u1�<��?7�-?��>Ŏr�1�ɿc���y¤<���?0�@�}A?=�(���쾝�W=���>�	?N�?>0C1�(S�
����A�>�3�?�?F�L=پW��=	�Չe?��<��F�6޻���=A�=�=.��OhJ>Ma�>#c��QA�ܽ��4>I�>m$"�����^�W��<�]>��Խa��/Ԅ?�@\���e�г/�h'��d>=,U?'�>+3�=��,?�H�/�Ͽ��\�$sa?��?@��?�P)?�	����>,Mܾ�L?�5?oM�>֘%��	t����=��׼)&ֻ����U�(��=���>�i >m2-���RQ��_��W��=Dh �>^ÿ��"��{"�弜<D!=�.�a���D���Q�"����c��Vǽnm=���=�>>l`|>�~<>�5>hW?�n?�]�>�+}>�)�0Ȗ��aʾU@��G��w���e���a𽚪��N����ό�±�Ko���!=�D�=7R�n���8� �q�b�]�F���.?w$>p�ʾ��M��-<qpʾc���݄��᥽�-̾�1�$"n�c͟?��A?������V�N��X�����V�W?�P�ٻ��ꬾ���=����ˡ=%�>�=���� 3��~S��91?d�?�ǽ�H}��U>z�罝{='�)?��>��D<䇪>��?�'H�g�����a>vAB>�ݭ>��>�=y��� �Խoy?��Y?<�ڽ���H�>ҩ��c����[=�Q�=Z���I��N>X�,��ݔ��-����T��<HZ?��>WF9��������/I���=�*w?MI8?*:!?�"�?MLW?Ep�<!��u�|��g����=��?�Oc?��=�,|>Y �#�پ[�??�k_?<�s�㇪��EϾ��A��8���3?��q?T?X��=�[��򍖿M�E�]-g?k�v?ǰ]�ϟ�1���Z�߆�>)!�>O��>!o8��{�>�/??�)$��s��t迿1�4�Ğ?ft@V��?9��;�R���=�?r�>��S�v"Ǿ�E���ͱ��3�=e�>�͟�v��d�n/.�˽5?Gc�?$,�>�z~�w��=X����)�?%�?x���Q��<���<�l����G�|<u�=�"�vr$��J쾕27��Už�

�����n⳼u�>�@���X��>j�6�i���ϿX����ѾAGp�?[�>lý�����i�sKt�.G��H�s���>� �=6b%��Q��Cc��58O�j��=5�>�!�4��>�/��|#����!����>9Z?n��>�:��b�����?}�	����zu���O���-�?ȇ�?V�?ƙ?H�J=�$���!�3���e?b��?�n�?��>���� ="�j?B_���U`�ߎ4�YHE�}U>�"3?�B�>�-���|=>Ɋ�>Lg>�#/�w�Ŀ�ٶ�]���G��?��?�o���>d��?Hs+?xi�8���[��~�*��T,�t<A?2>ی�� �!�(0=�:Ғ���
?~0?6|�{.�e�a?��N�Z�
g�ݻW����>)���u���ף����#X�ڇ����9�S�?���?o~�?گ�<lA��HR?Wy�>#S��!ٺ��l��vV�>��>��E�H�漼�>�M���5�b��>�,�?	]�?+@?�t��1��9N,�A[�?��>��?3�>lEV>.v~>��Eb�j��>י�=�e��K�>��W?�E?
a�=z����\�ᶀ��[G���)�l�@�M�>�pR?�Z+?�:u>�G7:��ڽ�}����=�5C=d��+�W��hR=sXI��ǈ>�o�>�/>.7(��+����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�L	?���G��6G~�ۇ�'7��T�=��7?�2�,{>���>��=@vv�뽪���s�"ζ>�G�?�}�?N��>g�l?��o���B�BA0=W�>�yk?��?�!W����C>��?K��<���XW�� f?�
@j@��^?�㢿�bӿ� ���ʾ�K��J_>�A>_2m>ݖ��|0=��0��"�<Փk<��>���>C09>`&>o=>��>nn�=�ƅ�"�-�����_@��	�J�_+�������ϊ
�Qۄ��s��Z ��Cﱾk����潅�޽x=�H��V��+d>hY6? �D?�h?KF!?��ܲ>o����e��` ��?��r�=��/?&Q?��?�F<���uVh��Q�������@��R?0��=��>��>yJ�>M�h=F�>�[>=]>J>A��<��<]ۇ=;�x>�z�>��?p6�>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?�g>C�s>rg3�KA7�թO������~>�^5?�5��ϝ9�˰u���H�*(ݾ�N>n��>�<�*�����)�~���j�J�s=>~:?b~?㪽tư��9v�L��YR>#�^>t=UӬ=�L>hTa�6IȽ�I�w4&=q �=�[>�}?��+>Lv�= ��>r"��),O�L�>D�B>��*>{�??%?4�u��{#����-���w>c�>0A�>��>�%J����=���>W�d>�x��`������?�0�U>�~�e�_�,i�Z�|=�ܗ�0R�=�w�=h ��F:��(=_�~?L+��������?J��=?��0?�
>k%�+�"�����p�x�?�@ġ?)ZӾ1�?��D�>-�?�Nҽ@(:>-��>���>#���1`��>l�z��\���ڵ���?#�?�O�(��|�N������7?��߾Ph�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?��H>�đ?wjs?(��>��r��v/�;R��s"��m��=��u;���>4>�����E�Ġ��Zo���k����ǒ_>#�=�_�>�f�#:��ƕ�=/��^@��}�i��>7yr>��I>4��>�� ?3-�>���>=�p��$������K?
��?����/n�[��<���=�^��&?�I4?�3[�=�Ͼ�ۨ>~�\?���?[ [?�[�>���<���翿����ΰ�<g�K>�2�>fK�>1 ��nDK>��Ծ�/D�hn�>�ї>�����:ھ1)������G�>�f!?���>"Ȯ=-� ?��#?�Nj>�!�>YE��5���E����>8��>6J?*�~?>?SŹ��Y3�&
��"顿��[�%JN>�y?�K?�ӕ>D���������C���I��M����?�cg?x���?#0�?X�??��A?�%f>v���ؾ�r��,߀>
"?����mA�٪&�����?�C?�>�>o�����׽�Ƽ}6����[5?�\?X'?.��`�A�ľVy�<�r��"���`<��u���>jI>am����=��>V��=/�l��5��\<���=�>X��=��2�7�����,?�@b�����?�=sr�;�C���>mV>�Z��/_?ν+��Sz��M������'u]�)�?�-�?��?��ɽ��f��@<?��?��?��>�H��r�ᾒ�޾��t�@s����dZ>�'�>`$%�K� a��s���1���JȽ�������>:�>l�?
?�->L��>���#4��H�
g���c�����
!�R+"�c<���ľ��}�e��LʾgG�� �>���4q�>ִ?�G>�%k>�I�>��_=I��>�VM>r�f>,�>�Q>�D>|��=n4�<cY��NR?v���j�'�j���հ�^+B?&sd?���>qk�X���c���J?]��?�y�?S�v>�Oh�:'+��D?o��>d#����
?�:=���_�<�S������L��	c�?v�>�*ֽN�9��M��g��1
?6%?~E��WY̾��ؽ�ɱ�FKn=��?�`E?ʛS��Ve�a�\���o�R�U�]s=B^ž�u�����x�����GP��iE��ڦ��>�G?�i~?�	��B!���Jվ�g��7�'����=V��>��>#��=��>�?���E��`�˄*�~�q��>�>�Eg?�c�>߫I?��;?�SP?�L?߀�>���>����SD�>K|�;-�>�B�>F�9?ϻ-?= 0?LT?�S+?�[c>�x��������ؾC�?^�?�=?,?��?L�����ý�)��)�f�x:y�,%���7�=V
�<7b׽��q���X=��T>�X?�����8�����gk>h�7?��>w��>���+-���<u�>�
?G�>@ �~r�c��V�>���?����=��)>���=����}�Һ+Z�=����=�5��Dz;��e<���==��=�Nt��?��g,�:���;on�<]�?MH�>OI(>�}�>�%ƾ ����x��(�>�z�>���>�d?����}������'x��UN�>�*�?[��?:�E�e�=>^��s���M!��4�ݾ�ϫ��C�>;�)?��Q?�/�?O�F?��"?��L>�$�'!���q�a�|����>$!,?��>_��ѭʾ�憎�3�Ҟ?3Y?/>a����<)�H�¾��Խ�>EZ/�]-~�~���D�)��r��ņ�� ��?p��?��@�p�6��w�¾��7Z��~�C?��>nW�>M�>��)���g��%�'(;>���>�R?�X�> P?�0u?��Z?rrs>�c2��°��暿>Ԥ�X�>&�8?Y�}?���?D�y?���>A�>Ҩ<����;�;m!��d��@��.	=�k>��>f��>u8�>A �=ۘӽ>��'�p��=�_>���>!
�>n�>K�q>b=�wM?f�>������J�Ҿ�����>�$o?,{?�?�:W>���=���y�
_�>%(�?1�?U�?Fž}Ĩ=�����Ե���2��2x=6N>�k�>[=>�>F*�>�!? �B>E`��F#���c��ͽgs�>��H?��ɽ�ƿ��r��|��颾�+<�����X]�aޛ�7�J�F@�=�A��="�Q���XV��}������ƀ����=��9W�>�q�=�g>�>Fr<�����<�['=IC<Q=��m��|�<����ػ�ɉ��8>��x4�^�>=i��A�⾨��?�wJ?2G�>��u?�tF>���\>�??Ê��?:�?�4�>�ɾ+Č��Ҧ�tL��ի����������)�ڒS=|�<9�=�y>?��>�#��b=ޱ;����=}��:\"Z��k9��=b��<[�$>n��=+?B>uex?6�z����@L��\��=4?_��>_�=�t��Oi?�=�쐿XV����쾝!�?���?]G�?Y��>&���#�>���AM�4�
<��=�0�>c7>��߽ș�>�X>
ݾm��&�x�e=�?�@��2?�s��A׿Lj>��:>=�>�eR��1���^�,�^���W��f!?�-:�ə˾m�>yv�=��� Ǿ�_>= �;>��=���\����=;�x�rC=F��=��>'2B>4״=𓴽R1�=._P=��=;.S>Q2����F���I�"-=���=�ce>��%>��?#A�>~�?a�V?��>*6�����z��d��=�^� O>��k=.�'=���>��S?�a?ZOD?	�U>Z�A>~�>zl>��ć��'��宾�3�>���?���?��>{q>/����}_��<h��k���&?N%O?w�	?~2��#��]tԿ^�b�	8���z;�;�>��8=|�{��bC>��ὟH���=�3>�9�>�Г>���=:PE>Ƈ
>�;*��>ۙ�>+�=��><MV
��T�=����ց={��=��=�����+���\�i������<؂�<n�<;���	W��"�=���>/>���>=��=C����L/>������L��w�=N��,B��/d�v<~��.��;6��B>HX>�����0����?��Y>ӹ?>͇�?{.u?��>U"�*�վ�F���Ye�[$S��и=��>>'=�^|;��V`���M��zҾ���>�ߎ>���>N�l>J,�h#?��w=��(c5���>��A����4q�Z>�����i�^Tݺ6�D?/F�� ��=3!~?2�I?�?\��>)$����ؾU+0>	D����=��s)q�\����?�'?��>�$�D��챾��ݽ�<.?���=�����F���p��w��|���?�:�J�ξ��I��Ǒ�ͫ��3(I�r�����>(--?���?��A���SY�W�ܾH�����?��l?w�k>}W ?���>�5������pJ��iw>�u�?���?D[�?qz�/d�=֘н?�>b�?��?�~�?�	s?O�;�3l�>�{�>�=�Խ�d�=Ǖ>x(�=U��=�?�9? $
?A�}�T��i������z�C�O=�Db=��>>c�N>�s>�!�=� f=ЖA>΍�>�l�>V��>�A�>h��>�p��ѹ�\0?��>���>�-?�.�>=|�ý�e�ԧ۽�;s�~�y��c����Y�<��0��(9<-�����>!齿��?ތ7>�W� "!?U��ȼSSo>��=O4��J��>�G>��O>�>ߣ�>�g>N��>�j`>�FӾQ>����d!��,C�Z�R���Ѿc}z>�����	&����w��OBI�zn��ug��j�Q.��X<=��˽</H�?l����k��)�W���L�?�[�>�6?�ڌ����̯>���>�Ǎ>�J��i���Xȍ��gᾥ�?E��?=o>��>��Y?�?�@����P�S�j�x�d@��7k�I]��Ì���{����\�����]?�os?��8?�=q�>C�?�4-��p��c�>�^(��
N��Pp��)�>
ީ��+�����2���꽍�h>��l?�J�?ͩ?� *����fkl>�0?�(?�!�?S�0?]['?U@�x�2?�|�=г?�$?�8?",?�7�>K�<�8i=�hK=���=R��.q��8k��7����?��"=�d�=���
��=�� >�����G�� �=��=c6�<G�:Һ�=K�=���>�S?��>�۹>�w0?��½�9�a����H?PBW<�v�K�r���ž����#��=��a?���?��N?��!>;�8��s<��P3>���>�.H>�O<>S�>òνe�T A=~�=Y%p>�X�=���N���l}�9]��>11>�?k)>���ӟU>�J��X��8O�>5���k��&����>�9�>��(��Y�>NY8?o�?D1�<�1�U�ϼc
W�{?�K(?h@�?���?�oڽu�辄�)�eW����+>!�y=q] �L���fN���Z0�~�'��_�=[���۠�	Ob>���o޾d�n�J	J�r���M=��V=J�� ־ 4����=�"
>>���l� �S��|֪��/J?ۦj=�q��H^U�xu��P�>>��>ٮ>K�:��.w�,�@�ꪬ��#�=���>�;>,N��m�yG��3��M�>pE?*H_?EY�?���^r��C�G�������Vܼo?���>C?2�B>ׯ=x��0���d�̛F�0�>Q��>7���PG�p������>-%�d"�>�?J�>%�?3�R?�6?8�`?�j*?H3?���>�綽%(��B&?���?F�=��Խ+�T���8�dF� ��>�)?e�B����>��?_�?��&?�Q?S�?��>� ��?@����>}Z�>w�W�)a��d�_>ԫJ?t��>�AY?�Ճ?��=>1�5���}����=�=�>8�2?l8#?��?���>���>�l�����=l��>Q|b?���?\�o?�D�=cX?I!2>O�>���=>���>(?�O?&t?�OJ?p��>�C�<g�������q���J�#e;��)<�jy=s����r����T�<g"�;�*ǼK���Փ�~LA��Ay�;
<�g�>S�s>&���,�0>��ľY1����@>���o��@���:�Ϝ�=Ũ�>�?�ʕ> 
#��C�=�j�>G�>���FB(?��?�*?D;_�b���ھ�K�4�>��A? �=��l�{�����u��Mf=��m?�i^?/�W��E��PMW?�<k?ϻ���9������{C�+>�T�P?��?�[�{�>O5�?��|?�I�>�����j6��_9W����V�0;^r�>�mݾ�
i����>y� ?)�>���>�ku���׾Fw�r�Z�`��>��?�!�?@�?qn�=��i�a�ݿ�e�������U?��>O ��8��>[�&��Y��b��*?��ežC�ľ����S)�����~�M��ؐ�<H��U�*=�/-?V�?��?�f{?#���<)��W�����
d�@^&��Q1�_1�4�#��->��lp�v��o�^k����>�K��o/��~�?��?�s��q�?^g�������s)���U��4G��׹<6��P�=�ɓ=��z��_^�~���x�?O��>���>�=?�EP��X�~ N�_U�J`��`e�=8R�>ǣ>�!�>do�=G����fi�~N����@�b�>E8v>�vc?j�K?ӵn? A�3*1�����!�x0�mk����B>�]>r��>A�W�̚�U4&�>X>���r�����y����	���~=խ2?H4�>���>�J�?��?2x	�^��bx���1��+�<t$�>i?�5�>�>��Ͻ�� �n�>�m?�q�>/ϛ>pӈ�¨���x��v��)��>�ƨ>�?�q�>P����Z������~�<�
��=�Hm?/��çH���{>fB?1��<mc�<���>�t�x�%�����|4^���>��?F��=5�D>x�ƾ۾�Dm��j��� p)?�?����)��*|>��$?I��>Ԭ�>PE�?Q��>��������?4�]?1J?BB?�}�>��=��Ƚ�Z'�ت5=��>ѻZ>�)W=]��=����c��5�P�4=���=ĀƼ��½����2���oc<�n=��6>:&ۿ�yJ�\�־@��#Y�-��;/��������}�66ܽ�˭�7����x��W�ߍ;�K6W�wD]�Ű��w�t����?��?�n��i�����F�s���^�>+��ƺҽf����F��Y����N�����jR�5�e��\�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�{A?��(����,�V=���>V�	?��?>w:1�HI����MR�>9�?��?2M=��W��	�2�e?��<��F�i	޻���=2B�=<p=���!�J>3[�>�{�AMA�"ܽ~�4>Yڅ>df"����?�^�Ǎ�<��]>Xսk;�����?kh\�	�e��"0�V^����>$DU?(��>�Θ=r�,?�;H�P�Ͽh]��+a?  �?�z�?�N)?)s��-��>�aܾ�}L?��5?�>�0&��Ut���=��aŻ13徸OV���=��>�">�*�dh�էR��^�����=�8�Y�ÿy�)�Fv ��u�<�۽\焽ᔽk�˼�?6=%���Z"p�a�-�9=A��=�
4>q��>tY>e`&>�OV?@s?;;�>�dF>2����4��ܾ��u�	ʑ�u�X�!���[b����?~���پ6����5��X���~!=�5�=17R�X���� ���b�%�F���.?x$>��ʾ$�M��-<=pʾ1���*ބ��᥽c-̾��1�*"n�R͟?��A?p���i�V�V���R����ԮW?�P����ꬾ���=����g�=�$�>��=��⾢ 3��}S��/?#� ?n󛾰�T�o�E>iFW�N^~<H�1?1\�>/
��"��>��?�ـ���	�ߦX>�M>m�>�e�>���=)��@M��{!?f�P?c�f�QP龲>>]�ľ��̾���!=̔��50�wA >�/��_���,�$&�<0=o�P?���>�=�=)�����.�,�E�9>4/�?�:I?�@�>`��?�Tx?�$3>�����Vw"�@nǼUe?_8�?Ý|=�a�=���yξN'?F�F? ؼ����)纾��,�.��>�j?ц ?��=BǛ�ܻ��f�?���2?��v?�r^�[s�����X�V��=�>�\�>���>��9�Nl�>��>?<#��G��𺿿�X4�Þ?��@Z��?��;<��J��=5;?|[�>ΪO�~=ƾ�x��Ӄ����q=�!�>~����ev�����O,�؈8?٠�?n��>䔂�������=�֕��Y�?��?�}��çh<w��Vl�Lt��ZK�<ީ�=�0��^"�^����7���ƾ߻
�,����ֿ�祆>X@��.�>%>8��0��TϿ����ZоQq���?愪>RoȽ������j��Iu���G���H�"������>�I>���W쑾���	<���i��-�>_�+��A�>`s_�/����㨾�zN�-��>uQ�>$�>��������P
�?����T�ϿTߟ�T���_?���?�a�?�X?ȳ<_���}�٣n��C?_x?}L`?�LP��BT��,�%�j?�_��xU`���4�tHE��U>�"3?�B�>S�-�a�|=�>���>g>�#/�y�Ŀ�ٶ�@���Y��?��?�o���>r��?ss+?�i�8���[����*���+��<A?�2>���H�!�B0=�TҒ�¼
?U~0?{�f.��WU?��Y��]��TG���f�	p�>���]���8���{����m�E���KV�v��?^�?/��?m;�0,4���=?���>Y��d�˾����dr�>�7�>��6=�_E�j�>1-���7��Uo>Iz�?x[�?��>���ɣ�ri|<��?��>��?U;>��x>��y>�6��`��t9�>�b$>�`�;���>��x?�+?�_�=K����%Y���k�oc>�w�#��B�cG�>	qW?�K?ål>�d\����v-�U�L��ו<��������ɢ[�C��>�C�>�+>��M����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�e�?!� �t/}�V�s�����W��S]>kx,?������>Ľ>�=Yp~�t���dW�Ҡ�>���?���?C�>�r{?�l��]��н���>(�?�%?�,X=^��i�>�?l��j���x۾6C�?cS	@1�	@�F?+哿5�׿m����2 �jZƾ�e>(��=�.>�;���R�=\�!>m$4�?�ּf��=�N~>e?K>͕%>Z�>��^>O%#>�$���(��+��+b����T�]A�����} ��Tھ��ѽ�����D0Ͼ�⿽����H���_��o�i����<��=�.?��N?k@V?�(?���YN>�
��Y罣����4�=W�?��<?�5?���=��>�q�6G���
��>����>��=��>~�?�0g>SϢ��ZK>�	>̭�>|�/>oH����M=�.>���>�?�%�>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��u�T�4:>9����j�5`>�+ �~l���)��%Q>wl?+�f>:�t>�2��J7���N��~���~>��4?:���Z=��+v��.I�Q�ܾZ�M>(+�>�*�j%��5���~��j�� w=�:??|���J�����s�Pl���S>8�`>�}=V�=)�J>5h��Ƚ�I��)=z��=s�[>��?�N/>u�=�E�>)H��M�J��]�>t0H>.p,>Yj>?�!%?�
�z������K-���x>Ц�>n9�>�N>0�J�t��=p��>��c>�4�i����)�-gA��CJ>�V��>�c���S�FOw=���T�=U!�=�v�&�5�� .=�Bv?����Ԭ��R�!��S��S?Z�!?��/=��սo'.�7y����оw��?�<@��?r ߾z!?���>xp�?E굽��>��>Y	�>��Ͼ,�L�0�>�$���W�#B���N��?��?���Y���NV�\��<փ??o�Ph�>wx��Z�������u�v�#=P��>�8H?�V����O�c>��v
?�?�^�੤���ȿ5|v����>X�?���?g�m��A���@����>;��?�gY?roi>�g۾?`Z����>һ@?�R?�>�9���'���?�޶?կ�?�I>o��?Țs?hh�>��w�W/�6����J�=�L[;@e�>�o>y����cF��֓�i����j������a>Fw$=��>�D�G/���Y�=�⋽sJ����f�睷>S#q>Y�I>�X�>�� ?�`�>-��>ա=�h��<䀾����0�K?���?����2n��^�<��=G�^��&?,I4? t[���Ͼ�֨>�\?&?�[?Db�>���*>��迿�~��{��<�K>�3�>�H�>�%���EK>N�Ծ	5D�q�>�ϗ> 	���?ھ>,��a���B�>:e!?Y��>�ͮ=� ?,�#?�+j>�U�>8FE��#����E���>CA�>fG??�H?�8��rg3�S���⡿iv[�J�N>vy?�?.��>4z��Ks����;��7G�}��qn�?E$g?����?K�?̌??��A?�;f>O3�&\ؾ̫�����>,�!?K(��MA�|�%��Q�UA	?��?�h�>�=��2׽�ʼ��r��#�?�X\?r�&?I��z a�E�þ���<"&��[x����;�$k�&o>a�>O����=��>���=?`m�H�7�.nJ<�ϵ=�-�>��=�$4�u���>,?2�A������u�=��r��:D�ƪ>��L>����u�^?�=� �{����l���T�q��?���?�Y�?@��N�h�<=?��?l?9�>����#�޾����Lx��x�]��	�>E��>�p�I<徬�������^(���ZŽd����>���>A�?	H?',
>^Y�>������-����ud���c�����$�I �s	�y"ľ�؂�oP�����&t��6�>����v�>��?7�P>r�f>"��>`9K=Vш>J�6>a�I>a��>��?>��>u�>���<�h��5R?)4����'��阱��;B?1Fd?���>T)p�(�����q$?ŝ�?���?�Tx>S�g�+���?���>�����
?S�A=����y�<�!������3��������>+�ӽ�s9���L���h��	? 3?�җ���˾�y۽��	 �=Yߋ?��6?��6��xM�]�v���`��pJ�P�6���{������nm���������� ��S�=��:?�n�?P�þ�U��opǾ�Sb��f"�1�?>9�>-�>V�~>��s>�!�,���R�w(�HU�l��>D�u?���>)�I?8 <?\zP?2`L?���>"�>d����>�X�;}�>��>��8?Z�-?00?Ac?R�+?� c>�`��?����ؾ1?�?sF? ^?�g?�����ǽWQ���t��kx��/��s̀=@��<�Nٽy�u���[='�S>�X?`����8�-���Ik>��7?�~�>���>a���-��Y�<�>϶
?�F�>{ ��~r�}c�yT�>���?*���=��)>���=	}��#�Һ�U�=7�����=bF���;��<���=���=U�s�Q�����:?�;�F�<!�
?��?���>Z�>�|��!�ླ2��^�>2|�>²�>�~?�[��y�������mv����>��?���?4�ͽ$�>�D�<����۶��������*v�=&��>{ P?nI?u��?IHI?�?i._<�];��e�#\x�!�^���?q!,?��>w���ʾ��F�3�	�?�Z?�<a����;)�Đ¾��Խ��>[/��.~����iD��Ӆ�����z����?��?�A���6�y�¿���[��ܓC?1"�>Y�>c�>��)���g�%��/;>���>{R?���>	??	^j?�_?b��>�����@᭿0
ӽ�ڸJ�?��j?�Ƒ?2�?�[�>`*1>�*u���޾
�c��� <��9���t��l=�=�>���>��>���>��w>.��;����-ʌ�c�>Ǐ�>��?�.�>� �>��C>���=��E?���>쿡��q˾:���	��=�@�=�w{?��?i?#6%>N�� �_�	�˾�4�>��?MR�?���>Xخ��
�=SLL�����L�J��TM>"h�>K�>s>�ퟻ��a>���>��>@�B���� sU�<L��?8�V?�,=��̿�����ؾ$���V=*L޾hN��������ӽ��Y>�yP������c���2�������r���P<�A�ǾD,�>�e�=o,>
��=�J/;_��[�{=y��=��=G}�=7U�;���<{�6����;[��|�;9Â;�����G�Rj��M�?��D?�%?��Q?��J>7~��Y���>�`���?"
�>�͔=(���%H��Ժ��ƻ�7ᾢZ���(k�:+��{��=�=�QR>�0>�0�=�̹���=�y=k�=���<�;=|�=���='>Lg$>2�>�(>0
p?aDp��Ƒ���\�5�t�1E?��?���<Zv���H?�^�=c&�����(�so�? ��?i��?R��>z@��ٞ>yľ�̽�j���&'���s>�j�=����� >4�;m6�����a��g��?��?��.?����o ٿ�>��7>%u>+mR�q"1��}[��c�tsZ�h�!?GX;�
�̾���>�κ=.�߾8�ƾy3.=��6>f+d=}*��T\�V^�=|���<=��m=ω>{`C>���=U
�����=��J=n�=?�O>V�����9�c�-�x3=�J�=�c>�w%>�5�>�	?߉)?�-_?�x?�9h=(о�.��8��>ïν5-�>�E�=on�=���>KU?��^?� ,?�O=>�->�{�>�F�>���DJH�/>����5�>��?�/�?�F?�ϰ>�q��gL�"�[�m����5?3W?���>�l��r� T忕�u��*^�����������@�?9>&e^>�ֽpw"��*>��x>�U>�z>�ys>!��>��=���>A	>J�<�%�=g{�=Z�X�̽��r<)8�<YP
=���='�< ;�=!T����R�!��=7�R=�g����=���>�>>���>Ⱥ�=?��/K/>⾖���L��P�=�T��
-B�-d��>~���.��>6���B>�	X>�����2����?Y�Y>rw?>���?�1u?��>���վ�I��Je��rS�f��=9�>�=��y;�sZ`�/�M��|Ҿ{��>�ߎ>l�>�l>;,�#?�Z�w=���a5�C�>�|����'�l9q�@�������i��/ӺàD?F��7��="~?N�I?r�?U��>c��*�ؾv90>�H��m�=+��*q�Eh����?�'?ܖ�>S���D�)ɾ�o�[?S��;?s�|뜿h� �h��pξh��>���_�ǾMG:�G����:���0I�<�8�x�>h�A?O��?l7��Q���B�f��b�+�ĽcR4?��o?;�i>��.?�	�>��̧��ᐾp�>�!�?;b�?��?t>���=�Ŵ�ZI�>�.	?���?|��?�vs?�I?��a�>>3�;�� >�꘽r{�=u�>궜=���=�w?��
?��
?�K��$�	�������R^����<���=ހ�>�l�>E�r>�j�=ׁg=�G�=��[>M��>�ޏ>e>�1�>I�>������
�f-?��=�n�>(�.?���>���<��ݽ�Pg�(ߤ�V4P�v�*��p���ҽ�ʷ<(ڼXR�<�n���e�>���Zs�?�VJ>'�?g"��ksi��	G>��">@ν �>�->��p>M]�>��>��.>sF�>�P6>�MӾF~>����[!�:.C��R���Ѿ�_z>�����	&����މ��{4I��q���i��
j�R.���9=�V�<I�?����ѳk�-�)�����"�?N[�>�6?#⌾C%����>���>Vō>@J������Bȍ��iᾫ�?���?�d>���>d7Y?N�?�R*�6�$�CY���u���A���g�W�`� �����P�zv��/�]?;(u?>d=?�-+<�}z>��?�&��܉��z�>K�*�
9>����<���>3(���MX���;y��&�J�Q>WNn?�ւ?�&?�<���m�A)'>�:?�1?�Pt?�1?��;?�����$?�l3>bE?Wr?nN5?=�.?�
? 2>5��=����ټ'=�6��$M�ѽ�uʽ����3=�T{=�����
<~=-�<�z��ټK;��gQ�<�#:=%�=>$�=��>� W?�?�*�>q2:?��9��2���|�(�?}jg��re���Z��[�U��,D�=�Y? ը?�8R?qd�=��<��W�->��>��>	��=���>u�����j��/.=k�>��)>rHe=(�н^O���_���g�P�T>���=K	 ?� >����
>�7��B�/��>z�����������rQ�o� �z���>#�???�"<�\7����	�U��':?	�1?/�o?Ȥ�?鹿��׾��"��L:���L���c>��ཊ�!��Т�!栿1�(TB�gl>�Ѿ�b����d>3�	�J�ھmi��_I����)�=���8�4=b��rC־�y���=�^	>�"���K"��`���w���F?�\�=�m��^�W�~곾�>�b�>51�>U�/�Hn���@�����Z}=ok�>�b6>������eI������>�_D?V�`?fb�?������o���C��� �~?�����?F��>?�D>���=�4���!?d�>E��\�>e��>���ZF��Κ����<&��>��?kF!>u
?.yQ?�8?�`?.�+?�?��>�i���ӵ��A&?���?"�=��ԽX�T���8��F�M��>B�)?ӺB����>[�?z�?.�&?U�Q?K�?R�>E� ��B@�+��>_Y�>��W�Wb��w�_>S�J?���>8>Y?�ԃ?[�=>̃5�좾2۩�QO�=�>�2?�5#?]�?��>���>������=$��>�
c?�0�?h�o?ۇ�=b�?�;2>(��>���=��>���>�?�XO?�s?��J?c��>L��<F8���7��"Cs���O��Ђ;5wH<��y=���7t�(G����<] �;g��GW������D��������;w��>A;i>w+��S�=>�)��]ܐ�;2(>�N���Щ�0 ���M�]��=�;�>8S?D��>4F!���6=V��>pw�>:k��-?�2?(�?QO4=v�_���Ҿd�H�5��>b�<?0/�=p�l����uv����<<h?��R?@�w�@Z �V[?y�w?!��\(�o���O^�Y���c?2#4?^�zw�>í�?��w?���>̬��^����)���hb����:;G��>X_ ��j���>�?�y�>!P>�rֽN�־���|��8�?iB�?٥�?�4o?���=�Y�P�ٿiK���+�� \?�m�>ݧ��.�?����Ѿ{F��Y[��Xs��/���3��q┾����	�-�8~���b߽�8�=�?��v?�Nt?�c?9y�Ag�[��&|���U�nW��}�@�C�H�D��mB��o��"�܎��&��T��=w�Q���1��:�?�*?0��Q�?fĹ�Ҍ��Ǿ*��=F������=xX��DL�=9�=�X{��J:�N���{?�ګ>�k�>B9;? �5�p!���E���J��bݾ��:>��>�f�>��>�I�=������<j͵��?k�r�ӻZv>1�b?S�J?|�m?\u�۾0��k��\�"�RSW�$����]5> >Ae�>,@N�����$��k?��t����0��G���z=�'0?�>)|�>�?A?���-��'~�@<3�I��;�a�>|f?Yp�>�U�>6y齃!�c��>*+q?w��>��>������nnz���E�Ȁ�>?��>�s?��>-��q\�ے�y֐���:���=�jl?�鄾7B���i>z�??h��<a��<���><Gf����@���x�{�U5	>Wn?1F�=�GQ>Vھ�x�������X)?&�?����*���|>e"?��>�~�>��?�,�>�þ�Y(�Y�?��^?W]J?PjA?8�>�}=�;��ŒȽ	�&�-=�a�>��Y>Z n=��=�w���\�M. �HkC=d'�=�xǼTe���<�꾼�C<~��<4>��ؿzz.���þ8^�b��L{�̣�A������1���m锾��:��l�k�������k�뤌�������?�[�?� ����J�6Ҕ��V��CF�>�2��F�ƽc���t���y����ྡྷ�˾��3���V�7j�v25�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�tA?C�(������[=7�>	t	?a"?>��1�m�x���SG�>�%�?���?@�L=ϧW����F�e?4�<�"G��,ợL�=�֤=�=�N�*�J>�6�>.'�) A� *ܽ�4>�>|k ���*�^��-�<�]>�Խ	̔��Ȅ?�v\���e�ԏ/�=F��hh>LU?�e�>*\�=�,?a!H�
uϿ�Y\��Aa?
�?H��?t�(?�翾��>�ܾi9M?�6?7�>�7&�%Dt��=L�	����J�A�U�	0�=��>uC>A-�԰�zP��H���;�="�����v�'��F.��W=��<|����F��ع�Eh�2m���Td������D=��=j�>>��x>
*U>p62>�yU?��y?�{�>�?[>#���k����Ͼ���9���*�oR����3�鼧���!����������rz��� =���=�6R����_� �>�b���F���.?�t$>��ʾ��M���-<�oʾH����ڄ��ॽ�.̾i�1�1"n��̟?��A?������V�����U����?�W?�O����묾���=忱�ߞ=q$�>�=���D!3�~~S��u0?mQ?C����\����)>H� �g�=��+?��?T�\<�.�>�9%?+�#��Xk[>��3>�>S��>�	>C��0۽:�?�T?7������>�|���z���_=@>�5���W�[>%F�<���WU�.��� E�<6�R?|�>���B���Ml���S�U\=�ф?�M?��>�?�@n?ϣe=ub�,ۀ�d��d�=MJ?�jw?�4�=��=N��1���{|$?�yR?N`�<7/c�܆��r\%�;(7��� ?�nt?/%?r��<.��������B���.?I�v?2h^��f��v��&%W��*�>r��>���>I�9�V��>�>?�7#��C�� ����W4�Þ?h�@��?�\=<6���9�=u9?�<�>��O�`Dƾ2l��&s����r=P�>�=���Pv����[�,�7Y8?���?�b�>�s��.����=�ٕ�bX�?��?�{���7f<��� l�px��L��<��=�����!������7�,�ƾ7�
�Χ��e𿼴��>MX@>7�v.�>�8��2�PϿ���P]о&Oq���?~w�>��Ƚ������j��Gu�˲G�"�H������>�]�=���������L��W�9�ƥ�=��>�ׅ����>�ן�r/׾B�Ⱦ_����>�R�>�V�>�����Ӷ�^-�?�^��^տR˞��辕'm?ۧ�?\�z?g?Rм�v4�R���W��Ԓ=?�?��v?h�>ĕw�����%�j?�_��xU`���4�uHE��U>�"3?�B�>S�-�g�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�VҒ�¼
?V~0?{�f.���]?�d��Cj�M{(�0���?�&�'d�m��w����+f�J��� _���?j��?UΫ?R~$�=F=�U/?�V�>y���j���(U�<��>#	?\=+>����	�>=�0���-�Z��=���?];�?���>Ri��/��� �f=�"u?�^�>{�?�N�=h~�>�֧>������^�>YA>i#7��x�>+Yr?�=?n�=����W��bm�rtO��1�F�c�>��b?��(?l�>��n���սȔ�5�������.��=VWx�^د�H�ֽv�>���>�!�=U��ß���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��z?�����{� ��B@���>C#6?����>/6�>���=�dv����hdp��J�>Q#�?���?#}�>3in?��p�`H��^�<�!�>�m?�x?0E�;Y4��u@>@o?%A�	R��Ȕ ��pk?��
@�b@1�[?O�� �ӿ����%ܾV+Ͼ�#>~^>Ɏ9>,����=U_�=��=���=�B>���>P�?>��j>���=;�)>�0>V8���'�2'��,����<O����������d��}�$�K��_����f����������A�?����󸴽��(=*K�=xaA?a&V?�G?~P0? ��=�%>	����Tᇾ��>�M.�=��'?53U?G?; ���������	V���~��A���K?���=1)�>E�?��>{q�=\x�>M�>�[e>D]�=�II��6���]�<�r>�<�>L��>C��>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?��f>NBu>�3��I8�5�P������^|>�6?����9�k�u���H�|6ݾo�M>ѳ�>�?E�π�� ��d���i�R|=ti:?6i? ���˼���Iu����\R>T6\>�]=�Z�=��L>��c���ƽ++H��S-=x��=�]^>-�?
'>!�=�4�>����|Q�*��>��K>�5>�u@?A'?�$�Ma��������3��!>���>��>;�>{�G�U(�=���>�Bb>�C�ZY���4�@�B_Y>����R��R� �l=[5�����=Lގ=uM�z:�oK#=�.u?����Y�~��;����J���s?a)?�Q=�&�<N5 �1c��"��&=�?ں@x��?:�վ�I=��4�>�s�?������=���>L��>��Ǿ�׾Il�>D|���T�h~����?�t�?e�Ƚ�ځ�l6o���	=��6?7ѾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?T$I>���?�s?co�>�
x�YV/�d4��ύ��F�=�j[;0l�>�>�����fF��ٓ�qj��/�j�����a>d$=�>�\�>���j�=S֋�P����f����>�q> {I>LQ�>o� ?j�>���>�=����m�S���J�K?"��?���S#n�Ie�<�b�=+�^��?n44?V�]���Ͼ]Ǩ>��\?���?��Z?-T�>��v?���俿d���Eۗ<��K>��>�T�>5���`K>��Ծ+D��n�>¶�>����Nھ *�������2�>T!??g�>=v�=&� ?$?5�h>��>UE���]�E�ÿ�>3�>�5??2�?�˸��3�@���衿^q[��M>�7y?X�?D!�>?k���Z���+�� D�pp���?�?��f?|�齲P?r��?ԯ??�A?��f>f[��%پ�]��W�>4�!?��n�A�+7&����:	?�w?6��>����כֽ�a��;�)�����?�F\?}O&?�o�Ea�o¾n��<��%�̧M���;	wL�u�>�>�D����=�U>$p�=^!l���3��z<N��=Ә�>��=ء6��u���2,?1�&�&Ɓ�Y�Y=��|�b'5����>2mz>7u����Z?H��z���O��f՘��A��.�?I�?m��?���(�\���6?'��?��?*�?�ė�X'�����)��)ž-���"S>��p>ɥ=�k����Gg��0ރ�u�ʽL��A��>���>??J�C>pt�>����%*������T���[�C!�w�/�&*��:�aߦ��;�^t���¾�:j��M�>�<��jO�>�
?�\m>���>1�>s�I�߂>�S<>s7j>}�>3=O>��+>�b�=���s�ӽ�"R?�����N'�c��.��y�A?�c?m��>x�o�˃������X?���?6u�?]Ev>�3h�$C+��?0��>遀�2�
?��;=�h��Ǚ<3s��s`��`������u�>Ffؽp':�FZM�eog�k�	?A�?{g��P&;��ٽ�Ҿ�Nh>��?,?� 4��-x�eJc�*�I�m.T�����h�M��#��)h�Ya����a\��j*��W-�$G>�<?j�q?(0����_�s���w`���PX>(��>bؾ>�C�> �U>ji���(�b>\���*���B�>�r�?P��>�I?� <?�tP?0pL?���>�W�>sH��CK�>�M�;��>���>h�9?��-?M20?�t?�b+?��b>ʻ�����RkؾL?|�?cP?�?��?�Ѕ��Zý[/���i�U�y�iځ�.��=r��<�׽ڳu���S=��S>4Y?Ý���8�����dk>ك7?���>���>����-�����<.	�>x�
?�L�>����{r�eb��Q�>���?���=��)>��=ǧ���&ҺH]�=@���J�=�[����;�J�<G��=���=�t�i��%��:���;�q�<��	?�a?|�v>�>�ק�N�����ۖ>OQ�>���>�v�>	���脿!D���d����>U��?�h�?�o=M��=׸U>y���r��Np޾�.����M��> �(?4�<?�ކ?]�_?�)?]>'�a��\�j��d����?!,?�z�>)��/�ʾ�憎@�3��? P?m<a�_���>)�V�¾Y�Խ�>�P/�-*~����tD��J��J���Q��n��?���?��@�/�6�{�辈����l����C?�(�>ki�>c�>��)�s�g�p#�b;>��>��Q?�˿>T�A?��?4t]?��>'6�\ȵ����� �ټ˒�=� #?��p?]�?&mz?���>�9Y>�[O� b�.yȾ-�����߽pL��Bn<]�>���>�g�>��>5��=�kB�屄���b����=."}>`�?���>��>��D>ѡ�<�DA?2�>K6��;��:���[���>M5�?�I�?J�J?��_>��9�UrE�α&����>�s�?=U�?��Z?TG��ۣ�=�z<�6�������]�<`�*>��>�>�s>��v>{?��X>RX��W.2�K�Q�.i�«�>��P?��=�ƿȷq�'�q�	���af<G���<e�_���m[�X��=Jo��q���6��k[�|���x�����X ���{����>� �=��=J��=�"�<��ȼ"�<I�I=n�<�[=�3s��q`<Q^9���ڻ�j������Z<l�G=O7��q+˾��}?�I?#g+?�D?�ox>?>�t6�Е>�����?O"U>�N�F»��L;��Ȩ�R���ցپ�
ؾZ_d�a�����>BBK��>g3> ��=�ɍ<'��=��s=޷�=x����D=��=0�=�4�=��=}�>|�>!pq?�O���L���	M���R��2?�.�>I�=%�ľ�`V?�d�=���A]��)e�!0�?7��?��?%��>��V��۪>�׭�d;��m�<���<H��>S�=��5��̰>o�s=4���7��B�޻���? 9�?)`??˵���Ͽt�y>O�7>>7�R�Bz1��\�}�b��EZ���!?�A;�~<̾d1�>���=C;߾��ƾ��.=e�6>��b=C��\\�!��=	�z���;=�Sl=�Ӊ>��C>r�=*H�����=�SI=��=��O>i����7�#�,��23=���=d�b>W&>���>���>�?L�d?�)?�
�����B���l;>�[��20�>����6�<�E�>f�D?޹X?��:?�A�>�碼��>��V>l#>�6���0�4�q�����>.��?[�?3 &?��>�vξ����`���)@?��<?.�,?��k>�e��/ҿ%�p�?8����:*�=?��Jh˾e������Ě�=�>H<�>��>�X}>u	>{Ё>�8�>��^>(�>p�M>��=��;'����c=TFM�K(=�V�<��#�7�ݼ��늼�b��{�<΂<�B�;{�.;	��XC�=Q��>�>���>�W�=���'>����O�M����=,(���@���i���y���)�>A)�?PO>�hR>J�ý����b�?�Z>��f>�8�?:�o?� >�>(��gᾖ��ϔj�2�3����=��>�OI��;�c�Y�C�L���Ծ!��>�Վ>9�>��l>E�+�	$?�Pw=~B�Dn5�*��>������Ļ��
q��/��k蟿�i���D?lC��{�=�~?��I?��?ow�>���&gؾ�,0>}9���=���q�F𓽢�?'?�Z�>�K�h�D��Bɾ4Є<V8? :=2E`��㟿x��?���k�Ͼ�?�)Ⱦ�]���*4��6z��̉�1#Z�"�|�x�>8!p?4�?g��vt���F��{�f��=a?~�G?�G�>�l1?�]>�*g��_�%�f�Lċ>���?���?&K�?ؖ�U۽=n���v�>�2	?��?�?�Qs?1�?��W�>qN};�R >4����A�=��>[�=�i�=�\?�|
?A�
?<����	�����񾲿]��<H�=M�>�p�>o�r>�F�=ohg=϶�=O\>��>�>I�d>���>�m�>���� *��,N?\n�=lW�>��:?^i>���;8�ݽ������)�(�5����j�a��{o�����Rμv_�1��>�E���.�?Mv�>���u;-?�.�D��W.l>�>_´���>��>��4>m��>>�>@5i>O�>�>�tӾ�>���<!��1C�P�R���Ѿ�$z>rĜ�Z?&�c��My���I�t��(q��j��/��y==�ɠ�<�H�?01���tk�H�)�h?���g?�a�>�6?k���a>��~�>Z��>�{�>�G��o����ō��u����?���?�g>{/�>0�X?�?�����%�x[�z9v���A��nh��^^�����Q���J{����]?�v?2�=?Df�;׆x>�p}?.%�7�����>��*��L=���<��>3ر��+\�O�ɾ�����}��M>uCn?�˂?��?��K�
�m��'>��:?˛1?�Ot?��1?e�;?�����$?Go3>zF?�q?4N5?��.?%�
?L2>�	�=x
����'=�6���N�ѽ|~ʽ`���3=�^{=��͸� <&�=���<,��ܣټO�;%��w%�<$:={�=4�=�>�>:CG?�b�>�F�>B>N?!v��=�1�˾?N�>�%#���P�+Qw�1����澑��=�]?�1�?"vK?.�=}�@�ګ����=���>��r>`\>1b�>h��2�=�WS�<��=�|>��>���������%�H�*a�=x�>���>�>7>�j�Z>�܆�!�����>I%��x��B�}�2�|��"�����>�_9?	?��=[˼�L&&��Z�S�2?X<5?��d?L�?�pʽˣ
���P���]�٤��b�|>a�>�=$�����0V���F%�����`ͅ=�Pپ*Π�+�b>��>a޾pn�rJ���羂�L=z���T=�2���վ,�e!�=�G
>Q����� ����Ԫ��
J?B�j=�K���cU�6b����>2Ř>�֮>�)<��Nw�/p@�޼���p�=���>��:>8~��N��G��Q�X'�>��D?8�^?S_�?�E��~�q��C�� ��{�����`;?�>�?�D>�ұ=Ū��Y9���d�`EF��>g��>��s
H��M��C��G%��C�>�Y?�?>�l?n,R?�?n�`?.�*?��?��>��(V��l/&?�m�? G�=K�׽�IS�H�8��TF���>+)?�C��j�>�&?}�?'?{�Q?��?:�>B� �C�?�V��>C�>��W�;��`�]>�aJ? �>�Y?��?�a?>�4��c���)��ߞ�=�>��2?�#?�u?�y�>��>0U��L�Y=|��>4_?�<�?v�p?��=u�?"�3>@��>BÃ=��>d��>6�?H�P?�Hs?ZI?f��>���<� ���ֳ���E�@;"���;��G<�Gr=���M�r��b�(�=��;��
��2�{� C���O�d��;^Z�>qu>'����7,>9�¾\��p�<>�4��u��v���F�:�S��=��>&L?x_�>���q��=Ed�>��>x?��(?=8?zj?jG�̻a��վ�,A��ò>�`B?���=��l��ᔿ��u�@=a=�m?+_?��V��?���r\?�>p?����&/�'�����`�ȥ�2R[?�x#?@�k�a7�>��?��?��>T������[��~xX����Ņv=�>����@b�S�>��+?��>.W>�E�<0���˹x�9\���v?pD�?�+�?�ǀ?��=S�e���ؿv��������U?� �>�ݙ�b� ?����E�ݾ�X��� ����Ѿ����2�����V&����g��&���D��>�1 ?�ۃ?X��?,�p?Ǽ�Uux��gZ�Z?u�ks\�+:��|"�N�C���B��]L�Zmq�!��X����HK�=�j_�k�<��B�?t�-?��ݻߌ?G�޾X���Ͼ{=���������=�7(=8k�=��=pن�ܒ1��ľ��?��>�A>��3?��4���y\�E�x��R ��׳=���>d/�>s�>���=�3�<"�Ƽ�>��4$�2�>�u>�c?7�K?�tm?�'���1�O����� ��4���C�9>�	>F��>��R�xi�N%��a>�w5s�'�����������=��1?nO�>�ӛ>֗?�?�	
�W��ZMv��k1���6<�?�>&vg?���>g&�>U�۽�5"�E��>v+o?H��>�Ϣ>,�����E�x�U痽�:�>�>�?h�>˵�AY�OD��eǐ���:�G��=\�n?q��K�R����>v�K?p��;�!6<-!�>qd�c�!�������<�$�
>$o?9��=�%<>�oȾ�@�HF|�(~���)?��?t"��ϱ$���Z>�!(?�k ?���>��?�̛>u!��H
�L�>z�U?��G?l�G?���>i=�����ŽP�"�Gx/=PI�>��\>��A=�=Z���mN�����76=z�>؜���_���1��g���<<!0�=ͅ'>>�ۿ��J���׾Ŗ����,�������¸���(��r��yޗ�y<s�ҥ�I�0���Y��g�W*���%h��!�?b�?:Ҏ�oV������^��sQ��ջ>Av���|��ݭ�������,^��q��6"�q/P�T�h��d�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���z¤<���?0�@�pA?��(�����X=���>Mo	?��?>��0��C�7��c\�>/�?�ӊ?��K=°W���	���e?J�<��F��7߻YD�=��=_=o��k�J>Ȏ�>�c���@�v�ڽs-5>M��>c1!�~�K�^���<i/]>'ս�Ɣ�Ӆx?m=m�?g�7;b��H�l�~>LCI?<P�>�񐽃M?�	2�?rҿK�K��܃?�q�?�3�?�4?�F�=[>�'ɾ�+?� ?�΅>g\����n�t��<�8��a�q=������I�Z>@�%?#� >��^�:�پ��߾�p�=�=����ƿ�"��n#�V�_=^`�=0r����&�����Ѳ��<k)���2�qi@='��=�/>n�K>��;>�*�>9.V?��x?�R�>�Z>av��5����Ѿ8�e�q���8<��_��H8��i���<����߾X 
�h� �a���ڻ�� =�~�=�6R�_���&� �P�b��F���.?)v$>��ʾ��M�f�-<�pʾ3����Ԅ��ޥ�U-̾�1��!n�;͟?^�A?������V����Q�}���m�W?�O�ϻ�k鬾���=뽱�v�=}%�>���=|��� 3��~S�"�+?��#?$�ƾ&�"�F�M>k�r�u�t=�+?'J�>^�~�>�[?Є������X>�X>G�>Ӟ�>,�<P!��EZ��j? `?ޏ�=����ʹ�=����9������_=gV=o�W���>P)��վ�j=�kz=�+c=-yJ?j��>(��듾����m����=�h?�
h?��?N��?���?H��>'Y�$��X]4�m�z<Ye?��p?U��=j;>�n�����A�'?�3?� \=ź���t���2�����,?�Ot?�o*?�o�<�݌��6��HW=�FDh?L�v?Ok^�Gm�����	�V��*�>6p�>���>��9��n�>g�>?�#��C������^4�连?��@׌�?��:<����e�=^3?�I�>֢O�m2ƾ���{}����r=�-�>@_���Pv�����W,��k8?�?��>����5����=(ݕ��O�?��?����ms<%��>l�;����[�<�/�=�-��L!����T�7�$�ƾ�
�9���<�����>nL@U��:�>��7��⿨[Ͽ�1����оa�q�,�?�m�>�jǽ�;���gj�)u�۩G�a�H�����Gh�>]��=��彜̧��-��X�B���=Y�>�<��ʹ�>P����gž�@�������:�>���>�y�>�'�� ���zp�?� �oAԿ�n��:�ݾ�tn?u�?Kt�?C$? V���ǽ�㈾;DʽC�H?z�?=Fd?_2�=sD~�d̎�%�j?�_��xU`��4�tHE��U>�"3?�B�>R�-�`�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>q��?ss+?�i�8���[����*�B�+��<A?�2>���H�!�B0=�VҒ�¼
?U~0?{�f.�c�^?[%a���o��L-��	½7h�>�H7�B�d�'���{"��cd��ś�Hbw�-�?ǩ�?[�?���@#�q$?�,�>�K����Ǿ��<�ߦ>3��>ϧF>��x��gq>�;4:�?�>w?�?{�?��?#	�������V>��}?H԰>5��?e�>ѥ�>Ϧ!>q�¾2໎g>�
�=����1��>��A?���>�X>c��j�!��E�!�R���
��D�?Γ>�fa?j-D?��i>�#ǽ����&����	���=��mF�h�G����W��շ>g'>Y�=T�}������?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��w?�G�p����$~��n�hB����=�36?��v�>4!�>���=�w�!r���Op�RY�>��?���?���>,m?.�n���G�w��<
��>�o?
�?C)
<M�(/>55?�f�h���rf���lj?>
@V�@�tY?o]��?�2��9}龓�ƾ���=T�>>r�|>BS+�S�=�T=�����;<(�g>�א>
�5>�S>8�'>o�>��!=�}�L �����n;���O�8�"��a�yho������h>���:��Ӱ��}ӽ����ݖý��*���F��e��J�={�E?T�^?٥2?�2?i�3�.dC>���#���b{��G �%>�4?CFH??g��=r�׾��|��Ս� m����Ͼ�`�>��>^/�>�?�\�>h�����5>�%>�7�>�D�=�0ں��WF�DS(>w�>n�>�T>�C<>��>Bϴ��1��c�h��
w�e̽.�?z���N�J��1���9��ۦ��i�=Lb.?8|>���?пb����2H?���y)�ٹ+�q�>{�0?�cW?V�>����T�Y:>G��Ӧj�`>�+ �pl���)��%Q>gl?��f>"Iu>C�2��W8�oP��}�|>6�5?g���:�B�u�0�H��zܾhO>�G�>-��T�
𖿲�~���j��|=�a:?�2? ��ȕ��,�t��(����P>�Z>�`={n�=c�L>]�h�gɽ��G��%=���=ϱ[>��?��>�'=t��>�����U�ՠ�>T|t>K~i>i<?�6?�����ԽhҪ���m��)�>���>�*�>S��=y�9�<��=,��>d�X>,����U����&��rB��_�>�ӻ���`���߿=�:��P#=c 5=�ڽQ}����<�~?�~��f㈿�'�ˤ��^eD?�*?��=�E<�"������W��o �?}�@!m�?�v	�֛V�	�?�<�?}$�����=��>��>9�;�L�7�?�8ƽ-�����	��@#�V�?e�?,o0��ȋ��l�(�>bb%?��ӾPh�>wx��Z�������u�v�#=Q��>�8H?�V����O�d>��v
?�?�^�੤���ȿ5|v����>X�?���?g�m��A���@����>;��?�gY?soi>�g۾>`Z����>һ@?�R?�>�9��'���?�޶?֯�?>I>���?E�s?�g�>��w��W/�i4��������=�W;�h�>{�>T����bF�dؓ�}k���j�"��vb>b{$=��>XH�z8��P;�=I����f�J��>`q>�I>S�>� ?�b�>̧�>�t=ؐ��〾=�����K?h��?S���n����<s��=
z^��?�)4?Mc��о���>��\?���?A�Z?@h�>}��[;��࿿����a/�<1 L>��>]%�>�"��/wK>ǾԾ��D�_L�>���>;���gھ�:���@��'$�>E!?u(�>?�=@� ?��#?�tj>z/�>RE��3����E����>\��>}I?.�~??����V3��
��꡿ �[��BN>�y?�K?dЕ><���h~����C��FI�-�����?�hg?L����?g/�?��??��A?Q$f>[��wؾ86�����>��"?��"�SA���/�X7��?��?���>S�ý`�}����̀/��(�c�?w�f?��,?pz���e���ƾ\��<�� �!滉:t<\���
>�>B Q�j��=�Q�=���=?���gݽ�/�=|�c=�X�>�(�=G;&�M�ǽ�<,?�G�Nރ����=��r��tD���>TYL>����Ϊ^?m@=���{�����x�� U�1��?z��?�l�?�)��ޘh��#=?�?	?�&�>�H��v�޾���"Lw��lx�t�Q	>���>Ll�徏������=B����Ž���>2 �>m�?�� ?K�K>(�>�򗾶0'�Y�����]�%C��[7�W�-�:��qL��W�#��H4¾��}��:�>��>�
?]Mi>��z>Wy�>��R�>�O>n�}>�>��T>�d5>? >~�"<�lӽ�.R?������'�Z�辳⯾DB?̝c?���>ul��������4X?兒?�w�?w>� h�
H+�r2?8}�>ֲ��l
?�t8=�:%��X�<�o��������'��>�lֽ>:��M��cf��
?�Q?�S����̾b�ֽy�����>�h�?��5?�g7�dc���p���[���R��l�nݏ���\�����v�17��d���P����U*��Q>�9C?k��?y`l���u��i�ǅ�>�'�A#>��>���>λ�=cw�=U��Ĳ>���Y��#�?RR����>��k?���>��I?��;?MP?��L?P+�>��>�0��3�>�S�:��>3F�>��8?%�-?4�/?2�?�q*?-a>C���et���\վ�Q?b�?��?R� ?<�?ef����ν�޶��֏�h=v�Eǉ���y=�<�mݽ�
t�q�I=�bM>We?՞� �8�����*�w> �/?F	�>�M�>��h����	V5=�_�>w?�F�>'���{�Z��rS�>#j�?[=#���2=��">��=�I��xŅ�˸�=�9��T�=����ᆽ�/�;�B�=�^�=�^<!�;!k��Rް�c=�L��>��
?�>��>8v��*��ƫ��!a>7�>�{W>�#�>����9;��퀘�mRg��"�>��?BQ�?�_���=��L=c.��8�ǾSJ��i��:��=K�>��B?�>d?l��?�&?��-?��O=&�Y�o���h�|6^��?t!,?���>�����ʾ�񨿿�3�ҝ?H[?~<a�1���;)��¾%�Խ��>�[/�/~����.D��녻����}��*��?쿝?�A�d�6��x�ҿ���[��:�C?�!�>�Y�>��>]�)�x�g�d%��0;>��>PR?��>K�8?�Vb?��O?�/�>)#�[A¿Q��������?��h?��?&��?N��>|kG>B��l�ھ�鮾�.;�+���A��{�ӽ*Y>�*Q>���>{��>��=�wŽ����\�U����=�o>�?���>�l�>�V>��>��>?���>>˾Am ��ש���#��=#�s?�ԇ?N�?=#H>z����G�!���Qk�>��?*�?Fa(?���dM�=�,��O������S]>���> �>� �=Vi>A�>:�?f��>��t����N�2�v�+-	?�H?�+����Ŀ|�q��d�笖����<䎾j�d�����>X�|=�=�}�����YЧ�#�V��埾ѓ���"��]���ʼ��l/�>�s�=���=��=R�< �x��3d<R'=A_u<}r=��h�<�~<��8��潻�V��f+��t�<�6k=�S������~?lyC?;�1?�xI?�df>�>MμT:�>:)ý�?_�c>���[���:�0����ng����Ǿ�ܾ�3d��q���s>d46�[�	>]�(>��=mQ�<��=��U=��=j�n9at�<H_�=�f�=hb�=�	�=�S>�u>�el?4����8Kd�a9y��=/?���>��=
�⾯�E?|��=�z���c���$���?���?�	�?´�>�	R�7�>֎������]<`Q=TM�>	��=��4���}>T=����X:��*��6�?Qi@�U2?}OY�Կޕ�=�;>�>BAR�?/���Y�q�\��R��0"?��8��ʾ���>�ٵ=�ᾥhƾ��0= �;>�q~=q��"\��N�=��}��-;=�|=@��>�@>]��=j����{�=fN=I��=�S>#3a�9DP�L���"=fi�=�}i>�`#>IU�>��?�?�u?�B�>l�ܽ�9�{�޾_>8���x_�>�;ϻ�>>&��>HH?$�Q?t�?P)M>���=Ѫ>�W�>w��/\c�b���	�����>٦?yd�?'�?ep>O3��L��G���\c?�J?B��>T�=�U����-Y&���.�'����o��+=nr��QU�w����l�#�㽙�=dp�>C��>`�>-Sy>��9>��N>��>I�>@B�<�r�=H쌻���<���5��=Z�����<�zż}扺�&���+�y����׍;x��;�]<W��;��=C��>]#>���>�:�=���1$/>����¼L�*�=@4���B�'/d��3~�o�.��96���B>�SX>܄�c+���?�Z>��?>
��?6u?(�>��{־�P���`e�!�R�tS�=ɔ>� =�$�;��:`���M��mҾV��>xߎ><�>g�l>�,�S#?�Q�w=��Eb5�"�>}������(��9q�@������ii�ːҺʠD?�F��I��=p"~?�I?X�?���>�����ؾ�:0>�H��(�=]��*q�\i����?'?Ǘ�>����D�k�⾱���6?C>& ������`+�(�C�a>��>:&?���b���6�+ώ�G����K�7����O�>1�Q?�߰?c?������7Y����g�(<">?7Q?Mt>p	&?=��>������ ���:�Z��>�o�?���?d]�?�սZ��=lᮽ���>W�	?��?n�?��r?�;���>"{�:*s!>����=*	>=��=q��=��?9N?��	?nU��j
��,�e��'`c�hM�<�m�=?#�>�K�>��u>q��=8�V=��=J�W>���>�0�>�b>�w�>�`�>�M������<;?���=:�>��1?��r>/�^=���Q�1������AC����f���=�̽*y�<㑏��ڴ��7�w��>���pA�?�<�>wP⾠�/?����?ҽ�d[>-�L>������>(<6>�f>k{�>龑>a�=>W��>0V>�FӾw>����d!��,C�[�R���Ѿ$}z>Ȝ���	&���Cw��BI��n��~g��j�V.��Z<=�:ν<1H�?������k���)�����?�[�>�6?�ڌ��
��a�>���>�Ǎ>K��i���[ȍ�hᾙ�?9��?�6c>��>��W?�?�X1�B�2���Z�,�u��)A�e���`��ۍ�c����
��ѿ�?�_?��x?pA?���<�Bz>p��?,�%��Ϗ��-�>�/��3;��v:=p �>�/���`�ϤӾ��þt��F>��o?�?�S?��U��0n���%>��:?�y1?5Yt?`
2?�W;?�w�Z�$?��2>{?�G?^35?��.?��
?��1>��=4���j"=����芾sҽ��ǽa��q�8=t�u=�]��l�<�%=�S�<��켊�ټש#;W?���ʪ<m<="D�=؎�=�4�>P�b?���>��><@O?��0���2��Tj��%?����5P���"�{�Ӿ�꾇g>4J?Չ�?�#b?��
>��A��.=�G�>�\�><{>~l">���>8���v���0=�>L�>�V6=����r���e���j����=��>���>>�[>�(|�ĳ�=&mr�ZH��PG>E�s�Ч��p���G��!�C�ս{��>�zK?u7?1�%< �۾����VS^��@?��S?֫\?�l�?�A��%־��&��-���p����=x�\>Ş�PD��#�*�2�f���{=>0㴾۠� _b>ĸ�Fu޾�n��J�C��M=�����U=& �־8�A��=s"
>A���X� �A���ت�*J?��j=�l��iYU��_����>Ƙ>kݮ>��:�9�v�l@�����9+�= ��>��:>P(�����_�G�8:��?�>V>E?Z_?�h�?�܂���r���B�M����p��$t̼D�?Wc�>��?ӬB>��=�n�����d�I�F�<�>Ѥ�>*����G����x/����$��> !?�>��?�R?��
?	�`?p:*?I?�>*뷽˥��}A&?��?��=]�Խi�T��8��F�r��>�~)?�B�D��>0�?`�?G�&?�Q?��?m�>&� ��@@�哕>V�>��W��a��=�_>�J?0��>�AY?�Ճ?�>>}5�B�
����=�
>*�2?8#?!�?0��>T��>�}��Yف=�6�>i&c?c�?�o?	��=��?�d1>5r�>�K�=�6�>X`�>F�?�AO?3�s?�J?3��>LT�<,��s��{t�(T�kU�;�N<p�w=tW�)�t�~��^�<���;���0]��UG��A�N8��R��;�%�>6�r>7Ɩ�Uc(>�¾�߅���8>Xȼ����c��؏=��=�[>��?��>���N��=t�>���>��g<&?AQ?��?�	��Ajc��T˾{>*����>��B?tg�=�n�ᖿ+�w�]eR=��n?�xa?~]�U����\?Q$k?N����l,�����b1d�;߾�`?��"?Q P�=��>�Y�?rV?ϫ�>����Z����e��V \����Y�<O��>8o ���_��>.�4?)�>PN>���;֏�J`r��i���m?�U�?�?�{?�S�=�d�?�׿���[�����R?֔�>,.{���	?�H��""��s���@V��ٕƾ�>���⧾�K�������X������j���
>��)?�=�?�ˁ?��s?�P��?a�ْK��b��s�L��־��%��E�/<��H���u����_�P̗�۬�=�E�!�.��d�?��&?��D��[$?uNʾ$�l�ؘ̾��q������,�*>�ȃ=O��=l�=|r��R �QVv�#T?i��>�t7>-�8?E�B�(�"��YU�<e�5�꾸->v�O>7�>:�?�4>^�2=���&̾�|�R��=�-v>�tc?�K?��n?�A�/1�v{��%�!��u1�⋨��(B>h'>ڣ�>�~W���<'&��T>��s�a	������	���=u�2?�]�>�؜>�M�?|�?	��+����w��{1�I!�<��>�i?@�>R݆>�н� �R��>%m?�E�>Z��>>,���S!�6z����TK�>�M�>�� ?"K>X9 �В[����D��N�9�7��=��i?�C��
�U�Z߄> �O?��<��<�&�>�n�y� ��F���t.�C�
>��?�v�=)-?>�ƾ���B�{��ቾ�?)?�M?������)�Чq>�� ?h|�>f�>:��?-��>�P��8�
?��]?��K?��C?���>��<%B���jŽ4)#�&!B=♎>��`>� S=��=��
�l�`�� �cV\=5��=�`�qx��h��cݼS��<��=sY%>O=ۿ�H�CMԾ����<��9
�K4��9e۽4@��]������e��c.x� ��h�4�{~_�>an�������]����?��?V�����o�|�����������>�u�R�W�J���b��,c��W%�	Ĵ��"��2R��_f�g|_�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@wyA?�(�R����W=_��>׌	?�?>F<1��I�f��:7�>�4�?�?0[M=�W��p	��e? <q G�U޻��=k�=�=C����J><g�>u���A��ܽ��4>;Յ>n�"����^�)T�<$�]>ս�0��T�z?jGU���]�<�0�����<>��Y?�x>��ν�2?��?��׿|P`���~?D�?���?*�&?� ���;>��־'�?o�?�u�>,	� �v�Yn���R����=U�1���U��-2>�(?�~�>�TQ�G�����ݾ���M��=�w��#¿)�"�G����=hZ&�`�½pU���d�ǡ��	#>�,�潴�g=y��=H�'>��l>D�@>��v>�<Z?.�|?m�>eX>���w����˾p�ý��<���I���T�	���������p�� *��&�~\��� =��=�6R�i���9� �a�b�D�F���.?�v$>}�ʾ��M�%�-<�pʾ3���+ل�)ॽ�-̾!�1�+"n�Y͟?��A?������V�H���W�d���a�W? P����Qꬾ���=Ա���=�$�>$��=T��� 3��~S��g0?"�?+���aL����'>�� �d�=�+?�9?$�d<�\�>��"?�V0�YNܽ�W`>�W:>p�>N)�>��>ot��1ڽE?E0V?����휾 4�>�9����o�_=�>��*�<BԼ��X>AXE<Ua���!����Bܘ<!�L?4T�>���_<ľ$/��z��@x
>?�C?���>�|�?��p?�>���Ȃ�� .�� �<��S?o�c?,��=d�>��ƾc���� ?��=?��=e7��W���L6�
�!�At6?�Wk?0!?='�Y̒�����ǭN��E?�v?�^�Zm��@��|TX�u��>� �>�R�>�!;����>�<?Q�$�����������2�TW�?��@h��?�(<����=�� ?l��>�kJ�����c��/w��-�W=��>�I����v�� �>� �l ;?���?%�>�7����D��=Е�,Y�?��?�`���m<���(l�Ao�����<�w�=3��!�9����7���ƾ0�
�k���9�����>!T@s
齈'�>`8�y+�VϿg���^о3=q�޿?K��>�ǽ�`����j�99u�k�G�Y�H��t��L��>RN>�����:�{�o�:���y����>�p��5�>G�S�ڭ���柾���;:?�>s�>ap�>�ڤ�
����r�?Y����οM۞���1ZX?���?[��?<�?U�g<��o�Ӟ���&��E?��r?	�Z?�����X�k�4�$�j?�_��vU`��4�rHE��U>�"3?�B�>M�-�]�|=�>���> g>�#/�x�Ŀ�ٶ�@���Y��?��?�o���>q��?qs+?�i�8���[����*���+��<A?�2>���G�!�?0=�SҒ���
?S~0?{�g.��^_?:a�8�o��-���Žj��>y�1���_������ ��e�t盿L�w����?��?Aղ?�����"�'�$??t�>Z����/Ⱦ��<S6�>v��>�8H>�7o��t>���:���	>���?EB�?,�?펿
覿,�>�}?_�>���?�M�=��>��>�y׾��M����>�G>,�$��?�x?��(?��<=K��w���r�H>�x�˾N�N�`:�>�+K?v?��>�+=�PD���#�yX�����ޡ��u���W �١��c(�>��">��=Z���&���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�}�	?�9���&����n�����x�]�T>{�'?18�{4�>��>��=ay���� i`���>��?���?��>
jx?��{�Dh��!�@P�>CH?��?���<���ѫj=nV?�`�_؊�X;��W�?��@@�@ȁI?4��M�߿���mp
�W����mu<-�q>���=��彷Y1>D�<%'=a3�<خU>HY�>�PD>N�0>�cY>��/>Z&s=�O��g�#�����y ���KL��h��c��:��W�f�S�#" �\Ͼӷ������μSH��Cs6�|����<\��=r�E?F�Z?��F?�$?y�����)>%v �]gF��U��� ���)>j�?$cD?I?��>_�����}�/}��OE��/�Ǿ b�>t,p>�j?�$?�!�>�-w����>7�d>�%�>��>���=�x<e�=�k2>=֖>a�>M��>�C<>��>Eϴ��1��j�h��
w�h̽0�?}���R�J��1���9��֦���h�=Ib.?|>���?пe����2H?$���y)��+���>z�0?�cW?/�>��O�T�<:>=����j�+`>�+ �vl���)��%Q>rl?��f>0�z>�.�r�7���L�8!��kMz>�Y1?��ʾH��x�[�H�?�ݾ_�P>�M�>�?���?�����un��Ҧr�*7�=V;?a?�����ꦾ��d�T֚�BAB>�8j>��^=ѫ=J&G>�q��˽�CA�1�/=��=��L>y?^-)> ?�=�>�"����O��֬>"EH>��2>��??�Y&?�_�F����ކ�b 1��z>���>�V�>�s>��I��i�=�b�>�Dc>�g��䌽��gO?�,)Y>�����U��c�{/u=�X���[�=MF�=:���6@9�Ł!=ǖ~?U���㈿�뾸h��lD?�*?���=�pF<�"� ��J����?J�@&m�?*�	�z�V��?]@�?������=�|�>A֫>Uξ��L�T�?ƽ�Ƣ�E�	��-#�sS�?��?��/�Aʋ�
l��1>�^%?��ӾPh�>yx��Z�������u�s�#=R��>�8H?�V����O�d>��v
?�?�^�੤���ȿ5|v����>X�?���?g�m��A���@����>;��?�gY?soi>�g۾>`Z����>һ@?�R?�>�9���'���?�޶?֯�?��H>Y��?��s?�
�>��t�k/�/9���e����=T�I;+��>�>�W��MF�_Г��|����j�����ea>u�"=:��>}�����~�=�$��Z��h�䁷>(8q>h�I>e�>� ?�4�>��>�=7����Ԁ�FŖ�m�K?�?p��B'n����<÷�=ב^�?(4?Fe�0о���>'�\?���?#�Z?�d�>���=E��a�H�����<�$L>V*�>��>���A�K>��Ծ�zD���>��>+���3ھ�-��c!���G�>�R!?�>�>[�=I� ?��#?��h>0�>93E��&�� �E�<��>���>�?�?��?�>��}^3�70��M��i�[�A�M>�2y?��?쀖>yT��3F����-�XbA�/ϔ�Ji�?g?���&0?�"�?[o??ثA?�\f>�J�A�ؾ�Ѳ�$��>�!?���El@��$�+�M�4��>�U?1��>�����vν ��|
/�[�	���?��g?��:?�Pپhn`�r�¾���<!Gʺ'�#:�=��9�ͣ=Oh>�B�=�`�=��T>�
>�[��u���a'���Y<�ԍ>��]>�~.��f/��<,?�XH�z؃�
�=)�r�YuD��>}xL>����r�^?�=�~�{�T���z���:U����?Q��?�q�?B"���h��"=?S�?�?	�>X����޾�ྗAw��`x�f�;,>$��>�Ak�e���������A��|�Ž��� �>�b�>��?t� ?�5>�-�>4��+�:���;�ˇ]����Q1��*���ˍ���H�T��?GȾ�'j��2�>�zu�g��>1?)py>�v>3(�>�'�<�w�>�K>@zu>�>��P>q�:>���=\�8�21��R?fN���V'�i�����P�B?��b?8k�>�m�����b���&?��??��?Fy>ߵg��~+�;'?k'�>�~�C
?&�/=��7�6�{<Co���n�#������>��ս�3:��1M�g�#�
?�m?\���g8;��ؽ	�̾�>�&�?�>?.E/�3�U���h�SOj�-�F��m=�x��@��w����l����W�����yj#���t>}cK?3�?�Ջ���R�5p�I�d�$�W<h>+t�> w�>*0>�M>��Y/�2�`��9�=L��)�>Ђ?T�>�R>?�<8?�f?�X?
�~>b҅>⮐�P��>�8��<�>���>:�#?�&?�o,?-�?�|.?��I>-IQ�*����CѾ1�?�o"?�( ?>�?���>-F�����ǽh��_fr��i�<H�8���-�5J(<�8>�^>�X?����8�Y�����j>M~7?8}�>���>���\,���X�<;�>ݷ
?�B�> �A�r�>d��R�>	��?@�4�=H�)>#��=_H���κgO�=����|�=N����;��<,��=�=��r��o��
9�:z�;�\�<VX?��?��_>$^�>,��j^�D_����w>�*�>��>��>綾�������%�v�bԍ>6�?��?Cʘ�.ȼ=�6>�8��ˍ����߾����I�>��?-LK?:Ԏ?O�^?Iq7?y�1>�� �o��� Ob��䘾�E?$!,?m��>���ͳʾA���3���?�Z?�<a�1��_<)�T�¾;�Խ��>U[/��.~�x���D��������K{�� ��?���?�A�;�6�6w�x���z\����C?#�>�X�>��>�)��g��$�1;>��>MR?��>��C?h�q?tLZ?��>�|
��۷������l�LBv=A�"?[r?޸�?��?��>Lv6>�$k�tZž��PD�WDƽ^l����q;R�Y>��?>T��>�К>�%�=<zT�����1D�u��=�%>b#?t��>�k�>��8>�2:=�uA?%��>9���b=�2t��ٞ4��͊>�A�?���?��4?�G>,�v&:�̑%�w��>q͟?9�?ѕW?�>��L�=,�#�觾�V��3_>v�\>�o�>A4>F��>�g.>T{)?�#�>U6:�����]Q���e=���>}E?�Q>�Xƿ��r�\zu����x�P<cۏ�I^f�|v���-X���=a������J��4�Y�������Q����I��4�z����>z�=Co�=@��=Z��<iPμc��<�G=��<��=&�p�)eg<�a=��_ۻ쁅�b#��?G<�II=�r����ɾ�~?r�H?`1*?ѐD?!zr>��>�]�9��>�)���?�'[>�^>�����4X>��Ƭ�9����[ؾH0ؾ��e�l���p�>[J��/>�t1>���=��Q<,=�=q�u=�F�=k^����
=S��=��=�='�=�>�>�o?�Ys��v���(S��3�-&?���>b�)=��@?/��=7�����Ŀ��
�ns�?���?���?e�>6�X�1�>\��������=^؄�rǬ>4�>O���a��>�*>�����������?�@�JQ?%y�	�տ-�=�8>?>ظR��m1�&�\�Pb���Y�w�!?B;�f.̾B�>*�=�p߾�7ƾ��1=҄7>jd=���J\����=3ez��==0�o=r��>S�C>ϰ�=M㮽���=� K=�Z�=�9P>����3�8���.�ML2=�8�=��b>�9%>1U�>!�>�?z�L?]t�>e<���㾨Mξ�v>�����>K >=�'9>��>��;?e�6?��4?�4�>�~׼�;�>S�A>9�4������9��"¾�2?<��? 2�?�>?Ǭ�>6ľQ�0��
e� ｦ�"?�,?z��>A>]�����i�W�Li�t��R�>۩���%��4>Z�;�O*��r���J>Gּ>R�>�U>g>�B�=�l>�ӛ> O!>�]�=*�=yq�=b�ȼI5:=��d=5���<r�<Ȩ+����<݊�RH��]<�W�nB�G��<�/�=X��=�'�>��>���>qܗ=ռ����.>2��P#M�.�=�	��'B���c��z}�r�.��E5�n.A>�S>s���%��1�?x�[>��?>��?�`u?$�!>��H<־;���h�a�JS��G�=��>��<���:���_��N��Ӿ(��>��>5�>�l>2	,��#?�&�w=�⾤b5�t�>���c���%��5q�k>��H����i�Lܺ"�D?hF����=$"~?��I?��?��>���P�ؾ9+0>0A��Z=+��)q��i��"�?�'?��>��g�D�ٞ��wQ=d�"?�jJ>�������\�R��ç���0?3��蕾\�8��c��eb��K5=�X�Q���>Qcr?�(�?�1���9����Z�9��z�Y���?��n?�O>���>#M�>v�1�w���wR���L>4��?x�?���?k��̤�=�K��Wu�>��	?�ǖ?��?��q?\?���>���T�>�*��t�=�>�g�=���=�?#
?T�?Y���'	��m���G�a�9�=bП=a��>�t�>y�p>D �=��j=�S�=��Y>�Ν>N]�>(Eg>�>Ċ>c����H�u�I?��=�I�>רG?�rn>������7���G��.C`������Ի�آ�tG=������
�&ý�m�>N��z�?���>�:
�<?��f� �c�>���=2@����>�i>ü{>���>z"�>�`Q>��>̥>OӾ��>j���]!��)C�<�R�*�Ѿ�Yz>���A&�ԝ��p��;CI�br��Yh�Fj�x/��(;=�5i�<�I�?G����k��)���/�?[�>Y6?B،�>̈��>,��>č>�M�������Ǎ�k���?��?)sc>C	�>
�W?��?GD0��2� kZ�`u�v(A��e���`���������gv
��y��a�_?�x?jA?�M�<|z>ߌ�?��%��폾�ފ>��.���:�Ǡ9=�T�>3���`�i_Ӿʶþ���n�E>
^o?g"�?2{?�BV��,k�)'>ñ:?*�1?�wt?C�1?p2;?]C�8o$?a2>n�?E^?M�4?��.?j�
?�$2>��==~��p""=~b���ӊ�Zѽ�ʽ@���5=�u{=�q�<G�=8 �<�X�t%ݼ���:���L��<H=>=!|�=$(�=�0�>?V?��>F��>��@?	
��7�R;��^n?��,;@Љ��g{��ê��P
>wGd?�b�?TU?�J>מ<�ln9��>��w>�}>)�f>Br�>����"�K4V=��>$�%>��k=J%��pΊ����cj�!f�=�>Q��>X�M>@ے���=pԅ��*��4�=�,V��޾�����Z�0,,���d��;�>�E?�#?}=��	�2���^���/?��V?1�R?@��?�7��5о�[%��^�W�S�o��=�+�>d���!���U�����I�S�~�	>���6_���R>��mnо��~���H�ԕ̾V:�=�L��~�=�������5�26=���=)�ξ�J ��R��r���5:S?�>=�Eھ�3u��\;U�>X1�>�	�>5�j;��H���M����ӷb=�@�>��>�� ����Z�A�����>aC?uK>?�#�?+��+���zz>�@񩾄������$?o��>�B�>꣚>�Q>b����2$���O���,�$3�>9I�>���M�2��a���)⾝� ���`>;?e�>��?��K?��>�<??��?��>g�n�f[��R�-?N��?\���܀ƽ;E���c���>1�N?�Oᾩ�>�?�o�>(�Z?��$?��> ū<`��we�����>׬�>����������mn?U J>ML	?굈?*��> �N��T�r��x|�>L�^>p�	?n?�i>WW�>v_�>5X����="X�>��W?xp?-fr?6[��?���=���>�	�=��=�R�>���>��:?�*v?,�J?�;?Eݶ<��#������彃��7�𵄼��7=��+���,��M���/�=d�=�n�<�I��=��D����^>�1�>�Sv>�Ε��
8>O����ƍ�~e=>�l��>���?���o4���=>f?��>#{'���=�j�>���>f��\1'?�}?��?5�;G1b�! ھ�HH���>qHA?��=��k��u�Ηa=n?J^?�!W�[;��X�a?ֈ^?C��r;�Ez���zb�͓���*H?�=?�C�9�>�?0!q?:�?gBl��Lk�U�����a�o-\����=�ϛ>���Ee�Ǚ>w07?�D�>Ja>�.�=?�ݾ|�t�5t��r�?���?Z*�?gI�?޸4>q�p�u�޿o�4���D�a?Z��>�瘾�%?�rź����%Ϟ�L��6��������t�������0������Ž��N==#?'�?��h?k�b?�>�bqi�#�b��*z��dG�@u��-�=<E���>��B�t�l�R�kP�ə��b��	�Ӿm�:����?�!?[�X���?�*����x�=F�)�>�VQ������>��վu��<Hd>}Mg���U�r���5?=z+?t��>n�=?��l���k�a�%�B�+�վ^�u>��>�>F}>�W;��/�
o��b���tо�
ԉ> �_?6�&?H�o?�օ=h�C�ë��U�"�<�~p��3p>m��>;��>�-B=Ԝ>��2��rV���N�lZ�|ׇ�6�����=�I?j�>}�=1�?`2?�a8���ľ���<�O�}���>��x?��;>uU;�I$>&��&��>��l?n��>L�>͂��rI!�N�{�o�ʽ� �>�ʭ>P��>)�o>�,��\��j��R}���9���=Ҭh?|���U�`��ޅ>�R?�E�:PJ<L��>��v�w�!����ӛ'��>d?�˪=�;>��žI$��{�+9���J)?�?j����@+�Z~>�
"?¹�>�r�>AD�? ڜ>�+þz�p�$?�C_?�J?Y�@?*t�>d=�Τ���ǽ��&�(=ON�>v�Z>�Sy=a��=�&��4\������G=�Y�= ��l���|l<���Y3S<<m	=5>4gۿ�bK��&پ�����N�	��ވ������߇�aF	��@��i���wv�_3���&��vU�6rc��w��];m��t�?T>�?lK��Of�����m|�����ʡ�>*r�߱����g��������0謾yZ!�D�O��Gi�6�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��6�"���8�� >_C�<-����뾭����οA�����^?���>��/��p��>ߥ�>�X>�Hq>����螾}1�<��?7�-?��>Ŏr�1�ɿc���¤<���?0�@�=A?�(������U=���>��	?±@>s�1�;�����X-�>�*�?�؊?�,L=��W�N]�Ae?>�<�5F�M���=�c�=��=���5K>�Z�> ��FB�X]��5>��>#"��,�a�]�C�<��\>!�ҽF���5Մ?&{\��f���/��T��U>��T?�*�>t:�=��,?X7H�a}Ͽ�\��*a?�0�?���?#�(?9ۿ��ؚ>��ܾ��M?]D6?���>�d&��t���=:6�����z���&V�v��=S��>M�>��,�܋���O�SI��>��=�/��Ϳт'�8�-�p��;��_>�$�e+���o]�����K�(�L��Y��=�����$>ܰ>�/~>��>�!m>�O[?��f?�
?ϝ�>��j6�m8�P�=��c=��D���'���%�C�0�$�ྎ]�R�C�  .��X��=�8
�=2R����� �U�b�ɈF�+�.?�>$>��ʾ��M�"�(<�Sʾͪ�����?��z/̾W�1��)n��ϟ?��A?��e�V�x�����۸�ݰW?-$�}����%i�=2����c=��>�٢=V���3�uS���+?-$?�;$�+��g>�=S�2'�<!'?*!?u:����>��?�J��)$�`�>ĝ�>���>�&?Ie�=0�����(�^_%?B�X?��-�$Lm��9�>�F�j^����=e_\>��8��g�=���>�G��<:��\���;��r=T�V?�G�>]�(�m�[���p�\E=}�v?ɂ?C��>jOj?�oB?��<�����T�_�	��S}=AW?�i?�I>*���Q�ξ���F5?�e?�EP>J�i��
�:�/����ӫ?�So?$?7�ü�`}�o���F����5?��v?s^�ws�����E�V�c=�>�[�>���>��9��k�>�>?�#��G�� ���uY4�%Þ?��@���?e�;< �D��=�;?p\�>��O��>ƾ�z��������q=�"�>����|ev����R,�f�8?ܠ�?���>������+>_I��_��?���?����7p��3���&6�D��l�r��T�;�{�<�N���Z���F>�ii����p�����W�>?k@;(����>|0�w<࿈1ٿ[ɜ�t�������%?ӥb>�5�%M�$��� c��&B��B�V4(��V�>�&�=+j������D��q?�F�=�Y?ϛ5�ȴ�>����������s̽�i>`Te>�s7>S{�!��5V�?� ��^߿�J����㾸�`?Q�?�D�?)?Ɂ(= Ծ0~��1��� U?�R?'�m?���<��Q�ǹ)�#�j?�_��uU`��4�pHE��U>�"3?�B�>R�-��|=�>���>g>�#/�x�Ŀ�ٶ�;���Y��?��?�o���>p��?rs+?�i�8���[����*��+��<A?�2>	���I�!�>0=�OҒ���
?S~0?{�g.�\�_?�a�H�p���-�}�ƽ�ۡ>.�0��e\��K������Xe�
���@y����?I^�?`�?ݵ�� #�p6%?�>_����8Ǿ'�<���>�(�>$*N>	H_���u>����:��h	>���?�~�?bj?���������U>�}?�$�>8��?���=���>��=�a��c�H�
�%>�z�=6[L���?�$M?���>��=74�0T/���F���Q���e%C�~O�>��`?ML?g�a>�H��	t1�) ��Cǽ��0�B�輟�?�`�,�W�g�3>��@>Z�>�E�PxҾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�c��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?HQo���h�B>��?"������L��f?�
@u@a�^?*n|ݿW���3꾑��-7�<�>��>W�����=2kZ=~ܫ������O=�}>D\�>o��>�|>��7>��e>`���/i&�]К��l���J�/����/ﾊ`B��_˾�BQ����� ���[���<���ƻ��;�!�D��Ψ�8R�&�=��S?��J?E|u?��?=G�t�>٬��`V<��>��2�=�>��,?�dP?El/?�W=V�����`�z�{��j��̗����>�M>߯�>�|�> �>L��;��d>��?>#́>��>f$=�"���\<��l>���>Ak�>뜺>%ml>�W�=�����髿T�y��oM�ך"<٨?�����T0��<���پF��J�$=�?P�>ӂ���:̿L9��;wH?����$��_L���D>�0?G�L?��=�?b�
͍���=p7 �[�H��b>N�ؽ ����5,�lY1>�	?
8�>�h4>>�e�1_=�m8�����F�>�qY?�n��������z��Rx����=<�J>���=��3��5�����ZS���=�B>?�{�>��X�*+���ˣ������ �=�:>�-m�4`!>���<[Ě����a������*�M=��'>f?�>��=�z�>�ډ�?E7����>��_>��%>L�C?�c ?ώ黟9��H�h�E%�\�e>EI�>��>��><�>�aK�=�?�>�a>���Ȥ��r��:�,��#X>.���y�z�颛�i�|=�썽���=��l=�k��A>�U>=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾOh�>yx��Z�������u�]�#=U��>�8H?�V����O�m>��v
?�?�^�ߩ����ȿ2|v����>S�?���?g�m��A���@����>:��?�gY?{oi>�g۾<`Z����>λ@?�R?�>�9�n�'���?�޶?ԯ�?yg�>Q�?�]?�!�>��=�?�i���=$��4��<��^>KNE>���>$���G��6{��AP��;f��t��v�>8-=:��>%L�;뾵�1>hk>��.�$��?t�>!�5>���>�� ?o:	?�o�>�I,>#+�;a
��l�?���K?���?r��M2n�r��<Ut�=�_�l?�N4?��[���Ͼ,ڨ>�\?�ǀ?�Z?t]�>���?��*ٿ��v��-h�<��K>��>�>�>����gK>2�Ծ?KD��>���>)"���Mھ ��Y왻�-�>[S!?&��>�=| ?*#$?��b>���>2B��K���iF�}y�>+��>�
?6�?~�?E���S0��M��ʚ���[�jO>v�x?dX?'K�>�����板~ƼL��xJ��/�?�Nk?���Ob?_U�?^�>???r�W>�u���Ͼ#~��y{�>q(?���<C�<���O��Z��_?}�>��>��=䑱<
l��u7�2l���5?]�t?�?A���[�r�սt��<<���`|$���7�v�<��y>�[>�-i<��>�.>>���=N���������)�*�'>�(�>��I>[��<��)��<,?^]F�hჾ��=K�r�RyD���>�UL>T���C�^?k>=��{�|��^w��a�T�H�?��?o�?x����h��=?\�?�?|#�>jD���a޾���rw��jx��l�{�>���>�=i��#��������A��a�Ž7bƽ�X�>K��>X�?��>��>A��>��ξ�&��'��}�(��%=��T
�1`(�y�,��+��sm�u��i�Ⱦe�����>�'��W?��?j��>�l�>fa�>A�)�%�>*N�>��>���>I��>q��>	��=�Q,>����_?R?V���'����e���B?�d?���><�e�q�����P?�`�?���?ɺv>=bh�$+�(?�m�>���OT
?�h:=� �tr�<�趾��i�����>{׽Y:��VM�]f���
?�?�6��_7̾Iս�͟��i}=]s�?/?��2��S�1\g�c:�2ka�ӣ¼��4����� .���9�|��v2����x�y�/��Fѽi:?G��?V&�)[�ܿ��Y���*�e?>���>�H�>�t>���=���#�=�i���6������l�>�Ok?�>\G?�5?��T?�P?{��>&r�>nu��ܞ?�/K=ci�>��>)�!?�t'?_!?;l?AH?�
�>xνc��[�̾q�?:[?�?��	?/|?�����޾�4�(=�����dQ�A(=9��<RTý����;�<�G�;�E>?���12����O�}>R:?j`�>���>�����Ɠ��C%=D��>x?�	�>�� �i�p�h2���>��?Q!��s�<�&>9�=�C��d6;�x�=T�߼�w�=�9��,���D<���=j �=��1<%ޔ���:�t�<9��;vl�>N�?k��>�7�>3 ��(� �Y��K�=�HY>'S>��>h7پz�������g�˄y>�t�?�p�?�g=Y�=X!�=#���R������߽��4�<��?�$#?�2T?;��?��=?�m#?t�>%0�C���b�������?>5+?��i>�[�,����
������?#��>Dh���<T�a���������w���5���|�򆧿t�d�兾O���H�a��?!�?y�<�z2��?�������Ⱦ��O?\�>�Y?�#�>${�A?C�{�C��Ћ>,��>�<-?��>d�S?E�V?�<?�C�>k:��E��1������*Ԇ=�4*?��?W�?{��? U�>N�&=_���g��*d��<�L�����Um���{>�YN>#�>BT�>t�>"�T=,�k��,C����L�+>.�1>���>q��>]\�>��>!^���J?1�?P���#s7�3i<�D�FZ��~o?1V�?�;	?���=��6�����y@?��?�@�?B(?"���mi=Ѫн�����">Y�>���<�e}>��>�s<��?�k
?�?����o�X��M	��s>�w:?=�?j4��igſ�q�?5l�<���-v<uޑ��Rc��Ҋ���\���=iG�����Ĩ���X�vG���ړ��j���w��� {����>�Յ=���=�b�=�J�<�ɼ@E�<yV=Һ�<HY=�y���@<�;��v���腽b%[��\<�yH=	���k˾�j}?�-I?�s+?L�C?�Iz>��>76�؅�>�V��G?�V>�R�i���|;�|䨾~���Dؾ[P׾�c�9���w>�4I���>r:3>	��=�:�<���=M�t=l�=��\��l=��=�=O�=?}�=��>>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�??ti��d�>M���㎽�q�=L����=2>p��=w�2�T��>��J>���K��D����4�?��@��??�ዿТϿ6a/>�8>�>��R��0��Z��g��	Z��&"?�;�7 ;iQ�>�=?)޾�`ľ��8=�4>��R=}��a�[���=3�z�C;3=An=�?�>	B>�= ���] �=�I=N�=�DP>�K��_;�W 4���@=��=_Nb>�&>Q��>re?\�$?m?���>�蛾��վ�ժ�(�>��k=K�>O��=�3>���>��8?��:?�9?_ʮ>#<�=�ͽ>�<�>u�)�O]l��[�����x��}?�x�?=/�>?��<uA�����8>�܂��e?h4?iG	?;׫>�J����R�L�	�b�������I>�Zw>�&��vꞽ�����<�R�[���gc\>�?�8(?��>!(�>#�m>i>�>M+
>�<=��T�9C	=Bݵ=˻����=��C})��a�=�@����=>��q&���}�ZԼ��=�6���!�=���>W>p�>���=:c����/>�����L���=�����A���c�U.~��/��6���B>�`X>�������?��Y>�?>j�?2u?�f >po��3־Y���Hd�`GR�ƹ=L8	>@=���;��I`���M�nҾ���>�}�>��>p��>@i9��@��@�=X~����8�=��>�t��{RF������o�N2��7����>f���p���*?S��<��=�J~?n�F?{I�?@o�>�C��n5ھ��C>��k���<s@�,�a�Y^Ƽ�?��#?��>�wо:$:��C̾����߷>�)I�D	P�QÕ�|�0����۷����>[�����о73�0h�������B��[r��ں>D�O?��?B=b��^��,XO������h?:�g?�"�>7J?m.?�<��x�W�� Z�=�n?���?�5�?>��=��;���>˽�>A��?Ś�?�{?w�z��>s�K�c��>��=����qŶ�2P뽒쒽@�+?2�;?�2?
�ƽ.�۾0M����ھֆ[���=dT>���>$5b>��&>⎀<N�k��m�j=�>z�>��=�u>�(�>�0d�/}��L?��>�(C>8?m��>B��=�o��<�>��r>pӉ��|F;nٽT�(=��!��ٯ<�G��b��>j&��/s�?!\�=ز\��?{����`>`��=���>��>�*?���>�e�>��>i> m�>J��>IK�>�CӾYx>���GE!��FC��R��Ѿb�z>�͜�_�%�����Z���H�����k�6j�I*���C=�X�<O�?,�����k�i�)�T_��Ap?���>�#6?�����)>M��>���>��������ō��c����?���?�;c>��>A�W?�?��1�3��uZ��u�H(A�e�I�`��፿�����
�_��&�_?�x?1yA?�T�<:z>C��?��%�hӏ��)�>�/�'';��?<=b+�>3*��6�`�h�Ӿ��þ�7��HF>��o?#%�?ZY?TV�w��B�=�H?�i+?ذl?;K0?l(6?S�м	Q
?̸�>���>��?��0?� 1?���>j��=��=�3l�ݥ7=EL�C��n��q�� ���[={=y;���=w�9=C�+��*Z�~�̽!�%�f�=��<� �:�+�=ow=\^�="��>:�M?���>N�>�V:?aHý4���&6��O<?d�=n9�P(G���ʾsľZ�
>8�O?5��?ޓi?��>NhA�di��dj>o�>��X>��>A��>��w�C������=F�=�W^>(Ԟ>?*�9I;�"���.)�hL*�e)#>���>�+|>����K�'>�v��\#z��d>��Q�Gĺ���S��G�A�1���v��T�>5�K?��?}��=[龠��=Df�H*)?�Y<?�JM?%�?�=�۾e�9���J�#O���>��<���f����"��1�:�Rt�:��s>u+��h�n>H�$�,��e7��6@����Yq�=�"���Q>�C����2]��h�>Gs}=m�,�Aw��5��SFH?��O<4���t��v�����=5��>��>��8�����O>�	M��I_$<��>� =�/�=)��|�?��1�y�m>{�7?�P?���?�������,G�Pm����ݾ�_ �.�,?��x>DP�>8�7>�P�=�婾���v�c���*���>��>���bC�Sg���۾~�����=�V?�%�>��>�.9?v!?@N1?��?$�?p[>a9 ���@�OB7?Q��?�b��m���~�m5��>���?�5?!�����>��;?�?17�>1�?��??�C�>���ڞ(�?�>��>0�E� 2��2E
>���?cI�>��7?�?�BK="�k��j�\6ݼ��=%�A��M?��"?&�l>��	>9��>�%��5s|����<�	G?�ww?Ye?H,-�.53?\��=���>{�y>Ok =���>�?��?IPE?=�W?�*?8�q�u^ּio�T�y��Zy=�ż\7�<Tn��D�=���=�߾<�Y�<ކ���>J�<>�>�;����<�0��*�>+t>ᤕ��2>Vľ������@>�z�����������8�'O�=��>��?J��>$����=v�>���>w��A�'?\�?��?�M�:�b��Aھ�J��d�>�A?���=8m�p��F�u���e=L�m?�!^?�X�/A����b?�^?s�=���þm�b�g�龆�O?b�
?}H�Iڳ>��~?k�q?_��>�If�xn�O���KHb�Q�j��=rz�>5S��e��5�>�7?K�>F�b> L�=�|۾�w��}���?&�?M�?��?�*>+�n��.�L3��R��^?)p�>�����"?$C�76ξM���8<�����᪾&�������Х�3$����>�ӽi,�=�?&�s?�Zq?��_?�7 �
�c��]^�5��t�V�з�k���D��<D��ZC�sdn��=�I��������AG=���U��o�?��4?������>�����G��{+�Id�=��ScS��6�>�X��b4�=-�ڼ�坾6�=����F?Ͷ)?��>Q4?��0���y�<�"���#���0��e3>���>j��>ͪ�>5��>Q^�U����1�Tžl��6�V>��X?��;?��?� �=��R��&m�%/�%�>���瑮>�B>�=> ���@h�4?5� �ȟO�����n������<�##?�>Y�>��?�� ??"��M޾�o�k�]�3�Y�}��>K?W�>��0>�m̼��	����>Ҧl?���>dС>Zҋ�3�!���{���Ƚf�>�ʬ>�3�>�to>�C-��[�`E���y��i�8��B�=YMh?�c���]a��ǅ>�Q?�����4<�̢>f�r�n�!����
'���>,?�/�=Z;>Bž�/���{�㍊�~�9?'+?ZҾ+�V��N�=��?�n�>���>�Ǆ?��1>���4g�p��>��2?VYR?s�]?Q�>�,�`�V��ʽ�H	��EC=�߬>BDb>2O�4d�=�`���A/��:㽒Q>Qs;=�-�3$����=������<���=��G>�xۿ�bK��پ��<��?
�\䈾� ��f���������
4���x��i��B(��V���c��K���Qm�\��?�:�?���找n���:���N���C��>r��{��.�J�������Wr��Y!�G�O��i���e�Q�'?�����ǿ񰡿�:ܾ2! ?�A ?8�y?��-�"���8�� >=C�<H,����뾪����ο>�����^?���>���/��m��>᥂>�X>�Hq>����螾<1�<��?1�-?	��>Ȏr�1�ɿ^����¤<���?-�@!�E?���V���׻���>�j	?�*>�m�ǥ���¾=��>�C�?�&�?��=��]� �j=��f?��?��NF�mK��1�=YT�=^��.n���~>�m�>�����L�{���=��M>`!���>�y�T�7�<��6>.]�#���CՄ?4y\��f�ߤ/��T��mT>�T?<,�>?@�=��,?�7H��|ϿW�\�*a?�0�?ڦ�?�(?iۿ�iؚ>��ܾ�M?�C6? ��>d&�O�t��=!Ἴ;����㾯%V���=}��>A�>}},������O�/�����=����ܿ���L���O=g2>�E���,ֽ�d=AS��}6Ǿ�Y��Ğ;&�/4 >��>�|�>�T>@R?\�\?�?!G�>p���?�������k>�Ǿ#��Ғ��'X�w�ƻ�Vྴ���ʗ�7*�AGþ�����<�}��=tHR�^���p� ��mb��kF���.?'&%>˾��M���:<��ɾ�������&����˾e�1��n�褟?�A?\腿�8W�s��(*�����xhW?f�4������ ��=�ݵ��f=8Ԝ>)d�=��⾯,3�bS�~2?6>%?u4Ҿ+����>ֵ��-�=Kd0?�:?R`�*�>�?7�J��*�On�>j�H>���>ߏ�>((>W+��v� �@?��`?�T�;Ń�y��>��ɾ�v��<F�>�xT�Ϸ�*v5>M�{�ؾ��u<4Ƽ< e={�V?��>�)�`C�i��n���:C=�3x?$�?�ϝ>l�j?�"C?H�<K����wS�A�	��=�tW?!lh?�B>�����Ͼ�ͧ�2�5?H/e?K�L>	%i�I��,�.�%����?�xm?Δ?e���k}��\��P#�n6?�eu?,]�ğ�1�v�P�p��>��>�i�>��7��>�=?��
��DX����2�ퟞ?մ@�q�?`�Y<J-�4�=1?^��>�CG�$Ǿ�Zý90����}=V\�>�!����u��� ���0�&7?=��?(�>���r��x�=+���ߣ?F��?i�q�[�u�G93�����U�f��:�K>� �=+k�<������)���X�MT���1.�3;:>#@[��8%�>�	�MCɿ�п�u��!۾�髾x ?�>54�<%��4}�[/Q���8��N��+�p�> ��<��n�h�w�[����H�0:0=6��>�nq��! ?-�f�XN����Ս>&e�>b¶=���b۽ty�F׫?���Б�����*U�fp\?���?���?�7?�6�>����I��ob��!?[B?��T?yfN���*����=$�j?�_��vU`��4�rHE��U>�"3?�B�>P�-�A�|=�>���>g>�#/�x�Ŀ�ٶ�5���Y��?��?�o���>r��?us+?�i�8���[����*��+��<A?�2>���J�!�@0=�[Ғ���
?W~0?{�c.�j�_?��a�f�p���-���ƽ�ۡ>��0��d\��H��c���Xe�����@y����?1^�?h�?2��� #�>6%?��>0����8Ǿ��<���>)(�>�)N>nE_��u>\���:��h	>���?|~�?�j?���������V>��}?��>c�?���=\��>��=����B/�:�#>U~�=�i@���?חM?O2�>�m�=%�8�n/�0NF�s<R�h!��C���>_�a?ioL?��a>������1��� �t�ͽ�Y1�C��0�@�H�,���߽�5>��=>8�> E�%Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��a~����I 7����=�7?�/���z>o��>&�=�nv������s�˹�>�B�?�{�?5��>Ӯl?��o�3�B�&�1=M�>��k?�s?�Jo���ٲB>̶?��������K��f?�
@ru@X�^?(׿���U@����¾D��="��=;�E>X�׽��=Uԥ<���<���w̌=SFv>x�g>���>ޓL>�Zq>3�Z>���Ɏ)�Gs��������?����;4��!T����5�=j���ž�tȾ҉�rL�caܽ��~��l������=rU?��Q?3p?e ?Ƀ�9�>g���a�<k�#�^�=�h�>z2?�L?��*?�Α=~z��g�d��C��X���u����>;#H>�e�>�(�>J˭>��;��I>{]?>̀>%P >��(=�lo��6=IO>�l�>&��>볺>cI`>N3>�B��R ���\j���V�����;�?�h����E�㳕����Bѳ���=�0"?�j0>�*��z�̿�M��_QA?���x	���<�T3�=��)?�S?�x>_������q�>�r5��q�1u�=�ͽ�	g��,���c>r ?P��>��:>s�e�n�K��q�&��DK�>��4?Y�����a�\Ё�'>i�O�8�>�M>�Ӫ=�I.����(脿T�q���=x�,?CK?�	��8����u�Up�����>ɯ>����� �=}�>��&��6��:e��ͺ��#��a�>�?�$>�m�=J��>h���Q�E��Y�>�]M>H[+>�<??j"?J��'��������"���n>��>��>nV>w�M�Ҍ�=D�>L�a>�ۼ4l��oO��<��*X>ʓ��V���y���S=�s��A��=��=��&j9�U�A=�~?���)䈿��=e���lD?T+?n �=^�F<��"�E ���H��E�?r�@m�?��	��V�?�?�@�?	��;��=}�>׫>�ξ�L��?��Ž7Ǣ�ɔ	�0)#�gS�?��?��/�[ʋ�7l��6>�^%?�ӾOh�>�x�}Z�������u�۶#=Y��>�8H?�V����O��>��v
?�?�^�ө����ȿ:|v����>;�?���?d�m��A���@����>9��?�gY?�oi>�g۾`Z����>��@?�R?�>�9�܎'���?�޶?���?��3>ۍ?S�n?�/�>�(�<'m#���� ���~t�<�y =O5�>zI>
-���/�\���r�q��\e�BJ$��j^>���<��>���ڳؾ�˽=u)!�HF���a���s�>?Ճ>}:>볗>?��>�E>M��=�3ż%���&y����N?��?̺��s���;�=6V�]B	?*�6?]�ܼ!�Ծ:��>{W?7$y?��^?�ǡ>�c��ɘ�Iܺ�($��.�<��M>%H?���>f����P>�˾v<�eT�>�[�>]P����־TA���c;,�>�� ?$��>l��=h#!?Y%?�yH>�=�>]V>�����כ>����>ɞ�>y?W��?�C?ݢ��Y6�=ዿ����I N�r�[>��u?:�"?��>����e������~=9n�4�y?�}?��c��>�?�AB?�4?3�>���l���������q>L4?�aN<j`�ҺZ��ԇ��B?q��>'c�>��_�e����3�yW����C
�>�s,? �B?C0���`��{Ծ�ے;�H޼uz�G����JU�;�d=��'>����-�=��&>�C=i ��&�I��^��J>�I>�`�7��~=T��'?��N�\ℾ�t=�1g�&K9�HҌ>`F>�U����P?�8�)�n�����ћ�U�D��?���?�!�?�S����f�W�3?���?�?�\�>�ܲ���뾚9��^�
���$�-��=���>_��������M֭�U=��VP�������&�>�3�>�]'?���>=�N>U��>d�G��ܡ�� &�ظR���*�ێ�|a4�� =��qr�6	�|!=_ξ��¾➻>���X��>TV:?.�>-6�>���>�r�go[>�
J><>���>�nj>y>^�>aZ>l�$�|KR?D�����'��辇����2B?Tqd?F1�>�i�����{���?4��?s�?�<v>8~h�c,+�vn?|=�>
��q
?�P:=�@�O=�<,V��C��r3�����>�?׽  :�_M��mf��i
?B/?@����̾�;׽�梾fq]=BŅ?N�)?
�)�9>S�Un�%�V�1iU� 
���a��ՠ���!�_l��H��/���K����'��<;�,?p2�?���Q���(����j���<�߅h>���>���>ǁ�>kZC>	���/�V�[�$6'�Mp��8�>T�x?��>�oI?��;?#�P?��L?���>P �>�m�����>�;�$�>kM�>�8?��-?`0?�?�*?w�a>���τ��|)پQ?�?�??
"?��?z���GUͽ�ȼ0���~�9���sq|=Ś�<��ݽ�kt�)�k=�oV>5�?[���*��x��F]�>�d9?��>Ŋ�>�8���o��C�:qo�>��>4rx>q۾s�f�P����>��?��E2h=��->��=���3p���7�=�Q�̕`=���<��_�],���=B��=$�P9C��>�3�m�s<" |��;�>a�?�W�>��>�ǅ��l ��m���=g�Y>�Q>�>��ؾ慊�]"���g�U
y>M��?�}�?,�f=��=�:�=nk�������� �����<�r?lU#?�T?]p�??r=?�#?�>���Q������Ee����?aE%?&��=��6������¿E�;�օ?���>� Z�1|=.;m��� �|1�u�*=�Ni�U�u��u����j�}7�(� ��������?T��?�p�=@���!�^;���ľ�? 7�>�A
?���>�F��\H�H�<�)��=�E>qbn?��>��o?�sn?l@.?�h�>�Y(��~ʿE���m �X+�>�??o·?�V�?s��?���>P,z> �(;|�A��� ���7�����&��<R>	�B> by����>���>�"=��S�uai�p���
���G�=
$?>]y=c�>$�~>6�ü��@?�^�>pA�����5��_���8S�=�5v?�Q�??�6�<�"���8����D�>��?��?B>-?���\S=�-��k���ǯ���O�>50�>_�>�l�B�ý�/>.��>��>�{�a������<?$�D?`k�=��˿�z�Ery��֞��ps<#����Y��B���*T����=��� x��?��ܝ��k����w��(�������-�^��U�>�~=��=vv�=�q<���{r<�:�=�T�<��D=6�(���>�2��jGb�3P��J��<%:=�l1=ni��5}ʾ�L|?d�H?�P+?�iD?5�x>V�>CC���>�����?�8W>�&U���eO<�虪�$e��v�վ�MӾ��a������	>Z�Q��7>��1>W�=�|�<�~�=v�=�e�=
��$=2g�=Q�=y��=���=a><�>�6w?P�������4Q��Z罥�:?�8�>�{�=~�ƾd@?^�>>�2������xb��-?���?�T�?2�?Cti��d�>L���㎽�q�=c����=2>���=p�2�J��>��J>���K��_����4�?��@��??�ዿȢϿAa/>�C>.>��S�>v5�iQb�N�Y���W�'�!?�^7�%�Ͼ�O}>�ȷ=y*ݾ;ž�]=��H>D4g=Ď%�^[�q�=c*���� =E�J=z4�>��?>F�=:���)\�=�X=���=;y>>L4��=��:���=A6�=�f>��*>��>�?>�?��g?���>�'Ⱦ������Z/K>�l=���>EM}=d�">I"�>Z�7?�i3?��6?��>���=���>��>i�2�;�k�$T���m��5�&�y?���?Ii�>�MH���s�s��z�F��9�$,?�??Cb?O�>�p�&���S&�n�.�N:��":��+=�\s�M�T����A����ġ�=Ϩ>Ʒ�>�<�>؍y>�:>ԲO>!�>�]>h��<QЅ=К��<�,���l�=`ᑼU��<�0���4#�EX��v-�n����;K�;��Z<�<�;���=�f�>`�>�>P��=Mү�n5>����E�I��7�=綦���A���e���|�$.�+*=��FK>��^>j�t����W�>��_>��D>N��?��u?>u!>QN�8,оP�����k�k�V�{}�=�%>&DC��5<�5�^���K���ξvڴ>HT>T�>�>��9�IP�v�p<<a���E�4b?:��>���Ө���b�P���t���d|��l-�KY4?�Ӏ��F=(�y?�8?/!�?4��>�	��b���>fA�ο=#s���O���=��!?tr?D��>�Δ�[
(���˾�
��p��>�8G���O��Ε��s0��t�(A���Ա>&���о��2�Z4��Tя���B��0s�YR�>��O?���?��a�\>��7PO��}��I���z?�vg?�Р>H<?�)?���Z�쾦��DU�=]�n?���?�>�?ـ
>�Í=Њӽ�E�>Z�>̓�?R��?�pp?��c��_+?@��d@�= N�<d����=�\�e?��'?�R?=��U��⚾���
���T_=�4/=c�s>gR$>�Z�>�I�=��=¡h>\�=
ً>��>d�=��>�B�>����/�{�%?��M>gn>&-?���>��>�Y.�d,V>��8��s>�7�޽�K�<6Gf��;-,Q�i�(=S���>����?Z�>M�ƾ�F?Д��g{9>.q�>n�#>�3�=,�>��>��B>���>�`�>.Y>��>rR�=�%Ӿ��>*���5!��C�X�R���Ѿ$�z>ɜ�X&�t�_����TI�q[���;���i�|)���:=�<��<gA�?FM����k�m�)�7a����?�M�>��5?O����퇽ԋ>��>Iύ>����'���C���">ᾤ�?*��?�;c>��>0�W?,�?��1��3��uZ��u�W(A�'e�,�`�z፿	����
�>�� �_?�x?yA?�S�< :z>?��?��%�tӏ��)�>�/�';��@<=�+�>�)����`�+�ӾF�þ28��HF>��o?7%�?vY?TV��I5�t^=�'3?�1?�j?@
2?�2?:�@�}�?]�I>�h�>��?"d!?�5?B�>Y!�=���=���=�|>Кk��~k��j�^��%K����<B��O%Һ������=��=C.���}켉`�<ؠ<���j?.=c��=�k>�C�>�]O?���>�O>��6?n��������� ;1?��LQk��`<���� �"v>��l?4��?�	g?��u>�a_���i�Wn�=b��>��h>�)>�d�>0o.�i�.�b�;���=S�>��<�_�|)������ž��7S�>u ?�;�>�l�PZ>F.���)f���w>�q��Qą��Qx�N�0�>�-�]F����>�~D?�x?�Q>Sݻ�F:��zg����>�C?��k?�'�?3�I>ړ���uD��i?���8�&��>{G���-�.g���Ȫ�\[Z���>��>T�@�c4��$�h>����n־#j�+E��E�7=�Z�:Y}=�C�q��!?B�l��=�>|����#��0������:Q?m �=�$����\�CӾ��=:G�>k��>2�R��(���=�4B���9�<?��>
i
>��g��R�PI��
�lr�>��??�N*?��?yM��̂��+1�ʦ�6�|���-?ӗ�>Xs�>*~>�Y+��^���RѾPA�L�4�'�>�s�>c�
�>�I�����q�ԯ8���>��<?�Kq>n��>Ng�?�z@?�;?�A?�x(?��>��F2���y6?�m�?�l������`����J��cD�7L�>�{6?�GA�,��>u�6?&�5?��?�?958?#�j>�b���+�g�>iٴ>�MA�E�ÿL�y=Tky?��>��8?�{?<�=s�B�i|��zeѽ�;=T�>�+,?X�>�M�>�C�>�z~>����Ƈ�=��=X`?W��?��j?�v��'?���=b�> �D>.<����>J?�K7?'s�?`)`?QL(?p�������⽊d?����:7i���+h�M+���`8������%�cp���y	5�m1��U�7�G�TJҽH�x��>X{u>�$��1�5>�D¾)���A>�����.�������R4�P�=.,y>wa?a��>�d)��S�=܉�>�f�>����&?��?z�?W��;#b��&־	H�'ˬ>z(B?���=q�n�4�����t���R=��k?�^?�aQ������b?�^?l{��8=���þ�Nb����b}O?��
?M7H�O³>r�~?�q?''�>sgf��m����s;b�Yj�J�=���>�H���d��<�>[�7?��>X�b>�Y�=4�ھ��w������?�?x�?���?�+)>�n�<࿮���ɔ�=�c?�&�>�ט���%?E������f뒾��1���Ͼ���Qq�����H����O��&n�{�d��=OE'?���?z��?��c?t_����b��T]�<�|��g�~��O
��08�U�6���9��S��6	����\�����=H4Ⱦ_�O���?1?�X����>7���z=�{���?�I���sn��,�>�_���.�>�D�rB��.O��U��#�;?��?/+z>�?�8��?�SN!����z�0�?�'�<g�>DWd>��>t����a8����m�d����6���[h>2b?�f*?q�h?�x��q�H���z��,��}5���	��f�>��b>Xt>w7��?�����(����Pf�<��%}��������"�@?���>�c>��?��'?p�D��款��ƽ�N���߬��R>C.6?{&�=�>ޕn>1������>��l?��>��>����N!�s�{�E�ʽ��>Y̭>��>��o>2�,��\��f������9�p^�=ǡh?ᆄ���`��х>�R?_��:��I<�>�lv��!���(�'��>	j?�_�=#�;>ӌž1)�Ϛ{��=��ٯ'?��?H����)-����>��!?\��>���>�'�?S�>Tr��l�ͺ�]?`j\?�G?�9@?���>�)=&��� ҽ�+�2~==և>!a>�Af=v�=��$lX���#�y�,=$k�=�vԼ
�˽ �<|���~�;���<��0>��ۿj�L��4��~m���g��g��T����$��Vj��񃨾�0����A�"#?���0���c��d�70����{�]��?)�?[�y���x��Ǜ���_���Jֹ>�|���.������RJ
��嘾=�׾$���*��L�#�k��G`�Z�'?^����ǿ�����:ܾ<! ?�A ?%�y?��=�"���8�� >@�<�1��c�뾦�����οD�����^?��>���/�����>ӥ�>��X>�Hq>����螾�0�<��?5�-?��>юr��ɿV���/ä<���?"�@��A?��&����RiG=M]�>�4?��;>��3�ܭ�����*z�>�?�ъ?:�I=�X�J�ݼ^e?dd�;IF���һd�=���= !�<���tT>B"�>� �@�#�ܽ�1/>��>q�2�Y�!�Y��R�<�T>�@ٽ^���4Մ?{\��f���/��T���T>��T?a+�>1:�=��,?~7H�e}Ͽ�\��*a?�0�?���?��(?tۿ��ؚ>��ܾr�M?KD6?���>�d&��t���=::����D���&V�i��=;��>�>�,�����O�?I�����=z�	���ֿ�)��>�%`�=9�>X�1���x�<��3>x�[������=�H�����<A�>1�g>�ݶ>F�#>�)l?x?��$?xy>���R��^�__�=�����鼈4{�/�h�|�k���qd��[o�.������̾1�:���=�|P�U����� �G`�~�F��+?��>oWȾ��J�T�&;-3Ǿ�H���������#�ξ[�1�U m�Ѕ�?&�@?�Y���0W�c	� ��Y��Q�W?[#����A^�����=^��q�=��>� �=�v辺62��&S�?$1?��?�ɾRs����(>���Ze�<��(?�[�>�{^�6��>�]!?�X4��f���r>��">L��>w��>���=�w��q����?�oZ?��\������>:o���u�;�U=I�>��/�S�ʼ��b>�E�;-���B�A_����<�b_?(��>U�2��{A��$��%<�<b���B?v?���>�a?�7?�=Ճ� �L�;��� =��2?R�W?�c�=|C�;0�̾���12,?�?�Z8>\��P�j�!��`�4ю>�(?�  ?��t=��~�s:��͞�D$?��v?�r^�ks�������V��=�>\�>���>��9��k�>�>?�#��G������nY4�Þ?��@|��?��;<o �휎=�;?Q\�>�O��>ƾ�z��������q=�"�>%���tev�����Q,�B�8?Š�?���>���Ʃ��/�=؏�����?��?#p��@̼���%�_%�@������
3>�v�=�=������;�Sl�?5!��<B����=">D�@X2�����>�� >�UؿVdп]垿/�����+�?e��>ش�j��き�t���tE�O�R���;E��>@R!>�Zd�(�g�𖐿��H���<��?�/��·>�:N�@���&������7�=���>���;2��rU�8�?�gɾ��ֿMk���\��L?�ʸ?[
�?	�.?�C{������q����n?h�N?�;l?��ھ���&��$�j?�_��xU`��4�tHE��U>�"3?�B�>T�-�Z�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ss+?�i�8���[����*���+��<A?�2>���H�!�B0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?ֵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>bH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�A�>��?�+�=�b�>���=K|��R�4��[">�
�=0�?�pB?m`M?ԧ�> A�=�8��0/��nF�"?R�b2��C�r��>^b?rL?v�b>%1����1��+!��̽=1�/P伩M@�7.�$ݽ��3>�J=>��>�CD���Ҿ��?Mp�6�ؿ�i��p'��54?7��>�?����t�]���;_?Fz�>�6��+���%���B�a��?�G�?=�?��׾�R̼�>4�>�I�>>�Խ����X�����7>1�B?S��D��q�o���>���?�@�ծ?li��	?���P��Ta~����7�{��=��7?�0��z>���>��=�nv�ܻ��R�s����>�B�?�{�? ��> �l?��o�M�B�|�1=5M�>ʜk?�s?�So���p�B>��?������L��f?�
@~u@Z�^?,Bhֿ|����M��������=���=l�2>��ٽ7`�=O�7= �8��:��U��=��>��d>�q>1(O>Ab;>��)>���#�!��q��"�����C�������Z�
��rXv�z��3��r���A��S5ý�y��|	Q��2&�=`��~�=�U?|gQ?1�n?X��>��[�>�N��7�=N�xD�=<��>��2?*L?ˋ*?)��=q�����d���j��������>�tI>A��>��>��>���_K>(D>h��>Q�>�8=�s�;��=;yO>�>E7�>��>$<�>0]>3_���y��#Ɇ�p�e��.�=�E�?ʔ���Q7�#����{о&���AR>�'?kݠ>~����iпs|����N?3(���� !T���>'-?�O?�!7>���[/U�a�ͼj�K��ey��2D>2]v�+�
�K�oSR>8� ?G�>H9�>�Z��H=���t�����v�>�/?;=��������UIN��@޾�u�� 1�>؀=E�E������ ��Z����Dҽ�g?��??���z[����ة��j�	>���=ƍ�='�>�y>�н�s����r��O��,>]>��?[�4>�5�=lI�>�����L�B�>`4>
�">�;?#�"?^�B�Tࡽ�Ny�F7��h>�N�>�>���=y:Q����=���>�N\>��"�&o����
�~�;�ffc>��ü[S������=�v��� >�w�=�m���:��Rg=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>zx��Z�������u�z�#=R��>�8H?�V����O�e>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?�cX>n�?��N?О�>���<��1�|㾿hł�i�b=E�e�II�>V5�>�h���xf�裿eI9�CKl�Ś.���>�G=?d�C�o���;�S=L����V���z���>�Z�>p�s�Z�>�g#?h��>1��>M>B�8��Z���;�K?��?���1n���<uf�=t�^�X?�B4?^�Z�i�Ͼ|ި>H�\?\��?�[?�h�>(��{9���ܿ�π���ە<D�K>VA�>�3�>����K>��Ծ�#D��~�>�ڗ>�W��ھL���P���,�>�d!?߅�>D��=�G"?��#?��.>��>��7��}���?�+��>��>��
?��?��?H?��l:#�UЛ��ĕ�>P@�oT>�Fc?��%?P�>���������%�)�k��O!�QFq?�%�?����VJ�>��?�V?�I"?�a>[��;<ʾ�y����{>	V4?ޏ�=��^���t�fm.��L(?Z��>7ۮ>�˘�B�K��2��n&�d]�`Ӕ>W�I?�h?�`��?O��0��u��85r��ҽ5��=AO�=���=��2>j�A=(=�=���=� �k�i�;H\��K ��Y>H�=��j=@b����!=,?K�G��ۃ�z�=K�r��wD���>=IL>���g�^?l=���{�����x��	U�� �?���?Sk�?���4�h��$=?
�?=	?;"�>K���}޾1�ྫྷPw�'~x��w�
�>���>Q�l���F������F����Ž�T����?��>��9?�Y�>.���=�>����n�8�%�������.l�]Q�6��
J7�_	^�%���rp�*�p�Q�׾������>���� <}>��
?���>b�=��>'�>P�>��=��>8��>�ش���>���>U�A=)s7��KR?+�����'���辝���16B?�id?	!�>�h����f���z?v��?�n�?(/v>�vh�$,+�Vk?[A�>����n
?�!:=���ջ�<(C������%���2���>�s׽|$:�M��yf�l
?�'? G���̾�^׽e{��λp=��?}�)?J�)��wS�nap��_T���X�j��f�V���������r����G����m2+���<%�2?�"�?M�	�����þ�0k�?�6�^t>a��>7��>���>bRF>���G-�q�a�m!�P!�>X�s?��>S6?g�*?�e??8!7?@�|>i�>�����,?�ے>��>[~�>%p&?&�?�02?qu
?�	f?��>%e��x����{��>3��>�W?�*�>46�>pn2��� =;G�=�J�=,K8��c ���>'6>5���I�=��>L=�>�?K�-���0�����5�>ZgG?���>Ŀ�>qic�s��"=P�>���>\u�>s����:x����nA?��?��{Bc=a.>Cp=�E^�ʶ<~�>�~&;�ӑ=��<-�X�-�˼�K|=+��=�s�<��5=^^_�j��S�=7r�>�?��>]O�>�5��E� ���)]�=��X>�S>�$>�Lپ�~��U ��-�g��9y>pw�?kx�?S�f=�"�=���=�{��UQ��m��A������<s�?�H#?tYT?Г�?f�=?Tl#?O�>\-�VI��\�������?j3?��>R�"�����V���,A��I?��?�xI��E�?�C�������W�<��Yl[�������I�)|"���7�c~�����?>-�?��滏�:�y����ا������?|��>Lv�>")�>�&��LW��=�2>��>|�,?g��>��[?��W?�.?�1]>RP�]�ƿ\ŗ��~�=W�Q>hT3?!�?x��?�z?���>#|�>��,�E��8;���-1ٽ3�2�X>�2�=r�>���>�i>�0�j5]�`/�={�:��@d�e��>��>А5>'`	?���= ���8�G?�>������%���x����>�uju?���?w+?�=:p���E� ?����>�h�?M�?*?.�S��g�=<zռF綾C\r�,.�><!�>�$�>�ѓ=L�E=1>��>>2�>���%a�YI8���N���?tF?@n�=
�ſ��q��ap�������m<`���7�d��{���lZ�Zl�=�x���c�����gA[�B���6E���Ե��W��v|z�{��>/?�=��=b�=.�<��ȼc�<ZjK=�l�<�4=Ao�6]o<��6��Q㻆󈽧�D�maa<�I=���Ⱦs�w?>�E?I%?�D?e^�>a�*>Hv�����>�����?CcS>�?n�׺�fH����n����;�Ծ��k�ܠ��>�XY���>�>���=d0�<��=0��=�u=R.<gSO=��=j-�=�#�=��=">��>�6w?V�������4Q��Z罥�:?�8�>X{�=��ƾp@?��>>�2������xb��-?���?�T�?=�?=ti��d�>K���㎽�q�=A����=2>q��=u�2�Q��>��J>���K��X����4�?��@��??�ዿϢϿ3a/>Y>8(6>�7Y���A��-X�x�'�Y�`��z?�0��+Ծ��f>,1w=���Tھ�΃=�!>]�<�!��oV��y�=͕�M(�<#�=�>I.>1��=�m�y=�=l�=)0�=�M>%Ϳ�����+���<�i�=�Y>ܟ>̉�>%,?�[.?"�d?���>��v�Ͼ�?¾�6�>���=3��>��=��D>���>{:4?l;D?�L?v[�>���=@��>W��>�g,��n����A˦���y<t�?���?��>Zk<��6�	7�M�>����eW?kp0?U�?,ݞ>���P��:K�S�6�*����)=�>ڼar��2=m��[���Ͼ�9�u>��>L�>���>i�>>�{>[� >�F�>s�"=v��=���=-$=��f>6 <=>���<5yt>�U�=����<�u�-3��N=�?=	Y	>n�:A��=d��>P�>���>qގ=���+ '>i꘾sJ�~�=�4����@��@d�gn|��i-���7��T9>c�S>�i��'z���?)X>-@7>��?Bnu?A�">9��|־K����Fl��Ae�?w�=m�>�n=�|<�y�_���I�	�Ҿ�8�>��>r�>�>�-��sB��k=���/��8�>�n��Ш��.?�m����@󞿄�i��1����.?~����O�=��?�~E?g��?�)�>��O��⾕�C>�z�`��<%����~�qY��Y{ ?�s?�� ?��Ǿ�h;�H̾����޷>3/I�h�O����0�;q�uٷ����>&�c�о�!3��f������$�B�WOr��>�O?_�?57b��X��SO����E2���u?2}g?�>�J?=?4���~��l���R�=��n?M��?�:�?��
>�Մ�$�k��#�>l&^>�d�?��?>T?+��C?tl����I>�(>=9��c��=����Σ��E)?�xE?�kK?I������Ou�����=�Y�=]�>5�d>KLB>�HW>�,>��f==�(>�9�> ) >��!>@�>eG�>Qk��}+���U?f�7>���K�?jC�>ߌ>�'�=êV>��sΈ���p��ũ>��软a�=,�����۽U*3��;r>)�ÿK��?G�l>��ǽQ?��پ�=�>�j>ý�>�gN<Q��>	K�> ��>i��>�^>F��>ԓ�>�U�>�DӾs~>��	`!��.C��R���Ѿ�lz>Ȥ����%�5��z����6I�Qo���g��j��.��Q?=�1�<�G�?������k�C�)������?1e�>�6?�ь������>���>O��>p8��
����Í��iᾏ�?���?�;c>��>��W?��?��1��3�euZ���u��(A�/e�1�`�`፿�����
������_?��x?�xA?qN�<�9z>��?��%�ӏ�.)�>/��&;�*;<=9+�>�(����`�ͮӾ �þ(7��FF>a�o?%�?Y?ZTV�ȑ�̓>4g2?�6?9s?�'?8�3?��%�ӈ!?w�>��?m�?��!?,},?�>_�L>�k�=W��<I	>�Ͻ#)��<
Ž�4"�2��<�ĳ<�;;q�:�c
�<rL<�6�<2���5<��~Y�\Yϼ�f=��Y=���=⠥>xs\?��>e�>��7?-���R6�~����/?��E=v2�eڈ�r��Y����>rj?��?�OZ?\i>1|D�-�E�>�}�>r�'>��[>�J�>sy�+E�s�=_�>��>�
�=�gB������'	�2M��.޷<v�">Ө�>E��>�6��4�5>M���݆��-]>ۇJ���z$f���D�|�/�0��E��>�{J?��?�d=��澳ů���h��#?_u@?��O?��~?�ׂ=�yվ�<��BH�]��3��>��<��
��ѝ��ҡ���<�BԔ<Z>�霾J���d�Y>������۾��h��zB���徦��=�<�'Ҝ=��.V׾
2e��=f>����!�%���l˩��J?B*�=�j��xaj�Zy;h��=-��>o]�>
-C���6D��¹�mu�=��>>�@>�9>�[���F�F�� �5�>��@?��_?T%�?s�R�^v�U�M�$H��a����漕?���>7-?o�>���=|����&�>a���;��K�>J�>O����:�m"��a���TY3�F,E>��?,5
>� ?�,O?��?�X?k� ?�:?�>s ������&?���?Q��=3jٽ�GU���8��9F��P�>~+?h�D�\��>��?k}?��%?�]O?��?F�><� �L>����>�ߋ>�W�dװ��+^>�K?U�>DY?�A�?L�;>q5�����|��Rq�=�j>#3?#?V�?��>�r�>;P�����=��>��b?w�?�o?�%�=� ?In6>�:�>kE�=�D�>Ɛ�>2�?��N?"s?"WJ?;�>wԍ<୩��ൽ��s�6�Z��)�;�}W<"��=�f� !}��!��n�<�T�;5\���[�Ei�bE�|r���f�;�$�>��s>ʕ��1>o�ľx爾o"A>����t��A�����:��P�=>��?�~�>=�"�i��=��>���>=���$(?��?�?�S�:ְb���ھ�K���>@�A?~�=Ƴl�C]����u��>i=x�m?^U^?��X�s���T�p?,Ur?��8�s�h���lt��/Z��l�!?�X2?�����>�r?+<? u�>�"�6�U��j�>U[��`�0��=��~>�g�����a�>ߎT?T<�>�x>�!���������Μ����>X��?0f�?i4_?&� >�&9���㿎��]����\?l�>*����,$?�P��Tо����*���RY�h%��V���s��~��q�"�w����(Ž�"�=�?@�s?�ns?8�_?�`��b��h_�".~�V����F��v�D��gB��gB�&k�UC�F���Az��|f4=D�Ѿ�+�;��?L�6?���=��?iТ�����L!���>݉���Z��"�>�����>
OF>Gsy��f�=iľ��	?o�?"��>���>sQ�c F��X<�[⾑ϓ�"�V>���>��>-�q>�� ����9=0��AܾD\����y>��_?��B?xm?C�@�8 ��=}���)���������	Y�>-�.>j7d>��H��ｨ�$�`9�Ĉa�T���k��������m?ZƐ>e��>껟? ��>�T�R�s��#����L�ܶ;�ſ�>��*?��}>��>3|�����>.�l?lB�>x9�>�[��>� ��7{��νu��>�w�>�g�>`o>�.�p$\��>������/�8�NV�=bgh?�T����`�8�>]^Q?/�:?	S<D�>o�y�ח!�,��r(��M>�1?,?�=��8>�Qž�����z�x����9?]�!?�0̾v�b���>�~Q?���>�>ƣ�?�HU>`��m��Y=�>��W?�&?�r?�!�>�|�<�ˇ��Խu� ����=6.�>\�	>%\�=�!>A��k�i�0������D��=]�J=���\%>���<b�=��(����=�cۿ�5K� Rپ���k��9
�N����m�����[��"$��� ��r�w����IU&���U��uc�~����&m����?Z/�?衔�/S�����������o��ƶ�>y�q�R�}����'@����]Kྚ����t!��P�/i�?�e�Q�'?�����ǿ񰡿�:ܾ5! ?�A ?8�y?��:�"���8�� >C�<�-����뾬����ο?�����^?���>��/��y��>ݥ�>��X>�Hq>����螾~1�<��?6�-?
��>��r�/�ɿb���j¤<���?0�@#�B?�
"��j��<s�>q�?c�8>��/�^d�㲾v�>/��?Z��?.k=��X�1�4��?d?d}t;�7F��� �B'�=�җ=9�=='�_DP>�>�����E��oӽҷ>ǧx>4�!�τ���U�=�{<ng^>-j½
��Ԅ?�w\�Nf�U�/�MW��W:>��T?�8�>�F�=�,?�7H��}Ͽ��\��)a?�,�?%��?��(?f忾�Ӛ>3�ܾo�M?WG6?g �>�b&���t��_�=ae�Gk����㾳"V�k	�=��>,�>>p,�̌�:�O�vu�����=�$��Y̿�L���ܾ
=��4>d�a>�{�O�*����l��sC��Rq/������ͽ�ώ>�f�>ē?��>�GH?䲅?��#?{��>ٯ�=C`x����'W��1����������d>/��K�e��b޾[`B�����TӾZ7<����=+PR����� ��a�N�E��.?\�%>Q.ʾ2�M�l�<u%ʾ����G���h̤�� ̾GU1���m���?FA?�߅���V��t�B�����NfW?�C�8���������=�F���M=��>�إ=�`ᾑ�2�
T���8?�v$?�k��`���>lpk���4>] ?~?IՈ��ˑ>w�?��ξ8����ڊ>k4�����>o�>��%>�Ѿ��"�V&?ft?��̽�L��,�>_�ھ��=��k>���>�����mL��#�>�fN�������Ͻ��a=~��>�KY?�J�>v�)�G�������J��;�<��p?|.?�	�>�j?*�H?��C��*��p�V��=�T�=�=O?8$m?�i>qV���Ҿ=��d81?uj?SD>�T��q龅,��m���?�j?ٕ ?1�>�q��Ȏ����ȕ,?��v?s^�ys�����M�V�g=�>�[�>���>��9��k�>�>?�#��G������{Y4�$Þ?��@���?W�;<��_��=�;?j\�>��O��>ƾ�z��������q=�"�>���}ev����
R,�b�8?ݠ�?���>���������=a��G;�?��~?M�e�5]@����)I�F��WO�< }�=�=�4�,=�����z��<�v���H��]>��@s�I����>$����ݿ��ڿ�����Ҭ��+���.?Sz�>����[���j���<�=�I�9�8���b���o>���=<��Qm��噎�%QB���=�
?��&����>Lz�<��]����+=_u�>K@�>G����ܽ��ž��?�fپS�׿����9�9��C?��?Fxv?�U2?��=n��1���ĽK�Q?vs;?��X?��A�����ֵ=#�j?�_��tU`��4�qHE��U>�"3?�B�>P�-�3�|=�>}��>�f>�#/�v�Ŀ�ٶ�7���V��?��?�o���>p��?ts+?�i�8���[����*���+��<A?�2>
���G�!�?0=�TҒ���
?P~0?{�].�0�_?��a��p�/�-���ƽ�ܡ>~�0�yU\�����l��|We�&��Ay����?v^�?�?���� #��4%?5�>Z����9Ǿ+ �<�~�>%�>#N>
V_�бu>��F�:�Rg	>ѭ�?�|�?0j?֓������R>��}?
;�>4�?D��=�p�>��=�Ȱ�G[$�?@#>���=i�B���?�M?F�>+��=��8�~O/�@F��R�7��n�C�-ׇ>~�a?�EL?�yb>���@�3��� �>�̽�>1���=@�;�+�mN�&�4>Y�=>_~>D���Ҿ��?Gu�I�ؿ>h���o'�C44?+��>��?q����t�2��8_?Vt�>5�+���#��J&�
��?�E�?��?�׾"�̼~>��>_M�>#�Խ�t�����7>�B? %��C��L�o���>E��?1�@�ծ?� i��	?�!�=Q��?`~����%�6���=M�7?�-��z>6��>��=�nv����@�s�并>7C�?\{�?���>��l?��o���B��1=HL�>��k?9t?�o��󾝮B>Z�?��s���UL�0f?��
@u@��^?�5�ٿ�"���I׾�z޾Ky/=�.u=T�>gE�,t=^�=�M�<���P�f=��:>'%=>�Ʀ>�>�y>Z�>���7~'�Y������I���~��hD��{�Ӿ��ҽ����䶾����Rx��?���1�[�B�-���7����=8�!?��X?�?���>Vß�)�>�B���N�I=�D��ǟ>��?sY?7�?YQ�:8��x2��Q�_�{��DҾ��>#�)=��*?r��>�K�>�d=U>�O�>	�v>��>C���{�<�$�=���>5��>a�?�;>�A>�>T���Q��s�m�m�m�Ϣ���?���8�B�ez���B��0 ����=��-?t�>0,����̿7���%�G??������7��>�y6?K�T?J�>���z\����>Ɵ轷{v����=8��7=����:�D>�? �>��b>9p(��/���x���I���>��?1�9���� ��l4p��斾f��=ce>�)>�־)C��9�l��wn��M=�{C?[|I?e&'�"c*�6wD�����O,>V�H>��>	�<3>2>���v=��-���<�F��$�>p�?D'>�T�==�>�����=�fZ�>FY>C�>�<?A�"?@%��ѽ!m|����xaO>�&�>��p>��>wK�dz�=��>{r\>x=�^�s��"��3�X7Z>�>��"�\�}�����h=xΥ�HE�=v�=��!�8���=�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿi�>�u�zZ�����B�u�h�#=w��>c8H?U��S�O�>��v
?F?�]�����k�ȿ�{v����>��?[��?�m�sA���@���>��?}gY?�oi>�g۾�^Z����>��@?[R?^�>^9���'�Z�?�޶?��?<^I>^l�?�4s?]��>��p���.�zг�,�����s=\�(;=�>�%>�����F��ԓ�#h��*Bj����Sb>�%=���>���������=�����a���ch���>��q>F�H>�	�>�� ?��>`��>;�=-)��-8��O���~sL?r��?���22p�ȣ�<ѥ�=��\�`�?Zd4?\摼9@Ծ#+�>�Z?��? �Y?���>_��͏��Z߿��泾*�<�N>i��>x��>�؋��GM>�<Ҿk�D��_�>ŕ�>�䫼� ؾآ����w9S��>�i ?�"�>��=��-?ti4?��>�e�>��"�q6��r�(�Z
�=p�?�k�>��|?�G??���lQX�l���ҝ��%���Z>�#�?��-?��><3���U��ie���\=�h��K�?�D�?�8��c�>��?�?|�C?KD3>�p;<V\��ǰ>��v�>=h%?D����F�Y�J�@:���\+?@d?3?&��f�.�-Y����(�]�Ҿ�?#�"?�?�R��A��|��S=龼�j,���{�-R�<Js>��r>� �=r�D<L�<
y��7�̯:�;���2�=��>� ^>�e��*c�=,?p�G�;ۃ�<�=j�r��xD�+�>�NL>�����^?Wn=���{���x��yU�� �?h��?8j�?����h��$=?>�?�	?�!�>`L���~޾a�ྻQw��|x��v�o�>{��>,�l���)���|����F����ŽA�i�p�?�$�>W
?��?��v>�:�>�Ⱦ��$�Ab�[��U�G��@%��O�˲.�j�5�r)����ѽ��;=�����Ê��R@>Q`�����>@C�>���>}�>r��> h�=�f>l�=T�e>��=���=,��=�o2>�*(>�y���R?S ��O(�4K�[���o	C?�jc?���>�'Y�Q?���f�|�?���?�{�?�/q>�h�d�)�b�?��>���ܨ	?M�5=3��8��<�`��q�唀���Ʊ�>�)使�9��TL��Nd���
?�&?�z��m�ʾX������=�<y?�h-?�g���K���Y��.b���_�@�*��I��A��v�$��{��8��Eڄ��=u�� �#�=��+?�?�?�{����ؾ��־�r�9�1��l> (
?s��>-��>*"�>23�|�3��M�DI��}����>�`}?,��>hI?�W;?��P?L�M?�2�>�_�>���JY�>ʽ�S��>vK�>�&6?�+?�0?��?wL&?}�\>F��ʊ��S&׾�k?�3?�W?r ?��?^↾ �������N�� ���\Y[=*K;�����]�5Oc=O�T>�5?5��(/����T5�>� ?�1�>���>1�]�_���LF>s��>8�>8ӆ>b�Ѿy��Ö�89?	،?^N�$�˺��!>�6�=^s�;[�q��t�=�@$���;=�-��zA<r�2=���=�E�=j���B;<��N��k�lT�=
Y�>�?��>�4�>/����� �� �_��=�T>90R>#;>�0پoX��IN���.h��u>� �?&��?+o=5��=Ĝ�=xh��}������S�����<͂?�L$?��S?� �?��>?�P"?�(>,���풿��Tn���
?|�$?m��>����hw��K����E���?k��>S�Z�Z����Y0��}ؾ�.����*>���k�"��>[�(�I�G��ؑ��c�?�?l�<-�v�����cǾ7,4?��>���>ݿ�>���A�T��10���=���>��B?���>%~S?��m?G1?ۗ�>��H��&ο!���RC>h����>E?�:�?zD�?��T?:?s=e?Ʊ���<����.�W�K����]�C�f=�:>9!�>EC�>RD>K�[=9W�����8�S�ټd�����>���=<��>��I>�~o�+�G?���>�˿�$��'S��U˂���:�l�u?��?�D+?�=x����E�'�����>�8�?T��?�)?xwT�+	�=��ڼ�涾A�q��>�<�>�[�>@��=cD=8>�`�>�K�>�u��L��?8�:AI�W�?m�E?�b�=��ſJ4t�zz��̔��׃<�>���4X���i�Y��k�=Kі�_J�F1���X���㐏�tʪ�� ���~q�!�>^��= ��= R�=8�<���U^�<Ç[=�F<�F�<��{���<�9�D�M�裃�.�<�ڎ<C�m=��Y���9|?��E?xv*?�J>?�x>�$>&�"��ě>�����?�gV>ýVľ��2�����\����Ѿ;�¾��j��'��;g>p�^�l>��?>��=7�-<R��=�Vi=��=,ۻS�,=L��=1ç=٨�=���=�* >��>�6w?X�������4Q��Z罤�:?�8�>r{�=��ƾq@?{�>>�2������xb��-?���?�T�?=�?@ti��d�>L���㎽�q�=N����=2>o��=w�2�T��>��J>���K��A����4�?��@��??�ዿТϿ7a/>/KC>N�
>+WS�g�5���e��C�HL�#?A�6���˾�Co>A�=u�ݾ1Jľ��=z�5>nn=��^��=�m���K=�M~=���>��@>+�=�s��诨=�B"=G�=�I>�,��M�z�
�&�Y :=���=�^>��>[^�>��?B*0?
Dd?j�>��m��|ξ�-¾:H�>��=ݙ�>ԅ=@A>�]�>.+7?0�C?�DK?l��>;9�=���>��>!X,�<m�.6�"���6��<,K�?���?�E�>{5O<!�@�;���}>���ǽ&�?q$1?Kw?<�>� �5��O�^��������?O��SW>���n�>�B9>^��`���<=�v�>��=�ui>��?��>��>x��>| =w���vJ>@�:<k��=���=7�A>=]<�a>�����~%��sh)��֣��K�=��'>��>��`�-�=q��>:]>^��>��=T���	/>�얾�L� W�=���nB��d��*~�]�.�"�6��cB>s�W>�r#����?9�Y>�H?>�s�?-u?�^ >I��P־�.��[e���S����=�&>�=�i�;��)`���M�/8Ҿ���>t܎>��>��l>q,��+?��x=3��^5��>�����-�V!��$q�,1����"i�&��܌D?wA���E�=�~?S�I?/�?���>��ӯؾ�0>�B���3=���q�M4��,�?��&?�j�>���ŴD� !̾X����ʷ>�H���O�������0���%���{z�>Y�����о�#3�$o������,�B�T'r��޺>��O?W�?��a��N��=O�D�����$e?�og?Xu�>�D?�/?ɳ��"��l�����=ڹn?��?~5�?�`>@v>�� �7Z�>���>���?���?cX?OkS�Ƃ ?��4�u�V>񌣼߬̽_���kM>0�H�0�>!Z??�8?f��m�JQ���ݾ3�8=�]ƽ1e=�O->�}>>e[R>��g>�->�� >I �>�9�>�;&>�a>�9�>H��>�p������/>?�>�͟>n?��s>W�,=:(>�+�>,nȽ�"ܼI�,����<�G4<^�>=�ѽͺ�< q�;���>[����?�l�=������-?+D�rtE>��=�Ǫ>�<T�>��?>{�l>���>'p>"11>s��>E=">�@Ӿ�>����Y!��"C��~R��Ѿ_z>)����&�������/I��o���b��j��,��J8=�-�<�E�?������k���)�w���ύ?�t�>�6?����}���G�>8��>�>B�������ȍ�_�
�?���?�:c>�>.�W?z�?�1�A3�gtZ�k�u�|)A�we�ǹ`�
፿k�����
�p��|�_?��x?XxA?ic�<�:z>���?�%�ҏ��&�>�/��%;��><=},�>�&���`���Ӿ�þ�=��EF>�o?�$�?9Y?�NV��X(��V�=��I?b'?��q?�/?�1?�R����?��>���>_?�+?�8?�H?��>'B�=G@l��49=�}�|�y�1���*�꽞�����=�=4��=;\�:���<���<��ܽM���f�<��(=C�:R�f=�7=E�=٦>w�]?R��>�}�>�=8?�R���8�.����.?��)=*��k���|���m���B�=ϟi?=P�?i�X?1h`>CSA��D�Ŀ>^�>A,&>Q�Z>8ײ>cW��AH����=�\>��>��=�A`�̀�\	�����^��<�">A�>�'p>||��b_>�@ؾ�.���~y>e3�rr������nJ��:�p�E����>jF?�<?zc=�c�n轃�d��� ?�E?�&P?��z?{
H=��\6`�aS�SC����>�f�=ݩ���%���ǔ�e'O��'����.>#✾B������>�z�n�+pk�y?��⾶o=��֖A=�:��۾�ჾ���=���=��ž�`�KF��>���
AB?�N�<������D�5.�� �>�Ř>�F�>�Qv�aM��)%H�Z,���#K=~`�>��B>ඍ��i߾�:�)X
��;�>?�E?>�_?jۃ?be~�I�s�t}F�$3 �7���ݨ���?>�>c�	?�L>���=Ź���L�I�e��E�h��>���>|���G�?����&��,�>V�?��#>u?j2S?:=?�Y\?� !?�T?K�>LIȽG�E�'?�у?C�Z=��߽H!U���:�qF�c��>�-?@����>�.?b!?��'?^9M?�,?tH>F����Y;����>;�>W��h��XU_>ݰN?�U�>��T?҃?�\D>�!4��n��w���^>��>�3?�!?b�?k��>�ı>t��|���!=�(}?�*x?Ɋ?M�/����>�N=��>��>5�_��(!>!?C{5?'/G?}CZ?(�+?di����>�8=ͽ1����?=Hu�<�JY=(��=�V���������q�Nm�ԅ�=:K=D-=Dc}�u'��г� ��>�t>�l���0>sEžZ눾��@>��������Ǚ���J<�/ƴ=V>�?���>6�%����=`ܼ>���>@��7�'?3�?��?5�k;.Yb���پ�{J�8~�>RcA?���=8�l�#���D�u��Pe=��m?�]?�V������o?ENv?�����f�}~��~#3�����u?d�5?=9�ч*>�?�>?��/?ܸ����c������R��V1���=��>��rډ��Ћ>�~?�>$�=�֖<����^�!� ��)�>e_�?�;�?�?>�F|��d¿�y�����(�S?���>����_?t0 �L�оy}��Í�����A���N�����Iپ��d�j��g�iI�=��?3�?���?=�t?�� �&}P�.�d�}+r��_�z4�s��]N�I�$�PN���b��� ��o���]���]�;��	34��@�?�};?ľK���?�첾�Fl��7�}�
>�$=8��Ӭ>���nzz=��>֟���<�P߾��/?���>z�>�}?
u���8�����Đ��[���4�>�+�>\ >��>��&=8���!m=��L�I�X�<e���x�>!s_?`;9?�y?�`����I��~��Ϟ��S6�C��I��>"��={�q>U����m�����2�Y���i)���o����v��"?�)=_n�>�K�?M7?5�4��o~�H!���NJ��ϖ�UЂ>��5?>p��<�A=^��P��>X�l?��>�y�>ֆ��n!�8�{��`Ƚ5I�>��>�c�>>o>@-��\��V��|���9�oJ�=�=h?�f��r�`�'��>��Q?�` :@�K<��>��u�
�!�����#)�XY>�?�1�=�3;>��ž�+��k{�J���54?��'?Ä��p�W��H>�3?���>(|>>�؇?Hi�>O侍\p<��>�l?��?L�#?��>�dʼ��� �νM*4�xq<�h>��>�d�=��>26��hY^�)m��m};�OS< ��o��U/=V�_��}=�j%=2fo<doۿ�LK�rmپ�����#
��舾� ��䟇�f	�Ev��1��8x�����)��V�o	c��v��?�l��y�?�;�?֓�O���b���?���r������>�r��%��髾Vz��䕾���Dʬ��K!��P���h�p�e���'?ݹ����ǿ9����Hܾ� ?�@ ?3�y?��w�"���8�� >�h�<�ڜ������7�οߡ��e�^?���>��0��
��> ��>��X>�;q>	��c瞾��<��?]�-?��>>�r���ɿ5���پ�<���?|�@�IB?X$���I=�_�>��
?��9>c6�����!��>���?�)�?�Vl=LmV�"[?�h(e?�<�;@�G����t�=7;�=65=a���G>�/�>D����A��gܽk~->�=�>��J{���V��K<	�a>�=ǽ�#���Ą?%U\�O�e��W/�O{��A>M�T?b��>���=�,?H���Ͽw�\�I2a?x�?��?�k(?�s�����>��ܾ�{M?Y6?�>A)&�G�t���=<鼥���l7㾥V��@�=0��>��>Hg*�>���hP��퟼���=�[�l
ѿ��1�bS*��w�=6��=�L�<˓l���� ��5b�B 6�~%��V���fH}=Z�r>�`�>���=��>��K?<�q?+?��> &U�b�������F<����a��m�侇S���z�Dʾ����L���҅Ͼ=����;�i�={�R�����+!�>�`���E�4.?��&>q�Ǿ�O����;� ʾܧ�嘼�T���~˾��0�S�m�� �?�@?(f���dU����G� 0��RKW?���O�������=�q��{=��>�3�=�@E1���T��7?�&?�yݾ�v����=���b=��?XE?���帽=�F?kt��T����o�>���L�>=��>B���o���V��?*t?5�/��P����>�}��S֐�������>a4�OXS����=o:����5�J��<�;=:�F>cFW?8�>�F*��U�0�����(��D4=�"w?v�? ��>&qi?��B?;�<
��ɔS���
��p=%�V?�Oi?'�	>9Lt�$eϾ1֫��45?[Bg?�PJ>G�i��辿�-�7���K?��m?7p?}ǳ��T{��e���Q��5?��v?�r^�s�����3�V�'B�>�_�>��>��9��j�>�>?J#��G�����pX4�VÞ?��@P��?H�<<����=�;?�Z�>��O��<ƾӀ�������q=��>c���Zbv�����V,�Ǉ8?Y��?���>]��������>I�����?`]�?����֋��g+�n���þ��I��=����_&=c]-�#r�k�����'�#���5g��<I>�#@BFs����>��\�/�ٿ2e�}+��
���پ��?\��>�5=�s���d�)wf��nu��=p�𬼾"F>�Ԭ=�6�Ӈ5�>K��bcP����<ܥ?��D��!?h	�ٚ)��)<\%���SA>Z�?�;�=\ō�!����[�?).ľ�l࿌���r"8���
?"��?Ln?�*?��>���GӾ�o�A�d?�,?��D?�X��8�_�ED�>�j?y_��*U`�͎4��GE�U>#3?~B�>�-�߯|=1>Ê�>e>�#/�5�Ŀ8ٶ�����N��?͉�?wo���>J��?Us+?�i��7���[����*��V*��<A?Q2>�����!�}/=�@Ғ��
?D~0?�z�^.�/�_?�a�\�p�c�-���ǽ	��>��0�A�[������S��Pe�a��pGy���?Z�?��?D��v�"��/%?�ӯ>A����Ǿ�O�<L��>��>�N>�T`���u>��e�:�"�	>��?v�?�|?ߓ��@����>O�}?'�>*�?L��=م�>�$�=�����/�6�#>���=��A�]�?J�M?��>��=E9��#/�gNF�OWR��*�ίC���>��a??fL?	�a>^���Q0�Z� �,ν�?1�3��`~@���.�e�߽V�4>��=>�>{�D���Ҿ��?Cp�6�ؿ j��'p'��54?0��>�?��_�t�V���;_?Fz�>�6��+���%���B�\��?�G�?;�?��׾�R̼�>5�>�I�>A�Խt���]�����7>+�B?Y��D��s�o�s�>���?�@�ծ?ei��	?���P��Sa~����7����=��7?�0��z>���>��=�nv�޻��U�s����>�B�?�{�?��> �l?��o�L�B�z�1=2M�>̜k?�s?�Mo���f�B>��?������L��f?
�
@}u@]�^?'˥ۿ2P����Ѿ�*��FR@=5�m�t@�=��M���=R��=@��=W��;�p=���>�Ǖ>*�>���<�<">J�>�r��O�)�>4��'ᑿ\�H�\��D���G���3 ��s4����|������.����>�xq�����WĽ ��=�0?FWa?��?B[�>�)��K> ��D�����=�$ƹy�Y>�<<?�c?h�D?� ������Hb�U�y�e���Z���d?�f�=l�?���>	C�>l8>2� >U>n��>�fT>m�3=.e��1Љ���P>\n�>��>���>	^<>1j>�Ĵ���&�h�+�w�0˽��?1���q
J�H1��] ���Q�����=�.?c�>��(п�­�d:H?����+��+�5W>��0?yW?�?>
�b�V��->o����j�c>Q� �ǂl�Ws)�Y�Q>]??�(�>d�Z>59�E�-���q�խ��pC>{O?�ϒ����Ës���g�ɾb��>2d�>�!��M9�Hsx�eap���I�+�v=]3?,�?-�ֽ%&;B�������6�f>	�->i}1=�b�=��=F�2�0}�=�����:ʼ�=�A>KF?�0>�=�P�>�ڪ�y&@�Vݬ>��v>r�[>x8?.�&?ڽ[6���X����h>��>�b�>>ɹ=�]\��S=-��>ʾX>�`�:�q��t�ѽ��/��\>ы���G�˼=7@�<c	Y���>�%3>O�4� ��>�~?���(䈿��/e���lD?R+?q �=ԝF<��"�E ���H��F�?q�@m�?��	��V�?�?�@�?��C��=}�>׫>�ξ�L��?��Ž7Ǣ�ʔ	�.)#�iS�?��?��/�Yʋ�=l�6>�^%?��Ӿh�>lx�WZ������u�}�#=��>�:H?:V���uO��>�q
?z?�Y�}���i�ȿ�|v�~��>�?J��?F�m�U@���@�Ճ�>��?TdY?�ri>sf۾�fZ�䈌>w�@?`R?��>�:��'�1�?2޶?D��?4�L>���?��t?���>�Ӷ�oW8�cn��j>���W^=�Q5��I�>u$.>�ׄ��|%�������������#�A�M>n�=���>:w˽$�ȾYg�=(�A�iC������>Z�>��*>�V�>"B?;��>�m�=��c=�ߘ<�B���۔�C�W?�%�?1(.�/Ԋ������J>(����ۿ>NkB?���L�5�a&�>�y3?�Pw?�A?�ݼ{Z��B����ǿ&Ξ�[x�C�R>��#?���>�
;>	��KM�l�N>��8>- �S���,��!�=���=t�#?�L?(dʽ�.?�a5?�4�=�M�>�d0��L���*��ڢ>���>	Q�>�&1?޿=?�s��+����?%��<�;�MP>R�g??5?{��>�C���E��:�_�����|A��~#?c�?A�>��?`�?Q�L?�U?�>�ၽM����޵=i��>U�+?���;>dN�SO��Z�F?S=�>% �>��=eI ���(�� �����^?f�'?,�
?:���Q�������<�S���x8���>=�X����=/�>ʾ����=��=�ƺc�y�S9���-�5�8>"��=��>.������=,?]�G�!݃����=��r��wD���>�WL>������^?Jp=���{�$��wv��� U����?1��?�j�?���P�h�#=?��?e?�$�>�K��h{޾ ���Qw��zx��u���>���>[�l�g����)���F����ŽɄ�< o?WU�>�?G(�>B|�>��>��ý���S!�w��j�9N�,�7���C��Z����JE���ug������;��4�>�9m��|�>sV�>�.>�?>c��>���=���>��\>��>r�D>�#">�T�>�t>߿2���=��R?�]��GT(����Ű�~B?��b?�Y�>��O��ф������?���?��?H�p>r8h��/*�p4?.��>�����	?�57=5����<(����}�a������ƍ>#cٽ�W:�Z[L��$g���	?V,?}����˾�p�B_��t��=Q�w?#�,?� ��T�96M�jY.�\�`�;/��o��+J��lK9���y��.�����x���Y�1�ǣ:=UP+?*��?	�
��羜����j��n(���>�a?4س>R��>���>��r�+���C�i�,�rd�x?�z?=�>*B?Ҕ/?��H?��C?1�>ƴ�>�������>��<v�>�]�>��?̏?��,?��?��.?o��>T趽F����׾��?!�?�w&?!T?0?��p�	&�yn�jTۼ�G�[f
�M��;3�=��e�ཇ�=l��>�\?�]�O�+��y��з>@/?���>�{>����M��đ�=7��>c�>>�R��
N��
�`��>�.�?�	4���=�,>b�f=��@"��D��=�iн�6c=��;�4����=v�!>"�<̣Q�SGr���#=�W�=Hο<�u�>N�??h�>L�>ㅾ�s ���H�=�SY>�cR>�!>hGپi{��^��*�g�7[x>�l�?�a�?l�e=�}�= ��=���:�����rS����<_`?gC#?L�T?衒?��=?��#?1�>������CI���Ƣ���?��?�;h>ȩ��|��y���nP�G��>��?IhL���>�$����;7��+�>�����R��u���G%��:�;g�	��:��?��?�tK>c� � �¾?��xL�/�;?�b�>�r?�?+���R<!�z�0�_!1=v�<>A?�7�>��e? l�?~,?:|>
�W�Vkο5�����<R��}j?�E�?��?E+L?֡`�2�q>b�>;�s�+m6��w��%}�$Ni�9#�=<\�=��C>�X�>_��>F�>1�����\�O �?����r��r��>jk>Rx?�!=Nv(���F?%��>�e¾%��#���b��B.��4w?o��?��.?}��<�J�JC�����>-��?��?B�)?�%M���=h"���p���q��¹>��>Z�>��=�==z�>��>���>r��P��8��\�0�?!F?i��=��Ŀ9q��ju��e����\;T���7�a�������\�K�=����� �R����FX�W ��Nj�����KҚ�\w�H�>jW�=D��=n��=�V�<Z���(�<��V=�m�<N�<�sq��;{<�<��v���v��0*����z<��X=+) ���ƾz?��E?T-(?��E?pWr>�">;N��p�>jÝ�N�?+�]>O7~��¾�4��i���	����;&W˾Ib�x@����>�X���>6>�#�=��<��=X7o=��}=��<mF3=	��=�Ұ=�*�=>��=�Y>�g>�6w?W�������4Q��Z罠�:?�8�>�{�=��ƾr@?|�>>�2������tb��-?���?�T�?>�?>ti��d�>H��x㎽�q�=T����=2>f��=w�2�U��>��J>���K��L����4�?��@��??�ዿ΢Ͽ9a/>�FL>���=�tP���&��Զ�$�v��31�s9?��:�bA��>@	��˘�����
sv�x�z>�|B�\ ��~E����=q����y=T��=,Ӏ>��X>��O=VU+����=��<���=˷O>��� v]���r���=���>a6�=��>��?-�4?Qzd?�u�>t*x��dȾ����>mv>e� >�߭>�=�uO>2�>e1;?s�??bD?Z�>�h�=�Ҷ>�i�>0%���o��Ծ:=���p=�?��?K�>~�<�x;��G�A�M�Ƚ�{?��2?�?ᾣ>��!:�==�JK7�0�?��=���=�-̾��^�����U�����V<5`=�7�>#��>mר>��>�D<F�>LP�>��N>
`�=�@�<W��=��=���vv�=|hʽQ����2����<��;��k�8���iͽ�5+>�6=BV���e>t�>A��=A�>Id�=4�����H>�i��uoB��r=l7��x@��$m�ԓx��4*��Dt��,W>�j>�˽�>����>h>�W>f�?3Pr?/>go���F׾������I���w���=�=^d`���2�pZ���G�	1�����>���>�#�>��m>(,�l!?��_x=N��$5�AY�>B����������p���B퟿Y#i���ﺮGD?>7����=�<~?&�I?���?s��>4��.gؾ$D/>ab��m�=Q����p��=���?P�&?��>'�뾉�D���˾?i��RϷ>�5H���O�\����X0��g�N��԰>XO���о\W3��x���ޏ� �B�ɬr��t�>��O?A�??Ra�hX��Y4O�Q��lY��3?�g?��>>t?9.?�X��|�H��[$�=�dn?���?�a�?C�>��>���N>���>�Ü?�/�?�#�?Bj��B<�>�|}�5�>�]>�G������
Pw=sS%>���>8UO?�W<?�.��;W�"�ľ�v��/GV�Y�h@�=V�C>SY�>o��>)��<,[==�8=>���>��t>,�>+"W>Q>�܉>^���[�XSg?I�5>IY>ޱ?�>i/�>p�.�͹M>��<�X9�>��E�P��=��=ώ����=p�� ��>�����t�?r��=ꃎ�I�8?)ؙ�&�>�n?��<=iҼ �y>Y&>�	>@g>M`�>i�b>`��>W!�>f�;B�>= 
��5��A���R�!s˾њ�>sw��+(7���
�� ��Z������Q!j�Ң����?�� �<�	�?+R�"�j�D�(�k ��?5|�>�j2?�d����d�e�>��>�F�>{���n���6��V�޾�"�?|�?;7c>��>R�W?:�?&�1�3�uZ��u��(A��e�d�`�5፿X���t�
������_?��x?AxA?0+�<�:z>���?��%�Dӏ��&�>�/��%;�lQ<=+�>c%����`��Ӿ�þ�8��LF>��o?%�?�Y?�TV��6[���> l<?%V.?ݙp?c�1?�=?!����$?rT=>�,?��? �6?��-?*\?�z<>bZ�=ڜ�;;LR=aM���r���۽Gﵽ����O=|�{=�	�;�<��<M7<W8���J�귯<P5����<U�p=�=&��=z�>�Z]?~*�>6"�>{�7?5��&�7��c��&0/?��3=~^�����.��g�񾃥>d�i?��?��Y?c>IaB��dC�9:>�<�>��'>�	\>�ͱ>���9F�T݃=ņ>l`>���=��R������?	��ɑ�'��<�� >`��>�J�>"�_��r>񽽾�|���_>�Y�k�ʾl
�7J���1��h_���>^�T?l��>�S�ݾw����b���?E�I?��O?n�?�Z�=T����2B���[�n")�PH�>��S=����蘿)(��"W:���d��/> ���肯���x>�ڮ������X��F^z�mu�S{=�5�U�9=�q�8�ӾU88��=�#�=,X���&'����r�?�b?���=6뎾d�+�Оž_x=a��>���>��������r(=�o-����q=�ܼ>�4>�-���o�2�A�f� ��"�>bnE?E_?�[�?��$�r�0�B�yu��� ���̼�?j��>�U?�A>v��=�㱾� �#e��-G����>�i�>����G�W���^����$�t��>�?i�>2�?�R?��
?t�`?e*?Y?�A�>���績�A&?��?��=��Խ~�T�M 9�F����>�)?��B�q��>�?y�?��&?хQ?ϵ?H�>ڭ �lC@����>SY�>c�W�wb����_>$�J?蚳>�=Y?�ԃ?��=>T�5� ꢾTԩ�cV�=B>[�2?�5#? �?���>֩�>O������=Ş�>�
c?�/�?��o?xz�=�?�42>G��>@��=ݙ�>���>�?�WO?��s?:�J?K��>Ʊ�<�+���=��/Is���O��)�;\�H<��y=.���8t� X�F��<���;y���R�����2�D����'�;���>I�d>.���->Y#þ�Ԇ�n�5>f�+�v����X���8A�ꂲ=�р>�L?�Е>���ޓ=�J�>�P�>�-�m+?f?U�?�6�<�]_���۾��G���>�=?���=�l�𖔿��u��W=UJh?�Z?�4V�m����b?�^?�T�k=�Y�þ�Zb�Zu��O?��
?��G���>`�~?��q?���>xLf��Fn����h?b�v�j�0O�=���>�Z���d�|?�>�7?�"�>��b>%�=�۾��w��w��N?��?}��?��?��)>�n�00�^�������g?h��>#(��7	?`�Լ�H̾�ג�؎����f��)0��,��yP���j��ʈ���
�)�=�Q#?��x?��z?"�e?��	�^�r��0W���s�]�S�w;��@���E��A��eA��ie��U�8A��ա���)+<(}��*>�,��?��(?5���>������q̾#�>>S�������:�=�n�t_R=^�i=t�o���8�a����$?�_�>�
�>t�A?��[��A�i0���5�v�����5>0�>���>��>���;� &�E��O�˾���:㽅P>m�t?�`H?�e?����8K+���z
���Ǻ�R��/�M>#d>܈�>��x�WS��*4��HF�a�|�p"$�ܶ���T���=�6?��)>!1K>���?��?ո��f���z<�t;�}2�=߯�>�`?��?��>m�������>W�e?Z�>|��>��X��H���_�qq����>�;�>��>��>iS��XW��y���ܑ��
3�s�>�a_?�ܔ�,�ཾgd>	�6?<o�<c�:=l�>�]ŽQ�����)~���X=��?c+�=��>>c�־�S,�ޟ��Q�y�*)?�?����>(��8�>��?���>l	�>�}�?���>o&ƾ=�H;|�?ۛ_?$/J?��@?�R�>��=�K��"�ý�H.�],M=0�>�![>�Ar=�$�=Tw#��Q�KQ�N:f=���=y
�������G<1��L�+<�i=Nm;>��޿�5:��\]����y~����&��T���װ��gt��ž�xr����i	�ò��ÈC���p������$3�׊�?+�?;��=W�d<�Ϣ�o)����p�>�٣���o����u�*�̹y��Aᾆ���"<���Q�ɛv���r�Q�'?�����ǿ�����:ܾ-! ?�A ?)�y?��4�"�Ò8�� >�E�<�*��v�뾤�����οJ�����^?���>���.��w��>⥂>�X>FHq>����螾,3�<��?;�-?���>�r�-�ɿR���Ĥ<���?(�@�aA?��(�V��`Z=�V�>W�	?�N>>;T3����t
��sr�>� �?Ĵ�?��O=3]W����[ie?UJ�;G�F����̱�=!�=��=�����J>q^�>�u�f�A��I߽��4>l�>8�%�6���x^�oƾ<�\>��Խ���Vӄ?�\��~f��/��)���>�T?7��>z�=��,?�UH�c�ϿW�\�~�`? $�?[��?�)?vd���Ϛ>�ܾ1M?��5?��>�/&��~t����=*����=����~�V����=�n�>�>{�(���-NR�?������=T(���ƿ��$�t��+�<07l�:]���ѧ��E������k��.�;�f=��=)iP>p܅>�qV>�U[>�W?W�k?ܿ�>�x>�߽ѧ���Ͼ�s��ꁾ���e�����/��������޾	�ft����o�ɾ��<��K�=*9R��u���� ���b�%oF�x�.?O�#>˾��M�Y�&<ٌʾ���Ag���E����˾��1���m�Ԥ�?�B?6��V����S�	�E����W?@�������T��=�K����=���>]K�=��&3�]�S�AN0?��?t$��h��wf+>���'S=$u*?�� ?@�<+�>C$$?�(��߽� [>�3>_d�>���>��
>���_�޽��?��S?��� ��J_�>;a��]Cv��2_=��>N�0�񙭼f`>\j�<���큄��鍽�3�<AU?�P�>?<�� ܾI�K�5�=}�>�q?>w?Y��>\�r?�]?��'�����
n�2��3/>�Bl?C6P?��==��;����9�RS+?�Y?��>�m��,麾�D�9��'�?HY�?t�)?�$i����Tt���.�NC??ABw?V^��m�������l����>5�?"U?Y�4�Vc�>�E9?��^��M��"ƻ��,�2��?��@���?�*�<�����!=�a�> K�>8�.׼�����6���o=-
�>O㝾'�c����Z�(��>?�y�?Q�>pV���\��V��=#ԕ�uY�?��?d~��u�g<}��sl�j��-��<1ѫ=���YA"���)�7���ƾ{�
�S����ƿ�ϟ�>�Y@9c��"�>�=8�03��RϿe���[о*]q���?f{�>&�ȽL�����j�gOu�ʴG���H�t����Ƿ>���=������_[i�Y���� =�2�>���el�>� ݽ�wپ��о͜D;܈�>�v�>sM�>��E��ɼ����?���T������8�/���&?�)�?�K�?�d?v�f>17���&ھk7j=Sp*?��b?�]?猽���A����=$�j?�_��wU`���4�vHE��U>�"3?�B�>O�-�r�|=�>���>%g>�#/�u�Ŀ�ٶ�<���V��?��?�o�"��>q��?us+?�i�8���[����*�#�+��<A?�2>���J�!�D0=�^Ғ���
?S~0?{�d.�(4b?�o�B:�� H,��yܽw>��-�BY��Y��=}�j�z���Λ�K��s�?V@Å�?���*��+?�>�Ά�#	��-آ���O>?q�>��>e콇�w>�/@�)?e�'��>*��?�@��?䁞�k�����=���?C��>ߓ?_ >��>�]>��56�"�(>r�z>C���μ�>�IR?}�>3�����;e$d��d��~b�����R9�䧾>C8?؉?Fb>�V��49�F���]�̽�&��vR)�����(��ݾP>��0>���=�����	��?�'�e�׿�X���c$���3?2؂>�?���v�>4��h]?���>�	�u3��HD���'�B��?��?�A	?�Eؾf3���O>Ņ�>G��>��нy.��/���?9>�CB?����Z����n��t�>R�?U�@R�?Y�h�1�?=��!܀�����'F�s�:>>?����}��>�Ǩ>c����s�82��Z<i�4v�>8�?T%�?���>!j?M�t��fX�ڶ�ĝ�=�(A?��,?O�>�������>�q	?���ca������?�@�@��>?^����׿)���e��S���w��>���=�!��>���=>">р�=Q�G>�Pk>0�#>�*Z>��v=r�A>�g >�{�e�%�d��$U��(�c��o�k�˾;al�h�񾂏�$C����	�� B�����	�)t}��1۽�K�=e��=L�U?��Q?��o?8^ ?��z��>���#y=x�#�:O�=!ʇ>�c2?KEL?�0*?�ؑ=T�����d��R���.������}�>�J>�(�>�>?	�>\ja8��H>(�?>	��>�� >L-+=H�u�Kj=�~O>n�>|��>Bz�>�C<>��>Eϴ��1��g�h��
w�o̽.�?����S�J��1���9��Ѧ���h�=Fb.?|>���?пc����2H?&���v)���+���>z�0?�cW?�>����T�.:>-����j�@`>�+ �wl���)��%Q>wl?�m>~"u>)34�M�6���K�T��6v>��1?+���q�D�$u�/�G���پl%N>&�>Mv/�;k�>"�� �x�7Bd�D�b=�~9?�;�>n3��������� ��2�V>�.S>m
�<���=9�`>N?�]&��b�@���<D��=v�a>e�?�D->
Wy=��>꾔�C�J����>?8>֙(>\�;?'4 ?>��+��N���=�6���m>p�>%�z>�>1�K�R�=���>��V>.m�R���M���/�/cT>JY��Qj�[ٖ�@�{=���o��=`l=��>�H�pb�<]s?� ��q_����/�������+?{�>?uu>p�
=DA>���ſ�F�����?�e	@���?�7ؾl�P���>��?�␽� >��?}cD>V< ������>}�}�V���Hr��	�=�f�?#��?Ն�������_��>��>�띾T��>�Q��� !��ȹq�@��<�e�>k�C?3���l�R�D�m$?�?4�򾓫��#ɿ�Fw�N�>>8�?U �?�gm�������B����>D|�?�YV?�{X>��۾�Z�"��>�t9?1K?z�>���d�#��?ɒ�?��?�">?��W?uL�>	�%=J��ˬ��>u�Q>��^��o>�k`>Ƙ���6G�����&���]���1�b�=���>��>X}Ҽ�c���ҺQRQ�l|Ҿ#��$`�>�>9�j>]Ԕ>3&�>rJ�>�H�>�֨=_�B��ڇ�X�ľu�K?y��?&���2n�WS�<x��=��^��&?dI4?{x[���Ͼrը>׺\?a?�[?d�>N��8>��迿~����<#�K>:4�>�H�>6$��EK>�Ծ4D�Jp�>�ϗ>	��>ھD,���4��mB�>le!?���>9Ԯ=P� ?�#?�j>>+�>�ZE��5��G�E�E��>u��>�J?��~?g�?JϹ�OZ3�{	���硿ܒ[�>:N>g�x?�O?�֕>w���ǃ����D�_I�A��옂?�ng?�q彼�?�-�?��??5�A?�'f>����ؾK���>7!?;����eC�Y"������>���>'��>s
��R�������e�����?�M?xa ?� �K\�����4��<���<�T��@�8��QY���=��%>n�����=��>q�[=S�}�KN&��,<�$�=�}>
�e=�7� �ս�,?G	����V=:�j��m@���>k�u>���X�[?���n��1������`gl����?��?���?�׽N`���;?��?��?�l�>(砾�[�l��dYX�^�c�5'���=>��>l�<JE �p����=��}���5c��2r�>��>��>?�
�>�@>^�>����n%�Tk������\�pF�N�3��+�''��Т��*�¸�8`���Is����>��$�>�W?&�Z>�>[��>��O��ʄ>(=R>X"�>�>&e>��/>��=[� <�ͽ/?R?כ��q"(�}���I����A?	�d?�b�>;�e��I��gp�[;?H��?>r�?��x>t�g�{�*��?J%�>&1��t
?��G=�ǻ��<�;��0��wS�����We�>\V˽L!9��L���h�6(	?�<?�H���
̾��׽����:p=s�?Y)?A%*�c`R�'�o�}�W�S����H�h��k��_�$���p��؏�@Q��D'����(��)=a�*?b�?�t��^%��� k�z�>�bf>2��>m�>v��>��H>��	�u�1�u�]��^'� ���!�>S2{?��>�_H?�n;?GDP?b�L?崍>�u�>�籾i\�>�7�;�+�>��>Q:? �.?c0?6�?0*?�b>�A�����Bپ�,?k�?�?/�?�c?�x���ﾽ�k�' "��Ix��r�W��=�>�<H�ս�Is���W=đT>"x?j��7}<������W>�E!?���>�>�x��&|���������>�c�>��>#����b��d�>\�>wVx?w���=p.>�S=H��;�4� ��=�|]<���=�Fܼ2Zq�ӟ<�w>�e�=DP=�:���W���:<�@�<��?�?�?v>wQ>�Hh�����yɾ��b>�P{>-_�>�ު>�琾��]�����n�Q��>Y�?5��?��λ'�=�s'>F=�T 8�]�ܾ�߁�'������>��*?�L?~�v?�Y?R�A?�0�>F4�����Q��6�־#m?SO,?[��>��|�;�g��lf2��f?R?y�_�H��z)*�7[��ұý��>�,�w|�5?��Z�C���L;���폽l��?���?��(�-(6�y��P)��]���u�C?���>���>Tl�>��*��0i�H���!?>�7�>Z�P?�t�>#͗>}�??���?��>�!�N����Y�����=#�ļ.��>%�(?���?�Š?�?�[�>sh�j ��o�$>��z��T�St���=�&#>u�O>@��>x�>�!�o:Z=�q>�5���7���q>.#�>�Y>�=�>���=�e�[~E?�Ւ>t{ܾ�>������z�~��>��?t��?�&C?�p\>.:<� '��#�.��j�>�?�а?��j?�z���=��Q=&S���L��=�>��C>�z>һ7>����P*�l�?47?~]��F���^�Qw��d?�9�?E���ǿ=t��w�k뙾DlP��⏾3�]�f���GQ����=���m��E���U[�����?@��Ǹ��u��Ϗo�v��>�
�=�;�=yA�=7�=��Ѽ�Z�<��==l!�<Ԋ(=����g�<?J��û��z�OȻ*l�<�8=恻z!�W�?��F??�?z�$?\=�>f#>��>���� f��D?�?�>9p�=ځﾆ�ľKO⾭6$�1T߾dVA��V��0��d�C=�h��_>�AF>�s>X��#�C=�y=��f=2-��,�<4 �=>��=���=jJ>\X>�O,>�z?�K���1���X�y�֊?�P�>+[>Cl����Y?�a�=�ד�}���,	�bC{?w��?���?A�?? �b�>�+���:P�P!>�O�`��=8}��q���N��>�j�<�f;���@��<���?��@�lM?˪��@ſ�+>�qI>�>�GS�PX,�d�J��{��;Q���?�s6�o�Ӿ�HZ>�^p=��վۢ���s=��.>5˸<��%��%O�g��=�x�����=�w�<�+�>��0>�gR=dF��ד�=�$	=��=R0b>p_=�a;�3�<�J=�k=��`>��1>���>6�>&
?��X?q�?���<ɴ��h ���e���!��a ?E3�<M�!��*�>ըA?�;?(Q?�x�>��H�A��>�/�>ǡ�F�����Ř��O{�>�ȟ?�(�?9X�>z��9!������@�!ƽI�?�4?ɛ?ݐ�>*W����� �d:2�ae���ta=��=����	[=V
�>�z%���=�=���>�%�>u|[>ձ>�+>`2�>ң�>�$>�2�=�Q=��>��<��)��o��Y#�=��9�4t>2������Ћv=��ʻ���=Bw ��0I=I>���>^$>�&�>�+�=�!����5>�5���4:�YG>)���_p-���V���y�9�Q~�L�>׿H>��+��ې�Ӆ?�1'>C9�=���?��p?n3�=c�QӾ�M��򚈾wHz��͌=�M�=��-��y9��zi�Z^��ݾ��>���>>�>om>eD*�i�<�2|=i\ྲ�3����>����b�������p��`���4���_i�m�4�ED?16����=x�{?�CG?ri�?��>v�ԥؾ�v.>7m��q:�<�[�z�q�q>���[?͕%?q��>����D��)����Ͻ���>9���y'�i��4D$�U}Ͻ�Už�;n>�\������1,$���{��Ó�CV�6$��o�>�[?X�?����q����%]��׾��>w��>��C?�s>?> ?u�?>D{����Ϯ<�(P�=�>q?Z�?���?3�>�ý=����2�>,	?���?M��?8zs?��?�~t�>6�;B� >�Ø�!W�=��>���=8�=�m?׍
?�
?�g����	���s��^��Y�<���=ބ�>�i�>�r>���=�zg=2t�=�/\>�۞>��>�d>a��>L�>�{k��a��z�?ay&=��>�?� >�>s�[x�E2��2	#�Ae$�f��
�;������=F�˽��<IGv=��>���Gi�?�I�>�,Ҿ�?�� �z�.����>`xU>�i��g-?6�>��>��>���>��=�>���>ʎ���� >g�5�.rپ~b�K��ꇺ�[�g>v$��m>�����n5��XS���¾0��6q�oU���G�Afk<�~�?l�Hp����N�]^?>��V?;U�>��>?D�Ʋ� _>d��>���=D�2H���Ր�*���+�?`��?�d>+�>�;U?�r?��!�-'&��Z��x�p�E��ye�?�\�~8���S�����*��W�^?�x?��>?��;��v>���?��%������Ɉ>�}-�*c7��T=ߨ�>X����]�P=ξF�ƾ��&��A>�vm?ɐ�?G?�[�Qeb�0!">��9?)�3?Ʊr?߬/?�7?$S��k$?d)>�?4?e26?�p0?z-?�r6>���=�L��%�S=�̑�t���νCGн���Y =z �=r;�mT;�Z=q��<j�m�
�+�,;�P��K��<�1N=�9�=!�=<��>	�\?p��>�Ç>_s8?|���8����r�,?�,=W���i��c���7��H>�j?b٫?��Y?�u_>@A�e[@�s�>h�>�v%>�\>g��>��]E��Q�=�> �>/�=�+]�����Z	�SR�����<{>L�?��ػؼ��T�p>�Y˽o�)�D^���)����̯�d���n���0���?V�C?��?�
T>�޾�<=��2�eO?(�?(F?��?Q"L>b� �y#C�t�]������>C2���Y���舕�Qg�f�=�P>���þ:y�>��t��aݾ-�~�[���F��>C�.��=x=m� ��^� �,��^�=V>&�Ͼ�����u���0h?���<�J���S�Eo���=�i>�w�>���5�=k�5�������=��>
�>&g=���
��#E�Z���=�>7RE?W_?�j�?A!���s���B����Hd��s ȼ�?�y�>Lh?�B>R�=d������d�)G�b�>���>�����G��9���/��p�$���>9?8�>r�?U�R?.�
?��`?�*?iE?�'�>������B&?)��?��=��Խ%�T�� 9�)F����>r�)?�B�͹�>3�?̽?�&?�Q?��?��>� ��C@����>�Y�>��W��b���_>��J?˚�>q=Y?�ԃ?��=>M�5��颾�֩�KU�=�>��2?�5#?C�?鯸>���>񵡾���=T[�>|�b?�ς?��o?���=��?�b3>D��>L�=�ƞ>V��>�4?v�O?��s?�J?-��>捌<����/b����w��!0�W:�;��9<g}|={��}+r��v���<㊝;a�ǼR$��2f�j3C�Q���[��;F�>�z=2�i�
�>�;��k��,�>�L������4��Q��p�D��>wQ%?y�>�3c�Ն>,O�>�~�>�+�� ?k��>.5?�[齫�]��0��E�S�ⳟ>;|!?��n>1J^�������N���={U?4�j?�U�����b?�]?�i�R=��þ[�b����8�O?j�
?|�G���>��~?s�q?���>:�e�f7n�;��jCb�W�j�&ʶ=Vg�>�S��d��>�>;�7?�N�>��b>.*�=&u۾a�w�.p��??F�?���?���?V0*>��n��1�#!��I����^?�w�>�����1!?[�O�Q�; ��6B�����5Ԫ��e��a3��������"��U��j޽���=Ä?�u?�s?$�^?/��q,g��8_���}���X�������\H�<�C��XB���m���1���p��<2=�>]��<�-�? ["?�9�E�>�'¾�<��־�?*>�y���S�Չ�=����Jp�=��=WV��4����u�?�s�>���>�aN?��`�]�=�Z�4�%,(�Ko�L�>e�>R�W>�>�>���=��Խ���ܞ�_�z�����p>�df?��K?��l?x��-@0�Ǡ��Jv ��vY��T����H>�g> K�>�uW��})���(� z@��Nt��,�2͔�����>h=��1?S�>�>��?4P?F��D��A�����.��؟<�U�>[j?���>F6�>�ٽ�#��Z�>\rk?��>w�W>3eJ�(��to_�nڵ����>݌�>�?�>�6�`rZ��������ԕ>�=;�=>me?yO������>~B@?��2���";6�>W�뽊����q�'I>8�?V��=��U>Ԙ�W�.�����S$j�E�*?�L?C��!"���j>@�?�r�>`q�>z��?�e�>cѾ��ټ�?}
]?zkC?o�<?���>�`�<Y�6�)Ž��Y���=sn>b?e>P��=�m(=�]:��`a��J5�j�=h۟=��ܼ�u��ܣ�<�P�;�v=4 #=�7>��ٿ��1��<����^�ML��5ľ���$~�7{M��}��,��D$&�� �!��;��7�A�V�%G���f0��E�?\K�?�E�=�+/����_�#)�L�>ÿ�2�����¾��ξJ�x�'�ƾn^��6��Hj9��(=�yn�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >cC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾t1�<��?7�-?��>Ŏr�1�ɿc���¤<���?0�@�@?Ӥ$�g�i��=��>��?iu.>�QR��F��Lþ���>�z�?9��?\�=��T��7żX�e?�r�<�qK�|{3����=��=c
=$��]#J>p��>hP��9����"�0>�>�OC������`���<�xU>�m��э��ӄ?F�\�]_f��0��`��j#>��T?у�>gW�=~�,?H�H���Ͽ�=\���a?�)�?W��?S�(?�����p�>��ܾ�M?�+6?��>��%��ct��c�=�ܼ����w�V����=՛�>{>�z,��f�IQ��(���'�=o(���ÿN.�65%�de#=
�X==�g�ŌĽ�h�2,��Ꮎu�:�5��H.`=�	>#�O>5v>_)>�Vm>�JX?y#q?��>Do>X��6���\�ξ
`5<�+����9�����g�n�K���P�⾴Jվ����������=��9!=�{�=�5R�O����� �)�b�ϗF���.?at$>L�ʾd�M�0�-<�oʾ+���Gل��᥽�-̾�1�&"n��͟?��A?������V����b�؆��l�W?�R�D��jꬾ΢�=���à=�$�>ˆ�= ��� 3��~S��P3?M?��̾�h�\�>Z����=D�#?Ww?�=>-�?���8��aT>Z*>�!�>���>�1>`W���٧�� ?��O?[� ��$��K��>����KM����=�Q�=��J�p�3=�(a>q
ܻ�T��t���긽��=�cV?��>\�%���0i�yT�;샐=L�w?��?���>_�?�{Q?Jj�*i�j̄�S���xD>ꇂ?ȯX?ٽ =�>�����hþ��K?�^(?d�=�j��]�P���A��D7��B?)aW?�B#?��w�0���`��;^O���?�v?�Y^��s������qV�[�>�*�>l��>�9���>Ί>?A�"�P��7����K4�5��?�@��?:�4<4���I�=�8?�-�>w�O��cƾ�=��O2��2�s=5�>����DQv�����L,�j~8?+��?���>�x��������=�ٕ��Z�?��?}����Dg<R���l��n��`�<�Ϋ=���E"������7���ƾ��
�����࿼̥�>EZ@�U�x*�>�C8�\6�TϿ)���[оSq���?K��>Y�Ƚ����A�j��Pu�a�G�2�H�ť�����>�>�5��̉��t���7������>�3:�z>�oG�,��`����٫�փ�>���>n~�>d�	�g¾ڀ�?���u�ÿ(���g���)F?�Ƣ?���?\+.?+��=z�K�����:=�/=?�m?d�X?ӸͼV�b�&�0;��j?G���P`��4�R;E��U>3?�8�>��-�{�|=X/>��>�U>�$/�ǐĿ�ܶ�l�����?х�?͂�}��>�~�?%p+?j��1��Y��*�*�{l0��5A?��1>�s��Ȱ!��&=�9���,�
?e0?���&�je?2j���%��A~��Pݾ��>9!?=�;��b�^�T$���F��{�����m��ڹ?�E�?���?�K=�"���?�c�>j#�EA��Am*�OO>v�i>(x�>���=�%>��ľy�1����=���?{f�?}Y?I&{�=q��3�����?0��>/5�?�o>�ġ>;��=���/���f;W���TN��Q%?�K�?��>V��B��Ќ���>���Dq������d��a�>��C?�5?�"�=���	���3�$Cܽ�k�\Th��9M�d��=م�<F�>'u>c_�=����\���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��� ?C����\�Wx��b־�ş�X��My5?-�\Dx>���>#hm=0����	����t�L��>��?���?��>�؆?��j��0��h��=|��>9
�?�?��������h=E��>Q�!�����Nþ�A�?�@!�@�\�?N���ݫ޿�r���]���4Ѿ��=�=�6>��N>7�T=���` "���>��>u[>��J>�{*>Z�	>�,>�U��if��(��#�����7�n��i(j�b���sV��������J����ڽ�X����L����������=��U?��Q?��o? ` ?�`z���>�i���=#���=�V�>�j2?�XL?,*?"��=�S���e�Q:���g���D��'(�>�CH>\y�>�;�>��>��8%J>��>>��>�� >_�'=�����=�^O>�n�>y��><�>�C<>��>Fϴ��1��k�h��
w�p̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?~h><�t>��3�b�7���P��l����|>?�5?���K�6�n�u�-�H��cܾ[�M>�}�>��A����AՖ�\~��j��Ix=fC:?�+?�|��駰�P�t��c��3QQ>��\>I�=p}�=�N>}�`�?4ǽv#H��+=y��=�k^>ѡ?>��T��?�>@0����{���>� >��D>x�N?ݳ�>�н�����H�߽Ӑr>�>c>�O^>��m�Y��<�9�>v�>�¢9h����ᢽ �O��^>qɄ��f�����%>vT?�w:�=2�>=����^/�A7=���?���� ���޾6���^VC?U�f?"��=KϽ R�~/��������?k�@r��?L4��7�V��A�>�N�?�Hؽ�~h>D�?֫�>0鋾�����
?;�=�8��P��y�:�8�?�&�?��;��fb�|�K�I{�K�?y&��Qh�>{x��Z�������u�d�#=S��>�8H?�V����O�n>��v
?�?�^�ߩ����ȿ5|v����>W�?���?i�m��A���@����>:��?�gY?moi>�g۾>`Z����>л@?�R?�>�9�y�'���?�޶?կ�?YI>��?��s?Ej�>� x��X/��3��̔���=QHX;jj�>�q>����1dF�	ؓ��i��}�j����i�a>�8$=	�>I佯)��&P�=����'G��O�f�e��>q>�I>TS�>�� ?�a�>���>1�=2N��〾�Ŗ���K?`��?���2n��L�<���=!�^�g&?{I4?Y[���Ͼ ը>��\?]?�[?d�>M��4>���翿
~��h��<\�K>y3�>�H�>�#��0EK>!�Ծ�4D��o�>�ϗ>����~?ھ�,��G��tB�>�e!?���>�Ү=ܙ ?��#?ҕj>5(�>�`E��9���E����>g��>�H? �~?��?�Թ��Z3�����桿��[�,;N>��x?�U?�ʕ>2���у��rE��BI�����(��?<tg?dS��?12�?ډ??C�A?�)f>Ĉ��ؾ������>٨"?�����@�Q� ����b?�}?)�>#�z�5���tpP��'������?X?��"?����j_�+��7��<.���k<	��C���� >NB>�����=�H>h��=S�h��~*�7ٖ<��=~ߕ>H��=i-����e,?��=�0:���7�=�Wr��B��Y�>i�V>=���`?�,�3y��¬�$����M\�
ߍ?P��?��?����e�.>?��?�'?�#�>�\��O.�T��/���o��^��1�>�Ľ>/��f{�&𤿩���s��^���]~�,V�>�D�>�?���>�N>x�>>���zK&�'�����]��#�Q,7�j�-����0
��KU#�	���: ¾>3���>������>��	?�i>�	y>B��>�黟x�>��P>�G�>�8�>�V>У4>t� >�9<~#ν]�V?�=��'����h�޾�;??�o�?Z��>���9�e��N(�}�?L@�?��?/#�>t�C�	4�$��>R�?`�z���?y����)�@���ž�ɛ�Uѽ�`�=w��>��=���s�,���R�>�?�7�=����:2�� �-Eo=���?YQ(?:\*�4tR�>!p���V�]oS����<�h��g��@o$�$�p�؏�%����$��Ȩ(��(=��*?��?n���c�7��D�j�b�>��
g>y�>+��>���>�K>K
��2��r^�-^'�䜂�q�>��{?p��>�nI?��;?7tP?JUL?��>�S�>�I��[`�>��;SΠ>���>�9?��-?d-0?�s?SV+?h�b>h���������ؾ?�?�:?�	?B�?���ý1�����e��y�*��[��=�<t�׽at��T=3T>�?�?�^9�Wm�sY>�H.?��>���>&���@Q����,�>�?%��>.c��� l����M�>,�?j�(�u��a5>�n�=��}����:d��=c�ζ�=�`���������;�R�=�1�=A��Hg�;�Ŷ;�R	<�Z�<٨?��?�>>P�>�/4��,Ҿ�����&=�\\>~�<Q�">�����������^�K��ϔ> �?H|�?h�p�,��=�G�;�O�k ��? )��~���T>�3?��N?�{?hć?�"?�$?Y��=�����}�e�e�{o��*�*?0!,?���>:����ʾN憎��3���?�X?�:a�а��8)�ׇ¾��ԽQ�>�]/�1~����2D��m�����lq�����?�?�1A�k�6�2w�¾��Z����C?��>�Y�>��>�)���g�f$�!;>u��>�
R?�m�>��B?Qjv?j�_?ȽF>_�3�`㭿V����ռR>9?@s?�5�?�|?d�>�_'>k��޾��ھLq=�)��>dm�i��=�7#>-ń>u��>aT�>a؏=��(�F���[�=�{=�2>�-�>[�>���>�u>I���B?�X�>�C����/3������� k>X��?�V�?�B�?cՆ>����hkB�6���>���?���?��`?���q��=�$m<�]�j��Ҟ>��>��>�
>�>�I�>/B?`��>�P���l��i�PΘ��>��@?��>>��ƿ�r�Cuo��ך�X�]<4���f�o��+CR����=�����O��榾�Y�%��X��w⵾U���,�|����>���=�%�=���=��<����%ݼ<?�G=�$�<��=>)f��C^<��8�W	�;���7�FfZ<�xD=�̻g��~�?X2�>�?tO{?�*�>��>�KY=\̗>���� *?xʿ>��M<��ʾ�X���d��y���K�������n��/IȾ� ==��; >W)<>��="\���r>��G=�A=Ʉ7�"�<˹�=�>5�>��!>G�1>�R>�Lj?� t�!��ژ/��ȴ��z<?!�g=��y�y��#\�>�J����1R������>i? 
�?�n�?G4?�	���U�>�����W���Ⱥ��N��@m�>TR�>3������>��	>\�EԤ��s=ކ�?�;
@05:?:���o�ܿ�>>��7>`Q>��R��L1�Z�[���a��Z�aM!?=K;���̾�3�>�.�=�y߾��ƾN�.=�6>ʾc=���Dk\����=��z�]I;=2k=���>L�C>�?�=�>���Ʒ=�I=�W�=r�O>&m�� �8�r0,���3=���=ac>I&> �?<M�>�� ?��?01,>�+��M.b�� ���jb>���<��>���`]<G��>�A?	M?O"e?Z�>���rB�>��>�l��Sj���ԾRic>�z�?bh�?�H?���<b6���H-���4�ļ���?�p?A��>!�L>���lҿ���PNH����ο=rO�����r^>�=��_���=�@>%��>'��>�c�>�>ȗ=�"?=�'�>�0>��=}n�;����!��Z�,���=$;U�u<.�(<T&Y<�&;W�k�kʏ<���<=���2%Ҽ˚�<�z�=���>��>���>�G�=8���->G��o�L��0�=S`����@���d���}��/�~6�dD>)�Y>�ԋ�(#��q?6OS>H[=>���?�Su?&>�3�5<׾�v���]f�X�N���=0�>j?�B�;�)�`���L�R�Ҿ�k�>T�>�A�>{`>k�(���=���~=���v�4�	��>�(���e������p�� ���7��T�j��/2���D?̈��#�=��}?�RI?�5�?+�>�m��j�ؾsm/>J��f�=��,�k��Ћ�iE?�/$?�U�>õ�!�A�ދ¾4�ý)K?�{���S��*��o�P�9ւ>�0�pb�>��Ҿ����\�'���������W�o��:_����>VP?lܹ?����3��}p2�Sf{���;:Xj�>;8?a�><��>y�>�P��3/)��Q��7�L<���?v�?���?��>+о=_���3��>�3	?Т�?䝑?@Ks?o`@�E7�>
��;i >����;/�=}�>"��=�p�=�9?l
?�
?MW����	�Q�+��]�u�<�0�=j�>���>�'r>:�=[[g=��=\>�Ȟ>��>�Be>2�> V�>dYL����=D?̚�= �y>J�?�m~>�ۓ���ټ���=t��v)k��1ϼV��:����"��=dWf����;6��=Y��>��Ŀ� �?��V>޾�?���$�#�ti�=���=̾�<�V�>��>�>��>��>�E�>�7�>+�H>��㾱�>C��*���l��ą�HT�e_�>X���g`����+9�܅���Ѿ5����ߧ����C��7ؽu#�?���W�YQ$�t�YX?��>F�7?)�w����e^V���?�S>��'�%ؤ�����d���X�u?g�?�hh>\�>��O?�8?������6�Z��tz��LB���k��\��D���V���c��ջ���^?�My?�aC?�B���q>K�?Ҏ'�	���V��>�+��\:��9=�i�>ǵ��^��h̾��ž S'�2<>]Ck?���?��?�DQ�cD�R��>�(A?Bb5?�,�?�>?��?ߏH�^�??��=��?>t?Z3'?^�?[T�>��>>�n�=��A=O��=�ԣ�*l`�s���4��i��.1=R8�=�$=���<��=�t��������h4<���<�j�=ϼ>�#:>��=�߮>3X?Iί>>��>�C?�
��9�<��r��c�?e'��W� h�ީ޾�{�Q��=�ae?��?�?e?Uh�=m�?�� �f��=��j>��>?<>f��>����Z ��s�<��=b60>�=��ܽ$m��!c�m=���=#64>�?��=���붳>.�C�V�1���4>�?V���h���S����ה��_ƾZ �>��A?�[0?,��>�K���#��R�0A_?�\�>�e7?s��?�͟>�z/���Y��F��-�����>tK�=� !�ᤫ�����R2��1L�ӎ><~Ծ�W����>@���Ǿ9x�fYl�m���F��=v3�4>�P���徐pQ��m�=>�
>}�Ͼ&W�k~���⥿s�L?b��<&s��w�u�0ĺ��H�=�>���>�������<�G6��PH�� �=]�>��2= ���r���Y��%��{<�>mQE?4X_?�j�?�$���s���B�Ĭ��Vg����Ǽd�?Lt�>�g?�B>���=Q�������d�hG�g�>G��>f��y�G��=���1����$�ō�>�6?��>/�?r�R?��
?M�`?�*?�B?h#�>�$�������A&?6��?��=��Խ��T�` 9�4F�m��>h�)?��B���>>�?۽?�&?�Q?�?"�>� ��C@����>?Y�>��W��b����_>��J?Ú�>J=Y?�ԃ?X�=>=�5�5ꢾ�֩��U�=�>��2?�5#?A�?ү�>yG�>�d���.�=���>�*c?�,�?��o?�"�=�	?� 2>���>��=�g�><m�>�?�DO?�s?X�J?%��>�F�<_��;��H�s��sL��]�;�I<Y*z=\x���s���?;�<��;+��Y�����D� 
�����;�>�dp>�ݑ�B->3�þ������D>����䝾1����x=���=v�>�}?��>ˢ$�	�=1��>��>���O'?�?�9??d�;�Db�a�ݾF�N�)d�>��B?]M�=*^m�妔���u���v=��n?��_?1�O�j����j?�8?�L�׾��¾몾���w+�?7U/?(����  ?��?)�?��1?�;���Y�W���q_������M��n�>Q(վ�@��ґ>;Q�>4�	>t�=�D��C��Ќ�҃˾�>%�~?�a�?vZq?#�=��c�T��0�4�����d?]�>����!�?ڌ����ݾ�3���ؔ��~���Ͼw���'���%�����%,V�
���.�=7�"?��?mT}?~j?�����q���g��w�&b����(�N��3E��5K���Y�D
�4%ؾ����=����F���p�?`n?�U��5��=�%�]�Ӿ�P%���X>}�׾@Q޾��R=E���/>Q�W<��N&�����ˮ>?��>���>��;?+���7f�:-"�]���C23���>���>�>��>-T��Hi��<~�F�߾s���*��5v>�yc?��K?�n?Vj��)1�4�����!���/��e����B>�m>+��>��W�t���8&�Y>�w�r�-���x����	�۠~=ͯ2?~*�>���>�N�?\?2z	��n���lx�W�1�菃<?+�>Zi?�>�>��>��Ͻ�� ���>f�l?4��>���>����"G!���{���ʽt�>�­>���>r�o>��,�A \��j��P��39��x�=[�h?����"�`�x�>FR?�$�:��F<�|�>� v���!����&�'�7>d�?֪=Pu;>/�žG*�>�{�E��t)?zF?1Ӓ�oo*�b%>�"?�6�>�c�>&�?V��>}�¾bI��+�?��^?�WJ?>A?&��>�.=����MȽc�&���-=�x�>�([>�Lk=v�=�	��!\�iR���F=�/�=gѼ�ι�ʗ<�����~F<1k�<��3>{�ڿ��B�An����ƛ�

�/9��9p�H���V���ľ� ӾZ�}��r�����8�����v�k�h��e�?��?X���ʎ�����3����g����>#����=�����t�p� ���Z��p�����-<���Z��YZ�M�'?�Ǒ��ǿc���J<ܾ5' ?O ?��y?��3�"�4�8��� >>+�<߮����뾆�����ο[����^?���>��>�����>n��>��X>V;q>P���垾j�<\�?�-?̓�>�r��ɿ���u��<���?��@{A?�(���8�S=���>��	?@>�11�5K�n鰾��>�.�?��??�K=��W��I
��be?j�<��F�:��=#��=*7=i���J>7Z�>�m��iA���ܽ�d4>ۅ>'�"�B?��%^����<�]>��ս෕�5Մ?+{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?'�(?5ۿ��ؚ>��ܾ��M?_D6?���>�d&��t�ޅ�=i6�����|���&V����=W��>^�>��,������O��I��P��=�#�Gǿ��$��~�U4�<=Wͺ��Y�;F�S��E�H������n�'R彜n=���=��R>�c�>F�U>��Z>,�V?��k?�~�>x�>��Խ}���}�;�1��Q���������9z����W�뾢s߾� 	�Pf����S�Ⱦ�=���=�7R�昐�1� ���b�ەF� �.?Gu$>1�ʾp�M��u-<�oʾaŪ����\ߥ��,̾�1�9n��˟? �A?���/�V����;��z��|�W?�T�����מּ��=�ű���=�(�>ȓ�=6���3��}S��0?�.?�¿����y)>����=��+?�|?��d<��>W-%?Z�*�����Z>�}3>���>X��>�	>s'���#ڽ��?>�T?;�������>�K���{�K^=�7>u�4�̪��d\>QH�<⹌�E�P�v���~��<�]?7�a>��-��������CEýXG�=G��?��&?��>��?�qP?�V�=�����e�	�x	廔.?��m?�e>H�'�=���Z6�.�?hV?�9�>a����Ӿ&M5������?,��?�K?w��=��n�����,��$x0?�v?�\��3��MK��V�e�>���>�>�8�]�>�"<?'+�ὕ������2��֞?�H@��?%3<(�4�=?��>k�N�i�þw���a���b=�U�>�_���	s��s ��A*��9?|�?V'�>�<{�mL����=dٕ��Z�?~�?b���*Cg<����l��n��Q~�<DΫ=��RH"����7�r�ƾn�
������߿�ɥ�>7Z@�U�5*�>�C8�M6�TϿ���[о�Rq�f�?2��>c�ȽC���N�j��Pu���G�W�H������0�>;�>}r���둾�{�k�;��Y��kH�>v 
��>�>��S�6������)l+<X��>�9�>0��>u\��㥽�r̙?�|��?ο"���8����X?�k�?�_�?y?^7C<Bv���z�u�$G?0_s?� Z?��%�?/]���6�#�u?Q��'��p���N��>>�.?�>*�����>��=m��>�I5>b�\�l�Ŀl8������`�?M��?��ξI"�>�Z�?�z ?����������D7�0?�AH>$~�)6�|9��%=��19?VA)?�� ��N4�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�^�>�?�*�=Q�>�o�=@#¾��.�M�>���=�	���?�-L?�	�>3�Q>�%ٽ�H$���E�x�^�G
#�0�D�iw�>K'd?�
P?5��>Cмɵd��'���
���:����>�*������B�F�8>��%>��>�y��7����,?�2(���ۿ�����H�EJA?Z;�>�s�>���`g���ٽopv?�A�>X>�f ��:	���~4�D��?;��?�P ?9����>t;�=�ќ>��:>�fC�w�۽]}��)��=�B<?��o�kt��M�x�v�<>�B�?Ԑ�?�|�?:nu��	?E$��K���j~�n���7����=J�7?�&�{>q��>z��=�_v������s�^��>5�?�s�?Ƽ�>J�l?�\o���B�8�3=bK�>��k?jf?�-w�X���vB>Î?�������/��'f?�
@^p@�^?�⢿f�ڿ񮰿�ľy�q��=�_>(��>.�c��6>]y�>c�&�ԍ�=5�7>���>��K>B�>m;6>��
>��0>'Ā�~�&�<e��΁����Ut�
R�kn���ľH)��4�C#���4��鱡;�HQ���-��jI�3e����NP�=j�v?:E<?�,�?�� ?��$#����Ӿ���<w���W>�H�>"�?�i?��E?u�=�UӾϏf�,�����ʾ�:4��j�>M>�H�>���>��>��=D�1>vق���Y>�M�<Ŧ�<�����O=Z�\>o�>:6?J!?�C<>��>Eϴ��1��j�h��
w�_̽0�?����T�J��1���9��Ц���h�=Eb.?|>���?пf����2H?(���v)��+���>{�0?�cW? �> ����T�9:>6����j�;`>�+ ��l���)��%Q>sl?Gf>W-v>��2�c�8�,kP�[��h��>�U5?8���>@�c v�x6G�N۾��J>��>�g��u�?���j�~��j�j
h=o1;?��?�I�����e�r�#𛾯^Q>QX>66*=�y�=j�L>�U��\Ž�_J��-=�+�=��W>sR?s:>�� =~Ѝ>#���2@W��x�>'�E>Z(>tWC?6!?)�0��ڝ�^ᓾ�4A��r>XY�>>kb>��T��)�=q��>��w>�"ܼ�N,����ò>��gB>J6��`e����N�u�J=��(��e>���=J�ٽ�/���=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�Z�>Hv����E���a��f�=k�?&�E?'+ݾ�W>�pP���?�{?ͦ��ݦ�I)ǿ'a��>N+�?)Q�?Np�����R�c��6?ݜ�?O�?E<����jI�Y7�=V�`?��x?E(�>����rP���>�Q�?Κ�?�I>H��?��s?�r�>��w�7R/��:��N���#�=��V;)`�>�->����QhF��֓�Ge��K�j�0����a>'�$=��>>\��?��&�=0���@���Df����>�-q>p�I>)f�>1� ?�f�>��>��=�΋��퀾?���.>G?�?ĸ���>�yi��J���G���_	?��"?t&������'�>ʽW?�h�?Y�U?Y�}>�������=iϿ+;;x��= |>o��>�X�>�4ļ�/>S �_>��h9�>_�>�b<�����a->G��>M?��>4ܽ%[(?�?���=�¢>0�	��6�P����>�7?Y�?�W�?��?�����*��*������[YP�/�,>�Lk?��?� �=�
��^[����m����Mm]>��?0�p?�C�=��M?��?J�\?.$_?�h�=�-*�j�����n�\�>��!?j�]�A�UL&����~?�O?���>p;��UֽQּ���w����?�&\??&?���Z*a���¾I��<�&#�c#T�Po�;�>D�м>ڎ>�}�����=�>�Ѱ=UIm�$D6�C�g<en�=f|�>��=�47�c�����-?�z��S{���=�eg��4�Yf\>]4>�c���
O?9>5���y�3v��˺����A��܏?���?,�?�YƽPsb��:?�y�?�?�\�>E���L��n;P�f��nP��(
����=_�>��<�%��Q���Z���3\���Cm��P�v��>���>5��>���>�;�>���>�듾�y>�i��ϸ��TA�����R�0�� <�k
�������6��{����ʾ�(����>��h�Q��>L��>L#|>���>;�>��ҽ#�>�7t>��>ș�>V�6>��=��=©���r]�EWR?�|���'������2�A?�3d?�N�>@�c�儅�*_�h�?"��?�o�?��u>�ih��R+�F?�>P���W
?�O;=��r\�<������۬���F�O�>M�ڽ�":��M�T�e���
?�+?79��?�̾�ݽca��}A�=2�?�$?ݑ.���Z�no�HfJ��BZ�1Q�e_���9��� �r�p�b���XR��Y���T*��NV=�-?�̓?���쾬���_�n9�5Sf>���>k]�>���>�O>"�	��6�L�e�j�&��M��X�>Ѕ~?=��>�J?I�:?�P?�L?Y)�>���>�B��V�>b����w�>/��>K�8?��-?/!1?�\?Q�)??`>$��ܔ��U�پE�?D?}�?I�?"�?[섾�QǽY��&�W�N�~�&���r�x=�N�<�ν�k��{_=�T>�?�S%��J?����<X>��9?v��>���>����� h��\H;���>�:?�a�>��� [w�D����>6X�?Ӽ΃�<$>'_�=	�;�<Ⱦ�=�]�_�=�0�h��!r<�۩= lv=����y���/;�ү<��<�i?$?�09>�4�>tXr��l��d��-�Χ�>�(�<�i>%��@���ŕ��RP���>B}?��?�G�=�_�=�W=>g𡾔�xܾ��������	?+�'?Z�>?�av?Lz.?�8T?+�>jtL��D���ե��#�c�?.!,?��>U��ʴʾz񨿲�3�D�?[?�<a�޻��;)�̏¾��Խ-�>\/��.~�r���D������������?���?cA���6��w�D����[��_�C?"�>Y�>��>U�)���g�M%�}1;>��>R?��>��O?�7{?s�[?�sT>�8�[-��ϙ�{�3���!>2@?G��?'�?y?���>i�>�)��(��i��zK����}ق�Z\W=�Z>C��>4#�>V�>��=)SȽo��w�>�wQ�=Qb>E��>���>��>\�w>b�<h�H?�T�>t�̾�3���	�� mW�6<J���T?;�?e^?�l_;��%�cb�?����>k��?͵?��<?��l�W��=Nt󼚺��z&��ȣ>RΡ>|K�>�v�=!=���=�"�>�C�>�W�V��Q "����/?�AO?cz=�ƿ߭q���p�PƗ��d<9�e�d�7����Z����=����؍�h���M�[�l���hy��s�]���N�{���>���=��=X��=#H�<�ɼ^3�<�J=��<fz=�mo�P�m<�(9���λ������\<��I=����Ҿ�v?ޚ>?��&?�Q?��t>�v�=.M����>���@%?'�t>�Ո��J��(�ཁ���Z���-о!�˾�TT����r�>��"�]� >��+>�8>����#*�=��=1��=��k=ځ(=�=��="��=�>�G�=�;	>�6w?����鲝�r3Q�V�Ӷ:?O8�>t�=�ƾw@?^�>>3�������b��-?���?^U�?��?�ti��d�>L��B鎽�o�=*���&<2>w��=s�2�c��>r�J>؂��J�������3�?��@k�??Vዿ�Ͽ�_/>�j8>r�>H�R�^�1�is]���a�(TY��g!?Z);���˾���>�Q�=A�޾@1Ǿ�g'=16>��_=��[��=I�x�9�B=0�p=��><0D>�{�=����7�=�B=�@�=n2P>S;��N50�R�&��R4=a��=~�b>��$>t��>l�?rW0?>Zd?<�>l�m�aϾM��iH�>���=�5�>�v�=m1B>v��>T�7?\�D?��K?v��>���=��> �>��,���m��j�`ҧ�ܪ�<_��?�ˆ?��>�^S<�A����g>�u�Ľ�p?�M1?p?ٞ>�*����6z��$� ~���f�<�R�=�H�d�=�EU>uǊ�-8��J>��>0��>色>0v>	C-=mI]>x�>��~>�=e3\�M->��F�:���4>��y���ֽ:�=�EнG_�����(�<9+<�O1=2�=�!�=��L>h�>Qu9=f�= a��2`�!�>ѫ��$;U�p�B=%H���(��4>�^"t��#7���^7>��>(ժ<���.�!?��>��u>�J�?V�?꧚>ֹI�B�'��ʲ�*�Ǿb����nD>o�>&�=��*��^O��>\������>�L�>B\�>G�Z>#-��^>�ٻv=�q޾m�3����>$&��f)�.����r�~礿�e����f�x��;>^D?�Շ����=��}?��J?�ێ?��>��h׾��&>���YC�<����r���j�Nx?�'?S��>��Q�C�9'���똽�u�>P�M��b�J��q/�P�>�^޾f"�>��¾c�����%�B@��i5����^�m@���>�-V?�}�?8;��1�����X�2	�&">��?�B??���>��!?e��>+þi�zQr=�np?͐�?F,�?{~e>�ͻ=���&�>�#	?_?A��?�s?�>��!�>�|�:8!>A�����=��>	��=#��=�?�>
?�X
?Dٞ���	�;���l�N]��9�<���=.�>�>n's>��=-ze=��=�]>u��>�v�>Y�d>�D�>�R�>�������;�A?�������>uV=?�8�>��q=�ˎ�2�L���B��b���ؽ|�/�i������C��ϕ=�E&�cM�>�	ÿr��?-�>'���ʇ�>���K�սB��>���>�`��v�b>\��;TM>:9�>��>��>� ?�,�=�Ͼy\K>��n��o��`��,������P�>>g����=M3 �Ҁ�������ʾc�#���5jw���L����<�4�?O�P�o�p��t!�CN
�R�?� �>�g*?3	8�n���E�=8b?F�->~;"����N���T����y?L�?d�>jJ>7�F?�N"?~�<�=D"3�����z$�Y�I��o�Nq��CQ��c�u;���ň?���?�[j?�uɽ�d�>F�w?h�o�^ >��>��UJ>��,��(?����Ja �j
���.��df�kT�>C�?|&�?�5?��ٽ�֤��۴>gx�>^��>�	�?�)?�f�>��'��"?��k�Q�4?xt�>�ͻ>G�?�rC?1f�>ϋ����C�
_�<ʐ����d�3���U�=��=!c>Q�<�(�=B�>n�&��q׮�W��H����仌�=���=za@>6��>�g;?�F�> ݺ>��1?_U����'�]��O?��L�Z�{�5\پ�E�g�#���>�|�?B��?���?X�x=���HaN���y>oh�>-��=^�N>�D>H�<[�N�cO�=pp>{iz>���=�tJ����p��u���S >��>5��>h@|>J ��+�'>�z��� z�?�d>>�Q�3Ӻ���S���G���1��rv�P_�>C�K?��?|v�=�c�Nq���If�6/)?�^<?KNM?��?:�=��۾o�9���J�9_���>w��<������U ����:��D�:�s>f/���ޟ�,�c>4
���۾�n��$L����)B=
���?l=j�҉Ӿ?y�"��=*�>j���e ��ږ��調�rL?�
r=w���S�Ɗ��@�>G$�>��>H�	Ԁ��?�&\���ə=�?�>��4>-�����ﾫ�F��e���>EC?�\?(��?-1���	���T�����k������<X	?[�>�g?��M>ґ�=�箾����~d���N�Ò�>�l�>2-���B�YN���� �*�NǄ>"9?>��=M�
?JU?�	?%�W?��?�+�>�&}>&T��z:��B&?2��?��=��Խ �T�} 9�GF����>v�)?,�B�̹�>F�?Խ?��&?�Q?�?��>� ��C@����>uY�>��W��b��'�_>��J?ښ�>y=Y?�ԃ?��=>U�5��颾y֩��U�=�>��2?6#?P�?���>���>f�����=��>Zc?z0�?q�o?�}�=I�?�:2>���>^��=ך�>Z��>?�UO?��s?��J?:��> ��<A4���-���8s��O�Nʂ;�JH<$�y=��t��L�	��<Ȁ�;TS��;F�����5�D��������;G[�>�5>-���>tݾe;����>̚=�8���o�Ӿ�������<ȗk>]�?G��>�w�����=�Ȓ>Q�>���� ?��?M'?4�����U�Rũ�C+��F�>l8?�M>�Fb����C3e����g?��W?f�۽�j��¬b?a^?��� �<��þ��c�����O?�[?ÅE���>�_?hr?���>�sh�U�n��1����a���g��=�H�>���:�d�CC�>�R7?(�>��`>a��=?=۾(�w�ą��T�?S��?g�?>��?��)>�n�� �R{���%��*3^? ��>U!���?"?$u�]Ͼ�䊾�Ҏ�}�?�������!~���ҥ�\W%��烾�p׽g:�=}�?�s?5�q?��_?(a��Td�rB^�"d��xV���U����E���D�h
C�Xn��n������>��3�@=�!��m:�ٽ�?��&?�L���>n���z�-4о��X>�♾���F־=�h�Bbs=�6=Hf��:��L��h`.?���>���>�;?��W���C��(;�x�7�����<>�{�>7j�>�u�>��<m*�2�νE�ȾC���O����u>�d?,�K?'�m?5� �	�0����1$ � �5������F>D#>0r�>�AY�(P�P�&��J>�}sr�x��D����	�L-�=��2?洀>]�>��?�q?aM
��ױ�s{�O�1�-�X<;�>�i?Q�>�O�>"ҽN�!�<��>�mo?�T�>'��>�Qc�G|&���r�̦�o� ?j��>)�?�H�>���mV�� ��6���J�x��=� u?�h����k��>��??ŵ =j�O<x�b>�i����1����v[��G�=�w?=;�=�Bl>�����	��m~��h��*Q)?�8?�򒾪y*���}>�"?�e�>\�>Q!�?Pٛ>��þR���ӧ?e�^?vLJ?�]A?�A�>�=����4Ƚ�&� �-=���>��Z>��l=���=�e��B\�z�2�E=�2�=�wμ�=���$<%r��HN<���<��3>�Ϳ�G5����Y���B�m� ��ƾ��0�D�'�6�C��$�$��mƽЭ��v<w݀���f�l����.��\��?��?]�.�U௽�ݝ��e����'���>x��L->�₾�d�|�=8������j�8��\Z�Bk�X�'?ں���ǿ����?;ܾ+! ?�A ?�y?��!�"�ے8�ǭ >eG�<'��8�뾒�����οI����^?x��>e�/�����>楂>{�X>�Gq>����螾�,�<��?L�-?Q��>T�r�/�ɿV���+��<���?*�@�dA?$1(��6�Y�^=���>��
?��<>"7�[�������&�>���?�ˉ?��@=wqW�I���f?�U&<��G�������=�Ԡ=�=����M>N�>� �]�C�2�ٽ�4>ϔ�>У,�)����_���<��[>O�Ͻ!*�����?��a�br�W�N������u>�4f?p �>_��<sj(?�-`�5:׿��R��Y�?���?���?'�?Q"׾�s�>f�˾�j)?��?�+o>a�4��`����=r�<<Un>����\����>�f?�Cw>0`:�P�(�؊��+%��s��=R� ��Ŀ�b��B�J$&=����s��A0ؽ�������U ��g5�� ��Z2�=N��=N|B>��z>:�H>!Q>�\?�Pq?��>PS->4�(� ����˾[�Q<b��\8��鉾:�'��㥾
߾��վ��@�̑�Ѕľ!,<�X�=X=P��v���!�*�d�_II�1x-?C#>��ƾLL�B$\<�%Ǿ���f_��;���˾9�1�o�Ѫ�?z�A?�8����U�F����!��zǽ�\V?Mi�����W��Ĉ�=�S��>=ԛ�>1ȡ=߹�%W2�f/R�!s0?�X?*{���Z��(�)>�� ���=��+?Ni?>$[<���>�%?/+���UT[>�3>��>�k�>t9	>T��� ۽��?gT?������i��>7��Q�z�>a=�b>_�4��O缧k[>�Γ<<ߌ�W�l��So�<hR?���>����#��V��\�1'�=�O�?��D?���>u�?�/g?!��=� �T�z��H"����#�Y?{Z?&�n=;��=�A��w�Ծ��5?
H-?���<ߗ���߾�95�	�	�� ?�a�?W�#?3����a���a��u�Q��,;?��w?��\��#��l�Xg�IҪ>�9?�	�>��@���>�)>?�96��6������I2���?ɪ@�1�?P�@=St����S=n��>���>��'�Oܧ��4���Aʾdy<�4�>w�����"���ӒB?6��?z��>B��V)�����=�ٕ��Z�?��?}���pDg<R���l��n��r�<�Ϋ=���E"������7���ƾ��
����ῼΥ�>EZ@�U�v*�>�C8�]6�TϿ)���[о~Sq���?M��>T�Ƚ����A�j��Pu�b�G�3�H�ť�����>7�>󦌽N���f/|��>���&�A��>h�o�>u�O�ޑ��1v��yQr<h��>:��>�݄>5����¾lݚ?y#��+�ϿX���j����T?�&�?�|�?��!?ߛ�;�$s�o�q�8��pKE?�o?sX?�H<��S[�r'��j?�]���T`�Î4��GE�(U>'"3?lC�>ޒ-��|=�>B��>�i>�#/���Ŀ�ٶ��������?��?p���>b��?�r+?i��7��~\����*�&�/�D<A?s2>���͸!��/=��В�_�
?�}0?W}��.�2�^?T�Bf�l�"��:�U�>�e-����_G���`��ƃ��H���?T��ܰ?'��?��?W����z1?�N�>P/ľ��'���>�I�=�yQ>Ł<<�]���>��X���?�W>)=�?���?+?7�n���y�Dx-��=O?F�>���?���>Y�>��>񥷾����\��>�b�=�>3C,?%�b?�$?t)��M����W�`(P�iA@��F後ZF�r6�>��c?�MD?��*>|�=�B#=9�vWľhy��G�S�]þu��/���=I�>��n>z�V>*5~��&��?^o��ؿ�h���'��.4?���>{ ? ��7�t����:_?
v�>l8��+���$���<�t��?�F�?q�?�׾8%̼]�>[�>�V�>�ԽA퟽B���e�7>�B?�1�[F����o�g�>o��?��@;֮?	i���?���3����Xp�7�&�u]��Vj�>�W?��K0�>RF?j��=͒}�������r�hM�>���?~��?�)?�d?�ut�?���#,�
-�>j�?4YQ?�.ٽK�H��&�>��>��E��J��4��ΰk?��@M�@`�g?����\�ֿϼ����þ�D�`����=-��=��i�=O>�@>��E<��
>��>�>�V^>Hf>4r >˚�=J�#>H���!���뺛�Z�R�J)��p�Y5���ξ�|�W� ���r�>٨�c�ν3_Խ��� I�D�,��s5���=��T?�zQ?�)k?
�>~����*>�9��#�|<��!�Zyn=���>��1?�1J?k�)?iԒ=P�����e��*��HC��m0���=�>�4A>l�>���>Җ�>��A� �D>�G5>��u>��>S= �E;�9=X Y>�N�><��>���>�C<>��>Cϴ��1��i�h��
w�W̽/�?����P�J��1���9��Ц���h�=Gb.?|>���?пd����2H?*���t)���+���>y�0?�cW?!�>!����T�-:>0����j�5`>�+ �ol���)��%Q>tl?��>}��>>�!�9g4�(�C�%����4�>� ?�۾�/�Ljj�'N�v1ξ�34>�q�>�����t,��n��&pg�S;d�zf�<DI?f��>��^�K*���1�K�d���>�A4>n<=�5>���>G}n�����n�f�J=�p�=��>�o?�K->W*�=(��>N���ݤO�2Ϊ>��@>D�%>w�>?�=#?L�+�������	O+�w$v>��>GKz>*�>�\J�ګ�=
�>b
^>���������	���:�g�S>�}���[�~�i�A�=�%����=$�=�%��B�;��>=i�|?(��؎����������:?�#?߸=�|�<����F����ƾ���?'	@��?>g־|wH���>�֓?�T����=>f��>���>�>��A����|�>2@�P���KF���o�?2��?��:�?���8�c��d=�,?`�Κ�>PH�O���䆿��u�[L=�>�eH?���~O�e�<�Ę
?��?�k�⥤�/�ȿ�Tv���>���?���?bn�����0@�ݎ�>'��?�iZ? �k>��۾mZ��)�>�@?u	Q?\��>�Q�g!&��?v�?�̅?�I>+��?*�s?Wo�>u�w��V/�2��/���k<=�\;�i�>\_>�����dF��֓�|i��9�j�4��#�a>gm$=]�>15住1���B�=y�C���f�k��>&q>*�I>jR�>� ?�V�>���>Z}=�c���‾Ҷ��l�K?@��?��)2n��4�<-��={�^�M%?�A4?k[���Ͼ�̨>��\?}��?5[?]b�>Z��->���忿^z��. �<��K>�,�>;J�>k.���@K>4�Ծ�5D��i�>�ȗ>ͽ��*5ھ(��l���G�>/f!?��>�̮=� ?	�#?tj>��>�UE�E;����E�R��>1��>`P?��~?�?�����X3����|硿��[��:N>Dy?�J?1ؕ>��������C�m\I��"��O��?�^g?ը�W�?�+�?U�??<�A?�f>���L+ؾ�?��S��>�#?<�/���H�=1���9��>���>7��>���Y��yM��)���A��(?m?�).?L�ﾃ�k��x���ұ<�y���;m�=���b:�=�K>2�<3��=��=�>&兾Z�A�g}�<�#y=��>4>�>���ٽ>,?7G��܃�F
�=8�r��sD�,�>2~L>;�����^?e=�Y�{�����y��9U�M��?���?qq�?�紽��h�\%=?-�?�?��>�T���x޾Y���2w�Dyx��f�#>���>�[k��徂���̟��bK���Ž�����>I0�>���>�}�>@KS>�ڽ>�ǚ�U`,��z޾?��S�`�Uz�e�0���$��q������X���u��hm�z�>M˽~�>[��>=�}>��>�(�>�G�����>5�f>׽�>陸>z�k>��4>�_�="J�;v���9HR?F)���(���u^���}A?Wec?6��>�cp�O����s���?iZ�?��?Ŷy>�vg���*�m�?t1�>h���3
?zt3=�n����u<�������셽����>~�Խ��9�M�L���d���	?;)?[����̾ؽ�X����r=J�?��(?�<*��R�K�p��sW� �R�zP�g�����9 $���o�3���c,���D�(�R�=��+?��?���� �)����pk�A�?�<>e>��>a��>Nľ>I�J>�h	�Gm1���]�<�&�_'��9��>�z?��>0I?:�;?.�P?�WL?D��>=a�>(��<e�>P��;��>��>ٜ9?��-?-:0?z�?�u+?�0c>Tt������Szؾ�?f�?6I?�?��?Ѕ�[Pý�X���He���y�������=/h�<��׽S�t�:�T=��S>�R?f�nj8�q����#j>�B7?-��>�I�>����S���g5�<A��>W
?��>���o5r����8 �>�o�?���$=��+>�k�=7ڃ��>�p�=I���@�=�h��8���0<N��=�ϓ=��0�S��8tZ�:�xt;d��<*�?I�?+�=s��>8����Tu� ����>�?�>���>��>sy�𐿣H��P�f�o�>8��?�n�?w���`�=�L>*K?�D�t������� x�= �)?�P?E�j?���?�@W?M25?�>�=�)�ދ�5{�~���1)?q!,?G��>�����ʾ]�W�3���?PZ?H<a�$���;)�l�¾n�Խ��>�Y/�0-~�)��_D�U���.��q|����?c��?�A���6�/v�\����Z��|�C?"�>�X�>��>��)�b�g�$�<1;>,��>�
R?vK�>z�O?��z?S�[?oT>��8�!.��ܙ���>�# >}�??䎁?�܎?�Ly?;�>�>��)�gu�����d�������[\=f�X>)�>T!�>!�>u��=c�ɽ�u���@?�:p�=c> o�>�ܥ>L.�>��v>Rܬ<��G?tC�>N���n�B�s��d�/XR��χ?�w�?�$?5�k��_�e�c�%��J��>s�?1ղ?��T?t?b�yG�=�
a��˾|���>N>pދ>M0�>�!2>!�]>y��>�o?&r�>G�s;�4���;�=�x<pq?qT?\;>��ƿ@{s�ťv��#��(4M<������h��2��nyI��t�=���P�������U��ݜ��S���ɴ��[��=�~��e�>�Y�=�J>}��=-��<Z_ʼ�p�<Y�b=�Z�<�)�<���X<��7�Xa��ㆽv6��0<3�V=¥'�lԾ�p�?;�?��?��Z?��>�y�>�s>NZ� ǳ���?� l>*�<��������D:��1
���߾�#!���^�2���xs�;�Gy�t>Me >�؏=��l��P>�Ȗ=G�*=�"��6�`��=�H�=��>�$ >JP>a�i>�>{?Hy�B�i����YF?�?�<���t�W?b�>ͧ��Ŀ�]��u?�N�?�?(�?���<�4�>��T�ֽh�@�'�޼{ra>@��<������>
z�>�KV����2�<Q��?�`
@^�S?�n��#�ɿ٣�=��8>�8>�R�Hl1��:\�7�a�@HW�L� ?Ư;�%�˾��>�'�=�޾�-ƾ��0=��5>��U=�2��[�!�=Ǽ���J=?d=��>�B>}P�=ꐭ����=�E=�L�=��P>\ٺQ/6�]"�0�:=�6�=\c>��$>iw�>{i?Ձ%?\^?�r�>t@�x�پ�'��=}>�k=mޓ>Xq3=䷏=;��>�-?�u>?��R?x'�>���<S�>�>��#���i��& �"�ʾ79<=rs�?��??��>x��<N�X�d��*�3�f����v?ݦ-?f�
?���>���o�ֿ��?�84���F��d�<��]�b���>~/ �6�߽�)i>7��>C:�>�>��
>W 5<g���0�=Tֹ>l@�=�)�= D#>_�=e�I<�jۼ���=����z���μ൅�z�<;��;��!=ڢ<�*49Ӈ����$=p0�=B��>\">W�>K��=����2�.>c���V�L����=\ͧ��YB�Jd�U�}�(�.�st5�JB>�V>�t��5���?�;Z>�D=>tY�?n(u?a >B"��@־�ϝ���b��&R��=�>��=��u;��/`�h�M��[Ӿq��>9.�>�>/�l>=�+�!$?��@v=����.5��H�>2��On����)q�e=������"i��3���D?�B�����=�(~?ٟI?�ȏ?֔�>]Ø��qؾ��.>X[��A�=R�^q�gX��@?�'?`��>q쾩�D����o���x�>��9���T�������6����=����&�><݉�%w��2�'����=͐���@��J����>afT?:&�?PG��Sr�\$T���5==e�5?t?�`>�  ?�]?i��_��D����u&=��o?%��?���?]�a>̈�=萳�G��>	?���?3ԑ?�r?�jA��*�>��1;I >����	�=t
>��=�S�=��?��
?73
?�Ĝ�ˊ	��J�"�񾒴^����<�Ѡ=�*�>��>��s>�x�=�Sh=�0�=�\>�Ҟ>���>b�d>&l�>ݐ�>�[�1���%�.?�?7�FՌ>�?o8�>.~�:m�a�'�;���zw��|���HFp�kvB��:�=
������C
�ע�>5Hſ�2?�؀>F宾l~?Yu�]4E�J�r>{��=��x��a�>fqN>�z�>,=�>�Y�>&�c>��>��~>�W���!)>���Bb���@�ǈ���8���T>c��F���ӫ׾E�<p能@����~ �"�]��r�@�5���I�;}�?��h��)���J-�PrʽY=�>M�>̷K?�q���Y���N>�9�>h�>�`�䠿�׀�HǾ$֊?k\�?�8�>T��>cB?
b?M�q<[%a<	:U�P偿��I�(�o��O^�AV��S��K��+��Ru[?�;�?�Q@?�޽�Ua>��o?7�#������+�>!�O4�4̊�]�p>�돾��`�o���g׾��m��9�=r@J?o�m?�@?�#[��<Ƚ.[P>^WB?�Z,?�Hy?~3?��0?�}��G?�/T>�3?��?n/?`
#?��>Ơ�=�n�=�4&=��=�都��|�vm��A��t(���A=�K%=��a<�z�<�X�=͌,:a�Ӽ�Z�;E�<y-����<��=f�t=t=�=7�>G?��>A�>Be?m�>�7��=��y�>N���x���M��X�����	��([=)�`?�?�$Y?
g2<��/��g�)��=��<>�2>�f]>yԖ>؎���e��c�=0t)>ֵF>�xV<!߽�jv�)�I���a*�= 3>:�?,�=�f�r�
?���>`��Ȏ$>��S�$ߚ����#�]��VN�S��s�'?��@?��??��\>���_a�=Q�'��jQ?S�7?�R?Æ�?��>������N3�\�X<���>�[�:�9��@��b���&&���=!�1>�k��{��6B�>��U�<^�����bX����^=�=��8�{�>~h��͙��ߒ��:�=B >���2��_
���d���b?f��<�xžƦ�;Iܾd	�=恠>Ǡ>�j��P�:m#��1���=��>+G>����C����<��c��߆>PcE?��_?oU�?��҉s���B�2<���)���Ѵ�z�?���>��?��A>ꛭ=�����PGe��QG����>�C�>����G��i�������$�vv�>�?�>��?��R?\�
?aa`?� *?k�?!3�>���:鸾�L&?R�?�:�=f�ս�wS�Ȥ8�u�E���>�)?�C���>k?V�?�t'?W�Q?��?�a>-8 �x�?�HZ�>֤�>��W��`��i�`>�J?��>ܷY?��?WN=>�5�r����4����=�� >��2?�"?��?�z�>p��>5�����=Z��>Rc?0�?>�o?��=��?�+2>���>,�=O��>M��>�?�XO?��s?�J?��>���<�&���:��**s�[O���;K�G<��y=����Zt�3R�x��<���;����^���x���D�p����;���>�it>�B���3>O¾k��$<>>����4��o���q?�d�=B�>5??���>`!��/�=��>���>���m;)?,�?��?���;�b�پ�rC�z��>.MA?�k�=�/k�����@v�M�U=L�k?]?�+Z�������b?��]?se�=���þ;�b�F�龂�O?��
?��G���>��~?�q?���>��e�&1n�����;b�s�j��ʶ=rv�>�[�Y�d��C�>z�7?�R�>rc>b_�=�t۾��w��r���?���?��? ��?�*>:�n��3�o@��F��{�]?`�>Me��#5?����� ��mLP���K���˾v=���#��ܿ��x�����%�?Q���H�!4>5H?yo�?��? Ep?u羅j{��\�D�e�$�t����$�"�9*G�BX8�G�9��<d�fu��f�Ǿ*�<������cn�?�l5?g%����7>C׾��ƾZ���7��>�Z�����5�>蚔��>�<���C���\���̓�3�B?\?ō?;�%?<���Ru��I+��3'��-��ֿ>e�l>�Z�>���>��K=�^�G�^��i��[,Ⱦ.!���p>K�e?��K?�n?�b�/����}��
b�0�����K>�Q!>�Ƌ>�'Z�b/(���(��?�[r�=�����w	�s=K1?�A�>r��>L;�?��?���ѱ�S�|���.��<�<�ú>��i?�I�>\�>JB½u��`[�>��r?�9�>ص�>�9�����~[�o�/�1�>pϜ>$�?P��>�!&��QR�\��)x��}+���@>�^L?8���(Ľ0<�>R_-?:�T��>=n�o><-z�f[�ᑼ��� ���Y>^*�>'�=�9T>��ǾUy �ݡ�#���-?xF�>+�����2���>G5?�P�>���>왓?��s=�>)�jV����?�5j?=4�?вg?��=m�>J#���p���7���Y=��/>�<�=�� 9�l*�1������i޽�'=-�C�Xo�xx��T�=49�=3x�=氲�
�=]ۿv�I�SXξ��
���
~
�	��fæ�9��	-��rs��������m����T�.���V�C�j�l����RY�Uz�?E��?�O���'}��Q��Qق��` �v��>�#��؉'�����G��,����޾�����#�3M�z�j��6d�R�'?�����ǿ����;ܾ-! ? B ?/�y?���"�͒8�� >3E�<�)��l�뾜�����οF�����^?���>��
/�����>᥂>��X>CHq>����螾
1�<��?Q�-?G��>�r�1�ɿY������<���?)�@pzA?��(�E��q�V=��>��	?��?>�Z1��I�/��Md�>�2�?���?K�L=��W�y�	�$�e?^�<��F�]�߻�;�=�T�=eR=�����J>�:�>X��C@A�Xܽ8�4>]݅>|�!����^��t�<�W]>��ս�E���[�?�D\�zyv��K�ԩu�U�>^t?� �>*�7>��.?[�e���пk3L�k<�?��?�+�?{4?��b��>T�׾F�?�1?�?,>��@���~�D�$>��g�Y��N*����q���>��=?h�W>H)�J��!V뾂�4����=�������^��Ɠ$�����C=r���������=z,�<(�8�ٵ��������=�q�=$�8>�(>��P>�o�>*L?\�|?:a�>($>�F�a�þ�AԾ�g�=�Z���=�w	���Ic�[$��>��B�о�����,������=���=5R�)����� �N�b���F���.?�$>`�ʾ\�M��?-<kʾ��������ӥ�*1̾��1�En�Yʟ?��A?����~�V�_��Ya�g����W?�L�����㬾H��=cر�-{=j"�>L��=E��o 3�rS�� -?��?�Zľ��m��\3>�����=��3?|�?��_="��>�?��-�})��/I>�z+>�y�>B˾>��=�W������o?@uD?�X#�$Y���2�>;Ɍ�����O=��h>�� �	��}�I>������\�: ���h&W?Ҡ�>�)�(���M��;����==��x?ׅ?�>Gk?��B?���<x����S��>x=J�W?f#i?��>�[����Ͼv���5?�e?��N>�h�Q��g�.�S�#?c�n?]?II���x}���"��e6?��q?hJ�Sq��5��x�<�C��>�?��>�WG�=�>�JF?&�[��ՠ�d����'���?Q�@��?�M>�-�_��=�z�>lV�>�	��@�c���+K;M>�=���>Aހ���S���������M	?�?��	?k�x�׾'��=�ԕ�%\�?��?}����f<M���l��o��!�<�ū=��*"�����7���ƾ�
������������>=Z@��A)�>�[8��7�zRϿx��Eiо!7q���?K��>ĊȽv�����j�Qu���G���H�ȯ���ϫ>D��=8���ꟾ!Jq�^�*�|���n�>�+$<��b>k��anоH޶�j��<`�>���>�(�>��ƽx¾㋒?��Hɿ ��eF��KQ?$�?�e�?k�(?�>{��R������b8?k?��G?Gx��E���.=�j?2_��fU`�s�4�HE�!U> #3?>C�>]�-���|=u>2��>+e>�#/�^�ĿHٶ�����v��?���?�o�1��>R��?�s+?Mi��7���[����*��,�<<A?�2>����ָ!�0=��Ӓ���
?~0?{�Q.�ܷ_?�a�3q�{.�aȽw�>̲,�4�Y����_���te��@��{�V�?�<�?��?���e4#��%?sޮ>����ž�P�<c�>��>��O>ۈ]�)}u>EX���;��d
>��?BI�?'g?䒏�A��'l>J-}?ה�>�B�?�Ad>=�>��^>�$���*���RU>��:��ǽ�y?<�d?��>���ʾ��S���R�N��!��d:�#TY>�G??1�+?
�'>�׽�:���Y
�ln��p#��!4��� =9O�өv>tG>e��=�`������?Mp�7�ؿj��yp'��54?U��>�?$��_�t�����;_?z�>7��+���%��B�^��?�G�?C�?��׾�T̼�>`�>$J�>��Խ����[�����7>&�B?���D��Z�o���>���?
�@�ծ?Mi�&�?�y��ݏ�@݆�[�2��x�O��>��9?����	h>�_�>�U��4��d���`�%�>Nb�?2�?ʬ ?�xq?����~md�P�=/��>�ϐ?ZX"?��X&�	��=���>�>D�k����Ծ��e?J@{?@�7g?������Կ}���9�;7�ԾU5=�n-<��=�^$��^]>Jc�<�O.=��=�(R> �>6^>�bE>�>!>�!%>��>���v�"�"b��%���1V�%<%�����w�z+�yƕ�AA��`���씾���QѲ��F��K�K�q��{A߼�
�=ҜV?J\Q?��o?
� ?;�z�Ѓ>�\���V�<��(�ֿ�=�͋>��1?nJ?�(?^��=����d�;5�����������>J>���>�x�>�>��ҺEI>۷;>\|~>]�=ަ*=�~;�\-=w�S>9W�>���>��>�C<>ő>?ϴ��1��_�h��
w��̽2�?����A�J��1���9��ͦ���h�==b.?
|>���?пa����2H?/���j)���+���>v�0?�cW?��>0����T�J:>E��}�j�l`>�+ �Zl���)��%Q>xl?f�g>�fv>�M3�EA7�o�O����	!�><�6?x����6�C_t�$H��Rܾ�L>Ľ>��=� k��ܖ�4�~�U[h��Sm=�:?��?��������t��	���M>��X>D/=࿨=�O>kL��ýc�D���6=���=�]a>3�?��>>���=���>�,��]�P��>�F>�)>hD=?��#?S8�����S膾o�A��t[>Ғ�>��}>�A > ;Q�+N�=���>y�T>�=���w����kQ-��IH>��c�.e?��:�yx=����0�=�v=:i��S���<#:|?yߥ��Ӈ�z��!���w>?�T?pz�=���<Z��ZҪ��H�����?ʅ
@AX�?�����L�=�?R�?����=#�>��>�y���^i�V�>�y�Fت�'��1i��?�v�?H���w	��'f��?�=�+?���id�>jj��S��z����u��#=���>�8H?�]���5O�i�=��y
?�?�e򾠨��n�ȿ�vv���>��?���?�m��D��)@�O��>��?�fY?=si>�S۾B�Z�ӈ�>߮@?Z�Q?��>�=�tr'���?��?`��?%cP>̄�?�pj?ɜ�>�0�<�����z凿��)=3�;e�>�6>�ȶ���B��㘿�8���,b����@>@�R�!y�>1Ƚ�þ���=�a7�f0��x���m��>��D>�>�l�>��>9��>m�>�?,=(���@��
�K?C��?c��*n�n��<��=�^�.-?�F4?� [���Ͼ�ƨ>ɴ\?.��?p[?�f�>��G;���㿿�y��J�<��K>�'�>�<�>`'��\CK>6�ԾYGD��e�>�ԗ>RJ���8ھ����ޢ�LC�>�d!?ۄ�>�ٮ=ז ?�#?}�j>r�>`E��9����E����>^��>.L?��~?��?ѹ��Z3����?衿ߍ[��,N>��x?�T?�ĕ>鏏�����g�D�<�H�B㒽0��?Itg?d�彠?9-�?O{??&�A?f>�y�� ؾ]t����>��"?��G�A��$�[��E?3 ?M��>V�<�r	��eݽ�� ���Ҿ��?3�f?�<.?�;�[�N�*i��y/�<Q	��Ԑ;�0.������>V��=_Ҵ���=��>x�=#���IW����M�=��>D�>�~G�8Ɩ��,?ow�<�A���**>�P�9+�i�>@q^>��վ,�.?>B)���j�ʬ�ì������ȇ?=�?�z�?c�d�Ԫ^���:?��?��?b��>$ݭ���p��ze��A����N>���>��.<3N�J=��+K��"�y�#"�ir�U� ?���>>�?.�?��K>N̮>緜�1$�
�辅���jT�=h�>�6�(6��� �������L�u6ľ�v`�p#�>ĸ��M��>��?/�]>�{>s��>�]�<a�>�e>^~>ϣ�>35Y>p�>���=	���wWҽ��Q?p�����!�l��'��N�<?KZ?P��>�+��������2I?I[�?��?^x�>�EH��c1�`h?�?Lu�`?��5��"���m�=����_&��Hԣ=	�=��z>��`��3��jC��΂��:?͞?�U��h����B��ʠ�$�q=�{�?��(?&$*��IR���o��dW��:S�����$h�����$��jp��Ώ��^�����(��Y*=�*?��?�H���ֶ��0Ok��>��5f>�&�>>w��>��I>��	���1���]�K^'��e�����>��z?ы�>��I?��;?xP?�iL?���>�b�>�6���[�>e,�;��>���>��9?��-?�30?&y?�m+?�c>�D��I�����ؾ$?�?�J?�?�?����m�ý��&;g�e�y�13��Y}�=���<��׽k�t��U=:T>KN?�����8��D��[�j>N97?���>S@�>C��!ـ����<���>�
?[ �>����yNr��g����>o�?{��	t=4*>7�=����ƺĺ�D�=�X¼ �=�ǃ��8��{ <�$�=T�=*2j��-X��i�:�j;��<:�?�#?x+A>M��>����g�ʾ��վ�ͼ L@="6��8�>:��Ά��k-��o.��I
>(�?}{�?D�a<��=$�>��>,��SѾA^����z�aP�>�?\ d?��h?�G6?�:?�<�>@��̩��ɒ�{��/- ?�!,?"z�>/��b�ʾ�񨿭�3���?>[?4a�ȗ��C)�p�¾��Խ��>�N/�Z#~�c���D��������l��^��?n��?��@���6�Ƅ�\����`����C?��>�m�>�+�>=�)� �g�)"��;>ϔ�>�R?�q�>K�(?�w?��i?��>����%���L��h~콠��='	-?�s]?�:�?��?���>�)Q>�_'�	�¾ǮF�BԽ:K� ��0���+�% >CY�>�<�>ꂶ>�/>��<�ع:���j��?�=���>*{�>nh�>�>�d�>W����C?�>�ܾ~*�׽��ײ����>���?��w?V#?��=�o1���q�-�����>L#�?U�?�M?�����=g\�=�оmt�����>^��>��>��>�P)��N�={�:?�?eV��/4���S�@���i/?1r?��S>i�ӿW����zE���h���D�6�f�Uf���]>�"d>�`���=�2=��J����u�ݶ�%ɾJJ-�*���Ų
?cU�=%K&>�q\=؈#����=���=��=�0b=s}�=^��<@�U�s�̃߼)f+;u�T=�X�<�f�=yG�=�x����?V>?��R? �J?�H9>�<�=p�n>Y2�^ET�1?m�?��=鞻��K���#�(�>��4��Д�	���*Y�=Qk�=��>7>�B>྇=X�[=��~=�"�=�ɠ���=��>�e+>RW2>�++>��=�>"cv?3�w��;���BP��Xʽl�c?�p�>�'�=!򦾋�3?�t#>:����-¿e7��6_t?���?ϴ�?�o?�9��^>=���~��2d�=�����>F{=����]�?�#\>�Q2�����q�\=�-�?�L@��?�?��[7ҿ;:=�=>My>cQ�T&+��8Y��i�bv<��L'?��9���¾O��>D��=~ھ�aľ��=�x1>)=�W-� �[��V�=����n=�0Q=G-�>��C>/��=VJнDڃ=�=l��=�D>�$'<iӅ�:j��V=���=�X>\�->���>�_�>^|"?{�P?s��>3������k�m>�#ֽ�o>ǽ6�$��=O�>�i9?�C?�!9?���>��M��>.ڑ>8�\���0��b~�$�>){�?Wh�?I��>�<
�����-���Y"�E��<���>�+�>��?�B�>���5�ۿ��y�/��/����m��꫾d�>������:�	>�s�>la�>!?�>�`3>^=�=>�K>�&>��>�pK=6��=��7>�b��Ϗ=��<r{i;Z��=�f>��u^=vu���=n��;�<@pZ�g�ڼ��6�WZ�=W��>��>g��>���=�ֲ�M�/>P)��QL��*�=�Τ�D A�W�c��~���/�N�8��&C>t�Z>�E��D�bX?�\Y>E=>���?Zht?is>F`�B�Ծ�ꝿ>�f�%�P�'��=J�>��=�:2;��x`�1N��Ҿ���>b�>:�>v�l>��+��?�"�w=n� ]5���>�h���f�&*��5q�
A�������i�.˺��D?�D��<��=�~?�I?�ݏ?��>'A��vؾ@0>�J����==��q�w��y�?'?.~�>�&���D�������p��>�奾=�c��L����)���=��پF�>;���!�����,�5Ή�����Z��:Q����>~�`?�?�,��	���b�@�l�ᾡs�=�L?�CV?/�>h�c>�)�>���BY)���ȾDŻ�o�?U��?���?h�.>���=Md�� �>�(	?��?���?Ds?V�@��>��`;��>����$�=�A>s8�=�W�=�?�
?�?���\�	�F���)��b]����<��=���>/�>��q>�X�=6<f=�̢=5\>&L�>^��>~#c>��>P��>�J���澸�?�L>RE�>��?���>`�c�{��06=Fۼ11c��Rx��G[=؊���n�=u��,�8�>�M�>\�ȿ���?���>̡��Z�?�#��h־8�>�*�=����z��>��>&�?���>���>ka>���>��>�xžPAO>��5�$��3l��́��"�=�>���>�'�}H= ��(�����2�}�NFn���`�o�ж�?7�T���%;��i<��&?��>��(?%D��$q��A>OG�>o�<i�s'��t鈿ץ��$�?y��?ռi>.��>NV?�F?d��(�#�c���z�`)?��~l��d�Л��� ��]���s���_?�&x?K:9?����s>�	z?>W#��6���:}>�)�r5��M�<>�>w��I�Z���;��ľ<y �;�A>��b?C�?��?�Z�0�m��1'>3�:?��1?�Lt?<�1?Q�;?�����$?k3>�F?np?2K5?{�.?�
?��1>��=/ݪ�	�'=\<���t�ѽ�zʽ�����3=Ȁ{==���)
<�|={1�<����`ټ(V!;2$���^�<_*:=�ܢ=�&�=��>��M?m��>o��>&<?#�ͰL���Ծ�>?ax��6����������L�>��h?<ը?�LH?�=fV9��~>��	>݊m>�4�=��Y>��>3����#�Z�=D>f�>��f=�I���|����^m�R�=�V�=�?�f�=���~>Ԃ���tI�� �x��ZnK�$.x�ܤt�� 3�������>-G?��5?��&��Ϸ�y�=�mF��v;?��*?`�z?��?�Z���i!��E ���(��	���z�>��_>]B*���s�����7�7Fc=���=~��x񠾈�b>���J޾?�n�j�I����J=4��qzT=� �P�վqu~�ާ�=��	>������ �����Ϊ��J?Uk= 4���U�<}��/�>-��>��>2�:�C`v�Bd@��W��Cۖ=�~�>��:>�y����RG�X:��*P>�_?�I\?J,X?H*�(�c�J*������ɾ����`?2�>��"?���=D�t=�U׾��&�f���{�h��>R�>H����b��U���վ<e˾E�>���>4�[>s�?��|?�v�>#h?�<?��??�#�>-�x㲾H�!?�Z�?�>���aI;��Ay�k��>��?#\
��^�>��-?�o!?	f&?�%7?~�?k�=j��<�c���>��,>�%T��O��/�{>��P?�ݣ>��@?]��?:�>�	2�oL����>�z>��>?oF.?�J3?B:�>p%�>A���B9�=�i�>ܬb?t*�?g'q?��=9#?�34>̆�>
\�=1��>���>�+?TN?��s?ؒJ?k�>1�<[V���D�� s����w�D9K;Z�<"�=u���q�
���<Ig(��!ȼ-�����nE���f���<�^�>��s>����0>��ľ(M����@>����Q���܊�S�:����=邀>��?(��>tR#���=���>�F�>����8(?��?>?�#;(�b���ھ��K���>�B?}��=�l�e���z�u�v�g=��m?|�^?�W����,�b?�]?�g��=���þ�b����:�O?��
?�G��>��~?m�q?!��>��e�
:n���.Db�X�j�qҶ=.r�>DX�}�d�k?�>l�7?�N�>h�b>�&�=0u۾�w��p��/?��?��?���?�+*>D�n�(4࿠]־�@��T�O?\��>�I��^�-?��<�f������ᠳ�����������hz�K����ͽa	���;!�P=���>�"|?}�R?|p?���,���M�h�B9��O#e����������5��`g�Ӓs��$�Ҳ�]1���	>�I~�ƈA�[�?�p'?��/�ˁ�>A��c��~;(/A>y������P�=��p�;=lA]=�$i�K%/�8^����?GҺ>���>1!=?�n[�v�>���1�
<8��~����2>�H�>Dȓ>Y��>ȧ��7/��
�K�Ⱦx胾.�н�5<>�Zc?�~=?��[?���|b��y�Mv.�$ ���ZԾ{�>�s=�s�>I��]�P�?��=�0�~����cD���������=�� ?��8>�{�>m��?��?�`��xþ�A|�:�A��k?>�|�>ů]?�Q�>���>B"�XJ�2�>Pwe?�Կ>�H�>�̇��q�r����iҾ�)�>p~>�k�>��}>Uf��kY�p�������DF���>4�?䃚�\N��S>ޒ4?qC�<���= ��>5�=���p徇Sƽ��=dO-?,���[m>#|��6k��y��bZ���3.?n\?��v�h/$�0��=��-?��>^<j>Ӕ?�?y��:�b=��?��f?zB/?��8??��>��=_ �?$��3�:�
[P<j8�>��W>�O=��=j����� ���4o(>�K<O���}�B�P�)>�6�=t�=ȝ�>"�⿊�>��Eھ�P�"����	V�����틛�b!ս�ꭾS�����U�L���?5����n����=R���ӆ�K��?���?�R����>����v�`��@>�ͬ������[�r�an������Q���c.��J�
�c��Y�P�'?�����ǿ򰡿�:ܾ6! ?�A ?8�y?��7�"���8�� >RC�<�,����뾬����οA�����^?���>��/��q��>ݥ�>�X>�Hq>����螾l1�<��?6�-?��>Ŏr�1�ɿc����¤<���?0�@*A?<�(�e�쾎�U=���>5�	?�?>'1��B��ܰ�/I�>d9�?��?� M="�W�^Q	�B�e?0�<k�F��/޻���=~��=�=����WJ>gC�>����SA��sܽ�4>�Ӆ>S�"�����G^���<�U]>� ֽd:���,�?�m��m~��'���m��>�?�$�>y�A>2/�>�d�a����h�%�X?��@�5�?ѷ�>��׾�:�>�3߾օv?��F?W(R>I�H�-c�×;�\����ҽf^;���K�hr�pI�>�z<>M�J�����H땽y&�=��3>�N�����.���"�9Z���I`����M�ν�ƨ��ݕ�����+ag�/˽�j�=��>I�%>�(>*&>
� >^O?�s?��?�h>ԛH��͇��
��_R��������$n)�P�$�G���~�ɾ׾A����!��X ��̾6!=�\�={6R�D����� �-�b�M�F�#�.?ft$>9�ʾV�M�8�-<�pʾM���e؄�%ॽe.̾D�1��!n�)͟?G�A?b�����V���UU������W?CP����"ꬾ[��=@���N�=�#�>釢=��⾘ 3�~S���1?�'?�ʢ��<��s�=~2���1�=�"?��)?�Q>!A�>L�$?�����EM�5A/>շ>>��>C��>�>ɶ��U潑?&&y?�Ž+�e��>S��t~�S����A/>z�Ž�li�[�,>�O@=62��6�J�,��~g�=�(W?͛�>u�)����a��.���Z==��x?!�?�.�>z{k?��B?;פ<�g��\�S����ew=��W?*i?ٹ>V��� 	о���#�5?1�e?9�N>ah����g�.�U��$?��n?�^?�z��w}�]��c���n6?T�|?�h~�G���9�tx��;��>���>��?~���U
?��8?�4h�H�x�/Ŀ}�?�eP�?y�@[��?�j���,�3�罿0�>��>ܠ>����bJ���y���#=���>����@��7������>?�i�?��>��վ]�����=_���Ȩ?>M�?�妾X��;��'�e�y��<|A�F�|=ʏ����[�q:��o�9�j��]���_���	����>�'@���T�>W'$�� �D�Ͽ�'��U�澨#y��s?l�>M��$^����d�~�r�4X:��M9�F-i�3K�>�	>�l��X���o�{��q;�����>B����>��S����|���5<@�>j��>�>�������Ù?�\��{9ο������]�X?Pe�?�r�?�v?p:<��v��,{��;��2G?�s?1%Z??�$�$]�S�7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�b�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�8na?+e�_Gt�P,�'ᦽSU�>�h4���H������E���e�R���E���W��?t @�?
�%��m#��#?�I�>����� ���s=m֒>Ny�>x:N>��T���}>���=����=}��?�4�?di?&�������B6>8~?B�>��?��=br�>��=���,�E�">���=�wA�r?aM?���>�K�=}%9��@/��NF��PR�<���C��	�>��a?JgL?��a>⼹�E=1��� ���ͽ�/1���|'@�.k*�Y�߽?Y5>ܛ=>�>�D�4kӾ��?2r�8�ؿ�i��zx'��74?"��>;�?*��[�t��M�w>_?�u�>S8��+��-$��S5����?�E�?8�?j�׾Fn̼%>���>P�>��Խ�埽]���U�7>��B?���A����o�/�>7 �?C�@�Ӯ?~i��?>!�V����샿6P�Q�=�S>6@?�����Q�>5�>sE�>�/k�oW���r��`]�>Y��?7��?�?��?����M>��=>���>頁?��?�O,>��ɾTى>9�8?��߾�FK�	��*K?O�@�D@b,>?'���dfۿ�#��N���G,��P��f'1<9Q�>UZ�=��A=�t�<�Yr�����q�6>�Ig>[k>9|>�2@>4UK>#��=(���^��P��:N���?�����������پ��x�?������_�����8z��Fnl���8��3l�K��=�T?T?1�s?�%? gZ�uf5>�x��T:=xU��Ħ=*��>�86?]�Q?��(?�>�=�9���c�H����x���/���>;9G>���>e��>	\�>��%���<>�#4>��y>��=��q=N�P��<��N>E�>��>i/�>FD<>�>Jδ��1����h��w��̽>�?7�����J��1��<������e�==b.?��>����>п�����1H?�����(���+���>
�0?�cW?�>"��S�T��<>(��-�j�c>, ���l�`�)��$Q>(k?#�h>��j>��0���7�`N�zƤ��~>�8?$ٵ�H�>��Mt��>K��ݾ�O>r��>嶰�2��er��e�}���h�6�=�
9?r�?9��������t������LL>~�U>��=�q�=�)L>�i���Ὦ�L���7=���=N�\>�M?�<>¢�=KA�>(����,I��P�>C}E>�U>)C?
(?�]�����Z�v�b/�p�w>���>��~>��>'�P�䍤="��>h�>&ܼTSŽ/Lʽ� ���L>z۵��CQ���6�A��=�&��8��=�}l=V���w=�n�H=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�'�>f���V���&����u� �!=�f�>�H?���f|L�8�>���
?��?<��^�����ȿ�dv�pv�>m�?Y�?�1n��c����?��!�>���?pY?��j>r�ھ�IY�ی>@A?�Q?x�>)��u%�;7?dݶ?�}�? ��=+�?�@f?���>�@"�����u/��r�|��$>�l����iN�����B���7q���'��c<'�=�i�>c��+����,��ͽ�ȝ�����i�> ؖ>S�]>G�>G��>�*�>�Ԟ>P��=����<�b���߾�K?��?��i�q� �r�Z>��?����>mfI?Y��=Š�����>��Z?���?.�K?a$�>�����󐿁3��&(��ޏ�����=�?)m�>����2�=_��X���K��>�+�>����k�ξ��Y�����f�>]q%?P��>�i>�� ?;�#?E�j>D#�>�^E�V8����E����>š�>�D?��~?C�?�ٹ��W3��	��硿��[�MUN>f y?fO?�ƕ>A������F�UI�S������?�wg?�,�f?f3�?�??��A?�f>���ؾ�,��>Cs?E����j��.P1��{�=�*9?�`�>_�)?�~ｊ�3�T�i�[T�����3�>~*B?��=?����h��a��(�
=xɽ�"=5�=��M�~7�>�܂>L��=D�>��|=ǅ3>H驾RH�<�>�w��Q6x=�>�;	-�^�=,?��G�ۃ���=k�r�xxD�?�>�GL>���@�^?o=�+�{����hx��FU�� �?Ƞ�?5k�?����h��$=?�?_?�"�>�I��)}޾C�ྌOw�	zx�w���>���>R�l���=�������8F���Ž�c���>�8�>�g�>^�?A�6>#�>/T��Fe)�����A	
���`��!��5�����������>������H��P��f�>볽���> �?U��>D��>�h�>�a�=P}o>
�O>M��>��>�"$>��>nM�=�F�/c��KR?�����'���辵����3B?�qd?z1�>�i�3������R�?���?Ls�?�<v>�~h��,+�an?h>�>=��Sq
?-T:=�0�Q:�<"V�����4��-�&��> E׽� :��M�Lnf�Aj
?�/?	��y�̾Z;׽�n���@�=�|t?��?���]���y�n{e���b�o���(>�q���.��cd��Q��om��6��f-� 6��;-?,N�?�ɾgi�Z����\���%���O>�j�>�gK>��>�*0>=A �cL���k��o8� %��[��>��z?6�>�lH?D�H?G9�?�#!?��6=�u?��<�b)?q�.>�?c�"?�H?��]?��?���>��1?�� >����������-?�F$?0�3?���>�?p�����ľe��gG���Z��i>��>���=H����;=�T?��E�8�K���5k>��7?�}�>>��>=���>��=U�<"��>��
?�K�>q����er��g��,�>Õ�?��[�=1�)>�_�=׀���ٺE�=�(ü���=]B��mM;���<���=��=��\ٹ��:��;���<�Y�>�#?٦�>�Z>�����,�	���A�<��<��������ɏ�~���o�p��l�<_g�?�"�?fgY>@LR=g�>�衾;�Ͼ����8��?�۠>`�M?zX?@q�?��D?O="?{E>�:��ɔ�����"%���	?R!,?��>��{�ʾr񨿬�3�Н?�[?J<a�����;)�]�¾��ԽX�>�[/��.~����)D��	�����1{��Λ�?���?�A���6�Uy�����~\���C?$!�>BY�> �>��)���g�x%�j2;>&��>MR?o#�>��O?%;{?W�[?:aT>c�8�s.���ҙ�Qh2���!>�@?��?��?Iy?np�>x�>8�)��ྥT�����a�ނ��DW=!Z>���>v'�>l�>���=� Ƚ(N��K�>�f�=,�b>��>�>�>S�w>�b�<��G?mY�>�澾UT��Q��y�����=�cu?Ґ?c,?�M=i�zE��%��H��>�?�?�?+�)?��S�ް�=�8ټn��h^m����>ȸ>Iޙ>
�=j�G=z�>��>XV�>C��bu�~78�lO�-�?
�E?��=NfƿZ�p���r��ޘ�L<:쓾�Af������]�.h�=^͘��8�:��y![��p���n��	���Y��ؔ|����>4q�=Z >���=&�<�ӼH�<�O9=��m<��=��n�V8_<�]G�G��ʿ��5����!<��?=���%ʾe�|?��F?R*? a;?��n>�D>ږ���L�>4���?��5>������l�E�*s��fs2侗 ؾb�.֗���>J`7�y��=b�!>c�=&��<&��=�|=�sD=���%�d=D�=F��=Ү�=�=4�>��=�T�?\���c��f9?����>ir�>3%3=Q��>'5����O?�b�;r;�Z�����=$s?���?+u�?�l�>h���o�>w�
�j���B@J>ŵS�� 9;䙨=m(P�Hͭ>Pq.�v93��H��4o󾄾�?Z�@D
L?󀥿�Ŀ�g�>�8>>��=Q�%�1�G�P�A&a�s�[�c!?�X;�c�̾�>D��=-�z�ƾ�r8=�R=>�Y=:)���Z���=�����L=Cs`=E݊>�XJ>�$�=�����=�
k=���=%|O>�-D��D���>�+�,=Ž=��Y>t�!>���>�?�`0?�Ud?i!�>��m�b�ξ�;��|p�>���=�[�>#�=$�B>S��>5�7?��D?��K?���>��=���>��>ʍ,���m��b� ا���<���?RȆ??��>�IU<ߗA�K��He>�"�Ľ5i?#M1?�i?U�>W����ڿ��2�Yy4�� 콋�ȼIM�=��>�&u�yB �/U:�Ӧǽ{��=�ѣ>���>��>J~\>6>t=>�w�>d'>.s=Lů=@I<��w<i��������Լ��b=fq�?񔼒�ü�>�;�҄�-v;�'B�)S�9��7=�=�|�>�4>��>W�=a��^�.>c��z�L��=����>B�7Od��*~���.�D 5��eB>�W>�烽��&�?.�Z>��>>wu�?�Ku?R!>_+��{վ����BJe�9�R����=K�>|�=�P];�@P`��M��Ҿq��>}�>��>ڻl>,��!?���w=W�l_5���>�|��3���'�d:q��?��P����i��պ?�D?�E��z��=2 ~?o�I?�?T��>!��Ёؾ�-0>�L����=���q�1o����?*'?ە�>��a�D�bD�����v*W>k3ɾ'N^�"ȋ��$���r�}%¾-�>4vž�䔾t1�gs������ߢW�w]��n�?�~?�F�?�E��n��u�T�c��s8�=-?�X�?��>l�'?�T�>��A>E;���sE��H�<vz�?L��?�U�?ЎB>���=xD��|'�>��
?0f�?���?��t?��>�$��>X��;M�&>l���Q�=�h>Ί�=���=��?h5
?��	?@�Z�����p��`�v��<L��=T?�>��>BIr>���=�-M=��=�X>dQ�><��>ac>o�>1҈>���s����&?K��=��>2?��>'�_="���5�<��S��}A�8�-���F޽�R�<�����zG=�aʼ���>�\ǿ7��?�S>��FY?���$��T>�4V>�i޽�	�>�`F>��|>��>���>vM>�7�>��&>۟�/T>�C�8�!���=�~\�\l�n��=�پ�7P�ho��g��=C��1-پ���x�w�V����g0��6J=U�?r� ^e��-<�z�.�]j?���>��5?YT��E��l��<p�>ɋ8>�c������c��өѾ
��?���?-%u>�,�>��6?F�?���;q�׾=N���i����<��?Ca�V=��XS����&��b�ܙ3?�q??I?6�D>�_r>-��?��
�B�����>�$7�� ��:�i�G>ͯ��[���Y����i$p��K>VB?�E�?�:?K����<����b>'r?�*�?;A[?;�W?��?�����?}={>��?)�<?Jt?�v?��%?=ɵ=Ҕ�>W�>_̣:ᝏ��g�.�<3��M�ݢ=p�ʽ�6�=�:�=b<=p">��o|ý�~Z�3��=\�+��qX<U� >��=��>��[?k-�>�f�>�6?H�-�P+5�K����W'?9�	=�V���ˏ�4&��PS��=4~e?�.�?�[?gk>�U>��68���>�R�>t=>��[>�ݯ>I����-��ؓ=��
>�>��=!]1�˃����F����=%�>�<?>q���P=9�w�:Ѭ�᡻�ED�|ϾK��gkT�ޔS����]x�>4J^?��@?<5�=~Ⱦ}�?=�e��2?~Fa?��?bb�?��1=����2� i[��6=߻�>��]=i��oǦ�a���iD��E�<9�S>W��4٠�_�c>�^�b޾�:n�~+J�����;?=����V=���v�Ծvs~��a�='�>�F���!��&���Ϫ�[yJ?�Ak=8̦�cX�Z)���Q>��>��>t�=���u��@���z�=Ψ�>�9>�ڨ0G����9��>Z]?�Na?��k?���nU��7�6V
�I�������
�>��>-��>y?>��	=�h��VN�-�h���n����>��>f-�N�W��CᾀO侂��Gd�>�?6�>TD?�rG?��?:i]?��=?	�?;��>׼1��m�*?��?9��=�l\�Ir����*�	-C�M�>��5?ĝ��~�>m�
?߸?&?FYN?��?r�E>z����N���>�V>z)^��ӱ��ߢ>��??�'\>W_Q?���?��>v(�np����T��7*>�j>�1@?�_)?�?װ�>s��>&Ɨ��4�>�t ?�,?���?\g?�{>���>��D>}k?OC��x�?l�	?`<?�^0?�e9?-�S?V�>#�;M�뽯H��i4G��4�н��1�:�5�*�ֽ�;�<KV'>g*s�"�ټ��ڻV-�o�μMh�ë=�_�>j�s>+
��f�0>F�ľ�O����@>쇣�%P��$ڊ�9�:�c޷=5��>��?#��>�X#����=/��>I�>6���6(?��?�?k�!;��b���ھ��K���>"	B?T��=��l�����q�u��g=��m?s�^?��W�l&��L�_?>g?���Y�2���K#���6���.?qN?�T�\�>��w?�=n?��>��F���1����h��c���M�=ӡ>�	���V�9wq>�%)?���>��>��1=Tվ=�u������G$?���?Xȵ?���?�� >�+Y�����Ҿ!�����a?9�>����a1?��R=e־�ܦ��þ;������ƾ�d��3�о�KĽD������n��=?|�H?��\?;Q�?����W� �q��ـ��_��ܾr�۩L��%�P/��ʐ��;�Œپ����d<Ɂ���j7�Y��?�'?�1%��1�>���iM����˾z�/>�Μ��+��ڛ=�@W�1*=Ȣ�<y�%qW��幾=H$?��>�
�>��9?�7U���>�Y�<�X�G�����|S>�
�>$ѣ>A1�>7�	�� <�1��Ӿ�������>"�?�?j~Z?��9�ɞ(��[��Ω:���=)e��A���W�=N��>���Vze��'c��q'�Z%s��+K�֮��r��wD�>0}*?1�=�P�>V3�?�x?�uP�9��� ����b+����$>�b?��?�tB>��"�t�ɺ�>B�l?d��>�>�����Z!�0�{�!�ʽ54�>�׭>ǥ�>$�o>ǧ,��"\��k�������9�Q=�=ݢh?������`��߅>8R?��:�zG<F��>�mv�B�!������'�A�>M�? ʪ=?�;>c~ž� �2�{��I��	G)?�:?/���ڀ*�:~>',"?�j�>@6�>q(�?[|�>3þk�V��?��^?�GJ?�SA?�Q�>A)=�����Ƚ�&�,=㊇>2�Z>��l=I��=M����\�����<F=~�=�*μ�y��Ú<>,����K<o��<��3>��տ�>�nּ�����y�ھ�����JS���w��6�����s����r�mԽ��z��(~��`��(�����?�>�?��$��(���������z��-!>`��ŝu������𽿪��zYӾuU��s
"��*T������g� q8?x/z��῍r��5p����?iΪ>�ȃ?�03��ؾ��R�j����^�:5��7� 
��'�߿`�*%h?f�?�����)����>��2=q��>@hY>��u��/W��O��34?��:?4s$?1���<�ɿ�Yɿ>lT�?��@�|A?.�(����V=[��>�	?��?>:W1��G�����$R�><�?���?�M=T�W���	��e?vS<G�F���ݻ5�=G?�=�F=���6�J>�V�>��HWA�n@ܽA�4>hم>�i"�٨��z^���<Ą]>�սwE��5Մ?*{\��f���/��T��U>��T?�*�>b:�=��,?X7H�`}Ͽ�\��*a?�0�?���?&�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=S6�Z���~���&V����=_��>a�>ł,�����O��I��Y��=����f¿L/�2����A��j&��
j�e{q���L��ͽ_W��Wx��f��cc�=��=�v>���>6N>�R2>S�P?$�?m��>��I>��̒���� ���ټ�g2�x�"��j���d�z8ȾGE��m������� ����־��;�H��=�Q�P6�����fd�*�H��+?6�>z�Ⱦ��L��!�<�ɾ�^����ż1���>5Ͼ8�3���m��z�?6�??w뇿�Y�=���S�k���;G^?x���I��+�=��
��
�<���>��=�-�3�2�Z#Q�;?��,?��A�m��>���v�v;`�0?x�"?=U>�{�>��4?�@���޽�<i>�M�>���>���>���=��̾
G���?R�w?�K:���ľt��>�������ΝB�B��=��;"�>�c�>W#���"ܾ�S=�u�����<�(W?/��>��)�m�t`������R==��x?�?�1�> {k?��B?���<�g���S���!xw=k�W?)i?Ҷ>􆁽оK|��z�5?��e?��N>B_h���龽�.��T��%?��n?d_?�����w}�������Qn6?M�|? gC�윿���4վ�6�=���>1	?ʺJ����>��<?���#ә���̿�H��ؙ?��@|��?�w�=X����zK>��)?��>��y����QF�o���� �=f2�>��;����2?*��s�h?���?�?v
s����*o>h����?7�?־2*=�X�׿u��>�������jވ����ݾ-V�9�ɾ�0�.ɾ�:�<]T�>�@�:a�W�?|O��2�3ֿ.��� 0����W�!/�>}��>\$���� l�ԇv�� 8��ch�B$��혣>���>���iԾM�p�?���J�7z�>�cؽ�\�>����> G��&��x]���*>���>>������	��Z�?+@��F�ܿ����(��h�4?�ۏ?���?��%?�s>G�z�_�$�u�O!0?�gz?�:�?[�����+����=�Ep?���Irl�>�4���M�?��=��*?e:�>��;���<�E>|�?���=w�H�:_ĿB"��/�׾�(�?���?V �ix?~E�?�n$?'�(�� �Q���Zr)��<����C?��S>g�ݾ9�2�?
B�A���-O ?�UV?��M��#1�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�"�>T�?���=`d�>9�=$簾�T.��D#>��=]_?��?\�M?�A�>L�=�9��$/��TF��HR��.���C���>��a?uL?~Cb>�︽�1��� ���ͽ�p1�Pb�FG@�"_-���߽5>D>>�>P�D��
Ӿ�O3?��̦�S����E�1�?�FC>�.(?p���k���X�䫀?2�f>?k6�����G���C�c�k�?1�?���>�ޱ�1H>��C>"�==�޼�V=Tb��ʓ��<�=d�s?�2�ӯ��ԃ�\ۂ>�þ?uL@@��?��j�D�
?�r������}�r��}�D���=<�:?0����q>3�>:�=�'w�-��6u��=�>�Ư?���?��>�i?�k�|<�<�5=*��>��d?L?*��#���I>�2	?Z��᏿����?d?&�
@@/@��_?�᣿��ܿ\��ھ'վb �=h\<�Km;>:����>.�=��H=�0��I=A~>dY>�#>Z�>�;1>��>5�����ԛ�I�����A��,�cL���Ž0�澇7<����f8�@p��  �=aKl�<ǣ�^n����Z�pv;���=]�U?��Q?��o?A��>M7v��>c%��cH�<�$�4��=0Ӆ>2?!�K?��)?P��=E����d�憁�xk��������>��G>�5�>=��>�Ů>��:"dG>�=>�*�>� >Ć=��L�=�UP>F[�>v7�>���>@{l>�P>�L��J
��k�,�T0���/����?~#վw�5�@	����*�����{{;�A?-�>	C���ٿ�o����U?h���c�2�O$�OM^>NG?�vZ?�j>5��v��=��{=H�˾������=�TҽR�_�E�5��B >� ?�f>@u>U�3��d8���P�Q{���g|>x26?b鶾�G9��u�^�H�}cݾ�DM>�¾>HED��k�W�����ui�R�{=:x:?��?�;���᰾̭u��B��KQR>�9\>Y=Ul�=yVM>YXc���ƽ(H��i.=]��=��^>V#?�*>��='�>$���"�M����>�)C>�D+>�@?�[%?�������G,��v>��>�q�>�<>k�I���=���>z{a>6@�D����x��?��UV>�z���]�cq�au=�ؘ��3�=h��=�; �Ug=���'=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�k�>9z�\�������u���#=��>:H?;Y����O��>� w
?�?�a�M�����ȿ�~v����>�?@��?��m��?���@�Uy�>e��?�gY?ti>e۾snZ�ޑ�>z�@?�R?��>�9�6�'���?H�?���?U��>���?��?��?O��=��%�v�ʿ�@��C�?����([����~>����!��&@��}��ZuI��~P�h~�>5m�<�X?��^�lN$���)>d��<Td�������.�>�s�>TV�>�BE>W#?La?s�^>�c����=��&��YI���K?���?0��1/n��L�<O��=9�^�� ?FL4?��[���Ͼ6ը>`�\?���?,�Z?;Q�>���)>���迿^��p��<��K>76�>�=�>���/YK>�Ծ�ND�*m�>Η>�C��8ھ�,������G�>�a!?_��>���=�� ?�#?�j>��>q0E�_G��4AF�=Z�>�q�>��?J�}?h:?.�����3�����ʡ���[� ^L>Gzy?.?/��>ċ��>����X)��DD����em�?�g?�F�;?E3�?{4??�,A?[�f>���ݟ׾Y���'��>��!?��A��K&���&?�P?!��>�9����ս.�ռ���jz����?�(\?�?&?6���)a�j�¾�7�<
�"�\V�d��;L�D���>i�>9�����=�>�۰=�Mm�8H6��f<\e�=�>���=417��|��� 2?�)=u����;J<"�����j�]�{>mAY>޽�VC?{�-� _�������������n�?R��?�{�?�+���p�4,9?�A�?���>�?0򐾂^���$� 5~�&}������}ܼ@�>Ws�=BFᾼ���:��x���� ���ڽ��?�а>H5�>�S?��<>P��>����a�+�֠'�����k�l'0�wV?���/�Ά"�hw���������ʾ�܆�HǼ>;@Žs&r>��/?cv`>E��>��
??~���O>߱�>�P^>���>H��>E<>&=�����-��KR?�����'�y������f3B?�qd?M1�>Yi�6��������?���?Qs�?0=v>h��,+��n?�>�>D��Rq
?pT:=�9�i:�<V��s��3��[�3��>�D׽� :��M�2nf�rj
?�/?�����̾�;׽�N~��)�=�bc?��J?EQ#���q�r����ڎ��2��S�[�Ͼ�p^�t[�f�!���%��N5���ZY���>�4?U�?͉5�s���0���Iq��q��c >�?�N�>l5�=%�?b��m��87�ǟ�ܸz��́>�}?�i�>sXL?ئ_?�Zt?xe�?���>=?����`�>X>��>��)?:�6?F?��B?��;?��I?�s�>ω[�RD�@V��s�'?5��>�?�r
?��?����V)��3��K�=���,>y�=C�>PHZ�~���x�>o=�=wM?Ȧ�{�8�����	�j>ۅ7?,��>���>V��� ��$`�<��>�
?VR�>�����jr�:S��]�>��?��G=�)>A��=�cߺ=L�=������=����q:�|� <-�=��=tz��Q��-��:��{;z��<�u�>y�?���>C�>�?���� �T���h�=�Y>� S>m>�Dپ ~��j$����g�7ay>�w�?�z�?Y�f=a�=y��=|���R�����#���h�<(�?+I#?sVT?3��?��=?�k#??�>O+��M��X^��3����?v!,?��>�����ʾ��Չ3�ם?e[?�<a����;)���¾��Խʱ>�[/�k/~����>D�����_��6��?쿝?dA�R�6��x�ٿ���[��x�C?"�>Y�>��>V�)�z�g�o%��1;>���>jR?>$�>B�O?#8{?��[?�{T>ܕ8�b-���ҙ�'o1�h�!>q@?��?U�?�y?�l�>8�>��)����^�������Nւ�W=h�Y>���>l*�>��>���=��ǽ+^��V�>����=ɔb>Е�>s��>\��>��w>�9�<*Z?i�?�����5�\GH�f��	mz�^nD?��?��?��7<���4�z�԰���>���?�?��?���A�	>��׽�`��T�O=���>��>k8�> >��=6&�=T�>R��>�`���'���#�am�x�?�6?@�w>�ƿ�q��.q��2QZ<�����d�5����Z���=}���o���i����Z�&Y���z�����X�����{�.��>5*�=vp�=q��=�c�<�x˼;�<�'K=A�<�/=��p���e<� :��dԻ�䉽� ��X<��I=r=����Ⱦp�}?o?I?�	+?aA?!�z>[>i2@�zM�>�w���d?��Q>!�V�󂽾">����C�����پb�۾L�b���>� ^���>�,2>��=���<7�=1�g=���=�:��=���=A7�=��=��=z>�a>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?~�>>�2������yb��-?���?�T�?>�?Ati��d�>M���㎽�q�=F����=2>o��=w�2�U��>��J>���K��H����4�?��@��??�ዿТϿ7a/>��7>�&>w�R�E�1� �\���b��xZ�՚!?�H;��J̾6�>��=Q+߾�ƾN�.=ք6>T_b=Th�pV\���=��z���;=-�k=0Չ>s�C>�x�=.���=¥I=���=��O>�v����7��(,�Q�3=���=�b>&>!��>�?uZ0?G)d?_�>b�m��Ͼ�<���g�>���=�-�><��=qOB>T��>�7?1�D?2�K?�k�>�v�="�>��> �,�$�m�9.�ٱ��$]�<���?�ӆ?�M�>�U<I�A�T��VA>���ý��?�K1?w?k��>�^� ӿ�w(�y�Z���׾;[w�8w=e�鼵�=�%Xɽ��<{DM=�zM>�h?��>i�j>bM�>��n=��=���>��>^ݖ=��>�%D;���=4�ü�<~<K�o���ӽ`���=��=���~�/��S����=�Gw<���+>���>蔶=��;>��>׺	���>М�p�U.��|��ŕt�J��>z��b�O�`�+��]>��>���=)�����>�D>�~�=��?`��?@�>�-�A*�����4����@�t^�=bC�>"�<��L�艇��zc�2�˾Z��>g�>�>��l>�	,�#&?�8\w=��W5�0��>和�_��@@�@q��?��b����i��L�J�D?�C��	��=I~?��I?��?���>�H���ؾ_W0>E��6=g��4q�Ȏ����?�'?���>~��D��J̾�I���շ>�3I���O��ŕ�&�0�^*��﷾��>Dݪ��о�3�b^��������B��r����>A�O?���?B(b�j���xO�.��qB��Gf?�g?9�>�<?�?�Ġ�*��Ϣ�����=��n?s��?�*�?>t�=�X�)J?RI?sF�?&��?��{?̦����>|�N=�b>�5޽od>6�F>��/>;�/>(#�>+�?W>�> �����$����]�Wv��:=g�0=�Y�>`l8>N&>��=���<��=�a(>ߵ�>�L�>4�L>���>��>瞄�L��	?wq����>g#;? v�>W��<%���l�Ɓ��~�M�3桾-�񽋒�x��'D%�O46>ӮU=ѻ�>uͿ��?��>z�$�~(?x4����	���)>�Р>�H���>
��>(�>��g>��>�y�=��><RR>EӾ{1>�V��� �<uB���R�cwԾ!ur>N�$�K�h��(�G��9�����+j�P>���=�6g�<΋�?�a���m��++������?�Ψ>Xi7?��������D>���>'��>>�������e���r�྽��?�]�?�;c>�>P�W?�?��1�N3��uZ��u�.(A�?e���`�T፿ߜ���
��	��F�_?y�x?*xA?D.�<*:z>*��?n�%�3ԏ�w(�>�/�w&;��@<=�+�>P)��O�`���ӾB�þ:6�JF>��o?%�?'Y?�TV�c��=	K��{1?��#?i��> BJ?!\=?X�>1��>�V�>��U?��e>�N?�'?�/?x�g=��="'�>�{=h�v��OU�\y�Ԍ��7��g�9�^�=?W�=��=.gW�*ñ�^½Y4B����;����-���V�=��L��`}=>�>��^?.�>.Xt>�+8?����&9�jE��Ğ8?�H�=��x����+��<1�:E>��r?d=�?yV?1pS>FB��GC��#>�]�>Q6>�JM>�ݼ>�k��^/O�H��<ە&>��.>XS�=hܐ�r��Ob����k�=�b.>���>C1|>���r�'>�|���0z���d>��Q��̺���S���G���1�|�v�?Y�>��K?J�?U��=y_�J/��`If�0)? ^<?�NM?��?"�=�۾[�9��J��>���>�X�< �������#����:�m�:O�s>�1��4٠�_�c>�^�b޾�:n�~+J�����;?=����V=���v�Ծvs~��a�='�>�F���!��&���Ϫ�[yJ?�Ak=8̦�cX�Z)���Q>��>��>t�=���u��@���z�=Ψ�>�9>�ڨ0G����9��>Z]?�Na?��k?���nU��7�6V
�I�������
�>��>-��>y?>��	=�h��VN�-�h���n����>��>f-�N�W��CᾀO侂��Gd�>�?6�>TD?�rG?��?:i]?��=?	�?;��>׼1��m�*?��?9��=�l\�Ir����*�	-C�M�>��5?ĝ��~�>m�
?߸?&?FYN?��?r�E>z����N���>�V>z)^��ӱ��ߢ>��??�'\>W_Q?���?��>v(�np����T��7*>�j>�1@?�_)?�?װ�>s��>&Ɨ��4�>�t ?�,?���?\g?�{>���>��D>}k?OC��x�?l�	?`<?�^0?�e9?-�S?V�>#�;M�뽯H��i4G��4�н��1�:�5�*�ֽ�;�<KV'>g*s�"�ټ��ڻV-�o�μMh�ë=�_�>j�s>+
��f�0>F�ľ�O����@>쇣�%P��$ڊ�9�:�c޷=5��>��?#��>�X#����=/��>I�>6���6(?��?�?k�!;��b���ھ��K���>"	B?T��=��l�����q�u��g=��m?s�^?��W�l&��L�_?>g?���Y�2���K#���6���.?qN?�T�\�>��w?�=n?��>��F���1����h��c���M�=ӡ>�	���V�9wq>�%)?���>��>��1=Tվ=�u������G$?���?Xȵ?���?�� >�+Y�����Ҿ!�����a?9�>����a1?��R=e־�ܦ��þ;������ƾ�d��3�о�KĽD������n��=?|�H?��\?;Q�?����W� �q��ـ��_��ܾr�۩L��%�P/��ʐ��;�Œپ����d<Ɂ���j7�Y��?�'?�1%��1�>���iM����˾z�/>�Μ��+��ڛ=�@W�1*=Ȣ�<y�%qW��幾=H$?��>�
�>��9?�7U���>�Y�<�X�G�����|S>�
�>$ѣ>A1�>7�	�� <�1��Ӿ�������>"�?�?j~Z?��9�ɞ(��[��Ω:���=)e��A���W�=N��>���Vze��'c��q'�Z%s��+K�֮��r��wD�>0}*?1�=�P�>V3�?�x?�uP�9��� ����b+����$>�b?��?�tB>��"�t�ɺ�>B�l?d��>�>�����Z!�0�{�!�ʽ54�>�׭>ǥ�>$�o>ǧ,��"\��k�������9�Q=�=ݢh?������`��߅>8R?��:�zG<F��>�mv�B�!������'�A�>M�? ʪ=?�;>c~ž� �2�{��I��	G)?�:?/���ڀ*�:~>',"?�j�>@6�>q(�?[|�>3þk�V��?��^?�GJ?�SA?�Q�>A)=�����Ƚ�&�,=㊇>2�Z>��l=I��=M����\�����<F=~�=�*μ�y��Ú<>,����K<o��<��3>��տ�>�nּ�����y�ھ�����JS���w��6�����s����r�mԽ��z��(~��`��(�����?�>�?��$��(���������z��-!>`��ŝu������𽿪��zYӾuU��s
"��*T������g� q8?x/z��῍r��5p����?iΪ>�ȃ?�03��ؾ��R�j����^�:5��7� 
��'�߿`�*%h?f�?�����)����>��2=q��>@hY>��u��/W��O��34?��:?4s$?1���<�ɿ�Yɿ>lT�?��@�|A?.�(����V=[��>�	?��?>:W1��G�����$R�><�?���?�M=T�W���	��e?vS<G�F���ݻ5�=G?�=�F=���6�J>�V�>��HWA�n@ܽA�4>hم>�i"�٨��z^���<Ą]>�սwE��5Մ?*{\��f���/��T��U>��T?�*�>b:�=��,?X7H�`}Ͽ�\��*a?�0�?���?&�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=S6�Z���~���&V����=_��>a�>ł,�����O��I��Y��=����f¿L/�2����A��j&��
j�e{q���L��ͽ_W��Wx��f��cc�=��=�v>���>6N>�R2>S�P?$�?m��>��I>��̒���� ���ټ�g2�x�"��j���d�z8ȾGE��m������� ����־��;�H��=�Q�P6�����fd�*�H��+?6�>z�Ⱦ��L��!�<�ɾ�^����ż1���>5Ͼ8�3���m��z�?6�??w뇿�Y�=���S�k���;G^?x���I��+�=��
��
�<���>��=�-�3�2�Z#Q�;?��,?��A�m��>���v�v;`�0?x�"?=U>�{�>��4?�@���޽�<i>�M�>���>���>���=��̾
G���?R�w?�K:���ľt��>�������ΝB�B��=��;"�>�c�>W#���"ܾ�S=�u�����<�(W?/��>��)�m�t`������R==��x?�?�1�> {k?��B?���<�g���S���!xw=k�W?)i?Ҷ>􆁽оK|��z�5?��e?��N>B_h���龽�.��T��%?��n?d_?�����w}�������Qn6?M�|? gC�윿���4վ�6�=���>1	?ʺJ����>��<?���#ә���̿�H��ؙ?��@|��?�w�=X����zK>��)?��>��y����QF�o���� �=f2�>��;����2?*��s�h?���?�?v
s����*o>h����?7�?־2*=�X�׿u��>�������jވ����ݾ-V�9�ɾ�0�.ɾ�:�<]T�>�@�:a�W�?|O��2�3ֿ.��� 0����W�!/�>}��>\$���� l�ԇv�� 8��ch�B$��혣>���>���iԾM�p�?���J�7z�>�cؽ�\�>����> G��&��x]���*>���>>������	��Z�?+@��F�ܿ����(��h�4?�ۏ?���?��%?�s>G�z�_�$�u�O!0?�gz?�:�?[�����+����=�Ep?���Irl�>�4���M�?��=��*?e:�>��;���<�E>|�?���=w�H�:_ĿB"��/�׾�(�?���?V �ix?~E�?�n$?'�(�� �Q���Zr)��<����C?��S>g�ݾ9�2�?
B�A���-O ?�UV?��M��#1�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�"�>T�?���=`d�>9�=$簾�T.��D#>��=]_?��?\�M?�A�>L�=�9��$/��TF��HR��.���C���>��a?uL?~Cb>�︽�1��� ���ͽ�p1�Pb�FG@�"_-���߽5>D>>�>P�D��
Ӿ�O3?��̦�S����E�1�?�FC>�.(?p���k���X�䫀?2�f>?k6�����G���C�c�k�?1�?���>�ޱ�1H>��C>"�==�޼�V=Tb��ʓ��<�=d�s?�2�ӯ��ԃ�\ۂ>�þ?uL@@��?��j�D�
?�r������}�r��}�D���=<�:?0����q>3�>:�=�'w�-��6u��=�>�Ư?���?��>�i?�k�|<�<�5=*��>��d?L?*��#���I>�2	?Z��᏿����?d?&�
@@/@��_?�᣿��ܿ\��ھ'վb �=h\<�Km;>:����>.�=��H=�0��I=A~>dY>�#>Z�>�;1>��>5�����ԛ�I�����A��,�cL���Ž0�澇7<����f8�@p��  �=aKl�<ǣ�^n����Z�pv;���=]�U?��Q?��o?A��>M7v��>c%��cH�<�$�4��=0Ӆ>2?!�K?��)?P��=E����d�憁�xk��������>��G>�5�>=��>�Ů>��:"dG>�=>�*�>� >Ć=��L�=�UP>F[�>v7�>���>@{l>�P>�L��J
��k�,�T0���/����?~#վw�5�@	����*�����{{;�A?-�>	C���ٿ�o����U?h���c�2�O$�OM^>NG?�vZ?�j>5��v��=��{=H�˾������=�TҽR�_�E�5��B >� ?�f>@u>U�3��d8���P�Q{���g|>x26?b鶾�G9��u�^�H�}cݾ�DM>�¾>HED��k�W�����ui�R�{=:x:?��?�;���᰾̭u��B��KQR>�9\>Y=Ul�=yVM>YXc���ƽ(H��i.=]��=��^>V#?�*>��='�>$���"�M����>�)C>�D+>�@?�[%?�������G,��v>��>�q�>�<>k�I���=���>z{a>6@�D����x��?��UV>�z���]�cq�au=�ؘ��3�=h��=�; �Ug=���'=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�k�>9z�\�������u���#=��>:H?;Y����O��>� w
?�?�a�M�����ȿ�~v����>�?@��?��m��?���@�Uy�>e��?�gY?ti>e۾snZ�ޑ�>z�@?�R?��>�9�6�'���?H�?���?U��>���?��?��?O��=��%�v�ʿ�@��C�?����([����~>����!��&@��}��ZuI��~P�h~�>5m�<�X?��^�lN$���)>d��<Td�������.�>�s�>TV�>�BE>W#?La?s�^>�c����=��&��YI���K?���?0��1/n��L�<O��=9�^�� ?FL4?��[���Ͼ6ը>`�\?���?,�Z?;Q�>���)>���迿^��p��<��K>76�>�=�>���/YK>�Ծ�ND�*m�>Η>�C��8ھ�,������G�>�a!?_��>���=�� ?�#?�j>��>q0E�_G��4AF�=Z�>�q�>��?J�}?h:?.�����3�����ʡ���[� ^L>Gzy?.?/��>ċ��>����X)��DD����em�?�g?�F�;?E3�?{4??�,A?[�f>���ݟ׾Y���'��>��!?��A��K&���&?�P?!��>�9����ս.�ռ���jz����?�(\?�?&?6���)a�j�¾�7�<
�"�\V�d��;L�D���>i�>9�����=�>�۰=�Mm�8H6��f<\e�=�>���=417��|��� 2?�)=u����;J<"�����j�]�{>mAY>޽�VC?{�-� _�������������n�?R��?�{�?�+���p�4,9?�A�?���>�?0򐾂^���$� 5~�&}������}ܼ@�>Ws�=BFᾼ���:��x���� ���ڽ��?�а>H5�>�S?��<>P��>����a�+�֠'�����k�l'0�wV?���/�Ά"�hw���������ʾ�܆�HǼ>;@Žs&r>��/?cv`>E��>��
??~���O>߱�>�P^>���>H��>E<>&=�����-��KR?�����'�y������f3B?�qd?M1�>Yi�6��������?���?Qs�?0=v>h��,+��n?�>�>D��Rq
?pT:=�9�i:�<V��s��3��[�3��>�D׽� :��M�2nf�rj
?�/?�����̾�;׽�N~��)�=�bc?��J?EQ#���q�r����ڎ��2��S�[�Ͼ�p^�t[�f�!���%��N5���ZY���>�4?U�?͉5�s���0���Iq��q��c >�?�N�>l5�=%�?b��m��87�ǟ�ܸz��́>�}?�i�>sXL?ئ_?�Zt?xe�?���>=?����`�>X>��>��)?:�6?F?��B?��;?��I?�s�>ω[�RD�@V��s�'?5��>�?�r
?��?����V)��3��K�=���,>y�=C�>PHZ�~���x�>o=�=wM?Ȧ�{�8�����	�j>ۅ7?,��>���>V��� ��$`�<��>�
?VR�>�����jr�:S��]�>��?��G=�)>A��=�cߺ=L�=������=����q:�|� <-�=��=tz��Q��-��:��{;z��<�u�>y�?���>C�>�?���� �T���h�=�Y>� S>m>�Dپ ~��j$����g�7ay>�w�?�z�?Y�f=a�=y��=|���R�����#���h�<(�?+I#?sVT?3��?��=?�k#??�>O+��M��X^��3����?v!,?��>�����ʾ��Չ3�ם?e[?�<a����;)���¾��Խʱ>�[/�k/~����>D�����_��6��?쿝?dA�R�6��x�ٿ���[��x�C?"�>Y�>��>V�)�z�g�o%��1;>���>jR?>$�>B�O?#8{?��[?�{T>ܕ8�b-���ҙ�'o1�h�!>q@?��?U�?�y?�l�>8�>��)����^�������Nւ�W=h�Y>���>l*�>��>���=��ǽ+^��V�>����=ɔb>Е�>s��>\��>��w>�9�<*Z?i�?�����5�\GH�f��	mz�^nD?��?��?��7<���4�z�԰���>���?�?��?���A�	>��׽�`��T�O=���>��>k8�> >��=6&�=T�>R��>�`���'���#�am�x�?�6?@�w>�ƿ�q��.q��2QZ<�����d�5����Z���=}���o���i����Z�&Y���z�����X�����{�.��>5*�=vp�=q��=�c�<�x˼;�<�'K=A�<�/=��p���e<� :��dԻ�䉽� ��X<��I=r=����Ⱦp�}?o?I?�	+?aA?!�z>[>i2@�zM�>�w���d?��Q>!�V�󂽾">����C�����پb�۾L�b���>� ^���>�,2>��=���<7�=1�g=���=�:��=���=A7�=��=��=z>�a>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?~�>>�2������yb��-?���?�T�?>�?Ati��d�>M���㎽�q�=F����=2>o��=w�2�U��>��J>���K��H����4�?��@��??�ዿТϿ7a/>��7>�&>w�R�E�1� �\���b��xZ�՚!?�H;��J̾6�>��=Q+߾�ƾN�.=ք6>T_b=Th�pV\���=��z���;=-�k=0Չ>s�C>�x�=.���=¥I=���=��O>�v����7��(,�Q�3=���=�b>&>!��>�?uZ0?G)d?_�>b�m��Ͼ�<���g�>���=�-�><��=qOB>T��>�7?1�D?2�K?�k�>�v�="�>��> �,�$�m�9.�ٱ��$]�<���?�ӆ?�M�>�U<I�A�T��VA>���ý��?�K1?w?k��>�^� ӿ�w(�y�Z���׾;[w�8w=e�鼵�=�%Xɽ��<{DM=�zM>�h?��>i�j>bM�>��n=��=���>��>^ݖ=��>�%D;���=4�ü�<~<K�o���ӽ`���=��=���~�/��S����=�Gw<���+>���>蔶=��;>��>׺	���>М�p�U.��|��ŕt�J��>z��b�O�`�+��]>��>���=)�����>�D>�~�=��?`��?@�>�-�A*�����4����@�t^�=bC�>"�<��L�艇��zc�2�˾Z��>g�>�>��l>�	,�#&?�8\w=��W5�0��>和�_��@@�@q��?��b����i��L�J�D?�C��	��=I~?��I?��?���>�H���ؾ_W0>E��6=g��4q�Ȏ����?�'?���>~��D��J̾�I���շ>�3I���O��ŕ�&�0�^*��﷾��>Dݪ��о�3�b^��������B��r����>A�O?���?B(b�j���xO�.��qB��Gf?�g?9�>�<?�?�Ġ�*��Ϣ�����=��n?s��?�*�?>t�=�X�)J?RI?sF�?&��?��{?̦����>|�N=�b>�5޽od>6�F>��/>;�/>(#�>+�?W>�> �����$����]�Wv��:=g�0=�Y�>`l8>N&>��=���<��=�a(>ߵ�>�L�>4�L>���>��>瞄�L��	?wq����>g#;? v�>W��<%���l�Ɓ��~�M�3桾-�񽋒�x��'D%�O46>ӮU=ѻ�>uͿ��?��>z�$�~(?x4����	���)>�Р>�H���>
��>(�>��g>��>�y�=��><RR>EӾ{1>�V��� �<uB���R�cwԾ!ur>N�$�K�h��(�G��9�����+j�P>���=�6g�<΋�?�a���m��++������?�Ψ>Xi7?��������D>���>'��>>�������e���r�྽��?�]�?�;c>�>P�W?�?��1�N3��uZ��u�.(A�?e���`�T፿ߜ���
��	��F�_?y�x?*xA?D.�<*:z>*��?n�%�3ԏ�w(�>�/�w&;��@<=�+�>P)��O�`���ӾB�þ:6�JF>��o?%�?'Y?�TV�c��=	K��{1?��#?i��> BJ?!\=?X�>1��>�V�>��U?��e>�N?�'?�/?x�g=��="'�>�{=h�v��OU�\y�Ԍ��7��g�9�^�=?W�=��=.gW�*ñ�^½Y4B����;����-���V�=��L��`}=>�>��^?.�>.Xt>�+8?����&9�jE��Ğ8?�H�=��x����+��<1�:E>��r?d=�?yV?1pS>FB��GC��#>�]�>Q6>�JM>�ݼ>�k��^/O�H��<ە&>��.>XS�=hܐ�r��Ob����k�=�b.>���>C1|>���r�'>�|���0z���d>��Q��̺���S���G���1�|�v�?Y�>��K?J�?U��=y_�J/��`If�0)? ^<?�NM?��?"�=�۾[�9��J��>���>�X�< �������#����:�m�:O�s>�1���7��� b>M���gԾFW��B�����|���n#��A=���쒬�ߓw����=h��=����M.#��k�����/�H?�o�=_*��Z��ٛ��Q>%X�>$^�>}�ý�.＃�;��R���1|=PԹ>�ݼ=���b��D�����߄>�A?�g^?�B~?$U��n�Y�d)D�'�������~sμZm?z�>GE�>�!>˹�=rǲ�X�)h� B���>���>8��rI�zО�M��� ��ڗ>�^ ?�C�>��?B�W?��?�%d?n"?�?�ς>�P��hī��A&?.��?R�=��Խ6�T�K 9�MF�i��>Y�)?
�B�繗>=�?��?��&?��Q?Ե?�>� ��C@�ٔ�>]Y�>��W��b���_>��J?�>u=Y?�ԃ?��=>W�5��颾�թ��V�=�>��2?�5#?H�?���>�t�>��d�=���>��b?�-�?��o?I�=�?42>���>�K�=!��>�b�>�?l6O?��s?��J?ˍ�>|܎<_������Z�r��,R�i%};T�G<��y=k�b_t���wc�<�M�;�~����}�N���D��Ꮌ*��;fg�>d�s>������0>�ž>���A>e̟����#�����:��/�=._�>+�?h��>~)#�ϒ=k�>��>���;(?/�?�9?�+;µb��ھgL����>O�A?)��=.�l�P|��F�u�_�f=��m?��^?�W�G��r-r?Y�2?���B^�M	����ƽ!��?S�=?��>%��>��?�3�?UJ ?;,��H������Ja����:�yr=59r>o
羶�3���>��E?+ ?f�>�Q>��0�����c��J/?1֙?���?B��?ZϏ>��Q�0��!������KSV?,#�>�¢�p. ?�^�A�9���^���K߾Y�����I1��������O����"����=�)?@zv?2h?��i?�Y��f���U�����c��H���PV7�XbA��-�j��?
�۾{r���t=�f���I3��F�?�?T��"��>����#D��8��H{>���Y�����<6C�!r=�=�:��?�fP���y(?W��>W�>,�1?�K�Ʉ:�<�$�؈;�s���\=>�N�>���>b��>��=}H����빾鐾(�q�u>�Ec?$�K?�7n?�R�T�/����o�!�S�4��'��T�D>��	>ES�>C�Y��/�|W&��w>���r�d��P���E�	�6�=��1?�g�>��>��?�?x�	��ɬ��w�q�0�ة~<gݺ>-i?-��>#ą>:�ֽ{� ���>��k?G �>�Ǡ>\��������{��G���<�>~��>W� ?�_>tn7��I^��Jy��VG8�ћ�=h�d?|��pa��`�>�#G?������<�>�>��D�"��F�IT	�>��?���=��M>Doƾ68�?���X�2)??����-�*�U|~>E6"?e0�>8s�>��?P��>Ξþ�>�zs?��^?�KJ?^8A?��>V=Yc����ǽ��'�ܒ.=���>O+Z>�Op=���=����"\�L!�<�E=�S�=��̼����j�<A���!�J<���<s�3>��ܿ�1I�!Ѿ"�
���߾={���x�B���M��sת�� ��I~��I��%��OT�eVo������_� 4�?kM�?�v}��u�O3��ѧ~����L�>Ȉ��W�����ͽ����&�Ӿ�~��Wo �~�O��g�M�c�6�'?�����ǿ�����;ܾy! ?@ ?��y?��h�"��8�� >5�<M3��a��[�����οA���y�^?e��>�
��>����>���>�X>DIq>����䞾�{�<{�?�-?[��>�r�O�ɿ����Φ�<���?��@0}A?D�(��쾅OV=b��>"�	?w�?>�W1�E�����I�>�8�?���?�>M=��W��}	�v�e?��<�F�Y$޻k.�=>�=Y='��|�J>�S�>|�SA��Bܽ��4>
܅>��"�'��̇^�)�<��]>��սC,��o=�?�8�����K,�U>���Ң<��'?�\*?��&>�G�>9M���˿oB/�mv?'�@I��?���>�پ��?��۾!�h?4sL?[�&>,a���e�a�*>XԀ��B��_�z�Q�/�=ѱ�>��o> 2*��� ��O_��s�=��>��֬�� h�H�DZ�=Qٿ:�l��s��S���_���H�6�(����+=�.�=e=>��D>5-X>�qo>_e?|ч?;��>�N�>R�1=���ٖ���F�Qؾl�Z�;�n��_�<^�����R�پ$��}�+����P4þ=�E�=F3R�-���� ���b���F�B�.?4_$>��ʾ=�M��&-<�rʾ�������	ͥ�k.̾L�1� n��ʟ?��A?����'�V����*C��{��{�W?�W���x鬾ߩ�=�ڱ��Y=	�>xw�=��⾒!3�@S��`0?�P?^7���Ð�R+)>09�`=,?>�?t@<��>��$?��)�+|�5b[>�i2>��>0Z�><>����۽N�?[�T?���E��rב>���̀{�H�Y=4<	>~�5�F����X>}�<������H�]y���Z�<SY?#�>�*�D��X4��`���Z=�=n?�T?���>�)q?e�K?��=���{V�`�"w<z[Q?C�o?�E>�َ���Ծz ��;r5?ob?&h>�=|��'پK�,�?��� ?�Wo?m�?�z��Y�u�r䍿x���O5?z9w?��k�O,����
���\�6�>]��>���>k2��ʵ>��1?����ړ�����[:��4�?��@��?|�(������m�.	�>���>)�&�c���AD��Ц��B=g��>�����?������N�V�N?��?@��>������
���=�ٕ��Z�?i�?����VKg<���l�o��,y�<�ͫ=��_H"�����7�j�ƾ{�
����⿼٥�>.Z@�V��*�>�C8�P6��SϿ'��h\о�Sq�j�?T��>�Ƚ���'�j�\Pu��G���H�Υ��tH�>��>�I�����{�\(;�����>;����>�hS����:�����1<��>���>l�>����۽�A��?�]��G4ο����ӗ��X?�T�?j�?vn?��P< �v�e�z�:��6G?�Us?�Z?uT&���\�s6�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�e�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�d�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�F�c?cr�1�� 1)��o���>+�B�(���x꼧f-�_��$���x��v"�?eU @�_�?���(�u0?P �>�ā�lܢ���v<��@>��>u�_>K$T�&˚>=�#�V�A��'z=~��?���?<�?���$����=t��?�[�>(�|?	��=�?�N�=Q�ľ*�/>̓}>��N>I^6��y�>�{.?7_�>Ġ�=ג.�W.�"!9�~�s�c�$�F��>>h?d�Z?��>5A�<m��=v2�7.�N�h�I~�=4O�]!&�9����i=��=��<>�j�F�����?Mp�9�ؿ j��*p'��54?/��>�?����t�����;_?Nz�>�6� ,���%���B�`��?�G�??�?��׾�R̼�><�>�I�>>�Խ����\�����7>1�B?[��D��u�o�z�>���?
�@�ծ?ki�N�?������G�}��iT�C���l�#>7'3?ľ��k>[�>q�>>�'|�,����l����>À�?���?���>j�t?QA���Z����=7��>�ф?�� ?���������>���>�Y�oUU�i|����e?��@��@�pG?�i��p���Т��V¾�lо��=�s=��b>y��<��=	Z=���<w5�r%>$�y>)L�>�g�>�{>VX>�z_>�ق���"�AӜ��c���'�˾����ƣ�٬ھQf*�.��`>��ZU���a�������?�;�'��	������<�=Gsa?q�I?讁?�]?/]�[��>Aʸ��D>��W�1�1>�6d>OcO?�R?���>�B5�&"~�d�Y��,}�����Y.E�zv�>9.�>���>*!�>���>�����G>��>�ƈ>B�=>B]@>2�p>���=�>�S�>�T?&�>�G<>Pk>#ƴ��-��a�h�.�v�I�˽���?����m�J�1���U�������8�=�b.?�>����<п��o.H?�����#�y+���>Ŷ0?mfW?��>�$����T��->����j�e|>�P ��ul��)��.Q>�f?j�m>@�%>�����K��&������t>�G?��뾯���O����Q\�=��i��=�� ?��>��� ���AY�W0i����<�%+?H�?|�����0ua�b�c��q(>��>��>@Ƶ=��S>񰽽�J��W��ų�=m��=�I�=N?��+>3�=���>�L���O��j�>�B>��+>��??� %?���)P��қ��M�-�w>�,�>��>�>�(J����=\�>l3b>���[��0��A�?�pW>$�|�9_� �u���x=�{����=���=,a �;�<�=�%=e�~?߀���房��q��WD?�#?̝�=�nH<��"�=����g��O��?B�@�s�?6d	�y�V�~�?�F�?�7����=V��>Dë>�;�L���?�ƽ�ޢ���	�P9#�`K�?�?0�ȋ��l��8>Ib%?֯Ӿ�p�>�o��X�����W�u��#=E��>!1H?�D���N��=�`
?�?�b�Ω��M�ȿ�v����>z�?��?.�m��@��b@��}�>���?JkY?�[i>�X۾NjZ�၌>�@?�
R?&�>95��'���?3׶?��? G>�x�?��r?}�>�!��ҷ&��|��0����W=�2)�;m�>9�=U�ž H�������+�j�����\>R�-=l��>k{ԽY����Ц=[N��uO�����J�>��>�lE>�E�>���>���>嫝>�J=,���aB���3���FP?W�?N��{WP��ǽr����n%-?��K?�|F�B�׾l��>�h?o��?��E?\�>�$������Yÿ��;T�=���>.c)?a�>�rp�Q#u>p�Ⱦ�����>�D�>m3!����E'׾:�4=^;�>[�?֚X>"�>�1+?��?L�>� 8>�L\��χ���C���>��>��Y?��?*�1?BȒ�tD+�9����_��z|���C>��?J,?۱d>�u��53��0�t��]��D)�=�HH?[{?��<!?�9�?[�U?�#?yp��ʾվI��8��>J?6�1�Jd.�!6(�:��B�?-��>�Z�>�ƽH��)���B(�������>�o\?�� ?�����e�i��j1=����>|�<5o�=�ȣ���->j�D>�م�Z?I=.�>5N�=�v��GZ#�a�/=G4�<�}>��=�=��<�+?��D<���ˮ]>��\�,�a��=�r�=�(��Ѳ6?���W�v������������<�?�R�?�Ţ?�H�N�f�WYG?�&�?���>C�>
vO�a4Ǿ�G���������#\���4�=�ҟ>b��,���!����\��?�v���*�i� �H�>� �>hp�>��>���>��F>¾Ͼ/���
��U��o�X��#�J�����P%�D뻾�C���3�"������2M�>�\_�~%v>x�?ߎ4>DĲ>s_�>xN->uq�>)�>�">'�>hB�>�>>|Z�	Ղ��KŽ6(U?�9���&��𾧂��v�??;La?��?���<I/���B	�J�?��?�՞?R�d>�!i�ڝ+�Պ�> S�>�ǁ�z
?)h=� �=���<�ѾR�+����;F�W��j>G.�MF�ANN��*Q��_?4?��M��$˾X_!�F�-�=mNx?��N>E�⽖�1�VɊ�׶y�j��#�^>s!��e����f��qc�����le�1V��Rd0���� �9?og=?\~%�GX.�-�f�(�M�,�-��a�>��?k��>� -=G��\��I6��}h�/���~�p��>w�|?�H�>7�I?��;?��P?�L?���>�^�>	x�����>��;Pf�>Yt�>��9?k�-?��/?l?*�*?`>�q�����N{׾]2?.�??�)?y�?����ýβ��EU�11x��>}�ZY�=qS�<�ٽFWq�}q\=l>T>CX?֛�"�8�����;k>��7?�}�>m��>����-�����<�	�>u�
?�C�>����1|r�jb�oQ�>���?����c=��)>��=����Ϻ�_�=���*�=�0��[x;�?�<?��=���=N�u�b������:�Ƈ;Bk�<M� ?ZJ?Je>�N�>�R|���ﾙ���N=B"d>�)>��=�?�:��������j�]��>:�?��?���<���=�>s������Lb��������<kv�>�?3�C?6T�?�T8?��?�a�=��
��4���6��������?" ,?���>���)�ʾ�먿��3���?�d?� a�a��'.)�Ƈ¾y�ԽE�>�O/�['~�� ��+D�尌�����n��9��?��?y@�Z�6��8辮���>l��wC?d:�>p=�>���>��)���g�L��?;>1u�>R?W#�>i�O?�<{?~�[?�fT>�8�1���ә��M3���!>J@?���?��?|y?5t�>��>_�)�Z�eT�����3�8���SW=�Z>*��> (�>$�>���=��ǽ�Z��^�>�ra�=M�b>���>C��>��>��w>K�<.IH?t�>�ľ�Cτ�V�⾪R�Y-?�̆?�; ? ���/�-�gY�QfP>ܭ?��?8�I?YYþӳ>�j=ch����$��˼>�	?v�>y�$>��>n��>m�?���>�'�����I���=H�!?�S?_��=�uĿ~�\��\��-����=���X����F��F���}=��z���d�O-���(�����rX����ž���m/���?3��=V�;>i
>=�9Ӥ���+�<��g<3C��(�l=�)���B=���V,; ���t��-<����ݽ�ξ)�z?pjI?��*?ŭB?f��>�44>��N!�>��a�?�\>U�Լ�+��R�5��u���̓�k�;�mϾ��U�Շ�����=I!�<��=�-%>���=/�<�ں=��N=]n=�w��f��<�G�=�$�=��=9 �=*D&>`>�}?������B�M�5L=x�?<V�=o�>�w���5?'�>Gpn�08���x�o�p?�g�?��?�,?�����`�>�m�������G>�o����=Kn=��>G�>�SY=N��g�� =��?m�@o*?[��
"ֿ���>k�7>��=1�L��l4�TG���S���W�i$?��:��bо�m> ��=�ྀ^ɾ�=�A>UmQ=<6���W�ѕ�=z_��:�v=^��=멇>̾c>B��=:���~�=�=�>��E>���;�G�Y�e��y�<�]�=I\c>�s>*��>��?e60?�[d?%�>Ao�nqϾ~���3�>��=�K�>��=LB>u6�>q�7?P�D?&L?���>L��=�	�>��>�,��m��.�����m�<���?�׆?W4�> �S<L=A��l�Ue>���ƽ�?GZ1?{?#˞>p����(&���4���j����;�2=��3��FҼ�����Bܽ�m��">���>�o�>���>�Nn>�K>��a>�`�>l�=(��<P-=��y��<�;S�e����<����pO�<�2;�:�<��X=�y^��m伳�l<�,=�/�<�(6<�>�`�>��
>��>Pޮ=ҏ^��
�=,%Ծ��9�*[���}���8C��uY�󃿂z4��ZQ��z>S�>��������P>?uզ>~΢���?h�z?=i >��d�#g�L��װ=�mB�$o�<��=F�\(m������k��������>��>��>��l>�
,�8?���w=�⾨`5�]�>.w��&��/��:q��>������i���Ѻ(�D?�E�����=#~?h�I?)��?���>���I�ؾ�00>$E���.=/��0q�f�� ?Z'?���>[#��D�m۹�$Ԅ�OL>�߾79�������I���V�O���u��>��о�2����g�5G��)���i�?��֞�t�>��e?@x�?O���$����-��7v�Q���R?D;�?h�>��>��?��>PR��C��:K�=��r?���?�f�?�>�#�=�մ�CH�>Z	?���?���?wvs?c�>�\�>w0�;y� >kǘ�؈�=�c>o�=P��=	V?s{
?a�
?|��	�=��G���X^�V��<��=Yo�>m8�>�ir>0{�=�Af=t!�=;B\>;��>c�>��d>��>*8�>m!��X����!?FLl=N��>=;??�TH>L<�=@���S��"��fPu�(YS�c��."����<#W��eE�^8����>8���]��?m3g>E%��q?'B־1 ��RbE>P0�>��཭~�>��S>3P�>�Ŋ>�B�>���=��>Rs>�����>�-��v� �us=��6��Q��\^>^h��d��a�����&k�"ó�Vv �1�b��.��Ė<�?%�<���?� �Ils���-�������>��>�2?��E��o�=�X">�^?�.�>3�޾Ϋ��� j���?KT�?�N�>��
>�?<w*?�Xa��^��>��9Z��_��<���]�����d���ξF����Z?[t�?�;*?ش��q{>�s@?[��2ú�q>�UX��sm�Ғ���h
?܊����T��0O��bv��<��e? e�?�'?ܜ���A����4?6Z{?c�]?\/9?;'I?l�h?�����!?���>AfG?8� ?�o\?lN?K��>RXB���=�O>�.�>&Խ��q�'�ƽLB��A�<��'=�����گ<}Z���,=�hS<���<�4��|�	~�;#�=�ע<!�>" >���>�lQ?��>z@�>�M1?�3%���:�c��ޒ0?�X=����s���㡾�����z= 
t?�Ѵ?�h?t�#>��F�0�
��P>�#�>O�>�I�>�2�>�7̽�1G���*=��M>�+>v=Kj��������F��B8M=�`5>�i?d�	>�!��H"�����u9����N>>@���IӾZ羊�^��CP��B��'��>؈o?�)=?���<�9�f��=G]��7L?1�W?�?A��?&!L=����V&�'e���νH >x�.=��+��'������5��<��W=^���4٠�_�c>�^�b޾�:n�~+J�����;?=����V=���v�Ծvs~��a�='�>�F���!��&���Ϫ�[yJ?�Ak=8̦�cX�Z)���Q>��>��>t�=���u��@���z�=Ψ�>�9>�ڨ0G����9��>Z]?�Na?��k?���nU��7�6V
�I�������
�>��>-��>y?>��	=�h��VN�-�h���n����>��>f-�N�W��CᾀO侂��Gd�>�?6�>TD?�rG?��?:i]?��=?	�?;��>׼1��m�*?��?9��=�l\�Ir����*�	-C�M�>��5?ĝ��~�>m�
?߸?&?FYN?��?r�E>z����N���>�V>z)^��ӱ��ߢ>��??�'\>W_Q?���?��>v(�np����T��7*>�j>�1@?�_)?�?װ�>s��>&Ɨ��4�>�t ?�,?���?\g?�{>���>��D>}k?OC��x�?l�	?`<?�^0?�e9?-�S?V�>#�;M�뽯H��i4G��4�н��1�:�5�*�ֽ�;�<KV'>g*s�"�ټ��ڻV-�o�μMh�ë=�_�>j�s>+
��f�0>F�ľ�O����@>쇣�%P��$ڊ�9�:�c޷=5��>��?#��>�X#����=/��>I�>6���6(?��?�?k�!;��b���ھ��K���>"	B?T��=��l�����q�u��g=��m?s�^?��W�l&��L�_?>g?���Y�2���K#���6���.?qN?�T�\�>��w?�=n?��>��F���1����h��c���M�=ӡ>�	���V�9wq>�%)?���>��>��1=Tվ=�u������G$?���?Xȵ?���?�� >�+Y�����Ҿ!�����a?9�>����a1?��R=e־�ܦ��þ;������ƾ�d��3�о�KĽD������n��=?|�H?��\?;Q�?����W� �q��ـ��_��ܾr�۩L��%�P/��ʐ��;�Œپ����d<Ɂ���j7�Y��?�'?�1%��1�>���iM����˾z�/>�Μ��+��ڛ=�@W�1*=Ȣ�<y�%qW��幾=H$?��>�
�>��9?�7U���>�Y�<�X�G�����|S>�
�>$ѣ>A1�>7�	�� <�1��Ӿ�������>"�?�?j~Z?��9�ɞ(��[��Ω:���=)e��A���W�=N��>���Vze��'c��q'�Z%s��+K�֮��r��wD�>0}*?1�=�P�>V3�?�x?�uP�9��� ����b+����$>�b?��?�tB>��"�t�ɺ�>B�l?d��>�>�����Z!�0�{�!�ʽ54�>�׭>ǥ�>$�o>ǧ,��"\��k�������9�Q=�=ݢh?������`��߅>8R?��:�zG<F��>�mv�B�!������'�A�>M�? ʪ=?�;>c~ž� �2�{��I��	G)?�:?/���ڀ*�:~>',"?�j�>@6�>q(�?[|�>3þk�V��?��^?�GJ?�SA?�Q�>A)=�����Ƚ�&�,=㊇>2�Z>��l=I��=M����\�����<F=~�=�*μ�y��Ú<>,����K<o��<��3>��տ�>�nּ�����y�ھ�����JS���w��6�����s����r�mԽ��z��(~��`��(�����?�>�?��$��(���������z��-!>`��ŝu������𽿪��zYӾuU��s
"��*T������g� q8?x/z��῍r��5p����?iΪ>�ȃ?�03��ؾ��R�j����^�:5��7� 
��'�߿`�*%h?f�?�����)����>��2=q��>@hY>��u��/W��O��34?��:?4s$?1���<�ɿ�Yɿ>lT�?��@�|A?.�(����V=[��>�	?��?>:W1��G�����$R�><�?���?�M=T�W���	��e?vS<G�F���ݻ5�=G?�=�F=���6�J>�V�>��HWA�n@ܽA�4>hم>�i"�٨��z^���<Ą]>�սwE��5Մ?*{\��f���/��T��U>��T?�*�>b:�=��,?X7H�`}Ͽ�\��*a?�0�?���?&�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=S6�Z���~���&V����=_��>a�>ł,�����O��I��Y��=����f¿L/�2����A��j&��
j�e{q���L��ͽ_W��Wx��f��cc�=��=�v>���>6N>�R2>S�P?$�?m��>��I>��̒���� ���ټ�g2�x�"��j���d�z8ȾGE��m������� ����־��;�H��=�Q�P6�����fd�*�H��+?6�>z�Ⱦ��L��!�<�ɾ�^����ż1���>5Ͼ8�3���m��z�?6�??w뇿�Y�=���S�k���;G^?x���I��+�=��
��
�<���>��=�-�3�2�Z#Q�;?��,?��A�m��>���v�v;`�0?x�"?=U>�{�>��4?�@���޽�<i>�M�>���>���>���=��̾
G���?R�w?�K:���ľt��>�������ΝB�B��=��;"�>�c�>W#���"ܾ�S=�u�����<�(W?/��>��)�m�t`������R==��x?�?�1�> {k?��B?���<�g���S���!xw=k�W?)i?Ҷ>􆁽оK|��z�5?��e?��N>B_h���龽�.��T��%?��n?d_?�����w}�������Qn6?M�|? gC�윿���4վ�6�=���>1	?ʺJ����>��<?���#ә���̿�H��ؙ?��@|��?�w�=X����zK>��)?��>��y����QF�o���� �=f2�>��;����2?*��s�h?���?�?v
s����*o>h����?7�?־2*=�X�׿u��>�������jވ����ݾ-V�9�ɾ�0�.ɾ�:�<]T�>�@�:a�W�?|O��2�3ֿ.��� 0����W�!/�>}��>\$���� l�ԇv�� 8��ch�B$��혣>���>���iԾM�p�?���J�7z�>�cؽ�\�>����> G��&��x]���*>���>>������	��Z�?+@��F�ܿ����(��h�4?�ۏ?���?��%?�s>G�z�_�$�u�O!0?�gz?�:�?[�����+����=�Ep?���Irl�>�4���M�?��=��*?e:�>��;���<�E>|�?���=w�H�:_ĿB"��/�׾�(�?���?V �ix?~E�?�n$?'�(�� �Q���Zr)��<����C?��S>g�ݾ9�2�?
B�A���-O ?�UV?��M��#1�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�"�>T�?���=`d�>9�=$簾�T.��D#>��=]_?��?\�M?�A�>L�=�9��$/��TF��HR��.���C���>��a?uL?~Cb>�︽�1��� ���ͽ�p1�Pb�FG@�"_-���߽5>D>>�>P�D��
Ӿ�O3?��̦�S����E�1�?�FC>�.(?p���k���X�䫀?2�f>?k6�����G���C�c�k�?1�?���>�ޱ�1H>��C>"�==�޼�V=Tb��ʓ��<�=d�s?�2�ӯ��ԃ�\ۂ>�þ?uL@@��?��j�D�
?�r������}�r��}�D���=<�:?0����q>3�>:�=�'w�-��6u��=�>�Ư?���?��>�i?�k�|<�<�5=*��>��d?L?*��#���I>�2	?Z��᏿����?d?&�
@@/@��_?�᣿��ܿ\��ھ'վb �=h\<�Km;>:����>.�=��H=�0��I=A~>dY>�#>Z�>�;1>��>5�����ԛ�I�����A��,�cL���Ž0�澇7<����f8�@p��  �=aKl�<ǣ�^n����Z�pv;���=]�U?��Q?��o?A��>M7v��>c%��cH�<�$�4��=0Ӆ>2?!�K?��)?P��=E����d�憁�xk��������>��G>�5�>=��>�Ů>��:"dG>�=>�*�>� >Ć=��L�=�UP>F[�>v7�>���>@{l>�P>�L��J
��k�,�T0���/����?~#վw�5�@	����*�����{{;�A?-�>	C���ٿ�o����U?h���c�2�O$�OM^>NG?�vZ?�j>5��v��=��{=H�˾������=�TҽR�_�E�5��B >� ?�f>@u>U�3��d8���P�Q{���g|>x26?b鶾�G9��u�^�H�}cݾ�DM>�¾>HED��k�W�����ui�R�{=:x:?��?�;���᰾̭u��B��KQR>�9\>Y=Ul�=yVM>YXc���ƽ(H��i.=]��=��^>V#?�*>��='�>$���"�M����>�)C>�D+>�@?�[%?�������G,��v>��>�q�>�<>k�I���=���>z{a>6@�D����x��?��UV>�z���]�cq�au=�ؘ��3�=h��=�; �Ug=���'=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�k�>9z�\�������u���#=��>:H?;Y����O��>� w
?�?�a�M�����ȿ�~v����>�?@��?��m��?���@�Uy�>e��?�gY?ti>e۾snZ�ޑ�>z�@?�R?��>�9�6�'���?H�?���?U��>���?��?��?O��=��%�v�ʿ�@��C�?����([����~>����!��&@��}��ZuI��~P�h~�>5m�<�X?��^�lN$���)>d��<Td�������.�>�s�>TV�>�BE>W#?La?s�^>�c����=��&��YI���K?���?0��1/n��L�<O��=9�^�� ?FL4?��[���Ͼ6ը>`�\?���?,�Z?;Q�>���)>���迿^��p��<��K>76�>�=�>���/YK>�Ծ�ND�*m�>Η>�C��8ھ�,������G�>�a!?_��>���=�� ?�#?�j>��>q0E�_G��4AF�=Z�>�q�>��?J�}?h:?.�����3�����ʡ���[� ^L>Gzy?.?/��>ċ��>����X)��DD����em�?�g?�F�;?E3�?{4??�,A?[�f>���ݟ׾Y���'��>��!?��A��K&���&?�P?!��>�9����ս.�ռ���jz����?�(\?�?&?6���)a�j�¾�7�<
�"�\V�d��;L�D���>i�>9�����=�>�۰=�Mm�8H6��f<\e�=�>���=417��|��� 2?�)=u����;J<"�����j�]�{>mAY>޽�VC?{�-� _�������������n�?R��?�{�?�+���p�4,9?�A�?���>�?0򐾂^���$� 5~�&}������}ܼ@�>Ws�=BFᾼ���:��x���� ���ڽ��?�а>H5�>�S?��<>P��>����a�+�֠'�����k�l'0�wV?���/�Ά"�hw���������ʾ�܆�HǼ>;@Žs&r>��/?cv`>E��>��
??~���O>߱�>�P^>���>H��>E<>&=�����-��KR?�����'�y������f3B?�qd?M1�>Yi�6��������?���?Qs�?0=v>h��,+��n?�>�>D��Rq
?pT:=�9�i:�<V��s��3��[�3��>�D׽� :��M�2nf�rj
?�/?�����̾�;׽�N~��)�=�bc?��J?EQ#���q�r����ڎ��2��S�[�Ͼ�p^�t[�f�!���%��N5���ZY���>�4?U�?͉5�s���0���Iq��q��c >�?�N�>l5�=%�?b��m��87�ǟ�ܸz��́>�}?�i�>sXL?ئ_?�Zt?xe�?���>=?����`�>X>��>��)?:�6?F?��B?��;?��I?�s�>ω[�RD�@V��s�'?5��>�?�r
?��?����V)��3��K�=���,>y�=C�>PHZ�~���x�>o=�=wM?Ȧ�{�8�����	�j>ۅ7?,��>���>V��� ��$`�<��>�
?VR�>�����jr�:S��]�>��?��G=�)>A��=�cߺ=L�=������=����q:�|� <-�=��=tz��Q��-��:��{;z��<�u�>y�?���>C�>�?���� �T���h�=�Y>� S>m>�Dپ ~��j$����g�7ay>�w�?�z�?Y�f=a�=y��=|���R�����#���h�<(�?+I#?sVT?3��?��=?�k#??�>O+��M��X^��3����?v!,?��>�����ʾ��Չ3�ם?e[?�<a����;)���¾��Խʱ>�[/�k/~����>D�����_��6��?쿝?dA�R�6��x�ٿ���[��x�C?"�>Y�>��>V�)�z�g�o%��1;>���>jR?>$�>B�O?#8{?��[?�{T>ܕ8�b-���ҙ�'o1�h�!>q@?��?U�?�y?�l�>8�>��)����^�������Nւ�W=h�Y>���>l*�>��>���=��ǽ+^��V�>����=ɔb>Е�>s��>\��>��w>�9�<*Z?i�?�����5�\GH�f��	mz�^nD?��?��?��7<���4�z�԰���>���?�?��?���A�	>��׽�`��T�O=���>��>k8�> >��=6&�=T�>R��>�`���'���#�am�x�?�6?@�w>�ƿ�q��.q��2QZ<�����d�5����Z���=}���o���i����Z�&Y���z�����X�����{�.��>5*�=vp�=q��=�c�<�x˼;�<�'K=A�<�/=��p���e<� :��dԻ�䉽� ��X<��I=r=����Ⱦp�}?o?I?�	+?aA?!�z>[>i2@�zM�>�w���d?��Q>!�V�󂽾">����C�����پb�۾L�b���>� ^���>�,2>��=���<7�=1�g=���=�:��=���=A7�=��=��=z>�a>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?~�>>�2������yb��-?���?�T�?>�?Ati��d�>M���㎽�q�=F����=2>o��=w�2�U��>��J>���K��H����4�?��@��??�ዿТϿ7a/>��7>�&>w�R�E�1� �\���b��xZ�՚!?�H;��J̾6�>��=Q+߾�ƾN�.=ք6>T_b=Th�pV\���=��z���;=-�k=0Չ>s�C>�x�=.���=¥I=���=��O>�v����7��(,�Q�3=���=�b>&>!��>�?uZ0?G)d?_�>b�m��Ͼ�<���g�>���=�-�><��=qOB>T��>�7?1�D?2�K?�k�>�v�="�>��> �,�$�m�9.�ٱ��$]�<���?�ӆ?�M�>�U<I�A�T��VA>���ý��?�K1?w?k��>�^� ӿ�w(�y�Z���׾;[w�8w=e�鼵�=�%Xɽ��<{DM=�zM>�h?��>i�j>bM�>��n=��=���>��>^ݖ=��>�%D;���=4�ü�<~<K�o���ӽ`���=��=���~�/��S����=�Gw<���+>���>蔶=��;>��>׺	���>М�p�U.��|��ŕt�J��>z��b�O�`�+��]>��>���=)�����>�D>�~�=��?`��?@�>�-�A*�����4����@�t^�=bC�>"�<��L�艇��zc�2�˾Z��>g�>�>��l>�	,�#&?�8\w=��W5�0��>和�_��@@�@q��?��b����i��L�J�D?�C��	��=I~?��I?��?���>�H���ؾ_W0>E��6=g��4q�Ȏ����?�'?���>~��D��J̾�I���շ>�3I���O��ŕ�&�0�^*��﷾��>Dݪ��о�3�b^��������B��r����>A�O?���?B(b�j���xO�.��qB��Gf?�g?9�>�<?�?�Ġ�*��Ϣ�����=��n?s��?�*�?>t�=�X�)J?RI?sF�?&��?��{?̦����>|�N=�b>�5޽od>6�F>��/>;�/>(#�>+�?W>�> �����$����]�Wv��:=g�0=�Y�>`l8>N&>��=���<��=�a(>ߵ�>�L�>4�L>���>��>瞄�L��	?wq����>g#;? v�>W��<%���l�Ɓ��~�M�3桾-�񽋒�x��'D%�O46>ӮU=ѻ�>uͿ��?��>z�$�~(?x4����	���)>�Р>�H���>
��>(�>��g>��>�y�=��><RR>EӾ{1>�V��� �<uB���R�cwԾ!ur>N�$�K�h��(�G��9�����+j�P>���=�6g�<΋�?�a���m��++������?�Ψ>Xi7?��������D>���>'��>>�������e���r�྽��?�]�?�;c>�>P�W?�?��1�N3��uZ��u�.(A�?e���`�T፿ߜ���
��	��F�_?y�x?*xA?D.�<*:z>*��?n�%�3ԏ�w(�>�/�w&;��@<=�+�>P)��O�`���ӾB�þ:6�JF>��o?%�?'Y?�TV�c��=	K��{1?��#?i��> BJ?!\=?X�>1��>�V�>��U?��e>�N?�'?�/?x�g=��="'�>�{=h�v��OU�\y�Ԍ��7��g�9�^�=?W�=��=.gW�*ñ�^½Y4B����;����-���V�=��L��`}=>�>��^?.�>.Xt>�+8?����&9�jE��Ğ8?�H�=��x����+��<1�:E>��r?d=�?yV?1pS>FB��GC��#>�]�>Q6>�JM>�ݼ>�k��^/O�H��<ە&>��.>XS�=hܐ�r��Ob����k�=�b.>���>C1|>���r�'>�|���0z���d>��Q��̺���S���G���1�|�v�?Y�>��K?J�?U��=y_�J/��`If�0)? ^<?�NM?��?"�=�۾[�9��J��>���>�X�< �������#����:�m�:O�s>�1��.Р�\ib>��� x޾��n�XJ����,dM=�|�WEV=��7�վa*�ǜ�=e*
>b���S� �|���ժ�8.J?��j=x���rU�c��,�>��>�ڮ>c�:��v�l�@�6����G�=8��>�;>覙�����zG��:��>N�F?�AL?H�?�%����m���4��j྆�����*�b�?�g�>ɜ�>�>���=	޾=��Rz^�h�����>���>a�)��?`��嘾���1:��(�>]�?��j>[�?�`?�T?�^]?��&?��?���>��7���پЇ'?Nރ?�S=i潔�V��8�pXG���>b�'?�`C��P�>�?C�?�%?�1Q?Z}?�>����A���>���>�V��ﯿ)li>�H?-g�>7rV?��?��E>�I4�].�������=Uf+>�z4?�#?�??kX�>w\�>���n��=��H>�5r?��?F|?��->S:�>z�M>���>�/9>&*�>�{?��?o�W?��p?w�@?֣�>�ɟ<�뫽|��E�ѽ{���������;N.�<͛l������@<an�=,��:��ɻ��<���֏���9ۼH&���_�>B�s>�	���0>��ľ�P��)�@>�����O���܊�œ:��ַ=ς�>r�?D��>Z^#����=׮�>�K�>��\6(?��?$?�4#;1�b���ھǴK�u�>�B?���=�l�̂���u��h=��m?��^?�W��&��>�f?|d?(Z�J(��t۾sȈ����.b??^&?Y$��^}�>��m?ĊW?>w�>�9�n�T�Ct��Ζj�-�x�M>���>�e�7��.O�>A�+?Yi�>"^;>�-�=�m��U\H�6+���??��?@{�?\�y>Y_��鿲��z`����q?���>XН�4.(?�h<Ͼ�󠾿P'��Y������6������!��fV�0�=�j�=�t?�r?�d_?��f?�m�h�o�0�d�6gx�'�R������%@�l�:��V�F*^�~�)�&	�*Y�\:<v�p���F�t��?["?�z(����>����r�CDξF;\>������"�m=������4=�<f=S[��,�q.���L"?�޲>_�>v�@?4`���=�Rv1��<����>�(>G�>�k�>��>�;��D#�����iԾ>I9��͐>"]?��,??z?	�H�I"�s|��!�����)���O�>��=f�=G�W{ƽs<�lxX�C@O��f���	R�z+:>DM^?">|�>�?��?���'�#�|���"A^���Q>�?��P?�3�>4/�>dѽP����>��l?ۺ>C��>%���iE������I.��>���>A?'�w>栈���e�$,��t�����G����=��k?Fń�*P����>�)L?Y�Y��<���>�����a��p޽J��=�q?s�@="�~>��������$y��v��Vf'?��?�)��k1��d�>��#?���>u��>��?�>�P��d�(=��?��_?��N?7F?�g�>G<�:нۉѽ�R'���=	�>��Z>ָg=�+�=S�"���F���"��P=F��=��H�m��\��<9�u���;��x<S3->4׿��N�%ľE������|����3���m���v��"&��ir̾||$�:^Ƚ`�A�?����o4��X�����b��?���?S��x�V2��ex�����ZN�>��žNi��ݨ�B@����~���Z���4�Xw���`��&U��'?������ǿi����ܾ�?h ?��y?*��S�"��8�͖ >s��<�K���������4�οfA��H_?���>��ﾉ~��h��>kՂ>>aX>�p>�����ʞ�@ �<p�?K�-?6��>͏r�҃ɿĈ���8�<��?��@�|A?��(�����V=���>I�	?��?>7T1�nI�����T�>x<�?���?�M=��W�>�	��e?ej<��F�Q�ݻ4�=�;�=D=j��B�J>zU�>L���SA�->ܽ7�4>�م>��"������^�]��<2�]>�ս�:��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�����ȿ��1���v�=؜_=�mk="d�.͎:��G>'f�똯���X='�{>���*>V}?Ⴭ>Z5�=�U?inb?�t�>Mq8>o-��S�˾�y�}���$�j�\��i����W�۞��F���Z�p6�{c۾�y��q=�}�=7R�x���� �Q�b���F��.?w$>#�ʾ��M��-<�nʾ����܄�l⥽.̾C�1�] n��̟?��A?������V�#���K�����N�W?�K�q���謾/��=ǆ��J�=r&�>�=��⾷3�]S�B0?`�?�����ڑ���)>=Z�0�
=��+?��?��e<d�>x%?�$)�S��]>�5>�j�>�K�>c%>*��X"ܽKt?�T?�Q�����ٹ�>����Mhy���]=�s>��5��ټ�\>���<P����_������<i�^?T�E>,�3�k*�a���\n���=aȌ?�T?<��>�<R?��?;�Ӽ'���Cc�hH����}�K?V�}?eF>U��2�/A��3�4?�D?�=>W(پ�E���gA��2�EF?��?�6?Ϙ�{�}��B���U�6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������7�#>���.��?��?C����<�4	��m�� ���==&Ľ���<ڽh���6��0־<���m����W<���>��@�b��}�>�2~�ܑ꿠Aɿx�k�qž����0?��]>��i�p���Yr�����7�O���0�Q�=����>�>'������D�}�x�=�������>�����>�NB������ٝ��oq��k�>��>y��>*ߪ��A���?o��#ο�I���r���W?>ҟ?{��?��#?��;��y�q�v�{���pE?��p?�IZ?.�/�{W�����l?J*��5Lg�;7�b�M��4�=�?���>s*������=��>�VV=�4��Ŀ��ב����?�V�?���*�>�C�?�1?�B������n���C�BWK�a=,?��n=�ݻ�+�(�:�7��pT�>�L,?#o���c�[�_?�a�O�p���-�b�ƽ|ۡ>:�0��e\��L�����Xe����\@y����?M^�?j�?ϵ�� #�L6%? �>l����8Ǿ�	�<���>�(�>*N>cI_�Ӳu>����:��h	>���?�~�?`j?������U>��}?�-�>��?�3�=][�>=8�=Q��/��K#>��=<�>��?*�M?:�>��=��8�U/�o\F�[FR�/ �ؿC���>��a?A~L?Ib>'���1��!��_ͽ�Q1���鼓U@� ,��߽�N5>^�=>�>��D��Ӿ��?@p�3�ؿ�i���p'�[54?���>�?���޴t�����;_?�y�>7�,���%��C�]��?�G�? �?s�׾ Q̼T>g�>�I�>��Խ����t���_�7>�B?N��D��h�o�Q�>���?��@�ծ?Oi��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*��ֿ٠�|⾠9��g�>آ�=��>�ᄽX_�>�+k>��=�"Ͻ�M�=+��>�V:>̈->^�>���>���=��{�ǘ������r��j�VU��������졾)\̽���������=�/=�j��#}o��K��Q�]�w��/�=5^Q?�R?1/?+#?:x�=���>��d.�=͒��K� >��>[�L?�]U?�	P?:a�>�bQ�"8v�}���>w���ʇ����>��.>?aJ�>�F�>�~�=;+>��=3Ɔ>��	=��⽤M��jw^���>,�>�?묦>D<>M�>@ϴ��1��V�h�w��̽�?a���<�J��1��r9������i�=Lb.?T|>���?пc����2H?����j)�N�+��>j�0?�cW?�>
����T��9>���j�_`>�* ��~l���)�^%Q>=l?��f>�;u>�3��f8�K�P�~}��C|>�.6?-ᶾ�?9�ʷu�P�H�hTݾ�KM>tо>��B��h������/wi���{=�r:?�~?����ݰ�՟u�A���NR>C\>+	=K��=�lM>;c��rƽ��G��.=��=��^>�b?�f,>걍=��>@����HP��Ԩ>QmA>
�+>{@?,5%?��?���W���).�,�v>z�>IҀ>9>^fJ�eX�=ik�>�zb>���ͧ�������?�G�W>"}��M_��\v�\)|=8������=!��=\ ���<�hU$=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>ʝ��G������v�L�=�o�>��H?����M�2�<�?%
?��?C��ʨ����ȿb]v�w��>.��?��?1�m��?���
@��)�>�}�?�jY?��h>RKھ��Z��ŋ>`�@?!�Q?��>t��6'�i�?�Ƕ?���?&�>ȗ�?�G?�N�>s���!��9�������@z;T��<��>��><c����V�[���rւ���z��~�a �>�-�<Ǖ�>�h��$U����X=+�o�I��� �Nv�>�>�[�>�ʠ>�&	?��>e�>�(>�e��Eh���㧾*rI?�ǔ?*�(��a��9�=�� �~�Ͼ�q�>%�"?�qм/n}���?�?ڟl?t��?�b?03�=����0�������a���}>J��>��?�=d��>����*��Q�=���=)/�=��.<��/=kx�>J+�>q6�>oq>:��<�/%?�w?+r>L��>Q������9���>�h�>Y��>t\l?~��>g3�uZ@�T�������TgX��{>�2�?e�"?���>������X�:�d]�?_��~T?{�k?���\?�)t?��?]�?-�1>ڶ$�^��ˮ��d`�>V�"?m�DB���&�����?MS?g��>���i�ֽ�
���2�����Q?\?�!&?��Ša�?\ƾ���<Pf�p����;�t���">�>�݈�)�=�C>�ڧ=Z�h��M0���<s�=>�>#��=�?7�j%��0=,?̿G��ۃ���=��r�@xD���>�IL>����^?ml=��{�����x��!	U�� �?���?Zk�?U��?�h��$=?�?S	?n"�>�J���}޾9�྿Pw�~x��w�[�>���>6�l���K���ٙ���F��^�Žj�����>���>�91?���>B�&>���>�ⰾsF�� ������d���݃2������������Ͻh'�<f#оD2a���>�����{�>FT?���>b��>���>��'��>wɆ>���>�k�>X{>X�D>]NW> ��H�ʽ�KR?����/�'����󲰾23B?�qd?e1�>i�9������v�?���?7s�?�<v>h��,+��n?�>�>C��Nq
?*T:=6��=�<V������4������>7F׽� :��M�Lnf�]j
?~/?���|�̾};׽)1���I=E	�?a�.?B�2���V�|�z����k���]L���Q��.�*�H�f�7ℿӊ��'
u�ʲ��#=`??���?�o�J��7�ݾ���ۄ9�e�>�q�>�/l>�?�m{>�+���Y���h�Ѫ#������f>3t?�%x>�F?��D?��*?Aw^?ծ�>��>v�վ`�>�(
���>��?�D?W�5?dgA?r�1?�'?��=�އ��A��	GӾ<�?�9?L�?�{?X?ΐ��R½X⚼�剺������A�<�����z3�=x><nr>�Z?F����8�������j>tw7?�u�>)��>���L1�����<��>��
?�7�>� �$~r��f��W�>裂?���=��)>i��=p!����Һ4�=�ü���=�s����;�^ <�L�=�ݔ=H�u��d��X��:JD�;̅�< z�>��?B��>!Q�>{G��N� ����9_�=�X>`�R>�>�Aپ���$����g��%y>o�?�{�?�Yg=�*�=�=�����b����P����<ǣ?�C#?;LT?i��?��=?�V#?A�>�)��J���`��5��7�?c<,?�B�>_+���ʾ0��3�dG?�N?Ǿ`���M)��G¾��׽�O>g�/��M~�����ĆC�]������Ҙ��s�?���?`�;��6�3\�T瘿����0C? ��>s�> �>"�)��g�)�b};>/��>Y�Q?��>��O?j2{?�[?f�T>�8�� ��Jә��2�/�!>�@?0��?d�?}y?R��>J6>��)�G;�Rr���]�t*�ճ��'4W=�7Z>ܚ�>F8�>:�>���=v9Ƚl���>���=�jb>�^�>Β�>��>��w>|ή<��G?���>t^�����d菉�ǃ��=���u?x��?i�+?�b=i���E��H��CG�>�n�?���?�3*?��S����=*�ּ�㶾��q��%�>�ڹ>2�>���=!�F=�]>Y	�>f��>�,��_��p8�.UM���?�F?'��=��ƿ�t��pz��/��"��<�ᎾW�Z����:�E� ڼ=����
� ��?��řK�4���l������������a��>��=���=��=�M�<b꡼���<CP=K	U<�G=�pr�P&-<�"!��&��J���&��]�<�1=C����p˾ۄ}? 9I?w�+?r�C?��y>-�>�3�\x�>�Ѓ��%?>�U>��P�����S�;�%����8����ؾ�E׾=�c�C����C>Z�H���>�3>00�=f�<e��=IKr=�ݍ=m'H�[	=G�=P �=2v�=���=�>E�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>ԁ>>RO>/S�^ 2�v�\�]&d�U6a�ؑ ?��9�Z˾|!�>��=�ܾ�eľ�I=:>>wZ=�O �wL]��9�=�n�m�6=F�U=��>�4B>~�=������=QV_=a�=@�S>W	�:�'%�;<�6!R=���=��^>)� >_��>��?�f0?#Qd?�N�>��m��ξ�B��Q�>�~�=BB�>V��=��B>Q��>��7?�D?��K?Jq�>���=�>�>:�,���m��[�3����ͬ<���?ǆ?��>B�O<q�A����K]>�raŽci?N1?x?��>�����4LA��a�7$->gO>�F>�5��T�>�CF>m��՝����>�	?��X>��Y>�?�Wd>^۫<z��>��>Ω ���=Zb;����='�]=Ʌ>S1��Sk=I�k=��6�K�=R�d�&�����~=�= K��c�=(�=b��>sN>�z�>�1�=AU��K"/>�����L��6�=V:��[vB��d��n~�{�.���8��N@>/�X>g�|�?:��U^?0^>�@>ޭ�?��u?��#>�{�V�Ծ�\����c��9U����=�>Fy6�a�8�m^�ƘM�L�վ���>�e>]]t>�/U>��/���G���4<y��O]#��j�>�}�2�Ὧ���0��T���	���<�Y����=`�U?(�����=1��?�wR?�_�?�[?*>�<�=�P��<� ����$��_��/S��;?�5?N�?�$� ]��0��8+ǽ�a�>��.��s]�2���?���1>1����>&���z�ZZ$�6m���`����I���v��	�>�?=?�3�?��_��!��_�N�/%��/ѽ�?6k?Ʌ?9�>�}?�~� 2߾�������	s?�?X��?Esu>�=�Dx�8u?���>���?gڦ?�.�?b���FZ�>�TG�(��=�k~=��D>{��>&�!>uL�>: ?A�>���>���;�#��߾� ���>�s�U>C̺=g��>���=���>���<!>��c>?�>Z	E>-�->3��>	��>~1��:����E?ꬉ=H
�>��5?�F�>��=*a��Z2�=)�s���Խ4����+��I����= ��=��=�7=�q�>�0ƿj��?��M>Z�����%?�ɾ�37=�A>N��>/^'�E"?�d�>h{z>S<�>��t>��(>�O�>�y�>��Ҿ�C>��Zb!��OC�՜R�#�Ѿ��{>���A�%��g��8��}-I�y���Ӏ��j�%���=�o��<kD�?9���m�k�z�)������?�k�>��5?�K���Չ�t>5��>�o�>�.������s����p�@�?���?[<c>u�>��W?f�?U�1�O3�gsZ��u�L'A��	e���`�@፿�����
�����_?�x?xA?b��<;z>��?T�%��ӏ��'�> /��';�5C<=�-�>k(����`���Ӿt�þR6�HF>�o?"$�?tW?�MV�?i��M >�:?I�#?f�w?V�9?��??���e ?��8>��?�m?�3?��0?��?�G>r��=.��&=<ڎ�o��꽏�׽j���(=�n=b���0m<a#=�@=Q���+�ż|�;�y����<>�='t�=�Ƽ=+��>Q�]?�R�>
��>��7?����o8�Hʮ��)/?�f9=�������w�����K>��j?���?*\Z?�Fd>��A�C��>Y�>�y&>�\>�f�>C`�!�E�h�=_G>�>>=:rM�nف�^�	��~��`j�<�2>��>�4|>����'>{��:,z�ާd>��Q��ʺ��T���G���1��zv��Y�>��K?S�?��=�a��/��WHf��-)?�]<?LNM?��?Z�=�۾��9���J�YH���>�Z�<���X���#����:����:��s>[0���ߠ�QUb>���wt޾�n��J����IM=?�fZV=@�%�վ5�n��=f%
>]����� ����֪�j1J?@�j=�w��7bU��q��j�>���>?߮>��:�_�v�Ň@�߯��h7�=ص�>��:>�e��:��4G��7�Uؗ>_L?�8;?_v�?޻@��Sx�u�+��<�����������R?V�>�z?ڝK> G=��޾S8�v�C�J�'�>��> k�}E�0���魾!}���>��?x�>�	?+Ō?�4?��n?�5?-8?��>�0����׼&?ʃ?�q=I�˽��S���7��F���>44+?+wC�C��>E�?�?Ǟ'?
Q?1F?�Y
>{��8�@����>S�>.�W��#����_>unK?��>ciV?؂?�B><G4�����դ�|�=��#>H4?,�"?
?H.�>���>�K����=s�>$�b?to�?W�p?�-�=�A?�C4>�P�>��=�B�>���>p7?��O?rs?�AI?���>F=�<C0��9ӱ�5z�.�~��Z;��]<d�m=��׼�a� �3��C�<�5<���[�l�ܼrG��s�N3H< ��>��s>	9���0>��ž���
t@>����ܛ�X���GI;���=j�>q?���>��$�q��=�1�>���>�H�1(?0?�?�)q;�b���ھ��N��@�>a�A?�4�=�m�h�����u��d=��m?.<^?�cY�D�����d?�m?8��(��*����S�� �C�/?�y2?��U���>Õ�?�L?�?��'�=�wM���i�6��l��=�*�>.��F؊�X��>��I?��M>I�=�Y�=-�~��@W��f���� ?
ҋ?׆�?���?U6>�(���i�[=���@���"�?���>$̟�8�
?��<go۾�����c��_�O����z�鍃�f��=�ڃ�����!�=��2?��}?��c? j?k
���!�o�{�X�Ё�s��C�-�~8���>�����I����J��/'���e�>7�>�~o��dE�t�?�� ?��߼?H���-@�r&��?>���� ����C='����3=�c=��^�,�� �q� ?\:�>��>�M<?E�W�w�5�þ9�W�3�J��NG�=�ُ>�Hr>>��>�we�i�(��'�/B��E�xl��!hw>�c?�E?�Sq?��ݽ��/�L��TM�$0.���ƾ��T>�y�=y{�>@�V�p�)���D�8�o�T���R����	� �=��8?�l�>n��>d��?�?��;+���K��sT.��D=~��>��b?`�>Ip�>-�׽�3 �EW�>�l?�ѥ>�n�>��d���	��xn�����܏>K+(=i�?�K�=�u���L�#c��{����sj�#�>�uh?�*������jV>Q?���= �ƽu9�>X�pw����m�N��=��?�3�=YEy>c��oP꾸���z1��I)??x?���n�*����>&�!?�b�>��>�?���>�¾6��:##?�H_?ӺJ?��A?���>D�=a鶽>�ɽ��'�K�/=V��>�.[>��j=��=�� �\�����C=���=;�Ӽ'���r<aw���{H<گ�<~4>m�ڿ�K�STվ$�g�X�s-��>H��rY��ֲ��*��yΘ�C_p��
����pQ��|`��-����k�g��?��?�����"���a��љ�����]�>�
�X�[�G����	��放�x��F��o#��6O���g�}[`�P�'?�����ǿ𰡿�:ܾ5! ?�A ?6�y?��9�"���8�� >C�<,-����뾮���	�ο9�����^?���>��/��j��>ޥ�>�X>�Hq>����螾X1�<��?6�-?��>Ďr�/�ɿb���¤<���?0�@}A?��(����+V=���>�	?N�?>BS1��I�����jT�>*<�?���?�zM=v�W�~�	�]e?�<��F���ݻ�=58�=�A=���<�J>sU�>0���SA��?ܽJ�4>څ>�"����^�w�<��]>��ս�8��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�����nÿ�o�3> �;�<	e=E�#<J}��V��`��X܉��f��<��jζ=��">�c>�Ԁ>�>ˣ3>��T?.�h?�]�>I�>8�j�-c��p��t2��!��qN������}���3��_d���پћ��:���0Ӛ�N =���=�6R����,� �{�b�|�F�u�.?st$>:�ʾF�M��-<�pʾx���턼祽�/̾�1�t!n�
͟?��A?�����V���Z]�|�����W?�O����T謾���=������=�$�>���=���?!3�Y}S�k0?�g?j�����S*>[2�b=G�+?8r?f=<�g�>	%?/+��q位:[>_�2>��>܈�>1�	>�d���o۽�?I�T?���7����>b���z��A\=7�>�H5�P�伌\>�ؒ<M܌�!�K�x*�����<��`?XL>*�?�0(���׾n�9�ض�=H:�?S�?�h�>;hm?vv4?��<���[�������=��m?��s?��=�=����ዾ$#%?IE?�6�=�|T������?*�@D���?�NZ?g9+?�����)��c�����uP:?%�v?�r^��s��F����V�T:�>u\�>F��>��9��l�>W�>?�#�<G������Y4��?G�@b��?<<�N��=m:?�Z�>�O�\?ƾ+y�������q="�>
���ncv����oN,��8?ϟ�?��>���T����>������?9�?�Ϝ�^ا=���\q�Ս��h���@��h"���u����1�� ̾���9':�����E�>\@��U����>y^��/~׿�п�i�+�ྕ����?u>N@��犬��Lq�9~�iV��4�.O����>�E
>����Lb��b\}��Z;�$�\�ڵ�>q�����>�rM�}'������J-q�i�>@#�>��>�˗��	�����?�c��Bjο:�������U?�Z�?���?�4"?�6�<f�^�KXn��zȻ��D?�r?�1X?GI+�A�I��5*�0bm?d��k�e�VM4��AQ�Ո�=5
(?%�>��9�='�>��>��>"-3�"���zS��};־�٨?{��?����?�C�?	�+?���]W������G��4��R(?�A=*ʾK�2��h)�����{�>7�"?�u?����]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�+�>��?���=��>�U�=���c5��0$>��=��Z��?n�L?~��>u�=E8�.s/��2G�5�Q�)���C�WF�>�a?M?�8d>l��a�%�����Ƚ�5�x3��R@����ܽ�z5>��=>i>�:F��Ҿ��?Mp�9�ؿ j��"p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>B�Խ����\�����7>1�B?Y��D��u�o�y�>���?
�@�ծ?ji��	?v��O���^~����M7�T��=;�7?F+��z>���>^�=dlv�輪� �s����>�B�?�y�?��>��l?��o�n�B��;1==�>.�k?�w?�Na�!���B>'�?ç������J��f?�
@r@\�^?�颿O�ؿe���Q��[Ͼ]n=퀼=-�e>!<�[�v=���<}�=:����>��>��b>Ȣ�>�nw>��7>�4&>&����䨛��L��'�=�&d�i
	��8u��5��A`����?��x��ɷ½ZL���%���b.�uX��qO����=��U?@	R?>p?�� ?e�x�y�>���M=�d#��τ=x@�>�m2?F�L?��*?"�=�����d�Tb���E���·�ɇ�>�yI>�{�>A�>k2�>dh9F�I>�1?>A|�>�� >�7'=[�ۺz�=F�N>�H�>���>�y�>�C<>��>Fϴ��1��j�h��
w�s̽1�?���S�J��1���9��Ӧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW? �>!��s�T�4:>8����j�5`>�+ �}l���)��%Q>wl?[�f>Zu>%�3��d8���P��p���y|>:36?�߶�E9��u�K�H��^ݾ.MM>;Ⱦ>ɤC�$j�����F��ki�%�{=w:?��?m��T갾B�u��C��YER>WG\>�s=f\�=�\M>�_c�I�ƽ�H�Wl.=��=��^>h\?��+>Í=���>Ō����P�u��>��B>_�,>�@?j%?��e����ȃ��h.�ygv>�U�>�R�>��>�K�bv�=P��>�b>�|�(т����@��W>��~�]�_��kt��y=�K��n>�=���=�L �t�<�l�%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿqh�>`x�{Z�������u�g�#=&��>�8H?�V��l�O�5>��v
?�? _�ߩ����ȿ(|v���>G�?���?D�m��A���@�h��>��?�gY?�oi>�g۾`Z���>λ@?�R?��>�9���'�Y�?�޶?կ�?�L>	*�?�q?Rx�>��{���-��ٳ�����Jzh=!�׻t�>E�=�S����E�A���ĉ��ml��l��}c>� =���>������"��=�J���B��φl��Y�>s�p>�P>x��>0 ?�D�>�>��= Y��dp��.��?+H?QϚ?FO:��I����?S�>�?1��8?�.?�.>��ν7lG?"n�?ת�?7�?9/ ?g������IϿ�6־�� �%�a>.�>ʇ.?�fo�o��>CԳ����"+�>f$>�<Ъ��o��8�K>�֎>p��>SϤ>f�=B%!?��#?g�`>
�>��C��[��~G�|8�>y��>A	?��y?V�?.�����1�C�������]�`�:K^>�5v?l�?o�>��z(���JR��`h��n��~?kd?��߽�?1��?��:?>?��g>[���ݾ![ܽ�"�>��!?��*�A��M&�F�u~?]P?)��>�7�� �սnFּ����� ?�(\?nA&?��%,a�0�¾n5�<��"���U����;�{D���>ˎ>]������=�>zװ=hPm��F6�B�f<�k�=��>I�=�.7��u���,?�F�ċ���t�=Rs�� E��
>#:P>�����^?�=���z��n�� S���\Y��܌?��?e��?4>��i��5=?.�?�?�M�>}���>߾�]��x��y���� >G�>D]��8�\1���婿rC���ʽ�����Y?wƩ>\�?�`�>�5�=L��>�]��/��-�	�:+�)�`�]�(�#�3��I!�[$�w������w��	����Ke��>��=��>s��>�W�>Ϊs>Ƿ�>��:���>�R_>���>�4�>��>�C�>�v>�Pr<ۖ7�fKR?������'����ն���1B?RSd?�!�>[j���������h?+x�?�f�?�u>�h��B+�%w?>�>����y
?99=B�）<Y\����I�����B��>�vֽ�:��M�mhf��i
?$#?�Y����̾W�ֽ`�X�;7�=��?E�0?
�*�6�6�J�l�կ6��p�����5�����ʾ�� �%�h�c��
ތ��B���0�`�>�6?8g�?�� �|�žC�;X�f��+1�
�t>#�E>&> M�>_�k<%�#�~0B�Gg��jx<�����r�>m�|?C��>&�I?R<?XrP?jL?��>�b�>�3��fp�>��;m��>���>V�9?��-?Z50?}x?�u+?0c>"������ܑؾ�?��?tF?�?��?�څ�`ýNL��|�f��y��\��:X�=�|�<`�׽|u�L
U=�T>\?�e�å8�������j>x�7?TF�>���>n2���O��p��<���>�
?�,�>� �v�r��}��p�>O��?/1�}�=�\)>��=�$����溸��=�d¼��=]邼^�9�v�<|'�=Hٔ=��n��h�����:L'v;�7�<��
?�#
?9�4>`=>�1����
�F��%�'>�a>��t>XLK>�ھ񾄿����{m��:}>Q��?�z�?���=�<>/"�=y?�־}��&=ɾqC�=|� ?ĩ.?��M?ż�?H?GR$?Ղ>���ꐿ:���։\�){?� ,?]��>�����ʾ�憎	�3���?a\?b:a�����8)���¾��Խ��>uZ/��/~����D�脻���/�����?R��?EA���6�u�S����W���C?d�>�X�>��>��)���g�$��9;>���>E	R? $�>��O?.<{?��[?�hT>C�8�`1���ә��53���!>6@?��?�?�y?�t�>��>��)�T��T�����ႾE	W=	Z>e��>d(�>��>z��=��ǽc[����>�}b�=��b>+��>���>��>t�w>�A�<�>H?w�>*�������]�������(2��u?�7�?�~+?2=3��߫E������K�>�
�?���?��*?8P�y��=|��Mٸ��u�%9�>�!�>L8�>��=�\=��>���>CJ�>P��!��hZ7���S�X?/�F?㍿=��ſ-�r���l�bN��t�<�N���I�-D��F�H���=�ϔ�=���楾_�N��^����������;��F���&�>�ˌ=��=��=�a����2��H�;Rx0=�T<�@S=H2K�y�;�����ȻM�w�ԟ���r<�J�<��;R�˾��}?�;I?Ε+?z�C?Z�y>�;>��3�[��>�����@?�V>;�P�㈼��;�
���5 ���ؾx׾4�c�;ʟ�pI>�^I��>�83>9H�=FJ�<��=�s=%=��Q��=R%�=�O�=�h�=���=&�>"U>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>)�7>$'>��R��1�]�\���b�J�Z�,�!??J;�O̾Y6�>5�=o/߾��ƾ\T.= u6>��a=tV��Q\�$ܙ=��z���;=.�k=�׉>��C>��=�6����=��I=���=��O>������7��,�k�3=Ҹ�=�b>�&>}��>��?�a0?�Xd?D6�>�n��Ͼ?��yI�>�=(F�>j��=sB>⏸> �7?.�D?O�K?��>:��=�	�>��>E�,���m��m�o̧�̑�<���?�Ά?	Ӹ>8�Q<��A�b��Xg>�z/Ž�v?mS1?�k?�>,����0̿�M㾾 ���=Ƶ{>iU?�&��*��=�=ޮ�=˟��{���>�G?7�?���>�'>M�	>��k>�i���h�=}3�=8x"=��y=��G=���=�B�=�!�=*E �Cz�H�����'�s=�R�����c�<}�<�T>���>wJ>RN�>��z<��ɾ��>�y����=�;�=��Ѿ�@A��ms��q��i�<�T�t�}b>��c>`a�b䘿�S?_ �>�H>�a�?��s?@UU>��Z�𜺾0ˍ���W���T~�� >m��$�!��P�f�R�x���>�>蓠>��W>�D>�+�J�8�5�
<�־O �7�>�p��2:ڽ}����fm�в��Q?��x�Z�z�=FEN?�ˏ��
>��v?�@E?&r�?��>+z�<����Do>�~���������������f?�?�)�>�:�*F�^{M��U��Y�>vgĺ�`�s⚿�?
�}��+�+�3v�>~h�j6�w�/�,ed���8���T��Gw>��Z?���?W螾���d*^�Z3���>iX?��D?U?���>��;?�͢�����	���A���-�?��?wa�?B�<d!�=wýX�>*?�_�?���?lbt?�JC�A��>O�; � >,���#�=o>��= ��=d�?e�	?��	?is$	��}���^a�y��<6H�=�<�>;.�>�)u>9l�=C.^=F��=g�^>�ٞ>ͨ�>u9b>�l�>�-�>�8���n��<�Q?1P�=�i>�q0?Q.�>�T����=��>�����<�_�����ƽE�!�CNa=Ui->(>/H��O��>��׿~��?�H>��ž�A7?�־cų����=��=��6�>��y>L��>��>Ѧ>�=K�>?�>u�Ҿ�>M��@<!��&C�_IR���Ѿ�az>"Ԝ��&�^�����=�I��v���z��j�W;���<�~Ҿ<<7�?3��k�k���)�0���m?8G�>R	6?�挾휉�Xu>ï�>~�>�8������wč������?��?Ec>��>�W?؞?M�1���2��tZ���u�*%A�Ye��`��ߍ�������
�z��h�_?>�x?��A?R$�<.Hz>6��?*�%��ˏ��>z/��.;���<=w�>|>����`��Ӿ{�þrE��F>�o?7�?X?�0V�xm�á�=Eb3?��)? �q?�8?�eC?p(�!?S>A>L�?�
 ?�*?g|-?��?�UY>�>��ɻi��<�Q��f��G浽e}⽙rS�;��<�Au=����vi$=x=���Y"����:S��<m����<��=ѿ=�?>p��>��]?4M�>z��>��7?����w8��Ʈ��+/?[�9=��������ʢ�����>S�j?w �?�dZ?�ad>��A��C��>�X�>�q&>�\>e�>�z��E� �=�L>�Y>�ȥ=(XM��΁���	�f������<D&>8��>�/|>H����'>�Q=z��d>9�Q��Ⱥ���S���G���1��v��P�>��K?��?��=�U�����Kf�)/)?�_<?�MM?��?O�=��۾��9���J��=���>�ѩ<�	�Ϳ���"����:�OG�:�s>�9���Ӡ�k_b>B���v޾�n�VJ�u�羒!M=7|��sV=�A�վ�*�B��=�%
>h����� �����ת��.J?��j=�z��,hU�"n���>���>hҮ>��:�P�v��@�����$�=���>�;>J=��:�}G��6���>�*Q?NL?���?�䚾'�s�3&��^��Cz;�uB�b�?�I�>�H?�>���ۈɾe��N��(�Rh�>`ǵ>]�3��l[����Er�z|F�q�[>�_?Փ[>�2?<_W?��?��y?��>?��!?Iڑ>�紽�6��B&?<��?�ׄ=��Խ��T�� 9��F����>�)?x�B�˻�>��?��?��&?��Q?��?R�>Ѯ �E@���>�Y�>��W��a����_>ŬJ?���>+:Y?�Ӄ?��=>˄5��ꢾvҩ��^�=B>��2?"5#?(�?F��>�>?�о�+a;�6]>.�x?/ʍ?=`y?�x>�]?�>�7�>�	�;<r�>l?Pg?OO??C*�?z�>?2��>�<w�r�ǽs�ͽ&��:�M�<�c:���)>��s��V	�h��<�6v��<���J�=V�j=�o�����<�̧<�c�>%�s>���)�0>{�ľ,W��P�@>|���H���ڊ�r�:��=��>��?1��>X#�P��=b��>�P�>
��X2(?��?-?��';ڛb���ھQ�K��
�>6�A?Jr�=��l�������u�1�g=��m?Z�^?��W�����xj?��[?}��I-�����ľd����*?�?'�k���>�2�?��q?��>ћ?��PG��А�fN����Zs>ϯ�>���u}�/�>:oD?B�p>l.3=^ �<�#\�w�Q�H�ž	�?��?���?\.�?<:S>��u��J�����Ñ�O'g?�V�>�ؤ��#?�j�;d�;�ɛ�Rp�����RP��F8�����F������@E��s�����=4?:�m?��n?��`?5
�gHe���\���w��R�a.�����SA�v�=���;�7(o����RI�x�ެi=3j�MpE����?Cf ?<:��%�>�Mp��羼~����=Bd۾�"��`�������+���^=Sz���r�e<��4�)?8�>諯>B?�;o�CH���8���$���Ӥ�=)h�>a�>��>4�=��k�3;���6¾E_ٽ�Z'�HCv>�c?_K?)�n?�� ��#1��{��O�!��(+������/B>�I>sʉ>2pW��u���%�zT>�h s�����ɐ���	�Pۀ=��2?�+�>��>K�?O�?fZ	�K˯��mx���1�T�x<��>�h?$��>���>�#Ͻ�� �m�>�Y?��>�h�>Mdྫྷ� �<�Z��	>�>Z>^��ڇ�>�	*>�}����Y�RԐ�˛���S�ĳ�>�Bw?QQľ�kX�]��>�?g?"�&��V=��?m@߽)���M���we�[0A>�]'?|ȱ<͎�>����D�>�����x��?�J�>�����
A�Ӹ�>�b5?�?���>ߣq?���>Řľ��:�-?H7b?HM?�F?� ?��=Fe������)�<�z0I=��7>,:>Ó=vs�=�ec�ɮ�����4ȇ<Z��=�v���0�<�nW<�uy<�3=F>,�ڿL�P%P���	�+���?���ݾ�;����ؾӥ9��L����Ӿ�[#�:�>��c�=�Q8��f�G����ݧ��B�?D��?j��W��]���8���Pj��?�LϾ�j<8zy�J���4}޾NR�7,վ]nG��_l���`��aN�?�'?���x�ǿ������ܾ��?��?�y?���<h"�|y8��� >�F�<D	���뾑�����οs֙�W�^?�b�>�~� ������>m�>'zX>�p>�X���➾)f�<~S?"o-?0W�>r���ɿ�u���<j��?��@�{A?��(�<��c�U=��>��	?��?>�N1�H������T�>�;�?���?�M==�W���	��e?�<3�F�@,޻}�=�:�=,F=����J>GS�>w���OA��C֮ܽ4>J؅>�"�5����^�?z�<�]>��սQ.��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��=D��yKǿ5C��R���9<~�(�"�ݽ�gc�Y.�����#?j��J�v�	�� #=W�a>�ȃ>�>��L>�>e�Z?y�q?׋�>l>8�Y�����[����;YM���*D�����F	������s
���߾h��T�:k�3�ξf�<���=a,R�c���c� ��b��F�N�.?�e$>Շʾ>�M���)<'�ʾ
��|����N��J7̾h1�` n��П?t�A?��DW�������~}��$}W?eF�g��Y8�����=������=Rۜ>�u�=�⾦�2��CS���0?� ?unž�ˏ�$�+>{`��F�<~.(?�?A��;n��>� +?c� �E^⽗n>0F>>�>���>�j>rU���� ?�EV?�J�]d��6��>K��$p��&�<1��=�dC�:8���J>]�<a���[[ɼ/(���̶<�`?��Y>�1;���2�p;}����;6y?m�?M��>:�M?�l0?�C���y��G����ؗټ�'`?�P[?�>���FHܾڲ�x9?lY?�i >o&���ⶾ�9�=*�tm?˘F?׎?�����x�|-������Q�D?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?w�;<��U��=�;?l\�> �O��>ƾ�z������1�q=�"�>���ev����R,�f�8?ݠ�?���>���������=���Io�?���?YH��Ͻl<&r�`k�צ �Ϭg<(�=ɚ"�!>��է8�^ƾ�
�Yj���j��-��>cU@�������>[C<����]hϿ�4��[�̾+Qp��?�K�>�½E���j�m�t���G��^G�������>� >X���C��������qB�g��v8�>P^�U��>��(�����ͫ�o$3�q܌>C<�>w~m>~yz��+��b�?5-����Ͽ^O������Z?�>�?��z?�G,?qO���琾�?�]�N�)~=?0/c?	S?�K�`W��:���m?e$��yg���A�#G�]M�=%�?p~�>D���a|=�k=@��>�=;�6��x���i������B�?�w�?������>`͟?f0?�쾴y���T��T0�&V����+?/�\��<�����o/�� �����>.�5?8Rܽy:�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�۵>��?*�>�"?aF�=�y���<�6>i��=#Cǽ��>eH?���>V��=W.R��17��H��cJ�wr�E��c�>� ]?�oJ?��k>)�ֽƝ�:��$��曽޾,���k��y.��ʒ��Ľ�>��->82>#g�������?Hp�8�ؿj��9p'��54?#��>�?��{�t�����;_?9z�>�6��+���%���B�`��?�G�?5�?��׾�Q̼�>H�>�I�>S�Խ����b�����7>�B?T��D��m�o�d�>���?�@�ծ?Xi��	?���P��Va~����7�c��=��7?�0� �z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B�{�1=7M�>Μk?�s?�Qo���h�B>��?!������L��f?�
@u@a�^?*�hֿ����ZN��V���-��=���=�2>��ٽ_�=��7=��8�-=�����=l�>�d>4q>*(O>la;>��)>���J�!�	r��M���G�C�������Z�C���Wv�Fz��3�� ���j?���3ý�x���Q�2&�}?`�9�=$V?��;?]4m?!F?��� >'��ͫO>[S��%{<��>G"?�B?])?F0�>?q��|y��o���˾����<ض>T�=)��>A?1�>ݙ����=̉�>#��>���<�D>Gt�(�S=���>7|?�(�>�C<>��>Bϴ��1��p�h�w��̽/�?t���C�J��1���9��ߦ��vh�=Ab.?�{>���?п^����2H?&����)��+���>��0?�cW?�>����T��9>��˦j�3`>�+ �~l���)��%Q>yl?��f>u>ƛ3�e8���P�o|���h|>M36?�綾WE9���u�߱H��bݾ(HM>]ž>R�C��k��������wi�R�{=Ux:?��?34��o᰾Ӯu��C��PR>Q9\>xR=�d�=�VM>*^c��ƽyH��f.=���=>�^>M]?�+>:ō=��>�e���CP��t�>�B>�8,>U@?�%?iz������.�E�v>F3�>�$�>z�>�J�,�=8m�>��a>������(���@��`W>M�D`�9�u�j�x=���39�=F��='� �f�<��'=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>���U��l��'�u���!=��>�AH?.���cN���=��b
?��?�򾲙����ȿ�pv���>T��?��?�m�sD���@�Pr�>���?;[Y?$i>^۾}�Z��"�>3�@?��Q?��>gB�ѧ'�l�?sܶ?!��?b`F>`�?�qt?Sf ?G�ѽ��'�����J��ZGP=U���_g>�>����� E����G����j�a�0��>�=��>yh��q��$p>l�۳�M��>��>}�>�cG>���>�^?y��>˒>��=�-F����ڜ�iHS?���?g�]��V�m&��A��n��(�ս�p8?)��=�$A�=�"?��j?/}p?y��?��?R_��䭿�#����پ��=<4\>���>�%?��ڽx�>�m��w����<~��<��=>혴�0j�����>4��>�ǻ>�'I=z�>� ?��%?t@\>(�>��D�O���A�6��>y�>��?iyx?-c?�ﱾՓ0�Ã���g��m7Z��R>�t??K ?��>|���F��Ҍ��y��� ���{?zZi?ɸ�"�?��?v�??�/H?��>�ؽ�Ӿ��ZG>��!?'���A��S&�2����?^Q?2��>�?���ս�iּ���pp��'?)\?�B&?���H&a�?�¾;1�<#��bU�[��;��D���>�>gi���i�=k>|��=�Dm��A6��f<Iw�=	��>��=�+7�����=,?ΦG�%ڃ�Z͘=S�r��xD�N�>�HL>���ߩ^?d�=�Q�{�����x��U����?N��?�k�?�ʹ�q�h�"=?3�?�?@(�>mG��9w޾ܗྔew��}x��{��>���>��l�=����9���F����ŽK�'��!�>�|�>ʐ?�U�>�d>�.�>���KV5�r0�GD"���H��m3��gE��0+���!�6ʹ�9� �ܨG=�WԾ���K�>`PɽQ�>`�?��>I��=	�>)Ɏ���y>�=,>G>F~�>��">��>
��=�"��s��KR?����7�'�·辺���G3B?�qd?Y1�>ei� ��������?���?<s�?�<v>�~h��,+�|n?�>�>[��Rq
?U:=8��=�<�U��w���3��3�
��>�F׽� :��M�nf�\j
?�/?����̾';׽�O�����<�}�?�x(?�*/��,E�@fo�g5�u�p�;[	�����2\۾��3��q����
n�V�v�_�⾐��<�O?�9�?gg$��Z����ܾ���j@�u��>��?3Ҳ>: ?B6/>�o���V(�1g_��+�~����>/[�?��I>rM;?A?.t<?�BZ?qA�>M��>����_T?ݑj�C��>���>�`$?!F9?��-?�-?�?��=>e�����6���?�n?�*,?<�?�	?і�����Nvt>���=�ϾmL.��V>����'΢��!>��>�Ja>=�?�����8�;���5sg>=G6?���>���>�ێ�������<���>C+	?k;�>�� ��mr����7S�>ς?q���u=У)>�V�=�8��L���=򸾼��=�����7��}9<��=]��=/�4��*��'�ѺN�@;��<�d?6�?3�>7,�>�������g���=��>>�	>��=Qݾ�]���'���t�}V>I��??�?M>1 >��Y>L���1vþ����ľ�D=���?�0?�8I?���?q�4?@�+?�U>,{�H���3w���U��=z ?��,?;��>���;������3���?rG?��_�����)�?b������&>k�/���~�bS��E|@����;8���h��Ĝ�?ۗ�?�%�\6�7)�⊘�m��B?� �>���>���>-�(��Zg�%���g@>2�>�R?�(�>T�O?�,{?�[?�nT>{�8��/���ҙ�.(1�+�!>'@?8��?��?gy?9��>V>��)�Y1ྑR���6��*��΂��W=�Z>I��>�(�>0�>��=	jȽM�����>��&�=�Zb>���>+��>]��>�zw>�`�<��G?���>�k������⤾����ă<�3�u?"��?��+?6=�x���E��;��.K�>�e�?�?�7*?��S���=Y=׼d춾�r�4�>��>M-�>��=edF=�/>J��>��>�6�BX�m8��VM���?�F?Z��=��ſ�q��zo�3�����g<ƴ��A�c��v����[�=
�=.�����6;��y\��������嵾�\����{�R��>D�=s�=E��=P�<�ϼZ��<4�J=?F�<#1=�in���n<T9���û�	��A�����[<AN=� ���˾�}?�;I?��+?g�C?%�y>h;>)�3���>�����@?hV>ŞP������;�x���� ��C�ؾ�w׾+�c��ɟ��H>X`I�F�>U83>�G�=�H�<��=�s=#=��Q��=F$�=;O�=�g�=��=��>GU>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>۷9>�L>b�R�Q�1�r�^���c���Z���!?L�:��j˾��>�Z�=H�߾<jǾ��*=�i4>�\=[����[��~�=�Rw�E�5=;�f=�u�>�D>7V�=J����-�=�w@=p��=r�P>DZ���3��5��D,=���=(jd>'6(>:��>c�?�a0?lXd?�6�>-n��Ͼ�?���I�>��='F�>���=~rB>8��>Q�7?��D?��K?���>���=7	�>U�>5�,��m�m�Ņ���<���?�Ά?_Ҹ>�Q<��A���ug>��0Ž�v?eS1?�k?��>�1����9^���!�͗��
(��~��= *��[a��C4���:��~���>�>���>]��>�dJ>]��=4>���>3�=��"��"0>��0��%ν`Ѝ�z�=�9��mF�<��=���<���g4"�\�?�hY9=��-<�h�T��+�=�>��|>w=�>�R=�p���B>��}��\�"�=����/-�9p����.:/��&��gm>)1�>՞�=Q�����>H�q>,?d>�s�?[}?7O>Q^�޽Ӿ@8��ر&�G�V���g�ޞ�=G��<�#�]��Rf�=L�����>8`�>��>(	>>|@(���?�d��<�¾�I8�g�>4L�|)�+r��Dv�IV���͟��R�4�=��^?��ޝ�=���?	T?7�?���>�M�^�4h=����4��yp�$z��հ��&?A�?١�>�D
��'.�Z2��mn��X��>��,��|[� ���:��m>��侀f�>�x%�=��!]1�FL���|�K�D�H剾��>�0?m��?�%i�_㎿QQ��s��E����?��G?�� ?P?5�>��p=�T�^���8Ի�yZ?m�?>K�?��d>�&���ҝ�9�a>���>�p�?��?[��?;9��O��>�?�j�>�'þUí>�?^�ռ��S=GQ�?���>Q��>Fǽ��+���A�����P�'�,=6m�=�@�>KiP=0B^>���<<��=��>�ӷ=si>Iz=>#T�>�|>��>$����d��.4?o�=sX�>��7?]��>~[�<S�)�҅��M9C��O�󾛾��:�S��͑�<����\=��2����>%dſ}+�?�}Q>�����?5׾�r���94>H�>-���%'�>�8A>=\z>w�|>��> �>���>��=ãǾ��>z�
��!�эF��U�U�Ӿh��>#ڜ������+����W�:����w��hh�����Z]6��3�<�E�?�0��{No���+�:��n�?}�>�a0?/t�� ��/��=���><(~>���Hǔ��z����߾�W�?��?��c>�f�>� X?ð?O2�b~2��Z�Lu�IhA�('e� a�R�������6�
�)�ýk_?_x?�A?}�<��{>�ڀ?�A&�|5����>$f/�[�;���>=���>�����^�4�Ӿ}�¾8T���D>�o?Fу?�i?��S���n�<�%>�:?�1?HWt?/$2?��;?A_�R�$?� 5>�t?VQ?f�5?�/?o�
?��1>U��=���6'=����DL��ҽ�>ͽ�n�J$7="}=��Ӂ<!=ϡ<3X鼹�Ҽ3�;5���5�<��7=}��=��=2��>ܛ]?^?�>A��>s�7?Ȫ�3e8��ٮ�U1/?�8:=[����"��(â�����>�j?���?XZ?�<d>��A�)0C��>i\�>��&>_\>�j�>?I�d�E�R�=Z>�>���=f�L��偾\�	��R���N�<�->���>��>���L�U>���ѧ��_�2>>"S�>�w�xۋ��VG� ���GK�r��>��Y?�4?���<w3��Zܽ��l�i?�F?�OP?�s?�j>���$$)��9�Cā�Y�>���KP�|���Bj��4K4�m�����>­��ڠ��Wb>P��#r޾��n��J����\M=N��O�V=����վ�8����=�
>���g� �����Ԫ�3J?Иj=�}��OjU��q��,�>Ø>�߮>H�:�I�v��@�q���g$�=���>'�:>�/��^ ﾔ{G�T5�<��>b{I?�I?�Ƙ?2"s��p���B��@�61����;�Z(?b�r>�2�>fZ >��~�B������O�o{C�;,�>���>Qp"��q�����N���0 �e�>��&?��5>��?�`?��?���?"�?�?s�?>�q��}��t +?V��?����彠(^��95���P��>9�-?j�jo�>4r'?u>*?ܣ ?Y�T?�?�sr=fW��Q��a�>���>A�S�E���ӽ�>�H?�>N�Q?�V�?�>�T7�S!V��4��,�=U�t>V�@?g�?�}�>�2�>jC�>tˡ��D�=5�>$c?�(�?��o?��=?[�1>��>��=.��>�^�>f�?/HO?o�s?9�J?i`�>a
�<��������Ws���N����;UM<�4x=7��	�t� ���<��;a���O#�������D�PW���b�;bu�>݊x>n6��ìl>��þ�k�WZ'>���ܨ�������8���=q>1 �>4��>?F=���=�b�>�M�>����c$?b��>3 ?���<�7h�u�ʾ�O��ԭ>\jE?�(>��d��W����w��P=�]k?IZa?,������|e?)Ie?z
�ȴ�t�¾�֨�(u�J�V?�?��C�
��>�{{?��r?��?c:J���=�Cޝ��>S������>���>Tp6��L����r>Ox-?�PY>�p>��Z>e��`l�U`�=�9?mBa?�\�?�٣?�"=tV��t Ϳ8r޾~芿��t?���>������?Y�����;E����$���(Ҿ�|���᰾�#��x����9���꺱���=�?�x?8�Z?�qd?�:�dn\�M�a�;�y���m���= ��aE�6H� �D�!�q��s�dp�-=�X|�=>�y�@�y
�?�#?s>,��*�>���UW�~Ҿ��C>U ����A��=����Z)=�L1=o,T��V*�����c"?U�>kF�>�N>?�\�'L>�i�1��5�����1>KJ�>d�>�F�>�q�R�>�M,	���ƾ�Nz�2�ʽ��v>/5c?�9K?T�o?8��*)0�;q��7�!��:�*��c%B>'	>��>��Y�H���y&�ϒ>�,Jr�9������f�	��z=�v3?uс>�m�>�,�?��?m	����Ju�}1�K�<��>}h?gP�>�>�o׽'@!�p��>7	[?I�>	�>�W�����Ev���_��+*>Pƚ=���>OC�<G��D>�ḣ�S9��P�Z�8&�>�oj?����t�W���=��p?2��<�p�h��>�wL����p̎�����r�->��?�Iw��cw>h��� �FJ��wc���:)?re?������*� ^>�)"?�_�>hX�>�5�?���>��þ^�:��?��^?JJ?NtA?�>L�=�ᲽnȽa�&�o_/=�R�>5[>;�n=��=�
���\�U)�nB=�޹=�qѼgٹ���<c���AN<�|�<��3>4Կ�J����������;狾�mɼ���[�������7��Y�1������;<�B������c���eb�a��?���?�`����y����A��-��V;�>���jߔ=Ь���'��K��rr���gԾܶ;�΄Q�K�c�׀U���'?b�����ǿư���<ܾS  ?�A ?O�y?��Ν"�?�8�ߩ >0�<�=��E��Z�����ο����&�^?���>L�0����>���>��X>�Gq>����枾��<��?��-?c��>��r���ɿ����{ۤ<���?�@�|A?n�(�����&V=���>��	?=�?>V1��I�0���uQ�>z:�?'��?�aM=��W���	��}e?�<��F���ݻ��=�;�=`=���=�J>^S�>��tUA�D?ܽe�4>�څ>*u"����3�^�:t�<ǋ]>��սA=��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�}��=[��>c�>,������O��I��U��=�-��ż�� $�*�$=ʬ�+�=�	.=����ػ%�½ÞN���'�"*>��>�Zt>y�>���>��=+�@?�#{?iC�>'�=`�Ƚa_k�YT-�6㏽��[���h��J����0�������� �31��⩾������q��=�p�=/7R�˗��k� �b�b���F��.?�v$>��ʾ��M�A�-<toʾྪ��ᄼKॽF.̾L�1��!n� ͟?��A?������V�o��-K�����d�W?�I�W��M묾Y��=W�����=�%�>I��=b�� 3�4}S�"%4?K�?j2ǾQ����q�=b��R�<�b/? ��>%<=>�>yU?h�9�d��d�0>�"+>6��><&�>y{P>vd��Db���m!?/�O?��ὭП����>�þ�=}�:�	=PS�=�A�; ��67>\��^���=�}i�D)=^X?_L�>��*�d��d���ӗ:��?=� y?߷?7��>��h?[�=?�1<�����S�k�	��)�=�BW?Цk?NH>,Xj��0˾�T��v�5?Mb?�iD><$g�����.��7��]?�	m?�?N�����z�������FD7?��v?nr^�Ss�������V�<�>_[�>���>�9�bl�>��>?:#��G��ﺿ��Y4��?\�@2��?�#<<C$�❎=�;??\�>��O��>ƾ|������?�q=�!�>!���dv����WS,�Ƈ8?f��?l��>u���.���n�=�ҕ��W�?��?O�����e<>���	l������Y�<���=��|�!�I��"�7��ƾ��
������ɿ�'Ɇ>�V@MQ�.Q�>�8��5�JϿZ��y}о��p���?7e�>�$ɽﳣ�!�j��^u�[�G��H������l�> �>�ԭ�3㏾���,#@�{J���>\�uښ>�A����Hң��T�6	�>�9�>ݼw>Gټ�����|�?"$���:ο�㞿�t�C�Y?=B�?�σ?��%?|�+;J���[���Ġ⼃�C?a�l?�QZ?V
A�3�B��мzxl?PЖ��I[�F�3�}�K�uo>X&?�}�>,&���=�0�=�V�>Q)�=�q9�V������� Ⱦ���?M<�?^^�s��>�?�?j�&?�j��S��D���
�0��˼�-?��A=� ���!��>��I����>�$4?2����n�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�-�>O�?�}�=}��>�'�=ī��q�1���">���=�.@�;�?�xM?�#�>~*�=�9�)/�$_F�-/R���L�C���>z�a?��L?Q�b>'���K1�� �ͽB�0���),@��#+�?.�I�4>��=>�>UrE�(3Ӿz�?�g�Бؿgg����'��!4?���>+?���Zt����r_?Y�>B<��'��o���@����?{D�?��?R�׾�̼��>���>'J�>P,ս+ꟽkl��c�7>��B?��1;����o���>!��?��@�Ԯ?s�h�	?���P��<a~����~7�}��=�7?p0�;�z>p��>��=�nv�û��J�s�O��>WB�?N{�?���>ٮl?$�o���B�,�1=�M�>��k?_s?�=o���r�B>�?��������K��f?��
@hu@��^?���Eѿ�ϝ�Z��������&>�H>��>J���b�;�-^�T�>>֗�<ؠ>3��>�4.>�eP>[�r>���>��>dy��%�k	��p�t��91��1��'��h�m�m�S�^����I3��1N���sT��ֽ�NϽ�e��@v �a,�2��=��^?Y�F?�h?��?�4���'>����:c>*rQ�.�2=y&�>\[F?WTm?`u=?	�Z>
���:bm�'Om����Z,����?�">��>q�?���>Y^X� m>8e�=���>g�3>e�߼)�ܽ�e˽�0>ޚ�>_8�>�'�>yI<>��>bϴ�1����h��w��/̽� �?|����J��0���0������i�=Gc.?��>��?п�����0H?9����(���+��>"�0?�aW?��>����T�I2>�����j��\>j ��sl�Ō)��Q>�m?~�f>Hu>&�3��e8���P�}��+n|>�66?涾9�X�u�}�H�jݾT+M>��>ED�wh�'�����ki��{=�s:?�?W����ٰ�Y�u�m>��XR>@\>v3=e��=�ZM> �c�k�ƽ3�G��/=���=(�^>�	?h�(>(�+=n-�>�����^��M�>�]>H�#>
�B?�?n!u�&e��������A��o>5f�>4��>�6>�J��G�=��>b�\>��%�#抽����@�َR>�&��8l�	�g�ք=9���^��=���=[u��K�d��=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�>	����������;x��0�<��>��H?�\�����t�:��n?�B?���l�����ǿK^v����>�[�? ��?hm�ҩ����@����>�N�?��X?��j>&�Ҿ�v`��l�>>?O?�>�Q����u'?��?c��?MW>��?�Mk?��?#[]��n"��;���Ռ�ĴV;��c�M�>�c�=䏽��AI�Kx��Eg���Bb�w��kO>_o=kϿ>.���!����=��������8�>���>�(�>/y�>�)?�z�>K9s>BEt<MaJ�W��yݚ�cJ?Sh�?8�9�~�3�Ym�>v���f�sD3?��r?}�+��[���@?���?o]w?M�?>�0?�p;����U����$þ����蒩>s<�>�?YNJ����>�s����ֽQ^�>O�=^�����Ⱦ��=�m�=��>��>���>+�>D� ?U!#?^F`>+��>�G������C�6��>S��>=?�?�N?c|�� 02�?��0f���XZ��C>Քt?�: ?%O�>ǅ������{���+k6�`�}��I�?��k?g[�@�?��?�;?��B?��^>!'���۾V.����}>�-"?���6�A�[b&�:��?8=?t��>����ͽ�Bټp��(����?�[?V�%?^M��E`�����[�<�|�*�L�$��;����1>�i>v���ֿ�=�2>��=�i��4�<�S<~��=�>J�=
3�0���T�.?u�<R�q�<�)=ϳw�t�I�a�m>��Y>�K��{�\?V�����h��������P��^��?�)�?��?=	=Ysk��h2?��?�'?9 �>����c����5\�������/�;�=���>�$��v�ݾt���a̢����Ջ���O��>���>�B?��>&�>�q�>=X��<�$N޾�=#��c��U*��GE���2���'�����ꁽ��=�i��Q���>����B�>� ?Nhd>�T�>��>M��=��>tE>{��>9��>I"D>\]B>x��=�+W�kЂ�6KR?����G�'��辍����?B?mZd??�>��i�D���R��ml?r{�?�l�?[v>Ոh��7+��z?L�>���dh
??�9=��
��R�<�[���������W���>J׽�:�M�&�f�m
?z.?������̾{׽�֏���=(�?7e,?�\?�w�o�K�b�Z/��v�I�6>�������_u�@}m�aQ���6��D�m���+�I�d=�ZP?	!�?�@"�#�Ⱦ��꾔Uo��R���E>�U�>_M�>þ>��=��6�o�=��{���.��о��>��u?}��>�gP?�|??�MM?��Z?���>�̭>�ž�?�"b��&�>��?�eC?��<?��6?fI#?� ?�(�=y��&�����Ͼ�%?� ?uE?l ?�{?k~%�\� ����)&��ݹ1�r�ν��K���u�TW���߁<�5�=�
3>	U?���0o8�����	�E>)�1?̃�>�>M8��N�h�M��<���>�C?��>p��u[n��p	���>�/�?`w�H =�'>Ƙ�=�*�:A,��c�=�ί�)��=�H��H�̆='�=V{=;8e�{:;@��<Ќ�<�"2=q!?�Y?��>���>�g����"��2��>��=�G�=�������"n��;Gk���>�S�?�^�?��=��=�Q>k���te��{������f3���?J�?��I?�C�?�`(?��?��C>vd���������c�gM'?�$,?ۈ�>���]�ʾr��3��?O_?N7a����7)�2�¾ սv�>�\/��(~�`��D������`�����?\��?��@�%�6��z�Ҽ���X���C?�>tl�>�>z�)�^�g�T#�&X;>��>^R?�#�>��O?4<{?�[?�iT>c�8��0���ә��3���!>�@?˱�?��?Sy?u�>��>ں)�K�4T��`��M�N߂�xW=�	Z>���>U)�>Z�>���=�Ƚ�U��\�>��_�=��b><��>��>y�>�w>I�<b�J?%?�>�GǾY��2+��Vx�����I�v?�;�?��/?(�=U��(�F�y� �^�>hϣ?��?�@)?�/"�\F�=��x�񮮾��m�!��>��>V�>�V�=F2]=%�>���>C��>�4����?�2���(���?MvH?6��=wkſ#Yr�\dp��*��c��<0cX�����(S��ħ=����X��ϱ���mW�����&폾ݣ���C��A^~�v�>de�=x��=A(�=4�<.��6B�<e�3=�Ć<^�<WKp�I<��!�����݌��b����<R�K=�7��F�˾.�}?�<I?k�+?��C? �y>�<>��3�?��>E����??#V>�P�j���b�;�I���;��V�ؾ[x׾8�c��ʟ�\K>]I�x�>�93>�F�=�D�<��=�s=?Ȏ=��Q�=� �=zL�=|f�=3��=8�>�S>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>BQ>[h�=�9S�`r2�� ��'�k�*�I���$?�P6����?��>�zW=(��[�;�<��1>��c=�����K�!ޛ=K�R�n[E=�I=�S�>�E>�֒=𫫽w)�=#h�<~�=/%j>�M�;�+g�{u��Hf=�5>4�}>AjB>i��>t�?_a0?nZd?�5�>�
n�GϾA���F�>��=F�>�څ=qB>댸>#�7?׳D?w�K?��>n��=�>.�>��,��m��k�fϧ����<C��?zΆ?Ը>n"R<A�A�ß��f>��6Ž#v?�S1?�j?��>9���k�п���U.�<>']'=���>�i~�]��=m�=B�&>�ռ0�=��>���>N�>��>�db>�8=��>���<���:965<4�C���d|�<pA>�qн�I>���8�ѽ�f�3��@]>l�H=��j=���(A"�bJ>3�>%�>#`�>�X߼���eO4>�Yо��@���>���a�4��{w�[���5�;�t���k>�	e>���=�/����>��>�p.>��?���?�]>����1�����%疾n��{6���>�
�F�.��u�)sA�"O����>Ò>��>ʀ�>~�*��$�1�<t���:��>����Y����1��0p�����͟��Jl�=��B?�����=l?��Z?��?jw�> �м�׾��">��N�;�=wa
��C�QL
��Q?S�'?��>�a
�"!M��j�!��� M>�ib�(.{�pH������4�=��Ҿ�!?�Cn�D�A�6��an���u>�f��m1�>�#S?�̪?�B��h���iZ�������=�	?V?��>%�>�ɯ>Y#�r���F`Y�W�=�q?yO�?�d�?�\�>�Y�=^h��Z��>)�?/��?���?Ws?�@��s�>�k�;� >ֽ���>�=}`>�L�=��=o�?@v
?��
?������	�L2�=���]�K#�<��=�=�>�>ڝq> :�=�(g=���=u \>���>̏>Ue>��>2�>aB����
�]�D?7�s=�K�>��=?�.�>��<ϑ�
�&=%���I�:!w�4�2&���8��=�<��d=�߇��%�>� ��]`�?Z�S>���"�?� �]��jǳ=l��=�Y=4S�>4�G>z�>a�>d��>�z>^ �>�d=�ξ�_>zg�2��S;F��VV�<о]~>�ť�=�	��?�"+��fM�/w����8�j�|���$=��D�<�x�?���0o�c*�a���K?�m�>vq4?�Q����|���>�Y�>��>����	�����b��{p�?;��?tt�>c܏>r?��?@D$�Z�k<
lN��7���N��{�2�]��Ë����[��EL���3?��u?��R?B<�<��>��?pg4�\{_����=)���V���"�[��> ��0&a����B�����|�o�=��-?�dT?�'H?��<|�l�ZZ<>@?Qt-?�_y?��6?>9<?�3���'?\J>�3�>u�?�m7?1=.?)�
?�aN>��=�X���<Xx��g������u��������=%t�=B1=}W�(=�6�;l.�����o��w>��m�<7b=CM�=և�=Vɦ>6�]?�U�>���>��7?.l�>|8��ڮ��/?O8=R����2���٢�:��>A�j?��?1xZ?��d>4�A�q�B���>�O�>aK&>!\>>I�>�9ｗ�E���=FT>fY>�=�L��ā�E�	����2/�<QN>i��>�9|>��@�'>~���"z���d>��Q�%κ�Y�S�X�G��1�сv�zA�>��K?>�?z��=�R龋�Ff��*)?�[<?�RM?L�?�Ó=#�۾��9��J�s'�%�>��<�����������:�/Ǵ:P�s>t5��L����:F>H9ھ3��H~��Z��W�� b9�S ��Ȇ>���vX�@�]�O��;{�>���.��W≿$:����f?����a���B@�ut��QW>rj�=%�>�c��q�=�s'�df�����>.>*׼:V���O�C��C�>�HE?^K_?�n�?&'��6�r��B����4����!ʼ��?H6�>Hd?��A>�1�=��������d�3G��%�>��>�����G�A��LG�� �$����>�:?E >��?��R?��
?-�`?t�)?TG?h�>^﷽$и��B&?L��?�܄=��Խ��T�X�8��F����>*�)?ȷB�I��>l�?�?Y�&?#�Q?R�?!�>Z� ��B@��>�Z�>��W�9a����_>֫J?O��>�;Y?1ԃ?-�=>��5�
颾Dө��N�=<>��2?�5#?g�?宸>�~�>n��� =�q�>��k?�h�?��w?C�.>N��>�4>�L�>L��=V�>���>́?��N?�{?��F?{�>`b<n�����ͽ�F������u��;�<ʜ�=wQ8��T�⭩���=щW<�j*����ᡧ�#�a��xV���/:�g�>��s>�����0>=�ľ�J��~�@>����D���ي��n:�y�=�>b ?̣�>�I#�|��=���>�C�>����7(?�?�?�#;q�b�/�ھT�K�&�>�B?2��=��l�5���u�qWh=0�m?�^?�W�G!����v? &K?��0��z:���˾+?������_?��&?�10���#?�Ё?X7[?{�?+����|:�����y6�@!7��DY=>m�>�	��/�P'c>U�M?��>���:�)6>@����'j������?��y?�c�?O��?(�->\�~���̿[�޾����m_?��>Y犾��%?�=�� ��V���a�`}���¾�]۾��	��f%��!�~� �w��>�)?)�`?�Sb?f?G�5�v�g�Yjg��f��C�F��`�]�Ց4��_��Nb��O��8<�G@��y��i#�=�}�ϔA��$�?� '?�p3���>����@�p�̾�)F>�������u�=@.���1>=�H=�i�~+�����1s ?�4�>a�>��<?�[���=�9�1��7��k��6�3>L��>�Г>���>6�#�4,�0w�˾�Ղ��˽�sw>�]b?f�J?Do?�Y�ia0�4{��r� �X8������C>g>$
�>4�Y�~(���%��]>�+7q��������	�U�=�3?l�>���>+�?��?oo
�(²�rCv�
n2�"�<#�>¨h? ��>D�>'�߽�R!�A�>�,[?\��>-@�>5����@���{���-����>��>H
�>\�%>���E_�������u�G���l>��a?j葾�S���M>i1L?bC<d�=���>z*=[�&������1 �<��!?�>�Q>-/��>[ھ۪��y����c-?:�?�ά�DD'���n>a�#?��>>��>��?�u�>>����v=�?÷^?-PD?#B?J�>'J�;F@��h���W�b�.=���>�t]>��&=�� >�����_�r)��'�d?�=ϓ��Ƽ����=ʯ <�Y<�{�:K�+>�lֿ�*�M���9��j��O,�����2%U�&�~�����i��볒��t[�歖�ʜ>>�K�,� ���[����?�R�?eI��ע�O�������*���>�a��h>�7����k�@�N���۾��˾��K��7��[?��
{���'?z�����ǿ����;>ܾ� ?�; ?Q�y?c�o�"���8�|� >#��<}������?���`�ο������^?U��>���1��  �>���>��X>�Oq>"��?螾%c�<��?��-?K��>}�r�,�ɿˊ��*�<��?b�@�PA?=�(�t�fM=4H�>@�	?��@>**0�Wg������<�>V;�?V�?ۏP=�W��?�p�e?F<�F��ٻ26�=�t�=��=�4�H�J>C�>eB��3B��۽1�4>��>� ��y�	q^����<� ]>�սrʕ�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=���Gſ�{��)�;+=rYɼ��:�@�րؽM^�����ȬY�U��)py=�5>Z�`>�u�>��D>�J>>�X?0E?�>ڧ2>>����#��D;���x�@C$��@����G��u����Ӿ�Ͼ���FA�f���ݾ&�<�2ڒ= �O�>��B}!��d�s�F���,?2�#>C{žR�L����;��Ⱦ�䩾˩K������,ʾ+0��lp��y�?�@?�d��V�V��@�r��Ƚ�nV?���z] ��ꬾA��=�h��Ӹ�<�ؗ>�+�=n���23��uQ���1?w ?{oǾ����T�#>r��Ij�<�+?��?z�<ú�>��%?b(��fν��^>H�=>�˟>a�>;�>����Sͽ�~?�T?���-�� �>�����Y{���H=�[�=�3,�"��r R>�w=?����:�؜��d�<�+W?���>q�)����}��J��:�:=��x?ߐ?�N�>��k?�B?#Ң<L���S�B�WMu=ƮW?�i?��>>���
о�[��ҳ5? �e?+�N>��h���龸�.��L��2?�n?�S?gJ���W}�������p6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������Z�=�^���?��?e�)k<&=��m�`������<�+z=��;��܁��z���x7�ہξb|��{���
[�	Q�>s�@G�3��>��S�j4�%�οϲ��0"ɾ/n���?�S�>������;Ih�/t�,�I�z?�N���#�>s�>pM��w��o�{�n�;���U��>���@C�>��S��^���|��J[1<�ʒ>�4�>���>u>���N���͙?!d���)ο|���Գ��X?9�?\�?�U?)I<�v���{��r�}�F?�Bs?
�Y?�L'���]��y5�#�j?d_��IU`���4��HE�nU>�"3?�A�>�-�б|=>,��>�d>�#/�m�Ŀ�ٶ�����t��?ω�?�o����>,��?Os+?bi��7���[��Q�*��`,��<A?�2>a���¸!��/=�&Ғ��
?@~0?�|�U.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?S	�>75�? �=�h�>��=�Y���ut��3%>�r�=`xB�l?�M?��>7a�=B7��H-�1�E�0qR��y�~�C��>�6a?.�L?�c>�����$�� ���ν$�2�4	�8>�ȗ)��>���:>&x@>X>I�G��%Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?bQo���i�B>��?"������L��f?�
@u@a�^?*SKֿ���䷾xx����=U��=6�2>}ڽ|C�=[�8=g:@����&��=Ѷ�>Qd>�p>YO>�G;>�W)>V�����!�rU�������C�����u��X\�����v�Hi�O,��3���f����ýl���FQ��R%��_����=7|_?
�D?| h?�?���.%A>%Q��.�=]~���=뼘>_p5?��Q?V�7?|�2>�^�ͯl�4���dc������Yd�>�hA>���>�V�>�k�>��M<,>oE'>�	�>��=kLE=ޒ�T\�=��>�r�>��?]��>�H<>Ɓ>4ɴ�-0��X�h��w��]̽ ��?����˩J�/���F�������'�=�`.?*d>����<п����r3H?����(�U�+�#�>�0?�XW?V�>���=�T��=>����j��=>� ��ql�L�)�?Q>&v?d�v>�Q>�\&���7�ݹW�橽��{>�X'?���,���j���F�xK�eU�=���>��_�+���r����u��I�z�r=��)?*/
?Xu�s���=�q��T���F>�^>ӹ)=�%>G>W�ǽ�4���O�&�0�.��=`˩>l�?^&+>�=�$�>BR����Q���>�@>q�+>4�@?hx$?���R��.���۽*�S^s>�?�>5i}>]>�I��E�=@w�>�Ae> ����E�&�D��U>��y� q_�bGb��
p=-T����=���=�S��=���F=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ^h�>*x�QZ����x�u�{�#=���>9H?TX��O�O�O>��u
?�?_�������ȿ�{v�y��>�?���?�m��A��@�݂�>���?�fY?�oi>
g۾�\Z����>�@?tR?6�>;:�B�'�"�?�޶?௅?�Q>��?;q?*��>�֙�L�-�u���D���=}b/;[u�>Nd�=B�ξ�vH�ן��$���S)m��L�^Jg>��%=�%�>�v�]�`��= h����	e�S��>[g>c�V>���>ID?��>�c�>��K=v���V��Mi��^�X?r��?��[��6��%\;� ���ނ�HU�>�iB?����N���Q?�\?T�~?7iB?^2 ?G���y�����ݴ���?"=/޸>a��>��>B�9��>v�P)�V�C=ϟ��3><V��
�'�y S>��>�R)?]��=��ݽ}22?>q?�<�f�>G�9��K���mF��L�>���>��>���?�X�>��޾���'թ�@����aH�	��>8\v?(�#?��>/I��]I���^3�/ޠ�E�T���T?G�?�'�=2�T?\l�?[�?�:}?��e>6�3>����k�0l>�L"?��<B�C�%�F��}�?r?N|�>�����Sн�+��0��Ǡ��߯?Tb[?f�%?!��O0a�=3¾�	�<�⻂�^�(&N<��"���>gA>퍽I��=F>?�=Ԧi�56���"<�r�=�>/�=�9��.=,?��G�{ۃ��=��r�:xD���>�IL> ����^?fl=��{�����x��	U�� �?���?Uk�?l��=�h��$=?�?T	?o"�>�J���}޾/���Pw�$~x��w�R�>���>��l���J���ԙ���F�� �Ž�+!�Ӏ�>&��>�$?4�>_�>��>�m1���G���������|���C|;�6P5�!g%��i���6#�faۼ~h����|��Ro>L�h����>�?%4M>63�>w��>�o�y0�>HK�=���>衳>E�d=�>Bq�>{3q�Q���6MR?������'���r����1B?ild?O2�>��h�ۈ����`�?��?As�?6v>�zh�6,+��k?�:�>����r
?ZV:=E���9�<�M����F����Ȩ�>XW׽m :��M�Vsf�?m
?�0?獼9�̾�;׽t�<���2���~?��??ob7�H'3���a�y�R��>��䒼6彾�bʾM�N����x������5}��4��l�=�.?��?���W��iS�D�j���I�Ό>�Q�>�*�>�I�>���>(�$��U'�0�U�����;��?	>a?�>S?��H?i�?�4t?���>�<?��,�vh�>�+�����>��?��\?ĥH?� I?��8?�{S?��#=&`^��W�| K6?�3�>��?W[
?��?�o.�����ܼ	�<�M���Ƚ�ah����qEu�.$`��r�>_�>�S?���\�8�����%k>�7?Ӎ�>��>�#��2'���U�<}�>?�
?�Q�>�����pr��Q��S�>���?H��~=�)>��=�Յ�k�Һh�=
����Ȑ="��Q;�p�<��=���=P
u�79`��[�:�;;\�<��>'J?���>H�>�E���������=�X>>,>\�>T1𾿽��얿q�m���O>8q�?��?CT�=�">ܹ�=KŮ��ξ܀��_Gʾ��;�:?�4#?��\?�J�?��@?�r?�X>�%�/g��i���s���̼?Ԓ(?��>~��Yžgb��{�9��|�>��>~�Y�"��W�&��鱾���6�Z=5w�dƀ�����C�@����=ki��,i�y��?◘?뭫;�:3�������x8����A?��>7��>mD?+�.��Gu�r� �(^�=���>�b?�#�>2�O?_<{?^�[?fT>o�8��1���ә��G3�i�!>�@?̱�?��?�y?�t�>��>ɺ)�,�[T�����b�BႾ�W=�	Z>��>�(�>;�>���=Ƚ�Z��2�>�6_�=��b>1��>!��>��>��w>�`�<c�G?���>�]��V��R줾Ń��=�ٜu?���?�+?�U=����E�QG���J�>o�?r��?Y3*?m�S����=��ּbⶾ8�q��%�>�ڹ>q1�>�ē=�sF=�b>��>K��>�)� a�q8��OM���?F?A��=��Ŀ�(q���n�"����}<瓾4Ci��`����[�|�=����	��
���i_�����U���۵�흾ǋ~�	��>��=R,�=��=�N�<=v��db�<2u@=���<�=�j��9�<ЂQ��+����4�ߺ�A<�n@=��:��˾͎}?�<I?�+?��C?��y>G>E3����>�����@?�V>2�P�A���ր;�ݧ����
�ؾ#t׾T�c��ʟ��A>QcI���>�93>�C�=t�<�/�=�"s=�Ɏ=�R�)�=�!�=uL�=�c�=I��=l�>�Y>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�;><%�=ѶO�#�1��%j�ii�MEi�0-?�F:��{����>���=1J��ʾ��I=�,>wXG=��"��[��u�=[��^�'=K��=���>��B>ۮ=?Dý��=�nS=��=I�Z>I����^��d�%�-=�=��]>F�<>b��>��?_0?[d?�0�>+ n�Ͼg3���3�>���=�B�>*��=sB>-��>i�7?�D?�K?���>�ǉ=��>��>��,�v�m�Ad��ӧ���<e��?�͆?k߸>�AS<�{A�:��Gc>��`Ž?w?$O1?�j?��>7�����^�(��O;����<�|=ٗ3>���OI��j5���������:>pݲ>�)�>eQ�>H�>�E>���>���>���=�l^�V��=B�h<�mټv���>��1�� Ļ �ƽ!�c�='A�/w���Y;u=W��=�W=vr'�%K>e��>��	>.P�>�:���݁�=�}�#�Q���;Tr��ƚT�ۉ^��Hv�M"*� �L���/>H�\>MV�X���S�>�\>3g>�u�?�Bu?L�f>ؖԼ5��N<��Usi�����GgS>�K>�|I�� B�8�2��3X�c˾Z�>Ij]>��>C�t>r�*�Ya;�|k<�V1��b>�tz!?J�ؾH��Ao�wᅿ�ۘ�駱�����z3=�y`?�
��_��=VHp?��+?9,�?�p�>TO�>�B�� ��=`Rھ���A�+�\Τ��C�<�(�>�'/?n�#?�3���dD���˾)�����>t�F�&�O�en��s�0���&S��z�>�ꪾ�Ҿ�2�(^�������B�I^q�}˺>�O?RЮ?�a��j���O��^�U���0�?EEg?0g�>�?x�?�i���N���3U�=~�n?�O�?��?|m>>��;�1� ��>�O�=��?xߨ?��?�h=4�>�r�<Fj>�x�=�~>��>�G>)kH>�G?��?2(?ˊ#�] �.%����6�3���j>��=���>ީ��ޤ>!
D=)*>4+<>�?> �W>[�>ҤK>G=j>U>�>о2��9.?3�=G��>�|5?�.�>6σ=Uu�<���=]�%��c_�>�s�r ���f��<�%�<s��<e���b��>H׿�;m?υP>`پH�?] �����P>F�]=����ľ>�=�>��>ێ�>GL>�!�>��=W���(:	>�?�M�WnF��OT����lWM>䴗�����\������1j���ž�J�7$j������<��~=���?��ֽ��b����
����K�>ux�>�?f���t����=ˎ?��>�P�ɏ�������J��?]�?�sc>��>��W?0�?>2���2�MlZ�>�u�b!A�)�d���`����������
�p���z_?\�x?K�A?�Γ<fgz>��?�&�o֏���>�/�:&;��;=�6�>�����&`�FjӾ	�þe���E>��o?+�?qM?�U�*���o�=>��F??0'?�>�?S�:?��Q?�&����6?R�<=?�Y?�w/?��,?\�
?<�l>%>>c==��=�* �����E�%�F�ʽ!X`<M�=@�1= /q=J�>��=�R�=;����%������D��;	�)=���=|Y">y��>��]?	M�>朆>��7?���;u8������'/?��9=-���F���Ţ�:�Y�>i�j?���?PbZ?^d>��A�
C��>W�>�v&>�\>[f�>q�(�E���=�H>qT>�Υ=amM�Ӂ�*�	��������<4.>Z��>w{>��1X&>y����|���^>��S�V3����M�vEG�G21��sx����>J�K?��?���=�	�g����f�7�(?��;?�JM??�?�H�=�پ�;��XJ��g�ڷ�>���<�(��u���㡿`;��h���t>7�������xd>�J����Om�#�I���龃ne=".���=h���ԾG�����=���=��¾H?#��떿�~���xK?��`=|꫾HX�����>AQ�>�>x:���E�E
?�Y��t��=+��>�_D>�%���
�#�F�
���p�>�D??�s^?@]?1-����m��82�_������DWi=�?&?ˇ�>��?�+f>���<�ϓ�:U��KJ=�M��]�>^{?}@���N�i	ؾ���]��=*��>��">��?�FW?z�?YG]?�'(?_*?�D�>�Ǽo���Ig$?�y�?�g�=�6½�m��9���8��%�>��?�,,��֪>�@?��?Ϻ*?u�E?s4?�K>H��hY<�[��>�W�>.�Q�No���(]>�;K?>��>�R?�?�
>�i1��+���&����=�>O�>?G)?Ax?���>A��>y魾1��<�*�>�?U�?)=m?d��=$->?�&*>r��>c�>��8>X�>��?H�E?j��?�xO?s�?O\�<}�ӽ9�ƽ���|�=�}�=��k�����[Ȓ��e�Õ{�t�Y=�)�=�/1��챼;��<���<��:;�9�>/�s>����M1>l�ľ�S��NA>�o��������k�:��2�=桀>Y�?힕>��#����=|��>o�>/���(?��?b?�.;�}b���ھ�K���>L�A?�3�=��l�Ny���u�P�g=�n?d�^?�W�9�����b?��]?�o��=�Z�þ߱b�����O?��
?�G���>��~?4�q?^��>��e�g9n���Eb��j��=kk�>�Y��d�b:�>�7?Y�>��b>#+�=�j۾��w�av��h?`��?O�?r��?29*>4�n��2������p���#]?��>3å���"?<���Q�ϾK���H����T⾹����򫾝"��2a��]1%�HЃ�/H׽u<�=� ?�r?A�q?;{^?H����c��r^����|V����I���E��_E��C�Y�n��������󇙾�:=X�o���E�K��?�0?z�ҽ��>�Ȋ�TG��� ���7>��x��!r�d�<=`k�� D�tH�<�wa�� �8g��F�?0��>��>�j)?`� �J��2�I�f��R&U>�*�>�u�>�?/B=-���Nc� &��K�%���P�v> ic?o�K?$�n?�r�#1��z���!�}/��K���CB>=>&ω>5�W����K&�-P>���r�*���|����	���~=��2?u:�>L��>\I�?s?�j	��\���px���1��)�<�3�>�i?�?�>���> �Ͻ�� �2��>��l?�`�>�/�>���U!��z�<6����>�ޮ>�� ?$Ao>N�*�1v[���/�7��>�Li?-����}_�儆>HQ?P�;&��<���>�'r���W���H*�Y 	>)�?,o�=t=:>�(ƾ��
���{�Yh���)?R�?΅����)���>g3#?��>��>n҄?�ћ>y����$�;��?4}^?�uI?�A?w�>��*=�W����ǽ�'��+=}��>'c\>��y=���=c����\����3&C=�8�=�
���(��7{<�즼cEX<Lz�<�l3>>�ۿ:_T�0J����d�о����Uʾke��x���A�� ����0�ҙ����f�$,ֽi	���L��)g���k�ҋ�?�y�?@�k��ݮ������.��R�>�Ѳ�؊��KeX����m0���Y�� �0$��z��������P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��q��>ޥ�>�X>�Hq>����螾x1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@�{A?��(� ���V=���>d�	?��?>�\1�
A�����&Y�>E<�?���?άM=��W���	�ւe?��<��F�J�ݻV�=4�=�.=�����J>�R�>���MA��Lܽ]�4>م>@�"�4���~^�g*�<G�]>��ս����Մ?(z\��f��/�U���X>��T?9-�>�6�=�,?�6H�]|Ͽ��\�R,a?�0�?���?'�(?�޿�Ԛ>]�ܾ��M?�C6?���>We&���t���=�XἸ����㾊&V���=���>}>fz,������O�2]�����=���cпa/���!�|=��k=kٮ��J�,|��쒫������7��R ��2�=N7>�P>�Ӄ>�q>�T�>��Q?ωp?S)?eR>��K��/����ƽҩ�yg�������:.��Ǿ!3��y�k�#��m6�[�)�� �]<����=.nL�*���c��Uh�{5Q�Yn+?�I�=g达-?����<����%Ⱦ	圽L�սn[�jW3��Jo����?a�=?=J��f�T�YW�uĮ�-�<�Y?'ϳ�c���������=8{N�:�=Ka�>�#�=W׾�~0��2E�v�,?�&?���y����7>Q��ܛ�<bMD?��?�b{={�>=?�W�
���2>��>�c�>c�?�`>�>��S�Ƚ�~?�)J?��m��Hd�lӓ>�9������j�+\�=�?�/н9_>���;�ؘ����<1��޷�9ڞR?R,�>�����ꃾu���+�<���?b4
?�|�>P|?&�2?��R=s�[@L�<z����=C�j?4�r? ��=쐽�����H����+?�b?bZ>��9�8�����.�M��Q�?d Y?��?OB��B��Б��7����0?��v?s^�xs�����G�V�h=�>�[�>���>��9��k�>�>?�#��G������zY4�%Þ?��@���?��;<��R��=�;?l\�>��O��>ƾ�z������0�q=�"�>���~ev����R,�e�8?ݠ�?���>��������=B~���@�?R�?��G~<5��ig��������<t?�=�_G��s����+9�˥ƾs��8F��qC�Oa�>@d�5��>K�ܱ῕FͿ燿~QӾ�2a��?���>����u��k�e��on��"B���C��b�����>��<>�6z�=���y�ֹ9��t���d ?
�Žh�v<����^���<���0����=xB�>4��<v�e���ݾOQ�?����ѿ���#� ��\w?�*�?�M|?Ц&?�6>����ؾ��{<�?d��?{�J?�>�둾F�D�%�j?�_��wU`���4�tHE��U>�"3?�B�>R�-�j�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*�Y�+��<A?�2>���I�!�B0=�UҒ���
?V~0?{�f.�_�_?)�a�P�p���-���ƽ�ۡ>��0��e\�,N�����Xe����@y����?M^�?g�?ڵ�� #�a6%?�>d����8Ǿ��<���>�(�>*N>�H_���u>����:�i	>���?�~�?Sj?���������U>�}?�$�>��?Hq�=�_�>�d�=��-�r#>�,�=2�>��?çM?OK�>�S�=��8�?/��YF��ER��"���C���>�a?��L?�Ob>����2�!�)hͽ�f1�rs�V@�B�,���߽�%5>��=>�>k�D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?sQo���i�B>��?"������L��f?�
@u@a�^?*��ֿū������ѾD�4>��>�>��ý�1�=�5�=���"D�����=�{�>@Ma>.��>�t�>>�>t��>w�z��������It�{�B�
���%�Hţ��5'��u�ؗ��+оۛ�����c+üW�\�򐾘?۽�����=�RT?:1Q?\{p?���>P~��_!>-����=T_ �Fe=V�>ܧ2?�hL?��)?q��=�Μ���c���UΦ�������>&H>"��> �>���>�i�:�F>��>>_+�> >=�'=�k��� =ZxT>���>Hl�>�o�>4�>+a	>��I���6�n�dN*���B��h�?Wʞ��I�ܝ���Ҵ��H۾<�F>H�)?]�=&����ο�ج���J?�٢��c��x6�p6�=0;?KGd?ێ>/����Z�=�=7��h�?���f>���<�����	�	�>?�M�>h�>>j�P�OlJ��`��u����>��>?����B�:���d�@7����^#�>�)?tt�[� ����������\��>=L�-?�M6?k�O��!Ͼ^���꿾� �=$a�>�[�����><<{>�K�1�*=M� �	R����K=a��>�|?�	�>��=��v>`.����^����>Y�>�j>"�5?�|6? �
��+��Zqd��F��e�>E��>/��>tna>�M�LPp=\��>*eZ>[@u=�3]=��4��vD�>x�߈����&��TļV��B�=���=LI������"�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ&h�>�w�zZ�������u���#=���>�8H?�V��D�O�f>��v
?T?=_�ꩤ���ȿc|v�/��>�?���?N�m��A���@����>2��?�gY?pi>g۾_Z�V��>D�@?�R?��>Q9�T�'���?�޶?ů�?�I>q��?�s?�l�>$/x�oZ/�>6��Ȗ��gt=��[;~c�>\V>�����fF��ד�rh���j�����a>��$=��>6E�C4���7�=N���NH����f����>k,q>��I>W�>S� ?�b�>٦�>w}=Ck��]���������K?���?0���2n��M�<{��=�^��&?�I4?3j[�{�Ͼ�ը>޺\?j?�[?d�>=��P>��F迿8~��H��<��K>54�>�H�>�$���FK>��Ծ�4D�ip�>�ϗ>I����?ھ�,��LT��AB�>�e!?���>�Ү=� ?��#?D�j>e�>�^E�h:����E����>ў�>bD?��~?��?"ٹ��\3����"塿�[�>N>��x?MW?�ŕ>����	����=F���H�m������?�ug?�H录?.�?��??�A?F.f>���ؾ"���~�>�0?�I�FP��%;��UH���?��?���>Aۨ����p����#���
�w~&?��_?��?$M�~�j���|K>=���Ux:e�Y=4{����>��6> \���z�=`"�>� ={��i��R�<�k4>;V�>ah�=��E�%Й�/=,?�G�wۃ���=��r�?xD���>�IL>����^?>l=��{�����x��#	U�� �?���?[k�?��;�h��$=?�?P	?n"�>�J���}޾,�ྠPw�!~x��w�T�>���>��l���I���י���F��B�ŽB�L��/�>�e�>�x:?ҝ�>�h>>d�>^��������S���K��e��]��V��X��_:Y�hL���f1�ظ�9���Ȩ��x�>���/��>Ȧ�>�n>S]�>�>�>�� =_��=4Զ=��>=�>/o�=W\>3KA>��>s=~KR?������'�\�辕����2B?�qd?M1�><i�㉅�K���?���?As�?=v>8h��,+�(n?�=�>���p
?@R:=;��;�<vU�� ��b3��H�/��>�A׽t :�dM�Enf�Tj
?40?���Ӌ̾P;׽�+ؾ�	�=W�w?f��>/G
�1�_�F���V�H�E�o��S���M�D3��2������.��v� |����/�R�;�ח5?�?�n��� ��2���mb��^"����>=�>r�x>>�>_��=�����$��(V�� �Kl��Oo�>?�L?V��>�F?�pS?��B?��=?�/�>\�
>�wҾ�
�>������>gx�>�??�I"?��?�`N?�$?A�S>�x�=�Oھ��ž��	?�f ?�*?�ŵ>�s�>��Z�n�4[�<9i�Tn���A(>�E�<�(+>!�����㽄��X�/>�J?8��8��-��8�j>6?���> �>'t����~���	=�8�>��
?��>������q�m�����>�҂?��H�=��*>���=�us�V'�:,6�=���ڕ=wG��C<��^(<H�=��=;�m�>)I�ڷ�9#�6;�C�<B�?�b(?x��>,�K>Ǯo�4��G���J>nh�>�.�>��>*~Ⱦ$n{��<����]����>x;�?婶?h� >h� >�i�=�Ի�/�þr	��~��ҩF=Cz?~�&?��I?Lc�?j�?��?��=���9��lO����P��?��B?�zP>�%��8���X��&��G�?w��>��h�5��<�D�F�A���!����=��o� Oh�mĪ�;k�oP��<�"<���?�p�?�����O	��ԧ��8¾n�?���>Lv>��#?�G<���N�/57�]�/>�
�>��/?�_�>��R?�{�?�=`?M��>��@�����2�z=O>�x?��r??�?�l?!��>\`�>A���ǚ���7���`�b~���o_�^?����[>27>���>4ϣ>Œ�<�$�y)�z��Ȫ�<�c>{ �>��o>ٔ�>�>ep=ݜG?҇�>����ͬ�����Uą��|B�W�u?�5�?�0,?��$=DO�ѥD��}��~�>	(�?A��?B +?��N���=��ټu��i6t�Դ�>[��>,�><�=�:[=�>8�>ݔ�>R������8��rZ�h�?!�F?_,�=�,��E�y��,�:8N��B�=��<����n@�;�>P���=B���ݔ�5>���@]��߲��X��船��ݒ��b����>(~=\h>�H�=�I=�Fۼc�G��=��:�}O�p�<���<�r����	<e�̽n\1<qw�<��=�����˾�8}?XI?��+?/�C?�ry>s�>��2�>'�>�Y��?Y?l�T>�wM�}E��F�;��ĩ����Kqؾ�[׾d�,���>II��>5�1>�c�=�Y�<J��=�s=6}�=�V�?=��=f+�=㖬=2�=�>�.>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��7>��>׼R��n1���\��b��Z���!?�0;�� ̾��>mu�=
߾{rƾ֐.=�?6>!jb=e�M\��=m�{��;=�k==ى>GD>K��=Z6���>�=ɹI=BR�=#�O>/ɛ�e8�	4,�(�5=U��=�b>�&>R�>�,?�!B?jq3?^n�>XO���̾Y�� K)>}8 >�c�>��>�ו>�j�>!~2?�U?Z�]?�K�>V�1>B2�>(͌>b�@�潀�-G���ߎ�aR�= ˌ?$�y?���>蛐>D��@�0��2N��Y����>�+-?�]?E�>�U����\Y&���.�`����*��+=�mr�_RU������m�M�㽕�=�p�>���>��>\Ty>l�9>��N>A�>��>�=�<q�=�ꌻ���<���ɲ�=������<3yż�Q�� �&���+�����^͍;<��;��]<K��;1�=���>��>?�>H?�=�j��@]/>ʘ���L��r�=͘���>B���c��:~�?�.�8���A>�V>Y��f1��Ⱦ?lZ>�4@>U��?�,u?�E >�F�ĦԾd����f�R�T�	��=�T>Np?��~;�8�_�%M���Ѿ���>&Ŏ>g+�>�Do>>7,�v>�?z=��hw5�X�>Kj��H�(�+�!#q�����"����h�	Ŋ�2	C?I��$�=��}?ݷI?�?��>ϯ���׾l�3>�ʁ��5�<T����o�J����?h�%?@	�>�k���C�<�˾�ൽ[�>ؕO��LO�������1�Z�ջ_��}[�>i��hϾ��4�`ކ��r��Q�B��
{�)V�>rM?�/�?Xcb�f@��[�N��A��u���?��g?�Ң>?�?X-?=8�����Eu����=�.m?B#�?���?��>���=�w�����>�!?g��?ܐ?��q?#�'�t�?���<r.�=����2�=�->�a�=�r�=7L?)�?�	
?����
�Q��j��:�9�=&��=�r�>�^>�;f>�3>�m]=F��=WM>$ʑ>�>�e>��>(\�>}���V>�*�?��]>���>=�(?��>'�=�d���m�=��\V��gn�0�����;���J�!�V<��N��\�>���B�?A`>��ѾxZ!?P�پ�w���Ƒ=�c>�`�<＜>��r=�+>_O}>���>���=�)n>�\>��Ӿ�>�:��"�4B�FUS�ԍվ,Dz>�Ğ�;�.���SX�=O�y��y��8�i�o���lc=�7�<Wc�?O`����l���)�W��Q?cԫ>��6?.މ�����>>e��>��>L9���Ӕ��z��$'��V�?:��?|;c>Q�>-�W?�?�1�E3�uZ�j�u��'A�ie��`�X፿����9�
������_?��x?yA?'U�<�9z>(��?O�%�ӏ�;)�>Q/�';��8<=D+�>�)����`���ӾN�þ7�mHF>i�o?%�?�X?�RV���n��|(>�:?!�1?�3t?k�0?�:?w��a�$?��1>͞?�U?��5?� /?�?�%2>�m�=�����+=�����Њ��~ѽ#hϽ�e񼐁4=�+=&��:�	�;�5=I/�<��ټ���h9;�ɘ��N�<�D=�ՠ=F�=���>�^?:A ? �>��6?��;��07��l��sp-?��;=�v��q�~�~�7�ܾX�>h�k?�R�?վZ?I��>@�<���;�K9>8:u>^�6>��b>(��>�K��ܳB��{�<�r�=736>[bj=����g�����A��4*;�|%>s8�>tp>����8p>5�߾��:��Z>e���� ھ=0�W�A�'�*�����:�>ZMT?_R�>4gF;��~$=�sl�� ?4�??y<Q?�=�?Gw>����+�.��#�bm4��c/>ߡ�JϾ���Ui���E�+5�=�p�>�ύ�����xd>�J����Om�#�I���龃ne=".���=h���ԾG�����=���=��¾H?#��떿�~���xK?��`=|꫾HX�����>AQ�>�>x:���E�E
?�Y��t��=+��>�_D>�%���
�#�F�
���p�>�D??�s^?@]?1-����m��82�_������DWi=�?&?ˇ�>��?�+f>���<�ϓ�:U��KJ=�M��]�>^{?}@���N�i	ؾ���]��=*��>��">��?�FW?z�?YG]?�'(?_*?�D�>�Ǽo���Ig$?�y�?�g�=�6½�m��9���8��%�>��?�,,��֪>�@?��?Ϻ*?u�E?s4?�K>H��hY<�[��>�W�>.�Q�No���(]>�;K?>��>�R?�?�
>�i1��+���&����=�>O�>?G)?Ax?���>A��>y魾1��<�*�>�?U�?)=m?d��=$->?�&*>r��>c�>��8>X�>��?H�E?j��?�xO?s�?O\�<}�ӽ9�ƽ���|�=�}�=��k�����[Ȓ��e�Õ{�t�Y=�)�=�/1��챼;��<���<��:;�9�>/�s>����M1>l�ľ�S��NA>�o��������k�:��2�=桀>Y�?힕>��#����=|��>o�>/���(?��?b?�.;�}b���ھ�K���>L�A?�3�=��l�Ny���u�P�g=�n?d�^?�W�9�����b?��]?�o��=�Z�þ߱b�����O?��
?�G���>��~?4�q?^��>��e�g9n���Eb��j��=kk�>�Y��d�b:�>�7?Y�>��b>#+�=�j۾��w�av��h?`��?O�?r��?29*>4�n��2������p���#]?��>3å���"?<���Q�ϾK���H����T⾹����򫾝"��2a��]1%�HЃ�/H׽u<�=� ?�r?A�q?;{^?H����c��r^����|V����I���E��_E��C�Y�n��������󇙾�:=X�o���E�K��?�0?z�ҽ��>�Ȋ�TG��� ���7>��x��!r�d�<=`k�� D�tH�<�wa�� �8g��F�?0��>��>�j)?`� �J��2�I�f��R&U>�*�>�u�>�?/B=-���Nc� &��K�%���P�v> ic?o�K?$�n?�r�#1��z���!�}/��K���CB>=>&ω>5�W����K&�-P>���r�*���|����	���~=��2?u:�>L��>\I�?s?�j	��\���px���1��)�<�3�>�i?�?�>���> �Ͻ�� �2��>��l?�`�>�/�>���U!��z�<6����>�ޮ>�� ?$Ao>N�*�1v[���/�7��>�Li?-����}_�儆>HQ?P�;&��<���>�'r���W���H*�Y 	>)�?,o�=t=:>�(ƾ��
���{�Yh���)?R�?΅����)���>g3#?��>��>n҄?�ћ>y����$�;��?4}^?�uI?�A?w�>��*=�W����ǽ�'��+=}��>'c\>��y=���=c����\����3&C=�8�=�
���(��7{<�즼cEX<Lz�<�l3>>�ۿ:_T�0J����d�о����Uʾke��x���A�� ����0�ҙ����f�$,ֽi	���L��)g���k�ҋ�?�y�?@�k��ݮ������.��R�>�Ѳ�؊��KeX����m0���Y�� �0$��z��������P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��q��>ޥ�>�X>�Hq>����螾x1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@�{A?��(� ���V=���>d�	?��?>�\1�
A�����&Y�>E<�?���?άM=��W���	�ւe?��<��F�J�ݻV�=4�=�.=�����J>�R�>���MA��Lܽ]�4>م>@�"�4���~^�g*�<G�]>��ս����Մ?(z\��f��/�U���X>��T?9-�>�6�=�,?�6H�]|Ͽ��\�R,a?�0�?���?'�(?�޿�Ԛ>]�ܾ��M?�C6?���>We&���t���=�XἸ����㾊&V���=���>}>fz,������O�2]�����=���cпa/���!�|=��k=kٮ��J�,|��쒫������7��R ��2�=N7>�P>�Ӄ>�q>�T�>��Q?ωp?S)?eR>��K��/����ƽҩ�yg�������:.��Ǿ!3��y�k�#��m6�[�)�� �]<����=.nL�*���c��Uh�{5Q�Yn+?�I�=g达-?����<����%Ⱦ	圽L�սn[�jW3��Jo����?a�=?=J��f�T�YW�uĮ�-�<�Y?'ϳ�c���������=8{N�:�=Ka�>�#�=W׾�~0��2E�v�,?�&?���y����7>Q��ܛ�<bMD?��?�b{={�>=?�W�
���2>��>�c�>c�?�`>�>��S�Ƚ�~?�)J?��m��Hd�lӓ>�9������j�+\�=�?�/н9_>���;�ؘ����<1��޷�9ڞR?R,�>�����ꃾu���+�<���?b4
?�|�>P|?&�2?��R=s�[@L�<z����=C�j?4�r? ��=쐽�����H����+?�b?bZ>��9�8�����.�M��Q�?d Y?��?OB��B��Б��7����0?��v?s^�xs�����G�V�h=�>�[�>���>��9��k�>�>?�#��G������zY4�%Þ?��@���?��;<��R��=�;?l\�>��O��>ƾ�z������0�q=�"�>���~ev����R,�e�8?ݠ�?���>��������=B~���@�?R�?��G~<5��ig��������<t?�=�_G��s����+9�˥ƾs��8F��qC�Oa�>@d�5��>K�ܱ῕FͿ燿~QӾ�2a��?���>����u��k�e��on��"B���C��b�����>��<>�6z�=���y�ֹ9��t���d ?
�Žh�v<����^���<���0����=xB�>4��<v�e���ݾOQ�?����ѿ���#� ��\w?�*�?�M|?Ц&?�6>����ؾ��{<�?d��?{�J?�>�둾F�D�%�j?�_��wU`���4�tHE��U>�"3?�B�>R�-�j�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*�Y�+��<A?�2>���I�!�B0=�UҒ���
?V~0?{�f.�_�_?)�a�P�p���-���ƽ�ۡ>��0��e\�,N�����Xe����@y����?M^�?g�?ڵ�� #�a6%?�>d����8Ǿ��<���>�(�>*N>�H_���u>����:�i	>���?�~�?Sj?���������U>�}?�$�>��?Hq�=�_�>�d�=��-�r#>�,�=2�>��?çM?OK�>�S�=��8�?/��YF��ER��"���C���>�a?��L?�Ob>����2�!�)hͽ�f1�rs�V@�B�,���߽�%5>��=>�>k�D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?sQo���i�B>��?"������L��f?�
@u@a�^?*��ֿū������ѾD�4>��>�>��ý�1�=�5�=���"D�����=�{�>@Ma>.��>�t�>>�>t��>w�z��������It�{�B�
���%�Hţ��5'��u�ؗ��+оۛ�����c+üW�\�򐾘?۽�����=�RT?:1Q?\{p?���>P~��_!>-����=T_ �Fe=V�>ܧ2?�hL?��)?q��=�Μ���c���UΦ�������>&H>"��> �>���>�i�:�F>��>>_+�> >=�'=�k��� =ZxT>���>Hl�>�o�>4�>+a	>��I���6�n�dN*���B��h�?Wʞ��I�ܝ���Ҵ��H۾<�F>H�)?]�=&����ο�ج���J?�٢��c��x6�p6�=0;?KGd?ێ>/����Z�=�=7��h�?���f>���<�����	�	�>?�M�>h�>>j�P�OlJ��`��u����>��>?����B�:���d�@7����^#�>�)?tt�[� ����������\��>=L�-?�M6?k�O��!Ͼ^���꿾� �=$a�>�[�����><<{>�K�1�*=M� �	R����K=a��>�|?�	�>��=��v>`.����^����>Y�>�j>"�5?�|6? �
��+��Zqd��F��e�>E��>/��>tna>�M�LPp=\��>*eZ>[@u=�3]=��4��vD�>x�߈����&��TļV��B�=���=LI������"�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ&h�>�w�zZ�������u���#=���>�8H?�V��D�O�f>��v
?T?=_�ꩤ���ȿc|v�/��>�?���?N�m��A���@����>2��?�gY?pi>g۾_Z�V��>D�@?�R?��>Q9�T�'���?�޶?ů�?�I>q��?�s?�l�>$/x�oZ/�>6��Ȗ��gt=��[;~c�>\V>�����fF��ד�rh���j�����a>��$=��>6E�C4���7�=N���NH����f����>k,q>��I>W�>S� ?�b�>٦�>w}=Ck��]���������K?���?0���2n��M�<{��=�^��&?�I4?3j[�{�Ͼ�ը>޺\?j?�[?d�>=��P>��F迿8~��H��<��K>54�>�H�>�$���FK>��Ծ�4D�ip�>�ϗ>I����?ھ�,��LT��AB�>�e!?���>�Ү=� ?��#?D�j>e�>�^E�h:����E����>ў�>bD?��~?��?"ٹ��\3����"塿�[�>N>��x?MW?�ŕ>����	����=F���H�m������?�ug?�H录?.�?��??�A?F.f>���ؾ"���~�>�0?�I�FP��%;��UH���?��?���>Aۨ����p����#���
�w~&?��_?��?$M�~�j���|K>=���Ux:e�Y=4{����>��6> \���z�=`"�>� ={��i��R�<�k4>;V�>ah�=��E�%Й�/=,?�G�wۃ���=��r�?xD���>�IL>����^?>l=��{�����x��#	U�� �?���?[k�?��;�h��$=?�?P	?n"�>�J���}޾,�ྠPw�!~x��w�T�>���>��l���I���י���F��B�ŽB�L��/�>�e�>�x:?ҝ�>�h>>d�>^��������S���K��e��]��V��X��_:Y�hL���f1�ظ�9���Ȩ��x�>���/��>Ȧ�>�n>S]�>�>�>�� =_��=4Զ=��>=�>/o�=W\>3KA>��>s=~KR?������'�\�辕����2B?�qd?M1�><i�㉅�K���?���?As�?=v>8h��,+�(n?�=�>���p
?@R:=;��;�<vU�� ��b3��H�/��>�A׽t :�dM�Enf�Tj
?40?���Ӌ̾P;׽�+ؾ�	�=W�w?f��>/G
�1�_�F���V�H�E�o��S���M�D3��2������.��v� |����/�R�;�ח5?�?�n��� ��2���mb��^"����>=�>r�x>>�>_��=�����$��(V�� �Kl��Oo�>?�L?V��>�F?�pS?��B?��=?�/�>\�
>�wҾ�
�>������>gx�>�??�I"?��?�`N?�$?A�S>�x�=�Oھ��ž��	?�f ?�*?�ŵ>�s�>��Z�n�4[�<9i�Tn���A(>�E�<�(+>!�����㽄��X�/>�J?8��8��-��8�j>6?���> �>'t����~���	=�8�>��
?��>������q�m�����>�҂?��H�=��*>���=�us�V'�:,6�=���ڕ=wG��C<��^(<H�=��=;�m�>)I�ڷ�9#�6;�C�<B�?�b(?x��>,�K>Ǯo�4��G���J>nh�>�.�>��>*~Ⱦ$n{��<����]����>x;�?婶?h� >h� >�i�=�Ի�/�þr	��~��ҩF=Cz?~�&?��I?Lc�?j�?��?��=���9��lO����P��?��B?�zP>�%��8���X��&��G�?w��>��h�5��<�D�F�A���!����=��o� Oh�mĪ�;k�oP��<�"<���?�p�?�����O	��ԧ��8¾n�?���>Lv>��#?�G<���N�/57�]�/>�
�>��/?�_�>��R?�{�?�=`?M��>��@�����2�z=O>�x?��r??�?�l?!��>\`�>A���ǚ���7���`�b~���o_�^?����[>27>���>4ϣ>Œ�<�$�y)�z��Ȫ�<�c>{ �>��o>ٔ�>�>ep=ݜG?҇�>����ͬ�����Uą��|B�W�u?�5�?�0,?��$=DO�ѥD��}��~�>	(�?A��?B +?��N���=��ټu��i6t�Դ�>[��>,�><�=�:[=�>8�>ݔ�>R������8��rZ�h�?!�F?_,�=�,��E�y��,�:8N��B�=��<����n@�;�>P���=B���ݔ�5>���@]��߲��X��船��ݒ��b����>(~=\h>�H�=�I=�Fۼc�G��=��:�}O�p�<���<�r����	<e�̽n\1<qw�<��=�����˾�8}?XI?��+?/�C?�ry>s�>��2�>'�>�Y��?Y?l�T>�wM�}E��F�;��ĩ����Kqؾ�[׾d�,���>II��>5�1>�c�=�Y�<J��=�s=6}�=�V�?=��=f+�=㖬=2�=�>�.>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��7>��>׼R��n1���\��b��Z���!?�0;�� ̾��>mu�=
߾{rƾ֐.=�?6>!jb=e�M\��=m�{��;=�k==ى>GD>K��=Z6���>�=ɹI=BR�=#�O>/ɛ�e8�	4,�(�5=U��=�b>�&>R�>�,?�!B?jq3?^n�>XO���̾Y�� K)>}8 >�c�>��>�ו>�j�>!~2?�U?Z�]?�K�>V�1>B2�>(͌>b�@�潀�-G���ߎ�aR�= ˌ?$�y?���>蛐>D��@�0��2N��Y����>�+-?�]?E�>�U����\Y&���.�`����*��+=�mr�_RU������m�M�㽕�=�p�>���>��>\Ty>l�9>��N>A�>��>�=�<q�=�ꌻ���<���ɲ�=������<3yż�Q�� �&���+�����^͍;<��;��]<K��;1�=���>��>?�>H?�=�j��@]/>ʘ���L��r�=͘���>B���c��:~�?�.�8���A>�V>Y��f1��Ⱦ?lZ>�4@>U��?�,u?�E >�F�ĦԾd����f�R�T�	��=�T>Np?��~;�8�_�%M���Ѿ���>&Ŏ>g+�>�Do>>7,�v>�?z=��hw5�X�>Kj��H�(�+�!#q�����"����h�	Ŋ�2	C?I��$�=��}?ݷI?�?��>ϯ���׾l�3>�ʁ��5�<T����o�J����?h�%?@	�>�k���C�<�˾�ൽ[�>ؕO��LO�������1�Z�ջ_��}[�>i��hϾ��4�`ކ��r��Q�B��
{�)V�>rM?�/�?Xcb�f@��[�N��A��u���?��g?�Ң>?�?X-?=8�����Eu����=�.m?B#�?���?��>���=�w�����>�!?g��?ܐ?��q?#�'�t�?���<r.�=����2�=�->�a�=�r�=7L?)�?�	
?����
�Q��j��:�9�=&��=�r�>�^>�;f>�3>�m]=F��=WM>$ʑ>�>�e>��>(\�>}���V>�*�?��]>���>=�(?��>'�=�d���m�=��\V��gn�0�����;���J�!�V<��N��\�>���B�?A`>��ѾxZ!?P�پ�w���Ƒ=�c>�`�<＜>��r=�+>_O}>���>���=�)n>�\>��Ӿ�>�:��"�4B�FUS�ԍվ,Dz>�Ğ�;�.���SX�=O�y��y��8�i�o���lc=�7�<Wc�?O`����l���)�W��Q?cԫ>��6?.މ�����>>e��>��>L9���Ӕ��z��$'��V�?:��?|;c>Q�>-�W?�?�1�E3�uZ�j�u��'A�ie��`�X፿����9�
������_?��x?yA?'U�<�9z>(��?O�%�ӏ�;)�>Q/�';��8<=D+�>�)����`���ӾN�þ7�mHF>i�o?%�?�X?�RV���n��|(>�:?!�1?�3t?k�0?�:?w��a�$?��1>͞?�U?��5?� /?�?�%2>�m�=�����+=�����Њ��~ѽ#hϽ�e񼐁4=�+=&��:�	�;�5=I/�<��ټ���h9;�ɘ��N�<�D=�ՠ=F�=���>�^?:A ? �>��6?��;��07��l��sp-?��;=�v��q�~�~�7�ܾX�>h�k?�R�?վZ?I��>@�<���;�K9>8:u>^�6>��b>(��>�K��ܳB��{�<�r�=736>[bj=����g�����A��4*;�|%>s8�>tp>����8p>5�߾��:��Z>e���� ھ=0�W�A�'�*�����:�>ZMT?_R�>4gF;��~$=�sl�� ?4�??y<Q?�=�?Gw>����+�.��#�bm4��c/>ߡ�JϾ���Ui���E�+5�=�p�>�ύ��O����>������ؿi��R�v������<>��Ue�<���B����U�Y��=2�>�3Ѿ�_(�g�L+��B J?K��=�s��J�[�w�����=MT�>o9�>XP~�W|S���,��K�����<�d�>H>a�d�+���A��p�g>!I?��h?x�i?�K��Ɓ�.S�DU
�0A��u~��Ҁ?B��>��?��F>QC�=��Ѿ�$�o�s��Z��s�>4?W��aA��՞�H� �A�,H�>�B�>H�>��?ܻE?�;�>��b?��?Ka�>݈�>駾�W~��A�$?`u�?�U�=��'�_���9�	�=��V�>�k!?�3���>��?ʝ ?a�!?�L?�|?�  >�����C�*��>���>�>Z�B󰿻 �>�H?m�>�}Y?ۂ?��=>�2�@L���,׽�>m��=)�0?�;,?�M?2��>-��>Gڟ��~�=/@�>�.d?�t�?�_?l�=D?�S�=���>wk=��r>+��>�?�~Q?�xm?��<?��>�{�<�-���?���U��n�:���k<vB�r�=1M�0����V;�$�<X�<oy^�����q���7���b�j(�<�=�>�u>�^��*�1>biľ�{���?>X����́���@<�b��=M7�>�?F�>H� �"�=M�>���>�p��d(?}U?�v?_�;/�b��ھ��L��>A?���=��l�#��
�t�UMg=jAn?�b^?��R�Y���=�b?��]?�g�=���þ��b�ډ�Y�O?4�
?��G���>��~?M�q?.��>'�e�
:n����Cb���j��ж=r�>4X�d�d��?�>��7?�N�>��b>�$�=[u۾&�w�fq��d?f�?�?���?�+*>��n�[4�O<��il���]?ð�>F����"?J�+��/Ѿ�+���\��?�⾠���̫����m���ԫ$���)ؽ;�=�i?��s?W�q?o�_?� ��Rd��~^�6��d�V�eq�����iE�E�C���C���m��C���J�����1=� ���&�X,�?	4C?^�7����>�j��LKپ����U%=>����lm�i�`>:�U=�<>eIr=x��}[u��̾�?�??P�@?��c��]X�<D��E�����̈�Ar3>���>��1?���>Eb�=��$<�@��y�d=����@�x>�lc?K?�o?B��~u1�����6 �9�L�������G>�)>��>!`�oK��c%���=���q�����J��Y'�r=ă1?���>1��>���?=�?K��-W����s��4/�n=<*�>��f?���>�@�>\2ƽ\8!����>Rwj?Wi�>��>2:��j��3�y���ѽ�|�>S(�>8��>�0l>��#�x�T�SX��壊�R=/�c�>�o?6)��倾wa�> �H?&,="�=��>��u�����۾�A0�lK>\�?h��=>>D;ǾO���%��R鑾�_ ?�d?�F���_��S�>�)?�a�>���>E�?��>y��W���7�>>\?�]R?�TM?^"�>�v=C�,�Z���f5�8�=�~�>t�_>!��=2'@=�����ig�d�$��M=
>�<@B�����䀚���;$�k=���<�f!>5[ѿ��S��������������d��e�n�r�P�C�	�Q�yr`�t6�n���P�=�s-�����M1��o�|��c�?4��?)Ƚp,m�nȍ�@@��]�����>�����O��о�޽<ܽ��
��~�bG��B�P��u|�:u��S�'?�����ǿ󰡿�:ܾ1! ?�A ?A�y?��1�"���8�� >�B�<�,����뾪����οA�����^?���>��/��q��>Υ�>�X>�Hq>����螾�1�<��?.�-?	��>Ǝr�/�ɿ]���hä<���?,�@�:>?��#�*��㚖=�\�>��?Q�+><�)�	F�������>���?뺅?|[�=ϥU�u�!��6b?�	�E$<��a!�̣�=���=4�<�����I>�,�>I�<���J�@0a��u>rK�>Z��ȵ�EJZ�4D��6DA>���KI��4Մ?+{\��f���/��T��
U>��T?�*�>]:�=��,?Z7H�`}Ͽ�\��*a?�0�?���?$�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�ԅ�=i6�Z���|���&V�m��=Z��>j�>ǂ,�ދ���O��I��Q��=�����˿Ź#���$�y)�<�~=�	��DJ��r�;ܹ�=�5��������.��=��=�{�=��->�i>S�q>�]?^`^?u�>q�V>�D�p�g��*���B��G�O���;�1#���M���˾�\�F績��[��� ���<�B��=�Q�����x� ���b���F���.?Ys#>�ʾѧM�ؑ9<?�ɾ����u���N��~�̾�1�}An�u˟?hB??�����V���a���?��1�W?K����1����=͐����=#��>���=��⾔�2��fS�@x%?�7 ?2Ȭ�a#���R�>e����R=�/?j��>����D$>��?4�b� ��7e>��H=��`>�[�>mW>������u?�l?���=��P�H�>79ž:���>:�=Ya߻���1;���>LH>��W�����m=���=U?���>�Q(��	�;䊾Sj'���r=�^x?z1�>R��>��e?��;?��<;����R��N�Ɏ=��V?�c?f�>���EҾ�š�=^6?L�d?$5X>�JW�̚־�V*�-����?/�e?� ?8��	�~�J���%���R6?�w?�]�q����V�d�\�z��>P��>�K�>+�:���>�d??��'��
�������5��~�?�_@M��?� <ei �E�=x�?���>�P�x�ƾ�x���ϵ�Fx=�k�>�ը��7v�v��P�1��8?㜃?��>Sc��!��e�=�;r�j�?��j?ƻ��r�ɽ)0��u�30���ܼ�6���H=b�=M��f��������#�3uҾ,�	�̆�>@�G���z�>~��0'�i�¿�m��)��d���?HO�>$���؏���c�@{�%�I��WU��ݾs��>�>��t�j�냿WT��ᅽ��?tފ��F><�m=P�¾�҅���"�B%>��>>)Yu=1�~�Ͷ��+�?��徠A߿�%����D���i??	ԣ?#��>0�>�p=���1���/X ?&?Ik?~\�>�T=Ă��i�j?�^���U`�;�4��IE�	U>�#3?�D�>G�-�H�|=�!>L��>�e>,$/���Ŀ�ض��������?��?jo�@��>���?hs+?mi��7���[����*��)�S=A?�
2>k���+�!�U1=��ђ��
?n}0?{�4-���_?C�a�O�p���-�
�ƽ�ܡ>��0�Gf\��-��]��rYe�����Cy�U��?<^�?��?��8 #�36%?6�>�����6Ǿ,�<���>()�>�%N>�C_�T�u>����:�sc	>��?}~�?�h?��������"V>��}?V-�>��?���=���>���=-�����'�"M$>��=G>�L=?�^M?���>���=��8��4/��IF��R�0��ͰC�X��>l�a?	�L?��c>�&���0��!�l�ɽf�0����G@��1��ݽ�J6>�H>>�[>�wE��aҾ�?p�E�ؿ
j��Nq'�{54?w��>b�?X���t����~;_?z�>�6��+���%��BB�A��?kG�?>�?��׾�S̼>��>J�>6�Խ��������*�7>1�B?���D��\�o� �>���?�@�ծ?[i�U	?)��T��'f~���A7����=�7?�E�[�z>���>���=�kv�"����s�z��>�?�?u�?R��>&�l?o��B��	2=�8�>�k?%{?��o����B>r�?��I���)J��f?��
@bt@�^?�뢿��ؿ`����;��޾">��p��=��F��
�=~"�>m>��=��=�J>�>���>��E>8!>�1;>+�������ٓ�,kM�y��]���Q������p'���[�W�(uݾT�^�&��3����@�O�8�r����=�ZT?$�P?��o?o?^�_��O>�����=vo$�?!�=��>e1?�}M?�*?�*�=uf��v�e�I��������=���y�>݃F>���>���>	�>���I>bLA>^ځ>�k>�*=�?F�?�=N>I-�>��>�b�>�gV>9�,>�p��Ḳ�Нo��n}����v~�?�r���$D�[<��?#���n���`�=+&?V��=3(��S�̿����ĴH?[Ɨ�o��[M&��!�=25?�)_?�+>�G��{ ׼\p.>L.��j����=���SM������f>=i?��g>Q�o>�2���4��N�%��Ȟ�>17?林�R�,�,�r��1K�"�߾\�B>��>]���/��Z_��z�}�/&d��E =�[<?��?�}��Nr��$|��I�����f>�wY>3;�<?ϩ=U�E>�EJ��?��$;D�6zC<t��=mf>ة�>��8>kM�;���>����n�$�v��>��>�6	>�Y:?$?���n̽���������l>T^�>�	T>�y|=1�5���5U�>�bx>Rq�;��\��|B��!P��"�>,���+���v�̥�����+�>|�=Z��|�k����=�~?���䈿��Oe���lD?I+? �=�F<��"�D ���H��J�?q�@m�?��	��V�K�?�@�?�
����=}�>׫>�ξC�L�Ա?/�Ž7Ǣ�̔	�D)#�dS�?��?��/�Rʋ� l��6>_%?ѰӾ\h�>Sx��Z�������u���#=P��>�8H?�V����O�#>��v
?�?�^�ݩ����ȿ1|v����>I�?���?d�m��A���@�g��>:��?�gY?�oi>�g۾`Z����>��@?�R?�>�9�J�'���?�޶?ϯ�?��G>9��?��s?��>�x�H�/��P��E���g�t=>�:k��>��>�����E�fl���z��6"k�J��8^]>��)=��>����U��?.�=>�����`���>��p>4DL>aW�>q��>���>ט�>�=��� ��������K?���?���*3n�4�<���=�^��'?eH4?�][���ϾԨ>[�\?>?([?�c�>���>��P迿�}��f��<��K>!4�>bG�>j!���HK>��ԾI6D��p�>ZЗ>x���?ھ�,�����yB�>�e!?��>�Ю=� ?^�#?�k>�U�>IE��-����E���>���>�M?��~?��?4����I3����?ۡ��u[�o}N>�y?RK?ˈ�>�����{����>�#GE��B����?-]g?R�佋�?�+�?�??-�A?-f>����׾����'��>�D?P���5�jQ��\P���?d	?���>2�Y=�xz�Mq�W����
��O?As?}�+?C���SjM��h���^=�a<VPx=^��=��g�tI>��_=3���t3!=�!�=�ĵ�s9����&���=�h�<?��>P�0>(z������.?�[һ����$}={w�c8C�Z��>^^>֍ʾ]�`?m*�R������Sٝ��rg���?���?�f�?iν*�f���:?���?!]?l�>ˉ��������T?h�w�f�`�G� >��>�����ܾ�ǡ�2@������������܉�>��>�Y	?��>,�U>G�>]o��{�&�ݾ�W �T�Y�����L3�B/�Gp�����@[��>���I������З>�%�M�>�_?��Q>��q>��>k��:YTo>W>�3[>�ߤ>��_>��">ݳ�=���`���DR?u���*�'�t��f���7:B?sld?��>��g�����=��D�?��?�s�?4v>��h��2+��Y?#M�>����d
?��9=z���ۈ<�b��o���ކ��p����>I׽d:�#�L�:f��g
?:(?�/��mu̾P׽�X�����=�	�?Ev?@�$�n�\�ͤx��{Z�Q�U��g��j��W�����A�c��n��$#�������7��ϼۛ.?Ɔ?�!�U��鉺���c�QR3����>�?�>ɽ�><��>�#>Y���&�)@]�v�(�1-|����>V�t?�`�>�F?�9?qO?ټR?ꘌ>&u�>����l��>.��i>(`�>w�?��)?�8?�.?��&?Z�d>� W�w���� ھ�?�?�o?|�?��?ԑ���Ƥ����*��@�����s�=��=1S����ꦹ<_�G>��?�z��8g+��\���>��a?�� ?\�X>���=�¾��>4�?��>�!�>�b������6#���/> �?N�Й��=��4��oN�Ieʽ�s>�{�=��;�`�+�1=��P;�$>'�>ŀ�<���< �Ӽ��=\iK���>H�?C؉>Wo�>: ��r �yA��ʺ=�N>yI>��>�Xپ ����6��=�d�S�z>R�?g&�?��u=��=���=����鼾���+M���P#=aI?��#?^�R?��?Go;?�} ?X'�=���6g���M������O�?��G?�?�>g�����TĿ�&�{x+?�S2?c��s�O>�畾�7��>o=֑���N�p�%����ާ&��?\����.�"�ʺ�?.��?@ۓ=��4�G���ߒ�S.Ͻ	�<?7D�=�/�>O�6?ѴF�4�	��������.y�>l�F?��>S�N?�}?��^?v�L>f�6�*�������|Q���><�9?#�~?2��?�
z?q0�>��">S(��$Ҿ���2�e"սS�y��7+=&V>��>-��>�S�>���=�|ҽ�aƽ93��x�=��d>X��>��>���>�ex>:�<�9?$��>	Kվ�^��߬�=ϔ��O>l�}?5�d?�$3?��>5t&������3>t��?��?�?#?���K��=J�����ٽ�����>$�>��>7�>���=\�>a �>�-�>�聾�8���F�? �'�?��4?:��=�qʿ�샿ޢ��!¾�e=�br�D�]��@׽����g�>{{R�J��-6ɾ>L�i�Ⱦ��Ҿ�c���2`�Uf���?��<=��>6~�=���b~a=�r�����sAh���<����7�O�(<m��=י�<�{��w��E��=�����@˾X?}?I?#�+?8�C?��z>��>�y6�?��>q����$?7V>I�T�UE���;�;���h񔾞�ؾt�־k�c����V(>W.F�?�>�d3>L��= �<%%�=j	t=h��=�xR��a=�U�=���=E,�=<��=O>�c>�6w?<�������4Q��Z罉�:?q9�>�|�=��ƾf@?+�>>�2������}b��-?f��?�T�?�?�ti��d�>���D⎽�r�=����)>2>V��=��2�̣�>j�J>����J������l4�?��@��??�ዿ��Ͽ�a/>��>��T>�z��FG�[���I�c'=(�U?�k�)b���P?�� �x�߾16�����c">J�.>`��Fy�#̳=�5�+=�=���=4�>��b>G;>*<$��0�=��>4.�='�=lAż?N��b�&��=���=�5c>�>>84�>�[)?��a?;3O?�0�>�Ғ�D��yۥ�R8<>켆�R¼�
>Z�>��>Ԗ6?�Q?��X?y$?�'>��j>�&�>�t��/q�́�f$�:��<��.?�"L?�A4>�ʈ=X� �}\,��A'���%���?x.?��?���>�����l12�0jK�[����]d�I ڽ�|���=y=?%���{��%M>CO��>�����>�>��9>B��>I8g>�>Rm�=���>�<��6�w"�=4�H=oQ>�7>~�3R����,=�S�2� ��<��d�lZ�����N��;�=���>V�>���>�X�=�"��s�0>ǔ�h�L�3��=��.>B�%tb�YM~�u�.�ՠ5�v4B>��W>�4��
���k�?e�W>L�?>^��?d�t?v�!>\�ʣҾd�����d��P��{�=��>��<�A4;�{y_�6�M�/�Ѿu�>{��>L�>�s�>J�F�)hC��=�^���XF�m��>���޼-�/�=�r���t�������`�5I�!w?����M�">kPj?��P?�?�¯>�m����ھtMi>�������=Jʾy\y�' >Z?��	?��?�c��:�D���ɾi)���'�>F�N��LP�{�����0�kT��۵���Я>L��� оy�2�ǅ������vC���x�J��>2M?�(�?z�b�n���8�O�jb��r�Ӄ?�,j?lk�>�i?�?����.�󀾖i�=[xo?Ȃ�?�$�?��
>,c>�\�ܥ�>��?��?n�?��)?�d��9?e���y�<���=�ݽfӄ>1O=�\�<c��>ib>�k#?��E⾇%޾X<��N0�W=�=��+>��|>*��>��>P�=�!�>�n,>��=��*>8�+����=>��h=J�}�o5 �-?U]/>��>I�$?>}��=�� ���=Pܳ��:���et���нN�N��n�=�i����:m$����>#@�����?fZ�>�̾��?ٚ�k�#M�>��P>|���k�>3�:>}ͅ>�!�>ϔ�>�w�kgI>��#>��˾�
8>s���#�ߑ?�K\�J��:`>�����01�~1��h����E�����u �Q�t�����G�>��"F�?8m�Ҵz��>*��[B���?ʍ�>�E?vK����H�� D>1��>rl>!&��0���=}���PӾm��?�8�?��d>�d�>|�U?=�?��H�1�J&X��`o��:�@f�Bpa�1r��l��w��X�n�T�`?�v|?ſB?��=�{>W=}?�j%��P��{�>��0���7����<���>�Z����I���n�¾����>>9ar?�,~?�%?�0U�ɉ�;\�=9�?��.?<�r?��I?�? �����%?�W�=W�?��?%�>V8I?,��>��=o�="y:�@��='Ȝ�	Ә�j���1�� ����=��<��G<�=!�=�Ņ=1s�<x��^����'$=�/=j]=�.	>0�9>7��>hd?��?�jq>7?jވ��&�IC���(?���z���o�nz��������%>�x? �?�O�?�@�>���i�c����<�,>s��>~*�>:��>t�=A�=���g>^��>���<��<`���]ɾ�%�����:B9��2P>B��>i|>H��r+>yw��aYv��c>2P��	����Y�	�G�E�1���t�ql�>
RK?*?z��=���	��(e�/>(?�;?
�L?]i?�ڔ=F�ھ�9�	J��e���>���<�:��$�������:�Hw�;��n>P���Р�h@b>����}޾ْn��I�t��%vM=�y��V=����վkC����=�
><���M� ����GҪ�0J?�	j=^���aU�os��	�>���>1ή>:�:���v��@�����I%�=F��>�;>\����wG�Z<�y3�>�GE?J�_?T}�?�K����r���B�@6��b���˼�t?8B�>�?ҶC>~˰= e�����`�d�J,G�C��>�#�>���I�G��c��+�����$���>��?�� >�r?��R?C�
?|`?�M*?��?@�>d(��e��$&?\��?>q�=<�ӽR�T�*�8���E�fG�>�q)?لB����>�S?O�?��&?9�Q?U�?��> � ��K@��'�>O�>u�W�Uc��t�`>%�J?J�>%AY?�у?�.>>�N5��Ƣ�{Ъ�ȑ�=_�>��2?Ł#?��?���>�L�>��Ҿ��˽^6�>�k?҅?�W?$����>�`ܻw��>bk>�v�>�3�><��>)4M?��j?��?dI�>��l�W;��C)���>R�A[��
>�</�;-��;�.�=�V$�d���.�<�h�=�������Q�U�*���v!G=�`�=��>N�>��h�E�o>�I˾xd���>>����m0��0�����r�o��=Bv�>�?0��>(��:Mp=E{�>L��>����N,?��>c�?��K� :h�'���%[�T�>_�K?}.�=�%n�e����o�H�y=��d?��]?��޺�N�b?��]?Ah��=��þw�b����f�O?=�
?3�G���>��~?e�q?T��>�e�*:n�)��Db���j�*Ѷ=Zr�>LX�T�d��?�>o�7?�N�>/�b> %�=iu۾�w��q��f?��?�?���?+*>��n�Z4��Q�co����[?ڎ�>c����$?R?�a�ξ�C����9qݾ�­�oY��'���I᫾�O-�쯋��ű�i1�=@V?��{?��w?B<_?��e�3�a�_{���[�$�����%�D��?�uHI�Ϗr�mH�5W��\����<�=�f�����?��=?;�i�q[�>�o�Xq������<.�Ծ�d����>:oR>{'�=N'>�p��o<�-]��?A`?k��>{D?��Y�~�W��l6���b��=/���`>�@�=g	�>�?���=�K1>(�r�.I��������Ž5v>pc?��K?��n?j1�B)1������!��.��M��}�B>@�>�y�>��W��|� ?&�G=>�E�r����������	��=��2?QO�>�͜>cH�?��?
i	�$^����x���1��E�<��>2�h?�G�>�͆>�kн�� �叧>3F�?:`?�ɬ>.�v��<�`�� ��L�>��?Ý/?li>g���/�;��#m�}떿O ����>���?q����p����>�I?>�=̬�=���>�U�pa�����(�>�ئ>���<㗩=���4Ĵ�̭Q�}ٞ�\'?���> L��$46����>( 7?m��>x�>�v?�n�>Ȥᾌ��='�?X]U?�2?��@?���>��d��O��i-�b�<ء�>.~U>��=7e�=����`{�#�S�^ ��_=<��=���eļ��|�f�q�q�=	W>y�ܿ�L��6��ŀ��xھ��ǾF��=�ؽ�*���������ߜ���뎾������.�<���u�¾ӷQ�Py���?/�@�e�!:��"��U���_�%��/�>�Ӿ�ى�1�_��'����p��4쾭1��z��Ϡz���'?g����ǿ���L;ܾ#! ?$B ?f�y?#��"�,�8� � >vH�<�.��%��X�����οt���K�^?r��>��-�����>���>��X>�Iq>f��g螾A:�<t�?7�-?r��>�r���ɿR���?ͤ<���?�@Y�=?��+�e���/=���>Kj?�;C>��)�-�ͩ���(�>;u�?wa�?�=�U���%���`?�ȣ���?��!��� �=�Ŧ=H�*=�f�H`>>��>M:�vsI�5e��V,>��s>����o�yS�"X�<�Q>���61���݄?'W\�f�|�/�$b���	>U?�S�>�Z�=��,?��G��qϿS�\�N�`?��?��?��(?ӿ��r�>��ܾ�bM?�?6?�.�>Z&�B�t����=G��G���R^�:HV����=���>@>��,��n��qO�kU��HF�=��x�ƿ|�$������=��غ[�[�i���m����T��$���eo�{�轠�h=I��=�pQ>@n�>y'W>�8Z>�aW?f�k?_A�>+r>�2��o��fξ`��;�����������"�@�l�߾x	�=��z����ɾ�6��G�=�� ��Vx�z:&���R�ho��@'?��:�������$�ߘ��+�Xq�%��R�w�G�Qxv��÷?8�m?����S��KG�*g���N׽B|?�}�*���>����=��>��?=c�>)�>tJ׾U�O��t���)?,�?�<���ꍾ�c+>i�[v.�}<$?��?N"}<3�>m)?��N��o󽉯g>9��=�X�>��>P�)>W7����B?��S?uF��É���>\a�����N�.=��>��
�M�H���\>�û�}�u^üg6ҽ���<�V?��>�f)�����᏾��&�S�.=�x?��?aџ>XTk??+C?	�<?���S�����Y~=/X?00i?�>����QϾ�~����5?-�e?<�P>�i�3�$�.����E�?��n?�/?3o��N�|��ݒ�U"�
<6?��v?s^�ws�����6�V�n=�>�[�>���>��9��k�>�>?�#��G������sY4�#Þ?��@}��?��;<����=�;?e\�>��O��>ƾ�z������
�q=�"�>���vev����R,�a�8?ܠ�?���>���������=���hs�?86�?+ͪ�]�b<����Bl������ގ<�7�=;�����뾑�6���ž�
���ڼ~X�>@@���4��>w�9�q$��$Ͽ�V����ҾRFn��?�>�����u����h��eu�WG�ĨG�%q����>	5s>�/�3���3i�� *D�8Z �,?Z{x���-=���<�޾Aѽz��)��=��?"��n��^��j��?�Zʾ0p����.V$�ކF?V��?oz�?�(�>�KM>m0�gCžQ=��K?$`�?y?��j=����V���%�j?�_��xU`���4�tHE��U>�"3?�B�>S�-�a�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���H�!�B0=�UҒ���
?V~0?{�f.�\�_?+�a�M�p���-�|�ƽ�ۡ>��0��e\�N�����Xe����@y����?M^�?h�?ѵ�� #�e6%?�>c����8Ǿ��<���>�(�>*N>kH_���u>����:�i	>���?�~�?Pj?���� ����U>�}?&ٶ>��?���=K[�>2�=����:���">D=�=�B>��?��M?^i�>[��=�u8�Q/���E��Q����,�C�e��>��a?~�L?_�c>����	P-��� ��Mͽ�m1��4�!�?���*�c߽p>4>_�>>T�>��E���Ҿ�u?�N�I`ؿL[��e=$��?4?��>	c?��Q}t����8B_?�1�>���ݳ�2Ջ�HE�(�?���?�&	?ܮؾ�	ۼ�h>��>�Є>��ս�˝�m`��ȋ6>}B?�T�y����o�,��>���?��@bB�?�ii��T?��4�����)���;�"���=�q2?x�� �r>��>m`�=�Zw��S���1p�_��>-!�?Z�?�e�>��l?�#q�|"A�j�[<cX�>��j?4?���;����;�:>��?��	���� ����g?,�	@i@��W?�����bֿ��U��ɘ��0=�={'�=�~2>Xڽ(��=]�7=�8�q�����=��>g�d>U�p>8#O>"\;>��)>E��L�!�_s��T�����C�s��}�n�Z�}��_v�p�a*�������S��r�½�8��O�P�8&�L�`����=��U?4�Q?�p?�n ?�x���>�)��H=�`#��l�=�>B2?�{L?��*?��=X�����d��[��sw��е���.�>ծH>���>�R�>]\�>���9�J>�M?>ې�>�� >�%=�����==�O>�Ϋ>���>�>5ŧ>tV>�ʸ�����B���E�k���=��??<	�w�B��XP�OB׾s�0��
x<a%??и>V���I�ƿg��J�L?��*�!��h~X="�<?xU{?�l�<�2���<�=CY>����q���QW>Z��;`���{־��>��?���>�|>��9�nP�1�f�m��2#�>�1B?���� � ��=B�8yM�����t��=X3�>㛽=����������Ie�_�,<��:?��?b2۽�'۾�e��Gʾ�n>ô�>�G��m�>BR>�\N����� 8D����=�{�=1no>���>���>�@>4�>������5�>6>��g>'@?��+?0�;��U�f=��I���=���>&C�>G5e>c�L��\�: ��>�4>yh|���>�!�$��T�>�H�����`�J��;`�����4>콱=�f���S���r��~?���(䈿�뾸d���lD?P+?I �=ΝF<��"�E ���H��A�?o�@m�?��	�آV�:�?�@�?-��:��=}�>׫>�ξ�L�ޱ?��Ž9Ǣ�Ɣ	�)#�eS�?��?}�/�Wʋ�9l��6> _%?�Ӿkg�>�x�LZ��H��W�u�N�#=Ш�>�7H?�T�� �O�/>�w
?�?.^���k�ȿ�{v�k��>#�?b��?u�m��A���@�0��>���?�fY?�ni>�h۾�`Z�=��>k�@?�R?M�>�8�<�'�n�?m޶?N��?��B>�.�?��s?��>lp��(0�Q���������=�y=J�>yX�=Q�žңD�h���K���}�b�����ew>B* =�5�>ab�q��qs�=�I��?����
�q÷>#(d>�U>S��>���>��>�>E��<�6����t��'��dL?���?���@n���<���=�:^�h9? 4?%�[��ϾR��>�\?Y��?�[?c��>���I:��;迿�n���X�<��K>��>	2�>:I��~K>վ�D����>���>q���Gھ�<���~����>Ho!?N��>v�=4� ?
�#?=�j>�>RE�#8����E�a��>��>�e?��~?J�?a湾�R3������㡿�v[��N>$y?�D?9��>r����x��IE�ɢI�u	��F��?p_g?��?�1�?uh??��A?�f>���j�׾�x����>]�&?N�D�7�E��{:�]�ʽ�?�?x��>��ӽ�sý[�?�	����'?��K?)�+?���1Z^�Z�ξ#n=�g����<�4�<"|��o*>H7>�hʽ!Ҏ=�>�d+���R��П�Xc�<�{=�.�>���=_���.��iR,?\F�z�����=��r��D��)�>��L>�C��3�^?uP=�0�{���� ���� U�.�?]��?V�?w޵���h�>=?8�?�4?�
�>M���I�޾)��w��Hx�����3>k�>��x���侉~��R���WI��I�Ž�;'��?/�>��?~��>�8,>,�>�/ٽ**����8��Y�U�&��18��� ��r���zC�h'��lɽ�ԾF����e->��)U�>$�?�)�>"�3>�t�>�/1;:ȁ>��3>}4T><?�>��#���O>x��>4P=����ZQ?}¾{(�o2�*쩾�@C?��c?���>�Or��O��@��\q ?
�?{n�?�|o>g��`)���?zR�>�ʀ�l�?3)3=�^���D<I8���k�]���{D*��V�>�@۽��9�e�L�&�o�5�
?��?�z���ƾB�˽����j�p=�{�?��(?��)��Q�!q�V�V�#�S��9@�6�d�����'�#��q� ~���4��y���J/)��m=[+-?�(�?+�����Բ��<m�Е?�1bm>U�>���>Lr�>4}H>vN��B1�~�]�s�$�t􄾧��>Y�w?�\>p�??\�??��N?�(F?%�<>`>����?b=�:q�>�
?�U?T�?V�'?�:�>\)?t�>4�p<�C�#;�z�?�?N�+?�t?O
?�_u�h�^'ۻ�=��y����<�%y=�V��a�H��σ�@e>�[?ֿ�8P��2ʾ} ?`v?��>��`>��
�s���(��m@?$�?gg?Hu�"-��Uc�e�=��?����=	>:�_>UuɻJ�V�}>�a\=��<[l�����=�z7�Y��=�O�=�h��O�<�Lb��稽��"=�f�>��%?@ߘ>Ij�>T����p��H��{=ڿ_>fO�>�`!>�SᾶH������3]�LvZ>J�?���?+c�=�K�=}�=�q��Huþ�Y��_�����<?�?/F?AM?���?��E?�?
�=�.�&#��`̀�գ���>?�M?.i�>pM���ʾp���]F�0�"?�5?~d����M=��� ZӾ��.>f����]�0W�'���!P�n@J���'�>�^����?�?���<I>1�ި+�|2���[@�7=? ��;q��>�;?D�"��"�[�.F���wu>OQB?Fn�>�P?�{?�f\?E1Q>��8�eU������A��g">�>>?F�?��?lcy?��>3�>��'��3ݾ�����i#��j���j�U=��W>f�>���>/)�>H��=��>C����@���={�`>s��>q��>�I�>VT|>���<G�F?}��>�Z��ږ��ݤ��H���1#�`ev?�Ώ?��*?\�=9����E��-��S��>�٧?f�?N�(?��V��U�=�!�B����t�z>�>]��>�ś>���=�I=�J>��>�D�>y��?�X�9���E�|�?�DE?$V�=�iÿ!{q�՜x��Ο�s^�<E����ge��}��QT�Z�=�i��2��Q����\��������I�������u�x�(G ?�P=�c�=��=Z�<�)w�h�<"�^=��<<��=O��\s{<
�<��Z����?�;c��<]M3=ٌ��("ƾ}�z?��J?`-?��:?�N>U%>M=��ģ>GA���?_/`>q��>>��;�,�s���$Q��̺�������o�����Y2�=Dƒ�@�->�IP>"m�=GT�A�>�=5=�׾<k0�ѳu=�7�=�d=���=��=,g>���=G5w?^���~����7Q��=�x�:?66�>�t�=~ƾb@?�>>�/������a��+?���?eT�?D�?�si��f�>���l܎�p�=�����D2>���=H�2�<��>O�J>��CI���j��+3�?�@]�??����:�Ͽ!T/>��R>�	�=��S��<�8��|���1��?46���þ�ŉ>�=������}M=�'Y>&�=��-��YW�(�=ڽvVh=�!B=� �>'XM>��=O<Ƚ��=Ա�=�'�=��L>q<���i@�e�Z=��=�J[>M�>���>�a,?.&R?�u?�*>;�ݾ,־�N��J�>ߒ�>|����!�Öd>c��>$�]?�"?<5&?�%	?��s>mJg>���>3����i�ً��p�¾���?��}?�8?e' >����ӛ:��I[��U�U��>f?�E?ѽ#?c���x鿻����2�ҩ��S7N�[���ib�e:>̞�=�?t�,���`;��p�>�><�
>�R�>!�>ޡm>^ǽ>MH\=FV꼀p�=B���]�>�ަ��J��&Q�=es�=�N�,/����v�$�=_i=��*>.�Z=�wQ=V�i=��=�f�>�a>}%�>DH�=؃��M].>X5���FL��q�=?ܦ��A�O�c��~��W.�z�6�1KB>��W>�W���"���~?b
Z>��?>h�?~&u?m( >��q�Ծ^��*$d���Q�)�=��>0d=�k8;�ګ_�ЎM���Ѿ��>�>m�>���>�Z8� @���=�ӾV?���>ov���`�������t��������R�y�����~�.?�i��?>���?lQ?7]�?���>ں���;��>����H�h=��>.���<N={�%?�n?J�>?�;Eg8��?̾8��]��>leI���O�������0�Q��b���x�>�ު���о�"3�$b��������B��Ar�]ں>��O?��?[b�qW��cbO���������f?�yg?|��>6>?B?�硽���w����=��n?m��?�+�?��
>�n="����>58�>�ړ?�?_QQ?�p�]�>:��sm�=+?�=�>v'>�	P�<��>�2�>5?��n�+��i��C���-5�+m�=q=x�7>n��=ۯ>��	>I��<aہ��u�=��><$�>ci>��>ҜB>4���O�����>�$:<�j�>�$4?��>�aW=@�G=x������� ?��Y��-�.���l�ԏ>	>�� �V�����>�����>�?[3�=
�׈
?�)ξ�Y�1zV>��e<�a3�>d�=���>C�>:��>ko�:�B/>��yFӾȀ>z���d!��,C�i�R���Ѿ|z>G����&�����y���BI�Kn��8g�nj� .���;=��ڽ<�G�?a�����k�&�)�%���0�?�[�>�6?�ڌ��
����>i��>XǍ>=K��e���hȍ��g�t�?��?�"c>
3�>k�W?��?��1��c3��{Z�$�u���@���d�Ġ`��Ս�(���	�
�����_?��x?z�A?��<�&z>���?��%�Z׏���>/��,;��g==$@�>�4��T�`�T�Ӿ(�þf-�k�F>�so?-�?�T?�CV�Ld��>1�7?`�/?Ʉt?�}2?[�:?Xc���"?͖*>��?Cw?1~4?�.?��	?��4>�v�="d��N,=yn��4e��_Mӽ��ɽ0����w1=#�u=}�Ż��#<��=\U~<S��GӼ-&��A���+"�<W9='�=YC�=b>Cp]?�?j�M>�| ?R�Ӿq�c�c��kP?� �>�@�Z`7�v��iOʾ[��>�Z�>?�?���?���>esM�p;g��d�;�q;=�>>ً>(x>k���i۽�;E�y�R>�Æ>��t=�+��Uׁ�2l�>���s�<�>���>�H�>+��<�ּ>��о�p��3I>G,&¾�;I�` D���7�R|"����>�n?rG?���w��Z<�\y����(?߾(?��?*�?��=>����F����ھpn����>e�,�sQ>��F���0���u(��s>�T�>�)���O����>������ؿi��R�v������<>��Ue�<���B����U�Y��=2�>�3Ѿ�_(�g�L+��B J?K��=�s��J�[�w�����=MT�>o9�>XP~�W|S���,��K�����<�d�>H>a�d�+���A��p�g>!I?��h?x�i?�K��Ɓ�.S�DU
�0A��u~��Ҁ?B��>��?��F>QC�=��Ѿ�$�o�s��Z��s�>4?W��aA��՞�H� �A�,H�>�B�>H�>��?ܻE?�;�>��b?��?Ka�>݈�>駾�W~��A�$?`u�?�U�=��'�_���9�	�=��V�>�k!?�3���>��?ʝ ?a�!?�L?�|?�  >�����C�*��>���>�>Z�B󰿻 �>�H?m�>�}Y?ۂ?��=>�2�@L���,׽�>m��=)�0?�;,?�M?2��>-��>Gڟ��~�=/@�>�.d?�t�?�_?l�=D?�S�=���>wk=��r>+��>�?�~Q?�xm?��<?��>�{�<�-���?���U��n�:���k<vB�r�=1M�0����V;�$�<X�<oy^�����q���7���b�j(�<�=�>�u>�^��*�1>biľ�{���?>X����́���@<�b��=M7�>�?F�>H� �"�=M�>���>�p��d(?}U?�v?_�;/�b��ھ��L��>A?���=��l�#��
�t�UMg=jAn?�b^?��R�Y���=�b?��]?�g�=���þ��b�ډ�Y�O?4�
?��G���>��~?M�q?.��>'�e�
:n����Cb���j��ж=r�>4X�d�d��?�>��7?�N�>��b>�$�=[u۾&�w�fq��d?f�?�?���?�+*>��n�[4�O<��il���]?ð�>F����"?J�+��/Ѿ�+���\��?�⾠���̫����m���ԫ$���)ؽ;�=�i?��s?W�q?o�_?� ��Rd��~^�6��d�V�eq�����iE�E�C���C���m��C���J�����1=� ���&�X,�?	4C?^�7����>�j��LKپ����U%=>����lm�i�`>:�U=�<>eIr=x��}[u��̾�?�??P�@?��c��]X�<D��E�����̈�Ar3>���>��1?���>Eb�=��$<�@��y�d=����@�x>�lc?K?�o?B��~u1�����6 �9�L�������G>�)>��>!`�oK��c%���=���q�����J��Y'�r=ă1?���>1��>���?=�?K��-W����s��4/�n=<*�>��f?���>�@�>\2ƽ\8!����>Rwj?Wi�>��>2:��j��3�y���ѽ�|�>S(�>8��>�0l>��#�x�T�SX��壊�R=/�c�>�o?6)��倾wa�> �H?&,="�=��>��u�����۾�A0�lK>\�?h��=>>D;ǾO���%��R鑾�_ ?�d?�F���_��S�>�)?�a�>���>E�?��>y��W���7�>>\?�]R?�TM?^"�>�v=C�,�Z���f5�8�=�~�>t�_>!��=2'@=�����ig�d�$��M=
>�<@B�����䀚���;$�k=���<�f!>5[ѿ��S��������������d��e�n�r�P�C�	�Q�yr`�t6�n���P�=�s-�����M1��o�|��c�?4��?)Ƚp,m�nȍ�@@��]�����>�����O��о�޽<ܽ��
��~�bG��B�P��u|�:u��S�'?�����ǿ󰡿�:ܾ1! ?�A ?A�y?��1�"���8�� >�B�<�,����뾪����οA�����^?���>��/��q��>Υ�>�X>�Hq>����螾�1�<��?.�-?	��>Ǝr�/�ɿ]���hä<���?,�@�:>?��#�*��㚖=�\�>��?Q�+><�)�	F�������>���?뺅?|[�=ϥU�u�!��6b?�	�E$<��a!�̣�=���=4�<�����I>�,�>I�<���J�@0a��u>rK�>Z��ȵ�EJZ�4D��6DA>���KI��4Մ?+{\��f���/��T��
U>��T?�*�>]:�=��,?Z7H�`}Ͽ�\��*a?�0�?���?$�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�ԅ�=i6�Z���|���&V�m��=Z��>j�>ǂ,�ދ���O��I��Q��=�����˿Ź#���$�y)�<�~=�	��DJ��r�;ܹ�=�5��������.��=��=�{�=��->�i>S�q>�]?^`^?u�>q�V>�D�p�g��*���B��G�O���;�1#���M���˾�\�F績��[��� ���<�B��=�Q�����x� ���b���F���.?Ys#>�ʾѧM�ؑ9<?�ɾ����u���N��~�̾�1�}An�u˟?hB??�����V���a���?��1�W?K����1����=͐����=#��>���=��⾔�2��fS�@x%?�7 ?2Ȭ�a#���R�>e����R=�/?j��>����D$>��?4�b� ��7e>��H=��`>�[�>mW>������u?�l?���=��P�H�>79ž:���>:�=Ya߻���1;���>LH>��W�����m=���=U?���>�Q(��	�;䊾Sj'���r=�^x?z1�>R��>��e?��;?��<;����R��N�Ɏ=��V?�c?f�>���EҾ�š�=^6?L�d?$5X>�JW�̚־�V*�-����?/�e?� ?8��	�~�J���%���R6?�w?�]�q����V�d�\�z��>P��>�K�>+�:���>�d??��'��
�������5��~�?�_@M��?� <ei �E�=x�?���>�P�x�ƾ�x���ϵ�Fx=�k�>�ը��7v�v��P�1��8?㜃?��>Sc��!��e�=�;r�j�?��j?ƻ��r�ɽ)0��u�30���ܼ�6���H=b�=M��f��������#�3uҾ,�	�̆�>@�G���z�>~��0'�i�¿�m��)��d���?HO�>$���؏���c�@{�%�I��WU��ݾs��>�>��t�j�냿WT��ᅽ��?tފ��F><�m=P�¾�҅���"�B%>��>>)Yu=1�~�Ͷ��+�?��徠A߿�%����D���i??	ԣ?#��>0�>�p=���1���/X ?&?Ik?~\�>�T=Ă��i�j?�^���U`�;�4��IE�	U>�#3?�D�>G�-�H�|=�!>L��>�e>,$/���Ŀ�ض��������?��?jo�@��>���?hs+?mi��7���[����*��)�S=A?�
2>k���+�!�U1=��ђ��
?n}0?{�4-���_?C�a�O�p���-�
�ƽ�ܡ>��0�Gf\��-��]��rYe�����Cy�U��?<^�?��?��8 #�36%?6�>�����6Ǿ,�<���>()�>�%N>�C_�T�u>����:�sc	>��?}~�?�h?��������"V>��}?V-�>��?���=���>���=-�����'�"M$>��=G>�L=?�^M?���>���=��8��4/��IF��R�0��ͰC�X��>l�a?	�L?��c>�&���0��!�l�ɽf�0����G@��1��ݽ�J6>�H>>�[>�wE��aҾ�?p�E�ؿ
j��Nq'�{54?w��>b�?X���t����~;_?z�>�6��+���%��BB�A��?kG�?>�?��׾�S̼>��>J�>6�Խ��������*�7>1�B?���D��\�o� �>���?�@�ծ?[i�U	?)��T��'f~���A7����=�7?�E�[�z>���>���=�kv�"����s�z��>�?�?u�?R��>&�l?o��B��	2=�8�>�k?%{?��o����B>r�?��I���)J��f?��
@bt@�^?�뢿��ؿ`����;��޾">��p��=��F��
�=~"�>m>��=��=�J>�>���>��E>8!>�1;>+�������ٓ�,kM�y��]���Q������p'���[�W�(uݾT�^�&��3����@�O�8�r����=�ZT?$�P?��o?o?^�_��O>�����=vo$�?!�=��>e1?�}M?�*?�*�=uf��v�e�I��������=���y�>݃F>���>���>	�>���I>bLA>^ځ>�k>�*=�?F�?�=N>I-�>��>�b�>�gV>9�,>�p��Ḳ�Нo��n}����v~�?�r���$D�[<��?#���n���`�=+&?V��=3(��S�̿����ĴH?[Ɨ�o��[M&��!�=25?�)_?�+>�G��{ ׼\p.>L.��j����=���SM������f>=i?��g>Q�o>�2���4��N�%��Ȟ�>17?林�R�,�,�r��1K�"�߾\�B>��>]���/��Z_��z�}�/&d��E =�[<?��?�}��Nr��$|��I�����f>�wY>3;�<?ϩ=U�E>�EJ��?��$;D�6zC<t��=mf>ة�>��8>kM�;���>����n�$�v��>��>�6	>�Y:?$?���n̽���������l>T^�>�	T>�y|=1�5���5U�>�bx>Rq�;��\��|B��!P��"�>,���+���v�̥�����+�>|�=Z��|�k����=�~?���䈿��Oe���lD?I+? �=�F<��"�D ���H��J�?q�@m�?��	��V�K�?�@�?�
����=}�>׫>�ξC�L�Ա?/�Ž7Ǣ�̔	�D)#�dS�?��?��/�Rʋ� l��6>_%?ѰӾ\h�>Sx��Z�������u���#=P��>�8H?�V����O�#>��v
?�?�^�ݩ����ȿ1|v����>I�?���?d�m��A���@�g��>:��?�gY?�oi>�g۾`Z����>��@?�R?�>�9�J�'���?�޶?ϯ�?��G>9��?��s?��>�x�H�/��P��E���g�t=>�:k��>��>�����E�fl���z��6"k�J��8^]>��)=��>����U��?.�=>�����`���>��p>4DL>aW�>q��>���>ט�>�=��� ��������K?���?���*3n�4�<���=�^��'?eH4?�][���ϾԨ>[�\?>?([?�c�>���>��P迿�}��f��<��K>!4�>bG�>j!���HK>��ԾI6D��p�>ZЗ>x���?ھ�,�����yB�>�e!?��>�Ю=� ?^�#?�k>�U�>IE��-����E���>���>�M?��~?��?4����I3����?ۡ��u[�o}N>�y?RK?ˈ�>�����{����>�#GE��B����?-]g?R�佋�?�+�?�??-�A?-f>����׾����'��>�D?P���5�jQ��\P���?d	?���>2�Y=�xz�Mq�W����
��O?As?}�+?C���SjM��h���^=�a<VPx=^��=��g�tI>��_=3���t3!=�!�=�ĵ�s9����&���=�h�<?��>P�0>(z������.?�[һ����$}={w�c8C�Z��>^^>֍ʾ]�`?m*�R������Sٝ��rg���?���?�f�?iν*�f���:?���?!]?l�>ˉ��������T?h�w�f�`�G� >��>�����ܾ�ǡ�2@������������܉�>��>�Y	?��>,�U>G�>]o��{�&�ݾ�W �T�Y�����L3�B/�Gp�����@[��>���I������З>�%�M�>�_?��Q>��q>��>k��:YTo>W>�3[>�ߤ>��_>��">ݳ�=���`���DR?u���*�'�t��f���7:B?sld?��>��g�����=��D�?��?�s�?4v>��h��2+��Y?#M�>����d
?��9=z���ۈ<�b��o���ކ��p����>I׽d:�#�L�:f��g
?:(?�/��mu̾P׽�X�����=�	�?Ev?@�$�n�\�ͤx��{Z�Q�U��g��j��W�����A�c��n��$#�������7��ϼۛ.?Ɔ?�!�U��鉺���c�QR3����>�?�>ɽ�><��>�#>Y���&�)@]�v�(�1-|����>V�t?�`�>�F?�9?qO?ټR?ꘌ>&u�>����l��>.��i>(`�>w�?��)?�8?�.?��&?Z�d>� W�w���� ھ�?�?�o?|�?��?ԑ���Ƥ����*��@�����s�=��=1S����ꦹ<_�G>��?�z��8g+��\���>��a?�� ?\�X>���=�¾��>4�?��>�!�>�b������6#���/> �?N�Й��=��4��oN�Ieʽ�s>�{�=��;�`�+�1=��P;�$>'�>ŀ�<���< �Ӽ��=\iK���>H�?C؉>Wo�>: ��r �yA��ʺ=�N>yI>��>�Xپ ����6��=�d�S�z>R�?g&�?��u=��=���=����鼾���+M���P#=aI?��#?^�R?��?Go;?�} ?X'�=���6g���M������O�?��G?�?�>g�����TĿ�&�{x+?�S2?c��s�O>�畾�7��>o=֑���N�p�%����ާ&��?\����.�"�ʺ�?.��?@ۓ=��4�G���ߒ�S.Ͻ	�<?7D�=�/�>O�6?ѴF�4�	��������.y�>l�F?��>S�N?�}?��^?v�L>f�6�*�������|Q���><�9?#�~?2��?�
z?q0�>��">S(��$Ҿ���2�e"սS�y��7+=&V>��>-��>�S�>���=�|ҽ�aƽ93��x�=��d>X��>��>���>�ex>:�<�9?$��>	Kվ�^��߬�=ϔ��O>l�}?5�d?�$3?��>5t&������3>t��?��?�?#?���K��=J�����ٽ�����>$�>��>7�>���=\�>a �>�-�>�聾�8���F�? �'�?��4?:��=�qʿ�샿ޢ��!¾�e=�br�D�]��@׽����g�>{{R�J��-6ɾ>L�i�Ⱦ��Ҿ�c���2`�Uf���?��<=��>6~�=���b~a=�r�����sAh���<����7�O�(<m��=י�<�{��w��E��=�����@˾X?}?I?#�+?8�C?��z>��>�y6�?��>q����$?7V>I�T�UE���;�;���h񔾞�ؾt�־k�c����V(>W.F�?�>�d3>L��= �<%%�=j	t=h��=�xR��a=�U�=���=E,�=<��=O>�c>�6w?<�������4Q��Z罉�:?q9�>�|�=��ƾf@?+�>>�2������}b��-?f��?�T�?�?�ti��d�>���D⎽�r�=����)>2>V��=��2�̣�>j�J>����J������l4�?��@��??�ዿ��Ͽ�a/>��>��T>�z��FG�[���I�c'=(�U?�k�)b���P?�� �x�߾16�����c">J�.>`��Fy�#̳=�5�+=�=���=4�>��b>G;>*<$��0�=��>4.�='�=lAż?N��b�&��=���=�5c>�>>84�>�[)?��a?;3O?�0�>�Ғ�D��yۥ�R8<>켆�R¼�
>Z�>��>Ԗ6?�Q?��X?y$?�'>��j>�&�>�t��/q�́�f$�:��<��.?�"L?�A4>�ʈ=X� �}\,��A'���%���?x.?��?���>�����l12�0jK�[����]d�I ڽ�|���=y=?%���{��%M>CO��>�����>�>��9>B��>I8g>�>Rm�=���>�<��6�w"�=4�H=oQ>�7>~�3R����,=�S�2� ��<��d�lZ�����N��;�=���>V�>���>�X�=�"��s�0>ǔ�h�L�3��=��.>B�%tb�YM~�u�.�ՠ5�v4B>��W>�4��
���k�?e�W>L�?>^��?d�t?v�!>\�ʣҾd�����d��P��{�=��>��<�A4;�{y_�6�M�/�Ѿu�>{��>L�>�s�>J�F�)hC��=�^���XF�m��>���޼-�/�=�r���t�������`�5I�!w?����M�">kPj?��P?�?�¯>�m����ھtMi>�������=Jʾy\y�' >Z?��	?��?�c��:�D���ɾi)���'�>F�N��LP�{�����0�kT��۵���Я>L��� оy�2�ǅ������vC���x�J��>2M?�(�?z�b�n���8�O�jb��r�Ӄ?�,j?lk�>�i?�?����.�󀾖i�=[xo?Ȃ�?�$�?��
>,c>�\�ܥ�>��?��?n�?��)?�d��9?e���y�<���=�ݽfӄ>1O=�\�<c��>ib>�k#?��E⾇%޾X<��N0�W=�=��+>��|>*��>��>P�=�!�>�n,>��=��*>8�+����=>��h=J�}�o5 �-?U]/>��>I�$?>}��=�� ���=Pܳ��:���et���нN�N��n�=�i����:m$����>#@�����?fZ�>�̾��?ٚ�k�#M�>��P>|���k�>3�:>}ͅ>�!�>ϔ�>�w�kgI>��#>��˾�
8>s���#�ߑ?�K\�J��:`>�����01�~1��h����E�����u �Q�t�����G�>��"F�?8m�Ҵz��>*��[B���?ʍ�>�E?vK����H�� D>1��>rl>!&��0���=}���PӾm��?�8�?��d>�d�>|�U?=�?��H�1�J&X��`o��:�@f�Bpa�1r��l��w��X�n�T�`?�v|?ſB?��=�{>W=}?�j%��P��{�>��0���7����<���>�Z����I���n�¾����>>9ar?�,~?�%?�0U�ɉ�;\�=9�?��.?<�r?��I?�? �����%?�W�=W�?��?%�>V8I?,��>��=o�="y:�@��='Ȝ�	Ә�j���1�� ����=��<��G<�=!�=�Ņ=1s�<x��^����'$=�/=j]=�.	>0�9>7��>hd?��?�jq>7?jވ��&�IC���(?���z���o�nz��������%>�x? �?�O�?�@�>���i�c����<�,>s��>~*�>:��>t�=A�=���g>^��>���<��<`���]ɾ�%�����:B9��2P>B��>i|>H��r+>yw��aYv��c>2P��	����Y�	�G�E�1���t�ql�>
RK?*?z��=���	��(e�/>(?�;?
�L?]i?�ڔ=F�ھ�9�	J��e���>���<�:��$�������:�Hw�;��n>P���Ƞ�b>ߪ��m޾�n��J����'M=��FV=�#�b�վ��~�/��='�	>g���6� �����Ԫ�C/J?clj=u|��U�Γ���>xȘ>nخ>*K;�O�v���@�;���Ö=���>/';>4�����T�G� 2��ɞ>�2R?^�^?'�l?�^y�bgt�5ET����y��x)W�cJ+?'�>�?t}>��<����KZ[���4���>u�? �?W<�좘��6�ti2���o>��?]x
>;?UEf?cK?��u? W0?V�?��>��� s�*�?평?�ۆ>l����Ƅ���*���@��?Q)5?�xɾi�>�#?��?^S-?��D?PR5?ܑ>*U��RD�ۇX>�ς>�=�+ζ�a��>!H?���>,c~?a9�?��Z>�����Ͼ/v���#��:�J?�(?�0?��>�>�d־��=�?V�q?<�?��?e�U����>D!�>,�?��p>�@ �^��>UzM?d#?�<?Mw?�ߑ>�z+<�;Y=,�o�]8�;ų�=�=$<�i��{yZ��]�
�L�)�D<n?
��V<ऽuE�;#�p�@P����c=a�>��s>������0>��ľoP����@>���^e��㊾�f:�隷=�>
�?�z�>g#�Y�=��>a�>����H(?��??m�$;��b��۾L�~�>v�A?��=��l��{��T�u�Nh=j�m?o|^?�W��8���_?8?q?�0��Y,<�<�¾�b��u^ �G�:?�U�>Gr��P��>+l�?�{�?sa?�2����O�-+���Q�k����n)=��>����mS�N�>8�"?d�>T�;>��P>}�ܾ�n��<��+:*?�ԕ?�د?ҭ�?e
�>�ml�ܗ߿ذ��|!��;�]?���>Y�����"?ϵ���Ͼ�犾�x���(��r���b��|G��E���OY%��w����ֽLӺ=�a?cNs?Z\q?�`?A.��	d�%<^�6��G�V����W�r�E�m�D�`�B�|�n����_���F��z`B=(�q���E�,�?}�%?a7:�r
�>�Z��� پ�	־�#>2!��|l �'+�=�؜�=O�<�$=�'n�j!�W��z?\�>��>�3?�[�� =�?�4��H8��|��9�@>��>u�>���>܈�;$�^��~}Ͼ�<��]Ľfߔ>��m?�V?�O?�K=��	5��|��%��<͆��o�����=">���>�j���S��	�e�(�S΂�3�*���������o�=�}H?���=���>��?��>D̾���fž�~#��뽂��>�e�?�T�>���>�*��������>�Yl?���>��>���ǋ!��z��RĽ'z�>�S�>��>� o>F[-��\����E���k59����=��h?wo��e_`�e�>�Q?B݊9�M<i�>!mu�O:"��1��n�)���	>��?l�=�=:>
�ž$:�p!{�������(?�d?G����*��}�>}>"?p�>v�>�;�?32�>$���������?�]?�aI?��B?��>f�=3���mY˽��'��(=Ȝ�>Z%^>x�n=���=&Q���]�:����B=�s�=Y����s<'�Լ��<Q��<sm4>�XͿ�O5��̴��V�Vr��-��*��7+��A\�qF*����.h��Y���g���A��q��2㵼<\��5������?��?Άa���&�Û��4����sR�>F��㦉<�̾���Ay�v�W˾,(R��z��Γ�>�Z��H0?�=����ӿ�J���)���^?�?�^?����"�Ғ%�X�->cѹ���i��,L��t�ͿI���i?y��>�޾&<��T�>�դ>�O>�,�>�uY�;n��5|=��
?��+?�?*����O̿,�����;�1�?C�
@3zA?��(���쾡(V=.��>�	?��?>҂0��Z��9��nL�>%(�?A�?�M=`�W�c�
��_e?��<��F��=ڻ���=��=E=���fJ>��>����UA���۽��4>�܅>�!����z^���<w0]>u(ֽ���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=r6��{���&V�}��=[��>c�>,������O��I��U��=di��yR����%��X�����W���x��~�Ǟ>z&���Ⱦ�Ȏ������}��=ÊZ>b7?��>	{|>;jb?��l?m!�>�ܫ>�T���H�Ѿ�!�6>��>�Z�s�վGS���F��Wྏt��Vz��߾ͯ����e�6�R<�=��G�xe���/��_� I��� ?���=fd����^���D��淾�＾�<�]n��i���h>�kj��ۧ?��8?k2��l�C���%����f$���`?��o�!����s�ǟ�=��ڽl��=.�e>��<���.�A��CA�B0?#�?r��\v���3,>c����=h�+?
�?%tm<p-�>Y�$?@})�n:�%0[>��7>ss�>�?�>�/>���<8۽�/?�sT?�^���蛾Mѐ>5���`f{��4j=�Q>M�4�����[>Ձ�<7ߌ�_�e�7���c��<�%W?�y�>��)�X��Ch��٪�[�==�x?n�?W�>_sk?��B?���<�i��!�S�$���v=��W?.i?�>uB��T�Ͼ딧���5?��e?ۤN>rh�\�龆�.��F�'$?��n?�\?�͜��o}�������dk6?��v?s^�rs�����$�V�g=�>�[�>���>��9��k�>�>?�#��G������cY4�Þ?��@���?9�;<��I��=�;?w\�>-�O��>ƾ�z������)�q=�"�>���`ev����R,�^�8?ՠ�?���>������3�;>vǘ��*�?��b?� ����O�d
��T0�rg#����ʀ�=��)�M��=,���"@�d/��+��V���D>�>�2@�鵽̸�>N�^�ҵΏ��3q��K���?�J�a�?"f�>r�D�~��x�L��eI�7�@�8�S�����b�>��>�C���ڑ��:|�0�;�vj�����>ǂ�xb�>T�U�N2��'��� /)<�.�>D,�>uq�>δ�{7��%�?������ο|_��r���W?:>�?���?��?�#,<�ds���z�P�?��sG?�r?e�Y?�[2���^�C�1�D�o?|��vs�7��FM��^>A�&?"z�>�F��%>��>>d��>���=�-��\ƿq���z��k�?��?�����>x2�?�+?t���`���&���!���=,�3?m��=G?Ծ���4i<�� ���1	?�3?�*��~��]�_?+�a�M�p���-���ƽ�ۡ>��0� f\�N�����Xe����@y����?N^�?i�?ֵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>^H_���u>����:�	i	>���?�~�?Pj?���� ����U>
�}?�-�>��?η�=2H�>��=� ���M2�2e#>Y��=!�?���?��M?*s�>���=_�8�/�9SF�:IR�Y-�~�C���>Q�a?�L?�b>���D�1��!��>ͽ�Y1� ���@�˵,���߽Qs5>�>>�;>R&E��Ӿ��?�t���ؿn���'�q*4?���>��?����t����5_?�r�>�?�O'��t ����&��?�B�?��?T�׾��̼>��>�V�>j�Խ���k{����7>�B?,���@���o�7	�>���?�@�Ӯ?�i��b�>�g��Ƈ����z��ĒE����=m�3?����nr>�
�>���=��o�����Tdk���>�ײ?	t�?
��>��m?�_�f@�m-�=�`�>D�n?��?Ml	������%>\��>~r�����Bh��X?�\@�h@�W\?7F�����5⤿�ۭ������=$+N;��	>a�H��}��|	�e�G��<��Z�>e�>� N>��>>��~>��8>t >���)� ������Φ��9C��F��4�]�p����Kjj�{t��*��b;���aCF=��+��N���7��~(��"�>�4[?'�Y?�Hi?��>�4
��MX=����\�=�5��p�=�Q�>�o'?"\?�H.?9�>����r����1�]�G�>�;>Pl�>k��>�%�>Mk�=j�H>��=��>~��=�=j�����z��B�e>
?�>��?��>�D<>+�>fϴ��1��E�h�;w��̽� �?D���V�J��1���9������`h�=a.?[w>���4?п����3H?�����+��+��>-�0?�cW?��>N����T�Y@>�����j��a>H1 ��~l�R�)� %Q>�m?�f>�u>R�3�tC8���P�������|>K@6?�-����9�k�u�A�H��Gݾ��L>�Z�>K�M�|�������~�j�i�)�z=Qb:?�t?�����԰�"Gu�9.��KHR>+\>U�=5��=ѴM>bOb�Ieƽ��G��.=�=��^>�?�*>/��=�c�>s�� �L����>`A>#�->I�@?x%?����Ξ��)���(�0�w>p?�>���>"'>��I�&�=4�>"�a>���~��/�cB��W>�~�y]��f���=�w�����=��=_�wR=�`�&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�f�>����S��������u��<#=���>�RH?�����R�Ds>�AG
?�?nr������ȿ�uv����>g��?�?��m����@�RX�>���?�:Y?�i>�F۾{�Z�?��>��@?�R?�
�>��m'���?oֶ?ū�?�op>�1�?�+p?U�>��x���2��˵�8���VF�7���*'�>�	>e����?G�Dr�������bq���	am>J�$=�|�>K{�y���`M�=�6	�I�о������>�Jk>=�>���>�h?���>K��>�ҿ=(M���c��׿��gK?ҽ�?���I[i�6\<cMo=�u����>�1?�6Ӽ��Ѿ!_�>�3_?<G�?x�X?��>G��Y䜿�'��X\���)P<��I>C��>#�>�(���ZT>PԾ��1�qȅ>p��>��b�z`㾣�|�<]�<㙟>� ?���>���=�� ?^�#?�
k><��>�.E�~0��-F�Mu�>��> ?"�~?X�?�k���m3����ϡ��[�/aM>�x? 1?���>�G��X��0D;��\O��^��&_�?рg?8s�k<?]�?�??-�A?�f>�-��X׾���>��!?��¹A��K&�D ��?xQ?���>�7��N�ս�)ּh��ۀ��{�?�(\?;@&?���)a�c�¾�3�<Y#�!�V�]��;�ID�%�>k�>򈈽���=�><Ӱ=�Sm��I6��f<�l�=�|�>y�=j+7�8q��=,?<�G��ۃ���=x�r�)xD���>�IL>�����^?�l=� �{�����x���U�� �?��?Xk�?����h��$=?�?d	?<"�>�J���}޾9��Qw��}x��w�W�>���>��l���G���љ���F����Ž�Nѽ���>�I�=&2?��>�#!<�?���X�O��U�\�3�-,B�����v�A�[�W�W�:�{��z��a�=vȾb���ɏ>E+��ڻ�>��?�m�>W�~>x&�>Oy��wE>�R�=i��>�>��x>pv>���=�E�=�����N?�@뾁h��X־�Ѿ�o�=?��`?հ?��b������s?c�?c,�?�%>q�j��H/�5`?#�?�X�@�?ܣ�=]nؽ�KK�dľI������WQ�-f�>IMļa )�wl<�CR���?�P	?Mݪ��پ�7���{���A�=�?��?�'�HO�p�uN��lY�e]�=�P��׭�}��X2r�픏�n������J�(�;��=Vx(?�n�?G���(]����g�q��+R�C�+>F��>Nm�>���>Dw>��ë,�MW� l�.�x�vu�>Pi?%ho>�J?yA?,h3?5�`?���>���>'ݾ���>ԉ$=h��>B�>3�?#�?�D?p�I?ۉ?��>���]׾z���8�>5�?��>���>f�>�:���"��n�t�<��]���=��w>�30>L���#��]|=�/;>��?���+<��r��`Q>�,?��>;��>e��8-���zF���>6
?���>�9��	v�����>��?�+���z<��$>@��=���%8�?�=�+���L�=
+X���C�(剼���=���=oI2<�0�<v�r;�g�<0��<�t�>4�?���>�C�>�@��+� �_��f�=�Y>HS>~>�Eپ�}���$��p�g��]y>�w�?�z�?��f=��=��=}���U�����I������<�?>J#?'XT?_��?}�=?`j#?ҵ>+�hM���^�������?�4?�z�>|�.�A����ާ���-��Z	?$m?6�X�!!��!3��壾��׽�I�=63>�-J��o���<D��
>��'��� ��?Dӟ?�����NB�T�̾r5���4>�r�C?�)�>iҚ>���>��*�!j�{��īJ>�?�[?8��>#�\?͇�?�>?5=x�B����C���ZC�<ae�W�?F��?�ݎ?ˇ�?���>P�a>�N��nk(�,������^�P�d�!>[^�=Eea>���>>��>��E>�W%��好C���|aٽq�q>^h?u@�>�o�>�1>���@�B?�?�������K�����t�s_���ۀ?��?r�?*-=���E4�w���Ð�>�U�?�ߪ?�� ?��q��}�=H��������Z�ף�>�)�>��>�Z�<��B=ߔ>c�>r�>����(�c @��䩹��?[�7?���=��Ͽ܉y���{��_�ro����ξYI��_5p�� �<r�>7Ԩ������?��"̎��,���~�3,v�֊<�b9�n��>z)d=%�=ˮ�<��=��=G��<�2�=X�C=x[ݻ�w�F>t-<>E7����@����=!ֱ<��F�ކ˾�}?=I?�+?��C?��y> B>n�3����>َ��??&"V>��P�:����{;��������G�ؾ�y׾_�c��ǟ�J>�CI���>;3>�K�=��<|�=�9s= Ǝ=�fT�B�=��=�n�=�b�=z��=�>�J>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��7>�%>�R��T1��\�.$c��dY�'�!?o;��~̾ٞ�>�[�=��޾�ƾ(*=�w5>h#_=$��\�-�=>|��o;=m�k=G�>,�C>��=����n7�=�nI=�l�=j-O>
�~��6���*��|5=]��=D�b>�&>R��>)R?��0?��c?�k�>P�m��	Ͼ�W���Ҍ>�=}��>�R�='�A>TD�>3�7?�D?��K?���>o6�=M�>ڌ�>�Y,��
n�{㾆I����<���?㿆?���>�wR<��C�E{�ͮ>��Fǽ��?�k1?��?�>�>*��w�࿓����^���Խ�佽 �
������M�\����k���;u�,�*>"��>��>��r>f>��t>a7�>RY�>�e�=8C<�#%�~BP��^/=�E���?�=5�-=J�=�1=��+<RJ���ĽY˞�2Zb����C;�=�O�=�|>�n�>j'�<"K�>B��;�Lپ#.c>����W�=8J=+m׾��?�B\��I���eI��~�=K��=�
=q�����>n�V>Lͼ=�O�?��g?	��>�1��p������*������(	>+?�=n'[��#0���R�t�K������>���>��>��>��3���Q�o��=�Q��� �̊�>^����y��-^3�ϳq������٠��5d�\��}�\?R?��O��=��?��/?A��?�|�>�W�<ّƾߡj;Q�ɾ�]�y3��k����?Ab*?�O ?�P��W��	�H{�$x�>�S���sN�����F^0���;�#���R�>߮��6�;�w,�HO��኿A�9��*@�a��>�rO?��?q�P��W��F�D�D%	�hDμ�v?��]?�Z�>�~�>�?�����aߚ�[��=��q?�+�?���?��=�N�=�b1����>{�"?V��?�ę?�O�?až�)�>=��>�p�>@g�����eME>��>O਼6}�>%�*?��I>���3��ܾShž�s<�U`ɽ��=��>z�U>~��>���<ٍ�=�@��@>�I�>S�j���>u`�>>ٗ>V�f��8%�Y�>G�`>]�9>\?Tȼ>�J�>5��"�m�e�p���ؾY@�X�a�͝�}dɽ0d���R�=��>o��>̿0!�?��=�b�@�>?(.��>�k=>V��<��>��>���>�tX>$�>���>b2>i��>�>�Iw���=��C�����q���T��Z徻:�>���}e�'~���� ��jT��x]�[�|��;�`l����e��?G���������=����� ?�>3sU?���Nt����>L]�>|�>������X�q�W��PDu?�?�;c>��>?�W?�?��1��3��uZ�,�u�f(A�e�E�`��፿����
���"�_?�x?1yA?�Q�<#:z>H��?��%�Tӏ��)�>�/�';��@<=o+�>�)��6�`�{�Ӿ��þ8�IF>y�o?=%�?yY?5TV� ���*|v=�`?�[%?M��?��U?f�<?VdǾx"?}`c>:c?�d0?���>�>4?�E?Ġ�>=�9��Q>T�M<:G齢c���K�������AD5>l����
3q��53<�L���%M=ڃý���<�>�'>M>׾�<L;�>�r?;7?�%>��@?��0��,� �P�̏E?2>��%��k|�*�J�����>4�?���?eQ<?���=0FX�S#�2�>--�>g�>���>X`�>N���nbs�WF�>TY >X'�=/�<y��qԅ��(������I	I;��=��>�Y|>�ʍ��'>�k���#z�f�d>1�Q�ۨ����S�y�G���1�Aiv�UD�>��K?��?��=�U�'L��gCf��*)?�U<?�KM?~�?�^�=��۾��9�\�J�~��y�>� �<�������}!����:�U��:?�s>-���Π���b>���O޾zzn�( J���羂K=>����T=J���վ���.�=�M
>b���� ����gϪ�}J?5\k=@Z����U�ds��4 >��>ˮ><���y�\@�����4�=��>�9;>=J��x���_G�L`�غi>�	K?��I?��o?��u��\��M5�7����ؾ̶J��(?��>��
?'K�>�6>v������I�a�I�_�ע�>�  ?��ھ>�&��Ԯ� %��]D)��d>��?�>h�?��7?��?גb?u�6?��?�͟>�\��u ��?�0�?��=�5�)u"�Eu�P�g���>zf??R�⵫>�5�>��?ku@?�8m?�2?��^>J�
���y�#Ŕ>�T>DG�[����9�>\;O?fph>E�?&Y�?B�>��7�����l^�޾�`�]>=>?Z�?��%?:�>�	�>Mw�����=k��>&c?�2�?\�o?H�=3?��0>��>숗=�՟>���>�?BSO?��s?��J?���>$�<����ԁ��ڻr�f�O��ŕ;$�N<�z=�� �Q�u�}��`=�<k��;�Y��̚������~�C�1{����;�_�>��s>!
����0>5�ľ�O����@>1����P���ڊ�R�:�H޷=���>��?ક>�X#�۸�=8��>I�>!���6(?��?�?`�!;��b�Z�ھ��K���>�B?���=��l�����%�u���g=��m?�^?_�W��&���b?(^? ���<���þ�@c��/꾶VO?1�
?��F�L��>y/?[�q?�j�>��e��n��%��3b�2�i��n�= ��>k���d�%�>L^7?��>�^b>O,�=P�ھow�}����W?�?��?_��?��*>T�n����F������^?���>����\v?����q���ݓ�苾�&������������L��K*�^~�`=ؽ@��=��
?=1d?�g?.�S?�����b�fJ_�\�~���W�����h�L�H��D�
�B���q�H]�ݾ��㝾oZ�=��w��nB����?ll&?ҽ0�X�>ˀ��  �<@Ѿn*0>>����H�1(�=i����A/=-Sa=��[���"�������?r��>�c�>�=?&0Z�
=�}w3�~�8��I�@ ,>Ql�>�ڑ>2�>�3<މ'�Vｄ�Ǿ�����ƽ�f�>��]?��7?"�m?P���lW8�@�z��:�@�����R�b�>���>��S>�8�O��LP�>�� v�?��]��h���I誻c�?.�\>�h�>�?'��>�A�b2��y��5>�*[Z=c��>%EZ?�l�>�\�>�.��-\E�h�>��l?���>h �>�i��lc!�%|�$KͽL�>���>M�>\rq>?-�O�[��L���t��Zj9�B�=�h?Fc����_���>t�Q?`Ϟ:�B<⢢>lx�١!�o ���&�`	>@�?���=I=>�ľ���ȸ{��Q��e�?��?�r���;��̱>&3??/�>U�? x�?�9�>�����#=Z?�-Q?<�Y?W?��>�=�G]��8��2��6�=LS>��x>�:>��>�������B�ݽ�T�=x�8>!>�0��0ǽ�+��\�{��۳8��>;mۿ�BK�=�پ�*�w?
��爾ȩ���c��S���a��~��vXx�ʍ��'��V��7c�]���F�l����?�=�?����1��A���R������h��>e�q�g�������J)��[��=����d!��O��&i�5�e�s�'?ố��ǿ'����;ܾa  ?�A ?ͧy?
��"�w�8��� >sO�<K?�����̚��#�ο����f�^?n��>.�5��\��>F��>��X>\Jq>����螾�5�<�?�-?��>��r��ɿ1���8��<2��?��@z|A?	�(�ڽ쾈V=A��>��	?��?>�O1��K�� ��pO�>;�?���?�jM=��W���	��e?R�<��F��CݻH$�=ZF�=X=�����J>#Q�>����QA��Vܽ��4>]؅>#�"����G|^�6��<�]>��ս�;��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=Y�3�ƿ�$��|�r_=��ݺx�[��}�հ��<�T��#��fo�J��a�h=$��=݈Q>Tl�>{%W>M4Z>gW?Z�k?�N�>�>[6�
���ξ�x��G��f��4������W�bR��߾\�	�������Z�ɾ� =���=�6R������� ��b�ȖF���.?9t$>Y�ʾ��M�I�-<3pʾV����ք�M㥽�-̾�1��!n��̟?
�A?������V�_���S�p���ۮW?qR�5��O鬾���=ś��9�=�$�>"��=���? 3��~S��f0?�`?>w���t��>U*>ڢ ��Z=z�+??�?mZ<!�>�I%?��*�D�㽔�[>��3>=У>���>��>o���O۽ш?2~T?���Dݜ�Q��>�T����z�P�`=�O>i
5��r�-�[>�h�<�����\W�f_��ٶ�<�(W?{��>��)��ka��}��X==��x?��?.�>e{k?��B?.Ԥ<h��p�S���Law=��W?%*i?��>Ƈ���	оZ���D�5?ۣe?��N>�bh���+�.�MU��$?#�n?'_?O~��w}���p���n6?��w?Gk�+������,��>>:��>�h?C�3���>s4?��M��}���^��/�9���?W�?iU�?Ei�;� ��fe>4?�c
?��6�Ͼ�Mռ�짾1S=M��>�x����b��|,�y?a�I4?ԋ?�5
?h����m�C>Z/��3�?�փ?�u���?=m��7f^�������J���Ž@��"�־72���ݾ{���j��C�=���>��@��i��/�>Bc�ۛ޿��տ�Y�������j��A?��> �&�9���d������;k�S8=��Cb�@M�>��>Ѵ�����/�{��q;�*����>��

�>p�S��&��������5<F�>]��>���> *��^罾!ř?�c���?ο\������V�X?	h�?�n�?�p?��9<��v���{�x}�".G?��s?4Z?|o%�?=]���7�o�m?D�� Uh�z�?���O��"">H70?���>�0,��N�=��>���>���=�g4���ÿ�ܶ������%�?���?�����>�F�?�.?�Ae�������6��<N!<?�t>>�ᬾk+���>�O�{��S?~w<?z���}&�]�_?*�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�f6%?�>d����8Ǿ��<���>�(�>*N>`H_���u>����:�
i	>���?�~�?Qj?���� ����U>
�}?;��>��?�*�=-��>a��=�2��aU�P�>5;�=�����?&WM?��>Uj�=h1+�c�-��qD�άP�
��A?�)�>�<^?�F?�wT>Û���������K�L�w�f�mq9��ζ�	U�� �?>�@>�>��=��l�M;?�C�t��z���d,��1��>�A�>��?����E��ӽ����?d��>��+��ŷ�|����}���`�?���?_?�ƾ@��;�\>^%/>�	#>�_�Ն=mC ���>�2?�������^�c��>�><3�?°@���?�%����?��	�q����B����
���I���=}v9?���>n��>o��=�yt��Ъ�u�R�>ܦ�?�?�e�>T�g?Y
j���;�)\s=���>��d?l
?�	<+�Q�=>��?�U	��W��Q��c�f?:�
@_h@$�Z?rƣ�A?��������^���m�ypH>�>�)7>l¼�>�ڈ=m�<������=��>"�b>�I>&�L>E)�=��J>a�~�����ݝ�!-��q�n�
�I�L�)�/R��8)��������x�Ӿ'U�����> ��1Ƥ��b���=�<���=�,U?�YN?��l?81�>��t��>�@��R�<C#,���=x�>]m0?^�K?�#*?���=�뛾zKc����bƣ�����s�>��@>L��>��>̭>^,���:>�#>���>8q >�5O=���<�10={�K>Q��>�}�>� �>�C<>��>Fϴ��1��k�h��
w�r̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW? �>!��u�T�4:>9����j�5`>�+ �~l���)��%Q>wl?��f>�u>B�3��d8�O�P�2|���h|>�16?붾�G9��u���H�lbݾjJM>)ž>�%D��k������}ti���{=�w:?�?e:���ా��u��B���LR>X3\>Ic=�k�=�\M>UPc�y�ƽ�
H�bj.=P��=)�^>�M?��+>v��= ԣ>BU��AMP��x�>�3B>��+>��??6$%?@���嗽"l��S�-���v>?8�>���>�>3CJ���=b�>U�a>��|B��b��S�?�f&W>���#S_��u�GEy=����%�=4A�=#f ���<���#=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>�Vk�`tt��U�}����ko�>�>?+���=�=��@����>h�?Y���󨿏ʿz�����> ��?'�?m��㜿-�>����>K��?'^]?�y>�+ܾ ">��P^>�G7?o�K?��>)q��jD�y�?�I�?�{?Y>Z��?��[?���>��H��1��Y���ӎ��Q�=�=5f�>�؇>�V��>�����bƅ�������g�>�04=���>4	{�l��2�=׍���/���ʽe�>�>#�>��>g�"?O�>���>��>�]��MP��S�K?=��?����3n����<�=z�^�/?	T4?p[�T�ϾfΨ>.�\?p��?7	[?�w�>��9��迿%|��12�<��K>�$�>�P�>�숽TjK>��Ծ|-D��r�>Rŗ>Z���/ھ�7��gI���;�>�]!?W��>��=��%?�n?�Y>��>"H8��ҍ��^X�!��>�l�>��?*y?=I?�,�a�3�rl��N⡿��k��FW>,;v?�t?���>$܌���R�<Fo�����#jg?�t_?5����'?���?kK?+2?���>e��Ul����+�T-b>�!?1a���A��(&�2���Q?�*? 9�>�򔽟f׽_�м����I���?
\?I
&?!���a�g@þ-��<]�K�C��_�;UrJ�� >�>�v���^�=g�>���=+�l��:5�2(s<�w�=��>\1�=0�6��9��^�%?�콜���Bh=�5���Ba�^�>쎉>��ھ��c?l�T�l�y�H鬿���`U���b�?ƽ?>�?f���՗i��M?��?�-9?pD?�ǁ�d ��p����ڇ��壾��.�&o=-�>x�ü��`����������jg��^p�3��>XeK>�?5�>[b�=K� ?;�G���ľ��6��k�>�&�B�G� �;�Ñ ��ܯ�p��!�H=�.��y�z�.�>� �vX�>�r?v�V>>�>���>u�E=��`>��>�w�>#�>��>N�s=&R=M��<�xM��KR?�����'���辽���b3B?�qd?D1�>i�<��������?���?Ps�?=v>h��,+�}n?�>�>@��Xq
?�T:=�8��:�<	V����53��2���>�D׽� :��M�!nf�xj
?�/?�����̾�;׽P����I=6��?e�+?��%�� N��Mu���V�sL��Z�3M^��ۣ��g5�#�j�[���܆�][����6�=6c'?��?/���G�%�����n��J��wD>*��>�ݫ>PP�>�
�>�(�5�$OZ���(�c��AW�>�n?���>a�I?<?�/O?��L?}v�>,q�>�2�����>|W�;$g�>���>�v;?d.?��0?�?�/+?��W>z��T����)׾��?a?X?-?P`?����d�Ž)�K2���l���=��=���<o���QR�m�I=M\>&S?~���8�O�����j>�x7?�v�>��>5$���9�����<R�>C�
?�M�>����~yr��a��F�>.��? ��B�=4�)>���=���oɺ�Z�=�������=i���7
;� <J��=�2�=��m�%�R�g�:�҇;=��<.8 ?J�?�ٍ>��>����z��"���=��S>��D>��>�پ�W��������f�H�s>7��?�(�? �=�l�=,%>qΣ�������Eþ��"<��?�.$?x�U?c�?��<?��?H0>eM�S���2��C����??w!,?��>�����ʾ��։3�۝?i[?�<a����;)�ߐ¾��Խѱ>�[/�i/~����>D��텻���V��6��?�?JA�W�6��x�ۿ���[��{�C?"�>Y�>��>U�)�~�g�s%��1;>���>lR?��>^�R?r?�X?�D>��7�p%��x"��p޼��,>O�K?���?I�?�yr?:��>:�>�2[��}��V�7�c�Ͻ��k�i�i=�rM>���>���>��>",�=�������Y��6�=N�>.��>��>���>>�K>4C[��5G?���>>����A� ��fG��TY���v?�S�?��*? |=U��� E������=�>ନ?�u�?�p)?�vZ�f3�=T����i�s���>�H�>XA�>�n�=�^G=�>b��>Pd�>�	����<78�hO�J�?׻E?X�=Kſ�,q��|������,�;����Q��
���_[�y
�=ӡ�����Ԫ��	d���N"��_{������J,p����>@ c=A>��=u�<	i��dͭ<�=�J<p�=�B�a��<
��U��95�r��տ<`H\=�$���ʾY�|?��G?��*?S�B?��t>�Z>��K�3�>yȆ��?,�Y>�XQ��~����7������`��� پ�Tؾ~�b����{>H�[��U>}7>_��=��<m��=��F=�ڒ=v����~'=2+�=-�=Wl�=���=�>�>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾp@?}�>>�2������yb��-?���?�T�?>�?@ti��d�>L���㎽�q�=K����=2>p��=x�2�T��>��J>���K��F����4�?��@��??�ዿТϿ6a/>�v6>f�>3R�O�0���Z�j c���Y��?��;�й;8h�>��=5*޾��þ��6=Y�3>�5Y=��p\��[�=�p��3A=�e=\�>��E>j��=2���iL�=�-=z$�=QP>��X9v{$���ל9=u'�=�a>6�>�~�>�?(Y0?�?d?M�>p�m��XϾ/_��-\�>Qf�=�^�>�z�=�B>=ϸ>�8?,�D?�K?@&�>���=��>�	�>o�,�n�m��徢������<0��?>�?F�>�KK<YAB�z��UR>��5Ľ8�?�K1?�i?�Ǟ>�U�ȡ�VX&�r�.��~���$�*+=lpr�'DU�����k� ����=�p�>��>��>�Vy>��9>��N>p�>j�>0�<Ds�=����ص<��q��=�������<ż�����&���+�������;���;ј]<�R�;��=���>��w=�$�>r����Ծo��>���-�Q�2Y�=�a׾N�L�j@m�����=x;���,���6>�l|>Æ�������
?ەO>��>���?4��?��V>�wJ�UB���晿�A���q�]��=ԇN>a�9���>���g�g�G��~�����>b܎>l�>~�l>�,�]$?�y�w=C⾊b5�=�>�}��u��9/��:q�@��8����i�0BкQ�D?lF�����=�!~?�I?��?��>G���ؾq90>"J��z�=$�#*q�Gd���?�'?���>?��D��̾�½6��>h�G��O������V/��$�����m�>�Ƭ��Ѿ��2��c���᏿?�B��?s��X�>�O?ˮ?�d�����ްO��_�A����?ɿg?\�>s?
�?&a������&�Ud�=�|n?=W�?���?�M
>x�=�<��zU�>��	?U�?~��?%�r?�B����>��<���>�����A�=.�>Z�=(�=�&?�	?�?_����	�!\ﾚk�g�]�"�=���=�$�>�)�>	Up>��=bc`=֜�=1�[>���>���>�je>Jz�>q9�>�9��v�.�$
?�|�<8�>m�?�,�>^y>YR��*�=SL��g���(���|�L�p��Ɛ�O>Լ��o>��=��?�S��.�?�(=*��1?�� �u,<U���a��M�;�u�>�} >���>5d�>��>v�>|��>W�R=�	������&C�e:;��\C��{W�#�־x�a>�����<[��,���J�+�(⹾���(y��ꄿ�dV���*>�Ə?6���.���M�м־9O�>^��>g�?�';��=/�R=3\�>�+�>��0�1~���u��%�����?���?iׂ>��&>�%h?f^	?-^8�t $�d�2��Y�H�P�Ă�*y��Ç�Z��p�	�#V���P?���?2J?��|=��>'I�?����n��\_>l[$�O�����g�>�þ�t;�$����!�M���sm>��I?To?�?{y����т�>2?��?�d�?�W?��?5�	��B;?�۽73�>En?5	V?j$??��+?_� ?���>:h��t��<'���p��ɹ��2�=�=M=~x����=��Y���=9��FF]��17�����gv<j��P���,�=���<�+�>8�>��]?�R�>��>�8?V���9����1?oM>=s7��\S���`��G�A�>O l?oM�?,Y?}�Z>�B���D��7>�2�>��*>��`>ߵ>�޽M�F�ӓ�=��>��>�{�=�e�f��?�	�2X����<Z�&>��>�/|>����'>�|��m0z�,�d>5�Q��̺���S���G���1�ʅv��Y�>�K?��?���=�^�,��<If�Q0)?�]<?�NM?��?��=�۾��9���J��=��>�X�<��������#����:�!Ҝ:e�s>�1���]��O�a>'�
��ݾc�n�-�I�X�羃�C=^��*�U=߽��־�;��E��=��	>"P���[!�'��ͯ��9RJ?�)p=�̤��T�������>f�>�î>+�9��xv�ӄ@��|�����=���>P�8>���������G�Vl��ל>�xO?^K?�s?5\���p���^��5�е�c���0?*��>�?0�W>�<=���!�%���d�K8L�k�>���>R��D;2���B�
�Tj�y�g>�{?^S`>��?zRQ?6?�.�?�QX?J*?+��>��4�{�?`��?��=W���m
��1��k<����>n�"?C8�%�>�j?�o?�t@?M�d?�7?��=>_��[��؃>Fj�>X<�<�����x>_%d?PhY><�v?��?�xe><���0��!���۽G!Y>��O?ݵ2?xN?�>'�z>ڢ���/>}->BOl?���?�t?D��<eN2?����t�>��=;�q>J
?�� ?�U^?*gz?�?�$�>����q὎ �%%o�Z=��;*�=��	>��e<;?G�맑<��->FI=?۽��ř����3߼4Q=�`�>h�s>����0>��ľPP��i�@>�	��BV��ъ���:��ͷ=U��><�?آ�>wa#�*˒=1��>�E�>u���3(?/�?Y?��;�b��ھܯK�i�>B?���=��l�Ȁ����u�Th=��m?��^?J�W��&��E|b?s�^?,��5i;�.�þ��g�Yx��K?��?�K�Ь�>�e~?�kp?Β�>3�i�߿m������b�E�p��Z�=,�>���n�b����>�e2?Z�>c9^>O��=�OվS�s�mw�� �?ޜ�?X��?F��?��3>��m�l࿾��$����a?�4�>��þ<��>���}��>q��G/[�
���Ɠ�����@T��:����\��ϛ���ν�=F?!�t?�?g�s?��$���<���g�'t~��<C�yL�ן;��gT��=P�J5�YЄ���I�,tJ�X��Ԕ���ˀ��A�ɽ�?�'?vQ3���>%A����i�;A1B>"���_�CD�=���;K<=<�G=DIn��2��Q��ɀ ?��>&��>��<?C�\��~=��$2��;7�ž���F2>h��>��>��>�S>;+n2�^���˾Q���h2ڽ��>�rh?'�B?qZh?�\#��<8�]@��Z�%�ד������e>G_Q>d��>�� ��	���"�74A�G�p�� ��ғ��g�ȟ�='/?S�i>1U�>���?���>�O
� ��Mg��G!���=�.�>�t?�|�>( �>G���H#�־�>L�l?a��>2�>����{S!�"�{��ʽ��>;ӭ>;��>A�o>W�,�[(\�1k��ƅ���!9�X��=��h?e~��4�`�9Յ>�R?Q�:~H<�W�>3w�~�!������'�o>}x?>��==�;>(�žT0�w�{��(��Q}$?x�?�쎾��*�A0�>�% ?���>�\�>�q�?���>|����;��?�V?��K?��I?���>��/=�u۽?�׽��+�{(=�P�>��>��=��=�%�%+j��!E�#&<�
>�I�<�ZĽ]����oh��09��=�T>�jۿSK�R�׾���=����	�����u���ˇ�?Y�ʶ��U��k`x�Y��>���`S�d�`��d��!�i���?���?�#���Ά��Ϛ�����������>��u�Qzv��>��a���`�����}���t"�Z�P�bi�Ie�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >WC�<
-����뾭����ο@�����^?���>��/��o��>ޥ�>�X>�Hq>����螾z1�<��?7�-?��>Ďr�1�ɿc����¤<���?0�@�xA?��(�o(�7W=���>�i	?_�@>�?0��i�SJ��3,�>��?�ӊ?�]L=	�W�iu�9we?Ґ<L�F�@�ݻ:x�=�֦=\R=���ڵJ>I�>A� �A�� ݽb`5>B��>QY����o3^��J�<��]>�Xս���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=� ��l����X�6���9=<XRy��QT��Ϲ���:���O�CL���B�@>z��>�?�>ٗk>��y>�ZV?��t?�.�>��b>�5k��Ӿ�%Ͼ��?��gy���ϾW�c�����y�����e���F$�������!=���=7R�i���C� �f�b�O�F���.?�v$>N�ʾ��M�=�-<�pʾm���[݄�G᥽�-̾�1�#"n�i͟?��A?������V�X���W�񄹽K�W?4P�޻��ꬾ��=w���T�=%�>܊�=���� 3��~S��-?��!?���`;���gC>�,� ה<+?�?N�C<9��>3�$?�0�Y�۽�hh>�RN>�C�>��>��=$鮾FM�2�?h�S?PӽH�����>�dɾ�-��A����=����K�<��\>�Ĵ�98����̼�5����=��U?`L�>�G.��`������gO�Zr=�y?v��>P�>@�a?]�:?�_�FZ���3U������=�!X?-�b?�'�=�y�;о�ȩ�b�3?]�f?�i>��x��k���+��� �K~?r?� ?��Լm~�}�����{�1?C�?ӝb�+F���g�C��� {�=^�>I?�%�J7
?V�f?�����ڌ�v���#�I���?,�?6�?�v>=l����w>��?`?��z�����Ǒ9��?>2��>�Z����+���1�������B?G�?x= ?�[��������%>}З���?,�?���X��<u#�+]����?x�/Z6=����+�ν 8�n7@�X뾄��w8x�U[�� �>�M@T.�F�>�5�nJο�4ֿX�������^س����>F��>'������c`��!x�S|g��Q��LF�P�>��>ٔ�G�?�{�&q;�𿞼w�>>���>��S��(��y���'5<�ޒ>֣�>���>����㽾�Ù?�b���=ο����ɞ�`�X?�g�?�m�?�l?X�9<
�v�]�{��O��-G?��s?>Z?*R%�Q3]�/�7�Ux?m�ӾUǀ���T�z�W�t��=�g+?R��>��3��?�>�5�>��$>��=sT(�Jȿ�5��/VϾ�P�?F�?�ݾ��>�h�?Ƀ+?�#�I�������td���=�ZH?�k�>[@���3��/>��_V���&?wG?",��)�\�_?)�a�M�p���-�|�ƽ�ۡ>�0��e\��M�����Xe����@y����?M^�?i�?е�� #�f6%?�>d����8Ǿ��<���>�(�>*N>}H_���u>����:�i	>���?�~�?Oj?���� ����U>
�}?�'�>��?;�=��>�s�=!���$e`��� >���=��G��?>�M?f��>��=[�6��.��FF���Q��V	��QC�+L�>�a?X�K?�c>�ٷ�Z�(��V ���ʽ��/�z��^{@�(�,���ݽ�6>I?>Ur>�BD�p5ҾV�.?��%�E�߿�p����x���(?e)v>�z	?��
��轕fp=�%?/�b>w���IN��z���W�?�,�?^�?���l��>Y�=튓>��Y>K	 �ꮽ�ǚ�LPw>OIM?2g�T�x��jQ���W>���?P@-\�?�a}�qV	?�G�
z����~�A���~7���=��7?��w!}>)n�>��=K>v�����t�^��>��?��?��>�Tl?jCo��bB��-3=�f�>��j?�^?q9�pJ�USC>��?�m�2ǎ��X���e?�
@�d@@N^?㢿�׿p����򟾕=�>s�)>K>��_ϵ=�a�<Ey�ᛉ�6�4>&5�>,�>f�[>���=�)>_� >{����e-�t����S��G�?���1d��Ɩ�����j��/�	��u��5I��Moo<�K��̵��؅��-?�B�h�b�&>��_?�t<?�i?x��>�]���V�u���O���r�Z(>��>3�S?�Q?��"?�u�=����'J����䖾.�\�І>}BN>l��>ㄝ>�g�>��<:Y�>\�>t�5>&�<�ϼ��@=��3>A��>�J�>}�>�ȫ>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?J�f>|u>�3�^e8�h�P�{|���j|>�36?�鶾�C9���u���H��cݾHM>�ľ>rD��k�\�����vi�w�{=lx:?��?�7���ⰾx�u�C��GPR>
:\>nV=i�=YM>�bc���ƽ�H��g.=��=��^>5?��=�m����>=	����`�8#�>��><1V��T?D�?�������꒗�On��+��=��?~l�>�L�=�(��<)�$?=V�=�`*���ؼ�0��)�M��>J|�d��
iؽj >/��4'>4�/>@�	�"�����~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>/6@��^��59���`�� �Ƽ�>��P?�(���=@\��ڝ>GϺ>�s�����ƚ¿e�q�b?.�?0�?��s��y;r�p�>�U�?�L?�e�>���z"޽[�> ��>�{b?�?+�!�NOj�U?u��?-F?E1�>~��?5|Q?H��>�˿�����2��v����ӫ��%Ͻf�z>�>?�ʾ�jJ�������;[��y�s8>�=~�?XRܽ�#Ǿ�å=g?K�����m6�{�>�a^>>S�>� �>y?�]?%��>��>�uS�e���m���X�K?���?���n��k�<t�=t_��?Z.4?*]��Ͼ��>��\?%��?��Z?Sl�>����4��
꿿�u��Z~�<��K>�.�>�Z�>����WK>��Ծ��C�h��>��>�w��G6ھ�!����LG�>�a!?w��>(�=I� ?��#?�Ij>r>�>J[E��-��F���>sT�>I.?,�~?)�?����'l3��
���衿��[�|N>9�x? R?��>�������D���I�֓��J��?�ag?�.��
?80�?�??��A?5>f>]L�6ؾ.���q�>�!?���A�IM&�/��}?O?p��>l#����ս�!ּi��0�����?�'\?�A&?a��F)a� þ}(�<��"��U���;#D��>��>������=�>�Ͱ=Km�CB6�.~f<^�=x~�>w
�=�&7�h���,8?
�ܽ�����[�=��u���\�@X>�.�>�/���s?�i���z�4r��
e��ظ�n�j?�ٶ?��?8=���@Z�.�8?n�{?��3?��:?��)�%������`���̾c'G�a�e>�[>�7g�,b��v՝��@����~�����½z'�>_fw>�?5B�>�+ >aW�>(`E�9/�PT��İ�LPZ�{�&���2���9���+�F��+�����k���kn���>�v����>�?^��>�X>7��>q]���>�nC>���>Q��>
d>>�-> >���<[^ڽ�KR?����6�'�e��Ų��J3B?�qd?�1�>�i�������f�?���??s�?<v>h��,+��n?�>�>9��>q
?�V:=�@��6�<�U������2��$��>D׽� :�uM�Snf�rj
?�/?*����̾<׽;���Y�=h5�?r�<?(�S��59�h�i�v���+�H��D��K))�,�<O��v��.������gj���Th����]�M?�D�?�z.��1F�ȶ�ør��$����>h�>m�>��>�ͧ<.������]��R�jK�θ�>�O�?�st>?yR?{?�5?y?g?Qy�>�A>Lɕ���?�fG��dk>��?�Ka?x�?q-.?�?��(?��>ɖ���|?޾j�
?��?'?�B�>3�)?�O�������H}� 3���+�L'�=��4>�<�����A8����>Yz?fM�p;�̩���f>*�4?ܝ�>���>�=��$*m���<�>aJ?�,�>SE��t�3�	��C�>��?���\�<DM.>�U�=`x��;_F�=録���t=%������<���=!?�=O0m����;�51<8��;���<C��>��?�=�>��>���m� ��.��s�=�VW>U>��>LjپX������h�k�v>�Q�?�i�?��e=�=�8�=ri��򺿾C�����\n�<L?1�"?�T?[t�?ߏ=?r�#?�">���3��+"������1n?z!,?���>��~�ʾ�񨿳�3�ŝ?�[?�<a� ��a;)�.�¾��Խ��>�[/�Y/~�����D��������~�� ��?ȿ�?�A���6�z�忘��[����C?�!�>�X�>5�>d�)�3�g�f%�\/;>v��>(R?���>Tb[?G`?�F^?�>FD��é�c䒿��7��=��9?��?��?*�?��>N��=V�r�n4��4{$��z�5���<q�C��=0�p>)t>�5�>�;�>�v�=g'�)��,C��=�t>�?>.�>[u�>��f>=N���i??��?F;��w��Yk{��%R�8�����u?R͙?NA*?��=�o�mX?�����>uL�?���?@?�Õ�A<�=$n�!9��4tN�_r�>���>z��>}��=o>0G>�>�>'p�>p<'�?�!��1:��l�:?�@I?��,>O	ƿ��q���p�6㗾g4e<�В�`�d�������Z�W�=2������Z����[�@����r��B⵾���#�{�d��>"̆=P��=��=G��<�9ʼ��<��J=ӡ�< =�o��cp<��8��QһI~������^<�tI=���FEʾ؇}?]I?�o+?)�B?��v>U7>�]8�Dד>�G���&?1 Y>�$;�º�e9��	���ѕ��>ؾ-3ھ%Rd�ɼ���O>i�I���>�W3>�l�=�]�<��=��t=o׍=�� R=?�=��=k��=c��=��>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>X�8>�_>�!S�f�0�r�\���b�G�W�1�!?�};�{ʾCŅ>�q�=z�߾�ƾ%=p�3>��e=�%�,\�Y�=c|��@=�gb=��>3�D>m��=x����\�=	G=��=O>��M5�&o+��6=v!�=<�b>�C%>	��>�$?�/0?7)d?�,�>Iqn�>1Ͼ��"k�>�e�=���>)-�=T�B>���>�8?�D?a�K?��>�Ȇ=��>�	�>��,���m�����&��4ڪ<ᚈ?.�?��>�V<�RB�ɲ�*c>���ý��?�a1?�a?DԞ>F��y����[��6����i>��X>�|1��;��I�KQ����<x�F>��>ts�>��>xi>�F%>���>@��>Z�>!<�=p���C���'=��N��Z==9��<��6>�/�=�k>:���2!��}��)�<���=��#=�f���*>R��>ծR=n��>/V=b�ʾ1�2>����K�@{G>�����B�? y�q���1�8���u�LM>x��>��܋��� ?ڹ%>�J>��?\^�?r!b>\�n��� ����;��m�)����=��i>jq5���S�[�_���>��4ʾ��>�ώ>e��>��l>8
,��?���w=����g5���>�x���7�9E�
;q�;?�������
i�p<��9�D?7A����=8~?]�I?6ݏ?���>g���@�ؾ�.0>�a��f�=z��q��i���?B'?�k�>�쾂�D� ���&�k�[>Q�8=�^�ⴞ��#�͜J�����s�>Ӣ�0� ��[�����K'����N�r떾�#W>׫x?∷?�/��@����d����iM�����>���?[׫>��(?� (?�K�ѵ��?����;�d?ڨ�?'Y�?��><�=t��f��>+�?�Y�?���?�vs?��C��q�>ˑ(��>�ϐ����=�R>6�=o�>��?�2?��	?�@��0	�h��s�Y�Q+�<�N�=俒>��>xj>��=3�o=Ja�=K�N>]�>��>�N]>Gɡ>{	�>\���p|��3&?�=W3�>��1?�i�>Aab=II�����<NSG�@���+��+����作J�<�+�l�W=�ϼ/��>�Tǿ�Q�?O�Q>���(�?m����u0��R>*S>	h۽�D�>'�F>)�{>Ԁ�>T��>�o>�@�>
�&>QBӾ��>f��vY!�p/C���R�ƾѾ�bz>�����%��������`I�x��^k�bj��.���?=��c�<lI�?M�����k���)�B���|�?^�> 6?9Ԍ�ڈ���>���>�>�N��ɐ��^č��W��?`��?�;c>��>F�W?�?ߒ1�.3�vZ�&�u�p(A�)e�R�`��፿�����
����&�_?�x?2yA?�R�<):z>Q��?��%�Rӏ��)�>�/�0';�q?<=u+�>/*��9�`�x�Ӿ��þ 8��HF>��o?4%�?pY?3TV�z����>�iP?v�?�s�?~U`?k&k?���\�9?hb��#��> �,?w7?[�;?G)?���>t̑>e$"��>E[��<����=N���!���=^��<�#"�M��=�SW=-"Ƽ^Z�^w:�ޓ��cp=q�6>�>��=RQ�;q��>Y�e?U�>�A>qb=?�A佹�8�xgx�WI?�C�=��b�Au��۞����2�C>4y?r�?��L?�>g=K�ՉH���=
Q�>.S>B�`><�>�$*�k1|��C��}R=u>C�@>(6U��%���1���"= e>C��>.|>����'>y��O+z�֚d>�Q��ʺ���S���G�t�1�ւv��P�>��K?��?���=�U�u<��,Ff��-)?_\<?}NM?��?��=��۾��9�w�J��d�$�>ٽ�<������!��F�:�B)�:��s>�,��NȾ?;s>���J^��.��Xf|�(Dپk�5��f����=��O�E��TJe��L�;C�>������!��\T����O?�+>�,Z�R����Ⱦ�>�ex>���>R����T��/a����\�g%�>V_>�7g�L����{�V��>�E?�?_?)�x?tt��#�k�7�F�	z�ID���Mּ�.?@O�>��?�>�|i=e�þ(����V��<�1�>��>]R��YH�ճ��)���'v3�.8g>�?�cL>��?(aP?�/?�me?cr5?eA?��>���D��צ#?�?���<�Gۼ�Y�_� ���<�� �>%[?Ѣ�p��>^��>`L?�1-?�GX?)�?�|9>`�Ͼ��K����>�L�>�K�k'����L>��M?��>�p?��?�->O���?پ��&�U�ǽ>��H?Ad ?w�?J�>�Fg>�t��31s>Q�>H�|?�~o?9t?N�(>�S,?����L_�>��=P�(=��>�?�_B?^[?��?c��>>�!=bg�<�ρ���Ľ��ż��1=�>5�<��E����<�׽���=5�>�"]=���F�V��m�U:c�A=�b�>�s>���0>��ľJ���@>�����Y��+ۊ�o�:��ط=V��>�?
��>:i#�Ɗ�=���>�L�>^��=:(?h�?�?��;��b�[۾��K���>�B?`��=��l��~����u�*h=N�m?\�^?5�W�%.���`?_?����GE��M��w�������"? q�>*��"�>�*?�\�?q�>�_��j�i����<F�oH��^m�=��>��
�7cW�	�>ܖ?�q>�>�>�c����Q��]��>X"?�D�?ӷ�?�l�?E�>��w���P�ؾ�Y����[?Ky�>����q`?�Z==Ԥ�g?��ߙ��f���1�����u1���u����l�n^��u����@>~�?�w�?+�s?,�X?�>xZ�F�[��ȃ�Ā^�K�/B��DG�ZC���O��Lg�Z���2	��`���=z��<A��>�?�j'?�y4��@�>Η�;𾅔ξ��B>@(������3�=�ᓽ J5=��I=�wj�?.����>C ?�>���>E=?!�\�-�=���0�(�7������?/>1��>�}�>$E�>sd�۬*��h��Hɾ�;�� o޽ǂv>�}c?��K?_�n?��!1�T���C�!�b�2�.���C>Q�>[_�>��V��6�&�{H>�-�r�i��n��M�	�F~=D�2?^�>#��>�B�?��?I	�k[���Yx��g1�`rx<캺>�:i?���>ZO�>�ѽg� �U��>N�l?���>t�>|挾�a!�č{���Ƚ)��>-A�>��>u�o>ph-��V\��~��x����C9�z��=��h?MƄ��k`�*�>�Q?�!J:�0M<e�>&w��!�jj��C)���>�_?x��=��:>��ž*:��{�檊�[O(?�?X듾��(��ւ>�� ?�@�> ǡ>!΄?z"�>���Le;�!?�t\?�QI?3)B?�F�>��=�޺�!�˽C�'�]U7=��>��_>aqZ=���=iz!�AkV�i%�i�F=���=lRü�®�8�;lrмH<y��<��.>#�׿�gG�>핾����
�Q�:��h��֊���q�-IU=����:��
]���D���x��T���A�ދ������}�?-��?)�W�� �<�α�ց��yN޾'Q[>�������֨�;�߽�-���`�]/��W.���&������pv���I?~x��$ݿHu��uR����<?=��>�w�?'������9��s��=H�m>⤽� ��И��[Ͽ��]���j?9�>F�J)���>R^�>{����>ʻ�"Q���< ��>��?;��>�Rᾭ�ɿm��(M�t�?��@/gA?��)��z�"%U=.�>�	
?E>��&������F��>��?�Պ?*5S=�cW������b?�Sm<M�C��������=���=�8"=����sK>�>����M��o�k39>U��>�%�M��.X�N^�<�BX>�mɽ���2Մ?
{\��f���/��T��&U>��T?+�>�:�=��,?I7H�`}Ͽ�\��*a?�0�?���?,�(?0ۿ��ؚ>��ܾ��M?SD6?���>�d&� �t����=9�'��q���&V�<��=m��>u�>��,�ۋ�_�O�K��;��=#��9�ƿ�2��,����<�q��Zʏ���"��
����B���w�q�R��E�>�=2��=�vF>�w>�JQ>��p>T�V?<�u?^>�>l�>�%;�����
�����}p�^����������*������ݾ�H��e��J�qk��� =��=f6R������ ���b�ɗF���.?Rt$>N�ʾ��M�/z-<fpʾ���� ��好.̾��1��!n��͟?E�A?"�����V����`E�����W?�P���R鬾\��=������=�$�>`��=���f 3�J~S��.?^�%?��ľ����T�M>ݞ�����d%?�D?��<gФ>b?G�"�K�����`>Q�`>���>E��>��=|����
뽹�?=�W?(�˽2���b͌>{xѾxP�s=8>��������j>��j�Z��+f<V[���;�W?Q�>�j*��}��~��G�#���M=��x?�$?�U�>�-i?
!B?��<?����T���ز`=��W?,bi?�/>tk��ξQg����4?�fe?R>VJe��-꾢F0�p��b3?|�n?�?#���}���`���u5?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?p�;<��U��=�;?l\�> �O��>ƾ�z������3�q=�"�>���ev����R,�f�8?ݠ�?���>������<�>�������?�=�?���}�0=�A�"^�A��U����Q=�P��:$�'b�w�<�:��t�۸}��!�= X�>��@u����8�>p�~���ۿ�`ѿ�D��N�ƾx�B��`?>p�>@ˬ�ƴ��ؙd��k��CD���H�?a���0�>s�>*n)�����v���-���O���>~���V�>�e����
T��7�&;T,�=�$�>�>PI�ٔо�U�?�p�~������[���?�/�?k,�?j0?�X>��<�� �8޿=,2@?0h?fs?���U�	��ݪ<�T{?�
���,h�Y�&�IJ����=״?��$?%Z7�#�>Ԩ�=U�>ֻ�=Аh��Vƿ�Y��5�?�?�?}�?co�/� ?ծ�?U�5?@(�����їY�,&>�%��ɡ?]��<߲{��9�D�5�'aX����>�?M��y��]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?N$�>��?o�=�a�>�d�=3��-�\k#>�"�=�>��?��M?�K�>�W�=O�8�i/�[F��GR�Z$�3�C��>w�a?݂L?kKb>Q���2��!�Jvͽ�c1�NP鼀W@���,�l�߽(5>��=>�>;�D��ӾE�?t�^�ؿ�c���'��$4?	�>e?���@�t����f_?�s�>v1�2���%����׏�?)A�?��?��׾Ekȼj>V�>4[�>�	ս�㟽T��5�7>��B?���2����o��i�>��?�@�Ǯ?�h��	?���P��Va~����7�i��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�O�B���1=9M�>Μk?�s?aQo���i�B>��?!������L��f?�
@u@a�^?*h�߿����ּ�G�羱��=S�=�4o>�M��~�=��="z�<V6N=��";���>�_�>KKE>��/>�O >�&�=�˂��#��ޗ��񘿌�^�Ir��\
��Ͻ N�`_��y�ݾ�p���ξ#���a������"��|�X���f>E!V?D�E?j�v?���>���N��=j����e� U����=�3�>��'?��d?4�5?5ٸ=)񅾱�_�u���q줾�m���>�{R>-+�>@+�>���>�8=�+o>n�9>�/p>G4>=TE�� G�,ϔ<|.>�i�>B�>9��>tJ<>>Dд��2��e�h� w�i)̽~ �?򂝾%�J��0���9��죷�El�=�_.?'w>���V>п�����3H?����+���+���>8�0?eW?��>L���T�
?>F��[�j��^>�) ��{l�Ə)��,Q>[n?��f>�u>�3�8e8�>�P��{��Of|>�36?�涾�B9�U�u���H��bݾFM>�ľ>��C��j�1������vi���{=%x:?S�?�.��䰾��u�pE��;SR>�9\>�O=�r�=AYM>HYc�F�ƽ�H��o.=��=ά^>(J?��,>
 �=��>�♾�P�s:�>$BB>��,>I�??P%?�������Y���u-���w>���>��>��>�VJ����=np�>b>���g!���E�y�?�32W>��b_�G�s�3"x=����(Z�=���=�f �_t<��^%=Ֆ~?����㈿�ie���lD?�+?<�=�aF<y�"� ��uF����?�@Fl�?�	��V���?A�?���Z��=�~�>�׫>�ξ��L��?�ƽ�ʢ�	�	�%#��R�?)�?��/�Yɋ�el�N4>Z_%?�Ӿ���>�w� ������n�}�qm�=��>�_D?��r�H=�36����>5o�>Y�ܾD���dg¿�{�&a�>RI�?/�?��p�>ɞ���L�e�?�*�?7`?+�>�s��.�9����> I?�"_?!�>
4��ũ��W�>7��?�h�?l�[>��?q�s?2R�>�DýqN)��б�i�����<�B��jɌ>>˨����H��ђ�|⊿��o�>�� u>�=�s�>���ϷþS�=��ͽ�Ǿ����=&�>=�>��f>���>�0?3��>Lv�>1_�=jb���҄�������K?ٵ�?��� �m�#��<�O�=�_���?�=4?�AT��ϾT�>S�\?��?N�Z?���>g���/��Rۿ�A����,�<�K>�~�>��>b*��HK>�$վ�-C�=c�>>��>�֞�\ھ3Ձ��O����>�u!?�t�>h�=�]!?�s#?lv>O��>�7G�:�����E���>�v�>9�?�{?G�?�����4�ؐ��M[���s^���S>��x?NQ?e�>	��/՜�b���	Z��O�޽\L}?��d?���? 1�?�.F?�-B?�#z>W��,Gɾ���v�T>��!?����A��J&�x��}?�N?���>�3����սpּ���|~��� ?�(\?NA&?ԙ��(a�þB�<F�"�9�V��)�;�@D���>,�>�s��Q��=�
>vް=Tm��F6�;1f<�h�=f��>K�=W(7�l��->,?"�G��䃾��=E�r�nxD���>SL>`����^?�v=�s�{�����y���U����?A��?�j�?贽e�h�"#=?v�?p?��>=E���l޾����aw�v�x��}���>`��>(l�������י��SE��vƽ����>��>�!?*�>;8;>4��>�fe�+)��-��+9�ۣ^��h�F�8��>�8h#�1p��D��E�;����픾�©>������>g?��d>��>��>����l�>t2U>J׌>F�>�Ɓ>��i>��>��CZ½�P?��޾<�'Mܾ�骾��C?� h?/�	?��EX������f#?|a�?^�?"�J>�h��0���?h? �]�&6?��=}�<�B><�S���E2�$���>$��G\>�@��0�HD����?���> [��ץ����}����!�=���?�n0?n�H�J�|��>r��iW���O�@�g�L�����%�c�Y�禆�WD����u�2T���4��@�:?dqj?�U#�x�
�}�7��1�g���>��>�g�>j��>�Zk�M����'舿��M�=�о\?��a?GRE>I 8?i[?�JM?�]?Q�>�w�>\�̾��?$xI����>�] ?
	?/�?�,?R�?z+=?Ea�>�mR�}u�����$?G?�L?��?r�?B.�������B>�)j�,1%��C=3#>v�lЅ��5@��,>�t?d!��Z6�m����kf>h�7?�)�>0��>|j���
����<�B�>;?�l�>�� �{�q�����H�>�R�?���y��<$�7>�x�=�~� x�;��=�w׼��H=-^���
��I�<i��=�щ=�s�<�ỻ-ĉ;jڅ<:��<�t�>G�?���>�C�>^@��-� �n���e�=^Y>lS>�>�Eپ�}���$��Z�g�K^y>�w�?�z�?��f=z�=і�=�|��aU�����8������<٣?:J#?XT?S��?q�=?9j#?�>+�_M���^�������?�,,?�'�>y#�^�ʾ�ߨ�Kd3�^�?Y�?Oa��%�ʃ)��¾0�սc:>��/�^~����C���&����������?�?��@��x6�V���{��u����B?!u�>��>~�>ue)���g���? :>c?�>�Q?���>9Y?�FU?�2B?Xy���V�z뫿Iם��������>�.?v�u?O֒?X��?)�?��=>^o��:	�zs?�>�ƽ�̔��>�� 0�>���>Ti>�^�>�t�>T�>�Q���B���Z�����t�>3�?���>� ?MS8>=�v@?��!?"�ھ2��Z�To�F3H�Mb�?Aӎ?��%?�xG>�S�z�J�����>��?�g�?Y�?9��|��=��;�p����k���'?�f[>�=��,Q�>�> o�=:��>b�U�����@��O=��%?��?P>�eǿ��t��n��g��$�p<S�����W�R݊�)�V�Ͻ�=v
���#��g���~]�Wڞ��5��3����U���(|�к�>VJ�=��=e��=Nٽ<�ǲ�@ڃ<0�%=�6�<��=.vS���<�#��Kņ��䁻UgJ<Д�=O	;�d˾�H}?�I?8m+?�C?xky>z�>�+3�Rޖ>Z����?��V>Q��:��C�:����.��n>ؾ�c׾$�c�O矾�>�J�#�>�Y3>�m�=�k�<��=�t=z��=�lF���=�8�=��=1�=���=+�>�2>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�7>x%>�R�/l1�yE[�:�b�:�Y��D!?�:�8;3��>Wƽ=a�޾�ƾ�	1=�7>C�h=��/-\��љ=�{��%8=��m=��>ʒD>�~�=&�����=M=���=�PP>" ����6�"*��O0=�T�=��b>�D%>��>X%?��?f?ƃ�>,�L�X�ʾ�%��+�e>�2�=���>4���B�#>�)�>~@?��<?K@E?OA�>�'��G�>�X�>ƫ"���p�x�پ�=L��=��?ݐ�?T��>j3�=����F8!��LV�]���}~%?��(?��?���>�q�r;��#���6�v���! "��� >��G���B.�������l�I�=z�>�{�>��v>P2>W>��>��>:�I>E=sy/=p�0�ݽ��e�	��o$��}
�>r��=
j!>� �>cÑ��:<��]��$Q<���=_?>�>}��>KW�=y��>�ղ<�����sZ>V�s��O���>��þ��;�?�i�ᄿ@����4�=˫z>v��j�����>��s>�N6>��?.q?t�>��� 򾳖��>����i��
�=�&>'��JT@�+$j��]G����8?�>i�\>��=#� >��;���3�"�Z>��.�3-C�2 �>o.��н��[��~����01��|��3��=�V?$<z��2�<�*u?X?�Oy?~�>B�<[3��U!>��Ѿ+��#��ڙ���c>�(?)�#?���>��WkC��.Ǿ�$����>)L��PR���>%7�����ؾ����>k$����W4��n���%��ޓG���}���>�NG?���?��k����V������'�>_nf?{Q�>��?�o?$J�����t�ߴ�=yr?���?��?5]>��\=s��K(�>;?�f�?�?8�s?��J�J��>경�Tb>S��Cd<3�>r�>ns2>�
?�!�>Ð�>�|��,�
��dӾH� �gk���a����=�'�>ee�>�>yI[=DA.�@e=�C�=�'v>b%�>�:�>�7�>r�>ҧs�����?��=l^>�-?㧸>�N>���Ld�;�/6��8 �T���Y:��[���yK�F��=_��=�> 0ÿ��?no>O����1#?�����B����=��H>��9�� ?R�}>���>��?�г>Ly>O�>>�U>�>��gA> %�jB$��JK�uN�hj���wf>#5��B�ý����jg�NAN��Ь�
����r�#���?I�ْo�^�?����͂��:��O����?�`�><N=?�Ȋ�Ŋ�;�u�>�o�>Zn�>X��.H��%���������?3P�?�;c>��>?�W?�?˒1�3��uZ��u�d(A�"e�B�`��፿����
�=��*�_?�x?+yA?R�< :z>N��?��%�gӏ��)�>�/�$';�t@<=�+�>*���`���Ӿ��þ!8��HF>��o?:%�?qY?5TV�{����=#�-?|Z?��?#-;?�H?
AY�<?������>�]	?��>�z?~�?kM�>��>l=���,�q��Е�.��D�M��A���f	�R�i��t����x�m��W �R�8��=�M���@,�s$�=��=��H=#"�>�|�?�i�>̵>�IM?�4���A����p1�?�w>L<��̽�(�g��e�2>X]�?œ�?˚>?��A<
3\�<�T� �F>���>"�>��>���>�Pd��9��q�����=�
�>^T��*=�L9�.���z�_�X>��>���>�m|>XU��*�'>�\���z�^d>^�Q�靺�r�S���G��1�rv�RC�>+�K?��?4�=u[��Z���Cf��%)?^X<?SM?��?���=��۾��9���J��8�h�>���<���㴢�R#����:�zF�:`�s>�7��em��#�r>@���i׾�`��:�B����a<���������N־pMt����=�>����Q��[4��aز�#Q?��=3�o��PĽGZ��>;�n>�*�>�t�t�3�5�ޗ��6�=���>��a>�p�����V�0)���>U�Z?��l?-�w?7����~�JIQ�f󻾊_��@��=��E?�
�>���>hEL>����oخ�a�+�<F\����]�>I/
?�iʾo�������(2���]=�#	?�>��9?up?�O(?�a�?�
I?fG?�U�>���!��@?&?���?!�=�ԽݬT�+�8�F����><�)?��B�躗>ҏ?��?��&?ʇQ?�?��>Ϯ ��D@�>"V�>��W� _��G`>�J?��>J4Y?~ԃ?��=>��5�|颾bϩ�Wc�=�
>�2?�3#?��?���>��>Z꡾G��=l��>Q�b?F�?p?���=e�?�R1>8�>�X�=Փ�>"��>p?cO?ys?��J?���>�ȏ<(�� ;��@�s���_��s�;ų3<�u=��B�t����Ȼ�<���;�����q�����G�k��E1�;s`�>��s>"����0>�ľ�O��Y�@>qs���Q��܊�A�:��۷=���>e�?b��>�[#�F��=���>�I�>���s8(?"�?]?�o!;��b�,�ھ̯K�o�>K
B?*��=��l�������u��h=��m? �^?8�W�?%��9�b?3�]?g�r=�7�þϷb������O?��
?��G�(�>��~?E�q?��>��e��9n����Cb���j�@ж=r�>=X���d�W?�>h�7?�N�>d�b>�$�=�u۾��w�Nq��}?��?�?���?H+*>.�n�-4࿜�þB����7X?�R�>������?n��<�ڜ��N;&ͷ��������l��狾S�����3�T/���ʼ��>k�?��q?=B]?�L?,����H��l�vD��pb@�����7���&��~4��I��@��U}�����þ��@<�9���%��A�?S?V�]x�>�|Ծ�<�:Ծҹ�;�����#�&�=���2��=�`��u��ݥ��-���4?�H�>�M�>(]?Y?��؀2�^4�$5�����>�Y�>%��>·�>���n��"���9侘���LEn�k��>� m?N�N?3l?��9� -+�3q���W%�姽"���#�>��h>[M�>My�d&b��*��[A�%�i�nW�D���8�~b�K#?
 �>���>�H�?͐�>&�n���־�I,�<��<��C>��g?��>.�b>gr��I��p��>��l?���>��>՞���Y!�
�{��vʽ��>�խ>k��>��o>��,�h \�Hl������� 9�PX�=�h?�����`��>iR?F"�:I=D<k�>M�v�z�!����B{'�g>`?��=&�;>�pžL �/�{��3��vl(?[I?����(�)Ƅ>��!?fK�>��>���?y�>k&ž^�.;(�?_?�fK?n�@?���>Ւ=W���b�ɽ�J+�?M/=�9�>��X>kd=��=l���f`���'�c4=�!�==5ؼ���uIR<Y�����F<N8�<y�9>ݶֿ�=���Ծ~��4�˾��qA��n��.X`�J�`�xX¾�F���t����jcB��)���L�ʚ��s��˴�?jH�?7:(�����7����t���	�;�>������˽~�������Ǿ�����F)��Y�?���u�P�'?�����ǿ񰡿�:ܾ3! ?�A ?8�y?��6�"���8�� >8C�<-����뾭����ο@�����^?���>��/��l��>ޥ�>�X>�Hq>����螾o1�<��?5�-?��>Îr�1�ɿc���i¤<���?0�@�|A?@�(�y�쾚V=��>��	?��?>ZE1��L�����M�>�9�?���?e�M=M�W�2�	��|e?oE<�F�:aݻ��=i?�= >=���(�J>aK�>Ǘ��SA��Rܽ��4>"݅>�h"�?����^��G�<�w]>��ս<��6Մ?0{\�f���/��T���T>��T?+�>i:�=��,?T7H�`}Ͽ�\��*a?�0�?���?(�(?ۿ��ؚ>��ܾ��M?]D6?���>�d&��t����=�5�a�������&V����=C��>~�>��,����܇O��J��[��=��Y���o����V3>���>��'��e���>�>��U��S���������v��Ԫ��H$?r�;?�|�>s��=��&?�9? ��>L~s>,��϶l���>�VP���,�+�K�@���f ��ܮ���V���;�=�ľ@�̾�ȾG���1�=�O��=�eQ�Y2��*��&`��F�j,?�&>��ξl�M�/��;�ɾD쪾ɔ���:���ɾ��1���o�<��?ȰA?7�����R������
���½�mW?�D�_9�l��9�=����#�=l��>��=�御&5���S��u0?�Z?����j\��{(*>f� ��=r�+?0�?T=Z<C#�>�I%?q�*�;佣\[>��3>bգ>|��>@	>����Z۽M�?_�T?�������ڐ>(e���z���`=&/>�+5����̫[>���<��a�U��I��$��<n$W?�l�>��)�t���W��jg��?=��x?aa?�	�>�Qk?�B?5
�<
_����S�"�q�v=|�W?>i?�>�f��G�Ͼ����r�5?V�e?ѣN>��h���龜�.�nC�n6?'�n?�R?���g}�N��%��L^6?[�?`4}��������B�޾O`>�!'?j?���
?�'L?{W�>����H��
�/����?�?Y�?�G=n����=y;?J?���d!�xD��
����~>� ?���M�c�\�,�`<߽�TJ?ނ�?t�?���-b羵�>�h���5�?�0�?� ����=����\�ؾ�h���B=D�J����:�;vB�ԛξ#��h���"u;�Q�>NU@��ҽ��>��T��ڿ��̿E��_����`��?�W�>�0���ٲ���s��p� �L���N�M4��rN�>_�>����������{��r;�+:����>l���>ڹS��'��~���X5<��>"��>$��>4)��<὾�ř?�f��G@ο������� �X?Bh�?p�?Po?6w9<�v�;�{����-G?<�s?oZ?ъ%�-]���7���j?�ȫ�u`�|`4���E�I{S>5�3?l1�>��-� ��=�>�>�5>�R/�փĿ�ɶ�u���P�?X>�?���p��>8H�?�S+?���{ �������m*��х;�ZA?/3>达��!�Ir=�r)��S?��1?���z�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�#N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>iH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?� �>��?���=��>�;�=���#o.��#>�9�=G�@���?��M?���>a��=1(8�+
/�ZSF�v?R�6*�2�C���>\�a?7ZL?K�b>{=��c;1��� �_�̽��0�o��Y@���+�'�߽�]5>�E>>&>��D���Ҿ�4?��8��ѿ����G����Q?�s�>��?�!�����=�D!?#F>�l�p���飚��0�v�?��?���>�}�d\�<�=��G>��>�%�=}��13���>ó3?pϥ��nu���z��0�>�u�?�n@��?}���?���Mu��O�u�M���;M��\J>�??�����a�>%W�>�H9=��o�xܩ�fw��R�>,��?�@�?���>��_?��h�t�2�-��=S�~>��U?��?.�6<�y���&h>�t?1��|늿��	�X�l?@@�;@�S?� ��iп�Î����(�j�>�^�>�|�=����+>�@�=��=D导$~e>*�P>��S>��>f-k>#~>��<>�Ӏ��C����Pb��
�+��~���8��>���&�c�@�d�ྺ+Ͼ#!������Ǿ� ^=�v6�{�ӽ0�
��~1>�s?�c?�`?�>�>s��|�=z���+ὶ�����r>}:?��j?��Y?9�T?e�<�;��mmY�,�f� ���+X��}I>=��<�?K%�>1�>A��;�l�>�{B>s�=��>S2�=�z?=U�<�$B>Ξ�>(�>�vW>8C<>ˑ>*ϴ��1��`�h��
w��̽�?����h�J��1���9�������h�=Jb.?�{>���?пy����2H?,���L)��+�O�>_�0?�cW?6�>Z��A�T�7:>����j�`>|+ �%�l���)�7%Q>{l?S�f>�u>�3�}d8���P�5z���g|>i36?!鶾K9���u���H�bcݾgCM>�¾>cD��j�����@�qi�Ő{=�x:?5�?�H���ాޯu�pB��'GR>C8\>�Q=�x�=�XM>�Oc�_�ƽ�H�tT.=-��=Ů^>��?#�>(��="��>�P���L��3�>'�Q>N>�	<?�� ?n�7�����^ԁ�(�-���r>���>�y�>
�>>�F����=A�>��[>{�ʠW�v���NR��bP>dB���^�΍=�t�=F��l��=X�=�c���?��B/=�~?���(䈿��e���lD?S+?_ �= �F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l�6>�^%?��Ӿ
�>n㊾c풿��]�p���nZH�H�>��f?����[=�C�]$�>�ۧ>^v�Q���Bjڿ��� �?�>�?�R�?���k&����o�c�>�"�?��o?���>j��%�Q��)J>�B�>(�h?�̞>4y��?_��"?���?b�d?�+c>��?�@s?�r�>����wH.�N?���u����<�Y��"��>��>~þHA�3h���冿^mp����M�r>�J=��>,���9����a�='�������n��`�>M�>=��>@۱>�?� �>�O�>�*\=;_�C���~����K?���?B��K0n��G�<r��=_�^��$?�G4?H�[���Ͼ�ר>��\?G?[?(b�>����=���翿%~�����<j�K>�2�>�I�>�#���JK>��Ծ:5D��o�>|͗>�룼y=ھ�/��N ���C�>Ne!?t��>Ӯ=�y!?��$?��w>�o�>��E��F��0�E��>�
�>�v?�%|?�%?aͽ��H2�bS��l���n_�}A>}w?��?l��>�߉��d��r�܍�� F��/��?"ci?S�t��?W9�?g0@?j�D?�{>���Ծ��ýX�~>��!?m4�ӰA��F&�	��|?�S?���>.���>ֽL׼��~����? "\?�;&?���a��¾Fi�<y#���R�J�;v�E�9�>W`>�����{�=��>�ϰ=C.m��/6��>f<�3�=0t�>���=W@7��o����<?�5��(��!_+>jal�s�^�F��>	�>�����?6S��������&���LC�Q��?,�?��?�t<�_�kIU?��x?�N?A�;?vr�B�����
���,����9�qi���d>I �=�̾m���q6����y�����������>	-�>��?��>�� >1�>FZN��c=���w��)�m�2&���3���2��$�NW��'C���y�`�ƾ|*j��>HI��ԛ>ˈ?�=s>%>�e>&ӽ
��>�&�>r1�>Ľ>�0n>?�->��>0
=o6K�}KR?������'�p��$���=2B?�qd?�4�>�]i��������}?|��?�q�?�9v>�|h�s++�p?DA�>a���o
?�^:=~P���<*P��9��^����e��>WB׽�:��M�eqf��e
?a,?�u����̾;׽��Z��L~=�Ey?�r/?�?��/�8nw�޻<�o.\���۽��l�	�}�d3�5^������2������[8�'�2���<?�~?����5��V�۾�[����{��>���>���>�.?�e'>D�-�$��w��.���� ��>��?���>0v>?6"7?#}P?�|e?�p�>i2�>�mҾM??|oռ��:>���>e�<?��2?cK?��?8�?���=]<*"���⾣]?!�?	?��?�6?+�)���i��:�6����Q��ü�S;��i<�0���u�6a�h�>]?����<8��M���ij>�_7?d��>�U�>A���um��wp�<�[�>�f
?�0�>����8r��A�O��>��?����=�*>�D�=�2����,��e�=�Pּ�&�=�����Q;�~0<"��=Ư�=�n��Ǉt���9ܦG;#�<Wv�>^�?ꐊ>E�>�?��Ӫ �̱�]��=��X>�S>,	>�Mپ~���#����g�yUy>$u�?z�?�f=�	�=ߡ�=�w���W��>��U��<
�?-D#?1RT?���?q�=?�j#?��>�)�bL��b]�������?]!,?���>��\�ʾ:񨿎�3�|�?�\?(=a�����;)�X�¾�ս��>�[/��.~�Q���D��ꅻz�����ޛ�?3��?7A���6��w辪���?]��8�C?�!�>�[�>��>�)�O�g��$�E2;>h��>1R?��>�h?���?|�Y?�f�=��J�����D����
��qz>8
r?o��?H��?���?.��>+\�=Kv������"�����=��(�t=�#:>���>P�>{�'>�=�=]�z�d�N��f-���>��>�b?G^>r�>>+z>�����G?���>�]��v���뤾.ƃ��<��u?���?�+?�K=��t�E��G���H�>�n�?$��?Z4*?E�S�i��=��ּ�඾Y�q�%�>#ܹ>�1�>�œ=�gF=E^>o�>A��>n&�\`�(q8��TM��?4F?"��=Uȿ�m��ξ����)�v=z����~�e��hw��l�<�ͯ�tY=��ě��Ƥ�3~����׽���S�'$����>0n=s�>��=���<Pk=�:��< I�<��<8&������~�P�ڽ���?ʆ��8�;{<�\=�ք�%v˾T�}?�>I?[�+?ԹC?Hxy>�.>и3�{�>kт�tF?{yV>�_O�Zb���G;�_������%�ؾ y׾��c�Q���\>��I�\�>3>��=�&�<�V�=%Vs=�ގ=Y�T��2=c��=<@�=�n�=��=>�>�I>�Fw?}���ᘝ�L�P�ʿ�,):?Q֒>�=�ƾ}@?d+?>h.������|t���~?���?5L�?��?��h�7�>�<��:e��@��=ao����1>���=��2�jX�>��J>���ob��X����)�?�o@Y�??䋿9�Ͽ��/> �>���=�XW�YQ9��O���:�$W�	�?S1���Ⱦ��s>��c=��фپ�q�<f�a>�%�=� 潃FT��Y�=�(o�J_"=��=�E�>��H>wԡ=��[��=|��<��=�$U>d�=�Ю���E��=�w�=G)Z>��>+��>��?�a0?PXd?�7�>�n�pϾ&@��hJ�>�=�E�>l�=xtB>��>��7?5�D?Q�K?��>g��=��>��>�,���m�vl��̧�%��<s��?^Ά?xѸ>4�Q<�A�Ҡ�wg>�G,Ž�v?�R1?�k?��>��[ۿ2�,���8�٘y��D=��=�3v�'�<@�x���e�#��x��=�ē>(�>�E�>�u�>�^H>x�5>�	�>��=�Z�=�V�=XD��=��;�輅=}��L�<kcм����ٯ�:���h�`�����Ҽ��t���o�:��?>��>v�=c,�>�h�=��վET�>!6{�&G��A>dɾMXe�1&q�Wt���+�}-��>��>������t?�I>`��=��?G�v?P(2>�E��$�'����NC���/���=&�=�^z��jM���e�M;���Ծ=�>�>5�>��l>�,��?��Wu=���:e5���>�A��E���~(q��K��U響n0i����C�D?�+����=n~?ϐI?㼏?|��>�>���-ؾ�K1>�J����=���ap��X��k?�'?�T�>�4��D��ʾ����]�>(�F�N]P�'�/�0���y���]�>	q��y.Ѿ��3�m;��o���DC��u��m�>��P?��?ƺe�X����O��L��׉��?Q�h?l�>��?/?*j��ǐ뾵��5k�=Ɋm?��?���?c�>��=�I��')�>� 	?*��?d��?Гs?4y?�%��>%Ӆ;f�>F?��H��=؜>�i�=���=�P?ZQ
?=�
? 휽��	��.�ε�%p^��G�<�
�=���>B'�>0#r>S"�=�i=��=YT[>o~�>���>�?d>�̣>�6�>Vu��]�� ?q�>��}>�w!?��>�tM>R�n���bp���z�l$_�🥽T�߽�C�<w�;Ψ'>�q=���>���{�?��)>�]�])#?J��`U�iy+>��>�	�X?r�>*�>u{�>���>0�>�(|>��T>wϬ�q=�=�����,���3S�LL^���f�>"x������>�۾���3�������0���{��J��E�>��� >Tט?�b��"��	.���]��>'!�>�d?�ꋾ���Ot\>���>|~>\�従���%K�����?���?�;c>n�>;�W?�?�1��3��uZ��u��(A�0e�Q�`�|፿����
����_?��x?2yA?�V�<(:z>M��?��%�Bӏ��)�>�/�=';��<<=r+�>**����`�+�ӾX�þ+8�"HF>X�o?%�?:Y?3TV�̎<^��>.G/?�t?�?8�G?m�>?�SʾMse?�ܔ>�Y>N??�[?1#f?jF?�B>5y�=�dN�6ZL��3M�t.���$ս�׽�a��fN��)�ü�b�<��=S$>�N�<
����1>�FW��&S�=�<=<�)=ߑg>]�>
~]?q��>O�>H�7?#6�Ua8�����;/?�Y9=G肾���)Ǣ�P�1>��j?��?nHZ?��d>!�A��3C��>7k�>�s&>D\>&d�>���u�E�#�=1�>��>@�=:�L�J�����	��������<��>���>cg{>�O����'>�u��>�y���d>�Q��(��:.T���G�_�1���v�A�>��K?�?�8�=(��c��gf��)?@H<?�'M?ؚ?�ɔ=|&ܾi:���J����c�>�}�<���B���8"���:���92s>/(��ő��~ma>����<ݾ'_n�z�I�F��FJ=����R=1B�Rվ�~����=��	>H����!�N��������I?��o=(����9V��l���>!��>���>��8�8Aw�1[@�g��9��=,��>b9>L������CG�O����}>�)^?�Y�?ͼl?������v������	�������?l�?>�5�>u��>�(y>�Hھ�#���}�B�~����>�2�>z���f=<�Rَ�p�rD�ӄ�>f�?|T>]L0?�X?<�>�y?��'?�-�>��>�jżhY���a?��?0Q>LϽ�p��E�snQ��?�+!?�q�yǭ>�?w7?��D?�a?��>b�=����N�ZS�>A�>��@�~��&M�>�Q?�5y>�p?�)�?e�>�'��q�����?M>n�U>��=?d�$?1�'?��>|h�>џ������͖�>k�5?��x?bgs?_G>�4?کo>�}�>��=�͏>��?��?,�:?�AR?c[4?*��>��K=���<����=�ܣ�]0=U`�<g���|���x���N�%L?���N=��4��ս(YD��6p��t=�7�=�D�>es>6����1>��ľ�2����@>摤�Gޛ����c$;�:4�=x��>j?���>=*#����=5I�>\�>���%[(?��?��?��;U�b��@۾�#L�Y�>y�A?���=)�l�.n����u�͟e=��m?xJ^?�X�s��O�b?��]?>h��=��þz�b����g�O?<�
?3�G���>��~?f�q?U��>�e�+:n�*��Db���j�&Ѷ=\r�>LX�S�d��?�>o�7?�N�>0�b>)%�=iu۾�w��q��h?��?�?���?+*>��n�Y4�6���ą�O%?(R?0���k�?��<����ʮϽb=���-뾺|T���f�͋� Kp����H|��;��r=���>��?�Yz?�E:?'ݾsF`��!b����+}D�����������0��bJ��cs�NY�����ؾw�ܼ�|�JA���?@�(?)0�hb�>~R���O�ɾy�?>u������z�=���_1D=m�X=k�i���2����R�?2�>���>q9;?ҩZ��">�"02�v�7�V���2O->�:�>Ʀ�>���>R:���2�s�AUʾ�ن��ؽ��g>B�g?ѸU?"Or?Q��d/��L\�]�3��\����M���=6�>��i>D�}��.y���.���?�F�m��T�>��ҽ��?�=H�-?��>}Ҧ>�ڗ?p'�>���������˾PA�ab^=녪>7�z?>��>;p#>�u�
}��Z�>��q?��?�˩>��ξ�.�,�d�z�cu�>�D�>(??��>�lp�V#P�l^���v����)���f=��O?ZS����i��ǉ>=0_?V�=���=T�>1m ��8��K���&��-��=�X	?��<ɬy>�/������u��yo�?.&?�� ?�n���!���}>;�!?�o�>�4�>D/�?tC�>۫ɾ'Q;��?�$b?ӲI?z	??'X�>t�!=�k��Ƴ�>����<��>��E>�Fz=��=����z]���(��I=z��=�LԼN�ӽR������]�M<��=�h:>c%ۿ�MK��پ*{����Q
����!R��䯆�_c�6���^���T�w��E��%�N�U�s�c����l�<;�?1�?m������t���4����2�����>�yq�Ô�������F��1������
���m!�H�O��*i�®e�f�'?&����ǿ�����)ܾ�, ?�9 ?�y?���"�Z�8�7� >f�<����ĥ뾋�����ο������^?���>$��m�����>��>��X>(q>3���۞�ϕ<��?��-?/��>��r�ˏɿD�����<���?��@7qA?��(����FfW=���>��	?�?>r?1��-�|㰾c�>�3�?F��?��N=&�W�;�	��ke?>3 <��F�NXݻ���=��=zf=����tJ>�4�>����MA���ܽA�4>7օ>/�"�F��N�^��½<3^]>��ս�A���ބ?�P\���e��/�����sG>*7U?Zq�>���=�-?�H�V�Ͽ��\�S�`?x1�?Q��?�*)?���(��>t"ݾ��M?p[6?�k�>Z�&���t����=Y�C5��wh�v�V�3�=�t�>��>«,������P�쒤�as�=x��n^ƿ��&�i��=�=g��:�0�^�������'�N.��}gi��̽��=_��=z�T>�
�>�M>�F`>��S?s�n?���>�D>Jv���_&վ���;��#���Ɔ�Y6�����D������G�Ԩ���ʾ�=�"Ѝ=�6R������� ��b���F���.?P�$>k�ʾ��M��!.<�gʾӮ�� ����ۥ��-̾�1�Mn�7̟?t�A?X���	�V�� ��N�Kr��s�W?�?�����ꬾj��=�ϱ�W�=+�>Qz�=���3�"wS��5/?�?�j���O��b�%>���'�=&7*?.&�>���;���>�Y%?��1���ܽ-d]>��5>��>_;�>�>j���6B�(?9�R?���w���>Sʻ��7l�S�l=�.>o~6�(���;B\>���<8���^Q�A�}�d��<�(W?x��>��)�A�a�����yW==޲x?��?v-�>g{k?��B?T�<�g����S� �\w=��W?�*i?!�>&���	
о聧�G�5?:�e?��N>�bh������.�U�{$?2�n?_?R}���v}�Q������n6?)�?��M��򞿐��N�	�$��>y��>b�(?��(�5�>�2r?Ћ�(O��yK̿u��4�?��
@�U @z���*�����?i�?������	>���L�2�m1?=㢾������=��C�u�\?f3�?8/?�"��ѕ��>(N@���?{K�?�ݭ�f#���	�IUi�}r	��U��+�=珯<Ԅƽ ��́6�DK��?$���)��w�̼.�t>��@�s��q�>¤�h��=�ƿ$㎿�dྲc�%?�Q�>~zV�oO��t@w��d�IB@�KF?��TV��>��>X������:P{��9;��ܛ�&�>;T ���>mU� յ��!���lS<�9�>o��>���>���{���:ə?Z���qFοc�����X?�d�?�x�?H�?w�7<�w�dr{�b���(G?Zs?��Y?d�%�/D\���4�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�P_?��b�-�p���,�������>��.��Z���˼(t���e�y���v��5�?��?���?~�4�"���$?�;�>����MHɾ[7�<i0�>^�>�%Q>X�N��|w>�����:��>���?k�?K?U7�������p>�}?���>�v�?��=���>��=�ΰ���G��� ><�=��C���?�zM?���>�H�=e9���.��aF�:�R��,��UC�n�>
b?�fK?Sa>�R��{>�_� �%̽2������n?���0�� 彝1>��:>A->`E�q[Ҿ�`6?�p辎lڿ�ﯿ���<�P�?\��<�R3?~Ze���w�k>?�]?g�3?����Τ�7ӆ���b�4��?� @E�
?���sf<�&�<���>^n�>H� �7�P���I�'0{>��B?Q���kC��H��8ٝ>=^�?��
@:��?E̓�UT?Z{���<��� �����D+�g�z=Z�J?@�о�ZV>g�?ɖ�=�VZ�]p��k�N��>�?H��?Sy�>��e?�&t��3)��7�=1v�>O=?v�?�� =5�lDI>e?�6#��;��}���h?ɐ@�@RW?鄮�4O׿{䖿^얾����\}v>�~�=�7!>��۽Mi<l�M�N9B�d���>OĬ>�o>�Yj>�c>��
>8->����.!��&������?�=���{������T�����` �����Ծ�۬�?�ν�v̽�>U�t� �@]�;ӛ�='�\?�lY?�eb?5�>���Y��=�޾#��=N:=��s�=~Ǆ>+?T?jB4?#�=驝�UF_�4怿-���P�v�Q��>�">)t�>6�>�r�>16	=q�s>�V=>ݱv>1��=��T=��;��q=&�b>�h�>��>�d�>2C<>`�>6ϴ��1����h�=
w�}̽�?���{�J��1��=9�����]n�=_b.?M|>����>п$����2H?�����)�#�+���>k�0?�cW?��>h����T��9>N����j��`>�+ �;l�t�)��&Q>�l?e2e>8�l>�I2��a2���O����z%p>X�2?����Y�?�U�u�HlD�ؖپ��Q>S޺>fS��b���.�}��Gi��=�*;?�q�>�b���벾�H������^T>��X>7n=
��=��D>���f㽟�N�&R=Z^�=ka>J�?A>��s=޲�>\����8��Ƥ>�8>��/>��4?*�?�]��n����4h���\5w>�v�>��v>�1�=5�F��o�=s��>�zZ>�/���_������B��Ig>?G���US��xy�v�=�G��t�=RV=��	���<���E=�~?�����爿�����)fD?�;?7��=H�O<W"�I����,�����?z�@�f�?bo	�ߏV���?7�? ������=�B�>��>'5ξTlL�۷?��ŽŢ�K�	�#��@�?f��?��0�����l�;)>Y%?��Ӿ0��>�~� X������[I�(J>`Y�>��h?�?��U�H��Q�Jj$?FNE?�0ǾnH���(̿݁�4@�>J&�?
ː?��;�+����s��?@��?k�9?��>nʾ�E�����>gF1?�?�H�>z�����8����>���?���?��W>�ڒ?y-x?j�>�����I������퐿�`�=o�ýW��>��=���(m.�/����s�ˑ?�c�從Q>�L,����>9h�
�澿%K���s㏾�@Ƽ5�>�G�>^�=>Je�>?�>��>���<%���䑽�:��i]��K?���?R��R!n�m�<�!�=�*_�:?k\4?b�^���Ͼ�Ш>ԫ\?�΀?W![?�c�>���1���޿�s����<��K>���>X6�>�����%K>�Ծ^�C�Sg�>٭�>�|���ھ���Z��1b�>�d!?���>�a�=�]?�+ ?66`>|��>��D�q���Z�E����>)M�>Ċ?�4w?ϟ?�{��[3�;$��Z꡿�]���5>y?�c?<��>W��N���Cm����� �V�?�\?��9?��?IZH??�<?�]^>��,�eӾh�%��>� ?���C��"�&?�}?�`?��>u�y�oPý8q�{k����|�?͚[?^�%?"��2<_�����a��<��Z_��!�?<�����D>H�>����
��=�>P��=$m���4��<�H�=��>���=l"7�@���b}>?���]�u-,<�����'��t�>�Ǩ>��O�#�?�3������{���?��ض�=q��?�_�?���?�K�;�D��A�5?�Z?a�>?�I�>�!��U!	��4���҇� l���:�2�>�->�F�=��X��6;��c������|�?�,?�f?��?8>�y�>��(�F�Ӈ��f-��$N�B�	��&*�)�����g��љ�v���|���F�,י>&�dUz>�	�>/S>1��>�>�n�+@|>��=��o>P��>
��>KV>A��=�����.z�MR?�����(��N�dS���B?�td?� �>ua�1��N�UE?�p�?2p�?إv>�g�-�*�*?0=�>Ϩ��
?a?=���*��<R^��P��f���@���>�@ֽ��9���L��f��

?��?�.��l*;^7ؽ|���T4=��z?�f,?��&�"-O�yt�-�R���7�Nu�U\������8��b��썿<ހ� �I/�i=�<B3!?V[�?�r���5����c��;��Pi>h��>$��>��>�9>(w�}�9���b��)��Z��DT�>@~?gɋ>�E?�t7?c�N?mC?"�>+�>8���b�>�5�b�>�"�>��0?7,?ZH0?��?�*?�pm>{��K���y�۾��?O�?џ?xr?��>;����`��q���ﻎ���x��e=3��<�,߽qk{�B|=TXc>�;?�����8������j>�q7?���>*��>�w���À���<<��>�
?誏>�����5r��F�|!�>S��?�i���=��)>"R�=L����tܺX��=u�żpP�=8��c?;�0a<Gq�=c�=a���̈́n����:��;p��<hs�>�?ј�>VD�>EA��K� ����B�=�Y>PS>�>�Bپc~��B#����g��Sy>�u�?�x�?��f=��=ѐ�=/}���X��/�����J��<ݢ?�K#?6XT?���?��=?hi#?b�>/,�mL��*]�������?d!,?׊�>���7�ʾ��ȉ3���?I[?X<a�^���;)���¾��Խ�>�[/�S/~����KD�d������-~��*��?ʿ�?�A�U�6�y�ȿ���[��_�C?�!�>Y�>M�>b�)���g�w%�C1;>ӊ�>_R?��>�P?x|?kZ?��U>̽8�7���0��mj��(�>K�??�<�?�Q�?�Sz?W�>�>�U+�i����^ �<�|��y�C=��Z>��>��>���>8>�=0�ƽuᱽ,d>����=��b>���>�y�>��>�#|>��<��G?��>�_��O���ꤾ�Ã�p�<�ڜu?���?
�+?�B=
����E��B��FK�>�n�?��?Z3*?z�S�W��=_�ּ	㶾�q��!�>�۹>�3�>�̓=}F=`>�>���>�(��`��p8�NM���?�F?C��=b�ƿ6mi�<eK��<��i�]=���O���T�t�H��=�,���Y���|���(�9ޓ�C���䧾ڂ��[ D�k&?�/y���s={3>�ƺ=��3=��="&=��A����=�伽�,=\��;O^W��Sν&U�:ۚ;.��X6b�G�Ⱦ3~|?��F?�R+?-OC?f�u>�>13A�j��>B(���3?�X>�:u������!;�7�������j�ؾ�tھ�fe����t@>�-J��\
>.P4>v��=1�<�"�=��_=�#�=��^;��+=�%�=���=�1�=\�=�>��>�҂?�9q�C˕���W��tV�H�6?���>�^i>I'¾i�\?�@�>6ޜ�Is��<�4��,�?��@���?ű/?(���l> -�����=�i$>V���u�X=��>Mڛ����>�}�>�L�����Fý���?���?:2F?��(Ͽe��>v�>>� $>�J����-'�»^�C��B�?��\�*����i>в2>�=�BQ��A��<Fw;>Na�=�����a��I�<?���>Ede=5�3>&�g>�=]����>��<�B>Z��>��=�f�=R�0=ќ�=n��=j��>n}>>x��>x�?�^0?MRd?-+�>-	n�%Ͼ+/��#C�>z��=�A�>�
�=�XB>��>��7?.�D?~�K?(}�>t�=���>��>G�,��m��j�Ǯ���!�<|��?�І?PӸ>v�Q<�A�ϓ��]>�C�Ľns?M1?�o?��>~X
�y�����׾;�r�~=l"���3�����&�Xn����=:E�$�'=�P�>�k�>(_>��T>��=DÅ>��>��=h����=6�ܼ�+b<��>!�=��8��&�=]/*=����ѿ���������8�8=���~�Y<�d��nT>4��>��_=2f�><�f=���Y�`>��q���_��I�=�z���2@�3y�]�z��A�5S�
\[>;t)>4��5׍���>�˩=�L>i��?��Y?��=l����4D�������L�=s?�=��4> K��WL�"M���U�J��y�>�ԏ>N�>��n>{�+�?�O�|=�9�7f5���>(���o��n[��q�DD���矿_�h�"�U��D? ����=K�}?��I?��?(��>��&�ؾ�~,>�x����<��wCo��H��z�?��&?���>�X��D�nG̾���F޷>(?I��O�a�ɰ0�Ը�4ʷ�쏱>]���%�о�#3�lg������-�B�OPr���>�O?E�?6b��W���VO���� ��r?�}g?��>;J?�A?�!���v�=s���s�=$�n?��?.=�?
>���=g�	���>��??	ޏ?�pu?�&��|�>D�=�)>�冽z]�=�Z2>��=���=�>	?1&?��?�=y��)��]���G��mu�l�"=�w�=F˗>~t�>,�`>��={�@=XՐ=� L>�`�>5x�>#�a>,��>؍>G��0c<�Ԋ�>-�)>!j?��?џ�>���<cE;A]~>R9G��[�����,�>!!6=�'�=�=���+影�(?u7пY�7?;��>}t޾*?*n���>��	?9��>i
��栲>�t�>1h�>K�>�@i>MX�=sː>>�>Wq��m��=���p&�V�?���M�����5�?>UN�Jo�rV���u��.;��ն�f��UPi�ԃ�^kE�+�=���?�U��c��xP���潦�?�.�>1J?R㌾��N��v>���>"��>n�����댿�;�t�?��?�<c>� �>$�W?u�?��1�3 3�	tZ�?�u�Z*A��e�9�`�rݍ�蜁��
�t(��6�_?�x?ttA?�^�<�4z>���?�%��ӏ�)�>#/��);�c�;=K'�>4 ���`�#�Ӿ��þ�1��*F>�o?{!�?tU?�FV��{d���">/9?�m1?z�p?��2?�^:?�d��$?L7/>}7?0F
?��2?y|.?r?;�3>���=8d�9�%=r��������D�����
>��ȚC=��y=����\^<��=ζ�<�����s��[���Ӽ1��<5/=5k�=��=���>Y�]?��>z��>�7?�v��I8�]���L�.?�-7=|����Ȋ�V���8��,F>	�j?@�?~NZ?!�c>`�A��AC�8>�K�>m�%>t�\>6�>�(��D�43�=�]>�>cϦ=lM������	�js��R��<1�>e��>�->���Jz>�j��3�h��g\>�M�����KE+�^oJ�^z$���\���>�B?�O?��C=r�ZE���*\�
^7?��<?�>?(�p?�9�<l����<�E��5m��>�w�=����ܛ��㟿f�@�"�g���
>���Q���kB>>�еѾ�Kd�țL����QM;=���~8=	
���ǾDtb�v��=�D�=+�þv�#�m锿���K?�=*���B�,�X���8|>��>�ĵ>�&���Ie���<��Ŵ��1>=m�>�CV>>�����侎�A���
��+�>g}D?��^?y}�?�~�h�p��jB����������Z�?\�>��?��E>�b�=3E��=n��He�p�G�6�>�>m��ZG��ᠾ�x󾬐#�3��>�?:�#>��?[�P?�Y?��`?� )?gs?HE�>]����I��3�#?��?��=� ���O�6�8��v@�}�>�c,?�s���>#?vj?v�"?VKW?�w?Y>����H�?�q�>0��>�P�X���K$h>��A?`��>�Y?�\�?��I>�4�Y�������է=�?->�O,?V�!?4�?9ܾ>X?n�ʾ%��Љ?9�?h�?�ua?#>��$?lР>C��>���>!�>S�$?0)(?��1?�#V?�0?C�>O�=��ڼW*��N����⼡��<߿=��#>�.���սm*����=Wg�=���<�c������^:=��~=��=]�>��s>�����0>y�ľ7I����@>�w���J��`܊�Ձ:��ַ=��>��?���>lE#����=ʥ�>�4�>���2(?��??o�;(�b���ھ��K�X�>�B?��=��l�����P�u��Ch=2�m?ň^?�W���M�b?��]?3h��=��þv�b�ŉ�\�O?>�
?L�G���>��~?^�q?[��>��e�):n�(���Cb���j�-Ѷ=Mr�>MX�I�d��?�>l�7?�N�>6�b>�$�=du۾�w��q��k?�?�?���?+*>��n�W4����ِ��;?�9�>�T��[�?��$���ɾ�X�����"羝u�����07�����j2(�e�������n�<5�?�qx?U8y?��I?�����{S��3R�����a�T����A���-X�r�A��F��Cw�/��;Q�C}��j�=iNU�[)��T�?c?��Y��?���D���ǾR��=e����)�N�<���6�=R�>f8��򽞵���e?�Z�>���>�;?�P�50��4�j�S��Ծ�m>-B�>5�w>%��>q��=[���O�^�پOͽ�Gʑ<���>s:_?z;?�b?�k2�5'�� ��S�>�w��<X�mE����'>i�>���k�ŋ!��(�F�N��Yվ8�8��<�A����`?ru�>���>pԕ?�-?�v1�t?��׺�Q�񾟱>|�a=��K?#P�>dl{>S�e��w7�W��>�l?,��>�Π>�猾�<!��*|���ͽ�w�>g٬>�E�>�o><]-�F�[��A���r���9�~X�=ݠh?	@����a��h�>�(R?��:8LH<w>�>iEt�� "��򾤼(��7>M�?���=&J<>{Lž�ȁ{� S��Ol+?��?9l����K?�>^U"?���>̔�>��?5��>G[���XP=�?>b?p�N?M<?��>W�=ܣ��.�����^i�<�,�>�b>�)�=zM�=W����T��]*�e2�;�;�=�)3���������C�!�=�>n=a�I>�6ۿMoK�Q�۾����~���
�qȉ�.�������
�Ǽ��.���kt�@��S�3��vW���f��P��
@m����?�~�?`���U���y͙�)��$���('�>�<s�]*�����W��������E����� ��N���h��8e�@�'?�����ǿ갡��:ܾ#! ?�A ?0�y?��3�"���8��� >�A�<u.����뾬���	�οL�����^?���>��N/��j��>ʥ�>�X>�Hq>����螾K2�<��?.�-?��>�r�5�ɿ^����ä<���?-�@�A?`�(����k�Y=@T�>��	?��?>�.1�p��:8����>\I�?���?JR=�^W�˪��=e?A�;|�F���ƻ*L�=��=W�=�L�Q|J>;C�>����A���۽��3>Q�>q� ���BG^�.�<��]>=�ԽN��W�?��`�A�]��;0����L<>|�h?���>�p�=��>?c;�� ӿU2Z���F?tC�?���?�:?�ڕ��V�>ǧ쾅�U?��;?�Ǚ>;�1��sw����=�㱽��<�G㾸gn��w�=߲�>`U3>�^K���8Y��ˌd� n>Xb�h'ƿ�(�E���$=՞^��$p�l��B����*j��롾��b�3�׽T�f=���=ʯH>w�{>�BM>��K>��T?��k?bi�>_>��㽟����R̾]���M	��+�#��ۍ�ã2����$��Β�	 ��c�g���Ⱦ\�O�Sk<t�_�C[���P�n�� I���?�B>����ø>����=
>������C|�'�罺�TL-�g�J����?i�$?���W�6ƾ�8��>k��GU?�B���!����v<�`���ռ=/�>�I�=�@��ԏ%�i�b��f0?�e?g8���4���!*>�� ��S=,�+?B�?��\<�>n8%?��*��#佃�[>W�3>oѣ>N��>��>���)۽<�?boT?���Iќ�`��>nh���\z�#a=�>6�4�1�� �[>��<��T����oѿ<�(W?��>��)����D���q��k==��x?x�?�B�>+uk?L�B?��<�J����S����!w=ܿW?!#i?��>ϳ���о�n��B�5?9�e?q�N>�sh����;�.��W��(?5�n?�_?&3��+u}���l��(m6?q��?�dt������1�q��&B?�4?�'?�^%���_>_<�?Cі���r��ǿ�W,�怡?�Z	@��@����{��F�[�D��>�c?߳��_2��
=쟾�*>��6?w?���b����P��!L�9�q?n
�?w3?�g���y	�>�/���?��o?�߾���=cA�[?��A �����r�=[\���b���¾����������|���,\<�<�>��@����>
�L�3?翨������{�s��OK�p�?�xf>f!��|ܑ=�uY�䆿��F���^��?�x/�>�f>� ���ؑ���{��a;��f���>���J)�>P}S�ҵ�-U���I:<��>ʏ�>���>�p�������Ǚ?�����Hο�����y�5�X?�U�?�_�?�j?{w=<��v��7{�����+G?҅s?� Z?}�%��]�ݵ8�&�j?�_��yU`��4�sHE��U>�"3?�B�>T�-�-�|=�>���>"g>�#/�y�Ŀ�ٶ�8���[��?��?�o���>q��?ts+?�i�8���[����*���+��<A?�2>���K�!�E0=�QҒ�Ǽ
?Z~0?{�i.��_?ȭa���p�*V-��K½�e�>�K0��%\�@��~<�ze�0���>x����??�?�?V+���"�� %?�e�>�����?Ⱦ��<�Ƨ>��>�tM>j~c�#�u>�����:�_�
>pp�?%N�?o[?X����Ǧ�$�>��}?t1�>��?�9�=_��>#��=����1��,#>���=.?��k?�M?�0�>���=�C8���.��?F�gNR��B���C��$�>��a?SDL?6�a><��;61��� ��̽`�0���(0@��A*���޽)*5>�5>>��>��D���Ҿ\4?�'.�KjԿ�m�����E�c?���>�?���5\���R�>�lM?F�>"�&��n���N���?���)�?���?�??$þ,���F0>J��>$�>��@������D�=�{<�A?%�c��\���Y����~>Ѿ�?��@Iد?|�~�É?����������<���!����=��9?��Hj>l� ?�c�=n�q�B4��ωt�n�>��?y��?�)�>e*k?Y�m��Q@��{k=�8�>K�e?T�?E�:M��~eI>�?t��X1���d�,�f? G@�@=G]?ʩ��>�ؿ�鉿�໾�����G�j�E<Ro>��彣�= > �(�-��<��>�>&5~=ƫ=�>�=>�:=%>(>�_��c������^ԕ���K���5�v�$����S{&��˽[g���������l�9y��c�u���sٗ��T+>H�r>�8?$�H?�`~?'T?3>��>E����|Q�=�mU����а�>�?�	8?��=?��=�R���h����������9��>Q;���	�=[h6>l�>B�P>-Ѥ>�D�>C.�>�M�<���=|��=��=(X�>H��>���>cwu>`B<>ې>Uϴ��1��$�h��w��̽�?T���0�J��1��49��T���Oi�=b.?�{>����>п>����2H?o����)���+�B�>p�0?�cW?˝>A����T��9>���4�j��`>�* �8l�u�)��%Q> l?�H>Pfs>F�-���2��I�c(���fa>	^3?�wʾ+}7�'�u���I����c�/>o��>����&��f��Q{��\��W�=�89?���>�lɽ�N���ކ�w����U>"T>��<5��=Ǽ6>�9���ٽ�*L���<@M�=��w>�t?�A6>�ä=��>���K�P��>��K>l�6>rG@?�!%?���(��끾��-7|>���>S�}>e@�=�I����=���>�6^>�w߼��}��)���?��b>�Qq�ޖh���Y��z=�\����=>�=W���ڋ4�4-Z=!�~?�n��$׈����u㩽r�D?"�?h��=�<�� �����	_��C��?��@�m�?�	���U��T?8�?�Қ�Mq�=#��>b�>�t;��K�'�?*ݿ�����	�b�%���?�Ơ?�l*�����l�R�>7�%?MҾ�S�>m䅾h;��SД�=2p��n�=C�>R�o?�����=$p=���>��?1���?����ſ�;8���?�p�?���?�0e��έ�Tz�R(�>�_�?_�k?e�F>��������v��>�@?z `?f�>���k�7�@ ?P�?��P?+�X>Dc�?�6{?��x>5E��{� ��������E�>x��TkX>Z�����V�ƿ�~Vb��h��=�u��>
��<��>�N&�T ���A>ഷ�����'3���?<6�����=gt�>��?:W�>*:[>.���߄���(F�"�$�{�K?%��?���rn�l�<�j�=A�^�I$?"G4?[4Y��ϾXШ>׮\?Q��?o	[?�j�>=���9���⿿y���z�<8�K>{�>_)�>P���+QK>��Ծ��C��s�>�ߗ>5L���Kھ6J��"흻B�>�a!?~��>�=�� ?��#?��j>�"�>�aE�;����E�!��>+��>�L?�~?��?�й��[3�	��硿#�[��8N>��x?Y?�Õ>����������E�3�H�\�����?�ug?�X��
?�2�?�??D�A?27f>`����׾Lm��=�>x�!?�����A��B&����|?�[?���>�����ֽ�HּL��_u����?[
\?�8&?ٌ��a��Cþ<�<*�%�L1L�w��;`�K��>QG>�臽�=�>s|�=�rm�k6��-e<��=ܠ�>N\�=�6��K��^�5?=��	h��Л;A���r+���>��S>��y�kl?�'��Y�������������ɽdg�?���?�?�O�=����*rl?}io?�S?ό?���2��A��d����m�#���>*��>oW=�&��Ϊ��ů���v�q�e��� ��G�>�G�>�h	?@N?gL>)K�>�ǘ�fw*�$����y��"Y��A��6��E,����(\��!�+�����s����m��3�>񞜽���>�n?�Wa>b>�>���>��0��>�Q>��s>���>�Y>�n0>T��=���:�޽MLR?����̾'�ְ�٪���3B?Hpd?�/�>�h���������?5��?�s�?�Cv>}h��++��l?	=�>����o
?8:=���`W�<DT��۸��.��%�ʪ�>O׽�:�8M�3jf�Ai
?=-?������̾~5׽��þ�p=rTp?�Y?�����Z�\�v�,g*���r���'�RbǾz�˾0�7���v�����b腿���%g.��x�=V7?KOZ?kL���Ⱦ����]�ɩ4��Q.>(.�>�=�>q�>��*>�����p8�� ��!���'�{��>�Ƀ?�~�>�U?g�H?�C?|V?�Q>��r>ot�8�*?��X=r�D>�!?�C,? $?}ST?�f?m7?7�E>�<���������k�>�?�_/?�~?r ?u��\z�Y�,�|���hؒ�;�=1�>�1T����缍��+c=��j>�?Ql���8�i����l>	�7?(��>���>���WY��8c�<Y�>U�
?�6�>("��(Cr�}��1�>���?<W���=*>ץ�=����y�ǺsY�=�[��峏=�(��P�=���!<�U�=m�=�����y�x+;P�;L�<Ur�>��?���>�?�>E���� ���NJ�=�Y>�S>�>Hپ�}���#��
�g�hy>�v�?�y�?��f=W!�=���=�u���N����r�����<f�?tH#?�WT?���?��=?f#?��>�(�gM��^�������?1,?]��>���ˬʾ�y�3�[�?�Y?I@a�?���?)�)�¾Q/ս�>g^/�T0~����D�<������c���ޙ�?���?�KA�j�6�Hy�E����Y��#�C?�>�R�>�>3�)�%�g�I%�nN;>ˊ�>fR?���>��T?	�{?H�U?2;>5�{���U��2hj<�/�=�9?�2}?l/�? \z?��>\>� .�2a۾-��4X��l������u�=��d>��>{q�>�>�{~=H�Ͻ�eٽO�2��F�=�I>���>fݢ>��>m�l>0TI<��G?���>�2������ܤ�у���<���u?��?��+?�=�w��E�	5���q�>'i�?f�?&*?7�S�(��=c1ּY׶���q�m/�>�ӹ>e'�>hȓ=��G=�W>���>F��>5�W��c8�d�M���?�F?�%�=@�����b������t��� ~p�Gv����b6�GZҾ���>�n�ܛ2�#��B���u�*�9  ��`��iC�>mpH>��>~�=@_��T��z��;��>��`�O�O�Vi��D�*��8�%��ջe������6��<ű �žf�~?�7?��?6�A??Z�>tf>����u7>���?��S>��t��.ľk�O�o���ǈ����Ͼh����c�+Ɛ���=_ν(d�=��,>���=�=)��=M�(=�M=�%�::�=Lʬ=.�=Ǻ�=�!�=LH>��=��?����T;�N�ėI���@?���>8�T>�ϣ�2]? q�>����W���eV(�^;�?c� @��?�-?�E�<�i>~\���=�2�=�Ѡ�M�_=T��>�;��:�>u��>rtI��������p߿?���?^�G?;r���ͿG�>�n>��0>O\L���0�q�A���?���֞?�NB�ܾO��>�?�=Q�ݾNAо���<�B>{fF=�\�aEg�%3�=�쮽i�w=�<�C>w�Q>�8;=0G���=�]=��=d�!>d�)���l���ʻ�/�=z��=��>��)>���>2�?ۯ5?��`?���>{C{�|�̾�
��}��>P��=�	�>lwr=3&<>��>�w>?z�A?@?}��>׈~<t�>���>�����i��C׾'紾Q�8=��?���?@K�>)o==�[��"���F��j3��
?;�.?'?�z�>�U���࿫Z&�m�.����g�`�D+=Kkr��RU�%����m�	�㽐�=�p�>d��>��> Qy>\�9>�N>�>�>HO�<Er�=��]ǵ<�����=·��U�<d�żD���h!'�)�+�	���w��;���;��]<I<�;�V�=�u�>nر=	 �>DF�=+�r�܎>y���?;�g�hJ��Vt3�ûU���v�;>.������^>��>5�E�1���71#?;f.>���="f�?Ufd?1�=��W��(��R������k��=�`�=8 ;>7���zh�?`w��h��9�D��>���>��>��l>,�#?�C�w=)��a5�;�>�|��b��)-��8q��?������$i��ӺĠD?PF��!��=�!~?ǰI?5�?	��>���g�ؾ�<0>I���=��+q��a��Z�?�'?^��>��Y�D��!ξ0��n0�>��=��G�������2�-E�=d*��?�8�������7���'��5�\�V P��R|>�Jq?�s�?��wKf��vm����G���/?@G�?���>Bc?z=?J5|=G��X�O6>zB?ͣ�?lu�?g��>YL	>|/�!��>�^?��?4��?l�g?!o	���?��=��>b�*=��(>��u>%>{�>c��>
]�>7 �>�g�<%������8о��6�f�%= 	�<��_>�<�>���>���=�d>��=�P>Y�>[�j>>�Z�>���>J��~P�B�?m�=o"�>�~@?�k�>C�=�a3�
F*��w��:�ӽ
�'���w�_���'>n��<�=J�A�a�>t���t?�TQ>�6���?�h!���E��y�>bڅ>����!O�>�a�=s�>ܨ�>�r�>k�=��>"�d>Am��>tw���#�9C���R��{о�Pr>�]��:M�;�L^�#�?��<��u����j������k>�X}=f7�?*`	�Sh�/(���h�?�c�>��/?�����&t� �>-��>T�>S���ʔ��挿e�侭P�?�,�?Y�`>f�>L6W?{w?ç:�7���Y�>hu��@�Uhe�C^^�Bd��cZ���
�=���`?�Qw?��A?�;Y:|>w?B� ��?��?&�>(�,�(�<��<Y�>`'��ZW^��*վPPž����%I>�k?�??Y�E��	e�8�9>��N?H�C?�@�?�z(?�C?սl��}.?'eE>�}�>h?uP3?�!8?$�*?uL>��1>6d<N��=�_K�R��Up4���ʽ(v���7 >�*> �>i؂=�h�=WGx=4�g�f:::S�=*���U�=���<�Ħ=�D<Xw�>�0^?���>�>7?{�\�7��骾Gs0?gJ=GQ��Fy���,����ﾁ><%j?^'�?d Y?�c>��A��OB��w>�>9*>��]>��>z���?�A�	�~=w�>d�>|a�=�A����e�	�񑏾"��<X�$>���>�W|>c'��%�'>北�3�y�d�d>�0R�����a�S���G���1�Ǻv�v��>�K?G�?Ob�=���]9��Q\f� R)?^0<?�<M?�
�?2��=aܾ�:���J�1<��a�>b��<���g���Q%��5;���K9��r>ȟ��T����P>���\ݾ�&f��+B�����=�0�B��<!�>ھ5�ߴ=j4�=�ƾ��$��|��^Q���gF?�=H���W�W���4�>���>kֹ>���X�v�C�WO����=���>��>�������RD������>M�T?9�P?��2?��M�c�r�����?��Cg=#:�;y#�>�X�>�	? �>��>�,�����J�oL����>���>�Ͼ �2��b˾s@��i:�`�c>�!�>��>��-?	5a?gH?��a?�'<?��?�c>Qb��}��Pb,?&�?�=����Լ��)��l7����>�p7?NHm��j�>��J?�	<?��C?q?��?�$>�T���[����>�*>z��暐��³>�wQ?۳\>�o?ʏL?�>0�/�ۇ��Y�(�.Tۼ!�=V��>��>=�>�x>��?v(��nǽk�>l�?���?A�~?6�>��?�ت>��?Z>�h�>.
?�?n?/�[?�(?�$�>6�8�����оּ�Z뽾#��w�����t=è�<cK��)���ʽ0�9�=0�;]!½���>���Z!�4V��>|b�>��s>���=1>?�ľ�F��g�@>�ۣ�E���Պ��{:����=8��>-�?1��>�Y#����=a��>�F�>D��4(?��? ?8T!;`�b���ھ�K�+�>
B?���=G�l�b�����u��
h=��m?��^?=�W������b?$�]?�X�=��þh�b���龚�O?�
?��G�Q�>��~?��q?V��>��e��1n�����Ab�J�j��Ѷ=}i�>xV�;�d�]7�>+�7?G�>x�b>��=]q۾��w��U���?��?��?���?�*>O�n�A/࿶�����T�o?N"�>�	ľ��@?�5���V�K��ѻ�ƥ����n��K�¾�,���c�OFJ��(��3�!��?͆�? �^?�ӂ?���b�j���@�����*;�%�Ⱦ�G�IM6��!N�!d/�yo����\�޾ǅ���>�s�͠@���?,^'?�Z��.?���2�����ZI>{߅��O8�g�㼗���Һ�d9�=6�<�8I���0���c?O��>8�>��N?��]�p�B�j�#�0W@���� �d>{ t>/rg>�<�>����[��gԽQVɾ����T���_>s_?0cP?U�q?��0�g��qo�:.�b@�<,M��?�=�(>�s>8F]�p�/�e`/�XC�r,u�6��֋��:����K=L�?
ɤ>���>�ј?�J
?��
�hb¾���#d%�>	8<�>l?m��>+�>�u��-�Wκ>u^?�~?d��>v#оQ���p�
o{�(5�>�6�>*�>%�,>��A��KZ��������yT:�� D=�o?��.��gk>�7?4e=5��=�Ϻ>ͱI������s��^p�=�Y>
��>T��=rZ{>�M��
���{�	ߠ�0?W�?
��{��*��>�W)?���>�O�>���?�P�>�M����z=��?r?b?\N?�.?Fz�>��9�������P�*�O㤼��>*�n>��=V�>�+'�]���a���</=�	K���Iu�������
(�^~�=�Q�>5XۿP�K��V۾6��]�f�ϕ������n(�����9��W˚��z�h���d-��U��b�lY����n�<��?��?�9��H�������������*x�>'1t�|Ђ���v�>���gB�=>���>!���O�Vi��Te���'?������ǿ۰���:ܾ! ?�A ?�y?��;�"��8�� >2B�<�5���뾫����ο������^?���>v��-��p��>6��>1�X>�Hq>����螾V8�<��?��-?'��>F�r�"�ɿD������<���?"�@�AB?r&%�~6���=���>q?�o=>�c3��t� 茶�?�>z��?���?2�}=ZBR����*�d?�&w:��H��\R::�=�`j=$&=\���S>@�>u� � �L�����$>k�y>[nH�C���i�(�l<vkY>/ ���z���?1�]��se�U1��=����>`�Y?J��>��=�r-?�E���Ͽ��^��\?��?;@�?�-?�s��#��>�K߾�O?R&9?s��>��)�?{v����=5z�<�6ܾ�o[�'P�=���>ڪ+><�,�{��b�b������=����$ȿ\)K����/�=@�y>�H����~�F7�a���]8;�����z>��֞=�=��V>xX�>�d�=���=��_?̙}?y��>���=�0���ϑ�����^ؽEh���N����_��F��V���Ж1�nR߾��쾚`���6��M�1=�nZ�=�R�܂��	� ���b���F���.?�v#>_J˾��M�i&<)�ʾߪ�X���䦽�p̾��1��n����?B�A?�υ���V�D�?�r"��|�W?G�G���4��_��=ꬼκ=���>�V�='���3��^S�OE1?� ?�\��i����1E>�,�W��<ކ*?W}�>e	;r��>�(?a���ߺ�MXi>�#(>+�>�>�>U�>6,����ν?�?�L?��|�����>qu��,FS4=N#>�+�6{���JF>�'<3��C���z�{���,=gW?��>L�)�U��5'���k!���8=�x?{?�0�>�Zk?�
C?�s�<2����tS���
� �t=iW?��h?�>fq��-�Ͼ�I����5?�ge?�N>.�i�,/��.��#��b?�n?�x?����H}� ��p���6?(��?Cr����hj3�]�(�l�>/��>�*?Mo��[�>��a?���������ſު0����?�m@�'@��� �b�/P�ޒ�>��?8����_޾��=1����_��<�?�B�������,N������l?bٕ?��?�H��l�����=���4��?���?�N� S�=t�1���L$Ӿ�"b�	b�=C^���P�����B������辨Qz��/;�>/�@����h?�蒾F3߿>���Ǌ�P�þ� ����>$ A>�-�&9��^䂿sjJ���4��rD�/��Iw�>�/>�������Ƀ{��2;��0�����>Ӱ�`a�>*(S�ծ���$��ſB<�6�>,��>vӆ>p���D��９?�j���\ο�����E���X?fR�?BL�?�7?og3<��w��9|�j�#�#�F?y=s?�Y?�C%��v\�_�7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�x�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�\�_?$�a�J�p���-���ƽ�ۡ>�0��e\��M�����Xe�
���@y����?L^�?g�?ص�� #�d6%?�>b����8Ǿ��<���>�(�>*N>�H_���u>����:�#i	>���?�~�?Pj?���������U>
�}?�}�>(Ä?�@�=�L�>X*�=�尾�� ���!>���=*.�d�?yN?�Y�>A6�=Z3�!�-��E��Q�{�[[B�_�>0a?g�K?<Vd>�%����K�+l!�%5ѽސ4�Rx�q:�u1���ݽ�k5>
Q=>��>��>�iӾ��+?A>,���ֿ�c��1D$��X?���> �?�i۾:���<�>HWR?(՞>��&��4����j��Q�?|��?�?B�Ѿ�������=��>�'�>�mw�ڢ����:�<DI?i�v��ۃ��H���G>z!�?��	@"��?1{�^�?�$�m���R��V��]A��=��N?�ƾ:�@>�
?�Zh=Y�c������v���>�?~�?n�>��a?.g�S/1���'>� �>j�E?���>T�7=dZѾ�nQ>�-?�(���������c?��@��@�X?�௿��ɿ����]�XV����>��8��o�=9��X�׺K=�✽��'��]A=`�{>X�#>�M�=<`3>>AK>�vg>XW����#��N���"|�y5���+�b������=|_�� ��g�:���.,��?(�R��:��/��0�@��=<"O?%�I?��W?���>n2&���G>���^=-�i���J=�	�>D@?��S?��,?��B=�Ǿ�oc�=�q�}#�������%�>�>`>'e�>��>�S�>ړ'>=�>��?>���>�-	="�e����<,��=YmR>It�>���>zy>N?<>;�>�δ�j1���h��w�C!̽� �?������J�2��:������a�=�`.?x>����>п���12H?���V(���+�?�>��0?9cW?ٟ>�����T��6>i���j��Y>20 �܀l�e�)��&Q>Al?F9V>��m>%+2��v7��N�����p>�a4?%ں��cC��yx��QI���ݾ�>>7�>� üՄ �g���t~��(b���=��:?:?νDG���2n�����2+N>Wa>��=��=�S>V��k4�B�J�
m=qp�=Oa>�i?��2>���=<��>����S��>��I>� 7>��B?c�&?�a�� �f�Gr�18��~>��>+�v>�R>�5H��и=���>��_>Yx�v���w���*F��C[>I�}��S�X�5�f��=Ǣ��޾�=H��=F����E���=�~?���(䈿��e���lD?S+?] �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l�6>�^%?��ӾA�>�V����������q��²��C�>C�t?	���0�=f����9�>���>�#�z����пUW���
?���?Ϥ?��c������长��?�e�?*�i?��s>�C��=þ7��>��g?�uh?J��>2T ���*��K&?S�?/�n?�7>]�r?^�?�9?P>�D:�����5)����>=�W>R���	������ubM����9�[��Q��.��D�>�]���>��ʽA�����=W�f�MHR�8�=�x�>o�>�
�=t͸>���>3T�>oն>��W�@j��O���_����K?��?���@�h��K�< y�=�Y��� ?/�6?en�;B�Ⱦ�>�7_?��?�]?i��>|/����K
���/���<�*7>F��>���>D?@�̀]>�ξ�pL����>��>CA$�>ݾz䅾�2�����>�� ?���>���=N� ?Η#?3�j>�J�>.oE�k7����E��y�>��>�O?��~?2�?D̹��W3�X	��⡿L�[��N>��x?PJ?Gƕ>�����|��aD��4H�����呂?�zg?y��*�?P5�?�~??�A?�If>���
ؾ&*���ڀ>GM"?����A�&�{g	��`?��?���>���|-�>ں�1�����"?5B\?%?�h��`�������<���?�q��A�;�A��>p�>X�����=�m>�"�=��n��
7�,<#<'��=���>��=l�4�8L���z1?�H��h��Kӽ����+F��<?H��>v#���g?������������(��NO����?^r�?˵�?��=,���g�?��?��!?��?�I��ڨ���2����2�����$�M�>���>�=�r<��?������Y+��yDY�Q�B�DP?���>|��>a��>�j>��?�پE� �����^G��3/�������&��?�3G;81���`g��L��$"2���(>l�a�p��>Cғ>1�S>%d�>�>y�ܽC�>�b>O�>H� ?�;k>�1>�m>� ��v��qLR?Z���O�'�Ű�%���
4B?�od?�-�>��h�߇��{����?��?�r�?�Cv>[}h��)+�
l?
8�>7��Yo
?():=h!�1e�<RQ��T���4��{3���>
M׽� :�$M�3uf��f
?�,?
��w�̾2&׽*�׾B�;�k?b?�.���?���b��i-���g�NVֽH�پ!T���
��Ȃ�`Y���D������.�/���<�'?cc?<�SВ�����^m��Y �h�p>;ԧ>�1�>��?�w�=M�־��$��aQ�����,"���?�A�?��>�B?d�2?/�K?MnD?��z>Y�>�A���?��\>��>W�?�L??�F?ҺD?m� ?� ?�	$>���~о�Iž5�?Jv3?�)?�S ?؅ ?X���ߛ��s��<�1�<#�u��@U�W��2<���EҺ=W��=`Y>$� ?�Y��ͼ4�?������>b+1?���>\��>����_A���֖=�I�>�< ?Il�>(־��g�!����>�m}?C0�~�=T�6>���=L�)�Α-<�gW=>[��$u<!9��}�VT7�u�=�>=�X��{�������8�<��7=��>)�?�ь>�^�>0N���� �:��ʹ�="X>�SU>m">�ھ*b��h����h�c�z>���?�ֳ?�w=z?�=���=�`��
���ʶ�����&��<
�?��!?�T?<��?�<?�,$?
>��/���T>���8��js?�,?k��>���$�ʾ��3��?�Y?�>a�����?)���¾_�Խ�>A`/��/~����D��v������z��A��?p��?�wA�L�6��t����]����C?�-�>�S�>��>��)���g��#�0;>���>~R?2��>�\X?�$s? �&?2�<�a����Sc~��<>vP�>��7?
�?I �?_��?��"?�#�>�'����� ��q3���H�h[����=��>��>n%�>�� >�`W=���m
�=��fР=�4>��>�M�>���>�>��h�BH?y$�>Db��=���y���ہ�w9=���t?@��?}�+?�_=�����D�@��B�>�?;��?�K)?��V���=g���c����o���> ˺>)�>Q�=��9=C>��>8K�>�d�%��R�8��U�x�?�dF?-��=Hsǿ*n�P�־�����=%�"�ξ;IR�@X��:�����r���9���p����Ⱦ����q� ��=�>Dc>�a�>�<%(��s&�)r�=\'t>�⑼O�=(�b��Nt��.>w\�e[�y�� �R�k�X恺�%Ⱦ�|?��G?�*?��B?u|u>��#>�R��>Aύ�=?�IS>�gN�ܷ��,<����6��2�ھӭվ�a�
F����>�F�L'>�+>�u�=&n�<���=�]a=Tx�=#Dc���=�g�=ۍ�=�õ=�=c�>�>�N�?����癞�.qk���`���7?�'�>5'�>�2��&6?��>���������(�u}?[�@Y��?JE?��"���e>"�h�<��=p�(>�Nƾ0��<��>�8a�T��>�9�>)�N�}\��^o̽y��?��@ڷ>?�S���пQN�>Ǘ�>���>A�{Q-���Ⱥ��m�Uþ2%?s>��,�nʒ>��>��ܾ:���y�>S�>GA�<~08��:@��)�=��d�mɰ��H�À{>�ڂ>D�<zD��}߻-�;=�K�=�W�=2̈́�8��>^��|���a�;�0\>`��>@�>��?#�=?Q�R?h�>�M�8�׾EP����r>|������>g�>�q�=�v�>J7?*~'?.�D?��>Pb=���>�F�>��E�,W�y��������Ž�.�?���?`͟><��<CpýzT�`4<�m��ã	??1?��>3?<>{'�$d迊5G�*����?�;�Z=�&~�2з�M��c���ၾLe�=i"�>�G�>���>i�A>�Fu>��>B@�>ط�=��=S�x=���;��>>A����Zb=+�e>=b��-�Y�=�=��=�=RW�=De=|�U������=�P�>5Q�=��>��=���>�>l� N�s�<�ȧ���;�\|`�]�|���3��l��<�/>fL�>e��d8���m?\q�=�> ��?[_z?Oٛ=�v�����> ��:�"�߅�;�Â=-o>�.��� a�ߺY�ɰK��?����>��>��>y�r>��,��1>���t=���E3����>pَ��������q��2���埿]i�)���H�D?�ه����=��|?f/H?���?Ď�>|���G�־�1>�X����<|�2�q����V�?�a%?��>l�쾲�E�֓׾e��7�>|�(�z�T�'���n7�9�=�6�CR�>�ٛ�/�����.�R������+\�����/2�>@�n?̈́�?�h��[�}�HC^�: ������?���?-��>6.(?�''?t'�=N
��KϽ���>0a<?t�?���?��>%��=�3��"J�>�
?#U�?�?�r?M=�2��>IV<wP+>S����
�=a`>�Ĩ=��=�;?�`	?�=	?�㢽IK�����n�_Z��I =!��=p�>��> �v>]1�=�Y=�Փ=�MU>�T�>#�>�g>�J�>�%�>2Y��Q��h�?��@���s>�L?�mE>v#�="��_A�0Ȃ�?�=�����E9��hS���r=	>	/>g��3��>+	ؿr�?�H�>j�2��H6?J��A��a?�>gN�>��9>���>��9>�=p,�>�3�>1��=R,{>8;�=�ھٳ	>��
� m ���@���N���Ծ%�z>�B���64���$��uL�/轾v!	�8 k������>��A/<J��?����b�k�%�gc�.�?jF�>�c4?�t��5L���>3"�>���>ߘ �؀�� ���߾�9�?4O�?�_>-ݝ>�\?\�!?��l�\3���X�ր�^7��X�/^�Mō����N��an�n\?>�r?F�;?!�n=�{y>��?k��n�K�u>�z6��;3�(�D=��>9����u��ġ޾�e��/3#�'�>~Vm?e6z?�C?��.�� C>�]�>w��>��1?��?�'?�$@?��޼^C#?���>Ҧ*?�j?�E.?�K@?�?���=ȷ>c�<��#><��$�$��64>��_��Ow<�H$�*�<s��=pD�=ņ�=�T	>i5t<��K�1��a�<�'Y=�'�=��,>���=}�>@�]?3D�>
>�7?�E��|8�������.?��8=�x��$�������m��m�>��j?*ҫ?�Z?�ed>M�A���B�2�>��>aU&>��[>�>���E�?d�=>� >�Y�=QYO���)�	�����H��<�x>���>R�{>c|��6&>g����n{��g>��O�%����|Q�D�G�0!2��ww�#��>RkK?�d?/}�=r��^�����f��K*?��;?CM?lx�?6�=�Xܾ0�:��K���!�Gf�>\��<�s�������X#<�":F��Br>�Ƞ�E�Ծ��C>���!|��XE�6�A�%�ݾh����[��o���{0��J���;�,�<y,�=���g�@�ŕ�4N���XC?�w�=q�����E��=D�>�R�>��'��Q>�SK����=�]>�Y>���Q����?��d��D�>�oE?Gh_?oo�?O����r�-�B����������ʼ��?�B�>�%?�B>�<�=%���o���d��G����>��>֬�(�G�q����8����$��r�>�	?��>��?��R?1�
?y`?��)?�%?)�>$����㸾pA&?+��?'�=��Խ��T���8��F���>ׁ)?S�B��>Ċ?5�?0�&?l�Q?��?��>ݬ �|C@����>�W�>�W��a����_>��J?}��>�=Y?wԃ?��=>��5��ꢾ�ة��]�=>��2?�5#?��?C��>�!�>���Rfe=g��>�Xc?�?��n?��=��?�*>n��>0c�=펚>�4�>d?��N?��r?=�J?�P�>(��<�����㳽\[��]`�u��;n�< �=¼��r�$����ϵ<��;�[�A>��u׼��6�\U�0jg<�]�>e�s>�Ε�&$1>�ľ<���l@>d���Q��E���lF:�>H�=�>�?5��>c1#���=宼>|)�>����J(?5�?�.?A+;s�b�n�ھ�L����>��A?�&�=��l�9���2�u��+f=��m?�m^?��W�p��6�b?�]?�g�=���þ�b�%���O?I�
?<�G�~�>��~?'�q?��>�e�:n�"��
Db��j��ж=`r�>"X�T�d��?�>}�7?�N�>��b>#�=�u۾��w�r��L?��?�?���?�**>|�n�>4�.���
}��]?A��>d|o�b)?��0��ƾ��P ���Ѿ*����R��ٛ��ku!�et�,n� Ì��?�����z?v��?�o?[Qs?������j�)#;�(���&�L�s.�������C�lI�<�[�,�p��d��	�=ݾ�s�z2l��?<�w��?)$?G�6�:�?Ϯ���۾F�����>�[���$0�;f�=~���=C�V=�f�r���ݱ���?j��>�P�>��G?�&Y�i�?��w(��s9���f6>�5�>4�h>�>��1���M�����<�;����ཉ�~>��m?ʺP?<�?�?9��-#�R6��`Q���I>O���ܖ<A��>�Y>�	j�	&_�2	/�s<��`r���PB��Xh�h�=?Wս>"��>_��?L��>'�U׾�����d.�*b��þ>fb?^�>�k>>p!�Ƌ����>�lu?k��>y�>:8���I.�zm��]�
?4�>���>~��>�!��O�.A������5���4=.#[?����փ���_>P?eq� P'=�o�>2�ڽ)��������^�C>W��>Q�=9>>�{Ծl����r������(?�)?_���U*��\>�1"?Q��>W�>�ك?���>��¾��2:��?֔^?,J?@A?I�>;R$=�����ǽL(���3=?M�>MY>�Jp=�N�=XP�r/Y��~��'J=�=*vȼ�ݴ���%<�����NK<Y��<ʻ4>�1ۿ�J��r׾5���-�6�	�2d���ж��x�����K|��|^���]v����7 '�!V��,e�B���n����?���?M=��ƒ���)���8���K���D�>ʉt�|y��מּ-C��-���|�xY���U"�D�P���i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >tC�<-����뾭����ο@�����^?���>��/��o��>ߥ�>�X>�Hq>����螾p1�<��?7�-?��>Ŏr�1�ɿc����¤<���?0�@�xA?n�(����^V=���>��	?,�?>�\1��E����<K�>Q=�?���?�FM=��W�m�	��|e?��<��F�q߻�&�==#�=
"=�����J>�[�>`��vA��~ܽ��4>"؅>�u"�Ҙ�Vi^����<~}]>4�ս�0��kۆ?��Y���d���,��#���m�=�Wu?Vi�>Z3�=s�J?��8�
tѿhf�n�F?���?���?Ȟ9?���i�>��⾂R?��??O�>B�%��cq�>�=�5��	ed=Aξ4�c�|u><��>��h>�,� d�?)��?s��H�=$n��*�����s��=��	��н[�Խ������*�&)���,��Ǚ˻)�>�>vug>�q>%$J>��9>RGO?Mt?S��>��L>���`-�xzϾ��ʽ�ۓ����Z����#�/B;A������@����4���'�S
ھ+!=���=x6R�1����� �;�b�U�F�F�.?�u$>��ʾ��M�ɣ-<"pʾ=���߄��⥽X.̾�1�M"n�J͟?��A?����c�V�d��7Y�ӂ���W?Q�T��묾\��=h�����=�$�>H��=���� 3��~S�ƺ-?ȿ?F�¾A����:>�T���R:=��(?��>>RX;�U�>D�'?�=7������V>�t6>^�>B��>��=�������]?A-O?i���%����>s����x�mW.=�!>�>:�+���*�h>,�#=�����G��wk�g�=[(W?���>��)����`��J���[==�x?��?�-�>{k?#�B?�Ԥ< h����S���dw=��W?{)i?��>�����	о����s�5?��e?"�N>Yah����y�.��T��$?��n?_?{���v}�=����ln6?�Ӄ?m)e��#�����=� ����>���>��$?֨-����>+g?�ֈ�I����ſ�1%����?�i@�<�?��¼��1���<��>��?����~���">���du��v&?20���I���tR��m��mHd?�ؘ?L�"?�������>��I�ޞ�?�g�?\����[����}�a��0ƾ�?�C+�=Q�ǽ�ͽ ݾ�12�c)��o��Ŵ��8x?��}>�@��ս7)�>�0��\�z�������r׾etؽ��?f�>�F �0{Ǿ_
u���d�l�?��_J��j�GM�>X�>z���������{��v;������>�{�x�>�S��)������q4<�ؒ>���>���>�6��ֽ��ƙ?�h���Aο׭�����ʼX?`i�?�r�?7x?��8<;�v�ex{�C���1G? �s?�Z?�%�d]��7�;�j?�_���U`�+�4�.HE��U>�"3?OC�>@�-���|=�>���>�g>�#/�k�Ŀoٶ�����g��?Չ�?�o꾻��>\��?�s+?�i�8���[��{�*��+��<A?�2>q�����!�w0=�1Ғ��
?�~0?�z��.�]�_?+�a�M�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�i	>���?�~�?Qj?���� ����U>	�}?��>��?���=���>ۋ�=�����C �!>�>�=68>��9?��M?A��>�s�=��9�� /��9F��;R�2"�"�C��ˇ>�a?oAL?�b>!���,�g� ��Ͻ�I2�x-�+�?�KF-���޽&�5>e�=>�>��D�r�Ҿ��??s!��ۿҬ��{���mx?I�>�'/?^����s��G�>�We?��!?;'��ᦿ�Z��j�c��v�?���?f�?��˾�4c�B�>8��>��g>-����w���t)����=�=#?�[�tW��n�w��ډ>0W�?��@��?b�d���?>������	������)�!�*�=&�;?����r>��?U�=eCq��㪿�t�ݢ�>�?���?GP�>~�h?*An��S>����=�p�>Z�`?�?�(:]&�a�K>@�?��.5����L�e?�H@4�@ćZ?�L��jϿȌ�������I��2�>T�= ��=�ƽC>�>м�l<�ڽn��=q�?���>Tsk>�PG>�)�=#pi>+�}��!�1��'D��e5�j� �-n�_��������k�������ž�+�=�S�D�]��E������;=�f�=Ed?�ta?�o?!Z?[�l;N�R>/�өT=<mq�J��'?�>�? H?�?��<Lʾwt����}�������ư>��>��>5��>��|>+:=Q#>B�>kՠ>��">���=�2=�Ys=��E>$Y�>�o�>���>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��s�T�4:>9����j�5`>�+ �~l���)��%Q>wl?)f>�u>�L3�-+8���P� ���G|>��5?���7�8���u�c�H�Hݾg�L>E��>��M�B������J���h��F|=XN:?�s?Y&��QҰ���u��J���Q>�S]>� =�=o0M>Z�d�'�ǽ�#H���-=�="_>�?f�+>3ِ=~��>����zJ�v�>��B>�S.>�>?]%?�B�5�������X�+�� w>t��>�H�>��>��H��=�l�>��c>��
������H�H}?�\&X>[]��N�^�\(}�T�{=f&�����=4��=��=��I%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>|U�蛘��̌�\`���e�;`��>j�f?Q��Z�<��<��?,�-?a��|����ſ�gd�ϧ�>�5�?�Y�?�"d� h���'x��?!?�5�?�+I?̔�>4��/ֲ�G��>��V?IEy?X��>(Ծ$P����?/��?�sc?��t>�?	w?�/?����2D�Q�������&m>��=_��>�j�=��ɾ�1�����f��IR�|��wD>a�<u��>�^�^q����=����)���-?�g�>ܳ�>	>��>�v�>k=�>v�P>k��>��㥾�/$�y�K?���?���2n��P�<���=��^��&?}I4?�m[�}�Ͼ�ը>Һ\?e?�[?�c�>>��M>��E迿0~����<o�K>4�>�H�>%���FK>��Ծ�4D�Mp�>З>�����?ھ�,���N��EB�>�e!?���>�Ү=F� ?Ԑ#?1�j>F�>QtE�Y@����E����>d�>5S?!�~?�?=��� a3�=���衿^�[��N>�y?�h?���>���������G��oH�:��,��?�g?����?4�?^�??t�A?�6f>�k�j�׾ڪ����>*�!?�����A�#&����Z?�L?���>ˍ���8׽��ڼ�|�G�����?�\?06&?�Z�X�`��þI%�<��-�:�[�K��;?�D�&�>��>����_��=	�>�z�=&�m�`;6��x<S�=R��>_��=�96�M���#7?�[�g����К=�	��D����>2�v>�{���b�?�pe��!x��(��G���jH����?���?�b�?�9|�q��Q?a��?W7!?��?�j���'�Ǵ����A���=�Q��>iM�>���=� ����_���y����]����gm?��>�x?:?��w>-��>�������J���@���J�2��Z�)�e�#��x��䲾7�n�-	�������H\��%�>kn
�^��>�?�dA>���>�>,�r��u�>\��=�Wl>��>��v>U�D>��=L�.�2OKR?������'�d�辷����4B?;pd?�1�>>i�)�������?e��?:s�??v>%~h�;,+�~n?�=�>G���q
?�b:=#���*�<�V��<���7������>xI׽� :�[M��of��i
?"/?����̾[<׽�P�����=<�?�5#?�t/�/�X���q�<I]� |����&>ٚ��-	����nou����!���2{���C�P0��"�2?Y>Z?zr
�[�ԾkȾ�ia� 7���x>�9">�~�>9� ?8@>~����9��"v��)���#�>cҞ?�g�>�I?h;?�4P?rL?���>9��>����.��>�u�;?2�>��>��8?�-?r�/?�J?�@+?�Sc>v"��_���HtؾF�?�"??l?_?���1�½1w��H�W�Dz��ր�ӄ�=��<Bֽ�t��V=�xT>S;?�s���8�Gu����k>XZ7?g��>Ƞ�>aU���I�����<���>�`
?4��>G����,r�$�fJ�>�b�?����=tL)>A��=���U�ຒJ�=��� ��=}K��H�;��<]��=ғ�=����b�9I� ;�u�;Q��<�t�>�?m��>z[�>�L���� �/���'�=�#Y>�S>*>PGپ/}��( ����g��Xy>q�?�r�?B�f=��='�=�v��yI�������~��<Б?�@#?�_T?9��?�=?Ea#?ϒ>0�I���[�������?a!,?��>�����ʾ��։3�Н?U[?�<a����;)��¾��Խ��>�[/�h/~����HD��������2��'��?保?�A�P�6��x�տ��\����C?�!�>�X�>��>V�)���g�r%��1;>��>uR?#$�>�
P?�4{?��[?��S>�8���Qܙ�b���k">c�??�?�ʎ?E�x?6��>��>�*��>�H���h�~��;ނ�YX=�Y>e��>�s�>��>���=�Ƚ���>��Z�=lib>�s�>�>%��>��v>�D�<��G?���> _��O���褾�ă�g=�x�u?��?�+?�I=���S�E��E���K�>�n�?N��?14*?��S����=d�ּq඾��q��#�>�۹>�/�>f̓=c�F=�b>�>`��>7&��^��o8��MM�8�?%F?�=UĿe�k�A�R�㋐��)�<���Ŀn�l���ok�I�{=A���������$T^�����Ǆ��;���Ӹ���$��O7 ?��=��=��=�զ9��G=�D=���:{�=�Q��!�v�X�C��������Gwv�'����.==zڼ�c���'�?�X;?/%?zsG?Pȍ>��y>�M� qx>�� �.�>G|�>���$�{�eU>����$`�������!��%d��1x�4��=�SٽE�9>}��= ��=$>�I*�1��Ib">G�o=�=�=ο5>�c*>���=W�=�2>��L=0ހ?�+��+�� aL��m��*?)��>�_>Q~Ӿ��a?�'�>�V��k@���#(���?�]�?P��?��?Jg���>��h�b�+=c�>��x����=g]�>&T��R�>�'�>�D3�}����A��DL�?�Z@�>=?����o�¿�W�>c4>�5H>OTP�v7�q���tJ����1m?f�<��}־-J>�/>-��1����Y=��H>�ڪ=vȽ>0W�jDB=g𶽈�<�C)=�J�>�v2>��= ��:09�=���;��=�L	>O߼�!"=�2�=f��=,{�=}�>�d>b��>,�?�[0?�Ud?�9�>�n��Ͼ8��oD�>���=?�>J�=^B>M��>$�7?�D?m�K?T��>Ϯ�=��>�	�>��,�/�m�:j徜ɧ��N�<~��?�͆?�ϸ>0ZR<��A�$��`>�ŽZu?�P1?�j?)�>�)���ٿ{H��kA�L�>�H_�����P����4X=2C���!=�;J=m;�>�U(?>K�>!�>С�>A>�x�>�`�>}�>�.�=���<;������I��;��=�)l���b��U#:,��=��J>F&x��j�I�=�u?=
7>�����>=�>�C�=�X�>��=o��6�=�2���(���,>������@e�@q��1)���ݽ��h>��n>�5��c���?sE>�>�G�?0�l?�c�=�c���̾AJ��uo�b����f>3�>\��?�W���W�1P����%��>F�>��>��l>j,��"?�,�w=��`5���>e~��ܪ�+�-9q��?������9i�idԺ��D?)F�� ��=�!~?ίI?q�?���>?����ؾ�40>4J��w�=��I+q�kc���?+'?g��>��:�D�������z��>9��Y�i�����l�,�ƞ0�o����>����}�pi�3���^����Y���X4�>�Ie?�?�O�����e�o�2��Y���Y"?�I�?�(�>��>�3?��H=�>�����[��=@0\?K��?�u�?p��>iG�=K2����>��?���?ָ�?b�k?{a�~��>H�	�Cn�=�n����Z=�t>� �=�-
>ś?;�?� ?�����qݾ	'����^�"�q=�2=�M�>Fߤ>ɗl>K�#>���<t��=��>�2�>�2�>�l>W��>ܡ�>Џ�'��!�?�^~=S�>�K?`�>��>ُ�<4zh�D��=�*۽��.�>�==�N�=��=y)�=�~>�=����>�3¿�Z�?w�J>9��M2?u���#;���>~�$>jѷ=�bb>���>�Ħ>�>'�k>�ib=SkF>61>*hӾq�>���� ��0C���R�KҾ��w>�����+#�?4	�����)H��#��e���?j��T���=��ɮ<�3�? ���k�ɝ)�������?`H�>��5?����Մ��>�~�> �>����u���`����v���? �?�Cc>1"�>U�W?p�?�1��3�otZ���u�zA��e��`����.���.�
����]�_?^�x?sA?S��<R4z>(��?��%��2$�>�)/�� ;��|;=��>�����`�E�ӾW�þhX��F>Ío?��?�M?�CV�8/k��)>�:?��1?	>t?Կ1?s\;?.��x$?� 1>��?қ?��4?5�.?^�
?�0>@S�=L��y�=�e��Ԋ�ׇѽ˽�qI2=j\x=�AY:n�	<h=���<��tWм��[;�%�����<��:=�֣=��=���>�]?���>�w�>��7?�_�-�7�������.?�6=�΂��:��E����>�j?U��?Z?�	b>�`B��C��T>cr�>&'>DI\>GX�>�@�C�E��=�`>�>KL�=y;F�Fʀ�yw	������<!f>���>��|>{����()>8����y�@b>�wR��S��1kQ���G��S1�8Jx��[�>wPK?P�?���=��B���COf�K�)?S�;?VM?W+�?�B�=�Xܾӏ:�q=J�/�����>xh�<�|�3Z��k���r;���?�Yp>�A��۠��hb>}���^޾�n�v
J���`�L=�|��:V=��?�վ�8���=
>���� �����ժ��-J?k=�p���\U��t��ۿ>ߵ�>�Ю>�:���v�-�@�����T�=��>��:><������+tG�L2���>�<P?�"L?C!�?��R�(�V�[V�����Q.����V{?��>c��>��{>4��==�����ik�1�X��@�>��>�h��h*�?H۾�G�MV쾞�>>��>�3I=p�?G?�k'?B d?_=	?���>5

>��=�ϧ�M|&?ī�?�/�=3����AK���;��F?�p��>��*?]�F�!'�>��?�!?�*?;P?�?<�=�� ��D�C�>��>�yS������YW>ypB?*�>S�V?�׃?��J>��3�񤣾Ȱ�����=��*>{�2?a�$?�2?Wp�>pl�>����r�u=.��>��b?p��?��n?�<�='W? �,>�}�>Dɐ=��>~��>�%?��N?��s?�}J?F1�>rǂ<" �������u��zY�F�;�<޼o=t��[,v�� ��3�<�-�;�L��hj���@�埔��C<�L�>H�t>='��qV2>�þ8?��@>�����\���_���C<��R�=��>0�?��>�+#�VI�=���>N7�>\����'?��?�?С:w,b�M۾q�L���>A�A?�s�=�l��9��Xu��h=ܓm?;K^?��W�������b?��]?ie�1=�J�þϺb�F�龓�O?��
?+�G���>`�~?��q?¹�>��e�=9n����Cb�:�j��Ӷ=�r�>�W���d��;�>��7?DS�>]�b>�(�=]t۾k�w�pq���?��?u�?G��?)*>4�n��2�T�5ň���V?��>�d����?�����1D��S���VA;b��Ol���S��ք�9$.�ǒƾ�-r���d=|�?�Ԗ?F�{?�D?O�˾��o�&UZ������X��Q�������N���U�lfH�P�n� .����%پf���f�2�2�{³?�,?� ߽F��>/���b�*��=i->)7���� ����=&1P��<k=�;�<L�f��h'��a���;?���>��>�x0?ߝ`��)3���*�n�;���M�J>�Ҵ>t�>���> K꼇�w�4���f�ʾ�셾��ֽ�%n>Vf?(Gm?4�?�v��� ����?V���<Sr��^}����E>'l>��l1��X ,�؉3�;c�pc���� �׾�p�<��
?�p�>1x�>B�?�+?�'����-Ⱦ��+�#=�|�>	{?¹�>e�q>;�t�ƿ.����>B(g?�\?I��>�h����������f�&��>�n�>��>��q>��f��N�@���������2�fo�=U�I?\����Nr�/�>�m^?�I=:�U�1��>��#�5��6��`8x��o>e�?�>:Њ>��ɾ,��Q3f��s�J)?�+?���JM(�<�>��?`��>U�>��?���>�ľ���4?��^?D3J?.8@?�D�>�v=����x�̽�[)�6/=�E�>��\>�t=��=.��jzV�Q�T�E=�_�=Ք�;캽I�"<�T��rA�<���<\V:>m1ۿ,�J�?�׾�o��]
�xƈ��� )����	��"�������w�����_&�~�V���f�����m����?#��?�c��<*���Ȁ��0��
˺>{�r�8�s��������û�����$����!���O�li�5#f�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >bC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾r1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@wjA?��(��쾗�W=��>(v	?��?>T1�,t�V�� ��>j.�?hۊ?�L=�W�a!
�/he?|�<��F�Q��}��=��=��=J��ziJ>��>����A���ݽ�&4>�x�>_�!��Z���]����<��]>\�ս>����ۄ?�h\��f�}�/��]��g�>�U?��>���=1�,?��G�H�Ͽ��\���`?2�?���?�')?-
��>zݾ��M?�^6?�i�>|�&��t����=��§�I��R\V�p��=���>p�>Cn+����DP�"��i��=������Ŀ���ml�qD�<ˣY=�7�]���r����)љ�-H��-����=@H>% i>ߕa>y,>��v>4�L?i�h?��>o�5>��ν�N��KԾ�}!�����F��P��;s+��ę�����پ���1�!������¾!=�!�=7R�^���"� �Z�b�T�F���.?w$>T�ʾ��M�I�-<�pʾK����ڄ�᥽�-̾�1�&"n�f͟?��A?������V�U��.X�����@�W?tP�޻�}ꬾ��=������=�$�>���=���� 3�w~S��(?qi?`,Ѿ�	O���~>����}�u=�N?u�>q5���q>KO%?��V�����&�a>��>N�>F�>%��=�O���;�d?C~R?~�˽�Ԓ��R>��ؾL���r����"`=|�p�u�T�>���=D߆�՘�;r������=�%W?���>�)�����O��V��+{==�x?I�?C*�>�rk?��B?A�<�h����S���(}w=��W?$i?b�>_����о}t����5?Ϟe?m�N>!uh���龇�.��U��?��n?@g?ਜ��s}�I�����o6?��?(�P��5��'�3���J�K��>A��>��?��ؾ"�]>?!z?t�̾���#˿-�8�)�?7�@�,�?4߽~���ܽO3�>a�'?����]������=�U�� �A�?�`���m���sP��"���gp?�Ǒ?��?�S�������= ֓�V�?���?�(��@X<� �9k�s� ��ތ<��=��"��� ���t6�_Ⱦ���pk��]����>BE@^�Խq�>�M:�05´	ο�~���jϾX�f�r�?�/�>+-׽�I��|l�u@u�G��I�D����I�>D�>����|�����{� z;������>�#���>g�S�& ��ȋ����3<֒>��>l��>},���۽��ə?h���Cο��������X?�i�?�r�?Cn?ފ8<W�v�	f{�h�M+G?��s?�Z?u%�s]��7�,�j?�_���U`��4�cHE��U>�"3?�B�>,�-���|=i>���>^g>�#/�{�Ŀ}ٶ����b��?܉�?�o����>k��?qs+?�i�8���[����*�n�+��<A?�2>@���r�!�\0=�,Ғ��
?�~0?�z��.�X�_?�a�M�p���-�B�ƽ�ۡ>��0�f\��O��4���Xe�	���@y����?I^�?c�?���� #�d6%?�>^����8Ǿ�<���>�(�>�)N>�H_���u>����:��h	>���?�~�?Qj?���������U>�}?7��>.m�?�f>f2�>"�=-]��Y����	>��=��@� ?9�L?���>�S�=��;��0�lE��O����]D�Z�>��`?�0L?�f>�z���"&�E.#��н��5�J}/���4����]�����>>��;>�m>j�J�Z�Ҿ��3?�����ֿr}��6� �+w�?�Y>k�?�ꕾ?>ؾ�ȍ>�Q`? ?�/��e����~�S�M�l�?B\�?�q?r]���<'L<�j�>V�>������H����>��<?�2������D��䧇>���?��	@ר�?$$����?f��6���凿�;����z��j�=T�:?��ž�w8>�1?l�=�Fh�3���E�|�ȿ>m�?�D�?V��>s_?�~o��33�@�=�g�>{M?K�?NW�<5�O}V>�r?rD�h+��R��1f?B�
@��@oRT?:̦���ֿ���C������LM�=�ؗ=PY1>��۽x��=a�3=9�?��8��?��=��>~f>�Vq>>�O>��;>/�*>���۵!� D��ot����C�W���\�o6[�)��g9v��o���I����)����½pY���P�	^&�I}]���->��c?�NL?d?v"?���DM)=�yھߘQ>	,�F�Ž�}<>X�?̷D?}t2?7:���@���`�rl��T]��M瑾ҋ&>�r��VR�>�(�>�<�>ZQ>7��>O��>���>�X�=����l5�����<�e>���>�1�>���>�C<>��>Fϴ��1��k�h��
w�p̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?��f>�(u>!�3�QK8�ٮP�Vw��#C|>�#6?����j9���u���H�`aݾUQM>�Ҿ>�bD�)[���1 �~zi��g{=�v:?Ƃ?�A���ڰ� �u��C��=R>�\>A)=	 �=�eM>�ob���ƽ%
H�jK.=���=��^>o�?�m1>+��=�>D����O�R~�>/8>�>�%<?uJ ?��g���I���"(�L&r>���>ꈀ>;>��K�롪=ǉ�>�ea>d���u�����i�E�pY>烅��>b�3牽�ew=���}�=ک�=�����<��?J=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿِ�>;�̽�����Љ�=x��;��o&?9p?���Db����*?g�H?���޼����ο�|��ee�>A�?��?�������?����>az�?�o<?�}E>�e���7��9X�>��E?�6X?Q"�>��6����>SX�?ᴉ?�k^>y�?�K}?^��>�3�����oA��Sċ��,�1��=7�>��==뱾ڣ6�����j��4[W����eT$>�]<1��>%7���TǾ�c�p9�D��C���+�>�>/�T>
��>�>�Q�>��>�=�<�6��')t������K?:�?�I�q�j��y�<Ḋ=�U�{%?��5?�kG���ξ���>��]?��?��Z?�B�>����L������`����n<h�F>��>�#�>a����V>�Ѿ�7�3�>���>n��>Eھ]i��p.˺��>�(#?�>e>�=� ?��#?g�j>�#�>dE��<����E����>W��>QO?m�~?��?�Ĺ��]3�D	��j硿��[�4N>'�x?c?���>����b���@1F�m�H�l���P��?6pg?�m�B?�3�?��??w�A?�-f>2��mؾ�5�����>�!?m����A���!��z�tE?��?c*�>�������$~$�����;����?U�[?u�$?{Y�
�]��达7o�<���J ���5<�ϖ�NL>W*>�}�����=<7>��=�Cz�k�1�ߤ�<��=��>՜�=R6���Y�,�>?� �P6��'�=�ɘ��$7��x?lb�>c6�B��?Q�Ľ���@	�������=���?9��?��?r�=zӌ��Fc?X߄?$�+?��>�dʾ���l����q�J
ٽSN�SU�>�X�>LE�=u+��葨�����֜�����kX��� ?i��>�%?��	?K1>!�z>+A����5��
�A��s�T�`���K��{����@S�̲��tj<l����셾4�>yx�I}�>$\�>�!�=Y�_>�(�>6=<���>��>T܂>�P�>6WB>�=�=��={s��Hi½�IR?���޿'����ȧ��./B?|nd?`)�>]�i���������}?を?Cq�?=Dv>�zh��'+�ym?;�>Q���n
?V:=ǹ����<LS�����hP�������>jc׽~#:�M�EMf�ok
?�-?�Ѝ��̾Z׽��Ⱦa��=*!�?�?�2�;�e�~<f��EZ�}�R�G��<q���H¾���1]�%��f���K����K�v��\9?w��?�P��4޾sԾF^g���(�8H�>u�>mY�>���>w�">O���L�<o��{*���@����>��j?#��>
�G?�$)?
QM?�?R?FUZ>B�>N������>Ψ��dU<>Q��>~�)?0�,?6&6?��?8!?�L>� �����O��7�?
Z?n�?���>I��>��6�c,��t�8=�'�= Y��Q&�ܭ�<E��<J������� =O�J>��?�g
��8����p>�5?���>?(�>7�������1<`z�>��?Oǐ>�^����o������>X(�?���]5�<�.>�5�=����:�:��=H���'��=>F��~�R��z�4/�={��=-A�9�q�Ȧ;:�5;���<�t�>��?���>�D�>]A��٨ �x���T�=Y>!S><>Fپp}���#����g�DWy>ev�?ky�?��f=7�=N��={��[S�����)������<�?�K#?ZWT?>��?�=?�g#?$�>v*��L��^��v��٭?u!,?
��>�����ʾ��Ӊ3�Н?f[?�<a����;)��¾��Խױ>�[/�f/~����9D�����G��4��?꿝?pA�S�6��x�ؿ���[��x�C?"�>Y�>��>R�)�~�g�r%��1;>���>eR?5�>o�Q?�x?��[?��T>��8��r���藿$cݻ�V>m=?���?ڍ�?.�x?#r�>�>x_8���ᾴ(�B��G���,%=��I>��>�[�>�T�>���=�rĽje����?� ��={�o>U��>�m�>x>�>,�>U��<��G?���>�]�����Y뤾ƃ�.=�˜u?���?��+?3R=�����E�QF���J�>)o�?���?�3*?߻S�i��=��ּMⶾ%�q��%�>۹>"2�>�Ɠ=~F=�c>s�>M��>*�a�Nq8�INM���?~F?:��=��ſ"r���q�"v��*�Q<WP��d�a�/��XqZ����=�?��q������^HW��垾I����~���^����x��M�>��=ː�=�.�=���<�8��r}�<�K=�d[<��=�,r�}�a<H2��Z�+>����{�?�(<:�F=U���د�Z{?�N?��)?a5=?L0|>�Mi=���.�>��:Vs?|�">;�νꭴ�1�@�{����P�����b��R�q���Լ=�����=��>;SY=�T�<�{4>U��=��>G�;=�կ;���=� e=��R=x@�=B;>�>��{?T�~��Ϝ�B�P���0T:?,ܬ>^ >�^���M@?�4�>풎�t���Z{��{?�&�?�y�?��?�q��C�>:8��隸�V�>W�&��4�=��1>���>g��>F�"�Nu���)�����?�@�:?�܊�{�ɿ��_>\E;>�U>��R� �(��D@��=a�CO��C?/A�L�Ͼq�n>ʕ�=T�z����NX=E�1>Q��=_��Y����=��z��$=a��=�>�E=>#��=ٽ�l�=ܡ<搳=�P->�R�:�\k:� ���F7=�Q�=:\>6%C>�a�>W+?F�0?:Ud?���>ڑm�g�Ͼ�d����>V��=�g�>��=��B>�a�>�}7?��C?/K?V��>�h�= 8�>�6�>,,�ޜm�P�զ��u�<��?���?��>Rjx<"�@�9���w>�X�˽�$?5�0?��?E��>����ݿ�+��%��d����=��>r�x���G��P1�u�w�u>�E�=o�3?,'?P��>��h>��-����>Ia�>Tzv=��m<���=̸����=��=�`H>�K�������E�����=�
��~н{b�<Y���>�ܽ���C>���>��=@x�>q��=f����h>U���4�WVe>�_��|J���a�~��'�(X���go>��w>�F)�RI���s�>H�y=/�p>���?��g?�<=����H���4��݆l��3=�W�=
0V>�J�E�V�ɊX���@��=��y��>���>V�><Vm>c�+��?��u=*j�A.5�-0�>
{��m��C�C#q��2�� ���4i�/b�"�D?yE����=�~?4�I?���?�u�>Rʘ���ؾF�/>~m����=���@�p�����!?�'?|�>h$�-�D���˾�x�����>�NA��/Q��	���m/�ǼS�M���ր�>�,���о�k+�����/{���CF�n�����>.K?=��?�&f�r���S�N�RS�8����	?m�q?�Š>��?�c?�'9���Ӿ�_�����=Cwe?g��?�?�V5>�4�=�"�����>Nm	?ݞ�?�<�?��r?,�@���>�o�:/g>���
��=ט>��=���=˂?�[
?ɨ
?������	�ȴﾱ�d-^����<W��=f,�>S^�>�gp>!��=�[=1�=B�^>�'�>c��>�>e>�a�>f�>yꤾ&Z���%?; �=[]�>H�1?ڀ>?�L=/S��+�<s�^���@��,�䳽�!ٽ�Ҹ<>�ں�S=�u��{�>4)ǿ�3�?�T>�Z��E?k����i$��Q>��T>�Qؽi��>��F>��|>���>eW�>j�>�C�>v%>җɾ@T0>�-Ӿ���5�J��ep��ž�ڐ>�ٛ��d�V��C>�q��C>پ>��W�t��H����5��b=RC�?]�+�R���VG6�Eb6�l?��>v=\?�i��v��0�>Qf?�`�>CU�)���҇���̾���?��?ʤc>�u�>H�V?f�?}�.��D3���Y��pu���A�I e�a����� s����	�-���5)_?��x?A?n�<çx>2C�?*%�9%����>ˇ.��;��1=�E�>e�����b���Ծ��¾���LG>S�n?�?�?��Q��d��G�d>��/?�,?�w?�.?�WD?q�� �8?@mp>�C ?�/	?\2?^�0?΁?��8>�J>�ŕ�Us�=큾�R����ݽ$7�[U�;3Bq=�,�=����<2�=�P=����6��A
��)_���=�S�=���=h�>Gl�>~�Y?+��>�M�>9?����/4��·���?>ru�*���=����M���پ� >��^?.��?dWS?aMs>�rI�":H�"�C>ہ>_� >s�W>$�> a콱�2�|ǈ=j> �=�g�=9.�41t����꾏�H�`<A�>qU�>��>�d�J�:>�����w��D>� N�5ƾ�R\�V�H�.�1��cn�w�>�L?��?N��=�p⾷��Gec��3$?�t@?j�I?��z?�Ɗ=vO�w;3��AH����Ӫ>��<!d��埿�H��a:���Жg>�w��G�����'>�@���L��1�G��]�z�1��p�,�:<=�u%���S�AI�	��=i�>�C־�.�h���ޱ���U?n�6<N�;΂b�1[���b!>�VU>��@>��<��ϼOj6��㑾��˼�1�>�%>��e}㾪+��|�r҄>>�U?�[?b��?H#��<\��9�!���������t�q���+?|��>��?�̴>�^>_E��cJ���T��rU��K�>y��>���t�K���z�߾h�:��χ>��"?F���"�?��y?�F�>�u8?�y3?��>2c>�q�����3.?�.�?���=Y����I��0�C��t���
?�o?�d��m?�?�+?\B#?ӑo?1�?�� >��ھ<�P�>ʭ>0��>�"Z�zɿ��=�Kh?��=�6n?�8�?���>��	�q��U������&OG>�8@?��9?=A.?C��>&��>;W�����=9(�>�vb?�!�?�[q?���=M�?�K3>,,�>+J�=_�>^u�>�`?U�N?�s?��I?r��>��<;���I��|iy�0�k��Wf;L`D<.pZ=����i���� ��<�L�;����ׯ���	�CtO�ȝ�E�;��>Pt>�啾d�1>Ϥľ�&��Tw@>mʘ�iƛ�"S��A�:��4�=�"�>�3?��>d�"��W�=yּ>�^�>���(?x?8=?6K�;ob���پ��M��L�>�1B?���=��l�G{��Lxu�Dbf=[�m?Q�^?��W�	���G�b?�]?h��=��þ:�b����F�O?'�
?�G���>~�~?Z�q?3��>2�e�.:n�*��Db���j�Ѷ=7r�>HX�(�d��?�>\�7?�N�>L�b>�%�=]u۾�w��q��s?��?�?���?6+*>��n�W4�x־������O?M��>������,?�!>:ι$�DC���^о�A����ξ��;�{��\�K���c���ʽ|$��A?�}?���?jFC?^�þ�/l�.{l��n���c���V�:��f9� ��cb��L��5"���?,۾�=N�[��*73�)�?��'?�`8�ʇ�>>��3�i�� >��Ӿ{l�f>ۂ���;��;�߈��.��2dؾ��$??|�>�x�>��4?os0��,I�q�M��iL����r�>U�>1��>���>�QE=��ٽ����8��žj��)�>6h?�eD?�d?{Y�M���pw��.-��FE���{��h�=�~Ƚ���>��5�[��S+���C�2������e������v�;"�S?��>�C%>�[|?�4?#�u��0��t�M���nM>��?�~?�?���>�z���5��M�>P�q?H��>��> ��Q���r�� !�Tn�>b�>�c�>%p7>
�4�9�[�o��ȝ����C�{ñ=�l?��}�1�]�hx>~,S?�)&;���<n��>v{z�o/���ྦྷ����=7�
?�j�=�S>����m���3���图|h4?��?�9������W>k�%?R�>�#?}T�?��=A&���>��$?!ST?�N?�;6?���>SW�=�_�:��\]v�s�=j�>G'c>N=�.�=6�}쎾��P�������=��<��n��'�=ַ]�y��IA��IX>l(ۿjbK��`׾�X�Ћ��	��z��y¯�����ݡ��L�����bw�6	���)��+V���b�ӌ�P�l����?��?et��~Ȇ�ս���b���� �9һ>�9v����L��s������ᾄ,��5!���O��4i�اe�M(?�����5ȿ١��ھ�7!?�L ?��y?5��$��7�&�#>:�<�^���N�)�ο������`?���>݂�:���{��>�%�>�X^>_bq>2C���g��W�<�?-?Q��>�Nn�T�ȿ�����Y�<���?!�@
}A?�(�����V=��>W�	?��?>oS1�>I������T�>X<�?���?P{M=?�W���	��e?ڄ<��F�.�ݻJ�=Z=�=�F=���g�J>mU�>T���SA�q@ܽB�4>څ>,~"�۫���^�x|�<��]>?�ս#;��$ք?ny\��f�Ԧ/�.Z���\>��T?--�>,;�=�,?11H�H�Ͽ�\�a?�+�?��?��(?먿�Oǚ>�ܾO�M?GR6?��>�o&���t�k��=���qr����i7V����=@��>Վ>܊,����O�Z����=~���3�¿̵�r�� �I�E��B����-��꽽�B�<����o�>�"@Ľ�3=D��=J�3>�;y>��6>E?E>J�V?�r?��>��p><n��[j��$�12;�y��B�P���Ҿn�3�G����. ����_ �:8�g������ =���=�6R�N���>� ���b���F���.?�v$>T�ʾ��M�_�-<vpʾ}���|ᄼl㥽T.̾*�1��!n�m͟?��A?����V�E��EU�^�����W?O����鬾��=���:�=�$�>b��=���` 3��}S��1:?�g ?]뽾�LT�J��=^����_��bN?�?�<��ʃ>�:?�l�<�^�9���>;3>>��>��>ۮ3>e¾ڲ#��d!?L�a?����?��>���������>�e�=�xV���{����>^X�=�f���&=�39���#=p`\?$G�>v�(�������w�<����u�?��0?ylE>_�m?��J?`�>�[̾q���Ҿz�>��Z?A@K?�>t�������6���.?3n]?��>�G���U�P�$�>�1?Ȣl?~�?h˻���x��}���h�B%B?pK�?��^�ɯ��£��톾ʉ�>\�>'��>h�)�`��>�;B?�*���䧿lv���o�Z/�?H�@S�@N�M�V����>-�$?Uh�>*2����ޗ��^����g=�h?#־�Ԑ���Q�>Q9���S?��?�?�ǎ�<F*�4=>�g���s�?��?�X���1�<�
��n��G��XEν��;ڽtŽ���G�@���ܾa/�ė���z����s>��@�㰽��>�h �֣߿�3Կ��t��Y����w�f�>���>�9��2྾h;x�]�k�WWN�WCI���`�SM�>��>���������{�1t;�󧟼��>���>��S�i#��m���:�4<�ޒ>���>D��>�3���ཾ�ř?�\���Bο��������X?Ij�?r�?�q?�8<��v�2�{��!��,G?	�s?�Z?�~%�5$]��W7�%�j?�_��wU`���4�sHE��U>�"3?�B�>T�-�b�|=�>���>g>�#/�y�Ŀ�ٶ�@���Y��?��?�o���>q��?ts+?�i�8���[����*���+��<A?�2>���J�!�D0=�OҒ�ļ
?X~0?{�i.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?J#�>��?W��=xm�>+��=�����B-��l#>�&�=�>�
�?P�M?�O�>w�=��8��/�pXF�\FR�;&�C�C�u�>��a?�L?�Lb>T��p�1�!!�/�ͽUX1�v��UD@�*�,���߽�45>��=>3>��D�M	Ӿ��;?Ve)� #�����}1=��d?���>\�?<Ͼ,a���ݨ���_?'��>�����������vj�?^;@��?T���A�<N>���>�eD>��N�Oz��ޡ>�0??Dn���l�������>*�?��@���?�>��Qc?K
������F~�2�4�۽׺>QB6?*�羪W>��?��=��z�	���m��!�>42�?^��?��>�wa?m�c�Rp2���=�2i>�vW?a�?-Yw��N�8xL>'�?*#�Di������Ds?v�@U@�^?e|����ֿ9ʘ�wľ5��	'=5U��U\*>�Ͻ�M��3S>S�=�]ѼS�>9n�>
od>i>͒C>_�V>ۖW>p���;���ǟ��6���2�9���:��q��T7���#���_�����>�R�������!@��)������� >{ W?|�N?��?4X?�	"���=&�Ͼ�%�=͋����=y�>g;?yS?��?�Z�=�����\�,��M���]11�,��>5/�>���>~0�=?Q�>���=�2�<�m>�c�>m��>�V����=�)7>#ِ>��>G?mV�>�C<>��>Fϴ��1��k�h��
w�r̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)���+���>}�0?�cW? �>!��x�T�5:>9����j�5`>�+ �~l���)��%Q>wl?�f>�u>̛3�qe8�k�P�t|��j|>�36?w鶾CD9���u���H�}cݾ4HM>�ľ>D�l�}�����vi��{=Yx:?݄?�6���ⰾc�u��C���PR>:\>8U=:i�=�XM>�ac���ƽOH�hg.==��=�^>\J?E�*>9��= 
�>���.lN�.�>�A>�->*�??�7%?���=������� �-���v>w>�>�>O�>��I�1��=���>wa>�)��؄���� �@��@W>����`��x�7rw=K욽���=���=:��i=�w�#=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ	�>^wШ�N[����S�}�>��>��h?����p̾P)��?QA�>�Ѻ�P��)�ο���b��>ֲ�?h��?P�y�I����2�-�?��?�At?�>ڽ���D~�� �>�GC?�2_?'�?!���$� A?�:�?Y�?��r>Vٕ?Ϳl?A=��d��j��Q�������3���f�=>��=݌��˜�"�W�������������?���<@��>/��=���L!��q= `j�i��Ks>�z�>Qv>)5>�&?~\�>_^�>�M1��v��/e������K?ٱ�?���� n���<���=K�^�9+?�K4?k]�4�ϾMԨ>p�\?���?[?a�>���:���⿿�����J�<C�K>9E�>|N�>�w���WK>��Ծ�DD�4y�>;җ>6����<ھ���:��jJ�>e!?'��>J��=� ?X�#?E\j>��>�dE�
;��Y�E����>E��>�(?ѣ~?��?�۹�6Y3�u���顿�[��N>��x?[l?ȕ>����������D���F�
����?'qg?�j潉(?�'�?ׅ??��A?��e>|����׾���6�>1�!?��ֺA��L&�� ��?�P?-��><��|�սQFּ����~����?((\?5A&?#��k+a���¾�3�<��"�E�U�G�;.hD�4�>؏>a���є�=@>�ְ=?Om�F6�q5g<s�=��>��=�)7��q���<?ՙ������h4ּ����.2��w�>e)*>d���hi?>�ؾ}m��Y�̿���D�#�?\v�?�e�?��ܽ�v���L?�L�?'?�>�>~@���<��{d�|��]��߶C����>� �>B�.�~$���W"��⫤��9��W�Jo�>�>x�?�`$?���>]$�>�����A���I��$�_����n�D�@S$��g�%m����g�?�̽ �þ��O��ˑ>�6<4�>��?�~>x��>���>ߠ�<T �>��=QK�>���>�n�>C�n>�yC>�i�=�ጽ�OR?����'�ٚ������-B?Wd?�d�>��g�8������m�?���?�p�?k�v>kh�!+��l?e@�>-'��&]
?�;=	�	�R��<a��I��G臽��
��>%T׽�:��M�~f�r
?�(?����u̾�׽�{��o/=g)~?��?�'�HT�B����U`���S�罶��(�z���Ig��1��?����̓���=��K𽫹?c��?2�����5�����N�/k��b�>\�>nG�>ĩ>��;����o*��k����z~���m�>Q�?}��>۝D?�n2?��i?�k?x��>��>�*����>�sL�6�^>D�'?��E?�hP?_D?�$?��I?z�?>��=�3�F⯾6.?t�	?[:.?<��>�?������ռc�u>���=�7J�����^�<s/�����:8�g;��N�'1>�Y?�{���8������j>x�7?�w�>3��>���5��r��<��>�
?�B�>�  ��|r��b��Q�>���?����`=��)>m
�=t���-4Ѻ'V�=���� ͐=�s���;�r�<���=��=��q�[�����:���;��<�t�>7�?���>�C�>�@��-� �c���e�=�Y>/S>X>Fپ�}���$��}�g��]y>�w�?�z�?��f=��=@��=}���U�����>���s��<�?9J#?.XT?^��?r�=?Wj#?�>
+�gM���^�����Į?w!,?
��>�����ʾ��Չ3�ڝ?h[?�<a����;)�ߐ¾��Խб>�[/�i/~����=D�?텻���U��5��?�?JA�V�6��x�ۿ���[��{�C?"�>Y�>��>T�)�}�g�r%��1;>���>kR?��>Q�O?w6{?9�[?hVU>Ҷ8���������*5�'�">x@?���?�?�y?Tn�>*�>��)��0�?���O���ɣ���Z=��Y>���>U�>���>���=�"Ƚ���	�=�H�=��b>b��>8��>i��>�w>{.�<{K?��?ľ�8�L���R�e���M�/`�?�I�?{68?�i]>x{�8� ��QӾ�C ?�,�?�o�?6�2?���m�=� ?�F�ž�d���>���>���> �>||���Q�<�Ԉ>���>�0�����,Z2�8�����
?lCG?�W->��ſYhq���k�▾�9<����T�j�KҜ���\�٨=Jҙ��g��㧾�TZ��𞾙���$W��{Ҟ��*��_��>���=�P�=�3�=c��<˟��-�<N�B=Ѓ�<�&=y����}d<�>��[�����O�̻�B<;�H=(�����˾1�}?�1I?��+?��C?�y>�R>#�3����>}̂�i<?H�U>M�P�掼��{;�������Ӱؾ�x׾�c��П��G>�I�4�>�83>�n�=��<���=�us=+֎=>rP�I�=2{�=���= �=��=�>�\>�w?�~������y�Q�y��P�:?�A�>���=Fƾ\�??�>>ע���C����M�~? #�?j��?s
?�k��|�>5���.y���= 8��5�*>��=�h3���>��O>�4�By��>���w��?w*@��??�p��UjϿ�_->��7>,>��R��1��]\�abb�\_Z��!?�M;�:Y̾�3�>��=O*߾ݜƾFr.=А6>�gb=Ps��S\�^Ι=�{���;=�El=gމ>��C>���=� ��x%�=c�I=���=[�O>���g�6��|+��4=��=��b>�&>Ư�>�.?�G0?�td?8ܹ>/�o�zϾA������>+Z�=,�>A��=�WC>��>�$8?��D?�K?��>:�=�e�>(�>�,��.n�o��m䦾r�<���?E�?"�>b<?B�rV��s>�Ký�?YP1?�h?e��>��iۿR�"��zO�e۷�����_=&o��j����>�=����<�>W�>Ճ�>�08>�>��E=N��>+&�=�b�=:6>2�����>6�:O�=�=r<�Dʽ��x=U�3�h�C���Ƽ%8s�������Z����>N��>�>�=&�>��=@Py��xW>�z����R�����ف8��]g�;䏿*95�%$��T>}i�=��۽ł���	? �>��X>8i�?�w�?e|�=97�$���J�� "�;79�P1�>f*>�O �d�K�ho�`^�Qx޾���>�>π�>+�k>�,��u>�1�t=G㾁�5��`�>�@���C*�L
��q��>��T����fi�v핻�vD?<��˰�=+n}?�J?���?���>A���h~׾T�1>��!�=�;n�����P?D<'?C�>���v8E��̾�����ɷ>��I�T�O��ϕ�"�0��A������1�>���K�о=3�_��%���ްB�68s�_|�>��O?��?qNa������O����΄���?h?�y�>�? {?`����e�i���=f�n?�z�?6�?�>�ɧ=ނy�7#�>��?���?��?�et?��J�뚯>�̽Q�>�),�e=�t�=c��=R�$>A�?�� ?���>�W��b%���˾�˾� ��	c=�">���>��>7	�>9!>9��=Q��z�>��>Z
s>�}>�~�>�4�>dP��3S��/?��0>���>; I?_��>XЪ<����;ؒ�<6F�W�j����pk���4=O�(=n̲='I����>�̿{�?6�5>3��K?�̺�C�½�r�>�}>E�E�8��>\L�=g+R>S �>�-Z>O��=o>f{�=������>����� ��C��Ba�����k�>l�����E��p!�Q�ɽld�8�þ��:u��{���9� H0=}u�?��v�������B�����_?�;�>pg?��(��1����>�@�>�*|>���G��W9��4�پvY�?X��?�;c>��>7�W?�?��1��3��uZ�$�u�g(A�ie�d�`��፿���i�
�+����_?{�x?�xA?M�<�9z>x��?��%�~ӏ�t)�>�/�}';��A<=�*�>k)����`�L�Ӿ^�þ8�XGF>6�o?�$�?6Y?�RV����(��= �E?X�L?7�q?0<�>�r?a��=�%?a��>�?��%?!�B?֐c?¬�>@4�>�Z�>�w�<���=�����ɾ�Y8��L�k�)��H1����=���:�s��p�(><r��أ����ƻ+�6�N��!���*�=�t���Ŧ>��]?�@�>z��>��7?���Uv8������2/?j�9=s���_��綢�{��>��j?G��?ibZ?Sd>N�A��C�>E^�>�p&>�\>q�>7V�O�E�˧�=�.>�v>�ӥ= ?M��ρ�G�	�������<�7>J��>_2|>r����'>qx��O+z���d>��Q��ƺ���S���G��1��vv�H]�>F�K?��?���=3Y�= ���If�/)?_<?�NM?��?��=�۾��9�n�J�?0�n�>�F�<�������E#����:��ء:_�s>.������7]>�
��޾h~n��,J�x龉�A=Q��U�N=�l�r
վ�}y����=�>v����n!��떿�����I?�p=E����T�����?q>���>���>B�4��m{��e@��ܫ����=���>��8>Y窼���F�����>�)G?]]?xY�?����|Uz���;�?�޾ b���j�j�	?���>�?�p>��+>�ꚾ/���i�q�O����>��>�"5�W�m�}���$ ����>c�?�=��?+	V?ZB?zRV?&4,?h$?��>CN�������&?6׈?��=�U�;(z̽�W��6W�B� ?�O?qG:�	h�>�@;?��?�6?�i`?e�;?mK`>�X�l)9��e�>N�>^AK�������?=�N?��U>dLQ?���?B�>������'��t�����=i�8?n�/?0/?d��>���>9Ѫ�ǅ�=�>�'[?}y?)5�?�g�= V?�&�>�>���=��>�D?�l?s�Q?��s?�uF?@f�>Ӓ<�ȃ�}	����W��8�KkR��ԅ�K{=ƥ�_
�)��<� �=��<6纼5��i�!�c퉽}�.�2��[_�>��s>���<�0>�ľ�O��d�@>���P���؊�|�:�޷=S��>��?b��>@Y#�Ŵ�=���>�I�>����6(?.�?�?e�!;}�b��ھz�K�&�>kB?���=��l�I�����u���g=��m?O�^?��W��&��+�b?��]?h��=�,�þA�b�n��B�O?�
?��G���>f�~?G�q?)��>�e�$:n�$���Cb�_�j�zѶ=6r�>RX�'�d��?�>d�7?�N�>E�b>s%�=ou۾��w��q��o?��?�?���?+*>k�n�=4࿌P	��Ē�t
Y?���>�ڮ�M�0?}�N=�x	�1#�z��� ����^���ϖ��ᙾЎ��|@����>���<���>�d?9/d?E;'?�T澭t��Ig��9L���^�M��9��i�B��<#�\:=��Fp��')�� ���ž,�� �~�aB��+�?�(?2��Y�>�X��a'�%�ʾ�PA>�����e����=p���D=H�W=��f��N-�����?&��>G�>٣;?�[�a>�ۘ1�ҟ6�����̳.>6��>i��>`l�>[꺺g�.�ր��˾ј��ٽN�i>�{e?�\R?q�h?6�ֽל'���w�p ���k��Cg���"=�]="і>2~��v��=:%�:K1��x�D���7z�����	\���:?w��>a�>'��?��?bپP�ƾ�飽��;u>�?5.�?v�?�n�>Y۽��1�Ԝ�>��g?��>�ǒ>[ɜ����tJn���Y״>[�>���>��B>f��!�W�᧎�(���l�?�f��=��j?�9��,�A��>~aJ?�g����;�k�>#p����6�~M��>�S?���=o�W>䀰��� �Bt����4??��?5D���;)�g�h>�?�z�>���>A�?1~�>=�� �>#f7?�3]?��g?��5?�?���=���<�2ڽ�=��kK�=5j�>A�]>�<�=HE>�.��ᨾM�7�Ab�����=O�X��&G=���=a���գ$=��<�c>��ۿ�kK��ؾ5����/%
��O��#�#�����=.��H����v�sU���*��V��!d�ь�TRo����?���?F"��&�������6������ j�>��q��.��Y[���p�wÕ�ؽ྅����!�1P��.i�x�e�C�0?����/׿p西����rN?C�-?}z?�����<��M=�H���(2>yE��C��� Ŀs��j)t?n��>�� ��,���x�>|�>�5c>"^{=�]��s�Ⱦ��'>N�>%2?e>�꒾�O���إ�fV�=`�?�V�?}A?��(������U=O��>:�	? �?>�Q1��I������U�>^;�?o��?��M=��W�\�	�F|e?sx<��F��dݻ��=x=�=�F=�����J>P�>h��WA�]0ܽ*�4>b܅>0�"�l���^�T}�<&�]>��սl0��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?X7H�a}Ͽ�\��*a?�0�?���?&�(?7ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=t6�扤�z���&V�|��=[��>c�>,������O��I��T��=���ƿ��$��z��%=��޺��[�C��쪽�U�@+���]o��W�ܧh=B~�=�vQ>�_�>�W>�Z>�^W?��k?TN�>;o>�P�ˈ��3ξ!��H�������2��ꣾmU�w�߾��	�%������ɾ��=���=6�Q����!��b��@F���.?��">�˾��M���9<��ɾ�����ΐ�DZ����̾~1�"�m����?��A?�5���W�E��m���Kr���-X?�a ���J]��(��=���$�=Vz�>׃�=g�⾩�2���R�5?&�?���sㇾ�4>܂Žv�;L�/?b?L�=�;�>�{&?�\�}<L��x�>�;>��>�8�>9i->����9R"?i�^?"T��*��랢>vǾ�ތ�RX=a�#>��L=��1�e>7���˭���"%��>;�%�={G`?d��>���'��_�����,�$n��t~?�E"?���>�f[?>?�_�=�iҾ_'*��ľ�>|�R?�W?�D�=_��hھ����\�)?��m?�y�>����a/��@���*��r?�>�?'#?46Y<%U���͌�?-�XW8?0�u?|�l�H椿�D!�w���>�E�>h[�>���h�>
�Q?�0��w�����¿s1��ٝ?�y@`K@�o�;�"�L�>�#?,�>우�rX�᫰�|�S���>>�?����Z����C�L٪��@?ʴ�?�:(?���b0�4��=@v��]��?� �?�����@=s5	��Sp��c��x�S�!X�=�,��<��%����j2�Ҿ���Dy�����l݃>{�@��ݽZ��>8%�����Ϳ�Jv�U�߾+�m��??l�>����b����u�	�|��N��D������W>��=�c �7�پ�^��m(����=8"?E1�<P�U=�k��G��<;��]�=��o>4�>d:�=h=齥��� �?3��{��^{�� #Ѿ��u?�#�?�=�?�.?H9�_�<d��Ӧ�=tl?�5�?H{M?����w
�+�=�j?ۇ���c`�$�4��;E��:U>�3?F9�>��-�jO|=C>��>0>�/���Ŀ�Ѷ�q���^��?T��?oi���>v��?;i+?�k�R:���e��7�*���<A?�2>����p�!�G=�ظ���
?��0?���>�4�_?�a���p���-��ƽ"ܡ>�0��a\�LD��%���We����?y����?^�?�?��� #�_6%?��>2���':Ǿ��<v��>�)�>�)N>�L_��u>��X�:�bg	>+��?o~�?	j?���������T>��}?ʅ�>.��?�=��>��=nϯ�_'�+�>In�=�o��� ?�J?���>z��=��>���.�e$G���R��*��B�0܈>�b?�L?m>]>ί��\&-�k���˽S4�V�%��o>��8(�"cڽep5>@V<>��>-�D��־�.0?V�P��u�p���᯽�YG?�Ђ>�+�>� �@.�����=�.Q?�2�=Ti�͹��+�����޽%ק?G3�?���>6��,v�=_e�=flt>�,_=(BI��ȴ��/7��As>�6?�c^�Z���⎿��>d}�?gW
@o��?"Ys�c�	?0��a݈��>����b�3���=LU7?��w>�A�>�@�=զw�M����r�F��>6[�?�2�?c��>�j?C�k�N�?�p@5=�K�>��g?�
?��1;����qG>�[?����ߏ���H�f?��
@Ť@^/`?��ӿޤ����t��&����=Q�=�Y>>�h-�K��ݠ=��ýZ�<6�`>a��>��4>	5C>#�/>Fx$>%#�<v}����[\��	����F���]43��y����#��wX$�v��`����0 �K�I�F5���>�n��+v�u�=5�N?bF?��?Y�??�*�#Զ=�-��v����S:�㈴=���>��B?��a?~YJ?��>��� i��,��&ߑ�W<y�k �>6��><�?G|>�Н>��U>5e%>VZ<�!�>q�>6ww=�!�<
*>�ئ>j=�>�0�>ː�>m�L>ڼ�=��l��Y�c��"��H�<���?yD����a�	��������B���l$>��-??��=X����uĿT�����M?�̲��s-��0��WR>��>?�:J?R�=^Ƶ�h�^�K>WwA��k{��)2>���a=���"��)>��?Ƨf>�Hu>4p3�]T8��P��q���Y|>@6? ��8�x�u���H�OAݾ�M>��>��G�iu�J���:�~��hi�:|=�|:?��?�y���ⰾǖu�����)R>��[>�==�c�=?-M><yc���ƽ�+H�uU/=���=p$^>�u?v�.>��=�k�>���nO�Vè>��;>��'>9DA?�"?�]����ʔ��w^2�\q>�\�>2z>��
>�J��]�=��>�td>h���ކ��]��;��U>����f��mr�z�w=�c�����=���=�$���=�Qf=�~?���*䈿��e���lD?W+?� �=U�F<��"�A ���H��D�?q�@m�?��	��V�<�?�@�?����=}�>׫>�ξ�L�ޱ?�Ž;Ǣ�Ĕ	� )#�fS�?��?��/�Zʋ�9l�z6>�^%?��Ӿ���>O���z��}���2v��+=���>n<J?����z��r<���	?�?�S�Iq��~+ȿmsv��?�>�%�?�C�?|m��J��}@�v�>/��?�Y?��j>��پ~�^�5�>q;>? �Q?�ں>����#�3�?�޵?nO�?w�2>8�q?�t?�E�>����m�����B������`�>\f�]�Z1��fhR�;8���T��� u�h����>H�<p��>\����m��^4�<��K��'�M�����?>���>�i�=h�>u#�>��>K�>]�u=����X��b!��.�K?w��?{���1n��l�<��=Գ^�Z&?3I4?	c[��Ͼ6ը>�\?�?[?$d�>���4>��.迿�}�����<D�K>�5�>FJ�>�'���FK>��Ծ*5D��n�>�ї>�գ�f>ھ^+��\���]C�>]e!?W��>
Ю=Ș ?��#?�j>z%�>xaE�@8��0�E���>���>eK?��~?��?<Թ��[3��	��R硿��[�G6N>��x?�S?�ɕ>�������l�E��0I��ߒ����?�pg?]9��?E1�?D�??3�A?]5f>\��Sؾ岭���>�!?��r�B��2'�4��^?	?s.?�$�>�o�����p���C�F��B�?��[? �%?1!���`�
���L(�<����{��V�	<�~�W>��>m[�����=79>b0�=*0n��h;��h<D�=g�>�D�=�8�U����?}mZ��t��rd7<(���NA�
�b>X>�>Iu���U?����KZ�������^��X�)��Q�? ��?&��?���J�t���c?CE�?O�??�j�>����Ţ����\B��G|����4v:>�u�>���=x����&��[m����ڙ��2X�|�?��>�?�?��N>���>�D��R/���𾱓Ӿ\�Y��C�Z�;��/�����w��$�/��r���࿾c�o��>n����>��?}�>��>���>�
�>�߀>}�>�x�>�ox>��0>���=h����L	�K;P?�O˾
�5��C ��\��W�G?�j?~~?��(��f���}����?<,�?�ٜ?h�|>�%`��!/����>ͅ?�X����>G>�UL�<�k=�[���$(�����Ԏ�-�>u����8�7`S�B�W��\�>%�?Z��dϾ]���D����&�<M=?��?��!��FD��#i�A�S��/M�0-�����B��1d���t��k��T뉿𧃿��$�/�鼈#?ɐ�?3u�F'��{J��_�`��>;�P�>��>gM�>�q>_�>G���5��x���"��5��>��u?�k�>W�@?��2?U�Q?��K?�C�>nŨ>�����>S�=jM�>j ?�8?t�C?	\8?
�?,t=?��>Ng�:��	��u˾�<%?T.?�k?Q�>�l<?�T��,�M��=&��<��!�S�����3=�1� �ʼ#";�f��=��Q>C7?�#�uW8�B���AUj>nS7?Ш�>��>�O���F��L��<��>��
?�!�>m �	dr��s�N��>y��?��mF=��)>��=�����%޺�M�=eK��A��=�ׂ���>��<:��=�_�=4�L�Q�9k;��c;1N�<u�>:�?���>�C�>�@��/� �j��f�=�Y>aS>�>�Eپ�}���$��q�g��]y>�w�?�z�?ʻf=��=���=}���U�����4���s��<�?3J#?(XT?W��?r�=?bj#?ҵ>+�jM���^�������?`!,?$��>e����ʾ��É3�˝??[?�<a�E���;)��¾��Խ��>�[/�_/~����ED��ㅻ����~��*��?忝?A�K�6��x������[��P�C?�!�>Y�>]�>C�)�Z�g�p%��1;>ڊ�>*R?��>C�O?��z?��\?C�\>��8�����|阿 c>��4 >�u??]��?a�?�`y?���>�h>�3)�0��K����z����a����e=�]]>�>��>G��>���=}-Ͻ�s��RP5�7��=sb>��>���>���>�v>�5�<��P?۝?���������������o�`��?�v�?T3L?��:>�
�~V2�r��rE�><�?J��?cp0?�q���>r�:�$��e�¾EH�>D�>놡>�r�=����h>2�u>&�V>�d�1{��4�Ǧ9� O�>�;?��	>�P׿��n�)���-����6罤������v#��e׾J�b<�����������2����謹�M�뾟�;�$���� ?8�=\U>a�~=O�^�2��ܼ�J>�1=�ˀ����dDŻ��"��-�O�ν�y��bX��b�,=��վW1y?#<?\Y(?�J?���>2�H>l����t>�ý��?V?<>߃��|���0�K�m������dzؾ5I��b_��9���d>ټ(�>��S>K�>R�꼂>],�=�&�=Ձ�<��=y�>_��=,��=���=J�=�/>�6w?W�������4Q��Z罜�:?�8�>�{�=��ƾq@?��>>�2�������b��-?���?�T�?O�?Lti��d�>/��1㎽r�=z����=2>���=r�2�R��>��J>���K��I����4�?��@��??�ዿ΢Ͽ)a/>�h7>�E>h�R�hx1��,\�9yb��*Z�\�!?@N;��`̾oK�> ��=�8߾p�ƾ'�-=�6>;�b=[h�lX\�;��=fG{�q0<=�-l=��>iD>�ں=����4��=ٚI=^��=��O>ћ��k�6���+�+�3=˦�=-ib>��%>i��>b�#?�O(?Ow?`��>�*�F0����3�>yS�<$k�>[��>��d>���>�M?�\?U�B?��p>����N�>�j�>Ah#����m���2��.�۽�Bv?��?m`�>���=��a�[.���C���3I)?��=?=?�ѱ>�U����4Y&���.�2���L�4�W+=�mr��QU�a���Vm�.����=�p�>���>��>'Ty>	�9>��N>~�>��>�6�<op�=L⌻{��<�����=&���V�<wżP����v&�a�+�[���J�;��;z�]<~��;��=�[�>�Z�=݌�>���=����VB>��3F���;;�q�GJ�)�v�����S�-���~rk>�x�>����Pʑ��>
?z�J>��W>+}�?�Zr?�k`>�_��4�[_����!��� ���>�">�m�3;?��@t���n�6&�o��>W!�>�~�>��k>�,���>��nw=��oR5����>>Ō� �Y��aq�,��|៿�0i�_?K��D?����{�=O�}?�I?˚�?Z�>�H��~�׾�0>�M��A�=���-*p�>�����?�&?Yy�>����D���澕@㽯&�>�u_�b@T�Mu��O.�&ͮ<�����x�>ȠǾp����C-��΅�(⎿��B�[=��'â>�>C?�P�?k@�49��zR�a�	瘼�?~@z?���>_w�>�#?v���xa��\�Du�=g�h?f��?gD�?0�W>,y�=����G��>�	?h��?��?�t?�?A�:p�>6�;{!>2���и�=��>���=�N�=�R?�[
?l�
?i���r#
�y��$��_�� =�4�=RÑ>U��>>�r>C�=�Eg=�:�=X]>��>3��>��d>ۂ�>���>'о�&�H?Mč>��>�Y?�u�>�e�Ŧ�;]󄽟V�=/.��wf�Kt����_���S= ŏ=�=	Z<?��>p�Ϳ��?߾r>�2.���'?�޾$��fU�>�o>շ���>w�#>��@>��>�o`>�>��>�:�>���2�=�~��� ���E���U��p׾��}> ;���,� K�:-Ͻl�C�+.�����Wi��g��:�=���^;$�?�|ѽ�Ur���+�	�͍	?��>��C?�gV��C����2>Zw�>��q>����������zپ���?ĩ�?�;c>��>N�W?�?��1�43��uZ�)�u�g(A�e�V�`��፿�����
�����_?��x?yA?CR�<":z>N��?��%�Fӏ��)�>�/�)';�k@<=i+�>*��P�`��Ӿh�þ�7��HF>x�o?1%�?hY?oTV���N���>Nu3?;"?�k?s�%?K�\?�L��?�r>���>�k?%�@?�=?��>�T>�D>�=���=׫������~o��>���Or�.'=��<g.K:��a�=� ^�d�I����<�_=8C��o��<Xlm=Fo=̥=�ͧ>��]?���>Xم>�H7?�^���8�������/?�xI=-v��x��ء�^a�	E>�Xk?���?�YZ?��c>�$A�o�C�m >E��>&>co^>"�>����G�Tǆ=|�
>�>r��=G�G������Y
��Ñ�ݺ�<r{ >-��>1|>�	���'>H|��5/z�<�d>�Q��˺�(�S�v�G�=�1�ǂv�DZ�>��K?(�?���=�^��'��If��/)?�]<?1OM?@�?��=�۾u�9���J�M>�+�>w`�<��������#����:���:��s>22��*_���e>0X��� Ͼp�a��~K�c@����<���n�<�@�}Ҿ3$w��D�=��>	L�����B���b���G?���=�T��A�B��)��]��=$x>ϯ�>�d}�ڳ��64��Û��/Q=D�>�A/>�ۀ�����?�C�����>�gH?�P?$ȣ?9��<%q���#�����쾤b��@?���>�#�>Q0�>˯�>�v�:�
��j��N����>P��>���~p-�Z_���k�8�;�!��><�?�._>d�?��T?�?<K?��/?���>���>�Kf=�����(?A�?h�=��=���T�T��Lm� ,?�mX?#�<�Z�>�?e=%?NC*?!m?�l&?�y>L���]hZ���>D٫>�c?�	�Ϳ�l{���t?�gv>2t?%��?��>4W]�oZ�A
�=-�r=O��q�6?�$Q?�LT?&��>�^�>O���P��=���>�b?d*�?��o?Y��=м?U�2>K��>x=�= ��>���>T�?�!O?��s?��J?��>���<���'
���Uq�)�^�U�;�<=<��q=����Tu��
���<x�;5͸���c�P4��G��=�����;�f�>�t>7��j1>^�ľ�U��8�@>���l	��w銾n�:�E��=6��>	?Pە>F#��Ԓ=���>MC�>6��w*(?��?�'?�M.;��b���ھ)L�v��>W�A?�0�=�l������u��h='�m?m�^?B�W�����b?��]?�X��=���þ��b���x�O?��
?��G���>��~?��q?��>��e�7;n����DDb�?�j��ʶ=�m�>�V���d�o>�>Ø7?R�>��b>�5�=�|۾c�w�<h���?��?��?���?�0*>�n��3࿯"ܾ�k���\?P�>���@%?@;u,�ov��0����پ}Ѿܼ�=������[.�Pɇ� _�����=��?�?b?��q?i`H?��2�`��i��|�(G��3���YU��2(���.��ac�=�'���i���Áy=K���(1��?�c!?@B����>f{������1�K��=����"��=^ei�^�=i=�Fi�d�����;��?E��>E_�>�D7?�R��w<��o:�S�,�Z�>>np�>I �>��>�bH�x<��<���۾c~���@�5/i>�`?q�m?{�W?�������$}B����Aн��D��=5B>���>J��x����"��U>���������|�㾖��Վ[?x��>�|�<��?F�>��龹����#��{���^���>Z9v?Y�)?��><�h��EB�#��>|�l?��>g�>r��sO���z��hٽ(��>F²>� ?K�e>�����Z��~��tǎ���:��]�=�eg?*���Kb�֣�>�O?�E��Ghg<y�>��h��R���a$,�sC>�?�I�=�xH>��¾�`��z�c���zw8?�o9?�D����>��A�=��?�>�$?�y�?���>���T�x>aU?��Y?� Y?�@L?6^�>�N\>�ҷ������/��^7����>�LY>R:Y=���=��1�z�S뾂L���>Ԙe�fV���=?�G���@��D:�侃>ϻؿxE��%˾I�
�>�߾������b��Ȗ���3��T¾厞���m�"����]ͼ�FJ���X�$���̀����?���?G�[��'h����f{��,��
�>u�����@��=P��n��
PپCo���R#�G�L���n�_�k�ſ(?�o��I�ǿ�a���E־��$?ך#?�!{?�|�s'��8�{5>��$=�Y�:�%ﾔ*����Ϳ�˕��Hc?��>���T������>�Պ>o�]>��j>w:���ȟ��T�<v?�,?�M�>��j���ȿ�l�����<��?�@�}A?��(�l���V=4��>�	?��?>J1��H�4��Q�> =�?-��?t�M=��W���	��}e?a�<�F�mKݻX�=2�=V=�����J>"S�>���]UA��2ܽH�4>}م>Ʉ"����Ն^�S��<��]>��ս�)��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��=�����&���] �+v �Y�r=���,���_!���	�@ �N���鋃�n�ڽ�4u=:��=V�N>4�z>.�>"dG>��P?<�s?�6�>��C>�z��J$��)�ݾ̏���é��`��
�����q����yʾ�_ƾ���$���/)��[��"=��=0R�Z����� ���b�u�F���.?�]$>��ʾ'�M��-<�kʾ񹪾�����ॽ�*̾6�1��"n��˟?u�A?��E�V�Y����=���.�W?T����嬾���=����[|=$%�>0_�=���#3���S�N�1?�O"?�F��7ȁ�{C>�{��T<ʚ+?C�?�F�)^>� 8?�X���ļ�u�>N
s>��>���>�6>B"�����c�?
�e?�a���d��b�>��ﾽ	]��+�<��@>3�C��GC��'|>��=k;w����:�cؽQ|8= 3W?���>�)��T�T���Ŝ�߇>=��x?4(?�~�>��j?b�B?{Ϸ<�I��)S��
�`=y�W?�h?��>ڋ���о|���{5?O�e?��P>_/h�
�꾇	/��E�c�?8�n?�??���@a}�( ��+���6?`�z?n�U�k��] ��!���>�z>�_(?���l>�m?�ᄾB��VĿ�Z&�NԞ?"�@��?���y	��s>�M)?�o�>�*�"��u���@�����=?�ﲽ�҅��7�E�ɾY�@?�.�?%&?,�D���/�O>󱗾�K�?���?vs��I=9x��T�����x���HH=Ee6����S ����5��g߾�������hH��CG�>�N@B�����>�4H�_ڿ�oʿ��q��۾�|��w�?E��>�NC�������������TU�b^E��{�ġ�>r�>�����
���b|�w;��T��5�>H���Ƈ>��R�r���gȞ��a<{�>�|�>��>Y���,��\*�?n#����οA�������Y?,�?]Q�?h4 ?M�<�u�Hx��t���H?�r?�X?>p�yCU����ؿj?�b��"W`�̎4�EE�RU>r!3?E�>>�-���|=�>���>!`>#/��Ŀ>ض�]������?Љ�?yo�S��>��?Rq+?tk��7��_����*���,�G;A?32>���b�!��3=��͒�`�
?6�0?�p�D2�]�_?*�a�N�p���-���ƽ�ۡ>�0��e\��M�����Xe����@y����?N^�?i�?ҵ�� #�f6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?W�>%�?�n�=��>�t�=�ǰ��1�÷">���=�6<���?VzM?�m�>�_�=��8��</��bF�VNR���@�C�Ͼ�>�a?0�L?`%b>mv��*i/��� �̽_2���R ?���.�O�ݽ�&6>��>>��>��E��`Ӿ��@?YmF�}޿����@U>��\?䑝>��?��־��������z?`D_>����`��}D���%�ԕ�?�@�`�>���������<�)P>�� =3��7�p	`�q�>9�T?��jR��C���ߒ>���?F�@��?k��hp?�	�P���U|�z=��^d�d`�=��<?��龤�`>GS�>2'�=��y��D���r�y�>���?��?v��>1`?x\�=3��w�<��y> `?���>1�=���>9>�?z3�����&���Gi?�@'�@H^a?W���\�ҿ^�����Ӿ�	Ӿb�P>�6�=پa>�'���}>u��=����)�D�>m|�>'�> ��>�qz>��$>A7�=Nـ�9m �h��0�����)�����@��ԭc�����
=���	�(eվ}JӾν,���@�cV�{�ʽ�j�=�dV?{�M?��?��?/�]�_N>�e����D�s�=D�>�!?�WH?,�2?%�=�����p��T��1]��N��0Ӈ>�l�>�?�mh>ύ>��5<;u�=�t>���>;�>n�=�W=vP�=�an>;&�>���>�I�>�C<>��>Fϴ��1��k�h��
w�r̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?�d>�*u>��2���7�6FP������z>��5?����YS:�ܢu�$uH�cݾ�M>���>�{N��O����!C�{
h��C�=|:?qk?w��2&���Sw�i���Q>��\>p3=�̬=L>d�i�0|ƽƼI��l'=bO�=
%]>Ts?d'>�S�=S�>{떾lnF��!�>{7>�S*>KZ??Q�#?d�i��������0�,v>���>��>��>��E��=G��>0�a>pv��Ӂ�����J��k[>_ȉ��]��㍽u�=q���4�>�L�=���7�A��4=Й~?g{���숿��!����D?�N?�6�=P�F<��"�]����Ƹ��?��@rM�?�	��V� �?�S�?Pm����=�<�>��>Σ;�;L�N�?�ƽ�Ϣ��n	��w#��A�?��?�-/�mȋ���k��>aY%?�KӾK��>��pΔ����w�q��X]>h
?X�y?k���o���� �ֲ+?ё?.S���l���ʿ�Bi��y�>OU�?g�?u���
��ny��a?T�?�S|?�C�>r/��ڞ���P>�xZ?�d?�?5?8�:��I�B��>��?�=�?��`>���?8�?��{>�^��&f��D�������~�B}>���>�/��%$n���K�*ߜ��鎿����5��=�>|�{�I�>
�=�����A�� :��~��Ǩ=�
=>�A�>��8>�ּ>0S?��>R��>�(�<@�<��]��4:�}�K?��?�����m����<���="�^��O?��4?`�s�s�о�"�>��\?��?QU[?n�>�j��뚿��������=e�<1L>xO�>�I�>bȌ�GK>y�վ��B�c��>D�>�^��2�۾�R����,���>�!!?���>��=�� ?��#?��j>�$�>~bE�f9��H�E���>.��>�G?��~?�?�ҹ��Z3�����桿��[��6N>I�x?�W?�ƕ>�������ƢE��I�ڒ����?Kug?�]�{?�1�?a�??ܦA?�$f>��Jؾ[������>��!?���A��M&�'��~?�P?���>�7����ս)Mּ��������?�(\?wA&?Ӝ��+a���¾19�<��"���U���;N�D���>[�>���m��=l>Kװ=�Om��F6�$�f<l�=��>��=�.7�u���+?/�.��ZY�q��<ǒ��C4�w.�=� �>��y���h?��H>Zir����������^m��(�?(�??��i�i���A?g��?��'?�k�>D'ž�΂����|Ma���+�q|6��T>��>��=8�����]4������������>�^�>6�?��?��d>Vu�>����z�*���J@��xV�]K ��E?���7���N�����噂�˔��W����C�>��q�X�>��?=��>� >�`�>���<�&�>~rG>[��>Z��>��O>�>��=�O���J̽�SZ?�k�ۓC��?ܾfsW�t%k?z�w?��?@%j�p���?����??7�?�פ?�}�=Y�{��G+�a
?Y6?"?/�H�>(����+=�+>ɟ��XQ�hB=��m��6[�>�	$�Z�,��{J���f����>Q�
?C��������X<VV��d�=L�?{�?κ���N�1�~��3c�&�[�����e�pڷ���w�d���������*�B�cV����!?z߄?�lپ�}�Q���+R���1��>�Q�>|�>��>yh~>�ξ:O1���}��I0�U2��sL�>Y�m?r�>�iI?:P/?
�T?��A?y[>�X�>���i�?T�;��_~>�f?�d.?)�9?U�J?t1 ?nj&?0oN>�õ�����ž�V.?��+?e' ?/-�>� ?[�ľ-�,���F;�E='��Z�I�7�=9�:=�Y�gu-�sR�<{�Y>�X?}����8�Z���ck>�7?��>e��>:��.�����<��>��
?G�>� �~r��b��V�>���?��� u=��)>N��=Aw��J�Һ�Y�=&����=���x;��b<:~�='��=Ut�"G~��S�:��;�u�<�t�>�?���>�C�>�@��� �:���e�=iY>MS>>Fپ�}���$��[�g�^y>�w�?�z�?4�f= �=H��=e|��-U�����A���%��<��?(J#?�WT?5��?2�=?Kj#?�>�*�ZM���^������?w!,?��>�����ʾ��։3�۝?i[?�<a����;)�ߐ¾��Խұ>�[/�i/~����>D��텻���U��6��?�?MA�W�6��x�ۿ���[��{�C?"�>Y�>��>U�)�~�g�s%��1;>���>lR?���>��O?�h{?�}[?q�R>��8�I�+����3K���">(@?��?EՎ?��x?
J�>�	>9�*���H���О�>��L���\=��Y>�	�>���>���>���=�6ʽ$����<���=8�c>[,�>�٥>�>�3v>�5�<�SJ?�?|)��������ĸ���gǽt8{?�{�?�J?�R�����0#���ʾ��>�?�	�?T$5?s����7�=Kb_�<�Ⱦ����>c�>T��>u|�=��c���$>��>\�>N@��hM��5�V��T�?��D?s+>�¿�c�]�@��Ċ�v~�<K۠�DǄ��fͽ���N9=���i%�G����Q�d����{������������>��>37�=�G>���=�<�uP�(�Ѽ�\3=M�t�|R=�"�v�=Y����>����m�Q���ּ��<����5y���2n?��=?�x)?��G?�;�>iP>�����[>$1p�B0?r�)>����]ξ��������s��F���d�ھ1bX��ٸ��E>�����>$yW>�g>����O�>���=�`�=E�;y�
=i��=�� >r��=)��=*��=0�>�6w?W�������4Q��Z罤�:?�8�>�{�=��ƾp@?��>>�2������}b��-?���?�T�?B�?Dti��d�>G��g㎽�q�=a����=2>u��=~�2�T��>��J>���K��H����4�?��@��??�ዿϢϿ3a/>��7>p->�R�uz1�|\��b���Z���!?�O;�sJ̾x"�>5ݺ=Q.߾h�ƾ�.=!h6> b=���:[\����=��z�<=D�k=�Ή>�C> O�=�X�����=�J=��=f�O>~-28��p,�A�2=���=��b>&>���>v_?�3.?�.o?e��>�(���PӾ����fN�>A��=}3�>�1�=gF>�>�:>?jyC?
SF?V��>�7=(��>��>8�(���r��>�b핾������?��?�c�>n�����?��?�;�;s����?,r5?LQ?��>��-lԿpkH��5A�5x~=��>���>%�ھ�=ǧw>�� ����0:�:�>؏�>�1�>�k�>�e�={u3>.�>na>��=�[�<��#������\C�����'��~y=���=:˼'�<���Mݯ�����*��I�ܼ�5=�T�=�&�>��>`
�>��C=����Sq
>��r��=�y�L=UB����8��Fq��Ņ�z�6�Z(	�e>6�w>�Q�����L�>@�/>9�F>$�?k�v?$~w>�u�'������N����:���j>B�7>&�����K�e:n�V�<@ɾ���>��>d�>�l>",�?���w=(�ga5���>9u������5q�\=������i���ںs�D?JD�����=�~?ϰI?Vߏ?��>�����ؾsF0>�R����=J��0q��E���?�'?��>�쾗�D��C̾�����>�ZI��P�������0�m���߷�Bs�>;몾��о�3�'g����0�B�dzr��ͺ>&�O?I��?Rb�<_���\O����)8��,�?��g?C�>�5?�=?�ѡ�)A�C���=z�n?٧�?B�?q{>�_�=tD��AJ�>��
?�Е?��?G�t?IL�ˏ�>�&�<J�>������=ƚ�=ߒu=YR�=��?�	?Ǆ?u���6��}��j2꾲f�s�=�i�=�!�>��>1n>���=��3=�L�=�6U>�s�>�ٍ>~�Z>x�>�"�>&���l��J�?�@6>��>x>7?3�>9��*��!�w=l�B���J���r��7$���4�=	3�<wG|=��%����>��Ŀ"�?~U>R��[?'-��ǧ��׀>�>�s��
�>��R>T�^>q>�>N��>v1�=�xN>��A>�dϾ��?>#��=6��7M�3	Z�5R�(�u>�k˾_�O�Fu�a�F�7��޾�0羆~t�W��ĂA���ϼ�;�?1>$�y����:��Yj��G"?���>a{?���u.�Uf->�u�>���>~{��di���͈����b��?<0�?�;c>`�>1�W?4�?R�1�"3��uZ�C�u�<(A��e�$�`�z፿����
�����_?��x?�xA?~Q�<O:z>��?��%�(ӏ�G)�>�/�;';��:<=v+�>g*����`���Ӿ�þ�7�RIF>�o?�$�?Y?�SV�}k[�5��=�=?
5?��n?Z�!?wxa?M=#�j�??�8>v��>��?� >?�??��?Pd>�=aM�;!5�=%Rj�{���t꽧z�����3=�-�=�%_=	�溠0�<�̂<���ٗu���=���uY�<��d<�\=���="�>��]?���>���>Zm7?w��YE8�d󭾗�/?hoC=�%���+���衾PU�f�>&k?c�?ہZ?�Yc>]�A�xC�X">`��>�K&>�p]>�K�>���b�F�5Q�=L�>��>�֧=�L�8�����	��鑾���<{c >��>�5|>)��^�'>Cy��5z��d>��Q�Rú���S���G�=�1���v�q]�>��K?��?���=�^�*��3If��.)?�_<?�PM?-�?� �=�۾��9� �J�:�i�>�(�<��ྡྷ�"�� �:��v�:��s>�/�������i>�h��Qؾ�]m���M��G꾅�-=���1>=('�Z�Ծ��s����=�>-�þ��"�}����]����I?���=@�����T�������	>9�>'�>Q�C��'B=����iR�=���>O)5>]�Ӽ���P�D�E��>�y=?[
s?lЋ?�ys�i۔���3���r.��k���3�?�!?�?��v>�څ>�_���8�Z�z�mlv��T�>4��>�'�4�#���/����=�_�l��>�,?&���N�>eu?3!�>YT1?��?鬟>��=�~ɽ�d]�s�/?E~?k�+8�I㼛~��_�4��E��m](?s?F;�����>E"0?|�%?�p?ށo?YE.?u<>�î�s�1�r\�>ZӠ>wr�ң��R�=4iV?��>?�?�H~?	�\>փ3�������;<>�>���;K�?-?��??���>>��>p���Z�=c��>�c?�0�?��o?��=��?�92>>��>'��=���>ъ�>�?XO?��s?��J?���>��<C9��i6��>s���O����;AwH<�y=���K/t�JK����<��;a��.=�������D�������;���>m�t>R����2>
mľ��U�?>7����-��z����g:��=�>+�?X�>C�"���=��>E�>i%�;�'?ݫ?��?�F�;��b���ؾ�P����>D�A?��=a�l�Ԅ����t�7@h=T�m?fI^?m"V�����8�b?�]?�g��=��þ��b����I�O?�
?��G���>S�~?M�q?���>�e�+:n�0��Db���j��ж=Sr�>)X��d�O?�>G�7?�N�>8�b>A%�=�u۾�w��q��y?w�?
�?���?+*>x�n�R4��ƾ�X��۶l?�h�>��۾��(?Q>�� j>��b����꾔(��e:���ѵ�n۹�@�UY����,�'1ɻ�Y?�X?M3u?\�5?��� �O�ܥE�S\�
ub��J"�b���DJ���7�l�U�4u~�������}���|�<y��9�1����?�Q+?� }���>�W|��� �Ojξq<X>�aɾ�۪�w�>�#��
�=��;Ƈz�>km�[�¾m#?���>�P�>|'2?R��F�[�-��5�M����>V��>�Ъ>���>�˪���#�(�뽍�̾�����N�P�q>��h?$8b?��U?�0W������s�����ǧ��ž��0�=m	����><	O����t*�6N�J"w�>g!��q�,�	�A<s�J?vn�>Ɲq>0��?�V�>�Ѹ��n��9�1�'�
�z�<�}?�:d?���>
;�>��1=U��+��>�m?�>@��>Ҳ��Š�W�w�)@ҽ)�>W��>��>LA>��*��r]�D��������@����=?'f?E?��g�R�oc�>��N?��E�&�;W;�>�}I�Q5�%P��x�-�%?�=X_?�x�=��I>!嵾�q�HBy�a����k;?��?�־\#�e�>��+?��M>Ya?`/�?SE�>S 
�7��=� T?N�\?cKP?��*?�}�>��>�4�=��ͽb�|��v'=U�>4�i>��2=;h�=k\��2��3�W�nnO��
�=[�ƽT=�" >���⽟�%^轴��=H�п�yB�:��F��p��v3��E����T~���V���m~�J	*�5�c���a l��g_�e?��PO�*��?S��?w?K��0)�QZ���ሿa����>�7}�F ^�,'������W�z��ǔ�!%�%�M���r�j=u�T�'?�����ǿ󰡿�:ܾ5! ?�A ?>�y?��:�"���8�9� >�C�<�-����뾮����ο5�����^?���>���/��g��>�>D�X>�Hq>����螾�2�<��?8�-?��>ߎr�+�ɿ[����¤<���?/�@^|A?~�(����7V=���>?�	?��?>>S1�zI����aX�><�?t��?^�M=Q�W�*�	�;e?uc<I�F�b�ݻk�=�>�=v[=;����J>�T�>7��RA�n9ܽ��4>�݅>�v"�@��D^���<��]><�ս>:���؄?`8\�K�e�E�/�)m����>Y,U?�l�>'�=k-?ɍG�b�ϿQ+]���`?��?E��?�h)?������>�+ݾp�M?�!6?�a�>�&�u�e��=�伢ٓ��侰�V���=<B�>��>+�,����¥P�L���6i�=�����l¿v��`:�Ѧj<�򭹨�����v̳�vQ�������_�;�½�*�=���=�9>��>�SL>K�r>��\?qJr?>g�>�D>���ԣ�EXȾ�{���S|�uz��yQ��������*����Q˾ږ�������`�ԾS =�h�=�4R�{���{� ���b���F��.?ku$>��ʾ�M�C�-<-lʾ���{���n쥽�/̾#�1�"n�5͟?b�A?����n�V����~|�(�����W?�N����j謾f��=�����=s"�>��=���o 3��}S�^_7?ۇ?�H̾0qR��.>^��&�z�ŝK?��?�1H���z>N�?���$-L=~��>�:>c�>��>�L'>�
ɾ�-۽!�6?�l?��[���ȏ�>B ��Jo��o��<^�_>�.k�>�G�~n�>1�=�u�i&�:�"��=�;�[?��>�2.��s�ɢ�U�n9Ax����?Q)'?��>��T?5�8?�>I�;��6��d㾭f�=Ӝ`?�[c?o�>N|����ҾWG���-?~}n?t�>�������c�&�-Z���?qq|?(l?��~�����jp������N;?I�?.<X�����m*�J�h�+/�>N�?z� ?�8�'�>�Ё?��#�6Z���]ſ��ѧ?��@��?��=������(>��?0�>��޾�^��'��=Ё����=5�?VI��Z��gLA�	?�<C�W?t�?��%?�鸾��8i�=����ܬ??+���V��<e�%�l��G������Y�P=�_�6�T�P!��F�;�F�ɾ8s�`צ���(��l�>�B@1�ܽ���>�b)�v�ݿ�.Ͽ-^~�w۾aʆ�v@?�>�G��h˯���n��r��-I�]GF�S���M�>7�>����w�����{�Rr;� @��k�>�	�>N�S�p&������5<_�>3��>:��>=.��a轾*ř?'c���?οH������ �X?�g�?�n�?\q?��9<��v���{�\���-G?�s?�Z?+n%�p;]�k�7�%�j?�_��xU`���4�tHE��U>�"3?�B�>T�-�f�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*�L�+��<A?�2>���J�!�C0=�TҒ�ü
?W~0?{�g.�]�_?)�a�N�p���-���ƽ�ۡ>�0��e\��M�����Xe����@y����?M^�?i�?ҵ�� #�g6%?�>d����8Ǿ��<���>�(�>
*N>mH_���u>����:�i	>���?�~�?Pj?���������U>
�}?�Y�>��?s7�=�S�>�	�=����f�(�� >�z�=��;�.?��M?��>;I�=��7�J/�MF���R����9C��ш>!�a?d�K?Kb>뺻�݁9�� �a^ͽ�2�~�Լ1?��}+�E"�05>9>>	r>�E�ԬӾ�g6?�.#��B޿����*V�=�:?s.y>��?���B�]�ih�MWt?i�>� )�a��4���X(��0�?�@��?����]��=�>kG�>���>���Z�>��o��U�>�6?�Q*�����4���&�>�*�?��@��?�s�:�?��
�M��㥁��þ	����I�=c~=?��龘��>�>��>4{��>��-�r����>���?���? F?�LZ?��`��+�<5i=!H>�Mc?w�?m	~��D���dZ>�y"?G�y��ol
��rk?Ԅ@�@�J^?�Z��i�п벡���Ⱦ�i��n�=[��=��>���4��=C�'>�֊�A�4=�,�=���>b�C>>՚>��>�[�>tA>����!�0���;��@�7�~��Y����`D��
��G���g�ݽ����)�x��ؽ<Ի�V�xX;.ꏽ&�>?�P?b�Z?���?pk?0ͽ/��=L�Ͼ��'=A����>��o>m�(?��N?W� ?�";=ֲ����K���������#�>Kz�>�-?�U>G��>�%<!>jUv>�2�>�d�>�<�}5����=��>?��>���>n�>�C<>��>Bϴ��1��f�h�#w��̽-�?x���U�J��1���9��ͦ��i�=Ib.?�{>���?пe����2H?$���})��+���>w�0?�cW?<�>����T�0:>F����j�)`>�+ ��l���)��%Q>{l?�f>?�v>��2�Q]8���P��ܯ�Ks{>�5?����{9���u�>I�^�ܾ�HK>��>�Z���
����~�i��8{=�`:?k�?����]а�oeu������R>܂Y>8q=�=�JN>�\���Ľ�-G���1=�1�=�[>�%?	-+>R��=�c�>�𚾯�L�E�>��>>-�.>1�??�$?	��xԙ�Ҹ��&�-�S�u>���>�B�>|A>YH�c�=T�>7�`>�3�nP������TA��X>�`{���a�H΀��u=�J�����=渐=@K��&?���=�~?���(䈿��e���lD?R+?c �=.�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>
׫>�ξ�L��?��Ž6Ǣ�ɔ	�-)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ"��>UV���䖿-H����W�#�Y����> �u?���͆���$����?F�?E���K����̿�a��v�>6��?��?rЎ�����B�H���?4%�?�gq?T,�>HB�R��X�c>�AX?��2?e��=n�*���6�[�?���?�N�?I�U>9#�?���?d�[�U>B��L��n����\�G����,> �&>W㻾Nʭ���s�@���bϑ�g�����>�<��>��@ʦ>!�������<�8r�|�B�G� <�5w>�%�>}G>��>�>�H�>���>0E6=��ӽW�����v���K?֭�?L���n�7��<tܜ=��^�k??�O4?8�\��Ͼ1Ө>��\?�À?�[?�^�>����.���տ����.��<��K>�a�>�J�>����yuK>��Ծ�TD��`�>��>r����oھ�􁾏c���8�>e\!?.��>雮=љ ?��#?ɖj>(�>4aE��9��d�E����>���>�H?�~?��?�Թ��Z3�����桿��[��:N>��x?V?Yʕ>[�������lE��@I�����\��?wtg?�R�)?02�?Չ??=�A?<)f>���ؾ�'�>�!?Q���A�3N&�%��~?�M?���>�;��i�ս��ּ ���w��o�?�&\?>&?D���+a�'�¾�#�<U�"�hTT�C�;��D�%�>m�>����y��=>�Ѱ=�Qm��A6��Og<�w�=h��>��=�17�@�����5?aC<�u�������1q�҉*�T��>�k~>�����V?�+�$φ��#����� f����?���?�ט?�ރ���w�r�I?��Y?_�?��"?\�վx~۾Ш��μ�����%O����>:	?th0=�x�Z챿?��6���TW�z���	?|��>��>�8?37�>옽>���0pT�	���ξ�R�5�S�8�s�>�<���㢾.uu�\�(�������S����>ј�<)��>�{�>�T>�B>1��>)#>�c�>�,>/��>��>R�q>�C>��>�v=�E.�qMR?������'������w1B?bd?�G�>�h�Ɇ��M���?���?s�?	dv>ouh�s%+�'m?>�>����i
?s�:=�u�#��<t]�����R���m����>�׽ :��M�If�>l
?+?���ʄ̾�H׽;v�}��=G\�?O�?��.��P(��S���P���M��?��KD���ɾ��!��D��aD��#0������$2�,Z��R(?��?�H����� q���R��Af���>B�>�1�>Q^�>�>6%��7�a�i�^.�n֥����>��p?��>�BE?�M:? q?��R?��Y>�=�>8L����>Ve(����>���>{�2?Q?��I?�H?�1$?�>sP��������j�J?@�-?x�)?�d�>�?B/��S����l��U-���ۼ��=���ݡ<u�B=1LL=L�t>�n?���8�������j>w�7?���>�M�>zT������ŝ�<E$�>�?�p�>���dCr��<�hw�>���?.��W;=p�)>�Q�=['��vQ��Hj�=��¼-��=�l����=�<�$<�[�=�ѕ=�PT�����(�:�X;皮<�t�>9�?���>�C�>9@��� �F���e�=>Y> S>�>�Eپ�}���$��w�g��]y>�w�?�z�?P�f=��=���=�|��SU�����D������<�?_J#?+XT?U��?v�=?Yj#?�>�*�\M���^�����Ů?l!,?;��>c����ʾ�񨿯�3���?h[?z<a����;)��¾�Խӱ>�[/�O/~����:D�󅻸��)��*��?�?�A�N�6��x�Կ���[��:�C?�!�>�X�>\�>�)�I�g�O%��1;>���>(R?���>�O?݃{?�i^?%�\>Kv8�[���Ș�u�O��x!>[dB?���?_x�?�gx?���>��>��(��h�|�����������Ɂ��k=��W>�B�>���>���>k��=��½ԕ���1����=� [>���> U�>��>a}s>��<c�H?��>�Q��vt��q��1��m����y?"��?#�+?�'=.�8KA��}���t�>tv�?���?ɇ+?d�P�°�=���a����|�{ʵ>�0�>f��>��=:%4=�>-�>촼>8������9��sk��8?%�F?�~�=�ſueq�*�o�\&��CQ<Ca���c��%��5J[�
-�=L#��<"���3OZ��'�������ʵ��'�{�?��>}�=��=^]�=���<&�Լ��<��H=o��<��=%m�>z<��6�!}������*��}Q<�D=Ŭ��rʾ[+}?�UG?��)?��F?R�>B�>;GG�c�>;P���}?$�R>�f^�,�����A�4ɧ�2�I�ؾ� پ�c��鞾��>1�3��_
>�1>��=E��<o'�=j4�=��=�ںk�'=X��=s�=r��=��=��>��>�{?� w�'����7Z��nP�q�D?߯�>4\�=�ҿ�gK?�T�>$���Ŀ����q}?h��?��?=�?�#7���}>�M_�iR�:�z�=���γw=�>J�`-�>�Ma>�-�*ޞ�C��n�?�?�??"A���<ȿI>u7>�>��R�"{1�R
Z�Mba���Y� J!?�;��~̾b�>=Y�=�A߾��ƾs*=oH6>�]b=����\\�=9�=n�z�N1?=%n=�r�>��C>Ξ�= '��Ge�=��N=�\�=��O>�^���}6���)�k5=�l�=�c>�&>d�>�?wT0?�t?���>�Ԋ���h����>���=��>�8>zj>�>�>4�C?�6D?9�;?c��>��<{��>ނ�>��;� ������ƚ�Y{Խ)�?�E�?1[�>��*��G���9w;��E�m\?j.?�4?}��>�i��`�ؿd-�$��������2<шe>����Z �G��>����|�*�z9H��j?���>ۨ�>� �>�`^>_�>��>�cB>z�{=k�{�������=I�)���
�m@�;i$0=?s�<s�=p8�=<lw��f���O��������N<S>.��>��Q<C��>
�>	>���D�>훾)8j�Xj^��O۾�(�g�i��qt���3����P>�+>P%�}ᖿ �?3�+>�)>w�?�y�?�Ѹ<V��
���Q��S�����˽U�K>�W�=ճ��hrb�T���n��Z���>y��>�!�>�rl>,�?�!�w=�⾄g5�t�>~��|+�P��9q� :�����i����(�D?�?��«�=�~?��I?֏?zv�>$�&rؾ@E0>�a���x=%
�M�p�� ���?)'?p��>9���D�oH̾����޷>�@I�+�O���_�0����ͷ�폱>������оY$3��g�������B�Mr�:��>�O?��?�:b��W��[UO����'���q?�|g?�>�J?�@?B%��z�r��hu�=��n?ɳ�?W=�?>���=퇫�d��>�b?���?���?1xs?��A���>��;�v$>�M��/��=>��= �=3?�	?��	?�����	���<��bve����<"��=fǑ>�-�>v>*��={t=�ܥ=_�]>���>���>��e>���>�A�>� ��eľ��?4�=>?�>�A8?�t�>C�ĽR�I��H��l�!=M�����S��X���"�Fw�<ao=^V=��u���>9ƿ9�?��>,�F����>��������>�2�>L�9�5f�>�">�J>�:�>sa>[�X=6�A>j�>p���ˀ>}��J
��i$�׹�����B�>@��o����B�(���Ͻ�]e��־�V���$���K������?A�`���}���H�q��?k�>�k?��<����C>l��>��g>�F'��&��!ۋ�㘔�V��?\�?�;c>|�>��W?�?��1�D3��tZ�'�u�:(A��e�o�`��፿򜁿]�
����E�_?��x? xA?�E�<99z>y��?��%�sӏ�*�>�/��';��J<=�)�>5+����`�<�Ӿ�þ�9��DF>��o?�$�?�X?�RV��j��(>X�:?��2?��t?�1?;?����+$?CE3>�?��?}05?��.?�
?3>:#�=fEӻ�z=�Ց��;��m�Ͻ�Ž���6
,= x=�N����<�=X��<��ȼ�[̼9�+�뒼/��<�4=b��=�{�=���>֤]?qC�>y��>U�7?f��bs8�'���'/?��9=����������>��>��j?/��?^aZ?�Xd>��A�|C�� >j]�>�]&>�\>�f�>���|E����=%C>Je>L�=�:M��Ł��	�e���+�<�6>�>��|>�Z��*�)>�ࢾ]�y�%Xd>P������T�f�G��1�wAu�4d�>�CL?��?�F�==f辷Ӕ��cf�G)?�=?/�M?b�?��=�1ھC�:�̾J��X�A�>)��<���$R��|����S:�|:	;�s>����K����;>�پ���Vt�1�]����	=� ���f=�"�o�־E���A�=�>(gʾ�,'�M���轩�Ec?WB=����Ba��' �oz�=�Pk>�p�>����63��.��P��bJ�=��>�dR>Η�r��LJH����>B�E?v�X?���?�d�r�x��)��;��񖶾'��mh?�>ͷ?� �>���=�>��?���f�OxO���>���>��M�>��R���D���$�w�>+	?�#>�?h�V?@�?�R?x�&?���>.�>d_������1?��}?m�=i�D<��j���_�I��"?��:?�#�@%�>��?�?܃?��c?��/?�$,>��Ҿ^�F��>�X>2vT��ȿBZk>�2@?~G>�ˁ?1P�?��>P7����sJ罍b���=�=e?]?W�5?�r�>���>&܁��2�=R�>ҽl?�ρ?K�?�z�=��?( y>�f�>މ:=��>� ?"�?hV?o��?�<C?�?ĵ<T��)���U�����üe=��=$�R=a���l�o,"�!K����<<�Ro�a(7����3���J����<�\�>��s>r��61>�ľZ]���A>Y���W���Ҋ�c�:�Ư�==��>??h��>�8#��˒=֍�>�'�>6��]/(?J�?�?��;߬b�&�ھ&�K��߰>�B?���=��l�K���-�u�h�g=��m?��^?x�W��*��B�b?�]?h��=���þ�b���6�O?7�
?�G���>��~?a�q?<��>��e�':n� ��
Db��j�6Ѷ=?r�>_X�(�d��?�>a�7?�N�>��b>&�=[u۾%�w��q���?��? �?���?C+*>n�n�R4࿛lþ�×���j?G�?����D?%��=%Z�K�d�>7۾f ʾ<����侅��b���`��9��P����N�=)�?�M?~�i?yA@?y|��c�R�d�V�j��Ih�I��L��+J�E�F�j~6��h�AM����z�׾.s�<�n���8@���?9v&?�x1�nX�>+阾�ﾆIϾ3�?>�Ҡ�S��y�=|�����A=��B=wj��5�����"?��>��>$�;?��\���>�@�1�f'5�����%/>�)�>PE�>C�>t�;��,�I��!о��̢��]t>]�i?"nD?��z?�-#=g7Ѿ_z�U�=�?s�<JsR��O��*h�2N�>[�5��D�<�r����Y낿�� ��hH�	B�Y,a�mRT?|}�>���)�?��J?������+�R������*>	 ;?��?��?>|����3�u��>��l?���>W��>�����I!���{��_˽���>�ۭ>г�>��o>��,�6$\�n��=���k!9����=/�h?�}���`�`�>�
R?+u:V�G<�n�>��v�A�!�U��e�'�3�>M�?=��;>�hž��;�{��A���6?��?+M����,�ep�>4�>�=�	?Oy�?��>���؀ ?�O?CZ?�x8?��Z?B��>�b2>� s�<��/fK�P{?=�-�>��r>���=�H=������ҽU������%)>��=��;��>@-�M�Ӽ_x�@<R> �տD�=��V�����e�1��H���1�ý|1��V���ǾBe���4�a@�\���Th�#[������|�wr�?���?�c�V@�!甿�]��O��k��>U�̾�+���C��`1P��c��վ����?%�r�h�0s��x�~5?B��S�ؿۨ�m�ƾ͒G?v�?e^�?���v�l�'�\�L	�= ߧ=BK�<mzž:钿
Cؿ�U���;?݌�>$w ��w����>lz�>�S�>��q>>��C��a�>U�?��^?�[�>���S�ڿ�ּ��>��?c@@RyA?��(���쾙W=���>[�	?&@>�O1��N�o󰾬W�>]4�?���?��N=�W��	��|e?��;��F��ݻx�=(�=��=���nYJ>�e�>}k��yA��-ܽ��4>�܅>>�"����L�^���<L�]>6�ս�T��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��=����Ҿ���	�f���9^���k�����'�q-�P:��q����$P�ꫝ=
��=�sA>.Ƙ>m)>qrx>��W?��z?>��>��N>䆪�t���)ھvV9?-¾r��;�����o,����>�Ͼ�^�e�-��z)�>k���/�m9=q�G�oԆ��V?�.-q��F���-?jk=�]̾'�M��a��-�������G�<r�ｧv�E�����/�?�;*?*Ι��b�
S��K�< W��ހv?`ώ�I��ے����<����9Ee<�>�u�=�!�&����b���4?0� ?rȻ�4����x>,��s'��S�7?��?q�<W]s>M8M?�e\���(����>��>Q��>��>]'>x���{����u?�yU?�{4�XYy�B��>{�쾃�K�z��xe@>�~��o{���b>�u	=\!��*������w=�[?BP�>k�%�=$�0z���p���$��ك?N�?���>;C]?[Q?�Ȑ=	�۾�.<�������=x�\?��Z?�t�=���\���ٶ���}9?��_?�0>Xs�x��h
7�.��c�-?�Is?9�?���4z�n ���;
��.?�'u?�_^�P��<��{(��,�>�/�>W��>9��i�>��;?��'�(������3l;�,�?���?���?��==0g��^*>�z?k��>�g���Ѿ��罂W���r�=*\?4�ξOr�r�.��G$�L5?j�~?"�?f�������>a��\��?Z��?���=����j����t˽��0=V3��`G����@�9���^����>O׻l>|�@��P@�>�$�T�ֿ�]п��y�:��W�>�>c ?æf>NH��'h���u���v��<I�K�F�n�m�xG�>�
>ӑ��mf�����^+>�ax���>*2>��Ƃ>12\������*���:<��>�%�>��w>�`ڽ?�ʾ�Ӛ?@�����п�I��	\��X?2��?�χ?߬?L��_Fp�j�������2C?��s?q�Y?K�:�O�R�uх���n?s��EXq�}�G�7BK�6K�>�+?.V�>��,���V=�1�>�i?퓈=wK�����N����� �?��?�޾���>}��?p-?mE�����ݩ�"{.�Aw����?�ú�����"a�wRY������F?�xp?��<�q�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?Z$�>��?�o�=�a�>�d�=.�-�+k#>^"�=��>��?��M?�K�><W�=��8�}/�8[F��GR�:$�6�C�$�>u�a?�L?UKb>����2��!�yuͽ�c1�7M��W@���,���߽�(5>��=>F>��D��Ӿ��?TI���ؿޕ����'�S�5?�>??��|��;l`?��>R��,��qk��~���%�?�$�?��?vؾk�P���>�]�>��{>~uҽb���B���=�I>�{??Z�� ���B1r�y��>�#�?P@�P�?�Tf�"	?: ��P��Va~���J7����=��7?�0���z>���>�=ov������s�{��>SB�?�{�?��>�l?P�o�+�B�%�1=XJ�>��k?�r?��o��󾅹B>3�?Ʋ�t���L�mf?��
@gu@��^?!�tۿtާ�S���ͫ����=I�=�8v>�8�E>�T�<������!>獬>4�>Q֏>�XK>��">��I>�=�����J���Ԉ�#$O���$�l�߾Z�U/���,�`	���澜��o��J@��˘�\�4����닸��|>eXU?��??��?u!?�YT�q9�>#�����g�齷�>[�>�{,?p�q?fi,?>��=jn^�7�o�����*H�����1Ϧ>���>�؃>��c>(k�>2�g=��=�bF>�Z�>N,>�vܼ(�u=��Ҽ<�>I��>���>���>��>�E=\���\���������������|Z�?'���?���}�Y�:�����C=/m7?2��=:,���ǿ�Sǿ�N?�S��CC�ޠ����>M�b?<�N?[S>u�W�;~�jz�>�dA�`&����>l�׽X����4����>�;"?�f>�u>˛3�Ve8�X�P��|��sj|>�36?�鶾*D9���u���H�scݾ�HM>�ľ>�D��k�}����vi� �{=Px:?�?7���ⰾ��u�kC��9PR>}:\>=W=wi�=|XM>jac�&�ƽWH��g.=/��=��^>U?q&,>(N�=U£>u?��[fP��~�>��B>y,>�@?�'%?5�����������-�5Nw>X�>#�>[A>�eJ���=d�> �a>��9�������?��mW>�>~��N_��Gs��qz=M���f��=���=�� �d�<��}%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ"j�>l|�6[����� �u���#=���>39H?;V��)�O���=�w
?S?�]򾤩����ȿ&}v�k��>3�?���?s�m�#@��W@���>���?�fY?�fi>�g۾VZ�扌>ȼ@?_R?��><�ȏ'���?�߶?s��?��+>`�?&^�?��:>�Eg�}|����F
����۾k}�=��Y>m��<��*�AQ?�����Ñ��R���q+��O�>���<��>�{�U^��e�%��I�C���ՕY��Ө>H�j>1:H>�R�>�B�>�ʏ> ��>p�D>���<K0��Ѫ����K??��?7��<!m�jl�<ڙ=�g\��?v�3?K3X���Ͼ� �>��\?��?c[?e��>C��WH���俿�4��֙�<��J>F��>���>'ď��N>]�ӾS�G��J�>h[�>4¤��ھkǀ��ӻ��/�>ς!?hJ�>���=ڙ ?��#?��j>�(�>BaE��9��Y�E����>բ�>�H?�~?��?�Թ��Z3�����桿��[�n;N>��x?V?sʕ>b�������TkE�3BI�@���]��?�tg?jS�/?;2�?�??_�A?~)f>Շ�'ؾn�����>��!?���A��M&���;~?�P?��>t9����ս�Dּ������1 ?�(\?�A&?М�4,a�(�¾2:�<r�"���U�m�;ىD��>�>8������=�>�ذ=3Om��F6�4�f<�i�=��>�=2.7��u��d�+?�8��Xy�w�>=�����B��ej>K P>,a��|	r?&IL�8�o�;��Ͷ��󓂾�2�?G~�?.ݛ?��7�V�l�
N?)~?+�?e��>����Q�Ծ�_�Z^Q��P����"�/��=#-�>���w�þ�!��H/��}ˋ�N���g,���?�W�>S��>�?�/>�޿>Ӯz�aY��ʾ0Ҳ�eO�G")��]h���5�����܌�ٽjM������{�!��>�W�;#��>(	?A�>_��>7>�>���<$��>m<d>`��>���>�F>��	>��={V"=J���KR?�����'���Z����2B?�pd?�1�>�	i����(��M�?Ɔ�?:s�?�>v>~h�J,+�qn?�>�>���1q
?�T:=��"A�<nU��Ѻ�%9�������>~<׽� :��M��mf��j
?/?�����̾Q9׽�y���}l=$]�?~-?	l�oZ+��Gv��qX�F�W�UQ �a����徾;�,�X#h�:W��r􍿍����'�f��=S�?���?Vl�oT ���x�s�]�L��:%>eg�>���>QH�>�|%>�����)��Ek�L(�xo���h�>�yu?J	�>ҫM?O�?S-L?���?2&�>�t�>���6?B?�S�:��>��?�5?�=?EfM?	!?�S?��>���=_Z����
?~�?���>���>�/?Y�ʾ�(���U�=T��<���r��ޛF=��������^>��h=W�R>�X?O����8�`����k>�7?V�>���>���,��R�<��>�
?�E�>< �i}r��b��V�>`��?� ��=�)>���=|���l�Һ�Z�=k�����=�9���x;�@v<j��=E��=�"t��D����:��;!m�<et�>[�?0��>�C�>�?�� � ����*f�=Y>�S>�>�Eپ�}���$��w�g��\y>�w�?�z�?��f=��=ǖ�=p|���T�����������<�?J#?�WT?n��?D�=?�j#?��>�*�2M���^��g��T�?w!,?��>�����ʾ��ԉ3�۝?i[?�<a����;)�ݐ¾��Խӱ>�[/�i/~����=D��텻���[��5��?�?TA�W�6��x�ۿ���[��{�C?"�>Y�>��>U�)��g�s%��1;>���>lR?�>�O?(?{?��[?�BT>�n8�t*���ۙ���7�z">��??��?�?��x?^�>�Z>��)�b��b���K�&>�z-���2Z=�gZ>3u�>D�>k'�>�"�=��ǽ'���??�Q7�=SPc>8��>S��>L;�>�qw>�Ϫ<��T?q��>F�ɾOR����]���!�4��?�T�?��L?�=>! ��~)��4̾�1�>?��?��:?b�O��_�=��>�uC���!Ծ⓸>�<�>��>%�>�iB��)>MD�>1��>��3��;�ٲF�%�����?�4E?L�D>�ƿK�q���p��ȗ�y�b<����d�K۔�[� ��=ܻ��J������"�[��������f굾h�����{����>���=_��=��=�<R�ʼ�<�*K=af�<E�=�Ap���m<�y8��rлy����Y���X<�H=�z���˾��}?M;I?��+?��C?y�y>�;>L�3�י�>����@?�V>�P�����ׇ;�<���a ����ؾ�w׾�c�;ʟ�WI>\I���>93>�I�=�M�<j�=Xs=�Ŏ=��Q�%=�)�=�O�=\f�=<��=N�>�T>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�B7>7>�R��Z1��[��b�ڵY���!?Z#;��˾c��>+;�=�|߾�Ǿ/�*=k,6>�cb=���\��=��{��==�n=R�>D>糧=�m�����=�oJ=n��=�P>?�;���1�w�+���2=.�=-�b>��%>J��>�h?��?�Q�?�Z�>�׾�'Y����?%?>��">ߨ�>�y�=�W>D?q�??�3?�H?�Qh>L������>��>�� �QAv���
��$������ӌ?]�?�&�>�o�����<�-��b��S	=��!?s�
?� ?�!�>ca�n>�
��/�Q�v��]�)�b>g�~��=�	x=�}��Z�����=ӹ�>���>��>Av�>��E>�g�>|�>�>0>�s�=��(=��Ʒ�<��+��uo=�j!=-��<|6 ��ݒ����<����Z폽�1�.H<phE<�}��q<�=~��>9�S=绝>:T�۵z�"�1>ˊ��@}:���=�\�4F(��҇��m��05��]@���a>��>:�<ϒ��8$?��>�T>S.�?D!d?ľ@>P�����Qţ�Y���ٟL�ۙ(>��.��J7�+^a�m�h�"�Ⱦ���>�>0�>?�l>�,�!?��w=��a5���>|�����5�B<q��?������bi��(Ѻ�D?@F�����=` ~?\�I?��?ʋ�>u���ؾB<0>�H��>�=�� q��k���?l'?z��>���D��H̾M���޷>�@I�3�O���V�0���1ͷ�6��>������оm$3��g��������B��Lr�[��>&�O?��?]:b��W��KUO����^(���q?�|g?/�>�J?�@?&��z�r���v�=�n?̳�?T=�?w>0�=B���W�>!5	?�Ζ?>��?z�s?��?��8�>$�;�� >v혽4f�=�4>�-�=d�=w�?��
?�
?�����
�H�ﾸv�H8^�7�=	r�=�>���>NDs>���=r�a=&e�=c�\>R�>;��>>�d>݂�>�9�>�<���9�ϰ?�K>03�>xTO?�u�>��H<%V���J�7n�=��ڽ�1���"��H��ɨ��;��>��<`��>��ڿ�f�?ꪝ>k��>?a�žځV�l�>�N�vTG��'�>�1>e�>�j�>���=S��=�}>7�+>4DӾI}>����e!��,C���R���Ѿc�z>���&�����~��zBI�Zm��=f��
j��.���<=�ܖ�<�G�?ι����k���)�����x�?�[�>�6?�ٌ�����>#��>�Ǎ>�H�������ȍ��i���?���?�;c>��>V�W?&�?ޒ1��3�vZ�4�u�u(A�,e�J�`��፿�����
������_?��x?�xA?�S�<�9z>Z��?��%�Lӏ��)�>�/�?';��?<=d+�>�)��l�`���Ӿ2�þ�7�pHF>W�o?%%�?WY? TV���Z�#�8>;;?o?1?�{?>5?�}L?���3J,?6�m>��>6��>��7?�2?�F?� l>Jd>�h<�8�=�뒽g<���𾽕�ɽ���,~=��=����6	%��u�=�~�<]?e�(Ǽ�<�",��g<�!=r}G=N��=`��>�]?^��>�>M�7?�m��d8�:ë�q/?J�E=ݕ���|���Ԡ�f��8a>��k?�ͫ?�Z?JXd>H8B�2B�+4>!��>9�'>��]>��>�u��E��
�=�[>k>�ƪ=k�H�&��8�	��֑�n��<j�>�s�>�C~>�����y.>�=��P}��Ti>I	R��ӻ��R�>iG�W2�׎s����>�
L?'�?���=|0뾼Y��zne�aw(?�X;?�M?\�~?��=��־n8��aL�.\����>|U�<�p	��{��
ࡿ�:��6�;�4s>C0�����ɶ�=�>������W~�V!g���v��
]�=x*پO�z��Q3���p>�)>�|��[-�%ٖ�D�܁K?:��=
F��'�,��%¾��>�b>b�>:M�<v�ȼ4f1������"<~��>e��=�νz�ᾷF�d6�T��>P�E?��^?s��?����
�r�W�A����p���Ƿ��(?^�>�w?=.=>�X�=��������f��)E����>���>����|G�ᾡ���o#�J>�?*�">?H�S?��?�a?�)?�Y?�$�>���w���+&?�~�?n��=�uֽf�R��8��[F�2��>ԕ)? 1E�d��>{�? �?b�&?[�Q?4?Q>!B ���?�9o�>���>�W�@��əa>N8J?�ܲ>�5Y?���?m�=>��5����r$�����=-H>�2?h1#??r?3Ѹ>���>謡�a�=ɞ�>Cc?�0�?�o?���=��?>:2>���>Y��=��>c��>�?�WO?��s?j�J?Ԑ�>B��<�;���6��"Hs���O�/҂;dhH<��y=5��1t��C�D��<�;e`���E��R��0�D�����)��;�\�>��s>�����0>�ľ D����@>س��oO��a܊���:�辷=�{�>�?A��>zN#�{��=X��>�A�>����5(?�??�� ;��b�I۾��K�S�>��A?W��=!�l�ǂ��}�u���g=��m?Չ^?^�W�#����h?��\?�����;�
����)�[���4�?]��>|����j>b}�?8]�?}�-?>4��Gr���7���%9�-�l��d�=��[>xL+� Xf�?�>4�5?���>�ߏ>c�$>)㼾`����}��� ?�?���?͒?�&R>}�i����h$��ي�XX?�͸>�ʾ��/?-�:�!ξ[Ӄ�OϞ�4˾��ľ� Ͼ6���Ր��O�ڽ�V��zc�}M;=�?�k?-�?�j?�UV��Yq���{��EH�����e���S�-�G��<��^�%��Nݾ��n�y� =����m�A��2�?�&?
q4�M,�>r(���n�6iξ*�A>y����j��C�=�A��{J=��[=ңj���.�0{��0!?`��>d��>'5<?J�[��=��2�N�5�\����11>>�>��>�#�>o��;�-����ʭʾ)j��-�t4v>?zc?U�K?�n?�b��%1�������!�R�/�tc���B>�x>Xĉ>�W�S���;&�XX>���r� ���t����	�N=�2?I�>[��>~M�?|?x	�8i��BKx��1���<�:�>�i?�1�>݆>� н�� �,ŵ>��p?4��>�~�>��^�ve&�B1j�.az����>��>�Q?��,>���e�f��䚿����������"pF?Zn���!�i�>ƞD?��'�Q&P��f�>]7ٽ��Q�-UӾw��� 9>�.?��>ҕ�=@��I>�ml���'1��A)?n�?zԓ��*�D��>�x!?�!�>�̤>p�?ј�>��ž�a;�?|�]?<aI?�@?1�>�*=;O��Go˽��#���-= B�>I�Y>(�k=���=��+�\��.���S=ii�=y=ݼ;ƽ�Ԃ;��'��<��<,�6>?�0�L��"�����Vq��T��k��;� �Qܨ�I.��ߢ�Jx��(���ĽS$0<�G���s�������g�(:�?&��?� Y�|�l�����������\�>?G�#�����q�սr怾�f��D��~�	��GK��fa�l�j�K�'?�����ǿ��:ܾ-! ?�A ?0�y?��-�"���8�*� >wB�<�,����뾫����οM�����^?���>��/��q��>ू>�X>�Hq>����螾2�<��?3�-?���>�r�0�ɿ^����¤<���?/�@�|A?��(� ��cV=���>"�	?B�?>�J1��E� ����H�>�<�?���?��M=��W��	�eze?�� <r�F���޻�$�=P�=��=����J>�P�>���ZA�Mܽ5�4>�߅>UW"�}��d�^��g�<��]>��ս.���/�?}�e�e�p�#7G��Hw�\�>�nr?��>z��=��1?��c������Z|�8�2?&�@hk�?�-?�����>���!z?�::?��4>�A?�9O������S��>�����sK�W;�=�|�><F�>D�˽1�'����"7�=�s�����ÿ������X{<��'�����!$�"����0�t��O��,���i�=&�>�=>��p>۠O>�MT>^>Z?��n?�>K�>	��#m�����4������舂�g��̆���־�g˾���)�����þ�6=��q�=GR�]���$� ���b�J�F���.?#$>��ʾ�M�u�0<eGʾЗ��_���Cĥ�7?̾$�1�&n�Bϟ?��A?)셿��V�������%����W?�)���̬�}��=�岼j|=��>Kx�=���((3�4�S��g0?��??�ɾ���>X>s�̽�as=�#)?,.�>��	=��>e}+?��J��U����J>�$>��>g��>Q�=,C���B��jl?%�X?�=��Œ����>�z׾�����=��.>T+�_���2%>a�U�S�)E<S�5�P=�(W?���>��)����a��8��kX==ڲx?��?�-�>w{k?��B?�Ӥ<�g����S���'^w=��W?-*i?�>����	о偧�<�5?֣e?��N>4ah���c�.�yU��$?G�n?o_?*|��w}����L���n6?Y�?������(�
��A����>P?�L�>9E#��	�>ˋE?�B3�I쉿	����>��ڙ?ds@��?q�<��	<Ƕ�=��>G� ?�ju�q�ݾ�&�aꢾ�[��yO?���u���I	���콰=?xw�?ɨ?vL޾-!𾇠�=Zٕ��Z�?_�?؄��ATg<)���l��n���v�<tϫ=9�M"�����7�/�ƾV�
�����t俼ץ�>%Z@@R��*�>�C8�*6��SϿ��h\оUq�B�?;��>��Ƚ������j�/Pu�<�G���H�M����ʢ>H�>U��������j}��C;���<����>'���:h�>�aY� ���N��j#�8P��>�%�>%��>�����`���Ś?T�����Ͽ����D��_?�ݠ?��?��?���8�-h���f�)ɓ;lF?W�r?L�Z?��PM�-aY�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�O�p���-���ƽ�ۡ>��0��e\�>N�����Xe����@y����?N^�?i�?е�� #�g6%?�>b����8Ǿ��<���>�(�>*N>QH_���u>����:�i	>���?�~�?Rj?���� ����U>	�}?) �>с?u�[=��?�N�>���4�=f�=]�>����8�>�}t?_��>q�*>�BK��I-�dD5��:X�� ���<�Ex�>Q�z?�6k?�\�=?�ż������%�y�V��塾x��>w��q�}>�i�;��1>�/>z#�=&(�����Z?3r���ؿ�����*'�~5?}�>|7?���t�7ջdq_?�B�>���������nP��j�?���?'E	?�Tپ��cU>��>�I�>��׽�Z��E ���$3>8�B?�"�
E���so��{�>���?��@���?a�i�ۊ?�.��)��8���t4�0_?=k��>��?mV̾3}>"6?/5>��O�Z���v����>厩?�)�?v	?[�v?7����f�;V<>̹?Q�?���>B(�+���H��D�?�Ԕ��b�����5�E?�;@��@��m?)��EO�����|���5Y�����=���=�> �4�w=Ǩ�=ta�<�G%=a!$>S&{>h[,>�j$>&�>o/Y>yJ�=�����!�C|���<���5�t�4���_������ԃ�&���z�}Ծ�ҽ�B�63��e��7�Q��W��[��=��^?z+X?P�?��?a�6=fVJ>x��P�=L(i��;>���>��N?�~Y?:�?�ޒ��A���sX��nu����!�n�T�>ф�>rļ>�f�>g˜>��=��~>���=�"�>*��<��=2�=��}=��>T��>�v�>�i�>{C<>��>@ϴ��1��g�h��
w��̽*�?~���H�J��1���9��զ���h�=Bb.?�{>���?пc����2H?&���s)���+���>x�0?�cW?�>���T�;:>*����j�`>�+ �gl���)��%Q>}l?��f>\Rz>��4�VS7�qL�b���!�>��2?�:��
�0���u�E�E��ྵ�G>�>�]����'	��%~�{Yj�}uk=9?]�?�Cƽ�����u��N��[P>�Y>q�J=���=)�N>��_��Tǽ��@�E�M=���=)zh>-A?�+>G8�=4��>9x��,qO�3��>�<B>Z�+>�??~	%?	��[���c~���-��w>r8�>�>��>�J�e�=���>�Lb> �8��}Z���?��}W>V��}�^�lv�gw=����9A�=�(�=k ��<�xH&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�Y�>z��ٌ��}�����×1=���>�hD?D�����>��R�O��>.?=e�ju��Ȳ�24Z��8�>x�?�!�?\��z���'V�K�> �?UVz?ΠH>�ZѾ�¾h��>�p?�nQ?Hܬ>e���V��z!?��?��H?�:A>�:�?�o?�3�>F�]�F0��"���(��1���]�n;Oh�>��={8���F��Ǘ�����se�l`'��\>�j=� �>�d½!���	�J=����l���W���ף>>s�>G�i>�y�>)��>GH�>Z��>Qۼ����5y���h�0KO?D��?�-�dT��/q>ص=>����L?��<?�v=����&�>ԏ??�?h�C?��=*%%��n��I!��:�������N�>N\�>lN�>(t�kIc>`x6��.����>ς>e�ż�� �kq�g�����>a�7?�Q>�л=<�?��0?_�p>1E�>H�G�E����#�m��>��>?���?E�!?ڋվ)��+���0���,Sk�vFs=�~�?n�.?g&0>N9���(��Ei����=�:��B�?{st?M7����>Y��?�#7?t�v?�Ԉ>�oW��;��	h>b^Q>T}?�g�#C�Ђ&�c<�bA?��?�y�>-̱�
�˽5���N�����
?aR\?�%?+��XI^�#�ľ���<����8:�i��_��c�>��>�$L�8��=1�>���=J�l���,�ej�<A��=�d�>:F�=a0���c���,?��e�C���x��=Ss�S1C�{ǁ>7L>����?^?z8B���{�V����w���uK���?�%�?�]�?BU���h��x>?봇?�!?��>������ྖe�7^z�m�w����^>���>#���%�䤿�l��fL��fϽ	��N ?���=�p�>�^?���>��>�����Ka�������L�U�Oi*�?�R���e���얋��72��UL�-�¾{$5��$}>P�!�.�&>���>�2�>K�>N��>��
<��9>:�=/��>���>�|�>��Q>I>Eb�=����ZR?S��
(�o�辊���}B?7Md?)��>��d��v���(�<�?鎒?�?Ifv>�|h��n+�^�? �>g%��C
?vw;=����ʓ<�ƶ�S9�L���\
�魏>�'ڽ!:��"M�׊f���
??v?����E;�ٽl���r�)My?�S?݅.��ej��]�kOL�<�G�ј'>Oj@���v�)>C�F`����ʀ��ꃿ5a6�w�D>��?}�K?W��e̾]VZ��`E���־t�>7ѽ>R6�>E�>�d8=:F!��F���e�Z��X����?���?,�>1J?�;?r+R?�eL?vy�>>�!���j�>�;�)�>���>{�;?��.?�.?�?��(?�^>�\���d�� �־�K??�?<�?�|?B�?�������
��8yȻ)V~��.n�m��=���<��ڽ��t��f=d!Q>DY?��g�8�C����"k>�7?c��>���>���A!�����<��>�
?�G�>����{r�sa�`;�>���?�5���=U�)>03�=Y�����к�F�=�9ü���=ψ����:�!<3��="��=��y�jr����:f�;��<���>�S%?j�>U;�>r~O�j�_��<�>�>��Q>��	>����R���\���r�ɧ�>�ޔ?��?"��<*G~=���=ݨ���)��� 1ܾ��_>���>�>�LK?��?��D?Q?Y�<�6+����-���h��?� ,?_��>���B�ʾ�憎W�3�q�?�Z?{:a���<)���¾�ս �>t[/��.~����3D�B=��E���|����?���?�A���6��v������\����C?p#�>nY�>	�>��)���g�r$�6;>��>�R?� �>W�O?�={?��[?QqT>�8�L,���Й�\C2���!>�@?I��?��?�y?cq�>2�>��)��ྙT�����"�iӂ�y2W=Z>��>�$�>h�>��=!Ƚ�@��n?��Z�=��b>{��>噥>�>?�w>#Z�< 4G?���>�U��S>�K鞾0���!m��^u?J~�?��'?8.�<��;MD�Z������>Î�?�+�?FI*?TRQ��t�=��Լ絾i�7��>��>	9�>��=sQ=v�%>I��>�Z�>���Ku��'9�`rU�~�?�pE?�m�=�x����]�p(=�@�$ɾ�)��D�i�`�R�����=��^����<�tB�t��=!�&�	����	�������q?�>��=��K=u�s�|��t�c=��=qD=��ļڒ޽$+����$�Tސ�G|��iɼ�J=�r˾Z�}?
6I?�+?h�C?|�y>�f>� 4����>}΂��F?�HV>j;O�hX��Sf;������$����ؾ�׾ld�����!g>y�H��>�3>{f�=�Љ<{�=n4s=7Ў=��a�q�=^.�=�I�=�9�=�<�=	>pP>��?[��x���%O�����D?�h�>э�:���:U?$6H>!���:��rv�Zj?�P�?�^�?�: ?ή6�+�n>	ܨ��<y/�<+�b��d���++>R>��>��>��G�����y&=�1�?ߞ
@e�Q?�6��o�ɿ�H�>�}2>�>��T��<1� �U�g;T���B��D?�o>���ž�s>���=���5˾h=xI7>�Sd=T��̌[��ߍ=����l�L=*Z$=,lv>��<>"��=�o~��=%U=N�=�4H>���;y�Լ�`���b=���=��f>484>,l�>?�>1?vY?W�>hq�+�ݾ�z���>w+=t��>���<:JY>��>��:?H�I?�O?̸>�ь=�2�>�%�>��-�gk�n�Ⱦٮ���[s��x�?�Y�?�F�>@�ջ�t!��Z�z�;��ө���?�.1?��?M�>�����ݿ����'��ϑ�8���<у��ٓ�0`��jF�6#���@�=�?�>Z��>B��>�E>�E)>+�4>iڹ>�_?>�-a=Z�=��L��Ę�:���3Q<I���>�;vq"���عd�<���W�=+��<y�<s*���<���=,��>�)�=��>�=����Y0>N��{h[�ɸ�=����Ϳ=��Lg�B䁿��%�j�(�>�%>X:(>@鴽8���M?x�%>�V>��?�5l?G#>�l2����=Ú�3um��V4�\�=y4=��k��?� [���I�26㾒��> ێ>��>�l>�,��$?�k�w=���a5���>}��=���:�:q��@��~���'i�vAԺ��D?0E��z��=_"~?��I?��?���>Y����ؾ*:0>�B����=��M+q������?'?I��>���D���Ӿ�im�n�?��R��J�ﬢ�����ν�Q���f#?�ؾ���ҚI������6��8��~�gS�>i��?�&�?jJ���Tq��l�������=c�6?�o?�x�>��?���>��E�k�������BX>I�t?�
�?#J�?���>Q��=h�����>�?=n�?ˊ�?B�s?0�@�h��>���;�y>�ٜ�[�=��	>M=�=, �=�A?�Z
?g2
?e���O�	�)
���ߝ`��x�<�s�=���>K�>m�r>�i�=�$e=���=aQ^>4�>q�>�e>�>`0�>e��i���>�Ƚ��=! 6?7��>���<]���C=�E��n���/=����Y�<�)�=�'_=ժ=�=����>n�ƿ˨�?�4>����'?*��9��<��>8~t=S؅=�4�>h�>�=�>'k;>e�>�L&>m�>?�*>���]��=NT������rL�$�_��:�0D>����N��7�����d��룾'n�sf��F��m�D��Z�;��?���al\�kP"��򍽻�?�)�>�g%?Iш��p�<�	>��>�2>r�������3��K�Ͼ��?�:�?�Vk>!�>Kg?\��>:�s�p2L���W�foc��	7��x��]�C�����]�(��Gz==p?�bl?�CI?'^����|>���?4��������?6�L���i�.z�=��>����ޭ�Meپԁ;�=]����>�o?L�{?q��>�?����2�A��>�eT?[��?*�v?8H,?�3?��f���?�>=��~?��? �s?#(m?�~�>�)���I=���=�� ��Ń��p��������.�}�W=1����=�$��E}����#>��=s��"姽yO���<Vc=p�=ѱ�=d�>��>�g?i*�>g�=)}h?�xc������(s�?��b8 �����Ƚ0��D�>���?ิ?/rT?a�l>u�6� Ͻ|�<���>�=L�9>9�h>I��="�&���>gs>��i>O�+��C���>�/���q��A�-=݋\=���>��T>�&����<&���d5�o�>+|��~����5׽hwD���3�;���9�>V?A�!?��=rZ�������s�1L?Z�?��W?� �?�$>�&���e�%�{��O5��$�>n�=�۾e㲿Ʈ��x`�*�)�I$<��ھ>����u>i������}�Sv�Q���N�����#/>CI���n���p��mE>3>u���@:�*Ğ�1⶿��G?: >����y��p:���:=��>'��>�����f:=P|G��V��;J¼��D>��=�4��re���VB��7���:�>XE?2Y_?}m�?����s�J�B�����&v��!�Ƽ�?Us�>�W?@�A>�l�=���� ���d��G���>P��>���\�G��>��x;����$����>�B?N�>k�?��R?�
?U�`?�*?><?D�>�Ʒ�Hϸ��8&?�w�?�z�=0�ս �T�9��IF�`�>e�)?�0D�y;�>�?>�?�&?�XQ?��?�>o\ �I@���>�W�>��W�{Q��L}`>�zJ?U&�>GDY?�?�d>>ކ5��l��rn��4��=��>��2?	4#?V�?:��>f��>w���_A�=��>Nc?�/�?�o?��=��?xA2>0��>�=��>Í�>�?oNO?��s?��J?F��>�Ս<�0���L��is�yP����;)\H<�y=n,��/t��f���<�t�;u���%���u�q�D�b򐼿��;�V�>��s>�ꕾ+�0>m�ľ�$����@>r����Y���֊�/r:����=Jc�>�?崙>5,#�ے=���>�-�>8��O7(?��?a?��;��b��3۾/�K���>��A?J �=��l��v���u�5!g=P�m?ʅ^?�aW�-
��
�h?Q\h?#�	�|�:�"���j]�wc�ϝ�?�a ?T��n��>��?�6�?]�?����׆�d���~�9��v�'�>5��>�!5�]Ƃ�k��>!O?4��>�ޙ>�<����X������\?���?^��?U��?�Y�=�s�O�⿂������I`?�|�>"Ҧ�$p*?7"S�;a߾kꊾ�G��Y�ƾ:C��}��3a��\�����iE[��j�v1�=c?Go?�Dr?l\?eB�nhb�|�v�5u��G�;����"��"V���1��CC��Nq� ?��پ�tv���=�2x�f�@��ϴ?�|#?ɰ1����>�햾���̾ɓ=>-�������>=��9�4�S=Z�=3�X�"�/�cH���?�[�>.�>�<?�]���=�kK;�g,5��a�\�>P��>U�>؍�>W��E�=�k�������t�ò��5v>yc?��K?�n?�j��&1�C�����!�+�/�b����B>�k>��>2�W�x���8&��Y>�[�r�����x����	��~=�2?�'�>e��>�O�?�?~y	��e��gx�-�1��h�<�2�> i??�>v�>н�� ����>��o?��>=y�>�u��c"�+�~�t�|�ZO�>�N�>&k?*�6>3���Te�����V����'���=�bP?�Չ�z�Խsc�>)R?�4;��y`���>�N�.A�mW���U��\l>�?�s=	ì=Hf	���1�$4��z����U)?[?/,��>�*���~>�"?��>�>�-�?���>Z�þDfĹɍ?��^?�J?�$A?�>,l=.Ӳ�^qȽb�&�-=��>6[>zn=	�=�h��;\��4��uG=���=M�ϼ'�����<-��+HX<	��<84>j翟�G����w���x��a�%��Q�2�8��Zн$q�9�o�1h����;��|Qh��x�L����k��=#�?1��?j�Ͻϗ��A��	������`4>#@1��b�=����̜�������N��pYf�89��X�Tq��7��Q�'?s����ǿ鰡��:ܾ2! ?�A ?7�y?��0�"���8�l� >�B�<�-����뾦�����οh�����^?~��>��P/�����>ܥ�>�X>�Hq>����螾1�<��?7�-?��>�r�*�ɿQ���EŤ<���?'�@}A?��(�/��JdV=E��>��	?/�?>�)1�e@�k��I�>=�?���?�M=+�W��-
��re?�� <��F��u���=!��=ݪ=N���J>Y�>V���UA��dܽ-�4> ܅>"l!����'�^��}�<
�]>!pս���o�?�oz��\i��de��Z����B>`�J?�zP>Vt>��*?�}���ӽ�<y���C?V@{h�?�8?�vξX�?�W۾��z?�K?Pd�>_�@���B�g�&>"u	>K�=��龬=��L>|
�>��>�\���)F��k���<lV��x��&ƿ�,��$����=�	����V�Ќ�Ɨ������a�܉ֽ%��=@��=IU@>_ހ>��G> _>��T?ޑt?ߒ�>�>��=��⧾+������|���нa����1�����Ͼ��ʾ�A�����`�;��=��ߍ=��Q�Xk���� ��=c���F�q�-?W�">�ɾJ6M�M�4<��Ⱦ�q��c����G���̾K�1�j�n�ꯟ?�xB?!t���	W����;��I ���W?�y���]������=񖥼�s=�>ed�=�㾂P3�L�S��g3?�#?���Nk�|4{>gf���c=��.?��>L��o�>��7?G��j^!�?�>��=!b�>�̝>?��='A��~K�rS%?��q?)�� d���>'�ݾ���y�:�>�.�� >�=<�3>Zfa��{�[3==��	=�Ǌ=y(W?���>��)���Xa��] ��U==��x?��?�-�>W{k?��B?�ͤ<Vh���S����bw=��W?�)i?:�>ކ��<	оހ�� �5?��e?��N>�ch�����.�U��$?�n?_?ց��aw}��������n6?��{?��u��T��D!��j��)�>�:�>{��>��*��3�>=]B?B��Lܖ�b>ÿ�7��?@�@���?��<��<Z�4;D&�>i��>��ɽA|��&���qپ�X���?�E���퀿��	��M����.?b��?U�?]���U�H��=xԕ��Y�?m�?փ���ng<���l��m���W�<5ޫ=�+��"������7�/�ƾ�
�����_������>�X@@8��,�>�I8�54�lSϿH��_о�\q���?�x�>]�ȽD�����j�Pu�q�G��H�͛��c�>R�
>mᏽ����=}�R�;��5��|��>��ʼ��>��W�z}��Q�����
;�>�>,��>��> �[���?ó���Ͽs����Z��\?=I�?���?H ?+
b;��o�*}t�?�a�E?�s?~sZ?>D��(Q��P�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.��_?Μa���p���-���ƽ�ۡ>��0�j\��C��N��3Ze����;Ky�9�?_�?�?���� #��8%?��>3���	3Ǿ���<�z�>~&�>�)N>"_�C�u>����:��k	>��?�~�?_l?m�������1U>��}?�m�>/�?F�~=d�?�'>Z��=�_=ʓ2>J�=�I��!?�i?)4?Ĭ�=��p�]))���/���=����=�훘>`	z?�=_?	�=pÓ���=��-�����˲D�~�Q> Hӽ��=�V�=ìY>�H>ڨ�=*s��<2v���?Np�9�ؿ j��!p'��54?0��>�?����t�����;_?Oz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>>�>�I�>E�Խ����]�����7>1�B?Z��D��t�o�x�>���?
�@�ծ?ji�q?��,�����Ѓ��C����>�4?�>Jw?`�*���{>���>S��=ӿ���]��t�Y�G��>I�?o,�?�?q��?�8���s���)>}k?zv�?
�?>� �v���>��.?#���u��^���1?v@��	@O�Z?�4��ʴۿ�U��3��� ���ey>h���=�H�c��<?�<i�=��}�,�>��>�/>oLQ>��}>�x=>;�M=x����G#�b��C݈��e׾����/��.��������gC�jZ����˾:ۑ����j�����#�$��ļ���=]0W?j�P?R�r?�u�>A�;���+>v����=�.�y/�=�L�>z�2?��K?w8(?��={��a:c�=�}�3ۨ�������>�G>�u�>�	�>��>\y(�LO>�D>\�>�=�=x	=5�<�<=y�H>;��>5�>{��>�B<>Œ>ϴ��1���h��
w�̽�?}����J��1���8��i���ti�=b.?{>���?пW���d2H??���)��+�>�>1�0?�cW?�>���c�T�:>�����j�P^>�+ ��~l�
�)��$Q>�l?��_>k1|>�|3��L5��'K��ۦ���>��/?$�¾�q'�@�t��!I����<J>��>)8[��	��<���4��QIg���G=��8?PV ?��p���?�g��e��Q�\>�Y>�Ls=i��=NQ>ٖ&�dé��X7�¤q=U�=�X>(P?�+>,�=�ˣ>6O��۸O�	~�>="B>�+>Q�??2*%?Lr��?���S��Q�-�'w>�E�>�>[>&?J��=Ӎ�>+ b>�d�߃��P���?��W>Y��(�_�mw�6�y=�,���8�=��=N �i�<���&=�~?��䈿h��k���lD?t+?���=��F<*�"�V ���H����?a�@`m�?�	�}�V���?�@�?���ν�="}�>�׫>�ξ��L���?�ƽ1Ȣ�ޔ	��%#�HS�?��?��/��ʋ�Sl��5>�^%? �Ӿ$h�>�x�NZ�������u�ֳ#=A��>�8H?�U��:�O��>��v
?�?6_�Ʃ��|�ȿ�{v�N��>X�?���?[�m��A��@�(��>o��?�gY?�pi>g۾:bZ�Ӌ�>�@?�R?�>U9���'���? ߶?y��?�>>73�?Huv?	�?��)�i6�-�w;{��+���S=>j�=|�ܾ��J�_�������`�/��P�>x�Z=��>ྉ��m��f�h=��-�M�x�[��<�5�>��>�(%>���>�?
n�>�p>V�m�|�齢sK�f��/T?@�?�P7���i�>-.:>��>��F?�o#?n������>��>�K?�M_?�<?ܡ�=�#(�.ܝ�N���(믾��ڼLv >V�?Q��>�b
;�z>^t%�5q����>Q�>���<�c#��N뾰��%�>�h>?�c�>��=$�?�l<?/5�>�m�>�u7�`̑���E�X� ?u]�>�o?��x?�(?ா��$�����P��N5Y���.>��?$#,?D�R>H;��s�����彞;!>��<���?1�v?n�˾>��>k2�?�j?�c?�^S>�#G���Vb=>m>?k�ͽ#�@� ��Dܽ�?U	?&_�>s�#���^��*����!����?��[?��$?��	�t�g�%�۾q��<£#�Bw�;;��� ����>��3>Q���Ƒ>��>H�>��=�ǰ��pv=�>@}�>в>J]��ɛ�9�+?��$��F���!�=�r��xD���{>fO>����5�]?��;��{��0���]���ZV�fz�?mp�?Lb�?�÷��Bh�g=?Nه?$�?J�>����ܾ��]�}�`�v��)��5>���>�҇�	�<)���򪿭����ؿ�"�i%?JM�>�_�>�-?�X�>���>�CվeW��蚾���/Ue��>�b�'�%�������Ѿ����4��ƾ�M`��q>�A���>��>m��>r�>>(�>�_�=�5�>��>(�A>�#�>BY�>�c>�q%>^� ��1�zXR?�E����'����ca���&B?�Bd?)�>��g�_�����S�?Ǌ�?�l�?Fv>�h��W+�}!?���>���KZ
?M�8=	f�m6�<
��43��:�� ��2�>�ؽK":�P2M��.g�ƃ
?ue?!����;�d׽qE˾{	=��{?
P?b�C�x�o���d��dY�^�Q�Yk�=�+��������	��x���g��`���0�\_>f�$?Yul?�xپ_ǻ�K�����V�,u*��.,>�u�>Y�>o�>�2>���3�I�B*f�Wh�E:�.2?g��? ͍>dIK?�2;?%�S?+vI?�e�>z�>2���_�>6��o��>{��>��:?-�-?�^-?�	?5?'?Y>Ͽ�U����7Ҿ��?�?	? ?�?紉��e��^5���ͻ�8{��ď���=��=��۽�x��b=�.U>�]?!B��8�S����Ck>j�7?�t�>���>����9�����<�5�>$�
?�%�>`����tr�q]�l�>B��?-e���=��)>{&�=G܅�|S����=ɢļS��=/���9��H"<��=z��=#���S`���;��;$b�<���>IF ?|��>"��>y�S�����)�n;�>Y&�>=�>y�>b� �w��L����]�z�s>ڻ�?��?V�j�>�a=�'>>�}�!,սS���U���>���>�|z>��F?�ږ?��Y?pA�>w�=�>�����쐿i�侉�?=!,?9��>���S�ʾ�񨿥�3���?R[?L<a�����;)��¾�Խg�>�[/�G/~����WD��򅻒��a�����?���?�A���6�2x�̿���[��2�C?W"�>�X�>��>p�)���g�>%�d2;>l��>�R?�#�>N�O?�;{?1�[?�fT>��8��/���ҙ�!,3��!>�@?���?��?�y?s�>i�>��)��ྛQ������
��݂�4W=.Z>H��>�+�>��>���=G�ǽT���>��X�=H�b>h��>���>� �>�w>�\�<��;?�=�>����¥��@��,;���D���Ur?2�?{s�>MW��F��y��R��׎>���?A֯?��=?�@��Ag�=PJ�<z�����b�h�>l{�>ѥM>��#>p/>�ԋ>*��>�)�>��A^��/����c�?��&?up�=Q�ǿ�Dr�E�}�Y×�[��<g���T�p�"����b����=���%L��-���Q�����n��'#���G����~� ��>+�=c�>P��=5�<���Yԗ;�N$=�$&<*�=W?x�Iۂ<]�S������N����K�MN;ñ$=��;ROƾ��y?��L?��.?�LE?c
�>�6>Q���˦�>	���?�Ji>'̩��
���R8��2������׾tԾ��c��訾�;>9$M���	>��6>�9�=��<�P�=HA�=%�=�0X���=6�=J��=��=�q�=�$
>�	>��?����Ҳ��{Z���#�$�>?�*�>\�U��(���V?	��=��~��Ĭ�$'�^�^?�@k�?�(�>{��=y��>ΪH���=�#��|����Ҽ��U��/��	�>�C>��P�W*��)A�=�?~.	@x�W?0`����ܿ'b�>�<7>��>D�R�D]0�:V�0[�YaT���?��;��ɾR�>ri�=���`ž?=��6>xNM=�� �l�\�}ϖ=�����E=V�t=Y�>�8C>@��=A~���d�=))E=��=��T>M����:)��.!���F=K�=9�f>[J%>H�>�?�t0?�Kb?���>أn���ѾA�����>�]�=ɮ>��Z=L@>�c�>P7?��D?.nL?�r�>�{=㎺>{	�>O,�s�l�����驾��0<���?�)�?���>��;�@�Y�S>�r�̽�?Hd1?(5?�>+��p�࿓�0��L'��
�<�<����o;��[�=��tς���/+ٽ���=��>e��>;�>��z>Hz4>�/M>���>��>�MH=���=���R�eؽ"��<�}����<P��1W�;�C&�nHW�O���E���UB��%8��=���=���>b�>j��>ì�=Q*����1>HU����P��w�=�����B��vf��G|���,��2��2>^=E>IC��֑�ls?VlQ>Ώ@>U��?,Eq?`�>�����ؾ�p��>Sl�Է_��ј=A!�=�?��@:�^�_�O�N���վ���>�>��>��l>R
,�  ?�v�w=i�se5���>^�����5��8q��>��y����i�l1غ�D?IF��$��=6~?h�I?1�?:��>����ؾ�40>�B��\�=��F3q�Zw����?d'?��>�쾻�D��O��K�s�>�O��e�n�m������&��<���?C�򾦎ɾca=��ᠿ����3-�AV���>�$�?J!�?s��M`�����۾}-�>��4?�o?��	?;�%>?�>!}��d��'�1�>�Ђ?� �?�w�?�>_��=�ഽ�(�>�'	?v��?��?�s?o�?�ZJ�>%{�;&� >�혽~��=�>�=N�=�e?p
?��
?dS����	�;�����^�A��<eۡ=���>���>Zr>���=Qah=���=b]\>/��>��>�e>��>�N�>p����0����?�O�<Oˊ>"�=?���>�Ӕ��|Y�x=�=�s�=i�Q�k��Î�=��=78>���;����7����>����U�?^��=�����? J$�?@���E�>8��<zȰ=ھ�>I��>��>�qI>~�>�>=S�>�k>U��>b�پH� ��pp��Z~��s����=F|;>p6=����h��(�A�ľ2�	�\Wb�������b�}����?{�[�*BF��߾���2��>���>98?4(��U�=.6=�)�> �j>�4�>��뇿�Z�����?)�?�m~>Oӄ>��`?���>򣾀�	���k���U�?�	�9_��9�K�����T�B!���2�4�e?}�s?�B?�����	v>��i?O���{�web>��v�ڶq��O�>���>iv�%�ž�u-��m�8�Ⱦ0�=6H?e]h?��*?��n�ht�P6+>+ h?�t?^�b?U�+?�zn?���&�U>&��=_�W?��.?Cf?��C?�Թ>l ��B��D�>�l�	����T��C�N���\�$=����K�N���j<#�;%>�e�����v���w=o��:�H�<uY=g��=�*�;�&�>\J?��>;?�=��"?Bր�u�l�a���Y�?l�O��a���F�����*+;��v?�8�?\�h?3_=��,�\H����=ޢ�>9�>�3k>;­>��<C�`�>~M>�p>_B�����y���&���E�?��uw=q��=�?��M>=l��P��<���iS�C��>�о*���e��5E�e�%�2������>�k?o#?�'λr>����<���y��R?�(?!+e?�ؕ?�N>��!�L��4��y�����>8�һ����V���D��ըM�q4H�Ze�=)��/6<���>4om�!���Ny�]�����'�����pe=�yȹ>��Ⱦ6X��S�S>O�>Rf>�ݲ��<�Ϧ������T??a��=�sE�|`�h���*੽r�T>�:>�����H=�:�#В��=���>o�O<�����a	���9�S���R�>S�I?�uV?���?6���[n��@8����^㐾���̞ ?ù�>�/�>�E>���QӾ�_�h�c�b>�w��>���>w����<���ž�����"�`]�>�?�O>LH?W�Z?# ?v�[?e�?>�>A��>�����~(?�?�]=���MQ�x�5�F5F�k?��+?3�L��@�>��?w�?+U&?|�S?��?��>�����?���>�(�>vZ��⯿��}>��K?���>�QY?�G�?�B>j�;�����`����R�=sF">�Q3?�f$?�#?VY�>�I�>硾ѭ�=���>�bd?���?��o?�I�=�)?�}3>��>���=:�>߀�>�?�M?��q?�J?���>�'�<�L��k����gj���'���;��}<��=F�ż�}�(�5���<]�H<��������{%�Q�K�z5�����;���>w�u>	�����4>��¾b7��0~C>m���Ǚ����uo=�r<�=�,�>�?g'�>��%��2�=���>D��>��C�(?u�?�}?�睺#b���پܘL�o��> A?~U�=7�m�|���}t�DZo=2�m?��]?��Y�����яp?&xY?@��B�,��q��:C�#/��\�?>�??l�L�j�>�bl?zd?}�	?����\��(���wp�	�a���I>��>}�3��ٌ�Ǳ�>��K?8�>� ?RV<�n߾mN��w�M��?S$n?Q+�?�y�?��8>"�F�K޿����g��v�a?h��>~L��bU#?�����Ѿ�۔��E���r޾<���P���ꌆ�W��e���d��ᏽ��=��?��t?��q?+�b?��c�e���\��F��)�Y�*a
�����P�1@��z=��[�;����W�խ���IN=m����@�D��?3�?ԆJ��"�>鳣�-�����Ծ	�D>����?i���=��&�
�t=5G�=2�M�r������q"?4��>8��>��=?�G[���?��i0���9����K�>�S�>�'{>���>�h�<�D��ܐ��Jƾ�0��Խ��u>ޓc?hK?��n?Bh��1�\e���q!�hv1����8�C>��
>Ԍ�>�WW����,k&��f>�P�r�7��,(����	���=W�2?��>��>�=�?�?�	��x��&0w��	1�@3�<��>��h?�v�>���>��ӽ�� ����>��z?8��>	��>vE�W#�QAh��v�,�>P��>qg?���=&�=��xP��������"�4��>q�;?Khv�*2����>\�k?ǒ0�tw���>XN�x^�
q徺����0>	J#?��s>�B�=Q4���_(�����|C~�ux)?�?̓���*���~>�;"?|h�>��>�
�?7H�>�þ�vO:�`?p^?Z�I?uA?)�>��=򃴽��Ƚ�L'�vz+=9��> \>�(q=(��= ����]�7���B=�R�=�/ϼw���=_�;�ս��V<���<�A4>[�ܿB�G���Ͼ���G���z�����`7ѽV+�� ���4��զ����h��5�����|R���`��ߌ��x�;��?���?����7v���9��5�����>��|�	�l�ʨ��s��=���g�ؾ�����! �f�O�qXj�Cyd�;??EP��ҿ�F��l��c� ?s�??=�V?�w���G�0�1�>�*�>��A�N��m���������Ѿ��?տ�>?����S=��>���>��{> >>F��
J��K�,=���>(9?3M�>�B���\��ڀ���Q�=�*�?�P@�D?Q�!�����=9��>&?TF>�a�f�����k׸>&]�?��?Z�<�~S���_?S�W<�PG��O��T��=�?�=�f�=ν�:HO>U�>(M��"G�e� ��p>a2�>�;�<p�˽7Nf��H��A�P>87����ۼՄ?�z\��f�ӣ/��T���T>`�T?�)�>�6�=��,?�7H�e}Ͽ��\�v)a?�0�?��?��(?�ٿ��ٚ>��ܾҊM?D6?z��>d&���t��~�=}6�|ˤ�W�㾰&V�'��=g��>�>�,�l����O��U�����=h���ƿU�$�%z�d�=���^\���罶Ԫ��wT�����Go�\T�`�h=��=4�Q>l�>hW>MZ>�fW?F�k?�a�>]�>u�ъ���ξ�� \�����ݰ��M���أ�8�ύ߾�x	����u����ɾ=��Í=�;R����� ���b���F�0�.?n$>b�ʾ7�M���-<�Sʾ-���<N���ޥ��7̾�1�Rn�R˟?S�A?����p�V������Q{���W?}f���款6��=���-�=P+�>)��=��"3��|S���5?y�?\��
E��B`r>�s!��Cr=��2?B�>��<�,j>
Z@?�\	�i���=~0>�M�=���>�t�>.v�=����麽�\?�6V?%��:卾�ߙ>FԾ��`��������=���K�=2�>ŜY<%v�������a�	��=�%Y?^c�>{�1�-�og����:��b=q�z?��>���>J�X?�M?��%<�2���mQ����|ސ=֮R?�Z?}��=a���J4���䘾�Z/?Ɯ_?�jX>����辥/�[��a�?-�w?� ?`���{���g����<?�Zt?'�Z��{��p�!�����T�>~�?>B�>Hm$��8?ռ?����m���ŕƿ]2���?�@��?�>�����;>pZ?y~�>ਔ��[뾿�k�����
�5=gB?��о�ƅ���%���P���N?�2�?�?�7���g����=�ٕ��Z�?n�?����nFg<L���l��n���|�<�Ϋ=��G"�����7�Z�ƾ��
�����@࿼쥆>9Z@UU轪*�>ZD8�R6� TϿ#���[о8Tq�s�?Ѐ�>0�Ƚ\�����j�MPu�I�G�+�H�����K	�>���=�Iu��������OD��;���>���:�(�>�q����cy��r�Y;�un>R��>�	V>��������|5�?��@]Կ�����	��Fo?v�?rƄ?��"?������@r��33=>$??�7k?�VS?�� ��)>��Z��pAl?h�ľ��b�y�B��C�yr>�y@?N�>U�-�1��=��=�B�>�>|�<��m¿#լ�kFǾ&�?�D�?H�t�?kȠ?m??ɀ�����ܹ�-X(�P�8=��P?�'!>C`����6��C�w`W�\�*?3bQ?�Ϫ� :�?�_?��a�O�p���-�ݹƽ-ء>��0��f\�p������:Ve�M���Hy�C��?_�?q�?���Q�"��2%?@�>���><Ǿ���<^��>�$�>�N>b_�-�u>��{�:��o	>1��?�y�?zj?��������F>\�}?��>��?zx�=�?|>7p.���=|�D>�Ї>������>
MR?��>��>b���T(���4�-F�@�m.D�E�>�l?�C?~��=��"�ɧt�k$���+���RV>h��� ��4Wٽ߱T>�s>�D>)�]��$̾�-?t�7��ֿ�����K���2?�n�>[[�>��:3��Ō�I�S?w �>�: �7e������1��&�?��@rG�>����Q��=f.�=ᦁ>��Q>�Q����	��ׂ�W�>��5?�$i�	长��}��>��?-	@bB�?�n��a	?G��KJ����~�����4��(�=�7?q��|>n��>�D�=��u�aժ���s�rC�>�I�?�R�?���>��k?
/n�=_A�E@/=ź�>�j?�~
?Ţ���K�4�F>�D?��(E��Ԩ��>f?
@��@�f^?�]����忈���4���������=:�Ȼ��=_���>@�3=��P=�Fh;+� >f�4>o(>�o+>;O,>&�>\AI>A���C$�~И����f�P��:�mr-�S~��N�7�R����®�[7پ�v^�#�52̽Wne�� u�Z;�:z��=ǎX?<K?g^v?^��>>)���<>��X��=54��L�=e-�>T0/?��S?��&?0o=�ޗ��B`�j<}�W�����{��t�>01G>4��>��>6��>�'Z���.>lB>j�>H�=)�t�~!g���X=��V>
֭>���>d=�>��^>zn�=����.��|�k�C�i��� �6�?Yj��	B��N�����߉�;3�=�?y}�=Ь����Ϳb8��T/G?,���)��1�UlE>��6?s�L?��
>�S���q���+>�G��f���>p���_�_�׈ �j�>Cq?�	g>�u>��3�Sb8�`�P�J��j|>[F6?>۶�u9�߾u���H��lݾ��L>D��>dFE��\�2��Cxi�7�z=�f:?u�?�u�������su��x��W�Q>�@\>Aj=;�=�OM>1&d��mǽ�GH�!/=�(�=��^><O?�4,>v��=@�>$M��h/P�bx�>.vB>:,>@?1#%?\�B��o���=.�c�v>��>��>c>�=J��ȯ=�n�>�b>S��ZD�����@��W>��~��_��6t���x=[Y���q�='��=�� �Pw=��w&=,�~?����䈿���i��xlD?�+?�=��F<��"�5 ��qH�� �?�@Vl�?V�	��V���?�@�?F�����=�{�>q֫>bξE�L�\�?��Ž�Ǣ�>�	��$#��R�?�?�/��ɋ��l�7>W^%?B�Ӿ�D�>(s��[���64��.����t�:[�>�>?�<V�<J������>�P"?x�ԾĢ�T'���'��y��>��?*�?v���<Թ�ܯI���>j��?(3l?�sR>˾#m��)<�=�2"?[ga?r<�>L��k���]�>A_�?4�c?��E>1��?��p?a!�>T�~��.�VI��dw���lg=���;i��>�p�=�z��TB�%�����x�j�q��CjV>�b:=�~�>��ֽVԲ�u�m=�Σ��T��z'����>��f>�fW>IV�> K�>8�>y��>ڭ<Y/��\����j���W?�V�?��!�u�n�PNc=�E�=�PW�d06?&h;?`���VyѾR��>|�H?�l?�P[?L/�>���Ζ����Ѭ��0�����=���>�S?�bI=EX�>���᛾���>��$>\�=8���]��R���Ǎ>>�-?߀�>���C?h�(?V^>s��>ZG�v�����<�Xǩ>|?_X?�\�?�?47�����_�����0�U���{=�6k?^}.?�b>��������6��d�<VRX�}��?�S�?y]
�3K?��?�C@?%!<?(A�>�l�j�ž.��r�>[*?J��-�]�1�1��GH���?�?�P�>��7�
����ｱ����c�?.?C?z�?0}�	�i�T��FyQ=���0
�y�c;��=��X>$G�=B\����.=�k$>�tC>&cU�qK��<�$�=�Xl>C�=s�2�m<�j(?��-��`���q�L8z��\,���>�6�=���pl?/!��@8��)��~���l����?my�?�֑?ĔW=��n�q:L?O~?�m/?��>U=���j��ĨӾ��̾6�ӾQ����C>�B�>�i�뫾�Ŝ�����mv���E���@�D�>>��>�9?ͫ�>�uJ>S�>V;��&�6����Yk��ع[�M>&�|�F�&+�A���풾��yo~�t�žh����>�����4�>��
?��B>9��>�7�>�����>{�y>}��>G�>N�(>SM�=c2�=>*��20���P?�󜾋�.�?��.�h� �M?b�a?00�>��:9x|��}��r??f�?	ќ?�?>�Wf�r�����>>��>t���E�?#�>��>8)��`�������71ڽ���=��>���<`�[�lw2���c�%�
?�J?`4�O �>�*��ᾔ>>�N�?_C?*�;����}�q���f��'S�r>Xs��7@p�D���A������t����t�K����+?P&]?�,�S�Ծl���Q�d��R�����>�s�>5 �>:	o>�r�=�����#���_��U��sh��w�>9?��>'J?�;?�R?�AK?���>�8�>n��.�>��:�d�>��>x�8?�/?��/?�x?��)?K�]>�������5�־�?�m?��?=��>�K?"b����˽�F��].ιo�{���u=�f�<$нT�`��wj=��U>�!?��"�7�E�q��?��>�>?Ѝ�>t �>M��
9n������?�?�ņ>ӆ���r��,�w��>�r?��Q�$�p=<}_>e�,>I���>��;B=�=�X���6�=維�#�"�t�<�pG>�/Z>{Վ<;��b�
��9��=	��>�&+?�nF>�&�=�����ɾ��6�(Ae>��>�SJ>�bw>������/�����k�;�}>*2�?<q�?�3���(�=�04>����B=J ���S�|>���>��>P�`?坕?��O?t�?�zL>O�	�]ߘ�-��oʙ�i�?",?q��>����ʾE𨿢�3��?�\?�;a�����;)��¾� ս��>j[/��.~����wD�����m������6��?y��?,A���6�>v�%����]����C?��>\�>y�>�)���g��%�3;>��>dR?�#�>��O?�<{?�[?�gT>c�8�`1���ә�H3�m�!>B@?ޱ�?��?Ty?Et�>��>��)��ྍT�����J�Ⴞ�W=�Z> ��>�(�>��>���=ȽVY���>��`�=3�b>��>3��>��>Ӄw>�O�< a<?$
?�ڧ�Q%�l�<'��t�þ�U?��?��>w��*�*�[�@�j����>�M�?)��?rG?��S�+ׂ=�i�����~;���s�>��>���>��<S�>L��>9L�>�\�>Qhy��%(��{������Y�>?Th??Խ�ȿ��e���A����������	��׷���e�/��=6���]������=�I�ۚ�*�����������s���h?�=��>AZ�= 0< �J��P<�&=4�K���1=#^���*=щ�g�W<�y� ��8N��}3<��u��6̾e�z?��H?�-?^E?��~>��>�y9��p�>^��b�?I�V>-7g�"���=t/�_.��@撾��Ӿ#)ؾ�ec�~��k>��P�'�>!�/>��=��O<ǃ�=�݋=�B�=;���=<�=]�=>/�=�g�=��>�U>�5w?��������59Q�	���:?FB�>1Y�=Xzƾ$@?8�>>4�������k�s%?��?jW�?��?)Qi�bY�>��񠎽V��=Uݜ�^2>{��=}�2�Õ�>��J>��cJ������.�?Ņ@0�??�ދ�ڞϿLL/>d�~>Ǵ>}�a�t8-��j���b�;���3?�1��=���J:>�IO>
o�߾*v<��>�Ġ=�Q�� f�?	==�&ҽ��7=�(�=�{�>V�e>P��=��R�e�<[?B=��=$��>�L=�I�<�e���=�N�>�<X>Vq�>d?~D-?3�H?7X�>�r�h�~���2Cq>��
����>cJ��|�=z\�>Y�a?�uh?"V>?�	�>�A=B�>�u�>�0�� j��f��4敾���X��?��?�#�>ޭ�����	��GY�����.?E�(?f�>E��>�U����7Y&���.����7#4��+=�mr��QU�0���?m�4�㽥�=�p�>���>��>8Ty>�9>��N>�>��>�6�<{p�=ጻ���<� �����=������<�vż����bt&�;�+�J�����;W��;M�]<���;���=&��>%^>Ԩ�>2�u;�w���]Z>�#���Uj�ֿ�=*Ȿ�)C���t�����~�f����u~>�9>�G�����
?��>��>�?
�[?^�=����s оO����[��~8��iB�<'q>>B��ۻa�.Xp��L����y��>]ߎ>��>̻l>�,�
#?���w=d�>b5�A�>�|������(��9q�@������Xi��ZҺϠD?�F��6��=q"~?�I?5�?���>j���ؾ�;0>I��g�=��*q��f����?'?���>�쾑�D�"<پ�:��s)�>�'<��v_������E$��?���I����>������ƾf��;�v�_����E9��.��>\�>f0K?.��?�����J��}�L��=��ӭ=S�,?��s?���>��>e �>{�ѽ2w���͊��D�=K.^?��?ʦ�?��P>���=����f�>G�	?0�?`k�?6s?>��^�>�� ;�['>C��Lh�=�<>}4�=��=��?62
?�J	?jL���	����O���\����<��=ߖ�>s��>��w>�B�=>�_=f��=X7Y>!��>�d�>�8d>���>{@�>:����&��x?Eӆ�@�k>��,?��g>3qS=[�M�HV���Dϼ��G��h���G`<G���_̼��=��'>�r4��>̿P�?�!�<�p�^?�(�,4���i�>j�d>*ɽ�R�>�n>�c?�E�>s#�>Mgq>W@�>�m>�ܾ$�>�����@�0�I���c��EѾ��\>����̽H����q(9��S���1��hd�s����WB�N�=�z�?�z!���l��&�V�!��
?���>�>?,W�j-S>���>���>�9������q��E'о�y�?��?Z�>O)>��f?�Q�>�'�ט��)X���^���Y�¢��JJ;��5���L~�4�W�⓳>se�?V�c?�E>?R�ѻ���>
Y�?�|!��g-����>s[?��P�_��=�Ӻ>����Fe��������UeA�]x�>�.r?��:?6��>����Fⅾ�>��*?\Rx?��?��1?o�0?AM%��o�>�묽c�e?���>wE�>�5-?U�*?�*,��I�=��K>Fm<���ǽ ���%��(�����=���8����
G<x����>u�=X��r��=o��nւ<@ؾ<��<�Ѹ=�o�=M!�>�E^?�t�>�k>_�;?�i��@����^1?���;����G�� ڧ����Q�>Ws?��?�rW?�`>�>�`n6��5>�`{>E>nbb> �>�`�**�O��=��>W>�m�=�Վ�4��̥���t��tw=i�>���>R�|>8���A%>�š�>�w�o$c>�7K�˹���S�}�G���0�xJx���>��K?��?5��=XB龝:��J�e�zu(?�A;?I�L?�8�?wޙ=ܓھmn:�z�J�4X�d'�>{F�<\	�@�%.��k�:�A��;�u>����q.�̈�=?F���◾n���A����4����*�&��>޻�nEȾ"��� J>R��=ur�И/�;뙿W���[�F?��p=��t�h����W޾�<:�%?�O�>�=�y�Ҍn�9"̾��!>�h�>$���S	�L����z������>mvD?E�\?>��?�:{���p��JC�>����K��3���P/?=��>V�?1;>z�=IĴ����Rc���D���>���>����3G�8\���\�� #���>,�?@�7>n:?@*R?��?P�]?ڎ%?d� ?��>�����X���1&?��?���=8�ս��S��9��7F�U��>:�)?]�C��V�>[C?Б?��&?_�Q?b�?O	>�� �2(@����>~c�>Y�W�3L��Ɇ`>B�J?�C�>_JY?��?G>>�|5�7â�Z������=��>��2?D#?��?���>��>䣡�D�=��>	
c?X/�?��o?4��=U�?�.2>i��>}�=���>f��>�?�SO?��s?A�J?a��>�<�5���G���`s��
O����;��G<\�y=9��CJt�G[�F��<�7�;GE���e��W���D�u��A��;�3�>t>`>���.>�6þ����[@>�y}�k��#���k;����=���>9?Oǔ>8�%��#�=���>��>U��U(?@�?"d?�;��b��n۾8�J��6�>�dB?&��=E�l�@u��ܙu�|�n=�n?�3^?��X����9d?��[?�����=��7��N}J�ޮ���X?�Q ?NN'�Zr�>��}?��n?��?�j�z�o��ϛ���_��n�<��=њ>E+�Z�_�K8�>��+?��>11X>�J�=ޔʾ�My�槾0�?)ˈ?�/�?�V�?�->�Wm���ݿ�/
�����N,]?[c�>�7�?S�I[Ծ*��j���g�̾8)��^1��ת��u疾p=� �W�-1��Ȱ�=��?d�r?��w?O]?���-g��Gj�����!Q�C���?v���A��?9���D��ze�����)>侅鈾erE=+����?�b�?��#?J|A�Cw�>�6��0��`'ھi9H>�[��CU�]�=�r4�N�=��=B!V�o���}��r�$?f{�>�_�>�S8?X�Z�Ӑ=�o�1��n>��:��<>�:�>~��>��> ��R�8�i���̾Qދ�����w>ana?��B?��s?5�%�)�+��*����m�	����M>���=�Zn>�K������"��n?�O�v�/B��쉾<���TP=93?pu�>&ǟ>��?0�>^'�����})C�~�"�'��<�#�>D[?Ғ�>��h>A�ͽ�����>֫l?�5�>�ޡ>[���!��|�EʽXB�>}�>���>%�n>��-��[��(���P���9��]�=�0h?F��'�`��`�>(R?L׽:Ϗ[<2�>Yy�"J!�b�X%��	>�e?��=�=:>��ƾJ\��m{�H1���n)?a9?
⓾�w*��/>�!?w�>!C�>��?���>��þɏ��k?�_?��I?E�@?���>3�=����	�ɽ'�0=)v�>R�X>�Nh=6�={��;�Y��+ �P:F=�h�=�Լ[r����<�գ��C<	,�<��2>v���N��^��@V������j�1M,�*ڥ�b���冑�����Җh���c�	D�;K+�S�C�'I�ED���?��?��"�BH�s����₿��7DO>��m��"��趾_7�UJz��`�} �����OG��U�v�^�}j*?�)����ȿ�ܢ�F�侻p&?�%?�th?_����1=�'4P>���=`�ۼ³��Ϛ��3�̿ߖ�3q?��>K���e&�6��>RX�>���>�?>�)������x�<�?}?{�>�'z��¿*=��E��<���?�p@K}A?��(�/��jV=���>	?�?>�H1�AG�~���jQ�>}:�?+��?�mM=!�W�� 
�Xye?V�<��F�L�ݻ��=A�=�Q=T����J>�S�>Ԃ�$OA��+ܽ��4>�ׅ>~�"�Y��L�^����<�]>x�ս	E��5��?��\��we�}k1�Wဿ�U>�pT?�8�>b�=h+?�I�}�ο�\]�Zk^?���?��?>�*?����Û>�Qྣ�O?�6?�U�>�w&��u�hK�=S?ü�9�*�^!W���=���>�O*>Ŋ �����^���9��=�]�&�ſ"��b��ƛ<�i}���+���+�z@ؼR��� ��!�B��=e >?�J>ʰ�>B�d>��b>�\?��y?���>�@>t���ۯ�������Ƚ�ʋ�:z��і�#���˜��v�_(ʾV �/�5�)U��b =���=�4R�ٗ��2� �N�b��F�3�.?�s$>�ʾ��M��"-<�pʾ���� ����ѥ��+̾��1�'!n��̟?��A?�����V�=��]U�����=�W?�D����鬾W��=b�����=�&�>���=���:!3�`}S�n�1?�?y�̾3g~:>���	9=]�0?z�?��=Ě>O"?�B%�k�����Y>X>&��>�q�>���=�J��¡߽�?W?.#�[�����>�Ѿ)eQ��� =ύ>��H�Xg��nI>���<��s�V=��{�����<<��h?�i�>*����Tݾ���=�(>�@�?�&?��f>B�?,�x?4b�>��m��j�3j9��2I��DQ?���?y�<>o��vZ�8��]J ?��|?H�?ث���ۋ�ǩ��
8��%?2W�?��'?ճ ���s����~1���*?�f}?������\w���	�� ?�/?!�">���F�>>�"?�B�;99���:ʿ��O�q\�?;Z
@�?˓�WAŽ_h>c�?:+O>Qҷ�N)��wc������=n��kE�>�e���U���!��V��C�C?�r�?�?+G׾O����=�ٕ��Z�?��?v����Cg<`���l��n����<�Ϋ=���F"������7���ƾ��
����pῼƥ�>=Z@AV轑*�>�C8�H6�	TϿ'���[о�Sq���?f��>"�Ƚ����?�j��Pu�l�G�4�H�å���;�>��>Q������d�{�pw;�������>'��6+�>��S�����{��/�3<���>Q��>˘�>�i��q����͙?����Hο����X��L�X?�c�?�n�?�d?��:<o�v���z��I��)G?C{s?O	Z?�'%���\�m�6�r�j?a��uV`��4��FE��U>�"3?mB�>Փ-���|=�>���>�f>Z#/�:�Ŀٶ�[���w��?P��?Lo�
��>���?Vr+?�h��7��V[��@�*�/��<A?~2>n���[�!��0=�ђ���
?�0?�z�	0��_?M�a���p���-���ƽ�ڡ>h�0��d\��^�����TXe����By�W��?�]�?R�?'��� #��5%?��>	����9Ǿ< �<3��>�)�>;*N>OL_���u>����:�dk	>7��?U~�?�i?I�������S>n�}?���>!�y?kz�<b5?<�=x�m����=�H�=Yp>c6ۼ|��>�!?��>\ZL>I�E��8�m�O�T��b��6C�[�>�?c,O?��z=��V���=I>�!Ic��[�`ma>���^�A��Ky_=��=^/->���_*r���9?�=}����rx���;��dUX?��>?M>��H��(�=]�뽗1Y?���>��
���:j����� �?~3@���>����n����m>���>�Tt>-B��.Gk�������=�]K?���{��jjy���(>�?�'	@%<�?�����r?i��9����|�G����� ��>�1?�꾥 �>o��>�|�=Fft������qu����>?W�?��?�
�>�Li?��j�H>���/=È�>�`h?<s?�z�����G�9>�?̏
�����K��Ⱦb?�]
@w@��]?�⥿H�տ����_���������=yd�=k�>�C��y*�=�a=hR$=Η�Ih>S��>�RS>hi>�FR>!\8>�>͆�4(��饿p獿 2�H������ZB�s ��ɠe�����g��mཾ9��c� ��!W��0K��8��}����=v�X?�J?��?���>@y8�+Z >�@侇Y=j�"���!>���>B?(�F?�R?i�C<W��3I^��mu�?X��Go��|S�>�zk>�j�>���>x��>��R=$K>-�r>̜>q>�{|=\��<
vH=E3>X�>[��>�l�>�C<>%�>-ϴ��1���h��
w��̽"�?�����J��1���9��ݦ��j�=*b.?�{>����>пK���o2H?���e)���+�P�>g�0?�cW?�>t��d�T��:>���~�j�`>�+ �+�l���)��$Q>/l?ۂ>^+|>z�8�AK-���?�����J�>I�9?$��������q�}�=�ƔҾ�n>RB�>�Lļ�g#��i���)��G��+�=N=?|3?�� ��ծ���m�Mʾ�Hj>�\2>)��=��$=q9>ի��@�׽��A>�<��=QGU>6#?�->&�=�t�>,���2pO��|�>$)C>c'>�D??�%?T)�����@����-��s>̻�>��|>��>H�H�a�=�v�>�
b>��
��������/�;�2�U>>�l�_Y���g��	w=����M�=�>�=����F8�|�0=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾAa�>��þ�Ǒ���������Ew=O�?s%?n�����9>����|?=!?��۾�����[�x�/Ũ>���?ﳥ?扎�+Ǹ�7F�p�?��?t�9?��#>�N����V�L|$>��\?�_L?���>�����K�%��>U��?i�?�YI>
b�?��r?#��>u���.�z��	>��T�z=�;�ϐ>��>_��a�E�Db��S+���j�&Z���_>�l%=��>ɪ�Ѻ���=�㉽i����f����>��o>��L>�(�>ϲ ?)��>�D�>���<�~���e��xw���Q?�?��(���^��>�#�=���9�'?~�%?I��=�E���>�nD?め?kQA?>.>B��s���)����|��C�x�--c>o?@.�>����@e>��
��s��%9D>2h�>D�Z�ܾ�w��q�=�L�>��?C�>Cf:E%?�?㸁>х�>ق?�Yр�|'E�`�?�Ȥ>�;?��?��?A7ɾ�m�Ҍ�,N���<�G��>��s?�!+?1�B>�;��䭪� Ò��m=o��=�n�?C�w?	���#n!?��?KGr?`�d?��%<p��ή�a5�=���>ۅ"?�����B���%��4��?�F?�s�>@L��
�Ž����K�ί��F�?	Z?J�"?eU��a�Z�ľ�'�<v�E��׺K�n<�(}��g>>Nǚ����=��>�\�=��q�5<9��\<���=�[�>���=�R:�嚽�B$?$�����1�νKB���,)����>-<�=�cžq�8?1����,~��+���9�������?N��?;S�?����~�]�g?�Zz?��4?�_�>݀��~��"xȾy��?e��$~�\��=���>���=vkʾ碭�E%��F�~��"%�_r`�{��>�\j>�
?ށ�>BN6>��l>t����E�`�߾��
�?O�r�3��V1��a�A��uޒ��M�v�_�I ��RO��ET�>_�-�H1�>�G ?z��>O��>a��>u~Ͻ�T�>I^>wn�>c��>4�>�Q>x�M>��=Fs���q?�'���R������t���`? i?��9?h-�=�҄��1��-Y?�v�?�?Qk��֌�X$>����>[�?�ڃ�vP?�D���gM��
�>r�ƾ��ƾ
g<�)���@?om޾r�P�����F[�(�?@�?X>ϼ8�PȾo��i9�=NƂ?��.?��"��N�r9o�9�O�c;U��ɼ�EM�e�����%��+m��A���΃�Ӥ����&�	F=k!)?-�?
��J���䲾��i�kt;���>���>n�>:v�>(�R>���6�-��]�d>&�+i�հ�>sy}?:��>�K?��<?WQ?�K?�ώ>���>����_�>uR��	�>'��>��6?�f/?yA/?3�?<�(?߽`>�G�����)g־�@?�?��?�?>��>δ������`˼~(�� �|�p݉���=<?�<=ӽ�}��=�0N>5X?@�� +<��i��zL>��6?��>�^�>%㖾z�g�0><<]��>��
?H�>x����s�o9����>�c}?��3��N=c|(>�7�=<�?��᲼���=d��=�v/�������s�=\Ò=@��<�,�<_@ <�F�P�(��[�>��?{��>C�>i��#� ����m�=c�T>��U>d�>�ؾAm���Ɨ�Sbg��Bv>I��?��?��h=��=�'�=�-��=P�����c���
�<��?�+#?�T?��?B>?(#?�>�����������N��C<?p!,?F��>���c�ʾ��1�3�Z�?s[?Z2a�c���:)�ڎ¾�Խ}�>X/��*~�����D��u�����i��`��?ҿ�?�QA���6�Nu�����fY����C?')�>mR�>��>�)���g��!�D.;>"��>�
R?��>��O?(�z?f�[?�KT>�U8�k(�����)>��@!>o@?nt�?n��?~�x?GW�>�R>n�*� ��Q���,����h悾��Z=�8Z>���>݉�>
��>D��=# ɽ����Jg=��ϥ=��a>���>!�>�3�>Hw>�o�<�SG?#�>�M�����ɠ�����Y�#u?z��?Gf)?�>�<��5�E�L�� ��>���?��?t�(?��R��v�=eּ�����n�"m�>l�>Xڗ>���=g�Q=�e>kv�>��>�F��7���7��L��F?YCE?�O�=� ʿ��l��8�`��Z�Y�R���f(��O���s���=�׊��������;�Y���8��a)��M����:w�z?�C�=��>���=�2A�Y�?���<��7<\ =�th=c;��K�+=a�S�1X�񴷽���;ʽ���ܸ����׈��;oy?�~;?��O?r16?)%�>PNA>�#j��p>Q�9�'�!?9_>����S����Ck���ా_~�C޾���˭��@�O>��<��P>���=ii�=��>�~>X:>��P>iB<R��=k��=So�=�D<�P	>ÕQ>R��==Iu?�툿�t��w�i�F:�S|??��>��^�Α��ѠJ?ϼ=i�y��;��p�/���`?�?0-�?�?S�3�(�@> <���M=�<!�~��Ԛ�C�:�r+���>�"=?JA��(���Y�����?��	@:?�<��͑����_>F�7>j�>0|Q�-�a�W��6^��8`�Y�?��:�̾��>��=���bľ�"/=~>1>�EE=��!���[�8��=�򄽨8=�.r=���>D9E>-�=�ѭ����=W�;=�T�=V�T>�&���B��;��5=���=�eb>�#>�o�>L�?.?Űf?�ؽ>W�o��=վ?���R|>(��=N;�>�6n=!->��>��4?��=?hF?�x�>w�=�T�>�>��$�G>l�*�QC���k<�݊?�\�?���>>p�<�1��H��e:�E?ҽ�p?�)2?��?s�>�U����-Y&���.�A����7��+=�mr�RU�����8m�A�㽰�=�p�>���>��>1Ty>)�9>��N>��>Ī>u7�<�p�=䌻F��<� ��>��=ŝ��
�<wżt����p&�|�+�������;�;��]<���;�y�=��>5��=Ki�>;�p=U��2�=R.��Q,b�V#�=��˾��>��#p�v
v�F��73$�/!>h�">�9����?��,>/��>��?�%^?
h�=���@߾F;��5�*�ؽ��=hƚ=��6	a�Ǉl�<�W�� ���>�ߎ>�>Ժl>?,��"?���w=�⾌b5���>�|�����)�P9q��?������ci�q�Һ}�D?�F��m��=+"~?��I?I�?���>g��N�ؾ�:0>�G����=^�+q�ci����?'?���>�쾯�D��
˾�	��\��>:C��O��o���0�����Ḿ,��>|���-4о7�2�-�� ���̓B��us����>�O?���?��c�����pO��D�"�����?��h?�[�>i�?��?����i����~�ⱱ=�gm?w\�?�[�?�p>.�=M������>Sl	?}ʖ?ڄ�?�:s?�-<�bH�>W�:G�'>O뒽�u�=��>0z�=���=�4?�n	?�W	?P���K
�t�ﾧ	�a�`�Q@�<���=��>l5�>u3w>�0�=�#g=ܽ�=�Fd>Ϝ>�H�>�f>K�>�Z�>k���]�^L?<���}>�=?���>�OC�h'�����P��:��'�������*��ҽ��m�=׌3>�">�pY�%��>X-��d�?L ��� ��5?�T��̒��q<>Z�=�*�<��>q�	>���=.�>]L�>���>��>H�;>���,6=5Δ��m�:�o��ن�K�j��i�= ��h�;���ޥm��"�^]�����I�L�����l��}<ͺ�?��� ڀ���#�M9�Y(?�p�>��=?��2��ۣ=�	y>�5?*u>����R����{����8�?W8�?S�/>��>��X?
�(>ȕʽ֬G�o�]�,G\�Z�t�H-���U�#�����c���9�W��=_�?�k�?;N+?�Y�JIL> :�?J��4�9��>;�W��H���>(��>�ⴾp˾�H��u���o��U?��t?�?c�=>��ƻ�$m����>��R?�]?�!^?1�>��6?���=��>Ƌ�:a�U?�q?	?�X?ƃ�>Ә�i�]=���=M�m�m,� v�>>���L�n�=���<�rZ<D�=٢��@}=��vr<p���Kl�;:ˉ�>�"=Y�6<���=���=�l�=Fs�>��^?͌�>!U��#�`?�m־?������C?��� ��A����'�G5K?ʫ�?&��?��>��={y��uA��	����>�Aݽ�I>ab9>����]���>?�v>�A>�z�L�>S޾���qh����Xgc=��>=��>j㮽��->仩�'�j�	�,>�^��ξ��J�o
H��"5�>/����>�G?z�?�|�=MB޾e��Q�f��.?-k(? t_?�~?V��=7�ξC;��}H���!��E�>��=�f���{�����?�Z��G罉�>�]����*�e�t>ͻ���ɾL����o�'T����	׾�%���� ⠾1�[��z�=�d4>6��=4�m��Y�ǿ4J0?��=��_�s��޾,��>��>�E>�Ȥ=	���sli�\�iQI��>���=L�4�	��^R�iQپ��>iAE?��^?n��?������r���B�*���������%�ڲ?(��>��?�u8>0
�=U������qe�y�D�gS�>t��>6���D��b��F��B�#��&�>�"?�2/>��?alT?�S?�\?��)?�N?��>����۶��A&?���?
 �=_�Խ�T���8��F�e��>�)?��B�"��>6�?�?��&?ɇQ?�?(�>Q� �C@�쒕>�Y�>t�W��a����_>A�J?ٕ�>�<Y?xԃ?C�=>�5��颾Rש�\M�=7>n�2?b5#?.�?e��>gr�>�m��{�=�>.c?z�?P�o?]�=�?&�1>�A�>�t�=Q��>���>��? 	O?��s?�J?�'�>���<WH��Eõ�4/p���R��>{;p�T<C�y=js�C�x�s��6��<Z`�;e���� w�ke�|�@�7����;�]�>2�s>����6"1>T�ľPQ��\�@>x����e������:�׷=��>��?ٞ�>"z#�R��=(��>/G�>���a/(?��??(�';�b���ھ��K�A �>yB?��=��l�@���3�u��Ch=��m?W�^?�cW�����s?�dT?L���"LL�Qu����GP�#|�?�o;?K�z����>�\�?�ܚ?��6?��a�v	��������G�T&�p�/>�s
>�����q�t>M*Q?�%5?���>dg>����Ԏ�'re�!�5?U��?�~�?N�?��=�-v�ho꿎�ݾHĎ���c?|�>Zu���g/?i���r��X�����C��
Ͼ����Ծ4���B���l����]���꽏 �<n�?�z?]�q?��g?�x��Zl���h��d��r�R����h�/�� Q���"�E��0e��eԾ��վ�e)�+�=�Qy�vpB����?P�!?rs,��[�>�甾<	�k�Ͼ��N>�n�����-�Q=&~y�4T=��Z=�_�,v8�b"���� ?�G�>���>_�=?V�]�{>��3���>�d���S:>�ё>�(�>���>ݛ�R�1�'�ҽ=þ�Gq�ߐ���t>�uc?��J?D�q?����r1�*��h@�4ʉ��᡾��>>�a�=�1�>g:Z���(�PT)��I=���t���<��P�
��P�=`3?��>Z>N_�?R�?�	��Ρ���p��+���<k��>��h?��>1�>a"��1V��U�>��q?0$�>V?,׀�+�5���c�c8�=�E>�1�>�@�>�h�<� ��t�C��Y��ǜ��B�,�[����C?�GL���e����>��J?PĮ<;D={c{>�̆��Y�$8���-��k>+�?�'3=�K0>���%)��f��_�3��R)?&N?N�v�*�<}~>�"?6u�>�N�>x*�?J�>Qqþ�ڣ�!�?��^?BAJ?[5A?<4�>9�=$���Ƚ�&��+-=,��>��Z>�Jm=q"�=����\��*��tE=�=κмuҹ��}<G봼6N<���<�4>�ݿ��K�?BԾ�������f2�y����(ͽXh�����A���v��t9i�81�'����N�Fzf������l���?���?��y���wZ������k����>'�h��R�Y`��t
�̽��
4ھ�i���O�D8N��Yf�#e�Q�'?�����ǿ򰡿�:ܾ3! ?�A ?9�y?��5�"���8�#� >�C�<M-����뾭����οH�����^?���>��/��s��>٥�>�X>�Hq>����螾�1�<��?6�-?��>̎r�1�ɿa����¤<���?/�@#�A?�t(���wU=+��>��	?\�@>;�/���������>�?�?o��?��I=�W�$��MWe?��;��F��~���=�צ=�=:����J>^H�>�H�<�A��ܽR�4>\��>��!��]�5^_���<,�\> :ӽm���*g�?��t�c9m���K���~��R�>πT?:�">���=��??L%U���ƿ�dk�?�� @���?�S?Yw��Ip?E��8d?��Y?thu>�pA�y�g� �@���f>��<���6�G���)>)�>Y�>h}��[0���E���=Q?Z��j��0ƿ��"����^Z;�<���W�������S��P/e�0����i�)8ؽ��j=�n�=�_R>6́>�kW>`�[>�W?ϕl?�g�>�$ >B�As����ɾye;����f�������i��g��ܾ�*�i�v&�_ʾ�=����=�~Q�s2��D� �1�c�C�F��-?N�">�H˾4M�D|H<�Hɾ������֧��&I̾,f1��xn�Z��?�B?j����W�.���_ ����.�V?�����qA����=�eü�M=�T�>�Ƞ=�n㾈�3���S���9?b?����V�����M>pQ��cE->On3?}��>��=W8M>pyD?K)�=�������=�B<8�>���=A>��Ͼ�4��� ?���?2�������>0C�)䠾��=G�>�B���h�;�U�>;QM�4�� 佾n>xB�=@(W?R��>\�)���la������Z==��x?T�?.�>�zk?r�B?�<rg����S�  ��cw=6�W?�)i?2�>[����о�����5?0�e?��N>�`h�	�� �.�	U�%?��n?�_?���w}�������Rn6?�
|?合��˷����̝���>_k?=��>��&�4��>��?�+��W��ڸ��Q�S�p��?�@��?��=�~��K:�=u��>2T�>Z@8��G��	���龵5�=�?4ű�ܾ��_Y#��/��lK?���?�?�ھ�����=�ە��Z�?��?K�����h<A���l��r����<��=/_���"�Z����7��ƾз
�l���������>_Y@�:轒2�>pS8�(6�+TϿ����cо%bq�+�?�g�>�fȽ������j��?u��G�<�H�-���F<�>�n>������v�{�[w;�}�����>2��Y�>$/T�q ��¢��p).<{��>J��>)��>.Ԯ�s����ϙ?����Nο���������X?o�?Yg�?�c?�U6<Rqv�?�{���-G?�ms?`Z?��$�(�\��6�$�j?�_��wU`��4�rHE��U>�"3?�B�>R�-�z�|=�>���>*g>�#/�w�Ŀ�ٶ�8���U��?��?�o���>q��?ys+?�i�8���[����*���+��<A?�2>���D�!�70=�VҒ���
?M~0?	{�b.�]�_?*�a�L�p���-���ƽ�ۡ>�0�f\�IN�����Xe����@y����?N^�?i�?ҵ�� #�f6%?�>b����8Ǿ��<���>�(�>�)N>[H_���u>����:�i	>���?�~�?Qj?���������U>	�}?Y��>cS�?[��=�<?i��=�t���>�}>�4N>J*��k�>�=u?>?}kZ>�D9�t:$�}�C�GcG�X¾��;�-�>Y+c?�:?`%�>y,����0�����=#��0��;J~�a�	�����I�w>�W%>�����x��%��e�#?LM5���޿u��3���>?�Ӣ>���>�� �Qn�����X?>����=���M��+���e/�?)��?�~?0���<��!> ��>A�>)���K�%܆�!R�=}�B?Yn����[e�.a�>O*�?:�@zL�?<cq�5�?YB&��喿�����V�`�����A>)�?��<R>�D�>��=&�h�s2���Ѕ��C�>qG�?���?}�?�j?�}r��Q���=8U�>�b?��>���.!�AK>O�?�(��M���[��O]?�v@sO@<�P?V����Pۿů���9����žji5=
<=�>�=�= �2�=>���Db�=$T.�k��=�L�>*�\>�V>ʊE>t�0>wt2>3q��J� ��=��}���֖W�>�� �iy��%�#�^�������/����d���̽X�G�Ic�n?�M��k��=��U?'mQ?#3p?�l ?c�s�8�">zh��?�=�#����=���>w�2?i�L?*?ޏ=$̞��rd�Ω��ׂ��5��-�>�2I>��>2C�>%^�>�C9��K>]1?>˴�>s�=��=v%��2�=X�M>���>���>���>�C<>��>Eϴ��1��[�h��
w�M̽1�?p���L�J��1���9��¦���h�=Jb.?�{>���?пb����2H?$���t)�ι+���>z�0?�cW?��>0���T�;:>+����j�`>�+ �ol���)��%Q>xl?�f>�u>7�3�rf8�1�P��l��.f|>�+6?2Ѷ�z'9�۷u�k�H�qKݾe	M>9ƾ>n�F��]�� ��L
�Oji��7{=�v:?��?kϳ��ʰ�Q�u�T��_
R>�B\>#�=qX�=�'M>��c��pǽJ�G��.=��=��^>J�?�w1> =�j�> ��E�zR�>��G>x�)>U>?!C"?B���ۊm��~�c94�THn>��>�w>�>�P��N�=0Z�>�l>�/��4���H	��<�4`_>ER��E�^�I�8�:�|=-fc�o��=�M�=�n���5���0=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>>��I��Lg���o�����=��?GH#?�վ���=�X;�>��>T�Ö���K��\�^�ms?���?c�?��}���ƿ�I���?���?r�[?�ݲ=^��۾wT�>j2:?O�L?ev�>#)���ܢ ?4ʹ?%�d?ǭH>�v�?Xs?���>)y�Ju/����ŋ�c�f=,��;�ӏ>� >����#F�7ؓ�N���Yj�:k�b>�)=�~�>��u��᭷=�܉�fɨ�v�l�Ƕ�>��u>�5J>��>�$ ?�\�><=�>'J=�燽\��+����Z?�:�?:�+������^>�3=`�q��i/?W�N?�i�9"�-c�>��p?��S?��x?-��=�{��J���~ ����;��%=��=>S��>��>�/;���k�4��G}þ�%�>�W�>�=�A��2�mf�~��>+p<?�ђ>9^h> $?�,?^�?>��>w<.�A��\�+��4 ?�L�>WaG?`��?=5?[,����1+�����Q?�l�>�>y?��8?���>}��ÿ�#R���>c�=i�?��?�R��h��>+�?n��?Qn?�1>d!V�\U��;�o��>��!?|�B�A��1&�����?7?�)�>&@��;�׽S�ϼO���(����?��[? $&?_���&a�4�þ�{�<1w5��.;��c�;[�K��|>�|>/���Z�=L�> Z�=�Ym�Fm7�C��<�#�=В>��=�6��ٌ���,?x���<x��>�B=6�v�'�=�Xa�>��=>z޷�0W?�vS�u�z��K���4��ZQ(����?[��?K(�?3���D�l�pD?�*�?<�?[�>�H��8���پ���.�����
���>���>$̠;ټ���z��a���ό���O�3�(�?C{l>~��>u�"?��>� Q>U�ϾkR��m�x陾�U��J.�"�L�_S'�������E3��?"���c��b�]�n>qf�8�>�?�Ǩ>�ޢ>,��>��=�x�>ۄR>t׼<�R�>��>�Mq>g�>��<����xd?���N(9���E�qSL?Z\�?H�'?�fW>����[o2?ϣ�?G
�?w>�>a�m�t�1��>���>�	��)��>�f�R*���k>Y�7t���>�j��܈>��?��T�;�b�Fƾ� ?}?��<c���v����� �l=��?))'?��-�ڪT�ްj�x�S��WO�@�ü�Y��kܞ�؞&��2o�K�������넿m�+�lw=1(,?��?�,��?�後���:�f��5��g>�d�>y'�>�^�>:�k>	
��w7��\�G ��ii�K�>ف?�ڍ>�?I?);?��P?`L?i�>�9�>�㭾���>L�;��>�9�>�9?�.?�-/?F?	*?�a>���9��y�־�5?4�?;�?5?�Z?2����� (��B�a���t��-��	�=V��<k�Խ�e|�*&\=��R>2V?Y����8��0����j>�v7?ަ�>)��>�ڏ�\��K��<���>
�
?�k�>���Rbr�-[����>Ñ�?>���q=�a*>���=1p��=���l�=�����h�=V�����;�B)<�$�=���=�_X���<Po:�;ۥ�< ��>�p#?>�>*�>R�����$�N�>4�<��>{#	>�.�� ���͌��>Y��K>H��?l��?~�]=�z6=�T>˽ƾL&�����M��lT�>��>p%?x�8?��?�3@?66?0((>=;(�A���nN�����-G�>�,?䑑>��%�ʾ����3�;�? _?BAa�����8)�"�¾f�Խ��>>]/��2~�f��.D� ������������?��?�A�|�6�q{�I����r��͙C?�!�>>d�>g�>�)�i�g�? ��:;>T��>�
R?,#�>Z�O?B={?!�[?eT>��8��2���Ι�26���!>8@?���?��?)y?t�>��>�)�X
�qO��0����ނ��W=7Z>��>��>��>���=гǽ�F����>��A�=tb>���>0��>y�>�w>/o�<'iG?	�>�g���D�1[���r���__��u?���?�G*?��=����F����"@�>���?���?��*?�S��P�=��Ҽ�A���Cl���>���>O��>ɹ�=�L=a�>��>��>�
��]�8�%6_���?��E?�/�=��ڿm[k��ڽ�i��ľ"4&�l�⾼�d��C�.Q��?5���9;	��;�ӽQ�H�4,��̝�Z+��f*`��z?Ii�>� C>2q>�>�d� f4��5�s���.4���ʽA�>���<Ɗ�<�1��:Ob��{�<���;�{{�4����f?� /?4�'?CO?a~>���=�G=T��>��<nB?�v?>X�Z���ϝA�����'������Ś���e��;��8$>F�[�cc�=�|X>Ȓ=��A��8�=ٽ�=�9>9�=<�ͼM�=���=i=	��=?%�=#�=�?z������?�[�Nm���M?�>�]�S����;W?>�P=���Y����1�܌W?�@V9�??g�>a*����u>��ν0>j�=k������=�T�=�?��t�>�h�>��g���$.��?�	@A�D?�R��� ƿ̥�>�I5>��>	UR���0��cS��'W� �Z�dp?D7<�V�;!y�>:�=��׺Ⱦ��%=�U5>6�X=t��O]����=0��N==�da=�P�>��E>��=ڏ��=3�=�M=h��=��N>;�B�M��B���5D=��=f}b>>Q&>�<�>=�?9�0?�dc?�>"o���ҾA�����>���=�8�>��l=�?>v�>��7?��D?G�K?~�>,��=�չ>s�>�',�El��1��)���b�<Nh�?�s�?�G�>v<��?���z�=�`�ʽ?y?�1?^�?�j�>��1�߿F� ���1��	9�	
�bx�؋���<H���v��=ӽw�ܽ��=?q�>4�>G�>�O>�/>iH_>�]�>d�#>"�,=�Є=����K���qѼ�ā=�#�:ƪ=?ƻ�3$�;"�=}禼��^;)w =�Q!�/��<�'<��=qg�>�.�=�a�>��=�Ȉ����=���V���=H3���D��!d��${�M}-�`1�>}>�a�ҝ���
?��>��Q>��?��{?�*�=��E�S~�1h��ϯ"���K����=�̆�'���ɻC���l��tW�2w񾲶�>��>-�>��n>��+�r?��[t=�c�D�5���>c_��/������.q�=4�������h���1��D?$��W�="�}?ǫI?�Ϗ?�;�>���ԭؾ@`.>�-����=c����q����?e'?���>$�ƅD�;�ξ��E��?C���q�I������A��CR��ܾ��K?�������2�83�� ;��x?7�ȶ����>��h?l�?�t���{��wN�w���1W)=�(?-�*?�IX>�8?r�?�<~Ǐ��霾�2K�5o?��?���?>	�>5ܻ=죱�;�>��?���?�ؑ?��r?gW@�`��>J�D;݁">�l�����=��
>���=^��=��?��	?�	?pp��cV
�ڬ�? ��^�[��<���=`��>���>us>#��="�e=E�=/�_>�ϟ>�t�>��e>��>���>���x���?I�,�>�ZZ?�c�>��<��p�$>#=���=�X���.���<v��<I��=2��<b�Ľ�Q>�m��>�Ͽ���?��=����>��Ǿ��<���>[Q�>��V��N�>��c>	��>�<�>5�>�F>0ĉ>?1I>q�j�>�s�����]�]�O`��<ɾ��>��o�:�S�n,��r����	����e�e�����V�QZ���|�?�y��5=��9�6�K���>���>4�>?�~���q=7m	���?�} >S��	Ԓ�1݂���Ǿ�N�?��?���>��>sw?�y�>s�f�W�0�鵀�ʴd� �h�kj�-]������\��Bþc<>���?��V?)�V?wg��T�>>��i?Q��I������>n0/�}�[�E�>�sA>%�1|�E.���TJ����>�.Z?�AI?�`?���}�<���>��>�gL?�v?��>&|,?�� >g�:?�Ͻ�\?$O"?�?L�Y?w��>|���^B���ri>�����/�	ɒ�~�������=�(ü���^�'xR��ds��k>�:�c�ؼ�� :�1<w(�=|��=|�>3�~�T��>�!J?'v?()>/�"?��g�z�m�f�<�>�5�G�����0Ͼ��پ.�t>�^�?[��?�za?��>�>e�E���D�<���>%>M4>��>*�2>�\���^:>�(>���=J���U��þ�����N.=��B>�!�>�8.>~����=K�ʾ��0��9>sP������ߔ��N�X�1�k��n��>>�F?c�!?ِ9>4���w_��s/��jhR?(�/?�a?0��?��=�^���9�R	c�\!i��W�>R
=v�ؾ�����,k��Qp��=��� Xξ��=�依ӑ�[l\��Ma��b���]�$&�,���>������R����>�>����S�!��c���"���"O?��=`�N����Ƞ���j	>n�>1J�>(� �� ��u>������W�	�>�C��U��P�ͫT��l�>�|T?�TU?���?-T�>�a�+U�Z���3���"��?C�q>Z^�>S�d>�>Mܚ��(��Fk�%�O�F'�>b�>}��kg:��奾����	�yt�>�8 ?��>�<?uJY?��?4j?�+?�m�>`Ʀ>�˽�c˾�%?�_�?;3�=�ѽQ�9�I4�6S?�ڍ�>��)?�x(����>�?��?��)?��R?�^?��>[���C��X�>2��>;�S��ܮ��L`>.�E?���>W?檆?rxF>E+4�L���5X���-�=eP*>�0?ڒ$?�?�W�>���>�x���=�7	?¹m?ʵ{?��b?!n�=[j�>�V�>�ٳ>�Y`=8&�>���>*2?�Td?��?��/?F�?g�=�	�<�Y�'q	<��<��=�W���=���=ՠ����.=��<�ޔ����=���;��<����b�<Bk��6t�>N,t>�!��Ja0>�žX���GBA>���Ge��;Ԋ�#�9�ٶ�=���>B�?Oܔ>^i$�W.�=�ȼ>�o�>�����'?��?�D?}��;W;b��۾JNJ��>�B?���='!m��c��5�u��Kj=Yn?�%^?�X�����=�b?��]?7h��=���þŵb�r���O?
�
?#�G���>��~?G�q?��>��e�%:n����Cb�k�j��϶=)r�>(X��d�4@�>w�7?}N�>�b>�%�=u۾��w�Zr��@?w�?�?���?�**>~�n�,4࿵���k����M?L��>�ń�[k8?~��!��"��澹�����Jv�D_��$��Ͼ{�GA��R����½��=�#?�}?L�g?�vo?�(پĦ��	NI��i��\�ď
��0��4���:�3I�:�R��1پ�� ��;���/z�uXB�P��?��&?�-��Y�>�#��:���žR
4>�s��J��`I�=�N���nG=��_=�g� �,��B��E?�y�>���>��>?6Y�i@�)�/��.5��-��JF*>���>r��>���>67����(���нQ Ѿ�V��K���>�f?aTH?- v?87�6�"�����q!�����4�����.>a�=��?>r�O�[�����z�B���s���p���"���<��?Dҍ>���>��?�+�>���4o���YC���*��9�B$�>{Jw?ڽ�>��>�Zҽ[� ����>@�l?@�>�v�>�B��!��~{��aͽ���>9j�>��>{�q> ,��\�n��i���}9�y�=�h?oǄ�al`�\�>AGR?M�6;�Q;<���>A�x���!�=J��'��>@?���=�;>n�ľ]G���{�1u��v*-?��*?�$ٽ�s/���>kT�> %?g�>?j�?9�(?ҾS�ܽ�}/?�dt?�k?[?W�2?'����ҽ�ǽ�؆�^�=�F�>Ķ�=Ԝ#>	��=������پ?V���6��(��=j�T>�r ����<�뫼��=�tS�-�>lۿuZ�QξԃȾY��D����� ?�6����)�+��.̛��r<�C������;�	K�f�:�`�M����S�?,�?�+���T9����������K>��w>�ކ����g�˾�h�����ǆþe���Ȥ2�Vx�����z.���^*?H9���̿5 ��q����%?�,?2)�?�y����d��Hf>���=�軞�y��'̿ m�4f?���>2��F+����>K��>2�>�)G>TI��+7����<I?I�?�>��.��Yÿ�^���Y=���?�/@��A?�^(�&z��>7="'�>?T�C>Q.�`������>���?�ފ?��G=wdW����3+e?ч�<��D��6޻v?�=w�=�h=�~�a�J>�ϓ>���	�>�Y�཈�.>G�>�^�w���)_��.�<�v\> �ؽ��2Մ?{\�sf���/��T���T>��T?6+�>S;�=��,?97H�W}Ͽ��\��*a?�0�?��?+�(?)ۿ��ؚ>��ܾ{�M?YD6?���>�d&���t�S��=U4Ἵ���h���&V�6��=���>��>Ղ,���̇O��M��N��=�����̿�+����߆$<�<�Vͼ���Pp$���s�~�������U��S�=�`�=Q�u>B!�>�Jr>$�>>�WZ?5�y?.��>Xa+>6�K⟾V���'�C�0r|��� �	�5��o �Cȕ���2�ξ{-��n$����H��)#=�Bҍ=�/R�g���r� �g�b��F���.?;M$>��ʾe�M�
�-<�eʾA����؄�8᥽�1̾Q�1�4)n�.̟?��A?G���V����`:�Xr����W?�c�߼�gV��=���Af=�	�> s�=h��s"3�}S��0?�?���\����0>����$=�,?yb?��<�*�>�v#?+�'�9eֽ�Wc>�;>��>:�>��>�����߽E�?�LS?�������f�>�\��}1~�@�l=���=�"6����t\>8�<E���7Ӧ��.���y�<�V?ꌛ>�!&�7&#���x� p|�O2�=Ħ|?+�?/��>
�m?��9?�Z�<��޾q�B��J��1��=яU?�A`?�� >�}��1Iɾ?R��c�4?te?=�h>~�Q�Bz��%�5��b?��w?��?J߾� t}����t�� b3?'�v?\r^��s�������V�$@�>2]�>���>��9�mk�>_�>?#��F��e���dY4����?8�@���?*<<��E��=�;?"Y�>�O�H=ƾQu�����ҙq=� �>����2cv���3V,�V�8?Ƞ�?���>Z���5��խ>Z�j�m%�?��?Q����7<�X���_����-�s`�=S�#�%���C<�U�&�$צ�:���%��r�d�猁>w@��:���>��69��Ͽe�~�,Yݾ���Z�?a�>��(׉���u��^i�R=G�RnO��窾�r�>z>b���$V�����!jC��=f��>t꛼<u> XT����������{�<'c>C�>�Z>Q8��/����?�Z���ۿp�����/��f?$�?�?5+?���<b�%�.X���>�R?��?�K?�c���/�E ���u?��N�ȯ���Vr��q{��0?wRW?���>�ܾ{n���@�>vu%?fȥ>s&��ث�C>��^֝�Bϴ?��?�ݾ�?F�?5X?`����@����W���#�ȹ�>9�<;�.�P����.�:Pپ�>�>6j�>�m��8 �3�_?c�a���p���-���ƽPס>$�0�Z\��������Ue�b���?y�Q��?�]�?V�?!���"��4%?Y�>����#7Ǿ��<���>�*�>a0N>%4_�ӫu>�y�:�|e	>���?�}�?i?������E>��}?�&�>A�?�~�=}e�>�a�=���.� U#>�=�N?�#�?1�M?B�>�4�=0�8�r/�\F��ER� #���C���>��a?c�L?�^b>�+��~~2��!���ͽ X1��B��_@�8�,��v߽o5>/�=>�>��D� Ӿ�C.?���+U������W��x0K?<~�>�u	?|�Ӿ��]���#>q�6?Wܰ>�M�pv���b����ʽ�m�?s��?ޏ�>�o��2�<p]�=�é>���>�H�p[J�	����4>??�1��ف�@�f�D$>�?i@+Y�?�XW��	?���P��\a~���*7����=��7?�0��z>��>v�=�nv�ѻ��R�s�t��>�B�?�{�?3��>�l?x�o�<�B���1=M�>Ȝk?�s?3Yo�u�a�B>y�?������L��f?	�
@zu@N�^?\%տ� ��龱���pe=F�U;$�=M�-�Hd<0���+��e=^���(>���>i��>��>�f4>`�>� >�Z���(�С����w���6� $�D�H�@XB�����.��΀��4-��Wv@=�9E��@*�*�����%�VeT��k9>~O^?�@?#?j?�n?��q���N=m^�;k	�e�(�e�>p?� ?PCX?Z+?oE->4�^�|Fr�C6��W+�������>�ʹ<��>���>��?��=g�>n��>��M>��v>'��=ke�=Mj�= ��>��?�b�>5�t>�C<>��>Dϴ��1��j�h��
w��̽/�?����S�J��1���9��Ԧ���h�=Fb.?|>���?пg����2H?!���w)���+���>~�0?�cW?�>!����T�.:><����j�-`>�+ ��l���)��%Q>wl?۷f>�u>�3��c8���P�v}���\|>�06?���L9�c�u�_�H��hݾDM>��>�FD�[m�������%ui��{=Sy:?\�?�0��<߰���u��B���TR>�5\>�*=�S�=�JM>��c�-�ƽ�H��[.=��=%�^>��?A~ >��=�*�>�ҵ9�G*�><�A>a5>�$<?�$?/x��tC��������)�$Dv>-��>I��>>]FF���=eD�>�o>��
�!������<���R>���s�_�2p��o=G���g�=x<�=[��COH��A
=�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>��P�Ko��f$��E0��*ހ=Y?��|?}9��-$R�,P�<{o5?�e?�E��@���Ŀ�s��?���?	�?�xn�)���0�y��>��?:mX?�ԏ>�1��,�<����>)C?S��?�?uľW���"[�>v��?��v?~�>���?�^k?A�?5��=8F��������ѯ<L�R�'_x>{ݻ<�T��7���{�
�Z��^p���+��"d=-:=H}�>�a��`���o=>���ny��\���9U>���>e�P>�<b><��>��?�>�2I���˼�T��S����K?6��?���7!n�ߗ�<b��=3�^�b?UG4? �W���Ͼo��>1�\?�À?J[?�{�>[��w;��T濿�t��k`�<��K>��>=�>+���mK>��ԾO�C�傊>ְ�>�楼V3ھ=�������G�>7m!?���>JϮ=�� ?Ɣ#?<�j>�>nE��:����E�Ⱦ�>U��>@?��~?��?��o`3���+塿Ŏ[��KN>��x?c?��>Ś�������!N��!H�N��M��?�wg?�K�!?�3�?D�??E�A?��f>q}�� ؾ�t����>��!?C��v�A��C&�Ź�g�?�F?��>@����ս3�Լ����b����?y\?�9&?����a�D�¾���<�5&���M�(��;�*D���>�i>>A���ݴ=P�>��=>m��$6�S�g<��=Az�>��=�,7�m�2=,?=�G�uۃ���=k�r�BxD���>&JL>�����^?l=��{�����x���U��?���?Vk�?q��2�h��$=?�?>	?r"�>�J���}޾���Pw��}x��w�<�>��>O�l���F���ٙ���F���Ž��׽Ui�>C٦>�a?���>��>��>11��m��PcԾ����t^�w���a0���1��P�9��E��<p=\�ʾn}����>OH���?�>~?��G>��>��>YYn<�S�>8�b=�E>,G�>��>��>��=>��<���2�S?-�Ǿ�Z7�o0�����3�G?)�h?���>�|�O���U�N� ?KW�?'S�?SNi>�&r��#,��n? 2?O�l�8�	?�(=�4$=}:�=�ܣ��k=���7zY���>�꽳3E���L���J�m��>��?�Z�<f���F��6��69�Vc�?N�?��� UW�r�d�X�b�Cv��?	��8������o�>���|���`�����*4��{w�t~�>*eB?hH�z̪�rt��?G��Fp��_>	D�>��>�9�=�O�=�>��gy/��rJ�Q3 ��g5�I�?��?��>AG;?Qt6?�D?��Q?ت�>6�>7��=�> :�> Wd>$p�>�>N?+  ?�OJ?�d2?�B?�>{�i��뾎޾D?u�#?E?��?D��>�ӽ�䡁���=K��=�Ɠ��ʀ�׎"��@=Zy���`��ֹ='̞><`?W�0>�T%�>�X>�;?�d�>��>�Ŋ��}��D=E��>�\?+�>�A ��s�S��>��?�m��b$'=�/>d��=1��}*�;,P�=�r�f�=���c�e����<䝼=��X=������<�z�<Ӄ�:s�<u�>8�?���>�C�>�@��1� �a��f�=�Y>IS>�>�Eپ�}���$��p�g��]y>�w�?�z�?Ļf=��=��=}���U�����E���*��<�?<J#?)XT?]��?x�=?`j#?ҵ>+�iM���^�������?�",?ɍ�>
��ƽʾx��3���?O?{8a����B3)�No¾Q�Խ�>�^/�k4~�7���D��h��
���i��f��?���?$W@���6�a��Y���hk��X�C?��>L�>�>�)���g�}��;>�s�>R?p��>AT?�zt?��\?+�y>-2��Ъ�*^��5���� >`�D?���?�?�y? �>�%)>s$'�G����*�5����L�{���<ѐP>�0�>���>���>7>/�&�������㽄��=��t>�>^�>���>�m>;�*�V[G?��?�\���k��}S�輾��� ��?溝?r�:?��c>����T��I���D�>� �?��?�9?�ph�3��=4�g<�ø��kþ���>���>�f�>�w�=�0H;U��>t�>��>1����
�����˼���>�(?�*>�ſ9q�ԋm������C<!A��5f��|���F\�[��=�ՙ�����.��G�^�ܡ��ړ���Ŝ���z���>~&�=c�=��=Lw�<Pͼ���<�|M=�_�<��=�Ms�gSs<�'A���� ��韑��b<lM=-��2Ǿ�}?pKI?1�-?�C?��t>iL>T�B�u�>⤖�V�?{;Q>łh��5���>��&��s�����۾�gؾ�a�x���Ü>�O��>��6>Ю�=(�r<��=}ς=n+�=ѐ�}=P�=�M�=+ȧ=���=��>�d>�6w?����ڲ���4Q�)X��:?�8�>�~�=(�ƾ�@?%�>>�2������b�.?u��?�T�?_�?Ati��d�>1��䎽�n�=Ҷ��g>2>}��=��2����>��J>ă��J���|��^4�?|�@@�??�ዿϢϿ�a/>��7>�> �R�`�1��\�|b��{Z���!?�C;�eJ̾�9�>���=�(߾�ƾ'�.=��6>]b=�^�9Q\��=\{���;=�l=eԉ>��C>�c�=�)��%��=J{I=/��=��O>=P����7��+���3=��=L�b>��%>�	�>@?�"?ɰ??��?0��P���p�<�O8?
�D>���>�n<Ma>�?�H?�WR?�f?��>�����> ��>5���+W��l�����V����?�!�?��>�>Υ���C5�V^2�oc���?c+?8KG?)��>Yo�����<����鲆�h�B�lV;�l}��l������}���L�_F>!��>�7�>W�>�>q�A>j>�ϧ>��>�J�=A�>u�_�d� >c��=�k�=�ܤ�.�=+M>@Y=SP���}�{iE��>�<Z�o>MS�=����a��=	��>�6>1��>#��=���OF/>ļ��m�L����=jE���(B�O1d�2H~�w/�7_6���B>e<X>�m���3����?��Y>�u?>���?�@u?F�>��,�վ�N���Ee�4kS�o��=��>Y�<��q;��X`���M��xҾ���>o��>ŋd>E(>�{0���Vw�=`N��35�RA�>�R�Ce�=ꟽm�d�:����ڟ�Ta��!�=��??�K��N��=w$j?�.[?���?x+�>Bs�S�z���>P���ݝ��E=�#�}�B�<�?+�Z?@h�>m
�n�,���о�y��I�>{C��N��ٙ������0��᯾|�>:m���̾��S�]���<���P�����Tt�>qw]?L��?�&c�.���*�r��?���>�$?.�?`e�>��>��+?�j�� �������^�>L�X?읻?r@�?fv>���=�_�"��>8��>�??�e?\	4��[�>�I<v�/>�_��b�=3g>�=P�=�?�>r�
?=?�"��3���Ӿ:� �G�,��b�=�=p��'>�֯>�� >b� >j��=4Du=�C�>�`�>�߇>:@�>���>�>J��A�Bp?�� =,�>��W?��N>���<�<P�<�^Վ;Z���S�d�Q���ѽ�;史<�>��L< ��>݄ſX�?S8�>����?���.=����i><t�=Ϛ�����>Jn#>P��=!��>��>n��=�}@>�]-=��Ӿ��>�L��� ��C�T�R��Ҿ�@x>�8���Z'��������-J��$���z��i�h)����=�'��<~�?����p�j��*��t���?U��>��5?������=6>���>�f�>�����ƕ�o�����Ὰ�?L��?s>c>l�>U�W?i�?ۋ1�93��vZ���u�&A��	e�k�`�f��������
�u
����_?��x?tA?2�<9z>���?��%�`Ϗ�t+�>�/�*;��1<=�'�>�(����`��Ӿ��þ�/��8F>t�o?g#�?MU?�ZV���W���(>+:?�1?f�t?m�1?l;?#��o�#?ѨD>��?��
?Ig6?bH.?��?'�<>6��=De�y7=v���~狾{�ؽ߈��óμxF=�i=]�8A}�<�D�<��<�	�������<�x��Ű<7xD=f�=Y��=f��>�a`?���>��X>>:?.�:��g+�?)��R�8?9-�=z�O������$��X۾!�6>n)p?���?*?X?��Y>�=>�#�D��J>�{v>�5>	�o>~��>P��M�Y�v!�=���=�>K�>+���u���	�x������'3>���>�7|>@ō���'>?a���*z�z�d>��Q�Ҽ��D�S��G���1�iDv�I�>3�K?j�?[י=�Z����� ?f�))?rZ<?VM?��?���=O�۾�9���J����#�>X�<�����������:��؈:ٞs>���0���oT>��
�ѾU�g�ZL�A"���,��(%��>E		�s�о���g>�8�=TR�����<�������RD?��=����k�%� ����=���>��>����E�W�6�>��r��U��=]��>�h�=�PN����x�G��>��xN�>�G?�_?��?˴|��Fs�x�C��B ��/�������?\O�>��?�0>'��=��������e���G�n��>��>���F�%۞�-��f"�Z׉>�\?($'>Q�
?�LP?�	?��_?�&+?�?x̒>A������K&?n��?��=hԽgT�;�8���E���>(�)?^�B��ܗ>��?��?��&?�Q?b�?�>
� ��6@����>��>��W�hH��Q�_>�J?���>)Y?B̓?�=>>��5��f���֩�B��=~>+�2?�
#?��?�ϸ>�
?k�6���]�H�>#Dq?с?�ZN?~t/=�x?D�J>Z/?�Y6>�~>!?��1?7�f?	(�?�?��>Y�=[+��i~��6��<����=^���½�i��.�����;R߄=��9<����|�a�]�,Q��+.%��m��>P�>1t>k��^b0>��ľ2s���A>����ߛ�	�����:�\ŷ=��>��?�0�>��#�3Ɛ=���>"��>�����'?�?��?mDS; Hb�1C۾S�K��>zB?�N�=�l���P�u�sTk=�n?��^?�X����&�b?�]?�e�$	=�K�þl�b�}k龏�O?��
?��G��ų>�~?��q?S��>&f�q:n�����2b���j���=Bf�>Z�$�d��r�>0�7?;H�>O�b>���=�۾��w�\����?���?.��?���?�*>��n�.��Ͼ���V�X?B��>\Sp��%(?D���7ݾg�<�G���i��k����ɾN��������D8�5�Z������=#�?N�p?wj?���?Aw��{�]�r[d��_�>�K�4I�I{���/��+0�	�L�˝{���"��r���ξ���<�4���/�h��??�+@�B��>$�Ǿ�/��� �"j�>(��֌3���>��n=4�=<��=�={��9n�F5��?=&�>ަ�>R
6?qcA�j&2��5���&�����e��>�X�>��>+��>�>j�謚�����'žaY��D��~{|>- v?�RU?�%w?�����C�0��'��$�<�$�����=�uC=��3>|�d�P�<;+��h����X�����!$�=D�+?:�M> ��>��?m2�><Q��9�2
��D1����<`?Q_?A��>�ۦ>ᔽ����>ӽl?���>a�>����Q!���{��˽h�>�ŭ>��>h�o>��,�8\��j��6����9�l�=��h?f���ޏ`��Ӆ>�R?���:2�H<_V�>z�u���!����Ѭ'��j>p�?�"�=�g;>dDž��A�{��L��/yH?���>����P����>ٞC?���>/�7>��??��᾿e|>��?��V?��Q?ЈH?�?��˽<E��c+	�'-=�8I>� >��=��=Z��Ìo��C��8�<�C�;[r=�<ƽI�.=�)K=ay=�7=�l>zxڿtrK��׾_��0o�(
��^��󬿽DK��S)�ݵ�����7m��w�/c��R�G�e�2���$9t���?���?��/B���B��w�~��%��s&�>��t�q�P�q���U�k��c�����4��_M�k�f�TMg��9?;N����']�� a�],'?k:P?%n?q7�ƃ�����K>���<+n&>����\ɛ��Jп>�<N�?�K�>!̾x���>J=?�F�>n��=�0����޾���Ǹ>�F�>ڱv>R���ο�KĿ�'5>���?���?��B?8t'�F��^=���>[�
?�A>}�.���ce��t��>,�?�)�?��n=>mT��R޼�Uf?Y�;HE�S E;��=AB�=�z=����.O>-�>�!�\/9�p�½X�">�H�>��+��2���]�R�<�8Y>�P۽!��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=7�󿨪��������F<Ĭ��6�����DC�����^C}���i��ǥ=��o>`I�>�?>=�>zҪ=	��=��Q?��x?���>P�:>dڽUZ��8?Ӿ��>�D���������׋��Η�g���z8�;�美�	������W =��=�6R�S����� �R�b���F���.?ju$>��ʾ.�M��-<�mʾ���O����ߥ�.̾��1�?!n�-͟?��A?����	�V����O�$�����W?R����/묾���=�����=�$�>_��=	��< 3��}S��B0?a�?젾����S�*>@$��l#=�5+?��?{v[<��>��$?�k,�.�0,[>�g3>��>�b�>�J	>�q��t�ܽ��?U?U� ��������>�侾j�y���`=߂>�x4���^�X>4Ƅ<���� J�y���.�<,�U?�"�>�%�������bA��p-=��?2?I��>i��?@}/?b◻�Cľ��%�_�ؾ��
>�j?�c?��=�x���ݾ\�ɾ??�0h?��|>L�2 ��+�\�o?}��?��?�5_��_r� ������B?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>��������>5�v���?d{�?��Z����=�}��r��LپŽ�~�=�K�������	�b�D���վ�� ��]��a�;݉e>�@/���R\?�����׿�m˿�ۀ����&Q��$!?S6�>a$j�%-���9z�O�]��kN�l)H��?��JW�>%�>���ba�uә��F%��%>�C5?�|�%��>����K��F���:�����>S��>�e�=� ����N�|�?�W�i������;�Ԩ~?��?�(x?�$?G�{�s��5u�8�S=�@s?��?|�S?����w�CH>p�i?�^��<�x�+�R���k����>��?D�>7s־�3��p��hF?��>IY�G���οҔ����?d��?��_�?T��?^�9?��$�����-w�'d%��f�>�E"?Kv�<�Ჽ���GL�K��\�>�?4���
��.�_?��a�k�p�..��ɽݡ>��/��A[���������De��蛿3Vx���?KY�?Y��?�E�N�"��:%?e�>�͕���Ǿ���<�t�>nS�>r�N>�Z`���t>�=���:�vn	>P��?�w�?�?i���A���;>��}?Q$�>��?�o�=b�>�d�=N��-��j#>�"�=S�>��?s�M?�K�>�U�=�8�c/�-[F��GR�X$�&�C�>�>q�a?ӂL?kKb>���� 2��!��uͽ^c1�9S鼗W@���,��߽X(5>C�=>�>��D��Ӿ��?�n�L�ؿk���p'�V84?�>��?�����t��T�7_?v�>|.��*���'��FU�|��?AG�?y�?۷׾\�˼;>�>�M�>��Խ���n��g�7>ĜB?#�^@��?�o�Q�>���?��@֮?��h��	?���P��Ua~����7�i��=��7?�0��z>���>��=�nv�ݻ��W�s����>�B�?�{�?��>!�l?��o�N�B�x�1=8M�>Μk?�s?�Qo���m�B>��?!������L��f?�
@u@`�^?*�¿^��� J��xz���l>�}�=(n�=�%���5��Ȅ�<���=w���bY<��{>� �=���>�#>ϊ>�>�:����%�Oe���4���6���6=&��'�I�7�U����8	�:A������]K�ڃL��X���(�z�&ט���>=Pf?4D[?��p?&�?��-y�=�{�r>'c���>M+V>�?��=?��3?�MZ>��̽$ s�#��귕�µ�(a>K!=C�>�r?a�>�-�=\/�>d�&>�
�>rx>��>�;>��=�b >�;�>���>P��>Q�>>A>Ƿ��"˱�p�j�T�t��W���u�?u����	J������l���������=�w/?a�>k@���8Ͽ�Ӭ�B)H?Ԙ������+��	>"1?�aW?��>+\���)y�6>u��Kn��>P�����k�Ir+��P>�?��e>�t>�a3�\@8�ʮP�S����j{>�5?PA����7�Țu�<�H�˅ܾ��M>���>��?��^�J얿>,���h��4=�:?�?�K���尾�&v�VN��M�Q>�']>c=և�==�M>�d���Ƚ�G�H-=X��=��]>^�?o�>��=%"�>>.��R���>�0>��=>�g9?�y)?��Q��ϽP��(F#�ap>��>7~>S2>J9��d�=��>���>�j��i�����$�&OV�~�Y>^4c�cq^��M��U�=佮)�=ZF�<,1�cfW����<��~?�~���䈿g�8y���lD?8-?�	�=3?F<~�"�L����E��(�?��@kl�?��	��V� �?%A�?������=�z�>Uث>�ξ��L�C�?ƽ�Ƣ��	��'#��R�?
�?
�/��ɋ�ml�2>X_%?H�Ӿr�>;�g_�����-�u�\.$=߻�>�6H?�]��x�O��>�Gt
?4?xG�W���s�ȿ�}v����>��?�?��m�N<��\@�uz�>��?�eY?Fi>�U۾qzZ�]��>[�@?�R?�>8�*�'�F�?�ݶ?���?e:b>L��?uct?tV1?�A>`A$�J���#������=6���%�s>���<��¾�?��PJ��L�$�B�>�U�/�3��<�һa�>�뗻T���	y�<�����ჾ5��;K7�>���>�;=�9�>X7�>��^>���>�0�>̨�:ᚗ�2=����K?H��?2��*0n�T��<ʬ�=�^��$?ZJ4?D[���Ͼeը>��\?N?H[?�f�>���=���翿a|��ҩ�<��K>4�>D�>5,��eFK>��Ծs+D�Fq�>ϗ>�����>ھ�*��"���|B�>�f!?M��>!Ʈ=��?�y"?��z>�O�>��F�̒��jF�b��>�"�>~/?��~?ɛ?X񱾃!8��Ғ��m����X��L>H�u?��?0'�>�F៿�sO��c�� |��g�?�Mn?�gٽCz?�C�?�E??<6C?xG{>���Ծ|ʉ�^V�>�!?���ʎA��%�����=	?�V?�%�>����LYڽ��ؼ��[���w?3_[?��%?���`�\�����<�Ia�}Tź<O�;l�1���>"">���"��=T�>s��=�l�Y9��}L<�@�=�!�>���=c7��A��(=,?�G�Rۃ���=f�r�xD���>�IL>�����^?�k=��{�����x��	U�� �?��?Lk�?$��%�h��$=?�?~	?x"�>K��
~޾N�ྷPw�8~x��w�X�>���>1�l���L���̙���F��d�Ž�����} ?��>��>��>���>X�>9��l��Cb������d��G�����2�������U��v��=k�������͆>�9��I��>�.?0N>۫u>4�>�%���>a*�=@��=���>�ň>%�>��>>B��
�I��%R?����-�ih���о��??�xl?���>O���u��������?#��?�{�?bܑ>.d��Y3��z?h�?��l����>iE���L<�H{==���8��;f����*e>��Խ��5��S�3�T��8?�?1���u�ž�⢽�u����=���?�/?�2!���w�����:�#���cM>�����Ӿp�=��~|�ar��a:k�Gsp�g�=���X?"_?�9e���賩��P�������>`=�>'�>���>yc�=����O�cC���O�(��`�>��?&�>![I?��9?�aN?�VN? M�>7j�>z��a?�ץ<���>F��>��;?��/?7p0?f�?��0?@>oC!����XԾ�?�?��?J��>���>�>����m���A;ֻ�9S�m�h�*���='s�;�,���������=O�=>�d?S���8������j>�7?��>Ӫ�>I���*���k�<a��>��
?$o�>� ���r��o�ı�>�?3%�o�=�F*>;��=��Ā�����=�iż`T�=����D
;��@$<�=5��=���#!X�� ;:Y�;uΰ<�t�>-�?���>�C�>�@��#� �]���e�=�Y>7S>�>�Eپ�}���$��m�g��]y>�w�?�z�?޻f=��=ז�=�|��`U�����O�����<�?;J#?!XT?Y��?u�=?[j#?��>+�jM���^�������?",?���>
����ʾ��p�3�,�?�X?�<a�K��;)��¾S�Խ�>�\/��1~���`D�w�������y�����?H��?�+A���6��s�'����R����C?& �>�Z�>��>^�)�+�g�]&��8;>��>R?$S�>�W?�~?�8b?Cr_>��>�PB���*��X�;��$>�w9?�2o?:��?/�l?���>�9>;T������l��3R�smv��qE=�W>R̚>��>�ҩ>�d�=혽*�6��'���=��>}��>��>���>�N�>G�(��kF?�Q?׾�������Z�ؾViw�z��?�(�?Tp?�~�>nT���V���?�ө?dR�?��U?(�^��I>�e#=���d6Ҿm�>�ف>Tɍ>��>���K�>6��>���>|+�����e���@��>��I?��>�Mѿ��;�I�U�(��'>TΌ����,�>��¾�n=�Q�T������
�i�k�`���k�a�������p�>���=.�	>iԈ> S����n=l�>�
���L.=5A�=�5)���ݽ� >~Bl=��;�����f�=Ӕ�=pʽ��˾��}?<I?G�+?1�C?#�y>�6>��3�<��>����@?�V>��P�����lz;�W������ �ؾ�|׾��c�"͟��C>�wI�|�>�E3>S�=8k�<B%�=�s=�Ҏ=�O�:3=C.�=�X�=�c�=���=��>�Q>�6w?W�������4Q��Z罤�:?�8�>q{�=��ƾq@?��>>�2������xb��-?���?�T�??�??ti��d�>M���㎽�q�=F����=2>t��=u�2�S��>��J>���K��;����4�?��@��??�ዿТϿ:a/>�7>_>x�R�M�1���\�I�b�YtZ���!?�C;�E̾D4�>��=))߾V�ƾɰ.=��6>�b=�h��R\����=�{�@�;=�l=�҉>�C>�l�={D��m�=|�I=��=C�O>���m�7�^5,�$�3=x��=ҩb>d&>s� ?�� ?�?ɧR?�}�>�j��=썾�z����?�5>��?�M>�2C>3r?J�??�XY?��?�I�>]!D����>IA�>w)�V+2������>�<�?���?�X�>�E��'��O��!�7g�<,��>�� ?ŧ5?\�>>�S|࿨�K��,���G����<����z(��L�c-8�0 ��a�>�v�>���>E�>G�!>&>,=:>���>�>��l<L�8�V+��_s��,)�!�Y��n׼:E=&�%>3bM>\��>�D�=���=&��;D-��d���:	M�=���>��>�}�>}e�=We���1>������J��ø=�%���@��'b��{���/�ӌ>��;>��Z>"Y_�ڑ��Y?)jS>�B>2s�?]�v?CG>����־ҹ���Hb�V�d�lm�=g>?�<���6�?�^�óM�/Ծ���>o%�>({�>�+<>��:��a-�">=���������>ƾ�9�=��?���Z�k�������c��k�=a+[?.�����4>�gS?��N?�-�?���>�D�q^�I�<�������=.KW��Rн��)>��>|kI?b��><���M���ƾμ���i�>��N��M�������?�O-�<��߾�h�>���7�Ծ����_��D<���bH��,{��4�>1GA?l��?DX��䄿gX`�����&�;,p?I�q?���>N�?��?RK�����g�)�>�a?vu�?���?4V>^��=r���>�5?Ί�?�ܓ?N�n?T8���>�[V��>�<�uԭ=�/(>K�=3y�=�'
?,�?�r	?�pK�W����u��W�0{=��=�9�>�>볐>��=���=6�3=�O3>m��>�k�>��>xi�>��>����?����X?�B�=���>QfK?\��>6_(=gԼ���'oI<��t��$��P(�I���:=�y����y=ջ<P�>�ſ�?C�U>p��#��>n�Э��wt>hJ�>]n�=~W�>G>���=�̵>4�>���>�>i>:>q=^JӾ��>@���H!��$C�śR� Ҿ�8z>�����[%�8��&.��>pH�ߠ���}��j�?'���@=�ĥ�<�;�?na����k���)�`�� y?�G�>�$6?���∽�>���>���>�q������>ȍ��:���?���?�?c>�E�>��W?��?D51�F?3�K{Z��u��A��e��`��Ӎ�Ӗ��.�
������_?��x?�NA?�9�<�z>Ԡ�?��%��֏�0�>c /�;�V_<=�4�>� ��e5a���Ӿ=�þvT���F>�o?��?�2?X�V�B�r9>��8?^�0?'�t?3�3?'6?̷�5'?5'8>Լ?�n	?g�7?�/?�?��K>A�>��˼�`.<~O���"��Ӕɽ�E����!�AC=[G�=7/���7�<�Pf=�� =HR����ѻ��O<O�&V�<o)�=��=h��=��>'^?���>��>��7?	z���8�S���to/?��&=>����u��\�����򾤟>٠k?�m�?:�W?�\]>��@�2�A�E�>�щ>u�">�W>��>��뽿$E�y��=>�T>�'�=3�'��L~��	����$
�<kf>���>�{>؆����'>;W����y���d>�R������S���G���1���v�#6�>�K?��?���=D������+f�&)?!f<?�tM?��?,Q�==�۾#�9���J�-R�$�>��<���<���h ����:����:�&s>4/�� Xξ��=�依ӑ�[l\��Ma��b���]�$&�,���>������R����>�>����S�!��c���"���"O?��=`�N����Ƞ���j	>n�>1J�>(� �� ��u>������W�	�>�C��U��P�ͫT��l�>�|T?�TU?���?-T�>�a�+U�Z���3���"��?C�q>Z^�>S�d>�>Mܚ��(��Fk�%�O�F'�>b�>}��kg:��奾����	�yt�>�8 ?��>�<?uJY?��?4j?�+?�m�>`Ʀ>�˽�c˾�%?�_�?;3�=�ѽQ�9�I4�6S?�ڍ�>��)?�x(����>�?��?��)?��R?�^?��>[���C��X�>2��>;�S��ܮ��L`>.�E?���>W?檆?rxF>E+4�L���5X���-�=eP*>�0?ڒ$?�?�W�>���>�x���=�7	?¹m?ʵ{?��b?!n�=[j�>�V�>�ٳ>�Y`=8&�>���>*2?�Td?��?��/?F�?g�=�	�<�Y�'q	<��<��=�W���=���=ՠ����.=��<�ޔ����=���;��<����b�<Bk��6t�>N,t>�!��Ja0>�žX���GBA>���Ge��;Ԋ�#�9�ٶ�=���>B�?Oܔ>^i$�W.�=�ȼ>�o�>�����'?��?�D?}��;W;b��۾JNJ��>�B?���='!m��c��5�u��Kj=Yn?�%^?�X�����=�b?��]?7h��=���þŵb�r���O?
�
?#�G���>��~?G�q?��>��e�%:n����Cb�k�j��϶=)r�>(X��d�4@�>w�7?}N�>�b>�%�=u۾��w�Zr��@?w�?�?���?�**>~�n�,4࿵���k����M?L��>�ń�[k8?~��!��"��澹�����Jv�D_��$��Ͼ{�GA��R����½��=�#?�}?L�g?�vo?�(پĦ��	NI��i��\�ď
��0��4���:�3I�:�R��1پ�� ��;���/z�uXB�P��?��&?�-��Y�>�#��:���žR
4>�s��J��`I�=�N���nG=��_=�g� �,��B��E?�y�>���>��>?6Y�i@�)�/��.5��-��JF*>���>r��>���>67����(���нQ Ѿ�V��K���>�f?aTH?- v?87�6�"�����q!�����4�����.>a�=��?>r�O�[�����z�B���s���p���"���<��?Dҍ>���>��?�+�>���4o���YC���*��9�B$�>{Jw?ڽ�>��>�Zҽ[� ����>@�l?@�>�v�>�B��!��~{��aͽ���>9j�>��>{�q> ,��\�n��i���}9�y�=�h?oǄ�al`�\�>AGR?M�6;�Q;<���>A�x���!�=J��'��>@?���=�;>n�ľ]G���{�1u��v*-?��*?�$ٽ�s/���>kT�> %?g�>?j�?9�(?ҾS�ܽ�}/?�dt?�k?[?W�2?'����ҽ�ǽ�؆�^�=�F�>Ķ�=Ԝ#>	��=������پ?V���6��(��=j�T>�r ����<�뫼��=�tS�-�>lۿuZ�QξԃȾY��D����� ?�6����)�+��.̛��r<�C������;�	K�f�:�`�M����S�?,�?�+���T9����������K>��w>�ކ����g�˾�h�����ǆþe���Ȥ2�Vx�����z.���^*?H9���̿5 ��q����%?�,?2)�?�y����d��Hf>���=�軞�y��'̿ m�4f?���>2��F+����>K��>2�>�)G>TI��+7����<I?I�?�>��.��Yÿ�^���Y=���?�/@��A?�^(�&z��>7="'�>?T�C>Q.�`������>���?�ފ?��G=wdW����3+e?ч�<��D��6޻v?�=w�=�h=�~�a�J>�ϓ>���	�>�Y�཈�.>G�>�^�w���)_��.�<�v\> �ؽ��2Մ?{\�sf���/��T���T>��T?6+�>S;�=��,?97H�W}Ͽ��\��*a?�0�?��?+�(?)ۿ��ؚ>��ܾ{�M?YD6?���>�d&���t�S��=U4Ἵ���h���&V�6��=���>��>Ղ,���̇O��M��N��=�����̿�+����߆$<�<�Vͼ���Pp$���s�~�������U��S�=�`�=Q�u>B!�>�Jr>$�>>�WZ?5�y?.��>Xa+>6�K⟾V���'�C�0r|��� �	�5��o �Cȕ���2�ξ{-��n$����H��)#=�Bҍ=�/R�g���r� �g�b��F���.?;M$>��ʾe�M�
�-<�eʾA����؄�8᥽�1̾Q�1�4)n�.̟?��A?G���V����`:�Xr����W?�c�߼�gV��=���Af=�	�> s�=h��s"3�}S��0?�?���\����0>����$=�,?yb?��<�*�>�v#?+�'�9eֽ�Wc>�;>��>:�>��>�����߽E�?�LS?�������f�>�\��}1~�@�l=���=�"6����t\>8�<E���7Ӧ��.���y�<�V?ꌛ>�!&�7&#���x� p|�O2�=Ħ|?+�?/��>
�m?��9?�Z�<��޾q�B��J��1��=яU?�A`?�� >�}��1Iɾ?R��c�4?te?=�h>~�Q�Bz��%�5��b?��w?��?J߾� t}����t�� b3?'�v?\r^��s�������V�$@�>2]�>���>��9�mk�>_�>?#��F��e���dY4����?8�@���?*<<��E��=�;?"Y�>�O�H=ƾQu�����ҙq=� �>����2cv���3V,�V�8?Ƞ�?���>Z���5��խ>Z�j�m%�?��?Q����7<�X���_����-�s`�=S�#�%���C<�U�&�$צ�:���%��r�d�猁>w@��:���>��69��Ͽe�~�,Yݾ���Z�?a�>��(׉���u��^i�R=G�RnO��窾�r�>z>b���$V�����!jC��=f��>t꛼<u> XT����������{�<'c>C�>�Z>Q8��/����?�Z���ۿp�����/��f?$�?�?5+?���<b�%�.X���>�R?��?�K?�c���/�E ���u?��N�ȯ���Vr��q{��0?wRW?���>�ܾ{n���@�>vu%?fȥ>s&��ث�C>��^֝�Bϴ?��?�ݾ�?F�?5X?`����@����W���#�ȹ�>9�<;�.�P����.�:Pپ�>�>6j�>�m��8 �3�_?c�a���p���-���ƽPס>$�0�Z\��������Ue�b���?y�Q��?�]�?V�?!���"��4%?Y�>����#7Ǿ��<���>�*�>a0N>%4_�ӫu>�y�:�|e	>���?�}�?i?������E>��}?�&�>A�?�~�=}e�>�a�=���.� U#>�=�N?�#�?1�M?B�>�4�=0�8�r/�\F��ER� #���C���>��a?c�L?�^b>�+��~~2��!���ͽ X1��B��_@�8�,��v߽o5>/�=>�>��D� Ӿ�C.?���+U������W��x0K?<~�>�u	?|�Ӿ��]���#>q�6?Wܰ>�M�pv���b����ʽ�m�?s��?ޏ�>�o��2�<p]�=�é>���>�H�p[J�	����4>??�1��ف�@�f�D$>�?i@+Y�?�XW��	?���P��\a~���*7����=��7?�0��z>��>v�=�nv�ѻ��R�s�t��>�B�?�{�?3��>�l?x�o�<�B���1=M�>Ȝk?�s?3Yo�u�a�B>y�?������L��f?	�
@zu@N�^?\%տ� ��龱���pe=F�U;$�=M�-�Hd<0���+��e=^���(>���>i��>��>�f4>`�>� >�Z���(�С����w���6� $�D�H�@XB�����.��΀��4-��Wv@=�9E��@*�*�����%�VeT��k9>~O^?�@?#?j?�n?��q���N=m^�;k	�e�(�e�>p?� ?PCX?Z+?oE->4�^�|Fr�C6��W+�������>�ʹ<��>���>��?��=g�>n��>��M>��v>'��=ke�=Mj�= ��>��?�b�>5�t>�C<>��>Dϴ��1��j�h��
w��̽/�?����S�J��1���9��Ԧ���h�=Fb.?|>���?пg����2H?!���w)���+���>~�0?�cW?�>!����T�.:><����j�-`>�+ ��l���)��%Q>wl?۷f>�u>�3��c8���P�v}���\|>�06?���L9�c�u�_�H��hݾDM>��>�FD�[m�������%ui��{=Sy:?\�?�0��<߰���u��B���TR>�5\>�*=�S�=�JM>��c�-�ƽ�H��[.=��=%�^>��?A~ >��=�*�>�ҵ9�G*�><�A>a5>�$<?�$?/x��tC��������)�$Dv>-��>I��>>]FF���=eD�>�o>��
�!������<���R>���s�_�2p��o=G���g�=x<�=[��COH��A
=�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>��P�Ko��f$��E0��*ހ=Y?��|?}9��-$R�,P�<{o5?�e?�E��@���Ŀ�s��?���?	�?�xn�)���0�y��>��?:mX?�ԏ>�1��,�<����>)C?S��?�?uľW���"[�>v��?��v?~�>���?�^k?A�?5��=8F��������ѯ<L�R�'_x>{ݻ<�T��7���{�
�Z��^p���+��"d=-:=H}�>�a��`���o=>���ny��\���9U>���>e�P>�<b><��>��?�>�2I���˼�T��S����K?6��?���7!n�ߗ�<b��=3�^�b?UG4? �W���Ͼo��>1�\?�À?J[?�{�>[��w;��T濿�t��k`�<��K>��>=�>+���mK>��ԾO�C�傊>ְ�>�楼V3ھ=�������G�>7m!?���>JϮ=�� ?Ɣ#?<�j>�>nE��:����E�Ⱦ�>U��>@?��~?��?��o`3���+塿Ŏ[��KN>��x?c?��>Ś�������!N��!H�N��M��?�wg?�K�!?�3�?D�??E�A?��f>q}�� ؾ�t����>��!?C��v�A��C&�Ź�g�?�F?��>@����ս3�Լ����b����?y\?�9&?����a�D�¾���<�5&���M�(��;�*D���>�i>>A���ݴ=P�>��=>m��$6�S�g<��=Az�>��=�,7�m�2=,?=�G�uۃ���=k�r�BxD���>&JL>�����^?l=��{�����x���U��?���?Vk�?q��2�h��$=?�?>	?r"�>�J���}޾���Pw��}x��w�<�>��>O�l���F���ٙ���F���Ž��׽Ui�>C٦>�a?���>��>��>11��m��PcԾ����t^�w���a0���1��P�9��E��<p=\�ʾn}����>OH���?�>~?��G>��>��>YYn<�S�>8�b=�E>,G�>��>��>��=>��<���2�S?-�Ǿ�Z7�o0�����3�G?)�h?���>�|�O���U�N� ?KW�?'S�?SNi>�&r��#,��n? 2?O�l�8�	?�(=�4$=}:�=�ܣ��k=���7zY���>�꽳3E���L���J�m��>��?�Z�<f���F��6��69�Vc�?N�?��� UW�r�d�X�b�Cv��?	��8������o�>���|���`�����*4��{w�t~�>*eB?hH�z̪�rt��?G��Fp��_>	D�>��>�9�=�O�=�>��gy/��rJ�Q3 ��g5�I�?��?��>AG;?Qt6?�D?��Q?ت�>6�>7��=�> :�> Wd>$p�>�>N?+  ?�OJ?�d2?�B?�>{�i��뾎޾D?u�#?E?��?D��>�ӽ�䡁���=K��=�Ɠ��ʀ�׎"��@=Zy���`��ֹ='̞><`?W�0>�T%�>�X>�;?�d�>��>�Ŋ��}��D=E��>�\?+�>�A ��s�S��>��?�m��b$'=�/>d��=1��}*�;,P�=�r�f�=���c�e����<䝼=��X=������<�z�<Ӄ�:s�<u�>8�?���>�C�>�@��1� �a��f�=�Y>IS>�>�Eپ�}���$��p�g��]y>�w�?�z�?Ļf=��=��=}���U�����E���*��<�?<J#?)XT?]��?x�=?`j#?ҵ>+�iM���^�������?�",?ɍ�>
��ƽʾx��3���?O?{8a����B3)�No¾Q�Խ�>�^/�k4~�7���D��h��
���i��f��?���?$W@���6�a��Y���hk��X�C?��>L�>�>�)���g�}��;>�s�>R?p��>AT?�zt?��\?+�y>-2��Ъ�*^��5���� >`�D?���?�?�y? �>�%)>s$'�G����*�5����L�{���<ѐP>�0�>���>���>7>/�&�������㽄��=��t>�>^�>���>�m>;�*�V[G?��?�\���k��}S�輾��� ��?溝?r�:?��c>����T��I���D�>� �?��?�9?�ph�3��=4�g<�ø��kþ���>���>�f�>�w�=�0H;U��>t�>��>1����
�����˼���>�(?�*>�ſ9q�ԋm������C<!A��5f��|���F\�[��=�ՙ�����.��G�^�ܡ��ړ���Ŝ���z���>~&�=c�=��=Lw�<Pͼ���<�|M=�_�<��=�Ms�gSs<�'A���� ��韑��b<lM=-��2Ǿ�}?pKI?1�-?�C?��t>iL>T�B�u�>⤖�V�?{;Q>łh��5���>��&��s�����۾�gؾ�a�x���Ü>�O��>��6>Ю�=(�r<��=}ς=n+�=ѐ�}=P�=�M�=+ȧ=���=��>�d>�6w?����ڲ���4Q�)X��:?�8�>�~�=(�ƾ�@?%�>>�2������b�.?u��?�T�?_�?Ati��d�>1��䎽�n�=Ҷ��g>2>}��=��2����>��J>ă��J���|��^4�?|�@@�??�ዿϢϿ�a/>��7>�> �R�`�1��\�|b��{Z���!?�C;�eJ̾�9�>���=�(߾�ƾ'�.=��6>]b=�^�9Q\��=\{���;=�l=eԉ>��C>�c�=�)��%��=J{I=/��=��O>=P����7��+���3=��=L�b>��%>�	�>@?�"?ɰ??��?0��P���p�<�O8?
�D>���>�n<Ma>�?�H?�WR?�f?��>�����> ��>5���+W��l�����V����?�!�?��>�>Υ���C5�V^2�oc���?c+?8KG?)��>Yo�����<����鲆�h�B�lV;�l}��l������}���L�_F>!��>�7�>W�>�>q�A>j>�ϧ>��>�J�=A�>u�_�d� >c��=�k�=�ܤ�.�=+M>@Y=SP���}�{iE��>�<Z�o>MS�=����a��=	��>�6>1��>#��=���OF/>ļ��m�L����=jE���(B�O1d�2H~�w/�7_6���B>e<X>�m���3����?��Y>�u?>���?�@u?F�>��,�վ�N���Ee�4kS�o��=��>Y�<��q;��X`���M��xҾ���>o��>ŋd>E(>�{0���Vw�=`N��35�RA�>�R�Ce�=ꟽm�d�:����ڟ�Ta��!�=��??�K��N��=w$j?�.[?���?x+�>Bs�S�z���>P���ݝ��E=�#�}�B�<�?+�Z?@h�>m
�n�,���о�y��I�>{C��N��ٙ������0��᯾|�>:m���̾��S�]���<���P�����Tt�>qw]?L��?�&c�.���*�r��?���>�$?.�?`e�>��>��+?�j�� �������^�>L�X?읻?r@�?fv>���=�_�"��>8��>�??�e?\	4��[�>�I<v�/>�_��b�=3g>�=P�=�?�>r�
?=?�"��3���Ӿ:� �G�,��b�=�=p��'>�֯>�� >b� >j��=4Du=�C�>�`�>�߇>:@�>���>�>J��A�Bp?�� =,�>��W?��N>���<�<P�<�^Վ;Z���S�d�Q���ѽ�;史<�>��L< ��>݄ſX�?S8�>����?���.=����i><t�=Ϛ�����>Jn#>P��=!��>��>n��=�}@>�]-=��Ӿ��>�L��� ��C�T�R��Ҿ�@x>�8���Z'��������-J��$���z��i�h)����=�'��<~�?����p�j��*��t���?U��>��5?������=6>���>�f�>�����ƕ�o�����Ὰ�?L��?s>c>l�>U�W?i�?ۋ1�93��vZ���u�&A��	e�k�`�f��������
�u
����_?��x?tA?2�<9z>���?��%�`Ϗ�t+�>�/�*;��1<=�'�>�(����`��Ӿ��þ�/��8F>t�o?g#�?MU?�ZV���W���(>+:?�1?f�t?m�1?l;?#��o�#?ѨD>��?��
?Ig6?bH.?��?'�<>6��=De�y7=v���~狾{�ؽ߈��óμxF=�i=]�8A}�<�D�<��<�	�������<�x��Ű<7xD=f�=Y��=f��>�a`?���>��X>>:?.�:��g+�?)��R�8?9-�=z�O������$��X۾!�6>n)p?���?*?X?��Y>�=>�#�D��J>�{v>�5>	�o>~��>P��M�Y�v!�=���=�>K�>+���u���	�x������'3>���>�7|>@ō���'>?a���*z�z�d>��Q�Ҽ��D�S��G���1�iDv�I�>3�K?j�?[י=�Z����� ?f�))?rZ<?VM?��?���=O�۾�9���J����#�>X�<�����������:��؈:ٞs>���0���oT>��
�ѾU�g�ZL�A"���,��(%��>E		�s�о���g>�8�=TR�����<�������RD?��=����k�%� ����=���>��>����E�W�6�>��r��U��=]��>�h�=�PN����x�G��>��xN�>�G?�_?��?˴|��Fs�x�C��B ��/�������?\O�>��?�0>'��=��������e���G�n��>��>���F�%۞�-��f"�Z׉>�\?($'>Q�
?�LP?�	?��_?�&+?�?x̒>A������K&?n��?��=hԽgT�;�8���E���>(�)?^�B��ܗ>��?��?��&?�Q?b�?�>
� ��6@����>��>��W�hH��Q�_>�J?���>)Y?B̓?�=>>��5��f���֩�B��=~>+�2?�
#?��?�ϸ>�
?k�6���]�H�>#Dq?с?�ZN?~t/=�x?D�J>Z/?�Y6>�~>!?��1?7�f?	(�?�?��>Y�=[+��i~��6��<����=^���½�i��.�����;R߄=��9<����|�a�]�,Q��+.%��m��>P�>1t>k��^b0>��ľ2s���A>����ߛ�	�����:�\ŷ=��>��?�0�>��#�3Ɛ=���>"��>�����'?�?��?mDS; Hb�1C۾S�K��>zB?�N�=�l���P�u�sTk=�n?��^?�X����&�b?�]?�e�$	=�K�þl�b�}k龏�O?��
?��G��ų>�~?��q?S��>&f�q:n�����2b���j���=Bf�>Z�$�d��r�>0�7?;H�>O�b>���=�۾��w�\����?���?.��?���?�*>��n�.��Ͼ���V�X?B��>\Sp��%(?D���7ݾg�<�G���i��k����ɾN��������D8�5�Z������=#�?N�p?wj?���?Aw��{�]�r[d��_�>�K�4I�I{���/��+0�	�L�˝{���"��r���ξ���<�4���/�h��??�+@�B��>$�Ǿ�/��� �"j�>(��֌3���>��n=4�=<��=�={��9n�F5��?=&�>ަ�>R
6?qcA�j&2��5���&�����e��>�X�>��>+��>�>j�謚�����'žaY��D��~{|>- v?�RU?�%w?�����C�0��'��$�<�$�����=�uC=��3>|�d�P�<;+��h����X�����!$�=D�+?:�M> ��>��?m2�><Q��9�2
��D1����<`?Q_?A��>�ۦ>ᔽ����>ӽl?���>a�>����Q!���{��˽h�>�ŭ>��>h�o>��,�8\��j��6����9�l�=��h?f���ޏ`��Ӆ>�R?���:2�H<_V�>z�u���!����Ѭ'��j>p�?�"�=�g;>dDž��A�{��L��/yH?���>����P����>ٞC?���>/�7>��??��᾿e|>��?��V?��Q?ЈH?�?��˽<E��c+	�'-=�8I>� >��=��=Z��Ìo��C��8�<�C�;[r=�<ƽI�.=�)K=ay=�7=�l>zxڿtrK��׾_��0o�(
��^��󬿽DK��S)�ݵ�����7m��w�/c��R�G�e�2���$9t���?���?��/B���B��w�~��%��s&�>��t�q�P�q���U�k��c�����4��_M�k�f�TMg��9?;N����']�� a�],'?k:P?%n?q7�ƃ�����K>���<+n&>����\ɛ��Jп>�<N�?�K�>!̾x���>J=?�F�>n��=�0����޾���Ǹ>�F�>ڱv>R���ο�KĿ�'5>���?���?��B?8t'�F��^=���>[�
?�A>}�.���ce��t��>,�?�)�?��n=>mT��R޼�Uf?Y�;HE�S E;��=AB�=�z=����.O>-�>�!�\/9�p�½X�">�H�>��+��2���]�R�<�8Y>�P۽!��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=7�󿨪��������F<Ĭ��6�����DC�����^C}���i��ǥ=��o>`I�>�?>=�>zҪ=	��=��Q?��x?���>P�:>dڽUZ��8?Ӿ��>�D���������׋��Η�g���z8�;�美�	������W =��=�6R�S����� �R�b���F���.?ju$>��ʾ.�M��-<�mʾ���O����ߥ�.̾��1�?!n�-͟?��A?����	�V����O�$�����W?R����/묾���=�����=�$�>_��=	��< 3��}S��B0?a�?젾����S�*>@$��l#=�5+?��?{v[<��>��$?�k,�.�0,[>�g3>��>�b�>�J	>�q��t�ܽ��?U?U� ��������>�侾j�y���`=߂>�x4���^�X>4Ƅ<���� J�y���.�<,�U?�"�>�%�������bA��p-=��?2?I��>i��?@}/?b◻�Cľ��%�_�ؾ��
>�j?�c?��=�x���ݾ\�ɾ??�0h?��|>L�2 ��+�\�o?}��?��?�5_��_r� ������B?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>��������>5�v���?d{�?��Z����=�}��r��LپŽ�~�=�K�������	�b�D���վ�� ��]��a�;݉e>�@/���R\?�����׿�m˿�ۀ����&Q��$!?S6�>a$j�%-���9z�O�]��kN�l)H��?��JW�>%�>���ba�uә��F%��%>�C5?�|�%��>����K��F���:�����>S��>�e�=� ����N�|�?�W�i������;�Ԩ~?��?�(x?�$?G�{�s��5u�8�S=�@s?��?|�S?����w�CH>p�i?�^��<�x�+�R���k����>��?D�>7s־�3��p��hF?��>IY�G���οҔ����?d��?��_�?T��?^�9?��$�����-w�'d%��f�>�E"?Kv�<�Ჽ���GL�K��\�>�?4���
��.�_?��a�k�p�..��ɽݡ>��/��A[���������De��蛿3Vx���?KY�?Y��?�E�N�"��:%?e�>�͕���Ǿ���<�t�>nS�>r�N>�Z`���t>�=���:�vn	>P��?�w�?�?i���A���;>��}?Q$�>��?�o�=b�>�d�=N��-��j#>�"�=S�>��?s�M?�K�>�U�=�8�c/�-[F��GR�X$�&�C�>�>q�a?ӂL?kKb>���� 2��!��uͽ^c1�9S鼗W@���,��߽X(5>C�=>�>��D��Ӿ��?�n�L�ؿk���p'�V84?�>��?�����t��T�7_?v�>|.��*���'��FU�|��?AG�?y�?۷׾\�˼;>�>�M�>��Խ���n��g�7>ĜB?#�^@��?�o�Q�>���?��@֮?��h��	?���P��Ua~����7�i��=��7?�0��z>���>��=�nv�ݻ��W�s����>�B�?�{�?��>!�l?��o�N�B�x�1=8M�>Μk?�s?�Qo���m�B>��?!������L��f?�
@u@`�^?*�¿^��� J��xz���l>�}�=(n�=�%���5��Ȅ�<���=w���bY<��{>� �=���>�#>ϊ>�>�:����%�Oe���4���6���6=&��'�I�7�U����8	�:A������]K�ڃL��X���(�z�&ט���>=Pf?4D[?��p?&�?��-y�=�{�r>'c���>M+V>�?��=?��3?�MZ>��̽$ s�#��귕�µ�(a>K!=C�>�r?a�>�-�=\/�>d�&>�
�>rx>��>�;>��=�b >�;�>���>P��>Q�>>A>Ƿ��"˱�p�j�T�t��W���u�?u����	J������l���������=�w/?a�>k@���8Ͽ�Ӭ�B)H?Ԙ������+��	>"1?�aW?��>+\���)y�6>u��Kn��>P�����k�Ir+��P>�?��e>�t>�a3�\@8�ʮP�S����j{>�5?PA����7�Țu�<�H�˅ܾ��M>���>��?��^�J얿>,���h��4=�:?�?�K���尾�&v�VN��M�Q>�']>c=և�==�M>�d���Ƚ�G�H-=X��=��]>^�?o�>��=%"�>>.��R���>�0>��=>�g9?�y)?��Q��ϽP��(F#�ap>��>7~>S2>J9��d�=��>���>�j��i�����$�&OV�~�Y>^4c�cq^��M��U�=佮)�=ZF�<,1�cfW����<��~?�~���䈿g�8y���lD?8-?�	�=3?F<~�"�L����E��(�?��@kl�?��	��V� �?%A�?������=�z�>Uث>�ξ��L�C�?ƽ�Ƣ��	��'#��R�?
�?
�/��ɋ�ml�2>X_%?H�Ӿr�>;�g_�����-�u�\.$=߻�>�6H?�]��x�O��>�Gt
?4?xG�W���s�ȿ�}v����>��?�?��m�N<��\@�uz�>��?�eY?Fi>�U۾qzZ�]��>[�@?�R?�>8�*�'�F�?�ݶ?���?e:b>L��?uct?tV1?�A>`A$�J���#������=6���%�s>���<��¾�?��PJ��L�$�B�>�U�/�3��<�һa�>�뗻T���	y�<�����ჾ5��;K7�>���>�;=�9�>X7�>��^>���>�0�>̨�:ᚗ�2=����K?H��?2��*0n�T��<ʬ�=�^��$?ZJ4?D[���Ͼeը>��\?N?H[?�f�>���=���翿a|��ҩ�<��K>4�>D�>5,��eFK>��Ծs+D�Fq�>ϗ>�����>ھ�*��"���|B�>�f!?M��>!Ʈ=��?�y"?��z>�O�>��F�̒��jF�b��>�"�>~/?��~?ɛ?X񱾃!8��Ғ��m����X��L>H�u?��?0'�>�F៿�sO��c�� |��g�?�Mn?�gٽCz?�C�?�E??<6C?xG{>���Ծ|ʉ�^V�>�!?���ʎA��%�����=	?�V?�%�>����LYڽ��ؼ��[���w?3_[?��%?���`�\�����<�Ia�}Tź<O�;l�1���>"">���"��=T�>s��=�l�Y9��}L<�@�=�!�>���=c7��A��(=,?�G�Rۃ���=f�r�xD���>�IL>�����^?�k=��{�����x��	U�� �?��?Lk�?$��%�h��$=?�?~	?x"�>K��
~޾N�ྷPw�8~x��w�X�>���>1�l���L���̙���F��d�Ž�����} ?��>��>��>���>X�>9��l��Cb������d��G�����2�������U��v��=k�������͆>�9��I��>�.?0N>۫u>4�>�%���>a*�=@��=���>�ň>%�>��>>B��
�I��%R?����-�ih���о��??�xl?���>O���u��������?#��?�{�?bܑ>.d��Y3��z?h�?��l����>iE���L<�H{==���8��;f����*e>��Խ��5��S�3�T��8?�?1���u�ž�⢽�u����=���?�/?�2!���w�����:�#���cM>�����Ӿp�=��~|�ar��a:k�Gsp�g�=���X?"_?�9e���賩��P�������>`=�>'�>���>yc�=����O�cC���O�(��`�>��?&�>![I?��9?�aN?�VN? M�>7j�>z��a?�ץ<���>F��>��;?��/?7p0?f�?��0?@>oC!����XԾ�?�?��?J��>���>�>����m���A;ֻ�9S�m�h�*���='s�;�,���������=O�=>�d?S���8������j>�7?��>Ӫ�>I���*���k�<a��>��
?$o�>� ���r��o�ı�>�?3%�o�=�F*>;��=��Ā�����=�iż`T�=����D
;��@$<�=5��=���#!X�� ;:Y�;uΰ<�t�>-�?���>�C�>�@��#� �]���e�=�Y>7S>�>�Eپ�}���$��m�g��]y>�w�?�z�?޻f=��=ז�=�|��`U�����O�����<�?;J#?!XT?Y��?u�=?[j#?��>+�jM���^�������?",?���>
����ʾ��p�3�,�?�X?�<a�K��;)��¾S�Խ�>�\/��1~���`D�w�������y�����?H��?�+A���6��s�'����R����C?& �>�Z�>��>^�)�+�g�]&��8;>��>R?$S�>�W?�~?�8b?Cr_>��>�PB���*��X�;��$>�w9?�2o?:��?/�l?���>�9>;T������l��3R�smv��qE=�W>R̚>��>�ҩ>�d�=혽*�6��'���=��>}��>��>���>�N�>G�(��kF?�Q?׾�������Z�ؾViw�z��?�(�?Tp?�~�>nT���V���?�ө?dR�?��U?(�^��I>�e#=���d6Ҿm�>�ف>Tɍ>��>���K�>6��>���>|+�����e���@��>��I?��>�Mѿ��;�I�U�(��'>TΌ����,�>��¾�n=�Q�T������
�i�k�`���k�a�������p�>���=.�	>iԈ> S����n=l�>�
���L.=5A�=�5)���ݽ� >~Bl=��;�����f�=Ӕ�=pʽ��˾��}?<I?G�+?1�C?#�y>�6>��3�<��>����@?�V>��P�����lz;�W������ �ؾ�|׾��c�"͟��C>�wI�|�>�E3>S�=8k�<B%�=�s=�Ҏ=�O�:3=C.�=�X�=�c�=���=��>�Q>�6w?W�������4Q��Z罤�:?�8�>q{�=��ƾq@?��>>�2������xb��-?���?�T�??�??ti��d�>M���㎽�q�=F����=2>t��=u�2�S��>��J>���K��;����4�?��@��??�ዿТϿ:a/>�7>_>x�R�M�1���\�I�b�YtZ���!?�C;�E̾D4�>��=))߾V�ƾɰ.=��6>�b=�h��R\����=�{�@�;=�l=�҉>�C>�l�={D��m�=|�I=��=C�O>���m�7�^5,�$�3=x��=ҩb>d&>s� ?�� ?�?ɧR?�}�>�j��=썾�z����?�5>��?�M>�2C>3r?J�??�XY?��?�I�>]!D����>IA�>w)�V+2������>�<�?���?�X�>�E��'��O��!�7g�<,��>�� ?ŧ5?\�>>�S|࿨�K��,���G����<����z(��L�c-8�0 ��a�>�v�>���>E�>G�!>&>,=:>���>�>��l<L�8�V+��_s��,)�!�Y��n׼:E=&�%>3bM>\��>�D�=���=&��;D-��d���:	M�=���>��>�}�>}e�=We���1>������J��ø=�%���@��'b��{���/�ӌ>��;>��Z>"Y_�ڑ��Y?)jS>�B>2s�?]�v?CG>����־ҹ���Hb�V�d�lm�=g>?�<���6�?�^�óM�/Ծ���>o%�>({�>�+<>��:��a-�">=���������>ƾ�9�=��?���Z�k�������c��k�=a+[?.�����4>�gS?��N?�-�?���>�D�q^�I�<�������=.KW��Rн��)>��>|kI?b��><���M���ƾμ���i�>��N��M�������?�O-�<��߾�h�>���7�Ծ����_��D<���bH��,{��4�>1GA?l��?DX��䄿gX`�����&�;,p?I�q?���>N�?��?RK�����g�)�>�a?vu�?���?4V>^��=r���>�5?Ί�?�ܓ?N�n?T8���>�[V��>�<�uԭ=�/(>K�=3y�=�'
?,�?�r	?�pK�W����u��W�0{=��=�9�>�>볐>��=���=6�3=�O3>m��>�k�>��>xi�>��>����?����X?�B�=���>QfK?\��>6_(=gԼ���'oI<��t��$��P(�I���:=�y����y=ջ<P�>�ſ�?C�U>p��#��>n�Э��wt>hJ�>]n�=~W�>G>���=�̵>4�>���>�>i>:>q=^JӾ��>@���H!��$C�śR� Ҿ�8z>�����[%�8��&.��>pH�ߠ���}��j�?'���@=�ĥ�<�;�?na����k���)�`�� y?�G�>�$6?���∽�>���>���>�q������>ȍ��:���?���?�?c>�E�>��W?��?D51�F?3�K{Z��u��A��e��`��Ӎ�Ӗ��.�
������_?��x?�NA?�9�<�z>Ԡ�?��%��֏�0�>c /�;�V_<=�4�>� ��e5a���Ӿ=�þvT���F>�o?��?�2?X�V�B�r9>��8?^�0?'�t?3�3?'6?̷�5'?5'8>Լ?�n	?g�7?�/?�?��K>A�>��˼�`.<~O���"��Ӕɽ�E����!�AC=[G�=7/���7�<�Pf=�� =HR����ѻ��O<O�&V�<o)�=��=h��=��>'^?���>��>��7?	z���8�S���to/?��&=>����u��\�����򾤟>٠k?�m�?:�W?�\]>��@�2�A�E�>�щ>u�">�W>��>��뽿$E�y��=>�T>�'�=3�'��L~��	����$
�<kf>���>�{>؆����'>;W����y���d>�R������S���G���1���v�#6�>�K?��?���=D������+f�&)?!f<?�tM?��?,Q�==�۾#�9���J�-R�$�>��<���<���h ����:����:�&s>4/���Lƾq6>��߾����f�XkR����伇��]5��P�=0ξ������ؽ�_�=��=�^��J��������CH?��>�|�F�I��7þ���=&JZ>	�>�0����=>9@����-k뼣��>(��=	@@�8"�3U]���g��>�E?z�_?��?�\u���n��WA�M����*��v.ؼ�?ъ�>R�?<>ͥ�=<��}I�@c���F�h_�>��>E��� E��ä������#�k��>N�?�##>�k?f/Q?d4?)�`?]`,?W�?���>���J3���&?w�?w�=f�ٽ��Y�_:�«D��d?k�.?�8(��z�>>�?9?�h?�T?�-?�"5>�����D�c7�>��>��X����&G>��@?��>�;]?	ԃ?�z:>!3�R����g��잋=+N>1 :?��?��?�U�>vz?�R<����=;?��n?�Nr?�42?D}��d�>2��=��>��d>���>�+?f�3?�&K?�*{?��?�݁>?��<
��i���)�������X���Q=tC >_�<�]����W�t=JĖ=U�;�WW<��w���˽0��=:�=��>�݄>�,���
G>E���`�u��/s>����Ρ��F��y{��D=K;�>���>ge>C$��?�=ݫ�>���>�/�0�?��?#<?�/�<��`��	��!^��q�>
�P?���=Fn������f���">��|?�\`?wO��M�b?��]?>h��=��þr�b����c�O?7�
?E�G���>��~?d�q?P��>�e�-:n�)���Cb���j�Ѷ=`r�>LX�O�d��?�>m�7?�N�>@�b>%�=ou۾�w��q��i?��?�?���?	+*>��n�X4࿷:ؾ�����[?-��>򁐾Ŗ+?,����Ҿ�.}�ҳ�(U�$����뾥 ���!���.��l�{"R�o�=@�?:�?�]?�ZL?�����R��o<���o���f�� �8���3-�R��mc�:ǃ�PB�IH+�����摽���O A�D%�?��?�m)��>�>s��������>�e���C��O�=�/���>=�=��.�Dua�5\پ�?�5�>���>T3?� T�%�.��*��O=�����[L>2i�>�~>f��>2j�9�n��*�����sǾ�[����r>4Dd?iL?��o?�ū�Iv,��|��,����.�䍯��SK>ć>�z�>�l[�O� ��> �Yu:��p��/��ꏾ�
�]h=a,?��z>��>H��?Dh?��3��q�{�l�-��=�1�>��[?���>�>�	�7��i�>݂l?rK�>�>!����� ���{�� ̽i�>�#�>�K�>�jn>2/���\�@y���a���A9�3��=��g?1Y��?e]���>�R?��;}m<�١>�z�W"�ݫ�p�&��>�?7\�=U{:>�ž���F{�wq�� �,?���>�8��J����>��?)��>�ϑ>~�m?جY>���#�Z>u/?��q?�a?�F?z��>B���󼵽�ꏽ#�H�c��<�Ơ>$�9>iT5�"�`=K�^����HA�Y�=?=�4I�E�����:��<#�=��<=~>��ٿ2�N��ξIL
�9_��!��s~���ν�X����Q�g���=��w�#��`��1���M�	1��(���^���\�?)��?�}3�A�<�H����u�N�
��l�>
á�� �
[���h�1�{�1��]e��.�!���V�pЁ��r���V7?E�޾=��ꙿ�O��I?Ba+??��?jr޾���h����(k>'��=F%0��:ʾ�s����˿֒0�u��?���>�����	�e?=?ꇴ>^�>σƾ�M���j>�?_�>�l�>&)�|Aſ����C1>���?���?&�A?��(��e�:�p={��>	?�y<>��1�����,�����>Yg�?ڊ?�7b=m�T���7�e?-ȃ;-eF���޻[��=���=�=s[���G>�>���HA�̞׽�6>'�>�C�m���@c�FT�<�Z>�Jѽ�ݛ�5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=v6�����{���&V�}��=[��>c�>,������O��I��U��=�����Ŀ��$�%g%�� I�'����<@<����/)�"�߽��y���o+��$�=��=[�X>���>��V>��->��P?�b?��>ЋZ>����|�Mj��dཛྷPƾ&HH� �Js������v��������v���W7�� ��!=�Y�=r5R������� �2�b��F���.?)l$>0�ʾ`�M��V-<klʾe���E܄��᥽!,̾Ƙ1�D#n�͟?;�A?k�����V�"���\�����W?�T�͹��謾��=����C�=o"�>:��=����"3�@�S���1?��?χ���۔�w��=23?�B�<��5?й?�g=.M�>�t?��l��ö�>�c>]��>���>�2�>w>�ѧ��R��/?O`?d����UK���>(n�+3����=�>�,���<R��>:�):at���Q`�\w.���[=�8V?b��>��!��������Us����x</�?�*?���>]�f?@�:?�]=����?�F�)��r¼=;�K?y�`?���=j�ؽ�eپ�
��$C0?��`?�S{>-���d���(�U����?��v?��&?-R��]~� 𒿡1�hl<?��v?s^�ws�����L�V�g=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�%Þ?��@���?��;<��V��=�;?k\�>�O��>ƾ�z������)�q=�"�>���~ev����R,�e�8?ݠ�?���>���������=u䁾�!�?o�~?:ߚ��g}=�K���b�����dȽ�@$=TT��~��`	�8w@��M;����|���	��r>v�@����`��>����>ܿ.�����~���p���?�{�>��u�vk��qt��X���F�Ǫ���>C?>>l�ؽ����(��#uL�+�ι �?���T��>k�&�`����ξ�H�:C7>-И>(V�=��Qٙ�ˠ?\�A�����.�2\z?��?�^�?�D?ǃ��n�k�����C>�>;?諅?"�U?���<��*�[/V=��n?u�ؾxv}��dL�a�r���?�>?��\> !����c=;(�>��>��>b�%�y\̿�˿{���H�?�Y�?���?O�?/x?X�(�(�����|���f�m[>ԛ?�5�(7�������M��x�����>?`?�����T�_?��a���p���-���ƽ�ڡ>��0��c\�H=��c��4Xe�����?y�m��?^�?x�?���� #�:6%?��>ٞ��%9Ǿ��<���>�(�>+N>�M_�\�u>����:��h	>���?�~�?�i?���������U>'�}?� �>\�?:�=�t�>�i�=��8<�K@#>�Q�=�s@���?k�M?m�>-I�=��8�z
/�[ZF��-R��"�e�C�w�>�a?͆L?�b>3ĸ��1�C� �̔̽�d1�"~�c@���,�X߽D-5>��=>�'>7�D�)�Ҿ��?]y�t�ؿqf���'�N4?�܃>e
?����t�5�
��%_?�x�>@"��+��71���x�џ�?K�?��?��׾ZfǼZ�>���>�P�>�Խ�Ҡ�qX����7>��B?�5��3��m�o�ٽ�>���?��@��?��h��	?���P��Ta~����7�b��=��7?�0��z>���>��=�nv�ݻ��W�s����>�B�?�{�?��>!�l?��o�N�B���1=7M�>͜k?�s?�Qo���n�B>��?!������L��f?�
@u@`�^?)��ۿꏪ���Ͼ]���Sa<�(X=�r^>;'� ?=�6� <�B���x�9�e>���>��2>�%�>�%>��>��/>���30!��ޣ��s���XB����yվ'�W�ܾ1/��j;�;վwˉ�~��<9@��悄=Kc�(A���<���=GdS?�Q?Fs?'�?ڎ%�I�
>�C����=)O*�0��=>|�>\j,?E�D?x`#?���=tՋ�~�c��E~�����ˆ����>"5Q>x��>�N�>9��>m��;��D>��J>Qy>��>@�=�/<	�?=ՋZ>O �>Wk�>sݪ>D<>H�>Vϴ�2��Ӝh�r
w��̽\�?���T�J��1��(9��t����h�=<b.?J{>����>п1����2H?�����)���+��>��0?�cW?��>�����T��:>]���j�`>�* �Jl���)��%Q>�l?`�f>�u>��3�d8�H�P�7}��^|>t26?<趾pF9�{�u�<�H�XcݾAM>�¾>D� l�����Z�lti��{=�w:?̃?!3���㰾#�u�B��xRR>`;\>}f=�y�=^YM>�Rc�O�ƽ�
H��k.=)��=o�^>��?I">�@�=�=�>��P�@�'��>YN4>v1>.�<?��#??
�O�˽ry���w0>��>(��>,��=S�A�I��=���>�fH>8�'��S�����=���S>����ej��x�P_Z=���� ��=��@=��!F'�3�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>9�~���� ��w匿�U=7^�>s�m?�ƾr;���N8��?�f�>@�ݾ�ݔ�8���H��,�>�.�?%��?&G���A��mA�8��>���?��^?:ə>�����s��yޖ>�WI?"1h?ֱ�>R�����2�?� �?uk�?q1Q>^�?`c?K��>x�)>O��_��8q�	a�`9���5?����n��@��+\r�܈Y���r���p���=��>&Ƚ�_�+�2>�P�����՝ݼ�X�>�Kv>0AQ>�)�>�h�>���>^)�>_;>��/]��t���K?~��?���2n��O�<ş�=�^��&?�I4?�k[��Ͼ�ը>��\?d?�[?ad�>��>>��&迿~����<Y�K>^4�>�H�>$��GK>��ԾH5D�Cp�>З>+����?ھ�,��[���A�>|e!?���>lҮ=8�?��#? �k>8d�>��E����?;F���>��>E8?&�~?�?>���3� )���⡿5M\�n�J>Q^x??�?
�>�؏�����\)����@��؇���?O�h?��꽚?ׇ�?�}??�vA?��g>�<��P־���s�>I�!?@��K|A��%�����]?q?JS�>񙓽��ֽ�P˼�X�{���?�D\?MX&?n'�[a��þ���<�h��`S���;�E��Z>�.>`��~��=5�>H�=��n��7�K>P<���=�!�>p�=J16�<g����+?���䴁� W�=O�q���B��Zz>��J>�]��I�]?d<��3{�K�������^�R�:{�?oo�?�O�?�f��ץg�C=?|��?��?��>�Ь�97ܾᾩ�z���~��F�u�>��>!t����VX��KŪ�����~н	��5X
?��>[?��?:.O>LD�>i���r,����[��?Y�����@�6=��A��������<�cž�w�7�}>f$�� �>���>R��=��>M�>L&=��v>��>=��w>Ӧ�>�=�>�h�>��G>���O2��s�Q?ԃ���'����U���B?e?���>�zr�~����2��|?�V�?��?�r>V�h�P+��w?|��>b��j
?v|6=ܕ��*�<�߶����B��v��č>��ս;��sL�^�e��3
?V�?h�����̾s�׽n#Ӿ)�>T�y?���>:p(�W~�}���r�֍�^��>�~�HF��X.�ډT�Fi���y�4:�������S�}�)?s&�?O�Ѿ�3&�;�����T�I�(���l>���>�G?O��>6^3>��G���i�^���D��[Ҿl�?�h�?�P�>l9?�)?��I?#�A?�"�>
�>O�^��6?����|>�n�>��5?R?��3?ي.?0�6?�/:>K ڽJ��K]���$?5P'?� R?�uM?0��>����ns�7��o?��&=����`n1>>��ѽ��=�h=*��=�?A��)�7�@�����k>�"7?���>?�>ꦎ��S�����<Q
�>Fi
?S<�>1�����q� v�s��>	2�?U���e=Bb(>b��=]��kT�~��=�V���F�= 7����?��e)<A�=M�=��}�(�s�/�����;"��<%t�>�?�>�?�>�>��j� �H��uu�=�Y>�S>�>}Cپ�~��k#����g��by>�w�?Ry�?��f=7�=%��=�|��YV��1�������$�<?�D#?%QT?���?Z�=?4l#?z�>�.�}L���_��P��[�?]!,?1��>�����ʾ�񨿔�3��?V[?�<a�����;)��¾��Խ�>\/�i/~�����D�(҅���������?῝?�A�N�6�,y�Ŀ���[����C?�!�>mX�>o�>T�)�2�g�%��1;>Ê�>:R?j�>�qF?�t?�l^?Шl>�+0�R�yϕ�ܬ(���>!A?Gb�?��?��x?��>��1>���;�l!�����������=�O>��>�Z�>ҟ>��=a����d����Y�dJ=`S?>���>�G�>���>��o>�*�;b�B?�?œ_��4�CG��gg�� <3�~��?��?��(?%�(>�o���L��~���>���?���?>L?.�v��W�=c,�6�߾����B|>��>�}>v\=hs=z��=�ڄ>)`�>v��=�M�7A��Iغ��>�n?3�u>Cƿ>r���r�o|���M<A��>d� -��M�Y���=ۘ��X��Щ�<�Y����������r��oݛ�n{���>\��=�,�=���=I{�<��ȼ���<`R=�O�<��=��y���e<��6������G��=pC�1Ub<��L=g��1Ӄ�Y�?�O?6�=?�cb?��*>9�����Ad�>8Q�K�?"�q>�g޽�ԾɝK��Z�5�����i���I����`1 >�n�=PE>,ŏ>�*�>7�<в<>�/�=`�$>���<\Vl=�<>���=#$>p��>b	�<�=�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>|8>[�>˥R�aL1�Y\�Mob��Z��r!?n.;�g7̾Q�>�s�=y߾�_ƾ�0=:�6>&d=�p�H\�8͙=�jy���;=d�j=,��>*�C>bJ�=�+��bI�=`�J=�"�=<O>1���eF8�e�-�62=y��='c>��%>���>�?�>?�Q~?$��>NW��¾I�m��M�>�f�=2?�,<>併��M�>�uG?�I?�A_?C%^>B�,�'��>Yh�>���m��������
�J�MI�?i�j?�>�L>F��Q�+��H9��ƭ<� +?��&?��?�~>(E����'�I��TX�B���j��)�y>��j�d���C�l>e�����	`�>�]�>%)�>lx�>��T>��Z>��>y��>ѧn>�	P=?ͺ=����` �ă�:]>\�d���˽�T=�$���7��}c�W������=/ŋ=󘵽���=ha�>�M>�I�>��=̏���,>����L�zѰ=�Z����@���d�<~�L/�͟8�U|@>��Y>F���ቑ��8?�X>�?>v��?�ls?
�!>
S��پ�H����d��(T�7~�=^��=�-D��@;���a��N��}Ծ�<�>u�>�t>D�	>'-���W��>���R0��Uj>�����>��S�b�g"���ڧ�=�[��Z> d?r�����>�H?�+9?�ǣ?��>鹼=����\�.�T�Ͼ�D��$>��6��iS=<C?~wG?t��>˸��2��n̾u+�S]�>1���R�Q�����98��h\�ܻ̾J?�����!�t G���Ò���H�E1��tg�>3lE?�a�?�
d�W���b�^�֢%���ټ�?��{?y��>R�>B�?�=�sо��Y��-�=G�f?���?�}�?�6O>|��=eț���>��?�?�*�?��h?#A���>�C%<�+'>U��\�=?'> ��=��>�?ޑ ?�^ ?�w\��c澏���t�~b�<�F�=n,�>13�>��e>�;�=�
�=[o�=@Cn>H��>���>�ga>t�>�*�>����s���?	g>k�>+?���=21�<�e�<��>�_<����p��~%����Լ��6=Z{�=��>c�G>�g�>�	ʿ+M�?.>�>����
?�X9�������>��>
�=���>~�+�Ku�>�?qI�>�Ϭ>���>]xT<�[Ӿ&>|���!��)C�C�R��=Ҿ��x>�q���"�:z�֐��B�J��n��̝�j��Q���~=�{Z�<�B�?���ؾk��4*������n?]��>�:6?:̋��ׇ�>>�=�>Q?�>Q���zr������!��%�?���?��b>���>�W?��?�00���2��iZ��Zu�$�@���d�U�`�ԍ�פ���x
�����Sn_?�x?�]A?���<,8z>#4�?�X%��܏����>ζ.��l;�ζ<=�c�>꧰�mb_�` ӾgľK.�D=G>yVo?�?w?�W�(T�=��2>��$?܊3?�r?X�3?�?!�*�5�?�v>�/�>��!?�E*?��A?DH?Tx>i1>P0�f�����L��|���"�!�������&2�<No=��~<�8����Q=L��<k�=!Ķ=���=-=8�<�ܻr�U=�
>�l�>1zW?ѽ�>=̈́>:"5?#<���8�2<���0?��T=��|�U�������ni�3_>��h?8+�?%�W?dMa>�!;��Y?�֐>�*�>�m>��e>�F�>S&��)M��dQ=���=�}>j�=��5����!��C�����<��>7��>��s>(����0>����u��d\>I�S��¹���V��$D���.��w�9}�>�7L?[?C9�=�����<Od���(?��:?l:K?�(}?��=�vپ�9�z�I�0���>�1<�}
����Ѝ���	:����"t>�ɡ�Zܠ��Sb>����r޾z�n��J����M=���nV=�� ־�2�^��="'
>-��� � �8���Ӫ�1J?��j=}x��@UU�yt����>A��>��>0;�:w�)�@�$����?�=5��>);>�<������~G��4�3�>�C?E�^?���?����9�t��V@��|��D��<����I?�ۦ>�F?��S>�=�N���\��c���A��r�>�&�>�Z���C�gş������$���>$�?�w>J?�WO?�	?�zb?��(?�^?y��>4e˽Ax����?�y?+hݼQ%���=f(g�Bfb���?�?ӓ��6@>Ia�>���>�?9�?��S?5b>M�N�����[>浕>��B��㠿0��>hh?�#սa`?�p�?^��=_����Ua�э˾���>�8?f#?�0�>��a>���>í�� 7�=��>fc?�+�?��o?2$�=��?�M2>v��>0��=	��>���>	?�OO?�s?.�J?'��>6��<�?����#s��O�yc�;��G<=jy=���
�s��0�
��<�p�;醷��L��/�D�������;�g�>��>l[���8�����vg���z�>t�O���ᾥჾ,C��	�����>�X7?L!�>e������>�D�>�pB�[�7?V�?JG�>��>�Xu��ݾ�䟾�>ӡ?ǋ�>�P���ʦ�.�h�͋�=��w?��p?��;�E#��nc?�nZ?$���=��k��OiL���C�O?��
?t�<�P�>"~?�q?f��>�lo���n� ��)ba���i���=��>�7��`����>ى1?�y�>��]>a8�=�Ͼq0t�#ǧ��1?a�?ee�?��?��4>��n�Gl�t�.�Ρ����e?F��>�����X�>阽����6���Gm�A �����󯾲e��q��G���h��U.�ƌ�=��0?>�{?�J}?��Z?�� ��m�|Rw���N3P�VuҾ��$�D���?�,;�� G����2�U�݄���<�s.�T�%��v�?/p�>`m�;�;\>6fr���߈��>@�Ӿ�����g=)��=_D�=���=����2���]���%?x��>*�>QuQ?��z�_�X�ſ�����$V�2���~�>yԦ>	�?-�>=�@=�7g��+a�p�����=t-v>
yc?�K?�n?`z�E%1�-���L�!��/��i����B> {>���>F�W�����9&�X>�?�r�G��+w����	���~=Ϯ2?)&�>|��>-N�?�?vy	�{i��gx�4�1�k#�<�)�>�i?�?�>i�>��Ͻ�� ���>��l?���>4�>����Y!�K�{��ʽ�"�>�ۭ>&��>�o>��,�R"\� j��܂���9�Ex�=Ʀh?B�����`�[�>�R?8*�:�G<<z�>J�v���!�����'�R�>�y?j��=�;>�ž/$�ʣ{��1���&?-�	?����E-���>��?���>h�>!'�?���>�ž�N��%?��[?��F?�&<?x��>m�:=,Z���S̽�W)���X=)܈>5�b>��T=��=� �hg]�-����S=M�=�����Ľ�[J:���v<Ӹ#=��9>��ۿ�K���׾���9����	�C3��պ���?���o����t����y�#%�{x,�ѷV�Vc����/k�5&�?ߦ�?fm�������M���Z�������L�>l�s�7�v�8��ؗ�������߾�{��� !��HO�o�h�:.e�V�'?�����ǿﰡ��:ܾ>! ?�A ?9�y?��<�"���8�{� >�D�<�-����뾬����ο�����^?���>���/�����>ߥ�>>�X>�Hq>����螾<1�<��?0�-?��>t�r�%�ɿf�����<���?-�@�~A?*�(������U=C��>ґ	?��?>�81�!F��谾Z�>�7�?���?;�M=7�W�$+
��je?�L<C�F�$�໹;�=�<�==����QJ>g]�>�o�3]A��ܽ"�4>���>B�"�8��7U^�Mֿ<;�]>z�ս礕�2Մ?A{\��f�r�/��T��U>��T?�*�>�9�=��,?Y7H�]}Ͽ��\�+a?�0�?��?�(?fۿ��ؚ>v�ܾ��M?^D6?���>�d&���t����=�5�(���j���&V�m��=ʬ�>Յ>��,���]�O�2I�����=W��{ſ�"��a��|A<Iw������3н�CK�w��E��^����`�<�E=��">p%j> �'>�xt>�S?O�U?�;>��)=I���cZ��,�����=�X����J:���(��ϓ��v���Ϸ�����t,���D�.��w=��)�=	2R�ʔ��ź �U�b�2�F�+�.?�W$>>�ʾR�M��+,<�oʾ~���*����a!̾A�1�`n�ȟ?��A?������V�X����ӹ���W?�� ���ꬾ���=����=�9�>	٢=���=$3��|S��-?��?���A^���>d� �ߟ��^22?|��>��<r\�>��?>e���ὴ�V>
_>�ϳ>ɤ�>��=� ��`m���>?,Fa?�EP�����"��>O���䁾�kM=k�=� /�i�3�(�J>�;A������g��x����[V=�Xo?���=��"��7/�p���~�9>�>Zy�?��?�:���?-�?�:�>�)��@���.$�����8�?��?H�O>قžQ��J쏾C�P?�'�?�<��nU��4��N'����o�"?�hm?,](?
D�=)ԃ��=���ƾOUP?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?p�;<��P��=�;?m\�>��O��>ƾ�z������3�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�ٕ��Z�?{�?m����>g<G���l��n����<`Ϋ=���E"������7���ƾ��
����{޿�ӥ�><Z@3V轂*�>	D8�Y6�TϿ��\о�Sq���?6��>Q�Ƚ[���/�j��Pu�P�G�4�H�����<�>���v�=�:�J����*�Tss=5'�>��۾U'?u����)�q�&>y�)?>�)?z�/>GM��ڍ�?7��L�h�}������?"��?���>�p�>*��<pBۼ��s<M�;�\I?p!u?�S?��3��t����,>�k?o�����`��{4�`�C� \>��2?RP�>6�+���{=�>�q�>�D>�.�LĿM|� �SS�?1(�?�k�]^�>C��?Gs*? 2�;ۙ�7j��n~*��Me�HLB?g=1>��þI�!��s<��ɐ���?��/?|w�qG�%_?���m��e��Ξ��6�>y�O�����`뽔�">��\�md���I��ۃ�?�~�?vɥ?�#����B�B�?�`�>#�$���W���̽��7>C �>��>g�4��P�>��Ѿ,�l�A��;��?���?e�?����*��߱�=bt?���>��M?s���lq]?�β=��N=;��>7B�<,��>|lK<�1&?��,?]�>s�M��Y���x-��(Y���A�r��uw���?�`9?rLQ?�Q�<��$�����F'��=�<�ǾҸi���Eʰ��NI�Q>�>�/�>E��1�����?Hp�5�ؿ�i���o'��54?9��>�?��R�t�����;_?mz�>�6��+���%��&C�P��?�G�?#�?j�׾�R̼�>F�>�I�>��Խ����q���:�7>&�B?���D��g�o���>���?�@�ծ?�i��|?å��������d��#���>�l/?Z:�����>?��>s��=Cw�W����{n�Z��>
հ?�0�?�j�>�2r?�x�L�M��J�=�N�>JOo?>?�N�k��
7>'�?em��v������|Mg?��@�A@v�X?�a���hֿ����,N��/���-��=#��=h�2>��ٽ�_�=�7=��8��;�����=�>5�d>�q>X(O>(b;>L�)>���8�!��q��Q���:�C�������Z�X���Wv�_z��3�������>���3ý�y���Q��2&��>`��>�=��U?!Q?<	m?FH�>�,O�V&>�a�� �=>�4��=��>��3?�1H?��'?�n=�O��m�`�,)��B������Dq�>�R>$��>���>��>��;��G>�>>x�x>2�=D&�<�S�	!�<e�U>0�>e%�>�H�>�C<>��>Eϴ��1��e�h��
w��̽1�?{���T�J��1���9��զ���h�=Kb.? |>���?пd����2H?%���y)���+���>}�0?�cW?!�>��L�T�1:>9����j�*`>�+ �|l���)��%Q>ul?\�f>��t>�\3���8�qUP��m���|>O�5?z��k`9��u�3�H��Gݾ{kM>Ѿ>23H��K�Hږ�
�~��i���z=��:?^g?�ɰ�����u�'����^S>��]>b�=�"�=�wL>&.g�)�ȽZ�H�T,=��=�^>f-?Z�@>�R�=��>9�����S�u��>R�a>�
>9�9?3;?с|�|�齟&����)��z�>�>�>G7�>$_�=*#b�B��=���>�_s>sA� ���n��1��N>Ef����n� ���q=/=��<�=���<���JH�EB�=��w?v��œ��������S?8�?LXQ����PV���I�������c�?#@oЖ?�����U����>� �?q*��̙>��?�o.>�P���9����>��x<�f��m�;�������?�V�?�|�젒�1�k��X�;�c?�0U��o�>�y�3Y��B����u��$=���>*;H?�O��3P�h�=�5�
?r?=b򾵪����ȿ>|v����>��?���?C�m�e@���@����>£�?�`Y?P^i>�_۾1fZ��}�>ѹ@?fR?�&�>�3��'��?ݶ?t��?�I>c��?.�s?Wx�>�x�>L/��,�������=�~P;Q�>*>����h\F�ӓ��_��1�j�\��_�a>^�$=��>��GH���F�=�L���7���g�|��>�q>m�I>N�>�� ?L�>�m�>�=�k������z�����K?娏?���f*n�H��<��=��^�_1?cG4?��Y���Ͼ�Ҩ>�\?b��?x�Z?X\�>����=���ڿ� ���7��<�K>�K�>�N�>�Љ��ZK>��Ծ�D�\��>	��>e��LNھ�=�����W�>�o!?���>M֭=�� ?*&#?8fm>~ó>h�G���Z`B��w�>d��>`L?.l?�h?;�����3�}�������u�W��1[>��w?"�?Z��>3I����P:��LGD�[#d���?�gg?��ӽK?4��?{�A?�/>?��\>����ԾỊ��b�>g�!?�K�
�A��R&�/��)?
�?Y#�>�H��?Zؽ�ؼV�������?�x\?A�&?T��wa���¾�<�$��#W�Aw�;�J6��->��>����>]�='0>�)�=p)m��P6�FR<�ɼ=�d�>��=��6���-)?s��<�-��E�>��q���@��_>��o>�d¾.YX?��G�ơy�/���yИ�N:O� O�?���?��?��㽪�i�ʀ;?���?Zg?u��>�G���Iʾg�ԾD�n�Z#�������=r��>�
�vA뾢g���§�(.���y������Լ�>=��>�`�>�i�>�>�-g>lX����������b!h��@"��T�X�����Ӝv��	Ľ�h�鮻����H��>�����>`��>K�&>�0>&�>�ʃ=���>@5,>hQ�=�fi>��?��t�=)P�=	#�=,�<U`?�d龺G�VN��,K���{g?��I?���>�\�=��H�������=?���?1��?u�~=���a�g����>MA3?{���8?l+�=!�?�Z��=J}����h�M]�N>G�D��>L�h��Ox��l=��{]���?��3?A|@=���� ���7�t=Cp�?��(?��)�1�Q�ӵo���V���R��Y���h�N"��Yb%��Ap�\�]������J�'�3z*=�}*?
��?�(��7ﾄӬ��5k��e>��e>-��>[�>s��>��I>��	�1�1�YU^�߸&��a�����>	P{?���>��H?��;?�
O?�L?6��>Ҧ�>b&��R��>��; ��>�`�>v�8?-?��/?��?�*?6c>(w��J����bؾ�k?�*?��?x�?�?b���P��<Jj��f�By�����x=��<��ٽUpz��\=��U>�,?��k�9�����n>�0;?K��>y��>�Ʉ�oV���9.=q�>Y�?t��>���[v��I��"�>K��?v �ߥ�<7�>�~�=W�d�Y����=�μ�Y�=>�8�9.u�')�3��=Ս�=2T�;����u,����T��f�<lG?�Z?�е>� �>��ݾ�L	�پ��w>~p5>�>�n>M������͏���}�|�V>\^�?>ó?Qe�=��>h"z�i��%ݾh"�@(�����>�x�>�#?��P?�Ұ?_�f?
�7?)�H:֭#������YW�3�x?`!,?���>v���ʾT�w�3�Ν?[?<a�Z��m;)��¾r�Խޱ>�[/�>/~����D�� ������~����?ڿ�?�A�I�6�ix辪���7[����C?�!�>�X�>��>U�)�K�g�2%��1;>��>�R?�Y�>r�N?��z?�|[?��R>ë9�zQ���i���縼��!>��>?A΀?���?�Bz?F�>��>��&��߾I���/��o��#���uf=��W>�>+��>�j�>�8�=�νW���G�@��!�=�kh>Һ�>�E�>�x�>t�q>���<��4?�?$:þ/>$�jI>���;��6�?C�?CF�>d�ۼ*��X�?�����/?͸?��?�Ew>ļ#�< �<�w�|n�C��_�K>���>�8�>�b=�Z�*��>I��>��b>W�8�d�侰e^�7���>?�Uj?�z�/�ҿ��w�
�R��ɾc��=������d������F ���>���$���\����j���bT��M���[�;+�
�Y��>+�|=hv>�l#>a��<7ཀޙ;�����5���>���9��<b!��Z��/ƽq�~<+?O=��F<�FW�A]����?�n?]!?�{�>�1?��|>��<�o!?����I@?�r�>:�>��ľY��8���S�c�V�]��	��\����=>�F?�9.U=q��<y��=j�=ค<�m�=���<�0������.�=D�=[��=1O�=O�.>�J>��a?�g���(��W%�so���*B?�"?d�����d?��>��[�~h����޾�	v?*��?�N�?�}�> @�d��>�>�U��� �>�C>��<h+=�oH����>��=b�ѾE珿����mY�?�y�?{�?����?iĿ�z�=��7>8�>�R�S�1�R Z��&c�tq\��!?l�:���̾ⵅ>7�=�>߾0�ƾ�17=�7>��d=��y�[�Q�=�{�,G==D�i=2$�>U�C>C�=�Q��?��=�Q=��=�/O>����<��y/�2= ��= dc>m�%>��>ժ�>T?��V?�[�>F���������`5�{t<$�}>��轂/>t`.?g�7?�pG?Մ??R1>>��>{��>F�9�PS�R����˾)Zս���?��?`�<�%�=�:��O$���-�)O�<�7?L�?P�h>�A>K��L�ۿ�{�u-�1!T���P��i-�i[�b�<dSX����㒚���D=��r>�!�>�u�>/i�>DE�>�s>��>uQ{=Y��<.^�:�`����=<Q=���=��ؽh�<�6�������;�K�;#ǚ�cgʼ�j�������<;'�=SO�>_K >���>��<������>��M��*G��Ρ=�䱾}$B���g�<�v���&�0���%]>I�P>�GȽ
򐿯� ?|��>�,>E��?uEi?p�>�F��:mȾ�y��F{��Y��#�=^��=�q��VE�^�(H�
������>�>��>`Vl>��+�r�>���y=M��u@5�T-�>X*����һ��q��7��B�(i��G���zD?%D��4�=V~?��I?�ُ?��>"��Hyؾ��/>����K�=����q�9���~?�%'?���>����D�e/#��%���R?�:,���h�H���ڨ`�N��<I����?RZ��v��v�g�~y��
(u��-߾�il>%�&?X	?f��?��ý�^6��;��@�s�.�C�>�E?�U>}M*?uo ?m��d�þԯ���y�3�u?���?o�?y�<˷=.޼��/�>0� ?��?��?�n?��Z�6��>�I�<S>�yǽG��=��>5��=�
�=��?χ
?XY	?N���M�8g羈����Q�f\�<
 �=~�>� ~>з�>i��=D�s=ݍ=��S>8?�>��>#�g>䳥>���>�]����	��(?X��=�B�>��+?�x>bM�<%�����=�2����Z�"�5��g��(����o<�$λ=?������>�pÿ�-�?��U>S� �	�?.?�UgY��@>�n>�xν��>��5>Zqq>�Ş>�?�>˔>|��>A�2>�CӾŀ>g��Zd!�8)C���R���Ѿ�wz>ʙ��V&�b��+����II�=l���f��	j��,��B9=����<�F�?����m�k�n�)�G�����?�Z�>�6?wԌ�3�a�>���>�>L��Ɛ��Ǎ�Bg�[�?���?��Y>�&�>`A\?
/?xȼ���I�U�T�	�t��X9���K�^�\���3��/3��M��S?�l?�T??'$ =���>1o?��������D>չ3��(���=��%>P��Mai�l���dܩ���ƽ� E>�o?̀?b�?e��mv��p_>�c9?�c%?g^b?jL1?"0?��N*?��
>��?�?.l6?�� ?^�?��=�n�=�˰<�}��ㅽ|l���U���L��d8y�I�<`��=�\����}�0=�^=i�;2*��2�<zb'�x��<[B\=�+:=F��<1 �>�VU?z�>�.>>nw??��H�Z�n�9ZV��k?�׻�Y���?��`V���뾰o�>��~?���?V&?=
�a�
%F�:�;>Ν�>!�нkBm>E��>�_ͽ�����n@>��=��=�R6���<4�����t[_��o>k�=@��>�O6>Qp'��}���7�{��~�;>�}ܾਮ������A���L�^�7�oJ�>k(I??Ǎ�=��˾@/̽m�_�v�?u�I?�?�Џ?��>�NؾU������7�z��Ņ>�Ĉ�9�.��j��+)��Kc>�_zO��ch>��L���_�[>������n��0H�W��(|=���SYM=
{�&վV�}�Y��=��
>�$������������I?Z8z=���IZ�'����>���>��>�EP�i?}�pB��7��?��=���>�>>㳈��_쾃�G��r���>��C?�s\?��?����Sv�)=C�� ����*�?�s�>�??^X>��=�l���5
��Ya��H���>?��>2��D�䒾�4���B"�/r�>�� ?a�>�8?��Q?�{
?aa?{�)?�?OǏ>���t8��� "?�v?�Ge=4�	�Q��f�e�^�^����>��>/��C��>��>��>� ?'n?��A?<cm>���:�4����>\Z�>b�:�d񭿦'�>�F?��c>�e?G<�?ހG>b���?������Y�C>ދ#?Y�?w~�>\��>���>Н��o'�=ؖ�>�
c?�/�?��o?{q�=��?�2>��>o�=a��>�|�>T?PO?��s?��J?���>��<+���=��.�s�>�Q�(�;J<��y=͹���s����&�<�9�;�r���"��W-򼈫D��2��C>�;�~�>��b=��Ү�� ��|���ɝY>�0��������3��-�;�(�>ʁ'?Ǳ>[-�(��=)�?�?�S��e?�D,?S��>�z�=6�������f���?7�*?8е����Nɛ�������m=�`?�ʆ?��+�%!y�L�l?8]??:�<�e�8�����`>gV��A>=??G(?�f��{��>5��?3mm?uN�>���J�y�7���\_q��E=�	u�@��>��g@$�"9�>�?���>�����r�=+�ϼ�e����<�>l�h?�'�?�f}?qɉ>IZ��m���(�"�I�v�]�V?��=�&ԾM�>d`�۵���Xƾ��������`ɾ�����M��􅴾��_.^��9���> m'?k�y?�?��m?,b���u�!y�n@��~�j��(��@�u�U���I��kJ��v���n�n�c~=��>r�S��A��m�?��>:�����>8Ⱦ�d���V徶��>9����{�D��=_���w�<����"��x{�;FZ��?,�>���>��7?��Y��d7�U^"��0�wg���;�=���>L�?>���>$��1{�����3̾g#d�K#�a:v>	xc?��K?ĸn?�j�#(1�����h�!�/�/��_��C�B>�o>�>;�W�~��M:&��Y>�a�r����w��d�	��~=�2?(�>���>�O�?�?Q{	� n��Wkx��1�Rq�<�/�>� i?�A�>.�>��Ͻ[� ����>N�l?��>�>�����T!�4�{���ʽV"�>\ݭ>���>��o>e�,�m!\��i������9�Ly�=��h?N�����`�6�>�R?/��:�eG<h|�>��v���!�_���'�V�>1w?���=��;>�yž"�W�{�B9���J)?<=?�Ȓ�ȩ*��n~>r"?�N�>+#�>�%�?�;�>�|þS�h� �?��^?$<J?�JA?R�>��=�ͱ��9Ƚ�&�&-=���>��Z>��m=y�=���j\��A�iLF=T>�=�3мL���!
<����o�I<�<�3>�ܿr�F���ξ�'&� �s �=$w�}R�V����k�����t�����p�h���
�A6G��
f�--��!h����?���?�>k��������<����@0q>혥�I2��a_˾(�)��٘��A׾�Ƿ�Ɋ�=�B��P��<N�Q�'?�����ǿ򰡿�:ܾ6! ?�A ?9�y?��7�"���8�(� >�C�<!-����뾭����ο>�����^?���>��/��r��>᥂>�X>�Hq>����螾N1�<��?6�-?��>��r�/�ɿb���9¤<���?0�@u�A?�(�t[�T=V �>j�	?"f?>*1�������nb�>e2�?I�?�yL=��W�GO�O�d?���;��F�(>���=&��=�k=b��5�I>r��>Dt�MuA�hܽB4>�k�>s&�����-]�D*�< �]>ջս�.��4Մ?0{\��f���/��T��U>��T?�*�>7:�=��,?X7H�a}Ͽ�\��*a?�0�?���?"�(?>ۿ��ؚ>��ܾ��M?[D6?���>�d&��t���=�6�򇤻y���&V���=q��>{�>̂,�����O��I�����=%���ſ�#�D~!�$�<�����&R�P@ڽ�����R��=����n�kU�j b=&��=�O>F�>6YO>�8W>vIW?��k?Yv�>�x>iq�&�����Ͼ�wc�D���'��O������������6߾����������~ƾ3�=�fɋ=�Q�r����� �+`b��	F��//?��#>��ʾ�M�H^$<$ʾ�M���o�������˾س1���m�+��?��A?Zʅ���V�$���'	�y&��q�W?c����� ݭ����=`����=d�>aG�=i.�B3�B#S��L0?z�?_������QB3>�m� c�<�M,?� ?[T�< Q�>~$?��/�����`>�;>č�>u��>�?�=u����޽��?��U?,��ƚ�.�>m~���q{�0�s=F>��4���� kX>Zn<����=P��~��(�<x�f?")�>��?��J:��ז����=�N1��N�?�	?��D>��?�+�?���=QJ����{�6��lD���W?��?�Q>V�E��#��ʾgYb?�l�?J�o<�V��h=��l�%?r8�?p5&?WRb<��m�<D���'��mX?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?x�;<��U��=�;?l\�> �O��>ƾ�z������3�q=�"�>���ev����R,�f�8?ݠ�?���>��������=�ٕ��Z�?��?����,g<����l��o��k��<ʫ=���H"�!��0�7���ƾ��
�è��Rӿ����>�Y@CX轙*�>E8�6�iSϿ����\о�Uq��?B��>�Ƚ?���k�j�eOu���G���H�Ϧ��$e>˽�=$�<jh|�����-�4o3=Y]>�i>�8,�>fv�4�>�뾯��y	�>��"?�$?C���芞�*�?�:���k9}�Nf���Yh?��?t�y?�W*?�t>i�u�RKm���phn?��?ov?�9����ܾ��5���j?G7��/Ka��k4���C�"Z>w�1?���>��+�XUw=`>a��>G�>M�.�8�Ŀn����B ���?	��?i����>�ۜ?޶*?"��1}��p��[�+�]����B?�@.>�����!�IX<��ْ���
?�h0?�y�Bg���_?F���w��C1�*�<��"�>�g�=��۾-��}��>�X�����*����)�?zQ@[�?�Eƽ�.��T�>���>h.����Y�>��>%L�>sÑ>�gؽƂ�>�n �"5�C��=���?�
�?�v�>u9��"����>f��?���>T-M?�L���@F?�
B>X3>rqb>@������>S�=�?�5_?�,�>����ҾT��MH�R��A�O�J�/�<�>��R?7X??K�L�#��{5>	���_��ǆ��d���,���Yb����{>�,D>�C�>K̽Ka��I�?�o�>�ؿ�i��n'�64?�>��?9���t�)��}<_?N{�>�6��+���%���F���?�G�?��?ֺ׾[̼[>u�>J�>��Խ���\���2�7>\�B?!�ZD����o���>���?��@�Ԯ?qi���?��0؇��(~���O�7�H'�=�7?X���Yz>p��>8ԥ=��v�խ��f�s���>�R�?�Q�?���>��l?T�o�N�B��5:=#�>�sk?.�?�����sD>�?���ꎿ����$f?��
@8t@#^?�Ƣ�q�ӿ+v���a��4����.�Q=8ō>H<���=��>���<�H;���=T}a>��:>2�L>�(t=?��=��=M����v������O�C�(���V0������𘽄\*������߾�OԽ�Iӽ�K�����"�J���
�=�PV?��P?�2q?�>��k�k�!>K��,�=�g%�&֐=��>č1?ǨJ?��(?��=᜾�e��e��XV��>6���,�>#�D>T��>�\�>��>���;�L>Di<>	��>,�=��0=a��3G=-"M>B��>���>��>t><>ȏ>�δ�/2����h��	w��̽W�?����J��1��w9��y���Ng�=b.?9|>����>п+����2H?�����(�0�+���>��0?�bW?Z�> ����T��5>���q�j��`>�* ��~l�0�)��$Q>Hl?��f>u>��3�vb8�{�P�:����(|>�66?�춾,J9�z�u�r�H��eݾT=M>rվ>-@�iW�8���!�u_i�w{=�p:?��?>��dڰ���u�G=���>R>�Q\>��=8[�=�>M>��c���ƽ��G��v.=l��=�^>Hb?Gn.>i��=��>�(����\����>m�Q>�Y>�;?�� ?�M��׽�ȉ���/��,u>f��>䗈>�"�=ϔO����=8��>F�Y>�<<�0�>�'�#+��][>-�ý��V�� ��~:H=�ꜽ�2�=*� =m�� .���N=��?HAÿ`b����~�ꏾ�E?�^?0l����[�U������-D�p	�?�@i��??�2�L|Q�[?�!�?�k�h�=�k�>sfr>/���П��@�>B/O>���;iX�J#�����?���?:H�󒿆��Y�=m�`?6_���y�>�h�[��Q����u�zm$=���>;BH?�=���1P���=���
?�?b�欤���ȿ��v����>}
�?^�?�m��@���@����>���?=\Y?_di>�H۾܃Z�(z�>�@?�R?�%�>E-�%�'���?Yж?���?I>{��?Йs? {�>�.x�4S/�c1��ϕ��W�==�X;xj�>�c>���jeF�|Փ��f��5�j�j��R�a>�v$=��>�7�F5��T<�=���L����f����>,q>��I>�M�>M� ?AW�>秙>�i=�u���ڀ�װ��� L?�n�?�����m�f7�<c��==^���?w4?�w(�yξ���>�a\?�f�?��Y?��>\ ��k��y࿿�e��w�<��K>�5�>q�>�G���M>�ԾJ�D�h��>^�>� ����ھ�ԁ�pN���>#!?��>��=�!?�M#?U$i>���>�H�A����B�v[�>��>��?��?��?�w����5�����P����U�#�`> x?/�?��>�葿�䞿�닼������=h~??^e?��ս�??���?Q8E?�5??e�O>{]&�u��e��i�>��!?����A�bR&�$g��?=�?1�>�b��dֽռ������Z�?_9\?xe&?�F�D>a�}CþAH�<��(���J�9{<�NG��>ܟ>����=�>l�=~�l��6���Z<�I�=�Z�>���={�6��,��3�+?B��%C��Z5�=�o���D��tx>�RQ>�f��,t]?P[9�P�z�/�����ЕT�.��?�s�?��?W���4h���=?^0�?�1?޵�>jꪾ��ݾ�i۾o�o�>2�����7�>��>;�q����2դ��ʩ����˾�"@�5E�>"x�>>?H?8L>1h�>�����
'��Qݾ`,�M_�ޙ��}6���*�[��֒�
��E�k,����p�1K�>6���.�>��?Y�P><_�>7G�>���<��>�T=>Mf>ы�>?#:>��>���=��;~ս8P?<����#�Hؾ� ���?�`?+Ԛ>���ږs�U�)��(>?�Ү?���?�Y>Ђt�קG���-?��?<}����M?�[>�*��3�j>��'��꓾P(����ǾX�>L�Լk�F�KyC�i�����?B�4?�A=`j�������s���}m=�W�?��(?��)�Q�Q�>�o�˫W��S�Ć�Ych�������$�3�p�k㏿�Z��0���j(�sa,=�v*?F�?�j��A�Z���0k���>��^f>$��>cϕ>���>8�H>��	�	�1���]��*'�!���jb�>@{?у�>��I?1<?�vP?kL?���>#[�>�(��_h�>+�;-�>U��>1�9?��-?�30?�w?�t+?�7c>l�������c}ؾt?!�?�G?C?ۧ?3Յ��oý�ۘ��g�	�y�������=���<��׽�Zu���T=HT>�`?����>��0��6y>Y�;?��>&��>�~�����I�X=���>\�?�ψ>�]�*�u�=�����>�g�?^��~I=3y>���=����<E�=��W���=��9;7����B����=-�=��;Ez<�\���
6���x9�L?.�?�D?D~�>�����-�����Q?K/;>6D�=�{U>j���"?���6��,9X� '8>!:�?�k�?���=J��>���<��c׾]�=�h*`��/w>���>+�-?2%H?��?��_?��?�z�<N�6�����$e�}7ƽ�/"?u!,?���>�����ʾ��ω3�՝?_[?�<a�����;)�ڐ¾��Խұ>�[/�c/~����3D��녻���N��2��?꿝?=A�J�6��x�տ���[��u�C?"�>Y�>t�>W�)�w�g�l%��1;>��>cR?'�>��O?�{?�[?�rT>��8�3&������2�F��� >5�??���??֎?$3y?G��>��>�(��ྴs�����W�*�ܲV=��Z>86�>���>�v�>::�=A
Ƚ�[��)�>��v�=cb>H��>Aå>���>�hv>��<��??_��>蝾��G�<m��J�����?z�m?�m�>�8%=�5�I�F����+�?U;�?YH�?�5�>������= ����o��]�����>��>�D�>ϭ�=���=��>�I�>���>�D��b"�n�+�2���/?;�5?��`��ѿ:�j�|. �2�������ٜK����(�=��G`>2���^T�T蛾�f����]ɂ�����e����r��g�>3I>ߧ�=�������y�,��ż�?7�=r-�6`��v��ꏽ�L �<��&�t]�<-"�<=�E��>@<�Ⱦa�?��?��)?�#?ܲ?�6�>����f�N?����d?�|>��=S��Qaf����W
о_�q�#վ�E8�\@;����=��y���=�%A=�Ep=�%>6�@=屭���=Ӟ��ҏ�= XC=�p>޶m=��b<�&�>9I8>�]j?��i]���;�����/?]��>�w%��{Ӿ��a?�yX=������&Ծ���?\��?�I�?"]�>�o��2�>�����M��=ԘT>o�b>�`�=�m\���>%�>HEu�⹘��rн,~�?��@r� ?E��b ſ�+�=��=>i`	>;�O�L�1�T�<�Gx��Po�|�$?��9���ξeԄ>֋�=�X��$ƾr��=�hM>5��=��&�`�\�|�=7����hB=��z=���>�4K>�޺=\E���	�=e�=�l�=��Q>^H-�m�s�e�2��i&=��=Ɲ`>�n>,�>�z?p�?��J?$��>]�����^���P�x�ʽ}�>�m��qr�=Ol�>��J?�b?�)U?�C^>�(���>ɮ�>���[�{�E�#a������l�?���?�>R�=�۴���
��U�S�C=�Z?Nh?
�>N�>���qwҿ�-�<�*�	X�9;���@�C�S�E5=���=��"���ǽ��^<K<�>�o�>`!`>ɭ�=b�+>��=Tޭ>�2>ʿ�<����R+=q:�=u���,=�,��8V�������X��(�;�O���	���ނ�J��=�%I��/�� �=�=�>�v">A��>���=����t�>2����J�2��=�0����@�EWe��'}���,���-�kJR>�a>h���OCn?x�h>�w9>�@�?�v?�=>�c���g;eڝ�*"`�5kP���=�^>RvF�? >�A�^���J�M�;��>���>�5�>��k>��+��?� �v=U�e5���>،�V����q�=$���៿��h���b�a�D?�5��^w�=�~?ΞI?֏?4��>VB��I7ؾ�0>������=4�%�q�&��;�?��&?���>h(쾡�D�ɓ���l�!�>9w���l��9��OB��������>��ܾ����<�?Q���T��X����e���>�BD?�V�?v)����V��C�� ",��S����?)�/?Ŏ�>i�?�h�>��M��+�S�^���==��?��?���?Tt�=�R�=l������>�?��?n��?G�r?�?��d�>���;Cw >�������=B�
>i��=�S�=�2?W�
?в
?��	�u%�	��՜^����<��=���>��>[s>�-�=�Sf=�=�[>�!�>��>�Id>nj�>�D�>�[��M7�ȷ)?���=ݽ�>c�.?,r>�1-=�-½�2=���%<L�!�{��4jѽE�<6u<ha�={��7��>�eĿ��?̹U>��K�?d0��
q��{W>�4d>�A��(�>D�->f�`>Q��>HZ�>>z�>��>{KӾ�{>����g!�-C���R���Ѿ��z>眜��	&�^��0{���AI��m��gf��	j��-��==��Ž<H�?ǥ����k�"�)�������?�T�>�6?4������(�>���>{ō>�I�� ����Ǎ��eᾰ�?|��?K8[>?>|�l?\��>�����ھqkV�Pu���l�\G��D��ҙ�)'`�uY�� �<3V?��o?��P?b;=�qs>$��?ITJ���(�݆+> }b���~�]:?8�<�I�ULY���i��ǟ���>���>���?��e?FL<>���\� �3�>�N,?�q?<fi?��8?F�5?��$�_�0?��j�?(8�>��/?_�?)��>lp�=�()<�s�=�G�=[&�]6���<��b��ȓY:k=y��<-�}�n���x=�j�<�.p��4���ڳ��㯽퀈��t'=:
�<T�=o�>6�7?v��>Ы>�FN?SkϾ{!`��� =_��>߂>n�.��m���8����!n�>�Z}?¡�?�E?����V:��F��茍>>w�>�����>�T�>X�����1&�<�m>C��=)]n������羂��ࢃ��P�>�Bl>���>�M->�*=��n=�(w��Tt��#>-p�j�ɾ��*\�$35��j9��ܯ>��D?e?Q
>㟾"*[=�yW�~?<T;?�C?d�}?�p>,�	�b��b+�T_!��>d���J��{���М��J:��ȯ�m>�z��Zܠ��Sb>����r޾z�n��J����M=���nV=�� ־�2�^��="'
>-��� � �8���Ӫ�1J?��j=}x��@UU�yt����>A��>��>0;�:w�)�@�$����?�=5��>);>�<������~G��4�3�>�C?E�^?���?����9�t��V@��|��D��<����I?�ۦ>�F?��S>�=�N���\��c���A��r�>�&�>�Z���C�gş������$���>$�?�w>J?�WO?�	?�zb?��(?�^?y��>4e˽Ax����?�y?+hݼQ%���=f(g�Bfb���?�?ӓ��6@>Ia�>���>�?9�?��S?5b>M�N�����[>浕>��B��㠿0��>hh?�#սa`?�p�?^��=_����Ua�э˾���>�8?f#?�0�>��a>���>í�� 7�=��>fc?�+�?��o?2$�=��?�M2>v��>0��=	��>���>	?�OO?�s?.�J?'��>6��<�?����#s��O�yc�;��G<=jy=���
�s��0�
��<�p�;醷��L��/�D�������;�g�>��>l[���8�����vg���z�>t�O���ᾥჾ,C��	�����>�X7?L!�>e������>�D�>�pB�[�7?V�?JG�>��>�Xu��ݾ�䟾�>ӡ?ǋ�>�P���ʦ�.�h�͋�=��w?��p?��;�E#��nc?�nZ?$���=��k��OiL���C�O?��
?t�<�P�>"~?�q?f��>�lo���n� ��)ba���i���=��>�7��`����>ى1?�y�>��]>a8�=�Ͼq0t�#ǧ��1?a�?ee�?��?��4>��n�Gl�t�.�Ρ����e?F��>�����X�>阽����6���Gm�A �����󯾲e��q��G���h��U.�ƌ�=��0?>�{?�J}?��Z?�� ��m�|Rw���N3P�VuҾ��$�D���?�,;�� G����2�U�݄���<�s.�T�%��v�?/p�>`m�;�;\>6fr���߈��>@�Ӿ�����g=)��=_D�=���=����2���]���%?x��>*�>QuQ?��z�_�X�ſ�����$V�2���~�>yԦ>	�?-�>=�@=�7g��+a�p�����=t-v>
yc?�K?�n?`z�E%1�-���L�!��/��i����B> {>���>F�W�����9&�X>�?�r�G��+w����	���~=Ϯ2?)&�>|��>-N�?�?vy	�{i��gx�4�1�k#�<�)�>�i?�?�>i�>��Ͻ�� ���>��l?���>4�>����Y!�K�{��ʽ�"�>�ۭ>&��>�o>��,�R"\� j��܂���9�Ex�=Ʀh?B�����`�[�>�R?8*�:�G<<z�>J�v���!�����'�R�>�y?j��=�;>�ž/$�ʣ{��1���&?-�	?����E-���>��?���>h�>!'�?���>�ž�N��%?��[?��F?�&<?x��>m�:=,Z���S̽�W)���X=)܈>5�b>��T=��=� �hg]�-����S=M�=�����Ľ�[J:���v<Ӹ#=��9>��ۿ�K���׾���9����	�C3��պ���?���o����t����y�#%�{x,�ѷV�Vc����/k�5&�?ߦ�?fm�������M���Z�������L�>l�s�7�v�8��ؗ�������߾�{��� !��HO�o�h�:.e�V�'?�����ǿﰡ��:ܾ>! ?�A ?9�y?��<�"���8�{� >�D�<�-����뾬����ο�����^?���>���/�����>ߥ�>>�X>�Hq>����螾<1�<��?0�-?��>t�r�%�ɿf�����<���?-�@�~A?*�(������U=C��>ґ	?��?>�81�!F��谾Z�>�7�?���?;�M=7�W�$+
��je?�L<C�F�$�໹;�=�<�==����QJ>g]�>�o�3]A��ܽ"�4>���>B�"�8��7U^�Mֿ<;�]>z�ս礕�2Մ?A{\��f�r�/��T��U>��T?�*�>�9�=��,?Y7H�]}Ͽ��\�+a?�0�?��?�(?fۿ��ؚ>v�ܾ��M?^D6?���>�d&���t����=�5�(���j���&V�m��=ʬ�>Յ>��,���]�O�2I�����=W��{ſ�"��a��|A<Iw������3н�CK�w��E��^����`�<�E=��">p%j> �'>�xt>�S?O�U?�;>��)=I���cZ��,�����=�X����J:���(��ϓ��v���Ϸ�����t,���D�.��w=��)�=	2R�ʔ��ź �U�b�2�F�+�.?�W$>>�ʾR�M��+,<�oʾ~���*����a!̾A�1�`n�ȟ?��A?������V�X����ӹ���W?�� ���ꬾ���=����=�9�>	٢=���=$3��|S��-?��?���A^���>d� �ߟ��^22?|��>��<r\�>��?>e���ὴ�V>
_>�ϳ>ɤ�>��=� ��`m���>?,Fa?�EP�����"��>O���䁾�kM=k�=� /�i�3�(�J>�;A������g��x����[V=�Xo?���=��"��7/�p���~�9>�>Zy�?��?�:���?-�?�:�>�)��@���.$�����8�?��?H�O>قžQ��J쏾C�P?�'�?�<��nU��4��N'����o�"?�hm?,](?
D�=)ԃ��=���ƾOUP?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?p�;<��P��=�;?m\�>��O��>ƾ�z������3�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�ٕ��Z�?{�?m����>g<G���l��n����<`Ϋ=���E"������7���ƾ��
����{޿�ӥ�><Z@3V轂*�>	D8�Y6�TϿ��\о�Sq���?6��>Q�Ƚ[���/�j��Pu�P�G�4�H�����<�>���v�=�:�J����*�Tss=5'�>��۾U'?u����)�q�&>y�)?>�)?z�/>GM��ڍ�?7��L�h�}������?"��?���>�p�>*��<pBۼ��s<M�;�\I?p!u?�S?��3��t����,>�k?o�����`��{4�`�C� \>��2?RP�>6�+���{=�>�q�>�D>�.�LĿM|� �SS�?1(�?�k�]^�>C��?Gs*? 2�;ۙ�7j��n~*��Me�HLB?g=1>��þI�!��s<��ɐ���?��/?|w�qG�%_?���m��e��Ξ��6�>y�O�����`뽔�">��\�md���I��ۃ�?�~�?vɥ?�#����B�B�?�`�>#�$���W���̽��7>C �>��>g�4��P�>��Ѿ,�l�A��;��?���?e�?����*��߱�=bt?���>��M?s���lq]?�β=��N=;��>7B�<,��>|lK<�1&?��,?]�>s�M��Y���x-��(Y���A�r��uw���?�`9?rLQ?�Q�<��$�����F'��=�<�ǾҸi���Eʰ��NI�Q>�>�/�>E��1�����?Hp�5�ؿ�i���o'��54?9��>�?��R�t�����;_?mz�>�6��+���%��&C�P��?�G�?#�?j�׾�R̼�>F�>�I�>��Խ����q���:�7>&�B?���D��g�o���>���?�@�ծ?�i��|?å��������d��#���>�l/?Z:�����>?��>s��=Cw�W����{n�Z��>
հ?�0�?�j�>�2r?�x�L�M��J�=�N�>JOo?>?�N�k��
7>'�?em��v������|Mg?��@�A@v�X?�a���hֿ����,N��/���-��=#��=h�2>��ٽ�_�=�7=��8��;�����=�>5�d>�q>X(O>(b;>L�)>���8�!��q��Q���:�C�������Z�X���Wv�_z��3�������>���3ý�y���Q��2&��>`��>�=��U?!Q?<	m?FH�>�,O�V&>�a�� �=>�4��=��>��3?�1H?��'?�n=�O��m�`�,)��B������Dq�>�R>$��>���>��>��;��G>�>>x�x>2�=D&�<�S�	!�<e�U>0�>e%�>�H�>�C<>��>Eϴ��1��e�h��
w��̽1�?{���T�J��1���9��զ���h�=Kb.? |>���?пd����2H?%���y)���+���>}�0?�cW?!�>��L�T�1:>9����j�*`>�+ �|l���)��%Q>ul?\�f>��t>�\3���8�qUP��m���|>O�5?z��k`9��u�3�H��Gݾ{kM>Ѿ>23H��K�Hږ�
�~��i���z=��:?^g?�ɰ�����u�'����^S>��]>b�=�"�=�wL>&.g�)�ȽZ�H�T,=��=�^>f-?Z�@>�R�=��>9�����S�u��>R�a>�
>9�9?3;?с|�|�齟&����)��z�>�>�>G7�>$_�=*#b�B��=���>�_s>sA� ���n��1��N>Ef����n� ���q=/=��<�=���<���JH�EB�=��w?v��œ��������S?8�?LXQ����PV���I�������c�?#@oЖ?�����U����>� �?q*��̙>��?�o.>�P���9����>��x<�f��m�;�������?�V�?�|�젒�1�k��X�;�c?�0U��o�>�y�3Y��B����u��$=���>*;H?�O��3P�h�=�5�
?r?=b򾵪����ȿ>|v����>��?���?C�m�e@���@����>£�?�`Y?P^i>�_۾1fZ��}�>ѹ@?fR?�&�>�3��'��?ݶ?t��?�I>c��?.�s?Wx�>�x�>L/��,�������=�~P;Q�>*>����h\F�ӓ��_��1�j�\��_�a>^�$=��>��GH���F�=�L���7���g�|��>�q>m�I>N�>�� ?L�>�m�>�=�k������z�����K?娏?���f*n�H��<��=��^�_1?cG4?��Y���Ͼ�Ҩ>�\?b��?x�Z?X\�>����=���ڿ� ���7��<�K>�K�>�N�>�Љ��ZK>��Ծ�D�\��>	��>e��LNھ�=�����W�>�o!?���>M֭=�� ?*&#?8fm>~ó>h�G���Z`B��w�>d��>`L?.l?�h?;�����3�}�������u�W��1[>��w?"�?Z��>3I����P:��LGD�[#d���?�gg?��ӽK?4��?{�A?�/>?��\>����ԾỊ��b�>g�!?�K�
�A��R&�/��)?
�?Y#�>�H��?Zؽ�ؼV�������?�x\?A�&?T��wa���¾�<�$��#W�Aw�;�J6��->��>����>]�='0>�)�=p)m��P6�FR<�ɼ=�d�>��=��6���-)?s��<�-��E�>��q���@��_>��o>�d¾.YX?��G�ơy�/���yИ�N:O� O�?���?��?��㽪�i�ʀ;?���?Zg?u��>�G���Iʾg�ԾD�n�Z#�������=r��>�
�vA뾢g���§�(.���y������Լ�>=��>�`�>�i�>�>�-g>lX����������b!h��@"��T�X�����Ӝv��	Ľ�h�鮻����H��>�����>`��>K�&>�0>&�>�ʃ=���>@5,>hQ�=�fi>��?��t�=)P�=	#�=,�<U`?�d龺G�VN��,K���{g?��I?���>�\�=��H�������=?���?1��?u�~=���a�g����>MA3?{���8?l+�=!�?�Z��=J}����h�M]�N>G�D��>L�h��Ox��l=��{]���?��3?A|@=���� ���7�t=Cp�?��(?��)�1�Q�ӵo���V���R��Y���h�N"��Yb%��Ap�\�]������J�'�3z*=�}*?
��?�(��7ﾄӬ��5k��e>��e>-��>[�>s��>��I>��	�1�1�YU^�߸&��a�����>	P{?���>��H?��;?�
O?�L?6��>Ҧ�>b&��R��>��; ��>�`�>v�8?-?��/?��?�*?6c>(w��J����bؾ�k?�*?��?x�?�?b���P��<Jj��f�By�����x=��<��ٽUpz��\=��U>�,?��k�9�����n>�0;?K��>y��>�Ʉ�oV���9.=q�>Y�?t��>���[v��I��"�>K��?v �ߥ�<7�>�~�=W�d�Y����=�μ�Y�=>�8�9.u�')�3��=Ս�=2T�;����u,����T��f�<lG?�Z?�е>� �>��ݾ�L	�پ��w>~p5>�>�n>M������͏���}�|�V>\^�?>ó?Qe�=��>h"z�i��%ݾh"�@(�����>�x�>�#?��P?�Ұ?_�f?
�7?)�H:֭#������YW�3�x?`!,?���>v���ʾT�w�3�Ν?[?<a�Z��m;)��¾r�Խޱ>�[/�>/~����D�� ������~����?ڿ�?�A�I�6�ix辪���7[����C?�!�>�X�>��>U�)�K�g�2%��1;>��>�R?�Y�>r�N?��z?�|[?��R>ë9�zQ���i���縼��!>��>?A΀?���?�Bz?F�>��>��&��߾I���/��o��#���uf=��W>�>+��>�j�>�8�=�νW���G�@��!�=�kh>Һ�>�E�>�x�>t�q>���<��4?�?$:þ/>$�jI>���;��6�?C�?CF�>d�ۼ*��X�?�����/?͸?��?�Ew>ļ#�< �<�w�|n�C��_�K>���>�8�>�b=�Z�*��>I��>��b>W�8�d�侰e^�7���>?�Uj?�z�/�ҿ��w�
�R��ɾc��=������d������F ���>���$���\����j���bT��M���[�;+�
�Y��>+�|=hv>�l#>a��<7ཀޙ;�����5���>���9��<b!��Z��/ƽq�~<+?O=��F<�FW�A]����?�n?]!?�{�>�1?��|>��<�o!?����I@?�r�>:�>��ľY��8���S�c�V�]��	��\����=>�F?�9.U=q��<y��=j�=ค<�m�=���<�0������.�=D�=[��=1O�=O�.>�J>��a?�g���(��W%�so���*B?�"?d�����d?��>��[�~h����޾�	v?*��?�N�?�}�> @�d��>�>�U��� �>�C>��<h+=�oH����>��=b�ѾE珿����mY�?�y�?{�?����?iĿ�z�=��7>8�>�R�S�1�R Z��&c�tq\��!?l�:���̾ⵅ>7�=�>߾0�ƾ�17=�7>��d=��y�[�Q�=�{�,G==D�i=2$�>U�C>C�=�Q��?��=�Q=��=�/O>����<��y/�2= ��= dc>m�%>��>ժ�>T?��V?�[�>F���������`5�{t<$�}>��轂/>t`.?g�7?�pG?Մ??R1>>��>{��>F�9�PS�R����˾)Zս���?��?`�<�%�=�:��O$���-�)O�<�7?L�?P�h>�A>K��L�ۿ�{�u-�1!T���P��i-�i[�b�<dSX����㒚���D=��r>�!�>�u�>/i�>DE�>�s>��>uQ{=Y��<.^�:�`����=<Q=���=��ؽh�<�6�������;�K�;#ǚ�cgʼ�j�������<;'�=SO�>_K >���>��<������>��M��*G��Ρ=�䱾}$B���g�<�v���&�0���%]>I�P>�GȽ
򐿯� ?|��>�,>E��?uEi?p�>�F��:mȾ�y��F{��Y��#�=^��=�q��VE�^�(H�
������>�>��>`Vl>��+�r�>���y=M��u@5�T-�>X*����һ��q��7��B�(i��G���zD?%D��4�=V~?��I?�ُ?��>"��Hyؾ��/>����K�=����q�9���~?�%'?���>����D�e/#��%���R?�:,���h�H���ڨ`�N��<I����?RZ��v��v�g�~y��
(u��-߾�il>%�&?X	?f��?��ý�^6��;��@�s�.�C�>�E?�U>}M*?uo ?m��d�þԯ���y�3�u?���?o�?y�<˷=.޼��/�>0� ?��?��?�n?��Z�6��>�I�<S>�yǽG��=��>5��=�
�=��?χ
?XY	?N���M�8g羈����Q�f\�<
 �=~�>� ~>з�>i��=D�s=ݍ=��S>8?�>��>#�g>䳥>���>�]����	��(?X��=�B�>��+?�x>bM�<%�����=�2����Z�"�5��g��(����o<�$λ=?������>�pÿ�-�?��U>S� �	�?.?�UgY��@>�n>�xν��>��5>Zqq>�Ş>�?�>˔>|��>A�2>�CӾŀ>g��Zd!�8)C���R���Ѿ�wz>ʙ��V&�b��+����II�=l���f��	j��,��B9=����<�F�?����m�k�n�)�G�����?�Z�>�6?wԌ�3�a�>���>�>L��Ɛ��Ǎ�Bg�[�?���?��Y>�&�>`A\?
/?xȼ���I�U�T�	�t��X9���K�^�\���3��/3��M��S?�l?�T??'$ =���>1o?��������D>չ3��(���=��%>P��Mai�l���dܩ���ƽ� E>�o?̀?b�?e��mv��p_>�c9?�c%?g^b?jL1?"0?��N*?��
>��?�?.l6?�� ?^�?��=�n�=�˰<�}��ㅽ|l���U���L��d8y�I�<`��=�\����}�0=�^=i�;2*��2�<zb'�x��<[B\=�+:=F��<1 �>�VU?z�>�.>>nw??��H�Z�n�9ZV��k?�׻�Y���?��`V���뾰o�>��~?���?V&?=
�a�
%F�:�;>Ν�>!�нkBm>E��>�_ͽ�����n@>��=��=�R6���<4�����t[_��o>k�=@��>�O6>Qp'��}���7�{��~�;>�}ܾਮ������A���L�^�7�oJ�>k(I??Ǎ�=��˾@/̽m�_�v�?u�I?�?�Џ?��>�NؾU������7�z��Ņ>�Ĉ�9�.��j��+)��Kc>�_zO��ch>���ɠ��Gb>��Z{޾{�n���I����p�M={��V=�'�վ#*����=�
>����v� ���XԪ�R(J?�Hj=r��@8U��a���>;Ø>�ծ>m;���w���@�����"��=Ц�>)/;>�9�����f{G��@��-�>�NE?V?_?�~�?*0���s�p�B�Zp��rS��%�ʼ��?��>�5?��A>���=����`���d��G�7��>ک�>Ƶ��G�V+��Z��ĥ$�s��> ?�>�?��R?g�
?4s`?
�)?�?��>�����׸�f�$?�?
�=��ཾ�F�s�8�I�4�>e�&?F�T���>��?O9?d'%?4/Q?n?7�>+����TB��>�>���>��U�sկ��xj>M�I?\��>:9Y?	؃?�A>j6�´��1D��Nְ=1>j�1?<6#?��?7�>��>պ��,��=�>�>I9c?%��?b~o?T��=l�?�2>���>�@�=�>�C�>M�?��N?�>s?��J?���>XӇ<Â��������v�n�H��*�;̦<Z.x=���ul����!9�<"�;�C���={���Q�J�*L�����;��>�2i>����R>8���l���?L>��%������2���nY�`Gy=�j�>�_?�$�>>K� q�=��>�3�>�0�%�'?�6?�N?ka�<�G]��n۾��3����>�a=?Zz�=.j��u��2x�zz= �f?��_?==E�k-���b?v�H?m��|>��B|�ŕ�:Ҿ�L?��?�	��&]�>#��?�r?��>Ӌ�rkn�}e��H>u�]�C��Z=�Z�>f�	��\� ʣ>��?�>n�$>Sq�������i�7���^��>�x?l0�?�Ȉ?M�^>L����  -��N��H	r?��>�V���?����[5���P��ѧc�>B�%���E��󑃾�)���x$���u�\ۈ�G�=8z ?'܋?��t?�PQ?)����l���l�s'���W��ؾu�����8�57��R�}�x����U"־nXk��]B>$�{�1h?���?��!?Hf"���>^�����nN˾wDI>�)����!�k�=�G��?pF=:�:=Dh�wx&�d<���+?cj�>�2�>�r>?f�\�y�?���/�&8�����0/3>[��>w"�>��>p�:�&,���ͽjm����r���ǽ(8v>7xc? �K?f�n?�m�$*1�ǅ��ɘ!�(�/�!c��,�B>Bm>E��>�W�u��{:&�Y>���r�&���v����	�Ҭ~=گ2?|(�>�>�O�?r?>|	�"l���gx�[�1�'t�<�0�>Wi?e?�>�>�н�� ����>~�j?���>t��>֣��u�+��w��	����>��>V�?`�U>��@��,\� 捿nK��)R+�6��=�Kd?R����"o�Ԭ�>"�J?S=����)�>ƣ���:���Z���,>�F�>�9>&X>�־��	�Gق�(qx��3(?��?�됾�8+�*_�>A�!?!��>ڰ�>*t�?~��>lľ��ݻ�a?��]?�I?��??l��>3t=U驽U ʽ]'��/=���>�6Z>�}=s�=����6\����/�W=���=Q\Ҽ������<Q�xd<�u�<7.>xۿOK�j�ؾ�����0*
����������f��B��s��w����x�����(���U�&(c�ބ���l�|v�?a=�?g������(���������a0�>�q��
�Qͫ��(��4�����d���p!�g�O��i�te�P�'?�����ǿ񰡿�:ܾ5! ?�A ?9�y?��7�"���8�#� >|C�<-����뾭����ο@�����^?���>��/��q��>ޥ�>�X>�Hq>����螾I1�<��?6�-?��>��r�0�ɿc���c¤<���?/�@��A?I�(�i[��P=�z�>k�	?4�?>�&0���%��`�>�)�?�Ί?e]O=�W��_���d?弙;��F�*�軄��==�=У=���n�H>m�>��(B��9߽})4>Bu�>+b/�����[�~F�<
�]>X׽�f��ʶ�?�\�̷e��x/�^����>U?`��>�=A,?@I�TϿ�:Z���a?�?�S�?h�'?�¿��>'ݾ�N?��5?��>�e%��qu��(�=��лN���U����=e��>�E>��,�-���!O��Ņ����=�����ƿ�V�������<L{<�JV�����Ve��#�+�+ا�?�]��g���3�=6��=u�U>��x>�T>|y2>|
U?~Dn?��>��D>����,���ܾ(���-��9c#�\����4�/h�����Ɖ��������+��C9��8=�&�=w4R�U���½ ���b�ʚF��.?$w$>{�ʾq�M�{Y-<�qʾ����:ʄ�ſ��9%̾Z�1�D#n�(˟?L�A?������V�$��jW�Tx��Y�W?0D�����笾H��=�򱼝i=��>���=��⾂3��{S�z�0?�C?��¾���(6>���1=gE+?6F ?mN<�]�>�7%?Վ-���߽[>F�)>ʢ�>C��>I��=D����^ݽ�?�xV?�� �����3�>p���w��1=s�>"V6����YFV>���<}���EcA����F�<e?Z?��$>f�.�r��4:̾kĽO��>�A�?i�>�-?>���? ΅?)��>��B����H�c]���R?	,�?Ƶ9>uGٽH���}Ͼ*@U?&͗?�T>B�)�H��a�L�@�L�Gm?�$z?�q?��.>]Nu�/��Hg��W?q�v?Zs^��s��u���V��>�>�^�>��>��9��p�>��>?�
#�H�������Y4��Þ?��@ۍ�?p�;<r����=o8?�b�>o�O�=ƾ���%���׌q=i �>Ћ��&ev�*��O,��8?⡃?��>�������z��=�ٕ��Z�?X�?*���UFg<P���l�vn�����<�ͫ=��F"�����7���ƾ��
�ʪ���ݿ�ͥ�><Z@�U��*�>�D8�Q6��SϿ$��(\оrSq�e�?��>K�Ƚ�����j�DPu��G���H�����kD�>�>�ؒ��y����{���;�ȯ�����>V��Qu�>�R���M���.<U��>}A�>A$�>=>��Ƚ�]ə?���=ο,���S��f�X?qi�?�+�?Oc?\�B<�s���z�g��{�F?D�r?�Z?DQ%�s[��5;�r�j?[���X`���4�[3E��iU>@3?�O�>*�-��8|=�6>T��>z�>/�+�Ŀ�ڶ�������?���?jn꾜��>z�?�a+?7[��1���]����*��H�=UA?&�1>Ѩ��s�!�&=�ϒ���
?uz0?|��{A��d?�΄��땿�����i-=�Y}>򇧽�-Ⱦl�t�t�=�WY�	n����Y���?�2@֛�?>wӽA=1�� /?���>.�}��^`��2�f�7>0Ȧ>>"V��Ķ>�@��W�_�*m�!��?G��?��>e������.2�=i�?,�>�8?�W�OO?�vS>�}�����>J/�_y>�_S�|x�>�iX?��`>��>���&4�[��/��d&�F�1�[h�>nC?k�_?3���n@ʽ�h�<Ȉ(�_ښ=d������;O��=�v��a:�=\^>�n>���F���?Mp�9�ؿ j�� p'��54?/��>�?����t�����;_?Qz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?[��D��u�o�y�>���?
�@�ծ?ji�L�>�p��Y�������a<�!���	�>#O?ɴ����>v��>}�=*���S����z����>�D�?�s�?�t�>�"�?�ⅿ����(ب=Q�>Q�?ՁJ?8�����Ͼ<�c>x7#?�����|� i��.=?��@��
@>�8??���ܿ%6��¤������\��=�->�A>+���X=?��<5@�;�:�)A�=��> &J>	)(>�>'�>oZ�<F����H&�:V��!ˎ�I00�o����"ހ�x���މ����*ʾ3wԾ�[G��?&����1/w���|��=2_?��H?�݁?���>�s8��uD>Q� �=�8w��f�=�}�>53?uA?�f ?� <�`��#m��v�w��|M4����>�_>�>E�>��>L@�=?�G>�
>��>���=�0�=�!���I=98>5��>p �>���>�L<>Ӌ>�δ��0��R�h�(�v��̽���?#���G�J��.���2��㤷�Zn�=�_.?|m>���?п����#/H?����'���+���>ۼ0?�bW?��>��� U��5>���l�j��X>� ��{l���)�o Q>hf?��i>��q>J4��7�]WM�r签��}>C�5?�򵾣:���s��F��޾�L>��>X����a��|��g�~���i�$�{=�e:?o}?=M��hձ��oq������4T>E�U>�'=6��=ԷH>��h��>��'�F� 11=���=`�[>��?P�*>� �=���>Ѡ��U�P���>�|C>{p+>��??~�#?� ��������5�-�1�t>/C�>M��>%�>8RJ��H�=y�>q`>�;�/O���"��?�UVU>=�n���X�A�o�rZt=�E��e��=K�=�4���=���=�gv?�Ǭ�EՇ�t�پX@��gC>?�*?���������^�`�������?J�@�?����~�L���>	N�?���C��>�?�1>]���|���?4�w<y!�ʽ��Z����?�f�?�_���V\���)�P�`=g'?���Dq�>`u�AY��Z����u�$=���>S@H?XQ����O�?�=���
??=[�ԩ��|�ȿr~v����>g�?��?��m�R>��{
@���>���?W]Y?Uai>�S۾'�Z�$l�>}�@?�R?B#�>_/���'���?Vض?筅?aI>���?`�s?�n�>�3x��Y/��5��疌�ty=̍Z;be�>�Z>�����fF�nד�ah���j�J����a>ߐ$=��>�A��3��;�=. H����f����>4)q>��I> W�>�� ?�`�>]��> r=7k��}߀�����L?a?�?�`�i n����<���=z�]�s&?��3?v@���ξ��>[9\?(��?�IZ?�ђ>�P�]�������8N��i/�<�5K>*��>!W�>�Ѝ��L>��Ծ�aE��D�>�6�>�Z���rܾEb��/�s���>�*!?nj�>T�=� ?�??�|>�:�>�fY��s���3�V��>�m�>?���?��?g�Ѿ�/�5���Ú��QB���v>�Je?�?U>&���י�&kē�R����l?��d?��ϽƔ!?睉?L�F?M�0?�<Q>�-�����r����Έ>��$?e���-H�_*(���+�ӓ?a ?���>�u���P���,�;�>���龦�
?��K?6�?hV��Ls��)оX_/<,7��{�:y��=F�<�f�=�/->����S�Q=o`V=%�=���1���S�K��Y8>4 �>���=m >��2��(?�/�<JTj����=%�w�,YL��V>��>l���(�\?���x����>՜���b��و?=��?T�?Ђ��	0d�b/?p��?O�?�K�>�Ǿ�\Ⱦltþg����r������>��>y1K=	N�Q���Vͧ�z��fB�����>�K�>�4�>Μ?}L=>}ϲ>M򃾘��kԾv"�`Id�X�t'����z�㙾4��21=�ɾǁ��ӏ�>���p�>_ ?���=��>�
�>���=�(�>P�V>�[>��x>k@>�ǰ=~IC=��U�»�j�W?�8��X�6�0�۾�Q\�,�]?T?�a�>�ك<wUn�H5Ͼ7PE?�b�?��?��>kdr��lN�h��>��$?������?��F=�ʧ����=�iľ�G6�N`0�7m�.t?�8�n�T�̒D��v8�
G�>0,?N�(=���p��||��=r�?b?.+��tO��T|��pW��"R�2�H;�0��Ɖ��M�'�"q��Ԓ�y���u��;�G�=�{8?�U�?�[־]��fǦ��z�d�H�� A>#Ǚ>�>��>�\�=iX��F���Q��_"���a�e�>�?t}�>�{I?k�;?�_P?noL?T��>�f�>r&��,e�>C��;�ܠ>/��>�9?i�-?10?�p?Fh+?6c>s��������ؾ�?C�?�F?�?��?w���{/ýA���a��y�>���ng�=p�<5ؽ��u�KCT=,�S>�E$?��&�F�@�J�F�>| H?@��>���>G��D��4��=��?6??��>^� �����L#��M�>Sd�?]�� �X<��>�>��8=V4�=`u~= �۽}>u�뻔�����1�=�>�M:=H�;t�cg��dSۻAL�>2P&?�2�>ދ�>W�ϻR��;���?�d�>��>9��>��˾UJ���I��k�q�( p>䁑?iۦ?�N��b >fE'�8b������8�\���B>W?L�>�?)�?�V?���>��\>+������x�g���b����>z!,?>��>�����ʾo憎�3�ܝ?HZ?<:a�Z��:)��¾� ս��>Z/�/~�����D��݆�r��	x�����?��?t6A���6�*t�?����W���C?V�>�X�>��>(�)�t�g��#�5;>���>�
R?��>��O?D7{?)�[?<hT>��8��.���ҙ�m�3�W�!>+@?���?k�?�y?6y�>X�>B�)�N��X�����h��߂���V=�Z>���>��>��>��=dOȽ@����>��a�=�b>X��>��>7�>�{w>�h�<#�5?E�?�F����!�I�z�t"��ׄ{��\?0�?��?ՒL������C�����b�>ӊ�?vP�?�$?.����>�t3�؞����X>��>�:�>�g�=���=�PH>�a?KѠ>j�6��P��+�q�@�+� ?ۦH?D��=�I���Gh����<MʾŢ>��B�[��g,��WdB�X��=ǧ��n�?���-��Y|��|���-����K����>q��=��>;�=�)����Ar����8-�]R�=2��d_-��0R��μ�\���ɼ�	=���=�����ܾ��?�SC?C�\?�b?�?�>?N=?�Z'�x9?�i�>��>�A��l�=P���N��p��nپ��y�"�þ�>�=R�T�Z�>�	>M�k�1{�=c
�=O-�=;2�=׈?�L㸼Z�<��>�J�=�Ԩ=~{�>��P<vn?� ������#
�F�����2?���>�m�|%�do?���=A c�[s��$��!c?�n�?���?���>f|E�;��>�`�5&m�"��>�>��={<��E�c�m>�<��������<�=�v�?%@m�@?����s~ۿ�(>d;>��>��R�D51��ZO��]�ǾY��	!?��9�2>˾�>�a�=F߾��ľ�4=�1>��G=2�"�_\��V�=�@~�a�E=���=�>�T>>.Ǽ=��� �=��)=���=K)L>h�S�I&F����1=F��=�a>� >j��>S?�3*?>TT?ߛ�>x4��H�u���9}>6��<�`�>�=	�>0�>��7?7�K?�TM?\�>v�;�l�>f��>�>&��o�s(̾�]���s��Æ?X��?�r�>Z�V����C�c���6?a�.?)��>�u�>Z�y�޿6����:� ���ۏ=3�X=�������Օ׼/�V���d��<4�>�>��>biX>vb�=��[<���>*��=��l>P,���6� ��<`Ґ�E>3ؽj>|�
�9�<]%���<
�<��]>�L�;)^j=�WF>���=���>>9[�>���=����o.>.0��gL����=�D���B��d�x~�3�.���6�D>�[X>���v摿?[>�}>>�F�?t?�!>��
���ؾ�ҝ�L�`�$�O�iw�=KA>��?�}�;���_��N���Ѿr��>ގ>R�>�l>�	,�� ?���w=	�a5��>�z��̮��&��7q�T?������si���׺�D?�E�����=� ~??�I?��?���>�����ؾ�30>I��W�=B��4q��k��+�?3'?W��>	���D�6s�PD�+!?t�v�{Z�K7���	D�dO
=	� ��Y?��ȾIѾ�D��ㅿO��%�/�ȃ��^�>fP?ƺ?-4w�3ϕ���>�o`#��Ax���D?��x?jSF><�"?�Ӵ>��P��[�׽��>��n?�:�?�I�?��;u��=��½F��>�P�>E֖?n��?E�n?��4�:#�>�Ab<�>�Խ��=.�>��=Y��=�k?:V?�?�ϲ��	���� ^���P���]=�g*=J͑>�ȅ>��>��>ru=���=^F>3O�>k�z>�kG>�a�>��u>����&��&?���=�!�>�+1?FI�>�]=�H�����<wf^�8�E�p,��ҳ�67۽m��<������T=�l��R�>ƄƿD�?�TO>�C�)�?�=��9�*��4R>B"[>��˽���>E4C>I�w>$-�>�F�>Η>��>�!>�FӾ9>����d!��,C���R���Ѿ�}z>霜��&�����w���BI��n���g�tj�+.��<=��ͽ<"H�?����k��)������?�[�>�6?nڌ�k
����>���>�Ǎ>�J��N���Iȍ�hᾒ�?#��?1/I>�ʹ>��5?)��>��<�<��V�k�=-^� �?��W��I��3���?]������(>gZT?�Y?5oS?��ݽ�K>+�X?0���A��k�>O5��ZL��T�=ƙ[>~#��D�JP��������?�[>Ё�?�w�?np�>PJ��+��,�8>}�7?*?�Zp?�5?�l.?���;T)?���=7�?�9?Y�-?Cy!?�'?c��=Zjv=�Ѽ*�S<���e:��+�Ƚ��߽:���`�H=�t�<G�(����9��i=3�=w�X�| ��#m7﫞�^�o<�Y;=z �=e�=��>�t?|9�>N���,�?ۉ���G���MU���N? �<n��*ΰ�,޾Z�9����>�?/e�?��9?u⑾�ܽJ��!�>�@>�#��N�=>�>$�f=$�3>�>s�P>s��=��=�S���� �ؾ������= �j>�,�>�t�=J���Δ�:��G�������>%(���L�����&|��<N�t׾<a�/?�xX?�?g��<_~��l(>h�W�G?}]=?��>���?WE�=�b����������<޽!g�>����.VY�Z����2���_-���C>���>�sO�rܠ��Xb>���\t޾u�n��J�����FM=R��`V=g�K�վy5�L��=�!
>4���� ����֪�0J?��j=Rw���_U��n����>���>��>��:���v�;�@����Q.�=յ�>-;>LM��i��JG�d9��'�>=GE?x�_?�a�?xO��;�r�isB��-���U��9Ҽ,�?��>��?��@>	'�=���F�ȉd��F�*��>Y��>N��9pG�����?��#$���>��?�>ƈ?a:R?�_
?�&`?h�)? �?4ޑ>(S��O���O$?��?\Z�=7ս���Y�:��G�D�>�@?��}��j�>'l?j�?��?U�T?�W?�O6>*���]H���>Ӂ>�[S�����C�j>�G?��>�bR?.��?ZZ>��6�Ǖ��ỏ��c�=,Q/>��5?.&?�%?��>�y�>�⠾��=���>�b?^�?�0o?ܢ�=R�?�>4>���>��=�D�>X�>��?��N?�Ms?^�J?�S�>��<􆮽�}��)an���Q�Lo�; �/<�qz=�!���w�,��	��<�ܳ;�>����_����E�������<3�>W[>����>��r����r^�><4'�J�Ͼ����9�=�A�>��)?Y�>�����!;���>N.�>i��x�I?V�>V�?��>��A�o�Ps&��g�>/W-?^��=��t��Z��8�x����c8_?�l?�ֺ�����,�b?��5?��T�R���m�)K\=���?p8?# ?�Q1����>�t�?\�`?Y��>m�Ӿg�y����pƁ�'�v>��T�.0�>����5��>0�?���>����5�;z�=�|[�X��{�>0�?_=�??�~?�2�>�政��=�����=a?�b�>R��(s�>`�#� E��m���#M���+Ѿ���B�о+|��I.��r_���p�,�T���>�!?��?}��?�Y?���'pu��a��҇���W�n���x��+�B�=l�Ͽm��;z����]'��ˡ3���,�F�}�P�@����?�'?D/��@�> \��ъ�nqξ�kC>c����k�J͙=�ݍ��5=��Y=��d���-��c���	 ?ݘ�><y�>�<?�w[�$�>�?�0���6�Va���2>��>�ƒ>��>|�.;T.����V�ǾN=��̦׽�1v>�}c?�~K?�n?���1�q��ˎ!���/�.�����B>�V>w��>��W�;���"&��:>���r�v���v���	�?~=c|2?�]�>Q��> @�?�?�~	�����w��d1�ٚ�<H �>�i?�,�>6 �>��Ͻ+� �ʚ�>@bl?ǹ�>��>����&� ��1{�Ɂƽ�>�c�>�G�>n�o>g,�A�[�a������k8�8b�=��h?cӄ���a�k�>A�P?i�d:J	t<���>'nd�ҿ �����#�!�	>��?&A�=M�:>�žPa���{�_Ċ�)�(? 	?�4��G�*��Z�>��!?��>5{�>Ժ�?T�>Z(¾g�5�R?fn]?�?I?�(@?״�>�*=����TOȽ�
'��2=-��>S�Y>C8p=���=��B�[���ީI=�,�=�^Լs���	��;1ῼlCK<�T�<��4>fsۿe1K��ؾ���	�Z
��ꉾ�Ա��Ç�j�	��㴾oř��y��u�6�(���T�Y�b�!+��@bj��A�?S�?��l@��
T��Z���M��"�>��s�F�w��Ĭ�y����eD㾾��7� ��2O�T5h�i�e�Q�'?�����ǿ򰡿�:ܾ5! ?�A ?9�y?��8�"���8�,� >�C�<-����뾭����ο?�����^?���>��/��r��>᥂>�X>�Hq>����螾E1�<��?6�-?��>��r�/�ɿa���C¤<���?/�@�0D?�x2�[����=p��>��
?�(B>�4������˳�>��?�;�?
B>��O�(G��VZ?w=�rL��qü��>|�=ڄ=�B�ԾE>��>A���2e<�4�!��>x�>�Hn��f��H`��	�/,^>oo�����-Մ?y{\�$f��/��T��^U>f�T?�(�>74�=�,?�6H�m}Ͽ2�\��*a?@1�?/��?��(?ܿ��ך>w�ܾ�M?D6?���>�c&�9�t���=%�Hf�����B&V�a��=ϭ�>ʋ>��,�|���O�gY����=>��B�¿�]����Ҙ~<� $�A�Ͻ���2���.��^>��m
Y��R�t�=3�=rsM>�'v>|OH>x>�AX?�Pz?���>>�>'ƽyy��'�Ѿ���_撾���퟾�34���־�
������X�պ�|O̾q =�<�=�6R�9���J� �<�b���F���.?0v$>Y�ʾJ�M���-<wpʾ.���Hۄ�jߥ�-̾��1�"n�͟?�A?������V����W�����f�W?O�����鬾��=���]�=G%�>l��=j��!3�r~S�� &?K�?آ��o����t>��hr*�f�%?���>�j�=���>�Y?��\�� >6��='@�>Me�>U�F>���O��hd?ŧJ?�����;����E>5%�����}�!�=$2�ATm��,>Rkpk�J1��[!�E5.=�V?Bj>U�,��/B������߽�.�;�P�?�'�>��O>�
�?��?�ԝ=,��J�����D��xo�qD? �?fY=>� ��J��P���}?/�?�tR�U��� ����U�g�(�Z�K?EZo?lZ?&��=fc�	L��W�-��(t?!�v?�p^�fr�������V�9�>�Y�>���>C�9�Ik�>��>?�#��G������rX4�LÞ?}�@��?E�;<� ����=�;?`�>��O��<ƾDq��<����vq=�$�>����Jev����O,�G�8?���?ԓ�>h���������=Cؕ�{Z�?��?�����Bg<����l��m���{�<(ʫ=�PD"�_���7��ƾ�
�w����Ŀ�\��>Z@XP轎,�>fB8�=6�hSϿK��
]о�Wq���?��>��Ƚ-���k�j��Nu�C�G���H����̍w>�o�=b�s������$�B���>[��>x���?Ȼ�h�辪(�8�	��=IN?�?k��=�s��A��?!|2�e����7��P8��r�?�ҷ?�}	?R�?�g]��E���%��0��Z?�A�?�)�?̉�<8׋��J8���j?2+���d`�6�4���D���U>|�2?G2�>A-�K�}=��>�"�>6�>Z/��ĿGѶ��G��ǯ�?���?H�꾔��>�`�?�:+?:�{��������*��{����A?�`1>0�����!��<�Eڒ�Z�
?b�0?�X�b��9!e?_�����T`�H3=n��>I�D6����u����=��C�����q���U�?�U@sR�?��7�2�>�s��>���>����V�d�ӈU>��>ua>�K�=.~��i �>3����*��CG=�4@j�@G�>~��uh���:'>�A�?)j�>gP?��^��><?A9=^	=lD>i`�w`�>����n�>QWF?^�l>?Y�=5���}3�ۀA�	u��(n)�quX�K�>7�+?�X?Cx���޽m=B}���T5����������[�,Q:�pQ5���X>��>�= �=�ه���?Fp�5�ؿ�i���o'��54?��>�?����t�^���;_?Zz�>�6��+���%���B�V��?�G�?7�?��׾0S̼>J�>�I�>m�ԽL���H�����7>�B?f��D��d�o�~�>���?�@�ծ?bi�H�?���8��vq~�:���D7����=U�7?����{>���>���=�v������s��>4N�?�j�?B��>�!m?�o��xC���0=�7�>�l?�?�ɮ�q��9B>��?M���莿^��?f?j�
@3_@rU^?rҢ�
a߿-���)��uEʾ9�=���=�Jx>ʊϽ��>=��?=�S<Е��5��=7��>�Bp>�&~>B4>�9>X
>���#�س������=|E��S�Ms��"�$����u�ܡ��P������䵽������ɽ��O���	�܁J����=JW?#�O?��p?<��>��5�[�>j����5=�R4��U�=�+�>�1?�PH?H )?��u=�����d�K������邾���>�5>L��>A�>�Q�>5I<�A>��3>|~>��
>��J=ȣ����)=��G>S��>M�>-��>�C<>��>Fϴ��1��k�h��
w�q̽1�?����R�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��|�T�4:>:����j�5`>�+ �~l���)��%Q>wl?�f>�u>j�3�V_8�y�P��s���n|>�06?�޶�g@9�W�u�p�H��bݾ�FM>쿾>��D�/l�������/}i��{=�w:?��?�c���䰾{�u��I��'JR>J'\>�=/V�=GPM>�c�0�ƽ+H��S.=���=w�^>%?lT;>�ז=���>�pz�vC�Ȩ�>E�L>��'>��;?:�?��(�$����}4��l`>K�>�'�>�+>J�K�n��=��>3b>`��zX��N��C� ��E>������T�8K���"=�ѽ�ʅ�=$"�=َ潬C9�G�=��~?�ֵ��B��E������=}�7?"߮>��;z>����M��	[���5�?e�@9k?'���3H�[�?�h?�Lڽ���=�߳>��*>�G��6���;�>�@�>Kٻ���E�\�>��?���?�E�"c��)����>#�R?��{z�>�h��W��4����u�
�#=a��>MNH?�7���lP��=�ݖ
?�?�]�����ȿI�v����>��?��?��m�o<��G @���>1��?DY?�/i>w۾h�Z��W�>o�@?9R?�#�>��?�'�q�?ƶ?ǵ�?�I>���?V�s?t�>�x��U/��1�����~=�[;�^�>4@>���0eF��ԓ�4d��}�j���S�a>�v$=��>�>佽/���_�=�勽�@���f���>Qq>=�I>�U�>z� ?~_�>!��>[I=3,���؀�RÖ�}�K?�s�?"�8"n�ץ�<c}�=;|^�D?NI4?�����ξj��>eW\?ģ�?��Y?!�>�������5����Ĵ�a|�<6RL>�q�>k��>ǉ�anL>��ӾG�C��t�>x\�>��`�ھDt��!]#�<�>:{!?�+�>�Ũ=��!?	�?R(l>�6�>�]��M���~2����>ʃ�>r�?���?�?R⿾�6�Bf��J���*H��W�>El?U�?��>����1���h�<G�<+����u?�c?0��#?5H�?[iJ?�w5?��D> o��b�@����e�>��!?�W�O~A��=&��~��A?/"?غ�>R���p�ֽ1Iռ"���f��l�?��[?�#&?�]���`��Zþ���<%r(�d"Z� �;��=�ֽ>�>}���3�=��>��=&m�k6��)d<�Ž=���>S��=�7�^x��_� ?6�=��ӽ�>̓x�ǡS�|�> �a>@Ǻ��$k?����ң��ծ���)��PՇ����?���?HX�?/?0<�}U�O�?�|�?o�8?N�>n:��l���&�ʾ����4�Qy���&= ��>�@�=�+��ʝ��*��K`��Žf<c�ѽ��?�=?�?g�>`��=�~y>%+��5�)ͧ��g򾡵W�4��m>3��`,�>��h\/�*1�X�=\���)c]��>��S	�>��?�>{z�>v��>*���f_?Epq>�9>�0�>;�:>�=��Z>�5�[4D��xS?X{���2�̐l����I ?��?�1Z>��g�~�%�8�z�??�ߧ?�9�?X�U>�e�.�2���?J�>Mž��E?��F>�3����|��h�h�=n�n���þ���>��-��@�;�B����?}\A?�.�sd۾Yk-���ľ��K=z��?}� ?��(��Y�MӀ��X��
T����n�e�k���6�rYx����ʉ|�xx�z�
�@=B�2?'�?i�Ǿ�ܾW箾]�z��_A��{A>I`�>�f�>�M�>�1;>�����F�2Ie��)�R�9����>��e?��>~I?h�;?��O?A�L?!�>�:�>v���05�>CY&:Y��>Ԩ�>a8?�-?��/?}?(q+?Mof>��W�����׾��?�:?�V?G� ?�"?�؃���½�����C���w�l���1�|=�K�<�Mн4�e�@>=�xN>I:?g���93�mB�=(�>��9?Dc�>N��>{�w���d���J=���>��?���>����@cp�µ����>�!�?�J�R��<��3>��=۽c��g�;'@�=�]'�1�7=v��i7���^����=���=�3N��tк�mZ�"�^<��=���>?(?.��>&<�>�پP40��׾餥>|^=B/�>��>(���p���e��_y���Q>�e�?)�?�3�<�Fs>2yN��n�TCľ	2��z辀;�=!�?�a3?:�L?}��?s�\? ?��=���;���l��tf����?c!,?���>m����ʾX��3��?�Z?{;a�8��;)�r�¾��Խ0�>�[/�D/~�����D�4������~����?�?M,A�Z�6�kw����\��ܓC?@ �>X�>o�>:�)�y�g��$��0;>Ȋ�>�R?�U�>
�O?��z?^D[?��X>��8��u���>����w�JW>\�>?�Ȁ?���?�x?r4�>V�>p�%�s�ܾ���A��ʳ�p肾��N=Ԅ\>��>�W�>���>���=��ҽF7��X>����=x�a>��>���>���>�-q>�no<�A?#n�>�E���r������%��2�����k?���?,?'��~���F��i��0�>ۨ?�Q�?c*-?b�V��u�=[�����0�B�s�>�p�>�~�>aݣ=��<G�R>;l�>(i�>B@��H��/�}�ּՊ?��D?���=D<ƿ��q�{�p�����R�6<���/�f�1Ύ��PY�JΤ=
Q���� R��)fZ��.�����j���|����z�J��>&��=��=S��=���<jkԼ�ɵ<�
J=�<b,=�vp�x"y<��9��"ջ�2���k��x&e<z�@=>A���z���;�?`C ?^?�=?��;?�>�5�=]6!?`����yD?�^�>��F> 5��>���%���Ӿ���
��/�˾8Y>B4R�:�f=��1>Ǌ�<���=R`f="�>��>tB��Z�==Jw�=�� >��=M�=Q�g>���=s�k?�?��I��kM�S���D?���>���x`�2`?g5j<�.���@���/��Ȇ?��@�U�?�l�>"�]���?�#�����ၒ>n��>��,>P�߽�p^���>�>��H�ˀ���j=�.�?kA@��G?�����g׿W��=^k<>J$>�M�0�.�D�?��<o�YY��?1�:��/վ&Ђ>��=�a�/ľ΀X=��?>�;�=O��^�ҡ�=)⇽y�$=��6=狌>ScB>R�=�����m�=
r8=�n�=��P>U���*s]�هܼ�%`=�k�=SK>��">�n�>��?,�?�@?��?3���`�̾%ū�~i*>ϙX�od>h�����=u��>��5?�D?̽J?xr�>���V1�>�Ǚ>Ǽ���a�򮬾�=����彋K�?*��?W��>��.=8�S���LU�9n��Ot?	0?���>E�>���Kӿ���X0�؂����<�Ž%��=��<rf��tl =L�u�=��>&�?�}W>��=	1>���=�.�>�^>��n=C-�=ϭ��r���>L6��`�=�ԼEq@���}���9�o��q#F��kA���v�VQ<|0�( �=� >�/�>�'�>L��>K�[�־� >x�c��/b�I�I>˾��T��`��kr���4��½�}>P�?>��=ڛ���T�>!�>��!>U��?|j?�Z�=�숽����V������&��A�=Vp>:g2�OHP�qT���G��oȾ��>��>G�>>fl>�+�?���v=}��]G5�!�>�b��P����&q��;����i�jQ ��D?b@��H��=]~?Q�I?�׏?m�>�И�Z�ؾ��/>z��2=%��Aq�Y�����?@'?L��>0��D�wE���@�RX<?����N��$���U�r�u=�S"�l.?2���u���_�?C��m���x� �V=8G�>�u?�ɻ?�Qx�ʘl��;���5�׊����2?�Bn?�Z='�$?{��><��@�þ�n����!=�@Y?x�?+��?Px!=?��=���/&�>�?l�?5�?�p?v�;����>��<��> ޕ�qd�=�h>~ȗ=�l�=�
?�	?�?�ߥ�+	���쾯5��k�\��=P�=�)�>z3�>T�v>��=q�= ��=Y\K>}�>�̊>�#d>oԞ>K�>_��������&?k��="�>u�1?ׁ>��_=ǧ�c��<�MD��=>���*��X��d^��1�<ʩp�GS=Shü�T�>�Hǿ�ܖ?��Q>�j�?.����&�7mS>�.U>�"ٽ���>�E>|>o��>C!�>��>��>�'>/DӾ(�>���3[!�t,C�R��Ѿ[mz>Ғ��0&�����d��<>I�po��~g��
j�
.���?=����<AD�?����Q�k�u�)�����;�?RX�>n6?[׌�_&��α>���>cɍ>�I��c����Ǎ��e���?h��?�8�>���>S?`=?��;�q�P��lS��;��r`��P�%݀� d���󈩽guM?>�d?�P?!珽j�R>K�l?�:	�X""�xأ>JE>�N��1��+� >0>��^,�^���������㧏>-�r?.b{?��>UZ�ޞ�L&V>F6?vg?	Hb?��9?�*?#J��{*?$�> ?vE	?$�/??�?�?�$�=2~�=�H <��_=����2k���̪�R
�[�C��Gb=ȳ5=�K�����C�<���� �<x��<hH��a ����<�8�=��>�\>)Z�>�Q?k �>v�F�?N?�����T��: �d:?�X ��ھ����g�ھ�E�{N>Ң�?j��?/�N?~�3�
�V��'I�DL�=���=�7���(=np�>�L�Ӽ�2�>F@�=1�L��§�	��	��&���#�Ľ�^=�'}>���>	~>[9���,>>tl��{�?�w>�5���?ž�^N�s`Q�&�0��05�:��>�jG?H�?��=S���b"���_���2?s�-?<9?�q?�a�={	� �"�"�B�׽�>����d������!��y0��q�=n�{>��c���ƾ��H>0���Ѿ_h�9-U��+�\G�<Å	����=�_rǾl�d���>��#>��ʾw���f���<���4M?)ʄ=0����`�����=w�>-L�>�a�+�;�^�5��ா�(.=9v�>��>�^�����C����L�>͞>?z�d?Z��?�w��j9n��0>�q=��٣�Jiy=3`!?Bm�>��?#;>o�	;+Ӿ{R�v�Z��<��y�>QD�>���3;J�غ�����8��[�>bD?V��="X?e`L?�?nBT?W�"?R��>���>�@�����<=&?K��?���=�׽ڄR���8��!F�r��>�*?��E���>�R?1m?6�&?z�P?f?��	>I�}RA��>��>��W�x믿)�`>B�J?�ĳ>��W?��?�F>>3X6�A�� ����V�=� >�3?"�#?�y?��>`�>�ҡ�^m�=�^�>2c?c/�?��o?	��=��?T2>?�>OL�=J)�>�E�>� ?9+O?��s?�J?�U�>R׏<�������%nt�h�Y��0l;�(G<��x=,b��w�A��c�<���;�����~�m^��b0C��팼6��;9�>!�s>�蕾��0>��ľ������@>f���o���D�����;��`�=�A�>w�?I��>�2#�ڂ�=2��>�v�>���Y�(?D�?�?v�;0db�"�۾�xK�z��>�A?P��=G?m��f��,�u�4�d=��m?+v^?E�U������RZ?�c?�ީ��.��(���ɮ�'��:�y?�"?v���d��>�E�?a�[?���>Ӣ��c�X�������]�5Ӿlp=	��> �-��.e�K �>��A?�G�>��&>���>$��m���0�*f�>�ԉ?��?�R�?t�|>|�(ڿr���؈�1�K?K��>����z$?3�<ThѾ������I���窲�>Z���舾=؋�+'�hҀ��߽��=��?()�?lk?ϭS?.���V�Ae�4nn�v�P���b���vX�g�0�H�1��E]����ʾ^
5����=�<��j.A��^�?&�'?�"/���>Ko��v�.K;�bD>R�������{�=k���==t&T=��h��/��=��� ?��>��>}<?u�[��Y>��1��57��a����2>��>J�>���>֪�:��-���뽀;ɾb�����ӽ�~s>2�c?�0K?�p?][ ��?0��5��ٔ"���>����@>�>W��>�[� ���l&�hF=�b5q������	����=R�2?�X�>T؛>�ۘ?Ƿ?#�JS��~,r��/��u�<'��>�Ah?��>�F>V~ֽ�9 �S�>��o?X��>��>}�u����[�f��)��Ԭ>]��>B]�>kTs>i�>�Q\��l�����e.��
>��N?vU����c�U�j>�`?�� ��2���>@��G`3������yF>��?���=n�r>�&��e*��5w�e���SA)?[?ӣ���d*��E~>A�!?���>j�>�S�?�K�>�RþPCx:õ?��^?��I?�BA?�M�>�=�j��3�Ƚ��&���.=��>l6Z>��m=���=F|��*\��U�H=U��=�"ɼ,s��N�<Mb��C&Z<��<�N4>.��@�G�O��@��֨�X��H~���"�P��8����zs��n��f�5�cnϽ�|�<��I�FF��&��������?�,�?�9�M\�����i�����]_�>&^v�
s������ ����˾�I����(��DF��v�L�p�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >[C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾u1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�|A?��(����eV=%��>��	?H�?>=S1��G������S�>�<�?���?�M=?�W���	��e?�@<i�F��ݻr�=I>�=RS=���7�J>�U�>~�� SA�8ܽ��4>Eڅ>�t"�w��r�^����<�]>��ս�7��bՄ?�|\��f���/��Y��Td>��T?!�>�>�=��,?$;H�.zϿD�\�*/a?0�?o��?3�(?dӿ��ߚ>�ܾ	�M?�A6?� �>E\&���t� T�=�S⼋N�����<$V�:��=f��>-a>]�,�=��O�k������=έ�	���uM�֦���<I�H�J�޽��I�<����B���);�swO��W��aͬ=+�+>��Y>��>o�,>"�;>��W?��v?!8�>x�5>�N��#Ͼ�O�๎��G��Jؽ��[�SC#��m��H�۾��¾w���j%�f��"=��=?5R������� ���b���F�#�.?�u$>�ʾp�M� �-<�nʾ���������㥽�,̾�1��"n�O͟?y�A?�����V����Es�K���ܮW?uP����鬾��=���r�=w#�>	�=6��W!3��~S�'0?W�?ƙ���q���V,>D�=�<��*?�?vn�<�˨>d'?��%��ݽ�V>�6>�>'0�>��=s���9ܽ*�?*tU?�h�f͚�B�>/ ���x�ju�=[�>,2�@����SX>�q�<������޼��`��<�(W?u��>��)��ya��|��Y==��x?��?$.�>m{k?��B?Oդ<(h���S����aw=�W?3*i?��>����	оX���C�5?�e?��N>�bh���=�.�\U��$? �n?4_?4~��*w}����p���n6?��v?@s^�{s������V�M=�>R\�>���>m�9��k�>�>?:#��G������"Y4�Þ?��@���?��;<)�ݘ�=�:?�[�>V�O��<ƾ�w�������q=�"�>�����ev����!P,��8?
��?<��>>���
��4��=*ו�AZ�?��?@���1Cg<���l��o���Ġ<�ԫ=���D"����}�7���ƾb�
�W���0̿�8��>Y@M��'�>:L8�\5�PTϿ����VоVq���?�~�>֡Ƚ����}�j��Nu��G�7�H�Ƥ��kM�>��>¸�����y�{��r;�����{�>��
�>�S�� �������4<u�>S��>���>����ܽ��ƙ?Fj��WBοu�����k�X?�h�?�m�?p?~-9<t�v�)�{�0"��+G?�s?5!Z?�%%�'']��8�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.���r?K��󖅿7K����"!�>%j�g>���³=��6���Z��!��T2���?+�@��?�)�:J
�B�"?�E�>�O��_H��H}�<��F>+��>ڿS>tۆ9�hN>B�@��Q�O��;���?̔�?7Y?r���;��c��=~_�?�8�>+�?���=�&�>�|�=���F�H��U#>m��=e�=�?�>N?m;�>K��=
�9�.p.���E���R����m{C�4e�>��a?��L?Ҳ`>�T���g-�e!�F�˽(�-���ڼ�4?��M$�η߽�'5>ْ=>3>�^C�%�Ѿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji���
?k� �s�~� ����*��y�.z?>؀c?�H���3z>���>�/>1���Q�����R��;�>)J�?��?� ?<%�?�������=����>���?�f.?������о�j>�X�>^��GI��o���ف?,t@�h @�^Y?>A����ӿ���8�������A >���=+�H>� �N3�=�=�HH=yH<��0>ٗ>zp>DEx>�[>*�O>��9>�����#������>��\�>��,�\�
��4s���Њ��%��w��˟������k���:Ze�5�L��#�A��>��V?MDF?��h?���>�r���ȅ=7��1=�>a�&�AN�=��>��8?�s??�w?��=@�H�1�j�$����^�����W`�>c�>�Y�>}�>s��>6s��WF'>�ڐ>�f�>I�>��>�V��9��=.L.>�Z�>�d?7"�>�C<>��>Eϴ��1��j�h��
w�t̽1�?~���S�J��1���9��Ӧ���h�=Gb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>��q�T�/:>8����j�6`>�+ �{l���)��%Q>vl?��f>g�t>��3�O8���P��(����|>�6?�����'9�I�u�3�H�Xmݾ\M>ֽ�>�D��c�$��~��7i���{=�:?vo?�ճ��ⰾ��u��B����Q>!�[>x�=��=#:M>�b�Сƽ�H��*/=�F�=W�^>�5?c�+>4>�=��>���O��y�>2�A>�,,>�@?]�$?Y��T����o��S�-�o�v>��>Ұ�>�>]J���=~��>��a>�	��0��w����?�1�V>�?� _�}dv���y=�O��=�E�=	# �H'<��}'=�V�?֭�����!���վ9�]?S�I?F�o>B�=n[������-ؾfc�?�@��?]1ʾL+G�)�$?X��?�,��jm>�Z�>��>K�)�懾`??S��۾��׾.���.�?�G�?�b�s|� xI�;g2>�?񉞾Jh�>�x��Z�������u��#=N��>�8H?�V����O�Z>��v
?�?�^�ߩ����ȿ0|v����>X�?���?h�m��A���@����>;��?�gY?�oi>�g۾A`Z����>ѻ@?�R?�>�9�f�'���? ߶?կ�?;>�o�?�(u?�H�>H)��)�����G���}�<�n=�l�>�*>����F����)+��Am�f����j>q+@=�̧> �Žv^���=����������*�>�|>�n>P��>��>P?�>�e�>ӌ<����az��Ԓ���B?��?o{����T���=���<z���
�?kf?-����۾�R?˂C?�Vs?C�-?��>'�sv����ǿ����=8v���/>��	?�7�>��<*�B>���jcK���>�Zq>���;����d��݂<���>G7?G4�>�'>��?�.!?�v�>^?�>o�J�w�����Y�i��>�&�>+0?Zj�?c&?`̓�m,4�!��u��"�j���:>l�W?'
?�`�>�9�����|3=0��y;���?��y?�h����>L͂?Ak/?�e;?Ĭ�>��M�l׾[{��V�>F�!?�n���A�b6&�&Q�Q�?�T?$��>�擽$�սWۼ��������?�\?�"&?���a���¾���<\�"���%���;�-M��[>�E>�눽Ȩ�=�%>�V�=Ćm�s86�o�i<�c�=D�>Dx�=$�6��.���;,?+0G�'׃�v��=��r�XvD�^�>FL>a����^?p=��{�x��Ix���U�\ �?���?�j�?����h�`#=?��?�?\�>�J���u޾F���Uw���x�-t��>���>��l�L�吤�8����F��a	ƽ�T9��g?$S5>r/$?y?�	�>��>@eؾ�N��7���ݾ�X�etӾX*�Ԛ"�� �{��M�u�c@��Hw˾WĖ�侵>�2���>�_�>�D<>>>-�>A�H=���>z��>ݾP>���>�e>��=�l�=T;ɼ�#5�&�T?�̾<,���$޾��B?-n?g�>0(=�>��Lr�DG?G��?r-�?��>��]���&��V?F�?=(����?�`=��<c�a<��(#�������ZV�>%Z���6�[QU��󊾳��>�8?4�ӻۙо�@ؽ�i��&��=Ȏ�?w�4?�W��AO�/�X���Y��M����=-ѽ�#g����@+j�5�������~��=�$���Q=Q(?�>o?���e����0!k�I�M�q0�>���>j=�>	��>7�X>[���+�I�S��"�	�e����>¡o?�(�>�UJ?�;?_S?GF?���>a^�>&K��DC?�� =���>zQ�>=E;?��)?%�)?HX?�,?��O>���Y����9־��?/,?�??N�>��?�;���?ؽ7!�j�r<�Mm��j)��Ry=@'=*d���b���=&@O>�&?)�V�8�^�����k>w�7?���>g��>36���쀾���<��>�e
?��>ϓ���@r��W����>��?+����=��*>��=3h��"����=�"ļɨ�=I����b?�'�<$�=hm�=ڊn��G%�P6;�G�;�׵<֍�>#!?�܏>��>��|�p���{��B�=��U>�W>��
>��־3Ɋ���2�h����>�ߐ?��?0��=�I�=�C�=^%��qN�����ڊ���[=���>�?.%L?�^�?��B?�&?�I�=ȟ��̔�{���K ��?u!,?��>�����ʾ��͉3�ޝ?a[?�<a����;)��¾��Խױ>�[/�a/~����;D��녻���(��1��?쿝?�A�S�6��x�ؿ���[��w�C?"�>Y�>��>W�)�~�g�p%��1;>��>cR?G+�>a�O?��z?�[?��R>��7�򠭿;R��I�0�CZ'>��??&T�?���?Mx?���>�>��#���ྒ:����#�5�� ���l&g=T3V>'�>�k�>D�>3�=0������=�Lk�=��`>�`�>��>���>��z>�V�<��G?���>�?������ɤ�����>�͓u?Q��?4|+?�=���1 F�\@���%�>gn�?O��?�B*?$�S�ժ�=F�׼/Ŷ�!�q��4�>���>�+�>)��=)G=��>���>���>0<��Z�ru8��`L�m?�F?T��=r����b�������&�=����F]�P`��g�,>1]�4f�ew��=� ��$R�͜��d8���۾�派S)?*�=�X>��'=��7�^i���|=3��=��˅�4廽ߑ'��r��٪���[����>�;ڙ=��.=n�þ��r?��D?��I?�%:?=tt>p\>Z��#�=��<�2?F�[><�<o�ξ�����þ?Ⱦ#PɾVS��J�`��ƾ�vS>�{��I�">+>��=�4�;�{�=K>��1>*�=q5=|��=ۑ���Z�<�7���=4�J>�6�?Ռ���ӥ��Ji��n�8�B?���>vx1>�f��]�F?-��>��o��۶�����?���?Q��?�?V��9��>w���ID�(�e=f=Y<���>���=��u�
�>? >�(��n��!��=�h�?��@u=?]甿�̿|9>�F7>��>ҭR�Q\1�|e[��ga���Y��`!?�C;�g�˾繅>"��=�8߾Qyƾ�V/=Cm6>v0`=���G(\�h�=��|��@=�j=�t�>]tC>'-�=	H���X�=��F=���=ȇO>�D����6�+�NN2=C��=B�b>�y&>ݎ�>��?`0?HUd?�3�>p�m�W!ϾY<��@�>`��=7:�>���=)`B>��>I�7?d�D?�K?���>Mԉ=��>��>��,��m��f��ͧ�@�<#��?s̆?MѸ>��Q<�A�
���d>�HHŽ�w?iU1?�m?Z�>#V����DM&��.��Q��P�08J�*=�r��jU���:4�3��HE�=�m�>��>Q�>�Oy>H�9>��N>H)�>��>���<F��=�M�����<����O��=�䒼�6�<�Cż�Ӕ�M�-�i�+�4��u�;��;MaZ< ��;�
�=���>���=-�>�=�=�֚�p&>>�ئ�ώT�N�=����0K�62Z��<v��+��	#���>-9>:��̷����?ӂK>�q>څ�?�l?�9�=g����ݘ����gdU�|��=o��=�e���8���`�0cL�Qܾ��>�ߎ>��>ʾl>|,��!?���w=g�/c5�J�>�|�����'�59q��?��`����i�;gӺ��D?RF��]��=W!~?�I?&�?���>B��ؾp70>vH��a�=i�>(q��k��9�?�'?V��>��w�D����������>�p���4��ܡ��u+�#3�=<��w��>V27��)��B	5�[툿�����bb��@5��j�>J
l?���?� ��|���'�Y�����n�=H9?߀?D&�>h��>��>����S���	��j~{=��|?L;�?���?o>���=�崽{0�>�?���?"��?��r?S�?�_(�>�{�;��>�m��O��=t�	>m�=��=\*?�b	?��	?����
�F^�{��^�jw�<���=|n�>PV�>ʕr>�-�=]Iq=Rڛ= +\>aB�>��>��e>
�>͉>�[��ƍ�>�?ϣ�=63�>bV<?�z�>�=�� �Zrx=���(2Z�3'>����%�����&=.�n��B�ʋ����>^�ſI��?_/�=�S���
?yN˾�+�͇>��\>+�H��?�>���=��}>u��>���>��:>�6�>nI>�e�!%�=N�ʾ���A�1��p�&�Ͼ�O@>����Rj�������ܽ��A�*����?)��,iq�A�M���ؼ�@�?���JY�[])�W�����>��>��;?���S�H��� >0��>��6>"��g���h���˾$��?h��?��C>�'�>�x:?G*?M�	��t��լ\���E�*�D�&=��#�f��|���y�(ﾆճ�=�A?��e?�eS?8�$>�+(>�|?��о>��;�>��"��G��k>U'�>l�x�s�H�����羅5��B�Zzi?]W�?p�.?c����k�tY'>�]:?Չ1?��s?W�1?�;?@a�\%?�5>�?n�?z5?�l.?@u
?/�1>ˋ�=u׻��=x������d̽�Ƚ���U�1=p�}=żw�h��;�n=�^�<�����Լ��.;����{Τ<*;?=>��=���=�G�>`if?\6?J�R>�QC?���1�L�e~��i�>�� >���aH;�v���3����?E�?v?��>�]H��yR���>tI�>g��=Pa>j��>+'L��ڎ�=�A>?�i>�=�>K�>_���d��~����� ݽ ��=B ?{�>���=���n1ؽ�8�>H��x7ݾ1�X�o�a���>�h���y�> �D?HN?�!8<��þ�=3�w��IT?�?2Ae?�]�?~�<���=8��l��]m&�@��>�J��+�(�;���7᱿%�%������=����������>�����վ��g��>�\���t���(��<T=�߾Xľ��7��5�=�=��ھ$�-�L��kݱ���R?�e>�y��i���v���p<Y��>B�>�OE�Պ��};8������=���>>�>o6�3��G�S�����E�>~�O?>z?f�u?�_��@�o���T���Ͼ�H��jd=�~;?H�>���>*�	>L5�� ��o,��]��w���>��>gx��A�P:�?�1����L��>bT�>�p3>�w?���?g��>d�f?jP?z�?R E>z�Ƚ��㾱�?նz?V=���<G�ֽ� O��F�]H!?;>?�ý�o�>�F?��?I?�3?T�?���=�����`K��o�>->e���#����F>�?UT�>��s?Kd�?�]C<�#�DAl��2)�S��=�=\9C?�b?��?D#?m��>����h�=ɇ�>�c?/)�?��o?���=;?�z2>���>��=�ß>���>� ?�RO?d�s?�J?�b�>+J�<!)��������u�C�T��'�;�-B<y=�S��iv�-}�?��<cG�;�S���+��|��0E���UI�;���>�u>qF���1>��ľ&����QA>�����ܜ�!x��I0@�H�=ǀ>�M?�Օ>u�#�.v�=S��>��>Nv��w)?X�?r�?�v;�Mb��E޾��K��;�>��@?g��=�m�h@��:Qv�O�O=�m?��^?� V�T���3�b?�]?9g�=��þf�b�#��\�O? �
?.�G���>��~? �q?I��>��e��9n�)���Cb���j�\Ѷ=�q�>�X�O�d�J?�>ܛ7?5O�>/�b>�'�=Wu۾��w�}p��?i�?%�?���?�+*>��n��3��þ�&t���P?2;�>�S�Y�/?ʾB=����Q��̴{�O	�/׵��k��:y�Y�b��.��𜾌٩�6">5�?ʣ�?�Xg?��W?�����\Z��b��S�h���U��>&��'�)U��6�m�9���g�����"��(�B�nf>4�v��?�aN�?�j%?�x$����>
@������;�rM>-3������=�R�i=�9V=�Os���.���T~?��>���>	9?0�Z���=��5�t8�����k>�Q�>TȒ>\2�>� <�(�[p���ž��z�� ���*v>yc?��K?J�n?�x�'�0��V���Z!�DW,�����,�B>|v>>3�>�Y����o&�U>�har����0��c�	��{}=1A2?��><��>(�?]�?]S	�\�����v� �0���<�>]�h?��>Jb�>N�ѽ�� �|�>�Lk?�$?��>�V��@���9k�t�\��>��>�-�>[�->��[�ig�ƍ�����r�2�l_>��(?D�p���:���S>�n.?k���f�=ݫ�>�S+��������df��:D>�?�Jm=W�>��¾s��Z�h�M���#(??����m'�cE�>�?���>��>�΅?�J�>�����<^�?\?�\E?ʨC?���>jU�<�������*h$���<�h>'wU>Ek~=���=�!� #O��6+�7:=D�=�����_����y� �p��o�;�=��C>nzؿ�BP�L�ɾ3#�d9�eR��%���|'F�����t�齫̀�/*��bW/��Q�O�e��f��Ƌ�)�������?P��?�AF�����9����8v�u���{�>�٨�(!{��H���ǽ����;o�*n��η5�GtQ�ߒy�t���N�'?�����ǿ򰡿�:ܾ2! ?�A ?5�y?��8�"���8�� >OC�<4-����뾮����οF�����^?���>��/��m��>᥂>�X>�Hq>����螾b1�<��?5�-?��>ˎr�1�ɿc����¤<���?0�@�|A?��(�L�쾉V=<��>��	?y�?>�R1��H�'���6T�>:<�?���?�M=��W���	��e?�t<��F�#�ݻ_�=�;�=�?=���<�J>aT�>���SA�0BܽX�4>)څ>�}"�~��ق^��~�<�]>��ս�7���Մ?�z\�	f���/��X��Ia>V�T?Q!�>3;�={�,?�=H�{Ͽ�\��/a?�/�?;��?��(?�ۿ�5ܚ>H�ܾ��M?�C6?;�>g^&���t�^\�=�1���c�㾍V����=��>B_>ȟ,����xO�:�����=Y� �hmÿ(����|��=��9;I��%J�8��2(��7e��.l����Z�=���=��y>=}F>�34>ĝ�>sZ?L�d?s�>�H^>o!;�X]������Ե��/񽼊�0�����A�޾�����@�$���!�Rd��%=��={+R������� �%�b���F��.?$>5�ʾF�M�w�-<lVʾ˾���)���6��B̾i�1�.n��͟?��A?	��V�N��<W��X��d�W?�_�f��7款ې�=���!=U�>c�=���7,3���S��f*?��(?�5���A�	�=F����?���-R?�_,?U:�.�>�`?VJ�$iǽW�W>�x�>q�>���>�z=����N���*? �S?{�K��Y7��S>���*�-�%]�=��>F����g>��/>��=�^�q��=!g��Sd;�'W?���>g�)���L_��A��O==��x?��?�+�>J{k?��B?��<�e����S��jw=9�W?�(i?�>�����	о����`�5?�e?%�N>ah����e�.�gT�6$?!�n?&^?9����t}�<��R���n6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�%Þ?��@���?j�;<��R��=�;?k\�>��O��>ƾ�z������3�q=�"�>���ev����R,�g�8?ݠ�?���>������j��=�����H�?y�?�=����p<Q��zl��x��V��<�0�=3z�)"���]�7�v�ƾʼ
�Ƈ���ƻ�ō�>`X@ω��N�>X8���-cϿ�����|о�"r�˕?ݩ>�ɽ~���:�j��5u��gG�רH����3�>��>���Ev���v{�g�;�e���;�>�\��>�LS�����j����;;!�>���>J��>��s�����?�e��<�οU���\I��Z?�ӟ?�H�?\(?-T<akr�	�y��j(�8G?1�t?��[?�T"�P0[���C�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.���t?��v�^���h�p%=���>{0=^�=�->nW�^Z�4����7��i�?��@uն?�lI�����D(?C�>U^l�C�x�Φ=�_>���>�m�>�A����>E�L���pH�=���?_�@?6~��<Ѵ����=�{?;��>v�?P��=�Z�>]W�=�ү�,0��� >�>�=�{5�Ƈ?�M?�P�>�J�=m,=���/�bUF�}pQ�"�\
C��>��a?U�L?K�e>�N��*9�� �ñԽ)�5�uڼ=><��&��ڽ�<5>@>ؓ>;�D���Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��?��KS��ٸ��0`��H��$�=�^c?<Xľ3<>��>q�=�
���:����P�V��> �?4�?���>D�?(�t�.�������rY>l)�?�>?���=�Q��TV>[)?��߾q�������)j�?Av@f� @c|b?In���%׿�|��#m��ȷ��_>@
>/(X>S���c�=Ё�<,�R=1�=]� >j�>;Y>n��>WKq>��>UP>�)��.%�˟����ǁ0��n��/:�N��� ��j���F�k\������G<��	�}�Ҽ� ������R�=CZ�=b�U?q`Q?��p?�� ?k���D >xt��UO=}�'�=�7�>�33?!�K?s�*?n[�=a�����c��=���<������w�>�$F><��>�c�>[ʮ>���;*ZI>�>>k~>_E�=�$=4���=��Q>�é>���>%�>�C<>��>Fϴ��1��j�h��
w�o̽1�?���S�J��1���9��Ӧ���h�=Hb.?|>���?пf����2H?&���z)���+���>}�0?�cW? �> ��x�T�4:>9����j�5`>�+ �}l���)��%Q>wl?_~f>JAw>��3��O7�;6O�z��
x�>m|5?�D���9��u�)BI�ӝܾ�L>��>1@�������f�}��^k�H��=�":?#+?E���|E��]u�x����V>fX\>�(=��=��M>kje�uʽ��F��,=���=��[>;	?3>���=l�>\�b[��أ>��T>��<>L=?��$?��x��
$~�\�%�L�}>���>&�>��=cH����=ZH�>
g>���,y��5�)H���V>\���8�a���L�ֲ�=ܼ��L��=ʔ=j�;63��N@={�?4w��c�����.�X����c?=P?�>�F>6�`�E7��V]Ⱦn/�?HH@�?8�徎�\��?Kv�?'Y ���f>8��>J�	?�Q6�*ގ��n?�մ�r!��i���/{��Wٚ?ߜ?@���ʊ�e�T�WQ>���>�w��Ph�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?eDK>�R�?A�|?\z�>�5�ܾ�u����c�X]!>��H>�"�>�)�=X��l`�מ�������k������q=᱑<���>��4��|ž�ԗ=���˙h������kz>��>�$�>v	�>)$�>]�>>�}>~�J����n��چ�/�K?i��?
���1n��U�<��=ز^��'?5J4?ƀ[���Ͼ�ר>b�\??[?Ge�>����=���翿4}�����<F�K>�1�>�G�>�"���DK>{�Ծy0D��n�>�Η>�??ھ�,���|���B�>�e!?���>�ۮ=�� ?֡#?�k>TG�>��E����b�E�
��>D��>7F?ش~?��?�ٹ��m3���_졿x�[���M>��x?e6?���>Cy��Ώ���N���H�UO���?[qg?���?7�?	p??�sA?�e>g��!ؾ�୽|��>�!?/��7�A��"&��,���?�c?v��>u����ս�ؼ����3����?��[?#7&?2���4a�Խ¾���<�p#��|M���;?a=��>�,>����!�=�>ܓ�=im��6�_Cg<qл=�u�>~��=��6�J;���<,?xG�*׃����=��r�wD���>{FL>��2�^?�m=�P�{����kx��U�g �?��?tk�?)��Q�h��#=?Z�?�	?�>GI���{޾|�ྵOw���x�u���>#��>��l���,������XF��~�ŽV�нH	?�E+>"?;�?���> ��>��R��J�s'ʾ�P��p�)��<0�Q`�����#޾i���HG6=a�̾�c����>�yؼ���>��>O@5>0ѫ>@4?Es> �>�m.>�ck>�Nr>���=D�$>oc�=ag=KW���S?\/ľ�_*��-�jžV�B?
k?�v�>�.]��邿k����?�N�?$�?�6�>��b���)�L%?S��>k���?(-a=ݶ=���<�q��\}(�!;ǽ���A�>������9��O������>'G?0�����Ͼ�-���������q?XX�>����oPg�!K[�gal�d�]�m�0��尿�����
�Uk��4���ؗ�����m5b���^��}/?f?����������7C����!��>]��>G,5>��>�9=XX-�CC�4Lg�c;����Z[?��?Î>3I?#5?�mY?��?$�;n�8>oR~�Z\*?<DU>x`�>C�F?��U?�g?�(?(� ?M�:?��v>N����ys���R?d�?� ?A�?�c?"��w%.��=�<��*p ����=�go=�@�=�"]���ý=���=�U?�����8�����wk>�7?φ�>0��>q���(����<��>3�
?�F�>����sr�Xd�t@�>���?/��=�)>|��=��W�Ժ�/�=�T��P(�=���oB;�Ԝ<��=��=��v�Z�p����:k�;x��<�5�>�E&?���>E��>E[��ԋ龊�+�W0�<|5B>w��>n�_=�9׾����7����v�
Tu>5;�?[�?"n=Ǥ=���= ���{�v��K�����p��=���>��?�@,?���?܌-?�a?��=D+��X���$H���3����>�S,?3ǐ>�4�˾�3��L�2�K?��?��`�s?�	�)�ɨ¾��νOk>�.���}��֯���C��$J����N����i�?b �?6�;��7����L�������D?F��>驤>}��>�K*�hAh���Z�;>>��>�R?�^�>��O?K"z?��\?��V>�8�H���'꘿S�i�Ь%>��@?��?��?|w?R��>�a>��$�S޾���^2�'S�چ�4;L=Ǭ`>��>�L�>��>���=D�Ƚ�D��RF��x�=�[_>�R�>�H�>�+�>eo>�"�<��G?v�>?�����}���΅�P�E��Rv?��?��*?D=���O�E�τ�����>�@�?���?�*?P�S�]�=��Ѽ
o��p2o��.�>ɗ�>E��>,��=��Q=�>���>��>�Z��L�4*8�E�p?��E?��=g�ſ��q�_�p�×�>�b<��m,e�d���~[���=���������n�[���������w���ޜ�A0|����>�1�=�,�=p��={N�<*�̼�<�lJ=�7�<G=�hp�7�l<�69��Ի�Έ�S12��eY<F�G=a]��ǚɾ/5}?��G?"�+?�MC?�[{>8">�	0��\�>�}{��!?��P>��J������:>�٧�	0���aپ"�վ��b�򙠾A
>�|7���>g�1>�b�=��<�c�=�<�=U��=�����d=���={¸=ӏ�=���=r�>�|>Z{�?�߆��Φ���w�H}���	,?\�>�O�>�7���9?��v>cx���ſ����S�?��?��?^�,?�	u���>����QD^�0��<S��=�V�>�m>6�q����>hN�>!J�$Н����=���?>@t�P?���=c޿�1>=A9>{>��Q�)�0�[]�'Xh��[��#?�9�̾���>���=��߾��žL�0=�99>�f=0g��[�!��=��v�p�7=�t=33�>�D>%N�=�Q��g��==�I=��=VCQ>L��)�?�r1��>=!T�=Z�c>�0(>G��>3o?O�/?�d?���>r(o�;�H��f��>���=A�>pL�=�;H>q��>`�7?SD?�cK?�Z�>�k�=��>h?�>U�-���m��F�벥����<�ǈ?_O�?O�>8�<�XF�����=��Cͽ@?�%0?��?�2�>����dܿ��<�]�#��:c>�;#>���=4���S�/�����;Ƚ[���Z>1��>,7�>�>��>��i>-�?�ۥ>S�=�2=ҭ�=.񼓳G��ة��p.��ͫ�5tz=*=�Y��z�������D&<�I�<J����Y����=S�=Fn�>�>�-�>倥=2y����?>�ř�f�R�Ӛ�=-���YD��yb���y��+���2���0>��<>]�H��/����?޵V>=>>-��?��s?��>���6ӾӸ���=S��[�[��=�h�=0�G���9���_��L�'�׾��>���>�1�>˿l>�/,��?��w=Z⾀<5��8�>fX��<���*��Eq�T?�������i�͓պ}D?�9��߸�=�~?íI?Nݏ?q�>�9���zؾ��/>����"=Z����p�>-����?�'?��>���e�D�у��[.��>�q�����C����7��P=���4�`>�[t���߾�S��3��Zk����q��������>�:G?��?;��KL����T�������<�~�>.�?K��>ZU?�l�>�ͽ1��-����>!��?�7�?S��?�_�>���=gޯ�L��>�R	?i�?���?C�s?	�<�59�>�X5<?�>#+���N�=M[>C��=���=N�
?��?Q�
?��T#�,���R��]��=g�=ʏ>%Q�>X�u>���=��}=���=xk]> ��>iV�>�\e>oʤ>6��>8���n��9��>��1>M�>�dI?^�>��=�4 �M�>�쁽�C�����]�������İ=�߻��L`��X踚��>�ÿ_��?���=����?�Ͼ�G�"a`>�D>�h%���?�\>}K�>���>��o>��>��>ٮ�=-|Ӿ��>~C��v!�9�B�B�R�^�Ѿ	w>�/��X�'�a�DY���I����[��w�j��K��#�=����<�(�?LI����j�(�)�Ky���Q?�S�>136?�Ӌ�����,�>K��>{�>P�������э�n��5�?b��?��{>O�>�wT?�3#?^	��o�λ
Wk��Y��.B��~~��
����(�c�C��P�5���5?Nr?��=?Uʉ>H�Z>�Q?7��	-��&>a.�M�Y����=/]�>��F���i�X���R��X{�����q`?(�?�!?wg����{`>�$1?3�>?�;m?�?��.?��+�x�*?
H>oC?�?��C?��!?w�?�*,>Jf>��E��v��`�� �v�9:?��z�w=E�=.��=i�|=<s�RS�<a�%�B��{ �U�>�i� ۙ=�[u<� <���=e�>/�]?�?o�>�s"?���Y}Q�s�'I?>酱�%B��EӾf\񾛅 �Ϋb?��?wXi?�u?>%yA��tV��?>�à>+�=�e	>sD�>)d�֢���?>*��>B�o>���<b��~���k�����ì=��=5�?�r(>_����>qƾ*��T�>��Ǿ]��Mޔ���q�l;�HZҽTx�>ʺD?I?4�R�Kb��|J>�r��v_?��!?J�w?���?�g=����J�Ɋ~���Ͻ-i�>�FG�p�A� i��ſ���L�A8F�2pq=��n����s>Z���־Y�[�~�>�7��c'<�}�7�n=)}
�E��'Ј��t�=}*>N�ξ!�"��O������=�C?b�Q=s՚�}�N�N2��!�>-x�>��>	��oܨ�9C:������=:�>�J>-^;��徵�I����<�>�66? ;\?I>x?����}�s�Ϳ����0Y��_�G=h�?G��>c?�t=/��z���<�ĽO��)�A?>&�>�9�N�'���׾�����3���>�6!?˕`>�?5�y?T��>��]?�"?��>��>n�C�I�Ծy�.?~?Ӫ=Q���y�u���8��>��?g�/?$pH���>j�?�a?u7&?�xD?��?�T�=)���V���>��>��N�������>�I?W��>�T?+�?�6>D�*�Du�������=43>S�/?�?�?)�>{��>D�����=���>vc?�0�?E�o?��=��?I42>���>��=d��>���>�
?�TO?�s?{�J?���>���<93��@:���Hs��;O����;n@H<��y=c��T$t��8����<��;v���N�����x�D��쐼��;GJ�>��s>� ����0>��ľ�7���	A>^M���V���ኾ��:��s�=�~�>Y�?خ�>0<#��~�=���>Xk�>���?C(?\�?�#?/�;��b��2۾��K�<ڰ>[�A?:�=z�l������u�\�f=2�m?6�^?RW��*����m?�Q?�Q���T�^^�4����$�%�]?'�?e�齌q�>1��?�ps?���>h�����U�����Y�T�*Eоp��=Yx�>���r]��y�>à6?�٭>�e�>�j>+X�u��3熾]��>�Y�?KM�?�ȉ?B�>]P[�����;����J?��>��h��u?%�2������RF���y�����2��6Z������g�)���'��;QP>w ?��o?3�j?b&r?/���o�8[l��G?�+�O��N�)���֙R�So?��BJ��h���ѾP�������{=
�z�u;�XL�?FG'?��*�0L�>&����I��hϾ9�7>�,�����v�=�.�����<ޟ=�D��G>�Wݧ�C$?�V�><m�>�<>?��^�F>���1���6�5��;>Q�>{�>��>}��;-���Jϼ���s�g�н~=v>dwc?ďK?E�n?����!1�����
�!��R/��j��`C>۱>�̉>ՊW���0&��O>���r� ��Zz���	�K�~=7�2?�-�>F>�L�?P�?�p	��`���ix�J|1�2Ä<G)�>�i?��>�؆>g(н'� �j��>�mg?���>A��>ɏ� �*��}��	ٽ䅇>�nX>��>W^>��=�K]`���������g>T/m?[����D�$R�>�j:?*�[=����l�>��f��Y���^�A�¡�>N?�<�=��,>[���)x�B�s���[�|?+?D�?�j���'�;1w>_�?=M�>�>�}�?�>�Ǻ�oʋ<z ?i]?F=G?�@?U��>��.=�|ʽ��ǽ�D!�v5=���>�`Z>�&}=;��=���X��s�F�l=Uf�=�]�����@<�피�u<�w=%f@>!lۿ�;K��پ��o�9
�������o��Ɩ�1c���!��Bjx���L
'�0-V��Cc������l���?�;�?���*&�����
���V���Ҽ�>��q��~��㫾���+��ٚ�/Ϭ��f!���O��#i�v�e�O�'?�����ǿ񰡿�:ܾ5! ?�A ?7�y?��7�"���8�� >hC�<-����뾭����οB�����^?���>��/��q��>ܥ�>�X>�Hq>����螾y1�<��?7�-?��>Ďr�0�ɿb����¤<���?0�@��A?|�(�|��}+V=ո�>��	?��?>�	1�l2�����u\�>�<�?���?ܱM=E�W��x	�	oe?��<�G���ݻ�%�=�:�=>=?��ҞJ>-R�>�z��DA�Kܽ��4>ۅ>��"���ok^�ξ<��]>�^սe����Մ?�\�bf���/�R��.�>��T?$+�>Ɛ�=£,?�BH��xϿe�\�1;a?\1�?���?��(?�ۿ�k��>��ܾt�M?�K6?d�>�k&�E�t�f��=Κ⼅���J��E$V���=k��>��>�,����~oO�+Q���.�=����ƿy�$��y���=�0ٺ��[���罦Ҫ�ܳT��$���xo�����h= ��=�wQ>�d�>YW>�8Z>aW?8�k?ZE�>�>D�5���
ξ ��O�������������T��߾��	�u�������ɾ[,=�)�=G9R������ �6�b���F��.?�/$>:�ʾ�M���)<k�ʾ����:����@���-̾5�1��n��ß?�A?F�����V�t��ȏ��T��1�W?_g� ���߬�9��=α��<= �>A��=���? 3�`�S�V�K?j"?4j8�^�8�c��=E�+���f��H?'�,?�����3�>#NL?�!�C?���%>���>�+>3R�>m�=�Н�Ƹ���?(�:?z�$�{�>�3�>�_�de��=j~�>U���ȗ�<�1_>�~:=4��	�P=�\���>�)W?{��>Z�)���U_�����O==��x?ٔ?�(�>q{k?=�B?���<Td��C�S�6�IKw=��W?�%i?&�>8��оm~����5?}�e?2�N>�ch�R����.�GQ��#?�n?�]?aZ��s}����g��[s6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������ƕ�=ٕ��Y�?��?Ă���9g<;���l��o���]�<hǫ=##��O"�S��_�7���ƾ��
��ϟ��q��>�Y@@M�Y-�>�K8�6�%TϿ,��n\оqTq���?m{�>��Ƚޝ���j�Mu�#�G���H����ng�>�X�=��߽8���3�}��E��h���3�>�Vɼ/��>:�U�����B�����
�ds�>��>��>�ʹ<��6��?���1տrx��6��^?˜?���?��?���=ڟ.���TҴ;�F?�z?I�g?�����s���%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.���p?�n�����Ǥf�b�g��>9�3=9��{u�=�w>��v��������!�?�,@0��?�R���.�T�&?�͠>N��j���Y�=X[>��?Mٱ>;-|��?�KW��Yl�:�>5{�?Io�?�A�>�0��uU����>A&�? )�>���?���=���>+9�=�<��j���P�&>��>��B�p�?;�O?���>���='�7��*���D�jPO����JB�i�>4�`?�DK?	\>%��-�/��@#�2�ֽk�.�ݠ���8�xR
��7ٽ\3>g=>�>��E�OԾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�|�>(�'��s�(?���F%�d�ؾ���=�5?�ԩ�K�=�%�>Mg�=�@��=p��
=�?��>s��?��?I��>��o?1L��c�����_��E�>HPC?��?��D>?��S��>4�?���눿QJ��s?O@�@\Q?���⩿=�����L�|S����>�x=��Z>�����[/>�"��q<˞V=�T�=3N>��j>R�C>k��>��>b��>
��N!�`���� ��%�h��9O��c���4�>���s�7�Ze��(�)��f���<W�E��檺&�<=�n��o@
>j]T?�Q?�l?v�>5X�k�>��𾁉�=�0��=HF�>�3?cJK?��#?�*�=mZ���h^������§��,����>��H>���>&��>7#�> E�;�R>Xr2>�n>{��= =]k�&J=ZZ7>yJ�>I��>�P�>�C<>͑>7ϴ��1��`�h��
w��̽,�?b���I�J��1���9������i�=8b.?�{>���	?пn����2H?!���l)���+���>|�0?�cW?�>�����T�;:>��Ʀj�`>�+ �=l���)��%Q>rl?��e>cUu>[�3��A8���P��L���8|>�6?A.���H9�Ԧu��H��Fݾs�L>Κ�>�:K��x����J��h��y=�r:?�~?Cd������ZRu�[��$�R>N�[>��=�Ԭ=Z_M>$c��Ž�hG�O�.=A~�=��^>��?�6>�ģ=Dƣ>kϚ�f�P�ቡ>�`K>{�=>G�;?��'?��4�1�����{��?,�V�~>]�>a��>�C�=0�J��;�=}?�>� e>[5�ŭj�����S��QM>:�u��WM�+�R��K�=������=n(�=]���&<��!=AS�?���V�ƛ$��1x�%�l?7s[?���=F9>��9��"��x�վ,7�?A�@�[�?�\��"�L����>�Y�?�����>%�?���>������eF?���� �و��Y�WY�?���?�`=)C���D����>q�)?Ǚ��Oh�>yx��Z�������u�t�#=S��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>W�?���?h�m��A���@����>:��?�gY?qoi>�g۾;`Z����>һ@?�R?�>�9�~�'���?�޶?֯�?�>9>���?e�q?�R�>�Gt�K1�ޭ��-䉿�>=l��BX�>��=�!����F��*���)����g�����j>  =f,�>Iܽ�;��6+�=ɋ������Ĥ��`�>��u>��@>tF�>�	?���>��>��<괶�P�������KXV?"��?����_�Z�ў���|�<�E^�OH?��;?A;,�����%�>��V?}v?�OG?'�>O��럓���ȿ�2�����<1�4>�d�>#o�>m;��.�L>��������e>&��>� I;#����)��<�Ɵ>}[?���><C)><m"?�+"?�>|>a@�>]H�p���.k@��w�>y�>�-?\?8�?�/����2�Qɒ����<*[�B>[�q?��?#2�>�����b5����	L̽�+�?�Kj?����N?}i�?�;?�pC?rt>������ǾP`��ҧ^>�"?����1A���%�m����?�?'��>4ˎ�5�ֽ;Ҽ�����	�?��[?F&?@����`�/�ľ&��<����`�@=�;eP,��r>K�>Kӆ���=�>.�=R�l���7�`=\<��= ��>lT�=@15�cO���<,?Z�G�,ۃ�e�=o�r�OxD���>�IL>b��m�^?<l=��{�����x��\
U�� �?��?Ik�?�
���h��$=?��?5	?_"�>�J��B}޾���Pw��~x�Fw���>���>�l���U���Ù���F��5�Ž�6����	?�R�>7I�>��
?��)Kk>[�y7Q��޾���8�C������<���M��QL�)1羳�x�I�|=�e}�DZ�fz>�X�	4�>�\�>��>#t�>N��>��=�ck>�8w>~�>��e>آb>Ʀ>f�
�U�ݖ(�/GR?'���~�'���農���7B?ϧd?`�>4i��������c?��?���?��v>q\h��+��g?L�>*G����
?5�<=V��І�<����V��0W���4�ێ>ֽً
:�b"M�Phg� .
?�?�?���n̾�+ؽ:/����w=���?��(?�(��7P�M�j��5T��#R�_���c�7��=� �W,p�Y�������^��9y(��2=�,?H��?� �BS羭߲�yk��?��_>Zy�>�>�&�>A�\>g���$/�p�[���%��B{�~��>Q�w?�>�yJ?`C?gcH?T�?��>=u>�婾W?�͐���?4f ?g=>?��/? <?]�?��?�?>�6r�c� � �پ:7?��?6�?��?��?�t��a�^�2�q)���8���L��{v=s;�`����H <�sB>9d?g�%�8�=�����j>�n7?�m�>��>�ޏ�0>��B�<W*�>��
?	F�>����Nir��a��g�>��?����=��)>��=u����Nͺ�=�ü@��=t`����:�HX <�J�='�=��n���h?�:��;	��<s��>NX!?7/�>���>C��IT��#���=�m>�9L> 9�=���_Y���I��t�i���n>�]�?#��?vƇ=�y�=���=Z��I$��N'����þ��r=!�?�?��I?��?FN7?�q?PT >c�"�[����w��꡾�
?:!,?���>�����ʾk򨿲�3��?�Y?D;a���1>)�ߐ¾!�Խq�>�W/�-~�}��PD�dS��E��=i����?��?�A�"�6��~������`��'�C?j#�>�X�>w�>\�)���g�8%�R4;>j��>rR?4ս>3P?({?�Z?J�K>7�LY���ǘ���|�ƹ>9!B?(Z�?#��?IXx?5��>8�>��'���ݾ������-�K��*����d=��W>��>�]�>{j�>N�=��̽�z��s�<��=Z(c>N��>�*�>��>/}r>�J�<��G?���>9:������ߤ��̓�*!=���u?���?z+?�Z=2W���E��*���2�>)c�?c�?�-*?�&T�z��=B�ռDҶ���q��.�>6Թ>�'�>O�=��F=>>$.�>h��>7|��X�HY8�X�L���?f%F?�L�={�ÿv�(������_`�d�q>�(�� [�����K�꾷#�=zɟ��	������Zt�2㓾��ؾ���e��U�>L�>���L>@�>`�f�����R�=i�= ��=K�q�=����">Z�<IA'�o�¼Y(�=I�.<M<�x���ϾY�v?+F?��#?k�J?�d>�%>HS���~>*u�a�?��T>�-P<%��� l�{o��!f���>ܾ!%ξEy?�V럾�y	>�AA�n�>�KO>�>�/	=�<>�=�"}=�=���+=)�=G��=L
�=�W�=s��=�>�q?�d�������J������?�I�>)<>Z�̾sR�?��N>�v�K�ÿ{2�d��?k�@���?�?���Ċ�>c�۾ŧ��U�<=���=n��>H�>-<�<�>s��>5R�l����.=e�?M@F[?���j �mI>	�I>�>cM���-�R]�Dg��Y�,%?��3���˾Y�>���=��ؾIE��Fi=x�5>\�:=G��ž`�7��={j�\m6=�]=,��>�F>2��=�����ܿ=�	2=�4>
5Q>B���jQ����caH=�0�="�r>n�A>-��>A�?q]0?POd?�#�>�n�� Ͼ>��>W�>���=�F�>�,�=�eB>���>��7?ŭD?�K?���>&�=k�>��>�,��m��S�w������<\��?�Ȇ?�ĸ>��T<R�A���R_>��"Ž�p?�L1?/u?;�>�U����9Y&���.�"����k4��+=�mr��QU�L���Hm�3�㽱�=�p�>���>��>8Ty>�9>��N>��>��>�6�<}p�=3ጻ���<� �����="�����<�vż�����u&�<�+�8�����;w��;U�]<���;�B<&]�>*��=΍�>�>4���oo�=i�оO�S�;J$>�ɱ�
O�G�e�Whl�k,"�R�d��
>�x4>`F���^���3?8��=��j>���?��`?8��=I�ý��,���V�Pn��<g=�'w=�T����I��9^���J�������>�ߎ>��>_�l>,�<#?���w=�⾷b5�e�>�|�����)��9q�@�����3i�n�Һ�D?^F�����=�!~?<�I?N�?\��>���H�ؾu90>H��/�=���(q�8i��<�?T'?��>�쾘�D�VD߾�7�G��>�Ve���Q��Ζ���*��ﰼ����I�>W:��+Fþ�<=��W���x��h�;���)����>L�O?��?�����烿�a��w��F�6��>�3g?\�>���>x�>��ὸ�
�O͒�u��=��m?���?���?^��=���=�
���<�>H+	?���?ݷ�?��s?u?�z�>�;{� >б���X�=��>�z�=I�=3q?�
?�
?d��m�	�������C^���<�ԡ=+��>�l�>\�r>���=�g=t�=�+\>�ٞ>��>��d>��>=R�>��ᾗ��f�?Ы>�~�>I�0?�>�>�I��}:�}�<E���dMx����r�����x�h�]����(��;߼��>�����ܛ?T�>W��ւ?�����+佑�>�23>���u	?E�E>�LQ>�~p>��>C	>;��>�^�>�_Ӿ�>����T!��C�lR���Ѿ�z>������%�E������RI�7j��eb��	j�-���;=��S�<L=�?�����k��)������?J�>�6?�׌��鈽��>i��>M��>�F�������Í��`ᾟ�?���?	�=���>L�D?g1?�n^�� Z�6~�$p��aG�N[�e�N��0��>�t�$$��\��3O?�a?�E;?�H}=��>�܃?���hț����=�,���G�©3>��>,W����y��^󾷶��qW����=�L?���?��*?�)������2p�>�A?R�3?c��?�S?���>�[�;�7?�m�=r�B?�y2?$�O?��?��>e`=�=�>�%�)(j���w���5�����fmֽ3.>��;4=8��$��ޑ�=cu=.o ������:��eRF��$O�7a>w�=���=� �>�Z?տ�>!7�>��?�!g�4!S����LH?��\=E䈾m`��~����<O��/R?��?v]?�:n>��1���2��|>��k>�'>F*>���>���K�F�3=�	D>�J>18�=�L��h��3��sG���ȼYX>"��>H��=BB+��q���pS��T!�>=zоD�ɾ����q��o0�T=�)i?�^?~4?\_K=�����>��}��dT?��&?_W{?�Ց?��o���Y���q���j��m= �>z4M��<�.��뷸�"C�UP�"�>A���U���a>��� ޾�m��WI��c羫�A=���mV=�1���־9��U��=)
>�.��G3!��<��֟����I?}�`=FS��S3U�(к��>�ޗ>���>�P6��!y��e@�#�P*�=���>�:>? ���H���F�����<�>�JE?`Y_?m�?�*��7s�*�B�@���W��QOƼ��?U��>n`?��A>k��=6���?���d�G��#�>���>����G�=���,���$���>�>?�>5�?��R?�
?ϕ`?�*?�B?��>7��<��g�&?i�?�.�=�ཆxQ�b8�N�E��d�>q�)?�S?�f��>y�?6�?�L%?�O?�2?�7>TG�D��ӓ>_?�>FrW��}����c>[�J?�ñ>3�U?���?@�A>y6�����*>���r�=Y >�r2?��$?�7?.T�>".�>��?��ɗ='��>�_?I��?&
r?�c3>� ?���=]?P�$>Wm�>1��>2��>n�4?�h? �S?�c�>]��<�i��K=.��1�%<lH|�[5Ӽ�Œ;Ba��y�ý%���H<�w =!�v=���<A4��K�8�hO=�ʼ9B�>��o>�-��AW,>�ʾ�Y���TA>����M����$���F����=mg~>�5?ѕ>9	'����=��>d�>�$���*?x�?r�?&����}a��fܾ�.M��-�>\R@?���=�Rl�K����v�A�U=ǁm?oW_?�'M��A��Kc?��E?Ɵ����*���ʾRָ�������z?�c
?�J̽�h�>��v?��i?���>iċ��{W�A���?Dy�*�վ�`�=km�>��#�m�{����>1h)?0�>>��>k{=�-��xފ�2շ���?1�?zֲ?ܭ�?i3>4�R��V�J#�}���uQ?a��>�û��(?�>a�ݗ���D��ˮ������ļ�����v�v����a��T��&9�t؇=��?"q?�Tq?�XM?�1"�mg��Z�Gh��M��o��h���O�'�7�}MH���b����d�žH�=�G��=��~� �?����?<m'?B�/����>����p���Ͼ=FB>����������=�l��%�:=!7=?q���/�B����r?YK�>LC�>��<?ڿ\�޺=�+80�Z�6��=���Z3>�F�>A8�>eb�>t�~��/����qƾ��~�m$��(Ms>}c?ΡK?�o?�O��x�0����Bt"���L��ħ�I�>>2�	>���>��[�����&�Y�>�>.q�'�����I
�ʫ�=�3?��>��>:2�?�d?Y��o����_}�E�/����<�#�>��h?��>�z�>�Wֽ� �Zu�>�g?4��>Ɗ�><�����!�%p���4�jRl>~��>}�>qU:>E3��Kc�����튿Ū2��">��8?=���L����|>/Fj?*�=�&==�>�.U���%�߷���q��m+>�?��>dݐ>�5޾�z:�s�H���?�(?l�?�����f)�V2�>z� ? ��>���>�]�?U@�>��Z<h?T@]?��G?yH@?Nm�>�a$=�����Bɽ�$���.=��>s;Z>��w==n�=q���Z�� �0�I=C,�=:��s3��d��;	c��3�Z<J=j�7>���B�U��E��=7�߷����I�������f���ㅽ�I��M�����w��9/�� ���G����U���������?"�?Ӛ0�*W��䰕�`���D'	���>������<>5þ�g�����e����ľ0<�1lQ��:i���k�G�'?�����ǿ��:ܾ2! ?�A ?%�y?��3�"���8�� >�B�<I,����뾬����οP�����^?���>��#/��f��>���>�X>�Hq>����螾	1�<��?2�-?��>Ŏr�+�ɿ\����¤<���?-�@�vA?��(����V=���>�|	?0�?>�0����
��$_�>:<�?��?��M=B�W�R�	��ue?7�<T�F��l߻�@�=�P�=�u=��HaJ>X�>���XA�S�ܽ.�4>��>+L"����b�^��C�<��]>h.ս\��'ӄ?��\�~f�6�/��g��}�>��T?��>���=��,?�RH�~pϿ�\�'Ga?�/�?>��?4�(?Vÿ�V�>��ܾ��M?=A6??@�>r1&���t���=b|���_㾝V��E�=�5�>��>d�,�_t��?O�O✼���=n�ڹƿ~�$�/~���=K��\��罧ઽ��T�"���ro����oih=n��=�mQ>T`�>W>�Z>zdW?�k?YW�>3o>(Y�b���}ξ��V����� ������}��Y��߾ɉ	��������ɾ�!=���=j6R�6����� ��b���F���.?�q$>��ʾj�M�Ao-<�pʾV����䄼�楽/̾��1��!n�͟?X�A?2���C�V�����c�����(�W?lQ�B���鬾<��=溱���=�#�>[��=����3�k~S�(�$?��0?��u�ꤷ>񃾔W>i�?��<?������>H�f?�/�s����p_���M>~��>�>��>�栾��W<γ>�??U-b���;��>?@�� �*��u��l�>�]f���C>��/>��O�����B=)�<]�>&�V?r��>`*�r�Ս��2#��~A=�Lx?��?¯�>lvk?UC?쯶<�|��r�S�L�
�3q=�6W?��h?{d>�;���Ͼ"��B5?\Pe?̍O>Ee����e/�M�PA?[o?��?�����}��͒�^W��v6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������ٟ�=>ٕ�oZ�?��?����C9g<��.l�No��t�<�ū=��I"����R�7�b�ƾ�
�����O޿���>Z@�P轣+�>+I8��5⿴SϿ���7[о^Tq��?�~�>ϡȽʜ����j�4Ou���G�,�H������=>>a����t<N�þ�%q���h�?_<���3?��]�d�>�l���\�����m�LN�>	�>�?���>)����ү?#-���;e��'�Jz?���?%�{?�]Q?쒽0:��0��W�Y��S?(�?d��?뇃=<@�����<#�j?�_��uU`��4�pHE��U>�"3?�B�>M�-�*�|=�>���>'g>�#/�x�Ŀ�ٶ�7���Z��?��?�o���>r��?ss+?�i�8���[����*��+��<A?�2>���F�!�?0=�QҒ���
?T~0?{�d.���t?���с��;T�� ���?�s"<��½��=pI��/]�I����|��t��?=@1��?�#�h����?�s�>ͥ<�H~��pЫ�4|>mr?���=��8��_�>��U���d���R>l��?Y@���>����W~����&>9��?�>(�?B�=���>2��=�ɯ�X��v$>R��=��G���?4�M?�>���=�:���.��{E�6Q�`��+C�:��>�a?|YL?��a>�㷽~�0��� �L0ͽ1����!?@���'�A�۽l5>i�<>��>��B�0JҾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�E	?W$��J���]~�P��+7�9��=��7?J6�R�z>���>��=sv�5���u�s�泶>�C�?0}�?S��>��l?2�o���B�â1='B�>��k?�y?�Rg�o��_�B>1�?�������NE�'f?%�
@Ru@�^?V颿�ܿ�D��A���X���@�=L�>���=?�����+=N�[=��="m����>�ہ>K�X>�q{>�,>BY?>�$>_���\�!�/��6p���ca�dR.�C-������{E���1G��оX��@�g����z�����������=��U?�R?"p?� ?��x���>0���e#=�X#��f�=� �>9\2?��L? �*?�^�=�ʝ�E�d�LX���9���݇���>[�I> s�>o5�>&�>Ǎ�8O�I>�e?>�e�>O>&0'=H��8A=�N>�2�>h��>o��>�C<>��>?ϴ��1��^�h��
w��̽2�?p���H�J��1���9��Ŧ���h�=Bb.?|>���?пj����2H?���w)���+���>z�0?�cW?��>	��$�T�:>��Ϧj�4`>�+ �fl���)��%Q>nl?]7>�P~> �:�o�1��s=��j���`�>�#?�2ؾ���!s�2�Q�U�ھ�CD>�\�>w��ş&�����ѯt��]k�2�?=��7?�
�>��b�I6��W)�� _��l�j>8�2>jw�=���=��=>��N��j����N��G=�/�=�O>N�?��F>��K=���>F7���B2����>&F[>:g>�5?v�*?fԏ;� �������I�m!u>/�>m��>�[*>WAC��V�=L�>�y>�����j�����{i:���c>BS���\��Ql��)k=O�+N�=P~|=8������,�<$�?�L���0���zH��4���?�6?�	>%�<��Y��ծ� R �EA�?@6��?E߾{j]�(�?���?.�$�LF�>|��>���>I��YM���?[�D��w���!���Х���?B�?�wнs����'W���2>���>�/��Ph�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?pYF>� �?&t?��>�l��8/��p��i�e�i=4.�;���>��>/׿�{�F��V���O��uk��V<b>�
#=�+�>{�ڽ#ָ� 3�=�)���r��l��g�>Pv>� G>"6�> ?	
�>j�>C�=0=���끾�����O?��?����V�i�ࠈ=�'k<{)�� u/?q�??¦�=�1���D�>�D?��W?5�9?�z�>�{�#����ѿ�
��Zp�=%��=qջ>�s�>�g1�	V>�6��5\���>�]>�ML>����5c��P���>#??�S?.�>T?T?J��>���>��Q�@|���\K�Z�>�-�>X8?(,t?�$?s���:�E�](�������i��?�=�i?�c'?��{>�Z��g���,��7����8��}�?�0k?u��[I?�Zv?�;?�6?�?S>à}���Ⱦk��7R=h�!? �W�A�H&�|��(Z? ;?L �>�r��g7ս�Qּ����=���?6�[?�1&?���G'a�T@þ���<�!��_����;��?�N�>2~>3T���|�=bY>x:�=�{l���6���d<�	�=�~�>���=��6��A���<,?��G�ڃ���=i�r�6xD�^�>�HL>L���^?�l=���{�����x��3U�� �?Ӡ�?Gk�?Z����h�Z$=?��?�	?�!�>WJ��|{޾Q��-Rw��}x��v�*�>u��>6�l�P�R���򙪿qF���Ž$�u�p{�>U�M>ʰ?{(?�JD>,E�>�� R������@�h�g�+��%H �"�����AP��̾�pDK������g����>���=Qu�>BJ�>���=V/�=[m�>*�<`��>��>�0>yo�>.X>Ϛ�=M��;�׾��e.�I�R?P�˾�+����MҾ{E?�l?��>��nP��tH�2|?��?�?p�>�a�!7)���?�I? ���y�?�w=)�6=�dx=PȾAx"��:�[����I�>
;۽,�0�W�]}��ʂ�>��?��V�\)پ��ؽ�߾q��<D��?��G?(����[�rYX�A�`��S��'Q>�����o�Z��x$u�L���?��w苿Z�-�\�X=Mo0?�IN?�˾��޾��;;[�]�2���>D�?*�>�(?�o�>��[�2�_�c��`3���5��z�>[/X?hw�>��O?��:?�"P?=D?���>>�͢�(?��T��	�>�F�>��B?�#+?��?�?�,?�Φ>��p����zھ�|
?3�?v
?9�?���>Ŝ��P�!���;�
�����ݴ��)x�=���=�{z�?���~ ��>��?_�=;��Ǿ�\�>Vk?~l?�/�>
Լ���?�`>DE?A)?�d>[d	�͐M��0��w^�>��?{�L�Ջ��Y�Q>���=���=]�>(j=�+ >`>������v��=��=���V�<=ZT��!a=z��=�A�> &?���>��>�������5�O�_=��>��>CU�=��׾����Շ���t�?�> ��?���?��
�0	e=���=�c��-��yR�m�����Q>���>��>}T7?!.�?5�3?`)?�*�=wg⾢]��)����	��Z�?� ,?2��> ��f�ʾl�J�3���?CZ?�<a���<)�)�¾�Խ��>M[/�M/~����D��������z����?���?�&A�Z�6��x辑����[��ғC?� �>X�>��>a�)��g��$�2;>��>SR?7#�>��O?9:{?S�[?DlT>��8��/���ҙ�Z�2���!>�@?ձ�?�?Sy?`q�>	�>-�)�i�lQ�������&߂��W=uZ>7��>1(�>e�>m��=�Ƚ
]����>��m�=-�b>2��>��>���>*�w>Ep�<�MH?�:�>g4��P���;��s0����L��u?���?%.?��=��pG�s���U��>%Ѧ?���?K�%?�!p�$��=�ت��ܸ��e�NP�>�G�>'��>��L=6�[=�S>���>-��>�i&��¿6�+?;��\?EkF?��>���f�#!j���h`=��u���W���"懾hc�=��~�7�%豾A. �W"��-ݩ��Bо����*���2�?RN�<=�g>>�=?����2���jU<�]?=�<4<���B0-=�����:�����Y6����<#>�}=/�žZz{?�C?<.,?|�@?z�w>�&>�)'���>ꍅ�b�?�`>�����\G�����1���)Ѿ��Ǿ�l`��۟��7>_ ޼�d>	E>�Z�=a\�<&*>o(�=2�=�3�;'/=aĿ=u��=à=��=?>�>�x?���������i��EH��-!?���>oZ�>/q���.H?�
>U_������b��l��?S @���?��?��v����>����dҥ��=�#F=��>�/>`Yd�>���>���;a����$;�\�?J� @��I?]���ٿ��>\:>t�>.%R��V1��V��[d�CY���!?l�8�&Ⱦ��>�r�=v�߾��ž�#=��8>�/_=����\�ʏ�=�"y���3=�lq=0)�>,p?>��=q>��	�= J=���=�%Z>�h-��j6�e�0�L�3=�v�=}e>+^.>%��>��?�`0?�Od?f+�>�n��/Ͼ]<���?�>��=�.�>W=�EB>倸>W�7?�D?��K?Z��>Y�=��>��>1�,�y�m�W微֧����<P��?�ˆ?�Ҹ>�Q<;iA�P��Af>�vŽ v?Q1?0k?b͞>�U����9Y&���.�$���_v4��+=�mr��QU�O���Im�3�㽯�=�p�>���>��>7Ty>�9>��N>��>��>�6�<zp�=dጻ���<� �����=%�����<�vż�����u&�;�+�5�����;z��;a�]<{��;�o�=���>��=t�>�Տ=[��r�C>>͠�X�R�{�=�8��XLG��j`�2�w�R-�;^5�1$>��1>)>.�_���M?�CK>��@>U�?t�n?��>\��3 ؾ6���P�:��r�h˶=v��=�R��*8�Wa�>�L��bݾ���>��>O��> �l>��+��?�ox=�/�r5���>�������a)�[2q��6�����i�p�ݺX�D?�@���r�=�~?ݵI?hߏ?~�>⶘�e�ؾ50>]&���v= �9�p�PZ����?d�&?M�>����D���,��׊�8o?y�u�R�1��e��EM�_��=ZQ���?�&q�;�SKO�[y�������7d��iG��h�>v6?7,�?6,���oQ���K���{�(��d�>�V�?ae�>��>��>��B��R���҃>:�?_��?���?�bM>���=�}��#n�>��	?�Y�?�F�?ۏs?��7�i��>-�2�i�'>�Ӈ�~��=^�>�Î=��=
�?�?lK?na���������=]��w�<��=騎>�	�>hn>}��=ƺ\=c��=�Y`>�Q�>��>.6f>7%�>�D�>�<��� �_�?���=i�>O�0?�^V>y����2�<�ུ&{�;xV��{��.��'s��ӽh�=���h��>��ƿ���?>`4���?;㾀V�&�o>�H$>;x6�M?�#>Uu�>/+�>�}>͘>�n�>Q�@>X�Ӿn�>���f!�fC� zR���Ѿ��y>��7�%�����K��8�I��_��Y��'j��0���Y=�ѽ�<�G�?]���Wk���)�]���9?"/�>�6?����w��I>���>�x�>.j���}��P����+ᾶ�?���?{�Q><E�>��I?��?oؾa���t��vg�
�A�w�M���o�o:���/�����Dݮ���Q?kzn?#�:?����U�]>~rq?��ž����v�>@� �RNc�:�<>>ѡ>v�H�ƫH�+ڇ�cuᾊ���,f<��u?�V�?�j?��Ծ��;]�>�w?��??�v�?��@?fb?����!?��޽�Z?�*? �T?d?)gw>�d>��>��<�>B0�����m�Ƚ͈��9��8�t|�9=��~���9���Q=0�=ψ�����D0��K�<Yaؼ�0�<�i���B�=؁�>)[?�v?�O>ɶ"?�Ё�Z]h�:ҭ��?T��<0�����.~ܾ���Ƽ��s?��?�)b?�b*�7&;�D��qu9>{W�>4�=;>�.�>����=��4�=��>]�U>�|�=6��񯰾����"���Ԅ=�֪=�H�>��>������=O
о�"�j��>3�������ĸ��o��:���c��>`kH?�X?s+ͺ���">�2q�F�s?�?PyY?hH�?-����;�IZh������>�Џ�ǭ)�R��(��[�G}��s<b����ʢ�TF_>�p�~#ݾX�n�q�I��>�qE=��zN=���Ծ��~���=��>�$���� �-ꖿ������I?;g=t���wW��緾'�>j��>*n�>~a?�Ju~�4�@�����D��=���>��=>�ʙ����G�]��s�>Nw,?� f?>�?��	��@��^%��ݾH?ʾK�d>�F%?w��>V?F�e>m���8�����Ys�dU?��=?��>�c$��@�"���>	��
X����>U(?�Q=A�+?*:E?���>xyG?��?Sd�>�_3>*���*����1? �~?8G�=7Fb�Ɇ���8��@Y���:?�T?� W�BŜ>�'?3t+?�=?<�>?�/?6�=^� �o�P=s>��>P�V���锆>��f?ta�>�:A?�ސ?tv�>�=:���-��8z<�{a���.>�Q?ʁD?m�-?O�>0O�>5D��Ѯ�=S��>�c?D2�?��o?�u�=�?Ka1>*��>�Ǘ=�"�>cy�>!�?�$O?�s?l�J?��>���<�����j��͆p�[��\�;��4<�{=(d�
	y�(���<l_�;���a�s�Gn�h>���+�;��>��j>pY���*> jľmn���AM>[��L&��������E�S�=O�>ҟ?1��>v�"��Ԉ=̣�>X��>�F� y*?��?�?�?g<��a�Z.۾�UV���>�4D?Mf�=<1j�!���'|x��K2=�7l?U�\?jBZ�r���ێc?KQT?�e;n�0�u1��!t������,Z?�	?n�G�$�>ʊ�?�jh?��?��`� �v�j����l�l��XA	>��>���*�x�UC�>��E?o��>�Q�>0l�>EA��Wu����7E ?�ԁ?�?1�?:>�`\�F�ܿ���4����X?0'�>�6��b� ?�@S�akپ�'��oI��xv־�˛�*姾w���r����&��
���ӽL�=�?Y�g?'�i?��\?m)��@]�U�_�^�y�$=Y��:�-Q��jH�'?�~t?�s�j����c��5k��޶i=�S~��<4��?�K)?.������>����v)��S;ܾӇe>�ٛ��d�!��=!<W��=��;o���X�#D��ܑ!?ڮ�>�)�>��;?��V���F�*�6�P+(���/Sd>��>��>���>�;_�N�<���iP¾~v�^3���eL>��e?�]Q?�s?�D���/�ejm��q#�������Ѿf_>.�=�߈>�s��; ���+�{�:��p��
�A������uh�=s#!?}��>'u>8�?��>��ʲ�p���q,�G�U=�]�>�i?]�>��>Ns�3�1�16�>�n?��>�ݾ>
���6�Q�s�(�����>+�>�
�>|�d>�;:���[�2���N���O%��S�=,�_?YX���D��?]>BT?���;G臽�d�>���'����b��[t>�?]`�=�}>������(��`�����!`)?;`?VT��_+���>�� ?��>&��>]�?u��>ہ��|'_< $?�+\?��H?��@?ā�>��6=��ɽ��̽ׯ#�V)=^�>�>Z>�M_=���=[��h�`�%�tM=B<�=m��}#��X��;��üR:�<b�=��;>�kۿ�BK�ؖپ���-��@
��ڈ�SƲ�\�����,N��6	���Ux�����'�V�@>c�������l�Z��?�2�?�V���9��9�������9���ΰ�>|�q����. ���.��A��"��E���Q]!���O��$i��e�V�'?�����ǿ�����:ܾ>! ?�A ?8�y?��8�"���8�� >�C�<�*����뾨����ο>�����^?���>��u/��n��>ʥ�>�X>�Hq>����螾�0�<��?2�-?&��>��r�/�ɿc���J¤<���?.�@}A?��(����
�U=:��>2�	?u�?>8J1�sE�f���VT�>�<�?���?ZpM=+�W��	���e?��<O�F�J޻��=.8�=�R=m����J>xT�>Ӈ��TA��1ܽ��4>Z܅>��"������^���<Z�]>غսf/��<Մ?O{\��f���/��T���U>��T?+�>I;�=��,?#7H�X}Ͽ�\��*a?�0�?��?�(?ۿ��ؚ>_�ܾm�M?VD6?���>�d&���t���=�9�|��E���&V�%��=V��>L�>��,�֋���O��N�����=����ƿ�$��\���<���Z�����v��|�U�u֟��o��o�nf=��=�rQ>=8�>s�V>3�Y>�\W?��k?���>+�>S������;b��N���=��ˋ�!���F���7�B߾�h	�>�������ɾ�#=�e�=?4R������� ���b�5�F�g�.?�v$>��ʾN�M���-<�lʾ�Ū���ܥ�j-̾=�1�mn�̟?��A?����V����T��Q���W?�K�W��笾�]�=9q��]�=f-�>��=����3��}S�e�(?Ix3? |��8���F�^>s�N���\��<B?d`.?�g>3>�>? e?$L��\���6>��G>D��>@��>�"�Y���y�˽�

?�6i?P�i���i�>Z�þ�K��/3ӽ�W9>/.��)Ṽ�a>��<Ԍ��U��q+ս[I>>'W?��>��)����\��6#�e==p�x?S�?\3�>�zk?��B?�	�<kj����S�B�ʟw=��W?�$i?��>�����о�u��{�5?��e?��N>Idh���|�.�R�Z#?V�n?�\?�b���v}���{���o6?��v?s^�xs�����L�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?d�;<��T��=�;?k\�>��O��>ƾ�z������6�q=�"�>���ev����R,�f�8?ݠ�?���>������{��=k֕��Z�?��?���Wg<����l��n���^�<o̫=i	��U"������7���ƾ��
�m����ƿ����>�Y@�\轷-�>�D8��5⿍QϿ���\оVq���?���>��Ƚ���}�j�KRu�Y�G�r�H�ڥ��c�>x-<����,Vľo:n���N�{x�=�p?��<y">!8�
�ھ3�پ���m��>���>;�>Ţ�=��Ⱦy��?jT�j�
���m��Ӌw?���?v"�?N�?c�
>�6���ž���Y�/?O��?�[?Y�=��,�p	�&�j?�_��xU`��4�uHE��U>�"3?�B�>R�-��|=�>��>6g>�#/�p�Ŀ�ٶ�>���V��?��?�o�&��>r��?ys+?�i�8���[����*�+�+��<A?�2>���S�!�K0=�`Ғ�¼
?S~0?({�a.���v?sM������WZ��T�=�A
?\���ޱ|���N>H����/��ޛ�O����?�@\`�?#�5�&G�=�?�)�>�ⅾR`x�ʁ�<���>"R�>1�6>L��d�>��$�ͮ^���>�*�?)T@���>���P��֕D>M3�?���>J+�?�y�=4��>��=�l������">]s�=v�3���?s&L?Z��>h�=Ќ9�0�.�?eF��Q�����C��V�>�Ia?w�L?Ub>���&d;�ho ��f̽v�/�g¼��@��e(����4>,>>V�>��E�RbӾ��?Mp�9�ؿ j��"p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>B�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji���	?J���(��%��� �?�ɨ>#�:?����u>R�>x�=�w��B��M�k�nĸ>��?C��?���>Ӓo?#�q�Q
J����<�ƫ>�r?�?|J�;���&�Q>�?��ɍ����yj?�%
@=x@+1X?�O��������@���`Z"�)����ы=k>B0���>�>�E0>��*>5v">�%>���=�>�,�=B/�=U�l>,�}�����Q��x]~�;䆿�c�M���`¾A����b��K�|�[O��g����F�轇T����j��=<�r={�T?�`?Z}e?R�?�7��7�>�������u/�s5���>��!???�>?��J��Xgq�Ք|��݁��*��E�>�:>���>!1�>���>�=�qW>TY�>졛>��|>b�="�n=�켬�J>t3�>>��>�+�>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?Էf>�u>v�3��c8���P�)}���m|>�16?�趾E9��u�*�H�}cݾBM>;��>P)D��k������kri�o�{=%y:?�?�)��{䰾�u��B��MR>7\>�R=�^�=�RM>�ec�ÿƽH��h.=R��=�^>|�?�d->��=��>�g���~N�@��>��A>B#+>��??V�$?�^���\����-�nv>���>��>:�><�J�:�=�!�>�Lc>6H�ك�Խ���>�!V>�i�d`]�ܳw���y=@ܙ�Dv�=�4�=�! ���<���#=�9�?H���T��UT8���x��o?�1?m>`��=7�B��l�� 1󾼁�?s@�Ǧ?������P��!?���?����>�-�>���>Z���G��D\?�<���%
�w+ݾ����`$�?�~�?#�>��Z��]J�W2>��?{�Y�Ph�>{x��Z�������u�w�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?��H>w��?�s?׈�>dCw�cZ/�$��-����|=P�&;��>�0>1���)TF�#ē�#p��εj�����Ja>5{$=�>���OM��@ض=�����䧾d�g����>�nq>vI>p^�>�� ?s��>%��>ë=Lԋ�~���ٖ�utL?��?I�
���p��=W��=�㍾�	?y(G?͢�<�����>F5b?�s?�pS?-H�>m�z	��g¿&����!=A�0>K
�>�)�>(����7>��Y)����>��>��=�/׾�P��ſ�����>^�1?���>?��=ΐ ?Յ#?k>�R�>;6E��M��2�E���> G�>q?u�~??�b��A+3���������#�[��TM>L�x?�o?���>�������KtS�YrJ�������?��g?���{ ?�!�?�\??h�A?�Ff>|\�ؾ����o?�>��!?��4�A��M&�2��~?�P?��><8����սiHּ��������?�(\?mA&?���,a���¾[7�<{�"���U���;f�D���>+�>�������=�>ذ=�Om��F6���f<�j�=��>L�=�.7��u��*5,?�\E�
���P)�=�r��lD��>)=L>��'�^?tr=�v�{�B��xv���"U����?s��?�f�?-ٴ�#�h��!=?��?d?��>*V���I޾p���Zw�$�x�g���>� �>'m�o����������J����Ž��I��?�t�>��?�?��)>���>}��;�7�6 ������RT��= �!Z"�%��".��þ�`�8���6��������>�l?��&�>��>j�x>��O>ɕ�>AX�=XZ�>?	B>0�x>Og�>	�O>[F�=;8D=֝���	A��U?i]˾��)�7��Չ����??�*i?k;�>��������/~?H��?I"�?��>7b��)�K�?��?ʉ����?�=ɾ= ,=
�ƾ;��� �O�^����>zԽY�-�6�X��+�����>��?�ٲ���Ѿ(YŽ�M��]�v=�t�?�>)?��'��XR� 0m��pW���S�@Z�K�f�1���"�G�n�n~�����ʃ�܎)�wr(=	�*?E��?���&������fl��.@�7j>���>��>k�>%/N>����0��o^�,�&�L�����>["z?|j�>h3I?�<?o�P?ThL?SM�>���>8A��L�>���;*c�>�)�>�A8?#~-?¡/?��?��*? ob>T��:���C�׾xq?��?��?�??����F.ӽ�ɼ�I��J�z�5҄�ك=��<�սW8[��Nb=�HT>MX?8���8�!����k>i�7?q��>��>���+��I�<n�>ص
?hF�>3 ��}r�0c�V�>���?.���=��)>���=�����1Ӻ}U�=������=�,��wj;��Y<S��=0�=�ct��Q����:|x�;�a�<��>%�$?�{�>�ۂ>�7P����$�(�͝�=�E�=��=�u�<�Ծ�e��F���οn�N��>�c�?�6�?@o�=�A)=�">�����ڠ�͋�?����H>;л><6
?�)7?$��?$�??�3?��=��߾���������p.?L",?��>&���ʾ_��3�=�?>Y?�;a�A���<)���¾��Խ�>�X/�.~����D�h������o����?��?-A�:�6�|x�g����\���C?� �>JZ�>��>a�)���g��#��2;>T��>hR?��>��O?�;{?"�[?�{T>R�8��+��,ҙ��5�/�!>@?}��?+�?�y?�r�>��>ެ)���%C��;�����fт��ZW=N�Y>>Y
�>�>aD�="FȽ�����?��@�=5�b>���>w��>�>q�w>���<��G?���>?举���k���Y[�����k�{?F�?W	4?�9=�����1�0-�����>�3�?��?�m(?����3�=-��/����U�&˶>H�>3%�>�h�<�-=�IM>NR�>}��>��*����[5��?��A?�aJ?l��=$ǿ�fe��ě�p��=��*��澊[��au��yW�6e��=���y�J=�����߾��)�E	��n���<Ǘ�~zB�g?``=�?�>��ֽ��~>	�=���>!y�=1������,r ������f���	7=��>�̧=��>�=��5���޾U�?�d?�;?�NH?�*�>g�>-)���=+>׫#>�I%?��ֻig��N�ž/BJ�Wݤ��ľ��Q۾}g�2wC��夾�q>=u���&>��=>y\X�t�5�ZP>�L�=���=�� >(1;; ��=鳺={�>���=��=g]�=~?�#���ä��q�[�)��X5?Ce�>�t>�,��Y9?���>>g��u���(���?��?A�?���>�������>V�ݾ�p���T<��%>H�?�Q���i6�#'�>6��>}���M������@��?4��?4fG?�7��yp׿�h>V�7>$>��R��1���\���b��~Z���!?D;��C̾�9�>��=6'߾ЕƾHd.=ˊ6>�lb=�f�2V\���=o�z���;=l=�ى>��C>n��=%3���ݶ=H�I=O��=,�O>�ܗ���7�v,���3=.��=q�b>G&>�s�>z�?_�0?�d?iº>�h�;Ͼ9������>	��= Я>�s�=k�>>jd�>��7?	D?��K?��>���=HQ�>��>��+�C�l�Z�徹@��n�<���?Au�?���>'�<��G�6���=��#����?%B2?W�?���>�U����:Y&�g�.�Ë��f�:�#+=	nr�QU�	����l���V�=3p�>���>��>�Sy>��9>o�N>��>��>�;�<�n�=�Ό����<���� ��=������<vżU��&��+�����8��;���;>�]<���;�=�^�>�>1�>f�="+���JI>h����JI�`��=V�����@�So[�)�j���%�J1E��8#>R(C>�%=�ڏ�6�?` >p҈>Ɉ�?�Y?��P>�g���ž�Г��*���r��W5>�i=��8���@�#�g�1H���ؾJ��>���>m΢> �l>��+���>��Fy=+�G^5�	 �>9|���n�g;��"q�43��C퟿�
i�.̺e�D?�E���=��}?=�I?�֏?kv�>�F��6ؾ�?0>�>��S�=���p�!����?T�&?^�>R��D��Ҿ����v�>�lV�w�K��홿6)�P�.�l��,z>�â�P[Ͼr>�! �������3�A�Z���>O�A?J��?$jl�Ov��$BT�����[U��?��x?Mo�>��?]r?0�%��4�QF��vN>�Gf?��?.��?]>(Ը=�«���>p
?7Z�?<��?�wq?��D��>�߹��>p ��2�=52>�z�=2��=��?��	?��
?�������(	�
��֒a�I�=�L�=G��>�,�>�g>�X�=f�G=\�=��[>�`�>Rߏ>�!o>Qq�>W��>�֨�����d�?�_>\��>�:?z�s>h�����|���=Ȱ<x��r�;��{s��8ݽ�j�<�����x�<���=)[�>Z1���p�?w�=>2&��C�?vZξ	�Ž��2=�}I���{��?X��=3p�>-}�>�(�>���>v�>%>�-��dH�=�������W���M��
����->�}�� ���6�{�p���$�n�Ǿ���S�e����.�7��N�=a�?$^H�c�m���ަ+�D�?�>��&?�3�������!�=��>02�>^)��3���W�����Z�?0�?c-Q>,�>��]??���;kE�<ǩl�)],��i�/�f��G��a���;l�dؾgQ���q?�6�?<j?�A�=��>.�P?S�����po}>Fk*���I�%�\>uƂ>N;��W�پ	�	�th˾��p�������?C��?E(3?پ�,p�(>ڧ:?��1?>t?�2?yA;?7���P$?��2>�?�_?�4?�.?w�
?��1>P"�=���I'.=�,���V���Rɽ��ƽ�����8=�et=[D�7�;�0=��<�<3�ǚ~;����s��<<hG=?�=8��=\,�>�TZ?+_?���=�;?pڽ�w`��A��?񱗼���bp�Br龻U���g����?�S�?֨�?	}�<��D�H;)�X>�֓>���=&�S>�o�>uB>�=u"� ��=|e>}�]>�C�3w��_Ÿ�|	��y�(:6��y>{�?3!>�_�-\�=*e���A/�>E�پ��׾I0��ˌ]���+����t�>G�:?$ ?�i�<��ž6�0>/�p��d?��(?,W?�o�?�x�=Q�ؾX���O5�G�=W'�>=�A//�p���kң�{J$��xy�q6=>�m�}&����=o6��y�����V���U��l�>�Խ�@��Q�=�+��mپ�	��,�=T>#����%�!t��[���K�??ݑ�=�c�.�x�z���Uj>�g�> А>�o
�.��>D��\����I=��+>���=������!\�C۾0��>�OD?��T?�݂?�v���5Z��(c�RD��ԾMl=�8o?V��>4�>Z�>_�W��u��������J��]����>P�>�����*�o��]؊�
��>��?nO�<_F?�%?�_�>�I�?��>�ǋ>��u>�M��\8�*+?_Ł?�*>=����ҾΈ+�ء�r�*?�:?��g�[�>h�	?�&?0QB?�2(?^��>i�C># ľN�7��b�>JƳ>��Y�"i��L�=>_!?!��>��\?�~?����H(��F��G��!
�=o\�=�7?��*?��/?���>#��>ಟ����=;��>�c?��?}o?�"�=6N?�Y0>8��>m��=G��>M��>��?w?N?,!s?ƚJ?��>:T�<-±����Öp��bP��D�;Tj<�~s=�o���q�hI�H��<���;+C���G���y��2�B�/������;i!�>p{m>�����Z>:ż��W�pw/>�A�~���Ƈ����^��O�='[�>@?�>�O�z�8=f*�>x?�>��� �%?.�?B�?�G�<#Z��%¾��0�(�>Ը>?Cb=N�o�5F���v�6�d<6�b?�@U?�V�i� ��a?J�_?+���I<�0�ɾ�j�p뾥)Q?�
?N�h�9w�>��?xKh?�?�M�=�n�0㝿��b��sY�U��=hъ>�d���_����>�:?�Y�>�b>��=��ž��q�sB���C?',�?Z�?��?�49>�Gj���ۿw���sґ���]?��>ꃤ�7� ?�Q;���о!U��V��{Z�u窾*J������ȥ��M$�f���'����=JL?ŏq?D�p?��^?`\ �onc���\�A�~���U��#����0�E�T�C���C���m��y�����j���,G=�fm���"�1F�? �>��<+��>�6ؾ�u�h;���>�W��R��/|C�-���A���"�<yJ� ;;�b?Z �>I}.>YGA?r~\�gK'��u[��EU�����=��>�t#>8�?\��=�ܽF�s����s�� \Խ��>�b?t�F?km?0��6�+���������-��6���lK>��0>{�~>�G�ŧ��)� @�=8p�/���H������{j=F�.?�[>�k�>�B�?�?���0��]����Y-�.C�<���>
%b?^��>�E�>�[������>��l?T��>��>�����b!�5�{� xʽC�>�\�>c��>�p>�-���[��V���p���"9����=��h?�p����`���>��Q?��:��H<�R�>H�s���!�I����'�nT>q?]�=y�;>vzž�6��{{��)���(??�%���P �"u>�0?J�>ַ�>-J�?���>n7����c=;�?f�Y?��G?8"2?���>࿀=J���_ǽP�?�C�=#��>R't>�Ƕ=$�=�'8���t�c�0|�<�J�=�;��޽��=?ڲ�,���|U<7KK>q޿l$K�*�Ҿ����
�h�������[���S��ġ��.���3T��������8V�=�t�����ww� a�?���?�3��.<��#5���}��|�3�>�Kx��ؚ�1ǩ�
'�߬������AҰ�ס!�I�O��<h���[�ʳ'?�����ſw��m���?�?u�y?���5%��Z4�û4>��<�;�:�f߾]����Zο�͠�?j^?y��>���y���hV�>8��>�k>mGm>�ߍ������,>=̶?�%,?8�?�e���ƿ�Թ��J=���?,�@�yA?W�(���O�X=fJ�>��	?�o?>^�0�Y�����J;�>z2�?7�?��Q=tzW��z��8e?��;�F����wn�=�W�=��=R�C.K>�-�>���IA�qyڽ��3>Od�>i� ���$^^����<3�]>�Խ���rl?�q]�:a��V�龵nG����>�))?���>,;�k�G?�yb���Ϳ4X����>{��?=��?�7?��t�=M��@Ԉ?b�4?�f�=�. ��q��2���<��V�>��h���AZ3�t��>���>"�U�"��ƽ:=�X�Cdm>п��8ſ�{!�׫���<�Ց��xl�<��TA���
>�t���#v��=���D=���=	�J>B�w>1>׬K>�iV?��h?�p�>C>J���nt��1��IE�����%�����#�V��ht �&�� 
��x�@4�M����=�p�=�Q��o��"e ��c���F�
.?�R$>��ʾ��M�8�)<�eɾ ����J�����$O̾)�1�n�x+�?PA?������V�գ�J���a��W?fS����O����0�=ơ�1>=�>a��=�?��i3�eyS�a�*?��4?	����Ɖ���=U6��ow�8�l?^�+?��9�Τ�>�\F?:�<�n�=�s>2�O�%�V>й>��>�읾��,�+�?d?���=`�=��>.�¾�ڥ�֙g>�'���K;���(�����N;>�샾���=�T��Ĩ=;U?���>J�������9�/�EUQ=��?w,?��=��Y?�7M?� >M�L���:�3����=VL?iZc?X0�=�z��� �RѲ�+*J?>�V?#<�#q�+���3��'�޾=.;?��k?���>\"w=�WN��b�� *��@?E�c?n���ڻ�i����{�G�E?�f?!�J>c-��T�L?cB]?�þ͒(�������i�hw�?$=�?,��? \">R�=7K�=��>}`	?H3F>{�9�F���񴾆�4=��?)F��Jl� x$���E���v?���?�|p��#۾�����=	����&�?X��?򼓾�3;�� �%Um�v�	�/�;�x�=��@��񦽌��_�5�O���W�
�e��<W�ʳ�>��@�.�ML�>ALJ�$,ݿRϿF
��Ӱپ��{�"�?hߒ>��ݚ��_�"�m��>�7C�䤔�o��>p�>qt�������	|��D:�i�Ѽ���>� ����x>.BH��N��>�����<�ĕ>���>�+w>~�½����~��?���U�Ϳ�t��|\�ӏY?=P�?ǀ�?�O?R	=��m���l��8�<a�E?C�p?�T?��R�ٶ6�%�j?�_��wU`���4�tHE��U>�"3?�B�>S�-�c�|=�>���>g>�#/�x�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*�^�+��<A?�2>���I�!�C0=�TҒ�¼
?V~0?{�f.�[�_?�a�G�p���-���ƽ�ۡ>�0��e\�M��>���Xe����@y����?K^�?_�?���� #�g6%?�>u����8Ǿ��<���>�(�>*N>�H_���u>����:�i	>���?�~�?Nj?���������U>�}?� �>4�q?/N.>�|?��=��4�%�J��Q>.z+>60��n"�>��Q?���>�"�>oY��\�E�k�3���J��}׾O�-�[|w>��`?n<?bۙ>9��$���>+��fB�·<��=w�i�%|=��)�[��;� >2U>��l����?�p�?�ؿj���r'��54?��>�?���c�t����g;_?�z�>*7�.,���%���=����?G�?t�?�׾@c̼�>��>sK�>>�ԽG���������7>��B?��eD���o��>���?�@�ծ?ai��D?��&�D�����D�+�0h
��l�>p�6?���6�>�?�z=�SD�����]��B�>h��?���?o��>��v?㭈�ȍX��޿=Ě>PD�?�F(?�cA���:�t}N>�l"?�X۾O~s�٬޾�?L��?D@O{f?���e�Xܑ��,��xB����=�bؽ0*E��P����<�V麝@��<�=�$�>���>�k�>w�>(��=:c�=���=�R��()�	���,c��u�6�!;��� ��!ž�v�,�[��������������ѽ�*v��`��Mž���}>�LO?ӦO?Y�p?�/�>�3<-b�=�����B=�k�!I=�m�>Vr/?8�N?�.?�������<c�=�{�=���fy����>Y�E>���>	��>_�>�c'=n5I>��A>�V�>��=S�=�M:�r<}<K>�͢>���>D�>��<>��>����
���h�2w�:�ͽR��?�Ĝ��	K�啿�ދ��鷾�E�=��.?�>�#���"п����H?����_�su*���>�1?f'W?��>���IbH��>Cy��)f�)>����]m��(�p�P>1O?��e>�pt>s�2�y�8��bO����o{|>O�5?���iL9��+u�.AH��`޾F}L>n&�>m�M�܏�u���o�pi��v=ϥ:?�?�����=�� �u�*���AXP>��\>'d=2�=��L>�Ud���ƽ�PJ�ʝ.=��=�^>59?�8>t�=ZT�>��h�B���>��Z>�MA>�7:?�?Jok����Sp������]>%��>�1�>I�>��I���=x(�>��_>�\Ƽ����%���k:���R>�/t��s�V�}�+k=G9��F��=U�=���;��x9=�~?;���㈿4뾞g���lD?�*?&�=�F<��"�����G���?`�@m�?�	�ޢV���?�@�?c
��!��=�|�>2ث>ξ�L���?\ƽ�Ǣ��	��(#�S�?��?D�/�8ʋ��l�M8>�^%?g�Ӿ8ֳ>��F������k��8G��&�<���>�G?u�	��<����>�??�{��������mBY��� ?�e�?��?2Et��L���I�[o�>-�?l/y?E1�>J����Ru�>�JF?]R?!�>mp*�3F���,?0�?�a^?dc]>�X�?]�Z?6��>�4��-�G�M����L��3�<�;�4�>�p�>\�,���U��Db�z�s��񁿪�:�\>l�z=Rw�>J��H���(er=���r�a���>y�>�但w�=��?X��>�5�>u��>:0�<�͇���P�Qc���K?���?&���n���<Ҝ=��^�C0?G4?��b�џϾ<�>ޤ\?�ǀ?9[?���>N��6������N]���x�<��K>�]�>IF�>����K>G վ�D�V͊>�ח>! ����پ���aū���>"p!?�p�>g�=�?ep*?óp>�}�>.lG��珿c�D��"�>P|�>���>��w?�g?C�ʾ$�����?c��gwc�/>S"u?�?�f>�֏��O��O���e�;o�c��G?C�]?�[=��I
?[Ј?'IN?��<?$vz>Jv0�xC�������w>��!?F2�pA���%�iV��o??���>
���v�׽�׼�C��J��$#?�%\?��%?*����`�|¾-��<�0�^V^��<T�?�x>B�>�:�����=�o>ǝ�=�8m��g4��lf<%��=eё>[_�=�7�����%?�ô����7�=Vf���@��lf>%S>�����gJ?������L�����p���q*�?;��?�?�w��٩e�\/??�g�?�&?��>W�оZ�־U��73�`c��D��N�	>�Q�>k�/��K	�&꡿����f5}��ƽ$�B?�>��>�M�2?��<�ʘ>n+���\쾿-澰��IT���5���=�6g.��׾����5�ǽ�#���Q���j��#��>ݷc<X��>�?�҆>>�>I�L>?�=l�>z|�>�l�=8�>
`^>�R2=2�W�	����&�O?�5��!~ �PE̾k��q�C?�Y?R8�>G����Hz�b&"?��?J�?.��>(�j��L*����>��>�Ԁ�r?���=�@����=����]>��M�`�9�$��=�>h��">�:�F�Y�����>�?�GO�:�þ�q�j�¾�B=���?Ml"?��(���U��Gh��VY�A_P�N���S�)æ�:��{�q���������tg�4�g3=��)?���?����龺̱�h��1��m>E�>�p�>z)�>�2>ܤ��/:�x�]��&�����2�>�{?B��>dF?��,?�yT?|�??P��>3װ>߄ �2�>�LX��L>� ?aW7?f,)?/�??S5�>��?I�m>�}>ڻ�N���g ?�@?.�?��?��>���I	�!^Ѽ���eFX��q=F,=�Տ=�d6�Я��X����=q?���O~6�<���t>i>��7?S�>@��>&U��ux��R�<|��>�[
?69�>,����r�/�+��>X��?1	���=z�0>z��=`�Q�g���d�=����=�=�1��
O�9��:q}�==��=��6������;�N�7d�{<؛�>ZC?(k>�N�=IBC��3����⹺uՎ>�>W)��a����ߋ��8���$c��ח>��?~:�?t�<.��=��=�b��n�y�۾��ľځ-<]��>��?"H?� �?�wQ?�#?��0=��*����%������t�>H+,?��>1��OIʾ�ܨ��23��,?Xl?Ӷ`�����(����rfӽ�>��.�7S~����+D��C�M���s��08�?���?w�=���5�W辍ј�������C?�	�>\�>���>�])���g�R��[=>}{�>��Q?Ga�>6�K?p�r?Q�^?��;>��+�=H��RŔ���Y���=tJ;?�h�??��?Pa|?��>���=R�<���⾿㾄�C�>��
�s� P�=rf>��>�p�>z�>��=3Ĥ����@�e����=(X>>��>�2�>�A�>�ۅ>)4����E?��>2澾���e���Ն�z):��Er?�M�?p,(?P�<V�V�E��6��"�>���?�ӫ?3t*?�@Q���=����߉�������>�޳>��>�m�=��a=eD>.�>��>ޕ�Lh�Z�<�7�e���?;D?�$�=���C�P�<a>*�ھ�'h>\�p��$�+�
`k��H�=\���6�������Ծ�ƺ��h��@�	���������@?�>L`�<SK�>�fZ>�LY��g��Z�<�>�}����=�D>.+ =�q��{����6�n�I�"�s<d9C>X�>��þ�y?eFK?6)?�NE?4��>�F	>ppX�Nޔ>T~k��2?�o\>b�U��&��QC�P|��
��?I޾s�Vz_��q���&>�5��z>��+>n�=�f�<V�=��=l�=��;]�\=s��=pj�=㭣=���=B�>ʢ>(v?����\���X�,����:�]?/��>*8�=����n?�_�>�.��u���{���Fz?'��?�K�?\�?�h��[��>~\��������=d9��f��=�g��~��=��>��>�g��m��(T8��F�?�� @BC?�v��º�G
���3>%>>��N�X�5�K�K�94e�!U�gI?�h8���˾��>vd�=�R�g�Ǿ��=1�7>YD=*����]�b�=?���FX=|O�=�b�>;�K>��=�۩�P��=8e=6��=��R>�7B������'=;��=�oY>��#>��>�?! 2?b�b?���>��Y�n�ɾS����>y�=��>�8�=��n>{��>�+?�1?I�B?���>q�<��>1��>�.��n������ƾO-�=+{�?�p�?n��>�)L=�fj��:�9'�¿۽D%?�	9?�n?龡>�U����9Y&���.�"�����4��+=�mr��QU�<���Hm�5�㽶�=�p�>���>��>7Ty>�9>��N>��>��>�6�<wp�=:ጻ���<� �����=�����<�vżH���eu&�G�+�5�����;o��;�]<x��;�E�=��>t�>MG�>��=ϗ��C�*>�Ԙ�)�I�@�=Q�z�B��d�+�~�/m/��+0�=A>_[>�2����! ?��c>0�7>D��?`�s?��>z���־=��V�[�;�H���=]�>��;��;��/b��EM���Ծ&��>��>a��>��l>S,�[?��?w=B�pY5�)��>(h������ ��q��2������li���ԤD?�@�����=�~?ʹI?�ߏ?���>_"����ؾB0>%��m=����p�Ɖ��-�?�
'?���>p���D��&�ץ���>��P�u�)�W��ӎ��{��<��_�>�Qǽ�!�Bu���5���W������y���>��_?o��?$敾�ۙ���@�X�I�%>���>p]?�R�>U�?�o?�(=��žM1>��u���l?�"�?���?�:>�=qT��Q��>�7
?�ŕ?P��?,%s?�-�ޮ�>+\^��>ڈX���=8i>�ξ=��=�1
?�D
?ǻ?�ǜ����Fm��2�gvO�H�E=�ڝ=y>�> �>p�k> ��=�.{=���=�_>���>뭐>�[>���>+˂>ꢾ����(?:�=gN�>\,?�G�>�Ge=-*���Ȁ<�?���8�:G�HG��!��T<��ּ�%=B1���>��ÿ��?b{k>�3�\"?}���1��;>wJ[>8�ƽ)��>�G>�{>2V�>p8�>G�>Zu�>l�,>��>�������A���T��Lξ�w]>�V���#���_m��)�nS���(���f�2���
QF��^�<�g�?�P ��6`�
�&���
���?�#�>\74?�Ñ������>l��>կ�>�,�H��\�����?���?�a>��>kW?�y?�V-���4�0�Z���u��A�Xwd��s`�p������S�
�����cD_?rx?<�@?C�<�y>o��?�\%�xҎ���>`/��;���)=‥>ɏ��?�^���Ҿ����+���A>c@n?9��?�t?gfX���=xa�>F?�W?H�~?��D?��?�*$��3?Ap=���=��G?j�M?��'?��H?��<�5
>��= ^�>�����(p��}5�ó�����=@�=���Ӆ�=�Yt=���<P���m��=O���Jҫ<5g�=�w�=+$H;%%�>~�Q?+C�>I@�=�R8?� l��.�����0?���;�Q��㬪��߹�����;�=[d?R\�?U8V?�>m�:�(�S�H��>Y}
>��U>e�?>5��>�睽ٵZ�K�a=+�N>��n>/V�=�O�������wɾ�^Իxq=��>Z_t>���5">�U��.���E�,>�쐾@�������v��rR�ꌾ�1�>�vP?�,?X[>@2��� �b�^��<(?��V?e�?�z?���ʐľ��/����8��ۤ>��=w����!����=�.���N>b?��A���y�Y>�����۾�Qh��L����2'�<�"��p=�
��UѾ!���@��=���=ѻȾ��"�v��󸨿(XM?���=�9��b�������*>.�>_F�>lS:��Ȁ��FB�x#���#�<M��>@7.>����b\A�����N�>��D?��f?=ׂ?�1a��c���8��Oھ(/�� ��<�>aM�><o;?�0^>b�=v���B#��_��bJ�1<�>��>'&�V
0�9	����/��}�>�T?ço>��?!-?��?ag?�<?��?�\�>���;�r���&?C�?�`�=���=@��/�B�c�*��_?WT3?'ȑ��Ҏ>��?�Q-?�l?��I?̈́?�G>��^��2�y>e�>�.V��i��_$�>?	?�l>��f?1%U?��ӽ���x�>��O�]���v>�,?�?cj?�j?���>e������=S��>�c?J-�?��o?��= ?��1>��>�J�=���>ה�>�?rFO?��s?��J?�u�>͸�<nG��T���s���M�Y��;t8J<`fy=b��nt��y�=�<��;��j���v�jYE�L%�����;Il�>�_�>}*��Uu0>P¾�`��?=1>�-�;�����ِ�,�8���=|�>l�?�>A�����=�>�j�>��sF&?�.?m�?�O�<�]a���߾��S�!G�>��B?F��=�Nh�`k���Ex��r�=��o?9�[?�t^������a?��]?��lT<�> žJa�mY��DN?��?��B��`�>,M?�p?��>�Ei�?�m����]b���b��@�=�q�>x^�C8d�F��>J�7?z�>�V_>�Q�=dc۾�w�qy����?몌?�k�?o��?#�+>a�n��d߿f.����,^?+�>���(p"?*��2оX���(9����ᾩ���ؕ���(��������%��V��+�ٽ���=��?��r?q?[�_?�o ���c�x3^�?��oV�Z������E���D�"\C��n��\� ��7���C=�.V�v2�C��?A��>�t�=+0�>^o�����0��\�5>�@���)_��<=�˽�O�w�ѼC������V\����
?�U�>k	�>�FZ?�9i��M���/�(L#���コ>���>x��>�k�>�j���X>����ҍӾ�{|���)>~p>��\?rr=?�o?x���J�2h�as���%����XA>Z4�=R��>�%��cIS�-/��L����\��si�r�ؾ,rG>X~?�k�>�(&>��t?w��>�0�o6���,�����!-�=�~>S�Q?��>��d>[�)�jF'�}Ų>��h?�Mh>��>f?����׾��}���@�a�?���>	jO?��>�vr�}\��W��ۍO�YZN�c�z?{!M�]CT��YV>֛)?==�=MC>���>[��ՍN�I���������*��>_��=���=k%��|ݾ<�x��F���6(?4�?����{�(�l�>6�?���><�>v�?sՍ>d¾�1�;ē?�%\?4eK?��A?���>!�%=D���\ZϽ\A)��yJ=x;�>�k>}Fy=Z�=Q!��S�2�Q:I=	_�=���\ɽ.�<�D��`WN<�$�<�v&>��ۿ��I�$Ӿg�����b��>����ƽg�ʣ�������v�G��B;���\���i�������l����?e��?����1ˋ�eh��f[}������'�>qm�΀������=��K�߾����� �2�M���g�d f�=�'?�����ǿ�����:ܾ! ?�A ?#�y?��7�"���8�ͭ >�@�<�.����뾦�����ο7�����^?���>���/��\��>���>��X>Iq>d���螾�2�<��?"�-?��>�r��ɿO����Ĥ<���?-�@��C?�LC���M���>7�?���>����A�7��-��?o��?g+�?3�B�� [�G�=���l?���>8�?�\�C=΋_�+b<?�->6&}��h>Ψq>��"\ὰR��Ο�>�>��>=�?���7��<� �>���)`�e��?�'K�U$i�ү	�k�t��o�>��X?��>BҢ�φL?%�e���Ŀ��/�0l?��@;��?n�9?5���>M* �,I�?r�>�k}=����\���m���H<ND���5�-}{�z�_�	m>��w>�0j=z0$�.q�B��=H:�}���3Ŀn� ��0 ��:=�|ﻔj���r����Ž�����o��Tj��޽"�Q=9��=�%8>�<x>+{K>�p>WmU?%�j?\8�>�F>E������T̾0�����|�
��C������������eᾗT	�N���������6$?���=leO�_���Hj�t�`��F�[�'?��>�,˾D�L���2�_�Ҿ�����Լ�B½âϾ
!2��Bm�2�?�B?����h�Z�AO��{���"���W?���d���ڱ��`�=��"�� �<��>p}�=>e۾|�*���N�L�&?�p1?�K����D�|8T>�p��Sq"��Q?� ?�П�W�>�)9?����5�#:~�>A�>�Ĭ>��>��>�=��G+�7:!?K|M?���)l�%��>����'q� �#>_VA>K������@>�̲�������<G���sH��v�V?�>(�)���B��,W&��!3=�x?�.?tG�>p�k?�PC?�ɞ<n���^S�H��t=�W?(i?��>��|�HIо����X6?ge?�$K>�zf�{(龐d/���\?dPn?uQ?FY���|������"6?�&�?	K�������`����ܾn!?�7N?��
?�7M���6?~�s?����Pl>�Qg���`�8ː?<@ir�?��D�Τx=B=�?�Ȳ>L<���L�mQ��x��^t<�ʂ>�7��S�{���G������.�>�?j�?3���g���=K��ƫ?���?����#�<�����m����(K=���=� μ�V*����2v:��Ǿ���{���N弸��>/@���!� ?�<��9��?ʿ�x|��Һ�އ(�j�?	��>���m(�� �h�lk���@�uG�r�G����>�><B���j���{���;�w��۳�>�*��Q��>N�S�����՚��L�<�R�>�B�>��>3b�����M��?�����fο����?
��hW?�b�?a�?
�?T2�<��p�y������NG?�r?A�Z?i'��lU�d��%�j?�_���U`��4�|HE��U>�"3?�B�>\�-�d�|=>���>Qg>�#/�v�Ŀ�ٶ����b��?ډ�?�o����>k��?}s+?�i�8���[����*���+��<A?�2>���D�!�40=�YҒ�ü
?a~0?${�f.���_?��a���p���-�W�ƽ��>��0��h\�����v���We����@y���?^�? �?ή�y�"�A6%?��>=���#9Ǿ��<%~�>�$�>y!N><4_���u>y�W�:�[d	>���?b~�?m?��������KZ>s�}?" �>�ހ?���=,�?zy�=�
�������Ѐ=��<�X����>��*?�F�>go>�^���"B�TP��m�F����'�$.�>�sh?�y_?��9>�nL��C������罅m۽�Ⓗ(���4T�����n>uG�=��=k� ��˾S#?�y�Y�ؿ�I��PQ,�=�4?L�>��?���s�n��k��(_?'��>[��$��UƋ�}���D�?W�?@�?'�پ-�ܼ��>ԯ�>\��>��ֽ��������7>E[C?0��Ʉ���1n�g��>�n�?��@�{�?!�h��?\�� �����w4�'a����>�/C?��U��>Z��>��C:�"b�>���+[�dQ�>>�?Z*�?�g�>C`�?�/���L�h�3>��>&ӊ?�?�{-<'%��B�>FL?#�L���'��3� ?�l�? @��?qۢ���ݿ0��(����Ͱ��8>XN�=k^`='´��-�=�fN�s���ְ��N�<�2L>�k>}x*>sa>�hR>��b>����"�y��ɖ��4�	����v"�@U���O��;���Ͼ�#޾&)K����x�Z�Q3��x�D�hqa���=��T?_�V?@�q?"�>�/ֽ��=�)�7�=۹B��30=�w>�F??��K?A�!?Q��<�;��3qg�FC�ܕ�F�p�w6�>IiV>z��>9��>)ѥ>�3=7E>J@<>�W>�!�=���:�	��5-=i>���>��>�>�<<>}�>�ϴ�c3����h�w�N̽$��?؀��ɻJ�+2���<��N����V�=�_.?�v>3��'=п=����3H? ���r*��+��>ֽ0?�fW?
�>�����T��0>���:�j�>Y>�! �Osl�ߊ)�P/Q>go?��i>j?r>��1�/+9�a�J��ε�E�q>iw.?�Z���$C��u��+L� P�Z�5>��>�)����DG���~�]j���N=r�=?7��>�������b����Z>n�N>�N`=#^�=�wT>I�9��n佢�F���<Ќ�=.<J>�.?O�,>^�=�+�>����;R����>v�?>��+>�>? a$?���̀��c��ڪ,��Xv>� �>M`>�:>�;J��ܬ=M��>��a>rF��i��4�	�6.A���V>�F����]��&y���{=YC��P��=�ǒ=p���;�!�=�~?���(䈿��e���lD?S+?b �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��L��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>�R���������x�^B=���>��H?�����	���8�=P	?��?�,��������ƿ{�p��W�>r��?�A�?Y`r��l���>;����>&��? Y?|_>��޾� K��)�>�D?v9V?��>q��'��?)	�?概?�7Q>?��?��M?���>۳н�(�؎��?��#sl>���=_��>
�d>4r��f�����8��+t�t�&���>�=8;��>�⠽a꾄�\=���<�艾QY��\��>x�J>�,K>��>�
?��>X��>���=��̽�E��p����K?:ӏ?�p���l�,~�<뢍=�d��t?3�4?;���Ukξt��>I�\?p��?s[?\�>i���f���������{��<^I>���>9��>���hkD>��־�O?�e،>�0�>d����ھ"���qnߺ��>Ũ ?O�>���=�?od+?TzZ>� ?H'Y��[���K�y�h>,>?m�H?[�?z�)?:�׾�0��/��6&����H���P='h�?8�>��>a��� 6���S�T�м�G@���j?W��?�eR�[�.?��?Ӿ�>�Z?x�>�㍾oV������eB�>�� ?]��ԝ<�P5'�<����?_	?���>#B��67����g��������?�\?��&?���R_]���˾�F�<�y��7�/<54�;>_-���$>��*>ꑌ�I�=�>F��=;ub��7>����<���=���>+;�=�}3�%��W�)?��;�˨�%6�<�Qe��>?���J>�j�=��ᾤO@?)���U��/?��H9��wҼE�?��?�~�?h(ǽ�,b��z3?D�?X��>{G?&�ѾǴ�6�Ѿ1�c����|־���=2��>�,���n ��ڥ��T���E<�yq��<�>���>B�>�4M?،�'�>�p	��ʾ3_���$�c,^���]'����>~Ⱦ�`��`���SQ����������l�>(���=	�>���>[5>�4:>�H�>��=\>*�>�n�>�q�>WZѼ���½��#<V�9��=R?�ۿ��'�%I�׾����A?�c?�l�>ke�$���/����?�}�?^|�?��v>|h���*�pa?�M�>���Me
?�8=`5���<
���GW�呇�Q�b�>� ׽�G9���L��`h�|
?�l? X����̾�ֽI����f�=��?��%?&	��7H��k�i�[��LP�:&v=�2?��{���{�uVn������z������_&�ͮ<L�(?{*�?D%�>Oy��x��q��*��l�>��?]I�>V��>S��=�)�&���Q������F����>XO�?�}>��P?�p6?�TK?�G?j��=�5.>dN�<��	?p�����>3�?�?ޖ>?&.?��>�V?�C>tuӽ	����ɾ�`?|j�>?SW?	�?'���U��:����(�'����<7�>��s=�B}�.H���z�=:�=>I?��2�8�2<��E>h>�7?�:�>��>P֍�0����=�5�>�
?@*�>�d ��ir�������>_ɂ?�_��3=џ)>���=c\��x��9���=BDм��=�����w;��|<���=��=ç2���:�;��;H�<�o�>U�?p��>p'�>q��z� �����=vY>��R>1�>]Pپ�|���!����g�VTy>pq�?�r�?p6e=���=O��=ne��XP��M���������<�?�K#?�ST?g��?��=?#n#?D�>�:�FO���]�����ʟ?x,?ƣ�>-��~>ʾ6ܨ�Nn3���?j6?�;a�5���#)��¾��ԽZ4>�o/��9~� ���8D��>��h���;��p��?�ʝ?�bA���6��h辵����c��f�C?-��>��>z��>;�)�ϻg��.�6�:>��>��Q?Pw�>�N?�}?�vT?�M>�6�[���\��`X�<d+�=�/?6z?���?�v?�
�>���=5d_�20�W ���O��ƨT�)��=�F>�'i>��>��>R'?=$+��r�㽯�V��~�=/�>|��>���>�,�>��T>D6���G?��>P(��\y��𤾒��9�<���u?��?�3+?v�=�n�0�E�~���Q}�>bU�?�۫?q*?v�S�LU�=�~ռ뜶�r�!��>���><�>G.�=��F=�>���>,�>�4�LR��T8���M���?�F?K�=�տ��W��r�����\���}Ѿ<���|X��B��";��N{�Q���9��4�P�x1��о��澇����ͷ�_?9ZS>��>��=�����/��[�,l5��/���=�0�<~9=1�<=�K��d-�*�9����w�I-ؽ�rȾ�}?H�I?k�+?�fD?3s>�{>�;ݼ�M�>�&��s�?/�_>��S�����[1��������G	վ��־��e��%���
>+}T��s>��:>���=;́<P��=B�m=L|=��ʺ?P3=�=a�=tK�=��=�>��>o��?x~���Δ��L(�_�L�$%�?l�?�V������g?��X>�l��l����<�E�F?��@���?Z?P��=U'�>�\-�}��=)U>�g@�CT�>BN�=�e��QX�>��>B�,�#�v�q�=�#�?H	@)(9?ș��轿��T>�*<> O>�\O��3��I��rs��x[��s?@�6�hVо,�v>oh=>���o;Rf=��@>�a=���~\�7�=� ���Q�=�I=es�>!�:>�(�=n
Ͻ&��=<�=̶>d�H>�0�;�輦�_�I�;=1ޑ=�ab>KF>m�>V?]L2?��h?��>>傾˰Ѿ����|"�>N�=���>J=f�p>���>�4?L�??�D?<�>�=�<���>���>Cb3�[?g��s �v<���w:=�?���?� �>lG*=�Y��#��1�Ǥ���K?�l9?��
?�?�>Ⱦ�Eֿf#��u>�7d=h(�=V�?�$9��=ѽ����K��S&��j�=-�f>�٘>�~>�}�=�b�=�È>*C�>J>j�,=�$"=e��=��<��߽Ɔ'�����q������F�q=?۷=&F=�j��'���=�J�Z��=��=7��>�_>�D�>���=�����;->�����nH��7�=믾kE�Zae�i7~��(��(��/D>uZT>cp�����+��>��l>G�3>��?]n?�:>�c���ƾ��$N��ZH���=LR>�]�G�<�g�a���K�nw׾���>9��>y��>�	m>i,��?��Bw=�⾻\5�d��>�f����i&�^q��=��Q���ki���ҘD?�=��a��=�"~?�I?Qۏ?Op�>W�ԃؾ�20>D��s2=��%q��֓��?�'?M��> 쾱�D��g�e"�x��(�&��|'�&�����̾��ڽ�V��a�>�	��h��p]�!{��Fm�ۯ2�Y����u>��(?�?�����?F�df%�a	��^?oы?�>Y?�C�>/0�j˿�Q�Ǿ'`+>NCf?8P�?�^�?�	�>b��=D5��܍�>�	?ȼ�?q��?�Gs?�?����>zb;� >s���ĕ�=�>���=6w�=J;?�l
?��
?F��� �	�U�����Yc]��}�<Vr�=�T�>!p�>�r>���=r�h=�=�\>X��>��>�	e>r�>d*�>��j��6�'?���=�f�>��/?��>��0=r���*g�<�Fn��!@�i�-����s�彅Ӵ<-��>M=p4���>k�ſ7��?+�S>.C���?S��a�.�@�F>�\[>m�ӽ(��>A�A>f�}>�/�>{9�>�>έ�>�[+>��־�R>�g�O#���@��QQ�3�Ѿ�{m>�����)��	��{��U��@��è�/�i�߁��
=��Շ<x�?eX��p�<�,�Y���z?��>[�6?mϋ��h����>���>��>����ғ�e��anܾ�s�?�]�?%Ac>}�>��W?އ?�O1��.3��eZ���u��A��	e���`��⍿͜��<�
��ؿ�1�_?c�x?wqA?�<}"z>���?#�%�-я�|=�>�/��;��;=)/�>�&����`���Ӿt�þ!��E>�o?��?�P?�uV�%����S�>+|k?�=!??�J?�A�>��>�/A?G���,bE>4�P?�6/?*wR?��??�	-����<�)2=vے=�1��N���������xɚ<� >,:�<�.�O}>P��<)���L9��N�L���a�<c|��� ��S;��=� �>�pV?���>)�i>0�9?�1��n0��t��,�*?d��<����岛��l�������>V�h?���?wWT?̚4>�HC��(M��?>�_�>��;>�'\>vj�>J�)j;��h=��>W�>�=�!��������fP��-��<�R >�;�>&>N>�yk��H=�K4�:����b�>a����K���b���K\���H�����ɰh>6�L?�|?Tc�=���{�m��R�;?L@?�x'?]I�?���<W��It/�Ϥ	�z�I�K�>~�=P��oÓ�=���(Z��#̽,��=(4˾����u�a>}�0H޾�qn�k7J���群SL=�4��TW=nQ���վ�#~� !�=&	>z����� ���$���@J?��h=iv��$�U�֨��s�>��>o�>Z�?��t��X@�[ì�Gt�=�_�>��;>r��Jo��gG�/ ��,�>�L??�U?�(�?�#��`�v�p�E�T0��tk����=b�?	�?�?�,�>ڨ
�#e�����9�W�����E�>C�>}ܾ��
�T����D���)���g=$�F?�#?�|�>/�V?���>���?�g?*E%?���>�#4ھ��?+��?&�:=��-�Jd"�rI+�B�X�Lu�>l�2?�/���Is>hP!?l� ?��9?��5?��?�kF>6�'���]�K��>�v�>(WL��������>�aD?��>�aT?-f?�Xv=ô-�Y�ھAQ��P��'>]�?�4?�?�M�>?��P���"�I)�>��U?EI�?�Y?�ڳ>���>�Я�O.�>DF�=��Q>�?H$?�}b?7I�?}JO?N��>���<�N�#��/O/���<|�=�Qn�z��<@���b��<���=��=�=�@㽷F���Ŋ��_;���=Aj��A��>%pr>�j��h->>�þ>ň��E@>j����Y�����̀;��r�=h�~>�|?��>��"�"�=�D�>�4�>a����(?��?�?T��:b�a�Ɖ۾ȦL���>g�A?g��=��l�����p�u��k=�m?�^?��X�������b?��]?AE��<���þ[c�����O?b�
?'�G�;�>D?"�q?���>,f�!n�\	��VOb���j��Ҷ=gs�>�T�Z�d��I�>*�7?��>d�b>^�=y�۾˺w�I[��c?���?��?���?z�*>&�n�19࿁��"�����^?ʟ�>@����!?��%���;�z���ی�-\����웫�Z���G��w�#�^_����ν���=�*?BLs?q�o?Sya?�x �Pkb�B^�����T������ �E���B��	C���l�^#�D�D��^�*=�KV�&���R�?_^�>�}=|��><�ԾIk���@ξ�'�>6IS���)�2$q;Eq���^����=�p��E�.�����>��?�G7>�}?��W�+�S�3��6�#���ˎ�>�|�>0e>�Y�>�I;���L�Xˇ�����&�W.v>��c?�3K?�n?r���� 1�V{��A�!�0<-�%���t~B>��>ਈ>c�U�����%�b�=�зr�s&��:��(p	��ȁ=�d2?yՀ>�>I�?�Y?4 	�&M��W�w�(1����<���>4uh?�t�>���>y�н�3 ����>6�l?��>�٢>�S��j!� }{�Żͽ���>�(�>��>t>��(�gf[��R��Z	��t8�#��=��g?����ZZ��9�>�R?����[0;��>���U����v(��e>��?��=�7>`�þ���}o|�Uǆ��4?��?[dȾ����%>��$?@�?sS�>2i?m��=T%���Q�6 �>�7r?��T?��Q?۹?a+�=����mν8漽��;�π>.��>�a�=�C>��k�![�HV�����<k�7>dȓ��2�ȑ�|+=T��=�M�=~>Erۿ`8K�ogپ~�����N
�3숾�ⲽ 9��%��E���>��Dx������'��OV��Zc�������l��{�?R+�?d��k���Z���.�������F��>�yq�¤~�p���9��������Ԭ��Y!���O��i��e�~�/?��"�fԿ<^������'UZ?6�Q?qRJ?�aL��oܾ�&��a���Q�F���=l������?(ƿqz�d�B?���>� ����� ��>���>t��>kp> ̄���ݽw>��a�=��?+8?K�K�8Gʿ}K����=>c�?��@eSA?�(�d&��Z=<�>+
?��@>��-�z�����p��>�)�?��?�*M=�W�� �/�e?P}G<��F��:����=Tn�=�s=f���K>\>�% �d>���ֽ��6>8ۇ>�"�����B`��;�<�sW>PpֽA施Մ?n5\�
Df�VE/��e����>��T?���>���=�A,?0�G��iϿc{\�dua?2	�?�|�?D�(?����X��>�Xܾ^M?ڛ5?��>i�%���s�%�=2`ؼ�P����侬6V���=���>�>�+-��t���M��a����=���ƿ��$��z��M=!���[��o��~��V�T��=���Wo��n�\�g=�Y�=�fQ>�X�>�"W>�Z>�aW?��k?�O�>i�>CX�ʅ���ξ95�>=��+������� ۣ�!W��߾�|	�+�����P�ɾ�͇��ȇ=��B�������YY�NF�֫K?q�>����i����R<Ox����Ҿ~�D����;"�'�4'\���u?��D?�v�ɢF�-���W��G�E��*?�S�h�"�$2�����=���,��a��>���=A���+���6���!?h�)?����1���o�>�ͻ;X�I��D,?d��>I}l��ŷ>�\?�]��4=,�>�K&>�?4�>+��S�����P�t�9?�J?�Ҁ�{xs�	�`>�W��ᨾO�>/�G>�W�=���=@)=P�$<���6���m��=)��=�#W?�{�>2�)�}��S`��Qa�)�>=�x?lp?��>Xsk?��B?^G�<���%�S����x=��W?Ei?D�>�H����ϾN���+�5?�e?#O>D�g��龎�.��Q�!'?�n?�Q?����h`}������zY6?��v?�r^�vs�����<�V�k=�>�[�>���>��9��k�>�>?�#��G������tY4�$Þ?��@���?}�;<( �L��=�;?g\�>��O��>ƾ{������@�q=�"�>����vev����R,�_�8?֠�?���>�������y�=u/���ë?���?@m����Z<��(	k�?i���n�<���=��	��������7��ƾ)&
��{���-Ѽ�>��@xw뽔��>JA��⿸�Ϳ����|<;��m���?e�>9v��JО���j�kkt���F���H������җ>���N���^Tc��ۘ���*���r>�e�>�D����>ʭ �G��
=�I�G�>>��>��|>6R-������?��5�A��G2��z�+�D��?��?P��?���`�;y�=h�����<�T?xO�?U�D?�Ђ�o
���S��E`?4�cz��!��Q��z�>�!7?TjV>�2>���>���=�la>	?��@�+������_�����?!��?��ż??2�?<v?����m�������m(����>�@?�82>�]�;��7�b�|��.��i#>w�<?����7\���_?�a��p���-���ƽ�ߡ>\�0�a\���������Se����gAy���?�]�?u�?	����"�25%?��>�����9ǾL�<r��>�+�>S*N>O_���u>��
�:�od	>4��?i}�?�g?͔��	����]>��}?���>b�?B{>�?7�>Z0��ï��ՠ=_}�=�?��?�=M?t�>@��=�|�0�n=�T:H�C�s�9�y_�>�4a?��N?U�L>��޽Ѕ���l+�XΡ�Z�8��;6���#���<�����g>(FI>�>�~�L8����?Op�7�ؿ j��p'��54?4��>�?��|�t�����;_?Uz�>�6� ,���%���B�_��?�G�?;�?��׾1R̼�>5�>�I�>d�Խ����W�����7>+�B?C��D��v�o�r�>���?�@�ծ?bi�	?< ��O���b~���7�O��=�7?�0��z>���>�!�=�ov�_���*�s�㸶>�A�?Q{�?���>$�l?�o���B���1=�K�>Μk?�r?gho���\�B>δ?>������cK�)f?��
@7u@1�^?��� ׿;����(��s�Ծ!��=&�=ˢ�=�=��k>�k<����`�<�>
�e>�^a=D��=ɢ6>�- >��>s��B�������㚿�gJ�L�+��}�Dʃ��¸�i5���>�9m����� :��ny���b�����`Zr�oY��\� >-"\?5�E?��f?��?!����KP=���9ڜ=4�^�O~ =��> ?�PH?��!?sX�=�����ag��$��Ő����q��l�>��&>�]�>�d�>�:�>���<��P>H�>�q>�N�=��<�챼CL@=.>v��>��>�0�>��F>\a�=�u���꯿6�p�T1Q�����#�?�i��Y�6�[l���)��i=��.ׇ=��:?^&>پ���<Ͽ@���H?�.��݁��d�8!>�8?f;R?�u>4���P V�f�U>�@4�������/>����Dx;�9�5�z�T>��?��f>�v>��3��G8��[P�KC���({>�6?�*���x:�:}u��sH�C�ݾ0�M>e־>K�F����� �bVi��Vx=b[:?=�?}���尾�u�(��_�Q>�G]>��=~ʪ=QXM>Q.b��'Ž$~H�},=��=�j_>��?�a->\%�= '�>����G�ٺ�>"�D>$> �=?�$?
�ɼ�Z��j8��x+-�l"s>��>>�=>��H��"�=�;�>C�p>M�!�i'������I�cX>N$\���Y��O��i�=����_�=o��=}>��mA�m=�}?�ۧ�.x����leѽ��O?{?��=o��Xo�v	��*dо��?��	@�L�?*P���Y�o�"?�F�?�\��A�>���>�A�>��ξخT���>�콏񖾽���"�J��_�?GD�?+橽ㅏ�:c���>K�?�t��ao�>u��O]��C����u���$=~��>�1H?i���O���=�?a
?B?�K�����9�ȿ�~v����>'�?�?0�m�s9���@��v�>��?�[Y?�Yi>�W۾>Z�)k�>��@?2R?��>rE��z'�o�?�ڶ?���?��H>Q0�?rs?��>-x��0/� ����6��hs=��<��>p>m��2\E�.��Ɉ�ӈi����N`>�*=5��>��ཋj��у�=͎�����lz�h5�>�[n> �E>���>4Z?>?�>>��>=����֫���(���2K?s܏?�%�YPl����<s�=Jh�(?T�4?�孼�$о٩>��Y?դ�?�Y?�Z�>m����%?������y��<��I>���>�,�>�$��9�M>��о�D�,��>>�>���0[۾�9��]zD�(̙>t�?�Y�>�ݲ=$�?��#?y�l>]�>g�D�V\�E�¹�>�4�>�?G~?�?����B�2������b����Z�Z�N>��w?-�?C��>󭎿N웿ꟓ��}m�&.��gt�?��g?����?{��?-�??�rC?�b>
F�0�׾�ѽ�r��>P�#? Ҿ)�c��#�����Hv#?�3?���>�o�����=���>9�X�?3�>?�]�?pO9?~x*���_��ؾ��=?���U  �V!>E��=��[>ۦ�=@c���?�=h�I; b�=*������1 >����VZ�=��w=�n<��ͽQ<,?�B��܃��]�=��r��2D���>F�L>���f^?��<���{�o���qa����T�`�?���?Gt�?�����h�"	=?'�?��?�-�>N����n޾k����v��w��A���>��>cMq� )�񚤿�����5��Dƽi��4t�>.��>~G�>�l(?Bb�=F"�>O���ʃ��c��ʻ��:�z�C�/ZF���4��:�泾���:VH�=c���{پ��>� ��C��>Z�>!��=�E�>���>�m ��R�>'��>��>��>y�=��x>&��o#�)�OR?n}���&(�ܢ��Ѱ���B?��d?	��>��o��W�����^�?r��?�]�?pEu>rIh��L+�%�?k��>J��S�
?�o<=O�Yf�<�(��;��T��Ҷ���>��ڽ��9�#L��]g��	??�����7̾=tҽ&1���wp=��?��(?�(��eQ��>o�XW�lR��=��o�e�VП��,#���p�|���ú��t����d'���"=�`*?[��?C!�d�����ʮk�m�<��e>O:�>]<�>W�>j�K>s���/���]��'�9�����>c1{?;ڍ>ǭF?�(0?$XO?FL?VQ�>�M�>L���~��>�G����>f��>�	?�T ?� 2?g�>��'?�K�>�"����[�ʾ�!?$� ?1�?���>�g?m��7����=��<xq �f�<p3<<�f��ð'�0�4�i9�<HGe>
?���7�����2	m>l7?(E�>-�>b��䀾���<z��>;�	?���>& �E1r�̑�b �>��?���	=�	+>7\�=[����ց8���=�˼���=e�a��!B�EM$<o+�=ӵ�=��R��;7�?;��;Rت<'��>x�?Eԋ>�ʉ>����U��+��D��=eS>�/Z>��>�վ�N�������Yg��Bv>$5�?�{�?��V=���=a=�=P���۠���B
��¾�a=�:?��"?�rS?>��?NB>?:$?5.>���Β���������\�?�$,?�Q�>9
���ʾ�먿�X3�֭?O?�Fa�#���3)�:�¾��ӽ"�>�e/��!~�e����C�-sn�@��2䘽��?���?ȫA��6�)��q����;��'�C?���>��>�R�>��)���g�>��H;>Tb�>�R?�'�>־d?$�c?5]g?Y�P>A�4�>{���k��@�h>��<U��>�C�?<�`?K�?��>�!�>ұ�<�F:�h�+��a���[�<��Q�b~���|L>q��>�	M> ��>!�>8Ж��)�����1�<])c>��>��>�"?�,#>�)O�!M?���>��۾��������C��t�<J/�?�?�?�O?�=qT�U�<��<��b��>?�?r��?�=(?��9����=�r:����([�H�>�0�>�>E��=�~=�h�=�Ǿ>b�>a������t1��W �?�?��??��=}Sſ#H�{%*>~H��E��;�*��`)�������=^q�=��
�?彄���߾�������	��v����?��[�c>�Q>Tq�<��J�\r> ���a�Ŝ�>}�\=$"�]+>�y�ά�/�'>zc<���*F�=b����'}?޿=?G?��G?��z>��=,�A����>4����s?�]>����6���Gv"�����;}|����df��X�Y�[N���T�=�Ƽ)p�=��>�>w�=���=� �=w��=�x��_=���=5D�=��<���=`W >�V->r(w?��>����;Q��&���:?���>��=��ƾg:@?�?>Z@��^z���W�X?%��?� �?�?}qi�Z��>�4���b��H��=����w�2>���=�3�#=�>�J>E/��N��ٴ�Q4�?}@I�??@��Ͽ��.>[�;>��&>l�M�M.��6��V�.�u��2?��-�jV޾/H�>E7�=���{���&Y>=�6>���=��2�$&a�!��=�E����3=uJ=RĆ>�e@>Vh�=������=}*`=q��=�T;>k�Z�e�#�������w<���=�Pu>��9>Z��>��!?(E@?,Wx?��>���g��.�޾��>+\j=���>sH
>��>��>!lD?B�U?��\?��>�R�<\��>�q>y�?�jIS�)Q�������!>`D�?CeW?�λ>�	)>���כ�Gx)�i���>�?��.?h�(?���>�U����9Y&���.�%�����4��+=�mr��QU�M���Im�2�㽲�=�p�>���>��>8Ty>�9>��N>��>��>�6�<{p�=#ጻ���<� �����=$�����<�vż�����u&�=�+�7�����;[��;=�]<d��;_G�=z��>��>>��>΂�= �����C>�P��
�I�3E�=�e��Z�?�qLf�9c���*�	m�؍,>�4x>3w�f����N�>z̀>W�>��?Gj?$}�=������Ѿ_���F�q���J��\=��(>��J� +���X���N����ŷ�>Y�>.�t>�->�'���-��e>��I.%���?��k��G���<^����쓿���Y�	8>�n?�ր��e]>F%�?K�?$�?�@�>�c(�`K�H�>�^��)����3�Ӿ�����D?N�?�Q�>b?��y�`����4�	�}�>K��R�H��\��1W��p��򥾕��>zų��Bվ�2��Ɖ�����>��A�>�	I?~��?u����}�a\���"�XO'��q?��n?�\0>�?��?|i���Ͼb����>�*X?p��?.�?��>�8�=�����>2/�>�ț?kB�?��\?���W��>|;�hc3>��<��="B>��=x%x=Hj?3^?n	�>�?���M�u�Ӿ�����Lc�@�=�/`<V!p> K~>�_>r�<b��=s&�=��_>qW�>���>H2I>#�>dHb>��C��[+?�½�v�>��?�hj>@U�=أ��t�G�I���y���T��0��h�$��?��Ņ��>�	R= ��>s���?:��=6���?����E�<`�>�ڂ>�
��~�>�*H>5�>e��>�<�>��=�i�>C;>�mӾ�>.��/I!�LC��R�TqѾ��y>O���l%��������]�H�����T|�� j�*���$=�A�<D�?Ҍ��8�k���)�0�����?���>l,6?�-��u퇽ķ>c��>z�>f%���p��[�������?���?�1c>��>�W?��?�i1�3�PqZ���u�J$A���d�ι`��ڍ� �����
��*����_?!�x?�xA?KW�<:0z>Ť�?n�%�Ϯ����>�/��*;�7�;=Y+�>����`�O�Ӿ��þu9�WQF>@�o?�#�?�L?wV�߅O�=/'>��;?$�'?=Cv?��6?&�.?9<��{,??T�=[8�>n�?<�)?)�0?io?�L*>�\>V=���<Iǃ�Е����ы��s뾼��<�Xx=�Z1:<$=G�:=>=�;����s_��#7=Ȓ�`ƕ<2=P;�=&>�4�>�_?;�>�_�>��9?gu���7�Cە�ǲ+?C
��/g��	p�P����Ѿ�>�a?���?��H?�>y`H��
M���6>���>"�&>�<W>�3�>��c�H��&�=�h&>�
>��=����rd�x\��8�����=o�1> ��>{|>#���5�'>�J����y���d>�KQ������]T��G���1���v�؃�>n�K?d�? ��=S�^����.f��)?tV<?�LM?!�?#��=|�۾��9���J����n�>BW�<��������
��|�:���j:Z�s>�	���P����W>.��rپ��_��FK�4�}��/#���<	w
��{Ͼ9�n��U�=�� >�󶾼:#��L���S���G?F�=�?���T�̤���>>
�>'Ш>٫���ٽ�%5�9���(��=���>K�%>���� ��AC�����]�>�#O?�wV?֙�?�^X�4d��3�����>���,?��>�"�>6��>�T����Ǿ��þ�k��~~�"��>�t�>2����=�쳾	��6$���>�?�>��+?�R?D�>�SL?�h?w{?>�5ֽ�Ǿh"?l�?;�=�S��)S��*�Z�C�!�?�K2?xeE����>�F?�-�>?�(?�)\?��?[>���ȯD����>u��>�,M��$����[>�i:?x�>��e?��?�(0>6�5����n�>��A=h�J>��7?P�?|�?bs�>���>�u�� �>;��>�_?�؅?�GC?�#>y��>��>�o�>��μ��;>n�?�)?�p9?��v?~?�>$�;�G��'.=NC�U	���=л�:9�9=oҌ�*�n�t��EC0��W�<�99��h�Ԕ۽�=M�>�[l�y��>�t>�����6>ޮ��ֳ����:>��������找�D7�W��=�`�>�a?�]�>�NӉ=�$�>�Ƽ>�3�B0(?`
?7?i���`���۾�MS����>��??{�=N�n��Ò�̌u�AW=~<j?�e\?)�c�D.��Ƞb?��]?�C��V=��¾�a����%O?��
?(AG�+P�>�	?��q?��>g�f�m�m�����a���j����=�֛>��kd����>�7?�>�>�c>��=�/ܾ�w������?-Ԍ?l2�?��?��*>5�n��	�24߾V���zU?-}?��_��>��=�z�U��wJT��ؾ�ﰾ9�]����]ŧ�u
E�����
��i=�5?��[?�Be?9�V?�b��qOY�8h+��jr�SiN��������H�l�@�9NN��s�7'���!����,=�^���B�?AT#?ɢ�����>D'��J:����f >�8��,畽G�E>�ҽ�̼�f�<W!��s������>�5�>璘>�K?77\��?�+p����?����o�>�>�>2@�=1�?D����`�@���ԁ�uؾK�S=�x>�<n?R�7?�NU?��������u�����	��&޾��>z��>e�Y>n���,�x�!�.f[��Uk���Z'v� ���4��H�"??�>%��>%��?k�?#���W�����Z��>[�=!��>�fM?\��>��>g���b"��H�>�f?[�>�:�>6��lc��z�:1ڽ���>♷>NW�>��k>6%
��X�]�����,�<�֙�=��a?����"Q�Z�>�8X?�p��*l;'(�>;I�������������=y"�>���=��.>سʾn�E{�"-��A�?���>�
��
�-����>��%?:�>�P�>V?;��=��}�=Ȅ�>�{S?�-O?�
G?"��>�E���=�s;����A�e�5=�'�>S�?>���=u�:=_,���j���3��&<`-"=?��Uڞ��X�C����=���=7$>��Կ��:�/ƻ����������^�����L�=���=I���M��U��J���q��e���ܽѪ]�+�W�M�?�J@b�	��q��Tt��Nz��$0�1��=�p������I��"6,�RSԾ&���,~�������N� `�_�P�h�'?ɶ����ǿ����ܾ� ?�- ?Бy?��X�"���8��� >�~�<������铚���οB���m�^?ô�>�Ja����>W�>Y�X>�q>�񇾡螾k�<��?;�-?_��>�cr��ɿa������<���?�@�)??Գ$���۾y=�<_#�>�6
?��G>?�2����b�����>5�?�y�?��{=�U��0��?�\?1��<��D�����=�="�J=-V��L>O�>����.F�1���R+>y�>P2�J���YH����<=�a>1$�ᙯ��҄?�q\�c	f�A�/�JP��Q`>��T?kD�>}��=�,?$>H�:~Ͽ`�\�Y)a?�0�?1��?��(?�ܿ�ٚ>2�ܾ��M?@6?���>^&���t�ّ�=w�༴P��a���&V����=��>�u>��,�`���O�8V��|3�=����ƿ�����
1^=������,��gҽ�8{�u�{��W��?,��KL�Bh=���=�*e>�5�>��I>��5>� [?ͫ?�s�>u+�=���eY��EX׾��Z���V�4���e_�@���F���bE�r��/a���`�
�U޷�>)7��0�=�]��\��p��g���R��]?_d�=��� �G�+�<�x̾�5��Zؘ�#(�*}Ǿ}-�|ph�8��?.~6?�Q����I�&��}G�!�սIE?��v�B!�Ԑ���?�=�;*G�=���>�㚼d\
�
�4���G�l+?��?���d����Xh>����[6�;��)?hC�>��ּ^�>��-?k]�'�����S>��P>k��>3��>$��=�}���˽��?�NU?����r��y�>����q���Q�=>�>�X��N�<��C>r�U����b^{��<����=�TS?V�>
�"���$����T�9���=Ayq?E� ?Ψ>��d?5<?6�n���W�&�=�k=��\?P>e?�>�=[۽�3�� _���=?��f?5^`>���P߾/!,��e��9?�n?3�,?$@E���q�ih��B�߸,?��v?�r^�ss������V�Q=�>I\�>���>��9��k�>!�>?�#��G������Y4�Þ?|�@���?6�;<!����=�;?t\�>4�O�+?ƾ1|������ߕq=�"�>���_ev�����R,�c�8?֠�?���>]�������[�=�����0�?a��?99��h�G;�Q�/}f��� ��<)=5O�=�E���N�	��S9���ؾ5��?�������>��@Cѽ��>6hH���ݿ��Ŀ���t@޾3ɉ�ǩ?��>W�����ʁx�9D}�y�6�"rB�{D���ܡ>޴>_�ቾn!���A�<������>;�⼁��>�G��
Ӿ}_���мڀ>��>��>���殮�N��?<���5Hѿɣ������_?�'�?"��?�?���=�0_�< w��lq<��I?��g?��T?�����$=��j�<K��?�H�>���~��������>3�?���>O���:@
?K��>��A>�?;lT�%Fȿ����-������?ؿ�?���\?�1�?2`?2/%��{��d/�ג���"�=tE�>��5=��Ľ�K8��c�`!�)?�r�>Z;��7���J�_?ёa��p�c�-���ƽ=ޡ>4�0��$\����۶��^e�����qy�\�?�]�?��?k��) #��5%?��>ݤ���3Ǿ���<��>� �>q,N>�0_���u>v���:��r	>y��?�w�?�_?|�������R>]�}?7��>�~y?O� >Sn?}~>�Ӫ���U�h>R�=:��%��>��E?��>{�>�[N���9e=�ȕN����
2�P|�>+�R?�$Y?�$>!ô���a����Γ��� z��{���+н2�)�:}>�4>�,1>�?���Wݾ�:?{3�� �u���ﻆ��&f?{p?�C�>�M,�F�i�c��=�C*?�R�>r�����ߏ�����fc�?�c�?!� ?����*�q��6>J��>��>����
��&>\�!��=�OF?��_�~�}�K�K��Ô>P�?�Z�?>��?Hȁ��	?���P��Va~����7�h��=��7?�0� �z>���>��=�nv�ݻ��X�s����>�B�?�{�?��>"�l?��o�O�B���1=9M�>Μk?�s?&Qo���e�B>��? ������L��f?�
@u@`�^?*��࿿f��*�Ӿ%�ž�h�=�c�=5�>|D����=���=����X�f�E&�=!ƀ>t�u>�Z>G��>�FQ>��n>����4�*������8����;�*0	�z���2���羋���ܾ���x�������\R��e�DUE���?��|:�h�>,�H?4{<?1�^?�t?��ڽi��=F���]<�@���>>��>Ν'?��`?��?液= ӧ�M[�đz�$?���M��ߕ�>���>�ޤ>�X�>�C�>�M$=t>��>��=ނ=�L�=}ď=�O%���>���>{z�>݊�>F<>u>�ി%���Gh�vw�:�ͽOˢ?�Ɲ���J�������1���_��=r@.?0r>����&п�⭿�&H?�,��^�6�+��q>{�0?�mW??�>�]��
�Y���>�Q���i�1�>�2 � \m�j�)���P>h?,V>_Kd>�z6���4�h�M������j>�,?8ʹ�� =�wkt�tE�X�ԾBZ>Z��>��Ӽ���?���?�}�G0h���=  <??~?,'����lx�j͕�+�O>6_>*�S=��=�#D> B���ɽ�3R��G�<�=��Q>H��>�F&>���=#W�>�����H�M��>UF>��>+`??-a?��l�kl�&yy��D��^>�>\�w>�6�=RE���=N/�>�j�>�s����������O�X>����0�K��j�d)e=)�ɽN,�=�̄=D� �P�o�6�,=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾYE?J ��0{�����˰�����=Zy(?V&-?fj�;?��ҽ)�=IH?���H���/�ÿ�TL����>}��?뎧??Ԁ�F�ǿ?-E����>��?ਊ?���>/�<�D)�����>�V]?�9V?"��>t[��.����?!��?��y?�
J>��?K�e?�x#?e
���V��¢�q�a�ϛ��>��d�?%��>������Zt��%���B6�L�f=�&�<���>�}=� ��(�*>k�<+�9�Cc��M�>K��<�?�=���>Gm�>Т>\��>С>v���X<-��i����K?G��?ȥ���m� �<כ=��^��!?�
4?W�f��'Ͼl<�>4�\?�ɀ?��Z?�q�> ���6���п�PI���c�<��K>r?�>C��>� ��HOK>�վZ�C���>rL�>Mݰ��Nھ)��������>y�!?���>n��=n� ?z�#?�k>mj�>�=E� <����E��z�>�j�>�?��~?"?����L3�����䡿��[��M>H�x?�4?�>#z��z���?�KI�L��Ӏ�?�g?�0���?*.�?F??g�A?[wg>���W~ؾ殽�+�>&
?���M8���(�4��	?�F ?�a�>ż�����r��o ��-�~?�2a?Ax(?�����q_�w���� �<�J���'���<+D�(>��">ހ��=S�>2ԇ=�w�*A��0,<��=�B�>�	�=�@3��S#�́,?3���{��'�=$�t��+F���>	K>_����,_?j�?��lz��z��LН���Y�Q��?���?Q$�?���C�h�7�>?rw�?W$?�W�>�Z���T޾�p:o�F�w����>�S�>���fᾗm��[!��K���\�̽�������>��>�'�>#�>b[�=Ǿ�>vOɾ��T5�����I�*����0�;�6�ҧ#�zȾ�yx�t���>���y��*=�>�{��>�c�>-D�>�P�=f��>�䍽PE>!Jh>%�>ꡫ><�/>X�W>�xͻ�#�9e� �R?F�����&�c������lJB?�+d?N��>sl��e������?=�?�4�?��t>Uh�2+���?RM�>���B
?�7=�廈�}<�������!�����_�>�4ֽ��9�f[L���f�QC
?9�?շ���̾6l׽�ǎ�f�a"�?��]?�C
�`p�����O��%�P���ts��6��`�Ծ<%��L��6l��⤌���&�{�<5Z?�2`?�Θ�!���->��;�i� ����=j��>ϣ�>g�>Jy�A򾜴�uw��W�7���X�g��>'-c?M�>��K?�n?N�.?��F?�ڙ>��5>Y5���?�VG�'��>� ?'P?�Q8?��T?i87?�&*?��N=���<p���J��>���>��>�?�&?&ϳ��rI�vN�G�T=�c��8?9�hs>��<�τ�+��cF{�߻">A2?`����9�����
�>ڈ7?���>�#�>p"��hJz��C/��:�>?
?���>�@���l�6B���>I�{?q�_z�<y�">u��=w�������&�=�.�b�=�\��b���T<��=Ŵ=%Dj���(�%q���ɻ�,�;it�> �?:��>�=�>[=��!� �)��g�=1Y>ES>>�@پ�|���#�� �g��Ty>Zv�?�z�?��f=E�=+��=z��=S��5��.���X��<g�?}G#?�WT?���?��=?�j#?��>+�.M��e^��v����?,?fZ�>I���Gʾ�ب��3�Ϋ?{ ?<a�`��n@)�W�¾!Խb�>0Q/�� ~�X���D�Q��|��㙽���?밝?D+@�c�6��1�񷘿�F��BhC?���>�>���>��)��g��E���:>�i�>��Q?�b�>��S?׃h?&�P?D<�>l)��c���#��!�o�I=�E?�d�?�?�?q?n��>(��=ʒ|��󾟍�M���/"�E�}�%��=��T>pl�>���>;��># �=�ꂽ�����Y�n��=$M�>��>~��>�?��S>Um����0?�I6?
����)��؅���l�T�����?<��?z`�>�;.J�F���BL��O�,?A&�?p��?���>�k����=2vӽ,s���kս?��>+�>d):>��=��=�2��$p���h�>R >�E!�Wg �*'=ԡ>�5?6ܩ>h�L�@���h���<���h-������>ND�#Ǽ���%T��sv���Z=��#��Ե����8�n������"�>�c=�7�>�5�>��<���q�X�/<���<U��=< +������FB�~������v���:=�fH=������06u?l�L?� ?VdB?E�z>�o�=E��ப>�hƽ�*?V�G>�vսA;���������퍾�K侰"Ծ�X�4*��ٮ�=s���6�
>��6>6>1�!=�d�=s�=�k�=󶤼\��<�Q�=��=v	�=��=�4>H��=96w?����{����4Q��X��:?�7�>���=Eƾ�@?j�>>�2��ϗ���a��.?4��?�T�?��?�ui�id�>���厽`m�=���<2>���=�2�I��>��J>��cK�����4�?m�@v�??�ዿo�Ͽ�a/>�C�=��z=��y���6��7:�P�Q��My����>�<���J�z>��b>4���A��W�
=o�>a�`�M*�j�7��N:��n>���=�>�ǃ>Ǽ8>�J/��?>���=�`s=�sM>qm�<��x��\ỡ�2=�H>O�>"P>R�>��/?�!?�!,?hXR>�B���оcȽ�0�>Wh=�Z�>��=��Vn?p�X?��U?Հ?�>J������>�B�>>U���x���վ����V�K���?]G�?2��>���<w��(bh��NC����>#�=?)B	?�	?�\�>=������@9��:.�O��<3
>~+4��S7�d/=^:��;��{����9>G �> ��>b�a>~w�<�=0�>�>*V>:�=D�=:ˋ<����2=�m�=R$x=��=�F<P��=t��=��߼`2���#=�����������V�A>��>�G�=�#m>���7����vs>k�u��0���>?���h*�ǜ`�r��,�;�Ch���o>�g�>f��=����#q�>�c�>��O��?aY�?Ri>z�	��ɲ�5R��FA۽A_-��^�=i?g�x��%Q���T���	�9f꾺��>��}>�}h>��>,2d�I�Z��_�=�ø�v5)�BQ
?�煾�x'���,������W���Ԑ��A�U%�=��T?�ׄ���>��g?L&??t�?�L�>;���N���}�>�\{�������Rľaㆽ4z,?q��>͈�>�W޾��,�d�����'��>P���{K��b��Ak���C�9D���"�>3�����4�s?��L����5F��������>��V?zA�?p~K��Ӈ��rp��O�7ۉ<�L�>��~?>�X?W�?���¢�wK ����æf?���?�7�?���>4�>A���X?>��>�S�?�?p�T?�n�%`�>2��vwA=��f�G�=7p�> �=���=��>� ?5�>�0-���ܦǾ?�� �@��=8n=qX�>�(�>P�>����d��<��">?<C>�ş>��>�>l7�>��=�8��W��-?�%�7��>߁(?,<�>��4�D����=����ՔὩ���b�q�1��ƺ�]�����">�$ �G�>�4��b�?�`>�aȾÖ?���}+�u�%>Uv�=B�#�MN?_Dj>/�>���>V��>Z��={?>�=�E̾�F>6))��$��L(��}P�]2�f�)>Zq���
e����5X���*9�:d�����R[�l����8�]L�:���?��2�<�o�lH#��[2��{?���>&B6?�ם��N+�x�<>�6�>��>��Ҿ,���V��>뾹��?�z�?�&c>�%�>��W?��?1I1��2�gZ�.�u��A��d� �`�l֍�
���Qu
��p����_?,�x?%PA?V�<'z>���?�%��͏��>�/�;��<=��>_#��6a�A�Ӿ��þUZ��KF>+�o?��?B?ۏV�J���v7�=�F?�}?��i?��;?�+?w���L?f��=�,�>���>��>4�8?B ?�UB>H*>��ֽ$��;Ird�0����`ǽg���m��K)�=�>�=ed�=9}��|�=iq�3s���=uĜ=�!� �T��=EŘ=a|C���>pI?�Y?�i>�??ai�;d�0���=�,h?�6��E�&�ُ�4Q�kK��``�>�V�?��?���>�1w>}�7�����h1>�a�>-�;>�> 'Y>n����H�>���>�B�>.L>��2;�r�����sś����>W��>��>HE��L>ڋ�t�p��i[>��(�� ��G�s���F�z�+�R${���>�oC?_!?���="�����ƽ�\��&?�57?��K?�q?[��=��Ծ!B�>G��FB��>�1¼�Q��쟿�5��E�:�{h2=?�O>����ˡ�j�d>t���侄�m�tK�����K=�
���X=#z�R޾g\��u��=�>����L� �𲗿Ѕ���J?6�=���ܑO��{��D�>O��>p/�>�p0��xf�uK>�t���+��=�f�>s�1>�N�����&�H�����>�o ?W{|?�3t?d�)�ڃa�����F��!��
6=�5?��M>��J?a��>���=0P�����̩N�Mh/����>���>��&�|��L '�?���?�)�?]��>�(>�+?c�?.?�>���?$�?��E?e��>�B��r���(?:q?���<�������E��/T��
/?�6?x�p�b�>�K�>�$�>fS?=W?Z�.?�<��o�	�-T����>���>}�s��eʿ�O�>LuU?�m�>\o�?���?�}�;^)�3��Fվ��<��>�=?#3�>�J?���>���>գd�u�>�� ?�"|?�Ή?6SV?�~=���>]�%=���>֓=[E>���>;w*?��D?Y7f?��5?ߓ ?s�=�Ͻ�`���~ �=?�={�x�k�=�o���-�� ������=���<�󌽸����h�=_��Q+o=X:��m�>�ey>^��"�1>[񽾧r���2>����难�f���]?���=U�~>�R ?+F�>G�)�C��=O �>E
�>����a)?d?tB?��L�;
a�Ěվ��?����>{�D?��=çm�#[��{�v�
�+=g�j?� ]?�WW�����b?��]?pg��=���þv�b�ԉ��O?��
?��G���>��~?T�q?��>&�e��9n���Db���j�.Ӷ=�r�>�X�T�d�r>�>o�7?lN�>��b>|'�=v۾��w��q���?��?�?���?u)*>,�n�14���������^?���> 렾`�#?���nξ~��;	������x��W���(���7ڠ�v�$��2��@sݽ��=j�?~?s?Bgq?�^?�l�:�a��^[���{�P�S��� �S����E�7�D���E��Oo�-h�if���A��g�3=D}E�G1$�(��?��?���<���>_��	��p��־�=����`��:�v>غ�*��=m�=�g���&���?"��>2��>�?��X�bJ�ޓ(���'���ھ�A>�3�>nr�>�<�>?[�<7
!��e#���߾I�����$��d>�Xa?��N?���?�t���^*�)�q���fH�=h��?��>]�f>#��>f;�����eP|�
�J��vN��@־��d�#

��>��?�U>@p>�?���>�־�ɉ��3������g����=c�B?�a�>CS�=Bd�%�ľ��>Өe?� ?Ͼ?,G��.�h�m�W�Ā�>�ˍ>� "?ԛ�>(�c�Qc4�����.����A�&�=�!Q?�7��߃�Sl�>=?�<}=IG�=��>63���3�����B:�!=T��>c,���:�>�꾱��JnT�h,E��d?�,?��������>G�?�n�>*��>�S?St'=�0��J��=]�>�e?�_?`8?���>���D��=���v��=��>��>ߓ>'@���ͦ�����%DǼ�6>JB=֣g=���=0�U�5=�4�=���>�&ؿ�>�	�־���TX�|��T|�Y��3bu���@������ ����d��)���=�&�k�O�\���X}��5�?``�?&@��/������Ä�C��4��>�w��-��P���ޗ�e�۾wG��k�f�#���Z4�[`d�)/k���'?������ǿ����9ܾ ?_C ?M�y?���"�/�8��� >���<sl��Q��ƙ����οg���"�^?���>c�~(��m��>-��>ȠX>�Jq>��z랾|g�<��?��-?Ǣ�>r�r�Ζɿe�����<y��?%�@*^5?����¹�����?���>���=�����;�*ȷ�{��>
��?���?��=m�R�B�X��M?l�J=��]�9bn�� >)b�=��7<����a�=?�0>~c\���]�qm�on>�f�>�m;=�ԙ�8KC��uV=1�>��<��c�5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�ޅ�=u6�����{���&V�~��=[��>b�>,������O��I��V��=~���¿��"�y���G=q��;R�D��.���%���Ȗ��0����f��(����%==I	>~�a>��u>7>X*S>$�U?�*z?:��>A-�=�&��,��j�Ⱦ:�#�M���|A����$&������A�<�þZj	����&�
�Y7׾H?D�k��=k5U�`+����-�1b��U1�C$?K�v>��� gw�k�A��F��m�ƾxW�=;�=��¾��@��
m�|K�?��T?Y���Tj�U$��v-�����-\N?R =6b�����-�9�<T��`�����>��d>���$W_���M�x�#?�L?�&ɾ>��v��=���K8����?b+?<�i��l�>e?Υ
���)>���>��>�4Y>1��>��>� ����\�?F>i?Eպ���վ@x�>{�̾>���$�>��=<
�b��=Kg>ļ~v��y@0>�>�w��=�V?�]�>!I*�͖�'�������/=�y?��?�t�>��k?��B?⟁<���}R�
�	�"qo=ЀW?ţh?a9>���OCϾ]g��c6?�d?d�G>Li���/����Z{?2o?j\?3��}��Б�����6?_D�?�̐�Y{�������R�3?�e	?�^�>5����B?b�p?2P����7��ٳ�Gp���V?��@z�?\����1���>��>G�)>�?l�ᚾ;��Y�_�]<=��>�?���/��#�F[����?�q?��>�H������W�=�̔��ʫ?˅?�餾��+<�~��Sm�'���I	�<��=���� ��쾹�7�Frƾ8%
�嚾��� ��>��@�Jݽ���>�;?����A�ο�����Fоlm�0,?��>X~�����5ii�1�r�`G�;$I�nO��!�>�9>�����J��_�|��	;���hO�>|����l�>��N�ў��>��
ͩ<֓>���>��>���Ҏ���\�?�����PοkR��C����X?CĞ?���?+� ?�G�;�u�� {��t��#G?f�s?��Z?��<�"7Z��6C���j?,���os`��}4�~^E��sU>+;3?I�>y�-���=3�>�r�>��>�./�p�Ŀ9ض�Pv��6	�?at�?2M���>�v�?9�+?�K�w1���ת���*�fZD9�5A?��2>�z��Ž!��=��i��6�
?�0?���z��_?��a���p�X�-���ƽ�ۡ>��0�Ye\�K������Xe����3Ay����?<^�?P�?s��� #��6%?�>T���
8ǾM�<l��>!)�>�(N>�J_��u>����:��h	>a��?Y~�?2j?󕏿�����U>��}?���>��?h��=� ?"�=�����<D��M>)��=<-���?C-M?���>���=��;�_�8��G��iM�:-�R�=��,�>��_?u!J?�f>������-��V�u3��tEA������I����4`�]7>̦&>q�>i�A��D̾��>?��E��Y޿�%��G	���;E?~y�>��>�bR�*�=j��=�*@?>�>�/*�`���5Ñ��X��*�?a��?ٯ�>�A˾c	�<���>��>�w>T4ǾK��sم<�4>�Ul?�)�������*��~�>�9�?g@�۷?���<�	?�웈��H}��=� �3�i��=�7?��;"�>l��>�e�=��t�󜪿�t��U�>�T�?���?���>��k?�o���A��dA=�Ѥ>�Pj?m�?�ú�ﾤdE>�t	?�R��Ď�3��^f?��
@�@�^?k{���׿�S���0��_Y���/�=���=g�>� ��$*z=o��=�Y��ꅻ�2�=bsz>�[:>췜>S�S> �,>0W]>D���w&�vি�ט��C�N��ʂ��Ar��P�\�������U��sH���C �`R\����<T3_��V�,P�<q%�=S�U?ҏR?d�o?Y?58e��>E����V4=�R.�Mj~=u��>V0?[�K?��'?K�]=ET���d�{�}��򤾅������>�IJ>;�>;��>��>��<�/N>��C>�c>�y�=E�=	KH�=c�<6�R>�0�>&�>+�>��=��:>����.���(c���#�ܽ5��?��8�@ 5��ܠ�nO��L5 ���G���1?L#�>G����Կ�Z���tJ?2���H������D�.>6��>��N?���=Eī���%�2>��J�j�v�m�=��G��獾��)��j�=2 ?�y�=%'m>�3���L�	1��6�	��>��>�$�D�ｭF������چ2�0�%����>i�>��+������] ��{��Ja?��?�=�B��8
>%��Dy�T^(>��<X0M>��I>no�>=��Y@ھ�eX��\7>�l�>��?TH9>��=Yͧ>�ɔ��KQ�E��>�)R>c�4>��=?��#?�������A{��l ���{>���>f7x>%!>�xQ�	�=�#�>�]>�����t_������H��b\>�5��s�f��b� O=�Ʃ�J��=g^�=-u���F���#=�~?���(䈿��e���lD?R+?^ �=�F<��"�E ���H��F�?r�@m�?��	��V�?�?�@�?��N��=}�>	׫>�ξ�L��?��Ž5Ǣ�Ȕ	�.)#�jS�?��?��/�Zʋ�>l�}6>�^%?��Ӿ�{�>�4��_�������L���w<�;`;?8[?�dU�Nغ>᜾�h�>��?�(F�1l���$��=�D����>���?0�?C���TK��=�����>���?T�:?8t�>;TC�kڽ��>��j?�;�?���>_<��%��˺?�b�?I�?\�C>	�?��;?Z?F��z@�~-��}�����=�f�=�e�>�f>4���� ��2��K���~^T��r�*s?=5)���/�>�Z��RC���U=%��X����v�=�v�>���=�_e>6[>+J�>��>��>P�v!轡�]�����K?���?<���5n��I�<��=s�^�g?�f4?yb�XVϾͬ�>]t\?�Ā?�
[?���>���r#���ҿ��w����<�/K>z��>�h�>Z���N�J>��Ծ�%D��A�>��>,��_ھ�n��0����&�>Jt!?/��>�B�=(h?�Y%?�b>�W�>�D�����hdM��K�>d��>T�?z�|?֐?�찾�5,�-,��*j��lgX�΍9>;�r?�?3�>����q�����c�#∽�Ӏ?�;^?�� ���?�#�?P�3?O*H?Ώ�>��H�z�۾�>��?��>W}!?WS	�]A��J&������?*?���>S����޽����G�����fc?v\?�&?����`������+�<WQ��@\��-�;�0�@_>�>,����=�L>Ә�=Ti��B5�c;<8�=*@�>Š�=[;3�XJ����,?�E�<������A=��C�,�l��>ZL�=��վ�Ia?%��B{��w"����񀪾^l�?�5�?Y٠?Jm���s�M�;?b�?`�?G�*? ��d�e��"�>Iwt�	�8���Q��7�>c+O=<����k�������J�Ξ_����>{�?�$?��?��3>c:�>��ξ[
�9���˰�˪7�϶��I*��i��A�����'C��^<Y¹��p�2�>��o�2ɧ>�p�>��>C�>�b�>�H�=;]>�GS>-B�>!G�>�>��>���=��ٽ����(JR?����!�'���&����2B?�ld?�,�>hi�≅����ɀ?��?�q�?�=v>W}h��++�pl?�:�>����q
?/m:=w���<V��3���)������>7׽�:�$M��tf��f
?�+?�$���̾�B׽ω����=�|?o#?�x�FVM�	�x��a�JGM�wO#���7t�K���b������Px�u�&�����?�ʊ?�U�y#��f���P^�+3�jq�>sO�>H�>��>�-=�n��@���j��?�d'e�h�>�p?~5v>5RN?��?��F?L9I?�w>:��>��3���?�uf�w>��>Y��>B�1?[v??�F?��?��=Ш�=�����;�K�>�>�&?\�?Nt�>*_ž0�缰+���7����P���ɼ^��=���}<�锽�9>�T?�&��8������#k>4u7?�.�>��>p叾"i��$%�<Z�>f�
?a�>�����`r�rW��]�>(��?MB�<T=��)>�Z�=x�������,�=b��D֐=wˀ�J�<��~<�#�=@Ŕ=Pq��a߹R(�:�2�;�X�<�t�>7�?���>FD�>�@��h� �����a�=GY>�S>M>�Eپ�}���$����g�]y>nw�?�z�?z�f=[�=җ�=�|���T������������<�?`J#?TXT?P��?P�=?j#?�>�*�=M���^������?ui*?���>ϻ�X̾)�����5���?�=?=8_��j��{+��Ⱦ.��B>*.���{�g���}�E���)����$G��ߕ�?�1�?�;5���5�Q;������xwB?��>)o�>h��>U�)��h�����8>��>�6R?Hî>�z+?���?�O�>�֦>[��f��#C�����ڸ/��kE?��?d'�?Ct?��$>��=Rn���˾��2�>�F���桷�y>>fo�>��>÷�>�V�=��q�~��� ꣾ����7�=���=���=aH�>力=�:>�FE?�3?G3׾�2�����;���i�K��?%��?�T?�A+>�����V�QN�����>6ʪ?�M�?j%?x�J��\�=�#�<X,̾���P��>IO�>���=؈_=H�/����=���>��>�*#�i_"�˟7�m��^�&?��T?H�^>� ƿ��q���p��ė�&�e<�ޒ��d�|�����Z��]�=v������-�����[�����Tx������٩����{�"��>��=��=��=˨�<)�ʼ�Q�<�K={�<�=�p�9�k<�H9���ԻS����l�P�]<DaI=%������x?��_?��%?��@?��>�?+>o��<ן>���Ҋ?��a>�|A��"��-�S�����ƭ����߾FD���^j��˥����=�$]����=��>�]>@�μ��>&��=h��=��Ղy���/>��=��%>P�>_�>���=�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?��>>�2������yb��-?���?�T�?>�?@ti��d�>L���㎽�q�=M����=2>q��=w�2�T��>��J>���K��D����4�?��@��??�ዿТϿ6a/>�58>g�>��R���1�Z\\�T�a��>[�{"?m�:���̾cц>���=��߾��ž��2=<�7>�t_=�����[����=W�y���;=�vl=�S�>wRC>�͵=�4��\-�=�VE=��=̡P>��X�A\:�9Q.��~-=m��=r]c>)'>���>��?'�9?R�U?�D�>�c
�wmؾ�R����>oC-=�[�>��=�`�=�Q�>�>?p,?��7?���>%�=Y=�>���>���[bY�������	7�=��?va�?N��>��=�_V�p#�b�G�I�	��>C�(?`��>���>�	�4�ҿg7�P�-�y?��۲>;��=���;r��=�4�=��62$�qȭ>i4�>n��>���>�y�=\>�f�>Y�>Mܯ=�r�=�D> ��:g�<êT=�"=��<1��=��; o���U�=O�R�X78����=�h���4ནh_���>���>b�>�>�@>"����">O���0����=8~¾��G�wBS��䀿��2��7���]>?H�>.kH����u�>���>%��=H)�?��u?��)>�5w� 7���X��M����qT=tW�>��>@T
���U�'��G6W�[	��d��>2ގ>t�>��l>5�+�/?�Z�w=r��\5����>Q~���i���X2q�=��b����i�պ$�D?B��a��=~?V�I?
܏?̊�>b󘽀�ؾ�'0>D?���=�
�q������?I'?D��>��l�D��̾pT����>�eJ���O���/��2�)㷾��>C�@�Ѿ�33�"���4���OuB�@mr���>��O?��?F�d�$_��HO���K4��`i?,�g?�&�>0�?��?iܞ��X뾷���%��=Y�m?��?�T�?6>��=�ݴ���>��?��?_��?]@]?�j�[��>zo�����=r&!�ߥ,�&q=>�?>���=�B�>a�>aV?5S��~����侯p۾��G�~=�Xy=�f>���>s�A>Kw_=ɓ=��={t>���>˒>��W>mN�>^w>L���,f
�q%?w�=��>Y�1?z��>4v*='F���<������6�-9%�~����ݽ���<���*�j=���_��>�8ſ�a�?�KA>�� ���?-���i7����G>`#J>5+ӽ-s�>�PU>���>�F�>Qy�>{�	>���>5�>��̾c�=̐�_�)��>0��w���	�H�=�y���հ�1��Ǫ�)ѫ����=���_U�(.y���P�݄�<NN�?�c��q'W�wt%�	_����	?-��>�3H?�J�p]*>��{>���>y��>Yd��Z쮿ꄓ�U�5���?���?0;c>�>��W?�?}1�53��sZ��u��%A��e�Ż`��ߍ�U���Ŕ
��꿽�_?�x?�vA?<H=z>��?��%�^я��*�>/�A%;��8<=�&�>'����`��Ӿ�þA�SCF>}�o?-$�?bY?7TV�Ƅ�9���>}Z<?�8?�?�+T?��?NK��H:?�����o>-Z�>h��>��7?�90?|>v�>����r>E���rR��%Y �CO����="��=ʂ�<}���:=R=4���gn��m�54U=���=?8t<�)�=���=Ԩ�=.1�=�Ɲ>iX?3I�>v�~>�A?Ѫ�3 <�����%?m�@*��2[�������ƾ�,Q>�Ek?�M�?��I?��>��&�Q�7�^y\>�Y}>v�>�{>��>p
�)pA��n�=��=;>��=:ٽZ�x�����J����<0$>�B�>�y�>�O�v�#>`���\��M>�K�����',i��I���*���{��>�uN?�~?3��=���4�^���^��*?��>?FuJ?��v?n$�=B�Ѿ�@1�O�C�������>(�<�	��������A�L�y�i>7���x񠾈�b>���J޾?�n�j�I����J=4��qzT=� �P�վqu~�ާ�=��	>������ �����Ϊ��J?Uk= 4���U�<}��/�>-��>��>2�:�C`v�Bd@��W��Cۖ=�~�>��:>�y����RG�X:��*P>�_?�I\?J,X?H*�(�c�J*������ɾ����`?2�>��"?���=D�t=�U׾��&�f���{�h��>R�>H����b��U���վ<e˾E�>���>4�[>s�?��|?�v�>#h?�<?��??�#�>-�x㲾H�!?�Z�?�>���aI;��Ay�k��>��?#\
��^�>��-?�o!?	f&?�%7?~�?k�=j��<�c���>��,>�%T��O��/�{>��P?�ݣ>��@?]��?:�>�	2�oL����>�z>��>?oF.?�J3?B:�>p%�>A���B9�=�i�>ܬb?t*�?g'q?��=9#?�34>̆�>
\�=1��>���>�+?TN?��s?ؒJ?k�>1�<[V���D�� s����w�D9K;Z�<"�=u���q�
���<Ig(��!ȼ-�����nE���f���<�^�>��s>����0>��ľ(M����@>����Q���܊�S�:����=邀>��?(��>tR#���=���>�F�>����8(?��?>?�#;(�b���ھ��K���>�B?}��=�l�e���z�u�v�g=��m?|�^?�W����,�b?�]?�g��=���þ�b����:�O?��
?�G��>��~?m�q?!��>��e�
:n���.Db�X�j�qҶ=.r�>DX�}�d�k?�>l�7?�N�>h�b>�&�=0u۾�w��p��/?��?��?���?�+*>D�n�(4࿠]־�@��T�O?\��>�I��^�-?��<�f������ᠳ�����������hz�K����ͽa	���;!�P=���>�"|?}�R?|p?���,���M�h�B9��O#e����������5��`g�Ӓs��$�Ҳ�]1���	>�I~�ƈA�[�?�p'?��/�ˁ�>A��c��~;(/A>y������P�=��p�;=lA]=�$i�K%/�8^����?GҺ>���>1!=?�n[�v�>���1�
<8��~����2>�H�>Dȓ>Y��>ȧ��7/��
�K�Ⱦx胾.�н�5<>�Zc?�~=?��[?���|b��y�Mv.�$ ���ZԾ{�>�s=�s�>I��]�P�?��=�0�~����cD���������=�� ?��8>�{�>m��?��?�`��xþ�A|�:�A��k?>�|�>ů]?�Q�>���>B"�XJ�2�>Pwe?�Կ>�H�>�̇��q�r����iҾ�)�>p~>�k�>��}>Uf��kY�p�������DF���>4�?䃚�\N��S>ޒ4?qC�<���= ��>5�=���p徇Sƽ��=dO-?,���[m>#|��6k��y��bZ���3.?n\?��v�h/$�0��=��-?��>^<j>Ӕ?�?y��:�b=��?��f?zB/?��8??��>��=_ �?$��3�:�
[P<j8�>��W>�O=��=j����� ���4o(>�K<O���}�B�P�)>�6�=t�=ȝ�>"�⿊�>��Eھ�P�"����	V�����틛�b!ս�ꭾS�����U�L���?5����n����=R���ӆ�K��?���?�R����>����v�`��@>�ͬ������[�r�an������Q���c.��J�
�c��Y�P�'?�����ǿ򰡿�:ܾ6! ?�A ?8�y?��7�"���8�� >RC�<�,����뾬����οA�����^?���>��/��q��>ݥ�>�X>�Hq>����螾l1�<��?6�-?��>Ŏr�1�ɿc����¤<���?0�@*A?<�(�e�쾎�U=���>5�	?�?>'1��B��ܰ�/I�>d9�?��?� M="�W�^Q	�B�e?0�<k�F��/޻���=~��=�=����WJ>gC�>����SA��sܽ�4>�Ӆ>S�"�����G^���<�U]>� ֽd:���,�?�m��m~��'���m��>�?�$�>y�A>2/�>�d�a����h�%�X?��@�5�?ѷ�>��׾�:�>�3߾օv?��F?W(R>I�H�-c�×;�\����ҽf^;���K�hr�pI�>�z<>M�J�����H땽y&�=��3>�N�����.���"�9Z���I`����M�ν�ƨ��ݕ�����+ag�/˽�j�=��>I�%>�(>*&>
� >^O?�s?��?�h>ԛH��͇��
��_R��������$n)�P�$�G���~�ɾ׾A����!��X ��̾6!=�\�={6R�D����� �-�b�M�F�#�.?ft$>9�ʾV�M�8�-<�pʾM���e؄�%ॽe.̾D�1��!n�)͟?G�A?b�����V���UU������W?CP����"ꬾ[��=@���N�=�#�>釢=��⾘ 3�~S���1?�'?�ʢ��<��s�=~2���1�=�"?��)?�Q>!A�>L�$?�����EM�5A/>շ>>��>C��>�>ɶ��U潑?&&y?�Ž+�e��>S��t~�S����A/>z�Ž�li�[�,>�O@=62��6�J�,��~g�=�(W?͛�>u�)����a��.���Z==��x?!�?�.�>z{k?��B?;פ<�g��\�S����ew=��W?*i?ٹ>V��� 	о���#�5?1�e?9�N>ah����g�.�U��$?��n?�^?�z��w}�]��c���n6?T�|?�h~�G���9�tx��;��>���>��?~���U
?��8?�4h�H�x�/Ŀ}�?�eP�?y�@[��?�j���,�3�罿0�>��>ܠ>����bJ���y���#=���>����@��7������>?�i�?��>��վ]�����=_���Ȩ?>M�?�妾X��;��'�e�y��<|A�F�|=ʏ����[�q:��o�9�j��]���_���	����>�'@���T�>W'$�� �D�Ͽ�'��U�澨#y��s?l�>M��$^����d�~�r�4X:��M9�F-i�3K�>�	>�l��X���o�{��q;�����>B����>��S����|���5<@�>j��>�>�������Ù?�\��{9ο������]�X?Pe�?�r�?�v?p:<��v��,{��;��2G?�s?1%Z??�$�$]�S�7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�b�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�8na?+e�_Gt�P,�'ᦽSU�>�h4���H������E���e�R���E���W��?t @�?
�%��m#��#?�I�>����� ���s=m֒>Ny�>x:N>��T���}>���=����=}��?�4�?di?&�������B6>8~?B�>��?��=br�>��=���,�E�">���=�wA�r?aM?���>�K�=}%9��@/��NF��PR�<���C��	�>��a?JgL?��a>⼹�E=1��� ���ͽ�/1���|'@�.k*�Y�߽?Y5>ܛ=>�>�D�4kӾ��?2r�8�ؿ�i��zx'��74?"��>;�?*��[�t��M�w>_?�u�>S8��+��-$��S5����?�E�?8�?j�׾Fn̼%>���>P�>��Խ�埽]���U�7>��B?���A����o�/�>7 �?C�@�Ӯ?~i��?>!�V����샿6P�Q�=�S>6@?�����Q�>5�>sE�>�/k�oW���r��`]�>Y��?7��?�?��?����M>��=>���>頁?��?�O,>��ɾTى>9�8?��߾�FK�	��*K?O�@�D@b,>?'���dfۿ�#��N���G,��P��f'1<9Q�>UZ�=��A=�t�<�Yr�����q�6>�Ig>[k>9|>�2@>4UK>#��=(���^��P��:N���?�����������پ��x�?������_�����8z��Fnl���8��3l�K��=�T?T?1�s?�%? gZ�uf5>�x��T:=xU��Ħ=*��>�86?]�Q?��(?�>�=�9���c�H����x���/���>;9G>���>e��>	\�>��%���<>�#4>��y>��=��q=N�P��<��N>E�>��>i/�>FD<>�>Jδ��1����h��w��̽>�?7�����J��1��<������e�==b.?��>����>п�����1H?�����(���+���>
�0?�cW?�>"��S�T��<>(��-�j�c>, ���l�`�)��$Q>(k?#�h>��j>��0���7�`N�zƤ��~>�8?$ٵ�H�>��Mt��>K��ݾ�O>r��>嶰�2��er��e�}���h�6�=�
9?r�?9��������t������LL>~�U>��=�q�=�)L>�i���Ὦ�L���7=���=N�\>�M?�<>¢�=KA�>(����,I��P�>C}E>�U>)C?
(?�]�����Z�v�b/�p�w>���>��~>��>'�P�䍤="��>h�>&ܼTSŽ/Lʽ� ���L>z۵��CQ���6�A��=�&��8��=�}l=V���w=�n�H=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�'�>f���V���&����u� �!=�f�>�H?���f|L�8�>���
?��?<��^�����ȿ�dv�pv�>m�?Y�?�1n��c����?��!�>���?pY?��j>r�ھ�IY�ی>@A?�Q?x�>)��u%�;7?dݶ?�}�? ��=+�?�@f?���>�@"�����u/��r�|��$>�l����iN�����B���7q���'��c<'�=�i�>c��+����,��ͽ�ȝ�����i�> ؖ>S�]>G�>G��>�*�>�Ԟ>P��=����<�b���߾�K?��?��i�q� �r�Z>��?����>mfI?Y��=Š�����>��Z?���?.�K?a$�>�����󐿁3��&(��ޏ�����=�?)m�>����2�=_��X���K��>�+�>����k�ξ��Y�����f�>]q%?P��>�i>�� ?;�#?E�j>D#�>�^E�V8����E����>š�>�D?��~?C�?�ٹ��W3��	��硿��[�MUN>f y?fO?�ƕ>A������F�UI�S������?�wg?�,�f?f3�?�??��A?�f>���ؾ�,��>Cs?E����j��.P1��{�=�*9?�`�>_�)?�~ｊ�3�T�i�[T�����3�>~*B?��=?����h��a��(�
=xɽ�"=5�=��M�~7�>�܂>L��=D�>��|=ǅ3>H驾RH�<�>�w��Q6x=�>�;	-�^�=,?��G�ۃ���=k�r�xxD�?�>�GL>���@�^?o=�+�{����hx��FU�� �?Ƞ�?5k�?����h��$=?�?_?�"�>�I��)}޾C�ྌOw�	zx�w���>���>R�l���=�������8F���Ž�c���>�8�>�g�>^�?A�6>#�>/T��Fe)�����A	
���`��!��5�����������>������H��P��f�>볽���> �?U��>D��>�h�>�a�=P}o>
�O>M��>��>�"$>��>nM�=�F�/c��KR?�����'���辵����3B?�qd?z1�>�i�3������R�?���?Ls�?�<v>�~h��,+�an?h>�>=��Sq
?-T:=�0�Q:�<"V�����4��-�&��> E׽� :��M�Lnf�Aj
?�/?	��y�̾Z;׽�n���@�=�|t?��?���]���y�n{e���b�o���(>�q���.��cd��Q��om��6��f-� 6��;-?,N�?�ɾgi�Z����\���%���O>�j�>�gK>��>�*0>=A �cL���k��o8� %��[��>��z?6�>�lH?D�H?G9�?�#!?��6=�u?��<�b)?q�.>�?c�"?�H?��]?��?���>��1?�� >����������-?�F$?0�3?���>�?p�����ľe��gG���Z��i>��>���=H����;=�T?��E�8�K���5k>��7?�}�>>��>=���>��=U�<"��>��
?�K�>q����er��g��,�>Õ�?��[�=1�)>�_�=׀���ٺE�=�(ü���=]B��mM;���<���=��=��\ٹ��:��;���<�Y�>�#?٦�>�Z>�����,�	���A�<��<��������ɏ�~���o�p��l�<_g�?�"�?fgY>@LR=g�>�衾;�Ͼ����8��?�۠>`�M?zX?@q�?��D?O="?{E>�:��ɔ�����"%���	?R!,?��>��{�ʾr񨿬�3�Н?�[?J<a�����;)�]�¾��ԽX�>�[/��.~����)D��	�����1{��Λ�?���?�A���6�Uy�����~\���C?$!�>BY�> �>��)���g�x%�j2;>&��>MR?o#�>��O?%;{?W�[?:aT>c�8�s.���ҙ�Qh2���!>�@?��?��?Iy?np�>x�>8�)��ྥT�����a�ނ��DW=!Z>���>v'�>l�>���=� Ƚ(N��K�>�f�=,�b>��>�>�>S�w>�b�<��G?mY�>�澾UT��Q��y�����=�cu?Ґ?c,?�M=i�zE��%��H��>�?�?�?+�)?��S�ް�=�8ټn��h^m����>ȸ>Iޙ>
�=j�G=z�>��>XV�>C��bu�~78�lO�-�?
�E?��=NfƿZ�p���r��ޘ�L<:쓾�Af������]�.h�=^͘��8�:��y![��p���n��	���Y��ؔ|����>4q�=Z >���=&�<�ӼH�<�O9=��m<��=��n�V8_<�]G�G��ʿ��5����!<��?=���%ʾe�|?��F?R*? a;?��n>�D>ږ���L�>4���?��5>������l�E�*s��fs2侗 ؾb�.֗���>J`7�y��=b�!>c�=&��<&��=�|=�sD=���%�d=D�=F��=Ү�=�=4�>��=�T�?\���c��f9?����>ir�>3%3=Q��>'5����O?�b�;r;�Z�����=$s?���?+u�?�l�>h���o�>w�
�j���B@J>ŵS�� 9;䙨=m(P�Hͭ>Pq.�v93��H��4o󾄾�?Z�@D
L?󀥿�Ŀ�g�>�8>>��=Q�%�1�G�P�A&a�s�[�c!?�X;�c�̾�>D��=-�z�ƾ�r8=�R=>�Y=:)���Z���=�����L=Cs`=E݊>�XJ>�$�=�����=�
k=���=%|O>�-D��D���>�+�,=Ž=��Y>t�!>���>�?�`0?�Ud?i!�>��m�b�ξ�;��|p�>���=�[�>#�=$�B>S��>5�7?��D?��K?���>��=���>��>ʍ,���m��b� ا���<���?RȆ??��>�IU<ߗA�K��He>�"�Ľ5i?#M1?�i?U�>W����ڿ��2�Yy4�� 콋�ȼIM�=��>�&u�yB �/U:�Ӧǽ{��=�ѣ>���>��>J~\>6>t=>�w�>d'>.s=Lů=@I<��w<i��������Լ��b=fq�?񔼒�ü�>�;�҄�-v;�'B�)S�9��7=�=�|�>�4>��>W�=a��^�.>c��z�L��=����>B�7Od��*~���.�D 5��eB>�W>�烽��&�?.�Z>��>>wu�?�Ku?R!>_+��{վ����BJe�9�R����=K�>|�=�P];�@P`��M��Ҿq��>}�>��>ڻl>,��!?���w=W�l_5���>�|��3���'�d:q��?��P����i��պ?�D?�E��z��=2 ~?o�I?�?T��>!��Ёؾ�-0>�L����=���q�1o����?*'?ە�>��a�D�bD�����v*W>k3ɾ'N^�"ȋ��$���r�}%¾-�>4vž�䔾t1�gs������ߢW�w]��n�?�~?�F�?�E��n��u�T�c��s8�=-?�X�?��>l�'?�T�>��A>E;���sE��H�<vz�?L��?�U�?ЎB>���=xD��|'�>��
?0f�?���?��t?��>�$��>X��;M�&>l���Q�=�h>Ί�=���=��?h5
?��	?@�Z�����p��`�v��<L��=T?�>��>BIr>���=�-M=��=�X>dQ�><��>ac>o�>1҈>���s����&?K��=��>2?��>'�_="���5�<��S��}A�8�-���F޽�R�<�����zG=�aʼ���>�\ǿ7��?�S>��FY?���$��T>�4V>�i޽�	�>�`F>��|>��>���>vM>�7�>��&>۟�/T>�C�8�!���=�~\�\l�n��=�پ�7P�ho��g��=C��1-پ���x�w�V����g0��6J=U�?r� ^e��-<�z�.�]j?���>��5?YT��E��l��<p�>ɋ8>�c������c��өѾ
��?���?-%u>�,�>��6?F�?���;q�׾=N���i����<��?Ca�V=��XS����&��b�ܙ3?�q??I?6�D>�_r>-��?��
�B�����>�$7�� ��:�i�G>ͯ��[���Y����i$p��K>VB?�E�?�:?K����<����b>'r?�*�?;A[?;�W?��?�����?}={>��?)�<?Jt?�v?��%?=ɵ=Ҕ�>W�>_̣:ᝏ��g�.�<3��M�ݢ=p�ʽ�6�=�:�=b<=p">��o|ý�~Z�3��=\�+��qX<U� >��=��>��[?k-�>�f�>�6?H�-�P+5�K����W'?9�	=�V���ˏ�4&��PS��=4~e?�.�?�[?gk>�U>��68���>�R�>t=>��[>�ݯ>I����-��ؓ=��
>�>��=!]1�˃����F����=%�>�<?>q���P=9�w�:Ѭ�᡻�ED�|ϾK��gkT�ޔS����]x�>4J^?��@?<5�=~Ⱦ}�?=�e��2?~Fa?��?bb�?��1=����2� i[��6=߻�>��]=i��oǦ�a���iD��E�<9�S>W��4٠�_�c>�^�b޾�:n�~+J�����;?=����V=���v�Ծvs~��a�='�>�F���!��&���Ϫ�[yJ?�Ak=8̦�cX�Z)���Q>��>��>t�=���u��@���z�=Ψ�>�9>�ڨ0G����9��>Z]?�Na?��k?���nU��7�6V
�I�������
�>��>-��>y?>��	=�h��VN�-�h���n����>��>f-�N�W��CᾀO侂��Gd�>�?6�>TD?�rG?��?:i]?��=?	�?;��>׼1��m�*?��?9��=�l\�Ir����*�	-C�M�>��5?ĝ��~�>m�
?߸?&?FYN?��?r�E>z����N���>�V>z)^��ӱ��ߢ>��??�'\>W_Q?���?��>v(�np����T��7*>�j>�1@?�_)?�?װ�>s��>&Ɨ��4�>�t ?�,?���?\g?�{>���>��D>}k?OC��x�?l�	?`<?�^0?�e9?-�S?V�>#�;M�뽯H��i4G��4�н��1�:�5�*�ֽ�;�<KV'>g*s�"�ټ��ڻV-�o�μMh�ë=�_�>j�s>+
��f�0>F�ľ�O����@>쇣�%P��$ڊ�9�:�c޷=5��>��?#��>�X#����=/��>I�>6���6(?��?�?k�!;��b���ھ��K���>"	B?T��=��l�����q�u��g=��m?s�^?��W�l&��L�_?>g?���Y�2���K#���6���.?qN?�T�\�>��w?�=n?��>��F���1����h��c���M�=ӡ>�	���V�9wq>�%)?���>��>��1=Tվ=�u������G$?���?Xȵ?���?�� >�+Y�����Ҿ!�����a?9�>����a1?��R=e־�ܦ��þ;������ƾ�d��3�о�KĽD������n��=?|�H?��\?;Q�?����W� �q��ـ��_��ܾr�۩L��%�P/��ʐ��;�Œپ����d<Ɂ���j7�Y��?�'?�1%��1�>���iM����˾z�/>�Μ��+��ڛ=�@W�1*=Ȣ�<y�%qW��幾=H$?��>�
�>��9?�7U���>�Y�<�X�G�����|S>�
�>$ѣ>A1�>7�	�� <�1��Ӿ�������>"�?�?j~Z?��9�ɞ(��[��Ω:���=)e��A���W�=N��>���Vze��'c��q'�Z%s��+K�֮��r��wD�>0}*?1�=�P�>V3�?�x?�uP�9��� ����b+����$>�b?��?�tB>��"�t�ɺ�>B�l?d��>�>�����Z!�0�{�!�ʽ54�>�׭>ǥ�>$�o>ǧ,��"\��k�������9�Q=�=ݢh?������`��߅>8R?��:�zG<F��>�mv�B�!������'�A�>M�? ʪ=?�;>c~ž� �2�{��I��	G)?�:?/���ڀ*�:~>',"?�j�>@6�>q(�?[|�>3þk�V��?��^?�GJ?�SA?�Q�>A)=�����Ƚ�&�,=㊇>2�Z>��l=I��=M����\�����<F=~�=�*μ�y��Ú<>,����K<o��<��3>��տ�>�nּ�����y�ھ�����JS���w��6�����s����r�mԽ��z��(~��`��(�����?�>�?��$��(���������z��-!>`��ŝu������𽿪��zYӾuU��s
"��*T������g� q8?x/z��῍r��5p����?iΪ>�ȃ?�03��ؾ��R�j����^�:5��7� 
��'�߿`�*%h?f�?�����)����>��2=q��>@hY>��u��/W��O��34?��:?4s$?1���<�ɿ�Yɿ>lT�?��@�|A?.�(����V=[��>�	?��?>:W1��G�����$R�><�?���?�M=T�W���	��e?vS<G�F���ݻ5�=G?�=�F=���6�J>�V�>��HWA�n@ܽA�4>hم>�i"�٨��z^���<Ą]>�սwE��5Մ?*{\��f���/��T��U>��T?�*�>b:�=��,?X7H�`}Ͽ�\��*a?�0�?���?&�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=S6�Z���~���&V����=_��>a�>ł,�����O��I��Y��=����f¿L/�2����A��j&��
j�e{q���L��ͽ_W��Wx��f��cc�=��=�v>���>6N>�R2>S�P?$�?m��>��I>��̒���� ���ټ�g2�x�"��j���d�z8ȾGE��m������� ����־��;�H��=�Q�P6�����fd�*�H��+?6�>z�Ⱦ��L��!�<�ɾ�^����ż1���>5Ͼ8�3���m��z�?6�??w뇿�Y�=���S�k���;G^?x���I��+�=��
��
�<���>��=�-�3�2�Z#Q�;?��,?��A�m��>���v�v;`�0?x�"?=U>�{�>��4?�@���޽�<i>�M�>���>���>���=��̾
G���?R�w?�K:���ľt��>�������ΝB�B��=��;"�>�c�>W#���"ܾ�S=�u�����<�(W?/��>��)�m�t`������R==��x?�?�1�> {k?��B?���<�g���S���!xw=k�W?)i?Ҷ>􆁽оK|��z�5?��e?��N>B_h���龽�.��T��%?��n?d_?�����w}�������Qn6?M�|? gC�윿���4վ�6�=���>1	?ʺJ����>��<?���#ә���̿�H��ؙ?��@|��?�w�=X����zK>��)?��>��y����QF�o���� �=f2�>��;����2?*��s�h?���?�?v
s����*o>h����?7�?־2*=�X�׿u��>�������jވ����ݾ-V�9�ɾ�0�.ɾ�:�<]T�>�@�:a�W�?|O��2�3ֿ.��� 0����W�!/�>}��>\$���� l�ԇv�� 8��ch�B$��혣>���>���iԾM�p�?���J�7z�>�cؽ�\�>����> G��&��x]���*>���>>������	��Z�?+@��F�ܿ����(��h�4?�ۏ?���?��%?�s>G�z�_�$�u�O!0?�gz?�:�?[�����+����=�Ep?���Irl�>�4���M�?��=��*?e:�>��;���<�E>|�?���=w�H�:_ĿB"��/�׾�(�?���?V �ix?~E�?�n$?'�(�� �Q���Zr)��<����C?��S>g�ݾ9�2�?
B�A���-O ?�UV?��M��#1�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�"�>T�?���=`d�>9�=$簾�T.��D#>��=]_?��?\�M?�A�>L�=�9��$/��TF��HR��.���C���>��a?uL?~Cb>�︽�1��� ���ͽ�p1�Pb�FG@�"_-���߽5>D>>�>P�D��
Ӿ�O3?��̦�S����E�1�?�FC>�.(?p���k���X�䫀?2�f>?k6�����G���C�c�k�?1�?���>�ޱ�1H>��C>"�==�޼�V=Tb��ʓ��<�=d�s?�2�ӯ��ԃ�\ۂ>�þ?uL@@��?��j�D�
?�r������}�r��}�D���=<�:?0����q>3�>:�=�'w�-��6u��=�>�Ư?���?��>�i?�k�|<�<�5=*��>��d?L?*��#���I>�2	?Z��᏿����?d?&�
@@/@��_?�᣿��ܿ\��ھ'վb �=h\<�Km;>:����>.�=��H=�0��I=A~>dY>�#>Z�>�;1>��>5�����ԛ�I�����A��,�cL���Ž0�澇7<����f8�@p��  �=aKl�<ǣ�^n����Z�pv;���=]�U?��Q?��o?A��>M7v��>c%��cH�<�$�4��=0Ӆ>2?!�K?��)?P��=E����d�憁�xk��������>��G>�5�>=��>�Ů>��:"dG>�=>�*�>� >Ć=��L�=�UP>F[�>v7�>���>@{l>�P>�L��J
��k�,�T0���/����?~#վw�5�@	����*�����{{;�A?-�>	C���ٿ�o����U?h���c�2�O$�OM^>NG?�vZ?�j>5��v��=��{=H�˾������=�TҽR�_�E�5��B >� ?�f>@u>U�3��d8���P�Q{���g|>x26?b鶾�G9��u�^�H�}cݾ�DM>�¾>HED��k�W�����ui�R�{=:x:?��?�;���᰾̭u��B��KQR>�9\>Y=Ul�=yVM>YXc���ƽ(H��i.=]��=��^>V#?�*>��='�>$���"�M����>�)C>�D+>�@?�[%?�������G,��v>��>�q�>�<>k�I���=���>z{a>6@�D����x��?��UV>�z���]�cq�au=�ؘ��3�=h��=�; �Ug=���'=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�k�>9z�\�������u���#=��>:H?;Y����O��>� w
?�?�a�M�����ȿ�~v����>�?@��?��m��?���@�Uy�>e��?�gY?ti>e۾snZ�ޑ�>z�@?�R?��>�9�6�'���?H�?���?U��>���?��?��?O��=��%�v�ʿ�@��C�?����([����~>����!��&@��}��ZuI��~P�h~�>5m�<�X?��^�lN$���)>d��<Td�������.�>�s�>TV�>�BE>W#?La?s�^>�c����=��&��YI���K?���?0��1/n��L�<O��=9�^�� ?FL4?��[���Ͼ6ը>`�\?���?,�Z?;Q�>���)>���迿^��p��<��K>76�>�=�>���/YK>�Ծ�ND�*m�>Η>�C��8ھ�,������G�>�a!?_��>���=�� ?�#?�j>��>q0E�_G��4AF�=Z�>�q�>��?J�}?h:?.�����3�����ʡ���[� ^L>Gzy?.?/��>ċ��>����X)��DD����em�?�g?�F�;?E3�?{4??�,A?[�f>���ݟ׾Y���'��>��!?��A��K&���&?�P?!��>�9����ս.�ռ���jz����?�(\?�?&?6���)a�j�¾�7�<
�"�\V�d��;L�D���>i�>9�����=�>�۰=�Mm�8H6��f<\e�=�>���=417��|��� 2?�)=u����;J<"�����j�]�{>mAY>޽�VC?{�-� _�������������n�?R��?�{�?�+���p�4,9?�A�?���>�?0򐾂^���$� 5~�&}������}ܼ@�>Ws�=BFᾼ���:��x���� ���ڽ��?�а>H5�>�S?��<>P��>����a�+�֠'�����k�l'0�wV?���/�Ά"�hw���������ʾ�܆�HǼ>;@Žs&r>��/?cv`>E��>��
??~���O>߱�>�P^>���>H��>E<>&=�����-��KR?�����'�y������f3B?�qd?M1�>Yi�6��������?���?Qs�?0=v>h��,+��n?�>�>D��Rq
?pT:=�9�i:�<V��s��3��[�3��>�D׽� :��M�2nf�rj
?�/?�����̾�;׽�N~��)�=�bc?��J?EQ#���q�r����ڎ��2��S�[�Ͼ�p^�t[�f�!���%��N5���ZY���>�4?U�?͉5�s���0���Iq��q��c >�?�N�>l5�=%�?b��m��87�ǟ�ܸz��́>�}?�i�>sXL?ئ_?�Zt?xe�?���>=?����`�>X>��>��)?:�6?F?��B?��;?��I?�s�>ω[�RD�@V��s�'?5��>�?�r
?��?����V)��3��K�=���,>y�=C�>PHZ�~���x�>o=�=wM?Ȧ�{�8�����	�j>ۅ7?,��>���>V��� ��$`�<��>�
?VR�>�����jr�:S��]�>��?��G=�)>A��=�cߺ=L�=������=����q:�|� <-�=��=tz��Q��-��:��{;z��<�u�>y�?���>C�>�?���� �T���h�=�Y>� S>m>�Dپ ~��j$����g�7ay>�w�?�z�?Y�f=a�=y��=|���R�����#���h�<(�?+I#?sVT?3��?��=?�k#??�>O+��M��X^��3����?v!,?��>�����ʾ��Չ3�ם?e[?�<a����;)���¾��Խʱ>�[/�k/~����>D�����_��6��?쿝?dA�R�6��x�ٿ���[��x�C?"�>Y�>��>V�)�z�g�o%��1;>���>jR?>$�>B�O?#8{?��[?�{T>ܕ8�b-���ҙ�'o1�h�!>q@?��?U�?�y?�l�>8�>��)����^�������Nւ�W=h�Y>���>l*�>��>���=��ǽ+^��V�>����=ɔb>Е�>s��>\��>��w>�9�<*Z?i�?�����5�\GH�f��	mz�^nD?��?��?��7<���4�z�԰���>���?�?��?���A�	>��׽�`��T�O=���>��>k8�> >��=6&�=T�>R��>�`���'���#�am�x�?�6?@�w>�ƿ�q��.q��2QZ<�����d�5����Z���=}���o���i����Z�&Y���z�����X�����{�.��>5*�=vp�=q��=�c�<�x˼;�<�'K=A�<�/=��p���e<� :��dԻ�䉽� ��X<��I=r=����Ⱦp�}?o?I?�	+?aA?!�z>[>i2@�zM�>�w���d?��Q>!�V�󂽾">����C�����پb�۾L�b���>� ^���>�,2>��=���<7�=1�g=���=�:��=���=A7�=��=��=z>�a>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?~�>>�2������yb��-?���?�T�?>�?Ati��d�>M���㎽�q�=F����=2>o��=w�2�U��>��J>���K��H����4�?��@��??�ዿТϿ7a/>��7>�&>w�R�E�1� �\���b��xZ�՚!?�H;��J̾6�>��=Q+߾�ƾN�.=ք6>T_b=Th�pV\���=��z���;=-�k=0Չ>s�C>�x�=.���=¥I=���=��O>�v����7��(,�Q�3=���=�b>&>!��>�?uZ0?G)d?_�>b�m��Ͼ�<���g�>���=�-�><��=qOB>T��>�7?1�D?2�K?�k�>�v�="�>��> �,�$�m�9.�ٱ��$]�<���?�ӆ?�M�>�U<I�A�T��VA>���ý��?�K1?w?k��>�^� ӿ�w(�y�Z���׾;[w�8w=e�鼵�=�%Xɽ��<{DM=�zM>�h?��>i�j>bM�>��n=��=���>��>^ݖ=��>�%D;���=4�ü�<~<K�o���ӽ`���=��=���~�/��S����=�Gw<���+>���>蔶=��;>��>׺	���>М�p�U.��|��ŕt�J��>z��b�O�`�+��]>��>���=)�����>�D>�~�=��?`��?@�>�-�A*�����4����@�t^�=bC�>"�<��L�艇��zc�2�˾Z��>g�>�>��l>�	,�#&?�8\w=��W5�0��>和�_��@@�@q��?��b����i��L�J�D?�C��	��=I~?��I?��?���>�H���ؾ_W0>E��6=g��4q�Ȏ����?�'?���>~��D��J̾�I���շ>�3I���O��ŕ�&�0�^*��﷾��>Dݪ��о�3�b^��������B��r����>A�O?���?B(b�j���xO�.��qB��Gf?�g?9�>�<?�?�Ġ�*��Ϣ�����=��n?s��?�*�?>t�=�X�)J?RI?sF�?&��?��{?̦����>|�N=�b>�5޽od>6�F>��/>;�/>(#�>+�?W>�> �����$����]�Wv��:=g�0=�Y�>`l8>N&>��=���<��=�a(>ߵ�>�L�>4�L>���>��>瞄�L��	?wq����>g#;? v�>W��<%���l�Ɓ��~�M�3桾-�񽋒�x��'D%�O46>ӮU=ѻ�>uͿ��?��>z�$�~(?x4����	���)>�Р>�H���>
��>(�>��g>��>�y�=��><RR>EӾ{1>�V��� �<uB���R�cwԾ!ur>N�$�K�h��(�G��9�����+j�P>���=�6g�<΋�?�a���m��++������?�Ψ>Xi7?��������D>���>'��>>�������e���r�྽��?�]�?�;c>�>P�W?�?��1�N3��uZ��u�.(A�?e���`�T፿ߜ���
��	��F�_?y�x?*xA?D.�<*:z>*��?n�%�3ԏ�w(�>�/�w&;��@<=�+�>P)��O�`���ӾB�þ:6�JF>��o?%�?'Y?�TV�c��=	K��{1?��#?i��> BJ?!\=?X�>1��>�V�>��U?��e>�N?�'?�/?x�g=��="'�>�{=h�v��OU�\y�Ԍ��7��g�9�^�=?W�=��=.gW�*ñ�^½Y4B����;����-���V�=��L��`}=>�>��^?.�>.Xt>�+8?����&9�jE��Ğ8?�H�=��x����+��<1�:E>��r?d=�?yV?1pS>FB��GC��#>�]�>Q6>�JM>�ݼ>�k��^/O�H��<ە&>��.>XS�=hܐ�r��Ob����k�=�b.>���>C1|>���r�'>�|���0z���d>��Q��̺���S���G���1�|�v�?Y�>��K?J�?U��=y_�J/��`If�0)? ^<?�NM?��?"�=�۾[�9��J��>���>�X�< �������#����:�m�:O�s>�1��4٠�_�c>�^�b޾�:n�~+J�����;?=����V=���v�Ծvs~��a�='�>�F���!��&���Ϫ�[yJ?�Ak=8̦�cX�Z)���Q>��>��>t�=���u��@���z�=Ψ�>�9>�ڨ0G����9��>Z]?�Na?��k?���nU��7�6V
�I�������
�>��>-��>y?>��	=�h��VN�-�h���n����>��>f-�N�W��CᾀO侂��Gd�>�?6�>TD?�rG?��?:i]?��=?	�?;��>׼1��m�*?��?9��=�l\�Ir����*�	-C�M�>��5?ĝ��~�>m�
?߸?&?FYN?��?r�E>z����N���>�V>z)^��ӱ��ߢ>��??�'\>W_Q?���?��>v(�np����T��7*>�j>�1@?�_)?�?װ�>s��>&Ɨ��4�>�t ?�,?���?\g?�{>���>��D>}k?OC��x�?l�	?`<?�^0?�e9?-�S?V�>#�;M�뽯H��i4G��4�н��1�:�5�*�ֽ�;�<KV'>g*s�"�ټ��ڻV-�o�μMh�ë=�_�>j�s>+
��f�0>F�ľ�O����@>쇣�%P��$ڊ�9�:�c޷=5��>��?#��>�X#����=/��>I�>6���6(?��?�?k�!;��b���ھ��K���>"	B?T��=��l�����q�u��g=��m?s�^?��W�l&��L�_?>g?���Y�2���K#���6���.?qN?�T�\�>��w?�=n?��>��F���1����h��c���M�=ӡ>�	���V�9wq>�%)?���>��>��1=Tվ=�u������G$?���?Xȵ?���?�� >�+Y�����Ҿ!�����a?9�>����a1?��R=e־�ܦ��þ;������ƾ�d��3�о�KĽD������n��=?|�H?��\?;Q�?����W� �q��ـ��_��ܾr�۩L��%�P/��ʐ��;�Œپ����d<Ɂ���j7�Y��?�'?�1%��1�>���iM����˾z�/>�Μ��+��ڛ=�@W�1*=Ȣ�<y�%qW��幾=H$?��>�
�>��9?�7U���>�Y�<�X�G�����|S>�
�>$ѣ>A1�>7�	�� <�1��Ӿ�������>"�?�?j~Z?��9�ɞ(��[��Ω:���=)e��A���W�=N��>���Vze��'c��q'�Z%s��+K�֮��r��wD�>0}*?1�=�P�>V3�?�x?�uP�9��� ����b+����$>�b?��?�tB>��"�t�ɺ�>B�l?d��>�>�����Z!�0�{�!�ʽ54�>�׭>ǥ�>$�o>ǧ,��"\��k�������9�Q=�=ݢh?������`��߅>8R?��:�zG<F��>�mv�B�!������'�A�>M�? ʪ=?�;>c~ž� �2�{��I��	G)?�:?/���ڀ*�:~>',"?�j�>@6�>q(�?[|�>3þk�V��?��^?�GJ?�SA?�Q�>A)=�����Ƚ�&�,=㊇>2�Z>��l=I��=M����\�����<F=~�=�*μ�y��Ú<>,����K<o��<��3>��տ�>�nּ�����y�ھ�����JS���w��6�����s����r�mԽ��z��(~��`��(�����?�>�?��$��(���������z��-!>`��ŝu������𽿪��zYӾuU��s
"��*T������g� q8?x/z��῍r��5p����?iΪ>�ȃ?�03��ؾ��R�j����^�:5��7� 
��'�߿`�*%h?f�?�����)����>��2=q��>@hY>��u��/W��O��34?��:?4s$?1���<�ɿ�Yɿ>lT�?��@�|A?.�(����V=[��>�	?��?>:W1��G�����$R�><�?���?�M=T�W���	��e?vS<G�F���ݻ5�=G?�=�F=���6�J>�V�>��HWA�n@ܽA�4>hم>�i"�٨��z^���<Ą]>�սwE��5Մ?*{\��f���/��T��U>��T?�*�>b:�=��,?X7H�`}Ͽ�\��*a?�0�?���?&�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=S6�Z���~���&V����=_��>a�>ł,�����O��I��Y��=����f¿L/�2����A��j&��
j�e{q���L��ͽ_W��Wx��f��cc�=��=�v>���>6N>�R2>S�P?$�?m��>��I>��̒���� ���ټ�g2�x�"��j���d�z8ȾGE��m������� ����־��;�H��=�Q�P6�����fd�*�H��+?6�>z�Ⱦ��L��!�<�ɾ�^����ż1���>5Ͼ8�3���m��z�?6�??w뇿�Y�=���S�k���;G^?x���I��+�=��
��
�<���>��=�-�3�2�Z#Q�;?��,?��A�m��>���v�v;`�0?x�"?=U>�{�>��4?�@���޽�<i>�M�>���>���>���=��̾
G���?R�w?�K:���ľt��>�������ΝB�B��=��;"�>�c�>W#���"ܾ�S=�u�����<�(W?/��>��)�m�t`������R==��x?�?�1�> {k?��B?���<�g���S���!xw=k�W?)i?Ҷ>􆁽оK|��z�5?��e?��N>B_h���龽�.��T��%?��n?d_?�����w}�������Qn6?M�|? gC�윿���4վ�6�=���>1	?ʺJ����>��<?���#ә���̿�H��ؙ?��@|��?�w�=X����zK>��)?��>��y����QF�o���� �=f2�>��;����2?*��s�h?���?�?v
s����*o>h����?7�?־2*=�X�׿u��>�������jވ����ݾ-V�9�ɾ�0�.ɾ�:�<]T�>�@�:a�W�?|O��2�3ֿ.��� 0����W�!/�>}��>\$���� l�ԇv�� 8��ch�B$��혣>���>���iԾM�p�?���J�7z�>�cؽ�\�>����> G��&��x]���*>���>>������	��Z�?+@��F�ܿ����(��h�4?�ۏ?���?��%?�s>G�z�_�$�u�O!0?�gz?�:�?[�����+����=�Ep?���Irl�>�4���M�?��=��*?e:�>��;���<�E>|�?���=w�H�:_ĿB"��/�׾�(�?���?V �ix?~E�?�n$?'�(�� �Q���Zr)��<����C?��S>g�ݾ9�2�?
B�A���-O ?�UV?��M��#1�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�"�>T�?���=`d�>9�=$簾�T.��D#>��=]_?��?\�M?�A�>L�=�9��$/��TF��HR��.���C���>��a?uL?~Cb>�︽�1��� ���ͽ�p1�Pb�FG@�"_-���߽5>D>>�>P�D��
Ӿ�O3?��̦�S����E�1�?�FC>�.(?p���k���X�䫀?2�f>?k6�����G���C�c�k�?1�?���>�ޱ�1H>��C>"�==�޼�V=Tb��ʓ��<�=d�s?�2�ӯ��ԃ�\ۂ>�þ?uL@@��?��j�D�
?�r������}�r��}�D���=<�:?0����q>3�>:�=�'w�-��6u��=�>�Ư?���?��>�i?�k�|<�<�5=*��>��d?L?*��#���I>�2	?Z��᏿����?d?&�
@@/@��_?�᣿��ܿ\��ھ'վb �=h\<�Km;>:����>.�=��H=�0��I=A~>dY>�#>Z�>�;1>��>5�����ԛ�I�����A��,�cL���Ž0�澇7<����f8�@p��  �=aKl�<ǣ�^n����Z�pv;���=]�U?��Q?��o?A��>M7v��>c%��cH�<�$�4��=0Ӆ>2?!�K?��)?P��=E����d�憁�xk��������>��G>�5�>=��>�Ů>��:"dG>�=>�*�>� >Ć=��L�=�UP>F[�>v7�>���>@{l>�P>�L��J
��k�,�T0���/����?~#վw�5�@	����*�����{{;�A?-�>	C���ٿ�o����U?h���c�2�O$�OM^>NG?�vZ?�j>5��v��=��{=H�˾������=�TҽR�_�E�5��B >� ?�f>@u>U�3��d8���P�Q{���g|>x26?b鶾�G9��u�^�H�}cݾ�DM>�¾>HED��k�W�����ui�R�{=:x:?��?�;���᰾̭u��B��KQR>�9\>Y=Ul�=yVM>YXc���ƽ(H��i.=]��=��^>V#?�*>��='�>$���"�M����>�)C>�D+>�@?�[%?�������G,��v>��>�q�>�<>k�I���=���>z{a>6@�D����x��?��UV>�z���]�cq�au=�ؘ��3�=h��=�; �Ug=���'=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�k�>9z�\�������u���#=��>:H?;Y����O��>� w
?�?�a�M�����ȿ�~v����>�?@��?��m��?���@�Uy�>e��?�gY?ti>e۾snZ�ޑ�>z�@?�R?��>�9�6�'���?H�?���?U��>���?��?��?O��=��%�v�ʿ�@��C�?����([����~>����!��&@��}��ZuI��~P�h~�>5m�<�X?��^�lN$���)>d��<Td�������.�>�s�>TV�>�BE>W#?La?s�^>�c����=��&��YI���K?���?0��1/n��L�<O��=9�^�� ?FL4?��[���Ͼ6ը>`�\?���?,�Z?;Q�>���)>���迿^��p��<��K>76�>�=�>���/YK>�Ծ�ND�*m�>Η>�C��8ھ�,������G�>�a!?_��>���=�� ?�#?�j>��>q0E�_G��4AF�=Z�>�q�>��?J�}?h:?.�����3�����ʡ���[� ^L>Gzy?.?/��>ċ��>����X)��DD����em�?�g?�F�;?E3�?{4??�,A?[�f>���ݟ׾Y���'��>��!?��A��K&���&?�P?!��>�9����ս.�ռ���jz����?�(\?�?&?6���)a�j�¾�7�<
�"�\V�d��;L�D���>i�>9�����=�>�۰=�Mm�8H6��f<\e�=�>���=417��|��� 2?�)=u����;J<"�����j�]�{>mAY>޽�VC?{�-� _�������������n�?R��?�{�?�+���p�4,9?�A�?���>�?0򐾂^���$� 5~�&}������}ܼ@�>Ws�=BFᾼ���:��x���� ���ڽ��?�а>H5�>�S?��<>P��>����a�+�֠'�����k�l'0�wV?���/�Ά"�hw���������ʾ�܆�HǼ>;@Žs&r>��/?cv`>E��>��
??~���O>߱�>�P^>���>H��>E<>&=�����-��KR?�����'�y������f3B?�qd?M1�>Yi�6��������?���?Qs�?0=v>h��,+��n?�>�>D��Rq
?pT:=�9�i:�<V��s��3��[�3��>�D׽� :��M�2nf�rj
?�/?�����̾�;׽�N~��)�=�bc?��J?EQ#���q�r����ڎ��2��S�[�Ͼ�p^�t[�f�!���%��N5���ZY���>�4?U�?͉5�s���0���Iq��q��c >�?�N�>l5�=%�?b��m��87�ǟ�ܸz��́>�}?�i�>sXL?ئ_?�Zt?xe�?���>=?����`�>X>��>��)?:�6?F?��B?��;?��I?�s�>ω[�RD�@V��s�'?5��>�?�r
?��?����V)��3��K�=���,>y�=C�>PHZ�~���x�>o=�=wM?Ȧ�{�8�����	�j>ۅ7?,��>���>V��� ��$`�<��>�
?VR�>�����jr�:S��]�>��?��G=�)>A��=�cߺ=L�=������=����q:�|� <-�=��=tz��Q��-��:��{;z��<�u�>y�?���>C�>�?���� �T���h�=�Y>� S>m>�Dپ ~��j$����g�7ay>�w�?�z�?Y�f=a�=y��=|���R�����#���h�<(�?+I#?sVT?3��?��=?�k#??�>O+��M��X^��3����?v!,?��>�����ʾ��Չ3�ם?e[?�<a����;)���¾��Խʱ>�[/�k/~����>D�����_��6��?쿝?dA�R�6��x�ٿ���[��x�C?"�>Y�>��>V�)�z�g�o%��1;>���>jR?>$�>B�O?#8{?��[?�{T>ܕ8�b-���ҙ�'o1�h�!>q@?��?U�?�y?�l�>8�>��)����^�������Nւ�W=h�Y>���>l*�>��>���=��ǽ+^��V�>����=ɔb>Е�>s��>\��>��w>�9�<*Z?i�?�����5�\GH�f��	mz�^nD?��?��?��7<���4�z�԰���>���?�?��?���A�	>��׽�`��T�O=���>��>k8�> >��=6&�=T�>R��>�`���'���#�am�x�?�6?@�w>�ƿ�q��.q��2QZ<�����d�5����Z���=}���o���i����Z�&Y���z�����X�����{�.��>5*�=vp�=q��=�c�<�x˼;�<�'K=A�<�/=��p���e<� :��dԻ�䉽� ��X<��I=r=����Ⱦp�}?o?I?�	+?aA?!�z>[>i2@�zM�>�w���d?��Q>!�V�󂽾">����C�����پb�۾L�b���>� ^���>�,2>��=���<7�=1�g=���=�:��=���=A7�=��=��=z>�a>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?~�>>�2������yb��-?���?�T�?>�?Ati��d�>M���㎽�q�=F����=2>o��=w�2�U��>��J>���K��H����4�?��@��??�ዿТϿ7a/>��7>�&>w�R�E�1� �\���b��xZ�՚!?�H;��J̾6�>��=Q+߾�ƾN�.=ք6>T_b=Th�pV\���=��z���;=-�k=0Չ>s�C>�x�=.���=¥I=���=��O>�v����7��(,�Q�3=���=�b>&>!��>�?uZ0?G)d?_�>b�m��Ͼ�<���g�>���=�-�><��=qOB>T��>�7?1�D?2�K?�k�>�v�="�>��> �,�$�m�9.�ٱ��$]�<���?�ӆ?�M�>�U<I�A�T��VA>���ý��?�K1?w?k��>�^� ӿ�w(�y�Z���׾;[w�8w=e�鼵�=�%Xɽ��<{DM=�zM>�h?��>i�j>bM�>��n=��=���>��>^ݖ=��>�%D;���=4�ü�<~<K�o���ӽ`���=��=���~�/��S����=�Gw<���+>���>蔶=��;>��>׺	���>М�p�U.��|��ŕt�J��>z��b�O�`�+��]>��>���=)�����>�D>�~�=��?`��?@�>�-�A*�����4����@�t^�=bC�>"�<��L�艇��zc�2�˾Z��>g�>�>��l>�	,�#&?�8\w=��W5�0��>和�_��@@�@q��?��b����i��L�J�D?�C��	��=I~?��I?��?���>�H���ؾ_W0>E��6=g��4q�Ȏ����?�'?���>~��D��J̾�I���շ>�3I���O��ŕ�&�0�^*��﷾��>Dݪ��о�3�b^��������B��r����>A�O?���?B(b�j���xO�.��qB��Gf?�g?9�>�<?�?�Ġ�*��Ϣ�����=��n?s��?�*�?>t�=�X�)J?RI?sF�?&��?��{?̦����>|�N=�b>�5޽od>6�F>��/>;�/>(#�>+�?W>�> �����$����]�Wv��:=g�0=�Y�>`l8>N&>��=���<��=�a(>ߵ�>�L�>4�L>���>��>瞄�L��	?wq����>g#;? v�>W��<%���l�Ɓ��~�M�3桾-�񽋒�x��'D%�O46>ӮU=ѻ�>uͿ��?��>z�$�~(?x4����	���)>�Р>�H���>
��>(�>��g>��>�y�=��><RR>EӾ{1>�V��� �<uB���R�cwԾ!ur>N�$�K�h��(�G��9�����+j�P>���=�6g�<΋�?�a���m��++������?�Ψ>Xi7?��������D>���>'��>>�������e���r�྽��?�]�?�;c>�>P�W?�?��1�N3��uZ��u�.(A�?e���`�T፿ߜ���
��	��F�_?y�x?*xA?D.�<*:z>*��?n�%�3ԏ�w(�>�/�w&;��@<=�+�>P)��O�`���ӾB�þ:6�JF>��o?%�?'Y?�TV�c��=	K��{1?��#?i��> BJ?!\=?X�>1��>�V�>��U?��e>�N?�'?�/?x�g=��="'�>�{=h�v��OU�\y�Ԍ��7��g�9�^�=?W�=��=.gW�*ñ�^½Y4B����;����-���V�=��L��`}=>�>��^?.�>.Xt>�+8?����&9�jE��Ğ8?�H�=��x����+��<1�:E>��r?d=�?yV?1pS>FB��GC��#>�]�>Q6>�JM>�ݼ>�k��^/O�H��<ە&>��.>XS�=hܐ�r��Ob����k�=�b.>���>C1|>���r�'>�|���0z���d>��Q��̺���S���G���1�|�v�?Y�>��K?J�?U��=y_�J/��`If�0)? ^<?�NM?��?"�=�۾[�9��J��>���>�X�< �������#����:�m�:O�s>�1���7��� b>M���gԾFW��B�����|���n#��A=���쒬�ߓw����=h��=����M.#��k�����/�H?�o�=_*��Z��ٛ��Q>%X�>$^�>}�ý�.＃�;��R���1|=PԹ>�ݼ=���b��D�����߄>�A?�g^?�B~?$U��n�Y�d)D�'�������~sμZm?z�>GE�>�!>˹�=rǲ�X�)h� B���>���>8��rI�zО�M��� ��ڗ>�^ ?�C�>��?B�W?��?�%d?n"?�?�ς>�P��hī��A&?.��?R�=��Խ6�T�K 9�MF�i��>Y�)?
�B�繗>=�?��?��&?��Q?Ե?�>� ��C@�ٔ�>]Y�>��W��b���_>��J?�>u=Y?�ԃ?��=>W�5��颾�թ��V�=�>��2?�5#?H�?���>�t�>��d�=���>��b?�-�?��o?I�=�?42>���>�K�=!��>�b�>�?l6O?��s?��J?ˍ�>|܎<_������Z�r��,R�i%};T�G<��y=k�b_t���wc�<�M�;�~����}�N���D��Ꮌ*��;fg�>d�s>������0>�ž>���A>e̟����#�����:��/�=._�>+�?h��>~)#�ϒ=k�>��>���;(?/�?�9?�+;µb��ھgL����>O�A?)��=.�l�P|��F�u�_�f=��m?��^?�W�G��r-r?Y�2?���B^�M	����ƽ!��?S�=?��>%��>��?�3�?UJ ?;,��H������Ja����:�yr=59r>o
羶�3���>��E?+ ?f�>�Q>��0�����c��J/?1֙?���?B��?ZϏ>��Q�0��!������KSV?,#�>�¢�p. ?�^�A�9���^���K߾Y�����I1��������O����"����=�)?@zv?2h?��i?�Y��f���U�����c��H���PV7�XbA��-�j��?
�۾{r���t=�f���I3��F�?�?T��"��>����#D��8��H{>���Y�����<6C�!r=�=�:��?�fP���y(?W��>W�>,�1?�K�Ʉ:�<�$�؈;�s���\=>�N�>���>b��>��=}H����빾鐾(�q�u>�Ec?$�K?�7n?�R�T�/����o�!�S�4��'��T�D>��	>ES�>C�Y��/�|W&��w>���r�d��P���E�	�6�=��1?�g�>��>��?�?x�	��ɬ��w�q�0�ة~<gݺ>-i?-��>#ą>:�ֽ{� ���>��k?G �>�Ǡ>\��������{��G���<�>~��>W� ?�_>tn7��I^��Jy��VG8�ћ�=h�d?|��pa��`�>�#G?������<�>�>��D�"��F�IT	�>��?���=��M>Doƾ68�?���X�2)??����-�*�U|~>E6"?e0�>8s�>��?P��>Ξþ�>�zs?��^?�KJ?^8A?��>V=Yc����ǽ��'�ܒ.=���>O+Z>�Op=���=����"\�L!�<�E=�S�=��̼����j�<A���!�J<���<s�3>��ܿ�1I�!Ѿ"�
���߾={���x�B���M��sת�� ��I~��I��%��OT�eVo������_� 4�?kM�?�v}��u�O3��ѧ~����L�>Ȉ��W�����ͽ����&�Ӿ�~��Wo �~�O��g�M�c�6�'?�����ǿ�����;ܾy! ?@ ?��y?��h�"��8�� >5�<M3��a��[�����οA���y�^?e��>�
��>����>���>�X>DIq>����䞾�{�<{�?�-?[��>�r�O�ɿ����Φ�<���?��@0}A?D�(��쾅OV=b��>"�	?w�?>�W1�E�����I�>�8�?���?�>M=��W��}	�v�e?��<�F�Y$޻k.�=>�=Y='��|�J>�S�>|�SA��Bܽ��4>
܅>��"�'��̇^�)�<��]>��սC,��o=�?�8�����K,�U>���Ң<��'?�\*?��&>�G�>9M���˿oB/�mv?'�@I��?���>�پ��?��۾!�h?4sL?[�&>,a���e�a�*>XԀ��B��_�z�Q�/�=ѱ�>��o> 2*��� ��O_��s�=��>��֬�� h�H�DZ�=Qٿ:�l��s��S���_���H�6�(����+=�.�=e=>��D>5-X>�qo>_e?|ч?;��>�N�>R�1=���ٖ���F�Qؾl�Z�;�n��_�<^�����R�پ$��}�+����P4þ=�E�=F3R�-���� ���b���F�B�.?4_$>��ʾ=�M��&-<�rʾ�������	ͥ�k.̾L�1� n��ʟ?��A?����'�V����*C��{��{�W?�W���x鬾ߩ�=�ڱ��Y=	�>xw�=��⾒!3�@S��`0?�P?^7���Ð�R+)>09�`=,?>�?t@<��>��$?��)�+|�5b[>�i2>��>0Z�><>����۽N�?[�T?���E��rב>���̀{�H�Y=4<	>~�5�F����X>}�<������H�]y���Z�<SY?#�>�*�D��X4��`���Z=�=n?�T?���>�)q?e�K?��=���{V�`�"w<z[Q?C�o?�E>�َ���Ծz ��;r5?ob?&h>�=|��'پK�,�?��� ?�Wo?m�?�z��Y�u�r䍿x���O5?z9w?��k�O,����
���\�6�>]��>���>k2��ʵ>��1?����ړ�����[:��4�?��@��?|�(������m�.	�>���>)�&�c���AD��Ц��B=g��>�����?������N�V�N?��?@��>������
���=�ٕ��Z�?i�?����VKg<���l�o��,y�<�ͫ=��_H"�����7�j�ƾ{�
����⿼٥�>.Z@�V��*�>�C8�P6��SϿ'��h\о�Sq�j�?T��>�Ƚ���'�j�\Pu��G���H�Υ��tH�>��>�I�����{�\(;�����>;����>�hS����:�����1<��>���>l�>����۽�A��?�]��G4ο����ӗ��X?�T�?j�?vn?��P< �v�e�z�:��6G?�Us?�Z?uT&���\�s6�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�e�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�d�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�F�c?cr�1�� 1)��o���>+�B�(���x꼧f-�_��$���x��v"�?eU @�_�?���(�u0?P �>�ā�lܢ���v<��@>��>u�_>K$T�&˚>=�#�V�A��'z=~��?���?<�?���$����=t��?�[�>(�|?	��=�?�N�=Q�ľ*�/>̓}>��N>I^6��y�>�{.?7_�>Ġ�=ג.�W.�"!9�~�s�c�$�F��>>h?d�Z?��>5A�<m��=v2�7.�N�h�I~�=4O�]!&�9����i=��=��<>�j�F�����?Mp�9�ؿ j��*p'��54?/��>�?����t�����;_?Nz�>�6� ,���%���B�`��?�G�??�?��׾�R̼�><�>�I�>>�Խ����\�����7>1�B?[��D��u�o�z�>���?
�@�ծ?ki�N�?������G�}��iT�C���l�#>7'3?ľ��k>[�>q�>>�'|�,����l����>À�?���?���>j�t?QA���Z����=7��>�ф?�� ?���������>���>�Y�oUU�i|����e?��@��@�pG?�i��p���Т��V¾�lо��=�s=��b>y��<��=	Z=���<w5�r%>$�y>)L�>�g�>�{>VX>�z_>�ق���"�AӜ��c���'�˾����ƣ�٬ھQf*�.��`>��ZU���a�������?�;�'��	������<�=Gsa?q�I?讁?�]?/]�[��>Aʸ��D>��W�1�1>�6d>OcO?�R?���>�B5�&"~�d�Y��,}�����Y.E�zv�>9.�>���>*!�>���>�����G>��>�ƈ>B�=>B]@>2�p>���=�>�S�>�T?&�>�G<>Pk>#ƴ��-��a�h�.�v�I�˽���?����m�J�1���U�������8�=�b.?�>����<п��o.H?�����#�y+���>Ŷ0?mfW?��>�$����T��->����j�e|>�P ��ul��)��.Q>�f?j�m>@�%>�����K��&������t>�G?��뾯���O����Q\�=��i��=�� ?��>��� ���AY�W0i����<�%+?H�?|�����0ua�b�c��q(>��>��>@Ƶ=��S>񰽽�J��W��ų�=m��=�I�=N?��+>3�=���>�L���O��j�>�B>��+>��??� %?���)P��қ��M�-�w>�,�>��>�>�(J����=\�>l3b>���[��0��A�?�pW>$�|�9_� �u���x=�{����=���=,a �;�<�=�%=e�~?߀���房��q��WD?�#?̝�=�nH<��"�=����g��O��?B�@�s�?6d	�y�V�~�?�F�?�7����=V��>Dë>�;�L���?�ƽ�ޢ���	�P9#�`K�?�?0�ȋ��l��8>Ib%?֯Ӿ�p�>�o��X�����W�u��#=E��>!1H?�D���N��=�`
?�?�b�Ω��M�ȿ�v����>z�?��?.�m��@��b@��}�>���?JkY?�[i>�X۾NjZ�၌>�@?�
R?&�>95��'���?3׶?��? G>�x�?��r?}�>�!��ҷ&��|��0����W=�2)�;m�>9�=U�ž H�������+�j�����\>R�-=l��>k{ԽY����Ц=[N��uO�����J�>��>�lE>�E�>���>���>嫝>�J=,���aB���3���FP?W�?N��{WP��ǽr����n%-?��K?�|F�B�׾l��>�h?o��?��E?\�>�$������Yÿ��;T�=���>.c)?a�>�rp�Q#u>p�Ⱦ�����>�D�>m3!����E'׾:�4=^;�>[�?֚X>"�>�1+?��?L�>� 8>�L\��χ���C���>��>��Y?��?*�1?BȒ�tD+�9����_��z|���C>��?J,?۱d>�u��53��0�t��]��D)�=�HH?[{?��<!?�9�?[�U?�#?yp��ʾվI��8��>J?6�1�Jd.�!6(�:��B�?-��>�Z�>�ƽH��)���B(�������>�o\?�� ?�����e�i��j1=����>|�<5o�=�ȣ���->j�D>�م�Z?I=.�>5N�=�v��GZ#�a�/=G4�<�}>��=�=��<�+?��D<���ˮ]>��\�,�a��=�r�=�(��Ѳ6?���W�v������������<�?�R�?�Ţ?�H�N�f�WYG?�&�?���>C�>
vO�a4Ǿ�G���������#\���4�=�ҟ>b��,���!����\��?�v���*�i� �H�>� �>hp�>��>���>��F>¾Ͼ/���
��U��o�X��#�J�����P%�D뻾�C���3�"������2M�>�\_�~%v>x�?ߎ4>DĲ>s_�>xN->uq�>)�>�">'�>hB�>�>>|Z�	Ղ��KŽ6(U?�9���&��𾧂��v�??;La?��?���<I/���B	�J�?��?�՞?R�d>�!i�ڝ+�Պ�> S�>�ǁ�z
?)h=� �=���<�ѾR�+����;F�W��j>G.�MF�ANN��*Q��_?4?��M��$˾X_!�F�-�=mNx?��N>E�⽖�1�VɊ�׶y�j��#�^>s!��e����f��qc�����le�1V��Rd0���� �9?og=?\~%�GX.�-�f�(�M�,�-��a�>��?k��>� -=G��\��I6��}h�/���~�p��>w�|?�H�>7�I?��;?��P?�L?���>�^�>	x�����>��;Pf�>Yt�>��9?k�-?��/?l?*�*?`>�q�����N{׾]2?.�??�)?y�?����ýβ��EU�11x��>}�ZY�=qS�<�ٽFWq�}q\=l>T>CX?֛�"�8�����;k>��7?�}�>m��>����-�����<�	�>u�
?�C�>����1|r�jb�oQ�>���?����c=��)>��=����Ϻ�_�=���*�=�0��[x;�?�<?��=���=N�u�b������:�Ƈ;Bk�<M� ?ZJ?Je>�N�>�R|���ﾙ���N=B"d>�)>��=�?�:��������j�]��>:�?��?���<���=�>s������Lb��������<kv�>�?3�C?6T�?�T8?��?�a�=��
��4���6��������?" ,?���>���)�ʾ�먿��3���?�d?� a�a��'.)�Ƈ¾y�ԽE�>�O/�['~�� ��+D�尌�����n��9��?��?y@�Z�6��8辮���>l��wC?d:�>p=�>���>��)���g�L��?;>1u�>R?W#�>i�O?�<{?~�[?�fT>�8�1���ә��M3���!>J@?���?��?|y?5t�>��>_�)�Z�eT�����3�8���SW=�Z>*��> (�>$�>���=��ǽ�Z��^�>�ra�=M�b>���>C��>��>��w>K�<.IH?t�>�ľ�Cτ�V�⾪R�Y-?�̆?�; ? ���/�-�gY�QfP>ܭ?��?8�I?YYþӳ>�j=ch����$��˼>�	?v�>y�$>��>n��>m�?���>�'�����I���=H�!?�S?_��=�uĿ~�\��\��-����=���X����F��F���}=��z���d�O-���(�����rX����ž���m/���?3��=V�;>i
>=�9Ӥ���+�<��g<3C��(�l=�)���B=���V,; ���t��-<����ݽ�ξ)�z?pjI?��*?ŭB?f��>�44>��N!�>��a�?�\>U�Լ�+��R�5��u���̓�k�;�mϾ��U�Շ�����=I!�<��=�-%>���=/�<�ں=��N=]n=�w��f��<�G�=�$�=��=9 �=*D&>`>�}?������B�M�5L=x�?<V�=o�>�w���5?'�>Gpn�08���x�o�p?�g�?��?�,?�����`�>�m�������G>�o����=Kn=��>G�>�SY=N��g�� =��?m�@o*?[��
"ֿ���>k�7>��=1�L��l4�TG���S���W�i$?��:��bо�m> ��=�ྀ^ɾ�=�A>UmQ=<6���W�ѕ�=z_��:�v=^��=멇>̾c>B��=:���~�=�=�>��E>���;�G�Y�e��y�<�]�=I\c>�s>*��>��?e60?�[d?%�>Ao�nqϾ~���3�>��=�K�>��=LB>u6�>q�7?P�D?&L?���>L��=�	�>��>�,��m��.�����m�<���?�׆?W4�> �S<L=A��l�Ue>���ƽ�?GZ1?{?#˞>p����(&���4���j����;�2=��3��FҼ�����Bܽ�m��">���>�o�>���>�Nn>�K>��a>�`�>l�=(��<P-=��y��<�;S�e����<����pO�<�2;�:�<��X=�y^��m伳�l<�,=�/�<�(6<�>�`�>��
>��>Pޮ=ҏ^��
�=,%Ծ��9�*[���}���8C��uY�󃿂z4��ZQ��z>S�>��������P>?uզ>~΢���?h�z?=i >��d�#g�L��װ=�mB�$o�<��=F�\(m������k��������>��>��>��l>�
,�8?���w=�⾨`5�]�>.w��&��/��:q��>������i���Ѻ(�D?�E�����=#~?h�I?)��?���>���I�ؾ�00>$E���.=/��0q�f�� ?Z'?���>[#��D�m۹�$Ԅ�OL>�߾79�������I���V�O���u��>��о�2����g�5G��)���i�?��֞�t�>��e?@x�?O���$����-��7v�Q���R?D;�?h�>��>��?��>PR��C��:K�=��r?���?�f�?�>�#�=�մ�CH�>Z	?���?���?wvs?c�>�\�>w0�;y� >kǘ�؈�=�c>o�=P��=	V?s{
?a�
?|��	�=��G���X^�V��<��=Yo�>m8�>�ir>0{�=�Af=t!�=;B\>;��>c�>��d>��>*8�>m!��X����!?FLl=N��>=;??�TH>L<�=@���S��"��fPu�(YS�c��."����<#W��eE�^8����>8���]��?m3g>E%��q?'B־1 ��RbE>P0�>��཭~�>��S>3P�>�Ŋ>�B�>���=��>Rs>�����>�-��v� �us=��6��Q��\^>^h��d��a�����&k�"ó�Vv �1�b��.��Ė<�?%�<���?� �Ils���-�������>��>�2?��E��o�=�X">�^?�.�>3�޾Ϋ��� j���?KT�?�N�>��
>�?<w*?�Xa��^��>��9Z��_��<���]�����d���ξF����Z?[t�?�;*?ش��q{>�s@?[��2ú�q>�UX��sm�Ғ���h
?܊����T��0O��bv��<��e? e�?�'?ܜ���A����4?6Z{?c�]?\/9?;'I?l�h?�����!?���>AfG?8� ?�o\?lN?K��>RXB���=�O>�.�>&Խ��q�'�ƽLB��A�<��'=�����گ<}Z���,=�hS<���<�4��|�	~�;#�=�ע<!�>" >���>�lQ?��>z@�>�M1?�3%���:�c��ޒ0?�X=����s���㡾�����z= 
t?�Ѵ?�h?t�#>��F�0�
��P>�#�>O�>�I�>�2�>�7̽�1G���*=��M>�+>v=Kj��������F��B8M=�`5>�i?d�	>�!��H"�����u9����N>>@���IӾZ羊�^��CP��B��'��>؈o?�)=?���<�9�f��=G]��7L?1�W?�?A��?&!L=����V&�'e���νH >x�.=��+��'������5��<��W=^���4٠�_�c>�^�b޾�:n�~+J�����;?=����V=���v�Ծvs~��a�='�>�F���!��&���Ϫ�[yJ?�Ak=8̦�cX�Z)���Q>��>��>t�=���u��@���z�=Ψ�>�9>�ڨ0G����9��>Z]?�Na?��k?���nU��7�6V
�I�������
�>��>-��>y?>��	=�h��VN�-�h���n����>��>f-�N�W��CᾀO侂��Gd�>�?6�>TD?�rG?��?:i]?��=?	�?;��>׼1��m�*?��?9��=�l\�Ir����*�	-C�M�>��5?ĝ��~�>m�
?߸?&?FYN?��?r�E>z����N���>�V>z)^��ӱ��ߢ>��??�'\>W_Q?���?��>v(�np����T��7*>�j>�1@?�_)?�?װ�>s��>&Ɨ��4�>�t ?�,?���?\g?�{>���>��D>}k?OC��x�?l�	?`<?�^0?�e9?-�S?V�>#�;M�뽯H��i4G��4�н��1�:�5�*�ֽ�;�<KV'>g*s�"�ټ��ڻV-�o�μMh�ë=�_�>j�s>+
��f�0>F�ľ�O����@>쇣�%P��$ڊ�9�:�c޷=5��>��?#��>�X#����=/��>I�>6���6(?��?�?k�!;��b���ھ��K���>"	B?T��=��l�����q�u��g=��m?s�^?��W�l&��L�_?>g?���Y�2���K#���6���.?qN?�T�\�>��w?�=n?��>��F���1����h��c���M�=ӡ>�	���V�9wq>�%)?���>��>��1=Tվ=�u������G$?���?Xȵ?���?�� >�+Y�����Ҿ!�����a?9�>����a1?��R=e־�ܦ��þ;������ƾ�d��3�о�KĽD������n��=?|�H?��\?;Q�?����W� �q��ـ��_��ܾr�۩L��%�P/��ʐ��;�Œپ����d<Ɂ���j7�Y��?�'?�1%��1�>���iM����˾z�/>�Μ��+��ڛ=�@W�1*=Ȣ�<y�%qW��幾=H$?��>�
�>��9?�7U���>�Y�<�X�G�����|S>�
�>$ѣ>A1�>7�	�� <�1��Ӿ�������>"�?�?j~Z?��9�ɞ(��[��Ω:���=)e��A���W�=N��>���Vze��'c��q'�Z%s��+K�֮��r��wD�>0}*?1�=�P�>V3�?�x?�uP�9��� ����b+����$>�b?��?�tB>��"�t�ɺ�>B�l?d��>�>�����Z!�0�{�!�ʽ54�>�׭>ǥ�>$�o>ǧ,��"\��k�������9�Q=�=ݢh?������`��߅>8R?��:�zG<F��>�mv�B�!������'�A�>M�? ʪ=?�;>c~ž� �2�{��I��	G)?�:?/���ڀ*�:~>',"?�j�>@6�>q(�?[|�>3þk�V��?��^?�GJ?�SA?�Q�>A)=�����Ƚ�&�,=㊇>2�Z>��l=I��=M����\�����<F=~�=�*μ�y��Ú<>,����K<o��<��3>��տ�>�nּ�����y�ھ�����JS���w��6�����s����r�mԽ��z��(~��`��(�����?�>�?��$��(���������z��-!>`��ŝu������𽿪��zYӾuU��s
"��*T������g� q8?x/z��῍r��5p����?iΪ>�ȃ?�03��ؾ��R�j����^�:5��7� 
��'�߿`�*%h?f�?�����)����>��2=q��>@hY>��u��/W��O��34?��:?4s$?1���<�ɿ�Yɿ>lT�?��@�|A?.�(����V=[��>�	?��?>:W1��G�����$R�><�?���?�M=T�W���	��e?vS<G�F���ݻ5�=G?�=�F=���6�J>�V�>��HWA�n@ܽA�4>hم>�i"�٨��z^���<Ą]>�սwE��5Մ?*{\��f���/��T��U>��T?�*�>b:�=��,?X7H�`}Ͽ�\��*a?�0�?���?&�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=S6�Z���~���&V����=_��>a�>ł,�����O��I��Y��=����f¿L/�2����A��j&��
j�e{q���L��ͽ_W��Wx��f��cc�=��=�v>���>6N>�R2>S�P?$�?m��>��I>��̒���� ���ټ�g2�x�"��j���d�z8ȾGE��m������� ����־��;�H��=�Q�P6�����fd�*�H��+?6�>z�Ⱦ��L��!�<�ɾ�^����ż1���>5Ͼ8�3���m��z�?6�??w뇿�Y�=���S�k���;G^?x���I��+�=��
��
�<���>��=�-�3�2�Z#Q�;?��,?��A�m��>���v�v;`�0?x�"?=U>�{�>��4?�@���޽�<i>�M�>���>���>���=��̾
G���?R�w?�K:���ľt��>�������ΝB�B��=��;"�>�c�>W#���"ܾ�S=�u�����<�(W?/��>��)�m�t`������R==��x?�?�1�> {k?��B?���<�g���S���!xw=k�W?)i?Ҷ>􆁽оK|��z�5?��e?��N>B_h���龽�.��T��%?��n?d_?�����w}�������Qn6?M�|? gC�윿���4վ�6�=���>1	?ʺJ����>��<?���#ә���̿�H��ؙ?��@|��?�w�=X����zK>��)?��>��y����QF�o���� �=f2�>��;����2?*��s�h?���?�?v
s����*o>h����?7�?־2*=�X�׿u��>�������jވ����ݾ-V�9�ɾ�0�.ɾ�:�<]T�>�@�:a�W�?|O��2�3ֿ.��� 0����W�!/�>}��>\$���� l�ԇv�� 8��ch�B$��혣>���>���iԾM�p�?���J�7z�>�cؽ�\�>����> G��&��x]���*>���>>������	��Z�?+@��F�ܿ����(��h�4?�ۏ?���?��%?�s>G�z�_�$�u�O!0?�gz?�:�?[�����+����=�Ep?���Irl�>�4���M�?��=��*?e:�>��;���<�E>|�?���=w�H�:_ĿB"��/�׾�(�?���?V �ix?~E�?�n$?'�(�� �Q���Zr)��<����C?��S>g�ݾ9�2�?
B�A���-O ?�UV?��M��#1�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�"�>T�?���=`d�>9�=$簾�T.��D#>��=]_?��?\�M?�A�>L�=�9��$/��TF��HR��.���C���>��a?uL?~Cb>�︽�1��� ���ͽ�p1�Pb�FG@�"_-���߽5>D>>�>P�D��
Ӿ�O3?��̦�S����E�1�?�FC>�.(?p���k���X�䫀?2�f>?k6�����G���C�c�k�?1�?���>�ޱ�1H>��C>"�==�޼�V=Tb��ʓ��<�=d�s?�2�ӯ��ԃ�\ۂ>�þ?uL@@��?��j�D�
?�r������}�r��}�D���=<�:?0����q>3�>:�=�'w�-��6u��=�>�Ư?���?��>�i?�k�|<�<�5=*��>��d?L?*��#���I>�2	?Z��᏿����?d?&�
@@/@��_?�᣿��ܿ\��ھ'վb �=h\<�Km;>:����>.�=��H=�0��I=A~>dY>�#>Z�>�;1>��>5�����ԛ�I�����A��,�cL���Ž0�澇7<����f8�@p��  �=aKl�<ǣ�^n����Z�pv;���=]�U?��Q?��o?A��>M7v��>c%��cH�<�$�4��=0Ӆ>2?!�K?��)?P��=E����d�憁�xk��������>��G>�5�>=��>�Ů>��:"dG>�=>�*�>� >Ć=��L�=�UP>F[�>v7�>���>@{l>�P>�L��J
��k�,�T0���/����?~#վw�5�@	����*�����{{;�A?-�>	C���ٿ�o����U?h���c�2�O$�OM^>NG?�vZ?�j>5��v��=��{=H�˾������=�TҽR�_�E�5��B >� ?�f>@u>U�3��d8���P�Q{���g|>x26?b鶾�G9��u�^�H�}cݾ�DM>�¾>HED��k�W�����ui�R�{=:x:?��?�;���᰾̭u��B��KQR>�9\>Y=Ul�=yVM>YXc���ƽ(H��i.=]��=��^>V#?�*>��='�>$���"�M����>�)C>�D+>�@?�[%?�������G,��v>��>�q�>�<>k�I���=���>z{a>6@�D����x��?��UV>�z���]�cq�au=�ؘ��3�=h��=�; �Ug=���'=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�k�>9z�\�������u���#=��>:H?;Y����O��>� w
?�?�a�M�����ȿ�~v����>�?@��?��m��?���@�Uy�>e��?�gY?ti>e۾snZ�ޑ�>z�@?�R?��>�9�6�'���?H�?���?U��>���?��?��?O��=��%�v�ʿ�@��C�?����([����~>����!��&@��}��ZuI��~P�h~�>5m�<�X?��^�lN$���)>d��<Td�������.�>�s�>TV�>�BE>W#?La?s�^>�c����=��&��YI���K?���?0��1/n��L�<O��=9�^�� ?FL4?��[���Ͼ6ը>`�\?���?,�Z?;Q�>���)>���迿^��p��<��K>76�>�=�>���/YK>�Ծ�ND�*m�>Η>�C��8ھ�,������G�>�a!?_��>���=�� ?�#?�j>��>q0E�_G��4AF�=Z�>�q�>��?J�}?h:?.�����3�����ʡ���[� ^L>Gzy?.?/��>ċ��>����X)��DD����em�?�g?�F�;?E3�?{4??�,A?[�f>���ݟ׾Y���'��>��!?��A��K&���&?�P?!��>�9����ս.�ռ���jz����?�(\?�?&?6���)a�j�¾�7�<
�"�\V�d��;L�D���>i�>9�����=�>�۰=�Mm�8H6��f<\e�=�>���=417��|��� 2?�)=u����;J<"�����j�]�{>mAY>޽�VC?{�-� _�������������n�?R��?�{�?�+���p�4,9?�A�?���>�?0򐾂^���$� 5~�&}������}ܼ@�>Ws�=BFᾼ���:��x���� ���ڽ��?�а>H5�>�S?��<>P��>����a�+�֠'�����k�l'0�wV?���/�Ά"�hw���������ʾ�܆�HǼ>;@Žs&r>��/?cv`>E��>��
??~���O>߱�>�P^>���>H��>E<>&=�����-��KR?�����'�y������f3B?�qd?M1�>Yi�6��������?���?Qs�?0=v>h��,+��n?�>�>D��Rq
?pT:=�9�i:�<V��s��3��[�3��>�D׽� :��M�2nf�rj
?�/?�����̾�;׽�N~��)�=�bc?��J?EQ#���q�r����ڎ��2��S�[�Ͼ�p^�t[�f�!���%��N5���ZY���>�4?U�?͉5�s���0���Iq��q��c >�?�N�>l5�=%�?b��m��87�ǟ�ܸz��́>�}?�i�>sXL?ئ_?�Zt?xe�?���>=?����`�>X>��>��)?:�6?F?��B?��;?��I?�s�>ω[�RD�@V��s�'?5��>�?�r
?��?����V)��3��K�=���,>y�=C�>PHZ�~���x�>o=�=wM?Ȧ�{�8�����	�j>ۅ7?,��>���>V��� ��$`�<��>�
?VR�>�����jr�:S��]�>��?��G=�)>A��=�cߺ=L�=������=����q:�|� <-�=��=tz��Q��-��:��{;z��<�u�>y�?���>C�>�?���� �T���h�=�Y>� S>m>�Dپ ~��j$����g�7ay>�w�?�z�?Y�f=a�=y��=|���R�����#���h�<(�?+I#?sVT?3��?��=?�k#??�>O+��M��X^��3����?v!,?��>�����ʾ��Չ3�ם?e[?�<a����;)���¾��Խʱ>�[/�k/~����>D�����_��6��?쿝?dA�R�6��x�ٿ���[��x�C?"�>Y�>��>V�)�z�g�o%��1;>���>jR?>$�>B�O?#8{?��[?�{T>ܕ8�b-���ҙ�'o1�h�!>q@?��?U�?�y?�l�>8�>��)����^�������Nւ�W=h�Y>���>l*�>��>���=��ǽ+^��V�>����=ɔb>Е�>s��>\��>��w>�9�<*Z?i�?�����5�\GH�f��	mz�^nD?��?��?��7<���4�z�԰���>���?�?��?���A�	>��׽�`��T�O=���>��>k8�> >��=6&�=T�>R��>�`���'���#�am�x�?�6?@�w>�ƿ�q��.q��2QZ<�����d�5����Z���=}���o���i����Z�&Y���z�����X�����{�.��>5*�=vp�=q��=�c�<�x˼;�<�'K=A�<�/=��p���e<� :��dԻ�䉽� ��X<��I=r=����Ⱦp�}?o?I?�	+?aA?!�z>[>i2@�zM�>�w���d?��Q>!�V�󂽾">����C�����پb�۾L�b���>� ^���>�,2>��=���<7�=1�g=���=�:��=���=A7�=��=��=z>�a>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?~�>>�2������yb��-?���?�T�?>�?Ati��d�>M���㎽�q�=F����=2>o��=w�2�U��>��J>���K��H����4�?��@��??�ዿТϿ7a/>��7>�&>w�R�E�1� �\���b��xZ�՚!?�H;��J̾6�>��=Q+߾�ƾN�.=ք6>T_b=Th�pV\���=��z���;=-�k=0Չ>s�C>�x�=.���=¥I=���=��O>�v����7��(,�Q�3=���=�b>&>!��>�?uZ0?G)d?_�>b�m��Ͼ�<���g�>���=�-�><��=qOB>T��>�7?1�D?2�K?�k�>�v�="�>��> �,�$�m�9.�ٱ��$]�<���?�ӆ?�M�>�U<I�A�T��VA>���ý��?�K1?w?k��>�^� ӿ�w(�y�Z���׾;[w�8w=e�鼵�=�%Xɽ��<{DM=�zM>�h?��>i�j>bM�>��n=��=���>��>^ݖ=��>�%D;���=4�ü�<~<K�o���ӽ`���=��=���~�/��S����=�Gw<���+>���>蔶=��;>��>׺	���>М�p�U.��|��ŕt�J��>z��b�O�`�+��]>��>���=)�����>�D>�~�=��?`��?@�>�-�A*�����4����@�t^�=bC�>"�<��L�艇��zc�2�˾Z��>g�>�>��l>�	,�#&?�8\w=��W5�0��>和�_��@@�@q��?��b����i��L�J�D?�C��	��=I~?��I?��?���>�H���ؾ_W0>E��6=g��4q�Ȏ����?�'?���>~��D��J̾�I���շ>�3I���O��ŕ�&�0�^*��﷾��>Dݪ��о�3�b^��������B��r����>A�O?���?B(b�j���xO�.��qB��Gf?�g?9�>�<?�?�Ġ�*��Ϣ�����=��n?s��?�*�?>t�=�X�)J?RI?sF�?&��?��{?̦����>|�N=�b>�5޽od>6�F>��/>;�/>(#�>+�?W>�> �����$����]�Wv��:=g�0=�Y�>`l8>N&>��=���<��=�a(>ߵ�>�L�>4�L>���>��>瞄�L��	?wq����>g#;? v�>W��<%���l�Ɓ��~�M�3桾-�񽋒�x��'D%�O46>ӮU=ѻ�>uͿ��?��>z�$�~(?x4����	���)>�Р>�H���>
��>(�>��g>��>�y�=��><RR>EӾ{1>�V��� �<uB���R�cwԾ!ur>N�$�K�h��(�G��9�����+j�P>���=�6g�<΋�?�a���m��++������?�Ψ>Xi7?��������D>���>'��>>�������e���r�྽��?�]�?�;c>�>P�W?�?��1�N3��uZ��u�.(A�?e���`�T፿ߜ���
��	��F�_?y�x?*xA?D.�<*:z>*��?n�%�3ԏ�w(�>�/�w&;��@<=�+�>P)��O�`���ӾB�þ:6�JF>��o?%�?'Y?�TV�c��=	K��{1?��#?i��> BJ?!\=?X�>1��>�V�>��U?��e>�N?�'?�/?x�g=��="'�>�{=h�v��OU�\y�Ԍ��7��g�9�^�=?W�=��=.gW�*ñ�^½Y4B����;����-���V�=��L��`}=>�>��^?.�>.Xt>�+8?����&9�jE��Ğ8?�H�=��x����+��<1�:E>��r?d=�?yV?1pS>FB��GC��#>�]�>Q6>�JM>�ݼ>�k��^/O�H��<ە&>��.>XS�=hܐ�r��Ob����k�=�b.>���>C1|>���r�'>�|���0z���d>��Q��̺���S���G���1�|�v�?Y�>��K?J�?U��=y_�J/��`If�0)? ^<?�NM?��?"�=�۾[�9��J��>���>�X�< �������#����:�m�:O�s>�1�����(b>����m޾��n�7#J�@�羚oL=
k��+V=�(�վJF��{�=(
>̰���� ����hЪ�S5J?k=�E��|�U�z����>��>��>4�9�jw��y@�&����і=֏�>��:>n ����FdG�'��?�>�OE?�V_?�j�?� ��s�%�B�����wg��+�Ǽ�?�w�>�i?�B>$��=]���H���d�tG���>���>�����G��;���/��h�$�捊>9?^�>��?j�R?��
?��`?0*?�D?$�>
��a���;B&?���?��=��ԽW�T�� 9�,F����>ـ)?ֶB�=��>E�?�?_�&?�Q?\�?F�>\� ��A@�Y��><Y�>��W�eb����_>ݫJ?���>0>Y?�ԃ?��=>��5�'좾�ީ��Y�=�>��2?�4#?��?�>0��>T���s��=R��>�c?�0�?s�o?���=��?�:2> ��>q��=���>u��>�?�WO?�s?7�J?ԑ�>���<?5���8��gEs���O��m�;�vH<H�y=��I+t� K���<�;�t���L��E���D��됼�0�;�m�>��q>��mf >^5����4���'>��<f�w��
������Ї��f�>;?"<�>A��B�=���>6��>)��[�*?۝�>V?JG =d�y6�m� 3�>�xE?��=C�c��`��y�w�={w=��^?(K?��J&ž*+c?s�H? ��H�<����|�ڽ[�U�$v?��>�聾9�>,�~?[dO?��>+���!ҁ�}����o��=���Ħ=��>G�#��]W�G��>��+?�ߢ>w}J>�����|�I�U�+�����>�n�?Ӂ�?O�?l|�=0-���^�(���hD��^^?��>G<����"?=<��ϾVF��x)��?�8���#���?��n��Й$��ꃾ�U׽�ż=��?�s?_q?�_?� �sd��%^�����^V��'��#���E�'E��C�e�n�(^��$������ H=�#�_�&�A.�?�?	ԽK]�>���k2#����5D>^��Bׯ<�P�>-�=��=��M��؋�V<�!�����,?B�=�T?.nh? BK� �<��2�(ZN�!�9���<>���>pL�>�F?R܄=Mm��j�;���i�`�	��8v>$xc?�K?"�n?�l�+1�ㆂ� �!���/��c��G�B>Kh>���>�W�����8&��X>��r����+w����	�d�~=�2?/'�>粜> P�?D?-{	��k��nx���1�^y�<�-�>�i?�>�>��>��Ͻ�� ����>~�l?m��>�ޞ>��0� �g�{�~�̽j�>~�>(��>s�o>�\*�6�Z��	��fÎ�n�7����=��h?����Fb��ڇ>�9Q?3QF;@�:<��>�j���!�ˊ�[)���
>6�?|�=dM=>�4ľ��P|�VQ���)?�N?�A���l*�o5>A�!?���>��>���?7�>�?ľ�����?��^?�J?��@?pb�>d�-=@{��X�ɽ��%��-=fІ>_CY>j�b=���==8�6�\��(�F�G=&u�=BӼ/ ����;<q��ݼ=<��=n�5>�ۿ�J�)Y־;��Eo�[��t���<��5����Z������V�z�ї�
�-��-U�_�h��쏾{�p����?���?�#���ލ��왿����������>�id�5z��Wb��D��Iw��*S��Ʈ������P�q"f�v(c�H�'?�����ǿ鰡��:ܾ5! ?�A ?$�y?��2�"�8��� >�C�<�)��j�뾧�����οߦ����^?w��>��/��e��>ѥ�>��X>�Hq>����螾P4�<��?!�-?	��>�r�&�ɿ^������<���?*�@F�A?O(���x�K=Ұ�>�#?7B>�-��]�hl��]>�>t*�?���?y�S=ȓW�Ľ��c?�1<�%G��o���l�=k��=��=���]K>��>;&��?�Q1޽�f5>��>p�L�n�a�O|�<V^a>�Jٽ����'Մ?�z\��f��/��T���U>��T?�+�>�:�=n�,?7H�c}Ͽ��\��*a?�0�?Ħ�?�(?�ۿ��ٚ>s�ܾ��M?�D6?���>>d&���t��|�=FM�LD����&V�c��=ة�>܀>,�����O�xS��A��=T��ƿ��$�
�H�<�/����X���U���|Q��ߟ�p�>~��sg=��=y�P>3�>S�T>��X>�NW?f�k?/�>�F>��ub���.;r�$��� �G~��*������쾫�߾!3	�-�����ɾ� =���=�4R�ӗ��F� ���b��F���.?�z$>��ʾa�M�Y�-<�nʾ$��������諒�-̾~�1��n��̟?X�A?����+�V�f��ew�����z�W?�O����謾��=���9�=e#�>���=@���3�_}S�n+?��?d�Ͼ).���>x�v���+=��$?l��>;R>8J�>��?
��=(�Zx�=w�f>CN�>n��>�t<�����̽%�?��K?���Î�k�>�澩�e����=�C�=߽���<tSF>�$�����E�	=����ck=7X?�+�>�C�����ľ�CQ����=?w�?p?�^�>��l?oD?+C�<_��f�4A��j�<��K?�hj?|_>�ǽj���W��&k(?0Xk?� h>���9$��7xL�����Q?�h?�+?4�⢃����P!�O>?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?o�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�ٕ��Z�?y�?Y���=@g<{���l��n���}�<FΫ=���G"�����7�@�ƾ��
�����࿼���><Z@�T�h*�>�C8�K6�TϿ-��:\оUSq�U�?a��>I�Ƚ뛣�D�j��Pu�,�G� �H��������>u�=��<����	��c�;�4�>)bS>q��=\g�> C��{�/�׾9����!�>�?B�>~c���~p���?�	��οՑ���׾���?@ �?�t?͔?�����ǾM������>�g?E�?�[d?����t��!�r=۹j?GS���Y`���4�GAE�U>3?/<�>�-���|=��>�|�>�h>Z/�F�Ŀ�׶�Y���x��?r��?7n꾻��>h��?k+?pm��6���X����*�lX)�>A?92>t�����!��2=��ג���
?�w0?�v��'�32Y?q�i�R�h��悿�o�0 �>��e�FF���\�>ZB���k��3���߶�|ߤ?�	@q��?ѓJ����d�A?�	�>9_�ޫ����>+?�P?y��><U>6~7>g�!�(G,�P�=[��?:Y�?e�%?����O����A�=��e?jѵ>r2�?��=ux�>�1�=����%���0�%>��=T0�ʛ?O�N?�3�>ɤ�=Q;��(-�]�B���Q����h�C����>�a?�RL?��_>q���b3������ͽ��8�d���@�D�1�r�۽bC8>:�9>�>��D���о��?�o��ؿ�i���o'�~54?ָ�>��?�����t�����;_?wz�>�6��+���%���A�a��?�G�?M�?ͻ׾F̼�>r�>}I�>O�Խ4���Ԃ��<�7>ҞB?@�cD���o���>���?��@uծ?si�	?<�I��e~����'7�� �=��7?e�7�z>r��>��=�qv������s�¶>@�?�x�?B��>��l?�|o���B�1=�@�>��k?�u?�tr�K��6�B>"�?�������C��$f?��
@�u@�^?{梿S˿������Ӿ�bU�j�P>쐻�1�>��伆��;Jξ=���� p��b�r�H>C�~>6v�>i�E>nB>#��=��w�i�"�����N��ɺ(��!���[�Lh1�! ��]e�pӾ����*o3�%:g�
  �H�C��;����1�0��=�U?�R?�p?č ?F�x�[�>P���#�=(�#�%�=T2�>�]2?��L?�*?��=����.�d�~^���C��J���w��>KuI>�z�>GC�>�"�>ʼ|9��I>�?>Hv�>�� >�A'=���7=��N>�O�>���>�x�>�s<>�>@ȴ�"-���h�v�v�ei˽��?����|�J����8��)���4ɞ=RM.?�i>�� Cп�����#H?ݔ�!%�ӡ+�Q>�0?FW?q^>�	��N-S�Ҟ>����j��)>�����k��m)��Q>??A'g>�&u>��3��[8�q�P��6��ƽ|>Q6?�ᶾ�"9�^tu�y�H��cݾ��L>���>�Y;��p�����rti��|=�b:?��?����˰�<'v�[}��eR>�]>��=�9�=�M>�e�L�ƽx�F�!�1=���=Z�]>���>DV�><X����>�����>��>)�>���=Տ^?y�C?��\>�S��r!ݾ&�����>���>�H�= �T���g�P>2�>	��>�2ѽ�Q��A_����f�+>�E���Ⱦ
=�Cb<��9�˹E>S�~�w��8"�)-T>7~?�~��f^��d���]ޒ>�v?]� >C[>�@>S�'��읿_˾��?��@��?�jD��At�"89?��?�ؼk�>��>@��>"�Ǿ\X½TX%?�'%�~����׾��8x�?Ȯ?���x:��X(u���V>��?�x��h�>�v�Z��m���u�v�#=#��>69H?(U��4�O��>�w
?�?_�������ȿ�{v����>�?e��?;�m�eA���@���>��?EgY?Jpi>�h۾�eZ�ˊ�>޻@?�R?��>9��'�A�?�ݶ?���?YI>u��?s?^h�>�4x�QY/�=6��]���#u=�b\;w`�>�U>����deF�3ד��h��@�j����B�a>O�$=��>�5�u5���9�=�싽,F����f�Ȥ�>&+q>��I>�X�>h� ?�`�>\��>�n=�c��䀾�����K?���?���An�*ؾ<f �=�|]��?
�3?��E�GYξtݨ>4\?#Z�?�Z?�
�>����U�����fh��p��<�`K>Z�>���>�ሽ}�I>"xվ`�C����>�Ș>�k��$�پ�2��ާ��d�>��!?W��><Q�=��#?p� ?�>�B�>��S�<��\m+��T�>��>��7?�f�?�?_���q@�bp��dܚ�=N���d>R*y?w?Q�c>���8 ��OꂽI�<�5���ن?��X?iJ)�/�?�B�?)�D?��H?܋)>Y/x������8��Vo>�M+?ւǽ�4�ї��A�U�?E?E[?q���!�_�=JX���㾬��>�D?�:?�f�b�u��ܾ�l�:!K�=V<�<�=���=��.>�4J<L���n�.>^�>ƕ�>�|���n�'�۽�Y�=`�?B�>��8��K~�=,?v�G�{ۃ�O�=u�r�xD���>�IL>�����^?{k=���{�����x���	U�� �?��?5k�?���5�h��$=?�?Q	?"�>1K���}޾�ྍPw��~x��w�u�>���>�l�U�;�������|F���Ž�N����>���>h�?n ?�=N>��>N���^M'����r�N^^���� 8��).�=�Yq��1F ���������$�y�{��>܈���>Xj
?Ѵk>�]|>���>
��l��>]�Q>��~>h��>R
U>&�3>{>�ZE<QϽ(�P?��hF�x"���ȏ��f2?�{G?�ޑ> -�����6�$��A�>7�?��?���>XCJ�[����?���>m����1?ˆ�"���O'���������]*>�d>W>�uJ�0�W�[�s�a�/���?��?�8�=��;�4<�=����I=;Ƅ?g�#?�f*�`	Z��li���W��#J�u'1�+�`�𐜾v/%���m�|���%���O����)�+l�<�-?�ɇ?������鱾7k���9��GQ>P��>��>�z�>O<I>0�Q&3�`_��B#��������>~�z?���>��I? <?DwP?�iL?��>b�>!2���i�>q{�;��>��>��9?0�-?�50?�y?ru+?�.c>z���;����ؾ�
?��?�I?�?;�?y܅�[uý8���Vg�ٱy��|����=�&�<E�׽
<u���T=
T>x�>(K�<��J�F9 ��Z7>��?
�b>H0�>��2����:�5����>���>�0�>��ྮc��{ξ��C?�P�?�#�%�q=l��>�z����R����=���;�=�\u=��:�u�= �	>�WԹ�B��O�ѽ�<�<a�w���`J�>6X'?��>�ܒ>�D�����þȅ�=HV>�J�>��>l�о-#���C��5�d�G�>�S�?l��?[��=��m>g�������Z	߾+�4��F��UPL>��2?�+E?��?�?��B?�C1?2�:��2�]u��
�x��m����?!,?���>n����ʾ��Z�3���?�[?E;a�X���:)��¾��Խ��>>Z/��-~����D��݅�G���v��(��?���?xA�1�6�iy�o���HZ��|�C?n$�>�W�>	�>�)�Z�g�!#��3;>j��>m
R?8��>�?�b|?{�g?�YL>Gu=�����x㧿�����>l�?�fs?��?��}?P��>� �=�������u��V��<�6�\%����\=Ѓ6>�s@>H?P�>�=V=� ֽ#]B=�B���s=��f>p��>ch�>��>�|�>�@>��G?(d�>���0[�l����)v���� w?NL�?�t0?6J�=JG���C�F� ����>P'�?L�?ۼ ?ouy��/�=V)ü�\���Z�Z��>k��>��>v1=� Y=r�6>���>�8�>����>S�!�7�G�
� �?�EI?XϷ=��пT�k��PY�eNS�XjO�w�"����j��dJ�=R�q�!�:�������M�񢏾u��b���I�Ѿ�>��lO?�/>���>��<�5�����vӉ=kҽ)3a>���;:#����=Ÿ��F���`)��I�<M�;�L=��<�־�D�?J!8?Z?�5+?�	w>F�>��>q=I>���4j?h�>� z����V��;�+���4>y7��&$�3�#��{W��)<>��q=���>,��=�CӽWU=�nD>5����Pf=�c����?<�LH>M��<֥2��=~w�==t?Ȕ������X��
��27?y��>��t=�����??K1>�M���繿�|
���~?��?�?��?9Y��/�>`�����ƽ�`@=Ͷt�`�W>��=*���>�?@>!,���߾�����?�@�%??Cy��rο�D8>�T>��>t�O��b,��V���8��;��G'?�4��Q���.�>���=3�ھs�پj:;z�s>&��=3H��<k��U=&Y�Q�4=�t�=���>:�F>ժ�=���M�=%~�=1a>?]R>/e�<�:�KY~���=c >���>-f>�w�>��?��>?^?ݖ�>Ӕp�G�о��ɾ�C>;c=��>a4�<�`�=�w�>��,?H�??�I?���>"»=G��>S��>��!�3�c� ����2��^b>�'�?�_�?�_�>j��=.�<�o:�@�P�Y���*?�`3?�?3��>���S\忔TA��g����=�4�A��j�9�M:R�RLa���潉�6�}�s<35i>�>c��>�rU>�W>`t�=ᆙ>�U>�^=�>w5J=z`��}$��Mߏ<å��=��<���=v��<���N����;<�Г=���<w�<���=���>>>v��>ဖ=���G/>ݵ���L��ǿ=rA���&B�33d��I~�r/��P6�v�B>�2X>�����3��g�?��Y>�q?>K��?�<u?.�>�/�վcQ��[Ee��US�ĸ==�>|�<��y;�X`�Q�M��xҾ��>��>���>n�l>.,��?�T�w=�	�D]5���>K���L�����1q��<��)����	i��˺Z�D?KA���}�=#~?��I?��?���>w#���ؾ�0>�E����=�{q�<J��� ?�'?���>�$���D��[��z��� ?4綾�bf�,���!0��<i��덽��r>���W ��*$E��~�X���<�r����>��3?���?� 0�xQ�vkw�aw ���#>�?a0'?�۴>��?���>�d�����sn���={��?VO�?�z�?�y�>��=������>��?~��?ځ�?mr?(?���>y�h;�#>HV��yP�=,�>�j�=���=��?��?D??F��#	��p���o^�-a�<�1�=译>Aׇ>��t>���=��]=(w�=�X>A1�>G�>;�b>�W�>�D�>����ﾩ�?��/=4m�>M>&?�CM>�QM<�Y���}h=�;���,ٽ-�����|����=��=�g=|�>�5Ŀ��?�Aq>{(�7Y?6N��2��ʩ=g�->�5����>�`�>�E�>e��>�>(,>u�=��=e־��>��
�o!��?C�\U���Ͼ��s>�k���'�ʥ����L�ه�������h�c���b$=�9ȥ<af�?�����h�%M+���G%?�>��3?�����a�>[i�>���>��������컌����A�?[K�?��`>��>��d?�?���N�B��h�,�v��I���c�X_���������c����Z?�cm?�z7?Q5=�M>�n?�{�~�����e>�J�-���d�=\՛>�Ι���z�eʾI.¾3���*�=�7V?�V�?�6'?��,���m�71'>²:?��1?�Nt?��1?7�;?�����$?ml3>�I?�q?FI5?=�.?H�
?W2>�=�s����'=�1����ѽ�xʽκ�t�3='B{=&���f_<�x=[�<h���ټY�;�����<i:=��=��=�>4]?���>�u�>�=6?}Z�g1:��.��-7(?��3=�#��� ���_������j>H<e?�E�?�l]?'Do>2�E�� 1��a&>뇂>�z>��R>���>�L��T=��=}�>L�>�۝=�U��%刾��	�"V����(="�&>�?��t>O��=z�\>�遾�D{�^hJ�6t��H��෎�(�2�>.6�?ݞ�?�>j�\?s:?,�\�T` �ƍ��/^���;?��M?C7?�ol?�vw���`:^�XjO��7��u>,'>�A*��K��A��.:�e6>ƍ>����ꟾ�a>ڄ��3޾in�p�I��\�otG=���P=���վ24}���=��	>���<%!�
�������4J?\8g=����^T�ꉺ�R&>�f�>��>��:�i�w�g@�6g�����=\��>b;>1?����G�� ��>�>�OE?CW_?�j�?2"���s�%�B������d��;ȼi�?�z�>@i?�!B>g��=)�������d�G�I �>X��>��8�G��<���/��J�$���>�8?^�>��?w�R?1�
?��`?*?JD?:%�>w��V���B&?5��?��=��Խ�T�� 9�JF����>{�)?�B�޹�>O�?�?��&?
�Q?�?��>�� ��C@����>�Y�>��W��b��8�_>��J?ך�>r=Y?�ԃ?|�=>\�5��颾�֩��U�=�>��2?6#?P�?���>���>���9�=���>�c?x0�?�o?���= �?;2>���>,��=���>@��>�?PXO?&�s?��J?Z��>���<�6���7��X@s��O��ǂ;�nH<��y=����4t��I�H��<N�;�j��=O�����D�B���5��;}؄>��C>���Lh�������y�$r�>�#��g�`��������&�4t�>:?Ž>���ɨ�<�G�>I��>M�(�y*T?W��>{C!?�X'>��Z��ݸ�0��)�^>a?1�==@A���뎿I�s��Y�<��n?��K?	�k�ֽ��x?��D?� � �H����DW0=Tȟ��LO?��?��!�Ar�>��?�H?��>(�����x�r7��0��k�d��>�J�>K��-��^�>��?׈~>���>r��������B��D��>O�?pr�?T�?�H�=�^��i��hm���A���^?���>�1��
�"?.����Ͼ�N���2���"�X�����M/���j��w$�؃�i׽JA�=��?^s?�Zq?��_?�� ��d�7)^��	��"iV�z����E��'E�7�C���n�c[��������G=��C�'�?�'��?��?�:<�=��>H�侾�-�U��j}$<������=8��>��=�ֳ=u#������"2��xD���:?��=�d�>��2?��V�('�ĭ<�&,�p�޾/l=]0�>��>��?�">�->��:�}!��k�0m_��6v>�xc?W�K?��n?�n�:+1�����s�!�6�/�Qc����B>Qj>e��>�W�����9&��X>���r����w����	�c�~=]�2?<)�>�>�O�?�?r{	��j��}kx�1�1�.��<k/�> i?�@�>��>�нs� �6��>��l?ߧ�>&�>����6Z!�\�{���ʽ�$�>;�>ֶ�>��o>:�,�4#\��j������9�=w�=x�h?����I�`�(�>�R?qW�:|�G<*|�>߲v��!�����'���>7|?���=x�;>�ž�$��{�8��j?)?;E?
��s�*�� ~>�"?���>�-�>�#�?84�>'�þ�{��3�?G�^?�;J?rUA?F@�>E=�w���UȽh�&�_-=���>��Z>�l=.�=���\��w���D=O��=мӓ����<P���tN<o��<�4>mۿ-BK��پ�
����?
�爾⪲�d��x��ib������Wx�{���'�QV��6c�������l����?m=�?f��O0��粚������������>��q������|���(����Ῥ�&d!���O��&i�M�e�S�'?ֺ��ѽǿ߰���:ܾ! ?�A ?�y?��S�"���8��� >�J�<'����뾪����ο(�����^?���>��0��i��>���>ܡX>�Hq>H��螾�/�<u�?�-?.��>o�r��ɿS������<���?'�@t;B?��(�����O_=���>7�?��%>Du9����2����l�>��?	͋?9}=��U���'�iYa?�B�;Y2C�mԹ\f�=�_�=�e/=�]�Y/E>lP�>,�)�;��ݽ�'>`�}>z9�=�
���`��3�<V>����Ǹg�4Մ?+{\�yf���/��T��U>��T?+�>�:�=��,?^7H�[}Ͽ �\��*a?�0�?��?	�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=Q9�(���k���&V����=7��>0�>ق,�ʋ���O��J��T��=���[�ſD�%����"�=B�޻��O�j���ۮ��\H�=ҡ��s����Ǒh=a��=NS>巆>C [>5i_>ݗV?�7k?o!�>�>s��*ሾ�uξ޻Q�}����?��B���Y��/����7�	��+�4����Ⱦ�=���=|6R�Ɩ��	� �F�b��F�W�.?�~$>��ʾ��M�ہ-<Xtʾ�����z祽:7̾"�1�- n�ʟ?i�A?����?�V�7��Ӏ�g�����W?�b����ܬ�cg�=�걼P�=�-�>���=��⾻3�h�S�H9?K?�ϾL�x�fj�=ـ¼� �Pb=?�
�>]��=�l�>c�"?�`����T!>(�;>-I�>�B�>��=>¾`Ci� �"?��V?�8��������>����Q˙= o>�Ai��-`>�GԼbˑ��ȴ<]p�<��>"�l?.g>=��J�6�<���|w>A�>�8h?�]1?�P�>��a?�l?HJ
=ML��r��p//�ۂ^��:?mU?�=r>J���O��=پ��D?O�?���>:.�得/@�h���?�i\?3�>?��;%�|�\k���Q��,?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?r�;<��U��=�;?l\�> �O��>ƾ�z������3�q=�"�>���ev����R,�f�8?ݠ�?���>��������=;ٕ��Z�?��?ڃ���&g<���/l�'n���o�<Fɫ=��wH"����E�7��ƾw�
� ����п����>Z@?Q��*�>cA8�6⿾SϿ+���\о�Pq���?d��>��Ƚ:���t�j�
Pu��G�i�H�m����]�=_��� d=�b�Z��9M%�~��=�¢>�d=2��>_�[��O ��7�O���A��>�G? �>xOn�f�~P�?��+�2\Կ^�����|Ty?R�?N?b?���>n�>}^�:��Ď̽�q<?�ǆ?J^?|/�)笾v��=%�j?�_��wU`��4�uHE��U>�"3?�B�>Q�-�k�|=�>���>g>�#/�x�Ŀ�ٶ�>���W��?��?�o���>p��?ts+?�i�8���[����*�Y�+��<A?�2>���I�!�A0=�PҒ���
?T~0?{�e.��J?6҄���{��AR�oҾ�TO�>8S�݂ܽw�d>�p�� P�GP���ƾ(g�?�@#�?���X0��h?l��>�G��n���#$>o��>� �>�!��h�.=(F�>W��$Z��nY>G��?���?W�	?�ѧ��)��H�,>��^?�)�>�3�?fܶ=aR�>�)�=�a��[�&�&hK>���=�����%?s�G?k�>�q�=\4W��U/���-���I���	��DM��ڙ>�]Y?��A?=K�>	?@���%��
"���	C;��v����Q�x6�'޽%�F>� #>�v�=g�7�վ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Y��D��u�o�y�>���?
�@�ծ?ji�5	?B��L��a~�����7�}��=1�7?�$�y�z>���>��=�ov�����ǿs����>JB�?�y�?���>��l?��o���B�G1=�;�>�k?�u?3q��󾜱B>R�?�������6K��f?��
@�t@G�^?*ꢿun��wԀ�-Gս����1+I=��:��t�==�����{>%��=(�
��t���l�<]O8>�}+>�s�>:�x>��R>J%�=e^z���є��񤿇+w�j�8�js��D���Hj���#�����������ˁ��7�>jd���ǽ�ß<'��=��U?�R?�p?׏ ?4�x�Ԓ>����h'=p~#��΄=�.�>�f2?ߥL?M�*?�֓=ؤ���d�	`��uC��?Ƈ���>�sI>x��>E�>�$�>�0H9�I>�1?> �>� >]'=���]=��N>�N�>���>mx�>��<>�>�ʴ�
*��ډh�wv��̽ �?b��[�J���� /��������=�U.?�Z>����Hп>����&H?�放a(��_+���>ѧ0?�>W?��>�*���MT���> 	���j�XG>����
l�5j)���P>�6?Vm>G
u>̔4�js7��^O�����}�v>u'7?.,����2��r�W�G���ܾ�H>�W�>��������(h��j����=��9?Y!?¿��u9����v��s��.9Q>ށ]>&M=#��=H�N>��h��νE�D��]=��=��^>�?Òs>&8�;���>𧼾}-���F>N)�>���=g�H?��;?� Z=5P���ʔ�s���^:>>�A?�OC>� =�䷾v�e>���>�ل>�`ֻ�(i�x䶽V�����=�D�����/������<���>��=������j���i>��l?����ԙ����(J/���K?���>�$�=���=QS��	��x�����?�n@��?���7�X���?D��?�&��p�>6C�>���>���xV���r'?�0,�]��{��⿾�5�?XЩ?η�<�Ϙ�T�x���->��<?�/ؾv�>�~��R�������u��$=e��>[.H?M=���O��=�d~
??f_򾪪����ȿ�uv�{��>�?r��?�m��C��O@��>��?gY?��i>�_۾1vZ�<��>�@?R?s*�>�:���'���?Ӷ?㰅?HI>���?�s?�k�>,0x��Z/��6�� ����o=:�[;�d�>�W>n���qgF��ד��h��_�j������a>b�$=2�>9E�F4���9�=���H���f�F��>�,q>:�I>W�>i� ?�a�>t��>Ix=[n��,ှ�����L?��?X���!n�F��<�c�=�^�n<?�=4?�W���Ͼ�Ψ>8�\?�?��Z?�e�>���@���꿿鄴��7�<l�K>�A�>J�>��u0K>��Ծ:D��}�>a˗>7����ھX$��� ���8�>gu!?g��>�M�=/!?p#?�tl>�>6F�	��BRE��r�>�'�>+E?~?�t?o����4�8e��Fs����Y��JS>3�w?�@?��>�����1��tA<�ޯ��Ƌ�F��?�_f?,��?�S�?l?@?��A?��]>k��%�۾�������>GTC?$ν��I����u�U�(?��>��?٩��h��c�=��{��Q��>��D?\?���l�����9j�<3{D<�Z� :�=Z��ǀw=�u<��<�!��_�(>(�;>�ל��l�q܂�}I>���>��>���!���$1,?�&?�~����=��r�a>D��?>7�L>�����^?�<��{�����Mj���hU�N�?Ù�?�S�?"t��7�h��8=?E�?V�?=6�>����5T޾g���ow�R�x�l����>{��>��j����u���t��� 0����Ž1GD��!�>5 �>�?A��>Q>h�>����Cn%��}پ=^���_����,/��Y(�R�t��������=ִ��wj����>P��5h�>jf?�I>�Dq>)��>Nr/�o��>�]>�Yo>	��>�6>i>|J�=X�2<eʽٸN?en2�kG�����7���T�>��`?�j�>�?������
�5���>�}�?q%�?�?��a�Bk_���?�A#?�5G�&M?k_���$=��F=fߏ��>�$>n/>�F�>���<� ��eU���=�?5L?�!A����뾽�h����m=�J�?y�(?j�)�g�Q�R�o���W�S��J�Fh�R3��p�$�pp�_叿�^���%��f�(�B�+=S�*?��?���50���k��	?���f>��>n
�>|��>3I>��	�8�1�Q�]�cF'��΃��i�>]X{?���>E�I?^<?�{P?�jL?*��>�S�>�A���c�>���;��>���>)�9?"�-?e30?�|?St+?�-c>�`�����wؾ�	?o�?vK?�?��?yޅ��jý�嗼4(f���y�������=8��<a�׽�t��U=�S>nV?���v�8������ k>�}7?7��>��>����+��}��<	�>��
?AG�>�����|r��a�Z�>
��?���s�=K�)>+��=Ʉ��!qѺ@W�=���1��=�j��li;��<z�=���=)�t�����?�:�F�;�[�<}U�>�h?���>堠>BK��lT�-Y��߯<�x�>���>Ĺ=�����ȉ��
��Ѣb��w>P�?�?�	�����>f8<��Ծ�J6��s0��p*�ד�<�"?E .?p�_?�A�?�PH?�&?	�:=�B��U��Uم�2���1�+?�,?��>���y�ʾD憎ۊ3�x�?�X?�<a����=)�ޖ¾"�Խƶ>�V/��'~�;��~D�ra����(e��R��? ��?�A�1�6�z�켘� P��ÑC?,�>U�>:�>��)���g�V"�`9;>��>�R?硿>�aG?�y?��X?�uG>X�8�0s��ﮛ�lw���#>�:?`�?
j�?�e|?TM�>��>H+9�?�ھ�o꾱���q�k@��6xf=I>
�>1H�>�=�>�W�=��Խ��ս)�T����=/6g>�^�>�ˠ>8\�>G؃>?n	=�]H?ۚ�>�\��u��ݤ��e��BJJ�*&v?q7�?��+?j	!=��AYE������>��?=�?��(?�X��_�=�μh?���Wn��>g�>�>��=�C=��>���>T�>�4����g�8��iN��b?��F?���=������=���ž�Ud��=0=�u߾��/gS��vT��Q>�3Ѿ���>��S>�Vў�ߩ���섾k#�����;7$�>A��=�r>K�>��<�Ѕ<���=�C�=��ӽVi==.J�=(6ڼ�h�:L����,��N�?=��Ӽ)�F�:�?023?U-?ݢ�?�Z��9�;�禽������q>��[?A�>�����
1����6F�=��̾=�4�i�"���`��Ӄ>��6�I�>�Ӝ=~f�<[���V>#j<#�7��<��<���=v�&=��=v�$=j=�=��=��m?˒���!�� \�Y����<?�9�>���=�T��F?w4>][�����
�w��?z�?��?���>��R��'�>�r��b7���=�����	d>~6r=ێ�L1�>��:>����䖿�����}�?5(@&U1?0鍿�ͿΦ >���>�h>��_��r��G�dZc��Е�L�<?�v#��脾��>��Y=psԾ��վ0t�<�AR>�.�=>����q��N<b�ة=3�>��>��>�=��мB�=���=���=�t>�W�=�X��/����Z=�M�>���>�C>l�>	N?h�@?��?��>7��� ��q���X�>���=a?m>�,;<�t=|�_>�f)?�3??�R]?m��>���;��>\��>����-e�\��J�u�v�=Rp�?��?*�>��=�	��*���]���Ѷ�>�U)?��?]n�=YU�*��ZZ&���.�����s���+=]lr�
]U�*���s�׹㽕�=�o�>���>��>MUy>�9>a�N>a�>��>	W�<{�=�͌�Gµ<q��s��=�Z����<(cż�����0'���+������T�;eȆ;.�]<l��;T$�=�N�>��>-��>7%�=-	����%>��|L�_��=�?���l>�:b�b|��O/�D0>���N>"S>M֓��Ӓ�3m?6�Y>�b<>�]�?��j?��>�D�7վ͜�iJs�D\X�$޳=E�>��2�:���^��
K�7Ծ���> �>���>��l>�
,��?�-�w=$��Fb5�N�>�d��v��.�15q��=����ni��5պ�D?hH��D��=r~?
�I?��?�c�>���/�ؾ�(0>%J���7=��&q�n���?�'?��>&�"�D��4Ѿ|�ý�μ>LP�T$Q�猕�Pg0��(��ϯ�.�>З���qվ�m4�"��C܎�H=�Pe��>�5M?���?WQu�;0��W�T���K����?��c?�>�D?�m?����\��M����
�=��q?oK�?�Z�?�P>|��=N��;�>=,	?��?Ƿ�?x�s?#~?�cy�>��;� >]Ƙ��C�=��>f��=/�=&t?��
?9�
?h��9�	������^���<$С=���>fo�>o�r>���=?�g=9s�=B)\>�؞>�>r�d>0�>�M�>�A��pyھ�?c�=�v>�7�>��w>t"���<��$Q�d���a#�毌�,<����Ľ	c̺��2�.�>86>~e
?թ��1��?.2>r��Q?q��8���A�`=9��<J{r=�?�Z�>_X�>w/�>^w�>�$G=̣p=��Y=;�;�>=;
�����B�:5R���ؾ��e>����3��y�?�ڽ�3��������Vj�aA��j?;��A
=�J�?�v�p�l�_�'����v�?�8�>�*8?=z��t搽��>Ch�>�
�>����.y��zӌ�A_㾘%�?F��?p�?>�{�>7�c?��0?�M��]���2[�zB��W2�*Z�{�a�뢄�p�}������ý�D`?�v?Un4?��c=u�?>#z?af��I�M��>��"�|��sF=)R�>Um��fo����Ծ]���B">ʰQ?^��?N~%?�첾n�
,'>��:?q�1?[Ut?l�1?K�;?����$?p3>�H?�q?^K5?B�.?R�
?a2>J�=�����'=�)��t튾M�ѽ=uʽ����3=={=%����<��=��<.��yټ�+;F��9�<K#:=��=r(�=�>N[?��>�>c5?&
8�#H1��R����'?l=�u��q%���o��X8���>��i?��?��[?R�{>,#?��4�j�%>/E�>��!>��W>8g�>��ɽY���n=i�>��>	�~=5���e�����
�H����+=��>]��>ɯ/>�U�=��>w������Kݯ=j���<Z��j��B�Z���D�\���>NQ?B�*?������=�_��WB?06O?tKX?�x?*�ͽQ��%#i�~9Y�K��;NQ�>�a�=��iJ�������� w�>�d>�����(b>����m޾��n�7#J�@�羚oL=
k��+V=�(�վJF��{�=(
>̰���� ����hЪ�S5J?k=�E��|�U�z����>��>��>4�9�jw��y@�&����і=֏�>��:>n ����FdG�'��?�>�OE?�V_?�j�?� ��s�%�B�����wg��+�Ǽ�?�w�>�i?�B>$��=]���H���d�tG���>���>�����G��;���/��h�$�捊>9?^�>��?j�R?��
?��`?0*?�D?$�>
��a���;B&?���?��=��ԽW�T�� 9�,F����>ـ)?ֶB�=��>E�?�?_�&?�Q?\�?F�>\� ��A@�Y��><Y�>��W�eb����_>ݫJ?���>0>Y?�ԃ?��=>��5�'좾�ީ��Y�=�>��2?�4#?��?�>0��>T���s��=R��>�c?�0�?s�o?���=��?�:2> ��>q��=���>u��>�?�WO?�s?7�J?ԑ�>���<?5���8��gEs���O��m�;�vH<H�y=��I+t� K���<�;�t���L��E���D��됼�0�;�m�>��q>��mf >^5����4���'>��<f�w��
������Ї��f�>;?"<�>A��B�=���>6��>)��[�*?۝�>V?JG =d�y6�m� 3�>�xE?��=C�c��`��y�w�={w=��^?(K?��J&ž*+c?s�H? ��H�<����|�ڽ[�U�$v?��>�聾9�>,�~?[dO?��>+���!ҁ�}����o��=���Ħ=��>G�#��]W�G��>��+?�ߢ>w}J>�����|�I�U�+�����>�n�?Ӂ�?O�?l|�=0-���^�(���hD��^^?��>G<����"?=<��ϾVF��x)��?�8���#���?��n��Й$��ꃾ�U׽�ż=��?�s?_q?�_?� �sd��%^�����^V��'��#���E�'E��C�e�n�(^��$������ H=�#�_�&�A.�?�?	ԽK]�>���k2#����5D>^��Bׯ<�P�>-�=��=��M��؋�V<�!�����,?B�=�T?.nh? BK� �<��2�(ZN�!�9���<>���>pL�>�F?R܄=Mm��j�;���i�`�	��8v>$xc?�K?"�n?�l�+1�ㆂ� �!���/��c��G�B>Kh>���>�W�����8&��X>��r����+w����	�d�~=�2?/'�>粜> P�?D?-{	��k��nx���1�^y�<�-�>�i?�>�>��>��Ͻ�� ����>~�l?m��>�ޞ>��0� �g�{�~�̽j�>~�>(��>s�o>�\*�6�Z��	��fÎ�n�7����=��h?����Fb��ڇ>�9Q?3QF;@�:<��>�j���!�ˊ�[)���
>6�?|�=dM=>�4ľ��P|�VQ���)?�N?�A���l*�o5>A�!?���>��>���?7�>�?ľ�����?��^?�J?��@?pb�>d�-=@{��X�ɽ��%��-=fІ>_CY>j�b=���==8�6�\��(�F�G=&u�=BӼ/ ����;<q��ݼ=<��=n�5>�ۿ�J�)Y־;��Eo�[��t���<��5����Z������V�z�ї�
�-��-U�_�h��쏾{�p����?���?�#���ލ��왿����������>�id�5z��Wb��D��Iw��*S��Ʈ������P�q"f�v(c�H�'?�����ǿ鰡��:ܾ5! ?�A ?$�y?��2�"�8��� >�C�<�)��j�뾧�����οߦ����^?w��>��/��e��>ѥ�>��X>�Hq>����螾P4�<��?!�-?	��>�r�&�ɿ^������<���?*�@F�A?O(���x�K=Ұ�>�#?7B>�-��]�hl��]>�>t*�?���?y�S=ȓW�Ľ��c?�1<�%G��o���l�=k��=��=���]K>��>;&��?�Q1޽�f5>��>p�L�n�a�O|�<V^a>�Jٽ����'Մ?�z\��f��/��T���U>��T?�+�>�:�=n�,?7H�c}Ͽ��\��*a?�0�?Ħ�?�(?�ۿ��ٚ>s�ܾ��M?�D6?���>>d&���t��|�=FM�LD����&V�c��=ة�>܀>,�����O�xS��A��=T��ƿ��$�
�H�<�/����X���U���|Q��ߟ�p�>~��sg=��=y�P>3�>S�T>��X>�NW?f�k?/�>�F>��ub���.;r�$��� �G~��*������쾫�߾!3	�-�����ɾ� =���=�4R�ӗ��F� ���b��F���.?�z$>��ʾa�M�Y�-<�nʾ$��������諒�-̾~�1��n��̟?X�A?����+�V�f��ew�����z�W?�O����謾��=���9�=e#�>���=@���3�_}S�n+?��?d�Ͼ).���>x�v���+=��$?l��>;R>8J�>��?
��=(�Zx�=w�f>CN�>n��>�t<�����̽%�?��K?���Î�k�>�澩�e����=�C�=߽���<tSF>�$�����E�	=����ck=7X?�+�>�C�����ľ�CQ����=?w�?p?�^�>��l?oD?+C�<_��f�4A��j�<��K?�hj?|_>�ǽj���W��&k(?0Xk?� h>���9$��7xL�����Q?�h?�+?4�⢃����P!�O>?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?o�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�ٕ��Z�?y�?Y���=@g<{���l��n���}�<FΫ=���G"�����7�@�ƾ��
�����࿼���><Z@�T�h*�>�C8�K6�TϿ-��:\оUSq�U�?a��>I�Ƚ뛣�D�j��Pu�,�G� �H��������>u�=��<����	��c�;�4�>)bS>q��=\g�> C��{�/�׾9����!�>�?B�>~c���~p���?�	��οՑ���׾���?@ �?�t?͔?�����ǾM������>�g?E�?�[d?����t��!�r=۹j?GS���Y`���4�GAE�U>3?/<�>�-���|=��>�|�>�h>Z/�F�Ŀ�׶�Y���x��?r��?7n꾻��>h��?k+?pm��6���X����*�lX)�>A?92>t�����!��2=��ג���
?�w0?�v��'�32Y?q�i�R�h��悿�o�0 �>��e�FF���\�>ZB���k��3���߶�|ߤ?�	@q��?ѓJ����d�A?�	�>9_�ޫ����>+?�P?y��><U>6~7>g�!�(G,�P�=[��?:Y�?e�%?����O����A�=��e?jѵ>r2�?��=ux�>�1�=����%���0�%>��=T0�ʛ?O�N?�3�>ɤ�=Q;��(-�]�B���Q����h�C����>�a?�RL?��_>q���b3������ͽ��8�d���@�D�1�r�۽bC8>:�9>�>��D���о��?�o��ؿ�i���o'�~54?ָ�>��?�����t�����;_?wz�>�6��+���%���A�a��?�G�?M�?ͻ׾F̼�>r�>}I�>O�Խ4���Ԃ��<�7>ҞB?@�cD���o���>���?��@uծ?si�	?<�I��e~����'7�� �=��7?e�7�z>r��>��=�qv������s�¶>@�?�x�?B��>��l?�|o���B�1=�@�>��k?�u?�tr�K��6�B>"�?�������C��$f?��
@�u@�^?{梿S˿������Ӿ�bU�j�P>쐻�1�>��伆��;Jξ=���� p��b�r�H>C�~>6v�>i�E>nB>#��=��w�i�"�����N��ɺ(��!���[�Lh1�! ��]e�pӾ����*o3�%:g�
  �H�C��;����1�0��=�U?�R?�p?č ?F�x�[�>P���#�=(�#�%�=T2�>�]2?��L?�*?��=����.�d�~^���C��J���w��>KuI>�z�>GC�>�"�>ʼ|9��I>�?>Hv�>�� >�A'=���7=��N>�O�>���>�x�>�s<>�>@ȴ�"-���h�v�v�ei˽��?����|�J����8��)���4ɞ=RM.?�i>�� Cп�����#H?ݔ�!%�ӡ+�Q>�0?FW?q^>�	��N-S�Ҟ>����j��)>�����k��m)��Q>??A'g>�&u>��3��[8�q�P��6��ƽ|>Q6?�ᶾ�"9�^tu�y�H��cݾ��L>���>�Y;��p�����rti��|=�b:?��?����˰�<'v�[}��eR>�]>��=�9�=�M>�e�L�ƽx�F�!�1=���=Z�]>���>DV�><X����>�����>��>)�>���=Տ^?y�C?��\>�S��r!ݾ&�����>���>�H�= �T���g�P>2�>	��>�2ѽ�Q��A_����f�+>�E���Ⱦ
=�Cb<��9�˹E>S�~�w��8"�)-T>7~?�~��f^��d���]ޒ>�v?]� >C[>�@>S�'��읿_˾��?��@��?�jD��At�"89?��?�ؼk�>��>@��>"�Ǿ\X½TX%?�'%�~����׾��8x�?Ȯ?���x:��X(u���V>��?�x��h�>�v�Z��m���u�v�#=#��>69H?(U��4�O��>�w
?�?_�������ȿ�{v����>�?e��?;�m�eA���@���>��?EgY?Jpi>�h۾�eZ�ˊ�>޻@?�R?��>9��'�A�?�ݶ?���?YI>u��?s?^h�>�4x�QY/�=6��]���#u=�b\;w`�>�U>����deF�3ד��h��@�j����B�a>O�$=��>�5�u5���9�=�싽,F����f�Ȥ�>&+q>��I>�X�>h� ?�`�>\��>�n=�c��䀾�����K?���?���An�*ؾ<f �=�|]��?
�3?��E�GYξtݨ>4\?#Z�?�Z?�
�>����U�����fh��p��<�`K>Z�>���>�ሽ}�I>"xվ`�C����>�Ș>�k��$�پ�2��ާ��d�>��!?W��><Q�=��#?p� ?�>�B�>��S�<��\m+��T�>��>��7?�f�?�?_���q@�bp��dܚ�=N���d>R*y?w?Q�c>���8 ��OꂽI�<�5���ن?��X?iJ)�/�?�B�?)�D?��H?܋)>Y/x������8��Vo>�M+?ւǽ�4�ї��A�U�?E?E[?q���!�_�=JX���㾬��>�D?�:?�f�b�u��ܾ�l�:!K�=V<�<�=���=��.>�4J<L���n�.>^�>ƕ�>�|���n�'�۽�Y�=`�?B�>��8��K~�=,?v�G�{ۃ�O�=u�r�xD���>�IL>�����^?{k=���{�����x���	U�� �?��?5k�?���5�h��$=?�?Q	?"�>1K���}޾�ྍPw��~x��w�u�>���>�l�U�;�������|F���Ž�N����>���>h�?n ?�=N>��>N���^M'����r�N^^���� 8��).�=�Yq��1F ���������$�y�{��>܈���>Xj
?Ѵk>�]|>���>
��l��>]�Q>��~>h��>R
U>&�3>{>�ZE<QϽ(�P?��hF�x"���ȏ��f2?�{G?�ޑ> -�����6�$��A�>7�?��?���>XCJ�[����?���>m����1?ˆ�"���O'���������]*>�d>W>�uJ�0�W�[�s�a�/���?��?�8�=��;�4<�=����I=;Ƅ?g�#?�f*�`	Z��li���W��#J�u'1�+�`�𐜾v/%���m�|���%���O����)�+l�<�-?�ɇ?������鱾7k���9��GQ>P��>��>�z�>O<I>0�Q&3�`_��B#��������>~�z?���>��I? <?DwP?�iL?��>b�>!2���i�>q{�;��>��>��9?0�-?�50?�y?ru+?�.c>z���;����ؾ�
?��?�I?�?;�?y܅�[uý8���Vg�ٱy��|����=�&�<E�׽
<u���T=
T>x�>(K�<��J�F9 ��Z7>��?
�b>H0�>��2����:�5����>���>�0�>��ྮc��{ξ��C?�P�?�#�%�q=l��>�z����R����=���;�=�\u=��:�u�= �	>�WԹ�B��O�ѽ�<�<a�w���`J�>6X'?��>�ܒ>�D�����þȅ�=HV>�J�>��>l�о-#���C��5�d�G�>�S�?l��?[��=��m>g�������Z	߾+�4��F��UPL>��2?�+E?��?�?��B?�C1?2�:��2�]u��
�x��m����?!,?���>n����ʾ��Z�3���?�[?E;a�X���:)��¾��Խ��>>Z/��-~����D��݅�G���v��(��?���?xA�1�6�iy�o���HZ��|�C?n$�>�W�>	�>�)�Z�g�!#��3;>j��>m
R?8��>�?�b|?{�g?�YL>Gu=�����x㧿�����>l�?�fs?��?��}?P��>� �=�������u��V��<�6�\%����\=Ѓ6>�s@>H?P�>�=V=� ֽ#]B=�B���s=��f>p��>ch�>��>�|�>�@>��G?(d�>���0[�l����)v���� w?NL�?�t0?6J�=JG���C�F� ����>P'�?L�?ۼ ?ouy��/�=V)ü�\���Z�Z��>k��>��>v1=� Y=r�6>���>�8�>����>S�!�7�G�
� �?�EI?XϷ=��пT�k��PY�eNS�XjO�w�"����j��dJ�=R�q�!�:�������M�񢏾u��b���I�Ѿ�>��lO?�/>���>��<�5�����vӉ=kҽ)3a>���;:#����=Ÿ��F���`)��I�<M�;�L=��<�־�D�?J!8?Z?�5+?�	w>F�>��>q=I>���4j?h�>� z����V��;�+���4>y7��&$�3�#��{W��)<>��q=���>,��=�CӽWU=�nD>5����Pf=�c����?<�LH>M��<֥2��=~w�==t?Ȕ������X��
��27?y��>��t=�����??K1>�M���繿�|
���~?��?�?��?9Y��/�>`�����ƽ�`@=Ͷt�`�W>��=*���>�?@>!,���߾�����?�@�%??Cy��rο�D8>�T>��>t�O��b,��V���8��;��G'?�4��Q���.�>���=3�ھs�پj:;z�s>&��=3H��<k��U=&Y�Q�4=�t�=���>:�F>ժ�=���M�=%~�=1a>?]R>/e�<�:�KY~���=c >���>-f>�w�>��?��>?^?ݖ�>Ӕp�G�о��ɾ�C>;c=��>a4�<�`�=�w�>��,?H�??�I?���>"»=G��>S��>��!�3�c� ����2��^b>�'�?�_�?�_�>j��=.�<�o:�@�P�Y���*?�`3?�?3��>���S\忔TA��g����=�4�A��j�9�M:R�RLa���潉�6�}�s<35i>�>c��>�rU>�W>`t�=ᆙ>�U>�^=�>w5J=z`��}$��Mߏ<å��=��<���=v��<���N����;<�Г=���<w�<���=���>>>v��>ဖ=���G/>ݵ���L��ǿ=rA���&B�33d��I~�r/��P6�v�B>�2X>�����3��g�?��Y>�q?>K��?�<u?.�>�/�վcQ��[Ee��US�ĸ==�>|�<��y;�X`�Q�M��xҾ��>��>���>n�l>.,��?�T�w=�	�D]5���>K���L�����1q��<��)����	i��˺Z�D?KA���}�=#~?��I?��?���>w#���ؾ�0>�E����=�{q�<J��� ?�'?���>�$���D��[��z��� ?4綾�bf�,���!0��<i��덽��r>���W ��*$E��~�X���<�r����>��3?���?� 0�xQ�vkw�aw ���#>�?a0'?�۴>��?���>�d�����sn���={��?VO�?�z�?�y�>��=������>��?~��?ځ�?mr?(?���>y�h;�#>HV��yP�=,�>�j�=���=��?��?D??F��#	��p���o^�-a�<�1�=译>Aׇ>��t>���=��]=(w�=�X>A1�>G�>;�b>�W�>�D�>����ﾩ�?��/=4m�>M>&?�CM>�QM<�Y���}h=�;���,ٽ-�����|����=��=�g=|�>�5Ŀ��?�Aq>{(�7Y?6N��2��ʩ=g�->�5����>�`�>�E�>e��>�>(,>u�=��=e־��>��
�o!��?C�\U���Ͼ��s>�k���'�ʥ����L�ه�������h�c���b$=�9ȥ<af�?�����h�%M+���G%?�>��3?�����a�>[i�>���>��������컌����A�?[K�?��`>��>��d?�?���N�B��h�,�v��I���c�X_���������c����Z?�cm?�z7?Q5=�M>�n?�{�~�����e>�J�-���d�=\՛>�Ι���z�eʾI.¾3���*�=�7V?�V�?�6'?��,���m�71'>²:?��1?�Nt?��1?7�;?�����$?ml3>�I?�q?FI5?=�.?H�
?W2>�=�s����'=�1����ѽ�xʽκ�t�3='B{=&���f_<�x=[�<h���ټY�;�����<i:=��=��=�>4]?���>�u�>�=6?}Z�g1:��.��-7(?��3=�#��� ���_������j>H<e?�E�?�l]?'Do>2�E�� 1��a&>뇂>�z>��R>���>�L��T=��=}�>L�>�۝=�U��%刾��	�"V����(="�&>�?��t>O��=z�\>�遾�D{�^hJ�6t��H��෎�(�2�>.6�?ݞ�?�>j�\?s:?,�\�T` �ƍ��/^���;?��M?C7?�ol?�vw���`:^�XjO��7��u>,'>�A*��K��A��.:�e6>ƍ>����ꟾ�a>ڄ��3޾in�p�I��\�otG=���P=���վ24}���=��	>���<%!�
�������4J?\8g=����^T�ꉺ�R&>�f�>��>��:�i�w�g@�6g�����=\��>b;>1?����G�� ��>�>�OE?CW_?�j�?2"���s�%�B������d��;ȼi�?�z�>@i?�!B>g��=)�������d�G�I �>X��>��8�G��<���/��J�$���>�8?^�>��?w�R?1�
?��`?*?JD?:%�>w��V���B&?5��?��=��Խ�T�� 9�JF����>{�)?�B�޹�>O�?�?��&?
�Q?�?��>�� ��C@����>�Y�>��W��b��8�_>��J?ך�>r=Y?�ԃ?|�=>\�5��颾�֩��U�=�>��2?6#?P�?���>���>���9�=���>�c?x0�?�o?���= �?;2>���>,��=���>@��>�?PXO?&�s?��J?Z��>���<�6���7��X@s��O��ǂ;�nH<��y=����4t��I�H��<N�;�j��=O�����D�B���5��;}؄>��C>���Lh�������y�$r�>�#��g�`��������&�4t�>:?Ž>���ɨ�<�G�>I��>M�(�y*T?W��>{C!?�X'>��Z��ݸ�0��)�^>a?1�==@A���뎿I�s��Y�<��n?��K?	�k�ֽ��x?��D?� � �H����DW0=Tȟ��LO?��?��!�Ar�>��?�H?��>(�����x�r7��0��k�d��>�J�>K��-��^�>��?׈~>���>r��������B��D��>O�?pr�?T�?�H�=�^��i��hm���A���^?���>�1��
�"?.����Ͼ�N���2���"�X�����M/���j��w$�؃�i׽JA�=��?^s?�Zq?��_?�� ��d�7)^��	��"iV�z����E��'E�7�C���n�c[��������G=��C�'�?�'��?��?�:<�=��>H�侾�-�U��j}$<������=8��>��=�ֳ=u#������"2��xD���:?��=�d�>��2?��V�('�ĭ<�&,�p�޾/l=]0�>��>��?�">�->��:�}!��k�0m_��6v>�xc?W�K?��n?�n�:+1�����s�!�6�/�Qc����B>Qj>e��>�W�����9&��X>���r����w����	�c�~=]�2?<)�>�>�O�?�?r{	��j��}kx�1�1�.��<k/�> i?�@�>��>�нs� �6��>��l?ߧ�>&�>����6Z!�\�{���ʽ�$�>;�>ֶ�>��o>:�,�4#\��j������9�=w�=x�h?����I�`�(�>�R?qW�:|�G<*|�>߲v��!�����'���>7|?���=x�;>�ž�$��{�8��j?)?;E?
��s�*�� ~>�"?���>�-�>�#�?84�>'�þ�{��3�?G�^?�;J?rUA?F@�>E=�w���UȽh�&�_-=���>��Z>�l=.�=���\��w���D=O��=мӓ����<P���tN<o��<�4>mۿ-BK��پ�
����?
�爾⪲�d��x��ib������Wx�{���'�QV��6c�������l����?m=�?f��O0��粚������������>��q������|���(����Ῥ�&d!���O��&i�M�e�S�'?ֺ��ѽǿ߰���:ܾ! ?�A ?�y?��S�"���8��� >�J�<'����뾪����ο(�����^?���>��0��i��>���>ܡX>�Hq>H��螾�/�<u�?�-?.��>o�r��ɿS������<���?'�@t;B?��(�����O_=���>7�?��%>Du9����2����l�>��?	͋?9}=��U���'�iYa?�B�;Y2C�mԹ\f�=�_�=�e/=�]�Y/E>lP�>,�)�;��ݽ�'>`�}>z9�=�
���`��3�<V>����Ǹg�4Մ?+{\�yf���/��T��U>��T?+�>�:�=��,?^7H�[}Ͽ �\��*a?�0�?��?	�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=Q9�(���k���&V����=7��>0�>ق,�ʋ���O��J��T��=���[�ſD�%����"�=B�޻��O�j���ۮ��\H�=ҡ��s����Ǒh=a��=NS>巆>C [>5i_>ݗV?�7k?o!�>�>s��*ሾ�uξ޻Q�}����?��B���Y��/����7�	��+�4����Ⱦ�=���=|6R�Ɩ��	� �F�b��F�W�.?�~$>��ʾ��M�ہ-<Xtʾ�����z祽:7̾"�1�- n�ʟ?i�A?����?�V�7��Ӏ�g�����W?�b����ܬ�cg�=�걼P�=�-�>���=��⾻3�h�S�H9?K?�ϾL�x�fj�=ـ¼� �Pb=?�
�>]��=�l�>c�"?�`����T!>(�;>-I�>�B�>��=>¾`Ci� �"?��V?�8��������>����Q˙= o>�Ai��-`>�GԼbˑ��ȴ<]p�<��>"�l?.g>=��J�6�<���|w>A�>�8h?�]1?�P�>��a?�l?HJ
=ML��r��p//�ۂ^��:?mU?�=r>J���O��=پ��D?O�?���>:.�得/@�h���?�i\?3�>?��;%�|�\k���Q��,?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?r�;<��U��=�;?l\�> �O��>ƾ�z������3�q=�"�>���ev����R,�f�8?ݠ�?���>��������=;ٕ��Z�?��?ڃ���&g<���/l�'n���o�<Fɫ=��wH"����E�7��ƾw�
� ����п����>Z@?Q��*�>cA8�6⿾SϿ+���\о�Pq���?d��>��Ƚ:���t�j�
Pu��G�i�H�m����]�=_��� d=�b�Z��9M%�~��=�¢>�d=2��>_�[��O ��7�O���A��>�G? �>xOn�f�~P�?��+�2\Կ^�����|Ty?R�?N?b?���>n�>}^�:��Ď̽�q<?�ǆ?J^?|/�)笾v��=%�j?�_��wU`��4�uHE��U>�"3?�B�>Q�-�k�|=�>���>g>�#/�x�Ŀ�ٶ�>���W��?��?�o���>p��?ts+?�i�8���[����*�Y�+��<A?�2>���I�!�A0=�PҒ���
?T~0?{�e.��J?6҄���{��AR�oҾ�TO�>8S�݂ܽw�d>�p�� P�GP���ƾ(g�?�@#�?���X0��h?l��>�G��n���#$>o��>� �>�!��h�.=(F�>W��$Z��nY>G��?���?W�	?�ѧ��)��H�,>��^?�)�>�3�?fܶ=aR�>�)�=�a��[�&�&hK>���=�����%?s�G?k�>�q�=\4W��U/���-���I���	��DM��ڙ>�]Y?��A?=K�>	?@���%��
"���	C;��v����Q�x6�'޽%�F>� #>�v�=g�7�վ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Y��D��u�o�y�>���?
�@�ծ?ji�5	?B��L��a~�����7�}��=1�7?�$�y�z>���>��=�ov�����ǿs����>JB�?�y�?���>��l?��o���B�G1=�;�>�k?�u?3q��󾜱B>R�?�������6K��f?��
@�t@G�^?*ꢿun��wԀ�-Gս����1+I=��:��t�==�����{>%��=(�
��t���l�<]O8>�}+>�s�>:�x>��R>J%�=e^z���є��񤿇+w�j�8�js��D���Hj���#�����������ˁ��7�>jd���ǽ�ß<'��=��U?�R?�p?׏ ?4�x�Ԓ>����h'=p~#��΄=�.�>�f2?ߥL?M�*?�֓=ؤ���d�	`��uC��?Ƈ���>�sI>x��>E�>�$�>�0H9�I>�1?> �>� >]'=���]=��N>�N�>���>mx�>��<>�>�ʴ�
*��ډh�wv��̽ �?b��[�J���� /��������=�U.?�Z>����Hп>����&H?�放a(��_+���>ѧ0?�>W?��>�*���MT���> 	���j�XG>����
l�5j)���P>�6?Vm>G
u>̔4�js7��^O�����}�v>u'7?.,����2��r�W�G���ܾ�H>�W�>��������(h��j����=��9?Y!?¿��u9����v��s��.9Q>ށ]>&M=#��=H�N>��h��νE�D��]=��=��^>�?Òs>&8�;���>𧼾}-���F>N)�>���=g�H?��;?� Z=5P���ʔ�s���^:>>�A?�OC>� =�䷾v�e>���>�ل>�`ֻ�(i�x䶽V�����=�D�����/������<���>��=������j���i>��l?����ԙ����(J/���K?���>�$�=���=QS��	��x�����?�n@��?���7�X���?D��?�&��p�>6C�>���>���xV���r'?�0,�]��{��⿾�5�?XЩ?η�<�Ϙ�T�x���->��<?�/ؾv�>�~��R�������u��$=e��>[.H?M=���O��=�d~
??f_򾪪����ȿ�uv�{��>�?r��?�m��C��O@��>��?gY?��i>�_۾1vZ�<��>�@?R?s*�>�:���'���?Ӷ?㰅?HI>���?�s?�k�>,0x��Z/��6�� ����o=:�[;�d�>�W>n���qgF��ד��h��_�j������a>b�$=2�>9E�F4���9�=���H���f�F��>�,q>:�I>W�>i� ?�a�>t��>Ix=[n��,ှ�����L?��?X���!n�F��<�c�=�^�n<?�=4?�W���Ͼ�Ψ>8�\?�?��Z?�e�>���@���꿿鄴��7�<l�K>�A�>J�>��u0K>��Ծ:D��}�>a˗>7����ھX$��� ���8�>gu!?g��>�M�=/!?p#?�tl>�>6F�	��BRE��r�>�'�>+E?~?�t?o����4�8e��Fs����Y��JS>3�w?�@?��>�����1��tA<�ޯ��Ƌ�F��?�_f?,��?�S�?l?@?��A?��]>k��%�۾�������>GTC?$ν��I����u�U�(?��>��?٩��h��c�=��{��Q��>��D?\?���l�����9j�<3{D<�Z� :�=Z��ǀw=�u<��<�!��_�(>(�;>�ל��l�q܂�}I>���>��>���!���$1,?�&?�~����=��r�a>D��?>7�L>�����^?�<��{�����Mj���hU�N�?Ù�?�S�?"t��7�h��8=?E�?V�?=6�>����5T޾g���ow�R�x�l����>{��>��j����u���t��� 0����Ž1GD��!�>5 �>�?A��>Q>h�>����Cn%��}پ=^���_����,/��Y(�R�t��������=ִ��wj����>P��5h�>jf?�I>�Dq>)��>Nr/�o��>�]>�Yo>	��>�6>i>|J�=X�2<eʽٸN?en2�kG�����7���T�>��`?�j�>�?������
�5���>�}�?q%�?�?��a�Bk_���?�A#?�5G�&M?k_���$=��F=fߏ��>�$>n/>�F�>���<� ��eU���=�?5L?�!A����뾽�h����m=�J�?y�(?j�)�g�Q�R�o���W�S��J�Fh�R3��p�$�pp�_叿�^���%��f�(�B�+=S�*?��?���50���k��	?���f>��>n
�>|��>3I>��	�8�1�Q�]�cF'��΃��i�>]X{?���>E�I?^<?�{P?�jL?*��>�S�>�A���c�>���;��>���>)�9?"�-?e30?�|?St+?�-c>�`�����wؾ�	?o�?vK?�?��?yޅ��jý�嗼4(f���y�������=8��<a�׽�t��U=�S>nV?���v�8������ k>�}7?7��>��>����+��}��<	�>��
?AG�>�����|r��a�Z�>
��?���s�=K�)>+��=Ʉ��!qѺ@W�=���1��=�j��li;��<z�=���=)�t�����?�:�F�;�[�<}U�>�h?���>堠>BK��lT�-Y��߯<�x�>���>Ĺ=�����ȉ��
��Ѣb��w>P�?�?�	�����>f8<��Ծ�J6��s0��p*�ד�<�"?E .?p�_?�A�?�PH?�&?	�:=�B��U��Uم�2���1�+?�,?��>���y�ʾD憎ۊ3�x�?�X?�<a����=)�ޖ¾"�Խƶ>�V/��'~�;��~D�ra����(e��R��? ��?�A�1�6�z�켘� P��ÑC?,�>U�>:�>��)���g�V"�`9;>��>�R?硿>�aG?�y?��X?�uG>X�8�0s��ﮛ�lw���#>�:?`�?
j�?�e|?TM�>��>H+9�?�ھ�o꾱���q�k@��6xf=I>
�>1H�>�=�>�W�=��Խ��ս)�T����=/6g>�^�>�ˠ>8\�>G؃>?n	=�]H?ۚ�>�\��u��ݤ��e��BJJ�*&v?q7�?��+?j	!=��AYE������>��?=�?��(?�X��_�=�μh?���Wn��>g�>�>��=�C=��>���>T�>�4����g�8��iN��b?��F?���=������=���ž�Ud��=0=�u߾��/gS��vT��Q>�3Ѿ���>��S>�Vў�ߩ���섾k#�����;7$�>A��=�r>K�>��<�Ѕ<���=�C�=��ӽVi==.J�=(6ڼ�h�:L����,��N�?=��Ӽ)�F�:�?023?U-?ݢ�?�Z��9�;�禽������q>��[?A�>�����
1����6F�=��̾=�4�i�"���`��Ӄ>��6�I�>�Ӝ=~f�<[���V>#j<#�7��<��<���=v�&=��=v�$=j=�=��=��m?˒���!�� \�Y����<?�9�>���=�T��F?w4>][�����
�w��?z�?��?���>��R��'�>�r��b7���=�����	d>~6r=ێ�L1�>��:>����䖿�����}�?5(@&U1?0鍿�ͿΦ >���>�h>��_��r��G�dZc��Е�L�<?�v#��脾��>��Y=psԾ��վ0t�<�AR>�.�=>����q��N<b�ة=3�>��>��>�=��мB�=���=���=�t>�W�=�X��/����Z=�M�>���>�C>l�>	N?h�@?��?��>7��� ��q���X�>���=a?m>�,;<�t=|�_>�f)?�3??�R]?m��>���;��>\��>����-e�\��J�u�v�=Rp�?��?*�>��=�	��*���]���Ѷ�>�U)?��?]n�=YU�*��ZZ&���.�����s���+=]lr�
]U�*���s�׹㽕�=�o�>���>��>MUy>�9>a�N>a�>��>	W�<{�=�͌�Gµ<q��s��=�Z����<(cż�����0'���+������T�;eȆ;.�]<l��;T$�=�N�>��>-��>7%�=-	����%>��|L�_��=�?���l>�:b�b|��O/�D0>���N>"S>M֓��Ӓ�3m?6�Y>�b<>�]�?��j?��>�D�7վ͜�iJs�D\X�$޳=E�>��2�:���^��
K�7Ծ���> �>���>��l>�
,��?�-�w=$��Fb5�N�>�d��v��.�15q��=����ni��5պ�D?hH��D��=r~?
�I?��?�c�>���/�ؾ�(0>%J���7=��&q�n���?�'?��>&�"�D��4Ѿ|�ý�μ>LP�T$Q�猕�Pg0��(��ϯ�.�>З���qվ�m4�"��C܎�H=�Pe��>�5M?���?WQu�;0��W�T���K����?��c?�>�D?�m?����\��M����
�=��q?oK�?�Z�?�P>|��=N��;�>=,	?��?Ƿ�?x�s?#~?�cy�>��;� >]Ƙ��C�=��>f��=/�=&t?��
?9�
?h��9�	������^���<$С=���>fo�>o�r>���=?�g=9s�=B)\>�؞>�>r�d>0�>�M�>�A��pyھ�?c�=�v>�7�>��w>t"���<��$Q�d���a#�毌�,<����Ľ	c̺��2�.�>86>~e
?թ��1��?.2>r��Q?q��8���A�`=9��<J{r=�?�Z�>_X�>w/�>^w�>�$G=̣p=��Y=;�;�>=;
�����B�:5R���ؾ��e>����3��y�?�ڽ�3��������Vj�aA��j?;��A
=�J�?�v�p�l�_�'����v�?�8�>�*8?=z��t搽��>Ch�>�
�>����.y��zӌ�A_㾘%�?F��?p�?>�{�>7�c?��0?�M��]���2[�zB��W2�*Z�{�a�뢄�p�}������ý�D`?�v?Un4?��c=u�?>#z?af��I�M��>��"�|��sF=)R�>Um��fo����Ծ]���B">ʰQ?^��?N~%?�첾n�
,'>��:?q�1?[Ut?l�1?K�;?����$?p3>�H?�q?^K5?B�.?R�
?a2>J�=�����'=�)��t튾M�ѽ=uʽ����3=={=%����<��=��<.��yټ�+;F��9�<K#:=��=r(�=�>N[?��>�>c5?&
8�#H1��R����'?l=�u��q%���o��X8���>��i?��?��[?R�{>,#?��4�j�%>/E�>��!>��W>8g�>��ɽY���n=i�>��>	�~=5���e�����
�H����+=��>]��>ɯ/>�U�=��>w������Kݯ=j���<Z��j��B�Z���D�\���>NQ?B�*?������=�_��WB?06O?tKX?�x?*�ͽQ��%#i�~9Y�K��;NQ�>�a�=��iJ�������� w�>�d>�������2b>���v޾P�n�J�{���L=Jq�/&V=��־9:�~M�=v 
>ϯ���� ����rΪ��9J?}j=�b��\uU�p���>���>�֮>.:�/�v��@������)�=���>�!;>����Z��nG�}4�:=�>�PE?mW_?vj�?� ���s���B�����Ig��GGȼW�?�w�>�f?�B>:��=𘱾M��d��G��>��>�����G��<��`0����$����>f7?�>�?`�R?�
?Ǚ`?�*?�D?�%�>�������A&?2��?��=<�Խ�T�� 9�ZF�7��>S�)?,�B����>D�?ν?��&?�Q? �?��>� ��C@�ה�>dY�>��W��b����_>��J?��>�=Y?�ԃ?�=>J�5��颾�֩�mU�=�>��2?6#?N�?ů�>`��> ���Yπ=���>uc?�.�?��o?Un�=��?�I2>���>(�=)��>��>�?�PO?�s?�J?%��>�{�<'M�� ���as���N���;�9H< �y=(n�%It��
�ݙ�<$�;-~���~�������D�HN�����;��>�G?>��˾�u�>�a�,�u��=Kľ�jK���Ҿ6(����8��>�s*?a}�>z'���<s(�>�W ?�	H�m�F?�?�C�>D��<�<�V�B��d��ͺ�>
L3?�5=1.?�;ͩ��\��NN�=�<;?3�|?�����,�b?��]?��=���þ�~b�U{�=�O?��
?گG�F�>��~?m�q?��>ڽf�4Pn����N>b��[j��׵=-��>�>�q�d�ם>q�7?�?�>=�b>��=�۾��w�����M?E�?���?���?�*>r�n�I.��s���<���]?9$�>�����"?<����о�!:���⾷/���ޫ�H�� �����$��ă�}�սV�=�?S�r?�q?��_?�� �md���]�b�� vV�1��e�S�E�bE�:HC��In�u�s(��_���F=O���9�x��?��?j�K�>�|���R�=���)�e����)*ܼY�g>@�->D&%>��Z=8���'%���s��}?TKt>���>B�P?�(��`6I���'���,���5�$�I�A*Z>>�?dd�>��'���;���Q.Z�}:�=I/v>3{c?�K?��n?Ue��*1�ц���!���/�y[���B>�j>���>v�W�9���6&�2S>���r����#y��M�	���~=�2?�)�>}��>�N�?�?�z	��g���fx���1�я�<**�>�i?TE�>���>9�Ͻ�� ���>�k?���>G��>�����B�s:z������*�>��>�c ?�t>:0��Z�S���i��k:�h��=Ti?SI��
�W���>i�P?��*�3<��>ݜ�����<��8D*�h >f�?��=�>>�ȾEk��~��`��o(?��?^>��	*���~>�"?���>�]�>4��?��>|^ľ]m����?�w^?�kH?�u??%V�>��.=q�����ʽ,*�b�8=��>�_>�d=6
�=����,Y��R ���X=/�=O<ü���%��;�d���I0<ԑ�<]�0>����U�_���3%6�.��h��,��;���J�
��,����JV���i�,0$�j�(<$_�?Yw�����gU�Y^�?�0�?��7�=@ƾ#4���݄�yaҾX��>����mP��?����½�n�����4�Ҿ�M �y�Y�6�G��B=�O�'?ɺ��ƽǿİ��);ܾ�  ?�A ?��y?��t�"���8�?� >�M�<�"��k�뾌����οƦ����^?���>��
1�����>���>١X>�Hq>����螾�8�<��?��-?^��>l�r�'�ɿA���c��<���?0�@N5G?�9E�c���=��>>G ?щ>(@�B~��LȾ�>9A�?Bϔ?^?�=�ES���ս.[?�Gy=�L;�ےмc>@��=ۭ�<�k�Ջ�>���>�n1�M�(���*��+@>&=�>[ܔ���B�t��zvR=Z,�>�����0�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��=p���iƿ~�!�-e!��g�<3Q � g��;��ܨ��!V��f��=Zu�Y,�Y�[=�x�=�K>`�>~lP>�V>�Z?sm?@��>���=LX��J��,̾K���gn�֜�����&I�eB�����޾i	���������žL'=���=�*R�7����� ��b�t�F�t�.?Ñ$>��ʾ��M��+<�oʾIĪ����ӥ�.̾��1�Dn�{ϟ?{�A?�􅿨�V�������b��Q�W?�F����מּ��=߲���=b+�>w��=��{3��xS��,?�?Ͼ�o�>����9�K=E�%?��>7׳<j��>:� ?&!���Ƚ�nM>=�>��>N�>g�>b��Lڽ�Q?d�Q?��-#��Uy>-���!DR�\�=�>��)������PI>�T+�5���.W�(?����<.dw?o5M>w�U�nx���=�6_>�>6�?���>c�>��?ٖa?n3E�+$��~����Ҿڌ2>��j?N�J?E�<�D�<i� ��喾"|0?�c?���,�羂R)��r �J[?�X?m;C?6�6�������a�?���`?p�v?�q^�/s��`����V��?�>�]�>���>\�9�1m�>��>?i#��G��3���aZ4�TÞ?��@���?�;<y�	��=`9?b[�>.�O�c;ƾ������niq=��>-���8av�����N,���8?���?���>B���y�����=�ٕ��Z�?z�?�����>g<R���l��n���z�<CΫ=#��D"�����7���ƾ��
�誜��߿�Υ�>9Z@�U轆*�>=D8�T6�TϿ"��.\о�Sq�y�?J��>��Ƚj���/�j�}Pu�d�G�#�H������Y>>���<ڨ4>�����]��>�<���_���>�\$>��x>Q��L���dӾY����?=j>?��>b�f�yȾUO�?M�
�+:οD��[㦾o`?0��?~��?�W?��->S."���оD傽�D?���?�D]?9c�=�	���Ҿm?�?��k��Q3��P+��X>��%?��>�[!���=m7J>EK�>a}�=u<(��9ȿ���d���x�?P�?�S���?�a�?d�)?r%�e���2���'��}6;�G.?��>�Kɾ����O0�|�n���>��!?p�����#���S?�Xo�$Z�n�g�?0��?��>H����80�t`G>��m��LX�2��DBf�P�?"@N"�?�M������?G�?&	�F���ÿ=�"?~�?z��=�m�=��=��꾟�)�;�=1�?�	�?���>�"��瞛�$�J>s?�1�>݄�?sC����>N�A>g�����%��ɑ>��<�<uS#?�v?��#>�k��:�Ѿ�sh�=�N��5����
�c��H?��n?�T?� >��S���¼���=�B�S��;��x��2���bٽ���_�>��{>���>lx���:�2�?�o���ؿ�i���l'�c54?=��>��?�����t�����:_?{�>6��+���%��A�0��?G�?��?��׾�(̼�>o�>!G�>��ԽN��S���c�7>T�B?!�)D����o�]�>c��?r�@ծ?4i��	?���P��Ua~����7�a��=��7?�0��z>���>��=�nv�޻��W�s����>�B�?�{�?��>#�l?��o�O�B�o�1=7M�>̜k?�s?Qo���g�B>��?"������L��f?�
@u@a�^?*xhֿ����|N��M���I��=��=��2>I�ٽ`�=D�7=��8��=��5��=x�>��d>�q>G(O>�a;>�)>���J�!��q��[���5�C������Z�7��OXv�>z��3�������?���3ý�x���Q�$2&��?`�e��=iV?D�Q?��o? � ?Xz���>1����<ף!�a �=d�>��1?9)L?>D*? �=+���+e��u��8�����-M�>�H>�L�>pe�>�ԭ>]O9��I>R�>>d�>�#>�S'=5��=A�O>)��>96�>�F�>�C<>��>Fϴ��1��k�h��
w�p̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�6`>�+ �~l���)��%Q>wl? �f>�u>b�3�Se8���P��{��Ni|>�36?v鶾�B9��u�L�H�cݾ�FM>ľ>�$D��k�X������ui��{=xx:?A�?�6���ⰾ�u��C���PR>`;\>LW=Vf�=YXM>"bc���ƽ�H��d.=z��=�^>��>7�>R`	� l�>9Ԋ����g�>��=���>�A?\��>z	�Z�K�[:'�o�_��~�=Yw�>,�>�~h>�`���-ջ���>�!>J�=��ٶe�?t����>�/%<4T����~�]��=�ĺ�e��;^��<{�������;]ـ?}м��
����徍G�=�<c?��
?N�=�!m=t{ ����O]׾���?+k@�;�?��XL�M�.?�-�?<x�P��Z>��?�����8�3|?sq-�s�̾�W�SY��0Q�?Q�?��G��{��"^��:]�>7$+?/�վQh�>�x�~Z�������u�T�#=:��>�8H?�V��$�O��>��v
?�?�^�ة����ȿ4|v����>V�?���?Z�m��A���@����>/��?�gY?�oi>�g۾�_Z����>��@?�R?��>�9�o�'�p�?�޶?ӯ�?�I>���?�s?|j�>v$x�5Z/�_6�������e=��[;�e�>fW>���lgF��ד�[h���j����~�a>&�$=��>Y?��4��+7�=b����H���f����>�.q>��I>�U�>� ?pa�>���>�s=�o��=���񸖾��K?���?,���2n�O�<T��='�^��&?�I4?�j[�y�Ͼ�ը>�\?j?�[?d�><��Q>��G迿8~��?��<��K>)4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,���R��HB�>�e!?���>�Ү=� ?S�#?4�j>t(�>�`E��9���E�p��>��>�H?��~?��?�ӹ��Y3�����桿�[�<N>��x?�U?�ʕ>6���v���gE��BI�����F��?tg?]Q彼?�1�?��??;�A?�(f>���ؾs����>G�!?,� �A��I&�		�
}?Q?��>�?����ս/oּ���9x��C?�&\?�?&?��)a� �¾��<��"���U�ɑ�;FD���>��>����Ӓ�=>�ڰ=Qm�wF6�"�f<Lm�=��>8 �=�37��|���<,?��G��샾��=	�r��kD�S�>HL>"���ѩ^?�b=���{�R���u��&U����?���?�n�?x����h�-=?/�?(?2�>4��~�޾R���?w��ux�;e��>���>w�l��}�������}C�� �Žg3���>^y�>��	?�:�>��T>-��>����@�vؾL5��V����W/�2�-������������`�ƾ����N�>�ԫ��¿> �?�
G>�7b>�7�>�|�<��>r�C>��>���>�6>w{&>O��=�⸼�n�.W?
��6��=�=�8�&�?��?>k>��о͉�eS(�ƒ(?�m�?��?_�>6f���K���?J�2?�-��ƀG? �
��{c=�|;��@������JMV>	q��Ҡ>b�Ž=�<�iON��a	�i��>@ ?�<��aT=ђ���n=VM�?L�(?Y�)���Q��o�w�W�aS�z��3:h��i���$�=�p�B쏿k^��:%����(��y*=|�*?��?��#�����%k��?�y[f>
 �>0#�>�ݾ>RvI>�	���1�w^��L'�����*Q�>�Z{?h|�>�I?�;?UrP?dL?S>�T�>j0��*t�>?*�;G�>���>b�9?��-?x*0?�k?�v+?�Tc>�F��6��ÌؾE?4�?�M?G?��?O߅�Eýo[����d�x�y��Y���=N��<y�׽mwu��T=��S>�??�Y�r(;�����1m>�N5?�R�>Ұ�>�Ã�
j���<���>2Q?�)�>7&�6�q���
����>�u�?�J ��֧<�/>x�=%���q뻫��=�����ߜ=�¼r���B˂��9�=���=��ƻ|׃�VͻK�y���<���>a�?�"�>��>����f �Pq���=�5Y>�S>m�>��ؾC{��R(��H�g���y>���?醴?~!e=���=�l�=۬��l/���������7��<�?��"?�T?Ѧ�?��=?Ol#?�>gJ�*\��tc����*�?!,?�>���u�ʾ>�c�3��?�U?�=a����<)�ߌ¾��Խ'�>JY/��+~����D�;������w����?+��?bA���6�Ws�.���T]����C?��>oT�>�>d�)���g��#�$&;>���>R?F_�>Ik:?:�q?xy[?Ѧ�=�J� '���`��wį�0��<1�*?�z?_��?�i�?/A�>+�'>urg�ϐ���9ž2M����9ۚ��>k*>t'�>79�>X��>�Z�<ӌ���d����V�KF>�rh>�]�>9ѡ>$�>��>��	>_�V?�ϰ>V������ ž���d�>�o�?�F�?��]?��
>}-%��`�W�*���>䧷?�'�?P�6?wľ^�k>*����O���!?u�>�P�>܃I=�ď�	o�<��g?�|�>�����c���b�l}���
?D�w?)��=~�ҿ�]���_��׾Y/��b������F����w��Y��<�]��\�#�� ��繾U�Ǿyn;j[�]慾]r ��F?�Q=6`v>���>6�=��>g�=�f����4;^����#����}}��Eu���&����='a�=<�>C��;��ؾH�u?��E?��>�V?��U>�۽�}�>�����>.�P?�n�>6X������<���R�=��?��*,�	V����Ǿyp->t���F= ��=2�� �<��=�+Y;���Tq<{��=�fz=�ӣ=��>^p4=�7O>��[>�6w?W�������4Q��Z罢�:?�8�>?{�=\�ƾ]@?Q�>>�2������ib�.?���?�T�?6�?7ti��d�>e��b䎽Uq�=����{>2>k��=H�2�K��>��J>���K�������4�?��@��??�ዿɢϿJa/>Nx7>�X>�S��1��\���b��@X��3!?��:���˾�>�9�=�v޾)�žJ-=��4>�{g=�c���[�`�=w*z�<6>=�%q=0��>aD>4�=*U���{�=CNP=���=�P>I+��&=���1�(�-=��=�a>Fx&>�8�>�?�!;?�Ic?ߣ>쑉�
A��h�>>���=遄> Sa=��>x��>��5?��W?��O?��>s�=Ԛ�>�ɉ>r0�wwj�W��x��9f>�t�?˪�?�k�>�s*=+�O���_A��Խ�?9�5? �	?Hh>�V���vV&��.�.���S8��R�*=�jr��PU�
���*k�\���==m�>u��>t�><Ry>��9>��N>&�>��>Z�<�H�=���<���m��=q%��g�<��żS����%���+�����3�;��;ǜ]<K��;)��=k��>h�>ޥ�>���=����z/>�Ɩ�5QL�$�=p§�X�A���c�7�}���.�%�6��;C>�Y>R��t'����?��Y>�?>�p�?�.u?Qi>�y���Ծ����	d��S��V�=Fc>f�=��o;��*`�jN�JXҾ���>��>�ў>�j>�*�� >�e�t=� ߾[4���>i���Q��*���p��_��,=���gi��R���C?�h���x�=d~?�I?~��?��> ����ؾ��,>M���ł
=}%���p��?���W?3'&?O��>(���)F�j ���@����>&�4��g^��񐿐S*��=��~"��S��>ޭ�u��B�0�t������2��9o�q>�>�)A?/��?�gh�MIc�p�Q����S�?��^?���>�:�>���>"(��*�K!;�&^>J�?U�?�ʼ?ÿ�=�<�=Ԩ��Q�>��?�9�?,��?׮m?!XE����>TO�<��>�����t�=��>@4v=���=��?T?�8?-���1��S�澣i��3�E�G�<��=!��>C�>�g>Z�=�e>=���=�@Y>���>,�>�Z>*��>`ˁ>�_���S	�)u?��-=��>�R?#2|>�1���9�='��<ѷԽ�Mj�3���M%��5��84�R��<��">�S<$��>����fͣ?E61>B �yr�>nƺ�+�_��n=�!��y��8%�>Ē4>ݔ�>=i�>_�>�Ǐ=^�^>�k�=T�Ծ��>�$�;�!�D�G�S��(Ҿ�/w>I���3'����Wg���uG�5﴾�/�i�i��B��7�<�l��<L�?	���k�2�(������?y,�>N/5?����s�����>��>��>����󖕿�������鳋?��?=8>���>�g?4s!?l�\���e�{J��W�����[�Z�f��d�h���z���@�6=�e?�~r?��?/ˋ<�UD>\�[?\�ߣ�`��>�,������6�.>}Dk��t�����cܾ����0��=d\m?��x?'��>yL��Fq�*�'>%�:?�1?$&t?o�1?�:?lh���$?W�4>jW?m?��4?%?.?B�
?�(2>��=��λ�'=k�������Y�н�dʽ�X�bm3=�"z=�>��<4=)��<	�R�Լ0GB;3Ѣ��p�< K7=h�=���=iӤ>9\?.�>L}�>^�5?�I�|�9�����V!.?�#C=�(��H���ͤ���>�ii?TB�?~�Y?�/f>�jC�D�F�v�>�T�>.>�]Y>�x�>|���?�!�=��>�0>c��=��Z����9�`5���<��>R�>-�>�D$�FiP>�7��~�s�(�>q�}��l���Hk��EI�C�,��A{�u�>8�N?�N$? ��=�Y޾|4���f��r'?�rE?��9?���?;�G=5_�qC�zM����J��>C �<Q3��a�����=�$��$=�yM><ɼ�Z
��_C>I=m��mR��J�� 6j��0���*]�����/�>����s�F���I(�=<q�>����u ��ț�J���*�M?�2�ϭ;�t���(��g=�31>o�>ؑQ�(�F��9�v�I>��>��#>.Z�Z5�z�?��Ѿt�|>-�C?��f?_Ĉ?��U�Z?_��\J�:xܾ�c�����'!?E^�>�q	?�O>b= u¾��	�z�Z���8�A|�>U�>:2���@� ���Ɂ�A&�n�>^F?p�>�a?�W?N?�k?��,?H�>�1s>UGw��n��*B&?��?��=�Խ��T�- 9��F� �>ۃ)?��B�̸�>~�?=�?*�&?�Q?۵?N�>� ��C@����>QY�>��W�zb���_>��J?V��>�<Y?�ԃ?m�=>c�5�ꢾ�ة��T�=�>��2?"6#?ï?`��>g��>G���u�=���>�c?�0�?�o?���=&�?�:2>R��>���=���>S��>�?OXO?(�s?��J?Ǒ�>���<�7���8���Cs���O��ɂ;�pH<Y�y=����3t�.K�,��<d �;�g���H�����l�D��������;g��>�cy>z���K�.>��������dF>�4����M~��U�5��=��>�?�ђ>��)����=��>=��>Y* ��B*?s�?�?���;��`��j׾�=W���>��A?���=;6j�V��R�u���a=y`m?�~\?Mjb�����,6k?z�B?IT����$���־|+M��)��߭}??t�/��>���?6�?[� ?)�
�,(p��謹��@�Y�����5>�A0>xNP�<�q�JuU>�=?�U?���=V�>J 辰����L���?2�?��?��?�{�=��~��׿�]��4��MU?fH�>[>��Z�/?�'�9u־�r��3@�Ǿ<ޱ������l�������w�����9������<�?*9n?Դm?�]?���]�%ae��r�VN��M�K�$4F���D��1?��b����ei۾ �q��[�=����&�4�?�U2?㹾��m>�������Ꮌ��d�>��s�Hf���O�=״;�&�>LU<O�<� �o������x6?b�>fg�>� -?��f��]=��0���;�%� �G��>"]�>���>L;�>�=��㒅<��'_־G8���q�N�k>(c?��N?@q?Y���S(�ń������t����dL>5z>��>�sh��e0��^&�)�:��-n�����<��c��Ϧ=��5?w��>ݚ�>"��?"u
?>�&r����b���0�b׶<���>�Cg?�|�>F҉>�ڽ+S!�c��>�ol?��?.�#>>�߽b������#	���>�"3= �?7',>�	L�n�r�nў� ����$��c�>q�g?t$���^���U�>"�y?|��|>ft5>�;> 6��{�x� �҉�>F��>ς|=�ō>$���tVƾ��q�QӴ��O)?�K?J꒾�*��6~>$"?R��>�.�>I1�?�(�>qþ{�@�ұ?0�^?.AJ?�SA?H�>3�=���aAȽ�&�Ф,=���>��Z>7m=�}�=����t\��v���D=�p�=�μ�M����<�����K<���<��3>���QI?�����s�Ӿ^����
��Yn��Q�3q\�b�������Qv�OD\�=w���g�0�h��o*��w�����B�?i��?>�Ƚ���+\��W~������u>])o�}��='Ɛ�jȽ�����q"\�M/���2��`�&�m�U�'?�����ǿ𰡿�:ܾ*! ?�A ?<�y?��4�"���8�Z� >D�<0+����뾠�����ο(�����^?m��>��Q/��f��>ѥ�>ǡX>�Hq>����螾m/�<��?,�-?��>��r�*�ɿc���9Ĥ<���?,�@�A?��(�y����T=���>2�	?`�?>@�0��4����<O�>�:�?M��?*ON=�W���	�xpe?l�<� G����#,�=:i�=<a=H���SJ>Z�>r����A���ܽ�4>�҅>�#�d��(�^�@E�<P�]>�sԽ������?�u����q�K�o~n��Ӑ>Ի_?���>��>��?PH:�����B���I?��@ǁ�?Z�?�
&���>1�Y�<??��3>n�@�H;v��CK><����=\��3y�f{�>���>St�>�ɽ�x�\^���Ľ���>Z��3Ŀ��.����D=�8����?3��u���]�󢏾�nR���ͽ��=�g�=��'>��>�QZ>�~E>�"[?��}?��>4J>�*�WH��:`ξr����|�#潞so�F�Ľ�&������cھ� �B��mm���!=���=7R�f���C� �c�b�J�F���.?�v$>U�ʾ��M���-<pʾS���rۄ��ॽ�-̾�1�*"n�k͟?��A?������V�]���W�����K�W?P�ͻ��ꬾ��=x���V�=%�>ኢ=���� 3��~S�N�1?`5?F
��ƹ���>�A.�i�n=��C?g��>l*���>Ȍ8?�d=B�0>���=��<�A�>L?Ls�=�(�0���&?[K?/;�)�;���>����ܿ��?C=���=��V�dU">{z�>�]$=G8ھ`v�<�*<T�j>�!W?���>@�)��
��P�����V�<=��x?r�?��>�yk?��B?��<>k����S���Pw=��W?�!i?��>p�����Ͼ.���q�5?u�e?��N>]hh�u�龡�.�EM��-?o�n?�X?x��� y}�!������n6?�K�?��w�"㞿T�������>�Y�>\�?c!=�{��>��i?�M>������~���P'���?�x@��?��=�N���|O=��>���>��_q��`e��G����=9]�>�KL�Z|`�Z�(�Q|��jH?��?�~�>�Ȏ�yE-����=�ٕ��Z�?|�?v���wHg<M���l��n���~�<�Ϋ=+��F"������7���ƾ��
����9⿼ͥ�>BZ@�U�w*�>�C8�Y6�TϿ'���[о�Sq�u�?,��>t�Ƚ����7�j��Pu�L�G��H������k�>��>�X��؛��	w���9�_j��tC ?����_>,2%�^✾#&���G=^3�>-s�>�R>c���*q��� �?.g ��*ҿϤ�������Q?���?댄?a�'?����ݑ��r�a�}4=�<P?hs?�\?ܞ��I@d��$���j?W_��xU`��4�FHE�<U>�"3?%C�>D�-�°|=�>���>�g>^#/�_�Ŀ�ٶ����R��?͉�?�o���>m��?~s+?�i�8��B[����*��+��<A?�2>����!�0=�+Ғ���
?>~0?�{�O.���_?<�a�d�p�R�-��ǽ '�>��/��[��H���-��e��	���ly�ԭ?>d�?�?d��&#��$?Ւ�>C���=Ǿ���<X��>��>��N>÷`�U-v>1�M;�ڟ	>J��?�a�?�g?D���� =>�~?氒>!h�?��<��?��>vپ:[>�e>��=A���*��>��U?�?�ܤ>TGW��b$���!��{(��׻�0�f����>��T?�|r?�i�>�!n��M5;��Q�f�G=�@˽�*�Jی�� ��找��>�I�>p�=숾�ͤ���?Pp�8�ؿ j�� p'��54?2��>�?��z�t�����;_?Jz�>�6��+���%���B�`��?�G�?>�?��׾�R̼�>D�>�I�>Y�Խ����Z�����7>3�B?V��D��r�o�|�>���?	�@�ծ?li���?y�5��p��]���Z��@�'��>�9?R�
�p��>���>�C�y�u��	��Ad�v��>�s�?���?̞?p��?B��-i���c�����>�:�?/	?�)>���N�=T#8?�&��F������k�N?u�@@�MN?ű���hֿ����_N��P�����=���=Ն2>�ٽ,_�=��7=��8�B=�����=t�>��d>"q><(O>a;>��)>���Q�!�r��\���S�C�������Z�C��Xv�Xz��3�������?���3ýy���Q�2&�)?`�z��=b�U?t�Q?i6p?� ?}�y�o$ >s���e?=%�#����=>�k2?��L?y*?+��=䱝�L�d��=���o��xӇ�gm�>p�I>�t�>1E�>�	�>�<9��!J>a�>>�.�>>Z�$=1���e�=5O>�>&��>�m�>�Y<>�>[ϴ�1/��>�h���v� �˽��?>i��k�J�K3��*��׏��
��=�c.?��>���n=п����.H?����-���+�">��0?\W?�>����O T��'>���j�8U>�# �TKl���)�fQ>�e?��c>m"t>�q3���7���N�_���A�>#_4?i���?6��t��LH���YLI>yý>_�	�L[�Eܖ���~��&i��Lk=�:?��?����Cn����y��V����T>0�]>α"=tq�=LrO>?:Y�W�����F�ˎ.=u��=��W>&&?/c+>��=���>���_N�{��>��A>RK*>H�??*"%?fU��Й�B����-�O)w>��>P��>%�>KJ�x��=��>�kb>I0�����^��\�@��W>Qp����_�I<x�A�v=���c�=�D�=����*<�<'=�~?���(䈿��e���lD?S+?a �=!�F<��"�E ���H��G�?r�@m�?��	�ߢV�?�?�@�?!��P��=}�>	׫>�ξ�L��?��Ž7Ǣ�Ȕ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ\h�>ux�{Z�������u���#=J��>�8H?�V��q�O�'>��v
?�?�^�ة����ȿ9|v����>P�?���?i�m��A���@�n��>2��?�gY?�oi>�g۾�`Z���>λ@?�R?2�>�9�7�'�p�?�޶?ȯ�?�G>m��?Zs?��>�cl��..��Z���"�����=�����>���=�p����F��4��{��+�i����I"b>E�#=��>�t὞i��㰴=׫��N5��Ǆc���>n�m>�DJ>Ӥ�>?� ?yH�>.\�>�q=�:��EI��i���;[?��x?�LA�Oi�3-�=��>�cJ��Z.?ݔm?d���4F뾢��>'f?)��?KJ>?
�>�:��⓿!���־s�#>�l >�֏>
�?�7�Q����j�e�þ���>��>���� � �`H���o�
�;>��M?�+?�Ȑ=�?�J?�m�>��>k8"��|��|K���	?�~�>�\�>�X�?a�?�KL�7��A"��]ҧ���U���k>��k?xvB?Ѹ�=%ݝ�с���u'�ѣn�"�A>i	�?��w?�]��Z��>,Ԍ?1FT?|F~?���>-]W����3���8">� ?el�T-A�9�%��&�@�	?�W?P��>��y-ӽ�Lü�����<?7p[?�/&?2��a�k�ľ���<�q.�BB�{�<1q��>$C>���mF�=L>��=H�n�6&6�W�h<�Z�='>�F�=�83�Yb��=,?�G�_ۃ���=^�r�(xD��>�IL>���y�^?m=�0�{�����x��(	U� �? ��?^k�?k��.�h��$=?�?9	?p"�>K��~޾��+Pw�g}x�qw�!�>��>�l���G���ə��~F��*�Ž2�6��>ȥU>C��>C?��>�i�>���0�Z��aϾ�˾W�G���?�N3��9%���ʾz񭾹��%uO�R۾��t��G�>[Gw��<>��?�9>�&�>���>�>���>��R>39X>��e>��p>���=t�{=�#:;&u�MX?������2�z�p����W>?��d?*?Vj=�J����i(?��?�&�?Q�>ٜV�L[<���>im�>�U{�B�?�H˼X$2���=�F��;j0�^��T=>��>����`6�qP���o��w?�o)?i�0=11쾨��O�׾<��<`�?��A?EB]����2Ae��*j�״'���>ٵ��
+�>�־J�d�p�i�\������.?��C=�?$A?�׾��˾��W�6C@�*����>�D�>?e>��>��=N� ��Z��m{�C|����?�?*�>,K?�):?��Q?FwM? -�>�a�>�=���?�>g��;ޟ>���>� :?�[.?�i.?�?Y�)?{Ga>��s ��b׾&T?��?�8?]�?�?�Ċ��ٶ�)���W`���u�b��Tv=��<(н�S��e�V=h�T>�X?���8�m���Gk>�7?��>���>'���.�����<��>D�
?�I�>2 ��}r�qb��X�>0��?��|=�)>R��=H����kԺ�c�=����L�=�"���y;�><捿=� �=��s�Y������:�d�;R��<]��>h.?z%�>�J!>���r�ݾKs6�^��<��>��=%V�=v�&���t��R��o�w����>���?� �?�A�<5��=���=O������������l���>��?xJ;?Lך?�
I?LA0?/=
�2�c��Hi���ck��
?m!,?��>�����ʾ��щ3�۝?�[?g<a�����;)�5�¾��Խ��>�[/�b/~�����D� 䅻���'~����?߿�?�A�M�6�@x�Ŀ���[����C? "�>�X�>��>�)�0�g�P%��1;>��>5R?y�>9�O?�A{?��[?�vT>�8��2��w̙��5�p�!>�@?m��?���?	y?�^�>q�>��)��ྜྷB�����4�ׂ�LgW=�Z>~��>M0�>��>���=��ǽ�����>�:m�=d�b>s��>͏�>���>ހw>ҷ�<I�G?���>�Z��<��&夾)Ã��C=��u?��?�+?�=��+�E��F��E�>�n�?���?6*?}�S�L��=m�ּݶ�"�q��%�>|Թ>*�>Bϓ=�F=0m>2�>M��>���`��s8�O�M���?F?t��=.ſ�>p��l��"����B<�썾N�a�E��;�a�z��=W����#������Z�b蝾w퐾�I��/6������0 �>�X�=�*>wW�=��<�7ȼ��J<:2=Q�t<��<�y�r~F<+�<����"�}�p�J��ti<�EW=���
Wʾ~?-OH?I�>?U�H?�Ƃ>���=rsԼ��{>T	��~?v>O�9ݗ���N]�h%���G��/�˾K����`�^0���'>������>��3>�r>�{=n=�=bK=gj�=E!<���<�>��=po=J��=�J>{��=���?tȑ��ϗ�ud�9@=k?2/�>�\>'�Ͼ@�_?��>�	���<�������?7S�?K��?���>�վ��p>�H��������&>���br=�K�=�q�‾>�>Z)/��^����=&g�?�@@��0?J���Eտ�p�<#�3>{�>�R���0�FDR���T���P�Me?�=��hʾ'�>�ή=例Gƾv�#=j
;>��K=v>�t�[��3�=�z��M=��r=k{�>�E>�
�=rl��ڸ=�W?=�=W_M>�#�}�H�̽+��2=\i�=��d>�">-��>~�?�b0?sYd?E8�>�n��!Ͼ�:���B�>��=�G�>^؅=�pB>Ŋ�>D�7?z�D?s�K?H��>t=S�>��>��,�ֲm�k��ѧ�G��<$��?+Ά? Ѹ>�R<s�A�G���b>��%Ž�r?�P1?ll?��>{���߿�!�l>)�}x�'�/� �H=%J���,���������ٽ|$�=Q�>�-�>�җ>Gw>�=>o�P> �>`{2>n�K=�ڮ=��q<��Ѽ6GR=`i��_�=�
z�Z��<R�;�������2�������;F7߼X��=���>�>"�>ն=���*9>l����Q���='����A�Hf�L|�?�.���*���<>ұI>�� c����?^U>� =>���?�s?��">h��e�Ӿ\ɛ�ll]���G����=+��=�I�];:��_�+L��xѾ���>S�>F�>F�l>�	,�� ?���w=�a5�g�>�x�������:7q�o?��9���i��CѺS�D?SF�����=�"~?n�I?f�?���>�����ؾM/0>PD����=��#q�ah����?�'?�>u�n�D�d�׾�+y�x?�e���Rg�ʠ�[]�w+��~��E�?I̾�몾R�%�鉚��悿ɴ`���ǽ忪>Q~?�5�?݁���у�������̾6Α=O&+?E��?�=�@?k��>޷��l�$�z��a$=d��?��?t��?��>�j�=�����+�>�*	?��?#��?ys?cw?��P�>���;�� >����Q��=��>U�=l'�=a?�~
?��
?V\��E�	�S�����e1^��I�<̾�=�>w�>��r>�;�=0�g=���=8W\>H�>ӏ>g�d>��>I0�>�ʦ��~��5?�y=+�>]3I?���>�o	��G�=]�=��;=Nhf��쎾��߽�;��H~�=�M��-m�FJ:�l��>�{��}?�?Sl>�%��?xW�uX�A->�
>-�d�(Ũ>��>>�>/��>�W�>Q�>9?�>�ϩ=ޯپ��>J ��P���I�i�X��־�8X>c|����	�n�
��FսQ40� ��������n�������@��<<�ۍ?��#f���%�ei��?R�>S�6?x��'1��
=�=��>�>2�^E��w�����ܾ~�?7*�?`!*>��> p5?�: ?������<�^M�?|p���:�hy��`�����	���f�]�̼�*t?�Dg?{�;?\�ýBw8>%��?�.�ssy�!G�>�S�̑X�aDs=;��>�Qھ[�Ծ��3��:���2�+r=��S?S��?�0=?�{5��+4���>���>\[?h<?��>�M?l�U���F?%E�"��>��6?�'4?`�I?Y��>ײ>�ӹ����:��p>����Ő��<��~ac�Oɽek->%2�=��ߞ�=��<!.=�k���κ���=!��<q%~=Q]���=�#>dO�>��`?��>��=>U
7?�@�xyM�N��Z5?���ä�m���8���ۧ ��:�Yb?9�?�Bq?B�;>��;��+�C�,>�j#>o>,>ޮ!>��b>� ���ݽ�>�7Z>a9> B>�ս-������V��)`n=��'>l��>���=��K��S�;ͯ��J���>�sp��]�pBg���V���/�,�����>�;[?�,?���=<)
���J=����\�U?ȯ?��H?�?���=(Ѿ�.B��+���o]����>#����.�YF��^ܶ��������St>�ϾZ
��_C>I=m��mR��J�� 6j��0���*]�����/�>����s�F���I(�=<q�>����u ��ț�J���*�M?�2�ϭ;�t���(��g=�31>o�>ؑQ�(�F��9�v�I>��>��#>.Z�Z5�z�?��Ѿt�|>-�C?��f?_Ĉ?��U�Z?_��\J�:xܾ�c�����'!?E^�>�q	?�O>b= u¾��	�z�Z���8�A|�>U�>:2���@� ���Ɂ�A&�n�>^F?p�>�a?�W?N?�k?��,?H�>�1s>UGw��n��*B&?��?��=�Խ��T�- 9��F� �>ۃ)?��B�̸�>~�?=�?*�&?�Q?۵?N�>� ��C@����>QY�>��W�zb���_>��J?V��>�<Y?�ԃ?m�=>c�5�ꢾ�ة��T�=�>��2?"6#?ï?`��>g��>G���u�=���>�c?�0�?�o?���=&�?�:2>R��>���=���>S��>�?OXO?(�s?��J?Ǒ�>���<�7���8���Cs���O��ɂ;�pH<Y�y=����3t�.K�,��<d �;�g���H�����l�D��������;g��>�cy>z���K�.>��������dF>�4����M~��U�5��=��>�?�ђ>��)����=��>=��>Y* ��B*?s�?�?���;��`��j׾�=W���>��A?���=;6j�V��R�u���a=y`m?�~\?Mjb�����,6k?z�B?IT����$���־|+M��)��߭}??t�/��>���?6�?[� ?)�
�,(p��謹��@�Y�����5>�A0>xNP�<�q�JuU>�=?�U?���=V�>J 辰����L���?2�?��?��?�{�=��~��׿�]��4��MU?fH�>[>��Z�/?�'�9u־�r��3@�Ǿ<ޱ������l�������w�����9������<�?*9n?Դm?�]?���]�%ae��r�VN��M�K�$4F���D��1?��b����ei۾ �q��[�=����&�4�?�U2?㹾��m>�������Ꮌ��d�>��s�Hf���O�=״;�&�>LU<O�<� �o������x6?b�>fg�>� -?��f��]=��0���;�%� �G��>"]�>���>L;�>�=��㒅<��'_־G8���q�N�k>(c?��N?@q?Y���S(�ń������t����dL>5z>��>�sh��e0��^&�)�:��-n�����<��c��Ϧ=��5?w��>ݚ�>"��?"u
?>�&r����b���0�b׶<���>�Cg?�|�>F҉>�ڽ+S!�c��>�ol?��?.�#>>�߽b������#	���>�"3= �?7',>�	L�n�r�nў� ����$��c�>q�g?t$���^���U�>"�y?|��|>ft5>�;> 6��{�x� �҉�>F��>ς|=�ō>$���tVƾ��q�QӴ��O)?�K?J꒾�*��6~>$"?R��>�.�>I1�?�(�>qþ{�@�ұ?0�^?.AJ?�SA?H�>3�=���aAȽ�&�Ф,=���>��Z>7m=�}�=����t\��v���D=�p�=�μ�M����<�����K<���<��3>���QI?�����s�Ӿ^����
��Yn��Q�3q\�b�������Qv�OD\�=w���g�0�h��o*��w�����B�?i��?>�Ƚ���+\��W~������u>])o�}��='Ɛ�jȽ�����q"\�M/���2��`�&�m�U�'?�����ǿ𰡿�:ܾ*! ?�A ?<�y?��4�"���8�Z� >D�<0+����뾠�����ο(�����^?m��>��Q/��f��>ѥ�>ǡX>�Hq>����螾m/�<��?,�-?��>��r�*�ɿc���9Ĥ<���?,�@�A?��(�y����T=���>2�	?`�?>@�0��4����<O�>�:�?M��?*ON=�W���	�xpe?l�<� G����#,�=:i�=<a=H���SJ>Z�>r����A���ܽ�4>�҅>�#�d��(�^�@E�<P�]>�sԽ������?�u����q�K�o~n��Ӑ>Ի_?���>��>��?PH:�����B���I?��@ǁ�?Z�?�
&���>1�Y�<??��3>n�@�H;v��CK><����=\��3y�f{�>���>St�>�ɽ�x�\^���Ľ���>Z��3Ŀ��.����D=�8����?3��u���]�󢏾�nR���ͽ��=�g�=��'>��>�QZ>�~E>�"[?��}?��>4J>�*�WH��:`ξr����|�#潞so�F�Ľ�&������cھ� �B��mm���!=���=7R�f���C� �c�b�J�F���.?�v$>U�ʾ��M���-<pʾS���rۄ��ॽ�-̾�1�*"n�k͟?��A?������V�]���W�����K�W?P�ͻ��ꬾ��=x���V�=%�>ኢ=���� 3��~S�N�1?`5?F
��ƹ���>�A.�i�n=��C?g��>l*���>Ȍ8?�d=B�0>���=��<�A�>L?Ls�=�(�0���&?[K?/;�)�;���>����ܿ��?C=���=��V�dU">{z�>�]$=G8ھ`v�<�*<T�j>�!W?���>@�)��
��P�����V�<=��x?r�?��>�yk?��B?��<>k����S���Pw=��W?�!i?��>p�����Ͼ.���q�5?u�e?��N>]hh�u�龡�.�EM��-?o�n?�X?x��� y}�!������n6?�K�?��w�"㞿T�������>�Y�>\�?c!=�{��>��i?�M>������~���P'���?�x@��?��=�N���|O=��>���>��_q��`e��G����=9]�>�KL�Z|`�Z�(�Q|��jH?��?�~�>�Ȏ�yE-����=�ٕ��Z�?|�?v���wHg<M���l��n���~�<�Ϋ=+��F"������7���ƾ��
����9⿼ͥ�>BZ@�U�w*�>�C8�Y6�TϿ'���[о�Sq�u�?,��>t�Ƚ����7�j��Pu�L�G��H������k�>��>�X��؛��	w���9�_j��tC ?����_>,2%�^✾#&���G=^3�>-s�>�R>c���*q��� �?.g ��*ҿϤ�������Q?���?댄?a�'?����ݑ��r�a�}4=�<P?hs?�\?ܞ��I@d��$���j?W_��xU`��4�FHE�<U>�"3?%C�>D�-�°|=�>���>�g>^#/�_�Ŀ�ٶ����R��?͉�?�o���>m��?~s+?�i�8��B[����*��+��<A?�2>����!�0=�+Ғ���
?>~0?�{�O.���_?<�a�d�p�R�-��ǽ '�>��/��[��H���-��e��	���ly�ԭ?>d�?�?d��&#��$?Ւ�>C���=Ǿ���<X��>��>��N>÷`�U-v>1�M;�ڟ	>J��?�a�?�g?D���� =>�~?氒>!h�?��<��?��>vپ:[>�e>��=A���*��>��U?�?�ܤ>TGW��b$���!��{(��׻�0�f����>��T?�|r?�i�>�!n��M5;��Q�f�G=�@˽�*�Jی�� ��找��>�I�>p�=숾�ͤ���?Pp�8�ؿ j�� p'��54?2��>�?��z�t�����;_?Jz�>�6��+���%���B�`��?�G�?>�?��׾�R̼�>D�>�I�>Y�Խ����Z�����7>3�B?V��D��r�o�|�>���?	�@�ծ?li���?y�5��p��]���Z��@�'��>�9?R�
�p��>���>�C�y�u��	��Ad�v��>�s�?���?̞?p��?B��-i���c�����>�:�?/	?�)>���N�=T#8?�&��F������k�N?u�@@�MN?ű���hֿ����_N��P�����=���=Ն2>�ٽ,_�=��7=��8�B=�����=t�>��d>"q><(O>a;>��)>���Q�!�r��\���S�C�������Z�C��Xv�Xz��3�������?���3ýy���Q�2&�)?`�z��=b�U?t�Q?i6p?� ?}�y�o$ >s���e?=%�#����=>�k2?��L?y*?+��=䱝�L�d��=���o��xӇ�gm�>p�I>�t�>1E�>�	�>�<9��!J>a�>>�.�>>Z�$=1���e�=5O>�>&��>�m�>�Y<>�>[ϴ�1/��>�h���v� �˽��?>i��k�J�K3��*��׏��
��=�c.?��>���n=п����.H?����-���+�">��0?\W?�>����O T��'>���j�8U>�# �TKl���)�fQ>�e?��c>m"t>�q3���7���N�_���A�>#_4?i���?6��t��LH���YLI>yý>_�	�L[�Eܖ���~��&i��Lk=�:?��?����Cn����y��V����T>0�]>α"=tq�=LrO>?:Y�W�����F�ˎ.=u��=��W>&&?/c+>��=���>���_N�{��>��A>RK*>H�??*"%?fU��Й�B����-�O)w>��>P��>%�>KJ�x��=��>�kb>I0�����^��\�@��W>Qp����_�I<x�A�v=���c�=�D�=����*<�<'=�~?���(䈿��e���lD?S+?a �=!�F<��"�E ���H��G�?r�@m�?��	�ߢV�?�?�@�?!��P��=}�>	׫>�ξ�L��?��Ž7Ǣ�Ȕ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ\h�>ux�{Z�������u���#=J��>�8H?�V��q�O�'>��v
?�?�^�ة����ȿ9|v����>P�?���?i�m��A���@�n��>2��?�gY?�oi>�g۾�`Z���>λ@?�R?2�>�9�7�'�p�?�޶?ȯ�?�G>m��?Zs?��>�cl��..��Z���"�����=�����>���=�p����F��4��{��+�i����I"b>E�#=��>�t὞i��㰴=׫��N5��Ǆc���>n�m>�DJ>Ӥ�>?� ?yH�>.\�>�q=�:��EI��i���;[?��x?�LA�Oi�3-�=��>�cJ��Z.?ݔm?d���4F뾢��>'f?)��?KJ>?
�>�:��⓿!���־s�#>�l >�֏>
�?�7�Q����j�e�þ���>��>���� � �`H���o�
�;>��M?�+?�Ȑ=�?�J?�m�>��>k8"��|��|K���	?�~�>�\�>�X�?a�?�KL�7��A"��]ҧ���U���k>��k?xvB?Ѹ�=%ݝ�с���u'�ѣn�"�A>i	�?��w?�]��Z��>,Ԍ?1FT?|F~?���>-]W����3���8">� ?el�T-A�9�%��&�@�	?�W?P��>��y-ӽ�Lü�����<?7p[?�/&?2��a�k�ľ���<�q.�BB�{�<1q��>$C>���mF�=L>��=H�n�6&6�W�h<�Z�='>�F�=�83�Yb��=,?�G�_ۃ���=^�r�(xD��>�IL>���y�^?m=�0�{�����x��(	U� �? ��?^k�?k��.�h��$=?�?9	?p"�>K��~޾��+Pw�g}x�qw�!�>��>�l���G���ə��~F��*�Ž2�6��>ȥU>C��>C?��>�i�>���0�Z��aϾ�˾W�G���?�N3��9%���ʾz񭾹��%uO�R۾��t��G�>[Gw��<>��?�9>�&�>���>�>���>��R>39X>��e>��p>���=t�{=�#:;&u�MX?������2�z�p����W>?��d?*?Vj=�J����i(?��?�&�?Q�>ٜV�L[<���>im�>�U{�B�?�H˼X$2���=�F��;j0�^��T=>��>����`6�qP���o��w?�o)?i�0=11쾨��O�׾<��<`�?��A?EB]����2Ae��*j�״'���>ٵ��
+�>�־J�d�p�i�\������.?��C=�?$A?�׾��˾��W�6C@�*����>�D�>?e>��>��=N� ��Z��m{�C|����?�?*�>,K?�):?��Q?FwM? -�>�a�>�=���?�>g��;ޟ>���>� :?�[.?�i.?�?Y�)?{Ga>��s ��b׾&T?��?�8?]�?�?�Ċ��ٶ�)���W`���u�b��Tv=��<(н�S��e�V=h�T>�X?���8�m���Gk>�7?��>���>'���.�����<��>D�
?�I�>2 ��}r�qb��X�>0��?��|=�)>R��=H����kԺ�c�=����L�=�"���y;�><捿=� �=��s�Y������:�d�;R��<]��>h.?z%�>�J!>���r�ݾKs6�^��<��>��=%V�=v�&���t��R��o�w����>���?� �?�A�<5��=���=O������������l���>��?xJ;?Lך?�
I?LA0?/=
�2�c��Hi���ck��
?m!,?��>�����ʾ��щ3�۝?�[?g<a�����;)�5�¾��Խ��>�[/�b/~�����D� 䅻���'~����?߿�?�A�M�6�@x�Ŀ���[����C? "�>�X�>��>�)�0�g�P%��1;>��>5R?y�>9�O?�A{?��[?�vT>�8��2��w̙��5�p�!>�@?m��?���?	y?�^�>q�>��)��ྜྷB�����4�ׂ�LgW=�Z>~��>M0�>��>���=��ǽ�����>�:m�=d�b>s��>͏�>���>ހw>ҷ�<I�G?���>�Z��<��&夾)Ã��C=��u?��?�+?�=��+�E��F��E�>�n�?���?6*?}�S�L��=m�ּݶ�"�q��%�>|Թ>*�>Bϓ=�F=0m>2�>M��>���`��s8�O�M���?F?t��=.ſ�>p��l��"����B<�썾N�a�E��;�a�z��=W����#������Z�b蝾w퐾�I��/6������0 �>�X�=�*>wW�=��<�7ȼ��J<:2=Q�t<��<�y�r~F<+�<����"�}�p�J��ti<�EW=���
Wʾ~?-OH?I�>?U�H?�Ƃ>���=rsԼ��{>T	��~?v>O�9ݗ���N]�h%���G��/�˾K����`�^0���'>������>��3>�r>�{=n=�=bK=gj�=E!<���<�>��=po=J��=�J>{��=���?tȑ��ϗ�ud�9@=k?2/�>�\>'�Ͼ@�_?��>�	���<�������?7S�?K��?���>�վ��p>�H��������&>���br=�K�=�q�‾>�>Z)/��^����=&g�?�@@��0?J���Eտ�p�<#�3>{�>�R���0�FDR���T���P�Me?�=��hʾ'�>�ή=例Gƾv�#=j
;>��K=v>�t�[��3�=�z��M=��r=k{�>�E>�
�=rl��ڸ=�W?=�=W_M>�#�}�H�̽+��2=\i�=��d>�">-��>~�?�b0?sYd?E8�>�n��!Ͼ�:���B�>��=�G�>^؅=�pB>Ŋ�>D�7?z�D?s�K?H��>t=S�>��>��,�ֲm�k��ѧ�G��<$��?+Ά? Ѹ>�R<s�A�G���b>��%Ž�r?�P1?ll?��>{���߿�!�l>)�}x�'�/� �H=%J���,���������ٽ|$�=Q�>�-�>�җ>Gw>�=>o�P> �>`{2>n�K=�ڮ=��q<��Ѽ6GR=`i��_�=�
z�Z��<R�;�������2�������;F7߼X��=���>�>"�>ն=���*9>l����Q���='����A�Hf�L|�?�.���*���<>ұI>�� c����?^U>� =>���?�s?��">h��e�Ӿ\ɛ�ll]���G����=+��=�I�];:��_�+L��xѾ���>S�>F�>F�l>�	,�� ?���w=�a5�g�>�x�������:7q�o?��9���i��CѺS�D?SF�����=�"~?n�I?f�?���>�����ؾM/0>PD����=��#q�ah����?�'?�>u�n�D�d�׾�+y�x?�e���Rg�ʠ�[]�w+��~��E�?I̾�몾R�%�鉚��悿ɴ`���ǽ忪>Q~?�5�?݁���у�������̾6Α=O&+?E��?�=�@?k��>޷��l�$�z��a$=d��?��?t��?��>�j�=�����+�>�*	?��?#��?ys?cw?��P�>���;�� >����Q��=��>U�=l'�=a?�~
?��
?V\��E�	�S�����e1^��I�<̾�=�>w�>��r>�;�=0�g=���=8W\>H�>ӏ>g�d>��>I0�>�ʦ��~��5?�y=+�>]3I?���>�o	��G�=]�=��;=Nhf��쎾��߽�;��H~�=�M��-m�FJ:�l��>�{��}?�?Sl>�%��?xW�uX�A->�
>-�d�(Ũ>��>>�>/��>�W�>Q�>9?�>�ϩ=ޯپ��>J ��P���I�i�X��־�8X>c|����	�n�
��FսQ40� ��������n�������@��<<�ۍ?��#f���%�ei��?R�>S�6?x��'1��
=�=��>�>2�^E��w�����ܾ~�?7*�?`!*>��> p5?�: ?������<�^M�?|p���:�hy��`�����	���f�]�̼�*t?�Dg?{�;?\�ýBw8>%��?�.�ssy�!G�>�S�̑X�aDs=;��>�Qھ[�Ծ��3��:���2�+r=��S?S��?�0=?�{5��+4���>���>\[?h<?��>�M?l�U���F?%E�"��>��6?�'4?`�I?Y��>ײ>�ӹ����:��p>����Ő��<��~ac�Oɽek->%2�=��ߞ�=��<!.=�k���κ���=!��<q%~=Q]���=�#>dO�>��`?��>��=>U
7?�@�xyM�N��Z5?���ä�m���8���ۧ ��:�Yb?9�?�Bq?B�;>��;��+�C�,>�j#>o>,>ޮ!>��b>� ���ݽ�>�7Z>a9> B>�ս-������V��)`n=��'>l��>���=��K��S�;ͯ��J���>�sp��]�pBg���V���/�,�����>�;[?�,?���=<)
���J=����\�U?ȯ?��H?�?���=(Ѿ�.B��+���o]����>#����.�YF��^ܶ��������St>�ϾL���>�m�3�K��^q��[�)��B�������2<C���u�E:�3&>G>�����Q6�󄛿	�ȿ(vC?��=�
,��ȽG����>�B�>��>�׻=�0{��/)�f�Ǿ�ٰ�"�=u8'>0�P����I�s:�7Q�>F�>?u�w?�&{?y���]�T��#t���e��L��υ���X'?+��>;�?��=��\=K��H(��}���7�`H?�\�>��1���S������'���0����>��/?���=���>X�?��3?��?�5?��?Xxs>!ώ����N7?�h|?���<�Q��;�lF�M[�͗=?_?�D���Q=�?��Q?38?9�Z?�z	?� ���i�u�R��R�>J��>~�����}o>��V?:��>{e]?y��?�]z>+gH�ҫ���.���#->c&>D%Q?�,??S&$?I��>5��>l����i�=���>j
c?J�?`�o?��=׻?��2>&��>���=�&�>���>��?WO?�Us?B;J?'��>���<ŗ��WԲ��s�̲X��;t�<��x=f��r����6��<E�;~��:%��k�D�`���;\_�>T�v>lڕ���0>�þ���2�C>����Κ����{;�B��=4��>Cq?���>l%��b�=��>-_�>}E��p(?1<?��?�͚;Da��Yھn�R�$��>�vA?���=g�l�������t���e=An?ۣ]?�[��~���a?�[?њݾ�6�^ܺ�~z�����mX?�?� X��*�>��~?�py?���>{�E�ǭk�9ٜ�lb�v����$>B��>a�$���p�*��>w�*?6��>"��>�r>��ھsP���A���?.�?!�?�"�?&�,>Z^��*ܿ�\־f���:?��>����G@?�{��,�о�Ҿ�wm�X���&�徴��q���Ƭ�V*��ȍ��D��Lz&�/T?|�w?�%n?D%N?����\M���h�wh��ؤ<�+.����i�*���A�W�h�����-�#a�����?3�<�}���b<�C��?P5$?4�9�5f�>و��)��f�ܾ$�> 6���	�)��=*(꼐.=��b=�.h�z�;��"ž0�"?5��>:��>��@?�|[���=���2��B>���=�N>Ϡ�>ݽ�>}�>nő<Ƿٽ�����پ�.��H�g� �e>��Y?�.V?��k?k�Z�������^���\��"���=0>]/=$��><ż��\}��:���K�DGw����wь��>�1ol>��1?w�O>om�>���?ȣ?.	-�R�l�j�X�63��i��s�>�^y?��>]��>�e���$�9��>tr?���>��z>ⷡ�l)�0��YՖ���>��1>?���=��������/���ʎ�;�P�n��=�LI?�j\�
���`Ț>GY?�3�{� >�(�=x��=c��B��6������=a�?t �=:�j>�����
��wx�Ju���+?*�?\����,��P�>G
#?Ǌ�>�#�>�̈́?�$�>ߪ�� ��<Jr?\?xuG?�j@?
w�>mn�=fܽ�HԽI&�S�?=�؋>��V>�Dr=U}�=��"�l-n��U$���=���=�(>�ӎԽ�/$���f~<�Q�=�/5>�~߿�[G�V���������5��V����O:����(O�)G�� ���d�J�ټ��Gz���=5���R��χ�6�x����?n�?��X�w"�`Җ������r��:q>�tz�{b*�6���;��`D�����ގ��9�E�N��[f� ��P�'?�����ǿ򰡿�:ܾ4! ?�A ?7�y?��7�"���8�� >FC�<-����뾭����οA�����^?���>��/��p��>ޥ�>	�X>�Hq>����螾�1�<��?7�-?��>Ǝr�1�ɿc����¤<���?0�@�A?��(���ejU=A��>Β	?/�?>g1�K8���IM�>�=�?���?��M=M�W��}	��~e?��<!�F���߻I
�=�Q�=y�=���N�J>�_�>T���rA��Yܽ��4>f�>�#�j��Ў^��ʽ<&�]>7&ս� ��:b�?����T��D�T��4��_>wom?\�>�:�=�H?���?����k6���y?��@�m�?�a
?�O|�>!!ݾ�_?�?��=�bC��nf��IQ>������=���qX�1��>��>�u�>O]�\� ��襾R`�.ү=	Q�m&ÿ,%��'���/=�I.<Sa����E�y1�՟�-���!}���ֽ3a�=zX�=��e>V܂>��@>�5t>(�W?���?���>W�f>c.[�A���Ӿ(8��z���T�Z-�_�/��
p�u�ؾ_ �	��n�����DG�@!=�<�=c6R����� �\�b�`�F���.?�u$>|�ʾd�M�٫-<�oʾ{����؄�gॽ.̾�1�o"n�G͟?��A?����\�V�r��XY�m�����W?�N�s���ꬾ~��=^���f�=4%�>���=���� 3��~S��{<?�>2?���:���G`�>��4��عK�\?�`?R� �@Ό>��~?�N�=vx=:�j>��A=���>��P?;�u�_T޾~����?�c_?��>��"㾉�1?� ��̡�.r��3n=������X�>:�<�Cľ���9<½z_R>�(W?ݞ�>�)����]�����G==��x?�?�*�>�yk?��B?� �<)d����S����ow=w�W?�&i?ͳ>����оz���5?V�e?r�N>~ih�#�龨�.�OT��#?k�n?�^?�s��x}�g�� ���o6?�*}?�ix�᥿r���LZ�r�>���>:Y�>��N��r�>=_?*)�P���?a�� �.�0��?YS@=��?��=k��)B�<!��>��>#\9�R6��E	3������?=�R�>w��4��k-�!���^K?�1�?���>����
����=�=�����?Y@�?�U��HI�<s��W�k��x��,<sK�=�G>��J�1�X�8��@Ǿ���&�����Q]�>�Q@�߽d��>J<�����ο�x���Z˾�7~�?�>{W׽�g���l��u�-9H���H�ϵ��ڨ>6>bT��r��Kit�!`@��������>hz~���z>AA�M��FĄ��r�<>:c�>�7f>�zܽP�Ǿ쏚?�#�`п����q����M?�y�?9]�?��4?������=;t���D=�*T?��v?��b?g��@A��ݏ�#�j?�_��vU`���4�sHE��U>�"3?�B�>T�-�8�|=�>���>g>�#/�y�Ŀ�ٶ�A���X��?��?�o���>q��?ss+?�i�8���[����*�m�+��<A?�2>
���F�!�C0=�UҒ���
?V~0?{�a.��a?��c���r���.��ӽ�>Ay%���K�a7��M���e��圿7y�H�?�; @�³?B��-#��%$?�8�>�i���|Ǿ�K�<��>���>~X>F~�y�>g^�v�>�[{
>���?a>�?-x?Ù��-�����=v2|?��>>ӄ?�E�=^��>|;�=x���	�Y��%>n��=�}��� ?>�O?ԟ�>���=�]2�ҿ.�`)A�uUL�Æ��QD�K��>q�a?r�M?�`f>�쬽�4�/%�����,����SJ����ï׽�'2>�:J>@6>o�O��iξ��?Op�9�ؿ j��%p'��54?1��>�?��{�t����;_?Kz�>�6� ,���%���B�a��?�G�?>�?��׾�R̼�>@�>�I�>L�Խ����_�����7>2�B?]��D��t�o�{�>���?
�@�ծ?ji�� ?�K6�Jl��cB���;%�o[��5Š>�K?�n
���?�]"?ǥ>����7	����n����>`7�?��?��?R�?1I���e��e�	=�I�>��?ve�>\�=n�3�|�=��L?t��Z����ܾ��X?yt@��@�*r?#x��5�ܿ����C�����"�Z>>ү�=6�G���=R>��!��������=G�>�NX>���>GH`>�[R>�Ro>����C!$������֙��|.�R. ��[�F��0��c ���j#�{>ɾ�ɾnۻ�n#�8�4�9S佼[���a����=�U?�R?Vp?ڐ ?�x��>_����p=��#����=4�>�i2?Y�L?A�*?�̓=����d��]���A���Ƈ���>�zI>3~�>�H�>� �>qWH95�I>�,?>��>� >0Z'=t��}c=.�N>�G�>���>�z�>�D<>j�>2ϴ��1��&�h�2w�b̽W�?=���+�J��1��m9��¥���j�=^b.?�|>����>п[����2H?�����)���+�9�>��0?�cW?�>����T�H:>b��{�j�c_>=, �v~l� �)��&Q>`l?5e>�n>�7��K9�8E�)̟��
�>��-?��ƾ`"��pt�(=O�RV꾠*D>�c�>�\��H��_���y�B&q���]=Z�5?]5?�ə�����g�{��U��G�J>��k>��f=㾥=m�D>8Py�-�t'D���=\��=��S>J?��&>Q-x=���>纖��rE��@�>�TA>X�>~D@?��$?R�4��g���{��Β(��|>c��>0�>g� >�H�;H�=tQ�>��c>g�l
_��Z��E�FR>�H��iT�<߅���=*��'��=}=���2i5����<)�~?���7䈿F�h���lD?�+?� �=�F<I�"�[ ���H���?l�@+m�?@�	���V���?�@�?����=)}�>�֫>�ξm�L���?�ƽ@Ǣ��	�)#�gS�?��?��/�Wʋ�-l�6>�^%?�ӾLh�>�x�pZ�������u���#={��>�8H?uV���O�z>��v
?�?_�ک����ȿ�{v�
��>R�?���?~�m��A��@�x��>;��?�gY?�pi>�g۾�_Z��>�@?�R?'�>�9���'���?�޶?¯�?�<B>Xx�?�QN?urw>����.�����e�c�5XؼV�v�j��>x�軆�־�|p�ࣿ��y���^���	��>8��<}R�>=;=�U]�+��=~R-��̾x��=L��>F\�>���>�n�>z�?4>5>`	v>4g��C��������:���W?�X�?q
��us�� �=��=�Ʃ���1?��S?��<�����>H�l?��x?�S?}�>d6辐������u��l�n=�=f�>���>�ק=#�>ְ�e��~��>���>?�">��4�������>�68?�?G͛=�� ?�#?�l>GC�>�E�)/���F�/��>P��>��?��~??|���L53��ǒ��衿�[���K>Ox?��?���>̹��d���M�4�!1T��1��C��?�ph? H��X?�L�?U5@?�dB?�g>[���׾�x��ӿ>�?�e�cZ�Ξ'�����$?3�?��>�{��$�=�M˽B�6��� �k��>6I?��!?��u�]��˦�����g�����<��ǹ������=.^�;RƆ=�I�=h�>�U>K�����񽀲/=��>n��>�>�ѽs	���<,?y�G��ۃ���=��r�3wD�c�>FIL>����^?�j=�.�{�{��ux���U�� �?���?"k�?����h�e$=?'�?F	?k!�>�I���~޾���Qw�U�x��v�:�>���>��l���Z�������KF��N ƽ�t
��;�>�>Ϟ�>���>miu>�԰>朔�2�2���̾��r�i�����4�UT%��{�����ծM�iJx��;¾��m����>��*����>?�?�oA>}	�>��>��!=j�>�\>�/\>���>6DS>��->>�=_{4�ؑ���DR?.�����'��辘���sB?kpd?�.�>x�h�s�������?��?dp�?�Dv>syh��+�{y?)�>)5���u
?�[;=n�	�Pe�<�;��9��SZ��K����>�׽�%:�G�L��Hf��^
?�9?�ɍ�\�̾O�ֽL���<�<�z?�*?��t�V$�}]I��]�Q�/������r0	�/�8���p���w� ��oB���\8�$����?.�M?'������u�� DZ���a��>x��>��=�i�>��<��
���N��af��m,���'����>ue�?4��>��W?�`#?�Q?�>Q?9�>2��>�O��5(?I�����1>�?̮C?y�7?v�#?r>?+�$?�ލ>�VF��c��D���?�G;?z.?�-?��>q;�2�<V��=��\���ĺ�.u=���;6ې:���ti�h�t>@P?2����8�:����+k>�7?0��>԰�>>��s�Wh�<��>��
?�0�>U����ir��]�F/�>9��?cr�rI=��)>W%�=;^��ʺj��=	���E�=�����w:��"<�i�=�Ӕ=� t�
a����:�߆;N�<�s�>�?/��>�@�>&?��Ъ �=���]�=>
Y>�S>�>�Eپ�}���$��r�g�Xy>�u�?ky�??�f=��=���=Wy��=R��!��T�����<�?�J#?�XT?O��?��=?�j#?֮>�)��L��1]��M����?0!,?E��>����ʾa�n�3�b�?�Z?�<a����0;)���¾��Խϯ>	\/��.~�����D��ⅻ����|����?���?�A�/�6�Ly�w���[��o�C?m"�>�X�>��>R�)�m�g�Q%��1;>���>GR?�#�>��O?�<{?�[?�gT>&�8�K1���ә��?3���!>�@?ݱ�?��?y?Pt�>U�>��)���T��i��M�����W=;	Z>c��>i(�>��>���=Ƚ�X����>��_�=�b>7��>0��>x�>n�w>dO�<ɓI?�N�>�'ž��'���4�y�_/����y?��?C�*?��<���=��K��u�>�?���?tu*?�~b�7��=�d��}Ǵ��mj��4�>�>{�>ݼa=��<�K>���>#+�>2�"�Ə��19�V�^��h?�=L?^��=r�ſ)`q�D�p�v�����c<�Ғ��d�?a���O\����=/Θ��G�Sש�iB[�V��l3��:��E뜾�}�ɠ�>bІ=���=�O�=���<yȼK�<(�J=5�<��=��m��Yp<AV8�"j�pw��ۭ4�p_O<�:G=���L˾Fy}?�RI?�+?�C?Zz>hv>��1�@1�>���?w~U>��N�{���S�;�8����R���ؾ/e׾��c�s����>�I���>��2>_J�=E��<���=%�s=���=]uF���=G��=�H�=���=��=V>�5>�?�i��Wj�J��,D\?а�>qd�>����R?�>����4ſ���5�?���?���?��#?^���I�>	�ҽb��;X�=vG�]�%>0�=S��?�z)>pjj�}̧�Wl�>XD�?�\	@��*?gA��{�忋��<�4>c3�=��V�խ2�9�<�6�<�d�7���?5@�������t>�, =}���㿾Ľ^=�qF>"<J=��"���U�e�=�o����=��}=��}>.?K>�h=]�����=��F=f>�uO>-�F<aA���W��(9=���=�@n>�_>a��>��?�a0?�Xd?q6�>�n��Ͼu?���I�>��=�E�>�=�rB>8��>Z�7?��D?��K?6��>��=c	�>��>@�,��m�Um�I̧����<���?�Ά?@Ҹ>�Q<�A����g>��/Ž�v?RS1?�k?��>>��K,ΐ��n�+�H���\=^�������]���39�<�]���-!�=�O�>���>���>6�>WK@>�dx>�ĺ>Av+>��=�r=�˽�H��H
=O�z=箯��*ݽJŝ��vr<�ݺ\t޻��l�g�������߿���	�/��=�~�>>-�>���=	Ʋ�sT1>m���97M����=d;��H�B�Hqd���}�G�.��5���A>t�V>Z,��H��s�?�3Y>�A>Jm�?-.u?�v>j=��վX�����c�X�T�G)�=Q�>��?���;�^`��sM��Ҿy��>��>I�>��l>5,�"?�˹w=:��a5��>0z������)�.:q�@������;i�n�Ժ��D?�E�����=0"~?��I?��?���>���N�ؾ080>{D��[�=�U%q��g����?~'?r��>��G�D��庾�T��}�>vaI�c8x��S���j��N~
�#ۋ����>vN���Ͼ��9��T����*�o�� ����>�ip?9�?A�����������Z����(�~QF?c�?�O�>lyh?� ?[1D> ˾���=S�=>q?�D�?�2�?S�->~9�=�T��&��>��?h��?��?�js?��?����>��;��>#Й�+��=E>Н=/X�=�?9�	?��
?����	��ﾳ��y^�ܿ =ǁ�=�"�>{/�>)r>���=J�k=>��=y�[>�?�>�r�>[�e>ҵ�>�<�>����n��I?��4=���>�3?���>�#h=T�#�G=�=�
���p{�>^��皽���p_�=tM?;�9R=�����>Sb��8K�?^�O>�[���?rp��e�V&'>��
>����|�>���>\5M>��~>��v>y��=�Ф>_*�=�־R	>F�������E�bkQ�HҾ#�o>�0��WV7�	�	�ݐ���N�Cp�������k�`ق��>��;���?���8�i�Ė(�UK���?�0�>��5?��������Q>\�>u�>\{��zϔ�(����"�?A�?�;c>��>��W?u�?�1�3��uZ��u��(A�Ue���`�t፿���<�
�R��|�_?	�x?�xA?O�<�9z>���?_�%�ӏ�c)�>c/�R';�@<=�+�>2*����`�A�Ӿ@�þ[9��EF>�o?�$�?Y?�PV�~Б����>��?Y�}?�-�?��*?QC?E1����S?*=*��>c�/?�FC?�2M?��G>׈w>L�>fU�=��>�o������M=e�d�]w�����=͂=�����p��`�=��=z�߽�xF�zм�y<�-B�=Y�M=�*6<ڧc=��>��]?v �>�X�>��7?���8��^��j9/?�7:=ݚ��w����|��l���>��j?���?	tZ?6�c>��A�#C�6>dz�>�f&>�[>c��>I����E����=�>1�>�٤=�oN�hہ���	�P|��&��<	9>��?
>�m���n �p���V#����>�v��>�+E�j�h���?��ɸ�cu�>�qb?�n ?jr8=/Q�����5�n�9IE?<g&?��I?���?'�>��x7���f�nʽ���>rf��(E�����>��!D��μ�j�>%俾Z
��_C>I=m��mR��J�� 6j��0���*]�����/�>����s�F���I(�=<q�>����u ��ț�J���*�M?�2�ϭ;�t���(��g=�31>o�>ؑQ�(�F��9�v�I>��>��#>.Z�Z5�z�?��Ѿt�|>-�C?��f?_Ĉ?��U�Z?_��\J�:xܾ�c�����'!?E^�>�q	?�O>b= u¾��	�z�Z���8�A|�>U�>:2���@� ���Ɂ�A&�n�>^F?p�>�a?�W?N?�k?��,?H�>�1s>UGw��n��*B&?��?��=�Խ��T�- 9��F� �>ۃ)?��B�̸�>~�?=�?*�&?�Q?۵?N�>� ��C@����>QY�>��W�zb���_>��J?V��>�<Y?�ԃ?m�=>c�5�ꢾ�ة��T�=�>��2?"6#?ï?`��>g��>G���u�=���>�c?�0�?�o?���=&�?�:2>R��>���=���>S��>�?OXO?(�s?��J?Ǒ�>���<�7���8���Cs���O��ɂ;�pH<Y�y=����3t�.K�,��<d �;�g���H�����l�D��������;g��>�cy>z���K�.>��������dF>�4����M~��U�5��=��>�?�ђ>��)����=��>=��>Y* ��B*?s�?�?���;��`��j׾�=W���>��A?���=;6j�V��R�u���a=y`m?�~\?Mjb�����,6k?z�B?IT����$���־|+M��)��߭}??t�/��>���?6�?[� ?)�
�,(p��謹��@�Y�����5>�A0>xNP�<�q�JuU>�=?�U?���=V�>J 辰����L���?2�?��?��?�{�=��~��׿�]��4��MU?fH�>[>��Z�/?�'�9u־�r��3@�Ǿ<ޱ������l�������w�����9������<�?*9n?Դm?�]?���]�%ae��r�VN��M�K�$4F���D��1?��b����ei۾ �q��[�=����&�4�?�U2?㹾��m>�������Ꮌ��d�>��s�Hf���O�=״;�&�>LU<O�<� �o������x6?b�>fg�>� -?��f��]=��0���;�%� �G��>"]�>���>L;�>�=��㒅<��'_־G8���q�N�k>(c?��N?@q?Y���S(�ń������t����dL>5z>��>�sh��e0��^&�)�:��-n�����<��c��Ϧ=��5?w��>ݚ�>"��?"u
?>�&r����b���0�b׶<���>�Cg?�|�>F҉>�ڽ+S!�c��>�ol?��?.�#>>�߽b������#	���>�"3= �?7',>�	L�n�r�nў� ����$��c�>q�g?t$���^���U�>"�y?|��|>ft5>�;> 6��{�x� �҉�>F��>ς|=�ō>$���tVƾ��q�QӴ��O)?�K?J꒾�*��6~>$"?R��>�.�>I1�?�(�>qþ{�@�ұ?0�^?.AJ?�SA?H�>3�=���aAȽ�&�Ф,=���>��Z>7m=�}�=����t\��v���D=�p�=�μ�M����<�����K<���<��3>���QI?�����s�Ӿ^����
��Yn��Q�3q\�b�������Qv�OD\�=w���g�0�h��o*��w�����B�?i��?>�Ƚ���+\��W~������u>])o�}��='Ɛ�jȽ�����q"\�M/���2��`�&�m�U�'?�����ǿ𰡿�:ܾ*! ?�A ?<�y?��4�"���8�Z� >D�<0+����뾠�����ο(�����^?m��>��Q/��f��>ѥ�>ǡX>�Hq>����螾m/�<��?,�-?��>��r�*�ɿc���9Ĥ<���?,�@�A?��(�y����T=���>2�	?`�?>@�0��4����<O�>�:�?M��?*ON=�W���	�xpe?l�<� G����#,�=:i�=<a=H���SJ>Z�>r����A���ܽ�4>�҅>�#�d��(�^�@E�<P�]>�sԽ������?�u����q�K�o~n��Ӑ>Ի_?���>��>��?PH:�����B���I?��@ǁ�?Z�?�
&���>1�Y�<??��3>n�@�H;v��CK><����=\��3y�f{�>���>St�>�ɽ�x�\^���Ľ���>Z��3Ŀ��.����D=�8����?3��u���]�󢏾�nR���ͽ��=�g�=��'>��>�QZ>�~E>�"[?��}?��>4J>�*�WH��:`ξr����|�#潞so�F�Ľ�&������cھ� �B��mm���!=���=7R�f���C� �c�b�J�F���.?�v$>U�ʾ��M���-<pʾS���rۄ��ॽ�-̾�1�*"n�k͟?��A?������V�]���W�����K�W?P�ͻ��ꬾ��=x���V�=%�>ኢ=���� 3��~S�N�1?`5?F
��ƹ���>�A.�i�n=��C?g��>l*���>Ȍ8?�d=B�0>���=��<�A�>L?Ls�=�(�0���&?[K?/;�)�;���>����ܿ��?C=���=��V�dU">{z�>�]$=G8ھ`v�<�*<T�j>�!W?���>@�)��
��P�����V�<=��x?r�?��>�yk?��B?��<>k����S���Pw=��W?�!i?��>p�����Ͼ.���q�5?u�e?��N>]hh�u�龡�.�EM��-?o�n?�X?x��� y}�!������n6?�K�?��w�"㞿T�������>�Y�>\�?c!=�{��>��i?�M>������~���P'���?�x@��?��=�N���|O=��>���>��_q��`e��G����=9]�>�KL�Z|`�Z�(�Q|��jH?��?�~�>�Ȏ�yE-����=�ٕ��Z�?|�?v���wHg<M���l��n���~�<�Ϋ=+��F"������7���ƾ��
����9⿼ͥ�>BZ@�U�w*�>�C8�Y6�TϿ'���[о�Sq�u�?,��>t�Ƚ����7�j��Pu�L�G��H������k�>��>�X��؛��	w���9�_j��tC ?����_>,2%�^✾#&���G=^3�>-s�>�R>c���*q��� �?.g ��*ҿϤ�������Q?���?댄?a�'?����ݑ��r�a�}4=�<P?hs?�\?ܞ��I@d��$���j?W_��xU`��4�FHE�<U>�"3?%C�>D�-�°|=�>���>�g>^#/�_�Ŀ�ٶ����R��?͉�?�o���>m��?~s+?�i�8��B[����*��+��<A?�2>����!�0=�+Ғ���
?>~0?�{�O.���_?<�a�d�p�R�-��ǽ '�>��/��[��H���-��e��	���ly�ԭ?>d�?�?d��&#��$?Ւ�>C���=Ǿ���<X��>��>��N>÷`�U-v>1�M;�ڟ	>J��?�a�?�g?D���� =>�~?氒>!h�?��<��?��>vپ:[>�e>��=A���*��>��U?�?�ܤ>TGW��b$���!��{(��׻�0�f����>��T?�|r?�i�>�!n��M5;��Q�f�G=�@˽�*�Jی�� ��找��>�I�>p�=숾�ͤ���?Pp�8�ؿ j�� p'��54?2��>�?��z�t�����;_?Jz�>�6��+���%���B�`��?�G�?>�?��׾�R̼�>D�>�I�>Y�Խ����Z�����7>3�B?V��D��r�o�|�>���?	�@�ծ?li���?y�5��p��]���Z��@�'��>�9?R�
�p��>���>�C�y�u��	��Ad�v��>�s�?���?̞?p��?B��-i���c�����>�:�?/	?�)>���N�=T#8?�&��F������k�N?u�@@�MN?ű���hֿ����_N��P�����=���=Ն2>�ٽ,_�=��7=��8�B=�����=t�>��d>"q><(O>a;>��)>���Q�!�r��\���S�C�������Z�C��Xv�Xz��3�������?���3ýy���Q�2&�)?`�z��=b�U?t�Q?i6p?� ?}�y�o$ >s���e?=%�#����=>�k2?��L?y*?+��=䱝�L�d��=���o��xӇ�gm�>p�I>�t�>1E�>�	�>�<9��!J>a�>>�.�>>Z�$=1���e�=5O>�>&��>�m�>�Y<>�>[ϴ�1/��>�h���v� �˽��?>i��k�J�K3��*��׏��
��=�c.?��>���n=п����.H?����-���+�">��0?\W?�>����O T��'>���j�8U>�# �TKl���)�fQ>�e?��c>m"t>�q3���7���N�_���A�>#_4?i���?6��t��LH���YLI>yý>_�	�L[�Eܖ���~��&i��Lk=�:?��?����Cn����y��V����T>0�]>α"=tq�=LrO>?:Y�W�����F�ˎ.=u��=��W>&&?/c+>��=���>���_N�{��>��A>RK*>H�??*"%?fU��Й�B����-�O)w>��>P��>%�>KJ�x��=��>�kb>I0�����^��\�@��W>Qp����_�I<x�A�v=���c�=�D�=����*<�<'=�~?���(䈿��e���lD?S+?a �=!�F<��"�E ���H��G�?r�@m�?��	�ߢV�?�?�@�?!��P��=}�>	׫>�ξ�L��?��Ž7Ǣ�Ȕ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ\h�>ux�{Z�������u���#=J��>�8H?�V��q�O�'>��v
?�?�^�ة����ȿ9|v����>P�?���?i�m��A���@�n��>2��?�gY?�oi>�g۾�`Z���>λ@?�R?2�>�9�7�'�p�?�޶?ȯ�?�G>m��?Zs?��>�cl��..��Z���"�����=�����>���=�p����F��4��{��+�i����I"b>E�#=��>�t὞i��㰴=׫��N5��Ǆc���>n�m>�DJ>Ӥ�>?� ?yH�>.\�>�q=�:��EI��i���;[?��x?�LA�Oi�3-�=��>�cJ��Z.?ݔm?d���4F뾢��>'f?)��?KJ>?
�>�:��⓿!���־s�#>�l >�֏>
�?�7�Q����j�e�þ���>��>���� � �`H���o�
�;>��M?�+?�Ȑ=�?�J?�m�>��>k8"��|��|K���	?�~�>�\�>�X�?a�?�KL�7��A"��]ҧ���U���k>��k?xvB?Ѹ�=%ݝ�с���u'�ѣn�"�A>i	�?��w?�]��Z��>,Ԍ?1FT?|F~?���>-]W����3���8">� ?el�T-A�9�%��&�@�	?�W?P��>��y-ӽ�Lü�����<?7p[?�/&?2��a�k�ľ���<�q.�BB�{�<1q��>$C>���mF�=L>��=H�n�6&6�W�h<�Z�='>�F�=�83�Yb��=,?�G�_ۃ���=^�r�(xD��>�IL>���y�^?m=�0�{�����x��(	U� �? ��?^k�?k��.�h��$=?�?9	?p"�>K��~޾��+Pw�g}x�qw�!�>��>�l���G���ə��~F��*�Ž2�6��>ȥU>C��>C?��>�i�>���0�Z��aϾ�˾W�G���?�N3��9%���ʾz񭾹��%uO�R۾��t��G�>[Gw��<>��?�9>�&�>���>�>���>��R>39X>��e>��p>���=t�{=�#:;&u�MX?������2�z�p����W>?��d?*?Vj=�J����i(?��?�&�?Q�>ٜV�L[<���>im�>�U{�B�?�H˼X$2���=�F��;j0�^��T=>��>����`6�qP���o��w?�o)?i�0=11쾨��O�׾<��<`�?��A?EB]����2Ae��*j�״'���>ٵ��
+�>�־J�d�p�i�\������.?��C=�?$A?�׾��˾��W�6C@�*����>�D�>?e>��>��=N� ��Z��m{�C|����?�?*�>,K?�):?��Q?FwM? -�>�a�>�=���?�>g��;ޟ>���>� :?�[.?�i.?�?Y�)?{Ga>��s ��b׾&T?��?�8?]�?�?�Ċ��ٶ�)���W`���u�b��Tv=��<(н�S��e�V=h�T>�X?���8�m���Gk>�7?��>���>'���.�����<��>D�
?�I�>2 ��}r�qb��X�>0��?��|=�)>R��=H����kԺ�c�=����L�=�"���y;�><捿=� �=��s�Y������:�d�;R��<]��>h.?z%�>�J!>���r�ݾKs6�^��<��>��=%V�=v�&���t��R��o�w����>���?� �?�A�<5��=���=O������������l���>��?xJ;?Lך?�
I?LA0?/=
�2�c��Hi���ck��
?m!,?��>�����ʾ��щ3�۝?�[?g<a�����;)�5�¾��Խ��>�[/�b/~�����D� 䅻���'~����?߿�?�A�M�6�@x�Ŀ���[����C? "�>�X�>��>�)�0�g�P%��1;>��>5R?y�>9�O?�A{?��[?�vT>�8��2��w̙��5�p�!>�@?m��?���?	y?�^�>q�>��)��ྜྷB�����4�ׂ�LgW=�Z>~��>M0�>��>���=��ǽ�����>�:m�=d�b>s��>͏�>���>ހw>ҷ�<I�G?���>�Z��<��&夾)Ã��C=��u?��?�+?�=��+�E��F��E�>�n�?���?6*?}�S�L��=m�ּݶ�"�q��%�>|Թ>*�>Bϓ=�F=0m>2�>M��>���`��s8�O�M���?F?t��=.ſ�>p��l��"����B<�썾N�a�E��;�a�z��=W����#������Z�b蝾w퐾�I��/6������0 �>�X�=�*>wW�=��<�7ȼ��J<:2=Q�t<��<�y�r~F<+�<����"�}�p�J��ti<�EW=���
Wʾ~?-OH?I�>?U�H?�Ƃ>���=rsԼ��{>T	��~?v>O�9ݗ���N]�h%���G��/�˾K����`�^0���'>������>��3>�r>�{=n=�=bK=gj�=E!<���<�>��=po=J��=�J>{��=���?tȑ��ϗ�ud�9@=k?2/�>�\>'�Ͼ@�_?��>�	���<�������?7S�?K��?���>�վ��p>�H��������&>���br=�K�=�q�‾>�>Z)/��^����=&g�?�@@��0?J���Eտ�p�<#�3>{�>�R���0�FDR���T���P�Me?�=��hʾ'�>�ή=例Gƾv�#=j
;>��K=v>�t�[��3�=�z��M=��r=k{�>�E>�
�=rl��ڸ=�W?=�=W_M>�#�}�H�̽+��2=\i�=��d>�">-��>~�?�b0?sYd?E8�>�n��!Ͼ�:���B�>��=�G�>^؅=�pB>Ŋ�>D�7?z�D?s�K?H��>t=S�>��>��,�ֲm�k��ѧ�G��<$��?+Ά? Ѹ>�R<s�A�G���b>��%Ž�r?�P1?ll?��>{���߿�!�l>)�}x�'�/� �H=%J���,���������ٽ|$�=Q�>�-�>�җ>Gw>�=>o�P> �>`{2>n�K=�ڮ=��q<��Ѽ6GR=`i��_�=�
z�Z��<R�;�������2�������;F7߼X��=���>�>"�>ն=���*9>l����Q���='����A�Hf�L|�?�.���*���<>ұI>�� c����?^U>� =>���?�s?��">h��e�Ӿ\ɛ�ll]���G����=+��=�I�];:��_�+L��xѾ���>S�>F�>F�l>�	,�� ?���w=�a5�g�>�x�������:7q�o?��9���i��CѺS�D?SF�����=�"~?n�I?f�?���>�����ؾM/0>PD����=��#q�ah����?�'?�>u�n�D�d�׾�+y�x?�e���Rg�ʠ�[]�w+��~��E�?I̾�몾R�%�鉚��悿ɴ`���ǽ忪>Q~?�5�?݁���у�������̾6Α=O&+?E��?�=�@?k��>޷��l�$�z��a$=d��?��?t��?��>�j�=�����+�>�*	?��?#��?ys?cw?��P�>���;�� >����Q��=��>U�=l'�=a?�~
?��
?V\��E�	�S�����e1^��I�<̾�=�>w�>��r>�;�=0�g=���=8W\>H�>ӏ>g�d>��>I0�>�ʦ��~��5?�y=+�>]3I?���>�o	��G�=]�=��;=Nhf��쎾��߽�;��H~�=�M��-m�FJ:�l��>�{��}?�?Sl>�%��?xW�uX�A->�
>-�d�(Ũ>��>>�>/��>�W�>Q�>9?�>�ϩ=ޯپ��>J ��P���I�i�X��־�8X>c|����	�n�
��FսQ40� ��������n�������@��<<�ۍ?��#f���%�ei��?R�>S�6?x��'1��
=�=��>�>2�^E��w�����ܾ~�?7*�?`!*>��> p5?�: ?������<�^M�?|p���:�hy��`�����	���f�]�̼�*t?�Dg?{�;?\�ýBw8>%��?�.�ssy�!G�>�S�̑X�aDs=;��>�Qھ[�Ծ��3��:���2�+r=��S?S��?�0=?�{5��+4���>���>\[?h<?��>�M?l�U���F?%E�"��>��6?�'4?`�I?Y��>ײ>�ӹ����:��p>����Ő��<��~ac�Oɽek->%2�=��ߞ�=��<!.=�k���κ���=!��<q%~=Q]���=�#>dO�>��`?��>��=>U
7?�@�xyM�N��Z5?���ä�m���8���ۧ ��:�Yb?9�?�Bq?B�;>��;��+�C�,>�j#>o>,>ޮ!>��b>� ���ݽ�>�7Z>a9> B>�ս-������V��)`n=��'>l��>���=��K��S�;ͯ��J���>�sp��]�pBg���V���/�,�����>�;[?�,?���=<)
���J=����\�U?ȯ?��H?�?���=(Ѿ�.B��+���o]����>#����.�YF��^ܶ��������St>�ϾZ
��_C>I=m��mR��J�� 6j��0���*]�����/�>����s�F���I(�=<q�>����u ��ț�J���*�M?�2�ϭ;�t���(��g=�31>o�>ؑQ�(�F��9�v�I>��>��#>.Z�Z5�z�?��Ѿt�|>-�C?��f?_Ĉ?��U�Z?_��\J�:xܾ�c�����'!?E^�>�q	?�O>b= u¾��	�z�Z���8�A|�>U�>:2���@� ���Ɂ�A&�n�>^F?p�>�a?�W?N?�k?��,?H�>�1s>UGw��n��*B&?��?��=�Խ��T�- 9��F� �>ۃ)?��B�̸�>~�?=�?*�&?�Q?۵?N�>� ��C@����>QY�>��W�zb���_>��J?V��>�<Y?�ԃ?m�=>c�5�ꢾ�ة��T�=�>��2?"6#?ï?`��>g��>G���u�=���>�c?�0�?�o?���=&�?�:2>R��>���=���>S��>�?OXO?(�s?��J?Ǒ�>���<�7���8���Cs���O��ɂ;�pH<Y�y=����3t�.K�,��<d �;�g���H�����l�D��������;g��>�cy>z���K�.>��������dF>�4����M~��U�5��=��>�?�ђ>��)����=��>=��>Y* ��B*?s�?�?���;��`��j׾�=W���>��A?���=;6j�V��R�u���a=y`m?�~\?Mjb�����,6k?z�B?IT����$���־|+M��)��߭}??t�/��>���?6�?[� ?)�
�,(p��謹��@�Y�����5>�A0>xNP�<�q�JuU>�=?�U?���=V�>J 辰����L���?2�?��?��?�{�=��~��׿�]��4��MU?fH�>[>��Z�/?�'�9u־�r��3@�Ǿ<ޱ������l�������w�����9������<�?*9n?Դm?�]?���]�%ae��r�VN��M�K�$4F���D��1?��b����ei۾ �q��[�=����&�4�?�U2?㹾��m>�������Ꮌ��d�>��s�Hf���O�=״;�&�>LU<O�<� �o������x6?b�>fg�>� -?��f��]=��0���;�%� �G��>"]�>���>L;�>�=��㒅<��'_־G8���q�N�k>(c?��N?@q?Y���S(�ń������t����dL>5z>��>�sh��e0��^&�)�:��-n�����<��c��Ϧ=��5?w��>ݚ�>"��?"u
?>�&r����b���0�b׶<���>�Cg?�|�>F҉>�ڽ+S!�c��>�ol?��?.�#>>�߽b������#	���>�"3= �?7',>�	L�n�r�nў� ����$��c�>q�g?t$���^���U�>"�y?|��|>ft5>�;> 6��{�x� �҉�>F��>ς|=�ō>$���tVƾ��q�QӴ��O)?�K?J꒾�*��6~>$"?R��>�.�>I1�?�(�>qþ{�@�ұ?0�^?.AJ?�SA?H�>3�=���aAȽ�&�Ф,=���>��Z>7m=�}�=����t\��v���D=�p�=�μ�M����<�����K<���<��3>���QI?�����s�Ӿ^����
��Yn��Q�3q\�b�������Qv�OD\�=w���g�0�h��o*��w�����B�?i��?>�Ƚ���+\��W~������u>])o�}��='Ɛ�jȽ�����q"\�M/���2��`�&�m�U�'?�����ǿ𰡿�:ܾ*! ?�A ?<�y?��4�"���8�Z� >D�<0+����뾠�����ο(�����^?m��>��Q/��f��>ѥ�>ǡX>�Hq>����螾m/�<��?,�-?��>��r�*�ɿc���9Ĥ<���?,�@�A?��(�y����T=���>2�	?`�?>@�0��4����<O�>�:�?M��?*ON=�W���	�xpe?l�<� G����#,�=:i�=<a=H���SJ>Z�>r����A���ܽ�4>�҅>�#�d��(�^�@E�<P�]>�sԽ������?�u����q�K�o~n��Ӑ>Ի_?���>��>��?PH:�����B���I?��@ǁ�?Z�?�
&���>1�Y�<??��3>n�@�H;v��CK><����=\��3y�f{�>���>St�>�ɽ�x�\^���Ľ���>Z��3Ŀ��.����D=�8����?3��u���]�󢏾�nR���ͽ��=�g�=��'>��>�QZ>�~E>�"[?��}?��>4J>�*�WH��:`ξr����|�#潞so�F�Ľ�&������cھ� �B��mm���!=���=7R�f���C� �c�b�J�F���.?�v$>U�ʾ��M���-<pʾS���rۄ��ॽ�-̾�1�*"n�k͟?��A?������V�]���W�����K�W?P�ͻ��ꬾ��=x���V�=%�>ኢ=���� 3��~S�N�1?`5?F
��ƹ���>�A.�i�n=��C?g��>l*���>Ȍ8?�d=B�0>���=��<�A�>L?Ls�=�(�0���&?[K?/;�)�;���>����ܿ��?C=���=��V�dU">{z�>�]$=G8ھ`v�<�*<T�j>�!W?���>@�)��
��P�����V�<=��x?r�?��>�yk?��B?��<>k����S���Pw=��W?�!i?��>p�����Ͼ.���q�5?u�e?��N>]hh�u�龡�.�EM��-?o�n?�X?x��� y}�!������n6?�K�?��w�"㞿T�������>�Y�>\�?c!=�{��>��i?�M>������~���P'���?�x@��?��=�N���|O=��>���>��_q��`e��G����=9]�>�KL�Z|`�Z�(�Q|��jH?��?�~�>�Ȏ�yE-����=�ٕ��Z�?|�?v���wHg<M���l��n���~�<�Ϋ=+��F"������7���ƾ��
����9⿼ͥ�>BZ@�U�w*�>�C8�Y6�TϿ'���[о�Sq�u�?,��>t�Ƚ����7�j��Pu�L�G��H������k�>��>�X��؛��	w���9�_j��tC ?����_>,2%�^✾#&���G=^3�>-s�>�R>c���*q��� �?.g ��*ҿϤ�������Q?���?댄?a�'?����ݑ��r�a�}4=�<P?hs?�\?ܞ��I@d��$���j?W_��xU`��4�FHE�<U>�"3?%C�>D�-�°|=�>���>�g>^#/�_�Ŀ�ٶ����R��?͉�?�o���>m��?~s+?�i�8��B[����*��+��<A?�2>����!�0=�+Ғ���
?>~0?�{�O.���_?<�a�d�p�R�-��ǽ '�>��/��[��H���-��e��	���ly�ԭ?>d�?�?d��&#��$?Ւ�>C���=Ǿ���<X��>��>��N>÷`�U-v>1�M;�ڟ	>J��?�a�?�g?D���� =>�~?氒>!h�?��<��?��>vپ:[>�e>��=A���*��>��U?�?�ܤ>TGW��b$���!��{(��׻�0�f����>��T?�|r?�i�>�!n��M5;��Q�f�G=�@˽�*�Jی�� ��找��>�I�>p�=숾�ͤ���?Pp�8�ؿ j�� p'��54?2��>�?��z�t�����;_?Jz�>�6��+���%���B�`��?�G�?>�?��׾�R̼�>D�>�I�>Y�Խ����Z�����7>3�B?V��D��r�o�|�>���?	�@�ծ?li���?y�5��p��]���Z��@�'��>�9?R�
�p��>���>�C�y�u��	��Ad�v��>�s�?���?̞?p��?B��-i���c�����>�:�?/	?�)>���N�=T#8?�&��F������k�N?u�@@�MN?ű���hֿ����_N��P�����=���=Ն2>�ٽ,_�=��7=��8�B=�����=t�>��d>"q><(O>a;>��)>���Q�!�r��\���S�C�������Z�C��Xv�Xz��3�������?���3ýy���Q�2&�)?`�z��=b�U?t�Q?i6p?� ?}�y�o$ >s���e?=%�#����=>�k2?��L?y*?+��=䱝�L�d��=���o��xӇ�gm�>p�I>�t�>1E�>�	�>�<9��!J>a�>>�.�>>Z�$=1���e�=5O>�>&��>�m�>�Y<>�>[ϴ�1/��>�h���v� �˽��?>i��k�J�K3��*��׏��
��=�c.?��>���n=п����.H?����-���+�">��0?\W?�>����O T��'>���j�8U>�# �TKl���)�fQ>�e?��c>m"t>�q3���7���N�_���A�>#_4?i���?6��t��LH���YLI>yý>_�	�L[�Eܖ���~��&i��Lk=�:?��?����Cn����y��V����T>0�]>α"=tq�=LrO>?:Y�W�����F�ˎ.=u��=��W>&&?/c+>��=���>���_N�{��>��A>RK*>H�??*"%?fU��Й�B����-�O)w>��>P��>%�>KJ�x��=��>�kb>I0�����^��\�@��W>Qp����_�I<x�A�v=���c�=�D�=����*<�<'=�~?���(䈿��e���lD?S+?a �=!�F<��"�E ���H��G�?r�@m�?��	�ߢV�?�?�@�?!��P��=}�>	׫>�ξ�L��?��Ž7Ǣ�Ȕ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ\h�>ux�{Z�������u���#=J��>�8H?�V��q�O�'>��v
?�?�^�ة����ȿ9|v����>P�?���?i�m��A���@�n��>2��?�gY?�oi>�g۾�`Z���>λ@?�R?2�>�9�7�'�p�?�޶?ȯ�?�G>m��?Zs?��>�cl��..��Z���"�����=�����>���=�p����F��4��{��+�i����I"b>E�#=��>�t὞i��㰴=׫��N5��Ǆc���>n�m>�DJ>Ӥ�>?� ?yH�>.\�>�q=�:��EI��i���;[?��x?�LA�Oi�3-�=��>�cJ��Z.?ݔm?d���4F뾢��>'f?)��?KJ>?
�>�:��⓿!���־s�#>�l >�֏>
�?�7�Q����j�e�þ���>��>���� � �`H���o�
�;>��M?�+?�Ȑ=�?�J?�m�>��>k8"��|��|K���	?�~�>�\�>�X�?a�?�KL�7��A"��]ҧ���U���k>��k?xvB?Ѹ�=%ݝ�с���u'�ѣn�"�A>i	�?��w?�]��Z��>,Ԍ?1FT?|F~?���>-]W����3���8">� ?el�T-A�9�%��&�@�	?�W?P��>��y-ӽ�Lü�����<?7p[?�/&?2��a�k�ľ���<�q.�BB�{�<1q��>$C>���mF�=L>��=H�n�6&6�W�h<�Z�='>�F�=�83�Yb��=,?�G�_ۃ���=^�r�(xD��>�IL>���y�^?m=�0�{�����x��(	U� �? ��?^k�?k��.�h��$=?�?9	?p"�>K��~޾��+Pw�g}x�qw�!�>��>�l���G���ə��~F��*�Ž2�6��>ȥU>C��>C?��>�i�>���0�Z��aϾ�˾W�G���?�N3��9%���ʾz񭾹��%uO�R۾��t��G�>[Gw��<>��?�9>�&�>���>�>���>��R>39X>��e>��p>���=t�{=�#:;&u�MX?������2�z�p����W>?��d?*?Vj=�J����i(?��?�&�?Q�>ٜV�L[<���>im�>�U{�B�?�H˼X$2���=�F��;j0�^��T=>��>����`6�qP���o��w?�o)?i�0=11쾨��O�׾<��<`�?��A?EB]����2Ae��*j�״'���>ٵ��
+�>�־J�d�p�i�\������.?��C=�?$A?�׾��˾��W�6C@�*����>�D�>?e>��>��=N� ��Z��m{�C|����?�?*�>,K?�):?��Q?FwM? -�>�a�>�=���?�>g��;ޟ>���>� :?�[.?�i.?�?Y�)?{Ga>��s ��b׾&T?��?�8?]�?�?�Ċ��ٶ�)���W`���u�b��Tv=��<(н�S��e�V=h�T>�X?���8�m���Gk>�7?��>���>'���.�����<��>D�
?�I�>2 ��}r�qb��X�>0��?��|=�)>R��=H����kԺ�c�=����L�=�"���y;�><捿=� �=��s�Y������:�d�;R��<]��>h.?z%�>�J!>���r�ݾKs6�^��<��>��=%V�=v�&���t��R��o�w����>���?� �?�A�<5��=���=O������������l���>��?xJ;?Lך?�
I?LA0?/=
�2�c��Hi���ck��
?m!,?��>�����ʾ��щ3�۝?�[?g<a�����;)�5�¾��Խ��>�[/�b/~�����D� 䅻���'~����?߿�?�A�M�6�@x�Ŀ���[����C? "�>�X�>��>�)�0�g�P%��1;>��>5R?y�>9�O?�A{?��[?�vT>�8��2��w̙��5�p�!>�@?m��?���?	y?�^�>q�>��)��ྜྷB�����4�ׂ�LgW=�Z>~��>M0�>��>���=��ǽ�����>�:m�=d�b>s��>͏�>���>ހw>ҷ�<I�G?���>�Z��<��&夾)Ã��C=��u?��?�+?�=��+�E��F��E�>�n�?���?6*?}�S�L��=m�ּݶ�"�q��%�>|Թ>*�>Bϓ=�F=0m>2�>M��>���`��s8�O�M���?F?t��=.ſ�>p��l��"����B<�썾N�a�E��;�a�z��=W����#������Z�b蝾w퐾�I��/6������0 �>�X�=�*>wW�=��<�7ȼ��J<:2=Q�t<��<�y�r~F<+�<����"�}�p�J��ti<�EW=���
Wʾ~?-OH?I�>?U�H?�Ƃ>���=rsԼ��{>T	��~?v>O�9ݗ���N]�h%���G��/�˾K����`�^0���'>������>��3>�r>�{=n=�=bK=gj�=E!<���<�>��=po=J��=�J>{��=���?tȑ��ϗ�ud�9@=k?2/�>�\>'�Ͼ@�_?��>�	���<�������?7S�?K��?���>�վ��p>�H��������&>���br=�K�=�q�‾>�>Z)/��^����=&g�?�@@��0?J���Eտ�p�<#�3>{�>�R���0�FDR���T���P�Me?�=��hʾ'�>�ή=例Gƾv�#=j
;>��K=v>�t�[��3�=�z��M=��r=k{�>�E>�
�=rl��ڸ=�W?=�=W_M>�#�}�H�̽+��2=\i�=��d>�">-��>~�?�b0?sYd?E8�>�n��!Ͼ�:���B�>��=�G�>^؅=�pB>Ŋ�>D�7?z�D?s�K?H��>t=S�>��>��,�ֲm�k��ѧ�G��<$��?+Ά? Ѹ>�R<s�A�G���b>��%Ž�r?�P1?ll?��>{���߿�!�l>)�}x�'�/� �H=%J���,���������ٽ|$�=Q�>�-�>�җ>Gw>�=>o�P> �>`{2>n�K=�ڮ=��q<��Ѽ6GR=`i��_�=�
z�Z��<R�;�������2�������;F7߼X��=���>�>"�>ն=���*9>l����Q���='����A�Hf�L|�?�.���*���<>ұI>�� c����?^U>� =>���?�s?��">h��e�Ӿ\ɛ�ll]���G����=+��=�I�];:��_�+L��xѾ���>S�>F�>F�l>�	,�� ?���w=�a5�g�>�x�������:7q�o?��9���i��CѺS�D?SF�����=�"~?n�I?f�?���>�����ؾM/0>PD����=��#q�ah����?�'?�>u�n�D�d�׾�+y�x?�e���Rg�ʠ�[]�w+��~��E�?I̾�몾R�%�鉚��悿ɴ`���ǽ忪>Q~?�5�?݁���у�������̾6Α=O&+?E��?�=�@?k��>޷��l�$�z��a$=d��?��?t��?��>�j�=�����+�>�*	?��?#��?ys?cw?��P�>���;�� >����Q��=��>U�=l'�=a?�~
?��
?V\��E�	�S�����e1^��I�<̾�=�>w�>��r>�;�=0�g=���=8W\>H�>ӏ>g�d>��>I0�>�ʦ��~��5?�y=+�>]3I?���>�o	��G�=]�=��;=Nhf��쎾��߽�;��H~�=�M��-m�FJ:�l��>�{��}?�?Sl>�%��?xW�uX�A->�
>-�d�(Ũ>��>>�>/��>�W�>Q�>9?�>�ϩ=ޯپ��>J ��P���I�i�X��־�8X>c|����	�n�
��FսQ40� ��������n�������@��<<�ۍ?��#f���%�ei��?R�>S�6?x��'1��
=�=��>�>2�^E��w�����ܾ~�?7*�?`!*>��> p5?�: ?������<�^M�?|p���:�hy��`�����	���f�]�̼�*t?�Dg?{�;?\�ýBw8>%��?�.�ssy�!G�>�S�̑X�aDs=;��>�Qھ[�Ծ��3��:���2�+r=��S?S��?�0=?�{5��+4���>���>\[?h<?��>�M?l�U���F?%E�"��>��6?�'4?`�I?Y��>ײ>�ӹ����:��p>����Ő��<��~ac�Oɽek->%2�=��ߞ�=��<!.=�k���κ���=!��<q%~=Q]���=�#>dO�>��`?��>��=>U
7?�@�xyM�N��Z5?���ä�m���8���ۧ ��:�Yb?9�?�Bq?B�;>��;��+�C�,>�j#>o>,>ޮ!>��b>� ���ݽ�>�7Z>a9> B>�ս-������V��)`n=��'>l��>���=��K��S�;ͯ��J���>�sp��]�pBg���V���/�,�����>�;[?�,?���=<)
���J=����\�U?ȯ?��H?�?���=(Ѿ�.B��+���o]����>#����.�YF��^ܶ��������St>�Ͼ8���sH>�
�h_�KUq�5NK�h޾�$�={���<��1�̾�����.�=j,>�о�H!�������G?���=eߒ���G���'J$>��>�Ԣ>ᾋ���o�a�=�@>���ٟ=�^�>��,><#���"��d�P�����1��>cF?��^?��?�l��|r�tvD�����᣾`Ļx?'m�>m�?͡;>ٓ=֗���_�/8d��F�6B�>��>ۉ���I�����}y��'�$�݊�>9�?��>P?�S?��?�`?�T+??���>�D��I߷�_&?���?gc�=-v̽�9L�r�9��E��@�>��)?\yI��>��?BS?�(?��Q?��?�>Jf ��5A���>A��>��U��ᮿ֚O>�J?�W�>�xU?�B�?�%@>�24�Ձ�������=��'>E�.?�B(?)�?�N�>�p	?����D8�>#f?|{?�.�?=��?C��>�I�=	���R>��!=�h[>�`/?�IX?K�?.A�?&m|?��>���<c*����=h� ��;5��;��<�б=B�v�0.>C�<f�8RP=�A�=(�=�%$>΂��)�޽�
9�y^�>E�s>5��}�0>�ľD����@>4Z��lN���̊�g�:����=D��>U�?���>[V#�y��=I��>?C�>���&(?=�?�?�q+;W�b���ھ��K�P�>�B?<�=2�l�����h�u�1�g=��m?o�^?ˀW������c?��T?�����^��ZӾ\�d�T ¾v�T?���>vz�8�>E=a?s��?�N�>�O��1Xs�X���Ld���f�y��=�|>�����g���>O�>?�E�>��v>�	�=��徍�M��������>j�?3��?�Ѕ?k;>��c�ڿ(���=}���$_?,"�>�o�� �$?����J;"㈾�8��|Sھ�ǧ��B���r��E᥾0"�r���1�н��=d�?�s?��o?4a?s����c��]�򅀿�V����U���+E���C�C���n�K�5����}����L=NA� kS��ҿ?�?9M����#?�����tžɭ��l.>e٦������[�
�f<�(�<�r�=��[���Ƚ$1��1I?��>~޻><�Q?`@H�(�6���<�<iB�v�徖]/>���>r�>4��>n�l���?�9K۾[9|�����Ţ>��s?@�0?+U?@�>S=G�]&����־$��=#�<&7>��j>5��>� 	���~�ɾ�I���i����lTu��a�pM'=5�#?k�<�Ę>��?Qu ?[p����O�c��1�w�.=��?��`?���>|�?�@��v��P��>��l?�f�>k��>O@���w!��]|�{�ͽ��>J?�>���>W�q>��+���[�<-��K���Q9�pr�=,h?fY��(�`��>��Q?�}�:�Q><��>l�m�+k!��9�/�'��]>�~?\;�=4�<>�xľ����{�ս��4�-?M�?\Z��%7�/\�>?�)?7^?j�>	?qk�=����">��#?$�`?6�R?mZT?>�?��>'���s����G� �=�%>�j>Iѽ=(>֔'�}��B�� >��>'歼L��f!��&!=B����^g�g
j>Ǝٿ%iQ����E���g���s�M�Y�d���7��:ɾҠ���ۏ�L4�H�較.|�g�Y�Ռ��f��u�?{��?-!a��>���%r���߾�̮>� ��kk���)���f׽�p��Á㾽"��-�(���V���n��2\��I3?K���� ʿ����N��YG?��*?LR?b	'��$�&�E�-�y�p>������#�䖿G�ƿ��8�i?^w�>�Y�NkC��n?��>���>��m>|ë�M���|Eݽ�i�>��?�(?#�9���"�����~�?�@PzA?٢(�R�쾈�U=��>�f	?Le?>��0��,��>���=�>&�?V��?�P=�W�c7��Le?��;s�F�؇���=�j�=�=���+K>5Г>�?�
�A���ڽ�5>s��>+�#�p��r�]����<��^>��ս����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=s6�䉤�{���&V�}��=[��>c�>,������O��I��U��=����\ſ��W�_�(�����Q���@ �����=��>�ņ��&ξ{L�lC���l&�3>���=5�`>��=�0>��S?�Z?^��>BC#>ZT��$���T��aC�=4E��mW��ν�S����鮾��
�Ⱦz�2��N!�1q	���d�Q^?�q�M=}JR�#䏿$�-d�.DC��X/?ʲ->�PѾ��O��Z�<u�о垰�'uT��ǽ��˾}&0���i��[�?��A?W�����R���h�߼
�����R?�8�>��j��<�=LY��¸�<{�>�g�=�46�#O�'1?9$? ��������5> �׽�~x=�:4?�|�>�KûT�>��'?���×���p>L�]>�Ϯ>�)�>/�>׍������=�?U�T?����hܑ����>Uߴ�p!o��n�=>r�A�KQ�~"V>dT7<!n��.���|<
'W?ٍ>`�)����x����?=�x?��?E��>Nk?WC?ެ�<���_�S�B�
���y=��W?�i?��>W����оy�����5?��e?�N>�h��A�?�.�u$��I?��n?[c?h���G}��#��Q���|6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������6A>}-}��%�?�6�?Ciھ��q>�C��$��1�;=�I>��?�X��*���̾�B�x҃�6h��'�����=>H]>�	@.ꮾ�0?�,<.�G�ƿ�j���d����=�s�>���=��Ҽ�+��R��Jx��QS�0�T�ʡ��d�>�'>���,���F}���;�)��a��>��*���>J]Z�uķ����K��;~��>+k�>`,�> ���q-���ܙ?�8����οI8��*�)QY?��?�5�?ZV?Pu�:[�{�D`x�&>h��K?8s?��W?c�'���]�ͼV�A�e?���	=[���,����HyB>��6?��l>$L�v
Q>`��<���>�ԙ>XB�Ejǿ����!��d�?��?��a?ki�?~v#?x�3�W3��@��>l��L��ΈC?�6@> )�G%����F�o�fF�>��*?�!���.�\�_?)�a�L�p���-�f�ƽ�ۡ>��0��e\�_N�����Xe����@y����?N^�?i�?õ�� #�f6%?�>d����8Ǿ��<���>�(�>
*N>mH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?/�>��?
��=�$�>���=����;���">���=�z?�K�?r�M?�U�>���=��8��/��ZF�*%R��$��C�E��><�a?1lL?��b>c���U2�� �x�̽�1�����@�s+� �߽��5>�%>>g�>��D���Ҿ��?3p�/�ؿ�i���o'��54?e��>��?'��}�t�^���;_?�z�>7�,���%���C�/��?�G�? �?m�׾�N̼6>}�>�I�>��Խt���J���(�7>��B?���D��U�o�w�>���?�@�ծ?(i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*�wȿN0���8�^Q˾#��=c��=��|>�x�<��Ҽbw7=�[=�Җ=�H�=>$�>aFf>!J>V�>b#{>H!���N���Z!��$��TY����B��X��"-�V➾D����_�_��yM��^�e��G��r�"�ϙ��r�E��1� )	>��S?�KM?�bm?|E�>@�P�*>~��m��<�C:�g��=�c�>��.?�|T?/�,?/��=�ƅ�v$c������f���@��L��>_t>ɀ�>�%�>|g�>�Q0;��'>q�M>��>�{Y=�g��9�,� `�<��/>=<�>t��>�>��J>'\>����a[��+�f��Pt��y�� T�?|��t�D�C0�������H�� ��=_%?9�=W���Ͽ������E?�B�����R'���>�H1?��T?�p>����Y�w�`�/>8]���u���	>�I��Ya�a&%��E>��?�a>*Fe>٩5�Y?�NRO��Z����>&4?��2�-��%q���E��BվNCM>F�>م!����f���L�w�K>c���]=��3?ݲ?I��㤾@�o�yD��)bS>j�Y>!u=�*g=U#3>�\���hݽ4�=��Z=���=�6i>�T?��+>��=��>r0����O�Й�>q�B>>�+>��??�%?�R�����J���~-��Ow>Qd�>��>�2>U\J�|L�=�]�>�a>7�PI���C��e?�QEW>_�|�dp_�'�v�x=�O��(��=ה=�y �|�<�4�%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾC�>�M��Ǉ���������ң+��p�>,�B?'���pr=ᓋ����>�$?���}K��< ǿ ���ڝ>���?ף�?Kwi�����m���?T��?�'l?r�>�뾭枾��O>��/?�YS?
V?j���)��b?xw�?�#Z?�J�>��?}\I?��>��">��M��ɿ�{��+?X>��߽a��>d@�>���Sq.�\=|��uj�ǀc�z��P�½:��<UY�>�����"�>	u�l���|v[����>AA�=����#>��?�=�>\�>s>�=�2�)�߽�H��|�J?u�?r
�?�e�wr�<k�L=mc����>�)?[]Y�TOþ�f�>6}^?���?�Y?��>���ka������w��/w����Q>^f�>���>�n=<���>�����Z�͒�>��>�k��V꾭�h��<��>�3?���>�{=w�?J�<?��{>/�>�K������Z�c��h�>@?��?���>�)���y?�m��R��PTU�u3�=6\M?xX-?���>���R�����<U���g�����?�!H?�uԾ~�n>~��?�?�?M?l=�>e����%�d��=��T>�&?<��NGI�=�I��u?Lk? �>�������|���$�/�ξR�?�C?@?�Q��e��ž���<�����hA=؂=[�+>T�>�޽�m�=
>��>e�����]�B`��Tv�=���>���=�&I�tL7�/=,?�G�ۃ���=��r�?xD���>�IL>����^?ol=��{�����x��	U�� �? ��?Zk�?b��?�h��$=?�?S	?l"�>�J���}޾6���Pw�~x��w�\�>���>�l���K���ڙ���F��]�Ž�N����>���>MT	?���>�CA>���>�A����#�;��N�	�3aX�G���7�;�+�[9 ���a�9�@�̼��Ǿɹr�^��>Dq���&�>?�b>��|>	�>!	7����>�8>�g>���>���>�&>q'>b�P=�<��%�R?R�6�)�I���a���L;@?.d?���>B�-v���9�e�?��?5�?K�f>��h�`,�2?��>?m|���?&@=P?Z���<l���n�G���^T��h�>�:���;��,N�rb��	?��?��Y�az;ޡսN��%y�=Cɇ?��)?����S2�.%R�C�[���j�@�o=`����'��f�����t��"��M���
�"�4X��B?���?���� �D�-�}��e�A�Z:�=�3?�l?C0?���>�^ �#�+�Lň�S���P,�-�>�?'�>9?K�*?��Z?�;5?�4�>���>eO2��7�>�f�����>2K�>t�?�G<?Yj5?�8?I�7?�S3>~�b��t���?�?�/?H�?yp#?�4?�O����!��s=�Կ�V�ܾH���!��>�S��Bνd۟:n�>M^>�"? ����B�h�
h�>�=0?
�?��>����jS��[���{r>�++?�g�=T{!���O�>]&�WT�>?�?�9��U�u=��v>:>��<�왼���=���lf�-��=Ň归ĭ=K�=��d='�g<��#>����p=��=u�>d�?L��>RE�>�@��7� �Ҷ��Y�=�Y>\ S>P>�Eپ�}���$����g��[y>�w�?ez�?r�f=1�=���=1~��iV��6������e��<��?�I#?�WT?[��?y�=?�i#?��>�*�TM���^��8��B�?.�0?"O�>rC�٬ھG��S��8=? �>�jh��X��y�%��l��f=~��;�!H�*�l��o��$]I�%"r>�3
���,�ZQ�?�Ǚ?��ؼ�U.�\5�o����<��k{>?���>���>�m�>��(�)�U�����HL>���>�WP?���>�7d?�c?�|7?���>B�;�C��������>�'c=ej1?ts�?�<�?G�Q?��>�>ԓ��\#�����e����|�N�a>��a>���>g��>���> m=�A*�B+�u�ʌ!>"Y>"��>�w�>���>0`d=ˀ�=jH?'l?�։�9�Ɓ����W#�=u��??5�?�''?�`��t��)5��ϵ��`?|�?��?DZ?�Ź��Z�=�Q=�A��G���>�w�>lR�>#Q�=�k�=f�)�?ʒ>W��>K��<���P1�%���?�ng?	C>����߮S�jvi�/�I�����Ӿ� �]�<�0>#�>=~#���>5"�������dD��uP��e�^�����>>��'>��>(X >�(�=�[����:�+������=��'>Bg��#��= ��=�ط�F��=�p�=�J>L�.��6˾�)}?�"I?S�+?��C?0�z>�>P�/�S:�>����4?*�T>�T�c'��@�:�8j�������eؾWr׾�d�a����>��H���>ww3>���=�-�<�R�=h�s=��=B�f�'=��=cE�=���=d��=�G>�>�6w?O�������4Q��Y罨�:?�8�>B{�=��ƾ`@?V�>>�2������db�.?���?�T�?Y�?)ti��d�>L��X㎽�q�=!���>2>���=}�2�0��>��J>����J��
����4�?��@��??�ዿɢϿka/>[>�(�=�hO���8�ֵ����k���8���?g�.��4���e>�۪=��;濯���<�:�=/|=��A���M����=����=�<�1�=���>��T>���=�\��6�=z�=��@>��%>×�9��E��i�L�=�v>>~k>�X5>�^�>ֻ?W�2?][]?�Q�>(&$�������I�6�>'��>X��>8
C� �d>�m?�+T?�g?��R?0��>��z��>,�>V�<�Oj�F�ھ.����=c�}?t(�?��>r5��Y�+�}�!��f6��J˻�(�>0D?H�?N >ڽ��lۿdg9�3�)�]�Z���4��8{������o0��&��݆&�?yE��r��*�>���>p��>{7�>��U>�ޡ=���>T�=Y�=}��=�=�;~� a�<r(-=���%������ͽ�0�=ߑ��ԽX��>։=�Q����=@��=j��>�?>��>/��=h��,</>�����L��ɿ='X���#B�'d��G~��/���6���B><X>Bc���2����?�Y>�W?>��?X@u?��>�c�վ�N��Re�gbS����=+�>]�<��z;��N`�W�M���Ҿ���>|H�>6'�>��C>d����I�q�.=�澐{D�Q?��׾��=��d=$Oq�Z��������Y�=�}�<=V??�� f4>��?0=&?�:?��>�VF��������>Y���z�(�ɾ����j8¼ňh?�{v>n3?N��`o�'�̾����M�>W�I��*P������R0����w���Y�>��IϾ�d3�?J������B�%r�6�>Y�O?���?ݽa������N��r�������?��f?,�>�?\�?���������~��ظ=D�n?���?�?�?n�	>��=������>�?ޕ?�?�?�Hr?�a3����>c���>Ӓ���8�=Rm>�V�=���=v�?m�
?A?�j��h�	��꾠VS���=��=��>��>��u>��=B�H=/?�=5�Z>���>c�>�^>�.�>�C�>r�&J�}�H?6/ =MA!>��b?i�>+��=�UӼ���<&I>x����?�=7����(�8��<�^;=�.=#?��ֿW��?�bn>kU=���\?߾]$6= O>��=;5'>GO�>q�.�E^�>"8t>;S�>ɦ2��J�>}`>O�Ѿ�>~���!�C�_+R��о��x>A��:1#�@��I���?F�o���}	��j��(���=����<��?\�����k��7)����V;?el�>�Z5?�Ì��(��h�>,��>�P�>�������i���Q�ᾇ��?��?�<c>!�>��W?��?��1�U3�ZuZ��u�6(A� e���`�c፿������
�����r�_?��x?yA?�@�<:z>9��?�%��ӏ�S)�>&/��&;��@<=�+�>z'����`��ӾݸþA7��JF>��o?�$�?Y?�TV�x0�'� >
�C?�>?0p?g�=?>�2?��/�L�?��>�6�>I��>�s?�g8?O?��d>2:>ҝ�;�����#_�Z�꒻��⽼W����=^1F�!�*��<�q�=�BQ=|;�<�V><X8=4�'=A
p=�G�<W�>Y�|=ߪ>��Y?���>�Y�>��??q���)�g�����$?'�<˻�����������߾@+>��p?#��?ʠd?p�`>�9�E�E�	e>��>e*>��o>F�>�j�� oY�ξW=�#>F)>���=y{��?v�q�� ��+F�;u8>b�>M}> j����*>����w�d>�JR������}U���F��m1���u����>��K?Ug?l��=ڋ�T����e�U�'?�J<?U�M?X5?圡=�bؾ��8���J�w$�ß>��Z<�&
�墿�����Y:�	8 ;Քw>䄝��䠾2\b>�����޾O�n��	J��Q�5EQ=��!�Q=��
־E�}��2�=j(
>����'!�e���q����$J?��h=����U�]���7�>�=�>+��>_�>�Ղv��T@� i��?�=���>'�;>�������G�99�D�>$eE?Mf_?of�?ؕ��5�r�#C���������T���Xm?s#�>C�?�,B>Am�=�����(�q�d�GHF�4��>Y�>�����G�vl��ɬ��0<%�F7�>�h?m8>8t?��R??�`?��)?��?��>�!����A&?���?�Ӑ=��ܽ��4��6�dI��#�>bR/?�2���>�u?G?�i&?��N?�{?���=����0A�X��>1Ǉ>5{W�<'���xb>��I?1�>�gS?l��?RO>)�6�ei��޵���> |B>x�5?��?�7?�ϩ>�,?r��o�>�!'?Ͳ�?�-�?
dh?��#=��>��?&�>f�>�Q���>A>l�?G|>?��??Wp?�N>*�x=��&�T��<�cڽ<Q��R�� ��<��,���1�5�p=�����h>�t�=a3�=�0=��=��F>�6>#�>9��>N�n>�Ǜ�8/2>��Ⱦ���JfH>����u}��R���	4����=/߀>�� ?qӊ>�+���=�G�>s��>���&?�Z?�,?2ƅ;�b��0��T�b��>�	A?¹=}�g��rxw�� x=��h?�K^?CM�Ғ�	�X?lXw?�Ĵ�_'$�+#e������P��!?2x,?���y�g>�n?@�o?���>�U���]�������8��Ñ���=x��>�&��Py���>�.?rD�>!B>- �=dI��fC�����T?��?_��?�5�?�M�=񇆿��ԿV����d�X?���>mԾ�3(?_ṼL����zb��{��1�Ǿ!���Nj�����������iW���f���2>�&?t^�?Qzj?�Qt?0:�Dl�O������Z�xc���Ծ"�@��oW���?�7�|�\�3����>���:<�>i�f_�"��?�#?ʇt��%?C���z��o��.��=(�����&���=�q�<�#/=�R�=�TD�d&��~7��ǅ?���>j��>Q?ʈQ���.�»��Q@�� ��]>���>{T�>��>?�=�n�$����оͤ������v>޸c?fK?�[n?(���81�ፂ���!��'��䧾y0A>DK>X$�>2�V����&��N>���r����7��w�	�F{=�52?�)�>;�>O3�?�?4V	�譮���x�2�1��b�<�Ժ>�Hi?Я�>v�>�ҽ� ����>��l?���>��>�̋���!�f�|�ݬнN��>��>�P ?!s>�,�ī[����+B����8����=�Ch?�΃�fu^��Ą>�P?���;U�O<���>mt��( �t���*�Y+	>��?�Ш=6j;>��ľ�Z��Vz��H����*?td&?���E|���>]�?2�>���=�S�?�-�>�{ᾡfм:+?(I�?c?�;;?�h�>�ˠ�Cc�!��6W4�h�G�GJ�>'*<>t0=���=�=����M��^�,=��=O"���hG�=t��=�7<F钽t&M>�tݿ�&M�e޾�������p�����;���V\}��"�R6��Q���b���R����9�l���n�v����LA�nS�?��?��l��f�5z���Ɂ�'(�~�>�2��B�������a"��%�����޻��-��U�&�c�m2`�n5?KA��;�̿x��gԾt?N~%?�Tv?A�}�$�pB!�F�=���<��74޾72��ο�X����\?�{�>r��zʽ4��>���>�va>��>�K���燾/=$�?��?�O?��<�P�ſ�����=E��?j,@6}A?^�(�����6V={��>Y�	?8�?>�P1��G�����U�>i;�?>��?
uM=��W���	�b�e?�@<:�F��sݻ��=�@�=C=����J>iU�>Q���UA�R7ܽ��4>Dڅ>�e"�ѡ�x~^�eh�<6�]>f�ս�5��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=s6�󉤻{���&V�}��=[��>c�>,������O��I��U��=����ſ,k;�YY4�!��E�Ƚ�we��>`_'�Wu�������FK=���=�H"���V7>�J>�W>Ƹ�>��F?�V?���>�z�>/��+���W��p�P;}����Ұ�oڷ�W����c3��߾���|�#����x�U�e�?��{=��R�{���!�(�a��:D���0?Q�#>~}о �N�m �<�Jþ�C��k਼g����X̾hl0��k�g|�?�0??�䅿qoT�����(�����V?� �~������d��=�����W�<B��>���=����2�oZP�l|0?�e?&^��[&����*>�� ��/=�+?\�?7�]<���>Q;%?+�*�4�㽴�[>�N4>��>lq�>�>����	[۽��?~T?���+휾,ߐ>f-��� {��_=>�N5��R�[>��<vÌ�U�0Ґ��G�<�(W?���>��)���aa�����[X==��x?��?.�>m{k?��B?U֤<h���S���7aw=�W?(*i?��>�����	оo���C�5?ݣe?��N>�bh����-�.�oU��$?�n?4_?|��w}�w��w���n6?o�v?�h^��l������V��>�>G^�>���>�9�y}�>��>??#�I��ﺿ��P4��ƞ?��@ߋ�?l1;<8��=�<?�X�>E�O�D3ƾ�l���}��^Wq=�>g~��bhv����:,��~8?z��?��>>���ǥ�˿�=&Ϝ��ȧ?��?�F��>%p󾃥��Tf޾�1�=��>���wꕾD؎�\"I������Ͼј����%>��k>TG@2[R����>�Wɽ������|��`����sx=] ?[�>6�s�}�޾��_�}����0I�XH�ilL���=>����a�2 ��wV�g뮽�~?���ʕ=\AJ�. [�n� ��}ٽ�$>�ʫ=c{�=S8���T��O�?���}ڿ�X���ʾ�@a?���?Ղ�?�?x���ru���o ��J�=�>e?*"�?|�~?����b�A���7�{*f?OI���Zd��2���E�7�H>}6?M��>=4���y=��>���>m[>$�%���ÿ�.��h	��n�?i)�?�����>m��?�W3?/���}���𸾴�*�\�
��GC?��">��� �#�I�@��]��9 ?�0?����.#�]�_?)�a�M�p���-���ƽ�ۡ>�0�f\��M�����Xe����@y����?N^�?i�?յ�� #�e6%?�>d����8Ǿ��<���>�(�>*N>YH_���u>����:�
i	>���?�~�?Qj?���������U>
�}?Z$�>��?�m�=�a�>�c�=���-��j#>M!�=L�>�ˠ?�M?�K�>%X�=��8�`/�[F��GR�G$�&�C���>��a?�L?�Kb>���T"2��!��sͽc1��W�%W@���,�1�߽�(5>��=>6>��D��Ӿ��?Np�9�ؿ j��&p'��54?2��>�?����t�k���;_?Vz�>�6��+���%���B�]��?�G�?<�?��׾�R̼�>8�>�I�>R�Խ����Z�����7>-�B?R��D��v�o�u�>���?	�@�ծ?di��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?lQo���i�B>��?"������L��f?�
@u@a�^?*!�׿����	ھ��}'�+�>:]�>!g>&��=�������\>�b>�m>��=���= �G>�;F>�H!>=������������b�n�!�(_��1ϼv��������G?�
����=�MB���t��+G������탾���=��W>ӝZ?�H?6o?W?Y�Ͻ��>��׾ �b=t�.j�<xW[>�<?��??�@?��N>�5O�F�g��������T����d�>'�>-��>8�>��>���=>�e=�/G>�ح>�W�=��X�![	��y�:>GT�>�:%?��>���=��=���������a�bߐ����=�-�?jf���]��ꂿ5�Ӿ@Ep�=V�<��!?�sM�F����꼿�
��!z=?�z����5���
��ʩ>V�A?8.H?2�= 𾈺�<_)q>$G�� �(>>�lB�hyɽ�54���޼<%�>1_d>��q> 6�֨9�JP��s��9-�>rX6?l���?�=�l
s�	J�W�۾�XM>(��>� ������疿�|��xf�5�y=>W8?�?>�������Hu��מ�8?R>��^>�+=�A�=�$K>�]��ѽ��H���E=���=o�`>�?�d->�ȝ=|w�>[u���L�Ę�>M�=>��(>8oB?�$?o��m���/����#�ȃ>�Q�>ޒ�>+��=�wG�F��=��>�:[>[W�%���Y�w�;�1�X>�r~�/Y��.q���r=AH�����=Y��=���
�9���-=�~?���(䈿��e���lD?S+?] �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l�6>�^%?��ӾxK�>�k�_W��H����u���"=���>�9H?�`��P���=��t
?�?4e�襤���ȿ�wv�;��>-�?
��?��m��C���@��t�>���?�xY?��i>�K۾��Z��u�>��@?u
R?�3�>*�SQ'���?�׶?���?��p>Ex�?q�}?�!?�S/��5�nW��?��N�>�q�|?1[�>�����A+�K���Do��'Q���-�>Jg�=�>�3F���޾��>�[�����P�Q�	?ȓ>�������>��?�y�>��>�PD=���	$�B�޾.�K?Z�?䴾ی��I�>���ξ�p=T#k?Y>�=��)�p9>*�O?�\�?bt�?�
?� ��W��Mm��A-`��܎�8�3>���>?�m>/��٧>l�/�C殾p��=|1�>���ZKҾa���C�<�]�>��?8�>�-½�?��+?W%�>%_�>�xA��6���fX�d�K>���>9	?���?X?�1ؾD\�!b��@ߖ���`���a>�Tv?��?���>w��	��%ZO>���Bh��i�?��l?tq��'Z ?�@�?�/C?jo?o>[|2�Y��X�H>�v8>�K?*��+,S���0�Bf�\�?;�?��>[��+���e<�d'� �޾qy?Z�L?��?;j�s]a��Y����=�k������_�)=�;G��r0>J/9>ai���Y�=�>���=�]~�(����/N=�=��>�G>H^%��ݔ�D,?b`D������[�=7�r�gbD�H�>�OL>������^?p
=���{�����x����T���?4��?�h�?;����h�_=?��?w�?��>5��!l޾s���sw��ox�/b���>��>�f���􉤿� ?��bƽ��Y�DI�>2U�>��>f��>@>|Ҷ>٧U��y�������_�Z��*<�x�$�80�,��<ˇ�UB	��J�$�;S��IW�>�_�+R�>Q�'?�L>(�>�V?W��$E�=l�>+	�=*�>fO�>qZ�>y<�={>��)�4DR?������'��������Z,B?�zd?P7�>V8j�������`?���?br�?��u>Kwh�V++��\?JT�>���l
?��:=Ku�9��<�i������$��@r����>�X׽�:��M��vf��Y
?J?�j���̾{a׽+��*�\<�m^?���>� 9��3~�7���z�b���C�Sڤ=�:��r�����ꯐ����p�KC��V��)t>��+?�,�?t�O�ι��)����K�tJL��<�n<�Y�>���>�/\>�D����t�<�^�R�-F��r�>�1@?/�>I?��8?��T?h�S?d��><ݨ>� �����>GF;b7�> )�>�+?�)?��6?�??G�*?�<I>��=������澻#?��?�}?��
?��?�i��r�!�C;�T<CZ����½86C=�-.�U�Q�B�Rk>C,�>�� ?��+��!v�N� >D�#?zQ.?���>���N���:7>:#�� ?%��>��9Q����p_1>��?�T <l�=A�r>�π>��,��ꏻ�>7����,<�4�<�Ľ�Ȳ��v>��#>h�<�<��>�]�����=-w�>\�?��>�F�>�=��]� ����e�=Y>�)S>%>*Dپ`~���$����g�_ny>y�?6z�?T�f=��=��=�z���T��������.��<E�?�G#?�UT?���?A�=?�i#?�>�*��L���]��J���?�^!?�]|>�P"�X�Ⱦ�飿g�+� ?H�?k�s�,k��Xb��� �n�$�A	B>_Q<���u�#���@�K��'�=��-�`�f��??ե?o�Խ	�I��Q�Ф��R:��=�I?�B�>�ܭ>F �>��8��O]�1w%�4vj>=K�>��?v��>�\?��o?7�I?
�>�1�3�������ܴ=�YC>�&?��s?�{�?�3w?��>̌>�nE�� ־������i,�A�����<�Y>Ǝ�>���>��>�u�=��J�d콿�`�(�=�\�>�a�>T%�>�»>��'>Z�����H?6H�>7̴�iN�Ӝ�q���9O���n?���?d�/?��=N�_G�qa��2��>��?8;�?|A+?Ya_�'�=�1t�n���PXv���>!��>ͭ�>'��=�Jc=�>M6�>2�>�<�y��'6���ټl�?�C?�s�=�ǿe�r��݀�䠾&Y@;�R��a�X�x�=�M�S�R�L=�1����ѽ���y^�����t������+^���Yq����>��V=>��=���=�̆<�x'���s;��I=�͠<���<�r��8H�<h���c�����Y9�;<�W1=�}<�˾ُ}?�;I?˕+?��C?/�y>4;>�3�I��>䆂��@?3V>��P�ڈ��م;����u ���ؾVx׾��c�?ʟ��H>baI���>�83>�G�=�K�<F�=s=|=/ R�d=$�=�O�=�h�=i��=0�>]U>�6w?S�������4Q�|Z罣�:?�8�>n{�=��ƾv@?��>>�2������}b��-?���?�T�?@�?Dti��d�>I��u㎽�q�=J����=2>q��=x�2�I��>��J>���K��5����4�?��@��??�ዿ̢Ͽ/a/>ƻ�=H��=�h`��<��nG��{>��B�4o&?z�>����*�F>]������o���1<�=K�=�B���9�+N��j�=�ǽu�R���@=mC�>�9�>�k�=�4ƽ� >��=�n>��%>�j<]o»�ڪ�c��=��>��\>��r>�Z�>�[?��/?�Ca??�>�OZ���m�ľ��>�ER>`��>���=d��=c��>�;?�+R?�c?m��>$<'$�>ޱ>�#)��h����d�����<]��?$f�?��>0s	=ɾ�í�+>D��}ʽ&?W+?R#?b(�>�U�����Y&�d�.�ʎ���6��+=�fr�JU���(s����P�=,o�>���>��>�Ry>��9>u�N>��>k�>�&�<�v�=���;��<Z,�����=e���m�<6�ż���[�%�u�+�D����;�{�;ڌ]<M�;�:�=A��>ٓ
>���>�<q=����5>U:��O�K��:�=Ӫ���E���e�`Gy���-��J��A>�G>^�ͽ�����>�:s>5>@��?B�v?��>��׽n1��랞�p����!��c�<$>D_ɽr}1��)Z�"�=��d�(��>�s>�N>���>}�2�m�D��G�=��ؾ�K���>�9y��H�;��< ]��K��	�����N������'?�ꇿo�=�k�?/<L?'d�?^~�>+�%���־�>N8���E���վg�ɾm^(���,?��?��>�,��:�u��� �鈉��T�>�����/Z��K�Mj�ۉ��>��u��EY��$��͑������g�à|��2�>�AS?�*�?�!*� w��7c�y��+�3�?���?`��>_x�>��>����̢�����G*>6T?m��?Vt�?>�=� >�B��%�>w�?>Θ?T�?�[r?�0,��P�>��<��(>�og����=�a�=��=fO�=[�?M~?�?:��<I���پ��8=k��@5=ʤ�=#��>i2j>��u>18�=bK�=/��=�	q>r�>�Ӈ>��>9_�>�p�>k7���<N��
?jWC<>�=�uY?�z>�Ɛ>+؜={����R��1������~߿�T�[=�"2>�~=?*s>�6���>MS���:�?�{M>�E�l�E?�侫=�^t>,3X=1�L>���>� �>�q�>��8=�>��=c�_>�a?C�Ӿ+Z>����!�/&C��[R��HѾ�i{>����cQ'���#6��8FH�g���i���i�$&��'/=�`��<��?R���טk�E�)�،���1?й�>6�5?U���ֈ�j�>7��>���>�n��cp��ᝍ���� ݋?���?�@c>\�>-�W?Z�?��1��3��qZ�!�u�r&A��e���`��ߍ�`����
�=𿽟�_?G�x?�xA?z��<�6z>Y��?(�%��֏��%�>/�8%;�5M<=P/�>p*����`���Ӿ�þ�@�KF>��o?$�?�X?OV�D�k�cK'>��:?t�1?+Pt?��1?~t;?�����$?{�3>G1?�i?�;5?~�.?��
?9Q2>��=qǡ���%=���抾�ѽDsʽ���,<4=�R{=T�J<��=��<%�aټ��#;�u����<�U:=M��=���=#>�>�X?�?m��>\	1?{㸽�e�;ኾ.e?q�t>���bjs����J����7>��?�B�?�[?a2>��/�O� ��U8>��p>M�>�i>W��>�f���s�>~{=zM>��*<���=���=�@��P��5����:�~>(��>7^|>�ď���'>�Q����z���d>u\Q�}���vS�r�G��2�1�u��t�>�K?W�?4�=��������f���(?js<?v�M?x�?��=��۾�9��J���^��>X�<�4	����Qn�:�J�
;)t>z���4D�uĂ>H�O�T}��#���u�^�#�f�$��h�.m��p����OU��7�>�>�>�Ծ���@���;ҿ���F?zE8>\��f������X֗��>E�?)`���#-�I�/�qn��Ҵ�=Aj�>0tA>�k�<,~о�:�~c��B�>�E?�d_?L`�?vpr�ӊB�����t>����Ƽg�?�y�>L4?>C>���=Vȱ�f���pd���F����>��>H��jH�iX��������$�B�><b?d!>��?�mR?g?k�`?�)?$?���>����\I����&?�S�?�D�=��н�g\��b8�h�B�UY�>M�*?��.�O��>�{?�V?�b'?�^R?��?�>f���Ho>�!��>�0�>��Y��y��P]>AxG?K�>��Z?�݄?�=>8��e������?/�=<�">7{4? �%?O�?��>#g?uѾNŉ=�?�"n?T�?K��?�ͳ��߽>��>bl�>�>8�>>{?�^?ͫ5?6�?:@^?��?Uo<H�����A�ս�pՋ�nd���G���A���<��w��R���1�=��2��|�=#����0������Vg�>�t>�땾�31>��ľ�Q����@>����E��)����:�-[�=\��>%?F��>�#�ɀ�=!n�>��>����(?!�?�5?Y;F]b��sھ8L��>�,B?(G�=\�l��o���u�#�g=�m?ɷ^?bW�R ����b?	^?=���<���¾gd�bO�e�O?V?��K���>��~?�'q?�%�>zVe��m�l���b�1Ij����==ٛ>���d��H�>�N7?@w�>�Sc>D~�=��ھOlw����L?��?-�?5܊?E�*>��n�V�߿y���I���	^?���>K1���#?������Ͼ1S����f�I'��y&���:��5|����$��Ń���ֽ���=)�?�	s?�[q?��_?ɬ �t�c��*^����I_V�+-��#��E�^"E�r�C�+�n�`���f�K�G=?�O��$~��2�?t>(?�(`�o ?�������雾�5>v����r5�}�>6��=ʍ�-eo>H�pe��T���?�[�>�*�>�!B?gyL�Ð$��t<��LY���ʾ5��>�_?ٟ5>���>>�=��\��kü�̾������=�>O�h?�	)?�:S?ʛ��җ5�����,ƾ귻=�	�Ʋ.:�x>�%->'H7��<�]��GUK�	�k�`�����_��r�?��=fS?n�=S��>���?.��>}�8�hf=�B���>�ӳ>��%?�b]?���>o#?�$S�����3�>�[u?��>���>XsC�,9&��ہ����T�>J�>ߑ�>㹕>Yu���g��s���^����C��<�=,cR?$�`�}�g��Ra>ƹF?/���J�;s�>���=ߤ�3�	�q�o��V=���>a��=3m�>����`������Z����1?ڿ?꒠�>�$�8�>�Q ?X��>�>=��?��>�派�W�=I?(B?�0P?�2Q?|��>�>�W#�OSŽ$&�N=ď�>��>B��=!=/�D�X\V�22�%1�=���=Uߏ�}I��^B=W�;�N���@�Ͱ:>4@濙�@�q]���
�N��̴��d���ϙ�vx�� �7V��tƑ��q����Ľ�M��i����V���1�����?}��?AP!� l���ƕ�fy�Mi��>�K�L�Z<�`���;�:~��'Ӿ�������	};��ȅ��V���$?D��-dɿ}��վ<1?�� ?,:y?�1���$�Gr4��Q�=vɡ��<_�0���t���cϿ6R���U?v��>�,���f�.d�>@�_>�dZ>�1�>e����՟�_K�<�?SR"?e�>�x^��ɿ�J��f)��l�?�|@XEA?g)�%뾕V^=��>r
?h@>w�0�L��@�����>ٞ?�?�T=��W��/��ue?|�<amF�G⻘W�= k�=zQ=���8�J>we�>3��"g@�Z�ڽ27>ܸ�>|� �Zv��^���<0\>]�ӽ�ݑ�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�퉤�{���&V�}��=[��>c�>,������O��I��U��=��ƿy�$��|���=;�p \�?F�g���HU��#���ro�\�轚�h=�D�=]OQ>�Y�>��V>�Z>�eW?��k?b`�>*q>6}�����ξ6���.�����d�������裾NT�ɂ߾j�	������vʾ�i>���=��O�2o���m"��gd��F��t.?�>�+ξ߃M�"�?<{1ž�奾	R/��$����;h�4��q�x��?|@?yŇ�,X�������|��V?����i������^�=�ޠ�a��<��>A��=_����0��P���A?+G?�pѾ�t~���
?`� =���<��4?�N1?��=�.�>��D?%���s�S���>�e�>��>��?қ�>����c�,��?#S?��l<�����>2Wþ�
�X�L>A7>����v��=���>��ȼr����v<��9����=y�W?1�>�)�����k��}�k|J=�\z?��?��>�i?�+D?ʥ�<�;���JP�h���=\Z?�ah?�c>�z���mϾ�u���):?�ne?�PA>��m��&込D1�)� �{8?3�l?�n?���E{����C����4?��v?�r^�gs�����>�V�}=�>�[�><��>1�9�`k�>�>?W
#��G��ﺿ�Y4�3Þ?t�@z��?��;<	 �3��=w;?d\�>��O��>ƾ�|��˃���q=n"�>ь��,ev�����R,�r�8?٠�?W��>��������& >�-�1ȭ?�l�?�A˾�yV>��&�e�q������Q>V�>�l���7=6�����^��b���Ѿ(g=�� �>E&f>�@�;h�?�>ъ"��F��ο�g���-���d���?�>����cN��Wt�|أ��f��p$���2����>Z�>3𓽧���O�{��L;������>�/�Lz�>9�R�}����P���!P<���>�
�> �>Q���p���_��?E*���JοӬ�����g�W?�Z�?�?R  ?yJ<Yly�i�{��*!�0uF?I�s?'xZ?{���k\��7�žj?_���U`�0�4��HE�(U>c#3?AD�>y�-���|=�>��>1k>h#/�L�ĿRٶ��������?0��?�o�b��>���?
t+?�i��7���[����*�+��<A?z2>����9�!�`/=�fҒ�^�
?@~0?0y�.�\�_?+�a�J�p���-���ƽ�ۡ>��0�f\�3N�����Xe����@y����?L^�?h�?͵�� #�e6%?�>`����8Ǿ,�<���>�(�>�)N>rH_���u>����:�i	>���?�~�?Qj?���� ����U>�}?�%�>�?�n�=�\�>�j�=������-��k#>a:�=sE?�ߜ?�M??E�>�5�=��8��/��\F��ER��"���C���>��a?��L?�Fb>���X2��!�z�ͽgm1����2\@���,�)�߽545>t�=>�>f�D� 
Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?oQo���i�B>��?"������L��f?�
@u@a�^?*���8�������}���K�<����@
>��:��*}�|>!>쩼G��=Lҥ>�>4[q>��c>�Ր>=<o>2�a=����0����\���B���-�\L�j��q�����}����K�)k</ؽ_����S�J�A�Ѝ����=}�U?�R?p?�� ?+�x�d�>o���:+=%r#����=�)�>	g2?�L?v�*?��=�����d��^��>?��[Շ��>E�I>�s�>[�>�:�>\��8c�I>�[?>���>�� >�q'=�M��(=��N>Bi�>���>rx�>JĀ=��G>�ʼ�Y����7����rhӻ.$�?���Q����'7Ͼ?R7�=��/?�1�=�Ɇ�4bǿ�
��iA?3蔾ެ4��kQ���@>I=?��^?�W�=�!��F����O>�E��/[�g���e��W�5���%�U��>� .?�2>��J>4U^�wAZ�`%B�� þ�A�>rtA?TW���c���d��{��̝��3�=��E>s\�fqC����@K^�1�\�u=(Y=?T�?�{��K��y����oA�I�f>��>�u����=��>i�=hW���J��x=�em>n,4>U?g>�S�=�Z�>~����5��;�>��3>�N!>��>?��!?)m@�{p�����x�*���~>���>I߂>e�>x|M�O�=�.�>�V>��`L��
�=���]>����g8R��BS�a/V=�����V�=��i=����2��O-=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾQh�>Yx��Z�������u�i�#=���>�8H?�V��B�O��>�`v
?�?�^�Щ����ȿZ|v�d��>#�?���?&�m�RA���@�ȁ�>��?�gY?�oi>rg۾�_Z�-��>��@?�R?K�>�9�{�'�y�?�޶?���?���>�Y�?�	E?A�>q�=�p2�3v��z���Dk�>' ��2?ͅ?Ah+�菃�E������Hh���@�Fq?�=$��>�Mf�����]>�xF��?+�d�_=�@�>U�%��>����q>�>�\>�H�>��>�B�O���Ӿ���K?�r�?8��6k��̪<AV�=`��E?�3?�G:�|�Ͼ��>��[?+�?�?[?ִ�>��r������F����<�VM>��>a@�>�~_���Z>7�پ�_T����>�I�>��߼:�־Kf}�v��NV�>X�%?�;�>���=ʺ?��#?�q>�y�>�'E�3��4�G�J��>�$�>+�?P��?_K?�g��fd4�/���n����Z�`R>�{?F,?��>�鎿����fy��Rw�����S�?�)e?���d�?�e�?��;?=?��`>��x+ܾd5��z�>�N!?��u0C�us'�����?�?ah�>���� l޽���!1�V����?�oZ?��$?~���a�۲¾:��<H��8sv��?<`���>�G>Yq���l�=~>(
�=�Ho�`�1��n�<R�=৐>iQ�=��3�؅�K<,?ԃH�KӃ�B&�=��r��nD���>�;L>���X�^?�l=���{�����u���U����?̟�?sj�?Z����h��#=?A�?	 ?^!�>�F���~޾8��w@w�ψx��q�U�>R��>,_k��9������_A���ƽ��C����>!�>#
?a��>&�>�`�>���38� �6]��+W��(M�ѻ�52�<z�L񋾘�=�� 3�1,ܾ-����Ӯ>�<�! ?�&?��>0��>���>���in>3F�>���<ԩ�>2�,>Y��=��>}B>��
��KR?o�����'�ж�򲰾,3B?�qd?�0�>ci�͉������?r��?'s�?"<v>�~h��,+�yn?�=�>#��Jq
?�W:=�C�E1�<�V��N��2�����>bA׽: :��M�{lf�8j
?M/?���Y�̾X9׽!���cُ=0��?",?��)�%J��t��;Z�RG�ë,<�V�����D%��p�լ��^�����P���=�@%?�?W*��8������u���A��f>��>27�>%��>�{>�^�=���^� &1��K���P�>��v?z�>�vA?�-?�K?�"d?=��>��>Ж���>[2�=b�>��>:b>?=�)?5?^�?�3?�s�>�)����h�ݾ��?��#?�0?��? �?o;���h��:$=��<��4�=�M>0Z�����!����<�;2>\�?�h���:�3����'f>�5?q��>+v�>�?��z.��
T�<�U�>6�	?Jz�>O` ��.r��w�e,�>���?gp��	=�y.>���=Rhм�-�g��=F<��/9�=�\9��VQ���<[R�=��=��k�u���Z=�;�<�ƪ<�q�>_�?��>Bf�>�?���� ������=s�X>S>�>�Bپ�~��R����g��Wy>v�?�w�?Ċf=���=��=�]��7���������;��<s�?�J#?�HT?Ö�?T�=?�h#?W�>��TQ���_��>�ä?K�!?R6x>��1d�1����4�=v'?j�?��^��U>��E3�9����>�2�=�=�Hsu�.��,�$�)�"B������?i�?�`�b��yb�m������fE?��>=o�>��>{��o�D�7����x>9��>�W4?@*�>J�O?�2{?Q�[?>^T>��8�t+��4̙�f�1���!>@?���?��?�y?#v�>8�>��)�"ྕK�����@�ւ���W=J�Y>4��>,:�>�ة>�D�= fǽ>8��W?�咥=��b>���>ƥ�>�>�gw>��<�4U?�N?��ƾ�*
������b��=9T�?-��?��G?x�����='�!%žm_�>�X�?��?��A?�ƽ�}>*)�mb߾��} ?��>��>Н=nU'>�*�u�>%? y���.���0�H���"{?R_k?&�">C{ſ߶o�R�k�H�����<Tː�#�_��ɖ��]�W�=`ٜ��+�1x��܊U��D��R��* ��=^��
:}�[^�>�y=WW >2��= �<�t���B�<� f=��<���<#������;�Q���I��✽N}����<��e=H�����˾4�}?C;I?�+?r�C?Ѷy>�6>��3�Ǜ�>����??�V>��P�U���\�;������!��ɵؾ}w׾��c�ʟ��G>�]I��>83>�F�=~j�<��=J
s=,��=f�R��=S$�=�U�=�k�=`��=��>�S>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�??ti��d�>M���㎽�q�=J����=2>q��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>$>�4+>�x���p`�wޱ��������G��>KDQ�9�Ⱦ��=��)��џ�q����;��>�H�7I��V�k�&��=�½�T�P�U=��>jq>A��=��i�׏H>� <2� =�Փ=)���I���)齻û+.�<K�l>�k�>K��>p?-?�?S?p�Q>����5��:<}�M��>���>�L�>�_#��@X>�"�>� 5?�+?*x<?��>��=���>+C�>_9Q�b�v�m����C��=�>�?�v�??�c콐������<�3�< �=�9?�C?m��><y�>�U����9Y&���.�"����m4��+=�mr��QU�L���Im�3�㽮�=�p�>���>��>:Ty>�9>��N>��>��>�6�<|p�=ጻ���<� �����=!�����<�vż����u&�8�+�;�����;���;T�]<i��;�J�=UL�>{u>?��>�7="����T>�9��`�Q�b7�=y��+�A�P�a� t�O](�k>Q�>T>�^9>���-���>�>H�l>; +>�G�?Wp{?��>�_���ݾ;f��X�\���-�|趼�}>����8��N�[]M�̀Ǿv��>*��>#��>`3K>U�B�O9;��*>�����9�xy�>毘����"ļZ�X��ԝ��Ǚ�˒i����W+?����~�=�H�?#C?ȭ�?�[�><��aN �Ej�=�����V�=7�̾"dݾXG�ϱ7?|-?)0?z��M2�|H̾N���޷>�@I�.�O���F�0�Ȭ�<ͷ�+��>������оh$3��g�������B�Mr�L��>�O?��?W:b��W��AUO����I(���q?�|g?0�>�J?�@?&���y�xr��lv�=�n?Ƴ�?R=�?t>">�#���?��*?�,?ץ�?GRk?誐�	��>���:e�'>⋽#�뼓v|>��=�V�=�g?�9?���>��ͽ9�������(�H�:�Q3��Ć*����>]��>��c>J�r>�r.>.?>���>�%�>���=s�=���>��>�b���$X��>?fN�>�H�>dx]?�ȍ>�_>}��F;���f�lϡ�q�z�e?>s����"�s>��3>ܵT="��>�;��2��?)l9># �(h?{�����=Q��>[=�=�h�>N��>s�>#X�>h�=�?D+�=|�>��<>�оo>����#�m�A�`R���;��>�:���,��.�8	�>LM�����ؕ���i�fȂ��E=�(�<�z�?�T��p�h���(�=P�[?�٬>��4?$֍�|��2�>���>`:�>�6�������/�������?���?��c>�u�>��W?�?��1��#1�t�Y���u�A��d���`��ٍ����%q
�z�~�_?��x?[hA?^:�<{Zy>�}�?Mm%�	C��*�>;�.���:��;=g�>柱���_�c�Ҿ��þJ@�4DF>��n?���?��?�WV�m�l���&>H�:?4�1?�/t?	2?s|;?)���$?+�3>bL?=k?|.5?��.?��
?��1>�#�=2K����'=�쑽5����$ҽ�̽�;��p�/=�hy= I:ҟ<x�=�O�<��]�Ӽ�40;䡡�l��<�98=�a�=��=�k�>4�[?���>�ml>TBM?��˽ܵ.������@B?�v=?�r�^���Ӕ�nW ��W>:�}?��?O�^?uu�>��A���O��a#><��>&?>��p>I��>����w�s�=��>��>���=�t��t���C0p�*pԼ�N>(�?�V>Uk޼�K�>t�����%��B�>2�����оZ�Ӽϴ9���2���5�Ķ�>��=?gR,?�U>0�F���&�O�m��>Ո8?Jaw?�\?u��>����<���U�3��� ��>�N�� ���*��������g>'5�>�wE��ʞ��g>��
�c}�Ɏm���J�_.龠�Z=:���za=�8��־����$�=+=>�ƾ��"�n`���쩿��J?3�p= ���$b��Y��\>�ޝ>s�>-;�a�g�]�?��8���o�=b��>��B>a��}��GG��c�<Y�>+I?�Z^?ƈ?H�Ⱦφ��h~]�N����]�8�ŽI�)?�Ŧ>9��>◝>|b�|�Ⱦ*]�0/W�T�M�M��>�o�>"E-���X������3��~!���>�;?���;�#s>k�U?�K�>��@?'�;?��?�*>6.�a��_�$?Cj�?��I=7 ���!���M�_u`�ӵ�>�P??�=��3>6�?���>o
?H[5?�M?��!=*���u�D�|B�>j�>��Z���d�>6?�%x>��E?�=�?*b>�C��g;�l�=*��=�^t>�~,?�B#?��?/�>�P?->�ťv=w�>�i}?���?�o?�k=��>��>�Z!?VY�>���>߫�>uY?`�L?y<o?Gs?%@;?���GԽ~D>bb�=�.�
5���<�+�i�v�<�=��>��=�U=5C�1��<8�U��[�qR��9a�<�>rt>����x0><�žL;���A>n	��Vl��������:����=.�>n6?9<�>��#�%Ǐ=r#�>���>�%�v�'?�;?��?30�;c+b���ھ~�K����>�@?�{�=�8l�ح���v�S�r=��m?��]?f,U�ZF��ӟb?�^?��򾷔<���þ�e��a꾤UO?�
?��H��l�>�z~?oq?���>�xg�=n��
��_2b��vl��t�=x��>(n��e�q�>�?7?���>�c>�I�=��ھ 'x��'��R*?���?��?��?�)>�n���߿���@V��M~V?i��>�/��Us?�Wv��f�%������;�ƾfB���ߓ�6̧�����*1K��m�hB���O>DB?��?��x?B1]?�j��	e���f���r�#K�s� �V'���A�Z�F�K!V���x��a0����jSѾ�s��l���V�^�?z� ?�T|��b?���L��1���f>����RM�͜�=��<�V=��=\>�/鴽߯b���?���>��>-�B?1Ui���8�k�5�/�C�����=�n�>��E>5��>5��<0{v������C�Qy���ؽ��>
ni?~@?�'a?�E۽8�j~���#����<N-��8>V�=L}�>Z)�%��;�!���A�2.p�"���������n&=&l!?��>"�>�N�?���>� �8ƌ���.�?�4�2=�+�>�N`?Hn�>�=�>�+��� "�ǹ�>L�l?"��>��>����HV!���{���ʽ�"�>F�>���>}�o>}�,��\�,h�������9�Ʉ�=Ũh?������`�Uޅ>$R?߈:v�G<�z�>��v�p�!������'���>�y?�=�;>�žv$���{��<���d)?�?�:��+�,ő>?���>���>�1�? =�>A�̾��(��N?!�`?�QF?E<?"��>!]=v�ｕѻ�#$+�\h3=Ӻr>I�=>�M�=P��=.�+�c�ܟ#�gi=B��=�0�v�ʽp)=��7�����/�<��#>�)ڿqcJ��Tž ���l�[�	��#���'��љ����R����皾KZr�U;8����k�x���h��=����^�ɶ�?K)�?�{�ņ������4ۀ�X����>\m�Y��L������a����۳�rd,���[�9Fs�g�q�=�"?��g��Aҿ����$9���>�W�>4��?\2������j�zc�=�,���c� �힩���¿�J �k�2?���>�߾�(���;�>fv�>�2�>�J>�/9�w�����{'�>;z�>�%A?�Z_�G�ۿ쩬��� >��?�@=yA?��(����H�V=��>3�	?;@>�b1��>��찾�l�>~8�?��?T�L=�W�V	���e?Ti<��F��ݻ��=�]�=�=����J>zQ�> ���PA���۽��4>��>9H"����~^�fż<�f]>Heսq���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=a� ���ſ���T�i�<��.<�w���L��`�hC�e��Z J��x�	�c=O5�=��]>��>Z�p>�Ƒ>N)Q?8�l?_w�>")G>O�VՏ�9c��s������>���9����fk���M�[������
|��;��Ѿ56����=��@������#6���r�yI���0?��=M����D�R[�=������׾3��DWC��x�1H�'Tg�;�?��4?N���ſr�,���[�;9�=�s?~J#�I�
���پ���=�_ɽ��%>M��>��0>2Ӿ�G�n=V��z<?$� ?�f¾�����G�>׷�=k�=z�-?��?���b<�>B I?�F�n}{��#�>َ�>T*�>O�?*��>ߥ��et8�U�*?��N?��@�[�l�w��>����|�=·> �=����o2�.d�>�35;I���(���.��i=5�X? *�>b�,��F��a�e�+�@?=��w?�?LՁ>��h?�C?�=y���"UK��r�K�=)"c?Gg?>�5��;�;�����5?x�f?��d>4}�O��̆,�! �r�?	�k?Ϳ?Wk��y��]�����?xA?��v?�r^�vs�������V�s=�>�[�>���>��9��k�>�>?�#��G������pY4�%Þ?��@���?i�;<��@��=�;?\\�>׫O��>ƾ�z������^�q=�"�>���jev�����Q,�_�8?Ӡ�?|��>��������>���
�?F�?�4�v\�=��'��f�^�ɾ��4><K�>��W�K0=�����T�Ҿi�:>��q�[�>Vڊ>�R@E m��?�c��xb���ǿཧ�꘷�ڮb�D96?!��>�ڰ�aꤾ�%����k�j>E�P�_��ܾT��>�z>�ם��E��������B�J�,����>hɃ�i�>�z^�ǜ���z��A�߼s��>?�>�'[>����þ^Ҝ?����!Կ����-���V?�L�?Q
�?�X?��-�����C~z�i��=7N?��v?�]?��0��K�����9j?%���'a�" 6���C��U>�~3?@)�>\�,��yh=�z>_k�>,S> C.��6ſP�������VD�?��?G?龲J�>��?�*?�d��ʙ��~��O�)����G�@?�}1>`���Zm��M9�둾#I?��0?i��ְ�]�_?+�a�M�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?0�>W�?_�=y^�>K�=�����+���#>���=�=?���?��M?�H�>L��=N�8�`/�(_F��?R�����C�V�>��a?��L?O�b>T����2��!�[9ͽa�1����YB@�d;.�f/ཏk5>-�=>��>��D��Ҿ��?Hp�9�ؿj���o'��54?8��>�?����t�6���;_?[z�>�6�,���%���B�S��?�G�?8�?��׾�Q̼�>�>�I�>��Խ����N�����7>&�B?���D��Y�o�k�>���?�@�ծ?ni��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?eQo���i�B>��?"������L��f?�
@u@a�^?*��ٿƹ��$�̾�������<��>S�>(\���
�-�u�\Z�=�w�=.7.>=f�>���>��>�(y>}>Z>�����!�k���򗊿�XD��6����%����:�֒���\��g��?`����=�	��GM�{'�90-�iױ��E�=�V?�O?.El?� ?����0>N� ��7=�|���]=LSx>�0?^�M?��'?^H�=�ڞ��jc�����!��Uʅ��>:�<>���>�X�>Q߭>
��WjK>�oK>�Ӏ>��=jG=d�<,U=�)P> �>d��>;S�>D�P>,,>�c��9��XlY��N��.�i�x��?Z���4�����w��/��̻<Q�A?<d><@q��m�ݿA���tV?^]���?�3�'�$e�>��8?��@?V�	>9Ï��#�=��̼Y�%tI��K?=��$��_b�R�5dQ>�p�>U�n>p>�G7�)�>��5O�F���>�^;?[�+�:�wy�I�Q�jž	`>��>�m&�u6�����z�
�h���=��9?�?u+�s*����h�㙾�E>Pr>L�s=zU�=�`>*��,뗽 Q+���Y=vW�=��7>�?�K6>q>���>��{�����>�>|>(*R?��A?J��?5���y�n
���'>,�>�U�>hA>K�;�'�=u��>��Q>�O�S^��<��A%.���@>�[	��q��7ͽ-�=̽>�=w�L="-�tj� T���~?���)䈿��6e���lD?X+?� �=��F<��"�F ���H��F�?p�@m�?��	�ۢV�2�?�@�?#��a��=}�>׫>�ξ?�L��?��Ž7Ǣ���	�)#�eS�?��?��/�Rʋ�.l��6>�^%?�Ӿ�~�>�m�as��F4���Tu�+�#=c�>hH?$\���DN�\D?��>
?o
?	��¤�_	ɿuv�N*�>t��?�ʔ?̸m�S����?��D�>ׄ�?�lY?,di>�ھ�x[�s��>�1@?�*R?x5�>�w��>'��?�¶?���?�Um>[8�?(�d?��>����P��g��rZ���p$>�F,��>~p!>Ͼ(������r�r��q�,����=�T4=BM�>�_g�Q���#�p>���΢�臑�\��>ֆ->o��&-n>-��>���>��>V��;���#Z��㓬���7?�c�?���l�O�Ű�=��+�
�|PT>j?�2��
��u��D[?��u?3h^?�ț>,�4�PB������/�{��8��>^a?�^�>�^�k�>yt�JrI�?����P�>P�>Z����Ҿ�k�=��>?��>?�0>c�?�\$?�Lx>C�>x�I�
*���&I�Z�>���>|�?VӀ?�?_����?+�}唿�����Z��^E>�r?��?���>�揿�<��^�<����ǣ����?��e?|�U??�?�k6?��@?љt>/��K�ؾ���Ic>�M!?B� ���@�B�&���	�Wk?�?C��>(k���ĽZ���A�Cf���?�kZ?��#?��8Q`�ɾ���<�f>�,ݲ�LB;�ga�j>��>շ��'�=W3>�Y�=��l��0��Sc<���=�!�>s`�=�=4�V!��/=,?��G�zۃ���=��r�<xD���>�IL>����^?el=��{�����x��	U�� �?���?Yk�?h��?�h��$=?�?R	?l"�>�J���}޾5���Pw�
~x��w�U�>���>2�l���K���ٙ���F��a�Ž�{�}��>g��>|p(?�?��D>U��>� ��+���$�$1��;XV���)�p(:���������s��+����>Ծ���3��>�{y����>��3?��>2>���>�JE=���>���>��>��>m�>z�>��>�j�<(��;�hO?$���G/�"���{���"<?sg?U�?�f�%���f�P� ?�l�?��?�,>}�l�M�&�HI�>���>�y�q		?&�=\�D;����C�Ⱦ���6Hf�ɾ3�/��>�����a5�8��R��>K
?�z?��<^Cƾc�1��R쾐J=.r�?�w?4y8�;b��u����h��ka�8N�=�3\���~�(�%�����q��0����A���9��Fн��=?���?y��b�|۾�bh���5�6_�>���>�>���>A��>@_�����#���<��)��=��/?d!�>_$D?�c8?��O?�N?�.�>f�>���^��>oW=���>+�>�F4?��,?�_1?pO?�],?̔x>�������aԾ�,?lQ?`V?H��>�>����ڣ�:\<�=�o�r�����=������/�d��I�=T>��?�{�X�^��
3�-Ģ>(?n �>�?둾+���s�V��*>W/?���=��E�L������]>=ހ?���0 =x�v>��=x�>�k�<�Y�>wz_�"k >*���p�����L�GHZ>(`�>�ݪ�B��=��=�5����s�>��?��>FN�>4��� ����B�=u�X>S>�$>>پ�|���#����g�Oy>�v�?�w�?f=,�=��=�s��)R�����l񽾣�<r�?�G#?{XT?��?
�=?Jf#?��>)�[L��L]������?�!?�Ŋ>��"�F��]��ّ@��$?d�0?7�M��g��s0����|>��>ʩO��~v�������H�4;��7��k&<7��?�J�?�?�DhS�J�2���~��(�-?�,?�R�>�*�>˒��{ 羪i���30=A	?��,?�>t�S?�bt?� T?��W>:G;�~��ԙ�����<.>%>�4?�u?7�?�wy?�_�>+�>�0B��S����� ��/꽢{��%��<��X>_��>t��>xڞ>W�=*���5JŽE�d�K��=@\�>���>e�>`��>�,w>�n;_�Q?ޗ?;K�6��F7���d��@�9�?�$�?b�?�i�=f9ྪ���
�<F�>�v�?܃�?��B?\����=�M�7�о�c��+?�)�>��>��=u=AY����>3��>�GD��� ��/1�>��;�;�>�Xv?(�x>*�ſ�oq�0�o�g���-M<Mܒ�ed�ٓ��D�Y�N'�=Jt������,���LZ�����hq���r��O�����z��v�>1߃=x�=
��=�<\�ʼ=ұ<�bH=�`�<��=�Dp��Չ<�6�߮����|q���p<��K=a[�fo���o?�AR?�08?�E?٬�>X�^>,�����R>�ڼ��?G�>�����DH��9��hS^��Ҿ���C�A�:��4��=ga��l�=�/>ps�=��<�\!>i��=���=侏=�Z�=��>g	�=���=D%�=�s%>��;>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>מ7>�)>i�R��}1�F\���b��-Z��!?$%;��`̾��>�)�=�"߾ZsƾN/=�m6>��a=mm��@\����=A|{�Ɋ;={k=ŉ> D>�>�=����m�=8J='�=��O>������7�;�,�@q4=���=��b>�4&>k{�>��
?�*?�f?���>O��S�����ž�j�>N�C>b�>�L>
f>{�Y>��?��*?��L?���>Ի���>���>]�Q�E<�����{���W����^�?G˟?�>�)4����	�C�.��ڐ=~b/?�1?��?Oxx>���p�鿸��K������kk�==P>�����X��7ڔ��׽�9���z=#��>���>e��>ZQ�>���>�%W>>N�=n��=᷷=� =*�<b�V��h�=1�<>J`�<�����d���<<`L��(����3<zn�;�U>���=�^�=A��>jG>�:�>d��=q��h�0>Д���L��=�����A���c��R}�.�-��-7��a>>��W>�S���7����?�%\>�1C>[��?%�u?ka!>����ԾW�����e�TBS��ܩ=��>��8��:��z_��iL���о��>��>��>J�r>�84��P�	��=�姾u�0�X��>����R~�n���2K�?���!O��g+l�j�B��]2?�ފ���=��?�ic?�i�?�}�>ו��a�ʾJ> 徒%�;f�����ؾ8\��v3?J�?0_�>�z���X$��̾>��B$�>HI�>P��Ε���0���$�d
��'�>�ê�SyоD3�����;돿}�B�5Ns��:�>�iO?��?Ha��l��U�O�	��l��j�?E�g?�>W?j?	ՠ����c��DK�=��n?��?��?�#>���=j���,�>��?��?;��?�.z?=W*��,�>w�a<��w>م�	�<��=u��=a��=��?	�?�J�>f�w��q��nD徇���q���.=�}'<w'I>�j�>pޑ>3">32=Μ	>�7S>"}>Y��>�/e>xr�>���>�ɣ��
2���C?%]�=�V �!�3?��?>���=�!X<'�=/���_��;�I���>}��<�ʼ�  >�kI>�r>֯�>����yg�?kC>�����??6b侻�@>k8>���>?���-^�>�t}��]>��>s��>k�A>n�m>nt><�ҾY^>AS�s�!�D�B��[R��Ѿ��{>+��h$��	��b����J��K���D�Pj��:���=��`�<�?�)����k���)�<,����?���>&�5?u$���뉽(>���>(�>�F��ĕ��ɍ�k�ྻ�?c��?5Dc>�>��W?Ț?��1��3�sZ�O�u��"A��e�7�`�ߍ�ٛ����
�������_?��x?ZwA?��<�@z>(��?��%��ߏ��!�>� /��*;�b�<=�9�>S*����`�&�Ӿ�þp9�>UF>��o?�%�?�W?�VV�^���z&>��>?Zn<?��p?#2?oA?x31�b�?��q>��?!�?E'?Y?P?�>�5>��<1=
pd��z�����jH���e��
�<�#=�B2�{�=�St=�uл��;��<��Ự�r��q4=�BX=���=�2�=�j�>�]?y&�>ot>�	=?������0��a��Ś5?��;,\a��n�����	���?H>N�n?2w�?W3d?X�p>h�;�>	>�~>���>�:>=
y>C��>��N,a�Uy9=%�
>%>A��=ɑ@��3}���
��H���X>=OE[>���>"n�>+$�ؕ>� 1�������N>&�w�;ަ�:RξVn7�F�e�q�d� >��B??*"?�>����J�X���W��k�>JqW?�1\?��r?1$w>᳈�Mi)��=���;G�?��>�H:�H���}�����^�S��œ>��>�Q�����Orf>��}��p�@P����6�=&�&�$<��0|���a���>>*�Ծ^$��L��r���MM?�y=�귾��P��Ŭ�n?>�g�>��>�%��km����;�RK���>�=W��>�jV>j���޾.L�B�	����>((B?�`?S��?�:s�u	o��|<��+��F>���z�Nt?��>��?�m;>H-�=���N���`���G��p�>�{�>����G��&��p��]*��p�>�	?M�#>��?�$V?��?��d?�P*?���>|B�>]W�"*����%?i#�?襁=���w�T�:�9��(H���>U�+?�;��M�>�?��?�v'?+�O?Z�?�e�=�� ���?����>aw�>��W�
��W�`>��I?��>�rV?�x�?+�I>�Q5�hѤ����#4�=��)>�2?i�"?�?8��>��?谁���?�7?���?	��?���?�-���>�K ?c$V?��>��>͎�>ZJ6??O?Qv~?�*o?�^ ?�rͼ>��$Խ���L}�b�������E����=\�M<��Q=}�=U��<,��<
`����h��7˽���<kxӽ�a�>e�s>���J�0>f�ľIM��,�@>�e��OR���ъ���:��=���>t�?ح�>CW#�XȒ=���>|D�>%��H1(?#�??M�;�b���ھԫK���>�B?a��=T�l�ၔ�|�u���g=��m?�^?��W�D!���E\?�i?����m?�6
�������;���0?O�?����/�>��^?��m?�?�)X�>Wh��?��i�\�Si��J*�=m+�>���Yg��Ğ>��1?���>�6*>ڣ>�����r����7?�ܔ?HԱ?	-�?pp1>:u[��ڿ~m�g���kd`?���>U�����'?�L��ݾ�nJ��1�۾=Ԯ�H��������þ�)�u���佣>�8?�Cn?K�p?��d?����N�c��U�G�z�AV��M뾥��eYJ�uD?�?�B�F�p�Z��D����;����=�ks��U�>q�?��0?��z�*� ?����3��(����D>#��4����\=�@���*��a]F=�H��u7�G�|��=?F&�>\F�>s+F?W�ְ8��H$��2��~����z>��>{]>���>)���\�v�O�ӽ�NžϾp�x�.���>Cj?�f/?�R?�ɽ��D�ş��_X�#� =l���Ml�=U�={#}>��<��75<1��h�G��r����d阾����#>��I?��.>��>���?�N?cJQ���[�o/���U�)�z����>�@?^��>:s�>�=3?/����>l�l?���>}	�>d����_!���{���ʽD2�>0ҭ>��>��o>��,��&\��j������ 9�G�=�h?v}��o�`�yօ>�R?�l�:U�H<b~�>[�v�%�!�(���'���>�}?o�=ò;>�lž�#��{��:��3)?jh?Z�����*�H�>�h?���>};�>Є?<�>jFľ$<�a?�_?t(K?zm@?�q�>=�=�ײ�\|½�R'���8=�>ĠY>Ua=c��=r_	���b�p?'��!?=*�=�7	�vlýOY�;�հ��0�<T�<p�6>��ֿ��A�^���g~���wf�r쓾�ս�0��ph�����'��g%��O�Q��O�������\����2����?V��?]M���ڧ�N���e���ڶ���?�2��-[����w�4�O�1��I��}2����E|��ݑ�ƃ�K�'?�����ǿ񰡿�:ܾ#! ?�A ?3�y?��>�"���8�˭ >}B�<(-����뾭����ο_�����^?���>��F/��W��>ť�>�X>�Hq>����螾+1�<��?(�-?��>̎r�+�ɿ]������<���?+�@4�A?B'�$��'�K=%^�>��?��@>�/��c��ⰾ���>�p�??�zI=rTV����qe?U�9<��D����<��=�g�=�h=SU�X�K>�ڒ>��`B@�/�ؽBr6>�J�>]3 �r��O�_����<��b>��˽sݕ�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=� �6�ſ��=��1���L���t���ʈ��P`�������d0��+�v�\;m�d��h*>��e>>?>�Z>NV??n$X?�>�C>����n�Z����|�=q�H��!���~�uI�n�ܾ�K����U������Ӿ*Y��G�>���=��C�����K�!?x�4:�s�@?��A=,�Ӿ�m�a���C%��r]��vѽ��P�!]�F��r��8�?��>?�
��+�H�n����ͷڼ:�?�(k��������P;�o��=prR>q�>+�g۾pQ{�N����hK?�m7?���l��;�b>��f<]�e>A�n?U"�>ȑ����>mX?Ԁ�> ���l��=Ł�>'%�>�4?$+?9���ͅd�J�P?�4?j��ۇ��[�>��ʾ��о�C�>���=����{��.�>��~=DUƾ�v
=A�3<`V��4c?�7�>r H��F��K\���;D�>3�?R�,?qd�=ͮH?�oh?f�=��G��7�|�����>5�v?�j�?O��=Y��ާ׾bp���A?O�Q?��>+��������p��:��AM$?���?YJ�>�����@�2_�����)�M?��v?�r^�os�������V�e=�>\�>(��>��9�jk�>
�>?#��G������lY4�'Þ?|�@|��?�;<I �ޛ�=�;?d\�>0�O��>ƾsz������ْq=�"�>����yev�����Q,�R�8?Š�?v��> ��������=��ԾMɫ?�R�?99��zi�<{��(�������;�8&>��T�� ^�GNо��{�����j�����6>Qb>��@���t�>�Ү���,�ѿ�f�@ƾo_[��i+?�f�>>��lB�%hS�����l�]���V־��>��>�����쑾�{��{;��
��\�>p��ke�><�S�w���џ��=< �>���>�Ȇ>{Ů��轾���?����Lο��������hX?�F�?�l�?c�?=zI<_�v���{�P�$��F?]s?�IZ?{���\��p5�(�j?=_��eU`���4�WHE��U>�"3?=C�>7�-���|=>���>�g>�#/�`�Ŀdٶ�����]��?���?�o꾿��>y��?�s+?�i��7��8[����*��b,��<A?�2>[���L�!�0=�2Ғ���
?;~0?�z�i.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?9%�>��?�q�=�_�>�j�=���V-�i#>�+�=��>��?o�M? L�>�[�=��8��/�[F��FR��"���C���>��a?��L?�Mb>����2��!��ͽ�g1�z?�&W@���,�Q�߽�%5>��=>�>��D��Ӿ��?jp�3�ؿ�i��[p'��54?1��>�?2����t����;_?3z�>�6�,���%��eB�L��?�G�?2�?O�׾DO̼>*�>�I�>��Խ>���}�����7>�B?#��D��=�o���>���? �@�ծ?\i��	?���P��Ua~����7�e��=��7?�0�!�z>���>��=�nv�޻��W�s����>�B�?�{�?��>"�l?��o�Q�B�t�1=8M�>͜k?�s?�Po���j�B>��?"������L��f?�
@u@a�^?)B_ڿ����&�о��G�ֽ$��<�#>�ٺ�=�&\>�4����f��[���U�="">W��>�qQ>�q�=�q�<�w���'"����'���isa�����C
���j��- �4>@��O�oþ���\�۽���^>��q��w�"ż!*�=��@?&�T?�n?!+�>?�+�lh@>���r����|O��ܕ<:_]>��?��1?E�1?--2=/1���@c���3��P��ar�>G+>�1�>��>�d�>�s<��]>��=�!�>�Y>�f�="��=!��=na>��>�x?��>�>�>���栿��Y��^ݾ0�1�=j�?8� KD����^��Os���k>ݴ ?�"�:���nؿ�n��ER?y���5��渽���>��+?�E?h&�;������_�+R�>����O����<�Ų�Ľ�w�w�f>�5�>��t>8�>ңd�;�R�o�
�L��O*�F\*?C7����ݾ����[{����&�=m�x>�e���<��$��>ό��"����=�G?H._>�`G�w���B�ľ�
~>XH>T@��N镽6;�>����Um���x�-�ȼ��(>�(�>j
?�Y)>+�=��>����M!�p��>�-j>��>*F?�?������1z�/�"��w>�B�>\?�>��6>e`���<�� ?��>�Po<�������m��߳<>�����[��O��t�F=�O��P.�=H;-=��
�GL^�X_y=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾOh�>|x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?roi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?�r>�ȟ?	�E?��>G�0�.2g�U�Կ�����Z�>%D&��F�>�N>tp���f�Kn���0��8��\�EJ�=aj�=��>����i�(>;�<uk����;���>���>��q�����e?��?�)?�:�>���	�����۾��6?'ϙ?XL���o��ג=��7���pk�=��?۠S>�����>�?��?�gx?tʈ>k�K��Ӌ�ջ���jk���P�;�9>P�?IQ�>ݱy���t>��9�]��iqL<�_Y>FN>�־S���Ly�=8Z�>��$?Q�>im >(�?�(?:T�>dz�>�@I�S���dD[�{O�>���>Q ?~��?Ɏ?��ƾ�H�L��������b���A>j_q?��?�u�>�[�������<������T���|?Y�z?�Z
���?4�?~�7?�)?%�>���
8��t����+>ؗ!?̈��7B�Do&����d�?�S?|�>`���N�ڽ�鼝@��m����?f�[?R?%?���2�a��Nľ��<��:y�,�;�S��X>��>�[�����=:�>�|�=�m�=�6�/�T<sֺ=���>���==�6�<����=,?��G�Oك��=}�r��vD���>pOL>1���^?�k=���{�o��
x��DU�{ �?]��?�k�? ��Ɲh�"=?g�?{?@#�>�G��U}޾֗��Qw��ux��w���>~��>f�l���쏤�6���jF���Žt��M�>�� ?e�%?��>�`4>���>�P��Q0J�p��_f �; T�@a�j2��&������oǾTq���?��_ξ�Ʀ�i��>�q��|o�>6?�&>��1>d�>��1�%�>"`�>+BU> ��>�7�>y_�=�(>��=�qy��KR?`����'���辀���L3B?�qd?l1�>�i�*��������?���?<s�?"=v>�~h��,+��n?�>�>9��,q
?�V:=_3��8�<�U�����2����X��>�D׽� :��M��mf�dj
?w/?�����̾�;׽������=�օ?501?�.�R�V��u�ʗ`��3N�pDo�Z$�M+���'�Փx��m��󨋿����;#�x7�=�'?
U�?�c�M���w����z�0@X�ق_>) ?���>���>�{�>���J%=���T��/�Y霾,��>�zc?�^�>��*?�F?�O?��I?ZR�>n(�>��]�{��>�c>Ĳ�>W��>e<?m?�� ?={?s)1?�˱>��B=r���Z� �?-�(?��$?�U�>�S�>�E���L��Ă���jJ=UE�J�s��g@=X�(��	��� ��Ჽz�j>^�?"���:��x����w>u6?CE�>�6�>͔���X��R(�<UU�>�
?�u�>7�����i�7	����>�׃?���Ť=�,>[/�=ʸ���Ԏ��R�=Ъ����=Og��(�:�Zg<ɣ�=���=�_����E;�H;�p�9s��<u�>5�?���>�C�>�@��+� �\��.f�=�Y><S>~>�Eپ�}���$��p�g��]y>�w�?�z�?��f=��=ۖ�=}���U�����7������<�?=J#?XT?]��?~�=?bj#?˵>+�gM���^�����®?�?`��>���d^
�"����-�0v�>gZ�>&�I��8����t����>���=Q�?�W����ڦ�Z�Q�pO�|d�Kf*���??��?�0�_2"�{��������i��ZS?Q��>?�>��?<�
��IX�����>���>�@?�&�>�J?�m?�J?��;>�_5�s�������������S>q�C?`!z?�D�?M~?���>�w>6��BK־���h�
�95�[����&=TQ>���>���>�ڬ>��=�H��og�*��Ԝ=~WH>C(�>	��>1��>;�>E�#<`�Q?��?,�־B��t���[���L�<Ќ�?���?��>?۸�=���
�h��O�\?�>��? �?��:?0�	�	�>��;�>�v﮾O��>6��>Kn�>��J>�Y!>\ϯ��̭>���>5����8��K8����=<8? |k?���>ǶϿT�����x��A%��߀��E�-�C=�����q����������r��аr����]庾޻���h\�#3C���>]|�=E�'>/�=y��=���=xX�=��|/��{�����M��<K��;QQ>F$�ѳw<�
>��^=xMȽ7˾\ }?�ZI?��+?�C?��x>�(>F�4�r��>�9��|�?LT>n]Q������|:�W���J��b�ؾaؾ�+d�H�����>8�F�J\>�	4>���=f��<�'�=��j=���=*���=0:�=�f�=� �=���=v> O>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>~7>�
>�Ug���1�0d�o���s��F�*?(9A�l�־�x6>b�ڻ�׾�=��9�`=K��=�e������q��M�=m�����p==�<֫�>��L>�=�h��>�D{��{�= /,>h!��s��-T����==���<3/{>�sY>ws�>ѝ?��(?�}U?P�v>jE^��Sx���e�I'Z>Yu\>5��>�>��=8��>n8?�T?�N?9ǿ>J���q�?u�>��d�N����:���|��=��?��?�s�>w텽:,p��A;��,I���f�@?�U?�?w�>�l�ӨϿ655�,w+��z��+��^��圾�d��'u~��ݽUe&��M����>2K`>�N�>�J�>ʠ�=l&5=���> '>�e�=��>�G�=�{��G����q<d�)���ݽ��}f0�V�9>��f���<��O����<��<�:>���=Q�>(
.>]��>�L�=XP��$�'>�ޥ��L��!�=�#��A�@�~�b�!vx�,'� �/��Y>i ,>��K��xY�>�f>��X>��?��y?':'>%�&�r�޾x.���^/���4�Q_)=�>�����6�7�X��L��[Ⱦc�>���>7��>#�(>��A� �6�� =d����.*�i��>�Yپ�5�HGE���]�A���y����w�E��F�?x���r�c=��?$g?݁�?�?����X�b�=�Ρ����>3`Ⱦd��i���6@?�#6?Xo�>�<��V!�F̾A��ݷ>&@I�c�O�W��0��W��ʷ�*��>����о{%3��f�������B��Er����>�O?b�?�3b�wX��bVO���&+��q?�}g?H �>K?�??G)��}�@v���o�=��n?���?:=�?.
>��>����ED	?;?_�?���?
?g?�"&�r�>�+�=��>��/=L��=��:>1�2>�~=3J?X??y
�>P(�m���޾�+�*gj��mc=R�y�Y��>���>D�>i�7>�b>�Y<��>D��>t'
>F�w>�Q�> ��>i��w%���)?Q�>�>�B5?K�*>w^5��vȽ�󐾛 {��)~��������=�4�b�Z��,���>�p7�=tj?Mbҿl��?�!�>v0���-?GJ��<|�r��>�є>�$�<p��>T(�=�ql>>x���"�>t�>��h>��>DӾac>���m!��C���R�&�Ѿծz>���� ^&���U_���}I�4j��k^�	j�+���D=�W{�<=<�?eW���k���)�����k�?�j�>`6?���������|>���>͕�>�G��Ћ��"ō�)e���?���?V:c>�>2�W?q�?�1�3�AuZ���u�h(A�Ye��`�_፿����^�
�`��y�_?�x?xA?XL�<�:z>���?��%�ӏ�)�>�/�g';�/B<=-�>�)���`�s�Ӿ��þ�6�cFF>ѕo?_%�?gY?KPV�.E;�U>9$??!�7?��q?L4?�=?,�ܽ��?���>v�?>�?�*$?$�4?�Q?A�
>\��=�#4=ɏo=1,�������i��Oڽ#�A�D���qM=��÷�\��4Q�=�(���f�WM��&<�<o�U<E����Ee=D&�=�6>K�>�]?���>t8�>�8?H�ca7��r��'A/?�{&=��`#��伟�T��BD>X�k?���?ͤZ?�hi>��A��0B�?�>N��>�$>��[>�y�>�����E��^�=�`>?>\��=c4>�]��n	�������<@�>�x�>He�>�����>����IȘ����>�@-����JN��:���?�D�|�D��>�tI?Bl?��K=���c.���d�2?��L?(c?�l?�lG>�Q���#�U�r�P}E�r�>������ک��3��Li"���=3&�>����VھR�=R�'���3���<5��{�l��=��6�=�3��oԾ�Wѽ�6>�>����Id��5��4x��<�O?���=�ȥ�X6d�����=���>[�>��G��i�*�=���ľ��l=`��>pE>sWh=�ʾaW>���;w{>�K:?�h?��?�`j�W�W���>�o!��a��U���hc?x��>Pb�>��=��;Z�׾���|�f��!5����>щ?�<$�k��8�����= ��u�>IJ?,z>c�> �A?��>,mA?��'?Ӗ?�&�>�]�=
d��<�'?�̈́?�h=v(�իK���8���G����>�z-?�iG���>|�?��?��?��K?�N?0h>���^�;���>��>�'Z������d>K�I?3c�>�X?$�?#E>2�*��N��5A���̴=��*>J�3?l�&?�r?��>b<�>۳��Q�{=\��>'�b?ac�?�o?�K�==�?�2>`}�>p��=��>��>:?��N?�s?WIK?~�>��<yɮ��嶽�n�%OJ�\r�;mU<$t=����X{�p���5�<��;T����1��f-���G�>e��tg�;Q��>X�t>�����2>��¾�@�?>�+μ�͛�����7�H�=��>�]?���>�$���=)	�>��>���'?}�?��?�_>;�b��r۾�3N����>��@?v��=}dl�h���Cu���`=R�m?�m]?IwY����5�b?/�]?h�=�B�þ,�b���龝�O?��
?A�G���>��~?.�q?��>^�e�:n�>���Cb��j��ж=-r�>X�
�d�@?�>.�7?;N�>�b>�'�=Yu۾��w�cq���?Z�?��?w��?
**>8�n��3�7���̑���]?���>�����e"?�[��^�оڻ��0`�����^=��I-�����uv��1%�X����ؽ�I�=KI?�r?��q?<�_?]2����c��^�g����U��R�E����E��@E��C�o�n� W�J9������CO=�
���W����?362?�W�����>�ȓ���뾞�����>4?w�F���;E��<��=(|�=�䐾�ɾ��<���?o�>�a?-?��X�zZ������.��߾#IU>;.}>W��>�?�41����L�+����a�mi�=�n>ڭ[?�O?"v?������*��
����h���ͪ��~j>W�>�m�>f�j�m�4���*�5<��p�����!�1H�=�04?��>˞>f۔?��>q�h����2s�o�6��	<�c�>E3a?q��>V�>W���w"� ��>m{?��>�K�>�a����#�J<��I�t>+ B?�K,=�S�>��
?�	|=޲_�汍�ˌ��,u��+;c�?D��)���w�>1FT?F	���*;��>�㷽��)�72��@i�=���}E?>٬e>�Ͼ�]�� �V�fѿ�%*?I�?"����*�ͻ>�$?�%�>���>�@�?��>���dH;O�?��\?��I?�&??2��>��B=99��Ƚ~)��Q*=�\�>{�Z>3�z=���=$���R_���#�ϧF=���=�hü򋮽ڂ<%)Ƽ�2<<��<�3>|K��^c��7��G�Z��xu�خ�A;<�!�������eɾ&����m4��ż0Nݼg�\�ނ������NL��}�?VB�?P�̾�(ľ>#���i��dp��c�>�z�����x����Q�B�v�+�̾,ֵ�,	���4��[b�vT�K�'?�����ǿ񰡿�:ܾ.! ?�A ?3�y?��2�"���8�� >�C�<�,����뾬����οG�����^?���>��t/��n��>ꥂ>	�X>�Hq>����螾41�<��?4�-?	��>ߎr�2�ɿc���N¤<���?0�@3�A?�3'���AR=}x�>��
?�?>Y�3�r���~��{��>�$�?���?��D=��V�,�Ze?�b<�)F��x�g��=j��=��+=���-�G>�"�>2�"��V?��_�Q+2>C�>91�,a�5X`�5��<; X>D�ܽϓ��ʇ?Hj�)`m�t .�{�d���=0KY?�c�>X(�>9�?ŁY��ѿ����|?z@���?E�3?�eX���d>UԾ,48?̃??��>�����"��Y|���z>�=��5�W�񾏦�=���>�_�>�t?�����7a�:$�<蛑��|��}ο�%������;K��<�<�(S��/ɽ耼4�����M�T��;���=�U>�6>�!R>JY>a�[>g`?kr?O��>T��=e4p�����j��3o%=�����5�ȥ��%�����@�߾���P;��x�϶��i��0q?�`\x=�T��ڐ�D�"�0�`��A�0/?$>�FȾ5fN��<�þv^��kl�������Y̾2 1�ŋl�'ڟ?�B?�兿m�V������
�钠�q�U?U��:��qC����=�
����=>�>溮=ٱ߾�2�R�!�@?��&?���:q��#ƀ>�S<>e�=���>v��>��Ȥ�>/�6?5!��z�%���I>@�<pO�>L�?*��=pN��v�*�_^?�f?�W��^y��s�W>��y2�G���=vL=���%�NXy>�ɴ���,�5��WG��=�e?�e�>�6���+��<+��Z> ����t?2�?ծ�>8�w?�vJ?erl=&�^&����
ie>��~?�Q;?ھ>��ʒо>�}�oF?]m�?ᕯ>Fս�����i��o��̃�>�q?�3?5U�=m�v� �R���Ӿ�9?��v?{r^�ps�������V�
>�>�[�>���>��9��k�>7�>?�
#�tG��캿�4Y4��?w�@���?Y�;<  ����=t;?t\�>��O�%>ƾ?y��������q='"�>񌧾2ev�����P,�:�8?���?`��>���������=/���fp�?y�?ސ���CS<�����k�Q���
��<�S�=�9�&r ����7��Vƾ�/����x�&��>�@l��k:�>��:��+�0�οhy���о<o�1�?V�>&v���	��a�k���u���G�2�G�����F�>��>M�]��Ԫ�6�a���F�6�7=;��>�>&�~�q>�}����RS���^|���>��?�@�>-��=K˩����?o3���Ϳ킚��澩�j?0h�?�Pg?g�L?h�J> �Ⱦ��F�6�w���U?��?&#�?Eʨ=mtv�@ݑ<$�j?_��lU`���4�HE�VU>�"3? B�>7�-���|=�>��>
g>�#/�J�Ŀuٶ�����R��?���?�o꾤��>q��?�s+?Mi�8���[����*��%+�<A?�2>����m�!�0=��Ғ�ͼ
?�}0?&|�:.�K�_?t�a���p�g�-�j�ƽݡ>ز0��r\��5�����i\e�f���Sy�2�?�^�?
�?'����"�05%?��>#���!5Ǿ@d�<Vw�>�$�>�$N>m_���u>\���:��]	>c��?�~�?7l?�������V>0�}?5M�>��l?�G>�(?�C5>�ˑ�w�Ľ��=Φ=]"B��G?l�O?D��>�5^�Wr�$7�D�8�p\N�$�̾Mm>��~>ɔh?�{d?�h>~������=5������4�����u{[��]6�(��X�=��c>��'>Ь������?p�*�ؿ�i���o'�~54?���>-�?�����t�����;_?:z�>7��+���%��B�^��?�G�?=�?k�׾�U̼n>C�>�I�>��Խ'���8�����7>=�B?��D��n�o���>���?�@�ծ?^i�>��>���%�l�t�r�N��v������=��&?Q� ���Y>X��>�v��P�}�樿��q���>��?b{�?���>mtk?��g��$D���W=���>,u`?��?���=-�ʾ�3>8��>�f�BZ��](ľ|7q?yb
@H@��S?�y��cT�������O����x�$l�=Dl>�bT>�p���=� >�G�=��@;8 H>��>�ۅ>��l>�>I>N+�=T`��Mp"��➿{����[D�qK��E��:�l��#��`q��2+��ֺ�g"���Q��Ҥ������ian�d|M�eg̼	r�=R�T?Q�Q?�p?}H?q�c���>5>��� =
_#�?E�=��>�1?RxL?��)?��= �����c�T���?���;��cj�>F�G>a��>�\�>���>�;�G>��A>3��>���=�3;=�q�:�"=ӰO>��>`�>~��>:7>aT> ��@4��Ni���u����c΢?J�����I�)8���\��M�����=�-?]�>�Α���ϿႭ�-eH?�������6,���>�0?S�W?�U>�����P�~>W*��Lj���>O���^8i���(���O>?̣=�}�=v�A�LNH�Y���� پL��>��.?6�;�K�<��w���>�F�C�o��>2��>���=�d
�1����;g�9��.�V>hZ?�. ?y;½�	�SC��!�¾v>V6�> ^�>�;>�y�=����ro⽾��!����X��|>��?l.>9�=�>Ѯ��e�I�P�>T�?>9�*>�>?י%?Q��c��hރ�-�s�s>���>9ڂ>ڐ>�cK��u�=.��>O�d>՟����������B��4W>�}����_��&q�D�n=(���=a�=���=\�`�>��&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾQh�>qx��Z�������u�f�#=M��>�8H?�V����O�a>��v
?�?�^�੤���ȿ4|v����>W�?���?e�m��A���@����>:��?�gY?voi>�g۾;`Z����>ӻ@?�R?
�>�9�|�'���?�޶?֯�?�SR>B�?j?zG�>b{���&)��������t�=�NV�"�>�R>bӮ��J�䖓�����DNn��4�,�>�0=}��>&������Ϛ�=�U��䤾��U���>|�I>�">���>lM�>�z�>�i�>8��<$��7�e�Jم���K?���?-���2n��N�<[��=)�^��&?�I4?1k[�}�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��G��<��K>*4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��_S��GB�>�e!?���>�Ү=�?�6?Y�n>@�>�u�&���.�\��?�(�>0��>�=Q?tI,?Ud���D��C�����Z�E�3>��?�r?���>�6��퀟�Li�=B�����K��]�?fބ?�3��&?���??'��>�>T�Ź��{J�=�9�>��?|S�� @��T#�T��r�	?3�?���>o��+f۽�߼���~���u?63[?�g%?g��&fb�z�ʾt��<����6���<CD����>P�>-�y�{��=��>ㇾ=�U`��N1��t<怾=�я>&�=,I=��D��.=,?>�G�oۃ���=[�r�2xD���>�IL>���k�^?�l=��{�����x��TU�� �?���?Nk�?���N�h��$=?�?a	?�"�>�J��~޾L��MQw�@~x�w���>���>C�l�	�N���˙���F����Žw�;����>�`�>m|?�?��>��>�砾J�!�A�󾢚�V�e��#����r%�ܭ�iɈ��a��*���Ѿꃈ��8x>�t�s��>kC?Z�N>�n�>_��>n'=L��>��,>pDZ>���>P(1>Lu�=�s =�c佅�A�MR?h���Q�'��辄����AB?�bd?���>(Di�ϐ��%��Y�?�}�?g�?�#v>xzh��+��v?�-�>�*��mb
?;�;=�|�p`�<yb��z���퇽�g��a�>d�׽:��M�Vf��U
?2?$S���̾i)׽�U���=�Q�?A?����U���R��Q7�LJ@���=��g��c�~t��FK�ΐ��m�F|����-����=Ѭ?��?(���Y	�l$�VI�;[���>"-�>R�C>��>]��>A�J�T�b)v�o�-���a�"6?�?�?+#�>��B?��<?F�U?�uT?���>o\�>�
��P��>�Ͻ��>���>I^*?H?�?��>f�?$�>���MV����ݾN�?��?�n?���>���>�3t����t��=� �������K�<+�>�]=����zU	���=\�2>�<#?�`���=�� ���{>�UI?���>ߑ�>>~����X����=O_�>�j?Ryl>�u��p��,��e ?�u?�@(���к�� >��>�@�
p�<�G�=ͦ��b�=@7��e����<�i�=y5�=*�����L��2��f6����<�v�>�? ��>�?�>3>��0� �P��4~�=oY>�S>(>@پ }��6%��L�g�[y>�v�?�z�?S�f=|�=��=����X���������R�<��?�I#?�WT?U��?��=?Ni#?��>t(��K��q\���	��֬?}:?�e�>P���@վ������@��[?-^�>��b�����;!�� ���V��;>�X&�Ms��M��E%M�Q�y���J���S��?0�?�"=��5��V�3��Ua��N�6?��>/��>�n�>��7�/Zq�?�'�*$>���>�W?��>��M?]�{?�_^?��r>��+��Ī��<� >��@?�'|?�|�?��o?�9�>���=��)�=JѾ����8����4{��=�]>��>v+�>�K�>yҚ=�13���н�V{�_Y�=]C{>:��>�ǚ>/��>�?x>�(<��L?'A?i�Ⱦ'��ʈ�0��N �/˃?��??O�*>f辒�:��'����>��?^�?��:?[B�K8>{7<S�վ��Oи>�o�>#L�>
p�=e�,=�VX>�]�>���>��нm�	�΅�E�Լ܋"? �W?�gF=�����p��hž������ �UK�;�\<�O<K���=j�=�0ľ�Rd���?��A���u�D�U��/��k��Ɛ��?��X=_i>ɒ�=<�����Ul=궆=m=z�=C5���9j��	>���=�r�:轛=�[�<Y�9�7+�p疾G`?	1X?~X?��A?���>�T<]ŝ�P0�>𧞾�|,?��>C���f�;����0þGo��?ھ����nh�@�w�4DM>M<'��O�=[�>�Y�=w�U��_>�#>��������<��
>�Q=��.=�4�=~�>0��<�yu?:7���Ν���o��"���Z?e��>AAҽ�\��9D�?�o�H��С��t �u�?���?�o�?� ?OW����>�ᾲsV���<O�۽P��>�]>�'���>�>u�>�(�Ÿ��>��T|�?�?�?�P?���޴�O(>��)>-z�=y<O��+��yF�p�G�b�X���?�7�P3˾���>��=�A� ̸��+R=�f7>۴s=�+�a��=�E����A=�9x=l�>��C>Xn�=�t�����=��S=>�=� a>�Ib;��)�
q���=pH�=pP>��>���>aV?��/?yXa?��>�n���Ծ���g�>�=o��>���=@�=>�ߧ>�m0?W;?�ZE?8'�>��=&��>Y�>s�1�t�w���޾����
�;��?H��?c�>��=\�-��c� oA�3����k?I�2?��?�"�>ݙ�� ��&��,.��w��B�:3�<=$�m�XZ����k#��]�x�=���>=
�>���>6�u>��9>h�N>7�>a'>�'�<�2�=%�I��}�<�t1�!ڊ="������<Hq�\U"������+��<ļP;��W;�;<]�;#L�=�C�>#�>�,�>�J�=Tɪ��l)>%��e�M����=_���]TD�:�d�B9t�Z:(�|�#�m{K>@IQ>�b��M������>ѼO>�p@>���?*`{?>�
��ZԾ'�����H��RU���=���=Y�R��M@�b�`��7R�Q�پ#�>q�>>��l>��+�pG?��s=���a5�7��>������� ���(q��+��Y矿U�h�~F�B�D?���� �=O�}?8�I?B�?�V�>,͘���ؾ��->�O����=JF��s�������?��&?�^�>�g뾂�D�.��8�<��>�Ά��uH��Q��J5!�+Ҷ������>�A��P��#�M~��%���8���R��+�>�D?�Ӝ?��N��Wi�w)/�5�|��<� �>��j?2�H>좬>�C�>��W���@���þ8��=vu?m��?y��?Q�$=Wz�=�����\�>u�?�	�?�[�?�d?h,��2��>���;�i>>����ٸ>L/>K�=�m�=��>ZI?���>}���l�l��>I�$�G�Ʈo=���=�T�>�{h>���>��>��<��>W;�>p�>Y8�>F[:>g��>�z�>�������v?��>�y�>��6?�+k>`�=���|�;Tt�:�`�#�[����]����=�`6��Y��G*
�3Y�>/�ÿ��?��]>���_]	?*�[Yd�k=R>=�V>퓟�W��>M0x>w�S>�l�>=,�>-�=�*y>�>� ߾��">�\���"�ZaP���\�(���$�S>�1���N޽n� ������r`��{��Hd����<�B����<ӈ?�F��|�S��#��pڼ�?%�k>�@&?D`��B�����'>*��>�h>Nw��S��i%��Kg�4�?"��?�_]>!��>יW?s.?�71��+<�*Y�h/t�w�C��d� �_����#��=��Mǽz�^?l�y?�;B?�<w�~>G�~?�\&�"+���ڋ>�E-�8�tX=�(�>U��/�e�N�Ҿ��Ǿ����N>�Yq? =�?��?��W��z2���=��F?pl=?��{?�6B?��/?��+���)?gv>-,?���>�>?�M<?׷
?�>Jz�=k�;����������������ν~�,�̷=Q �=�2�<��/��g�=�Ks=�_�e�C=M��=�������<�<��\=q��=�W�>`�]?Љ�>�І>��7?���-8�����P�.?[�+=����IO��Q��� ��
>��i??��?�pZ?��b>�TB�mPC��V>m��>H&>"W[>��>��E�DЈ=̓>��>{z�=��F�|���r	�ޑ���x�<�>eS�>�4>���9>�r�����b�d>���:﴾�����S��\A�ӄ����?'�Z?٘4?�<>�涾�c;���z��$?�4?�G?/��?r�>����`9���b��,�%p�>�Q�=1j��I��<K���k��y���h�=O����ݠ�SQb>���o޾�n�cJ�����RM=��SMV=����վ�=�2��=�'
>������ ����fת�s/J?|�j=ds��T[U�0p��8�>���>+ܮ>ٲ:��w���@�z���3Y�=���>Q�:>~�����|G�5��ǅ>R8?��m?R�?���hd�wI��B˾מ��.�D�?c�>��?(\&>g����VK���^���3��0�>*�>�4"���W�"ݢ�H�ľ�"�S��>�=	?t�%=D��>`�;?�<?��Q?�.?���>.բ>pٟ<�T��R)?�S�?1�]=���Be�1�6��M�E�?ME0?}]�cg�>|?X�?R�?{xA?�?N?>�n󾫾&�&�>ݪ�>��[�qe���5>�@?��><xL?�;�?��>#���]��-��zf�<�,5>�g=?��+?�^ ?�0�>��>�����aN=���>Ra?�3�?�7m?�C�=D�?Y�+>t�>R՞=�}�>���>~�?2CM? x?��N?C�>B�K<�Ժ�,8��|��`���Ļ=g<�T;=t �6|��-�<�AG�<�q�����h3L��v��Y�đ���E��n�>�t>v����0>J�ľF=����@>mS���1���ۊ��Y:�]E�=ف�>��?G��>�P#��@�=���>.7�>z���+(?v�?F?g�;I�b���ھ\�K�z�>�B?e��=�l�—�*�u��.h=��m?��^?s\W�8-��+�b?+�]?�g�=���þ�b������O?��
?��G���>��~?5�q?��>}�e�*:n�	��eCb�v�j��Ѷ={r�>�W��d��>�>�7?dO�>{�b>f(�=Vs۾^�w�$q��J?F�?��?y��?'+*>��n��3�R
�,͏�ʅ[?$w�>�C��gR?d��.ܾ�����A��]�Y����璾��q��7����O��e�0�/1�=�?�d�?٣u?�KM?����y��a[��%}��e`�ؚ�#%%�K*A��:8��/V�]Ą�M�&���	�D���>�4f���?�2@�?S%?�2��?Kf���2�Go¾/�
>��w�N�����=����˓=1�r=��[�Y9m�o޾��"?�ٷ>�]�>?[(?�Y��A�N�9�W�?�q��#W>�"�>X��>=
?6D��i~����o��U����:u>\_?��L?�Xp?����4�����
B��s�d����K>��1>�Ē>هc�1�=���,�}�A��Uv�$��2�����t�=��6?aF�>�ҕ>Ɣ?8��>b��i����c��Y6����<�>�`?�*�>��>i�׽��*�a��>IƂ?��>��-��[����Kx����d>G�5?%TC>S�T>hc?/�U>�{I��F��𧖿P{t��� �.ڛ?�'Y��M���Wn>��\?�J�����G��>->p��1�J�ɾ[�ý6MC>՟�>�G�=�.>_p���ƾ�n�K2���*?�)?�<��n�*�+Yz>��$?I)�>��>���?C�>8٭�ǣ<T�?f�X?�D?�`=?c�>���=�I��t#Ƚ�;3�w�	=���>��j>m��=� �=Fh-�K�s��[.����<B�=�߼ZM*;$��þ=�=�E>fۿNYK�N�Ҿ<�f��]
�4ʉ�T�Ľ8����I�����Ę�ȣn����(!��)T���e��ߒ��.i����?���?s���䊾H���ł�C���ox�>zɀ���L��L�����G�꾐��&��R�Di�2
^�N�'?�����ǿ񰡿�:ܾ2! ?�A ?>�y?��9�"���8�:� >�C�<).����뾬����ο3�����^?���>��~/��R��>ԥ�>�X>�Hq>���}螾(3�<��?6�-?��>��r�,�ɿ_���¤<���?/�@��A?�w'��s��T=H��>;c
?g@>f�1�S���{��e>�>���?mm�?k�I=�FW��@�1if?�y<�G�*��4 �=-�=��-=ݝ��lH>/�>	2!�:D��9ά0>�T�>��2�?"���]�n*�<�a>8(Խ<+��0|�?�	B�3Lr��w0�5ߑ�Q`=��d?ċ�><�=��9?��Z�*+ڿ2錿�V_?�D�?�l�?1?��K��l6>��输 C?��Z?	��>�t �rav�!L�9��=c�<9��}hB���=P�>{a�>��	������PC˽Z?<���ƿ��$��d���=��<���Y����n���"S�$���n�6����m=���=��Q>//�> �V>��Y>mJW?�k?!h�>��>̥㽮r���ξ|���7��o���:���<,��:[�V�߾n	�D������ɾ�=��=;6R������ ��b���F�#�.?�x$>w�ʾ��M��-<Doʾa���]䄼[好�-̾��1�� n�&͟?��A?������V�����U�����S�W?�J�	��X謾��=����l�=>%�>C��=���R3��}S��4>?D�&?ۃ߾�����:">@��=��J=��?.�?���=�?J�?O���w@4����=��/>O�?h1?L
Z�Jϔ���B����>S<[?��<���N��>�<�w����#��xv�<�F��@㽉&�>$l�˿��?>�}=S!7�O9X?��>T:'���!�w�����%���<�Mv?�]?��>��v?9�@?�=�!����K�җ��"�=��^?��_?��>M���!iӾ�y���?5?�4l?�o�>�$��f�뾾$�{7��+��>n�j?�\(?)��xo�ǟ��*��?E$?��u?NdX�Z=��%	��Rh��(�>+?���>�D����>L&;?�:X�'ݕ�W��� j1���?@H�?\�e<!��9n"=zW�>�&�>.,%�"랾�}W�Ռ��jځ=�W ?B՝��ew��v!����ۘF?ه?���>oz�Y���{��=����?0�?g�?o۰�>g=���i�r.����;��>����௼[�ﾁG0�6Y¾4.�N���������>�$@�H��JN�>�$�'�˓ӿ�^v��Kݾ~ i���?]Ƣ>bz(�-���u�0x�-�O�׾?���!��Y�>��>���������{�7o;����B�>(Z���>,�S�;�������O2<�ْ>Ԓ�>[��>o+��ɽ����?�A���=ο譞����X?�a�?[k�?�x?��><�v��f{�����G?Y�s?� Z?�{$�3�\�Ũ7��j?i_��dU`��4�jHE��U>�"3?C�>>�-���|=�>���>Mg>�#/�u�Ŀ�ٶ�U���N��?��?�o���>n��?ts+?�i�8��b[����*���+��<A?�2>���>�!�)0=�OҒ���
?N~0?&{�b.�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?UȨ>{Br?Ig>`?u�=����Y���<>*�;c����$?l�S?���>�_�<i����C�UkN�VCe�͙Ǿы8���>>�`?8�P?�۔>/����NB��p8��B���ǽ�P༃_��o��Y���:�=��W>�I+>FJ������?Ep�5�ؿ�i��(p'��54? ��>�?����t����;_?Pz�>�6��+���%���B�]��?�G�?=�?��׾:S̼�>2�>�I�> �Խ����O�����7>4�B?S��D��u�o�z�>���?	�@�ծ?hi�f?��ྡ���e���	���þ�A�>��(?<#��ے>��>�ҽ���DЮ��q�m��>�@�?:��?�O�>�?`�p�^���=���>ő�?7�B?j*<���8��>�O"?�3���n�ھ�;�?z�@�
@��p?Z1��Qڿd쩿����e����=fnd>4n�>�i���>B�,>�9��A���\�>��?e��>Ϥ|>:�>�m�=���=�@���!��&��*��ggW����(q�!m����;�]��8Ҿ�ZʾEbݽ��Pݼ��!���&B=���=�~R?��S?�,s?RT?m�R��>U^��h�<��C�	�m=Z=�>�1?��I?�r)?��=�����Ua�!�eЦ��_��M��>q�F>���>Y��>P�>9+f�s >>�I@>��u>�>.�l=�B��<�=I>y�>ں�>J�>}C<>��>Aϴ��1��_�h��
w�)̽,�?����B�J��1���9��ꦷ��h�=Fb.?|>���?пh����2H?+���s)�߹+���>~�0?�cW?S�>	���T�L:>����j�$`>�+ ��l���)��%Q>ml?^f>��t>�3�nE8�*jP�Y����%}>�>6?�a���a8���t��H��޾i9M> Ѿ>�%C��;������Z���i��w=�I:?5�?�'��GN��{�u��4���tS>:CZ>hV=Ź�=8�M>",d�9�ǽ>�H��(2=΍�=�(^>�?�8>��-=ͭ>����2'����>6>>�$>t65?��#?���󤭽�σ�T80�>��>�?���>���=T�O��=`��>�q�>M�*<|����q�'OW���H>�6����T������m,=�{9�=i>�=�����G��MI=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ}h�>�s��Y�����\�u�r�#=���>�9H?�T��P�O��>�aw
?�?�_�Щ��t�ȿS|v����>�?<��?��m��@��.@�.��>ˢ�?�fY??oi>�c۾ZZ����>��@?�R?��>�9���'���?�޶?��?��P>d��?6q?���>ά�/�&�=����ay�ک=�YټyG�>��@>�	��l�C�'A��{≿o�m��o�/{>�5L=%4�>�w������ ��=zUϼ������c����>r{w>�->���>.4�>���>	�>��^<-���3F���y���K?���?,���2n��N�<[��=.�^��&?�I4?j[�m�Ͼ�ը>�\?f?�[?d�>8��L>��C迿3~��P��<y�K>$4�>�H�>�$���FK>��Ծ�4D�ip�>�ϗ>�����?ھ�,���S��HB�>�e!?���>�Ү=#�?�R-?Edk>�\>����{��>q�X?���>v�}>a�P?g$?�q��*9����Dқ�E�S�ܨ$>�q?uB?ڦ�>����ꛧ����y+ <V���Å?6E�?��=�/�>;�?9�%?o�?4�D>�����`��!�=�k�>��?3���R@��&�!i��V
?��?��>�ν�n��޶=����~�&�?��Y?<#?4M��"d�ֽԾ�@\<�־�xF�>�v<A>��t*>�6>\����=���=���=Z[��)��P�;ñ�=|��>+ �=��1�p����+?`���m����=�ru��H���>� Q>-Qľ\�]?�S��f��mO��i���P[(�35�?�.�?/l�?�nϽk��>?8�?�D?���>v!��r޾�WܾE��9�k�w-�՛&>���>�,�\���樂�ڪ��s���x�\����>�Q�>Ԕ?�?��`>s�>:楾�*�����{���Z� �� �0��$�>��f����n2���v���¾X���r!�>�������>�?�Xr>��o>r��>}�j�Ʋ�>A�n>V��>n��>��A>܈>�p�=�B�<cm��KR?�����'�}�辥���c3B?�qd?[1�>�i�2��������?���?@s�?�<v>�~h��,+��n?�>�>A��=q
?hT:=H3�X;�<V��3���3��:� ��>!E׽� :��M�%nf�gj
?�/?�����̾Z<׽b�����=�|?���>�v1��_�*�e�'�J��\�_�	�O.���?p��ξ�Xh�����x�������F���>z�5?�,�?`̾��#�ѽ���~��]���>�>ٞ:>B9�=�Q>��:db����"F�����u?%E�?�4�>��%?߰6?�'�?�#�?y�>XOk>�����>���y�>~8�>��?
�?�&?�?��2?Ž�>e@�4���qѾ!�3?�i?$%?���>[�>�夾08�ݭ���]�*;U��b0>u��=d��=`3������,�㲦>�[?>c�(8�����j>�u7?���>���>�e���π����<1:�> �
?Q�>� �#yr�a�/�>���?f��*\=X�)> �=�^��q�׺$��=�ȼ2�=��}�Ph=��"<D-�=�Е=X~��V��.��:��|;vv�<�u�>6�?T��>�9�>�8��H� ���� ��=�Y>�
S>�>�7پ�z���#���g�Jy>�s�?y�?��f=V�=\��=�u���X��z������<ܠ?�N#?�YT?��?��=?�i#?��>)�/K���\�������?n!,?��>��q�ʾ��ى3���?{[?<a�Q���;)���¾3�Խ��>�[/�k/~����CD��݅�������(��?�?�A�N�6��x�ӿ��6\��x�C?;"�>�X�>R�>2�)�g�g�l%��1;>���>&R?7�>�O?�y{?��[?m�U>�{8�	������[?�w�>-�??���?���??wx?DQ�>ϛ>�*�h�����	1����U���3JR=8QZ>��>>N�>3X�>���='˽K��>�h��=�bc>���>��>���>��x>l��<H�J?�W�>�+�����&7���~��͖Ͻ<!�?�K�?_n(?�O�=����6�(��>���?٤?��*?��&�*��=�G;T���E�����>29�>u��>�aἺ�=E��>�N�>��>��������)�pH;��?H�P?��=�ſ��q��p�J���3f<�ْ�?�d�����"[��R�=����$��fɩ���[�����k���c�6����|�S��>TP�=���=~�=,U�<$wȼ�z�<�J=�e�<�U=�Zp��+o<�8��GлH���	@�;\<#�I=Ve�*q¾�v?��N? �2?��A?�S>[��=3ns�]Y�>O梽�?\�i>Y�K�0�����^��`��픠����Gվ�U�3���>�`�T�,>bI>���=��<C��=��<0K,=sA���{�<�t�=��=��=p$�=��%>h��=�x?o�g�n���2[�t7=�'�?� ?��E;���s.b?���=���g���}���|?u��? ��?�"*?}T6�9_�>�l�����<�=�T�Ey>��<�sE��*?8�X>�,$�w9��Y�����?�7@�/>?/����Ŀ��g=�%>Ġ>��G�f�(�M���ٽ�����%?�E�e����Y?ӡ{�Di�&/��R�={%>�==?틾ޚz�ǣ<��Q��=��>�P�>/�l>+�j=�ϧ=�\P>��Ͻ�C�=P�>��k==m���lɽI�*���4>��u>��=��>s�?�0?w:c?[��>��o��Ҿ�����>t�=�X�>�x�=d�E>�R�>$=5?>#@?l�H?�&�>��=
��>ʎ�>�/���p�|��¡��n%�<�?�?�>��}<ə7���L�?��ܶ�7`?��1?s�?���>D���)��g�%�M&��Б�7�(>%k�>�*����g>��e>�s��z2׼*ء>��,?��$?E�>;">��+=��>+�>"M>���=�m>�%�=����<��)�=mO��]ǽu�=D�2=�.�������vK�<�Թ<����v����= ��>�=�k�>���=�ͭ�	S>����?Y��k>旀���G�]k�l�r{����">��>��K��D�>�mF>Q�>\f�?U.�?h>_��o�־�2��(Ӂ�0[���>9&�=����G��N^��.[�t����>�)�>!��>ޞn>C�+��]?��p=�P��<5���>�t���y��C���p��#��H��0i��Κ���D?� ����=)~?g%J?���?J��>�R��ʍپ+(,>u�����=��]t������?��&?��>��<|E�Ėɾ(=��(��>e$���Is��馿�g!����5���՚>/1 �\ZվZ'�(����]��JmI�����"��>+IU?���?�Y�����e�R��)�*}��wP%?R u?տk>�?u�?�����-��I��^�0>��?���?���?{5��ƽ=�l��eK�>.?���?K_�?�q?2)G�<�>V;�:�>����4��=�>3n�=�/�=�?�	?��	?�b��=���7��eBd��m�<��=��>i�>ws>G1�=��=Ο�=�&[>�a�>�>�>�`>�ѣ>�<�>�������a�?.�'>�ǚ>J&D?@|�>*�*>:����װ�כ=a�O�;5��M��-ڠ����<�F=�0�������>[(��MC�?&��>tE��P'?�m���)m�!5>���=����c$?b��>��9>�I�>Sߘ>�=�^>:]9>��о�	>���!��A��|Q�zB׾u�>ל���-��3���/0F����0V��j�B-���n<�R��<T��?Y���wj��B+�HI��b�?B��>ׄ7?h��"����e
>j��>!�>�y��Z�������Uᾶy�?���?�;c>��>6�W?+�?W�1��3��uZ�-�u�b(A�5e�;�`�x፿����
�����_?�x?8yA?�P�<�9z>A��?��%�$ӏ��)�>�/�';��><=Q+�>*��K�`�g�Ӿp�þ�7��HF>|�o?,%�?gY?5TV�s��NpK=�v?��n?��?��>?�?�Ͼf�?}=�=�>2��>�C:?�e? �?�M>b�=}u�<��<�6N���L��"��Z��2y|�P�I�<,�.>7	>+>`�=�l�=��=�@�=�6=�(����L=�?��I��>ZoX?���>�d�>�b6?[���.��8��G�'?��=,�l��z���S���y���=�f?�?��a?�0>v�J�e-D���:>Y��>.�>>^?>;�>n��F1?�-_m=�>;��=7�=Y���ic��}�A�����;%>�o�>6*~>�νU�>�����v��t%�>�--��T�8�ԽV<��}H��'̾�o�>_�\?N�)?".�=��ؾf�)��q���*?5"/?�8?_=�?��=>�ھUi/���Z�-K׽W�?�|*>����� ��y����Y��M����<�ϾѠ��kb>��Ya޾?�n�J����s�L=�w�/�V=8���վ�����=�
>8����� �.���Ъ��'J?��j=vh���QU��n��\�>���>��>W�:���v��~@�ߘ���+�=>��>�:>\?�����xG�D=��T�>�C?��?��z?W%���{�g�c��<���.��!�>SP$?�À>��>��P>PK=��ϾH_��uz��]��?�>%�?�����d�WUԾ�������A��>��	?ێ�=J�?l&^?�X�>~-l?�,?�j�>ʗ>If3��B���B&?��?jm�=t�Խ��T��9�'F�K��>@�)?�QB�|˗>�?޹?A�&?QsQ?l�?�>� ��1@�>�\�>&�W��^����_>ɢJ?���>�:Y?�̃?�=>��5��Ӣ��a��֍�=�>��2?**#?f�?I��>�	?6Oľ�>r?��?���?�a?`i�>�e#?��X>-�>e`߹6>��?�o=?8�p?$�?�4?e�<>��=]V	�U��3�<�/o=5�»�S輵뤼U�ۼ
 >�ѼD�A>�ȥ=߈>� A=W�qN$�?rս�ע<�a�>�s>$��\�0>4�ľ�d��W�@>����Ed���Ȋ��X:��>�=nG�>��?um�>�=#���=�Ǽ>�8�>��b(?��??��#;v�b�a۾��K�r<�>-B?�f�=��l�w����u��i=D�m?@f^?��W�X,��n�j?�1p?A���dW�1��d��C��P?��#?Zd��q>�}}?F��?��>
��3�z�WI���}\�=���^��=�?�>��(���_��Z�>�aV?;��>ʃ>`�2>�!վ㈿T���@%?�Ԉ?�%�?f�?���>&r\��Hѿk����Z?��>Ȣ��ѽ?��!<�8ǾuƆ�ݺ~�;G򾐟��Հ��3��������2���!Խ3�==��?�%r?:Zu?XGV??���n�e�u�W��=}��4R���۾����?A��~B���M���s����p�[,ƾ��<�p��C�!Z�?9�(?`U$����>ʯ���ܾ���h�U>������S�h#�=�BX���=�ݣ=3Mg�K)"����K?z��>��>��7?��W�VUA�K,��_<�!
����c>m�>S@s>�,�>5���Q8���ٽv��xh����ٽ�m�>g�[?M�`?�T[?ʘ8�w�K��뒿�.�k��D�L�n>É2>x��>N�Ƚ+M��%w���C�)��,�����8'%��*�=U�I?���>���>Y��?H��>}��8,��xJ�7s�R6,�b�1>/�6?WI�>xϰ>^ H<�����>�3k?�U�>���>�&��o%���y�nK��@u�>���>:d?3�o>%�E�8m\�|͏�q����2���>�e?Ñ����k�Mڒ>r\O?Dvo<�
`=��>������d�5V;�7> d?J�=�_>6ʾ��)\}����t�*?�??/j��i�,���>4$?��>�i�>���?�$�>V�Ǿ$�"<�4?�g]?�G?�m<?���>�R�<+Y���ɽ��&�B�8=BF�>�1]>��t=¡�=bR�.\�9��4<=�ƾ=�m���L�h<�B���V%<�S=$�9>�ѿ4�D���Ǿ�����Q�P�������S�2O����C����^.R��dD��?��x��X�%��Jp��;��m�����?L�?g�4�n����ؑ��gz��` �g��>LuA����<�\����Y���9��`P�A�@��vd���|���r��'?(���@�ǿ�����6ܾ5" ?�A ?X�y?��Þ"�Q�8�>� >���<.����뾦���6�ο����!�^?���>�
�R��� �>���>n�X>�Gq>=���螾�)�<��?)�-?���>ܐr�8�ɿ����ȳ�<
��?��@P}A?��(����V=���>|�	?��?>�Q1�eH������R�>i<�?
��?�{M=?�W���	�-e?�c<y�F��ݻ�=DA�=2R=����J>\U�>w���SA�{>ܽϷ4>[څ>ކ"�ʫ�W�^�2�<�]>��ս�7��5Մ?,{\��f���/��T��U>��T?�*�>U:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?$�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=�6�"���y���&V�v��=Z��>`�>Â,������O�J��T��= �뿬?������5ȾW=���>��=} ��񦾔��.�����KŽ��>��>�H?@9�>��>X=σ4?�wB?��y>Fe>�]��{���J����?�ﰾ������g�`��-9�����(D���i��k���bo���!=���=�5R�s���� ���b��F���.?\r$>�ʾ��M�м-<�pʾ@���tʄ��إ�,̾�1��!n��̟?��A?����K�V�I��d�r���g�W?pM�e���謾���=~ñ�j�=�"�>��=i�⾹ 3��}S�"[2?�"?O�ž鏘��.>ժ���g;=ǣ+?��>vM<��>|k'?�(�T���:m->MX
>���> �>�
4>䕴��l��](?�U?�F�9O���}�>.Ǿ"�d�m1�=��>��&���1��V>�|�<�ݍ�%��������<�6Y?�Π>�#%�� �����2q>��e�<^�x?�	?��>�Uf?��D?ʁB=E�UV��}����<�JM?5;n?g>��-�h-�h����=?͸n?��L>T�e�[о�}7������?Z�w?��?v�d�̂w�퉌�bO�x�.?pv?r<\�����0�͔=��ӥ>���>?(�>��3�:�>�C?�@.��I��t9����0����?��@�3�?�5�O&#����=�x?>�>TA���ľ	��%񮾚O<=&g�>�T����w�^�!�
Z&��-9?��?���>�ކ�Ś��D>������?;o�?�&�������hL��Y��$.>�r�~~���K��7��l���⸾�� ��ľy���Ʒ�>Lt@y�K=�I�>[G��V2ܿU�ٿ�c���Bƾ�,�F?F(�>�9ܽ��ʾ�>��~��ywZ��Zg�����IH�>��>2�������e�{��r;�ZL���
�>���Y�>:�S�(��ᘟ�/q3<�ݒ>���>���>�7���ڽ��ę?�Y���>οѬ�����&�X?j�?mn�?p?"�9<A�v���{��X�A-G?U�s?�Z?PR%� ]�u7��c?��8� b���M�@q?��n�t+?��?�JV�b�]��ԉ>Q&�>@曽�MT�ZgɿJ衿}R��eK�?�^�?���L��>��?6?�\� m���o�6��Ʒ >o�f?4��>H����|F�-��S%k�4�?O�D?�G4�=�%�]�_?+�a�M�p���-�x�ƽ�ۡ>��0��e\��M�����Xe����@y����?N^�?i�?ϵ�� #�e6%?�>d����8Ǿ��<���>�(�>*N>oH_���u>����:�i	>���?�~�?Qj?���� ����U>	�}?SZ�>��?Շ�=s��>B�,>��l��<\$>i�W>س��NJ�>i+_?�|�>�
�=�#Z���@�@�C�0 I��_��C	?��z">�?�a?x�I>.��������$��q&�T3���B=�>X�QP��~�0�>a>N>]b>^A�5Ѿ���$?Ąܾ�F��Ŧ�4����3?���>?�*��B���<"$X?�5�>R�:�1x��ꙉ��	H�%T�?��?���>a�����ͽ�>s��>�4=ۆ�����=��Ծ�(�8�K?�N������h�|r>�D�?��@�A�?�S��_	?A��Q���b~����7����=U�7?�6���z>)��>|�=�nv�f�����s�.��>xA�?�z�?,��>��l?7o��B��2=7N�>��k?go?��n�+�}�B>�?;�����/J�af?��
@Au@�^?�տ����LR����G�pn�>}]�>��y>!4��'8>9	Ͻ*#���G=.f�={`�>�~>�=�>DP~>��P>*��<����3�!�����B�����=����߾�K��>���'J��d�-�W�Ѿa�������É�=�*½ۥe�ӎ��>�EH?dud?�w?\��>��aӻ����߈�;z���r�=��>��&?�;?�?�U�<����h(p�D�s��� *�>�~�>���>���>"�>2��8�O>�Ո>Gb�>^�=�)�;L'��}Rü�sY>��>�]�>�ڶ>�C<>��>Fϴ��1��k�h��
w�q̽1�?���S�J��1���9��Ӧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��u�T�3:>9����j�5`>�+ �}l���)��%Q>wl?(�f>�u>4�3�d8���P��{���h|>^36?0趾�A9���u�ݲH��aݾIM>�ž>��C�ok�����`��ti���{=�x:?ʄ?�6���ⰾz�u�>D���OR>�<\>,F=�d�=�WM>�lc��ƽ@
H�P.=��=Ŭ^><�?�&>�y=�I�>H��fp]�}�>z�]>s>��=?��!?y�Z�g�Ž����Q�6��&p>�k�>Z �>V�>P�Ih�=M� ?��g>շ��m����:V�Y�k>ఆ�Nvw�5Ӓ��&�=�ڇ��>{��=���(j_���<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿˈ�>�!��l璿�I��Z��:�s<�5?F:(?K�޾�xB�Fy�>y�?@�;���,���%�}�J��>�f�?�2�?�fJ��а��"U��@�>]��?*�?hҪ>z^�9`þ{�X> 	? �]?@��>�_ ��@��/?���?�V�?�%Y>���?�*~?F��>p�׽9�<��C������&��=3Т=���>��>�m���o6�\B�������gl��'��|Y>tY=���>"��`�ƾ���=����@D��N$���>nn>�rS>�Ǵ>�<�>���>T֤>S�=\�	�H��J����K?:��?w�[�m�	�<Ϝ�=�b��?t�3?��J��ξ���>9�\?��?^�Z?_��>���Q�������l��\>�<&rL>O��>(��>.`��5L>��ԾfWE��&�>-C�>M:��(ھ ͂��Ա��*�>�b!?���>�y�=�e(?k�0?��>ԓ{>�j9����!p:�¼�>���>C@?�r}?�`?������M���2����U���G=�$z?l�$?G��>����@���p�=�d=�PȽjڇ?=�b?�Y־R��>z��?	nK?zB?=D��X��@����<��>�!?���A��B&� ����?O?��>���A�ս�k׼.���a����?"\?}6&?��&a�~�¾bk�<�g%���I��y <��D�O�>��>.������=;>�P�=dfm��-6��5g<y˼=ƚ�>9��=�E7�����Y+?�A�<����'="�m���M���g>�p>]�ǾϹ[?X�	�p�23�����O����7�?i��?.C�?����Yh�J�2?L@�?�?���>�C��.�����}<���F����*>`��>�L<��¾Q���4��Vބ����Rs�L�>գ�>�� ?���>?:q>�w�>� u���r@پo�о�dU�L����1��&�H&#�2ڌ��Ľg5!������L���]�>;b*=�>��?+��>�ʃ>su�>ŸI��q>s��=���>X��>�>ʀA>��8>�α=�Q�PR?&�����'����됰�U:B? kd?�4�>�g�胅����w�?X��?�j�?v>��h��)+� [?DU�>P���c
?;={����<�H������w���8�Ĥ�>�6׽�:��M�hf��h
?�)?E��u̾R�ֽ7���Ö�=vs?3#?й9�p�S��j�=�Q��8B���3� 2���2=Z���������Qi��R��-y:����G�&?h�?{0��0-�i���Ra���%���>�?���>5��>Ā�>P��H�Q�<�V��j?�嵾��3�>^�?���>JkI?�&<?y�P?UNL?"f�>�˨>GC����>9��;��>��>D�9?��-?V0?�K?<+?Pb>����y�����ؾ��?��?�l?9-?u�?�r����½}���b�d�y��ˁ���=�2�<#׽�tr�4�V=)T>S3?Fi >�F�̨&�d9�>�P?���>�9�>7qg<����q�9�ܶ?�A?0ދ>@����w��f���W>�c�?~lz����k>�H�>��G=ط�<��E>�w��Y��<��T��c-�'S�=�Y�Xf<�z=?�<X���u��=�>���>��?u�>��>�Y��� ���ױ=b>X>S>��>pپ����$���h��y> l�?�r�?��g=V�=�H�=v֟�d������὾���<�m?�p#?J~T?!��?r�=?^P#?}H>���9���G��	:����?1",?���>����ʾ9ҋ3���?�^?�:a�����2)� �¾�.ս��>a/��+~�v��"D�5:��������Z��?ɾ�?A��6�Ձ�;���(H��ƙC?t#�>�U�>i
�>�)��g��!�e3;>R��>�R?�>�?W?��?֒G?�v�=|�T�BF������٢�<���>|[=?��h?���?��t?s>�>)�=\��7��}b���L�E�.�<��웒=� I>Ɇ>b��>�>�+=�{5�a佬�)���=�;^> ��>�U�>~̺>�x�>�O��ZE?_��>eS徛?پҞ<C�ֽz�9=�'}?_Q�?�xP?�e�>�	�K"b�Q��Ġ�>��?���?0�W?��߾���=��k�p;��f|�z��>��>1��>�ő>�eX�o�>h?C��=D���g�����Ӡ:�?��B?rW���xƿ��s�p�y+��TK��匾[�N� ֽ4a�h�?=���\�'��+����?�9E���h��{���5����|����>M҈=	��=��=kk&<�1ؼ%�{<��v=�	=�n=ǘd�'e:=ɽ/��WŻ
T��=t����<�Ga=�f9y����jh?7.Q?0/G?��9?��J>�S�=����L��>G�C=�?g�4>ߨ>�~�����>����ᖾ�a�}�̾��U��훾���=�h��N�=�K>]*=>��7� >�~�=d��=�E*���Y=&�>j�==�==�>��I>��>�,q?��m��%��e�!�u�>L�5?_��>�\�>��\�(�@?�U�>��U�ſiI�*K�?K��?�!�?��!?m�׾��>�"��N��<j >��<��5>�>��0���>>E�<�����bK���?0� @�?b&��H�п���=X�6>��>��R��%1� \���a��MY��V!?�;��5̾�>�	�=�a߾^lƾZD-=�E5>�d=;�,�[��(�=~�~��w<=5�n=hL�><}D>"�=UЭ�kH�=��H=t_�=i+O>��m�i�.���%�?95=�q�=E3c>0�%>���>q\?>C1?��d?�ŷ>�o�c�ξ�`��9[�>K��=g�>�3�=��A>���>Ŋ6?��B?��I?�Э>�r�=ꓻ>���>��,�Kp�|W�)����d�<��?s�?�>k�{<4�;���Լ<�P���:)?3�/?�?���>D��=ؿa������{u���(�=�*>����l��W��߼پvf������c?� ?V�?��>�*�>s��=��>p��=ł���_=�P���0�wiq�|�0=h��$Ov;� �<���D�=��=g�<w�=���<OVX=�	=� >9��>j��=Z�>�M�<ވƾ,6�=y�O�"~F�1�=� S�)�(���`���}�[�6�{ {�3�3>��]>W�H�_W���մ>m�>T3�>P��?��?xb>bv������拖�~!��!�s�
QV>��>A�<��3�Jl^���N�c��1��>M��>��>�Lg>+�+��y?�2vm=�+߾:I5���>	|���3�f��o?q��$��Ì����g�T�&:��C?�7���r�=�D~?ċI?-��?ɹ�>h���׍ھ��2>~���H�<%����j��D��@?��%?ē�>ND��D�T�˾�5�����>�3J��P�h̕�A�0��%�y綾Cȱ>}��W�ξ��2�`ᆿe��ܝB�/Au���>��O?/�?�E`����1-P�Ee�9����?�Pg?�W�>�?o�?����E뾺�}�i�=��m?;H�?�3�?�>��=	h��At�>*?�n�?�n�? yo?U0)��s�>���:>�!>2�ɽ"�=[�>��=K֥=�	?=�
?Z?�2����O�U�ƏX�K�=���=0j�>�z�>�ii>��=�,=5��=?Y�>W��>zR�>k�t>�ɦ>�4>Z����
�f�?s+*>��t>S.?i�>��>�O��5��m;�U��� ���[#<��;U�g<��~=��>������>�ٿ�lT�?aJW>�����>�Lվ\f�<~��>�ߠ>�v�>wJ�>�Ȁ>K�?��?��=?.>���=6�ľm�3>܎�Q���O�c�Y�b�־�_^><>����ڽ
����@��T�=��������ujh�����`;;����=�?�Ď���q�}h@�<eI���	?ۿ�>�28?�"W�Ⱥi����=�P�>��>�*ܾ�Ò����z�ɾlƍ?7�?p:c>0�>�W?�?J�1��3��uZ�5�u�`(A�?e�z�`��፿	�����
����_?�x?:yA?�P�<*:z>.��?��%�dӏ�s)�>�/�';��B<=�+�>�)���`���Ӿ6�þ�7��IF>l�o?+%�?`Y?�SV�Dg��@&>��:?.�2?+t?*�1?�:?�"�ސ$?�H7>H�?��
?��4?M�.?:�
?��1>�:�=���W�!=����X����ҽt˽�����[5=bh�={��9D<g =w6�<���94ؼf{�;֟�b/�<�l==��=��=�ڦ>]?���>��>/�7?���E8�\-��N/?� <=r����U���1��
�T>�	k?F�?��Z?|8c>��A���B��;>W��>��&>��[>�h�>�c�6F��i�=�l>�d>�i�=d�L��}��Y�	� ������<��>H��>R�{>^5����'>�n��,z�=}d>��Q�湺�5�S�v�G�X�1�{Mv��T�>�K?<�?�:�=�b龏����5f�s)?�c<?QM?��?�ԓ=��۾�:��J������>N�<��P���X��0�:�^:Rs>O��m����AZ>D"��AܾH�l��pK�����P�=�D��:=���S�ܾB����S�=�[	>'㾾���5▿-���5G?2MU=��� �R�B���T>k�>y��>$Z�6���;�󊨾A��=���>�k->���,7�4�F�eL�n)�>S�D?��_?���?* ����q�k(B�L �¤�{ռ��?81�>��?�?>�5�=�G������e�$fE�$T�>��>{m��uH��y��Uj��%����>a�?�i>̈?�}R?�H
?"$_?�*?�^?��>J��rB��T'?���?��|=�|ܽ�WT��89�AG��v�>R*?��9�b�>�?�H?�"?%�P?W�?�V
>qa��>>��F�>|C�>��W�h=���c>��H?�ɲ>aRX?~��?O�J>Q62��~��7���"�=�!>�3?��#?n#?��>���>Sd���ؔ=��>0bb?ָ�?m�m?�}�=��?E�C>�K�>��=��>�� ?�8?�=K?�qp?�F?�>]�<V����e��#R�`c���׊;��<k�_=3/�9
����¼�#=5<Sm�q�(�JT�j������f�;>Q�>��s>������0>��ľ`W��d�@>�᣼&=��Nˊ��t:�(��=Fx�>��?���>�@#�$#�=���>�/�>b���'?F�?8�?�:��b��ھ��K���>�A?x^�=1�l�掔���u���f=��m?+�^?�W�K��M�b? �]?<h��=���þ~�b�ȉ�j�O?@�
?�G���>��~?d�q?5��>�e�(:n�(���Cb���j�.Ѷ=Qr�>GX�F�d��?�>j�7?�N�>�b>�$�=Pu۾
�w��q��`?~�?�?���?1+*>{�n�T4�Y������)Y?SO�>3g���&?_�_���;]-���,��}gӾf��������՗��c���Z��6�������3=�,?��t?ɭn?�\?�� ���g��lf��-}�'V��a�����;�+�1��A��s��D�k�wĂ����=V����/L��D�?<P?7�*�#?����;�0�ݾ�5->���w���)=w���60_=��{=	��%�����ѾX�(?ڄ�>���>+S8?D�U��H@���A�3x;���p[y>d�>|��>�^�>zz���g�zJ8�����?�r=��Q>S)\?iwN?�~q?h�i�*��~�]�)��C��S���q>mn>Hϕ>�bt�EJ6�,+�u�<�Ӛ}���ԯ��*7�U��=�:?ş�>V��>��?���>��S���r��OD<�ߐ��A��>�Za?>��>���>d1�dp"����>�x?���>��>BDZ��}��E����=�E�>^�=5*�>�r ?Կ�=��Q��╿綏�K�~��7<訋?m�O�ғ����d>�w_?�>�|m��j��>
���X'�ѕ����ƽ��<>@��>z���Fe>�A��9���'�~�R���E�??��?`M��/��z�>�H8?���>C�>ձ�?�D�>
������=0?�J?��>?ݫ(?�V�>c�>��x�c��1`��Þ<o��>6�E>���=�X;>��F��ˊ�`����W�<��=�м�ӽz�=3���+�= �=�U�=Yۿ�bK��1پ������	��������ض��.d���������gx�_����&�N�U�M�c����o�m��n�?E*�?����ԉ�P���㠀�l���7�>
%r�[R{��ū��y��d��h�ྦY����!�P���h��e�N�'?�����ǿ򰡿�:ܾ2! ?�A ?7�y?��7�"���8� � >~C�<&-����뾭����ο=�����^?���>��/��j��>ݥ�>�X>�Hq>����螾z1�<��?8�-?��>��r�/�ɿa���&¤<���?0�@�A?`�(�M��
V=���>�	?�?>/X1��F������T�>�;�?p��?Z\M=��W���	��~e?5y<g�F�]�޻�=AO�=ȓ=����J>�T�>ތ�AWA��lܽV�4>lՅ>G�"�3���~^�ڈ�<��]>��ս�E��3�h?��j��o���@�.���;�>��e?km>��K>�,,?7[`�ԇԿ�ɀ�x"f?��@|��?B�5?<����a>
�Ծ��Q?�sG?���>���"!z��M���o�=���vϱ��X4��:=�Fl>~��>$)��y�@�:�VT����ü��1�ƿ�$�|S��K=t��8�0Y���潯���=W�F����:o���齒�f=�=�=�Q>�>��T>��W>ҁW?b�k?��>�>���ys��P�ξ��)�^���0W��ڋ�Y���梾:W��߾��	�}F���Q�Ⱦj�>�4y�=p{Q�짏��F �r5d�A[D���0?eo>��˾��J�[��
?;1-��	S��j���ɾ��1�w�o�­�?	�??�΄�`�T�����P�7_��b�X?�&����Tx�����=)y���� =�"�>��=2��xF3���S�:�Y?3$?L@龟��K-X>���=��=���>��>���=�>�>~r1?0泽{�J�EQe>��=$��>��?��>�W���N�Le?��f?f���^��޴v>�9�t����ȅ��	�<׷n��p����=rh���R�}�����8���[�s?6H�>�+��h.�l�6���<����r�n?+�?�B?�^f?%rD?��W=����L}-�+������=�th?u�d?��">�&��E1Ӿ�ғ�s-?�R}?֊�>ha��^u߾��|���ZE?QV?J�@?[�h�H`�o�^��c侺a ?�v?�^�ȉ��2�l[W�4å>���>�O�>��9��M�>�Y>?��#�5W�������14�'Ϟ?{�@���?��8<Rc��D�=R�?Y0�>o?N�)�ž�T�����j�q=��>�f��mkv�����&+���8?ļ�?O@�><���{����=��]N�?�	�?K�����g<1���l�����l��<!8�=`3��K"�����7���ƾ��
��ǜ��]¼�ʆ>vZ@Y!轱�>28�/5��^Ͽ���eoо/Cq���?a��>��ǽ������j��ju���G�!�H�-��S�>j�>�]������{�ƃ;�{��F&�>����>�+T�g����D���-<�X�>m?�>E͆>c����^���D�?�����cο�������߰W?��?�J�?)H?�LL<�[w��|���_�7�E?a�r?9_Z?����X���7��j?r_��hU`��4�lHE��U>�"3?�B�>J�-���|=�>���>Yg>�#/�t�Ŀ�ٶ�Z���H��?��?�o����>o��?�s+?�i�8��h[����*��,��<A?�2>(���C�!�90=�7Ғ���
?g~0?h{�o.�C�_?C�a�m�p���-���ƽ�ۡ>��0��f\��J������Xe����Ay����?N^�?�?��� #�A6%?�>���?8Ǿ<�<��>�(�>Z)N>�F_� �u>|���:�uh	>��?�~�?}j?ߕ������U>��}?K��>?�?-��=Y�>��>쬜�<J��xG�=�'�=+6��D��>ËL?�)�>ޝ�=�.�Q,�R�<�6�H����� G�Mr>CXh?�^S?�L�>��н�l��$�������d��?u�UM�+�!��ף���/>�8>>ȯ >Th�A�ľ��?7p�3�ؿ�i��p'��54?��>�?��<�t�w���;_?Sz�> 7��+���%���B�_��?�G�??�?��׾�S̼�><�>�I�>�Խ����P�����7>/�B?L��D��k�o�}�>���?�@�ծ?ei��3�>��up��ʋ��-O:�)���H�> ?6O��4�l>�>�>�>漗�|������vd��M�>�]�?���?��>�H5?0T���.��3U8�R�>�):?�?�ѽɺ�D��=֢>_�*�ͧ����!���J?�		@	]@��f?�.��*���3�����!���?=iZ�=�%�>��ڑ�= e�=�=4�y�/�>��>�Ls>JE~>��f>^�A>� �=QW~���H^��b����y���8�DTܾ�"/�9��C{n�g�'���ؾk���Z���`�|2[��r��h
���J�z[�=5T?�nR?��q?֙??�y��z>� ���=�_1��n=OC�>�1?,�K?t�(?]��=3t��-)c�$K�������1��>�7H>��>���>c�>�ԣ;�LO>G�C>�t�>��=&�4=�<��<��L>p��>KK�>i߸>�5<>R�>rδ��0��*�h��w��̽��?󂝾(�J��/���=�� ����l�=Ca.?|>����>п����1H?����*(���+���>h�0?�bW?b�>���f�T��>>޸�ɡj��Y>�/ ��l��)�!Q>2k?��=2L>H�/�s�.���J���׾��>�iD?C�ھ[TR��][��X�x��g�k>V��>�������?�����������=��4?t�?�/�<,��[O�ƹV�Y�}> f#>ա.>��Z=�o>w���T�A��	��$�=>?p=�>��?��.>�T�=���>ʒ��U�G���>��<>��(>�>?�$?2B�{'��V���7+���r>&��>�@�>�8>]O��X�=���>��i>]߼����+��v�D��T>oi����a��ʁ�~Bt=R���j��=�ҕ=�O�J%C�a�!=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�g�>�v�QZ�����I�u�ȴ#= ��>�8H?�V���O�H>�w
?�?�^�穤���ȿX|v����>5�?���?��m�cA���@�p��>��?IgY?Zoi>�f۾`Z�;��>ٻ@?�R?�>�9���'��?�޶?�?g>��?�X?��<>-���p�6rU�Θ�=?��z�K>8<l>M�n�/?5��̚�����:Ӆ�������>�5�=���>�q���ý��̅=Cn;�)S�kK���?�l>�٦=�6�>/p?@ �>I��>6 �;d�S�E|����=��K?���?-���2n��N�<Z��=)�^��&?�I4?k[�}�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��H��<��K>*4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��VS��GB�>�e!?���>�Ү=y#?w�%?X�]>S��>�-@�6���,CL��e�>���>E>?��g?d�?cڢ���<��ӌ��e���X�g�N>��u?F�&?C �>�P��9i��� <�������f�?"hr?"s��e?�8�?�-,?u�,?<M�>t����ž��<�q>U�!?��4�A� N&���?3P?���>�2���ս�4ּ���j~��h�?�(\?�@&?��*a�M�¾>�<��"��U��/�;��D�R�>�>����߉�=�>Nװ=�Nm��F6�%�f<�k�=1�>�=�-7��x��:�+?QoR��!�����=��r���D�~G�>>\L>����Z�^?�V?��|�x'��&��g^R�!�?ր�?�=�?�ַ���h�.=?���?j ?�e�>A��޾�y߾��y�Oy�e��33>�n�>J�}��6ͤ�I����8��Ez˽��3�~��>#8�>nh?b7�>��=>1��>IV����,�b-��

�	gV��'�&6��[.�j�1�����a�_JD������q���>��5����>�?Fr>�'t>��>xڼ��>�0*>l�j>a�>q�D>82.>g�>�:<���LR?	����'�¶�ڱ���3B?rqd?50�>�i�'��������?t��?�r�?=v>�~h�R,+��n?h>�>����p
?�\:=�TF�<.V������5���t��>DG׽� :�UM�Pmf�7j
?z/?���7�̾D;׽�4��+�=�,s?m"?����-�ߞ`���?� ���`���`�I�1�ҾȘ\�돍���}��
w��1�`��=�D?�_�?
�n[�dKj�:Y���z����>`��>a�P��5�>'8�>Ɖ���X��dJ�^&��V���
4?�{�?���>*�4?�1?{�c?��^?�f�> �y>=e����>!�y�P�V>='�>+?j�?s?���>�i?G>>�n�Nn�4�̾a4?Ќ)?�	?L��>/~�>@1��/T�<���M��H���?R�#4f>��O��������]� �!��>�s?LP�.S9�����|o>+1:?hs�>���>�ً�4<r�],=V5�>�W
?X�>�(����p�������>M��?����4+�<E�'>pD�=m����ZE�9��=���.�r=����bM��<&{�=5c�=�|����c<�1j;�1#<z�>��?=��>m=�>�>��̪ ���oy�=Y>�/S>�>�?پU|��%��N�g��Yy>Yv�?�z�?��f="�=���=�}���V��_������E�<��?�H#?�YT?���?��=?kg#?�>�)��K���[��{��ǭ?i,?,��>���[�ʾ��߈3���?�Z?�;a�����;)�ً¾��Խ �>%\/��/~�g��{D�J�����׉��қ�?B��?A���6��r辢����^��4�C?f�>Q�>��>@�)���g�\$��=;>l��>�R?�޻>;�O?qM{?J�[?�'V>/�8������ș���VL>�??���?�̎?o�x?Z��>)�>��)�9�߾�r����<��
��n
T= �X>㯑>H�>|!�>�R�=l�Ľ�!����?����=�oc>���>�^�>b�>��w>_�<V?ab?udǾ���"��𘝾����Fy?�z�?݋E?�S�<'��vD1�N��ݦ�>�3�?�=�?4/8?�r��r>9Ɓ=L��?8���F�><,�>��>�!<=;/�=UӖ>���>�e�>��B���۾��&�`���6�?��F?9��=i�̿�f�oM�WPa�NWy<ߒ���畽A">������t<�:ݽ�̦��%ʾ�3+�&G�����8;������^��)�>L�B���>���=8��="XB>0��=�d)���=��;<����Wz>֧�<79
�L���)�<�j�<|S�N��U�ž�Sx?�M?�p1?O�E?�f>҃>�˗��h�>'n����?��O>*��������D�?H��Gꕾ�mӾ>;T�_�;Z����>u�g���>{z6>�>\��<���=7�=J[�=��e�|/m=0��=?��=��=���=Η	>S�=;SI?i.������vo����0�>�w?�'��ľ�%?dt��:���¿�4쾡��?���?k��?��.?��p��"�>�JM�TD.;X��=��w]�>bOt=�M�"�>�3w>і�R�������"W�?�@R�Z?�h�����(V>`�>���=مP�Je.��K[��8x�	 I���)?�#;�6Ͼ��>�@`=[Y徫����Z)=X4>+n|=�&�W�a�\}�=�Y���D=�f=�A�>̨V>���=D4�����=�;;=��>��\>�};|�����!/!=��=�U>�>���>�f?��.?�^b?5U�>Oto�lҾs���~>_��=��>�U�=��E>��>�s6?�&B?�BI?��>�h�=��>���>!.��o���צ���:<wو?N��?���>0�<{�;�!@�y�>�ۡ���F?��0?�?���>�U����4Y&���.������1��+=�mr��QU����'m�:��q�=�p�>���>��>0Ty>��9>��N>��>��>z7�<�p�=r㌻���<�����=����O�<�wżi}��=l&�w�+�����+�;g��;B�]<>��;�w�<��>NZ�=�`�>u$0=8��-H>��Y��Na�}��=�Ǩ��O���j�2�]�������W>�0*>Y4�ꓗ�U��>�h>��r>�*�?�>a?	�=�j�%(ϾM���� ��Rtq�6	->B(�=a���W�*
]���S�(������>(��>�>%t�>�%�M\)�&i�@��w�2�,��>�o��yr�=3��U�n����8Ɵ�r�h��F��M?%b���q<c2�?ьc?��~?ڧ�>o��=�e#�hCM<>x���۶��0@��ט��Ȉ�V�?��?[�#?R���	M�پ������ �>4�IH�w{��f�6�ل=d��@E�>�о^b��\������Y���Z9����4g�>��I?5�?������%�t�)�����#��\�>�nu?�q�>�� ?�?�L��h<�K����>>oj�?�Ӽ?��?�;�=�ݽ=i輽J�>�R
?iۖ?m��?�lr?e@�F-�>�lO;�%>:퓽�g�=[C>��=�%�=��?�N	?+�	?�$��yP	�iBﾄ��:�^�{��<�u�=m�>:�>�r>^��=�Aa=���=�_>t��> V�>�0b>|R�>�5�>��M��[z?���=�1�>.#8?@��>B	>O�߽�	P�	�w=Q�S���p��	ѽ�|ʽ�*[=�i�<����I%X�y�>B���_͏?�PE> � ���.?���g_Y�[8>�O]>�>��?W��>5�!> ��>(H�>X��;�4a>��>�Ҿ�.>����!��
:��+R������>�T��:�@�)��3�ƽ��=�@M��ژ���j����V3��=e�?�x{��fe�7x/�;νe?��>u�5?�o_��\���=�=$��>��>�쾦������ �辜~�?}��?�;c>��>J�W?A�?(�1�3��uZ�6�u�J(A�Be�V�`�o፿�����
���� �_?��x?yA?8U�<:z>G��?��%�Uӏ��)�>�/�';��A<=�+�>�)����`���Ӿa�þm7��HF>x�o?%�?tY?TV��G�$�y?=n?��?Z�(?�<?H��G?C�_���?;�>|�F?��z?���>�R�=v��<��ǽ�]���䰻�k���2K�Zt9���ȽN/^>���=V��=��*=�	D>��==GsŽn�>,
>�4V�ɼ<����<:P��*9�>ͤ]?`��>���>]�7?����n8�����>/?�;=�����e���W��\���>o�j?ë?�RZ?U�d>��A��KB��I>�>�=&>"�[>٧�>_���D�V~�=>�>���=�nE�J⁾	�	�P3���n�<"�>u�>�n!>�	�u*�=Hؾ��̾;K�>��$�U�־�����\��LL���ھe`�>wsi?�T7?
�)>��ľ�3���w�Bs1?,4?q�L?�v�?ɛǽ�����Co�AV����>���=���񂙿�j��!�m�MW���>y �}ܠ��Rb>t���]޾^�n��
J������L=8���iV=��c־�$����=�
>N���� �)���Ѫ��.J?A�j=	v��jeU�]n����>ε�>�ݮ>��:�<�v��@�ݶ��E@�=���>C;>���m��rvG�4��>�$4?��l?��?[Ď�F_�z�<�Q7�Y�ľ�/�R��>�sM>�??�>U�=���\N��h����:�>�?g�)��o�j?����оi�2��&�>��4?w�F>q�?��h?���>�uE?`�@?Kf�>�=�>!�*>Pb���l+?:X�?��=�L<��k�a%���K�r�?�lE?�]м��>�W+?d?M
?�P?��>l�=x_Ծi��E�>qV�>}p[��b��s"�>��S?=��>��H?Q�?ĭ�>���_�P��Qd���>J#2>\�(?�'?3_,?���>}�>
���ާ=X��>X�g?Q�?{bn?)>i�?PP>h��>�%�=!�>f�?I%?ǼP?�,q?��A?ع�>�B�<-�ý	ؽ��#�O;�j<�/q�+�w=(��M&��i�Ҽ`@�=Z�U<숼��ӻ9����°�O�<^h�>)�s>�
��c�0>9�ľ�A����@>q���/���ኾxo:��k�=���>��?ꠕ>;f#�fx�=9��>JT�>���{((?��?V?�� ;+�b��ھ��K�>�>`�A?�~�=N�l������u���g=��m?��^?#�W��4��U�b?��]?g�=���þ
�b������O?S�
?��G�o�>(�~?�q?���>��e��9n�!��Ab���j��ж=�p�>[W���d�F?�>�7?�O�>�b>��=�t۾]�w�r��??��?Q �?R��?�)*>��n��2�*�$�&8���X?j��>��u3
?�������Wb���M��j�������w������l�ч��3k"�Z�=�8&?K�?[r?-pP?��8�h��D?����X~`������@���E��w%���^�D����'�!�
�����9>�����F�Xǩ?�.?�^�����>�ce���ؾP"ؾ���<��������}<����M>�n�=$d<��N�2�ܾ�w ?EW�>�I�>��+?ud�� ?�A-�d&F�4z��pQ>���>��>¼?5�.��E~��`
�����ʸ���=H�W>=)H?[�T?��^?;��#!�"�r�h��Ø&��K��_#����>wK�>_��&�=���/�(g:�6Ո�x�ƾ9���f����e>�f?I�,> ^T>ӟ�?_ӌ>�K ��l����� O������>6_B?���>t��>qQ2��<���>^0n?_u�>Ѳ>��>�}
�1����%����>�0>��>]��>��K�9�K�4Z������R����o�?�t��������>�Q?�����:����>��[�5�'��)Ծ�4E�@~>a��>F #�<Ax>s��������������G8?�)?ȍ��}�O�ʉ>ŠM?�7�>$^l>��?��>D׃����=M�!?\�l?|�8?�?���>�S�=��=�g��QRC�]����k>�^>���=��+>.@�V}�z���ᙫ=.��='p3=w#���/�������S;��>[	ܿ@rL���Ҿ������`	��P���A�k����y��G˶�����C�t�q"��}��R�ĺh��ю�`�k���?��?؇���8�����v���k����
�>��~��{��u����Ƒ��G�`'��=$���P�H�h�E:^�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >^C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾w1�<��?7�-?��>Ďr�1�ɿc���z¤<���?0�@�A?^�(�}�쾩BU=���>��	?��?>�=1�H:��谾~e�>�=�?���?�)N=!�W�
��ue?Ry<|�F��޻���=\.�=W�=����TJ>9I�>�m�|6A���ܽh�4>��>��"����~�^��*�<�p]>"ֽ�@��\Ʉ?��[�9wg��.��[��	>KAU?�4�>Q�=1<,?��E��EϿT�^���_?�x�?C3�?5�*?_��>�zܾ�M?�7?��>(}&�L�v�z.�=���Ґ;����U���=�\�>�%>T�+�V���R���ѼV��=��-	ʿ%Z�V:��=�=��C;����^���	�Z<����}�\j��ܽ�`�=��->;�\>!�m>��B>�E4>�vZ?��z?��>�>�A6��%���ȾU��w������ѿ�T�c� ���9��|��}@�%u���9y��!=��=7R�g���3� �a�b�U�F���.?�v$>}�ʾ��M���-<�pʾ~���'܄��ॽ�-̾�1�%"n�e͟?��A?������V�?��)W�򄹽[�W?�O�Ի�}ꬾ��=o�����=%�>���=���� 3�y~S��x9?��"?�}Ӿ,��*B)>�k���2=��#?��?M ��z�>URH?�ё�.泼0�7>���=�\>���>�z>�g�����C�?�R`?<5���Ծ�=>�^���O�P�b�(�T<�D4��+�%��<����<��z�W"�ȁ��X�[?Ҁ�>~����2�K�向=G���+j?B&?5�?�a?p�F?O[�=�����,�d%�\T�=.9R?l?b�>��L�Ҿ�����l5?�u??�>�~��%k��2G�3B��d��>��`?q.?�i���'v�.+����2"?��t?-�S��q�����՜c��N�>j>?�D�>��Q�k��>7"d?U������ ���I���?7@��?�q��P�<�Xe=�G�>�e?� Ȼ~�^���.���a��0>u`?�
��h�]�T�'��ֺ�!�s?/��?���>r��Ⱦ@L�=�嗾��?4ǂ?}���t��<�	�L�m���	�.n�A/�={��:A�)���{�(���J��"��e[��(�>�V@��߽)�>�54��Tؿ
�ԿB���a����s��0?��>��	��;*cx��Gt�HU��J����Y�>9>�C��P����{��k;�����$�>�/��>��S������s����4<���>��>R��>�=��9������?���X=ο沞���'�X?�U�?�t�?F�?�;C<�<v��z�Y^�GG?J�s?0 Z?j�#��\��7�C�j?M]��iU`�8�4��GE��U>Z"3?�B�>=�-���|=3!>O��>k>H"/���Ŀٶ�O������?���?~o�K��>��?t+?li�18��\���*�q+�O9A?�
2>S�����!�1=��Ғ�ͼ
?}0?_~��.�[�_?,�a�J�p���-�n�ƽ�ۡ>��0��e\��M�����Xe����@y����?O^�?i�?е�� #�c6%?�>e����8Ǿ��<���>�(�>�)N>eH_���u>����:�i	>���?�~�?Qj?���������U>	�}?z��>��{?��=�=�>��=�ߗ�PI��{�>5h>�B;�9i�>r�[?��>��=�c@�|{#���B�Sq>�B4վ�]?�c,,>�x?8�Z?�[o>����П�k3�l����2�:5	�b�����-�����>�>��">#cA�)s���?Mp�9�ؿ j��#p'��54?0��>�?����t�����;_?Oz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>=�>�I�>A�Խ����\�����7>1�B?Y��D��u�o�z�>���?
�@�ծ?ji�R\?(*��n��+M��u�>�6Ӿ�c�>�j*?��%�F�">v?������Lы��#�>e��?7��?��o>�w?�`��5��=��=
?�g~?7�?���=�Ҿ��[>�@?N о�|��}D ���_?��@.�@�|�?(�����ο������O�/����=%y�<�)�>�X�~7A>M�=����r�e=�[�>u@?/e�>"+�>	0>���==4 y�[��!l���Y��D�B�������0`�����	�U�aT4�A�Ǿ����$���������؅e�bhS��K;���=H$R?n(T?9iq?;\�>2tn�x�>� �a��<�K$�l4Y=D��>�/1?:�I?os%?�/t=9Ϟ��e���}��:��*���>��T>~��>rg�><¬>�f���A>J�B>��>3��=6�=�<��=��D>ߦ>���>�;�>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?�f>xu>��3��d8��P�B{��;j|>*46?�鶾�F9���u�ƲH�&dݾFM>8ž>��C�_k�+���R��ui�֔{=Sx:?��?[4���᰾��u��C��%QR>�9\>hT==l�=lYM>l\c��ƽ�H�we.=���=��^>�b?K8,>�v�=A��>�2���O��j�>�tB>E�,>�@?�(%?����_��*-�� �-���v>2�>'�>��>SJ��[�=-a�>ORb>4���愽M��P�?�!xW>����Hm_��Ev��Dw=t���g>�=�L�=� �{<=���$=�~?���(䈿��e���lD?S+?X �=(�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��H��=}�>׫>�ξ�L��?��Ž7Ǣ�ɔ	�-)#�jS�?��?��/�Zʋ�<l�6>�^%?��ӾPh�>xx��Z�������u���#=Q��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?roi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?-{M>T�?�|U?�64>V��=���E¿��Z�b�=k�Q��ԝ=��G>�[<�L:4����H�~�H*z� �����>I�=崹>�"׽РѾHW&=|��L־]��=f��>*�>":w=x�4>��?jq	?�ur>#�b������:I;��K?���?���2n��O�<\��=(�^��&?�I4?�d[��Ͼ֨>�\?Z?�[?�c�>/��%>��迿$~��}��<��K>'4�>�H�>�$���FK>��Ծ�4D�p�>�ϗ>����?ھ�,��{Y��B�>e!?i��>kѮ=?� ?�"%?�q>8��>�D����;G�q�>@��>!;?�t?�,?�ڭ���/��{������c0X��@F>U9w?�8?��>�#��=���C�仮�	�CF���?6r?��~�œ?))�?3�;?'7=?��p>^\�ƾ�N�=�>��!?�	�ιA�O&������?*O?���>y$����ս��ռ��/x����?'\?�<&?��&a���¾�6�<�N#��U�~K�;+D���>��>ƌ�����=��>�ް=�=m��<6��Fg<�n�=�~�>*��=�-7��q��r�+?C�J�;0;V�&>�8`��=h��!�>�ǋ>j�{�+�C?�:��_w�ӓ���x����	à?�R�?�Ϛ?�M��5e�7�2?�J�?�J�>}�>�۾W����8¾C ���������8>ԃ�>�d���� �پ��ó��)����Z��r8����>G��>�?h�?��<>;�> Oa���1�������}�e�m��/�8�G��˖��d��E�R�t�������m��C�>�d����>0^?�J>6f>���>MO����>��>E4�>-%�>�B�>�>>!��={Ί��c��s�R?ܾ���'��꾬���^B?��c?�C�>vpW�ꄿ�&��k ?��?vi�?N�u>u/h��*��C?q�>;��!�	?��:=i��ܵw<U���w��7������>ؽ�9�U�L��$j���	?e??�y��Κ;8&ٽ��ƾ�T�=�*�?��?gn4�sH��}X�&��L�J���ҽó���O��B�����o�����ts�>E��G�5����=ʐ-?@��?C��ZS�ح�Y,h��3��c�>��>��2>�}i>�\�=�p��I�-�?�x��n:���|���>杇?��>��@?��>?g�K?٤F?��>�>�)��b�?��A;�>���>��4?�(?�!?<�?a?$�K>�#��k���]ܾ_?�Y?� ?�m?���>F���U н��<�@�`���� 뽿>ݖ<���B�#E{=X�>�*?Pb=q�1���+���>V�i?�>zُ>h��\����=���>�#?�>ό;�n�
��R��>�^�?���lD�@��=S��=��6�|���G��=��=��=|��1��=��$>*@>{}=�`�;�Fl=���Nμ�[Y=�t�>6�?���>�C�>�@��/� �e��f�=�Y>5S>y>�Eپ�}���$��v�g��]y>�w�?�z�?޻f=��=���=}���U�����G������<�??J#?)XT?_��?z�=?_j#?յ>+�jM���^�������?]!,?���>U��<�ʾ��ǉ3���?D[?�<a�����;)��¾N�Խd�>�[/�a/~����dD��慻������*��?���?^A�E�6�Ox�ڿ��\����C?"�>nX�>_�>+�)�d�g�K%��1;>���>+R?kػ>u�O?�n{?d�[?�T>8�n���֙���I��">��??�x�?ێ?��x?��>g�>�>*���������=���D����,Y=�Y>�^�>o��>�]�>�A�=�\ǽ�~��A�9G�=��b>|�>�B�>J��>v�w>���<��G?G��>�!�����`פ��L���|A�_�u?�Đ?<	,?�M=v��RvE��������>Q)�?�ū?�0*?kR���=j1ϼz��Zs�f�>w��>�c�>�=סH=4q>4Q�>%��>Z������98��6O��?F?��=�3ſ��p���i�Y����}<����/Cc�Ǜ��^�q��=�C���:�Nr��]�\��࠾���е�{O���z�D��>Ą=@�=�"�=���<��Ƽ�E�<0s>=�@�<b�=��s��6	<��.��Sq���k�8��L<��Q=��"�Ǿ:Tu?VML?*2?n@?�m>��>�$�����>@(����?�?G>�-�'r��7/C�M��o���^�чѾ�K^��w���;>Y�ռx>�3> �=�\һ�j�=�V�=���=�w?��kA=7C�=��=y��=���=f3>g�>�x?Жy�j���G�7��Oͽ8-?���>N!*>�;n�=?��>�p���Q��Ry��}?\-�?�8�?�+?�����G�>�o����=��=B��ſg;�=Pv�d��>-C>�k�7���yN��?�v�?��1?�}��vǿQ�=>�R�=(�='L�C&�6���t6�K���:?`%;��(��_ɰ>n(�����۾@�=r&K>��=q��1t�P�D=�`Ƚ���=�؄=Xȱ>P�>���=� ���.>NS�<+��=d*�>�0�<r��<<Zd=��5=d��=q�<>�>���>D�?iC0?ׇ`?|�>�q�EӾ�����ڍ>/��=v��>�h�=�H>|��>ȶ7?h4???G?/x�>���=l�>~��>TC/�t�q��j�k֡�oH<J݉? �?�O�>"='�������;�U��gc?7j2?��?�x�>�Q���B&�:���#̽��6���>ѭ��^�㼏�w=�~v����Y>���>�w�>[��>��Y>�>I�4>��>>�>�ֺהA=�y�˧B=ql=�Ԝ=��
�͠�=������u�*�_0���}�����<JƓ<:y�;��<D��=��>l�^=�]�>��=9ؾ9>$��ttY�%m;�d��mW��eq�TZ��1���s���> N}>㽊��������>e{A>�
�=/��?�A�?&�=�h;m5��⬣�0��-���g>�T;���1�I��[f�C�Y��h�����>�ڎ>f8�>D�l>�+��?�f�v=����d5����>����CQ�;���.q��/��J2	i��$�I�D?;8�����=*%~?g�I?�ɏ?O[�>F����ؾ'�/>�遾��=�+��+q�������?�'?H��>�쾞�D��m龷E���*�>T<Y�󒈿�*���5 �a������f��>SY�,3���Y���h���ZJ���h���>�H?���?�Q�u��+8p�-��4���j?��?[fM>n�>z�+?��jH��l����=�@y?���?���?</���=Z����p�>64?�?�?�?�Ds?�h!����> �=B)<>�ꔽ��>�|<>��>/�>:?x,?�G?_}���D
�)��1+㾐�H�d�
=�[=oՏ>X��>��c>�]�=�A�=]��=�?\>�͠>�G�>�7g>3S�>ཋ>>[����?�>���>
_<?���>�)>����~��ze�<��d��|��j�2x<[&�=�=�ZV=�Z��E�>پ��?�? �n>e�r?P:����J>��0>��*���>��>eّ>��>�}�>���=P�M>FQZ>��ӾR>�M��� ��kC���R�g�Ѿ~�v>�Ŝ�(�%�^	�{r���H���������i�3���C=����<\>�?�V��ybk���)�cX�(�?���>^6?�F���V���>�9�> ��>�t�����1Ӎ��9��?���?�:c>Q�>�W?�?a�1�3�puZ�`�u��(A��e�ͼ`�u፿���q�
������_?�x?�vA?ah�<�;z>*��?�%�C֏�R(�>'/��';��U<= -�>|)���`���Ӿ��þ�5�{NF>O�o?�$�?rZ?SV��C�E:2=)E?��J?�Kx?�;?�\(?E��c�3?*>��?0?@$1?K�R?�?��
>Yw�=����d�Z�d����N琽��	���=��>�G#=B���w�1��[��ʴ=M�X=�!#�`�>"'<�&��E+K<�>���=�Ʀ>ب]?{A�>k�>��7?1��v8�����83/?��:=U������Ϻ��f�>��j?���?�aZ?rd>��A�>�B�~
>CH�>x�&>�=\>�l�>7���E����=^G>�7>gإ=~�L�Kρ�0�	�3���&1�<>���>�)|>-!��o�'>�~��]Qz�X�d>��Q�#ʺ�>�S���G���1���v��R�>��K? �?�Ι=�P�;V���Jf�?.)?�]<?�IM?x�?�$�=��۾u�9���J�N�}�>�<���I¢�{"����:�f��:&�s>&?��Q:辶^> ���࿾`�K��g��/�B�=���n�3�]�$����Z�Ѿ	�!���=���G�:/��#����>?-�=�
�uu�¾׾�I>$�>���>�gϽf�g���m�r޾�k=m��>&�F>�ٳ�H��W�3�|8�Sk�>�gF?�K[?E�?�"��h�v�h E�Z���������CH?�K�>C�?D�2>
�=�{��HU���c�gfD��J�>eE�>����H�h���1w�$�2@�>�q?}
>S?�|N?��?B�a?u,?�O?��>hDԽ�g��K�%?-"�?WK�=U3ڽN�i,9�4G���>f_'?�P�k��>�?�?̜%?פO?�:?og>yo����?�귔>N�>��V�c-����Z>'J?�T�>�Y?�?��<>i�5�9���y٫�:��=W+>�2?*1$?��?rƸ> &�>)֢�u|�=�"�>D�c?Lރ?��o?J�=��?�4>���>2h�=���>���>I?��M?j�r?��K?JB�>�K�<�g���e��ؿk��S���ĥ:r�)�l=Ò �և��3���<��;w�ԼB��������$�=x�2�J<q��>}�9>o�����>�G����f��w>�#�����`�}��猾v�V>�v�>:N	?�,�>Kܽoh>9@�>�*�>JX"�Z�J?e�>Λ-?�z�=��q�#��ф3�QŊ>3�&?�o��̅��ڍ�H�{��g=�R?�m??�9��o�Ҿ_�T?$[d?�[�[��Ⱦ�NvT��I��jx?�?�#���=�>I*r?��O?Ԃ�>Vt�
/e�jT���[g��^��R�>K}�>%Y� ��X��>�V?~t�>��>���=�⸾�Kn�'���jR?k��?�j�?92�?H��=��d��V޿MS �,!����[?�\�>X}���"$?�����Ӿ���������۾�����p���]��Pȯ�����,���@��=�?�s?�t?�^?ϛ��]8Y�
�b���i���R��6� )���N���C��MB��	b�x�3�������>w�U>��Gr7�IG�?VR&?D�-%�>� ������
ܾ��<>�k¾U|P�8Q}=D�ֽ�ܕ<ܺ�<HG���T�%���*?"��>��>8;?�;U��	<��f,�Ԅ5�E����D>jr�>�@�>6t�>㦁��9J�^�ѽ����&�K����1v>�{c?sYK?��n?K-��S1�����3�!�..�U���LC>��>��>	 X����4m&��S>���r�L�� <����	��@~=qk2?��>���>]4�?�3?V	�G���.x��{1�U�<|p�>�(i?�^�>�>Wѽ�� �$��>dkr?���>�}?{�ͽ��P�4Kq�֒�=��>b�>�# ?G��>��3��aj�󮐿朑��' �D>k�n?�0��:��[j>N.N?'h�=H ��	�>����"N��%־��p�g�>��?�x�=�=����y�������K)?sN?�ݒ���*�I~>g"?n�>j?�>�/�?�3�>�_þurA���?d�^?(FJ?+NA?9�>+U=Ј��\dȽ �&�e(-=���>��Z>��l=���=3��hj\��X�T"E=+W�=�)ϼ�o���~<�ǵ�V�M<C��<t 4>�ڿ,I�jEվ��Kr�5��B�oaǽ;���O������k@����*�NC���S��]f�����n�L��?���?��������$��w�|�����zp�>�"v���������P���꙾�(�����!�]xR�X�h�-h�M�'?�����ǿ𰡿�:ܾ6! ?�A ?6�y?��4�"���8�� >TC�<&-����뾬����οC�����^?���>��/��n��>ݥ�>�X>�Hq>����螾�1�<��?6�-?��>Ǝr�0�ɿa����¤<���?0�@��A?��)����t	P=��>^K?&%I>w5����e��)��>�;�?-��?9"z=��V�i��xXc?+�<��E�w���:��= m�=M]
=?o��6K>�n�>dz�B�7ݽ�c3>0��>�(�8���}b�b��<\�`>��˽J̙�5Մ?.{\��f���/��T��U>��T?�*�>k:�=��,?X7H�`}Ͽ�\��*a?�0�?���?$�(?9ۿ��ؚ>��ܾ��M?]D6?���>�d&��t���=�6���������&V����=g��>x�>ɂ,�����O�>I��O��=�*���L��$���'��b�<���<�o����K�~��������G���m��&����<BNW=��P>בm>��=��N>ǷT?kp?�9�>8^>i�X�{5p�[��u[�<���48f���оzFu�r���a �l/ݾ�
��*�x����-%=�}�=m+R�۔��f� ���b�8�F���.?cf$>8�ʾ��M�6,<L|ʾZƪ�y���諒25̾�1�
"n�˟?q�A?&��V�b����I���³W?@a�տ�����D�=l3���Y=% �>O�=��� 3���S�4�.?=�?�6��]����P1>��	�#��<_w,?a#?�|�<^ʬ>ؼ"?C�0� ��A%o>�3>I��>���>���=�ձ�L�ͽH�?O�U?'����X��M3�>F�ʾܹz���o=`!>'�.�p��0`P>���;(#��=�0;�̐�;�L=�#W?x��>U�)�����X��Q����<=Ͷx?�?Z-�>�{k?��B?w"�<|u��"�S���
pw=�W?�+i?��>Wq��3оe��K�5?|�e?��N>Mzh�M��@�.��G�U+?r�n?�[?,̝��|}�������7f6?��v?s^�vs�����I�V�e=�>�[�>���>��9��k�>�>?�#��G������{Y4�&Þ?��@���?��;<��V��=�;?i\�>	�O��>ƾ�z������F�q=�"�>���|ev����R,�c�8?ڠ�?���>���������=�ٕ��X�?2�?�d���|k<���l��k��A�<�x�=u��Z�!������7���ƾ(�
�{��Y������>�W@|~�z0�>?d8��6��[Ͽ���D_о2�q��?�Y�>;�Ƚ�����j�w3u�+�G���H�%����j�>�~�<Dı��u¾=���+oS��6a=���>�$�=�}?�]�8tҾ=챾�*�	l�>��?@ �>s��:~K�V��?%���ܿnk��e��{K?�m�?A�{?�e?�OE>_~�M�C�����Pxi?g��?=o?]H�=g+����$���j?�_���R`�8�4��EE��U>e"3?QA�>̓-��|=8>��>Qk>%"/�ݍĿ�ض�i���s��?T��?�n꾨��>���?Ds+?j�8��b����*�!T-��9A?<
2>ߎ���!�0=�uђ���
?�~0?Rs�C-�)6p?�7���p��UzK��!���l�>�g�=���C�>���=q�E�*X���f��\��?2�@�շ?��F��$��9D?Ai�>�wԾݖ�����=�"?�"�>r.�>�k+�p��=i�U�2�-�h��>���?O;@��?�N��Z�����>3�\?P+�>9f�?&�=!��>h0>�L����9��)>2w>�[u��?�H?5@�>�ͼ=�����)���?�ӳS�t���;C����>e�b?��M?
w`>NG����P�)�%A۽�S1����;EH)��_"�$G��L�>��+>��.>��A�d�����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�b��=��7?�0� �z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�Q�B�{�1=6M�>͜k?�s?!Qo���l�B>��?"������L��f?�
@u@a�^?*��׿���5½�0-���_B>=�n>>��x��Ӳ=#�!>�Л=Q�=�_F\=�$�>j!>�uK>R�u>��>�D+>+q~���Q���ʺ��� B�V+�O��57��6��
:�������������D��Tֽ�,ҽ�����r�M�=SLX?,�J?d�e?$�?�h��J�.>�9��=0����"
>�a�>XQ?�4>?cm.?�Z=�R����c���{�US��f<�����>��]>1G�>���>/e�>����J%,>�>m��>>~*>X�@=�Q���ɏ��r2><�>�X�>R��>�C<>ܑ>;ϴ��1��]�h��
w��̽9�?d���Q�J��1���9��̦���h�=Qb.?|>���?пj����2H? ���m)�$�+���>v�0?�cW?�>��1�T��9>U����j�4`>�+ �<l���)��%Q>_l?V�Y>��v>��,�H6�|�O�h��8�{>o�5?ˉ��;�+sw�xJ�.�ྀA>�%�>���V�!��H�����;�b�Fww=~�8?I�?�⼽�[��(�d�d���q�L>�f>0<=�}�=�8T>��n�
ν�.D�56=��=@o>ȋ?��.>&R=Q�>Mؗ���U��˪>�Y2>�>�9>?,�?S)��{�1C~�6"+��Ym>�O�>1��>x�=!+Q�~��=��>�i>+(F�bl� �
���4���G>�+^��WN��⚽?u=j#���_�=׍s=6K�4+C�3�=���?�o���L����[����H?l4?�)-�n.���5�N𕿇l��J��?�@ë�?�d�wQA��t"?ET�?74��Η�=s��>+۩>޾�6{�j!�> X����#���佼_�?Tٲ?ed��Xo���w���=9%@?'l�Ph�>{x��Z�������u�y�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?L:>��?��Y?�R?�o��(lS�*���c��V��=Wi�<��>J>�Ǿ��P���������`����h>`��=L�>�a콋@���	g<��J����)���c��>�+>�C>��{>E��>��>_z�>)=řϽ����o��+�7?��?���aPm��Y�=c>�=�����mN?@K?��f=`�?��>O{+?	~Y?�z�?N��>�������7Iοa緾�ā<X�>]�>|��>M}(�	=�>���-
����>��g>�I��'vྈr���<�L�>��*?�>�K�=�?��+?g>>|��>��6������3Q����>���>��>,G�?�7?�lȾ2�5�o���#���Y��C>�rg?�)?}�>�9��LW������4�=����7�?a_?�68�%?aw?.U6?�4N?`��>l#����n ��j/>a�!?
��(�A��m&��E�Ǧ?�?0
�>�!��z_׽�ʼ�q�����[�?J�\?%/&?����Ha���ľ�=�<�z&�*�'��0�;*�'���>i�>������=Ԓ>�ȭ=3=n��#6��2j<�:�=*+�>P�=-�6������;,?`�F��݃�9�=��r�ixD���>�dL>����ڪ^?va=���{�h���x��U� ��?#��?�k�?�ڴ���h�b#=?��??�'�>*S��x޾���Uw�!vx��l�%�>���>2Am��徴���k����F���ƽf�
����>Å�>�'?$��>�|L>�>������4�l�ɾ����S�y����!����\��%����Y!��8�La���������>�墽�9�>��?j�>�t�>��>#p�=S۩>j�'>��y>��>+y3>��>�XV=q8�G�m���e?e��g����s��{�Y?C��?��D>��1�q�z���R�i?'1�?���?(L+>�+I���
/	?�g�>,+���#H?N�{=##������>D�lKU�?vԽAA&=�в>8�'���/���s���¾��?��?	��=�R��L�����T�=���?.?G�+��q)�mI���@���p����RLʾ�(����x��a����|�-w����,�v6�=�0?#�b?y�ܾ|�Ծ����Pb�ƝL�Ί>k.�>�ߋ>�;�>w�]>5־R&���W��x�ӈ��U?�p~?Mv�>�[N?��=?�GL?��J?��>y,�>� ���| ?	�=���>���>��-?VH$?�2?��?��(?��,>����%D˾��?��?�?�?��?�/���o۽�.�7�=LyP�
�E�j�'=��2��ܽ�����==*1�>�U?Y[���8��`���k>,c7?���>���>�H��H�����<
��>
�
?�Q�>����dwr�Z��_�>텂?��i�=u�)>b��=��~�U#��v��=ʾ�~;�=����8��<�M�=+W�=�}u��P�X�:��p;#}�<��>-�%?�:N>�$.>G=��L ޾w9%���>�˔>�P>A�=Ř�T���Hk���o��:�>Mu�?��?N�>��=�#>�Գ��E��ܾm�CN`=��?Lc�>�mR?��?W7N?z�?�-S��u�S����-���~���
?[,?5��>����ʾ+��3�ҝ?�Z?r<a����%=)��¾��Խ��>F[/��.~�����D��?��I��;���%��?���?�A���6�Cw�y����]��@�C?W"�>YX�>#�>��)��g��$��1;>���>�R?4#�>��O?�4{?ۢ[?�vT>F�8��0��Wҙ�a�4�R�!>�@?���?��?'y?o�>��>פ)��ྐྵV���������䂾��V=k�Y>���>�!�>%�>	��=XȽ Z�� ?�U�=`b>΅�>���>��>�nw>X%�<6�@?�U�>uG�������7������g?�ދ?ћ?��
��<�;����ଔ>JN�?@�?Z~9?*�݉�=M��������9��5��>`=�>S4�>ݏ+>*E�=N�V> ��>z?�>cGR�r���*;�򫰽s�?�kC?0>����]����S���\伝�J�PD�Pg0�퐂��d=��;��x��F���݄�a(����������9¾c^����>J.h=�v�=�� >�2c���3����=���<h"����=}y��)��;�S�<�ﰼ(��U-<8D<eP�=�*�=��ľek�?�qf?�3?ՄW?`�>��]>k̽���>`v|�3bK?���>�½�¾o��s���� ��w
����3ၾ�+����2>6ha=�̍>��>���=����=K����)>j�z=��\=���=}�%=t&>���=q�>��>�ww?�偿򈝿�DR�)1�V18?-��>���=-����C?�=>����y���i�%R�?���?���?x?R�_�F��>�(�������b�=OȄ�Z:>.v�=7�2��V�>�G>W�������h^�?$�@Ň??=F����ο�[0>#=8>��>9�R���0� �[��c�1(Z��� ?[;�e3̾�Q�> �=�޾��žrn-=�v6>wlc=B���>\�cY�=�z�G�;=�nj=|�>��D>lŻ=����U��= L=�>�="N>���6���.���/=eM�=�`>Q�%>��>�?'(?��U?1��>n���b���lþܠy>�@�<氛>	=��G>�I�>��,?�Q?�O?��>_�O=X��>?c�>�I)���n�M�羕L��c��<S�?�X�?���>����9�N������:���	�oc?#7?^�?��>���c
ҿ�H*�v�A�k%����P;$=�@���Ww���=�����ߨ�E����>⭗>m^�>z��>$�>s>�v�>� 5>?U��My���G���\�=ր�_�<�䒽#[<�ȁ=&���E�J�g�*���H�=6�P���A �;�z>c�>9��=ߜ�>o�=������9>�m��hJM�FC�=�"����:���T��7s�۫)�˩B��;>�n>����ӏ��9 ?_�R>��K>!j�?�?r?��%>�$ݽ1�޾"t��Ɵ2�	o�N��=�c>�.>�_�<��ca���O���о���>X�><�>��l>�,��!?��"x=y��c5�y�>=��������-q�-:����?
i��º)�D?:D��"��=�~?�I?9�?q��>7����pؾ�0>9����=��"q�cZ���?�'?u|�>� �۾D������Kнg�?�= ��b��܈�B�1�Ge���|�7��>�(ž�� �#��ۈ��m����0��y���ʢ>�Q?��?�&��3\����_���>��o��Y�>j�Y?u?��?P�?8L<���s���u>B�u?`�?ǅ�?��->��>��{��>?D�>��?�M�?�v?��1���>,v=e��=� ���U(>�33>U�=V�= �?
&?t�?��������ᶾt�K���%�<-����{>��>��>� �<ܔ�<��=w�#>�m}>u�>�S�>��>��>c�j��D��V?�>E��>�e;?Q�>'
=�9�:�>��q���uۑ�퍭<��k$g�#`��[�=���]
�>�nĿsâ?��X=��ʾ]�+?�Ͼt��<u]�>)�:>K����>�\7>�Yd>��~>��>��I>��>���>�,־��>���H�eC�t�M��h˾Yjy>�����w$�]'�t��X�L�	2���j��i�N����>��H�<~n�?�� �çh�>�%�p����?Ш>gl2?�Ő��1g�l8>�/�>��>#����0��� ���޾��?���?N	�>ϣ�>�C?.�	?�?��o�l�cao���F��q��R�a�����L�vӾ!ݛ��Fw?�r?bTb?=5;�Q8'>��?)2�/<��t">kWI�imN���<4�><|��;��N���ƾ�PL�R�9>Iy?�n?�3�>[���dNu�->%<?A=2?Vu?�2?�@;?�9�X]%?+g3>��?��?k�3?mc-?F
?B3>���=q�I�ʺ-=Tʔ�?"��B�Ͻ�I½p￼h�7=Es=����V�;=���<rL��Ҽǯ�;K0��揾<��3=�s�=Q��=ʩ>b�X?;L�>/>��/?f"���D�ɇ���*?gi��2{���,��u➾����=tT?d��?��h?;cp>�9)�m7$��>�fQ>�׎=I>��>�_�<�Ž��>�L�=��=a������L��]	�?�H�T{�=M�v>ް�>�D|>���rM>�u�������Su>������C��%L�ы!���B��n�> �C?��?�Ϊ= ��������e���.?>�,?D�T? ��?��e=�޾��*��\J�\��[]�>����Xe��n��� =���1��ei>����ܾ g>�״�(f޾��x�G�5���Ҿ?�F=Ί�jM�u7�ٷ�����<���=���=�|�������KG?pr�=88l�_�G�tо���=q��>$��>I���?ʼ{C�:���(^=%��>3��=s��|F�"�K�����A<�>XE?Z+_?={�?k��Vs���B�w����)��Ȑ̼��?�w�>�8?%�A>P��=౾���d�OG���>�q�>����G�5q�����$�?Ҋ>v??M>ļ?��R?�
?��`?-*?�@?��>���Ѹ��C%?��?K�W=���/�?�:��K���>��?�FR����>g�?�?�(?�0[?�b?�`>�����3�-/�>�}�> �R�����v�f>�M?�ͷ>j�^?�U�?�lU>D�1��V���mҽLÌ=0�>��0?f�#?�?o�>N��>����D�=��>`?o�?��n?,W�=�s�>L�.>(�>��=�:�>��>\*?�6M?�{s?B�M?5��>�^�<=D���w�������a����T���3=|a	�l�̽D���|�<�[ <�E߹j2�5O�����5'9�.|<`��>�^>��׾Q!9>�`������(�>�P����徟�˾� ���^!>�^�>H?%�>���X�=p	?�ͪ>K#��w/?�P�>̘?�mU>�\����2��j� Q�=�,?:�$>�Cw�U����`�OM3>6I?� "?n\��h�ƾ�W?�f\?�㾭}(�s@��[!g�ЍǾ��x?��/?̾��>�ym?��>?$�>���Q]h�

���G~�}�ž	,>{)9>��Ӿղ���9�>�*?W�>�s�>�b�=�|���.���/¾�p"?�u�?pX�?Q0�?+�=d)\����L���鑿k^?��>�
��X�"?7�.о�Ջ�H鏾�⾝��æ��Я��@ԥ��&��#��S���,�=�e?Rot?��q?h�^?_Z��xc���\�mx~��U��g�+���E�fE�InC�O�n�������M��n_6=ؕ}��,A��$�?��&?�@1���>�k�����RTξ��?>�Ġ�z�A��=\���%A=L�^=�f�i�*���m�?�9�>��>�=?[�2�>��g2�#,8�F��>10>\ܡ>Y��>;�>�\+;4�(�vs��
ɾ�m����ҽs�u>�c?��J?�Uo?������1��l��q�!��*��z����D>��
>wy�>Z����k�&�rF>��nr���F)��R�	�'�=�2?��>���>��?�r?��X-���w��1���s<��>^�h?��>�ԅ>}Ͻ�� ��I�>�~?�|/>�T ?�- =~]�V�w��܍�B��>���>b�?\Lj> 	��t~�����{m��6�e��=��C?W)��Ƒ��0�B>@�Y?���gtZ�%a�>����� ���>�����>�1�=�7'>/��b�0��x[��.��WK)?a@?�ᒾ�*�S1~>"?8z�>��>]#�?�(�>�eþ�y2�A�?��^?�2J?�JA?8L�>̍=�ﱽ�DȽ/�&�NE-=a��>>�Z>r�l=g-�=#���u\�J��N$D=�w�=]μ����P<Pd���#N<E��<�4>_fܿ#[B��͔����X���W�È��������V�;���̾l񶾄����8�b����~��2���Կ��Vl�B��?�K�?��սc�v�7,���n��-ʾ�W�>\�a�hy���+^�]
��+�x�þW�/���k����\Oi�@�'?����޽ǿ찡��:ܾ+! ?�A ?1�y?��4�"���8�� >2C�<7.����뾮����οL�����^?���>��/��n��>襂>�X>�Hq>����螾�1�<��?6�-?��>َr�+�ɿ\����¤<���?.�@-�@?/-���v륻̘�>r�?�V_>��B���Tڪ��c�>EÞ?�׈?%I�=�R��˦��Nc?Rk=�8��a::�i>���=ҽw< bN��X6>���>�2��=�g�&�[�=�Њ>�<�a^���L�K�c=j�s>JT���]��7Մ?5{\��f���/��T��'U>��T?�*�>�:�=��,?V7H�\}Ͽ�\��*a?�0�?���?�(?Cۿ��ؚ>��ܾ��M?VD6?���>�d&��t�Å�=_7�|�������&V����=���>��>ʂ,���ÇO�EH��u��=�{�Y&ſ���t�8<?Խ<����;!�ȝٽ@,O�����z��ٽ#$=d9>K�@>��>o�W>c>E^Z?�y?"�>�{>�,��[��Ӣ����ּ	���[B��Ǻ���3�����i����N־����(���$�$Ӿ�!=���=�1R�떐��� ���b�|�F��.?Jt$>��ʾ4�M��-<�sʾ�����������{3̾�1�x!n��̟?7�A?!�����V�O �]�4x��!�W?�O�����מּk��=����ڢ=� �>E��=���z#3��~S���)?8%?;��u����Z)>7?��:=�a8?{	?ʨ�=z�>�R?��D��~��>>ֆ'>H՚>:�>C�	=ݺ�j0���%?�{[?%ỽ������>������t���>�>eg������3>�~��Us����=�����>�W?�ڍ>��)�_���쏾i����7=o�x?�?t��>�Mk?[C? A�<������S�z&�Noz=��W?_i?=0>�h��FUо6�����5?m,e?��O>��h����;�.������?M�n?� ?�K��Ğ}�*0����ށ6?��v?dr^�Js�����p�V��=�>�Z�>U��>t�9�4l�>Q�>?N#��G��ۺ���Y4�HÞ?��@X��?n�;<{���=�;?s\�>�O��>ƾ��������q=u#�>����dv����bS,� �8?y��?���>����������=�֕��V�?�?����d�f< ���l�cv���m�<���=V���"�����7���ƾ��
�7����Ŀ����>Y@7r��4�>I68�&8��UϿ����_оfkq�t�?�z�>n�Ƚ摣���j�^Eu�D�G�%�H�դ��Է>��d��ԙ;��7� &#L�zN=���>f�n<��?D���ҧ�������ɽ0
�>�?�g�>N��*�C�(.�?\�*����R$��Qm*�6sb?:׿?��t?w#y?�K&>�m���Y,���,��$i?fم?�Qx?���<�\�.y��j?�`��U`�C�4�"HE��U>#3?QA�>��-���|=�>���>{i>K"/��Ŀ�ض�����Z��?���?o���>+��?s+?Hj��7��_\����*�H,�R;A?�2>������!�l/=�[ђ��
?8~0?�y�@.��p?0�����-�/�Z�F�<+�>��<4Q��.O�=�ˆ=kU�X�������D�?�" @���?�=� �7��� ?��>`����1M�<�b?D��>i�(>��7�ݧ�=dE;��B.���Y>���?BU @���>����䦿��>Yn?ޣ�>�܄?T��=S��>[��=�m���w��y9>gY>�q��??gLC?�D�>�O�=>t<��,��A�M�X�
�A��#�>�4a?JM?��^>�Vн�5���!�̗ѽm����ݪ:�!j.��(��H$>T�3>Â+>�<��O����?Np�9�ؿ j��%p'��54?2��>�?����t�����;_?Uz�>�6� ,���%���B�`��?�G�?=�?��׾�R̼�>9�>�I�>D�Խ����\�����7>1�B?Q��D��u�o�w�>���?
�@�ծ?ki��	?���P��?a~����7����=��7?�0�W�z>���>`�=�nv�߻��V�s����>�B�?�{�?.��>*�l?��o�S�B���1=M�>��k?�s?iAo�O󾞲B>��?!�������K��f?�
@u@T�^?'MW޿6p��S������[{�=UA>�;>���S�=x���
=8(���>��>�q�>p�>*�`>�}�=�*�>����5��,��y?����2�E��5��遾!��T���=�1N���
��%����r<? �ý>���a=V��=N�U?cR?>�o?7� ?r#y�(�>�b��V=�3#��ȅ=3�>,W2?�L?>�*?(Ó=�����d�bZ���G��(Ǉ�l��>�I>��>�U�>s�>�)�8شI>`?>�~�>�� >��'=0�ʺ�=��N>�K�>���>뀺>1H<>ʖ>�ʹ�2����h�
w�̽C�?�y��o�J�)0���7������n�=�`.?�y>��?пk���G1H?~����'��+�0�>:�0?�bW?ߝ>���,�T��6>
����j��b>�$ �Xrl��)��)Q>g?ŏg>I�z>�1�tg:���N��5����z>�7?簾�_4�7q��TH�3;޾�CF>?�>�hd��y��.��ײ����k���=}�:?)T?���GŰ�`�q��C���dK>L�j>�z5=��=��J>����ͽ��D�%e=���=��m>�?\ZD>ݝ`=2��>r�����d��,�>�;>�G&>t?? [%?��=���W�~��)���h>�\�>���>h�=:8X�\^�=��>�Xx>ك;���,����7�Q�>>ƕ��F��CA�2�=�w�/�=��=�<��i�?����=;ފ?I��'j����ҾQ�O�Z^L?GS?� �.����������挽�[�?Cx
@�x�?k��#}A��?��?���E�">�?{�>n6 �����>R�������wh(����?1|�?g��Ab���>}���>5?C?3���$h�>�x�kZ�������u�j�#==��>�8H?�V����O��>��v
?�?�^�ᩤ���ȿH|v����>R�?���?^�m��A���@����>3��?ogY?oi>�g۾�_Z����>̻@?�R?��>�9�W�'���?߶?ׯ�?��?>
��?��W?2X
?�����K�%&���n����=��9�O[�>���=��پh�P�2W���ɏ��g� 
�M�>�H=��>��ʽkj���2<Ea�G�����n��y�>FC>�E>�M�>���>(
�>�.�>Žƻ�ֽ�Pp��B{�bOE?�ц?6���t��V�����R�$���6?':G?���+�{�u�E>c�0?��Z?��=?Sw>z"�p��5wؿ򳱾�o=��h>lJ�>��?�����>S��b܃���>&D�>v��9kᾨ,����I�	��>,?�?S��=�?@/?��>�3?X�0�ވ���~;���>� ?�_�>�΂?�@?c<��t?�B���W#���Y��X>�FY?�x?��R>�Bz����K_��n�=@g��ؓ?N�j?�#�,��>�b�?��6?�P? \I>��Y�f#̾E@m���[>��!?x�T�A���&�`���>?�5?	C�>����+�ֽV(Ӽ���T����?�\?�!&?���a�n�þ�=�<�N!��9A��5�;��8�6>�Q>�V���x�=�>���=W�m�.�6�-�\<�;�=X��> :�=!M6����=,?�G��ۃ�{�=��r��wD�J�>%OL>F��>�^?�l=� �{�����x���U�N �?��?-k�?s���̝h��$=?�?
?U"�>M���{޾���^Pw��x�<t�t�>}��>)�l��徏�������F����Ž�:��W�>��>S.?�P�>�->���>���K�%�������%GY������5���*�9������
��V9�8뻾
B��s�>�߇��4�>H�?�uW>��{>wN�>y-�;���>;LS>h�k>���>�TJ>5g+>��>i�>�ʽ�t`?����N'����6�	��]?L~?L�w;� H���j�L�O!�?���?��?Ϥ->��(�f5ܾtZ'?rn�>����MW`?	=�;��>�/>/M��	Ӿ��7� ŵ�P�=Ǆ���EQ�F�S�������+?S�?>��� ��nR���8۾af�<�Ə?��?��F�}�9�Z!B���,�H�h��ª��ž���	���Et�K����������h4�M�=a)?��N?02վ`<���(�g�4�t=�d��=�w>1�>Kа>��{>�r��Y|1��C�zL	������-?�{�?ͅ�>$�I?��<?�RO?�J?ұ�>�>�ާ�Wa�>,�<Ĕ�>ʢ�>A�7?�,? <-?]�?�%+?��`>���6���վ�[?j ?.?<�?�/ ?Wֈ�cw��W�
��_ܻ�y�V�i����=��<|�ڽ0 ���X=�P>%;?�����7�Z���0)k>o�7?r��>���>[��rm��jM�<���>�f
?.H�>�����p��
�~��>�P�?:�p=	,>Ҳ�=�׷��w���˽=b~׼�4�=�ȶ�(4Z�o�"<�_�=֎�=�/�`�s;TZ�;�Z�;�V�<m�?��&?��=>�[>U�.��/¾P�S�.�>/e�>���>�H)�m�W� z������ k���P�>S�?�ͭ?yK�=wX�=�>�M��3�O���ؾ5����o;te�>��?Y�-?���?2?��?�ļҷҾ3���֍��/X���<?',?���>�����ʾF먿��3���?d?�*a�˪��+)�~�¾Vս��>XU/��&~����D�3Đ� ��V�����?���?��@�Z�6��o�/����^��ϝC?�-�>?T�>Y	�>��)��g�O��e;>ϊ�>+R?�ʿ>1G?g^c?̜L?��>�BJ�룰�=��d���I=n2%?M�~?>��?���?_�?Sr>g�L����ʾ�;�$�������a<撟>^ʄ>�T�>���>��!=�F�V��|!��|`=�>͎�>�M�>sſ>�W>�S�=�=?�5�>�o��wP/�����>��*7�2�n?�/g?]�&?�M�&�ﾎ#Q�����
ܫ>�G�?���?��4?�����\>@)$;�	��(��h�c>�'�>���=O�>F_�>���>��v>���>�ꆾZ�6�I���ý�|5?֊4?� ��/ÿZ\��w��њ��h˽����`:G��jj��w��F�=����뀾uϼ�GZ������-w��a��4���>C��J��>bG�<u >̙�=�؆�&_��-W=��=\j����=p�!:<��r;謨�R�P���+���.Ӻ=�1M=�U��Q&u?��Y??7�7?��e>��<>fv>�D?D}���_?$�����<�^�yC��h��{������1�{8��n���:#>P	>�<W>�õ>RD�=σ&���=����'>���b�=�(>&�=�� =|�</�>#g�=�b|?K·�����VcN�7mk�9?(�>��=����Q^?�>�͂�� ��eB��h�?��?��?%��>iPD�X�>�¾�q�VZ<G���{8�>��>����#��>�S&>�����\����޽e��?c@Z�4?������ʿ�/>(�8>D>TS��L0�'\��d�"�Y�W�?g�:�Y�ʾXɆ>Z��=t�ܾ�ž�s1=�&4>D�X=S���\�F<�=>���g%L=��o="Ì>��@>���=�}��\�=�i=6O�=SDN>��Ի�O<���4��1=(��=��^>�	&>���>]�?�� ?��?{�?�;��)y���̾n�H*��>��)>��6>���>6��??vi?v=??�>\�>�ڛ>A�>����Qh�1��k���6�>�?�{�?���>?��;|�j�,%1��__���;�g�?�C4?�@�>蛉>�E�|Qݿ�]���$��fG��j�<��E�6v��w휽wջ��ݽ������=hK�>�>_{�>��>y�L>��>�9�>aY>�ݡ=� 5=䠃�G��<N����=��ۼ�� =8�!�#h�<Ӓ��`w��{	�<��.�=W}�s�����u����=��>r>���>/��=��� />���Q�L��ڿ=�7���"B��-d��F~��/�zi6���B>�EX>�P��^1����?�Y>r�?>��??.u?��>�?�a�վoM���e��eS��ڸ=��>�<��y;��Y`���M���Ҿ���>�ߎ>���>�l>�,�|?�ryw=�⾸c5�Y�>�z��W��@ ��:q��=������,i�a�ɺ��D?IA�����=�~?8�I?�?�{�>�6��ɒؾ�'0>;���V=.�.q��~����?p'?U��>�쾾�D�:ԾjK��??�<���C���{�r�=��#�����rG�>O��|���f� l��������:��;��F~�>z�q?�C�?����\��]�xd�Tv���>��F?���>>!0?uj�>������.���R>���?`��?��?}[�=z��=��ý�.�>�j?�Y�?�b�?�r?�aB��#�>���;Mm>��DM�=��>�i�=�	�=�G?0V?<�
?�I��;T	�Ϛ�����\Gf��t	=>�=!��>�߈>Z,f>1�='�u=C�=r?b>��>��>yk>F�>b�>1n^���
����>�L�=1A�>J�!?F�|>�߽F�z���=G��UŽ3����,>=�h���J<(ۧ<��>��y�C��>�gſyW�?[	��Ƚ��� ?�����4�=M+=>�>>�A��4��>���=<�>W�w>Uʾ>�z>qZx>��>d��S{>���+����M��QM��!��u�z>޵���@,�M�8 =�XbT� x¾.B�?o�K6��(mK�L�<t�?��]�)���"۽'a�>���>��+?����U9\��>#��>=4�>`1��"���������پz��?9��?dFf>J��> �U?E^?�3���5�ӐY��w�4#B�6[f�La�P�������7����)`?p�x?�bB?���<�w>+��?�&��\�����>@�2�8O>���=\�>������_���Ҿ����G���U>}�o?�9�?�h?
�T�V���>-H?�S;?��y?�f^?l�$?˲���;?��<YGR?�]�>e?�?�b�>Sk�=ٺ�=��S����2�'��^��_	�>zt�y�}�meY=xx�=�f�Wnj���.;�Dϼ�d=S�;��;�<3�o<?�=�<4r>��>��[?���>j[|>C:?4�)�b^=�ҭ���&?:;=���2H���1��=#�ml>=n?�R�?9�Y?��k>y�>���:�3L>V �>Xf3>��[>Z��>>:��G>����=_�>0$>Xڋ=+`��	����^	�G���<��(>��>z1|>�T���(>P���${���b>��V�E���VV�~G�31���r�?�>�L?`�?)t�=jc�^u�e�M�(?�\;?d�L?��?$A�=��ݾ<9���J��V�K��>˒�<���p��jh��9:��[:o�p>������̾� >��о�"��p$j��27��վ��O=����͖�2|��, �����v=5�_=��׾�f*�����ͫ��}L?k	>��_�K�Z��+ξɆ�=AѪ>�N�>+e-��i�JkJ�L˲��#=�V�>�<>!F�������O��X���>��D?"5`?r��?0~�[�n��C����,�������9?~.�>eY?��*>���=_9��]^��c�6�B����>�~�>����%E��m���,�R�%�N��>�
?�5>��?ʢQ?�_?�_?�)?�z?\(�>f੽����2j%?9/�?PyD=�Aݽj�(���<��;E�#��>b�?wpo��e�><�?��?_a+?z�Z??�� >���1��.�>���>��U�Y뮿ko>7]E?�T�>'�U?6�?we!>�D0�؏�����f='L>s�0?m�?�i?�O�>���>�����=ן�>Rc?�:�?��o?��=�?"2>���>p��=殟>ˑ�>,�?�;O?��s?��J?B��>?#�<c��x�����s�JQ��s;{�C<i2y=�%��qt�j��4{�<��;k����~�b��̭B�ʿ����;��>P�b>�v����H>a�|���4�>���Q���@*��˭��%@>rS�>��?g�>��Ͻ��>�R ?x��>?�6�T�q?=��>'�?��
>��s�Z��#�<�ш>3?W �:���wȑ�� Y���=>�`?�JD?�Si��p�c�Z?�g?����sgn�Fd%�[}�9�Ӿ8Uy?|?���&�>�p?{�$?�>&�g���y� ���W���S�ӻ���>���^�v�#�>k�+?���>� > Ƈ<�����t�~��0S?��?/U�?9��?/��=�)����n���<���]?	X�>[즾!�"?����=оV0���ԏ�aAᾹ����(���V���k��%�����cNٽ�[�=�K?ts?(}q?�w_?x�o�c�/�]�ѳ~��yV�CN�ɕ���E�l0E�ZC���n�5��z������f:=�^��KA�3��?��'?K�0�`��>����}��-';u/C>:���{���=]捽�l;=�yU=kyi�6�/�s���i ?y �>d�>�<?��[���=���1�Ȣ7�=�����4>+#�>���>��>*�:zG-�� ��ɾN#��G�Ͻ�+v>�tc?��K?��n?�S�E"1��}���m!�?�0��0��؛B>��>u��>�QX�>4�7T&�=>���r�.���o��(�	���=�2?�*�>VŜ>�6�?s�?�n	�c7��
�x�>\1��!�<Z�>oi?S�>���>�.н� ���>�ji?�z�>�4�>`lr���$�;�h���-<��>%{�>Wq�>>E\>"8o���q��������f��]=�??�+���*����>:(?@=5r=���>IC	�.B�@�ؾ6 .�Fm>���>�/=R�>���?���k��t��\&)?q�?ڿ��+*�z��>��?R �>��>���?8��>g�þל;��?�~_?9L?�C?�,�>* #=���˽��%��=kW�>�_>�q=o��=!����X�)d"�H�?=��=��ԼiYͽ��<Mح���b<�~�<c4>V�ؿ�K�m���V��)$�EX��q���^��؜����Y�S��.���^^���I'�����o|���w�ؤ��я���?B0�?c*���l������l��i־�?�>2����r��]�ZlK�"���TYվ�����u)��N�u��6t�O�'?�����ǿ򰡿�:ܾ5! ?�A ?7�y?��6�"���8�� >LC�<-����뾭����οB�����^?���>��/��o��>ݥ�>�X>�Hq>����螾�1�<��?7�-?��>ǎr�1�ɿc����¤<���?0�@{�E?��1��B��ߎ�<���>�$?���>W�H����$��l�>?J&�?��>SpZ��W����Z?��=ϱB�e�����=T��=��Y�2�o��E>�F�>vU���$�37�� j>Z>!���n����i�)p;=�4x>����	�5Մ?*{\��f���/��T���T>��T?�*�>F:�=��,?Y7H�_}Ͽ�\��*a?�0�?���?%�(?6ۿ��ؚ>��ܾ��M?]D6?���>�d&��t�څ�=6�q���}���&V����=\��>b�>��,�ދ���O��I��W��=�� �@4ÿKi��v�S�='qJ�d���b$,��@������-��o��.���b.=ͭ�=o�C>�l>��5>��G>�5Z?�^g?��>��%>H^�D፾��¾���=�����@��ͣ�`�@�����o�	�L)�*��d��ྪ"=����=�0R�;����� ���b�W�F���.?�m$>n�ʾ8�M���,<)rʾ]���m�������/̾��1�'#n��̟?��A?����V�� ��]�bm����W?eQ�w����׊�=�۱���=� �>*��=��⾙$3���S�K/?��?�I��q����=>W����-:�y/?5��>���ߜ>7� ?
:3�j�����b>�=W>U{�>b8�>��>ᒰ���ڽ��?^�W?�h�eY����>�õ�E�]���=#> m@�..)���N>�EϻG��z�,;�Z��D/<O#W?G��>	�)�����g������==�x?ց?!�>�fk?��B?�<�U��:�S�#�Q`w=2�W?�'i?��>������Ͼ�~���5?k�e?��N>%h����X�.�eM�5$?��n?�R?�!��q}�|�����	^6?��v?�o^��r������V�<�>�R�>���>��9�;e�>��>?�
#�G��V���W4��Þ?n�@���?�<<�+�ᘎ=�;?�a�>��O�};ƾO�������q=�'�>����Xev���� R,��8?���?���>����a��;��=aٕ��Z�?~�?c����Gg<A���l��n�����<-ͫ=�	�QF"�����7���ƾN�
�y����ڿ�ƥ�>.Z@�V�6*�>#D8�V6�TϿ��v[о	Sq���?��>,�Ƚ�����j�Pu�C�G�
�H�b������>Ɏ&���	�e{���d���Gs��k��u?nMi����>vž/v �-��Se��Iԣ>��?2��>�׽�[R��½?rB<�����*���|��k?�h�?L
�?B+r?l�=O��M�Q���<���?�M�?��w?>���͚ɾCP���j?!\����_��)4�y�D��1W>�3?[*�>�-���z=D>t��>�9>6�.��tĿ������O�?_�?X�M�>GX�?�+?H���X��{����*������@?n�1>s���G�!�Q�<�ő��?��0?
E���,Qj?Ҽs��r���`C���y�)b�>�r;Uϑ�c��<�a�;��f��@���;t�Fǭ?O=@��?�+���3���7?���>��վ>�
�� 5�#��>!?.˵>+�����>�����N>S�?B @��?O���`����r>�7�?��>���?��">�ܞ=���>�Ѿ�Rh���>a1�>��>?�n'?�;\>��<xռ��@�T�%m��ZV��
T�#�E>�OZ?��e?��*=�7�����=��F��F����v�v��=�L3���=k����=N�>@�>���\���?4p���ؿmi���n'��64?ٹ�>�?U��>�t�H���;_?${�>6��+���%��@�e��?&G�?�?�׾K@̼D>N�>,H�>Uս����z�����7>T�B?&��D���o���>���?��@�ծ?6i��	?4�jN���_~����7���=>�7?O6�M�z>%��>0�=Tnv�������s�l��>iB�?�z�?���>m�l?o�x�B�V�1=aJ�>��k?�s?��l���w�B>!�?ޱ������I�!f?,�
@�u@O�^?����ֿ����:��L������=�k�=ە1>JKܽ�W�=K�5=�/�~*��V�='×>0�d>�eq>��N>��:>��)>����"�!��V��΂���C����a���Z����<w�l��Q��`���V淽.��������OP�Қ%��K]�a�=�ZW??�R?��m?��?�����D%>d��^AD=���w��=[�>��.?�kG?�(?�)�=�䞾i,c����|�����7�>\�]>��>���>��>�(?���R>��&>H��>=\�=��#=�$�¸=R>卭>37�>��>�C<>��>Eϴ��1��i�h��
w�q̽1�?~���R�J��1���9��զ���h�=Hb.?|>���?пf����2H?&���y)��+���>|�0?�cW?�>!��l�T�0:>:����j�5`>�+ �{l���)��%Q>vl?vZf>�u>n+3��i8��?P�q�����{>c!6?#���8�+[u��H�)rݾ�L>��>`'K�f����5k���i�Q$z=ш:?��?�d���˰�t�t������Q>��]>�=�Ϫ=mjM>@�c�_Sǽ[�G���0=4b�=�(_>L�?�r9>�2E=�7�>�n����K��q�>��;>��>}x;?X�?eG��k�'���M/�fza>ON�>�N�>L4>�;Z�%�=���>5�b>�~��d)�V����*�.�B>����,�W��j�Vs[=k3��*a�=�<`=e3���K��27=�1�?8��)���=�����3�T?l|X?
�z=�Zͽ��徵d�����D_�?T�@��?�Rݾ�{'� f*?��?���D�=���>h(�>\��}�<��?���3Iپ�0;�{�F=�h�?���?��c��쥿����;=��_?�e*�lh�>�u�HZ��X��)�u�|�#=���>�7H?�W����O��	>��v
?�?�]�J���x�ȿ${v����>��?���?�m��?��@�˄�>7��?fY?si>wh۾{`Z���>w�@?�R?��>:��'�U�?�ݶ?ή�?�G>8Վ?p�u?Q)�>�:K�U8(� I��.T�� g�<��=}G�>��>c�Ǿ�SP������{���w_�?o�6
b>_T=���>�/ѽ-מ���=�W-��Y��gU���.�>���>WkL>�>��>{B�>�%�>ª=+����t�|�x�7�I?�<�?���K�r��s=<B�=�	_�/r?�R6?/-;j7¾?Ҩ>��S?_)z?�Y?��>8o��Ĝ�"����W����;	�W>�}�>�,�>U����H>]�ܾ
;���>�>�ۼ��˾4���I}��W�>��"?N��>k�=v?��&?`7p>���>���Y����SO����>��>�H?��y?y�"?��f<>��҇��1��TZY�m >�n?P`+?��>U9��nϷ�k?=Z
�?��ڌ?��?��5�s�P?P�f?P�	?�pR?�^L>��º�11����I>-�!?n��	�A��&�\�%�?t�?Q��>͔��NG۽��ݼ�g��2���S?
�\?��&?����`�1���n��<��"��<����;`�"�S�>dI>�%���~�=�>�1�=��l��@6��8<�b�=0|�>��=҃7�1@���,?�B-��򃾰"�=�wr��WD�}{~>��L>�(��ǅ^?��=�ٛ{��ᬿPf��)�U��?���?�:�?�F��B�h���<?}�?�?p�>����Gݾ �ྺ�x�fw�t��->D��>d����z徳��������B����ŽH�����>�׻>�?��>�J>4��>������'�es����95P�+~�
9���/�yB#�������$yI���¾�����|�>�6H���>f�?>$G>��|>��>A/�9��>�k>CCg>Σ�>�N>ć>Ӣ�=Ki�T|���d?;��>�B�JA�E&*�bPp?D�?�iڻG$5�X�����о	��?�Į?�n�?u �=
nH�+���h=?�Y9>�¾vQ<?lZ=��{=VL�a���0��[�4�1	�J�`>@Ml��1D�0um��l�h�?�u?��=Ԛ��q�;���r�x=�r�?]�?{�?��3 ��sN�=I�)\����|u��qoܾc�!��2l�j���!���M���6�&	�;�;-?}cn?Nm̾�@ھ�ϫ�%�L�bEO��>��O>�>QH�>Y�g>�N���r3��WP��1���н�,?P��?�ˍ>λI?�:?�O?soL?�A�>? �>xį����>bJ;,Π>���>�@8?�).?x�0?Vg?��*?��b>&��-F��Ne־�O?t�?�?
�?:J?�ބ�2���(ϼ6��yw����BIu=��<��ͽ�=y�J\?=UU>%�?:/���2��T�ןp>��B?=��>��>�!����}�/����>{?��>����7r��4����>P?L�żn�<�5E>�٩=�ϻ�@�>�=��Ѽ7E�=�g��Iソm.�<-�=�=k�==�`=�h=�/=X,�>3�&?�e>ذ�>ds�0������â>>�$�>H=y>%��=��ھ�爿N��6_�p�>I!�?�5�?��=�9[<���=#����d�>M��Ǿ(`P>a��>b]�>[p\?���?�9.?1?���<P�����|;��s־�*?D!,?���>����ʾf�}�3�ӝ? [?<a�\��q;)���¾��Խ>�>p[/�'/~�v���D�������/�����?���?�A���6�Sx辈���>\��-�C?�!�>�X�>.�>4�)�E�g�q%��0;>���>-R?dF�>�O?�z?i[?�U>��8�j	��R����L��>��??���?���?�Zy?���>�0>BU(�hg߾�<���[ ����X����R=�]>%+�>�b�>$ө>���=7�ʽ����T=>��;�=��a>K�>�7�>m'�>�u>�~�<��??���>WD;����,ԕ��N3��6w?�v{?���>��i�J� �$z<�ĝ �B��>!U�?y��?RO,?޵�~�=�������6�D3�>2(�>�>��G>�,>+^`>��>+G�>�C�@�(��	G�@GO��?9D?�A���n���N��L%=�v�����ړ� {�}��"�v�H�½�����j��¶վ0���ʾ}A�����-n�����?�4�=�Z>[��[�E�9���k�=��J�4CϽ�^&>(@���������q�����Խ��;F����<Q+L=�'��ִ�?�[?B�o?��h?��>��>v�I�0�C?�J>ϱ�?�e�=����͑о��1��(����'��eU����Ⱦ_��=�s�=��N>�R�>�?�p춽��,>�;u<OUB>&����ɜ=���=3ʯ=���=��=���=|hB>�5w?H���v����1Q�H[�q�:?�5�>�z�=f�ƾ(@?
�>>1��앹��\�/?���?aT�?��?�ii��a�>F���󎽆i�=����02>���=|�2�f��>^�J>���WI��u���G3�?n�@Z�??�ዿ$�Ͽ�`/>LL8>�$>�R��g1��Z�@d�Im[��t!?Z;�@c;$j�>�C�= �޾�ož~Y;="~9>��g=o���r[� F�=��z�o8=|�e=g�>�D>��=)����/�=��E=��=�bO>뎥�\B���,��n5=�c�=�a>R�%>sI�>^?��?=�H?�>60���ھP���Pr)>��A�CӀ>�5�=�#>˅�><�Q?��[?u�N?��>�'>tO�>J�>�)�u�k�CS���(���J?��W�?vz?R�><4<��-�����H�W�|�d?װ ?��>5G�>����ο��%��I;G�a=\=�pY�ɩ>�iA��=J���=�Ӈ>�>�^�>���=ڋ'=x�>���>9�=���^�`={->��	;� M<�f	=�nJ���b�z������s2�=7!��P99L��k`�ֺ����9��E
>���>��=�O�>�@�< d��/)N>��� �C��m�=Ѯ��J8�tL�Ѝr�!�+���Z���[>2��>���������e�>��>f�2>+��?��t?Ũ>�ġ�\h��T��^�A��=���=^��=R$a��>H��Qf��N�wWž3��>���>T��>�
m>d,��>��y= ��c5����>ڕ���������q��0����8�h�������D?4A���<�=*~?ޚI?�ݏ?���>GS���3ؾܼ/>Q��0�=���Mq�����z�?�&?�E�>M!��D�<�Ǿ�C���?&TQ��"T�{P����J��� �� ����>B|�����ۻ%��C���ٗ���?��E��%�>�`?வ?�T���ho����5��y¾F�>gTw?��'>7%?:��>��j����Z���g>���?q�?���?��>o�=
�ݽV��>t�?ޛ�?�&�?ŵp?iF����>�3�;�=�Ϫ���>��#>�P<&Ԃ=k?�??�k?X>�(|���ξ�n��[�9��J�<���>m��>�![>\��=;�_=_I=?�>��>uC�>��>�?�>�>Uw�R��^�?��D>�$\>t�H?h�>�f�=&2>�e�����P%��:�҆��'�z�뽽�	�/�*>�<��>vп�-�?��>Σ�m�+?Z"�R�j=��>�V2>���a,?�">`��>�Y\>��>�(>�H~>6��=j�׾s�>�w�����&F�dDK��˾��j>/��0s$��	�
���\W��.���r	�Ii��J��V�A��:��܎?�轮�c��(��:��?�>��.?os���O��>��>E��>���S���͋�'pؾ.��?���?��y>^��>�L?��?��G��tT��P�X�f�r�A��`�db�Y��ӄp��J׾�3���\?dÀ?/�N?��==T>9Ђ?�$�ě�=Q�>T0F��tA��6=��>�ƾ�2��1Ծ~)׾������>�Ӏ?k�n?���>d�A�
����@>>��<?޽:?��z?�a=?j6?E�5�-�.?�sA>aF?D?�/?j#(?bH?��?>
�=�ƼKx�<�M��5���jؽ�vս�B��j��=���=S��T�ka<,�M<&&�#ʀ����<��M�;��<�2=�P�=�l�=�u�>H�S?���>��$>�dJ?"߂��W�`;]�?�>��y�������?����N������>�	�?_�?�cL?�<�>Z�u�����]�=��>��=ޅ<>�Q>l�8�E<�<�.@>���=0=��'��{�޳��z�B��Q^z�Ѫ�=�1�>L;�>`A���6>�����z�\@�>7�R�:���zgH���H�3�,��XM�+m�>bE?��?�E�=��ƾ��<���j���*?�9?fpJ?�.|?���=�Yھ�(�t�G�x��9w�>�-B��_��@��IꞿΎ>��/Ƽ��N>]6���k	� �v>�����ؔ���eK����P�SCݾc���b=5�~��$ ���'\�T.h�^���J��Q��u鯿�:?��'>��7�܅��kȾ�����>��>�h꽜8�Dua���¾���=\�>HJ=�v�侴�:�3��76�>iRE?v`_?�u�?6 ����r�{�B�����U����ü��?�Y�>vX?��A>�x�=5���|����d��F�,�>E`�>���R�G�e9�������$�Oʊ>%?��>0�?q�R?�
?�`?�*?�/?�/�>C���B����4&?H��?���=��ս�;T�2+9�!*F��v�>�B)?2�C��c�>v?�?W�&?t�Q?��?(>�~ ���?��o�>CZ�>h�W��I��p�`>�J?�&�>�#Y?���?��=>�Q5��Ӣ�+B�����=y�>�2?y�"?0k?S��>ow�>?a��y��=��>%c?�/�?�o?���=�?]�1>'�>�v�=���>kf�>��?5O?O�s?��J?R��> �<����"W��s�r�/�N���t;��E<1�x=WW�Gs�O��/�<`�;����#�{��u�*�C�ֲ��s�;��>��%>������=ȴ�-c-��	}>����.��c~�ۍ��Oia>Y�>�E ?W?>����	k>�f�>��>5�&�4O?���>�! ?�oe=a�����on�*�>�4#?�ǽ΅������e���7�<b]?�oF?}���k���<c?p.\?����?@��ָ��^��澗7T?�S
?Z�J�)��>�?�+n?\�>��h�ӑo�x۝���^���i� �=�%�>ɕ��`�;D�>(�7?���>��[>���=��ܾoOw�%i��i�	?BK�?��?x��?��$>��n�f�߿!�a���o![?���>�{���#?P �:ھ��������&S޾�٩�����(������� $��~�����u
�=?}?OK}?qw?AKZ?'����e���\���v���O��%��y�Z�F��*C�u�H��	l�C��:��ାVD4<�\�k A����?F�'?��0���>O���I��ov;�JC>O����`�4>�=jȏ���9=_�U=�h��:.����� ?��>�F�>�<?Nu[��=���1��a7�������4>��>!|�>k��>Z��:'�,�L���Ⱦ��O�н6v>�~c?8�K?/�n?�n�	1�qt����!��'.�i��C>C>�>#LX����&.&��3>��r�o���\����	����={�2?n�>��>�=�?�?��	�`Ӯ��x��_1�u�<�=�>b�h?���>=��>gMн�� ����>qm?i�>���>er����N�w��۽y��>���>�e ?~�`>�8.�`'^�q(��s���J4�e�=3=c?%8���i��ˍ>��N?��;���<���>��Q���#��@޾���2>�,	?L��=#�/>�Ͼc��y�-}~�;D)?�T?'꒾ʫ*�[�~>��!?��>Vۣ>��?��>qþ�"7�'�?�^?+�J?9tA?y:�>�=4����]Ƚ}�&�I�,=���>�[>J�m=\��=��D\���O�E=�=¡μ�칽/<g"���7L<���</�3>�ۿ��E�w���-C��[���C�?o��v1����G;����Ps��;����a6�?:���`�灾'd����u����?w�?�p�������E��pу��� �q��>@ J��������ANZ�ĩ��7���������)���e�E }���s�K�'?�����ǿ񰡿�:ܾ0! ?�A ?5�y?��5�"���8�� >XC�<�-����뾭����οH�����^?���>��/��q��>ू>�X>�Hq>����螾q1�<��?8�-?��>ώr�/�ɿa���r¤<���?/�@�N?��M�pm���!�Z��>�0@?��>�ܪ�Mw�sm��䂯>p�?uȧ?��|>�uL�R]����]?(�.=�v��S:�ۣ>�h>���΅��bƑ>Pf`>�4���Iy��5R��`�>DJ�>�ټ �8��}���=E�>�ߒ��g�5Մ?,{\��f���/��T��U>��T?�*�>R:�=��,?Y7H�`}Ͽ�\��*a?�0�?���?%�(?7ۿ��ؚ>��ܾ��M?_D6?���>�d&��t�م�=�6�N���}���&V����=]��>e�>��,������O��I��V��=R���ƿf="�9?��6�<���;�Uy�M��[���f�i�0��u�n���,�]=�l�=�KN>E�>�Q>�\>"�W?yto?��>�H>���Ps����Ͼ�g��S*��%"����#��ߤ���������	�oj��i���;�'=���=Q$R�H����� ���b���F�9�.?�j$>�ʾ��M��+<�vʾ`Ǫ�>H���
���:̾�1��$n��ʟ?��A?D���}�V������|��ɯW?A���u��Z_�=�����q=�>�6�=��⾊'3�@�S��4?��?�J���������>�Yؽ���<`cA?�\�>�<��,��>�)?F0X�{Wнm�M>rS�=��C>
(�>���=b����?����?�[?.m6�с��>�O��p��t��=u=�=Ǥ9��6����!>�N�=�b��)�;*
�R���se?�c�>( �I�a�"k���.�K��=��?�>'?���>/Ƀ?�J?�W�	���
6^�7� ���%�R�^?�P]?�Ĵ=�]����LM߾�j?k�_?Q��>�=򽮬���p��Qվ�?��L?�"!?���=І����w_�F��>��v?�r^�ls�����O�V�V=�>�[�>���>��9��k�>��>?�#��G��ﺿ�sY4�!Þ?��@���?��;< �휎=�;?V\�>5�O�?ƾX{������ȓq=�"�>���ev����4R,�k�8?栃?���>쓂�������=�ٕ��Z�?}�?���Dg<Q���l��n��=�<�Ϋ=���E"������7���ƾ��
�����ῼ̥�>DZ@�U�o*�>�C8�]6�TϿ(���[о�Sq���?B��>_�Ƚ����9�j��Pu�_�G�.�H�����-<�>9����B�7�ѽ�����:I���=���>�=��� ?�ð�����3о.��nG�>Y2"?�ٶ>�|{<.m�?�D�ot�E����
��KZ?G �?�	y?_�y?G	>U�9��|Z��`��?�u?c��?xLj?s4��e��=�p��j?]_���T`���4��GE��U>�"3?�B�>�-�s�|=�>���>�f>�"/��Ŀٶ�M���W��?h��?�o꾰��>C��?s+?�i�48��6\����*�Dw,��;A?|2>����z�!�x0=�Lђ�^�
?+~0?�x��-�c�j?K�x�����$'���^�hb�>��=S@2�Ɩ:>pg�=��a�C@���`�����?E:�?�3�?���0���6?<�>�r��8���P���?S��>Ɛ=>)޶�]@�>��ҋ(�N=S>���?$@^%?�[��򮥿��>� }?Ԋ�>�c?q=�l�>�Ԧ>������=��{>o�=�@'>�/?�*E?,��<.�,�����>�:��w���C�AZ8���O�{��>�C?l]?�`�<H�A��1>�"P����G���h,��?X��y��c��x�M>���>
�v>k+F�d陾��?Mp�9�ؿ j��p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>D�Խ����\�����7>0�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?��?@���C~�H��J-7�Tb�='�7?	Q�{>��>���=Ahv�*�����s�bö>r=�?�|�?u��>�l?3�o�F�B�2=�.�>��k? |?`�b����\�B>�?��[����7�E-f?i�
@Ys@��^?뢿h�п"]���༾������=D��=*Z	>s�ٽmH>�Q�<��<��3���>	�>��f>�q>P�n>.9>Х>�w��B�"�����鐿iE�MQ������I����/!���J�2��7	��������7����l��X������L�=�/W?��N?��o?�??�HL�~8>����l=^����=�q�>˘+?�F?m[(?/�p=�ۤ��.b����ݫ�c�z����>R>U�>��>=W�>��<�)g>jB>�O�>��==Pv=�-<vl�<n�T>��>���>��>}C<>��>Aϴ��1��m�h��
w�b̽/�?����R�J��1���9��Ԧ���h�=Bb.? |>���?пf����2H?&���x)��+���>{�0?�cW?�>(��_�T�/:>6����j�(`>�+ �{l���)��%Q>xl?j�e>.3u>�L3�2a8���P�@�����|>K6?���
?9�(�u�b�H��Pݾ��L>K�>eTP������@��i��1z=�\:?p?7���ϻ��P!u��<���gQ>n\>�L=Z��=�oM>B�d���ƽ��G� .=k�=��^>�?q/>��=Ux�>����XJ��>[�?>'�)>&C??�#?\G��#��\���Q�0���q>�E�>�>�>��J���=|��>�}`>� �kO��d_�LK<��oQ>��k��^��x�v=���H��=J�=?����:�#17=Q{�?\������tϾ�V�ƧJ? �??G�2�!	�=y龽眿������?��@w(�?���a�<���
?S�?ֳ���r�<�>�>�9�>۔��S6���>������Ӯ;���E<���?���?~=Ο�D�����l>o�.?�4�Rh�>xx��Z�������u�m�#=R��>�8H?�V����O�\>��v
?�?�^�੤���ȿ6|v����>W�?���?g�m��A���@����>:��?�gY?qoi>�g۾F`Z����>ѻ@?�R?�>�9���'���?�޶?ԯ�?�H>	��?��s?Q(�>��x�q%/�n�������=V��;p|�>��>����&�F��͓��W��߂j�n��m�a>�$%=
��>�����A�=���,����c����>�Vr>* J>`e�>�� ?Kn�>e�>�P=9������;���K?��?���+4n�&&�< ��=J�^�^-?H4?��[���Ͼ�ڨ>�\?���?%[?zW�>���;���濿T���P��<��K>�:�>>�>S,��?K>��Ծ6D��u�>�ŗ>M���Aھ�/��j���yD�>d!?<��>��={�)?Te?��~>#T�>?�(���jfB��.?	0?�N?I	�?l?��ᾍ
/����ې��Q/�گ>��z?��6?�eC>�ך�Py�����<6�m��=�<П�?�&x?d�*?��?��+?I�9?�Y >m)�Ǘ�oa�<�>hE!?���S B��%�q��X?��?���>諛�>ֽd�Ҽ3��T:��.O?5[?�D%?�3�L`�]�þ��<g�q���+��;�G�o>S'>#s��eu�=�)>Ō�=��h���3��!�<�F�=7��>q��=l�7�����6,?^�D��̓� �=��r�"xD�>�"L>O���Y�^?q=���{�����r����T��?q��?�i�?U���̗h�7 =?�??�>�H���h޾���T?w�Xzx�)a���>���>HYo�0��̋�����nG����ŽI�IO�>Yv>�< ?T��>N��>�[�>��w��X7��㹾��= R��Ѿ�� �D5��E���@1����<Zպ����U,�>Rh����>ƻ?�>��>�Av>���=���>�)>��s>��>��U>��0>��="�#�*,-��
_?��+0�����,�q�?�H�?�) >�3�r��bgѾ�y?>Ъ?S&�?_E>ڃV������>;�>xή�ٷ@?�z�=UIa=���=�7	�s]6�$B�=Q��Ə�>@s���([�Ww�$�ew?�>?���;���O	:>7�Ѿ�|�=V�?���>�%@��{I��:F�5�E� k����>�ξ�L۾�?��s���F���Ɔ�m����I7�b��<m%?��g?�ɾ=���Ǡa�O�4��;��c�=�o�>gm>0�>Ƌ�>n�о�5�<F�G����0�6"%?e�p?�]�>ŧI?M�;?:�P?v@L?���>�C�>�I��en�>*�;�c�>���>�J9?n-?�0?*@?S0+?QWb>�D��b����Pؾ�?�?@?� ?�}?;���ýyl����R�Vy��S~��x�=?��<;ٽ��s��S=�T>�C?v��#9����l��>��4?u�>���>�����)����=N��>8?��>� ��[u����
�>ZMw?�5d�eX<��)>�>B�w:�%�<
Z�=_{�֩W=11ϼg	���[l;%r�=Ŗ�=��!=R�I<=X�(��*�'�1��>�+?�p�>�.�>�i���I�z��s݄=�4�>l/*>2t)>85�	���/Ԗ�HX�Kt�>�k�?P�?0%�<�>�=+:�=�G��)�O���𾬾�$>��>��?�t\?�6�?�R,?�,?/s�<���阗������ƾ7�?x,?܊�>w��Ҵʾv�-�3��?N[?&<a�}���:)�l�¾�ս��>�[/��/~����D�����s���|�����?l��?TA���6�x������]��2�C?l�>Y�>��>��)�$�g�6#�Z2;>ً�>R?`�>�O?�z?�*Z?n�W>);9��9��Ù���b�ˈ>��>?�G�?z��?�gx?�s�>�c>_�'���޾�s���g �$,��t��e�V=X2^>�ʒ>���>^��>�J�=;�Ľڷ���>���=S�_>W�>s�>.��>?t> �<f�E?� �>�$����p��Ӆ���ފ���s?k�?r('?���<�1��|E�����)�>�M�?2S�?��(?�P��g�=�W������3�e���>�н>��>�^�=��~=,f >8+�>��>�Y&�L��I<���f��??kE? ��=|3ſ�k�q�S��
��lH3�o}��3�\��ș�{_��8�=���@/��Щ�v�e�G���Q���\���2��e���>b[{=�(�=}��=j��<ɂ���=��F=d���`|"=7W���/X<����ɗ����5�����'<~Jl=���;�阾��?S�0?�A?^A?&�>D�>֣=�#?%}P�^m?�>)�ͼ�쎾NsV��n��*��Z������?�����0��=I���|�=s;>o�l��o>�u(>�u���Ԝ=���!�->���=�gL����=s\>�>6��>j4w?���������+Q�]�v�:?�Z�>�f�=.kƾY#@?b�>>L2��-����^�O1?4��?�N�?d�?[Ni�`��>���"����=�b����2>Hz�=��2��й>:�J>�t��B���`���5�?M�@c�??S㋿��Ͽ��/>ng8>̂>tWS�u�/���R��?\�`�U�~$"?Ph;��ʾ�a�>cV�=�۾�_���&"=��0>-rR=j���7\��t�=��p�I=8c=��>��D>�µ=����Oi�=�Q=gR�=v�T>�;����/�|h<=u/�=,�]>�1>���>#�?kx5?x�g?��>6�I�S�پ���C�>I�>0d�>�V=��+>���>�t/?�9?¤L?���>h_�=���>�-�>�Z(�-n��{�}y��9!�[�?bZ�?i��>���<Bd2�u&"��?2�j6��?Ն/?�M?�/�>���]��p(+��K����J�=�:������1[>����vs8��4��<׼>�	�>�U�>wx�>�8�:5�<�>���=&p�=�W�=��<�`>9ז�����g�v:=J�=bb<�C���M�V؈���ڽ�Q�/�<9��<��=�	�>���=��>�@�=	٥�s$9>�����K�Η�=��a&=��R��p���/���T�QI>��w>����_��U�?0BG>P�h>i3�?źo?���=?h���پ�"���N��Y���Г=�T~=��I�@38�sx_�
K�{�ʾ���>D�>���>O�l>��+���>��_x=9��kn5����>Ô��ܦ�u��'q��7��z�h�D��ΙD?KA���[�=J�}?ҼI?�ߏ?���>ܙ�O/ؾ�/>����
=B��'q�-┽��?��&?v^�>2��МD��ž<��M�"?��\=d�P�INm���.�O����pz�>��þ�3��K��??��H<(��M;�+?�Z?��?�Ʒ�g�j���	�M�р�"l�>HN]?���>'/?Q�>����³��۽P��>�?���?��?���=��='F�����>� 
?�,�?�z�?�mr?�<���>-Q�;9J!>P���k��=�J>Kp�=h��=��?2~	?�	?�9���z
���B�%^�:=��=@[�>5�>lt>A��=�lv=Ǜ�=qPa>���>��>�#g>�=�>�8�>� n�]�ϾX] ?Ћ�>�/�>o�B?(Jt>W8�=0Z�|J#>o��Z��VǬ�rG=2$�?��]�=oq�;��� e�>3<���ݔ?��I<���X�?�}�$�^=&ut>"�>�L��3�?���=x��>�ӛ>�t�>��>!�>*�Y>�F�0�">RqȾ��%��S�f�S��'���|^>����a+����o�=�I�tKӾ�,�M'n�Q����Z�G��䯊?v��WjX����ս�m?�i�>�A%?|G��2�qr>l��>��>z;
�j����g��UݾWy�?Vk�?�z>Ǔ�>ԽA?��> �Z�9ڸ�KJ��;s�y_<�|`�b�e��i��e��Mƾ�H�:�s?l��?�f?�c=�#>���?u1 �����P	�>�T�ףC���� G>nr
��K9���:���t!M����>c2~?GG?�h�>�d��0����n>4�,?��2?�2p?��1?��2?u����1?���=.�#? ��>/ .?��?���>�>�-�=3~<�N�=���~���������2���{)=��c=n16��)�<��1=e&;,�?���̻]䢻U�{�4f]=��~=�=��=�ϓ>1b?�6�>[�6=�h[?:x��f��U�����>��ܾ-����q�'���1y��u@?Qc�?Ɇ�?<�'?�Ĩ>�b��y}� XB>��>Bm�=V�>vY*>��=!�s=��u>І�>[�0<���J i��������)���x�.�}���>^{>�
Ľ;�(>���ƙu��	l>��S�(ཾ�
S���E�=�-�6qc�m�> yD?[f?#��=.*پ��r���i��.?EQ5?RQ?�?ۭ�=���!/��#H�\��=�>z̼�D
�g����u���:��� ���k>qS��rݠ��[b>���q޾o�n�EJ���羖BM=��uTV=���վH/����=##
>3����� �����ժ�G0J?e�j=ts��eaU�m����>�>Yޮ>��:�?�v��@�>���7�=˶�>�:>�y��2��
G�48��?�>&RE?�U_??��?���o�s�q�B�K���z���߸�	�?��>�\?%0>>�|�=T³��p�*e�B�F��f�>x��>1���+G�bZ��)���N$���>*�?wx#>�F?��R?��	?��_?P*?.I?��>o㰽����A&?���?���=k�Խ��T���8�#F�)��>u~)?��B�F��> �?l�?`�&?�Q?ϸ?z�>c� �R?@�Ԓ�>-Y�>��W��a��1`>a�J?3��>l?Y?xԃ?#�=>C�5�)䢾�ǩ��?�=l>&�2?�3#??�?���>R��>蟾P�n=�;�>9^b?�?�%p?�S�=�e?��0>w��>J
�=7[�>��>Y�?U�N?qs?[K?��>#Ʉ<�?I��9�p�}*A��
�;-�[<�5}=��r��!�9��<ܭ�;CR���Յ�f���B_I�ޘ��ʆ�;�,�>�d�>�о���=�9˾��"�r�|>��ֽ!��Ɖ���k��K>�ޔ>֓?yx�>����=>:�?�k�>�c$��QP?-j�>T"?:��=˦Z�8����(���G>�?+ϧ=�z��k���Iz�o�'=�Q?{OH?����-��jPh?�(]?�MҾ0_G��᜾-���$0�����?�v=?��?��A�>�ݑ?��C?�c?����OX�ȧ��P]�,O����=�Ņ>��hN��N�>;*B?�B�>���>+�d�,{��S���nʾZ�.?; �?Ě?a�?E?�=��h����>�	����E?�< ?��s�&-?B�y�����D¾�g۾⬭�
���r�������A��LE�ϳ�Za>�;?x
}?���?�I?R}��M�F9��5d�D0M��J���6���8��V�<�G��탿�8����
h���L>]�v�-�@��6�?.J$?:,�o&�>ɋ�������ɾ)|G>yj���.
��B�=��Z�[07=��g=gv\���!��)���?~��>���>�]=?,�^�ܲ?��`1�8\9��s����#>�D�>�}�>��>�`�-�+��սE����p�"�����u>�c?SZK?GTo?>��1��T��w� �0�>Y���{C>˛>��>`)Z��� �\�&��c>�uss��������h�	���=S�2?_%�>�>���?��?��	������w�R1�r��<%��>�h?�h�>A8�>Vѽ&| ��m�>Y�q?s�>�j�>���|�u��=V��>~�a>���>�^�=O�}� Qq������N���.���`�B?
v�+�b��C{>G�U?�!E=������>a�`��$��K��+�S���=F?v�>��5>C���*�����0����(?�x??:���~)�p�z>�]!?40�>�ܡ>m�?`��>�þ�1��z?��]?3vI?�1@?q��>.�0=J���̽BH#���6=k��>p�\>|=J�=���)�]����z�A=��=�?��U���?��;�;м�<��<IC,>{lۿ�BK���پ�����;
��舾�Ĳ�,g����@^��1���Ux�N��>�&�YV��2c�ܢ���l���?�<�?1w���,��ڰ������U���M��>��q�ŵ�@���7���,��\��Ǭ��c!�f�O�%i�˻e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�A??D(�r}���1=���>��?G�<>�-��"��˫�n��>��?E�?;w�=x�U����vue?��<��C���»{q�=/��=F�4=�y!�D�=>:/�>Z5(�m�A�4��ֻ->�x}>�sA��6��]��� =�cg>S����z���Մ?[|\�of�Ҥ/�BU��a>��T?2*�>^`�=M�,?'5H��|Ͽ��\�+a?J1�?i��?��(?�ݿ�Qܚ>��ܾ�M?:A6?���>�^&���t�̈́�=��P�����A%V�w��=��>�>�y,�9���O�������=W���7ƿ�$���@=$�:�)f����������_�f͝���p���{?b=`�=g<O>]�>�*T>��V>[�V?Fl?�>��>A�ݽ��4˾�7�LԄ�Z�!�j��pg��*����Z�ᾋ���3���R�ž!=�,�=7R�l���A� �f�b�H�F���.?�v$>e�ʾ��M���-<xpʾ\����ۄ��ॽ�-̾	�1�"n�h͟?��A?������V�N���W�r���W�W?<P�һ��ꬾ��=������=�$�>���=���� 3��~S���/?�:?5	ľ�����'>� �q.=Yc*?;( ?+�2<$�>�$?��$�#��1\>�3>�h�>���>
�>����{�ҽ�*?#�S?�]��P���̵�>�_��X:|�d�e=�>��3��Mļ�AW>
I�<����%����F��R]�<�$W?ઍ>O*�� ��`��Q��>�==t�x?~�?j#�>�qk?r�B?K�<_����S�h��ew=��W?s(i?g�>烁�.�Ͼn}��g�5?��e?\�N>lLh����d�.�'R��#?��n?&[?�����s}�O�����\b6?��v?s^�ws�����G�V�f=�>�[�>���>��9��k�>�>?�#��G������{Y4�%Þ?��@���?G�;<��T��=�;?n\�> �O��>ƾ�z������>�q=�"�>���~ev����R,�c�8?ܠ�?���>���������=�ؕ�Z�?��?c���v]g<"�� l��o���Z�<�ǫ=���V"�����7���ƾb�
�q���Ϳ�n��>�Y@oK�S*�>sD8��5�eSϿ���A\оRRq�*�?}�>��Ƚ����\�j�}Pu�X�G�3�H�����6~�>��)=8;Q�H���F��9CA���=|��>o��<�:?�C��7�!о�)��m�>�4?g(�>T�g���a��y�?*�$�3B�6���%�)��h?m��?k�~?��`?5�B>�Ӝ�fB�Z�#�l8?��?e�?<�w>)��8^��j?__���T`�ю4��GE�'U>�"3?B�>ԓ-�4�|=�>4��>i>�!/�ˍĿ�ض�!���V��?|��?Go�z��>��?vs+?zj��7��O[����*��W-�0;A?�2>���%�!�R0=�Ғ���
?`~0?2v��-���o?�Ap��&���=��!�����>��>Gq�=�X>��q=N�F�s���eq��}f�?R[@��?��μ�6'��2?�i�><R��W,��=��=���>��^>�k=>c���=�NZ��#5�5�p>���?t@���>��������F,�>�(|?-��>?7q?&1�>G��>#��>W�Ӿ���u�a>9�B>�"#>��?��,?VO�>��=72�;""�C�M��e��e�x���@�,V�>�KH? \l?��%>��C<�Ä�a�#�l ���޽��>����0��Т?�ib�=���=.�>�K�i{н��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��a~�߃��7����=��7?�/�P�z>b��>6�=�nv�ۻ����s�m��>�B�?[{�?9��>��l?�o�L�B���1=�K�>�k?�t?�o�7�!�B>Ѷ?ٱ������K��f?�
@xu@��^?��ſ�M����n��վ���=�B0=A��=T���#�=�:>�>yn=+t=?�>��=�JF>�[>m >��>��z�X/��.������-]��9�k@�l䊾G�%��>��`}�.�վv�۽�d��w?c�P���e�V<���=�_Z?|�S?i�r?�B?A�q�f%>	��Vm�=`��>ę�>(�+?��;?[,?��b=+����h�)G���~���[T�j�>��]>	��>	$�>��>�=�<}i>>p">{"�>I��=!�P=�&6���!=
�T>���>!'�>�!�>�C<>��>Eϴ��1��g�h��
w�j̽1�?|���R�J��1���9��Ц���h�=Hb.?|>���?пg����2H?(���v)��+���>|�0?�cW?�>"��R�T�.:>>����j�2`>�+ �~l���)��%Q>ql?Ȋi>��u>�1��g8�<ZN�͓��ў{>�D6?�����3�c�s���G��!ݾ��K>2�>qKX�c����������}k�xw=j�:?�?%��O௾/�s�}}��:�M>��`>�
=炬=
�J>_a���˽��K���6=�u�=�(_>�?1�6>��F=eT�>a]��2�L��Ӯ>s�<>��$>��<?�V"?���
n��ǁ�*)��5u>&V�>���>c�>�cM���=��>��a>����p�u��)9�dBP>N�s�;y]��q�{��=����5��=@"�=+���J�u��<L�?o榿$���:N��9B�n�!?�;P?}
�=Y��'�sv���] �js�?Zs@y�?N(��eS�nD(?�ϐ?�$����=��>���>vM��x1���?%����T��E����?�w�?k8���G��Nk��QP=�f+?����Jh�>�w��Z�������u���#=���>�8H?�V��u�O�|>��v
?	?�^�˩����ȿ!|v����>E�?���?��m�cA���@�ς�>=��?^gY?�oi>�g۾�_Z�y��>׻@?�R?N�>�9�}�'�n�?�޶?���?��F>���?ƙp?���>E���F.�]�����l=���wN�>���=�����H��w��ha����i��&���N>�H=J��>Ҷ��h����=�s꽶����oŽ6��>��>��C>�˘>p�>�U�>>,�>�a<01���A���ے��lO?d$�?��ɱ|��@>W����=�C?X\=?Ņ+��Lv�.�>��A?(�V?)]?s��>��1�=����Կ��������ȏ>}��>�	�>|/�`!>D'��݀���>�6C>�x@�4�⾷m��:�^=L�f>� ?��O>E�{���?�"?�٥>e?nG��4����;�%x�>�e?�+?��?\�,?�(��+=���{�L��z�m��W�=o�r?��+?�n�>�7�����Ё�3�=c�=��?��?�s�uy$?{��?#{#?C�U?h�>e�+�7������d�>г!?6��]B��&�����@?�?�X�>���n�ֽ�ټ����D��I�?a�[?��%?$e��`�%�¾��<h���B��2<�z8���>h�>b�����=H�>!�=3�l�}�4�m@`<2!�=���>�a�=L9�a葽�<,?J�G��ۃ���=��r��wD��>�JL>����^?�l=���{�l���x���
U�� �?���?Dk�?�	���h��$=?��?~	?"�>�J��`|޾���HPw��|x��v�"�>���>N�l�6�M���㙪��F��8�Ž������>'�>�4?�>~�M>���>������&�82�9���\�.���7�i�-��Z� ���� ��O�J����z�`��>���=�>~�	?f>�
z>��>C�:�>�QS>���>¦>�ET>%�,>���=�- �/ݽ�/_?dfо��E�S��.��g9?���?��F>w�5�HMq�[���7n?�?��?Afw>�4��J	���
?Z.�>.����>?��_�G>�<��=�|���:̾��q��[y=�و>���]?�wo�! ��
��>
�
?-�#>�,���|��C���V�=���?��]?Ӿ�L��_���X�� a���ܽ�[s��⾢�D�S�z�!🿹���e=�6�+��Q�=q.?,XL?=>�量�q��a���8��� >���>^j?:��>I@R>�����Ո����m���P?��d?B��>�I?��;?tP?|jL?H��>�_�>�1���d�>���;:�>��>9�9?p�-?�80?�y?�r+?~5c>ks������g�ؾ^?��?M??^�?ׅ�gý����g�
�y�@j���=��<�׽�Bu�{\T=,T>_?,�˼��Q�N��&5D>s�,?��?�A�>�������_}"�_P�>@�?�ņ>���fa�������>��}?aY�K^�<H~P>♵=�,=椋=8��=�ڎ<�R�<˸v<��A�U�A=v�>^�=ڞ��B>4�J�5�G1���s��:�>`6-?<�>?��>3Y����w8�8�>�Y|>K��=�P�<���)���f��L���dN�>Fr�?�s�?j��<s9=��=����l�
��9 �&Ⱦ�>�n�>^�?cL?��?�0.?�{�>�Ȼ����T��KY��=�T�?�!,?H��>���E�ʾ�䨿@�3�M�?�]??*a�����.)�@�¾�ս�>LI/��&~����")D�6�������|��k��?>��?˒A��6�tm辂����`����C?_
�>�W�>��>��)��g��'��8;>^��>�R?�"�>��O?�<{?��[?pT>��8�0��ҙ��2���!>D@?B��?��?y?�v�>��>
�)����Y�����[��₾)'W=Z>D��>p(�>��>k��=n
Ƚ�5��~�>�"e�=�b>@��>Ѡ�>��>0�w>S��< ]F?צ�>�����2=����}�����t?�	�?"?�5J<R��$eB�Xs���s�>�5�?���?�I+?�QP����=��м؄��\
f�M�>IY�>0C�>G�=!t=Ė >��>7��>����=�� >�e�^���?u�E?9�=��̿瀿��C�Rl��ad���-���y��]�9�|���=��7��B�"۴��Y�[����6�����A���H�dM�>Ř�=�>�;7>4}=N�=���=ˊ�<�k�� �Z����YY������W���^�c�#;~0�<�K"�L奾vҍ?)6F?.�H?�m?3��>��=b��=�?v���9a?x6>�#�<a���&<����-��y�������T���z���*=��\��}>z��>>�<$:<��J>�ܽN�>rk��[r=��[>�==���=��*>*`C>��>��{?�?�����ϗ[������6?�x�>�Λ=�Y�al?��>�Ą��T��h���v?�\�? ��?���>l6�x͹>�;���f��,h9�Ā<	&�>��J>6��py�>��>��;g���ղ��m�?;@�-B?M����˿>_.>�8>��>GrS��1���\�>�a���V��� ?�-;��]̾�j�>K#�=�dݾ�ƾ+�0=h56>��c=�J�:f[���=(w���?=][l=-�>2E>q}�=���Bh�=ѺK=���=K�O>��/���9���.�.=��=#~^>Z7#>�1�>�T?h0?�za?Q[�>nbh��8Ѿ�{���>V�=���>��s=V�A>o}�>Br8?�'F?1M?���>CP�=ۢ�>,��>�+�E�l�^�䱦�aD\<�s�?`��?��>��<e|>�gw�'�>�Cн5#?<�0?]�?B��>�m��8ο���ܐ��L��8�>����q�é*��
�<�a�=R�����=��;>|�>>i;=���=��u>���=]��>FM�=��ὩJ|>N9�<wþ=UZƽiuټ�[����-<Xt1={���t�=Gؼ���=����vJ�=,}�<���[�=���>/�>�"�>�K�=+���s1>�����L���=�a����A��oc���}���.�t�5���B>nZ> �4���J?�IY>��?>"J�?��t?�@!>�r��վ����ɶd��NT��~�=F->j=��a;��#`�3 N���ҾW��>?��>��>��l>_,��"?�g�w=w�Bb5�l�>�|��l���'�(9q��?�������i���Ѻ�D?gF����=�!~?��I?>�?$��>����ؾ�90>�G����=B�N)q�k��a�?g'?Җ�>��l�D��Ǿ������?:���?oA�u����=.�ci���i��W�>@=پ���@>�߻��X���9F�Sp�F��>��X?��?*F��|�x�0�\��&;���&�6�?;n?*��>{J7?�ߩ>(���Ѕ��Q�b�NL�>���?�1�?��?�4>�=�N���=�>=	?���?hő?@os?w<?��b�>*�;� > ͗�ں�==@>�i�=	;�=xt?C�
?��
?*����	�.m�w�񾧀^�?��<{ʠ=�R�> o�>�Vr>��=<�f=|��=�!\>m��>v��>�Ke>3A�>�Z�>�d8�MgϾѹ�>�<|����>w�g?!��>}m�=/�D��2�=^3T�-��<�̺=�!>�����"{��oG����<�7�<=v�>Ɇѿݗ�?Ӏ<�����5?�o1��G=1$�>Z0�>Ί��]��>�.)<"2�>�rd>�a�>��>��>4��=�FӾ�>���xd!��,C�p�R���Ѿ}z>֜��h	&�Ɵ�zx���BI��n���g��j�M.��g<=�˽<#H�?�����k���)�������?�[�>�6?pڌ��	��F�>���>�Ǎ>�J��D���Rȍ�hᾠ�?.��?3 �>���>��K?��>��n��E�� �A��h��{]�|f�Ԩo�XԆ��G�R���H�=�Lw?�,�?3,{?��>Qh>_>z?�8������>�X1���@�@���=(��>�ɽ���ў�?�����>aa?id?[��>��w�v5r�7>�i:?��2?��w?h�1?��7?|��t�(?�*>�
?��?�M4?m�-?�G?l/>ޚ�=V�P��E=�������coս0
̽�Ǽ��U=��_=�O�o�;��<�6�<�/켘!��(�;������<��I=��=�e�=A��>�c?��>��<i�:?C��W�b��<5����>������PLξ1�j�\��k��<��?ٸ?jh?K)>�� �E���!>�U�>1�G>�� >� �='<>3�
=��>\�]=z�>b��[�K�������9��
2=g+�;@��>{�>��սO� >sâ�%u��u>��T�UM���Z��ZF�0*/���h�G�> �I?C?h��=��ؾӍM��Of�~�-?58?_sK?U ?���=�Ѿ03��\I�e�S�>�K;�f��֢�B��Ð9��U��'�e>�����ּ���;>������X/k�/YK�?���n=EB�ؓ�<%� �C�Ǿ&F��ˌ
>��>�����+�����5����E?Y,=����,6p��sþ/��=]��>�W�>��Q��C���:�8����� =�\�>DL>΀��.�2�D�q�`e�>*cE?@`?x��?�o}���p��D��V�DD��n���z:?�>6�	?Z�D>D@�=%���>�)2e���F��M�> ��>�6��dG�G����-�$g&��ʅ>�l?2G>��
?-5R?ii?��_?=&?�
?�>��ý�*��F&?Q|�?��=x%ӽ2'T�Ǿ8�<<F����>Y�)?C��l�>��?��?s�&?)FQ?˨?��>	� �L@�Qy�>�$�>k�W����YZ`>dJ?'�>�UY?�Ӄ?�<>��5�̇��!��[�=� >G�2?�F#?�(?�|�>�F�>����G��=p��>�%e?�c�?qUl?(�=�h?�]>(��>�ޕ=�z�>m��>�>?�#N?��r?kN?�o�>؞�<�2�������Ō�X��}�O<Y�<�-J=h}I�����Ƽ� �<ٸɻ�޲�>%��������Bm�:�,=Ec�>�s>���1>�ľMG��I�@>đ���@��vኾ��:����=���>�?���>CA#�fђ=��>G�>����1(?X�??�/';G�b��ھ��K���>7B?��=��l�p�����u��zh=��m?��^?�bW���O�b?��]?=h��=��þx�b����e�O?<�
?0�G���>��~?f�q?W��>
�e�+:n�*��Db���j�(Ѷ=[r�>LX�R�d��?�>o�7?�N�>/�b>%%�=hu۾�w��q��g?��?�?���?+*>��n�Y4���U����I?��> �ƾY�%?��=�aо�I�Q��v�Ay����Ⱦ��k����:*��tu��u��=��?�iv?W��?�6f?��ǾZFh�c�h��Sp�Z�m\�E��E��q*�(	;�U�������T����$������B�mɲ?��?K%�XV�>X���u���NN߾	�g>�x��V�e��=�9=U%�<�U�=���I�?����x�?3�>���>
'?�%T��H��_7��|'�~����O�=�>�̭>ȡ�>U�=���������������"��3w>�hc?��K?�n?�Z ��t0�!�����!�-�A����A>�>��>2T�����%���=�h�r����폾Y�	�Єt=��2?M�>}!�>�&�?�L?����h����x�{�0��?}<G��>�'i?f?�><a�>V*ƽ z ���>%�l?��>�>�����Y!���{��ʽ�&�>�߭>���>M�o>�,�#\��j�����*9�Bs�=֩h?������`�S�>R?��:P�G<�|�>ئv�ѻ!����!�'��>
|?�=o�;>rž�$�N�{��6����0?q�?��u��y�~�>D�(?� ?�,�>��?S��>]Iݾ+Za��?�NI?�[4?&T?W�?�7">��=p�ܽ�o���t=�>dR�>N��=��U>��;�c��	$��#K�ڟ�:h��?�j� -�= ��=�\�=�c=��=|LݿjJ�dẾT���K�S��U�����&��y �����h����[�8���ӏ���x=��g���Ė�5�����?�7�?��ľ���04��1`������>W�F��`��A��V���1�����ɉ�j�0�"A��^��`_���'?鼑���ǿ���Aܾ7 ?�A ?l�y?J���"�{�8�Ҭ >��<[���뾏�����ο������^?@��>F����)�>��>j�X>Q<q>)��螾/ޕ<T�?�-?��>ۇr�`�ɿ7���)��<���?�@I|A?+�(�՟쾑OW=���>��	?)b?>�q1�5+�T���*�>.;�?���?�*N=ǼW�\���te?pE<��F���ܻ���=�n�=��=Т��VJ>�z�>� ���@���ܽ�`4>ׅ>�"��,�9^�5��<��]>�ӽZ)��0Մ?{\�af���/��T���U>��T?�*�>W:�=��,?�7H�n}Ͽկ\��*a?�0�? ��?]�(?�ڿ�3ٚ>r�ܾZ�M?;D6?���>�d&���t����=�<ἶ�����㾻&V�Q��=-��>x�>U�,�	����O�H��y��=N�ȿ|�#�����,�<t�
<V������4���g��V�j�M����=��=%]K>WA�>ݿR>|Y>;W?�ih?��>H#>�o��!��_}ϾT��脾p(���Q
�P��_G�iݾ�/��E�&��âʾvyO�C��.�I��%����<�򉆿t�D�y7>?��`�'���?���<?羮�(�C��=��˽=��Q-��t����?��#?����=	[���6��N����=���?R���0���ľd���&��]�/�J�>�Z��YJ���[��sG�6�3?$?�r��q����>�Ͻ_�=�,?�0?��;���>��?����b��w�:>�L>��>��>v;7>��������K?�YR?V��|���ʘ>�b���4��
�\=_��=^�a�cP~���m>9)=�̄�T���Ӝ��n<�CX?z�>�)��7��Y����	�@Z3=��w?}
?���>O�h?��>?
y�<����[!U�;��#�=[�X?2k?�>��d�CX˾�����1?�vd?��L>[^��a�q�,�����v?R.n?@?�7��x}�����:��4?�v?�o^��r�����"�V��=�>�Z�>���>��9�zi�>�>?�#��F��h����Y4��Þ?G�@��?��<<��譎=^:?S�>k�O�H>ƾ����n}��]�q=?%�>�����gv����Q,��8?��?���>b���W�����=d^��#�?JA�?F�\��"=�?��)l�X��-Sb=}=�(�=�Ì�5SϾ}��������P���粽�φ>9�@sky=���>m;�<,�ѿ mۿ���b�ľz&��3�>J��>V{>v_���2b�)X��5�,�-7M��CԾ-"�>+�>J��n��[�{���;�Q ���,�>���߈>�S�(��u����@7< ��>X��>���>-[�������ę?�P���Cο��������X?;f�?:u�?q?44<�	w�-�{���� G?�s?�Z?y�$��)]�SO8�%�j?�_��wU`���4�tHE��U>�"3?�B�>R�-�a�|=�>���>g>�#/�y�Ŀ�ٶ�<���Z��?��?�o���>r��?ss+?�i�8���[����*�]�+��<A?�2>���H�!�B0=�UҒ���
?U~0?{�e.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?\$�>�?)x�=�a�>f�=M�"I-�f#>E �=9�>�C�?��M?�M�>\�=b�8��/��ZF�HR�($�:�C��>��a?�L?qIb>`���2�*!�/xͽVa1��5��X@�0�,�P�߽�&5>�=>�>��D�d	Ӿ��?Lp�8�ؿ�i��p'��54?.��>�?����t�����;_?Nz�>�6� ,���%���B�_��?�G�?<�?��׾�R̼�>?�>�I�>9�Խ����X�����7>1�B?Y��D��u�o�z�>���?
�@�ծ?gi��	?���P��Ja~�	���7����=��7?�0��z>���>�=�nv�׻��T�s�Ź�>�B�?�{�?%��>�l?��o�C�B���1=RM�>՜k?�s?�\o��󾌲B>~�?"������L��f?�
@|u@`�^?!e����Ix�Ԡ:��l�f�>��=�*#>��.�t�G���f>�&�=�뜽�z>�ɗ>�� >���>��=�<>�}�=N�}�\��op�-���dQ/��z-��	9����T���ꃾ��F�>��g��98>��!����<�]��&���6��U+�=��U?�R?pp?� ?=�w��>����G�=�E#�y��=BO�>$w2?}�L?)y*?�+�=j�����d��T��� ���ć��b�>ΎI>�f�>Y�>��>��9d�I>~5?>��>H� >G^&=�r��i�=�O>�'�>O��>ǎ�>y >��;�Cÿ	��cg��hp�6 W����?7N̾�{������~��7)�)B��(�>?g^�;<o��j�����7;??��l��[	�V�(���=��.?�K?T��=������� ���6W�;�2����<n���Z���3����=�I�>�"g>J�4>��G��@H��Fa��־O[�>�C?��Ӿ�f��1���F4��e��
>uo�>�(��E�"�SO��\ˆ��T��ԏ=�O@?�?G�����qt�����&.>1g�>�>x=\�n=7��>. =;��8���d��`=�^=�M�>(�?�/>��=Lܢ>Q����M�4A�>�@D>��1>�c??�$?*!�U������(�/�fy>�s�>O�>�{
>�&J�C�=W~�>!b>��dK��/V���>��V>/�{�M`��Ń���|=����R�=\�=#{ �?>=�p!=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ,h�>�x�tZ�������u�6�#=(��>�8H?�V����O�_>��v
?�?_�����ȿ.|v����>:�?���?8�m�iA���@���>C��?xgY?�ni>�g۾�_Z�:��>��@?�R?��>�9�f�'���?߶?⯅?߶G>�^�?���?���>=�p<Z��Ѵ�GД�t,O=ss=oQ�=�G�>8���=�0�������K�*�.�XǶ=��=�o�>F�e�N�������������WY���R�>)��>�ak>��O>�:�>z��>%�">w�=L���	:��X�4�v�K?o��?����1n��Y�<���=�^�9&?�I4?�[���Ͼ�֨>�\?I?V[?Yd�>����=���翿�}�����<�K>:5�>�H�>g&��"IK>(�Ծ93D��n�>�Η>�����?ھ^.���C�>�e!?��>�Ү=ۙ ?��#?��j>�(�>BaE��9��Y�E����>آ�>�H?�~?��?�Թ��Z3�����桿��[�o;N>��x?V?rʕ>b�������rkE�3BI�7���^��?�tg?vS�/?;2�?�??^�A?|)f>Ӈ�'ؾc�����>6�!?���A��M&�i��|?�P?!��>
��>�ս��ּ���D}����?�$\?XA&?ۖ�_$a���¾�&�<	�#���S�D��;�C���>�>P��� a�=�>W��=�Ym��=6�;�g<~�=��>��=!-7�I����=,?��G�nۃ�v�=��r��vD���>�JL>P����^?�n=��{����{x��y
U�!�?��?sk�?N���P�h�h$=?��?M?� �>�I��/}޾��ྱLw��yx��v���>���>}�l��B���s���FF����Ž)6��ˈ�>�N�>���>�d?Y\h>׳�>�}��P�x8�������Z��%��dL���(�|� �&�h���s�����ƾ_R���y�>I���0�>�k!?Q��>�Ij>w��>) �=T�>�+>=�{>�?�>�>�>�U>�`'>S�'��7��KR?�����'�>�辇���`3B?�qd?B1�>�i�5������m�?���?Bs�?=v>�~h��,+��n?�>�>?��7q
?�S:=@0��>�<�U������2��	���>�E׽� :��M�}nf��j
?�/? ��>�̾�;׽K�����n=M�?��(?f�)�2�Q�}�o�@�W��S���z!h��d����$��p��돿n]���%��p�(�?D*=�*?��?h��B��F ���%k�n?�]hf>��>=�>e�>&wI>S�	�!�1���]�4N'�ഃ�4P�>@X{?!r�>��A?�9$?pU~?An[?�X�>"m�>dC���%�>��%�.>�?56?�>?*�C?��?d� ??3�>wxt�Ոݾ����iy�>�n(?G<?,o�>�B?�U��'=�׍���=�ǎ�mA�� 0���>�����Լ@e>
!�>P\?�t�$�8�U�����j>��7?�z�>R��>����Z-��!�<��>��
?�<�>� ��rr��X�$_�>���?F�xt=�)>(�=������˺Av�=����.ߐ=D��u�;���<|��=��=W�o������"�:�}�;��<Ez
?8�&?��g>)�c>��m��9�l�����=�@�>��B>�
>7T;�q�����ȶm�!�>tӓ?�ҳ?.�>,�>*6>����V0�+�Js���m���?9�=?�dR?�ɇ?��?��"?6�	>����Ñ���{�vF��;�?,�?q�->EJ�����⡿�Y��K?_?�{r���8��%������-o���g=��9��:�����׉H��5
���	��A��?���?�>E>s��������i��&.X?x3?e�2>	j?�6��}�������]>�x�>�?�0�>=�W?�"�?G�9?�S>��ɾYW�����d=c��Os>h�?��p?�͐?���?,)=?�׼UH��O)���� ��<�@�Ȼ��']>RS>5�>��>w%�>F�P>��{���p�.�����;b{>��>��?�F�>L��>q9�=�$J?e��>쨾����c���Ӿ�=	�j?C��?HO ?��Խ�<�*)����'w�>su�?���?� ;?���=����,���?]����>��>�+�>��������w>�#�>��>~�[��Ɋ������j?��>?�`�=�dƿ�s��y��G����<h�j�&["�b�ý�9:���2>U[l���(������H�"�_��ˎ�Ӭ��xt���v����>}���&�=[!�=��*��3��<;5=��<ri�<!�5�p�c=Mi���mE=fz���ռ������<Kk��B�˾$�}?�:I?��+?��C?��y>G9>��3�T��>����>?eV>^�P�㉼��z;����������ؾ�s׾��c�>ɟ�SG>B_I�$�>�<3>�N�=p$�<t
�==s=�؎=ȔR�p =�&�=(P�=h�=���=�>�c>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�??ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��B����4�?��@��??�ዿТϿ6a/>�m7>��>݈S��#2��7a��Qe�InX�5G"?%k;���;� �>=��=_Z�w�Ǿ�~8=e�3><�X=�T���\���=ҝz�*i>=Y5l=t�>a+D>�k�=9���z��=�R=8u�=�Q>Mq���2�-l0�ZN(=�0�=�a`>��$>B\�>|�?�e
?wb?��>��Ͻ^����͸����>-Ί�Dk�>��o>6�9>؇W>S�?�z\?��T?��?�X�>Yo�>��>U�*��߁�s�������<9G�?Ԡ�?�:�>?����_��(�+-9���W��a?g3=?D5�>M	�>�����޿�)���0��`�����<�̜=�t�f��xߛ<����l��w�=>��>���>uǓ>x�z>ΰ->��L>lI�>��=�ʀ<?x�=�w��M=<�7�69=B�+���%=�D��M�<�(9����@��d������;�<���<���=8��>t9><��>g��=�	��:A/>Զ���L��ÿ=$:���+B��3d��J~��	/��^6�<�B>�9X>�z��]4��h�?��Y>q?>,��?�Eu?��>y)�ͺվ
O��18e�SS��ʸ=�>�<��x;��S`�:�M��uҾ��>��q>-9�>��5>�s���G��0=��¾	�C����>Hz���t���@4�''z�;㭿����k\_�נC���4?H��� >{2v?��I?TD�?��?X�����Iw>��!�+%>����~J�@���?�3?�|?D��A~�<L̾�*����>�VI�M�O�ۿ���0��G�$�����>=U����оj 3��n�����)�B��Tr��޺>"�O?�ͮ?X�a�CB��o(O���Dp���w?Cg?2Q�>�V?�S?����Z����]��=�n?ż�?=�?��>$g�=��P���>"?p�?��?��f?'s=�gw�>`/(�(L]>�.2�Bù=��=�;K>�=�	?��?��?Bp���D�C'�L
���{���=Ü�=��Q>_p>��R>���=Q�=M=�KO>�͔>.��>� �>���>�*�>�tվ	#/�FM�>-G=/�?>��:?���>q�m<�&4=�r>�]<�j�L�V����0"��#Ib��4=���<��";� �>��¿���?g3�>/+�c?�;�A��>D>WI0>PȽ��>i��=Yk�>Ulw>N�>E#\=a\>��>�EӾ�q>���e!�1+C���R�j�Ѿ�z>ި��D
&��������JI�p��l��j�K.��y;=�Dr�<D�?Ǥ����k���)�c�����?2V�>�6?Gӌ��2�>���>Rȍ>�P������ō�CV���?/��?c=c>�>��W?ݚ?�1��3�]uZ���u��'A��e�ջ`�	፿ʜ��'�
��	����_?d�x?�yA?]n�<�:z>N��?��%�bՏ�(�>�/��&;�5J<=�-�>e(��<�`��ӾԹþ�7��EF>��o?'%�?�X?�SV�N�L�V#.>
49?]#7?s%v?��1?�~9?�����"?z�(>^�?�?��3?1+?��?2>�p�=�!<��O=	��������н��˽�мT�M=ω�=����i�8�-�==$dݼ���u�;n)���<�mL=0��=x��=�"�>E�^?Y��>�94>Cd,?<���V4[���N?�2=�����U�L��T��\�=[�|?�߮?�0m?��>?41�I�D��
.>��>�Q7>���>.z�>G��zm�8>��=^�<y��=˲-�����h�Ȋ����6<^�="��>0|>�����'>�{���/z�ަd>��Q�t̺���S���G�/�1��v�Y�>�K?��?=4^龆*��XIf��/)?�]<?�NM?��?��=U�۾��9��J�n<�-�>d�<��������#����:���:��s>�1��V����A:>�!�d����|�9�E��Aؾ_�%>>�3���Su��ڨ�M����U�=�f>t�о�p�@���!��CLF?6a?=���"aE��6��x�,>Y��>2�>&ª�^p�T�C�����S�=�W�>�>ں������!O�/* ��:�>�OE?LX_?9k�?����	s��B�����g���pǼ��?�|�>�j?�B>!ѭ=Ҟ��6�1�d�DG���>��>�����G��7��D*����$����>9?Ɲ>�?P�R?�
?��`?*?�C?�'�>x���������&?X��?��=��ӽm�S��M8�|�E�G=�>� *?�sC��ݗ>�?+]?�J%?��P?�Y?O2>���o�>�-��>��>�jX����\�]>Q�J?�9�>�+Z?TL�?,�7>�4��`����1�=q�>��2?v�#?�?�Y�>���>x��8�|=�v�>�\?�&�?�q?�2�=�V?B�R>��>��5=���>���>;?��O?��l?}0K?���>��={����%���(V�S���D��3����=Ud�O��L}�J#=�$=�'^�ʶ�����<`�������2=z_�>K�s>���W�0>A�ľ"N���@>դ��LP���׊�_�:��ڷ=T��>x�?���>�S#�b��=u��>'J�>n��<6(?f�?�?<�!;P�b�&�ھ�K���>WB?F��="�l�ゔ��u�ch=��m?6�^?:�W�x#��O�b?��]?@h��=��þz�b����g�O?=�
?3�G���>��~?f�q?U��>�e�+:n�*��Db���j�&Ѷ=\r�>LX�S�d��?�>o�7?�N�>/�b>'%�=iu۾�w��q��h?��?�?���?+*>��n�Z4����������\?#�>l��8h#?�c�bϾ����������!���Ŭ�8������p#����oyԽ���=3�?��p?.�q?8`?]� ��Pd��_�(����U��� ���e�B�IFB�_B���m�~��7����K��8�L=�$���j���?S�%?O�]���>��T����M����v�>��'2��S%=�u뽉C�=��f=�3Y�ez�#a���U"?���>4�>��A?��G��AE�<H��F��F �>�f>Ӝ�>�[�>�c�>
*8=�t_�����>Ͼ󝟾�����CK>�
X?N|G?+w?�]�<r�.�4Ɖ�:D(����|��d�>��`>�,�>��������%��3�ʦ[����yLc���?�Ȕ+?�Ts>~Q�>#��?��?�ɽ�}����)�.7�N�1���>���?E�?�)i>��=ݮ�D��>Z�l?���>��>����`]!�(�{��ʽ*�>��>���>Ip>�,��%\�Nn��]����9��:�=1�h?;{����`��ׅ>IR?h��:�dG<�t�>^v�:�!�y��-�'���>Hv?*t�=��;>�tž�!���{�d6��I�H?G@)?�4˾��+��o�>
UQ?���>� �>�e�?ҋ��S־�@��_^0?OrK?(	?{�q?�7=?S��>�黰����!^��B>t��>~
�>W�>oJ7>�~��o�-"��z���
V="&�B6>
 �=�(=,��=O9�<�z�<2mۿGCK�{�پ�
�m��?
��戾����b��&��c������[x������&��V�
8c�����w�l�e��?Z<�?ǂ���1��z������0������>�q�$��h���	���+��~��b����d!���O�%'i���e�:�'?����ݽǿ𰡿�:ܾ! ?�A ?8�y?���"���8��� >�@�<-����뾩����οu�����^?j��>��.��x��>���>�X>xHq>����螾�1�<��?�-?0��>!�r�)�ɿX���[��<���?/�@e}A?��(���|V=���>Α	?��?>R1�(H�����T�>D;�?���?yM=�W���	�f�e?�<\�F�|�ݻ��=�<�=@J=���@�J>$U�>���TA��?ܽv�4>�م>7u"�1���^�7��<Έ]>�ս<��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=v6�����{���&V�}��=[��>c�>,������O��I��V��=����uǿ:�#���i�<���;��4�M2�'���@�@��4��pns�����pP=	#�=3P>�L�>mqV>�Z>��W?�xh?�g�>�_>���4���0}оB�y�PĂ�v��ĉ�f�$��`Y쾊�޾m	�M�ַ��;Ǿ_fY�n�G�߾@�9~���A�\���Z�/�HX=?>�:��(P��y�>S�
�j�c<���=?�F�,���� ��H��ѵn?��?����k���E��A�u6ӽ��?�"������\F¾r��=B���G1����>���j現�nR���w�\�0?̔?��������K+>vF���I= �+?��?{�3<}��>2H$?z�(�m��!�Y>�6>��>L��>��
>oƮ�(ܽ%a?^]T?���.图��>�_��Z�{���]=݀>�p5��(༏]>�5�<�B���sG������Я<X�Z?q�>Ψ-�8� �>�� �6��W=��u?��?��>�f?�1??U+=�����uS�������=�\?,m?��>up���Ѿ�6���8?�i?k�]>5X�cv� �/��z��?��o?�?��ļWt�
f���-���+?>�v?�]^��a��r����V�&��>+��>.��>{q9�tس>A�>?�#��$������EO4�_��?��@�{�?r�Q<��k��=�%?.5�>e�O��Mƾۨ�������p=���>툧�A1v��|�a+��s8?�ƃ?��>�����r������ ��j�?�/�?�j��Ϲ�<f��z������=��>&��v�=W$ܾ��;��Fɾ�
����c�<j�>[Q@\��<��>I==��Ϳ�пw���G��$���L<?}��>z��=� ��򊁿����0D��iI����kJ�>��>����������{�nq;��2����>����>t�S�� �������5< �>-��>��>�+��K齾Eę?�`���?ο��������X?jg�?�n�?o?&9<p�v���{��7�#*G?�s?�Z?Q%� ;]�b�7�<�j?;l��HM`�A�4��;E��dU>�?3?)V�>e-���~=`>6?�>�`>#/���Ŀ�ɶ�;������?^��?�M�=��>�t�?�d+?�d��2���s��S�*��5�g,A?:�1>$x����!�=�麒�e�
?�}0?���4�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?L$�>��?`o�=�a�>d�=\��-��k#>,"�=U�>��?��M?L�>
W�=��8��/�G[F��GR�S$�<�C��>��a?�L?�Kb>�� 2��!��uͽ�c1�P鼭W@�!�,�ޞ߽2(5>��=>�>>�D��ӾP�?Up���ؿ�i���o'�64?���>k�?��o�t�ڐ��9_?�y�>)7��+��Z%���@�I��?�G�?"�?��׾�T̼�>��>H�>Hսk ��������7>"�B?X��C����o�X�>e��?��@ծ?i��	?
 �UP��`~�H��|�6�,��=6�7?3*���z>���>@�=�mv������s���>�A�?){�?���>e�l?�o�_�B���1=J�>I�k?�q?�p�q�@�B>�?������I��f?@�
@�t@��^?�좿I��燿7,��P����T>�o�=��Z>Qǽ�
>&�<��q<'QX=1��=a�>aBA>5Y>�[->Ui>��@>��\b��a���i����`���E����v��y{ﾝ���os)��M��v� �$=p���r��#��N����t��
�=vU?�Q?�Sp?�� ?JJw�@>5�����=��$���=��>� 2?P�L?�-+?�3�=_֝��d�?��u���������>��I>���>dK�>n�>Ŝn9��H>h[?>� �>e;�=�"=�@�:b�=_ZQ>���>K��>���>z>�֢=V���o�����X���p����?y�þbRK�Pu��:������=�3E?x�K;��}�n�ȿ���f=?�·�U�?X�5>�h"?�jP?P�=h�ƾ%��=�<�EO�˻{�7IO>��-�[d��55�2��<Jq ?�,>�j.>@<�2G�2�c�wTܾ�q�>�GH?a� ��\��1e����.���l�>���>.ͽ�@0�� ��IQ��Ýy��=�0W?��>{G�.ڵ�v�M�`��Ԑ�='��>���=�#�T2�>�$���|7���F���݄�=T!�>vp	?�m>M:f= ��>&ӕ�+9!�N|�>H�N>��R>quH?d?'?�*����J�� J1��w>�t�>{��>��=>r�2���=ĺ�>J�V>9�G9��1X(�y�S���O>��t�i�f�W�I�l�=O���=�>�t½��<�
Ӆ=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾQh�>~x��Z�������u���#=W��>�8H?�V����O�_>��v
?�?�^�ߩ����ȿ3|v����>X�?���?f�m��A���@����>9��?�gY?qoi>�g۾7`Z����>ѻ@?�R?�>�9�o�'���?�޶?֯�?%A�=�ɏ?gӉ?+��>~7�=3�����4���*ν\�(>�\�>�>gނ�Q�L��W���a���P�g��d>B�=���>��1	>��r�=
e������=��>p�?>�m>.��>�v�>*U>��>D�M;^��H��$g���K?���?-���2n��N�<Z��=)�^��&?�I4? k[�}�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��H��<��K>*4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��WS��GB�>�e!?���>�Ү=ڙ ?��#?��j>�(�>@aE��9��X�E����>آ�>�H?�~?��?�Թ��Z3�����桿��[�q;N>��x?V?qʕ>b��������kE�1BI�/���]��?�tg?uS�/?;2�?�??_�A?�)f>͇�'ؾf�����>�"?�
���A��?&�N�Z�?�?;V�>s܌��
Ͻ��ȼ�7������r?�[?��%?
�I-`�q���=[�<�_ �ZH����;*J��>�n>�/����=�>D�=��l��3�X�<��=��>"��=OE7��F��0=,?��G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?a��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>�l���K���ڙ���F��`�Ž$w9�"��>�1�>&�?:��>5�6>e�>.Ð�(��������`�v����6�Y�,�0�T��+4�����Y̾��t�/D�>��5����>}?��s>�-g>���>wG�5��>kO >Ҕ�>&~�>�H>ǂ7>j�6>��z=\���LR?�����'�c��O����3B?rd?G1�>�i��������?���?,s�?�<v>�~h�n,+��n?,?�>��#q
?�U:=�3��:�<&V��ս��4����E��>(D׽� :�PM��mf�rj
?�/?�����̾�8׽���异=vڅ?x(?��&��}P��Kp�5�Y�u�R�fW��^�V���=�!���o�+_���L���ރ�F�(�D�)=�)?�^�?7� ��2ﾴ����8j���?���^>�7�>�Γ>x�>��Q>l���1��_�ݝ*�����Np�>��x?B_�>�E?Kp4??N?(VU?�`�>�B�>�K��n��>��@�P��>��>��:?L/4?�W0?j#?��0?�J�>�⦽�P��`��o�?��?��?��>�?�8���#���=��2=�f�4�ƽ���<�l=�ج���ܽ�X=��>��?�3��x8�����5�i>��7?���>:��>����p{�\, =~��>EF
?�{�>|����q�fY�h��>���?���M�=x')>}��=�؎�ŀ��^�=�2ؼO��=	N��!�?���$<$�=�`�=(�4�6p<~�;�~b;P5�<u�>?�?���>�C�>�@��� �X��9f�=$Y>S>�> Fپ�}���$��q�g�^y>�w�?�z�?J�f=��="��=#}���U����������<��?AJ#?	XT?V��?Q�=?\j#?Ƶ>+�^M���^�������?�l?n	v>�?�#쾰����C���?
G?��|�J�>��+����T�N1>@,���x�Aj��h�Y��ϕ�9
���	����?-��?��=�#�|n羬��(ܑ���7?3~ ?w�Q>v�?�m=�c�e�="����=�O?V�l?�~�>��N?�y?��\?�]>m�7����^���j`�� >��A?H��?^��?st?P��>ݠ>�R-���޾���q���� ����vm=Y>�o�>�o�>*�>{�=�]ؽ��9�D���=�m>6?�>as�>zt�>d*�>�I�<�CX?ME?O侧�������r��Rg?Ls�?���>���=�#�8k�<4� �>>v�?目?�4??�����%�=���;i#ҾY���>���>��>1b>��=���<���>m_,>��0�oG�j�6��u�x�?ǨR?��_=�kƿ��r�eq�8���TSr<����M�V�7A���+R�'X�=I9��Y��S��:o\�ٹ���z��]Ҵ�Қ�Oy�#o ?��O=XS�=>��=�g<��鼒�<�<=��<T�H=���N�<N�;���f��?���Aܻ��2<�B=���|�˾�}?_?I? �+?�C?�y>�	>�4� ��>f���E?+V>�7P�押�[�;�����>"��9�ؾan׾_�c�ʟ�[B>0!I���>(3>�,�=YȈ<��=js=6Ɏ=qN��=J�=�J�=�r�=���=�>�T>�6w?W�������4Q��Z罦�:?�8�>{{�=�ƾt@?��>>�2������yb��-?���?�T�?@�?#ti��d�>J���㎽�q�=M����=2>S��=��2�O��>��J>���K������4�?��@��??�ዿ͢Ͽ>a/>�6>y�>�wS���1�y�`��!c���Y�sY"?kQ;�r-;ǂ�>TK�=��྾xƾ-�>=��3>u�c=�~�']����=��{�7�6=�2l=H��>&E>[q�=aQ��ǋ�=aP=���=r�M>	����J.��_0���0=��=6�^>Z�$>�m?b?�l? 	m?�Ѭ>�#6����ؾ�=�>��+>3�>��=�\�>ICY>��9?reP?��>?ͺ�>�:H>q��>��>��<�깏���޾|Z��Ϧ�� �?�?��=�M<�re�"�(��7D�A\d��?��`?-�?��>!U�!���V&��.�k���Õ=8pp+=Mir�`U������s������=i�>���>��>�Ny>.�9>��N>%$�>��>ځ�<���=)D��#W�<]��"��=ѽ��k�<G�ż1wz��d%���+��z����;��;�C]<2u�;R��=���>�@>���>a��=�
��s@/>f����L�|̿=cI���,B��3d��H~�u/�A\6�&�B>�/X>,w��G4����?��Y>{s?>���?�Bu?Y�>�&�Y�վ�Q���0e��cS��Ը=k�>� =�#y;��T`���M�wҾr��>^|�>4��>>�*>�-��3C�~q,=�2þ��>�D��>"���佽1��j��ڜ�k���tt������><?�'���`�=�t?'yK?pȓ?���>�eN����	�>C���>�~&��E8��(��К?2�?N}?6�����*�b�ξQ���O��>`kK���O�h|��0�����r˸���>c����Ҿ��2�
���Xy��L�B���w���>�+O?�2�?��`�⛀���L����*zb�"�?-�e?5ʦ>>�?��?�T��Ԃ�â��-�=��m?k8�? ��?�t>��>�����> �>���?�V�?D �?�}����?�}�=�I`>��!����=cЌ=�0J=�{�=��?��?�?��K���������%���ת��D=E�~>�;�>+-�>�=`W�=��>s�m>ج�>���>+�>E��>��>����`�5���
?:
�=Ʃu>�yF?��>��P=�U�<�O�;��?����o�C�$�k�=�(��<e<���|=�Ni7��?g;ɿF��?��>���~�>�z��Cxؽ�2(>��>���V;?r�8>���=�@�>܋l>�p�=��W>�mM>A{ӾSj>
���u!�L9C� �R�z�Ѿ��z>n����$����c����I�ə���S��j�L��:a=��k�<$��?C����@k�I|)�Jv����?-�>��5?曋�s��K�>���>�&�>kw��~��ש�����H-�?N��?V<c>��>�W?�?��1�3��uZ��u�(A�e��`�m፿񜁿�
���>�_?�x?.yA?0X�<a:z>S��?�%� ԏ��)�>�/�';��D<=,�>�*����`�ׯӾ��þi8��GF>�o?G%�?�Y?�SV��7��E��=~�'?#�Z?�@j?��#?G+?����,�>g:>`�"?U�>z�$??".?/ ?�W|>$�C<���=י=HK;���%�_��;�$���4	>��k>����*��gik> B��eE��ƨ=7I^�t��è1>!�1=T��=�m->�`�>D^?%�>9/u>�\<?/Ͻ�,�._��A=2?�6������O��������޾7��=X�r?q��?'�`?��w>��A��P�x�,>�Œ>C>>SEc>��>cc�$qV�[�=�>H�>w�=b�)�ڧg�����䑾Y'�<�9*>]��>x/|>w����'>L}���4z��d>��Q�aк�8�S���G���1���v�YW�>��K?��?��=�`龉(���If�6/)?L^<?�NM?2�?��=��۾K�9���J��?���>��<�������#����:�(��:^�s> +���� ��y�=4潷����(���q�ף����W�H�����̣�ʧz<'��p	?D��=��Ծ�'8�����&ʴ�|<?�&�<;���è����ܾ���=�>oN�>��?��&6�̨<�0Q��
�����>�J�=��>�n0��*��a���>.(A?��]?�l�?�X;��g��9�t��/u��̉ͽU�?$x�>#?��V>�	>K�������V���=�~��>2?�>���G�A�
P��m���%����>���>*=�L?��M?^X?��Q?͍ ?Xt�>*�>Q��(Թ��g(?�`�?>�?=��ɽv�=��4���F�x��>A�0?�H�'�>��?'�&?��?�8I?l!?-G3>����6�d�>2��>�_�F��0;>�L?h��>�T?ӑ�?.�Z>��7�|����P��=���=�|-?U+?� ?�}�>�� ?��<�UX����>�QN?Ɍl?-�?��>
i�>���>�'?�+�+�
>�f=h�>3�(?��>??�^?��?a�=���%�����<s�=0�Ȃ�y)=��W=M~�=�����+�=ƾ':�Q�<t���M�
Z��Ⴝ���_�>��s>1����0>��ľ)M��$�@>����+O��vي��:��ڷ=��>�?6��>#R#����=�>pJ�>W���5(?y�??�� ;��b���ھR�K���>�B?y��=W�l�����$�u��h=��m?��^?`�W��&��N�b?��]?Ah��=�
�þ��b����g�O?=�
?6�G���>��~?b�q?U��>��e�*:n�*��Db��j�2Ѷ=\r�>NX�R�d��?�>p�7?�N�>7�b>4%�=ku۾�w��q��h?��?�?���?+*>��n�Y4�3�ؾZח���C?G��>Ⱦ"�?�ׄ<�j�U('��H���"Ⱦ�y�����ޏ��u���-J�� �������=]!
?�l�?_�l?�i?9���ڀ]��j�4���t�a�E�!�[\�h�0��uQ�g�>�F�}��e��叾ŉ����߾Q�3�FV�?d�(?���"��>d�Ǿ�� ��E�:��=K!�������<1��=Z�"=^;8j���i�����ӧ?�.�> 1�>Q8)?j)M��xF���0���+�Zi����F>���>��>��>$(!<P4+��7�bU��C#������ s>�g?X�W?{i?5\���oO���|:�\�Ӽ�qz��0c>�h5>��>�R ���5�T>"��+��q�f�
��ӂ� &�;�H��|>?i�1>�ܔ>ZR�?
w?fd��%�������d0�x�<��>{y?Y�%?���>Ó𼷿!�ײ�>�l?��>��>n���R!�O�{��H˽��>R�>��>Y�o>��,��\��m��愎��9��,�=�h?�|����`��܅>TR?QS�:8VF<�~�>�6v�N�!����\�'��	>�{?�\�=ʬ;>Xnž>�W�{��J����6?-k,?���w}T�� �>�>?��>0��>�?%��>���{ �O& ?H�<?u�>?�-n?��N?I-�>��F>a��P`��v�Y>{H�>2�v>��|>m�>8�s��"���{�k`�i�=0��,x��'��>���=f#�=C^R>� >�H�`E��k���p��^�о4��`ә����~둾�w:�9������2���4��EH�2�r�c�~����{���!��?x�?�"��I�s���Z�B����>��n��U��֛� u����)�������h��;���v��}���-?���{2ǿr�����B����>p�?�H�?@%���h`�p�#%>/��T�>�a7�������CƿA0¾�C0?#(�>G7ɾ�z�<p.�>G-�>=��=���=~Ǹ�v�����>p?��?��?�����4ֿZ�Ϳ���x��?�@�/A?Fk/�l������=���>Q�?��i>/����E���5�>e^�?�Z�?�$=�,T�^����b?���<B�;�jF<�I�=xx�=��|=��+�8�>`��>4����8�V����>}��>�kὦ5ӽH�J�T����>����н�Ԅ?�v\��f�&�/�PR���g>��T?:)�>30�=s�,?�9H�k}Ͽ�\�(a?�0�?���?��(?�˿��ݚ>J�ܾ��M?&F6?���>�a&���t����=Ξἱu������V���=���>�r>ׂ,����[�O������=���r�ƿW�$��>�^� =�B��U�W�Ǒ����@pO�4����n�/�轙qg=0�=IiQ>�c�>KaW>RsZ>�RW?G�k?4�>�>�B鉾Q�;}q��n��*���ǋ�ZB��������5߾Kz	��������Aʾ�2����=�C�5ꏿ�$9�E�y��tD�	3?w��=�]̾��T����=�
	��
����y=}ϽȜ�!�<��z���?N�G?�<��b�!�2��.c�u�D=[�v?�7�;δ	��T��ݼ���� U�<���>��=s`����#�F�[��t0?sT?�t��9w���*>!k��7e=S�+?wt?�\<�h�>�$?�*�A���4\>�5>���>�n�>Jg
>"���.ܽc�?��T?h�h���ߐ>����{��Ta=!]>4���９�Z>�<,ь���c�4揽�C�<��T?*�~>�+��{��?y���{��Ώ=�x?_�?Qߞ>��m?_%<?d�^<&�����U�����=�X?7h?3G>�-��Y�Ӿxʠ��3?�$]?A@>��b��,1��.���?��k?+K?Q��ղy�����>� �5?O�v?tz^��q�������V�i>�>4u�>��>6�9��o�>��>?N�"�lC��˳���T4�_��?ǐ@L��?V><c����=�2?�f�>��O��ZƾZ��Km����q=K
�>�����Ov���{,�B�8?a��?M[�>�������4�=S�f�hɟ?y�?�����B<R�Hz���`�=��<q:�=�T<�Y��Z�@��Fʾ�6��𰾏ɱ���D>�@__g=s��><0L�	MͿ�"ҿ7��������C?��> �g< y�9^�g�z��U���g��2��x9�>��$>�]h������B�U�%����8�>����Sf>苾4SX�-辪W=6��>�@�>�^>�U2����2�?{���#ڿ�c��%=/�c<J?�ѣ?�?l4?�yI��������sw���7?��?-h=?*=J7<�Ž���j?K~���X`���4�'hE��Q>˞2?Ǥ�>��-���x=r>���>�>:�/��Ŀ2��`���cĦ?[�?Ӽ�w��>��?�+?+�5˙��g����*�)5j���A?��4>jT����!�==�+���2�
?�_0?�+����]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?}!�>��?���=�d�>bi�=BﰾZ�-��P#>M�=?���?\�M?bP�>\�=�8��/�=ZF�!GR�q#���C���>m�a?�|L?~Qb>M��Hi2��!��ͽ5d1����qW@��3,��z߽�5>�=>�>��D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>D�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?�Qo���i�B>��?"������L��f?�
@u@a�^?*e޿`y��I����w�`==p�=?94>��� �<�#��C�X<��ؽ�/�=��i>5�p>ʴ�>9E9>C�l>�1>LP����#��������~x]�o]�4��z97�\������:	�]}��pŨ����	C�Z���C�'-���O�����=IqT?�zQ?R�r?���>PTr��Y>FW��ڠ�<'�"�R�=O�>�O5?�J?�X+?�ҧ=����a�p���ǣ�q��~�>��I>J;�>�d�>�׬>�q�<zB>��/>��~>��=aVK=�a˻{8=M�Y>pj�>��>
l�>��q>[7f>م��?���� �������!���?�;��`W�������A�y~�]�/>fU?C/�=�|����̿k췿@yE?o�zF!��n6��(=�^N?��Y?`)>�^��4:�~�#<X
[�YP��%�=)�l��\�����|>��'?��f>B$u>x�3��g8�6�P��u���x|>�66?�޶��S9���u�ܴH��gݾ&?M>C��>f�D�"k�����d��ui�a�{=ht:?z�?�7��Zٰ�Şu��B���ZR>�7\>~=�c�=�rM>�rc�.�ƽ�H�<[.=���=��^>�	?o��=��<�9�>�S����:�(A�>z�O>B�;>[�:?�I'?}|9�)��v�Z�-���k>%��>e:�>V>h���=���>C}>�����
�o?Խ��I>Q圽iNy�e۹�-Y#�t#*;��>|.�<v�H�&��^u��~?���(䈿��e���lD?T+?a �=3�F<��"�D ���H��F�?r�@m�?��	�ߢV�@�?�@�?��K��=}�>׫>�ξ�L��?��Ž5Ǣ�ǔ	�2)#�iS�?��?��/�Yʋ�<l�6>�^%?��ӾQh�>qx��Z�������u�,�#=N��>�8H?�V����O�w>��v
?�?�^�ᩤ���ȿ7|v����>V�?���?f�m��A���@����>8��?�gY?boi>�g۾`Z����>ѻ@?�R?�>�9�}�'���?�޶?կ�?$�>`��?��?�{>Yj����J����!��Mx��lFw>��>�p�=�u�TkҾ�U����)x`��-1��mq>�G=a��>zL�=�^��:��=RE�r�پ�غ�]�f>-E�>Xx�>S��>wF?w6�>�S=j���&�=a�h�߃ �}�K?���? ���2n�iN�<p��=:�^��&?�I4?h[�t�Ͼ�ը>�\?f?�[?d�>3��L>��A迿3~��8��<V�K>54�>�H�>�$���FK>��Ծ�4D�dp�>�ϗ>�����?ھ�,���N��rB�>�e!?���>�Ү=ۙ ?��#?��j>�(�>BaE��9��X�E����>آ�>�H?�~?��?�Թ��Z3�����桿��[�s;N>��x?V?rʕ>a�������~kE�>BI�:���^��?�tg?pS�0?<2�?�??_�A?{)f>ׇ�(ؾq�����>?$?;�:���C����PD�z?0�?�[�>��d���˽ 1Ż���ܱ ��?pX?0 !?6�YY�,��`=��)�N���)C<���8>�9>�7��A��=
�,>_ut=��f���0�߰U=%x�=���>͸�=�;�f���<,?�H�oك�,�=��r��iD���>?L>����է^?.s=���{�k���v��e�T�8�?`��? m�?�ô�=�h��=?1�?@?�>�M���u޾���Jw�tx��h��>���>%n���������OD����Ž�:W�`�?���>�T�>���>��>���>X�	�.��5���������*�68�0�6���&������=_��ڇ<t.վ�|U���>�Q��A�>�B?�K�>-�g>$!�>�z�<�_�>���=�º>�}�>\Kk>���>�%>�U��`���LR?-�����'�3��䧰�X*B?�zd?�2�>��h�܁�����.�?ny�?�m�?`-v>fth�"+�cm?�<�>h���i
?K:=n��鄈<�c��f���	��C��7��>Q�׽�:�(M��"f��j
?�!?榏�!�̾�׽ �ž5O�<x�?�q?Lj"�H1c��"z���S��g���d���p��!��3��K�|���$p��܊��8:��(��U4?�8�?�U����k�uG(�wҹ>V:�>R՝>!�n>��>���>�<�B�K�!�KXp�@��>��d?���>��9?��2?0�r?2`9?�y�>&��>�nž"G�>SA�=��>��>�4;?�r?��0?ǫ"?�i?p#I>|(�y5־������?p�?��+?=s�>���>�ö��J���5s��׾=3�a�Bg=�3�=��=�n���r���6�=dK>�d?&��l><�i[����>d1?�?X��>�e��}e��OF>�&�>��>=�|>/(�~W�����35�>�}?��X���<x�>$�=���� ���=
b�\�F=&�_J����=;��+>f�>��=óA=m64� o� "�<n�>��?��>nJ�>��{x ����	�=z�X>4S>#>�Gپ�o��=(����g��y>,y�?>��?� i=h��=��=�R��&�����@�����<�?�7#?�KT?��?P�=?4M#?hb>�7��G���]���&����?9\/?���>!��9�農����F��� ?^?�_R��x���-D��̓�[�L�R�Ҽ,�O�O����ֲ�7+�D�=�'�w�z�vU�?\��?D�/>��+�X�����������i?]��>�Ǩ>���>�4��Sa����%A>�m�>ƦR?-\�>x�S?Zp�?~X?Т9>z� ��k��c���F� �\>�K8?��q?�/�?�3g?���>���=\��Hk��꾪,
��b�������>,�1>��~>�?�8�>Ȳ/>���Ͻ�?��_�=¹>ǖ ?՞�>���>
�>dL�N�N?�i?tu��%��9����P�c���m?���?o�?bΟ�#M0����v���<�>�s�?�z�?z�5? ������='/<��پ�澺��>���>4��>��=�?>�aN>	�>�h>J+n��6���/1�x�㼩?�D?v�A>��ӿ1�L�/\H=��ཽ?�=RO���X��3(;�n���u�r<P%�����J���v���to��˶��g��y�޾z���>�F�=�4>�*>���<47�����<9!=������4�=�v>;3�p~>��������L��:~�:����˾��}?+I?Mq+?ΨC?Mz>��>b�1�ֶ�>�	���&?V&U>�?Q�����;�����+�� �ؾ:H׾�d�ᴟ��%>LI��>>33>��=�;�<��=[�s=��=EM���=0�=�s�=c��=,��=��>Yj>�5w?���ǲ��C0Q��P�I�:?�@�>5��=�|ƾ�@?��>>\0�������a��)?���?HS�?��?�ii��f�>��k厽M��=7Ҝ�C)2>���=��2����>��J>@��H������4�?w�@��??㋿�Ͽ!R/>,8>2>��R�JR1��m\��jb�zY�_�!?�;�N+̾�[�>Ky�=�T߾�Sƾ�.=�r6>.fb=�&�&&\��)�=��z�h�;=Y`l=j��>�C>$D�=���z��=V�J=���=�O>�I����4��*���2=3*�=�:b>-�%>��>[�?gX!?�Yo?�k�>a�|��
޾Ju��%�j>��m��ٮ>�!�=ʥ�>��U>�C3? I??�F? ��>�J�<�C�>c��>6hK�,��n�)�m�,�νG}�?�ܜ?���>���<��\����f���P�D?ǴT?�"?&�>�U����/Y&���.�����Hk2�+=�mr�+PU�7���1m���㽱�=�p�>���>��>Ty>�9>��N>��>��> 8�<�q�=�֌�"��<*�� ��=f�����<�wżЍ����&���+����O�;*��;<�]<w��;�z�=���>�P>Fd�>NS�=�⳾�/>r�����L�rC�=VS��v4B�^7d��E~�L/��6��XB>�W>.:���5��7�?�Z>�y?>Fw�?�lu?v� >����Sվ:S��ٴd��UT�Fc�=�	>�<�bD;��`�{�M��zҾ�K�>���>�|>�ļ�j#��%9�K�[�<h��E��>�ʾ�C�矧�����3���[���r�_D^��<?J������=�v�?w�)?��?�~I?�ػ=b����}>�;^��]�>w�Y�V� �dN�=|�?t�@?��'?l!��~7�@L̾0��l�>z@I���O��Õ�a�0�`��Է�[��>������о�&3�e��Z���j�B�^r���>ðO?��?�(b�cX���WO����=��~r?�g?s"�>�I?�:? >���v�����=��n?��?[;�?�
>UX�=mc���>u~?lM�?���?��t?=Y�����>TT��v>�y�����=��d=��4=�l>%?�L?�C?A���U��`��uw�[��;�Q�<�\p>ց>3QK>�u>Y2O=!i�=[W>�*�>��>]�+>H5�>(!�>�g��e	���?31��֗=��%?>PS�=�i(>I��>�H�;�w���������5��p�9mƽ����y1\=;`�>��ֿ�Ny?f;�>>���>�>1���v7��T�&>�P�>i�ǽ�?e�->�q�>���>���>��C>��>q�s=�Ӿ��>���y!�XC��R�МѾ�z>[o���&�	�������I��D���T��j�M.���K=�}��<=�?+���+�k�T�)�W��� �?@�>�5?Ō�l���>��>��>�}��휕��Ӎ� |�l�?��?�;c>��>F�W?"�?��1�3��uZ�(�u�j(A�'e�O�`��፿�����
�S��/�_?�x?3yA?MS�<!:z>N��?��%�Pӏ��)�>�/�#';�@<=e+�>%*���`�u�Ӿ}�þ�7��HF>��o?6%�?rY?5TV��[O�]->��8?�(9?��n?�I.?��4?(���Q#?��;>+/?�D?W6?�e)?�M?/�K>Z�=�f�I�=:������̽EN���;�;���<+��=�<W<ȼ�'K���=�5����{�lL;���� �<��$=�-�=X��=,��>z]F?F�>�Q> >9?H��=6��9駾./?��x=����UǾ�GQ�����4�>���?`Ҳ?�?���>��q��{u��$�>3��>J?_>��5>�ԗ>��V�pLF�@��=B��>@��>T\9���o�&�ľ%*����Ӿa�<��8>T��>�8|>���X�&>���I�t��Tf>hUR�Z���&S�	H��2�[lt�x��>�DL?G�?���=���61����e��c(?��<?#�M?F�?���=��۾D?:�ISJ�{i����>�v�<�'	��Ң�D+��_:��)�rs>+䝾����i4>�U���6&c�W�W�G���ɒ=��Jӗ=*����򆦾�9>�U&>����h6'�(��a{���nL?�(*=����$4n��ٱ��
>�S�>o�>P,<�����vA�������<?��>�y.>����󾊔A��T��r�>?IQ?��b?ï|?���5�j��EH�R���C��"����"?�\�>}?��>�%�=��ɾ�&��g�-@I�
^�>�?^� ��;@������*ܾf2���W>?J�>c�?'�5?�J?�Wt?օ!?���>�x4>uǂ�Ŧv���&?I��?��x=:,˽�Y�F�6���F�(=�>��*?��M��z�>�E?�?��#?��M?��?�?>9��r�:�TҔ>��>�8W������*Y>�K?'?�>�H]?��?ݝ%>�3���w��U��=��>H�1?8$#?��?���>�<�>G���k��=�>�>G|�?���?)��?�b�=��>u�=zs
?��	���t>�q�<��>�:?���?�xn?B!?^U=���4�ս<������<��k�S��#�=Q�<A2=�К;uښ=�l}�i[#�����S�$��&��6����⽇^�>8�s>畾5�1> �ľ-����@>����!������u:�^y�=I��>��?���>�"�G�=�¼>�d�>��((?��?�?i;�b���ھ�K�R��>sB?	��=��l�uk����u���g=H�m?��^?�JW�/��K�b?��]? h�=���þx�b���1�O?.�
?��G���>��~?w�q?A��>$�e� :n�!���Cb���j��ж=Br�>NX�C�d�n?�>]�7?�N�>��b>�%�=�u۾�w��q��`?m�?�?���?z+*>Z�n�F4࿪�������L?Q��>�s���n?��@='�ѾI��p�:�.���>��汾����u�����°��^���.4=���>��q?�nr?��X? ����g�n���q�(zm��m���� ����F����F�8��;�>꾉��ٳ��E�R��?�?N4)���>菉����~�ݾ��j>�K��#|Խx;M=���P-=��F=�Q��.�4�����V?
�>���>��>?M�P�J���9�;�2��[����E>���>+]�>�5�>�˶<���0Խ/<վɮ��DEK�Ђ>��a?aE?�s?%����,�P݃��2'� �1ؚ�X�=>�a>��>kVM����OF!���:���i�s���y���$=��)?y�s>�a�>>��?�?�q��=�Ǿ����;I/��
<�ī>T�q?�k?�z�> u���w�Ը�>��l?���>x�>����Z!�A�{�Ǭʽo%�>��>5��>R�o>�,��"\��j��n����9�.t�=�h?����|�`���>vR?7�:��G<�|�>��v���!�U��6�'���>�|?y��=М;>Fž�$���{��7���$5?\�>?U���>E���!>��,?x�>��?
Q�?����Bｾf�޾9T,?=#A?bX??�>?�?7��>M��=�J��7�r�&>�a>�c>���="��>�蟾������=E=+=�B=�}����)R>V΂��W�=���,>�E�&ZQ�絾�?�P=�\>�6ɑ�V�]��+H��պ������Ą�R��IzT��:N���w��ۈ�-$����?~��?��p��/\�����K&���@����>�z��(+Ѽ�Ԟ�蔖�������ľl?��S�J�S�5o�]kw��(?�O����ȿ�⡿8'�'�?��?R�z?�����"�S<��#>ǃ<��o�WY�@0����ο�٬[?}��>�_�d���<��>���>�R>�gn>�����l��Gkv<#?hQ-?�A�>��{���ȿ��"�<���?��@�fA?)�2���@V=�i�>��	?e�A>#�0����#�����>��?sߊ?w�F=��X�-	��e?��<v!F���һ��=�!�=�U=6?�1�I>#��>���_�>�xOٽ�4>�Z�>�&��f��_�$x�<��\>srؽ�+��2Մ?{\�vf���/��T��6U>��T?+�>�:�=��,?P7H�e}Ͽ��\��*a?�0�?��?1�(?ۿ�ٚ>��ܾz�M?aD6?���>�d&��t�~��=�9�?���5���&V����=6��>�>Ղ,�ϋ���O�;J�����=B�E�ƿ�S �],�:�<��y+r�ud��8��� �*��Z���8f�;�񽍁�=@�=�`O>~m�>�RR>;P>�U?�
k?;	�>�>��9���;
Ծx�o�������V ��w��;졾�r�E�۾؂���n��
Ծ�26���,<�g?�S.��Y�0��$~�E�I��X3?lJq=<�¾��H���(>v}�jԒ�W�=1�K�s���u-�BJt��ҥ?�"5?M?��	�l��]B��=�̐=��s?�m���,����|��<�"��"�:Џ�>��=�^��Ӯ$�OW�dd0?�<!?�f������8Y&>�߽{�/=X�,?�?̀e�ʦ�>\�??������Hb>��@>���>�E�>0v>�����뽚�?��T?�f�6y����>eƾc����=g">z�#����mIK>'�)<�=��+�f�����C�<��Y?EΞ>��)�%_��4���*̼uB�<�O~?�0?��r>kye?��3?�k3=��EKV�E���A��=��Z?��j?Ӥ>�Io��uξb3���5?�`f?R�e>�C��iھ��-���3�?S�j?�?�5�Pk���c��a� �gy(?�v?y�]�$P��d~���M�L'�>�6�>	��>�}4���>�X??�%�S���<���7���?�@��?lգ<|��}<�=�n?>�>;fV�aǾBD������ފ==f�>�7��==u�$�#�QE,�.�:?��?í�>Յz�O�Al�=�^��L�?!�?݈��I�������d�������ؽ�~;�y�=�䅽�̾s���zپ��
�վ�2�\�m>�=@j��<Q�>H���vοT�ֿ�B��4˾��w���?��=�+��m�FvA����R���B�i���*�>���=Ċ�Y�+>���Q��ه��?�z��Xo_>�|��Ql��Ѿ=p<�>�o�>e>�S�����Hj�?$,۾�/ݿ���D�*�> _?�{�?��?�!!?�_¼*Y�����J�]��>?�kp?ќL?9N�=;��U�r�j?�f���S`���4��>E��/U>�'3?aC�>��-�/�|=1>���>m>i%/�ސĿbԶ�Ⱥ�����?��?�g�l��>�~�?�k+?�i��5���T��9�*�ul�n<A?
2>�����!�R.=�Iɒ�K�
?^y0?r{�[/�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?5%�>��?Os�=�c�>c�=�ﰾ��-�b#>��=��>�:�?��M?�M�>e�=E�8�!/��[F�`GR�y#��C�c�>N�a?��L?Kb>v!���$2�?!��pͽU`1��\��S@���,�n�߽�$5>��=>�>��D�5Ӿ��?Sp�!�ؿ�i���o'��54?���>�?���ֳt�w���;_?Gz�>7�,���%���A�T��?�G�?5�?,�׾HQ̼A>��>�I�>V�ԽD�������
�7>�B?���D��Y�o���>���?��@�ծ?di�/	? �)P��`~�ڀ�J�6����=&�7?�)���z>&��>��=�lv�������s���>cB�?�z�?k��>�l?�}o�G�B�V�1=�H�>��k?�q?dHm� �0�B>�? ������OK�� f?3�
@qt@�^?����ӿ�1��Z��k�˾-��=y��=Gqr>������=��=
�X���t�=`|�>�>�D>=B=>x_>��M>����"�ym�������:���.�|�)��y���A!���S�A��䇖�!K�ԨR=�?�����M[���Æ��"����=��V?�R?ro?�H�>��|�A>�. �El =<���ƈ=S��>��1?Q�N?@N*?��=Y��ye��F㤾n����>MK>��>'r�>_�>q\�<H>NF>���>P��=��P=ۋ�;���<Y�K>�~�>��>�a�>E��>�\V=ܗп-g���r���a���ȕ�LM�?����?�3������5�X�_�y>'�'?u�������Pο�3����@?e�����*���\��W>�"?.C?X��=���@��즎����H2��n	>\E������:���J��� ?#�n>��l>"�9���:��,S�6��$�|>��8?����>�BI{���D����5\S>+ܸ>`����������{�"�e���=f:?C�?c�������hu�����R>��S>�L=m�=M9S>�֔�Jv׽Y�M���<��=`n> ?�� >$7�=g��>�����<�i8�>F~J>�.;>'�@?�h&?�x%�����G��[DD���}>���>E�><�>�yC�8E�=p��>1R>��(���� ����0�{�_>�!^�l�_��х�_t=C���~	>Ξ=���7�2���<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?��D>�z�?�w?��>������*�����G����RV=o�$=෎>�N�=�x����'�'�������o��N��u@>��X=���>�J�����#~�=#{+�ż��᩽*��>���>�rl>��>�Q?��>��>*��<�����f��*G���K?���?'���2n��N�<f��=:�^��&?�I4?&l[�w�Ͼ�ը>�\?i?�[?d�>7��I>��@迿7~��թ�<��K>"4�>�H�>�$���FK>��Ծ�4D�Yp�>�ϗ>�����?ھ�,��:N��RB�>�e!?���>�Ү=ޙ ?Ŝ#?�j>b)�>�`E��9����E�7��>��>%I?�~?��?sӹ��Y3�����桿��[�k:N>{�x?�U?�ɕ>L�������hlE��BI�����+��?Gtg?�S��?#2�?�??��A?�(f>��Oؾ𥭽��>��!?t�Q�A�JO&�(��?&O?���>�ᒽֽ�ּ����s����?*\?�B&?N�� a�P�¾�#�<_"�/�T�Ơ�;?D��>]�>Fy��*��=�>麰=�[m��B6��zg<`��=�q�>s	�=�$7�g���*=,?=�G�bۃ��=o�r�xD���>�IL>�����^?&l=��{�����x���U�� �?���?Yk�?��6�h��$=?�?k	?�"�>�J���}޾r��HQw��}x�fw���>���>��l���:���͙���F����ŽY����>>���>� ?#�>���>�K�����.;6&��0t����+��Q�����J��3���슾�����h׾�%T���>����_�?�@?1�>�ސ>��?��P�A�S>'>nL?
��>�� >x d>�=K>���KR?����ݾ'����䱰��3B?`qd?\2�>��h�9���_���~?���?�r�?y;v>�}h�++��n??�>{���p
?a[:=�F��7�<U�����c4��/�9��>�D׽h :��M��mf��j
?f/?�
��H�̾�:׽M�����<=��?Ks$?E�$��V�-�q�10T�_�V�"����a����l(��Yh��7��V�������)�Z�<w�-?|R�?������q���?Pj�S�:��w>Y��>��>΅�>��S>"
��z4��6V��*�|0�����>�Ry?U�>�8?B�%?�l]?�O<?r{�>+)�>Ĺ����>2l�퐃>���>R<D?��?a�M?s2#?�:?���>��$�ݬ���*�4?TT?u?�?\�? P������:�Qm���}�@;b�(e�<K��=���;��ܼ���=	�>jY?�Z��d8����l�>�A?b( ?��>��c�
�U�w�=J�>ל
?�2U>u|�1c�DV����>$[�?��_�=J�3><��=0�޼4����>h!�<f�	>�H=���ӻ���=V�=�f{�6=!y
�L���w��u�>��?���>�A�>T@��� �����k�=:Y>�S>�>dFپ�|��V$����g��dy>�w�?�z�? �f=��=̗�=�|��kV���������R��<��?�I#?�UT?���?'�=?yh#?ĵ>|+�.M���]��?��L�?V�2?
�k>B1J��q/��f{L��x?t!?V���V��x��'D�]֜�
�+=��,��Ѓ������[�d[���� =v��?��?`i<)�*�nž�[���[侠�D?v?a-�>�%�>��l�iG4�� ��
�=�+�>�bT?���>�W?�@Z?-t?)�7>B�۾�׸�5Ϩ�C�#�B��>�3?�dI?���?f �?�K�=����֑Ҿ�������F='�p��븾G!]>${>�u>S�>��{>��=��4�A-�ȵ��a�>�C�����>7��>��>B��>��=�#P?��?�����D������x,�;I��Z�~?Lx�?��>�cF=�j(�W
����m�D>`�?Eũ?h%<?_�l<o'> PS<�G���P��8-�>Ί�>ۊ�>cg}>  >�=\=U�>@pS>}�?�ӿ�<C.�~�Y��K�>=�@?9��<v9Կ%{\���(>�V�N�D=G� � ~�z�>�أ���g�>fR+�m�>F⾺=�=������b�H��[7Ծ�;��O?&�=C'�=�8m=�=���\a��=Ő��Y{t���+=���=��u��̱;n~��𶨽���-0���F���˾͎}?�;I?��+?��C?�y>p=>��3����>���A?�V>'�P�����J�;�������*�ؾ�v׾��c�˟�F>~dI�{�>j73>�B�=�?�<��=�s=�Ǝ=�IQ�=~$�=8P�=sd�=>��=��>0W>�6w?E���𲝿�4Q�7Y罱�:?9�>8{�=b�ƾL@?��>>�2�������b��-?}��?�T�?X�?�si��d�>D���㎽�q�=Ḝ�>2>���=�2����>:�J>���K��i���x4�?��@��??�ዿѢϿH`/>�f6>�>�R��S1��[��a��X���!?`�:�s̾���>aD�=�M߾�Ǿ62=�r6>��`=.�V\����=��z�H:=�\j=�X�>5C>~�=�鯽�:�=�-F=z��=�P>�#Ϻ�{2���/�Nr2=�&�=�cc>A�%>��>��
?�!?�8w?-	�>�;s�6G־�6׾ݾ�>��:��>� z=��>Hg>>O?�.{??PI?��>\�_>���>���>�)�{���/���ľ����؏?�x�?s4c>f;Ł^�oؾC�� ���"?& Y?WI
?zh�>xU����X&�!�.�S���c�2��+='nr��JU����Im�^����=�o�>��>��> Sy>��9>��N>�>�>�F�<Yt�=�}��<`���ⴄ=Թ��!�<�ż�����d'��+������"�;E|�;��]<%��;A#�=���>`$>���>��=������2>|7���M�U�=���oC��	e�K�n}-�(�7�{|A>�Q>o����7��*)?��Z>*2A>���?�Yw?Ф%>�	��<Ͼ�X��=�^���[��&�=��>z�8�޵8���]���K�
о�@�>#��>8�C>�6>�L3�=��	�=���`�X���?M�n�,3��X���d���Ή�q����`�W�@�i?���y��=nB�?��U?��?��;?_2�='/��c=>DB㽁Y�>D�P�
1_�ʽٽ��?6�=?j�=?�t���| �|K̾�#����>�CI���O�Bĕ�)�0��n� ҷ�ۍ�>������оp'3�xe��2���ďB�~_r���>f�O?K�?�5b�TZ��WO�����&���s? �g?�"�>rF?
:?S)���y�x�� ��=u�n?���?�<�?��
>�>$��>�?���?�s�?�_}?�=�2�>/�~:j�>�½{�>Y`:�qjɽ}�U>�P?Xz?0�?e�&���ɾtxƾ�q羂����漡�= M�>�F�>���>��=��ᚽD�%>���>�*�>OhJ>(�j>w��=��ɾL�#��>�e�=2�$>��?ǅ�>�C�i�=Θ;>|=D^ҽ�iz�/���W���������F������M�>]ֿk�?�6�>�P�Gۻ>��7
&�֐�=_]�>p��|(?_~d>, �>�ї>�R�>o;�=1�^>���=�`�	��=�C���93�e�`�����j>R����&�� ����Bу� ���?���Xi�>턿l3?��*ͼw�?߯��r��'� �E�,��>
��>_B;?|�]��GؽB3�=+.�>��o>͌����菿O����?kb�?�Ec>�	�>+�W?��?zl1�b�2��iZ���u�yA�4e��`��ٍ�d���ؖ
������_?��x?�wA?4ߓ<[8z>��?z�%��׏�w�>9./�6$;�J�;=."�>���#�`��ӾY�þ<<��$F>��o?Z(�?�W??V��ģ����=��3?�}B?NEy?��9?�S1?&�u:"?���=f>?��?�0?f%?w�?��b>z�>#z_=���=IW���ě�j���O�e뼋�%��!1=��=��j�S�n=�wS=�hj��8����1�9<1w=��L=Z�=��>�9�>^�\?��>�J#>�!.?Z�;.&�S���g�*?~��</�p��Ym�����Q�=Q�l?�m�?�/l?��>�!Z�]��K�R>3��>�d�>�c>���>0֌� �ƾ��=�R>�ͫ>��<f���¾�. �[:����>j��>N��>��>bb��[�>�⡾�p�5(j>FSM��ﵾ#,R��mE�݁3��o�d�>M)L?��?�׭=��Y)��d�e�}&?o<?нN?�?T،=s?վ�
<�{�L�W@�n��>�=[���ݢ��a���8��I����s>�\��G���:2>���җ�l�+�E�
eԾ��=�q�����E���1������0�1>�S?=
��P�"�1U���V���98?�Q�<����,58�*P�����=6/e>�Ǒ>��0�bk��e>�hé�t
3=�� ?_�3>u��8��^bQ����+�>�.F?��_?[�?~1��e�q���C�����9��g����	?f�>��?M0H>wB�=�ݴ�<B��d�;F���>���>B��c%E�?��'y��$��w�>�?j�>Je?�dP?%~?${`?'�)?v�?v�>����� ��i�(?]r�?��=�|��C�]�à3�2�B�r��>�7?�cG����>;�?�R?�:#?07Q?�?�B#>��辉�,�Ѿ�>�>�X�ш���=>�IO?-+�>7�]?
�?4�%>͠2�S���g��t]�=i�> �9?�@?��?�>�?2���Fƣ=�W?n�?-Y�?	�z?-`���K?e�?(%!?)�޾()�>X�V>X��>�_B?[��?�g�?]{Q?�Cn��$`��'����=�xK=ׯ���=̋�J�2�&�C<�:����=������P�.��$���VWĽ�Ԏ� \�>��s>����0>'�ľ�O��R�@>)���WO��Uފ��|:��޷=���>^�?&��>�^#����=r��>|D�>]���2(?��??�%;t�b���ھQ�K�j�>4B?���=��l�8���[�u�"h=��m?��^?f~W�8��!�b?M�]?�e��=�v�þ!�b���u�O?��
?m�G�e�>��~?A�q?ɹ�>�e��:n����Cb��j�+Ѷ=�q�>zX���d��@�>�7?�M�>@�b>d*�=�u۾Y�w�]r���?h�?��?0��?�)*>��n�4�b޾����K:?ZN�>�쯾�"?��=j����\���d,��_�Zz��!�Ѿ:>e��N���7����q�<c��7�>��?e m?�:?�'W?�q����f��oi�Rv��	�V��� 
�9
�|	A��~*�����6�	�о�ؤ��s�=����"�D�@]�?'(?W�$�>C�>�(��}?���W��3>�J��`�w�w��=�rc=$K��=�Ϝ���S�`���?�p�>�>
E6?�L���@�H/=���3�'���T>{�>7�>���>���/�}c����پГ�����e�>��i?�	D?"[^?�xc��i#�ܬ��(��-�e�ꑀ�,}E>k�=�?�>^w��K&��4��t6��%_����K���z�
�.��SH?Mq�>��>���?Z0?�m߾�� �&B�������8<=NGb>��T?e�
?���>�#�����x��>�m?"�>�>�ƍ��� ��{��ν$��>�4�>|*�>�!r>�d-��\�.!��1����%8��&�=��g?�ă�z�_�Ք�>�P?� 6��@<���>��m�|�!���� t)�Q�	>&g?	��=��=>��ľQ�
u{�⤉��^)?a.?���**�]>~>C0"?TF�>�y�>�x�?�ٛ>'�¾x�a�w�?ل^?�RJ?�A?���>��&=�5���Ƚ�;'��+=��>G[>�'r=���=���0/\�`��0+F=7�=(7м7總�;
<�ΰ�G�L<���<�i3>��ۿ!MK�\i׾�m�g��y�j��P,������;�	��յ��镾��y��X��4:�N%T�j�j�齍��o�5\�?���?Iޖ�p;���Ӛ�2؀�kY��A��>��j���s�֭�O��Y���y�2Ū��� ��
N�Q�g�bSe�G�'?����߽ǿﰡ��:ܾ�  ?�A ?<�y?��6�"��8��� >+?�<T,����뾳�����ο������^??��>�-�����>���>0�X>#Hq>$���螾�2�<��?�-?b��>F�r�%�ɿ\����¤<���?(�@{A?*�(�?��R�V=W��>��	?;�?>�V1�>������]�>?8�?���?IqM=��W���	�zue?C�<��F�Η޻���=Q�=�-=���/�J>uV�>\b��<A���ܽ6�4>���>"�"�W��Rh^����<��]>��ս+ޔ�5Մ?-{\��f���/��T��U>��T?�*�>R:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?$�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�ۅ�=�6�.���{���&V����=X��>c�>Ȃ,������O��I��X��=4k���ƿY%����0��<G*\;%$;����eد� D�s��$p������o==��=��S>���>�8T>��Y>=W?Rfi?��>�|>���A���ξGw.�l���~��c΋�*�����`�꾃��f�����3W�}&ƾw�W��'�<�+=�`���~�2�c釿�-���-?�B�=�
���]��n>ӄ�<sT��P׽�#��v����%�7�y���?&�C?�ۗ�n1n�e�0�~�<��d>��?���&��9k��=>F=�N��+�I&�>�L>8�Ͻ���j�K�&O0?>�?+�������1>HF �A��<+?�?k�<4��>��%?N)'�Z-体vc>]G6>�}�>�5�>�
>���]�ܽ1p?H:T?~��Y<��0P�>�t��~���e=�~>�O3�+F�hw[>���<L��B)�ꡄ�d�<z(W?q��>,�)�`�qb��Q��\==2�x?��?�,�>�zk?��B?���<Oh��+�S���?dw=��W?s)i?�>����|	оe���>�5?��e?��N>mbh���� �.�iU��#?��n?d_?҃��w}�g�����Ln6?��v?�r^�ss�����!�V��=�>\�>���>��9��k�>�>?#��G������bY4�#Þ?��@���?��;<8 ���=�;?h\�>��O��>ƾ�z������c�q=�"�>󌧾lev�����Q,�c�8?͠�?���>������M��=�����? [�?΀�\�
=�g�S�i�����Cؼ`F�=v�#=Um�23¾�qr�ܘ۾�e�������<h�p>S�@��g=d��>�Խ�VпP�Կ�����Ӥ�Sx���B#?j|>��>�Ҡ��Q��z���K�X">�nñ����>�G>QR�񌬾�쁿��G��({;Z�?�è�)
k>u����3��7V����I��v�>Z��>�%�>a߽�'�ξ���?~�߾:ѿx���=y���_?�ԡ?O��?�?��9�:�[�ۖv��	g��2?��p?��]?n
=L�E�)肽%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�W�_?'�a�S�p���-���ƽ�ۡ>��0��e\�@N�� ���Xe�
��Ay����?G^�?c�?۵�� #�Z6%?�>g����8Ǿ=�<���>�(�>�)N>�H_���u>����:��h	>���?�~�?Rj?���������U>�}?�&�>�?���=�B�>�%�=u�~0��[#>@��=�S>�/�?��M?�H�>�4�=H�8�2$/�$UF� KR�L�*�C���>�a?}�L?$\b>� ��22��!��Aͽ�f1����c@��1,��R߽�05>�=>>��D���Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>A�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�	?\�?P���_~�m��+7�|��=��7?�/�4�z>x��>^�=hnv������s�޸�>!A�?�x�?��>�l?�o�7�B���1=qO�>��k?]w?)�n�e��B>_�?W��8����L�?f?��
@�t@��^?�좿��Ͽ� ���w{�-���Bn�=y�<� >�N���鼐`��	!��Q#r=Mq>J��>���=[m0>h� >qF>�X�=���s��Ȋ�y6���?��*�ѝ�x&��ئ)�$O;�?��.���K�_�=>lh�����������`����=aWV?�P?S�n?��?<y�N(>����G4=���e�=^Մ>5?ML?8�*?�	u=! ��h6b�����(���(���ؽ>Z>8Q�>�Y�>�>���;��L>&$>/�>�X>��%=����H=u6_>E�>߯�>�2�>�'_>�#>y�ĿԵ������	����<�i�?�_����g�����������"��@���5? �>sn��|���x���@?�윾�-��5��u9>��1?�N*?oU>~ƾ�����|=�A�Vc�4�R>��4�yf���#���C=�Y�>��>�[T>�X��P�Q�W�\:׾'�>6�X? ��q���ڍ��Z8�����,�>�>+ߺ�����3������3�_���=aJ?�:?}���)�پ������ƾ�W9>�V�>�|ɽ���<��>�5;�J��/Ⱦh�<�;�k�>�U?�,>�ގ=���>�V����O�(s�>(aB>`-,>�@?�!%?������ɍ���-���v>�W�>��>>�=J��t�=?b�>�a>��;׃�j��9�?��@W>��|��f_��\u�Ty=Ǘ��v�=�ۓ=} ���<�s&=�~?���'䈿��e���lD?Q+?Y �=�F<��"�E ���H��G�?r�@m�?��	��V�?�?�@�?��I��=}�>׫>�ξ�L��?��Ž5Ǣ�ʔ	�,)#�jS�?��?��/�Zʋ�<l��6>�^%?��ӾOh�>yx��Z�������u�e�#=P��>�8H?�V����O�i>��v
?�?�^�੤���ȿ5|v����>W�?���?g�m��A���@����>;��?�gY?loi>�g۾<`Z����>ѻ@?�R?
�>�9�z�'���?�޶?֯�?h��>���?R��?�c��}R�����L���2n�xIP�ɱ�>�\>�'V>8<��� Q��"k�Eь��F+��S���7>�=-�>��='����ܽ�9��$=��?�R=[�>>zJ�>4h=Ut\>d\�>��>?��>ky;�m�m�����|�A�K?uƏ?-��AIm���<3�=0Ad���?��3?7�
���ξ1�>{p]?3�?��Z?J�>r��E���Wq���ڳ��ʉ<�F>L��>pp�>����I�I>�gӾl�@�`�>���>�"v�-�־%�������D�>�`!?��>~v�=�� ?+�#?�j>�#�>�aE�9���E�ͯ�>R��>|J?\�~?l�?Zҹ��W3�����桿1�[��1N>��x?-U?�ȕ>����F���;<E�<I�����?�tg?DO�0?&0�?Չ??צA?	+f>��ؾ/���o�>r�!?�����A��L&���>�?�s?��>�r����ֽ�Oؼn��������?n\?�E&?'����`��þ�O�<��0�M�X��a <|%H��>
>�$��̍�=�->yʯ=�l�A�5�o�v<bt�=?D�>��=g�7�����-=,?��G��ۃ�c�=��r�6xD���>�JL>)��k�^?�l=���{�����x��6	U��?��?Hk�?h��"�h��$=?�?C	?"�>�J�� ~޾0�ྲPw�~x��w���>���>͚l���K���֙���F����Ž��Q��*�>��>O��>��>vRT>T��>'x����� ��Q���~Q�=���R��!�U��{y�� �TӠ�m[Ͼ,���	<Q>� =G��>��D?��>��A>��>e��=��>�=->m�T>s��>g/�>�e�>��=����KR?�����'�b�辔���U3B?�qd?'1�>�i�*������p�?���?Ns�?U=v>h��,+�tn?|>�>>��>q
?iS:=m0��@�<V��f���2����̪�>ND׽� :��M��nf�kj
?�/?
����̾o;׽� ־cb6���?�`%?f&�#\�gj|���Z��X��=���vd��o;�K	"���U�c���>�s�����,���G���2?��?9x�"��q3����w�$/�a�>�+�>�J�>���>`�7>us���8��%N������^�(�>5g?T7�>gh@?!.?�p^?#e?�x�>�H>pn��� ?�f�����>��>�<?�)?��??H�?�9?<)y>�ɽ���޾�]?��?qR?{��>§	?�Y�24�߸f�"q�<�%���R=ج>"�L��w<�>�s�>�W?5��-�8�����Uk>&�7?���>���>A��C,����<p�>�
?DF�>  �}r��b��V�>)��?����u=o�)>���=�����"ԺcX�=v��� �=�,���x;���<��=���=��s�A�|�q��:�_�;��< u�>6�?���>�C�>�@��.� �b��f�=�Y>=S>|>�Eپ�}���$��u�g��]y>�w�?�z�?ѻf=��=��=}���U�����G������<�?>J#?)XT?_��?{�=?_j#?е>+�jM���^�������?	�"?�F�>-��� �n���'M����>c6?\���V��yk��^���[d�0?>)!�[燿Jd��{�S���Cz�۟���!�?�'�?^�w=�N��������xξ&�2?�?BR�>e$?48���f�qa/��!>�
?�a?�[�>�]?��n?t -?�xf>�$� ��������=��>��/?��:?Zߊ?�Tz?>��>7O½��v��þ�1ݾ][׼3�@��~��&��>_��>��h>�4�>��r>��P>G̖��g,=�(��E0>0�<> ��>㧘>)9�>�� ?1�˻��M?��>K>���>�����{2��t)��I�?Zm�?��?�P=2��$-��xվ�w�>�x�?��?zi2?9��	m�=U�8�B�˾}����(�>_��>#�>�6�=<=���=;�>eP�>��:��7�+�����	?�D?^I��ӿaw������$�bH�;���iɈ�]A�,ﹾ��n�en��*�`=iJJ���=�{¾��Y���	��c�����?M�a�77�=�^�=9ȻB�D�i��[d=��0�&_(> x0��>"bm�&�����!��=���c�E�`Z�=6�˾G�}?_8I?ْ+?��C?7�y>�G>ȏ3�4��>�����??�V>R�P���-�;�9�������ؾ�w׾��c��ϟ�a?>YI��>�M3>[�=�D�<�!�=�_s=7��=��T��=A3�=k�=�l�=���=��>S>s6w?���u����5Q�/b罼�:?�8�>p��=�ƾ�@?M�>>#2��	���b��,?9��?PT�?W�?1xi��d�>_��r⎽�r�=z���;2>f��=f�2����>��J>i��K���}���4�?Q�@Ŝ??�ዿ��Ͽa/>�p>>�.>��\���9��Z����j��u>�w�.?qY;�~�޾��p>8�=����$Ӿb=�Aa>��=�&��Ma����= *���"=�JB=���>V�U>��=���I�=%��<n�=z8>�R5������Մ���<#�=�}B>� >��?�?�?%?�w?��>�-{�sEӾG������>N�<}��>���=W)�>���>�+g?F6?�[?7%?�,�>	�>�=�>U~��:w���6�5*l�=P�=U�?赛?�·>3�G�I��c�`m�v����?!�#?��?�? ��rT࿧^'��y-�Ӝ�}3<IxL=��o�rY�e�q��q��c��=*%�>���>F�>W�u>�p:>��M>���>��>6��<�ψ=���P<mO�����=`¹����<�Ƽ"�;�ΰ�6C�QG��p�;4�:	��;��=<���=���>�7>��>T��=;���C/>����8�L����=KB��~*B��1d��I~�&/��d6�ޭB>�0X>�����3����?��Y>E?>��?[Gu?� >U'�y�վ�N��e�`ZS��Ƹ=��>+�<��o;��O`��M�QvҾ_��>�+�>�:�>�{4>N�&�M�@�44�<\Uɾ��7�<a�>XE��p�_�v��4Sl�&�������,�c���.�2J.?����m�=πv?r�S?5�?.?V!=���F>پ���c}>T �`�7�@��$�?H:4?[C
?|�����'�-����72�>3�N��M��Q��s+5���[�>l���Q�>ݸ��̩�
Y4���}�����&�9�ܗ�9o�>v�=?<��?C���憿�[�B�	�ӽ\#?b�x?�ʻ>��?���>��A����Ū
>3e?�n�?^�?Y�=τ�(�%�r��>c��>-��?�Η?+;�?�v�ӣ�>�x�<��>�na�<0<;�U�	L
>?p�=:?���>��>勽K'���m۾�ƍ��T.>�_�=�-m>��|>��>.�h<7�I+>��>�%�>o�>h[�=sZ�>��>����(�X��>���=�PQ>�qC?���>K?�=��̽���=@��������!
�����<��=틺��Md=���O�>�ѿ����?�Hh>�w��s�>[���Լ��=��x>����a�>Y<�=w��>톆>�ţ>�=-D>��v>�FӾS~>����d!�L,C��R�H�Ѿ |z>M���o&�֠�do��CI�cm��Ih�tj�t.��u<=���<�F�?մ��8�k���)�u�����?�[�>$6?�،������>$��>�ȍ>2M������Ǎ��c���?G��?�;c>��>G�W?�?ڒ1�23�vZ�(�u�h(A�+e�S�`��፿�����
�v��.�_?�x?2yA?TS�<-:z>Q��?��%�`ӏ��)�>�/�$';�.@<=�+�>*��1�`���Ӿ��þ�7��HF>��o?:%�?uY?=TV��j�|'>�|:?K�1?}�t?\�1?��:?��C�$?�2>��?��?H5?M�.?�/?��2>�i�=9��ɣ)=DՑ�����kн�Ƚ���H2=B�=�:9��;i�=�e�<���|�%;/n��~(�<z>=���=%��=��>��\?�(�>���>[�8?�<��a8�}⬾��/?�1"=/�y�bt�����������>��j?�&�?&2Z?�Ef>sX@��;C�y�>���>��">�|Y>?�>���D5J�
R�=r�>#�>s��=`eH��wz�3]	������0�<�$>���>A|>���b�'>�}���$z���d>��Q��ͺ�C�S��G���1�y�v�xX�>6�K?u�?}��=�]�3"���Bf��-)?�_<?sOM?��?2�=a�۾��9��J�)R���>	4�<������8&��q�:�oX�:�s>
(��n㠾��a>����޾&[n��I��D�AfP=�W�.X=o�`�վ���C��=�9
>����e%!����a����J?"�h=�ڤ��=U�R��1�>�Q�>g®>��<�Kv�`@��h���Z�=-��>Z�:>�������^(G�{,�(?�>e�F?�5Y?�!�?���$ ]���\������&��+����E?���>��?�I3>/�=h賾�9	�[\�_�m�n� ?���>ĵ!���
���ھܒ$�������>U��>���>�>1?�6?&��>�N?H�7?���>�؟>������	���1?��?WΚ�-+�=�ݰ��<X�=�1���'?a[E?���	?EN,?�?�?��=?t��>�[	>K�ľ�Dj�ݪ�>��>Grl�_�����>8�"?�)?��?V*�?z4�+M�@��<+簽��#���j=}�+?��$?>c&?��?��>�����=$��>�c?�0�?P�o?w��=��?=2>���>���=ᜟ>p��>G?;XO?��s?��J?[��>��<�4��V4���?s���O��Â;��H<��y=����9t��P����<)+�;�f���C�����1�D����_��;�1�>�{s>�����a0>�ž�$���%@>0)��u��4
��b�:�=��>��?�Օ>4�#����=�`�>t��>ܩ�G�(?E}?�/?e;��b��۾�KM�}6�>!A?T�=km�Vc���u��c=��m?��^?�tU��j���b?4�]?�h�&=��þ
�b�݉�&�O?6�
?��G���>��~?��q?���>��e�9n�����Cb��j��Ͷ=Hr�>�W�U�d��?�>/�7?N�>�b>i"�=u۾��w��q���?�?��?9��?�**>\�n��3�%d
��s��a&W?�̫>A(ξB^ ?�A �����$��'������0��HȾ�r���_���yw�9J��q�&���= �>1lU?2�]?�m?�$���f��f�;爿�:o�~�$��^��Z�j�7�� 0��Yg���
81�1�&�/Q&>�%~�L�@�Xٴ?h�$?�P3�ʙ�>����뾋�̾0@A>~���M�R=��sE=�N=�;n�[�.�gP��� ?G��>V\�>m�>?��\���<��2���7�R����'>���>�	�>N*�>;N.;8:,��潓����f}��L˽Z�q>4`c?G>G?n�s?y��7(��x��4��驘��N��j>i0>F�>B*p�j!9�;_(���>�]ks��	�7����z�=�1?��>m6�> e�?.;�>�p�����~W|��p6�꜅<��>��j?��>n��>�ꈽ4g$�K�>�e?i��>�d�=�}��w�Ѿ6��%��=N�2?�4�@c?.M?��#�IF��/�������7�?�@�ަ�?~�4�UvM��>�?��c<�:�>�p7>�����-���=՗�<��?3У�t�Y>ZǙ��������S��u)?�h?s�����)��ǀ>�?�~�>VϨ>A��?�]�>c����}b<�b?Ǐ\?|8I?�:@?47�>��=5"���Ͻ�Z#��0=(w�>�	]>�{t=`>�=9����[��,�nN8=���=�b��$d����<}ͼ�N<���<��2>&mۿ�BK�o�پ2�E�K?
��爾�����c��ò��a��;��nXx�ۍ� '��V��7c�(���n�l����?�=�?���D0�����(���������>~�q�(����{��{)�����u���`d!���O��&i�h�e���'?ٺ��~�ǿ����W4ܾ�( ?O> ?��y?>�'�"�C�8��� >���<��ő��@�ο����Z�^?���>�����\�>��>O�X>�q>~���󞾇ړ<��?�{-?Q��>Y�r���ɿ������<���?��@x}A?��(���쾘V= ��>1�	?��?>�C1�{C�����4W�>|<�?��?܎M=��W���	��~e?��<��F�ny޻Y$�=�:�=m3=G��-�J>LO�>y��NA��6ܽ�4>xօ>�#"����,^���<��]>7�ս#+���̈́?,]��d���+��O�Y�>�V?	 �>�N�=bA.?��G�)	ο�[U��fe?N��?K%�?]�&?��� �>#�ܾ��O?'�4?���>�^'�I&r��-�='���%?�h�龙kU���=���>�>�D(��RR�Uv����=M��ƿ�$�$}��`=8�ݺ��[�~���~�T��#���fo����`�h=���=��Q>�k�>�$W>Z4Z>�fW?J�k?@N�>�>�5����ξcv��G��o��襋�������R��߾e�	���������ɾz=���=�7R������� �;�b��F���.?Yx$>�ʾP�M���,<5pʾi���oW�������8̾��1��n�`ɟ?��A?�����V�X��\�������W?�M����a⬾)��=#���S=o�>�q�=	�⾥3�K{S�>4-?�0?Y��H�����d>�_��+(<�yH?��#?胜�Ĳ>� X?s��<b���{O>2�9>z%�>Y�>5>�������XX?�f8?!6������azo>t�ھB�x��R=XW�=�.����<�L>"�<�P��q�:�C���2:?W?��>0�3�q'���k�Ӛ���$>=oڈ?z� ?��l><ki?0d?��=�U���8E����N�=�K?�M_?�
�=濢�!]ӾF���i�>?C3_?܀0>icm�;�Ⱦ�D5�<���?FVx?F�?�鼻�j�%����~��F?��v?s^�xs�����N�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?r�;<��S��=�;?l\�>��O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������"��=Gٕ��Z�?W�?	����hg<i��,l��n���p�<�Ϋ=��JK"�'��y�7���ƾ\�
����Y׿����>*Z@qU轌+�>�C8�<6� TϿ`���\о�Uq�<�?X�>:�ȽH���
�j�\Ou�ܱG��H�����E<b>5�{�T"(��PV�i�����.�">C�>ǴT��Y�>�����.���g����� �.>X�?�R?��n<g>о���?��+���׿؉����Ҏ?z�?m�u?��	?�H^>���X��T��V�?r�{?>h�?Bk��F�����=$�j?�_��vU`���4�uHE��U>�"3?�B�>S�-�Q�|=�>���>g>�#/�x�Ŀ�ٶ�?���Y��?��?�o���>q��?us+?�i�8���[����*���+��<A?�2>���H�!�B0=�VҒ���
?V~0?{�d.�O_j?E5���q��s=	��:�>�b�>�YT;+���_�0��>�O��ٛ���3���?j�?� �?A
�=�1�#��>5�>�����3d�=��:>���>���>�7�+�^>���D�N�,,K<���?]��?H�>!��X������>Ǭ�?�\�>��?Z��=�-?���=������d�Q�Q>m!>)�ɽb?�D?�C�>��<iip�d2�[F���S����>�b�>��^?�E?H�>�$�Ҵ;س.��^����*�y�E�����6�G(���%w>6&=>D
>�Xݽ\���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�	?�'��E���P~�8��"7���=��7?�E���z>I��>Qת=hv�����`�s��˶>gH�?�t�?��>��l?h�o�� C�6�1=<,�>�k?�?t�j�J��5�B>Ʒ?\��x���"I��f?^�
@�o@��^?n⢿�^��$�~�K�>��7�)�>w�=hFb>����i=��%=8p���A�=% >��T>�	(>�>͙_>=^n>���<ө~�I���/��v
����7��F�.����a۾цC���_� 5?��Q�8h���CW�@z��\���B��3��mN���=H�U?R?|p?� ?$#x��}>����J_=R�#���=�)�>�g2?&�L?w�*?��=������d�{]���@������>�\I>`��>	G�>N!�>^B�8�I>9?>�m�>x� >>'=��׺�=��N>�H�>2��>�d�>��;>�Z>
���D2���qh��Lv�b˽���?Z\����J�R"��;,�������Q�=�N.?��>J���6п׭�JH?���I��y�+�ͪ>��0?Y"W?a�>�"��}mT�Y>�Y�0�j�6�>�P ��5l��n)�݁Q>�C?� >E�_>��=�p�Q�	�1��yH����>�8?S������_�#C��FоA�>r'�>T��M�C��{��#jG���[�sȽ��O?���>���f��$B����'�=N�=>-�f=�Z>"G�=o���
�g�AQ�\��:
��=;w�=zX?DI,>Rj�=�ã>W$��XuP��l�>9UC>��,>1�??�%?���Q����ƪ-�vw>[*�>�׀>3�>�zJ��n�=Rb�>,�a>���6��C��
@��5W>���_��u��z=� ��K��=���=uQ �-=��0&=hg�?�𦿶�n���G����SB8?ض;?���A/���"a�����׾�{�?#@���?&G����C�{��> ��?-੽<ȑ>;�?���>ɐ!���;�?�-r�mk�0�;�)��;��?�d�?�y���tM�-�7�H��ր�>� |�Oh�>{x��Z�������u���#=R��>�8H?�V����O�g>��v
?�?�^�ߩ����ȿ5|v����>W�?���?h�m��A���@����>;��?�gY?roi>�g۾<`Z����>ѻ@?�R?�>�9�~�'���?�޶?֯�?+�H>p�?es?��>�=r��|.��'�������=X��:J��>Y�>a����E������n���dj����Ee>�%=��>+|�?���6�=$�������^��
�>³r>#N>���>�� ?7%�>���>k	=�Q��$��������K?س�?~��
1n��~�<���=I�^�X)?�K4?�[���Ͼߨ>��\?���?V[?�c�>f���=��9濿:�����<��K>�0�>�G�>� ��ZCK>��ԾE5D��o�>�͗>���h<ھ�+���1��?�>�d!?���>�̮=�� ?��#?s�j>��>/OE�k.��-�E�Υ�>&��>�3?��~?�	?۹��Q3�Y��6桿��[��fN>�y?nL?��>�����u���bG�.�I�G"��ך�?�qg?0彦?�2�??�??�A?{�e>���5ؾr����>V�?�ʽ�T��9�`�����?�f??��>)�������u���'��u�
�?��]?��?�G��e�閖�#��eč�9���=P;6�<6"%>֤>�GV�=ֽ >���=��x�T�O��vz�٬�<k�g>gx&=�[a����0=,?��G�}ۃ���=��r�>xD���>�IL>����^?ll=��{�����x��	U� �? ��?Zk�?a��@�h��$=?�?R	?m"�>�J���}޾6�ྼPw�~x��w�\�>���>$�l���K���ڙ���F��]�Žx����>4F�>z�	?��>%�P>���>`����%�����7��'^�����7�G-�f��|�{)*��/��ݛ��l�~�\f�>�[��#��>2�
?�f>�|>y��>0�/�0&�>h�T>�5z>&��>��R>^4>H��=
�2<�l׽;�S?��ʾXh��dϾ� ̾J=?/Rn?�o�>�Y����w�����?��?Ң?�H�>� V�fB(��,�>�?9e��V�?� �<:/���U���㰾τ"��5�-߼4>c��6=5��XU���z�J?�?����Ѿ���Š��~n=O�?��(?��)�b�Q���o���W�-S�����wh��b���$��p��j_�����&�(��~*=�}*?��?l�җ�J���&k��?�#)f>���>��>�Ӿ>LPI>��	�-�1��]�+H'������W�>vZ{?҇�>�I?[<?�wP?hkL?m��>�a�>M/��@o�>�w�;{�>��>%�9?��-?�60?�y?�s+?i0c>�z������ؾ�
?�?�J?�?O�?�����xý)b��Qg��y�,{����=�<�<O�׽�Bu�/�T=�T>k?����1;��� ��3m>��6?��>�>4����|��`�<���>(�?��>����[6r�l�O��>�9�?����4="h(>���=��c�>��:�4�=�'��D��=�9i���-��^�;롴=��=��8���v�%���z�h��Xl<�=�>�)?�L�>9�=��,�T����-�k+=#W�>nM=0~�=3����(��JP���lq��1K>�G�?�Ǽ?ig>��=r�X=�~�g0þ�������&���Q�>�*?*/Y?W�?�P?�(?�?�=�r3��L���������&?,?��>&��!�ʾ�𨿎�3��?^]?�9a�L���:)�'�¾I	ս��>'X/��-~�����D��������u�����?x��?�YA�c�6��}�W���a���C?$�>�Q�>��>��)�n�g�l#�?D;>Ð�>R?�"�>��O?><{?`�[?�eT>a�8�V1���ҙ�`3�"�!>F@?��?��?�y?�r�>��>�)�O�UV��~����;ႾPW=�Z>���>�'�>��>\��=�ǽO��(�>�b�=��b>��>���>��>J�w>��<u�G?���>�Y��N���������N�H�g�t?�J�?�*?�	=@a���E�l���؛�>�|�?Ы?_�*?�R�-0�=_�̼���l�t��׸>��>���>N
�= �\=�>��>��>�r�����8�j�U�3�?;F?�=�п��E�_#+>}-��|WK>k-�	�ɽ�dz��C߾DG�<J���1��*���Ⱦ��߾�ؾK��t� �)B�&��>���@�>�K��Ot<�<$�𽼼�<��|W�=�����������\�=�?�=�>]�r>9~>:��"���,�|?p�H?��>?S�-?@��>>�����=���>�`8�y�?H�J>�*�=�ɾ	Hg��%ʾ������ƾ
�ھ
�;��ւ�WZ>g&�@>�i�=&������y�=��>Ԇ<t�=�&5=$�c>>�N>�\�=�!>��H>�[ �Ps?��Σ�*�������C?�B�>�"��~(��v]?0�|>��c�k���r>�A}?۶@c��?�v�>�Ԥ���>{����X��o�=�x�>�su>b#��u��z�>d�>%�[��z���p(�l��?��?sw�>���87���y�vX0>u�>V�R�~n4��V�ssV�\eN���!?�~7�r^ƾ�}�>��=G߾�þ�>G=}L)>��=�(��X�ڥ�=ȅ�#`=�a=��>,M>��=�9��A��=��Y=;��=�5O>��G�\�<�l�F���-=0�=�b>�b>:��>Z?�A0?�>d?̌�>j?n��sϾ_���|I�>��=�z�>~T�=HB>l�>��7?��D?��K?f��>�?�=O
�>B�>V�,���m�����ɧ��<���?��?�q�>�DF<�@�k���P>�IuŽub?mS1?�?๞>�U����9Y&���.�#����}4��+=�mr��QU�K���Hm�2�㽰�=�p�>���>��>8Ty>�9>��N>��>��>�6�<yp�=ጻ���<� �����=&�����<�vż�����u&�9�+�0�����;t��;I�]<R��;���=���>2>��>5��=����E/>����G�L����=�H���,B�|3d��G~��/��Y6��B>�4X>�p���3���?:�Y>Fh?>E��?C@u?/�>����վ|P���?e�YS�Ƚ�=w�>0=�7{;��Z`��M��|Ҿ|��>*�>��>��l>�,�I!?���w=��_5�a�>w��|���#��9q��?������Bi��պ�D?F��d��=�!~?�I?�?ю�>��M�ؾp,0>^F��
�=���(q�Hg����?_'?���>���D����T�����>�S*��=�D�����%�kNʽϸܾV�>��žC���1����Q݊��2�[2��3��>, *?���?D���f���;`7��!�& �=�?�S?_��>��? �>�.y���ľ_9c�#*�=�Ny?O��?�A�?�]�=`��=����9�>�)	?�?���?`�s?�y?�z�>h��;p� >���E�=!�>���=('�==r?��
?/�
?�h��c�	������=^�8��<{ʡ=���>�l�>I�r>*��=C�g=�u�=�-\>u؞>��>x�d>R�>�O�>W���&=	��p?I=���>_�4?�H�>N��=� ����4=����1��`A������RʽKc6h��dYJ� O��&�>r:��9��?�P>�S�?gT����-��d/>kK>s�ӽ���>��*>��>�?�>ڻ�>�%>鱛>��>CӾox>����k!��&C��tR���Ѿb�z>U����%�������pJI��f��:^�j�"0���?=���<0C�?ݴ����k�{�)�������?@F�>6?�،�l
��@�>_��>ն�>=G��l���oč��_�w�?���?��d>D7�>;�C?��	?�ᮾ�	��i�[�P�jY>�5Jv��B�XH����{�y�Ѿ>����c?��`?�zN?��>�@Q>�+�?���2��}}�>��(�z�,�k7��`�>޾�A��
U����,��,�=�*�?���?]�-?�I��m��u'>r�:?ۛ1? At?8�1?�c;?`��$?�3>�F?Rl?GK5?��.?��
?��1>Pq�=Z[��� '=�����銾SMѽƵʽ�=򼦦2=s�y=�P���;<D�=��<�I�pؼ��0;!����ǫ<��:=�֢=hu�=�`�>ۍc?�/�>�p�=&?�m��?�1����&?p}�t۬��獾�����Kپq�=wr?b֦?�9y?\�\>a�)��(��2>���=�ua>�o> �>�3����<��=	��=$��>}c�=�R�2�;eP'�C䎾*��=��>��>�Q>)��Zg��	߾E�%��̺>�qW�=���2S9��M�23������?��j?��? ?��t	����=:�f��W?�ν>9X�>��?��t=�N����O&�"�_��B�>㐯�< @�Ͷ���k����N�;r˽Y�2><̓�ϴ��5�b>ʳ�a޾ �n�0�I���羠�N=�a�T�T=��_�վ� ��V�=q�	>L����� �������J?��k=�7��g�U�0~����>���>��>�,9���w��v@�n����q�=R��>��:>I��%���vG�:L��7�>^�5?�[?h�?U{��e�f�W�6�������]�=�)7?�O�>Z�!?�=	�0��h׾�����_��a�E4 ?[��>2@'�r�(��QϾ]��LW%��P�>���>W�>�c?78>?�U?tD?^�?��?a�t>_�A=pc��C"?O�}?&��<B��������W>�C1;��A?�s+?G���?�<#?V?�y?�~.?)�?��=�žy@��>(J�>��b��ি�7I>g�L?�̱>�xy?�S�?���A�z$��J1����=;�>�~&?�1)?A.?y�?�h�>J��A�=�H�>�3c?�B�?�jo?�O�=�?��1>��>�Z�=營>�7�>�?�N?�s?|J?�&�>�T�<c����H��~�u�P	e�38A;�?<4�x=!����w�������<�(�;�۳��@��h���<D��4���j�;�R�>$�x>j����>�Ⱦ{����7>� L�ؘ�a,��^�>���=-��>�G?�ݖ>G�'�m؈=�!�>�^�>�2�f)?�?�?�ܢ���_��ؾ�8>�Fӱ>p�>?{�=+m��{����t�Y�4=l^k?ϙ[?/�T�������b?Q�]?/i�=�/�þ*�b��龷�O?/�
?R�G��ҳ>��~?�q?^��>f��5n�.���Gb�q�j����=�q�>�N���d�VE�>ϝ7?k�>��b>0I�=ׂ۾B�w��k��W?6�?��?1�?�B*>��n�`5��� �r��.e?P��>M�"�P��>�� ��c��]��>�!ǾL���I���J�Ǿq#оog�X��$d�=-F?��P?}1}?@mq?O������ʉ�����`���T��P%�wEg�~�0�ު,��慿Vd�3��{<��9>Ty��)�zֲ?.�&?W�����>!����U쾁\��t:
>H����9�����=+��]�ȼ�\�����``��ʾ��?�,�>�ǹ>��>?��U�RmK�8@1���D����x�>
h�>�>,�?���>�5�c�q���ƾ��5������y>f�[?2&@?g<s?���-�����
�
�T��bfȾ)>�k�=0l> ��f�X�j�#� �F�&{����E��H0�3l�=�z?J��>��>�|�?#��>�	�����ǃ��0��	ϼ>A�>Z�R?P�>;��>�7a�98?�؅�>?V?���>��>����������u-�=��>�����>7�}>Ȉ��ؓ��`�z�,���:�h�m�3>��w?�
n�Qw��4`�>fCY?���">O~�>�烽����)����<Ǒ+?7
>A}=�h��&�A�����¾�?� ?jC�&�9��E.���>��>�a?��?��>߇g��.�>��>w�F?B�M?܆?��
?����掾����r2/�*D�=b��>�Y�>ܠ�=�܁>�������P��=y>�j<�y½p��>B��!;5��=��r�
kۿ�?K���پ�	���';
�+ꈾ�����[��z��$^��/�� Sx�E����&��V��+c�楌���l�M��?�;�?�y���1��H���ޕ������ﴽ>_�q�q��!�h��*�����:���`a!���O��!i�νe�<�'?+����ǿ|���[=ܾ*" ?@@ ?%�y?��՜"���8��� >Ug�<������������ο������^?���>��*��> �>P��>��X>�Bq>�
���㞾V�<��?p�-?���>W�r�i�ɿ	������<(��?}�@�HA?Ä(���nT=-�>�	?Ƨ>>h1����尾)��>�F�?�݊?�M=wcW���6�e?��;��F���ͻ���=z��=%=�a��H>�ϒ>+X��\@�]ݽc�3>%Y�>�."�����}^��O�<"\]>��ս���[�?�9]�Zeg�k'0���~��A>�T?��>`m�=�B-?p-G�s�Ͽ�!\�c?���?�`�?r)?a��f�>t۾�-M?��5?9C�>�%��Ot��&�="�����x�ྦྷ:V�Z�=B��>��#>2�-����LR� 䍼���=���ȿ3�'��I����<B��;�.���x.�G�ս0=����Z^�5����&S=���=��a>Ѻt>yrd>��Z>�]L? Ik?���>}/=����C�nʾ��=�A:�	~�_�]����ľP־�~�������Y�������<��u�=jR�����*� �b�g�F���.?�&>~ʾk0M��BM<^ʾ�����x��{��r�ʾ��1�=�m�X��?)�A?l�����V���\���2��y�W?��r/�-I���2�=؅��؃=pҜ>��=9��2��TS���?_�7?!ߕ�m�����˽��ɼ{��?PP?j�E?�gg=�?��Q?�b�����J�t>ovj���?G��>�������}�# ?�?K�A�~�6��(><����T꽊<1>�����R;���Q=b�
=
����r=��M�B�d�T?赘>�*����(ږ�w�$�z�=#�{?�O	?+�>v�m?ݠC?!/<��gvP�]����=�4X??+e?f��= (<��$;Un��?�7?>g?&J>�-c���ݾ;=-�4F�$?L�f?�n?�)ü�~��!���s��S:?��v?s^�xs�����L�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?e�;<��T��=�;?l\�>��O��>ƾ�z������+�q=�"�>���~ev����R,�f�8?ݠ�?���>������+��=�ӕ�FZ�?��?�����fg<R���l�Wg���u�<lӫ=���P%"����"�7���ƾv�
����*���>�W@VZ轏-�>�N8�6�SϿ����cоh q���?�>�\Ƚꛣ���j��Iu�ڱG���H�������>��<(���ž�l�D|�ƙ>�>Ʊ��sQ�>V�~�)�<'��rp���x>^]E?9��>���=I���6v�?J���u�f���9�U*�?��?�҆?�u?ʊ8>\j���ܾ�B���pP?>�?؆�?��R=OB�T>����j?�^���U`�8�4��HE��U>�"3?OC�>N�-���|=%>���>�g>t#/�<�Ŀuٶ�������?��?�o���><��?�s+?�i��7��[��2�*��0*�W<A?i2>����5�!�e0=��Ғ���
?~0?�{��.�k�?{��P���FU�d�>��o>���<������ž�3�=d�0����"R��F��?Ta�?O��?���=Z�Ǿ�7?���>[p�:־�6>k�>�3�>���>ad���>Y����z	�ƔR>��?���?�)�>R����m���B>�o�?���>T�?���=���>�_�=�=�����h�>>G�)>��-�1�?�P?4z�>B��=K�3�S�3��:���P��4��Y?�h�r>gD`?��G?9s>f���ug�Fe$�IK��� ���ɼ�p3��Uu��� ��P<>h8>~d>��U��,ھ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�K�?�������i1{�ץ�ʿl��)>22?T�����o>��>1s=�-t���QJt���>��?;��?	��>�r?(�m�}JL�X�;�Ϗ>aai?��	?"3=;���DM>v?��C���_���q?�*@P�@+eW?z���ο-ٝ�r���&��l�=X��=s��>f�\��U��(��>�vK=�o��n�>2�>�n>�M#>	�==5�=c�C=v����H$����V���'�x\�v����pH�*�4�myĽ��)���������X��\ 1��ð<�K�y�����T�=��M?{O?��Z?ʵ�>�^��./�=�����=+��6W>���>�V/?�F?�d?���<��V��jh�v"���'����}����>�'>"�>(��>琎>+ޞ���V>�d�>Y��>��>���=���<��,=d%5>/N�>���>���>"S<>�x>�̴��-����h��Xu���ɽP�?nY��-�J�mA��/�������=�:.?G�>����9п	���x�G?B����yG*��S>��0?�/W?X>���[�r�>�t���k�0C >n� ��Gl�X)��ZP>��?�Ha>s��>�5E��F��NN�����>��J?>E���a�
����I�Sæ��}M>��>�xѽ?-�3G��2�J��m��D��aB?�?~�>�ߓ����_���i�>Cs�=x2>z�X>;d���&���	�8{:���;_�>|�r�`��>�t>��=u��>�P��A���vs>)j�>�W�>>',?�*?���=3x���Ho��[�1�B>���>v�[>ѷ�=l�9�Q��=���>n�?>�HA�Y�l��)�H(4��
[>���!Ո��⦽���<U]����=�� =�ڨ�|�I����<@�?^���O��Z\�����#�>Do?S1���½?�{�򩤿ˊ�p�?�@�Φ?-A�V�r���?Vp�?�󽅧�>�?�3z>`'����Bi�>��A>s/��G�[Lվ�9�?W��?�1o�m�=�L�V��.u�S"�>A6~�0h�>�u��Z�����3�u�)�#=s��>.9H?�V����O��
>��u
?2?�]�a���]�ȿo|v���>c�?��?��m�HA���@����>���?�gY?�qi>.e۾�bZ���>��@?R?��>:���'���?6޶?��?��H>�}�?=�s?�b�>��w��/����s����=�/;!0�>�>�����HF�QƓ��n��#�j������`>��$=Gָ>~��|ϻ�HO�=e>��K����j�S��>o�r>��J>S��>�?{�>瀙>)X=mq���������֗K?���?���In�{��<G��=�R]���?��4?��T���ξ3�>�@\?r��?��Z?��>53�r�������(��?͍<�eL>AW�>f!�> ��,,L>vvԾ�B�j�>��>����{5ھZI�����G��>�� ?K�>;��=F� ?(�#?��j>�+�>�bE��9��Z�E�ǳ�>R��>G?r�~?��?¹��W3�S���⡿�[��6N>��x?/T?:Е>���������bF��,I�풽���?azg?>���?�.�?�}??|�A?L-f>�i� �׾v�����>*?�`���*J���3��s�'?\#?Ze?�ᠽ����\Uݽ�M!�F;�&?�2R?�?���Ge�潌��jF;f�b���c��M�=(K<��.>��<>&����5>��y=�,�=��1���P�&<��)=$'�>ܐ�=@Y]�k)�-=,?��G�wۃ���=��r�5xD�p�>�IL>����^?_l=��{�����x��	U�� �?���?[k�?C��8�h��$=?�?F	?w"�>�J���}޾#�ྦPw�%~x��w���>���>�l���I���ҙ���F��b�Ž�I���>�?J?��?��=��>�f1������q�K��T�0k&�q]���6��ݾ�q��sZ�}c���[?�m��>��/�Ǻ>t�>��>�z>��?L�>�ɉ>�9z>��n>̾>� I>m'>�6>��=�����N?����V/�Y_���Ҿ�d??e�b?rm�>��ʽ��p�/����>��?���?�j�>dQ`�_-0���>?���]_?{��<�Ȕ����u���~:�|u"<[<~�-<H>�½C_1��TL�@ݛ�`7�>3��>=�����۾r����ϾˍC<T<�?P7=?�N�4�r���.��op��k�Lqͽ2���{Nž���,i����Uφ�e������|�A=Q.-?��l?T٭��4�������9z�(���,>Np�>��>o��>�5U=O�޾��O1h�6������z�>8�_?qT�>�E?i�9?\cD?�:?9��>���>����?��=�7�>��?�"1?��$?Q(?�?��0?�<3>��r�8\�h�Ӿ4?1?r ?*�>�r�>s��8!ѽ����̼ҩv���n��=7cм�xҽv*�~�ټ� (>?�q	���9�����x^f>a�8?z��>�V�>H���3��l�<�-�>!�
? ��>"���Wq���
���>\H�?����=��'>��=:Ҽ�ͽ�T�=����ϯ�=��ݼ�DX�2j+<�X�=c��=+�G�;�*�:�Ҳ���j<_��>(?X�y>y�b>�?�$<��0�W��=��->���)j=�ӹ�t��^���QJV��h4>c��?���?>��=��>�$<�����e+�^���=����,{�q�?�.?��,?S�}?��=?ұ#? ��=���n��Ì������B?�,?�>O�a˾
稿�!3�Ô??x?�a�����[)�f�¾i�ӽ��>�)/�~�����*D��X��������}z�?��?�Z?�E�6��b�1����۫� 7C?f;�>5p�>V��>,�)�!�g�U��_�:>SU�><�Q?�ջ>O?xHz?�|Y?�T>G(6�P����$D��$>�uA?��?`ǎ?�x?��>&p>{��K��>� ��� �r��.��;#F=�k]>��>���>7�>h��=�ƻ�5����;�(��=��d>�`�>�`�>P|�>}v>ɐ�<��E?���>z�'��⍪�W;��H�|���s?�?�[$?t�=Qh�/G������>�¥?�|�?�,?��T��|�=�浼�ӳ�'Vy��A�>?a�>�
�>5�= �:=�H>3�>�r�>z�S��6�mu��{?	�F?X|�=��ݿ�藿'�����>>��/=�)]���������$����>�����6���Jǽ�
+�f������ه��D����-����>]z>&��=J	>��Q���
� �8; �����=���<��f����=��>�̽,����
=;I�<�e>�u�=�����j?-U,?{�?Y?=��>������5=��?��;�Q?O1�>	*a���Ҿ�S����w���&E��K��Gyc�N`þ���=U�2<增>��>0t+>M��� �3��K=��>����ѭ=�_1>� >�>�\�=�\>���=\Ev?�b��砛���\����s�'?a��>}��=�]�2A?J�>�߈��*����	�ς?k�@���?oE ?��W�c�>V,ľ�E�@�'= 7 :���>Σ�<}�Y�s̷>z�>>K����������I��?b,@�5?���}Ϳ��1>G�:>JH>)�N�o2�<�t�gW��te�)�#?��.�5�ľ�.�>���=�۾�k����l=BG0>�ߣ=|� ��Y�ҝ=]�P�F�d=~�B="�q>�3>�
�=�k����=�/R=5q�=�DM>:��Z#���
�Rh8=��=hb>Ls><�>T�?�#?��R?�>��H���޾�b���Ȥ>xĴ=��>�=Y�?>]��>�I4?��7?�L?,��>RE}=���>�a�>D��*�i�0��K�����W<�=�?ܡ�?ܝ�>':��t�����/�����?�a*?�?ٞ�>��q�ϋ&�nN���椽#v;ŋ�=�O�����>�5����z�f>���>Tp�>BO�>��@>�3�=4>��>�>S�4<��b=ZbL8�
=.����'<�:
<�3;�i�pa<=p�i=��r�|��<<K<<�ڍ=�,�=�=���>�o>i��>��=����->���ݺL�
Ż=1�����A�Zd�1~��/�"7�jA>$�U>!󅽾��
�?O�Z>�o=>�q�?�#u?T�">��0FվSG��Ane��S�:��=��
>r�<�<�;��_��N�ZJӾ���>4�>;��>�km>�,�y�>��Qq=�V�U5��6�>sŌ�=�o��1q��$��֟��9i���H��oD?B/��,T�=��}?!>I?ď?� �>P����*ؾ{�/>~����=,�1<q������?��&?���>����4E���T����!?�,���<��d����۾R��7��4=�>]5����c�7����i��������}?�<L?��?U�K����
tx�| ����#��>p3v?Z`>��>ؽ�>����;k���6��J�>��?�e�?� �?{�=���=�l�����>��?�˗?���?j�g?��;���>(v����2>���y��=�H>��=4
�=��?1d?E�?��������P���Y]��q�Ϻ	�=i�>�J�>/�U>��=[F=�6�=��`>���>>Ï>��_>�g�>�	�>�挾&�+�?�h=�=�>�U<?�?W>SF�=�F]���ɼ갳�b�S�8;H�{��{쿽,)P���-��O������<��>��ȿ���?��>1X��H,�>���º#��u�=��>��b=Z#�>�5#>`��=�Q�>é>`5�=0]�>��>)Ӿ��>��{�!��BC��ER�՗Ѿ��z>�Ɯ���%�q��y���+�H�V���B�yj�1���?=��I�<�#�?P���λk�ͳ)�ڶ����?�C�>�,6?�w��}Z��@�>���>���>֖��ϖ�������}���?���?ۜ�>�|�>rI?�?9խ�D���\�X��Lu�����Ry��RE�銿;������N��%N?�x�?G�e?�J>A�>>���?G��\vϾ#��>�F���C�՗=<��>�پ/Ԛ�������K)�5ۨ=�@?�&�?�g?��I�˿��5`>��?�n?'�?��\?2��>_h����??l�t>��4?,#=?�[?��?;,?� =�I�>��>�"J2�����Db��y���3�@��a��<89��R�c1N���9���=���=��=���=E�ʻ��<�K�:\�]=��7>�?�>.�h?k��>j��=��+?E[�	+Y������?�dg�d���Q	���
���TN= L?��?��?�>f���M���=�a{>�ړ>$��=ךo>!3������z�Q�U�=���>�c]�y7?��r�������'�=���=�?���>fc6�#����ľ�=,���>׾Ͻ�.޾K����n�B�;��P�̕
?WI^?��>������?>��z�\r]?��	?#�?؟@?A�W>��%��|
��?E�������>�G!��'�fw��mШ�H�A��B��F�=��w�b٠�/mb>���R޾=�n��J������M=p�Q�V=���־hP��/�=�
>������ ����fѪ�O&J?z�j=x��TU��`����>�ɘ>Qˮ>��:���v�|@�R����R�=��>9�:>���s�~G�>6�>��C?A�Y?�K�?2|k�V�>����dِ�Dg�<�V?Ȥ�>�c�>,#>)�=z績`��Cg�&�A�8,�>T��>0���*E�K���<��s�!��>��>�LX>��?�mH?q	?��Z?� ?�7�>p%�>�0G��G���[?^#�?��=ʑ�ڱ�]�%��\m�9�o>��>����>��>�t�>{n ?��<?�#q?��?�L<�g����l/�>Ξ|>R�T�������>'�L?���>y8?yi?k�?>�K��K޾�Xp�?=>�
�=N'B?�?ڢ?�w�>���>MW����H=w�>$�b?n�?eUn?���=��?�z.>t��>Q�= ��>�n�>�!?�nK?�Ms?K�L?�J�>%Ȍ<@���J���h����M��:p�C<f�}=*���uj�����i�<��;y�P�C��MƼ��4�$���@B<�>��D>�޶�QB)=�#��27���@>q����ȾS-���8��g�Q>l:�>g]�>t�>ؒ���+>[��>j{>1W'��O?$;�>��?�� >dSC��� �-��}�>UGC?o�ýjH��UŦ�@)���(�=��p?l�H?~�d=Yӷ�xdc?)�_?I���M�5��g�{���ݾ� r?��%?0�/e�>��]?��M?���>��T��@H�I�����l�����<n=�+�>�-��|���>ٳ[?�b�>�u>���=���7ل�#!�8�	?ws?Y-�?WP�?���=p l���ѿ�Y�{�zhc?U�>�����?���;3 Ծ�۞��؎�q���ŵ�2��������о}�=�*���V�>���>�M? 
f?Z�R?���lSX���I�����_��A	�,#&�F�>�ѧ6�|�>��&w����M微\}�2�=�D�����6Ь?0}??^�#$>�W���Q�����o�=�~޾�2w��[�u��X�:타>�;=���=��!�h/?/�>���>��,?ig��!�bvB��7Z�+�#QW>vC�>�1�>H�?�O�=~�=�	=F����׾UG=}%v>wc?2�K?��n?����1�܀��r�!�m�.��J����B>�>>���>e�W�'���;&�XT>���r�*���{����	��m~=ݫ2?T;�>���>�M�?��?\m	��[��Vx�i~1��ȃ<�-�>�i?��>�͆>�Qн� �Ĕ�>�<k?6�>^��>噾���b�t��늽C��>�u�>a��>׍J>�"E�L_�O����k��^4��x�=ߊ]?�	����F�<�x>]CQ?fЮ<���ŉ�>�����j�ߌᾑ8��>� ?�Q�=l� >W?ܾ��}�}��镾�k"?Y�?!����wR�Ʋ>�g?[��>��L>�A`?��q>�m�������\�>:�h?�V?y@M?���>$��=I&U����<� .=Q��>��c>�Z�=h��=����=�^��l�E��=9R�=��&�x$���że�{=�P=����Ź!>�lۿ�AK�1�پw	����>
�p舾�����c������b�����[x����'��V��5c�����l����?T=�??���{.��%���`���ǿ����>�q�pi���%��z)�����T����d!�~�O��%i��e�c�'?s!��l�ǿ���فܾ�4 ?� ?O�y?���w�"��-8�� >���<wq��(N뾿v���ο�Ț���^?gx�>����B��(i�>'��>��X>s�q>#���4ߞ���<
?�c-?�b�>�r��uɿ�u��;&�<���?n�@��f?�����D�m��Q��>%1�>G ?P吼����=ھ���>`;?�?Y��>�=[��h��?�R���Ĥ�Ue���>��1=[Ǌ����b��>C�K>�h�Q���#(����>8�>Ϡ�=�EB��q�����}�>��l�k	b�Մ?�{\��f���/�T��;V>��T?*�>}9�=��,? 7H�(}Ͽ7�\��+a?�0�?h��?��(?Gܿ�Jۚ>��ܾ.�M?�C6?S��>�c&���t����=�+�eG��u��E'V���==��>��>�,����W�O��+��F��=���ƿH�$��v��=���u�[���B����#U��-���so�s���]h=�x�=L�Q>rv�>�CW>3Z>�eW?��k?�W�>ŀ>SV佼����
ξ����O��&���������D棾�G��߾�w	�������Z�ɾMw<���=)R�����9"!��b��aF��k/?��&>%xʾ�M��p+<�Zʾ�����݃�u��m�;3�1��n�x}�?3B?���"8W�w�~��ƺ��_W?�N��<�~������=�Ȝ=�ܝ>��=���83�FYS�E*?U[6?MZ�_�eq�;s�c<�d�;VR?��?�w3�V�>a�?7#>�o0|�EFW>b>.>�>gx�>y�Q>�q���~z���?��f?���\g��$��>�~���;�φ�=x >ܸF�	����{>�h��^����>
�B<��>!'W?���>��)���b���T����<=D�x?Ҟ?!�>�}k?��B?P�<���}�S����vu=��W?�i?!�>���о�s��u�5?�e?8�N>�Sh�b�龧�.��M�$?��n?�W?	���h}����y���m6?��v?s^�xs�����I�V�f=�>�[�>���>��9��k�>�>?�#��G������xY4�#Þ?��@���?"�;< �\��=�;?l\�>��O��>ƾ�z������L�q=�"�>���ev����	R,�d�8?ܠ�?���>��������>�	��8�?���?w����
C;V�&��oq�~���3���b=�Z�r�:�ƾ2g��Ǡ�T���(f�oj9=�c�>A@ѽ��^��>0K$���ۿ��ڿ�Ň��ݾ�ʈ�v�?gj�>Î7���x�P�@��fg��[��I��E��B>�����$�=�=���Um��pN����=[qU>]�t��^�>�"�����ٮ��\q<��>}�?�>Ǧ��}�U��?�0A�$�Ԯ���%�N�?���?�O�??:�X>ʶ��� v�/<⧆?���?��? �4�Ѹվ�~b� �j?n_��yU`��4�yHE��U>�"3?	C�>>�-��|=>���>
g>�#/�p�Ŀ�ٶ�C���Q��?���?�o� ��>q��?ws+?�i�8��q[����*��+��<A?�2>���@�!�40=�ZҒ���
?Z~0?{�[.��Y?�0��?h~�.�>��'��ؗ�>���=�|@��ݽ�t>�R�_�������O=�?�?o�?[�	��&4�)�%?���>D���6e��*:>;A?��>�sp>�E�<���>�5���#�A'�=L��?sl�?5˾>9���P�����>u̓?�~�>,ً?A>=�� ?e���\U���'=H�>+�~>�#�e�?V5>?UB�>ڠ�6�2�����]?���K�@7Ӿ�~B����>Zw?i�=?\d>ݻ�SA=iT*�K�SY������&��!���O�o��>>Rl>e#J��ؾ��?Mp�9�ؿ j��p'��54?0��>�?����t�����;_?Qz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?W��D��u�o�x�>���?
�@�ծ?ki��	?���P��Ta~����7�^��=��7?�0��z>���>��=�nv�޻��W�s����>�B�?�{�?��>!�l?��o�N�B���1=6M�>̜k?�s?SPo���e�B>��?"������L��f?�
@u@`�^?)��¿�Ӏ��i�f����=s�<�aY>����0�=E��=�&���O�h�=��7>�?�=��>K��=�9�=�sH>`<��U��e���U��x�(��*����ʾ1�D�l��.4��-پCoܾ��8��Z����<�⌾�K�2�<���=�U?dR?_p?э ?��x�[�>)���)T=�{#�lՄ=�.�>g2?¥L?�*?{ӓ=����G�d��_��#B��Oɇ����>ppI>Ѐ�>�H�>�$�> �@9��I>#2?>��>>�d'=���o_=h�N>�M�>���>Oz�>�I>�L0>ó��
���ck��g���ٽ���?��6)G�0	��i?��y����E=(+,?�\>̲���п!���'�A?HM����]�(�a�>Ui5?><Q?�b>�F�������>Υ��_�
!>��1�k�\�"�h�\>0?ؾh>H�x>��3���8�~VQ�y���ƻy>MK7?�:J9���s���G���ܾ�hG>%��>��'�u�����a�~�� j���=�8?�`?r���e����u�	E���.O>#Y>s�!= ��=�.M>�4^�}�ý\�H��,9=ޕ�=FGa>?�E>咃=���>����9�S��>�L`> �C>G�=?�6#?��K��J���R��2�8�f]h>B�>8c>�Z>|�Y����=N1�>��r>����5����Ͻ�kM���h>�~��a�Z��}���=G�����=���<����dpO���<�c�?���Ԍ�i�����=��?�J2?�:p=*��<0�;��Ǣ��o��|`�?C�@p��?��ӃZ��+�>U��?؝�<��=���>���>!�L�7Ka�+�>�z=r-�B8��\�)�?�z�?i���喿y���>��H?���Ph�>{x��Z�������u�y�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?1uH>�t�?]Vs?~��>�,{���.�����;B��)�=}��;�"�>�?>��$dF�����ZU���j��&��Q`>�#=�޸>�3������I�=����ߧ���j��j�>�q>�XJ>�5�>� ?qy�>|��>�X=������ǖ�U�J?�C�?K����q���D����=jj��?�:?ȼɜ����>��N?�bc?�jT?=�>1�!�ٳ��y���Q��a�Y=��>)i�>8>�>��'�<>:Ѿ��Z�k>���>�<[p̾��g����;��>|$?o�>�>F&?�C#?�"w>�x�>��{����b�"��c ?ł?Bc?>H�?c�>�'����>������N���Fa���G=��L?��(?�O�>7o��>������Q��E/���$�?-gY?Gw��;?��z?f,?N�?�>�޼=7; ��tݼqRV>�	?j툽��8���M�m���w?���>�/�>Z������<�������?��d?�5?�[
�`�C�"���Br�<�T���:w�l=0�@<��X>�}>|jS�0Bi=���=�d
>),>�9f���Hs��l=�>-}> �x�٦R�/�+?��3�_ꂾ�"�=\�r�M]C���}>�WN>�2���I^?]=���{������j��'�U����?|0�?�ʕ?ky���h��]=?��?ю?���>�b��~�۾n�߾?-t�!s��"�~� >���>{�)����E��C��;r˽�3"� �>�:�>A�?��>�Y>�u�>O'~��g��cӾ�^�AY�$���7�[,��;�m��K�!�����Z;���{�"+�>�64�CC�>2c�>c�|>'^>�;�>܈<���>�.>!(g>X�>��:>2��=�=H��-߽S�P?���ȍ/�w���ɾ�O?�eb?��>���i�������S?��?���?�r>�e~�����#��>zZ�>�Ҡ��l:?��>r(B=���=���+x��Z0��gjý���>N睾!�O�I/]�FY��ѿ?-!?8����YG�ma;�C��`1�=1�?��3?f�$���J���^���D�l�8�ϴ�=�j.�����A%���o��b��{C�����3�~{D<?O3?O�}?�����]ܾ�s|�X�3��{b>	��>��>���>�3>A��^J#���Y�v���t�CA�>5�v?���>I{I?J�;?��O?T�L?c�>D�>~�����>&��;�Q�>*��>�D9?+�-?fY0?��?�D+?3^c>�3������+�ؾ�?�?84?�M?�\?zk���鿽����o^�
:x��2��$�z=���<�Tֽ"�r���P=�[T>'�?���ϑ@�	��*�u>f2?���>jg�>=���4����Sf��:�>�?au>����Tm�.���>�Nk?�-�mG�<.#>ӵ>��<�f���=�̻���=|V=��]��hu��܁=�ۼ=�忼2���-�����G��<ܿ�>��?��>�<�>����'Z��D���z�=��Y>��S>8�> �ھ1p��^���Zg��+y>�ʏ?�?tOe=:0�=vC�=���=���]���6��r�=�?3�#?�U?!Ñ?%P;?S�"?T� >\��|���ᄿg���8?*!,?���>���?�ʾ=��3���?�]?9a���68)���¾ս��>�Y/�N,~�<���D�
}��r���s�����?C��?;+A��6��q�W���LZ����C?�!�>�T�>��>��)���g��&��7;>W��>%R?d/�>lqI?�af?�vX?�>a>xoA��8ƿ�ܚ�DU�˹�y�)?"ef?Ն?�}?�o?�:>ӓ���0�GՍ��8�`(�;�-����?���>s�y>XϘ>�c�>	�=Z��2�=I������=��>�r�>ʕ_>�L>�+�>�A�j�F?��>m����H���Nn��8��s?(>�?�G%?�q!=&I�;�F�����s�>I_�?|��?�&?��H����=���[��AW]��>�>
��>�>v��=~KG=l4!>	��>P�>��������:���~���?�1B?>��=80࿃�E�C>{%�U��>(�	�}%?���;�Ѿ��]�B� ��*��C����ξ�^��^���>��7x=؎H��2�>�1�=�1>�L>{:�=Q"��g���5=�X�;���kֽgP�\}��8w<_��=p��>�Wo>�	'>�C���p��4e}?ԜB?�`$?K�Y>Gդ>�\>��>��M?�)>�8!?d�{>~	��+���P�=.��Q�~��$�'	J��`A��9��^�>�[�@>8��=���=��A��L=���=�Ϗ=b*�<_O���>�D�=˯'�MR�<;�=:��=a6w?z���鲝�R5Q��_罄�:?:�>�z�=�ƾ�@?��>>�2������aa��.?7��?|T�?S�?�si�|f�>R���$p�=r���|@2>���= �2�h��>_�J>ׂ��J��쀳�5�?Z�@��??�ዿt�ϿKb/>A� >2>4>�Ja�Й*�~]$����ec(��*?��o˾���=&��=kЬ��MȾ�}=5��=��=n��<��R�Zӹ<�Ƽ飤:��>D��>y�^>S�=�M��y+>q�=��>�K�=�m��]=?�X����S=��=I�{>�0>���>��?�"?Q2?#?�U>��M�ξ�>�5����>� �=ϫ��6��>�_?}My?2*?贈>��H>Kæ>��9>zT��Nf�����MB�� w=>+�?�0�?��z>ن	����FL��m���?!�>C?)��>딄>�U����=Y&���.�����6�4��+=�mr�sQU������m�V�㽘�=�p�>���>��>\Ty>k�9>��N>w�>q�>Y8�<wp�=�݌���<� �����=U�����<�uż����5z&�	�+�3�����;��;��]<��;�G�=���>GK >��>ۢ�<ۊ��^!> ΁���?�i1�=�졾zBD�e�d�u��x�0�Qa<�V<>��(>���JՐ��?�)E>�Q[>!�?Ze?�eJ>������Rh���[���V�阼=9}�=��]��/I��^���Q��d߾o��>)�>S�>��l>y,��?�P�w=��ᾰY5�<�>�y��u"��=�I;q��>����(i��l�$�D?�E�����=J~?��I?Wޏ?7|�>0˘���ؾHZ0>6��:�=D�u!q��x����?Q�&?���>�!�7�D��*�ؽSf�>��&�,�Iї��(+��GȽ��gϞ>U¾��ھ��9��Y�� ��ա0��%\��v�>��G?9է?����u���C��'��)%����>Kg?�L�>��
?;�?����f]���Dm�G/�=Y�t?B��??Ȼ?k��=�	�=^ ��J�>'.?�_�?*Ώ?.q?'�=�C%�>Z�;�?>ơ����=B�>�ʙ=7�=��?[h?!�?�і�@'���t���S�?>�<JJ�=���>3&�>~Nr>��=��V=��=�*l>W:�><�>ok>��>�.�>�z���u���?oE�=�G�>	?FU�>Bs=�����lu<�����K�����yܼ��ٽ��;�>R�W>�����>ӓ��)̡?ÀU>�|�3�?�}�?u����=@:>��k�>CkG>��>ʐ�>H��>�E>u�>_��>)Ӿ
�>ؤ�� ��	C�XR�a�Ѿ�z>m&����$��j�;�����I����zx��j��-��f=���<2C�?�����~k�*�)�����?�6�>��5?�݌��􅽙->���>��>~�������?����Cᾯ�? ��?{&c>g�>7�W?�u?b1�2�2�;uZ��u�H A���d�Л`��ύ�����ts
��F��4�_?�x?<|A?�e�<lNz>f��?��%��^���Ċ>>�.��>;��+;=N�>� ��B�`��\ӾӒþ����XF>��o?��?�&?��U�U�n��]'>�i:?�w1?�t?T�1?�v;?�4���$?	^3>�?NM?i5?�.?ӹ
?N@1>���=�L����&=v5��E4����нxʽX���#3=g�{=Y�Ÿ��<��=���<��Jۼ+�S;�v��>;�<��:=�E�=�_�=�|�>�#U?D��>&C>�;G?`
{��NI����??�MK� 4�F���y��82վe;t>(�~?sΜ?�H?�j�> ~)�E]��5>ޕ�>9�=A�z>���>���<*6ڽ��<=Y��=��.>���<<QD�qy��������j�iGF���>���>:�>N`���`>�K���Žl=�=?�ѽى���h��5��o.�6#-�>�^;?�x%?���=PX�����\�#A,?��&?c`?¹8?3�0�ltg����F�.�s�D=�L�>�`���G-��F���[k�Ȝ]�u�><6��4Р�\^b>����g޾�n���I��羈�M=Fr���V=��i־M,�H��=-
>F���� ����KӪ�l)J?�Xj=�\��	TU��v��l�>s��>�î>q;�s�w��@�(����o�=���>d;><������{zG�<8�FÌ>.yA?��Y?���?� ��(@k�5�T�u��(ϣ�'Z@��?A�> *?Bt>�>D��������Y�~C�}��>K-�>�	��2�/M����0�/�#�>e�?PA,>1)?��V?�?�T`?Z�$?�:�>�k?>�h,��䧾c�%?�c�?�؆=�ҽ\�O���8��PG����>W�(?D.G�֔�>?�0?|(?�HR?B�?��>����L�@�#>cF�>FV�̂����a>Q�I?�A�>G-X?�@�?@�=>_�5�A���ԫ����=7X> �1?��"?��?4��>!��>қ���d=�^�>^�b?�?��m?���=�1?!_1>���>W�=(��>]��>Yj?��M?��q?��I?@��>���<kT��|����X~�	�%� �j<�`w<sd~=�X �|�s�"�����<�4<~c��t�� �����/�s暼ux�;��>B=�=~`��(ަ>�ȾԀ��j<�%��|�پO?x�~t����c=c*>+��>P"?�> �Ge�=�e�>
W�>o��
�??�2?��?z{,>�AT�?����T>��N?�8%��m��s��Tq��m�/>��I?J.?�E���,�Rc?�\?Tr��]�=�w����3P����ՌR?�R
?hyA�^��>~?7xn?!�>'q��n�C���yrc�B�_�̮�=YO�>����^����>��4?���>��U>�H�=�sվ�3v�9���M+?ތ�?�?w��?e�,>nnr��T߿��'�JZ����[?:�>�BA���?��=�о����Δ�(a����׾=ʾu���^þa�p��ל��<���=�(?[�u?�X�?�+h?��׾m���};8��b��Æ�����H��|X��@���B�Z���xh��.�W"��*F>8�$���%��Ƞ?�<.?�|M�V��>��߾ț���>�=�����O� �>��=�>U>GM>�8���E�����0�!?�>2�>޵W?��X��HT��r��R��*�"h>u�>�t�>���>D�1>Ic�=���=���'�j��
�<r8v> xc?��K?|�n?�]�!*1�퇂��!�'�/�Pg����B>&j>ٸ�>��W�����9&�Z>�=�r�{���v��W�	�R�~=[�2?1(�>ǰ�>�L�?�?�x	��b��oqx�܉1�訃<3"�>�i?G<�>n�>i�Ͻ-� �#��>�l?�k�>#��>q���-2!���{��ɽ��>�>p��>��o>B�,�9\�-b���|��K9��=_�h?�~����`�,�>�/R?��]:_�@<���>Nx���!�D��_�'�e8>3]?��=��;>kdž��{��B�� ,&?�?c���7�)�L��>o�?5��>RȘ>¶�?	�>���L����?V�Z?qI?o;?���>��=�﬽S����t/�ϧ-=5҄>��O>]�=!��=���_�\��+���8=ծ=�^���'��d��;d̼�^�<E|�<�B>emۿlBK�s�پ�	��==
�*戾i���Cc��s���a��S���Zx����
'��V�j7c�����1�l�2��?{=�?_z���*������b����������>��q�R���������+��n�ཱྀŬ�#e!���O��&i�ξe�|�'?�����ǿΰ���;ܾ�  ?�A ?B�y?;�Ԟ"���8��� >2e�<B��G�뾃�����ο������^?��>��b7��)��>��>��X>�Fq>���l瞾l �<��?l�-?D��>�r�#�ɿL���ത<���?��@�'Y?]�u�y�:�S�����?>�?j+j>�Q��R[%�"��_,�>W�?���?>,?�[���'�Ȗ[?�3g=2.F����Ί>z)_>+$�Y�͔�>SA�>4R�<_��1v׾��>8��>d`����$���+�����>�_����5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?:ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=z6�扤�{���&V�}��=[��>b�>��,������O��I��S��=��ݸƿ�$�h����<�H�� Z��;�����aQ��<��Q�n��f��f=�\�=5R>�ޅ>eW>�EZ>vHW?X�k?{}�>�>����D���ξ���nŁ��������Et�9����,�p߾�x	����U���\ɾg=�N�=�7R�떐�?� ���b���F�7�.?�y$>��ʾ(�M��4-<mʾ����pʄ��⥽�(̾��1��"n��˟?�A?C���z�V�����$�h��ҫW?{Y�w���ꬾ^��=�t��K�=V%�>�w�=W���3��|S�T&0?_/?߿�:���T)>�����!=�	+?U� ?��< �>w�"?�,�G9޽z?Y><�.>|�>��>.�>�ԭ�=ݽ�?'�U?�8����֑>����Fy�}�q=~}>>:�����'X>�f�<-���.�dɡ��ܾ<�gg?f��>�k5�J�S�X���# >8�>�ϡ?�4�>���>�	�?kn?�G-�QX������&��>�=Y%??�9J?�m�=�>����Ņ�t�%?.��?��	���(�'2��Q�0�n��ƚ?e}?&�9?j��<�(��\1��?�E�v�]?��v?�r^�ns�����q�V�;=�>'\�>��>��9��k�>,�>?�#��G�������Y4�.Þ?��@���?��;<��|��=};?\�>�O��>ƾ�{��?���/�q=0"�>ӌ��>ev�����Q,�K�8?Š�?1��>򓂾��� T�=�Γ��p�??E#��O�b<w����m�-H��u�q<��=����)������3����Ԏ	�O��X�ּ��>��@ ܽ<
�>�A8�W��Ͽ�+��>b;|�k�5?�&�>�qƽ�x���h�Hs�uJ�-F��n���p�>�Σ<hfP>�[��Z���o��q$=Ҭ�=�޾)�?��ˎ��"?���;��d>��.?{+�>й'� ��O��?_��$��9���%�.��P?�.�?�Dk?��:?R�=�A=a�;>T��>5��?�K?�%?��=n�Y�Y�;�m?+�����h�OI1�7�-�>�t1?�?2��5�=�X>��>�S�=M�!� ¿�������w?�?|b�?�8�V��>��?�TI?�!�#��k!��?�7�rF=��A?��>�8�����G(�d�*��?~<-?nu��r�+�AW_?�]a�:p���-���ͽ�՞>��/��*`������q�e��؛���u���?���?�Ӳ?���"�vf%?�_�>΄���̾k3�<�Ф>�a�>X<S>	�[���x>0��:��?>2-�?ɐ�?��
?i돿2����T>��}?�`�>BI�?~@=�_"?w�齋������=�>��g>������>��?���>(�f�i����Ֆf�5 ��0��'U����>Kl^?>�?n��>�o���c=��X�S�K������!�҇��������j>�!�=>�=���=j���?Qp�9�ؿ�i��	p'��54?-��>�?����t�W���;_?_z�>�6��+���%���B�_��?�G�?=�?��׾cR̼�>A�>�I�>A�Խ���V�����7>1�B?O��D��q�o�v�>���?	�@�ծ?ki��	?��P���_~���7����=z�7?�0���z>^��>T�=�nv�ӻ����s�Z��>C�?�z�?���>L�l?C�o���B�$�1=^L�>؛k?t?�m�Z��B>5�?e������CK�'f?��
@]u@�^? ���h����̷�Oa��Χ�=�=">�d���5�=�iX=_������<�=(��>�W0>�z�>i�=��+>��A>�X����#��#���9���I�n��+���9��J.��RZ������a�&?�$��C���(�xi�>��
�=��U?��Q?��o?�� ?��x��M>�k����=�$$���=�:�>�,2?�L?U�*?�Ԓ=���d�LZ���<���Ǉ����>�`H>���>��>�ӭ>%�08�I>G�?>��>s >�&=�2�q>=��N>�]�>6��>���>�C<>��>Fϴ��1��g�h��
w�j̽0�?}���Q�J��1���9��Ҧ���h�=Gb.?|>���?пf����2H?'���x)���+���>~�0?�cW?�>%����T�0:>6����j�@`>�+ ��l���)��%Q>ul?:lj>��t>i�3��%6�cMQ��S���~>�<7?�U����3��s���H�_n޾��I>�Q�>B\F�C*�W���}���l����=K�:?4�?����8��]r����2\U>kY>L=��=mK>�Tw�����B���&=ry�=m�T>(�? K0>¶�:�[�>g̾/��E״>3�>�Q>BZ@?�r'?(���	�������P��xg>5��>DG�;�-�=���K!>�?d��>!�"
Z�/ƽ䏾|�o>�ݽ�r�������X=N��X8>U}�=�@/�Fzm��z���?�y���\���U��Zu�"?��?�ӽw%g�Yc�uo���/���?3�@q�^?��j�E�u�?�~u?�C�<�P� M>�ߐ>Q�=dV��j>��=�ń����>��*p�?@��?��=zꋿ��q��>=W�
?ڹ��\�>Y<��ߘ�4���ٲ��W�#<��>ֽ.?��	�!ރ��}��?��?�b�����g����{g���>��?��?VSx�����5��1�>c��?�V?VɃ>�����������>��J?��g?2L�>��"���k����>���?��w?�ZI>rU�??t?g��>��o��D/�����b���%u=�;�6�>���=Fh����F�o��$��si��R�c>F�#=�>�+�;o���=���i7����m���>�3p>��I>���>D_ ?��>T��>D=�/����� *����K?��?���.n����<yM�=�!_��?�<4?:�_�I�Ͼ4ި>
�\?�ŀ?�[?M�>���.-��㿿^v���x�<��K>���>�:�>�Q��[+K>��Ծ|3D�~�>̣�>Ɍ���.ھ�\�� y���6�>Ba!?݀�>˭�=�� ?��#?*�j>�(�>�`E��9����E����>��>�H?{�~?��?Թ�fY3����q桿,�[�2@N>��x?�U?+ɕ>��������qE�'SI�쒽>��?sg?oO��?@2�?$�??��A?�(f>+��^ؾ����[�>��!?aN�C�A��0&�r�Wd?)�?ip�>~瑽!1ս��ۼ]�������?�[?�%?`[�Ւ`�%þT�<�*�7F��w�;��A��>��>~q�����=Tg>��=gm�5~5��y<$��=��>���=y�7��{���G,?2�F��ڃ�M�=��r�VxD�>"�>��L>�����^?H�<��{����kz��"�U���?w��?�n�?�~��M�h��=?r�?[�?��>���"�޾~(�c7w��jy� W��>b��>��l�2徒���7���R4��j�Ž0�ӽ��?i�>XQ�>)��>�"�=�E�>:���ޮ��F!��}��%&��&O�Y<����A彷�H�b^սHۗ��h����>�Ԗ�� �>�?��V>��>|��>X�=Zy�>�A>��o>ڈ�>��u�S6>��C>;��6+`���P?
����K@�mI"�Pm1��#3?k^L?Z�>iI�=#������J?7��?^	�?���=Kj���Ҿ%�>��>8����M?z�=��0>$��=o:��|���s���ܰ��r�>�u����@�_:W��پ#(9?�7<?�� ���r�R��2�о��=���?\�1?����MT�?Q��lL��lW�-ƪ������ھz�)�ڽo�O얿�Ԇ��.����/����=�-7?+]w?����ʾT图����f+�N
 >�;>>�0�>���>��	><�*6��Ed�$V�[�i��E�>�M�?�ɍ>sH?>L<?&@L?��L?���>;��>)u��Q��>V:Xm�>V�>!s8?��-?�1?��?�(?�Vm>- �������ھ�?�?ҕ?��?�?,����&��k(��o��}܁��l�lX=���<��ս�Om���^=�/_>�Z?�<�<�8������l>�O7?4��>�f�>���
��R}�<|��>#�
?$��>���>sr��W��n�>��?�w��;=o�)>Q�=Z��U;?�-�=󱽼���=�i��z5:���!<�ڿ=2t�=��z���d�V);�};2�<�F ?�?Ƨ�>_�>�冾�� �����M�=��X>9�V>؝ >��ؾ-Ċ��7����h���>�U�?��?�.[=�`�=z��=�4���F¾H�����y��<� ?��"?�Q?��?V%??;�"?�>�=�1d���ą�?d���U?�{,?�:�> ����ƾ�ר��,1�q�?�?��^��N	��&�R[ľ(޽�=>�/��|��K���$G�R����A��Z��#�?���?Y6b�$�8�����嘿}&��M�A?$�>��>��>�1*���d�T��,8>���>t?N?h��>��$?��Q?o?k]�>W���\ؿ#��З@��,5�v4G?�-?��I?�/�?ʌV?��1��h꾗Ȕ>XТ�=*�l�9�!^��A�L$f>�" >�(�>�z>�w=#k�=A%���퉾ֶ��@�<�>�JD=��]>O,�>��>-/T?�c�>�?�����:u�������Vr>k"�?+z?��d?�n>���7D\����3L�=�9�?���?-�*?R	����6>RZ��;�'>�O��>�X�>L]�>D}�>�?�=9��X?�?����������=�*Lͽ�]�>��o?�g�;�ſ�Eq��Op��8��h�r<AŒ��lf�ٖ�v�Y���=��������69[�礟�RҒ�\���R͚��z��k�>M��=�F�=���={0�<v�����<��H=pj�<:=��o�c5]<]5��R��+
���u2�Pqb<2�F=鸻x�����?�n�>GJ�>#�?��2?6�>�v�>��o?2xŽ=h-?��[>�3о-������S��d摾q̾���6v� ց�u�=W-���=��N>w��=�<׽��=�l=�f=Ö�<���<
��=�Ӌ=ݛ�=��>-T>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>q��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�T$>��#>ɧZ�ޗ%��_�4*A���F�J�?p{"�o����5>T��<w�ʾ�μ��Q�=�=(>���=��t��3e�=�=o����=��(=�> ��>6�=Q���B�>3�=�={�%>$�D<Eۨ<����/�h<2�>vC'>>���>?�1?|oU?���>��y�����ھ�w>�>/�>��Ż	M@>2��>��;? K3?;.6?(p�>O'\>R۸>x �>"�$�
A�Xhݾs(¾���=�^�?��l?ͥ�>�ª<�^��M�+�E�1��}ν.�?�'?L��>���>M|�@�#�n#���ξ�����K>�L*�k:��]B>.����C���>�F>a�>!�?y'�<�	o>��n>���>2�6>���=�S�=k��<W��<�ȫ�26�<H�
>�>�׎��5������齚:�7�;=����i��u=���=�;�>�^>M
�>�=�ɾ��*>�y��q[M��a&>�����Q�rf��Ă�e!���>�H�i>��>e|h�� ���A?��^>>��=�<�?e�|?E�>8𽡯ɾB���nzz��_�����<��n=���m�7�6�K�DnD�՛ �)��>���>���>0�{>��+��7>��{=C�ݾ˯3�z��>�҈�X-6������n����B1��ϖg�5ȃ��VF?~���
�=R~?h�J?�k�?`��>�\���~ؾ�m,>6�~��$�<w�2s�B ����?~E&?+��>v���F�5i۾ ̽1n?��2��d������=���VO��B�>�U�v���-�f���G̗������>���r>�[P?r�?�ګ��P�w
(�����[�]*�>��,?��=��2?�?YT-�a�x������F>�5�?�s�?Q߸?B�C=^8�=s>�����>��?���?�G�?��q?��<�<R�> �;��>�>��A��=�$
>���=�Y�=:�?%Y
?w�?�z��G�	�&���PC\���=�'�=r7�>�B�>�Sp>ʊ�=��g=C�=Ea>���>���>7�e>�5�>��>G���r �8�> ��<G�>�:?�r>9^=����WP@��5F���n� ?�6D����)��T"���&>�3�=�)B��+�>\׸�A��?=K>}'���?���%��¨�x4,�9��i<�>WG�>S�>Ĵ�>�>��f>��C>�E1>1Ӿ�6>/���a!��6C��}R�q�ѾR�y>�ɜ��%�>��[{����H�"$��S���i�#��!=���<�H�?Ֆ��Q�k�h�)����}�?�j�>i6?����#���8�>��>��>�,�������ȍ��o�3
�?���?QvS>|��>�^?)1?���\�)�T��Cu��	H��fX��e��i���&�����?ڽ&#`?��u?>F=?�=�}�>�0|?|;!�I����!�>��*��=��a=>!�>���8^��yվkr������y_>{1r?�p�?�T?�[u��νE��>�f'?=??J�`?z)K?�K5?��P�=�@?zE>�
?%!?u�?�?[N ?x�9>�k=�'���l=�}V�Df�����Ps���-<}�=��R=����r�<�=�D�ϳż��!���<ٯ�<���<t7,<�̠=�<�=��>�	R?E��>Du]>��6?�Y&�MD�W)����$?��5=�|�>6���ѓ��y߾�5>Q�W?�0�?�fa?��z>g3��U��e>aH�>�n>KNa>T��>�@Խ`�,��8�=��>��=�Ϡ=�!H�����Z���`΂�
�<EdW>��>OO�>�k)=�Ј>~ӟ�4���c�\>m�h�L�ξ ��>M��=��[���o>ҠN?,?���=C:��b�< �_�ȱM?�O4?q�?��n?��$>�+���A�"�*��|�-7>������t���ȣ�c�1�d�=V>g��⠾Rb>���W޾��n��J�n���L=}���V=�"��־�P�6X�=S	
>ĳ���� � ���Ϫ�.J?�j=(l��M=U��]����>Ƙ>KԮ>�7;�vw��@� ���58�=���>�;>@h��W��7xG�r4��C�>��C?w^?l�??g���Zq�1�E�ch�$-��;d�+�?V��>�+?F>Ύ�=�h�����9�\�W�B����>w�>�`���D�"��j�꾴"#�i�>^+?�& >d?,X?Co	?��a?��(?W��>���>w5��,���A�?��?E�=�*�5�P���(��c�,a�>�f?j���>��!?�?�}+?(ME?CW?(�=L���)�-���j>A͆>�q>��鬿b>�|'?~5�>��7?�?h?�J�>��J�o���[<���.>�=V+,?��?=J�>=��>��>������={��>�c?/�?��o?u}�=�?�62>���>9��=6��>���>y?VO?�s?��J? ��>�ҍ<9>��$"���(s���O����;\H<��y=ٟ�ft��.�ڨ�<��;*\��p��Ƚ񼋶D�T��q;�;_�>GuF>�Fվa�G=5����?��O>�w��K�׾�����~�zD>���>w��>��w=QSӽ��>x^�>�jN>��-�>�:?\�>x��>1$F=�Ur���۾;�V�>W/?��p���i����%����N=ql[?�H?�(�h,|���a?�:]?J4��L�s���\���Ǿ�\?f>.?Ɠ��o)�>Y�j?5�X?,8�>CQ�Ɩ`�壿��p��G۽��4=�%�>���85�ɩ�>��?��>ؘG=��=����r��ož��>�D�?A�?@�?�F�=g���i㿙�+�Z��J�g?:��>�ҿ� �>I�ڽ��Ҿ����6Vl�wM
�1�����?d���@��v����_�����C�=�A?�r�?�=�?l�q?E��;����n-� ��$�a��ힾ<�L��b�oF��2]�*Ɣ���o���C���;�3��O���?�'?��l�&$\>��þ#�	�K<羮6W>[ɾ�;5�H-�<�@���=��X>7c��ߞ���v���%?7*�>Ӏ�>��??��I�z��OL5�DRU�c/%����=3q�>@�>�"?�T>��=M�=�z��G���ٿ��iv>�Wc?��K?�n?�� ���0����՚!�A�/�����8B>��
>z��>��V�D ��&�Y]>���r�2���W��%�	�4+�=��2?���>��>.^�?�'?)�	� ���x�!t1�g5�<���>hi?-��>a��>��нM� ����>J�l?VJ�>Z��>�w��_!�
�{�*�ɽ3m�>���>���>��o>�,�U#\��X��fy���29�f�=R�h?������`���>�R?Ĕ�:0�C<p�>�6y�T�!����(�Ì>ci?@ѫ=��;>a]žb:�U�{��\��,�?&�?E�n���E���>�j?aʈ>X+>i7]?[�>�8�����k�>Ci?MI=?�/?�F�>�>�<?��5W�G=�s>�&�>g��=�!�=�|�A��L��C�:O��<������V����<5����ͻ�k���S>�yۿ�1K��ؾk��q��
��<��/��8+�����埵�j����y�2���r!� vT��c�w���V�k�0r�?*2�?T��Ј����Ā�nf��yѻ>��r�]N������ej��K���:�~��W!�t_O���h�f�e�Z�'?񺑾ڽǿѰ��^;ܾH! ?%B ?�y?��*�"�˒8�Ʈ >M�<$'����뾪�����ο%�����^?���>��0��\��>���>r�X>�Hq>���,螾�+�<��?7�-?��>F�r�+�ɿc����¤<���?�@��h?1�d���4�P�>�V?���>��?H�=���0!���!?��?޷?X�?^+���K��,�?&�F�.����������>��r��ݽ��P��o=�=�>����������M>�iK>۴½� ��h����?>l��>#)p�vZ��Մ?�z\��f�,�/��T��#V>=�T?4*�>$6�=C�,?x7H�}ϿZ�\��*a?�0�?��?@�(?ۿ�ۚ>u�ܾI�M?�D6?r��>e&���t�3��=ἧN�����&V�	��=H��>�|>��,����O��O��N��=2���ƿ��$�fJ�M =���	�\��N罎z���T��D��x�o��&�f=^��=R>+2�>��V>MAZ>�W?�k?�!�>Y�>�W�D"����;�.'�ɘ���H��p���k�7e��-���=�NR	�ߣ�����ɾ�=� �=�9R�����~� ��b���F���.?oo$>R�ʾ�M���-<�kʾ��������Hߥ�/̾C�1�� n��Ɵ?,�A?����V����H[�o���U�W?�2����묾�}�=ư����=�&�>���=��3��wS�e*?�?҇�����B�>�>���ѻ?��?�}��d#�>�?C�(:���^Q>ƻ9>�\�>�Ƽ>�n�=�����y��޻#?#3W?Q7"��@þ�_>�]ѾǸ����=95�=n�h��ޗ��)�>�R~=�"T���º�V
������X?>j�>�>��R������J�>���=ǿ�?9'?6s>B��?b� ?��R;��'�����-��g$?&es?s�=���=Q��Cg��.":?�^?}">/�]����=��w�a�޾�!?���?K�?� ��2��F���_n>��m2?*�v?4O^�)`��J ���V���>v*�>���>��9�X�>Tu>?-�"�]4��P����L4����?6�@��?6�8<'���=�[?���>|�O��jƾ�״�����;�o=\�>Gg���?v�$����+�ҽ8?���?eu�>�����b����=��P�?_�?욪��Ic<��Ol�gv��D�<ƫ=Y�M"������7��ƾE�
�ys��C�����>�Q@���D�>pR8�b��KϿ	���о��q�q�?/ͪ>�Ƚ�O����j��Au���G���H�󖌾.�>Kj�=^�=��$�17����?�+�O<X�>>��X�д�>��,��;dS��+�=�\�>EY?O�<>���l���?#��f�Կ{����)�j�t?'��?e��? �?�
:����D�?=v$�> qI?j�7?[	?����sN�U�]=��j?�U��HW`�W�4��CE��4U>�!3?�I�>��-�Pa|=�*>
��>:`>�%/�>�Ŀ	׶�S��� ��?���?%p���>?�v+?nf�a8��(V��G�*��,.��7A?72>˔��N�!�H&=��ϒ���
?z0?u���5��"B??�I��%�.�����ƞ>��I��2�sb���w<�\~��=���8�s��?N��?���?�S�,��d ?���>lK��]����A�@@�=�$�>d�P>?<<UQm>p
��W���m�>�j�?�S�?3�?����2���"�=��}?ۖ�>Ḧ?|�I�?0�>����7B��^�=%�>̲�>�Au�e ?pM
?�B>al�S����j�`�ш��d���M��Q�>V?��F?�~2>'9������ľ6�J��z$�w������:�ȽO�p>���=�`�>�Pǽ����?{p��ؿ�i���n'��54?���>�?��9�t�����;_?�z�>6��+���%���B�Y��?uG�?+�?x�׾iR̼M>��>uI�>= ս���/����7>p�B?^��D��9�o�	�>���?�@�ծ?�i��	?���P��Ra~����7�:��=��7?v0���z>���>��=�nv�λ��J�s����>�B�?�{�?���>
�l?q�o���B�c�1=M�>��k?�s?Io��󾰲B>��?�������K��f?��
@ku@7�^?����ڿȸ��0����$�����=�K9���a>��`�GF�=A�>N���4�S�h�o=A�?>��!>}�P>dJ�=r�>�>�����)�L������03�X���iӾ�{�PsǾ�������H���r��.�0�yiD���;C�r���<�	n��.�=6V?gIQ?��o?�( ?	q��W>�����=}}$��U�=4-�>؂1?(nK?Y�*?���=������e�>2��y����i��`�>-�F>~g�>���>R�>g�A;�fI>�a@>Q��>���=1)=�	��=�1N>�N�>�v�>@�>�C<>J�>:ϴ��1��B�h��	w��̽-�?р��^�J��1���9��馷��g�=6b.?�{>���?пI���u2H?����=)�$�+�}�>3�0?�cW?��>:��f�T��9>����j��`>m+ �/l���)��$Q> l?�u>�Ԍ>�3�V-�b�L����o%�>>�5?���}_f��c�� G�]���<.>�ͺ>B-�>�'�����2z�����ǰ={W9?�?ս�h˾p��(����>X\e>���9��=�7>�z�������G����=Z+�=�&>A�>�">�Y,=��N>������t���|>[�8>u>w4-?ו?�&����ϋ��#���>7h?�ʲ>�=��罝r�=ƽ?��>M "�>Q��FFy�Gpw����=�="�qIO��
X���=��M��{�>&� >���}5��>��?��������]��I(��}L?G9.?$�t=�DQ�"��7�����]�d@�?�p	@W��?�}��XT�3d?���?�KB��F/<̬�>to�> 3ƽ  1�]q�>��=݃D�����v���?�=�?���<	ǈ��^w�dk,>�8?\�3��>v�v�X���f�Oʓ��;�=Z_?��?�z� C)��_����?#_,?����֜��_f���cn��T�>�a�?���?����胡�ٵ)�sX?��?T�q?�>����� �����>�M?�`?�w�>�.@� ���@	?��?�c?iJ>�!�?1�r?��>-�b�rE.��N������i|r={��;f�>�$>����C��̒�'ш�C�i�*��[�c>�]%=Ӧ�>߆߽�!��Y�=�b��Y���m���>O�r>��E>ӥ�>b ?��>O��>J�=K����&�������K?���?����m�c��<�C�=�+]��I?��4?8��Wξ��>��[?�M�?P�Z?�-�>�n�܈��V���:ᴾn�<چM>*��>J��> |��(�J>�xվt�F��<�>���>�����۾`���|����>tj!?b��>�	�=� ?�#?�j>�"�>|bE��5����E�l��>L��>bF?#�~?��?�չ�OZ3�d��K⡿��[��FN>R�x?T?[Е>ɏ��w�����D�t�H��������?]ug?ޣ彗?/4�?�??��A?� f>K���ؾH���#�>L}!?��
�r�@��A'�>�
��t?��?���>�푽�yԽ�Mż�]��|���p?1`[?�%?���U_�h#��=��<)qJ��@~���F<Lj"�j�>:�>�)�����=�>:?�="o��r5�� �<j9�=z��>��=Hw:��팽q),?�D�����L��=W�r�y|D�zo~>��K>/���-n^?�v=���{�5笿�Z��n@T�@�?���?>k�?�P��4h��+=?X�?�K?Z��>�-��0߾�9��x���x�Y/��>��>w[V�S�㾅W�����|*���!Ľ��*�I�>�
�>sv?Q��>�q	>�4�>P����$���� ,���`�jj�S�9��^,�A��'v��������ض�[�q�Ӆ�>s���>��	?#i>geu>��>w����>4�@>��|>f<�>��c>4W>�>^�h</��(�W?P�羪S.�Xξ�9��
A?a`k?��>t���V��|��\:?R�?��?<�=�~p� ��yH?c��>��h��o	?�}_;v���2�e>��᾵~�������-�:%V>Ȅ��11�t�T��qO�`�>�-�>�b�=Z���_�>����8S=���?)/?�0�++^��i�c�[���Q�*�;B���T)�Ju�I/���,���$����'	=D41?#�?�k�?�׾�ũ��s�K�,��:>���>;��>�ɠ>�>>����0��^���&�lu����>��q?���>��F?:?�PA?��O?hi�>���>���[h�>_�<�/�>�;�>�83?W�3?,..?��?�##?��q>e���#���ݾ��?�"?�?�5?���>�{���n���ҭ��肾K�m�1�=�'!=�.ٽ$����={�g>�:?�j�����5/�\(�>hO?��\>�>><²��Yh���=Fɬ>	��>�E�>�w��xjM�P��qh?�w?�K�RW��f�V>/�'>��=@�=�i'=<]A�,gq=�o<!�����7�=���=�!��Lݐ��TY�����\��܊�>��?Ks�>�Ո><����_ �����q�=��X>`#T>��>�Pپ�z���#��a�g��hz>j�?�_�?�h=���=���=���+���W����y�<��?�S#?��S?��?�
>?��#?Ї>���B���Q������? ,?g��>���ˢʾ�訿�p3�B�?�]?Za�R�")�ě¾�ս&�>�K/��~�	���8D�����&�����?�ĝ?'B�H�6��h�d���8��=�C?���>WO�>?��>��)���g����a;>>W�>X�Q?;3�>A�5?b�P?5�"?�Nm>H� �ȸ���$j
��嶽-�G?��x?��R?S�x?Kw??��=�UX��-ʼYހ�y�9�!:Ž��_�Y��<-wd>�ϡ>i��>5X�>u�R>\��\;���z��[=��>�e�><�>
�&>�;>Un�<�G?%^�>�_����`+����Mϊ��<�?x�?4H?ɏ�="��X�d���>n��?(7�?�h$?�d��(/#>�f�=���$ľóV>DY?�۳>64_>B�G>V��=$��>^�?�-���=��oB����9�?��(?ƃ�=��ƿمs�Z�*�Y
L����p)���d%���w^[�]T0>G���|;������w��i����������F��n<a�E.�>7O�=�@> ��=c�`=��p��<Y%�<�1��6�<oL��֒<-O,��:��d���;Cj`<b_�=��B�S���:�?���>�1�>K�&?R{�>��=�2?��l?�K���!?��G=�[��3�(����>B�����Sz�� f�]3e�����o2>�w�m�>�[>
Ϭ={�˽��=�h= P�=I=.ܱ�w�"=9��=/�2='O(>��e>Hr>�6w??�����4Q��Z�[�:?�8�>N{�=j�ƾR@?)�>>�2������yb��-?h��?�T�?[�?ti��d�>����Ꮍ�s�=����p=2>���=K�2����>j�J>����J��<���x4�?��@��??�ዿ��Ͽ�a/>$�>��>�Rb�lOX��:��e��6�����>�����
�9=M/�={Ȯ�=žo󈾕��=���>I�=�:M�%�5�hD�v~>��:=ѹ�=��>6�=�^=ї>s�k>��*>� �=P�1�wBݽQ((>6�=�Ez��o�>!n>���>3g�>	1@?�B?��><�����Х��-�>>S�e>ˇ>z��@�Ƽ��>F?��K?�?�1�>��{>[!�>�%A>�M1��V:�"��_L�j��>�~�?�MU??���=ܞ ���
��)W�:�<���&?��?m��>6��>����ۿ�{���оHy;��T�R��>����kv=�a?�>�*���ݼ���=ۂ~>���>�ռ��)>Q�7>��>s>&�>��>oN��.c=a�|���]F#�Ur=��R=������5�{=�|>�o�<�=gE>��K=���=���>m`>���>	R�=b��% />z���$�L����=ZH��y%B��*d��>~���.�c!6�g�B>yHX>W��s-����? �Y>�U?>p~�?�7u?��>4��վ�Q��q	e��6S��w�=��>D�<��s;��T`�B�M�j�Ҿ���>��>��>ψl>L,�D?�� x=$��B5����>c��>3��?�#7q�7��v퟿Ci�ԯ ��D?LC�����=�$~?��I?؏?CU�>����֜ؾ-�/>�G��'b=9�Hjq��ޒ�j�?�'?���>�0���D�����ѽ��>㑽�@T�n8��Be��8ֽI�Ǿ�D�>�P�1K����9��
��`>����8��a�F��>s�>?�֪?�Y_��di��7��׽��?!�O?r�f>?)�>s��>�����Ѿl4�i׽=x$k?�&�?���?��=Ƅ�=�����>.?`ږ?~"�?��o?a�@���>���;��>e������=Gs>��=���=
?�o
?%a?�ŗ���
���1g�e�]�8�<}_�=R��>�H�>/)v>[��=tZd=���=�[>�>P�>�a>cK�>�>�p���t�v�&?:��=g.�>G1?MZ>r"=K}����=m�^�}SK�mK,��0u�C����H�<�Zk�R=r=s\��c�>��ſ
��?%�i>��!D?���b��{�[>!�_>�q���0�>�t?>��y>g�>{�>h
>�?�>�@;>�˾g�>�	���.�K�R�O��ž#�`>c���O��(\�9
ֽU�)��/������@g�������<�w"=�ё?�(���q�xy'����o�?���>�M=?I[��w�����>mL?{ܞ>UW���9������ھ^ �?���?�N>�>E~�?x 1?�]�����/�0��\J��G�W*�� ��v㝿�Z~�U��+x�xv?�W?5S/?+�h=u �>�gD?�6
þ���>���ƢT��g���PG>��������Q�ž?@˾Ih=���>�|r?F'f? "�>`m9���^�.->�9?�+?9t?�y0?�5?g��a�!?hT3>�?!�?��2?T�/?Q}
?6v->c{�=��G:pC=�t��#���Ľȵ�᰿���:=��V=z���6�}<f'.=�c|<`����Ƽ#��;(鐼V\�<�[;=3��=��=�B�>:V?	S�>̆�=^$'?�['��>M�/�Ǿ�?�a=�BX��M���)��̃����#>��\?�B�?Zb?�ċ>��-�e�r�&2�=��H>&�N>��`>]��>�]��t@C��ɻ=�c�=�ڨ=+�*=A�Z��V��{����|sA<4EL>� �>[�a>D��=�>�$����%�pv�>����^۾��c�E�G�2=�n�a�^ǩ>�IN?w�:?��<o&޾�ӿ=9�X��n1?�I?-#3?�Y?���<W?���\վVP�A�u�hޟ>��W���h��|v������b�=6�t>���m����
^>$�	��۾�Am�M&I�à�ب4=�����8=a��57Ծ$�~��0�=�<>ql��x!�cC���Z����I?�{=	���Q�U��ջ�K�>z=�>�:�>� V�\�}�>'@�H�����=��>%6>7w�X�� G��W�*u�>ڤD?�G~?�P�?�����To���3�8���>����<��?���>�>2?>H>@�������+��]{��0��k?���>�1�
E$���������7�xJ�>#�6?1�>1m$?�v'?bs0?C�{?}Q?4?L@�>]{v����̘2?��t?��p=�E�$����B�wI�0�"?A,?8_�G�>��?�j5?��8?�)8?��?&�d>�2���Q�zR�>ƝJ>Hg��i�����>t�6?��>�+p?�?Wh>je8�Wҗ��o-�x.�=�E>jH4?%�B?�D??٨r>��>�'�����=���>��m?R��?&΀?��=�?>��>pxN>���>��?��?�G?,e?_E?���>��=�	���T����������<��W=���=��������=jw�=.��=��<{�<��s��x���.SۺZ`�>�s>���B�0>G�ľV���@>�ߢ��N���Ԋ�O�:�߷=ǈ�>��?���>b#��Ւ=�>9>�>����4(?��?n?�U%;��b�n�ھ�K�p�>	B?K��=��l�儔�T�u��h=E�m?��^?�wW�n#��P�b?��]?h��=��þ��b�ω�t�O?2�
?�G��>��~?t�q?q��>-�e�(:n����Cb�0�j��Ѷ=*r�>_X�S�d�q?�>b�7?�N�>��b>�%�=Fu۾�w��q��`?��?�?���?x+*>N�n�W4࿉���9���U?/{�>�R���?"?�<ռ�CоOg��(���4Ͼe���󘾼΀�ܪ��������/�A��p�=�v?��r?��o?�U^?D��r&^�N��v�\ h��0�L���!��?���E�Txn��~-��I�)���ϼ�B]�%H�k �?�?
���+7?e���muξ>�����'>��~�`�G�<`y=�v{��t�=�o�=�u��K�3��I�?��>��>��L?A�[�!&@��l0���2��3�rC
>�N�> H�>�F�>h�h��5��_�R�37žʈ�~&�g�>�$a?i�X?���?2=�=�f&�b^t�^�ݾ�$$���-w>AH>�c�>	t��9��m�A��ZD�%&j����gN~����2�>�d?=�=:[�>\<�?u�?�W�AФ�M����FZ�E�=�i?/�d?���>i�m>��н;�A�>��>�? m�>Ж�>�ϯ��(?�F�� ���:/?��>��:?�a�>�2��&_]���U����P�z�=Zր?)]�/-��L.�>��W?��=��=Xά>�� �#���+��}w�vM��,�>ydF>���=��ž����(l�����{)?t�?�ؑ��)��"�>p�!?q6�>_�>1ǃ?�ڝ>Wn���z�;�/?�_?��I?۹@?���>��/=2����Ƚ��$�6�.=�1�>�[>H�y=���=���
Z�3����Q=�9�=�~̼�Q��( <ט����N</��<�>4>|�ڿ�K�l�վ���ba�3�	�Ҝ��	0���q��n��8���
���H�v��d���/��WU��e�����y�m��0�?M_�?�ޏ��.��Z♿�*��i�����>{��d������������ྋ¬�z5#� Q��i���d�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >VC�<�,����뾭����οA�����^?���>��/��p��>ݥ�>�X>�Hq>����螾k1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@ҨA?�f(��H쾇\Y=u�>�	?|�@>u|-����(P��I��>�:�?G�?�U=|WW��)
���e?��4<��F�[�6�=R<�==��K>��>����@�A�ٽ��4>�j�>�*'����	x]�*��<ql]>oCԽMӓ�oS�?�@!��T��~��V~��ǳ>**?�>��ؽA?Vl�6Lпn�V�|Ed?�?@���?�2?
��6�2?�Ǿ��'?�4>?���=m'2���6���"<����;��ҾaJ�'��>g<�>$n�3!��6��g�iO�=VM�=�J��c�¿����3!@=��мC5��y�$�1�P��k�����H��G,��~/=P�=�Nk>�4x>s�!>/P4>tO?��v?q��>~�i>�eĽbʙ�g��%��(��=��`R�g�پ�@��Rܾ�����%��z(��J¾� =���=�6R�:����� ��b��F�v�.?�v$>��ʾ��M� �-<Rpʾ񿪾�ل��ॽ�-̾�1�#"n�P͟?j�A?������V�d��pU�����m�W?�O����Uꬾ���=]�����=�$�>\��=\�⾓ 3�5~S�N�B?%A?�L��ʗ_��|�>H��P|ɺ}�H?{�?��>�s�>o�4?�����s
:��>��u=7
?l�?�}P<�ʾՁ<[�(?��O?�۪�	�b�>�	 ���W��-��de>�z��%���Ga> ���z�Q�&�{�T~�<��<��W?A��>��)����#����/���4=v�y?A[?b�>l�j?�C?�<�<���KBS�X$����=&/Y?�g?��>��y��$ξL�����5?�?e?�O>S�m�it�d.����s?�Cm? �?���y�|�)���6?�v?�r^�\s������V�d<�>Y[�>��>��9��l�>�>?�
#�pG������PY4��?��@���?��;<7!���=�;?\�>ݪO�{>ƾ]z��-���ؕq=�"�>)����dv���GR,�@�8?���?0��>ޓ��>���V>�ם���?=�?�.վ5��=���wd��n��Kٔ<�BM>4婽Rd���9ܾF�-���Ӿ������0� �w8g>!�@@�۽��>h�׺������ɿ�Ԉ�L� �~Ma���-? �?��I�l*�!�����{���S�j�!���w�.Е>�]L>Kp�쇾K�����B���`�_��>&�w����L��;���-Ož�.�<��>��>�Q�>'��=]U���c�?�����'�� ���p?[��?:k�?V�?�~����� �l��y�e?2s�?zՙ?�	Q>�f�dh�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�h�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�Wa?�nP����-m?�e�OP�>=�(�&��n^��qü6}b�Y���S������?gl�?��?"���5�s�6?�ƭ>Q���FW�����+ʿ>|�>��=g�i�[7>8�辽q4���>��?���?y�?I+��c��m�=��t?)l�>�Ã?#>�"�>u}�=+���?`�4>�@W=�G���W�>&.H?e�>
��=��I���4��nG��R���	��m=�:�>��^?>WG?��J>�~ֽuu�9m"����k�ｘ�����f�_����P?>�,>��#>�^]��]¾��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�-	?7�,P��X`~����7����=��7?�0��z>���>��=9ov�ܻ���s���>�B�?�{�?f��>a�l?ڀo���B���1=�K�>e�k?t?8�n�B󾯯B>��?������K�� f?8�
@yu@J�^?����ҿƥ������o���#'>DtG>���>1��`�=�;��w�;��<QpV>�%�>W�_>a�p>��>Vg>,�=*��c%��?��;,��]�;����Κ��m�!�-����pޮ����$>�������Į��޽�0:)��=�MQ?3�H?>iq?�
?D��m4>�����<�M���<=]q>Ҕ#?��??o,?��=�֪�GLd������������u�>�K)>4�>���>�-�>"�}<17D>�.Z>TF�>��>)y={C=��{=�V>��>���>JT�>wC<>��>;ϴ��1��<�h�W
w��̽�?Y��� �J��1���9������mi�=Rb.?V|>���?п]����2H?S���a)�^�+���>��0?�cW?̝>�����T��:>���s�j��`>�+ �nl���)�s%Q>�l?�f>�u>D�3�
_8�}�P�d��Z||>c!6?�涾:$9�"�u�αH��kݾ�@M>�ʾ>H3C�:n�D��� ��li��J{={r:?�|?�E��wϰ�@�u� 1��yXR>�,\>w�=N�=�YM>��b���ƽH��A.=���=U�^>�?P2>�q=�9�>u2���Ss�̜>��>Bx7>�(J?!?�o�P��0�i�s�-��[>���>�ԡ>�9�=�U����=���>-g>F'���/�I��/v�?�n>�'~�eT�I���B=x���9�=o��=_2��BQ�v�x=�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?�q>�^�?�U[?��>�V�=p�J�f����Z��ʎ>��=n-?L��>ֵ��f����ᕿ`���4u����_9�>��%=?s�>&��G ߾&��='E%���z=#��>���>\��=u4�>�:/?*�>q�`>�a=�Hm��;~�<;����K?���?*���2n��N�<X��=&�^��&?�I4?6k[�|�Ͼ�ը>�\?j?�[?d�>=��O>��F迿5~��@��<��K>'4�>�H�>�$���FK>��Ծ�4D�gp�>�ϗ>u����?ھ�,���R��EB�>�e!?���>�Ү=2?C&?�+s>���>)r>��j��Y�J�<�>|��>k?Ē�?��?����4�8�3��9����<]�ȰS>\�v?vO?�1�>���mќ���<������Ͻ�_�?%�l?����R?'V�?ό>?Ql5?eN>�����;zi�4݆>�_ ?^�
�b�A��
&���~	?��?U�>VԒ���u�����J���?"Z]?�-'?�2�!v`�J�þQ��<j�[��0Q�7(� ��<5#>� >�pZ�$X�=�@>��=�r��2����<=���>L��=�R4���b��F,?�F�ڃ�.ɘ=Ϭr�l}D���>��L>m����^?�e=�q�{�����i��.�T�O�?���? s�?�D����h��%=?��?�	?��>)��DQ޾(����v�2{x��f� >��>xUl��ǅ��W���zI��W�Ž��n��>��>��?Y~?�$�>���>�ھ�&��Ǿ����U��A�%!6�c�� �,0Ǿ��j�	�B�þ�J�p>985��3�>���>��b>��Z>&}�>X��=��>,�q>�
�>�;�>�σ>�FE>�&>�=j��KR?�����'�Z�辙���H3B?�qd?�1�>�i�$��������?���?Rs�?�<v>�~h��,+��n?X>�>6��Iq
?�S:=;��=�<�U��2���2����K��>E׽� :��M�fnf�tj
?�/?���g�̾�;׽�V��R��=�{?'� ?����BB��6O�H4S�cZ�%�Q�����wb�k�CVm� ۊ�ꏌ��醿�g!��Z=�@?��?O�侭Oܾ�#�l����a�[�8>.��>�s>s��>+lv>���K�J���e��~��p;�JQ/?�ac?���>�QK?:�>?#*b?�x_?AJ>�=�>򧇾S+4? 4�=WN�>?��#?�&:?�?aY�>��#?�S�>�Z��a������Ϊ?]4?�?�U?!g?N���Ƽ�m���<�2~�}��<��w=(��="�<�O���=�|a>�X?�����8�����Gk>;7?�}�>*��>!��u+��l?�<C�>��
?�C�>� �i|r��b�"W�>���?���|=��)>���=������ҺI_�=�����=A"���l;��<M��=���=t�s��1��"��:Fe�;Rx�<�u�>I�?O��>�C�>H>��� �߶�bn�=�Y>�S>�>1Cپ�}��U$��$�g�Zy>�w�?{�?˸f=|�=r��=�{��U�����y���^��<��?K#?vWT?Õ�?��=?�i#?��>�*��L���^��#����?(!,?Ћ�>����ʾD񨿿�3�O�?<[?�=a�Ⱥ�7;)�'�¾�Խկ>?[/�Q/~�]��^D�E��Q��[}�����?���?�A�3�6��w辸����\��
�C?q!�>�Z�>��>4�)���g�>%��1;>���>�R?�#�>y�O?�>{?Y�[?�nT>^�8��+��LΙ�Y�5���!>o@?���?"�?�y?bg�>��>4�)���V��A����ق��
W=f�Y>Z��>�&�>��>3��=X�ǽ�N��L�>�ٍ�=��b>3��>��>�>�nw>e��<@\?Q��>�VǾܼ��|�mҾ(��|j�?�o?�pI?�=���,<�޷��!��>�Љ?^,�?�W?��վ��=�s�����������>ؖ�>�	�>2%=c��1�>�W|>$Y�>��;ZN ��w��ߥ�N�#?X�f?zV>( ����c������W��V��*j��/����Jw���(�
��LK���ʢ���y�s���s��< ؾɼ׾]3 �>@?>�->�S�=ua�ˈ �$X�= �m=�{����|;�����;b����,��0�"��w��?^�<�-<����N{? @N?� -?�>?�s>��>s
���`q>�����8?\O>����h����M����������ھvS޾�{]�����s>�`��E�=�G/>���=4Ǟ;^��=��= �\=�R<��k=��=x��=�ܚ=��=���=��>čo?ۑ_�����b�_�<���]g3?���>3 >��ž8F!?o�칲S������@�ݾ�;�?���?�T�?���>�2~�Wy�>䕻�
k��H:=#�=#��>l'=�0��[�>�B	?R6���1��I+��E�?� @W^9?᪈�s�ѿ{�>+�C>1.>C R�h&0�X�S�˘n���]���&?�p9�����Mv�>���=��ھ/>����%=�0>��==����]�J�=�m�	�==�e]=8u�>KoC>��=�8ý�ܴ=�e=���=կW>,S���N�Yu��{"=6��=ng>ei/>'�>��?��/?$d?>c�>�o��MϾ�Q���z�>?��=�i�>n��=|�D>`��>�7?�:D?��K?4��>)ǃ=sm�>:�>� -���m���侥V����<�?�Ն?���>c�J<Q6B�����=�`½i�?`�1?+	?˝>���1�뿰�2���9�"���>���>��h���U�����Ո��AI�=��>i��>lyj>�W�>؟�>�C�>ު�=��>t�A>?�!>��=���'��&���Y\=���<�FU=�q���.����=���Cӎ��s=Oߔ<�tp�-GûT�=lK�>��>T��>w��=襾�?=>�����J�%�=o���C���f�&�~�+�'��+*�4&>ɩ?>�+���������>��Q>�n>c��?1p?�*>��"�[�Ѿ	ܚ�`�\��7;�u�=@�>�B�B�7�_�_��]J�ȸ�
��>��>�>��l>,�	?�&x=:⾖a5���>�����-9��9q��<��9��i��ٺƘD?F�����=�~?�I?��?9��>���?�ؾ'60>�D��I�=��#q��f���?�'?I��>��Q�D���۾����Դ�>���o�G�;��U�6�ҽ`Ͼ�a�>=඾��Ͼq�:��ʉ�Ɓ��A`N��
]� *�>�i=?���?W!���l�d:����H�H��>�T?��>F��>���>�N�;���ń�ņH>��?���?�y�?��=qP�=s*9���>%�>h�?�?{p?�ʨ����>��>��=8�<��>�4A>��?>,*�>���>�Ϸ>�{S����7��U ��^�����=��U=[��>¬�>��|>J�s>���I�=���> ��>.!�>{Do>���>e��>�������?If���$t>W5f?A�>���;��=��>ڦs�G⫾�q��Ҫ�=IT�=�U>2g���I�M���	�>XͿ@�?�mJ>��E��8?T%�e�i>��>97�e�>���>��>~.�>��>��8>~�>W�G>K˫>��Ӿ�>��� �>C�N<R� �оMdx>X���7(�������v.I�~����h�H%j��9��B�=����<8�?�]���6k�S�)�� �L'?S�>��5?i⌾�刽��>@��>BV�>���׉��捿����?���?��@>齟>�lY?��?C�6��Xc�9]�ޝw��y@���b��`�:v���ǃ�=��'���O?h�s?s�D?r�<�r�>�F|?��#�\8��U~>~�-�J�3�6ǀ=~t�>h���漖���쾨�оO���W�>�5�?y
�?}?\���
���'>c<?�0?��|?
�0?��P?�����'?�a�=��???�
F?�/?���>j@>���=�ܛ=[7=`�O�7���|ѽ1���ڃ�S@)=��=��<���Ǝ=�x��_m<wa=�\�<��x<t�^<�I=qr�=v<><��>C�Z?��>W��>��8?�Q1���7��0��D-?�1�=4�~�����h����辉�=g7d?D�?��a?�'M>�E�IL5���$>�[�>��,>A`>�ٱ>�]���2��F�=B�>F�&>P��=�5T��g}��F��ٔ��ge<��/>d�>���>.�����;����&�Ūr>ʽ�Yо���#�n_��E���о��=>�(`?%?� ��S/�<[�x�2�?ߨ@?���?�?���=da���a���"��6&�~4�>^&>$N�,/��F���y�8�Z{����=H�:�m����
^>$�	��۾�Am�M&I�à�ب4=�����8=a��57Ծ$�~��0�=�<>ql��x!�cC���Z����I?�{=	���Q�U��ջ�K�>z=�>�:�>� V�\�}�>'@�H�����=��>%6>7w�X�� G��W�*u�>ڤD?�G~?�P�?�����To���3�8���>����<��?���>�>2?>H>@�������+��]{��0��k?���>�1�
E$���������7�xJ�>#�6?1�>1m$?�v'?bs0?C�{?}Q?4?L@�>]{v����̘2?��t?��p=�E�$����B�wI�0�"?A,?8_�G�>��?�j5?��8?�)8?��?&�d>�2���Q�zR�>ƝJ>Hg��i�����>t�6?��>�+p?�?Wh>je8�Wҗ��o-�x.�=�E>jH4?%�B?�D??٨r>��>�'�����=���>��m?R��?&΀?��=�?>��>pxN>���>��?��?�G?,e?_E?���>��=�	���T����������<��W=���=��������=jw�=.��=��<{�<��s��x���.SۺZ`�>�s>���B�0>G�ľV���@>�ߢ��N���Ԋ�O�:�߷=ǈ�>��?���>b#��Ւ=�>9>�>����4(?��?n?�U%;��b�n�ھ�K�p�>	B?K��=��l�儔�T�u��h=E�m?��^?�wW�n#��P�b?��]?h��=��þ��b�ω�t�O?2�
?�G��>��~?t�q?q��>-�e�(:n����Cb�0�j��Ѷ=*r�>_X�S�d�q?�>b�7?�N�>��b>�%�=Fu۾�w��q��`?��?�?���?x+*>N�n�W4࿉���9���U?/{�>�R���?"?�<ռ�CоOg��(���4Ͼe���󘾼΀�ܪ��������/�A��p�=�v?��r?��o?�U^?D��r&^�N��v�\ h��0�L���!��?���E�Txn��~-��I�)���ϼ�B]�%H�k �?�?
���+7?e���muξ>�����'>��~�`�G�<`y=�v{��t�=�o�=�u��K�3��I�?��>��>��L?A�[�!&@��l0���2��3�rC
>�N�> H�>�F�>h�h��5��_�R�37žʈ�~&�g�>�$a?i�X?���?2=�=�f&�b^t�^�ݾ�$$���-w>AH>�c�>	t��9��m�A��ZD�%&j����gN~����2�>�d?=�=:[�>\<�?u�?�W�AФ�M����FZ�E�=�i?/�d?���>i�m>��н;�A�>��>�? m�>Ж�>�ϯ��(?�F�� ���:/?��>��:?�a�>�2��&_]���U����P�z�=Zր?)]�/-��L.�>��W?��=��=Xά>�� �#���+��}w�vM��,�>ydF>���=��ž����(l�����{)?t�?�ؑ��)��"�>p�!?q6�>_�>1ǃ?�ڝ>Wn���z�;�/?�_?��I?۹@?���>��/=2����Ƚ��$�6�.=�1�>�[>H�y=���=���
Z�3����Q=�9�=�~̼�Q��( <ט����N</��<�>4>|�ڿ�K�l�վ���ba�3�	�Ҝ��	0���q��n��8���
���H�v��d���/��WU��e�����y�m��0�?M_�?�ޏ��.��Z♿�*��i�����>{��d������������ྋ¬�z5#� Q��i���d�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >VC�<�,����뾭����οA�����^?���>��/��p��>ݥ�>�X>�Hq>����螾k1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@ҨA?�f(��H쾇\Y=u�>�	?|�@>u|-����(P��I��>�:�?G�?�U=|WW��)
���e?��4<��F�[�6�=R<�==��K>��>����@�A�ٽ��4>�j�>�*'����	x]�*��<ql]>oCԽMӓ�oS�?�@!��T��~��V~��ǳ>**?�>��ؽA?Vl�6Lпn�V�|Ed?�?@���?�2?
��6�2?�Ǿ��'?�4>?���=m'2���6���"<����;��ҾaJ�'��>g<�>$n�3!��6��g�iO�=VM�=�J��c�¿����3!@=��мC5��y�$�1�P��k�����H��G,��~/=P�=�Nk>�4x>s�!>/P4>tO?��v?q��>~�i>�eĽbʙ�g��%��(��=��`R�g�پ�@��Rܾ�����%��z(��J¾� =���=�6R�:����� ��b��F�v�.?�v$>��ʾ��M� �-<Rpʾ񿪾�ل��ॽ�-̾�1�#"n�P͟?j�A?������V�d��pU�����m�W?�O����Uꬾ���=]�����=�$�>\��=\�⾓ 3�5~S�N�B?%A?�L��ʗ_��|�>H��P|ɺ}�H?{�?��>�s�>o�4?�����s
:��>��u=7
?l�?�}P<�ʾՁ<[�(?��O?�۪�	�b�>�	 ���W��-��de>�z��%���Ga> ���z�Q�&�{�T~�<��<��W?A��>��)����#����/���4=v�y?A[?b�>l�j?�C?�<�<���KBS�X$����=&/Y?�g?��>��y��$ξL�����5?�?e?�O>S�m�it�d.����s?�Cm? �?���y�|�)���6?�v?�r^�\s������V�d<�>Y[�>��>��9��l�>�>?�
#�pG������PY4��?��@���?��;<7!���=�;?\�>ݪO�{>ƾ]z��-���ؕq=�"�>)����dv���GR,�@�8?���?0��>ޓ��>���V>�ם���?=�?�.վ5��=���wd��n��Kٔ<�BM>4婽Rd���9ܾF�-���Ӿ������0� �w8g>!�@@�۽��>h�׺������ɿ�Ԉ�L� �~Ma���-? �?��I�l*�!�����{���S�j�!���w�.Е>�]L>Kp�쇾K�����B���`�_��>&�w����L��;���-Ož�.�<��>��>�Q�>'��=]U���c�?�����'�� ���p?[��?:k�?V�?�~����� �l��y�e?2s�?zՙ?�	Q>�f�dh�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�h�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�Wa?�nP����-m?�e�OP�>=�(�&��n^��qü6}b�Y���S������?gl�?��?"���5�s�6?�ƭ>Q���FW�����+ʿ>|�>��=g�i�[7>8�辽q4���>��?���?y�?I+��c��m�=��t?)l�>�Ã?#>�"�>u}�=+���?`�4>�@W=�G���W�>&.H?e�>
��=��I���4��nG��R���	��m=�:�>��^?>WG?��J>�~ֽuu�9m"����k�ｘ�����f�_����P?>�,>��#>�^]��]¾��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�-	?7�,P��X`~����7����=��7?�0��z>���>��=9ov�ܻ���s���>�B�?�{�?f��>a�l?ڀo���B���1=�K�>e�k?t?8�n�B󾯯B>��?������K�� f?8�
@yu@J�^?����ҿƥ������o���#'>DtG>���>1��`�=�;��w�;��<QpV>�%�>W�_>a�p>��>Vg>,�=*��c%��?��;,��]�;����Κ��m�!�-����pޮ����$>�������Į��޽�0:)��=�MQ?3�H?>iq?�
?D��m4>�����<�M���<=]q>Ҕ#?��??o,?��=�֪�GLd������������u�>�K)>4�>���>�-�>"�}<17D>�.Z>TF�>��>)y={C=��{=�V>��>���>JT�>wC<>��>;ϴ��1��<�h�W
w��̽�?Y��� �J��1���9������mi�=Rb.?V|>���?п]����2H?S���a)�^�+���>��0?�cW?̝>�����T��:>���s�j��`>�+ �nl���)�s%Q>�l?�f>�u>D�3�
_8�}�P�d��Z||>c!6?�涾:$9�"�u�αH��kݾ�@M>�ʾ>H3C�:n�D��� ��li��J{={r:?�|?�E��wϰ�@�u� 1��yXR>�,\>w�=N�=�YM>��b���ƽH��A.=���=U�^>�?P2>�q=�9�>u2���Ss�̜>��>Bx7>�(J?!?�o�P��0�i�s�-��[>���>�ԡ>�9�=�U����=���>-g>F'���/�I��/v�?�n>�'~�eT�I���B=x���9�=o��=_2��BQ�v�x=�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?�q>�^�?�U[?��>�V�=p�J�f����Z��ʎ>��=n-?L��>ֵ��f����ᕿ`���4u����_9�>��%=?s�>&��G ߾&��='E%���z=#��>���>\��=u4�>�:/?*�>q�`>�a=�Hm��;~�<;����K?���?*���2n��N�<X��=&�^��&?�I4?6k[�|�Ͼ�ը>�\?j?�[?d�>=��O>��F迿5~��@��<��K>'4�>�H�>�$���FK>��Ծ�4D�gp�>�ϗ>u����?ھ�,���R��EB�>�e!?���>�Ү=2?C&?�+s>���>)r>��j��Y�J�<�>|��>k?Ē�?��?����4�8�3��9����<]�ȰS>\�v?vO?�1�>���mќ���<������Ͻ�_�?%�l?����R?'V�?ό>?Ql5?eN>�����;zi�4݆>�_ ?^�
�b�A��
&���~	?��?U�>VԒ���u�����J���?"Z]?�-'?�2�!v`�J�þQ��<j�[��0Q�7(� ��<5#>� >�pZ�$X�=�@>��=�r��2����<=���>L��=�R4���b��F,?�F�ڃ�.ɘ=Ϭr�l}D���>��L>m����^?�e=�q�{�����i��.�T�O�?���? s�?�D����h��%=?��?�	?��>)��DQ޾(����v�2{x��f� >��>xUl��ǅ��W���zI��W�Ž��n��>��>��?Y~?�$�>���>�ھ�&��Ǿ����U��A�%!6�c�� �,0Ǿ��j�	�B�þ�J�p>985��3�>���>��b>��Z>&}�>X��=��>,�q>�
�>�;�>�σ>�FE>�&>�=j��KR?�����'�Z�辙���H3B?�qd?�1�>�i�$��������?���?Rs�?�<v>�~h��,+��n?X>�>6��Iq
?�S:=;��=�<�U��2���2����K��>E׽� :��M�fnf�tj
?�/?���g�̾�;׽�V��R��=�{?'� ?����BB��6O�H4S�cZ�%�Q�����wb�k�CVm� ۊ�ꏌ��醿�g!��Z=�@?��?O�侭Oܾ�#�l����a�[�8>.��>�s>s��>+lv>���K�J���e��~��p;�JQ/?�ac?���>�QK?:�>?#*b?�x_?AJ>�=�>򧇾S+4? 4�=WN�>?��#?�&:?�?aY�>��#?�S�>�Z��a������Ϊ?]4?�?�U?!g?N���Ƽ�m���<�2~�}��<��w=(��="�<�O���=�|a>�X?�����8�����Gk>;7?�}�>*��>!��u+��l?�<C�>��
?�C�>� �i|r��b�"W�>���?���|=��)>���=������ҺI_�=�����=A"���l;��<M��=���=t�s��1��"��:Fe�;Rx�<�u�>I�?O��>�C�>H>��� �߶�bn�=�Y>�S>�>1Cپ�}��U$��$�g�Zy>�w�?{�?˸f=|�=r��=�{��U�����y���^��<��?K#?vWT?Õ�?��=?�i#?��>�*��L���^��#����?(!,?Ћ�>����ʾD񨿿�3�O�?<[?�=a�Ⱥ�7;)�'�¾�Խկ>?[/�Q/~�]��^D�E��Q��[}�����?���?�A�3�6��w辸����\��
�C?q!�>�Z�>��>4�)���g�>%��1;>���>�R?�#�>y�O?�>{?Y�[?�nT>^�8��+��LΙ�Y�5���!>o@?���?"�?�y?bg�>��>4�)���V��A����ق��
W=f�Y>Z��>�&�>��>3��=X�ǽ�N��L�>�ٍ�=��b>3��>��>�>�nw>e��<@\?Q��>�VǾܼ��|�mҾ(��|j�?�o?�pI?�=���,<�޷��!��>�Љ?^,�?�W?��վ��=�s�����������>ؖ�>�	�>2%=c��1�>�W|>$Y�>��;ZN ��w��ߥ�N�#?X�f?zV>( ����c������W��V��*j��/����Jw���(�
��LK���ʢ���y�s���s��< ؾɼ׾]3 �>@?>�->�S�=ua�ˈ �$X�= �m=�{����|;�����;b����,��0�"��w��?^�<�-<����N{? @N?� -?�>?�s>��>s
���`q>�����8?\O>����h����M����������ھvS޾�{]�����s>�`��E�=�G/>���=4Ǟ;^��=��= �\=�R<��k=��=x��=�ܚ=��=���=��>čo?ۑ_�����b�_�<���]g3?���>3 >��ž8F!?o�칲S������@�ݾ�;�?���?�T�?���>�2~�Wy�>䕻�
k��H:=#�=#��>l'=�0��[�>�B	?R6���1��I+��E�?� @W^9?᪈�s�ѿ{�>+�C>1.>C R�h&0�X�S�˘n���]���&?�p9�����Mv�>���=��ھ/>����%=�0>��==����]�J�=�m�	�==�e]=8u�>KoC>��=�8ý�ܴ=�e=���=կW>,S���N�Yu��{"=6��=ng>ei/>'�>��?��/?$d?>c�>�o��MϾ�Q���z�>?��=�i�>n��=|�D>`��>�7?�:D?��K?4��>)ǃ=sm�>:�>� -���m���侥V����<�?�Ն?���>c�J<Q6B�����=�`½i�?`�1?+	?˝>���1�뿰�2���9�"���>���>��h���U�����Ո��AI�=��>i��>lyj>�W�>؟�>�C�>ު�=��>t�A>?�!>��=���'��&���Y\=���<�FU=�q���.����=���Cӎ��s=Oߔ<�tp�-GûT�=lK�>��>T��>w��=襾�?=>�����J�%�=o���C���f�&�~�+�'��+*�4&>ɩ?>�+���������>��Q>�n>c��?1p?�*>��"�[�Ѿ	ܚ�`�\��7;�u�=@�>�B�B�7�_�_��]J�ȸ�
��>��>�>��l>,�	?�&x=:⾖a5���>�����-9��9q��<��9��i��ٺƘD?F�����=�~?�I?��?9��>���?�ؾ'60>�D��I�=��#q��f���?�'?I��>��Q�D���۾����Դ�>���o�G�;��U�6�ҽ`Ͼ�a�>=඾��Ͼq�:��ʉ�Ɓ��A`N��
]� *�>�i=?���?W!���l�d:����H�H��>�T?��>F��>���>�N�;���ń�ņH>��?���?�y�?��=qP�=s*9���>%�>h�?�?{p?�ʨ����>��>��=8�<��>�4A>��?>,*�>���>�Ϸ>�{S����7��U ��^�����=��U=[��>¬�>��|>J�s>���I�=���> ��>.!�>{Do>���>e��>�������?If���$t>W5f?A�>���;��=��>ڦs�G⫾�q��Ҫ�=IT�=�U>2g���I�M���	�>XͿ@�?�mJ>��E��8?T%�e�i>��>97�e�>���>��>~.�>��>��8>~�>W�G>K˫>��Ӿ�>��� �>C�N<R� �оMdx>X���7(�������v.I�~����h�H%j��9��B�=����<8�?�]���6k�S�)�� �L'?S�>��5?i⌾�刽��>@��>BV�>���׉��捿����?���?��@>齟>�lY?��?C�6��Xc�9]�ޝw��y@���b��`�:v���ǃ�=��'���O?h�s?s�D?r�<�r�>�F|?��#�\8��U~>~�-�J�3�6ǀ=~t�>h���漖���쾨�оO���W�>�5�?y
�?}?\���
���'>c<?�0?��|?
�0?��P?�����'?�a�=��???�
F?�/?���>j@>���=�ܛ=[7=`�O�7���|ѽ1���ڃ�S@)=��=��<���Ǝ=�x��_m<wa=�\�<��x<t�^<�I=qr�=v<><��>C�Z?��>W��>��8?�Q1���7��0��D-?�1�=4�~�����h����辉�=g7d?D�?��a?�'M>�E�IL5���$>�[�>��,>A`>�ٱ>�]���2��F�=B�>F�&>P��=�5T��g}��F��ٔ��ge<��/>d�>���>.�����;����&�Ūr>ʽ�Yо���#�n_��E���о��=>�(`?%?� ��S/�<[�x�2�?ߨ@?���?�?���=da���a���"��6&�~4�>^&>$N�,/��F���y�8�Z{����=H�:�m����
^>$�	��۾�Am�M&I�à�ب4=�����8=a��57Ծ$�~��0�=�<>ql��x!�cC���Z����I?�{=	���Q�U��ջ�K�>z=�>�:�>� V�\�}�>'@�H�����=��>%6>7w�X�� G��W�*u�>ڤD?�G~?�P�?�����To���3�8���>����<��?���>�>2?>H>@�������+��]{��0��k?���>�1�
E$���������7�xJ�>#�6?1�>1m$?�v'?bs0?C�{?}Q?4?L@�>]{v����̘2?��t?��p=�E�$����B�wI�0�"?A,?8_�G�>��?�j5?��8?�)8?��?&�d>�2���Q�zR�>ƝJ>Hg��i�����>t�6?��>�+p?�?Wh>je8�Wҗ��o-�x.�=�E>jH4?%�B?�D??٨r>��>�'�����=���>��m?R��?&΀?��=�?>��>pxN>���>��?��?�G?,e?_E?���>��=�	���T����������<��W=���=��������=jw�=.��=��<{�<��s��x���.SۺZ`�>�s>���B�0>G�ľV���@>�ߢ��N���Ԋ�O�:�߷=ǈ�>��?���>b#��Ւ=�>9>�>����4(?��?n?�U%;��b�n�ھ�K�p�>	B?K��=��l�儔�T�u��h=E�m?��^?�wW�n#��P�b?��]?h��=��þ��b�ω�t�O?2�
?�G��>��~?t�q?q��>-�e�(:n����Cb�0�j��Ѷ=*r�>_X�S�d�q?�>b�7?�N�>��b>�%�=Fu۾�w��q��`?��?�?���?x+*>N�n�W4࿉���9���U?/{�>�R���?"?�<ռ�CоOg��(���4Ͼe���󘾼΀�ܪ��������/�A��p�=�v?��r?��o?�U^?D��r&^�N��v�\ h��0�L���!��?���E�Txn��~-��I�)���ϼ�B]�%H�k �?�?
���+7?e���muξ>�����'>��~�`�G�<`y=�v{��t�=�o�=�u��K�3��I�?��>��>��L?A�[�!&@��l0���2��3�rC
>�N�> H�>�F�>h�h��5��_�R�37žʈ�~&�g�>�$a?i�X?���?2=�=�f&�b^t�^�ݾ�$$���-w>AH>�c�>	t��9��m�A��ZD�%&j����gN~����2�>�d?=�=:[�>\<�?u�?�W�AФ�M����FZ�E�=�i?/�d?���>i�m>��н;�A�>��>�? m�>Ж�>�ϯ��(?�F�� ���:/?��>��:?�a�>�2��&_]���U����P�z�=Zր?)]�/-��L.�>��W?��=��=Xά>�� �#���+��}w�vM��,�>ydF>���=��ž����(l�����{)?t�?�ؑ��)��"�>p�!?q6�>_�>1ǃ?�ڝ>Wn���z�;�/?�_?��I?۹@?���>��/=2����Ƚ��$�6�.=�1�>�[>H�y=���=���
Z�3����Q=�9�=�~̼�Q��( <ט����N</��<�>4>|�ڿ�K�l�վ���ba�3�	�Ҝ��	0���q��n��8���
���H�v��d���/��WU��e�����y�m��0�?M_�?�ޏ��.��Z♿�*��i�����>{��d������������ྋ¬�z5#� Q��i���d�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >VC�<�,����뾭����οA�����^?���>��/��p��>ݥ�>�X>�Hq>����螾k1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@ҨA?�f(��H쾇\Y=u�>�	?|�@>u|-����(P��I��>�:�?G�?�U=|WW��)
���e?��4<��F�[�6�=R<�==��K>��>����@�A�ٽ��4>�j�>�*'����	x]�*��<ql]>oCԽMӓ�oS�?�@!��T��~��V~��ǳ>**?�>��ؽA?Vl�6Lпn�V�|Ed?�?@���?�2?
��6�2?�Ǿ��'?�4>?���=m'2���6���"<����;��ҾaJ�'��>g<�>$n�3!��6��g�iO�=VM�=�J��c�¿����3!@=��мC5��y�$�1�P��k�����H��G,��~/=P�=�Nk>�4x>s�!>/P4>tO?��v?q��>~�i>�eĽbʙ�g��%��(��=��`R�g�پ�@��Rܾ�����%��z(��J¾� =���=�6R�:����� ��b��F�v�.?�v$>��ʾ��M� �-<Rpʾ񿪾�ل��ॽ�-̾�1�#"n�P͟?j�A?������V�d��pU�����m�W?�O����Uꬾ���=]�����=�$�>\��=\�⾓ 3�5~S�N�B?%A?�L��ʗ_��|�>H��P|ɺ}�H?{�?��>�s�>o�4?�����s
:��>��u=7
?l�?�}P<�ʾՁ<[�(?��O?�۪�	�b�>�	 ���W��-��de>�z��%���Ga> ���z�Q�&�{�T~�<��<��W?A��>��)����#����/���4=v�y?A[?b�>l�j?�C?�<�<���KBS�X$����=&/Y?�g?��>��y��$ξL�����5?�?e?�O>S�m�it�d.����s?�Cm? �?���y�|�)���6?�v?�r^�\s������V�d<�>Y[�>��>��9��l�>�>?�
#�pG������PY4��?��@���?��;<7!���=�;?\�>ݪO�{>ƾ]z��-���ؕq=�"�>)����dv���GR,�@�8?���?0��>ޓ��>���V>�ם���?=�?�.վ5��=���wd��n��Kٔ<�BM>4婽Rd���9ܾF�-���Ӿ������0� �w8g>!�@@�۽��>h�׺������ɿ�Ԉ�L� �~Ma���-? �?��I�l*�!�����{���S�j�!���w�.Е>�]L>Kp�쇾K�����B���`�_��>&�w����L��;���-Ož�.�<��>��>�Q�>'��=]U���c�?�����'�� ���p?[��?:k�?V�?�~����� �l��y�e?2s�?zՙ?�	Q>�f�dh�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�h�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�Wa?�nP����-m?�e�OP�>=�(�&��n^��qü6}b�Y���S������?gl�?��?"���5�s�6?�ƭ>Q���FW�����+ʿ>|�>��=g�i�[7>8�辽q4���>��?���?y�?I+��c��m�=��t?)l�>�Ã?#>�"�>u}�=+���?`�4>�@W=�G���W�>&.H?e�>
��=��I���4��nG��R���	��m=�:�>��^?>WG?��J>�~ֽuu�9m"����k�ｘ�����f�_����P?>�,>��#>�^]��]¾��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�-	?7�,P��X`~����7����=��7?�0��z>���>��=9ov�ܻ���s���>�B�?�{�?f��>a�l?ڀo���B���1=�K�>e�k?t?8�n�B󾯯B>��?������K�� f?8�
@yu@J�^?����ҿƥ������o���#'>DtG>���>1��`�=�;��w�;��<QpV>�%�>W�_>a�p>��>Vg>,�=*��c%��?��;,��]�;����Κ��m�!�-����pޮ����$>�������Į��޽�0:)��=�MQ?3�H?>iq?�
?D��m4>�����<�M���<=]q>Ҕ#?��??o,?��=�֪�GLd������������u�>�K)>4�>���>�-�>"�}<17D>�.Z>TF�>��>)y={C=��{=�V>��>���>JT�>wC<>��>;ϴ��1��<�h�W
w��̽�?Y��� �J��1���9������mi�=Rb.?V|>���?п]����2H?S���a)�^�+���>��0?�cW?̝>�����T��:>���s�j��`>�+ �nl���)�s%Q>�l?�f>�u>D�3�
_8�}�P�d��Z||>c!6?�涾:$9�"�u�αH��kݾ�@M>�ʾ>H3C�:n�D��� ��li��J{={r:?�|?�E��wϰ�@�u� 1��yXR>�,\>w�=N�=�YM>��b���ƽH��A.=���=U�^>�?P2>�q=�9�>u2���Ss�̜>��>Bx7>�(J?!?�o�P��0�i�s�-��[>���>�ԡ>�9�=�U����=���>-g>F'���/�I��/v�?�n>�'~�eT�I���B=x���9�=o��=_2��BQ�v�x=�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?�q>�^�?�U[?��>�V�=p�J�f����Z��ʎ>��=n-?L��>ֵ��f����ᕿ`���4u����_9�>��%=?s�>&��G ߾&��='E%���z=#��>���>\��=u4�>�:/?*�>q�`>�a=�Hm��;~�<;����K?���?*���2n��N�<X��=&�^��&?�I4?6k[�|�Ͼ�ը>�\?j?�[?d�>=��O>��F迿5~��@��<��K>'4�>�H�>�$���FK>��Ծ�4D�gp�>�ϗ>u����?ھ�,���R��EB�>�e!?���>�Ү=2?C&?�+s>���>)r>��j��Y�J�<�>|��>k?Ē�?��?����4�8�3��9����<]�ȰS>\�v?vO?�1�>���mќ���<������Ͻ�_�?%�l?����R?'V�?ό>?Ql5?eN>�����;zi�4݆>�_ ?^�
�b�A��
&���~	?��?U�>VԒ���u�����J���?"Z]?�-'?�2�!v`�J�þQ��<j�[��0Q�7(� ��<5#>� >�pZ�$X�=�@>��=�r��2����<=���>L��=�R4���b��F,?�F�ڃ�.ɘ=Ϭr�l}D���>��L>m����^?�e=�q�{�����i��.�T�O�?���? s�?�D����h��%=?��?�	?��>)��DQ޾(����v�2{x��f� >��>xUl��ǅ��W���zI��W�Ž��n��>��>��?Y~?�$�>���>�ھ�&��Ǿ����U��A�%!6�c�� �,0Ǿ��j�	�B�þ�J�p>985��3�>���>��b>��Z>&}�>X��=��>,�q>�
�>�;�>�σ>�FE>�&>�=j��KR?�����'�Z�辙���H3B?�qd?�1�>�i�$��������?���?Rs�?�<v>�~h��,+��n?X>�>6��Iq
?�S:=;��=�<�U��2���2����K��>E׽� :��M�fnf�tj
?�/?���g�̾�;׽�V��R��=�{?'� ?����BB��6O�H4S�cZ�%�Q�����wb�k�CVm� ۊ�ꏌ��醿�g!��Z=�@?��?O�侭Oܾ�#�l����a�[�8>.��>�s>s��>+lv>���K�J���e��~��p;�JQ/?�ac?���>�QK?:�>?#*b?�x_?AJ>�=�>򧇾S+4? 4�=WN�>?��#?�&:?�?aY�>��#?�S�>�Z��a������Ϊ?]4?�?�U?!g?N���Ƽ�m���<�2~�}��<��w=(��="�<�O���=�|a>�X?�����8�����Gk>;7?�}�>*��>!��u+��l?�<C�>��
?�C�>� �i|r��b�"W�>���?���|=��)>���=������ҺI_�=�����=A"���l;��<M��=���=t�s��1��"��:Fe�;Rx�<�u�>I�?O��>�C�>H>��� �߶�bn�=�Y>�S>�>1Cپ�}��U$��$�g�Zy>�w�?{�?˸f=|�=r��=�{��U�����y���^��<��?K#?vWT?Õ�?��=?�i#?��>�*��L���^��#����?(!,?Ћ�>����ʾD񨿿�3�O�?<[?�=a�Ⱥ�7;)�'�¾�Խկ>?[/�Q/~�]��^D�E��Q��[}�����?���?�A�3�6��w辸����\��
�C?q!�>�Z�>��>4�)���g�>%��1;>���>�R?�#�>y�O?�>{?Y�[?�nT>^�8��+��LΙ�Y�5���!>o@?���?"�?�y?bg�>��>4�)���V��A����ق��
W=f�Y>Z��>�&�>��>3��=X�ǽ�N��L�>�ٍ�=��b>3��>��>�>�nw>e��<@\?Q��>�VǾܼ��|�mҾ(��|j�?�o?�pI?�=���,<�޷��!��>�Љ?^,�?�W?��վ��=�s�����������>ؖ�>�	�>2%=c��1�>�W|>$Y�>��;ZN ��w��ߥ�N�#?X�f?zV>( ����c������W��V��*j��/����Jw���(�
��LK���ʢ���y�s���s��< ؾɼ׾]3 �>@?>�->�S�=ua�ˈ �$X�= �m=�{����|;�����;b����,��0�"��w��?^�<�-<����N{? @N?� -?�>?�s>��>s
���`q>�����8?\O>����h����M����������ھvS޾�{]�����s>�`��E�=�G/>���=4Ǟ;^��=��= �\=�R<��k=��=x��=�ܚ=��=���=��>čo?ۑ_�����b�_�<���]g3?���>3 >��ž8F!?o�칲S������@�ݾ�;�?���?�T�?���>�2~�Wy�>䕻�
k��H:=#�=#��>l'=�0��[�>�B	?R6���1��I+��E�?� @W^9?᪈�s�ѿ{�>+�C>1.>C R�h&0�X�S�˘n���]���&?�p9�����Mv�>���=��ھ/>����%=�0>��==����]�J�=�m�	�==�e]=8u�>KoC>��=�8ý�ܴ=�e=���=կW>,S���N�Yu��{"=6��=ng>ei/>'�>��?��/?$d?>c�>�o��MϾ�Q���z�>?��=�i�>n��=|�D>`��>�7?�:D?��K?4��>)ǃ=sm�>:�>� -���m���侥V����<�?�Ն?���>c�J<Q6B�����=�`½i�?`�1?+	?˝>���1�뿰�2���9�"���>���>��h���U�����Ո��AI�=��>i��>lyj>�W�>؟�>�C�>ު�=��>t�A>?�!>��=���'��&���Y\=���<�FU=�q���.����=���Cӎ��s=Oߔ<�tp�-GûT�=lK�>��>T��>w��=襾�?=>�����J�%�=o���C���f�&�~�+�'��+*�4&>ɩ?>�+���������>��Q>�n>c��?1p?�*>��"�[�Ѿ	ܚ�`�\��7;�u�=@�>�B�B�7�_�_��]J�ȸ�
��>��>�>��l>,�	?�&x=:⾖a5���>�����-9��9q��<��9��i��ٺƘD?F�����=�~?�I?��?9��>���?�ؾ'60>�D��I�=��#q��f���?�'?I��>��Q�D���۾����Դ�>���o�G�;��U�6�ҽ`Ͼ�a�>=඾��Ͼq�:��ʉ�Ɓ��A`N��
]� *�>�i=?���?W!���l�d:����H�H��>�T?��>F��>���>�N�;���ń�ņH>��?���?�y�?��=qP�=s*9���>%�>h�?�?{p?�ʨ����>��>��=8�<��>�4A>��?>,*�>���>�Ϸ>�{S����7��U ��^�����=��U=[��>¬�>��|>J�s>���I�=���> ��>.!�>{Do>���>e��>�������?If���$t>W5f?A�>���;��=��>ڦs�G⫾�q��Ҫ�=IT�=�U>2g���I�M���	�>XͿ@�?�mJ>��E��8?T%�e�i>��>97�e�>���>��>~.�>��>��8>~�>W�G>K˫>��Ӿ�>��� �>C�N<R� �оMdx>X���7(�������v.I�~����h�H%j��9��B�=����<8�?�]���6k�S�)�� �L'?S�>��5?i⌾�刽��>@��>BV�>���׉��捿����?���?��@>齟>�lY?��?C�6��Xc�9]�ޝw��y@���b��`�:v���ǃ�=��'���O?h�s?s�D?r�<�r�>�F|?��#�\8��U~>~�-�J�3�6ǀ=~t�>h���漖���쾨�оO���W�>�5�?y
�?}?\���
���'>c<?�0?��|?
�0?��P?�����'?�a�=��???�
F?�/?���>j@>���=�ܛ=[7=`�O�7���|ѽ1���ڃ�S@)=��=��<���Ǝ=�x��_m<wa=�\�<��x<t�^<�I=qr�=v<><��>C�Z?��>W��>��8?�Q1���7��0��D-?�1�=4�~�����h����辉�=g7d?D�?��a?�'M>�E�IL5���$>�[�>��,>A`>�ٱ>�]���2��F�=B�>F�&>P��=�5T��g}��F��ٔ��ge<��/>d�>���>.�����;����&�Ūr>ʽ�Yо���#�n_��E���о��=>�(`?%?� ��S/�<[�x�2�?ߨ@?���?�?���=da���a���"��6&�~4�>^&>$N�,/��F���y�8�Z{����=H�:��ڠ��[b>w��[޾5�n���I���{M=���4V=8�s־����=t&
>���� ����Ϊ��,J?t�j=�l���AU�_�����>���>�ޮ>��:�-Hv�І@�󮬾\�=��>_�:>��?��ˁG�v/����>�E?�@0?4��?$��P^�9�	����)A��4�=p!?�W�>��"?�A�>�%=�ԡ�w!�&�������>'b�>�~ �9F�%���~R����^��>��>ý�>�4?h25?��?�{Z?'W?�]�>�N�>��t�y�Ͼ��3?^��?.��y��~%v�%�c�x��d!0?�:?<;���> ��>�� ?~I?��@?}X? �=�����+�n[�>s�w>[5`������ՠ>]w=?�r�>��~?q�p?l�D>i�"��8ľ��}�R�=��@>�X?L�E?(tP?�S>Ky�>d������<���>q�U?녁?�@k?(l�<���>ҟ5>���>>�1�>L+�>?��T?�g?�XE?��>7a�<{+���?ܼ2-r�vټi�<��#��C=��ǽ0�0�s���Qs=���<<Ð��8�c����ǼA��8l�=hu�>'�s>h��^1>-�ľ�!��zA>�����[��
⊾�;:�r�=���>��?정>^;#�=���>��>����((?��?p?�f;̕b��۾��K����>�B?�l�=�l�Ur��X�u���h=��m?�{^?�tW����h�b?��]?�g�@=���þ�b�e��V�O?��
?�G��>#�~?��q?W��>X�e�9n�����Db�A�j�ն=�p�>�X���d�q=�>{�7?xN�>��b>#+�=1s۾��w�@s��c?]�?��?=��?�.*>��n�>3�+�
�aǔ���b?���>_:��I� ?�� ��1ž�I������v��$ѷ�c����l���ࣾG@��j��2۽��=c?�v?�jm?	AX?^����\��#V�`r�a�J�e��;�C�@�&L�h�D���l�#�`~��b���#<�`�V@���?�6/?߱I��v?��������u���O*>?�7�r���g�=~��<�-�=@8@=/If��%e�x����� ?��>3�>x�W?z�d��I<�fC6�����˟���J>��>��W>��>��6=���h�6�1������ �Z1v>�o?T�2?��b?A�$>��+���u��}���<�\���a>�b>0{�>;kýg�{�e�G�S�V��	z��S���@��G&�n`�=�)?.�%>w?N�?3F�>:K8�nT���w���L��)��A?�k�?g�?G>U���ƾH��>��m?���>�=�>�.��Κ"�E |�@�Ž4��>Z*�>c6�>�ds>�c#��]��֐�ꎿb!;���=��i?&��Z\�1V�>ڛL?_�'<��<h\�>&Ꮍ*�}�:�3�2��=s�?�X�=�9>�CǾG���{�M����)?@K?�$���(��K�>�j!?���>�:�>7�?��>�u��2�W<�O?�_?2J?@L@?��>f�$=2����ȽB�%�x==�z�>4}\>#/~=͚�=���T�Z��
'��9=��=2���T��F�<����F�S<��< �=>��ۿ��N��̾����G�>���A��˩�
����	$�D_��L&��ޓ|�a���;=�,Da��Qg��J��ȝp����?��?$䍾�����(���#~��������>��j�)U�������
��u�����찾�g&��P�Oj�b3f�P�'?�����ǿ񰡿�:ܾ3! ?�A ?:�y?��5�"���8�� >SC�<�,����뾭����ο@�����^?���>��/��o��>ߥ�>�X>�Hq>����螾y1�<��?8�-?��>Ȏr�0�ɿc���w¤<���?0�@�&D?g�����o��=�V�>�?;�E>�<L�[���iľ�q�>�^�?��?48~=J�R��1��fZ?���;E�п�:"��=� �=%h@=�D�^�%>(�v>ڔ-��G������V>[c�>�x��{���R��'<ʕT>�?��N���Є?�f\�V+f�P�/�]��(p>��T?�!�>1��=��,?�SH�xkϿ��\� �`?p,�?���?1)?\c�����>P�ܾ��M?�U6?��>�]&��t�z��=V��~���㾘V���=$r�>��>��+�9����O�`ۚ��>�=.j�L�ӿ~8ξ���u�Y<�ж=��d����S�
���맠���H�*s�="�=ז'>yJD>f�9>�܏>�X?��v?:[�>R�>0�)��9b��8��s�]��﷾F�׾L�h��R�����0�@M*���/����$��!=���=�6R�f���?� �Y�b�=�F���.?�v$>P�ʾ��M��-<{pʾU����ۄ��ॽ�-̾
�1�#"n�f͟?��A?������V�W��X�r���\�W?P�ϻ�|ꬾ��=����y�=�$�>���=q��� 3�s~S��m2?BU ?��ľ9T��P�3>����w=�G1?ƞ�>ɫ =#U�>��"?w'�U䩽!�]>E�'>�m�>_a�>zS>�����ֽE� ?�hO?�콕��jŌ>�8ž�.[��i/=D >bv�q���K>���<ǭ��t׼�O���
=kVW?i�>Vn*�M;�Î���6�X�S=�Bz?�!?#�>]sk?��A?&��<s%��S�^�9}=kpW?��h?�>��~�+;s�����5?u�e?�fN>�l�͗�-l.�!��~P?u�m?�?�ڗ���|��Ӓ�6��;a6?��h?5D�]���f"?�Œ �}ʥ>�?~�>l��;�?�Ӫ>{H�q����Gǿ�~��&�?�w@�#�?<�o�zǸ����=|��>��?�x����}�.��	ؾ��=�=�>�iľGO�r�9�-'s��@i?��K?���>�bA�]&�_��=���%��?DΑ?�4־^��=,� ���9��~�<^�;�/�>�_��㜽����C
E��8ž�R�lM���vI�}˃> �@��V��?�X����q��E��������n��_�?�&�>@/ �"j�����Sx�b�^���;��t>�/Nv>�K�=����ܾt��'�B�b��;��>Q��=�vc>�E��7��"��t䄽���>p?zE�>�>�8{��r�?Y��=��/z����B�jUI?���?�0�?��R?���>3�k��Q9>p�z>�%?˲??Jg??��=#����r�<%�j?�_��xU`��4�qHE��U>�"3?�B�>R�-���|=�>���>g>�#/�w�Ŀ�ٶ�:���Y��?��?�o���>r��?rs+?�i�8���[����*��+��<A?�2>���G�!�C0=�RҒ���
?R~0?{�c.�W�_?'�a�I�p���-���ƽ�ۡ>��0�f\�O�����Xe�
���@y����?K^�?i�?µ�� #�f6%?�>l����8Ǿm�<���>�(�>�)N>�G_���u>����:�	i	>���?�~�?Mj?���� ����U>	�}?��>4�?;��=pA�>�`>枝� ;[t>7�=Hޣ�_�?�M??$�>���=tL8�&,�'CE�$�Q�P��t�<��f�>�A^?��J?��F>t3��H�������H���K�(�-��B��ϴԽ�58>9�5>TX>�xV�����?3p�{�ؿ�j��Wv'�,54?���>��?����t�
�>;_?y�>h7��+���$��>=����?/G�?I�?w�׾9t̼�>)�>K�>[ ս���.�����7>��B?M�JD��K�o�)�>g��?ȶ@�ծ?*i��=	?��T���8ꀿ���?�4��>E�8?St�3�>��>�=r�u�����s��ɺ>���?w�?��>l?^n��:D��J==��>�k?��	?�7e�`1��&�D>&J
?=�����(�XKc?(
@�@�]?5E��lɿEϝ�G�v��ؾ��=_�*>��C>��S���=1񄽂r�<v�<��g>n�>W|�>��l>�$j>�>5>)y�>a��J(�*S������6�4��^ھ\�a$�E�־'���_�g�Ѿ՟�4X����n�wD̼�T��)�ֽ�K���:Z>�dK?��7?k	c?)�?�+�u��=����	��~*���@>�>�>��A?}�O?��'?���<�����[�aE}�ǚ�J+���H�>0>���>J�>r�>j\�=ɱh>��H>4�4>�4-=�=�[�=<�>J��>�]�>z��>*Z�>�C<>��>Fϴ��1��i�h��
w�Z̽3�?����N�J��1���9��Ҧ��i�=Gb.?|>���?пe����2H?$���z)���+���>}�0?�cW?'�>��h�T�/:>7����j�.`>�+ ��l���)��%Q>vl?p�f>�$u>��3�?`8���P��}���}|>66?�궾�&9��u�k�H��_ݾrRM>�¾>" D��g�������hui���{=�v:?Ѐ?�,��Nݰ�z�u��B���QR>O?\>K=�=)MM>qc���ƽfH�a}.=���=:�^>I�	?S&_>>�Z<���>*���:���]��>�e�>o">8xM?�{&?i�K�����W>�����]>�$�>�	�>$,>��`�D�=�W?�hK>쬀��������O�p�/��>GĽ=Q�ͬ=|s=��߽+W>�҆=&z���}t�=�~?���(䈿��e���lD?S+?] �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>}x��Z�������u�d�#=[��>�8H?�V��l�O�y>��v
?�?�^�ީ����ȿ-|v����>V�?���?g�m��A���@����>;��?�gY?moi>�g۾,`Z����>ֻ@?�R?�>�9�{�'���?�޶?ԯ�?�J>2��?-�*?d�>#5�>�[��8��*4V�7k?8�E=�p�>�*�>a"�<�{R�����!㞿S������
G�>}�/=��>�}�7�¾,ɜ>i���ŀǾ�6_�\B�>��B>��B��i�>m�?�:�>Z,b>��I��은��Ν��IL?��?�M�Km��u�<�h�=�Z��U?�l3?b�'��F;�-�>�N\?e�?_�Z?Ȗ�>8�Ӛ�5~��")����<�K>+��>
��>j���g�M>2rӾB�bP�>J��>U���#�۾C���N}�{��>�W!?nX�>�r�=2�?�N(?Ɓ[>!��>&�6�EC��x�G�oh�>�h�>�P?�3�?X�?�¹���8�TQ��-Q���_�u�.>�\u?�?�ŭ>����<��c��=O��֠}��kv?�r?�ý�9�>���?�_B?�! ?A�D>��(��Ѿjvv��Z�>p;!?�s��*A���%�%����?�?Q�>�R��.wѽ7�ӼW,�����>�?b�[?�&?T+�/i`��þ��<B)�L���;��f�4�>!P>�c����=�\>��=Vm�Ƒ5����<G̿=��>rz�=�5��;����"?�z�<8վ�Gݽ�E�����[r>iE>ڂ�<�o?bپ��W��Ƕ�|}��\��=\h�?�[�?ӛ?����a�d���0?4[�?B?�?�x��M������E���������o��=��>� �=t)�-ݜ�=���8��]����N*�l��>$�>��?GE�>e�>GG�>�";CL0�&�˾��5O���
���?���u���"���<��w�P"ǾB>���}>ݷ�a��>��?��{>��f>�̍>G��=SЃ>�O>ǥ�>R��>x�b>��>P� >v9a=q�d��kR?v1���'�П�,e��5/B?8$d?p�>��k�6����0���?+}�?�N�?v>#h��+�P?�R�>Z��)<
?�U<=����l�<nv�����o��G�6�>��ӽڸ9���L�̦e��d
?��?Ix��j�̾`hٽ���z�<4B�?��)?9&��E��|k�H�8�#�D��4�����G���2&��_�)쎿=��C샿�k!�0�>f�?+�?+���y
վ�b���|�ؼ=��=(��>Ϯ�>�>��A>5�
�+�J��cD���c���?8�?�*�>?R??K�+?cEJ?�aJ?
i�>�8�>�쳾q��>�y����>s�	?�!??�w:?[;?��?C�?E	L>�!�����z۾V�?��?f�?<� ?��?��n�蜝�۬��H�ռn��4��2��=�,�=��üo��-�s<�K�>a"?z�ݽ	�/�8�Ѿ�>/	C?���>���>�=����¾;�`=Wi�>l?l=�>N���K�_�>K�[��>�o?zY�p��=�2>n>����;ł=��W���=�^��8�8�<�~�=ҹ;�F�W��O3�����E�RS���t�>�?���>yC�>�@��� �0���e�=$Y>HS>%>�Eپ�}���$��J�g�`^y>�w�?�z�?��f=��=ӕ�=�|��QU������������<�?	J#?�WT?R��?t�=?gj#?�>+�jM���^�����î?s",?���> ����ʾg憎�3�f�?�`?J:a�����7)���¾�սj�>�Y/�.~�a���D��o������y��u��?｝?��@�a�6��u�ǿ��WT��ǑC?��>�`�>A�>'�)���g��$��);>��>�R?7;�>%�H?٢a?��Q?+�c>T�,�jk���×��&��� >I�L?�.�?�Ȓ?�u?|N�>"��=�n<���޾���^E�lp�&iv��<�W7>ڱ�>�\�>u'�>2 >~��2	��QcB��x�=`�>���>�ѭ>�ݽ>3�>X��=�~I?y��>����2��v�X��u�>��?�T�?Q_Q?�s)�����5��຾��>ə�?gU�?��2?͟���>83���ﾝݏ���>�1�> B�>��#���C=��^>t��>�9?��;�8�<���1�F(��3�?��g?��=��Ŀ�&y�S�p���������xe�`5T���n����7�:-��m;^�\����yf�������ԾD�ξQ��0<���?z�3>#�>4�=	w���_x���*N6�֒�=�m�=�S��3<�-��)���#���9���T5����<B��=��Ǿ�|?bH?�~,?��E?�ɀ>�f>�I�	��>�Ȁ�Ɇ?�J>��:��޴��s5�D?���3%ྡ7Ѿ)6_�6ӟ�l�>�'�<� >{�0>���=2B�<
��=��=�zg=Vw�z�C=)��=^o�=�>�=���=т�=��>NGv?�����(	R�����x9?:C�>^��=�����PB?g">S܂�kb��(�����?0��?�k�?��?7�r�/<�>e����YP�'�=���6z.>V�=H�2���>]�D>��n����7Ƚ�?.@~q;?zM��klͿ�#>��/>#�>��Q���0��^W�AKQ��qD��?K�:��F���9�>rK�=�۾��Ǿ��S=��F>]��=���E_�Dq�=�+~���T=��+=��>Y�A>�y�=`���G��=p�Y=JP�=KqR>9�(�������Ȇ= ��=Du>R�H>7�>q�?m0?zd?���>9Nm�yξ�v���ҋ>���=���>콅=�nB>�9�>��7?*�D?��K?+�>�K�=�Ӻ>�ަ>�e,�S�m�{��֧��p�<&��?o��?�ܸ>$�[<PMA�����=�#(ý��?��1?�? ��>���]��8���0��a����v=�')=�'��_{<{@H=�����W���0>.��>�$�>��>}��>�;:>NLk>^��>�=Ǉ=�� >�Í���<]T��\P8=2�ٽw�=���
렽:�<�:�5Q��1�<�ݫ�j0x�0��=l-�=
��>'�=�x�>ű�<30���h>m�ξ
U;����=�f���=5�(oZ�m������s{���6>J-M>N]��T�����>3Q>�C�>��?[>y?SW|>�g���!�z����K
�h�2����>eK�=�,���
5�B�w�t�R��M���>�ߎ>��>��l>,��"?�,�w=V�!b5��>|�����T)�Q9q��?������_i��Һ��D?gF��ٛ�="~?��I??�?���>O���ؾ�90>mH��H�=i�L)q��h����?!'?e��>a�D�D����d
���>vV��J�r2��V�?�Y�T����Z�>�����}�-BA�HҀ�}����L�S���>�[?J��?g2#��De��8�;��S�����>v�L?<�>{�>�?m`��x	��m���X�=�w�?���?��?���=��7=���Y٬>H��>��?kK�?[ot?��]@�>���=ν�=��y�kB�=F�Z=<~�=!�Q>yp?b�?��>�O��A� � V˾8��{���<?�=R��>�5�>g��>�q>�Й=Ɵ>=�Y�>�{�>�C�>�Ƹ>
��>m��>����jR?���=aaD>iUE?Ѷ�>"�:=�Ƕ��/û�&@��������Ю��;�?>M��=�`�=�+�=e��>��Ŀ`?�?���>Eb��3,?�&���g>z�
>��N=��=1�>R%O>iy�>�|�>�Q=>up��/�<�9>]NӾ'l>j���c!�,C�3R��Ѿm~z>����� &�w��ߋ��`KI��n��hh�}j��-��<=��ٽ<�F�?�����k�@�)�R����?�O�>6?dь�m눽��>���>n��>�K��7���Ǎ��e�1�?_��?���<�?>�K�?�C�>��M�k�c��6u�Mp��y<��y���)h�b���7H��!���졽URO?�M_?O3Q?y��=;��>[�f?̪��r~��?>U��/����`=�_�>x��0��ʣ�I����2�q�a>7z�?S��?�8&?Y戾�H3>��>[�>8?Of?8�6?�-C?��#�:��>�IE�Ϥ?-$?}3?d�Z?j
 ?V�H>_:�<^g�~�=��7�crt��f��s���t~z����=ѱ`��R)�NF��mo��=��1=)	F=�꼆W;���=�O�=7�d�C���9ʐ>�S?�`�>h2Z>,?��ν��&��u���?�X�=U ��ˀ��ԡ�(L���#>C�t?��?�{]?2�_>Q�<���U��[H>�ɘ>��>�A]>xx�>l�o����S��9�>t�>^=�=�q�~����W�S��|���8e>��>�U|>򀎽Rf'>4�����y�ve>��R�����;S���G��1�0�v����>�K?y�?7�=2龊���Kf�`�(?�K<?�YM?0�?
�=P3۾�:� 7K�5���X�>2��<�l�,���))��4�:��?��ur>�o���ڠ��[b>w��[޾5�n���I���{M=���4V=8�s־����=t&
>���� ����Ϊ��,J?t�j=�l���AU�_�����>���>�ޮ>��:�-Hv�І@�󮬾\�=��>_�:>��?��ˁG�v/����>�E?�@0?4��?$��P^�9�	����)A��4�=p!?�W�>��"?�A�>�%=�ԡ�w!�&�������>'b�>�~ �9F�%���~R����^��>��>ý�>�4?h25?��?�{Z?'W?�]�>�N�>��t�y�Ͼ��3?^��?.��y��~%v�%�c�x��d!0?�:?<;���> ��>�� ?~I?��@?}X? �=�����+�n[�>s�w>[5`������ՠ>]w=?�r�>��~?q�p?l�D>i�"��8ľ��}�R�=��@>�X?L�E?(tP?�S>Ky�>d������<���>q�U?녁?�@k?(l�<���>ҟ5>���>>�1�>L+�>?��T?�g?�XE?��>7a�<{+���?ܼ2-r�vټi�<��#��C=��ǽ0�0�s���Qs=���<<Ð��8�c����ǼA��8l�=hu�>'�s>h��^1>-�ľ�!��zA>�����[��
⊾�;:�r�=���>��?정>^;#�=���>��>����((?��?p?�f;̕b��۾��K����>�B?�l�=�l�Ur��X�u���h=��m?�{^?�tW����h�b?��]?�g�@=���þ�b�e��V�O?��
?�G��>#�~?��q?W��>X�e�9n�����Db�A�j�ն=�p�>�X���d�q=�>{�7?xN�>��b>#+�=1s۾��w�@s��c?]�?��?=��?�.*>��n�>3�+�
�aǔ���b?���>_:��I� ?�� ��1ž�I������v��$ѷ�c����l���ࣾG@��j��2۽��=c?�v?�jm?	AX?^����\��#V�`r�a�J�e��;�C�@�&L�h�D���l�#�`~��b���#<�`�V@���?�6/?߱I��v?��������u���O*>?�7�r���g�=~��<�-�=@8@=/If��%e�x����� ?��>3�>x�W?z�d��I<�fC6�����˟���J>��>��W>��>��6=���h�6�1������ �Z1v>�o?T�2?��b?A�$>��+���u��}���<�\���a>�b>0{�>;kýg�{�e�G�S�V��	z��S���@��G&�n`�=�)?.�%>w?N�?3F�>:K8�nT���w���L��)��A?�k�?g�?G>U���ƾH��>��m?���>�=�>�.��Κ"�E |�@�Ž4��>Z*�>c6�>�ds>�c#��]��֐�ꎿb!;���=��i?&��Z\�1V�>ڛL?_�'<��<h\�>&Ꮍ*�}�:�3�2��=s�?�X�=�9>�CǾG���{�M����)?@K?�$���(��K�>�j!?���>�:�>7�?��>�u��2�W<�O?�_?2J?@L@?��>f�$=2����ȽB�%�x==�z�>4}\>#/~=͚�=���T�Z��
'��9=��=2���T��F�<����F�S<��< �=>��ۿ��N��̾����G�>���A��˩�
����	$�D_��L&��ޓ|�a���;=�,Da��Qg��J��ȝp����?��?$䍾�����(���#~��������>��j�)U�������
��u�����찾�g&��P�Oj�b3f�P�'?�����ǿ񰡿�:ܾ3! ?�A ?:�y?��5�"���8�� >SC�<�,����뾭����ο@�����^?���>��/��o��>ߥ�>�X>�Hq>����螾y1�<��?8�-?��>Ȏr�0�ɿc���w¤<���?0�@�&D?g�����o��=�V�>�?;�E>�<L�[���iľ�q�>�^�?��?48~=J�R��1��fZ?���;E�п�:"��=� �=%h@=�D�^�%>(�v>ڔ-��G������V>[c�>�x��{���R��'<ʕT>�?��N���Є?�f\�V+f�P�/�]��(p>��T?�!�>1��=��,?�SH�xkϿ��\� �`?p,�?���?1)?\c�����>P�ܾ��M?�U6?��>�]&��t�z��=V��~���㾘V���=$r�>��>��+�9����O�`ۚ��>�=.j�L�ӿ~8ξ���u�Y<�ж=��d����S�
���맠���H�*s�="�=ז'>yJD>f�9>�܏>�X?��v?:[�>R�>0�)��9b��8��s�]��﷾F�׾L�h��R�����0�@M*���/����$��!=���=�6R�f���?� �Y�b�=�F���.?�v$>P�ʾ��M��-<{pʾU����ۄ��ॽ�-̾
�1�#"n�f͟?��A?������V�W��X�r���\�W?P�ϻ�|ꬾ��=����y�=�$�>���=q��� 3�s~S��m2?BU ?��ľ9T��P�3>����w=�G1?ƞ�>ɫ =#U�>��"?w'�U䩽!�]>E�'>�m�>_a�>zS>�����ֽE� ?�hO?�콕��jŌ>�8ž�.[��i/=D >bv�q���K>���<ǭ��t׼�O���
=kVW?i�>Vn*�M;�Î���6�X�S=�Bz?�!?#�>]sk?��A?&��<s%��S�^�9}=kpW?��h?�>��~�+;s�����5?u�e?�fN>�l�͗�-l.�!��~P?u�m?�?�ڗ���|��Ӓ�6��;a6?��h?5D�]���f"?�Œ �}ʥ>�?~�>l��;�?�Ӫ>{H�q����Gǿ�~��&�?�w@�#�?<�o�zǸ����=|��>��?�x����}�.��	ؾ��=�=�>�iľGO�r�9�-'s��@i?��K?���>�bA�]&�_��=���%��?DΑ?�4־^��=,� ���9��~�<^�;�/�>�_��㜽����C
E��8ž�R�lM���vI�}˃> �@��V��?�X����q��E��������n��_�?�&�>@/ �"j�����Sx�b�^���;��t>�/Nv>�K�=����ܾt��'�B�b��;��>Q��=�vc>�E��7��"��t䄽���>p?zE�>�>�8{��r�?Y��=��/z����B�jUI?���?�0�?��R?���>3�k��Q9>p�z>�%?˲??Jg??��=#����r�<%�j?�_��xU`��4�qHE��U>�"3?�B�>R�-���|=�>���>g>�#/�w�Ŀ�ٶ�:���Y��?��?�o���>r��?rs+?�i�8���[����*��+��<A?�2>���G�!�C0=�RҒ���
?R~0?{�c.�W�_?'�a�I�p���-���ƽ�ۡ>��0�f\�O�����Xe�
���@y����?K^�?i�?µ�� #�f6%?�>l����8Ǿm�<���>�(�>�)N>�G_���u>����:�	i	>���?�~�?Mj?���� ����U>	�}?��>4�?;��=pA�>�`>枝� ;[t>7�=Hޣ�_�?�M??$�>���=tL8�&,�'CE�$�Q�P��t�<��f�>�A^?��J?��F>t3��H�������H���K�(�-��B��ϴԽ�58>9�5>TX>�xV�����?3p�{�ؿ�j��Wv'�,54?���>��?����t�
�>;_?y�>h7��+���$��>=����?/G�?I�?w�׾9t̼�>)�>K�>[ ս���.�����7>��B?M�JD��K�o�)�>g��?ȶ@�ծ?*i��=	?��T���8ꀿ���?�4��>E�8?St�3�>��>�=r�u�����s��ɺ>���?w�?��>l?^n��:D��J==��>�k?��	?�7e�`1��&�D>&J
?=�����(�XKc?(
@�@�]?5E��lɿEϝ�G�v��ؾ��=_�*>��C>��S���=1񄽂r�<v�<��g>n�>W|�>��l>�$j>�>5>)y�>a��J(�*S������6�4��^ھ\�a$�E�־'���_�g�Ѿ՟�4X����n�wD̼�T��)�ֽ�K���:Z>�dK?��7?k	c?)�?�+�u��=����	��~*���@>�>�>��A?}�O?��'?���<�����[�aE}�ǚ�J+���H�>0>���>J�>r�>j\�=ɱh>��H>4�4>�4-=�=�[�=<�>J��>�]�>z��>*Z�>�C<>��>Fϴ��1��i�h��
w�Z̽3�?����N�J��1���9��Ҧ��i�=Gb.?|>���?пe����2H?$���z)���+���>}�0?�cW?'�>��h�T�/:>7����j�.`>�+ ��l���)��%Q>vl?p�f>�$u>��3�?`8���P��}���}|>66?�궾�&9��u�k�H��_ݾrRM>�¾>" D��g�������hui���{=�v:?Ѐ?�,��Nݰ�z�u��B���QR>O?\>K=�=)MM>qc���ƽfH�a}.=���=:�^>I�	?S&_>>�Z<���>*���:���]��>�e�>o">8xM?�{&?i�K�����W>�����]>�$�>�	�>$,>��`�D�=�W?�hK>쬀��������O�p�/��>GĽ=Q�ͬ=|s=��߽+W>�҆=&z���}t�=�~?���(䈿��e���lD?S+?] �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>}x��Z�������u�d�#=[��>�8H?�V��l�O�y>��v
?�?�^�ީ����ȿ-|v����>V�?���?g�m��A���@����>;��?�gY?moi>�g۾,`Z����>ֻ@?�R?�>�9�{�'���?�޶?ԯ�?�J>2��?-�*?d�>#5�>�[��8��*4V�7k?8�E=�p�>�*�>a"�<�{R�����!㞿S������
G�>}�/=��>�}�7�¾,ɜ>i���ŀǾ�6_�\B�>��B>��B��i�>m�?�:�>Z,b>��I��은��Ν��IL?��?�M�Km��u�<�h�=�Z��U?�l3?b�'��F;�-�>�N\?e�?_�Z?Ȗ�>8�Ӛ�5~��")����<�K>+��>
��>j���g�M>2rӾB�bP�>J��>U���#�۾C���N}�{��>�W!?nX�>�r�=2�?�N(?Ɓ[>!��>&�6�EC��x�G�oh�>�h�>�P?�3�?X�?�¹���8�TQ��-Q���_�u�.>�\u?�?�ŭ>����<��c��=O��֠}��kv?�r?�ý�9�>���?�_B?�! ?A�D>��(��Ѿjvv��Z�>p;!?�s��*A���%�%����?�?Q�>�R��.wѽ7�ӼW,�����>�?b�[?�&?T+�/i`��þ��<B)�L���;��f�4�>!P>�c����=�\>��=Vm�Ƒ5����<G̿=��>rz�=�5��;����"?�z�<8վ�Gݽ�E�����[r>iE>ڂ�<�o?bپ��W��Ƕ�|}��\��=\h�?�[�?ӛ?����a�d���0?4[�?B?�?�x��M������E���������o��=��>� �=t)�-ݜ�=���8��]����N*�l��>$�>��?GE�>e�>GG�>�";CL0�&�˾��5O���
���?���u���"���<��w�P"ǾB>���}>ݷ�a��>��?��{>��f>�̍>G��=SЃ>�O>ǥ�>R��>x�b>��>P� >v9a=q�d��kR?v1���'�П�,e��5/B?8$d?p�>��k�6����0���?+}�?�N�?v>#h��+�P?�R�>Z��)<
?�U<=����l�<nv�����o��G�6�>��ӽڸ9���L�̦e��d
?��?Ix��j�̾`hٽ���z�<4B�?��)?9&��E��|k�H�8�#�D��4�����G���2&��_�)쎿=��C샿�k!�0�>f�?+�?+���y
վ�b���|�ؼ=��=(��>Ϯ�>�>��A>5�
�+�J��cD���c���?8�?�*�>?R??K�+?cEJ?�aJ?
i�>�8�>�쳾q��>�y����>s�	?�!??�w:?[;?��?C�?E	L>�!�����z۾V�?��?f�?<� ?��?��n�蜝�۬��H�ռn��4��2��=�,�=��üo��-�s<�K�>a"?z�ݽ	�/�8�Ѿ�>/	C?���>���>�=����¾;�`=Wi�>l?l=�>N���K�_�>K�[��>�o?zY�p��=�2>n>����;ł=��W���=�^��8�8�<�~�=ҹ;�F�W��O3�����E�RS���t�>�?���>yC�>�@��� �0���e�=$Y>HS>%>�Eپ�}���$��J�g�`^y>�w�?�z�?��f=��=ӕ�=�|��QU������������<�?	J#?�WT?R��?t�=?gj#?�>+�jM���^�����î?s",?���> ����ʾg憎�3�f�?�`?J:a�����7)���¾�սj�>�Y/�.~�a���D��o������y��u��?｝?��@�a�6��u�ǿ��WT��ǑC?��>�`�>A�>'�)���g��$��);>��>�R?7;�>%�H?٢a?��Q?+�c>T�,�jk���×��&��� >I�L?�.�?�Ȓ?�u?|N�>"��=�n<���޾���^E�lp�&iv��<�W7>ڱ�>�\�>u'�>2 >~��2	��QcB��x�=`�>���>�ѭ>�ݽ>3�>X��=�~I?y��>����2��v�X��u�>��?�T�?Q_Q?�s)�����5��຾��>ə�?gU�?��2?͟���>83���ﾝݏ���>�1�> B�>��#���C=��^>t��>�9?��;�8�<���1�F(��3�?��g?��=��Ŀ�&y�S�p���������xe�`5T���n����7�:-��m;^�\����yf�������ԾD�ξQ��0<���?z�3>#�>4�=	w���_x���*N6�֒�=�m�=�S��3<�-��)���#���9���T5����<B��=��Ǿ�|?bH?�~,?��E?�ɀ>�f>�I�	��>�Ȁ�Ɇ?�J>��:��޴��s5�D?���3%ྡ7Ѿ)6_�6ӟ�l�>�'�<� >{�0>���=2B�<
��=��=�zg=Vw�z�C=)��=^o�=�>�=���=т�=��>NGv?�����(	R�����x9?:C�>^��=�����PB?g">S܂�kb��(�����?0��?�k�?��?7�r�/<�>e����YP�'�=���6z.>V�=H�2���>]�D>��n����7Ƚ�?.@~q;?zM��klͿ�#>��/>#�>��Q���0��^W�AKQ��qD��?K�:��F���9�>rK�=�۾��Ǿ��S=��F>]��=���E_�Dq�=�+~���T=��+=��>Y�A>�y�=`���G��=p�Y=JP�=KqR>9�(�������Ȇ= ��=Du>R�H>7�>q�?m0?zd?���>9Nm�yξ�v���ҋ>���=���>콅=�nB>�9�>��7?*�D?��K?+�>�K�=�Ӻ>�ަ>�e,�S�m�{��֧��p�<&��?o��?�ܸ>$�[<PMA�����=�#(ý��?��1?�? ��>���]��8���0��a����v=�')=�'��_{<{@H=�����W���0>.��>�$�>��>}��>�;:>NLk>^��>�=Ǉ=�� >�Í���<]T��\P8=2�ٽw�=���
렽:�<�:�5Q��1�<�ݫ�j0x�0��=l-�=
��>'�=�x�>ű�<30���h>m�ξ
U;����=�f���=5�(oZ�m������s{���6>J-M>N]��T�����>3Q>�C�>��?[>y?SW|>�g���!�z����K
�h�2����>eK�=�,���
5�B�w�t�R��M���>�ߎ>��>��l>,��"?�,�w=V�!b5��>|�����T)�Q9q��?������_i��Һ��D?gF��ٛ�="~?��I??�?���>O���ؾ�90>mH��H�=i�L)q��h����?!'?e��>a�D�D����d
���>vV��J�r2��V�?�Y�T����Z�>�����}�-BA�HҀ�}����L�S���>�[?J��?g2#��De��8�;��S�����>v�L?<�>{�>�?m`��x	��m���X�=�w�?���?��?���=��7=���Y٬>H��>��?kK�?[ot?��]@�>���=ν�=��y�kB�=F�Z=<~�=!�Q>yp?b�?��>�O��A� � V˾8��{���<?�=R��>�5�>g��>�q>�Й=Ɵ>=�Y�>�{�>�C�>�Ƹ>
��>m��>����jR?���=aaD>iUE?Ѷ�>"�:=�Ƕ��/û�&@��������Ю��;�?>M��=�`�=�+�=e��>��Ŀ`?�?���>Eb��3,?�&���g>z�
>��N=��=1�>R%O>iy�>�|�>�Q=>up��/�<�9>]NӾ'l>j���c!�,C�3R��Ѿm~z>����� &�w��ߋ��`KI��n��hh�}j��-��<=��ٽ<�F�?�����k�@�)�R����?�O�>6?dь�m눽��>���>n��>�K��7���Ǎ��e�1�?_��?���<�?>�K�?�C�>��M�k�c��6u�Mp��y<��y���)h�b���7H��!���졽URO?�M_?O3Q?y��=;��>[�f?̪��r~��?>U��/����`=�_�>x��0��ʣ�I����2�q�a>7z�?S��?�8&?Y戾�H3>��>[�>8?Of?8�6?�-C?��#�:��>�IE�Ϥ?-$?}3?d�Z?j
 ?V�H>_:�<^g�~�=��7�crt��f��s���t~z����=ѱ`��R)�NF��mo��=��1=)	F=�꼆W;���=�O�=7�d�C���9ʐ>�S?�`�>h2Z>,?��ν��&��u���?�X�=U ��ˀ��ԡ�(L���#>C�t?��?�{]?2�_>Q�<���U��[H>�ɘ>��>�A]>xx�>l�o����S��9�>t�>^=�=�q�~����W�S��|���8e>��>�U|>򀎽Rf'>4�����y�ve>��R�����;S���G��1�0�v����>�K?y�?7�=2龊���Kf�`�(?�K<?�YM?0�?
�=P3۾�:� 7K�5���X�>2��<�l�,���))��4�:��?��ur>�o�����;>�=���Ⱦ��\��J�9��G)�<���Ƕ<Σ�J𭾈zF�)�>*z>�︾5 '��љ�{��|�E?��=ua���d,��7���Z>�>��>,O��f���+H�^��w7�< !�>��/>li*�?��ZEN�����ϕ>�DM?�?��~?KQ���&*�L�a���۾?����־=s?uE?�>W,o>�7b=��8���N����Y���>-?��;�t#�f،����~���i�>�@?b��=���>��V?T+�>�:�?�\C?M�?�Q`>�T��}�ᾱ�)?��?�q�<��½ٷe���<���C��?6 9?�`����n>�?6�?�{4?�T?�m?�ė=c����N�zG�>�!�>�Gd��Ѱ��[j>�s@?U��>��W?4\�?ReQ>T�?��_���'i��C�=��4>�B7?3{!?�A?��>��>j롾3�=#>�>��b?��?��o?�$�=2�?w�1>��>ω�=�?�>3s�>�?�O?!`s?��J?M�>��<F����1��|�s�$%U��\�;S�I<��r=�]�s���r��<l��;bt��B�]�6���G��`��x�<0�>�s>i����6>�鮾V녾�L>����X��Hsa�:0�w[�=�Rs>�v�>@l>i��I�j=�!�>��>����%?�R?qi?�;��];[�1�����E��>9?��">64p��+���o��`�=��h?�*_?��+�$� �n1`?#�q?4޾͉��vϾQ$��P�J�U?|�1?��۾���>��}?�eS?O�%?�L⽧c�8Y���t��^�ؾ)uO>��>rX��hq�q�>h��>�	?��>ݰ�>zX��<�!��Q#?�?��?v�?a�=R�a�~Mҿ����둿"�]?g��>����!?ǽ�9�о�T���^��^^ྜ������?���i��U5#��k��Fj߽�
�=�?�@s?Rq?a�_?;� �oc���]��~�ѮV��%�H�kSD�(E��B�w�m����Ο��{���7=.ہ�C�>��`�?�?нֲ�>�s��H����3Ծ��?>Ĺ���0��v$>�y�c=B=�fp=Aǉ�f�V�����9?^��>�|�>��=?�U���8���1���*��|����=��>[ɝ>lX�>�R�$I'���ؽ|�ľ�h��Ҵ!���{>QY?�!a?Sd?OU���HQ��k���J�N����<>Dc>`��>�.l��b���@��J��Iw�����⓾j���(>�l?uo> ��>���?��>��Ҿ�S�����+?	�U�X��4?~`v?D%�>dVW>��#�C�$����>�Iu?��?��>/ ���3�M.��(x�=�Vq>�̚>�Y?|E>�v���p������]���� ��ɐ=�4K?�{��:�
�>���>1�=�K>�K�<�*�G���ki0��(��"G�>��2?A3�<�T>���WWC����C�Ҿ�p(?>0?�㏾�$)���>$?Q�>dB�>FL�?��>c�¾�Ȣ;�?q�_?�@J?<6??g��>ٹ"=���)Ž��)��6=��>��X>�6f=:��=�U�K�b��!��T=�=p�������C�;��м"~?<��<ez?>�Kڿ�K��ؾ�X�_�ﾕ�	�Z>���˾�_�����v�����4j���	���lsS�4�g�ũ���o��~�?[R�?�����F��1ә�[�������(�>X.t�����%��v��ެ��3�ݾ���'C ���N�n�i���d�L�'?�����ǿ򰡿�:ܾ4! ?�A ?4�y?��6�"���8�� >]C�<�,����뾬����ο@�����^?���>��/��p��>ܥ�>�X>�Hq>����螾�1�<��?7�-?��>Ɏr�0�ɿb����¤<���?/�@tyA?ۙ(���YrV=�S�>�e	?�@>c�2��q������>|�?��?�F=��W��*�>e?��<��F�!�׻�O�=�g�="_=h�k�J>�>�>�w�5B���۽Q6>�i�>�(�[�_�]��p�<��]>zeԽ:[��>Մ?�z\�tf�R�/��T��ZV>��T?*�><9�=β,?�7H�z}Ͽȯ\�H*a?�0�?&��?��(?�ڿ�^ٚ>��ܾ��M?D6?��>�d&�j�t�'��=C5�T�����8'V�3��=��>ƅ>ہ,�����O��R��U��=�i�Pv����g
���=��#�z}��:���Ҫ���¼N�h���b��<�C�=T�:>��6>�#>J�>Zq%>�&P?�<x?֊�>��=׽���GY�p�#������IX�t�<TI]�|�о�������e�d�"�������@�&�H=�T�����_�$��6`�
�G���'?r�*>�ƾ.�N���<��¾����G�A3���̾��0��"k��Λ?��@?d�����Y�b���jѼ��Ͻ?-S?h�?��[���'!�=ۑ⼦�=L�>�f�=)S޾�p1��#L��*2?��+?|ܾ��Z���P>G4.����=��??��?�i���?�>v�%?���]Έ��Ђ>c>>��>���>$Ķ=#mž�'2�g�&?~�Y?�x��&X��E�>�u���N�����=�;">[K�8Y='E>zc&=����<�o���r=(W?��>��)�����b���>��C===�x?�?�/�>�zk?��B?:j�<�k����S�|��rw=��W?�(i?~�>6���о����5?��e?��N>�_h���龤�.��S��'?.�n?�X? ����v}����i��{k6?��?�@�4���5$ȾFg��'o?E�`?�em={5x��{,?�f?��ڬ4�����3R����?'{@E��?0�K>���^r>��?��>?�Ͻ�ݯ�`���q��>��>H`-��lw��75�����P?�(�?z�?�/����۾ �=핾)F�?��?\8����b<���ml�[t���$�<]R�=R��! ������7�ǹƾ;�
�>����ü﹆>N@0m��O�>J�8���,@Ͽ����zоo�q�;�?�>Reɽ]h���j�*u��G�9�H�1���>�[>�o��	����{��
D�Cx�;��>l��Z�>-�)�O����"��lG���*�>J��>���>� H�q>���e�?����[п!���
n�i[V?۩�?�q�?�:?=0=<�o�(N��q�=a�2?��W?CS?ڷ#��3-�^��:5�j?fY��K`�p�4�S>E�5U>�"3?!.�>�-��}=�>���>\g>�(/�j�Ŀ6Զ���� ��?���?Qh����>>~�?|y+?�q�l4���m���*���=��7A?t12>Y���_�!��.=�>Ȓ���
?�~0?�e��.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>n��?��E=��?�w>"�Ծ(=�>U�?>#a��:��>kXO?���>WɆ>�2�<��"��.���8�S��oJ��R?>�|?e�J?t_�>KYB�.��<l��yé�/��������Ж�HO�>��2>�uP=����׾"C=?uL)�Ľ߿B+����x�[�P?�!�>E|�>:$�[*�Iw�=ʛ/?�?GX ��ڻ�It������?�6�?�b?ΒϾUJ�3��>^��>�<?G�	�s ���ص��4N>��+?>hD�;���B����>+�?d4@���?s���]1	?�!�SW���I~�т�/�5����=Q�7?�t��F{>��>9�=6v�3���o�s���>\J�?��?,��>}�l?�No���B��_3=>\�>��k?`h??������LC>�?���i	��7T�f?��
@�{@]�^?Q�����п��W�Ut���T�F ]=��$=	K��0>�3�=���݇��r>�q�>��{>�/^>j�>�`>���=c���U����z3����B��6*��sԾ�2ʾ�N��
�/�ʾM믾V&Ҽ� ��V��S�I�]M��̖=��=�]<?J�Q?��o?uD'?��?����=?o=����=��i�q����?�>$U�>SI?`�??���_Ѿ�Et��rw��������Pw�>�qB>6��>���>���>)�>�[>��A>�#M>�Xh�g����
½��=Y.�>~ ?�?�>�}?>�u>ʹ������Bh�!�y�U,̽8#�?�P��p�K�~������������=��.?�y>O)����п�y����G?U瓾u���/��	>�I0?�nX?��>��)bG��s>~�� j�E��=�O���yh�u(�݁U>�?��f>_u>�3�{V8�
�P�u��~H|>�+6?�ⶾ�[9��u�o�H�DdݾgLM>�־>��D��k�|���W	�aUi�Q|=o:?p|?I_��e�őu����,AR>$R\>��=��=M>Boc���ƽ�H���.=��=��^>�?��4>��=�6�>�Ƌ��CQ�] �>��>��>�SA?��?b5K�z^���-��"HU��2u>��>{��>-�
>3HB���=�>��>-����o�ve-�W�!�*v@>������5�ք����<<�����=���=��0�/��#=�~?���'䈿��	e���lD?R+?] �=;�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��H��=}�>	׫>�ξ�L��?��Ž7Ǣ�ɔ	�,)#�jS�?��?��/�Zʋ�=l�6>�^%?��Ӿ<��>���~њ�,i��z��Ϋ���g?1�P?h3	���>�m�3M�>	�8?�]�伨�L����R��^? |�?��?Uꑿ���k8�뢱>���?�*�?��>��%��暾��4>�?2_�?f�*>�N��L½5��>̙�?JȒ?m=K>�K�?x?8��>M剽��'�V��¥��3~=���x�>�>�R��͘B�!'�������k�6a��N>��4=��>�Eٽ.���8°=�w�*���������>��S>9SF>9d�>u[�>�*�>h�>�",=�v�����(8����U?��?�[F�a	9���f=�1νl޽�4?���?�Ğ���Ý�>u9*?V��?,{d?��s>���>B��-̿&1������cK>� ?�?u���Ȍ�>#���9���>Qw�>.$P=F�Ѿ�������\EO>UK6?kA?3	�>�� ?5�#?I|k>�M�>�tE�@E��<�E��n�>���>\7?U�~?�x?����3�����ġ��[��QN>�x?��?�A�>�A���k����2�#�E� `���Y�?vTg?����y?<�?��??~�@?��e>� ��^پ�,���>�!?#���bA�'&����d?�&? ��>8'���[ֽp�м����r��I�?�/\?%&?k��.a��¾���<N���ni��;�;��H��%>�Q>Yl���r�=>�ӱ=�Sl�]6�{b<�?�=���>� �=O�6��H���cH?R)�=�R��q->x:U���[-�>we��+žq�x?��S��������=���Հ��ϸ?`[�?�?�Y.>%Mg�D�H?�̃?AT�>f9?fn&�vӾ���6��D���W辛qs>�R>�m�=x�̾A@��F�����e��~���>tT�>���>�}?��>���>vcȾ�V)��v����$�J�N��7A��uA��������۽�%�7���|���ȕ>�]�>9�?�t7>W�O>4��>���<���>� �>)w>��w>���=X�>��-�q��<��]��KR?������'�@��Q���N3B?Zqd?�1�>�i����������?���?Rs�?�>v>�~h�u,+�Cn?e=�>g���p
?�\:=��K>�<�U��*���1��}����>�A׽" :��M�[nf�1j
?/?����̾R5׽�L���n=�;�?l�(?]y)���Q�rvo��xW���R�"$� Rg�_����$��kp�Ѵ��/��
	��;u(�o�*=c�*?��?\~�28	���>k���>��\g>Ͳ�>�ٖ>�l�>��G>��	��1��^�='���0�>1#{?�֍>�J?�:?��R?B�Q?U��>)@�>���tN�>��=<q��>=i�>��6?Tn2?)\5?��?��#?}�T>����K��<
ھ �?g�?_�?��>���>P���Q�Ž ��!ջ&no��[��u�]=�<ֽ�n�=�M=�?]>:E?L��-8��S���
m>p,7?`��>�;�>�����P�����<���>�
?��>. ���q�9l���>я�?���]� =X�)>��=_���Xc����=�ֿ�K��=�����6��|%<���=�ӑ=us�3��9\$�:��;��<�?
�K?��>�R?���$���F3>[x��j��>|M�>d�%��	��Qg~���y����=-ƒ?;ڨ?T��<�e�<��J>[��i���R��v������cv?�?ZA?Z�l?�A?��?�|>�2'��{p�%�ξ��.?~!,?N��>���V�ʾ��ɉ3��?Z[?a<a�ܸ��;)���¾��Խű>�[/�5/~����D��򅻵��U�����?�?A�0�6��x辩���\\��u�C?W"�> Y�>K�>F�)�J�g�X%��1;>��>bR?.޻>(�O?B7{?�[?.�U>�8�J�� ���r�+�-�!>��??5��?��?	y?���>3�>�1*�+��s��I��U�e��UcY=��Y>Og�>)X�>��>���=��ɽQ��2�>��O�=U�a>$9�>� �>&��>>w>�S�<��G?���>~O��V���󤾤ȃ�O=�.�u?p��?��+?2�=�� �E�MJ��{<�>�k�?���?�7*?%�S����=��ռ�޶��q�8�>�ӹ>g*�>q��=�F=�Q>B�>k��>J7��V��m8���M���?pF?H��=�m����`��쩾�6�Vt5�G맽&	о������=w���19�^�5>�h�}^%�!*l��;���I����y��a= b�>mhR>��#>~Q�= �=�#콇�^=��4>��o.�=< �=(��<ĥ	����ؽ܏����C=`��=�q�B�;m�b?*WH?{�"?w)I?�|>�>.�(<��>z����k	?L�P>4ӱ��x��.N@��A��a1��G|ھ$�پ�[��Ӧ�K�=����R4�=�D>�'�=ѹ�9�Ҭ=�r�=��>󒏽c��<��	>�}�=m��=�H	>��~>��0>�Kw?���)����Q��k�p�:?F��>��=+�ƾtB@?��=>UL��'l��3��u�~?���?i�?��?Qzh�f�>����hč��V�=����:�0>$D�=.�2��Q�>=J>8���A�������?�{@|??OӋ���Ͽ7/>��1>m�=��O��K0��iT�0�^��W�(- ?�:��˾ɖ�>�/�=]�޾ �þ�|D=�4>ǷK=��^Z�c�=�w��M{)=��e==��>��B>�'�=�뿽�=:.L=���=t�U>
9@�
�<�����G=��=D�a>��+>6��>i3?m:+?g5N?��>������Ⱦy���V�[>P��=���>G�=�@�=�C�>��4?o�1?��0?�6�>�i�=���>g��>B�)���^�&����� 2�=́�?=Tt?D?jd�=X��`:�U�9�C�����>��9?�Q1?)&�>&�ι��B��l��b�����=�S�ۉj���9>s�ͽꄒ���=X�=H�>���>l��<=K�= !>h1�>sދ>#V!<���=L٠=u�=�8=�_l=��>7�����j�7��;R	����<�T��'�=Et�=�倽{?��K6��»>cf�>�+>�Y�>���=g��4?>$Ȣ��0N���=�����%E��s\�at��LL4��I'�	�X>�`d>N,���L���_�>LCj>\>N$�?�0n?�>���h�ξ���xG��`��-��=�F>Ck���G�K�q���E��<Ҿ���>�H�>R+�>�n>�[*��%>���l=��ᾠ�5�c�>�����ʹ�pr��]��X.����h�sպΒC?����iG�=�p}?t�H?�*�?���>�>����վ�v.>�兾ۥ=����{t�xԋ��)?A�%?���> ��hE��ݲ�F�Q�H��>��;��wC� Й�s��U�<������>zBd�iξ&�.��2���~��3�}AP���>��I?�$�?t�'�c�����L��7�D��a?�8l?{�>� ? 
?[jb�o�������Ɨ޽�V?�b�?^4�?md:>�|=����a��>���>�+�?�G�?�ad?:�,�-�>8�.���>�r��)�=rD>�T�=qܲ=���>5U�>�	�>2&��(��������Dp��7=��=KM>��W>�~>��6>V�=�
�=�T>r��>B�>@o;>;F�>e��>�¾j���?x�a=���>l�%?]�P>3��=�c�� �]�F=y�4���E��0����T
��#�=}5U��:�>�O����}?6�>-M����?�6��W��A>@�x>�5���/�>��{>�Ɏ>~�>Pq�>���=-K�>��=?�׾H�	>ӳ�ϔ#���E���P��iӾy�n>Bٗ�����I�����HdC�������4�g��Ԁ��;��Q�<���?�N��k�%�*���??	
�>�/5?b~��y����o>��>@Q�>H���������4{ܾ���?S(�?�ڗ>�c�>$r^?�m$?ܷg�ۺJ��dC���a�Q�X)+��"�_Ə������]'�{�b���O?��g?�T?�bD���]>:�?)
��"%�lO��#�9?���>���>rRҾ��������&�<H�u>�#=?�ƍ?"h$?��|���:o0?�?��?.�
?4�?�[�����>7�=��?��?��>Lp*?��@?�	�=��1���弻�a=���響�3Q:�	ʆ�L��7�[=�]=H^:�;�\�C=�~�,�>гc=���6��=�y�;C��=On[=�)O>��>$]?�I�>�1�>��7?�2!��N4�o����*?�^=岃����� �������^�=*]h?KS�?o�Y?��d>xLB�hEH�R0>�\�>!~*>�W]>���>z���$E��4�=��>hS%>��=e�W�#���9p	�2����^�<#�&>l��>#F|>�����'>Gn���;z�I�d>��Q��ƺ�]�S���G���1���v�lR�>��K?^�?
��=�V�X9���Ff�O()?P\<?�KM?�?S��=B�۾��9���J�;,��(�>��<���ܻ��0!���:����:0�s>+*������Ti>�_
��Bپ�l�NI�����^=�����0=��
���Ѿ�7z�J��=
�>���a�!�5�ڪ��I?�uj=I˨��pO�M컾��>-��>���>�*�#r��#?��ӫ����=�g�>�D6>Cw����{�F�����>�XT?�PV?�b�?P�"�эV�j
G�`��a��� F��,?�Z�>R�?�D7>�)*=��Ͼ�0�5~����`�p��>P��>��(�Pr��ܾcv뾦�����>~*�>�
�=���>=�5?C�>h�c?G�?���>�9�>tR�������?�5�? !�=5`���\�9�!�ֺ5�'K?�t8?�W?��Ѡ>�=?�/"?��%?�I?�%�>���=�\پ��)�c��>��>T9Y�J����2>��@?U�>,�U?T0�?�I>>7<�����L�=А7>�2?UU!?<�?���>f��>�ݟ���=���>�b?"�?�o?���=
?�V2>T��>�`�=�>RS�>N;?L|N?�s?5�J?_�>G��<J����2��S:|���F�o�;�}1<+�|=[l��s n���(�ۤ�<MD�:�\üK|g��伞D��	�����;���>�ut>Xٓ�3.>PžJ��G?>bɼY2���Y��Rf?�B��=p�x>[7 ?,2�> M!��Ս=x8�>0��>O���v&?|R?̏?�]��b�|�ھ�8H���>*�@?���=0n�jR����s���Z=��m?��^?�(U������b?�^?�*�s�<�j�þ��b���[�O?��
?�H���>i�~?o�q?���>{f�f-n�h�� �b���k����=�E�>i��Ɲd���>Ij7?��>z�b>���=j7۾��w��R����?E�?�ί?��?Fu*>�n�<�	��?n��� [?sA�>
���}�?�s�־O菾�'����������0���N��������I�����ڽ���=�?c�i?$8u?-|h?�8� �c��[��v���S��\�ڵ�XpM�OF��L;�S`l�2E��/��i��h�=��z�Nm?����?[�&?id5�X4�>�뗾���(Gξ�<>B:��~�!�f=�=t��"�6=�h=֝g�Zm.��9���:?��>($�>rA?��[��y>�ߥ0��5�i���z3>�Q�>i�>���>�>�;�0��ս�¾����S,��n�u>�fc?7L?�Pp?GNǽj�.�l,��t���T�Rȭ���N>�K>F�>��R�o�.�2�&�jD���z��_��l��G��aA\=�)?���>�ח>�L�?�A?� ��ں��Ѐ�C**���<���>�}e?�z�>�s>N���2"�7��>�'c?�
?lf?����M^&�.�s��k��i�>���>�b?k��>�a|�`^\�>B���݉�4�,���ݼC`?�E��e�)�='F>�]?�W�>��=~��;M���hFپ����].���>��F?>��^>�ָ��6�[0���6ľ>�"?%�?R_�]W)�	&�>_	)?5��>c��>�5�?ic�>E�ʾ�.~=�a?��O?݇K?��)?�p�>x=���ý���n��=>��m>��=��7=�;���E��V���J�K���Ľ���w�`<�l�;���M;r�IV�=��ڿ�J�L�ھz��bN�F�������������a��˂��rW���5u��<�^�,�Y�L j��&����d����?Ͳ�?O(������o~���(������s6�>'�l��h��۰��A��;)�����*
���~ ��qO���i�OHc���'?�㐾�ǿ����pھ ?�m ?��y?�4��8#�3�8�n#>��<�䃼"�^���̶ο�����_?���>>��jܪ��E�>g%�>m�W>��q>/���3N�����<��?��-?Y5�>��p��ZɿXm��,ީ<q��?z�@�aA?ߨ&�M��GK=���>)�	?�SC>+(�'�z`��c�>���?��?�v=�@V�̓(�Ӄc?ce�<� D�������=4i�=:�=�r�5F>Mu�>u���zF��@�/�2>�a�>���z|���_���<� ^>Q�ƽl|�����?�GT�D�n�Y�N�Ǌ��t��>'`?3�s>��H-?z?�oN˿A�S�6�L?�W@,r�?��!?�Ѕ�T0Q>l���Ua?X�>?�V>�W/�:芿�hӽxE>ۨ.��m:�B�g��rw=�ϯ>�.�>:�M���!�MK���_�����=����oÿ0-.����� ��@���2��g���
o��dŻ�]�J�!�w��һ= Է=��=�X8>��>�eL>,WL?.�r?^װ>��&>�^r�����*ݾ�Ȝ�$]���OH�MJ�������r���ݾǏھ�[�cq�:��z���r=�b�=�3R������ �}�b��F�$�.?�q$>��ʾ��M�n2-<xqʾ7ê�lЄ��ݥ�|0̾��1�5n�Wʟ?N�A?��V����n�s����W?T>�����謾��=t���B�=��>n^�=����3��{S��i-??�?>q��떾T�M>.	����<��2?UH?)4�<��>��#?�n�|Ƚ�Nu>�%>��>��>_>J@���ѽ%�?�iS?�0н�팾~F�>�����*r�(w=g�=`~s���@�Q�F>5T<�4��g��U'ڽs��}�V?ֵ�>|^(��p�/������D�N=�x?o.?�ʘ>��g?�zD?� 	=4�w�Q�sM�; g=�X?��i?�D>�P����Ծ\����4?<b?��T>uMZ�ѧ�/.0�i����?�'p?f�?��*}��ˑ�����n5?���?�Pk�J	��l%�1���d+?}v@?C^>>��`�.�?�dP?�]��Fw��ο��/��g�?3@�,�?%�s>NL=і�;���>�k�>QMt=�F�\�<�-L�D�1>�?�����-C�~�	��v���W? ��?$y�>�vt�_�����=�ԕ�[�?}�?&���i_f<U��Ul�xk��\��<8�='���"�h���7���ƾ�
� ���䊿�r��>�X@IZ� ,�>E8�4⿯SϿ���3QоiMq�8�?���>ȽU���$�j�MSu���G���H�柌�/�>"��=�+S�@G���{�ܡE����=y��>�툽z��>�)�m�Ծ����27�!+J>�>T��>[���$0ʾ�A�?.s�0ӿT���r:'�8Ey?Qo�?='�?i��>5��=�ǽ�������='�2? �m?�d?�0=d�M��7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�^�_?*�a�O�p���-���ƽ�ۡ>��0�f\�WN������Xe����@y����?O^�?j�?е�� #�c6%?�>Z����8ǾC�<���>�(�>�)N>�G_���u>����:�i	>���?�~�?Tj?���������U>�}?{%�>�W�?��c=�<?��.>O����B���y>���>c(S����>��P?��?���>�ڢ�EL'���.���K���r���w?
>�P?Q��>�K(>�L<N"���	�\�Z����=�">ݸ��,�l=��ҽ6Q>h��=�>�->½���?Dp�8�ؿ�i���o'��54?:��>�?����t����;_?qz�>�6��+���%���B�c��?�G�?>�?��׾�S̼�>?�>�I�><�ԽR���X�����7>/�B?U��D��h�o�r�>���?�@�ծ?_i�7?�d�N�~�����/��
����>x$?+� ��'�>��?���OGU�����$x��d�>��?�>�?<x�>E&�?-E����s��Y�=�"#>!�?��F?�/��1�� ?��*?������E��R��]?�@" @[�<?�D\�yؿ���&ʺ��b¾���=��d���c=�창�Lw=���;�H��Ϙ=��=��>)�>��>���=���=Y>'=S#���.�{>��m ���yP��6�$���6�r��ś��s���Bw�����ID��Z�����O�z�	���U�s`��`>��X?��H?�s?Ţ�>jׅ�z�>��澎'�=(�:���=��>b2?�J?�:?9.=�1��8f�}����ҡ�X!���ſ>B8>���>���>'V�>�4��Z6>�Q>[ �>qz>�7=g6;8=��F>3��>���>oĺ>D<>�>ϴ��1��$�h�w�̽�?����}�J��1���8��I���cj�=�a.?�z>���,?пe����2H?����)�Ÿ+���>5�0?�cW?ۜ>���y�T��9>+��Цj�a>\, �a~l�<�)�u%Q>7l?��^>\r�>K�&��V;��
C������w>��?���r@�3����JM�����A>�>��	;���i���0>w�{�J�-�q=!?@?k?hH�y`��8��������:>�,>��=lS	�� �=�ɼ5��O�M���=l�>� Z>[)?�z->7�=Av�>5M���BN�=�>!�B>��,>ą??�)$?K��p��Z#���,�ցv>n��>�Ԁ>zz>�-J��7�=Y��>�`>u���l�����Ђ?���W>cw�~^��v�[r=,���!�=!��=���p<���"=j�t?1��G�w�	N�bӢ=4>C?Ў?��\>iV��E�	����
����?��	@f?�?H����J��tA?
T�?�����C==�">\!f>�����;u�3�?��= �ݾ�p��� �?�ߣ?=�����j���$>es;?ﱾLy�>���L������u���$=���>�IH?�[��eS�kp>�~�
???���&���8�ȿ�lv��1�>��?��?i�m��K��@@�0��>���?�fY?��i>��۾1�Z�z�>��@?�R?V,�>�7���'���?�ݶ?���?��9>�ψ?`=z?��?�h>�N��#��$Bg�V�f>=����>�@Y>�S��=�)�j���Qz�M���IM��2�=�S�<�>jUƽ �¾��>A�=�4���Ą�Ab�>9|�;T>x=d`�>���>���>���>��=�ߧR�w̾�J?�?��" [��a�<1��=@�^�4L?�s8?�zM��	ȾW}�>��X?�P?tO?�>�r�%c���N���ɪ�d�g</>���>���>��s��lV>�־e69�I�>6��>�)���qԾ�=w��vؼ��>�}"?l��>c�i=w�?#�#?UVx>x�>l�G�d֑���D�<E�>%��>&�?%g?��?�����4�~���j��.�X�'iM>�y?�?�f�>���������9��(������?9g?sV۽B?Ft�?�E?z=?��b>�%!��k޾G���=�y>�4 ?���O?���&�.r
��?�Q?�I�>/Ɛ���׽��Q�;2�Ƒ����
?lLZ?�%?���_�`$þX�<�����2�;3��;~���>�>L���0|�=�>\�=�y��8@�JV�<ϭ=�c�>t_�=	2�����C�+?&w:������=��q��sC�2 �>�G>�bþ�^?��A�-�{��ڬ�xq��$S�	�?�4�?�ܕ?@��.Fh�e�<?���?י?�2�>4����ݾ�ྙ�p���v����L>���>�ĥ�"羬���s���O@��4�ƽ]��#�>�Ķ>w�>���>1OL>�ڬ>�?��i"��۾�!8�!_���!��D�����}򾖊���RM��"�'��͋8�硷>�mڽ�	�>c�>�%3>ɐn> ?CK$�z)�>k�	>_L>'D�>���=���<O%:��e<_�&�2�V?+O�CtH�04���T6=�=7?n�i?�:G?ޓ=��7��#���_Q?2P�?���?�J>D���a���M?ee'?�i�0��>�)Q���$����=�$����ݽ4!>k�y��W�=�׼����<�^%�>'�>]:_=)%�:g���Ee=	��?i�&?��(�#�T��Vo���Y��P���=d����t�!���o�����F����`���#(��$F=)/)?�ԇ?�X��!*�e����i��+:�.�S>Y�>ä�>#��>��9>Z���1��_^���"���r���>�6y? ��>*�I?~;?�K?�L?�œ>��>�������>��$<��>;3�>�	8?�l,?7/?�s?}�&?��_>���2���آԾ�?+�?7�?~? ��>毆�ν���N������r�<Fi=���<�ҽ����;=3=SE>H�?W���;�z�����>4�6?.��>���>u������J��<���> ?ژ�>����wnt���
�q�>%��?������<>O��=w�>��*���վ=�Z0�J8�=�}��E�2�3E�;>��=��=������ֺ��;H݌:9��<�?�>r/?;b?�s	?5.߾VJ�K��b��T,=�%�>K��>5��������w�u�z�hx�>쓅?߄�?�g*>�j�=��Q>P�~��Bm����,Ͼ�w½�]�>d�.?�=?�*�?��?ܽ?�3+�z���7��0_s�t씾�%�>@,?���>�����ʾ"娿�o3���?/?\7a����L)��¾LֽK5>�K/�~������D�I�����p�����?՝?��C���6�ր�㣘�'h��<uC?!R�>�Ȥ>I��>��)���g�)��Z�;>#t�>�R?�ݻ>n	P?!�z?9L[?n�Z>�7�ő��h���঻+>??���?�s�?�#x?R~�>u>�1���k9��U����𽠝��O�P=�W>�D�>T��>y=�>O]�=@ѽ�c��,�<��Щ=�id>�|�> ��>A��>w+z>k�<��G?��>�e��>���X��䧃�#�5�zgt?�܏?�c+?��=��A�F�҉���B�>\�?\ѫ?lS*?q�O��w�=̪¼������r�r�>���>�	�>M�=I�?=N- >\��>���>r'�D����8�D�T�b�?��F?�b�=�к�<.c�����IO��2D���e ��]���\�l�N��8a=����U
��OE��7��>���7þ���
$��]m�����>l��>��>Wq�=�3=��;��'Z=�iV��?��9=���{���r<OR5�v�j��mR;Z���E�<�=�k���/{?�rZ?'�"?']L?��>]��<�o:�x�>�M��N�?��>�{=IV��+Q��j��P�ʾ}�ݾG^��d\��җ�{!>��q��>!�J>M(�=���4��=��=Bl<�_����=zXn=w�>W��=?�=�6">��B<9��?`���~J��SG������|?�Z?�/��������?wk>̹�������K�0j�?Q@��?{�?�f$���i>��@���(=o����9
�@�N=)��:��?�n�����N9���_¾qq�?Hx@/?y�����ĿL�2I7>�y>T�Q�t1���Z���`��Y�=2 ?�:��)̾K��>�ʴ=��߾�Ǿ��.=Ʉ6>g>W=lX�Q\���=*Tu�f�E=(�j=?͇>d�B>�d�=�د�ƒ�=E�A=��=6IJ>%;�4d1�5���(=���=�jc>��#>oG�>>�?�0?��a?H��>'�\�[ʾ@V����>��=���>~c�=��R>��>Z�4?<�;?��D?�Z�>�m�=�]�>� �>�-/���p���A���?�"=��?��?h��>:I�$�5�� ��Z:�om����?`u1?=�	?+�>���.��B�܅Q��}��fE�a�.��0<�dw=y��=���<��_;!���ё�>R��>u1>��>��t=�>���>¨/>X����Y?>ȶ����=�j������<.u>!'>T���X꼍ز�㰌�[����VѺ)�;�%=��=#��>�n	>!��>�=�e��_c4>-D��4EQ��%�=AMþ�$C�Mc������%�����B>��@>d�W�O͎����>�]o>�+>���?5�j?�>����W���ۘ����	�4��<�=���=z�\�F#C��Vf���M�u�־[��>`�>x�>��l>,�'?�q�v=��(T5�s
�>(e�����B*��4q�j>���🿆i�����D?�>�����=\!~?D�I?^�?�x�>�?��ÀؾJ0>�S���l=(��q�
1��
�?�'?���>\쾁�D�$��*ƽ��>aw}�k���|��l7�E���>���8�>Qe��M9ھ;�'�	[��PH��Ş%���ν�m�>��@?�%�?�[��X+���V�y��^/�+(E?�zc?d>F>��>�J�>�־�'!�ے��j�<,�?�)�?�A�?݌ ����=����H�>JV�>��?Y?�?�f?ٜ����>����;�=��;=E�Z>�Ts>���=�<6��>B ?>	?�����-���}���[�C:F�Q(&>*�>�P>�V�=�׻���=��Y>V��>�(�>d�G>��^>14�>n�|>�j�����&�&?��=t��>~3.?T)}>I!=ʽw7<W&����a�c�K�pܽ��佻)�<�`I��/<=�2⼅�> ſ۞�?A}�>:C�|b?}�����ڼ��C>-�L>fx���N�>
�,>*H�>��>��>*�->Rr�>�KD>cAӾ��>���b!�H&C�a~R���Ѿez>활�P&�����L���(I��a���d��j�L-���5=�sP�<�F�?ʽ����k���)�q�����?�a�>M6?�⌾�0��՝>���>�ύ>�@��8���#Ǎ��a᾿�?���?E~o>UB�>vm?�0?<񠾴�a��%9�ky\���:�j�N���k��$���猿�x�ڐ�pk\?�.^?�U?b{>S%f>��J?�p��AD�=��@>��#��9��ܐ=��>&����<q����о�����+=�[s?5��?DR!?R���"=���>o�J?��?��o?��9?	��>N�>�GR?!�=>J�>��?�6?��?��?�z�<�:�:=�5�1�r��Ӥ�";����gy=_D�=���=�;�;�r>�w�=�ƽ��
�өQ�
ԯ<V�	=^��=�̖=ɻ�= g=[|�>%�\?�u�>��>�06?�0�5�6�8�����,?@?>=�ӄ��捾)���%�u >�k?�[�?$UY?��g>�A���>�>&��>�'>�Z> ��>5e�z�@��z�=�V>N�> ޜ=��O��g���
�1��_��<�|>���>�Yg>l�&���<�&ž+9�.�~>B��]�$���Q��q��>M��*�����>��m?�E?8�q>�ж���纪g���,?V1?@]L?��??��=9rܾ��Z�(�����=>/�N>����ǻ�:���.�v����=��k��n���b>t�
��ݾ��m��vI�]��G5F=�@�(�L=��9Sվ������=�V>_*���0!��!�������I?;�k=���Q�R�M����V>hM�>$�>5�<��u���@�Ԭ���=f�>�8;>Hg��)h�G��]��I�>3@??�e?��{?�/]�]t�^�?���ľ���í@�^�-?���>%��>�N�>R{��������F�����}`��?j��>��	�5��߾��H�TW����>gg�>ܚ>�:?�8?y�O?�]�?�k?�[?��C>'�;(���&?g��?�]�=�F˽�@Y��9���D���>()?��F���>$?�?�5(?�O?_�?kd>���B�آ�>MЋ>�#X��Ԯ��d>�K?u��>yX?)�?��9>236�r����,��R�=!�>#�2?�$?s�?w�>���>E���T�=���>�c?�0�?�o?Z��=�??;2>��>���=K��>���>�?MXO?)�s?��J?���>���<�7���7���Es��O���;�jH<d�y="���3t��L����<��;	d���L��B��Z�D�� ����;@��>��s>QV���0>�ľA���>>nw��'�������E9���=ni|>w?7R�>@#�\�=���>��>����'?��?��?����h�a��:ھ÷F��T�>"�A?�|�=�Im��v���t�z�c=J�m?��^?��V�i���Gb`?gr^?���xL��;�׾q	Ҿ}o_?�`�>H9����>nx?��?qB%?Tː���a�a���lk������w�=k��>�)�º=��v>f�<?Z��>ur�>?��=P,߾��}�۸�H�?��w?ok�?��?{�>��g�̯տ���g��N�J?��>��7^?��a䲾�оO՛�`%��>����������^]��$tP��˔��D��B>F� ?_l�?~�?��f?�\�PV���l���P���|�G���6)�/8m��?2���l��Mp������˾���u*>\x�55����?s>?�����>`Ϟ�4� ��BW%>�댾���\�<D�����<>�%=~=v�Dd	�����?d��>��>�K?=Dg���2�1-�*���@	�&HP>dH}>�er>S��>{��m�C���ӽ;⳾�a��U��}f>mH[?2;F?OZi?�d�����{���=�Ȼ\�ɾD�p>u*>�0c>W)9��?u���2�&L�h���V�؊��{�q��=q�*?,��>�u�>�9�?J��>�����Ѿ���i�3�'~<���>�3x?���>Oh>Z_��a�8���>�&e?*�>�5�>�%��%n��x��6�0	�>R�>��G?�>�A���>��ʦ��މ���Q�b�_=
7`?�i��n簾%��=N�J?O�=8%>�[�>R����(	���޾{���]=Tv(?�=�=�>����,�4����¾�K)?�F?�ᒾ5�*��[~>�!"?�{�>)�>�*�?�#�>�Wþ�X�0�?��^?�:J?fPA?C�>?�= .��:Ƚt�&�g�,=5��>�Z>�Mm=�G�=F���~\��v��D=�κ=<μ:4��"><>̵�Z-I<��<��3>nIۿ�K��ؾ^������	��҉��������P(	��Zn����x�	�&�f�V���c��׋���j�xX�?��?�����ω������x��ֱ�����>4s�Z�w��>��H:�E���l:�O���Q!��wO���h�Ee�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >[C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@C|A?9�(����Q�W=��>�q	?p@>��0�s8�>����<�>�6�?(��?�6O={�W��
��ae?���;>G�� ��S�=�=�W=�k�x�J>�U�>9��{.A�u۽5U4>�>�#����jc^����<�]>JԽλ��1�?D_;���R�N�W��R�����>��j?�#�>:	>��F?��V�/�ɿ�x�>2�>�t @i.�?(	?��=�M�>Ь�@�=?_6?�ߣ>@F�斐��}k=lq�=*n�XU���1�[�<��=r\�>qk > 3=��_=��Y>�|��<��c�¿�L*��E'��5>���=��W 2����<�B׽{����OK�<��#��==<>�c>a�?>hL�>.,V>F�P?�1u?��>d��>b�+���a�8�ξE`��Q	�yc�.�Q��כ��?�hB��־�����>N��!=��=�6R�b���)� �]�b�S�F���.?�v$>g�ʾ��M�ˢ-<�pʾK���l݄�>᥽�-̾
�1�$"n�a͟?��A?������V�c��[W�����[�W?~P�����ꬾ���=������=�$�>	��=V�⾻ 3�o~S��s0?~\?9��8]��M5*>1� ���= �+?�?� Z<�)�>�J%?��*��&�nU[>8�3>�ѣ>Բ�>r	>���:I۽�?��T?
��V���d֐>qa����z��@a=O&>!-5�T���[>.*�<�����V���ּ<:%W?.��>��)�Y��n�����k8==��x?��?�(�>�xk?A�B?v��<�j��e�S� �$~w=��W?�+i?)�>ﻁ��о����5?G�e?�N>�Vh�>����.��L��'?.�n?�Q?y%���p}�������ee6?�
}?�Sb��C���"
�(��7��>Yr&?�z>w�'��;?ȋ?o<����w���Ŀ`c$�C��?G�@��?��%>�F�<��<6 �>H��>'�?�Ԝ;���.�J��ת=
U�>������H�I��9����@?�؀?���>����V���g��=�ؕ��Z�?\�?����Qg<D��ql�n��zk�<�ϫ=�
�QQ"������7���ƾ��
�\����࿼饆> Z@�S�O)�>LD8�6⿷SϿ����Zо�Rq���?f��>$�Ƚ������j�DPu�W�G���H�⥌���>� ==�	<NOž�d����3�
V=..?�7���>Tc���| ��3~�Ͳh��Q�>��>�B�>#׵<��%��i�?�d�lܿ�[��%�.���N?���?8�3?�%C?gM�>`4���o���H.>��!?b^?Q/�?�x]>�Mm�r��<%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�j�_?"�a�P�p���-��ƽ�ۡ>T�0�f\��L�����Xe�
���@y����?A^�?v�?���� #�d6%?��>���~8Ǿ!�<���>�(�>�)N>�D_���u>����:�h	>���?�~�?�j?핏�����U>��}?�*�>��?���=��(?{�/>��Ͼ���=Mk>�j5>��b�q��>�~a?s�?Ȧ>s�^7�m�-�,(B��,5��S<�|�>�*Y?�u;?�҂>�n��@D��d$�} 7=>S�0Oĺ���*5�<g�b��_>.G�=�N�=(��=��;��?Mp�9�ؿ j��#p'��54?0��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>=�>�I�>C�Խ����\�����7>1�B?Y��D��u�o�x�>���?
�@�ծ?ji���?�
�m*����y�_� �p���w}>��3?=W�K��>]r�>V?;�}_�����_�P1�>��?��?8-?��o?k�k�ƺZ���=�K�>� {?�?^~2��1Ѿ�N�>X�?%7����]7��R?%A@^	@n�X?f����ſ�t��á���-u��]�>� W�.�=�(�6�=����>��=d(>��X>�>'�>w�(>�� >kUN>�v�=��z�|�)�w����<���|�pt2��4�A���L�Q�˾�6����˾U�m��ox�e��� Kh��6G��/^=��=��\?��L?w�y?��?𛰽.�/>���o5�=���l�=�ǧ>�\<?,�L?�;?>L�<{ۡ��Q[��~��l��n�����>8C>��>Y�>���>kA3�7�d>o�;>8?�>{�>VW;=ڷ��.w=UDT>Zp�>6A�>���>�C<>Ց>?ϴ��1��l�h�w�X̽3�?s���U�J��1���9������ii�=;b.?|>���?пl����2H?���)�Ĺ+���>��0?�cW?%�>����T��9>����j�`>�+ �[l���)��%Q>il?��f>u>��3�le8�0�P��{���f|>06?�궾�F9�۾u���H�meݾ
GM>1¾>y"D��k����� ��si���{=x:?	�?B��5᰾T�u�qA���HR>h;\>�>=�l�=�XM>�\c���ƽH�Sd.={��=1�^>�??,>�N�=� �>uP��N�O�,¨>��>>�(>�d??	%?���>��O����.��{v>?��>�V�>ŝ>�EI��*�=�P�>j�d>,���������Ì=�MjU>� |���`�:!t�ԋv=z����_�=��=������;�;�,=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?-�E>��?81t?�I�>:��%C�҇��J���m$�=%>�����>#c#>|�ؾ�/����RǇ�N;k�9��/~\>�x=#�>��ʽ������=R]��K��yp����>+jZ>�oC>��>w�?���>�&�>���������J����:J?�&�?��E�Y＝4��j����)?�U?6=�
7��bj�>�kq?x8�?�^?oPC>.��u���Y�ӿ�7��6
�=X��=�.	?�m?(�[=�%�>��ҾW�/��(�>��>�@=�{�����_�軇�D>_�??�?9>�=*�?�O&?\'|>��>˻D����oJF�k��>(��>�v?�?JU?/�ľ��/���������QY�8Y>��x?6?3��>;�������Aa��w�U�������?�g?��޽�?~c�?��E?>8?�F>;�#�̦�-﷽G �>��!?����A�0\&�Œ��|?�L?�x�>zq��H�սԼ}��|�����?5\?,>&?��1a�þM��<��"��H��m�;��B�p�>BB>ӈ��<�=d�>Y��=��l��26��i<q��=�f�>@�=�'7�ێ��:,?}�G�@؃�Й�=3�r�ixD���>�2L>-����^?�=���{�����s����T����?���?�i�?}����h�~#=?��?�?�@�>�D��f�޾s��\w��x��e���>���>?m�x/�ۏ��i���6D��Cƽ[����>X�>{��>�?�8>cf�>�'Ծ C'�g�򾷍����X�R�-��-���#�H�	󛾿��~ٽI���G&l��t�>�nL�K[�>$M?�!>�l8>���>�t��`A�>�>�by>�<�>|-�=k$>fBk=~��<б��KR?�����'�g�达���T3B?�qd?\1�>pi�9��������?���?Ss�?�<v>h��,+�fn?j>�>F��Uq
?TT:=�5��;�<�U��^��3���4��>NE׽� :��M�Snf�rj
?�/?s����̾�;׽�?��!l9=�{�?��?0��ŰD�H x�JG��1\���7�ͳ��)���=�#�I�s��A��(.��j>��qL����=��.?5Ň?�,Ծ���;�d�4�F�(��>�>��>��>s�=K���A��[���!�ɮ_�c/�>��r?!�>bJ?r�;?hQ?�XL?o��>"��>g������>=�;��>���>P:?2.?�n/?��?;*?g(b>P����m���Nؾ��?ln?\�??U�?���?��9��sLS���w��!�^��=}�<,2ֽ�v���Y=�>Y>�X?���'�8�5���Hk>�7?g�>��>��q-����<��>�
?�F�> ��}r��b�7V�>��?k���=��)>���=����֪Һ
W�=���F�=6���};��<7��=���=��t��Y����:���;Nl�<���>P�4?�\�>�>�O������_P�!�=kb�=xq�:��> w��o栿�_��Br�5�:>�Ȅ?v��?_�$>.��=&i>`]���������Sא�YN����>"�W?�?&F�?��s?�A?$$�<���ގ��*���(��|�?\!,?���>J��[�ʾI�ˉ3���?S[?B<a����<;)���¾��Խ��>�[/�/~�m��AD�\~�����9}��ݛ�?ۿ�?�A���6�6x辥����[����C?� �>�X�>��>a�)� �g��%�P2;>���>�R?�>��O?�'{?�[?��T>a�8����������%�ٙ!>�@?�?���?2y?�I�>�1>*�o6྇Q�����e%��Ƃ�<�V=Z>륒>;��>p�>�,�=EȽ峰�t�>��*�=�xb>?��>���>c�>'rw>៰<�&L?�Z�>��ݾ%3���Ծ+
9����=�J\?ɘ�??D?(瞻�]#��0����п>䷫?��?��-?I@� �>��M���ྒྷ�]��>�>>�>�j�>����+Yx=�`@>���>�F�>T����Vg;�4�S=�V?�<?H��=�k����l���p�槾��=Ŗ��l{�X��t��� =>v��V�{�����E������~��$���ˇ���՞�>^�==�6>���=B���%-���8�7�=�����6}=�.Ž���<d��W�	��\Խ�~���6I<�S�=�H=�b��c~?I%F?*0?҈E?	Z>>��f��>~%��)?��>��=:����7<��k������UѾQ�׾��e�5k����>�$�ה>;[3>gr�=�զ<c]�=�0c=���=^��<�=F�="�=�N�=�P�=��=��F>��?�ŀ�ox����o�ߍl�U��?~�?�h�Ӈ���$�?�i���DZ��V�9���L?���?���?L��>:�<��>ҍ�E�=1s���Zs<�->��漪��<�I�>��=�:�5�n���uF�?���?��"?����b.���'M�`
4>��>�N���3���>�'^`��X�{�?x�:�f";�ۏ>c��=��羠�ľ��&=��3>aL=�9��"]��K�=˜~��"d=G�x=+��>�G>�G�=A*����=<�>=�1�=V�c>k޷:E�%���f���=���=��b>�>�^�>��?��0?%Yd?2ʹ>M�m�u�ξ�'��:ۊ>���=Ű>��=`x?>3o�>6H7?E{D?/�K?�߲>#��=�>�x�>�7,�-m�����g����<�~�?y̆?��>0�[<�@�ͧ���=�]ƽ�-?�11?�Q?Ae�>u�����a�t�-���h>�('�����Ҿ���Q�������= �>#Ϻ>a�>�>��	>��[>���>��>�!>��=�'�����<t��=T><<�Q��<�<��>�5�����Ĝ�;�-׽�.==,�!=��<�;|��!�h��=R�>
>���>��0>ù���CF>[L��B��eM=���;I���p�mWo�ٵ����y�I>��a>�T���Ί���>�(f>⵿=��?��v?&��=w���־򐿹�l=�|ܽE���z��=Ϫ��=�Q�g�҆U�B��m��>��>(�>=m>��+�]�>��rt=]��
5��4�>�q�����`��p�^L��#����:i�O�q��vD?)��*)�=�~?ԈI?�ݏ?��>����ٌؾ��/>���Lr=f���p��9���[?+�&?�2�>���s
E�iT߾IB�7�?oxl�$�;�Vz|�M�d��`k>����>�c��	v�xh#�����
�r�]|:���@�1��>�Q?0#�?8%w�ɭV���U��,=�,a�?l�y?@��>A�?�&�>�EZ�NH���՟����=>{?�j�?fʫ?��	>О�=W򴽊>�>�	?"?���?Kws?ҽ?�h�>�ǈ;�� >�Ƙ�@��=��>�r�=��=ui?��
?�
?�c����	�ݽ����^��<ώ�=�w�>W�>͍r>|��=�eh=˜�=M)\>6��>Jۏ>��d>��>�I�>>������'?���=ӥ�>��+?�Sr>����P��&2<�ļ�B��K� ������}�<*@���z=ҊW�U��>����]��?��>�"���?���W���$>Bf]>��f�>��F>Ƶv>�>i��>��>���>��7>FӾn~>����d!�+&C��R�7�Ѿtgz>Ԥ���&����w���|OI�5p���f��j�-���6=����<�F�?6����k�}�)�'����?S�>�6?�ጾ�숽ݢ>a��>Ǎ>4L��4����ō��a�@�?��?h�`>�E�>"7[?j�#?.�4�v.�8�>�h�[�q���/8D�"CA�گ�������־�d`��??�f?�7?k�5�>�o?�-�u�>�d�=��VZ�cf~>}֢>.�Ⱦ�?���������\j�<Z�E='�\?��? �?� ��5���>ũ=?�i?i!p?���>]�?���<�ot?�,>��?�W?~�S?��:?�(�>�&½a69=��r��E>
��D����yм�oL��F=k�>h�3��=w>�=!�;�6�z��>D�<T~�=tv��T��=�.>qxp> a�>k\?,��>���>�N8?6�K�6�$���C+?�=ʺ{�2#��\��4�����=��h?���?�6Y?=P\>�.@���=��  >���>��!>��\>�i�>V/�A��L=U�>L)%>�U�=SA�mS���{	������8�<��>U��>G�Q>�Kj�>
=v������ܥ�>��^��e���j���]�>�~&��D�>M�c?"�?�$>�톾��꽫�e���(?��0?��/?/X�?bo|=�e�C�L�8}E�Hӂ�'��><F�=��6�d���BE���CO���$����=3�;8����]d>2
��,ݾ��m���H������K=T�L=�
��Zվ`}��x�=�>�¾�u!��=��NŪ���I?A�f=�񥾱{V�����˜>�Й>Ϯ>Rp3�[&v���?�-+��LP�=���>�T;>����^�m�G��R�l�>3D?��x?�uj?yE��"�Q�);�5��&=���!�%?Jڜ>7�?&u�>^�ޢ���-��0x���O�9�?h��>0�I��$�)����� ����#�G>�(?§�>�?)2>?I=?�i?�?{��>��>j4�����0�'?�x�?�
7=j�˽c�^�4;�]5?�s��> +?_�R���>��?��?�.?�N?~r?޼�=���G���>��>@<[��C��'�d>�F?�j�>f�X?Vy�?+)>�6��[��1kٽ+��=�d->{2?��"?��?uv�>��>cG��-��=/	�>bvd?���?�Rn?�m�=��?�m/>pM�>�|�=�>�d�>$�?b�M?(�r?I!J?�v�>�a�<ˬ��D����}���T�V}�:�'<�ـ=;��Bh��
�k,�<.��;�ʼ� ~����p.�]_��(��:de�>�t>Vĕ���0>�;žN���I@>�S��si��R���B;�#��=�u~>�?ɕ>ɮ!���=�\�>N��>����!(?��?Z?Q�;�b�Ӈھ� K�\�>�B?���=4�l��]��:v���a=��m?
�^?��W�����f?��]?��޾�i����xz��ߜ���G9?80?W0���>{c?�Z?	�:?�)���Tw��ࣿ����A����	>Y�>i�[�4F�;a{>}`?6
�>�ּ>e�>�,�?�s��������>��?�,�?��?k�/>�]��̿����5���JT[?R��>넡�q!?Z����Ҿ{`��쫏����{���O��r�����?M'�,����ɽ}��=�a?�|v?��p?>�\?�q�$�i���[�
�{��S��8�����$�I���A���B�Mq�9?��U��fG��;�=�h��-�k�?�?�O	���?�
��}6�7�ʾ��=�w���m����=��m���~d4��ы��X��T�6�?���>�z�>�S-?ux\�	NH�����1�ܾ9De>\	�>�ʞ>���>='<�l�������Ҿ1z���Lͽ�/t>q�c?*M?��m?�p���,�%䂿���m5�����D>��>���>^�R�� ��('��o>��5s�*�:ˏ�|O
��}�=S�,?>݃>��>`Ֆ?��?p�	�(����r���.�T��<�}�>�g?��> �{>n�������>�m?�I�>{5�>5���Q���}��Vν�`�>�~�>���>l�f>y8&�T�X��؎�d��]�7��A�=��a?f-+a��^�>�E?�<�@A= F�>к?�գ!�E����G���>.
?u��=X�=>��ʾ(J�2*���s����(?7?�w���*�Իx>sJ"?u\�>	�>�*�?P�>I�ž�V�]?�m_?P�J?D�A?Z��>N =X	��tƽh�&�L'=�̈́>Z>�	~=_W�=W��ʞ[�����S=[:�=j�򼀒��q�<6��` <��<��7>��׿(�D�{�����
���оa�e����!���u��˽K*��+���b�(���d�� �g��rU�6}Q�A<ͽW�?��?)L\��|�󨿌,����־l��>�K�� ��=i������r�i��:��������fT�pvL�4g:�R�'?�����ǿ���:ܾ)! ?�A ?8�y?��9�"���8�8� >vB�<�+����뾬����οN�����^?���>��/��u��>ݥ�>�X>�Hq>����螾2�<��?1�-?��>�r�*�ɿ_����¤<���?0�@�|A?��(�����V=���>��	?��?>�Q1�]I�'����S�>�;�?^��?@�M=9�W���	��~e?�B<��F���ݻ*�=�@�=�8=\��]�J>�T�>Ձ��RA�@ܽ��4>�څ>F~"�P���^�^|�<�]>#�ս0:���g�?dhM�ʎg�2:N�ːr��-�<��M?ő ?�UG:��B?�^���Կ�W��7?�9�?���?z�+?ۣ/���>w�5�X?��I?�?UO!���{������>�G=�+�*�b���>���>�W�>���=I�:�q���;K���m�����Ŀje"�����'=Գ�:_���a1 �X�����k�	e��Cg��@ǽye=8��=�3H>��>.�Z>fci>�X?�Yp?d��>#�>�"�z���<j̾������U�ߌ��m8�DI�����.��I)�~�Ј�B߻�=��=7R������� ���b���F��.?-z$>��ʾ\�M���-<�oʾ�����ք�E襽0̾{�1��#n��̟?v�A?a�����V�4��F^�򁹽��W?vI�ļ��묾��=�ᱼ�=�&�>'��=��⾼3��|S�0?�?P��߀��8�&>��W�=
d+?j�?V�G<�q�>�%?-0��NܽJ�[>J�0>��>A��>��>!���Z�ս�?�T?�-��D�����>s���$v�u�k=��>{�8�S�׼�}U>�r�<k.���F��M��,��<�(W?��>��)���pa��'��7X==��x?��?.�>c{k?��B?Nդ<!h��~�S����aw=��W?#*i?~�>���i	о���I�5?�e?c�N>�bh���?�.�SU��$?�n?9_?0~��'w}����|���n6?��y?�h��[���?�
���T�>�6?�b�>��m�>�>�ƀ?Ꞿ�����iȿ�xV�K?�?�@#T@ %�<���:P�<���>��>����X����\7��d�H�n=�?��V���2��>䍾��@?Ho�?���>��ƾw�����=����aU�?��?͐��afg<���l�|b��~�<���=8��bb#�"����7���ƾb�
�P����㾼D��>}T@G��A�>B 8�R0⿧NϿ��0Cо�Oq�t�?���>N�ǽ˦����j�xju���G�
�H�4Ռ�u��>u�>P͏�)��sw}�b�@����z��>���O+�>
�M�����W���"�}�>�d�>��>
���2����қ?_C���οiß�X|�sV?���?7��?1?�e�<�j�͢��В0<��A?�l?��V?z�%���Z��S$�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�d�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*��+��<A?�2>���I�!�C0=�VҒ�¼
?V~0?{�f.���_?��a���p���-���ƽ5ݡ>��0�܂\���������\e�]��_dy����?�[�?��?ݥ���"��2%?��>����8Ǿ���<}�>�1�>�0N>�_��u>T�'�:���	>���?{�?k?���W���GX>2�}?V�>��?	�[��'?�C�=+M��΄=<h3>���>h��]~?�$Y?���>Zo�>��4=��<��M�dI���l�=�L:D>&�~?��8?���>��;�B��a���U��A����=�߳���>�@��.q�=&�>�(>)Z��s�����?D� ��[ؿL���?x�sS%?���>=??��(�+��<=�M?J}�>��&"�������?����?���?�h?-�龪����=���>��>PO\�5v½뉫��y?=�Y?�Q��훙�v�d����>V{�?'	@h�?_�}���?B� Ȓ�������p�>�2>?Xn��8�>_�8?9��<n�a��$������}�>��?�%�?'�>�<c?��k��A3��Ø=�'�>P*l?ґ�>ф��3� ۓ=�-?|�h���Q��\?	@�U@Wq?�3���cٿnȤ�����+r��1b >�'C>��?>�O|�_7�=E��=�J:�3�}YF>>�8F>�(:>!ɀ=v>�Cz>���%/��O���m����@�]&��5����
�?(����Ǡ���Eʾ<�1�1iɽ�^�;S�z�rv��6���v�=�+e?{�N?� c?�G%?��1�b���Ʊ�w>ZO��'">P��>��;?[#@?�8.?��Ƚ�Uƾ�R��K��sh��������>~�>i�>���>GN8>]M����S>���>�I�>�o=�w<LG9<|�=�_->卍>��?��>��<>�[>Q̴�3	��ߑh�*�w��ʽ��?�᜾/�J�	��b�������g�=�L.?7�>���vGпF��r�G?#���T���+��?>Ւ0?�,W?��>�[��c�V��v>�M��k�^� >����?�k��G)���Q>ɣ?'�j>�{>��4���6��lP�T����p~>�6?*<���/<��Ot�A�E�.߾ԕT>$��>����r��ϖ�q�~��7j�I��=�%:?�p?Qɰ�����2�w��ߠ��wV>�`>9='��=/
M>1�~�(M��%�H�`�0=e��=rhg>ȵ ?ok	>[��=;Η>�<����!�$�j>F�o>�^h<$�5?�:�>#7���5�������o�0C�>EM?`ߜ>]��=�;�,�=N��>G��>� ����9�5���g�LT^>h���us=�@����=�tE���=i��=Ύ����B�P�H=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�
�>�G4����������H���
�Q?�OX?�P��n>��սM��>m5?���[�������M^`����>��?�ơ?ɿy����-�f��4�>۶�?�&�?ܺ�>,�Ѡ��=��>�:?<V3?�Њ>�M"��>&�of,?�}�?iS?��H>V1�?�eu?W��>&k��+��)�����V�u=����}��>5�>�]��:�D������^����j��U��*\>~.=�>�۽V�����=�l���E���`i�x=�>�qs>�<K>�O�>8 ?*��>7��>?=mU������핾a>R?�Ð?86���F��F��R���]&���?�J?��:�>�����>�?1H�?��K??>�[&����&i���q�����=���=��>uQ�>:��}��=�@ھD�7<
��>	*A>hݎ=	'���������=B7�>��?$�?��>y� ?n�#?5Nk>G�>�RE� )����E�k��>��>2?��~?��?Q����43�����塿ţ[��M>w�x?�d?yЕ>����0n����R��jL�Y	����?Pyg?��� 
?�$�?�??��A?f>֛��ؾ�y�����>��?Z�s�����;�,~���?�Ű>C&>-������>��N���6���&?ff?��A?!�۾��<��C�NZ=�q��x��f'�<Y�Լ�Y>V�i>g+����=�Ғ>�+>��B��A���+���� �wL�>��W=��h�
�#>�+?[�-����F�=�q�;�B�Vyz>�H>�¾}r]?}rE��F|��Q��������V�ԍ?F�?�2�?W��~g�[R<?QӇ?�0?~��>J����&yھ*2l��z�F��y�>���>rM����;l���v��5����� m���?���>��?R��>��>�E[>����B!�G_
�gn�P�S��
���$�$-��S�M����fi�����[���]�����>�W=����>�k?(S>Z�>`D�>��*�]��>Qd>2�~>|7�>	42>%�>SM<ܳ��hڽmLR?���o�'����崰�
-B?iqd?�5�>j�h�=�������?���?�t�?$?v>�~h��.+��g?�/�>���q
?F':=���]�<�T��;��3��&��Q��>O׽�:�M�uf�k
?�.?�⍼��̾�׽�⚾�ݔ=*e�?h�#?�"��E�a�q�KXQ��HM��悽�oQ�]כ�T��e��&���D��b��-�-��<i-?f�?e����澖�ľ٧u��c.�6T>et�>�$�>���>��H>+����*�:�_��$�_������>Y�q?+�>��I?�)<?�kP?�M?"��>�Ʀ>-��0�>ô�;�+�>���>qq9?��-?��0?��?7�)?�~a>I�������Oؾ8�?|�?�z?��?� ?�����YŽ����v���y�����v~=���<�׽?�t��Y=��U>"V?���ޡ8�����Dk>�}7?ck�> ��>D��\��7/�<���>��
?�/�>) ��nr��R�HZ�>���?U��}�=V�)>���=G��h�Ǻ�;�=�0¼��=`a���;���<넿=K�=рw�K��@I�:�S�;�ۮ<��>!�?�b�>؞�>�'��������=�=&�O>|�U>,>��ھ����&���?�g��r}>��?��?�i=���=��=(���D@��P	�z���c��<�(?��"?S?�m�?�:<?��!?{%>������؂��ޡ���?n',?Cȑ>9���ʾ.稿��3���?X?	�`�+��'()��=¾w�ս`1>�3/��+~�X��nD�M���������"��?}��?��@�x�6�݂�����9����C?B�>��>	�>��)���g�:��$;>��>�R?���>�O?k5{?��[?�~U>�}8��#������L!�A!>�@?׳�?ގ?��x?S��>��>�I*�:�_���I�����ႂ�2�U=z_Z>���>���>,m�>���=�fƽ���s?��:�=\pb>�}�>�o�>+��>1x>�G�<'	F?�/�>K����>�Q���N=��̈́O�.�t?��?^�*?���;<���F����E��>�5�?�֫?C�*?�cD��K�=t�����J`q�q��>H��>���>_�W=��G=0$>E��>�w�>���:��0?�o{��N?�+B?�A�=�ſ'�q��Fo��Q��K�t<�ܑ��f�&����[��Z�=]���|U�7��2�[�u���Y��#����Z\{��<�>�T�=�2�=Ī�=���<��Ӽ�h�<(�H=q݅<(�=;{l�*Έ<)�7��jƻ���l�:���b<LGH=ڟ������J~?�S?��%?�	V? �I>a�d��j(= ��>d�	�.�?�W�>u׫=��v��/����۾���@��p=��S����y�Q>:��4?L>��r>�N�<��)����=\Й=e��<�<k��=Ť�=��=�ŉ=�=It�=��=,|?�À�༥�H߀�&��&L5?61�>)����X�if?j9>_J������s�<���I?�	@)��?5�!?X)�:�Q�>�f��3�;�g�=��"��=��+�r���c� ?ynY>�d�Ϛ��z"�v�?9�@J�??�z��u9ҿB�q>X*;>�x�=$dM�@.�y�W��S]��b�/!?�=���þ��u> }�=��徣�˾q9�<H�B>}�=	���X���=z&o���x=��r=Z��>�N>�=����
�=N�:=\,�=4�F>�ϻ�*B��V�Z�=�8�=�}^>] >�x�>��?��/?x�b?	%�>��e�I�Ͼ�ľI��>kv�=�0�>�|=34>Wi�>8?b�E?u�J?.�>�J�=҄�>I~�>�+�w�j�C��nڦ��q�< �?-��?�>�l�<��A��T�[�>�j3ѽT�?!1?F�?�S�>d���߿�=�������;�g���g<�.�P�	���=�bo��i=8U�>�C>�#�>�+>��V=Z`�=@%->�N�>�x>
��=�S�<6�T=��=����=>�׽�<���l=�r2>��={��=�dD<�D�oa.>FP=��< � >�?��l>�1?K��<@b��#"�����&�3��5[�W���i�9��U�� q�E8� o���v>ߓ0>�E�������>P�>�J'=���?��t?��˻ߝ��=�Ⱦٚ��ѽ�̫���>��P>K�L��)q��R����O�
�����>���>��>��l>,�"?�F�w=@��a5���>�{������'�9q��?������ i��EӺ��D?SF��ƚ�=�"~?��I?u�?Ȑ�>d��لؾ80>)J��=�=���%q�w_����?�'?��>��p�D�#	ܾ��½�:�>A0U�#�U�˛���G&��L��e=��w?�7���⾏��߂�r��J�9�{u�h��>uka?�i�?Q=�-���=[���N���� >?�,|?�>��+?�	?��h�m��>ʧ�V=���T?�#�?���?71>K^�=�U���1�>��?���?hӒ?ddq?�B1��w�>J�˺@>$	�����=�	>�4�=�l�=QD
?ʓ	?�
?0�� .	�f��A��4j\�Zi�<���=�G�>S�>)o>1`�=�`=�P�=�Z>���>ֲ�>@�r>x�>��>ǥ��y���'?DM�=��>!*3?��>G�Z=b.�����<�YE�Ţ?�D*�����\��<�0޻h>=�+ݼ~��>S;ǿ1@�?�WO>g��!?�[��(.�a[R>X5T>�۽r��>�E>K\~>��>kb�>_l>
�>u'>fӾ~�>�q�:I!��sC�JMS��CѾ�}z>	���BU �c9��l���F���������i�� ��w�<����<q��??���l��i*��d�k+?'V�>2�6?�?���킽��>>)�>��>Z�������@���m�Lŋ?���?48~>�F�>�wM?��"?�{�������\�z)]���G��d��3��ӝ��Clz���پ^���b�p?S�?8%?��=��2>6
v?��3?m��=��Xa(�{�G�ھ�>M�������䌾�\Ծ��R>�T�>ҐO?��&?[c�>W��J%��E>��??Sm
?{�?��`?��>��>feW?��=�Ͻ>V�P?��G?B��>��?ӹ��T�u�
��อ�^�=3<���"�\;	��E�5Z��.n�=��V>3��<,r=�������	�=���S>ʼpj�=��>>=< =R�=���>lL?���>��u>ʏ?(�罸�8�i$��,�?L�4�"��3����ھ .;>�>�o?� �?�N?�Ui>�K5�/w0��:$>��0>{�!>2��>]�>D1%�	['��+�=�t^>�"0>�B��U"�_ۇ��;�]٠����<�Z>��>/�n>�.|�^z�>�侺J`�u��=�6Ѽ'+�~FB���d�E�:� ��಍>��:?��C?���>�����RX>��G��
?C�#?�F{?De?	}/<�.޾a#�Ѹ,�pA��p�>�>�=?(���ũ�OS����Z�me>��/>|����ޠ�Xb>X��	v޾��n�yJ�����8M=��]V=_�U�վ�;���=�$
>����5� �����ժ��0J?8�j=]v���^U�wo����>���>�߮>i�:���v�h�@����d8�=y��>��:>�[�����X~G�&7�R+�>�RE?�\_?kf�?������r�2�B�����eH��V6ʼ��?(��>�`?�B>�f�=����>���d��G��>ׁ�>��!�G�K6��72��a�$��~�>a@?��>L�?��R?��
?s�`?�*?G5?�>�.��O��� B&?6��?��=��Խ�T�� 9�JF����>{�)?�B�ڹ�>O�?�?��&?
�Q?�?��>� ��C@��>�Y�>��W��b��=�_>��J?ؚ�>r=Y?�ԃ?x�=>\�5��颾�֩��U�=�>��2?6#?O�?���>�(�>�R�����=��>�fd?w�?]qn?�R�=C2?�!0>%�>(�=N��>Bw�>0?��M?%�r?�VJ?��>�|�<7����s����w�Y�P��u�;f.<�=�!�|�u�o]����<���;rʦ�Y����e�&�?�������;#w�>#�5>�p���SN=�׾�T˾��>�!n��.˾�ܐ��}��I:j9��>	?�>Qڽ�k5>�Ѷ>	�>��+��+?,	?"��>�ٌ=��O���R#��S<�>��9?�;>7�P��Ƥ�.������s?��I?*U6�紺��vn?�p?2.!�gZN��u�������þ�˄?W�"?��̾b�?�:�?�1�?NN$?˖��vp������y����#6�=0��>\�#�U�L�W�>�MF?��?��>"�8�q���v����8��>���?�i�?�?,H}>[ߏ�Ϝ�Q�G�˕���V?B��>�����X?�����r7��\~9�ײﾽә��Ծ+���4����*����YսU=*>Gc&?w��?�n?�R??y����k��<M�����e�(����Z&���o��L��"_���s�S���sپ#
I��v�>��yA��v�?�b'?i�/��v�>�Й�S��wL;��A>����������=px��-:==^=��h��~-��"��r�?ܹ�>���>ŧ<?�~[���=�'41��J7�����T3>L�>���>}.�>��B:��.�v齂�ɾ7�����ϽR1v>�xc?̏K?z�n?Rg��(1�W���ޗ!���/�Xh����B>m>c��>�W���;&��Y>�1�r�)���w��-�	���~=��2?-�>s��>�L�?|?>x	��o��2kx�;�1��σ<w.�>�i?c=�>��>Bн�� �T��>�l?�L�>L$�>�֊������|�қƽ���>��>)� ?��o>,3���[�Jf��Z]���R9���=g?Մ���a��~�>�rO?���;/*`<Y�>�|���������!'���>ZV?��=��<>+�ž���{�w݊�>�(??�7��8j*��H>�>"?�7�>��>��?���>�oþئ��$ ?��^?��I?�A?��>#=럮�>Ƚ��&�[�/= �><�Z>Q�p=���=@��d\��x��!D=b��=�μS���� <O���Y�S<(��<�3>�ܿ� L���־\ �r0�F�	�㳊���ƽ���[[��6���{��[*|�]M��?,� V���c�c9��"�g�/�?t�?5_����Κ�H����\���U�>a*w�Qi�S������[n������殾�j � �N��:g��5b�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >_C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾~1�<��?7�-?��>Ŏr�1�ɿc���}¤<���?0�@+}A?��(�]��TV=��>��	?��?>�O1��I������T�><�?���?rtM=�W���	�
e?�?<�F�r�ݻP�=<�=�^=L����J>AV�>0���SA��4ܽU�4>�ׅ>Q�"����*�^�m��<*�]>��ս!2��v,�?��x�����?�D��y���[>��f?p�>Rԉ��T,?|�U�¿h
�3�J?E�@�\�?�,?iƃ����=�:� b?�&?��>��x<���6�=��>��˽S�M�>�S����=�>�>�+?���RWS����˯�=��y��>ʿEe��f��ը=��<�ϯ�60���c���A�;X��viK�k8F����=[��=�->�k>RG>��J>�uU?�>j?5@�>4V>�F�� ���辎���ˮ�8��K豾)�,�Hي������p��������l�h���� =���=�6R�q���D� �w�b�L�F���.?sw$>Q�ʾ]�M�d�-<Spʾ,����ᄼS᥽(.̾�1��!n�X͟?��A?������V�x���V�����h�W?�O�����ꬾ���=������=�$�>���=���� 3�c~S��`0?5l?����@��,�)>� �	#= �+?3 ?+�]<Jܪ>�%?ճ*�����Z>��3>���>'�>�>v���ڽ��?��T?R��?���&(�>�T��|�z�nFd=)Q>��5��4�7�[>¢�<�茾�#M�0K�����<�(W?;��>��)��]a������Y==��x?��?8.�>\{k?��B?=դ<+h��f�S���cw=	�W?'*i?��>�����	оq���K�5?�e?:�N>ch����.�_U��$?�n?_?l}���v}�v������n6?Ty?f�h�Vo��*���������>�{?�J�>� 5�A �>�S6?4MQ�˻��b-Ŀ{�(���?�@���?�<��<���E�>���>�G�{kp����پa�M=�?i�����l�z�lG�%#4?�D�?�{�>�8���:�ҙ�=�֕�[�?N�?�~����g<W��zl��k��a��<]�= ���C"����3�7���ƾ�
�臭�Q޿�٧�>IY@ii�j'�>�I8� 6��QϿ���eVо�Jq��?���>P{Ƚљ��;�j��Pu�@�G�G�H�)�����>���=�ֈ�A���޶��O*D��r=���>�h�`�>��J��iǾ�����g��5��>7��>!��>��=K���r��?����3ֿ����p��k?F�?x?S�$? �>HO4�a/��d��=�t3?�m?��m?��'=��S����%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.���_?��a���p�~�-���ƽPݡ>��0��W\��Z������Xe� ��m>y��?_�?��?ܳ�w�"��2%?��>����"3Ǿ/�<�}�>!�>f*N>p_��u>����:�Xj	>��?��?ei?H��������\>y�}?��>��?P���:?�+>�T	�4>vIP>�R�<ʷc=��?&A?M�>��m>�p��=k=�R '�y���zT��8��6�>��j?��u?{wT>jeO�kd	>|<��*>^'ʽ�Ľ�~�� ������=�><?�=�c�=�""����;��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji���
?�I������d�������p�6Ǎ>*�7?���i�>FA�>� ��TL��6���X����>㒷?�y�?��>���?�F��l�j�ϼ1���Y>�?��,?�1˽i=ȾԿ�>�?��Y�j�����GW?��@�@��:?����w�ӿ�֘��2��3ۣ��v�=���=v<>�e:�=;p=%���阹{�=U��>[�[>H2O>�DE>��5>��>(܅�z)��.���쑿`�>�%d�������Ϊ��ge�U"�t�ؾU˹�gx罒u����'�b���3�� ��"��=�U�?��J?��?�-?N|C�go�>AR�-��=<���>��>��7?�jQ?[[�>z@ƽ�ü��.o���u�������y�>���<�>Rt�>�k0>��/�8[>wS}>`0�>��>6]�<��ɽg�=��>��>~V.?	��>�D<>~�>Jϴ��1��-�h��
w��̽\�?_���~�J��1���8������j�=b.?�z>���&?п����N2H?f���E)���+�E�>E�0?@cW?ߛ>�����T�&9>(��5�j�[^>�* ��~l��)��%Q>�k?: f>�hu>FB3���8�b�P�7԰� �{>2n5?C�����7���u��H�H޾��L>��>���ܽ�(����2~�֍i��{=wr:?�1?E���2��uv�ui���WO>ث\>��=S��=�N>�}f���˽�#G���/=��=_>@2?+>7�=$]�>Ͳ��[MB���>@�1>�h>�f=?֯?���.؛����/�,��?�>���>��>�>U�C�β=��>^�d>rz2�<�F�l���=���U>%��ˌG��Tf��(w=ۯ��aq�=iC�=h�����5��x%=_�~?�ƥ������[ٽl'>?5\?[��=�3�:9!����OL���4�?��@���?!��ddP��P?bΊ?'�ý���=���>p��>��ʾ��i�L�?�������4
��'��?kn�?@� ����)�j�yQ)>W"?V�;Qh�>wx��Z�������u�d�#=O��>�8H?�V����O�_>��v
?�?�^�੤���ȿ6|v����>W�?���?f�m��A���@����>:��?�gY?yoi>�g۾;`Z����>һ@?�R?�>�9�}�'���?�޶?կ�?'>g��?�Ƀ?���>��:=�B�\���A�u���=�Id����>��>�P�nO;�v\���S��h�u�����'>`[S==��>bЁ��Ӿ�m>f���7Y��-ө�ֳ>[$>��>���>l� ?'C�>��b>���8�QK�@>J�/2d��p[?p�?I�C�mvg�~�<�=l�U��'S?4��>�{h�w/3�d��>�U?�h`?Pe$?��=T.�&{����ݿeT����"��R,>L?S�?�����4=�
��Z¾���>(>ai�r�پԲྌ���c�>��B?��>���cF?��$?	�b>��t>�-�����\�e�>�	?��>[��?�m ?��ٽ2��%���Ѥ�����X�H>�g?l7?��>����Ҟ��`H;$��,>V�?D�}?���<\��>L�?��Q?��Y?�
�=�&.���޾��'���[>`l!?�[�'6A�rb&�A�-1?C�?�i�>�6����ӽ-���8�+���[?��[?�&?Q���u`�@����h�<�����(��O<7�K�h�>�&>:���Yݳ=�>H��=�m�V^6��X<��=��>��= 7��،�1�+?a>�Xb���ߗ=��r��,D�+0>l�J>c���i^?Ty=���{����J��2�T��?�u�?�X�?�h��hh��<?���?"?U�>�殾��޾��߾��v��x����z�>:*�>�9k����^���f���:����Žc�+����>���>n�?~��>h>Ӧq>�Ǌ����bI�Qg۾!�S�G&�'�4��W1�q�� d����&��E �p���x-���X�>��	���>R	?g�>�Y>~��>L$���π>{�t>㟈>ΐ�>]\>�>��g=����M~콏>R??����'�c%龘z���A?��d?:D�>9t��Z��zO�w~?$Ò?峜?fRz>��g��I*��S?��>1i��;a
?Y"A=�����<t�������򍽩����>�]ؽ�"9���L�	�g�:�	?��?�n��4̾�
ֽPʾd��<�?�?�2���>���}���Z��h@�y�ͽ$A �zč����/kl�����}U}�A���u�R�=2�/?޼�?!���,Ѿ�v��2 �mVV>�B�>�_�>��>��7>e*��6�/�x�c��(�z���a�?\G|?/8�>oI?��;?]P?ەL?J��>��>��p��>���;�'�>|N�>�_9?.?%0?.?�A+?պc>���.�����ؾk�?�v?NK?!*?C�?�؅��ýXl����h���y�`
��*��=���<�׽��u���U=>�S>��?�^�q8�]W����m>��7?8C�>G^�>�K���d���8�<2��>3�	?���>Cm���vr�mJ����>%��?�� =�R*>,��=��y���H����=̼��=uN��K>�L�G<j(�=���=�g��~�����4;OB4;���<���>;??�>Oϟ>s~��;j���	��i�<�3�=�2>�C>�������N'����a�ȶ>���?,`�?��%>$ �=�p�=�z��w�`��۾W����֓=i9
?-�?�6?B �?rRR?�<�>!YD>�$��Λ��;��(B~�X��>�!,?o��>����ʾu�ފ3�Y�?�[?�=a�	���=)�c�¾�Խ:�>[Q/�'+~���WD��������	p�����?���?_A��6�<u�#����e����C?-�>T[�>��>��)���g�q"��C;>���>�	R?��>(�O?�;{?��[?VmT>ԛ8�x.��Gҙ���2��!>�@?���?��?�y?fo�>]�>�)��S�����4'�uނ�>�V=aZ>���>� �>��>���=k�ǽ#0����>�T[�=y�b>S��>���>^�>��w>�ܯ<��G?���>ǳ�����a���N��8�A���t?g$�?�]+?-d	=���=�E�~t�����>��?�׫?�*?E�Q�4C�=`+м\;���sp���>Q�>�Ԙ>���=^5E=�>ݍ�>3J�>?��x%�]z8���L�f�?�E?l�=6ǿ7Mp��-N�D���x�;����$�q�%x���n���=���F|%�~e����{�>*��~q��JP�����r{P�� ?��=s�>�J�=���<>�(�RU�<~��=x������<�_�������&�g�B��YX��9=�c�=Li��(ɾ�kr?��H?�,?>O?Uf�>���=-���͌�>�$����?䈆>W����.��)�:����������Ͼ#LɾP^�ez��>��3�'>�d0>�(�=x��;�2�=�^d=!7'=cw-��=�ŵ={�=g��=m�=�U>��>1;�?�����ʤ��hd��	�R?M�?���O�Ǿd��?r�=������}�"J��;t?rc�?6_�?���>�ڽ)��>we��'#���=s��=|q>���K���J�>tX>
<����}lt�nx�?��@9�=?!l��TԿcb�=B~6>�)>ʚQ���1�`^��hb��3\��?.Z;��?ʾ��>���=�t�D�ƾ�+3=��<>�m=�O�#}Z�qD�=�p��&C=�v=�>PyF>U�=�!���L�=A�N=�M�=��K>罦�\�?�w%B�!�8=/��=�za>��'>�n�>��?�V0?�;d?��>$�m��6Ͼ�E��U�>3\�=���>m��=~JB>�A�>��7?8�D?��K?���>��=��>���>܁,�şm��[�����
�<4}�?�ǆ?���>�Z<�9A�9��Y>��tŽ!p?�;1?�X?�Ϟ>�|�e��r�%�,@.�~��/�9:p'=~�s�/$Q����� ���ὕ��=�}�>+��>V1�>�dx>\�9>�.N>Qk�>g�>cZ�<�Ê=�=���@�<���f8u=�Ϭ����<��ۼڋ��'��>�/��Բ�d��;���;��O<�A<0ґ=�>i��>��?�ѻ��N��z[</5�� @�5�U3B�a�-�z�|�ϜZ���F�M.#�}�>A4�>u&�9�Ո�Z�>^��>�
D=���?\�H?{c��ν�~vؽM���F�>`>��Ǽ
#�=��V�z~~�m��O�e�\6����>Kߎ>R
�>V�l>�	,�7?�	�w=�	�	`5���>�o��X��]=��7q�@��>����i�?�Һ%�D?�E��#��=L"~?�I?��?`��>@D��W�ؾ�K0>@R��T ="�u*q�Mo��`�?�	'?i��>@�O�D�&(��Vd�#�?�;����4�������)���/��~��ԯ>bNϾa8��"�&q����u��)1�S[�7*?�a?���?x�6�p�d��|=��(�E%�x�*?n
�?�Ò>}�>�`?�=)��㖾�3[�1߅>��I?���?[��?2��{��=1q��<[�>�?�*�?e�?�nf?P�A�}��>�M�}#&>�;���=2�!>���=#�=�"?�?$1?澘��t
��:��K?R�b=�.�=4܇>7>��i>���=��=��=�)P>��>���>�-d>��>��>�N����_-&?oc�=��s>p�&?}�g>��(=���֌m=V��h�s�6YF�k�սu Խ��=���<�Ě=.�<0D�>=�ÿ>�?�q�>pL��m?H5��M΄��Y-> �E>��z��>�sj>��a>�/�>��>;�>|ē>�95>z�Ҿ�(>��
��� �bSA�NQ���Ծ�y>솛��J-�Ċ���:�G�U����H��	j������<���<!�?���,Al�xs)����M?�ҩ>�a5?�u��.ꀽ�}><��>���>���:���}�����⾫
�?.��?�?4>��>�WE?s;?�D��v�ѽy�W�� Z�%V�~�(�fh��?{��aP`����e�Ľ�j�?zp?I<?U>o> OO?�I��{{�0>�6߾�4�����T8�>�?���8̽F��U��\F�c��=\?X^?�6�>�L?�.�ѽ.=y�{�?��=?DR�?�p?�*�>,����?���)�?HJ^?Wz>�s!?�M�>Q��z�=��>�L>%2�嚭�󝽕����
�F<�=��h=ֻ�=��<���<�2����;��<��-=N��<�~�;�Z�<�\%=�Rj>��:?��>�
�=�|�>x�ý܌0��Ѿ�v�>>���a��=ؾw)�Q��=�q�?}��?_�??���>xn�l���!m>S�?u<y�>��{>�	�:�:����=� >-��=�#�=�_T��\Ǿ�оT:U�tb�==U>K��> r.>9��Py���þ�� <�>�叾���a�<��Z�7@��=s�E��>�	q?��?�s>W��`�V���b��1?M�6?V�?e?���=����7@�٬%��I��>�>�%���;�z[���?���UھP'3��F>rƽ�A����d>��
�4�ݾ�m���I����� @=�g�$pI=Y��ģؾRLy����=�H	>���� ��C��8h��~�I?�uz=�ަ���S��:����>���>�6�>�7G��僽�>�r���qʛ=���>�C<>$��F;ﾐ$G�|���T>DG?��L?ήi?/te��n�q�e��S�0�ɾG���d�>Fx>� ?\I�>�#=�+��l��j"y�Ni:�b �>���>u�������c��8���"���d>�٫>��u=�~"?�;V?��>B�v?�?{\�>�o�>K�?����>&?g��?s�=�Խc�T�9��F����>�})?��B����>y�?۾?v�&?��Q?[�?��>�� �uC@����>*S�>�W��^��2�_>a�J?8��>�=Y?<Ճ?��=>��5�M䢾wꩽ�E�=>��2?�7#?'�?���>�B?#6�Z��:�H?��u?��?�<l?w�;��>� r>��8?�ͣ>uTѽ_�=,�>a�E?�w?;�r?�?��=6�9R�s�<��0=��=�_=Gܵ�7
"��,�����<KI`;�K(��7�!R�<������:�r��q�>�=s>������1>V�ľb܈�G�A>�馼����h��y�:��	�=ʜ�>�?�Ք>x�"�ʒ=��>�D�>D��WD(?s?��?�`;�Pb��#۾ jL��d�>W�A?���=�
m�,���˸u��h=o�m?�k^?��W�����O�b?��]?>h��=��þt�b����g�O??�
?&�G���>��~?f�q?U��>�e�*:n�)��Db���j�$Ѷ=Xr�>JX�P�d��?�>o�7?�N�>1�b>%�=fu۾�w��q��h?��?�?���?+*>��n�X4�p���œ���[?b��>�z��'�$?=�[�>K޾e�'ۄ�������춾_c���|��d�X�-�=b?�ˆ?5�g?�NT?������_�w�`�\X|��hC�K���^�S�K�*���:�c�e�Z��������{�M����P�8��?g�!?�+�ڗ�>mA��՗��;l62>����0�K�o��=R1w����<��=�8m���P�����q�?���>˹>�6?��W��!B�?y7�֥3���I>�ܞ>f��>ߥ�>��u<4a��]ݽ�Vؾ����@:�t>�c?��D?�Tk?�񽐭2��h��*q'��옽0)���u5>���=���>��'��"��%�+p<���t��]�,Y������]=6%5?�y�>Xޚ>!3�?R�>&N	�����@���&��O#<���>w�d?���>�e�>;���ٯ"�ٯ�>N�n?���>I*�>�i���c�/Py���>��>���>e��>�U>����V��c��&����1�B��=��j?Ԃ�w�r���>�wS?��<�Z=%��>��M���!����Ä
�d��=��	?�N�=ĺ=>�ƾz�F}�ʘ��L`+?�k?`�w��$�e��>�F&?���>��>Χ�?,�>ߧ��Rr��U?!�T?�C9?h�,?��>'�<�p0�=ҽT�/�=<��>���>%B�=ʲ�=���1���(����S�=��=!����2���=@���v=����W=>�ڿ�K���־)Y�Ȃ�'	��~�����V���+��+��ϋ���x�!�n�8��VT���a�7:����k��}�?���?2f��y��ly��툀�$0 ��z�>�m���������U��n�~���<� ��Q�W�i��f�iP?������ӿ������R?X�L?��?�����B��[�8�[��(�=�н1������oԿhW��p�;?�>�>ѕ��/L�=m��>�弲�>>���>�`"��~�I�>�W�>��B?�3/?'����:�<L��p�t��?2�@'�A?q)�EQ�EZa=|`�>h�	?B'B>��0����������>�%�?#��?��F=,W�L*��re?�.<�F�¡��r�=�k�=@1=C��D�J>�;�>T��xEA�T�ڽ�2>5��>:E'�v���]��J�<�+]>�`ֽ�ӕ�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=dO ��ǿw���#��"=3�g<���d����Ƚ��M��"��d�j�C���;�=ǿ=} U>i؇>=bR>U0_>K~U?zlq?r�>R�>�w彨^���Ҿ9�輭�}�34�N\���%�n2��/���Ᾰ����6��c;׮|�BM>�fB������E��/���P.���5?�>���U��}t;�����2FL>�r��g��"�9�⎿���?�?���9����1
��ܽ�x>L>o?�ԩ�ϱ.�����W�=/����J�����>G5d>�]��IG���f�J�1?~$?B8��:l��[�A>����(e;F,?_
? >a��> 8?�R׽̽r�A>R�	>f��>N�>]�<>8 ��pm�#�?T�X?�A���݇��h�>��������Ս=#I<>u�#�^N��\>��/=�e���-�<w>置���W? ��>b��y�!�Ĉ}�����;�d?�3?IG�>qN?nN(?%��<�`��5K�F ��R�=��a?�l?o��=%���)��.挾~O/?�Hv?�0>��B�vU������Ծo��>�\�?�8?��:�����W��2&$���0?�?w?3�^��&��2��J�S�}ͧ>PM�>5x�>e9�ɉ�>)�>?{��)��_����34����?�e@!X�?<c<R �z��=� ?@�>7�P���ž���t괾G�n=��>{駾�u��f��,�t�8?�-�?�'�>�,��� ��3�=.܈��4�?1�s?N���	�,=��$�7Fk�>���o\(<YO,���'�dʺ��Ծ�9�8���up�@y��	�F��z>f�@���g�>�=w��$ڿyο$r��첐�R�?D�*>-�a=(���N�E�k[��]��FZ�+T��KD�>��>�Ӕ�l����{�Eu;�y�����>H
���>!�S��$��������4<��>��>���>�?����3ƙ?d���Aο���#��\�X?i�?en�?To?Q�8<E�v�Ǝ{��j��(G?a�s?pZ?��%�zG]���7��f?�Y����`��6�z�N��#A>��7?�<�> e*��Ƈ=t�=�?�UO>�!*�g7ƿ|赿�
��Σ?і�?.Z�Ke�>B��?ڎ)?SY��ؚ��e�9��&�-�K?��>>h��ge%���5����6Q	?�@1?�Q��H�\�_?*�a�P�p���-���ƽ�ۡ>��0��e\� N�����Xe����@y����?N^�?h�?۵�� #�f6%?�>c����8Ǿ��<���>�(�>	*N>NH_���u>����:�i	>���?�~�?Nj?���� ����U>�}?�'�>��?e��=eb�>`��=�߰��u/��>#>n"�=�
>���?��M?�Y�>A��=��8�]"/�XKF�;CR�I!���C���>?�a?)L?�Rb>%���2��!�E�ͽ}R1����v!@���,�Ћ߽�K5>�=>�">��D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Qa~����7�v��=��7?�0��z>���>��=�nv�ݻ��W�s����>�B�?�{�?��>!�l?��o�N�B���1=7M�>͜k?�s?�Ro���j�B>��?#������L��f?
�
@~u@`�^?)	�ѿ� �н�^����"=��:щ=2��,6=���<�H�=�:��Yܣ=��>��>� >_	>m1>��3=�>���f�4�������}��K�d������������-+�e��r6������ʻJ(��J�ݾ�ΐ���v��=V?��C?H�i?�~�>�Q�#�S;�4%��n�O<�B�>�y�>��3?�x?w ?��μ`���-�b���������Z��KE�>hJ6>��>��>��>�:�<��N>�YH>i��>;�V>�̼�i<:Z�=zq>�C�>���>-��>�K=��= �Ͽ"��:Vg��@��E�=���?V;����k��x�������;��2�x{?*�>����Sӿ%���֔c?����S��~���%>>N]?�@a?�Ib>+$���8ͽm:>ŷ��hv)��P>1{ؽ����T�J�(�>C�G?Z�f>�,u>�3�1[8�t�P��{��V�{>S6?z򶾦`9�P�u��H��4ݾ�BM>X��>�D��l�p���a��[i��|=�c:?z�?���i2�u��I��(R>�[>=c��=�bM>6ab��yƽ�H�D.=ʘ�=n�^>?44><��=ţ>|���F8��M�>�C>�9E>�	D?�=$?��<m��S~��p/��m>���>}l�>�>y9H��̞=�A�>�j>iM�#�_�6��ک>��?F>?0^�;J��+��z=� ���D�=
��=U�߽�qA�x=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾOh�>zx��Z�������u���#=V��>�8H?�V����O�l>��v
?�?�^�੤���ȿ6|v����>W�?���?f�m��A���@����>9��?�gY?joi>�g۾2`Z����>ӻ@?�R?�>�9��'���?�޶?֯�?z:>�"�?J�r?���>����%.��嵿������B=�,$��T>:�=�ë�zH@�����oǄ�n|h�8�ƏQ>��@=g�>3�f1�����=��ƽS������ւ�>��Q>q8V>sǞ>a�?X��>���>gq�<J��������˓�P�K?��?q��B(n���<���=��^��?�=4?=*\�λϾ�ͨ>ռ\?nƀ?Z�Z?�S�>r���=���濿�x��<5�K>�5�>�E�>���eIK>��Ծ�6D�2s�>�ޗ>�p��*BھV��4砻c7�>�f!?��>{��=ݙ ?��#?��j>�(�>5aE��9��T�E����>��>I?�~?��?�Թ��Z3�����桿��[��;N>��x?V?Tʕ>X���ポ�iE�AI�F���X��?�tg?	S�4?.2�?��??l�A?v)f>��,ؾ�����>��!?����A�>M&����~?%O?C��>$��|�ս�7ּ=��3{����?'\?�?&?[���*a���¾'3�<�#���T����;�(D���>ۋ>툈�c��=�>�=�Om�DC6�8g<On�=H~�>�
�=w47�vw��R=,?��G��ۃ�x�=I�r��wD��>�IL>m����^?�k=���{�����x�� 	U�� �?��?ck�?�
���h��$=? �?(	?:"�>�J���}޾ה�nPw� ~x��w��>1��>��l�_�F���֙���F����Ž���s�>���>֭�>I��>�_>͝�>~@�G�>�M��?!��m�Vw��:�;�ٛB�;.9�OzӾ?:h�m���־�����n>��!=߄?�q%?ㆉ=5wh>��>ac�r�>���=r��>���>D	�>�.N>�V(>e�=�*���IR?����_�'�߸辿����-B?�rd?-�>'i��������N�?���?�p�?Hv>�~h��.+�m?.=�>E���p
?̴:=)�����<Z����ln���}����>�=׽k:��M�tif��e
?�-?�����̾�V׽6����.o=<M�?��(?�)��Q�8�o���W�dS�^���Oh�j~��S�$��p�ꏿ�Y���"��ަ(��A*=\�*?~�?���� ���(k�S?��Tf>���>o�>��>�iI>��	���1�v�]�I'�:Ń�?�>�Q{?Sv�>�@?�
8? H?!H?(�d>��z>n衾-��>�1*>�l�>�G�>��/?��-?��&?8j�>�M4?tke>/E��nV�d��O?��?�?չ?J�?'E��>/ӽ�!=���=�r�AQ�/J���8<+$Ƚ�U��^�.>�M�>�Z?-���8�c����
k>Ɂ7?�w�>���>s���,��[e�<$�>��
?�C�>����wr��X��W�>���?���S=��)>��=����3|ɺ�:�=Ij���ѐ=�����5;��^<C��=!�=r�s�pws����:��;yi�<��?�K??<~�>^@0>�p�3�B��p�>G�>�Ӗ>��>a0��>u��H����^�f��>'1�?"�?>\>ī>,�#>�>��U�������G�=� �>:�2?�h?��t?��?&� ?�\>-�\����܉�q\����?N$?b8�>�q��a��Q����'���-?^�?�"M�����q6�#�s��>�>'bF��.��ר���'����={?�d���tN�?�'�?
�x���G�����s���r;@�p?UT�>��>0��>����?���W�alw>��>ރ;?�Т>#P?@�`?�~R?�U>,S��꥿)!��[L�}=#3+?6Mp?t�?;��? ��>0U�=����������ӝ^�W����'�n�=�F'>D�.>_	?Ҩ�>1a?>M���-�;I��i< r>Ro�>~p�>�?*%�>~��=�G?���>_ν��5�
����ք��F��Eu?��?��+?+:=�z���F�R����h�>�Ũ?��?��*?�P����=\Ž�
]���w��+�>�ĸ> B�>g�=�a=�� >���>'��>�����2�7�'Mg�l�?��E?��=Ͻ��Wy�k�-�:���^��<�����e�;w�V���s�\���蘾�6ھ�6K��~��������e����1��Q�>˒	��\1>(�>"i=�fD�E�c�����<��>�����G=!V;���=�H��->��l>4n=�@�=�ʾ�.}?DI?M`+?�1D?|>N�>�1�P��>��h� �?fV>jC�j�����9��h��:7����׾4n־��d��u��=\	>RC�Ǌ>�02>��=�xa<��=�Yn=���=�<���=��=�=�4�=�n�=�&>�>�6w?X�������4Q��Z罦�:?�8�>b{�=��ƾp@?��>>�2������zb��-?���?�T�??�?;ti��d�>I���㎽�q�=I����=2>w��=u�2�R��>��J>���K��D����4�?��@��??�ዿϢϿ3a/>17>��>�R��|1��\�Rb���Z�`�!?OG;�&b̾G5�>Nl�=��޾
ƾ�P.=� 6>�!a=����D\�ɿ�=#|��;=�m=��>J�C>��=��N�=�J=���=�O>����Pc6���*�Uq4=$e�=l�b>��%>^��>T�?mE.?6�N??�>60���!��D��l��>D�>\�>��>hF�=��>�u?��{?��Y?q'�>��w>mj�>��?�A�tu����ܾx@ɾ �� ׌?"m�?]��>������g���-���\���(?�f=?�?�'s>�K�i��e��2*�}���<cǢ<B.r�Qs���� ���?Lɽxf�=�+�>*��>�^�>q�|>�e6>F�\>T��>D>J3=�}=k�<�c�<�i5�x��<��ἜU&=>;�c��<k��;˂ݼ�;�^�<+��<��6<=�u;���=�,�> \>�.�>h��=}��)�3>����^N��I�=`©�^�A�|c��}�>%1�N�@��s9>��P>n�����ы?PhZ>��B>���?A�u?�w><g �f�վ����s]Y�.c��Q�=Z�>�5�)�:�W'^��8M� Ѿ�y�>���>��>��3=��V�!I���*>��Ͼ@L���>iLϾ4�>Ig���UK�����3���{w���B"?���Xf�=�{?+K;?��?[7�>�Q;�k���YW���ݾ��>#�H�����l��S?Y?Yh ? ��˳>��H̾[���޷>�@I�0�O���K�0�0��Aͷ���>������оj$3��g��������B� Mr�I��>�O?��?y:b��W��>UO����(���q?�|g?4�>�J?�@?'&�� z�~r��w�=�n?ȳ�?O=�?}>L>k/��>4�?��?��?GNn?�@=�_��>ZT�<��i>0�n���m=U�>�M�=�g>;�?�U?k?R�� �	����ܾ��d�
�=#�f=��p>L��>j�O>�T�=�4�=Evb=	�/>Ib�>C��>�p>���>�Hy>��Ͼ'��:f?&�=��>��4?W�X>lV�=�-�3�)�=���Hx�ݍ6�)��{O但����$��=��E;0��>!N¿�p�?12P>#�;�?��� w�TmU>�j>Mdɽ���>��!>��>w�>��>��>(c�>��/>FӾ`>���Ve!��,C���R�7�Ѿ�z>圜��&�t�����AI��n��)f��
j�}.���<=���<H�?չ��/�k��)�����X�?]�>�6?bڌ�!��d�>o��>�ȍ>zH�������ȍ�?h���?��?;4c>[�>`�W?��?�}1�3�KuZ�{�u��!A� e��`��܍�E���
�
�L����_?@�x?�wA?�<>z>���?@�%�i���M!�>' /�2);���<=�<�>r#��:�`�óӾ�þ�S�.=F>�o?,#�?�T?�VV���/��\4>��6?3?��n?�'?*�'?��0��?�j>��	?w?5�$?f�+??f�>�G+>�)=�h�=do���l��������-�I;���=�= �>���C;�P4=-�=6������l�;`��ۃ=u��<��>r-*>�1�>:c^?���>w�y>S8?!�ʽ�7�.���<?a >��T�ؗ��,��$J����=�=W?L+�? N?k��>�1C���d�Er0>z��>�Q>|�_>�a�>����,t�-�=�K@>6�,>nf�=j�^���V� ���ms�Bm�8��=���>�0|>e���'>F|��1z��d>��Q��̺���S�|�G���1���v��Y�>��K?��?m��=�_龻,�� If�0)?�]<?�NM?��?��=*�۾��9���J�]>�=�>�\�<��������#����:��i�:��s>2��n�׾�Z>�%��A�پ�Ct�PD\�A�"���Q���[<��	�.�ľp�0�.%>O�>�þ�}"�z]��[�K?���=������y�˷׾TT�<ZЍ>�s�>�N�C횽�6�`{�����?��>Ƈ>�ɞ�����>�!=����>�HH?��]?u�?m�t�8�m��yH�A���ٟ��oȼ1�?���>%�
?[O>PA�=g���\��#c�_�K��>�N�>�����F��ǜ�������i8�>Y��>8'">=-?��T?�c?�Hd?	y-?�?I�>Ƹ�E�¾�B&?��?>�=I�Խ�T�'�8�8F����>"�)?]B�շ�>!q?4�?H�&?��Q?��?�>œ �+B@�B��>Cz�>f�W��k���_>�J?���>]>Y?�܃?�7>>�s5������R��-�=�>��2?69#?��?���>A�?k¾���c>u�3?Y�j?��w?��A?�Z�>�>�>;�1?¢�����8?��%?,)D?�
�?��L?jr>�M>=D���[�~�<<�/����<�I<OB/=����=�⁼/.彗���g��=�	,=5���'�a�l=R��;�_�>i�s>�	����0>��ľ�N����@>ۊ��BO��Iي�Q�:��ܷ=��>j�?���>�U#����=|��>kH�>h���6(?��?�?n�!;n�b���ھ)�K���>�	B?���=��l�Q�����u��h=�m?q�^?��W�m&����b?!�]?pg�=�t�þJ�b����~�O?��
?��G���>��~?�q?���>c�e��9n����Cb���j��ж=2r�>!X�.�d�2?�>m�7?�N�>��b>D"�=�t۾��w��p���?��?
�?���?�**>��n�;4�n��u��f�[?9x�>j���K� ?�5T�iZ��~�D�R��7���CZ��, ��쩓�6�D��h�L��ɨ=yo�>�Tu?��U?�h?p����y�(�d�3�t���C�	Z���<0A��O0���I��P�{t���@=۾��ɽiH�SKC�i_�?�'?V�0���>�혾���+k˾@qB><a��tD���=,V���Q;=�rf=��f��
0�a|��k�?胻>1
�>[l=?h�Y���>��m1��7�����?�1>�X�>_��>��>�rr��S,�{���/˾�
����۽+�s>Md?�9K?�Jm?G/���	0������N#��P5�ǜ��d�@>O>�]�>��P�n��Wr%�0>�5�r�������� ���y=��0? �>�ܝ>���?��?$�	����N�s�B�.�t��<I�>�i?���>���>��߽+�!�~1�>��l?7�>l�>+ڌ��!�(�{��$ʽ���>t��>]Z�>�o>��,���[��[��Г��9�> �=��h?�U��P�a���>��Q?� �9C�P<��>�Iz�-!�	�b�'� o
>!�?7�=�	;>��ľ����L{��K��|Y+?��?+j����&�H0�>�?���>^�>��?���>h�����<�?��L?�wB?!??t��>�Qt=����ڽ��>���u=�,�>l�h>$V=��=x����g�]�l�D�y<��>�kV<2ӽx�5=4z���%ż��"�I�#>�[�{�U�0<�����S�d�V�辔{��g�ľ�	��������Zʻ�0�=�]x=>9��U��@��xV��O��? &�?N�&�Pg���������z��l�> �¾u$C��⠾�ǩ=8�L¾�O���67�BB>���~� �u���3?ȑ���i�\ ���������>j�e?RD�?���.9��y9�.i}>�U6>�HĽ��⾙
���ɿ����_�h?���>���//��?��= e)>-^/>�N�������_>#�?��?h�!?q���޿�̴��g��Y�?��@�{A?�(�8��yV=5��>��	?w�?>�Q1�;F�^���|K�>_<�?���?�kM=��W�u�	��e?:|<��F�~�ݻp�=AJ�=�v=����J>U�>}�<QA�7ܽ��4>PӅ> �"����}^�P�<��]>��սjJ��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=s6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�8���ƿm^$��3��D=�ߺ��d�����߬��WY������gq�����Rq=�<�=!�Q>�k�>p�S>��X>ʯV?b�k?q��>�H>lK�N����ϾO�7��n������N�����He�5J߾�	�T�����v�ʾy^>��؏=��P�rK����!��zd��(G�tb-?�>��ʾPYM�;>Z<�Ⱦ�����n�����O;�3��n��ş?��A?�����W�����Z����X?6f���a�QN��*�=B�Ҽ���<�l�>M��=O��v2��	R���1?Q0-?hI��ۆ��S>t���
�����?	Y'?���=1�>�u0?b���#���v>��j>�Ǻ>-��>��C>[L��d�6�!m?��X?��ƽ� Z�ݤ>O�Y���c���~4>��u��Ŕ��g >��'=�Vh��Ox=�������zX?ө�>�!�� �N���7)����/=ݿm?�?br�>[�b?�k0?�3��u}�8J��r�$�=�T?��d?L�=N5���ɾ����=+7?Z?�>EZ��$��ʇ6��U�'j?�.c?��?�c!<pr�k1���$�w=?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�n���^�?t�?�i���jżn����`��f̾�ጽ��L�-��c3��v8!��<��ɝ��l	����*y��N>~�@�I���>g_�@)ڿp�ſ���G�߾�օ�1�+?(�>�\�+���O�c��5���Y�e:8�\殾a�m>��<>]��G�=7����_��V);��?Mt��}6r>`ţ�����0��Ib��m�>Ͱ�>���=�$t��]���ң?�侞�俱֭�#���6�?���?<�?6-?�H��ež�o��i�9L�=?�zo?�~??Y�^�S0Ͻ�n�<�Qf?�6Ͼ%���b�?�\�َN<�Q?#�?�U�q��=�	ɼ�d?d<�>ַE��߿���)l/�ԯ�?wx�?+��q�>�9�?O�D?�@��Ώ�]�T�N�"3ﻲ.J?9�6>Ż���hW���/�����
?*��>��ؽ׊�Y�_? �a�?�p�}�-��ƽ�ۡ>��0��e\�M��B���Xe����@y����?K^�?f�?���� #�h6%?�>n����8Ǿ��<���>�(�><*N>eG_���u>����:��h	>���?�~�?Nj?���������U>��}?�$�>$�?�t�=S^�>Mm�=��-�c#>�9�=��>��?}�M?	N�>T�=��8�a/�rXF�
FR�/#�`�C���>��a?R�L?�Hb>���T2�z!�]�ͽ?l1�r5��J@��z,��߽�+5>��=>�>��D��Ӿ�?*]�;�ؿ6g����'�b/4?^��>��?���6u�����1_?t�>>3�{(��{*���X����?�A�?�?��׾W�˼;�>nҭ>"V�>Q	սQ���W����7>t�B?���3����o����>C��?��@�̮?i��	?���P��Sa~���n7�L��=��7?�0��z>���>\�=�nv�ջ��Y�s����>�B�?�{�?��>�l?��o�0�B���1=1M�>̜k?�s?�Uo�f󾫲B>[�?	�������K��f?�
@}u@H�^?%��տ�]���Σ�����W>�5A>��@>����"n�=���▙��KN�G"�=�s�>��>즇>��>��J><�	>�����1�㹗�H����]4�	 ���&���������v��	�T�ɾ��I�˼�)3��}�����#ל�)؍��C�=�(T?��I?�Do?�o?�܋<L�κ���C=�BD��T>؆>ya ?�p-?�%?��W>O��p/q�.��Y�����I�>�l�>�O�>��>�.�>�/>]z�>Exc>Ȱ�>o'��q!�(0���i:2��>�M�>��"?`v?�L>�X2>�#���8��A]�XW��<}=��?�q���Y�������3��*��d��<��7?��B=!���� ̿wϣ���T?-+��a)I�{�P�6ؑ>F�C?tQs?��?>/��`�4��	>��[��7B�i:@>k������,�N��>p??��f>�u>ʛ3�se8�o�P�y|��j|>�36?�鶾6D9���u�ʲH��cݾ#HM>�ľ>�D�
l�w�����0vi���{=Mx:?ӄ?�6���ⰾx�u�lC���PR>�9\>�V=�i�=�XM>sbc���ƽqH��g.=_��=��^>�J?Ґ;>YP�=�Ҟ>�*���!I���>�)@>��?>C?}�#?�r
�g����-���K*��u}>C��>tw�>��>��I�hO�=���>��g>ڠ���!�����`E�Q>��h�b�3�9���=e��s >og�=���cB��?=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�n�>n��q䘿!↿��u�b�'=4W�>�DG?�9����t���2�/�	?�8?��'a��M(ɿ��u�5�>���?�6�?�on�lI��N�?����>���?��W?lMc>?m־��[�dZ�>>�B?;�R?�	�>������C
? ��?c�?��>yo�?��g?���>�<<�&��K��O���5ˀ=XȽ��>�>(�Ǿ�v>������w���Y��@���=���<F��>5ݽF�߾P��=\Q�:4N�����}�h>�i�>Eb>6��>��?�'?i��>&�T�#æ�t�p��ھZ�K?���?
���-n�w~�<-��=W�^��?�E4?�\���Ͼܨ>л\?���?O[?[g�>����?��s鿿�z����<��K>�7�>�I�>J��DIK>��Ծ�'D�m�>�З>�t��OFھ�2��8�IK�>�g!?��>cծ=@� ?�#?�j>�!�>�`E�C7����E����>d��>7@?��~?=�?�ع��Y3����衿�[��CN>�x?)S?\ĕ>����"����nF��.I������?�xg?���?�4�?Q�??�A?tf>���	�׾�����>��!?2� �A�M&���V~?P?���>�*����ս�Eּ;���~��i�?3(\?�A&?C���*a��¾�5�<��"���U�
F�;�eD��>��>7������=�>�ְ=�Lm��E6���f<�k�=�>���=Q/7��s��g=,?\]G�Dۃ��=��r�ewD���>.JL>���խ^?yj=���{�k��Jx��#	U�� �?���? k�?s����h� $=?��?8	?�"�>J��o~޾��ePw�1�x��w���>���>v�l�4�܏������F����ŽGYy�o�?W~�>"��>f��>��I>	��>�Mb�m�H�)��y-��ʒ{��b1���3�U�)�`�H���־�ǃ���%>v���7�"��)>���<�`>��?#�=p�b>l�?Y��Z��> ��>�'�>ә�>F)>aR�=���>N�>\�"��KR?�����'����Ų��h3B?�qd?M1�>Ji�9��������?���?Ps�?=v>h��,+�~n?�>�>>��Kq
?�T:=#7��;�<V��y���2����9��>lE׽� :��M�Mnf�wj
?�/?�����̾�;׽\kپ��=�K�?�? U;�\�q���z��W�?^��˭�Fe`��Y��H����`�C(��R9��}���B���x�yA1?�Ʉ?�v��1)�c���'�q��c-��_�>���>)�>@��>
��>ue�3�N��DO�J|(�㑟�S��>R{?-N�><B?yy3?�$G?'E?���>�U�>����S?cX=���>��?#$?ޕ?�)?��?�85?��U>��ս�u�G�ܾ��?�)? ?nL?�F?��w��]C�+�(�5�=������	�=�+=<K�����<֬�=0>�Q?}��8�"�����j>�}7?�w�>���>��u;��>�<�	�>��
?^>�>� ��r�Rb��[�>Ȣ�?����=��)>K��=��2&̺�J�=�l¼T#�=�1s;�!�"<.��=`��=T�v���"���:>*�;q�<� ?{�?�Y�>���>�6��]R ��D��D�=F�]>v4Y>j�>�tھbG��}ߗ���g�ðz>��?8g�?o�f=���=���=:���r ���z������Z�<Z?�,#?��S?�:�?��=?�"?n>�J�����T�������G?+�,?,�>�����ξ7���<�3��??۠b��W��S)�UR���{���2>�1�"����r�@��E<� ��ܜ���?խ�?"X����5�)��%��D⮾^'D?���>�:�>�j�>~�)���j������5>ѓ�>|bR?iW�>��`?Ag?� =?l.n>���G�������ൽ��\=�-!?+�?SB�?R�s?_%�>�5>w'[���$��B���̼+b�S�a�=�>�]>Ձ�>���>ؐ�>��=� �k�;ȸB��bS=ܠ>!�>PC?MZ�>P�=���@#K?��?�ޡ��Z�S��HJr���#���p?ܟ�?'�]?��h=��*��~7��|�	��>�ʡ?���?kW:?��M��x�=c��=3���{0¾}!�>뷴>�L�>�T�=��>��> ֿ>X�>��Y�����jD��D׽�H�>RJ*?�]>�ƿ�q��p��Ǘ�@c< ��me�ߔ�b
[��=ǘ� ��@�����[�8���4����ଡ଼���{�D��>p��=8��=m�=�l�<
wʼ��<&+K=�)�<y�=�/p��l<W%9��Jӻl������s`[<�RI=[����ʾF}?�I?��+?1�C?��z>��>q5�`�>�~��ud?�U>P N�����Ͱ:��n���M���aؾ�m׾��c�q��o�>��E���>�/3>��=(�<���=��r=�؎=����I&=+j�=�6�=/�=��=f�>Wy>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��6>�>��R��1�~^]�c"b��XZ�rw!?>4;���̾��>4��=7߾��ƾ�K*=�.4>Hj_=�:�j�[���=����;=G=h=5�>�_D>J��=;鱽��=E�F=���=�%R>3�G�S�5�D%.�X8=���=��b>)6%>�(�>��
?�k?�b?�ռ>]�:�;ؾV���%�>�*�>7-�>K����>,S�>:�@?hR?T?ā�>9(�;��>�T�>Œ�����ƒ��ݯ��+k=%�v?�<�?�w	?�|=\�]���)���2�����>��/?#t?T3�>�U����9Y&���.�$���"z4��+=�mr��QU�M���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=$�����<�vż���u&�:�+�0�����;w��;C�]<^��;�3�=y��>�h>���>BdZ=�a���^9>�����[�Sr>3ٸ� M�?r�u}�U6/��Mg�܄><D>����W���f
?K]7>T�@>�]�?N�}?��>3۰�.tо�@���
A��푾t�=AY>);ȽE:0��K��H��վ*��>BD&>Pp�>!�	>^�^��S�d�>���&:\��Z?��!�F�.;辞+v�;����˦�׌��Z�{=�_?� ���-W>�u?��2?�\�?v?����Ᾰ�>=��W�g���O�C��ƾ�,���\?��?Ē?�*��=]�Q}̾��*ŷ>��I�>P�Zϕ��0��*��Է��O�>�����nо�3�h��v䏿3�B��r�ڋ�>g�O?��?�Vb�_���O���rv��D�?��g?v��>�'?&?�퟽B�w��F�=��n?��?�)�?�Z>��=`Tx�~��>˨?e�?j1�?ǵa?�5��$�>����zV>�豽�@�=�A$>{��=S->k�?C�?u?���*8
��Jﾙ߾<�T��L?��q	>���>���>�W(>^�<(Pr<Q��=�W�>W��>sb�>��o>�&�>��>A��"&�l�	?$q>�=��<Ǯ5?�	/>���e.���t?��궽F��=���BԽ�'�����������>��=�/�>H�ӿJ�?y��>�c���X?��Ͼ򻁼4��>��>{}�*z�>��^>]9>q��>��L?J��>G&q= �;���� �4> �羭/%���Z�.���{��PIS>�鮾 ��C0����ڼ�Q���־���xdh��^����V�-�<�#t�?(dʽ��s�1E���?:X�>VtW?r��t�"�w=�%?�I`>�t�悿�h���bݾՇ?�	�?�;c>��>%�W?G�?�1��3��uZ� �u�3(A��e�#�`�t፿ٜ��ח
����6�_?	�x?yA?`O�<V:z>M��?��%��ӏ��)�>�/�';��?<=�+�>_)����`�P�Ӿ��þ8�"IF>G�o?*%�?xY?'TV���&�>�2?)9?T�m?��1?r�'?�Z��MY#?�1'>
�	?��>��6?�?��?�N�>,H>S<�˔:�M�񧙾�	�����$G��=V��=�߃=��A�@jQ=�^Z�X����^$=#�=������<5��=�.>�>�>��d?W#�>�Pd><i2?YK��3�=��=?xz�=L�y��?���������>��g?S��?V?+�w>(�A�XK�=">��>�%4>��X>�V�>����L�f�(<�Z�=,�F>���=Y�Z���f��t��띾�@!�x)>c��> +|>����'>�{�� /z�8�d>h�Q��ʺ�w�S�X�G���1�΄v�WW�>B�K?��?q��=-_��,���Hf�X1)?�\<?AOM?��?k�=?�۾��9���J�L@�T�>�M�<�������#���:����:>�s>E3���A����d>��
�4�ݾ�m���I����� @=�g�$pI=Y��ģؾRLy����=�H	>���� ��C��8h��~�I?�uz=�ަ���S��:����>���>�6�>�7G��僽�>�r���qʛ=���>�C<>$��F;ﾐ$G�|���T>DG?��L?ήi?/te��n�q�e��S�0�ɾG���d�>Fx>� ?\I�>�#=�+��l��j"y�Ni:�b �>���>u�������c��8���"���d>�٫>��u=�~"?�;V?��>B�v?�?{\�>�o�>K�?����>&?g��?s�=�Խc�T�9��F����>�})?��B����>y�?۾?v�&?��Q?[�?��>�� �uC@����>*S�>�W��^��2�_>a�J?8��>�=Y?<Ճ?��=>��5�M䢾wꩽ�E�=>��2?�7#?'�?���>�B?#6�Z��:�H?��u?��?�<l?w�;��>� r>��8?�ͣ>uTѽ_�=,�>a�E?�w?;�r?�?��=6�9R�s�<��0=��=�_=Gܵ�7
"��,�����<KI`;�K(��7�!R�<������:�r��q�>�=s>������1>V�ľb܈�G�A>�馼����h��y�:��	�=ʜ�>�?�Ք>x�"�ʒ=��>�D�>D��WD(?s?��?�`;�Pb��#۾ jL��d�>W�A?���=�
m�,���˸u��h=o�m?�k^?��W�����O�b?��]?>h��=��þt�b����g�O??�
?&�G���>��~?f�q?U��>�e�*:n�)��Db���j�$Ѷ=Xr�>JX�P�d��?�>o�7?�N�>1�b>%�=fu۾�w��q��h?��?�?���?+*>��n�X4�p���œ���[?b��>�z��'�$?=�[�>K޾e�'ۄ�������춾_c���|��d�X�-�=b?�ˆ?5�g?�NT?������_�w�`�\X|��hC�K���^�S�K�*���:�c�e�Z��������{�M����P�8��?g�!?�+�ڗ�>mA��՗��;l62>����0�K�o��=R1w����<��=�8m���P�����q�?���>˹>�6?��W��!B�?y7�֥3���I>�ܞ>f��>ߥ�>��u<4a��]ݽ�Vؾ����@:�t>�c?��D?�Tk?�񽐭2��h��*q'��옽0)���u5>���=���>��'��"��%�+p<���t��]�,Y������]=6%5?�y�>Xޚ>!3�?R�>&N	�����@���&��O#<���>w�d?���>�e�>;���ٯ"�ٯ�>N�n?���>I*�>�i���c�/Py���>��>���>e��>�U>����V��c��&����1�B��=��j?Ԃ�w�r���>�wS?��<�Z=%��>��M���!����Ä
�d��=��	?�N�=ĺ=>�ƾz�F}�ʘ��L`+?�k?`�w��$�e��>�F&?���>��>Χ�?,�>ߧ��Rr��U?!�T?�C9?h�,?��>'�<�p0�=ҽT�/�=<��>���>%B�=ʲ�=���1���(����S�=��=!����2���=@���v=����W=>�ڿ�K���־)Y�Ȃ�'	��~�����V���+��+��ϋ���x�!�n�8��VT���a�7:����k��}�?���?2f��y��ly��툀�$0 ��z�>�m���������U��n�~���<� ��Q�W�i��f�iP?������ӿ������R?X�L?��?�����B��[�8�[��(�=�н1������oԿhW��p�;?�>�>ѕ��/L�=m��>�弲�>>���>�`"��~�I�>�W�>��B?�3/?'����:�<L��p�t��?2�@'�A?q)�EQ�EZa=|`�>h�	?B'B>��0����������>�%�?#��?��F=,W�L*��re?�.<�F�¡��r�=�k�=@1=C��D�J>�;�>T��xEA�T�ڽ�2>5��>:E'�v���]��J�<�+]>�`ֽ�ӕ�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=dO ��ǿw���#��"=3�g<���d����Ƚ��M��"��d�j�C���;�=ǿ=} U>i؇>=bR>U0_>K~U?zlq?r�>R�>�w彨^���Ҿ9�輭�}�34�N\���%�n2��/���Ᾰ����6��c;׮|�BM>�fB������E��/���P.���5?�>���U��}t;�����2FL>�r��g��"�9�⎿���?�?���9����1
��ܽ�x>L>o?�ԩ�ϱ.�����W�=/����J�����>G5d>�]��IG���f�J�1?~$?B8��:l��[�A>����(e;F,?_
? >a��> 8?�R׽̽r�A>R�	>f��>N�>]�<>8 ��pm�#�?T�X?�A���݇��h�>��������Ս=#I<>u�#�^N��\>��/=�e���-�<w>置���W? ��>b��y�!�Ĉ}�����;�d?�3?IG�>qN?nN(?%��<�`��5K�F ��R�=��a?�l?o��=%���)��.挾~O/?�Hv?�0>��B�vU������Ծo��>�\�?�8?��:�����W��2&$���0?�?w?3�^��&��2��J�S�}ͧ>PM�>5x�>e9�ɉ�>)�>?{��)��_����34����?�e@!X�?<c<R �z��=� ?@�>7�P���ž���t괾G�n=��>{駾�u��f��,�t�8?�-�?�'�>�,��� ��3�=.܈��4�?1�s?N���	�,=��$�7Fk�>���o\(<YO,���'�dʺ��Ծ�9�8���up�@y��	�F��z>f�@���g�>�=w��$ڿyο$r��첐�R�?D�*>-�a=(���N�E�k[��]��FZ�+T��KD�>��>�Ӕ�l����{�Eu;�y�����>H
���>!�S��$��������4<��>��>���>�?����3ƙ?d���Aο���#��\�X?i�?en�?To?Q�8<E�v�Ǝ{��j��(G?a�s?pZ?��%�zG]���7��f?�Y����`��6�z�N��#A>��7?�<�> e*��Ƈ=t�=�?�UO>�!*�g7ƿ|赿�
��Σ?і�?.Z�Ke�>B��?ڎ)?SY��ؚ��e�9��&�-�K?��>>h��ge%���5����6Q	?�@1?�Q��H�\�_?*�a�P�p���-���ƽ�ۡ>��0��e\� N�����Xe����@y����?N^�?h�?۵�� #�f6%?�>c����8Ǿ��<���>�(�>	*N>NH_���u>����:�i	>���?�~�?Nj?���� ����U>�}?�'�>��?e��=eb�>`��=�߰��u/��>#>n"�=�
>���?��M?�Y�>A��=��8�]"/�XKF�;CR�I!���C���>?�a?)L?�Rb>%���2��!�E�ͽ}R1����v!@���,�Ћ߽�K5>�=>�">��D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Qa~����7�v��=��7?�0��z>���>��=�nv�ݻ��W�s����>�B�?�{�?��>!�l?��o�N�B���1=7M�>͜k?�s?�Ro���j�B>��?#������L��f?
�
@~u@`�^?)	�ѿ� �н�^����"=��:щ=2��,6=���<�H�=�:��Yܣ=��>��>� >_	>m1>��3=�>���f�4�������}��K�d������������-+�e��r6������ʻJ(��J�ݾ�ΐ���v��=V?��C?H�i?�~�>�Q�#�S;�4%��n�O<�B�>�y�>��3?�x?w ?��μ`���-�b���������Z��KE�>hJ6>��>��>��>�:�<��N>�YH>i��>;�V>�̼�i<:Z�=zq>�C�>���>-��>�K=��= �Ͽ"��:Vg��@��E�=���?V;����k��x�������;��2�x{?*�>����Sӿ%���֔c?����S��~���%>>N]?�@a?�Ib>+$���8ͽm:>ŷ��hv)��P>1{ؽ����T�J�(�>C�G?Z�f>�,u>�3�1[8�t�P��{��V�{>S6?z򶾦`9�P�u��H��4ݾ�BM>X��>�D��l�p���a��[i��|=�c:?z�?���i2�u��I��(R>�[>=c��=�bM>6ab��yƽ�H�D.=ʘ�=n�^>?44><��=ţ>|���F8��M�>�C>�9E>�	D?�=$?��<m��S~��p/��m>���>}l�>�>y9H��̞=�A�>�j>iM�#�_�6��ک>��?F>?0^�;J��+��z=� ���D�=
��=U�߽�qA�x=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾOh�>zx��Z�������u���#=V��>�8H?�V����O�l>��v
?�?�^�੤���ȿ6|v����>W�?���?f�m��A���@����>9��?�gY?joi>�g۾2`Z����>ӻ@?�R?�>�9��'���?�޶?֯�?z:>�"�?J�r?���>����%.��嵿������B=�,$��T>:�=�ë�zH@�����oǄ�n|h�8�ƏQ>��@=g�>3�f1�����=��ƽS������ւ�>��Q>q8V>sǞ>a�?X��>���>gq�<J��������˓�P�K?��?q��B(n���<���=��^��?�=4?=*\�λϾ�ͨ>ռ\?nƀ?Z�Z?�S�>r���=���濿�x��<5�K>�5�>�E�>���eIK>��Ծ�6D�2s�>�ޗ>�p��*BھV��4砻c7�>�f!?��>{��=ݙ ?��#?��j>�(�>5aE��9��T�E����>��>I?�~?��?�Թ��Z3�����桿��[��;N>��x?V?Tʕ>X���ポ�iE�AI�F���X��?�tg?	S�4?.2�?��??l�A?v)f>��,ؾ�����>��!?����A�>M&����~?%O?C��>$��|�ս�7ּ=��3{����?'\?�?&?[���*a���¾'3�<�#���T����;�(D���>ۋ>툈�c��=�>�=�Om�DC6�8g<On�=H~�>�
�=w47�vw��R=,?��G��ۃ�x�=I�r��wD��>�IL>m����^?�k=���{�����x�� 	U�� �?��?ck�?�
���h��$=? �?(	?:"�>�J���}޾ה�nPw� ~x��w��>1��>��l�_�F���֙���F����Ž���s�>���>֭�>I��>�_>͝�>~@�G�>�M��?!��m�Vw��:�;�ٛB�;.9�OzӾ?:h�m���־�����n>��!=߄?�q%?ㆉ=5wh>��>ac�r�>���=r��>���>D	�>�.N>�V(>e�=�*���IR?����_�'�߸辿����-B?�rd?-�>'i��������N�?���?�p�?Hv>�~h��.+�m?.=�>E���p
?̴:=)�����<Z����ln���}����>�=׽k:��M�tif��e
?�-?�����̾�V׽6����.o=<M�?��(?�)��Q�8�o���W�dS�^���Oh�j~��S�$��p�ꏿ�Y���"��ަ(��A*=\�*?~�?���� ���(k�S?��Tf>���>o�>��>�iI>��	���1�v�]�I'�:Ń�?�>�Q{?Sv�>�@?�
8? H?!H?(�d>��z>n衾-��>�1*>�l�>�G�>��/?��-?��&?8j�>�M4?tke>/E��nV�d��O?��?�?չ?J�?'E��>/ӽ�!=���=�r�AQ�/J���8<+$Ƚ�U��^�.>�M�>�Z?-���8�c����
k>Ɂ7?�w�>���>s���,��[e�<$�>��
?�C�>����wr��X��W�>���?���S=��)>��=����3|ɺ�:�=Ij���ѐ=�����5;��^<C��=!�=r�s�pws����:��;yi�<��?�K??<~�>^@0>�p�3�B��p�>G�>�Ӗ>��>a0��>u��H����^�f��>'1�?"�?>\>ī>,�#>�>��U�������G�=� �>:�2?�h?��t?��?&� ?�\>-�\����܉�q\����?N$?b8�>�q��a��Q����'���-?^�?�"M�����q6�#�s��>�>'bF��.��ר���'����={?�d���tN�?�'�?
�x���G�����s���r;@�p?UT�>��>0��>����?���W�alw>��>ރ;?�Т>#P?@�`?�~R?�U>,S��꥿)!��[L�}=#3+?6Mp?t�?;��? ��>0U�=����������ӝ^�W����'�n�=�F'>D�.>_	?Ҩ�>1a?>M���-�;I��i< r>Ro�>~p�>�?*%�>~��=�G?���>_ν��5�
����ք��F��Eu?��?��+?+:=�z���F�R����h�>�Ũ?��?��*?�P����=\Ž�
]���w��+�>�ĸ> B�>g�=�a=�� >���>'��>�����2�7�'Mg�l�?��E?��=Ͻ��Wy�k�-�:���^��<�����e�;w�V���s�\���蘾�6ھ�6K��~��������e����1��Q�>˒	��\1>(�>"i=�fD�E�c�����<��>�����G=!V;���=�H��->��l>4n=�@�=�ʾ�.}?DI?M`+?�1D?|>N�>�1�P��>��h� �?fV>jC�j�����9��h��:7����׾4n־��d��u��=\	>RC�Ǌ>�02>��=�xa<��=�Yn=���=�<���=��=�=�4�=�n�=�&>�>�6w?X�������4Q��Z罦�:?�8�>b{�=��ƾp@?��>>�2������zb��-?���?�T�??�?;ti��d�>I���㎽�q�=I����=2>w��=u�2�R��>��J>���K��D����4�?��@��??�ዿϢϿ3a/>17>��>�R��|1��\�Rb���Z�`�!?OG;�&b̾G5�>Nl�=��޾
ƾ�P.=� 6>�!a=����D\�ɿ�=#|��;=�m=��>J�C>��=��N�=�J=���=�O>����Pc6���*�Uq4=$e�=l�b>��%>^��>T�?mE.?6�N??�>60���!��D��l��>D�>\�>��>hF�=��>�u?��{?��Y?q'�>��w>mj�>��?�A�tu����ܾx@ɾ �� ׌?"m�?]��>������g���-���\���(?�f=?�?�'s>�K�i��e��2*�}���<cǢ<B.r�Qs���� ���?Lɽxf�=�+�>*��>�^�>q�|>�e6>F�\>T��>D>J3=�}=k�<�c�<�i5�x��<��ἜU&=>;�c��<k��;˂ݼ�;�^�<+��<��6<=�u;���=�,�> \>�.�>h��=}��)�3>����^N��I�=`©�^�A�|c��}�>%1�N�@��s9>��P>n�����ы?PhZ>��B>���?A�u?�w><g �f�վ����s]Y�.c��Q�=Z�>�5�)�:�W'^��8M� Ѿ�y�>���>��>��3=��V�!I���*>��Ͼ@L���>iLϾ4�>Ig���UK�����3���{w���B"?���Xf�=�{?+K;?��?[7�>�Q;�k���YW���ݾ��>#�H�����l��S?Y?Yh ? ��˳>��H̾[���޷>�@I�0�O���K�0�0��Aͷ���>������оj$3��g��������B� Mr�I��>�O?��?y:b��W��>UO����(���q?�|g?4�>�J?�@?'&�� z�~r��w�=�n?ȳ�?O=�?}>L>k/��>4�?��?��?GNn?�@=�_��>ZT�<��i>0�n���m=U�>�M�=�g>;�?�U?k?R�� �	����ܾ��d�
�=#�f=��p>L��>j�O>�T�=�4�=Evb=	�/>Ib�>C��>�p>���>�Hy>��Ͼ'��:f?&�=��>��4?W�X>lV�=�-�3�)�=���Hx�ݍ6�)��{O但����$��=��E;0��>!N¿�p�?12P>#�;�?��� w�TmU>�j>Mdɽ���>��!>��>w�>��>��>(c�>��/>FӾ`>���Ve!��,C���R�7�Ѿ�z>圜��&�t�����AI��n��)f��
j�}.���<=���<H�?չ��/�k��)�����X�?]�>�6?bڌ�!��d�>o��>�ȍ>zH�������ȍ�?h���?��?;4c>[�>`�W?��?�}1�3�KuZ�{�u��!A� e��`��܍�E���
�
�L����_?@�x?�wA?�<>z>���?@�%�i���M!�>' /�2);���<=�<�>r#��:�`�óӾ�þ�S�.=F>�o?,#�?�T?�VV���/��\4>��6?3?��n?�'?*�'?��0��?�j>��	?w?5�$?f�+??f�>�G+>�)=�h�=do���l��������-�I;���=�= �>���C;�P4=-�=6������l�;`��ۃ=u��<��>r-*>�1�>:c^?���>w�y>S8?!�ʽ�7�.���<?a >��T�ؗ��,��$J����=�=W?L+�? N?k��>�1C���d�Er0>z��>�Q>|�_>�a�>����,t�-�=�K@>6�,>nf�=j�^���V� ���ms�Bm�8��=���>�0|>e���'>F|��1z��d>��Q��̺���S�|�G���1���v��Y�>��K?��?m��=�_龻,�� If�0)?�]<?�NM?��?��=*�۾��9���J�]>�=�>�\�<��������#����:��i�:��s>2��MJ���k>z��C_ھ3o��JK��E��=+��b"=�e�K�־o.y��F�=�>tk����"���i2��X�H?�^�=����w�Z������}>8��>�}�>24�.����9�P��V�=���>Q$;>�����澹�F�߂���;>C~D?�u\?	�w?2�����{�]�R����Č��yc����>���>W?C�o>���=掗���\$g���Z�>��>sl?O��.'H�����j��@f����>���>�[^= u!?�??���>�i?�8?@ �>_U�>~���"���1?�i�?���=�a�%"*��E��zG�2�>ٖ^?0e���I>�	?�w!?T"?�1?�;??X�>���!��1�>N�>�	L�d����԰>1<]?��>��u?�8�?�	->�1�Rξ�8I��ţ>p~<CG?�� ?o��>��+>Q�?�7��>�>2l�>��?�x�?�O?���=r`?�x�>�K�><Q>��>O1
?��?}VZ?G�}?`<?���>�z�=[H���e;n���ƽ.Z�o�};i���-�2�J=��=���=R<"��6��#E=�ʉ����=�a�=j9>O�>۪s>1啾�.1>�ľ�8����@>&����R�������u:�6u�=���>��?�Ǖ>#��a�=2��>mS�>,��RC(?	�?�?�;��b���ھ�K�}!�>��A?q��=��l�fx����u��=g=F�m?�^?uW���P�b? �]?6h��=���þw�b����i�O?H�
?�G���>��~?f�q?`��>�e� :n�#���Cb��j�,Ѷ=Wr�>LX�Q�d��?�>x�7?�N�>F�b> %�=bu۾�w��q��h?��?�?���? +*>��n�X4�8���M��� fR?�'�>����2*-?�x�<ĝھJ���1��q�� ����羺K���Ǜ����X}g����[�=�n?��K?��k?<�i?�>¾� T���C�~p���N����,*�*T���1�~�O���D������Ѿ���B�潜A���PV��K�?�l+?"r�S+�>H'������Ҿi�>�{���S�Q��<�����=B�=�O�Oc��$�?�?{�>K2?��E���Q�3U@�ޣ6�ah�����\�>�a~>n/?�0�=)���\��VkľB����m��v>�{c?��K?ұn?���4-1������!���/��n���B>	G>��>:|W����b1&��N>�[�r�s��pj����	�\=w�2?��>��>�O�?�?y	�3f��/x�;�1�t�<�7�>�i?�9�>���>н`� �Զ�>Y�l?��>3�>���>]!���{�رʽ�"�>��>۹�>��o>
�,�-%\�uk��F����9�đ�=��h?G���>�`���>�R?C��:)rG<R�>N�v�-�!�'��#�'���>	w?L��=ߪ;>!wžG"�v�{�	<����2?�?6�t����]�>�3?A��>���>Pؓ?�F�>��O{��e;(?�$`??�<F?�#�>���;�89��`��i�`�d�f��߀>�k�>��E>-<>��#�t"�G�\>��>H.=�S%�A���I���Ւ�#�D<&�>�Vۿ�/K�Fپ������F
�'#������#y�����ݵ��?���x��{��8&�k�U�VEc��͌��vm�qe�?nC�?R���E��ݮ��ꡀ�������>/q�F|��x���|��ȕ�8ླ���Z!�7�O��i���e�t�!?�S���Qֿ����������>��7?_�?�B��]�"��0_<���]Tt��B۾-���Lѿ��6�1�K?^]�>�оQCN���>ne>�E�>���{��f�~�;�=l�>M�8?wy+?�Ք��5ݿQ�ʿ�q>���?ir@)}A?c�(�
��y V=���>A�	?��?>LN1�2E�-����T�>�;�?L��?@�M=u�W��	�=�e?�<��F�`�ݻU�=T>�=�F=<����J>�S�>݇��UA��=ܽ��4>&܅>�~"�%����^�>p�<��]>x�ս}1��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=D��D�ƿ��$��3���<in���HY�\�轂쪽��K�����o�����d=,�=&�Q>�G�>7~V>�IZ>KW?�pk?��>��>�"⽝�����;�t�҃����s>��'M�*���|����޾�������'�ʾ��-�
v�=W�����	�-��\��#���:?�c>�Q߾j�R�7����ƾ-N����=�Uv�$AԾ�I�5Eb�g*}?�'?5<��w�s���������P&^?axE��W�n����'G=0�޽�1��{�>><c� ��R7���P�}0?�S?^o���C��4�*>Bv �+=��+?'�?��`<�;�>�R%?�\*���㽾[>e�3>�>f��>l	>>��w۽�?�wT?�������3��>)���3�z�ӳ`=�K>b�4�&7��[>4��<����z`T�����$�<%)W?i��>��)�N�MX������E==}�x?��?�1�>�uk?%�B?�K�<�X��~�S�x� �w=q�W?�$i?E�>�����
о�����5?`�e?��N>�Nh�����.��R��?��n?x_?0ڝ��s}�]�����qg6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=����b\�?V��?{\���lD�����t��� ��y�<�_	�vt�����)�@�(�$���lG�����Oo��)�>��@Zm����>P�[�X�῞RϿ/���⽾J����?�/�>=�ռ` e�8]�[*m���@��A�/�P�>��>�ܔ������{�.p;�(���=!�>0����>��S�_'�� �����4<(��>���>���>�����⽾���?e���Aοs���E��>�X?f�?0p�?f?M�6<j�v��{�п�g"G?�s?�Z?��&��V]��98��U?�f��A�x���H�:�V�V��=?�> � ?��>�W���=��>/">�y^��Ͽ�3¿� ��j�?p�?�^ھ��> �?I?pO-�P8�� G�} Q�&Ә=�xf?��>=�n��L��� �� ����?Q�?~�3�[�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}??$�>��?�o�=�a�>dc�=i��-�Ck#>["�=��>��?��M?�K�>�W�=��8�~/�1[F��GR�r$�.�C�1�>��a?قL?jKb>���Q2��!��uͽ�c1�WN鼙W@�N�,�R�߽Q(5>��=>>`�D��Ӿc�?p��ؿj���q'�O54?ݸ�>:�?���t�����;_?{�>67�,��&���D�\��?�G�?��?b�׾�9̼<>��>�I�>
ս� ��􀇾��7>.�B?��yD����o�b�>d��?��@�ծ?ti��	?���P��Oa~���~7�[��=��7?�0�F�z>���>��=�nv�ػ��R�s����>�B�?�{�?��>"�l?��o�@�B��1=7M�>Ɯk?�s?�Ro���w�B>x�?*������L��f?�
@{u@P�^?*�����a|��ۥ����jeW=N+>,��>��s���=�M�9[�����1	>À>O��>���>�|>#��=:">œ��**��(�������q\�W�/�jr̾R'�����%�)%�����H�Ѿ�9Q�*�=uq��Y޾|!���K������-h?��r?tW?*��>Zݽ�0���)��8���Xz���=Q`/>K ?��e?�.?��7>(|׽�Jf��3���J,�0~�����>���>��>���>J��> �=��>��[>�>_@&>UJ=A�Z<��4>��|>��>7�>��>C�>�F�=�:�������gb��Q��-<>}��?�P���e�[Q���ѻ����3��jG?���=UG��4�ҿ\&����.?�v���s0�`4��"_�>�|?�9?�<>�j���'��>I>�R.�k��B$=�s;���Ծ��K����>x�?�~f>�Zu>�|3��R8��P�G���G�{>6?�඾ǋ9���u�u�H�vJݾ�{M>�>�XC��]�������Ii��|=�x:?Pm?ǖ��ΰ�Qu�O*��ER>\>�=U�=�EM>�b�K�ƽ��G�=�/=�g�=B�^>��?�n)>^�=�>����mAN���>p�>>�*>b@?}�$?J�J���(��;�)���y>���>���>��>��G��J�=���>�]a>���B���S�?�LY>�Kz��z]��|���y=z-�����=���=hr���n;��"+=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ3E�>`Y�^W������u���#=��>Y4H?AX����O��=�bx
?�?�U�7�����ȿwv�y��>��?v�?��m�;���@�cb�>d��?
\Y??i>�D۾�Z�2u�>5�@?�	R?!�>�9�Q�'�B�?"ݶ?k��?��G>�}�?'�s?�H�>�;��գ/�/��O���M~=g��:v�>�>6#��f�E�/���M���Jj���D^>��&=��>L�����Q�=]׋��M��0"d��t�>?|o>�GL>���>� ?�#�>�{�>�=����������}�K?���?b���,n�X�<溜=2�^��+??R4?42Z���Ͼ�Ȩ>��\?aÀ?�Z?Wj�>!��;��W濿�x��LP�<��K>�-�>�V�>�ƈ�aK>;�Ծ�9D�*o�>Uӗ>����2ھX+���ꤻ/@�>Ca!?��>���=� ?#?��j>�(�>.aE��9��^�E����>]��>�H?��~?��?GԹ�yZ3�����桿P�[��;N>��x?V?�ʕ>T���񃝿�fE�+AI�{���p��?�tg?bS��?2�?ŉ??��A?�(f>ԇ�<ؾ˩����>��!?��[�A�@M&�V��~?�P?���>f-����սGXּ����}��" ?�'\?�A&?���+a�K�¾�=�<��"�B
V���;YID���>Ӑ>K���=q>�ٰ=Om�MD6�8�f<i�=��>"�=V/7��x��0=,?ĿG�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>#�l���K���ڙ���F��_�Ž���H?/Ф>I��>�K�>~_D>��>�a�� D�.�������W����0��l$�< ��>)��4��e�V�V<�p���u&�g�`>;��G2�>�i?��o>���>���>[0��S3�> �i>;�>��>�>���=uJ*>~@�>�i;�KR?����#�'���辿���f3B?�qd?T1�>Ki�;��������?���?Ts�?=v>	h��,+��n?�>�>G��Vq
?qT:=9�W;�<V��s��3���1��>E׽� :��M�Bnf�vj
?�/?�����̾�;׽�ޠ���p=�3�?��(?��)���Q��o���W�S�����Tg��w��b�$�*vp�c⏿Y��^��_�(���*=�s*?�
�?�|�̫�E?��8�j�L?�x�e>�N�>3�>:о>��J>i�	�O{1���]��8'�����a�>n`{?9{�>��G?�<?|�N?-�N?Uޒ>n��>�款y��>�W�<K �>��>��8?�>0?�,?yD?�2/?��j>Zm��������ھE?�?<O?:�?36?M���;�佐���w:�߀������x=�e�<�cν�NX�S�Q=��T>�X?g����8�E���Wk>��7?��>���>���,���
�<��>H�
?G�>N ��}r��b��V�>|��?���?�=��)>���=?����Ӻ&Y�=�����=�6���x;�"s<Ɂ�=;��=�:t�����cN�:P��;�r�<u�>7�?���>�C�>�@��<� �d���e�=�Y>RS>y>�Eپ�}���$��e�g��]y>�w�?�z�?L�f=�=l��=	}���U�����P������<�?]J#?XT?S��?g�=?Sj#?�>+�bM���^�������?h ,?){�>J��j�ʾ3憎�3�;�?�b?�:a�����:)���¾L�Խ�k>�f/�V:~���|D�H1z�D��y[�����?���?�B���6����h���*I����C?R�>�`�>h�>��)���g�#��4;>���>TR?�>?�O?q|? \?��V>W�5��������T��Fq>�?? ;�?�T�?�y?��>� >G#����k���4��Uv��&���
}=��^>�>>��>	�>�3�=9���̾��D�9�2ߣ=o<a>��>/¦>���>�mw>p�=jH?���>����}��B"��g�C�7)v?��?��+?Ze�<����A����}��>O֧?q��?�)?��V�E��=�f�
Ϸ�s����>���>ą�>�z�=�<= .>���>d��>�6����{8�'M��?�FB?q)�=%Aſ��q���l�I����P<W捾��^��×���_��ϰ=m��H�����ۈ]�nҠ��U���������&w�M�>�n�=�+�=R��=ւ�<�/Ƽ�2�<��8=��<M=!����>r<���P�ܻ������;yue<�==����˾6�}?q0I?�+?�C?��y>t/>t�3�dY�>���K?qpU>��Q��j���s;�8���x����ؾ�׾?�c�q���`3>��I��>�o3>�M�=#�<�;�=��r=��=��M�PZ=�X�=�,�=�<�=m�=G�>�j>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�'>v�>4hQ��0�*�W���]�X�W��-!?��<��;g�>>S�=f�ྮ�ľ�=~a*>F�T=/��_�Y�b֙=��t�μ+=sK=���>��G>PL�=Z���G��=6uc=���=�_>T�'<�#���M�XJ(=�Y�=?�e>��1>��>� ?�E2?pxm?��>l3��,tƾ�Ͼ�C�>�=>�P�>h�?>R̔>�Zw>tu7?ZJ?�a?���>	G>M�>H2�>=C���Z�2�b��u ��/��?�ښ?JA�>�~��(5{���
��k,���S�=��>�?��>�R�>�U����0Y&���.�!����2��+=�mr��QU�����nm�/��u�=�p�>���>��>:Ty>	�9>��N>�>��>7�<�p�=�ߌ�f��<� ��W��=Ҟ��g�<=wż�����q&���+�㏦���;���;v�]<���;z�=��>��>�z�>|5�<�n¾�>q����*Y����=�&i���B���u�9y�6(� �e��Y	>�=>Nv�����?)W>��@>���?S�}?�R>��D���u ��CF�Ap���i�=N�O>0Dֽi"1�>=�zcW�Ա۾4��>�x>�qr>��->#^D���^����`9��1��v�>�v�����=�ǽ��u|�3����қ�$w�V_>�|>?�$���>�s�?ЕR?p��?\Խ>I˛=���)͓�ݕ�&��=�$��i��u'�=�=?�2?�7?��#��2O�}J̾����ݷ>RBI�^�O�����w�0�\��η���>����Q�о$3�8g������P�B�aMr�G�>A�O?�?4;b�iW��UO�����#��Iq?y{g?f�>�K?@?����v��p���o�= �n?���?=�?Q
>�t�=6�ǽ���>9b?}{�?&
�?�Lo?��@��+�>7A<p�!>�ރ��I�=�->�9�=�}�=�}?"?��?|���R�4q��G�n�Z��<=?<�=A��>���>o>R�=���=��=w�L>|�>��>{�a>?��>�:�>�w����K�>��M�=(%<?��r>����wͽ	^9>��=���=.�$��E=a��E"��vh�C�$>���>��>��ſ1��?Z�>U�$s?(vɾj|8���>�=�>������>�y�<H�>k��>��>��+>��t>^��= ,���9>�^
��M!��R9��EE���þ,>�񩾀�-�B�ؾ��צO�p����
��l�!�|��'8���q=��?Y��M,e��(*�����I?�|�>05(?�G�����3	>|d?X�>��⾮9���|���پ�e�?B�?R"c>��>l�W?'�?6�1�6-3��wZ��u�&A��e�}�`��ߍ�(����
�>�D�_?��x?EmA?��<�8z>W��?:�%��؏�A�>U$/�|*;��2<=�,�>B��O�`�šӾ}�þc��=F>،o?i!�??R?gV��5�n���,/?N�I?_u?�R4?[�?�]���?+;>�^�>��?�5?Ń2?>#?r�>.�.>�����ټ���<*t����\�w�>���7�=��!>�=Xq�Π3=N޼���=ļy��aC(�r^~=���=K9)>��V>�]�>��^?ݹ�>�ƅ>�8?�'�Z�6��ڦ��|3?p�Z=ჾ�"��ћ�����=��j?��?D�X?�m\>->���C��>�5�>٭8>�q>R�>��ڽ��F���=0�>��>u8�=!�5�4׃��c�����q�<\`>���>0|>���{�'>,|��m0z���d>z�Q�(̺���S�w�G���1�Ӄv��Y�>-�K?��?쟙=�^龂,��If�T0)?�]<?�NM?��?��=s�۾b�9���J�`>���>PS�<��������#����:���::�s>	2��%?����a>:�?Vܾ�gq�k�O��3��R�<�-��\e=T�	�Ï¾Q�{��6�=�x>{﻾f�!�Q◿S����N?}γ=������n���F��=�(�>�9�>:�N�1y��E����ꎝ=���>l�)>�0����=G��E��\y>�@?PJ?_E|?Q���`n��YM���+�2�����s�?q��>�,�>��>�sq=w��5
��"Y�iT����>N_�>�1 ��%�����S���#����>#��>Sh�>��+?�7F?��2?�,n?��C?&�?@t�>�̵���Ӿ.&?H4�?1��=�н��N�!�8�G�I�pL�>y2?1r4�攕>��?SB?�?�%O?�z?D0>�����9�P֕>���>��U�M���T>��E?��>BCW?��?��E>p�6�MӚ������=)>�(?� ?��?� �>A?��׾�=կ?��M?�?z�{?\U>F.�> P���?#b���=��"?(�%?�I?�?�
2?��\>��ǻ��7��摽��<宄=�DZ=�=ך�<Nf��Hvr�q-�������������<��=Ǎg=\r=N��:6]�>;�s>����0>��ľ�L����@>6%��S������[�:�|Է=���>&�?q��>�a#�|��=��>�C�>4���8(?x�?W?�}!;�b�� ۾W�K���>�B?���=�l�4���c�u��-h=��m?Ɖ^?��W�'*��N�b?��]?=h��=��þ}�b����c�O?;�
?7�G���>��~?f�q?V��>�e�*:n�*��Db��j�%Ѷ=]r�>KX�Q�d��?�>m�7?�N�>.�b>.%�=gu۾�w��q��h?��?�?���?+*>��n�Y4�"[ؾ�w����V?	P�>N|Ӿ5�*?���=c��h����'��kUԾ�/��ߦ�����Z�ɾ:�P��h��]��<Q>n�	?=|�?6[Y?zfh?�B���^�ܶR� n��d���>�$�vL���7���"�/�N�����")��۝�K���S�|�ݩE��T�?�B%?��5����>-Q���o��ɾ�?>'؛�ɻ��~��=�I���� =?�Q=�Dc��&"��4��F?��>�A�>��<?�Y���=��A/�h�8��)���N3>�י>�T�>�	�>���;�~*�O����Ͼ�7��>w�� v>�kc?�{K?�n?����>1�����z�!���0�ih���eC>Ǘ>9H�>�V�����%�AG>���r�"��P����	��t�=��2?2Q�>*��>/�?t?�3	�P��x��A1�'K�<�1�>�)i?�p�>L�>��н�� �:��>��k?M�>z�>������"���y���̽(�>Bo�>��>t�k>fa5��5]��܏��F��'�8�{S>�h?�{���wa��+�>PR?�$;'�~<���>��{�8�"�����+��X>\=?Q��=K;>��Ǿ����|�����$K*?#%?hjW�?S ���>f)?Xq�>��>�8�?;�>��;@7y�x"(?�N?�<?�:?|��>-v����;ҽ�\3��=���>��>U[>��6>�%޽d��nnN��k>�s�=e�j����Ὠ=S���E�F�����0)>�]�	�C��"��0���a��;��Ӂžt������{̽rؠ�؜�C{�IݽE	�=�	�n��H;컾2��?�%�?Mh��C��f��.���#�(��<�>�r�a޽�fվ�2��$Z]����t/������yT�`*g��Sb��^+?&�H�a�ῲ�����뽑��>@)?uȐ?�1��A�[�d��>�yH=�߇��ݽ�v��aݿ����yg?��>��ﾆ����>�m>(>�_.>@N�i-W����=�%?F	H?�?b�������V>�0�?V.@"UA?2)�Q_�W�T=�N�>9�	?�R@>�W1�2"��氾�I�>dP�?�ߊ?kM=(�W�#O
�_e?� <>�F���ԻSM�=��=!�=9����I>�Q�>P�p�A�0�۽�3>B��>��"�-P��6^��ͼ<�\>�ս����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=d��ʿ���-��1]<�Y����k����#L��9CH��K"'�n�����=�b#>2_Q>��>+#>%�>E�M?o]v?x�>D�>���Q��	�����Ԋ���K��������ۋ����澊���?���+\�xE ���ž#�K���=�!7�^��{�5��F��7Z��(?�K�= ݳ���X��U�=����m����3=�ؽlܾZ�J�l�z����?r�??nڑ��a����x������=Do�?�%�@����V$D=+l���Ы����>A��<�8��T�2��)��M0?�?6���NƏ�8�1>����ml=",?��?�6Z<�8�>�U$?(�!���߽e8]>��5>��>g��>|�
>�>��v����?�T?�5����l��>�����у���N=m\>��1����_�\>��<�匾Z�H�Xŋ���<�&W?���>�)����a���g�<�<=:�x?�?K�>�fk?�B?���<%g����S���R�w=��W?�$i?�>�����	о�y����5?��e?��N>�Gh���龉�.�eV��?-�n?�c?����'}}�������d6?��v?�r^�`s�������V�i<�>\�>���>��9��l�>֑>?�#��G������Y4��?g�@���?
�;<!���=�;?�\�>��O��>ƾ8y��׃��z�q=x#�>)���^ev���[Q,�.�8?���?.��>2���	��r8�=���K�?���?����s!i=�L�H_w���Yӎ�k��<�6���B��.�Ҿ��:���ݾ-����{��4���z>��@Wf�;/�>����ܿ��ο;����ɾ˚���?�?>;׽���i�I�+�i��FQ�cT�wH���a�>�>Q��r���"}��4@�� �9�>E�$���>C<q������q���#�:%��>�X�>#�{>���þ$�?�p󾪍п;����� �_qY?�j�?4�?��?�Y��y������0�I�[C?|�s?�LV?�}�U�a��Aȼ�m?`�j��2{��R���D��˾�D&?$��>�u(�Z�>D>)�q�>=��x��Hȿ�������j�?���?�0ʾq��>�e�?��R?�KN��ώ�E3V�>3�M�$=І�?RP>:���h�����5Ծ�%?}�=?�'d=P�D�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�!�>�?v��=�e�>?F�=�����'/�pP#>�	�=��>�o�?��M?fa�>;��=��8��/�WF�SGR��+���C���>��a?�~L?2ib>㸽�R2�!��@ͽ�_1��<��V@���,���߽�<5>7�=>�>E��Ӿ) ?�����ٿLt����!�k�/??�>E�?X��:�t�ӏ��f"b?�=�>�������܌�����?� �?#�?(�Ӿ�����7>�٠>��}>5�ܽa���ip�� NO>�B?|j�������n�+�u>˛�?8�@�?�e��	?���P��Va~����7�g��=��7?�0�#�z>���>��=�nv�޻��Y�s����>�B�?�{�?��>!�l?��o�L�B���1=3M�>̜k?�s?Ro���r�B>��?"������L��f?�
@~u@a�^?*T#߿pw��>��a����=���=�e�>������=�)B>	
>P��;�	�=pm�>X��>�v>�=>�"P>C��;f}��Ģ��R��6���xGB��O(����;��������v�E�F�Q\о�Yv�j��;�����n��ۀ�.K�'�=^�F?\�d?p�l?�Z?���(��A�=�����=ݡ>��T?�O?|{6?�<>�Z��*�x�,�����nۙ����>�bB>7�?�!?:ڊ>N�<bh�>=u>�o >8��=�q#�.j�>�=�Jy>�҈>0��>)��>��>��W>�ε������J[��2��~Rh�^ε?UF����H������!��>ݰ��V�<L=?v��=�����ֿ�]��v�]?�쌾��Q��ϝ��Q�>�}G?��?c�>סǾ�}$����=Yx[��у����=֕������%sQ���u>��(?��f>�u>˛3�ae8�o�P�i|��j|>�36?�鶾�D9���u���H��cݾJHM>�ľ>D�l�s�����!vi�͚{=Nx:?ׄ?'7���ⰾӰu��C���PR>V:\>�V=Qi�=�XM>bc��ƽ�H��g.=���=��^>�B?� +>#��=�ޣ>D���$O�4��>�B>�Q,>-�??"1%?s��O��t%���-�A&w>�d�>�#�>s>B�I���=F�>��a>.C�����mP��?��W>\'~���_��v��y=�e��H��=f��="� ���<���#=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�k�>�x��\����\�u��#=���>�9H?�W���O�#>��{
?I?�i򾑩����ȿ�}v�_��>��?"��?��m�h>���
@��v�>͟�?�bY?�^i>Ze۾�IZ����>�@??R?��>T@�<�'�(�?�߶?���?�C>,�?#j?%��>�-���(�
ͮ����+ƴ<˳����{>G��=�ľ�U9�x���������q�A�8�->��"=���>9�dצ�]��=�0X˾���ٲ�>{3i>UY�>{=�>�?�W�>�F�>5�=�U������ϭ���K?d��?}���(n���< ��=�^��*?V4?O�Z��Ͼ1ͨ>#�\?J��?[?�g�>���;���޿�Cz����<-�K>$B�>6I�>�ሽ�hK>B�Ծ-�D��[�>��>�����>ھ,��)���7�>�]!?�|�>�Ӯ=ۙ ?��#?��j>�(�>DaE��9��V�E����>բ�>�H?�~?��?�Թ��Z3�����桿��[�z;N>��x?V?rʕ>a����KkE�,BI�8���]��?�tg?uS�/?;2�?�??`�A?|)f>܇�)ؾ������>k�!?=���A�?L&���?�P?(��>v3����ս�!ּZ����� ?�(\?uA&?P���*a�S�¾�@�<Y�"�V���;��D���>��>����^��=�>�԰=?Qm�kF6���f<8j�=���>��=�,7�8w��J.?�t�:Moq��^8=�}��Q�[��>ߑ2>#�����}?Dc���v��y���x��� �����?q�?���?0�;��&e���/?���?i�?�i�>� ��܏����ݾ<c��u�H�W���>k1�>�e;n�׾%���y����!�����	H��P�>	),>���>���>��>�G�>�����;���ھ� Ǿ���0�8�3�<[���D�U�E��x��}��=_����|���>~4��;>X�?C�=�w>ٔ?�ǽ� �>�^�>T�c>�EO>�׎>��>{�O>��=���+KR?R����'��辈���C3B?/qd?�-�>�!i�3��������?ʅ�?�r�?�8v>�~h�-+�sn?s=�>���gr
?�O:= �@�<�W�����0;���C��>gD׽!:��M��kf��j
?�.?7���̾E׽x̠�Ao=�I�?7�(?��)�C�Q�n�o� �W��S�����*h�j4����$���p��ۏ�CT��+#��/�(�Y(=Y�*?��?΂����$1��u3k�M?��f>|��>+�>���>EeI>�	�o�1� �]�KR'��Ń�0!�>!<{?ʭ�>¢N?��7?R�C?�?Y?�˟>
u�>Yy��n?�W;v*�>�H�>M�C?"?�t,?��?9L*?��>�������^h?�?L� ?U?$;?	V���;��Pِ�=��=U�G�d�ϽW)�=�G=�m�0�R6�=fL2>?S��~I8�����J�i>�7?µ�>�k�>�ӏ���Q��<� �>E{
?��> �~Er�"���>���?\���e=2�*>��=R��H*�$��=��ͼ��=��}�eB��a!<JN�=i�=dd��Jӹ[����֓;i"�<�w�>��?>�<�>"M���� �C�� [�=FY>GPS>; >�Fپ�~��y%��6�g��Ry> u�?�{�?��f=-�=���=t���L��3����Y�<i�?GB#?]WT?��?�=?�e#?��>~(��M��I^��q��Ч?"#,?���>���L�ʾK�I�3�W�?.\?
:a����d>)�¾&�Խey>N`/��3~�����
D��U~�������J��?��?&�A��6�`t����BZ��6�C?s�>$X�>�>��)�~�g�F ��J;>���>�R?Ơ�>�tM?!!i?*�V?^}�=��E��)��)@��>玽���=�hJ?�w?���?��?��>p)'>I F�i�Ӿ-�����M}��J�/4m=��>�/�>Xo�>P5�>-|�=�"������#@>��p>�\?���>W��>�>�O���G?��>���$��΢����i����s?L�?:�*?�=x}�s@����pF�>��?!|�?'8)?�M���=`񴼋ѷ�^����Ŵ>��>���>W��=qj�=� >.�>}c�>W	��c��u8�J���p?}SE?�=��Ŀ3t�7l��)����<�A���y^�������X��y�=й��Yj�$��A�Z�*;���p��#䳾q=��Ut��c�>G�=���=���=���<��伪��<Nj*=�6P<��=�߉�EEw<s�6��Õ�!]���S���*;��O=ÛT��~˾=y}?dGI?/�+?��C?�z>��>24���>z��Q=?�:V>3�O��u���/;��v��
����ؾ5k׾��c�l؟� >c�H���>ˏ3>���=3�<g"�=�s=���=7�[�xy=,)�=��=^F�=QC�=L>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>R�7>�->��R���1�{�\�K~b��]Z�[�!?zI;��E̾�9�>���=2<߾7�ƾϻ-=�Y6>��b=mX��I\�Eڙ=QO{�43<=םk=���>�D>�3�=E6��n?�=�I=���=�O>P���qX8���+�]V4=���=�b>��%>XH�>|� ?�*B?��^?Xm�>I�#���/G��*��>���=�x�>�嬽p*�>�,�>!�.?�t?>X?��>ǃ=���> �>Q����~���������Q+�?�k�?�>6!���ٽ�T����[��-�C�?�n>?H�?\Q�>�c���࿌C&�tr.��ҙ�T_��Y�*=/�r�}5V��`�����F����=���>a9�>9ן>V7y>k%9>��M>�>�>�k�<��=T|��.ĭ<;)����=����~�<��ͼ�d&���7���,�����ٚ�;`\;�H<���;"�>���>"��=P��>r6�իѾ��>�w�	)g��v�>�&�ĳM��}�����t�U���ƣ=Rǀ>��S=�����z�>�F=磓>���?��?�Q?>+#�����]���`��(Z��~�>��>��.��Q���.�i�p��ǽ���>��>MΖ>�DY>�S/��]A���=I�ؾ�;�R?�̜�윽�M��Qu����蠿�e�va�<mE?�G��<��=?�m?1KK?p��?���>ܙ_�D/̾�X�=4͠�!�V=�Y���\������?E�?in�>���)�?��H̾7���ٷ>q?I���O�տ��H�0�y���η�.��>B���Z�о{&3��g��s�����B�"Fr����>1�O?��?Hb�U���UO��������n?�{g?i�>I?�A?�����t�v�����=J�n?���?�;�?h>�!�=�֪���>�D?{�?�Ԓ?6�i?-�G��y�>m����L>����[k�=��->r��=n�
>?R?�?	�}��`����V�-���e�*;��=���>�Հ>�V>��=[Z=���=\�j>g��>�ƚ>U�y>��>_�~>����p(���?���<�N	=1�H?���>�;�=;m�����H��=pI�f��9�3��c�������=DN>:�=���>4˿��?���=����?�������~Д>��>нj�<?�u�>�H�>���>���>vW�=�V�>E,)>�Ծ��>�~��u!�anC�"�R��Ҿtgy>�����%�����r�>KI�2~��f���i��!��O�=�r��<�b�?S9���k���*��:���D?M�>I�6?,㌾�����>~\�>̪�>s��U��0���|ᾏË?���?�3c>=�>��W?5�?yg1��2�@pZ���u��A�
 e�h�`��ߍ�♁�/�
��ؿ�J�_?��x?�mA?֑<Bz>���?U�%�ӏ���>'/�� ;��g<=�1�>�(����`��Ӿ��þ<:�:F>@�o?G$�?�S?}JV�A������=��J?%#=?ߓ�?��K?�?b�A��J#?��e>J�?�t?>�?Y� ?c�?� �>���=#����+�<��F�
J����g���Ō�FL�=4nU>���UW`�� <io.>+�"YU�6Z>�L��>=�d0>��->CZ�=���>[�v?<��>��>�O'?�,�݂P�{fW��w?��>wU���]��]�\��Ͼ�>s?��?R�D?�:o>d�|�5���_=|T>��w>$Q�>�H�>P���o޽�R�=��=�>o��=^��=�����H*��Ͼ"C���� >��>s0|>���޷'>|���0z�C�d> �Q�o̺���S���G���1�Ʉv��Y�>9�K?��?䝙=b_龼,��oIf�50)?�]<?�NM?��?�=��۾��9���J��>���>NX�<�������#����:��<�:��s>2��z����/b>�Y�z�޾�Wn�5�I�8羙pL=���%�T=�/�`Q־�o�����=��
>����V� �����ڪ���I?Cg=T�����T�Q����>�w�>ޚ�>R�8��sv��g@�yz���>�=
�>�):>������20G����>��>�8J?��Y?���?�;���si��G�e�b6�n����?���>��?�tA>6�p7��Ȣ&�NY�e�/�-��>�&�> 	��
r�L�̾?���$�ܣ>���>k�>'?eV?3?<�\?j�9?N�>��4>h�L���LP&?���?;��=o0Խ��U�In9�{8F��;�>Z�)?(�C��1�>��?5=?+�&?ׅQ?s?�
>�q��8@��4�>��>�gW�.���:`>�{J?_��>.Y?���?J|>>@�5��뢾�Ū�r��=!�>3?�\#?�?���>$k�>OD��}£=N �>�ed?E��?�'q?�$�=]��>��K>���>W0�=뺮>Y��>t�?P�G?{l?�H?��>\�<�������yU�Lճ��E^<��=�2}=&z� ��	��#��9>�;R �y�׼��~�k������uǼH\�>f�s>���	�0>��ľ�F����@>�Q��z\�����L�:��ݷ=��>��?䦕>N#��ڒ=���>�5�>����0(?��?R?��!;��b���ھ��K���>�	B?@��=C�l�=���@�u�Qh=��m?H�^?��W�4#���a?��d?�b��� ��.㾰�����eL?�)?������>�>�?��?3n?�L�6�k��d���'��"�T�@I�=�d�>G�
�ĺU��mp>��?��>�p�>�%>&~վ@pd���&�@�?2�?Hϳ?��?�#M>,ⁿ��̿mo!�.���
�K?A0�>��1�'?�#������.��ǔ��Lnվ�0¾���'���M�����0����!����=�?�mq?�da??D^?�(߾��R�9�a��\y�f�R�����+�}P��+���Q�8s� r	���־��[��=�&y�� @�^�?�a$?�3���>����
��qm;g$=>g��w8�T|=~|���lD=��O=�qh��I5��R����?��>q��>� >?DzX�i�;�B'0�5�8�����2$>�(�>��>�/�>���I6�x��l¾��u�נɽ�
z>X�c?�J?��n?}���
3��G��,���_���V���IH>^�>�E�>�^L���`l$�_m>�k�s�io��鑾��	����=qE3?fu�>N��>�?�T?|6	� ?xs�#~1�l��;��>ޡg? ��>*��>vǰ��E�Q.�>6u?��>��?,v_����4�o��pn�e��>��L=���>�Ä>MD��[G�N/w�݌x�e�/���1>��M?���Kl��ѩ>Pkz?�����<�%�>�j>�'�Tľ/��#��>�2?�]>��y<?�� J������R���H)?�E?�Ԓ�I�*�"H~>�%"?`��>(�>*�?�2�>`gþ��0�V�?��^?�@J?[LA?�>�>°=�����Ƚ&�&�52,=$��>�Z>�<m=��=F���m\�)��b�D=�!�=�μ�j����<� ��̺K<՚�<�3>��ۿ��J���ؾ~��_����@���B��uJ���F�y`��^���u������9���W�1�c�*֋�T�g�/�?3��?�P���ֆ��Q��?{��O� �vh�>�8p�ϱ���6��
|�t퓾
T�ۆ��?`!��O�Dh�Je�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >[C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾u1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@�nA?��'����RX=r��>�Z
?��?>��7�,�������c�>���?�^�?`tA=��W����)f?PRM<u�G��6лԒ�=z��=��=�r��J>n�>ݩ�6�B�?Aڽ%(7>}g�>�V#��f�v�\���<��`>8�ѽ<f��@��?(f��n�?�O������=ƨ~?�>1?e�>��X?m�y�~u̿�g4���d?��?��?�A?;���
?����\?�?���>C�Ѿ#a��ʐ��T�����')���9���A=��>��>��=�� �����eݻz�=���-*�����	=�.�=#&�=�w��O׽XB�{��A���� �����<���Te;<"�>��B>�p8>��>��]?��s?Կ�>��w>8J¼�T��� ��7�򃾒b��-˾U|@���`�S_�o���i���x�������#=�?:�=P4R�����7� �y�b�(�F���.?�g$>-�ʾ�M��+<vdʾ�ͪ� L���0���7̾;�1��n��ʟ?)�A?����V�� ��w�������W?>=���� ܬ�ܖ�=�ܲ�q^=A%�>���=���/3��lS�q0?�g?�d��!3��j*>t� �<=]�+?C�?sgU<%�>�=%?�+�,��b[>�z3>$��>���>��>t*���۽>�?��T?|��眾v�>L��R�z���a=�;>��4�gs�A�[>��<�Ԍ���]��䐽��<g(W?ɞ�>��)�+��_��:���3==��x?�?o)�>&yk?��B?���<�g��q�S�� �pxw=L�W?.(i?!�>Ň��'о*����5?e�e?��N>�`h�j����.��S�G&?��n?"^?�y��>u}�������fn6?/�w?�b�)1��G�����j�>���>d�>>�3�7]�>��:?�[(�r8������'4�uf�?�@�1�?�F\��!߼k=8��>Ԧ�>�p6����Y������u�=���>NǾ5mx�H�����u??�_�?�*?)Y��;����=�ؕ��Z�?7�?􄪾gg<���l�,n��nd�<��=�$��i"����{�7�7�ƾ �
�����?��{��>�Y@�]轇,�>i?8��4��RϿ6��b]о�Zq��?��>��ȽƝ��M�j��Ou�!�G���H��v�>�,>/����Y��%|�%<��%����>����-�>�eQ�%޵�5H��� <�ɑ>D�>��>#���ԣ��(ݙ?�E���IοZ���sE���X?By�?o5�?�I?��B<�u�`�{�-����F?9Es?t�Y?�I�d�Z��:�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�nc?L�z���p�к9���T��ۇ>��v�C��.�=���m�t��}��2�h��?g/�?!�?���(��<?�a�>x���X&ȾZ~2=uA�>wW�>��>X�i��>���}7�A��=��?Xc�?�Q?�덿�V����>��y?&˶>AЄ?��=�6?��=����s���Y�>�A>�+���1 ?�mN?���>hm�=MA���)��WH�ȭQ�c� �2�A�ṁ>=�_?M�N?+ya>T	̽��'��Q��N�����'W����3�u����s����>�)4>n�
>�W��yξ�?hp�?�ؿj���r'��44?⸃>[�?�����t�m���;_?~y�>!7��+���%���A�]��?�G�?m�?a�׾K^̼�
>v�>�J�>��Խ����4�����7>��B?��yD��m�o���>���?�@�ծ?�i���?� ������i��W�A������=�tB?#���zA�>��?�o=�}�6���9v���>�>�?���?�H�>�>h?���0C�����m�>M�?"r$?ԡG�pR��#�M>�7Q>D��h$q�����v=o?y��?Y:@��q?>��Y�ؿK���fw��+1ʾ<��=��(>1A>��1�=a>i��=j<���=�\~>`�S>E*>�y>�f�=Q�=� �����֖�5����3�A�����X�J�J+	� ���"�\�ffԾ�����.��o���^���(������>�8O?�[?Իp?���>��$�_I>����	�=I꾽��M>U�>�]9?C9H?�3?�	�=�Ȳ�uu]��Os�!���ܗ����>��)>:�?��>��>4�C�1Ŷ=�ҙ>�v>�=Wx�����bǄ<�H%>�J�>��?��>�C<>��>&ϴ��1��Q�h��
w�c̽�?����@�J��1���9������h�=Eb.?�{>���?пk���}2H?v���?)��+���>n�0?�cW?/�>���6�T��9>��ڦj�`>�+ �;l���)�*%Q>Xl?��q>�Cc>9_Ծ.�L��.�H\��Z�>(9	?Y�ݾ�:��%i���K�W�,�$�=���>������1��0���b�k��,�ЦO?y�>��ڽ�@W��>B��x�E�n>1XF>�ϓ��p=�Y�=�����K���w���ރ=�:>�Q?u,>�#�=�ģ>zV���P�-t�>�;B>�+>��??%?�V������~��,�-���v>O#�>EՀ>��>1^J����=J��>`�a>Eg�J���Ñ�x�?��}W>a�}�{_��t�Yy=�X��&�=D�=�� �W=���%=&�~?/��刿P�#���CgD?!.?*�=��F<�"����P����?G�@�p�?'x	�O�V��?B�?���JA�=�w�>J�>��;}�L�٢?�}ƽe㢾��	�\#��R�?��?&�/��ǋ�>l�B>^%?��Ӿj�>�|�.[�������u��E#=ߣ�>C<H?Q���O�K�=�ku
?p?�a������ȿ�xv����>�?d��?R�m�`B���@�r�>��?�iY?>ei>�d۾ZZ�T��>��@?ER?��>�6��'��?�߶?�?S|R>��?�h?ֱ?�+:�����/��R���Pn>�夽�>�??>1���Hn2��ߒ�f����yl�k���~>�_p=(�>�G3��hȾ^�M=���CJ���<漦ə>ب�>7�>�i�>	�?�>��Z>������Hr�jҭ���J?CĎ?BD��B�O��c�퟽O2����	?��C?�������ى�>3�q?�?��Y?T��>�Y������ö��ȹ������r>u<?�j�>5R���w>
��ЁN���>\߈>��ɽ�r��+D�G� =!(�>&n+?�\?=�=��!?=�'?�=�>���>�@�����I���>4p�>�U?��?��?�B���v#�b
���Q���d���">h�i?+?���>h���`a���F�������ǽʑ�?Z�c?��4?�B�?Q�R?C4E?�C�>��43޾_.��,p>��?Ea���;��Q(�&���^?J�?���>�o���սR#�3w�9V���?�[?#]#?����c�/�ξ"l�<E��QG�<�.<49~��N">]�>�s�����=P>�%�=��k��t=�ʍT<��=n�>�#�=��4��#��@=,?��F�Pۃ�R��=��r�uvD�B�>T8L>���^?t=���{�����w���U�1��?ӡ�?�k�?���[�h��"=?��?.?V�>jM��7޾���9w�5{x�9u�
�>���>ʆl��徱�������E��<�Ž���x�>]��>/�?�E�>��L>��>�o���C'��)�� ��]�Le���5��h)����FȞ��-��+s���þ�$����>=}��7��>�?~�m>�v�>���>��;��>�4X>uv>G%�>UjQ>��3>���=n
l�p�Խ�KR?����	�'���辊���c3B?�qd??1�>1i�%��������?���?Vs�?e=v>�~h��,+�zn?�>�>-��Qq
?R:=�2��;�<�U��O��L3����>�D׽� :��M�Unf�_j
?�/?�����̾=׽z��}j�=�x?��&?���uAW���t���D���I��&���fu��������q������� ����{#�`z�=��-?�8�?F?��˾b��w��6?��Y�>�1�>^)�>���>"�b>�"���/���Q����� g��D�>��{?�1�>�j@?��J?SZ?��8?.j�=�>1v9��f?a��=���>��?DD9?�V-?_@?�?�\�>�
>G�-�����dӾ�}2?��?�7<?��!?e�*?����KV���> -=*0�-q���;��ԽA��:s�=��'>[X?2����8�l���mk>��7?���>���>���#+��g/�<l�>��
?�H�>u  �j}r�hb��V�>~��?b���=@�)>���=�����Ѻ^]�=�����=�4���n;��|<l��=��=�^t�T��t�:���;p�<Y
?�;?�S3>޼>_O)�
����&�Z����?>�I/;y�b� �w=���Ǉ���B���>��?�+�?9`3�-�=X�=��G��Փ����P�����㽍��>Q�F?� ?��y?�6?���>5�
>/��������������F�#?g!,? ��>e��гʾ�񨿧�3�͝?=[?�<a�/���;)��¾�Խ��>�[/�;/~����ID�@�������+��?Ϳ�?A�8�6��x辳����[��X�C?�!�>�X�>M�>d�)�z�g�p%�N1;>Ԋ�>BR?c�>��Q?��v?�GW?�_8>:�A�z2��@���i��<1V >R�A?���?	T�?�tx?n�>�>�I������A��@�@�(����p� 8�=s�b>���>A��>|��>s��=����>˽�H���w=Օl>�F�>s|�>�>���>)v�;�G?���>�\������椾����=��u?$��?
�+?�"=W����E��H���F�>|n�?3��?�6*?��S����=��ּ�߶�|�q��>�ι>�*�>�ߓ=z�F=�c>
�>���>�4��^��o8��|M�!�?F?Ȼ=_�ÿ�I#��iɾ~˥���z>�ԇ�o��ӳ�=ό��o/�����/ѾEսʯ��W�Λ!�7�����&�sa�>H.B>d��<{�]=݀�;kUk�QN���B.>rۅ=�o];-��_=/(��,��<��#��b3��`f���B<L�=8ǾN{?fL?�>*?cC?�!w>d�%>�`�m�>@Q��W?e�g>/!E�=����+�ӫ���B����ھI�ھ| i��!����>�'����>��:>94�=�к9U��=�n�=Xjf=���I�3=Z��=��=�R�=_��=�>#�>�y�?7���K��_��{�dc5?�!�>no>�L=nZ?g�.�_ ~��ݪ��?���]?��@{��?X?ܷ%��>������U>���=I>��A�6>+��>���=M?7�>��\�M��*��="W�?���?��X?c���m��4#�>�8>>�)Q�� 2��Q\��`���U��� ?#L;��˾W�>况=��Q�žtm9=o 5>Z�Z=���vX]�A��=#����O=�ah=$�>I�D>�?�=������= `N=ơ�=MO>�;滘�8���,��17=	2�=�3`>��$>���>�??��/?!d?�v�>�fl��DϾz¾R�>J#�=+-�>�ρ=W\@>���>E�7?��D?3�L?���>7K�=���>��>�,��l�a�>]���:�<D��?w�?H0�>F2G<��B������=��Ľ��?W01?�+?N��>�U�z���X&�g�.�r���+��F+=�lr��TU�����m�.����=Oo�>���>�>�Ry>W�9>��N>��>6�>B�<�s�=sҌ����<j��N��=ꪑ���<��ż�5���O&��+�j����ݍ;q��;��]<}��;ʑ�=�.�>�	>�G�>��=mڳ�2%/>$喾��L����=O_���4B��Bd��~���.�`q6���B>��W>(���U*��L�?/�Z>ȋ>>dZ�?W
u?�� >���nVվ�����d�:�R�^ڷ=�d>ŗ=�f{;��|`���M�i�Ҿy��>�ߎ>�>��l>�,��"?�'�w=���a5�v�>�|��E���)��9q��?������Si��*Һ��D?�F��z��=X"~?O�I?*�?���>]��υؾ�;0>�H����=���(q�>h��o�?B'?���>��+�D�Uħ��C��|�|=�
ཌྷ�L��G����Q�x�>��q�5 �>J|�zj���#E�p ��Bߒ�8r��������>��k?�5�?�Ծ��{kv� �}�!�(�?t�T?���>@�?9�E?M��=�� �,.P�9?�<�P�?�`�?�n�?��>^u�=.������>wV�>� �?ߐ?~�r?�X7����>�'=g�.>�����>�';>JH�=X�=*�?��	?w$?v,w���g���4�.�c�1=���=`~�>�Ӂ>՜T>�ͷ=���<#��=�VA>���>\/�>'an>�ל>��]>)Ԣ�E�
�hc&?4��=ba�>�0?���>y�K=����:��<s���F�O�=�A`���@̽`h�<�8�+�=�aC���>�Iǿ�&�?ߞQ>���?W���*�T��lT>%�U>�2潎u�>��8>�y>5�>d�>=�>��>�+'>�HӾ$�>^���\!�Y"C�5R�&�Ѿ%{z>ښ��f#&�ԣ������OI��y��i��j��+��A8=���<QE�?T]���k���)����K~?�C�>v6?�֌��2��K�>���>i��>�O�����⾍��K���?,��?�߱>���>q&?o��>��e=>�j>B��9���np���Æ�Xfn�g/m�cZk�������76?���?��^?�W�M�c>ca?��@�������>����7���y�KV@>kB������#���7om��&�jһ=��I?�E�?�{/?V�#���s=�?t?�>�>�ޅ?��4?Fk?|�A�I5>��,?�@?��O?�Z?�qv?c?�=7��)��*c>�Gx>&v��"m��Տ�ku��9?s�W,>��=UQx��h���<Ms�=��Z���L=�^>
�T��m꼤��=�=�=#iW>#̮>�ua?���>O�>A3?H��M�=�3�þ��+?�P;�_��D⓾+帾����=F�Y?�?�?�/b?��H>�>��k9��((>���>�v>��o>]��>�7�d["���J=��>��9>���=/@��aw�'|	�hk����;�'>��?lf�>-�n�[�"=������F��Kf>����p� ������Y�\
G����_�?�Lt?r�?�?>r�x-�h�]� k�?��\?/@#?�/�?���=��RNU��d[����Qi�>��=�e9�V��_ǰ�;�k�띒��>!�:��Р��Ob>��oe޾�{n�e�I���羅tN=
j�	�W=��g�վ�"�<��=j
>0���&� �i���Ӫ�J? /j=�k����U��n���1>ô�>fծ>�8���v���@�𥬾�=A��>��:>�E��4��HpG��:�ӊ>�??�d\?7ޅ?ܬ��bh�x5?�8 ��⚾�Mt�k�?YE�>�?�0>$��=г�������a�VX=�fL�>���>�����A��e��g���c�)�Q��>o�?�g0>M�?�eQ?Ls?jpY?S�'?�4�>Pō>�j��Ɇ����?��?z`=���� ��d��x?��A�>;S1?��<�>�4?�)?��H?@O?q��>���<�I��M���>:��>�R�cTʿY>�V;?��>��Q?u�}?a�>@X�6OѾ���~>�A>l<?F�?�?0��>���>M���n�=���>mc?Z1�?��o?sk�=�?�q2>Y��>�k�=���>!��>>?�EO?Y�s?��J?��>(��<}`��},����r�8`N�uF�;#�H<y=�����s���η�<4��;�m��ǉ�����iFD��я�ώ�;)��>Ԡu>Ey����5>ž퉾qO>>�£�.e��0S�� �0����=[т>��?k��>��!�Ǝ=�K�>k��>���'?�?��?G=4<�a��־d�M�yǰ>�B?4X�=
l��ڔ�u�u��e=��m?F9^?��O����Jb?] C?��۾R��r��z���5�!9P?�-?w��"?^��?Z�?{�?�A�]�v�N$���f���1A�p�=u��>�"	��GL��G>�"?�D�>��F>S�=@��`OF�j0��Q,?!��?��?��?�}>Tk�	�ֿTW�����h�X?V�>:~��^?�&>�/�ݾ1瘾�	w����������#����ƴ� 2�Ħ��D��Sa&=���>�^?� [?cU?��ᾗ�Y��Y�G�~��Y����Y���?���G�SzE�#�y�ǎ��1�"���ڐ;��D��wT�e׷?
(?�[���>��g����w�ľ��Y>�E߾�B����)H��a
=���=�BD��7��	޾<
?�x�>V��>8R?]w,�{7�6D�
^�iE$��<:>I��>��>�س>lE���7���(�į羈���@M�ANw>�Tb?�FK?��o?d/���/��ρ��
"���2�s{���&C>
e>Z8�>��U���أ%�wC>��q�(�ܫ���	�R�y=*�1?��>hM�>3*�?n?���W����}��	2����<6��>�h?b1�>�Ƀ>��ͽ�N!���>�~U?���>�
�>���$�^z���&�U�>���:��#?2�>&<��_Zo�C*��,�z��[�}�>V��?����
��6s�>�e?�a%=�q7>���>��D=�����6����.�>�.?�p�=�@>���|�3,R����>V_G?YD��,������>5�t?W�:?O��>]�r?f��>���q�!>WD?\��?(d?�%�>�;=1ܫ�c�v�/}��H���}j=@R0>��=w�;+B��?35���d�͐��=��=�s=	
�1�պ�I=߫�<HϞ���>Vmۿ�BK��پ}
�^�A?
��ꈾW���^d��e��{b��K���Xx�p��'��V��8c�:���<�l�;��?2=�?/���:0��ղ���������7��>��q����O�����'����¾��d!�3�O��$i�R�e�L�'?�����ǿ񰡿�:ܾ4! ?�A ?5�y?��5�"���8�� >C�<-����뾬����οC�����^?���>��/��q��>ۥ�>�X>�Hq>����螾71�<��?5�-?��>Ŏr�/�ɿb���{¤<���?0�@4zA?��(��쾨}V=���>�	?��?>nV1�G�����_�>�9�?}��?̖M=g�W���	�kwe?��<	�F�2�ݻS?�=��=N�==����J>�T�>���CA���۽��4>Hǅ>{@"����pd^��þ<�]>�ս�H��6��?Z偿�σ�y�3���
-���3?A'?1�>�
=?͚G��ֿz�L��2S?�r�?1��?�BE?�K��6�>�1��{?G�m?�0�>�*��Z�cὓ���9ԾF^�@�U��J����==M>DZ=J������>�
��j��ƿf�$�Tl��;=rXֺ[�\��<��&�T�sM��0no�M�轆�f=ŕ�=7(Q>{Q�>�V>��Y>�UW?�k?�4�>"f>��es��= ξ����K���3�������������@���߾��	������S�ɾ�%=���=~8R�䔐�� ���b���F���.?Pl$>I�ʾ��M��5-<�lʾ)ͪ�v��
���0̾�1��n��˟?�A?+����V��3��Ͱ��r�W?AG�z���ܬ����=���Y=21�>ez�=��⾵3� mS��k0?e?=p��6T��*>D� ��t=�+?;�?�\[<'\�>�]%?�*��$㽼�[>�3>S��><U�>&	>����=۽��?�T?nN�朾��>�m���z��:b=u*>�I5�ll뼷^[>�e�<�ǌ�ijR��%�����<(W?>��>��)�q��a�����9Y==B�x?��?�*�>�{k?�B?(Ȥ<�f��i�S�c��Yw=��W?m*i?и>͈���о%���r�5?�e?�N>H[h�l�龄�.��T�S%?;�n?�_?Y����u}��������m6?��v?٫^�F���/���cW�E�>G�><6�>�q9�j��>,f>?D�#�;��F����.4��מ?��@2��?'@<���`k�=�G?�U�>��O���ƾ�[���	��vs=��>뜧�_iv���˙+�'�8?���?�&�>%���&���a�=�|��"��?O�?���O�A�ܲ�]zr��_ �F�x=%�<Ze\��;]�F,����-�N����#���k��]��|>�P@�����>L		�)aٿ�`���X������&���./?�n�>F�L��;���h���g�b�/���#�Ç$����>�F�=�oW�+l��Aℿ-�$�����ߜ�>� =���>J���ˎ־���X-��m>��?��	?�3+>dמּ}��?ʽ4�ߒ޿����#���8?i �?oz�?V\R?
�>��8����5����J?cl�?��z?G��=�"����&=%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�\�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�^�_?/�a�R�p���-���ƽ�ۡ>��0��e\�NM�����Xe����@y����?L^�?j�?���� #�g6%?�>a����8Ǿ��<���>�(�>*N>LH_���u>����:��h	>���?�~�?Rj?���� ����U>�}?�ҷ>M�?�I�=��>��=���uA���#> ��=KG���?r�N?�{�>���=�S3��l.�>BF�-�R�=��1jC�눈>�Va?��L?,ef>ⰳ��#��a!��:ͽ,�A��}�?��u5�ޅ�j�6>��B>��>	�>��%Ҿ��?�k���ؿ{e���a'�(4?Y��>7�?�����t�f��-/_?Ps�>D>�@*��J%��\J�s��?�F�?F�?D�׾))˼k�>���>@Q�>ޤԽ���M����7>�B?�S��B����o���>���?@�@�ٮ?>i�P�>e�۾2�}��Do��n������$<A�?;� �]a>��>�_��*i�r��pz|��i�>ܛ�?S��?�O�>3�?J`��C����9E]>��b?�f4?��=�U���&�>���>U �#����þnYU?��@8�@��P?�|��J6׿of��}y�U���,�W> 
�=�߫=�G<�y	Q<'��=%* �a���
D�=�H/>�>�#>|�>)8I>��>!���*��� C��r�I���I-�����[��Jl���1>���辒��>c��X���o�9�Im��熾�C�7d>��S?�.F?6{t?u�>O���� >P��c�=��/�We=>ú�>!�<?��G?�e3?���=I���ld�
�y�r:��,4e����>po>�+ ?JJ�>���>�h�F>ä�>��^>��=�D�������<�js>@=�>�?.=�>�A<>k�>�ʹ�+3��i�h���v���˽ �?y��Y�J�0���4��7���t��="e.?#{>��>п���]/H?�����%��+���>o�0?�cW?z�>���J�T�.<>�����j�OI>� ��pl�o�)�>Q>Ck?��f>�t>.�2�ė8���P�,毾�*}>�g6?Wf���8���u��iH�c7ݾ�KM>7�>l�9�r+�h֖���~��i�W�v=cX:?�?q���fϯ�T�t��e���#S>��[>��=ݭ=�FL>��`�m�ǽ�G��P,=y�=�^>D�?ud>`|�=���>����I[�/�>�U>�u%>*�>?�n?�"D�ʃ���愾�s-���x>���>�F>�E�=q�N��b�=��>ߓa>�\��,�����
?�dk>p��ʩZ���7��D=�b���V�=���=3���B��(�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ1h�>�x��Z�������u���#="��>�8H?�V����O�g>��v
?�?�^�੤���ȿ2|v����>V�?���?Z�m��A���@�n��>0��?�gY?�oi>�g۾x`Z����>ʻ@?�R?��>�9�}�'���?߶?ٯ�?�I>�x�?~�s?���>8�w�D/��������}=;4�>�w>T����XF��ē�!_����j����#Ob>�5%=\�>e_�w���G�=���]����e�G��>�Tq>�MJ>U0�>�� ?���>�ř>�=�苽ր��Ė�#�F?�݌?�	
��_���1;���=H�G��?��2?���?M��~^�>��f?��}?~`b?���>����j��Pw�������D=s|T>�� ?���>Ƽ�VXl>����F�jɞ>��>-Ȼ��߾b����"=���>�?-�>�U�=�M%?;��>��>0?v�.������UP��\�>��>w�>�\�?*~#?tp���$�C�{�����w�i�:N�=I[|?T�?
>
������($*�뢯�sUU�%R�?Ljc?W׽��/?�?�?ʵm?:X?TH^>�.��);U{�h 7>\�?V���@�h�9���ƽB?�?+�>�%˼BГ�z������ѾP�?@�b?�*?����}d��;ؾbY�<��Y;��r<��ںj6G��>۔9>[����6=;>S�=�8��yP���Y���>��>��)=Ce[�g�_�=�)?S�(��+�X�F=�s��V��X>��>�־X?>��`ς�����<�����2���?dk�?��?׭ٽ�Ib�d�*?�Ϗ?�4?s�>����L���1���\�@�r������X>�w�>`	Խ��k������e9}�ٔ��+����>ӷ�>�S?TA�>'c>���>(j��&�#���W�
�U*6��a�/�#��������L��u$���=殾L����s>�g�3G�>b�?�]>�N>@��>.}=��>\�>D|�>A�]>v!j>�z�=LЇ���O��gh�
DR?����]�'�.��q����8B?�td?e7�>�h�������{?O��?�v�?�Xv>zh��++�c?�>����g
?O�9=	��E�<>C�����m��u��E��>��׽�:�UM��ef�f
?Z+?3>����̾U׽'Ⱦ́<��i?�##?s�[�?�G�y��Z��I�N ��~�����S��Ѷr�U�����������&�)0R=Ǧ-?��}?�n�O�־5���n�v�Q�&�>2�>��m>���>�(�>wƾ�Q8���?�E "������>@*�?���>��I?֕"?q9l?U�K?Ƶ|>�&�>'���+�?K�4=�?P�?>Y=?�[?5�8?�(?8��>��
>I~����v���?�%�>��L?'?l�G?\<�Bx��rT�>h_F��>��J�/S?>*��*%��/��] >|��=��?�q��)8�#���l>�8?O��>���>ok���?��4�<�>>Z?LU�>���t�q�}w����>�6�?���y�<q�)>�j�=*��k�'��N�=��ǼPV�=�Å���6��<D[�=6��="4��y^��;{�;-a�<�B?�-?5��>6�>�,���D$��9���(��L������	>�n�UɈ��ؔ�7
Z��M>Z��?#X�?a�f>;z+>��o��p�煾$j9����D�m��3?�S)?K71?�u�?h#?^$�>���<���Y]��݌���I�_?q!,?ي�>Z����ʾ����3���?[?�<a�˸��;)��¾��Խ��>�[/�"/~����D�H󅻻�����7��?ۿ�?�A�$�6��x辶����[��Y�C?"�>fY�>^�>j�)���g��%�C1;>���>1R?�g�>|�M?��u?��[?�;>U9�ʄ��LY����-;�0	>3G?'��?�T�?uw?x%�>�q>�7�Yc�����5��̽X{�+��=�Re>PT�>��>�Қ>h�=�Y��yc����5����=�iX>���>υ�>��>P��>~�<��G?S�>�������5���L��M=���u?�c�?�+?��=ޣ��F��M���>�R�?b�?�*?�7T�L��=Wzݼ�c����q�t��>�_�>�R�>oL�=�L=%>�>�>���O@���8�5�O�X�?��E?���=p����m��(9��UL��м>�:&��m�~���T%���=d=R���◾B޾%x˾ޏA�%"���ʾ������o
?�e>C��=��h;63�(�� =�?u=I��<�؀��?�qP����<A�o�+����2���u/���<,˾� }?�1I?��+?uC?	{>�j>��<�ܴ�>V��� �?AV>T�S��]��r�;��먾�ו�.�ؾ�2־3dc�͟�է>vH���>�
4>�~�=��<���=4vu=L��=�I��ڌ"=0��=��=��=�M�=�X>0�>���?x2��u	ɿe9Q�����%A?A�>Mp�>ZD>��H?�{�=��������<���ZZN?� @�O�?�07?�F�����>5�1����Xu=z�ýX�սy��=�M�=���>�(+>r'��h��!<B�?U��?��(?g���)�~LI>�7>T�>x�R�z�1���\�N�b�N/Z���!?�6;�U̾V��>�e�=�.߾�}ƾ�/=��6>C�b=z��U\�bp�=�|�ϙ<=>/l=ż�>�cD>���=�1����=�_I=���=##P>������7��-���3=�x�=lNb>E�%>d��>�~?�0?Ad?���>�k�=ξ �¾l7�>�t�=���>�ڃ=�0A>��>��6?7MD?�(L?{��>#��=���>�t�>w�,�5`m�n������,�<�J�?�Ɔ?Q��>��L<}cD�1o�|�=�����r�?��0?�J?�:�>�U����7Y&���.�눙�qG4�O+=�mr��QU�P���^m�:�㽘�=�p�>���>��>.Ty>�9>��N>|�>��>r6�<qp�=�������<� ��y��=Y����<�vżS����x&�:�+������;ﮆ;N�]<���;:�>���>yNf>��?���;�?��\��=�I���p@�cB�����D�ǂc���r�N+�~�.�*�>8B>$n�=Gڎ���>��>>��4>���?�z?#xw><�t�;��y!����;yJ���\�=¤�>���W�6��Ff��C��U��U��>�̎>��>@ �>��-�(�=�6sD=�E�;�3��8�>�ꀾ2* ��"�bq�j@���Y���]e��;��eL?/懿�@�=�ox?�|H?cR�?��>~�K�bF�s�@>�\|�fd����ac�A)ټi?"?N�>�1�HNF����lϽ;>TA��U��
����u�\�����y��=W ��8��h�g����a��OJ�1�y���?L�j?�͡?����-���8��Z\���<��?l:<?��+>Ⱥ>��>O鏾UZ�ƀI���,>`+x?Y��?�*�?�/8=f��=i� ��R�>��?��?���?�cx?�N.�W]�>s�!=`�>>S*�a>A6>V��=9�=���>4�?�o�>�ט�k{����1���[�z
i=f��=)��>=�>y?�>c�N=��;�`�=�q�>�R�>&�p>P>�T�>0k>������!�:�??�̌= ��=S�?�?e>�Q>���~�p=LI_��^��Tĥ�  ѽ'�罩��=��=�v=t�C�/��>�V����?�9�>0JӾ�'?�-��hv�E1�>u	Y>�"��j�>��/=��>�&�>��>�!�=d&B>g��=���F�=����M�����3L�� �9>�㟾����`	�v���'M�LrѾ���z�j���}�28��yH=8�?�0���g�$� �N�=��>��i>�:?�lu��3�q4>O��>��>����'���پ?� �?y��>���>��[?S)?h=���T���&��-�� ��U醿�0�E�g�'wy�3 �����D?��u?!|Q?Vݽ��>�?��@�f峾�Η>�4ʾ�.�<uv>В����0��&侷����)���v=�d>?���?�"V?�0�����<�~�>)�?U>տ^?��2?�h?
yJ�cv�>٩�>p�?�0?�At?,+]?��5?+ý8��>��르=0�U�%���9<-�=�<�R|=�t<�X�q�2�E8>���=t/>�2j����	����ʗ���>}�>�!�>)�]?�S�>Jˆ>d7?�<��8�W���8�-?{�,=K������4΢�Lz򾜩 >��j?��?��Z?��b>��@���A�42><S�>��%>�<\>ĺ�>'���/D�nh�=�o>�>�(�=��M��>����	�ΐ��8��<! >"��>$=1>���lR�=�׾6~ʾ>n>���{ϾK�rw`�MR�����xܷ>W�R?C�7?�6,>U��ӥ��Ʒ`�k�+?}gz?�J?�?>e=�j¾*�)���Y�g�E���f>��=���ZF��� ���`��@��^>1����پ��T>Z	����6�M�a�f������k=@��3˥��H߾�
*���b���\>i/=͸Ҿ~F&�Ȭ�gx��_�D?og�=fR���a��@��[�>�:>��>}��rC���r2�.^��|#>��>FWf>�eԼ��ξ_�7�-5�˸�>�<?J�d?���?{XI���C��GF�/ d��=��$���#?8s�>^w?'ȇ>B�1>����-#�,0R��R�p��>�/�>��_�;�����dI���Q�s�>�\�>��K>��]?�M�?GNX?�?\�8?^�>jy�>�`�=�}{�DE&?���?�?�=��̽�.T�'�9���F���>��*?�J�㔛>�?z�?�H(?�R?��?r�	>N6 � u>� ��>}[�>9�V��{����^>H?^��>-�X?0W�?Җ6>��4�6����������=�">��1?t�"?�?Ot�>� �>(~����=�׾>�^?؅�?��q?�w�=��>R/>���>/,�=��>���>�?�J?�~m?�F?���>�Y�<J�Že��� ��,s��u�����<�݈<"�ʼJ6�����i<�	6��2��y1ݼ��2�����C�����<�^�>z�s>����z�0>��ľ�O��b�@>���FE���ފ�#�:�t۷=���>j�?g��>�N#�峒=ʪ�>yC�>Y���1(?D�?�?��!;a�b��ھ��K�S�>$B?o��=��l�͂����u�L�g=��m?��^?�W�_��C�b?��]?�:�<�<�&�þbNb������O?��
?�H�(۳>��~?k�q?���>M)f��/n�����Bb���j�8,�=[y�>Z�y�d�-z�>��7?�`�>0c>��=L�۾F�w�檠�[?��?m�?��?��)>�n�S'��Ͱ�뚇��Z?���>-b��K�?H�>�����j����"$�]q�� ������$���M���1���ҽ�'�<(J�>.?"W?~Kl?�-ξ82T��S��ۿ?�N�	�n��	�-��� ��P7���l�7�!�ƶҾ-��m�=��t��=�q۳?�'(?�u(�F��>���IL羟���^.>w���� ���=�ɒ�E==��}=�ap�%4�Qȯ���?���>[a�>c�:?�Z���?�$L3���7�����nF>�>"~�>��>s�<<��*����7¾=E����@�>��Y?�wC?���?�5��z߾Ggu����k=>Y�b��=�A�=/�S>p��1�O���#�U�K�n���������Ⱦ��?�T�	?���>o̖>j��?(G?݌龒��=���V��ͥ=���>}M�?ļ�>�s >@��	�
�w
�>c�Z?�?j��>����ؾ�t�����z?��>b=?�>�c���d�����G���6�(�a<6�c?{���ɔ��u>�T?I>��=�?>�Kٽ%�������W��5>�?Ya�=��
>P֘��A;�]y��Ծ/�%?@� ?��w���$�+�q>��"?P��>��>.|?YO�>x�۾ �����>�,T?�+B?�g??��>u�a=���p����E�w�=��>��V>�FN=�=�D`��(I��'��=uW�=�߅�<L��+J<i8�� �d�q+�<��Y>gX߿$BK��P׾����<$�����b���`�邽��f� �K�[���SRR����Y�z���m�����Oܽ%��?53�?ȓ����J�����`���0�([b>R�Q�j<�����s��<4��`Z��s<��w.��4]��燿`�|�(�'?s����ǿ鰡��:ܾ! ?�A ?�y?���"���8�'� >vB�<-��۝뾱�����ο|�����^?���>��/��n��>ू>ǡX>VHq>���v螾�4�<��?	�-?��>�r�*�ɿN���A��<���?+�@{A?(�(���쾺2V=��>9�	?�?>�_1��H�%���L�>^;�?��?8�M=��W���	�_}e?�(<b�F��oݻ3�=�G�=}=����J>�W�>���JA�
9ܽ)�4>Xօ>��"�����^�_[�<y�]>V�ս['��z	�?#�s�M�u���4���d��<�\?�>$�<�e?\�%���ڿ�!`�z\?6��?��?f
8?T:k���>jR��q?1tk?��>"��8r`��|������҉����^v��e=N/�>��]>7�ؽ��C^��ߜS�iM�@���˿V�=y(��\�<�}[��ݼ,0��������7Y����Q��뽠w�;��>��L>���>��_>ڋ�>��^?�u?���>�Q>����[��3��%�U�H����W��B������ܾT��� ���������+�L	ɾ�1L��/�=TcP�w̍��5�2�y�6�P�S;?qQ>�¾�.�X�=x¾ӕ��
K��4����߾H��_m���?�KD?�'����C�$��{"4�wB���E?��a��E(��q(P>ʔ+=�!>d��>8�=�r��Q�ft��/?�\?�黾Ь��U(>;���w=˰,?,/?.�<q6�>�I#?��.�[M��[>��5>P��>^y�>C>٩������??g�U?�P ��2��\��>#V���t���K=at>�3�_��bNb>�1�<�/��g<�)��˯�<�(W?�>$�)�s�qb������U==r�x?��?�-�>d{k?��B?�Τ<�h����S����`w=��W?R*i?b�>����	о�����5?��e?!�N>�bh�*�龨�.�U��$?��n?_?Ń���v}�������sn6?R�}?��l��Z��28	�;ؕ�K�>�8�> �>�(�-�>�\B?��G�n��j���f�.��?w�@b��?�%~=!�X;�8�a��>�Y�>׈I�;ɾ:I'�Sx�ަ\="�>�s�����aI,�l۽/�_?�Ȓ?�� ?VY���̾�=�Ώ�)3�?���?c����<ؕ���m��8����[_;=<0r���������7�JȾ���g؞��fݼ̵�>vn@�#⽏��>�40��gݿ�+Ͽ�ą��8վBR���?�?�>E岽[��h�O%s�&�A�3�C�#���-O�>��>�]������{��a;������.�>�I���>ET��9�������2<�ޒ>n��>��>]��������?[e��37ο霞�����X?�f�?zi�?7�?V�4<A�v��x{�6v�5<G?�zs?SZ?��$�I.]��]7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�q�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>c����8Ǿ��<���>�(�>*N>jH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?���>瑄?���=%@�>c�=`��Q���g�!>�x>��S�ߐ?[.M?=��>�1�=M�:�#.��F���Q�:���/C�E��>g`_?�2L?�i>J����)�=q �sFŽH�,����l�G�Lt(�r��2>Ҽ;>��>�'D���Ӿ�e?6��hؿ�"HN��l.?�!y>Im?'��VH�-k��(�X?�c|>�������j��c$�����?&�?m?�<ܾX�,����=��>Q��>��%��}�0���3�;>ްA?rn�id��&6k��˄>�?Dh@�t�?]�j�fO?���x��@s���P�OY���">3R1?���9��>���>XL)=��n��t���@��Kvt>o�?r$�?�c�>��e?z�����Q���U>H�>�Oq?��7?L(+�W*�U�{��/	?Xv�M������e??T@N@F?ޖ��h߿�ޙ�8�������9k�=W%=}�>�"���>}�=C�O�����> �>@�H>?+v>l��>5+;>�A�>ܩ��ZB��T��[C����+�x����-��񾴹��4�ɢ̾�������1��@�k���e����=�-�=U&?]z9?�j?�#?��4����>+,'�
�,6�=�R�:/�>�Dh?@Hf?~ A?n�W��}W�\)m�X;c���� �>�j�>�M>�:?1�>�:�g�^>DE�>EOY�.�=P�x�X��;r1=�T=s��>���>���>i�:>`�>9������ngh�-�x���Ͻ�΢?8���ݬJ�a���ǃ��]d��L��=	.?OK>����Qп���H?Cn�� ��!�+��>F�0?Q$W?>�>�谾JQ�t@>g�	��Tj��� >e ��'m��[)���Q>�R?#T>%w>�\3�ա7���L�Tظ��V]>k�1?"ﶾ� >��q��A��پ��U>�ζ>�'�;������w����`���=	�7?M� ?e$���Ъ�3�n�� ���ZR>d�f>	�(=���=�UD>#僽�|ܽ�Q�V�*=rm >"f>�?B�!>���=�8�>�T����E��߫>��A>e�)>H�<?<�?� :�ݖ��*���8,�~�x>#��>���>#��=5�H�"�=͑�>�[n>���Ҋ����N�xFW>��{��g`�T*��~`=}�����=i��=����@�7�>=�~?���%䈿���d���lD?V+? �=۝F<��"�D ���H��G�?q�@m�?��	�ܢV�:�?�@�?��6��=}�>׫>�ξ�L��?��Ž/Ǣ�Ŕ	�D)#�fS�?��?��/�Xʋ�:l��6>�^%?�Ӿ���>�L������~����v���=��>��I?����%���<�F	?6?�����㤿�ȿw�u�a��>��?� �?*m�����nB��b�>�Q�?jw\?��c>W`۾��S�L�>��>?�FO?�u�>�|��e!��{?��?Z�?��4>GW�?��j?Kh�>��>���/�0C�����+?�=��#<�_�>i>	>�鿾v�B�C���Ί���i�t��,O>��0=a�> �ڽ���Ui�=���, ��)n�Oʼ>
�>}A>t+�>�$�>��>Z�>W[=�Θ��~�:�����K?���?+��r-n�mB�<�}�=:�^�X(?�L4?p�\�{�Ͼ�ب>�\?yÀ?l[?3f�>���<���俿C��}��<��K>�6�>"F�>v���LK>j�Ծ5D�bu�>%Η>���$@ھi-��k���L@�>�c!?Ƒ�>$Ʈ=}� ?v�#?��k>���>�E�����~F����>��>�e?�~?��?�"��l�3��������[�=�L>Sy?��?nM�>�H������(�W�I�D�yCP�?�h?�mݽ�?jV�?& ??{�@?دc>����ھ�B���>= ?W��Y9�"��
�,
?�?��>�f��{B��%!�������b�
?��W?��%?�0��;[��@ž�Z�<|Ƽ��_A�v��<�E���>v� >���;��=n>>��=:�l�?@:�Q�<)�=�!�>�x�=�:�J8]�K�-?Ƿ��21����=% u���C����>�;V>ˀ;�:Z?�D�0���"�����~�;���?k�?Iє?����:h�ݒA?��?�?��>#ؤ�N�������/Qw����S>�p�>9%���^���+᩿�Ӄ�����hܼ�h�>���>B��>*��>b�>{�>@P�n����	��3E�l�g��,�ߝQ������ᾗ���-���]n��	���w���>���8Ք>�b�>K�>*�>�?�}�<3�>��H>�<G>2��>��3=햎>��9>b�=��BKR?����!�'����s���J3B?�qd?	.�>(i�C���,����?ņ�?Ms�?>@v>�~h�{,+�Sm?�<�>���_p
?
]:=��M+�<"S�����~5��[����>�M׽� :��M��nf��i
?�.?���.�̾m5׽ج�ū=} k?*5?d��;W��(}�~Y�2�=����<��?����E�rgc��~��ʷ��դ����4��WX=9t(?��u?d� ���žQ���i�l��@���>���>e��>�Q�>��=����00��b� �����ɠ�>	F�?8>�`?4�e?��b?�k3?�9^=�d=>�R<��7?uy��9??޽N?�B?�A?�O?��>��G>�?	������)�>۷�>� 5?wQ"?hp)?Nپ)ݾ�6l>a7��ӗ��mA�D����7(���Ľ�g��N�=?� �vV?����8�����k>t�7?���>���>���;*���e�<��>��
?�H�>����$xr��`�Q�>��?V��pz=��)>]��=N|��q׺�`�=�¼��=F��B{;�<ꅿ=J��=k2u�������:O��;���<�_?�`F?л�>���>�7Ծ��������6����7\��=��F�=�`��S!��U�����l�fL>'��?t�?��>�\>`+��U��@_�q9���H��N�0?��N?��??�ȟ?�Jg?�n?u�'=[�߾�K~�����`�d�3? !,?%��>f��ϳʾt񨿢�3�S�?[?�<a�׸��;)���¾��Խ��>�[/�J/~����/D�<*���������?���?"A���6��x辞����Z����C?�!�>�X�>*�>e�)���g�w%�91;>̊�>*R?��>IX?6?,]U?��4>�I��2��nWu�r�4>�C��mY?�_�?��?��?Kz ?�OF>w�I��qϾi����Q����G�*Js���=֡5>Ǐ*>yD�>�ũ>���=�#�U���g�)��k�=��|>���>���>_h�>�gg>g�%>�wG?t�>����8����؁��#2��v?�?�*?�)�<
���_F�2����P�>��?���?=�)?�Y����=7&�Ŷ� j����>�ù>~�>=��\=x�>[p�>mU�>P�q����7�tu=���?�8E?�e�=lj���Z�@�������=�>���P����:�M��ۛ==\���k׽�����;�����I��TľSǾ�a����>�[R=�U�=�>��!=>�+�,5ٻ�=�6(=�4�=�7�Cvp��E��K�̡ݽ�?B�$tỸyx=���=��ʾ�r}?�mH?�q+?�/D?Mk|>�_>�.�!<�>y)�� �?�2S>YI��;��p9�*2��M͗�8sپ��־��c������>-%]�N�>n�1>���=�ѩ<<�=�%w=s�=�Z���-=��=C"�=�8�=́�=�S>B\>��?E���j6���%R�W���v,?�	�>�'�>�q��W?7ؾ>���������e�u?� @\��?��A?ʹ�=1~>$ߤ����=Q~T=4�Q� �˽Z>�d ��u�>>y6>��<���=��?��?�T?�,���v���j> <�&T>*@O��5�8m%��Ⱦm6پjk�>�2+�G侾�I�>pD>_���7�]����G��]2���Z;L0��[s�=j o<Н=S+�<쉫>�*|>��=̉`���>�G'>�s>�C4=%Oݽ��(��$B�d&���L�=ݬ�>�>���>v?�t0?aKd?�.�>�cn�G.Ͼ�������>��=��>�Ά=�C>KӸ>w8?��D?A�K?{i�>T�==Ǻ>��>��,���m��5�5㧾]��<a��?ӳ�?kw�>�hP<jA�q��:>��Ľ�X?x<1?�S?�*�>*��-��S�!�L����?�<��H=`ѽ���;���<N��A��yy
>�ԍ>4Y�>&`�>sN�>�cf>���>�u�>�f=cE�����=4s\���F��|=��>	6�����=t��=y
�=vG�;����=��@�m�m�<�<���^�=���>q@'>���>�'�=�����#$>�!����I��x�=�8��kA�IQb����|�-�� :�.�2>�2L>6o��?��L4? X>RY6>B]�?Y�q?C:!>X���	sɾj���Οv��o\��:�=�Y>��7��M9� �]�PJ��վ��>��>rR�>��n>�,���>���r=� ��4���>#��eg�Z��:q��7���ϟ��(i��i2��>D?B���O�=�}?z�I?���?D��>���	ؾD�/>6L���
=m���o�j��F;?D�&?��>����D�gh���9���=뼧�%�F������U�9�>��(_�>yҔ�"�����%�'M��{v��J~^��þA��>�p?-r�?�+]�\1t�e~�omW��J>��8?�Jl?�<�>s0?t��>	R����D+��t�(>�N?��?���?3C>��=ŉ�����>mO
?�9�?��?o�t?:l�:�>�=�>ʶ�3� >�>Q��=���=X?��?�)�>�e��ݑ��t�G��:�3n<i��=g �>��s>ad>�j>N��=l.�= �^>�>q��>�y^>�n�>a�>;���E����&?Ȏ�=���>��2?���>�=E�>�@����4�e��#b��Ƚ|ʽ'�^=S�<҂=/䭽��>ڹ��XI�?���>)n��D�?��Ҿ����lg>�=(>A,ǽ��>
#�=�֜>�&�>��>>�~>aO>��پ#�+>j'���5��/qi��F�W2>��m��5 �j}ؾ^�߽��C�������.��Iw�ߴ��8�E����=�	�?���\d�X@�1�G�k��>7�u>��X?>�?��tV�[��=�տ>��t>Z�
��Ǐ��w��lܾr�?��?���>��>�AR?4�)?����,���i2����ֳP��i�R��L���~��c���a�~?�(j?��0?�|��s>ﮆ?+>������<>���<m=��FP�])�=�}��ͧ������½��A�'�)=>�N?�mz?��H?1�C�Ȉ#���=!u?��?�A�?ЛW?�{?V�P�>�?�2�>�qM?��|?��Q?��4?���;���7�V=�r�<����xi��XY���]���A<��=���=ȝ=���=X�=��0>T�=��=�-;>5��<�d�<Tk=bk�=ϲ>p��>��]?���>���>Q6?8w��86������=+?��=��*���������>$�=[i??��Z?ڎ[>��>�.mD��!> ��>� >�o[>��>���M�B��[�=W�>�_>i�=U�?�����Gx��V�����<5�">�t?p�;>�`����=�bѾ�e�Nr>�_���4�m��fZ�(\�I����x>Y?[?��1?�_!>`������~#d���C?2̈?��*?]��?�&u>���_6��rQ�R���c�%<��>�=Ѿ{��`����r���{
�Hz&>�5�󬣾Y�_>��jI޾g�l��kH�S���>=��"�Y=qd�=:־,���`��=3>¾�� ����Ϫ�ƗI?`!k=�h���3W����D�>��>No�>d;�-\w��`@�( ��Y��=��>� 8>������~G�Op���>޹8?��Q?�4�?��پ�`��^�z���_��Ф����O?p`�>�p?pK�>)y������~E��zy�0�M��l�>��>����N�E�����i*��4J��}�>z�>HѤ>3F?�}X?�D?�;x?�?��>���>�wp���ܾZ&?|M�?%��=�\ν�W�=~9�g�F�a^�>�*?=�A�p�>��?�E?�o'?�Q?x�?7!>e� �� A�]e�>���>{W�Hï��>b>�IJ?)��>K�X?\փ?7�@>F�4����+꯽�D�=Ŵ>�g3?��#?Ps?��>�0�>����̿c=o��>�]?�=�?�{n?���=�F?�X>��>��>>�>u/�>ˎ?�B?��f?�*K?���>���< ý���̆��<���N=lϔ<��<= > ��@O�u'���u�=:��<~��j�y���`bw�\��)6f�v{�>�^v>	����<>��ƾL��<�5>yG��Y����憾Q'����=;K�>ª?��>�( ����=�L�>���>.����&?�?�C?9�<]�`���о��E�Y:�>B?���=��m��K\v�ic=�~n?�*]?�L�����r�b?�]?�$�x�<�f#ľ,Sc�=�龂�O?\�
?�H�^:�>B�~?Wr?���>��e�@n����M\b��uk��ٶ=�T�>Q���d��,�>�u7?M7�>�c>!��=�"۾8�w��F��=?��?���?w�?��*>��n��.�fZ0�P��}S?v��>�+���9?`���jо�R���?�����IN��*}��3+���*��B�� sS����,J>��?]p�?w�R?��`?24~�L�S�$h�6���6=�-���W5�Y:���\�Z��0����A��ᾘa���C��
�l�^xL�P�?��?4;3��;?�Ȑ�v�SF׾�*>���r��x��={z�?��=7��=�N���V��B���?�}�>���>$�>?�O��Y8�>8'�a�;�7���'>�F�>j��>���>/:7�ؿM����?���ت����ڼ�pw>b�b?aIJ?M�p?����j1�ɞ��.7����V𫾩�K>��>��>��O�J���z&�r�>�Gq����|Q��Z	��z=��2?���>���>GÖ?N�?��x����g��0��<�ϸ>�g?�+�>���>BoŽ�i�jI�>Xz~?N�>���>G!������|u��0�׼�>�>$��>�b>�n���k�*���䑈�k�(����>��9?�ڱ��A��o>��i?���=��<H��>"����������O��,>��?ue>,	>�
߾#�M��R������=<(?�w
?F���`*��x~>I�#?]R�>�ơ>m݃?L��>�о�<�?�R^?LJ?�>?%��>�?=����y����(����<9�>��Y>vڑ=Ȇ�=cA�/?]���ehn=���=�ѯ�鼽�<`���<��=�n,>��ܿ$K���Ծ��'����Ð��ؽht��&����倾5�%���p��%a�d�g��ˏ���p�!R�?+��?����8������q�y�>>qv��/U��p��6����0���#�\aO�lti�Mh�C�'?�����ǿ찡��:ܾ(! ?�A ?/�y?��2�"���8�� >7C�<.��뾭����οE�����^?���>��/��d��>Х�>�X>�Hq>����螾d0�<��?2�-?��>Ŏr�+�ɿ]���ä<���?0�@ekA?�$(����eGX=��>�6
?I?>�O5�{���ұ�x�>A	�?��?�K=�hW��� �_�e?e<��F��RۻO�=ϡ�=Ź=����I>�ʒ>���]@�B�׽X�2>A�>���v��_� �<�^>o�ֽ朖�E�?O:����}��)N�A򜿔�<P��?��?=�>�@P?�GH��[ۿ�~>�"�i? '@�P�?a0?�ӷ�5�>�u¾L�c?�sC?ۢ? J־��S��4\<�H+���þ�f⾕n�AOs>U*)?1�>��ƻ=���k��:}#���=�����ſ�^"�����.=��;�*��}�������U�䛡�`�p�!���"=���=��D>%�>��M>+�T>ġX?'m?��>� >]$Ͻ5���Y׾�����������]�!�ɴ��FP��� ����Z������$о� =�c�=�R�z���� ��b�8�F���.?c�#>��ʾ�M��#<;�ʾT���Uゼ�ϥ�\̾r�1��n���?��A??څ�hW�
������*��l�W?b�����֬�ާ�='��X�=��>�J�=���&3���S��s0?Ue?:Y����!�)>!b�w=(�+?#�?3�Y<\^�>I%?��*�W�F$[>E3>w��>Y��>k�>�@��^۽,w?�T?��|؜��$�>eG��oz�F!`=y>�=5�)d�t[>T��<3ڌ���_��Z����<�!W?@��>��)�
���]�������<=��x?�?.%�>�lk?��B?R��<�n��k�S�6"�c[w=�W?�i?r�>@����о�Q��J�5?�e?��N>�ih���龅�.�H9�0?��n?�[?/P���u}��!����P6?n�w?��`��Ǣ�hR�`Xm�oo�>'��>���>�3�Oӻ>��=?��$�)F��U1���O3�2-�?S�@h��?��<=мF7=��>��>�=��0���R��V:��s��=���>������w�1��Ab���=?���?�?�o�������=ܕ��Z�?
�?*����%h<����l�8n��&��<���=�&�bZ"�N��]�7�%�ƾ7�
������r�����>�Z@�f轹*�>�:8��3��QϿ����^о�cq���?O��>!�ȽB�����j��Nu���G�V�H� ����S�>��>Pؔ�n��7�{�Oi;�_Ӟ���>�m���>�S�0������w�4<��>���>���>����潾ﾙ?�k��9ο����@��j�X?�d�?_m�?�t?��7<h�v�u}{��z��.G?�s?6Z?�V%��P]��#8�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�x�_?Tb��q�<.���ͽ�A�>�_-�T>Y��$���O%e��8����y�Sҭ?�f�?�2�?w����"�"J%?}��>�����ž���<
�>�{�>��N><a��s>R��US;�LS
>(��?nZ�?��?�y��������>�}?�i�>ޯ?�2Y>��"?M�=��2<=aGz>�U�>�%<��.??VE?��>�>����A\��XA�[<���/��cW�^a�>�Q?�?<��>c�:��x>X+��r��_>�f!�iFC�1����KJ>Ó�=A�����ꂾ��?pm���ؿ�h���j'�C04?㯃>��?��ٽt�Q	��8_? x�>\8�3,��p%���C����?2H�?x�?ڷ׾8M̼� >��>�G�>~�Խ�퟽q�����7>$�B?�*��D�� �o�[�>���?�@T֮?i�Kk?���ۛ��2x���:��ž]>[�E?r�Ǿy��>�W�>�: �"�ͧ�o�w��c�>�?���?���>�N�?e����;y�6�,��T�=��r?��5?P��=�y���>��	?:�Ѿ�e���tؾi�?T�	@p�@RX?������ӿ����Ʃ���̾�S�=� �=�?>������=��=G�R<v��<�)>G�>3�p>��T>IeM>;P>&6'>����\#��N��X:���<��k�&L��u-�y�� ey��V�F�M���Ç���q��%��.~B�T���^�@�=�,V?��P?�Gh?���>�\!�?"N>)ȼ����=Y½H~>��>�-?�I?�#?�<0�����^�����oƾ:�_��P�>��=2�>��>�a�>�>=���=��'>^�K>� �=��;&|�ѐ=9�>�Z�>)2�>/��>�C<>L�>�δ�"2��Q�h��w�]̽8�?�����J��1���:�������i�=Vb.?6|>����>п^����1H?����(��+���>��0?bcW?h�>���|�T��9>�����j��b>a+ ��}l�c�)��#Q>�k?��n>�b>c� ��O�nRN�x=o�#�v>��A?�_���@���r�8UP�����oM>SC�>�S�:Vs�tg��L怿���jȶ���??�F�>�ͽ�o��X��D����>e>=�=J�8>�{F>�'=`v��z���e�<�V=�$>C?��,>��=Px�>|���lS�9U�>X�D>��0>��??�&?��䀘�����Q�,���v>ƀ�>���>ٺ >�bM��5�=5e�>�a>V%ݼK#������&?��V>�|���`�'x}�9�i=�ם����=�=[����<���+=0�~?���1䈿��5h���lD?y+?�=�F<W�"�I ��/I�� �?l�@5m�? �	���V��?�@�?v����=+}�>�׫>�ξ��L�K�?ƽPȢ�!�	�p)#�YS�?��?��/�eʋ�8l� 7>�^%?;�Ӿ
h�>jx��Z�����t�u��#=ߨ�>�8H?�V��b�O��>��v
?�?�^�橤���ȿ3|v����>U�?���?9�m�uA���@�D��>��?|gY?�oi>�g۾�`Z����>��@?�R?��>�9�?�'���?�޶?߯�?B!H>Vn�?s?:��>��t���.��r��RL�� �=n������>x(>�k��w�E��m��gT��B8k�5���]>�'=ᶶ>�_�ڵ���:�=P����sf�-�>��o>~�R>Ц�>�� ?��>�>��=�[��"������.�K?��?���^+j���h<T��=�tg���?��5?&��A?ƾ���>)n]?��?5�Y? ��>�U������{��n��4r�<I>��>���>���d�T>�Ҿ��;����>3z�>��̼r&޾遄��jK�|�>1"?�:�>䠬=�� ?}�#?��j>�/�>�aE� 9��}�E�װ�>u��>�D?��~?��?�Ϲ�`X3����桿�[��/N>�x?�V?�ȕ>2�������o~F�b�I�������?�rg?�A�b?d2�?,�??ߦA?I'f>h���ؾ������>|a?l@���4��U&�nw��?&�?���>���N��S�4��o�����?��[?�*?]�����c����pl=$��3�<���<2����=>�#>U���X�=��>�G�=��p�
�0�?=¼��u=!a�>���=t�7�O���m=,?�!G��׃�,ј={�r�lsD�ݺ>�JL>�����^?�t=�(�{����Ww���T����?~��?�h�?���h�a"=?��?H�?m�>X<���w޾È�oDw�:�x��s���>F��>�4m��徰�������F��Wƽ��6� ?q�>Ʀ	?��>�wJ>[�>�����&$�����*_� �X����X5�B(�GL��b��0x,��M��߶ξ�샾���>�ȓ�M�>��?M�w>@�}>G�>�Ƽ���>�]>x>%~�>L�L>]�#>Kɵ={�6��8뽨KR?����þ'�p��*����3B?�qd?�0�>�i��������?���?%s�?.>v>�~h��,+��n?�>�>����p
?�K:=�;�oB�<T��ʻ��3������>F@׽�:�"M�nnf�j
?W/?w���̾L=׽I+׾y�<�fZ? #?,��6�O�_�}��6V��:K��u+��ʕ�灡�)�&�Ct�FP�������Y��1���-=*-?$Z~?���A	Ծ���W=s�h?��,�>6��>�
W>T��>z�2>�罾#'"���R������f�I�>���?O��>gH?�<?�W?}NC?�b>��>�6���?��<�O�>r�>.�7?v�-?��+?N�?�K!?]cR>�6����r�ž9?
?�W%?!�?�?�M��ñ�ԯʼ!�����Jý��=�p=/Jͽ`շ���<�Rb>W�?NM�=6�<����Xp>o5>?�g�>��>�c��hdR��)O=��>�%?ﻕ>�G���m��R�4a�>�U�?{��4߮<0>��=����B =}��=?���,\=�O-���E��D=t�=�R�=�f�]x�9��jy;�;w?��7?~ψ>"�m>l_��5��p���䦼k>z�C>�F�;�߾��������$]�8Ԉ>`f�?�$�?u=�9�=��=�Ml�0���D�d��`M9���&?ʒ??kX ?��?�R?�%�>܇#=>���S���ጿ�H4�tZ?v!,?��>�����ʾ��ԉ3�ڝ?i[?�<a����;)�ߐ¾�Խձ>�[/�g/~����>D�����^��5��?쿝?:A�U�6��x�ڿ���[��y�C?"�>Y�>��>S�)�}�g�q%��1;>���>kR?T��>JD?�Qq?��`?�P=�M�����wV����>��>bsa?�ǂ?�ݓ?��?��>U_x=�X��� ���$�l����	�����թ=Tݒ>��>�k ?X��>PP>�G=��?��*I�Z1 �O�0>�9�>��>A`?��>#���G?���>�Y����夾3����A=�U�u?>��?n�+?ݨ=���m�E��O��$?�>�o�?���?I4*?J�S�L��=(�ּ�Զ�%�q�"�>ɸ�>(�>}2�=h�F=Kw>��>$��>M:��f��q8��M��?F?���=��ҿR�O��b{�l<4���>�r:�)�龼�þ1��!�>�M�v7�&��E��{ ��a�m}���O����?�\�=�qݽ��='�w=ݰW��+</d�=;A�ع�<�r�f�����e��ј=�PA�9zü�ܰ���޼7�x=�¾�?�&J?��2?�(0?�L�=i�>����.~> �S��F?�d�>�p=�k���t�;W�'� �4�޾|]Ӿ�ᇾ)���6>�<���=��>�2F<��s���=��5eB=�X8:pn�=��>�J=�K<e��=�L�=��>���?�ٛ������ن��ɾ�?ֱ>�r�>SL�<�"?�C>����������g?p��?Ȑ�?��'?�#罐�w>	�Ҿ}��=+��VY�TJR>b�:>az��I�>���=f�C����p���?}�@�=?����ڿ=��=��7>�>$�R�ˮ1���\���a�RZ�ޯ!?�\;�'F̾p��>���=�U߾�pƾ��/=͍6>�b=����_\���="�|��x==�j=���>�XD>��=�ݯ���=�gH=ʹ�=6SP>.˒�g5��,���4=<��=�Tb>g�%>���>??? �+?2b?�>a�Q��Ͼ��վ�yx>�H�=%T�>�p=?�<>խ>v�2?'5H?��O?3)�>8�a=���>��>+'�G�i����m3���RH<��?��?���>��J�
d�V%��A����v�?]i/?�?��>�U����9Y&���.�$���Zm4��+=�mr��QU�N���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<{p�=ጻ���<� �����=!�����<�vżЗ���u&�=�+�6�����;p��;A�]<|��;]�>���>+�>�Z�>�D�=|����E">�ጾpM��=­��;�@��\b�iz�.H'�w9�43>�DP>��������9��>V�t>˂!>��?-�t?��<>���Y�ɾoF����o�$8�G��=��>O{A�N�9��c�&eS���ؾ���>���>��>��l>�,��!?�V�w=v�5Z5����>|y��Ϟ�H,��8q��<����i��/ɺ%�D?�F�����=� ~?3�I?��?_��>i����ؾ�90>�N���S=��
q��'����?~	'?�t�>�,쾿�D�W6��z<H��=V:E���i���>�d�d��=
;�R/�=�5��K/Ծ�.�������9�C��΂����>��?ŷ�?y���Q��X��]Z��<㽟�?Уd?4/>�[ ?e?,^w����-rT�8�9>1��?�c�?*\�?��=���=�䶽r��>'�?xȕ?㔑?e�r?��@���>M@<�!>u9w��2�=��>,��=I=�=��
?�8?��?k���If	�͗�s���\�p4"= �=Jq�>�H�>R�r>!��=�J�=~�=4�W>�(�>Z�>�
`>أ>���>m߄�:#�Ҋ+?`��8&>��O?�kh>��;>Rm�V[���6�D�t�Jp��=�9=BB>��A=�8���=h�>��˿�N�?�3�>�Ǿ&�?oPѾ��F���>��>^��\�?	̘>v�>�Ԏ>7~�>��,>��C>�!�>������=�R�,��CL#��&V�.���|P> ��O�7�o����Q�9�˾�L��pm�I����B=���^=A��?� ��6�c�.#��C�G��>^:�>FoA? cz�O����a&>]��>ϧ�>�Y�[^���x���ž.k�?���?qĢ>�?H%'?rt�>޸,<�/�>�%�����0w��鄿N�t���]���S�E�����Q|?ƿ�?'�&?�g�<�tA>��v?T�4����C�p>�s/�d|2�,>��M>jQ���
>��'��$������D��� 0?k=v?��,?ܩ���6��T >�+?�N�>]�g?#�?h�L?L �� ?��?��>�Y?��?�ZT?]�?�]����	���e>Yy�>5(=��������нAQ���l>!8�<��z�8?�=lW�=u���X�4<#�=�:�:�9=�;�=�Xp=�p�=�.�=�T�>e�a?D��>�^�>�.9?�Ħ�K�4�NU־��?�b������o��󁣾M��-��=�yn?�٬?��X?H�Q>�;���;��@�=�ʎ>��>û<> �>�����2����=6�=i*�=㣼=p��?���! ������<��>��?���=6q�3�=����ԔF��H>�2T��.���b��R��[�?���VL�>�`? �1?��B>%�׾&��Yh�`�=?!�g?g��>���?ވ�>�������Vd���v�'_�>�V�=�6�2���Mϯ�Z+^�8 P;w�>-��z����/b>�Y�z�޾�Wn�5�I�8羙pL=���%�T=�/�`Q־�o�����=��
>����V� �����ڪ���I?Cg=T�����T�Q����>�w�>ޚ�>R�8��sv��g@�yz���>�=
�>�):>������20G����>��>�8J?��Y?���?�;���si��G�e�b6�n����?���>��?�tA>6�p7��Ȣ&�NY�e�/�-��>�&�> 	��
r�L�̾?���$�ܣ>���>k�>'?eV?3?<�\?j�9?N�>��4>h�L���LP&?���?;��=o0Խ��U�In9�{8F��;�>Z�)?(�C��1�>��?5=?+�&?ׅQ?s?�
>�q��8@��4�>��>�gW�.���:`>�{J?_��>.Y?���?J|>>@�5��뢾�Ū�r��=!�>3?�\#?�?���>$k�>OD��}£=N �>�ed?E��?�'q?�$�=]��>��K>���>W0�=뺮>Y��>t�?P�G?{l?�H?��>\�<�������yU�Lճ��E^<��=�2}=&z� ��	��#��9>�;R �y�׼��~�k������uǼH\�>f�s>���	�0>��ľ�F����@>�Q��z\�����L�:��ݷ=��>��?䦕>N#��ڒ=���>�5�>����0(?��?R?��!;��b���ھ��K���>�	B?@��=C�l�=���@�u�Qh=��m?H�^?��W�4#���a?��d?�b��� ��.㾰�����eL?�)?������>�>�?��?3n?�L�6�k��d���'��"�T�@I�=�d�>G�
�ĺU��mp>��?��>�p�>�%>&~վ@pd���&�@�?2�?Hϳ?��?�#M>,ⁿ��̿mo!�.���
�K?A0�>��1�'?�#������.��ǔ��Lnվ�0¾���'���M�����0����!����=�?�mq?�da??D^?�(߾��R�9�a��\y�f�R�����+�}P��+���Q�8s� r	���־��[��=�&y�� @�^�?�a$?�3���>����
��qm;g$=>g��w8�T|=~|���lD=��O=�qh��I5��R����?��>q��>� >?DzX�i�;�B'0�5�8�����2$>�(�>��>�/�>���I6�x��l¾��u�נɽ�
z>X�c?�J?��n?}���
3��G��,���_���V���IH>^�>�E�>�^L���`l$�_m>�k�s�io��鑾��	����=qE3?fu�>N��>�?�T?|6	� ?xs�#~1�l��;��>ޡg? ��>*��>vǰ��E�Q.�>6u?��>��?,v_����4�o��pn�e��>��L=���>�Ä>MD��[G�N/w�݌x�e�/���1>��M?���Kl��ѩ>Pkz?�����<�%�>�j>�'�Tľ/��#��>�2?�]>��y<?�� J������R���H)?�E?�Ԓ�I�*�"H~>�%"?`��>(�>*�?�2�>`gþ��0�V�?��^?�@J?[LA?�>�>°=�����Ƚ&�&�52,=$��>�Z>�<m=��=F���m\�)��b�D=�!�=�μ�j����<� ��̺K<՚�<�3>��ۿ��J���ؾ~��_����@���B��uJ���F�y`��^���u������9���W�1�c�*֋�T�g�/�?3��?�P���ֆ��Q��?{��O� �vh�>�8p�ϱ���6��
|�t퓾
T�ۆ��?`!��O�Dh�Je�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >[C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾u1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@�nA?��'����RX=r��>�Z
?��?>��7�,�������c�>���?�^�?`tA=��W����)f?PRM<u�G��6лԒ�=z��=��=�r��J>n�>ݩ�6�B�?Aڽ%(7>}g�>�V#��f�v�\���<��`>8�ѽ<f��@��?(f��n�?�O������=ƨ~?�>1?e�>��X?m�y�~u̿�g4���d?��?��?�A?;���
?����\?�?���>C�Ѿ#a��ʐ��T�����')���9���A=��>��>��=�� �����eݻz�=���-*�����	=�.�=#&�=�w��O׽XB�{��A���� �����<���Te;<"�>��B>�p8>��>��]?��s?Կ�>��w>8J¼�T��� ��7�򃾒b��-˾U|@���`�S_�o���i���x�������#=�?:�=P4R�����7� �y�b�(�F���.?�g$>-�ʾ�M��+<vdʾ�ͪ� L���0���7̾;�1��n��ʟ?)�A?����V�� ��w�������W?>=���� ܬ�ܖ�=�ܲ�q^=A%�>���=���/3��lS�q0?�g?�d��!3��j*>t� �<=]�+?C�?sgU<%�>�=%?�+�,��b[>�z3>$��>���>��>t*���۽>�?��T?|��眾v�>L��R�z���a=�;>��4�gs�A�[>��<�Ԍ���]��䐽��<g(W?ɞ�>��)�+��_��:���3==��x?�?o)�>&yk?��B?���<�g��q�S�� �pxw=L�W?.(i?!�>Ň��'о*����5?e�e?��N>�`h�j����.��S�G&?��n?"^?�y��>u}�������fn6?/�w?�b�)1��G�����j�>���>d�>>�3�7]�>��:?�[(�r8������'4�uf�?�@�1�?�F\��!߼k=8��>Ԧ�>�p6����Y������u�=���>NǾ5mx�H�����u??�_�?�*?)Y��;����=�ؕ��Z�?7�?􄪾gg<���l�,n��nd�<��=�$��i"����{�7�7�ƾ �
�����?��{��>�Y@�]轇,�>i?8��4��RϿ6��b]о�Zq��?��>��ȽƝ��M�j��Ou�!�G���H��v�>�,>/����Y��%|�%<��%����>����-�>�eQ�%޵�5H��� <�ɑ>D�>��>#���ԣ��(ݙ?�E���IοZ���sE���X?By�?o5�?�I?��B<�u�`�{�-����F?9Es?t�Y?�I�d�Z��:�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�nc?L�z���p�к9���T��ۇ>��v�C��.�=���m�t��}��2�h��?g/�?!�?���(��<?�a�>x���X&ȾZ~2=uA�>wW�>��>X�i��>���}7�A��=��?Xc�?�Q?�덿�V����>��y?&˶>AЄ?��=�6?��=����s���Y�>�A>�+���1 ?�mN?���>hm�=MA���)��WH�ȭQ�c� �2�A�ṁ>=�_?M�N?+ya>T	̽��'��Q��N�����'W����3�u����s����>�)4>n�
>�W��yξ�?hp�?�ؿj���r'��44?⸃>[�?�����t�m���;_?~y�>!7��+���%���A�]��?�G�?m�?a�׾K^̼�
>v�>�J�>��Խ����4�����7>��B?��yD��m�o���>���?�@�ծ?�i���?� ������i��W�A������=�tB?#���zA�>��?�o=�}�6���9v���>�>�?���?�H�>�>h?���0C�����m�>M�?"r$?ԡG�pR��#�M>�7Q>D��h$q�����v=o?y��?Y:@��q?>��Y�ؿK���fw��+1ʾ<��=��(>1A>��1�=a>i��=j<���=�\~>`�S>E*>�y>�f�=Q�=� �����֖�5����3�A�����X�J�J+	� ���"�\�ffԾ�����.��o���^���(������>�8O?�[?Իp?���>��$�_I>����	�=I꾽��M>U�>�]9?C9H?�3?�	�=�Ȳ�uu]��Os�!���ܗ����>��)>:�?��>��>4�C�1Ŷ=�ҙ>�v>�=Wx�����bǄ<�H%>�J�>��?��>�C<>��>&ϴ��1��Q�h��
w�c̽�?����@�J��1���9������h�=Eb.?�{>���?пk���}2H?v���?)��+���>n�0?�cW?/�>���6�T��9>��ڦj�`>�+ �;l���)�*%Q>Xl?��q>�Cc>9_Ծ.�L��.�H\��Z�>(9	?Y�ݾ�:��%i���K�W�,�$�=���>������1��0���b�k��,�ЦO?y�>��ڽ�@W��>B��x�E�n>1XF>�ϓ��p=�Y�=�����K���w���ރ=�:>�Q?u,>�#�=�ģ>zV���P�-t�>�;B>�+>��??%?�V������~��,�-���v>O#�>EՀ>��>1^J����=J��>`�a>Eg�J���Ñ�x�?��}W>a�}�{_��t�Yy=�X��&�=D�=�� �W=���%=&�~?/��刿P�#���CgD?!.?*�=��F<�"����P����?G�@�p�?'x	�O�V��?B�?���JA�=�w�>J�>��;}�L�٢?�}ƽe㢾��	�\#��R�?��?&�/��ǋ�>l�B>^%?��Ӿj�>�|�.[�������u��E#=ߣ�>C<H?Q���O�K�=�ku
?p?�a������ȿ�xv����>�?d��?R�m�`B���@�r�>��?�iY?>ei>�d۾ZZ�T��>��@?ER?��>�6��'��?�߶?�?S|R>��?�h?ֱ?�+:�����/��R���Pn>�夽�>�??>1���Hn2��ߒ�f����yl�k���~>�_p=(�>�G3��hȾ^�M=���CJ���<漦ə>ب�>7�>�i�>	�?�>��Z>������Hr�jҭ���J?CĎ?BD��B�O��c�퟽O2����	?��C?�������ى�>3�q?�?��Y?T��>�Y������ö��ȹ������r>u<?�j�>5R���w>
��ЁN���>\߈>��ɽ�r��+D�G� =!(�>&n+?�\?=�=��!?=�'?�=�>���>�@�����I���>4p�>�U?��?��?�B���v#�b
���Q���d���">h�i?+?���>h���`a���F�������ǽʑ�?Z�c?��4?�B�?Q�R?C4E?�C�>��43޾_.��,p>��?Ea���;��Q(�&���^?J�?���>�o���սR#�3w�9V���?�[?#]#?����c�/�ξ"l�<E��QG�<�.<49~��N">]�>�s�����=P>�%�=��k��t=�ʍT<��=n�>�#�=��4��#��@=,?��F�Pۃ�R��=��r�uvD�B�>T8L>���^?t=���{�����w���U�1��?ӡ�?�k�?���[�h��"=?��?.?V�>jM��7޾���9w�5{x�9u�
�>���>ʆl��徱�������E��<�Ž���x�>]��>/�?�E�>��L>��>�o���C'��)�� ��]�Le���5��h)����FȞ��-��+s���þ�$����>=}��7��>�?~�m>�v�>���>��;��>�4X>uv>G%�>UjQ>��3>���=n
l�p�Խ�KR?����	�'���辊���c3B?�qd??1�>1i�%��������?���?Vs�?e=v>�~h��,+�zn?�>�>-��Qq
?R:=�2��;�<�U��O��L3����>�D׽� :��M�Unf�_j
?�/?�����̾=׽z��}j�=�x?��&?���uAW���t���D���I��&���fu��������q������� ����{#�`z�=��-?�8�?F?��˾b��w��6?��Y�>�1�>^)�>���>"�b>�"���/���Q����� g��D�>��{?�1�>�j@?��J?SZ?��8?.j�=�>1v9��f?a��=���>��?DD9?�V-?_@?�?�\�>�
>G�-�����dӾ�}2?��?�7<?��!?e�*?����KV���> -=*0�-q���;��ԽA��:s�=��'>[X?2����8�l���mk>��7?���>���>���#+��g/�<l�>��
?�H�>u  �j}r�hb��V�>~��?b���=@�)>���=�����Ѻ^]�=�����=�4���n;��|<l��=��=�^t�T��t�:���;p�<Y
?�;?�S3>޼>_O)�
����&�Z����?>�I/;y�b� �w=���Ǉ���B���>��?�+�?9`3�-�=X�=��G��Փ����P�����㽍��>Q�F?� ?��y?�6?���>5�
>/��������������F�#?g!,? ��>e��гʾ�񨿧�3�͝?=[?�<a�/���;)��¾�Խ��>�[/�;/~����ID�@�������+��?Ϳ�?A�8�6��x辳����[��X�C?�!�>�X�>M�>d�)�z�g�p%�N1;>Ԋ�>BR?c�>��Q?��v?�GW?�_8>:�A�z2��@���i��<1V >R�A?���?	T�?�tx?n�>�>�I������A��@�@�(����p� 8�=s�b>���>A��>|��>s��=����>˽�H���w=Օl>�F�>s|�>�>���>)v�;�G?���>�\������椾����=��u?$��?
�+?�"=W����E��H���F�>|n�?3��?�6*?��S����=��ּ�߶�|�q��>�ι>�*�>�ߓ=z�F=�c>
�>���>�4��^��o8��|M�!�?F?Ȼ=_�ÿ�I#��iɾ~˥���z>�ԇ�o��ӳ�=ό��o/�����/ѾEսʯ��W�Λ!�7�����&�sa�>H.B>d��<{�]=݀�;kUk�QN���B.>rۅ=�o];-��_=/(��,��<��#��b3��`f���B<L�=8ǾN{?fL?�>*?cC?�!w>d�%>�`�m�>@Q��W?e�g>/!E�=����+�ӫ���B����ھI�ھ| i��!����>�'����>��:>94�=�к9U��=�n�=Xjf=���I�3=Z��=��=�R�=_��=�>#�>�y�?7���K��_��{�dc5?�!�>no>�L=nZ?g�.�_ ~��ݪ��?���]?��@{��?X?ܷ%��>������U>���=I>��A�6>+��>���=M?7�>��\�M��*��="W�?���?��X?c���m��4#�>�8>>�)Q�� 2��Q\��`���U��� ?#L;��˾W�>况=��Q�žtm9=o 5>Z�Z=���vX]�A��=#����O=�ah=$�>I�D>�?�=������= `N=ơ�=MO>�;滘�8���,��17=	2�=�3`>��$>���>�??��/?!d?�v�>�fl��DϾz¾R�>J#�=+-�>�ρ=W\@>���>E�7?��D?3�L?���>7K�=���>��>�,��l�a�>]���:�<D��?w�?H0�>F2G<��B������=��Ľ��?W01?�+?N��>�U�z���X&�g�.�r���+��F+=�lr��TU�����m�.����=Oo�>���>�>�Ry>W�9>��N>��>6�>B�<�s�=sҌ����<j��N��=ꪑ���<��ż�5���O&��+�j����ݍ;q��;��]<}��;ʑ�=�.�>�	>�G�>��=mڳ�2%/>$喾��L����=O_���4B��Bd��~���.�`q6���B>��W>(���U*��L�?/�Z>ȋ>>dZ�?W
u?�� >���nVվ�����d�:�R�^ڷ=�d>ŗ=�f{;��|`���M�i�Ҿy��>�ߎ>�>��l>�,��"?�'�w=���a5�v�>�|��E���)��9q��?������Si��*Һ��D?�F��z��=X"~?O�I?*�?���>]��υؾ�;0>�H����=���(q�>h��o�?B'?���>��+�D�Uħ��C��|�|=�
ཌྷ�L��G����Q�x�>��q�5 �>J|�zj���#E�p ��Bߒ�8r��������>��k?�5�?�Ծ��{kv� �}�!�(�?t�T?���>@�?9�E?M��=�� �,.P�9?�<�P�?�`�?�n�?��>^u�=.������>wV�>� �?ߐ?~�r?�X7����>�'=g�.>�����>�';>JH�=X�=*�?��	?w$?v,w���g���4�.�c�1=���=`~�>�Ӂ>՜T>�ͷ=���<#��=�VA>���>\/�>'an>�ל>��]>)Ԣ�E�
�hc&?4��=ba�>�0?���>y�K=����:��<s���F�O�=�A`���@̽`h�<�8�+�=�aC���>�Iǿ�&�?ߞQ>���?W���*�T��lT>%�U>�2潎u�>��8>�y>5�>d�>=�>��>�+'>�HӾ$�>^���\!�Y"C�5R�&�Ѿ%{z>ښ��f#&�ԣ������OI��y��i��j��+��A8=���<QE�?T]���k���)����K~?�C�>v6?�֌��2��K�>���>i��>�O�����⾍��K���?,��?�߱>���>q&?o��>��e=>�j>B��9���np���Æ�Xfn�g/m�cZk�������76?���?��^?�W�M�c>ca?��@�������>����7���y�KV@>kB������#���7om��&�jһ=��I?�E�?�{/?V�#���s=�?t?�>�>�ޅ?��4?Fk?|�A�I5>��,?�@?��O?�Z?�qv?c?�=7��)��*c>�Gx>&v��"m��Տ�ku��9?s�W,>��=UQx��h���<Ms�=��Z���L=�^>
�T��m꼤��=�=�=#iW>#̮>�ua?���>O�>A3?H��M�=�3�þ��+?�P;�_��D⓾+帾����=F�Y?�?�?�/b?��H>�>��k9��((>���>�v>��o>]��>�7�d["���J=��>��9>���=/@��aw�'|	�hk����;�'>��?lf�>-�n�[�"=������F��Kf>����p� ������Y�\
G����_�?�Lt?r�?�?>r�x-�h�]� k�?��\?/@#?�/�?���=��RNU��d[����Qi�>��=�e9�V��_ǰ�;�k�띒��>!�:�5ߠ��Vb>#��It޾T�n��J���pEM=��}[V=��u�վ�5���=�$
>������ ����֪�o1J?�j=�w���aU��p����>���>�߮>��:���v�[�@�����)6�=ݵ�>R�:>ae������~G�B8�t:�>�RE?	V_?#l�?[���	s���B�a���aS��iKȼn�?B��>k?�B>���=M���}��d�G���>[��>I����G�H3��|/����$�P��>�;?V�>?�?�R?��
?`�`?*?�B?
�>4E������C&?Ȉ�?~؄=2ս�T���8��F���>�)?}�B�:��>��?�?��&?�Q?�?�>?� � J@����>/_�>��W�Ec���(`>��J?���>^4Y?�҃?�
>>�5��뢾��D��=>��2?�3#?9�?3��>��>������=[��>vc?/�?G�o?�j�=!�?(G2>1��>��=���>S��> ?�SO?B�s?��J?|��>�G�<6��!���:s���P�+H�;!�H<3y=���+Et�Ȋ����<�d�;r��ᓀ�\j�ݰD�~����;�9�>��t>�T���2>p�þ˱���WA>B������|��X79�^��=���>-�?�Օ>��#�]=�=�?�>���>����y'?Y?�??U8�yb�apپ�}N�"��>�B?8��=Q�l� "��	xu��rj=�im?�B^?�@V������r_?>Z?�о���7������0��C�x?q�3?��R�5��>�(t?~��?�� ?R#>���\�� ����`�M��%�1>��X>Y��_���ߐ?i�M?�>2��>���=~�ʾ)����)¾�?��?tҦ?�d�?!��=��R��\�����&ُ��0M?���>'����?��J�_��b��i�¾����ા(��}I����j�/��ɔ����3fR>i-?'�v?�w�?ۼH?�Dƾa�k��
M�Y��ek�KX��5���Q���_���:�T�ܳ#����ƃ��]��=êu��@�>�?�<$?�^+� ��>�s���i쾴PؾN>;����K%�te=�v���4a=v�~=qe���(�����E_ ?%"�>���>��9?�X�|T9� �5��X6�!$��9Tk>��>�v�>s�>�vP�Y�T���׽�ȯ��SO� v��v>�c?�xK?�n?=� ��1��y����!��n.�~u����B>,>�>�>W�lQ��&��<>�,�r�8��w����	�J�=]�2?��>ma�>�?�?��?�h	� ��+�w�ԏ1���<�-�>�i?s��>�ņ>a н�� ���>kpZ?��>KH�>/��DE��{1�d�[;�Ͽ>��?j?6/�>��K�Ch:��}��/5����)���X>�po?r��o+s�~;>V)l?�
�������>�A��پ�������1n>�?Jo��?�>9Y̾=4'���r�#D�l�%?H�?�Z����1����>��:?���>���>)�?��t>'PϾ#�=��?��Y?dx4?9?D?@s�>Hy�l5�]q��]!�9<���>�D>u��<���=�Dd��Vf�CK���=�w�=���<�����U�sܼ�Il=��ٻҎ|>�lۿ�EK��iپ���$!�(7
�I򈾟ʳ�0j���-	���������x�o���P'�6V�Nlc������l��x�?�1�?E���&������?������s��>�0r��O}�5Ы��l��s�����Y	��I{!�n�O�Mi��e�O�'?�����ǿﰡ��:ܾ8! ?�A ?7�y?��:�"���8�6� >D�<�,����뾨����οH�����^?���>��/�����>ե�>��X>�Hq>����螾;2�<��?4�-?��>Ǝr�*�ɿc���ä<���?.�@E#A?��&��[��"X=h8�>_
?
�;>#�-�:(�"±����>�I�?���?�S=e�V���td?�ȯ;�UF�+��K+�=��=R�2=	��H�E>�>|���^G�;,ͽ��7>琄>C��%�Y�3|�<�9`>�u̽T����W�?k�e���T���(��R��ٍ=-�f?(?7�;�}q?�&��ڿE�n�{Q?�� @�	�?"�M?ӯo��^�>caFw?�B?٧�>4�,�_�Z���b>��=<�ZE��:��l�X��2�=xc�>)0Z>�W�Y>�Xm��ν�Jt<U��ĿN�!��G�Ϩ9��P9<���Z;������d��仾q�c��p�aה<�V�=�L>��w>'H>+{>��O?�i?���>י>�c���P���ƾ�p;
����*��C���vC�S%˾x����美�
�E��0��D��!=���=7R�k���6� �[�b�?�F���.?�v$>c�ʾ��M���-<�pʾm���ڄ��ॽ�-̾�1� "n�a͟?��A?������V�S��X�T���P�W?�O�ѻ��ꬾ��=����ڠ=�$�>u��=���� 3��~S��7'?�,?�NH�0�>�%:#6ϼC+)?P��>S���Ӣ>ݮ9?�|�;ɢR��^>!�>�>q֠>���=zl���0��&?D�n?�V��dþ�z�>Z���7�����>j]>�yh��h=`P+>��>�����=n��=hE�=��V?+�>P'�N���i��9��:�=*{?�  ?g9�>�)z?~�5?�~J�1pѾ��c�� �t�=�g?��n?Kl�=`�F���p[�[?�CL?mX>)�Q�W
���;�K{�#�,?�^n?4�?I�������䙿z�#�^:?��v?=r�������V�/��C?��(?��>E 5��=->`��?���𧏿�N���H%�Х�?۠@�4�?���=�N&=ۜ�=5$�>	��>��P>�F���9��4#�>y�?'����k�Z��m����s?<��?�v�>S�l�n�Ҿ���=�ٕ��Z�?��?�����Ag<@���l�mn����<�Ϋ=�
�xE"������7���ƾ��
� ����࿼���>@Z@jU�w*�>�C8�S6�TϿ%���[о�Sq�y�?H��>�Ƚ����5�j��Pu�b�G�6�H�����>H�>��>���������{�8r;��흼e�>�+���>�vS��:�������,1<潒>Ҋ�>�ˆ>%����罾}˙?����Hοڪ������X?mk�?�l�?Db?�&9<	yv�w{��C�!G?�~s?EZ?�_#�W]�U�8�~�j?xS��gO`�x~4�9KE���T>�3?�G�>�-�Ns}=�:>��>�T>�/�T�Ŀ�ڶ��������?���?u����>bz�?+?�f�w7��~J��n�*�u�%�x/A?;�1>tx����!�V3=�ᾒ��
?�o0?r��I.�_�_?0�a�P�p���-�e�ƽ�ۡ>��0��e\�wO�����Xe���Ay����?N^�?l�?���� #�h6%?�>N����8ǾM�<���>�(�>**N>�G_���u>����:��h	>���?�~�?Tj?���������U>�}?'�>�߀?^��=��?���=$͝�#=Zۮ<`�E>�������>��Z?Y2?�o�=ƿ�Fs�}�%�Q'@��R�2C��q�>B�e?�?G?��a>�(�i�νj$����=�?��A��.*ܽ2��������6>?�H>�lk=�r��s�ܾW�?����ؿ�i����'��c4?^�>��?���2au��h��f+_?%U�>�X�6$����%(����?�/�?	?:�׾�<ͼ�>��>Ԅ>sս�j�����1
8>8�B?��\C��ϼo�ŀ�>.�?˥@�ɮ?�h��i?�v#������z����*�<ڒ�|.�>
.3?	t#���P< 5?�=����c�YF��D���x4>�͵?(��?��>Ԥ�?�s��<�r����<���>"O�?n2?,Z�W��8�>b}-?>�I���Z�^��9a?8�@@U�X?Ty��I�ؿ�c���i��փ��O3m=�?�=�F�=ouT� ��=��=�ˤ�ݼ�3->�Ü>\�@> cW>��,>y�>C� >͂�eK&��5�������P�*��P� �J%�Dc���y��W��Ө�#���������zyȽk�C���>�;��{��f�i?�Cq?د�?U�.?5Ǻ������r=���>(���Q\�Nq�>Z�I?PM?��?��=�`������|�S}���7��kj�>�P�=�Q�>��>��R>�P���Hm;���=/G�>!�@;1<��@�<�;�=�b=��4>6��>���>�C<>��>@ϴ��1���h��	w��̽&�?'���b�J��1��9��F����i�=b.?�|>����>пS���|2H?6���f)���+���>6�0?�cW?5�>�����T��:>Ϳ�1�j��_>[+ ��l�a�)��%Q>�l?e�W>�5>C�� '&�x�,�ʋ����>��2?�����*^��o��+h�Fq���=� ?-&�=o���ɋ�۷j�]ے� v�<Q�S?y� ?����a̾=0���E��ҘR>�ڂ>>E�=�V>��>6��I���{�4�Ľo��=\��=��?�K>�1S=lx�>y_�������>J�/>��+>�wE?�� ?|P�<�$������A�V�>:�>nӄ>Q/>��h���>C��>G��>U��4ͽ��ӽ)����ǔ>�Dؽ���,%����=Z���Y>��=��+��6>���<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>����Y������u�ٱ#=��>�9H?�_��OP�W�=��p
?:?#g�5�����ȿ�qv����>�?��?�m�ID���@�~w�>��?�lY?bi>e۾�aZ����>T�@?
R?4�>�5�W{'���?�ݶ?��?�yI>��?�	s?��>�΅��Q0��O��88�����=�W�;��><�>,��kF�غ�������j�
���e>�%=�x�>���ev���'�=}4��=�����h�o`�>�<m>xfK>Z�>��?���>y��>��=c���ᓾ�>@?���?��0������� ?�� ?�N���?��L?̚�=���r�>�P\?��?FB?�~�>J�7�Q�����ſ�v���=�=�=�ñ>׆�>*��=�3�=���U��q�*>�>>�=+U��Sy��؏���z>�S?�I�>�:'>�5?_�1?65h>�?6d��O���(�C�>�/?3�	?��x?�$?��y���,�����^䪿Io��c<>�	�?ؑ?�pi>��y��A���X���>�������?`�c?�iQ�eq?�l?mvq?�Y?o��>��ü�o������>��!?!��̼A�N&��F�P�?�T?���>Lֽ�ۼC�������?=+\?�K&?2}�a��þ���<,����K�>c<-^F�g>�>�臽�=�>س�=}�l�E*6���^<���=��>�.�=��7�q��7+?
j���t��E	�=�>m��@�	}�>��M>�$Ǿ�oY?��I�q(�N�������;�呍?o��?×�?������h��<?Y��?@�?:��>v7���C׾��ݾQ�^�r�G�{>ш�>.�ּO`�p��.C��������۽�2����>$�>�h?B ?<N>��>�A��~V'�L5����L_����[�8�\j-����f.����#�l��¾(�z�/�>)��a�>��	?_g>`�z>�W�>>���&�>�OS>�>PV�>$U>	U2>�(�=gI<D�ҽGR?������'���辴���	3B?4fd?�1�>��i����������?���?dn�?�Fv>�vh��$+�
e?�1�>���Y
?l�:=��
���<�a��]�����}b�fю>S�ֽ�":�MM�ff��o
? ?���j̾�׽���0����?'o?�0�.`_�Y�aO`�w`���ļI밾�ξ)]5�׏o�"������l���$�9�p>`N2?gXn?�l��� � CZ���k�j�
����>��q>��>��>P� >�������l�5��n�u�>rW?a�>7+G?3'?<�Y?�1@?T��>~�>��¾��>#b_=F�>l�?��N?`%?��)?v	?��?t�'>�(�
���!���[$?_i?e��>�]�>���>Y�̾Z�=�
*�a���	e���f��`�=L��;�I��L�,a����=�X?���1�8�{���
k>��7?�z�>{��>U��l-����<�>��
?�G�>�  ��{r�c��S�>;��?��π=Z�)>p �=X�����Ӻ�\�=T�����=hi��br;�؀<���=��=.�t������:�_�;��<��?ؗ�>5��>��r>�O����	�_���^.7>�m>�u+?��Z>������!̆��y�x�g>�
�?CV�?�/�=SA>��>���-[���d����p�i=A6?�	A?�C??6�?]%<?�0*?lG�>�t.�hޜ�&p�-�3�(�*?�,?���>����ʾ�먿h�3�?�?�Z?�:a����;)��¾q+ս��>YN/�f#~����VD�YЈ����=������?���?�3A���6�܀�\����g����C?�!�>h�>��>ѿ)���g�!�81;>���>
R?�׻>��O?bI{?V�[?#U>��8����ә�٧��R!>��??���?���?�y?���>��>��)����r���� �_�򽉋��{�V=19Z>�^�>���>ܺ�>{��=��ǽ�쯽��?�QG�=��b>=��>�J�>j��>��v>h�<t�G?��>���q���餾�ԃ�8=�؉u?���?#�+?�=f����E�*b����>�g�?^��?�I*?3�S�K�= mԼ�Ѷ�µq����>[ù>���>�S�=$�I=�>|�>X��>�9��F���8�˲M�}?A=F?U	�=wƿ�q�9HJ����?�T�y���L�h��G�qg� ��=������{��>�j����R~���ù�����V�z� ?��q=}U>qڮ= |�<G� �/(=�FZ= @<�|�<�Ӈ��ى<ьX�
7�44��p�R�"DH< א=��F<yBϾz�{?C�O?]�3?:wI?�s>)��=����7�>���^P?��u>3�ڼ0(��9F9�������)_�^�ݾ81q��Z����>a3X�I�=S2>��">E<���=Ab=�r�=��U;Ԅ�<��=�=�=�G�=�X�=#�K>�
8> b|?m���=�����U��*�=�G? �>s�>p���JM?�=�>����P���Ս�M*�?>\�?���?�C?+/ɽ'�>�H���nD���@=���;<!���<�Œ= )'>��g>�S�Z[����ƽ'�?��@֒D?��{�:�ɿ�KB>�8>��>��R��q1�9I[���a�^�W��|!?`P;��R̾1�>㷵=Y�߾&�ƾ=M6=ɥ7>K�c=~��o\����=��w�A�>=x_m=bo�>�B>bS�=����{ع=aJ=}n�=%�O>�(���;�)/�`-=D�=r0a>��$>��>�?|g1?��c?��>5Do��Nξ�~��[��><N�=��>��=q�=>���>=�6?��D?�+L?=�>��=	�>�u�>��+�F�l����J�����<�k�?%�?a�>%t<�cA�j���q=�CҽQ�?S�2?(7
?*��>Ub��W˿b�N
���ܩ�\�9����]��O%=p�+�������˔�>�I>�ơ>@>�Y
>N�=A|>h;�> �Y=]���9!�=\v��fɶ=�(.=�1��)6�<|q��|�֜��{v��>��V=� �<y�7�m�=�m�=p)�=���>\>*D�>M.�=�;����3>����'M���=\��EC��d�E~�P<-���2�qDD>M�V>���4#���?�tY>��>>���?*Wt?�!>���	�Ҿ������e�AR�#��=��>�P>��;� a�g�M��ӾD�>�a�>$��>`2s>ۋ,�;@��=f�߾�t4�Bc�>�㉾f�
����Cp�B���;���ah���3:�D?R��!��=j�|?�J?/�?)�>ZN��v	ھ��2>�;���}�<���+�o��[��p-?��%?� �>���vD���Ѿ�Q�1/?׀�_�/�>|���a�5���:<�rcA>����v󾶺<�E����V���pK�{+E��`�>K(J?[�??vm�e�����R�I�%��<�=��>�?�h�>�ѱ>v�8?�^�ø�`���I�;��P?%D�?r�?�^�����=�˴�Q �>v0	?���?��?�}s?�j?�	]�>h4�;]� >�b��f��=�>缜=�	�=p?�
?e�
?j����	����6��R^���<�I�=�W�>�x�>e�r>���=a�f=	��=@(\>�ޞ>ޏ>��d>��>�G�>�����	��./?��=��>a�?���>ٲM=��0���C=�Ͷ��5u�DX������c��Z=�񚼥�=F����5�>�ʿ�Ne�?�]>��� 	?j 	��Gͽ��=�i�>�И���>],>��5>V.5>�s�>��v>=r�>9>�PӾ�g>H��a!�*(C�0�R���Ѿ]z>����H�%�ʡ����=XI�uv���n�oj�.���:=���<�F�?����-�k�j�)�������?�a�>�6?�ٌ�I����>���>ˍ>"J��5���ƍ�^_���?���?��g>��>X�]?ܢ?3p2��=���S�P�o�mD�j�S��]������Ӂ�U9�C̽~�]?��x?2�C?�<<u�>�s}?��q��"V~>��*���>�3 r=l��> ���A�M�[Ͼ��ƾ�?�>�j?T��?@�$?��?�9�m�K*>UY:?TD2?3t?gA1?��:?����$?��3>��?i�?��5?�.?9?�0>�2�=��	�؅=D㕽�Ŋ��t˽ 9˽������2=�{=�_����C<
�=]��<�V��;���9@;=�R�<}�8=<��=�5�=q��>��]?�6�>Y��>?�7?K��zx8����:&/?&X9=ܮ��������_���>{�j?���?XZ?$Pd>��A�9C� >j�>(c&>@�[>	q�>���еE��
�=Z\>�Y>Dݥ=d~M��Á���	��~��/�<K1>���>g�%>轂��=�Bv��E_����>2x۽\2��Uc��8�G���T�G��ވ>��c?�/?5�C>K�˾�l5���f��@+?n)?��1?n�r?Y_�=�߬�}qB�[$�$�*�NDB>�cb=̙
�����J��F������ >�㶾>ߠ�OWb>ý�Xt޾G�n��J���羞HM=@�� XV=����վ�6�٠�=8#
>~���� �-��z֪�r1J?ګj=�w���bU�p����>ſ�>G߮>2�:���v��@�篬�5�=��>��:>~t����~G�08�~5�>�ZE?K_?�r�?�����r�)�B�W���jh����ɼp�?8��>�o?d�A>�=�����W�d��G���>��>���W�G�����"���$�-��>B+?3~>8�?k�R?��
?�`?*?U=?��>����}���B&?3��?�=��Խ��T�V 9�1F����>��)?n�B�ȹ�>B�?�?�&?�Q?ŵ?��>� ��C@����>�Y�>��W��b����_>��J?A��>B=Y?�ԃ?��=>J�5��颾Yש�.U�=
>��2?�5#?=�?���>B��>�����=��>�c?�0�?.�o?���=8�?�92>���>2��=盟>R��>�?DXO?�s?��J?ߑ�>ܹ�<�7���8���Bs���O����;�yH<��y=����3t�eL���<��;�d��`H�������D�1�����;oZ�>#�s>���0>n�ľ�6����@>uY��~N����V�:�.��=Uf�>u�?ͱ�>kD#���=���>F�>+���(?%�?U?J;Νb��۾��K����>o�A?��=��l�˄����u���f=!�m?.�^??.W�e���y(k?�H?����t�=�^_��(���i�?2�?��X����>Q`?ǵ�?�m-?�=�����5u����9���̾�X>���>#,�\����n?P�C?��>º�>��X>�X,�"�\�w�XL?;��?*�?�-�?x&>��W�Ql�D���"��B6_?>�>o!����>�Ͻ�+Ǿ����ŕ�ϲ����uH������a���$�a���_�#���G>?�?ک�?R(}?��L?n���F�h���C��[�B�~�� ���&���C�_�G�HNI�����$������]ʙ=~��uA�}�?��'?p/����>!N���s��̾��C>�ȟ����e�=�$��TA=��Y=��g�9.�y̭�� ?�G�>�4�>��<?��[�*>�$�1��7�4
���3>��>ޓ>zz�>)A��.�.��[Ⱦ�Ճ�?iн5v>fzc?�K?��n?Ib�W(1����l�!�e�/�g����B>x>R��>��W�<��9&��X>���r����`w��~�	���~=l�2?X'�>D��>SN�?W?�y	�2h���kx�*�1�ٚ�<�/�>�i?g>�>&�>�нG� ��!�>�J:?fO?g��>��;L��$��Ñ�s?�}K?+̈́>8�>T����7V�R����� $�9y�>>�l?�$��Q���	�>��>?��=N�=9A�>��<��9�����h���iQ>L	?4G>�>Ę��s���p�4d$�vF)?�g?y}��ט*��>�:"?��>�h�>��?��>$þj&��?<�^?{(J?�A?���>=�����Ƚ='��.=�ˇ>��[>xNl=���=����\����)�E=���=GRԼ���t�<�C����S<���<�A5>KMۿ�#K�Nl־ɻ�%o�cR
�h����2���,���	�C����:���y�r�݁/�V�U���d�B��kmf�.��?\j�?�ː�����8������#�����>��|������.�����᝗�K��	䰾D"���O�5�i�WOd�H�'?�����ǿ簡��:ܾ6! ?�A ?!�y?���"���8�ȭ >�B�<�*��r�뾠�����οP�����^?~��>��.��c��>��>�X>VHq>����螾M1�<��?E�-?��>��r�'�ɿS���lä<���?,�@nzA?�(�8�쾴/V=@��>e�	?��?> 	1�bK�s���`�>�<�?6��?x�M=��W�I�	��_e?��<G�>;⻻��=^M�=X�=���7cJ>�^�>a���A�+ܽo�4>Յ>��"�^���l^�Hż<�q]>c�ս�=���?�a�xr�M�I�XP��,>�+?U�>W�����>��g��Qӿ"�ᬎ?�@���?d�'?.7Ծ�¼>�~ݾ`�X?�C1?d#x>�3F���a�ſ�>+߂<p`H����Ao���>h
�>6$����r���bP��N�$u(>�� �nĿr��nw����<L|����ӽ�����m�h0��ʔ��wX�K{���S�<���=�K>Mlp>1�S>d^~>8�T?I�w?<(�>�,;>,�ý�Ȅ�_xľQ�::���b�[J��.�	���"C���`�@��m��£�!=���=7R�p���C� �f�b�S�F���.?w$>e�ʾ��M���-<}pʾY���܄�᥽�-̾�1�-"n�k͟?��A?������V�Q���W�̄��T�W?,P�ӻ��ꬾ���=����2�=%�>芢=���� 3��~S�://?�o$?;پ�����k>a���ɉ��q1,?��>E}�??�>�!,?)��FȽN�X>��>	��>���>#�=k��������?��`?����Ȟ�AQ�>��ʾߪ��3�=��=��7��୼Q�+>~��<I\���u���d��w4�=>(W?i��>�)��� g����ON==ȯx?�?S6�>�yk?��B?��<j��9�S� �Cfw=��W?�)i?ƶ>����оM|��s�5?i�e?m�N>�hh����O�.��T�4&?j�n?^_?�����v}�R��'���n6?��v?�s^��s�������V��F�>�]�>ܿ�>k�9��k�>n�>?�#��G������W4��Þ?��@���?Q5<<��C��=�6?N_�>˟O��4ƾ瘳�V����}q=!�>*����dv�`���I,���8?`��?��>�������¢�=�ؕ��Z�?��?D���k�f<���l��i��]�<׸�==���R"�&����7���ƾ9�
�'����������>Y@�W�p$�>�D8��4⿗SϿ����[о�Xq���?=��>��ȽΚ����j��Ou�1�G�@�H�����]�>/�>�j��K䑾)�{�]m;��#��Y%�>��%�>��S�W��gu���N6<���>1u�>��>�Ӯ�Cн��ę?/I��<Cο!������Y�X?�g�?�|�?ya?��2<ϐv���{��y�`DG?��s?IZ?�p%�U/]�`�9�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�j�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�+�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�F�f?��p�F.���+����<���>'H�������CP�:�;�����9l���V�?�K@� �?c���%��"
?ͨ>��V�|���w�ҽ��K>G��=��>��=B��>+"���g��vv�q�?�J�?E?/E���w��t�2>̘|?÷�>��?�{B���>?y�>�g���=Qe������N�q
?e1d?�d?�~�<��q���M�<�w ��6���2�y��>��_?&g?"�@=���:J�;2�>�#�[���%�O������>�=�xJ���>�>7L4>y,G��yI���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�܃ ?x	�ph��'���6�������Ȯ>�f+?��rr>��"?�v��1u�~2����i�j�>���?�%�?���>�c�?ۇ�L�����<(�}>7ǫ?o��>}����qվ�?J>\�>?S��d��e��M.}?�W@ȱ
@�qS?q��Ahֿ�.��Ɔ�M�վ���G?ݽ�䴼o1޻�_�=�=�v�8Q�0<6=8=d"d>"(>�9\>�p> �&>x9>>�Y��hS%�aj������%�_�FR*�-��A9�S.��#�9���˾�Ǿh
��/�<�I嶽�q��Tk�wM���=�_?y�J?{?}
?3Z'���=O�	��F�<bR�ZO�=9£>�58?�JC?��#?��}=K����f���}�V5��>�y����>�>S�>�I�>�<�>��<k>#�?>��[>�Э=nY=),�;��6<��?>՜>f$�>�{�>D<>��>ϴ�y1�� �h�	w�_̽�?͂����J��1��T;������Tj�=�b.? |>r��!?п+����1H?/���p)�)�+���>#�0?<cW?��>Y����T�;=>���B�j�_>�, �=�l���)��%Q>k?OAn>�9w>�=�����+��_��A?��-?�ھB0K���s�
�d��1���p�>�?	E�5����u��w��ُ�=�l*?�ջ>��>rTn����ϴ���>�ި>��>`7>'HE>`༂�?�Xf� ����ك>Ÿ6>j�?qd*>�s�=_�>M���A�R��>�Q9>�!3>C?!?^�ܼ���������-8��9g>��>��>�B>�dL���=3X�>x�^>Е�I��6J�r�3�m:M>�����a�P�f� ��=�⚽7��=���=m��r�@���%=.�~?���0䈿`뾑c���lD?�*?.�=#�F<V�"�+ ��)J����?s�@Ym�?ǁ	�0�V���?�@�?��ٺ�=7}�>�ի>ξ��L�L�?��Ž�Ƣ��	�+,#�`S�?��?E�/�*ʋ��l��5>�^%?��Ӿ�h�>�w�Z��%��&�u�=�#=��>9H?wU����O��>�w
?:?�]�⩤���ȿq|v����>��?���?��m��A���@�؂�>���?�gY?8ui>h۾�cZ�Ҍ�>��@?�	R?��>�8���'��?�޶?쮅?%�I>��?4�t?8��>}��۲.�F˱����ᖊ=�<�>�>[|>a����F��̓��+���3i��`��hj>�*=���>��`ݾ�a`�=�������=6�E�>��f>d�N>Q��>}�?���>�=�>��<�>�����1閾�Q?Gِ?��>���o��s>[c�>(	�{J?slD?A�%��*�	��>M�i?�|�?B  ?��^>O�D�^`�Zd߿̠�� -�=y�;p�?%V?��Glt���&̾��'>��>�V�>ٞ�l1���z�=��>*?��>۔V>E|?��?���>V��>��l�����5)���>���>n�2?�wK?�#?�8q��
&����}e���c��Qg>��j?�K.?�>c���x-��۝��:尹S@'�D@�?/?.P��)�2?�GJ?]�?�h?w�[>���w������څ��� ?�
��AB���#�޽�m�?��?J��>1���ɽO�0�j9����d?��]?�#?�v���d�Hcƾvk�<�Ň;�(�6K�;�㹀�>��>=
��Y�=C.>OA�=��g�k�5���]<�P�=:s�>	��=4X-�u���2>,?W7I��i��ќ�=� s��D�!@>�K>;)��<_?�d=�W�{�����x����U��܍?���?�u�?c�����h��=?%	�?L(?,��>(���v޾��u�w�F�w�]W�f(>���>Лd���늤�����B���:Ž9�����>>$�>30?.* ?O>���>M����&�*�� ��7z^�	q��k8���.�^��й����"��M�b)¾��{��>�>j���!�>z�
?�g>��{>4��>#l�6�>#5R>j�>D�>��W>�[4>|� >��<K'нNV?���� g)�� �U����A?L0b?��?t�<�����_�vb?uD�?�Ý?G`O>#�h��X0�xk�><��>��z��?
=^�H�钜=]*��4͂�8׽4A�<�#�>Ut��r4��M��Ɂ��9?j?����t�ľ�o)��߾�Oy=�B�?2~�>���q�"^��<��m{�:�R���ž����VS$��s��]��J"��=�ܮ7��	,>ȩ3?6��?�겾&��
N� �`�s7
��w�=�u�>��>�1�>���=!�����-Z��fG��:i�m��>B�m?aG�>;�I?O�;?��P?8sL?��>w��>����(#�>��;�D�>�g�>b�9?K�-?I0?�X?�1+?Mub>z������k7ؾ�?��?K2?f�?�a?o�:ýA���fo�Xmy��À��̂=�-�<�%׽�
u���P=ͪS>�X?���ŭ8�����d	k>)�7?�~�>2��>���-��2(�<i�>��
?CF�>����s}r��c�U�>��? ���=`�)>��=�ۅ�.Ӻ�k�=� ¼w�=4���8;��(<~��=*�=�Ft�z��Ը�:e��;t��<�4?�[�>�s�>�a>+��q%�����>z�?s�?f#��p�Ѿ����J��H�f�M�>��?+�?Q=>�ͫ=s�q>D�����wP5�.��FW��v/�>��8?c�?�=�?�Ã?#�?D�>!�-����9���E�e�B��>Q ,?#��>F���ʾN憎��3�e�?�Y?s:a�Y���;)���¾ սӹ>�W/�<-~�n��bD�q����������K��?'��?k�@���6��z�����tU��ΒC?" �>4^�>O�>��)�;�g��#��3;>���>�R?8��>#ZP?��z?TK\?¥V>38�	���陿+�G���>�@?�ہ?���?�{x?�@�>jP>>j*��ྫྷ���$!����q偾UwR=ϣZ>�D�>�>�ɩ>�I�=h�ǽ�i���?����=�c>Һ�>�%�>�!�>iu>
[�<=�G?��>���A�W奾����5@�-�t?]�?�+?F��<����F��f��y��>f��?���?�+?�qO����=זҼ�@����r��T�>���>�6�>�*�=W�l=��>���>���>
�������8�S�M�.�?�hF?�H�=Aҿf%��?�'������+�ɾ騾8����!���;=�À�p��%��{eh��u��뀾Eά��΍��0���> ���~>Ϟ�=t?x=�/.=�(f=�
��M=ac�=aӽ���`Y��s���EX��q��ɿ3<��=e]�=�_��Zk�?��%?��p?�l?QPs>c"}�:�ƾ��Q>ȴ��yF?�z?_�>J@��dd⽽�V�*	��5��,�Ҿ�q��9��G�>�Ѐ��+>�1�=%�5>8R�=� &>PƱ=`�>}��=dͽp"�=5=���=o�!>��=ۂc>ܜu?����[h���I��R=B;�?2}
>�a��H�2�'?�z?v��w�����?JJ�?��?V?�%����>�c¾_�[���p>�@ >y��=ך������>�>L�&�<���:�8��?f@��0?�'��QR߿IOZ��Q8>��>�
S��21��AZ�a�@Z�s�!?QM;�:b̾�&�>	�=H�޾K�ž�$2=�6>��]=j���\��ۗ=��{��s<=@�s=x5�>^)C>���=����:��=HvL=ik�=��O>�䠻��;��-��.=���=�*c>�'>�	�>��?-�2?��`?�[�>��l��wϾ�Lþ�@�>iQ�=�_�>�sP=p(>nl�>q4?v$G?��Q?O��>��=�w�>�?�>G8*���j���n[�����<�u�?zu�?��>��w��RJ�& ��A�D��C?0�2?�K?�j�>��	���׿�g��8�*���R�{`�(��?��S$>�5O=���`[ý+E�=��$>;�?>�c>�9�=&x8>�Ə>-{�>�� >>�k<�'e���z=�"�=_�^kR;d��<�ظ=����U=�==F��Z=>�<�4W;��=�c�=C��=G �>�)>���>-І=Dq��|3>�^��i�J����=�n��
c@�3/d���}��/���:�xC>�[>e�t�^呿�2?]eZ>=0@>D�?�t?�h!>e��׾����סh�lQ�/�=�f>��:��;�Q�_���M�QѾ%��>J��>���>h�m>Nf,�&?�$8{=!��9�4�Lu�>����p[���#q��@�� ꟿ��h��v�^�D?W6����=h�}?��I?V֏?���>�_���ؾ�[.>X���	=6��q�p�J4��r�?�&?� �>�V�lD��^ᾎ��?����	�!�Tu
�]ж�Uz�0
�>�H���?Ҿv�7��L���]Wi�#�-��>fy?°?3���Dy��J�q���Kߟ= i?I<c?���>�i?|03?��ԧ�<9���d>��?�h�?v��?~��=��=���:�>�+	?7��?��?�s??�?��y�>!(�;� >f����N�=��>%��=,�=�r?
�
?.�
?j����	����Z��3^�9��<y͡=���>0m�>G�r><��=��g=Zw�=�.\>H؞>U�>T�d>��>�Q�>�ъ��,�+�?�G�=ˤ�>�}1?���>�F�����T��=����|�[L_�\�ļ꒬�c��<�>2<��<��ȼ/	�>&|ƿ��?h�g>�� �  ?2J�9S8���>�9%>;�ս�?5LS=к�=��:>跹>�Ϡ>W��>PƟ>��Ӿ�w>�@��j!���B���R���ѾF�y>څ��e '�����-����I�η�����[j�>/��LN=��4�<�>�?��$dk��)�����;Y?��>��5?�����1���b>��>�o�>d����f������r���?p��?���>Ul7>/(i?BY?��.�O��I�&<x��B2�@0��l�'���`��ݠ��X���f?ׁ�?w�I?���=��>�`H?�@���r�2���U<�3O0�Pʆ>
s�>w�������'�lGᾈy���]��D�x?�n�?XR4?�LȽ���9��>�� ?y�S?y�z?�?�>tV?Sx��>Z?���q?�&?�S?>�?��>��j>[j�=��^��j�=����L^���$u�}W��M���ꆽ� �=t�<�>ȷ�<�AD�,{c����=[� >k#�<�m�;��к�j�<P��=���>�]?O�>���>��7?����t8�jɮ�_,/?�&:=m�������ˢ�5��>u�j?���?�dZ?�gd>��A��C��>�Z�>.w&>�\>�e�>�r���E��̇=2C>�\>�˥=�[M�8́��	�������<�)>���>�Q8>�f���=᡾��?�VR�>�����־�n�P�l��L�Z=����>k�c?]!?Sf�=�����1���i��s6?*?��Y?�j?�L�=��x�F�IL�j���A[�>5ݺ<�!����>����JH��qv��,>��Sߠ��Vb>!��gt޾W�n��J�6���EM=���^V=s�%�վ�5�k��=&$
>����� ����֪�d1J?�j=�w��RaU��p����>���>n߮>b�:�m�v�`�@�̯���6�=��><�:>�a��N��G�!8�>�>�QE?jV_?4k�?^!���s�)�B�����b���ȼO�?"y�>+h?9B>��=)������d��G���>̠�>}����G��:��/��]�$����>�9?Y�>X�?b�R?��
?4�`?�*?�D?�&�>������� B&?6��?��=��Խ�T�� 9�KF����>|�)?!�B�޹�>P�?�?��&?
�Q?�?{�>� ��C@����>�Y�>��W��b��?�_>��J?ך�>q=Y?�ԃ?z�=>]�5��颾�֩��U�=�>��2?6#?N�?�>۩�>������=%��>�	c?z0�?��o?1��=��?{92>���>���=���>r��>y?�XO?��s?��J?��>cʍ<�:��`6���;s�cP�/-�;z�H<��y=A���&t�2@����<mu�;.���'��ݚ񼀱D�����"��;_��>�Y>����P]3>C�ɾO-v���\>`&ۼi������hU�"N�=P��>Y�?�)�>�����=��>b�>)q��&?���>�?A�j�|�^�yS¾��+���>�K??B.�=(dr�����el}�Őw=r:k?�Z?+�Q�w�g?0�Q?d!%�Cee�7)���WZ���?�,?��۾$M?2[�?A�W?�K�>��k�ft�����S2I�T�kU�=�L�>a��NMT�|�>��?�����x>�>v�νe�D�	������>IH\?�,�?��?X)>;q�A����'�~�W�Q?qe�>M�o��>�?����Ҿ�u������?����V��~ɾ �¾얾������������>Z<?�n?g.�?�@?ZI���X��
?�VE��������dF���H�]�E�V�]��놿�a�1��!x�{B�=��~�oYA�f��?�'?��0�k^�>.A���)��;��A>�h�����>�=�ꏽ\H<=0�^=��e��#,�c��� ?ƹ>���>�<?u5[�T�=�.1��'7��p��N�4>�G�>��>=��>�ƌ:��+�j��Ⱦ�&���Yҽ�!v>�{c?�K?��n?I��$1�������!�?"/��]��3�B>�{>��>}�W�Ψ��7&��V>�F�r����v���	�ѳ~=�2?W-�>���>�M�?�?C|	��j��Kkx���1�T�<�+�>3i?B1�>A݆>��ϽZ� �\��>�l?���>L�>����FZ!���{���ʽ0%�>k�>Z��>,�o>��,�N#\��j��+����9�q�=�h?U�����`���>�R?�Ї:O�G<�|�><�v�`�!�I����'�{�>�|?W��=�;>�ž�$��{��5���G)?�B?P㒾ե*�~>�"?Υ�>6,�>�#�?+�>!sþ��q���?�^?�@J?�AA?Y+�>|�=`m��&;ȽZ�&�fy-=凇>�Z>��l=v�=V��(\��{��E=���=�ͼ���m<���%�M<���<��3>�ۿ��J��-پ(g�Z �
�
�������)��e���մ��Θ��y����v��_V��d��B��eBj�VI�?"��?Yc��ޠ��޻���^��4g��Hʹ>Lsy��Ê�U���{��і�O��m���* ��N��h�sd�J�'?�����ǿﰡ��:ܾ1! ?�A ?,�y?��6�"���8��� >�C�<�,����뾫����ο?�����^?���>��//��p��>ݥ�>�X>}Hq>����螾1�<��?8�-?��>��r�,�ɿ\���]Ĥ<���?)�@�zA?e�(��쾃V=���>.�	?+�?>�1�;O�簾�h�>�=�?���?��M=ٺW��4
��le?݁<G�����&�=�F�=��=E��iJ>�j�>���wA�x͙ܽ4>kӅ>��"�$����^�2ڽ<"�]>��սs��|��?��[�V�k�'���$��=7�V?���>�&�=+?
eF���οDY^���X?E��?�s�?�(4?�Ұ�N�>�H׾�D?�x-?p��>�g/��-{�P�=.?��y�</'ؾ�M���@=T�>h�=Q{A����fGL�=A�;4��=��(|Ŀ�a#���e��<�J����l��"ؽ�I���q���x��Sg�N��M=[��=-LK>��>|�Q>�[>zOY?�wm?��>�!>��ν���E�;O������W.�����p!(������j�侙x��|�a��{ľ"!=���=7R�n���A� �m�b�O�F���.?w$>W�ʾ��M��-<�pʾ`���sۄ�
᥽�-̾�1�"n�f͟?��A?������V�J��X�����C�W?GP�Ի��ꬾ���=~��� �=�$�>��=���� 3��~S��0?*x ?	�Ǿ�v���;>�� �Y��<p�-?�1�>5�<�N�>_�(?BW*��ٽB`>�(>F��>���>xi�=l0��<qѽ��?��Y?��,��]�>�����Rs=���=0���ލT>��^<�z���h�tZ��#wQ=b�`? ��>aa6���"�{�O��=���>�8�?���>s��=�g�?D}Z?�ok>cJ�:��`�L�˟�<�?X\C?Q%�=���iD�A�w�T?lfX?8��=��5�;td��ډ�t��i�+?>S?��1?1�r��և�?ܱ���;���d?��v?s^��r��*����V�<�>�\�>��>�9��k�>R�>?K#��G������QX4�PÞ?��@6��?��;<"!�%��=*;?�\�>�O��?ƾ�|�����o�q=("�>����5ev�G��qS,�F�8?���?c��>����L��=�ٕ��Z�?��?2���\5g<���Bl�Hn�����<Cɫ=*�a"�W��c�7���ƾӺ
���������>	Z@�O轤+�>?8�)5�SϿ���xZоsRq�;�?�>��Ƚl����j��Ou���G�G�H������>-��!:Z>́��c�i���H��o<߀�>���><�?+���?˾�D���>ܔ�>ر�>B�<Q�9�䀩?f���U����l�1���?|k�?i��?�s?~�J>W��<.���56Y�a�W?��?�p?sv4<�D���^���j?�$��hr`���4��E��U>�,3?��>�Y-��s=%>l��>��>��.�f�Ŀ����PX��nަ?k}�?�5��>]�?3#+?�7��'�������p*�̎��1A?��1>%�����!���<�W���7�
?P�/?r���M��"b?�xz�R�}�Z�B�� �/�"?Z�d��&̾����>½<�2R���V���	�?�@�A�?�z�h澔q?-��>��$�wCɾ�y�=t�>�4>3X׻�52<���>��<bJ�*!�=�o�?�Q@���>�靿bB��؀�>tzP?>��>���?�h�͢*?�B�>�rw���0�:"�>g؅���t<�2!?�Po?��>�t&=���YQ��A@���f��1B�Ӣ4�gB�>�KK?uH?{�=��<�kT��+(�s->��Յ	�����T��<f���Ⱥ,�=Ij=Wl־~X�<��?Kp�9�ؿ j��p'��54?1��>�?����t�2���;_?Qz�>�6� ,���%���B�_��?�G�?=�?��׾�R̼�><�>�I�>^�Խ����Z�����7>/�B?_��D��r�o���>���?�@�ծ?ki��	?���N���_~�<��7�Z��=��7?3��z>.��>��=snv�����c�s�[��>�B�?;{�?l��>|�l?{�o��B�F�1=�J�>�k?�r?��m���Q�B>M�?��a����J�"!f?��
@?u@)�^?q��BϿ���+�����z�g<�ս~97>��!9�=P�8>��fj.=K$`=�<A>�S>�.>�'>W�a>-�$>�}��,��R��8��t�ʌ;��0߾������~�2��+�/Ց�����F轸����P��z���v�����=�hV?��P?��p?�� ?�(p��>�2���=�%��"�=}�>B'2?n�K?��)?@�=Kƞ�X�e�eF��򬧾-K��I�>ſF>��>�C�>G��>݌��ݫJ>O9>:�><�>d==++��F=�vL>fu�>P��>�V�>�C<>��>Fϴ��1��g�h��
w��̽1�?���Q�J��1���9��Ѧ���h�=Gb.?|>���?пg����2H?#���y)��+���>{�0?�cW?�>%��[�T�0:>5����j�4`>�+ �{l���)��%Q>tl?��a>�Nl>7�/���7�N�g֦��і>��3?U����g?�Br�|<I�4Ҿ��K>,��>9P񼑕�nU��#Fm��}h���=�X<?� ?�b������ⅾ12���`n>�O>�YF=΃�=T>|!��ҽ2P���y=��=�EE>U�?�>��	>@~�>tc���O�ڇ�>ln(>�n>uh7?L?��]���]���-4�za�>���>� �>��=�QY��J>��>�z>��p6�"Z��$��+�Bv>�i�H�?���]� ~�=�[ܽ�o�=�O�=��ڽ�'��y=e��?�ؠ��K��:��������u?�x?�)q��j�H	��򠿐����?�@-��?2þ�hR��?��}?ׄG�,�h>�?1��>F�T�����;?��>�$�q9��@}�Q(�?��?6YP=�Q��Jxe�k�=<�>> ڽ�h�>x�_Z��v����u��#=ک�>9H?�V����O��>��v
?�?_�ߩ����ȿ�{v����>�?���?#�m��A��@����>��?�gY?:pi>�g۾�`Z�_��>��@?�R?t�>�9��'�&�?�޶?���?��H>�?<�s?�>��v��T/�c7������-j�=	�X;f�>7k>l����]F��ԓ�Pb��g�j������a>��$=8��>�低+�� �=�!��aC��~�f����>ZFq>�I>n@�>�� ?�Z�>)��>��=�U��)ʀ�����|iL?ra�?O�:�v���7��>S��=��᾵�4?�y?��<�����{�>�K?BR?�??�/>>��&�k���=dܿK��f�=ܩ>mF(?�@�>���-`�>$���� ����>n�I>!��=�(��T;���Q=ً>c�2?���>�}*�u� ?ʁ#?��j>���>	�E����=E�r��>��>o�?O�~?��?7�����3�����ɡ�m�Z���P>wrx??b?���>���������!���D��l��
��?�f?n��.�?�K�?��??7�A?�7c>e�vؾ�A��Uv�>�{ ?�y��@��o&������?8�
?���>b��>ܽ�7�_�6�����?��[?�3#?Qe�*�^�M������<_�ֻ�h;��;�;��A>Z�>�^��;��=�'>I��=%d�BP3�C Q<�3�=#�>���=5�;�s��[�*?!�~^�~��>u���w\9��oh>��3>���e@?䀾��r�����n���H���?�(�?�z�?c��KpW���I?�xv?r�1?�S?Fd0���������Y4����8�>z{�>���~���C���;�a��(#���Cn�>v/�>�1?�e�>;C>w�>�O����*�����.�e(^������6�F*�3;�
��	�����8]u���w����>p�|�Zw�>�?��W>&�k>W��>dc�:�ۇ>]4T>��~>�)�>$V>8�/>�Z>�`<�)ڽ�K?u�ž���>�ʾv��??O�?�Ͽ>l~��.�v�MU� ��>B�?��?���>�mF��.��?GRK?%�����%?��=[�
���=�Ӫ��=���=C�|�!�>���L�+r���S!�m��>���>:Wh�im˾*㍼���Dgf=!چ?�%?�s'���U�\7m�'�Z���T�qS���c��p����'�g�s����͒���`��ͪ"���R=z.?ޅ?��_��x��� h��-8��	R>�t�>���>���>ql:>;��n�4��d`���%�ƃp����>}x?턍>B�I?�<?�wP?tkL?{��>i`�>5��o�>���; �>��>��9?�-?@60?�x?s+?P*c>���������ؾ�
?��?JJ?�?�?�݅��yý?��� g���y�g|����=�$�<k�׽�Pu���T=T>V�?�T�م3��f���/>Ga0?O?�`�>MJ��}1����t<B]�>(Q?@��>��߾߿s�`S�3t�>; �?]��&3W=AF\>��=����5_�4Җ��.ܽ�� >��B����Dߓ=D��=>��=�"=9bi��2k��f�����5�?Ӏ?���>)=�>���A%徖���:�>�_>���>�{>��ʾ!��Dy��)H\���>Ԙ?0�?g���\��>��F>iQ��B.�D�����jӤ>��O?���>�C?$R�?�2?	C?���=��%�����YX������w�>�,?�q�>%����ʾਿ^e3���?�J?�:a�+���2)�ڬ¾�\Խ,�>�(/��#~�����UD��[�����g����?F��?�@���6�=���Ș��ޫ��kC?���>-}�>�>��)���g�/�}�;>�|�>H�Q?�"�>��O?�;{?0�[?0iT>��8�G1��qә��3���!>�@?籁?^�?Py?s�>��>;�)�!�U����������:	W=�
Z>1��>K(�>��>t��=dȽ�Y��@�>��^�=v�b> ��>*��>x�>u�w>@W�<��G?<&�>i�{�Jk�lh���à���J=�Im?��?w�'?�����1���U��_�-�>Y�?G��?��.?n�'�]]�=��!�����!���t>t~>�g>�J�=���=
>��>�ޞ>)����$vF��A<���>c�F?���}Aп
����W�����<�����ξ@�D������"�F4>����\,�
۪�Լ]�詛�-���W��w ���Np�y��>؏=>W�='>DYk=/�O�auu<e�e=Ʈ=�&=�������l�	7*�%�=]�3��X�<߶�<>3����ڼ������?���>..F?�?�?�7n=��=���c?܃Y=�D?dt�>#J��>5��ξ|����e����D���fS
��Τ����=VN�<-5=Ϸ�<�Y�=!፽�k#>jCJ>�N�;v��㟐�O�I=�T=�F=�C>���>B�/>�)s?0T��@1����l�^S��`?�1�>��<6��Bd?���=����N��`��Ά?:F�?A��?��>�zý�Ŀ>�־�RҾ��=�]>��?*�=U-Ǿ�J�>R�>��=�������ֽO��?k��?;,W?�씿�᫿�H< �7>E�>��R�Ty1���[� /b���Y�I�!?n];���˾�[�>��=��޾�+ƾas1=:�5>$d^=� �TW\��=y�y�0w>=|\r=߱�>�C>|ۺ=w±��:�=��I=/��=�>P>5���\6��-��1=��=C�b>N�&>��>���>pH?�+U?D�">���������e��Y��>��=޿B>L�I�o��=��>ڼP?��S?�[u?J�>"�
>���>XI>���&=��7!�	� ����=�?�?�(r?3��>���=ι�<��K���=�l1?�56?^��>SPh>w��~s޿�
�[�"�?s��щ�75ϼ���/򠼍�[=}Zk�[�j�ܶ���>�Ů>��>�9> ��>兪>���>�WQ�{zE>y��=�-6=��T�)V�=�dk���8��X
=�~�<%��h�C@�=�<o�4=A�>5=/��=��>6q>���>?�=����1}.>�ޖ�5sL�oT�=���� hA���d���}���.�t1�oE>/Z>ӆ� ���?�1[>�B>E�?ּt? �>�G��վ~ӝ��c�:�O��8�=�P>??��';�տ_�EWM��.Ѿ8��>ގ>��>�l>X,�I!?��x=�⾴b5���>�}�����J%��7q�n>��n����i�_�Һ�D?�E��{��=d"~?��I?r�?��>`#��Y�ؾ�A0>�H����=D��&q�ya����?u'?��>$�3�D���0���o:?OGC���:즿����n���%�Lo=���� ݾ�=C�6_��M���{���Y�[{ ?=NR?��?���R�#�/Q�r2ξ����&�?��N?U��=;	&?ƥ�>�2�L����6Q�؍U>U?-��?��?+�4>*1�=>o���c�>	?8��?i��?�vs?^s?��[�>߅�;�1 >����Xv�=��>��=���=�?�
?2�
?K�����	����s�񾪏^�aK�<���=<��>�k�>e�r>�'�=��f=�L�=��[>��>*C�>��e>T�>o#�>xF^�������'?��=Z�%>8? ��>������s���ShA�+Ad����(�=`��^���5�=t[�=T>O	?&��% �?�ќ>�?��R�?o��8Y��-�>��9>��7�wb�>2��=��h>��>I�>��
?�л>�J=YIӾ�}>����c!��+C��R���Ѿ�pz>3����&�����z���II�:s���h�[
j�;-���9=�n�<�H�?0�����k�M�)�/�����?�\�>�6?Mތ�S����>���>�ō>+N�������Ǎ��b���?���?SM_>�А>�;e?jW'?�~n��
H�/�J���j��R7�9�T��]��̅����qo���B�f?I4}?z�D?��<Ih>J}?d$��m���>��#��-����=�v�> ��pD-��
ݾ6̧��ML�<1<>��a?��?l�?=�(��0���*9>�2?}�/?�"s?~5*?�+?�=���-?iY>l�?��	?��.?��)?g/ ?�>q�=����(F*=�X��䄉�`0ͽ�3ӽX����=i�\=�%?�X��<�]=0�<��ۼ`i[�~�ڻ�ټ&��<l�c=S��=�=���>%]?r�>���>��6?�-�8�.�����.?dN<=I͂�p����Y~�{f>3:k?r�?�@Z?@c>B�1$@�H�>'��>I�&>��[>�6�>�꽣�B�k�=*�>��>�+�=c�W��ρ�|�	��鐾�R�<�( >�_�>�r>;䃽#=->�*��&n��et>dS�	���yU�8�H�~,1�KAq�(�>7�J?�?�=���[Y�p�e��3+?6n9?�I?Z6}?�=��о0�4��J�� �ם>�R0<=�d���􁠿3�8�
��P�j>�ܚ�Aߠ��Ub>r���s޾��n��J�	��(HM=|�UTV=����վ�3�H��==#
>������ � ���ժ��0J?G�j=9v���`U�2p����>���>�ޮ>��:���v�؇@�P���-7�=H��>��:>�]��O�~G��7�=�>HPE?�V_?|j�?�#���s�x�B�����	c���)ȼ��?\w�>�h?�B>��=G�����&�d��G���>
��>{��p�G�Q8���1��)�$���>[8?e�>��?��R?��
?��`?�*?9E?$)�>x
������ B&?0��?��=��Խ$�T�� 9�?F����>|�)?�B�Թ�>B�?޽?��&?�Q?�?��>� ��C@����>�Y�>��W��b��>�_>��J?皳>t=Y?�ԃ?��=>S�5�ꢾ�֩��U�=�>��2?�5#?C�?䯸>4��>����L��=>��>��b?�#�?��o?�w�=F�?�X2>F��>$��=Gf�>7T�>Y?c^O?^�s?��J?Tq�>�+�<�﬽�'���ms���L���~;��F<d$z=8����s�Wh�4��<��;za��>����w�	E����X��;��>��J>����6�>�tѾ�,p�)W=>!e	�����M����$O���}=�"x>�V?1͢>e��6��=/�>S��>̳�� (?}A�>�?��3[��沾����Ѻ>��G?���=��r�ג�x�w��K=J�p?��T?�[�����b?=�S?�"�#)G�e�V�4����!5~?��?��x��,?-Rn?D_`?�o�>�~_��!l����sO���,B=�>9� ������i>�-?f��=f�	<X!>dz���@��w��3�>U?��?J�?�� >��r�����Ud>�����Y?���><ޕ�;�>4���Ϋ��ᴾ�'����tUɾ�;���W̾oAK�t�;Ґ��u>�0.?W�j?�?y�W?�d���Y�z��3����f�!
��<B��V-��UN���T�@�~�Ð�=��X8X�x��=-c~�CSA��A�?�&?Y3����>q�!�̾ڞ?>���Q��a��=����J�E=:�U=��e�h/�H«��?R��>���>��;?-[�q>��U1�}77����f�2>{)�>�>F��>�#;��*�$�ҋǾ�ǃ�>�ӽ�7v>�xc?H�K?��n?!p�+1�����G�!�:�/��c����B>�j>5��>�W����N:&�qY>�M�r�o��w��2�	�ˣ~=}�2?q(�>6��>�O�?�?�{	�tk��lx�(�1�l��<-1�>� i?A�>"�>�н#� ����>��l?s��>��>����bZ!���{���ʽ8&�>�>���>��o>�,��#\��j��Q����9�Su�=%�h?���8�`�[�>�R?�:�G<�|�>��v���!������'�M�>b|?���=Y�;>�ž�$���{��7��2)?�?����Qj*��J|>�<"?���>�_�>��?���>�þ�Č�?�?��^?�J?��@?@��>�=Rx����Ƚlb&�}B0=&:�>ώ[>8�e=��=C_�)�\� �X�D=�r�=ʼ/Y��q�<�X��@[T<��<��3>��ܿ]�I�)Fվ���4D�6�z����Ž5����)��д�t����|�[���g@��W��qa� L���f����?4-�?������좚���:������><���͍��3������ՙ����s����|!���N���e���a�P�'?�����ǿ񰡿�:ܾ5! ?�A ?8�y?��6�"���8�� >�C�<�,����뾭����ο@�����^?���>��/��n��>᥂>�X>�Hq>����螾B1�<��?7�-?��>��r�0�ɿb���{¤<���?0�@~A?_�(�}���#V=;��>�	?8Y@>�0��O������>�A�?D��?XN=��W�\���Te?i}<��F�`E�pl�=9פ=��=b��IJ>�!�>�-�^oA�'ݽG}4>�܅>�#�A�+D^�?#�<y-]>�ս�,��SԄ?��\�pf���/��N��1�>��T?E�>v�=�,?I2H�=�Ͽn�\� 0a?p/�?��?��(?�ӿ��֚>y�ܾw�M?�46?���>GY&�Ѹt����=�߼\�����V����=A��>��>��,����m�O�T���=�;�S;ƿ�$$�'��`=@����l���/���Hd\� ӟ�!�n��i��f=��=ԹO>���>�>W>n�Z>��W?��k?���>�9>���
ʉ���˾��[�/���f�5}��El�������zᾥ�	��������Ⱦ� =��=7R�o���)� �:�b�C�F���.?#w$>\�ʾ}�M���-<Wpʾ?���ۄ�H᥽.̾�1�"n�U͟?��A?������V�L��RX�����5�W?OP�Ļ�yꬾ���=���T�=�$�>n��=T��� 3��~S�_[0?�p?r;���k���+>�� ���=x�+?�� ?�V<;��>�^%?d,*�#�㽊�Z>n�3>|@�>7��>^8><W����ڽ@?Y�T?}��ś��XƐ>$���{�ݚ_=��>�34�����[>"�<Q���TO�I׎�Tc�<�j]?���>M+�ht���	 ���=���>�N�?Й�>�q�>��}?��Y?5ǹ>2��&F���������Ug?��b?<6>ߌ鼅��dnd�%L�?傇?'׃>��Z�03Ӿۅo���i�_nI?;`?��O?�"��B[������95 �Jf?��v?s^�ts�����a�V�W=�>�[�>���>��9��k�>�>?�#��G������tY4�(Þ?��@���?J�;< �n��=�;?}\�>�O��>ƾ!{������x�q=�"�>���nev���� R,�\�8?֠�?���>����������=�ٕ��Z�?}�?����IFg<>���l��n����<ZΫ=���E"������7���ƾ��
����5࿼���>@Z@�U�p*�>�C8�[6�TϿ"���[о�Sq���?Q��>�Ƚ����9�j��Pu�Z�G�.�H�����Zit>5�9��_T>�$þ��u��K#�x˽��s>�+��]�>!�پ��Ҿ�ƾ@���>U��>�]?,��=^Ȝ���?F9��	�󗟿���Z\o?V��?�Տ?��5?��>)��4~��s�=�E?��?�a?a�? �� ����j?%N���T`�6�4�4E��NU>�+3?�i�>��-��|=TD>���>��>�/��ĿT۶�����`�?	��?Xk����>v�?�a+?1_�L9��������*�y��M1A?r2>�����!�1)=�������
?�]0?���-��h?�t���q��.��g��!�?��P��L��J�=���=-)R�Gf���h9�O�?;_@�S�?����x!���?jJ�>�|e��F��-Up>,��>�¬>�Z>9p��ʶ>���.����v<X��?���?���>c����W��4Ó>�Z?܅P>-c�?0���@6-?8�>�i�S X��7�>ծ��f߼�
.?;�`?���>pM��ETS�	�ʂG���c��P���C��d�>��D?FFd?�d㼷�&�/c��@�+ =�i��>C��u��g
���c��|<=�zr=���=P�ǽ r���?Gp�8�ؿ�i��p'��54?0��>�?����t����;_?Vz�>�6��+���%���B�]��?�G�?;�?��׾�R̼�><�>�I�>��Խ����Q�����7>0�B?r��D��t�o���>���?�@�ծ?mi��?��[!��g�}��I��)8�U�=6?���hz>�v�>A�=��v�l���4�s��(�>�{�?}��?�#�>��l? �o�r4B�Z�.=ţ>�Lk?*k
?���8�rE>V�?���%c����~uf?3�
@�~@�]?d�����׿d���o��J뙾'o�=�=�>>��~�>A�=J	A�uټ��=o�>ٟ7>~�`>�W=>�B#>	>�M��G�%�����d��1mL�� �����j��
<
��\�����
���fþ¨��H�ˮ����m��A@�͉�Te�=תU?.�Q?<p?�� ?i�x��~>���/�=�#�X�=�B�>�_2?��L?u�*?�j�=Ϻ���d��W��K��r���'��>�NI>���>g,�>���>������I>��>>|�>>Y�&=oA�;#=��N>qY�>��>k�>�C<>ԑ>Fϴ��1��I�h��
w��̽1�?k���K�J��1���9�������h�=@b.?�{>���?пf����2H?���p)��+���>y�0?�cW?ٜ>1��"�T�,:>5����j�6`>�+ �6l���)�l%Q>Nl?��<>=�C>v�!���$���^��U����>��5?�y��c�D�Wn���=� ��ݶp>X��>�k�����h��2O�����=;?��>������j��&�����>G�>��?=Y�>�r>V\Ǽ�렽��*��"�=G=�9>.�>�>x>xH�>�ܵ�9�P�R�>N�4>&0>�<?�4?7y����!����i�>mw�>ci~>e�=��e����=���>vW>L^<@J��/������68>s	��kt�+�5��%�=ߢ��O�=�X@=�j�wF?�F7L=N��?����������d� �oX?@7�>hc�<�#�>2t������_�,�?e�@q��?���]D���!?�-}?�sԽd->���>��=9��9�ʾ��>�%>8o�� 'T��L���?U�?xԍ=p����r��s>E0+?E%��`Y�>�-�wȘ������xu��=̆�>��H?7����)���8�N�	?�?�������nȿ��u����>�%�?8ܔ?4=m�/����?�T��>��?�Z?�>m>�۾^�k��>0B?yT?O��>&�#/�P~?ܭ�?��?%I>���?�s?�k�>&0x��Z/��6�������o=��[;�d�>�W>f���wgF��ד��h��n�j������a>��$=;�>E�\4���9�=���H��L�f�C��>�,q> �I>W�>f� ?�a�>c��>�x=�n��,ှ������F?i�?��5�k|�S�>��>����z?��?R�мp�"ĺ>�C?0W?_	3?�}�>�.)�.M����ʿR¾fC�=Y$>�?�G�>]��wj>�Ծ�bھmn>S(q>-H)=�P��\)H�e�i��e�>��:?qd�>�q��q ?&"?(�k>L��>@�E�ӌ��� ?� �>�N�>��?}?�5?���� 5�~������ɊX���g>��t?�4?
9�>cP��%r���=�;���E�H��3�?n�b?�>޽�w?rn�?U�G?�B?�I>�5%���ھU���L�>��!?�9���A���&����h?�?�n�>�k���Fֽ$�ȼ��������?��[?}�%?����Ia���¾^�<�w��zD�+$�;9�A��I>�K>�Ŋ��ٲ=�s>���=�m�O6��d<�L�=|0�>�@�=)8��Ԕ���&?[�/�iνJFW>��|��QO��"�>O8>a0�cVq?q��`����J~�������?bu�?���?��a�y�e�QD?D��?̽)?ǝ�>`���?;�����A�}6ľ�/��SR>b��>.Ի%�վ�Y���m���b�(�ԽK��/��>ܾ�>3l?���>��N>j˳>'����%��^��f�^�/��58�J�-�H2������"��*�-�¾\�w��t�>�2��5��>?I	?�e>Gt{>e��>��f��>tWR>��>z��>Y�T>�3>�y >�<Uν��??�ܾf����˾���=u?��??�i�>6Zk�:1x����b�?^�?~3�??oF>�ځ�VR�Q��>?16?��¾:zB?=�=�a�=�Ž+�H��i̽�x='�j��7�>��v���*���Q�N��H��>
&�>��E��D����<��Ѿ�YF=�5�?�&?M(���W��Cf�gPe�LY�v�ͽ{���t���X.���o��'���Y��cu��2��=Q�5?9D�?|�Ծ��[rƾ�6a� {#�v�>9��>��>�ʓ>�X>���ˌ5�l�Y��!�����f��>�fr?���>{�I?@<?yP?_gL?f��>�e�>n3��k�>X��;p��>7 �>�9?��-?�60?F|?�u+?�5c>@���A��$�ؾ[
?	�?�K?1?��?܅��vý�|���g�q�y�}s�����=T�<��׽[Ku�n�T=�T>[�?����_7�wH��p>/q>?+?���>�ӑ�-��QGl=K��>�G?pٕ>h~�i={����H�>�e�?.+8�\�h=�$>���=Z��<��L�AC�<}�;vH�=ڿw�L��F�#<ɢ�=�g�=���<�˼S��_����x=���>�X?^�>E�>h���{��U���4�=߭'>V^�>f�&;�vȾF�����=Z�᪬>"�}?��?:����1q>sP�=��	���f˾����	> �?,��>'X?%Ĵ?m�(?x�a? J>:E��֌�~��dŽI�?�,?�q�>����ʾ�򨿈`3��?_?�#a����D;)��¾YԽ��>�J/�p,~�����%D��-t����d4��1��?���?Aq@��6��辫���X_��rtC?��>�f�>��>p�)���g�E��:;>W�>J�Q?�#�>��O?={?0�[?�`T>�8��0��cә��o3���!>�@?��??�?�y?�v�>Y�>�)�*ྵO��n��;�$����W=�Z>ʎ�>n)�>w�>���=�ǽX����>��R�=Q�b>���>���>��>�w>?�<�F?	�c>�	[��y�5辨پ��H�>�i?ӵ?/�i?i^j��F^�_�S�1�G��>k<�?p��?+��>t6ݽ!��=��=���o<�X�>�zh>��9>��!=P
>��>Yz�>�>l����:���=�A]�<:��>F�J?�,U�OLǿ��i�d5.�����u�)���LiT�o���L|��9=Q���N���ؽ�Y[w�4C��J"���?��$�zO�
?qh9=��>Ct�=d#����P=m`<���<��1=T��ߣ=�:�� ���I{�=��+��<X�=c�˻a�>�G��?!�>�a?�%j?h��Z���!Z���<>�����?���>v����	þ����|�����pZ�e��Hf��E4dF>8�*����==e�=�9�=�����Xc>�5=RR�����@%=��,>ɒ�=��.=�>qh�=z#>"�t?势�����Ns�=-I�V�N?>K/-=`]��MAH?�=�=g&��z���� ��?��? '�?��>Ɔ;�KQ�>���Lס���=@B�=�
�>�h4=@�j��o�>�Lq>
���PV���:���?FR@;�8?O���ɿ��+>t;>��>ݺT�t�0���G�B�`�q,^� �"?U�<�S�ʾ��>�q�=[�ھ?�þ��%=�7>ٸE=b����`�=�=>q�Cy)=]��=���>I94>��= Ȯ��w�=N6==��=�-T>����C�=���3�m�"=B��=�h>rQ%>m��>�J�>1{:?z�-?�7>@�q��맾��=
p>�N�<�@W>�s4���>���>�+D?F?!�Y?o�>kP2>�X�>���>4�)���U�O��Ѿ:JN>C̍?լ�??�U�=�&ɾW/%�e^A�8r���:?�?���>n�~>�U����9Y&���.�%����x4��+=�mr��QU�S���Im�2�㽱�=�p�>���>��>:Ty>�9>��N>��>��>�6�<zp�=.ጻ���<� �����=%�����<�vż����u&�9�+�,�����;���;J�]<Z��;$��=���>	6>}=�>u�#=e�� �>>�j^F���=����:i?��i���|�N�(��P�ޫV>�'c>���C��`^?�e>|�?>oz�?3#r?�I>�	�@5׾�ś�J愾�^O��(�=�j�=��>���8�b�[��L�c_Ǿ��>�׎>A�>i�l>�,�(?�#nx=�\5�F�>Á�������0q��;�������i����=�D?�D�����=l ~?�I?Kߏ?�s�>@��A�ؾ�.0>M��A�=��q�R]����?�'?��>�쾺�D����r ���1?��G���=�?���j���~ݾT`���w:>����f����[��]���݊�I�0�T*����?#�7?p�?U�þ}K%�?�B���Ⱦ���=�>o>�rS?o�8>ǉ ?ì�>��a���\%��$t�>�)i?��?Gv�?������=�S���J�>�	?:��?���?trs?x�?��f�>��;� >���U�=��>�Ӝ=)�=�y?ڋ
?��
?����	������&2^��=�<��=b��>�e�>��r>G��=*�f=�=�2\>t�>��>`e>#	�>AE�>�P���-?�8����=?J"?xXE>���8Ƚ�-���A�I���c�Z��=�n�;k�u�$��=�bC��K>�T�>�ܼ����?<�="���>����g�"��=�C�=+��&�>���<�Z�>`��>Y��>�'�>��>|�>lMӾ�z>����]!�.,C�ՃR�O�Ѿ�cz>$���/�%����ex��YJI��v��vm��j�+��A/=���<�H�?c���$�k���)�v���#�?wm�>�6?�ٌ�G���>���>�э>G��ݐ���ƍ��j�.�?��?��b>���>�mX?3o?d6��2��`Y�$�t�*6@�F9d�Ya����� ���j	�q��oD_?�Ay?��@?X��<�z{>��~?*�$��q��1�>z�.��9�z�J=�,�>#���_�g�Ծ��þ�a��+G>�o?}��?Q:?��U�Q�m��'> �:?��1?Jt?��1?P�;?L����$?�g3>�C?�o?�N5?^�.?��
?��1>|��=�7��(=�;��{��ѽ��ʽ���ҡ3=F*{=�J�f�
<�p=���<�u�N�ټ��;���3�<I%:=r�=��=�>��U?֍ ?~F�>��'?��,���*�P}��J4,?*�=)噾C����׷�2����=^�m?_��?�nW?C>�E�|<'�c>!��>��>>'�D>9��>)�ǽ��@� �=k�>1�>�o�=���	���ҿ�ђ��VG=�Q>I��>Wv>�Շ�?m)>A+����s��a>U_T��F����T���G��0���v��J�>�K?۲?/w�=�&羓Г�&f�)*?"�;?��L?�n~?�	�=�ؾmE9�}^J���R��>&��<�{	�ܢ�吡�wk9�b::�p>�/��Sޠ�Tb>���t޾x�n��J�O��]TM=_~�JV=����վ�2����=*%
>����,� ����ժ��0J?Ĭj=vu���ZU�p��+�>f��>�ޮ>O�:���v�U�@�𯬾k.�=f��>��:>�#��f��+~G��9��;�>�SE?�R_?mm�?N���
s���B�}����j���ȼ$�?P��>�h?�B>�߭=d�����V�d��G���>ע�>����G��:���/���$����>�:?D�>��?�R?M�
?N�`?*?�A?�#�>�!������B&?㈃?��=�Խl�T�� 9��F�d �>߃)?�B��>��?}�?
�&??�Q?L�?��>� �C@�֔�>-Y�>	�W��b����_>.�J?ݚ�>�=Y?	Ճ?	�=>"�5��ꢾF٩�P�=D>��2?�5#?Q�?��>c��>譡��=���>�
c?i0�?��o?[��=o�?;2>���>H��=���>���>�?+XO?I�s?��J?��>��<f4��X7��@s���O���;|H<��y=m��h8t�SF�Q��<"�;*p��4Y������D�����t��;%H�>xl>�4��2�>��ϾнO���V>~��ϓ����5V��y=�Sz>�2?;y�>�;���=���>#�>0��[#?�+?�8?��u<?`_�.�ھG�籧>�>A?6�==�h��M��G,s��q=<j?��\?r4U����`?�]Q?��,�G�O�ӕ�<���a׾�C�?J0?u�þ4f-?�D?�d?�>�����k������{@�|7
�j�s=$�x>�F羛a�|{>��?}sm=��M=��=�k[�׈J�����c>�UU?��?���?��>9��a��X������Z??q�>�-���&�>�bh�>��~{���\���k�����{?��M)��C���'&�S{��ν���=�+?�(�?=܈?��I?�޾x�T�3�(���u���I��r��9���>�OqN�giR�0R���<$�o}�0��O)*>�C�	u7�u��?7&?.IO�Ȋ�>"���p��=<���e6>RѰ��9���=s;=} >��i=cn����7��(Y�ɑ*?�d>�>�o\?��=�/bb�ח2����u/꾢u�=2-�>�h�>�շ>fO&=�X4�j.�=�̻�z���B�	�I4v> zc?K?M�n?Wh��*1�������!���/��d��Q�B>Ct>d��>�W�6���9&�Y>��r�����w����	�٨~=+�2?Z)�>��>�N�?�?�y	�7k��6kx���1�$��<S0�>i?�>�>��>�н� ����>��l?\��>��>ŕ��GZ!���{��ʽ]%�>^߭>ķ�>�o>-�,�e#\��j��>���(9�	u�=˩h?�����`�]�>&R?�͈:��G<�{�>ǫv�s�!�#��n�'�Z�>�{?<��=W�;>vž�$���{�8����(?��?�����+�k�o>%%?Ƚ�>�>	R�?���>�`ƾ7���&?2`?*�I?�=?���>`-,=�(���vʽJU%� {O=ed�>�mV>.bS=���=���5�U����U=�X�=ǌּ�S��O^�;良׭�<?��<�F4>�Wۿ`*K�0�ؾ���~��l
�9�������oQ��p�	�2_���𙾄�w������&��IU���b��ߌ���l��S�?<�?vݑ�5��#.���<�����4��>Q�q����먭�8��ۖ��{ᾭ_��x�!�j�O�U�g�ܸd��'?͹����ǿ����;ܾS" ?�B ?L�y?���"�8�3� >J�<���ܜ뾮���x�ο����E�^?
��>N
�0�����>��>ӡX>8Iq>���T垾�3�<��?��-?i��>��r�ߕɿ���1��<d��?�@A?=� ��%��G]=Mt�>_?��<>�	���"������>���?A �?��N=$�U�M��hR_?�qZ;w�M�&X���r�=�D�=��=e��~GA>���>Q4��c\���ͽvZ'>m�>Q�����>�h�u>�<�f>�]���]��yԄ?�\�	f�Ϡ/�nO����>��T?(�>�=H�,?3H��Ͽ_�\�&a?p.�?��?��(?뻿�rњ>K�ܾv�M?�A6?��>q&��t�X��="�߼�v��k�㾎*V��Z�=���>��>�,�͟�C�O�����~Y�=�.�UDĿ�A!�������<��ؼT���0��ǲ�秂����If��r߽И�=x;�=v%R>hـ>ι:>�H>~�W?�'o?2Y�>*z#>XT����}�)���Rc�����$���W���Y?�Ň���i�Q����y���I���� =�s�=w7R�\����� ���b���F�#�.?Tw$>��ʾ%�M��-<oʾ����ބ��᥽;0̾��1��!n��̟?=�A?.�����V�#��;M�߅����W?�S�ݺ�dꬾ���=����=%�>���=M��!3��S��Z0?�%?{����]/> ����D=j}-?e�>�]6<)F�>�%?�U%��uὮyW>L�5>�r�>��>���=�+��_Vҽ��?	�V?j��\5��=�>tg��ә���h=�Y>�
,�ϸ��Z>�lR<2���F�[�}�Z�<6[?�ٜ>z�,��5����:�>iT�>9�?U�k>���>a�y?��C?*��>��޾�����0������}?���?��$>Cnʼ}���׊�ďx?o�Y?]ڷ=�b��vrȾ�dL��G����>�9�?!7\?֣��5�����ߢ�9�r?��v?�r^�cs�������V�Q=�>�[�>���>��9��k�>��>?#��G������[Y4�+Þ?��@z��?L�;<| ����=�;?�\�>�O��>ƾ�z������W�q=�"�>���Kev����'R,�E�8?���?}��>ɓ��������=�ٕ��Z�?~�?����KAg<C���l�gn����<=Ϋ=���F"�����7�{�ƾ��
�骜��࿼���>@Z@�U�x*�>�C8�S6�
TϿ$���[о�Sq���?G��>�Ƚ����E�j��Pu�_�G��H�Х��;��>r�<�F>`Ѿ����3$���&>L��>	Lv����>^x���oɾW���#	��@�>�l�>�L�>z�>�Ke�i�?p ���߿� ��!*%�&�?��?ڬr?�;?��{>u½�=����S)?_��?km?*C�T����e��ĥj?����a���1�%u>��MT>��3?Dx�>�w,��>=�;+>[\�>��%>C,�Ŀ��p���8�?�;�?���j��>w]�?J(?�[r��ɰ��S'���8<.�;?�9>��¾��"���;�2���
?
c*?�e�؀�O�b?�\{�v���-�A���	�
?D�2�Y6׾���=�=3>�EP�t������ĥ�?�*@Ȱ�?�� �(����?�d�>�.W����{�;���<�9�>�f�=�=���>��*��R[�9��;�?7� @���>� ��Z���S��>��{?볛>ZĐ?Y���4W?�>��]���(�>���%�-��+?}̀?�?��������ھs&6���Q�s6Q���=���>�N@?�]?��=[!��)G��Q<��R�=Q�8�S �����<�4��T��
>�rA:���=Wפ��T���?Y�0�ؿ�_��?�&�x$4?Nǃ>M?���Zu�@�
�'_?�>�(��*���,��7��ԗ�?D�?��?�׾S̼{�>W�>X�>ˇս�㟽EV����7>4�B?���G����o��5�>��?�@���?Ui���?���oЅ�#������0��>�p5?��ﾧ̓>`��>�=�x��l��:�o�~�>M��?[D�?}��>��n?	�p�L,G��[:=F�>�+p?ec?R�����$jO>*
?��%���i ���h?�T
@�r@�`Y?����0ɿ%���f����y�!�=�/I���>�*���C>�@>)�Z�K��=$�=_D>
�>�T>�

>�;s=D�>\�|���*�E���⟅�֡G�	x��
#��=���_�� >��q�����㧾�g0�7�ɽ�2Y��t#�fӓ�H����=�V?D�Q?J�p?�� ?q�z��>���ͬ�<�$�-;�=�W�>42?�L?!*?(�=�����)e�Eq��Jj��1^���b�>�H><��>���>���>�5Q���J>5w>>*�>���=�&=u?ĺ�w
=�7N>^�>���>@�>�N<>��>ϴ�{1���h�5w�R5̽� �?���b�J�8+���:������"d�=�^.?�y>���?п�����.H?;���J%�:�+��> �0?$bW?J�>��ѣT�8:>�����j��Z>�' ��fl���)��Q>�_?��f>Tu>h�3��q8���P��v���_}>��5?x����l9���u���H�xBݾ��M>�׾>A�R�tH� Ӗ�\�~���i��|=bi:?�\?�ʳ��Ѱ�K_u�ܝ�]SS>ܑ\>�]=��=*M>��e��ǽ=�G�¥/=9(�=�#_>�~?�a >�V>���>]Ѱ���m�J�>X�'>'dV>0ZA?R�?Q����/�������V>�>`��>���>]P>w\�+�>gd�>7N{>��ݻ"%���A�	�Z���B>(��dQ��8����=Yܽ20I==(s=T��r4�bU�<z.?�˟��vw��H$���]��l?l�?n\=�\(>/�	�&I�����G��?�@hL�?����z�.�j�?Y�?����8җ>߿�>�"/>���aq�|�(?��T>u�#�}�]�ր$�c��??U�>�%��JDt�C>���>}������>�"
�u:��0���6t���6=���>��I?�����8���,� �
?u?�����{���ƿ�r��}�>���?�Z�?�.k�Ü� �@�22�>���?y*\?D�y>�B��pU���>\�B?"oX?���>|W!��B��?��?1�?h�H>���?��s?~��>> w�7X/��5�����R=��R;Lp�>͓>����aF�iԓ��c��M�j�P����a>,>$=��>��=?����=��GJ����f�ĸ�>�:q>��I>�6�>�� ?�W�>Ԡ�>��=�f��$Ѐ�������J?�r�?��,��b��Jd>��=�W����$?��>Z=��3�E��(�>I�C?��S?�.?AO�>Tx&�� ���ɿ�&���>nEN>sB-?Rɦ>�a�<8��>Mߗ�qA��5�>+ی>��?>lÐ���T��j���`�>��G??T?���)� ?��"?�n>�&�>��E�$�K�>����>lI�>��?�X}?��?�����c6����m���LbW�ۺc>�u?��?կ�>�ڐ�����q�9D�����9�KT�?��_?h=ǽ
�?��?1�E?q�C?�H>�q%���߾Z!����>E�!?,E�	�B���'��?��??w�>�k���߽�Mr�$�������?BZ?c$?��K9b�G�ľF�<N���X(�Z�_<�.~��E">�v>q���队=��>d�=�(i�|-7���1<�`�=�b�>2��=�9�!���s�,?"me��
� ��=��~�W!@���s>U*->ڵ����o?�X����l��,��k��IB̽���?v��?6g�?�U� �^��K>?�6�?ZY?�>�>]z̾6���6���~����>���>���I���t���#��{^�}�:���"s�>X�>&�
?8
�>w{W>p��>r���m�&��]�z�q^_�X���6��x-�
�C��w� ������¾��x����>W����>Y>
?�Cj>�~>�[�>�҄�LX�>�]R>0O~>Kv�>3?S>r�2>
>�
I<�;ǽ�I?�o��~$����o���Ba?�h?"#�>����XJ��������>\��?�x�?]�>���+3��N	?vv.?&���,?iu�;��;2hP=������n����|�*I>��Z���@�\X^�:;ԾD��>��> u𽝞�����ⴾ5�>=NI�?�p?�� ��~W��^�D�]�y�M���'푾�ġ���'�0�k�9������Ii|�4U��ߕ=��7?��?:������]���d�U�"���I>Nd�>��>�M�>�8U>�4��T8�5,d��5�YiV���	?j?���>T�I?<?xP?�kL?m��>�c�>�3���l�>��;@�>^�>�9?Z�-?�70?�z?�t+?4c>�������ؾ�
?l�?�J?�?�?Jޅ��sý8g��� g�ϳy��}����=~#�<��׽�Du���T="T>�	?	νn�1�c	��0�=�;V?�(?8��>���.�ӿ0��ԓ>� ?�>u'޾�w�F��Z�>lЉ?�aE�&�;��u>��=�3�8��򈃻dmO=�[O>�=���<aZ�=���=�"=��Ѽ�j=�׆=�Y]��9B=]p�>�?P��>8��>v,��)G����j��<ku{>KJf>�=�ھ"7v��B����]�i�>�d�?Uk�?�q�<)?_>]� >K2��t;=uƾ���:�>��'?�5�>kNG?�)�?f�P?]?H'>��:������B��
�ǽ|�?�,?F��>:����ʾ���3���?]??;a�Ǻ�6)�5�¾��Խ��>�X/�9,~����aD�����������;��?9��?�A���6��y�弘�|Y����C?<�>{^�>0�>`�)���g�Q!�J<;>���>oR?"�>��O?r;{?:�[?�kT>�8�]1��Uә��o3���!>$@?<��?��?�y?ar�>g�>��)�}��V�������߂�W=hZ>퐒>�&�>S�>���=Ƚ�[����>�?^�=
�b>{��>ʟ�>��>��w>pH�<��O?��G>�&v��!�)a��&�����:�n?���?��3?���>R���g�5K����?i��?��?�*�>���>�c=2��H�{�ק�>�p�>I->�/O�Řμb��>��>�_�>e<���qP��,:�/�T�5n=?c?c
��ѿtqx�����z��3彮��W����*q��Ε<m��$��=��h�	]A�UCk�\C@�(�~�_kľx:��]��>�/>�>�UB=8��;x6D�߈<=�ǩ=˱�<D͓��9y�vÒ���A��B`=2��!g��
$�<8�6=�S�<���5�?��?�`�?���?�S��-y��m��K(>�ɧ�}�?�m�>��Q=(ѡ��ն������"�&���-�X|���Ā��*>v��Z.D>K��=G2>��U=@��>^� >N�	<�R�18=�>�)�=��=�>�"�>^5�>^t?7��"O��˒Y�o�ν-�e?��>cr�|���"��?���=p2z�{ÿ��/B�?�i�?n�?:��>h�E����>�������5>^P�>y��>��&�]����r�>��g><�t�O��\�Oz�?�b�?zH?6����տ ��<2�;>m�>iyS��50�$\R��Z_��qY�~�#?fm=��9̾��>�
�=\�ھ��ľRT"=�
9>3>N=�����^�,0�=S.d�/H>=��=���>�A>���=J��#�=�SQ=5u�=o�W>�:�G6���@�*e6=t��=�/k>�N%>��>�>�?F?�0i?~Q>_����~���DP�PV�>p<^�9>��G��b�=��>�FO?T?�<C?,|%>!S>!o�>�'9>�@��c�^U�>v��Q��=�7�?G��?��>ӿ<��4�� S$�1�K��5���4?�?Y��>R�`>~��;ǿ��K�|d*���V���)ྌ��C���@�L>�N�=GI>�k�>7��>�N.>�v�I�<��>g0;>�x_=��#=� �ObZ<�Ļ��=Ǽ1Á�W��<������a����<m��<ȟ�;'v���<6-�;W��=|��>Z�>D��>{p�=gJ��*o/>𼖾�=L�&��=dħ��3B��Qd��s~�=�.�ճ4�VD>X�X>�V�������?<Z>;@>�U�?I�t?�3 >v��-�վTI��-�d�DdS��F�=B�>tT>�YA;��;`�%�M��FҾ���>�ߎ>��>y�l>�,�"?��w=v��a5�_�>�z�����E#��8q�@��K����i��Kк��D?F����=�!~?v�I?,�?���>�#��O�ؾ�<0>�I����=b��+q��h��`�?�'?ޕ�>�}�D��*ھ�<ݽ�9J?��ɾ[%$��z�����/�;�������A>������tUW��+��i���S�M<Ἂ�?�L?�x�?��{@4���Q�,�	���=���>�~U?�2->b�7?k��>/7��|$�[g���>��n?���?GG�?�g�=���=B3��è�>�?d�?�?k�s?�?��%�>��p;
�>���3��=��>-�=���=�B?N�
? ?�ۃ	��}�%��^�<�<H��=��>���>�s>"n�=��h=+�=�cZ>��>�u�>�d>@�>��>�.��; ��t)?��Z=�<>�D?j5�>s58=k�*:��=�r��
�a�ͭ����<�O�Zi.�?5�=lځ=� �=2��>����!Ɵ?�A�>Z`žT�>����K��=HaM>JL���>��2>@��>�_�>
��>N�c>�S>Pk�=7�ӾV�>Ɋ��� ��B���R�Ѿp�v>�Ϝ�Ƒ(����� ���J���������i��避�c<����<W`�?L���_�i��'*����}�?�w�>Or5?��;����>��>��>�.��s����퍿v��P�?t��?�c>��>�JX?��?��3�G$5��fY��.u��?���c��`�����l���<�
����_?�!y?�TA?c��<�Ty>���?�P%�OA��� �>n/�(:�P�9=�U�>�.���{]���Ҿ�¾pZ�6wB>B�n?]m�?{L?��W��m�?'>��:?@�1?hSt?�1?�;?t���$?�j3>�F?Nq?M5?��.?-�
?D�1>0��=�����'=9?��]���J�ѽǜʽ6#�-�3=��{=�	��<~�=�<�d�sټà ;����Z��<�U:=��=�L�=���>�W?�� ?��>`�*?�10�y�/����R^1?�Xv=9���i��/ˮ�Ԥ�hO�=_�k?Gʫ?8Y?�e>) D����m>擎>�,>�tH>]߳>U\���E��I=��>C�>E��=F���)4����#s��;�$=��	>.�>�2q>IҐ���>͎����?�4�q>|Xa��A��9;c���J���3���o��)�>�MM?�?t�=#���^���f��,?�F4?��D?�z?�&�=9�ƾq8���I�"g���ɐ> ?�`C��g���Ki8��	`:.�x> Ջ�M���Qwb>���O�ݾ�)n���I�����UJ=�q��@Y=�����վ݂�+��=��>- ���� �	�����'
J?�j=�z����U��񺾲">��>��>��=�0�v��7@������=Y��>��:>~ɚ�!ﾅ0G�5&��&y>��B?>�b?
υ?��o���s���D����𸑾�:L���?��>���>��4>l�=����&�4]V�+�@���>p��>���@.A�ܵ���} �
�$��؀>�{?k+>�w?hVF?=��>MAW?:�0?�?� �>�x~��׼��&?�݃?Um�=>����P���7��K��0�>�/?�mU��G�>��?�O?e�?��T?D�?y�$> �N]:����>l��>�Y�|诿�%`>�I?~��>fZ?�2�?��C>o�2����x�0��=S9>�y6?�$?�c?�>y��>�n���g�=U��>>c?�(�?}�o?/��=F�?n�1>7��>�*�=u��>�P�>��?�4O?��s?z�J?&A�>�Ë<�t���޶��Is��SI�'|�;��I<��y=�]��v������<d�;qZ���6�����OB�i���A�;��>&N|>0��&/L>u��v���8>�Y�k ���拾�:����=�l>ve�>�n�>�F5�P�C=�~�>�'�>˂�4�(?�Y�>�n?gp��jUd�!7�J,l����>�@?��=�am������o�-J�=��i? \?��J�k��E�b?��]?vh�=���þN�b�<��N�O?��
?�G�/�>��~?h�q?��>��e�:n���Db�?�j��ж=er�>?X�L�d�Y?�>Y�7?�N�>�b>�&�=Tu۾�w��q��(?h�?��?���?�**>e�n�M4࿑:������"Z?O��>����j?��,�_�Ѿ�f��6�H��S��t��@Ae�Tf��쬾&�|�l����A����=rX?���?o\�?�Rh?pwپa�s��ʁ�@j��W�~iԾ�/��E��J�T04��]W�"�ξ�վ���폲<WW��Z� ���?�5?,g��p�W>]���@
�Ӡо��>v	��83��=Y;S���ڦ�=L =���
r!������J*?Ƿ?4�>I�4?E�C���j��Y�A;/�����<��>0�r>L�T> <漉ƻ<�>�g��F����\��Fx>{b?��L?l�n?O���f.�\���6 ��ټ�ԭ�=1>N��=G�>��E����mL"��p>���n��
�����d	��j=O�1?i9�>E�>��?q?�&�����m�Ǚ/���<갳>��e?4��>��>�5ϽCz$�V
�>��l?\��>��><	���� ���z�>Eν�X�>;̮>r��>�o>;U*���[�x0���r���9���=��g?�����:`��9�>@UQ?.��;GgO<6��>SWt��"�ui�RS#��}	>G�?t��=�P9>�Bž`�
�(�z�"Ԋ���(?';?Kۏ�=�(��|}>��!?x�>d�>�8�?��>e�ľ�E`���?~�^?�mI?t�@?�_�>XG=�*���E˽��'��%=��>��[>��s=݇�=��V�W���v8M=��=�j��݄����;
Jμ�T<7D�<\�+>
ۿ��K���վ)X��_�]��}T��O���釾ך�\��S7����u���
�Mk&�T`�1n�����Eg���?�-�?
�������l���������>��t��x`����2���u�� |�s���q* ���O��Di�B�d�=�$?\ޛ��vƿy����۩��'?��&?�7p?��
��T�]��b��=#��:�r<M]ξ����]l̿G���қP?-w�>���B��c�>o>�^[>�O>��������,�=A��>�.?��?ƫ~���Ŀ�Z����<N��?tE@YU<?��O�i����<?�"+?}e�>T��pH��)���??�ٞ?���?'\1��L�;?�(½f�8�ss'�'��=�_�=O2ݽϮ��p�>i�>� �,i�jY�n#�=��>��A]�ݎ��*�L=3Ɉ><1���-�Մ?�y\��f�x�/�TT���W>7�T?�)�>�2�=}�,?A6H�n|Ͽ�\�x'a?�0�?���?��(?�޿�&ך>t�ܾf�M?D6?���>ee&�r�t� ��=�/�ê��#�㾒&V�B��=Ԭ�>��>��,�ċ�/�O�$*��z��=�����Կ�)�C*��=�<a�N�O=�!��L��¿#�I��D����9k9>�>ռ=��<_s>DiK>�5J>�4E?�j?Z��>T?9>����&��Z�о�]�E%��X�1�^�������ٽ��m��̾���U} �]� ��y����;�Tg�=�R�Uʐ�l�!���b�پE�$0?: $>�
ʾ�rL���;-:˾̝��;0�������˾��.��`n�᝟?.IA?L+��MW�B��U��f=��5ZX?���j�Nì�80�=����=��>�.�=w���2��R��2?]#?�I��DI����=����V=��?Ь�>���>�ċ>*�?��8������e>UJ�>�נ>��>��<��Ⱦ���?#?�S?���[���i�>�žz���CuQ=��N=�(��V܉=���>�b�<����ޛ��*ә�h�=W;?��}>2$��a�N־륨�,�>Pʋ?.b�>�$_>�*X?eK?�=8����B���*��>�=BPc?R�:?�.*>a���j���xe���'?b�?x�>mdؽ�<�|'.�Y���<?*hs?�5?[�!���e��������0?Gu?��3�����'���þW�q>p�>�$?��$��-�>&V-?5��<�.���#���J�/�?h��?]�?�|�����[��=`#?.&�>B,����ܾ�3���9ھ�< >)?�Jƾ��h��6���`��e ?�T�?�:�>�A��f���6>d�����?�Á?�<��r�;=�(�%^�?w*�.dT=)G0��g����=�Ⱦ�t8�h1��g���+꿾�SO=�[�>fe@�L;�Q�>��h��{�Կ���̾�b��o�?��W>8�E�1Ā���A��D�g����,�؃�<�}>0e>�M�=�¾.������j�O?�~��Į%>ړB>i�ξW�����=|Ơ>F?m/d=�A�>�W��?��̾��ܿ�W¿/8��C�[?���?���?���>��3>��\�z
��TK�=��>?��>/��>�C�=�y>����j?�N��X`�U�4�>SE��U>�3?)h�>�-���|=�%>@��>R?>] /�2�ĿUԶ�չ�����?��?�g���> ~�?�n+?�`�73���W����*��`��?A?��1>A~����!��8=��Ԓ��
?9z0?���w*�\�_?'�a�M�p���-�y�ƽ�ۡ>��0��e\�uN�����Xe����@y����?M^�?g�?ڵ�� #�d6%?�>f����8Ǿ��<���>�(�>*N>cH_���u>����:�i	>���?�~�?Nj?���������U>	�}?<�>���?o�=.��>�f�=鎮��v ���>��=T?�`~?y�L?���>���=�i9��e/��AF� �P�ވ���B����>�`?:�K?��a>�#���O1�� �	Fн��.����/M?��DJ�L�ݽnR7>֛9>=�>MA�VkҾT�?7n��ؿ�j��=}'��34?ḃ>� ?h���t�ԏ�%=_?�u�>)6��+��]%��0=�r��?�E�?}�?#�׾�A̼>��>�I�>r�Խz��~����7>��B?�D����o��>	��?S�@�Ӯ?4i�)	?X�pQ��gr~�*��\7����=��7?(�1 {>���>��=sv�1�����s�3��>�>�?�x�?��>�l?�io���B�>2= Y�>��k?lg?I}�����B>��?4��4����X��f?��
@�n@&�^?C袿��ο7L���ܿ����H �=�b�=��@>��ܽQY�=��=[�<t��;�>.��>��1>R�Z>^@.>Zf:>�O>>2���&�h!���c��GO��!�?5	��SW��*
���v�.���/վ�����q�N���	���G�k����d�=��T?�
R?e�p?�l ?�`��@">����V>"=7��M2m=�n�>C�2?�VK?(�(?�=KꞾ�b��o�����!k���>F>?�>�.�>���>"=��%F>�=>T́>)">�o,=yX;l�
=��D>wU�>�l�>W��>>Q=>o�>�Ӵ��s��j�e���r�������?�3���7K�&���ZT��9���z�=�.?�>�d�� �ϿRͭ�ӉG?�����S���.�:�>�}.?zV?s$>a��8�W��>�Y
���q�o;�=V}��9�h��)���N>JX?d�x>�7[>.�9�_�;�4�:�����zx�>��-?Y�������c���7��ھ_$>�5�>]"�%#��1���Mx���x�O�>=�05?�
?�W�M�����c�����&N�>��Z>e�X��'==ɗE>J�����6G������>��>�G?U�>p��=v��>a4���
��C�>�v�=��>[�f?�>46��4G<�. ��g��uV�>7�>�M�=�A�<�����=m^�>�^�> �=�Tݽ������c�o�>��u�>j����� v�=r�>�����>������=y-�=�~?���(䈿��e���lD?S+?] �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��H��=}�>׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l�6>�^%?��Ӿ`�>���s���� ���-u�2=���>�MI?�Q��+2a�*z>�G�?�?	ﾫ��Hyɿ�u���>���?���?�mo�Կ�� >����>4�?]:V?&�e>}8ܾ`�W�'��>Lq@?��S?i��>B��<B)�j?�ô?O�?�'L>h�?�s?�%�>��w��-��Y��L��b�=��%<�-�>� >^���m�E��ɒ�����k����^>Z�=Y��>���Ϻ���=Ì�U쥾�(n���>"^n>+�O>�˜>G��>fk�>��>���<#ᄽ��u������K?X��?p���*n��a�<6��=Ԡ^�� ?�I4?��Y���Ͼ�Ѩ>��\?��?� [?fX�>���|:��C濿?}��Ɩ<�K> .�>M�>w%���KK>s�Ծ;D�Tj�>u֗>�֣��>ھ ��9��f8�>�e!?ʙ�>?��=�� ?��#??�j>@)�>�`E�48����E���>��>5I?�~?-�?,ѹ��X3�0��桿<�[��EN> �x?�T?�ʕ>?������.E��=I��󒽋��?Spg?S��?1�?a�??�A?%f><��O ؾ����M�>G�?�
?�"1f�����r> �?�6$?IP�>�滽4�G��$>;� �n����>��c?�j�>[�.��'i����~��<��k�>π�Z�����+�= ��=�>�<�+���3c>Vˈ>!}4���4��� =a�W=j�K>�9�=Y�	��6>�A$?��>�u���(���~�r�[�+lV>��>u���@q?YHk�o�U�|���x��]e��s`�?�+�?Aڑ?{E�a�y���	?@��?Ne0?�
?HZ���4����	�!.��x�j��t�Pp���{�>���=��S�􍐿V���s���=ϳK���?���>�?0��>�R>���>����ۇ��&����c���SF���־�)��Z#�����G��\`}�#=ӽ?w����Y�Gs>������>�:�>�1~>v�Y>�px>�H˽��>0Bx>��@>�0�>��=5�=�h>���=\F?��bH?��Ǿ��%��+Ѿ+�|��J?��e?�O�>�{B�������	��?��?���?�Hz>��l���2����>P��>!�K����>JJ��u�Pj��Ǿ�.����:�x���s>����k�6��R��M����?"?퇍�SԾN�������i=�t�?�)?I�(�A�Q�5�o���W���R����?%j�������$��No��|��0X���6����(�r*=�*?�ω?����
꾯�����l��A�7b>���>˨�>� �>�@I>a�
��,1�xj\�e%�s�����>�ky?�О>s99?��E?m]?`D?
^�>�Q�>�4ž~��>[�V��o>���>�Q?��+?;J�>
V�>��'?z��=o�ཚ��T^ྷ��>�7
?nj+?07
?���>�,l� \�e"�<j;p�
6��Z�=[MV>TF�=%����'����
�c�8=39?!\_�K{P�5
�SL�>��J?�?6��>��P�ֽĽOC�= J?�?�K7=�� �5�N��:��,>�lo?��W�R[=>�4>�*>��Z�Z��X��=q˒��p>{~=1�����C=x�>s�!��j7��b�=n�=�"1=�>�t�>"�?���>~@�>D��� �^���s�=Y>�S>i>,Fپ�}���#���g�@^y>{w�?{�?ˬf=��=���=d}��OT�����������<�?�H#?<VT?���?��=?�i#?�>�*��M���]��o��ݮ?�,?�c�>�����ʾ�Ϩ�%G3�.�?R?u$a�=#��)�:^¾�Խ�D>�8/��~�{����"D�1��5��<�����?��?wB�$�6�ld�����$��ȁC?���>^'�>/�>ۨ)���g�3���:>z�>�R?�>�>��S?bۃ? GQ?(�=>��2��Ь������G����$�
?!m?���?2/�?���>(c>y2-�&>��N^�Jp���-�=w�U�=7>C>���>$��>�}�>45=>˨�q`���!_�=y�=��>�A�>���>�K�>�-f>謃�wI?��?�;t�`���'W��12Q�O#X?W�?2�?���=��:�D��#�S�>��?VȨ?�&?)W�js�=�dŽ}ؾM��ں>�x�>v�>`f�=7wf��E�>�e�>b�>C�A��m=��^-�xT=���>���>+����ȿ�z�D���s��`�3<���{�Z�*c��4U���=�ڗ��{��ә���:�47���l���E������Po��<�>�A�=��>J�>@�=0����̻�T�<�{�;_��<��v�3�H=%��g�:��{�L?P���=г�=f�D��ɾ~7}?	I?��+?a�C?��z>X>	b:��y�>�����?�X>	H�.-��W�=��������4�׾��׾�fd�fx��{�>��G�`�>�-4>�f�=�x�<�D�=*5l=g;�=����=�
�=�|�= ��=QE�=�2>�]>w6w?隁�ղ���4Q��\�ܵ:?t8�>+}�=L�ƾ�@?��>>�2�������b�Y-?h��?�T�?!�?�ti�Nc�>����Ꮍ�t�=G����=2>��=��2���>9�J>@��K���}��D4�?��@/�??�ዿ��Ͽ�b/>:��>X�)>kf�J�a�B�ž�;����t�[?H3<� D���~�>���>�?��$o���\����7=���=�{ ;z/[�sbt=a��<�t=�>=\�>نT>\��=�$ɽk�>�>�ّ��t�>�o�D`Z�q�ý57#>�d�=DYg=ӳ!>�>��#?UO2?�st?���>������.����>x���5��>����Խ�e�>�![?�Z#?!D?E��>��h>���>3��>B%.���X��rľ>ž��x���Z?��u?֮G>1�)���O�~]��?���"=�*?@,H?�Z�>�"�>0�����%��g�W���!ŽpK=�͌����˹=/�?���s���=A�>鈨>Z� >ɸ>���>��y>�U�>^B�=ܯ�=�O�=�(�=Y^>�E�<�V#=Z�=X=�C�;ˆ>���*�����=�o<>u��=Ni:�����=��>�>Ƞ�>}����Ͼ�[>�rc��D��
>���r�=��xR��<p���p�Խf#�>p�f>G����폿�u�>
|F>$�t>~ڼ?Q�~?%!P>օ�����ZO��܅,����`>F�>y��YV��c�U;A��F��>��>�>m�>�@m>�+�<�>�ؼy=)�l15��K�>�~�����h�'q��+���럿�i�����._D?M2��m��=�}?�I?\�?{k�>o���*^ؾ�$/>:���pU=����_q�������?��&?]��>����D��J̾W����>z7I�3�O�NÕ���0��.��˷���>E�����о�%3��e��������B��Or���>��O?'�?�*b�V��zRO����FI��[m?F{g?��>�F?dB?���|�q��A��=V�n?f��?J=�?�
>X� >&��
��>h2?���?��?�h?}���+�>�cn��r�s�Q��4�>��>}��= ����>Aҝ>��>���� !��?-����H�1|�g��=�}�>I<�>�aA=*=C�B�^>�����=���>��>d(�A��>W>����nh�t}?��=)I}>�|5?uW�>=��=����2;�=v�+m��꙽W}X�y9 �F������t�==����0[�>K�ĿJ��?6CL>�� ��k"?ޖ�	ƽ���=,�|>��6��^�>Ȇ>Yn>�{�>	�>��=�$;>
�@>|�Ҿ�]>����!��+C��cR�tѾ50{>���x�%��l�5�����I��#���a�e�i��$����<��j�<9�?J�����k�X�)�U ����?KZ�>f6?�ی�����"9>��>Rҍ>{'������6č�--����?9��?b�h>%\�>�Ye?a�?��8��oa�	�q���s�K�W�V\^���Y�"����X�#�޾9Q���)V?K;�?��&?��	>/a]>-}�?���8��Q�>�~A���E�A�ȼF
�>+�߾��S�R3��$�ܾ��o�>e�h?`6�?��'?�^A�4	��YG>˩@?<8?��f?nF-?ͺ)?M=��/?�"=�q�>�m?j�7?�>!?���>��=�=���[څ=������u����W�_��4�KJ�<�-�=�}b��~�u�>�$g>͟D��j�r�����Q=�����P)<A�=�DF=�B�>��_??r7�>�
?y�ΩY���Ͼ$a�>n���+�o+�i:`�:�����i>o��?)�?"�?��?�N[�-�l��x>q,>@�>���>zl�>�C��fG���>6Ҩ=?�=EB���5"=���ޤؾ����M�d�9�>�v>�e�~]0>�<��y�u��$]>G�Q�����5_�WtH���1��}t��I�>�?J?�L?1H�=��澾*|��e��d&?>�9?�jL?z.~?Ǭ�=��Ծ�>8��F��.�w��>ٙ�<����2��ѿ��7;��<;;�q>�K���I��.j>����ܾ�Uj��AG���⾐�K=���6�_=9�	���Ѿ�{�e��=�>�K���] �jm��d��K�H?��U=3V��yja��%��W/$>�^�>�"�>�{P��N[���<��Ƥ���=J��>�c1>#0�����mK�B���>�^E?�_?v�?�����#s��ZC����٧�����#)?���>g�?�A>�k�=�� ��Cd��F�B��>�c�>����YH������,��#'%����>lN?�>>�s?0S?n�
?�O_?�a)?��?���>馷��߷�_�"?ۤ�?^P�=+�l�\���1:�@8G��>T�$?{�m���\>2#?*?���>a�P?�$?|>($����&��C�>�>1�Z��~��:�k>��L?V�>�S?�v?�c>(�&�cK���<0�=��=G�,?g.?���><�>AL�>Zz���rW=[�>�ec?$�?��o?J��=�?44>��>2i�=�n�>�y�>s�?��M?H�q?a"I?�m�>�7�<�����}��Ʉm�O���z<���<�4}=F3���k���!��<�|�:���X�u�Y8%��ӼlV�;��>��t>�
��1�.>cGž����~@> ��3��*u���3;�g��=Z�>�?*�>W(!�P��=�>��>$���'?o�?�?0I�;&�a�F�پ��L�2��>��A?���=�l�����u�z�n=�Qn?e�]?2�Y�I���G�b?��]?�h�=���þ��b�8����O?��
?(�G���>��~?-�q?��>��e�l9n���jDb�N�j�'Ҷ=�q�>TX�8�d��>�>Z�7?VO�>:�b>&"�=�t۾��w��o���?@�?��?#��?8)*>`�n��3���6���x�c?�B ?�y���j/?P�f�����E�e�����׾ξqR��f̀��~���l��O�h�j���&w=��?��q?Tx?�c?���q�l�[�k��w�n��L#�i���D�-E�t�'���Y�����(����F�х%>�V��#�c��?%�?��I��W>���U�[_��	��t����*�=�2 =&�Q����/ǈ��P>ē��?]2?D@?r ?�rO?@FI���Z���N�7���O5��ȼ>q?p7J>�+�> %�>k�0=���>'ob�����ώ�z�o>��b?EUM?�xs?"5��9�.��v�� �*�j�C��>þĉ>gO>�AW>@��ѯ���T���6��!q��;���O����0S�<Xa2?�A�>BU�>�Z�?��
?���QҪ���1��Y)��%;>��>�po?j�>�F>�ʙ�p�#�i��>O�l?U��>`�>����Y!���{��ʽ�'�>�ޭ>���>a�o>M�,��#\��i��փ���9�\^�=ɨh?���C�`��>�R?��:��G<$|�>j�v���!�]�򾔼'���>�|?���=��;>o�žB#�ؤ{��8��+)?.�?�	��P*�!�>��"?]6�>��>�ă?�2�>����&t;��?�]?QJ?�g@?	�>* =���ƾƽQk&���+=H��>�\>i}=|�=����Z����Y?=��=�ۼ�������;�k���y<�Z�<�3> ޿yO�wѾ�>����5��L��a�Ľ�؂�+:�H��x�������7�l!��� v�S a�maq���i�v��?��?oWR�aHP��뗿�)��t���8�>ẍ�;���꛾�4���|�������˹���[�Gea�zc���'?г��0�ǿ�����5ܾ�  ?�B ?%�y?�%�"�J�8�@� >��<Ͻ��]�뾀���K�ο����d�^?���>	�l8�����>���>��X>|Iq>����鞾��<�?x�-?A��>��r��ɿB���@��<���?�@G�=?.�����F��<V��>
�?�8i> �� ���֜�(��>q��?���?�e�<�bQ��"��o\?{Z���E�\g���r�=�n�=��=���R`{><!�>��QI�E�ʽ �,>�;�>G�N�xg>��~�D�w�Xi>���w���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=����Ϳ�*%�d�L�c4�; ۥ=��	=t��;��rZ��Cc��㘾(����ʄ�4ݥ�C,<�X�>ϗ>�A�>2�M?�h?�[�>i�U>��-��c��Ҹ������6��������X�]��i��!�޾pQ����3�n״���ǾfK;��K�=�R�r돿�a��a�J]E���-?ؿ%>�hɾ͞L���=<Ssɾ樮�(bI�����I�˾y92��-m�6B�?�@?�����W�ď��sҼ����W?���[H�-o��ޤ�=|����(=���>�\�=�\�?5�}�R���7?�?��پ�O��~'>�Oн�La>�4?SY�>jO���t>�iQ?�S�މ���0�>��*>�)l=��=]�7>|���8ͽ�3?� _?�@���6���w�>���/ɽ\	q=��1>bJ��BJA��Ɣ>:۸���о��9�븼+Iu��W?��>' ,����W���i�#�=0�q?[�?Ɵ>9�f?�@?���<Q����G�WG�@R =+�D?�a?�d>�H��پ�ಾ+�,?�Fg?��v>�xJ�뾳'�v���F�?Ro?v#?�x�R���0�������2?��v?ur^�`s��<��O�V�a<�>\�>.��>��9�4m�>ґ>? #��G�������Y4��?{�@t��?�;<;!����=�;?i\�>+�O�=?ƾ�z��V�����q=�"�>㍧�ev�$��DS,��8?���?D��>����3�����=Hې���?,ڊ?���|�<�{���c�����K����=B���O���xվ�/-�ߦ��ݲ��c�������̈́>~�@S���2�>����4鿦(ο��������O
?i��>u������dW��e��0��2��QB��ld>��D>�(�=�S���H��\kG�g>j��� ?x%����c>|�=j�@-�����=Z�<>-D?8��>OX>�sվ���?�xþSrֿGŢ�q�[���??#�?)�?�a?�U�>��ξϔľZ����f?LP ?�-H?M�^>�e�������j?`���U`��4�&HE�U>�"3?�B�>*�-�4�|=^>X��>h>�#/�Z�Ŀ�ٶ�����?��?���?lo����>^��?Ks+?oi��7��\��x�*���+��<A?�2>X���S�!�0=��ђ�ɼ
?�}0? {�d.�\�_?$�a�K�p���-�s�ƽ�ۡ>��0�f\�N�����Xe�
���@y����?L^�?g�?ٵ�� #�g6%?�>f����8Ǿ��<���>�(�>*N>.H_���u>����:�i	>���?�~�?Qj?���� ����U>�}?�-�>��?���=�?$�=Z����=7�>�Q>x,����>�cO?�W�>�jZ=��g]2�J�M�<]]�����#[9��Fh>�ob?�bB?"GP>�꯽�g���.��T����O=(�����<�3>=�=�;4>� ��ݾ��?�r���ؿj�� k'�K54?@��>��?H��ݴt��m��:_?�|�>�6�6,���%���;�N��?�E�?��?v�׾�@̼�
>��>�F�>�սI��������7>I�B?�(��D���o� �>���?�@%ծ?!i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?oQo���i�B>��?"������L��f?�
@u@a�^?*AQ߿�|����ӾѾ�5�=���=+kM>Mb��m�<\�!=?tR����dK'=�~d>���=}�)>SBG>YLw>�Ub>s�����)��㞿X&���HQ����5澤h'���
�᳚�g �(9��An¾�E���@"��Z��p/H�\��V���3>�3E?��??{�s?I;�>��=�&��>���1�g;�⬽���=ߝ�>O2?��@??i?GIb����g�ǩj�!k���2��8s�>�>a*�>n?t]�>�L�g��=`V>[f�>*=]���d�'>�E�NF>"ڹ>.�?d�>�O?>o�>r������~g�ϕt��[ŽT�?�:���~I��Q��#h���q�����=~t.?\>�ԑ�i@п�4����G?�����E�/�>� 1?�X?��>e���K~O�<>8 ��d�k�>�r�Ղq��)���I>� ?L�g>w�u>&�3�@8�vkP�6���y}>��5?w~��a�8�4�u�T�G�Biܾw�J>M�>9@�ӑ����֛~��~i��?z=�W:?�y?�.��?°��t������SR>B�[>W=���=	�M>N�`�ǽ��H��,=&@�=X�^>���>L[N>7u�=�WY>�E��<(���`�>2zl>�c>��G?��?����>�������(�>���>H��>�YO=�Ɇ���G=��>�,c>���=��<�P��:zh���> ږ�[T����rˏ=��˽.R)>�J2>��B�e���a>�~?���(䈿��e���lD?T+?U �=9�F<��"�C ���H��F�?r�@m�?��	��V�>�?�@�?��M��=}�>׫>�ξ�L��?��Ž6Ǣ�˔	�&)#�jS�?��?��/�Yʋ�9l�6>�^%?��ӾMh�>�x��Z�������u�ӷ#=W��>�8H?�V����O�X>��v
?�?�^�ݩ����ȿ:|v����>R�?���?b�m��A���@����>7��?�gY?noi>�g۾W`Z����>Ի@?�R?�>�9�b�'���?�޶?ԯ�?GI>c��?W�s?�i�>:�w��]/��7������$�=��N;tJ�>�x>�����dF��ӓ��^����j����C�a>+�$= �>AZ�	A���b�=V󋽱J����f����>�$q>8�I>�F�>�� ?�]�>���>��=9<��܀�������K?[��?z��?%n��q�<!��=��^�3?$D4?�"[���Ͼ��>�\?l��?�[?|U�>���0?���࿿�{��{*�<��K>�2�>�A�>x��AK>��Ծ|8D�qo�>Z֗>[���.@ھ����N��	7�>3d!?���>謮=�� ?��#?��j>(�>�_E�F9��P�E�۱�>آ�>�H?@�~?{�?�ӹ��[3�����塿�[��5N>��x?�U?3ɕ>k�������myE�6*I�^璽V��?9sg?:M�B?*2�?�??��A?�%f>\���ؾ%�����>
p?�i��)MV�~C$���\<@�"?\?}��>�S�M5r�s'>f?оd���;��>�Q?�8 ?6���N�O��H=vA���L������3=w��>M�>uh�6S�=��>��_=)1ս��+��Ũ��
!��w�>U?>���h��zL1?i��=C!��S�콐/����T���>~�>�s˾���?�:���&���Ø��#��}F����y?˳�?���?/޾�!d�	0.?jό?<�?;b?	{�����W�	�ʘz� T���1&���k>^?g�2��ӎ��)��XI���v���U�H����>l{�>�>?"�?Zp\>���>�ߚ���#�%?�\�{
\����3��H-�����*���a&��$����������i�>���ӭ�>�L?��`>k�~>�?�>��"�L�>��N>7#x>��>�Q>�6)>��=�\<H�ɽ�Q?��¾�R(�@��宾B?;d?U��>U�f��儿�����?Mv�?� �?Ot>�h�H�*�w(?���>,h~�+�	?�l@=�����<�����Z����O��/�>tW̽%:�C�L�n,e�D5?X?�<���̾x۽�����o=�O�?e�(?��)�3�Q�l�o�l�W�AS����Dh�{k���$���p��ꏿN\��G#���(�}l*=Ċ*?F�?����-��0%k��?��rf>p�>�>��>zcI>��	�?�1�� ^��D'�ܰ���K�>�U{?&ԃ>ͧG?�;?CF?RiD?*��>�O�>�;��58�>w��<!L�>f��>�DA?�$?� 1?ݯ?��'?�]>#����< �ݾ,?�/?T?p4?~h?�������@���h�<1a�u���=UD�<���� §����<�-n>Z�?Pm߾�{f�ޜ��w�>�:g?J$?��>#t˽��E=�N>��>k'
?��D>��D�T%|��B8��:&�� ?�{�W4��=Ŗa=A���:���\H=m���D�=����?Y�m��=aV���0���=�|�=N���[���Q���u�>��?���>AC�>�>��ǩ ����bd�=�Y>�S>�>�Dپ[}��	%����g�_ay>w�?�y�?�f=��=ē�=�~���W��2��J����(�<o�?!I#?XT?��?��=?wj#?W�>P+�M��q^�������?�+*??	�>���OؾF���� ;�l[
?e�?E�^�)���L�.���ľ3����=��0�<�r�������/��[Խ+q�� ��@��?��?Q�w<�.�^I�\���8S��դ/?Z��>]'�>
�?�{2�^4K�:o	��y>�<�>y+b?�q�>[iO?A
y?c�b?v>2g5��K��j����1м}ߊ=�E-?.y?I�?Z�{?27�>&=(>g�!���F-̾�5��D��ӓ��]�=��i>�A�>I�>���>N�=�F��·�C���=��)>�}�>��>$M�>k̓>΢`�b\P??��>s��?�I��h;�S��U퉺]L�?V�g?Zeb?.�=�]K�X�Y���7��C`=���?���?&T?�Q �;�>���=_���گ����>�S>p��>Yx�=	Us;֋>J�4>���>��r�-s�L3:���w����>u�6?0����ſ#�q�9Dr�LU��%�<�N��gCb�G���N�Y�y=�=�E���2��5���xZ�oO��^��w���O ��E�{�YC�>�W�=73�=9��=���<A�м���<G�E=��<10=�i�֤�<x�9�P�ڻ�����C���,Z<qK=�����˾�}?�9I?'�+?��C?��y>xI>%�3�B��>|���>?�V>�hP�������;�G����$��e�ؾv׾��c��̟��L>�eI���>�>3>]@�=���<R�=�1s=�ڎ=k�T��=�H�=EG�=DW�=���=��>�K>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>6�^>��>7NV�l�.��<��u:�U���?�/��Ķ��Ǉ>�>�¾l�ྴ�=�<<>!�;�f�q�O�+�=ӎ��:_<���<u�m>5GY>�`>�׎�F|v=#/=0^�=���>��A=����-X������dl=��6>\B>{�>P?1� ?�8w?g>�>�-;7��;���z�[>
I�� ,>BZ�=#�G�tU>o�l?T�6?��?�Y�>��w>W��>�X�>7�4���s��ƾhG��:- �up?��y?�o�>��q��P�u���ܜq��Tg�	"!?��?���>`��=�U����CY&���.�ވ���X2�/+=~mr��QU����m�!���=�p�>u��>��>,Ty>"�9>��N>�>��>^7�<mp�=G������<j�����=h���� �<�sż�����&���+�����5�;A��;��]<ĝ�;v4�=R:�>�>x��>�T�=�]��p�.>$Ӕ��L���=�R����A���b�f�}���.� Q5��FE>�Z>.���;��f~?�K\>@>��?V�t?dP>-=���Ծ�G����c��hP���=��>�7�N4:�Il`��M�`�ξ@��>V�>�'�>�5>��1���E��YP=��3@3�Թ�>����7I���0�_�o�gn��WD��{T���.=�'?q���^�=>�}?.5C?��?]d�>���HX�\�>>3�����=m��\U����[P*?�;0?�l�>R���ah�'�̾K־��K�>/�H�y�O�ɾ���0��C�F���"�>;J����о�3��C���돿ucB��r��Y�>_�O?��?=�a��R��2PO�7��[��O?܏g?�f�>=??L?c�����o��m��=��n?���?2�?͛
>Y+>z�5��)�>��?�H�?��?g8q?wЀ���>���=�F,>	�{�0�s��Ř>A/�<�]^�q7�>$�>���>����r������Ԅ<�M>�(�;���>%m�>v�!>	6�<d�f��i=@o6>�S0>��<��=ґ>��><���f?���?��>U�5>�6)?��>k->	�F>�)>7�=3����1�����~����E>�@e��B���m½�[�>����-��?�b�>eW��8;?��������>y�:j7�{2>o�6�%��>�~>8�;>��=�y*>H>	+Ӿ��>���a!�3 C��tR��ѾQrz>4�����%�8��k+��^)I��}���[�vj�P.���D=�Pֽ<WC�?9���w�k�/�)�����+�?�^�>�6?�ی�����>���>�ԍ>�4��슕��ɍ��n��	�?b��?��Y>�٧>�"f?�I-?�6���m�dPd��;n�*�<��tk�a�P��x���{��_�P���|`?�Gq?W�.?0�=Q�n>`�?�������U�>paS�u�J�� 8�c�>w��x���g;�����&?�`�S>��h?�Â?�?����l��'>V�:?֟1?�=t?��1?R�;?����$?��3>�>?yf?z@5?��.?��
?Ad1>� �=^����)'=�U��6&����ѽd�ʽ���n6=-�z=ޱ��
<j�=�ݧ<LQ�X߼�(;;������<��:=��=���=!˔>ݍ�?�&?|>�>�K"?ױɾSG��	>�M�C?�����9��%6�����۽I0�<څy?G�?�~?P&?�W"�oR��%>h��>��>��a>P8�>k�m����N[=*�->a^e��)གl1>����������̼�'�>��>nc|>�_����'>�}���uz��d>p�Q��ú�ПS���G���1�ʟu�+�>��K?4�?D�=z/�
���Df�])?G<?�9M?��?_��=
�۾>�9��J�{E��Q�>�Ы<���򶢿���i�:��9:
gs>/����I��.j>����ܾ�Uj��AG���⾐�K=���6�_=9�	���Ѿ�{�e��=�>�K���] �jm��d��K�H?��U=3V��yja��%��W/$>�^�>�"�>�{P��N[���<��Ƥ���=J��>�c1>#0�����mK�B���>�^E?�_?v�?�����#s��ZC����٧�����#)?���>g�?�A>�k�=�� ��Cd��F�B��>�c�>����YH������,��#'%����>lN?�>>�s?0S?n�
?�O_?�a)?��?���>馷��߷�_�"?ۤ�?^P�=+�l�\���1:�@8G��>T�$?{�m���\>2#?*?���>a�P?�$?|>($����&��C�>�>1�Z��~��:�k>��L?V�>�S?�v?�c>(�&�cK���<0�=��=G�,?g.?���><�>AL�>Zz���rW=[�>�ec?$�?��o?J��=�?44>��>2i�=�n�>�y�>s�?��M?H�q?a"I?�m�>�7�<�����}��Ʉm�O���z<���<�4}=F3���k���!��<�|�:���X�u�Y8%��ӼlV�;��>��t>�
��1�.>cGž����~@> ��3��*u���3;�g��=Z�>�?*�>W(!�P��=�>��>$���'?o�?�?0I�;&�a�F�پ��L�2��>��A?���=�l�����u�z�n=�Qn?e�]?2�Y�I���G�b?��]?�h�=���þ��b�8����O?��
?(�G���>��~?-�q?��>��e�l9n���jDb�N�j�'Ҷ=�q�>TX�8�d��>�>Z�7?VO�>:�b>&"�=�t۾��w��o���?@�?��?#��?8)*>`�n��3���6���x�c?�B ?�y���j/?P�f�����E�e�����׾ξqR��f̀��~���l��O�h�j���&w=��?��q?Tx?�c?���q�l�[�k��w�n��L#�i���D�-E�t�'���Y�����(����F�х%>�V��#�c��?%�?��I��W>���U�[_��	��t����*�=�2 =&�Q����/ǈ��P>ē��?]2?D@?r ?�rO?@FI���Z���N�7���O5��ȼ>q?p7J>�+�> %�>k�0=���>'ob�����ώ�z�o>��b?EUM?�xs?"5��9�.��v�� �*�j�C��>þĉ>gO>�AW>@��ѯ���T���6��!q��;���O����0S�<Xa2?�A�>BU�>�Z�?��
?���QҪ���1��Y)��%;>��>�po?j�>�F>�ʙ�p�#�i��>O�l?U��>`�>����Y!���{��ʽ�'�>�ޭ>���>a�o>M�,��#\��i��փ���9�\^�=ɨh?���C�`��>�R?��:��G<$|�>j�v���!�]�򾔼'���>�|?���=��;>o�žB#�ؤ{��8��+)?.�?�	��P*�!�>��"?]6�>��>�ă?�2�>����&t;��?�]?QJ?�g@?	�>* =���ƾƽQk&���+=H��>�\>i}=|�=����Z����Y?=��=�ۼ�������;�k���y<�Z�<�3> ޿yO�wѾ�>����5��L��a�Ľ�؂�+:�H��x�������7�l!��� v�S a�maq���i�v��?��?oWR�aHP��뗿�)��t���8�>ẍ�;���꛾�4���|�������˹���[�Gea�zc���'?г��0�ǿ�����5ܾ�  ?�B ?%�y?�%�"�J�8�@� >��<Ͻ��]�뾀���K�ο����d�^?���>	�l8�����>���>��X>|Iq>����鞾��<�?x�-?A��>��r��ɿB���@��<���?�@G�=?.�����F��<V��>
�?�8i> �� ���֜�(��>q��?���?�e�<�bQ��"��o\?{Z���E�\g���r�=�n�=��=���R`{><!�>��QI�E�ʽ �,>�;�>G�N�xg>��~�D�w�Xi>���w���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=����Ϳ�*%�d�L�c4�; ۥ=��	=t��;��rZ��Cc��㘾(����ʄ�4ݥ�C,<�X�>ϗ>�A�>2�M?�h?�[�>i�U>��-��c��Ҹ������6��������X�]��i��!�޾pQ����3�n״���ǾfK;��K�=�R�r돿�a��a�J]E���-?ؿ%>�hɾ͞L���=<Ssɾ樮�(bI�����I�˾y92��-m�6B�?�@?�����W�ď��sҼ����W?���[H�-o��ޤ�=|����(=���>�\�=�\�?5�}�R���7?�?��پ�O��~'>�Oн�La>�4?SY�>jO���t>�iQ?�S�މ���0�>��*>�)l=��=]�7>|���8ͽ�3?� _?�@���6���w�>���/ɽ\	q=��1>bJ��BJA��Ɣ>:۸���о��9�븼+Iu��W?��>' ,����W���i�#�=0�q?[�?Ɵ>9�f?�@?���<Q����G�WG�@R =+�D?�a?�d>�H��پ�ಾ+�,?�Fg?��v>�xJ�뾳'�v���F�?Ro?v#?�x�R���0�������2?��v?ur^�`s��<��O�V�a<�>\�>.��>��9�4m�>ґ>? #��G�������Y4��?{�@t��?�;<;!����=�;?i\�>+�O�=?ƾ�z��V�����q=�"�>㍧�ev�$��DS,��8?���?D��>����3�����=Hې���?,ڊ?���|�<�{���c�����K����=B���O���xվ�/-�ߦ��ݲ��c�������̈́>~�@S���2�>����4鿦(ο��������O
?i��>u������dW��e��0��2��QB��ld>��D>�(�=�S���H��\kG�g>j��� ?x%����c>|�=j�@-�����=Z�<>-D?8��>OX>�sվ���?�xþSrֿGŢ�q�[���??#�?)�?�a?�U�>��ξϔľZ����f?LP ?�-H?M�^>�e�������j?`���U`��4�&HE�U>�"3?�B�>*�-�4�|=^>X��>h>�#/�Z�Ŀ�ٶ�����?��?���?lo����>^��?Ks+?oi��7��\��x�*���+��<A?�2>X���S�!�0=��ђ�ɼ
?�}0? {�d.�\�_?$�a�K�p���-�s�ƽ�ۡ>��0�f\�N�����Xe�
���@y����?L^�?g�?ٵ�� #�g6%?�>f����8Ǿ��<���>�(�>*N>.H_���u>����:�i	>���?�~�?Qj?���� ����U>�}?�-�>��?���=�?$�=Z����=7�>�Q>x,����>�cO?�W�>�jZ=��g]2�J�M�<]]�����#[9��Fh>�ob?�bB?"GP>�꯽�g���.��T����O=(�����<�3>=�=�;4>� ��ݾ��?�r���ؿj�� k'�K54?@��>��?H��ݴt��m��:_?�|�>�6�6,���%���;�N��?�E�?��?v�׾�@̼�
>��>�F�>�սI��������7>I�B?�(��D���o� �>���?�@%ծ?!i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?oQo���i�B>��?"������L��f?�
@u@a�^?*AQ߿�|����ӾѾ�5�=���=+kM>Mb��m�<\�!=?tR����dK'=�~d>���=}�)>SBG>YLw>�Ub>s�����)��㞿X&���HQ����5澤h'���
�᳚�g �(9��An¾�E���@"��Z��p/H�\��V���3>�3E?��??{�s?I;�>��=�&��>���1�g;�⬽���=ߝ�>O2?��@??i?GIb����g�ǩj�!k���2��8s�>�>a*�>n?t]�>�L�g��=`V>[f�>*=]���d�'>�E�NF>"ڹ>.�?d�>�O?>o�>r������~g�ϕt��[ŽT�?�:���~I��Q��#h���q�����=~t.?\>�ԑ�i@п�4����G?�����E�/�>� 1?�X?��>e���K~O�<>8 ��d�k�>�r�Ղq��)���I>� ?L�g>w�u>&�3�@8�vkP�6���y}>��5?w~��a�8�4�u�T�G�Biܾw�J>M�>9@�ӑ����֛~��~i��?z=�W:?�y?�.��?°��t������SR>B�[>W=���=	�M>N�`�ǽ��H��,=&@�=X�^>���>L[N>7u�=�WY>�E��<(���`�>2zl>�c>��G?��?����>�������(�>���>H��>�YO=�Ɇ���G=��>�,c>���=��<�P��:zh���> ږ�[T����rˏ=��˽.R)>�J2>��B�e���a>�~?���(䈿��e���lD?T+?U �=9�F<��"�C ���H��F�?r�@m�?��	��V�>�?�@�?��M��=}�>׫>�ξ�L��?��Ž6Ǣ�˔	�&)#�jS�?��?��/�Yʋ�9l�6>�^%?��ӾMh�>�x��Z�������u�ӷ#=W��>�8H?�V����O�X>��v
?�?�^�ݩ����ȿ:|v����>R�?���?b�m��A���@����>7��?�gY?noi>�g۾W`Z����>Ի@?�R?�>�9�b�'���?�޶?ԯ�?GI>c��?W�s?�i�>:�w��]/��7������$�=��N;tJ�>�x>�����dF��ӓ��^����j����C�a>+�$= �>AZ�	A���b�=V󋽱J����f����>�$q>8�I>�F�>�� ?�]�>���>��=9<��܀�������K?[��?z��?%n��q�<!��=��^�3?$D4?�"[���Ͼ��>�\?l��?�[?|U�>���0?���࿿�{��{*�<��K>�2�>�A�>x��AK>��Ծ|8D�qo�>Z֗>[���.@ھ����N��	7�>3d!?���>謮=�� ?��#?��j>(�>�_E�F9��P�E�۱�>آ�>�H?@�~?{�?�ӹ��[3�����塿�[��5N>��x?�U?3ɕ>k�������myE�6*I�^璽V��?9sg?:M�B?*2�?�??��A?�%f>\���ؾ%�����>
p?�i��)MV�~C$���\<@�"?\?}��>�S�M5r�s'>f?оd���;��>�Q?�8 ?6���N�O��H=vA���L������3=w��>M�>uh�6S�=��>��_=)1ս��+��Ũ��
!��w�>U?>���h��zL1?i��=C!��S�콐/����T���>~�>�s˾���?�:���&���Ø��#��}F����y?˳�?���?/޾�!d�	0.?jό?<�?;b?	{�����W�	�ʘz� T���1&���k>^?g�2��ӎ��)��XI���v���U�H����>l{�>�>?"�?Zp\>���>�ߚ���#�%?�\�{
\����3��H-�����*���a&��$����������i�>���ӭ�>�L?��`>k�~>�?�>��"�L�>��N>7#x>��>�Q>�6)>��=�\<H�ɽ�Q?��¾�R(�@��宾B?;d?U��>U�f��儿�����?Mv�?� �?Ot>�h�H�*�w(?���>,h~�+�	?�l@=�����<�����Z����O��/�>tW̽%:�C�L�n,e�D5?X?�<���̾x۽�����o=�O�?e�(?��)�3�Q�l�o�l�W�AS����Dh�{k���$���p��ꏿN\��G#���(�}l*=Ċ*?F�?����-��0%k��?��rf>p�>�>��>zcI>��	�?�1�� ^��D'�ܰ���K�>�U{?&ԃ>ͧG?�;?CF?RiD?*��>�O�>�;��58�>w��<!L�>f��>�DA?�$?� 1?ݯ?��'?�]>#����< �ݾ,?�/?T?p4?~h?�������@���h�<1a�u���=UD�<���� §����<�-n>Z�?Pm߾�{f�ޜ��w�>�:g?J$?��>#t˽��E=�N>��>k'
?��D>��D�T%|��B8��:&�� ?�{�W4��=Ŗa=A���:���\H=m���D�=����?Y�m��=aV���0���=�|�=N���[���Q���u�>��?���>AC�>�>��ǩ ����bd�=�Y>�S>�>�Dپ[}��	%����g�_ay>w�?�y�?�f=��=ē�=�~���W��2��J����(�<o�?!I#?XT?��?��=?wj#?W�>P+�M��q^�������?�+*??	�>���OؾF���� ;�l[
?e�?E�^�)���L�.���ľ3����=��0�<�r�������/��[Խ+q�� ��@��?��?Q�w<�.�^I�\���8S��դ/?Z��>]'�>
�?�{2�^4K�:o	��y>�<�>y+b?�q�>[iO?A
y?c�b?v>2g5��K��j����1м}ߊ=�E-?.y?I�?Z�{?27�>&=(>g�!���F-̾�5��D��ӓ��]�=��i>�A�>I�>���>N�=�F��·�C���=��)>�}�>��>$M�>k̓>΢`�b\P??��>s��?�I��h;�S��U퉺]L�?V�g?Zeb?.�=�]K�X�Y���7��C`=���?���?&T?�Q �;�>���=_���گ����>�S>p��>Yx�=	Us;֋>J�4>���>��r�-s�L3:���w����>u�6?0����ſ#�q�9Dr�LU��%�<�N��gCb�G���N�Y�y=�=�E���2��5���xZ�oO��^��w���O ��E�{�YC�>�W�=73�=9��=���<A�м���<G�E=��<10=�i�֤�<x�9�P�ڻ�����C���,Z<qK=�����˾�}?�9I?'�+?��C?��y>xI>%�3�B��>|���>?�V>�hP�������;�G����$��e�ؾv׾��c��̟��L>�eI���>�>3>]@�=���<R�=�1s=�ڎ=k�T��=�H�=EG�=DW�=���=��>�K>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>6�^>��>7NV�l�.��<��u:�U���?�/��Ķ��Ǉ>�>�¾l�ྴ�=�<<>!�;�f�q�O�+�=ӎ��:_<���<u�m>5GY>�`>�׎�F|v=#/=0^�=���>��A=����-X������dl=��6>\B>{�>P?1� ?�8w?g>�>�-;7��;���z�[>
I�� ,>BZ�=#�G�tU>o�l?T�6?��?�Y�>��w>W��>�X�>7�4���s��ƾhG��:- �up?��y?�o�>��q��P�u���ܜq��Tg�	"!?��?���>`��=�U����CY&���.�ވ���X2�/+=~mr��QU����m�!���=�p�>u��>��>,Ty>"�9>��N>�>��>^7�<mp�=G������<j�����=h���� �<�sż�����&���+�����5�;A��;��]<ĝ�;v4�=R:�>�>x��>�T�=�]��p�.>$Ӕ��L���=�R����A���b�f�}���.� Q5��FE>�Z>.���;��f~?�K\>@>��?V�t?dP>-=���Ծ�G����c��hP���=��>�7�N4:�Il`��M�`�ξ@��>V�>�'�>�5>��1���E��YP=��3@3�Թ�>����7I���0�_�o�gn��WD��{T���.=�'?q���^�=>�}?.5C?��?]d�>���HX�\�>>3�����=m��\U����[P*?�;0?�l�>R���ah�'�̾K־��K�>/�H�y�O�ɾ���0��C�F���"�>;J����о�3��C���돿ucB��r��Y�>_�O?��?=�a��R��2PO�7��[��O?܏g?�f�>=??L?c�����o��m��=��n?���?2�?͛
>Y+>z�5��)�>��?�H�?��?g8q?wЀ���>���=�F,>	�{�0�s��Ř>A/�<�]^�q7�>$�>���>����r������Ԅ<�M>�(�;���>%m�>v�!>	6�<d�f��i=@o6>�S0>��<��=ґ>��><���f?���?��>U�5>�6)?��>k->	�F>�)>7�=3����1�����~����E>�@e��B���m½�[�>����-��?�b�>eW��8;?��������>y�:j7�{2>o�6�%��>�~>8�;>��=�y*>H>	+Ӿ��>���a!�3 C��tR��ѾQrz>4�����%�8��k+��^)I��}���[�vj�P.���D=�Pֽ<WC�?9���w�k�/�)�����+�?�^�>�6?�ی�����>���>�ԍ>�4��슕��ɍ��n��	�?b��?��Y>�٧>�"f?�I-?�6���m�dPd��;n�*�<��tk�a�P��x���{��_�P���|`?�Gq?W�.?0�=Q�n>`�?�������U�>paS�u�J�� 8�c�>w��x���g;�����&?�`�S>��h?�Â?�?����l��'>V�:?֟1?�=t?��1?R�;?����$?��3>�>?yf?z@5?��.?��
?Ad1>� �=^����)'=�U��6&����ѽd�ʽ���n6=-�z=ޱ��
<j�=�ݧ<LQ�X߼�(;;������<��:=��=���=!˔>ݍ�?�&?|>�>�K"?ױɾSG��	>�M�C?�����9��%6�����۽I0�<څy?G�?�~?P&?�W"�oR��%>h��>��>��a>P8�>k�m����N[=*�->a^e��)གl1>����������̼�'�>��>nc|>�_����'>�}���uz��d>p�Q��ú�ПS���G���1�ʟu�+�>��K?4�?D�=z/�
���Df�])?G<?�9M?��?_��=
�۾>�9��J�{E��Q�>�Ы<���򶢿���i�:��9:
gs>/���M���Qwb>���O�ݾ�)n���I�����UJ=�q��@Y=�����վ݂�+��=��>- ���� �	�����'
J?�j=�z����U��񺾲">��>��>��=�0�v��7@������=Y��>��:>~ɚ�!ﾅ0G�5&��&y>��B?>�b?
υ?��o���s���D����𸑾�:L���?��>���>��4>l�=����&�4]V�+�@���>p��>���@.A�ܵ���} �
�$��؀>�{?k+>�w?hVF?=��>MAW?:�0?�?� �>�x~��׼��&?�݃?Um�=>����P���7��K��0�>�/?�mU��G�>��?�O?e�?��T?D�?y�$> �N]:����>l��>�Y�|诿�%`>�I?~��>fZ?�2�?��C>o�2����x�0��=S9>�y6?�$?�c?�>y��>�n���g�=U��>>c?�(�?}�o?/��=F�?n�1>7��>�*�=u��>�P�>��?�4O?��s?z�J?&A�>�Ë<�t���޶��Is��SI�'|�;��I<��y=�]��v������<d�;qZ���6�����OB�i���A�;��>&N|>0��&/L>u��v���8>�Y�k ���拾�:����=�l>ve�>�n�>�F5�P�C=�~�>�'�>˂�4�(?�Y�>�n?gp��jUd�!7�J,l����>�@?��=�am������o�-J�=��i? \?��J�k��E�b?��]?vh�=���þN�b�<��N�O?��
?�G�/�>��~?h�q?��>��e�:n���Db�?�j��ж=er�>?X�L�d�Y?�>Y�7?�N�>�b>�&�=Tu۾�w��q��(?h�?��?���?�**>e�n�M4࿑:������"Z?O��>����j?��,�_�Ѿ�f��6�H��S��t��@Ae�Tf��쬾&�|�l����A����=rX?���?o\�?�Rh?pwپa�s��ʁ�@j��W�~iԾ�/��E��J�T04��]W�"�ξ�վ���폲<WW��Z� ���?�5?,g��p�W>]���@
�Ӡо��>v	��83��=Y;S���ڦ�=L =���
r!������J*?Ƿ?4�>I�4?E�C���j��Y�A;/�����<��>0�r>L�T> <漉ƻ<�>�g��F����\��Fx>{b?��L?l�n?O���f.�\���6 ��ټ�ԭ�=1>N��=G�>��E����mL"��p>���n��
�����d	��j=O�1?i9�>E�>��?q?�&�����m�Ǚ/���<갳>��e?4��>��>�5ϽCz$�V
�>��l?\��>��><	���� ���z�>Eν�X�>;̮>r��>�o>;U*���[�x0���r���9���=��g?�����:`��9�>@UQ?.��;GgO<6��>SWt��"�ui�RS#��}	>G�?t��=�P9>�Bž`�
�(�z�"Ԋ���(?';?Kۏ�=�(��|}>��!?x�>d�>�8�?��>e�ľ�E`���?~�^?�mI?t�@?�_�>XG=�*���E˽��'��%=��>��[>��s=݇�=��V�W���v8M=��=�j��݄����;
Jμ�T<7D�<\�+>
ۿ��K���վ)X��_�]��}T��O���釾ך�\��S7����u���
�Mk&�T`�1n�����Eg���?�-�?
�������l���������>��t��x`����2���u�� |�s���q* ���O��Di�B�d�=�$?\ޛ��vƿy����۩��'?��&?�7p?��
��T�]��b��=#��:�r<M]ξ����]l̿G���қP?-w�>���B��c�>o>�^[>�O>��������,�=A��>�.?��?ƫ~���Ŀ�Z����<N��?tE@YU<?��O�i����<?�"+?}e�>T��pH��)���??�ٞ?���?'\1��L�;?�(½f�8�ss'�'��=�_�=O2ݽϮ��p�>i�>� �,i�jY�n#�=��>��A]�ݎ��*�L=3Ɉ><1���-�Մ?�y\��f�x�/�TT���W>7�T?�)�>�2�=}�,?A6H�n|Ͽ�\�x'a?�0�?���?��(?�޿�&ך>t�ܾf�M?D6?���>ee&�r�t� ��=�/�ê��#�㾒&V�B��=Ԭ�>��>��,�ċ�/�O�$*��z��=�����Կ�)�C*��=�<a�N�O=�!��L��¿#�I��D����9k9>�>ռ=��<_s>DiK>�5J>�4E?�j?Z��>T?9>����&��Z�о�]�E%��X�1�^�������ٽ��m��̾���U} �]� ��y����;�Tg�=�R�Uʐ�l�!���b�پE�$0?: $>�
ʾ�rL���;-:˾̝��;0�������˾��.��`n�᝟?.IA?L+��MW�B��U��f=��5ZX?���j�Nì�80�=����=��>�.�=w���2��R��2?]#?�I��DI����=����V=��?Ь�>���>�ċ>*�?��8������e>UJ�>�נ>��>��<��Ⱦ���?#?�S?���[���i�>�žz���CuQ=��N=�(��V܉=���>�b�<����ޛ��*ә�h�=W;?��}>2$��a�N־륨�,�>Pʋ?.b�>�$_>�*X?eK?�=8����B���*��>�=BPc?R�:?�.*>a���j���xe���'?b�?x�>mdؽ�<�|'.�Y���<?*hs?�5?[�!���e��������0?Gu?��3�����'���þW�q>p�>�$?��$��-�>&V-?5��<�.���#���J�/�?h��?]�?�|�����[��=`#?.&�>B,����ܾ�3���9ھ�< >)?�Jƾ��h��6���`��e ?�T�?�:�>�A��f���6>d�����?�Á?�<��r�;=�(�%^�?w*�.dT=)G0��g����=�Ⱦ�t8�h1��g���+꿾�SO=�[�>fe@�L;�Q�>��h��{�Կ���̾�b��o�?��W>8�E�1Ā���A��D�g����,�؃�<�}>0e>�M�=�¾.������j�O?�~��Į%>ړB>i�ξW�����=|Ơ>F?m/d=�A�>�W��?��̾��ܿ�W¿/8��C�[?���?���?���>��3>��\�z
��TK�=��>?��>/��>�C�=�y>����j?�N��X`�U�4�>SE��U>�3?)h�>�-���|=�%>@��>R?>] /�2�ĿUԶ�չ�����?��?�g���> ~�?�n+?�`�73���W����*��`��?A?��1>A~����!��8=��Ԓ��
?9z0?���w*�\�_?'�a�M�p���-�y�ƽ�ۡ>��0��e\�uN�����Xe����@y����?M^�?g�?ڵ�� #�d6%?�>f����8Ǿ��<���>�(�>*N>cH_���u>����:�i	>���?�~�?Nj?���������U>	�}?<�>���?o�=.��>�f�=鎮��v ���>��=T?�`~?y�L?���>���=�i9��e/��AF� �P�ވ���B����>�`?:�K?��a>�#���O1�� �	Fн��.����/M?��DJ�L�ݽnR7>֛9>=�>MA�VkҾT�?7n��ؿ�j��=}'��34?ḃ>� ?h���t�ԏ�%=_?�u�>)6��+��]%��0=�r��?�E�?}�?#�׾�A̼>��>�I�>r�Խz��~����7>��B?�D����o��>	��?S�@�Ӯ?4i�)	?X�pQ��gr~�*��\7����=��7?(�1 {>���>��=sv�1�����s�3��>�>�?�x�?��>�l?�io���B�>2= Y�>��k?lg?I}�����B>��?4��4����X��f?��
@�n@&�^?C袿��ο7L���ܿ����H �=�b�=��@>��ܽQY�=��=[�<t��;�>.��>��1>R�Z>^@.>Zf:>�O>>2���&�h!���c��GO��!�?5	��SW��*
���v�.���/վ�����q�N���	���G�k����d�=��T?�
R?e�p?�l ?�`��@">����V>"=7��M2m=�n�>C�2?�VK?(�(?�=KꞾ�b��o�����!k���>F>?�>�.�>���>"=��%F>�=>T́>)">�o,=yX;l�
=��D>wU�>�l�>W��>>Q=>o�>�Ӵ��s��j�e���r�������?�3���7K�&���ZT��9���z�=�.?�>�d�� �ϿRͭ�ӉG?�����S���.�:�>�}.?zV?s$>a��8�W��>�Y
���q�o;�=V}��9�h��)���N>JX?d�x>�7[>.�9�_�;�4�:�����zx�>��-?Y�������c���7��ھ_$>�5�>]"�%#��1���Mx���x�O�>=�05?�
?�W�M�����c�����&N�>��Z>e�X��'==ɗE>J�����6G������>��>�G?U�>p��=v��>a4���
��C�>�v�=��>[�f?�>46��4G<�. ��g��uV�>7�>�M�=�A�<�����=m^�>�^�> �=�Tݽ������c�o�>��u�>j����� v�=r�>�����>������=y-�=�~?���(䈿��e���lD?S+?] �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��H��=}�>׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l�6>�^%?��Ӿ`�>���s���� ���-u�2=���>�MI?�Q��+2a�*z>�G�?�?	ﾫ��Hyɿ�u���>���?���?�mo�Կ�� >����>4�?]:V?&�e>}8ܾ`�W�'��>Lq@?��S?i��>B��<B)�j?�ô?O�?�'L>h�?�s?�%�>��w��-��Y��L��b�=��%<�-�>� >^���m�E��ɒ�����k����^>Z�=Y��>���Ϻ���=Ì�U쥾�(n���>"^n>+�O>�˜>G��>fk�>��>���<#ᄽ��u������K?X��?p���*n��a�<6��=Ԡ^�� ?�I4?��Y���Ͼ�Ѩ>��\?��?� [?fX�>���|:��C濿?}��Ɩ<�K> .�>M�>w%���KK>s�Ծ;D�Tj�>u֗>�֣��>ھ ��9��f8�>�e!?ʙ�>?��=�� ?��#??�j>@)�>�`E�48����E���>��>5I?�~?-�?,ѹ��X3�0��桿<�[��EN> �x?�T?�ʕ>?������.E��=I��󒽋��?Spg?S��?1�?a�??�A?%f><��O ؾ����M�>G�?�
?�"1f�����r> �?�6$?IP�>�滽4�G��$>;� �n����>��c?�j�>[�.��'i����~��<��k�>π�Z�����+�= ��=�>�<�+���3c>Vˈ>!}4���4��� =a�W=j�K>�9�=Y�	��6>�A$?��>�u���(���~�r�[�+lV>��>u���@q?YHk�o�U�|���x��]e��s`�?�+�?Aڑ?{E�a�y���	?@��?Ne0?�
?HZ���4����	�!.��x�j��t�Pp���{�>���=��S�􍐿V���s���=ϳK���?���>�?0��>�R>���>����ۇ��&����c���SF���־�)��Z#�����G��\`}�#=ӽ?w����Y�Gs>������>�:�>�1~>v�Y>�px>�H˽��>0Bx>��@>�0�>��=5�=�h>���=\F?��bH?��Ǿ��%��+Ѿ+�|��J?��e?�O�>�{B�������	��?��?���?�Hz>��l���2����>P��>!�K����>JJ��u�Pj��Ǿ�.����:�x���s>����k�6��R��M����?"?퇍�SԾN�������i=�t�?�)?I�(�A�Q�5�o���W���R����?%j�������$��No��|��0X���6����(�r*=�*?�ω?����
꾯�����l��A�7b>���>˨�>� �>�@I>a�
��,1�xj\�e%�s�����>�ky?�О>s99?��E?m]?`D?
^�>�Q�>�4ž~��>[�V��o>���>�Q?��+?;J�>
V�>��'?z��=o�ཚ��T^ྷ��>�7
?nj+?07
?���>�,l� \�e"�<j;p�
6��Z�=[MV>TF�=%����'����
�c�8=39?!\_�K{P�5
�SL�>��J?�?6��>��P�ֽĽOC�= J?�?�K7=�� �5�N��:��,>�lo?��W�R[=>�4>�*>��Z�Z��X��=q˒��p>{~=1�����C=x�>s�!��j7��b�=n�=�"1=�>�t�>"�?���>~@�>D��� �^���s�=Y>�S>i>,Fپ�}���#���g�@^y>{w�?{�?ˬf=��=���=d}��OT�����������<�?�H#?<VT?���?��=?�i#?�>�*��M���]��o��ݮ?�,?�c�>�����ʾ�Ϩ�%G3�.�?R?u$a�=#��)�:^¾�Խ�D>�8/��~�{����"D�1��5��<�����?��?wB�$�6�ld�����$��ȁC?���>^'�>/�>ۨ)���g�3���:>z�>�R?�>�>��S?bۃ? GQ?(�=>��2��Ь������G����$�
?!m?���?2/�?���>(c>y2-�&>��N^�Jp���-�=w�U�=7>C>���>$��>�}�>45=>˨�q`���!_�=y�=��>�A�>���>�K�>�-f>謃�wI?��?�;t�`���'W��12Q�O#X?W�?2�?���=��:�D��#�S�>��?VȨ?�&?)W�js�=�dŽ}ؾM��ں>�x�>v�>`f�=7wf��E�>�e�>b�>C�A��m=��^-�xT=���>���>+����ȿ�z�D���s��`�3<���{�Z�*c��4U���=�ڗ��{��ә���:�47���l���E������Po��<�>�A�=��>J�>@�=0����̻�T�<�{�;_��<��v�3�H=%��g�:��{�L?P���=г�=f�D��ɾ~7}?	I?��+?a�C?��z>X>	b:��y�>�����?�X>	H�.-��W�=��������4�׾��׾�fd�fx��{�>��G�`�>�-4>�f�=�x�<�D�=*5l=g;�=����=�
�=�|�= ��=QE�=�2>�]>w6w?隁�ղ���4Q��\�ܵ:?t8�>+}�=L�ƾ�@?��>>�2�������b�Y-?h��?�T�?!�?�ti�Nc�>����Ꮍ�t�=G����=2>��=��2���>9�J>@��K���}��D4�?��@/�??�ዿ��Ͽ�b/>:��>X�)>kf�J�a�B�ž�;����t�[?H3<� D���~�>���>�?��$o���\����7=���=�{ ;z/[�sbt=a��<�t=�>=\�>نT>\��=�$ɽk�>�>�ّ��t�>�o�D`Z�q�ý57#>�d�=DYg=ӳ!>�>��#?UO2?�st?���>������.����>x���5��>����Խ�e�>�![?�Z#?!D?E��>��h>���>3��>B%.���X��rľ>ž��x���Z?��u?֮G>1�)���O�~]��?���"=�*?@,H?�Z�>�"�>0�����%��g�W���!ŽpK=�͌����˹=/�?���s���=A�>鈨>Z� >ɸ>���>��y>�U�>^B�=ܯ�=�O�=�(�=Y^>�E�<�V#=Z�=X=�C�;ˆ>���*�����=�o<>u��=Ni:�����=��>�>Ƞ�>}����Ͼ�[>�rc��D��
>���r�=��xR��<p���p�Խf#�>p�f>G����폿�u�>
|F>$�t>~ڼ?Q�~?%!P>օ�����ZO��܅,����`>F�>y��YV��c�U;A��F��>��>�>m�>�@m>�+�<�>�ؼy=)�l15��K�>�~�����h�'q��+���럿�i�����._D?M2��m��=�}?�I?\�?{k�>o���*^ؾ�$/>:���pU=����_q�������?��&?]��>����D��J̾W����>z7I�3�O�NÕ���0��.��˷���>E�����о�%3��e��������B��Or���>��O?'�?�*b�V��zRO����FI��[m?F{g?��>�F?dB?���|�q��A��=V�n?f��?J=�?�
>X� >&��
��>h2?���?��?�h?}���+�>�cn��r�s�Q��4�>��>}��= ����>Aҝ>��>���� !��?-����H�1|�g��=�}�>I<�>�aA=*=C�B�^>�����=���>��>d(�A��>W>����nh�t}?��=)I}>�|5?uW�>=��=����2;�=v�+m��꙽W}X�y9 �F������t�==����0[�>K�ĿJ��?6CL>�� ��k"?ޖ�	ƽ���=,�|>��6��^�>Ȇ>Yn>�{�>	�>��=�$;>
�@>|�Ҿ�]>����!��+C��cR�tѾ50{>���x�%��l�5�����I��#���a�e�i��$����<��j�<9�?J�����k�X�)�U ����?KZ�>f6?�ی�����"9>��>Rҍ>{'������6č�--����?9��?b�h>%\�>�Ye?a�?��8��oa�	�q���s�K�W�V\^���Y�"����X�#�޾9Q���)V?K;�?��&?��	>/a]>-}�?���8��Q�>�~A���E�A�ȼF
�>+�߾��S�R3��$�ܾ��o�>e�h?`6�?��'?�^A�4	��YG>˩@?<8?��f?nF-?ͺ)?M=��/?�"=�q�>�m?j�7?�>!?���>��=�=���[څ=������u����W�_��4�KJ�<�-�=�}b��~�u�>�$g>͟D��j�r�����Q=�����P)<A�=�DF=�B�>��_??r7�>�
?y�ΩY���Ͼ$a�>n���+�o+�i:`�:�����i>o��?)�?"�?��?�N[�-�l��x>q,>@�>���>zl�>�C��fG���>6Ҩ=?�=EB���5"=���ޤؾ����M�d�9�>�v>�e�~]0>�<��y�u��$]>G�Q�����5_�WtH���1��}t��I�>�?J?�L?1H�=��澾*|��e��d&?>�9?�jL?z.~?Ǭ�=��Ծ�>8��F��.�w��>ٙ�<����2��ѿ��7;��<;;�q>�K���I��.j>����ܾ�Uj��AG���⾐�K=���6�_=9�	���Ѿ�{�e��=�>�K���] �jm��d��K�H?��U=3V��yja��%��W/$>�^�>�"�>�{P��N[���<��Ƥ���=J��>�c1>#0�����mK�B���>�^E?�_?v�?�����#s��ZC����٧�����#)?���>g�?�A>�k�=�� ��Cd��F�B��>�c�>����YH������,��#'%����>lN?�>>�s?0S?n�
?�O_?�a)?��?���>馷��߷�_�"?ۤ�?^P�=+�l�\���1:�@8G��>T�$?{�m���\>2#?*?���>a�P?�$?|>($����&��C�>�>1�Z��~��:�k>��L?V�>�S?�v?�c>(�&�cK���<0�=��=G�,?g.?���><�>AL�>Zz���rW=[�>�ec?$�?��o?J��=�?44>��>2i�=�n�>�y�>s�?��M?H�q?a"I?�m�>�7�<�����}��Ʉm�O���z<���<�4}=F3���k���!��<�|�:���X�u�Y8%��ӼlV�;��>��t>�
��1�.>cGž����~@> ��3��*u���3;�g��=Z�>�?*�>W(!�P��=�>��>$���'?o�?�?0I�;&�a�F�پ��L�2��>��A?���=�l�����u�z�n=�Qn?e�]?2�Y�I���G�b?��]?�h�=���þ��b�8����O?��
?(�G���>��~?-�q?��>��e�l9n���jDb�N�j�'Ҷ=�q�>TX�8�d��>�>Z�7?VO�>:�b>&"�=�t۾��w��o���?@�?��?#��?8)*>`�n��3���6���x�c?�B ?�y���j/?P�f�����E�e�����׾ξqR��f̀��~���l��O�h�j���&w=��?��q?Tx?�c?���q�l�[�k��w�n��L#�i���D�-E�t�'���Y�����(����F�х%>�V��#�c��?%�?��I��W>���U�[_��	��t����*�=�2 =&�Q����/ǈ��P>ē��?]2?D@?r ?�rO?@FI���Z���N�7���O5��ȼ>q?p7J>�+�> %�>k�0=���>'ob�����ώ�z�o>��b?EUM?�xs?"5��9�.��v�� �*�j�C��>þĉ>gO>�AW>@��ѯ���T���6��!q��;���O����0S�<Xa2?�A�>BU�>�Z�?��
?���QҪ���1��Y)��%;>��>�po?j�>�F>�ʙ�p�#�i��>O�l?U��>`�>����Y!���{��ʽ�'�>�ޭ>���>a�o>M�,��#\��i��փ���9�\^�=ɨh?���C�`��>�R?��:��G<$|�>j�v���!�]�򾔼'���>�|?���=��;>o�žB#�ؤ{��8��+)?.�?�	��P*�!�>��"?]6�>��>�ă?�2�>����&t;��?�]?QJ?�g@?	�>* =���ƾƽQk&���+=H��>�\>i}=|�=����Z����Y?=��=�ۼ�������;�k���y<�Z�<�3> ޿yO�wѾ�>����5��L��a�Ľ�؂�+:�H��x�������7�l!��� v�S a�maq���i�v��?��?oWR�aHP��뗿�)��t���8�>ẍ�;���꛾�4���|�������˹���[�Gea�zc���'?г��0�ǿ�����5ܾ�  ?�B ?%�y?�%�"�J�8�@� >��<Ͻ��]�뾀���K�ο����d�^?���>	�l8�����>���>��X>|Iq>����鞾��<�?x�-?A��>��r��ɿB���@��<���?�@G�=?.�����F��<V��>
�?�8i> �� ���֜�(��>q��?���?�e�<�bQ��"��o\?{Z���E�\g���r�=�n�=��=���R`{><!�>��QI�E�ʽ �,>�;�>G�N�xg>��~�D�w�Xi>���w���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=����Ϳ�*%�d�L�c4�; ۥ=��	=t��;��rZ��Cc��㘾(����ʄ�4ݥ�C,<�X�>ϗ>�A�>2�M?�h?�[�>i�U>��-��c��Ҹ������6��������X�]��i��!�޾pQ����3�n״���ǾfK;��K�=�R�r돿�a��a�J]E���-?ؿ%>�hɾ͞L���=<Ssɾ樮�(bI�����I�˾y92��-m�6B�?�@?�����W�ď��sҼ����W?���[H�-o��ޤ�=|����(=���>�\�=�\�?5�}�R���7?�?��پ�O��~'>�Oн�La>�4?SY�>jO���t>�iQ?�S�މ���0�>��*>�)l=��=]�7>|���8ͽ�3?� _?�@���6���w�>���/ɽ\	q=��1>bJ��BJA��Ɣ>:۸���о��9�븼+Iu��W?��>' ,����W���i�#�=0�q?[�?Ɵ>9�f?�@?���<Q����G�WG�@R =+�D?�a?�d>�H��پ�ಾ+�,?�Fg?��v>�xJ�뾳'�v���F�?Ro?v#?�x�R���0�������2?��v?ur^�`s��<��O�V�a<�>\�>.��>��9�4m�>ґ>? #��G�������Y4��?{�@t��?�;<;!����=�;?i\�>+�O�=?ƾ�z��V�����q=�"�>㍧�ev�$��DS,��8?���?D��>����3�����=Hې���?,ڊ?���|�<�{���c�����K����=B���O���xվ�/-�ߦ��ݲ��c�������̈́>~�@S���2�>����4鿦(ο��������O
?i��>u������dW��e��0��2��QB��ld>��D>�(�=�S���H��\kG�g>j��� ?x%����c>|�=j�@-�����=Z�<>-D?8��>OX>�sվ���?�xþSrֿGŢ�q�[���??#�?)�?�a?�U�>��ξϔľZ����f?LP ?�-H?M�^>�e�������j?`���U`��4�&HE�U>�"3?�B�>*�-�4�|=^>X��>h>�#/�Z�Ŀ�ٶ�����?��?���?lo����>^��?Ks+?oi��7��\��x�*���+��<A?�2>X���S�!�0=��ђ�ɼ
?�}0? {�d.�\�_?$�a�K�p���-�s�ƽ�ۡ>��0�f\�N�����Xe�
���@y����?L^�?g�?ٵ�� #�g6%?�>f����8Ǿ��<���>�(�>*N>.H_���u>����:�i	>���?�~�?Qj?���� ����U>�}?�-�>��?���=�?$�=Z����=7�>�Q>x,����>�cO?�W�>�jZ=��g]2�J�M�<]]�����#[9��Fh>�ob?�bB?"GP>�꯽�g���.��T����O=(�����<�3>=�=�;4>� ��ݾ��?�r���ؿj�� k'�K54?@��>��?H��ݴt��m��:_?�|�>�6�6,���%���;�N��?�E�?��?v�׾�@̼�
>��>�F�>�սI��������7>I�B?�(��D���o� �>���?�@%ծ?!i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?oQo���i�B>��?"������L��f?�
@u@a�^?*AQ߿�|����ӾѾ�5�=���=+kM>Mb��m�<\�!=?tR����dK'=�~d>���=}�)>SBG>YLw>�Ub>s�����)��㞿X&���HQ����5澤h'���
�᳚�g �(9��An¾�E���@"��Z��p/H�\��V���3>�3E?��??{�s?I;�>��=�&��>���1�g;�⬽���=ߝ�>O2?��@??i?GIb����g�ǩj�!k���2��8s�>�>a*�>n?t]�>�L�g��=`V>[f�>*=]���d�'>�E�NF>"ڹ>.�?d�>�O?>o�>r������~g�ϕt��[ŽT�?�:���~I��Q��#h���q�����=~t.?\>�ԑ�i@п�4����G?�����E�/�>� 1?�X?��>e���K~O�<>8 ��d�k�>�r�Ղq��)���I>� ?L�g>w�u>&�3�@8�vkP�6���y}>��5?w~��a�8�4�u�T�G�Biܾw�J>M�>9@�ӑ����֛~��~i��?z=�W:?�y?�.��?°��t������SR>B�[>W=���=	�M>N�`�ǽ��H��,=&@�=X�^>���>L[N>7u�=�WY>�E��<(���`�>2zl>�c>��G?��?����>�������(�>���>H��>�YO=�Ɇ���G=��>�,c>���=��<�P��:zh���> ږ�[T����rˏ=��˽.R)>�J2>��B�e���a>�~?���(䈿��e���lD?T+?U �=9�F<��"�C ���H��F�?r�@m�?��	��V�>�?�@�?��M��=}�>׫>�ξ�L��?��Ž6Ǣ�˔	�&)#�jS�?��?��/�Yʋ�9l�6>�^%?��ӾMh�>�x��Z�������u�ӷ#=W��>�8H?�V����O�X>��v
?�?�^�ݩ����ȿ:|v����>R�?���?b�m��A���@����>7��?�gY?noi>�g۾W`Z����>Ի@?�R?�>�9�b�'���?�޶?ԯ�?GI>c��?W�s?�i�>:�w��]/��7������$�=��N;tJ�>�x>�����dF��ӓ��^����j����C�a>+�$= �>AZ�	A���b�=V󋽱J����f����>�$q>8�I>�F�>�� ?�]�>���>��=9<��܀�������K?[��?z��?%n��q�<!��=��^�3?$D4?�"[���Ͼ��>�\?l��?�[?|U�>���0?���࿿�{��{*�<��K>�2�>�A�>x��AK>��Ծ|8D�qo�>Z֗>[���.@ھ����N��	7�>3d!?���>謮=�� ?��#?��j>(�>�_E�F9��P�E�۱�>آ�>�H?@�~?{�?�ӹ��[3�����塿�[��5N>��x?�U?3ɕ>k�������myE�6*I�^璽V��?9sg?:M�B?*2�?�??��A?�%f>\���ؾ%�����>
p?�i��)MV�~C$���\<@�"?\?}��>�S�M5r�s'>f?оd���;��>�Q?�8 ?6���N�O��H=vA���L������3=w��>M�>uh�6S�=��>��_=)1ս��+��Ũ��
!��w�>U?>���h��zL1?i��=C!��S�콐/����T���>~�>�s˾���?�:���&���Ø��#��}F����y?˳�?���?/޾�!d�	0.?jό?<�?;b?	{�����W�	�ʘz� T���1&���k>^?g�2��ӎ��)��XI���v���U�H����>l{�>�>?"�?Zp\>���>�ߚ���#�%?�\�{
\����3��H-�����*���a&��$����������i�>���ӭ�>�L?��`>k�~>�?�>��"�L�>��N>7#x>��>�Q>�6)>��=�\<H�ɽ�Q?��¾�R(�@��宾B?;d?U��>U�f��儿�����?Mv�?� �?Ot>�h�H�*�w(?���>,h~�+�	?�l@=�����<�����Z����O��/�>tW̽%:�C�L�n,e�D5?X?�<���̾x۽�����o=�O�?e�(?��)�3�Q�l�o�l�W�AS����Dh�{k���$���p��ꏿN\��G#���(�}l*=Ċ*?F�?����-��0%k��?��rf>p�>�>��>zcI>��	�?�1�� ^��D'�ܰ���K�>�U{?&ԃ>ͧG?�;?CF?RiD?*��>�O�>�;��58�>w��<!L�>f��>�DA?�$?� 1?ݯ?��'?�]>#����< �ݾ,?�/?T?p4?~h?�������@���h�<1a�u���=UD�<���� §����<�-n>Z�?Pm߾�{f�ޜ��w�>�:g?J$?��>#t˽��E=�N>��>k'
?��D>��D�T%|��B8��:&�� ?�{�W4��=Ŗa=A���:���\H=m���D�=����?Y�m��=aV���0���=�|�=N���[���Q���u�>��?���>AC�>�>��ǩ ����bd�=�Y>�S>�>�Dپ[}��	%����g�_ay>w�?�y�?�f=��=ē�=�~���W��2��J����(�<o�?!I#?XT?��?��=?wj#?W�>P+�M��q^�������?�+*??	�>���OؾF���� ;�l[
?e�?E�^�)���L�.���ľ3����=��0�<�r�������/��[Խ+q�� ��@��?��?Q�w<�.�^I�\���8S��դ/?Z��>]'�>
�?�{2�^4K�:o	��y>�<�>y+b?�q�>[iO?A
y?c�b?v>2g5��K��j����1м}ߊ=�E-?.y?I�?Z�{?27�>&=(>g�!���F-̾�5��D��ӓ��]�=��i>�A�>I�>���>N�=�F��·�C���=��)>�}�>��>$M�>k̓>΢`�b\P??��>s��?�I��h;�S��U퉺]L�?V�g?Zeb?.�=�]K�X�Y���7��C`=���?���?&T?�Q �;�>���=_���گ����>�S>p��>Yx�=	Us;֋>J�4>���>��r�-s�L3:���w����>u�6?0����ſ#�q�9Dr�LU��%�<�N��gCb�G���N�Y�y=�=�E���2��5���xZ�oO��^��w���O ��E�{�YC�>�W�=73�=9��=���<A�м���<G�E=��<10=�i�֤�<x�9�P�ڻ�����C���,Z<qK=�����˾�}?�9I?'�+?��C?��y>xI>%�3�B��>|���>?�V>�hP�������;�G����$��e�ؾv׾��c��̟��L>�eI���>�>3>]@�=���<R�=�1s=�ڎ=k�T��=�H�=EG�=DW�=���=��>�K>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>6�^>��>7NV�l�.��<��u:�U���?�/��Ķ��Ǉ>�>�¾l�ྴ�=�<<>!�;�f�q�O�+�=ӎ��:_<���<u�m>5GY>�`>�׎�F|v=#/=0^�=���>��A=����-X������dl=��6>\B>{�>P?1� ?�8w?g>�>�-;7��;���z�[>
I�� ,>BZ�=#�G�tU>o�l?T�6?��?�Y�>��w>W��>�X�>7�4���s��ƾhG��:- �up?��y?�o�>��q��P�u���ܜq��Tg�	"!?��?���>`��=�U����CY&���.�ވ���X2�/+=~mr��QU����m�!���=�p�>u��>��>,Ty>"�9>��N>�>��>^7�<mp�=G������<j�����=h���� �<�sż�����&���+�����5�;A��;��]<ĝ�;v4�=R:�>�>x��>�T�=�]��p�.>$Ӕ��L���=�R����A���b�f�}���.� Q5��FE>�Z>.���;��f~?�K\>@>��?V�t?dP>-=���Ծ�G����c��hP���=��>�7�N4:�Il`��M�`�ξ@��>V�>�'�>�5>��1���E��YP=��3@3�Թ�>����7I���0�_�o�gn��WD��{T���.=�'?q���^�=>�}?.5C?��?]d�>���HX�\�>>3�����=m��\U����[P*?�;0?�l�>R���ah�'�̾K־��K�>/�H�y�O�ɾ���0��C�F���"�>;J����о�3��C���돿ucB��r��Y�>_�O?��?=�a��R��2PO�7��[��O?܏g?�f�>=??L?c�����o��m��=��n?���?2�?͛
>Y+>z�5��)�>��?�H�?��?g8q?wЀ���>���=�F,>	�{�0�s��Ř>A/�<�]^�q7�>$�>���>����r������Ԅ<�M>�(�;���>%m�>v�!>	6�<d�f��i=@o6>�S0>��<��=ґ>��><���f?���?��>U�5>�6)?��>k->	�F>�)>7�=3����1�����~����E>�@e��B���m½�[�>����-��?�b�>eW��8;?��������>y�:j7�{2>o�6�%��>�~>8�;>��=�y*>H>	+Ӿ��>���a!�3 C��tR��ѾQrz>4�����%�8��k+��^)I��}���[�vj�P.���D=�Pֽ<WC�?9���w�k�/�)�����+�?�^�>�6?�ی�����>���>�ԍ>�4��슕��ɍ��n��	�?b��?��Y>�٧>�"f?�I-?�6���m�dPd��;n�*�<��tk�a�P��x���{��_�P���|`?�Gq?W�.?0�=Q�n>`�?�������U�>paS�u�J�� 8�c�>w��x���g;�����&?�`�S>��h?�Â?�?����l��'>V�:?֟1?�=t?��1?R�;?����$?��3>�>?yf?z@5?��.?��
?Ad1>� �=^����)'=�U��6&����ѽd�ʽ���n6=-�z=ޱ��
<j�=�ݧ<LQ�X߼�(;;������<��:=��=���=!˔>ݍ�?�&?|>�>�K"?ױɾSG��	>�M�C?�����9��%6�����۽I0�<څy?G�?�~?P&?�W"�oR��%>h��>��>��a>P8�>k�m����N[=*�->a^e��)གl1>����������̼�'�>��>nc|>�_����'>�}���uz��d>p�Q��ú�ПS���G���1�ʟu�+�>��K?4�?D�=z/�
���Df�])?G<?�9M?��?_��=
�۾>�9��J�{E��Q�>�Ы<���򶢿���i�:��9:
gs>/����/���Q�>�!���V������^��"'�O)��r��Ǎ=��F��)��#5콄��<3E#�J�1�3��K녿����&Ld?�f	>���h����ľH�=g�=��>�h]<��>��/�jʟ��۽=�
�>�T?C��>T"׾��O�����Ɗ>hP=?7RV?�2V?����xP���<�3�ԾX�����k&�>Nj�>G'>:'�>�z>6�4� ]*���v�Cm,�o��>O%?eԾi�=��Ϭ����E?O�d��> �?s������>�CC??��>@G:?DX2?U�>o@�>`�����$? _�?L�">	�0��D!��-?�?_[��l�>�� ?֣T�0X<d"�>�b�>���>�M?�u8?Y�<�(!�}�<�O�>2ؘ>I�5�އ��G�0��>�-�>?-$?E��?z&�>�!A�wf��>3�R���%�P?�?Ģ?���>μ�>Ώ��QY>�*T>�y?/ۉ?��>?���=�)�>��f>+T�>m��|��=l��>�!�>��?�6y?�[?��?�������kt]>�� =V��-3��	�e�a>*��<]C��C���:�<  C���;���:X=� ,�;"'A�bɻ����>��^>6'��s�5>'��'/����c>�w��	���7�_���L�_��=o}~>�4?��>��2�>3\�>��>&��	*?�?�J?�a�?e�&Y��@R�{�>��!?�<6Kq�{����\`�n3(=�s^?�Of?V���l�2�b?u�]?�e�=���þL�b�+����O?�
?��G���>��~?�q?���>��e�E8n�����Eb���j���=�s�>�T��d��9�>O�7?�N�>;�b>��=�z۾j�w�de��?��?1�?m��?6*>��n��1�V�����)P?�P�>�d���$?����B�����?��NȾ|�������
G���|��2(�'��qS���>F5?��q?�8r?N?;n�~�d��`f�і�,U��E��	�qoJ�A�4�`�A�gi���	�U�	��H���͋<�>���3��`�?u�-?�=��>�d����
]��(�>�8m�+��~=��@��=�y>�d���6-�P�R���?�	�>��>�1(?��M��hF�֪&���5����A��=��>A�>l��>:U�<ȏ+��1)����*_�� ����>�mX?�� ?r,e?�<�^�J��3����о�fW���ھ!_�<,;�>1@�>���99�8�.��L?��Pm��9'�r򒾓7��Q�=��1?�t�>R=�>ڭ�?#�?�h����
�̎n�G"�������>��a?�h�>�G>i�f��tھ8��>רl?���>8��>�狾 � �{{�Ͻ���>�ҭ>;i�>6�m>8�-�F\��)�����E�8�\��=lh?{S���$a�1X�>@R?$_
;d�D<1T�>d�v�^�!�����"'�p�>^�?�P�=W(<>sOž9��� {�����8'?T�?��|�ǳ'�
�}>U�?���>�7�>a��?_z�>l���,�O�?��R?ZM=?�E?ޮ�>*�/=ݾ���H˽��=���f=�ւ>�=l>�p�=B>���f>����|=���=�6̼�ν�-ż��t����<K�&=�7>Kaۿ<>K��پS����08
����֑��`w����!B�����x�����'��-V�t~c�䐌�3�l��v�?s;�?�q���3��A���ĕ�����x�>W�q�������z��*��l]����V!� �O��/i�|�e��'?���q�ǿ㥡��1ܾ�" ?�O ?��y?p�Ս"�r8�
� >�c�<j���nq�����t�ο��^?r��>��c����>辂>.�X>J/q>!@��_鞾^��<��?u�-?F��>��r��ɿ7���c�<���?5�@)@?�%����~=���>E�?�d>_M�(��k�����>u��?�%�?�Q=-~J��K2��d?5|_=H\7��b�hI>)��=�j!==����=0�t>���V�Z���&��?�=�0e>��v����tzd�@�FL�>k����&Մ?�z\�2f�p�/��T���T>|�T?�+�>�>�=ò,?H7H�U}Ͽԯ\�D*a?�0�?٦�?��(?0ۿ��ؚ>A�ܾM�M?�C6?���>�d&���t����=�4ἀE��$��f&V�c��=S��>>�>�,�֋���O��F�����=a���տV����]�֏i<u�%��6�=t:�t�侊���]�=��	����>�t7?���UX�L�?yX?��G�_�A?~<X?'�=��>|��<PR�3Ӿ�ѯ��K�"�t=qݽu�j�zξm{����������V����-�t���]��B�D�۳��zh��B��,� �"?� ����-�%YT>*9�=�8Q�au��ߦH��!��U
��֟|�Mʎ?nJ?T����h/���8�`^���<>��J?��C�_��/�y���H>�>v�>]d�=*���L�<��kn�5U/?~�?�浾�<���&>���$i"=�%?j�?�Ƅ<���>�K!?f2�g���BW>�vH>丟>�Y�>�,>�Ī�� �?�P?�e��ᐾ�>Nž��{���*=@>'R2�
���|rY>CF��≾%1�9E�\����<�N?�n>��'�-�Oꅾ�1E=�{b>��W?�	?���>�a�?�g=?9ʼ��
�Ph%��������pG?�J�?l[�=������ξW%��{jB?4f?��
>�U˾l��$ ���̾A?�^j?я?�x��*���2���羈F8?��v?�r^�ns��|����V�=�>E\�>��>��9�&l�>Ǒ>?~#�tG������Y4��?x�@���?[�;<<�ǝ�=�;?&\�>&�O��?ƾ�~��������q=_!�>̍���ev�����P,��8?���?;��>󒂾���]>�T��lI�?��|?�P��'Q<Op!�3>�i�����<�v>\��(�L��㾱9 �[��w�0�����ij:=~>�@|ڈ��k�>+���<ܿd+ſ(���;������>[�>��#�+�3��I;�r�T���/�i�e�ERҾ���>j= > ���r�z�ab~��A<�X�ϼ�s�>����͒>�dv�)���ڏ���=��$ۏ>(5�>�,e>~B併ٻ�p��?��c�ʿX���k
�I�P?FD�?�s�?�`?qi�;�:��vL����<?�|?�a?q�Y��&]�JR�{�j?0_���U`��4��?E��U>�$3?�6�>9�-�\}=S>���>�j>	/�-�ĿY׶��������?+��?j꾴��>��?ho+?h��8��j��#�*�W�C�~/A?	�1>H���^�!��'=�;Ӓ�m�
?�0?�R�n1�\�_?)�a�K�p���-���ƽ�ۡ>��0��e\��M�����Xe����@y����?M^�?h�?۵�� #�h6%?�>c����8Ǿ>�<���>�(�>*N>ZH_���u>����:�i	>���?�~�?Sj?���������U>�}?@�>���?�?�=;s�>���=R�������#>�B�=�wJ�?�eO?���>���=%o5���.�W�E�!�R��P	�$B�*>Za?sK?p�e>I���
�%��x�ҐĽ��6�������:���0��ϽK>9>A�9>�>w�@��4Ͼ�W�>T#;�� �k��FKٽ�;?ͽ�>�'�>�5#�Ud��l�=�sP?���>p�ǝ��<���9Ɯ�f�?���?��?̲��X�=�>�"�>m19>�ؽS� ��G��LT�=��-?V��������8���0>Rg�?6X�?���?4=Q��	?���P��`a~���[7����=��7?�0���z>��> �=�nv�ӻ��`�s�y��>�B�?�{�?���>�l?w�o��B�i�1=�L�>��k?�s?\Wo����B>��?�����-L��f?�
@vu@E�^?"��п�l��g���=�v�F�cp.>�M�=C�;=�F�;�T!�p}�=�E�=��)>�4�>�$n=X)A>O�Q>�z>/>S���p)�i����H��������;����:��^0�΋�'��]Q���6;�W*����K����������=:?���>�->?8q/?�Fe?+��>����D�,=�^��3G��N(��%|�!��>�?�B?�6%?�h%�cV��` _��Ro��Ҭ��zξ��>��6>��	?B??0��>�ҷ��*�>ߖ>]�>}�:'��F��<���3Si>���>c@�>)?2T<>|�>�Ŵ���Q�h��w�U�ͽ5�?�����J�$/��ʌ�	����̞=R.?�>����8пz���/H?����"�:�+��>��0?�iW?�>9Y��SNW��>;@�ݘj��>�@��llk��V)���P>�O?��g>dw>?3��X7���P��/���u>C�5?���9�8�'Su��}F�59۾�J>�C�>��W�A�Tݖ�6=�=�g�Z2y=K>:?��?.���v��R�r�'���@S>��Y>�=���=�
N>��X��jŽ��E�� =+G�=|�_>��>X	>���= O�>�:��a=��=��>hJ�%9>��?P�?�?�ǖ6��u���ȼb��>�H�>��>�7�>���!�V>� ?��L>���$߽�ʄ��^��n9<�5���]��:��R�E<�D
��Z�=֮���w��\/�$Ro��~?���(䈿��
e���lD?T+?U �=7�F<��"�D ���H��F�?q�@m�?��	�ޢV�A�?�@�?��O��=}�>׫>�ξ�L��?��Ž8Ǣ�ʔ	�6)#�iS�?��?��/�Zʋ�=l��6>�^%? �Ӿ�c�>��Z�������u���#=���>�7H?�W��E�O��>��v
?�?9[�򩤿u�ȿ�zv����>Y�?q��?5�m��A��|@�ރ�>ޢ�?�gY?fmi>�g۾baZ�ي�>��@?R?8�>�9��'�`�?�޶?M��?�I>XW�?�s?�~�>��z�C�/��糿�4��+it=�X;���>^,>�P��*�E�<������9�j��)�B_>��%=�^�>ཇ̻��ʶ=2��c���N`�G��>�<n>�H>��>�~ ?}��>��>[=������𖾒�K?=��?���n��<���="_��?�,4?0-d���Ͼ��>Kz\?���?��Z?;��>|���-��ſ�XT����<�K>���>�G�>5o��1$L>n�ԾW>C��>���>aj��$$ھ���8���I�>�Z!?H��>�¯=�� ?Ȝ#?z�j>�(�>�aE�:����E�ڱ�>D��>I?��~?��?Թ�_Z3�����桿��[� :N>��x?VV?cʕ>Y��������zE��CI�2���X��?�sg?YR�B?;2�?i�??��A?-f> ��bؾ����s�>��?��
���5�����=#�-+
?Ѓ? ��>���}w��(%=��������>mW`?]'?�	���V�r��<}�<vr�,�1�C����,<	�>�>ǟ���=��,>�O>�p�[-��������=B�>�:�=���$��6@,?��%������=��r���C���>��L>j¾���^?JV>�"|�����7��P�T�x�?��?�?���/]h��v<?�<�?�?�w�>	����-ݾ}��{�m�y�?)�JY>r(�>��l��H徍����L���,���a½�Un���>�~?�D?=��>ᬖ>���>��ξ�;��(ƾ�����[���oDH��v���㾡vǾmE�s5�=3*�����5�>�cX<�ё>�U ?@�><�>�V�>�Rt�v�>:=>-�>�8�>��>4e>���pW����̼�eP?�I��W['����#���@?\a?��>q�n�1������} ?�~�?C��?��z>dyh��R)�}}?�]�>��OO?�G5=� &��D�<vr�������~k�*�>�/νI-<��XK�5�b�a�?�%?~S�|Ⱦ����Dþ��=�?�??L.���`�ԕd�:�]���_�ޚ'�q+~�P����B�_�{��䤿͢���zo�%M�
�'���5?�?�@��ݾ"���wd�w1F���P>�?C��>��M>��|>�����#}O��8��þ+��>�6?���>I�/?>�8?P�?�<?eӚ>a�>Jξ��?�xg�M��>��>�R?.�?���>GN-?��?�^4>����K5�������?v� ?��?�?JS?`�`��E��gp����;pp��Oa޼�J^���F�նg�nvN�PԔ=UJ>(?�}!�pZ4�de���>�D?���>ڲ>=��.!��>��>�u?_�f>�R㾳gf�  � ��>ρ�?JA���=�2>kZ�=���<�z<��/=`����s�=�ؓ; �������g@->N��=B�ż6/ռ-��<һ<�|:1u�>�?Ҙ�>�I�>�<���� �2��M�=�Y>�!S>�>:Jپ}��}#��/�g�sdy>7v�?�w�?��f=��=��=#r��_F������`�<v�?B#?�RT?T��?��=?@i#?N�>Z(��K���^�����d�?|,?���>S����ʾ�쨿�}3�B�?X?>.a����#)�O�¾hLս,�>�I/�e#~����\D��F|�N�������?���?HR@�$�6��u辞Ř�.]��՚C?,/�>�k�>��>��)��g�a*��);>��>R?ļ>2O?�u?��X?��C>��;��~���ɖ���޼�+>g�9?��?iӍ?�pt?:��>�>m�2��|����\����mv�%�d=�_>JƓ>X�>��>�L�=mཆ��M4�L[�=�k>��>�f�>���>�	|>���<��C?z?�T���[	����L[[��B=��?Tݲ?�aS?yy���W���?���
�O^?i�?u�?)Q�>t@f�_`=��`�I[t����d>��>�|�>�Қ����=���=�
?Cf�>�����þ?C���v�Ob�>[#%?�W�>��ƿ+�v�3
��;����\����^_�fj�����Z�=�{��f��wO���?\�?������n����z�|��}3�>[��=�96>߼�=����po��ґ;64>=�[=ʓ<�[K�`	@=�:���7�<��\�$��<Р2=Em�ϸ����žP�{?K�J?2,?��B?�z>}�>S`��u�>ȱ��E�?EO>�xf�{Y��VW;�G��I㕾�#׾�Ӿ{sa��١���
>�%2�5�>0�;>t!�=ѣ�<U;�=�`^=�ޑ=���&=���=�<�=٥=��=�D>c�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�lc>o�t>4�L�b���ž$��~Ѿ?\�V�2�����=ƈ�>���iMԾ�9=���<Ǻ/=�����x��}�=K1���>qj�=Ϭ>�_>��>�O�O�<��<����=!�{>���=RV�<LM;��M�=�Xϼ�x>I�a>	+�>h�?��-?(�d?���>7dS����]v�����>�>ex�>$+��x>v��>�8?�EE?�K9?���>��=�$�>���>/�-�=�w�m���<��VN5=s��?q-�?�Z�>�p�:(�V�<v�%U4�k���??�4?˟?�Օ>�U�o���Z&�Z�.�����V�\��
+=xr��uU����f�]���=o�>���>]�>�[y>^�9>b�N>��>Ӫ>f��<Xy�=���ǚ�<���ﳄ=�f�����<Onż�~���'���+��z���Q�;�`�;�\<	^�;H��=CK�>Q�>���>6'�=���0H2>����FJ�^��=
(���_B���d���}�8).�b�1��G>tYS> �r�灑�Lk?�a>�M>��?Wt?��">�7���ھC᝿�^���N��ӿ=��>c�=�v�:��}a�r�L��ѾB��>8ݎ>U��>��l>,�@"?��vw=��ᾷa5�"��>&���2���)�=,q��6��A����i�toܺL�D?�C���H�=�~?W�I?g�?)��>�瘽�|ؾ�T0>/Q��c�=`�(Aq�BA����?)'?3��>�쾄�D�)B̾�¾�0ѷ>�I��P��ŕ��0�<��|ɷ���>5����о;3��b�����A�B�br��ݺ>m�O?��?2&b�~X���LO�o��pE��Bh?�g?o�>�L?>?�ˡ��v�"l��W�=/�n?x��?/.�?��
>��P>y����>E�3?��~?O]�?�Jq?������>��0>q�>��=�A4�:�0ǉ>�>*��=�Ps>��@?��R�����שξ&�ؾL�j@i��1>=N�>��n>[�>�큽y���̚=�\>��M>7�}>QD7>��>mɢ>���4����?�o>ڢ>��2?X�x>���=H���?����@���+�1�.��ڕ�����o:5<\B��[��<<��;�$�>�!Ŀ?a�?� G>wu����?�Y�k@J��{X>�C�>(D�����>�O>�L>gΙ>���>���=<�>�Z>�QӾaI>1���\!��&C�,{R�G�Ѿ*�z>d���H&����6��� I�KO���`�2j�o(���/=��ȼ<>�?� ��	�k���)�IA����?fb�>+6?�Ɍ�3��k�>���>��>�@��㊕�Uč�[᾽�?Z��?�Wl>���>��O?�?����8���S�ާw��=��}_��a�,�����}��S�r�����X?�t}?�J?��=��w>?����ˍ�Z�>`+�9�A��=���>�!���n�NLھ_�¾b����?>�Bk?���?O�?��\���X�nU'>�:?�E.?�s?5�0?��9?�&���%?��*>�?��
?_�2?"j-?�[?=�;>�=��Ż�X!=攽�č��Ƚ5s��?غ��d=`=�=��պ��@<HY=>�<�E���ټJ�Z��k���̱<#P=_�=���=(Y�>�G?��>�x�>��?h}������D?��'?�M�=�[������ï�0�վ���=ML?S�?�H?+�>�1B��@�8��>�B�>��>�y�>�D�>Ϫ�����I�<:��>�31>�">��Ƚ������l�����*>���>�=�>�bJ��h2>᰾k�6�8�v>A�@�xr_�ey�h 9�4:�&G��M\�>6.<?��?9�.>�5�e�/�4�[��a?
�I?��h?C?�e#>˧�&\S�B�h�ȧG�<�>ӯ�==��]V�����֖?�+�7�	�1>��z��Cc�=�>����iv�
\����{��Y㾭0��C�G��Z~>2����k��홽��">Ih}=.��Z��������c��"�G?3I_<�����p�:���ϑu>F̻>&A�>�^_��ј���>��);;@���r�>X>"�ʼV���H2�Z�(�,�D>R=>?g�c?_ф?]���~���k�X���%��w�3�>�D0?G� ?�?��->H��|�W���~��5N�*�?���>'�2�u�.��uɾ�K��]龑��>���>*D{>�7�>Y@K?��?�U?�2?ʁ	?��>
�P�S5뾊�!?�9�?��=ea���_<]�Oc��q�>�o,?��w�>4;?6�>?*?{�?�8�>E�=#�X5���>.Ɏ>��P��姿�w�>� ?o
�>�n?�=�?!�>��e�������W���P�tu�>M�?�-F? ?���>���>㞾���=�:�>,c?�5�?;~p?� �=	�?h�0>�+�>��=Ŝ>ur�>��?�O?�r?�J?��>�o�<�D��7o��:�i�и3��><�)]< is=�Kv��l#�hb�<�'�;�%���U��P��1�W�=}q�F��;M]�>��t>�����/>Sľ�3��E(@>�㠼Q̛�c]���F;��չ=�ր>��?V��>�}#�z��=@��>�
�>[���'?��?�$?1�;&{b��<ھibK�d+�>�B?\0�=-�l�ř���v���m=��m?Ld^?uV�����b?9,^?�/�=�<���¾�b���{TN?c
?�fL�(ӵ>�?,br?�;�>��h��m�+��!�a�p�m�X��=�f�>F��[e�~�>t7?���>Cmd>v��= n۾��x��x��#j?�?v��?:?��/>Oo��߿����(ޑ�{�]?�?�>Jç��5!?�3�0�о�K��b�����ᾦ۫��ޫ�x�����ʷ(�Z>#ݽڕ�=�k?μt?V!s?a�`?F&�3�e�a��"��x-X�C������C��JC�4$C�f"p�n��	��������(=kZ����K�T��?�"?��A���?;����P��m����j<�S��%nL�3s�=m髼��=C5>ja���a�3p�� *?�j�>�S�>ψ/?p�_�ӔE��|C�G�P�����L�/>�J�>�g�>��>F�>�x�h���|+ƾ�T�A�C���t>�h\?�,C?�~i?��� 4��<|�<�s������J�4>%'>w��>Dy�;���U&��9�9�u����I��6��)f�=30?���>��>�Ց?Բ?"�۾u ��
Ja��$<��	4=�ƴ>E2j?���>�qQ>ރټ��
�-��>>�l?���>Z�>锌�<Y!�F�{���ʽ�$�> ߭>
��>��o>�,�L#\�Xj��c����9�r�=*�h?*���J�`���>�R?P�:<H<
�><�v�V�!�$��J�'���>}?0��=��;>уžx$�
�{�29��i�)?�M?�����	.�TC�>��?���>G�>T�?���>`�ľ�	<�:
?U?/?H?g�A?�"�> �k=J���֬˽�+1�p�3=�3�>X�W>��x=%M�=)�_gU�1����<��=��6�ֲ ��=�@��F�Ϻ�%D=?�B>��ڿ#VJ��_Ӿ{�Bz�3�
��{���9ǽ̄�{�J���XE��.�x������V�5�_�Ěd�sa��s�i�a�?���? ��fy�����|���O��Oi�>�υ��Kj��v���F��8̏����HԷ�%��P�Gn�Ddg�G�'?�����ǿ򰡿�:ܾ2! ?�A ?4�y?��2�"���8�� >C�<4-����뾫����ο;�����^?���>��/��q��>饂>�X>�Hq>����螾"1�<��?0�-?��>��r�0�ɿa����¤<���?/�@��A?FQ(����a=V�>o�	?3F>��2�G���������>I��?\�?g�l=��V�����ce?Jb1< �D�יͻ�H�=6A�=|=E=��'L>V��>�%�O�B�����	3>��>�&������[����<��_>|�սyᠽ6Մ?{\��f���/��T��%U>��T?"+�>�:�=��,?M7H�Z}Ͽ�\��*a?�0�?���?!�(?ۿ�
ٚ>��ܾ|�M?YD6?���>�d&��t�ԅ�=�7�r���o���&V����=]��>�>��,�֋��O��I�����=�����ǿ�H/���0������g�㏽�*@�6~B���7= ﴾�ט�y�S�@��<I��=��>�Kg>$U^>} p>�4F?�Y?8�>L@�=v�ܽ�ׅ���Ѿ���:5d���ڽ��&��Š�ޝ���R��z־�L��+8�$�<���[L=��h�=x@R�d���b� �)�b�%�F��.?��$>�pʾ��M���$< �ʾ�Ǫ�{!��;B�� ̾�x1�z�m����?b�A?b�f�V�!������Y�W?M,�.��������=�)��A�=���>�ԡ=�X�23��^S��,1?�o.?�ŉ�3����?�޼��=C8?��'?����lV�<�F?�&��I���5�>`��>�J�>���>���>����w�[�b?hČ?�h]�k˾֖�>��þ�0����.>���=\�=�P%��wc�=�_�=�����㾽�,���\���HW?�E�>�&*�jP��������A=��x?�?&�>$k?�+B?u�<����.S���	��|{=��W?(Oi?#M>��v�Ͼt���Ǹ5?��e?C�N>]i���龺�.�%Z��E?��n?;�?�4����|�o<��{��Ns6?��v?�r^�vs�������V�n=�>�[�>��>��9��k�>�>?#��G������bY4�,Þ?��@~��?��;< ���=�;?w\�>ȫO��>ƾ�z������Γq=�"�>���`ev����CR,�Z�8?֠�?J��>������Aa�<�e���?��r?�������,~0�`�l�X ���_�GU�>{t�=�=n���dI�$沾�RB� +���8���>��@�z�=���>Qf���꿿Pٿ�֬�~S$�W1��H?u?u�#>: ����m�#����0���\�05��0�>g�>��������{�J�;�ϝ�����>Κ	��g�>TpS�����|B����4<�>�b�>d��>�h��0!��R��?I��}Aο����(��~�X?B`�?�l�?�H?L 0<o`w�Ŧ{��-� &G?��s?yZ?,�#��B]�'�:�%�j?�_��wU`��4�jHE��U>�"3?�B�>M�-�s�|=�>��>^g>�#/�r�Ŀ�ٶ�$���Z��?��?�o���>o��?hs+?�i�8��u[����*���+��<A?�2>���D�!�F0=�JҒ���
?X~0?'{�o.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?kٵ>vڂ?�M�=���>ky�=������f>���=��:��z�>��N?w��>���=���Q/��UC��.T����-�@�f!�>T}c?>�J?�Wt>�����Q�-I�?ӽ�/�0�G�H�2���	W޽��?>#3>�I�=<���ž��?Mp�9�ؿ j��!p'��54?0��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>@�Խ����[�����7>1�B?X��D��t�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?gQo���i�B>��?"������L��f?�
@u@a�^?*C�ҿ��ݾ�P�����;�\=I�$>N烾 8�={�>|����;ཻ�L>�y%>���>���>�$�>=04>-���/<�Q��X-��OЀ�%�0��+�j���mվ���<:�������o9N����¯g�K϶�jc�����f�=`�>?�J?i~m?���>���l��=K,��@���7ٽ�e=�e>�0?�t"?{�*?�_<�r��C�_�{T����о���i�>Ī�>�@?}� ?�l�>�ڱ=X��>���=���>ϕ��F;=W�S='0�<e�b>N�m>�J?$^�>�C<>��><ϴ��1��u�h�^w��̽�?ၝ�7�J��1��v9������i�=0b.?�{>���?пp����2H?���n)�!�+���>y�0?�cW?�>+��,�T�2:>X��ަj��_>�+ ��l���)��%Q>el?��g>�ev>92���4���P�U\���0u>>r3?e�¾=;2��Vs�6�D��پ��C>�2�>u︼[������ڍ��n%k���v=��:?�?c���e����s����2�W>��Y>�i&==�=}XM>�ȃ� ��r�A��9=[>N�i>�B?]->t��=1�>u˙��R�v��>\oB>�?%>�??|&$?�Rb��MB����,���u>���>�|>n�>��K��(�=��>|�d>M���t�
�	��?� X>��!�]��X��I��=pf����=a�=�K�(28�Y�*=Kz?>\��j����"��ؓ�=�\?��3?�H���=��־iz��+�� �?�(@�ۅ?k�*���CgD?#!�?Bż-�=D�>`)�>�7�͙u�2�?A����=��D��� w��ޫ?�?�?��)�dh����4�V��>���>)��Ph�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?[:Q>1ѐ?չo?'��>�2(��*�47��m䎿��=1 n�̲�>!�1>ؑ����9�.���@���s��3�|�1>]EO=/��>�t��^ʾ��>k���섨��`����>e6T>
t>V5�>\�?���>�&�>n�=yD�����������I?�J�?fC�x�o�μ^=ȍ�==�q��-?3�4?"LX�ǡѾ��>f�_?R�?U�U?L��>e
������t��5��q�,<e<>x�>3��>������`>��Ǿm7�cg�>	C�>����W�G����u�<.��>�#?���>�s�=˙ ?��#?�j>�(�>aE��9����E�ɱ�>J��>wH?}�~?�?�ӹ�?Z3�����桿�[�T;N>E�x?V?,˕>S���烝�YE�vDI����2��?�tg?T��?2�?�??H�A?)f>��Lؾ�����>��!?����A��c&����Jy?�R?�G�>�b=ս��ּ���=���5�?x\?��&?c�0�`�ST¾��</�(��LI�Jy	<y�;��5>Og>t����=8�>�گ=d5l�,�5��*U<g��=cb�>��=�6�(5��A,?i2>�{����=}Wr��KD�! �>o�L>���4�^?�e=�֟{��� r��b�T�e�?���?�D�?Gk���h���<? A�?�V?yE�>Ѯ���ݾK6�Cx�]y��X�Bi>n��>tU��������1^��z9��F�Ƚ�����>�t�>�L%?���>��X>翮>� >��'��*־~�پ�X�>%��+����������-R�M���ξ*������>doR�n�>w0?9�m>m#�>�1�>U��b�>���=]k
>'��>��=�>�z�<�J�=��%�_nW?E�¾��$��L���g���[?ީ�?ZX�>I!\�`.�
�$���?{�?k��?%#�>6j��޾��?b�?�W�K�?�==n"�ʇ�j�\$Ҽ}��<�Mؽ-E=y?��,���*R�ec��M�
?��?�X�=���������'��Rc�=D�?C�.?�*��\��v�k�c��PW�<o���U#�i���Ƈ���i��C��3���L샿J�4��@�<��1?�n�?����yӾʎ���Ut��#C�B�N>��>&;�>��>sA�>Q�꾻F*�OT��� �P�~���>nf?`E�>�[??��V?��Z?8J?:o�>���>��@�>� �?�M>n��>=N ?�?��?��?m� ?EF7>	����"��H̾!�+?��'?��>�B?��?���"��<��0<��t��,�= pi>Xeؽb����ݽ̺�q=�?���M�8�n����$m>�8?���>��>�����@�����<f��>?yƖ>g����r��u	����>l�?� ���	=��*>2��=������':���=����a4�=h�ȼ��6�f1w<mo�=}�=y�"�,VS;��;��;0�K<+u�>3�?V��>8D�>�?���� ���xg�=%Y>ES>>�Eپ�}���$��&�g�_y>�w�?�z�? �f=e�=˕�=�{��QT�����p���!��<@�?�I#?�WT?(��?'�=?�j#?3�>X+��M���^�����,�?l,?��>����ʾ@�^�3�v�?0W?�Da�y���8)���¾u�Խݞ>JX/�2/~����pD�j\�����P}��6��?���?)�@���6��t�C����P��N�C?�!�>UL�>�>�)���g����;>��>�R?~�>�T?��r?��M?tj>��1��ˮ�cS�����Ѻ�=�E?M��?�{�?FWx?@ԩ>Wy	>&�H�x�~���!����ʇ�U-$�ey>q��>K��>��>�.>��Ͻ��>��>��
�=	�p>���>r4�>��>��L>(k=M�^?x~*?|3�kC�-�-<�M�Pn�� �?���?�f-?�S>[.�n2y��*�F�M?��?1��?�+?�S%��T�=u~o���Ծ������>�a�>;J�>!w�=��=�u=\�@>i��=����:оBA-��u=,��>_�;?YV>�ҿ�𖿻�'�T��U	��{��+���YN�����>�ھ�ҧ�+��q���_�
��ˁ�Y2�q~��%��<���>���=oz�=	<>��\>��<��=n��=���<�h�v�ܽ ����>�qf>o�R�Q�.�����	=Z
>h�ʾ�}?±I?g�+?˭C?�Q{>Û>�32��ѕ>gނ�0�?
qT>�O����7�<��ਾT���5=ؾO#׾d����ʴ>ĦJ��A>��5>PJ�=���<���=��q=@֍=�3��a�=q
�=��=���=�J�= y>T�>�6w?R�������4Q�XZ罤�:?�8�>�{�=y�ƾo@?|�>>�2������}b��-?���?�T�?@�?!ti��d�>N���㎽�q�=,����=2>v��=�2�M��>��J>���K��2���4�?��@��??�ዿˢϿAa/>��S>�%>L�D�������bt˾�l��F�>k$��Ɗ�RW1>�G>����Zֶ��x]�̾{�� �=)⾙N����E=(�ۼ�=(�ʼ�U�>Y.i>��<bG��P=�=b�>b��=�Y%�����$�;���<�W(=/K�>�k�>���>��?�P5?H�U?�@�>�i���\Ҿ����͖>����O�>���>�V>��>�6?��?O{P?�Ț>{o�<�>���>|G�ꀿ��	�]Ƞ�g��H'�?)L�?#�	?�^>=U߇����Úl�\w���G?!A?�h�>3w?*��Z�ۿ��9�+�9�Jz�����m�9=���ic�<�<"�4�!5����<��>�F�>q�X>���=̒>>�v�>��>�D>U>�=M��=��=m!��̜:.>�䲻}o�=Q�;=,�=4�X=yè�um>*�W=��=u�O�l���EL�=��>�>c��><�=����p0>:��^L�V��=3��_�A�}�c��~���.��55��PC>1mW>r���W��Y?�\>�A>g�?�ou?׹!>-����վ�6��M�d�*�S�B�=��
>�P?���;���_���M�P�Ҿ���>W�>�ݢ>{m>e,�5?�~t=:^��*6����>qB��:�����.q��Ť��ß�J�h�͇��xC? 3����=�6~?Q�I?1ʏ?�A�>ǻ����־܄4>n<��yn=ó�4Ro�ե��`4?t'?I��>��龇�C��H̾����޷>W@I�(�O���S�0�4��;ͷ�0��>������оZ$3��g�������B�Mr�+��>�O?��?�:b��W��FUO�����'���q?�|g?:�>�J?�@?�%��z�or��w�=�n?���?L=�?q>d�A>��׽�o1?1w?�u�?�|�?9�?s#���&�>�#S�?|�<z삾��<R>8���=��U?0I?F?�P��}��z	��O��5�e��=���M��>@��>�IR>QI�=��<-��<}&�>*��>�r�>*YM>q�>�\�>������"�G$?7�N>��>8�??�
[>��>Hɝ�B���w�=����Z�2��Č���O�=0�<�ܘ�<�C��ӏ�>꙾��x?��L=!��:?[Ӿ1�=�w�>�(0��XN=�=�>=�=a)�>L��>�$?\�=�a�>ږ<>�DӾ�}>m���a!��,C���R��Ѿ�yz>����;&���o���>I��n���f�`j�-��4>=��M�<pF�?������k�&�)�<�����?+Y�>�6?�׌�O��Բ>���>ō>;M��Î���ƍ�h���?��?�;c>��>I�W?�?֒1�03�vZ�*�u�m(A�,e�U�`��፿�����
����-�_?�x?1yA?�R�<+:z>Q��?��%�[ӏ��)�>�/�&';��?<=u+�>*��-�`���Ӿ��þ�7��HF>��o?;%�?wY??TV�r0��"+>ϪA?�6?e�r?�5?�]A?�?�,?^?*>e� ?�?"31?�Q,?I4?)�">�=��m�"6*='y���M���aӽ�Dѽ2�ּ��=�Ē=|?<�����0=�3<0�G��L&����<\���Y�ú�=䡵=!N�=���>z�\?$��>�a�>��:?�4��<)�by��kf1?i�L=)B��侌�����%���0>u:p?��?)�V?}�~>b]D�պJ��>>w��>B�>	4s>t7�>os��}Z���;=+�=l>�=�?+�툉�V�����j�<�}>;)�>�I}>h|���2+>�]���y�d*f>��N��K��4}R��]G�1�A�v����>_K?B?�|�=���cƑ�#�e�:F(?'�=?8N?�~?x�=��ؾT�:�RK�Q����>RX�<��F����4���<�M
;�8p>����<v��Z[>���=��q�ݩK���Ҿ�ڀ=�
��1�=(���Ͼ(�}� J�=�>����F�v���1=����F?�7{=P���m�Q�i1��?�
>3?�>5��>~c��Џ�:����]�=e��>��R>��-}�2E�����Cv>�/?M�p?�?h�A��JU�?\�O���j���T�8�0?s�>`�6?��>5T�����'O*��Pu��NH����>ѵ?N�;�&P�B(��
�a�߾�5l>�?�j�>k*�>�K?�Ǿ>F?�'?�?�L�>S.2=B��PJ&?l
�?3�=� ��WIO��47�bE�	{�>� '?�H�0> �?�:?�`'?�N?>�?�u
>���Y�@�dʔ>Ov�>�,W�_����e>QH?��>'X?���?�5D>��2��l����Ľ�b�=�b>�n1?K�"?�?1r�>b&?��[�/��=���>��i?Ӆo?��;?Tb�>�1?i�¼ {�>5&��}S�=w܇=��?�O?6Qg?D.T?��?��a=�(��ת���%Ƚփ�=�qe=�_��=>0v>�S�;֏=*�e=#�F��/��C�d=bF��d *����=�j�>�t>�񕾓1>s�ľe=��Z�@>����,��.�3�:��/�=2��>#�?���>�#��0�=俼>9�>����+(?�?`?�L);̆b���ھ�LK�8�>�B?��=�l�Q���4�u�2�f=h�m?M�^?��V�����L�b?��]?/h��=� �þz�b����^�O?5�
?<�G���>��~?h�q?^��>�e�$:n�'���Cb��j�2Ѷ=ar�>OX�K�d��?�>i�7?�N�>�b>*%�=Zu۾�w��q��\?��?�?���?	+*>y�n�S4࿁ ��&9����X?}��>l���R?�ݲ�#�վ���i2��~eܾ�m��󟪾�F��C詾�):�}���+�����=nE?�u?yNv?9d?����U'g�fea�{�~���W�������eRH��C�EPA���u�FA�Ȳ��$'���N=��`�j>�;B�?H�$?�4(��?���Mf����&��<�!"��	�ļ5>�Eм�Lٽ".K�d`��%]��ܙ�Qv?�L�>�<�>Y�B?��M�%A���K�k�=���߾�2>D8�>{�><��>t��=f-����j̾T����&'�q}o>�Ib?�DL?mn?1���(�2�N`���U$���~�HX����K>�d�=aϋ>�F�z�$��(�09A���u��x��"���$�O�o=�F3?@�}>&[�>Ö?k�?G=�v
����o��0��D<Ge�>�.k?�2�>���>Н��1"����>l�l?o��>��>؈���`!���{�Ni˽���>�	�>��>�|o>�s,�w \��o��K����.9�V��=��h?om��ͧ`�1��>�R?��:�<G<��>:�v��!�ܲ�U�'���>�?��=��;>�hž��պ{�fl��p,?ӗ?iM��d�#�s�>í"?\N�>���>EV�?�2�>��������Y?"rO?RYC?�A?B��>�?X=�	H�8з�Q��S�<㿀>R�Z>ݣ�<�5�=�J�O(V�i(�#��=q|�=]k��)���O��0⼻!�<Z�/=7�7>�^ۿ�K�KAھ�^�S!�G�	��:���b��pS�� ���������oy�����Z!��_U��d�`�I�k��H�?��?�򔾥
�������r���$��G�>Xnq���������3��┾/s߾A3����!��}P���h��e�m#'?�A����ǿAˡ��Pܾ� ?� ?jIy? ����"��y8��`">�M�<	���U���p����ο�֚�r�^?��>w���$�>���>9YX>��p>����Þ�_�<��?4+-?�/�>c�q�#Nɿ�y���L�<���?��@
oA?P�(�'f�xzW=%��>Q�	?�?>��0�>��G��O�>�0�?� �? �M=h�W�6i
��Ue?+1<��F��[ٻ��=R,�=i1=�����J>��>k<�2A���۽�	5>o��>�<#��f�b�^�+K�<$�]>IԽ/���4Մ?({\��f���/��T���T>��T?+�>]:�=��,?Z7H�`}Ͽ�\��*a?�0�?���?%�(?<ۿ��ؚ>��ܾ��M?_D6?���>�d&��t�΅�=?6�U���}���&V����=P��>f�>��,�����O�J��?��=<���
˿+I��M�ɐ��� >�G�>k)|�hݴ�F��<�R��=����Ͼ|<h;�>�K�>
ݔ>6�=�V>4�<?�$G?ڇ�>;O+>�E`�i���'��T����H��5��H0>d4�x)_�}vþ���OH�$J�6GJ�Ϣ>���=w�T�������"�4\�3�I�(?�� > �þ
�M���A=��;ݖ��j4�;Ý��
�ξ~�0�yg�ޜ�?�@?zV��7Z��m��c�*7���fT?o��^�'t��M=�=���;�1v=K��>��]=JN��/��&I�]@?�(?�@ξ��T�z��>��輗����C?]Y/?��<.�>���>ML�tx~��>iI�>pe�>��?���>-/����5�!?�&-?� ���o��p0>����ZN����>b�z>$S�=�z��
>�1W���v�S�=+�=
)=�rY?a<�>�����m�b��"��f�<��s?�?��>�.l?�>?3 p��
��L��� ��=#z\?ڕl?U��=`<>��ݿ����gb*?7�n?C�>�g��ﾕ�0���`x?݆p?��?�⪼.��j���� ���8?��v?�r^�qs�������V�]=�>�[�>��>��9��k�>�>?�#��G������mY4�#Þ?��@y��?��;< ���=�;?\\�>�O��>ƾH{������1�q=�"�>ጧ�Qev����2R,�P�8?Ѡ�?���>쓂����^o�=$󘾛�?��?ܩ��(�T=�4"���V��6�i#��;G\>y����=����P�P�)� ��w%�W���Nd<��>��@�*���!
?Qt���޿�̿S勿&b��ZI��gq�>ӱ�>��;��B���I�UMU��40�78S��־��>m�9>�Nf�yK��N�����T���y=���>i��n�>�뙾���GkF��6;���!>.�>N�l>�>�u�˾���?��̾&������� hB��F-?���?d�?�M?É��ؾ8��u��<t?$[K?*d|?UEN>�@���ｏ�j?�_��U`���4�HE�	U>A"3?�A�>T�-�ܱ|=�>1��>9g>�#/�|�Ŀ�ٶ�N���3��?���?�n꾤��>���?�s+?[i�8��[\����*�f�-��<A?K2>���ڸ!��/=��Ӓ�D�
?�}0?[}��.�7�_?�a�+�p�l�-���ƽ~�>�H0��z\�<k�����Re�J�dPy�{�?�Z�?��?����#��5%?��>����IǾN��<�y�>��>�N>/`_���u>��d�:��=	>8��?y�?7n?���������[>�}?90�>?	�?�G�=���>���=�����9+���#>�o�=�=�uh?�fM?��>���=��7��/��3F��{R��t��C��߇>��a?�sL?q�c>O���_n3��3!��ͽ�j1�0A���@�ξ(�4�޽��4>�=>R>fND�h�Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�c��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?�Qo���j�B>��?"������L��f?�
@u@a�^?*2�п8v����;7��ؽL��=��>C��H�
>��7=5\c���@>���<E��>�W�>0Л=|�>�nD>�t�=3���0)��c������.�k���#�]�$�d/��2k��\��<�)�㯾��Ǿ%Ē��<��a���ν������>��S?^xF?��r?��>gB`�Bp�=� � �ø:�,��T�=��>��)?�[U?T*?:��=4����V����<ס�ҫ��7�>�>>G7�>Q��>V��>i1�q�A>f`>�:j>`�=�Z�<��*���=�e>*	�>���>�4�>2��=2�X=q���������c��fD���M=C�?r&��%iA�A~������¾�:�=S8?~l>�Ò���ȿ����C@?��k�����~�4�=0x$?#�J?Z>ٽ��N�z�f�2>��NK�u�8>uZ�������<�2�K>�?X�>p�>b���w�������6����>��c?0B��	�<����w�:��R侍ީ=���>a6�=`Ⱦ$j���ꏿ��V����Fr7?l%?U��=阍�������B�Խ/͐=�
>���=a�V=���=*&�=Eۿ�@{Ž�)޼I=輋�?��2>1d�=��>�M��?R��,�>�	J>0>v�>?��"?� :�瘽 ����+��{y>� �>�ك>��>RdF���={��>wb>�c�C̓�;���7�x�W>�D����Y���p�kK==~s��|8>ĕ=�R��;
=�9$&=�~?���'䈿��e���lD?S+?Y �=�F<��"�E ���H��G�?r�@m�?��	�ߢV�@�?�@�?��J��=}�>׫>�ξ�L��?��Ž4Ǣ�ɔ	�0)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�f�>?y�MX��^����u�:�#=l��>�8H?�X��x�O�� >�w
?�?C^�4���1�ȿ�{v�/��>�?���?	�m��@���@�h�>��?YeY?xpi>�i۾`lZ�Ҏ�>-�@?�R?�>�:��'�E�?�޶?R��?�* >��?��v?���>�wB�_7�p��ƹ��"r�����=A��> <ͼl훾�b!��t��|���
{��-��n>�z�=���>T���3���ך=�E���Q���>�6Q�>�R>�Ak>�>�^�>�H�>��>6�C=�釻 ��r����K?���??��(+n�'M�<���=��^�$?E4? �[���Ͼvר>x�\?f?�[?�d�>���/<��\翿K|�����<n�K>�.�>ZM�>!���yAK>��Ծ�1D�Ak�>�Η>��%?ھ�+��$:���A�>c!?���>��=n� ?0�#?�j>�)�>`E�+:����E�ܭ�>���>�J?��~?a�?�ѹ�=Y3�����桿ɒ[�.+N>�x?�V?Wɕ>��������F�SI�jҒ����?�wg?\U���?2�?��??��A??f>,t���׾r�����>��!?�*�}�A��+&��0��m?�!?O�>�ޏ��ֽ5�ؼ���i��&�?��[?�G&?AR���`�Ml¾Z�<!�!�Cnr����;YA���>��>�t��:�=�>1��=�]m�4,6���l<D��=�=�>8��=��6�Y6���<,?�G��ك���=��r�E}D���>cL>6����^?X}=�o�{����w��'�T����?B��?�f�?�1����h�� =?��?*?9"�>>J���޾\�ྪhw��x�Ds���>���>�k����琤�����MF��H ƽ=��O��>�a�>_�?�3 ?��R>-�>�q��$�'�`!�Vo���]���<�7�M�/�< �쳡��q"�������9A~�i��>�2�>'�
?��c>O{>9��>�-.�ፍ>�&Q>�t�>��>.U>,�1>N+�=�7<
>˽7KR?����ü'�-�辆���t3B?�pd?31�>-(i�����^��9�?���?�r�?E4v>�~h��,+�An?�<�>���@p
?�T:=1	�;@�<�U������6��5�ɩ�>(=׽k :��M��gf��i
?�.?!���̾�:׽�±���=CQo?�?�3�{
Q�t v�M�a�a4K���;w�;����3��Z�g�я����5؋����?�R>�(+?�Z�?6��� �7ߕ�Irx��IK�
<>�I�>H=�>���>�̩=���m| �r�~���/�B�� �>�g?n��> ]H?��'?�(P?�)J?���>wT>�<��>�>�N��5��>d�>��&? �9?�*?Y�?�H?�r�>&�����Yqƾ�^?:��>Q�?:8?/��>����Џ��D��>�g��2�� E۽�2X;2&�=l{�6�@��=��>��?7���M9�B���rx>=�7?pi�>f��>낾:���<s�<���>��	?�b�>����$m�E��H��>�Ђ?�@��ձ=8�!>�<�=c�F��MK�}�=����f4�=v���J�r�a;��=�=q�P���۹h�M;��<�i�<�7 ?��?�/�>���>�������O��r�=�=^>��R>��>�
ؾ�_���l��:g��g{>_�?�<�?׭u=���=,d�=��������܇�.#���P�<�?�v"?�CS?GU�?g=?��#?�}>b�� M���F���5����?A�*?�>����P��	��0�9��?��?�a�b,���(�rpľ#ܽOi>�'�.!}��F���H���{�]뛽��?3@�?eh�$�-�)N�i_��@é�γ??K�>��>�K�>��%�cg�e��3�(>���>��M?YR�>��M?'e??�h?�CN>��)��������3hd���=0�6?L��?@h�?��?Y2�>.W>YJ������W� ݸ���弾�=�ۛ>w�>S��>�y�>��=Z�o��D���]�!��Z�}>-�>p!�>p�>���><��=��G?�H�>JԺ�8��`z����������K:|?��?:C%?����6�og7�]��>�?m�?��?q�>�Յ�=���O�����p����>\�>Ƃ>�8�=�^=]n>�\�>�9�>�S6�¡�-&���e��,?��8?��=��ſ�Mu�����D'��v�::
���1�3�����I�Z���=ڠ��!��ί�fM�dޏ��X�����u���n�YY�>�b�=�J�=p�=�Y�<�M���<�U8=U��<΄�<�kp�[�;ѱ���;	!E�'m$�,�^���==�J�;
�˾Ϗ}?�:I?v�+?��C?��y>D9>��3����>銂��@? V>h�P�ވ����;�ê��X����ؾdv׾/�c��ɟ��G>U_I���>/73>�F�=�J�<��=�s=]Ŏ=�KR��=$�=�M�=*h�=���=d�>�U>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�7>�1>x�R��u1��]��b��ZY�e�!?A�:�d̾k��>{��=��޾@�ƾO�/=��6>Jc=��!\��=��y���:=�k=Rĉ>8^C>�n�=�#��е=�tH=Q��=�O>����\5�X)�0=2��=�fb>Z�%>���>�c?,Q"?Ұ]?Y�>�<�W�Ⱦ_ް��щ>�3��>�#>�w�>:|�>E6?w�A?F�@?�ȵ>�P�=�դ>e��>���EZ��¸��3���2>���?E~�?���>��7���g��x
��M��'T�I��>�M@?��?�b�>d
���念oZ�0�u��l^����=K�>���̯���L>Z�:�����A�A>���>��>�5�>��>��>�<�>4y>2ۼQ�M=���=P�?>l�>9��<D սR�r=kD��h����.���<utd>����yu����<
�=���>]>˸�>��=jI���H/>���,�L�F	�=�V���)B�Y+d�^3~�d�.�~s6�ŰB>�W>�����.��C�?SZ>&�?>0��?�Gu?�>�x�c�վ�H����d�yS��J�=��>`=��r;��Z`���M�JyҾ]$�>�K�>�r�>͚b>�X��J��`ͽ �H��?U;�n�>�<1���4���I���0Ј�����Q�Y?.�\���i>ٌ?��[?��t?Y��>\���!Ͼ��\�;훽��=�??�!8����>�X?��?��>�7�Qr� #���u���>6^!�<FN�ʤ���(��!���Ǿ\t�>�,��4�aU"�N��7Њ��D��5��Ț�>3~=?'Y�?R�J���~��wZ�ؘ4��ǽpj?�I�?/��>��>[%�>�����zʾUX���վ< W�?�B�?R�?o��=e��=������>�?���?�0�?i n?B�'����>ȴ��� >�#���u�=/�=,A�=Q�=�z?X�?�E?�̍�5%�\�����uM�=��=�_�>�j�>�\>�Z�=y�j=B�=�YE>��>��>�aY>�8�>¥�>eؙ��
���3?��	>���>��=?Oe�>���=��+�%�׽P5=/���s�BA����s�W|�n���1f=]~�;��>Dm¿��?(�X>���0�?Ag�� ���)>N��=@������> \l>lX�>�k�>��t> ��=2r�>��D> fǾ���=�Z��W�|$�{�"��!��P��>r~����p�DZ޾����B��������w�Bc��@{�	l0�CE¼}I�?ł�B�W����~hԽ�<;?*t�>M<2? �þ�u����l>�n?�ֳ>a�ƾA>��S������ꊊ?���?�=c>��>��W?,�?؍1�3��tZ���u�x&A��e�z�`�፿����
����"�_?��x?ryA?f�<�9z>���?��%�Cӏ��*�>�/��&;��I<=�-�>�)���`�O�Ӿ'�þ\;��FF>�o?�$�?XX?RV�FI���H>;U0?�1?�.q?�4?�9)?��T�ɟ?���=���>�'?�_2?��9?�8?�7h>[�=S��;��<SC��i���R�������{�9��<�=�/=��4=�mB��o��;����q=Ft����P�B<�<�=�n�=��)>l��>4�U?��>�i>5�J?��%��<�A���G?�I�=� �O�T�Y���F��?Ǟ=X�a?;��?;�e?G�>��,�J���{>�">ܢ�=PǨ>2��>��+���W��#>A��>��=3��<jm�w����X��镾�F >��l> �>�ց>o�9��%>>d`�������a>�k1��~ľ]�<�2F���1��%v��I�>�7P?�+?���=�n �g5
�c�d�cr"?<??��I?ss�?w��=�Rܾ��?�
C�������>��-����Nl��w ���4��mü1��>�j���/���Q�>�!���V������^��"'�O)��r��Ǎ=��F��)��#5콄��<3E#�J�1�3��K녿����&Ld?�f	>���h����ľH�=g�=��>�h]<��>��/�jʟ��۽=�
�>�T?C��>T"׾��O�����Ɗ>hP=?7RV?�2V?����xP���<�3�ԾX�����k&�>Nj�>G'>:'�>�z>6�4� ]*���v�Cm,�o��>O%?eԾi�=��Ϭ����E?O�d��> �?s������>�CC??��>@G:?DX2?U�>o@�>`�����$? _�?L�">	�0��D!��-?�?_[��l�>�� ?֣T�0X<d"�>�b�>���>�M?�u8?Y�<�(!�}�<�O�>2ؘ>I�5�އ��G�0��>�-�>?-$?E��?z&�>�!A�wf��>3�R���%�P?�?Ģ?���>μ�>Ώ��QY>�*T>�y?/ۉ?��>?���=�)�>��f>+T�>m��|��=l��>�!�>��?�6y?�[?��?�������kt]>�� =V��-3��	�e�a>*��<]C��C���:�<  C���;���:X=� ,�;"'A�bɻ����>��^>6'��s�5>'��'/����c>�w��	���7�_���L�_��=o}~>�4?��>��2�>3\�>��>&��	*?�?�J?�a�?e�&Y��@R�{�>��!?�<6Kq�{����\`�n3(=�s^?�Of?V���l�2�b?u�]?�e�=���þL�b�+����O?�
?��G���>��~?�q?���>��e�E8n�����Eb���j���=�s�>�T��d��9�>O�7?�N�>;�b>��=�z۾j�w�de��?��?1�?m��?6*>��n��1�V�����)P?�P�>�d���$?����B�����?��NȾ|�������
G���|��2(�'��qS���>F5?��q?�8r?N?;n�~�d��`f�і�,U��E��	�qoJ�A�4�`�A�gi���	�U�	��H���͋<�>���3��`�?u�-?�=��>�d����
]��(�>�8m�+��~=��@��=�y>�d���6-�P�R���?�	�>��>�1(?��M��hF�֪&���5����A��=��>A�>l��>:U�<ȏ+��1)����*_�� ����>�mX?�� ?r,e?�<�^�J��3����о�fW���ھ!_�<,;�>1@�>���99�8�.��L?��Pm��9'�r򒾓7��Q�=��1?�t�>R=�>ڭ�?#�?�h����
�̎n�G"�������>��a?�h�>�G>i�f��tھ8��>רl?���>8��>�狾 � �{{�Ͻ���>�ҭ>;i�>6�m>8�-�F\��)�����E�8�\��=lh?{S���$a�1X�>@R?$_
;d�D<1T�>d�v�^�!�����"'�p�>^�?�P�=W(<>sOž9��� {�����8'?T�?��|�ǳ'�
�}>U�?���>�7�>a��?_z�>l���,�O�?��R?ZM=?�E?ޮ�>*�/=ݾ���H˽��=���f=�ւ>�=l>�p�=B>���f>����|=���=�6̼�ν�-ż��t����<K�&=�7>Kaۿ<>K��پS����08
����֑��`w����!B�����x�����'��-V�t~c�䐌�3�l��v�?s;�?�q���3��A���ĕ�����x�>W�q�������z��*��l]����V!� �O��/i�|�e��'?���q�ǿ㥡��1ܾ�" ?�O ?��y?p�Ս"�r8�
� >�c�<j���nq�����t�ο��^?r��>��c����>辂>.�X>J/q>!@��_鞾^��<��?u�-?F��>��r��ɿ7���c�<���?5�@)@?�%����~=���>E�?�d>_M�(��k�����>u��?�%�?�Q=-~J��K2��d?5|_=H\7��b�hI>)��=�j!==����=0�t>���V�Z���&��?�=�0e>��v����tzd�@�FL�>k����&Մ?�z\�2f�p�/��T���T>|�T?�+�>�>�=ò,?H7H�U}Ͽԯ\�D*a?�0�?٦�?��(?0ۿ��ؚ>A�ܾM�M?�C6?���>�d&���t����=�4ἀE��$��f&V�c��=S��>>�>�,�֋���O��F�����=a���տV����]�֏i<u�%��6�=t:�t�侊���]�=��	����>�t7?���UX�L�?yX?��G�_�A?~<X?'�=��>|��<PR�3Ӿ�ѯ��K�"�t=qݽu�j�zξm{����������V����-�t���]��B�D�۳��zh��B��,� �"?� ����-�%YT>*9�=�8Q�au��ߦH��!��U
��֟|�Mʎ?nJ?T����h/���8�`^���<>��J?��C�_��/�y���H>�>v�>]d�=*���L�<��kn�5U/?~�?�浾�<���&>���$i"=�%?j�?�Ƅ<���>�K!?f2�g���BW>�vH>丟>�Y�>�,>�Ī�� �?�P?�e��ᐾ�>Nž��{���*=@>'R2�
���|rY>CF��≾%1�9E�\����<�N?�n>��'�-�Oꅾ�1E=�{b>��W?�	?���>�a�?�g=?9ʼ��
�Ph%��������pG?�J�?l[�=������ξW%��{jB?4f?��
>�U˾l��$ ���̾A?�^j?я?�x��*���2���羈F8?��v?�r^�ns��|����V�=�>E\�>��>��9�&l�>Ǒ>?~#�tG������Y4��?x�@���?[�;<<�ǝ�=�;?&\�>&�O��?ƾ�~��������q=_!�>̍���ev�����P,��8?���?;��>󒂾���]>�T��lI�?��|?�P��'Q<Op!�3>�i�����<�v>\��(�L��㾱9 �[��w�0�����ij:=~>�@|ڈ��k�>+���<ܿd+ſ(���;������>[�>��#�+�3��I;�r�T���/�i�e�ERҾ���>j= > ���r�z�ab~��A<�X�ϼ�s�>����͒>�dv�)���ڏ���=��$ۏ>(5�>�,e>~B併ٻ�p��?��c�ʿX���k
�I�P?FD�?�s�?�`?qi�;�:��vL����<?�|?�a?q�Y��&]�JR�{�j?0_���U`��4��?E��U>�$3?�6�>9�-�\}=S>���>�j>	/�-�ĿY׶��������?+��?j꾴��>��?ho+?h��8��j��#�*�W�C�~/A?	�1>H���^�!��'=�;Ӓ�m�
?�0?�R�n1�\�_?)�a�K�p���-���ƽ�ۡ>��0��e\��M�����Xe����@y����?M^�?h�?۵�� #�h6%?�>c����8Ǿ>�<���>�(�>*N>ZH_���u>����:�i	>���?�~�?Sj?���������U>�}?@�>���?�?�=;s�>���=R�������#>�B�=�wJ�?�eO?���>���=%o5���.�W�E�!�R��P	�$B�*>Za?sK?p�e>I���
�%��x�ҐĽ��6�������:���0��ϽK>9>A�9>�>w�@��4Ͼ�W�>T#;�� �k��FKٽ�;?ͽ�>�'�>�5#�Ud��l�=�sP?���>p�ǝ��<���9Ɯ�f�?���?��?̲��X�=�>�"�>m19>�ؽS� ��G��LT�=��-?V��������8���0>Rg�?6X�?���?4=Q��	?���P��`a~���[7����=��7?�0���z>��> �=�nv�ӻ��`�s�y��>�B�?�{�?���>�l?w�o��B�i�1=�L�>��k?�s?\Wo����B>��?�����-L��f?�
@vu@E�^?"��п�l��g���=�v�F�cp.>�M�=C�;=�F�;�T!�p}�=�E�=��)>�4�>�$n=X)A>O�Q>�z>/>S���p)�i����H��������;����:��^0�΋�'��]Q���6;�W*����K����������=:?���>�->?8q/?�Fe?+��>����D�,=�^��3G��N(��%|�!��>�?�B?�6%?�h%�cV��` _��Ro��Ҭ��zξ��>��6>��	?B??0��>�ҷ��*�>ߖ>]�>}�:'��F��<���3Si>���>c@�>)?2T<>|�>�Ŵ���Q�h��w�U�ͽ5�?�����J�$/��ʌ�	����̞=R.?�>����8пz���/H?����"�:�+��>��0?�iW?�>9Y��SNW��>;@�ݘj��>�@��llk��V)���P>�O?��g>dw>?3��X7���P��/���u>C�5?���9�8�'Su��}F�59۾�J>�C�>��W�A�Tݖ�6=�=�g�Z2y=K>:?��?.���v��R�r�'���@S>��Y>�=���=�
N>��X��jŽ��E�� =+G�=|�_>��>X	>���= O�>�:��a=��=��>hJ�%9>��?P�?�?�ǖ6��u���ȼb��>�H�>��>�7�>���!�V>� ?��L>���$߽�ʄ��^��n9<�5���]��:��R�E<�D
��Z�=֮���w��\/�$Ro��~?���(䈿��
e���lD?T+?U �=7�F<��"�D ���H��F�?q�@m�?��	�ޢV�A�?�@�?��O��=}�>׫>�ξ�L��?��Ž8Ǣ�ʔ	�6)#�iS�?��?��/�Zʋ�=l��6>�^%? �Ӿ�c�>��Z�������u���#=���>�7H?�W��E�O��>��v
?�?9[�򩤿u�ȿ�zv����>Y�?q��?5�m��A��|@�ރ�>ޢ�?�gY?fmi>�g۾baZ�ي�>��@?R?8�>�9��'�`�?�޶?M��?�I>XW�?�s?�~�>��z�C�/��糿�4��+it=�X;���>^,>�P��*�E�<������9�j��)�B_>��%=�^�>ཇ̻��ʶ=2��c���N`�G��>�<n>�H>��>�~ ?}��>��>[=������𖾒�K?=��?���n��<���="_��?�,4?0-d���Ͼ��>Kz\?���?��Z?;��>|���-��ſ�XT����<�K>���>�G�>5o��1$L>n�ԾW>C��>���>aj��$$ھ���8���I�>�Z!?H��>�¯=�� ?Ȝ#?z�j>�(�>�aE�:����E�ڱ�>D��>I?��~?��?Թ�_Z3�����桿��[� :N>��x?VV?cʕ>Y��������zE��CI�2���X��?�sg?YR�B?;2�?i�??��A?-f> ��bؾ����s�>��?��
���5�����=#�-+
?Ѓ? ��>���}w��(%=��������>mW`?]'?�	���V�r��<}�<vr�,�1�C����,<	�>�>ǟ���=��,>�O>�p�[-��������=B�>�:�=���$��6@,?��%������=��r���C���>��L>j¾���^?JV>�"|�����7��P�T�x�?��?�?���/]h��v<?�<�?�?�w�>	����-ݾ}��{�m�y�?)�JY>r(�>��l��H徍����L���,���a½�Un���>�~?�D?=��>ᬖ>���>��ξ�;��(ƾ�����[���oDH��v���㾡vǾmE�s5�=3*�����5�>�cX<�ё>�U ?@�><�>�V�>�Rt�v�>:=>-�>�8�>��>4e>���pW����̼�eP?�I��W['����#���@?\a?��>q�n�1������} ?�~�?C��?��z>dyh��R)�}}?�]�>��OO?�G5=� &��D�<vr�������~k�*�>�/νI-<��XK�5�b�a�?�%?~S�|Ⱦ����Dþ��=�?�??L.���`�ԕd�:�]���_�ޚ'�q+~�P����B�_�{��䤿͢���zo�%M�
�'���5?�?�@��ݾ"���wd�w1F���P>�?C��>��M>��|>�����#}O��8��þ+��>�6?���>I�/?>�8?P�?�<?eӚ>a�>Jξ��?�xg�M��>��>�R?.�?���>GN-?��?�^4>����K5�������?v� ?��?�?JS?`�`��E��gp����;pp��Oa޼�J^���F�նg�nvN�PԔ=UJ>(?�}!�pZ4�de���>�D?���>ڲ>=��.!��>��>�u?_�f>�R㾳gf�  � ��>ρ�?JA���=�2>kZ�=���<�z<��/=`����s�=�ؓ; �������g@->N��=B�ż6/ռ-��<һ<�|:1u�>�?Ҙ�>�I�>�<���� �2��M�=�Y>�!S>�>:Jپ}��}#��/�g�sdy>7v�?�w�?��f=��=��=#r��_F������`�<v�?B#?�RT?T��?��=?@i#?N�>Z(��K���^�����d�?|,?���>S����ʾ�쨿�}3�B�?X?>.a����#)�O�¾hLս,�>�I/�e#~����\D��F|�N�������?���?HR@�$�6��u辞Ř�.]��՚C?,/�>�k�>��>��)��g�a*��);>��>R?ļ>2O?�u?��X?��C>��;��~���ɖ���޼�+>g�9?��?iӍ?�pt?:��>�>m�2��|����\����mv�%�d=�_>JƓ>X�>��>�L�=mཆ��M4�L[�=�k>��>�f�>���>�	|>���<��C?z?�T���[	����L[[��B=��?Tݲ?�aS?yy���W���?���
�O^?i�?u�?)Q�>t@f�_`=��`�I[t����d>��>�|�>�Қ����=���=�
?Cf�>�����þ?C���v�Ob�>[#%?�W�>��ƿ+�v�3
��;����\����^_�fj�����Z�=�{��f��wO���?\�?������n����z�|��}3�>[��=�96>߼�=����po��ґ;64>=�[=ʓ<�[K�`	@=�:���7�<��\�$��<Р2=Em�ϸ����žP�{?K�J?2,?��B?�z>}�>S`��u�>ȱ��E�?EO>�xf�{Y��VW;�G��I㕾�#׾�Ӿ{sa��١���
>�%2�5�>0�;>t!�=ѣ�<U;�=�`^=�ޑ=���&=���=�<�=٥=��=�D>c�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�lc>o�t>4�L�b���ž$��~Ѿ?\�V�2�����=ƈ�>���iMԾ�9=���<Ǻ/=�����x��}�=K1���>qj�=Ϭ>�_>��>�O�O�<��<����=!�{>���=RV�<LM;��M�=�Xϼ�x>I�a>	+�>h�?��-?(�d?���>7dS����]v�����>�>ex�>$+��x>v��>�8?�EE?�K9?���>��=�$�>���>/�-�=�w�m���<��VN5=s��?q-�?�Z�>�p�:(�V�<v�%U4�k���??�4?˟?�Օ>�U�o���Z&�Z�.�����V�\��
+=xr��uU����f�]���=o�>���>]�>�[y>^�9>b�N>��>Ӫ>f��<Xy�=���ǚ�<���ﳄ=�f�����<Onż�~���'���+��z���Q�;�`�;�\<	^�;H��=CK�>Q�>���>6'�=���0H2>����FJ�^��=
(���_B���d���}�8).�b�1��G>tYS> �r�灑�Lk?�a>�M>��?Wt?��">�7���ھC᝿�^���N��ӿ=��>c�=�v�:��}a�r�L��ѾB��>8ݎ>U��>��l>,�@"?��vw=��ᾷa5�"��>&���2���)�=,q��6��A����i�toܺL�D?�C���H�=�~?W�I?g�?)��>�瘽�|ؾ�T0>/Q��c�=`�(Aq�BA����?)'?3��>�쾄�D�)B̾�¾�0ѷ>�I��P��ŕ��0�<��|ɷ���>5����о;3��b�����A�B�br��ݺ>m�O?��?2&b�~X���LO�o��pE��Bh?�g?o�>�L?>?�ˡ��v�"l��W�=/�n?x��?/.�?��
>��P>y����>E�3?��~?O]�?�Jq?������>��0>q�>��=�A4�:�0ǉ>�>*��=�Ps>��@?��R�����שξ&�ؾL�j@i��1>=N�>��n>[�>�큽y���̚=�\>��M>7�}>QD7>��>mɢ>���4����?�o>ڢ>��2?X�x>���=H���?����@���+�1�.��ڕ�����o:5<\B��[��<<��;�$�>�!Ŀ?a�?� G>wu����?�Y�k@J��{X>�C�>(D�����>�O>�L>gΙ>���>���=<�>�Z>�QӾaI>1���\!��&C�,{R�G�Ѿ*�z>d���H&����6��� I�KO���`�2j�o(���/=��ȼ<>�?� ��	�k���)�IA����?fb�>+6?�Ɍ�3��k�>���>��>�@��㊕�Uč�[᾽�?Z��?�Wl>���>��O?�?����8���S�ާw��=��}_��a�,�����}��S�r�����X?�t}?�J?��=��w>?����ˍ�Z�>`+�9�A��=���>�!���n�NLھ_�¾b����?>�Bk?���?O�?��\���X�nU'>�:?�E.?�s?5�0?��9?�&���%?��*>�?��
?_�2?"j-?�[?=�;>�=��Ż�X!=攽�č��Ƚ5s��?غ��d=`=�=��պ��@<HY=>�<�E���ټJ�Z��k���̱<#P=_�=���=(Y�>�G?��>�x�>��?h}������D?��'?�M�=�[������ï�0�վ���=ML?S�?�H?+�>�1B��@�8��>�B�>��>�y�>�D�>Ϫ�����I�<:��>�31>�">��Ƚ������l�����*>���>�=�>�bJ��h2>᰾k�6�8�v>A�@�xr_�ey�h 9�4:�&G��M\�>6.<?��?9�.>�5�e�/�4�[��a?
�I?��h?C?�e#>˧�&\S�B�h�ȧG�<�>ӯ�==��]V�����֖?�+�7�	�1>��z��Cc�=�>����iv�
\����{��Y㾭0��C�G��Z~>2����k��홽��">Ih}=.��Z��������c��"�G?3I_<�����p�:���ϑu>F̻>&A�>�^_��ј���>��);;@���r�>X>"�ʼV���H2�Z�(�,�D>R=>?g�c?_ф?]���~���k�X���%��w�3�>�D0?G� ?�?��->H��|�W���~��5N�*�?���>'�2�u�.��uɾ�K��]龑��>���>*D{>�7�>Y@K?��?�U?�2?ʁ	?��>
�P�S5뾊�!?�9�?��=ea���_<]�Oc��q�>�o,?��w�>4;?6�>?*?{�?�8�>E�=#�X5���>.Ɏ>��P��姿�w�>� ?o
�>�n?�=�?!�>��e�������W���P�tu�>M�?�-F? ?���>���>㞾���=�:�>,c?�5�?;~p?� �=	�?h�0>�+�>��=Ŝ>ur�>��?�O?�r?�J?��>�o�<�D��7o��:�i�и3��><�)]< is=�Kv��l#�hb�<�'�;�%���U��P��1�W�=}q�F��;M]�>��t>�����/>Sľ�3��E(@>�㠼Q̛�c]���F;��չ=�ր>��?V��>�}#�z��=@��>�
�>[���'?��?�$?1�;&{b��<ھibK�d+�>�B?\0�=-�l�ř���v���m=��m?Ld^?uV�����b?9,^?�/�=�<���¾�b���{TN?c
?�fL�(ӵ>�?,br?�;�>��h��m�+��!�a�p�m�X��=�f�>F��[e�~�>t7?���>Cmd>v��= n۾��x��x��#j?�?v��?:?��/>Oo��߿����(ޑ�{�]?�?�>Jç��5!?�3�0�о�K��b�����ᾦ۫��ޫ�x�����ʷ(�Z>#ݽڕ�=�k?μt?V!s?a�`?F&�3�e�a��"��x-X�C������C��JC�4$C�f"p�n��	��������(=kZ����K�T��?�"?��A���?;����P��m����j<�S��%nL�3s�=m髼��=C5>ja���a�3p�� *?�j�>�S�>ψ/?p�_�ӔE��|C�G�P�����L�/>�J�>�g�>��>F�>�x�h���|+ƾ�T�A�C���t>�h\?�,C?�~i?��� 4��<|�<�s������J�4>%'>w��>Dy�;���U&��9�9�u����I��6��)f�=30?���>��>�Ց?Բ?"�۾u ��
Ja��$<��	4=�ƴ>E2j?���>�qQ>ރټ��
�-��>>�l?���>Z�>锌�<Y!�F�{���ʽ�$�> ߭>
��>��o>�,�L#\�Xj��c����9�r�=*�h?*���J�`���>�R?P�:<H<
�><�v�V�!�$��J�'���>}?0��=��;>уžx$�
�{�29��i�)?�M?�����	.�TC�>��?���>G�>T�?���>`�ľ�	<�:
?U?/?H?g�A?�"�> �k=J���֬˽�+1�p�3=�3�>X�W>��x=%M�=)�_gU�1����<��=��6�ֲ ��=�@��F�Ϻ�%D=?�B>��ڿ#VJ��_Ӿ{�Bz�3�
��{���9ǽ̄�{�J���XE��.�x������V�5�_�Ěd�sa��s�i�a�?���? ��fy�����|���O��Oi�>�υ��Kj��v���F��8̏����HԷ�%��P�Gn�Ddg�G�'?�����ǿ򰡿�:ܾ2! ?�A ?4�y?��2�"���8�� >C�<4-����뾫����ο;�����^?���>��/��q��>饂>�X>�Hq>����螾"1�<��?0�-?��>��r�0�ɿa����¤<���?/�@��A?FQ(����a=V�>o�	?3F>��2�G���������>I��?\�?g�l=��V�����ce?Jb1< �D�יͻ�H�=6A�=|=E=��'L>V��>�%�O�B�����	3>��>�&������[����<��_>|�սyᠽ6Մ?{\��f���/��T��%U>��T?"+�>�:�=��,?M7H�Z}Ͽ�\��*a?�0�?���?!�(?ۿ�
ٚ>��ܾ|�M?YD6?���>�d&��t�ԅ�=�7�r���o���&V����=]��>�>��,�֋��O��I�����=�����ǿ�H/���0������g�㏽�*@�6~B���7= ﴾�ט�y�S�@��<I��=��>�Kg>$U^>} p>�4F?�Y?8�>L@�=v�ܽ�ׅ���Ѿ���:5d���ڽ��&��Š�ޝ���R��z־�L��+8�$�<���[L=��h�=x@R�d���b� �)�b�%�F��.?��$>�pʾ��M���$< �ʾ�Ǫ�{!��;B�� ̾�x1�z�m����?b�A?b�f�V�!������Y�W?M,�.��������=�)��A�=���>�ԡ=�X�23��^S��,1?�o.?�ŉ�3����?�޼��=C8?��'?����lV�<�F?�&��I���5�>`��>�J�>���>���>����w�[�b?hČ?�h]�k˾֖�>��þ�0����.>���=\�=�P%��wc�=�_�=�����㾽�,���\���HW?�E�>�&*�jP��������A=��x?�?&�>$k?�+B?u�<����.S���	��|{=��W?(Oi?#M>��v�Ͼt���Ǹ5?��e?C�N>]i���龺�.�%Z��E?��n?;�?�4����|�o<��{��Ns6?��v?�r^�vs�������V�n=�>�[�>��>��9��k�>�>?#��G������bY4�,Þ?��@~��?��;< ���=�;?w\�>ȫO��>ƾ�z������Γq=�"�>���`ev����CR,�Z�8?֠�?J��>������Aa�<�e���?��r?�������,~0�`�l�X ���_�GU�>{t�=�=n���dI�$沾�RB� +���8���>��@�z�=���>Qf���꿿Pٿ�֬�~S$�W1��H?u?u�#>: ����m�#����0���\�05��0�>g�>��������{�J�;�ϝ�����>Κ	��g�>TpS�����|B����4<�>�b�>d��>�h��0!��R��?I��}Aο����(��~�X?B`�?�l�?�H?L 0<o`w�Ŧ{��-� &G?��s?yZ?,�#��B]�'�:�%�j?�_��wU`��4�jHE��U>�"3?�B�>M�-�s�|=�>��>^g>�#/�r�Ŀ�ٶ�$���Z��?��?�o���>o��?hs+?�i�8��u[����*���+��<A?�2>���D�!�F0=�JҒ���
?X~0?'{�o.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?kٵ>vڂ?�M�=���>ky�=������f>���=��:��z�>��N?w��>���=���Q/��UC��.T����-�@�f!�>T}c?>�J?�Wt>�����Q�-I�?ӽ�/�0�G�H�2���	W޽��?>#3>�I�=<���ž��?Mp�9�ؿ j��!p'��54?0��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>@�Խ����[�����7>1�B?X��D��t�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?gQo���i�B>��?"������L��f?�
@u@a�^?*C�ҿ��ݾ�P�����;�\=I�$>N烾 8�={�>|����;ཻ�L>�y%>���>���>�$�>=04>-���/<�Q��X-��OЀ�%�0��+�j���mվ���<:�������o9N����¯g�K϶�jc�����f�=`�>?�J?i~m?���>���l��=K,��@���7ٽ�e=�e>�0?�t"?{�*?�_<�r��C�_�{T����о���i�>Ī�>�@?}� ?�l�>�ڱ=X��>���=���>ϕ��F;=W�S='0�<e�b>N�m>�J?$^�>�C<>��><ϴ��1��u�h�^w��̽�?ၝ�7�J��1��v9������i�=0b.?�{>���?пp����2H?���n)�!�+���>y�0?�cW?�>+��,�T�2:>X��ަj��_>�+ ��l���)��%Q>el?��g>�ev>92���4���P�U\���0u>>r3?e�¾=;2��Vs�6�D��پ��C>�2�>u︼[������ڍ��n%k���v=��:?�?c���e����s����2�W>��Y>�i&==�=}XM>�ȃ� ��r�A��9=[>N�i>�B?]->t��=1�>u˙��R�v��>\oB>�?%>�??|&$?�Rb��MB����,���u>���>�|>n�>��K��(�=��>|�d>M���t�
�	��?� X>��!�]��X��I��=pf����=a�=�K�(28�Y�*=Kz?>\��j����"��ؓ�=�\?��3?�H���=��־iz��+�� �?�(@�ۅ?k�*���CgD?#!�?Bż-�=D�>`)�>�7�͙u�2�?A����=��D��� w��ޫ?�?�?��)�dh����4�V��>���>)��Ph�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?[:Q>1ѐ?չo?'��>�2(��*�47��m䎿��=1 n�̲�>!�1>ؑ����9�.���@���s��3�|�1>]EO=/��>�t��^ʾ��>k���섨��`����>e6T>
t>V5�>\�?���>�&�>n�=yD�����������I?�J�?fC�x�o�μ^=ȍ�==�q��-?3�4?"LX�ǡѾ��>f�_?R�?U�U?L��>e
������t��5��q�,<e<>x�>3��>������`>��Ǿm7�cg�>	C�>����W�G����u�<.��>�#?���>�s�=˙ ?��#?�j>�(�>aE��9����E�ɱ�>J��>wH?}�~?�?�ӹ�?Z3�����桿�[�T;N>E�x?V?,˕>S���烝�YE�vDI����2��?�tg?T��?2�?�??H�A?)f>��Lؾ�����>��!?����A��c&����Jy?�R?�G�>�b=ս��ּ���=���5�?x\?��&?c�0�`�ST¾��</�(��LI�Jy	<y�;��5>Og>t����=8�>�گ=d5l�,�5��*U<g��=cb�>��=�6�(5��A,?i2>�{����=}Wr��KD�! �>o�L>���4�^?�e=�֟{��� r��b�T�e�?���?�D�?Gk���h���<? A�?�V?yE�>Ѯ���ݾK6�Cx�]y��X�Bi>n��>tU��������1^��z9��F�Ƚ�����>�t�>�L%?���>��X>翮>� >��'��*־~�پ�X�>%��+����������-R�M���ξ*������>doR�n�>w0?9�m>m#�>�1�>U��b�>���=]k
>'��>��=�>�z�<�J�=��%�_nW?E�¾��$��L���g���[?ީ�?ZX�>I!\�`.�
�$���?{�?k��?%#�>6j��޾��?b�?�W�K�?�==n"�ʇ�j�\$Ҽ}��<�Mؽ-E=y?��,���*R�ec��M�
?��?�X�=���������'��Rc�=D�?C�.?�*��\��v�k�c��PW�<o���U#�i���Ƈ���i��C��3���L샿J�4��@�<��1?�n�?����yӾʎ���Ut��#C�B�N>��>&;�>��>sA�>Q�꾻F*�OT��� �P�~���>nf?`E�>�[??��V?��Z?8J?:o�>���>��@�>� �?�M>n��>=N ?�?��?��?m� ?EF7>	����"��H̾!�+?��'?��>�B?��?���"��<��0<��t��,�= pi>Xeؽb����ݽ̺�q=�?���M�8�n����$m>�8?���>��>�����@�����<f��>?yƖ>g����r��u	����>l�?� ���	=��*>2��=������':���=����a4�=h�ȼ��6�f1w<mo�=}�=y�"�,VS;��;��;0�K<+u�>3�?V��>8D�>�?���� ���xg�=%Y>ES>>�Eپ�}���$��&�g�_y>�w�?�z�? �f=e�=˕�=�{��QT�����p���!��<@�?�I#?�WT?(��?'�=?�j#?3�>X+��M���^�����,�?l,?��>����ʾ@�^�3�v�?0W?�Da�y���8)���¾u�Խݞ>JX/�2/~����pD�j\�����P}��6��?���?)�@���6��t�C����P��N�C?�!�>UL�>�>�)���g����;>��>�R?~�>�T?��r?��M?tj>��1��ˮ�cS�����Ѻ�=�E?M��?�{�?FWx?@ԩ>Wy	>&�H�x�~���!����ʇ�U-$�ey>q��>K��>��>�.>��Ͻ��>��>��
�=	�p>���>r4�>��>��L>(k=M�^?x~*?|3�kC�-�-<�M�Pn�� �?���?�f-?�S>[.�n2y��*�F�M?��?1��?�+?�S%��T�=u~o���Ծ������>�a�>;J�>!w�=��=�u=\�@>i��=����:оBA-��u=,��>_�;?YV>�ҿ�𖿻�'�T��U	��{��+���YN�����>�ھ�ҧ�+��q���_�
��ˁ�Y2�q~��%��<���>���=oz�=	<>��\>��<��=n��=���<�h�v�ܽ ����>�qf>o�R�Q�.�����	=Z
>h�ʾ�}?±I?g�+?˭C?�Q{>Û>�32��ѕ>gނ�0�?
qT>�O����7�<��ਾT���5=ؾO#׾d����ʴ>ĦJ��A>��5>PJ�=���<���=��q=@֍=�3��a�=q
�=��=���=�J�= y>T�>�6w?R�������4Q�XZ罤�:?�8�>�{�=y�ƾo@?|�>>�2������}b��-?���?�T�?@�?!ti��d�>N���㎽�q�=,����=2>v��=�2�M��>��J>���K��2���4�?��@��??�ዿˢϿAa/>��S>�%>L�D�������bt˾�l��F�>k$��Ɗ�RW1>�G>����Zֶ��x]�̾{�� �=)⾙N����E=(�ۼ�=(�ʼ�U�>Y.i>��<bG��P=�=b�>b��=�Y%�����$�;���<�W(=/K�>�k�>���>��?�P5?H�U?�@�>�i���\Ҿ����͖>����O�>���>�V>��>�6?��?O{P?�Ț>{o�<�>���>|G�ꀿ��	�]Ƞ�g��H'�?)L�?#�	?�^>=U߇����Úl�\w���G?!A?�h�>3w?*��Z�ۿ��9�+�9�Jz�����m�9=���ic�<�<"�4�!5����<��>�F�>q�X>���=̒>>�v�>��>�D>U>�=M��=��=m!��̜:.>�䲻}o�=Q�;=,�=4�X=yè�um>*�W=��=u�O�l���EL�=��>�>c��><�=����p0>:��^L�V��=3��_�A�}�c��~���.��55��PC>1mW>r���W��Y?�\>�A>g�?�ou?׹!>-����վ�6��M�d�*�S�B�=��
>�P?���;���_���M�P�Ҿ���>W�>�ݢ>{m>e,�5?�~t=:^��*6����>qB��:�����.q��Ť��ß�J�h�͇��xC? 3����=�6~?Q�I?1ʏ?�A�>ǻ����־܄4>n<��yn=ó�4Ro�ե��`4?t'?I��>��龇�C��H̾����޷>W@I�(�O���S�0�4��;ͷ�0��>������оZ$3��g�������B�Mr�+��>�O?��?�:b��W��FUO�����'���q?�|g?:�>�J?�@?�%��z�or��w�=�n?���?L=�?q>d�A>��׽�o1?1w?�u�?�|�?9�?s#���&�>�#S�?|�<z삾��<R>8���=��U?0I?F?�P��}��z	��O��5�e��=���M��>@��>�IR>QI�=��<-��<}&�>*��>�r�>*YM>q�>�\�>������"�G$?7�N>��>8�??�
[>��>Hɝ�B���w�=����Z�2��Č���O�=0�<�ܘ�<�C��ӏ�>꙾��x?��L=!��:?[Ӿ1�=�w�>�(0��XN=�=�>=�=a)�>L��>�$?\�=�a�>ږ<>�DӾ�}>m���a!��,C���R��Ѿ�yz>����;&���o���>I��n���f�`j�-��4>=��M�<pF�?������k�&�)�<�����?+Y�>�6?�׌�O��Բ>���>ō>;M��Î���ƍ�h���?��?�;c>��>I�W?�?֒1�03�vZ�*�u�m(A�,e�U�`��፿�����
����-�_?�x?1yA?�R�<+:z>Q��?��%�[ӏ��)�>�/�&';��?<=u+�>*��-�`���Ӿ��þ�7��HF>��o?;%�?wY??TV�r0��"+>ϪA?�6?e�r?�5?�]A?�?�,?^?*>e� ?�?"31?�Q,?I4?)�">�=��m�"6*='y���M���aӽ�Dѽ2�ּ��=�Ē=|?<�����0=�3<0�G��L&����<\���Y�ú�=䡵=!N�=���>z�\?$��>�a�>��:?�4��<)�by��kf1?i�L=)B��侌�����%���0>u:p?��?)�V?}�~>b]D�պJ��>>w��>B�>	4s>t7�>os��}Z���;=+�=l>�=�?+�툉�V�����j�<�}>;)�>�I}>h|���2+>�]���y�d*f>��N��K��4}R��]G�1�A�v����>_K?B?�|�=���cƑ�#�e�:F(?'�=?8N?�~?x�=��ؾT�:�RK�Q����>RX�<��F����4���<�M
;�8p>����?���Ջ>|D��x̾� P��	K��<�7>��!����=% ���徯(%��Rl>��=K��%�(�-����M����=?K����8���\n���;�&;>��>%�>��A��zݽZ6D�������+=K��>�?v>� <=��^4����I͆>7sE?i^?�E�?�Pr�ԣA�V���Ef���ۼ�
?E0�>ƹ?��@>$K�=襲�����d��<D��y�>���>@����H�S�������$��Ӌ>n?%O(>��?�T?J�?�`?��)?W?��>Gý���7&?ᇃ?�[�=�tԽ��T���8�DF����>�})?s�B�c��>n�?��?��&?��Q?Q�?G�>ͱ �>@�T��>�W�>��W�0^����_>��J?9��>K.Y?�ڃ?��=>��5��ע�h⩽��=�>n�2?�2#?��?ۻ�>��>�G���\�=UL�>�Ya?���?��r?J��=X�?�3>j��>�}=yV�>e��>�1?�O?�ar?_�F?���>lF�<�⠽\���Ҏ�u�b��׻}�h<��S=�f������m
��l�<��:�,��mh����XI�������;Q�>T�s>╾��0>�ľ>��A>A>�������Ԋ���:���=`h�>W�?���>#�G�=�>��>(��9=(?e�?�?�&;]�b��#۾ qK���><�A?ī�=@�l�f~����u��h=��m?'�^?�W������V?K�k?����-�ޚ	��ؼ����a?&��>r�%=�\�>,x?�,�?2?�t��l'k�V���Ņ�R[^�L,>{�>�K
���H�[%�>�4?ui>΋�>)�2��=˾��S�n��~�>��?2ƙ?�?�1Z>�j�w���ֈ������^?m��>襾*�"?J��hҾ �������`�˯��{������3��j ��|����ս4��=�r?�&s?��q?�^?�� �&�c���^�̈́~�FV���=���`E��D��XB�[m�����q��%��hdJ=S|z���@�-t�?��#?��&�IL�>E��������A��*]@>�졾���"�=�њ��+V=R�=�a]�~�+�Rw��J�?�w�>|$�>L8?��Z��>�c4��3�ik���a!>��>��>�n�>��'<l�"�ޤ�4)þ��h���ɽ�8v>�gc?�vK?��n?��X1��t���� ��$6�dI��W!C>WK
>�Q�>�
V�����)&�i>�~�r��������I�	�U=�=��2?^�>g��>P.�?&�?�L	������x���1��"�<⫹>[�h?��>ߕ�>Fн5� �.�>F]o?-]�>ǳ�>H�, ,�ĺ2��
�8n�>n`q>�7?�?�>�y]��G7��I�������*��n>�Hk?ٌ�"�I���>q�_?,�T���=�{�>��L�9�b��r ���0�����>�5=�pD>)ݚ�Q�&�ڋq��i����!?���>w_���u#�$��>��$?�?q|>��?���>l�ξ����? 9L?�F?�fC?�{�>��<*��y�ƽ���q�=T�Y>��P>�[�;�!>�fW��K�F+��|=R��=�@+��Fv�+G`;.A��3����=�E)>	��
�>�O2��L3�����˾�7��������!�1y��D��)����ӽ�Kɽ��r��X��&���Qq�_��?bs�?FI���Ӿ����l�x�����d݈>yB|�thw�t�پ^����u޾�J��˾��B�9>[�Ad��8O���'?������ǿ����\;ܾ_  ?�A ?�y?����"��8�֯ >�>�<k@��I��ݚ����ο連��^?���>0�2�����>���>)�X>Kq>����螾�9�<%�?G�-?���>�r�ʕɿ.����ͤ<��?�@�A?�)�a��S=���>��	?�\@>J�0��J�����E��>�?�?�ڊ?8�K=d�W����֐e?��<F�F��nػ?T�=��=�p=l��T�J>�a�>&�'�A��!ܽ~�5>Vȅ>�$����9�^����<0]>�&ս�����I�?�a�WV�4o�q9n�� N>�lY?���>��V;LkW?�v-�r%��[��yo.?yk @�N�?�;>?�������>)��+m?M2?C�?�@����{k���9��ߨ=_���^��:ɼMB<?��P>��}��s�Jnu�
����p>v�l�ƿV�$�,|��]=wXຟ�[�]�罔�����T��"���fo���N�h=L��=x�Q>+j�>�!W>O0Z>ygW?m�k?gS�>1v>�L�򀉾�ξ����G�����(���(���mT�J�߾��	���������ɾ�=���=�4R�R���G� �z�b�.�F���.?�h$>)�ʾ��M�m-<lʾԸ������諒d1̾G�1��#n�]̟?�A?.�����V� ��H�?x����W?�M����8��=Ա�v=~$�>$��=����3�D}S��_0?/`?z����#��N�(> c�R�=�+?(v?B?b<�`�>}N%?
�*� ��<Z>>�2>���>��>�~	>����m۽{�?a�T?�r�g���x8�>^���d�y��_^=*�>�j4��u�q[>��<�%��C:m������<T?1F�>�*�+������&���t�=ȼx?���>8h�>�o?&�@?��<TZ��!Z��|�ZĆ=� Y?��d?vs>2j��[#ľ�G��;�%?G�`?�{`>��o�5aԾ�.�l� �1=?W�l?�o?�?�ZR���$��H�	���8?[\�?��k����A��-<=�?�?��>�>�0b�>�yt?�b�<R��0Ͷ�]�#�1B�?���?M��?/v=�\�?3=̈́�>b�>q�'�{�¾�N�^�ʾ\���?�<�Jx��S2��?���>?�+�?�>\�W������=�ٕ��Z�?o�?^���lEg<!���l�Nn���~�<8Ϋ=���F"�����7�g�ƾ��
�𪜾M㿼¥�>?Z@�T�Z*�>*D8�Q6�!TϿ��\о�Sq�w�?/��>��Ƚp����j��Pu�D�G���H��������>p1�=�N������X�|��6�i~�ɘ�>rbֻo��>ɧU��˯��	��L����j�>I��>���>�!c�e�c؛?����lͿ���e��*�b?�H�?�.�?m�?^U=@d��=y� �J�3�G?5Hr?��_?��*;��p�z0B�!�j?�_��sU`��4�zHE��U>�"3?�B�>Q�-�`�|=�>���>g>�#/�y�Ŀ�ٶ�?���Y��?��?�o���>q��?{s+?�i�8���[����*���+��<A?�2>���B�!�@0=�OҒ���
?L~0?({�`.�]�_?+�a�M�p���-���ƽ�ۡ>��0� f\�N�����Xe����@y����?N^�?i�?е�� #�f6%?�>a����8Ǿ��<���>�(�>*N>~H_���u>����:�i	>���?�~�?Oj?���������U>	�}?�3�>pW�?|��=7�?�J]=�����J�!>���=�1<���?ML?�Y�>"�=�a��l2�DE�0qF�����lA��~�>�_?*�U?7{i>�U��-<���O"ڽ	�J���>�=g�j��`E��~6>"�I>��=��[�-m���?�M���ֿ`N��\�,�z�1?*�>��>�z��z�|��	0a?���>�� p������qu��}�?+s�?�<	?ѥ׾@�Ǽ�>Q��>d��>�=ʽ�����E=>/�B?�����7\m�+��>���?E�@®?��h���?��1��Rx�o��7��ҫ>�A�>�??ܭ��b˳>���>w2�>�l��͘�T+F�oԝ>O��?f�?<��>�?�҆��z���Y=�A?/"�?���>p�3>S~�z�b>��>?k ��CB��Ȼ��[�9?�K@!@�?��?�!���o�@���V�¾ӝ��~'>^�C�X⮻ͨ���d�=���=J����e>o&�>�ە>��=>�S0>�dV>��=�$��E�� ����"��^Q�����'��v��e�����z�-|ؾ�g��jΒ< �'�	��S �������"��=�??Pb�?\y�?݃�>�� �����ӽƶ�7����>�lE=�f?H�q?��*?c�R=w���,o�g�r�C3��ʱŽ�r�>�݉>�t�>��>p�>�#B� ��>��x<R>�>݅�=5In��=5q>fA�>�� ?�m
?�r<>��>�ƴ� !���th��8w���̽+�?|���J��'���^���^��O�=�L.?�Y>g��gAп��+H?E ��l�*�+��l>��0?DW?�z>�e�U���>0��Եj��C>4c���l�щ)��CQ>�K?J�}>tn>� )�6t(�wa7�$�����)>=7?Sع�ڷ��nn�.G�H`��#�>���>p�<K �@����≿��b��';��K?��>)f�pK���%b�#派qly>C>� X=���=�K>߫��q��#>��n<{�'>�c>H9�><�=�$^=5j�>ś�&e�i�>=��=�z{>��:?"	?����޽�;��`���.�>Ǟ�>�+D>Z�=��I����=+�?��>��ȼ�ؽpؖ���{�S�f>���s;�� P��a�<<?5�A��=k��=V$�hy� 7�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿı�>D���(����Q�u�MY=���>a�G?�]���V��D?�N�
?��?�� ����
ɿ��v�1��>���?D�?��m��.��%�?��E�>�{�?��Y?�5i>�T۾ngY��+�>��@?a�Q?���>#���t'�N?���?Ɩ�?��:>O5�?pf?N�>j�����)��.����<�v�����>��=�ѭ��@��q��0����j����֐>aN=�q�>�����־�x�=�V��B��H^���>��}>��'>¸�>��?��>�5�>H��<�~Խ�F��:����rG?Չ�?���V����<D��<�;��%�?w��>��;��Ͼ��d>�Yd?��?�G?q��>\$"�X���ިɿI�������6�>���>K^�>*��<��=GʾwX�I�X>�g�>��D<�ƾ�f�=x%�>%�?ѷ�>��=��?/�.?�>���>�o7�D*���Q%��f�>�E�>�}?�pW?�+?��7�z��OI�����m�=gZ=��?P� ?��>�V��X��ɠ>��'�k���?NJU?O�^>��?�M�?d�Y?�d?+x>bE2��Bܾ�Β�ZW	>3�?Z����A��e��u��?U��>re�>�E��ۗ�7��<������?F�T?n$?���p�d�R7ؾ?<�g�6='�/����">��?>?s齇�>��%>,�=�`��I�/�<|��=�r�>�[E=ci0��μ�<9,?�iL���P��=
�r��RD�X�>D.L>D���{�^?��=���{� ��lp����T����?���?�V�?�����h�D=?�
�?b�?77�>�����v޾��྅�v��}x�Cm���>�>��t�h>�v�������8D����ƽz��W��>�o�>m�?} �>�tW>Q7�>�X����g+�ۭ�a��!
���4��],���=]��6���<�(����t��x>��/����>�	?�bb>X�G>7�>��<Y�g>��O>&�{>�ݏ>�K:>�D>�=�$��hq���KR?����Y�'�������1B?\od?�4�><i�"���L��H~?���?�s�?�9v>+~h�w-+��j?�6�>���Eo
?�c:=Un��<�R��޾�M2�� ���>�N׽� :�M��lf�Ak
?C0?�$��S�̾�J׽����߭|=�0�?�%?�.��U��n�O4^��N�#Z��O�z��G����$�%m��Q���@��� ��F�)�[�
=;�/?�"�?�U��x����G���f�!0��2h>� �>��u>w4�>
\>����#;�~]�kc1�Ɛ���Y�>{?���>��I?��<?�P?��M?�}�>�Ӧ>?���ȟ�>�1�И�>#�>��:?��.?=d0?V[?H)?WY`>��뽄�����־�k?�?��?��?I�?�#���Y�� ᧼\Ka�Ёr�4/��T�l=���<�0ս��e�ޘ`=��W>{J?�A���8�����j>zl7?�w�>i��>X&��!_��Na�<���>�
?�/�>� �Ozr��h�i>�>���?o���M=��)>*�=����ysú�X�=3¼��=����r)<��x!<-ڿ=�=L�o�7����r�:D�x;2԰<QO�>H�9?�>�iS>�]�>{�*#��G�=GO�=��o>��t>����{m��z���n{�?��>7�?��?��/5>�k�=�J��萾�P�u���+>WH?�0N>f�a?Sb�?N]T?NF?`�>A5M�����ۇ��⧾�?� ,?�>���ިʾ騿c~3��t?lj?�Ba�6��S6)���¾�IԽ�'>H/��~�.��'$D�����x���Й���?*��?��A��6�'�����YH��"�C?V1�>�\�>�	�>i�)�H�g���=E;>x��>�R?�>��O?yM{?ë[?��T>�z8��������&\.�cb!>G@?U��?i��?.-y?ښ�>��>N+*��,ྡྷ1��,��b�t߂�<�T=�2Z>C��>"��>_��>���=��ǽB���q>�l7�=Nb>i�>b��>��>d9x>拵<��E?@��>�ɺ���C����a���l�)lq? �?�'?��<����3F�������>��?���?��+?p�U���=����(E���p���>[�>a��>��=���<K�$>���>��>Ư������=�Up��z?}D??��=��ſ��q�Nq�7q��m<����Xc�r0��}�X�=��=�I�������]��#������2��@�����|��9�>-%�=�}�=�u�=f��<�ϼg�<r=D=��<�=�m��o<��;��彻������4K<��K=[���'˾��}?"�H?�H,?F�B?_�w>P>�05���>S����?US>��K�;G��0>�u0��=Ǖ��/ؾ=PվO�c�򖟾/b>ߖQ�%�>�R4>�T�=9�<�A�=�i=2��=e�����=L�=�P�=;ج=̌�=|>�Q>x�?�$��t���8f�I9�=(�g?�B�>��6>���?k?���>	�Y�0���Ҧ�LG�?��?r\�??�\���@�>�y0�3��=� #>ŏ��A�m���=�rn:_��>���>�ZD�@g��rv����?t@E?Ϟ{�G(ſ��=�x8>e��= �R��a,�I�T���J�(V�^�?��6�/ǾJ�t>�,�=��ݾ��ʾ��F=X�>>+
�=�x%��\��l�=]����9I=��=bu�>yoH>�O�=�^½���=�9~=ͅ�=KKO>^�3���I��>���=1l�=R>}4>M�>��?��0?�c?=�>3m���;�¾�*�>���=Pu�>�(�=I�A> �>��7?	�D?��K?p�>�0�=基>K�>��+��Km�.S�Oʧ��q�<���?#��?�>��G<׊A�%����=���ý�0?$M1? 	?%�>����߿c(�<.�鑂�Q*����4����@Q|���<M�%��H
��>��>�X�>o�>��n>î9>��G>�'�>P�>RNT<U�=<��� 7=��?�T�<��<tծ<�%<���)�B�%�����+�ʯ��B=���=>�>�=>���>/�=�)�� t0>k>���K����={�����B��<c�D0~�;�,��..�G+J>�6S>�Ŋ�Ñ�� ?�UV>��7>w�?]�u?i>D����о#���Gb��P��ָ=���=�>C��W;��[`���N��fվJ��>A�>��>f�l>,�O#?�)x=D	�[\5����>�l��9[�C��3q�@������oi���Ǻ��D?SB��'��=~?0�I?�ޏ?���>���Y�ؾ�#0>�V��]=���q�Zj���?'?ބ�>�쾤�D�
���<�)�М�>P�߾5V��F��1Ua����_۠���л��Ǘz=kB&�<6���8���`��聑�U	?��Z?��?C����?M�3
�mG;�U>4Q?�_b?5�>�+?V��>���c�(�mfN>a:q?+��?�ǽ?�%<��=��ݽp�>��?���?䄏?Ц{?Y�s�
�>2N�<���=�TȽɧ=���=��=t4>��?h�?E��>ᙽ0�v̾����l�\��޻�*�=#rz>�c�>3SQ>��=��d= �=��h>+��>�7�>U?[>��>(��>�t����O�%?���=ر�>2?}ي>@=����i�<�j��>E��T0�X�Ž�zֽ�A	=p>:LG==K�
�{��>�Ŀ���?�QI>�����?��kO�I-O>��K>�N׽�p�>�U?>�r�>��>�o�>�u>���>�e&>L���)>�p���D�J�P�Z�d�iξ��X�h����gϾA���f!<�s��fھ"��䂿����);>�w�=�Տ?m��o2U�U�$�vs�S�>D�>�@!?I*��u���S�<�?Kώ>�9+�E��'��E?徰>�?� �?�/>H{�>��u?�B�>�j/�^-ӽ�9�r�k��ՙ���X��Ad�}����S|��e���=x�k?�Qt?��Q?�ĳ�T@>۴�?n�
���%�*�>�0����� �>�v>>����U6����:'Ǿ��^�p=~>?���?�@?����V��9ƨ>�5T?(�L?���?�,?���>�&�gMz?q����:?q/?�HU?-�??��?T��>V�>����
}>�ǽ@����qNY�&0>)X}=ͻ<y�����=);I=ᬪ=j�?>��b���2�*�s�c�B��=Q��=a�0>�+�>�]?2)�>.��>�
6?���9��ۮ��0?�M=�넾mؑ����������>�zk?��?R[?��^>Yq=���;�_�>��>��'>=7S>�I�>���g�Q�UC�=��>jb>��=��\��:��hV
�ᄍ��q�<�?>�}�>y7>@��Nn�>����a���m>i�@��w���]G� �\���>����Z�>WjQ?�.?9�z>��ؾe���_<c���?L�?�z;?:�|?zCj>X�Ͼ_�1�|�%��zY��l>�B<�P��o%��lm��0�5�]�#����= q羱�þ�~>�»�9޾�4f�r�R��K����U�C.'�"���bb�|�Y�X�=�>`�̾5�)�F���ρĿ�TS?�x>5���-��$�_v-=�?�>�I�>�`{��� �/0�A���~٘<m�>�==ݶｺ����K�I}��P�>c�G?��\?e8�?�O��7p��sB�M
�]e���6���>?y�>��?r,:>�&�=BR��@��Wf�)�=�H��>���>����<��T��T����� ��W�>��?G&>e�?P�P?�?�Qe?�h*?9?Q��>@�߽������&?�o�?��=9o����N�`�9��@��� ?@)?9�6�
3�>�~?�?-3? QJ?�x?�?�=<n�`�H�j��>5h�>�SU�ps����x>C�D?0��>��\?q)x?�y'>t"0��a��9��>dQ#>I]2?'�'?�q?���>���>�r����=�>��\?��?!s?�ɵ=��?
�+>e�>i�\=���>T[�>�?��P?�Pr?_�G?14�>�U�<����I4��u|�M�z<� :<���<��=[M�<��kg �Q��<�`<�p��hֻ�G��=�	�;1$��&\�>?>s><ؕ�Ra0>�ž���^9B>����ܸ�������>;���=�&�>��?���>X"����=㫼>$B�>,���(?��?g�?�[#;̲b��.۾�L�z�>��A?��=P�l��z����u�~�c=��m?M^?��W������W?�m?�����ƾM�ľh9����,�M?�#?8���T�>N�M?\�?��?W�g��/]�C����#��hSy���$>f߉>�01�Z :��L�>dV?���>���>�6G���þ �K�F���>'��?:D�?,��?xg�>��a�����2��<���*^?��>�즾�"?%`ܻ�Ͼ�r���p���F�I���.��u=�����C�#�䓃�Luս�D�=Z�?�s?�>q?��_?� �q�c��Q^�S����V�N�n��~�E�H�D�UkC��n�����r���E�E=KP���,@�u=�?UA$?�+�V��>�J��m4���};R�5>ö��!a��{�=�;���j]=��j=��e�]�+�I���H^ ?蕿>� �>�.=?:SZ�8L<�'�2�ч5�>����2>�>|t�>_��>��H���3�=��C�˾\���9Eｘ3v>׷c?�4K?,wn?��$1�XD��{� �U(��,��B�C>�^	>-W�>��W��* �&��?��r����dq���]	�L��=�]2?�"�>|�>B��?��?؄�g3���w��s1�D�s<��>N
i?���>��>]�н,� ��X�>`~?���>ir�>�-���}9��V�u����>�h ?�! ?���>6ʸ���P�{��������[��B=+Y?m����%J���>%,=?��ս��>'>�V��f�"���j�篰����>Х=�"Q>�þ��7�ل����k���"?#�>�cW�q�1���`>T=??$Dn>v�?\s�>�ؾ׆�g�>��H?k�L?�E?.��>txT=�t���줽����=r�>o�>˺�=�`�=F+��<~��"�>��/#=�R[=�b<��6��?�<+8��������=W�	>�׿<;�1�������Ѿ��
��v��K�G�F0���gr���Ͼ�/$� �9�.н�6=�[��!c���0_����?���?�T׽"�`�~q��̒y�tc�ezu>q�����������+='������.��c,�	�c�ݙ��]���K�'?�����ǿ񰡿�:ܾ-! ?�A ?0�y?��3�"���8�� >=C�<�-����뾮����οD�����^?���>��/��l��>ܥ�>�X>�Hq>����螾32�<��?4�-?��>ӎr�/�ɿc����¤<���?1�@}A?>�(����RV=Y��>q�	?k�?>�S1��I����T�><�?:��?�sM=�W���	��e?П<��F���ݻq�=�:�=�<=���ߕJ>�R�>5���SA�Fܽl�4>�م>ل"����5�^�՛�<Z�]>�սL:�����?!J�e�|��*����WΦ>&�n?:�>fa�z�(?��N��0���Ih�IK?n�?�.�?Z�H?6�X�D��>O����2j?��??���>�g�HV��^�>񤥾��̽����s���7>Kp2?[=�>� ���:h���轇�>�� �������1%�u�~=���:9����d^������U���r�{����;�=�a>h�9>_��>�,K>��E>��V?�[n?���>��+>	� �몃��\ɾm���⌾_{��o`�e���l��q;��Ǿ���ۉ���!���&=��#�=R�ϒ��?� ��b���F�i�.?G]$>��ʾ��M�j2<�aʾ̸��V*��V���5̾J�1��7n�-͟?)B?�셿}�V���(�ψ����W?�U�����ᬾ���=�g��p�=��>�9�=��� +3�z�S�h0?�G?�����V���)>�� �=�M,?n� ?j�<<n�>�"$?p'�A$ܽ]Z>i�3>��>���>�?>�-��G��>?�T?	���̚��Ԏ>�t����x��J^=��>:�1�($¼>U>�<)����j;�yX����<��Q?A]�>"�%�T�T��q��q�"=��{?�j?/��>xwp?�\E?��������kka�
��Hg=�:^?j?���=v"l��ҵ��m���G?ۦ_?D:>>o���[ݾIz����&�?l�?8q?���m%��u��������B?��?�t���p���N9�+3��-?��>9w�>�Hk�f��=�ρ?�=�<���������-3�P�?a�?���?��=H�3<��6>���>O�?��f�N���k�"�BS����<W�+?���6̙��A��DR�ת�?�,�?\^�>!Dr�<>�}��=�ٕ��Z�?m�?o����?g<f���l��n���{�<�ͫ=w	��E"�����7���ƾ��
�&���迼��>AZ@�T�Z*�>�D8�P6�TϿ!���[о9Sq�{�?e��>��Ƚ����;�j��Pu�v�G�G�H�:����X�>ъ>埔�����{��g;�^&����>���WY�>��S����G����x0<�Ғ>b�>б�>Iq��z���̙?�����Bο嫞������X?�l�?�x�?oi?��:<a]v��{�Jo��4G?�ws?�Z?��"�D�\���7�%�j?�_��yU`��4�sHE��U>�"3?�B�>V�-��|=�>���>g>�#/�x�Ŀ�ٶ�7���Y��?��?�o���>p��?ss+?�i�8���[����*���+��<A?�2>���K�!�C0=�NҒ�ż
?T~0?{�f.��_?<�a���p�]�-��ƽޡ>7�0��h\�Z����pYe�����Fy���?�]�?��?e����"�N5%?��>����.Ǿm>�<х�>�'�>�/N>h{_���u>�
�#�:�Tj	>��?E|�?�i?���������V>��}?�$�>6p�?��=R��>�S�=ڬ��h���.>e��=����3?�G?Ku�>��=�|5���*��F�?�P�G�/�B�e�>�
d?�0N?sR>�����L��!������xF�
����5��м�4��g�P>}\A>��>��9��ʾ��/?�D�}߿/P��9�D��gl?2.�>�u?�l��о��[>ˉ�?_)>���s����"�����;�^�?�@�?�c�>]��}&��� =�T?F�>�1r�^�H�e�ξG��d9m?O�;�Ik����i��Q>E��?N��?w��?�+N��	?���������_��	=0�b>�=�8?x���w>��>���=�;v�����a)t��c�>V%�?(`�?��>�-l?�uo�kPC���(=��>s�k?��
?�f���3���$<>n�	?���A ���V�ee?z�
@�@@e!^?҉��~@ؿi��R3��Ԍ��0�S>�K�=��<�|����<��sN���� >p�>LJ�>'[R>~o>?�>w�F>r���/�����;��>�X���!�T�筸�EJ��;>����%���4���.5�4�����Ž:����"�G���T@>��A?q�@?my?w��>����4���G����so�^$>ps>�UK?QVH?��?��==c���JV�aLf�6������6�?淸>�z�>��>�C�>�{;�]�+>{'W=�B$>	?4>l�<>�'��8>�in>b��>��?��>�C<>_�>;ϴ��1��>�h�Dw�x̽8�?H���1�J��1���9�������k�=,b.?�{>���?пr����2H?"���f)���+��>j�0?�cW?��>G����T�:>[���j��`>�+ �l�l�)��%Q>Il?O�h>�Nw>x3�%�6�bWO��y��T�y>-�6?��AU5���s���H���۾��R>a��>�}8��x��ٖ����Di���h=� ;?su?�Ϻ�M��*�w�����WQ>��\>4�=jp�=��O>%~��`Ž��E���2=%��=֖b>�k�>���=���=f=S>BA���jH�./�>�H���>�(?iO�>Ţǽ Z)����%ٽ�Į><�>��c>q$	>�pP���y=,
?���=���<Ҫɽt�5��E��i�>�����pE�eݴ�s�<6����B*>1�<YT��W!�:�<�~?���(䈿��&e���lD?U+?Z �=t�F<��"�E ���H��E�?q�@m�?��	�ܢV�@�?�@�?(��R��=}�>׫>�ξ�L��?�Ž;Ǣ�˔	�0)#�iS�?��?��/�Yʋ�;l�|6>�^%?��Ӿr}�>�F��+)�� ���L݆��&>o>?|e?��ʾ��>f��}4?v@�>Kx��Q���˿�|?�?�?�w�?�1�?f������^�j��M�>���?��k?��>���B�澹�?�e?�o$?���>��%���c=�sF?�"�?�
f?�6>Kj�?M n?P��>�*�u#"�M����g�]�Y>�
E����>�+<Ę��ΝG������x��^Ʌ��5�k��>,�=���>{����^z��N�=M��<Q٥��v=��>]�}>z�8>=>�{?HN�><��>�h=�q��_��}o���G?��?�Y���!�5�=<pu�)�Z�X�??��?߄<��<��7>�E?�Ơ?��3?��i>���	ݤ�`�ȿ)@�������>�w�>e�>6ש<t�=���ď��G^�>�lY>��u���ʾ�����Ǻr�>n{?��>��>�e?��*?!�x>�>yC�����;E�\��>J��>}6?�*z?�5
?;Ǔ�1�/�?���Р���h�� >g�|?7!?�`�>�{��ށ���ɛ��䟽ak���Fz?{[?e����?���?��M?NaM?�H�>����˾�8
�\>�T!?*f�&@�In%�����D?��?��>�O����ҽ<��+������?p;[?�.&?@!���`�uľ���<y@H�Ùg;k��:�π��>�>�Ss���=4�>ǚ�=�o�z|5����<��=��>��=�0�'���N
)?���%�u�ddN=��q���<�ck�>���=��̾&�R?K�Y�@�v�KԪ��z���^H��?���?�\�?-����e��5?��?P�?_��>T���b��޾Z�&�u�S����~�=+ϩ>�;ԼB1�HР��<��6^���J̽���?'�>���>'E?��>BwG>z��>=*��}#��y�����]��N�CV8�f,����I���v�"��?ݼ�m��2,x��M�>oה�)�>�V	?!�b>0�>Y��>]����>�F>@�z>��>G�^>�X/>d0�=p=D<C�ֽ�KR?����'�'�j��ڲ��e3B?�qd?61�>i�1������k�?���?Ps�?�=v>�~h��,+�on?�>�>_��Jq
?*V:=�6�T>�<V��:��;4��@�窎> E׽� :�xM�Unf�_j
?�/?�����̾�;׽%s��x��=bS�?0� ?�+���T��`o�?Z���P�ZG=�gx��镾yX!�an��<�����2����.�8z׼0H,?�b�?Q� ���|���g���2�U9o>GD�>�/�>7�>��->%����4���_�&�+��&����>��?�>�FB?A�L?�n?I�>?��>��>�(�����>�D�����>���>�R?��,?�<?�N?�s?��>�������:���]G?�.?+*.?Tj�>��?����m�R;h��\{g� �c���=/�;��н���F�=��>�X?���Z�8����]k>�7?��>���>T���,����<u�>��
?�F�>  ��}r��b��U�>]��?�����=!�)>��=:���k�Һ�X�=���8�=17��8{;�I[<���=��=�
t��Q��N��:���;�o�<��>:6?��>�y>3�&�2%��ھM�>��q>k�>⽒>�O�{)��r��8����x�>�T�?jM�?`<�	�=
�>뮾M���֍���d��"�6�?�QO?ǟL?4��?,hr?7J?kB>_� �����|�x<z�*$?m!,?���>4����ʾ�쨿 �3�(�?�`?m9a�T��4)���¾k�Խ��>JX/�D(~�����D�ټ�����a�����?��?��A���6��|辴���IV���C?x�>�[�>��>��)��g�`��6;>���>�R?E$�>E�O?4{?T�[?�_T>k�8�,��rș�.2���!>�@?Q��?n�?cy?�s�>��>Z�)��(྄X�������Eނ�%�V=y'Z>ō�>t'�>��>h��={'ȽO����>�5�=��b>���>���>�
�>�w>�t�<��D?��>���	�@��W���U�Gkq?=։?�*?\ۢ<5%�{�J���	�>#�?~��?p.?��L�A��=PX$<,��Jn��?�>I�>��>���=%�=w)>���>�*�>�{B��B@������?�E?�v�=
�ǿ5�s�*�s�~J��$��<���� 6��p�½f'W���=�䡾`��
��1"G�^���6����������z�
b�>6�z=�
�=�1�=q<\E뼼]�<�j=���<�T�<�̈́�ߪ�<�K%��A�X;���O��ec<vt"=NZ[��jʾ�M{?�I?U-?O�G?��w>�?>�O�u�>�K���?�b>з�ޱ��͞8��p�������xپ3ӾA!d���}�=�af���>��4>`�=�C<��=_�d=�0�=�d�:��=r)�=���=���=,I�=�>1�>n�?�Յ�Z�����Z�s43���P?d�>�5>�����C?��l>����:Ŀ�(��?���?t^�?�;?�kW��
�>o��/)<�A>������<��0>9�R�>w�>��S��5��#�C��(�?��@610?ƛw���ǿ�>��8>��>�zR��1��[���b���Y���!?$�:���˾:'�>w6�=��޾Wž�>/=#�6>Y�_=� ��e\�n�=*��AC=�j=@��>==D>8�=>5��9~�=C�K=:Z�=�O>/���8�=�Đ*�I24=�3�=h�c>l�&>���>��?�)0?�d?b��>�,m�r{ξ�����l�>}C�=�T�>^u=�!@>��>Ճ7?L�E?��K?��>!ވ=���>kD�>�,-���l���ζ��+��<(��?׆?Ꮉ>m<<2A��+�f�>���̽N<?�r1?�c?qҞ>�K��lο�A��R#�a�Ǽ94��aھ�fd<��G������H@���>��>sw�>�g�=K�[>�z�=��=�з>�><�W=�+��α�"V�=�
>��<��_��ҿ�^��<z�O=iE�O<5ҕ��ļbk��P�����=���>�H>_��>)O�=���q/>7Ԗ���L����={S���*B��5d�/G~�!�.�-!6���B>�5X>�d���.��o�?A�Y>�H?>��?)4u?f�>r����վ�J��;e��bS�5��=S�>.�<�v;�L[`�}�M�!yҾ���>:�>"�>1�l>,�(?��@w=�	�UO5�?�>^��7��](�E3q�ED������Ui��I��D?!A��$��=:!~?�I?s׏?��>_9��Xwؾx40>x~��Ͷ=��dq�sn����?x '?,o�>�#� �D�h������;��>�T����V�񴐿C�3�F�
B��=��>�6ܾ�E��KS"�dd���8��_�k�P��+�>�1R?�?��Ծf���~JE�R��>j�!?Il�?M<�>��&?u?+}�k�վw@1�	��=�L?ey�?��?�]�>�۽=����ys�>��?���?t��? �s?�}@�5��>τ;��>�ٙ�v��=
>�	�=���=w?el
?��
?�^����	�9%���c\�'��<�*�=c��>}S�>�r>���=bf=f��=�Z\>�ў>a��>��c>s+�>W�>�q�����&?~�=|�>\�/?E+�>S+Y=H�����<�Z��lG�ţ*�⎯�4�ҽ���<�ِ�LH=g��g��>�vſdX�?��Y>�H�6�?)����,�bH>�'M>JI߽���>_P>( u>�Į>�ף>J�>�ˏ>U�&>�ݾ��5>;g���(�N�J���a�zEؾ�as=��������J�@���C��Q��	�P�{�,���M� R�/B�?�Wu�V�����h���>���>@??�w�ʖ�=b�=�c�>z]V>����ڏ�[�����Ծ�.�?,@��>��>��]?�
�>gҽ���M���X�%�d��=L���W����$(m��\�BSB�t�?��i?pT?F#��'r>���?�==���W=�>La��Y����>��>����K������)�о5��qF��%�q?,
s?4?n%�=q�[r|>̘X?�l?�߬?7|?�"?��?��gI?fj�[� ?p�?r�T?U�1?Z[?�>�=΋�=$qL�\:>#�Խ�r��%�R���L!�>,5s=+��=}5����1>�g�=�F=�o�=�C,�]�Ҽ�4���9���0=90<+�=膦>z�[?	m�>�4�>6�5?*8�e�5��±�;'/?�g7=Q���t���ा9��0d>y3k?���?KOY?�6d>��@�@B��� >b�>��+>��Z>�>����8@�DǄ=:�>Ű>Sڥ=�(=�_�~�V	�LR�����<-v>�`?�!>Bװ����=��¾x�ce	?Až�
��?���X�S�&��Qx�Y�>mZg?�X@?�W�>'ۚ��a<G~b����>��U?S�?n?!k��ڻ�\�O�/-�^��E�>����y� �����1�����p��;^KT>�m���U���z>����Zؾ[Nk��L�M����=�Z�:�=�V���ܾ@_u�>� >ҵ��[$��P�����1WG?q=yV����k��ڬ�jm>�i�>�:�>S�`�eJ����>�
B���X=��>$yU>]���X���*E����-�>��F?8�]?��?�v��>�q�@iA�r���H���f�S��L?�B�>=	?2H>�š='��Q����d���C�7��>:�>]�ZG�kD��'P�Qv(�*��>}R?�f!>�;
?�HP?\	?!�`?׽*?�j?�9�>�սɁ¾2'?Ӥ�?a�E=��ؽ�QO���;���G�� ?6�? (��5�>�
?9�?oT/?��N?�?���=�}
�xtI��%�>(z�>K'R�oͮ��!u>%�G?`��>�_?��?y�(>�&0�������Ľ)�>m�=>ܩ2?/�$?��?�W�>���>�����4�=ɦ�>�c?�.�?��o?�Y�=?	�1>���>T��=ƣ�>M��>?,SO?��s?`�J?��>��<�Ƭ����.t���N��O�;b�G<��x=Ԏ�G�t����,��<�;񪷼�Z~�8��)E��3��`��;P-�>r>�链G�.>m�ľF����D>�9Ƽ|ś����;�=����=�P~>�� ?=O�>r�!�b>�=���>���>©���'?�D?�?�&;��b��پЄK���>P�A?��=� m�U����t�$Bh=�cm?K�]?h>U�Ѥ��|�R?z�u?��;�m���Ծ�j���}�2�F?O(�>�:�=�g�>
� ?b~`?	�?�q��V�q��У�Q���,���^>>B�s>�[���\����>J��>
z<�u�>��`�a���l��<��+��>�E�?�~�?`�?�
Y>�+������R�����z]?���>�̥��y"?���X�о��� ������Cu��sq������Aۥ���#�i��{�Խ���=�6?��s?� r?F�^?���c���^��~�DpV�������xF�:D�V�C��mm�Z�H��������D=�Ml���;����?�w%?MC@�4&�>Bǟ���pѾ,a>!����J��U�=��`�}��=�No=�c��p@�5���& ?`l�>��>��>?f�V���;���*���:�C�TR>I�>�ʖ>DH�>��a�3�	��Tӽ+�þ�v��>��v�w>��b?�GL?�{n?[���.�T������=IE�����'�@>ϵ>�7�>&CR�,G���$�*~=�TGs�(��j���=	���=��3?l��>��>Z��?�X?b�e޳��s�0��W�<bu�>B�i?Q�>ͩ�>Nnʽ� ��>n�s?D��>��>T[���(���Z��:k���>#��>-?{!�>Zؽ��C�mᔿ
��,?F���=?�?�����vJ�x;�>�,U?5�"<��=kM�>փ�h����;�o�(>��?�=�=���>�'��I���|���W��H)?.?NC����)�`Ry>�"?��>�ܥ>h!�?��>w�þ�Km�`�?��^?�$J?v�@?o�>(�=:���:�˽�)�U%<=�z�>
�V>s<p=8��=d0��\��B�[�B=g��=�c����½��w<H��Gab<��=�<6>-�ҿ�^?��c���/�F�־]������������T5|���K����뇾�.�9Փ�Z�W��-���ן�?ň�16�?A��?B�<�)��Ü��ـ��k�(��>r���r=z��I|��!�W��T�|Ъ�EM5��d�(~��W�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾x1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@�fA?k�(��J�7�T=$\�>�z	?�A>��2��o�O�����>�?eƊ?�+H=��W�����re?Y%<��F�s�o{�=됧=�=F���cI>Mo�>D3��@���ܽ�q3>���>�I!���O^��=�<��\>�Խ嫖��.�?�)[�>Ah��?0�d��>�T?Q-�>�X�=�,?�/G�P�ο�`�}CU?z��?��?�~.?�ͱ�n՘><�Z R?�6?ڦ�>��*�;�u�t>�=��"�أ������Y�N��=\)�>E� >�����
���N��! ��f�=Wh���~��������{=b�<���gf����^�WX��;�,���C�=p��=�?>��s>�M>�� >�T?�x?5��>��	>�#��ӕ�'�뾓F��������U�����lk�r��Hn��q0ƾ)e�я�"U�����=��b�=�4R�J����� ���b���F��.?{M$>n�ʾl�M�Cs+<�fʾO����˄����%<̾�1��)n�Yɟ?��A?(�����V�4���y�Cm����W?�Z���묾l��=m���9k=Z7�>j��=�⾞3��S�q0?�D?Ğ������~�(>�����=,�+??�3�<̟�>Y�$?��)�����\>��3>���>R��>4	>�;��+�ܽ��?3�T?�I�ؽ��c�>���v�z�ň^=�>�3���ؼ��Y>r��<������P����h�<�R?͗�>��;���2���JȠ�.�=�*�?n%?��?��|?<>?��JḾ�w��a�(��lռ�<?�z?#��=�k��~q������?&�d?\K�>[���������p�=?+p�?��*?<e�<X������N�A��_�?�?Ql��ҫ��"7�Qn��'�?ŕ?x��>x�,���>��W?�i��F��-Ŀ"��>)�?j�@(s�?NK�=�ު�<ub>���>Y�?ʚ��74�LH���w���	<g?b�����CP�1Y	�*�?���?i?�|7������=bٕ��Z�?��?����-Lg<����l��n�����<�Ϋ=��?"�\��/�7��ƾ��
�b���Y࿼B��>%Z@�U��*�>,B8�=6��SϿ)��([оVq���?���>��Ƚ������j�Pu�H�G���H�٥���N�>+�>�,���l�{��q;��Y��q�>~� �>��S��)������̾4<s�>̬�>$��>���?F]���9ο����Ě�?�X?Of�?�l�?�u?�N:<D�v�՛{�9Y��.G?^�s?Z?@i%��+]���7�(�j?E_���U`�Ў4�RHE��U>#3?C�>�-�2�|=�>��>g>�#/�v�Ŀ~ٶ����;��?��?�o����>`��?�s+?ii��7��|[����*�r_,��<A?O2>����!�P0=�mђ�ڼ
?.~0?�{�(.�X�_?�a�$�p�y�-��ƽ�ۡ>s�0��e\��P��[���Xe����@y����?A^�?\�?е�� #�\6%?��>v����8Ǿ	�<���>�(�>.*N>@J_���u>����:�]i	>���?�~�?hj?앏������U>�}?!9�>Gz�?8d�= �?�<F�۾S��=�G>Ց>C�>*"?G??��?e�%>o����S�ј`�"�N�����=�s�u>(h?	*B?�7Z>8�<��:��\�G��������;�짾��ؼ�J��ϛ>B>���=�_��$�Z.4?�_-�udؿ�;��8s>��Xk?M��> Y?�޾�蜾Z�*>�9�?C�j>y~
���Љ�����y�?�y�?È?£Ծ9Ȩ��BU>��?�d�>�h��i���0���p�'=iD]?o���S㏿��h�b�>���?�@�5�?܄b�v�	?��!�����~��v�/���=U8?���bx>��>��=�Nv�ˊ���s�-�>,Z�?eU�?��>�)l?�n�@tB��=<=�K�>,j?�a
?Ǒ�����U�D>�c?����R�������f?@�M@5^?c���q�տ�{��{ Ծ�v��� >�=}�=`勾E5r=o᫽̤ҽ:?@;G��=:�>V�>_C.>7->\L+>�=�V��o�'�$螿n��$�]���!�����r����/�Dyp�R��_���N0����^�`u�%0%�80@��ͽn᷽.B>h�C?�k?[�?�=�>�E�=��̽[��n~ϻ��^����=P�">�_?=6?�M?l�>A2���Iu�5�F�α�<t��_�>��>�
?|u�>Hq�>�x�q+�>�"��	�p>�v�>��4>��%�Ӝ�<h�t>�>�`�>*�>]Z<>�>>˴�,��=�h� -w�Ta̽s�?� �J��-���G��V���B�=?_.?_k>����@п����y,H?����f$���+�>g�0?�]W?�>����U��5>S����j���>�����]l�Ā)�?'Q>�`?�|�>WP�>E��!���H���m�/�c=�H?�Ӿ~���Q�e���S�O�����>�>��<<'��	��6�m��Fq�gj���>?T��>cDT�D�b��HN��˾�>]�>���;��>�ח>�K�f���г6�^R�=5��=�˞>��?#8>�\�=��>~i��[Y,����>��#>q[�=�a5?�?�~B�w���Ӕ����� ҁ>
��>��s>~�=�^�a}=��>��`>4a���1�⽢ym�#g>Ӂ��	�j��,K��=�P���>NR�=[��q����<�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>��{�����f��|k��;�>M�>C�^?����O>�����i?��>-�������H̿��P�|�>���?qn�?�[�����Vt4��@?���?�N�?&�x>!��b��y�?1
t?̴)?1�?���Ռ�'F?�?8T?t�Q>�;�?@�f?��>-�����*�#�����w���'>�+9=S�>�a=H���.��_���}����y�-���"�>�J$=~]�>z���+�[t=�S�"�Ͼ�w �yf�>吃>�C>{TP>j��>E�>A��>D�^=�����:k� �ھ��K?ҥ�?����OW>����=ʂ@�[�]�W?���>��>簾 �=�,?��?�L?Y�j>��� ����ſ�����	���>IK�>�Q�>ra>�k?=�����;�^r�>]�w>X0���z¾�����V����>�h?��>�?z>�� ?�{'?
�S>�>�\D������@���>���>6y?M�?�/?�q���l.�������q�V�g�P>~v?��?��>�G��An���F��Z'������Q�?��f?���3�
?E2�?��G?�HD?Z>M8�`��"����>7�!?6w	���@��]%�����?ӳ?��>Λ���Ƚ�7޼v���%���^?m~[?d�%?���>b��ľP�<�f��3���;ƛw�&( >�G>Jr����=X>#n�=Jk��v3�ͷ0<`��=�]�>2��={4��t��
7?j�f��P���T��.$������7�>��(<|�����"?���\�J���ܬ��~s<��?5m�?1��?��K��?f��?.�?��?�&�>䖇��3� �"��������q1Ծ��x>Nt�>���=����0���᝿{jk�-y��a+����>,��>a��>K��>�1>���>gؾ%�)�������P��t�n�F�s $��(���<t���M��uԽ��žAti����>,C׽s�>���>��>aC->xH�>��b��8�=��>k-f>Bڲ>�@L>>���=�=�n��KR?
���۾'���ɲ��3B?�qd?71�>�i�������1�?���?3s�?<v>"h��,+�An??�>'��!q
?�T:=(J�9�<�U��_��3��a�J��>-E׽� :�tM��mf�yj
?�/?�����̾�>׽���KPf=���?u?�-)�αO��t�Y[Q��[�]��\��O-����!�y�o�s���a����?a+����;�1?e#�?��~������Mbk��p6��߂>R"�>${�>L�>��8>5m���K8��4e���2� ���>jnx?��>�B?|�I?jc?}�??�u�>��]>���]��>�Ϯ�7k�>D��>��O?��%?��F? *?��?ʠ�=7���+��inþ�w�>�8?��&?���>u��>�B��0}+�����M��=c�O�5���_�=���=�跽�rȽ��=�aH>FR?����8�N���5�j>�d7?�>���>J؏������<<��>�
?iE�>� �o�r�nx��'�>׭�?j8�G>=��)>���=����^��p��=�N���d�=�#���+;��<TL�=��=��h���n�P�:k�;��<�?�s5?G�">��>�T�i�L���\�6>�>��W>�v�>�Y3�rk��yɈ�����cQ�>[��?V=�?��V�>���>_Hھ�#�����b�׾Cf˽��#?
l�>�?&N�?�F?�>7?X�>�-�����W��� ��!?�#,?}�>���O$ʾ֨�Rs3�>s?�q?_�`��o���(��J¾�RӽJs>�t/��)~������D��R�����ۃ�?a��?�.B�YT6����0ǘ�:Y��0[C?¤�>�ȥ>;��>�)��?g�a ��:>���>�%R?֏�>jM?'�}?�^?��M>Y�2�x��쩖�n���>��=?t�{?A��?��v?��>��*>��,�(k�@��SN���ѽ�ρ�%k�=�!r>��>\��>�ɛ>/�=���m-��ǻ7���=ǟO>���>7��>��>5�o>{=Y<�F?J��>�����������4���w�O�n?A'�?�"?%P�<T{%�}pP��| ���>8C�?Z�?`R3?ge����=���;aƾ?
2��D�>��>W�x>h��=�l ={�+>�>%��>.E$��[�L.C��8���?/}B?=T�=$ƿ�Fs�b�w��t��QŽ<$?����d�1����]�6�=�ǖ��v�CF���T��_����������$2���b�>��=U#>מ�=���<6�輻�]<ߢ!=	�$;��3<2L���-�:�:(��������DM�5�<G==�3�p`˾�e}?"I?��+?�C?��y>`�>M�2�n�>/*��Q<?��V>Y<N��!����:�����%��v�ؾE@׾�c�X����2>��H���>)K3>$�=�τ<M��=<�r=ğ�=X	h��=1#�=*[�=�W�=8��=��>
�>{Lw?ޏ��o����:Q����y�:?�i�>���=jeƾ�@?]G>>�=���������3?X��?�d�?�?! i�v>����j�����=6;���<0>
��=k3�r��>�J>_��F0���3��S�?&z@w??F����Ͽ��.>y8>�M>�R�q1��\���b��7Z�$�!?@Z;��J̾��>�=�%߾KPƾ��.=h�6>G�a=���h\�<�=��{�R>=�{j=A�>��C>���=�(��U��=\AH= ��=�O>��56�\�*���3=6��=M	c>t�%>z{�>��?�l0?aPd?�<�>P�m���ξ�Z���T�>�]�=-0�>a��=��B>,~�>C�7? �D?&�K?�i�>���=�޺>���>�,���m��B��맾�6�<���?�ֆ?���>��M<G�A�J��E>��fŽ�a?�41?Yg?�̞>��;ؿ��E�ސ�&¾=ö�=I��c��v���w=�V�|->Ў�=M(>�yt>��=� 	>0 �=�<���>�=/>�?�==\�<��m=�4�=�E�;oO>6��<.<<&�<�GK=��IW<�]����9=X��R�z�rq���>7��>�}>'�>6��<Sԣ���h>'W���NT���=�^���:���e��A���-*��+���`>�Gq>VR���ې����>9ā>�*?>(�?rYg?1>��7�O�̾{9��P�K���J��)�=Q�>bWi��:9�I0a�A[@��a�L�>J��>[�>��m>$�+�J>?��}=�Tᾷ�4����>�ǋ�j:�Q��/�p��M������Ci����qE?&����=�%~?v�I?h��?m��>E���q�ؾF�/>ɖ���U=	��:�n�G���E?Ǻ&?���>�v�7;D�� ��[����X�>���I[������=(���z=�Ծ�ſ>޹�$�Ǿ����b��J���/a����a��>�W?)}�?�塾ژ����A�^(���$=Dt.?�s?D�?�M??�?���<OZӾo[�<Z����R?���?���?���>a�=!���¶�>�S
?/�?ʨ�?G�q?C�B�x��>�);[�%>`�����=�>R�=���=�
?C"	?�
?uԠ���	�n�!���Pw\�N��<��=���>}�>��t>.��=�c=;��=z?`>�؝>���>��_>/��>�ǈ>�Ș�1���G'?C[�=��>�$3?�W>�ף=P�ֽ$ч=G�r�a�X�!4"����[ȽŬ�<���͠<w{�`�>��ſ��?� T>>#�
?��辣K���L>Q#e>/o�>Kd>��Q>���>�՞>X0>�|�>��=>Np׾��>T�x�}B��BD��?R�J �Άv>n�����:���(�T�2��޾���J�|��y��9�\�����?6ʽ��P��w@��f��?��>�S�>�rF?��O�xw�=��=���>�ܩ>�_�V栿W3����۾���?��?Մ�>�U>6�{?�"�>e�v���۾'�J��[���^ھZ�s�	���D���^��&�'�V��-�q?F�q?F�x?T�^�8�u>*׉?Kg��D�=Њ�>�,��G@�$~�>U_�>��"������V����O� �惽9l?�a�?P9?'J�	Ž��U>m.?k�,?!�?��?��\>s����?�6���?�J?�fH?T�3?��6?��m>���������+=0Q��"u�� Խ�Kc�9�=������A=5�\=_k�=&3�<Fn}�$06=��dV+<x�������@(=���=��	:-Ǧ>RQ]?u��>�F�> q7?e����7�/����.?�J6=9��'J�������<���>��j?�ݫ?VZ?�Mc>��A��B�9>HD�>�J&>9�Z>Yj�>�A��C�=܈=��>��>P��=L�H���P�	�iz��s��<��>6�>�x>dυ��c'>�ѥ�O�s��sf>��T�Ҭ��pV��#F�,1�q�w��Ѿ>��J??��==�mږ��f��A&?ѷ<?3�L?x(�?�j�=�Yؾ8�:�|�H���&���>ps�<����a��l���us9�9M���t>�H�����mo>^`ݾ����[�� _� +���ۼ�>�n+��c��S��탾NL�=���=�eξ��%�޶��Rկ�2pO?�y�=o~���g����%�=Eٝ>4+F>���=f��=�]9�8x��/�<=��>U+>W8⽛D��D:��Z���>8Q?�7P?�u?'�u���J��$W�K�ﾝ`���7���z?z=�>D�?(NL>sߞ;�E�|r<��f}�C0��`�>4�>�*��.�Y�6�׾���797�K-�>hk�>�݀>���>>�c?���>着?Ǹ;?t�?!ժ>�Λ�����&?%5�?�o=2�н�4^�N�7�=�H�da�>��?PH���>4*?��?5,?�4M?^�?7�="���G��B�>���>�+Z����9(p>�C?�V�>:`Y?_�|?�)>9i2�.2��T����=)] >��5?��&?�?�8�>4��>VZ��5L\=���>�&J?qف?7ok?���=�E?�8o>�4�>�?�;Ӽ�>�a�>��"?��Y?Cl?*�J?t��>6A�ghK��t��a��&J<+�5����=S��:������'���Y��F{�<��㼝j��%.�����d�3�q\�C��>��v>�,��:'5> �����3>���Km���v���{3�8��=]��>R ?P�>�&���=ѯ�>ϊ�>�����"?f?�?�&x���^�}�ھTK�"`�>+�A?^��=��i�aǑ�_�w��}f=�]l?�s[?.'X�.vﾲ�]?�bd?��۾�/�Zξg�f�5�	���D?�j�>��B���>rwy?.�n?�	?��W��-i�e'��z&{�B������=���>����h���>�* ?}��>�׈>=�<��Ѿ�k��	����?�i�? I�?Ef�?��s>#�l�.��U������U
^?��>~{��ǧ!?D�Ի�eѾx鋾����%��ի�k���uC��[Z��p�!�A�����׽;��='�?�?s?l�p?��^?IE��%�c��8^��!����V����q�ܻE�	kE�aMC�Яn���RT�ߘ�WF=Ȁ��SA�
v�?�X'?��/����>�ژ��'�Ʌ;s�A>�㟾hg�X��=�؋�E�@=�[=��h���.�Ů�� ?���>(��>Sw<?�)[��0>�Yu1��8�|Y��64>���>��>vu�>�KF:��-��W�Xɾ�ڄ��EԽ,�v>R�c?�ZK?H�n?���=1�����V!��#3�ah��0C>��>��>uCV�{s�E)&��d>��As��%�[D����	�3�z=m2?�f�>Qb�>�M�??��	�r����Sx�/Z1�eD�<M�>��h?~��>8G�>�Ͻh !�倷>�]|?�ȣ>��>�@��S}����"��oͽ
�?1}>�$?���>�;�<.@�4����>����Q�V�>d#�?�|�\h��I�>��E?�r�=�C=>1��=2ֹ�%��k���P��b����>��=A=|>vX��2��"ⅿ)�)?u?�a��7�(��H{>�"?Ui�>N��>���?O��>|ľ&k���?F1]?o}J?�A?$a�>e�'=�w��I(˽+�$�/=U��>X]>�Qh=��=�����`��^��U=�u�=�����P��_�;t��BhD<��=d�1>85ؿ�<��Ǿ��A�辳���崾K����ƾf��;���S8u��K�Ӱɽ�����ZW�Q��	���U��?j��?�w-�讏�+	��t������M~>�D��3:=ZD��iBv�T�Ⱦ�,Ӿ���� Y)�r�H��Kc�-dc�Ԕ'?p���f�ǿ����/:ܾ5  ?B ?.�y?^���"��8�� >"I�<�9��M��Ț����ο������^?;��>��-�����>��>ǣX>�Lq>���C螾�9�<��?�-?.��>ʐr��ɿ���Ф<��?:�@w#A?PD'�Ŗ�U\=��>��?N=>�}+��@�+����>/Þ?�Њ?�q=F�V����d?���;�F�����=j��=i�=����CK>���>� �ݹB�Fֽɜ->Z�>���XX�q�[�e��<u/^>�ӽ
����?n�x��.�zS�������>ڡC?�?D]�>xhi?zwW�nҿ�����\?���?�~�?�O5?mݾ��>��Y�X?�V8?k
�>CB�O$|����4oU��J>���&0��y�>B?��
>������s[��U�>���>�V�.�¿�!#���"�Q�<@c��/��\�սd�ӽ�V����#	T�!�����=-�=DK>TKz>��>>��8>��W?�}n?G��>b��=�dĽNt���Ҿh��d���}\�8勾HRC��E��lg�A�ؾ�s
�m�����_˾N�>��q�=CQ�ʑ���h ��b�T�F���-?��>��о�aM���x<�UǾwm��F��<���(^̾��1�\n�@�?��B?d����V��a�=%�/ ��ќU?0a	��'��Ь�6��=;�缰r=s�>�ʗ=W���2�"S�ɀ*?��"?��Ͼȝ_��Wi>_���bD��]7?�`�>T�<��>� ?Rz����=�;>�e�=Sٜ>,��>G��=\!���8��	!?
�N?�.�E|���n>ZI��M|��g�=�]=ڀD�w�=�>;>��2=aS�����<# ���>GIM?�V�>�0�'�����-4��mf�=�&_?��?� �>�"?%�Q?���<[��Zi�~g��=P=�{?O�f?�,�=�MI��-��ק���n?��e?��N>kmI��,��E�U�����&?�	s?5V?���<	���C��%o
��9?/�v?fv^��t��c����V��K�>]�>���>M�9��r�>`�>?�#�LH��׺��U4��?ڕ@E��?#H<<��S��=�5?L_�>U�O�h9ƾ+���F����bq=I"�>���fv����yF,�*�8?L��?��>w������ߠ�=ٕ��Z�?N�?����)Fg<����l��m���n�<U̫=U��B"����}�7���ƾ�
�I���p޿�ॆ>�Y@>S�k)�>�B8��5��SϿ���\о�Rq��?ā�>�ȽȚ����j��Ou���G�2�H� ����I�>��>RN��g��a�{��p;�8���>ʍ��>��S��������1<�Ւ>ۓ�>x��>»�������ș?�����:ο����m����X?te�?�x�?vk?�><��v�ϥ{��<��G?��s?)Z?�N#�]�z�7��j?�^��\U`�ǎ4�fHE��U>�"3?�B�>�-��|=g>��>~g>�#/�n�Ŀ�ٶ�7���Z��?ԉ�?�o����>p��?~s+?�i��7��f[����*�`+��<A?�2>�����!�:0=�Ғ�w�
?�}0?�{�.�F�_?,�a���p�E�-�L�ƽ�ۡ>�0��e\��H������Xe����Ay�m��?>^�?f�?0��� #�6%?��>򝕾�7Ǿ���<���>�'�>*N>O_��u>���:�fh	>p��?�~�?�i?ݕ������6U>��}?er�>f�x?G�u>8�?&�>�֚�6���{Hv>I�<��<˄?��A?��? �C>�"�>� �!�+�',@��ʾ7K;����>�2w?��p?c��>R�l?��¥%�;X�=��6�T��=�"&�k�	<�i*�"4>"6@>���=�U������?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>B�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��"?�-��Nk�F��2����}=��>��n?���p��>4ʫ>*і=�W�K��NJ��[�>�ڸ?d>�?k#?�n�?j8��<b��y�<�>u'�?��s>�,F>���o�>g�?�?"��@��A�ݾ ��?��@.�@ʯ?������ٿn���3;�^澫�F=���<���=���i{=���=�dv��=I>#��>�L>�,>'>�I>�V>��Ck��ۛ��8����c�j�5��;����+�*�s~E�ّ�{3s���þz׽͡н�=߽��a�!	B�2����=<�U?��N?~�o?�?�����>�&�^��<� �(��=Z܉>��2?�~O?�?'?-�=�̚�v�a��K��z���b��,��>`U>kD�>���>G��>��ֺ��H>-�=>�5�>�z�=��@=�	<)�=9qG>��>��>�н>YF<>M�>cδ��0��y�h�w��$̽� �?�����J��0��Q6��d����|�=(a.?�y>����?п����}1H?O���f*��+��>��0?AdW?I�>�����T�n9>���j�:a>-+ ��wl�~�)�P*Q>gj?ܫf>�u>��3�]8���P�!���AJ|>7(6?q����G9���u���H�jTݾ�UM>�¾>��C��e�u����
��_i�m�{="|:?Kw?�&���갾�u�zY���^R>+=\>d�=�?�=�FM>��c��ƽNH�w'.=Γ�=�^><��>�E>$ ?=�>UQ��$6���>��p>.�/=y�9?@�?1���w�
�����)p�Ǭ�>*��>�%�>�>�]���<3�?�D*>G�˽���hm��憃��_/>*�7������ٽ1_�=q���=B��=�0���K��n�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>B�Ք���b���ts�C�<v�>��D?�S���Q���D�3�
?�?�󾫉���ɿ�w�]c�>�y�?��?%o�p���VO?��4�>7�?�G\?qIu>�bپ�T�VF�>� @?f�Q?xհ>�����$���?f��?��?��G>�_�?H�g?�`�>d/�z��E7��A����a�=.�#��'�>��=Aު��B�x?�������t���,�y>�#\=�ȵ>��ʽ��+�=��ɽ����Cu�8��>��>��,>b�>���>��>P��>�_�=��[���{���C?�?���e�G��wc=��¼�v��f�?���>�A�E:��	�>�LN?;
�?�2?-_>P��)����ȿ����%��Z&=�{�>�/?�j�3Y�>q���a+�Gv>���>�ûY��O�8����l�>�-?��%?J� >̘ ?��#?X�j>(�>�^E��7��]�E����>ߣ�>�E?��~?��?�Ϲ�hY3����O桿�[��CN>K�x?oT?Aʕ>����ׂ���3F�E:I�P��O��?.pg?YA彥?_3�?��??�A?7/f>.�� ؾ�ĭ���>��!?l��^�A�Ӏ%�����?ɸ?���>Ӌ���ս�����/�������?��[?�%?����`�J�¾^�<"M�5����
<��Y��/>v�>�4��R#�=�J>@j�=Dn�@�3���i<ͽ=��>���=��5��!����+?H����$��r5�=(jr�%WC���>��F>�����J^?PE�xx|�1��q��*�I�*@�?]�?%�?0[��`�g��<?�#�?!�?��>N����ھ��v��倾�[�#g�=��>��(��Z�j棿�㩿�񃿎YĽ|��)�>QZ�>mV?� ?�>S>A�>����%�Q��	����^��,�&�7��/��������p#��߼i�� ({�o��>����b�>Bf	?�Me>�	z>$�>�	���J�>�yR>��>b��>��Y>��5>���=�	;P�ٽ�R?3鿾��'�4�羾���]�A?O�c?��>ޏt��D��B�FW?u�?���?��u>�Nh�%�*��*?N'�>=��e�	?�@=4k��Ng<�����y��A�����>�ݽy :��sL��g��G
?�?ω��C̾�н�e��Rԝ=O�?��?$/!���_�4Mx��Z��V��讽z@z��5��>;!�Dba��������I��~�0��pq��/?�s�?����+�����f���,�>8?w��>6Y�>[X<>��}G2�ݪS�.�狾�b�>�:m?B}>��B?Ã_?�&q?�p[?Zu>�Z>Z��L�>c�=���>.��>~�K?@�6?Έ?���>��?�fS>O⏽/��:t��$?R8?,�5?
��>ƪ�>�����W�=C�˽Jw�=,�B��<�cn:=1�*=��a��v��|��=���=�?c�;���.��鸾�)}>�*4?N��>��>��~�����}�>��>�?���>��
0�[�`�>hy|?M!���ȼ�<!>O(�=<��~���=W��}`�<8�<�U��|�/;S
>�T=��z=��P<T?3���/W-����>7-?U(�Wo�>�x��A��tQ��T�Ɋ>��>�h#>���6y�������}����>_��?�B�?2��;��=7��>/����T�s�����EVܼ*�?d ?�d;?�7�?]݂?�$?�>��N�c����yr��2[�O��>� ,?s��>v��M�ʾ���3�^�?�\?M>a�"���9)���¾	�Խn�>Z/��-~�����D�D|����5���p��?���?[;A�M�6�x辯����V��@�C?��>X�>>�>{�)�O�g��"��.;>]��>qR?>JeP?��y?��Z?��Q>I:8��������mQ��Jc>��??�v�?Ҏ?��y?Z��>��>��,��u��p�����p����TM=K�\>��>���>��>���=3̽)����=�ɾ�=֣d>��>Z�>)��>��w><ْ<��D??�>�������j���m�*��m?�ˏ?k)?����1�gD�a}�a��>��?g9�?.�*?�Y�ܣ�=,��䯷��sN����>Eh�>���>|F�="�<��=>��>���>�H���b�8��Bd��N?!TE?v�]=��ϿLb�c�x��׾�8��i���;](��ؾ�����M�|�%>9�� ��������j�`����������D�?�>��=�7=�,̽��n��0K=Sp>���=`���a��tM=��<%�^<�����Y<�@�m�����V�0�ʾ# t?�JO?Ҡ3?��e?={d>r��=�-~�m�>DIӽ?�x�>��������)�q ���8��SP־Ŋܾ,�O�������=&����>��D>��F=m�,=��>"76=�-=�W<g{=��=?�={d�=�>�=Jx
>�\>�[�?0Ś�ê��DFb��/�̭�?��>X�>��Y�w?�k=>8����^ӿ�"�d �?��?l�?݉�>9L���>$Rb�wk7<Ֆ>�3r=�X�=B2�=�)���J�>��r>a��h���y�d��?��@I�C? ���S�ȿ�l�X�V>��W>�V��r����Uch�Dg�I*?�M@��ľ�S�>j�>¾�p�v��<��>F�==�c-��*c�:�[=�]���i#=u*�=xu�>�U>@�=�dc���L=I��=8<:>�,>��<�=�����L��">98�>��~>A��>�?<90?�Nd?b�>a+n�=�ξލ���	�>li�=Iذ>Bă=��A>��>��7?=�D?8�K?���>{�=���>O�>ۿ,�>�m���M���˦�<���?�Æ?.*�>4zV<bjA�?��_l>���ƽ>f?9W1?s?�֞> ~��`ӿ�i���<�f齮������оJ#��a_�JL��1�<��=﩯>�[�>�>i�>�B�=�>�ϯ>�>��=x�=��<�m�=�=��6=�����A���{�j�)�m��8���JD���6=��<�֏<6��A��=��>�>r��>2��=x	��\�/>wۖ���L���=׌��W>B�� d��>~��.�L�5� �B>�PX>�Մ�+(����?XAZ>p�>>|�?�u?��>���~�վ�\����e�jS�~��=��>�[=�
x;�dH`��M� eҾ���>��>�	�>�l>�	,��?�c�w='�r^5���>vt�������2q�#>�������i�1�Ϻr�D?ZD�����=�"~?~�I?.�?܌�>� ����ؾ@0>(M��2=��_#q��v����?K'?w��>�6�D��@��uw
��R�>x`��"u/��ג��@����L�g�z�ڵ�>�;þtK����
��P���\��"ES�S���X��>oAh?*:�?�ᾺVf���H�!�!�c�I>G ?��?�R�>i**?�?U�ݽ�K۾���+�X>=�?���?�t�??�V>8?�=#���;��>�+	?9��?s��?�:s?�d>���>��;��!>C���a�=�:>ꈜ=tG�=5_?Ku
?ܮ
?w̝���	�8c������^�Y��<�+�=:V�>��>K�r>(i�=�oe=:g�='�[>bޞ>{ҏ>O�d>r�>�ԉ>,��~�	�$?�\�=�s�>�0? w|>��=-�ƽa:�<�0�`;��� ����޽�՛<���\�M=��s��>]�ƿ�3�?W�V>9���(?4�����2�+R>KYZ>���h��>m�G>7�o>sm�>���>}0>�2�>&�2>ž⾻4>�H��nI>�#�'��y�~ڲ���w��D���>h�Bq��|	���������z�Z	���9�.���T�?�l���IG�5�>=9��?�e$?�v(?^ԽV�=L��=+��>#��>��c�������Zs���ʗ?�}�?5l>�^>��L?8�?�Q��I0b����!��5[0�F]���v�������z���&�Zܖ�(�~?I�t?5n5?��<�>V��?2J�����>�#��,�:�=��X>?�X��s���˾z�~������i?o�?��?����OF�x�~>�.t?5{?�v�?<�?�M�>*�ý	�N?�[�;�s%?m5$?8KQ?��3?�B�>/(>/�;��;���ὼ���bU�5����+м�=>�_�;Ѵ�=Y�������*9B=f�����x�כ=�ۼ�,a=z =wƦ>�L]?�>2�>��7?�O��68�T����/?)�;=|傾"C��{���-��>�k?��?$VZ?�c>�B���B��?>�_�>U�&>ќ[>>���bF�gʈ=`�>�>IC�= %O��ȁ��	�y��7��<��>���>/s�<��=8N>=��Z3�4�>��3V������ugQ�����NtS>Jyh?�MC?��=0���5�<��FU�\P?-.?d.?JJ�?2g�;�����=��/�]v��]�>�9=��ؾ/Y��P��������<�>~;ھ��s>����;`j�U4F���辸��=�N
��J=����;�b��!>���=l|���#��L��������H?�vл�)���i[�D-��4 >�h�>H/�>*���qX��=��䠾���=*��>DL>��<s�ؾ[?�v_�t2�>(l]?��L?d�o?I��ZPY�(/?��̣��}��^Ն�:�7?��i>ߜ�>�2>*N�S��n�5�փ��TU��!?lP�>�F�JQ)��6���Ҿ������>ʊ?k��>���>��T?9O?/�?�7?i� ?$�>BV	��\6�<A&?���?�K�=�cԽٶT���8�$F��*�>�q)?ĬB��ߗ>�?D�?6�&?;hQ?�?ّ>C� �jm@����>��>ſW�IZ���`>��J?���>�7Y?hЃ?��=>�}5��Ţ�P���^��=:=>h�2?M7#??�?�y�>g��>ԉ�� ��=�P�>�}e?�?��m?�g�=�?#Q#>nu�>HK�=J��>���>��?�tL?�*s?��H?��>]�<���)L��u�q��G���,;�g<�=�u��vPf�����<�k�;(tӼs���ü��C�)����<e�>Z8s>"ߑ���8>v�¾U^��`O<>{p��<1���Ɖ�O�1��ޭ=!�}>�? u�>�9 �)��=>.�>���>~�Ag(?(�?�?f};\�_�ݾ �Z��Ω>�>?���=0!n�����Tv��p=Yl?�^?wVC��쾓�`?_?�ݾ��,���Ⱦ,�m�[���V?�?V\7� ��>|�q?��l?5�?p�'�g�Oӛ�ŵn��n��^��=b�Z>K�� �\���>�y2?��>V�>6��=0�˾2s�tҏ��C?�Y�?���?��?1lH>��c��޿/e�T��*�[?4�>�I��a�?�,��hӾy񎾘^��K�ھb��D����T�������s�`���	ǽ���=˒?�rt?��o?��`?�G���m\�^(a�m��Z Y����Q�m�I��D���F�O�m��F�$��2�}�t�=~��FA�~��?��'?>�/�"��>� �����K;�}B>E���9��f�=�����?=�\=�g�� .�bc����?/>�>���>4�<?tf[���=�׬1�^�7�d,����2>Bb�>��>�!�>F:U�,�bN�D�Ⱦn�d`Ͻ$�]>��h?~I?^�j?���x3�'�z��c��0P�� ��p;[>X7�=cRt>eۃ��wY�2y2���M��vt����'����~�%c�=y�,?�ȟ>+��>�?b�	?�W�g���/�F��5>�����O�>� j??��>�#�>��ot%�'̊>�	�?�N�>�v>����/�I�wYA�����F+�>���>��?Ԟ�>P"��8�m��ԟ������b)=�Q�?-gy��yw�[��>O�H?��">���=�r>�#�����J� ���h;�=^�>��=�Y>-���t���,��+�u�w&?w�?#H���1!���K>�K?�< ?>�d�?��>f׾�Gz��	?�oY?�N?-`C?�!�>��<+䯽k�ݽR0���=�ފ>��c>��k=�a�=��I��eb�5g��=b=�2�=���'Tǽ�䁺-�ڼ)�w<�=Y�>��濨�;��ɐ�j%�p�վ�����������3�<ှ����,����O��~��S&��JN�m�]�����)[��zo�?��?��?�F>��j٠�ȿ��|Q��5V�>_ڛ����9��u�ʽ����}d��2��j�4�įM�8\L���N�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾}1�<��?7�-?��>Ǝr�1�ɿc���u¤<���?0�@�~A?��(����h�Z=G��>�a	?�
?>�g0��"�y���P��>���?/͊?[S=��W�7���e?���;�MG����=+�=��=u2��J>��>Y/���A���ܽ73>A�>lM%������]����<#�^>Cн�=�����?ed��ߖ��D�������=��v?��>c�>��*?Ŧ����пt΅��Yx?�:�?_b�?��	?Hξ.��>^����M?B)?OJ�>j�>�`7t�"!�=�=�=�I>�F���B\�H��=p�&?J��=�������Ϫ�J8[�d(�=�U��`Ŀ���'�%�x}G=�����3���;1���F�� ࠾�m���Ͻ��,=
�=��R>�y>g(>�6>hW?	lp?q��>�>�������۾�_K�LЕ�1?�ܧ����,�j9��pؾ�OѾ ���M�>���Ⱦ"=�/�=�4R������ �q�b���F���.?�n$>��ʾ��M���-<�oʾK����ㄼ�楽�.̾^�1�f"n�}͟?}�A? ���c�V�����j�y����W?"N����鬾?��=�����=P"�>�z�=���  3��|S�}�0?��?_����ގ��c)>
�����=I@+?�� ?-�X<?��>7B$?�Z*�Љܽ@Z>��3>E\�>*�>?>�쮾�!սŨ?�U?�^ ��ڛ����>�4����}�g�W=Q>�9�`l���U>W͘<L׋����v��w� =��L?��>�,��*�N�����ս�&�=�Mh?4?n��>�9k?FC<?�=�3��\�r����;��Z?�~s?�u>��|��ɾ�j���(?��W?�Z>�j�Ubʾ��/�2���-!?8o??�W�rW~�Q��?��Q??��v?s^�s�����n�V��=�>\�>��>��9�l�>	�>?�#��G������`Y4�$Þ?��@y��?V�;<��曎=;?�\�>~�O��>ƾU{�������q=�"�>댧�wev����Q,���8?蠃?~��>W���é���=�ٕ��Z�?l�?B���GBg<G���l��n���|�<�ͫ=j�kF"����7�,�ƾ��
�����ῼ���>4Z@U�*�>}C8�!6�TϿ��E\оMSq�b�?���>��Ƚ⛣�X�j�sPu��G���H�m����[�>��>�U���ۑ��{��f;��5���8�>���>6ZS�k���v���;<*Β>���>��>L���;����?c����1οͤ������X?�e�?Pk�?�q?Ȣ:<��v��^{���2G?ăs?�Z?>Q$�!]�ش8��j?)_��qU`��4�HE�:U>�"3?�B�>+�-�1�|= >���>6g>�#/�z�Ŀ�ٶ�����J��?��?�o����>r��?ys+?�i�8���[����*���+��<A?|2>���F�!�60=�JҒ���
?-~0?�{�\.���_?;�a� �p���-���ƽJ��>W|0��4\�h	���b�Xe������y�u�?�^�?��?���.#��.%?)ԯ>����ǾH��<�R�>��>�PN>�\_���u>���;�K	>���?��?�i?H���(���B3>�}?�u�>�'�?���=z��>���=�ܭ�u\i��!%>��=K�:� 
?��I?���>8^�=� :���+�{C�XQ�j��TA�|��>��`?�N?�d>����lN[��j%�g�轤�7���*��S��HO�����4>�?>K�">�9$��ɾ���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�(
?��'��0������S��@)�e��>�R?��˾�j?X�>c1��\��Ǭ��S�՚>�]�?��?V�>\W�?EG{��g����>{��>���?�?�݂>�E���>yQ?���1P��n����?�H@��@ �?u��V^� ��KȾ�M�m9>&�<���=)Y��?k>ƒ�<Ն���ĕ9�l>�%�>�}�=� A>t�U>���=��c=���?�!�@J���$��א`�q���_	���h���,Zc��&�nȭ�~��æ��ͮ���������E�Sb��c>:B?[�a?�x?���>賈���7�r��=�C��C^����='��>O3&?	�K?�L?"!�=N���u1]��p�������{s�.%�>�U>)��>⇷>MPX>�c����=�W>�[~>���=&H���μ��<�(>��>���>-��>�E<>��>�δ�@1���h��
w��̽a�?뀝���J�1��49������r�=�a.?�{>���&?п����q2H?F����(�E�+��>^�0?�cW?y�>���T��8>���ɦj��b>V) ��{l���)��%Q>�k?>�j>��Y>�K4���$�**\�{���&�>+{N?V8��E)�Ӂ�XbH�0�ܾ$�F>��><�[=~��f����5n��"~�>�&=m�@??�?"b���Q��:B%�O���VZ>�W>X�==�1'>�*S>�Y��c* ��O���-=l��=�%>m?�|2>�S�=��>����;�>���>s`%>n�>f56?|�$?��{��얽Sae���(���z>V��>�˂>���=%[Q�&�=��>���>��μb�M��E3�.�n���">�d��+Jv��z���r�=��̽M>
ը=yڴ�C_��Hb�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�f�>x�Z�������u�<�#=��>�7H?�W��V�O��>��v
?�?+`�ԩ����ȿ�|v�	��>>�?���?��m��A��>@����>��?YhY?�pi>�f۾�[Z�W��>κ@?�R?��>�9�)�'���?2߶?ׯ�?��,>q�?��l?|�>��u���+��Y��������;�2�����>[��=�{ƾ|L�ԓ��M��7z�Y/$�|[�>Ng�=�ά>�s�`����\>��@�\����H���>1�>�,�>U��>��>��>Gؿ>xj�=����p��fȾ&�O?P��?6���N�g�<���=@T��@?Ս&?~�;d(���(�>�mP?:'�?�2D?�,�>n�
��}����ʿ���\I[� oJ>X��>Q��>����>>����4M���u>Gh>i:��!�ܾ	7���j<d�>|5'?�U?oHC>� ?ħ&?��`>?Ʈ>��F�����sC��/�>%4�>LT?��~?�?wﶾv�4��k��~��PO[��W>�Iz?��?x��>ޖ��ʜ�1��*uS�,儽�A�?�ag?�����?�*�?~�@?F�A?�<\>L���:ᾖĽ\��>\�%?���:4�֭���i^?��>��>B�����Ž�~�<=��xo��"?o�P?�?��_�k�R��2=�|�E�6�S��;%��<cv(>�*>���_C�=�n>�*�=��\���=��<V�=�#�>`C	> {�a/�(=,?,�G��ۃ���=��r�4xD���>JL>�����^?m=��{�����x���U�� �?��?Qk�?��2�h��$=?�?j	?M"�>�J���}޾۔�$Pw��}x�rw���>���>��l���C���ə���F����Ž�) �ڈ?��>U?#��>��<>pB�>w�����'�Ԧ������\]�"��Ǡ:��	2��H ������;���˻�V��Ley��>�ʏ���>�?@�a>�b�>X�>m�Һ���>E�7>�|>D�>�r>��?>0>��лRf	�LR?d�����'���ֱ��q2B?Xpd?�0�>�i�������B?Ѕ�?s�?�:v>�}h��++�m?�8�>&��Kq
?Ea:=����E�<eT��)���D��'���>�M׽�!:�FM�sf�j
?D/?�獼��̾�$׽������=��?,?)�(��']���p���]�L\�h���3m��6��;� ��g��k������Ȃ�v�*��b2;8L2?�~�?@���t+���{��p+m���5�' w>��>��>�չ>��M>&��ˎ5���_�=�3��砾rl�> +{?o��>��5?�Z?�#{?�:-?�S�>-�=��پK�1>"���ۦ>I�>S�1?)	$?ݛ?&�
?,�&?Cɋ>�)ϼz��ͭ�p�?��? �?��>ݬ�>7�z��-Ƚ�J�'O!�E�f>�v=�I=v���������<8�>�O?/��s�8�I����8k>��7?�y�>E��>����=����<V$�>ż
?�M�>�����sr��W��P�>���?�����=<�)>���=Yv����Ϻ9`�=�¼+��= \��-�;���<�n�=,Ք=~t�d���F��:?�;l��<D�>R�S?E�>�i�>������8��Ѵ�=3s�>�Ƈ=��2�~��䣿�g�jsx=�~?�#�?Y�\=�%�=r��>%$�*����E5�r��W_>�I�>�b2?@0q?Į?�\?K�@?;�J>�D����Z��4�Ծ��+?�!,?���>���y�ʾ����3��?�[?�8a�#���9)���¾�Խ-�>+Y/��+~�����D��U����Bv�� ��?쿝?�
A���6��w�X����]��}�C?��>�S�>0�>6�)��g��#�7;>���>�R?Df�>�;?�:�?��r?,j�>���߷�Rܚ���<��"=�16?��t?	�?o|l?�\�>�">!I���Y���̾5�j���+�ͫ�;����>5��>�V�>&�>ډ>Gd��zQ=�D
=>�	 >�S�>�!�>��>���>���<`�G?*&�>Q�������?�������^/�Ov?(��?�?+?:=e��b�E��������>2c�?���?]s)?��R���=Xݼ�:��ݔo�32�>��>�ә>�L�=�vF=�N>���>��>Q��P�L8�l'O���?۷E?��=��ƿ��q��#p�����̗�<�x���=g��B����]�o��=�Ҙ������� *\��ܟ�Ng��ɘ��_ڝ�1N}�a��>xu�=��>~J�=�I�<L��Z�<�}9=��K<�z�<�z���G<�^8�K^���7��Yk��[<}K=q��m��ss?U�U?d8?H3B?r�i>���=����P�n>۴ �h�?��_>�%�������4�=N��2����վ{�Ծ�Cb��b��n�
>T�^��q5>��>a6�=l5��EȞ=��=��=m�;�G�Mp�=���=�f�=���=�>V�>W��?|��t����X�s0
��Qs?Z��>�p�>M�E��||?h*>4/����տ�c�:͇?Y��?f��?���>��[���>Z����e	���a>�R>�?7>���;�
��봵>����u��!���־f��?�7@b�X?����~�̿��=�;>	�>~qQ�C0���\�L�a��Z���"?�s:��6˾I߇>�!�=l�ݾYR¾�+=?6>uMW=�$�
t^�֚=L����;=�m=��>��D>�D�=�.����=�I=��=��N>Ǧɻ҈;��O$��_<=K�=]�e>�_(>��>�p?��6?}ia?J��>�M8�����^Ⱦ�kJ>�,Z=���>��B>���>��>�k?��6?УD?;��>JT=i��>��>A�=�jv����վ�h��4�.>���?,��?*��>���<E�$�M��P�5��@ý/?5�'?���>ڛ9>W���^T&��.��g����*=�r��U��Y���s����w�=\f�>}��>��>�Ey>O�9>C�N>�%�>��>�?�<�|�=S����ܴ<����o�=�ɒ�E�<@Ƽ�p���&���+��P��:��;^��;
�]<r(�;Y��=u��>�@>��>J��=���I?/>����8�L���=qF��,B�J3d�vH~��/�FV6���B>�:X>Cw���3���?��Y>/m?>E��?�@u?��>��M�վ�Q���De�+SS��ϸ=%�>��<�z;�=Z`�+�M��{ҾC��>5��>�[�>�[n>�>,���?��n=S��D�3��v�>mb��4(�����q��y��9h���<k�����r�E?�x��#�=~�}?�KI?��?zY�>Ǹ��ԂԾg&>���=�[�d�t�0'��4?��&?���>�&�G�D��d�V��o�>��þ�L�  ��w���ؽ�f�����>g޽��XӾ<��玿�󎿎�\��������>�"^?�ٲ?����
��$�0�����Ӛ=@�9?�u?�+�>\�6?���>��c�;�Ͼ�]�����=��z?��?��?[�/>ڌ�=Ct��(m�>hq?0ߖ??n�?T�l?I�<�b�>(����*>F�B�m*�=��>/��=W�=3�?R
?�?P�����X�����5s^���=�'�=mi�>�>��w>/��=���=�=@W>��>�>v{f>��>]}>�C���v�q�&?���=X��>d/2?c[�>�Z=@N�����<I�t0?��+�z��~"�5 �<fr����O=�lм �>9�ǿ�-�?��S>���!?�9��$�0���S>�0U>��޽���>^�E>JK}>�u�>3*�>�g>�t�>�(>�	��&>>y����L���?���v��~�8�=J3�P�-�2��s��
�<��0о���vy��牿Z�@�0�y<�֒?>�W��c�%�#�g�-��p�>���>j�.?I�a��1.>˷�=q�>Ф�>˲#��͗��{���h��b�? ��?�:>%�>�F?�n
?�/�m���M���x���D�*E��d����X����7�Sh�
�T?��\?8@q?8�=QE_>�5�?3@��ҙ�M>>Te�4�<���>�^>󶉾Fw������5}��X� ?0?�.�?m�9?�or��u���2;0�>>+?F.�?�#h?��>�.5>�o�>�é��$?|y?�%`?p�$?���=���=
|�>���=z����$�<0��(�w�&U-�9�(=���<���=Q�=`E�<�U<z�@<P^ɽz�\�;�ѽ*���ż�������딃=���>��\?c@�>���>+K7?�[���9�4Ӱ��+,?@o)=j����������ﾅO>Sj?�c�?"�Y?��d>lC��kB��>�n�>rj)>�/\>|��>�𽠮E��ـ=Ƈ>H�>w�=5�N�4ှ����������<�~">wX�>�,= �t�>�.>�vǾ���&�>�_��ٷi����#`�!�Ṡ���n>��h?��/?8�;9ľp����D?���?SgJ?Ii�>{�?Or=�-��Jw��M���0� �>f>��!��2������$�?<��>�78�����Db>{��+۾>(n��%J���辇^=O��i4J=��
�־��|��8�=o�>�����H!������C��D�I?�l=&����BW�-���>4��>?�>&9��_m���@����_`�=���>�-8>�Ԥ�?��zG������>�)E?P-_?�s�?�F��	s�`�B�����7���Joμ��?��>As?dA>��=����3���d���F��2�>���>v���G�������$��Ê>}?� >J?h�R?H)?D;`?�)?��?5-�>?���bշ��A&?-��?�=��Խ.�T�� 9�PF����>^�)?>�B�Թ�>9�?�?��&?�Q?��?�>� ��C@�֔�>�Y�>��W��b����_>��J?Ϛ�>n=Y?�ԃ?��=>e�5��颾uթ��U�=A>o�2?�5#?-�?2��>��>1������=g��>�c?�/�?��o?X��=j�?=2>6��>6�=.��>ψ�>�?pYO?t�s?��J?��>N��<�5���=��SFs�(4P����;�+H<��y=1���4t�(W���<���;X��><�������D�g퐼Κ�;g��>�t>	����@3>\ľ`���I�?>y3��0�>�����;�l��=\�>D�?jޔ>�+#�W�=|�>��>����2(?bk?�?$/3;�=b�9<۾R�L�P��>>�A?��=��l�Ɔ���v��Ik=)sm?��]?��W�����h?Ť_?�����P��Ǿ��X>f����g_?��>���/N�>8/?�>�?�?�ɾ��e��-���ks���^�W�x=�-�>�+'��f�Z�>��%?��>���7M>  �Hv7��ܾ�{>|w�?-1�?��|?O�>ߌ��WܿO�D����qUh?��>\��?VMk��"����۾�þpM�&N��Pз� /���|��cdl�Y{m�_逽i4:>�30?��x?�{?hX?[+�V+���A�R�J��t���b�v*S���d��+�[�a��/z�Ar$����q�+rN>���}+A�Z�?d�'?�0�ٹ�>I9��A��Sh;ioA>0ǟ�߲��j�=�C��A'<=��T=��h���-����U�?fl�>./�>�V<?��[��=��P1��h7�7���R4>ζ�>v�>O��>�����.����Kʾ���#ν�*O>�(\?mA4?Om?�����I��2~��0����X'����>��>�C>�[t�,F��?,��C8���\���	�^����O� ��=�9?�ry>!�>EN�?�V?%�^����
L�A�N��>�Q�>�%r?��>��/>�9V�-8-�ML�>��c?��x>�b�>9x���V����
J�<A8�>c>�+
?t��>a��}+M�����y��Z!%���=�l?��U�H?���ޏ>G�0?8X��+�L1�>�S>�N%������5޼��=aI�>�L���3C>����I� �M�]@�zM)?�Q?����*�u*~>�'"?%��>4�>I*�?o�>�Jþ'��˧?��^?�6J?�@A?�,�>{ =o�����Ƚ�&��=-=c��> [>%}l=40�=���1=\����?<D=�պ=��μâ���s<ﵼ�J<���<�3>�ܿ�1K�·־(%���h�	�$ы�Հ���T���V��õ�����_y�mK�l-*�j>W��fb�LЋ�k�i��.�?	��?�������㙿,!��� �i��>�!|�Un��Rܯ��D�2l���E㾞ʮ���!�IO�X]g�7�c�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾w1�<��?7�-?��>Ŏr�1�ɿc���z¤<���?0�@�|A?��(�>��&V=P��>(�	?�?>�Q1��H�H���HT�>S;�?���?��M=��W���	��~e?L<u�F�F޻% �=<6�=�G=l���J>�T�>V��6SA��Bܽ$�4>�م>F�"�&����^�yf�<[�]>Y�ս�>����?�i���n�4%�ـw�x6+>;Q?�9�><ܢ=~�2?�#A��]ͿG]�zM?"��?�D�?u�1?���l(�>��?PO?�\1?��>uz6���`��=|���~m=��˾֞K�.��=z��>LG>[�2�����`�Z>.;_�Q=8��A�Ŀ6O�s��㸹<�
��c���`������Q���7��l�f�?����8?=��=BlE>�{�>~UT>Z�]>�Y?T(l?�1�>�l>��׽���ܾ)>���V�����΋��m�4�n����������.��u�����f=���=�4R�p����� ���b�ԖF�d�.?�}$>�ʾ��M��o-<rsʾ����H센�إ��)̾��1�� n��˟?R�A?����t�V�C��"e�����A�W?�Q�d���笾���=������=L�>���=��K!3�|S���+?i�?jR���<���x">BC����<��'?e�?�R�<x��>S�"?�@#����`:>�79>x��>��>m��=Vy������z?� X?��˽ݟ��D��>�F��cɅ�o-@=1�>Vl$�$���Sj>T2�;
���';��Z��� =!W?���>��)���9i���6��==�x?+�?�(�>�tk?��B?���<d���S�F��5w=`�W?�i?��>s��5о?{���5?Ȥe?��N>[h����x�.�M�  ?��n?^`?{[���q}�*��a��l6?ԯ�?��������J����=�2�>�*?���>@�;���?!�!?2���8�r�GL��i�����?~z @�i�?}�Y=>Ž�,S=׆�>V�?*������&,��ξ�'>̗>��g�<V[�����G��U�2?đ�?��>�����������=�ו��Y�?��?R�����f<����l�m��%y�<�«=���T"�����7���ƾ��
�����п�٤�>�Y@%Z�F'�>bC8�.5��SϿ���1[оTSq���?��>=�Ƚ�����j��Ou�ĳG���H�S����E�>l�>j����	����{�h;�0����M�>�Z��G�>εS�I��[p��M�0<^��>�[�>̞�>yw��'���Jՙ?,����Bο����Ŧ���X?ck�?�v�?Lj?L�E<?�v�7j{�`���+G?�bs?�Z?�T#���\���7�%�j?�_��yU`��4�sHE��U>�"3?�B�>T�-�g�|=�>���>'g>�#/�x�Ŀ�ٶ�C���U��?��?�o���>o��?ns+?�i�8���[����*���+��<A?�2>���N�!�=0=�LҒ���
?W~0?0{�k.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>dH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?Ѣ�>#D�?4�>S��>A#�=�课�h-<c��=��=��o��>ylJ?��>�� >��ê.�L�G�.TW�W_���E��u~>Xh?s�S?�?>*`��E��O���'�(v.���.������Ҽ�6ƽp�>�%>U�>�M,�������?Wp�9�ؿj��'p'��54?:��>�?��H�t����;_?Hz�>7��+���%��`B�b��?�G�?B�?��׾BS̼>e�>�I�>��Խ����h�����7>0�B?!��D��u�o�h�>���?�@�ծ?ci���&?n�1�T����}���n!������5>�2h?������	?�i�> ꘽��b�����E�a�jH�>�?��?}��>��?Ԓ�qk��X���?a�z?��-?8�;6D޾�Gg=�?��C��i��&,��z$?��@�2@GK<?aߗ�qhֿ����`N��ܗ�����=��=s�2>��ٽ_�=��7=�8��>��5��=K�>}�d>�q>T(O>�a;>�)>���;�!�r��U���?�C�����)�Z�9��Xv�Tz�4��"����@��j3ý@y��'	Q�62&�[=`�{���G�U?x�y?1�1?�.�>"�ټ<�>΢7���<����p�=�� ?�&?v�o?�O?��M���
�[��\Hp��0Ծ@��m�>ԇ>���>��>$Q�>�޹5p�>��L=��J>ԁc>b��/_<$
�<�Ũ>���>��?���>�C<>֑>Fϴ��1��b�h��
w��̽+�?���K�J��1���9��¦��Si�=?b.?�{>���?пc����2H?���t)���+���>r�0?�cW?�>����T�2:>8���j�I`>j+ �ol���)�%Q>gl?ϲh>���>��.��B>��I�<��\��>�e+?�b��`*L��q��C��վ�]>���>H:���R ��d������}�eX=�AB?��?6>�9Կ�g���.Z����(> �J>g�2==�=�wQ>�wq���ʽ>�N���=��=c�c>D�>0�%>L�=f�>8���9v��A�>:y<>��9>'�5?��?S��|��+���R�I�A�q>���>BZ�>i��=��[���=���>�x>C�z:	�n������E���,>G���"l�Mf��ւc=�Z���*�=�?�<���@>2����=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�!�>)�t�F����}�@$}���=�{�>v�m?�����V=eo߽���>Na0?�Ѿ�q���0Ŀ%���吴>�]�?'��?�GJ��T����P�*�>r��?-��?�fh>�����ɽJ��>��'?�Gt?a�*?�1'��"����>�
�?y�}?9z�=���?��.?1��>�A�=�8�.����p��v��=d��d%>�c�=r��<�{#��gp{��sI���߾$��>�=�m�>a����پ!�=AQ���ľY$�=���>͆�=�Ѳ>��>�>��>kL2>�s����T�lV��<�ɽ,
C?ȇ?}\$�����W;>��>�F_>�v�>:v ?2޽��)���v=��2?R	�?�pe?k�=�o�.�����(0�l���\�>r��>���>Ϧ��`T�<<���rH �,�T���'$H>�׾b��/��>kt>P<�><�>*�ֽ�_?Y�!?�hm>��>�H�H�����G����>{ȹ> �?k?/U?q]��_�2�������d���2>�#y?��)?�G�>+��#���L���=�=s6=��?)bM?�h=�?UD�?��O?@�Q?��=3!�~�ܾoF��:<�>�$?*�½E�G��s1�����2?)�?<��>����\�Ƚ�_�<���-���9?�R?�U?����j��Ǿ�?<�>�F�: ;�h(<�7>Wg">�]��oj�=b�>T�=Mg��rd��l=B|!>^~�>e=�=V�@��׽�>&?(U�������L�>�R��,���*>���>-p�=Um?�Z��0�]��,���g��R��;G��?ab�?Er�?W���M�n�f�q?�X�?ȅ�>�22>H�L϶�R���	��2ʾ�{���5>��r>@dH=]�Ҿa�����=�\�W�_���2����>g��>��%?��>T��=�d>�.��������g�?9R������0��v'����p��9�̽Z���H���Tf����>P��^��>�a?(��=e!W>�ߟ>Z"5�ZH>Ŗ�=��>�S>?l>�1�=�Q߼z�����_S?�i��E�*�d��N��o<H?s%g?B��>�����a��������?��?Jm�?f�_>7\g��G-��x�>I2�>v뀾?�}�<�}���<<ѷ�h��-̽P�]��[�>#Ƚ�<;�.PU��K���?��?��;;@ھ�A�*����N=���?#%#?�'+��S9��g�D 7�tGt����5F��.�Ⱦ7��Rs�����k����Fw��Q��vY>�6?Z��?s��'�Ѿ�2����_���@l#>CT�>�B�>�
�>]�>�ָ�u�2�C`�pm����� �>>��?f�>�H?�7:?�Q?qK?㾇>F �>S6��"�>
}�;�>���>�Q7?=�+?{�*?��?=D+?�g>���������
Ӿ�?L�?;1?�R ?'q?4χ��Խ垷�����h{�͘����=��<4P�C҉��k=�\>uY?�w�h�8�*���G�j>��7?���>���>���3*��"�<-��>�
?IT�>9  �9|r�vd��:�>A��?� ���==�)>��=)��9Xغ�d�=�¼T	�=x���h;�m?<�>�=��=`~h���x���:���;_��<��>�o?+ч>���>p꘾�
�f���2�=ϡ�> �@>�[�=��ܾ𔇿���� �a�Y~�>
��?��?�ې; �=Y�>bl��ro����� ���U���_�>r?�;D?o��?�>?�,?��=��$��#��Z������9�?�G%?!��><����	ݾߡ���/��Y?w��>��U�j ;���!���������Qq3>�M��wy�����hM��A������r��?6V�?^�ٽ�/<�F���AÐ�>�Ծ��7?5��>H��>C�>o��7i�
z�N�$><�>�RT?��>!�O?�?{?+�[?�dT>͕8��&���Й�s4���!>�@?ȭ�?��?�y?R}�>~�>��)�l4��]��"R��?�kۂ��AW=�Z>x��>��>�ǩ>���=>Ƚ!�����>���=��b>���>���>U��>PVw>8�<PE?� �>!���|��·������dP�)Kr?Q
�?��(?\��<u��
�E�������>��?ag�?�)?�a�il�=Wo��Ӝ����t��u�>1��>�G�>>E�=�	=�>���>��>�ｼ��/=��h��)?�m??���=%�Ŀo�n��\p�2��(�<�P��E�h��S����Y��˟=������L����,]�J����s������c���w��K�>EÌ=�p�=P.�=H��<�ѽ���<$�3=C�n<�=э����<��P���u���r��n��;	�;=ל:��ʾd�}?�K?B�)?ܣA?��r>�>�f�G��>�����?��]>GA&�����/�HJ��cP���2ݾ��־ҙg��ӟ�X>%d@���>=U1>���=Ƴ*<�r�=��w=�@�=I����$=�`�=U��=���=�l�=%�
>��>=��?,���>�����1�8��<�21?�e�>|v�=e׾5�L?��Q>cg���ݫ�*��~Tm?���?�b�?;�?{G�tq>Ŵ���wؽn�>4�]��r�<��<���3V�>ܡ>�g������d�C��?���?18?J��ɾ��m7>�4>��>�3P��4.��f`�Lj�1�`��N ?��7�gʾǃ>H��=:�ܾ&uǾ��=E9>�w=���\����= Dm�AF4=7 =��>�ZG>O��=�:��u��=<�I=*��=�HU>ɇ/<�(�u	Y���<�X�=��^>-�+>�a�>O�?}C0?�jd?
?�>�Pn�=+ϾL\���D�>��=�>�_�=��A>H^�>��7?��D?;�K?ד�>�߉=��>s �>d�,�(�m��T�r���sB�<�{�?O��?K��>D�N<#�A����v>���Ľ�Z?$1?�H?��>�U����9Y&���.�$���|4��+=�mr��QU�M���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=$�����<�vż�����u&�:�+�1�����;r��;B�]<_��;#	�=w��>ψ><I�>쮤=3�¾��>�ԓ���@�dɮ=Hu��-	:���]��u�Ί2�u�-��cR>�6g>c.��&���q?~MC>�Y>C��?�&l?Z>�� ��=޾b���;j�@#`�@��=�:�=��*�X=�"�_���C�Д��ڳ�>��>E�>�m>�,��B?��v=����W5����>d;��i\�b���.q�[7��j�3i��/Ǻ��D?�:��c��=~?ٷI?�Տ?k��>����\ؾ�/>�A���K=9��Op�x'��{?%�&?�H�>���T�D�)����&����>�Q}���V�x���#���<Q�$��>�W��ϋ�*T	���������FH�ä�����>�?n?���?z5����swv������	�z�>~ل?��?*ʁ?=H?��2�B ﾲv��R�>>�^?	��?ؙ�?b
�`�=������>kN	?��?SN�?|�r?�5B����>K�j���>EΎ��=�N>�Υ=���=??l�	?!`
?oG���l
��]𾘤��n\����<�d�=䕒>B��>Or>*��=�d=!*�=�X>dG�>�S�>�e>��>}C�>�b��%M�j�&?=�=_��>4�1?���>�]=̑��<��<R�D�+�?��L+�.總b὞�<vp���sQ=�Ѽ��>�qǿ�'�?g$T>��,?�G��9.��R>�~T>�߽	�>i�G>�|>݌�>9̣>K{>(�>_b(>Usʾ�� >���������?��-T���»�>����SA9�(�����������þ��m�O���pX1�L�T=mݍ?�N���sX�{�7�/�7�>�?��>��7?����|nG=��=˂�>)�>'\ᾧ������������w?U@�?�4T>���>dpO?'{?�$��VE��X��Xt��v8�ֳ]�1hd������U���2
��PӽFZ?�u?�G@?�L�<��k>0�~?QE$��
���[�>H�*��=�8��<H>�>҄��K8d�s\־�w;i�3��?>��e?� {?�l?Z8��6Ⱦ��=)�^?T?	�?�?>�?�f���]b?��`�Z�8?
��?jA??�%e?��O?7{>V��O��"�7=.��/�m�p��O��ۆ�= �b�'��y�=v��=As>��B3��W<=">��L����Du<:XV>.^H>��=�h>@b=?UZ�>g�>[�?j���04�)��6)?|�%=�&��ܚq������DE��orO?e'�?�F?4��=#䀾0l�KyL=��>�~�>�%=>�`>r:��ؠ���<��>�>>l�<���9R��A%�K^��A�9=�T�>d��>��x>��x�zR">�����D��"�_>+�R��G���R��II��/�e~��X�>�H?+?
�=Ox㾉�̽��d���(?8�:?b?I?�Z{?B�=8޾z6��AK�-�"�`l�>Mq�<�]�[����c��o�9��x�	rb>O���o���k`>�>�IZ޾�nn� J���羏�M=�6�"Q=�|�S�վ4c���=�	>$M���� �U����ʪ�Y�I?�&k=W�����T�-a��0>!
�>�)�>�3;� �u�7@�5����4�=���>��8>΂��Eg�*=G�y���$�>�yE?a�_?�q�?~.��*}r���B����ή���ټ|�?H'�>�?uiC>���=ɚ��70�3�d�ԔF���>S�>u)�b�G�>㟾ʹ�}�$����>��?�">C?R?��
?��_?@�)?5�?/;�>��"���@&?x��?��=�Խ��T�F�8��*F�?�>Ji)?�B�֗>�o?ͪ?��&?�nQ?��?��>�� �N0@�5��>�Y�>��W�(c��E�_>��J?ϕ�>�BY?(ԃ?�)>>�y5����������=��>��2?�>#?ک?���>k��>ޭ����=���>�c?�0�?��o?��=Y�?t:2>5��>���=���>i��>�?.XO?�s?��J?���>���<q7���8��#Ds���O���;�sH<��y=&��44t��J���<�
�;9f���H��1���D�� ��)��;f��>�w>�Ñ��q9>����m����9>1�����_���� 8�#��=�y>t� ?��>�M*�bq�=F�>��>���=<)?K�?��?Ur��\6b��ܾ��A�+�>��@?F�=мk�Ӕ���u���m=J	l?�O[?��c����D�b?��]?�g�=���þ�b�Љ�W�O?:�
?��G���>��~?/�q?&��>��e�2:n�'��Db�w�j��ж=�r�>+X�T�d�@?�>A�7?�N�>~�b>�%�=?u۾.�w��q��8?m�?�?���?�**>��n�J4�}���7����Y?��>x��m?�<��,�ξ�g����������a������Gr��]���%�ci���6 ���=�?�en?5r?�Z?�9��8b���_�`�v�qmV�:��M��^J��OA���G�L�m�����ﾧ�����j=�lA��:��^�?�?�-��H�>�M���n����4d>%@̾Vm�S��=�/�J�2�V��=��M���7��>ھ,%?�B�>
��>_�2?�T�.Z�����DJ�#�
���)>�ɽ>���>˂�>w'�=���ڼ e����9"��e�`>��z?%_?��n? _��ՒD��q����#���=6k�����=V��=m3i>�:���+��v=�t�N��;��_/��<���|_=��4?�b3>���>u!�?8�B>��۾��g��iɽ�%��>���>�p?`@ ?�[> �=�/:�7�>r!d?���>P��>³޽R@��}^��u���"�> �>�<?b�s>i&��9�` ��v>��c�&���=�sh?R}��t�+����>��R?��=��7=�K>i�1�ռ5��<.����1�"=Խ�>��={	>>��ؾa-,�C�������
)?O?*<���_*��>�'"?w�>�.�>a<�?���>�%þ��P�C�?_?�J? �@?�K�>��=�V����ǽ��&��@+=)9�>oZ>d�m=�(�=Y&�H9]�H ��6G=�2�=5�Ƽ|u��f�<Y���$�P<��<A3>�&ۿ�KK���ؾ���H���	������m��L���M��d������1Mu��B�+�)��:V�#Sd��d���l���?<��?宒�����NR��K�� �����>h�r�Hlr�s���?�+[��{�⾷���!���N���g���d�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@O{A?��(�e�� �V=���>C�	?��?>L1��C�U��UP�>�5�?���?�NM=:�W�e�	��ve?��<f�F�)�߻�8�=�w�=�O=Q��ʘJ>C�>���YA�pܽH�4>:Ӆ><�"�ѧ�Wt^��_�<�e]>��ս�*��x��?2Rt��|\�Am�07���#�=��e?��>0(=_=?�rI��OͿ��-��?l(�?<H�?��G?�����?C����|M?.L?ߦ�>�1��}���#=��=�����y��dS�a^->�Y�>'F�>ҹ�8� �Q����޵��qV�X���Ŀ�W#���"�܀�:���:�喽�� �R=н�m��bs��>��B��Al�<-J�=�8/>�Xf>��8>8 M>��R?B_?g��>��>KĽd�u��IȾ`� ����$�mT��4���o���0����ھTm	�
@�c��ھ[&=�=L-R�󒐿�� �Y�b���F���.?�R$>"�ʾ4�M�_.<�dʾ�ժ�����T ��.̾�1��n�UƟ?�A?�텿��V����Đ� e���W?qa�!��Tլ����=�(���=��>�b�=���J3��zS�DU0?��?�]ž"���m/>u-�sp�<�/?f-�>��m=���>�/?��G� �Ƚ�->7�)>���>bZ�>W�>�y��d��fb!?��V?b_��Г�U��>��ľ*ꄾ8��;0'>�VC�Q�滝�e>��	= ]��$�@��Ͻ���<��V?��>��B��D�$UA����t�=��?�n?�>)?V�?c�:?�X�{xѾO�L�� �8�9>_?y�k?�X�=@mӻuZ��Wz����??!�8?t�m>�ۡ��~�tE8�)���
��>.t?yb)?��u=I߉�В��'.�M4?z�?kn�'����G���O���>��?3@?��=��[�>�t.?Sy�����
��c6�Dx�?S8@�N�?�^	>��7��;2=?D;?�Ȗ�%���Xy���þ��u>9(?a�v鎿���ep���!u?[��?���>�L����G��=�쐾�?g&�?g¥��D<��#�i�=����.<��=�=���D�˪�T�6���ɾ������Hj�Ń>�-@ک޽G
�>sN?����c$ο5܃�|ʾ`k��A?Gɧ>K�ܽ������h��
t��G�ѧK��!����>x�>�ǒ�h��E�{�� ;��b��>����>�zR��޶�o��T� <7��>*��>�n�>h�������j��?8����Bο�Ş�����Y?�ޟ?w�?�"?�`<��r��x�-�軯�G?��r?��Y?,���IX��#+�=�j?`���U`��4�4HE��U>M#3?-C�>��-��|=�>���>0g>�#/�p�ĿHٶ�+���`��?��?=o�o��>\��?�s+?6i�+8��B\��x�*��[+��<A?�2>'���f�!��0=��ђ�o�
?�~0?sz��.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?}2�>K�?��>`�?�FF>���@d2�Z�>'��=����,?�E?m�>�G�=��@��:���C�v#K�~�ݾ��A��E�>CLn?l1:?S�*>����(> ����Y��0ei�D���G��+�8���J<>��>�x%=ZÓ�B�ξ�T6?m;�f8��t����V��ۊ?�B$?c?��'������T�=�wf?�Զ>Y�Ӿ�ֱ�c�g�)
m=q}�?H�?��?��/tʽ]��>	?Kdw=vU�٘���:���=J�?�r��U��JF���>���?N�@(-�?�Kb��?<H��2x�� x�\� ��5��t�=p2A?Y�mH�>��?�Ԣ=�~x�|G����v��f�>A3�?���?���>�Ek?��l���A����<��>�g??�?r�¼C�վ�?>� ?����@���8��n\?��	@�@%^?�|���CֿE^���`���v���M�H��ގ�<�پ��<({�<`n���=֜�>J5�>�>��`>��:>��J=�������+����������g�B�2�$�7���n��"�-T����J,;�};�s����H������R�R[������Z=��j?*�^?Բo?�h$?]JX���&>��H�@:>��P��>���>`M=?�\? N?��ｐj�c�c��r�̠��T�26�>K�=ӫ?|�?x��>k޽��$>�f�=X�u>TO�=ȃս�.��J��>,\�>�zQ>z?M�?zC<>��>Dϴ��1��j�h��
w�x̽.�?����S�J��1���9��Ц���h�=Fb.?	|>���?пe����2H?"���w)��+���>z�0?�cW? �>#��g�T�6:>:����j�)`>�+ �{l���)��%Q>ul?���> �1>�����/���E��b�!R>95?��_�W�-�	�\�h���:3��>Wz=�������;'���v�$��=ZT?�5 ?G�۽�����|s���%��/u>�U<>��C<��=��>z�<�¢n� �t�Ԑ�<:=��6>��?�U>�=T��>�l�8qt��+t>�4�>8t.= 8>?3�5?$_�� ��� ��1D9>���>�.�>�@�=��A���V=+j?-��>ko}=I��'?t��Wm�zI�=}AG�A&Q���1�Rz>J���͠>>�5=;P���=�@-�;�~?���(䈿��e���lD?S+?] �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>�74�0a������ ��>��?#FR?,X#��	�=�hѽp"�>z�'?$W�eV��U߱�0�R��}�>E��?�ر?u�}��M��@b����>�L�?�ї?���>Y�ľ1�k�R�>��a?�([?��7?�/�D����3?x%�?�9�?� l>�{�?�y?V_�>�*�=C7�Js����U�|�=r���T+>h�=V���2�GN}����THi�V�B�y�g>I.c�v��>p�J�F�Ͼ�d��kX�Ms��b����0�>��>^�=ٯ">��>uD�>���>5{�륽Iľ����r�K?���?���2n�P�<?��=�^��&?�I4?!m[�d�Ͼ�ը>�\?l?�[?�c�>E��L>��@迿-~�����<g�K>4�>�H�>�$���FK>��Ծ�4D�Op�>	З>�����?ھ�,���L��JB�>�e!?���>�Ү==� ?�n$?�_d>�ϱ>�=@��|���]J�l��>���>h?�?��?º��>�0��ʒ�����@�U�D=Z>��y?d^?��>*%��*ߝ�;��;WO�&�v����?�Vi?F7��F�?�׊?�E9?k�:?��Q>w��$�Ǿ#������>O�!?��ҹA��M&����}?�P?���>=1��-�ս�Uּ����~��u�?�(\?+A&?���+a�n�¾7�<��"���U���;^�D�a�>3�>�����=�>�ٰ=�Nm��D6�w�f<�h�=��>��=�,7��s���X-?�6Ľ>z]����=�t���H�Fx�>�+i>?{���1=?LS���瀿*���h��P�����?`�?�؈?�;0�̭c�<(B?o��?۲�>�?9�ɾ�]0ܾ����	[�����%�=O�y>{e���8�S3��������ߴ���4潥^�>�=�>��?���>�o�=n��>5�V�����>�#���i�����6��?/�R���MO�e�|����k���>p7��+�>
�?R@>��[>/1�>G�мcͅ>�!7>���>���>M�O>J2I>�C�=Y�*=��Z��JR?
�����'���^���0B?,jd?(,�>�i�������?P��?p�?c5v>]�h��-+��i?�C�>l���s
?w�:=����<�W�����2����D��>�׽f:�SM��xf�Li
?8,?�����̾ <׽�?��T3W<��z?k?(%���E���s���D��\[�d�Ҩ������
3��쁿{Ʌ���x�ރ|��S5��9q=��2?=$�?FQž���D�ľ��^�Ƿ&��	�>i.�>r��>tT�>H@*<m���<�5�P�k�$�Z]N��t�>WPq?�>��I?�4<?�@Q?o�L?=ݍ>��>�ѯ�[P�>��;�k�>�h�>��7?=�.?�F/?l?��)?BRc>\���?���"9ؾ8c?�Z?[?�<?�U ?�υ� ����u¼�����B���y�WPt=)v�<�UԽlw��G�c=�%R>�X?�����8������k>��7?1�>���>��z*��''�<�>��
?�G�>E �W}r�b�cW�>8��?�����=��)>���=vz����Һ W�=n���7�=HJ���s;��U<B��=���=�+t��ڄ�~�:�.�;�w�<�6?�'?!0�;�l�>��9��2� ��q�>C�7>C?=��>���������<b������>G�?��?i[5����=塜=��C�Ծ�lľ�6����=��2?�?t�w?p�?ǣ*?<*?]�>,�����U �xQ���s9?�,?+z�>9��A�ʾ~쨿��3���?a?�$a����aH)���¾Rս[>'[/�~�����D�������x����?���?=�A��6�vk�)���P����C?�>�X�>�8�>��)���g�'�I0;>�{�>cR?
��>��P?��{?%!]?,�_>��6�����	a���5�,�>��??�u?}��?P�x?���>O`>�1�%߾����''�[(󽡤��U?=�^>]�>ok�>mL�>�=q&ǽ�!��L�A���=��Y>�/�>�K�>��>Z��>�=��O?���>��ܾ�7 ��ꋾ�:]��n���?}g?;�P?��p>U* ���b��D��<�=f3�?Э?�<K?C�!�z�4>����/þ�|��W��>���>��>lm齿X�>+k=puU>U�>��B��� ��Z�k��=p?�39?������ȿV(|�E_ž�w��b���������T���_����M@�����pJ>��~Ո�B�1EϾ#�ݾ����/ƾ���>#q@>R�>+b_>&|��X���D={�{="���oS=г;������y��h�н�%�,~c<�LѼQ���0o/=P#ʾ�T}?�I?_�,?:D?x>��>	3�/��>@��j�?}	N>&�V�<����|:�����
;��*�վ��־»b�ǌ��=N>��S���>y�3>���=��<5j�=c�r=�U�=����Z�=l�=���=�ή= y�=��>4�><w�?�ꉿ�R��- A��LD���;?��>@�>򟻾��J?���=����J���3�Cr?r�@/��?��
?ω��%Ӆ>����r�"=@��=��n��44;l�=v\G����>�Ɗ>��$����������ܵ?Y@�D?aB��	4ѿn Y>W]B>�>b�R�d�0�]W��[���e���!?ʯ6��ž>W��=s���o;T�<��A>=�=(����Z�P�=�׉�Cb*=M�d=��>�;>�]�=��ƽ�1�=�&=V�=��T>��/���7����K&=�G�=Q1\>�%>R��>��?�$?R�n?���>H��G�+����!�P�>���>j�a�c�=�	�>J��>��?��B?�� ?q��=_��>)ҵ>P�D��'��/���O���H��[�?�:t?P?�Ȅ=$}�<�A"��%@���L��Q	?��??�&�>]��>�L�l�Կ�M�P�PX����6��REz��н��ӽ]����P�̴\>݇>-1�>�9F>���=]{�=V�>2�>�%>��,=��>�*{=�j�=��L=�'=��5���=����t�=B߼�k;�F���6G���ܼ���=���=uA>��>�>��>t�>�з��T>�t�	�L��'�=q�H�t8�S]\��}`�Y\2��=b�X�C>� f>1���	勿O_�>F�>�U�>��?��m?Ad=h7M�"��Ք��뛒�}���A@�=K� >>a��8���j��DO�47־���>�\�>���>N�v> �(��=�װe=��߾G�4�4�>jf���o�x4���n�nt��������g�����D?k������=��?��H?	��?�M�>6߫�<�־�J.>�~�����<U#�v�����B�?8%?#�>Dtﾗ�C�{
ľ�3��ֆ�>�	R�z�M������6�*?�=iX߾�#�>����,߾L|(�F���M$����:�}�_�鵝>�wN?���?�����}��^�kv"�o�'=þ(?��x?���>]�?�$?�����nѾ�D���g=��[?���?���?f(c>���=4��[�>�		?��?�?��m?oz����>��";�>�n����=)� >˃>�G�=��>$�?g�
?������U�����#R�X�9=�J�=���>�E�> �>Z��=P�=�ߴ=^�p>;l�>8
�>�5a>띣>�>�>0,�����YG)?/]�={��>��-?4t�>�>x=�᝽:�<��p�/wH��S+��2ɽW�뽴��<��h��ED=�m��e�>^�ſAݖ?��U>k�t?[_��F�w<M>�]Q>�ӽ���>��R>F~>;F�>���>}:>���>��->7Lվg>��	�4� �i�C�e�Q��վ��w>W!��t,&�,�������B��������h�KP���>����<�'�?@.��h�q�+��w
�Ͱ?��>��8?x���dE�o�>���>�F�>�J��L��O��`�۾3��?�?]ā>W�>V�[?�G,?aA_�����=��_�P��V1�ކ>��of�8P���Z��h�E~d�y�g?+�r?��@?T0��6>���?MC���y=�\�>�<�����9:�r�o$���eɽ�>�����*O1>Iچ�f�7?�l�?��>?�S#�q�Ľ�w�>��>?�B�>�]�?��K?_l?�i4�Vi�?0-�֗�>L�B?�Re?��?�m�?�	�B��5|��Ԧ=��4;m�
Y����z�o�x�b=���<^"�=��=~�v�Zt�b�N=t">$��=����;�=��>Fml<��9��>k�Z?�[�>���>�4?�����8����
'?��J=$�n�۶������W�I�=��g?;L�?d�]?��L>�;��j?���>v&�>�7+>��R>��>����+�R�z=��>�N>�=(�g�
Xs�;\� ��Lh=�/>�?��=��1�fE>6*�Q��+ǂ>E���
����y�laZ��YA�����zn>eD?r�=?��>�a��d�>�1?�p2?R�?�?N�	��@�Q8������Oa>-�<���ؠ�� G���2W�� -�k�>q
�8̠���a>Y��*z޾E�n��J��l羯M=����'V=v"�9־e����=�e	>������ �����Ҫ��J?a�j=����!U��0��*�>���>���>�8���v��{@��ʬ����=���>]:>����M,�i�G�y>��5�>�YE?5S_?�i�?]��zs�U�B�����ZI���ȼM�?[y�>@b?�B>�*�=�������d��G��>-��>����G��#���*����$�^z�>�;?E�>v�?|�R?e�
?�`?�*?�@?)�>C淽"���A&?/��?��=h�Խ.�T�� 9�KF�{��>��)?ܷB�~��>3�?ν?��&?��Q? �?��>߭ ��C@����>�Y�>��W��b��[�_>~�J?���>v=Y?�ԃ?v�=>=�5��颾�ש��U�=a>z�2?�5#?n�?ǯ�>��>џ���B=���>�Ya?���?p�k?G� >*?\^/>���>���=�~�>��>��?�N?is?�bM?�F�>ͦ}<����G���\~��q��TA;��<��z=K����|K�l��9��<�<�=��6#�m|�==O�!a���Sg<�G�>��s>h���c�1>G�ľ͍��.A>����A����U4:��[�=m(�>K�?7��>�c$���=V�>t��>���t(?1?��?&;;�b���ھw J��s�>p�A?���=S�l�w��r�u�M�f=Y�m?�^?&Y� ���H�b?�]?1h��=���þ��b����Y�O?9�
?�G���>��~?V�q??��>��e�0:n�(��Db���j��ж=ir�>=X�D�d��?�>a�7?�N�>�b>b%�=fu۾�w��q��c?��?�?���?�**>}�n�U4࿠�,���f�`?5��>+��(�?���<��ξ~H��\���"������/���n���̱���'� z�΀����=�?��m?��p?D�Z?����?_�msY��Tu��nN������i�q�D���A�l=�)�k�=F	�����묾��e<}��{C���?�N"?n�6�*��>;���>���о��;>V���@+����=������<˨*=|�d��%����,6?��>�>%??pT[��O7�V�2���;�$�����.>�q�>���>o�>���i��9�����>[~���½��_>T�j?t*H?��o?�ڄ�w�2����B�Z�<`I����6>�K�=��>��0��l����*�X�A��;w�f�h�����M�_=�(?�c�>�z�>�G�?/,�>`/�pL���Bb���6�u�=ۭ�>��V?���>
c�>�W���&�
��>�k?���>�>ᯇ��p ���x�˽F��>!Q�>(G?��t>&)��*Z������ꎿf8�8�=�Ak?�[���W�B��>�/R?�5!;��B<t��>�(��O�$��x��A'�~y	>4F?PV�=ez6>��ƾُ���}��C����'?/C?�W���*�ظ�>��#?�>�Ң>x(�?�̗>i}�����;G?;}_?�oJ?F7@?R��>90=�\���ǽg�'���-=su�>}�\>�[o=L��=Xn���^�!�z�S=���=�ƹ��p���W'<IBü~�F<�-�<h�2>x��(�B������	�9��.�������*�_���M;��������S��y!νx8>�0�0�>rb�/[���D����?y��?ϊM�A]��K����vf����xK ?���#�=^8_�`����A���9�ҾN�� ���!��G;�P�'?�����ǿ󰡿�:ܾ7! ?�A ?7�y?��6�"���8�� >tC�<�,����뾭����ο@�����^?���>��/��p��>᥂>�X>�Hq>����螾t1�<��?7�-?��>r�1�ɿb����¤<���?/�@R�A?��(���쾡�U=$��>^�	?{�?>�.1��@������V�>�6�?��?��L=>�W���	� {e?H<�F�.���S�=Hl�=�;=�~�P�J>�[�>�x�=dA��<ܽ��4>��>S�"�Bi��x^��y�<�O]>��ս�6��4Մ?2{\��f���/��T���T>��T?�*�>:�=��,?]7H�^}Ͽ�\��*a?�0�?���?&�(?%ۿ��ؚ>��ܾ��M?aD6?���>�d&��t���=V7�g�������&V����=X��>o�>��,���ʇO�I��8��=h����¿����b%��,=����0V���9���#���<�Pb��$�5��v�;Q�=���=~>>NW>���=�9]>��a?��~?4�>�S>��M.��K�۾3 =*�����c�P�J!,��ֿ��B��8����m��G� �8ξ�=�@ �=m4R�U����� ���b���F���.?�q$>R�ʾ��M��-<�qʾ6ê����ҥ��'̾�1�� n�@͟?�A?,���i�V� �mJ��u����W?VR�����款��=?챼��= �>��=
�⾡3�q{S��PU?�k�>��������U>7z<d���3?e�?��\>=�
?}v7?�ȥ�N��QcR>��=h;�>/
?�V�>��������?�M(?-�(�4�ݾe�>P�"����݇>_��=G�h�Iy:>��8>�>���٨+��~����d>�o?4�K>h�O�0*���jj�d:<�zU���j?D�?�I�>}v?��9?Z��u��V&����w>s�U?0�]?%~�=�ԟ=Lu���{��TQ?�W?S$�>|x��B�������A,?E�U?��,?�^R�A�g�D0��A��:?�?Ɨz��e������xF��5@�>,�?~�>��0�v��>v�3?&�]��Є����XO�I��?� @P��?B�<�E��A>,=��)?��?�u��!M��s���ԯ�f�->�O�>|�����R�#�EI̾&�<?Eٓ?LS?M���<�^��=ڕ��Z�?U�?�����7g<���l��n���~�<jͫ=��G"�����7���ƾ��
�જ��濼y��>,Z@_S�_*�>>C8�=6��SϿ����[оSq�a�?ۀ�>2�Ƚh���R�j�~Pu�j�G�u�H����ʢ>��>|��������{�>�9�~=�11�>���Ɋ>�MJ�<(������VT;s�>��>���>�n��	Z��b��?�`��U�Ϳ�מ��R��U?��?���?�<"?j�<�@m��$r�e��,�E?In?�W?����bU��fP�xTl?�3����f���4�VF�#�Z>G�7?�\�>�/����=�$>� �>!n>=�-��ſ�ò��A�2��?���?w5��P�>sZ�?��2?L�������~�$��<��@?��>��;n�$�BI��!���?^w6?N����]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�T�>>�?�9�=7�!? Xz>η;��;�G�<CT�=ɝ̼��?�;Q?�g�>�.�Qs���Y�r�`���r�Y�t���Z�ܐ?\U?��(?��>��;�l�0��C;�<>�腾�7˾�����_�����&�2>�pO>Vfg�N~���5�F�(?�K����JK��A���~a?�?BF�>/S-�`�!��=��O?�\�>�Җ�8��g��&�G�$��?���?~?���ҏ�>:�>�!�>����ǠN��X%��ࡽ>a>��F?%RP��
���݅���'>@��?��@� �?�؀�� 	?�2�*W���Z~������6�O[�=��7?8�F{>���>ͪ=�^v�ӳ��o�s����>�A�?rv�?��>դl?Yuo���B��3=��>�hk?)G?��i�
��F�B>�?>������s�bf?��
@�r@!�^?Y좿�hֿ����^N��N������=���=؆2>�ٽ_�=��7=��8�e=�����=p�>��d>#q>@(O>�a;>��)>���O�!�
r��\���O�C�������Z�E��Xv�Wz��3�������?���3ýy���Q�2&�O?`�4�����n?�*?��?4HZ?��/>�a?>c�+����>�Ǿ��>x��>��g?Wz?r�:?9�h��|'�%��3}o�.䳾�j��tHT>��U=�;�=��p>w��>F�,�{��g���Ⱎ>��>x��=�л���=(��=�zF>p��>T��>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?��f>��t>�s3�`8���P�������|>&6?����:9�i�u�m�H��jݾw�L>���>	�E�3b���b�:�i��{=��:?�?�㲽�۰���u�=$��X�R>}-\>ٺ=��=�1M>��b�(4ǽ�)H��-=n��= }^>�?.o$>��=Ч�>�	��0O�A��>�&`>a�>X=?*�"?k�n�lڳ��`���:%���x>C�>En�>z�>��O���=���>�Y`>���8�\�!�f�M�"oD>
����eL�)����_=�]���>�5�=���`B�FCh=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ]=�>�og�N��~y��'X��%Rs>1�?-D?��1�=p�<>t<�ҁ�>��?4��� ��0�Ŀ��^�U��>>��?���?3����c��K�O��� ?�g�?P�?�r+>]����:Ͻލ�>��a?Y?��?��%��Ǿ���>���?*�?^I>V��?#�s?Jm�>�x��Y/�%5�����X�=C1[;d�>�^>'����eF��Փ��h����j�B��h�a>�{$=��>@�A4��IM�=����J����f����>O1q>��I>(O�>�� ?Ff�>G��>v=�c��Uހ�����o�K?���?���2n��Q�<ڠ�=�^��&?�I4?ep[�_�Ͼ�ը>�\?n?�[?d�>E��Q>��G迿-~��,��<��K>&4�>vH�>;%��eFK>��Ծ5D�bp�>З>�����?ھ	-��LS��:B�>�e!?���>�Ү=ř ?v�#?��j>�(�>MaE��9����E����>���>�H?�~?5�?�Թ��Z3�����桿�[�;<N>��x?$V?{ɕ>[���򃝿JoE��CI������?�tg?Q�E?12�?��??Z�A?(f>���Zؾ����W�>��!?���A�'K&���~?�L?E��>�7����ս�ּ���ŀ����?A(\?A&?��(a�c�¾�7�<��"�tV����;LZD���>a�>S���Ս�=�>��= Km�5F6�-g<&n�=,}�>�	�=M.7��h����"?3��;�0��-�=��y��J=�e7�=^0�>��ǾM�K?g���Ju�
���/��|���*��?�Ҭ?��?i�.�Zt���?��?�4�>���>1�L��h������I��)����A	�/
��N�>L���	~��t���֦�VO��;�:`��xu�>
/?���>7��>4�>=��>�!��y
.��aվi��߬f�.����3�!]D�s�Q��K%����rm¾�z^�ۋ�>#��X��>��>�F�=C+6>���>��+��$>]��=��p>�ɲ>��G>0�>۞�=��"m��KR?������'�y��޲��l2B?�qd?)/�>5'i�܉������?��?�r�?k<v>�~h�.,+��n?d?�>/���q
?d:=T��K�<�V������2�������>)E׽�:�[M��mf��i
?o.?P8����̾�D׽Ή���n=�N�?��(?��)���Q���o���W�WS�M���Ah�<p��=�$�V�p�p폿W]���"��f�(�#"*=Ƅ*?[�?������'��c#k��?��if>��>y"�>]ؾ>�dI>��	��1��^�XL'�����RA�>U{?���>��I?��;?�O?��L?O��>�Z�>+Ű�%��>�w;n��>�.�>z9?
C.?��0?_]? �)?Ϧ^>�󽤹��QؾA�?��?"?�#?�?	���N������Qv���x�^₽�%�=���<t�ҽ'�y��T=�U>�H?����Y9�u����Nk>�8?��>4��>�q��:���8�
=0:�>Z�?�'�>c5���p��	���>K3�?�P�
�=��,>1�=�S?�T�#5�=ڸ���̐=�C�Uf4�B�/<T��=N�=`T���BL��1:�;c�<��?d?��<>���>�W����7��@���i>�e�>&��>��� $�t5���l���xs����>k�?!k�?�9�R�d=k��6�)�� ��� f�[d㽻�1?\?�cZ?���?(@?�'?P)>��������@b�b���p�>c!,?=��>G��U�ʾc�Љ3�ٝ?[?�<a���;)���¾R�Խ�>�[/�R/~�s���D�@ͅ�����|����?���?�A��6�hx辢���\����C?l!�>wX�>��>��)�a�g�s%�.;>g��>�R?*��>[�O?g:{?��[?�T>jz8��"���י��/��!>+@?���?{��?�y?���>Uu>�*�j*��Y��\����΂�<wV=��Y>�w�>��>{ک>m�=�ǽ⬰���>��.�=>�b>�Y�>G}�>���>��w>�_�<�s@?���>������������������?R@�?��#?���X2���a�}�%�#j=>!��?Hu�?�RN?����܇>�#�=����ݾE��>�/>��>�����=}�g=C��>�	?9�Ⱦ]�2W7�I�?�,��>�E?�R�cL����s������/`]�.��Z�?�����xo�q��=I����(E�K签`�d��Ϲ�������΍��d�����>Y�j=��>x�=�X�;�뻥u��׏<�%=Q=�͹�Ԛ:��ռ�\�<������;i��<>E|=%ܠ<��̾-�}?��H?+?�!D?�9y>G->�~>��͖>�a��d-?�-X>֌P��	��P4����������پ(־��c�.Q����>��T�%r>��5>���=v�<!s�=��j=&�=�V��g=���=���=���=*��=&s>��>9w?c���i����*Q�����:?q9�>y��=�xƾ!@?R�>>X2��ޑ��Bk�L?���?�T�?��?nXi��M�>p���K��4��=�ܜ��2>]C�=��2�E��>U�J>$��JH������=)�?�@'�??�ދ�m�Ͽ�/>	nY>x��=$U�Ei)��]���>��u�>'?�q0�K�Ⱦv��>�k�=�D��&оd�=W�G>t��=������S�]
�=`N���?=�"f=RZ�>CH[>���=�L���n�=H�Q=��>d�q> ֻ���!�T�=~ �=��d>�5:>���>�j?�$?���?���>�+��4�޾K����:�>"�>��={YL��#>
��>�_(?��`?��]?)?�>��<��>�>-D2���i���������7��	�?��?T1�>��U=~Yƽ�C6��J2������?_%)?[v'?�t>�V�ޡ�{X&�Λ.�����a�d�+=xr��zU��r��Ms�_��Y1�=�q�>U��>��>�Ky>=�9>"�N>�#�>��>���<_��=S������<�V����=����s�<<żR6����(���+�#-��:E�;�`�;�]<-��;���=���>��->�>��&<���&�G>�z���%W����=�0���JA���W���{���+��H"� �P>���>oÊ�!9��V?�H�>ތ>��?,�Z?�1>�ν�}ھN{���>��Qi���D=���=U�ً=��f�?�S�D6��Y�>c�>�ԡ>S%p>"H*��>�j^=;+�t5����>�舾
]���0�o�V��쟿�i���>�E?�M���`�=rK~?(lI?nώ?�Z�>%����־U1>lV����<����s�l����?�&?��>^�sD���Ծ=Ľ�X�>%�N�noQ�R����L/��ػR���~��>���Ծ�1������K����>�dHl�-ӷ>SM?���?J]����3R�@n��b��U?i?��>��?�E?�����$}����=V`i?�e�?�b�?�U>S3�=��z�.��>O�?���?�R�?�r?�H�$�>�P̼vy+>j�4���=\/#>��=���=�?�?�?=᤽TC�Y��D��,�S��{~=V�=q�>C��>!h>y!�=�ot=U��=`h>��>���>y�X>w�>p �>����ϙ��N*?lm�=�3�>�`.?#��>R�M=��ٍ�<e�u��G�19-����x�T{�<F��#O=4��w��>~uſ�m�?�(X>9����?[����a�u�P>e�R>���K}�>�TI>��{>_��>
 �>a#>_�>��*>Ng�Ns�=9)�~.��<S���H��X��⑄>�پV(,��j ��C�qF�嶩��b��j[��q�&�1�� �=���?�,�����(�F�]���4"?j��>�6D?_���;�=U�>�/�>x`�>Q`Ͼ�[��Q���Mؾ��?:�?�vA>tY�=ؾa?�H?���W����a=���o��z+�}�(��ӏ��񔿵�J��)�(����{?V�~?�6?"�ɽ�|>�p�?��M����=q>���peE�z֩=r?�O:�B;e򚾐��C��*�>�ō?G�?`=�>�����þ�n?�6?g#�>�&�?W�T?ry'?���0?ձ��f!�>��=?D:P?�>d?��d?��<��ľ<7��5~)<Q�l���g�4=�XK�U�=(#*>�e�;��<�=Ƀ�<͘��>���>�0>N#}���3=��?=X=*�X�,i�>EM?j��>{`�>��?P ��rN�O���?�=��o�H�ξD����
�>�">u�f?0�?�\?i�Z>'�@�* ?��\�=��>>�>D�>�K�>��N��\���`� kb>��=��=�?�Y�+�#E��Mj�ט�<��p>�H�>9^D>�p��M2>������|�K
v>��_��1̾�\���J��50���n��/�>YD?F�?8�=܊̾�Z�vIi�I�(?��>?�#>?8@�?��I=��ľ�|3�YM�9��J�>�1�<F��a�������->�q��Tt\>}U���a���a>j��?�޾o�n�J�(��A	L=7V��S=V��־#���=��
>�\��� �7	��aȪ��$J?x2k=O���T��Z���>�G�>WѮ>��<�Hlu�oN@��Ӭ��_�=kt�>]b:>�/�����/�G�9��Ć>�YE?Cv_?#I�?g��юr���B�2���ff��6Dּ�??iΫ>ȳ?ԜC>�+�=�ı�WI� �d���F����>�g�>�����G����h���$��-�>��?j�>�_?�R?��?�`?�l*?.F?�@�>ť��H���:&?�}�?�j�=��ҽm*T��9��5F�0j�>(�)?��A���>e?9�?��&?L�Q?�?:>�x �T�?�T��>3 �>v�W�LV���\`>@�J?��>�:Y?Ã?}>>>Z5��`��l>�����=*�>��2?�&#?<�?,��>	��>ʭ����=#��>sc?�0�?��o?A��="�?�82>p��>���=K��>Ƌ�>J?XO?��s?H�J?ё�>���<Y6��8���Ds�y�O�ǂ;7uH<j�y=���B5t�>G�+��<#�;�e���H�������D�#�����;\��>�qu>n�Q&/>f[þ{���ZB>��������|����6�ix�=D�>D?���>ş&��9�=���>lj�>$��I,(?5 ?��?N����b�t�ھ|HL�8ݲ>0v@?���=�l��N����v���^=�m?��\?V�[����$�b?��]?�j�M=��þĶb�̈́�"�O?z�
?H�G���>��~?3�q?h��>E�e��;n����YBb���j��ƶ=�r�>'V���d�5�>��7?�O�>�b>8H�=�w۾C�w��o��Z?�?F �?���?g*>��n��3��^�V���R?|��>P�ʾ�?�Gͽ�Ⱦ)Š�߯���K��[�ʾԙ���Pr�
'��l3�2k����[��e3=�??�o?~�u?
�W?.w�E#I�5rZ��t�P�^�u��~���<�~EH�y�J���~��r����u䉾�
�=�}�W(A�?�&'?T�.����>阾.#�_�̾�C>w����u�=����4=�$`=��f���.�|���-a?۾�>y��>�$=?U�Z��.=���1��7��Y��ڠ4>��>ʑ>EC�>�9;&m,����7UȾ������ʽ#�l>ȹf?:M?��q?2�a(� sy��'��z�<����r)>�P >p��>ē)�ð�=�,��^G��r����s������=�=%?=�d>J�>�f�?�/�>���ܪ��yZ��2*����=��>�Uh?�<�>�4�>�G�]�%��N�>!1m?�`�>�Z�>؎�~#��E~�sŘ�r�>���>h��>)�c>��9�_[\�-���_���4�z�>�xd?b7����e��2�>8X?��<t/�:(�>]z�3k�P���-�b�=pQ
?{n�=2�b>E6Ⱦ����x��ds���(?m;?������*��n~>~�"?��>��>`�?I��>^���jm;�t?HO_?R�J?9�@?�`�>B4=(@��);Ƚ�&��-=��>��Z>Rl=C�=lH�^�\�vm�˦I=rG�=u=��qY����<)⨼P[;<��<�1>�ڿ�L�.�׾�P�����	����k��
�_@�������Dz�(�	����e�P��>d������o���?�G�?]莾�i��
��
�|�Q�H�>q�Y0e�ä����W1�����L�����!�.�N��+h�Hc�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >ZC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾p1�<��?7�-?��>Ďr�1�ɿc���x¤<���?0�@�A?�F(��O���V=��>�B	?h�@>�0�]��Z�����>t�?���?UdX=@;W��U�*�d?�<��E�c��%��=�ǥ=$)=2j�`eI>�>4�L=��@޽�R6>���>0��B��MG^��r�<�rZ>7�׽�n��ք?-�\�=f�ݏ/��Y���@>��T?��>r�=��,?m-H��xϿ�\��`?��?4��?��(?������>�ܾ��M?0J6?��>md&�t�t�9�=�#༸p�����V��y�=?y�>c>�!,����R�O��y���{�=�U���	ſ�@����k�����C� �׽�Žη��oG��V�f���ɞ��Q��="/?>�{_>��\>�S�=,>_1X?Їd?���>�&>�
潁�B�ñ�91�����=Ȑ���v��PX�	�ľ1&�}��8���%�����1=�v��=1/R������� ���b���F��.?Hu$>q˾W�M�EH-<�Yʾ����	������3*̾ݓ1�t!n�aȟ?��A?������V�����T�ro���W?u<����¬�aI�=�ĳ���=�"�>���=q���*3�dsS�e�0?�� ?��ɾ���I>�D��d1=�S(?q�?�<�c�>Q�#?��������W>���=�g�>6��>])5>6���������?2O?�#��6��.��>����;7� ����� >��)� �����!>�v<��]�������%�;m�b?ѭ�>%e�K꾉�V=k����O�i-�?�>B�(?jp?Z\?�CR�w*���p?���-9�=�dV?o9�?C��=U[\�8`��!����e?�-?�>��B%�Q!_��<��K�>�&T?�>?c,`<u���*F���T2���A?B�?O���n��ڊ�����@?!�;?k��>�S2��9�>;�3?ж��Vb�t}���dD���?�7�?��?B�6>��2�k:�=#T?u�#?ϲ���.�p����
�>>w?B=�L��������^N?��?�P�>B ������=�ٕ��Z�?q�?h���^>g<9���l�on����<Ϋ=���F"�����7�x�ƾ��
�󪜾,忼���>=Z@�T�[*�>�C8�G6�TϿ&���[о�Sq�V�?-��>�Ƚ����F�j��Pu�Z�G�?�H�ڥ����>F�>�j����?y�Zj;��Eܼ�#�>��Ӽ���>�cR�����m��E<�d�>j��>b��>b��[H�����?���� �οp�������Y?�W�?��?�?F�<v�n�cWm�K�6�F?�lp?"�Y?�Q�5fV�A6:���j?�٪�ڣ`�F�4�!�D���V>�3?���>3�-�-�y=6�>���>fo>
�.��oĿ����͸���Ѧ?�t�?����O�>W^�?�+?�3�n^�� Ҫ���*����:�	A?�d0>D����!�/>�ɼ��J�?�Z0?��)~�]�_?*�a�M�p���-���ƽ�ۡ>�0��e\��M�����Xe����@y����?M^�?h�?ӵ�� #�g6%?�>e����8Ǿ��<���>�(�>*N>`H_���u>����:�	i	>���?�~�?Rj?���� ����U>�}?��>�p�?���=�?��w>���o)�<���=OV�>j�J�?�?M?�"�>�D�=-XN�;AY�s[w��jn��ء�&,;�'�>�y?QC`?�C>�MQ�,���-��6��Ʌ��K�8�B��c�|9���g=v >?��<��}�()��#.?R�:�#�ۿ����V�{-�?��
?�U?��>�^쐾��a>-�i?c��>��;�0���S��-=Cť?|k�?*?ɽ��ꌽ�+i>5r�>ވ\=k
<��ȹ��8z��B�=��0?T%`��J��k����%>MT�?z=	@�2�?�}a��Y	?;��*v��<�~��R�<�3��d�=��7?����y>���>W�=�!v����a t��q�>!S�?�^�?\�>o�l?4]o�\|B��:=���>�lj?�
?
ꧻN��2qD>�?/�� Ύ�xY�t�e?�@c@ʏ^?l����_ۿ�e�� >ľ%�����g=ym<r�=z�T���q�B��/=bLk= >7+>�"d>VU>��=��U=D�-<�����T&�S ������YX��"=��&�:���ʵ�����s� �Z0���Ɛ�<��	��3Y�&����9�v:���=+�W?�N_?�iI?o�?�E==�X=50���>�X¾�żI��>SO?�g?�x+?�wE���"�[\d��+^�B����x��>�(J���9>é�>&�|>�i��v�=���=���=�M,>-�=��=��q>
��>Y��>᥶>5�>�B<>�>7ϴ��1��p�h�"w�h̽�?e���Z�J��1���9������Oi�=Wb.?'|>���?п^����2H?1���f)���+�M�>m�0?�cW?{�>����T��:>����j�#`>�+ �pl���)��$Q>ql?.,g>�t>p�1��8���O�����ϳ|>��5?+��� M8�}v�%I��ݾX�H>�W�>Z[1�$��s��������i��a�=��:?=:?�կ��o���x�Uڞ��QP>�q[>E'=\�=/O>��g�g�˽��H��'=*��=d^>?Nz>է�=�c�>Ȼ��s&t�Ԇ�>JOJ>n�+>��;?��?�����ҽR���e<�s'�>6��>B/�>_|�=!�S����=�x�>�y^>b�:p���P/�k�M��k>ع��:��lO����=@x����=
�=���Lne���<	�~?�~��.䈿��2P���kD?+?�=|F<��"�_����F����?O�@�l�?�	���V���?HA�?d�����=�|�>8ի>aξL�ٲ?��Ž�¢�˔	�X##��R�?��?��/��ɋ�hl�r0>^%?�ӾU��>���+��M����c��>��#?{uN?%D� �D=��ݼ{d�>R?ZÏ�\˜��IÿB�U�å
?��?��?��������%T����>�/�?�0�?�ԧ>�k
�Cq�L<�>bǀ?�\?՜?�����Q��-V?��?V=?�H>���?ۡs?Ȍ�>�@v�%H/�h%��E���E�=n K;�4�>_j>?���<F��ē�Vd����j�����xa>� $=D�>���A5�����=YT���'��� h�g��>��p>eI>ZK�>�� ?g�>�Ù>��=����������=�K?���?���R2n��Y�<`��=��^�R&?�I4?�x[�9�Ͼ�ը>ݺ\?q?�[?c�>���@>��'迿;~�����<g�K>�3�>`H�>�$���EK>V�Ծ4D�rp�>�ϗ>���@ھ�,���F��IB�>�e!?&��>�Ү=� ?o#?��i>ޏ�>\'D�����FF�I��>I��>$0??~?�?ƺ��3�LY���X���tZ�R�Q>dy?��?�v�>�ۏ��k��8�E�d�8����(Z�?=�f?3�۽�|?���?q�>?�[A?r,b>����:׾톨��`�>�!?u���A��M&�' ��~?�P?��>k1����ս�$ּ��Kx��o?�)\?2?&?B��,,a��¾�)�<9�"��!U����;ٕD���>J�>�����=o
>}ް=�Nm��>6���f<9k�=��>���=I17��{��#0?]Zt��B��O�=��l��(-��> >;��CX?L+���m�[ԕ�͆���S��_�?H��?���?����EX�9VF?W�?��>Y[?��ھ���,�|�c����3��x����=�B>��=�ޕ�3ǝ�ԕ����d������ؽ��>�?[b�>NU�>�L�=.Z�>9���A`��Sʾ�U�L�e����~�D�[�8������
�"��d2�8��.�f�=�>�4N=o��>��?#	�=g^7>�ă>6|"=.�!>>�ϗ>�=�>�eO>�F>c� >_�=v�={R?�z��4�1fҾ�H ���$?�`?G��>x�<&�c�𰭾��?"�?N��?��>��/�/����>�?�����?�h�=�PԽ%���jɾ�.����{��z>�	>}�=<_?��'�U����>�.?�
a��W���[�B���t��<��?��!?F�2���E�1v��T�%Z[��}�x�V�7���(��f�m�����I����U5�� = �2?�?��ݾ����b����[�F�&�9�p> ��>�
�>���>R�=>SK��B;�T�j���2������?E߃?�>mrI?+<?� P?U@L?��>�G�>�Ѱ�٘�>�V�;��>���>��9?>+.?c~0?0-?��*?�>a>U�������oؾv�?rP?b�?f�?@�?�����JĽ�����b�U�x��)}����=�y�<��ս�iu���S="CS>K�$?9�R�b�D�_򾾖�?�"?'�>@��>�6��:����<0�>)�>Z?�>�=Ͼ�����Ti�>�o�?��j�X�<��A>u��=��>����%v>,��-YB>��ͽ��=�&:��ע>|�)>%��=bJ������*	�s���(�>:?b�.>LNB>S���<���&7E�$Ů>X%<+�>��\;��ܾBѩ��"���t���<�>X	�?�t�?��n��ܤ=t��=|'P�RR����(̾�����A?1�?�lh?J��?�1?�'?��=�3Ѿ�B������J�E�?o!,?���>���ճʾ/���3�ٝ?.[?�:a�����:)��¾�Խj�>c[/�q/~����D�᷅����,|�����?���?�"A�b�6�y辥���Z���C?!�>Y�>l�>�)�d�g��$�f-;>1��>�R?,��>�O?�y{?�\Y?��X>��4�����r���<Mc>�;?Ja�?)b�?ӑy?���>
}>�+7�l7�ӫ���F"�Z���􂾥�=U�G>���>�z�>�>-��='ݽn��ܚ-�R{�=��j>���>i�>�m�>�%z>KO�<�DF?���>�¾�þ�?J��~��+x �X`�?-��?�,R?�,�=l��ߚN����.�>���?��?�rA?�Ќ�V_U>g �<��t���/>M��>h@�>޹�=��;�A�>�#?��??�7����]O��`ػ ) ?bA?��=1B̿k<��
������3��8���HV��S�K��P��>���1�(
|�� -�-�d���y�@뭾A�dF�����>��=5�>��=>��4�-cu�A��=sw��ٹ=Q�=��v�ν�)�<1:=����\����̼\B=h����~?>�L?on/?��G?��a>���=�Ħ����>v⟽��?y�P>u�̼�!����1�Vt������辏��� m�i5����>Zx�/�>�,>�q�=h6����=Ej�=��?=�Eܻ�='��=�{�=��=(>(�>�h>�6w?����鲝��3Q�Ib�D�:?�:�>�y�=�ƾ.@?/�>>�2�����{c��,?���?�T�?�?|pi�Vc�>?��Nێ�\u�=���72>��=��2�x��>�J>���=J��ታ��3�?w�@��??�ዿ3�ϿY`/>�7>�>�R�5�1�͒\�$�b��sZ���!?�A;��=̾O�>	��=F0߾t�ƾ,�-=ɒ6>��b=�c��[\��Ǚ=��z�~\<=�Bl=ۉ>b�C>�*�=�E���ɶ=��I=���=��O>�L��л7��P,��3=��=q�b>�&>L��>`�?M�,?#�v? ��>,���T���x�H��Ƿ>�C>$��>���<G�=��>$E??L�5?e.F?���>�� >8�>%]�>��=���h�>곾�S�۰�=q�?�x?���>��j=	v9�����Q#���ܻ?��'?�?5�>���!ѿ)��E�o���Sh�\A(<Jƾ2������)�e�+=�#�e>���>��>_�y>'��=\����xP�>���<��=-�=RI ����:�����V�>�v\=䂲=H�>
?��%���=�	�<qF��A��<�v���=8*>J$�>�F>�߷>�*�=�XȾ%7F>�����<���=hް���G��a��Y}���-���dP>�\>+��_���	?&��>�)+>Z��?ee?���=ݷ/�Y��������z���\��7�=q�>�Fr�zR<�Ԇ[���U���ݾq��>�>���>.�l>\,�e"?�$�w=��FT5���>o������ �N1q��;������ei�Q+պ��D?�D��;��=� ~?��I?�܏?�|�>/+���ؾ&X0>�X��c�=���"q�z�����?�'?l}�>�#쾞�D�ڐξŜ��_O�>X�_��oW�U����+��9�;�N��S�>�����C2�����Dn����D�|0���v�>��R?���?e\,��~����\��`�u��<��%?~�r?�-�>�d?̢?��Q��m����E�,�~=�?Z?�a�?���?PAR>�:�=�2����>�	?TƖ?@��?Cfs?�v?��[�><�;'� >����P�=��>WZ�=�|�=�@?ms
?T�
?m����	�.�����v�^��%�<�==��>���>?Br>��=2Ng=��=\>z��>%�>JHd>@أ>��>�����8�X�'?�+�=*�>�+1?�[�>�W=HЫ��F�<�w[��'B��u+�D����,潧�<� g���N=���g�>Dǿ���?��W><����?����qp2�&�P>�SV>(MὙ�>IG>��~>�֮>���>�)>S�>�?,>C��Vn�=��ܾ�i� M�	D���羯&V>H�����=��� �E�ez���N�euf��~���B���y=��?���<�_Y���4�K�
�;�?�q�>��??�l���;<A�=���>�ɟ>*:��@{����R Ծ��?l,�?��t>U��>J�O?WHS?�� ���u���A��<R�3�)����m���Ӡ���a�i���y��%sw?���?:M*?qaa���p>�x?dp5���Žbޠ<�OҾx�!��}�;��A>럅��[G�[b���k$����g$v=�D?�s�?��!?.�{�����l>�[?ț>j�B?��K?Hy,?Zþ�$ ?$�����?��T?�|?5eZ?��s??4>snN��[���F�<FRt���,�tJ�9�O�U�=ͤ�<Ku=��1=@�`���v����=��4���=;n��s�Q=~7(>�̄=�}<'�=�A�>[?��?u��>_�"?2���JS���{|;?,�'>�6|��򬾊O��y�*>�O?ő�?w�W?eAu>)�s���>�.�>`-�>'K>>�Ƣ>%"���f���H=�ы=�.>�
>��<��9<���Y���΢�=0�>��>�%{>������&>P梾�|��Je>�CQ�q����S���G��)2�xsw�)��>c�J?0�?��=٬�K:��l�e��;)?��<?[�L?b}?3K�=�4ܾ'�9��>J�`��d�>ǥ<[��f��L
����:�j��SDp>�d���a���a>j��?�޾o�n�J�(��A	L=7V��S=V��־#���=��
>�\��� �7	��aȪ��$J?x2k=O���T��Z���>�G�>WѮ>��<�Hlu�oN@��Ӭ��_�=kt�>]b:>�/�����/�G�9��Ć>�YE?Cv_?#I�?g��юr���B�2���ff��6Dּ�??iΫ>ȳ?ԜC>�+�=�ı�WI� �d���F����>�g�>�����G����h���$��-�>��?j�>�_?�R?��?�`?�l*?.F?�@�>ť��H���:&?�}�?�j�=��ҽm*T��9��5F�0j�>(�)?��A���>e?9�?��&?L�Q?�?:>�x �T�?�T��>3 �>v�W�LV���\`>@�J?��>�:Y?Ã?}>>>Z5��`��l>�����=*�>��2?�&#?<�?,��>	��>ʭ����=#��>sc?�0�?��o?A��="�?�82>p��>���=K��>Ƌ�>J?XO?��s?H�J?ё�>���<Y6��8���Ds�y�O�ǂ;7uH<j�y=���B5t�>G�+��<#�;�e���H�������D�#�����;\��>�qu>n�Q&/>f[þ{���ZB>��������|����6�ix�=D�>D?���>ş&��9�=���>lj�>$��I,(?5 ?��?N����b�t�ھ|HL�8ݲ>0v@?���=�l��N����v���^=�m?��\?V�[����$�b?��]?�j�M=��þĶb�̈́�"�O?z�
?H�G���>��~?3�q?h��>E�e��;n����YBb���j��ƶ=�r�>'V���d�5�>��7?�O�>�b>8H�=�w۾C�w��o��Z?�?F �?���?g*>��n��3��^�V���R?|��>P�ʾ�?�Gͽ�Ⱦ)Š�߯���K��[�ʾԙ���Pr�
'��l3�2k����[��e3=�??�o?~�u?
�W?.w�E#I�5rZ��t�P�^�u��~���<�~EH�y�J���~��r����u䉾�
�=�}�W(A�?�&'?T�.����>阾.#�_�̾�C>w����u�=����4=�$`=��f���.�|���-a?۾�>y��>�$=?U�Z��.=���1��7��Y��ڠ4>��>ʑ>EC�>�9;&m,����7UȾ������ʽ#�l>ȹf?:M?��q?2�a(� sy��'��z�<����r)>�P >p��>ē)�ð�=�,��^G��r����s������=�=%?=�d>J�>�f�?�/�>���ܪ��yZ��2*����=��>�Uh?�<�>�4�>�G�]�%��N�>!1m?�`�>�Z�>؎�~#��E~�sŘ�r�>���>h��>)�c>��9�_[\�-���_���4�z�>�xd?b7����e��2�>8X?��<t/�:(�>]z�3k�P���-�b�=pQ
?{n�=2�b>E6Ⱦ����x��ds���(?m;?������*��n~>~�"?��>��>`�?I��>^���jm;�t?HO_?R�J?9�@?�`�>B4=(@��);Ƚ�&��-=��>��Z>Rl=C�=lH�^�\�vm�˦I=rG�=u=��qY����<)⨼P[;<��<�1>�ڿ�L�.�׾�P�����	����k��
�_@�������Dz�(�	����e�P��>d������o���?�G�?]莾�i��
��
�|�Q�H�>q�Y0e�ä����W1�����L�����!�.�N��+h�Hc�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >ZC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾p1�<��?7�-?��>Ďr�1�ɿc���x¤<���?0�@�A?�F(��O���V=��>�B	?h�@>�0�]��Z�����>t�?���?UdX=@;W��U�*�d?�<��E�c��%��=�ǥ=$)=2j�`eI>�>4�L=��@޽�R6>���>0��B��MG^��r�<�rZ>7�׽�n��ք?-�\�=f�ݏ/��Y���@>��T?��>r�=��,?m-H��xϿ�\��`?��?4��?��(?������>�ܾ��M?0J6?��>md&�t�t�9�=�#༸p�����V��y�=?y�>c>�!,����R�O��y���{�=�U���	ſ�@����k�����C� �׽�Žη��oG��V�f���ɞ��Q��="/?>�{_>��\>�S�=,>_1X?Їd?���>�&>�
潁�B�ñ�91�����=Ȑ���v��PX�	�ľ1&�}��8���%�����1=�v��=1/R������� ���b���F��.?Hu$>q˾W�M�EH-<�Yʾ����	������3*̾ݓ1�t!n�aȟ?��A?������V�����T�ro���W?u<����¬�aI�=�ĳ���=�"�>���=q���*3�dsS�e�0?�� ?��ɾ���I>�D��d1=�S(?q�?�<�c�>Q�#?��������W>���=�g�>6��>])5>6���������?2O?�#��6��.��>����;7� ����� >��)� �����!>�v<��]�������%�;m�b?ѭ�>%e�K꾉�V=k����O�i-�?�>B�(?jp?Z\?�CR�w*���p?���-9�=�dV?o9�?C��=U[\�8`��!����e?�-?�>��B%�Q!_��<��K�>�&T?�>?c,`<u���*F���T2���A?B�?O���n��ڊ�����@?!�;?k��>�S2��9�>;�3?ж��Vb�t}���dD���?�7�?��?B�6>��2�k:�=#T?u�#?ϲ���.�p����
�>>w?B=�L��������^N?��?�P�>B ������=�ٕ��Z�?q�?h���^>g<9���l�on����<Ϋ=���F"�����7�x�ƾ��
�󪜾,忼���>=Z@�T�[*�>�C8�G6�TϿ&���[о�Sq�V�?-��>�Ƚ����F�j��Pu�Z�G�?�H�ڥ����>F�>�j����?y�Zj;��Eܼ�#�>��Ӽ���>�cR�����m��E<�d�>j��>b��>b��[H�����?���� �οp�������Y?�W�?��?�?F�<v�n�cWm�K�6�F?�lp?"�Y?�Q�5fV�A6:���j?�٪�ڣ`�F�4�!�D���V>�3?���>3�-�-�y=6�>���>fo>
�.��oĿ����͸���Ѧ?�t�?����O�>W^�?�+?�3�n^�� Ҫ���*����:�	A?�d0>D����!�/>�ɼ��J�?�Z0?��)~�]�_?*�a�M�p���-���ƽ�ۡ>�0��e\��M�����Xe����@y����?M^�?h�?ӵ�� #�g6%?�>e����8Ǿ��<���>�(�>*N>`H_���u>����:�	i	>���?�~�?Rj?���� ����U>�}?��>�p�?���=�?��w>���o)�<���=OV�>j�J�?�?M?�"�>�D�=-XN�;AY�s[w��jn��ء�&,;�'�>�y?QC`?�C>�MQ�,���-��6��Ʌ��K�8�B��c�|9���g=v >?��<��}�()��#.?R�:�#�ۿ����V�{-�?��
?�U?��>�^쐾��a>-�i?c��>��;�0���S��-=Cť?|k�?*?ɽ��ꌽ�+i>5r�>ވ\=k
<��ȹ��8z��B�=��0?T%`��J��k����%>MT�?z=	@�2�?�}a��Y	?;��*v��<�~��R�<�3��d�=��7?����y>���>W�=�!v����a t��q�>!S�?�^�?\�>o�l?4]o�\|B��:=���>�lj?�
?
ꧻN��2qD>�?/�� Ύ�xY�t�e?�@c@ʏ^?l����_ۿ�e�� >ľ%�����g=ym<r�=z�T���q�B��/=bLk= >7+>�"d>VU>��=��U=D�-<�����T&�S ������YX��"=��&�:���ʵ�����s� �Z0���Ɛ�<��	��3Y�&����9�v:���=+�W?�N_?�iI?o�?�E==�X=50���>�X¾�żI��>SO?�g?�x+?�wE���"�[\d��+^�B����x��>�(J���9>é�>&�|>�i��v�=���=���=�M,>-�=��=��q>
��>Y��>᥶>5�>�B<>�>7ϴ��1��p�h�"w�h̽�?e���Z�J��1���9������Oi�=Wb.?'|>���?п^����2H?1���f)���+�M�>m�0?�cW?{�>����T��:>����j�#`>�+ �pl���)��$Q>ql?.,g>�t>p�1��8���O�����ϳ|>��5?+��� M8�}v�%I��ݾX�H>�W�>Z[1�$��s��������i��a�=��:?=:?�կ��o���x�Uڞ��QP>�q[>E'=\�=/O>��g�g�˽��H��'=*��=d^>?Nz>է�=�c�>Ȼ��s&t�Ԇ�>JOJ>n�+>��;?��?�����ҽR���e<�s'�>6��>B/�>_|�=!�S����=�x�>�y^>b�:p���P/�k�M��k>ع��:��lO����=@x����=
�=���Lne���<	�~?�~��.䈿��2P���kD?+?�=|F<��"�_����F����?O�@�l�?�	���V���?HA�?d�����=�|�>8ի>aξL�ٲ?��Ž�¢�˔	�X##��R�?��?��/��ɋ�hl�r0>^%?�ӾU��>���+��M����c��>��#?{uN?%D� �D=��ݼ{d�>R?ZÏ�\˜��IÿB�U�å
?��?��?��������%T����>�/�?�0�?�ԧ>�k
�Cq�L<�>bǀ?�\?՜?�����Q��-V?��?V=?�H>���?ۡs?Ȍ�>�@v�%H/�h%��E���E�=n K;�4�>_j>?���<F��ē�Vd����j�����xa>� $=D�>���A5�����=YT���'��� h�g��>��p>eI>ZK�>�� ?g�>�Ù>��=����������=�K?���?���R2n��Y�<`��=��^�R&?�I4?�x[�9�Ͼ�ը>ݺ\?q?�[?c�>���@>��'迿;~�����<g�K>�3�>`H�>�$���EK>V�Ծ4D�rp�>�ϗ>���@ھ�,���F��IB�>�e!?&��>�Ү=� ?o#?��i>ޏ�>\'D�����FF�I��>I��>$0??~?�?ƺ��3�LY���X���tZ�R�Q>dy?��?�v�>�ۏ��k��8�E�d�8����(Z�?=�f?3�۽�|?���?q�>?�[A?r,b>����:׾톨��`�>�!?u���A��M&�' ��~?�P?��>k1����ս�$ּ��Kx��o?�)\?2?&?B��,,a��¾�)�<9�"��!U����;ٕD���>J�>�����=o
>}ް=�Nm��>6���f<9k�=��>���=I17��{��#0?]Zt��B��O�=��l��(-��> >;��CX?L+���m�[ԕ�͆���S��_�?H��?���?����EX�9VF?W�?��>Y[?��ھ���,�|�c����3��x����=�B>��=�ޕ�3ǝ�ԕ����d������ؽ��>�?[b�>NU�>�L�=.Z�>9���A`��Sʾ�U�L�e����~�D�[�8������
�"��d2�8��.�f�=�>�4N=o��>��?#	�=g^7>�ă>6|"=.�!>>�ϗ>�=�>�eO>�F>c� >_�=v�={R?�z��4�1fҾ�H ���$?�`?G��>x�<&�c�𰭾��?"�?N��?��>��/�/����>�?�����?�h�=�PԽ%���jɾ�.����{��z>�	>}�=<_?��'�U����>�.?�
a��W���[�B���t��<��?��!?F�2���E�1v��T�%Z[��}�x�V�7���(��f�m�����I����U5�� = �2?�?��ݾ����b����[�F�&�9�p> ��>�
�>���>R�=>SK��B;�T�j���2������?E߃?�>mrI?+<?� P?U@L?��>�G�>�Ѱ�٘�>�V�;��>���>��9?>+.?c~0?0-?��*?�>a>U�������oؾv�?rP?b�?f�?@�?�����JĽ�����b�U�x��)}����=�y�<��ս�iu���S="CS>K�$?9�R�b�D�_򾾖�?�"?'�>@��>�6��:����<0�>)�>Z?�>�=Ͼ�����Ti�>�o�?��j�X�<��A>u��=��>����%v>,��-YB>��ͽ��=�&:��ע>|�)>%��=bJ������*	�s���(�>:?b�.>LNB>S���<���&7E�$Ů>X%<+�>��\;��ܾBѩ��"���t���<�>X	�?�t�?��n��ܤ=t��=|'P�RR����(̾�����A?1�?�lh?J��?�1?�'?��=�3Ѿ�B������J�E�?o!,?���>���ճʾ/���3�ٝ?.[?�:a�����:)��¾�Խj�>c[/�q/~����D�᷅����,|�����?���?�"A�b�6�y辥���Z���C?!�>Y�>l�>�)�d�g��$�f-;>1��>�R?,��>�O?�y{?�\Y?��X>��4�����r���<Mc>�;?Ja�?)b�?ӑy?���>
}>�+7�l7�ӫ���F"�Z���􂾥�=U�G>���>�z�>�>-��='ݽn��ܚ-�R{�=��j>���>i�>�m�>�%z>KO�<�DF?���>�¾�þ�?J��~��+x �X`�?-��?�,R?�,�=l��ߚN����.�>���?��?�rA?�Ќ�V_U>g �<��t���/>M��>h@�>޹�=��;�A�>�#?��??�7����]O��`ػ ) ?bA?��=1B̿k<��
������3��8���HV��S�K��P��>���1�(
|�� -�-�d���y�@뭾A�dF�����>��=5�>��=>��4�-cu�A��=sw��ٹ=Q�=��v�ν�)�<1:=����\����̼\B=h����~?>�L?on/?��G?��a>���=�Ħ����>v⟽��?y�P>u�̼�!����1�Vt������辏��� m�i5����>Zx�/�>�,>�q�=h6����=Ej�=��?=�Eܻ�='��=�{�=��=(>(�>�h>�6w?����鲝��3Q�Ib�D�:?�:�>�y�=�ƾ.@?/�>>�2�����{c��,?���?�T�?�?|pi�Vc�>?��Nێ�\u�=���72>��=��2�x��>�J>���=J��ታ��3�?w�@��??�ዿ3�ϿY`/>�7>�>�R�5�1�͒\�$�b��sZ���!?�A;��=̾O�>	��=F0߾t�ƾ,�-=ɒ6>��b=�c��[\��Ǚ=��z�~\<=�Bl=ۉ>b�C>�*�=�E���ɶ=��I=���=��O>�L��л7��P,��3=��=q�b>�&>L��>`�?M�,?#�v? ��>,���T���x�H��Ƿ>�C>$��>���<G�=��>$E??L�5?e.F?���>�� >8�>%]�>��=���h�>곾�S�۰�=q�?�x?���>��j=	v9�����Q#���ܻ?��'?�?5�>���!ѿ)��E�o���Sh�\A(<Jƾ2������)�e�+=�#�e>���>��>_�y>'��=\����xP�>���<��=-�=RI ����:�����V�>�v\=䂲=H�>
?��%���=�	�<qF��A��<�v���=8*>J$�>�F>�߷>�*�=�XȾ%7F>�����<���=hް���G��a��Y}���-���dP>�\>+��_���	?&��>�)+>Z��?ee?���=ݷ/�Y��������z���\��7�=q�>�Fr�zR<�Ԇ[���U���ݾq��>�>���>.�l>\,�e"?�$�w=��FT5���>o������ �N1q��;������ei�Q+պ��D?�D��;��=� ~?��I?�܏?�|�>/+���ؾ&X0>�X��c�=���"q�z�����?�'?l}�>�#쾞�D�ڐξŜ��_O�>X�_��oW�U����+��9�;�N��S�>�����C2�����Dn����D�|0���v�>��R?���?e\,��~����\��`�u��<��%?~�r?�-�>�d?̢?��Q��m����E�,�~=�?Z?�a�?���?PAR>�:�=�2����>�	?TƖ?@��?Cfs?�v?��[�><�;'� >����P�=��>WZ�=�|�=�@?ms
?T�
?m����	�.�����v�^��%�<�==��>���>?Br>��=2Ng=��=\>z��>%�>JHd>@أ>��>�����8�X�'?�+�=*�>�+1?�[�>�W=HЫ��F�<�w[��'B��u+�D����,潧�<� g���N=���g�>Dǿ���?��W><����?����qp2�&�P>�SV>(MὙ�>IG>��~>�֮>���>�)>S�>�?,>C��Vn�=��ܾ�i� M�	D���羯&V>H�����=��� �E�ez���N�euf��~���B���y=��?���<�_Y���4�K�
�;�?�q�>��??�l���;<A�=���>�ɟ>*:��@{����R Ծ��?l,�?��t>U��>J�O?WHS?�� ���u���A��<R�3�)����m���Ӡ���a�i���y��%sw?���?:M*?qaa���p>�x?dp5���Žbޠ<�OҾx�!��}�;��A>럅��[G�[b���k$����g$v=�D?�s�?��!?.�{�����l>�[?ț>j�B?��K?Hy,?Zþ�$ ?$�����?��T?�|?5eZ?��s??4>snN��[���F�<FRt���,�tJ�9�O�U�=ͤ�<Ku=��1=@�`���v����=��4���=;n��s�Q=~7(>�̄=�}<'�=�A�>[?��?u��>_�"?2���JS���{|;?,�'>�6|��򬾊O��y�*>�O?ő�?w�W?eAu>)�s���>�.�>`-�>'K>>�Ƣ>%"���f���H=�ы=�.>�
>��<��9<���Y���΢�=0�>��>�%{>������&>P梾�|��Je>�CQ�q����S���G��)2�xsw�)��>c�J?0�?��=٬�K:��l�e��;)?��<?[�L?b}?3K�=�4ܾ'�9��>J�`��d�>ǥ<[��f��L
����:�j��SDp>�d����پM1,>1������T�7���B�`�(��d�����!�=q:���8ξ�ج�`5=�sB�^�ݾ7���Ά��>����I?��L�\ň��U��9� �O�O>�#0>�m>��/�t��;3JJ� �
��t ����>��>�����Ӿ�3�����>�AK?��C?�?hP�VS��o�ξa�̾�Dؽfw>$()?Cb�>�
?/W�>�eM=m)%��2(�(	Y�@:|����>��>�þ�}\���g��T��M"����>�=�>�٧>�5?��C?u
?�m�?ɹ�>�s>tZ�>`���)iY�K.&?�Z�?�d�=��̽_X��-:�u�E�9�>J�)?�&?���>�G?-?��(?�P?�J?��>n8��@���>�B�>�aV�dF���a>fuL?Cd�>ްX?>��?[.9>�e4��L��E
���O�=�>��2?x�#?b�?��>��>׮����=Ҟ�>2c?�0�?��o?\��=��?�82>(��>K�=ș�>}��>�?bXO?��s?D�J?��>U��<%6��(8��<s��O����;��H</�y=���,t�E�*��<L �;�\���I������D�/���n��;���>_8}>K���P~b>�cԾ6Vm>(Ϗ��)��n���`kA��O�=��e>�1�> �f>Hg���f=E��>��>ͫ��?�b??6"?g��!�e���پd�"� g�>�B?!>�Sf��1����t�� >�Jr?TgE?+�����-�b?��]?�g�&=���þa�b������O?�
?^�G�>�>\�~?�q?G��>��e�0:n����Cb���j��϶=,r�>X���d�P?�>�7?�M�>.�b>?%�=u۾Z�w��q��Z?<�?�?���?#**>s�n�4�U������_�[?��>-/��E� ?K��(�ɾ�G���ޓ�@��̢���������դ�_��^���j�۽+0�=q�?h�q?/5p?��[?;����wb���[�҂���\�_����!HA���=��A��vq����\���8��l{�<�[���+>�sٳ?T�?��"�2
�>�L��?��/�˾�1?>�g�����tp�=���`�=x�?=��j��/��b���Z"?�h�>��>Rk4?�X���@���8���;�%7 ���3>NG�>��>aT�>�g����9�������Ǿ������q}>�`?�vG?��t?(� �;�0���v�Ց#��Y2�$����A>�}�=P��>��f����X�%�Ϻ@��
n��m�J��6O�6��=/?ɪw>#ю>�4�?�f?-3�:S��0e��c0�P!=_b�>*k?O��> .n>�T��_T(�>�>1j?R�>��>\�����p�5����>Y��>���>�i>��.�L�X�*!��\R����6�^�>�Mf?w��h�\�Sj�>�AU?L�� ����>�R;�"I�t�律��C��=�`?���=V�V>Z@���?����߽���J)?L<?���-�*�)k~>Q"?�s�>�F�>�&�?�?�>�gþ�Fx��?|�^?OJ?&]A?\�>rp=ve���EȽ��&��,=�}�>��Z>�m=��=����7\��O��E=��=Ϸͼa��|�<W��˾H<��<��3>��ٿjg<����e��dʾ�������!,�'Í�ܥ齳ז��W�'�ݽ/5'�-Ƚ�`���h�j����h��N�?<�?�G��Ӫ�Q���=���)-���U>�.������R���A��p~��oҾL�þH�!�s�G���Y�jNv���'?ຑ���ǿ�����9ܾ! ?A ?��y?���"���8�t� >A�<M8��ɝ뾄�����ο������^?���>��x.��>��>å�>�X>9Hq>���鞾�$�<R�?L�-?M��>}�r���ɿ%���Ǥ<���?)�@��=?����ؾҐ	>���>��?�ߊ>1萾W�M���ٞ>��?-�n?୽c�Z��Z¼uRl?<u%>j�+�J�]��jS> ǈ<l��=
C��1�q>U�>O8��#��$)+�/Q�>�ˢ>�P�5������-�7�?*�>��0=���ޑ�?߲��=����"�
��+���J??���>�L����@?Ϥ�[2¿�܁��l?�^�?�9�?��%?��˾&��>E5¾��c?V3?�[>b�c�Uf~��A>|��<ċ=���vp��S�z�>|�m��r��.��}��[A�=��������i��2���� ����=� =Q���U��F�5�4��z�������
��I;=���=��,>~�{>�H>�8>�Y?��c?��>�p�=�pڽ�2��*���H�սV ���Q�ՠY�|��'�������B��j��i�
���Ҿ^$=���=�"R�˗��x� ���b�ÔF���.?M$>W�ʾ��M�/*<�Wʾ�����慼�䥽�2̾��1��n�½�?��A?�酿��V����)g�F����W?�Y����쬾��=񕳼�|=�>O!�=���3���S��t0?}[?|���E���)>�� �7=�+?
�?vY<�"�>�A%?k�*���$2[>Si3>�Σ>���>RK	>#���\۽��??�T?N������}ϐ>�L���xz��Ha=kF>75���鼧~[>9��<�ٌ���W��������<�'W?���>M�)����g`��z����==Z�x?҄?w�>qk?��B?g��<�g��]�S�-#��w=��W?�-i?�>�����о�}����5?P�e?��N>�Sh�.�龿�.�9S�#!?��n?7b?�L���z}�S������n6?�v?IA^��b����,�V�c��>���>�9�>):�8��>n>?�n"��<��(����m4�_��?
�@��?��><Q'�ȯ�=&?.�>�O��;ƾ�4�����DFr=L%�>}p���^v����,�qN8?���?1��>FZ�����"��=qٕ��Z�?~�?����-Ig<���l��n���w�<xͫ=�
�&F"�����7���ƾ��
�ʪ���࿼���>6Z@V�q*�>�C8�-6��SϿ0��y\о�Sq���?U��>��Ƚ����)�j�{Pu�$�G���H����v߰>G@W=3������uf�Y�3�=ڞ���>o���[>�9�����4���^8����>���>r��>�5���ɾ�F�?����Nݿv��������H?'�?�I�?`~-?&ǚ=�#U�7�G�eu5��eS?���?A^?��<F����޼�h?7����S�0S!�A�B���b>��:?^�>�O1�U�f<�b�=���>ɞ�=��#�CpĿ�.���_��[�?��?]ݾ4!�>���?h4?���ǘ��9��l�&�=ΓD?��X>Eƻ����md3��Z[���?y]?�?\�'�'�s�a?3%g�|Zv���,����О�>��2��J�F�v�
�/�b����1I���Y�?��?�5�?7���"�8+)?M��>�퐾�꾾8�j=Cx�>Y�>��c>�Zu��Dg>>���W2���>�.�?�!�?��?{=���J���!�=/E~?È�>�o�?@3>z?�$�=�s���[4=��>��	>dM���?�F?���>��c=
�2��+�F�J�J����B���>�(Z?'�H?�$]>�����^輦��B��r��%�����@����C���f>>�e>ur�=��i�s���?Lp�6�ؿ j��p'��54?(��>�?����t�%���;_?Oz�>�6��+���%���B�`��?�G�??�?��׾�R̼�>:�>�I�>:�Խ����`�����7>.�B?Q��D��t�o�w�>���?
�@�ծ?gi�o��>�/�rT��҇���;�U��'�=��>����,�=�9>��ؼ&�?��<����l�M��>o�?w��?�й>	7�?�lt�!��jG?>{s=9`5?tb%?�U>�������=�ӄ>�,ھꑿ=z��ܑm?�^	@��@P\>?&����[ٿxϐ��׾�3־��e<h>�<��
>�ռ���=`IE>h��=��<�`>��>��I>S&>��0>��h>W��>lˀ����je���U���.�֦��b�#��Xh��9�ؽ-����n�f��)�0�{m��g�轀�I�(KZ�̞��O�=B�U?P?,m?ҹ�>��ν�>OR׾:�=y���4>��>��5?��\?�?|s5="����`�|c{��s��#����>�p?>��>�(�>A��>C��6Q>#>�Do>[l�=k�='r[�l��;l*c>א�>j�>/�>uD<>��>�δ��0����h��w�F�˽� �?v����J�T1��>L��ǵ���X�=�b.?�>���=п��,H?�����&���+�G�>��0?A\W?~�>>	���T��C>F��c�j�6Y>� ��sl�e�)�KQ>j?�wc>�ݖ>�tA�VC>��,��F��֓>3�@?+�����q��Mp�>����>	!�>�[i=�"�cД��{`�Q��Q5y=�\*?��>�FػE�k�����^���x>3��>���=D��=�bD>r�����9<������=��=�ZR>\?�8>3�=r��>�#���Z��<�>&�2>;n1>��9?�t&?9�c���`�q��@9�Z�X>�b�>�7w>�=�W��:�=���>�0q>�/ټ��C�Zf���1��?[>H���:U�W�����=d,Ƚ�Q>r��=��yB���$<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ h�>�x�eZ�����M�u���#=���>�8H?�V����O��>��v
?�?_�۩����ȿ(|v����>E�?���?[�m�{A���@�u��>%��?~gY?oi>h۾�`Z�j��>ٻ@?�R?��>�9��'���?߶?֯�?��I>'<�?��r?���>�,��\/��ʲ�zM����z=M�;�>�� >֬��%�F��咿����Kk�uv�j�Y>q�=�ո>��m*��~Q�=���7ਾ;�R�F5�>s�q>O�K>�c�>��?.�>"�>Ռ=�Q��l���l{����K?,��?z��<n���<F��=5�^��,?�L4?z�X��aϾ�٨>T�\?�̀?6�Z?C�>����<��,࿿�����.�<��K>T3�>�H�>�ꇽ�]K>��Ծ�C�J�>)ї>Nݥ��(ھ"���j��2W�>�k!?(��>&Ѯ=� ?h�#?`�j>�*�>aE�I8���E�r��>9��>F?��~?��?�ӹ��X3�	��d硿��[�_FN>�x?�T?Gȕ>���Q�����E��bI�����D��?Zvg?;@��?�0�?�??�A?-0f>��Y	ؾ<ĭ�K�>l�-?���S�f������
;���>��>���>�M����4=�닽�e��D��?I�~?A�N?a���H b���uR�;R�&���%=;x=7,�q>��>bn�����=�o-> K�=Փ�����s?C=F�N>��>O
<�AC�����0?E�,�G���$u=�:~�
�J�b��>O�W>ݧ����U?=0�U��_㬿���
�F�S,�?�J�?}n�?���q�h�cR?*[�?�n?�{ ?�����fо�~ɾ�cW�����V� ��$�=W�>\٨� ���%���Y���-����ɽ�{���>��>]�?���>��C>��>�3��(���<�\Z[�Yc���6��-�����죾�x
������ڿ��"m�AG�>��|��]�>�\?E�Q>�̈́>�J�>mm�<明>�H@>{x�>^*�>ԋu>o/>ϋ�=���+���*R?sK����%�p=⾦^��	9A?`ae?=��>4,���6�����?���?���?��c>��j�/)��,	?M.?`�}�rc?h4==2��;U�;/���p���Hb�2�}��~�>�W���8���K�R�e� ?�?�����Ӿ���I����<=��?��?�����L�z�u��Y� �O���ƼEKo�*F���n�`o��_��L��5\����'����a�+?CK�?5w �_%������b��-<��\>5�>��>���>�<2>��Xn2��qY��T ��T��]<�>�?2�u>��Q?��H?�Z\?�$?�b�>ә�>�	���?}���?�,?�DG?�??� �>���>|�?c}>��{U�/�{�S"?� ?��8?0O[?��'?�>���(���7my�c���"��y����!�=>����6���t�=�#�>R�?W�׽�o-���߾5`Q>n8?q$�>z�>�x��-����@�����>��?%�>�����z�w���n?��? ��9V�<�X%>xz�=�B�uy��4�=���<;�>Q&=�  ��5<�'�=�d�= �=����o򈽵%<�=E�; ?L� ?�9H>P��>���f�X���Y�	/�������_���ֻ����s�b���Ǌ�+݀=&Ԟ?���?�+f>X�>��=�mE�lk׾⾶WǾ�֠=���>��.?}%h?e�U?�(�>�?^\�>GX�dꚿ�o~���[�*�&? !,?`��>�����ʾ�`�3�`�?�\?R9a�A��q=)�)�¾�սw�>�X/�%+~�w���D��ӄ����o|�����?���?�#A�y�6��n�����9e����C?r�>_[�>6�>u�)���g��'�$6;>ߎ�>v	R?���>@�O?��k?�HT?xWm=��h����u���=h`>Zm?R�|?x��?�k�?�\�>��=���ӣ��:���$~�<Q��`����=�|p>&|�>Gպ>.\�>t,>�s6�J�=5\����=�q>î�>My�>ot�>���>��3=%�G?1��>�e��(��WӤ�ǎ����<�>�u?r~�?NJ+?}�=����E��l��!S�>Fc�?�۫?�*?�@S�+��=�>׼���-q���>���>2�>�^�=XED=Պ>,��>!��><u��Y�2o8��N���?� F?���=X4п,v@�(���xѾ�z>!���XS���	��X�<=�g>��c�0���V�
����!ɴ������ɚ�gž?s�><�P>�c���~">�N�=�e_��8K�2�엝�v)��pB���C���@������=u'A=�O�=�%�=�4о.��?D`?�sL?�SB?�5�>̟�>*�1>@�>Ā���?g��>�%>�G����?����۾� �����ʥu�n ^���=����\>t�=C�:;�2�=��=E��=֖ս��4=�ݤ=f(�= e >b��=P�F=t�=� 
>���?s��ı�xT�v��<4�?̉S=|�->����ZU(?�c�Z1O��ȵ���޾�?�	�?z�?��>����>5Ȳ��Ku���>��&�&w>?��>KU=�m�>��>�x`�O�M���w����?m�?��A?�"��s3п�`�>�u7>�f>�2T��k2��O�Zof��N��0#?{�9�2KǾ_�>Bw=&��ކƾ��X={Q=>�9=�{#�&�X�}�=�}���?=��Z=�Q�>��M>�Ԗ=|6��\b�=��\=��=uV>,u��^I�T�뼲�V=�V�=�R_>�1&>A��>u�?Ua0?qWd?1'�>e"n��Ͼ�-���R�>\,�=_�>g��=ÆB>���>��7?��D?_�K?�w�>���=���>{	�>�,�i�m��b�1�����<H��?Ĭ?$Ǹ>��Q<ƟA�֜�b>�!MŽ�v?,S1?�p?�ޞ>�R�ޮݿ�S#��2.��p��#�5<��M=�{a�ƅ���Ǽ�H�!ƽ���=Y�>Ga�>y.�>$t>��4>2�I>�~�>%�>�X�< �\=��:�ʘ<�����V=.	輣8�<Z���O��:��<�]�\Ѽ�2�;7�<q<y�U;�"H>�2�>#��7��>7���޾f�>$~��)�n/M;���D8g�P>~�w�i�g
�#
J���=Y�=u�:뭔��<?->�n/=�R�?j?�C>D�Ϻ_���닿,ʾ�Ѧ��ō�[A=���Ŝ3�+�i��kQ�a���/�>^u�>2��>l#�>Y2��7��i�=���T�,�}I�>J�L\1�$c�S�h�9<��e�� �b�!�<F|<?n:��"��=��s?X�S??R�?��>�D���꿾��T>��Q���=�	� _b��C���8)?��3?���>A[	��1U��˾2m����>�D������燿�O�x�ڽ g¾�U�>Oߴ�mr��!��4��h؍�(�;�f�|���>^bI?���?�|�c�r�o�7�Ę�3#���V�>9?H?y�L>&5�>)W�>d��u.������#w�=�Kp?o��?N��?��(>���==)����>5�
?Ʈ�?&P�?0l?������>��<*>l�ݼbd>5�
>���=WT�=[��>�?�t?s.��3~	�,i�������m���7<D�D=�Fq>��{>�7�>cd>I�=��-=�}>#(�>8�>d> ܠ>�zv>j�s��*W�>x���͈s>��?!�=3ג>^��=�擽���u(��Z��!�O����=��u>G����Ͻ�=�S�>H2ѿ��?��>��%��?4��� s�RZ>�e��䀾ߓ,?��>b�>�O>Ϸ�>�%D>�Y�>��V>[>޾��=�Yᾕ[9�)��#�=��z
�nJ>�E��%����)�h���G���ԾS���`��-}��2�b�����?�,�mQY�84%�<����?[>�>:!?%��:5����=���>�4�>\��ٝ����z�o[Ⱦ8B�?s�?��e>8U�>��V?�?O3�v�+���W��u��C��+g��a�L���j �����@ɽȐ^?��x?OB?�!�<�y>()�?��%��팾k͋>��,��48�_�
=��>�����W�nξ�s¾����=>m?r�?�E?J	W���u��(�>��A?�?`v5?\I>?��?��1<:J,?z�>�K?��#?�&;?�I?��	?gR>)J2�����=�伽�R�����A7��Lѽ����C��V��j	���;�O�<��
�PȞ��j(=H��(�=�M#>8�2>I�>n�>&�Z?�|�>���>.�+?U֊�*��`Ѿt%�>	�˽����tG��٦� W�nc=��\?k�?�vh?um>m�;��)���>}��>fp(>a�K>`�>����?�Ε=��>�\�=���=�F��5������V[�tC�=�&>C~ ?6�>�����[>�[�����'�U>��	��ѻ�����9b�,e�𑾗�>�I*?�?d(�=��¾n�$=��2�5�H?�U)?4 ]?�'^?��5>�.���z�5ƍ��;�����>�6>ax���r���ꬿ�VV��H>��>d����!���=_>��	�I߾Ѻi�tI�kL���'=Z���M=����WӾ8:y����={4>Կ��, ��ǖ�R_��KI?Ɂ\=s~���#a��賾&�>l�>�٫>����a���?A�򿮾�+�={"�>�0>�������9F�`�d�>9vP?d9??�m�?��*��b���C�P���O��2N�Ħ3?Z4i>���>W)�>��r=/����1��!o�����>�n�>$��!����ҾeJ!�r�g�Ԗ�>i�>;
׽wWg?�Je?aڕ>��s?���>��>���>��b�r�۾h�%?���?�h�=Y�=�9��Zr^�8sQ��z?��$?�ߐ� �?Gw1?	��>�!A?l?�>hԂ>����C[��$V>�J;>G�7�2S���^�>�sR?v�?�]A?��?���>��r ��\=b��=��=ʧD?O�?>'d?nx�>l	�>`F�����=[�>��b?�3�?I�o? ��=7?��2>���>�<�=���>�R�>?�?�O?mys?��J?	i�>���<4:���(��r9u��CO����;PZL<0dx=�?�Ss����v�<y�;vӶ�H���R����1E�l���s�;-��>�Rr>����Y�0>��ľY���DA>
���I���&���#�:��ݶ=�M�>=K?4L�>�\"�^~�=:/�>,[�>���A(?/�?`�?��9��b���ھϿJ�x��>�A?���=dm�����a�u�يe=s�m?]�^?��V�Z�����b?��]?�f��=�6�þ#�b���S�O?��
?~�G�1�>��~?C�q?R��>U�e��:n�T���Cb���j��ɶ=Er�>�W�h�d��A�>j�7?MR�>/�b>$,�=rs۾��w��p���?��?5�?���?S)*>��n�4࿆�������1\?��>�O��6$?k,�.Ծ(���Ƣ�%-��K���b���z����#��h}�s�ͽ��=Н?��u?��o?U `?�O��ݺ`���[��	��"�Z�F������B�|%A���C��Wr�;�r��ڳ���[>=+�f�kn*�w��?��-?�/O���>��R��Gоu÷�Z�->,馾ͩ����=��6>K=p_���1��"�Y�H�����"?�'�>bw�>x'A?bp�ѬI�m>��`2��}꾌�>Yk�>EOJ>���>��=�>5���3�\��֒�:�R����>��[?��@?kx?S�[��n��x�����z���Dc����>�FR=��W>�ܩ��\O�#�8�^�M�C�u������v��#=��?E�>��>��?�?`&׾����=�(���D>&N�>�Oy?�q�>�aP>��ۼy(:�FP�>B�g?+��>P��>��Ծ=t��À��B���|>�>>7�>?W>"Ԥ�?;n������*��
j4���=/)}?!�����w��l�>��H?�¼��f���p>C�������/�����`#�=ؤ�>1 �<B�]>å��v��.���'X�}I)?�E?"Ⓘ}�*�7?~>�&"?+��>.�>�.�?�2�>�mþ��F�-�?��^?�=J?%LA?�2�>r�=�ʱ�K9Ƚϼ&���,=8}�>�Z>�{m=W��=����e\��t�i�D=�r�=PμV8���z<Le����K<t�<T�3>�}ۿ,!K�bFؾ���@�D
��҈�JU������h�#볾˘�Ts��;���"�uT�ʴb��_���Wn�')�?;�?v���[$��L��`������r�>Hsp���Mū�{��󃔾RP�}t����!��N��5h��^e�K�'?�����ǿ󰡿�:ܾ&! ?�A ?B�y?��1�"���8�ĭ >A�<%-����뾡�����ο>�����^?���>��$/��c��>���>�X>�Hq>���r螾�.�<��?C�-?��>��r�%�ɿZ���"Ĥ<���?.�@_A?n�'�n�� �^=�$�>ܐ
?�>>�5���U��M�>Ѿ�?�g�?��:=�:X�DV���e?X�A< 0F��uȻ���=`��=0=���<JI>\E�>[��@�F��ܽ�4>:Յ>������<Le�u��<^�\>:�ͽ�����i�?s�o����^���,���f��hF?`��>�X���?)�$���̿b^�沁?�@�?���?k=?���57�>4辉�t?QO?��k>}=I�/ބ���=�\��!������%�h����>8�c\[����"�Ӿ��.=��=�ꟼ���,��s��	��H=g��c��`���==ǩ(>�p̽����)�=[��=�]1>@ٓ>��4>�z8=S��=�n]?�2�?�P?ʼ�>\;�5ȾP\��;4��В½�1�&���P�����ɻ<N��u�쾲�%��Ӿ-���SW�f�;��R�=�rR��W����,�b��E���.?�>'ʾ�_N�?H�:,v;�ث�*Sj�;S��s̾d�1��m���?��A?!셿X�_��(��@Y���=X?���.��.�����=�r���{=�ߜ>��=���W2�';R�.\0?Ғ?�׾�sA���T(>����=��+?�?�$U<̪�>'=%?�K*��߽PhY>3B2>ri�>���>�x>�$���cܽ~�?�$T?²��#!���B�>����1y���m=, >��8��tڼ�u[>��<3����`��È����< (W?���>��)�~��b���#�DL==v�x?~�?�+�>�}k?n�B?�<`_���S����w=��W?g%i?��>����)о���x�5?��e?��N>�_h����a�.�rT��?��n?]^? ����s}��������n6?��v?s^�vs�����U�V�o=�>�[�>���>��9��k�>�>?�#��G�� ���|Y4�"Þ?��@���?��;<��q��=�;?n\�> �O��>ƾ�z�������q=�"�>���zev����R,�_�8?٠�?���>������a�=ً��F̫?U �?s-����<�`�_l�ǌ ��[[<d�=����%����7��hǾP
��ݛ���Ǽa�>�%@�R�F�>��:����f�ο{Յ���Ӿ��s�`3?���>Xý�ࢾ3�k��"v���F�G H�p������>�>�`���K���pu�b�;�3$,����>d���>��^�A2���T��w�{�i=�>�7�>�W�>u_��	/���I�?����\Ͽ}����7	�swX?�J�?�x�?iA?�;�<g�r��t�����P�G?�x?��]?�G�W'l�o��9�j?�"��.;`��d4��TE�x2U>� 3?S�>��-���y=��>vy�>��>�3/��Ŀq۶�!������?N��?Vb�U��>�y�?{{+?�j��E������Ţ*����8�ZA?i�2>A~����!�a=�l͒�Ŗ
?�N0?���8��~?�B�����������O�=A�=>s<9�;��s���d�<y�K�F�K��䗾ퟒ?o:�?i9�?v'������\?;�>-谾۠���l>�`$>m/�>�J�>�>Ͻ *�>Eu��f���q>�J�?B��?���>����J��u3�=�Q�?���>ք?���=A�>��=F��:��[o)>dF�=W
!�G`?�/M?6B�>��=�L;��.�)�F���P�Q����B�%��>nH`?�TJ?�6b>4��e�9��l!��}ʽ��/��Vؼ�5���1��h�$�6>� ?>w�>��I���Ӿj�?�n��ؿ�m��P"'��$4?���>��?I����t��/��-_?�n�>j<��.��� ���$�̙�?�B�?]�?��׾i+ͼs�>��>nA�>}9ս�ߟ�����a�7>��B?�)��@���o�q�>���?��@�ܮ?4i����>�&��z��ˏ�+�Q��d��PH�D߽>����r=\�>������`��>��������>���?���?��>�Ã?�_��LX��O=VAW>�X?���>i�?>&���3�=���>�t�ù������ռ�?M�@��@M�e?	��fܿ��̪�n&��+=*�=�)�>Cཤ��=tuW>�ȏ�69W���;>��I>AQz>J2�>��;>gs$>�vG>���fu�	֟�d�����8�����i	�<2T�����:���ľM젾ZL۾�I��Y<���=!�e�2j)�$Cx��l�=��U?2�S?��p?a# ?�J�U�'>4����=O��m��=�Z�>�e3?LK?��'?��=�ܡ��|c��B�������ք�6�>�R<>�/�>�b�>��>� �9�N>��;>�uw>�>4*=�|"���=�'R>�$�>i��>���>Qd<>��>�δ�))��;eh�oIw�y�˽��?�ǝ�ȖJ��8��G捾H�����=l.?��>���.пn୿��G?�Ɣ�%���,��>��0?W?�h>zҰ���R�5�>���Dj�{�>.���8l�Mx)�=Q>�f?R�u>�r�>KS�b]N�����ž>�/>0�`?m�����޽�����*&��,�=\�>���=�������Q�)���c�r=g)?�F^>��ǁv� ������X��>�$>�,��l�/>@��>��=�p<(O߽���=q�+>��>?~eB>J��=ѕ�>Ok���u9��?�>oc>Y�;>��>?��)?B�C�ɊX�M�e��lC���e>l��>dG�>��=^cQ��s�=g�>��q>3C��	����R$/��@H>I51�/�q�*���=GR��N`�=�Z�=����0B��a=���?3���Mq��i޾�|���l9?��	?Ɯ�=9I�;c��`���㬾5�?	i@!Ԝ?a����T���?:�?�X����>��>U��>
޾�AA�=�?/悔�ϣ��X���(�pm�?Ao�?��=I!���-g�I#>��?�־Ph�>{x��Z�������u�v�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?��m>���?��d?z�?b�S���#����?��n�{��\���u>�"�=p���k�`�����-��[nl�j�)��{�>|X�;���> F��&��:!>驇<������,�E��>K.�>��=��=>y?�>ZN�>nU�=�g�t����m;k�K?���?����1n�:�<��=ܴ^�'?mI4?��[���Ͼ�֨>^�\?�? [?�b�>���+>��F迿!~��3��<C�K>P3�>�I�>� ��LIK>
�ԾM2D��q�>З><���>ھ�,���}��+C�>�e!?���>]Ԯ=6� ?\�#?j>�J�>mE�Z3��o�E�8��>�l�>,*?��~?��?����e3�[���롿q�[��IN>Qy?�G?n��>ނ���s���kG��J��E�����?-}g?[Y��
?s&�? q??�A?�,f>l��$ؾɘ�����>/<?z精-:e�x�lP��(k�>�b�>���>od�hV��[i½_1��sо<?��x?`�&?C��(Q������<��=a3��L��T��Ay�=k+!>���<t�9gy�=���=����.x��,l=(�=:�>�j=>]	l�&Yz��H2?żn�����=�t��~S��D�>Y�A>��Ͼ��L?p�F��Ǉ��Ȱ�`�$%!�5��?�m�?dF�?z�E�|m�=2K?M��??��?�Y��k7о⾯N�����Ư��:>�x�>Ͱ*��4�!;��w���͂�B��M����d?���>A�?���>U��>�@�>�w�ٟ ��8־][	���\���E�A�_��0�&����R>��f���־A<���>�	2�E��>e� ?0�>�{�>�;�>B*E<�%>�>N
�>��>6�>�x�>|m>	��=��ҽ\�R?�@þƩ(�'&�ӯ�&�A?�d?���>��l�����?6�?�Ȝ?��z>B[g��+���?  ?���_�
?�9=�H)�T�Y<�Y��D��>ソ�=��ȍ>plսj:��M���d��,
?�?`+v���̾�I�{��o�<JX{?V)?y���i�P��v��l��3��:��,����ۍ�[z���q��!���<z���t��/��/�3*/?�u?vT�����g�$f���5�|]>���>�g>�`�>O~�=���R'��f�|���I]����>��?1��>(=U?��A?C�_?V�?M5�>Y�>e��}?i!�=�?��>5?,�G?�Z�>
��>�?�K�>�5W�^��_ž�F?)�?�7+?�=?{T#?C�������t)>��[���ƾ�>���<�����z��.�=�W�>P�?�����8��C���*k>u:7?���>���>ُ�����]x�<���>��
?�"�>6����
r�	z���>ւ? F�M�=�B)>�#�=�V��s^�B�=����q�=Ƞ��S�<���<w��=�̙=pG���d�sG;��B;�[�<�P?z�,?��u>�ʿ>��ݾ��0�R@�;j-�%��1K��/o���E����~��+��I'��e ��ҋ?��?L�K>H�=�D=>�12����]� ��*��q�_?SM0?��o?��?X ?k!�>���=N�!�������T���
�&?A!,?<��>���J�ʾy񨿻�3�U�?�[?,<a����<)�ő¾�ս�>�Z/��.~�T���D�l���\��d�����?���?�#A���6��x辽����Y��F�C?"�>Z�>��>�)���g�4%��2;>��>vR?��>�oQ?�/y?N�\?<>*�<�y����C��%Y��>� D?4��?���?Az?{��>�>B�"�y���d �����������dLC=�j>�x�>^h�>i��>m��=/�-���^2�w��=ISc>9p�>���>�w�>K��>���<��B?DU�>j�;�������|���Zن�
%}?�~�?�?z/�2x��4O�E������>n=�?Y}�?��%?w�e��=���������_J��E�>��>݃�>���;S��=N@j=���>���>��������.�QT��O?�~F?ɇ�=�C��P�(���*=����D�M>#f���Dپ]1ԾD�����:>��6�|��=�˓<����^��qΉ�0�r���Ǿ_CԾ%j?�3�<K�g=���|�g>5�]����Xbҽ���(�L�&���4�����%Wv��i��T����B������<�����y?4[Y?l�4?�~'?�ҩ>�Y�>���=�.�>ǋY=j
?�8�>�H�=�*��x��/�����׾-�I�⾌�h��7f���=n&�ղ�=!���[>�.b=�n>�F<1㦽�Xp=����=>>�!>))>��=0>sx?m8��������o����=��?ļQ�+K=�	Ѿ!� ?1�Ot�X鲿nI���t?k @y�?�� ?��B��p�>^x��,۾N��>Q�m�çl>rK�>$u8>���>p��>.�ɾYY���p��i�?5�@�O`?5Ч���Կ���>�h8>{�>�S��2��JW��)e�7[���#?t�;��ɾ�L}>�h�=���e�ž>�O=��9>%�U=dB�gZ����=�{��}A=��H=�ʆ>�C>���=:q��>u�=X3=Z�=�dU>��Ⱥ�)�z��il==�d�=��e>�2/>Ҙ�>�?�W0?�Vd?���>dtn�}!Ͼ����'n�>���=q��>�i�=�jB>%��>��7?җD?��K?I��>���=:�>t�>`�,�T�m�g�&r��X9�<���?�ˆ?��>��Q<`.B��z�T>��{Ž|?�>1?��?=�>���.�ῦ�*���:��ͽ�00=�^�=�k��4��a�=���u�r����=���>TC�>n��>�X>��&> 9S> ��>��>{>zl>{5�<@0�<}��:ٝ=��8<��F=�@>1��=KKa�/ �<���PR-<Q(o�=��*���Z=>���>"z�;?�>��Z=ټ�^>Ja��>Y�m1�<E?Ͼ��f�	���&�u�|��F�ӽO�8>U�>�b�������?)��=���=Q��?]Gy?	Q�=�P(<[�Ծ�ك��¾%�J����=�蟻6����7�v�s���O��#뾊�>���>�
�>�\s>=�,��=�~^=�)�c�5�/��>5���c+�?���@r����j4���i�9r�ehD?�臿)��=[m|?��G?�͏?��>�W��vEվ��2>s ~����<���C�e�cz���??�8'?��>��V�E���Ͼ7�ɱ�>�;ƾM���r̕��aB�0�������c> �;-�ھ�)�n!��P���_�0�-}C���>:E?J��?Z�������T��|��O�.�>��G?[M4>���>7z�>x`$��\ ��(��k�=�u?�X�?cJ�?��\>�K�=}�����>r]	?x��?뱑?g�s?�=����>ޤ�;��!>Hژ�m��=�>-�=B��=?n�
?�
?�۝�G�	�"'��~�EV]���<lա=.1�>X�>s�r>|��= Qj=?_�=_�[>���>"��>-4d>O�>��>�q���o���� ?#���P>!�?|�;>s�A>H�5<�ؽM�h�<���Gq��'���!b=��=*��=Eܴ=��	>ȟ�>Pʿa��?ߤ>�\&�(?<V۾�i���Ҕ>���0x�;� ?��X>��>sa�>ˍ�>�w[>Om�>��!>4�־3�>�}	�J~%���6���R�E۾�`K>���.��W
�����C��7��:��P�f�� ��@t>�u<��?�l��Ro�O�.�g�ν�t?��>]	.?�D���[����	>Ϫ�>+s>����3X��;����ؾ��?���?h�o>���>�nP?u?_S�Ou̽��T�^[|�L�P��u�=`b�/����Y�����~����U?�Pz?�C?�|�<z{>�_�?�1�g�n�D��>�R&��1�U��<XiV>lh��g�]�����@ۭ�;/�T�=�(V?�@�?~�?�EJ���B�<f�>V�P?.w�>:9?S8a?��j?��0=�xW?�?"��>vH)?*X?�?�]�>�+�<��Q���B>��������j���\�(�\��>|<���=<�=ݜU��3�'�<G�g�R��=R:����J�7=�<)=v��=�}5<b~Y=GŦ>��]?�D�>��>�7?<���l8�0���E/?�8=�|����������񾏫>��j?E��?
fZ?~!d>p�A�o�B�9H>Y�>d�&>qU\>~��>qa�ՍE�i�=�1>,	>04�=�M�8���ݿ	����a��<(G>���>f��=w���b��=j��߅	�6+>J𕾽=������O�>@.�7jž��:>�wH?�?�sv>�����d&=Q�6��!2?�??��?!^A?HW�>����@}�bې�|������>*�>�Վ�u@��P���NG�C����>d�̾(�R�m>�(������+I�	�[�iB,�I%νbi�������^F����<a�����Ͼړ+�Ԙ�h����<?�����r���O��u������=��>в�>�E����v�!������ah{>�i�=��&�9Ѿ*�-�@���4v�>��4?o�F?5�?n�$�*l��hNྺվ���bm)��NN?n��>��D>�>��>�=�ʏ$��i����>�1�>(S� �
�&ho������P���C>��>S�X=B)?5K�?I��>Tr�?Y�B?��>�H\>���yԣ�0 &?��?f��=pUʽ�WU�rn9�jF�~��>�(?�b@�睙>-,?�?E�'?amQ?y?�>��^@����>��>x�V�����\c>E-K?��>UY?�v�?�RA>�D5����\U��RV�=X�>N3?��"?�~?r�>�2�>�j��{Ɂ=J2�>�c?t!�?߷o?v}�=�6?��2>j�>C�=&ҟ>Ҙ�>/7?[0O?�os?��J?ҳ�>IS�<?��kŵ��q�,K����;RO<)z=� �r)t�)��yk�<���;7s���䄼��QE�񒼄(�;Y_�>{�s>����0>��ľP��R�@>�{���P���ڊ�8�:��ٷ=*��>��?<��>�V#�{��=���>qH�>���/6(?�?(?6!;$�b�
�ھ"�K�U�>�B?���=��l������u��h=�m?5�^?F�W��%��<�b?��]?�g�=���þ��b�ވ���O?��
?"�G�V�>�~?��q?��>u�e�J:n���Db�7�j�6ж=dr�> X���d��?�>6�7?�N�>��b>x#�=�t۾��w��q���?��?��?���?�**>@�n�I4�}���G܏�c^??٦�>�^��*#/?J^>�	��Yվ���w���4ľ�߾gg����X����w�K���;��S=^?*��?2tX?Ag�?৾]�� >�
��1��B�A�u���+G�HR�*�wb���1������~��\�=Bx�C�ʙ�?�#?�=@��R�>�ٓ�>���˾7D>ɢ�����=�s���Uk=>�t=��O�)�"��魾�d?'R�>r4�>��??�eW���8���+���>���I�)>V�>>̑>l��>LR<�*�C���~Ҿ�|��XŽ�w�>��U?8�F?d>x?s�<���5���o���#��g� 2��,ge>S��=�Q>��{��XE�g�0��<�(q���8Ӑ��
���D=��9?�x�>��>ٲ�?��?�\��ӈ��m��=����=uu�>ۏd?�9�>��r>u�����4�9I�>��Y?ɂ�>s�>˾��,�+�d���)��>�>�k]>$��>�\r>�[��g�`�E��������[3�(aZ=�4o?��v�s���錕>Lj?��+�����z��>X�?��|�^C��a?��[`=b� ?���=w:\>���	�G��	ľ�<(?�K?�ʏ�^�)�2��>#?-.�>���>��?ğ>�I�����;�?5�^?12J?tz@?��>�h=G���]�Ƚ�&�0 =���>�\>�n=�/�=����\����A�H=S7�=o�������O<=}���<��<�6>��޿�A4�z����I]̾{�	����O�r�,��{�;��4Ӿ׸��r�'�م׼�U�7�@�!�o�������@�7E�?���?@��?-�r��רp����rU>���ҽ��ǾLL�w�����̾�;���d(��W������c�:�'?����޽ǿ�����:ܾ$! ?�A ?�y?��4�"�Ē8�ӭ >�@�<f/��Ɲ뾫�����ο7�����^?���>��%1��.��>᥂>=�X>Iq>����螾�0�<��?/�-?��>�r�'�ɿ_����Ť<���?4�@RkA?0)���p�T=\b�>��	?��@>��0�\L�j̰�PV�>��?<��?��H=�:W��C���e?�q<�F���Żt�=cĩ=>�=�����J>+ޓ>�� �+C�k޽��4>��>�.%���v|^�ٺ�<L,[>��ս����tr�?�p���v�u.�V�v��5=[�??e��>�=��%?/T���ο��]���G?�h�?���?��F?�����O�>�T߾�Q?#<2?�Ƣ>�XB��Bo���=O��wjP�6;�]MU��l�~�>�%]>jTR���@
>��g��;�=��ӍǿC��6*����<��л���`�$�)����R��p��:!�,�;� >/�X>m[>^ws>Fa�>'��>}[f?�{�?A��>H~�=��$��������X��㾲G����۾���o���k⠾��^�����)���^��@0=��R�=%�Q�Չ���� ���b���F��.?�@$>��ʾ1�M�6�%<Oʾ+Ԫ��m���_��;W̾��1��Kn�D��?W�A?p酿.'W�����Z���I�W?�$���E۬�IZ�=�>����=�>�D�=���D3�zJS�?N0?��?7&��˺���*>7�A�=,?�5?��N<Ԫ>��$?�=,�E�n>[>�45>V4�>���>m�>� ���%ܽ��?�:T?7��FĜ���>�)����y�^�b=<�>�'4�W�9{[>)��<���t=�%#���n�<Q&W?m��>G�)�+�`��=��u_==��x?��?�2�>�xk?��B?�*�<Fe����S���hsw=��W??&i?ں>����о�~��e�5?F�e?��N>�~h����u�.��R�0%?��n?�]?!:��^v}�������?o6?��?ף���~��*����9��{�>�,�>��?/!3�<�>�?������H����,�굥?;�@���?d�=u*<�q�<#��>�� ?>�����@��������= +?$�!�����O�B��og�?��?��?Z�����=�ו�L�?��?����]j<����*l�%������<��=��;x$���7�7�R�ƾ��
�6�������v��>�W@h��cK�>��7��+�qLϿ����о�r���?*]�>��ȽѼ���j��Nu���G�żH�r���lI�>0�>���c��r�{��m;��ʞ�i'�>-`����>a�S�P3��W�����2<�>��>Ά>�轾n��?q|��\1οO�������X?)`�?i�?�q?�|;<y�v�d{��)G?9�s?ZZ?�5$�]�K�7���j?�ɧ��_��23�<�E�4�Q>�(2?T��>�+-��|\=�O>���>S�>�/���Ŀ����k@���b�?���?S#龫��>�p�?�,?C��њ�ʓ����)�o�X<;CB?};;>�~���)#��;��ْ��?H�.?����g�=�_?}�a��p�h�-�!�ƽmܡ>��0�=e\�aS������Xe����Ay�L��?^�?E�?��] #�6%?J�>����47Ǿ��<g��>�(�>w+N>�W_�	�u>����:��h	>6��?~~�?j?������jU>��}?�&�>��?���=�x�>�"�=���(.��c#>%�=w�>�5�?R�M?PI�>?��=��8�; /�uZF��OR�%���C�b�>��a?/~L?2cb>5���]S2�� !���ͽT;1��Y�>@���+��t߽�5>�>>~(>'�D���Ҿ��3?>L@�����К�q�d��8P?�#�>e(?N{� ��n�=�n?_�>>�07��Hb{��Ɂ=L��?���?i9?^@����޽-��>��>�!�>�S1�7ӱ��Q��9~�>Ф2?�e�(;��(n���n>�(�?��@	S�?��d��	?�+���_�����0����=��8?����5s>���>�e�=�[u��8��[�t��@�>��?*�?�S�>)Ym?õo�εD��6J=�>��l?�(?���;����orB>�
?N6�،�\� �I[d?��
@��@��\?�;���Z�}꥿�M��U�Ⱦ�ڠ=��=,�,>�Lw��#,>��Ȼ�r�<�G<���=aT�>K�>Zã>�Pc>�y>��>]ƃ�"����^����)���%b��>����־W 6�\�Fp�=p��RE�'���r�r=�ݽ�:��Y��B�>��a?��R?m�?��>+���@�1>�9�����<i�D���>ʂ�>#�=?,�X?�,"?�Ù=I���Wo^�z"x�#���~���i�>�8l=���>�8?��>���=�@e>�ہ>U;0>^7¼j<]=���v����>c �>��>��>HB<>��>�δ��1���h��w��̽� �?M���M�J��1��#:��Ц��ag�=�a.?a{>���?пs����2H?-����)��+�,�>��0?�cW?�>�����T��8>�����j��_>, ��l�n�)��%Q>�l?�Zf>7ow>��3��{8�ZP���%�|>e�6?V��AG:�}du�T�H��Y޾ǬJ>[f�>o��v��ӗ����~��Bi��*w=N�:?S?����Bg����u�2۝�)mS>�\>v=/��=�=M>�b�h����VG���9=/�=��^>�A?z'+>F|�=c�>�[��P��֪>�B>(T)>h^??+�$?/"�����؃�Q�.�`u> t�>�I�>�>" J����=��>w.`>��"*��!'�~?�3V>��u�w�_��Sq��\�=D����2�=<��=�] �M�<���=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ܇�>��w�;������Xe[�8��=1��>�O?k��m0�d7�s��>|#�>� �:(���ÿTG�fW?���?�m�?Dp�~ݲ���Az,>�=�?��t?[� ?���&�t���?�f?��o?���>���sĵ��/Q?�à?t�q?.I>G�?�s?���>i�z��h/���������~=��U;ņ�>">[���YGF��ʓ�!n����j�����;a>�v$=F�>_��l����=�_��5R��Cf����>�Lq>��I>�j�>h� ?���>Dƙ>�)=Y���3���Ė�D�K?���?����0n��B�<]��=��^�t&?�H4?�K[�B�Ͼ�ר>�\?�?�[?�b�>���N>��迿W~��ê�<��K>�2�>(J�>���JK>U�Ծ�4D�<r�>ϗ>���W>ھ�.��Nm���C�>Ae!?���>�Ѯ=P!?��#?oi>'��>tG��N����C���>q!�>��?�0{?�?��ľ��4��.��s�����Y�WO>�{?ߕ?|�>��������t༲���\j��y��?-Fm?R���{�?k�?��7?�%B?*A`>y	1�\3پ�V�3�s>��!?��OB�^&� @��;?tW?_��>`���6�׽e*ټT$����Kt?B�[?��&?"���`��þ%?�<�� �U��9U�;�5j��u>k>[/��㓵=�>�g�=��k�"X6��]h<>�=�>�U�=y�6��Ռ���??��� v��69�9,�t�&.P��:>o#�>���,?����O���	��&r���H4�U�?���?�0�?��0�y��m?6om?lL?��?��1��C������V��<���J�Ͼy	�<�Ф>峢��T;�Й���$���|��&2��𮽆�>�`�>I�&?�3�>���=�m�>���t=,����]�޾b3o�����4���6���#�L����7�و�]����9�6 �>Z߶�� �>k��>rr>ya�>�>��C=��^>��&>A{�>���>W̓>�8>Q �=����qq��KR?�����'�U��ֲ��X3B?�qd?>1�>�i�5������o�?���?Js�?�<v>h��,+�vn?z>�>D��Tq
?�T:=:��:�<V��k��3��W�3��>E׽� :��M��mf�xj
?�/?�����̾-<׽:q��Fс=�K�?��#?%(���R���q�2oW��P�FUN��k�>V��[$�t�n�T����h��č��1�*�ҽ�<(�)?Y�?�� �E󾯠��n2g�FY;�IU_>�>���>{�>ޣ@>��B�/���[�g'�P?��X��>�bx?~>�OS?i�I?��`?�ZR?2P�>�s�>%W9��}�>G�q>�?*
?w�M?
3?+P%?��?��>�>�/������ϾO�?j��>π+?{�.?���>#�S��+��\�=�襼����q���ٮw���<����|E>�D=�=z2�>+X?O��۪8�F����k>ف7?A��>���>w���0�����<`�>~�
?B�>�  ��zr�~a�tY�>���?���(�=��)>O��=x����(Һ�V�=�������=�J��k;�֓<{��=��=�u�Ϙv���:���;���<�?Q22?�6<>�q�>ũ������xʾ0�X��~m�s��v��̿þ����˓��q�����=>E~g?�n�?�T�>���=2r�=�! �r[��_������ \��x?�{?gGO?���?�m5?긝>xF>���;���݉�a���?5",?���>���ѥʾ��F�3�/�?�Q?R6a�Z��6)���¾#rս��>Uc/��2~�n���D�K7����� ���ʙ�?��?RvA���6�n�J����@����C?�3�>YR�>��>ݻ)�J�g�0.��;>�f�>��Q?(��>Z�^?��b?��?cD=>�^�����_���%��l�(>n?��?���?䗑?³�> �ͻm�[�cb'��� ��	ȽR)��[,N�+��=H-�>+Ĳ>�v�>��>+P�<�c>��ܽ2����>p�>}1�>T��>�j�>j/�>�h�<��A?�`�>�hӾ�����㸅�v��E{?�Έ?�c ? ��<ή���K������>�;�?�\�?��(?��W��R�=�Y	���+i�&�>m��>��>U��=���=�?.>���>@�>1�񽨵���&��8^�;P?�D?a��=t�ÿ���H��j����O=�o˾�b �8ʨ��r8�s��u����,A�;]�U���������̌�b���ySξ	��>��.=<w.>�S.>N��
ؽ���<x�>�>��q=��<�aL=����T>��Lm����ݿ[�����ߏ_��ʾ�4}?��K?;�,?�D?���>Z�">�Lżd�>�jK�w�?�O>�`�"����<�����'_����ܾfKپҽd��O����>\�i��
>`;> "�=^��<��=߁=��r=n�C�k�$=ƫ�=+�={H�=�j�=��>˶	>��{?�N��j2��J�P��½i.?��>.�=� ž�A?n�>���=*��0A���?>�?B��?�?��k�R�>A����_��(�=����>���=�D$����>-&>�$�	z���?�=��?�@�%@?�V����ɿ+�->C�4>���>x�l�N6��e���a��P$<?�_A����z�?>�ƽL�����+.㻻��>�D&>�$���	T��<~򼝍 >wc�$s(=�.->ԅ�=�琽z�>�	w=Z�>9a�>��,���� �<>�j�=�9>��]>�{V>��>��?�b0?�Pd?)E�>��m�DϾ4���O�>a��=�M�>}P�=[�B>;��>�7?̩D?�K?�}�>P�=F��>` �>Q�,�۰m��M�䶧��r�<e��?�Ȇ?(ø>�aN<A����l>���Ľ�v?E1?q?��>�v����(�%��.��5��T�z9<\+=ȧq��
O�����D����ݽƪ�=��>��>̺�>��x>�<>��P>}2�>��>���<�q�=��?�=��<�#��f	w=Sn��c�<�[⼰#��a0��#�'����M;z ;�YB<���;%�>���>DIV�	R�>��>�9���C>Z�ҽ�M��n�<c�þ{`��Dc��f����@��Y��p�>�H{>d� �xc��1�?K�H>v��=Ǔ�?�u?$�b>P���GҾ?9��[]�������=��C=h;��,��Tr���N�nǾ� �>*�b>�>���>�gE�j9H�B�=������#����>��,��0������Bz��2���ܦ��3_�����{9?�gw����<0�`?��c?�7�?vµ>C_\=�ܬ��=�$��#п=��+�.F���<-�?E�?�>�>�p�f�m�%���T2
����>�0�����O����)��R������T$z>�۾o�羷
?��x������%�O��y����>b�Z?:�?򖉾-ښ��L��A+��|=�(?g��?�;>�V�>M?R����ž��W�{>�<��J?���?�k�?C�>;x�=�A@��y�>��
?d��?��?�3g?�f��>��=�G>�9ƼW1>>&>rh�=Q��=��>�?p0 ?G���+A�	����Z�J�1��D=�X����A>�\�>浐>w�=�� >5r�=7�D>�=�>�Q}>�.>��>eۗ>�<d�S� �:��>��|�>�;��)?B��>K��>�����ꔺ�6���s�w	���k�II�<9@e>ΰ�>>�8>]�Ͻ��>B8ֿ쩩?kt�>��!�FaB?�P�����l�+>���>u�J����>~ �>��>$��>��o=g\>�ʏ>)�&>��j�=�+Ծ��A�h���-I����=��]���h����W����,����ӾJ_��b��E~�vwH���ǽC��?)�E����GM�Z��=$�?I��>�	?x�D�E�!�w�p����>�=̂���懿!���o:���B�?�\@�Ǔ>�פ>��5?�_ ?��k�ᦠ��/�7>��q�v�#�����|�$(��Sφ��H��7A�E#:?h�t?�}Q?)=�	g>���?�� ��蕾eA�>)��8�<���<��
>�E��� �� ϛ��un���� :�?j?�T?e(?D��:��:����>�'?e%X>qg?�F?Kc�>9Ne<a�z?�],?fǣ>.?ɉO?}X=?�C?N)>a򳾨5��)��>XPD�����
�?���н��*�}^�=5�.=���=�B�ͼ�hn���ٽ����L3<�@ü%�=�8�=���=P��>0�]?y��>v�> �6?����<7�X�����+?S�=�q������U���&������=��j?.��?$[?`�g>:zA���?�f�>���>d8%>�\>`��>����B�΃==�>�>��=3`��恾`���s��7��<�}%>���>�t>@����s3>/����.m�D�p>�@i��Ǿ�i�'�I���3��􆾢#�>ִG?Qu?��=Va�7Ҝ�.�a���-?��6?$�N?��?K-u=B��<<�K�P��A�Y��>-sX<���߆��KO���";���+���|>~d����پM1,>1������T�7���B�`�(��d�����!�=q:���8ξ�ج�`5=�sB�^�ݾ7���Ά��>����I?��L�\ň��U��9� �O�O>�#0>�m>��/�t��;3JJ� �
��t ����>��>�����Ӿ�3�����>�AK?��C?�?hP�VS��o�ξa�̾�Dؽfw>$()?Cb�>�
?/W�>�eM=m)%��2(�(	Y�@:|����>��>�þ�}\���g��T��M"����>�=�>�٧>�5?��C?u
?�m�?ɹ�>�s>tZ�>`���)iY�K.&?�Z�?�d�=��̽_X��-:�u�E�9�>J�)?�&?���>�G?-?��(?�P?�J?��>n8��@���>�B�>�aV�dF���a>fuL?Cd�>ްX?>��?[.9>�e4��L��E
���O�=�>��2?x�#?b�?��>��>׮����=Ҟ�>2c?�0�?��o?\��=��?�82>(��>K�=ș�>}��>�?bXO?��s?D�J?��>U��<%6��(8��<s��O����;��H</�y=���,t�E�*��<L �;�\���I������D�/���n��;���>_8}>K���P~b>�cԾ6Vm>(Ϗ��)��n���`kA��O�=��e>�1�> �f>Hg���f=E��>��>ͫ��?�b??6"?g��!�e���پd�"� g�>�B?!>�Sf��1����t�� >�Jr?TgE?+�����-�b?��]?�g�&=���þa�b������O?�
?^�G�>�>\�~?�q?G��>��e�0:n����Cb���j��϶=,r�>X���d�P?�>�7?�M�>.�b>?%�=u۾Z�w��q��Z?<�?�?���?#**>s�n�4�U������_�[?��>-/��E� ?K��(�ɾ�G���ޓ�@��̢���������դ�_��^���j�۽+0�=q�?h�q?/5p?��[?;����wb���[�҂���\�_����!HA���=��A��vq����\���8��l{�<�[���+>�sٳ?T�?��"�2
�>�L��?��/�˾�1?>�g�����tp�=���`�=x�?=��j��/��b���Z"?�h�>��>Rk4?�X���@���8���;�%7 ���3>NG�>��>aT�>�g����9�������Ǿ������q}>�`?�vG?��t?(� �;�0���v�Ց#��Y2�$����A>�}�=P��>��f����X�%�Ϻ@��
n��m�J��6O�6��=/?ɪw>#ю>�4�?�f?-3�:S��0e��c0�P!=_b�>*k?O��> .n>�T��_T(�>�>1j?R�>��>\�����p�5����>Y��>���>�i>��.�L�X�*!��\R����6�^�>�Mf?w��h�\�Sj�>�AU?L�� ����>�R;�"I�t�律��C��=�`?���=V�V>Z@���?����߽���J)?L<?���-�*�)k~>Q"?�s�>�F�>�&�?�?�>�gþ�Fx��?|�^?OJ?&]A?\�>rp=ve���EȽ��&��,=�}�>��Z>�m=��=����7\��O��E=��=Ϸͼa��|�<W��˾H<��<��3>��ٿjg<����e��dʾ�������!,�'Í�ܥ齳ז��W�'�ݽ/5'�-Ƚ�`���h�j����h��N�?<�?�G��Ӫ�Q���=���)-���U>�.������R���A��p~��oҾL�þH�!�s�G���Y�jNv���'?ຑ���ǿ�����9ܾ! ?A ?��y?���"���8�t� >A�<M8��ɝ뾄�����ο������^?���>��x.��>��>å�>�X>9Hq>���鞾�$�<R�?L�-?M��>}�r���ɿ%���Ǥ<���?)�@��=?����ؾҐ	>���>��?�ߊ>1萾W�M���ٞ>��?-�n?୽c�Z��Z¼uRl?<u%>j�+�J�]��jS> ǈ<l��=
C��1�q>U�>O8��#��$)+�/Q�>�ˢ>�P�5������-�7�?*�>��0=���ޑ�?߲��=����"�
��+���J??���>�L����@?Ϥ�[2¿�܁��l?�^�?�9�?��%?��˾&��>E5¾��c?V3?�[>b�c�Uf~��A>|��<ċ=���vp��S�z�>|�m��r��.��}��[A�=��������i��2���� ����=� =Q���U��F�5�4��z�������
��I;=���=��,>~�{>�H>�8>�Y?��c?��>�p�=�pڽ�2��*���H�սV ���Q�ՠY�|��'�������B��j��i�
���Ҿ^$=���=�"R�˗��x� ���b�ÔF���.?M$>W�ʾ��M�/*<�Wʾ�����慼�䥽�2̾��1��n�½�?��A?�酿��V����)g�F����W?�Y����쬾��=񕳼�|=�>O!�=���3���S��t0?}[?|���E���)>�� �7=�+?
�?vY<�"�>�A%?k�*���$2[>Si3>�Σ>���>RK	>#���\۽��??�T?N������}ϐ>�L���xz��Ha=kF>75���鼧~[>9��<�ٌ���W��������<�'W?���>M�)����g`��z����==Z�x?҄?w�>qk?��B?g��<�g��]�S�-#��w=��W?�-i?�>�����о�}����5?P�e?��N>�Sh�.�龿�.�9S�#!?��n?7b?�L���z}�S������n6?�v?IA^��b����,�V�c��>���>�9�>):�8��>n>?�n"��<��(����m4�_��?
�@��?��><Q'�ȯ�=&?.�>�O��;ƾ�4�����DFr=L%�>}p���^v����,�qN8?���?1��>FZ�����"��=qٕ��Z�?~�?����-Ig<���l��n���w�<xͫ=�
�&F"�����7���ƾ��
�ʪ���࿼���>6Z@V�q*�>�C8�-6��SϿ0��y\о�Sq���?U��>��Ƚ����)�j�{Pu�$�G���H����v߰>G@W=3������uf�Y�3�=ڞ���>o���[>�9�����4���^8����>���>r��>�5���ɾ�F�?����Nݿv��������H?'�?�I�?`~-?&ǚ=�#U�7�G�eu5��eS?���?A^?��<F����޼�h?7����S�0S!�A�B���b>��:?^�>�O1�U�f<�b�=���>ɞ�=��#�CpĿ�.���_��[�?��?]ݾ4!�>���?h4?���ǘ��9��l�&�=ΓD?��X>Eƻ����md3��Z[���?y]?�?\�'�'�s�a?3%g�|Zv���,����О�>��2��J�F�v�
�/�b����1I���Y�?��?�5�?7���"�8+)?M��>�퐾�꾾8�j=Cx�>Y�>��c>�Zu��Dg>>���W2���>�.�?�!�?��?{=���J���!�=/E~?È�>�o�?@3>z?�$�=�s���[4=��>��	>dM���?�F?���>��c=
�2��+�F�J�J����B���>�(Z?'�H?�$]>�����^輦��B��r��%�����@����C���f>>�e>ur�=��i�s���?Lp�6�ؿ j��p'��54?(��>�?����t�%���;_?Oz�>�6��+���%���B�`��?�G�??�?��׾�R̼�>:�>�I�>:�Խ����`�����7>.�B?Q��D��t�o�w�>���?
�@�ծ?gi�o��>�/�rT��҇���;�U��'�=��>����,�=�9>��ؼ&�?��<����l�M��>o�?w��?�й>	7�?�lt�!��jG?>{s=9`5?tb%?�U>�������=�ӄ>�,ھꑿ=z��ܑm?�^	@��@P\>?&����[ٿxϐ��׾�3־��e<h>�<��
>�ռ���=`IE>h��=��<�`>��>��I>S&>��0>��h>W��>lˀ����je���U���.�֦��b�#��Xh��9�ؽ-����n�f��)�0�{m��g�轀�I�(KZ�̞��O�=B�U?P?,m?ҹ�>��ν�>OR׾:�=y���4>��>��5?��\?�?|s5="����`�|c{��s��#����>�p?>��>�(�>A��>C��6Q>#>�Do>[l�=k�='r[�l��;l*c>א�>j�>/�>uD<>��>�δ��0����h��w�F�˽� �?v����J�T1��>L��ǵ���X�=�b.?�>���=п��,H?�����&���+�G�>��0?A\W?~�>>	���T��C>F��c�j�6Y>� ��sl�e�)�KQ>j?�wc>�ݖ>�tA�VC>��,��F��֓>3�@?+�����q��Mp�>����>	!�>�[i=�"�cД��{`�Q��Q5y=�\*?��>�FػE�k�����^���x>3��>���=D��=�bD>r�����9<������=��=�ZR>\?�8>3�=r��>�#���Z��<�>&�2>;n1>��9?�t&?9�c���`�q��@9�Z�X>�b�>�7w>�=�W��:�=���>�0q>�/ټ��C�Zf���1��?[>H���:U�W�����=d,Ƚ�Q>r��=��yB���$<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ h�>�x�eZ�����M�u���#=���>�8H?�V����O��>��v
?�?_�۩����ȿ(|v����>E�?���?[�m�{A���@�u��>%��?~gY?oi>h۾�`Z�j��>ٻ@?�R?��>�9��'���?߶?֯�?��I>'<�?��r?���>�,��\/��ʲ�zM����z=M�;�>�� >֬��%�F��咿����Kk�uv�j�Y>q�=�ո>��m*��~Q�=���7ਾ;�R�F5�>s�q>O�K>�c�>��?.�>"�>Ռ=�Q��l���l{����K?,��?z��<n���<F��=5�^��,?�L4?z�X��aϾ�٨>T�\?�̀?6�Z?C�>����<��,࿿�����.�<��K>T3�>�H�>�ꇽ�]K>��Ծ�C�J�>)ї>Nݥ��(ھ"���j��2W�>�k!?(��>&Ѯ=� ?h�#?`�j>�*�>aE�I8���E�r��>9��>F?��~?��?�ӹ��X3�	��d硿��[�_FN>�x?�T?Gȕ>���Q�����E��bI�����D��?Zvg?;@��?�0�?�??�A?-0f>��Y	ؾ<ĭ�K�>l�-?���S�f������
;���>��>���>�M����4=�닽�e��D��?I�~?A�N?a���H b���uR�;R�&���%=;x=7,�q>��>bn�����=�o-> K�=Փ�����s?C=F�N>��>O
<�AC�����0?E�,�G���$u=�:~�
�J�b��>O�W>ݧ����U?=0�U��_㬿���
�F�S,�?�J�?}n�?���q�h�cR?*[�?�n?�{ ?�����fо�~ɾ�cW�����V� ��$�=W�>\٨� ���%���Y���-����ɽ�{���>��>]�?���>��C>��>�3��(���<�\Z[�Yc���6��-�����죾�x
������ڿ��"m�AG�>��|��]�>�\?E�Q>�̈́>�J�>mm�<明>�H@>{x�>^*�>ԋu>o/>ϋ�=���+���*R?sK����%�p=⾦^��	9A?`ae?=��>4,���6�����?���?���?��c>��j�/)��,	?M.?`�}�rc?h4==2��;U�;/���p���Hb�2�}��~�>�W���8���K�R�e� ?�?�����Ӿ���I����<=��?��?�����L�z�u��Y� �O���ƼEKo�*F���n�`o��_��L��5\����'����a�+?CK�?5w �_%������b��-<��\>5�>��>���>�<2>��Xn2��qY��T ��T��]<�>�?2�u>��Q?��H?�Z\?�$?�b�>ә�>�	���?}���?�,?�DG?�??� �>���>|�?c}>��{U�/�{�S"?� ?��8?0O[?��'?�>���(���7my�c���"��y����!�=>����6���t�=�#�>R�?W�׽�o-���߾5`Q>n8?q$�>z�>�x��-����@�����>��?%�>�����z�w���n?��? ��9V�<�X%>xz�=�B�uy��4�=���<;�>Q&=�  ��5<�'�=�d�= �=����o򈽵%<�=E�; ?L� ?�9H>P��>���f�X���Y�	/�������_���ֻ����s�b���Ǌ�+݀=&Ԟ?���?�+f>X�>��=�mE�lk׾⾶WǾ�֠=���>��.?}%h?e�U?�(�>�?^\�>GX�dꚿ�o~���[�*�&? !,?`��>�����ʾ�`�3�`�?�\?R9a�A��q=)�)�¾�սw�>�X/�%+~�w���D��ӄ����o|�����?���?�#A�y�6��n�����9e����C?r�>_[�>6�>u�)���g��'�$6;>ߎ�>v	R?���>@�O?��k?�HT?xWm=��h����u���=h`>Zm?R�|?x��?�k�?�\�>��=���ӣ��:���$~�<Q��`����=�|p>&|�>Gպ>.\�>t,>�s6�J�=5\����=�q>î�>My�>ot�>���>��3=%�G?1��>�e��(��WӤ�ǎ����<�>�u?r~�?NJ+?}�=����E��l��!S�>Fc�?�۫?�*?�@S�+��=�>׼���-q���>���>2�>�^�=XED=Պ>,��>!��><u��Y�2o8��N���?� F?���=X4п,v@�(���xѾ�z>!���XS���	��X�<=�g>��c�0���V�
����!ɴ������ɚ�gž?s�><�P>�c���~">�N�=�e_��8K�2�엝�v)��pB���C���@������=u'A=�O�=�%�=�4о.��?D`?�sL?�SB?�5�>̟�>*�1>@�>Ā���?g��>�%>�G����?����۾� �����ʥu�n ^���=����\>t�=C�:;�2�=��=E��=֖ս��4=�ݤ=f(�= e >b��=P�F=t�=� 
>���?s��ı�xT�v��<4�?̉S=|�->����ZU(?�c�Z1O��ȵ���޾�?�	�?z�?��>����>5Ȳ��Ku���>��&�&w>?��>KU=�m�>��>�x`�O�M���w����?m�?��A?�"��s3п�`�>�u7>�f>�2T��k2��O�Zof��N��0#?{�9�2KǾ_�>Bw=&��ކƾ��X={Q=>�9=�{#�&�X�}�=�}���?=��Z=�Q�>��M>�Ԗ=|6��\b�=��\=��=uV>,u��^I�T�뼲�V=�V�=�R_>�1&>A��>u�?Ua0?qWd?1'�>e"n��Ͼ�-���R�>\,�=_�>g��=ÆB>���>��7?��D?_�K?�w�>���=���>{	�>�,�i�m��b�1�����<H��?Ĭ?$Ǹ>��Q<ƟA�֜�b>�!MŽ�v?,S1?�p?�ޞ>�R�ޮݿ�S#��2.��p��#�5<��M=�{a�ƅ���Ǽ�H�!ƽ���=Y�>Ga�>y.�>$t>��4>2�I>�~�>%�>�X�< �\=��:�ʘ<�����V=.	輣8�<Z���O��:��<�]�\Ѽ�2�;7�<q<y�U;�"H>�2�>#��7��>7���޾f�>$~��)�n/M;���D8g�P>~�w�i�g
�#
J���=Y�=u�:뭔��<?->�n/=�R�?j?�C>D�Ϻ_���닿,ʾ�Ѧ��ō�[A=���Ŝ3�+�i��kQ�a���/�>^u�>2��>l#�>Y2��7��i�=���T�,�}I�>J�L\1�$c�S�h�9<��e�� �b�!�<F|<?n:��"��=��s?X�S??R�?��>�D���꿾��T>��Q���=�	� _b��C���8)?��3?���>A[	��1U��˾2m����>�D������燿�O�x�ڽ g¾�U�>Oߴ�mr��!��4��h؍�(�;�f�|���>^bI?���?�|�c�r�o�7�Ę�3#���V�>9?H?y�L>&5�>)W�>d��u.������#w�=�Kp?o��?N��?��(>���==)����>5�
?Ʈ�?&P�?0l?������>��<*>l�ݼbd>5�
>���=WT�=[��>�?�t?s.��3~	�,i�������m���7<D�D=�Fq>��{>�7�>cd>I�=��-=�}>#(�>8�>d> ܠ>�zv>j�s��*W�>x���͈s>��?!�=3ג>^��=�擽���u(��Z��!�O����=��u>G����Ͻ�=�S�>H2ѿ��?��>��%��?4��� s�RZ>�e��䀾ߓ,?��>b�>�O>Ϸ�>�%D>�Y�>��V>[>޾��=�Yᾕ[9�)��#�=��z
�nJ>�E��%����)�h���G���ԾS���`��-}��2�b�����?�,�mQY�84%�<����?[>�>:!?%��:5����=���>�4�>\��ٝ����z�o[Ⱦ8B�?s�?��e>8U�>��V?�?O3�v�+���W��u��C��+g��a�L���j �����@ɽȐ^?��x?OB?�!�<�y>()�?��%��팾k͋>��,��48�_�
=��>�����W�nξ�s¾����=>m?r�?�E?J	W���u��(�>��A?�?`v5?\I>?��?��1<:J,?z�>�K?��#?�&;?�I?��	?gR>)J2�����=�伽�R�����A7��Lѽ����C��V��j	���;�O�<��
�PȞ��j(=H��(�=�M#>8�2>I�>n�>&�Z?�|�>���>.�+?U֊�*��`Ѿt%�>	�˽����tG��٦� W�nc=��\?k�?�vh?um>m�;��)���>}��>fp(>a�K>`�>����?�Ε=��>�\�=���=�F��5������V[�tC�=�&>C~ ?6�>�����[>�[�����'�U>��	��ѻ�����9b�,e�𑾗�>�I*?�?d(�=��¾n�$=��2�5�H?�U)?4 ]?�'^?��5>�.���z�5ƍ��;�����>�6>ax���r���ꬿ�VV��H>��>d����!���=_>��	�I߾Ѻi�tI�kL���'=Z���M=����WӾ8:y����={4>Կ��, ��ǖ�R_��KI?Ɂ\=s~���#a��賾&�>l�>�٫>����a���?A�򿮾�+�={"�>�0>�������9F�`�d�>9vP?d9??�m�?��*��b���C�P���O��2N�Ħ3?Z4i>���>W)�>��r=/����1��!o�����>�n�>$��!����ҾeJ!�r�g�Ԗ�>i�>;
׽wWg?�Je?aڕ>��s?���>��>���>��b�r�۾h�%?���?�h�=Y�=�9��Zr^�8sQ��z?��$?�ߐ� �?Gw1?	��>�!A?l?�>hԂ>����C[��$V>�J;>G�7�2S���^�>�sR?v�?�]A?��?���>��r ��\=b��=��=ʧD?O�?>'d?nx�>l	�>`F�����=[�>��b?�3�?I�o? ��=7?��2>���>�<�=���>�R�>?�?�O?mys?��J?	i�>���<4:���(��r9u��CO����;PZL<0dx=�?�Ss����v�<y�;vӶ�H���R����1E�l���s�;-��>�Rr>����Y�0>��ľY���DA>
���I���&���#�:��ݶ=�M�>=K?4L�>�\"�^~�=:/�>,[�>���A(?/�?`�?��9��b���ھϿJ�x��>�A?���=dm�����a�u�يe=s�m?]�^?��V�Z�����b?��]?�f��=�6�þ#�b���S�O?��
?~�G�1�>��~?C�q?R��>U�e��:n�T���Cb���j��ɶ=Er�>�W�h�d��A�>j�7?MR�>/�b>$,�=rs۾��w��p���?��?5�?���?S)*>��n�4࿆�������1\?��>�O��6$?k,�.Ծ(���Ƣ�%-��K���b���z����#��h}�s�ͽ��=Н?��u?��o?U `?�O��ݺ`���[��	��"�Z�F������B�|%A���C��Wr�;�r��ڳ���[>=+�f�kn*�w��?��-?�/O���>��R��Gоu÷�Z�->,馾ͩ����=��6>K=p_���1��"�Y�H�����"?�'�>bw�>x'A?bp�ѬI�m>��`2��}꾌�>Yk�>EOJ>���>��=�>5���3�\��֒�:�R����>��[?��@?kx?S�[��n��x�����z���Dc����>�FR=��W>�ܩ��\O�#�8�^�M�C�u������v��#=��?E�>��>��?�?`&׾����=�(���D>&N�>�Oy?�q�>�aP>��ۼy(:�FP�>B�g?+��>P��>��Ծ=t��À��B���|>�>>7�>?W>"Ԥ�?;n������*��
j4���=/)}?!�����w��l�>��H?�¼��f���p>C�������/�����`#�=ؤ�>1 �<B�]>å��v��.���'X�}I)?�E?"Ⓘ}�*�7?~>�&"?+��>.�>�.�?�2�>�mþ��F�-�?��^?�=J?%LA?�2�>r�=�ʱ�K9Ƚϼ&���,=8}�>�Z>�{m=W��=����e\��t�i�D=�r�=PμV8���z<Le����K<t�<T�3>�}ۿ,!K�bFؾ���@�D
��҈�JU������h�#볾˘�Ts��;���"�uT�ʴb��_���Wn�')�?;�?v���[$��L��`������r�>Hsp���Mū�{��󃔾RP�}t����!��N��5h��^e�K�'?�����ǿ󰡿�:ܾ&! ?�A ?B�y?��1�"���8�ĭ >A�<%-����뾡�����ο>�����^?���>��$/��c��>���>�X>�Hq>���r螾�.�<��?C�-?��>��r�%�ɿZ���"Ĥ<���?.�@_A?n�'�n�� �^=�$�>ܐ
?�>>�5���U��M�>Ѿ�?�g�?��:=�:X�DV���e?X�A< 0F��uȻ���=`��=0=���<JI>\E�>[��@�F��ܽ�4>:Յ>������<Le�u��<^�\>:�ͽ�����i�?s�o����^���,���f��hF?`��>�X���?)�$���̿b^�沁?�@�?���?k=?���57�>4辉�t?QO?��k>}=I�/ބ���=�\��!������%�h����>8�c\[����"�Ӿ��.=��=�ꟼ���,��s��	��H=g��c��`���==ǩ(>�p̽����)�=[��=�]1>@ٓ>��4>�z8=S��=�n]?�2�?�P?ʼ�>\;�5ȾP\��;4��В½�1�&���P�����ɻ<N��u�쾲�%��Ӿ-���SW�f�;��R�=�rR��W����,�b��E���.?�>'ʾ�_N�?H�:,v;�ث�*Sj�;S��s̾d�1��m���?��A?!셿X�_��(��@Y���=X?���.��.�����=�r���{=�ߜ>��=���W2�';R�.\0?Ғ?�׾�sA���T(>����=��+?�?�$U<̪�>'=%?�K*��߽PhY>3B2>ri�>���>�x>�$���cܽ~�?�$T?²��#!���B�>����1y���m=, >��8��tڼ�u[>��<3����`��È����< (W?���>��)�~��b���#�DL==v�x?~�?�+�>�}k?n�B?�<`_���S����w=��W?g%i?��>����)о���x�5?��e?��N>�_h����a�.�rT��?��n?]^? ����s}��������n6?��v?s^�vs�����U�V�o=�>�[�>���>��9��k�>�>?�#��G�� ���|Y4�"Þ?��@���?��;<��q��=�;?n\�> �O��>ƾ�z�������q=�"�>���zev����R,�_�8?٠�?���>������a�=ً��F̫?U �?s-����<�`�_l�ǌ ��[[<d�=����%����7��hǾP
��ݛ���Ǽa�>�%@�R�F�>��:����f�ο{Յ���Ӿ��s�`3?���>Xý�ࢾ3�k��"v���F�G H�p������>�>�`���K���pu�b�;�3$,����>d���>��^�A2���T��w�{�i=�>�7�>�W�>u_��	/���I�?����\Ͽ}����7	�swX?�J�?�x�?iA?�;�<g�r��t�����P�G?�x?��]?�G�W'l�o��9�j?�"��.;`��d4��TE�x2U>� 3?S�>��-���y=��>vy�>��>�3/��Ŀq۶�!������?N��?Vb�U��>�y�?{{+?�j��E������Ţ*����8�ZA?i�2>A~����!�a=�l͒�Ŗ
?�N0?���8��~?�B�����������O�=A�=>s<9�;��s���d�<y�K�F�K��䗾ퟒ?o:�?i9�?v'������\?;�>-谾۠���l>�`$>m/�>�J�>�>Ͻ *�>Eu��f���q>�J�?B��?���>����J��u3�=�Q�?���>ք?���=A�>��=F��:��[o)>dF�=W
!�G`?�/M?6B�>��=�L;��.�)�F���P�Q����B�%��>nH`?�TJ?�6b>4��e�9��l!��}ʽ��/��Vؼ�5���1��h�$�6>� ?>w�>��I���Ӿj�?�n��ؿ�m��P"'��$4?���>��?I����t��/��-_?�n�>j<��.��� ���$�̙�?�B�?]�?��׾i+ͼs�>��>nA�>}9ս�ߟ�����a�7>��B?�)��@���o�q�>���?��@�ܮ?4i����>�&��z��ˏ�+�Q��d��PH�D߽>����r=\�>������`��>��������>���?���?��>�Ã?�_��LX��O=VAW>�X?���>i�?>&���3�=���>�t�ù������ռ�?M�@��@M�e?	��fܿ��̪�n&��+=*�=�)�>Cཤ��=tuW>�ȏ�69W���;>��I>AQz>J2�>��;>gs$>�vG>���fu�	֟�d�����8�����i	�<2T�����:���ľM젾ZL۾�I��Y<���=!�e�2j)�$Cx��l�=��U?2�S?��p?a# ?�J�U�'>4����=O��m��=�Z�>�e3?LK?��'?��=�ܡ��|c��B�������ք�6�>�R<>�/�>�b�>��>� �9�N>��;>�uw>�>4*=�|"���=�'R>�$�>i��>���>Qd<>��>�δ�))��;eh�oIw�y�˽��?�ǝ�ȖJ��8��G捾H�����=l.?��>���.пn୿��G?�Ɣ�%���,��>��0?W?�h>zҰ���R�5�>���Dj�{�>.���8l�Mx)�=Q>�f?R�u>�r�>KS�b]N�����ž>�/>0�`?m�����޽�����*&��,�=\�>���=�������Q�)���c�r=g)?�F^>��ǁv� ������X��>�$>�,��l�/>@��>��=�p<(O߽���=q�+>��>?~eB>J��=ѕ�>Ok���u9��?�>oc>Y�;>��>?��)?B�C�ɊX�M�e��lC���e>l��>dG�>��=^cQ��s�=g�>��q>3C��	����R$/��@H>I51�/�q�*���=GR��N`�=�Z�=����0B��a=���?3���Mq��i޾�|���l9?��	?Ɯ�=9I�;c��`���㬾5�?	i@!Ԝ?a����T���?:�?�X����>��>U��>
޾�AA�=�?/悔�ϣ��X���(�pm�?Ao�?��=I!���-g�I#>��?�־Ph�>{x��Z�������u�v�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?��m>���?��d?z�?b�S���#����?��n�{��\���u>�"�=p���k�`�����-��[nl�j�)��{�>|X�;���> F��&��:!>驇<������,�E��>K.�>��=��=>y?�>ZN�>nU�=�g�t����m;k�K?���?����1n�:�<��=ܴ^�'?mI4?��[���Ͼ�֨>^�\?�? [?�b�>���+>��F迿!~��3��<C�K>P3�>�I�>� ��LIK>
�ԾM2D��q�>З><���>ھ�,���}��+C�>�e!?���>]Ԯ=6� ?\�#?j>�J�>mE�Z3��o�E�8��>�l�>,*?��~?��?����e3�[���롿q�[��IN>Qy?�G?n��>ނ���s���kG��J��E�����?-}g?[Y��
?s&�? q??�A?�,f>l��$ؾɘ�����>/<?z精-:e�x�lP��(k�>�b�>���>od�hV��[i½_1��sо<?��x?`�&?C��(Q������<��=a3��L��T��Ay�=k+!>���<t�9gy�=���=����.x��,l=(�=:�>�j=>]	l�&Yz��H2?żn�����=�t��~S��D�>Y�A>��Ͼ��L?p�F��Ǉ��Ȱ�`�$%!�5��?�m�?dF�?z�E�|m�=2K?M��??��?�Y��k7о⾯N�����Ư��:>�x�>Ͱ*��4�!;��w���͂�B��M����d?���>A�?���>U��>�@�>�w�ٟ ��8־][	���\���E�A�_��0�&����R>��f���־A<���>�	2�E��>e� ?0�>�{�>�;�>B*E<�%>�>N
�>��>6�>�x�>|m>	��=��ҽ\�R?�@þƩ(�'&�ӯ�&�A?�d?���>��l�����?6�?�Ȝ?��z>B[g��+���?  ?���_�
?�9=�H)�T�Y<�Y��D��>ソ�=��ȍ>plսj:��M���d��,
?�?`+v���̾�I�{��o�<JX{?V)?y���i�P��v��l��3��:��,����ۍ�[z���q��!���<z���t��/��/�3*/?�u?vT�����g�$f���5�|]>���>�g>�`�>O~�=���R'��f�|���I]����>��?1��>(=U?��A?C�_?V�?M5�>Y�>e��}?i!�=�?��>5?,�G?�Z�>
��>�?�K�>�5W�^��_ž�F?)�?�7+?�=?{T#?C�������t)>��[���ƾ�>���<�����z��.�=�W�>P�?�����8��C���*k>u:7?���>���>ُ�����]x�<���>��
?�"�>6����
r�	z���>ւ? F�M�=�B)>�#�=�V��s^�B�=����q�=Ƞ��S�<���<w��=�̙=pG���d�sG;��B;�[�<�P?z�,?��u>�ʿ>��ݾ��0�R@�;j-�%��1K��/o���E����~��+��I'��e ��ҋ?��?L�K>H�=�D=>�12����]� ��*��q�_?SM0?��o?��?X ?k!�>���=N�!�������T���
�&?A!,?<��>���J�ʾy񨿻�3�U�?�[?,<a����<)�ő¾�ս�>�Z/��.~�T���D�l���\��d�����?���?�#A���6��x辽����Y��F�C?"�>Z�>��>�)���g�4%��2;>��>vR?��>�oQ?�/y?N�\?<>*�<�y����C��%Y��>� D?4��?���?Az?{��>�>B�"�y���d �����������dLC=�j>�x�>^h�>i��>m��=/�-���^2�w��=ISc>9p�>���>�w�>K��>���<��B?DU�>j�;�������|���Zن�
%}?�~�?�?z/�2x��4O�E������>n=�?Y}�?��%?w�e��=���������_J��E�>��>݃�>���;S��=N@j=���>���>��������.�QT��O?�~F?ɇ�=�C��P�(���*=����D�M>#f���Dپ]1ԾD�����:>��6�|��=�˓<����^��qΉ�0�r���Ǿ_CԾ%j?�3�<K�g=���|�g>5�]����Xbҽ���(�L�&���4�����%Wv��i��T����B������<�����y?4[Y?l�4?�~'?�ҩ>�Y�>���=�.�>ǋY=j
?�8�>�H�=�*��x��/�����׾-�I�⾌�h��7f���=n&�ղ�=!���[>�.b=�n>�F<1㦽�Xp=����=>>�!>))>��=0>sx?m8��������o����=��?ļQ�+K=�	Ѿ!� ?1�Ot�X鲿nI���t?k @y�?�� ?��B��p�>^x��,۾N��>Q�m�çl>rK�>$u8>���>p��>.�ɾYY���p��i�?5�@�O`?5Ч���Կ���>�h8>{�>�S��2��JW��)e�7[���#?t�;��ɾ�L}>�h�=���e�ž>�O=��9>%�U=dB�gZ����=�{��}A=��H=�ʆ>�C>���=:q��>u�=X3=Z�=�dU>��Ⱥ�)�z��il==�d�=��e>�2/>Ҙ�>�?�W0?�Vd?���>dtn�}!Ͼ����'n�>���=q��>�i�=�jB>%��>��7?җD?��K?I��>���=:�>t�>`�,�T�m�g�&r��X9�<���?�ˆ?��>��Q<`.B��z�T>��{Ž|?�>1?��?=�>���.�ῦ�*���:��ͽ�00=�^�=�k��4��a�=���u�r����=���>TC�>n��>�X>��&> 9S> ��>��>{>zl>{5�<@0�<}��:ٝ=��8<��F=�@>1��=KKa�/ �<���PR-<Q(o�=��*���Z=>���>"z�;?�>��Z=ټ�^>Ja��>Y�m1�<E?Ͼ��f�	���&�u�|��F�ӽO�8>U�>�b�������?)��=���=Q��?]Gy?	Q�=�P(<[�Ծ�ك��¾%�J����=�蟻6����7�v�s���O��#뾊�>���>�
�>�\s>=�,��=�~^=�)�c�5�/��>5���c+�?���@r����j4���i�9r�ehD?�臿)��=[m|?��G?�͏?��>�W��vEվ��2>s ~����<���C�e�cz���??�8'?��>��V�E���Ͼ7�ɱ�>�;ƾM���r̕��aB�0�������c> �;-�ھ�)�n!��P���_�0�-}C���>:E?J��?Z�������T��|��O�.�>��G?[M4>���>7z�>x`$��\ ��(��k�=�u?�X�?cJ�?��\>�K�=}�����>r]	?x��?뱑?g�s?�=����>ޤ�;��!>Hژ�m��=�>-�=B��=?n�
?�
?�۝�G�	�"'��~�EV]���<lա=.1�>X�>s�r>|��= Qj=?_�=_�[>���>"��>-4d>O�>��>�q���o���� ?#���P>!�?|�;>s�A>H�5<�ؽM�h�<���Gq��'���!b=��=*��=Eܴ=��	>ȟ�>Pʿa��?ߤ>�\&�(?<V۾�i���Ҕ>���0x�;� ?��X>��>sa�>ˍ�>�w[>Om�>��!>4�־3�>�}	�J~%���6���R�E۾�`K>���.��W
�����C��7��:��P�f�� ��@t>�u<��?�l��Ro�O�.�g�ν�t?��>]	.?�D���[����	>Ϫ�>+s>����3X��;����ؾ��?���?h�o>���>�nP?u?_S�Ou̽��T�^[|�L�P��u�=`b�/����Y�����~����U?�Pz?�C?�|�<z{>�_�?�1�g�n�D��>�R&��1�U��<XiV>lh��g�]�����@ۭ�;/�T�=�(V?�@�?~�?�EJ���B�<f�>V�P?.w�>:9?S8a?��j?��0=�xW?�?"��>vH)?*X?�?�]�>�+�<��Q���B>��������j���\�(�\��>|<���=<�=ݜU��3�'�<G�g�R��=R:����J�7=�<)=v��=�}5<b~Y=GŦ>��]?�D�>��>�7?<���l8�0���E/?�8=�|����������񾏫>��j?E��?
fZ?~!d>p�A�o�B�9H>Y�>d�&>qU\>~��>qa�ՍE�i�=�1>,	>04�=�M�8���ݿ	����a��<(G>���>f��=w���b��=j��߅	�6+>J𕾽=������O�>@.�7jž��:>�wH?�?�sv>�����d&=Q�6��!2?�??��?!^A?HW�>����@}�bې�|������>*�>�Վ�u@��P���NG�C����>d�̾�ݠ�NZb> ��\u޾��n�NJ�f��KM=�~�kYV=���վ�2���=A$
>������ �W��ת�1J?Ҥj=x���bU��o����>���>V�>�:���v�ǈ@�񯬾�4�=d��>_;>2_��R���~G�d8�i#�>��E?;\O?�͙?��f�\�}�1+&����R���sA!�� ??�>��	?�1>4*���ƾ̱�7&`�y� �/��>\i�>��$?��P ��"��d6��7>KQ?�L}>=:?��?d�*?�x_?"�!?H��>��s>�����4���B&?y��?��=��ԽU�T�U�8��F� �>v�)?ڷB�/��>4�?��?�&?{�Q?̳?��>�� �nE@����>cX�>�W�$b��j�_>��J?͜�>_=Y?<ԃ?�=>d�5��颾}ש�I[�=;>��2?@6#?,�?��>���>�����j�=̲�>�c?�-�?��o?ms�=��?92>���>j��=�ȟ>���>� ?iBO?Q�s?��J?�j�>�f�<� ���z��r��gJ�%�;=/F<C�x=�����s��j�a�<e�;����P����t�GE�F;����;�_�>q�s>8
��|�0>w�ľ�P���@>_���P��ۊ�o�:�hڷ=���>��?7��>�Y#����=l��>YI�>���6(?��?!?��!;ϡb�`�ھձK�8�>2	B?���=��l�'���-�u���g=��m?G�^?[�W��&����n?@{~?h�ݾK#;��*��厾��+���1?(5?�f�o��>H�w?�8w?%�?i^J�ȁ�R���xd��3�Ѿ��>���>(��\؉�Vݝ>�
[?���>O�>`8>x���������|�?b6�?���?Uk?T�>4�s�8�������䎿taj?_b�>YW��t	,?y�Q��F �����ɾ1�
��D����Ӿ�t��gᶾ/���F�o%�X�D<U
?ז�?�S?(�?P�
�g-q�L�3�󽚿�G�w��8�D�i0t�8B�+3�@9m�b�LB���Ծ�S=J�|��A����?�n'?�N/���>���1���uξX>>�ա��w�%M�=����c�-=��a=�De�.�����X�?�&�>\�>#W>?�e[�rV>��0���9�`����.>`a�>p�>"p�>���:{�.�����Ⱦ�ۅ�,<ѽ�t>i�c?8?5��?<}s��9�4i�����F���Ծ9z,>F��<��d>�GC�)�W�Ы1�ۯE���i�ѡ徛$|�"��y=�kP?���>'W[>���?��?	B.�sy���.��8O2��p�=��>�T?W�?D>�Z�m_'�c��>�s?k��>��>/\q���kH��M�-�R��>�L>>�>�}�=��=�¬=�-����)���-#�$��=Փr?�i>�5r��>G�?d�=Z�q�?Yq�=�)����Q�bX�<��?�و>1,>����{@��T���S��S)?�[?e����i*�MC~>`�!?�#�>��>�1�?�F�>$�þ�g����?��^?�ZJ?�A?��>m='��v�Ƚ�3'�!�/=Uʇ>��Z>7rl=G��=�� .\�]��&�H=/��=�м��<����9L<���<�H4>��ڿ0�K��k̾+��h���
��蓾Z���i��q
&���R���'�o�����6��ya��0s�9����{�]l�?~�?p�t��m��ؙ��^�����N�>4�R����b��]�C�^�����쾳ӿ���9UU�Uj�	P^�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�|A?��(����KV=���>c�	?��?>�V1�~J����yT�><�?_��?�lM=��W�t�	��e?,�<	�F���ݻO�=;D�=dG=���%�J>�U�>��RTA��=ܽ$�4>lۅ>�{"���Q�^�
z�<Ї]>�ս78��Մ?�N\��Lf�J�/��n��P>�3U?)L�>c�=v-?��G�%�Ͽk�\�{�`?���?F��?�)?T������>��ܾ/�M?!{6? �>��&�tu�@F�=�E׼C�b���㾗\V����=o��>�z>N�*�H���P�(˗�E�=0b�=ƿ�������<@��;P#ǽ��
��<m��@���"��j�B��Ͻ���=�4>�.>�s>"�->2.>�R?��r?���>��I>� �]��.!ȾМ���8���`�<����:u��e��ؾ�!	�������_��!=���=7R�n���F� �m�b�Y�F���.?w$>b�ʾ��M�8�-<�pʾ^����ۄ�᥽�-̾�1�)"n�n͟?��A?������V�X���W�����Y�W?+P�ֻ��ꬾ���=a���t�=%�>̊�=���� 3��~S��w0?�h?C\���8���*>�G��=��+?}�?�^<)�>I%?�U*���$�[>�J3>���>V�>K�>����ܽ��?��T?�������Ɛ>�U���z��]_=7�>4���Z[>x�<�猾D�W��)����<(W?���>�)�~��a��\��jC==[�x?̒?*-�>�zk?�B?ZȤ<�h����S�/ ��fw=�W?�)i?C�>Έ��\о���޿5?�e?�N>�ah������.��T�X$?�n?�_?���xw}�������Bo6?��?��_�Gƿz&$�sԾb�?��o?zL�>�W����"?s�Y?��������2�����Q����?>I @��?�?����o>*�?���>�����F���Q�iݏ���>%�?9'��� S���\�_-оȅ?_8�?� �>j����A��=7���M�?�ʇ?+���@ =���"#r���O��:��:=��K�uuT�6�^9����X�I1��Q��;'�>+@>A�n��>�8�c�⿃�̿ʈ��|Ӿ<����?⢜>ⅻ�������e��Tq���B��F��Ԇ�9L�>B�>/�������8�{��r;�#D���>:�,	�>��S�*������`5<��>���>R��>+��v佾�ř?�f��Aοy������ܽX?�h�?bo�?go?�@:<|�v��{�щ��.G?��s?�Z?]V%��*]���7�%�j?�_��yU`���4�uHE��U>�"3?�B�>U�-�i�|=�>���>g>�#/�y�Ŀ�ٶ�<���Z��?��?�o���>r��?ts+?�i�8���[����*�
�+��<A?�2>���J�!�D0=�SҒ�ü
?V~0?{�e.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�I�>�?P�=&��>�]�=�ʲ� ]�T>(>�B>�4�Ա?�=M?���>eY�=��2���.�#"F�ִR�Ğ���B��׃>�@b?�#L?W$b>�����'�I" ��Mν�;4������7��v7��~Ὥ�2>Q�<>K*>�B��Ͼ_!?�|%�7ݿ��"�]��C?nٯ>��?���|����=�YB?�B�>{
��黿C�����X#�?\��?,?D�׾������=@��>�G�>��賤�����>�6?'̕������s�|�Q>���?Q�	@u/�?��a�֑?���"��칃�h�v��?�r>j�6?���}�>�r?��H9�f� d��`���vP�>\�?wG�?���>2�m?�rc���F���=�ɴ>�n?e�?Ȉ<��%�=�	>���>���4���7~�Y�M?�@�@�^?]����ۿ��U������s'>�L���=�J�9Թ>���=V�<��]=��>=��>XF�=� $>�>��">�J>���������"8����A����V�z�<�����bo����\�����8�܊q= B+��<��V��t���I˽ɚ�>��6?P�Q?x�R? ��>f�l��m�=�g��ˡ>�������=�+?ru6?A_?��W?lB�!پ+�_��+i���3��^&�>9PA>���>m��>�8�>��?�	YR=�b�<��>�t>�Լ��}R�=�(k>"�>4Y�>��>^D<>�>(ϴ��1��x�h�W
w��̽&�?�����J��1��b9��&����k�=<b.?�z>���?п����w2H?+���k)�#�+�7�>o�0?�cW?��>$��W�T��8>u���j�v`>�* ��~l�d�)�\%Q>>l?�g>$�u>6�3�_8��P�0���(|>�?6?�����8�d�u���H��ݾ��M>��>�5H��l��������i���z=�z:?��?>���%����u��-���UR>��[>��=%	�=�iM>˃d�"ǽa�G�au.=�/�=��^>YT?�,>�ʎ=��>�I���P����>��B>�,>��??8&%?r�\Ɨ�#|���
.�a�v>Z'�>f��>�l>�BJ�ǯ=�m�>W�a>���ჽn��)�?�3)W>G�|�-_�5It�LDz=6��C��=�K�=0} ��=���%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿק�>h~Z��o���@���W��0	&=�3�>�I?.f�7��=���ő>8��>�پ���h���5o�eV?Ր�?&�?JQ�� ����U�^��>���?X��?�!�>�����x��kf>)�=?��`?��>P�%�gt����N?��?J�j?�SI>?�?2Zr?��>��g��J0�%����P��q=/����<�>X.�=�P���E����������j�Y����d>�j*=�>Nܽc����$�=l���9⦾�zp���>�y>��P>���>�^?�!�>�ԗ>u�=(!�����Z��XAZ?>�?����w�nY���T=�=x�6W+?b[?)��>U�V�_ �>U&f?B�?�mc?�?����
��M���oϿ���������1z>�	?A�?�B�'�q>WJn�o�I��>�:�>��v�-��_����5�= ��>���>'��>š�>�#?`�0?}�L>��?��R��h��@�I�`D�>��>�?��?mh)?B	Y��a�g5��T5��0~f�r)�=��r?EZ0?�Z�>hш�����(��/����/�i?b-�?�[ҽ��>M�?�}7?��U?�L�>Wf�� ־�+?��p�=��!?B�ҹA�EM&�C�F}?yP?���>0/����սnRּo��+}��� ?�)\?v@&?;��D,a�� þ�1�<v�"��U���;hD���>��>����=`>�ܰ=�Nm�VG6�c�f<�q�=m��>*�=�+7�Gs��l0?jp�<o,��ꪼ����BjJ�(	�>/T�>�"辆a�?��G�8|���m��p��1(���/�?�ֵ?�Q�?tc>�2v��XO?�B�?��?NF�>�.���+3��Y��q�.<�k���,�hs3>�`�>��#�(����^��D����8v���ᾛy�AK�>B�>�
?5�?p�;>��>�T����:�d��[Wھ/lV�i�.�C��z3�a�2�����q���c㱾�U����>��V�c,�>��
?x#|>A>p�>,Z�<@u>dT�>A{�>[7�>x$k>I��=]�>m���b����KR?����!�'��������d3B?�qd?U1�>5i�:��������?���?Ts�?%=v>
h��,+�{n?�>�>G��Tq
?uT:=9�N;�<V��j��3��3�3��>E׽� :��M�=nf�yj
?�/?�����̾�;׽�Kξr��=� ?��&?��1���m���t�j�g��OE�X*���C���Ҿ�����]��V����{�i����7��{��1�D?�t�?���G.׾�7쾏]g���0�6ߕ>DE�>��>���>��}�Wh��F�'Ձ�9���壾�q�>��?h$�>A?l�??R�M?a�R?�ԣ>�s�>�8��O+�>j ���b�>k�?�:?��.?�9?��?��?̎;>��������ӾZ ?De?��'?�?���>��Z�hX��aJ�'���|�d�����d;�:?н�#���=��X>�X?}����8�D����k>^�7?��>���>���'-����<��> �
?G�>' �~r�	c��V�>���?�����=��)>���=��6�ҺtZ�=�����=a3��y;��i<ɂ�=���=8Et�=ـ�6�:|��;"n�<��>��A?�¥>�����sj���ξq�(��9�ܣr>�k¼��r�Ǟ�T���җ�K�S��W@>y��?ի?�y�=�ޘ=
�=DỾ����*�	�럥�3EV��:?{�:?ysQ?�H�?�gB?��K? �k>UL/��O��iӖ������ ?o!,? ��>���0�ʾ���3�؝?f[?�<a�<���;)���¾��Խʱ>�[/�`/~����<D��酻���l��)��?违?tA�O�6��x�ҿ���[����C?'"�>AY�>��>C�)�n�g�]%��1;>ߊ�>_R?�E�>��O?L:{?}�[?Z�T>.�8�.���j���D:"���!>��??���?E�?r"y?���>ab>2w*��A�p���:�&+��������V=32Z>d��>>�>��>�r�=1TȽ�U�>�K��=��b>X��>Pť>���>��w>�٭<C�G?��>C\������뤾MŃ��=�u?���?��+?J=�����E�SH��RJ�>Yo�?!��?]4*?�S���=��ּ�ⶾl�q�1%�>�ڹ>�1�>�Ǔ=2�F=�c>~�>ؠ�>Q%�a��q8��VM��?hF?��=�}ƿ7�r�ާq�fS���rV<z#��x�f������Y�h��=_����v��&��|�W�|��'��s��6圾�Y|�Ǣ�>��=��=�<�=��<�XǼ��<��D=��<J�=�k�s�g<�u<��״��ɂ���2�EsS<\XI=(���T˾5�}?�2I?�+?�C?�)y>�)>G2�@��>R���-?�V>O�O��Q���e;������I��Z�ؾ�_׾��c�a⟾�>�,H���>��2>b��=�χ<��=N6s=֨�=�2@���=�&�=�r�=0ݬ=���=��>�N>A]w?dw���!��	?Q�N�ｑ;?�W�>��=��Ⱦ�EA?�B>Q��s���J+��~?]v�?�P�?t�?߉^��r�>TQ��|�����=�綠->'��=1��H�>��K>6��*6������Т�?%o@5??�ً�.�ο�#->$�7>�P>��R���1��\��Vb�qnZ��]!?�l;���̾�N�>�ƺ=wC߾��ƾW�,=7�6>rIb=���^\��ƙ=�|�{|>=�k=	�>=D>G޺=����Yŵ=�<I=�!�=$�P>
���^�5��+��42=���=Kwb>M&>͐�>{�?�c0?�Wd?�4�>Fn��Ͼ?G���D�>@��=�;�>Ҽ�=�WB>Ն�>I�7?n�D?*�K?���>�Ή=��>5�>L�,���m��h�>ǧ����<效?�Ά?�ָ>�5R<��A����f>��4Ž�t?�R1?vk?G��>���.�ٿ�84+��hɽ��o�NRj�	ǣ�1�<�xQ>����ݓ#>p��>���>�ע>��>�|{<x��Te���~�>,D>���:�ׄ�⼅�<n�=pE����<y��&L�<sݽ�[NнA�(���=	2ȼv�=F5�x���ȹ=���>u�Ὕ�_>��b=�ݬ�B��=/�{��X�a�<`� �d5N�Snt�_����0�E�:�vyf>{m�>˖�������>�3>�
>Yi�?`y?�I<����;�*������E��P�;ӗh>wau=Z�ӾH"=��PQ��dM�ZE� ��> ��>��>��l>,�e#?���w=>��a5�j�>i|��?��[)�R9q� @������qi��Һ�D?;F�����=�!~?��I?7�?���>�����ؾ�50>�H���=S�_(q�uf����?F'?���>D쾨�D�}<оh�����>��#�I�b��'��1�7��r������=��>��Y�R
�)j4��΁�QΖ���=�Tر�L#�>\�N?�̸?�ר��9����X�7�鸦=23?qp�?=�g>�+???/������7�� »�]?�C�?o��?�>���=����?�>�+	?���?}��?y�s?�l?��{�>�;�� >����Jg�=<�>窜=5%�={o?��
?E�
?q����	�Q��&��	^�O��<5֡=���>�j�>�r>���=.g=���=�'\>�Ӟ>��>��d>��>�N�>̓�K�	�rE?d��h1�>#�L?,g>��;��ھ>L����\�4��t���0���=���#=�_�=��=Qx�����>�ϿM��?V>w(���?6�žI�q>Sv�>cu�>����54�>��<��>�1�>��>vt>ו>���>�־x�>C���&��-G�8X�x�ھ=%e>{U����2��� ��@ �ET�t���"��PIh�������=�E�<�ϒ?}���s��+�g����	?��>��=?]����^��+>���>��|>H���X����;پ�=�?�h�?g�n>�)�>șh?�4D?�"� lS���=�=����,T����h����8��^Е��w%�����PZ?���?�3?o>��>�x�?6�����B�i>��,��4�[>�y�>�}����<C�ʾÞ���G�Ѕ�>z"N?��?[=?��U��v=+�e��f9?��#?�A�?�zD?�@7?y��>�?���=��?j�H?�V?Δ.?�K@?���<+�;��o���=�5�:�g�4��b���Y��;���N�=𾱽�� = �Q=�G��"�����3����������n3��0�=��=�>�Pf?2P
?Ѱ�>|�+?�-�+6��T��?&�������%������|�>n?�`�?�'a?+5�>��<�t:�,͗=��>c�>,f>���>tݽ�ئ���>�>�j,>�a>�����Ǔ�Nj�G�l�B=Nͼ=y��>=|>RM��3�'>>����Fz�]�d>��Q��κ���S��G�*�1�˫v�Z1�>�K?f�?_=�D龖#���Kf�./)?SS<?wEM?;�?PQ�=��۾��9���J����Q-�>ҝ�<���U¢��'����:�긒:H�s>�?��lޠ�59b>u���,޾/�n��J�û�u)L=1����T=!��վm-�B��=N�	>������ � ���Ī�JJ?,�i={����T�A���>�>���>?	<���v��v@�����2n�=	��>��:>��?�[�G��0��;�>�IE?�Q_?h�?\��s���B�����HK����Ǽ��?�~�>�i?�-B>�ǭ=Т��M ���d��G���>��>2����G��<��u"��=�$��w�>�;?d�>��?�R?��
?8�`?g*?�:?U�>����績�F&?���?�E�=OԽT���8���E�U[�>��)?�B�X��>J�?a�?��&?tHQ?�G?]>׃ ��J@�ڀ�>��>T�W�B.����_>tJ?&n�>pGY?���?d�>>�!5����6:�����=�G>z�2?43#?��?�*�>O��>m�����=T��>�c?�/�?	�o?���=F�?C2>?��>Q�=X��>���>�?�TO?b�s?s�J?��>���<';���:���Js�k�O��?�;�.H<}�y=d���t�^3����<��;�D��/���b�D�Cސ��C�;���>�gt>�ƕ��	1>�ľ�����A>w ������\����":�6��=���>U?K��>C$��~�=���>i��>����'?��?5�?%�:=�b��۾��J����>�A?S��=��l��n����u�.Dh=��m?̅^?ôV�������?@y|?�i�����~.�Z|>�g��v,?��+?7���t~�>"6n?���?@�>�g־ក�b��������ơ=֮�==³>����Z�@��>�F?- ?�;�=�v�<ͱ��K!��?�Ͼ{s�>r�x?�s�?�? S>OgR�P����\�@����*D?�Z�>d~Ծ�+C?��=�~���^��7�پ�b�����{�پ�2���-��i_� �2�w<l�?-�t?�!t?Ex�?���6�`��B�Q���jIB�?
�d6�j�K��� ��/��C}�S��Ҋ�	zb�+ޠ=�̀��?�,7�?��(?K7����>I�����DѾ��.>�٤�Kb�j�=�𙽼@ =TGF=��b�/�+�;n��	C?߷>{��>TA?2W���?��*�C6��D���V+>�*�>>���>��p<��/�4���Ծk� i��~Ot>I�a?��J?�no?$����v1��ꁿ�P!���H��A���*;>l�	>ꩉ>��V�]�!�LT&��o>���r�����;����	�d{}=��2?B3�>I1�>�A�?n�?�
�ӕ��eu��1�G��<ﲴ>�%f?�*�>2+�>�1�T; ��Ƶ>�U?(.�>��>����1� ��>t�׌!�׏�>\g>�j�>�cN>���xE�抿z]���0�,g�=�i`?"c�IY��x>�]?F  =ub~�9��> �= .���ھ5���=)`-?���=���=�����;�7���?�z�s�(?�t?����Z�'�&|>|n?|X�>��>�a�?��>�3fU<��?��_?�H?ʞ<?���>d$4=�b���pǽc�(��'=`n�>��\>"�}=��=Y���X����_i=��=k#��Pü����;�7��~<�~ =t�5>�lۿLBK��پ�	��?
�{舾b����d������b��2���Xx����	'�+V��6c�j���9�l���?�<�?7���P-����������������>�q�%�������%%��}������d!�}�O��'i�d�e�P�'?�����ǿ𰡿�:ܾ3! ?�A ?8�y?��6�"���8�&� >�C�<�,����뾭����ο?�����^?���>��/��o��>ߥ�>�X>�Hq>����螾�1�<��?5�-?��>ӎr�0�ɿ`����¤<���?/�@�|A?��(�,��1%V=N��>��	?��?>�%1�<�<����J�>�;�?_��?/�M=��W�Ch
�xte?��<��F�ݻ���=��=�`=P��`�J>�Q�>�T�pFA�Uܽ��4>�Յ>��"�V���^�eǾ<)�]>Rbս(Ҕ��m}?Ƶ����~���;������x=Wu�?��>{>=ɧD?���8տ�bq���?��?���?7�;?�
K��>�z�˽w?rD?�5�>:;��n��-n�<�i�M�h��������G=���>�aQ�]G�=�/����'�=�ρ<s�G�ƿ�%��o��8=��J���W���潱����W�@r��&.p����imd='<�=��Q>�L�>?W>�NY>�2W?�}k?׍�>�o>N�併Έ���;�m�����������Q��[D���w�Yྻb	����L����ɾ,"=��=�7R�{���y� ���b��F���.?;i$>S�ʾm�M�g/-<isʾê������إ�),̾]�1�m!n��˟?��A?������V����;�����=�W?>W����䬾���==󱼋�=� �>m��=���C!3��~S�Zf.?�� ?�
��tOB�IP>h���@_=lJ_?��?�t^<ϐ�>��1?l�R�B��=��P>�i�<r�>9�>ϪL=;������k?��1?H2�AӾ�T>�9z���.���,=X9L>$�o���1u>�!=[b��= �;��7=HW?��>Q�)����9K����!�R�<=�x?��?��>�~k?�	C?�p�<e���M�S��#��v='�W?6�h?�>mоx;����5?-�e?(:O>|mh�o�龣�.��&��5??�n?�>?�U��q`}��������[6?�8t?�!i�w���[���=��0�>�V�>�M�>�y=����>"H?� �HL��\��h�5�!۠?�@<��?(Y�<���I�
=Ȼ�>���>��G��a��.)н������=�� ?Ғ��Y{��$�wF��};?eۆ?���>{������u��=| ��CL�?P�?����-l<��,Fl�����T\�<M��=����n$����7�:�ƾǢ
�b���J>�����>�Z@�轓��>)8�g1�KϿ>(��u�о��q���?y�>P�ǽ�L��l�j�G1u�|iG�w�H�Rz��4M�>f�>V��������{��q;�D4��.�>����>��S��&��Ϛ��M�5<��>���>6��>*)���潾�ę?d��@ο�������o�X?Bh�?�n�?p?�9<��v�v�{�->�:.G?�s?Z?��%��A]���7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�w�>T@�?���=7	�>x��=˨��9�#�PB2>��>�A�D$?�N?���>O2�=.i3�c�.�`�C���N�k��j�A��e�>|g`?>�J?P_>�N���z<�KY ��ɽg/��(ɼ�)>��&� �ݽ�&2>�?>oZ>��B�HyѾ��?ap�<�ؿ j���o'��54?N��>	�?#��V�t� ���;_?,z�>7��+���%��SB�e��?�G�?I�?��׾wS̼>A�>
J�>m�Խ&���]����7>3�B?s��D��f�o���>���?�@�ծ?gi�~�>G�3�|%������PԾ��z�>F�.?͛��~�>"&?ծ�=�o����1�z���>�'�?���?|?!��?QY���Uc�0�>���>�[�?>%?� (���bV�>#'?樝�t�����d�T?�9@̷@X&?�a��>�¿�τ�0b�����W�=�O<�W=\��IU=��(=��9=�'��d >��m>��=m#�=/[�=��>m>�ԁ�bD��@�������OJ�+�)�.B���a��*����������H��w���ɾ�)�섏�~���oy�<.�9>u<A?��N?�an?��?��'�a>�˨��Ԝ=�+'��=d}�>f,5?VW?Fr!?�	˽+���V�x�����{�(�S��*�>d߆>YG�>��>�x>"�=<r5>U>q�>�;{=�u�H\�~�)�Z�4>��>�>�}�>�C<>đ>Dϴ��1��j�h��
w�p̽/�?v���M�J��1���9��ɦ���h�=Eb.?|>���?пf����2H?#���u)��+���>y�0?�cW?(�>��]�T�:>@����j�?`>�+ �sl���)��%Q>ml?,�f>�6u>n�3�Bb8�/�P�.|���f|>�06?�Զ�
69�=�u��H��OݾhM>/;>BE�>k������vi��^{=&z:?��?3���᰾�u�X>��8R>%\>^�=$��=m;M>�Zc�F�ƽ�H��.=?��=��^>r?nG>��=��>����ʜ�b[�>�|�>[�j>��2?#?IT�<�����(��v�cDA>3|�>�^�>m4�=��J���=a��>�S>q���#���&���I���T>f�g�'���'��`�=��B��a�==ŭ=
�㽜?3����<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>	w�UZ������u�Ȳ#=��>�8H?RU����O��>� w
??�^�������ȿY|v���>|�?���?��m��A��A@�*��>=��??gY?�oi>�g۾=bZ����>��@?�R?��>�9�`�'��?�޶?���?s�H>Tn�?��s?��>��u�0k/�d�������]{=-�V;�>��>�m��eF� ⓿W��m�j�l���b>�>$=���>�㽬.���x�=C׋��N��lg���>i�r>�J>29�>�/?���>�f�>��=�m��mˀ� >����X?��?���g�,�\;�;�=ŀ�h�?P�]?�<(>�p+��&�>k?-F�?�G?C�n:����ؠ�/�ο�����RĽiC�>��,?˙�>���%�f>4�Q�#�,���ؼ��>��=���97���A�=��->n?-E?ݰ�=&?�� ?��f>��>�o��g����a�[��>��? A?�bd?�?8G���q.�T��{{��F%m��i=O+�?_�8?]��>�v��4`��ԇ���Z�=�{�q�?���?Ҕ��.?Xz�?�?�^?q��=�9��(���_��x��>��!?�����A��E&����bv?�P?���>�ߒ�L�ս�Wּe���d���?�\?/&?���!a��þ�X�<<�#���W��!�;%+D�ִ>և>F)��_��=7%>c�=�Fm��_6�C@d<�;�=���>�3�=��6���T[?EM��Z2��3<�����	K��Ţ>��?>غ̾��O?~e�O��� ������>f'�[v�?�&�?d��?�%���v���W?o�y?[G?�?����pCi��������˾��M_>H�>e,���ݾ{���Ѫ�'�m��h���D�l�>\!�>��)?Ξ?��1=1�>�M��{�B�B ��	�D,J��{��;�ٮ<��U����G��B��t	���.q�$�>����Ѻ>��>f�e>6�v>[��>�lX>�ט>�,>� �>	T=�"x=�/>>r	y=b��݌��JR?���n�'�������E B?^kd?kQ�>��g����Y����?���?o�?"v>�h�_%+��g?\�>j���`
?<
:=SX�#�<�\������f����'��>"�ֽt:�.M�Пf�^Y
?-?��nJ̾�hֽ
2�����<�%?�4<?����)V�H�_�BO��iO�n�B=����ʠ�
���z��ɔ��{�0��26�k�>�+?�k�?�������#����W�U:I�{Id>�^%?Z?ex�>{��>lb�����
�E�S�9��q����>i��?q��>�FD?�6?&TI?�nC?W�<>9�>�]u���?q�,<���>�?6�8?�6?�(?6�?�u!?t>H��ŗ�W�׾	?q?�y?%
?F?�ċ�1�սAȼ��<~�1��B���,=�؅<� ���սAl�<5�Z>��?2��S�7����Oel>�(6?N��>"[�>Dی��{��G)�<ԧ�>��
?
{�>����{lr����� �>ޡ�?�t���<%V(><|�=�,���Ϩ�w��=����ܒ=�rL���+��<�[�=��=�S��S;���;Gg<\��<�_�>Ar?Uk�>$;�>H�w���۾*�˫y�I�,>/�=��3;��վu'������
.d�D�r>�^�?���?��{=� >@��t�����M�-W���ؾ�]>*�?7��>W�F?|?(�??R�D?}H]>���	���h���꾁2(?s ,?��>���v�ʾ��.�3�A�?�Z?=a����;)���¾��Խ��>h\/��.~�y���D�S҅���������?k��?k
A���6��v�򾘿�[��#�C?X"�>YW�>f�>��)���g�9$�;/;>9��>�R?*�>��O?~	{?�v[?�?T>��8��𭿡\������!>m@?u��?�׎?},y?*^�>p�>m)�z�߾/e��H��KZ󽡪��HuX=��Z>�˒>��>``�>)x�=TIǽe�����=��p�=5b>c�>�I�>ZV�>g�v>���<��G?h��>�Y��ʕ�줾wă�U+=��u?���?��+?2=����E�FD���F�>�n�?%��?�3*?�S����=,�ּ�඾1�q��%�>�ٹ>o0�>vɓ=C�F=�d>��>ϡ�>�+�b�zq8��UM�#�?bF?���=[�ſs�p���u��.�����<UK��mwa��Κ�c�ւ�=�2�����!��W`��U��$����״�ݷ������ƈ�>?�|=� >�z�=^I�<����أ�<B�B=^-�<�=�dt��Q�<��:�)�<���A6u��}Z<�j?=�f �=aȾ�|?L[I?�,?uD?Oq>y�>�m���>�|���?ҫ\>�/:��>����6�����Ɣ��־��־�a�.��G�
>6 K��C>D7>T)�=Fv@<aT�=��|=7�=z��bd="f�=Լ=���=X�=9L>&�>	�p?��������alf� ^����}?D|�>�*�=8�վ�\?7�
?��|��ϳ��� �tUM?̚�?�'�?��?[����>l����J+9=�h=�=��lz��$�R>-Ƚ\o�>�]�>�t��i��$�&���?K�@xZG?�or��}Ŀ��h>~8�:&�>��h�P/"�dQh��i������?M�_�Jg�f/�>�x
�M�����f�7>��n>�i�=g���yi�:�Z=zyU��g�=.Ż=���>�$}>���0n�X��<C����5�=�>6�6̼_B�1��<���=���=a=)=�u�>�?�H0?Bd?�
�>�m� �ξ������>8��=���>�<�='hB>�>�7?�dD?��K?wd�>K�=>޺>ѹ�>0k,��mm��循���69�<k��?Ǿ�?���>ri[<��@�i���l>��)ƽe?�W1?;�?Z�>�U����9Y&���.�$���{4��+=�mr��QU�N���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=%�����<�vż�����u&�:�+�1�����;r��;@�]<Z��;��]�n�>��u�-S�>�\�<�"����>�S�a�d�u�<*�Y�	/M�G�i����I7���k�[�C>s�>����D���!?x��=��r>�J�?��x?��=���,w�����`=�ֽ#��{�>蟾x;?���^�=E��Z����>���>���>��m>��+�c2?��!w=:⾽�5��]�>Aތ�ub�9��Rq��:��0⟿`i��"�gD?�-��+�=��}?àI?ݏ?� �>���w�׾�G/>����x=<�1o�$����?��&?���>��쾡�D�*IH��o]��Y>��Ⱦ�G������D���_=����>צ]����� �(�t����!���G1���u���?l�O?A�?7����L���up�����@%=�RG?�c?��>���>�?�B=����h����=oP�?%�?7��?��R>�0�=�=�� +�>[	?���?<t�?IXs?�=�D��>:�;h� >�x�����=+�>�C�=�y�={	?�a
?�X
?��S�	�?��'{�)^��y�<~��=Pf�>qv�>q�s>�8�=��e=ws�=ԦZ>��>,,�>j�e>
��>��>O
�'��(�>�\=>6�>;=?�>\չ�O¾[P���[�=Pwp�g׾
�8����=
��=QX�<4�L=�sT��%�>�9ο#i�?���=�;�a�?c�־�P�=8��>��>��M��_�>	�=Z6�>Is�<�>]>�=S�>�9�>�IӾ�x>����\!��(C�уR�#�Ѿvqz>ӝ����%����|��.I��t���k�f
j��-��<=��S�<�F�?Ѩ��y�k���)����'�?�P�>6?�Č�q�����>n��>Wύ>�F������ȍ�g�l�?���?��|�=#�>c�??C�"?�����3m��Bs�6�����H�s��� ;z������i~����W���a?tґ?��?	��=�e`>|Ё?�ժ�tʏ�7�v>>�����D�S�W>��>Tо������i���R��=�+�=P�K?���?[*?,�k��>���=�da?��O?.Ԅ?��>�?�(>�/?���>'z�>��\?&!@?8C?#�?��2�4t\�ο��M�%= ���|�p��<:=-�X��;�$�=��<�=���v>mI���@�a.�=,�="8>�V�=n�H��K����=��3>�fV?,?%�~>�?}'��sse��I
� 9+?(��8@�.�Ǿ7G۾�e۾ů�fu?9��?&b?�#>9q��ٯD�$-)>7PE>�\K>d&>\~�>�𓽗�/�y�O>�>��e>��u=�Ђ��Z��%s�򐊾��B>���<Y�>t {>T��_�&>����Q{�r�e>;'Q��J���T��G��2��pw�E��>�UL?Q�?��=	D辏͖�ӌf���)?��;?gGM?� �?藕=��۾�b9��-K�̂��+�>���<���w��U���+;��^��ws>o🾌���0�b>�y�1L޾5jn���I����?H=n�-zR=�8�0־�h��=D�	>a���M� ���b���(�I?S�o=����zV�1򹾺3>�R�>W$�>�A9�C�s�]h@�FB�����=��>�;>�����(�ÑG�S �F2�>�WD?<7\?��?Ga��G�m���>�U;�)`��%�;��(?m�>|�?�9<>�M�=�#��f��rza�K?����>9(�>`���5L��#��<���"�&���>_x	?g'4>4`?<4J?��?/�j?	�,?o��>	��>�)ͽu����A&?%��?r�=��Խ�T���8��F�z��>��)?p�B�s��>9�?��?��&?�Q?X�?x�>� ��B@�D��>{Y�>j�W�)b��&�_>٫J?{��>�<Y?�ԃ?��=>��5�&ꢾ'ϩ�d�=7>��2?-5#?��?���>F�>����{��=+��>�Ec?�)�?�o?�y�=��?fE3>~�>���=���>n��>�K?�1O?��s?ǈJ?���>���<����8��?�|�o�S�܂�;�kI<��{=0>�ѵm�>�����<��;鷼�k�����6mB��틼�[�;`V�>�t>�1>�ľ�!���q@>�%���L�������:���=�p�>=?���>�o#����=���>N5�>j��d'(?n�?�#??8;��b��ھ��K� �>y�A?�=��l��~��U�u�N�g= �m?�^?Z W����~�k?�	r?#9�Ja�B��揾�J˾>��a?�� �{��>�|�?�1�?+�?	p�vFy�c���}�u���+>C��>��̾�r���?%HN?�<�>��'>���<?���Hu��{6����>��a?9Y�?�]?�S�>淌����`b��H��s[b?a�>h���D�+?|����郾<����ʾs�f�����'���c���[m���K�N�ͽ ��=�?;.v?'gu?�P?Xb��
G��2K�vT�� �K����M:$��B�^8G��k4�Y��M���	��O�����=1�|��A���?,�'?�P.�� �>�7��z���M̾֋6>L���C��({�=�o���=6�]=żb�q-�ۧ���]?�I�>d��>�T;?�Z��<�3�/���;������K5>�c�>�׍>��>_8;6P+�Y��ξ缇��9ʽ`@v>�_c?�kK?��m?����V0�������!�J-�*Ԩ�V�=>��>R��>�%S�eq��&���=�7�r�}���[��_f	��|=�2?�͂>8��> ��?�-?h	��(��h�v��1���y<H�>��h?W4�>���>N�ƽe��g��>��j?�|�>�-%?I7���`��U8��r��-��>+tz>��?��=��ý$�D�����Jz�97�t�[=7�b?r��9"�h��>�L?���<�ZI�i��>��Լ��)����][!=��>�?�oX��>�e>�'�n�W�"�GA)?��?���fp*��5~>��!?x(�>is�>.�?��>~Kľs\�_�?�^?�HJ?ȿ@?؟�>j�=����ɽ�H'�85=�x�>a�[>�oi=���=J���\�j �R�G=���=��׼Sڻ��n�;)����M<���<�4>	ܿn-O�zI̾W� >��M@���z���}*z���ڽ����p:}��uy��
�򍕼�3c�adV�`'����L�;H�?���?@R�����
����݂�3~��A�>��L���������$.��虾�5�Ax��$��"H���W���U�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�yA?��(����V=-��>��	?��?>�Y1��F�����N�>7�?��?,M=��W���	��~e?G<�F�v0ݻ0�=_�=W�=���y�J>�Z�>i���\A�ܽ�4>3Ӆ>��"����^��G�<�c]>4�ս8����?y\���g�̪.�������>�^V?���>�ǝ=�D-?|F��Ͽ	_���]?�|�??��?�+?0��~j�>�޾*xN?�7?c��>�&�+Kw���=l�����.�_i後JW��_�=u��>#�>���g����Q�+�Q����=�	���ÿ�d��*��iX�'�$�,��]	��u�y�ǰ<���c����%Xr=��#>(�>�u>	 />3�j>COP?k�x?L(�>[b�<S��)�������<|�����7q���/��4��A��L�ݾq��I���߾�߅�!"=���=�1R�f����� ��b���F�P�.?�u$>@�ʾ�M���-<�oʾ?����Ą�'꥽�*̾�1�n�|˟?��A?�����V�&��Jn�󚹽��W?�K�����笾ԏ�=�(��a�=� �>��=��⾆3��{S�qb0?�s?Y3������)>����o =�N+?ԅ?U[G<�r�>:�$?|*�]�d�Y>�d3>�J�>�c�>��>M�����ݽ$B?01U?M� �"���X�>�X��l�|��i=�)
>DA5���9k[>��<X���v���������<�$W?О�>�)�� ��W��N��q==��x?��?�>H|k?#�B?$]�<�o����S����6w=��W?%$i?Զ>	x��s	о�w��k�5?�e?��N>vh����A�.�T��(?��n?Aa?S'���u}��������j6?��?@s��ſ\]�ԩʾ	{>?��X?��?�)��?q��?M��pĦ�⻿f�9�)��?��@]��?ͧ>J�<v�=���>�8�>�9�3<��x�g���~��>��>Ui��K�s��r�b��C�?�ϊ?`��>�� �ؾp >�k��wh�?z+�?ֳ����+>����e���R �Ϋ�:����I��f����5�������ݾ���&-�@^>��@ ]'�a_�>�e5�ٿ������}�2����U�>�5�=��;RB�� 5�g��WL�tRP� V|�gM�>��>��������3�{��o;��\����>����>��S�a'������J^5<�>Ȫ�>䶆>�+��/潾eę?�\���?ο0���,���X?+g�?Fo�?�p?�:<n�v�ȗ{���� 1G?��s?�Z?�~%�-@]�F�7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�b�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�3�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0� f\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>dH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?���>x�?���=l`�>��=����W��h!>��=Y�/��?��L?�*�>��=ʞ5�q~.���E��R�>e��C�I�>�b?��L?� e>�R����2�^� �4ѽy�4�g޼��<��y3�,���0>��=>>>ʲE���Ѿ��?2u�$�ؿsi���(�O_4?Vh�>A?�����s��%��J4_?�y�>0�I����������?�.�?!	?��׾!qټ�>��>�*�>Q.ҽt��?Շ��7>�B?�E��=��o�o�e�>��?��@�׮?��h���?���R���}���'��{v=Qe�>%�X?����]�>s#'?��0>CCU��)���Ƒ��ְ>隩?.�?�?�Dw?/�r�T�c�6 >-��>K�?�#?B`������~�=66?2<Ҿ���~�"�2-`?�@�7@�a?�'��6GɿZ枿j������N=�)�=��8>�񽗳����=��=�<��� �=��>\�>�ҏ>!�>O<#>�	L=n����˧����9��|�FC���ߑ���:��y��漾@};�M��νM什$�B��y,��ɴ��p:>� E?O�b?>rK?�a?�� �`舽Q|ϾL�H>p��9�F���'>�}?�JP?�*?��'�Ym��A�v�E�^�Q���GꪾIͷ>頴>�2�>�w|>��>I�=���� 3=\��>�>�i8=��=R"�=4+">�4�>4��>�!�>�C<>��>Eϴ��1��j�h��
w�o̽0�?|���Q�J��1���9��Ц���h�=Hb.?|>���?пg����2H?&���y)��+���>|�0?�cW?!�>!��Z�T�2:>=����j�7`>�+ �}l���)��%Q>wl?��f>��u>0y3�Hb8�ץP�hN��7�{>)6?w���5�8��u�L�H��ݾ��M>��>�FI��b�x�����f�i��{=~z:?/�?��������u�0G���R>K�[>�9=��=n�L>h�d���ƽ��G�,�.=���=�_>AW?u.,>U��=�L�>�e��A P�5{�>��A>V,>��??1%?�X�Dm���o���j.���v>�9�>O�>g>UJ���=x]�>?�b>4Q�e1�����}�?��V>~r{�W_^�j�s���x=C������=�|�=v��\=��.(=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�>�>��!�H	���p��ㅿo�;���>��`?V��_Ł=qWs�Q��>���>�f����p����u�eD�>HT�? P�?FCn�c����5�>��>Ǝ�?y��?YZ�>J�����j��>nzL?Z?� �>�+���p<?G��?]�g?��L>���?Z�m?��>Ӿe�^P �@�������^I=��q�e�K>9:6=�����b4����� ���]b�=�y�<>�S�<
o�>�S�ʕȾ�>Dե��8��_O���>�E�>J8>�K>�?�?�ӳ>�~<biĽ�3���`����R?;��?'�ӾR�<)`=f�j>mF����>�i?X<�>FyA�uC���l?oT�?q�i?����%"��������Կ����OŮ��)�>�
?���>�B�:"=�\��|U���>�B>/�/���Y.x����=��>�P�>Pk�>R�h>�r?�-?:f>.~?��D��?��� 쾱bi>���>�$�>��p?�N?3����X�V���>��؀�����=�m�?��?GQR>��󄳿��_�|��߯���I?:Ȕ?�>)D?Y�?&�U?�[?z��>�9�R����zU�Yh�>��!?8��A��I&���B�?��?�N�>���-�ֽZE޼A�^2���$?t\?|�%?E��v>a�3þ�T�<�����g�bb<��6�>�+>����1�=R>T~�=��m��H6���s<�Ƚ=���>Ц�=�p6�Qލ�e
3?R�������H<���NFN�~��>J��>��t�I?��� ������ڐ���%=S�?��?㳨?����}��#[?2B�?�g�>.'	??�˾�W#���@���߾�o�-ӾS:�f�> X ��z�?��o1����P��hr�x�W ?Z"�>�{?�#?�>@>$m�>PҎ��zJ�-� ���˾��;�J�!�L�=�*������#v��ܽ�O����Zv>$���-g�>�	?��Q>�`>->�>/� ��d>+5�>T�>�Z�>�as>W>�?>��b��搽�KR?#��� �'���辋���Q3B?�qd?�0�>�i�,������J�?���?Is�?�<v>h��,+�n?>�>1��@q
?[T:=�4��?�<�U��2��R2����X��>�F׽� :��M��mf�}j
?�/?�����̾)>׽P��o�=ɷ�?�?�p��[�%�}�J�P�ƾI�k�y��I�����ߝ�zi�I'�����C����#��>��:?�(|?�E �oJ�ݒϾV�U��	�"}�>5%�>���>O��>o�=�}�$�k'i�+@.�O���?�>��a?��>tI?�O<?�(O?�NK?\9�>N�>�����b�>��U<�V�>��>��8?9�-?��/?PR?�")?��R>Z���Z��X�پs?��?��?���>"�?DǄ�l�Ͻ?�̼����(r�u����op=��q<��ҽJ����H=�T>wT?����8�D���/k>�}7?�{�>���>t)��jD���j�<��>�
?\;�>�����{r��_�U�>���?�	��Z=ʾ)>��=n�i+Ϻ�M�=�����=�C��[�;�U <���=1�=��p�^�w��X�:�B�;���<9D�>�}4?v-�>4�>Rh��y���^A"�ν�d>fp�;�wº�5����t��	����^�|��>��?6�?�R�<�>
��=�����Du��4������>�E?X�?y�J?:��?}�&?�5?��3>i�����}Ƃ���ξ�?3!,?5��>���ԫʾ񨿱�3���?Y?�;a�v��:)�_�¾�ԽN�>�\/��-~����RD�������~��%��?A��?FA���6��r�h���C`��n�C?7'�>�Z�>�>j�)�^�g�r%�*#;>���>$R?���>��O?�{?9P[?^�U>�8���������X1��� >�??��?Q��?�!y?���>�<>?�)�
��+����! ��6�ۂ��]=<D[>���>V��>��>�{�=�Ƚ%��ܲ>�Y�=�a>E��>�>!��>C@z>�޵<i�G?���>�W��ő�@����d=��u?���?I�+?��= ��V�E�E���>�>�l�?F��?A1*?4�S����=�p׼s嶾�q�*�>8չ>CA�>�=KhF=w>�>��>K� X��r8��sM���?	F?2��=�W����K���2�����w����g��.�F;3�ּ��>l�z����<�E��x�����F.���Z^���!�&�=�� ?�F8>l">�<> ��=�����|���L������C�õ<�W�$KA=�����c��X<�����ń����=cNȾ�d{?��@?�	-?S<K?]u>�q>��2���}>�vн�A?�
e>�1��X���NO4�+}���K��u�Ͼ�۾qa�疦�+>� E���>��4>�?�=X��<Ì�=>
�=�ф=v^�;�Mv=���=��=5��=	� >HN>Ҫ>�Hw?����Vҝ�vQ�/����:?[Β>ٮ=Hdƾ2@?=@>�!��j�������~?���?�V�?	�?�i�DK�>�Ϣ�Lq��즐=|Z���1>�5�=8�2�?չ>�J>����@�������?��@$�??�ɋ�]{Ͽ />?�.>N>T��f%�ƣ�Q�^�)[B� e?�=G����Ŋ�>v��=��c�Ѿx|%=��">�*Y=&<��3�\���=޾���~=��=Ra�>{s@>��=p��ڪ�=��=g~�= �i>+�<�����¼�=Q��=��O>	�(>���>Q#?�P0?�*d?�P�>�.m�ֺϾ�¾�%�>:��=qy�>���=��A>��>��7?��D?&L?i��>Y��=(�>�O�>G~,���m�O澇������<#��?�ц?;|�>��O<��@��&�OQ>���ƽ�o?�01?�?�Ş>����LkξU�8� ���R�a�V>VLO�nDA���=�]��+IX��L>[4�>^}�>`��>)�=$�=���=�p�>��F>Y�<K/=�a=$K�=���;�>�>t=s2���>�k�<��#�# �:@޷���;�����g?=%F�={�>+�����>�;">�2���$>Kqм��}���G�C� ��gG�����	��$:!�[���j�=���>�G[�����g?%�N>j��>�x�?u9`?>�E>�ʾ֢��緿�F�W>�`]>�1>����_^��>�W�tY۾���>x��>d�>�l>�
,��!?�C�w=}�Hc5��
�>{��#���,�}9q��?��C���%i�ejѺ�D?�E��C��=�~?̰I?h�?��>1���ؾ(50>fH����=f��#q�X����?�'?���>:���D�)xƾ<Ľ��>�b��˚R��̕���2�u7=q���욽>�荾�޾��.�-)��cc��ZAK�1���}}�>�[?���?j�h�%����	P���.���=@�2?p��?ԁ|>k}?��?2h���ƾ��C��񎽬�e?���?9N�?��>e_�=Aj�����>[<	?wՖ?��? rs?9?�.��>�zE;~-!>�C�� S�=�#>ƹ�=u�=Wf?	�
?�
?3����	������l^�ai�<��=9��>���>�r>^|�=-h=Y��=4\>'��>A�>�Re>��>F�>L��a��.2�>q�V>�P�>�,?E�J>h5m>�����͖�=��<m�p��Vp�H,�U��;�X>?;>G�0�Ġ�>5�п1��?��=��:��p4?o;�Ǉ�1�?w�>�Vk���>,��=ׁP>�ث=a��>��`>l��=v�E>Ծ �>�i	�i.!��B��DS��kվ�ot>n��>�"��Q�����.K�ܶ�W����j�]
���<���=���?Ya����l��**��
���?���>_]8?����Q�t��>�<�>��>v���K����#��yTᾒ�?$�?Y\_>Ѳ�>]#B?J�?��=R�a=K�}��#��@,�5�z��Mq�?`��Cps�{C�_�"�!Y.?"��?�x3?�q#��m�>noq?o6�&�`��.>����� �\�5���>�7¾#SW�c/}�����ھ��$=$.h?��?�\7?U�O��n�;��>"yw?�R?f2�?D7�>c�?ܕ>�E?��>�`o>�	?� =?�4X?CT?�r=.c����K��_`=���ʿk��}>�7���,�=G�>4;�=�<,;��4=���=֔@<�.C�1���qƍ���8=TR�<-�`>���=���>M�h?��>V��>0?R��n�=�d�ʾ.?� ��J��qK��l�w��߾�<�`U?jp�?�&E?�2>N�'�F����q=g��>*�=��>Tf?4����e���X>(7�>P��=��#>/x�=��������;����g�M>���>�7>ˌ�R/>l{����v�u�b>��T������U��!G�j�2�-As���>�I?Y�?��=�d�r㕽�>e��q'?�p;?�*O?9'?�v�=�G־��9��K������>��<�������ޡ��$:�N�gko>����'ޠ��Xb>ս�Es޾��n�<J�h��BM=���YV=p���վ�3���=-"
>k����� �����֪��0J?�j=�w��-_U�Fo����> ��>�ޮ>w�:�n�v���@�����8�=L��>x�:>Fi��z�~G�68���>x�C?_?��?�"j��Lt�S|@��* ������{ּГ?��>�?`=>�H�=>H���a�!�_�eIB��2�>`�>�*���I������辨�%��w�> �?�/>�?-�S?�p?�_?�3(?��>���>����q���A&?��?��=`�Խ��T� 9�MF����>D�)?��B�D��>W�?0�?��&?��Q?G�?�>�� ��B@�e��>:Y�>��W�hb����_>�J?J��>c=Y?�ԃ?\�=>�5�颾�ԩ��O�=�>��2?6#?��?j��>r��>?���i�=���>�c?�0�?�o?Ѓ�=-�?j:2>N��>��=���>M��>�?OXO?<�s?��J?��>\��<�7���8��Ds���O�Wʂ;�tH<��y=��3t��J���<��;gg���I������D�����g��;#;�>�Ms>s�����2>�ž�򈾺rA>{;���n�����Ö:�dt�=�:�>]�?�2�>��"�m�=\�>A4�>����(?e�?�"?�-: �b��%۾��L�g��>��A?S�=`m�����4Wu��/m=��m?�^?OpW�b����t?�J{?k���o-��5ľ2��=C|��6?2N?O���?e��?~��??q$?j���怿'.�������[>%MA=��>�����c�	��>�F?�g�>"�>�콘����w����ž?��J?�~�?�1n?O0>�zX���ۿ�H�X����a?m��>F��:�?��?�r[����$�pƾA����J���㭾쾼�5AB��K���Tؽ��<�;?�d�?^m?Vu]?�"	�j`V�m�g�-a��n=����
�V���<�c�Y���)�!�e����־���=�kf���G����?PY2?i���?�W�w���	ʾ�=":�����

=�B��,�$���=/�G��-�D÷�pZ?q��>���>��Q?�Gn��D��7�@7\�P�O�m>`q><�t>v��>]t�<�>�����e��}���)�Q<F�u>Dc?'�J?�oo?=��:3�����!� �B�Zj���4A>p`>;�>x�Y��q!��:&�m�=��q���\��6�	�M�=�T3?�>j��>G^�?yI?�S
�
M��W�{�X�/���<޺>��h?���>�Ʉ>�Ͻ]���3�>g�d?^J�>��>j�WI���`�������>l�]>og�>!��=�P��`Z���˗��^y%��>�A?'���lDo���v>��b?zs�=R��R��>�6�LT5�Z����P���6>h�?��>�C>�_꾲j#�(hl�r�j��N)?M?�ޒ���*�`2~>S"?�y�>Z)�>�0�?�(�>Bvþd=��?��^?�@J?vPA?,E�>Ly=E���FȽJ�&��,=g��>��Z>��l=�r�=����j\��y��E=d��=�μ}g��j�<����ZK<���<
�3>8�ۿ��K�ϝԾ�����񾂲	�H��)r�����a�� ���v/���+w�AN�n/� �X�o.e�+�����m���?T9�?�U�������䙿9������>��o�v艽6����1�胘�	J澑4���7#�N�P�j�i�eSd�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�zA?��(����=dV=G��>�	?@�?>$_1��J�=���~M�>e:�?���?gM=��W�S�	��{e?h�<��F���ܻ��=�L�=B=���6�J>�N�>t���6A�`ܽ��4>&ޅ>F"�����^��@�<|y]>��սE���T�?��Z�΢z��'�M������=2�v?Ǩ ?��<4�N?�,>��JƿKyv��U??^��?޻�?[+?�cG����>�K���?Z?�VM?�M�>S�#��3��ّټ�c�=�V*<#_侵!s��倽���>	>&���A���č��P����x=>��^�ȿ������N@�<��K�y%���!ɽ��׽e�y������1�-"��ְ�=TU>nE>{Nk>^�n>F�C>�pW?�Tw??��>�I>u���V�����GᲽ�Di��p����m�'b4���Ӿ����X �S�����!K�'�Ͼ!=� �=7R�l���9� �f�b�Q�F���.?�v$>o�ʾ��M���-<�pʾu����ۄ��ॽ�-̾�1�)"n�i͟?��A?������V�L���W�����K�W?UP�޻��ꬾ)��=׭���=�$�>���=���� 3��~S��n0?V]?~���O��q:*>���z=g�+?��?��X<��>�B%?��*��c�dF[>��3>�У>]��>��>����D۽s�?ՌT?������A��>�q��s�z�m{`=rS>:5���鼟�[>9��<�����W��9��qL�<�`Y?Ѷ�>�&�dV� ����a6�9d<x�r?n?�J�>�cq?��H?�@4=��_�T�H���rT<��J?>bq?L>S1�?Ͼ�B��N4?��k?�8Z>9"��Z6�O5�����e?�Lp?{�?>4D�a�u��ґ�'�ǔ8?8�p?4j�t��@H	�gqz���>�I?�:
?=�?��;�>�3k?�3��-���c����,� �?F�@�D�?1Ť=�<m��<|A�>�P�>ƻ%�c��0�=���z>>XZ�>>����8o��LQ�5�н$_?ԏ?�>=���Y_��|�=���M�?�g�?[�����<�q�¡m�o�����<C�=�@�"Z(�?Y>8��]žѽ	������üÚ�>{@@�=�f�>>�?�2�Ώ�ο~��Ïо��n��\?ᴧ>:�˽�Ϡ�^�h��s�5<E�|iH�ԅ��{I�>��>��2 ����{��o;����5�>:�y�>�S��*�������4<\ݒ>��>Ҵ�>\�[ݽ��ƙ?Id���Bο^���"���X?�j�?Lp�?�l?�]:<��v��o{�}��E/G?܁s?Z?>�$��]���7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?*�a�M�p���-���ƽ�ۡ>�0��e\�!N�����Xe����@y����?N^�?i�?ҵ�� #�g6%?�>b����8Ǿ��<���>�(�> *N>`H_���u>����:�i	>���?�~�?Pj?���� ����U>	�}?�
�>ϱ�?� >��>��>5D��to(�z'>[�>�Ƽ8��>5DP?٢�>��=)*�S�.��/F�bwU�q��GSA�q�}>�,b?�Q?�n>8�Խ��_�������'D��q��>'�}�N��｛�2>�*>�>@7�欿���?-q���ؿj��v'�U64?�>z�?��L�t�|�o:_?�w�> 8�X,��L$��4:���? F�?Y�?׼׾A�̼�>��>�N�>��Խ��������7>
�B?��>E��d�o�M�>>��?�@�Ԯ?:i� l?���N=��Y��^���|��\:>zWc?\�A��>��"?��=Q#`�%�������>a��?�<�?���>f�y?�h�`�u��^�=��>#B�?s+A?��(��.��}�=!s"?,��U�������K?4�@�"@ElF?e�����ۿx𤿕���T���o>r
+>�E�>>;����=l��=]���%���H>�>L�>&->�>s >|�(>�L���q"���_����p/��I�B� �P'����XP��i��%��:ા1�hC!�������=�u�)�Jώ�g�@>{�J?�`W?��]?3?tͮ��y >�qt�Cۨ>�R =��t��?�W?��y?��B?@+:�\Bľ��j��J|��`������x�>!_.>�K�>�A�>pX�>�#��2�<,)9=���>"�%>� ��v=��8>dd>px�>s��>�7�>�C<>��>Fϴ��1��j�h��
w�n̽1�?~���Q�J��1���9��Ѧ���h�=Hb.?|>���?пf����2H?&���z)��+���>{�0?�cW?!�>"��t�T�-:>=����j�5`>�+ �|l���)��%Q>ul?u�f>+&u>*�3�Ye8�s�P�|��:i|>{36?�ᶾ59���u�ĭH��Xݾ�QM>ž>!�D��l�����3��yi�9�{="x:?8�?�,���氾įu�bD���PR>0\>uj=�t�=ySM>�oc�L�ƽ{
H��.=��='�^>�L?��+>��=�+�>,���6Q�=��>3�A>�|+>��??M%?����l��헃��f.���v>3�>D�>�(>
;J�B��=�i�>��a>d������z���?�
[W>�I|��_��/s�uz=����<�=1i�=�� ���<�W7'=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�O�>���0V������u��#=m�>lJH?d?���.N��=�Z
?2?�v�X����ȿ3kv���>���?`��?��m��U��@@��^�>���?��Y?�i>2v۾Z����>��@?S�Q?�5�>�B��'��?�?7��?{I>V3�?�os?
+�>-:_��/�����Jq���q=��+;俎>�{>NB��+�E�����0C���<j������b>n�*=�P�>S�߽8����L�=�����!��`&c�y��>�`t>��J>L��>zH?�a�>0_�><�	=� ���]�������R?�c�?��Ͼ�D��y��=��=^�ĽF?��??
M�>'�<���>LK�?�r�? d>?ǭ�;	�9�汫���ɿ^�I��%�>�:?�Ѥ>����=��Ҝ�y>:�	>@��6����9�ERl�NQ�>*?S�>�Κ��&?R?���>�Z�>(�5����
KC�p��>J�?Po?�a? /$?at�E��Ɍ�7���*�d�<8X>%��?f�0?[ҫ>�/���\��<�ྜh
>��C���m?/_�?�0[�	F?�"�?V?/?��V?�$>�]����{Ҿ��>k�!?y�G�A�6O&�Y �?�O?���>i=��:�ս�\ּ���{���?(\?:?&?]��0,a�� þ�,�<�"��V�?>�;HXD��>��>������=B>���=�Um�_F6��g<�c�=Q��>��=+.7�܏���&?]������5C=\7����D�\ڟ>܃�>8$��C�f?ŋ��	���8^��L�������?LM�?8!�?v�[��o�.*E?�ă?�
?v�	?@ۛ�����׾2o����ʾ� ����=���>�W���b��E��P��Ç�7����/ν�}�>�x�>pD?ab0?�yn���>>�Ͼ��R�!P ��
���C�*Cؾ{�&��n;����PA��d��9��=!���Ē��÷>&���{��>��"?&\�=�T>��>~�>�>���>�s�>1��>u�c>G��=��n<uH=���=ELR?������'�@��+���4B?qqd?d1�>Ei����w���?І�?'s�?�>v>$h��-+�'l?a=�>;���p
?wO:=�<�N�<V��ҽ��%���$���>X׽�!:��M�3nf��i
?�/?#���̾�S׽:_�e ;CU�?k�?g��	dE�3ˁ���G��:F�~���cb�?����B�&�y�y������_=���"��F=��2?�?�6�ܟ�:櫾�L���R��I>V_�>�̷>â�>�7� �	�G��V�������[��>j�|?�e�>?aI?]<?UWP?�{L?K-�>ߊ�>PK�����>J��;��>�z�>P�9?/|.?ͳ0?�?̞*?��`>�<�����-ؾG�?k	?�(?�?�k?�R���xý�6��sO��1x������=!9�<0�ֽ~
w�LY=1U>�X?��ͬ8�V���Fk>B�7?��><��>����-��Y�<?�>��
?DF�> ��}r��b��V�>e��?���܃=��)>���=㉅��~Һ�Y�=������=s7��y;�@d<ǁ�=c��=NRt�$���H�:ꡇ;�l�<���>�% ?��>8c�>X�N�����i4���=,5>$<'��=��
�
�w����W{�I{�>_ߔ?i��?>I��D�=ؕ=-������7�m��l�:>�g�>���>њ2?=ܐ?��?�B?�A�=�R�钙�"���ޢ�����>J!,?B��>T��F�ʾt�y�3�ѝ?�Z?�<a���y;)�E�¾��Խ��>\/�C/~�����D�h�����g������?���?�A�c�6��w�ֿ���\��c�C? !�>�Y�>��>��)��g�%�I0;>���>AR?@�>#�O?@;{?V�[?;U>�8���@����:'�aL">o�??���?��?�:y?��>��>��)�K�w���� �����ӂ���U=��Y>�{�>
�>=Щ>p]�=X�Ƚ&;���`>�݄�=8�b>p��>���>P��>��w>�C�<LAE?5��>������,,���J�������*l?��?�S$?V/<p~�d/F�ˮ����>�?N�?��(?�M��Y�=�E�����v��ʾ>�[�>X�>Ф�=��H=�>B��>Yj�><�	����Y:�k�����?�K?:k=�ƿ)�q�ݸp�������g<R��.e��˔��![��P�=���ͣ�󹩾6�[��Š��������e���ɸ{����>�j�=_��=V��=U��<>ɼ!��<Y
K=e�<�z=�o�Fm<TQ8�[ѻ�z���u�q�[<$)J=����˾��|?k)F?ا*?E?k�v>�k>�4<�31�>������?o�S>|�o����F7�4\�����%վ�nپ
�a�Ĕ���>{�A�ۮ>��:>l�=j1?</��=ߛs=d6�=`����`=���=M:�=���=�N�=�@>y>�it?fv��ON���E��Cc�s�J?[�?t�>�rʾ Y?x��>��o��8��Y� s?���?`.�?�(?�����4�>(�R�1}=�_�=4G�䷅��>VA½���>I�>V�K�`𘿐�p����?Pg�?ܖ1?a���5ֵ� ʈ=y��= �;>��S�3�����9�F�P�%��T?*�o��l��&�>Y�=��	�iB
�w�=��>.��=�zz�N�^��0?=��޼`�l=<�=Nj�>���>��[=:+q��.<)� �F�">��K>�>w�N�;X����4L=���=�#^>\Ӣ=u��>�?�80?�c?̶>��j�i�о��ľ��>1i�=N��>��d=#<>ȸ>�w6?��E?!�L?�̰>��=�ܹ>M/�>1�,��m����:����'�<�1�?X��?���>�s2<�~<�p5�I�>�νB�?��0?��?2�>{p�J��z�B�)��r�94�<$��=�ם���V��e=��Q��3����<>�۶>��>6Z�>�@G>dD>�C?>���>�k>e�=�n=��������A�s<�ݽ������<q9�=�#ǻeMg���=�ή=X@�<�>-ݸ;�ɻ=���>fw�=`�>-�=eH���?4>S[Y���X�+<!=:H��_�<���d�D���S����T�C>"Tc>�~��'����?vb>:�=>���?�l?XO>%B\��w ����������x�����=/yO=�)���D�54Q��`<�ޏ����>��>��>�m>	�+�b>?��Rx=T�li5�y��>�y��3��+�7q�=@���񟿰i�gvƺ�D?�@��=]�=\~?*�I?��?�n�>W{��<�ؾ��/>o.��k�=�����p������?��&?=u�>
�O�D�ڡ���;E�4�>����T�I��~�k z���=d'�����>R�0����f�����np���o=�X]���&�>E@P?�B�?���f����k�����==C�$?_��?y��>�v6?;�?�{�<�_���H��Z��<��?���?ط�?�A%>��=洽,5�>3	?�Ė?���?�ts?��?�E�>�W�;Z� >����}@�=��>bA�=���=Ai?�
?��
?�&����	�A��R�Y9^��1�<wi�=胒>ȥ�>�r>v�=H"h=k٢=0L\>KҞ>wՏ>��d>���>�e�>Hx��9���>��=�;�>L�N?�IH>`�<�7���Ј��a�=r06�+ϥ��k?�jF�6>�=$�~=B��=`�E�P��>G�ҿ���?a*�>�B�qF,?�(��V��_��>�93>�4>�y��>��>O��>�ג=�ܒ>^�={�=m[>+@Ӿ�>���!T!�/C���R�!�Ѿ\z>���^&����`j���*I��n���k��
j��+��Y1=��k�<�E�?߲��Ͷk���)�Y���?MD�>r6? �������>��>�э>�?������]ƍ��qᾊ�?���?��i>�.�>¬O?sb=?%z��	>��A�������.ρ��V�����s�}��6�Y� ��?E��?���>lz�>O<>�e?�	���ܾ��]>����4�3`z>b��>�PQ�D����'�p
����_���>j_@?_^o?�
?���1���'>�)L?�0?��|?bp?��(?!�ֽ0'(?%�_> ?�o+?��<?Ӊ<?sc*?~<W=��/<g��Xe����~X������d<��ڢ=��=9�YrI���v9G�g=k
�����¼�c��3F=~=f��==��=%��>Y?��>�/p>�?)?�C��&{G��b���)?\�4�{��Jܵ��A��w�����&=�yj?j�?��W?�)>^�'�q?��5>ƀ>��B>Q2>7�x>ۄ�5)S��]<�B>�>�y>�qB�����a�����˧>q}I=���>�La>�3��|>]@��d}|�,ql>��v�� ׾�R8�79�NK:�=����W�>��\?�h?M��=Jþ+�2�8mj�:|.?X�.?��>?�u�?��>L|ﾾ,>�_�!YϾ�u�>�5>,ھIã��E���W�&gѼ��7>;����ɠ� �b>%���޾gBn��FJ��V��pO=[��+�S=w��?־�����=�

>oi���� �����ت�V�I?��k=)	���U�RI���>)��>S�>�3�
�v�x@�^���m�=&8�>ݙ:>~���W�*�G�4)��7�>�?E?Z:_?p�?Z���os� �B������M�� �ͼ��?a̫>c}? =A>��=N籾
���d�]�F��
�>��>,��*�G��J�����s�$�$V�>e?,�>��?0�R?�
?��`?��)?>?��>�C��L����A&?/��?3�=��Խ��T� 9�YF����>J�)?�B����>�?}�?�&?ʅQ?�?,�>έ ��C@����>�Y�>��W��b����_>k�J?���>K=Y?�ԃ?%�=>e�5��颾?֩�]T�=>[�2?�5#?0�?���>{��>I�����=ƞ�>�c?�0�? �o?��=;�?�:2>M��>*��=���>g��>�?SXO?=�s?��J?��>F��<7���8��4Ds�W�O�2ǂ;�tH<��y=���2t��J�8��<��;�g��HI������D�#������;�U�>��s>���1>��ľ�w����@>����v���⊾��:���=w�>��?���>*6#�r��=è�>�'�>#���:(?r�?�?��-;x�b���ھҫK�8�> �A?���=��l��~��B�u��Cg=��m?z^?�W�E/����a?�Ex?���(�G�o<��@��қ���?jkB?skE�>�?�ԁ?n�
?&zb��|�����|z����=�0�=��>���MTm��o?��?)]�>�	e>y�2���7�*���}�ܾ2�?<�b?���?�q?��*>��u�+�����[G����f?uX�>�����&?8v�<�Oվ�3��{������	ҫ���������7����-�r����� ���=9J?U�m?*�o?O�e?�e
�_�a���[�=��q[�������8��@D�1�K9Y������Ӿ���_�=�h��H�GO�?��8?5�[��>��q�Vr���"Ǿ�/>w�����%���<y[Խ�D�<��<��i��}�oƦ��?�J�>�%�>�kH?�d��f=�gm1�"�c�{����=;�>I�>e��>e�t=�i���(���5��N1O��f�	:v>�sc?�K?��n?�	�[,1����9�!��h.�+X��.�B>.�>�ω>�{W�-u�;&��Z>��r�����t����	��=֩2?F�>ް�>�O�?��?_~	��V��RFx��r1����<�,�>\i?66�>��>�нi� ���>}tN?�!�>�^?�P����|v}�"?�����>�s>��>s�^>�y=LW`�����E���� ��X>��d?rd�C�b�W2G>|W6?k��<ܱ��vr�>	�.>0��o
����ټ �m>lV?���<x�>�˾��G�%�R��N|=�I)?u\?�Ē�˗*���~>��!?Y�>:C�>�7�?�@�>Z�þn� �?��^?5DJ?�A?���>^u=�=��ÓȽ '�ܱ.=ɇ>B�Z>�"k=��=��;\�E���#G=Y�=G�̼7��k�<V۴�6�L<�t�<��3>�ܿ$I�.���OR�d�پ~�����������g<�Rŗ�*T����C�p���>�Ǽ@&\��f��\��KSj�S��?|��?��#��u�����4�x�7S�_��>�MY��^C������h����U3�,ľK1��X�L�R�S T�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�{A?��(�7�쾵AV=���>_�	?r�?>�V1� H�� ��7Q�>�;�?W��?�TM=��W���	��}e??�<2�F�ןݻ�=3�=�6=����J>U�>t~��GA�	Jܽ��4>k߅>)q"�E����^��A�<$|]>C�ս-��h�?@�i���g��/�3����O�=�Dv?�>*W��(�\?j!4���?w�?8G?I@[�?�?k��%�w>�%���6U?�?�1�>�>��z�b�0:�;#==�<�'��}��L�>�X�>QXf>��X�x#��>u��a����?��ƿzO$��V��`=��
Kg�5\�Z���)�V����%�m�dK彜]j=�T�=��P>��>�V>t=Y>��W?�4l?���>E�>W�Hʉ�=�ξ%���`灾��A���w�ܠ����N྿
��K��\�[ɾ�=���=�6R������ ���b�S�F���.?th$>2�ʾM�M�C-<qʾê��ׄ��ץ�'+̾Җ1�(#n��˟?�A?������V�����:�
��j�W?r>�&���ꬾ˜�=*ܱ�m�=�!�> ��=v��!3�y}S�0o0?4_?Up���N��l|*>�(�:=�+?�?Pq\<��>�B%?��*���㽷�[>f3>���>B~�>�>K����۽�?e�T?X��_�����>g����z���_=!�>�5��z鼶�[>�<5쌾�RV�����?�<)$W?���>��)�C��+f��@L�T==��x?��?�>K~k?�B?��<^e��W�S�*(��v="�W?�6i?/�>#H���оp���ε5??�e?��N>�_h�T��>�.��I�
(?�n?�_?�Ҝ��n}������Ui6?��v?	
a�M	����_�e���>�� ?;�>+>���>A�E?1�4�Z~��(ÿ��4�
��?��@8_�?��=��3��L=��>��>��=�ѝ�� ��������n=���>/-����z�z�#��$��D?�8�?e��>}>���&���=�&��dd�?�1�?�|���5p<��-5l�x��:��<Q�=�B��h%�3���7���ƾB�
�I��<��F��>�M@��0j�>V�9���mEϿ�M��C�о��r��?k�>�ʽ;����Ij���t��G��RH�7���M�>��>����x���G�{��q;��#����>��	�>�S��&�������5<Z�>Ǯ�>:��>r)���罾<ř?�c��@οO���؝���X?Eh�?�n�?q?��9<l�v�ǐ{����-G?{�s?lZ?�m%�D=]�j�7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�a�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>��0��e\�"N�����Xe����@y����?N^�?i�?Ե�� #�f6%?�>b����8Ǿ��<���>�(�>*N>cH_���u>����:�i	>���?�~�?Oj?���� ����U>	�}?Ȍ�>i��?i��=���>��>xճ�3�}�#�%>��>E2�T3 ?�EM?n��>�L�=f2�c#/���F���R��8��.B����>"�b?]�L?6�d>��Ž27H�5��dɽV�7���m�Q^3��6���ݽ�t->F1:>ǒ>�cA� �Ͼ��?Mp�9�ؿ j��"p'��54?0��>�?����t�����;_?Oz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>=�>�I�>?�Խ����]�����7>1�B?[��D��u�o�z�>���?
�@�ծ?ii�_�	?P 	�v����-���� ��4����|>.B?K���W�>?��<`����^ځ� ��>{l�?��?�>�>��?�����~�	��=���>�ׇ?��9?�(�F'��;>�#?���j�����:U?��@N
@o�7?=#��a�οt��%���O��;��=���=UE�>��=���� ��=�>>�4)<J�n>H��>��{>�A>YW>@�>y�>��z����?��� ��r�L��7+�����+6�B%���_�4����#�L�s�ڜ����<����u齺#��"!>$"B?جb?��[?�vA?s��e>�=�c��N�>it����w<��>��G?��Q?7*?D�����5}l��9��Y��W�����>=Zx>�q�>��>��>!�<Y�:>�V�>M1�>N��<f=m�>�	+>��>�;�>��>RC<>��>3ϴ��1��8�h�w��̽,�?g���N�J��1���9���eg�=0b.?|>����>пd����2H?U���H)��+�l�>��0?�cW?"�>����T�6:>���}�j��_>�+ ��l���)�%Q>xl?}|e>��v>ck3��_7��DO��*�}>m@6?a��.�:�(Yu���H���ݾ�H>s6�>�7���������o���i�u	y=A:?9�?#��0���e�t�S��dX>��[>{s=��=-XK>�l���Ƚ��H��� =�U�=Z�]>��?V�,>R�=Ed�>��mGU�ߌ�>��C>�&>�??��$?�5������*��1-� �w>���>{Ѐ>!>��J��.�=i�>g�`>����7�����>���X>Y���_@^�iJz�QMr=�o*�=��={��$>��=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ.h�>ex�lZ�������u��#=)��>�8H?iV����O�>��v
?�?_�ߩ����ȿ |v�7��>R�?���?b�m��A���@�^��>6��?�gY?�oi>�g۾_Z�͋�>��@?�R?��>�9���'���?߶?���?e4H>
=�?V�g?o�>�.�� 2��)���Z���#3=�oz�*}�>stJ>iV���L�$����wee�0���>�(I=�K�>\��r5о�p=Z![��|��H������>5>~q>���>96�>�J�>v̍>�A��#���g{�
)pD?�Q�?f羰e��D�>:Z_���
��
?�]?3�!> z@�|��>Hn?��h?��E?�l��u9�)�������������]�>�)?=��>��#��H=�Yb�3���˛4>�{R>��d��Sʾ��2��˗=,��>��?�/�>��*�m?b�$?��n>_`�> 7��|�2�:�(я>B�?t�>�?��C?��ཌྷe�~����x��%�f��y@>���?�?���>{�q�������M���="j���SK?��?�0�=x:?�e?�_?��U?*��>�/�M��k_��wO�>��!?�����A��P&�����w?�M?k��>����o�սs�׼?���a����?�!\?�3&?+��S1a�þB�<��"�XR�zm�;�B� �> s>�W�����=>ao�=�Zm��N6��f<�i�=M}�>�={87������6,?��F��郾�=ξr�9�D�>�>>YL>� ����^?$g=���{�&���u��w�T�G��?���?�e�?+Y����h�
'=?��?�?�+�>�N��
w޾?��I5w�ڞx��n��>V��>]�o���Q���&���D��#4ƽ#U'���?R7�>�?X^?��	;�q�>v�����(�5"���b�����K�>��f���o���IU�u-k�����"��䌽>͕׽0	�>~�J?
�W>�'�>�� ?��V=�RY>+N>u�>>ēF>2">i�=�@<���e �LR?H����'�s������2B?qd?�/�>��h����X����?憒?�r�?-<v>@h�a.+�k?�<�>���hp
?]Y:=�?��o�<;V������*��W���>[_׽;!:��M��nf��i
?</?S荼��̾�Z׽伾1L3=�ą?�K?��$�"�Z�bx�kGK�PM�~bH�+�K�8�������_i�o���������/=��5?��?�Jݾ�<�(�վ�[\�?�9��l�>�$�>^�>�|�>�d�=��J�<���e�P�1������ ?��}?pt�>xqI?<?RhP?�L?&6�>�\�>J���C��>��;��>�q�>��9?.?�R0?�,?Q,+?~�a>�D�������Vؾ�?4�?�C?G�?�k?����q7Ľ,㗼�[�Bly��h���=�J�<�F׽�Xs�9V=��T>VQ?Ij�G�8�����k>.c7?d�>!��>B���J�����<�0�>x�
?��>; ���r��d�
U�>E��?n����=�)>�[�=�f���Fʺ9?�=��¼�Ñ=���w�:���'<�$�=	A�=(�t��۹2��:��;��<t�>��'?�?�>y�>F'��I����P��<=��z>-�=�Ľ?�����o������{�-FB>�F�?>��?Z�\�p�=�v��%��\K=��T^�~�=�*?��?�bK?��?�?�π?�F�<�[������������s�ۣ?v!,?��>�����ʾ��։3�ם?h[?�<a����;)�א¾��Խ߱>�[/�f/~����?D��򅻾��m��4��?�?AA�X�6��x�ٿ���[��r�C?"�>Y�>��>Q�)�~�g�p%��1;>���>gR?I�>j�O?�:{?��[?�T>��8�<!�������.���!>��??J��?��?w�x?�H�>{g>��)�$ྰ4��P��#�ɂ��W=�Y>�p�>aM�>���>��=U�ǽ�ԯ���>���=�zb>���>>ٶ�>JVw>kc�<C�G?��>�6��J��.Τ�r���O�>�Lbu?��?q+?�=�x��F��)����>�n�?l��?$0*?F�S�߶�=�gּ>ﶾ��q�O#�>��>��>��=e4G=�>���>e��>������s8���N���?xF?�N�= ƿU�q��p������e<�����d������*[��]�=�������ͩ��[�m����~��S뵾������{���>���=h��=���=���<@�ȼI�<��J=0 �<��=�p�ĝl<�9��Oһ�ˈ���y7[<CI=}�����ʾ}D}?�1I?��+?%D?�w> �>%}*����>������?�W>��K�A⻾�J:�u먾����9Vپշؾ��c����W5
>��E�pq>��5>���=�c�<���=��u=v{�=!B����= �=�ݻ=�g�=�r�=(�>�P>y2?ƈ�艨�X>P�c���gR?���><�
>�����q?o3�>����[7��{~#�&Hp?S��?�A�? �(?�<P�)�>�!��ZHY=���=��{�\�=Z��=/Խ>�X>q%�F��}�Q����?�a@\!?:D��F�пNg�=��'>�!>��S�i{���������'+��@!?+�L��\پ&�t>#�s<�� վ��;=rsN>`�=�'��c�G�-=�{���5�=��=��>�F?>�Y�=e�x�~�1>n��;d|�=\� >��I�q�����ɶ\<�F<Y�>�&�=!��>ߺ?�%3?��_?��>H�A�2eپ<`Ծ��>|��=`��>E�2=�>�E�>��1?�K?N?̲>�ې=�1�>wo�>��*��9q�־�᪾�cO<;��?�?<��>����-��;��_=�kwݽ!�?�#/?5K?'L�>�D����VR�q�I�^_�����~z9>�A�� ���B%��{0�6X=�54>�
�>��>n�>�r>	y�>y�Z>���>��>>�g=>8=�=�ӏ=T,�==JT�H��|}=M�����C�ރ�<
+�\k��a˽�H����=<b�=�dW=�O�=���>���=z��>���=V�վ�Y9>=$���aV� �~=4���ODD�g(`�?�{�,'����P>߽P>]�ݽᑎ���?M�f>�%.>���?�j?�o>[� ������ܛ���Y�tT_�HI�=Z�=S�O�_�7�Nb�DyL��׾B��>bߎ>�>Ѽl>�,�Y#?���w=h�Bb5���>�|������'��9q�"@������Ui�WҺ�D?qF����=
"~?��I?.�?���>^����ؾG<0>lI����=���*q�)h����?�'?l��>��T�D�]⾙ӌ���>7难V/d��7����@���= ���H0�>}�l��[̾U���쇿&+��+M��؜�y?�\?y�?�G�Ǆ����Z���'��d�=OVK?��s?>d�F?�t?#$�e��"�ɾ�\��tm?Pg�?�U�?��+>	��=����V?�>�)	?w��?���?|s?��?��u�>4,�;�� >\ǘ�('�=n�>�s�=&J�=�t?C�
?��
?�j����	����@�>^��a�<�¡=��>�n�>-�r>V��=��g=(}�=�\>�Ӟ>'�>	�d>�>L�>n��U��gR?Vq%>I�>N�D?���>>�8��6���q������fQz�n��B��g
:R��9,ܽ�0� �>#vп=��?C��>\0�rZ/?�:۾o���(�>':D> s�#��>`j+>���>:�f>END>�v>��	>ԏ>^=۾w5>�H�B �eB��)U�
ݾ��{>���~ %��(��*��#B��������@�j�k
��Q�8����<���?ڎн�oe���)����]�?[�>]�9?�
��8t ��j>���>���>�:��=�������+�W�?���?�v>hР>�%w?��9?����H�>�\Z��ӧ��7=��蕿'l ���w�
��|������l?��?��?b��=vnq>[p�?H'��k���u>�s���@a�L���#�>Q���ٽ5����龽��=�<�Q~?_�o?�8?t}�Yt+�!�>>7�H?��+?7	�?-0?�8?����X?�$_>��>�~*?d�D?�rK?'?�Ъ=f�=���[�<�MȽ	�~��HȽ�ʽ�7=�K<f�e��R�<���VV=t�=8���}���=�;C<@�)=�>g>��<>�t�>2�_?^2?���=w2+?�{�=��`�Gd!�-?��
�0	��HȀ�;���������y?��?!@J?��>�
-�����;�<�pP>�>>�A�=Թ%>�w�%Xz�n�W>U�P�P'�>-~>�/��b���ǡ(�)�-��.�=�>D=�I�>�hB>� n���R>I6���9ɾߚ>IK[��=	����ϫK��4�w6��� �>`�O?`�?��>�J���q%�B�`�z�E?��?e3P?e5�?l���I
��*���f�z@����>k�$>>E���f���񪿡4/�8+g=�5J>�о�Ϡ�!�b>U���	޾sdn���I�����{M=gq�.�R=��:+־��~�J��=�
>m���� !�^��!ת��J?_k=����jU�J����>�͘>?��>��8���x���@��[��h�=9��>�P;>���o�R{G����g�>��D?�^?��?�~���q�w;C��r��b���	�U?�>Vh	?4IK>l6�=
���>�οd���H���>��>^	��IG�'�����ﾕ	"�.��>��?��>��	?��R?Y?�^?�(?@�?��>ܱ���y���&?l?y?i����x	'�K	��V*��>F?�˾/��>���>��?"�?�G?��B?�K�>�&%���[��ї>Jɉ>5)j�筿�O�>m�Q?~1�>�Cn?�2{?�4>G�#�i�ھ{�ۼI��,�V=�#9?l??t..?˄>�	�>G�`�9�Z=��>c}?�و?��a?<�>,�?���>CS�>V�c��IG>���>=1?B`?�f?��4?�Z�>Mo�����M*�<D�G��T�9��<��=�q�=1災�����t=A�=p��;���݃=�Ӵ<����[lE�p�|=�_�>v�s>�	��Q�0>�ľL����@>أ�+L��/؊�ތ:��շ=���>��?���>"P#�뱒=���>zC�>���k4(?(�?�?b�;��b���ھ�K�1�>�B?I��=��l�ڃ���u���g=�m?��^?��W��!���:Z?[�a?!�ھ9=��i̾n������}:?ub?��ʽJ��=,J�?-��?�d?葛��~�Wq���^�h����=9�|>N%�W	J�pa�>��3?���>O^>�������P�I�־�&?�{�?�Ϻ?���?s��=I�w�ٸٿ���{����l?Z��>	Ж��F(?]�V=��d����s��f⾛x��Cr��R�_����E�9�V�{��;����&=�1
?�c�?��d?�/o?������q�E�b��zp�YyW������RJ��w>��TC���i�ot����쪾`'=�ZA�iYs��?:Q?e��y8?�l�����䦾ǙP>����]<�#�=�="��=�Ӵ: " ��۹��¾�c?��>���>P`j?��G���R�P� ���#��d���D>:c�>��>m��>I�=����9h�I;��X����b���>�LV?ʓ
?��s?{o	��D>��z���L��=��JŽZb=6cz=Cc�>�\9>X��=ػ5�)O�3��Y9��Y��� �X �=�r8?DȺ>��>��o?m��>^�/�B�����>�$]�bm�`ќ>dn�?��>��F>/��t1`�f��>h�l?ɦ�>r�>�����i!�D�{���ʽ;R�>��>�W�>P~p>f3,��\�-n��銎��9�+�=`�h?�k��m�`�V��>�Q?��e:<QJ<y�>Uou���!�:��^�'�]�>��?Sg�=�;>�ož��H�{��;���u'?R9?ȱ���	�A+�>�M7?��>k�>;Ҁ?b��>�f���G���?߫J?��B?UY?"��>pZ=3%����|���O>��>b�>j��=ߋ�=����5C�mƏ=-�o=��<�'�M�@i=@���ǧ��Q�=��>�ܿ5JL�
�ؾI����o�˜��G��V��ܩ�9泾^���ѭ����%�c���sM�G�o������g����?0��?����<M��#��X���JQ�����>�8\�I&-�Hݡ�����z��w���� ��*M�ݒe���`�9�'?�����ǿ�����:ܾ�  ?�A ?��y?��3�"�C�8�s� >�K�<�2���뾷�����οͦ����^?���>���0�����>]��>�X>�Iq>���K鞾�*�<��?L�-?v��>�r�&�ɿe���mȤ<���?�@V^A?�:)�`�뾜�Q=Y��>s�	?�A>��1����̰���>d4�?X�?�sQ=�W�
�	��e?�,<F�F�WIѻ���=7M�===���"I>#Z�>�����A�k�ڽ�}4>��>C3$�����O]����<1�\>��ս�B��2Մ?3z\��f���/��T��"T>*�T?�)�>�;�='�,?T7H�F}Ͽׯ\�x*a?�0�?��?T�(?8ڿ�Hښ>n�ܾA�M?oD6?���>/d&���t����=�:�0Ҥ�F���&V�6��=��>V�>�,�E����O�D@�����=w2���ſ�����J�>r�>��������ϽLv	��U¾���\j��[���J >�n>�+�=?h�=�_>�kM?�j?��>�ާ=e$A���S0̾��T��R�ʃٽ�����ný���|]
��۾�`��]�r?��l��� =���=�3R������ ���b�e�F�"�.?pt$>��ʾ��M���,<pʾ�Ǫ�!���諒j1̾��1�n�P͟?��A?y���� W�>����f���̳W?�I�˶��Ԭ����=Z5��b>=@�>f�=���y3��zS�X3?�?%?x��Lx����#>R��m�<�� ?��	?d�.<��>�k?��2����~f>�L|>>D��>�5>������Ľ��?��O?��h��B��9��>��ɾ�y���)�<,�=�Z��2�:k�}>�<=��}�k&���ֆ�
�8=-�W?�ߢ>���;�>y���]�u��<��n?1h?�h�>��f?_q7?ޑ�G�����G�u��h��=�Z?I�s?յ >W�k��7پƩ����7?��]?~�7>�~�}w��[M<�rd�_�?@�m?C�?�3F��k��������w/?��u?��3�
촿�"��!��f�x�T?2W?U���As�="�W?\J>Ս��SO��(�^��ă?��@�z�?b�<b��<k�?�:�>�)?����C�ξ�,#�0���$>�G*?�Ͼ7G_��/�Th#�?eI?��>Y��ᾖ>>,���¶?^]�?ɘ��V�����j�h�����Vㄼ���=��ݻ�$\�T�����%�H��y���A��W.佊�Z>��@bN��o�>��+���DCٿY�`�^쳾Yu��<?��>�����v�uXx�p�_�i�K��ӽ;R�>Y�>\�������)�{�)l;������>R�$
�>��S��������g4<7�>.��>���>���ν��?�T���=οh���&��̵X?�a�?<m�?bh?�6<L�v�c�{�8}�HG?ws?�Z?2�$��H]���7���j?r9��k{`�Ʋ4�΃E�89T>�W3?W��>t�-��u|=$i>��>�/>�#/�s�Ŀ�ɶ��������?nb�?�,�m��>Ml�?-}+?^u��&���ة�*	+�>֋�8UA?��1>�^��j�!�G=�n�����
?�0?�[�ZA��_?�a��p���-�ҽƽ\ݡ>��0��a\��'����?We�����9y���?e]�?��?���� #�}3%?��>Ɯ��7Ǿ���<���>�)�>|*N>�V_���u>��N�:��c	>��?�}�?[i? �������gb>��}?�M�> ��?hj�=��>��=du���iP���">z�=Lg:�kh?�M?ɫ�>�a�=��6�'/�ntF���R�AA�a�C�Rr�>c�a?��L?��c>�O��=2��� ���н�1��Լ
RB��1*�Z ߽��6>��>>Z�>�C�s]Ծ�>?ud
���ӿq\��lR���o?v_�>h�L?�0��"�����>�\?���>"���K��������+�?"J�?w6	?�`���焽�(�=�t>5k0>�d>/�^�����0�(>��2?&�Rr��
|U�;RO>���?�@�?�kv���?d��m��� 䍿1K%��-}��-�>�fL?yr0��$
>&t#?Ig>|�h�(b��͡��!Q�>���??��?���>��`?��V��?C��m�=���>f/?�?W ��%�;V�=�c�>J;��Ě�c���ZI?#T@�@Pi6?�ۜ�`�̿���I���!8���>>�TP>��p>�3J=?�=�u�=�o��f¼���='��>/��>��>'mF>}�=�-�=[����\Ɣ�/lx������پ������?1þ��s����ή��2̾Ɇ�AE4�i�J�����ˉ�=�>�lI?��;?j=�?�?�Bս�bC�=���{��e 쾦�i�'=MtK?NG�?r�?n��E��#z�����������H��M�>�;�=��>���>8��>�u��>�>�`v=���1�>Gʟ=eO>��<$�]>^bo>R��>>�C<>ґ>Gϴ��1��T�h��
w�`̽-�?b���W�J��1���9������i�=Gb.?l|>���	?пg����2H?���s)��+���>}�0?�cW?��>��P�T��9>f��b�j�I`>�+ ��l���)�&Q>xl?8c>j~t>c�2���7�ՌO�r���4�z>��5?�a��,;�k�u���H�S޾�M>eݽ>C�P�����f<~�X�g�֊~=��:?h�?�೽tp���)w�EI��{7R>l�\>�=>*�=�sP>��X�%�Ľ��J�ɒ"=���=��c>�?P�]>x��=�d�>�r��?�Y�?Μ>��;>Wqt>4�G?@)'?��8���
��ב�<��q͓>�f�>���>�U>��!�L!�=���>��b>�W���l�a��,]H�<�@>��
��<��i���G�=tr���@�=�C�=N9��}g�
�K=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>Q�$3��^0���l���x�C�>�g�?܊�n体0�;Y9?^a?!������Rɿf)b����>3��?.�?�T�߁����V�� �>�(�?6n?��>�� F��e�>��J?i�e?�w�>�(,�ڦ�^�?~��?;�j?Gl>�?�%e?J��>�߹���N�쪽��V��o�t>�wL=�k�<��>� S��T�k�������l��h����>��=�U�>�Eo�=����Ф�і � �����=
��>y��> �?��[�>V0?��?x�.>C�k�!�ݼ趑�kNB�[�K?�0�?C�	�k���=�ˬ=��\��?�c4?�����d;/4�>�3]?H(�?؅Z?�Ú>��
�:>��뱿��F��j��<�^L>m�>4�>�Gv��L>�־�=���>��>M���Ӿ��z�񘡻 ��>��?1C�>�:�=��?<$?|�s>�ó>'RA��뒿�/J��b�>:�>�X?.�u?�9?uX��c0�3���$o����\��ZE>�rv?�w?��>�w���:��m��Jgn�	r���u�?k?�y½�W?���?�/D?!�A?b�D>!�)���о������>W�!?1�
�u$B�%�b�	�� 	?��?;��>K����I׽*Ѽ-M��:���?�[?�Q'?���|`���ľ�&�<�����P����;�߾��p> >{t����=B'>�N�=v�n��4�@�q<���=��>�v�=��/�	���\1?�U�N���nf>8�����b�S�>�X\=j��h�?\��%?B�����Э�������n?m��?X�?�П�mk��?�-�?La)?0�?��E���%����t+$<!����#�I�%;�{�>����낁� 5���~����f����a��C��>���>�!?- ?pu>�H�>����<�^n����NFZ�n���2�e".�#���#���槽&4�4�žE�u�S��>b��!�>n�'?��^>��{>���>��輲Ș>Ly1>#�>� �>�@>��&>w�=Yx�;��D��KR?�����'�1��ڲ���2B?qd?a1�>�i�񉅿�����?���?;s�?I<v>"h��,+��m?/>�>���q
?<S:=�.�:�<�U��)��4�������>�A׽� :��M�mf��j
?�/?�����̾?׽#f�����=��?^�)?�m��R�ުo��8U�{=7��:��|t�״o�X���V�|U������օ���!�Dx�=��)?O�?���+��	ѯ���m�Q�U�pBM>�?���>T��>-ٻ>�ҾH4.��Kh��Q0���O���>ϙ{? �> wK?��&?��H?��X?��>�q�>R���y?��=�`�>�ݸ>NF1?�9+?�<.?�T?�.'?�f>��������Ѿ9J?�`?�m?�.?���>��x�t���mq=��A<����kP����<8M+="�ݽ{C����4=@k�>uX?���%�8�����]k>�7?�~�>���>���%,����<��>?�
?]F�>L �}r�xb��W�>i��?g��Zz=��)>n��=E|��� к�_�=U�����=�/��rx;��p<g��=C��=X{t��삹���:̓�;�}�<py�>�?7Ŋ>�׈>섆��� ���k|�=��Y>�`T>r�>�+پ�������g���y>et�?��?y�j=���=$i�=Tn���V����������<��?+I#?�T?�q�?c�=?28#?i�>�.��-��{F��.���?s!,?��>�����ʾ��Չ3�ڝ?g[?�<a����;)���¾�Խб>�[/�f/~����=D��텻���Q��5��?�?OA�V�6��x�ٿ���[��|�C?�!�>Y�>��>P�)�y�g�t%��1;>���>mR?��>L?K8q?c?�j>%�6�؎��.��U<�5_>�<?��p?�̐?�|}?k��>&�>�cM�xG�K��x�(��~�Lt��aQ=�!E>6X�>�i�>�>���=����6�
6:����=?>df�>�X�>p�>7w�>gEݼ��C?9�?�������>˾$������]?���?�H?1�>	��O�������>c�?=˥?��??+'����/>ʲ(=�$��W�e�x�>nɜ>uu�>~�<L˒=�7</�w>�e�>2��c��Ss/��:k��>c�$?��>��ſK�U�(����V���M>���1��5�ǐ�=|མ�վ�x�����+���2���;w�g��jþ@[���D?�*�=7��=���=Z�нk�ʽ}ݽ`���ݼNF�<}M�VH;=��<9%��TZC�5O$�����e��;	f�=��˾xi}?�%I?�u+?ȾC?]$z>�>��4�ܕ�>?���"5?F�U>ppP�s�����;�����m��xkؾ�D׾p�c��۟��_>�K�5�>w�3>~��=沇<˳�= xr=���=%.F�k=|�=2�=v�=��=�z>�Y>�6w?R���4���z4Q�yg罡�:?5�>�u�=Fxƾ�@?M�>>2������b�,?���?�S�?�?n]i�1e�>,���莽:}�=�����<2>���=W�2����>��J>����J���h���3�?��@�??�����ϿB_/>��;>:�	>�UT���0�ǟS��~X��sW��!?`�7��ξ>{�=پ^þ��A=E�C>�1�=��ٟ]�ͩ�=�o��v?=S�Z=o�>oG>�ɽ=����k�=�hv=���=IgF>��q;�i"�N�/�4�=g��=7su>��+>���>�?#� ?�pZ? `�>�/e��aӾOR��&�>g�=���>�#�=�{g>%�>�??��@?@n,?�5}>➐�_$�>LF�>#�2�%8_��T!������g=8��?��v?64�>��;>`���9�)�d�]���Ö;?{U?k�>4֚>I��ĉ⿙q�(�%���+�J��=��X=��4y���o��R�l��ul�=��>c,�>/��>e�L>��>�Z>3b�>��>�&v=�v�=�Y�<�j=�)<��$9�[�9^غ�VB��'����Ӽ�Z��O�����05�3�<�=4��=���>�wD>��>h��9�1��Z�>�N��l~E���#>�����I,��o]�z�}��g-����U�H>�&�>�8��������>�R�>��=���?b.�?�<����н�\��l����!�cJ��Ym�>�f>\����,"�n�h�͎@��������>e��>���>�6m>�,,��0?�>�x=Q⾧f5�1j�>^���A����?Cq�.3���֟�E�h�����~D?)M��S��={H~?a�I?�?�U�>1�Xgؾ�<1>������=J���o�G����?��&?ɷ�>��q�D�V�
��W��}�>]���5l@�YN���y)��(=��g��+�>?�u�����w�C�d��^]�����u}����>j�Z?���?�'��
p���^���)�V����>��g?�M�>��?<m?a(�?�ľX�U����<�
\?���?���?��>���=ꓗ�_	�>���>ٔ?A/�?]R_?�lW�NL�>M=V�<>���H
�=���=�;-=��>�?�h?�l?����q����Ⱦ`�	��(���>�>&֎>G��>��c>���=�=���=��d>�8�> h�>��S>셈>���>ԥ���!'�Yo??���޹�>QSn?���>lv����<u =iǽ�gս������+}<���=X�=� W>�c=*��>�-ֿ:n�?4�=�a
��N?�$�(�X�.�$>��!>gM��?xM>(��>���>��>�$t>|�=�
�y˾e> ��R� ��8��1H��~߾L�>�d��$���h�쾨�
��}5���ʾq��s|g�o{���7�-ڴ=�B�?���Zs}��jB�tEP�|�>"�>�#Y?�������F{�>�?6�>���������F̮���?b�?��c>O��>y�W?�T?/�1�N3�(]Z�ԧu���@���d� �`�j������
��\���`?2�x?qzA?��<��y>}��?��%�.���kq�>��.�,�:�LU:=U�>[6��ʑa���Ӿ=oþ�����G>��o?��?�L?DV��m��'>��:?��1?�Rt?2?�q;?m����$?��3>�I?/L?�B5?/�.?c�
?,.2>��=�З�U�(=KP������н��˽���g7=e'}=��(��F<�l=��<��zYּ��+;�.��k�<��9=�x�=���=���>f"j?(��>J�1> �?CY$���-��LǾ,?4��<Bʔ����uȫ��R߾��V>K�?U��?5�U?g��>l�E��� ��h>�
�>C�s>N�@>đ�>�Z�?�����<�J$=5=0Q�=�[�=��b�TþI�n��@�=��%>8��>�Q|>����'>fS��r�y��d>]�Q�2���t�S���G���1��@v�%_�>.�K?R�?��=T�&���a?f�5*)?e]<?KFM?��?t=�=��۾��9�U�J�#����>��<i����������:��:�t>'���Qhc>l�d�ݾ^n���I�cy�ED=}����[=�k�$�վ�t}�g��=X�	>A���v �z=��-�����I?h=`?����S�y���R�>��>��>��D�&�t�L@��Ѭ��w�={'�>G�<>B ���r��F��v���>qyT?�
y?9�?�Kw���k�f�S� �v~��^���3��>E4�>ԝ?>
x=Iy>��]�m�9�"�o�НK��L�>�x�>Ϯ&�R	I��-���MT���ƾ��L=h?(��>a�	?��'?�:?�q?�'?��?���>b��Y�ؾt)2?ޕ�?y! =��K�
��pȾ�?:���>��?������>R��>;�:?H?�\?b�?J8>���_�\3�>p$>b�������G�>���?�޴>�g]?`�y?f�>i+�8�޾�~�<���>獑�Qg?pZ?�@?ƶ�>-u�>_����T>��>�[�?�Qw?X�W?K�=S�>�6>Uk ? �=_�C>uS?tB?Z0Y?�O?��D?�?��=i2{�����V2�=��=^ѽm{�� X=�@1��棾�Ͼn�<<7�=�^½�?g���� i��e<��9ua�>=�s>7��U1>��ľ=S��_�@>�1��+P���⊾��:����=G��>��?���>V#�:��=럼>�6�>���44(?��?~?B);x�b�"�ھ:�K�d�>(�A?���=��l�	���w�u�Eh=�m?�^?��W������_?��j?ʆϾ��=�)Gƾ]������?f`$?6s۽��3>?�^l?�7?QP����v�����fr�������=�r�>!����F�RՅ>J0<?hA�>|�D>@"�3���R�F�@�¾V�>�ے?}ʮ?*\�?��x>ǥz���ٿ��Ѿ죥�Yv?U��>�v���_"?ʂ�=���Lm���:����u=Y�QM���-^�.�`�\S�ȑ��*샽�t�=�(?��w?b�Z?�n?Z����c�\�n������U=��d�,�Ird�/fJ��7��i��d���E��5���*;�fx�T�H��?��&?�f,�X��>Kf��~��m�Ⱦ� I>σ��_��+�=�n~�|=�;`=0h�]9&�\"��Q-!?�"�>+�>�d@?�]��*>�Q2�As7�7G��=6>\�>j��>!��>� ;{�5�� ��˾�'��N�޽x��>�5c?��3?O�j?Wpb��X(�a���+�:�漰�3�E��=���9��>Tߕ="����0��j(�G����9V��f�������=��/?&ܢ>;�B>+�x?I]?Gi�,��9����CD�<c��=ţu?��?d��=PQ��@�񾬺�>Y�l?"��>�	�>|����[!���{�(�ʽ/�>��>��>f�o>9�,��\�#k��Ƅ���9�	O�=�h?뀄���`��܅>�R?Nz�:�OH<<~�>0�v���!�?���'���>�z?���=��;>�xž` ��{�><���I6?�p,?-���w�)��� ?M}?���>���>	�u?gs�>�c��R����0?�HT?�#C?I�>?�5�>�ʂ=#^S��%�vQ���8">?_t>�G�>�@:Iϕ>���Osl��^l=�֖�R�>7oc��C=���=�ܥ=�ʽ	l>��>"fۿ:K��xپ����7
��숾���?_��ޙ�k�������x�����t'��HV� Gc�����Նl��}�?�-�?�}��$��!����������W̽>��q��`�oҫ�:��D��e��N����k!���O��i�l�e�L�'?�����ǿ𰡿�:ܾ+! ?�A ?:�y?��9�"���8�� >GD�<y-����뾱����ο6�����^?���>���/��O��>ӥ�>!�X>�Hq>����螾�/�<��?;�-?#��>Ɏr�/�ɿa���z¤<���?0�@�}A?)�(����`XV=O��>�	?%�?>wr1��=�߰��1�>�0�?���?��N=νW�sw
��ze?�I�; 
G�޻��=�7�=�=����|J>�T�>|M��A��ܽ2�4>�ȅ>"	"����d:^���<�c]>�.ս�I��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=p6�����{���&V�~��=Z��>c�>��,������O��I��V��=����@����� �f�%��w�=�m=5�>~��j��=�<y���4��P$�&�^=���=��O>�?0>�T.>҆q>�I?��b?#��>��%>�Q�� �������w�����s����K��ǩ+�@��tﾘ�������r�'���;��!=�#�=�6R�c���?� �a�b�[�F���.? w$>?�ʾ��M�n�-<~pʾ7����܄��᥽�-̾�1�'"n�f͟?��A?������V�]��cX�����[�W?qP�ʻ�aꬾȣ�=����b�=%�>~��=���� 3��~S���/?��$?v���^��V��>����=�
*?��?
e==���>-??��<��+̽ǈ>�eu>Ԛ>���>��>����}	���)?�R?A|E����T«>?C���>���r�<m�K>W�ڽb�ý��p>��=��|�3���Q����g=3(W?���>m�)���e`��`��>Z==_�x?��?%.�>V{k?��B?�ߤ<�g���S���ew=��W?�)i?͹>㉁�1	оށ��s�5?�e?��N>�bh������.�?U��$?#�n?F_?vt���v}�B������n6?�9�?�1��	���ƾ������=�3?��?QP��XO,>/h?�$e�_���ϿM>G��+�?k�	@�@��>��m;����?�q1?1��
W���c��{쾊��=��M?_�Ⱦ�y�#B�ҏ����"?�b�?�P�>7��Y���o>�2���ݭ?�L�?ڱ���	���������:Aʾ��0=�2��_"&�^&�"_ž�|1���㾲P$��׎���<?s>Z1@�|i�ǋ�>K[ ���ڿ���=��yL ��<��-i�>�Y�>����Ǿ�\������TS��6V��Wl�/_�>M#>r��˿����{�za;��ܠ�*��>}��ֈ>v�S����Xe��$�5<��>?��>���>j��������?n`��5Hο�������X?e�?,`�?�w?'�=<��v���{��B�=<G?�vs?;Z?K�"�\]���8�%�j?�_��zU`��4�yHE��U>�"3?�B�>\�-�"�|=�>���>g>�#/�x�Ŀ�ٶ�&���\��?��?�o���>p��?ws+?�i�8���[����*���+��<A?�2>���M�!�A0=�RҒ�Ƽ
?X~0?{�h.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>`ք?�;> _?���=ṾCXJ�Zr*>w�=�m཯��>�II?�(�>��=��2*�=:J�U���	��?�Y�>qe?31I?.�Z>��ý4�p��! ��f���C���"��k�ݝl�� ���!>8I>���=Gp5������.?����Y�п9���aW���z?�8�>\l6?�98��h�_m8>׍y?n��>�&��ᶿY)����)����? ��?��?�r���랽�L�=m/�=]�C>�,�>�����龩�=�jP?4h/=[r��
���$�P>4��?. @4˥?�|��5?���te��1ɀ�d.�\Ke��Ś>fcE?��*�ޥ>�!??�>��j������{��J�>���?�0�?s�>j?HZ]���8�@�>g�l>gU?y�?��_�価;t>X?���o���S��Y^?'$@�@N@u?�S����ӿP᛿����<߾Y��=�"Z<��L>�o�;8�>�rĻ� >5��=��2>�z�>���>�ٜ>��#>��I>��>A �����Ǳ��r���^]�k������&ɽsЏ�6;�Yt�?!���]��S6�Xԛ�O���c�>���vP��%>� W?x�S?��?(U�>�~ �|Hb��ľ � �R\��>^�=ҩS>�l8?"�'?�;?p-p=Εξ�p��0���!���nM���>�[>.��>;�>gn>�j�V�J>��\$6>���>� F�e�w�H��;�h�>�R>j��>� ?�C<>��>Fϴ��1��k�h��
w�r̽1�?����S�J��1���9��Ӧ���h�=Hb.?|>���?пf����2H?&���z)���+���>}�0?�cW? �>!��s�T�4:>:����j�5`>�+ �~l���)��%Q>wl?�g>_�u>dD3���7���P�KI����z>ޡ5?񁶾�x7���u�-�H��Oܾ�O>���>��]�>�H��ȏ�4i�
{=�D:?f�?ӵ�����u�K[��R+O><\>�� =�S�=��M>�Hi�pI½xH���)=���=K^>?�k,>��=���>铙��O�չ�>oKC>J�+>E#@?�%?���<���|�����-�Rx>�+�>R�>�>�K��Q�=�D�>��`>K��ƀ�����?�X�X>|�~�_�]�y=n�̲�=հ��h��=|C�=u��u=��x$=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>�$ �p�������Lv�tq��Ց>WI\?p����>���Ľ4�?E�?����Ѧ�ֲӿ�M|�}��>�a�?%(�?�AK�%ʞ��3_�7�> ��?{�q?��>�a"�k�ʾ9�>�&S?z&`?��>ږ!�R\���?%�?��?\m�>��?�0l?/�>$���*F�\:���8��U�>%�W�W���>M$^�����)��Zk��hS}�:�'�؅2>��=��>��e����՗`��b�Dy��d�=
��>�\�>��=Ə>��?s�?��H>�9L=��=�ؾAPȾL?�Ɋ?�D���?��j2�څ=�½����>.�1?��=�?�;�`>�\?��?2<5?t��=F8Ҿ�ݥ���ɿ����L_ټ/�,>D�?�3�>�V��e>���X�ž�>ꝲ>��Ƚ9���������;>�w>��?���>��j�\4 ?��#?��q>摱>��C��㑿��G�֏�>�>�>t�?�y?P�?^����2�E+��=U���P]���G>l�w?��?2E�>���Zx�������2m��Ҳ���? tk?����
?4X�?�A?�:A?�Y>���<վ�=|>��!?�R�׸A�oL&�\��-	?��?���>�g����ֽ�ͼ!$�;����0?T�[?/7&?���`�`�j�þ:X�<����r����;�� �>u�>2������=T:>���=�6n�6��#u<�=��>�M�=�x4�Gu����4?�A`�,+|�1��>�����>���=����{?A񽫡]�j���=Ŧ�5�uۋ?���?�#�?RzP�a�}�M.?�`�?r�?��
?E���o��l��������~#�<5��3�<#�>l�P=a6���Ơ�f���wh����#��k9���>r��>���>�u�>�m >X�>�8�40������PǾ�8���Z�"�6�G)��Ծ�dk��P���x>�վ���h^�>ݧ&�`�>ǝ"?�{>�P">�j?y�H�lR�>�/�>�>���>K�>;{3>��g=�A��5'� LR?������'��辎����3B?[od?�0�>i�|���u���}?چ�?s�?�@v>V}h�a++��l?�8�>����p
?�Y:=D����<�T����-��.�=��>RI׽�:��M�Oqf�j
?^/?�)����̾�+׽(�����?=���?�+?�>��L�ͱi�h�_��A��7�e=���흾�R8���b��2��=7��#�|��$ ��ؙ=��/?`ƃ?dg�\��4�վiy���G�o��>���>m�>u��>`>FV��>E�ϖW�4�7�K������> Qt?]z�>�tL?_"8?R;>?Z�e?��> Q�>�g�I�>�.=��>���>$�?��&?<2??�'?"W?�K>�;��&	����8#?B�?6B�>g��>�?{X#�r��-���ւ=��5��,���)>
��=LϨ�����{�L=IG\>aY?C��Ϭ8�;���;	k>N�7?�}�>e��>���D,��r�<	
�>6�
?�H�>����5|r�>a��U�>Q��?C��=��)>���=�D��j@Һ3]�=�����=���N�;��E<j~�=���=`t�[b��C��:\G�;���<t�>�?ѓ�>�C�> @��� �׵�i�=�Y>uS>>�Gپ�}���$��V�g��^y>�w�?�z�?��f=~�=)��=�|��.V�����K������<��?�J#?�WT?h��? �=?�j#?h�>A*��L���^��Q��n�?#!,?\��>�����ʾ憎�3�<�?�Z?D:a�����8)��¾��Խ1�>4T/�<,~�����D�|���(���u����?C��?��@��6�0y��Y����C?V�>�^�>��>��)���g���C!;>Ї�>R?��>.�R?!7f?"LO?�<�=T)��^���s��2]=$n>y?�X?l%�?�n�?7��>��[<{����x)��n8�s��g�t>]� >+z�>Hw�>���>X�~��۽�K^<g�m����=�>H�?��>%��>io�>�Ӳ���G?��>(���]��mQ��U�����>�X}u?���?YF+?�z=֟��lE�`����`�>_�?��?�*?S�T�Fc�=vvռ�򶾫�r�׸>��>��>���=�H=�w>[��>��>�����i8�5FN�n�?EF?]��=�W����G� �@Ŝ�)c�=Y%�(���D�X� �J�6>@���7��x���<����澬���l�־1h�����N�?X�>��\>�nq>Aq(�����J��� ���y��M��!@���
=�F7�н�k���n�)>�=Պ�=(	�� #˾ۖ}?7pI?Q�+?ΜC?rx>ܘ>��2�GK�>�݆��?�V>8TN�����Kp:�z}��������ؾ��׾��c�݃��k�>&I��>� 3>WI�=�<���=�t=Wz�=� -���=q%�=���=��=��=�	>@F>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>s��=v�2�T��>��J>���K��D����4�?��@��??�ዿТϿ6a/>=h8>�>=�R���1�xn[��]`��Z��!?�;�Z̾E��>#��=M>޾��žhp0=-7>Aze=�k��j\�;v�=��y��::=YVh=���>
�D>�x�=�쮽t��=y�N=��=x�N>�薻+�4���-��@2=|A�=�c>�&>[��>��?>T0?vPd?�4�>��m�/%Ͼ�5���B�>��=;M�>Z��={�B>��>��7?i�D?��K?�W�> �=���>���>֜,���m�+�����Z̬<��?Ɇ?J��>-S<o�A�a��.Z>�HYŽ�q?0T1?ns?:�>	8�u̿��}�;�w�7�ǽ�Y2>�^�>���>�W>A��=�4��uu�j,�=��>Ao�>�ְ>ݜ>a#3>m5v=�͖>�Z3>�,>��=�>� �=�d�f�Q=w�����=�0��XI���I��[��1��T���y��	���Aֺݰ�=�a�>�mA>y�>y�.;�} ��(\>�Ak�B[X�s)>#b���U����F�����5��#p����>�>��=����w��>G�]>��@�\��?E.�?��=��=N��8|����ͽ�����:r>ኚ>�f��M��h:g��=\�0r����>���>Z�>X�l>9,�|#?�`�w=L�b5���>:{��2���#�+8q��>��,����i�ʹԺ��D?VF��-��=�!~?¯I?��?��>d���ؾ7=0>�M����=)�l*q��y����?�'?ѓ�>C�q�D��J̾����߷>5I�=�O������0��8�~˷���>�����оj&3�xf������B�gOr���>��O?�?4b�X���RO����NF���m?,�g?��>LH?�C?����j�kp��(`�=2�n?���?`;�?�>���=�Չ���>2?�˗?�^�?��r?�;*�@�>~�<
�&>-Ҳ��E�=�j
>���=�?>�E	?�?��?�����
���ᾜ��J�^��=��=c֏>e+�>�R`>V��==���=%j>��>�;�>�X>�>��>�r���$��C3?s`=A�>Ư2?�/�>��~<���ƼP=�w�e9>�=��Qm��]~<(=>�A�J�> >?-�:�?1\k>ސ�3v?:�~/F���N>��2>+���h�:?�5>0��>"�?H>R)O=-Rt>E�̺�Ͼ��=����y{�p�C��RZ�,�<�|>�虾���^���)^�������w�}���z���+����=��?b½Tq��Y|9�{�o�g�>ˁ�>��e?�=��Ȅ
��>JZ�>H�?i,�Dڗ�i���	���9:�?��?;c>��>B�W?�?��1�3��uZ�C�u�\(A�e�T�`�|፿�����
� ����_?��x?yA?�T�<�:z>A��?��%��ҏ�o)�>�/�%';�5B<=I+�>*����`�L�Ӿ[�þ�7�DIF>J�o?'%�?NY?�SV��㙼��%>k�<?mV2?T�~?xT5?�@:?/�ýU# ?�> ?Q_?A�)?=F0?��?�fl>&��=���< r�=I=���:��q���O��=����<ȸ.=����	;b s;��F�$����<'Q<�*�넘;��=���=婽=G��>ȍ]?� �>9G�>��7?�W��7�0����.?�r>=o(��"�	p��1��>C�j?Aǫ?�Z?.�d>WB�tC���>�߉>��&>��\>���>{��)QD�{U�=�>�2>֙�=%~J�@π�[�	������Q�<x*>�L�>��>Z�u��79>�7��8h��vrS>��F��ߺ�� h��D���1�|'e����>��M?�?�ct=7NﾬѸ��d�k�'?�*>?��K?)n�?��=�ݾw7�A�F�}�6����>�=�U
��餿m���5������l>Y��\ꟾ��d>~�ә޾K�n���I��辞�==���U�H=C�
���־v]}�}�=�q>����3� ����n��2�I?��m=�����U�S��~W>��>Jۮ>��8�駀�,�@������L�=��>o>>���_��6G��A���>�e?�K?�m?_a���l���D���F�Z���'����?N��=O� ?U�>Mk��i��}	��a���n�χ�>�[�>���ZNQ�@���ܽ��B*��.=`�C?���<^�Q?6�?�r�>�MB?�*8?�?q	�>��ݽ��.�'?�a�?j_e=齺Ik��h4�5;E����>�6,?m�R��̥>H�?r�?*?��R?�?�>5��tH�r�>�9�>�W�1��d�Y>ŹH?n��>nV?�˂?�r&>��7�8w���M��<4�=��<>��2?=D ?/�?TǬ>cx�>_�۾�4�>}l?@pt?�?'�m?�->��>q.�>�F6>�n>�ʿ�>��>�QJ?�uS?`O/?�L'?��>�E><Z,3����u�;���#=��c�=���>�1+���5~.��a�=q�*>a#�=�O۽HP���;�?��h<��>��x>�"��� 5>��¾3{��ų?>�ا�U ������R,=����=j`�>�H?���>(�*�Rh�=� �>���>×�U�'?�?��?<�H<�Ob�dؾ�N����>�8@?F�=Om����E�s�?�W=�m?H^?�U�rJ���u?�Pi?b��gw��������Emh��S?H^5?� ��4���i�?qq?\T?D �ox~�I뤿@���	��<��=�*>��������=V��>9@�>�Jq<��Dد���X�iPھ��?��I?W��?ѕ??ns�>W�V��'ٿ�V�|떿�!a?���>I���t?�7�<��Ͼ�����։���޾�n��ͥ���|��󠾉�*�݈��]-��l�=D?��|?��_?%?_?�"����g��d��"q�S�[�,��4g�,�?���B���?�Xs�"4����Ჾv�{=\�q{o�չ?�?X�,����>|�`������&�N>A���3�ѽ'��=ut�<�Ę=u�=	4�6Z���N���e+?Z^�>l�>�TU?�k\��VE�3[+�e��|'��">���>�Ou>���>�	>�?}�؁��AᾫM����� �x>ԫc?,�I?ɮm?1� ��2�6/��ϸ �7@�p��,�9>�
>���>��R�T��'��s>�[/s��l���q��(�=f�3?)��>n˘>4�?�/?��	�n���)r���1���M<)?�>��h?�-�>=�>ڔɽ�"���>��l?x�>�$�>�Ԍ�5!��|�O6ɽ)i�>���>��>8{q>�y+�D�[��p������&J9��)�=��h?K}����`����>	R?�O�:�XC<��>��x�?�!�����'��>E}?0�=�y<>�žh���|{�����S)?`\?撾m�*��}>A!"?]p�>�>�0�?l��>�!þ8*��|�?x�^?-VJ?�BA?�>r^=uS��3Ƚ�&�_�+=r��>�4[>�l=��=|��W\�_���A=���=چμ����$=<B���B�K<���<524>�hۿ��J�=0ؾ���l��
�֭��ݯ���������"�T��?�x�(��X�+��V��c�d���/Kl�L��?���?�u��q������ea������˻>9[s�\e���o�������-���୾4!��O���h�%�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >jC�<�,����뾭����οA�����^?���>��/��o��>ޥ�>�X>�Hq>����螾Z1�<��?7�-?��>Îr�1�ɿc���o¤<���?0�@{A?��(����ѕU=���>�	?��?>�I1��C������4�>�<�?���?a�M=�W��_
��te?CN <I�F��6߻0�=�K�=9=����cJ>hf�>�{��{A�Mܽ��4>sʅ>"�T���=^���<~�]>��սX���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=`	�������
���q]=�$�����]�ǽ@�L����1*��XU�����k6=y��=�1>��M>V�>�e>��K?�{k?�><q:>[���7����ž��������i����y�M��7��ϴ�����-��
 #��پ< =�>�=c6R�(���h� ���b���F�X�.?x$>t�ʾ��M���-<:oʾϾ��Rℼ�好D.̾s�1� "n�͟?9�A?����;�V����RX��~��ĮW?�O�ܻ��鬾a��=���ٞ=v'�>���=7��i 3�S��}0?`a?꠿��)��7*>y� ���=�+?Ӓ?��S<��>�^%?U�)����8�[>ǆ3>ȣ>�E�>�t>�B���۽��?�T?{-�����*��>�н�PF{��(b=ĭ>yV5�g�ػ[>O�<�2���N��c��n�<�5b?���>	#�w_>������ �vD�(��?y�B?��>��*?-��?&!3>d�þ�p�v�*��"S�� &?�&�?��>c*�X�߾�d���P.?�U�?<Ȳ7�mƾ�?���X����p0?��N?��/?c�սs�X�����H��o4?Ibq?+a>��ſO��?L��r��>��W>C)?����#! �2gc?��������;Ϳ�C�Mu�?F@)g
@���=b�<��ͽӼ�>Z��>�"�! �>#E�se��z�=�%?!3��m�2�5�l�y��X�>Ed?��>м4���>�\ݾ���?m��?5����@����徛�]�9����1<Vxq=����;�A���f*��"ھ���������<��>�@K'[�}'�>rJ�/�޿�ؿ&Z�L׾�R��e�?�S�>VH��p׾�U}��c���\_��qa�(߽0��>>$>�씽�Ȑ�a%}�Q8��9��h�>r�{�_Z�>��'�����Ԙ�Ɖ�<�m�>cC�>�E�>��нV�̾&d�?
9����Ϳ
������>[?��?��?�,#?��A��a���}�k�<�!F?��{?�\?A|��og�3#��C�j?����cT`�V�4�pSE��T>�p2?q6�>�J-�N4~=��>��>��>��.�)rĿ�䶿�&�����?�`�?ft꾚��>$`�?��+?�N�X��W����*��H��TA?4;2>��K#!��7=��ᐾY
?��0?3�����\�_?-�a�J�p���-���ƽ�ۡ>��0�f\��M�����Xe����@y����?M^�?h�?ҵ�� #�g6%?!�>k����8Ǿ�<���>�(�>*N>hH_���u>����:�i	>���?�~�?Pj?���������U>�}?�W�>�b�?P�=`	??�8>�i�� �R��=�x<��<����>7)?iL�>4�(>n�:��;=��D�ŸT���OTC�Jƍ>-j?��??G��>VO���Sx�ɲ+�o����:���+<*�4��gI�t-e�;n=Y�U>� 4>;�%��� �w�?���٪ؿ���i7,�ǩ3?��>�%?R���y���Q�my_?�2�>��,������2���d�?��?�	?�E׾�J�6�>;ٮ>P	�>i�н�ڟ�1y����3>��B?���{=���po���>4u�?%�@��?�Oh� H?��¾�흿�+��oH�V�%�Sd>���?�D6���3��+V?��>�gs��`��K_��}ϻ>!O�?�_�?::?V/`?[�E�qZW�ņ�=�X�>�?%�?Rλq����z��]?i�	������{�gD?YB@1�@���?T$���^ڿ�T��:4��lJ��F:�=X+�="4>��Q=�p�=��Ȼ�� �U�=�X>3�`>�wS>'<>�+.>`F;>���=����i�����D5�Da�%�ᾟ�K�1���ཚ���!��n�Ͼ�<��㧽09׽�;��T��t���m>��U?%N?�߆?��&?�+��"�;>�3��ۘT�T�s=��]>}_;?LYT?(�*?��%<�J��U
X�yB�y��ȏz��J�>��>9��>��>ʻ�>�N<�I>Z�>���>[�=�ӱ�k湽b�T�ɦ�>OX�>Q��>`e�>�C<>��>Dϴ��1��k�h��
w��̽.�?v���L�J��1���9������i�==b.?�{>���?п_����2H?!���t)���+���>l�0?�cW?�>4����T�2:>O����j�`>i+ ��l���)��%Q>fl?��f>c+u>ʚ3��d8���P����&H|>�.6?a嶾�;9���u��H��Nݾ�QM>2��>sF��m�����2
�3}i���{=Dw:?��?/���Êu��B���*R>bE\>�s=�=�=_M>��c�4nƽeH�¸.=���=�^>9O?��+>S=Lң>�T���IP�4��>cdB>�	,>Q@?�%?�+��헽�����-��w>MU�>+�>�F>�kJ��=�r�>��a>���[��������?���W>ii~��}_�+�t��y=����&�=�K�=y ���<���%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�}�>�f��V��+���}v���={Ϳ>�H?���4{U��:�c�
?Ce?M��,���[�ȿ��u�F��>W��?��?sTm�ӂ��'T@��=�>�|�?��Y?��l>��ܾtc]�c��>/)A?S�Q?h �>�l���"�6?���?ܜ�?&�I>e�?:�q?k��>��G�Y�2�4챿c�����M=���;�B�>�n�=a˹�W?������ω���h����#H>�."=L��>��ɽx���}��=��K�؁������C��>۵q>0�S>�>���>��>Dh�>^�"=��~���y��$����[?1o�?'����;�!K���=�����R�q�_?gF�8�g�� ]>��N?H�?�Xx?ļ�>�������N�ڿl���ŽqL>9S?.�!?�'���z>f�
��Z�So>^:�>1c��
ј��Z���)�>��?+�>G��>Z�+?��0?b>"�">
�V�<����Fa�[�?�C?��?��?�[?4�����'��I��k���b|f��==�?�E?M��>G됿W��h��Y�l�F��?J��?ý�>���>�{?e�~?`�?T/�/z���;�"��I�>�H"?'����A���&�vE�Rr?BN?R^�>!��N
�vz��	~�����?��\?,V%?�D�L�a��ɾ2U�<�s���J8�;�'(�~�>�{ >����hֵ=��>�,�=nEh��5���P<h��=��>�+�=�8�ID��e�3?IJ��2����`6>����k� �L>&�m=p�
���t?w?�@q�ҷ��D�����ݾF�?���?�L�?���Ek���8?�%�?�?[0Z>2�9-����5��z�=9�=���`,b>�N?/�+=wҽ�8Q��O7��-ɯ����l�:��^?���>";�>[P�>|*J>���>���������������a�T^��SV��$3���S>R������}NϾ��k�-�>�q��~�>g�?��/>���>��>3���g>ܛ>&��>Ჭ>��>o�Y>o�	>�=	�ͽc�R?�A��3�'����㊱�2~A?S�b?���>��e�����-�y ?���?c/�?J"s>�i��x+���?d�>[x��z(
?X>=��͟�<F���x���ᆽ�O'�ܼ�>��Խ�y:���K��-h��?OA?�di�'˾�(��/¾$�=x;?|$?Y!��co���o��.�!�;����)�k�'���p3�~jH�?څ�ì���b���1�3�=�+?���?�����Ͼ%���q�e��+��I�>�L�>�Y.>��+>�J�>���A?�$:T���<��΅�L�><�?�X�>�d=?g>*?Lˁ?Z?�s�>C��>�ͣ��S�>t���n�>H��>O�I?�SK?	�E?��>\/?I{�=駖�x��oｾ��X?�X6?<�B?a6&?�&�>�Q���9����>�)�1��Ͻ�;�=�%�=��q��^I��_>���>Y?&��Ь8�����Ek>_�7?�}�>���>���u-����<��>?�
?DG�>� �3~r��c�nU�>���?�����=��)>���=����C�ҺOZ�=������=�3���};��L<���=���=�(t����ϴ�:�p�;\�< u�>5�?���>�C�>�@��/� �b��f�=�Y><S>|>�Eپ�}���$��v�g��]y>�w�?�z�?Իf=��=��=}���U�����J������<�?@J#?*XT?_��?{�=?_j#?ѵ>+�iM���^�������?X�0?�x�>��6}ؾ�I���/��(�>��?�X�L���9�Ȭ��;GD���>�/��Ă�3J���
J�ak<9����[��?���?@|L��5D��+���d��(Mξ�E?��>"��>%�?�+���D�����:X>��>'_8?O'�>��O?�({?*�[?K^T>��8�#��Gԙ��G4�.�!>e@?���?��?[y?�]�>�Y>m�)� 7� ������+��ֿ���U=�Y>P��>{�>F��>.��=�Ƚ
 ����>���=�~b>�>S��>���>�rw>�<��G?3��>�]��6��E줾�Ń�B	=�&�u?ᛐ?Α+?�T=G��.�E��G��iJ�>lo�?���?4*?��S����=)�ּWⶾ��q��%�>۹>�1�>�Ǔ=WyF=Mb>��>à�>)�a��q8�QM���?�F?	��=��ſ�=���F�i��ꈽ=!,���Iݾ��H��U�x?��u���Հ�Ė���g��ాG���ܾ��˾W���?�CC>�b>�>���LL��������4���
�o��7{4�#*	��W���P���ӽ�20�g�<�̝��˾�}?�9I? �+?!�C?��y>�/>v�3�3��>�y���9?V>�kP��x��؍;�����#���ؾ!�׾��c�ß��[>4�I�æ>�L3>N�=k؆<�M�=v0s=َ=�)O�k�=''�=0(�=Zo�=��=��>�2>�6w?X�������4Q��Z罤�:?�8�>i{�=��ƾp@?��>>�2������zb��-?���?�T�?@�??ti��d�>M���㎽�q�=Q����=2>t��=z�2�U��>��J>���K��A����4�?��@��??�ዿТϿ4a/>��7>")>��R�w�1���\�n�b�qZ�Y�!?nH;�2E̾Q6�>A��=b-߾�ƾ�r.=��6>^�b=�f�6U\�;ߙ=` {�#�;=�k=ډ>=�C>:j�=�)��)�=�~I=M��=�O>�L��1�7��+���3=&��=M�b>X&>���>��?�l0?$bd?�[�>��m��Ͼ:��Q>�>#v�=�O�>���=e�B>꒸>��7?��D?	�K?�v�>�=���>��>Ӓ,�k�m��k�W���G��<���?Uʆ?�޸>�.U<6�A���&o>��Ž��?�D1?,m?��>A2���Կ�
-�S=:�V�ź~Q����==`>������x�>ٜ_=5���9*=���><3�>��@>�0>KA >���=ƅ�>�*F>Z�@=�=�����<	<�4M�z����0=a!v=�k=���1���ӟ����}�Z�<����ü*��=���=���>�7>z�>��J�Uľꏩ>�Ǿ�A�`b�>f��6�O��y�z򌿓A@�[L۽��>�3>��i��圿2%?u~Y>��� X�?�|�?ט>,c�<RZ���ۏ��%�ف��>�dD��v˽��+��?�E�W��k��E�>��>�{>J�n>�-$�1[�]B����V�?�r�>x�n���Bj)>OY:�ʇ��7��*]g���?��� ?���k�*>�Dv?{�?lv�?�.o=wh>���vu��օ�^��>N�#���7d<��-?C�?���>;]���Pq�����q��ƃ>��e�R�k�>Ւ�z{1�I�=.�׾"�3>`Ō�8$¾U�E�Y׎������T�z灾�r�>�J?3I�?��L�.���o�o�C�<�=׊?f<�?�I>���>�2?��>[�}�B�Y��Alj?���?%��?Y
�>�Ѱ=�����>S�?���?�,�?,�r?�a8��m�>��a=*y>RY۽@��=��>��>�>i�?��?���>&���	��f��w�[3a�B�<��s=���>�>�6p>\�=$�~=C<=�&>p��>å>�Ya>w�>�j�>�	�����A?�硽[�>��?�k�>�dn�7�E��.V=6�`�T��R�x��\W�-�5��#>�>��;>lR�<� ?�翠(�?��>��g��>�ƶ�J�
��ܰ>��~=`hr��D�>8�>~R?z ?�y">�o�j��>&xw>�:پo�>MI�m�B�A��V���־�z>�f����?��A��h	�\?a�XT���#�N�k�|a���Q>�e�<0C�?Ȣ�d�k�H}'�����n?Ii�>��4?�^���P��7�=��>���>� �p��𯌿D�־�?E#�?�;c>��>F�W?�?Ò1�3��uZ�%�u�i(A�e�O�`��፿����
����,�_?�x?,yA?�R�<:z>I��?��%�\ӏ��)�>�/�'';��?<=u+�>,*��?�`�_�Ӿw�þ�7�IF>��o?7%�?|Y?'TV������n���}K?7WG?@�?[}?�FY?D5�<ci�>Xa�>2��>�3_>~�?�_??�P?���>�=���=kNB=بڼ�%a�R���o�H�.����"�x=�u�;��_=FX�<�8��B�S��P���z87��<�<�.=.Ϳ=Cٹ=Й�>1�]?�M�> h�>�7?c��O8�JŮ��/?:�:=����I��zԢ��V򾧽>��j?��?WZ?}Cd>��A��AC�U\>W6�>^�&>?"\>�:�>�1�znE��=�>��>y1�=�KK��b��ε	�刑�,�<?)>��>Y�>S����+>NO�������Bd>��Q�?鼾LS�\�G�'G2���p�]e�>�K?��?ؾ�=Ne���^of��(?��<?�6M?Y�?;\�=ǜھ�:�M�I�q�x�>���<,�
�K���1*���d9��,S;9�s>�ϡ�����G�`>�y�m3ھ��m��J����p+=�)���=_��`�ԾЫ�����=���=m^��-� �7Ŗ��N���J?0CP=�F����X��ۼ���>m��>�ϯ>�V����d�>�U>���d�=��>�K<>�Z��"���ZG�������>E�l?]OL?�l??�ؽ�7����h+��:�gq��v�?���>�T�>u�>ξ~=bh޾-���$d�-�Q���?���>�j*�f�'��c����$�GOq>`s2?�qn>S�9?��<?��%?5�?�Z5?#C+?%X�>q�~������*?��?<:a=k�����b�΄.���M����>��2?/��@�>/t?a�%?D�?�.G?�
?��>k#	�T?�u��>Cڇ>�[P��I��8ҏ>�A?�k�>n:?*�{?��b>��=��Ț�C�Ž�	=�:�=T}*?��"?�^?���>.�>��>��>�x�:¼>6O�?�4X?��>�:�>����1I�%�N�i
H>=d%>�??��[?�?�?}=�?��`?/F��˲���=v/*=�t������Q=h?H=��=eEҽ:\;w�==��>GA>ƌ�����>�ܽ���<~�.>un�>��t>mU���53><�ľ����@>�
��5̜�=����8�>��=���>�/?=6�>a%��Ӑ=ٔ�>��>j����'?�?o�?)0�;2b���پ��K�g�>�tA?��=Iqm�ȉ��P�t�t[=�m?��^?�pY�����Y
b?L�]?���|<�������q���	lJ?n?�B2����>VT�?��o?�X�>��l�_Fm�Kۜ�@�a���p�WV�=�
�>�0"c���>�8?���>X�b>���=?<پ,u�l(���p?�h�?|�?^��?f�)>>�n���߿�,	�ᅝ��L?!��>d�f��v?Π%>y	��%툾��ľ�{�WS��f\�� ���a���g��������"�ޤ���?{Zr?�DU?��q?����_o��#c�7Ev�2&����Ǿv����K�X���?�܃���O5��{��x�������i�Q��p�?�y"?@�#�]��>_�v�s'���¾��/>�s�����zX�=�O�+�V=9>�<)�y�F�1� ����&?�ϙ>ʌ�>��A?G^�p>=���+�4�3�{��g�E>�R�>'��>_�>��V<5S�V��(�;�;���`��ƃ�>*`U?"?h5P?}��&<� n�N6 ���c���y�>[,�>��w>��l��,3���.���l���"�3���ʾ��>�,K?�>C/�����?=B?��
��e��F��J�@�u�D��>��J?P�>gy>ġ�=%���w�>��k?���>���>t���j� ��}���ܽ�,�>*%�>��?� �>�9!�9'V�)�u����:�[I�=0Ke?6Y��
`�}}�>}�Q?猝�4�휥>��E�`�!�}c�'����=:�>zg�=��O>��ž+F
���v�$ׄ�ʻ)?�?l~��!����u>v!?�'�>i�>P��?���>{�������?��W?`I?d�=??��>�~x<�Ͻ��ý��6�{g�<*->� \>��<L�==�9 �U�5�^�]=�=W�/�-ǽ8�F�wJ�Ѭ�</��<Fm>>IVۿb�I�z*ھ��������b	���{����E��z{�� �y��1��U,�
^���k�	t��D�o�8�?S3�?�:��0j��H����J���`�j%�>������z����������*����> $� mP���i��e�I('?&���
ȿ����yݾ�r?G?8vy?ť���"�:�7�e�!>�\�<�����zɚ�m�ο�ꚾ��_?��>T�v�����>O�>׷Z>h-s>cp��]��R�e<EV?�-?	�>ˈs���ɿ![��N�<���?G@ϥA?_�'��R쾒hY=h�>T\	?v*<>�3��i��*���9�>���?���?T�J=�[W�<=	��e?ڪ�;G��ѻ���=粥=�=�7��J>␒>�L� �B��4ؽwT2>��>��$��j�']��w�<�]>�ս,M���D�?W![�-\e�^Z0�dM~���>�'U?T��>%�=��+?_�F��ο�#]���]?���?B�?�*?F����~�>��۾0L?�8?Ӛ>kR%���r����=��¼j�ݻ����V�d6�=�j�>�>s�5��=���T�|(���-�=�. �?����0��*N�3@�Y]�=�e�=�,^>c�=^p���۾��ξ^��<��>?��=��>z�=i>	x6>{�J?&$~?�\�>aer>㊕=Ŝ��]	پ�.(��sԾ�R�I���i����� �L�%��h��[�-�h'�<�B��C���<�Z9�= (R��鏿2s!�xac�+G�".?��>��Ǿh9K�J'<?�˾%�������W����;b�1�'�m����?�@?�↿^�V��L�@ �| ��F:W?7����P��y��k��=����=���>�:�=�@��T3�^�Q�<-?��?
��' ����#>w�/�%��=��+?|��>,��;a��>��?}�<�<����>�R>�%�>���>��
>���=�ѽ�L,?-xV?�����^y>
�������Ph�<�h=i��w<�;L>�~J�_˙��ԃ��P����=(W?s��>��)���C`������Y==��x?]�?!.�>�zk?u�B?�Τ<�g����S���nw=��W?(i?8�>�����о~����5?2�e?�N>`h�j���.��U��#?^�n?w]?����w}����w��\o6?�up?�	T��+������徑�>^�>{U�>�/l�p�z>2�W?X�U�K濿Ivֿ-O��2�?�@��@>��=�e�<�3ۼ��6?U�=?�*-�\����­�d��=��.?)����ւ�%"���뽚L)?�8�?��>bP��s�	���>��޾�ʪ?���?�ѡ�^E�x�վv�`������'��������$�GN��{�6�З�����o_��������>�|@Td�"�>�>��.��ؿ�xy�|	���cA���?���>	Հ���Ⱦ�쌿��x���]� >�����\�>{�>|&��5S���d{�/r;������R�>����ĉ>O�D����;�!<0��>�w�>hl�>�B����=̙?�`����οa~��F]�ʛX?�?��?��?i�K<��t���w�-���#F?(s?��Y?�v��A^�v�/�"�j?�_��}U`��4�vHE��U>�"3?�B�>T�-��|=�>���>g>�#/�y�Ŀ�ٶ�A���W��?��?�o���>o��?ns+?�i�8���[����*��+��<A?�2>���L�!�H0=�KҒ�ü
?\~0?�z�h.�P�_?ޚa���p�L�-���ƽ�ۡ>v�0�wf\��R����uXe����@y����?A^�?\�?���� #�6%?��>>���y8Ǿ��<耧>)�>Q*N>wI_�.�u>����:�/h	>���?�~�?Uj?ᕏ�����JV>&�}?^��>>��?+|>�_�>t4�=7����i�y>�L=�����?ݲH?MJ�>�>�;�T)0��A��8V�k�ݳ<��>�^?�H?�&]>�8���]�<����g���]�f���[�.U̽Nֽ[;>�4>��=��:�X��|�?��	��>濗ǣ����e�?��9>E�?���þY7>�a?=�&>�@8���|
���5�E�?���?̬
?D�����;��=�gS>عW>�4>7'��վ��;>�z6?�Z���퐿坎����>�'�?�K@t�?�s����	?���Q�������0�K�9��_>�_'?G����=\?<�p>#����\���o����>)��??	�?���>�0g?6�`��� �t�>P��>S=J?R@?i� ��	����R> ?����G����
�[?�@#�@��}?v���O࿲���Mþ�����=��R=_C#> JC�⠦>�8
>vD�<������>9Ѕ>Yϑ>vL�>b�2>���=��>0ƅ�E;�d���}��i;H������̾�N��֬��q?t���\:��^�ƾ��v����<r��!A�iʆ�57=T6c>�Qd?Oml?���?��?�T�=��>����}�px¾.�ӽ-�_���B?TzY?�T?D�h>�w��Y�<�	�������4��Ő>�u�=*�?�i�>��>��T>�>@r>�!P=��^=�X�=�AJ=�e��c$:>*�>,��>>�>�B<>��>7ϴ��1��A�h��
w�̽+�?����h�J��1��:��ߦ���h�=)b.?t{>����>п[����2H?����I)�N�+���>H�0?wcW?=�>�����T��:>J���j��_>v, ��l���)�:%Q>Ql?;a>��t>3)3�e�8��O�����b�{>�6?鼷�x=�1�u��I�Ԙݾ�L>�@�>{턼���L�����~��cf�6@�=��:?�!?����#�����y������!K>�'^>�(+="�=|jK>_mj�W�ҽ
�J�x/"=lN�=��\>�2?.s`>�a{=��>ߘ���!��"f>��>?y>>???L�ռ���<�Oj�LU��Lr>z�>�[">�z�=�h4��o=k�>�9P>�<�<�Z��x=R����ɡ7>��.;"끾�¨����=b
�Df=x�]=�淽y>�Yc=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>7�3g��l���E�}��?�;��~>�bH?��ܾ��U8˽�?q��>[u�謿�˿ަ{�Ի>��?؍?r�I����X�rM�>���?Q]?I��>g˾Td���o>�X??�9?��|>��&�NV��Z?�(�?yz�?h�>M��?�]?v�>��M<��f�ϴ�2���%g>�O�>-v�>@~?��ž���+`�������q��� ��~>"3�=D��>QHK��`ݾ ]�=����wӾm���c�>hK�>�+E>3��>9�?�,�>���> �$>��=�vl�����zU?�2�?������?��Wj9"��=�����>��>?Z�!>n�1��g�>�e?K�Y?e�@?���>�h�Mߛ�b+��+��Ҩ<��F>��>	��>%3��ey>�sﾚeg�mb�>E�>S���־����,�t�0�>2&?Hѻ>&9�$�?�#?mU�>/��>I�<�E���cBL�>��>�1?�jr?/($?�ݾ�v-�����랣�"zg���>�u{?;�?���>*���F�V�<@6὘�e��sk?5A~?{2��?���?=?S '?W�O>⥺�3ϻ������f@>t�!?"��LrA���%�C:���?�a?��>����5ʽU��qg��	��Q?L�\?'?#S�Z�_�þ��<�I���N��G�;[pq�gK>Ԣ>�/���x�=��>��=Еo�h7� �;k�=�א>�r�=�D7�������*?���vg�3c�>����Wo���X>t!=�߾��?��V���r����w5��CẾ���?]��?�/�?��p��4F?�מ?�%?ԏ�>~����9þ����%=î��^���� ?��=F��F#���)��	Q����߽j
\�Rb?���>��?�?��+>o��>$�9��t��9�����7x����5!.� +��(� ܲ����68�<_uԾ�̘���>,�$�?�k-?��>q��>��>�5��(Q�>0�>�>4F�>-K�>�T>F�s=x,�=�ӽ�KR?����j�'�8�辝����2B?Opd?�0�>i����������?d��?s�?=v>~h�=,+��m?i>�>V��`p
?�M:=�G���<EU������2��0�L��>�C׽H :��M�;pf��j
?A/?m��܊̾�:׽�Ծ�B=e�[?~
?�t	��Qa�&�W���6��\p����>.=��d߾ӆ>�<B�.��M���z��s�+���A? �i?�7�P"��v��
p���H���-d=t��>��?u0?
?�G���-<��f�D_پ|�=���g>ߴY?��>�OQ?��I?MW?��I?��>���>L벾ә�>�uӽ]H>a��>��A?@�'?�=?&�?ej?)�)>�������Mƾ��>.?�'?7��>�?�-����ǎ�iٶ�i>����/�47>�-=�Z���>��2�=��>�?k�۽�B2�{4��}�g>��-?1�>ᑵ>x����f�}�=���>6�?���>���wdr��3�OW�>�B}?8xڼ�}�<-�#>���=>�_�'�"�e�=2��R*8=�ַ��Q-��e<�?=��Y=(=�;���+2�X{˻:y=�t�>+�?���>�C�>�@��� �O��>f�=�Y>+S>F>�Eپ�}���$��X�g��]y>�w�?�z�?=�f=��=��=�|��iU�����D������<�?1J#?XT?Q��?w�=?^j#?ϵ>+�fM���^�����Ǯ?k,?N��>����ʾ�樿��3��?�W?/Aa�����7)���¾ս+�>T\/��4~�����D����~���d�����?���?�.A�8�6�p��
����u����C?:>�>�Z�>��>!�)���g�Y$�E;>���>)R?�?�[?��'?ߧ
?k��>s%�.ſG朿]G�=k<,?��<?)�?E@u?B�7?8e]=�z�G6��[h)�p&�f����啽�tW�Ɉ�<��9>X��>�p�>[-�>��x�nD�o�5�z�`��>!(>_��>e�,>�"�>�a�=��ɼ/>?/��>�9�>���|i�(2ýj�=QMe?+��?� *?��g<ִ��/G�f����	?(N�?���?n�0?��Q�ܞ>�:!�Z?�����9�+>�y�>D�>�Q=&
j��I`>��>�>r����7�]k�c_.;n�?��4?ZO�<�ƿ˰q�gq�5M���/_<E���;cd���DZ�?�= Θ��9��\��\�Z�򓠾M���� ��=X���o{�o��>�q�=���=��=[{�<��ͼ�Ż<0�I=�g�<� =�Qp��|d<o�8�Y�ƻ{���h�3�$�U<�I=�O���eʾ�R}?�<I?z�+?c�C?�Uu>��>�V3�/��>����0P?��T>�JV��5��]�=���������پ܊׾��c��ޞ�u�	>܏K�>�4>���=�`<(��=�m=���=cGҺ�d=�/�=Y��=�&�=���=o�>j�>�6w?J���	����4Q�9Z罵�:?�8�>�{�=e�ƾt@?s�>>�2������xb�.?���?�T�?J�?Ati��d�>F��S㎽ q�=���8>2>���=R�2�)��>��J>v���J��=���X4�?��@��??�ዿ��Ͽ�`/>�O8>Ԛ>��R�$z1��\��^a���Z��O!?��:�Ku˾+��>�M�=��޾!Qƾ2w1=�6>�tc= \��\����=��{�Ω>=�m=X5�>�C>�j�=��#}�=�0G=8��=ApO>l���	<�@�+�jw.=t��=-;b>�&>��>�"?D?�K?1 ?d8$�����`��;S�>ge=��s>t��<�u>Ā�>OoE?[N?�L?�,�>-�=�"�>�׋>bf;�r䅿���� ��X~=<Xn?��s?�A�>�&k<LoM�a�9�6�_��<�G"?s�C?�6?�K>�3�ؿ�,U��Ҋ�خ`�5�=#�p>wI�>�k�>��M��p����F7i>���>�8�>�>�� >��K>3æ>J �>T�=&wJ;�"=�QU��0�=�-�=�9>��bTĽB�� �!>�2i>���i>˽-\��Ԓ^>~�H�'�=���><*T>��>R㸻��о,�@>��Ⱦw�1�<��=S"�R�g�i�\��G���-9�MK�
�E>B>=m��	���r?�m6>��t��g�?�?�
�>�>,=��|�Yէ�4!��R����m�>FC~>�Ͻ��H�	M���v�����>���>O#�>ʛ�>�(���I�6�f=.�Ǿ:�q��>w�V�+�$��
^��퟿�i��{�e��X޼5?�������=%s�?�I?M2�?Vf�>������Ͼ>|~�����<C&�&��wr�>?_%?��>����&�F�]ξ�+Žy�> �B���P�\P���2�e;:��ݿ�p��>����fҾ9�4�z����H��*�C�#D���r�>'�J?Hp�?�j����+�L����[�����>(Ee?3�>�w?Z?�2n�C��}����=��m?���?7��?)�>�G�=�����>^�?�;�?`�?�u?}Ͻ\��>����=��ٽ,=>��V>t�>�0>ؔ?��?oI�>>n��wE���4���Ea6�u=3�T=�J�>��>RLu>9�>��=V�O<��*>2�>���>ﴊ>2��>ㅄ>8���%*���1?G;->���>VG.?�#�>A�=�����?m��6A��2��S,��᥼`ֈ<�*�iXu=�=.?�*뿜_�?Tw6>�S����>�O��?N�+@R>���>M��1c?\>Ǚ??#�>��>^�=? b>Z)�<�ž�n.=��5��L��!T��=W��?��n> ����ɽH����ʽ:�=�ϱ��)�"���r��ԃ��B�렎=�D�?��
�qَ�O�A�~�	��c"?CX�>�}9?f,w�(��-�)<�?���>�濾�蒿nk���¾��}?��@�=c>�>��W?�?�1�{3��pZ�6�u�y&A��e�i�`��������a�
�o鿽I�_?o�x?�zA?F<u2z>1��? �%�o͏��$�>q/�o';���;=�'�>�$����`�=�Ӿ�þ95��;F>�o?*%�?-Y?�CV�ު�;�;x>��?��=?N��?�<?UD?d+�=*�?�u��v��>Mk�>A�=?��Q?�`"?T�>[!>���<�<�uX���r���K��2�D%�<�˯���:�Pe@��]�<�L;e
a=���<�D��o�=d�=�!=\^�=D�_>�J�>)��>Ny^?�M�>�A�>��5?����K�B�=�Ӿ��&?5J@>����~��7��߾��	>��c?��?��<?���=�"?���6���?>k�r>�`�=_<>�b�>��s�i��h=A|�=��>m��=��!�3�M�F��w���MM�;D0�=���>R3|>�1����'>i�����x�`�e>O�ֺ�>"T��`G�-�1��/w���>�K?�~?��=�w��[��L�e���(?�<?�BM?�w?*�=�,۾��9�ΆJ��X���>�A�<I�����-#��!l:�wD�:�gr>�E���Qhc>l�d�ݾ^n���I�cy�ED=}����[=�k�$�վ�t}�g��=X�	>A���v �z=��-�����I?h=`?����S�y���R�>��>��>��D�&�t�L@��Ѭ��w�={'�>G�<>B ���r��F��v���>qyT?�
y?9�?�Kw���k�f�S� �v~��^���3��>E4�>ԝ?>
x=Iy>��]�m�9�"�o�НK��L�>�x�>Ϯ&�R	I��-���MT���ƾ��L=h?(��>a�	?��'?�:?�q?�'?��?���>b��Y�ؾt)2?ޕ�?y! =��K�
��pȾ�?:���>��?������>R��>;�:?H?�\?b�?J8>���_�\3�>p$>b�������G�>���?�޴>�g]?`�y?f�>i+�8�޾�~�<���>獑�Qg?pZ?�@?ƶ�>-u�>_����T>��>�[�?�Qw?X�W?K�=S�>�6>Uk ? �=_�C>uS?tB?Z0Y?�O?��D?�?��=i2{�����V2�=��=^ѽm{�� X=�@1��棾�Ͼn�<<7�=�^½�?g���� i��e<��9ua�>=�s>7��U1>��ľ=S��_�@>�1��+P���⊾��:����=G��>��?���>V#�:��=럼>�6�>���44(?��?~?B);x�b�"�ھ:�K�d�>(�A?���=��l�	���w�u�Eh=�m?�^?��W������_?��j?ʆϾ��=�)Gƾ]������?f`$?6s۽��3>?�^l?�7?QP����v�����fr�������=�r�>!����F�RՅ>J0<?hA�>|�D>@"�3���R�F�@�¾V�>�ے?}ʮ?*\�?��x>ǥz���ٿ��Ѿ죥�Yv?U��>�v���_"?ʂ�=���Lm���:����u=Y�QM���-^�.�`�\S�ȑ��*샽�t�=�(?��w?b�Z?�n?Z����c�\�n������U=��d�,�Ird�/fJ��7��i��d���E��5���*;�fx�T�H��?��&?�f,�X��>Kf��~��m�Ⱦ� I>σ��_��+�=�n~�|=�;`=0h�]9&�\"��Q-!?�"�>+�>�d@?�]��*>�Q2�As7�7G��=6>\�>j��>!��>� ;{�5�� ��˾�'��N�޽x��>�5c?��3?O�j?Wpb��X(�a���+�:�漰�3�E��=���9��>Tߕ="����0��j(�G����9V��f�������=��/?&ܢ>;�B>+�x?I]?Gi�,��9����CD�<c��=ţu?��?d��=PQ��@�񾬺�>Y�l?"��>�	�>|����[!���{�(�ʽ/�>��>��>f�o>9�,��\�#k��Ƅ���9�	O�=�h?뀄���`��܅>�R?Nz�:�OH<<~�>0�v���!�?���'���>�z?���=��;>�xž` ��{�><���I6?�p,?-���w�)��� ?M}?���>���>	�u?gs�>�c��R����0?�HT?�#C?I�>?�5�>�ʂ=#^S��%�vQ���8">?_t>�G�>�@:Iϕ>���Osl��^l=�֖�R�>7oc��C=���=�ܥ=�ʽ	l>��>"fۿ:K��xپ����7
��숾���?_��ޙ�k�������x�����t'��HV� Gc�����Նl��}�?�-�?�}��$��!����������W̽>��q��`�oҫ�:��D��e��N����k!���O��i�l�e�L�'?�����ǿ𰡿�:ܾ+! ?�A ?:�y?��9�"���8�� >GD�<y-����뾱����ο6�����^?���>���/��O��>ӥ�>!�X>�Hq>����螾�/�<��?;�-?#��>Ɏr�/�ɿa���z¤<���?0�@�}A?)�(����`XV=O��>�	?%�?>wr1��=�߰��1�>�0�?���?��N=νW�sw
��ze?�I�; 
G�޻��=�7�=�=����|J>�T�>|M��A��ܽ2�4>�ȅ>"	"����d:^���<�c]>�.ս�I��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=p6�����{���&V�~��=Z��>c�>��,������O��I��V��=����@����� �f�%��w�=�m=5�>~��j��=�<y���4��P$�&�^=���=��O>�?0>�T.>҆q>�I?��b?#��>��%>�Q�� �������w�����s����K��ǩ+�@��tﾘ�������r�'���;��!=�#�=�6R�c���?� �a�b�[�F���.? w$>?�ʾ��M�n�-<~pʾ7����܄��᥽�-̾�1�'"n�f͟?��A?������V�]��cX�����[�W?qP�ʻ�aꬾȣ�=����b�=%�>~��=���� 3��~S���/?��$?v���^��V��>����=�
*?��?
e==���>-??��<��+̽ǈ>�eu>Ԛ>���>��>����}	���)?�R?A|E����T«>?C���>���r�<m�K>W�ڽb�ý��p>��=��|�3���Q����g=3(W?���>m�)���e`��`��>Z==_�x?��?%.�>V{k?��B?�ߤ<�g���S���ew=��W?�)i?͹>㉁�1	оށ��s�5?�e?��N>�bh������.�?U��$?#�n?F_?vt���v}�B������n6?�9�?�1��	���ƾ������=�3?��?QP��XO,>/h?�$e�_���ϿM>G��+�?k�	@�@��>��m;����?�q1?1��
W���c��{쾊��=��M?_�Ⱦ�y�#B�ҏ����"?�b�?�P�>7��Y���o>�2���ݭ?�L�?ڱ���	���������:Aʾ��0=�2��_"&�^&�"_ž�|1���㾲P$��׎���<?s>Z1@�|i�ǋ�>K[ ���ڿ���=��yL ��<��-i�>�Y�>����Ǿ�\������TS��6V��Wl�/_�>M#>r��˿����{�za;��ܠ�*��>}��ֈ>v�S����Xe��$�5<��>?��>���>j��������?n`��5Hο�������X?e�?,`�?�w?'�=<��v���{��B�=<G?�vs?;Z?K�"�\]���8�%�j?�_��zU`��4�yHE��U>�"3?�B�>\�-�"�|=�>���>g>�#/�x�Ŀ�ٶ�&���\��?��?�o���>p��?ws+?�i�8���[����*���+��<A?�2>���M�!�A0=�RҒ�Ƽ
?X~0?{�h.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>`ք?�;> _?���=ṾCXJ�Zr*>w�=�m཯��>�II?�(�>��=��2*�=:J�U���	��?�Y�>qe?31I?.�Z>��ý4�p��! ��f���C���"��k�ݝl�� ���!>8I>���=Gp5������.?����Y�п9���aW���z?�8�>\l6?�98��h�_m8>׍y?n��>�&��ᶿY)����)����? ��?��?�r���랽�L�=m/�=]�C>�,�>�����龩�=�jP?4h/=[r��
���$�P>4��?. @4˥?�|��5?���te��1ɀ�d.�\Ke��Ś>fcE?��*�ޥ>�!??�>��j������{��J�>���?�0�?s�>j?HZ]���8�@�>g�l>gU?y�?��_�価;t>X?���o���S��Y^?'$@�@N@u?�S����ӿP᛿����<߾Y��=�"Z<��L>�o�;8�>�rĻ� >5��=��2>�z�>���>�ٜ>��#>��I>��>A �����Ǳ��r���^]�k������&ɽsЏ�6;�Yt�?!���]��S6�Xԛ�O���c�>���vP��%>� W?x�S?��?(U�>�~ �|Hb��ľ � �R\��>^�=ҩS>�l8?"�'?�;?p-p=Εξ�p��0���!���nM���>�[>.��>;�>gn>�j�V�J>��\$6>���>� F�e�w�H��;�h�>�R>j��>� ?�C<>��>Fϴ��1��k�h��
w�r̽1�?����S�J��1���9��Ӧ���h�=Hb.?|>���?пf����2H?&���z)���+���>}�0?�cW? �>!��s�T�4:>:����j�5`>�+ �~l���)��%Q>wl?�g>_�u>dD3���7���P�KI����z>ޡ5?񁶾�x7���u�-�H��Oܾ�O>���>��]�>�H��ȏ�4i�
{=�D:?f�?ӵ�����u�K[��R+O><\>�� =�S�=��M>�Hi�pI½xH���)=���=K^>?�k,>��=���>铙��O�չ�>oKC>J�+>E#@?�%?���<���|�����-�Rx>�+�>R�>�>�K��Q�=�D�>��`>K��ƀ�����?�X�X>|�~�_�]�y=n�̲�=հ��h��=|C�=u��u=��x$=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>�$ �p�������Lv�tq��Ց>WI\?p����>���Ľ4�?E�?����Ѧ�ֲӿ�M|�}��>�a�?%(�?�AK�%ʞ��3_�7�> ��?{�q?��>�a"�k�ʾ9�>�&S?z&`?��>ږ!�R\���?%�?��?\m�>��?�0l?/�>$���*F�\:���8��U�>%�W�W���>M$^�����)��Zk��hS}�:�'�؅2>��=��>��e����՗`��b�Dy��d�=
��>�\�>��=Ə>��?s�?��H>�9L=��=�ؾAPȾL?�Ɋ?�D���?��j2�څ=�½����>.�1?��=�?�;�`>�\?��?2<5?t��=F8Ҿ�ݥ���ɿ����L_ټ/�,>D�?�3�>�V��e>���X�ž�>ꝲ>��Ƚ9���������;>�w>��?���>��j�\4 ?��#?��q>摱>��C��㑿��G�֏�>�>�>t�?�y?P�?^����2�E+��=U���P]���G>l�w?��?2E�>���Zx�������2m��Ҳ���? tk?����
?4X�?�A?�:A?�Y>���<վ�=|>��!?�R�׸A�oL&�\��-	?��?���>�g����ֽ�ͼ!$�;����0?T�[?/7&?���`�`�j�þ:X�<����r����;�� �>u�>2������=T:>���=�6n�6��#u<�=��>�M�=�x4�Gu����4?�A`�,+|�1��>�����>���=����{?A񽫡]�j���=Ŧ�5�uۋ?���?�#�?RzP�a�}�M.?�`�?r�?��
?E���o��l��������~#�<5��3�<#�>l�P=a6���Ơ�f���wh����#��k9���>r��>���>�u�>�m >X�>�8�40������PǾ�8���Z�"�6�G)��Ծ�dk��P���x>�վ���h^�>ݧ&�`�>ǝ"?�{>�P">�j?y�H�lR�>�/�>�>���>K�>;{3>��g=�A��5'� LR?������'��辎����3B?[od?�0�>i�|���u���}?چ�?s�?�@v>V}h�a++��l?�8�>����p
?�Y:=D����<�T����-��.�=��>RI׽�:��M�Oqf�j
?^/?�)����̾�+׽(�����?=���?�+?�>��L�ͱi�h�_��A��7�e=���흾�R8���b��2��=7��#�|��$ ��ؙ=��/?`ƃ?dg�\��4�վiy���G�o��>���>m�>u��>`>FV��>E�ϖW�4�7�K������> Qt?]z�>�tL?_"8?R;>?Z�e?��> Q�>�g�I�>�.=��>���>$�?��&?<2??�'?"W?�K>�;��&	����8#?B�?6B�>g��>�?{X#�r��-���ւ=��5��,���)>
��=LϨ�����{�L=IG\>aY?C��Ϭ8�;���;	k>N�7?�}�>e��>���D,��r�<	
�>6�
?�H�>����5|r�>a��U�>Q��?C��=��)>���=�D��j@Һ3]�=�����=���N�;��E<j~�=���=`t�[b��C��:\G�;���<t�>�?ѓ�>�C�> @��� �׵�i�=�Y>uS>>�Gپ�}���$��V�g��^y>�w�?�z�?��f=~�=)��=�|��.V�����K������<��?�J#?�WT?h��? �=?�j#?h�>A*��L���^��Q��n�?#!,?\��>�����ʾ憎�3�<�?�Z?D:a�����8)��¾��Խ1�>4T/�<,~�����D�|���(���u����?C��?��@��6�0y��Y����C?V�>�^�>��>��)���g���C!;>Ї�>R?��>.�R?!7f?"LO?�<�=T)��^���s��2]=$n>y?�X?l%�?�n�?7��>��[<{����x)��n8�s��g�t>]� >+z�>Hw�>���>X�~��۽�K^<g�m����=�>H�?��>%��>io�>�Ӳ���G?��>(���]��mQ��U�����>�X}u?���?YF+?�z=֟��lE�`����`�>_�?��?�*?S�T�Fc�=vvռ�򶾫�r�׸>��>��>���=�H=�w>[��>��>�����i8�5FN�n�?EF?]��=�W����G� �@Ŝ�)c�=Y%�(���D�X� �J�6>@���7��x���<����澬���l�־1h�����N�?X�>��\>�nq>Aq(�����J��� ���y��M��!@���
=�F7�н�k���n�)>�=Պ�=(	�� #˾ۖ}?7pI?Q�+?ΜC?rx>ܘ>��2�GK�>�݆��?�V>8TN�����Kp:�z}��������ؾ��׾��c�݃��k�>&I��>� 3>WI�=�<���=�t=Wz�=� -���=q%�=���=��=��=�	>@F>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>s��=v�2�T��>��J>���K��D����4�?��@��??�ዿТϿ6a/>=h8>�>=�R���1�xn[��]`��Z��!?�;�Z̾E��>#��=M>޾��žhp0=-7>Aze=�k��j\�;v�=��y��::=YVh=���>
�D>�x�=�쮽t��=y�N=��=x�N>�薻+�4���-��@2=|A�=�c>�&>[��>��?>T0?vPd?�4�>��m�/%Ͼ�5���B�>��=;M�>Z��={�B>��>��7?i�D?��K?�W�> �=���>���>֜,���m�+�����Z̬<��?Ɇ?J��>-S<o�A�a��.Z>�HYŽ�q?0T1?ns?:�>	8�u̿��}�;�w�7�ǽ�Y2>�^�>���>�W>A��=�4��uu�j,�=��>Ao�>�ְ>ݜ>a#3>m5v=�͖>�Z3>�,>��=�>� �=�d�f�Q=w�����=�0��XI���I��[��1��T���y��	���Aֺݰ�=�a�>�mA>y�>y�.;�} ��(\>�Ak�B[X�s)>#b���U����F�����5��#p����>�>��=����w��>G�]>��@�\��?E.�?��=��=N��8|����ͽ�����:r>ኚ>�f��M��h:g��=\�0r����>���>Z�>X�l>9,�|#?�`�w=L�b5���>:{��2���#�+8q��>��,����i�ʹԺ��D?VF��-��=�!~?¯I?��?��>d���ؾ7=0>�M����=)�l*q��y����?�'?ѓ�>C�q�D��J̾����߷>5I�=�O������0��8�~˷���>�����оj&3�xf������B�gOr���>��O?�?4b�X���RO����NF���m?,�g?��>LH?�C?����j�kp��(`�=2�n?���?`;�?�>���=�Չ���>2?�˗?�^�?��r?�;*�@�>~�<
�&>-Ҳ��E�=�j
>���=�?>�E	?�?��?�����
���ᾜ��J�^��=��=c֏>e+�>�R`>V��==���=%j>��>�;�>�X>�>��>�r���$��C3?s`=A�>Ư2?�/�>��~<���ƼP=�w�e9>�=��Qm��]~<(=>�A�J�> >?-�:�?1\k>ސ�3v?:�~/F���N>��2>+���h�:?�5>0��>"�?H>R)O=-Rt>E�̺�Ͼ��=����y{�p�C��RZ�,�<�|>�虾���^���)^�������w�}���z���+����=��?b½Tq��Y|9�{�o�g�>ˁ�>��e?�=��Ȅ
��>JZ�>H�?i,�Dڗ�i���	���9:�?��?;c>��>B�W?�?��1�3��uZ�C�u�\(A�e�T�`�|፿�����
� ����_?��x?yA?�T�<�:z>A��?��%��ҏ�o)�>�/�%';�5B<=I+�>*����`�L�Ӿ[�þ�7�DIF>J�o?'%�?NY?�SV��㙼��%>k�<?mV2?T�~?xT5?�@:?/�ýU# ?�> ?Q_?A�)?=F0?��?�fl>&��=���< r�=I=���:��q���O��=����<ȸ.=����	;b s;��F�$����<'Q<�*�넘;��=���=婽=G��>ȍ]?� �>9G�>��7?�W��7�0����.?�r>=o(��"�	p��1��>C�j?Aǫ?�Z?.�d>WB�tC���>�߉>��&>��\>���>{��)QD�{U�=�>�2>֙�=%~J�@π�[�	������Q�<x*>�L�>��>Z�u��79>�7��8h��vrS>��F��ߺ�� h��D���1�|'e����>��M?�?�ct=7NﾬѸ��d�k�'?�*>?��K?)n�?��=�ݾw7�A�F�}�6����>�=�U
��餿m���5������l>Y��G栾'Kb>����x޾�n��J�X�羈-M=~���U=d�� ־�4�u��=
>I���$� �����֪��-J?��j=Yy��dU�`r����>��>�خ>�C:�Gw�<�@�y���1'�=��>��:>U����z}G�(2�S��>�3E?._?4G�?��~���q�/�?����������ɼ=0?3��>�q	?��J>�ȵ=����W����d��F�W��>�!�>0#�~E�)�������y&�@�>�^?��#>_@?��Q?�??&�_?�(???�S�>B����ж��A&?6��?��=��Խ�T�� 9�HF����>{�)?�B�۹�>Q�?�?�&?�Q?�?w�>� ��C@����>�Y�>��W��b��A�_>��J?ؚ�>q=Y?�ԃ?w�=>\�5��颾֩��U�=�>��2?6#?O�?�>0l�>瞡����=)�>yc?�5�?��o?���=��?��0>
f�>���=�B�>�C�>"�?�OO?��s?4�J?�>��<v���鶽m�q��XV���|;��F<��w=D��X�u����Wl�<���;S۵��}�Mf�1�D��d��m��;m]�>��s>1	��|�0>��ľ>K��.�@>jx��	P��ߊ���:�Rҷ=.��>*�?꩕>{T#����=C��>�C�>����6(?,�?q?�!;Ϡb���ھ��K��>�B?��=��l�E�����u�V h=��m?�^?��W��#��O�b?��]?@h��=��þz�b����g�O?=�
?3�G���>��~?f�q?U��>�e�+:n�*��Db���j�&Ѷ=\r�>LX�S�d��?�>o�7?�N�>/�b>'%�=iu۾�w��q��h?��?�?���?+*>��n�Z4���������'\?���>]���B$?�	�:��о���P�����+���A4��B����M��D�*큾5��Q�==?2Dq?�bp?F�g?���Ϣf��f]��K���Q�E������=���?�ӂ?��/m�H��L|��K����$v=>��$3�<��?i~?�X�R��>a�p�4���i����^=:žRC�=�<���ϫ=��=��e���^����?���>�p�>C�b?��e�d#Q��2�f<7�%�߾�"�>4�>>��>N%�;��a���\�No�߅��$�;�\8(>+Rh?B,L?�1�?/x=�b�ꮊ����h=(b��[�>��|>��>�����M�"�E��E�K�n��6׾�B����sC�=t�?��>!p�>MD�?��?l���J�&�v��Z�f<���>|�?���>s��=9�=�9���>�8n?���>z�>�^��p�#�c$}��*ݽ��>-M�>�r ?��x>�)��~[�np��P����q8����=�[g?�8���e�K]�>i[P?�A\;U$�;�՜>h>X��������-�@��=�?�n�=0�:>�Lƾǻ��y�E���i�(?@�?脒���*��'>�t"?V��>�>���?�Ι>u/ľ;�,��?�F^?d�I?FFA?3�>�=����N�Ƚ*�%�z\/=9g�>u�X>	'i=g��=).��jY����Z�==�ѹ=I�Լ1����l<+԰�[$B<LM�<�"5>� 迵;H�|����
�����z�����B���r���'�)�žg���<E�����"Nk�m�x�xx���1��3���[�?~$�?燫�����-%���er����3�>$5�F�"������t������aO׾����aJ��C`�b�O�O�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >{C�<-����뾭����ο@�����^?���>��/��n��>ܥ�>�X>�Hq>����螾d1�<��?7�-?��>Ŏr�1�ɿb����¤<���?0�@�yA?��(��쾓�U=��> �	?s�?>�H1��O�+���Q�>g7�?]��?#JM=��W��	�a|e?��<o�F���߻�&�=*'�=h�=���J>,]�>����.A���ܽ\�4>�څ>�"�.����^��J�<2~]>^�սpQ��"��?��a��m�� �y���#w�=
�I?<^?�U½�d? �q�u�Ϳ����ܚc?�m�?�)�?��G?����^!�>fH۾�76?݋[?"�>9���q���=��t>¤��<U��^J�A�<A�>�f�>������A��S+U<t������ƿ��$�6|��u=#�ٺͭ[�g������wU�q,���lo�l�轜�h=ϕ�=ÇQ>|f�>W>�Z>�dW?�k?CK�>j�>�a佁����ξ�z�t?�����K�������棾HP�"�߾E�	�������3�ɾ_,=����=X.R����A� �L�b�~�F���.?�w$>�ʾd�M�.�,<�cʾ乪��i�������1̾A�1�e%n��̟?��A?8��� W�� �])�㘹�ĮW?�����ା�g�=.U���=r�>��=h���3��lS��i0?S?�y���o��.@*>�� �e0=(�+?�?93T<��>E:%?�+�(S��Z[>2�3>�֣>��>�	>R��V5۽z�?'�T?�4���Ȑ>mp��M�z��a=�	>.5�t=�'�[>L��<쌾n5W�n���l{�<�(W?Q��>��)��da�����Y==��x?��?.�>b{k?��B?\դ<%h��t�S���bw=��W?*i?a�>����	о����P�5?�e?��N>	ch����L�.�MU��$?�n?_?̀��&w}�}��z���n6?�{?T!k�&몿-�'��䪾 ?���>h��>�>�0I�>�c?~hx��@���g����9��#�?~9@`O�?{͎=,�=\u8����>��>��c�7����|ս!Ծ'S\=V:?B�2��(�/���N�g�N?�W�?���>'������E�=�Oq����?�L�?$��9�»g�U;g�Evݾ!k{�h��<��U�2p�����3�I���x������0M�vD}>�@�ƽ�?��o�'��_�ȿq�������ΰ��(?Y��>�-׽�ء��kl�r����.G�f?H��MY��M�>��>5���������{�0q;�����>N�	�>	�S��&��Κ��2�5<W�>���>M��>]*���轾�ę?c���?ο[������c�X?3h�?�n�?tq?�f9<c�v��{����-G?c�s?'Z?op%�E>]��7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�^�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*�+�+��<A?�2>���I�!�C0=�UҒ�ü
?W~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�3N�����Xe����@y����?N^�?i�?ӵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Pj?���� ����U>	�}?n�>��?���=M��>���=��Z"/� A#> 7�=�>�Ѡ?بM?FX�>��=$�8�D%/��\F��HR�!���C���>��a?|vL?	Fb>K��jV2�_� �xͽOv1�]1�W@���+���޽�\5>>�=>��>*�D���Ҿ�?k���%ٿ�������k8?D�l>i?�s߾&4���-�=$QY?�j�>��f���5����� �?���?�?�b�U½���=�;�>��>�ni<`Z�V{Ҿl�>t�0?�L)�eY��'d\�Y�a>�n�?vK@凴?�z�k�?��p��Y��9]�7����>h�2?�k��|�$>+�?��=��c�����Q]y�O2�>cݰ?t�?c�>�Kb?o�l�g�6�q2=�<�>��f?�
?~B񽎅
��g>���>^�&�(m�����_V?7@G�@֏W?�§��=Կ����������-�>-��=?U[>B�����=w��������=];N>!ҧ>��{>`>^>&(?>_8G>9�	>l҄��+*��Ϡ�7���f,=��"�i��w�Z���l��n�r������l��|񽚑Ͻ$�a��,�g�d�EJ=9�L?Kj_?lv?6�(?�w߽fTW>|�Ⱦ��=���1�x=~y�>�XY?Ȳz?WVD?eā�o�Ѿ0�Q�G�f�����SK`����>j�=�@�>���>���>n��<�c�>T>>kX�=�4=>� �=�ء��>ۼr>�>��>l�a>�C<>��>Fϴ��1��j�h��
w�m̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?%���z)��+���>}�0?�cW?�>���T�1:>9����j�5`>�+ �}l���)��%Q>wl?g�?>�W>��$��:���9���}����>��)?%���Y���{���K�J�-�(>��>Z=�s�te���~�ŷc�-Ñ=p�8?(^?"��Խ�MZ������_x>k�^>�!;7ſ=��?>}6��r����@��$k;噤<�Y�>�N?V�+>�Ԏ=��>kB��	�O����>�B>~�+>��??�%?�?��䗽-���)�-��w>zE�>$�>@�>=tJ��*�=}S�>��a>O��/y��)��}�?�$�W>N�|_�W�t��lx=8`�����=^�=� �0=��w%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>?N��^���щ�p*��� u=��>�TW?j����?���ל�\�?>�?{� ��y���#��Q:{��_�>T[�?>��?~eh�����=A��i�>:��?vi?���>�� �Q/��X~�>sK?00?)��>(e�m��MX(?�D�?�v�?ń>��?�)Y?0�?�0P�=�T�ok�����e~8>s?�$?��>:���6Z�}n��ǽ����H�&iE�X��>��6<'�>�O��ֵ?�	�<>b2h������v�לe>�ω>�W>�j�>v��>AZ�>J�>�-W�]����D�;-���K?���?)���2n�CO�<W��=�^��&?�I4?*k[�{�Ͼ�ը>�\?l?�[?d�>=��O>��F迿5~��s��<��K>)4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��)S��GB�>�e!?���>�Ү=�� ?��#?�j>2)�>aE��9��P�E����>��>I?��~?��?�Թ�}Z3�����桿��[�|9N>q�x?�U?�ʕ>)��������jE��GI�����!��?Ttg?�P�]?82�?��??"�A?w(f>���ؾ�����>O ?P��&�@�� '��K
���	?�?\��>#ɒ������v�C����d?��Z?�(&?@�+�_�EIƾ=(�<�� �����:<����{>�>�𐽰K�=��>�z�=�lm���9��d�<��=��>s��=ӧ:�����h.? ��y��I�=S0n�j�>��v�>n�>	$����^?[׀�����ɫ���k��9ҍ?t��?�r�?R�ͽf�Ew2?!��?��?�\
?����[?ﾠu�Ad��'-l����u�>Ӈ�>�|�����\����������r��Q)�>WC�>r9�>�	?��>�>U�j��1�UE��� ���]����O6�(�#�eg ���*���^:���;�+��Nj>���B�>Ym?{A�>�/>Ì?s����>:�5>Y�>�c�>�wB>~�3>��=��)��Ľ�KR?�����'��������3B?�qd?E1�>xi�>������0�?y��?s�?�<v>�~h��,+�_n?�=�>u��[q
?FR:=�H�=�<�U�����4��H
�5��>�F׽� :��M�nf�Jj
?�/?���ċ̾�;׽����,�=��?ø(?�(��|Q��l�r�W�PI�?L���d�Yt���#�~ l�M̎�E���9��p�*�]=(?���?�� ��d⾟ڮ��k�>�?���V>��>�Χ>rX�>�l>d���1�A,^��Z*�|���D�>}{?hό>�lI?(;<?�P?��L?t�>��>ƪ��Y��>*�;��>���>\�9?�C.?n0?4�?v�*?��a>���������ؾ=�?��?�n?e�??t?b5�������o����g�A�w�"䁽e=�=�@�<C�Խ�tq��)X=Z;R>oX?���`�8�D����k>��7?���>s��>����.����<�>_�
?CF�>  �V}r��b�hV�>���?� ���=��)>Q��=�����*Ӻ�X�=.���z�=�@��ɂ;��\<6�=Y��=�'t��s~�V�:Fk�;z�<�s�>_�? ��>nD�>�@��?� �	���a�=Y>vS>�>2Eپ�}��Y$��L�g�@\y>w�?z�?'�f=j�=b��=}|��zS������������<�?J#?�XT?���?Q�=?�i#?�>8+�wM��}^��0���?k!,?n��>P��E�ʾ�񨿜�3�ܝ?�[?�<a�n��<)���¾  ս��>�Z/�z.~�M���D���������}��(��?ӿ�?A��6�iy辸���X\����C?�"�>bY�>O�>t�)���g��%��/;>ʉ�>�R?	��>e�P?Y�z?�-]?G_Z>��<�f����{������i&>Bu??�K�?��?Hx?�g�>�n>�c2�
�㾵���
�)�s �C�~�^^^=P�^>х�>���>1x�>���=&��~���m_D����=9/p>���>Or�>���>0�{>�@�<��G?���>�\������줾cŃ���<�Ȟu?��?��+?�-=�����E��C��/M�>.o�?J��?�4*?5�S����=�ּoܶ���q�o*�>sܹ>P.�>~��=gF=�`>��>Ġ�><�>b��r8�kM�/�?	F?���=��ſxRq�<,p�����Q�z<2���v'c��ѓ��nZ����=�s���/��?��GW\�-h�������W��;Q����}�J�>ro�=�_�=hc�=t��<��μ�y�<�D=&�<�=2�u�vQl<8�;�|���	���M/�:S<bjA=^̻|�˾�y}?�7I?e�+?��C?��y>J�>B%3����>����0?y#V>�Q��l���*;������"��J�ؾ��׾jd�YƟ�S6>&�I�ͯ>�m3>l)�=s��<8��=��r=�^�=�O��='��=Ɂ�=��=���=Ѽ>�:>	8�?�r��Ң�;=X���M�)�@?u�>Z��<����O�5?�=[���l��,B�ҽr?E�?4��?j�?l�����>Ӗ�����>Z>��$�$�m=�=Š;����>�+�=e������6��i'�?�� @��'?.܄�����{�>��#>Ѽ�=�I���6�V�/�d,!�7�(��@?7���꾗u^>!�D=�L�aʾ^=Y/F>⚆=�
�9c�h�\=��'�t�-=��~=]�t>��9>]��=<�P&'>M�;��w=@=>x,�`�������r=�<�=��=>V4>3��>?�?�a0?(Xd?�6�>�n��Ͼ'?���H�>��=�E�>P��=|rB>ʏ�>6�7?o�D?�K?�>���=	�>��>D�,� �m�m�9̧��<���?�Ά?xѸ>��Q<��A�����g>�C/Ž�v?(S1?�k?k�>�U����9Y&���.�"����b4��+=�mr��QU�a���Im�4�㽯�=�p�>���>��>9Ty>�9>��N>��>��>�6�<}p�=Aጻ���<� �����=�����<�vż×���u&�8�+�/�����;g��;.�]<{��;R$
>��>3�4>>��=s�t�U?>FH�0p�-�=s���H��TO���m�t��S�ֽ�gK>Idi>��-��=��[��>��N>���;i��?�,~?��@>�����找���=��k�2�>��<H��~�=�d�[�gZ����[��>Yߎ>$�>��l>�,�L#?��w=��Yb5�~�>�|�����*)��9q�#@������ni��kҺ�D?�F��f��=i"~?��I?^�?ݍ�> ��φؾM;0>�H����=g�*q��h����?'?���>�쾤�D�W̾~��kз>z\I���O������0�J���������>�T�о~3�^f������ƌB�
jr�c�>r�O?��?B4b�G_���WO����+ꅽ2t?$�g?�>tD?�I?�ۡ��f�$|��!T�=��n?Ӭ�?�@�? c>�n�=qO����>a?��?���?��s?h�=���>�C:�:>�v����=X�
>�p�=q��=w?B9
?U�	?��P	�i���T7^�g^�<(�=��>���>��o>���=�{e=s�=��[>3��>�&�>,�d>y�>5.�>���1��n&?���=!��>��2?�C�>��X=:!����<�e]�tB��.�[���(�߽��<�MH���N=����>C�ƿ��?b�Y>����?Gv����?���V>�T>~���W�>NKD>�w}>Xӭ>|�>�>�N�>{*>��(� >-��'#+��4���C�I����=-�����"��2���;���@��Jv�b�(��d::��5=��?�K�������=C��ʭ���?�|�>K�i?>����͜>���>b=�>|d��돿Knl��	޾���?�@�3c>6�>g�W?S�?O�1�3�oZ� �u��&A��e�+�`�+፿l��� �
�`����_??�x?�vA?ל�<�/z>.��?m�%��Ώ��#�>�/��#;�'<=�6�>b.��m�`�b�Ӿ�þ�2��HF>�o?#�?HT?IV������>�'H?33?�	�?i?,?Rp?1�H�a6'?�7>G}?�F(?g�/??n;?�w+?�S�<Z�E��$��d�Ͻ%����]�^ �w�����	f=J� >����O�[�=����~�0>�}=0�,�s�>���=�?�;,ĸ����>Ay]?k4�>�6�>F�7?t��?8�����[!/?�D4=�����M�������%�>��j?��?�?Z?�c> �A��B��[>�Ê>"�%>$�[>��>�����D�b�=x�>V>@|�=�xL�L���L�	�\����p�<1�>-�?�2;>��i�il>���M�u���]>��R���	�qO��\?��ʗ�s��>�pP?�K%?ɱ >����̽��b��(?�H?�51?.\�?��>�4�[�C���E�R�)����>���=�	���Z���k��eC�\���#>㲰�G栾'Kb>����x޾�n��J�X�羈-M=~���U=d�� ־�4�u��=
>I���$� �����֪��-J?��j=Yy��dU�`r����>��>�خ>�C:�Gw�<�@�y���1'�=��>��:>U����z}G�(2�S��>�3E?._?4G�?��~���q�/�?����������ɼ=0?3��>�q	?��J>�ȵ=����W����d��F�W��>�!�>0#�~E�)�������y&�@�>�^?��#>_@?��Q?�??&�_?�(???�S�>B����ж��A&?6��?��=��Խ�T�� 9�HF����>{�)?�B�۹�>Q�?�?�&?�Q?�?w�>� ��C@����>�Y�>��W��b��A�_>��J?ؚ�>q=Y?�ԃ?w�=>\�5��颾֩��U�=�>��2?6#?O�?�>0l�>瞡����=)�>yc?�5�?��o?���=��?��0>
f�>���=�B�>�C�>"�?�OO?��s?4�J?�>��<v���鶽m�q��XV���|;��F<��w=D��X�u����Wl�<���;S۵��}�Mf�1�D��d��m��;m]�>��s>1	��|�0>��ľ>K��.�@>jx��	P��ߊ���:�Rҷ=.��>*�?꩕>{T#����=C��>�C�>����6(?,�?q?�!;Ϡb���ھ��K��>�B?��=��l�E�����u�V h=��m?�^?��W��#��O�b?��]?@h��=��þz�b����g�O?=�
?3�G���>��~?f�q?U��>�e�+:n�*��Db���j�&Ѷ=\r�>LX�S�d��?�>o�7?�N�>/�b>'%�=iu۾�w��q��h?��?�?���?+*>��n�Z4���������'\?���>]���B$?�	�:��о���P�����+���A4��B����M��D�*큾5��Q�==?2Dq?�bp?F�g?���Ϣf��f]��K���Q�E������=���?�ӂ?��/m�H��L|��K����$v=>��$3�<��?i~?�X�R��>a�p�4���i����^=:žRC�=�<���ϫ=��=��e���^����?���>�p�>C�b?��e�d#Q��2�f<7�%�߾�"�>4�>>��>N%�;��a���\�No�߅��$�;�\8(>+Rh?B,L?�1�?/x=�b�ꮊ����h=(b��[�>��|>��>�����M�"�E��E�K�n��6׾�B����sC�=t�?��>!p�>MD�?��?l���J�&�v��Z�f<���>|�?���>s��=9�=�9���>�8n?���>z�>�^��p�#�c$}��*ݽ��>-M�>�r ?��x>�)��~[�np��P����q8����=�[g?�8���e�K]�>i[P?�A\;U$�;�՜>h>X��������-�@��=�?�n�=0�:>�Lƾǻ��y�E���i�(?@�?脒���*��'>�t"?V��>�>���?�Ι>u/ľ;�,��?�F^?d�I?FFA?3�>�=����N�Ƚ*�%�z\/=9g�>u�X>	'i=g��=).��jY����Z�==�ѹ=I�Լ1����l<+԰�[$B<LM�<�"5>� 迵;H�|����
�����z�����B���r���'�)�žg���<E�����"Nk�m�x�xx���1��3���[�?~$�?燫�����-%���er����3�>$5�F�"������t������aO׾����aJ��C`�b�O�O�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >{C�<-����뾭����ο@�����^?���>��/��n��>ܥ�>�X>�Hq>����螾d1�<��?7�-?��>Ŏr�1�ɿb����¤<���?0�@�yA?��(��쾓�U=��> �	?s�?>�H1��O�+���Q�>g7�?]��?#JM=��W��	�a|e?��<o�F���߻�&�=*'�=h�=���J>,]�>����.A���ܽ\�4>�څ>�"�.����^��J�<2~]>^�սpQ��"��?��a��m�� �y���#w�=
�I?<^?�U½�d? �q�u�Ϳ����ܚc?�m�?�)�?��G?����^!�>fH۾�76?݋[?"�>9���q���=��t>¤��<U��^J�A�<A�>�f�>������A��S+U<t������ƿ��$�6|��u=#�ٺͭ[�g������wU�q,���lo�l�轜�h=ϕ�=ÇQ>|f�>W>�Z>�dW?�k?CK�>j�>�a佁����ξ�z�t?�����K�������棾HP�"�߾E�	�������3�ɾ_,=����=X.R����A� �L�b�~�F���.?�w$>�ʾd�M�.�,<�cʾ乪��i�������1̾A�1�e%n��̟?��A?8��� W�� �])�㘹�ĮW?�����ା�g�=.U���=r�>��=h���3��lS��i0?S?�y���o��.@*>�� �e0=(�+?�?93T<��>E:%?�+�(S��Z[>2�3>�֣>��>�	>R��V5۽z�?'�T?�4���Ȑ>mp��M�z��a=�	>.5�t=�'�[>L��<쌾n5W�n���l{�<�(W?Q��>��)��da�����Y==��x?��?.�>b{k?��B?\դ<%h��t�S���bw=��W?*i?a�>����	о����P�5?�e?��N>	ch����L�.�MU��$?�n?_?̀��&w}�}��z���n6?�{?T!k�&몿-�'��䪾 ?���>h��>�>�0I�>�c?~hx��@���g����9��#�?~9@`O�?{͎=,�=\u8����>��>��c�7����|ս!Ծ'S\=V:?B�2��(�/���N�g�N?�W�?���>'������E�=�Oq����?�L�?$��9�»g�U;g�Evݾ!k{�h��<��U�2p�����3�I���x������0M�vD}>�@�ƽ�?��o�'��_�ȿq�������ΰ��(?Y��>�-׽�ء��kl�r����.G�f?H��MY��M�>��>5���������{�0q;�����>N�	�>	�S��&��Κ��2�5<W�>���>M��>]*���轾�ę?c���?ο[������c�X?3h�?�n�?tq?�f9<c�v��{����-G?c�s?'Z?op%�E>]��7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�^�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*�+�+��<A?�2>���I�!�C0=�UҒ�ü
?W~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�3N�����Xe����@y����?N^�?i�?ӵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Pj?���� ����U>	�}?n�>��?���=M��>���=��Z"/� A#> 7�=�>�Ѡ?بM?FX�>��=$�8�D%/��\F��HR�!���C���>��a?|vL?	Fb>K��jV2�_� �xͽOv1�]1�W@���+���޽�\5>>�=>��>*�D���Ҿ�?k���%ٿ�������k8?D�l>i?�s߾&4���-�=$QY?�j�>��f���5����� �?���?�?�b�U½���=�;�>��>�ni<`Z�V{Ҿl�>t�0?�L)�eY��'d\�Y�a>�n�?vK@凴?�z�k�?��p��Y��9]�7����>h�2?�k��|�$>+�?��=��c�����Q]y�O2�>cݰ?t�?c�>�Kb?o�l�g�6�q2=�<�>��f?�
?~B񽎅
��g>���>^�&�(m�����_V?7@G�@֏W?�§��=Կ����������-�>-��=?U[>B�����=w��������=];N>!ҧ>��{>`>^>&(?>_8G>9�	>l҄��+*��Ϡ�7���f,=��"�i��w�Z���l��n�r������l��|񽚑Ͻ$�a��,�g�d�EJ=9�L?Kj_?lv?6�(?�w߽fTW>|�Ⱦ��=���1�x=~y�>�XY?Ȳz?WVD?eā�o�Ѿ0�Q�G�f�����SK`����>j�=�@�>���>���>n��<�c�>T>>kX�=�4=>� �=�ء��>ۼr>�>��>l�a>�C<>��>Fϴ��1��j�h��
w�m̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?%���z)��+���>}�0?�cW?�>���T�1:>9����j�5`>�+ �}l���)��%Q>wl?g�?>�W>��$��:���9���}����>��)?%���Y���{���K�J�-�(>��>Z=�s�te���~�ŷc�-Ñ=p�8?(^?"��Խ�MZ������_x>k�^>�!;7ſ=��?>}6��r����@��$k;噤<�Y�>�N?V�+>�Ԏ=��>kB��	�O����>�B>~�+>��??�%?�?��䗽-���)�-��w>zE�>$�>@�>=tJ��*�=}S�>��a>O��/y��)��}�?�$�W>N�|_�W�t��lx=8`�����=^�=� �0=��w%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>?N��^���щ�p*��� u=��>�TW?j����?���ל�\�?>�?{� ��y���#��Q:{��_�>T[�?>��?~eh�����=A��i�>:��?vi?���>�� �Q/��X~�>sK?00?)��>(e�m��MX(?�D�?�v�?ń>��?�)Y?0�?�0P�=�T�ok�����e~8>s?�$?��>:���6Z�}n��ǽ����H�&iE�X��>��6<'�>�O��ֵ?�	�<>b2h������v�לe>�ω>�W>�j�>v��>AZ�>J�>�-W�]����D�;-���K?���?)���2n�CO�<W��=�^��&?�I4?*k[�{�Ͼ�ը>�\?l?�[?d�>=��O>��F迿5~��s��<��K>)4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��)S��GB�>�e!?���>�Ү=�� ?��#?�j>2)�>aE��9��P�E����>��>I?��~?��?�Թ�}Z3�����桿��[�|9N>q�x?�U?�ʕ>)��������jE��GI�����!��?Ttg?�P�]?82�?��??"�A?w(f>���ؾ�����>O ?P��&�@�� '��K
���	?�?\��>#ɒ������v�C����d?��Z?�(&?@�+�_�EIƾ=(�<�� �����:<����{>�>�𐽰K�=��>�z�=�lm���9��d�<��=��>s��=ӧ:�����h.? ��y��I�=S0n�j�>��v�>n�>	$����^?[׀�����ɫ���k��9ҍ?t��?�r�?R�ͽf�Ew2?!��?��?�\
?����[?ﾠu�Ad��'-l����u�>Ӈ�>�|�����\����������r��Q)�>WC�>r9�>�	?��>�>U�j��1�UE��� ���]����O6�(�#�eg ���*���^:���;�+��Nj>���B�>Ym?{A�>�/>Ì?s����>:�5>Y�>�c�>�wB>~�3>��=��)��Ľ�KR?�����'��������3B?�qd?E1�>xi�>������0�?y��?s�?�<v>�~h��,+�_n?�=�>u��[q
?FR:=�H�=�<�U�����4��H
�5��>�F׽� :��M�nf�Jj
?�/?���ċ̾�;׽����,�=��?ø(?�(��|Q��l�r�W�PI�?L���d�Yt���#�~ l�M̎�E���9��p�*�]=(?���?�� ��d⾟ڮ��k�>�?���V>��>�Χ>rX�>�l>d���1�A,^��Z*�|���D�>}{?hό>�lI?(;<?�P?��L?t�>��>ƪ��Y��>*�;��>���>\�9?�C.?n0?4�?v�*?��a>���������ؾ=�?��?�n?e�??t?b5�������o����g�A�w�"䁽e=�=�@�<C�Խ�tq��)X=Z;R>oX?���`�8�D����k>��7?���>s��>����.����<�>_�
?CF�>  �V}r��b�hV�>���?� ���=��)>Q��=�����*Ӻ�X�=.���z�=�@��ɂ;��\<6�=Y��=�'t��s~�V�:Fk�;z�<�s�>_�? ��>nD�>�@��?� �	���a�=Y>vS>�>2Eپ�}��Y$��L�g�@\y>w�?z�?'�f=j�=b��=}|��zS������������<�?J#?�XT?���?Q�=?�i#?�>8+�wM��}^��0���?k!,?n��>P��E�ʾ�񨿜�3�ܝ?�[?�<a�n��<)���¾  ս��>�Z/�z.~�M���D���������}��(��?ӿ�?A��6�iy辸���X\����C?�"�>bY�>O�>t�)���g��%��/;>ʉ�>�R?	��>e�P?Y�z?�-]?G_Z>��<�f����{������i&>Bu??�K�?��?Hx?�g�>�n>�c2�
�㾵���
�)�s �C�~�^^^=P�^>х�>���>1x�>���=&��~���m_D����=9/p>���>Or�>���>0�{>�@�<��G?���>�\������줾cŃ���<�Ȟu?��?��+?�-=�����E��C��/M�>.o�?J��?�4*?5�S����=�ּoܶ���q�o*�>sܹ>P.�>~��=gF=�`>��>Ġ�><�>b��r8�kM�/�?	F?���=��ſxRq�<,p�����Q�z<2���v'c��ѓ��nZ����=�s���/��?��GW\�-h�������W��;Q����}�J�>ro�=�_�=hc�=t��<��μ�y�<�D=&�<�=2�u�vQl<8�;�|���	���M/�:S<bjA=^̻|�˾�y}?�7I?e�+?��C?��y>J�>B%3����>����0?y#V>�Q��l���*;������"��J�ؾ��׾jd�YƟ�S6>&�I�ͯ>�m3>l)�=s��<8��=��r=�^�=�O��='��=Ɂ�=��=���=Ѽ>�:>	8�?�r��Ң�;=X���M�)�@?u�>Z��<����O�5?�=[���l��,B�ҽr?E�?4��?j�?l�����>Ӗ�����>Z>��$�$�m=�=Š;����>�+�=e������6��i'�?�� @��'?.܄�����{�>��#>Ѽ�=�I���6�V�/�d,!�7�(��@?7���꾗u^>!�D=�L�aʾ^=Y/F>⚆=�
�9c�h�\=��'�t�-=��~=]�t>��9>]��=<�P&'>M�;��w=@=>x,�`�������r=�<�=��=>V4>3��>?�?�a0?(Xd?�6�>�n��Ͼ'?���H�>��=�E�>P��=|rB>ʏ�>6�7?o�D?�K?�>���=	�>��>D�,� �m�m�9̧��<���?�Ά?xѸ>��Q<��A�����g>�C/Ž�v?(S1?�k?k�>�U����9Y&���.�"����b4��+=�mr��QU�a���Im�4�㽯�=�p�>���>��>9Ty>�9>��N>��>��>�6�<}p�=Aጻ���<� �����=�����<�vż×���u&�8�+�/�����;g��;.�]<{��;R$
>��>3�4>>��=s�t�U?>FH�0p�-�=s���H��TO���m�t��S�ֽ�gK>Idi>��-��=��[��>��N>���;i��?�,~?��@>�����找���=��k�2�>��<H��~�=�d�[�gZ����[��>Yߎ>$�>��l>�,�L#?��w=��Yb5�~�>�|�����*)��9q�#@������ni��kҺ�D?�F��f��=i"~?��I?^�?ݍ�> ��φؾM;0>�H����=g�*q��h����?'?���>�쾤�D�W̾~��kз>z\I���O������0�J���������>�T�о~3�^f������ƌB�
jr�c�>r�O?��?B4b�G_���WO����+ꅽ2t?$�g?�>tD?�I?�ۡ��f�$|��!T�=��n?Ӭ�?�@�? c>�n�=qO����>a?��?���?��s?h�=���>�C:�:>�v����=X�
>�p�=q��=w?B9
?U�	?��P	�i���T7^�g^�<(�=��>���>��o>���=�{e=s�=��[>3��>�&�>,�d>y�>5.�>���1��n&?���=!��>��2?�C�>��X=:!����<�e]�tB��.�[���(�߽��<�MH���N=����>C�ƿ��?b�Y>����?Gv����?���V>�T>~���W�>NKD>�w}>Xӭ>|�>�>�N�>{*>��(� >-��'#+��4���C�I����=-�����"��2���;���@��Jv�b�(��d::��5=��?�K�������=C��ʭ���?�|�>K�i?>����͜>���>b=�>|d��돿Knl��	޾���?�@�3c>6�>g�W?S�?O�1�3�oZ� �u��&A��e�+�`�+፿l��� �
�`����_??�x?�vA?ל�<�/z>.��?m�%��Ώ��#�>�/��#;�'<=�6�>b.��m�`�b�Ӿ�þ�2��HF>�o?#�?HT?IV������>�'H?33?�	�?i?,?Rp?1�H�a6'?�7>G}?�F(?g�/??n;?�w+?�S�<Z�E��$��d�Ͻ%����]�^ �w�����	f=J� >����O�[�=����~�0>�}=0�,�s�>���=�?�;,ĸ����>Ay]?k4�>�6�>F�7?t��?8�����[!/?�D4=�����M�������%�>��j?��?�?Z?�c> �A��B��[>�Ê>"�%>$�[>��>�����D�b�=x�>V>@|�=�xL�L���L�	�\����p�<1�>-�?�2;>��i�il>���M�u���]>��R���	�qO��\?��ʗ�s��>�pP?�K%?ɱ >����̽��b��(?�H?�51?.\�?��>�4�[�C���E�R�)����>���=�	���Z���k��eC�\���#>㲰���c>���W�޾��n��J�Q辈(G=���w�V=�����վO`����=��	>����� �g.��������J?�sn=�O���tW������>��>d��>Kv3�t|���@�H٬�af�=�,�>*:>�㚼���ɝG��(�(v�>�2N?A�^?{�?Ʌн��`��,�֒ ��fо9��� ?3�>j$?-�#>'�->��n�XO�B�a�؜]�r��>	�>�j��>_�����J���cQ�8��}?\@x>�`?wJi?�U?��p?�?W�?;�>CZ���ľSc!?s��?l��=8p��XJ*�h�3�Ί\��E�>�7?�V �
�>�>?69?�0?�P?��?.>z��qL��;e>Nl>6.R��V��f>)yG?�q�>%/[?��?��>�4��þ� G����=/N>b2'?�� ?�M?��>�2�>f����=�$�>t
d?�s?h o?S~>N�?:�>@K�>✬=@4�>V<?ү2?�| ?�cI?5�O?���>���<47���0���L�����ʼk�=�J�=�2�<'p��z|������D1=V��<���<9�ܽ6�����<���=a^�>0�s>���N�0>>�ľ�L����@>Sy��0L��?���a�:�3��=v�>]�?W��>kE#�Dђ=���>�>�>���74(?�?�?S$;'�b���ھ��K�}�>HB?���=H�l�������u�iBh=��m?t�^?��W����L�b?��]?2h��=���þz�b����f�O?=�
?�G���>��~?f�q?Z��>��e�(:n�%���Cb���j�Ѷ=Nr�>KX�D�d�}?�>_�7?�N�>�b>+%�=ju۾�w��q��j?��?�?���?+*>y�n�T4࿸����9����]?�P�>��h�"?����^Ͼm������,�j����z���R��f���D�$��h��!�ս�=��?�ls?�&q?d�_?�� ��Ud��^����eV�<��F���ZE���D��TC�<�n�1t�)��G�����H=gE}�O�@��=�?W�'?z�1��5�>}�����;/�C>���P��b��=6���r�4=syQ=��e��7-�!��_\?�˻>�r�>�[=?�[�(o>�_�0��8����'@6>	ǡ>0?�>]��>�3���.���9ʾY憾��ͽs=i>h�_?�>?.b�?�К�/����pw���I��	R��o��r$>&�o����> ��VS�ʆL���J��9n�Ɩ�ݖϾ��i�=#�Q?�A�>tG>���?{�?�0��S�e�پ1�/�t�����>��?��>(�?>K8������>p?R7�>*�>���t�2�i���2g6�o��>64�>'<?�)q>���l]�4�L��U�6��qE=B�\?I핾�b��}}>YtM?��=���~>ycs����|�����S�ܔ�=2�?�6>fh>�о�	��Mb�ؤ��7)?yH	?Fz��$�'��	w>e=?,��>�	�>��?yY�>5���o<�?(�`?�K?D;?=o�>�V\=�К��ǽ$U,�z�=�ˇ>F�K>uX9=Zյ=L�%�|�Y���*���>=B��=W=��X��>r<)`��]��<���<:�+>��пG�D�ȁӾ� �� ��F�������������l�s2��Rl���s��Ƚc<y��E��ɘ���OV���?'�@h�����	�������R�<������VG���=�!����� ���QQþ˚��0p���IE�䚐�/�E���&?7�V��Rֿ%8���+��X-?��?�C?���q�c��/��N��>��=���=3�'��̃��Kֿ&��^�?k?=���$��?(��>�@>H��=�&6�T�S�v>��?�T?���>ൾC����Τ�ν���?��@�|A?��(����3V=#��>��	?c�?>S1�JI������T�>�;�?��?�rM=h�W���	��e?r�<��F�n�ݻ��=�:�=vJ=����J>U�>ׅ��SA�&@ܽp�4>�څ>d{"�ª���^����<�]>p�ս�8��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��=i��^�ѿ
*������=R뱻4f	�<&����ս�a}��Bž�愾�>���=���=Ah+>�U>(�[>Z�I>9uk?L?b?G�>��M>��@�b��tj���T<�ܭ��@��^{��=8��r��۾����+�`�~G�nG���;���=�TM�8����/��e��I�I>?���=��q	?��W<�ɾ���ż 꼽�4Ծ<�-^j�=�?�I?�y��Odf�A�����<U늽'CK?�vz���
�*pþ�r�=�I)���=�>�S�=�@߾��:�8O��*?��?M����Ɲ��O>aiϽ���Q�%?���>`v��.o�>��?�p��.���>+%X>Y@�>Ä�>:y�=^Ϻ�-�뽎�?4FX?����s��w�>��P������=��=H5.���*}�>��s=;	��3�j�'m��C2=(W?f��>��)�b�.a��v��I==��x?Ғ?a,�>�zk?��B?P��<�i�� �S�(��kw=��W?#(i?,�>Ǒ��оq�����5?ͣe?�N>�gh�^��Y�.��S�=$?
�n?_?t���Yu}�����n6?���?��L�m٣�����Q��a5 ?�?�>#&�>�B��2�>��?^wR�a.��Bخ� d���?ii@;��?)g=�9�o�=M�?q�>V�˾�bԾS�(�O�`2��.�>1}L�㖞��5�����U?MË? �?�-k�g�s��=����%��?i��?�˯�=���`��Tj����U=oʇ=�ɐ��PĽ>@�Q8�gtξZ�������<9�M�>H�@�f����>�x3���޿JJɿ�1��uAѾ-,U���?�b�>�}�Iϭ�7_j�`�v��fG��KO�ڷt��P�>�2v>�M%�����F��2�*�#[���U>�ȼ�>G7{�����P��!8�=��C>�=�>y#
>�(��W�þ���?%H�0o����8�ݾ���?{�?��?��F?��s�g����=<^d`?N�?�<G?
�k���x�n$=$�j?�_��wU`���4�uHE��U>�"3?�B�>S�-�L�|=�>���>g>�#/�y�Ŀ�ٶ�=���Y��?��?�o���>r��?us+?�i�8���[����*���+��<A?�2>���I�!�A0=�RҒ���
?U~0?{�e.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?	�>4�?�V�=���>k�=�ӱ�c�P�g�!>�=�=@9���?�wM?�\�>��=z�9��U/��WF�wDR�;����C����>*�a?l�L?F;c>�H���2��� ��ͽ�2������@��^(��ܽ�G6>��<>Bb>Y�C��`Ӿ�a+?!������"���\?�a=?}�6>�?�>斗�������߽ڌs?��!>dӾ;���q{�u�i��ƥ?׶@[�?�G�-=�=�af>�O�>f�>��G4_���O��>�*`?}u����)I��4>W�?s@�y�?����/5?�� �%����~�N���Χ��\�=Yt-?��𾸼a>�>�f>[聿UTR��fN�>T�?I�?��?�j?��s���"�0G=u�>�ee?�	?���:� 	��v�>���>P��<��������B?�@��@��b?{����hֿ����\N��M���,��=���=�2>��ٽA_�=�7=u�8�=����=z�>��d>q>4(O>�a;>��)>���K�!�r��W���R�C�������Z�D��Xv�Sz��3�������?���3ýy���Q�	2&��>`�)��=N�O?�V?�]�?n??O,�_��=��ԾW�B��1T��ZD<�(>8?0P6?�0(?'"=QC���/e�:
��rh���5X�M�>�D�=���>��?�m�>�;��:>�e>���>��Z>r,=/�.�G�=]MP>b��>/v�>�Ĕ>�s<>��>䴿�[����h��ru��ʽ�Ģ?dќ��4K�l��Q���R����=��-?�;>#��LKп����JoH?¤�� ���+��>��0?�rW?�>�\���MY�O>%�v�i��G>���z�k�_�)�0�Q>�?��f>�u>,�3�ee8��P�mr���;|>616?඾�g9���u�q�H�"rݾbM>s��>��B��`�����͆i��]{=	w:?��?�C��}䰾�u�SW��P7R>�=\>�a=Fa�=<BM>v�b��ƽ�G��U.=��=��^>�?e�>�ǣ=F~�>l䛾=L�I��>V@>��'>_�6?r�#?J���ؽe��r�<�<~>��>\�>��=^lU�:�=���>u�w>R�+������3�w�Y�ʢA>���aQ[���o�ަ8=MlR�(�>oS�=1��s4@�3�9=�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿc�>�0�e��7-����u�B�%=]��>�H?���06T��1?�(Y
?-?���u����ȿ�{v�2L�>7��?I��?��m��X��� @����>���?bpY?e�i>�۾Y�Z�	�>��@?+�Q?e�>�m�R6'�X�?�Զ?ʅ?0>J�?Y+J?���>e���uW�ih���ʖ�8�M��;�>�1?�@>�y��9�d��?�z��8�?�/���>�ϴ�s­>�+���D�����=���T�����j��>�}�>RQ�>lR�>��?��>%4>�Kt<4'�Ǔ�����K?H��?����m���<��=�_���?��4?x?J�J�Ͼ^Ш>E�\?���?�[?E��>̤��'��y޿������\�<��K>m��>�F�>"��?L>XgԾ�C�x��>�>�ӧ��L۾'{���N����>/K!?���>A>�=� ?��#?�j>�E�>`E��=����E��&�>�1�>dX?1�~?��?�鹾5x3�^���᡿�q[���M>1�x?�3?w�>T���Xi���E���I�Bh��z�?�Qg?x��O?�7�?�??RA?�e>�p��ؾ�}����>��!?��f�A�J&�7���|?V?��>����}�ս�ռ���~l��?)\?�5&?ř��a���¾�<�Z#��bV��H�;s�E�?�>�>Ϛ���}�=L�>`Ѱ=r0m�56��!h<NY�=S|�>���=].7�@�����1?�Ak=��^��ͽ�
����$�Ѩ��H�>L@�^�?Ӑs��?���J������O&�����?��?���?FC&�la���!3?QB�?�?#��>�����ξ�����+��n�=���}�=A�v>+ <J�齎Կ�ţ��H���II�f'����>��>��?ZL�>�q>���>�Oy�q��{_��I���c�/j���9�I�'�B�O*��{(-��"��`ZѾ>����>�9m���>��?�X>��g> ��>����>�PO>
�V>LN�>ǔX>-�S>k>���;��߽YJR?C����'��������(B?�rd?�<�>b�h�Y���Ǿ� �?���?bt�?y^v>yh��%+�Qq?2:�>���d
?L�9=C?�{��<�_�����x���w����>�D׽:�;M��5f��j
??.?�+����̾JW׽O���"Ž=�k�?H�*?�-)��Y�f(d��fY�{eU�,S;;[ov�3妾;�/��q��r���s���xv���$��F�<��?���?M�
�b�о��hmc�66�>>�F�>d��>"��>L�>�оTVB�|�_��w"�ݸ���l�>��?A�w>��Q?�:P?��$? �f?i��>-$>g�о_??"�?���>J�>�-?0�4?��c?�#�>6�>Z(�=���*?��&߾W�?��?J�?xB?#C?#�߻�2k�i� � :%=�;��5��a(=��=K�9�l���x�>��>��?���,����2f>]t2?��?4�>>��u?P��:�=�R�>|�?�ų>z���on����'T�>�A�?��)��=�N:>�e�=v%(�*����.�=��S=ն>=�6��	����=N��=�M�=3����Ƽ��X��S	�;]���U�>��?;��>펌>w������P?
�9�=�54>ɣV>��>��Ud����g�f��JZ>Ts�?�Ӯ?�y�<���=� >���ޱ��8��I�Ⱦ֥=`��>��?D�T?���?qGB?�_$?�6�=�B��j�������?}!,?ي�>���C�ʾ��݈3�}�?�Z?�:a�����<)�0�¾��Խ��>v\/��.~���D�Ƭ����J�����?��?�A��6�oy�j����[��ȔC?�#�>�Y�>+�>=�)�U�g�%�l2;>���>�R?��>�DV?,v?�QU?n�\>�O4�Y޳�����HC=��>�=?ԅ�?���?�~?�D�>V�:>GT!��龅s��9��E�����6GO���^>�S�>Y0�>/C�>���>������	��:���C=]2}>o��>~D�>�0�>6�>��=��G?K�>����k��%Ԥ��H��4�F�%�u?`t�?��*?��=��w,F�5S��)��>�/�?Gث?�<*?��U��%�=%�fT����p��	�>q<�>w!�>O�=�'I=�>k@�>�V�>B������c8��F�h�?!�E?��=dǿ�]|�� ���l��b$=o󂾆�1����o�.�7=Vɭ���(�)�����P�+Z������1��Τ��Yqy�Ŀ ?��=�
>|E�=�?�<b���-:$��\=>O-���B=�O���<��޼�`��ͻ�@�;�/�<�F=�RP�m�ƾw[z?\J?�94?
UG?��W>1�>rf���>gX��?�?�e=>����T����*�Av��2��א߾r߾�Ei�w����>�����>�2Z>ȋ�=�<���=TՒ=��=t�<��%=��=��=��==F�=��>6>�6w?V�������4Q��Z罠�:?�8�>`{�=��ƾb@?��>>�2������~b��-?���?�T�?@�?Oti��d�>C��E㎽r�=o����=2>���=��2�>��>��J>���K��x����4�?��@��??�ዿʢϿ:a/>�o>>/
�=�QH��33��	[�Y{J�U񂾅�"?�0��߾��>�=ފ��ھ�j1:vbD>��=�^�]^��f0=E&���	p=��=1E�>�B>��=۽����=�0�<�G�=E�E>�Dd�
�7��$(����=/��=5�T>�c0>,�>.s?yZ/?�[`?@��>�o�wݾ�ƾ�>Bl�=wn�>퉏=<�^>Ե�>z�8?��C?xI?��>Ӱ*=[3�>�՝>�r*�q�n�33ݾ����.=�\�?3�?��>y�/<�P��*��?�������?ab/?�?ⵤ>D�p����F������<j>�>��g=̌���1�&�����O����>���>D֯>gH�=w}�=�D>?��=5�?њ>u8�<�Y>���=�)r=�f�=7��<�D|����#��b�ʽ�'=
��$j���ý�1���,e<Xa#<WV>~�>�+>��|>.��<�o���9�<H��5��ɸ=�����ZQ���r��܇�}�1�j@0���>3!�>�2��Z��K
�>Qj>��>v�?�+�?�	>fHk��;Z��ݢ�P�����b��=�� >�c���'�n�\�.pD���ؾ���>Q�>_�>f�l>�,��1?���v=�"⾎^5�;�>�S�����K#��:q��;�����
i�i񺒓D?�C���i�=i~?�I?`��?�y�>SO���lؾ�X0>nH���u=��L�p�Ӓ� ?�'?n��>��`�D��H̾A���޷>�@I�2�O���V�0�^��0ͷ�2��>������оn$3��g�������B��Lr�X��>!�O?��?X:b��W��GUO����V(���q?�|g?,�>�J?�@?�%��z�r���v�=�n?ȳ�?O=�?�>(�=�;��LY�>[0
?3��?�/�?�/t?�W�����>��=�}>����w��=	B >!7>�G�=�\?�?�'?Tp��$�,��l& �77x��P�<�3�=�!�>	�>��t>��=��
=�&�=�5h>�Ģ>b4�>s�h>H�>x�>�o��X�_�&?���=%�>(2?�2�>�Pb=�9��.*�<�]F���B��#.�� �����X�<u����W=�弔j�>�dǿ
�?�U>(9���?�*��YD��)S>R>֥۽�@�>H�D>��~>@��>��>��>(ȉ>�(>�ڷ��/.>��&���G�zHY��,�w<��HF1>'�W�`0��d�0�E���=*�w�k���Jv[�����ȱV��=.	�?�)o�񢉿�#%�8��<�R?�B�>6�C?Y�(��:��"���?+��>��վG���y�����@��?��?�Ec>I�>�W?K{?-�1�3��qZ�l�u��A���d��`��卿K�����
������_?��x?sA?�Ύ<��y>A��?��%�g��� �>�(/���:�5o9=��>�̰�g�`�a�Ӿ�þM��/WF>�ao?�?�/?��U�0;�=&�z;�eB?z?6�^?N�1?�u�?x�>�?�D>D$�>/?��?�cH?��D?��'=��<�>���=rt ���þBő���������V��ռ0$.<�����1���t;Z"z��(�9�4��%�=�(�=�Ģ=|_$<��>EX?>��>�@y>�3?��-;����p�-?y�<�z�� ���R��H������=��i?;��?;nY?�N>�M�mtL��E#>���>�0 >�U>a��>���I����=R�>lH>vޑ=����z���/����o�<�|$>���>'|>r����'>L���"cz�\{d>��Q��ٺ��S�;�G�W�1�cw��%�>��K?M�?��=&<�쵖�0<f�?:)?�C<?^[M?
�?�W�=ƾ۾[�9�:�J����_��>��<����������y�:����:C6s>���8䠾�Ub>P���B޾>�n��J�����L=�x���V=��]�վ�����=M
>������ ����(ժ��,J?[�j=�l��ULU��y����>���>Oخ>�7:��w� �@������=��>�5;>�v����G��>���'>��<?,�n?�ʊ?)"���b��D'����i�u����<t3�>���>\W#?�
�>�]�>���h�Amp��i����>��?���P.M�YW��N�뾘�G�/^�>��?)�=��>	�P?��G?ok? +5?�2?�q�>�8?���i�?�(�?��=�I��A�)�&�8�I�L����> +?'w.�a>c�?��(?��+?UGW?��?��=�	��DM�?Y�>@��>�SQ������!w>I?j�>"�W?��?IQ>�<2�G����Yx�.T>�>>2?"�#?ۓ?�Ǳ>���>Qŷ��<U]�>�b?���?�cf?���=q�?��!>%��>�?�=̚>���>ɮ?��D?��g?�NE?��>��<I���1\����ꏥ�v�B�J�F<A�?=�A�eׅ�~Eż��<<��i�����-��=��&���F�ڙ���_�>��s>
����0>�ľM����@>�o���N���܊�<�:��ٷ=ꃀ>��?ө�>;V#�»�=��>G�>���N5(?�?C?E]!;�b���ھ�K���>PB?��=��l�d����u�(�g=��m?��^?��W��%��N�b?��]?>h��=��þ{�b����g�O?=�
?2�G���>��~?f�q?U��>�e�+:n�*��Db���j�&Ѷ=\r�>LX�S�d��?�>o�7?�N�>0�b>*%�=hu۾�w��q��i?��?�?���?+*>��n�Z4����e��X"]?ZS�>򬧾�� ?��@:ξu���p��������C��E����꠾#��Jjz��ӽ���=�?:�w?� l?��\?�{�Pe�Z^�2���]P��#�/�K>���C��E�NCn�+m�����J��� v==�y��J;�Ю?�?@�S��O�>�<�����V��)��=B�����,�,��`���F��<��M=�� �nY �~����?b[�>��>I?D?3�O��`C�� (�`
6�)�߾�R�>Ә�>��>Ҡ�>��<,�%R���I����뷽�>san?�Z??��o?���S�7�R�!���\�9 n����>C�	>�u> �����Q�ŉE�=���j�C���&]������g�=S�?	��>��>Ip�?��?E'��~Ⱦ�ό�*XQ�X2�8��>�rw?�P�>��w>탄�wwF�?��>b�n?� �>*̩>3 ���'��w|��)�-'�>ͬ�># ?��~>�!*�2b[��y�����#L9�Q��=��h?т��\�mE�>��M?Å��<���>i�_��#��/�� �_|�=��?�a�=E?>�ƾ�B
�+�s��Ϗ��+?�q�>�`��ߢ��>Ș)?"��>��>�Ć?�ף>�aӾ]�=��?Ltf?�P?/	/?���>�H6=��Y�+���$(�$\�<3�}>��?>�f�<;��=�������#�=��=<V�=%�r�3鹽=�<���<U�;=~�*>L�࿽xG�H���p�t�޾o��ާ�~; �g����ƽ޸þ�ؕ��5V�'�L�����R��녾������Q�
q�?#��?β��$���n���9���o���G>?�*E���U�;z�]rѾE-�&d�y �tP��rh�XD�U�'?𺑾ڽǿʰ��E:ܾc! ?�A ?-�y?d��"���8��� >SF�<)&��!�뾙�����ο%�����^?���>��2��J��>{��>y�X>PHq>���g螾�0�<l�?�-?��>��r�#�ɿN����¤<���? �@�}A?�(�O�쾃AV=���>-�	?��?>�51�Y7������G�>�8�?5��?�N=ֺW�Q�	�ue?Ff<Q�F���ۻ}��=�=�E=���tvJ>�Q�>���[A��@ܽ{�4>Ѕ>b�"����i�^�ۉ�<F�]>סս�A��8Մ?({\��f���/��T���T>��T?+�>�9�=��,?X7H�e}Ͽ�\��*a?�0�?���?<�(?�ڿ��ؚ>��ܾ��M?fD6?��>�d&�/�t����=@2�ᗤ�M���&V����=-��>A�>V�,�����O�HK�����=�a���Ŀ-)�U��O=?!�;�s��WBҽni����,�/�����f��P���6�=��>tGH>D�l><�F>�}Q>��W?$t?���>4�>"�"��R��#$����"cz�/�
���t�o(��8��vR�- ��;��\�����.{��� =���=�6R�<����� ���b�<�F���.?fx$>�ʾ��M���-<.pʾ����~Ԅ��ॽ�-̾�1��!n�c͟?M�A?�����V�f���X�鄹��W?MO�̻��ꬾڣ�=歱���=b$�>ቢ=V�⾈ 3�9~S��h0?�A?"g��w����)>�� �H=��+?�{?O|Q<=;�>[(%?�N+�ͺ�� [>�3>��>���>g�>�����۽�?�|T?A��	�����>y���khz���_=�>3�4�����[>��<�׌���R����ue�<�'W?Ș�>��)����_������N==(�x?ؑ?�*�>zk?��B?k��<g��>�S�K��ew=�W?�'i?��>6����о݁���5?Z�e?��N>�jh���5�.�jR��%?}�n?C^?󸝼�u}�|�����5l6?L��?�[� .��mc=���m�;��>��*?�<�>�Q2�D��<��B?�O�������W����F����?_v@w,�?TP�0Mf��B�:|��>[�,?L,���Xҋ����u_�<^�.?��򵗿-�z~�XT?���?�"�>h���'uԾ:��=@�w����?�Yx?m�о�V����bu�*���~[=�8F=[n&�H�&����9�:8оET�͠���f���d>�@��	�G��>󂢽{mݿޛ˿����վ�E���?��>}�=�-پ �Y�pp���U��[�$����H�>��>g���!�����{�8g;�������>Rx���>7�S�/������p�6<��>٣�>���>R-��8ս��ř?vb���Bο}���P��4�X?.e�?m�?�q?�7<��v��~{�D���.G?Wzs?�Z?g%�S]�Po7�'�j?�_���U`��4�oHE�U>�"3?�B�>Y�-���|=+>���>�f>�#/�x�Ŀ�ٶ����\��?ۉ�?�o����>m��?us+?�i�
8���[����*��+��<A?�2>-���K�!�M0=�FҒ�ټ
?i~0?�z�w.�	�_?"�a�w�p��-�]�Ž[�>N�0�$\�^�t��Re��훿S�x����?KW�?1�?:��X�"�06%??�>,���V�Ǿf��<fH�>|��>��M>(�_�J�u>q �3�:�_J	>��?�j�?�K?����H���>��}?b��>{�?��=b��>��=f���M8�I�">F��=D=�B�?��M?	!�>�7�=Pa9��6/�([F�;MR����D�C����>�a?�bL?qb>����/�$� ��νC1�W��4�@�rY+���޽�O5>�{=>#�>�yD� 5Ӿ��)?�p�i�ؿ������V��1B?���>=v?��8���u>(e?�&:>��Ӿ`����6n��üXQ�?���?~?-���z�<\[>'
�>~ï>m�=7w���6˾|}�=�:?�J��@��gi�C]>���?{;@�a�?�N����?
��P�����������M>,�7?������L> B?V#�=�+t�U�����u�\�>N�? �?3��>_Kj?�o�@ =���h=6��>Y&g?�_	?!%��ﾢ�I>g�?XP�b&������&c?b@HG@�Q]?�X��M�pR�����D���Qh�=�>};<>a\н<�>�j�=�����<>>W�>��>�Uz>��>��>G`�>����%�������w
C�����$B���(C�Շ��ŵu�f�����vM�4�νX'ǽ�����A�3����<�A�K�U?�a?��T?h�3?�,��\P��m���j>�S�=u����5O>�Qs?v�]?V�@?(6,<'�����Y����h ��ΐ�L}�>aq>���>S��>��>�z��-��>�{�>�*0>k�>�̛>v4>rm�=���=�>�$?��>�C<>��>Fϴ��1��j�h��
w�r̽1�?���S�J��1���9��Ӧ���h�=Hb.?|>���?пf����2H?&���{)��+���>}�0?�cW?�> ��w�T�3:>9����j�5`>�+ �~l���)��%Q>wl?=f>^?s>��2��M8�6�P�Z���Kp}>D�5?ԩ����;��~u���H� N޾��K>bν>A�/�L��������~��pi�"�}=*Z:?d�?1q������ڌt��ʞ��R>a�]>�Q=Hz�=�L>�b`�D�Ž�fI�A�+=R!�=^^>7�?D�>��=%��>�����?���>]�=>�'>��4?:"?zUK���ɽ�ć��8��U>�\�>�4�>��=�J��7�=���>��l>6x-�Tu��d��5R�X>X\U��rh�O�N��U=A�����=
�x=�����a@���=��~?�ç�� ��GP�$���)G?�	?��=�!#=�Q���������y�?�@�M�?�����U��+?Z��?+[��$��=x��>�`�>P�ϾgW�L�?}�Ƚ�����o�8���u�?�;�?�f8��g��^oj��->�%?cоȵ>@)�$����>����}�kWS=O��>rM2?ar��Ǹ��Ӽ\�?S�>�\���������U怿�m�>���?z�?�#e�急�@�M�N�?'y�?D��?٧�>6��J �@T�>4ZO?�"8?.��>��%�����62?Q��?��f?��=Ò?�J?7�?�+/��\����펿m}�=�>���>9��>���E;e�qi���7x���E���D���>��<�ݮ>�-������Q�=vG��ژ��u,=�t�>�(>'�n>��q>ˈ?���>$�k>�v��2<N�p,S�������K?���?����1n��t�<˝�='�^��&?6J4?�8[��Ͼ�ը>.�\?�?6[?�c�>���3>��n迿�}��ɥ�<��K>+1�>EI�>i��zFK>Z�Ծ�0D�*q�>sϗ>���><ھ+������dA�>�e!?a��>�׮=٘ ?�#?��j>�&�>�aE��9����E���>���>nI?�~?��?�Թ�CZ3�����桿�[�9N>-�x?�V?�ʕ>��������fE�u;I��𒽂��?tg?t[�d?82�?��??��A?u$f>����ؾ������>8"?�~���A���#�����G	?�J?���>+����nڽ��ʼ��������?
\?�s$?�t��z^��T��Jt�<�����9���;p�r��T>S>���#|�=Ob>�ݳ=�k�"�8��a<�ͽ=���>OU�=L68��֑�q�4?�w]��{��d3<+����X�~�c>ʡ?2.��N?c�¾&��Υ�[���+�3����?�'�?�*�?�x���b��!H?W��?�,
?bI�>ξ�־�B���Л��:���־�U�=��>1�_=�U���ʲ��v���������Я>�B�>T��>c�?*��>� >4�>Kz���6��V�ѧ�
�_��5��=2�*����������H�`���T��� ���L�>���O�>��?Pކ>�O>���>�p.<T� >�;>'�J>A��>�ْ>o�Y>ĭ�=��Y�N�S??GɾH*�v�߾R��KD?�\`?R��>��
����X���?�W�?���?}g�>��f��*�w?���>�ry�ߡ?=�9���<�����I��D���KO�[o�>�ô���7�&�L���e�"�?��?�x�Հƾ�Mڽ��Ҿ�R�=6�?�?C,��K��8y�(�j�`A�=�}=� N�]��U~���i������J}����+�|/�=��3?���?U
���.��[1c�j�>�3>�u�>��>14�>��S>L��R�7���u��#'�m�����> �?{*�>'#F?��@?�%K?�ET?�M�>��>]��O�>��/=��f>8��>I�O?X<?��5?,4?��?v�T>�������Ծ� ?��?n?��
?��?�Ɇ�xh�5t�V��ܢR�&���Þ�=��G=���0aƽ�3[=�n~>�g*?�J�� �N� -����>(�??"�>\��>1:��yC�tw�=�9�>�� ?G��>�4G�YWZ��	�x��>5m?@�m�(�+=�dC>�b�<T�����C�=�{Q��C������Ȫ=-��=�;[Q;=�X�<z�P=��_=�
A�U�)����>�?��>���>�A���S��@
���=�W>`�F>�>�kھ����gr����g��%z>7\�?F'�?RG=��=��=Ρ���C��^d�(a��}z�<��?E�!?9GV?�.�?��=?>�"?X�>������k{��c���v?t!,?��>�����ʾ��Ӊ3�۝?d[?�<a����;)�ߐ¾!�Խű>�[/�e/~����;D�0���5��3��?쿝?8A�W�6��x�ڿ���[��}�C?"�>Y�>��>U�)�{�g�t%��1;>��>kR?4�>m6P?D{?�g[?P�V>I�8�$3���0�����t&#>�>?�x�?�D�?�&y?���>vl>m�*��}�,����!���������A=9�[>gP�>ւ�>�P�>w��=�ý�P��K�?���=��d>-��>���>�1�>�Yy>3ϲ<�G?�W�>�������������{<� �u?�C�?��*?s�=���F�˗���;�>�=�?�Ϋ?�*?v�T�w�=o~弋�����q�o^�>e��>�n�>#��=�N=��>2T�>�U�>�p�9e8��4L���?M�E??�=:�Ŀ��q���i�z��A�;Jˎ���]��L���Y��y�=YŘ�=a�ޭ�b[_���������h����m��>�>|�=EE�=�d�=W�<t�ȼ_��<K|-=T��<��(=�G��aǉ<y�:�ȅ^��G��p�e�G<}�?=\���˾og}?�5I?��+?	�C?&;u>M~>�;����>�B��@�?�T>��O�o���|�:�]ҩ�W���e�پi�־�4c��ş���
>��9��>�G3>u��= d�<�|�=W?{=(��=���8r(=,�=m��=,i�=	�=]�>��>�6w?N�������4Q�^\�e�:?�8�>M|�=ׁƾ_@?��>>�2�������b��-?���?U�?��?�si�Od�>����Ꮍ�t�=$����;2>X��=Z�2�W��>��J>ۃ�K��9���L4�?��@E�??�ዿ��Ͽ+b/>��1>���=RTF��k1���l�V�C�7m>���?�6��4�	��>T9e=sD�-�;v�N<�aL>�k�=(��J�[�t/�=.ߔ�?��=~��=�6s>{�U>S%�=��	��B�=��0=1Z�=/X>�8 �w�����U0 =���=_�N>�Q>F5�>Մ?0?�@d?%�>Ye���ξ������>.8�=�!�>�Ȍ=��C>�a�>��8?3�C?ȀJ?f��>�T�=��>�>�.�/m��X�����<���?yކ?fd�>Xq<}A�@��h=�>nͽ�?�0?��?���>�U����6Y&���.�+���&�3��+=�mr��QU�����Hm�;�㽒�=�p�>���>��>BTy>�9>��N>{�>��>�6�<�p�=/⌻���<y ��p��=������<7wżz����u&�)�+�!�����;v��;ҧ]<m��;�>W�>���=��>fC:3����B> ���XT�~`F=W����?X�*�_� �|��.��d��5h>%�{>��ܽʎ��E�>a�>�&�=�.�?{�?B&+>'�d���@�f}��4 �E���<ɳ>A����:�ٴ^��Q�Q���>�>��>S�l>�
,��#?�B�w=8�Nd5���>�x��
���*��8q��>��y����i��>ֺ\�D?}E����=u ~?A�I?�?f��>F����ؾ�40>2J����=���+q�tc����?�'?3��>����D�W̾ዾ�η>P�I��
P�������0���!��@��>�Ī�.�о�3��_��w�����B���r��ٺ>�O?E��?1b�de���kO���춅��?��g?`�>�$?�G?=����f��/��Mq�=�n?x��?�C�?W>==	>(ir�e��>��?'��?٠?B�F?�`ݼ(�?�=l��=?�=b[;>?�>��>��z=@Y�>]�>2w?V]�=^�w'F��Lھ���N[��x�;��]>�@�>��&>jz���,=|=�Be>�>�!E>v�U> ��>n��>2������)?m��<��W>BG-?^0�>�f	>`����E�/}#=U_���U���C%��03����=���=�)�=(h�R�>?ظ�N\�?D�s>�"�T!?�W��$(����>p�=�lH����>:��<Ms>��>�A�>��b>��H>i��=q���h}`>3���^2��)X�#H�o���f=�B �,0�<vٷ�/����Q��X��1�
�.�e�$Ȉ�A99�n=>��?|�26��ÖT��SP���?�"�>�D?�/��.�|s�>��?��n>���8����х��s��5�?Y�?��b>�F�>��W?�5?c�2���1��Y��wu��@��ae�ƀ`��ԍ������
�j�����_? y?VKA?Yb�<�y>�~�?�}%�	 ��yf�>��.���:�_6=�	�>�k���b��-Ӿ�þ����LF>[o?���?�?.�U�Y-�)t�=�t ?ɕ+?��z?YT4?��(?Zн}�#?�'6>���>�E?d�;?��C?��?>�=6n�=D���@2=em��C]w�ϒ=��ک����;�~H=I4m=bs����<�=��^»��o�d�к��;6��<l=;�:��=P5�>�\?w��>��>��6?^Z�1�7����3�.?6�&=Vт�Ë�o��<F��� >��j?B��?�Y?�a>��A� �A�>M1�>e�#>��[>���>��󽶺D��=�b>��>⹤=g8H��7��+�	��g�����<�>i��>��{>ˁ��?�'>���O�y���d>��Q��º��8T��G�j�1���v�a)�>E�K?��?F'�=�>�ǖ��7f�h1)?5O<?QM?��?ጓ=K�۾��9�	�J�����>᙭<J��R���L���:���O:sVs>� ��G栾'Kb>����x޾�n��J�X�羈-M=~���U=d�� ־�4�u��=
>I���$� �����֪��-J?��j=Yy��dU�`r����>��>�خ>�C:�Gw�<�@�y���1'�=��>��:>U����z}G�(2�S��>�3E?._?4G�?��~���q�/�?����������ɼ=0?3��>�q	?��J>�ȵ=����W����d��F�W��>�!�>0#�~E�)�������y&�@�>�^?��#>_@?��Q?�??&�_?�(???�S�>B����ж��A&?6��?��=��Խ�T�� 9�HF����>{�)?�B�۹�>Q�?�?�&?�Q?�?w�>� ��C@����>�Y�>��W��b��A�_>��J?ؚ�>q=Y?�ԃ?w�=>\�5��颾֩��U�=�>��2?6#?O�?�>0l�>瞡����=)�>yc?�5�?��o?���=��?��0>
f�>���=�B�>�C�>"�?�OO?��s?4�J?�>��<v���鶽m�q��XV���|;��F<��w=D��X�u����Wl�<���;S۵��}�Mf�1�D��d��m��;m]�>��s>1	��|�0>��ľ>K��.�@>jx��	P��ߊ���:�Rҷ=.��>*�?꩕>{T#����=C��>�C�>����6(?,�?q?�!;Ϡb���ھ��K��>�B?��=��l�E�����u�V h=��m?�^?��W��#��O�b?��]?@h��=��þz�b����g�O?=�
?3�G���>��~?f�q?U��>�e�+:n�*��Db���j�&Ѷ=\r�>LX�S�d��?�>o�7?�N�>/�b>'%�=iu۾�w��q��h?��?�?���?+*>��n�Z4���������'\?���>]���B$?�	�:��о���P�����+���A4��B����M��D�*큾5��Q�==?2Dq?�bp?F�g?���Ϣf��f]��K���Q�E������=���?�ӂ?��/m�H��L|��K����$v=>��$3�<��?i~?�X�R��>a�p�4���i����^=:žRC�=�<���ϫ=��=��e���^����?���>�p�>C�b?��e�d#Q��2�f<7�%�߾�"�>4�>>��>N%�;��a���\�No�߅��$�;�\8(>+Rh?B,L?�1�?/x=�b�ꮊ����h=(b��[�>��|>��>�����M�"�E��E�K�n��6׾�B����sC�=t�?��>!p�>MD�?��?l���J�&�v��Z�f<���>|�?���>s��=9�=�9���>�8n?���>z�>�^��p�#�c$}��*ݽ��>-M�>�r ?��x>�)��~[�np��P����q8����=�[g?�8���e�K]�>i[P?�A\;U$�;�՜>h>X��������-�@��=�?�n�=0�:>�Lƾǻ��y�E���i�(?@�?脒���*��'>�t"?V��>�>���?�Ι>u/ľ;�,��?�F^?d�I?FFA?3�>�=����N�Ƚ*�%�z\/=9g�>u�X>	'i=g��=).��jY����Z�==�ѹ=I�Լ1����l<+԰�[$B<LM�<�"5>� 迵;H�|����
�����z�����B���r���'�)�žg���<E�����"Nk�m�x�xx���1��3���[�?~$�?燫�����-%���er����3�>$5�F�"������t������aO׾����aJ��C`�b�O�O�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >{C�<-����뾭����ο@�����^?���>��/��n��>ܥ�>�X>�Hq>����螾d1�<��?7�-?��>Ŏr�1�ɿb����¤<���?0�@�yA?��(��쾓�U=��> �	?s�?>�H1��O�+���Q�>g7�?]��?#JM=��W��	�a|e?��<o�F���߻�&�=*'�=h�=���J>,]�>����.A���ܽ\�4>�څ>�"�.����^��J�<2~]>^�սpQ��"��?��a��m�� �y���#w�=
�I?<^?�U½�d? �q�u�Ϳ����ܚc?�m�?�)�?��G?����^!�>fH۾�76?݋[?"�>9���q���=��t>¤��<U��^J�A�<A�>�f�>������A��S+U<t������ƿ��$�6|��u=#�ٺͭ[�g������wU�q,���lo�l�轜�h=ϕ�=ÇQ>|f�>W>�Z>�dW?�k?CK�>j�>�a佁����ξ�z�t?�����K�������棾HP�"�߾E�	�������3�ɾ_,=����=X.R����A� �L�b�~�F���.?�w$>�ʾd�M�.�,<�cʾ乪��i�������1̾A�1�e%n��̟?��A?8��� W�� �])�㘹�ĮW?�����ା�g�=.U���=r�>��=h���3��lS��i0?S?�y���o��.@*>�� �e0=(�+?�?93T<��>E:%?�+�(S��Z[>2�3>�֣>��>�	>R��V5۽z�?'�T?�4���Ȑ>mp��M�z��a=�	>.5�t=�'�[>L��<쌾n5W�n���l{�<�(W?Q��>��)��da�����Y==��x?��?.�>b{k?��B?\դ<%h��t�S���bw=��W?*i?a�>����	о����P�5?�e?��N>	ch����L�.�MU��$?�n?_?̀��&w}�}��z���n6?�{?T!k�&몿-�'��䪾 ?���>h��>�>�0I�>�c?~hx��@���g����9��#�?~9@`O�?{͎=,�=\u8����>��>��c�7����|ս!Ծ'S\=V:?B�2��(�/���N�g�N?�W�?���>'������E�=�Oq����?�L�?$��9�»g�U;g�Evݾ!k{�h��<��U�2p�����3�I���x������0M�vD}>�@�ƽ�?��o�'��_�ȿq�������ΰ��(?Y��>�-׽�ء��kl�r����.G�f?H��MY��M�>��>5���������{�0q;�����>N�	�>	�S��&��Κ��2�5<W�>���>M��>]*���轾�ę?c���?ο[������c�X?3h�?�n�?tq?�f9<c�v��{����-G?c�s?'Z?op%�E>]��7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�^�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*�+�+��<A?�2>���I�!�C0=�UҒ�ü
?W~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�3N�����Xe����@y����?N^�?i�?ӵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Pj?���� ����U>	�}?n�>��?���=M��>���=��Z"/� A#> 7�=�>�Ѡ?بM?FX�>��=$�8�D%/��\F��HR�!���C���>��a?|vL?	Fb>K��jV2�_� �xͽOv1�]1�W@���+���޽�\5>>�=>��>*�D���Ҿ�?k���%ٿ�������k8?D�l>i?�s߾&4���-�=$QY?�j�>��f���5����� �?���?�?�b�U½���=�;�>��>�ni<`Z�V{Ҿl�>t�0?�L)�eY��'d\�Y�a>�n�?vK@凴?�z�k�?��p��Y��9]�7����>h�2?�k��|�$>+�?��=��c�����Q]y�O2�>cݰ?t�?c�>�Kb?o�l�g�6�q2=�<�>��f?�
?~B񽎅
��g>���>^�&�(m�����_V?7@G�@֏W?�§��=Կ����������-�>-��=?U[>B�����=w��������=];N>!ҧ>��{>`>^>&(?>_8G>9�	>l҄��+*��Ϡ�7���f,=��"�i��w�Z���l��n�r������l��|񽚑Ͻ$�a��,�g�d�EJ=9�L?Kj_?lv?6�(?�w߽fTW>|�Ⱦ��=���1�x=~y�>�XY?Ȳz?WVD?eā�o�Ѿ0�Q�G�f�����SK`����>j�=�@�>���>���>n��<�c�>T>>kX�=�4=>� �=�ء��>ۼr>�>��>l�a>�C<>��>Fϴ��1��j�h��
w�m̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?%���z)��+���>}�0?�cW?�>���T�1:>9����j�5`>�+ �}l���)��%Q>wl?g�?>�W>��$��:���9���}����>��)?%���Y���{���K�J�-�(>��>Z=�s�te���~�ŷc�-Ñ=p�8?(^?"��Խ�MZ������_x>k�^>�!;7ſ=��?>}6��r����@��$k;噤<�Y�>�N?V�+>�Ԏ=��>kB��	�O����>�B>~�+>��??�%?�?��䗽-���)�-��w>zE�>$�>@�>=tJ��*�=}S�>��a>O��/y��)��}�?�$�W>N�|_�W�t��lx=8`�����=^�=� �0=��w%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>?N��^���щ�p*��� u=��>�TW?j����?���ל�\�?>�?{� ��y���#��Q:{��_�>T[�?>��?~eh�����=A��i�>:��?vi?���>�� �Q/��X~�>sK?00?)��>(e�m��MX(?�D�?�v�?ń>��?�)Y?0�?�0P�=�T�ok�����e~8>s?�$?��>:���6Z�}n��ǽ����H�&iE�X��>��6<'�>�O��ֵ?�	�<>b2h������v�לe>�ω>�W>�j�>v��>AZ�>J�>�-W�]����D�;-���K?���?)���2n�CO�<W��=�^��&?�I4?*k[�{�Ͼ�ը>�\?l?�[?d�>=��O>��F迿5~��s��<��K>)4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��)S��GB�>�e!?���>�Ү=�� ?��#?�j>2)�>aE��9��P�E����>��>I?��~?��?�Թ�}Z3�����桿��[�|9N>q�x?�U?�ʕ>)��������jE��GI�����!��?Ttg?�P�]?82�?��??"�A?w(f>���ؾ�����>O ?P��&�@�� '��K
���	?�?\��>#ɒ������v�C����d?��Z?�(&?@�+�_�EIƾ=(�<�� �����:<����{>�>�𐽰K�=��>�z�=�lm���9��d�<��=��>s��=ӧ:�����h.? ��y��I�=S0n�j�>��v�>n�>	$����^?[׀�����ɫ���k��9ҍ?t��?�r�?R�ͽf�Ew2?!��?��?�\
?����[?ﾠu�Ad��'-l����u�>Ӈ�>�|�����\����������r��Q)�>WC�>r9�>�	?��>�>U�j��1�UE��� ���]����O6�(�#�eg ���*���^:���;�+��Nj>���B�>Ym?{A�>�/>Ì?s����>:�5>Y�>�c�>�wB>~�3>��=��)��Ľ�KR?�����'��������3B?�qd?E1�>xi�>������0�?y��?s�?�<v>�~h��,+�_n?�=�>u��[q
?FR:=�H�=�<�U�����4��H
�5��>�F׽� :��M�nf�Jj
?�/?���ċ̾�;׽����,�=��?ø(?�(��|Q��l�r�W�PI�?L���d�Yt���#�~ l�M̎�E���9��p�*�]=(?���?�� ��d⾟ڮ��k�>�?���V>��>�Χ>rX�>�l>d���1�A,^��Z*�|���D�>}{?hό>�lI?(;<?�P?��L?t�>��>ƪ��Y��>*�;��>���>\�9?�C.?n0?4�?v�*?��a>���������ؾ=�?��?�n?e�??t?b5�������o����g�A�w�"䁽e=�=�@�<C�Խ�tq��)X=Z;R>oX?���`�8�D����k>��7?���>s��>����.����<�>_�
?CF�>  �V}r��b�hV�>���?� ���=��)>Q��=�����*Ӻ�X�=.���z�=�@��ɂ;��\<6�=Y��=�'t��s~�V�:Fk�;z�<�s�>_�? ��>nD�>�@��?� �	���a�=Y>vS>�>2Eپ�}��Y$��L�g�@\y>w�?z�?'�f=j�=b��=}|��zS������������<�?J#?�XT?���?Q�=?�i#?�>8+�wM��}^��0���?k!,?n��>P��E�ʾ�񨿜�3�ܝ?�[?�<a�n��<)���¾  ս��>�Z/�z.~�M���D���������}��(��?ӿ�?A��6�iy辸���X\����C?�"�>bY�>O�>t�)���g��%��/;>ʉ�>�R?	��>e�P?Y�z?�-]?G_Z>��<�f����{������i&>Bu??�K�?��?Hx?�g�>�n>�c2�
�㾵���
�)�s �C�~�^^^=P�^>х�>���>1x�>���=&��~���m_D����=9/p>���>Or�>���>0�{>�@�<��G?���>�\������줾cŃ���<�Ȟu?��?��+?�-=�����E��C��/M�>.o�?J��?�4*?5�S����=�ּoܶ���q�o*�>sܹ>P.�>~��=gF=�`>��>Ġ�><�>b��r8�kM�/�?	F?���=��ſxRq�<,p�����Q�z<2���v'c��ѓ��nZ����=�s���/��?��GW\�-h�������W��;Q����}�J�>ro�=�_�=hc�=t��<��μ�y�<�D=&�<�=2�u�vQl<8�;�|���	���M/�:S<bjA=^̻|�˾�y}?�7I?e�+?��C?��y>J�>B%3����>����0?y#V>�Q��l���*;������"��J�ؾ��׾jd�YƟ�S6>&�I�ͯ>�m3>l)�=s��<8��=��r=�^�=�O��='��=Ɂ�=��=���=Ѽ>�:>	8�?�r��Ң�;=X���M�)�@?u�>Z��<����O�5?�=[���l��,B�ҽr?E�?4��?j�?l�����>Ӗ�����>Z>��$�$�m=�=Š;����>�+�=e������6��i'�?�� @��'?.܄�����{�>��#>Ѽ�=�I���6�V�/�d,!�7�(��@?7���꾗u^>!�D=�L�aʾ^=Y/F>⚆=�
�9c�h�\=��'�t�-=��~=]�t>��9>]��=<�P&'>M�;��w=@=>x,�`�������r=�<�=��=>V4>3��>?�?�a0?(Xd?�6�>�n��Ͼ'?���H�>��=�E�>P��=|rB>ʏ�>6�7?o�D?�K?�>���=	�>��>D�,� �m�m�9̧��<���?�Ά?xѸ>��Q<��A�����g>�C/Ž�v?(S1?�k?k�>�U����9Y&���.�"����b4��+=�mr��QU�a���Im�4�㽯�=�p�>���>��>9Ty>�9>��N>��>��>�6�<}p�=Aጻ���<� �����=�����<�vż×���u&�8�+�/�����;g��;.�]<{��;R$
>��>3�4>>��=s�t�U?>FH�0p�-�=s���H��TO���m�t��S�ֽ�gK>Idi>��-��=��[��>��N>���;i��?�,~?��@>�����找���=��k�2�>��<H��~�=�d�[�gZ����[��>Yߎ>$�>��l>�,�L#?��w=��Yb5�~�>�|�����*)��9q�#@������ni��kҺ�D?�F��f��=i"~?��I?^�?ݍ�> ��φؾM;0>�H����=g�*q��h����?'?���>�쾤�D�W̾~��kз>z\I���O������0�J���������>�T�о~3�^f������ƌB�
jr�c�>r�O?��?B4b�G_���WO����+ꅽ2t?$�g?�>tD?�I?�ۡ��f�$|��!T�=��n?Ӭ�?�@�? c>�n�=qO����>a?��?���?��s?h�=���>�C:�:>�v����=X�
>�p�=q��=w?B9
?U�	?��P	�i���T7^�g^�<(�=��>���>��o>���=�{e=s�=��[>3��>�&�>,�d>y�>5.�>���1��n&?���=!��>��2?�C�>��X=:!����<�e]�tB��.�[���(�߽��<�MH���N=����>C�ƿ��?b�Y>����?Gv����?���V>�T>~���W�>NKD>�w}>Xӭ>|�>�>�N�>{*>��(� >-��'#+��4���C�I����=-�����"��2���;���@��Jv�b�(��d::��5=��?�K�������=C��ʭ���?�|�>K�i?>����͜>���>b=�>|d��돿Knl��	޾���?�@�3c>6�>g�W?S�?O�1�3�oZ� �u��&A��e�+�`�+፿l��� �
�`����_??�x?�vA?ל�<�/z>.��?m�%��Ώ��#�>�/��#;�'<=�6�>b.��m�`�b�Ӿ�þ�2��HF>�o?#�?HT?IV������>�'H?33?�	�?i?,?Rp?1�H�a6'?�7>G}?�F(?g�/??n;?�w+?�S�<Z�E��$��d�Ͻ%����]�^ �w�����	f=J� >����O�[�=����~�0>�}=0�,�s�>���=�?�;,ĸ����>Ay]?k4�>�6�>F�7?t��?8�����[!/?�D4=�����M�������%�>��j?��?�?Z?�c> �A��B��[>�Ê>"�%>$�[>��>�����D�b�=x�>V>@|�=�xL�L���L�	�\����p�<1�>-�?�2;>��i�il>���M�u���]>��R���	�qO��\?��ʗ�s��>�pP?�K%?ɱ >����̽��b��(?�H?�51?.\�?��>�4�[�C���E�R�)����>���=�	���Z���k��eC�\���#>㲰�����->�ݹ��E���`�IXy��'�P�ț��s��x��0��n���>tI�>�Ґ��>��)���4���:?���=�*���i���H0��%�=_�>%��>c�=3>?>�^��\ݾ�\>�O?�ڲ>��>��d��X��ܾ�\�>=�G?�`?H��?+�|���n�xb@���������4�?ţ>u��>U�@>ɲ=�橾�2���_�J�5�>�c�>�����G�隣���龮L"���>ɼ�>S>��?�U?��?��]?��,?8�?7Y�>q����跾W�&?$a�?I�={�ͽ��O�zf8��RF����>�)?a=����>�S?�?�K'?60R?�~?'�>X���OH@��Y�>���>a�V��񯿺�c>#�J?\��>M<Y?���?Բ=>�03�% ��ڧ��8�=_>�^2?-#?�?y�>D� ?�L��!�=?��>Le?Hԋ?&q{?X�>X?�Z>O��>�ޚ�9�><?��?ΒU?)+{?�J?�Y�>1:=x飽2�ٽʠ⻽S�;U/[����<c��;#p+�=P�U���ߊ�<;�=�L=�X�;ewT������T�<��=�O�>KFs>wM����+>8~þ��� �H>����֗�� ��R2����=̚{>��?iv�>|#/�U]�=hF�>m��>��H�&?�?լ?FP:�;`��\־��X�/��>v�E?��=��l�I<����r�Iyv=kl?m�]?��N��-��F�b?��]?�d�N=�&�þ(�b��|�j�O?��
?�H��׳>��~?��q?���>�f�+=n�L���<b��j����=m�>)K�p�d�+U�>��7?�o�>�b>��=�۾�w�1^���?2��?+��?_��?=*>��n� 3�$S���L?|�>�x8�C?,�>�ﭾ-�ʾ�7ʾ~$ݾ������䨾�?������nK��5G��Y�=|��>�?B>?6WX?,0о<�n��-D�{t���WG�ֽ�XG8��b9��A��a.�f(m������	�(���J�0c�~�C�H�?v�'?h)�p��>�<��4"��ξHo7> 2��&!��R�=������?=�e=�b�Z5)�D����?G�>���>��<?�sY���?�"�.��7����=y#>�8�>�͋>�M�>�@V;h�-��%׽w�ƾ����޽�v>O�c?��K?-Ln?��q�0�&j��0"�=65��ȧ���B>��
>?s�>]�W���{�%�&>�Z�r��=��@���	���=X52?��>���>��?N?��	�����w���0��3�<�t�>Oi?��>���>�mн�� ��$�>�Ol?=%�>ָ�>֫��0� �n|���ý��>��>�y�>e�p>Q�)���\�׊������t9��L�=�pi?�τ�ODa�Q>��R?�F�:|�'<���>z�r���"�1O�A(�l	>� ?Cr�=@�:>�)ž�U���z��ʊ�Kr+?�>?���Y�%��҈>�3$?6��>?T�>�R�?�_�>���9'�;�?��^?�ML?�{C?Tg�>��C=��½�;ýh1%���*=A)�>x\^>�av=^9�=����N����W�P=���=q���ݏ���Q�;)��L��<l&+=,:>(�ڿ_�G���Ӿ�r���߾k������Ͻ�z��h�4�X������qo���]'���H�+x\�6���RȌ�1t�t	�?�k�?'Ն�e�x�G`��X݂�_����Q�>ZXu��$������b��M��I۾�2��\`��8O�u��i��*?,*N��ѿs2��e���S�5?֖�>W�x?qݰ������/��{�=�`7>�U���1��YͿ鈾MM}?���>\[�|��VE�>Յ>47�=+T4>v�Ͻ�q������9F�>?�C?K��>�@�om���б���=XG�?8�@�IA?�*�ݔ�`(Z=�0�>@
?�~D>�`0�R���E�����>lK�?
�?��J=�W�v���~e?h_/<� F��G׻�f�=Mߡ=s�!=�C�eH>S�>x����C��[߽?�0> ׂ>n&�+�K{^�̇�<��_>��׽u����Ԅ?r}\��f���/�#S��-_>:�T?+�>�4�=��,?|5H��}ϿƬ\��)a?Y/�?G��?�(?�տ��ؚ>��ܾۋM?A6?z��>b&�%�t����=`VἙU��g��7(V���=��>P�>E�,����O�p��%��=�����v����!��ﾬ)^>�HW�]D��Z���y���,��񌾾��C��g(�=��T>u_>��H>���>�v>�w>?bk_?/<�>�Z >�4��g�Խ�ϻ���5����4���78e�P�R�$��3���8�ҭN��s�����Uv=��I�=��Q�&���j ��"c�їF�Y�-?�">]̾�M��<%<�8˾�ڪ�y���_5��);��1��!n����?��A?C�����V�,��P��)淽�W?�M��j��F��̩�=�R��n�=�W�>�P�=@�5�3�mS��*?��?����zm��}�$>����H�=�,?u�?g�M�г>7k(?��/��½K>�+�=3D�>��>	k>=����b���?	mO?�q�@P���>�Bݾ�p�-'>+*a>�J��$ٽ%�m>�1="Ň��V�:�����n�<W?#��>��)���U_����a&>=h�x?{�?���>�kk?�B?9��<�]��`�S�%:���u=:�W?8,i?��>_�����ϾU��֯5?܎e?qO>��h���3�.����?f�n?�`?�H���f}��
������`6?��v?�w^�9p�����W�V�
C�>_b�>���>e�9�@l�>��>?�#��D��f����V4�;? �@a��?T<<����=@9?&a�>�O�7@ƾ�i��삵��Xq=�>5���hhv����{M,��8?e��?���>��������">�΃�꺢?�*�?�%m�e�4=�پ��p����JD�Q˶��\�+-��1����5�y/��ݾ�˓�۵�>�p>~�@�4�����>i�˽��ֿ1׿f����e��q���?2Գ>ܑ���5���Um�G|��
[��Q�({þȯ�>��>����鑾�{��;�U��"��>p��ȓ�>�T�	y���矾�H<Od�>���>��>ܐ���l�����?����hο������šX?�Y�?�[�?
�?5�W<�w���{����3G?�is?�Z?� �K]���4��f?�8���Hz�F�Q��*P�1n>4P�>o+?����@�=���=��>�@u>��H��ZĿ޻����Κ?�e�?U��j��>�ţ?o L?�/������*A���a�l���?��=�r��qp�'��������>'�/??������w�_?Қa���p�+�-��ƽ�ݡ>ɿ0��c\�]1�����eXe�C��yBy����?^�?o�?��, #��5%?�>5����8Ǿg�<9��>�'�>�)N>1P_�8�u>��Q�:��j	>Q��?�~�?Qj?��������W>��}?��>/�?�T�=�D�>�>�=�հ��R*���#>��=0O@�v�?�M?T�>�R�=�69�o(/��XF�v:R�����C��
�>��a?&}L?�gb>�ո��0��!���̽RC1�^���;@�?�-�#߽/#5>��=>$>�D�mӾ��?��pؿ�_����'��S4?P�>?B*�Rt�"���_?�#�>��h.��;C������m�?��?Z�?@�׾݊ʼ8>�a�>�փ>`�ҽ9梽� w:>��B?���gM��:o�'.�>b��?��@��?g�h��	?�!�fO��`~���)�6���=K�7?!/�O�z>���>��=�lv�Z�����s����>;B�?E{�?���>��l?��o�
�B���1=�N�>�k?�s?O�o�M󾤮B>O�?��������K�tf?��
@Vu@�^?P��8˿ѓ��ѹ��py���{>:?�Y_>l�:=l��=��<a5��zB�=!����>���>���>5�>���>��>�q��S��9���x�@2�W�1�z��k���S�-��3d�](/�W�d�x>���2�nU���"=�v7���S��	ͽiH�=�zV?�R?/On?���>f�}���>ˢ �X��<������=3+�>�4/?��K?��*?p��=DB��Gc�����L����Ѕ���>��E>�d�>>c�>���>4��;�'H>
 >>yv�>Ĺ>��>=;H"=3T>�c�>��>+7�>+�;>#�>������X�h�!�w��[̽��?�C��ÌJ�'���h��0���ʖ�=�t.?��>���Hпﭿ7.H?����A)���+��M>�0?`W?�E>ġ���8Q�.�>�]�tj��V >�� ��4l��W)�I7Q>ˌ?�->��}>��&��2��+]��PѾ�[>e�)?n����l�/q�>�I�M�վ��>���>1��<|��{	��R��j2�J>�=��&?�"�>�-
�J���$�6�;���q�>=��>��<n��=L�i>>[�P"�#l)��=���=�9�>��?�L&>�K�=!^�>%S����9�/^�>�9>�0>[B?׭+?k0���𸽎fu��.7���]>(�>�<�>��>�RE��n�=�)�>�T`>��B��\|����6��LL>5VT�x�P� R��ۉ=����~p>���=w_ҽ�+�rA=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�[�>(�v[��������(>ea�>�h;?Z���[{��j�:�>? ?e���`��$Yſe���|͹>���?7&�?�#i�B����C�"5�>>�?(9/?��>�������&�>&�??U@S?5x�>��sd�g��>���?b`�?/D�>^=�?¶n?�:�>���<� �&t��r���tX�����=�a>�N���[�%m/�����	{c��(<�����1��S=��>�b8�����,Խ#���M���6��Id|>�m>�M�>F&�>�=�>��>���>w�\=U�=��о��K?��?7���n�_8�<�=�^���?�64?԰S���Ͼ<�>��\?�ˀ?�[?��>|��=��鿿&u�����<UsK>@M�>��>͎���7K>��Ծ��C�b[�>ԧ�>q��yھ�����!X�>x!?CX�>���=�� ?j�#?��j>s�>�]E��4����E�!��>���>�C?P�~?Y�?չ��U3�
��#衿��[�AN>��x?�S?�ŕ>�����E�jI�+֒�ޔ�?2og?��佡?�-�?"|??�A?�-f>~����׾�}��x�>��!?�����A�C&�e���?�k?t��>I���hս��ϼ���S���h?q�[?�&?�����`�Y�¾���<�&�a�V�*C<�PI���>��>u5���!�=�>���=�em�g6�}�g<3W�=���>��=��6�/W���<,? PH�Z؃�>��=k�r��uD�t�>vIL>4��\�^?�n=���{����x���U�� �?���?�j�?����h�(=?��?7	?�"�>M���޾0��ZRw���x�=y�X�>}��>D�l�D徲���Ι���F����Ž� �� ?4��>!?��>"�F>���>7ĥ���&���5��Y�Z���6�4�w�,�h���ş�(-"�!�c�Oʾ��cn����>V���F�>�+
?{3m>�z�>���>�G���>3k>d2}>B!�>=�h>�}@>.~�=#�<�i�o�G?��b!"��H쾍���TA?;�g?R-?G�R�K#������?&?��?��?��>>q��,�a<?� ?qZu���?���<���;? =�.���=���J�<�$<�,�>�N<h�4��*]�	0�N�?�%? 3N�5���_潝���w,o=v?�?�(?��)�P�Q��o���W��S��m��sh��j����$���p��ޏ�BO���!��Ѫ(��(=ҁ*?��?�x�[���'k��?�A�e>���>d�>\Ծ>�II>b�	�#�1��]�>9'�vă����>K{?���>#�L?H'J?4�R?�2d?[��>�b[>��f�{x?�n�=3� ?��"?SC*?n�&?�
B?<�%?=�A?+��>��3�����ξN��>�?K7?���>��?��X���Ǽ�3���^��e����N=�)�Ʉ��ػć>�*�>��?9߽�],�*���L>P~<?��?�|�>1�0��
�����=$x�>:��>���>���J�}�F�
�d��>@\x?M�L�	n��o�>}�=�`��r=�E^>��ؽP�>#��=/>5{�:�w%�%q�=6=_=D26='�=c7�=�f��<u�>��?���>kD�>*?��� �5��V�=.Y>5S>�>(Gپ~��O$��I�g�C\y>Fw�?(z�?}�f=��=A��=�{���V������������<4�?�I#?�WT?"��?��=?ii#?��>�)��L��z^�����<�?L4,?��>���̾�稿�2���?��?CF`��2��.)�������н�?>9�/�0z~��
����C�zjC7а��X��r��?�ޝ?E|@�!7���羫]��â��C?ڈ�>v�>aL�>�)���g���.�;>��>��Q?+8�>f�^?�(w?<�D?��>T5�m��-��tWz��|�>�r;?П�?�N�?���? ��>:�w>%�h�4����e���>��$)��D�����=��>��)>YM�>�f�>�!{>&?��f�ܽ;T��Q=>��>ir?�l�>rM	?5;�=���<�H?��>����&9������g��ln@�]nu?{��?f�+?N0=���g�E��w�����>�p�?Z�?�*?�fT�D��=��Ӽ6���վq�{�>�%�>�6�>�j�=,L= O>�w�>\��>���L�3<8��3N�V?F?/��=��ſj0o��(n����iU�<Xљ�� n�'����d��YU=�����4��v����d��~���������n������M��>
�=�� >Z��=VV9��QI�M�<�=Jq�;;��<Ȩh�=%�;�*+�ۼ����y��~���;͋<�(BȾ�(~?�J?ho*?-B?d�w>�7>�3]����>�y� �?�<T>�m��ӻ���8��Q�� ���	ؾm>ھ�b�*:��EF
>�AO��n
>p'5>���=&��<���=��s=���=%sr;+^/=�%�=X�=0�=���=�,>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?��>>�2������yb��-?���?�T�?>�??ti��d�>L���㎽�q�=E����=2>u��=w�2�R��>��J>���K��B����4�?��@��??�ዿТϿ6a/>r�6>�h>ӈR�Wr1���]�΂c��HZ�1r!?��:�i ̾+ȅ>Z��=!�޾ �ž�p1=O�6>��_=�� K\�D�=��x���9=�Gj=fW�>pD>��=>0��r߸=f<O=���=mP>Y#���=�e0��f4=���=��b>�'>�V?�?K�9?.|p?0��>�	���ܾ�����]>�o>J��>Ooh>)+'>�1�>��L?V�Q?M�P?7ݝ>i&#�n̾>��>f:
��c���=��_�y�_�F�?�e?��><�`>��W=����''�`$Q=Vb?��?��?u<G>Ty�*pܿ=�-�����0m=T3�H�.<�Ø���Q��3�g����Zx>8��>7��>|�>E�>�Qu>3�&>S��> C�=6��9Z��<Wvb�8o>f����<�H�;X���ui=�+Ž%�=\0ѼXف=,�Խ�i)�[��=V}�=V��=<��>�7>���>(�=�����H/>���$�L�.q�=
N��4&B�$)d�uE~��/�%h6���B>c5X>�a��3��@�?d�Y>Bu?>H��?y>u?
 >/�T�վ�Q���9e��@S�N��=i�>��<��u;�`T`�S�M���Ҿ�w�>ɯ�>x�I>�Y�=�0�����=�<��K���F�l�l>?���+v=F��=1 d����p�����f�)�=F�Y?�҄�?�=|�?�u[?ZY�?"�>�6s>�C��5>��� ����ݾ��C�<I>��?{�&?2?�p���b��E̾���o۷>�CI�T�O�B���ޫ0��Y�Ƿ�2��>����о$3�f������Y�B��Rr�@��>��O?"�?R:b�1W���RO������=r?�ug?D�>YP?`E?�3��|��n��5�=�n?���?�<�?�>��=J������>�M ?v�?x�?F'}?�<�?�>�L=��t>떜���=�a>~o=�i=q�?+�?\_
?D���������~�о��Z���<(�=��l>�Y>��>
Y>���}m=��W>S��>�&�>���><ާ>�F�>~�W�ݶ4���"?�r�=��=5.M?��?���=	:�: �>C�>��v夽�h��½���J?s=�ϊ>�fI=���>!�п�\�?��>X ¾�?����)�	<g��=��3=L���tC�-?�>��=��>QU?)=�>��t>UM�=�j��>j4���6�oyw�d;>�����O��=�1��C=��!��j��!�; ��k�q�D��|�Xo�iPa=�u�?�����2����n�����\�M?77R>�\ ?����[��E=G��>��>I<����l�������?��?�c>,F�>��W?`�?Q�0��#3��SZ���u��A���d�~�`��荿U���H�
�{i��Б_?��x?�8A?�G�<h)z>^��?��%�������>� /�}G;��7=5Q�>t����%`��6Ӿ�ľJ��$F>�>o?J��?1?�W�0��<�@>��D?��C?4�j?�p'?R�A?�<���$?��p>�U�>��?799?^>?�v
?�V>W�e>�#�����泂�4f��>��x�����~���2Rp���q=���;;�"=�20;�m�;��;�w�/T׼�B�<�x�=�+>i��=��>M^?=�>�&�>n}<?��	�@9�I����;4?Rr�=�D��6\�������eZ'>�%m?�|�?�dW?_F>��<��<�T/>��>FC8>��j>���>D��K$�2�t=>*�%>	j�=��x�����J	�~T��{Z*=�4)>a��>_ {>܆����(>v#���ky��f>��Q�b��f�T�R�G�0/2���u�_��>��K?��?�_�=����N���f��)?�<?�2M?��?���=0qܾP;:�0�J��4��V�>���<j;	������"����:�,����2r>[Q��q쥾��e>����\ܾ)�m��"K��)���<Ay���$=m���pݾ2���p~�=m��=Gp¾��"��㖿1�����H?�=辝�SgW��#���F>S�>ߞ�>.->����>�=�8�� ԃ=©�>Hp.>��F�S�D�J�ֿ�O��>��c?�	k?;hY?���=]{�o5�n*�uE��k�<�?Xf�>G�>ȁ>�)�="���Q�_�z��<P�"��>��>0�Ӿ�K�����iھ�l��
D>o^�> �+>��5?��C?T>�>�XQ?ɴ+?v?�Ss>�ۇ��ľ�N&?�	�?���= hŽ�Q���7��&F�\��>��*?��<�D�>%*?�R?k�&?��Q?�h?��>w� �s'A�V��>�>�7W��\���L^>b�I?���>yZ?#}�?��;>k�4�$���ڲ�d��=�E>�P3?|h$?ޏ?��>_0?��w�W�����>)��?���?��?՛?c�?��3�ܞ?ځ>�2�=ϱC?�xG?��c?l�?\?���=�=�;����x� ��6K�릢��{�<�k=����=��<ލ��cqr=U ���=���P����z>�<,_�>:�s>	���0>�ľ�O����@>Ԙ��%P��eي��:�Eݷ=��>+�?p��>qY#�E��=3��>oH�>����6(?�?w?V�!;͡b�,�ھ��K���>B?��=&�l�h�����u�ch=��m?�^?.�W�"'��N�b?��]?:h��=�	�þ��b����c�O?:�
?.�G���>��~?c�q?O��>�e�(:n�)��Db���j�)Ѷ=^r�>HX�S�d�?�>m�7?�N�>*�b>%�=eu۾�w��q��e?��?�?���?+*>��n�X4�b	��_kM?H��>�#���1?���<��꾵^��&����羠S���@��s���6r}���`���M���ܽc�=�i?�N|?�kO?UN_?�H���q�a";�GEn��NQ���9�&E@��y9���R��}C��s�f+ž�����lﾟ����`��#W�9n�?�'?�tE�9��>e�b�.뾾ž�п>�J���+�2�>�������=c�<A0�x�Ʀ����?��>��>��L?�J�R,Q�!���?���=�>\!}>�*>Hb�>�4���D�$Y� C��u�ľ��ƽ�/�>}�v?\�`?�jA?h�K�˘2����h80���<���l�>Ɉ��J>W��Ϥ�>���4���u���������3�������5?�.�>�>yN�?wj?���Wl�������#��xV>��?��G??��>�Ǘ>3-E=������>9�l?E��>���>Y���KX!�~�{��lʽ"�>1�>=��>��o>)�,�c(\��i�������9���=ïh?T�����`���>
R?�]�:��F<҆�>^ w���!����8�'�7�>�w?ڪ=�;>�ž���{�!B���)?�$?3����(�=�>�~"?R��>�ަ>q�??��>Wk���;�?�S_?�lJ?��A?�_�>n:=�F����Ľ��%���,=��>]�[>hDf=vN�=T����^��j�`�I=�-�=Sx��_O��*<F<�4����M<!��<�44>�cؿR�E���ϾGM
�o��d9���������)�����y۸��K���g����R�[�e�\��k��w����o��U�?���?2��Iv��)F�� 4��y>��R*�>�"s�ʫ��������H	����ݾ�&���� �hS�	�k��Qf��'?������ǿ�����@ܾ�" ?�4 ?ԫy?��w�"�T�8�a� >6��<����Ф뾯�����οU���j�^?���>��B��M��>o��>��X>&q>k����螾$,�<s�??�-?ݝ�>��r��ɿ懻����<���?��@�yA?9�(�\��lV=��>	?��?>�X1��F�)˰��K�>s8�?���?I`M=.�W��	�\e?g�<��F��ܻ��=�Q�=�=����VJ>@X�>z���uA�)[ܽK�4>.҅>O�"���Pn^��s�<x�]>�Eֽ	9��5Մ?,{\��f���/��T��U>��T? +�>U:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=m6�މ��{���&V����=[��>c�>,�ߋ���O��I��U��=���1�˿� ���ʑ��y��U%�B8㽽۽l�6=��n������`���a�<Plf;��=_>�C>�\	>�I?{�Q?t&�> �4>�p̽E�T�c[澮�Q�#넾��<��G��<�x����I꾲=Ӿ!�+���>��� �����$=���=�*R������� �:�b���F�N�.?�M$>��ʾ5�M�GT*<��ʾ�ê�;������:̾��1�=n�{ʟ?��A?�h�V�m���mp���W?$M�w��Cꬾ���=BC��E�=O�>���=���`,3��wS�8w0?�X?s����X��2*>�� ��=��+?\�?sZ<V+�>�L%?k�*�a�{m[>�3>gݣ>���>�5	>/��FO۽�?��T?������ؐ>�f����z�7#a=H+>g,5��鼜�[>䞒<����QV�"U��=��<�(W?q��>��)��wa��G��MY==��x?��?.�>m{k?��B?�դ<h��{�S����aw=�W?2*i?��>����	о]���D�5?�e?~�N>�bh���;�.�\U��$?�n?1_?X~��%w}����k���n6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?w�;<��T��=�;?m\�> �O��>ƾ�z������-�q=�"�>���ev����R,�f�8?ݠ�?���>�������q>�L{�o*�?�Z�?`+[���ٽ�4澔�c�����Uoͼ(�7���;��)���L�~��Cᾥ䷾���k>6�@Z��<HO�<�����ۿ�Zο�=������;��)$?��E>77�����uz���N��i����\��x���N�>�>{~������R�{��t;�+F��I�>C��
�>E�S��%��+����5<��>"��>v��>�k���?�Z���:ο����c���X?�e�?�k�?�l?K�9<�v�{�����,G?l�s?�Z?�u%��R]��7���a?S�W�=���h�e��wG��0>�Z�>��?[��q��=ǭY��?�k>�-[�T��	���{
�*,�?� �?%���l�>Ω�?*�S?��������ؽ܊=��{[�jG-?K�>��%!�e�쾝U��)��>��F?��>��7�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�&�>Y�?�.�=<�>�k�=�����-���">��=��>���?��M?�.�>�4�=��8��/��TF�\R��.�G�C���>��a?tL?J�a>����92�0!���ͽiE1��弃H@��-�nF߽�Z5>l�=> >E��Ӿu@?�澗r�;�����g�OJ9?tյ�ȶ5?R�uof�3т��?я�>��I��T��������� ��?�}@���>�z�����=�>���>ar�=��߽��������t>�\)?�����҈���P�C0�>���?���?�?��V��	?���P��Ua~����7�l��=��7?�0��z>���>��=�nv�ݻ��X�s����>�B�?�{�?��> �l?��o�O�B���1=;M�>͜k?�s?kQo���h�B>��?!������L��f?�
@u@`�^?*�kؿ쌢���ɾ�4ž2ެ<4'�;%�->>}���8����9�'=b�<y��<�A�>0�M>o>�Bd>W:h>�_�=����w�2w�����ϙB��=.�nS�����9�ɾ^���W�0��Dվ���1������
`�gh��k���e�%2>>�5?�]?]�q?��>����"�="�,��������\>)�H>� ;?�KR?e�/?�=0>u#��T�����Y�r��킾3��>��>{��>��>҂�>)P���2>��z>+�>���>�*4>��F���>4h>q��>�S�>�MC>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?�f>�8u>��3�qd8���P�솰�Z|>�'6?ﶾ>9�}�u���H�kݾ�:M>���>��C�m��������ki� �{=7w:?��?�S���ް��u��@��5HR>*:\>��=�_�=SKM>O8c�Y�ƽ�H��[.=Q��=ת^>�8?�,>���=f��>�J��N�P�֜�>��>>D}+>�??Rg%?Q������⁾+�+�Nx>��>
H~>�>�{I���=��>@�c>� �6~���z��o?�GGX>�~���`�g�u��y=����4H�=8�=�&��2�<��=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾN�>�Mɼ�Z��Ş���y���q=Q��=�T?��u�'�齻�ھ�t?�)?d�9�������˿��?3�>�u�?5��?:�J��3���r�&m�>"��?�� ?N�?`��,��컢>-�p?�u?� m>;��!l����>�}�?�L�?�j>���?gu�?ٸ�>����n8��b��������U�!�O=,��>��=�w޾$�1��P|��?\��k^��rE�!��=�\(=���>�҆�?���E8�=��M<A;��f	;��`�>�A>�O�>��S>�'�>  �>'A�>H���;*��LB��!w���K?O��?���i1n��F�<�z�=!�^��?�B4?k[�D�Ͼ(Ѩ>N�\?׿�?[?�h�>���)@��*翿�z��<b�K>j2�>�A�>����9K>��Ծ�3D� o�>)ٗ>	��J@ھ!���W��*<�>Qd!?<��>Ӯ=O� ?��#?�zj>��>�aE��9����E�\��>���>�H?��~?��?�͹�A`3��
���桿ە[��4N>�x?fZ?�Ǖ>���v����QF��`H�;��V��?Uvg?B|彖?V5�?Ӓ??!�A?�0f>3��cؾ~����>��!?,f�=�A�WI&�2���a?PC?ۑ�>S���!�սM�Ѽ��� ���C�?.\?H&?ْ�Q?a��þn�<��"��O�W� <
�F�d�>�M>u���i{�=��>8��=�0m�W`6��\l<z�=�Z�>���=�7�sD��0=,?�G�}ۃ���=��r�>xD���>�IL>����^?ll=��{�����x��	U� �? ��?Zk�?_��@�h��$=?�?S	?n"�>�J���}޾6���Pw�~x��w�Z�>���>D�l���J���ڙ���F��b�Ž<�6�
� ?�I�>���>2%�>b��>(�>����H~��A�����H����v�2�?�=���+�����]�a*}�YZʾ�l��&�>@\<��>	?f��>a�[>��?���H�>#5z>��5>�2�>���>�{�>%i>��0���&��KR?���� �'���込���g3B?�qd?Q1�>hi�8��������?���?Qs�?"=v>h��,+��n?�>�>E��Tq
?�T:=�7�m;�<V��r��/3���+��>E׽� :��M�@nf�wj
?�/?�����̾�;׽�I��!�=Sat?��>ns?�tЏ��P��}W���k��+��\���@�	�z��Nq�����y�i����hl�8�^<�!??`?l
Ⱦ����d���AO��	���@>	U�>�?�>�c�=�@>���+fU��I9�:dƾa�Ͼ��P>3oK?x�>s2?�"8?��e?7�D?��>�X�>b����;?�=���>�@ ?�k6?mq=?Q7?��.?7QA?:� >��T����G�վ�=�>�6�>��"?�?4}+?$��Y4&�����,=���?嘾o/N>E� ���&� �>���T>zw�>*Y?����8������k>��7?l��>���>P��<-��g�<��>�
?�G�>O  ��|r�b��W�>5��?j����=Q�)>���=����AXӺCV�=������=�/���{;��\<���=Z��=/Yt������:cl�;�q�< u�>6�?���>�C�>�@��/� �c��f�=�Y>=S>|>�Eپ�}���$��v�g��]y>�w�?�z�?ϻf=��=��=}���U�����H������<�??J#?)XT?`��?{�=?_j#?е>+�jM���^�������?O,?K��>�5�Ek˾�꨿�m3��?|�?�%a��Tc)�����4ӽ?�>�n/�[n~�V�ձC��R���������?G��?�D�C�6�ZE�HИ�d?���OC?*z�>�O�>��>G�(�wh��4��<>��>zbQ?�L�>�HK?9��?�=C?Jئ<����/��7���jk��4w>p�M?�Z?��|?@�e?	,�>�o�>S�@��������L��L.�,�R�'�>(dg>9��>�Ȏ>綽>d؛>p�轻��2}�ı�=恊>���>^M>ʴ?�G�>]�<y�G?���>[����%餾MÃ�=�m�u?���?��+?ef=��^�E�B���L�>[o�?���?o2*?��S�*��=��ּ�ⶾK�q��$�>�۹>�6�>xؓ=�F=�]>s�>Ğ�>m1��^��p8�"EM��?�F?z��=�̿����CJ��x��},��Q���㘾��
���N>���g�j���о'la��h�����ro־,9����i����>�Q>�I>���=OȻ��������]��Ѵ�7�e�n����<�|���a��>ɽA�νo� �Ͱ�'�>�P�˾�}?�<I?*�+?޾C?6�y>v7>��3���>����A?�V>U�P�p����;�6���� ����ؾz׾H�c��ɟ��H>�UI���>�;3>:>�=!I�<��=ds=�ˎ=�jR��=~.�=Q�=�`�=s��=�>�T>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�7>�M>�R���1���\��b�j}Z��!?�I;��@̾�F�>���=�0߾q�ƾ��.=Ǚ6>N8b=O��W\���=e�z�:�;=� l=�ԉ> �C>�I�=p2����=ўI=_��=�O><���>P7��,�f3=���=��b>�&>�E�>*=?Қ5?!mk?��>�[�Dc߾<�Ͼ�7�>�>젱>Y>a�>��>� >?�J?eS?95�>d�'�ʕ�>���>Cj'���Z��ؾ_����=]��?'�?�E�>6Dݻ�P4�I|"�6�'�	xͽ�o?4B?W!?U�>!���'⿎�&�bN+�V׽o��<$I�[P?�۳���
!�O���9�<ZD�>�ʪ>�|�>��j>�b/>�,3>��><:>F�L=8�=�2�"Ϩ������sY=*LG=ه�=�|ϼpG���~ɼ �����o�8�W���������6��c��=���>�@>��>���=� ��EH/>*���[�L���=LI��3+B�d1d�#H~�{	/�\h6�M�B>NAX>�s���3����?��Y>-t?>u��?wAu?K�>&��վ�Q���7e��QS�z��=��>U�<�t;�cT`���M�j�Ҿ>W�>�z�>&�]>�Y=i4�fk�e�<����^�n��Xj>��ľ�΄�:���r��-�������VS�c�>c�W?(Y���$�=KV�?�c?Bz�?R�?��>ܥ ���>76��3!>��&�EΜ���>� �>q&?��?�"����#�̾$�����>Q}I���O����n�0�;�=�������>ַ���fҾ�!3�峆�Qj��w�B���w�X5�>OoO?��?ta����INP��l�gt��u?Յh?ڵ�>�?~>?LG����辞���F�=�5m?�]�?�`�?��>��"=�;�(��>���>�ؖ?���? yp?�6�er?�.,�v'>��e�4�=���=�=�=��?��?/� ?�aZ�����m��{���!�^ƭ=r�<���>�:�>;1�>��S>�*�=�=�=F��>y�?�}�>�_>닑>��>��������(?��=F��>��N?��>�/�=�7�=��7>��a����GN�;�Ž�<׼�0;>��<p�a>v�=�h�>�׿��?ރ�>�3����>�˺���彠=K�?h38��M�>�>�H>#s?��g>t�R>�x4>/�M>O�־�A>�����
�>��Qk��N����4>�����n	���:�p'b��Vh�i��m�1�33k����	^5��P�=1(�?�gڽ(���)�T�F,�o%1?Mo>��`?m���Lܽ�v�=��"?|��>���h��Ϝ���X��_ϒ?_��?�;c>��>^�W?Ś?Ǔ1�L3��uZ�I�u�X(A��e�ܻ`�k፿����ٗ
������_?��x?txA?�H�<:z>K��?d�%��ӏ�!)�>�/�';��=<=0+�>�)����`���Ӿ`�þ�6��HF>F�o?�$�?�X?UV�J� �˲(>m><?�6?�Jm?*�*?�V4?HU;���?��H>�?;�?6(7?%�0?��?�:?>�&>�	����W�Lh������R�ý�����
� �t=� *=���}O�;@�1=@�<��;E�:�eP�u����<&�X=T�=�o�=Ȧ>՜]?U�>Զ�>��7?h��o8�Yɮ�X?/?�u:=敂��􊾊���g��)>��j?���?tPZ?hd>��A��C���>�U�>?�&>+;\>
��>x���|E�,��=5P>�0>W�=[L�2с��	��������<g>K��>K"|>�卽�'>�z���3z�$�d>�R��к���S���G���1��v��R�>G�K?��?���=�e��2��HDf�p6)?+W<?�IM?��?Փ=�۾F�9���J��g�o�>O�<R��𼢿�#��R�:��(�:�s>16������->�ݹ��E���`�IXy��'�P�ț��s��x��0��n���>tI�>�Ґ��>��)���4���:?���=�*���i���H0��%�=_�>%��>c�=3>?>�^��\ݾ�\>�O?�ڲ>��>��d��X��ܾ�\�>=�G?�`?H��?+�|���n�xb@���������4�?ţ>u��>U�@>ɲ=�橾�2���_�J�5�>�c�>�����G�隣���龮L"���>ɼ�>S>��?�U?��?��]?��,?8�?7Y�>q����跾W�&?$a�?I�={�ͽ��O�zf8��RF����>�)?a=����>�S?�?�K'?60R?�~?'�>X���OH@��Y�>���>a�V��񯿺�c>#�J?\��>M<Y?���?Բ=>�03�% ��ڧ��8�=_>�^2?-#?�?y�>D� ?�L��!�=?��>Le?Hԋ?&q{?X�>X?�Z>O��>�ޚ�9�><?��?ΒU?)+{?�J?�Y�>1:=x飽2�ٽʠ⻽S�;U/[����<c��;#p+�=P�U���ߊ�<;�=�L=�X�;ewT������T�<��=�O�>KFs>wM����+>8~þ��� �H>����֗�� ��R2����=̚{>��?iv�>|#/�U]�=hF�>m��>��H�&?�?լ?FP:�;`��\־��X�/��>v�E?��=��l�I<����r�Iyv=kl?m�]?��N��-��F�b?��]?�d�N=�&�þ(�b��|�j�O?��
?�H��׳>��~?��q?���>�f�+=n�L���<b��j����=m�>)K�p�d�+U�>��7?�o�>�b>��=�۾�w�1^���?2��?+��?_��?=*>��n� 3�$S���L?|�>�x8�C?,�>�ﭾ-�ʾ�7ʾ~$ݾ������䨾�?������nK��5G��Y�=|��>�?B>?6WX?,0о<�n��-D�{t���WG�ֽ�XG8��b9��A��a.�f(m������	�(���J�0c�~�C�H�?v�'?h)�p��>�<��4"��ξHo7> 2��&!��R�=������?=�e=�b�Z5)�D����?G�>���>��<?�sY���?�"�.��7����=y#>�8�>�͋>�M�>�@V;h�-��%׽w�ƾ����޽�v>O�c?��K?-Ln?��q�0�&j��0"�=65��ȧ���B>��
>?s�>]�W���{�%�&>�Z�r��=��@���	���=X52?��>���>��?N?��	�����w���0��3�<�t�>Oi?��>���>�mн�� ��$�>�Ol?=%�>ָ�>֫��0� �n|���ý��>��>�y�>e�p>Q�)���\�׊������t9��L�=�pi?�τ�ODa�Q>��R?�F�:|�'<���>z�r���"�1O�A(�l	>� ?Cr�=@�:>�)ž�U���z��ʊ�Kr+?�>?���Y�%��҈>�3$?6��>?T�>�R�?�_�>���9'�;�?��^?�ML?�{C?Tg�>��C=��½�;ýh1%���*=A)�>x\^>�av=^9�=����N����W�P=���=q���ݏ���Q�;)��L��<l&+=,:>(�ڿ_�G���Ӿ�r���߾k������Ͻ�z��h�4�X������qo���]'���H�+x\�6���RȌ�1t�t	�?�k�?'Ն�e�x�G`��X݂�_����Q�>ZXu��$������b��M��I۾�2��\`��8O�u��i��*?,*N��ѿs2��e���S�5?֖�>W�x?qݰ������/��{�=�`7>�U���1��YͿ鈾MM}?���>\[�|��VE�>Յ>47�=+T4>v�Ͻ�q������9F�>?�C?K��>�@�om���б���=XG�?8�@�IA?�*�ݔ�`(Z=�0�>@
?�~D>�`0�R���E�����>lK�?
�?��J=�W�v���~e?h_/<� F��G׻�f�=Mߡ=s�!=�C�eH>S�>x����C��[߽?�0> ׂ>n&�+�K{^�̇�<��_>��׽u����Ԅ?r}\��f���/�#S��-_>:�T?+�>�4�=��,?|5H��}ϿƬ\��)a?Y/�?G��?�(?�տ��ؚ>��ܾۋM?A6?z��>b&�%�t����=`VἙU��g��7(V���=��>P�>E�,����O�p��%��=�����v����!��ﾬ)^>�HW�]D��Z���y���,��񌾾��C��g(�=��T>u_>��H>���>�v>�w>?bk_?/<�>�Z >�4��g�Խ�ϻ���5����4���78e�P�R�$��3���8�ҭN��s�����Uv=��I�=��Q�&���j ��"c�їF�Y�-?�">]̾�M��<%<�8˾�ڪ�y���_5��);��1��!n����?��A?C�����V�,��P��)淽�W?�M��j��F��̩�=�R��n�=�W�>�P�=@�5�3�mS��*?��?����zm��}�$>����H�=�,?u�?g�M�г>7k(?��/��½K>�+�=3D�>��>	k>=����b���?	mO?�q�@P���>�Bݾ�p�-'>+*a>�J��$ٽ%�m>�1="Ň��V�:�����n�<W?#��>��)���U_����a&>=h�x?{�?���>�kk?�B?9��<�]��`�S�%:���u=:�W?8,i?��>_�����ϾU��֯5?܎e?qO>��h���3�.����?f�n?�`?�H���f}��
������`6?��v?�w^�9p�����W�V�
C�>_b�>���>e�9�@l�>��>?�#��D��f����V4�;? �@a��?T<<����=@9?&a�>�O�7@ƾ�i��삵��Xq=�>5���hhv����{M,��8?e��?���>��������">�΃�꺢?�*�?�%m�e�4=�پ��p����JD�Q˶��\�+-��1����5�y/��ݾ�˓�۵�>�p>~�@�4�����>i�˽��ֿ1׿f����e��q���?2Գ>ܑ���5���Um�G|��
[��Q�({þȯ�>��>����鑾�{��;�U��"��>p��ȓ�>�T�	y���矾�H<Od�>���>��>ܐ���l�����?����hο������šX?�Y�?�[�?
�?5�W<�w���{����3G?�is?�Z?� �K]���4��f?�8���Hz�F�Q��*P�1n>4P�>o+?����@�=���=��>�@u>��H��ZĿ޻����Κ?�e�?U��j��>�ţ?o L?�/������*A���a�l���?��=�r��qp�'��������>'�/??������w�_?Қa���p�+�-��ƽ�ݡ>ɿ0��c\�]1�����eXe�C��yBy����?^�?o�?��, #��5%?�>5����8Ǿg�<9��>�'�>�)N>1P_�8�u>��Q�:��j	>Q��?�~�?Qj?��������W>��}?��>/�?�T�=�D�>�>�=�հ��R*���#>��=0O@�v�?�M?T�>�R�=�69�o(/��XF�v:R�����C��
�>��a?&}L?�gb>�ո��0��!���̽RC1�^���;@�?�-�#߽/#5>��=>$>�D�mӾ��?��pؿ�_����'��S4?P�>?B*�Rt�"���_?�#�>��h.��;C������m�?��?Z�?@�׾݊ʼ8>�a�>�փ>`�ҽ9梽� w:>��B?���gM��:o�'.�>b��?��@��?g�h��	?�!�fO��`~���)�6���=K�7?!/�O�z>���>��=�lv�Z�����s����>;B�?E{�?���>��l?��o�
�B���1=�N�>�k?�s?O�o�M󾤮B>O�?��������K�tf?��
@Vu@�^?P��8˿ѓ��ѹ��py���{>:?�Y_>l�:=l��=��<a5��zB�=!����>���>���>5�>���>��>�q��S��9���x�@2�W�1�z��k���S�-��3d�](/�W�d�x>���2�nU���"=�v7���S��	ͽiH�=�zV?�R?/On?���>f�}���>ˢ �X��<������=3+�>�4/?��K?��*?p��=DB��Gc�����L����Ѕ���>��E>�d�>>c�>���>4��;�'H>
 >>yv�>Ĺ>��>=;H"=3T>�c�>��>+7�>+�;>#�>������X�h�!�w��[̽��?�C��ÌJ�'���h��0���ʖ�=�t.?��>���Hпﭿ7.H?����A)���+��M>�0?`W?�E>ġ���8Q�.�>�]�tj��V >�� ��4l��W)�I7Q>ˌ?�->��}>��&��2��+]��PѾ�[>e�)?n����l�/q�>�I�M�վ��>���>1��<|��{	��R��j2�J>�=��&?�"�>�-
�J���$�6�;���q�>=��>��<n��=L�i>>[�P"�#l)��=���=�9�>��?�L&>�K�=!^�>%S����9�/^�>�9>�0>[B?׭+?k0���𸽎fu��.7���]>(�>�<�>��>�RE��n�=�)�>�T`>��B��\|����6��LL>5VT�x�P� R��ۉ=����~p>���=w_ҽ�+�rA=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�[�>(�v[��������(>ea�>�h;?Z���[{��j�:�>? ?e���`��$Yſe���|͹>���?7&�?�#i�B����C�"5�>>�?(9/?��>�������&�>&�??U@S?5x�>��sd�g��>���?b`�?/D�>^=�?¶n?�:�>���<� �&t��r���tX�����=�a>�N���[�%m/�����	{c��(<�����1��S=��>�b8�����,Խ#���M���6��Id|>�m>�M�>F&�>�=�>��>���>w�\=U�=��о��K?��?7���n�_8�<�=�^���?�64?԰S���Ͼ<�>��\?�ˀ?�[?��>|��=��鿿&u�����<UsK>@M�>��>͎���7K>��Ծ��C�b[�>ԧ�>q��yھ�����!X�>x!?CX�>���=�� ?j�#?��j>s�>�]E��4����E�!��>���>�C?P�~?Y�?չ��U3�
��#衿��[�AN>��x?�S?�ŕ>�����E�jI�+֒�ޔ�?2og?��佡?�-�?"|??�A?�-f>~����׾�}��x�>��!?�����A�C&�e���?�k?t��>I���hս��ϼ���S���h?q�[?�&?�����`�Y�¾���<�&�a�V�*C<�PI���>��>u5���!�=�>���=�em�g6�}�g<3W�=���>��=��6�/W���<,? PH�Z؃�>��=k�r��uD�t�>vIL>4��\�^?�n=���{����x���U�� �?���?�j�?����h�(=?��?7	?�"�>M���޾0��ZRw���x�=y�X�>}��>D�l�D徲���Ι���F����Ž� �� ?4��>!?��>"�F>���>7ĥ���&���5��Y�Z���6�4�w�,�h���ş�(-"�!�c�Oʾ��cn����>V���F�>�+
?{3m>�z�>���>�G���>3k>d2}>B!�>=�h>�}@>.~�=#�<�i�o�G?��b!"��H쾍���TA?;�g?R-?G�R�K#������?&?��?��?��>>q��,�a<?� ?qZu���?���<���;? =�.���=���J�<�$<�,�>�N<h�4��*]�	0�N�?�%? 3N�5���_潝���w,o=v?�?�(?��)�P�Q��o���W��S��m��sh��j����$���p��ޏ�BO���!��Ѫ(��(=ҁ*?��?�x�[���'k��?�A�e>���>d�>\Ծ>�II>b�	�#�1��]�>9'�vă����>K{?���>#�L?H'J?4�R?�2d?[��>�b[>��f�{x?�n�=3� ?��"?SC*?n�&?�
B?<�%?=�A?+��>��3�����ξN��>�?K7?���>��?��X���Ǽ�3���^��e����N=�)�Ʉ��ػć>�*�>��?9߽�],�*���L>P~<?��?�|�>1�0��
�����=$x�>:��>���>���J�}�F�
�d��>@\x?M�L�	n��o�>}�=�`��r=�E^>��ؽP�>#��=/>5{�:�w%�%q�=6=_=D26='�=c7�=�f��<u�>��?���>kD�>*?��� �5��V�=.Y>5S>�>(Gپ~��O$��I�g�C\y>Fw�?(z�?}�f=��=A��=�{���V������������<4�?�I#?�WT?"��?��=?ii#?��>�)��L��z^�����<�?L4,?��>���̾�稿�2���?��?CF`��2��.)�������н�?>9�/�0z~��
����C�zjC7а��X��r��?�ޝ?E|@�!7���羫]��â��C?ڈ�>v�>aL�>�)���g���.�;>��>��Q?+8�>f�^?�(w?<�D?��>T5�m��-��tWz��|�>�r;?П�?�N�?���? ��>:�w>%�h�4����e���>��$)��D�����=��>��)>YM�>�f�>�!{>&?��f�ܽ;T��Q=>��>ir?�l�>rM	?5;�=���<�H?��>����&9������g��ln@�]nu?{��?f�+?N0=���g�E��w�����>�p�?Z�?�*?�fT�D��=��Ӽ6���վq�{�>�%�>�6�>�j�=,L= O>�w�>\��>���L�3<8��3N�V?F?/��=��ſj0o��(n����iU�<Xљ�� n�'����d��YU=�����4��v����d��~���������n������M��>
�=�� >Z��=VV9��QI�M�<�=Jq�;;��<Ȩh�=%�;�*+�ۼ����y��~���;͋<�(BȾ�(~?�J?ho*?-B?d�w>�7>�3]����>�y� �?�<T>�m��ӻ���8��Q�� ���	ؾm>ھ�b�*:��EF
>�AO��n
>p'5>���=&��<���=��s=���=%sr;+^/=�%�=X�=0�=���=�,>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?��>>�2������yb��-?���?�T�?>�??ti��d�>L���㎽�q�=E����=2>u��=w�2�R��>��J>���K��B����4�?��@��??�ዿТϿ6a/>r�6>�h>ӈR�Wr1���]�΂c��HZ�1r!?��:�i ̾+ȅ>Z��=!�޾ �ž�p1=O�6>��_=�� K\�D�=��x���9=�Gj=fW�>pD>��=>0��r߸=f<O=���=mP>Y#���=�e0��f4=���=��b>�'>�V?�?K�9?.|p?0��>�	���ܾ�����]>�o>J��>Ooh>)+'>�1�>��L?V�Q?M�P?7ݝ>i&#�n̾>��>f:
��c���=��_�y�_�F�?�e?��><�`>��W=����''�`$Q=Vb?��?��?u<G>Ty�*pܿ=�-�����0m=T3�H�.<�Ø���Q��3�g����Zx>8��>7��>|�>E�>�Qu>3�&>S��> C�=6��9Z��<Wvb�8o>f����<�H�;X���ui=�+Ž%�=\0ѼXف=,�Խ�i)�[��=V}�=V��=<��>�7>���>(�=�����H/>���$�L�.q�=
N��4&B�$)d�uE~��/�%h6���B>c5X>�a��3��@�?d�Y>Bu?>H��?y>u?
 >/�T�վ�Q���9e��@S�N��=i�>��<��u;�`T`�S�M���Ҿ�w�>ɯ�>x�I>�Y�=�0�����=�<��K���F�l�l>?���+v=F��=1 d����p�����f�)�=F�Y?�҄�?�=|�?�u[?ZY�?"�>�6s>�C��5>��� ����ݾ��C�<I>��?{�&?2?�p���b��E̾���o۷>�CI�T�O�B���ޫ0��Y�Ƿ�2��>����о$3�f������Y�B��Rr�@��>��O?"�?R:b�1W���RO������=r?�ug?D�>YP?`E?�3��|��n��5�=�n?���?�<�?�>��=J������>�M ?v�?x�?F'}?�<�?�>�L=��t>떜���=�a>~o=�i=q�?+�?\_
?D���������~�о��Z���<(�=��l>�Y>��>
Y>���}m=��W>S��>�&�>���><ާ>�F�>~�W�ݶ4���"?�r�=��=5.M?��?���=	:�: �>C�>��v夽�h��½���J?s=�ϊ>�fI=���>!�п�\�?��>X ¾�?����)�	<g��=��3=L���tC�-?�>��=��>QU?)=�>��t>UM�=�j��>j4���6�oyw�d;>�����O��=�1��C=��!��j��!�; ��k�q�D��|�Xo�iPa=�u�?�����2����n�����\�M?77R>�\ ?����[��E=G��>��>I<����l�������?��?�c>,F�>��W?`�?Q�0��#3��SZ���u��A���d�~�`��荿U���H�
�{i��Б_?��x?�8A?�G�<h)z>^��?��%�������>� /�}G;��7=5Q�>t����%`��6Ӿ�ľJ��$F>�>o?J��?1?�W�0��<�@>��D?��C?4�j?�p'?R�A?�<���$?��p>�U�>��?799?^>?�v
?�V>W�e>�#�����泂�4f��>��x�����~���2Rp���q=���;;�"=�20;�m�;��;�w�/T׼�B�<�x�=�+>i��=��>M^?=�>�&�>n}<?��	�@9�I����;4?Rr�=�D��6\�������eZ'>�%m?�|�?�dW?_F>��<��<�T/>��>FC8>��j>���>D��K$�2�t=>*�%>	j�=��x�����J	�~T��{Z*=�4)>a��>_ {>܆����(>v#���ky��f>��Q�b��f�T�R�G�0/2���u�_��>��K?��?�_�=����N���f��)?�<?�2M?��?���=0qܾP;:�0�J��4��V�>���<j;	������"����:�,����2r>[Q��sj����>A8辡ʾ=9q���K�ȭܾD�=�>�#����=�	����Ņ�f��=���=%﷾����LŨ�g�D?�=�����[�OC־��=���>H×>L�%��>��Q@�gc��a�=!��>�/>�����YE�R����>�SS?��i?J�q?��Ǿ�ls���-��k�b$��"==h�>z�I>���>�Z>��=���������
n�^lS�vh�>�f�>	�#1�U�þT?� �!PB>��?�x5>_��>Ɩ:?4�?b?�?8��>%�6>P/���Ͼa=&?D��?�`�=�Խh�T���8��F�m��>�)?�dB��͗>��?A�?��&?�Q?�?�>[� �
G@����>�Y�>��W�1X���A`>��J?렳>�DY?3?��=>�q5��+��G$��͟�=�G>O�2?�I#?��? ��>��7?�T�m����Qh>5z�?IŌ?[�?���>��>�X�1�k?os0=(D��9�J?��??y*l?�ړ?��??��=���=?3��.�i���n���)�����<��7=F=�۰�B�<�s�<6}^<�t=���<�#����W��=\(�;�.�>?s>+s��12>tþ�o���yE>rE��7љ����O�3�*Q�=�;�>�E?�o�>ޱ*� �=��>f�>׽��$&?�?I@?� ��aVb���ھs-M�e�>��B?~��=��l������u�M�p=3lm?E�^?MQ��,��>�b?�]?_h�=���þ�b�m��o�O?�
?1�G�i�>��~?'�q?v��>��e�U:n�+���Cb���j�(ж=4r�>�W���d�e?�>�7?RN�>��b>�$�=ju۾��w��q��D?[�?�?���?�+*>p�n�Z4��%��ލ�k+X?i$�>�䒾f�?%�R���̾E���K�ʾEW��پ���dl��c�����܎���_h=$�?�i�?�`w?u�^?|���7�u�!z��I����6�F�������YA�^�I�>\~�%3(���:�Ծ}�j;��K�iC�Ԣ�?3/?���3�>�u��,�����= D>O$��?����>Oཽ܈+=��7=�j9�`�����P�?��>L�>�L?�M�+���$���1�Y����|�=�ъ>��>�n�>��=wm,�ϯ��cθ�Mذ�F1a�$p>��a?�H?1ub?~
���.�3�1�U���蝾}&>lc�=�s�>*Z�W�0��!�_<���p��x
�Au��X�����=nA5?S-�>b��>Ӈ�?~D?����ƾ`2�!�2�)��='�>�YZ?���>ȸu>��}�!�%��>��l?�t�>�&{> ��_�$�����D�p����>�9�>��>�b�>�G/��c�R����\���N>�{>�=�u?KV��W�[�ۥ�>׾b?��;������>�ޏ�����@���h����=p/?C�=�gM>_�������.�w��ة�T�*?��?�����)�tՂ>>�!?x;�>!p�>�T�?$œ>� ��K�:_�?��_?!�J?
�B?��>�H=� ��Ƚ��%�#f<=0��>d�Z>��p=qy�=�����U����wC=j{�=^����s��m��<N����4�;4�<��2>�ڿ�I��{;�
���� �
�+Q����½;���3�&��a���W�����,s�*�دN���l�:哾�Zv�f=�?��?�|���v�����悿f<���>zn�p�`��}���$Խ�+���.�r���)��
V���m��`��'?ΐ��ǿ���'�۾w9 ?�-?�~y?}p�<"�Г8���">��<nҳ���������οn����_?au�> ��������>꿃>�W>��p>"`��3K��3��<�?G1-?�z�>N�q��(ɿ?A��m��<�[�?��@i)A?�@)�w���=e=�@�>�:	?�B>�`1���D�����>8b�?p�?�)P=	�V����p=e?jB<b6F�����:�=wڞ=p�=�a�4�J>s��>TG���@��G�M�4>�G�>��.�Y���a^��;�<x�]>�ӽ4i��5Մ?+{\��f���/��T��U>��T? +�>U:�=��,?W7H�a}Ͽ�\��*a?�0�?���?&�(?6ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�܅�=�6Ἲ���x���&V�t��=[��>e�>��,������O��I��T��=@:��7ƿ�='�� ���<1���2�E�h_���O���Qs��Z���y�i��F�G=��=k\>H��>��G>��U>ĵS?)ri?���>��>�Y�(��� ̾Y�k�l����2��������S������O޾��k3����b���!=�W
�=87R�F���g� �A�b��F���.?Hx$>�ʾ��M���-<�oʾĿ��(ф��ޥ��-̾ʗ1��!n��̟?1�A?�����V�$���O�����W?S����ꬾ���=����ۡ=�$�>J��=W�⾠ 3��~S���1?^?r;þ�|����4>�)���Q=�o-?�� ?O��`��>֗$?�2���ƽS1b>��@>���>��>�{>	����ֽy�?eR?����J�����>#[���xn�� |=��>�A�<�ɼ�h>��=�ъ��I��s铽��<�W?H�>o~*�'�	��������,=x?�v?� �>)hj?4RC?�s�<���nT�X��nEf=+W?��i?7)	>�����^о\���W6?+e?�M>��e��꾩E.�Y��@�?ޣn?�"?;����|�[ޒ�����"7?b�v?�q^��s��t����V�}=�>9_�>���>1�9��d�>*�>?6#��G��g����W4�@Þ?l�@2��?v�;<� �e��=�;?ZZ�>��O�J>ƾ����b�����q=�!�>4���dv����L,��8?���?���>$�����N��=(I����?�(�?̲2��\b�����[Y���f;׼mҒ<lt�D��<���F������iؾy�N�{a���>��@�#5����>:\����п$�¿x�����l�"����>�5�>Kӵ�.rC��wV�	HD���D�����S�>��>�Ô�������{�+l;��_����>��;��>۫S�3%��	����_6<�>��>���>K����罾eę?�_��a?οj���\��R�X?�f�?�n�?�j?��7<l�v�^~{�^n��)G?րs?�Z?�o%��4]���7��`?��3���j�[j�&�.�>�i�>�g�>:+���>>�'<<e�&?��=P�H��@¿ʿ�Z����?ZN�?k3ؾ�?�>���?��M?�D��k���QҾ���!��=��,?���=��q��,��4��1(��Q
?~4?!���]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?u$�>��?Ak�=\�>�b�=!�V�-��n#> �=�>�Ğ?��M?�I�>1C�=��8�� /�n[F��FR����C���>t�a?,�L?Eb>�&���&2�4!�6rͽ_a1�@L�z[@��,��߽%+5>}�=>a>%�D��Ӿ��?�\���ؿas��pS'�(-4?>�?��unt����D_?&t�>�B��,�� ,��-�����?L�?��?��׾�\ʼ=>S�>X�>�Jս�џ��a����7>^�B?m��@@����o�,�> ��?��@�ʮ?��h�A	? �P���_~���>7����=|�7?F/��z>���>��=Nnv�����=�s����>
B�?U{�?m��>�l?�o���B�N�1=�K�>!�k?s?�Wp�F���B>��?-��R����L�H!f?�
@Hu@��^?���Ϳ�lw���R�|��3Y���W��i:>�d=�V�>�x!>��Žl��<7/>� �>dT�>N �>��B>nB>펾=�~�l��%�����"�<��a�zc ����nu��'���B�ȣ߾f����ֽ�W��y�d����Vt�u�M���*>&�.?�`?�xj?\�>iDY��hM<��߾i.!=U]p������>��d?�Wb?˦?;()>X4v�7QR�
���K���
gξ��>��>�?;��>�a>�R==���>�S=c��><�>ی=�~��]p�f�o>���>1c�>�(�>~C<>��>Fϴ��1��k�h��
w�k̽1�?���R�J��1���9��צ���h�=Hb.?|>���?пe����2H?%���x)��+���>|�0?�cW?�>!��p�T�5:>7����j�=`>�+ ��l���)��%Q>ul?�f>�wu>�m3�M8��P�����J|>x6?#7���9���u���H�tZݾ�VM>���>e7D�\�����\�qLi���{=�i:?�u?�ӳ��᰾@�u��J����R>5J\>��=U\�=��M>��a�ƽ��G�1�-=��=O^>�?I�>}�=`�>�`����L�9Ҫ>�+=>��&>Z�>?^]#?�43��<c�e���D.��p>g��>>%�>�~	>�H�56�=���>��_>��ռ�΀��7���@�SD]>��_��x{�e�q=ޛ���n�=Ĩ=�k�f6�n��<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>��n�� ������x����=`d�=v6?��E�';�1��C#?��>��髿��̿Ї��-��>%��?�w�?-�`��ꟿ�\�' &?���?&�"?��>�	��y���>w�;?mt^?��>�z ���[�pB�>= �?�R�?��T>hb�?�bv?���>� ��%3�!_��3���%"Z����<{�y>>d�=֧��zN9����6̓�z�`���#E">�1=���>jٽQ��ib=�u���ĭ��2�����>H~>��>A
�>M?E��>6�>CU=�Ľ@r� <���K?o��?��r1n��-�<)��=��^��%?GH4?Bb[���Ͼ�Ө>d�\?�?T[?4d�>���>��9迿�}����<��K>|4�>�J�>�"���EK>h�Ծ@0D�Km�>�ϗ>/ϣ��<ھ�*��9W���B�>se!?���>TԮ={4?F�%?q_>���>-I�[m���;G�xS�>]��>@G?�{v?��?q���O6��!��#���H]�ͲI>�Ux?�?_̏>k���=5��DC;�4��絽'��?�ba?�h���?@�?�B?3�=?yie>7� �f�ؾƯ����>��!?_��7�A�zA&��n�^|?uj?a��>���_�׽�fм������e?�'\?+W&?�X���`�sþ#��<��"���H��f�;�C���>�6>���F�=PN>��=��m�6��l<Ш�=���>�Y�=7:7�/c��/=,?��G�{ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U�� �?���?Yk�?h��>�h��$=?�?Q	?f"�>�J���}޾7���Pw�~x��w�\�>���>ʢl���J���ڙ���F��j�Ž�'�t�>E��>�]?DQ?d�e> �>/�h��)��)���ξ��I����~ ,��7�� �����Y9���$=�ž��a��=�>��ټ�M�>
�?j��>��c>Q�?�x;	��>�F>8��>�L�>�D�=7n=�O	> �*>�W���Q?N@¾d6'���'篾�A?�Ud?���>��h�r����Ͷ?]��?w�?U	v>�7h�ݿ*���?�%�>���1?�;7=1g�{P�<�E����z���3�C{�>?%ٽI�9�uM�J�e��8
?�p?�<��c�̾3�ܽ<��V^�>s�?�?|�F��Jy���g��Ð��,�Qr��&پQ����k�Z[���닿l�{�*쌿+�k�	G��?;?���?��򾔿��h���4)�E����o����>=�?�X�=aO>4��5�E�R�����I�]���_0�>n?w�>&�;?	~:?��V?̖M?6��>�ި>�訾��>��,=�g�>��>�3C?v�.?7�3?@q?��7?XI>6�,����vež�?eS�>�/&? �#?(�?���$��A:�x�<T����o6�|�{= <�=��(�ٹ5=L�>s�x>Ae?�)p��O�vv5��T>��7?�*p>�.�>�^ʾo))�Doo��?y[?�2�=���@���*��Q�>�?o�˼<�=�(>�48=�h�=�ǽ.�=�<%��=�A=@�4� =�=XC�=�R�<E�,�*�����|<��>u�>5�?���>�C�>{@��%� �L���e�=Y>S>�>�Eپ�}���$��i�g��]y>�w�?�z�?e�f=�=��=}���U�����O���S��<�?&J#?XT?Y��?|�=?Kj#?ϵ>+�eM���^�������?L ,?X��>B����ʾ�䨿�3�{?�a?a9a�u�>)�wQ¾��Խ@S>g/��=~�e���D��e�����\�����?���?M�@���6�*��r����:����C?��>�c�>���>��)���g���T;>�t�>]�Q?h5�>�� ?�r?�ok?+$>OW	�����ᕿ��E>_�>G;?���?��?��c?HD�>��>�l��'pӾ�|�ɀ���:������p�<0h>���>��>�c�>��>6�ý�	�=0�S��(L>���>�?�&�>�k*?g�>�RL�"I?`m�>�þ���	@��9!l����Nn?�5�?�� ?�=����vA����e�>��?��?�h1?�?X��>O�Ѽ�ƾ�m���>���>���>���=y�<�q�=rz�>{�>�F(�r���>�����w�
?�C?嵪=h�ƿ+_r��9y�Z3�����;���V_���u�ڼW���=�w�����
|����[��Ǚ����>ò�lN����x����>C\�=�>A$�=��<��ͼY�<�I4=~e<6z=��b��_<��E�N(�;]ᓽ�z��$�v<�QN=I�5���˾?�}?&=I?a�+?q�C?նy>�1>��3����>�o��k>?�V>�P�σ��D�;�襨����?�ؾ�z׾A�c�Ɵ��F>hI�ٮ>X83>�U�=Gև<�"�=�ss=^�=�_N�$=Y�=�b�=]|�=���=��>�V>/Vw?zH��B�����P�3��`�:?�N�>�<�=��žh�>?o�A>�փ��p��j��(?N��?�^�?�1?��i�@�>Y���sL���F�=����Z2>(��=73���>��K>�M��R���걽�&�?Ԇ@�M??mŋ�VϿ-/>�:>NZ>�S��D1�m�Y�1�`��hU��!?��:�\�ξoՇ>KN�=�߾��ľՎ0=:�9> �t=B$��	\�tՙ=W>z�HL==I�f=�j�>��B>��=���˕�=k�G=�(�=y}O>f	���e1����e<=���=�La>"l%>\��>=i?�G.?��d?���>�6N��>þ ��˴�>��=M�>Xw�=U>h7�>=+8?T�E?&"O?1��>��P=_�>� �>hA+�o�j�$پn2��+=�͈?e\�?cP�>vC�<��\�͝!���8�ه���?��4?�&?M��>��ҿ��X�V�@��F}�ޫ<g.�=��=>F�%=Ѫ%�m�c�Բ����;^KZ>R�?-o�>N�\>7!n�B�u=�P�>n�8>+KH>��=��<�	��R�<s��<�m�D!=堻=Jl��J@�k��:���+H��h�==�����=���=���>Q>���>�c�=5���[x.>jx����L����=�1��mB�$d�mJ~��/�a�6�
B>ףW>=����.��W�?�`Z>�@>�s�?�[u?S�!>�B��yվ�R����c�6.T�f��=�1
>Q=�F;�I(`��M���Ҿ�>3�>e�>��
>�#
���C�OV��@��;�@�b�>p9���C�=?��1���W��V����k�&���LRW?؅�Jc=��?�`y?���?{��>��>�M��y�=�˾o!H>;@���ተ=z�?��H?,?W�� 8v�_8̾)Q��j�>��H��P�d���
s0���*�V;����>�����оg-3� ]��3����B���r�κ>W�O?_߮?h!c�L��3<O�#��΅�/#?�Qg?�;�>�n?�?If��"��얹=��n?���?4�?��>�Z�=���=�>��
?*�?G�?�p?��M��>�>F=
��>QϽ0�>��1>% �==�=��?r�?�6?��c��(� �ܾ�@�Q~>�#�=i!>�`�>���>O�~>�7�=*!ż�PF�|U>ɲ�>O9[>��]>�l�>O��>Y���ޛ3�=�/??�>K�>3?o�>~h=��n��:�>-NW=
p��n���/�k�a�5����0�>�Ej>���>��ѿU��?dc�>���!�>��ѾzD�!�N=V|>6�Ⱦ�M>2�>P�;5�%?Xv?*`�>�L�>�A0=������>�! ���%�Kd��H�7�x`9=}.�К�{(�I`��
	�����U\)��-w�����@�8��=��?G�
��8��)sT�I�ǽ�'?�/2>�O`?9�9֪�#>�?���>C��G���"��ٵӾՕ?��?�c>�ݞ>\�W?(�?�"1�w+3�`Z�ޝu��A�- e�߰`�`捿ǅ���
��ѿ�&�_?*�x?�yA?2Ǒ<+z>S��?��%�0ُ���>� /��3;�4�:=��>���a�I�Ӿ�ľ���B'F>Փo?��?�?r�V��I��a>�~>?�9?7$l?N�.?@,?��>��`"?(!Y>5v?^�?r.?f)?@�??I>���=Z����7<�\���ȁ�gٽ$Ž�Xy�dLi=� �=� �<j=�>�=Ԥ�=��<����Ú�<�=:9�<��=S�=�Ŧ>�]?_G�>^��>n�7?���]l8�-���(/?S9=�������������� >9�j?}��?�^Z?u?d>|�A��	C�*>U�>8a&>�!\> a�>���G�E�/2�=�n>�H>�s�=F�M����	�ʎ���@�<�6>e��>�!|>rЍ���'>�p���0z�J�d>i�Q��ú�}�S�W�G���1�#cv��[�>0�K?��?���=�^�X���Af��))?�Y<?�KM?��?X6�=2�۾$�9�j�J����"�>ȸ�<�	����� ���:��G�:�s>�%��sj����>A8辡ʾ=9q���K�ȭܾD�=�>�#����=�	����Ņ�f��=���=%﷾����LŨ�g�D?�=�����[�OC־��=���>H×>L�%��>��Q@�gc��a�=!��>�/>�����YE�R����>�SS?��i?J�q?��Ǿ�ls���-��k�b$��"==h�>z�I>���>�Z>��=���������
n�^lS�vh�>�f�>	�#1�U�þT?� �!PB>��?�x5>_��>Ɩ:?4�?b?�?8��>%�6>P/���Ͼa=&?D��?�`�=�Խh�T���8��F�m��>�)?�dB��͗>��?A�?��&?�Q?�?�>[� �
G@����>�Y�>��W�1X���A`>��J?렳>�DY?3?��=>�q5��+��G$��͟�=�G>O�2?�I#?��? ��>��7?�T�m����Qh>5z�?IŌ?[�?���>��>�X�1�k?os0=(D��9�J?��??y*l?�ړ?��??��=���=?3��.�i���n���)�����<��7=F=�۰�B�<�s�<6}^<�t=���<�#����W��=\(�;�.�>?s>+s��12>tþ�o���yE>rE��7љ����O�3�*Q�=�;�>�E?�o�>ޱ*� �=��>f�>׽��$&?�?I@?� ��aVb���ھs-M�e�>��B?~��=��l������u�M�p=3lm?E�^?MQ��,��>�b?�]?_h�=���þ�b�m��o�O?�
?1�G�i�>��~?'�q?v��>��e�U:n�+���Cb���j�(ж=4r�>�W���d�e?�>�7?RN�>��b>�$�=ju۾��w��q��D?[�?�?���?�+*>p�n�Z4��%��ލ�k+X?i$�>�䒾f�?%�R���̾E���K�ʾEW��پ���dl��c�����܎���_h=$�?�i�?�`w?u�^?|���7�u�!z��I����6�F�������YA�^�I�>\~�%3(���:�Ծ}�j;��K�iC�Ԣ�?3/?���3�>�u��,�����= D>O$��?����>Oཽ܈+=��7=�j9�`�����P�?��>L�>�L?�M�+���$���1�Y����|�=�ъ>��>�n�>��=wm,�ϯ��cθ�Mذ�F1a�$p>��a?�H?1ub?~
���.�3�1�U���蝾}&>lc�=�s�>*Z�W�0��!�_<���p��x
�Au��X�����=nA5?S-�>b��>Ӈ�?~D?����ƾ`2�!�2�)��='�>�YZ?���>ȸu>��}�!�%��>��l?�t�>�&{> ��_�$�����D�p����>�9�>��>�b�>�G/��c�R����\���N>�{>�=�u?KV��W�[�ۥ�>׾b?��;������>�ޏ�����@���h����=p/?C�=�gM>_�������.�w��ة�T�*?��?�����)�tՂ>>�!?x;�>!p�>�T�?$œ>� ��K�:_�?��_?!�J?
�B?��>�H=� ��Ƚ��%�#f<=0��>d�Z>��p=qy�=�����U����wC=j{�=^����s��m��<N����4�;4�<��2>�ڿ�I��{;�
���� �
�+Q����½;���3�&��a���W�����,s�*�دN���l�:哾�Zv�f=�?��?�|���v�����悿f<���>zn�p�`��}���$Խ�+���.�r���)��
V���m��`��'?ΐ��ǿ���'�۾w9 ?�-?�~y?}p�<"�Г8���">��<nҳ���������οn����_?au�> ��������>꿃>�W>��p>"`��3K��3��<�?G1-?�z�>N�q��(ɿ?A��m��<�[�?��@i)A?�@)�w���=e=�@�>�:	?�B>�`1���D�����>8b�?p�?�)P=	�V����p=e?jB<b6F�����:�=wڞ=p�=�a�4�J>s��>TG���@��G�M�4>�G�>��.�Y���a^��;�<x�]>�ӽ4i��5Մ?+{\��f���/��T��U>��T? +�>U:�=��,?W7H�a}Ͽ�\��*a?�0�?���?&�(?6ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�܅�=�6Ἲ���x���&V�t��=[��>e�>��,������O��I��T��=@:��7ƿ�='�� ���<1���2�E�h_���O���Qs��Z���y�i��F�G=��=k\>H��>��G>��U>ĵS?)ri?���>��>�Y�(��� ̾Y�k�l����2��������S������O޾��k3����b���!=�W
�=87R�F���g� �A�b��F���.?Hx$>�ʾ��M���-<�oʾĿ��(ф��ޥ��-̾ʗ1��!n��̟?1�A?�����V�$���O�����W?S����ꬾ���=����ۡ=�$�>J��=W�⾠ 3��~S���1?^?r;þ�|����4>�)���Q=�o-?�� ?O��`��>֗$?�2���ƽS1b>��@>���>��>�{>	����ֽy�?eR?����J�����>#[���xn�� |=��>�A�<�ɼ�h>��=�ъ��I��s铽��<�W?H�>o~*�'�	��������,=x?�v?� �>)hj?4RC?�s�<���nT�X��nEf=+W?��i?7)	>�����^о\���W6?+e?�M>��e��꾩E.�Y��@�?ޣn?�"?;����|�[ޒ�����"7?b�v?�q^��s��t����V�}=�>9_�>���>1�9��d�>*�>?6#��G��g����W4�@Þ?l�@2��?v�;<� �e��=�;?ZZ�>��O�J>ƾ����b�����q=�!�>4���dv����L,��8?���?���>$�����N��=(I����?�(�?̲2��\b�����[Y���f;׼mҒ<lt�D��<���F������iؾy�N�{a���>��@�#5����>:\����п$�¿x�����l�"����>�5�>Kӵ�.rC��wV�	HD���D�����S�>��>�Ô�������{�+l;��_����>��;��>۫S�3%��	����_6<�>��>���>K����罾eę?�_��a?οj���\��R�X?�f�?�n�?�j?��7<l�v�^~{�^n��)G?րs?�Z?�o%��4]���7��`?��3���j�[j�&�.�>�i�>�g�>:+���>>�'<<e�&?��=P�H��@¿ʿ�Z����?ZN�?k3ؾ�?�>���?��M?�D��k���QҾ���!��=��,?���=��q��,��4��1(��Q
?~4?!���]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?u$�>��?Ak�=\�>�b�=!�V�-��n#> �=�>�Ğ?��M?�I�>1C�=��8�� /�n[F��FR����C���>t�a?,�L?Eb>�&���&2�4!�6rͽ_a1�@L�z[@��,��߽%+5>}�=>a>%�D��Ӿ��?�\���ؿas��pS'�(-4?>�?��unt����D_?&t�>�B��,�� ,��-�����?L�?��?��׾�\ʼ=>S�>X�>�Jս�џ��a����7>^�B?m��@@����o�,�> ��?��@�ʮ?��h�A	? �P���_~���>7����=|�7?F/��z>���>��=Nnv�����=�s����>
B�?U{�?m��>�l?�o���B�N�1=�K�>!�k?s?�Wp�F���B>��?-��R����L�H!f?�
@Hu@��^?���Ϳ�lw���R�|��3Y���W��i:>�d=�V�>�x!>��Žl��<7/>� �>dT�>N �>��B>nB>펾=�~�l��%�����"�<��a�zc ����nu��'���B�ȣ߾f����ֽ�W��y�d����Vt�u�M���*>&�.?�`?�xj?\�>iDY��hM<��߾i.!=U]p������>��d?�Wb?˦?;()>X4v�7QR�
���K���
gξ��>��>�?;��>�a>�R==���>�S=c��><�>ی=�~��]p�f�o>���>1c�>�(�>~C<>��>Fϴ��1��k�h��
w�k̽1�?���R�J��1���9��צ���h�=Hb.?|>���?пe����2H?%���x)��+���>|�0?�cW?�>!��p�T�5:>7����j�=`>�+ ��l���)��%Q>ul?�f>�wu>�m3�M8��P�����J|>x6?#7���9���u���H�tZݾ�VM>���>e7D�\�����\�qLi���{=�i:?�u?�ӳ��᰾@�u��J����R>5J\>��=U\�=��M>��a�ƽ��G�1�-=��=O^>�?I�>}�=`�>�`����L�9Ҫ>�+=>��&>Z�>?^]#?�43��<c�e���D.��p>g��>>%�>�~	>�H�56�=���>��_>��ռ�΀��7���@�SD]>��_��x{�e�q=ޛ���n�=Ĩ=�k�f6�n��<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>��n�� ������x����=`d�=v6?��E�';�1��C#?��>��髿��̿Ї��-��>%��?�w�?-�`��ꟿ�\�' &?���?&�"?��>�	��y���>w�;?mt^?��>�z ���[�pB�>= �?�R�?��T>hb�?�bv?���>� ��%3�!_��3���%"Z����<{�y>>d�=֧��zN9����6̓�z�`���#E">�1=���>jٽQ��ib=�u���ĭ��2�����>H~>��>A
�>M?E��>6�>CU=�Ľ@r� <���K?o��?��r1n��-�<)��=��^��%?GH4?Bb[���Ͼ�Ө>d�\?�?T[?4d�>���>��9迿�}����<��K>|4�>�J�>�"���EK>h�Ծ@0D�Km�>�ϗ>/ϣ��<ھ�*��9W���B�>se!?���>TԮ={4?F�%?q_>���>-I�[m���;G�xS�>]��>@G?�{v?��?q���O6��!��#���H]�ͲI>�Ux?�?_̏>k���=5��DC;�4��絽'��?�ba?�h���?@�?�B?3�=?yie>7� �f�ؾƯ����>��!?_��7�A�zA&��n�^|?uj?a��>���_�׽�fм������e?�'\?+W&?�X���`�sþ#��<��"���H��f�;�C���>�6>���F�=PN>��=��m�6��l<Ш�=���>�Y�=7:7�/c��/=,?��G�{ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U�� �?���?Yk�?h��>�h��$=?�?Q	?f"�>�J���}޾7���Pw�~x��w�\�>���>ʢl���J���ڙ���F��j�Ž�'�t�>E��>�]?DQ?d�e> �>/�h��)��)���ξ��I����~ ,��7�� �����Y9���$=�ž��a��=�>��ټ�M�>
�?j��>��c>Q�?�x;	��>�F>8��>�L�>�D�=7n=�O	> �*>�W���Q?N@¾d6'���'篾�A?�Ud?���>��h�r����Ͷ?]��?w�?U	v>�7h�ݿ*���?�%�>���1?�;7=1g�{P�<�E����z���3�C{�>?%ٽI�9�uM�J�e��8
?�p?�<��c�̾3�ܽ<��V^�>s�?�?|�F��Jy���g��Ð��,�Qr��&پQ����k�Z[���닿l�{�*쌿+�k�	G��?;?���?��򾔿��h���4)�E����o����>=�?�X�=aO>4��5�E�R�����I�]���_0�>n?w�>&�;?	~:?��V?̖M?6��>�ި>�訾��>��,=�g�>��>�3C?v�.?7�3?@q?��7?XI>6�,����vež�?eS�>�/&? �#?(�?���$��A:�x�<T����o6�|�{= <�=��(�ٹ5=L�>s�x>Ae?�)p��O�vv5��T>��7?�*p>�.�>�^ʾo))�Doo��?y[?�2�=���@���*��Q�>�?o�˼<�=�(>�48=�h�=�ǽ.�=�<%��=�A=@�4� =�=XC�=�R�<E�,�*�����|<��>u�>5�?���>�C�>{@��%� �L���e�=Y>S>�>�Eپ�}���$��i�g��]y>�w�?�z�?e�f=�=��=}���U�����O���S��<�?&J#?XT?Y��?|�=?Kj#?ϵ>+�eM���^�������?L ,?X��>B����ʾ�䨿�3�{?�a?a9a�u�>)�wQ¾��Խ@S>g/��=~�e���D��e�����\�����?���?M�@���6�*��r����:����C?��>�c�>���>��)���g���T;>�t�>]�Q?h5�>�� ?�r?�ok?+$>OW	�����ᕿ��E>_�>G;?���?��?��c?HD�>��>�l��'pӾ�|�ɀ���:������p�<0h>���>��>�c�>��>6�ý�	�=0�S��(L>���>�?�&�>�k*?g�>�RL�"I?`m�>�þ���	@��9!l����Nn?�5�?�� ?�=����vA����e�>��?��?�h1?�?X��>O�Ѽ�ƾ�m���>���>���>���=y�<�q�=rz�>{�>�F(�r���>�����w�
?�C?嵪=h�ƿ+_r��9y�Z3�����;���V_���u�ڼW���=�w�����
|����[��Ǚ����>ò�lN����x����>C\�=�>A$�=��<��ͼY�<�I4=~e<6z=��b��_<��E�N(�;]ᓽ�z��$�v<�QN=I�5���˾?�}?&=I?a�+?q�C?նy>�1>��3����>�o��k>?�V>�P�σ��D�;�襨����?�ؾ�z׾A�c�Ɵ��F>hI�ٮ>X83>�U�=Gև<�"�=�ss=^�=�_N�$=Y�=�b�=]|�=���=��>�V>/Vw?zH��B�����P�3��`�:?�N�>�<�=��žh�>?o�A>�փ��p��j��(?N��?�^�?�1?��i�@�>Y���sL���F�=����Z2>(��=73���>��K>�M��R���걽�&�?Ԇ@�M??mŋ�VϿ-/>�:>NZ>�S��D1�m�Y�1�`��hU��!?��:�\�ξoՇ>KN�=�߾��ľՎ0=:�9> �t=B$��	\�tՙ=W>z�HL==I�f=�j�>��B>��=���˕�=k�G=�(�=y}O>f	���e1����e<=���=�La>"l%>\��>=i?�G.?��d?���>�6N��>þ ��˴�>��=M�>Xw�=U>h7�>=+8?T�E?&"O?1��>��P=_�>� �>hA+�o�j�$پn2��+=�͈?e\�?cP�>vC�<��\�͝!���8�ه���?��4?�&?M��>��ҿ��X�V�@��F}�ޫ<g.�=��=>F�%=Ѫ%�m�c�Բ����;^KZ>R�?-o�>N�\>7!n�B�u=�P�>n�8>+KH>��=��<�	��R�<s��<�m�D!=堻=Jl��J@�k��:���+H��h�==�����=���=���>Q>���>�c�=5���[x.>jx����L����=�1��mB�$d�mJ~��/�a�6�
B>ףW>=����.��W�?�`Z>�@>�s�?�[u?S�!>�B��yվ�R����c�6.T�f��=�1
>Q=�F;�I(`��M���Ҿ�>3�>e�>��
>�#
���C�OV��@��;�@�b�>p9���C�=?��1���W��V����k�&���LRW?؅�Jc=��?�`y?���?{��>��>�M��y�=�˾o!H>;@���ተ=z�?��H?,?W�� 8v�_8̾)Q��j�>��H��P�d���
s0���*�V;����>�����оg-3� ]��3����B���r�κ>W�O?_߮?h!c�L��3<O�#��΅�/#?�Qg?�;�>�n?�?If��"��얹=��n?���?4�?��>�Z�=���=�>��
?*�?G�?�p?��M��>�>F=
��>QϽ0�>��1>% �==�=��?r�?�6?��c��(� �ܾ�@�Q~>�#�=i!>�`�>���>O�~>�7�=*!ż�PF�|U>ɲ�>O9[>��]>�l�>O��>Y���ޛ3�=�/??�>K�>3?o�>~h=��n��:�>-NW=
p��n���/�k�a�5����0�>�Ej>���>��ѿU��?dc�>���!�>��ѾzD�!�N=V|>6�Ⱦ�M>2�>P�;5�%?Xv?*`�>�L�>�A0=������>�! ���%�Kd��H�7�x`9=}.�К�{(�I`��
	�����U\)��-w�����@�8��=��?G�
��8��)sT�I�ǽ�'?�/2>�O`?9�9֪�#>�?���>C��G���"��ٵӾՕ?��?�c>�ݞ>\�W?(�?�"1�w+3�`Z�ޝu��A�- e�߰`�`捿ǅ���
��ѿ�&�_?*�x?�yA?2Ǒ<+z>S��?��%�0ُ���>� /��3;�4�:=��>���a�I�Ӿ�ľ���B'F>Փo?��?�?r�V��I��a>�~>?�9?7$l?N�.?@,?��>��`"?(!Y>5v?^�?r.?f)?@�??I>���=Z����7<�\���ȁ�gٽ$Ž�Xy�dLi=� �=� �<j=�>�=Ԥ�=��<����Ú�<�=:9�<��=S�=�Ŧ>�]?_G�>^��>n�7?���]l8�-���(/?S9=�������������� >9�j?}��?�^Z?u?d>|�A��	C�*>U�>8a&>�!\> a�>���G�E�/2�=�n>�H>�s�=F�M����	�ʎ���@�<�6>e��>�!|>rЍ���'>�p���0z�J�d>i�Q��ú�}�S�W�G���1�#cv��[�>0�K?��?���=�^�X���Af��))?�Y<?�KM?��?X6�=2�۾$�9�j�J����"�>ȸ�<�	����� ���:��G�:�s>�%��d���,�Y>US��!����j�&�X����+��v�CD�=����ԾdI^����=��=�Ǿ�|'��䠿�^����P?�T�=q����� `̾V��=��>*O�>���'���B������5=�Ο>�=Qf7����\�S��S�ߑ>�K?<�Y?�x?�{����q�1vZ��vܾ�Y�N2>���0?9(�>HT�>��=M�׺��о ����p�7th�dq�>]��>�:A�!�=�~m侦f����(�\��>�?�>���<�;?9V?��,?�u?l�?*�.?轺>��"��,���?'?���?�4��Uu���˾�h�S�`����>�6?Ir���/�>�)?�^?;
?1H?�� ?��Z>�w��Ul�eb�>�٥>t�;ף�K(i>>B>?:�>8C??2"�?'J�>�qW�)Ͻ��d���a>�6>�?y"J?_|6?{�>X�>�O���x=�[�>@Xi?�׆?��a?��=<@?�6>���>O4�=+\�>��>+?��@?(�f?��S?���>��<�A��E}��(���;���3���=����r����N��w<	r�;��h<��]9UE��\��ۇ＂�C�?��>��_>�Ë���5>��;�]�E3>ijҼ����	������A=y�!>ͤ?�Q�>�r4�e@k=��>���>7���p7?h/?(^J?S�=�#�V�G_��Ú���8�>�!?��#>@�T����^��R<$�r?a?�Q�)N��U�b?��]?�_��=���þ�b�`����O?>�
?	�G�L��>\�~?2�q?���>�f�7n�T���Fb��k���=�u�>^a���d��.�>��7? F�>%�b>�/�=w۾Ҽw��b��  ?n��?���?���?�E*>2�n��1��t���琿N\?�-�>7`����?��v�Z�Ѿ�Ō�+��8[�Nת�����敏�����'�q_��D�����=��?_�u?KLo?P�d?B���Pe�r�Z�߀�`�X�lD�A�q�D�lB�x.A��qo����������;�F=�;t�v=��R�?y�!?l)�yV�>k����q�y6˾F9Y>�J�����ψ=��`�h�z=8j#=J�u��5�����
�?$��>��>>�G?��d���<���(�"�<�, ��S'>�՜>���>j�>��;�.��Y׽b.���M��P����Ev>�~c?T�K??�n?"[��I1�gu��&{!��,��z��'IC>��>��>��X��F�,�&�$b>�#�r�c��Fx����	��"�=ņ2?�_�>$��>:�?-�?�N	�yj����x��1���<��>|%i?``�>y��>Mjҽ!�ª�>8yd?G��>h�>�f�xQ;�rp�fuٽ:}�>�t>*�,?��> �����j�n��`﬿��#���_>�lk?�*��6uu�x�> ;R?V�>����-��>$ ;�J���������ap���S�>���io�>@���$������;��)?�_?�˞�l�*�i�m>�C?hP�>��>�B�?�4�>�<����&<�g?�]?�2G?QD=?E5�>�,=�����ν˗ ��oA=	܆>��h>X7=T��=-�>�S��� ��#=Q?�=~c�hI½�Zu<���&Z<C�0=G+H>oڿ�F�f~���f׾�Ⱦ��ղ���`�ፚ�S��������}���^M��0J�M�мO�C��M��;�β�u�?ј�?RSS��Q;�����,�������<->������;�~Ծ�t�3��J���=���0?.��zO�C�����a�[�'?����^�ǿ#����-ܾ(  ?�< ?�y?/��"��8�=� >@��<�"��o��=���1�ο˨��-�^?���>���� ��>���>�X>�=q>e��=枾��< �?5�-?{��>��r�7�ɿ݉��O�<��?�@�rA?o�(�6�쾗~S=�1�>C�	?#?>m1�����-���e�>�<�?��?^M=��W��
��e?��<��F�y=�Q�=���=TP=�6�~�I>���>0O�b�@��۽54>��>)"�~��s6^�Ǿ�<�X]>\Խ�#����?hڃ�������P�yP���=(y�?�G?a�$�W?:�;�ܿ<p���ǫ?Q��?���?���>vOY�+|g>*Ͼ\?1�&?�d�=F�⾢�l����Ȋʽk�6��Ӿr�L��ڒ>H����ʽBDr��x��S;۽dA=�]�>���/ƿ��!��W���=4��K�o�e,�����P#N�uM����l�#Y꽁�s=س�=A!R>���>��M>i~L>6X?�dn?Յ�>-%>+��쮒�s�;"�|����G���s��$�!��r���`�G)�zI
����Z^�9�ʾ?=�Qэ=�7R������� �5�b�=�F�y�.? s$>*�ʾ��M���*<O�ʾ𱪾rփ��[O̾œ1��
n��ß?	�A?�腿^�V�\����3_��'�W?WM�Ĥ��鬾���="#���=v,�>]D�=���3�~tS���(?��??�U���:��N&�=l�&�N嵻�� ?�,?�E.���>6�L?�+0��]�I�$>/Q�=3t�>.�>m�=]������K#?TW?|W>����3��>�䩾�J���E?�Z�>���.{�<��=y�	>+i������g>�WV?���>��(������������߮=YQv?Jg?�c�>�cm?�C?�O<��U��Z
�V�=�=X?��i?��>��|� G;3|���-4?�`_?��K>ܧf���羏P+�(��\F?\nl?>�?��������뒿�!�z�5?��v?�r^�ps�����{�V�v=�>�[�>���>��9��k�>�>?�#��G������~Y4�'Þ?��@���?R�;< �|��=�;?0\�>�O��>ƾQ{��|����q=�"�>Ԍ��gev����3R,�J�8?Ҡ�?|��>����©���=�ؕ�=Z�?�?焪�.g<����l�Wn�����<5ϫ=���E"�X���7�A�ƾ�
�����j鿼+��>�Y@�R�5,�>G8�#6�	SϿ ��	^оOq���?B�>�Ƚ����J�j��Pu���G���H�/���O��>�UL<4˽ʍ7� τ��HJ��P�=���>�᛾�-{>�^�����Ͼ_�->e|�>P�?\` ?�= ��X��?��/�{#�Ԯ���!���?^�?�z�?�d�?��Z�<�(�deo���=>�ۀ?���?�8?�u���Ⱦ��{��i?ZF���(\���5��oH��n[>[�*?���>"(�u%<=V�6>��>@��=��-���Ŀg���i*����?E��?t�侉��>��?��,?�������������'�;m���D?��$>�὾�;�3�>�,T�����>)?�����?u?@�w������9�|1@����>>���=0����ng<WD��r��~/�uо?<+�?S��?�ˋ�Xr��%�>ҁ�>����۾�F6=�9?0r�>-e�>���/ф>\d�����.t����?o8�?h��>r�d�����~z�=st?Mٶ>�w�?A�=$� ?�>�*��J$��C�)>�>[>�6A��?��]?�F�>�?j=~��> ��T-���?�ˁ��n�?�6��>��x?�X?�Ѳ>�G���0ʽ(��X���������^��Aͻ�,���nt>*�>��D=��N�/�ξ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?C��N��]~�����
7�M��=��7?�6��z>���>{
�=�nv������s�鸶>�B�?;{�?��>��l?��o���B��1=�J�>M�k?�q?�'m��ͬB>ζ?�������OH�r"f?��
@ou@ϝ^? Z�˿i����Ա���~�/�!>�W�=4�U>ڕH����%?V>����ULv�y><��>�d/>�s�=+�:>���=cs=nԀ��f%�þ��^x�[0�`���������+�cǑ�;7%�	��6g��B�N�]�R!�t��KP/���ؽ[b�=s�\?�|S?+�r?k�
?{G���*�=J����=�JP��'�=���>��6?ۂB?�G,?K��=*~��v�Z���{��款�ƈ�v��>��?>&@�>���>���>�&�<�<M>y�I>+Bo>8Z�=Zt�<;w����m= �h>ʓ�>lf�>p=�>+g<>�T>&ʹ��/���Ph�A�v���̽4��?zb��ʗJ��9���a��~߷��Y�=-S.?�L>����+п�׭�WH?R���;�+�H�>�0?�.W?�>�鰾�?Q�>���Wj�]�>���P�l��w)��Q>�H?�n�>B&>P8���P�=���r���.#>r�??�\��p��ϊ���F������C>!��>{3��8�ң��>[O��67�Q�=�%;?�M?1s]�R�����N��NϾ�*%>���> �h<��=��I>yT=@Tm�j�i�z%�=���=ݡ3>N�?=g,>N��=輢>32���(H��o�>>>��->��>?��$?0�7A������R�*��'r>���>�$�>��>�&H�ot�=~(�>�b>���f~������B��7N>�߇�q�b�;�r�"*�=^������=1%�=b���?��=3�~?W������?�c���o|D?��?��=��><��!�n������ �?��@���?���?jV��?|	�?�B�����=V��>g��>�;�+M�H�?�KŽͧ��y	��L"�{�?���?��1���k���>%%?�9ӾPh�>{x��Z�������u���#=L��>�8H?�V����O�r>��v
?�?�^�ީ����ȿ7|v����>V�?���?h�m��A���@����>:��?�gY?ioi>�g۾(`Z����>ѻ@?�R?�>�9���'���?�޶?ԯ�?;+P>�.�?�?!�>���l�:�!q���&}�vk>����£>��!>�R�"�^�Sg��\ٕ��/l�KP�7!>�OH=�6�>�{Խ�B���+[<�Ҟ���ھ��ϼ��>��><+~>_��>��	? ^�>��>�W>�X�pƾ^��S�K?�Ώ?�r��n����<Q�=��_�/?W�4?��u�� Ͼ"l�>�\?(j�?}#Z?3��>�e��˚����r]���<�]J>���>�`�>����R�O>!Ծ��@��I�>ƻ�>mG��BAپ""���1��ۛ>h>!?]��>\�=�x ?��#?;�j>���>�KF�{���O�F�q@�>]�>�?��?��?�����)3��H������Z�8R>t�y?��?��>�Ў��#��.%�}�|��T���'�?-<f?Xֽ�]?ف�?�??I�??�~e>�1�3ھE���!~>��?��!��QO��.4���m�H�?���>���>��`��	���A�"�g��A?�HO?�?�'Y� v���ܪ<����[P=�-m�v��;$�K>�"�=+� �\o�=�d�>}�=�JB��r����=��>�bS>{-�=��u#���;,?]�F�kփ����=m�r�1jD�E�>7BL>b���͖^?b(=���{�m���r��`4U����?S��?^j�?�`��>�h�<"=?��??;#�>�s���v޾ʄ��Cw��Ex�=x���>���>ٻp���ǖ�������C��+ ƽ'��bv�>��>c�?�r?��?>��>`k���s$�I�������^�����4��.+���������8�������؃�[̓>2���eN�>*?�<;>M>K��>��?=�F�>�fK>�>�>e�>'S>�>(��=��<$��cGR?����ܷ'����\���)1B?�dd?�-�>>i��y������n?�{�?gn�?hv>uh�.+�Mg?"9�>����z
?�;=����"�<�[�������������>�?׽:�&M��7f�ef
?�*?L���ou̾��ֽt�Ӿ�R�<�+�?��q?F�/��'����>�{�G㎿g�F><�쾴%޾�<$�u�l�3�������d�������m䷽	'?�G?��Z�_��l�t��y�I�k�0;s>��3=`�5>�H>/�Z=8%��� �(�K�'����-�+L?M�?b��>�&[?�M=?��V?p$Z?�_Y>��_>�B���(?����˥>'�?z�A?,�?��0?y�?��?�;U>�������`̾��'?�f?��!?�Q�>��>b=E��h����6=t��)ᐾ̫��LB=���=\ػ������=��)>�6?|½�%�]����:�>�M?���> �>7\a��V����=�:�>�\?�=_>�޾�g���� ?h�t?�ۼ���;Q[7>-��=�ߨ��v�k�>M[�<OB�ɒ��U���&.���=#o)>{�=�G�2��:�%Z=tOW��N�>dF?�gK>gR�M����=��+�Z�V��1�>2˄�s�>|��������u�������>�Ԥ?��?�;�>�$�=�ϙ=�}4����J	��x¾�iν�k�>P�+?0}1?�?��c?�t�>w&>��<C���Հ�;�����>�,?�.�>���#˾���_*3�=d?�Y?��`�����)�H�¾ �ֽe>k�.��~���x�C� Xm�Ў�#��?�?�.O��6���;ј�����n<C?��>�Z�>.��>5\)�$g� ��g=>���>R?g�>��O?g:{?ܞ[?��T>P�8�
)��Tə��/���!>�@?�?C�?ty?��>m�>�)���߾PN����,�������V=m�Y>+��>� �>��>,��=P�ǽ�e����>�3T�=�{b>���>횥>}��>|xw>�i�<�gF?���>���� �������d�~C����f?���?��?�[�<���{�J��� ���>��?���?o.?�I#��K�=9�&����L����>�
�>G��> �=p��="��=��>s�>��׽;O��?��8��+?�fG?;�c=�[ƿ�5{�\���ƥ�N8!=�N~���P�K�6���`�ک�=5���h&������7a������)������Vr��*]{��!�>c�{=ub>C�=�?ɼlN��b�D=��=���<c>�Q�]|!<ү\�d��Vʭ��Sػ���D�x=���<�������?n�`?�?�e?�&Y>-�<�ʜ=$.�>/���?��>~��=z���� ��>��w����傾!<��rb�}Yƾ�@�=�`�^7�=�k>�[�=ޗ��W?�=��=nf�=Q�.==�;R=�=�<��[=!��=8E�=�6w?\�������4Q�T[罥�:?9�>�|�=��ƾp@?\�>>�2������Fb�.?y��?�T�?/�?�ti��d�>���g䎽�q�=���_>2>���=��2�t��>�J>t��K������4�?��@��??�ዿâϿKa/>;	=>�
>��T���2��JQ�)U^�X�_��T"?T�4���ʾ�iw>�	�=|]߾��þj'=,�.>��@='�G�X��ɏ=C߇��mA=�/O=6��>.0E>���=�<�����=�]�=��=<�S>c�9Qe#�{���	�<U��=Lg>��)>���>`�?�0?�}d?�)�>��l��Ͼ�����>Ƥ�=sk�>$L�=@�?>E��>&�7?�E?�L?��>˖�=С�>\=�>cZ,�`�m�@��嶦���<�x�?�Æ?�P�>�~}<b	@�H-�b�>��ʽ��?KY1?6�?��>��I῁��2���;h�l=���<��_�K	�6-��+Qa��=%��W�=��*>S�g>�8#>�iJ>{A�D�E=�7�>���=���=y5��g�f�%<�<�;��X2@>�R>�6���=|j>�4����#���=s+�=���`ļ�;��2C�=���>���= x�>K��=K���ܓ6>��y�T�H�`Ӆ=�Թ���A���g�G�z��=)�����s%>��J>c��U4����?*I>��J>���?l�s?�
><}	���ȾP{���d�[V�q²=���=
�W��>�.�d�c`P�ݾ���>I�>�
�>�>n>L�+��?��uq=���s�3��0�>+Ɖ����I����q�<��[��r�h�0,���D?쇿p��=�W~?��H?��?�	�>����n%ؾ��/>3���=��<(���s�-���?��&?��>G��,�D��z¾�T˽=�?ā>w�>���Nc��m����/�8I�>QQ޾�Eﾲ�*��ヿ�W����?��5��&��>j?�h�?�X��-X���4��:ھڗ���9�>B�2?׎>n)?ѡ?Ƿ�տž�7�r�O>Me�?nJ�?T��?S,��	U�=����s�>��>�h�?�ߓ?��o?�D����>=���3>���)>���=�"�=~̥=�J?�?v�?�[����w���羟�K�<�=p�l=�d�>�l�>�j>h��=���<��=�ig>�g�>Q^�>lSo>/�>��>����Y9��z?���=�>�>-1?�"j>y�=�����nX=�ӷ� "L�׮B������qȽ~O<4-���!=tf��i��>X6Ŀ��?��E>�	� ?���z�c�a�I>��s>���i��>��G> �>��>2ԝ>��%>-�>�!>�YӾ&V>n��J!��(C�R�R�[�Ѿ�y>�!���c%�B��t{��o�I�����ґ��!j��=���y=���<�:�?����?xk�z�)�(Q���?��>�6?�������	u>���>vf�>��l}���Í��(ᾛ�?Z��?�>�i�>��;?TO?�4������.�A��D��n3��Ge���y�H��(־H�H�d?7;�?�F?��>5�o>��h?��EH���D>�E���8��N�<���>D�����=qpo�r����D�����?��?Eٗ?�=-?.���(���ʯ>��3?��>���?G�I?(��>�<�|K?��'>Xj?�v?[>A?�t>���>-D>�e��h�>@=~\6<6�f��� ���۽�|�xX�=loi=��쐽��=l�J� .0�S� �߯�<�O�����OA��=zM�=I��>R}]?ä�>훆>�6?�;��]8���� /?��=���!����\���'��a >ˠk?\	�?gpZ?��e>��A�*'B���>���>�y&>H)_>�Ӯ>t�� P@��(�=͐>��>p�=�%V������	�����f�<�P>G�?
oC>l[M�>��������x��QI|>��<nQ���yx��j�E�1��jվ��>�E?�%'?��;<����+>�*e���.?�F?��Q?��??�(>!@оt!��B�S����>�V�=�+��Ү�􍦿��;��rB�5`�=馱�@���Z8`>�
�L�޾�m�GvJ���澯�W=+���[=i�Wkվ�]}��L�=��>����!�e��_-���sI?7l=0N���`Q�AԹ�<�>��>ܮ>2C�w�f��.@�%٭��i�=	��>��7>�۬�\���H��n�׮z>��H?�s[?紂?q�d��i�O�C��G���+��,���?�B�>�?��5>�� =UAþ�d���`��!8����>��>�!���A�ߌ¾-��2%7����>�$?�>Ny*?�+b?��>��L?�s"?���>qa>�����ћ��D&?_��?l�=.�սI*T��u8��9F�@��>��)?D�E�>��?<�?��&?��P?�n?��>O� �~~@�<C�>��>��W�cL��	�`>ʍJ?S��>��X?W��?C�=>��5�Sh��������=<f>љ2?�m#?7�?��>v��>R�����g=^�>�Mb?9��?��q?���=��?�4>��>�5�=�y�>���>�C?��K?��p?8-K?ݐ�>��<��Ž�����w���M��1�J<\Qj<�[t=F���ꅽ�&&��&�<i2���3���Č���ɼcdF��k�����;�H�>Υs>㾕��71>Až�$���A>[����S���㊾�+;��6�=�(�>h�?���>m#�(�=%|�>�^�>���D(?��?"K?�,;K�b�?۾o1L���>P�A?��=�l�����u��uh=��m?��^?.W�l���%~[?�ds?rp�w�,�﮴�.Sܽm���A?��?�/���� ?mc�?��r?�ܽ>zuξxo]����B�j��C���|�=A��>W�.��j�;�>��M?z��>��>-5�>����釿|�d�?�?]�?���?$і>�hG���ڿ	��Ƥ��9�X?��>��ƾH�?��T=g�о7��K���{�����媾����k��cj,��ц��%���=�:?&^q?�;^?���?��-0X��N� ��ZCb���j��WJ7���G��% �k7_����ʛ��o؁���@>Edu��=�ov�?KT?5�C�dn�>� �����ľ�0A>ھ�����"Zo=x\����K=]4&=>�n��(I������3?%��>n�><�O?��a�L�8�{Z(�i�J�'��K�	>A��>fb�>�&�>T��<G�9�߿�ۯ���l���)��6v>yc?�K?j�n?Jl��*1������!�0�/�oc����B>�l>��>ܰW�$��G:&�(Y>���r�����w����	�K�~=\�2?�(�>ʲ�>�O�?�?u{	��j��7kx��1���<1�> i?S@�>*�>�н�� �ƥ�>�l?���>��>�K��bB!���{�,�ʽ;O�>�­>.��>�Mp>�1,�@\��a��	~��19��Z�=��h?�����`�;�>�R?��:n�E<Ft�>��v���!����q�'��>��?���==x;>�{ž�*���{�����)?�"?3Œ���*���~>�"?��>�>� �?�֛>��þp���i?K|^?��I?]�@?@t�>=����Ƚ��&� �.=jm�>�:Z>~Ln=J��=lJ�$�Z�9��0E=_5�=3,ʼ����<�Ǽ�5mB<_�<�,4>_B߿�UC���;J���R����>��!�н�!��/� ������X��;6�&!1��?��u�f�\-��h����+^��A�?˘�?��o��U-�1���~#��d���>��-��>����$�O2����ھ ���I:�5�H��{�K�T�O�'?�����ǿ򰡿�:ܾ5! ?�A ?9�y?��6�"���8�� >LC�<-����뾭����οC�����^?���>��/��s��>ڥ�>�X>�Hq>����螾l1�<��?7�-?��>Îr�0�ɿb����¤<���?0�@CyA?�(���MoT=���>��	?�1?>y>1����(��kZ�>J�?���?�M=��W���
��Te?��;�G�=�㻜@�=� �=.�=�d�MJ>+\�>Z��[^@��V۽W34>�ʅ>=5"�9t���]��<n�]>k�Խw𔽐��?*��"n���T-�bwx�"�q=L1F?`]?� E��s$?m��v�¿; \����?'�?K�?3�?�ʹ��V�������Cg?t�:?���=��1���a��=ȖE�
(O�{˩���v���=E��>���>��E��\�u�@� ����>�(���ſ6$�#�C��<�"��`����rT��<xS��О�v�k��ݽ��Y=p��=-ZN>.�>?�S>M�Y>|EW?a�k?�r�>=�>����'��-; �-�W�����vw������A���쾣P�o��x�o����Ǿ�=��W�=��Q�栐�|� ��b�YXF�i/?o+$>��ʾ,�M�t}'<R�ʾ������Q��"̾F�1��n����?�A?zۅ���V����Đ�D����W?yb����tǬ���=�^��x=Lќ>{��=��⾞$3�euS�q.?4%?�Ⱦ�����A>a(�6�Y<wH(?R ?6��;n�>[�-?
�kh�_E>7>b�>���>�z�=V����׽�<!?�P?�^׽�d�����>�3����n�z��=KJ>b�8��꒼�{A>�U2=S;���*����d�4~n=r(W?A��>��)���`������T==k�x?-�?�-�>]{k?3�B?�ߤ<�g��x�S���_w=��W?�)i?��>�����о/���@�5?��e?��N>kbh�s����.�-U�y$?��n?�^?9w���v}�\��!���n6?v�w?��`����J���e�b�>��>u'�>�:�ˆ�>��<?e�.�#'���c���H2�/N�?mF@6��?pW<,ۼ�:N=i|�>�i�>�L5�����ʔ��.Ը����=ْ�>�ؤ�Ap�Q"�C .�	�??�Ä?���>F������]��=tF����?x�?	���� i<����k�^_��f�<�a�=ٍ�E�,��%8�Z:Ǿ��E���>��u��>n@��n��>�9�����UϿǅ�*�ξ��m��?�A�>�$ɽIC��Gj�8Ou��$H�7FH�S�����>���=Td�������2F=��SR�v{�>��T�	��>��E�?����������;u�>K��>���>�c������!�?b�� ѿ�C��T}��]?\�?|��?�?(��<'�n��Q��M�=<!^??hNq?�zd?'�׼��A��z�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.���_?�a�t�p�f�-���ƽ4ܡ>E�0�d\��N�����Xe����Ay����?M^�?w�?��� #��5%?��>۝��8Ǿ"�<��>�'�>+)N>e@_�q�u>����:�h	>w��?�~�?3j?���������S>��}?O�>��?�䌼��~>��>2�B��w'��:>��?Z���I�?%��?�?�x�Zv���/��qD���"�@�¾"aG��"V>�^r?]}I?+�>�"��g���AO����Ŋ=dP<���=��&�4J�>c- >cK��0��5�-���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�gf?,��\�� ,����=�)�i�jo�>��2?D��?ſ>��>�+�_A\�w��A�x�[�>A��?9��?4��>#��?����kD��%���9Q<>WH�?�~A?�1��#Y���q>�0�>��P^�
���t?�T@���?�j?Z4���yտ����n���<��U�=k'�= 4K>�ѽZ��=ah=�k<�cU�G�%>k��>E>�%Y>%$>7E>|9>����'�Qx��&4��dVC�g����G�k�9�	�evO�(U�}$�� 'о4�ֽ�����ڽ-�t��j?�(�x���=߬U?�R? p?ΐ ?�zx�֓>����P=��#�l˄=�0�>th2?��L?&�*?�ϓ=����	�d�`��B���Ƈ�w��>�nI>��> G�>W#�>DWO9<�I>�2?>Q��>� >�f'=b_�Cf=h�N>&J�>��>H{�>�B<>�>�δ��1����h��	w�/̽��?ۀ����J��1��G:��+����f�=+b.?E{>����>пN���(2H?�����(���+��>r�0?BcW?��>S��J�T�F:>��ݤj��^>�, �N�l�K�)��#Q>.l?�>|��=À���X��:�����o�>C�r?W������v���C�����>dc�>mkǼ�h�Q���ހ�s�Q��z�=�"?�?�@�RQI�T@��㟾�+f> �G>.5A=�-�=8eo>����U�2�:����,����Y<y�G>\!?!+>�y�=�Т>9䙾n�O���>"{C>G+>��??do$?���W왽3����,��w>��>�À>R6>lK�Ry�=�J�>!.a>���炽e��"�<���X>�^��_�)	{�/{}=7S���D�=Q�=����=���"=�~?���(䈿��e���lD?S+?\ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��L��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�/)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾLh�>{x��Z�������u�^�#=R��>�8H?�V����O�i>��v
?�?�^�੤���ȿ5|v����>X�?���?g�m��A���@����>:��?�gY?roi>�g۾;`Z����>ѻ@?�R?�>�9�~�'���?�޶?֯�?�<8>�~�?�p?k��>]榼}b'�q������\*=Fp�b��>��=����YB>�<m���͆��i�x;���T>��=>��>z���ž)-�=�����"��ڃ�Rؾ>i�x>!�>���>I��>C�>��>���;&����v������G?��?J`(���k�&��=�>� ��;>�>ɬS?<�������\�>�a?�mp?�'?�`N>w�����ʮ��P������<�gJ>�y�>Ș�>�� ���`>(2ɾ��B�>�j`>����xƾ��l�o!�=�]q>3�&?�U�>�>��?r�2?6\>��>�uL�������c��K�>���>N�?��?��?H胾Ց2�6����W��n�n���=~t?="?�
�>�p��\��龤�B��PQ���gu?��w?�k�ŀ
?g|�?�U-?ԛ?���=����z���8��u">*�?I=��>�)z(���
�m%?��?ϥ�>j͐���ѽa��1c��i����?��[?��$?̭�	�`�Y�ž��<l8�}���]w4<�k�C >��>������=��>���=W'm�v0���<���=zč>{N�=�<�7쐽��+?5���߀���=h�q���B�Iy>�E>�zþ1|\?��C��	{�s��6'��xQ��&�?���?���?���7h�/1<?�ȇ?�~?'D�> ����ؾoG޾��v�uuq���/p >�>M3������w��u��}��������Iy?ߌ�>=�'?���>[�R>� �>�~��|�'�7�����Q� ��#)��%+�ui�|���p�[���<�d�ʾ�0��/v>�5�|��>`��>��g>�i>�r�>��ܽK��>Na1>�>ײ�>A�=�X�=��qV�o���JR?����P�'�C�辕���^3B?nld?�,�>ʫh�2�������?U��?�q�?I-v>~h��*+�\l?5�>���;o
?�i:=e��bf�<�W��ε�0�� ����>�E׽�:�9M��of�l
?�,?@S�̾�!׽�ծ�Ti�=�&�?�(?�����M���c��I��nL��N��S�7�����b���b����o������dB-��U�=�)?�|?�*�ED澙�ξ�=h��I��j>�M�>��>gE�>q:�>��	��)��nK��7-������|�>�aw?�|�>��I? �;?u�P?=TL?Ϳ�>��>�J���"�>�y�;v��>���>h�9?��-?�0?WY?z+?�&c>E���L��Wؾ|?X�?�/?0�?�?}���$1ý�Q��+j�Ѿy�u5}���=ڽ�<B�ؽ�Ew��UR=�T>Do?���ɂ7�����4g>��A?�R�>��>(1y�~�n��=���>�?�h�>�����l���
�ͣ�>�ǀ?㻼�j�;��!>O�=�t��4�<M�=<ȼ�ۋ=��?�6�,�ha�;ٲ�={Ix=L�1��^<��Z�N����ީ<6-�>}�?^�>ӣ>���� �����X�b=f�*>��;>���=Жپ~ ��F���ܧ]�ўq>-ʑ?�ԯ?�ć=�h�=��=�]��ߪ���	��ż��ؔ=��?�f?4T?�?�=4?��9?-��=p�4`��*�����͖?� ,?��>���P�ʾ;���3� �?�[?);a�ʶ��;)��¾��ԽK�>�Z/�t.~�(��~D� g������w��%��?���?6:A�b�6�gv������]��L�C?@ �>�Y�>3�>��)��g�.$��5;>���>JR?2�>��O?�{?��[?t�T>�h8�m@���ҙ�p�5���>��??̌�?⥎?}#y?˹�>-w>��(��߾�m��:�g�ق���S=q�Z>�.�>���>h-�>w��=��ǽ�����">�F��=��a>a��>�U�>�>Ux>aҦ<��G?$��>W������᤾��j=�U�u?���?�+?�3=b��N�E�Q@���Q�>�m�?���?�4*?W�S����=q�ּ�޶�K�q���>�׹>5�>Oғ=F=oz>��>p��>8��d�up8��M���?F?���=�UοfF�P�z�?�(��!��q��\�>�wSɽ�1���K�>�򰾢����w���;�ؾ��Ǿ�Z���= �R��/Z?ю_<��>"k>�uD<J�1=��=}>_ȋ���,>��m�B�4�/_��˼W��6���-n=_�;U�>�̾]��?A�F?�q ?��f?)��>��=tH�]K�>5!��K?k՞>x�=��7a$����0��+�¾�ǿ�@Au�uT����>>#ӿ��\�=;$>)a>N=�6�=N,�=
=𵽥�#=�Ӳ="L�=�ϱ=���=-�>��=�/�?���ˀ���wG�c�ǨZ? x ?� =|Oξ��Q?��|>����)ѭ���%�V��?T�@���?h�L?ݱ��<�>��&���� r>X�=>G�>;�4��ռ�T�>�M�;�ƾ߾n�[K~����?�@?ߴ��(Cο"���2>���=N^N��~4�~|S���`�ñS���&?۱8�7"ɾskz>�=��ྂWľd�L=}�3>� E=&����\���=��y���C=*x=6k�>qcH>�R�=�p�����=��Y=��=ڹH>�9;%kW���>� �=}��=�2V>�� >�?�>;?�/?�Sf?[ �>��g��۾�Ⱦ�V�>�,w=�M�>��s=U�%>B+�>89?�6E?y�L?-+�>d�c=kj�>)��>��*��Mm�a�ؾ����Na<�@�?&��?K~�>G�<�2�U��<�=����>�?��0?��	?`�>����ܿ�1'���7��?Խ`w <�=\
-�15Ҽ<x������?���|
>,}�>��>^s�>�C>�\f>�a>���>C�>$6�<Xd$=zN��1`�<_ö�>3�=�8���<�J{<�d�<��=��4���C��"<��";�:�;LE;��=2��>TR>�9�>z�b=%H��y�>f��N�L�^�=�̾.�;��eL��s�I�%���>�A�m>��(>�3�U����?��P>ѳ>���?�^?�:[>=}��*���bE��bTF��R��r>��>�㑾�;�r�o�y�P��J̾G��>:ߎ>H�>"�l>�,�#?���w=��Ob5�$�>}�����)��9q�@������8i��Һ�D?�F�����=="~?7�I?A�?���>c��1�ؾ�:0>TI����=c��*q��g����?%'?
��>z�W�D�Av�4	$��g	?S0��a;����r)��=U@�s?pGɾ��߾��!���|��Y���V�j�ٽ�e�>J��?� �?y����h��fC��v�m�Ľ���>bX3?`��>R��>V�$?𦙾9�	��׽W]k=Us?�j�?��?*j��[�=���e�>��?榕?���?��v?c�Q���>F�E<�U$>h�a�9Z>�>"8�=wZ�=�	?��?25?l����	����ojh���8=ƾ�=Ƹ�>�>�[>E{�= �/=��{=��U>X�>�Q�>>�`>熣>��>�,���|���&?���=�v�>�/2?߸�>��e=���Jw�<�aP�1�?�S�+�䕹��i߽�^�<m���H=U�ܼ��>�ǿ��?��W>e���?D;�:EC� �Q>|T><޽�,�>G?E>�}>E[�>X��>@ >Fh�>��)>�Z�N�>�n��G�<��TW��߽��g�>k���W�۽gz�a��9<��]ľZ_��sn�(-����E�y�=�4�?��J�]�-�&�J���?��>8�6?m��h����b�=H��>�Aw>>�꾔_���Ӌ���ľ~r�?|��?�ko>!$�>)�I?7W?�Z��o.�cuT�j6��V�"�9ӆ���^�H�z�C����Z�I�=��V?#6j?��?2�/>�=N>V�q?m	�qý��>����=~���1<�S>��%��c;������k<"�>bb?�v?:�?뗜�.s�"�>6�?-?0�y?%NJ?��>?X(���:?'�>g�?�A?�/]?L!?R��>�I�zQ�]_O>TB)>�T#�zwϾ<�"]6�ѻ��F�0>A�>���=|�<�e/�D�8<��4��\w����w̐=���=k�-��J�<���=���>'`E?���>3x�>��3?=���^`��)ݾ �>��������&��w������T�>�{W?Ü�?3�V?�S=�T2�P�����>ۏ�>�m�<�X>��>0=��9׾B��>� ټ ��=E��>c���{�����F'�T���a>7e�>�%e=�ŵ��ƽ)����ݨ��{�>�r_��ؾJ�ڽV`���"�΂���?�K\?$h*?y�=g�Ⱦ�Ľ�r�*�??S�S?A?���?*�l>�Nɾ��Ҿ ���	]�M�>Y=�=���~`���c��P�C��Ԩ�N?Q>^Q�����#Q/>�&�Z�V�!WN�[��E���"���(��-�=�u�"���&(�r�:=��m��a辬(1��雿�_׿��E?�l>ҭ��8���2�����>{��>gYu>�m<��BU=;58���@�Z��*6W>�mT�M��@IݾժF�!fϾ��>�E?$�_?x9�?4����q�H0B�����.O���N���?n��>"�?�?B>�h�=m��`��Z�c�T�F�M��>��>3H��}G�2柾������$���>�B?�q>v�?_�S?� ?�1`? �)?�?��>�9��a���B&?r��?��=&�Խ��T���8�FF�:�>��)?�B�a��>��?��?X�&?F�Q?9�?.�>� ��A@����>Z�>@�W��a���`>�J?4��>n:Y?�Ӄ?��=>�5�颾/ϩ��M�=,>��2?�6#?��?���>ؐ�>����(E�=���>�c?5�?��o?3}�=X�?{�2>��>
(�=�ӟ>�z�>�?�3O?��s?��J?�b�>6�<�������Ss�MGS�3�v;�D<��x=�����s��t�e��<��;���ߝ�~x�vYD�������;�a�>��s>zᕾ�1>��ľ�q���CA>�����a���ފ�-;��I�=QZ�>#�?O��>t@#�=��=ߓ�>9<�>��O(?��?�&?��;��b��ھ0jL�tְ>��A?x0�=��l�����u�zh=�m?��^?PW�����k?WjX?����AP������y���YW?��(?RҾhA�>b�?RWV?3�?�Y��ʀc�wI��|k���y��:>3V�>X�3��w�<�>�I4?_v;>���>�>�-޾������q�E��>Eـ?
��?1��?�6'>�9����㿟�Ծ拿�_?s��>nS����?��=��������y��2�d�¾�q���Ϡ��������
���<1����=�5?��~?O?4Vn?����Qk�YA��W����_�������'�z>�bE�[GY�"��50��1e!��k=(�Y�mT&�R�?1?�ծ��3?��e��� �~Ք�v�>v���"J��>��3��5�=��<����w�������I|?u��>�˽>�	'?MV^��7C��'��N�����=]>4A�>=��>!(?�:<�QA�*�?ߛ�~�C���/?v>||c?_�K?ƶn?�Y��%1������!�l�.��j����B>E�>Vȉ>b�W�	��Q6&��U>�h�r����G����	��A=F�2?�K�>D��>M�?i?lw	�_e��PXx��~1�د�<�=�>�i?�7�>�Ն>нn� �S^�>t&k?(��>e��>�������x��ԽԵ�>d�>�U�>�o>	4��t[�@g��2���j/.��>`f?C���X:S��6�>�U?6��<�6�9�T�>�<F�u&��v����g�=O?
��=`�B>U˾�����w�荾z�(?p]?�'���E*�?̀>�!?T[�>��>�.�?�k�>?�¾#�9��?�j^?5J?��@?%z�>"�=�̰���ȽsZ'�XE0=Ц�>5Z> �k=���=w ��K]��M���B=���=�Ѽb1����<�Ұ��H<��=>e4>��ڿ�L������m�Ip۾��-���+H;�F��\Ҫ��R��p"����&��Ľ)Ľey���z�ۅ�������b�?�F�?$j5��C���ȍ{�`C׾�[�>Vq�����]V���9���X�澊�����
��W�5m��ɉ�r�'?������ǿ����5ܾ�& ?jB ?M�y?��"�0�8�� >��<&���>�������οQ�����^?T��>�E�����>���>��X>i8q>����O%�<Q�?��-?׉�>�r�>�ɿ�����z�<'��?��@�tA?��(����9�Y=�x�>�	?��?>%�1��C�����_�>,�?}݊?#�K=��W��,�g�e?>�
<�F���廰w�=��=�J=�[��J>���>���fRB���ܽ� 5>[��>�:��t�^���<�\>H�ս-H���#�?��h������8lf�/5�>c?�q`?-���Q?��꾜 ǿ�(��N�?��?2��?`wP?T������=�.��t7?�QM?�->����������=��
>s�us����[�W�*=���>%O�>�)������G噾zi�>Q=���ƿ_���7���>=N��E"�rzC�CI��T���P�.W��f>�C�=�_�=:݀>��Y>�_>��Q?Ge�?wS�>�9�>Ud�aj���پ~(��S���q.�wM���
�^��Z���L �����Z�H�J(=�Gҍ=9#R�T���B� ���b�}�F�B�.?L$>��ʾI�M��u-<�Wʾf����L������5̾(�1��.n�[ǟ?��A?C셿�V����~P��S��c�W?5N�����ାs]�=̬��F=�>��=���g 3��S�$<0?9=1?D�ϾIt��5��=���Y���+?cu'?v�����>X`+?�R���	�/>_	>��>Uh�>,�=��̾�&��12?��r?͌�<<����>�5���hW�n=�N>�Oh���/<�$a>4@�=<9���@w�t�=���=y$W?���>��)����m��g��5.==x�x?ǅ?��>^wk?��B?��<�k����S��'�my=�W?S#i?˘>�I��3 оGI��#�5?�e?�O>k/h�� �=�.�uG�7?��n?�Y?7^���z}�n$��{���X6?k�v?�m^�������	rW���>���>���>&�9��γ>Z{>?4a#��L������74�eҞ?W�@���?�@<���(�=�?+k�>~!O�v�ž�u��2~��J�r=,��><���Nv�� ��,�/�8?B��?��>ފ�������=׋��GQ�?���?���{<<��Ll�*����9�<�=TX��W���$�7�m�ƾ{�
����~ļЕ�>�A@F�罗��>gO9��s#Ͽ�(��q�о�q��?8��>=�½�k����j�_u�OGG��rH�VC���t�>u��=n��A���S���1@��%<>���>;Q����>\��i��4+¾V��G�@>���>�/�>[�=�����?�?���n���J���,���?'�?-4�?�lC?��>�����x������?�F�?���?���^�.�	�=�j?�_��oU`��4�sHE��U>�"3?�B�>Z�-�G�|=�>r��>�f>�#/�z�Ŀ�ٶ�"���W��?߉�?�o���>o��?ls+?�i�8���[����*���+��<A?�2>���G�!�60=�@Ғ���
?O~0?�z�b.�:�_?��a���p�P�-���ƽ-ޡ>��0�TZ\�x��x���Te���Oy�S��?�^�?��?թ�*�"�3%?m�>K����3Ǿ�7�<l��>�%�>�$N>v�^���u>����:��f	>?��?V�?�h?����o���E>��}?@B�>/��?'��=ޭ?p~d>>���&�9�>�>�y�>�S�G�?��U?9z?\�<>t�ܽ�|��l;��9�Ghھ��D��{�>�fl?�BC?��?K�V�y�<�
������i&���H<w"����;��=Wˏ>+�">��U<�Fx�˗���?Ip��ؿ�i��Jp'��54?0��>��?;��p�t�6���;_?z�>7�,���%��PB�X��?�G�?>�?��׾?P̼_>	�>�I�>p�Խ^���|�����7>T�B?���D��?�o���>���?�@�ծ?Ki��?�g�1Y��R�����0c��<}>P�6?!{���+�>qa�>��p<�Gw�w
��2'd����>�f�?u��?/��>B%t?t�i��_��=�
�>��h?X�
?��1<�����X�>���>+��H���d@�G�|?��@�M@��W?����0�ڿz9���þ��9>��=0�=VJy�~��<���=+�;v=�1E>��>ů3>�U#>]�0>�C>�#>:Є��+��뙿����WM<����g\��go�/�%� ������%?q���3�[���������H�p��=+c?TN?-i? O?SzS�tv�=��Ǿ�J*>KS�,��=6�>�:?8UT?�0?��^=M���`�� l�;̩���t���>xj�=۳�>���>�}�>���;U2>�BL>�wi>n��=D��=N�*�U\�=�Q>*Y�>���>�ȫ>�I<>#�>ϴ��1��ٜh�� w��(̽� �?|���J��1��5�����.y�=!a.?�z>����?пH����0H?�����)�w�+���>��0?�`W?�>���q�T��1>���t�j�v`>) �y{l�W�)��%Q>7i?jc�>|��=+A �j<6�av5��'���D�>uG?���#�v�}�U2N��%��J>��>�k=�5����?Ra�"�Y�a�=��1?��>���锾<.��5�֌>��>ޮ��G���V9>Y���e��p�Q��Ӈ��k�=��V>�?G�>�l�=�>�����]�N˯>HYb>�?!>w:?F�?��>�f���������#�V�y>Dy�>��g>�>,�L��Л=A�>�O>b�伶�&�ۊ��G@�N+y><���a�R�>�{�p�=o������=)�x=�)��F�A��<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�g�>�x�TZ��-��=�u���#=���>�7H?ZW��"�O��	>�v
?�?�_������ȿ�{v����>��?���?H�m�UA���@�A��>��?gY?!oi>h۾�_Z�{��>z�@?�R?��>�9�&�'��?߶?�?I>���?��s?���>ֲt��0/����A�����}=�t;T�>�n>G����fF�Dʓ�;c����j�Č�>b>�%=�ȸ>��㽇G����=����C;��&f��ѷ>#�p>�PJ>��>�� ?��>S%�>F�=u���t݀�:���-U?)@�?XSC� (�����/>���$,	?,�]?�B���߾p1?;mJ?�ry?�^+?��V>=�	�������_4ľ0�>#}g>a�>2��>@懾*ڤ=�־@��N�>c�>졼�	�j��!Ӿ M.����>mD?z�1?�>���2?�Z'?��R>>�>�J4��c��Y)��n�>L��>xQ�>'��?c�$?���ʋ���"y����^�@�5>���?��9?]F,>a-�����:���3�Wؒ��ǉ?�Ŗ?�y�=}�1?�S�?
J?}CU?��>#{�����&���>�K?��6���$��4'������>��?H�?y��j1�|9ܽN��v��D� ?��K?� ?(O��jm����u�<�RQ��%=Mwu�3�R;I=M>��=0H���=u�M>N=n���P�9�~p<��]=ݽ>Y<
=�$X��J���X+?��ݻ,6�����=��p���@��W>L�L>E�þ�HW?_?6�6eu�VF���e��_\`��H�?ix�?tU�?M��If���:?)�?c"?b��>=��IѾ��Ӿ������ʕ
�!��=�c�>�u���޾���(;���~���Q��=�����>���>�N1?��>�̗>Ş�>Ѿ��A�8v�V����^����mb��c�˿8�2��������2��d�Z������9�>��=�[�>�� ?`�=>,�>:�>�؞�$l�>�>��< ا> �+=���<D��=��y>�Wd>3LR?�����'�D�辎����3B?mod?22�>��h�O�����%�?,��?cs�?y<v>&~h�L-+�,k?Z=�>t���q
?�E:=V�=b�<;V������7��)�>oM׽�:��M�Clf�Hj
?p/?X䍼D�̾(E׽����sk=�s�?�+?��&�rS��&e��9Y���V��@м����λ�	���n��Y��x��Tу�� 2��bg�j�-?q�?=Z���$˩�.UO�t�*�OkS>���>��>Dq�>��/>9��+2�]�T�#���v�`�>	A|?鋍>��M?��7?z�N?JP?+�>�>����j?�H��F�>���>=?�G-?�b/?m?V�?� Y>~׽����^̾.�?*v?f�$?c(�>��?��t��P½5�]��c�>wd�=�}�lY�=30D=��Ľ�]��T=6\>rX?�����8�����k>j�7?��>Q��>Q���-��#��<�
�>.�
?�D�>�  �c|r��b�R�>���?N���u==�)>��=I����Ѻ>T�=������=r���u;��<�|�= ��=��t�
ς����:��;jq�<��?K?�mj>��>?O��P|���������8>��]=��=������(���Rav�3C>�Z�?t�?rK>뵅=�r��UE��s����޾"���S�=Z?���>j�4?u��?�=?�F?i�T>2�����"l�f)�J�>� ,?ʆ�>��E�ʾg�L�3���?�[?W;a�R��!=)��¾�ս��>�Z/��,~����tD��셻w��;x�����?}��?�0A���6�r�6����_����C?��>mW�>
�><�)��g��$�5;>��>�R?�9�>ߗN?O�|?b�X?ރX>��0������F��	_��^w;>�QE?\�?|�?�Zv?���>{Q>�W0���о���c�������èQ=��W>F-�>(P�><�>�f�=��!�Ľ��,��	�=��c>;	�>k�>f��>��q><=�-G?�8�>�[�����~����h��H��i&i?7��?��#?��;����#K���Q��>��?�G�?�&?ٞ+�vC�=a��:����q�6�>C��>�L�>|�=@7�=\�(>"]�>��>����� �>�٫~�^�?��E?�g�=��Ŀ>�i�mc;��ǔ�f:DΪ�a������s�짌=g������X����rN�@O��N���؎���/�����a�>E>\�!>�{
>�8;R�۽|x9=�VD=\e����;�V�W�(�����.�ͼ�����ڻl�ڔ�<�Rؽ&�����v?��E?�W?3�R?��[>P{�=���^6�>h�����?�ƅ>L4K=3����	�����s��9���%���a�O�@gվIN�=�@+���p=V!9>�h�=����IF�]�;>��=�\H���<���=�=�==�&�=|��=�]�=₁?�Lz��e��UF��>���&?mP ?Y*>ө۾��x?x�:>�Ɔ�&�ſ	f�R��?pR@)��?H6?�1:�g�>��!�9���>�x>���>�Pd��2���>I�ֽ�¾8��������a�?@�l/?ݛZ�d��� ��۸8>�2>�bQ��h1��	\�Db�4�W��h"?�:�
;�h�>6г=��߾�Kƾ�-,=��6>��Z=�>���[���=Ú�.�B=tc=<��>eMG>�*�=9�����=�:L=R��='�J>
����6�7e4�@�/=���=�R_>��$>��>�%?00?��c?ᱸ>��n�z�Ͼx�¾[��>T��=t��>ǃ=�=>�¶>p�7?t�D?�]L?9��>��=4ź>)�>M�+�L�m����hҥ�$��<%w�?��?:P�>�Ƃ<�?�T4�Y�=�=>˽�:? �1?�B?|l�>�W��i��G!�:|�\�(=<=�=��<�������ʽs�=�߽m���7o>�J�>���>�Og>ɀH>
3�>��>�\�>�4>��Z=�;��������<����fĵ=�g�  �3|e<W����鿽SH�<*�Z��s��o�<#��0#�Q�!>���>�v�=g(?){=����A>�����M�|!=���*^)���M�.vw��+1�߂��'��>��>�\���9����?kH�>��L>2_�?��:?��B>�v��8Kʾh}��1���া�ц>�4=�u���F�������=�I�ľ���>�ߎ>��>~�l>Z,�A!?���w=E�c5��
�>�|��1��*,��9q��?��v���Ri��zϺ�D?\E�����=W ~?��I?�?8��>�����ؾ�/0>�M���=���"q�0n����?�'?)��>��5�D��)��W��U��>��F�@G���f�=�Ⱥ�����;�>��v������6������=AQ��V�����>��1?��?��F�+j��@Y�Y��Eq{���?��z?�s>��?�.?��!���	�!DԽT��>`k?v��?���?���=���=�������>Ue	?s��?���?g�r?��@��>l��;��">������=
>�a�=E��=?p?n�
?�l
?f���K	����=��*�`�L�<?Ǟ=��>w��>R�s>��=��|=x��=,P]>�%�>��>�6d>Wң>��>Q����J��&?�z�=�a�>D�2?�
�>�OG=����Q�<�X�f�D��3,���Ž���q��<�GU��#Q=A�μO�>[�ƿa�?�}O>,t���? d��E�$��cN>�pU>��ͽH��>�"@>��}>�ƭ>-/�>�f>��>v,>{��-�=�p��<㾝;���0��%���p�=�qԾё�7|3��%���)���%%��j��悿m�\���N�"ؐ?R_A��4��l%��b����A?o�>js?��r���P���<.`?��=)|�zz��cԅ���u���?��?%�>�@�>+v-?�?�R��c�Ҿ�C!��y����<��{�2ʛ��v��ݑ���7�r�;�V?��|?)?dl�=��^>�b�?��|W���">w˾��m�oT��a��>s���T�(�D?(�)�}fB��]�=Z�\?���?�?�y=��<2��>��]?P�>_��?��B?G�?Ơz���I?�@�>��;?R�L?�fc?��>�S?���<����:a�>�=�=�(^�8u��[��s˝<omM��n>?B�>НýO�Ҡ>T|��ؽ���Ddʽq�T��׆<+X\=�KC>�}=���>]�^?6P�>G�>��?Ņ��q;��?Ͼa�%?�*�9�4���΅��'̾G���T�=H�k?_�?P?sɢ>\�7�`W�{]�=�ʉ>�3>���>�(�>�==�d��0��=�Pz>�pX>��!>!���ӵ�0��~.�m��=md>C?��>Ք�v�>�7��3�׾�г>��,=�S�ӱ��9�[�:)4���¾/y�>��P?i�#?�Ib>����۹�p_���?0Y[?��'?��n?YA.>�Ͼ\+��2��^���N>�
f>����~,�������>H�*1�A�]>�Ź������=�=��T�D�����k�Wui�����H���U�0��d.>������w��).�lN���ܾ]�*��e�������<?$�~=���r�1�)YѾ�\�=L.�>D:�>��=T_���/�.����P=��j>�Z>a.�<O��wE�DLӾփ�>O9O?A�Q?;�z?ἄ���d���F��ľ56�GVA���	?�a�>��>:��=�����۾��A�'<l�&8��p?���>��,��!I�(��ٔ����(����>�V	?;e�><N)?F�?Kd6?$t?�?Z� ?��>)���0�*?�b�?s��^�`������O��eV���
?6�H?OZN�L�>��/?�� ?�,?C�?,�?��t=l�.��r#���>@�>Z�\�X����,;>�QH?E�>G�Q?�%�?��>�*�u�����[�>-�h>�*?thW?��=?���>lx�>Υ��="��>��c?oͅ?��k?���=Na?m7>�N�>���=Cפ>��>�?q�K?C<q?�5J?1��>/�v<�����[����K������<�H<��|=d�	�9~��YB�����<�kp�����ܻ
�ļ44�������<���>77n>�/��e->�ȿ����PJ>����G�����5|H�"ƽ=�z>�?[��>!5��6�=���>>��>9�?t(?A��>Q?�#�;�`��s�tf��>��=?Fc�=i�����s�M-a=ޱl?�^?^+M�+[���b?�^?�B���<�҅ľ#�a�+4�k�O?��
?N�H�Oe�>�?�q?���>��f��m�=	����b��]k�c�=�Ü>����\e�Ƥ�>��7?h��>Td>2��=�ھ>Dw�躟��D?b%�?!�?= �?P->�rn�%�߿��������]?b��>�&���n"?֥�޻Ͼ�������}��k*����������P�#�7�����׽(�=��?w6s?#�p?�`?� �R�c�t�]����V�`�������E�E�D�@C��}n��!��c��(똾Z�D=�
����=���?�$?M�E�f��>���L��>�ܾ�\N>`����1�b��=����i�"=��=��o�� K��ɾ,�?4�>|��>�B?UXY�g�:�k '���4��/��!�4>�\�>!L�>�B�>��U;>SA�����¾����x!��u>�c?b�K?��n?'����0��n���t!�7�*�vn����B>2�>垉>_�X�˷�T&�2L>��r���҉��6�	�-��=�2?9�>��>E=�?v�?�q	�]B��(�x�>h1����<
X�>g i?��>��>�Oнf� ����>�k?���>���>�_x�Dv�\���m�����>�_>5��>h�>�R�U%c�"0��/��g��L�+>�2\?<��ir�!ŕ>�&V?<I);��:�f�>�����u�۾J\]�ю�=�?�뷺��c>k����$�{�N���+?�f�>)���Z<-���>"?A�>`�>d��?��>s�Ͼ��<R"#?w�W???'g3?N��>��x=�6��@ʣ���I�%�=�rf>��T>��!>e&�=�b-��u��pڽ�ם=`u�=�a��ac��� <;)���]C<(�<��B>׼ݿm�A�Aܙ�=���Hؾ*A�����'�4�����?�I?�����';�X1��I,���*�nrH�����B���R�?Y��?�C;��-*�xK��wD�Zо֍�>~`��p�=�Z��IAL�T;�Cؾ��۾(��{J�}c����Ȕ'?����a�ǿ�����;ܾ�  ?�A ?�y?Y�&�"�[�8�� ><F�<�;�����Ț���οR���t�^?���>���/��2��>���>��X>wHq>��S鞾G(�<��?C�-?d��>N�r���ɿ����Ӥ<���?�@MC?x�*�:��:^�^�?1?m�*>$�r��v��䉾QS�>t`�?b�?��=�J���u�V?%,=ɉ4��;�:�=F=n>�~=��C�D��>Us>6���g|��ܪ�6��>Js>n���!��5�7�
ڱ<��S>��ɽ�L-���?>P��Bn��ܙ.�B`�Wd�>��?>�U?z{=S8g?�l����տ��M����?ъ�?ʹ?��?���)+>���.�f?~�*?�Nl>�c��g����]�Z�=����?�1&����>N`?���=�	��(Ⱦڽ�ϼ_�>n_��h�����`:���=Lw{��-'��Q���(�2���k����o�oM׽uա<�>�b>�܈>�{>�+Z>��X?Ji?�*�>�f>>Y���
����ھ'Ȍ�UЫ��D��0<�X�����ܾ
rξ)����� 9���Ӿ�=�?�=6R������ � �b���F��.?t$>�ʾ�M���,<xzʾV��� q���¥��/̾�1�tn�ȟ?:�A?f���}�V�d���Q����ұW?hC�ĸ�謾�r�=������=��>j�=���+ 3���S�.�(?KC? �ؾ㾀0�=O�ȼD+/�L->?�D?�m� ��>-�>?{���|���>���=Fv�>Jn�>���>\���అ�?�a]?�&>�z���!�>V���f<��G�>�\S<~�<s/�r!#>ɟ�i����V<7�H=&W?L��>4�)�K"�ٻ������<=kx?��?�>�k?�B?Tb�<������S�s�w�y=��W?�i? T>pт��Ͼ_c�� �5?i~e?��N>��h��龇u.�_V��?F�n?��?����KU}��꒿U��0/6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?t�;<��U��=�;?l\�> �O��>ƾ�z������1�q=�"�>���ev����R,�f�8?ݠ�?���>���������=_ٕ�%Z�?��?�����6g<��l�n��Xm�<���=h�T"�����7�
�ƾ��
������Ϳ����>=Z@tb�R-�>�C8��5�TϿ���}[оIVq���?��>ѤȽꛣ�a�j��Nu���G� �H�X���3��>^G�<��a�֋۾�a���)6��>]�?3��a@�>�����þ$�¾�>���r> ��>A��>|=���t�?����������!���n?᲻?��T?�.<?�x�>��l������Y6�}�L?Ѫ�?2�?��½g����>�j?}_��sU`�ߎ4�mHE��U>�"3?�B�>L�-���|=�>���>�f>�#/�y�Ŀ�ٶ����W��?���?�o�"��>n��?{s+?�i�8���[����*��+��<A?�2>
���@�!�H0=�AҒ���
??~0?8{�e.��^a?��d��eu��-�|fν5�>�j�*�L���ݼ��0�^�����V6���?J�?���?{	��y$�V=!?Ϋ�>\h��FȾ�/=��>n9�>C�I>- �їw>K�E�;��8�=E��?.��? �?>8���+��{q�=�y?��>H�?Y��=U�>&i�>#�{������uI>�G�>���;H<?�i?TQ�>�=�ڙ�9�#��+�i:-���̾?�L��l>}3�?%�d?l��>�l����ν�18����Q`�<T�=.[!���/=�ɽ+}[>^u�=�Op���'������?Np�4�ؿ�i��p'��54?,��>�?��{�t�[���;_?\z�>�6��+���%���B�_��?�G�?=�?��׾>R̼�>-�>�I�>F�Խ����[�����7>6�B?O��D��r�o��>���?	�@�ծ?ci���>ü
��Ig�}�y�������C>��G?�=�/R>�	?��7=��h�ڭ��Gu����>%t�??�?��>_|?Cg\�	HL����R��>)_?��$?�"<�����fU�>�?.�������ҾY�y? Q@�@<dN?�~��+�߿9&������߰��#��=aB�<�]>%Q@��<6c�<�A��R�]<��>��>��F>�^O>��:>V�z>�UJ>���	��9��������F����e�ya����cc�������B�����ڽ��ｃY����;�ӊ*���m����=K�U?*'R?0*p?�� ?�v�&X>.c��O�=��!���=G�>�}2?(HL?۝*?��=
����Xd��[��z������0�>KJ>���>���>۽�>�A���F>�=?>졀>- >�B(=T�=)�N>T�>ɸ�>3	�>�C<>d�>.ϴ��1��2�h��
w�+̽3�?q���D�J��1���9��.���Ui�=Hb.?^|>���?п@���t2H?&���<)�Ź+�/�>Y�0?�cW?Ӝ>���T�:>���j��`>�+ ��l���)��%Q>Kl?b�f>�>�=-����S��k������y�>C�b?�,��L^��D���F�X&���>H�>��=eQ�q֒�H/�p���w��,H?�;�>.�X�P���z?��ξƠ=��=�U�<}H%>���>���=He-���~�g�=�J>���=]J?b�+>%��=��>�Ϙ��N�=�>A>^�->�i??ı$?׻����������[-�
Xu>���>B��>�u>QoI�խ=A��>�%a>ȹ���肽!� �@���W>:y��1`��|w��{=x��ǥ�=@g�=����s1<� �!=�~?���%䈿�뾞d���lD?O+?) �=ܟF<��"�D ���H��H�?o�@m�?��	�ڢV�?�?�@�?����=}�>�֫>�ξޔL�۱?�Ž9Ǣ���	� )#�fS�?��?��/�Wʋ�9l�6>�^%?��Ӿ�a�>)���V�������u�E�#=%��>K8H?a����O�O>��o
?s?d����.�ȿ&~v���>=�?!��?��m��?���@�@�>���?�dY?��i>sk۾�eZ�폌>��@?�R?��>�9�g�'�s�?��?��?��4>jԐ?��n?5C�>���<��+��V�������w�=�����m>/r�=��ȾmJ��e���a����x����:>��l=�x�>/���o���{�;���_�����9;���>
ed>��G>kУ>�� ?�5�>�H�>�Q=�-�eԟ�]i��pK?w�?���{�s��p��M,�=��m���?��=?�����nƾ�>�6W?��?~^R?�-�>b"��ḿ�:��%��<;Y@>#��>Oy�>���{�r>�ʾm/����>C�>H��<0�+r���[v��Ӓ>�O%?vi�>��=5?�%?��o>+��>xC�PD���9F�X��>���>R�?��{?CB?�����;3�sՒ��E��}�_��;>�s?O!?�ɓ>1���Q���i�C�ix#�1��/G�?�f?%{Ľ�|?j�?�zC?
�C?EUf>����WϾm��>�|>+�?����e:���)����$�?��?���>Ǆ��� �g荽8���N�� ??��Y?;$?_.�Ƽ_����V	=B۶8���07�<����>y>*L��h�=F>�D�=BW�ZA(��`=<�=��>F��=�(��ソY5,?nD��ჾUx�=��r��gD��S>�L>s����^?)=��{�(
��w��ztU���?��?�h�?����$�h�<&=?�?i?��>�@���Y޾���u^w�#bx��w��>��>3gr���������F��<ƽZ�\8?	��>6�?X)?U@>d�z>�B������m�Q����TF����1J�\�3��-����������S�Ҿvgh�`˰>[@ݽ�D�>�'�>�C{>�8�>_��>H{O���4>���=��^>m�>a^�>wG>��ý��3�^P��;�Q?����&���MD���B?5hb?.	�>�HG�Kك���2 ?�6�?��?��s>R�f���)�]�?�G�>�[x��_?ĳC=Ѣ0�q�G<�ί�N�s����
��)�>��ǽ}�9��8M� �f���	?8f?�d`��rʾ� ѽ�f� �}�r�?
�A?��I���p�oJ��O=�f�d�f=����Sf��q#���y����s5{�{%��xZ�� `��g?�]?�Ծj�	������T:�����ן>e��>���=�>1>]7꾂��_mA�2! �Nˎ����>^�p?�X�>?sU?O�6?�ya?��S?�σ>�6�>�%���e?��	>iH�>Y�?�l7?��?�/?�.�>Pd�>zZ�>��ʽ=s����)��>И?��>/z�>�?���q|ɾ��v�-|*�%yQ�cٽ�1�=��+=���-��ٙ>$��>?���P@6�d��6_s>�i9?���>���>����Ɂ}��=h)�>��?%��>���I�q���!�>w%�?���a�<У*>F��=������;�r�=T¼H��=�>����"��%<m�=�i�=ӄ4�+�;�z:!�N;�<ۓ�>O�"?FgA>gN>]T�T/¾�{*�֯��1S>u��l@>�Ɛ�� ��W���Ɇ�nq�>��?��?&V=!@;;��*=����2x��o��8���>%=�Q?�n�>A�,?��?��A?�?'�<<zc��Z��:o��Aˣ���?�,?^��>���ɸʾ憎��3���?�^?�:a�f��m?)���¾�սq�>�W/��*~�����D�R�����"������?8��?>A���6�v�k���]��K�C?�>{\�>_�>h�)��g��$�q2;>֌�>�	R?��>��O?:{?��[?��T>��8���ƙ�� ,��">�@?c��?.�?��x?�{�>�{>�)���߾M`�� ��~�dЂ���W=e�Y>�k�>m:�>�ĩ>��=_�ǽ���8?�w��=�b>��>���>n��>kyw>qx�<�DG?���>k�����>��HBu��Nx�n=r?�?��&?f8�<���,�D�R��Gܼ>�T�?���?о'?d�C�(�=^���/�����v����>���>-r�>��=M؄=7->0��>:��>_Q�Pf�)�6��Y���?[sJ?h��=eY˿��Y���>֮ɼe"�D���P��A��^���!>�X��`#���0��5����է�V���2K��~�r?�W-=��+>��>�X4�ԍŽ�T!=��4=�⼽r��=es=���޽ȈU�~�����A��ȶ��j���c1�i��,���x�?�9M? 40?a�J?��>��>�B�8�>mռ؀?/�>�\�������	�ƍ������p¾�>���Z��ܬ�}t)>�u��N&�=W>��%>ᄼ"?<�׍=>>�=Il�;{|=k��=�8�=���=h��=�3>e1�=�͂?+9���:��>|v��ᾧ�^?z%+?�|>�����:�?_��>:������hE�BZ�?�~�?扱?9
�>K����?p	���u�r>�fY>Z�?�?B��	�#� ?0ܞ>�ߺ�{h����l����?y��?/�?��W�ͿCc��U�7>˿>��R�v�1�eS\�O�b�%�Y�
�!?�2;��`̾���>�W�=�P߾�Bƾ؝/=��6>��`=���`"\�X�=�\{���==��l=?w�>��C>�u�=����r�=��I=��=%P>I���5��,���2=e�=}c>�
&>D��>%�	?7�$?�\\?%�>"Jd��a��3¾�~�>PUK=m{�>R��=[�~>���>�/?�&:?��;?�B�>�	�=}�>�n>=.�ɳq�c|�����O��I+{?�1�?�>�ר��m�����b�8��ﱽrY?�1?���>�c>9���JϿ����f�/�I�|��c7���b����:��i�u4e�iq�����=�zY>�C�>�K�>�~k>�Й>'�d>+��>��0>��=�iQ=�<����W*u��/c=+�~���ݻ�tƽM�G�ɽ6A���թ=�_�=,b=����9�4B�=�#?pj>l�>rp�=Kݐ�k/h=�B���8�?������ ��jZ�j�����@�x[��ɈH>%�j>f��瞒�59?�C�>�>=>[��?��V?lb>�A���6��/F��F롾9~�����=�ݗ=�S��V
6�'�~�7sI������>6�>�>��m>g�+�9�>��ct=���>5��g�>�K��(��
z��[q��B��5���o�h��ݤ��[D?�H�����=�*~?7�I?0�?�N�>?���0^ؾ�K0>gE����
=<"�'�p��"���?�&?a��>�.�>�D��pξ6kW��1�>��"�ff�$e��/a��nI>����L>�V�������W��F/���M^������>{�8?1ץ?]�t��1_�:BI�@&꾄�/f�><+x?��>)��>�*?��V>��(���}->[w?�J�?-9�?�?�=��>��!-�>Tj�>���?�j�?�]?q��V�>�#��&V>��=I��>!Y>[�=�==�>�z?i?p�'�$�&Mо�z׾��p�<C�=֯=�z>��>Ja4>�� >�����k/�g>$��>�4�>��Z>k�>��>��;��	�5�?H�=��>,?肀>FX�|�=`�=N�Ž����|��=hZ��N���J����ջ���=^<x��>:������?2p=�ͪ�?�?}|��-�<�>��>��E�iH�>B$�>�e>�Í>�>�@>�V>3�.=��,�=��Hq�y�U�5Y�ِ��0v>J���*�� �o�����@�����|y�����+C��Vu�牉?q�%���W�j0*���˽�"?^�>z:J?f 侓�)�ʐ>�W�>�>d�������p���b����?�F�?�>���>b=?��?�!:�蒰��P�-d����.G���Bt���k��N��&�������|?�t�?��#?��>�X6>�k�?����ʾ�?�>��Ǿ��{�g'���?c+Ծ�������$��p[q���:.u?�a�?J�?DC.��g(=���>`!?tyG?Dtg?9�?V#?�����?���>Tq>?�_M?�u_?��?P?+$|��~�_n�>���p���L���f��Q�彼v��Ӽ=N���v��;6�8�=����?��=�eL=�ܽ�=��<�U�= m,>襴>5�d?��>�8�<��0?T�=Ba�c��C2?i���_���H�u��	�׾�1��V�?��?�'W?e�~>e`u�����0>]oN>�ȓ>iK=�Ǎ>��<�l���,>Ǒ�>�Zi>f�M>]�I��������*��9>�e�B�?�K>A&��["�<��P����B�>���<����xT��'�|�����U	�/�>�vc?�aL?f��=�����>��v�vW?CZ?��?ݳw?Ҽ%>˪���@���	���������=�]D�G�Y�������?�s�">��b������=�=��T�D�����k�Wui�����H���U�0��d.>������w��).�lN���ܾ]�*��e�������<?$�~=���r�1�)YѾ�\�=L.�>D:�>��=T_���/�.����P=��j>�Z>a.�<O��wE�DLӾփ�>O9O?A�Q?;�z?ἄ���d���F��ľ56�GVA���	?�a�>��>:��=�����۾��A�'<l�&8��p?���>��,��!I�(��ٔ����(����>�V	?;e�><N)?F�?Kd6?$t?�?Z� ?��>)���0�*?�b�?s��^�`������O��eV���
?6�H?OZN�L�>��/?�� ?�,?C�?,�?��t=l�.��r#���>@�>Z�\�X����,;>�QH?E�>G�Q?�%�?��>�*�u�����[�>-�h>�*?thW?��=?���>lx�>Υ��="��>��c?oͅ?��k?���=Na?m7>�N�>���=Cפ>��>�?q�K?C<q?�5J?1��>/�v<�����[����K������<�H<��|=d�	�9~��YB�����<�kp�����ܻ
�ļ44�������<���>77n>�/��e->�ȿ����PJ>����G�����5|H�"ƽ=�z>�?[��>!5��6�=���>>��>9�?t(?A��>Q?�#�;�`��s�tf��>��=?Fc�=i�����s�M-a=ޱl?�^?^+M�+[���b?�^?�B���<�҅ľ#�a�+4�k�O?��
?N�H�Oe�>�?�q?���>��f��m�=	����b��]k�c�=�Ü>����\e�Ƥ�>��7?h��>Td>2��=�ھ>Dw�躟��D?b%�?!�?= �?P->�rn�%�߿��������]?b��>�&���n"?֥�޻Ͼ�������}��k*����������P�#�7�����׽(�=��?w6s?#�p?�`?� �R�c�t�]����V�`�������E�E�D�@C��}n��!��c��(똾Z�D=�
����=���?�$?M�E�f��>���L��>�ܾ�\N>`����1�b��=����i�"=��=��o�� K��ɾ,�?4�>|��>�B?UXY�g�:�k '���4��/��!�4>�\�>!L�>�B�>��U;>SA�����¾����x!��u>�c?b�K?��n?'����0��n���t!�7�*�vn����B>2�>垉>_�X�˷�T&�2L>��r���҉��6�	�-��=�2?9�>��>E=�?v�?�q	�]B��(�x�>h1����<
X�>g i?��>��>�Oнf� ����>�k?���>���>�_x�Dv�\���m�����>�_>5��>h�>�R�U%c�"0��/��g��L�+>�2\?<��ir�!ŕ>�&V?<I);��:�f�>�����u�۾J\]�ю�=�?�뷺��c>k����$�{�N���+?�f�>)���Z<-���>"?A�>`�>d��?��>s�Ͼ��<R"#?w�W???'g3?N��>��x=�6��@ʣ���I�%�=�rf>��T>��!>e&�=�b-��u��pڽ�ם=`u�=�a��ac��� <;)���]C<(�<��B>׼ݿm�A�Aܙ�=���Hؾ*A�����'�4�����?�I?�����';�X1��I,���*�nrH�����B���R�?Y��?�C;��-*�xK��wD�Zо֍�>~`��p�=�Z��IAL�T;�Cؾ��۾(��{J�}c����Ȕ'?����a�ǿ�����;ܾ�  ?�A ?�y?Y�&�"�[�8�� ><F�<�;�����Ț���οR���t�^?���>���/��2��>���>��X>wHq>��S鞾G(�<��?C�-?d��>N�r���ɿ����Ӥ<���?�@MC?x�*�:��:^�^�?1?m�*>$�r��v��䉾QS�>t`�?b�?��=�J���u�V?%,=ɉ4��;�:�=F=n>�~=��C�D��>Us>6���g|��ܪ�6��>Js>n���!��5�7�
ڱ<��S>��ɽ�L-���?>P��Bn��ܙ.�B`�Wd�>��?>�U?z{=S8g?�l����տ��M����?ъ�?ʹ?��?���)+>���.�f?~�*?�Nl>�c��g����]�Z�=����?�1&����>N`?���=�	��(Ⱦڽ�ϼ_�>n_��h�����`:���=Lw{��-'��Q���(�2���k����o�oM׽uա<�>�b>�܈>�{>�+Z>��X?Ji?�*�>�f>>Y���
����ھ'Ȍ�UЫ��D��0<�X�����ܾ
rξ)����� 9���Ӿ�=�?�=6R������ � �b���F��.?t$>�ʾ�M���,<xzʾV��� q���¥��/̾�1�tn�ȟ?:�A?f���}�V�d���Q����ұW?hC�ĸ�謾�r�=������=��>j�=���+ 3���S�.�(?KC? �ؾ㾀0�=O�ȼD+/�L->?�D?�m� ��>-�>?{���|���>���=Fv�>Jn�>���>\���అ�?�a]?�&>�z���!�>V���f<��G�>�\S<~�<s/�r!#>ɟ�i����V<7�H=&W?L��>4�)�K"�ٻ������<=kx?��?�>�k?�B?Tb�<������S�s�w�y=��W?�i? T>pт��Ͼ_c�� �5?i~e?��N>��h��龇u.�_V��?F�n?��?����KU}��꒿U��0/6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?t�;<��U��=�;?l\�> �O��>ƾ�z������1�q=�"�>���ev����R,�f�8?ݠ�?���>���������=_ٕ�%Z�?��?�����6g<��l�n��Xm�<���=h�T"�����7�
�ƾ��
������Ϳ����>=Z@tb�R-�>�C8��5�TϿ���}[оIVq���?��>ѤȽꛣ�a�j��Nu���G� �H�X���3��>^G�<��a�֋۾�a���)6��>]�?3��a@�>�����þ$�¾�>���r> ��>A��>|=���t�?����������!���n?᲻?��T?�.<?�x�>��l������Y6�}�L?Ѫ�?2�?��½g����>�j?}_��sU`�ߎ4�mHE��U>�"3?�B�>L�-���|=�>���>�f>�#/�y�Ŀ�ٶ����W��?���?�o�"��>n��?{s+?�i�8���[����*��+��<A?�2>
���@�!�H0=�AҒ���
??~0?8{�e.��^a?��d��eu��-�|fν5�>�j�*�L���ݼ��0�^�����V6���?J�?���?{	��y$�V=!?Ϋ�>\h��FȾ�/=��>n9�>C�I>- �їw>K�E�;��8�=E��?.��? �?>8���+��{q�=�y?��>H�?Y��=U�>&i�>#�{������uI>�G�>���;H<?�i?TQ�>�=�ڙ�9�#��+�i:-���̾?�L��l>}3�?%�d?l��>�l����ν�18����Q`�<T�=.[!���/=�ɽ+}[>^u�=�Op���'������?Np�4�ؿ�i��p'��54?,��>�?��{�t�[���;_?\z�>�6��+���%���B�_��?�G�?=�?��׾>R̼�>-�>�I�>F�Խ����[�����7>6�B?O��D��r�o��>���?	�@�ծ?ci���>ü
��Ig�}�y�������C>��G?�=�/R>�	?��7=��h�ڭ��Gu����>%t�??�?��>_|?Cg\�	HL����R��>)_?��$?�"<�����fU�>�?.�������ҾY�y? Q@�@<dN?�~��+�߿9&������߰��#��=aB�<�]>%Q@��<6c�<�A��R�]<��>��>��F>�^O>��:>V�z>�UJ>���	��9��������F����e�ya����cc�������B�����ڽ��ｃY����;�ӊ*���m����=K�U?*'R?0*p?�� ?�v�&X>.c��O�=��!���=G�>�}2?(HL?۝*?��=
����Xd��[��z������0�>KJ>���>���>۽�>�A���F>�=?>졀>- >�B(=T�=)�N>T�>ɸ�>3	�>�C<>d�>.ϴ��1��2�h��
w�+̽3�?q���D�J��1���9��.���Ui�=Hb.?^|>���?п@���t2H?&���<)�Ź+�/�>Y�0?�cW?Ӝ>���T�:>���j��`>�+ ��l���)��%Q>Kl?b�f>�>�=-����S��k������y�>C�b?�,��L^��D���F�X&���>H�>��=eQ�q֒�H/�p���w��,H?�;�>.�X�P���z?��ξƠ=��=�U�<}H%>���>���=He-���~�g�=�J>���=]J?b�+>%��=��>�Ϙ��N�=�>A>^�->�i??ı$?׻����������[-�
Xu>���>B��>�u>QoI�խ=A��>�%a>ȹ���肽!� �@���W>:y��1`��|w��{=x��ǥ�=@g�=����s1<� �!=�~?���%䈿�뾞d���lD?O+?) �=ܟF<��"�D ���H��H�?o�@m�?��	�ڢV�?�?�@�?����=}�>�֫>�ξޔL�۱?�Ž9Ǣ���	� )#�fS�?��?��/�Wʋ�9l�6>�^%?��Ӿ�a�>)���V�������u�E�#=%��>K8H?a����O�O>��o
?s?d����.�ȿ&~v���>=�?!��?��m��?���@�@�>���?�dY?��i>sk۾�eZ�폌>��@?�R?��>�9�g�'�s�?��?��?��4>jԐ?��n?5C�>���<��+��V�������w�=�����m>/r�=��ȾmJ��e���a����x����:>��l=�x�>/���o���{�;���_�����9;���>
ed>��G>kУ>�� ?�5�>�H�>�Q=�-�eԟ�]i��pK?w�?���{�s��p��M,�=��m���?��=?�����nƾ�>�6W?��?~^R?�-�>b"��ḿ�:��%��<;Y@>#��>Oy�>���{�r>�ʾm/����>C�>H��<0�+r���[v��Ӓ>�O%?vi�>��=5?�%?��o>+��>xC�PD���9F�X��>���>R�?��{?CB?�����;3�sՒ��E��}�_��;>�s?O!?�ɓ>1���Q���i�C�ix#�1��/G�?�f?%{Ľ�|?j�?�zC?
�C?EUf>����WϾm��>�|>+�?����e:���)����$�?��?���>Ǆ��� �g荽8���N�� ??��Y?;$?_.�Ƽ_����V	=B۶8���07�<����>y>*L��h�=F>�D�=BW�ZA(��`=<�=��>F��=�(��ソY5,?nD��ჾUx�=��r��gD��S>�L>s����^?)=��{�(
��w��ztU���?��?�h�?����$�h�<&=?�?i?��>�@���Y޾���u^w�#bx��w��>��>3gr���������F��<ƽZ�\8?	��>6�?X)?U@>d�z>�B������m�Q����TF����1J�\�3��-����������S�Ҿvgh�`˰>[@ݽ�D�>�'�>�C{>�8�>_��>H{O���4>���=��^>m�>a^�>wG>��ý��3�^P��;�Q?����&���MD���B?5hb?.	�>�HG�Kك���2 ?�6�?��?��s>R�f���)�]�?�G�>�[x��_?ĳC=Ѣ0�q�G<�ί�N�s����
��)�>��ǽ}�9��8M� �f���	?8f?�d`��rʾ� ѽ�f� �}�r�?
�A?��I���p�oJ��O=�f�d�f=����Sf��q#���y����s5{�{%��xZ�� `��g?�]?�Ծj�	������T:�����ן>e��>���=�>1>]7꾂��_mA�2! �Nˎ����>^�p?�X�>?sU?O�6?�ya?��S?�σ>�6�>�%���e?��	>iH�>Y�?�l7?��?�/?�.�>Pd�>zZ�>��ʽ=s����)��>И?��>/z�>�?���q|ɾ��v�-|*�%yQ�cٽ�1�=��+=���-��ٙ>$��>?���P@6�d��6_s>�i9?���>���>����Ɂ}��=h)�>��?%��>���I�q���!�>w%�?���a�<У*>F��=������;�r�=T¼H��=�>����"��%<m�=�i�=ӄ4�+�;�z:!�N;�<ۓ�>O�"?FgA>gN>]T�T/¾�{*�֯��1S>u��l@>�Ɛ�� ��W���Ɇ�nq�>��?��?&V=!@;;��*=����2x��o��8���>%=�Q?�n�>A�,?��?��A?�?'�<<zc��Z��:o��Aˣ���?�,?^��>���ɸʾ憎��3���?�^?�:a�f��m?)���¾�սq�>�W/��*~�����D�R�����"������?8��?>A���6�v�k���]��K�C?�>{\�>_�>h�)��g��$�q2;>֌�>�	R?��>��O?:{?��[?��T>��8���ƙ�� ,��">�@?c��?.�?��x?�{�>�{>�)���߾M`�� ��~�dЂ���W=e�Y>�k�>m:�>�ĩ>��=_�ǽ���8?�w��=�b>��>���>n��>kyw>qx�<�DG?���>k�����>��HBu��Nx�n=r?�?��&?f8�<���,�D�R��Gܼ>�T�?���?о'?d�C�(�=^���/�����v����>���>-r�>��=M؄=7->0��>:��>_Q�Pf�)�6��Y���?[sJ?h��=eY˿��Y���>֮ɼe"�D���P��A��^���!>�X��`#���0��5����է�V���2K��~�r?�W-=��+>��>�X4�ԍŽ�T!=��4=�⼽r��=es=���޽ȈU�~�����A��ȶ��j���c1�i��,���x�?�9M? 40?a�J?��>��>�B�8�>mռ؀?/�>�\�������	�ƍ������p¾�>���Z��ܬ�}t)>�u��N&�=W>��%>ᄼ"?<�׍=>>�=Il�;{|=k��=�8�=���=h��=�3>e1�=�͂?+9���:��>|v��ᾧ�^?z%+?�|>�����:�?_��>:������hE�BZ�?�~�?扱?9
�>K����?p	���u�r>�fY>Z�?�?B��	�#� ?0ܞ>�ߺ�{h����l����?y��?/�?��W�ͿCc��U�7>˿>��R�v�1�eS\�O�b�%�Y�
�!?�2;��`̾���>�W�=�P߾�Bƾ؝/=��6>��`=���`"\�X�=�\{���==��l=?w�>��C>�u�=����r�=��I=��=%P>I���5��,���2=e�=}c>�
&>D��>%�	?7�$?�\\?%�>"Jd��a��3¾�~�>PUK=m{�>R��=[�~>���>�/?�&:?��;?�B�>�	�=}�>�n>=.�ɳq�c|�����O��I+{?�1�?�>�ר��m�����b�8��ﱽrY?�1?���>�c>9���JϿ����f�/�I�|��c7���b����:��i�u4e�iq�����=�zY>�C�>�K�>�~k>�Й>'�d>+��>��0>��=�iQ=�<����W*u��/c=+�~���ݻ�tƽM�G�ɽ6A���թ=�_�=,b=����9�4B�=�#?pj>l�>rp�=Kݐ�k/h=�B���8�?������ ��jZ�j�����@�x[��ɈH>%�j>f��瞒�59?�C�>�>=>[��?��V?lb>�A���6��/F��F롾9~�����=�ݗ=�S��V
6�'�~�7sI������>6�>�>��m>g�+�9�>��ct=���>5��g�>�K��(��
z��[q��B��5���o�h��ݤ��[D?�H�����=�*~?7�I?0�?�N�>?���0^ؾ�K0>gE����
=<"�'�p��"���?�&?a��>�.�>�D��pξ6kW��1�>��"�ff�$e��/a��nI>����L>�V�������W��F/���M^������>{�8?1ץ?]�t��1_�:BI�@&꾄�/f�><+x?��>)��>�*?��V>��(���}->[w?�J�?-9�?�?�=��>��!-�>Tj�>���?�j�?�]?q��V�>�#��&V>��=I��>!Y>[�=�==�>�z?i?p�'�$�&Mо�z׾��p�<C�=֯=�z>��>Ja4>�� >�����k/�g>$��>�4�>��Z>k�>��>��;��	�5�?H�=��>,?肀>FX�|�=`�=N�Ž����|��=hZ��N���J����ջ���=^<x��>:������?2p=�ͪ�?�?}|��-�<�>��>��E�iH�>B$�>�e>�Í>�>�@>�V>3�.=��,�=��Hq�y�U�5Y�ِ��0v>J���*�� �o�����@�����|y�����+C��Vu�牉?q�%���W�j0*���˽�"?^�>z:J?f 侓�)�ʐ>�W�>�>d�������p���b����?�F�?�>���>b=?��?�!:�蒰��P�-d����.G���Bt���k��N��&�������|?�t�?��#?��>�X6>�k�?����ʾ�?�>��Ǿ��{�g'���?c+Ծ�������$��p[q���:.u?�a�?J�?DC.��g(=���>`!?tyG?Dtg?9�?V#?�����?���>Tq>?�_M?�u_?��?P?+$|��~�_n�>���p���L���f��Q�彼v��Ӽ=N���v��;6�8�=����?��=�eL=�ܽ�=��<�U�= m,>襴>5�d?��>�8�<��0?T�=Ba�c��C2?i���_���H�u��	�׾�1��V�?��?�'W?e�~>e`u�����0>]oN>�ȓ>iK=�Ǎ>��<�l���,>Ǒ�>�Zi>f�M>]�I��������*��9>�e�B�?�K>A&��["�<��P����B�>���<����xT��'�|�����U	�/�>�vc?�aL?f��=�����>��v�vW?CZ?��?ݳw?Ҽ%>˪���@���	���������=�]D�G�Y�������?�s�">��b�
`  �   *�>[���fM�"BG����Y� �ו�<D�?-����g>��d>�
>�'��
������_	��<J?��?��T?�{5?W���羋����=X>�>r�>�¶=p[�XI�>[��>^뾝�n�MX���?[*�?���? W?��m�௺�8�u��U��$���p�\=zW%�L^>X����^o=i�>���=�|��K��=�~�=�ʐ>!ٯ>Y�+>�3y>�c">����9�?,ɿ\$���)y�b3>���7f�<u�3�/_ȼ}���1��P �	y �{���ǋ�C�ž�|�/�<Pھn��>�??��>�<�>��>�+>�E�¦�`
�֌p�ᾥ-���(�mj`�@2̾�vվ��?�
)���mR������>5l��0�m>4�3?����#u>dJ>�0g��:�=/l>�P�>]�>��>̘>���=�xw>������4���鍿�u��K���A�]�E=�~A?*�<3�ƾ�_��4	�`�>YpY>y��>�->���;�u�N�>8'=C���۽;������u�=1��>-#�<s>��e<���:�=1݀����>���>�U��_������<�2>��>&�þ�>Al>=��?Q�F?,��>���=<k�>�ua>hb�>�Q���@�<�1�>8�H=�o�>5 ?�g?|��>�#>w���;��5�B�"�r*���=�B�=i�z��l$>3s7�B-���<���TL�����|=*�>N�z=�s8>�:	?A>5?�A?�o?�$:�2=�06��A��=�N�=F�>
�>�q?,~�>+J?�U>�|"��E̾y�Ǿ9u�>�=(pH��=U�{ی���>��>�SM?�<3?4#�������ڊ=w�=z]�>��>_	?`'�>��=��=�y�^�ѿk�&��3#���h�W��8;0(�\��lQ�<.�(��w"�!{�:1U>#�>��q>�1>�t5>68>�{�>i=>��Q=��=�D�<�n{<y^��$=H⼉S+<�en�p"M��X��1��"���TՈ�YJ����R�n�?<�$?���=N:�=Ȱ�ՙվ�{���*t>�T?d8?�=?�o�>Aܦ��N�h�[�]L���?�tR?�l�>.�����=��%�ϼ�t|�>���>���=%��'��d��Π�My�>��>Q�O>�	�r	6���e�����>pJ�=�_I����?��L?5�Ǿs�����A*M����#�ҫY��O�<����~&5�l��d��K^T��1>�`�>�ͬ?�E�<�P�>S	<��b���T��%g�7�=��=��>�5>�,��Ů�V!���a�JGm���1�u�=��,>=�>�;?gbM?���?�X$?�)�>�묾%�?�
>uY?�}P>�0?��3?��3>^A�>~�>6*>=���R�M�������<7�C=P�X=��>q�N>��e�f>UF>2����̸�����c=����\;>���>�+Z>U�>�?i�,���9��᰾}��=�R>duO>f����톾��N�Zb=i�?�7?�>��0>�z����������3C�>�A?e]?��>ql�x:a=Y��_���x�=�I�>n��˽�����4о����"�e��>�Q�=�]a>��w?�_?��:?�*�=��dڌ�q d��8�mo/�{�>_q�>U|Y>}z��� �X�7��rb��d�����K�K�c�=v��>�p>l��>��6>m#��j�ʽ�v�=��^=U�">�"�=���>,C>�a?��>�>u����;���A?����P
���Ծ:����*��JHb> �>~4��?�Ou�;Ԁ��頿-y8�dD�>���?'ֿ?��P?O�ý/��k �>
 P>�~>�I�5����	��l7�}J>��^�).U�ŐF�b�l>M۞>���>/-��6������"�n��a˿�U�vs�@��Yؾ��)�g'�K�>����L>�ɾ�x�n޷�3���L4 >�$2��L��C\��疾QRl?�?�aؼ��3�ϗξ�����(྄@)�Q�1�Gê���̾���<�u��I����Ծ����왾}�,�#d,�%�?���偿=K�	�)�۵=KM�>1�>c���������ͦ>�Ӫ=~T�=�������Z����v�V�x?G*?����42���P�=s�?:>��>1=�.8Y�N�>��?.m�>��=�Y��aᓿN�;}�?���?ԕc?�ɷ�,���ھiD��3(�>��?<Q>L_��Km��*r ;�(?Ƒ?.��>�Ѿ�A����G����>�4�?������>�$?1�>�뽿�䚗��r��4�Y�23�>.� �ɯ��o=q����'����>�%�=z��;?����>���f�K��cE��_���$�
9�<��>"����>@�r> �>�"%�l�\㊿y6��(I?��?�6W?�w3?4F�Q���(��[�=��>�o�>	g�=#\��D�>�>����(l�f��b?3:�?��?ҜU?�mo�xWпK���䫾X宾�;)>�, >E@>�3���ػ=&��=+�*��I�;}>½>��y>�$�>�&g>@V>�G>͉���(�Mz��MI���6��߭�-MN��?�tc��^��ƾ�۾�� ����)1Y�_81�C
��n�ģa�ai>zj?a��>1��>x�L> �=NV���	Ծ\���=���_k�筬��A�ÓǾ��z��5���Q�R�l��w���/��>�%��ā->vv�>�:���"�=���>��=���=l��>H>�kC>��>/�b>ᴽ=���>�>i=57�>��ؽ6䐿��j��{־D6�i]v>��1?�e���ɾ��ِ �0�R��� ?�}�>��&>��0�L.����X����>�8ֽδ}��b���,>|��>�G>����W �n����2ݽ��.�`�j�N�>�J>O����h���������=c�>����P��>X��>�L(?ꇄ?5�?O=e��>���.�>���>9��>u��=� �>��?�%?n�-?�ڻ>�K�=� ���0j��A��.�罿�I�ޘ�Hw��Q�=ێ���M���=�m>��~>]�F>B>b>�4�W���~?3M,?�c�>ێ?6m���x!���7/��Wcs>G�>�q?)�>��?h2�>/?���>�F�>��=�{��L�>���<G_Y�X�v�� ��D�>=В>�!?���>�(��FӾR�x�V�;,f?˅ ?�`?���>F��>/�ؽ��0����i�\����	�	�>.�s�(��<J �>�O�;=����;�t�;˖L�7�e=-��>ſ�>׏�>hq>��>$'>�86=턢=�ю�뎼��=�QE>B�=[���Ҽ���5����ELc��p�<|�b�vY@���;�� ?�?ܭ>�I�=a����	��;ξ��>�>�."??�9>>�}��
M�a�?�0�����>�
d?Yd?|�o�^�>�5�=MQ��/ƫ>xH�>�;�=ȫ�=Yǔ=N���)��P�>�X�>vh2>�	�V	7���I�H�Q(1>i�8=�����.�?�[?r��kwн�f�H�_��g���x=��At� ��j�&<����L�վ*�D��a>�{�>g�?bS�=i>9��<K����r���|/�=:�=�Ģ=��%�yU{�%�z7�H��q��l�D�*�="��=��>�Z8?�kQ?~�m?��?^H�>/���	��>>
.?M2�>�0 ?�{?h_?���>K�>wjS>�&�l��e������I����==+��=r��>&>�=6[A��l�=�>a�=hN�@��;*�o=:Q>IZ>�X�="��=.1?O�?�i�������>��`��QP�J>!b�=%ﶽȜо^PB�1^����>.�?��>&�>o�7�"�H�LD�=
E?9�5?Fc�>�1A���,=&"�������=�*�>��"�u���Z������:��>�)x>.E�>���=�sv?J�Y?��6?��=�|־κ~���E��6�=?�Խ��m>�>�>��>7�+���H��FV�%5��k��ͯ$=��8����CD�=z>I><�Y>ֹ�>D)=8����s=o� �� ;>E�>ؓ[>���>���>��>3-�=T��O��y�I?�������<��y_˾#�S�>y";>#X�l?�E�2�z�{��-�<��;�> ��?�U�?C�b?��F�8���\> �W>�S>#�;gA�,K��Ll��1>���=#�x�1���7�;sVd>�,{>Nս�Ǿ���~�Q�k��� U�Ҍ��[����@��;�L0>���5(��&���9��j���x۽0QK��^+='g���g�!tf�L��?^x�?�^��k����E��Q:�U]b�Rp�>p)��@"|;Dg�p��Ĉʾ��b�t���V�	���/��d�\���"�>F>=ׅ���!U�f�U��ڽ^#?e?���󱃾5���銽��=#���E��g_��H�����S?�[�>�`�X[���>S%�q��=V�>>K�>�vf��˸��޶>h�?y�0?�oN���Q���LF��� �?酢?�9?鎽��%�@����_��>��!?DU>$�ݾ�F�I�>��>��>[>�>���,M��:�J��	�>_�?�����M>P�*? ��>����־=1P��m�WyK��Z�>��<��x�!��=M��*�n��K>���>�"��� ��4�>���]�Q�'eF�e���,���=�y ?�ﾀ��=�]>>��-��5���9��>���VL?��?�S?c7?c���^��਽��=*5�>���>r�=�&�R7�>�?�>�&��r�J��\?>�?���?S�U?@$l���ֿ����&��oh۾2=�=�?�=w\�=�;�3�=��~�(\�!b�<��>�{g>�\�>��y>W~.>a�>�y>)���t)�K�$��G�)�lE����I%�����]�������þ�a��ƽ��k�#���%��3H���_ 2��=k,����>R�{>t��=w��>�Q�����;�����2�Cg*�i�?����C�
��i���P�����F����C?O!�d+�>�? Hi��/�>i�?Ύ_=�3�;�"��?�=j,�=��>�
�>}8����?�>�|�=��">~t�e�Z���]��%����>zuO?�Oᾰi��N��c����E��>`ފ=S I=��H�G+}�|Ʉ�<��>Ovn<ə��f���%$��=.��=��=Ɔ�=I�Y<	_�]��=�,�<���>�<x�=í.�clؽ��>��>q̾ؤ>?Ʀ=�1*?���?��k>�z�?�O�J>9�>\ �>����+	?�WN?eR3?�c?��,?�p�=�o������Ȍ��%��2D����6� >	G*�H���E���ܗ=:�=٫I���=w�=�W>�Bg<(01���>~1N??�%U?�J�<(!�����v�A;R>�)>��?��>��C?�/�>iQ ?�^�>n1׽���5�ݾ�p�>��l>�}>�Y�y�؈߾�_�>]M>��>�~?�9>�7���2�>ٛݽ)��=.=�>��?�W?@*>�e����7���*>"��RZ�*1)�^��<;f�;P@DK�f�ɼ�2޽`����/B=�kh>Ě
>�~�>��5><�x>���>��C>u��W2�=���s����U=�U=�r����i>#�=�	����[���ܼ����d���'�ƽ����<�&?��F?�r>|�B<P��M�����4�=Z]d?�{?]3s?ȑ�>x������@�M���w=�?�(]?Wy.?�go�9�Y�`?�=���=��?��>�<O=����Տ�":���>Eɂ>��?S}8>�"�a"�&u���ھ< �>Nq>!f��W�?��l?�3�:j����?���-�D?�n󼜶[�7�\$/�so���$�أ"��7B��J,�u`=桵>aw�?��;��=l�a��.��u���&J��ʉ�[R޽Zl�>1�?Н�Q��
M�NŠ��:B�����>�>h!%>k�y=�n?K��>��Z?C�%?,6�>�9̽�A�>�A��]��>,G?|@?	�7>/W	?.�?�R�> n>v;>>�ؽYً�� ����U��J�=@�=�y>��}=qYS�NA�+��O�V��$�'��!��<�@9��e:=d4�<3 �=�u�>3��>Mf>�βJ��W4��۾����!��>f���.'�<���?��=C�;N�>P?��>S�R<<��z�����̾2y�=��?�1W?���>s�b������p��F+*��̧<1�>����(C̼�L��'g�UҖ�������>�m�>��>���?a�f?�ij?ݑ@>
h�팔��	��%&��_���5?� �>���>gs��Ou!��Wb���m�{�����<�>-��dĽ��z���>d��>2��=L�>�|�=��ּݤ$<"�!>$c��A?�?�?�o>%->����h,�m�I?�'��J�����ݿϾ�+���>��?>�1��|?Y�
�d�|�x����W=����>��?�r�?Ҋc?s�C����{k]>�GV>�m>�<&�@����y!���M5>��=�9u�*���Ҋ�;�[>rQw>��ý�sʾ�`�qF��@ƿ�t�!��岰�9���⹾'��l6��ɘ����X��I.����x���赾G���O��Ź���
��m�?�ً?:�;>�ӿ=��%�\�0�������>�Ѿ�ae��ھ��ϾuԾ�����J����
�ƻ �qB�R1H��n|>, .������`�{)�ц���{>;m?oؽ�����e���dwx=���=+Lɾ%O��b���aR���C?vW-?z���7�ľ�LҼ�UK>U�%?��>z3�=P�`��Խ�l�>J�'?���> ����|�@ь��4[<�0�?��?V8?5k�����T��};�����>�n?w͠>�h��A��Ƙݽ@�5>k��>C+? q�k���=3�L�#>BL?��D�%(�=�� ?���>�#Y��逾gG�<\W��S��4�>@�=�\��y=l�+�l�,,~=t��>���/?�����> B꾝�N���H�~��F���e�<�?��k2>6i>0A>)�(�����͉�\���L?���?b�S?&j8?�^����P������=T��>9ά>���=��I��>���>�b込vr�v�)�?�J�?	��?i\Z?��m��a�����#��8�ܾ��=$ʤ=�N>=�$���=!�!=m�<��０n�=��>
t�>�T�>e��>�� >��>e@��.�%��=���
����^� �"����Y�M����鑾(��{z�����������I���Q��rŽQ+��)fO=�c�+�>�Ǭ>��>&=>sڡ��>ݯ��n�<�xQ��o}��`%E��4�(���'�a%̽a��W߾����jk����h�U?������>�i<?!�I/�=�
?����\?�ƛ>�n�>C�>�i�>��>�>L��>��>u��>֋=>��늿f���g�ֽ�+r�{�??���H��$y���!���2g��2>7d=Cd���>���dx���T�>�5�<+G,�jZڽ07�� �8=��5>8�K=��ļ/�L>��6
=9�;��L>��S>_�;��UV#�\]S��ً>�z����>���>m'E?��f?�g?�#�޽"?ֶм���>!T>�>��=C��>+Q<?I�#?�Lf?sI?���=���q��)T=	��@�Ž���ޔ�=,)��eF��l�B�,R��>1=-�=5�&<�{;=���=���=�o=K�>�'Q?},?��>��:<�׾��r������>:8n=��>�N?Z�=?�aA?n!?��<��4�Cߜ�~��.��>`I>�9��8�L�q��g>�k>J�2?�;$?��!>�T��F7<�w�< i >)�>MzA?�'�>	��>�.*�j%�G������5�2�_d>��8�ı���^���I�w �=vA��_�]�5�;T�[=��>�A�>��=��6>�TW>�=�>t��=#>m=��X>�-�>���=m����`�=��= �`����� is��<ʼ]+/<ޡ�xj,=&	�=R�_<����8?u�"?�o>��=|=ozؾ�O��ms> 
?�0?��'?��>��|�w�L���\�$�4�N �>N"t?�7+?�*ǽo�><����J��\>�I>�������ֲU<�_U�ۿ�=E 
?�v	?#��=.�]�w�V���m�_��tݸ>���=?n��^�?tfj?_Tؾ�G$�~��� <9����v���.���:�R�3��ں�'������]�:;>�i�=_��>}�?a��Y�;��W�g���㙿o/*�p���`X2>�r�>�;�>���6@���j��8���Ӿ�=@��L=���=���>YI?�b&?L��?�^0?���>V衾Ɩ;?V�>��<?2?oW?=�>:q�>d;�>0`�>�@�>�v>�G�fC�������=k2>�8$>���>5�=��n�z��<zX����S��C�-<�� ���OF[�gtZ>��|>���=�?��?���(E���xZ���z�����>�铼�ȁ>Qq��d���.>00?��%?2!B>�V��ͬ�v��O���Կ=V��>)�T?�N�>^[���%�Ry
��N��t�>~z�>�ڿ���<��ؾ�Z�|���<�Z>I�F>�W�>Fc?0_?��9?w<�=�@n���������>���>��>1�b>D�Ǿ��&��:��=t�Y�ϾG =(��^r=��(>`p+�'e=R�=�b�>������\��;Y=�[=���=���>?#6>��������.y��I?p����6����Ѿ�=u��">��[> ��(�?���^}��D���7�g��>���?�?F�`?'�A�s\	�x_>4�S>^%;>�N�;�zN�m4��݇��?>�ս=��l�6r��>��<��O>�Uj>�����Ӿ�&޾���s����SE�w��Ғ���qݾ��� �r�a��<s����=� ��A���]������!ƾ�3,�
l��⼙���}����?��?���$qj�*8�ͱ�3�'��B�>A꡾l����?��Ѿ23$�u���/��.=��C�e����C�t��>�mW�bD��3�{�(�(��ؼ^�A>/?LɾT��Ԑ���Q=�<">w:�<Ƕ�i���������U?��7?���g���ѽ�>�?���>�)>�B����轟��>ٺ2?Ӛ/?��� }���$�� .����?���?�w>?�B�7�B�����&�pV�>��?�	�>�g����Ⱦ����?�I-?B6�>��ۃ���w��>�TK?-cF��;]>ݣ�>K�>�����T���B�YВ�f4��2?>��溏��2�n���>���=ί�>�tn>
{R��v���4�>���]�Q�'eF�e���,���=�y ?�ﾀ��=�]>>��-��5���9��>���VL?��?�S?c7?c���^��਽��=*5�>���>r�=�&�R7�>�?�>�&��r�J��\?>�?���?S�U?@$l���ֿ����&��oh۾2=�=�?�=w\�=�;�3�=��~�(\�!b�<��>�{g>�\�>��y>W~.>a�>�y>)���t)�K�$��G�)�lE����I%�����]�������þ�a��ƽ��k�#���%��3H���_ 2��=k,����>R�{>t��=w��>�Q�����;�����2�Cg*�i�?����C�
��i���P�����F����C?O!�d+�>�? Hi��/�>i�?Ύ_=�3�;�"��?�=j,�=��>�
�>}8����?�>�|�=��">~t�e�Z���]��%����>zuO?�Oᾰi��N��c����E��>`ފ=S I=��H�G+}�|Ʉ�<��>Ovn<ə��f���%$��=.��=��=Ɔ�=I�Y<	_�]��=�,�<���>�<x�=í.�clؽ��>��>q̾ؤ>?Ʀ=�1*?���?��k>�z�?�O�J>9�>\ �>����+	?�WN?eR3?�c?��,?�p�=�o������Ȍ��%��2D����6� >	G*�H���E���ܗ=:�=٫I���=w�=�W>�Bg<(01���>~1N??�%U?�J�<(!�����v�A;R>�)>��?��>��C?�/�>iQ ?�^�>n1׽���5�ݾ�p�>��l>�}>�Y�y�؈߾�_�>]M>��>�~?�9>�7���2�>ٛݽ)��=.=�>��?�W?@*>�e����7���*>"��RZ�*1)�^��<;f�;P@DK�f�ɼ�2޽`����/B=�kh>Ě
>�~�>��5><�x>���>��C>u��W2�=���s����U=�U=�r����i>#�=�	����[���ܼ����d���'�ƽ����<�&?��F?�r>|�B<P��M�����4�=Z]d?�{?]3s?ȑ�>x������@�M���w=�?�(]?Wy.?�go�9�Y�`?�=���=��?��>�<O=����Տ�":���>Eɂ>��?S}8>�"�a"�&u���ھ< �>Nq>!f��W�?��l?�3�:j����?���-�D?�n󼜶[�7�\$/�so���$�أ"��7B��J,�u`=桵>aw�?��;��=l�a��.��u���&J��ʉ�[R޽Zl�>1�?Н�Q��
M�NŠ��:B�����>�>h!%>k�y=�n?K��>��Z?C�%?,6�>�9̽�A�>�A��]��>,G?|@?	�7>/W	?.�?�R�> n>v;>>�ؽYً�� ����U��J�=@�=�y>��}=qYS�NA�+��O�V��$�'��!��<�@9��e:=d4�<3 �=�u�>3��>Mf>�βJ��W4��۾����!��>f���.'�<���?��=C�;N�>P?��>S�R<<��z�����̾2y�=��?�1W?���>s�b������p��F+*��̧<1�>����(C̼�L��'g�UҖ�������>�m�>��>���?a�f?�ij?ݑ@>
h�팔��	��%&��_���5?� �>���>gs��Ou!��Wb���m�{�����<�>-��dĽ��z���>d��>2��=L�>�|�=��ּݤ$<"�!>$c��A?�?�?�o>%->����h,�m�I?�'��J�����ݿϾ�+���>��?>�1��|?Y�
�d�|�x����W=����>��?�r�?Ҋc?s�C����{k]>�GV>�m>�<&�@����y!���M5>��=�9u�*���Ҋ�;�[>rQw>��ý�sʾ�`�qF��@ƿ�t�!��岰�9���⹾'��l6��ɘ����X��I.����x���赾G���O��Ź���
��m�?�ً?:�;>�ӿ=��%�\�0�������>�Ѿ�ae��ھ��ϾuԾ�����J����
�ƻ �qB�R1H��n|>, .������`�{)�ц���{>;m?oؽ�����e���dwx=���=+Lɾ%O��b���aR���C?vW-?z���7�ľ�LҼ�UK>U�%?��>z3�=P�`��Խ�l�>J�'?���> ����|�@ь��4[<�0�?��?V8?5k�����T��};�����>�n?w͠>�h��A��Ƙݽ@�5>k��>C+? q�k���=3�L�#>BL?��D�%(�=�� ?���>�#Y��逾gG�<\W��S��4�>@�=�\��y=l�+�l�,,~=t��>���/?��_>�Y����]�ϾE�x=�ٟ���mb�\.?jf����>�8>�d4�\���	e� V��W1?�v�?��$?Q4?��"�۾_��<��<��U>yQi=<�=�[ ��^�>�4?���0��P"��a ?�?�?6��?Q<?��l���ҿm`���������~�;=�\�V�>��k>a��=�mҼ�>��3 >G�{>9�>a�_>hO>x�Y>qx�=�"��K�"�})���܇��L��3<��,"�>T��i�$6��J�	��G������凶�?�ْa�ѩ;��_���T��9�6=�T�>�@>�Ɔ>
`">*>�D��f�y�	������	������l�h��ԅ��u����{��L+�څ�2t?�B��q>R�>���=)	c=�w>�9$=���=�9>�S=���=M	k<�mn>��>��>�4:>QN=�+��u�|�ݱ?���Y�0ٔ��;=��Aj?��؝*��S���U��
�3]J���>�݁>=����W'� s��s�>V��o�@���>,^��%��=�Gz>�	)=�W�m>b���P���y>��>���<m��=A@~���ھ��E=�L
?sF߽&V�>�5^>�[?�n?�YD?�U��|�>�� ?U���`����>�A�>��=B��>�&1??Ul?F�>��5���K�c%K=�0(�i���b��2=�	>��m=�x�9�������<�<�l�=������6�=��漿n?��|?�"?$�?4�y=���&�wn��G�>w>>̅>?M?ԟ�>���>��?��>�ƾ�Gz��9!��v�>��=��C���V�*�c��%�>��>�QT?F� ?昕��롾�|9=I*�=>I>f��>;H�>���>~dU>��a�!�M��K�*�{g<�H�%��X<u\Y�`?4��D��ה�Hv+�(�������6߅>�Yq>��#=XH�=ͤL>,�k>
��>5`>��<>�gH=�j���%�=ݝ�D=x)=I��B�X����=��ʽ��/S >�%ս�!ٽu�e=kvg���?��?����������V��
�����.�>�h�>��>�P�>i)�=o���O�l7���Q� �> (i?�?�{+�ּ=9�L�촌���>C�>�=�8�~kֽ�^��}C"��7�>�[?�Ǭ>��'���S��.k�Z����>���=�g����?��u?��k�"񛽥�*��h��r��m>��E�����򇭾פ��7[��mپ;�"�~������=���>�7�?/Y�=�U~>����+����$���о
@=���<3�>v0	?��
>������.辠Z�=|8���>�a>kl�>��?�?�_m?�@*??-?�$	����>���=���>��>��"?�
?��>�	J>�xm>=(�=B�"=x�3�����<��2=�� >��>$U%>/`;% �<��=��)=2aý>������=����Լ���=���=�T0>�\?�?�z>��>�����5����׽Ƽ="��>��h���>��h>){?��?VH0�a�F�� �N�"�X�N=.)?c��>=�b?�K�>;��>�]�K�`�ߠ>�e7>|�!�Л���5�t ��\F���>P�>���>�H�>�ӆ?�R?��/?c���?%�=���4A����z��:� �>d��>��3> !�����Y�H����=��[,�j�#�+��=�ř=Є�=�d�==P��=B�=��0I��*d=}> ��>���>�?�[�>1&=����Ћ�4�5?-�d�Z?	�I����_̾k)A�E�=�> �8=Ji?�)��[��5����C����>�x�?:��?.nJ?�k��\h��%��>�	�>Z�)>&\���6Q��X�3�)�?�>��>z
V�tb���摽�m�=���>���Z������	5��tʿ5�h��l�l\�[���#J�������=�.�\圾U�ͽ����þ��F�`�}�� ������M3%�\���gz?�l;?�SþցW�`���~�X�����J>�A�䱸�T�<v�=�1��-8���Խ�kھ ��K4�R6���h�> oq�������w�t�(����=�3>�h/?ɳ��S�þ�O��oc=U�>��	=Mݾ����㕿��꽌�R?' 3?*9ܾ����}.�=�?~��>��>�|��*<۽�ƈ>2I/?�-?<y"<iㇿ���~���?��??7�Ľ�:	������n�?�??*
�>��⻎ƾ�6þW�?��9?_p?Ou��G���,U��?�t_?E�V���='��>��>������ؾ�՝��޾�)�=�s>�%��
�=�"3���R��Ab�0ښ>/^�>��e�\�[�G d>	��|p5��'V�T�����v.��?�H:�{�t�k�V>�m\>m'�&o��%���
�F�h?�
�?�P?�u9?�ô��,Ӿ��I�?i�=�Z�>��N>��>Ԅ��8n>�[�>�W�!Rf�`T�Y/�>��?��?��-?x��tb��r�m�s1˾�ھŉ�=3�=��%>W�'�b��xG=obx=g�����%> �><�>��e>��i>��=�����5�<߹��G��B$]�<!�Zz �c#@=�/ ��H�y�оG�����v�XI���$���b���H�o���R�޾�
=�ɵ>�>�S>]kz=J��=�i1�%��D&�����{������;�ھ�~��\޽�Pu��^����-��V�	`?R=I�>���>����Ⱥ�Z��>�U�=^��=XC�>'>�>():>�^�>[Y,>�'>!��>�:>1`�=���,p���a���U�K��^�A���b?����������۾�3���>S#>g���$�$V�� �}�w��>�<�B=M�>n��<T�<�� ?�{/�P�=�0Y>o'������>>Z?��c>��S��߾= ��A|>1�?o���a>`��>�I?ڕ�?ف`?�`��� �>�\?�.��"����>��8>��=���>�?��,?)�)?�o3>XO���GO��\<|0[�6�=��;�R-�<�Z�=ӻb<�� �7�5>9Y��s�t���H��^=�� ��=�J�=�Ӿ>�c�?��C?��>O�c=��;��Ŏ�Qw�'�>q?�<&{?�>?�w)?y?�>��;?��>��v�Q��X��M;�>z	
>��<��sR�ś�����>���>ol=?�[?���&&��.��=߽��`>~��>9�?��?��>�([>�;�������8���"����{>�|M��;wp<��ɽ�o�M��<�yS����=l�U>��>%�!�.��=R�!>>��>�k>>�K= �O>sq%�pm�d`J=�L_=�.�=-���a�û/3>��=�c�<\�	��	=�+.>?��=XY?5�?� ��Q��'�u����g붾��>n��>�k�>�o�>�m�=O�
��b�"wG��"	��?�g?���>c��ܮ�=Gy��� <<��>N��>Ⱥ>>��?<:�j�S���R��<Q��>��?l��>�I����L�or�v��G�{>J��;Ӷ����?�`?[/���A?�����̩e�:z�%=��=���0�P�C�S��U!�h�Ծ���j ����=���>m,�?��d��(>��I��k��V���e��@�U�?¿>Е��I��꾿MȾ�h��L7>����=��>,MW>�o�>�D?�
x?�U?�M#?nS���>�S�>���>��>�?n	?�߯>�?�=K�=�&�=�v�>]�@�o�ܽI�>[���O��=�
>��>w��;ɺ;�=���SB=���1t�=�Q=�s_�q�����=i�=�I�=�8	?�M ?�͟��{�0NĽ��p����<Z��=��=0�t<5e����߽5>�(?F?�Z�>����t
����Rg�[�$>h�?��?�?�N�=��=s����d��c,>	x>%�@;��ֽ�� v��D�4��'�>ִ�>��>zdT>N܇?Y�Y?�*.?EZͼ�X(�k�y�9�I��������o�>JD�>1�/>"������wZ���j�u^G�J�ͽ����=
2>��F>ĲS>��1�Q�ý���<~7���~�6n>�>>5�>�e�>�g&?>��>��<�&��:��/�E?�Α�_��v��WѾ9�=���=�z>���B��>e�ɽ*et�޵���E��E�>�^�?�>�?��`?����j����5>�K3>>�W�R� �{�X:��Ҽ�B�=I��=���\l���[�� i>ə{>�_���澺}�����G���,\A��~��+����<���zM;٫=����Ns�uԋ�l���I���R��	w)�OKv��W���8����X? @?P�=I�< *��齾������=m���I+����6�Qv�ki��;�]��#��a���>�f�̐��|x��,�)M�%�5>S�-?�˾,-�����I=� >���<���<��!H���)��O?�+5?�Ǩ�g�ʽF�*>Z?z�>|
>���+}�*��>N�2?��.?�٣�wi��|L���x��Q�?ā�?��?S����H�����R�1�>g%?L/�>\���o��载��?��4?��>bž��پ �	?��Q?X+D����>g��>tlF>�n����پ��+꛾>'>Vd��m�� ���Kxu�S��<��>���>]�q�����$�=B�E�s���E�����~���'��+?b���❽���>*�=�C)�&=�� ���z�(36?�P�?�*?�6H?*Y����𤏻ᒒ<�?�>Q�>q,>ni��lp�>�t�>�q��t���ZG��ò>���?�H�?!U"?)�~�L]��f��w���0�V���P=".�=��2>i޵���h>���<�n���0��>�<jS�>΁>Ԋ�>��4>���=���=33���$�j���5����w���.�֩>�j�T���Ҿ)�����侬鵾��ᾎ s����Q^�1f�����M���@���Z��=���>>�>0꾼`Z�bx�{����*���c0�xپ����*h���FҾ*�:�K�!=G�轹p��]������d?Wi�=�aj>�]�>��n!�(/�>��=.��&��=g�C>���>.�S���=�lg>�PK>;�s>qW0��������JQ5�"Q�����)��!�?�"��=/�1��n5=���Y��p���<*Y?�VC�Jõ�^᣿&�>�r=�k�=�l�o�(��}>�v�>�$ڽ�;��>�?��5�ݽ�.�>�`J>{Ϻ>FX�xʳ�I��9ZB>B.?9������>�|">&R`?��?��?�F��A?��/?��y�ν�?w�>v�c>=_�>t�D?�=?�Y;?B#=I	�����Q�����n��"���&����6=�q�}Ao��>�<�(>��=C��fr>���<����	�=���>5�s?z�"?��+?�����C�_,�1a��G>��H=���>���>b�?�{?5�?'�">��3��l����t�[��>#Q=��<�H� �$�/=��>ސ�>W�`?b�.?V��5���^�<����Yܕ>���>�k�>bɥ>���=�)ĽX ��>Ͽ�-#���%��ዽ�H��/�߼�>�6�_�(8W��P%�u�����<ޓ9>;n>�g�>��A>�>��&>vL�>%�H>���=��=A�;�X��G��;/=�{����<�LF��7�:��ټmh�Ɩ���e��c��~����W����>؟�>\�>����<��;H��3������>8]�>=�m>��>]|9>w���[3򾂨,�@�����(?]vb?�g�>Ri����=s�j�����o��>2?i��>�%-�������Έ>�*�>���>.��>^]���1Y��~��?Ҿ1^�>�#�=����˓?hTL?7X�?=_�����dM���.�[=������5�zb�������B��������/yb�欷=�_�>�~�?{Z	�3)>��������O��lͫ��o�;c����>�NK>��g��$i�'��A߾�]��K��;>�ƒ>���>_}E?�L?���?��>?��?��o�G?�A�> �^>�d[=��?^��>n8�>���<�>�x�>�MW>w����;h���Z�p���(=�A�>���>>ƽ�ә=�8�>���:��[��]���!���＞�>��>ï�=n��>�]=?r�o����=�����'���.��b��z>dfL;��b�Oі>�.>��>tO?��>�<5���ž�媾�H����=��?T�?�.?�w�dD=ZG˾��=�H�>}۽�k}���+4Ͼ�>義���T�>;��>g˨���>��?��X?j�?r����=���\���Q^��6��A8�3�>�	?�ؼ>Pʝ����U��l�9X2���潴S��
[>�g�>S��>�>�<����b�.=�$�;;"��bH�+�k>t�>��>��>uI?'��>#=˽4�ƾ5�վ�I?�����h����pfоJ����>��<>&/�֝?���}������F=�P`�>l��?��?�8d?��C��?�A�\>�NV>��>ј2<φ>����7���$4>jB�=��y��	����;f?]>�y>��ɽ��ʾ�(�ǑH��׽����/���5��=hؾ!�����d7=���<�(���F��|�\˟�㦙��̘�kW����zT��H���[y?�D?H�CY=[W��w-��ӷ��.?�`��<���O�0�1��.����]�P�ؾ?G �R5��:D��n
�>�.i���u��0����$�1�!=>��>��?��ؾ����,�G�m����Z>���m�ܾvBd� ����$��T?�Z?��0��ܾj���)B�>su!?-��= ���[���5�T�?��o?y#?e�v��w����a�u��;Oa�?5��?c?���i5����dHŽ>��>�;�>��#>V羶Ě�Ck.>o�M?�^�>���>�R���_���'���?l�W?�8�?3?���>I&>��=�h��?��
�����<�">-H9�ud=�S�6M)�)�->/K�>�"9>�Nx�ҍy��I�>�[޾�L�@Z���	��g��\�Ͻ��?�p����g=fƔ>��>���}������?=:1?K��?��?��P?��z@�ʡ�o��=ͣ�>N�Q>��}>�U;�C�<^�?���Xy��s0�nJ
?�&�?�|�?�7[?L�y�:Gӿ�� ��������=�$�=��>>��޽�ɭ=v�K=ɘ�vZ=�_�>���>,o>@;x>y�T>ě<>��.>n�����#��ʤ�-ْ�\B�� ���wg��{	��y�����ȴ���@�������BГ�O�G�I���T>�'��M�5>]?W�>��>In;>Z�>��Ͼ���!>��o=�'l��j���ҾEp���=�S��0'�iؾ�u�	?T�>Q��>�	?ol>�����ӗ>B�(>e�}=�L����=�ŭ>>��>\<>�诼��>�1�>ơ�=Ͼ�i���M\��$i�2����p��u�?_R��!+�az�=����쳾҄�>Ґ>*��<��v���4�>}�=?�����q�=1v>dYP>����iI�;�:>��I�t�jt�=�b?#lv>:��Y萾�i�R�>��>:�-�c:�>�D�>�5\?�k�?�8]?8g�<�>�?�����4>���>�&�>"�>J$�>�=?��?�V����)�{|�<q���<M��"%v���9=�='=�4k��$�:����4�%��=a�=��4=��=������>��c?V?@�潇�J��!/���B�e9���s�>��3>�u�>��>8:&?l^�>L��>C�>�Qz������_��K�>C�3>��N�$�;����)_�=����PQ?�z�>88 �>��=k�5�_����9>w�d=���>i��>EWq>?�佥����˿�+ �i5 ������>���xʼA�6��n}����:�r=����c:<L>q*d>��S>��!>�>�1>�.�>wN>�4�=��=Û�){�b�k���f=��0�Q��<i���T$��Լu��n�p��Z���������d��4�
?�d�>� �������H	�sѾ,�>*��>�9�>�B�>R~�<������+��3�qR��S?��H?�>�ڶ�]�P�Ƥ*����>P�>���>f?�>�7�==笾)���x��=��>�l�> -�>���;�(Y���P�mھ��>�ݬ=����?mu?����,��s�$Z�IF�b�>���nֽ�Y��du�S��c�����3��H@=��?N��?���;:#E<�оO���p��vȾ����)��m??b?M�J=�ڣ�����:��̏�$*��;�=���>�  ?�??Dw2?�?M�I?/-%?��ƾ܋>��z>�2=���>{�8?��7?~	?��7;��>H�>��>�ay������G�S�u=Xl>Q��>�!�>���>�I>5�>��"�0r��g3�����=D�=q03=�.C>���=7��>%�?���HCƽ �ɽ7g��u�=>�{�ƻ�>2q�<�Ľ��`�>׫�>5��>t�?c��>�7Q>G�¾�'m�\�)� >d>�%>?��>�?O�ȼ��}�t[�6���Tϩ>��>*P�L6���Tؾ.T�P���6N�>��2>��;J+n>�M�?�H?q4 ?EAͽbp.���t��i0�s�Q��F:<�>�k�>�=Užn_.���o���d�O�.�s?���>����=*v�=��=�C>tБ=>>'�8= ����q�<�Ɯ����>��>�E?� ^>���=�k������xY?&@r���bZ��z�Ͼ׬H���=�Q�>y�q�Й�>y�7�Q�X�j;��׺C�>઼D,�?�2�?O?Wn���R2��J	>��>⭝>l����ڀ�8R�>��j�&�����>����6���ǐ��ƛ> :�>���>W���S���=)��6�y�v�����Q׾dC�K��ߠ�;P���;���$�ƾ׼����;`�I��R޾���jx�J!����?N�?��v?�齢��=˿o�u�,�d�����>���-r��W <�Qf>�{�?� ��(��`��"7	������x��>1�Y�O��ċ{��$)��q��C�=>Ȁ.?�4ž����>����l=�0$>�d�<ߥ�ǋ�����	�?�V?��9?���7��y�ٽM�>�`?���>� &>��������>T%4?)�,? )㼑O���ዿ�墼��?�q�?
�? ���:tO�[3��ٞ�G?�?�	�>*hw���)�|��>3?��?7�?̩�<��{�aA���?�k?��P>_��>�l�+�#=�� �s8:�Qt�d�=>�	>�h����n=���=2o�u��<�J�>� �=�\%�B���b��>'���N�*�H�����S���<5x?�@�J�>n�h>��>C�(������� i�C�L?���?pS?U8?���<���,���ۏ=x��>0�>��=���4�>�
�>�H�pr��4�'�?8G�?��?�=Z?��m�V�ݿu����ƾ�B�5d'>2޺�#�=�@�Ƞ&>SH<=�����H��>�d>�C=s��>���>`��>�|�>3���~�.�aX���j��u��A���������	�1���E[&��g���TԾ�~߽��P�p=uc�����A{+=^�y��=��?���>|��>r�>I*>&v��-���4���9��J. ��z��);������u�\�v����ejo���j��_߾B��>�W=�K=.< ?�S�<�;���>��F�3�G>��	>6�	���L>�h>�>N�>;�H>�VG=�=7�����5�Z��[B���¾_��9�l?;_%��F
�G�>��b&,�ji��t�>LD!�P�<�d},�-*c�7��>�΍�����g>��=B��=��>�K$>r�?�;�=���M�=���=yo�>GR'�1=�����m�.>��?�I����
>!��=�P?�?:�^?���?)��>Qkþ�;M��t�>P�>��=J�>��Z?l[Z?.f?e��דx���@<'_'��6��E�����4=\�=�?:�����G�w>`�<ϥ�ʤ��c�<��A>h �=���?6�>M%�?��0?r2�>�>ڨB�f�O������>��_>�S>�	�>1:?���=	��>?��V>ϑ��p��i�>�iԹ!�S��>S�ߞc=w#�>+����%?5�?��=�����V+��nۼ�R�U�>>>?��>���>�ϴ=x���ڿ܂��V(��@��׶W��ù�!� �7������ ��#���D�<r[>2�> �6>X~L>��E>��`>���>7D\>W��=�x�="��<���<���J�͹.�z�T=9M��ױ���D������W��5*�XY�rCȽ�0I� �?cK'?1�=߾�=̛��ݾ�d��Jz�>���>f�?m��>���=(��/5W��p�P��=ҍ�>��F?yV�>�T��p���R��R>�,>Ө�>x��>B��=e�Z���(��)�;f�>�l?R`�>�����σ��#w�����AJG>$��=��ͽx�?�B�?�⾟��v���gs�8ƺ�I�=��d�q3ϼ�k������8��o���hԾ�h��������>�G�?pI�:ޫ>B�Q�����'���'��ܒ=�j?�n�>���<�^������Cأ��s��u���,�=�v�=(+�>b�?Sq?��e?h^?V�?��%�P"?��>2��>��>��?7�	?͉�>�J\>�Nq>5�<�Jj�!��r����
�(�ɼ���=�t>��>�����Z�<v!'=_��<j���$}�H��=k]~<���<�ן=��=Pr>'9?��#?����^�e߉�d�B��0[>�>շ> -��"�s=>�%�=���>�a?��>��;o��������!>!;A?���>��>�w���=�v#� Җ=���>(~�;�����D�#�}�N���Q����>��>\>ԇ{>ܷv?2O?�5?{kC�J&��ZR��Q"��������=s��>��>W�>�ھ�E.�	7f��^��8���(�-�+��˭��,�=D!S>�tk>�S>��+>v"[��~���Ƈ��g��(�ν<�>|��>�z�>$�=Ԙ�o�޾18�l�N?�V}�q���h�J�bI�H�&>��=!�R�?�y�=�n����[A����>�]�?��? �?)x�1D���I>+O�><{!>���=K���Ph�������M>t$�>04����ܾW#=FL<>�<�>�ȩ�_6���8��<,�Կ�3r���8���`ޛ�_���ӑ��ʻi�>���,�*.����վZ��k���M���I ��پ�X�	����?p�t?Q52��e�=�"D�-!ھΞ˾��d>����M��ƣ5���>�W���2��Ik���þ�!�����>� ��>�sV��Ǒ���v�ޘ)�y���y�;>:0?�OҾ�y¾B'�e��=	V>�[=��rŉ��0��m���P?��5?�N�H�)?��s�>e?F�>�8>�9��v��G�>��8?��1?v��:L��@��� ̼~z�?�R�??&���B�WL��p�c��D�>���>��!?m@���5��Q>ܣ7?md?M2?0�_�w^O��)����>�??|�@���>���>D:�<��<� }�9���k�]�t�x=��p>���K���x瑽[���%�>|r�>I7m>S���,����>�ؾNN@��a4����O��XR!=+��>7,����>~�S>�:>o��`�����C_���>? >�?�g?rO%?)����ㄾ�|:=�K��U>�`g>\�[�����ݞ�>�6�>��3Io�6|(�D7�>���?��?�OJ?"c�Y�޿ۂ��]:��X����	>�%��a$=Ww,����<�KH<	ǈ��ң:�%>�9�>R�>�Ƣ>d�]>��)>�[0>�����G*��ª��t��ͺ#���*����ɾh��63�_辴
���P̾fSݼ�%n<�.%� |m�IM�:������ T> 
??��?���>Va>F->(�Ⱦd̾e�=��¾ !h�Zhɾԃ⾞@6��h�{���B���Y�%=0E���^/����>l>+M>\�>��=���=���>�Kz<O��=�4�>���=�D�=�I > ��>�f�>;;�>h4�=W�M>3q>`v��|�rW��V̾�NR>�;k?6O�=�D��S��AA��X#�ם�����>�<�>m�t��ޞ���g�>��k=�+�l=���=�٤>/�
?�X>Jq��2��������=$��=��&>O��>�*�=d?��D�RE��
�>+��zc�=c��>�K?�b?���>�>H��>'�+>�z?��	l���=�ؼGǈ>�]?�$d?��>>��=���V��;p�E>B L�L�޼��=ڍ��a�N<�e)��r��W�?<I�*=<�_��q@= �-=8H�<�W=2��<Pr	?�?M?��>�7�>Bk����t�R2w�ٻ�Nw�>&��<��>0s�>U�>.B�>�?�s>��<8Z��'��h�> �>j|H�2<��ס�Cj>���9GZ?��d?� ռÙ㾋�m=���>��>A�%?m?NA7>1�޽��K:�F����_L�V� �� ��C���C���ѡ���=y
�=�y㼮�=�?�>V�+?�	?΄>F�\>�ǹ>��?�8�=_r$�}W<��F���4��+����>�����¼�0ͽ�q�==p���V; �.����i�<�И<��=��?l ?���=�W�=�^����EՏ����>b��>�j)?I�>����a������\�����$��>�^?�J?\���q�>�^>#������>#D�>7��=��{��x����0Ԁ�m=q?���>]�>D2��3b��NM�mom�b3>� ��#��?6�?�������0;��� h��_��Ƃ�>������"�ӽ�d9�we��C!�g�����>��>7�>%z�?�́��1�=B��"<��hSX�C(оu,B>��>Ҝl>,>�PI���˾,����,䕾f�w�xzg��f�>���>�0?�x8?���?1k?Y��>
��>ᝳ<
l:?�Y>Nd_?��?�:�>�v�>��?&�^>W=�;��g������{��=vg�=�D>���>���=m
�<�:�9}�{(l��x���3�=�V�4��]&*���=��>�d?�c/?���J��Gh�=:���料��>A�>�""���N=Δ�>���=�a)>M�
?y2?�0o>yٷ���������,��P
?e ?���>�>}HX��ƾ����r�=i�>ጾ=f%.�ӭ��I�۾+�1����>-��>�C�>���>�V?�^p?��7?�K��3�����`�_�<�`>B��<��>r[�>���I�}�~��WD ��L>�6'�7�l=�;�zρ;��>�(=b1��I�>�-k�"����>@�ɽ�R>��>���>Ql�>ʼ>�,���ʾ�F?������;����%þ�ܠ�-?>atY>����{�>s�����ե��@�c��>���?���?�|a?��<�F���>�m}>1��=�J��]![��ć�������U>*��=��V���=o=�vg>��>������۾����.��zᬿ$W��������C�0�%���2�(�p>ʾy�<�,������G�����ֽ8��h0?�"�����j�s���?���?|_ּ�z�V�5�����	��U8�>�Ft��Z�����!Q�d�ɾ	I��bLϾ�F¾�;a��8@�!�N���>a/T;R��6�b����g��>�`	?�h?D׿��ҭ�g����JZ>��>q�R>c�m�����(���j�;�}j?Xt?o�	�B��Z�>Ũ>_��>���>��ܽ�$��;�>���>q,?���>��&|��	ѽ��+e>���?���?n B?�c0��;������s��?�d?q�>섣�ԗ��"oֽ��?��2?D&�>�������E�6�?�Cj?
]�\�1>�=?���>�W!��̼��W�֬Ծ`��<��>�+��^"�ϣo��ژ��a����>���>NH#��1�����>�ؾNN@��a4����O��XR!=+��>7,����>~�S>�:>o��`�����C_���>? >�?�g?rO%?)����ㄾ�|:=�K��U>�`g>\�[�����ݞ�>�6�>��3Io�6|(�D7�>���?��?�OJ?"c�Y�޿ۂ��]:��X����	>�%��a$=Ww,����<�KH<	ǈ��ң:�%>�9�>R�>�Ƣ>d�]>��)>�[0>�����G*��ª��t��ͺ#���*����ɾh��63�_辴
���P̾fSݼ�%n<�.%� |m�IM�:������ T> 
??��?���>Va>F->(�Ⱦd̾e�=��¾ !h�Zhɾԃ⾞@6��h�{���B���Y�%=0E���^/����>l>+M>\�>��=���=���>�Kz<O��=�4�>���=�D�=�I > ��>�f�>;;�>h4�=W�M>3q>`v��|�rW��V̾�NR>�;k?6O�=�D��S��AA��X#�ם�����>�<�>m�t��ޞ���g�>��k=�+�l=���=�٤>/�
?�X>Jq��2��������=$��=��&>O��>�*�=d?��D�RE��
�>+��zc�=c��>�K?�b?���>�>H��>'�+>�z?��	l���=�ؼGǈ>�]?�$d?��>>��=���V��;p�E>B L�L�޼��=ڍ��a�N<�e)��r��W�?<I�*=<�_��q@= �-=8H�<�W=2��<Pr	?�?M?��>�7�>Bk����t�R2w�ٻ�Nw�>&��<��>0s�>U�>.B�>�?�s>��<8Z��'��h�> �>j|H�2<��ס�Cj>���9GZ?��d?� ռÙ㾋�m=���>��>A�%?m?NA7>1�޽��K:�F����_L�V� �� ��C���C���ѡ���=y
�=�y㼮�=�?�>V�+?�	?΄>F�\>�ǹ>��?�8�=_r$�}W<��F���4��+����>�����¼�0ͽ�q�==p���V; �.����i�<�И<��=��?l ?���=�W�=�^����EՏ����>b��>�j)?I�>����a������\�����$��>�^?�J?\���q�>�^>#������>#D�>7��=��{��x����0Ԁ�m=q?���>]�>D2��3b��NM�mom�b3>� ��#��?6�?�������0;��� h��_��Ƃ�>������"�ӽ�d9�we��C!�g�����>��>7�>%z�?�́��1�=B��"<��hSX�C(оu,B>��>Ҝl>,>�PI���˾,����,䕾f�w�xzg��f�>���>�0?�x8?���?1k?Y��>
��>ᝳ<
l:?�Y>Nd_?��?�:�>�v�>��?&�^>W=�;��g������{��=vg�=�D>���>���=m
�<�:�9}�{(l��x���3�=�V�4��]&*���=��>�d?�c/?���J��Gh�=:���料��>A�>�""���N=Δ�>���=�a)>M�
?y2?�0o>yٷ���������,��P
?e ?���>�>}HX��ƾ����r�=i�>ጾ=f%.�ӭ��I�۾+�1����>-��>�C�>���>�V?�^p?��7?�K��3�����`�_�<�`>B��<��>r[�>���I�}�~��WD ��L>�6'�7�l=�;�zρ;��>�(=b1��I�>�-k�"����>@�ɽ�R>��>���>Ql�>ʼ>�,���ʾ�F?������;����%þ�ܠ�-?>atY>����{�>s�����ե��@�c��>���?���?�|a?��<�F���>�m}>1��=�J��]![��ć�������U>*��=��V���=o=�vg>��>������۾����.��zᬿ$W��������C�0�%���2�(�p>ʾy�<�,������G�����ֽ8��h0?�"�����j�s���?���?|_ּ�z�V�5�����	��U8�>�Ft��Z�����!Q�d�ɾ	I��bLϾ�F¾�;a��8@�!�N���>a/T;R��6�b����g��>�`	?�h?D׿��ҭ�g����JZ>��>q�R>c�m�����(���j�;�}j?Xt?o�	�B��Z�>Ũ>_��>���>��ܽ�$��;�>���>q,?���>��&|��	ѽ��+e>���?���?n B?�c0��;������s��?�d?q�>섣�ԗ��"oֽ��?��2?D&�>�������E�6�?�Cj?
]�\�1>�=?���>�W!��̼��W�֬Ծ`��<��>�+��^"�ϣo��ژ��a����>���>NH#��1��&f�>�O�L�N�U�H����Ψ���<
]?��󾈧>]i>g�>t|(�u�������2���L?���?owS?�I8?s/��vX��\���*�=T
�>���>s�=S��ƒ�>:��>lw�%er�'��ߧ?�"�?���?�_Z?F�m��xҿ
5��v���~g��>���y�=���>�0��u����4`>Y9�,/���>�Ȳ>y0x>SD�>ۉ>8�.>�#�=*��bL%��7��>[����,��%߾�nh���3��ޑ��~-�����um������C��~��=��+�S���g>��v���=PvO?�S.?z_?R�w>^��=��о�q¾ˎq�Sx��ťL��k�񵦾�;��6�J����=�]H�� ���\��4��_�>��>c������>G�ܽ� ��� ?*�8>�#�>Pҵ>d��V00>3�(>��*>b�N>*�>���=�Ė>B��>Z�^�k�r�L�(������}G>c�J?UJ>�����Ծg����ܾ��>2?Ǩ�>q�=��[��Zڄ��Ӗ>Ǻ
=����e�>��	�;�T�>8�`>p����T>>��=T�[�V�}�B�=�:�>�=�{�>��O�-�|���ټu��>C�վ`�>أ?�e?�ֆ?���>O�f�2��>�8�>=�j>�&�=g>��>�ӛ>�?��n?��?�> K
>̚��q�=M� >�ط��gl=��߼FR�ym=��������g>cH�<��փ=�r��NV�]��s�!=� �>�??���>�ź> cD�ٮ=��*D��:ʽ�GJ>�|Ƚ� �>~��>8X?�@�>��>K�E>����_Ҿׯ����>,^/>��^���m�r���p>��>o�I?��1?�h����*�W\-=,�="�>��?5&&?�)�>؛>��ν���R�ͿM������x���yW�=�7�Է��U��<�w��<>���=7�>�XTd>�H�>p(?�f�>�(>9�>�}'>1F�=��~=�v�=؞�<�"���I>�|1=2��C^>]��=)�I$l�6��ir�L�B=���=�P��/�?i�#?nC=u6�)Ԭ:1��}���Û>Jo�>�/�>G�?!t^>�o¾�}H��ik��ZQ�>��_?�	?�e�������>�ۗ>��i>�d>M�����7�^�~��l<���>Q�P?�:`>ų����Z��J����͛?U��=åI�?Uَ?	得ؽ����|�Y���B{>Wz���ǀ�B��F$��E$�����ㅾ�xc����=p+�>6��?�D�8�sDH�ƺ��\����a��K�[�XZ�yp>?[�Q�.���þ�-�P�ʾ��f���V,�=&>Ǜ�>�
�>>�>�K?լ ?%C?���<3_$?��J���?n�>���>v�?I��>�h�>�Q>�B�ږ�f����G�l$<o5���"=���=�h>A>|�';��@����=�/���4r�=f?�;V�6�ɱ�=!H,>#�A>3o?�M?���R⟾Ɉ��?��=��f>��>�6?J�n��M�=b���F��?��??z�.?��G��D��Q4�~ô��#�=SW?�>R��>��ּ����¾�{ѽUҖ=�I�>HU}=r�V��)~��c�)�}�߆�>yߎ>RI>�ُ>�#w?�^G?��5?��M��W���e�������<�:� �>�j�>��>���T7F���i�d3����^�=��t���2=�r�>Y{G>�� >�>[.>�*��N��Ө���s�������>�f�>/?���>�">��þS�+�I?������#���>Ͼ���r>�[;>���Ȯ?�t�V�}������<�n��>�M�?��?r�c?#D���	�\>�W>#�>�<��=�Z��XD��Bi5>��=�z�}4��q��;�8\>�x>:�Ƚ#�ʾ�8��H�nP��7\D���6��~�þ���y��r��="����\�hvO���ܽ������о��Z�%	����I���R��`���@�?yĖ?el�ōھ�2/��7>������M�>o{ �r'~�I�����s�����8��#�c���,����==I�W��ʋ>��׽J6���l���(��c��Q-?�ߵ�t!���(�V�@>�y>�Tʾ��n������0��M�[?G?n�*���	��s>��>�a?�o,?T��=y*�'��=�>A+-?_`??A$]>�w��닿��Y=+ɼ?�y�?�C?Fѕ�װJ�<H�ǲ>_�>*�?���>K����>H�s��H�>@�>�t�>ٝ6�����'�PmD?N��?�s�z�g>	��>�d>�"?�
ټ��+>��;�@+=8�> ٣9�mW�w:k��&:����>{@#?�5'>�1��h�����>�ؾNN@��a4����O��XR!=+��>7,����>~�S>�:>o��`�����C_���>? >�?�g?rO%?)����ㄾ�|:=�K��U>�`g>\�[�����ݞ�>�6�>��3Io�6|(�D7�>���?��?�OJ?"c�Y�޿ۂ��]:��X����	>�%��a$=Ww,����<�KH<	ǈ��ң:�%>�9�>R�>�Ƣ>d�]>��)>�[0>�����G*��ª��t��ͺ#���*����ɾh��63�_辴
���P̾fSݼ�%n<�.%� |m�IM�:������ T> 
??��?���>Va>F->(�Ⱦd̾e�=��¾ !h�Zhɾԃ⾞@6��h�{���B���Y�%=0E���^/����>l>+M>\�>��=���=���>�Kz<O��=�4�>���=�D�=�I > ��>�f�>;;�>h4�=W�M>3q>`v��|�rW��V̾�NR>�;k?6O�=�D��S��AA��X#�ם�����>�<�>m�t��ޞ���g�>��k=�+�l=���=�٤>/�
?�X>Jq��2��������=$��=��&>O��>�*�=d?��D�RE��
�>+��zc�=c��>�K?�b?���>�>H��>'�+>�z?��	l���=�ؼGǈ>�]?�$d?��>>��=���V��;p�E>B L�L�޼��=ڍ��a�N<�e)��r��W�?<I�*=<�_��q@= �-=8H�<�W=2��<Pr	?�?M?��>�7�>Bk����t�R2w�ٻ�Nw�>&��<��>0s�>U�>.B�>�?�s>��<8Z��'��h�> �>j|H�2<��ס�Cj>���9GZ?��d?� ռÙ㾋�m=���>��>A�%?m?NA7>1�޽��K:�F����_L�V� �� ��C���C���ѡ���=y
�=�y㼮�=�?�>V�+?�	?΄>F�\>�ǹ>��?�8�=_r$�}W<��F���4��+����>�����¼�0ͽ�q�==p���V; �.����i�<�И<��=��?l ?���=�W�=�^����EՏ����>b��>�j)?I�>����a������\�����$��>�^?�J?\���q�>�^>#������>#D�>7��=��{��x����0Ԁ�m=q?���>]�>D2��3b��NM�mom�b3>� ��#��?6�?�������0;��� h��_��Ƃ�>������"�ӽ�d9�we��C!�g�����>��>7�>%z�?�́��1�=B��"<��hSX�C(оu,B>��>Ҝl>,>�PI���˾,����,䕾f�w�xzg��f�>���>�0?�x8?���?1k?Y��>
��>ᝳ<
l:?�Y>Nd_?��?�:�>�v�>��?&�^>W=�;��g������{��=vg�=�D>���>���=m
�<�:�9}�{(l��x���3�=�V�4��]&*���=��>�d?�c/?���J��Gh�=:���料��>A�>�""���N=Δ�>���=�a)>M�
?y2?�0o>yٷ���������,��P
?e ?���>�>}HX��ƾ����r�=i�>ጾ=f%.�ӭ��I�۾+�1����>-��>�C�>���>�V?�^p?��7?�K��3�����`�_�<�`>B��<��>r[�>���I�}�~��WD ��L>�6'�7�l=�;�zρ;��>�(=b1��I�>�-k�"����>@�ɽ�R>��>���>Ql�>ʼ>�,���ʾ�F?������;����%þ�ܠ�-?>atY>����{�>s�����ե��@�c��>���?���?�|a?��<�F���>�m}>1��=�J��]![��ć�������U>*��=��V���=o=�vg>��>������۾����.��zᬿ$W��������C�0�%���2�(�p>ʾy�<�,������G�����ֽ8��h0?�"�����j�s���?���?|_ּ�z�V�5�����	��U8�>�Ft��Z�����!Q�d�ɾ	I��bLϾ�F¾�;a��8@�!�N���>a/T;R��6�b����g��>�`	?�h?D׿��ҭ�g����JZ>��>q�R>c�m�����(���j�;�}j?Xt?o�	�B��Z�>Ũ>_��>���>��ܽ�$��;�>���>q,?���>��&|��	ѽ��+e>���?���?n B?�c0��;������s��?�d?q�>섣�ԗ��"oֽ��?��2?D&�>�������E�6�?�Cj?
]�\�1>�=?���>�W!��̼��W�֬Ծ`��<��>�+��^"�ϣo��ژ��a����>���>NH#��1��&f�>�O�L�N�U�H����Ψ���<
]?��󾈧>]i>g�>t|(�u�������2���L?���?owS?�I8?s/��vX��\���*�=T
�>���>s�=S��ƒ�>:��>lw�%er�'��ߧ?�"�?���?�_Z?F�m��xҿ
5��v���~g��>���y�=���>�0��u����4`>Y9�,/���>�Ȳ>y0x>SD�>ۉ>8�.>�#�=*��bL%��7��>[����,��%߾�nh���3��ޑ��~-�����um������C��~��=��+�S���g>��v���=PvO?�S.?z_?R�w>^��=��о�q¾ˎq�Sx��ťL��k�񵦾�;��6�J����=�]H�� ���\��4��_�>��>c������>G�ܽ� ��� ?*�8>�#�>Pҵ>d��V00>3�(>��*>b�N>*�>���=�Ė>B��>Z�^�k�r�L�(������}G>c�J?UJ>�����Ծg����ܾ��>2?Ǩ�>q�=��[��Zڄ��Ӗ>Ǻ
=����e�>��	�;�T�>8�`>p����T>>��=T�[�V�}�B�=�:�>�=�{�>��O�-�|���ټu��>C�վ`�>أ?�e?�ֆ?���>O�f�2��>�8�>=�j>�&�=g>��>�ӛ>�?��n?��?�> K
>̚��q�=M� >�ط��gl=��߼FR�ym=��������g>cH�<��փ=�r��NV�]��s�!=� �>�??���>�ź> cD�ٮ=��*D��:ʽ�GJ>�|Ƚ� �>~��>8X?�@�>��>K�E>����_Ҿׯ����>,^/>��^���m�r���p>��>o�I?��1?�h����*�W\-=,�="�>��?5&&?�)�>؛>��ν���R�ͿM������x���yW�=�7�Է��U��<�w��<>���=7�>�XTd>�H�>p(?�f�>�(>9�>�}'>1F�=��~=�v�=؞�<�"���I>�|1=2��C^>]��=)�I$l�6��ir�L�B=���=�P��/�?i�#?nC=u6�)Ԭ:1��}���Û>Jo�>�/�>G�?!t^>�o¾�}H��ik��ZQ�>��_?�	?�e�������>�ۗ>��i>�d>M�����7�^�~��l<���>Q�P?�:`>ų����Z��J����͛?U��=åI�?Uَ?	得ؽ����|�Y���B{>Wz���ǀ�B��F$��E$�����ㅾ�xc����=p+�>6��?�D�8�sDH�ƺ��\����a��K�[�XZ�yp>?[�Q�.���þ�-�P�ʾ��f���V,�=&>Ǜ�>�
�>>�>�K?լ ?%C?���<3_$?��J���?n�>���>v�?I��>�h�>�Q>�B�ږ�f����G�l$<o5���"=���=�h>A>|�';��@����=�/���4r�=f?�;V�6�ɱ�=!H,>#�A>3o?�M?���R⟾Ɉ��?��=��f>��>�6?J�n��M�=b���F��?��??z�.?��G��D��Q4�~ô��#�=SW?�>R��>��ּ����¾�{ѽUҖ=�I�>HU}=r�V��)~��c�)�}�߆�>yߎ>RI>�ُ>�#w?�^G?��5?��M��W���e�������<�:� �>�j�>��>���T7F���i�d3����^�=��t���2=�r�>Y{G>�� >�>[.>�*��N��Ө���s�������>�f�>/?���>�">��þS�+�I?������#���>Ͼ���r>�[;>���Ȯ?�t�V�}������<�n��>�M�?��?r�c?#D���	�\>�W>#�>�<��=�Z��XD��Bi5>��=�z�}4��q��;�8\>�x>:�Ƚ#�ʾ�8��H�nP��7\D���6��~�þ���y��r��="����\�hvO���ܽ������о��Z�%	����I���R��`���@�?yĖ?el�ōھ�2/��7>������M�>o{ �r'~�I�����s�����8��#�c���,����==I�W��ʋ>��׽J6���l���(��c��Q-?�ߵ�t!���(�V�@>�y>�Tʾ��n������0��M�[?G?n�*���	��s>��>�a?�o,?T��=y*�'��=�>A+-?_`??A$]>�w��닿��Y=+ɼ?�y�?�C?Fѕ�װJ�<H�ǲ>_�>*�?���>K����>H�s��H�>@�>�t�>ٝ6�����'�PmD?N��?�s�z�g>	��>�d>�"?�
ټ��+>��;�@+=8�> ٣9�mW�w:k��&:����>{@#?�5'>�1��h���]?Ȳ��Q'i�2�+�L��'�־B%#>�??Ӿ��>�7&?PO�"���Iq�꫗�q�Ru ?f��?Qp^?�Q?�]��if���%�=O2���]H?K�>���,�>e�"?C���bL���%����>�#�?�� @mV?�腿��߿׸�حϾ_��)=��=Ѡ8>a�9�-<;�q�=�L������=�G�>�@a>w�r>�C�>"3N>{�@>�͆����p/��pg����@���������E��A�l.R�>$�x#⾥jݾ�U���Kؽ`����Խ��q����eݽ��D>���>��>E.1>�S�>T$>�A��X��)�\�kgv�p=��۾&�Ծ^��`{D��-����ʾ�Ӿ���ʍ��I9?�׽N5>O��>V�T���u>��>Ҏ.�1z=�`j>� f>nS�=U��=��e=�h>8b>r�>��>�q>�Qq�a�A��T)��$>��=B�?����X���2��7�7,%��fo>���>FL�=U�3� ����.����>e̽@���.?=_�2���R> �/?����\����a�C�y�<���'�9��>��r>��=N�:���7��#�#�>7}���d�>�
�>�3?�-h?��8?x->��#?�Wx>î�>��y>���=E��>���>�$�>��'?�,?A��>T*>�6�A��=�g�>hT�����=�,T�ht�\�~�����>Ļq@Ƚ�|�>h�>�i��  >�Od�	���з=]?�>��<?� ?�L$?h��='o�c>g�П��p>�>���(?s!M?��0??e0�>���>Iȫ�Y�+��N̾S�>EE�=M�W���n���d>>��>��S>zg?%qR?Vá�h�����<���>w]q>�F?L�?��>+N�=[�|�ޒ
�Tȿ�@)6�����ν��#��L�I�������ö��﮽ִ >��>�H�>l��>t�f>�y�=��(>���>jvM>H:>�>�>%b�<{�Q<��	�	�=���M�>y�2�๽�c1�� b���󽾦i��*�������=���>�?�N�]��c�����3�ء����Z?�=?9�>?Q�?��m>�:#�m`~���	��2�1	�>��?|-/?�x��e4>2�Y>���=��B?l�>� ������a�>�����%��?>��>Yz�>�=�=�]�Bju�a��J��>R�>!ک�"��?g��?�_��ӽ,��7�'�\�͌���=X��<����8���b����U^о=������|/>�:�>�s�?������<)��Y���lڃ�YnR��s���jǽ��>�>Et���T�9�c��ھ���;��T�=�>*�>sOX?��A?7-�?n�f?�0J?��>���/?�>>8+2?�h:?_1m?-Xp?��=�(>�(,��ǀ���#��饾w�μx�½Šܼ�
>N S>�<�~Ľ��R>ֽ1=7Ö=�9��'��= o�<��m����<���=B7;>?��?P|�P#=�<4>|�>q�>�X��{Z=�k��1ľ�Ds���K>��>�2?V��>q��12�s�>�i߿�^I=��?[�>���>1i۹�H�=p��N���}�>-B]>ű0�ԥ�`朾�����l��Oc>`��>hW>A7>��w?2&?��>!ɲ�g����p~<��BZ�$ �����>[�x>������+�NV!��as�o�G�Y�!�A�=z�ֽ�Ё=H�_>D�=N9�~�>�;y=2�>z���6��i�='����>�;?*��>�l�>,Kg=�����*��K?|&1�pgu�Fح�5g���z��U�>���>.b6<,!P?��O�w�D��^ÿ?����[��?V��?��?N2R�s'�����>b	�>�)>SN>5��.m���+�<r�>�V�=A�������\~p���=��>�pJ���	�!� �l��<k����8_��u����� ͳ������&����.��nǾ}��g�!� ����ç9��PE�/�r��ݭ�֮;�@���W�?Cp|?��->��<u�2����O����=��۾�@���W����ϓ>�w!��s���0��͋M��1������>���I1p�M�k��.:�o�>�q~��R?$dپx�;tqﾘ�Ͻ@q>��w���F��x���%��[�?�y?�g?/�޾t3w�Mi����=>�'�>���>i�>sRE�ֈ|=?��>��?n?=-�����c�)��=��?R�?s9??\"�=lK�����*�U��>���>:�?yN������ޫk���?r+?�)>߽��@v�AS���??�]?�t��>J>��>�b�>y��/ѷ�.�������
���ZKo=p\:�i��R��پ��~q�=Vv�>��]>�Ѓ�<ܪ��CR>O�/�)�o�0jz���,���u���>&<&?t Q��2�>2�>Ǐ�>�
�RJ��o��[�	��u�?ѽ?�,@?s�?���8@��p߽�+x>�-���>'1�>��F�#����IC?�ei=�4Z��s)��+�=#��?��?[y�> �;�o�����}�7��{:��g=�*�=��Q>.l���[�=��<T#R�(m�c�,>���>��g>qr_>P�_>\u>��>�W���� ����}��A�_���T�ʛ\��;�<�����.���n�h,��4���x��ϼ��G���U�I�:���>�(rO��d�>��M>ب">���>�
�x#�n_��y��B��D6�9-���;�F�.����9=	�O2�] �R� ��>��=>�=�ݦ>l̙:>N)�>��=>>�*��i6i>��.>Mi�>��>��>��ƚ��I�=�]�=��w�;�x�2W�E$U�����0?�Vl���ξZ�R��W��u|���C >�$�>��>WB.�����C�l�߹�>U���G�@�u�=!��3R>��>E|)=^�����Tj���� �U֜<z/X>�D?>DJ�<���u,�Ջ޼���>�-�t�>�d!>��?��?��?��r>��	?�v�>�>���>�->>ʞA>��r>�?L�3?vv*?8��>���>O
ξ�C=�͊>����c�=�
6�Ж������=��8;~��)68>V�L>m��=l�*=�\�"���e"�s?�A?w[$?I?�;���w�󔌿3��af�>O���ؽ>l ?��?-Hb?�?�{�>:�<�u��!��`�>ܯ$=rYD�����*>:�����=<�i?���>[4�����a�g���>�G>���>�  ?�{>�$�=Q�����erӿ�f$�'"�4ς��	�H%�;ğ:���R�����+��,��{F�<�]>6��>�o>'�F>�~!>�54>	-�>?uG>�G�=S��=N7�;��X;!�E�-J=!���bZ< �P���ٻ)���Ł��.����I�AE���}�ӼKe?�	�>U�=�㍾ j2�>HJ���̾?'�>>c>?��?�Ŀ>�
��ow�\�X��sF�Dd?��_?L�?@˾P�>��>�C�=3� ?�� ?��G��g����s>��쾑�k��o�>��>"q>zc�=��G܌����ނ>�Ȉ=aռ)e�?��6?�i�������8�������J��K�o4���D�����AM羉�G��w ������5���>�C�?w"�ս[�\�~����!��9%�V��<��>�?RK�>����'��;H%�ҿ�����+--�L|�>[��>�	?�]C?�7K?e��?c��>H�>��=��G?|$[>�>?կ~>��6?��?��B?��??�\>ʑG<�k�����n�=��Q��0��=|��>E�R>CU�<F>"�]>�9�='��d������bP����=��=��C>��=�5?��(?�
>�v >��==Z� �[����=��>�p�<L�*�l}�;Ӹ�>�9!?@?�A?��>�ƾI��,%ؾ*�>:�"?��?)�>��	>t�>�z��l�2��h�=,Fp>�=#�A���bԾ�����?�:]Y>-H�>�lG>� �>�7�?�VM?T� ?�(��*��0��qT��,Y=�����=�>�/�>V =��M�*n�A�P��zR���/�Όн=AE�U�=�>���=�v1>�~�<��&;�=(=��Ӽ����@F��:�*�>���>��?j�N>Wڛ=�w��,.�x�J?������b����Ѿ}%Z�� >&�H>YA��?cx���z��`��Ȭ=����>���?̜�?��c?�@=��s�%�]>��]>h�>��3<�\G���@��	����8>"��=�X~��G��}w*�`"Q>_m>۞���jξ��ɠA��Ҷ�:l�����F�d��s���*,ɾĦ���b��󿰾��"�Lӿ�-���GOo�%���u����>��ھ����?�=N?>r��cQ'��$2�����˾q;ӽ2�j�,鈾�i������پe� ��/�����m(����M9���͵�g�ܽ�:���:��$vI�?G��T��7�>�Y��*�׽���9�� �=�dľ��"�����̏��p:=�}?=�O?����4/���{������=�>r��>��>,�$����>7c�=H-?��A?���=�x�����d0�d�?m��?'?q�̾W�����y�%��>���>���>i#۾7Ͼ�X��X��>�g?�ȝ>�
,�Cq���-�Mx#?��w?#�0�;�l>`3�>��>�Q��ϫ�6�^j����޽��;0$����� >�p���{
:>, >r�=�~������^q�>;*���a�Ӝ{��n%�~q �\B�>�"?� B�vĢ>oѤ>�J�>����4�����dϼ��T�?8o�?~hH?)?���Y�ž�G<�Y�>��?��>��1>��<����>k�>�.��9��<�Te?(��?( �?FiI?]�O��ӿ�y������L3�����=T.=U�>�����?�=��<��ʶ�<��=Aϡ>�w>���>(�W>�V@>�R#>���a�*��s��	����yE�L%��C�cу����T���P�
��y���������'A�Xo���LE�\�"�SAY��^���ޞ>��w>��>�Q�>}�>W�9Cd�%���Ѻ&��Y-���)�䒧��K �#t��m�����wк�ZѺ��"�9����?S.U>!�>�1?���<�,����>�rѼ%t>�{C>�y>�q^>گ�>EO�>�=n2>�� ���n>��!>�r��mg�f~�6�@��m��M�1?dBh�|0�Z�R��kپ�̾�/��՗>y��='�g!��K�e����>NO��)��T��	@ʼ�_�>&�>vv��B+���s�T4��nw(���L=3�B>�o>=E3t=�Tl�pT��%����>BXc����>�5�>!7Y?3�?$>4?*��<�m.?���>�i�>d1ļ�͉>u�l����>�?�G?��8?���>��i=������=��=t#��:����I��M� ��+4�p�7����=?�;>�9A>t��2鶽.d��c<�=D$
=�v�>�!? ?��4?�0B�m�a�	?�t�Ⱦ�<=�ѽ�x
?>��>Ih�>�?��
?ֹ>Hl��E�vU3��.�>|9�>�yE���j�;� >�~�<L:�=1n}?>�"?x��G!~��<�>���>��<?���>��=�`>�}r>L|�ar��� ��b>��
����=�ݾ���U�C�Xn��ž[�|����>� �>1&�>�>ͦ�>�H>/�d>���>t�y>��;3=RU=�I`=�}��$�<�.+=�d;=���و�N��=��m<�3�6����V��8�3�ܻ�"?�?%ۂ�OJ��̐6�k��U)=�b�6?;=0l�>Mr�>�ߏ>v ����@��I��S�2��>G>�?e�"?䝾:��>�j�=�=��>��(>�c@�v�D�?a">u߾f.�(��:?�6!>���=�h��7��"��R}�>־�=h���L�?�x_?�1���!�pw0����7e=.�F=��E��n�����ݦ#�C�;���E"�� Z��3l�>?�?O����>��$�tࡿ
����ĥ�0hw<��a�,b>0�'>��*���ƽ�y��V����3}����ec=�Ƥ=�Yj>��W?��-?o�]?�:3?&��>f@Ⱦ�RX?�ے>�?�>fj?�K)>`�#?Xl'?|h�>�o">#{��Wf��fV���.8���n�g�D;��=t�ƽ.
=
'%�j�> ) �j�a>�ٳ=an������ۉc=W%�=�ʀ�2<=s�>p�?�_,>fI�>�ܼ�����ٔ=?���>�ڼ���<ΟC���:Z��>�G?<�?�u'>+�� 3�D�ľ�|1�"4�>�8?�i�>�f�=�ݿ>�Zؾ?/	���>N�>��Ծ����{��u�p���'�d��>��9>�={�y>��{?ǎ0?�\?;G�C\3��,i�SV��)��V����>h �>��=��Ѿ]b1��9t�1�a��'���<�L����=5%>A�>�T�>2>�@=>�`]=�B@�ZA���&'Z� �>m�>T?�=�>=��=Qͷ����I?ʂ��Rs�u����ξFi���>}�=>�,�+Q?����{������<����>�r�?Σ�?�d?�D����Z>&dV>P�>D�<HB9�����i���95>��=��w�������=;�
Z>��{>�TŽl�˾G���B�����V�����p�M��Z��A��V��n����0
�<�<�([�������@%�֦��e�Ǿ��k��+���x��@�?�j�?�Ԁ��(l>����ݾH����>����n�Y�����7����c�-��uH������]��y�Fo�>�Â=G��)$��GQ0�;��.���W?!�����mcr���R������@��?��������%��U�W?=�1?s񮾱��� !����;�H>�)?��>�T��X2�>);�>��O?��[?�X<>�b����i���g>�I�?}�?H�;?���=C�L$&���<�$�>���>ѓ5?���7�'���X�<n?�I�>�V�>? �U��

��7?�?뻾��=��1?�o�>66��V�{�C������Kȫ=O-�tv8<I�<�h(����3)�=Bx�>�D>�v��WF�����>�9�O�N�_�H�S������Y�<7�?����0>i>�6>@�(�g��7Љ��;��L?ʕ�?�S?Bf8?�U�����pܧ�k�=��>zŬ>q��=t��"�>���><b�|r�X�5�?�H�?i��?�MZ?C�m�|�ѿ����`Ꞿjî��=f&�=^->K�����=}l<�������$�>�1�>;l_>��>.�M>��;>��'>����&�қ�Á���M�<2��t�3x�����f�y���X¾CH˾����~Ƚ��3��Y$�@���Z�=����h>#Q�>�J�>>�>T�=��s>Q����|žl�̾���^���Aվ�H����Ͻ��j��a��Jھ@؊=�zѾ�O�>!��<� >=��>�p�=��H��~A>��>�͋>&�	>MA�;���>�Ї>.>~�s;��6>N��=$)�>v��>$g��Y�V��=.����=��>ɱ����ؾ���%ľ������>�̟>s꾐��'<]��r�>�
0�:J[�7��b���X�=���>3di>�,��[,�������=��=���>~�,>�e�=ؿ	��Q����<�ў>��ž���>ժ�>Z-?�s�?[J,?�B	�w�\?���>���>���>`y>`�>t��>�~?�#?+P?���>Ϊ=)	���,>���>nz�����[�ie������D�,2���=��b=��>(�꽄����/�>�B���V�?%�.?x1?qTE?a>H���V�8�龜�>��=�?m� ?ľ>)��>p4?�W�=��3>Hy���ھ�}�>��E> �R�MR�	2�>�ӯ>�����?�[�>J;������I=�0��\�7=]�?ܞ?Q�=�,>1Ҽ���`��gP��>2��?R���F��ݽ�:ýC.<���=�~q�6��]Ӄ=��A>Ұ.>or�>�"�>}b\>3Q>P2�>��(>^��=K�<8p>�����ʋ4��䠽hJ�U���IԼ����*:�X�Z�$��|����F�`p��}Խ�%?�?T���U���X��3��{�����>��>W(�>���>'0�=ؔ��Q�Y�<�_9���>��b?���>��C�CR�=�μ�<� �>)Ϊ>��>nŧ�����|E��׺/=֏�>�?-��>�����V��l�=��z��>��>�d����?��?��*��9_�������Y��,ؾh��<�� ��X�����м��4�j���.���z�=��>�z�??
��u] �#�H�-]��nN��s�� D�A^��e�>b�>5�k� vԾ���7��/	J������>y�>�?�>#PS?�>?�N�?#c�>@��=V6M��� ?>'�>�J?+�>Բ?=7�>��?��>k3??ȟ>�zS������)�������=>>'�>~b�>E�>+�I��9\=@���i��3e�=����~�J�=P%>���=�G>��>���>��½D��F[�=zW���>>X>�>6�	>���S����>��=�y�=;^?��?�S�>�����D��϶=�h0?��>I�>���=ئ�=O���Ű>Ag^>$:>����;���6݋�Ԝ뽥-���[�>�>��>©5>�[�?�Y?��>�cW�N7-���n�<�O���ڽ�t߽%��>��>�/9����v���7H�O�J�E�)�J�&���f�J�9=Z�=�?>{��><��< �>��S�Ct���)�)�,>�8|<�u�>�	 >��1?Qj�>ʕ*�!A���?�F?C���x���<���@�����F�$>p-G>*�ͽ�P?M���x����U<�g��>���?���?<_?��J���>�X>}�l>�	>���:�&5����b�f��$O>?�=�<v�=n�����98�X>��q>7���ž(㾀 #�o@޿�݃���(��.���ʾ-1��:D�̈����۽���I��u���A�������:����	=:ሾ	������Jp�?H�?p��0<]��6~��{�6��=D|Ⱦ�8�F:(����-4�6q����m���x�ԚF�!���>��ӽ�꒿y�XsQ�E˪=��%> �T?�wD���y��о�B۾8h����d��2����]��N�/Kt?��)? �W�7��O"�&�C>{A�>f��>�7k>?���5b�����e
9?��R?��=Pi�������.,���?���?�)?���v�m�Z`�_JG�y/?M�(?ek?'�����b���a��=YCI?��>
J���g��<�c�OJ?T=�?�����>��-?y,=u�p�憟�Ș����ӽu%X;�}>�,�<��<�}u�����۴�<D	?�W�>Wt��W��b��>�D��_i�6V���vLd�B�->N	?H�����=�En>c3#>��ꦀ�����5~��?!�?�_?�2=?���,�#�B�a�[>��>z��>�,M>-�]��G�>���>!��ΦA�B���?�?�C�?�Yh?%w�K�׿�>������u�վF��=�vk=�a>�i��5 >$�@=d��Ez=r,>(�x>tT~>%>�>ow>r:>��)>������%�+���泞�7PF�U�"��}���d�er��t�
��ͺ��m��	'���E<�5�u�{�*�N,�h��h��u>z�G>�	�=�J�> ��=+f�^L��	�'PӾ��Pt�����n!��xɾ̂��1���t�'^�TK>��UY��6?��!>Vm=>�p>���hރ=p��>w�>�6�>���=�HM>�q�==��=2>�}f>c� >2�v�NXY>�fJ>��a��BP���U�␍��!�=��-?i�9��?���B��uX�����>��>��>�n%�־���@f�DS�>�{���.���)�īL��a>�T	?�,h>UA��$�<#���m7���罏��>��H>�;�=�!�3���e�z$K>���Q��>F�>!�7?��?k�?�(:��72?b(�>���>}ݓ>&�?Aa�>E�?��e?�΀?���>Ur=a�>B���<���>�־��q� d=�D;f�Yp�|j�>��(�O;���&��>آZ<�^��|�=V�<����S�>�	?C/	?�1?ь=�/F�� D�����.[>�.>?�>�p�>:�
?�?R��>%`>
U��$ݾS�>�pj=��K��\��d	����>��>�Qh? J-?r���5��^�$�h��<%?�&?��%?(�>oP�1M��,��e��a�!�Β0�r,彅#D��~���SD��;9	j=�˽$i����>=pW>N��>%[�>��n>�B�=c+>�I�><>`>�Z�=M�=Y�կn<�O��mG#=r�|P^�]v����Z�ý|���0͂�	j����鼌�W��G��M�?��?�0�������d��?��h��}��>mi�>���>���>��=e��.V���@���L���>��e?��>#�<�v�=�`�P����>:u�>��>λV�p��~���<{��> $?�w�>ow�j@Z�ZAn���
��!�>��=8ah�J�?0 �?Z�-���1��e��<Ǿ��>Of�j㚽�eK����*�7nX�бO��M�W��ks�>Ӭ�?�q���J��帨�v���������g\�<5�����>���=�-��A��~.��O���ТD��[�>�&>�Ύ>x�9?�Q?��~?��?A�>�1� D?�=9�?�4?2�Y>�RM?<?Y��>a=?�Q����p�8D��tM�D��]��>�>�f>���=�09=v�==�w�
�ٺ�=�����<>C�
�o�>uХ=�G=��>�?`�=�ǡ>,/>�N��i˒>Ъ>��>X���R�����~!����>��J?�1?)�>F�i����8��>��,?��>V4D?���>K/�1����>�{=3�>U�=z�?=�ܾ��t��>ɸ�=�y>v�a>>OG>�zk?V/?ט�>"")=u�� ���R=�{�p<���ǎ>���>��.�3�Q�3��^5@�:�����/�=|.�F��
5�j�>S-=�l��.2+=���>�Z���0�$)��i��_/>Ov>_�>�X�>�v>���HP��OF?�g���k�e1���D̾T] ��`?>`�4>�6���>���x�C����2���>��?��?ڥX?��]��`�ǂO>ݙ[>M>]�x���K�ʲ�-uh��/>�=�1��Q� �V<]W>Bs>Ch½9��U��5� �E�p%���=p�AJþAj�����< z��t��)��=>$�3��ӵ���u��E��U��7�ﾆ|��T�?�tp?���=3�>3�����ڻľn��<�Eھ�w|��r[��XL�Of���Ҿ�#��e(��w]�������}>�/н~�o�=�����l����<x*c���/?�ŷ���I��G߾���*2j� C$��,.��.���ꦿ� �=__r?��q?�7�Gw�阊�L� >�.?8>J?B}@>s�Ⱦ�b>w[�=�i<?�G�?�T�>����u�6I�N��?���?ĀJ?P�2�c����7F�%��� ?v�=?��?��$���>2��0�?O�>?��>��`�ǔ��٦��&?�=�?LcɾW >HC�>v3>GD��+[���}��ӥ�[��<ҽU����v�<v��z����3>{P�=[��=�b�2L1�@w�>Q��Y=��"��ߞ�㏊��@�۹�>v�Ѿ��=��+>���=�v���|Ӑ�+���x?'�?�E?��5?�Y�'?��ʽ=e_�>�?n$�>���>!��=�3>Ek�>����Q`��]��F?�@-@ȎL?<�W� mٿK>��;���F����=�o<hxt>�o'���=al�=Y�=��\=��>>1��>h�u>M%Q>�{�>�v>YM>}����	&�ɚ���ۚ��WO���2�S�!�������`S��>���`�y����p=��,�Kw��2����3���C@��s>���>%�>��>��=���=gUA�D��l�w������H�d&��5��Q;ұZ�`5�� ���>��佘Z�!��>jQ�=��g>���>�=��e=FV�>\���4>�j>��2>�؁>K�=�F>3()>��=rf�;=۵>Bӹ>���%Mn��������ܦ>	�?����]�� +��oپ��,��:?�>?�y���rZ����s�]�>;н��.�<�-׾���=ň�>I��>9�>?� >�f�=����̋
�*�&eO>\�5>I��*W�=_Z>��>Ժ�>�N��hP>S��>�R?	��?�$?��B>z�A?���=/k>���?�=�m�W�O��8?%�[?�L?7v-?�ꞽ?�l�%�=Dw�<F4޽�b��)��ȗ��?$�=�>��>w��=4�1>��=`��=�F��rн�)GA�1-�=0�>0�1?`��=t�?iY����4���6���ξ8`�T ,:b>�>Mk#?�Ҥ>���>�Ö>g������7���"���>2ɯ>4�r��v� ��C��>R��>0�k?Wk?�M����d�rH�h��>��?��?C��>�~�*��9��#���/���f��y�ғ�� ���Ц�����S�4�߽�½xO׽'N>v��>>��>�A�>)v�>��>67�>��>_9�=k�=>���!��� /�xP>���;h:G<��L���.����m=��h�(�ּ��^�̻u��;j%?��?�=��a����LY�D����D�����>�Ұ>��>�R�>,q=����U�@�>��#D��d�>M�W?e��>��3�R��=�Cy����<_��>�ԓ>'<K>j�@�3%�����|��Ѳ>�6?s�>_�N��nN���h��P�w��>��<�7[���P?�F?�����������H�5z)�2��>�e��ˊ><��J��U�������~J���8ƽcO#?\v�?	�󾑰9>������"Y��'�u�k��z>}<�>oN?����nS �i!����ܾD�b��qJ>u�?;`?��	?1�R??35?���=*
����-?��0���E?���>LL?0��>Zt?\� ?4"�>�z�>���,�0���9��=,&��P >�N>>�ΐ>��>�=:�=K�<�R�?xT���ı=q��(7�=$�:>ei�>@��>ԥ�>��������}��l��mD�=���>�M�;�[�=}�o�����6����	?�n.?>
�=� �">־��%�������;ؽ?�f=?q1?�����ƫ��s���پK��=Lz�>��:�W�<`����B��x#>���I�>d���sc�>q�m?�+E?3??��ݣ�?�b���?�%��]'��>�ۼ>ek�>����NN`�#K�v������\�=b��=�$A>��>�(>n(>�{ƽ0*&�˾��Vb��z�=!�<�A�>���>^�?BZK>�z�=��Q���7�I?�ǡ����v��m�ξ+���>��B>����[[?9
�r�|������;����>)L�?���?
�c?v�@����vY>�Y>ս>L�,<��>����:���\3>��=*�p�{~0<�lX>�wx>�BŽƼɾ�S㾕�B�Xa���%K���Խ�&��QΝ�\"����w��@E��!�f����������
��є�a�_�I���l�u��@r��k�?���?>Uj>��>B��>n�=+���f&�	-�w�Y=�4ξ�,-���"�9���A��;Q���U�;T�	� ��>S��0Y����l��-#�b�����>�W-?Ap��{���ռ�:�=�c
=V�2����i���,8�٦I?82?��Ӿ�/�����t>�!?w�>j�>>B�ξ�貼��>�#?Ҍ?�����␿P�������%�?���?��:?�e��M�#��p�*�m��>�)>?�T�>�ż��Ս�5�n�Ş�>s?�%U>E.1�ka���2>�;��>RZk?��-�-�>�g�>���>V���拾�Ɯ�85���� ���>��z���1�)���h��Ge�<?��>�.2>��������>��>�6�\�N�	�H�D��P�����<��?��1>4i>�A>�(�`���͉��$���L?8��?M�S?Tf8?�_��R��崧�O��="��>&ɬ>���=;���>3��>;W��or�|�)�?1I�?���?�ZZ?m��w㿁_���蝾�� �u=?؋=,=>�G���=����ޜӼ��@��/�=�->��:>lE�>�"i>�}>Y�e>s����'�>���i�I�����(�����b�O�X螾�������EUҾ��}ö<��=d���� ��STe�ɶi���>�J?ʧ>cm�>���=�+>�,B�q`�%�l�[כ�L����T���þ���}�ƽ�����T�H���*�"��x�?o x�X�x>.?�y����=+��>spE���>�5>�=HK�>�9v<�=Oj�>@q�>-��=�.�>�S�=Mt��+0(�b7M�y�M��3> �V?�*����m�o�
E�0����!?��?�{�����Zj��,+�>5�(=0 ��߾W����>R��>!�>�C>�����NC��b�BD>F�>���	�[=Nս��K>�l�>����&>�-B�"3@?#f?���>HY�>+7�>��>�G?�g�>��t>�87>g��=�?�j?ReI?��?M�=9�Ծw��c9>?C�D��Z��
b�=tN>O�>�.^;^HM>qs>T�o�v�|>Y=�-��f>k^�>qe�>�V?]"=�-?\�����O�`�Ra�����Kd�=�P�=��>��,>?�?HA�>aȘ�Wk��/
��B��l�>bՒ>8�Y���e���W�q��>��>g�h?�)X?;ό���Ⱦ6D��Rǽ$V?P��>w5?�6�>��q�#!��B���S�َf�3�8�΂U�?,�<�,��Q��m��Y*q����W�o<=�H=��>���>���=��$>[m�>g��>A�~>Z��=��JŞ�Ϣ,���T����<����=9!(�m&_=N��=a��3�<�TO�/-�]3V�q�9m?>�?��W<�{��N%����g�>P��>��>���>�u�;{���Cg�ϵ6�ķ3�fW>^p[?|�?�W��63>B�+�>J½��=�T�>�54>T9��k�� '��C;�*�?�q?b��>��>���a�"']��75��i�>��<�F-�L#�?!b?�����'���#�<�8���	��y>�/�<��=_hH�9	Y��4�G�	����򩌼/��=�i�>�S�?qᅾ�ES>\����0��@�z��_�A~H��q��L��>y�=�_�i!��3�#+�7A]��k�=��%P>��>o??�;0?Z}?r�<?l��=�4�h*N?;Lu>��?I��>��_?Z��>y�>=��>� ?&��>gG�=��#ܕ�~�B���=n>�X�>1�>��Z>t=�>��]=b����g�IBn�΃=3�=�4>��]>��%>�-�=�z�>(��>�г��;��7����t���s>���>{�>�c��
s�V7�9����>�A?�>�Y�=���J���o従">�/S?"�?">?v߱�p]�=zU�����C�GӰ>u�� ���c�������=������ ?�D>c�>2��?��p?&f+?�'�=������r�C�����>g?B��>*�>���/_q��]'�}�L��Wʾ��������=�,1>oP�=�r>���<q�����ڽ��̽�]>Nq>�0��'�?D�>n�?6d�>�,�={�������I?;>�����rˡ��$оUM�B>�`?>���?�
��7}��ߥ�̶<��k�>]*�?���?�c?�sB�r4��\>,MV>��>�� <��?�q��Æ�L3>�H�=L6y�?x����;�[>ay>+^ɽ|F˾�b�d�K��}��LMN�c�gq��D������e���c��I�޾ɋ�=�S߾.B���Bj�͓���N��Ҳ������4pľ JW��9�?>r?�9����J>C@��x�Y�Ⱦ��/�޾�U�=8+�����=�a��̥þ懹�i�I��2��MH��K��+�>�&T�X���J|���'��피�A>�>/?x�ž	���%��v�^=��>I�<���#���	������GV?�9?���=�����꽼�>��?E�>�Z#>g���vS���>�v4?�*?'�鼾���n<���#^����?��?$�@?��=�} ��C��kp�'q?A�W?�s�>��ý���v���4?&��>��>T���J��M��l>�w?�86���+>-�>b��>��;���ݾ�o���%����c�8T>�@=G7�w$
�(������;�>�`n=-G��E����>܁��G�r�E�y��	a(���;���>����=�?q>ك>��&�MJ���a��Q��bBH?�Ӱ?o"S?�k3?͢��]��I���D�=�ݫ>�;�>c*�=�����>eN�>֎ݾ(�l�ٳ��?�d�?@ �? Y?��n�+������Y� ��߇��'=)KM>�_>�½��P>�5>���=Mv=s�=M�p>b4s>�>��?>�8p>��>��|��*�p�п!��B�c���1��[���q�m����U��h*���¾�b�� �(���2��;���я�:m���!'�x��$8;>�?���>}t�>�~�@f�=q���'5�PY�d�(���Ͼ�c��N���^:�al�*��k%¼y�c�?㍽A��<�>��(���={��>Fϗ=o�>fo>r��>Z�z>�v�>B7>�ٗ;��=b||>���>]��>��u=H'>]=7v�|tW��;i�z�?��W�>��F?�o�����C\�	�⾫���p�>�?�hW>�s뾟᝿��V���>�T�=p�K���Ѿ�)!�}�?���>d��>x#>��� f��	I�=�Q<�7�,>��2=s1�=����R�<�U>��?���� �>�>��_?���?�@�>ơ=�?�ɱ>L7?̮�>Pz?��>�y�>P�5?��U?=QJ?���>�3>�.%�Ѫ�<���� D!��@��ް<�R >R�Ž�>=?��j&/�Q�<�"��;�>�M.<���g����=3��>h�!?>�?$?F㊻��$���w�#Y�L3*>�#�>-G?V�?��8?ڈ?���>Ik>��=�`���LվA�>�� < �t�R9"�G�=Cg�>y4�>�(H?�MF?���_���ǽ��>��>H?B<O?Q�>��>���6=��ݿ�"@����R;ý7������mE��[7�Q	��,�����̞��W>=�^>��>��$>�o�=aV�=(�>m$�>��>��=X��w~�\�IA����ǽ2�����z�5"?<�*�:7�Q��gN��rĽΈ��L�&�:�/y ?@i'?�q�k� ������羴&�Zũ>&�=�"�>���>�ü�:!�@�e��iL�)��s�3>jiX?��&?�}����=~���)7��|�>���>K�h>TM�<\@g��{�E�-=�k�>=�?ł�>��ٽ��k������2���?���<Dp�-��?�M?ƵϾ���(8�%�8����w=8�M���,�]���F��D��%���6���a> #�>�?Ja���s�=�o��/���ق��z߾�
>��i�>��U>ϣ\����6#.��c���8� ����5a>9��>�>;�!?v]?�?�3@?-�h>gΎ�j�@?�*>� ?V]�>%�^?��>#(�>m?�N?l�>��D<�#��qZ@�>mD�ٞ�sC�=r�!>~�>��>>R�=�-�=��=�ӥ�x=e�/�'= �m<;ka=��=r��=�f/>:V�>�
?|���料������Y>��?�ST>�<����ؾ�
B�q5?�`?.�>b�_>~��m�9����ЮJ>�e�>aEV?��?z؄�(�I��]��������>��H�+�B��8���0���c�y�"���=Eȸ;�eZ>�l�?��o?�2?��(=R�<��A���i�:���Gg�=>�?���>��=}��)�O�ڏa�w<������=l�4��T̽�qB>��9>�{>��">Ѱ��#'޽ІI=��H=�0�=��?>H�>;�3?���> �>v��>�_�H0��@?����]��]��qؾ(+�<�LX>�'�>T}���k?��0��т����1���>(�?���?�T?7�������h>�e>af�=��Y=��P����xaY���'>��@>�����d���5��3�>�l�>�@���������q��O���DEp��������F��/��7����x,��|}��C�/��$x�d.�����ǽe��n�{��pо����y?���?���>`m�=�qX�c�Ѿ��d�J-=W͏��)9�ɾ���9����_���M���$��v�mO2��,��$�>�m��[����r��r,�5?�=x�>E
!?x�-����8���==S<�8��ܾ�G���떿��R�9g?6�=?Fi��AѾ��T�J�\>f�%?�� ?mtL>q؅��k����!>�'?L*?�]�<d�|�썊��㧽�
�?���?�-@?B�ż@�����◾A?�??���>����B�����B��>%��>�}=��⾶Ԝ�z�E��9�>�Hy?o��^�w>PE�>3�?��
�4�J���9x��k��=�`&<���_�}�
�������=0�>Vi1>�\1�=��>��>�6�\�N�	�H�D��P�����<��?��1>4i>�A>�(�`���͉��$���L?8��?M�S?Tf8?�_��R��崧�O��="��>&ɬ>���=;���>3��>;W��or�|�)�?1I�?���?�ZZ?m��w㿁_���蝾�� �u=?؋=,=>�G���=����ޜӼ��@��/�=�->��:>lE�>�"i>�}>Y�e>s����'�>���i�I�����(�����b�O�X螾�������EUҾ��}ö<��=d���� ��STe�ɶi���>�J?ʧ>cm�>���=�+>�,B�q`�%�l�[כ�L����T���þ���}�ƽ�����T�H���*�"��x�?o x�X�x>.?�y����=+��>spE���>�5>�=HK�>�9v<�=Oj�>@q�>-��=�.�>�S�=Mt��+0(�b7M�y�M��3> �V?�*����m�o�
E�0����!?��?�{�����Zj��,+�>5�(=0 ��߾W����>R��>!�>�C>�����NC��b�BD>F�>���	�[=Nս��K>�l�>����&>�-B�"3@?#f?���>HY�>+7�>��>�G?�g�>��t>�87>g��=�?�j?ReI?��?M�=9�Ծw��c9>?C�D��Z��
b�=tN>O�>�.^;^HM>qs>T�o�v�|>Y=�-��f>k^�>qe�>�V?]"=�-?\�����O�`�Ra�����Kd�=�P�=��>��,>?�?HA�>aȘ�Wk��/
��B��l�>bՒ>8�Y���e���W�q��>��>g�h?�)X?;ό���Ⱦ6D��Rǽ$V?P��>w5?�6�>��q�#!��B���S�َf�3�8�΂U�?,�<�,��Q��m��Y*q����W�o<=�H=��>���>���=��$>[m�>g��>A�~>Z��=��JŞ�Ϣ,���T����<����=9!(�m&_=N��=a��3�<�TO�/-�]3V�q�9m?>�?��W<�{��N%����g�>P��>��>���>�u�;{���Cg�ϵ6�ķ3�fW>^p[?|�?�W��63>B�+�>J½��=�T�>�54>T9��k�� '��C;�*�?�q?b��>��>���a�"']��75��i�>��<�F-�L#�?!b?�����'���#�<�8���	��y>�/�<��=_hH�9	Y��4�G�	����򩌼/��=�i�>�S�?qᅾ�ES>\����0��@�z��_�A~H��q��L��>y�=�_�i!��3�#+�7A]��k�=��%P>��>o??�;0?Z}?r�<?l��=�4�h*N?;Lu>��?I��>��_?Z��>y�>=��>� ?&��>gG�=��#ܕ�~�B���=n>�X�>1�>��Z>t=�>��]=b����g�IBn�΃=3�=�4>��]>��%>�-�=�z�>(��>�г��;��7����t���s>���>{�>�c��
s�V7�9����>�A?�>�Y�=���J���o従">�/S?"�?">?v߱�p]�=zU�����C�GӰ>u�� ���c�������=������ ?�D>c�>2��?��p?&f+?�'�=������r�C�����>g?B��>*�>���/_q��]'�}�L��Wʾ��������=�,1>oP�=�r>���<q�����ڽ��̽�]>Nq>�0��'�?D�>n�?6d�>�,�={�������I?;>�����rˡ��$оUM�B>�`?>���?�
��7}��ߥ�̶<��k�>]*�?���?�c?�sB�r4��\>,MV>��>�� <��?�q��Æ�L3>�H�=L6y�?x����;�[>ay>+^ɽ|F˾�b�d�K��}��LMN�c�gq��D������e���c��I�޾ɋ�=�S߾.B���Bj�͓���N��Ҳ������4pľ JW��9�?>r?�9����J>C@��x�Y�Ⱦ��/�޾�U�=8+�����=�a��̥þ懹�i�I��2��MH��K��+�>�&T�X���J|���'��피�A>�>/?x�ž	���%��v�^=��>I�<���#���	������GV?�9?���=�����꽼�>��?E�>�Z#>g���vS���>�v4?�*?'�鼾���n<���#^����?��?$�@?��=�} ��C��kp�'q?A�W?�s�>��ý���v���4?&��>��>T���J��M��l>�w?�86���+>-�>b��>��;���ݾ�o���%����c�8T>�@=G7�w$
�(������;�>�`n=-G��E�����>A�0�N���H�������oƏ<��?��t>�i>L>�(�I��
щ����L?���?��S?�e8?�U��_��,���V��=u��>Nˬ>ݭ�=���F��>�
�>'X�6gr���`�?�F�?���?kbZ?X�m�[�Կ������5���r_�=�8�<�4 >�釽���=�S��
�Y�>��w>�$>TQ>�-r>9�>��>��>���^� �����K�1�7�$y*��R9��h@��:��᩾�x$�qi���q���F�Q<�~_=�_�ˡ��\;/=����W^�|x�>��3<��>�Iнt��>ʺ�-nӾ��n�J������վ�P��ž�2��ղ��r���i��zF�� ���?�	>{�_>���>Ն��=:җ>#?�=%U�>�\�>5�>��F>8�.=�>�>d@�>�#>S�]>ಮ>+��>۔l�0�n�o�a����}|L>�O?!�[�3����k����Z# �� �=�g�>�la��O��ņ���A�����>��B>�B���pi��ܽ�ǰ>��>�3`>�J�>�����y�8���t��GQ>y�=߉>vn=_[<��<�ѷ>r����?�7�>�$?)�g?�g#?��k>_??j�a>�3?�C�>ѱ>�d>�;0�W�*?�}|?t�g?�Y?�xM=/�g��\>Qmi>�r<����=��� |$>$]�=�_>wr����o��k��@=�'d�2�$�[=r��>�>d�>�;7?��?�c?$�C�����Y���#����>TD?Nw?_�3?���>��>6�F>51���ʈ�Z!��E�>Fs|>�;�uH�ڎ��j�>ْ�>ES-?�e ?Yk����C۽����8"=�)�>BA&?���>�=�6����׿u�:��C+��:)�Y3��chV�	Z�Xj�;�c�atd�yQ�P^����=�خ>��>,>D�!>�Lm>��>i�_>���>�_=�o���B޽w�<�����9$�[l���+��������Hٜ��ST�Hc��c�B�s��M&���
?:�"?w�<}��;�M:��ݣ��痾9�>g��>YK?�k?��B>_�ݾɻ_���4�������>e?��	?��)�	eT=�+5��>��!�>���>#�l>�ՠ����;vZ��
��>'�?`�>
�1�)�Q�C�m��T�+��>�t�=��/�nĕ?�p?j矾�j���!�C�=�f�ɾ"a#>�	*=$��;�Y��8_o�]���AȾ;x�<>vk�>��?��b��ko=#&̾�=���㡿S�F���8����={*?&?�5>�3þ�|�������tþ���>�ϰ=k˵>��(?n ^?��k?^*S?�}�>t;�By><�~=�G7?[^'?�2L?	Q�>���>}�>�>�ǡ>A�a>_?���H�`��=�@ǽ�j]>��>n�H>��>q}�=l�G<��,�\�`�*%��r��<]Fj>�۟���S>��y>�I
=�,?��2?����<�S!��{��Jӛ�2��=�\>A���������a��1���*?Y�-?����ð����վ���{��@�UA?ׇ;?,U,?� s���==�ͫ��9�p>��>��=���;Q"���5D�n�&��R�<e_?aZ�>�%W>i�n?Y(?��)?�J>�r?��p���	N�+{1�:�3>+�>��>9x>J�f�� �h+z�2�j��j����d�+���o=ޤE>�r~��>��O�%5>)Q�=�R��+A�<#R�5,����>��>�r?�	�>��ּ���q%���I?�����L����5о���@>��<>��y|?���4�}�����A=�x3�>��?��?9d?�C�E���\>�V>!>�S.<�K>����A��M 4>^��=��x��啾�d�;f]>�"y>�ɽ�ʾ��㾂�F�(~����4���I���ak˾���TG�^�9����DL������l��.�������(9v��d �j���g�-��?$��?H?λ�9a�!j���#�iH�����<s*��[�Ͻ�ƾt��<Zk�Ѕ���ֲ�k���;��(��k1�1��>M]E�����aa{�N+�Gּ@7>�y+?؅ž�7����N�9=V�>��<������i������O?��6?���2�vA��~%>kA?�"�>��>�Ù��d���o�>�5?�Z0?>釼�u��������ᦻ?��?��??��O��F?�x	�|��?�?��>}AӾ� ���?�5?Q�>�}��ꂿ(`�pB�>!�V?5fM��^a>�,�>C�>+g߽�ߏ���D������uo�7�;>f/~;��ô^�h<��s�=��>˧~>(#R��m��gp�>`Hվ�#H���1���iЖ���,<���>T@�m�@>�>Y>�K^=�8�lĉ�D?��̌U��yX?�۪?caT?�,?&&���־$v��h]>�7�>���>n��<%%���>5�>��޾$�E��\���>��?���?&Mc?�T�:Gӿ�����������=%�=��>>��޽;ʭ=șK=����Y=�@�>_��>�o>T;x>߼T>�<>��.>`�����#�qʤ�1ْ��[B�� ����vg��{	�-y�����ȴ���ȗ��#����ϓ�w�G�]���S>�������T>�?�J�>Cކ>@�<n>iݾ�vt��ߵ=�W���iI��,Ҿ�D�s˾+S ���=7Z���.���~��v����>�CQ�Y9>Jܷ>�^�=ZK3>Mz�>+	�;ı�>��>p{>��>^>�B�>��>㸨>�C;�>,��{���h��]��L\>���<�]T?W6Ⱦ��<��1�pz�9>�,|�=V5?��>�j8�'僿��V��>�s���$*��G	=�W���>�>i��=,�=ݠ%>KeȾ�&���^>���>,M]>��>Ϣڽ��%�����)��>ʏ���=DL�=�?`/h?�_"?����u&4>�k ?h�>)�>�>_0)�҉=��?�f\?��m?-�?ZX@=of�\�>!�D;T��3R��� �z-�^=3hY><�𽕱¼mȎ=������K>B�>��<�uc/>xzj=���>[�+?�?
?���T��58��`|���x>��<��?%ر>��]?W�-?'o?e��>�z1>�����5>�>�G�>����Wd{����=#��='�>�;K?Q�?���P��X2^>g�O>.��>,'?$:%?��>Eg�>��[����M��m�����b�<>�;��H��K�պ�<�	���W���x���:0w�>?/�>w��>�w�>��<>��=�>��D>��=�C%=~Ɍ�AzL=�Ѐ=<6�=S���#5�����k�R��ީ���O��?��<ԽQA���+��u�r�?Cw?R��� ��X��3��y��n�$>���>|�?7��>yS����3�g���=�bL���?��\?�?1�Ծ���=�]ٽ`�*= �>�[>��>;�:�����d�C�D="�>e=�>�g�>Z���3;X�v�[�(�;���&>��;	�9�j�?�YG?���X���EU	��Rm����wS=d,4����jD-�s�L�#�P��ܾ㲲�e&���^G>���>IY�?�pr���D>�*��@���4��i{����>`�#�0�>���=��x�Ѣw��&#��� �m�˾�-/��*�>�Im����>�a?v�h??<�?!Ή>ب?}��z�6?�?弭�?5a+?�?(�7?�?�e0?��	?t����;[��g��d��Q�=��=&M>��>bM>5Z�L=ʾ=����U��#��`_C���ɽ��y��暈=�3>Yc?���>�ZF�Yɽ�����J":S� >�O�>LB�=3AX��pW��A&;��'>�O�>i�D?��>l~�<J�Ҿ���_����$>6j?Z;?;\�>y����=��/�E9C�zKd�l��>��:=Q$��k<�p\��<)�>��>��?M13>1Ù?@mf?y�.?l~=>���j����K��B?�3=8�?0"�>g��=z��eO��~�97�Z�(��n>��k�E�'�7>�[o>. �u/g>���=L�%>�,o��4>��#���4�1�>N5�>�-(?�>�>,��=���ɼ�8>G?,�o������Kľ�Q2�K.�=��=�`��>�'?s_���	���ꑿl�Y�!߶>�-�?1�?v�}?*?ս̍k��f�>���>3�*>���b���`��PJ@���p>�2=�W��Y��~���(�>��">� /�g���vo���v������W���솾����j��6�p5r�:�>����uվ�{����=HH�����=�@�=�A㻢?� �=� $���F�?�y�?X嬾�脾.r������þ�i?�%$�[�G�w2���2!=z���v־쫡��.��.������C��k�>�̾��������&B�{�r>'>>|
X?m�����l�q���Z>h����x�=�� �!N��t
����=ƈ"?�n#?��*���>	���b?�"?B̻>x�P�����<G�����=���>���>��#�W���>���E�����?��?��A?0�꾓lZ��>�� �T� ? .4?���>6`���#&���ھ�v�>'e?Z��>���֥�,, ���?+�?����@�>�k�>$�|>��������Q�a�M�9�>$�D>��={��?7��ђ�;"�=���>Q.�>95��@,���)�>S�۾�	=��:�i���5��/�l=�-�>Ұ �
T>>���>�wC>�M�����P����P�9X?u�?[Z?�T&?�ᾏթ�*rƽT��<Dh8>3�~>�;��ô���>�>���򢃿L�K]?���?���?[�I?to�[9ؿȢ�u���@����%>��=t�=F����T>���=)��=6?�-�6<���>>Be>�6�>���>I�>P9�=��������Ϙ�F���51��$�������� �=�S�@g���Y�K}�r%����ě����a���j�鞽H��4�>�?.?!�?��><��Q������ޏ�f�i�Ō<��_�5���,z�?Q������mԼD��=�(ʽw�ڽ"g(�=U?���=��C<.I�>��7���`>�o@>��=�o�>�T>�4>���p>Z5)>�{>�cy>o��=r�>ۙ=ɦ��M`�ձ8� kd>�v�>�AP?����D�=�R�C���)$��*��>�(0?BM?��D�o
���4��{2�>�y��=���V½���<��>��>U��<�9����;G+�<�ᇾ��Px#>xǆ>���=Z������j_�<Xy�>�K̾���=-u>S�%?(gw?BW4?���=U�>w`4>�+�>Fi�=�2p>��c>d�v>�
?�x7?�2.?}� ?�<�=��y�g@m=�kD=Jn'��Küh���f��<��'�p<���O5=�I�=�<���0=��-=���;��<�>=p�>�?D?Q?ybQ?��>��_���]��g��?��M�J�+?�-?��$?��/>�?��`>�&�>�b�����r��>- S>����ǌ�x�$��Y/>��!>�Yv?�b?�����D��9e�>�4�>R�+?t��>�2u?U	?6R>>�W=y�����<?�������j�=�����r��?~�T8t>���ֵ@<�G@���X�ҘN>>�C>W�>�.�>�R[>�g�=�D�>ܣ>RhW=�܈�2�:���<���=�L�=Z�7�K���:���6�>��'>�}�;s�ż�^۽qM�k]�=�����A�>��?��K>O ��o$��N,����I��M\'>�7?�F�>ȸ�=��ƾWG_�sn�����s#?k�?8� ?[�ھ�d>����V�=��?+�>u�۽��=����̾�<*���>�)U�>��?_���R��t�bb�6)6>�p$<�R&�5��?�k?�(S��Iؾ}S:�btQ����M�2=�J���ݾ�b����R�%=a�s��T�����:�ZR>��>��?]�h=6�Q��|Խ�䈿n�i���	����;u���@}��֚>Uk۾ː��;��N������(�n�츮=Il�=5��>1�?�		?��S?�?#
?�e����?��=d��>$F�>�,?�?I�>Cne>�n>q&5�<���G�RȆ�̷��n�M��E�='�*>y &>�ǫ���^<�w�;�a<J����n9��Gq<Kxe<}��<\s=�
�=o��=��?$ ?�㸾)��Q�齊<Q>�i[>��>��>!x�=�����^�=\?�~0?Sq?�Ȩ��n&�5� �~+��Gr�>�4?<?�ć>�88��T�=�mʾ�x=+�,�}�#>�}�>���q�F�%�	�������=>mP�>w�>>�B>,B�?=�?��?:(�>�CD�H���U�z��])=M>�ZX>�䇼Ӑ1��U_���P��~(��.8�ݿ��ݽ1�N��N�	����>K䓽�t>~h.>�˻==�%�Y;=�"�>����>Wv�=�)X?}U>��`>(I��+��[�I?A���������k�ϾoS2��?>�l2>>��?�&��*{�����	�>�\��>8��?���?�f?B�<����]>,�^>��>��< :I�)=���)|4>:��=�ŀ�t!���	ػ��Y>q�x>�ν"}ɾD��F�R�Q���`E�_�7��L��͵徠�KM���9��8k��n㈾њ	�Ļ�"�-=�z�����=�G)�JH����8�?}{?��x��8<�O���&D��?��#�=}E����|��˽�����ƾ�ݔ���%�\���?���+��>�9;��D����\���R�Ul�<�+�>��9?)��'������}>W�>�P>��O逿�����!4?3?�i��㧾"{�z�>4�'?H��>i{>�+����A��x�>�R?��?HA=e�����������?���?�O?ľU;�W~��[���O?�c?��?��R�Ue!�D>�<?�6?�F?ˬ��̍~����6��>kI�?{��b_�=C�>���=L}>.^A��콾�ھ0Pƽf�?�E=��1�B1�� @��9�!���>���>r�=A�h�a��>;���6�B���3�t��p��PW<��>��L�1>�s[>�@�=�����������R����R?�J�?7sL??��Ͼ����g���:��K>f��>{{=�j[�=�>E��>[h���І�R�p�	?ʲ�?�I�?�z4?\Gy���W���
���ޱ� e�=D�t= x5>S����=��=,�<���¤�=�n�>��c>��>Q�>�W>��>zۄ�=�#��$��(&��s8I��������3��t��g���U��W�Ǿj���S�RĖ�mS���	�lw��|߳�^�>9��>C�>X�>�5=pI�=e�N�z�׾F0���U�r\<���|��p�Z��9J�R=\�I�~t�<)����u/����>Ն:��;r>I�?<��=�.�>�-0>�/=t�>�^J>z��>�$�>�=/�>�ʆ=Ѝ>�z�=��5>���9���)���^����֣o>�D?��!�������8�<۾�ݾ͢>ݏ6?�w>��?�Z	����o��?~ߣ=%\x��P&�f-T�Wx>���>��!;($>Tp�<�}|,���P>=">'a�= Cü�b��0Jw�Ө=i��>�پ�46=RBJ>�� ?%�~?�$2?�O�=!$�>!)�=�hP>ܤ>�Y�>{�>��`>���>��*?I�)?�P ?0H�=?W����<�E����L�PZ�z�^�}S���Z=���<��ZÓ=5�=��=�@q=g$�=`��<�(�<��<\j>"cT?�O?-.D?I=�=��t�:��ɀ
��HU>��>�@?_#j>f">��K=.�?ۥ?�Π>s�=��_�dZ5>�#�=1���'��=N�W,>E
�>�:?r4-?�rD���=�qW<=h>X�?R1? 
?e�?�E�=�,����
mӿ�$�m�!�G���xO����;��<���M�2�7`�-�J������<��\>n�>H�p>[E>�>�<3>�R�>�IG>�Є=[�=�E�;(z;��E���M=�
��LG<��P�����>#Ƽ�����k�I���>��;�q:ټQ��>s�&?��d=�k:
)?�M5�1F���[>�R}>�?&�{>Pj�#���~U�9C;�mн9?�w7?9,�>�Ӈ���;��F=�1m=}��>���>���=ĭ�<[ϱ�x��!(I���>ң?�Z�>�'d�r�q�C�W����*��>j7��/M�=p��?)ly?S�r�J꡾F�G���_������>Ц�=�/Ǿ��ھ�]H�}��F�԰��T�ʾ������>�*�?{��	!)>%D��]�������*�,w��\G�=	?�>J�پ��˾e��Uv��S/�X��	����<R��>h)?d�(?��^?Qe�>��>�46��?*�>lx�>��>��?�N?��?���>;��>���4�꽻V
��ĉ�F
 <����yW�=E>>~�2>{�<M'(=�p=��1=j���3�<<q*=��<^�%=Zc�=��=��">E�?��?s���7�~"\�1E��sf�=��y=� ?e�m��������Z����>��$?Q��>�+����E���z�b*? 3�>>y?�H�>6h��
���+\�Ѥ��L#�=/;�>_=���v���?���	�����W�=,ϥ>���>W�?>�w�?AOh?p�P?PI�=YTe������i��(+���>Q�E?�;�>bö��qC����Ͼ��/�8�=�/ܙ��;�!��'�z<8u@>�~�=J5�=�">���=��'�B7/��F�������>�^>�~�>V�=��3=$Qf�h���46?�&�i����|��߲��M��ɢ�=�W�=K_���?c��/�~��>��'>��=�>���? �?!�T?�BJ�aNL��Z>r�>�l=sڼ����)���g�zT*>�T>�ء����"�Ub>Ti>��D<#�[��3����T���rb��ii����L���CҾ[����O=�b��gP ��F¾ד��#��7�O��(k=��h����<�Ҿ���?�Mw?l@��yg���r�E�羵G�dQ�>cqѾ�F��3��@y+�\ӝ������<�:�ӊQ��fK���/���d>H�ľ�X���ah��&]��zg>��><�K?5(����߾J��L>t�>]�+>�U�����Є�A�н�y(?�*?şC�mE�t{����>80C?)��>ݑ(>��/��"оpؕ>��L?A?;�>$���3���6�=O�?,��?=�1?�_��C#�"u
��.�B�2?��?f�?�Ha�H��W�i���9?��,?e`.?�M��j������K?jtO?�락#Ո>���=�'�<�i=ze�$/���Z����=lϜ>��>����x^N���X�y��=#J�>��=�Qa�rZ���)�>S�۾�	=��:�i���5��/�l=�-�>Ұ �
T>>���>�wC>�M�����P����P�9X?u�?[Z?�T&?�ᾏթ�*rƽT��<Dh8>3�~>�;��ô���>�>���򢃿L�K]?���?���?[�I?to�[9ؿȢ�u���@����%>��=t�=F����T>���=)��=6?�-�6<���>>Be>�6�>���>I�>P9�=��������Ϙ�F���51��$�������� �=�S�@g���Y�K}�r%����ě����a���j�鞽H��4�>�?.?!�?��><��Q������ޏ�f�i�Ō<��_�5���,z�?Q������mԼD��=�(ʽw�ڽ"g(�=U?���=��C<.I�>��7���`>�o@>��=�o�>�T>�4>���p>Z5)>�{>�cy>o��=r�>ۙ=ɦ��M`�ձ8� kd>�v�>�AP?����D�=�R�C���)$��*��>�(0?BM?��D�o
���4��{2�>�y��=���V½���<��>��>U��<�9����;G+�<�ᇾ��Px#>xǆ>���=Z������j_�<Xy�>�K̾���=-u>S�%?(gw?BW4?���=U�>w`4>�+�>Fi�=�2p>��c>d�v>�
?�x7?�2.?}� ?�<�=��y�g@m=�kD=Jn'��Küh���f��<��'�p<���O5=�I�=�<���0=��-=���;��<�>=p�>�?D?Q?ybQ?��>��_���]��g��?��M�J�+?�-?��$?��/>�?��`>�&�>�b�����r��>- S>����ǌ�x�$��Y/>��!>�Yv?�b?�����D��9e�>�4�>R�+?t��>�2u?U	?6R>>�W=y�����<?�������j�=�����r��?~�T8t>���ֵ@<�G@���X�ҘN>>�C>W�>�.�>�R[>�g�=�D�>ܣ>RhW=�܈�2�:���<���=�L�=Z�7�K���:���6�>��'>�}�;s�ż�^۽qM�k]�=�����A�>��?��K>O ��o$��N,����I��M\'>�7?�F�>ȸ�=��ƾWG_�sn�����s#?k�?8� ?[�ھ�d>����V�=��?+�>u�۽��=����̾�<*���>�)U�>��?_���R��t�bb�6)6>�p$<�R&�5��?�k?�(S��Iؾ}S:�btQ����M�2=�J���ݾ�b����R�%=a�s��T�����:�ZR>��>��?]�h=6�Q��|Խ�䈿n�i���	����;u���@}��֚>Uk۾ː��;��N������(�n�츮=Il�=5��>1�?�		?��S?�?#
?�e����?��=d��>$F�>�,?�?I�>Cne>�n>q&5�<���G�RȆ�̷��n�M��E�='�*>y &>�ǫ���^<�w�;�a<J����n9��Gq<Kxe<}��<\s=�
�=o��=��?$ ?�㸾)��Q�齊<Q>�i[>��>��>!x�=�����^�=\?�~0?Sq?�Ȩ��n&�5� �~+��Gr�>�4?<?�ć>�88��T�=�mʾ�x=+�,�}�#>�}�>���q�F�%�	�������=>mP�>w�>>�B>,B�?=�?��?:(�>�CD�H���U�z��])=M>�ZX>�䇼Ӑ1��U_���P��~(��.8�ݿ��ݽ1�N��N�	����>K䓽�t>~h.>�˻==�%�Y;=�"�>����>Wv�=�)X?}U>��`>(I��+��[�I?A���������k�ϾoS2��?>�l2>>��?�&��*{�����	�>�\��>8��?���?�f?B�<����]>,�^>��>��< :I�)=���)|4>:��=�ŀ�t!���	ػ��Y>q�x>�ν"}ɾD��F�R�Q���`E�_�7��L��͵徠�KM���9��8k��n㈾њ	�Ļ�"�-=�z�����=�G)�JH����8�?}{?��x��8<�O���&D��?��#�=}E����|��˽�����ƾ�ݔ���%�\���?���+��>�9;��D����\���R�Ul�<�+�>��9?)��'������}>W�>�P>��O逿�����!4?3?�i��㧾"{�z�>4�'?H��>i{>�+����A��x�>�R?��?HA=e�����������?���?�O?ľU;�W~��[���O?�c?��?��R�Ue!�D>�<?�6?�F?ˬ��̍~����6��>kI�?{��b_�=C�>���=L}>.^A��콾�ھ0Pƽf�?�E=��1�B1�� @��9�!���>���>r�=A�h�a��>;���6�B���3�t��p��PW<��>��L�1>�s[>�@�=�����������R����R?�J�?7sL??��Ͼ����g���:��K>f��>{{=�j[�=�>E��>[h���І�R�p�	?ʲ�?�I�?�z4?\Gy���W���
���ޱ� e�=D�t= x5>S����=��=,�<���¤�=�n�>��c>��>Q�>�W>��>zۄ�=�#��$��(&��s8I��������3��t��g���U��W�Ǿj���S�RĖ�mS���	�lw��|߳�^�>9��>C�>X�>�5=pI�=e�N�z�׾F0���U�r\<���|��p�Z��9J�R=\�I�~t�<)����u/����>Ն:��;r>I�?<��=�.�>�-0>�/=t�>�^J>z��>�$�>�=/�>�ʆ=Ѝ>�z�=��5>���9���)���^����֣o>�D?��!�������8�<۾�ݾ͢>ݏ6?�w>��?�Z	����o��?~ߣ=%\x��P&�f-T�Wx>���>��!;($>Tp�<�}|,���P>=">'a�= Cü�b��0Jw�Ө=i��>�پ�46=RBJ>�� ?%�~?�$2?�O�=!$�>!)�=�hP>ܤ>�Y�>{�>��`>���>��*?I�)?�P ?0H�=?W����<�E����L�PZ�z�^�}S���Z=���<��ZÓ=5�=��=�@q=g$�=`��<�(�<��<\j>"cT?�O?-.D?I=�=��t�:��ɀ
��HU>��>�@?_#j>f">��K=.�?ۥ?�Π>s�=��_�dZ5>�#�=1���'��=N�W,>E
�>�:?r4-?�rD���=�qW<=h>X�?R1? 
?e�?�E�=�,����
mӿ�$�m�!�G���xO����;��<���M�2�7`�-�J������<��\>n�>H�p>[E>�>�<3>�R�>�IG>�Є=[�=�E�;(z;��E���M=�
��LG<��P�����>#Ƽ�����k�I���>��;�q:ټQ��>s�&?��d=�k:
)?�M5�1F���[>�R}>�?&�{>Pj�#���~U�9C;�mн9?�w7?9,�>�Ӈ���;��F=�1m=}��>���>���=ĭ�<[ϱ�x��!(I���>ң?�Z�>�'d�r�q�C�W����*��>j7��/M�=p��?)ly?S�r�J꡾F�G���_������>Ц�=�/Ǿ��ھ�]H�}��F�԰��T�ʾ������>�*�?{��	!)>%D��]�������*�,w��\G�=	?�>J�پ��˾e��Uv��S/�X��	����<R��>h)?d�(?��^?Qe�>��>�46��?*�>lx�>��>��?�N?��?���>;��>���4�꽻V
��ĉ�F
 <����yW�=E>>~�2>{�<M'(=�p=��1=j���3�<<q*=��<^�%=Zc�=��=��">E�?��?s���7�~"\�1E��sf�=��y=� ?e�m��������Z����>��$?Q��>�+����E���z�b*? 3�>>y?�H�>6h��
���+\�Ѥ��L#�=/;�>_=���v���?���	�����W�=,ϥ>���>W�?>�w�?AOh?p�P?PI�=YTe������i��(+���>Q�E?�;�>bö��qC����Ͼ��/�8�=�/ܙ��;�!��'�z<8u@>�~�=J5�=�">���=��'�B7/��F�������>�^>�~�>V�=��3=$Qf�h���46?�&�i����|��߲��M��ɢ�=�W�=K_���?c��/�~��>��'>��=�>���? �?!�T?�BJ�aNL��Z>r�>�l=sڼ����)���g�zT*>�T>�ء����"�Ub>Ti>��D<#�[��3����T���rb��ii����L���CҾ[����O=�b��gP ��F¾ד��#��7�O��(k=��h����<�Ҿ���?�Mw?l@��yg���r�E�羵G�dQ�>cqѾ�F��3��@y+�\ӝ������<�:�ӊQ��fK���/���d>H�ľ�X���ah��&]��zg>��><�K?5(����߾J��L>t�>]�+>�U�����Є�A�н�y(?�*?şC�mE�t{����>80C?)��>ݑ(>��/��"оpؕ>��L?A?;�>$���3���6�=O�?,��?=�1?�_��C#�"u
��.�B�2?��?f�?�Ha�H��W�i���9?��,?e`.?�M��j������K?jtO?�락#Ո>���=�'�<�i=ze�$/���Z����=lϜ>��>����x^N���X�y��=#J�>��=�Qa�rZ����?�[�`���ξ������h�H��>�o?O4�e9{�5w ?CB�>����E���M���=�Ȍ\?�߽?l�I?�/?%P��3����i:$�=�͠>f^�>J�����=�q
?�^?�B��c���%N���.?��?��@	{?�,��!J��ж�v���'��J�=�;�=X>��E��ґ=���=V-]=vcN��K">���>m�>�Ò>�hN>�h>��L>�H���8'�ˆ��O��\�+��H쾏�ܾH�O�����Z��+�0�;����X����A=H���J��8t�bb���t�=�Rv��?��E?q�?ޡ�>�V�An�����0���7��z.=�(���5�=��q����u����GF�;I龣� ���ƾq��>�g��16>�`o>���=�ę=�V�>j>H>J��>f�v>��>��s>_[�2b�=��=8��<��#>�z`=:�=�Ɓ�5������$�C�fz?5!(�@���\����Q��!d>aa?vy>ZX�}ߑ�2�_����>��s��O��/!�s�N����=$d�>q�>�I�=��;�iu�㓾q>R��>��=濼����P�w�e��=��>���y}�=��,>8.?*p?	*<?��B=��>��>0,�>�
�=52>A.i>��>U�?�+?��?�q�>A�=G%R�M�e=��1<��4���7��6j���������|�=?�ռ׹�<�<�PF=�[�=^�=�����1��K���>�F?�'?��?�3þ�[f�߿���޽�H>N) �.��>+;?n�?r��>��?�Yv>��ֽ�=�,���ў>���>�mv�ۘx�gsB>�Ɵ>_�+:�:?,aU?��=؃�S!���խ>�\�>(�&?,�$?�C�>��>�"�i~��̿�'�ρ#�$.���\��S�� E%��@������&\���e��MH=_~p>�/�>�)B>"!>y�>��+>BE�>	�>֧<��^=M�<�4<�
Y�7��=xO�� _�;+�.� ��<�y7��㽌����*��t�?�e�(�������>��*?e(�=g�=D���B���o�R���>�X�>���>� 	?JmŽ�5��sh�&�"�_q��"��>�Ua?�R>;9a��V>����M����>��P>۞�=�|����.��l���1E=]��>�z ?UV>;�\�чN�6�h�^����g>+A=�����?��j?Hs�J氾��%�#�8���)�Q���<����<��(��T.�NC������֧���� ����>ϔ?����j�=����~����g����R>�/�=tT�>�G�>�ݳ�UQ��a�� �����e x�k�>Z>lǹ>���>�w�>%�^?��?*?o(g���'?���>ou�>���>���>n� ??�E�>ǆF>/?�������(�����h�.��	�IQ=V&�=?�6>?N=�09=л�=��%=n���ֽ/��=�jp=gA�=H�=�s�:2O�`.�>��?$�����ɾ���>��A�x�=�n>c��>�M�>�L\�V����>/?�1J?E��>W��<Ap,��>���k�����=U�>ݲT?="J>a@��~���޼�'�'�z�X>v���c��[�E��~Y��b�=�>�>g߲=� �?_�|?ΥQ?�t|��J��lb���$� Vn��t�F�>D�=*��޹���9���5��A+�O���ξh���^!�I�>��P>yh��|X>ĭ�=m !=Ɓ�=�9�:#���"=N�>��>���>R��<�~��˾�W����h?׾�{$��!>�EV����VG>�?��މ�=$`
?�l>�+��%y��(L~��HB?�#�?��?�t�?oc����Ͼ��>b�>!�F>��*��*������S$@�"�O�_8���8t�1=��s>)�>�4�Q���'о3�@��qѿ2�A��ӾX�������]�(oľ��d=_[����Ǿ���`��=TC�9��)�L�;��������;��������?��~?8Q=����[�Ծ�X�������>�Z��\�R��(���k��N2�3���ʒ���ܾz�Ѿ��Wcܾ7`�>U��3p����l���޾���=�F>g7�?������t��IA��k�=v��>��=��'3{��"��=M����N?�i4?�:������)H=�m�=2Y�>ʆ?$��k�V��X��Em�>�d?!�?PWK��`��`�~�̈́$�ҍ�?=��?t?�:ܾo!Y�����X=�k{?�??��=Ŀq=^r��L׾k�,?�^?H?��-��{���Z4��ܠ>��?�RȽ�X>�>�kI>��=�:+���=J.��W�=\�f>04\>����I���a�=}��>O�f>�<�"��?+!�,%%���f[����P�m�>V�>'�i� ����>J��>�m�L���M�����7��g?ܲ�?��>?";?F�"��/��b9R<h%c<n��>z1 >�Zi��a��~P�>p.&?�ܾ�-��~7�`d8?U��?�^@K�?��h���|����o񣾚L�=@�=��=�����_�=��=!����~ݽ8(>���>l��>�{�>r�d>�ki>��J>G����+�6���.��������Õ���	��8��2E���5���9���fܽ!z�=���R�<��]O<���C>q�/?�?�>sv4>�">�]��S��0��eP������
��`ƾ�	���ɐ�i,ŽI�7���������P�>�i�=�����>U^>Rڪ>s�]>���<���=X�*>ehT>!5�>�	>(3=��=�f�<�r�=S�>��m=K2�����P����g���I�>� r?mk��r=`��`%�8w,�:X��[�?�n.?���>�˾#2����e�(3j>�jF��!�%�=�4�\��=]c�>+{�>~,x��f��4�j��H�����2��>O��=+i=z���Va�<�l=���>�۾͍(>�=�>G�?�Gv?E�<?cN�=r�[>_�&>ل>T�>��=�j">I.�>�b?��.?&0?8��>8��=,D�R=�[H> @���@����D��ry=[ ���^=}d�=~?����5=؍�=|涽Hd�՛5=�� ?�w:?w��>J��>�����-��4b�Հd;�!�>�k^>�� ?���>Y�?O5�><�w>�}�=r�:�EЋ���	'�>j*3>�s��wx�w�A<��>_6>�I?��&?���!'Q��'�=�X�>!զ>�?^K?F�>�N>��Ѽ�����I�"�R�'�%�<��1�=k#k�/lͽ,�ٽJ��=�.ҽ��T�=��><��>rQ�>��>��H>��[>��>�"O>_���I�Q��n=�&�= �=T�<�)l��e<���=h�V=$m�{W���Ҵ�)2O<_��ʺ�)�@�q?K�?X�=d�S=�`��re������>0��>�E?~�?M��=�+ܾj�7�:�:�@��v�>g5R?���>b5�P�=���mLo���>;M?%�=��>�t�=r�ݾe�:>Y�*?�|*?��>���0_��Wm��9ݾ��>D��Ca�=���?�y?8�;���c��ܹ��A�9�����=&�<�e��� ���(�9��e���N�.�g�o� �!��>Q��?Q���(��`�������&��;l�ܩ>C�C>N?觀<�k�mZ��7�髾a?����>�$�>Q���Y{�>��K?2�I?��?PK�>�.�>�-���!?���<��?d��>`k�>*?��>��>�o>�2R����{�˚�;�="��=i�=Y�>Ow>���=vu�<4  ��<�Aj�=��=�>hɗ=6�n=H[�=�#>R�(>�H�>@B?�;�^�۽dw~�~��K>�Q�>���>`r7>7�~�将�w>�>�,?gA?���>ﴎ���*�H��w����ٿ=�nP?�s<?�$�>���;hj>���n;$��<��=�8��I����پz�;�����'t>[.L>KLI�vَ=%��?�B?��$?Ɉ��ۭ6�]V��X�0��ϲ=�X�c>)?��>���=z,	�G�$�L�%�"� ��!���
�%����Ԯ�=C>�$[>��\;�D^<��<}�>�-�=[F)�\� ��#�>Z��>Ǩ�>�>�I:>Fb����ھZ�V?�Ͼ�.%������k:������=��N�� վ�M?��d�����b ƿ_v�G?�h�?���?};}?|�'��A(�>���>8�=bY�=[��񬽁���f�
�D:�=������u��<��>{�>��	�R��e����z�ƿNWE�ah�fC������� ���=����ꎾH!��щ�l���je\�Y��ч�;������h���ù�h��?��?��z�9ľ ���,��>���>�fD��*7����� �ٽN�y�
<"��G���	�9�D���E�M����>�&;�㖿~�����/��ץ>�~?�wu�v�뾦5�Z�>C��>�B>�=����u�ͅ�����3?:�C?�e��1%���P�;�;<>!�?-]�>h_h��Ȁ;��Q�f���Un?`�V?q�����Q������i�?���?]�?<\��sp��L�D��>�9j?�m\>�D==x 4<��L�)���4?�-D?3��>h�;���
08���?�}�?I.�����=��>�Y>� �y۷��i>ܯ:��ɽ�;C>K��=ò���l�>�<e�c>빣>�d�>�9������>���?��z7�F��J�5��3Ҽp�
?"����T��܌>)�>.��������T�l0C?G��?�aU?,�2?=�����i|l��<{>a��>�8>fo�ҴK��S�>Xk?�-���{��@��.?j�?R�?ѡh?/�U�3>пW&���u������
�=�w�=h�A>�����=���=i=2~Q�r�=�h�>1�>ұx>�d�>BF>2T.>�����+�{Ԣ��ŏ���;��@��}��X�L��R������վn���}��c�u�N�~����X`ڽԃ
�8�m��S>��?��? ]_>-�>ّ<8��ɏ��a
0�\����(���Ҿ��u�����ps�I5�B���%�E�p�ȾCٯ>M��bU>�/?�i;>�\���>V�>��?=S��>�9K>M��>�^0>yM><n�=r�>���=;yV>]�P>އ��4KZ���2W!��[�>$;?���>��-<� c�S��
y��Ed>��%?Y�?�W�|w���	��V��>>�z��-�עC>L`9�Z��>�m�>��x>���=N̗�3{�����|81��#m>n��>z=�_��>E%�.���s͖>>%ݾ��|>#��>�X�>s�z?��?ߥ	=G�>jï>�V>��='q�>�7�>��>���>�� ?Y�?��>��7>�#����=���= ������+Z�Et����$>���y==��=���T�<D��=�ß����<H�Ҽ?q	?�-?�L�>�Ǭ>���uLD��54��ܳ�*�_>6?��&�>L�>���>D%�>>�>Չ>>�<=��ʾ�d�����>�A!>	�U��,�J�<:��>��p=�! ?1#9?�T��lϽ�~�{����>j�2?��M?��,?��'>�~��^'���ѿ^gȾq͖�k�H��>W�>%�b>���=j�={�y�(��-l�#��>��t>m>�N�>Y=�Y���?b?��뽳|g�̂9=D7�=��>��>�= s8��"��&>#�=S<�_S�^5���� �����+=��?�?uM�=���=y���R5�#���5�>X34=H�>@�?��&%��x�J"�BXܽ�?J\f?B6�>�Z��>]q�~p�=i�/>#��>q�>�>T/�K�-�"�g������>�?�C ?�K>��#;�/�|�(��.�T>>6>2Q�˅�?�s?NHF�Ђ;� ��H�:��U��>���=��0����������>	��Q�徍򸾩Z�ܓ�>sƀ?1�<�"����������|�����t��=c&>����> ?��#��{��������B�ѽnƻ*H�>�ѥ=	�>t�G?0�5?:�?�R?�̍>ߨ����?6�e>�[�>�N�>ٷ?b<?��?|�K>ite>��h��/l�ֶ�l���Q
ּ��ѽ��=R�h>��>e q>� �<�6>��n=�>ѽ���=T�>�v&=x����=�B�=�df>��?�j�>�EA���=��%�Y�ؼ�#���>�`�>R�<�Z�tv����<���v>%Z?+Gd?X��:���9�Sx	��?��b?��L>q>2��>��6��a�\}u>ȩ�>t�ѽv�z�ڠǾޏ����	�=ul�>U��>`iS>�gf?�3k?3�8?0���қ#��Ƌ�ZQ���=qo���?~�+?�3>$w�� �!Y�,]_��S1�Dך���,���=I�>!0�=A#0>����e��s9(�=�i?<v�%=Jgd<��>�c�>T��>�*�>�>�J��v¾��I?Ml��[ʾ��ѽ�Lվ�MѾ�*���N>��K��1�>�e7>�^������HSr�d�?6έ?�'�?^�N?әx�.���� >���>"��=H_���d��GY<�<Jt����>{# ��a����㽟��=�_>@��� ���e����r��ʹ�55?�2P�����`勾Cq����@��s<�?����������vM�q�������4�nb��0������?O��?>̰�c���["�^���\�� Rt=�m��ff��0k�O
0�é�����`����̾�����p��3Ճ>ٯJ�����g�S���"��1�0?D�i?�:l��1�<O�fѾ>W;�>�aB=���Y�u�(���i����Z6?gR0?�,���a=�6����z>��?�冽�'>,b��.k?Լ�?5�Q?�9�XO���[v�3>�M�?*�?s�-?��>w��������g?�?��>�a����'�ݠ��	��{?N�?�J>~�l�?���--���_?g��?y`�k_�=�NM>]�z=I�;rm�Y>>�$F���2>"L�>+E��thT���#���=�Z�=��o>�f=A2����p�w[	?l'�gP�&3����O"��~��=j�>�]B����>j�>����Y���@ͥ�Ȕy�?��=�?�Q�?M�'?+HA?�����K�7哽�;E=$W�>�V?�ɾv8ѽ��?;D�>�!<�8�#����K�>���?lL@gV\?^�{�_����̿�Ѹ�+����>�c=X�>O�,����=_�<V�V�8����<�k�>��>�چ>`�a>0@I>�%>"��7�*��Ԧ�l暿��.��ӾR��������A	����G6�9J��a�ɾ�܆<8ej=�@�<�������}������D�>�A?�=C?�N��n�=�x>�&�w�x��	������pJȾ�gi��Ծ����;���;��
�����N7��5��Y��>�f=� >��>[�W=��=�=X�=>�U<�d�<8)>>�=�/>wt�<�0���>E{>� >
�=���H�i�:Y�Ұ��J�=�es?�=���쾺k��ξ3Ǿq�>Xif?��5>��#����c�u��2�>M���BF�l�:>Em1�9Ӽ�4�>3�v>�N�����l=Y�&�C��h�E>���>+"�=L����a/���}�%_�>�Ǿ�VL={�>�?�f?3^A?Gtm=��>�_~>i.Z>s��<y=V>�?>"`n>�B?U�5?ߘ?q �>���=��U��ނ= ��=x���������R�<e`�����<u�L<��c=�<=�B^=�\u=�=�,(ɽ�ܴ�FQd��q	?�R0?/��>q��>�Z�z�=��Kr���輺F�>g�ϼ��?�v�> �>N�>��>_<>���vJ��˾�_�>+��>ȃw�aሿ��&=��>B��=��H?��R?�{l<*��U�<j�>4�>�q�>iF?��>�>���=
���lӿ�$�!�!��KO��;I�<���M��_�7�-�����(��<Շ\>N�>��p>�E>p�>)<3>�R�>�HG>҄=�=�>�;};��E�ŚM=b��AG<��P�C����$Ƽ㟗����'�I���>��<��;ټ��L?9<?�g8<m�1�]"M��ƣ��7�Mh�>�j?��%?�?A+�=*���Hl=�6��/z����>@�?b�?��ؽ��8������q���>���>Z�>�K����	��*J�������>t�,?�E�>�jF��`��=n��� �ۭ�>>����zޖ?�<x?b�J����|�&��t;�6�����=Z=����76��������Õl�\��=�B��	��q�>��?���?r����J�L5������>�.�>0J&���W?b\?���s���o�����h��MH>\�>���� �?b}3?�/G?�2�>���>@�*?�+h��j??y��=z3
?�}�>t� >�y;?�Y�>�>���>�lB=�o ���ܽA�=����B���U:>�@>�$>W3�=�=��8>F�_>
C�;�V�=�(>w�=6��:���="�=��>_��>Q�?]m���>ZǺ=�2�� �>��>�U���Ż�Ȱ=R������,�>�6y?LŪ>������T��/��{R>PJ`?i�0? ϣ>$��9��zm߾��4�V&�=S��=��:��׸�\[�ز�!=���>��=�{>?I_=k
}?4�^?��5?�n�n�+�3;���c���H<>R���?sז>�g�*�I������+��?.���f�~g���G&��ޙ<��/>7=c���Jx�=57�=�JD><>�7���n�t�]=�p}>��>/!�>mC>�X�=LN�M�侢�l? M�1��[���g���r��]ق>(��B��^�?����9��)���sD��R$>3��?���?�0]?ޕ���?���X�>nӪ>���>����6�c��K;M�V��<��߽	X뾃J��# �����>��>��ż��3������sD��bϿf�N�hVu��о�v��35��*����TüL浽ǳ�s���]�웖���8=����X2�ɕ����Ǿ�?+-�?�Ӱ��P�c������"�W4L>sQ�<�,��V<��Bþ�͆��1��ԕ��I��.`� ��ˎ���aZ��|�ε@�}���x;=�2?!�� þ�޾q,�>zN��Z>�4A��_��ΰm��m9���K?�L+?�׾xG���ȾI�s>�6?��>y�	>m��[j>���=2@?�Pj?-�:������Q�K	>1��?A4�?#��>X����o��X�PK?
j?���=�?��<��ھ��׾a~v?t-a?;�x>%���+}��:I���?`�?A��:=q�d�*4�>G����F�����g�K>�=��=��=��P��п��8�>��>���=t��|� �-!?��� ����u-����^)�=W�>R�:�s޽/�>M�=SY�C��]Ԍ��Fn���?���?,�?��1?��4�@Ծ,s5:���g�>�g>�_�=6�S�e0�=_�.?� ���c���U���/�>��?�&�?�e�?XՍ�|H�&6��(�������J�D=S�=���=�+��Z=���<��v���=�z0>J��>�˿>I�>:2p>7�>�!>)����,�ݐ��[��H:�y�����D��&�.u!�B��ϡ�z�Ͼ�c5�X	纯R�\�N�:-���`�<�c�q��>��B?+�.?���?L:O��>�T��Y�NHᾦ���,*���ھ�þٳ��D:C������*�k{¼\�þ�ho>&�=9�<�*�>XM>��,>�o+>t~�=I��)�=�Ӟ>�k>��=G�>�q�=Ն�=9p=��>��=�R��$݀��=���T=>8w�� u?����ʀ�y�v���쾫�.=�iD>f��>��=L�&�Q0�����Z]?�L�����m���C��>4�?u�@>4�@>C�)u����<���<_�?P�&�0ǽ9�"=�ν<��=_�>�eǾ��.>�;�>QT�>Esu?��J?�*�<�=�>�=XՌ>I�=
>t��>ח�>�p?�2?Y�&?B��>.m�=+l��C��v�;����#%�.�����=@U��m�9>�T������/�=�u,��y�_��=u���/��<}��<E�>b�#?���>�*�>M����>���%�߹ٽ#�=>X�5���>jS�>���>�m�>{�_>���=�$���ϕ�g��� �>��?>�q����D>K�>�h=�D?�ds?t��=s圼�O>)y>z�>)�(?NG(?u�>���>��;���!��� ��V
�:Ů���S��!�� 1x���y��v&>�)�����̶�W��>��R?^2�>!D�>�g�=^tr>��>&�>��y=G@]<57�<:�=L*D=�$�=�o}��<w<n���f"Խ���<4q�����Ӽ��,�R��r_��C?1��>�/P<�6�6�e��_R�N��>4�1?O8�>5}�>�L�=�ޫ��F&��_3�V?����.>(s?�N7?�)��k�=(�Ⱦ4���y�>*�&?��0>����w�v�߆��j�yP�>��m?)�L>ʈ>�㔿5�n�|�-��>�>q`<�)�?�mi?�1�ڞҾۏ���E��L���J�7��糾�ӿ��|��@'���{�������
�=��=,�?T�?�-D�}��D�N0��Z������>����",+?%ܿ>R���{r��w���þ��[C^>L0�>{9���I�>�3?�o?�D?���>���>
U�<v�?�2�>T�.?ϐ?���>N�=?�6?g �>�V7>�+>�QJ>�����G^���=�߼t����S=�8='�<�s�=��=[է<="�<�H��Br�v��<���=Y}�=�Ѣ=E�^=���>Ot�>N�<��h�=�D��A��CI>5��;���=�y5>�������<H_?8C�>.)%>�SA=�����f��>�s:?2�l?Q��>.�������y���1���՞����=K�M����4��W�e$�d{k>T�s>��B>�>�qs?��:?��?��=�����G��R�!j+�u7�����>4��=��Fo۾E8��77�'x2�2�%�=������K��<��=\�P>�)~=�f7=E�%>}�>�<��M�T��6d�>���>K,�>��b>��=MC���sľL?�j��T���=�2�mR�WHJ�=g�=�ڜ�z'C�D	:=h`���a˿W�:��Q?]��?τ�?⚽? �ʾtgƾF� ?�<?E�>�P��I��tأ��hᾆ�:=$�.���#�p~�e�r>�� ?� >����L>��]F��}	>8��ˣR��&����ھGuܾ��վ��`�b+λ�)f��/;��#�ӟ��MTܽѵ9�f�S;��3��o�վ��ܾ�̪?2�?`� �I�U�4��������h�> ������_����3N�9w��(�f�;���$J��ta��t?�A<�>;~��š�z���s ���>B>>9j1?pʮ�7���2�3��b�;5�>�˽fg��������}��+���LL? �.?�� �Q^ľ5P��\I >d��>gZ>���dI���~=&^?9�;?�\�>���`5��Μ��#mS��(�?�?�&?;;�=O�~�X)���G?��1?���<z*
?��4��,�>헇��,W?c$Q?��R<��������k�>�ʽ��s?�"�=��=�B�>�K�>9�̾Q3>z��2
��e>]�=l�ٽ�V�$����މ=۱>�X>�����6�C�>����M��hG�d�G�'�p<ѩ?.��><�i>p�>Ӵ(���.̉�tn��L?���?@QS?9F8?(K��1�{���!�=��>��>�d�=�k
��>½�>� �EJr��-�)�?��?���?Z?m�(ӿ�����¶�v����#�=)��=|�>>�߽�=�N=�퐻bH7�8�>Qi�>�o>�x>U�T>��<>��.>o���5�#�����kÒ�^fB�"�r���g�Gf	�*�x�Ȁ�̴��󽾎Ϩ�M�������H�G�8t�\E=��J��oo?��5?��N?{?��>�r>�~��r���)=����0.��K��~��
"�=d=�6�=�,����/��=`C�x3�>BZ;����>�(?��=F��=��=�\��Rz>8-���� �Y>��>���>��+>�\<=`�&�>�\�7É��8{��ꇿ��;��,q??����>L�Z���JB���V���Z?�?�?q�@�cN���县M` ?���������F�j=��~>�)�>��_>��=�1(��̂=�E���/B=��>6���~"�q �����>uŀ>�w��w�=��Z<��*?�u�?�;E?O=��>��>�ɟ=y0S>���>˔> ��>̧?��N?5?���>Ÿ�=�����+=G�M�ш�o���U<�ǩ=�a��ͯ=�=�D3>���=
��=F_2>3Ђ���r�ƚ�<0@<�B�>�7?U��>P&?*,p��8.�d~h���<�8/>�)�>��>�T>���>���>9 _> ��>���<�r��vھފ?^�S>ͩ���m��h�^���<���>��^?z�#?m���)��?�>x�6<�t?ǝ�>��?Zq�>���=�
�	��������_�Ny�m�TZ>���s8���)}��$����ɽ���<~��>1�>�;�>?�[>���=�f�=J?X3 >$U�=lS.>�@�[�����r;[=F�����r>.�� ����8�\U<D�ƽ��<�� E�=~�.<d�$?��>��ս�����S���	�	8;��?��?�>A	?�">{S5�)lq��3���y�}ek>�k?��/?�<g��K�������鎏>R��>�
�>��>�o�;����g�y�>Z�#?��P>e�����*��J�u�,��Z�>�~]=*�����?$j?|&���m`���%��Q&�v�����>�m���j���˰��X���F����|:�����G��=�?��?^s���!�=������l���=��N>��5>z��>!\꼋��,��oH�"���k��z�>� ?�依��>'�&?��>t�?h?�?�'޾ �8?�=����{�>[��>���>��;?Y�>Lv+?�����������S���[���Y���J��y==,!>V� >�|�<�� ����</�;�(=`wżd������q�<n�==�w�=\��>D�?&����rX>���-p��GE9������1>��>H�ｔ@�=N|?l�|>� �>`,�>8�o= o����M�@�L���>]�R?%�W?�A?������/������M_>'9��H�������f!@��`\=q>�>�`>b9<��a>���?^l/?�-?��̽t	��}_�.@�Nɹ��ҩ���K>%�>�=!h��&#��^��A�39.��◽7��Uf�=�D=pQ}>N3>���=ҩ�=�#Ľf��<�"Q�}�˽t����h�>���>6;?���>J�X=���/(���I?����L��)��<]Ͼ�~,�1>abC>R'��0{?>��a}��M����<��\�>l��?9A�?�d?|�@�k� ���\>A�G>�>�۰;�S?��������]5>k�=�|�u�����;f�[>5n>��f�˾5�$&;������L��{B�I:]��D�]��_]徉����پ'*�=:��KZ;��ѾL��2.;�A���W ��s��N��\`�?�7�?U�u=;��=�^����[E��lý�G��؏��o����I�y����V��@��
.��S#��e1�V��A�>�Ɔ�,Б�e@z�qx,�������=!q<?[�Ѿ���~C���]�<�̢<�=�=�������}��d���م^?
�#?8m���o����=��=�u�>���>=���!ƻ�6@F>� -?՞?f�������c���V���G�?k�?KR?�"��Xmh�|�G��Q;��&m>�~�>V�?���jװ�}r�>���>���>�nD>*j澖哿�V�;V?!�m?��z��>�ؔ>���>�\=������m��vǦ=�8�>�f��=kf����6Մ>���>�8�>��d�Ez���b�>�hݾ�Xݾ_�	���j�<�ޥ�o��>������=4)�=A$6;�@I�M���*�j��9�<�hW?㺰?@+?ۚD?�V�F��4�������>r�k>iR�=��Խ|�2>�l�>l���f���i���_?P#�?b��?Os?+�H�->ܿ��������-���K�1>9:>K�>*/��`��<,>����c)>qȍ>��>��^>�PL>`|I>�0>��=�y��-�䯕��Ez�h�b�D�� �G����j��V����������D�� Q���o2�a��R Q�w��3�ɽGþ>ڃ>�IK?��?Fv?Q:�=��>�̀���A[�n~&�[FF�"A��?��oҾ6�)�}b���p��D�����o����\?�<��>��??�z�Ts��CDi>�F��US�=+kP>P4���7�>4�>��>=�?>��>7t��a<�>�h�=)߃��v����7�O�L�Q�e;�fA?{R������f0��_˾�䕾�В>�K
?�ic>�%$��Z����{�'�>���Kh��i߽�!/�<�>HS�>2-�=.S%��<�qt�*�콺i�=8�>�#>c��ٟ����
�Ms�=4u�>q�վ�(�=[2v>ӱ(?��v?�46?ɶ�=G^�>O�b>�h�>�=�ML>�P>g�>Y?��9?� 1?��>�;�= �`�i�=7=�U>�0SW�)7��9�ۼ�
-��܏<�o4�6�F=��q= <��^=��A=n�ļ���;��<0�?�?�ky>�L>hx4�R�p2���w��m1|>�;f���>���>V/	?^�
?���>�>���/�	�wd�H0�>P��>\<e��&��/�t�w�`>k��>ud?W�.?�� � ����n�>T��>H ?>2?�3?7y�>�%ӽ@�T��m����6��+��!�ս��<5��=�K��A��B��=�1Z�0n\�^�=�u>P�l>O�Q>�A>0��=)d>���>?BC>x�=/[>���o�C�죠�	!��^Ӽ�َ=��s�y�����}-ƽ��Ƚ�ڇ���ѽ~?����<� �?�t�>ޖu���.�>�������#?�p�>�3�>S��>��r�2����i�|�o�ߴ8�"�>�:?-��>�����A=HEm���|��T�>y/X>�*�=��a<�{y�Ȭ���#�=��=T�??��0>t�~�7o�ËR��&���>�/�<�~��T�?�_?���E"��~`�> Q����YV�=^л��u;�0z����Ug.����������.�+<�?���?#���֌��ӆ������Bt���u��c?=ߔ�=��?)�>�۽�ǅ�|	�>�Ѿ�$b�T�<@$�>樗�(�,?�=??w�?&��?ԌQ?�;?6�����'?�&>�C���ߤ>��*?��9?ZZU?X�>�I�>������VFL���Ǿ{.>��g}�>Co�>7H�>@�ؼ[IȽ��>���vY��-���<P<#�֯ɽ=ڪ<��;�%>��>��H?��X��V��8�"�#��Ֆ=��\>Q��>����(#-����>�9�>hMD?էc?ע?���=$��o]�N~��r�>ׁ0?/�e?k�E>9�K��@�6S����.�/�!=���=L�������^�^]��sE6�L�>Ƌ�>�tH>_Jg>�}?��@?d�!?���h/�<�u��i)����BO�)�>.Y�>J��=��ݾ`7�]Nr��_���/�)�.���F���<)��=>)>>&��=��>��=E白�&ӽ,<�������>%�>$?��]>�]�=�:��S:�40G?ç�����F�=G�����>sn�<��e�}煾�$�=��ξ8�����ɿ�vL�8�>�?bJ�?n��?��r�-�<�@S>@O���>�1!�J�i�C=�SL=\�@>��:=b�<�V����(>�
A>��������p��r���휼"�¿�[��A���ս^��
���Y�"����޾fS+>����gm=�����9����]����x�h���?EY�?]a�=#��=��`�_hL���Ѿܵ= A�� "��/B�ۑ+�����^߾��w�o�hf"��-�8�/���>P��F��t�=/D��u�p >��>+i,�
ݽ�<rǘ�GC>4��=�������鞿R�-�gg?�2?,ν�f4�pr��,��>�2?u2�>��>�T>�e�N��>���>)h<>J=Dь�P3��9{�5�?���?�O=?3ڊ�^0x�a�5�}���y>�_�<���>@��"~�@��>��>>c�>�[=>��tZ��_�P�_!�>;��?@��o�>��>���>��,�����U��R��Nl>f��>�7�!�=HL�
��Ⴧ>���>�)�>�F�����˳>��ž��I��z侚5�=���<�y>�H���8	��S����\��/����S>b�r�=��Z?-Ȱ?��0?4h\?rf%�w-�r';�)�=��>��>�q�<�H���>+Y�>��쌿n�&��7?V @��@�V�?�]Z�}�ݿj���_r���zľ'�>
�6>��>.6������j�>�`;�;m-=J�>jf�></�>�i>�G<>*1�=�	>�!��7/�a7��/���g�h��������4��8��7��U`��͟��E��������A3I��XC��J���=]���e�>�TR?.s5?���>���$��>�k��Ǣ��U��#��q�����W�����[�F�}�Q���g�$���B3���>?'��OCT>�E?�σ�%	=�b�>��'��0��ˮO>��=o��>,��>V��=t�=��_>�}>�n�>��=r�r�ǒv�1�?�'䟾����/?5��XmֽZ���I���C�N��>��?-u>��'�@��k��dv�>�h�������b��3Ǽ���>2t�>�5L>2�;�^�������u��=c�{>4�G>}:�=���c#��g>�T�>#dȾ{a}=�4C>C�!?q,x?|�=?k�>�o�>JhF>]�>��=�5}>��S>��>�a
?5�#?X�'?���>��=�K��h<%9�<ݟR�('Ѽ��7�D+���5�c	�������v<%�=<)�;�3f=�yf=�y�;mļ�'<,�?�Y ?�dU>!��='
�=�ླ�r���4�?�֗>W@?Ӌ�>��>�&	?�>��=�I�:��������>q�*>�,2�hσ���T<�$�>�+? �U?ۭ�>p�;� ξL��=�tu>��>�?�D�>�8t>Xh��x/�������ڿד�|
�׿L�J�>pkؼ@ރ�|̾
�>�4y��,@�o?�=v!�>���>��>��#>Zt*���>���>�&0>�f�>'Dq>��H>��t��ོф�=�x�K�=��na�<�ed<	�̽�K��i�q����<�u�<�ǽIx?�?D`>°{>���%�2s��T�>Ƽ�>���>��?^�p�:���9���`��ꤽKg?S D?���>�R^���S>����Q��nn�>-�=]���^��<5��򦽾O�>�%?��>�\ɽ5T1�ڷ|��!�+�=}�=="F�<!�?�n_?���9������uF��u
�-=�̽I%[�a���x!���9�&B�����k#p�PY�=�l�>EX�?EN}�H��=$���������#u=��d=-��>�>>,3�C���t����Ѿ��P�T<œ�>�>���>���>^��>��>?�x$?2(#?�xļDx?:0[=O >�ޭ>jG3?`?ta(?p�U>��=Bȫ�<�#�
�(�d�E�7��=�Fv��Z�<m��>��#>��ռM�=�\=����ͥ�l@�=��Q=S�<$�W=9��=���]c�=�i�>�X?�.���a��=B�P�6=�ͮ���>#,O>�J��.�>�U�>��S?p�L?��?~��<"Z3����F5��	>A ?��y?l�O>����yx(���ʾgNX�M�X>�i�>u��=o�Ծ�˾&��{?�o��>$�>�>��]>
�f?��>r�?r��=bO������,�,�=ݚ)�	;�>A��>��V=|"̾�a&�TBc��mM��^���)R��fO�V�=�2O�/}>�ҡ>eZ�=*-н����=!�> 4�=��=��<>xˀ>�}?eխ>�m��3͸�W�ܾ��@?y�z����=8>ae�^��>]0�>fF����ƾ�->:�r��'��N�Կ������>� �?�8�?�;�?�O�Sý�ex>�휽�s�=S�<{I���C���=�\\<�E>�AB�A�� d>�EZ>ed��(S��0��f
�����Ѳ�B�T�{��Jǩ��9ž/3�,�˾�½��
�?� >~Ϛ�A(�R�r��ҽ;ᱼ�	-�9tN����B�վ��?���?�4ʽ��0�Ys�{_T��{���R>�)R�����@��I��ّ��+P�о��	]��,0�����"�>bmf�F^��!�p���"�5_H�;�={�E?��5�T���M��(V>�YU=�_(=�kҾP�\ɠ��ƴ���\?�H?�^۾T���F�ܳ�>� ?#.�>���>�嘽澾��x>�w;?���>x{!�eᔿ(i��~B��8��?2@�?��6?-@s��T:�@|%�2����h>��?�Ju?��s f�L����*?��.?l�F� N5�?��+1�̯�>�-l?)����,>�,�>��'>N��:M-�X༩���!�?=67��\,�ћ�+\���>�J����T>�L�>7����̾��>+ݾ.���(þ�����=a�=��>����=�0�<0u����O�2Z��P$a��w���b?�G�?��&?�qU?����"�Y�½��>љ�>�+�>�!�=�`�'�>�f?K%a���qr��i�?��?Sk @fď?�DI�#��Z����=h��A���FM>�@L>t�>��� ����=ޑٽ����#�=�q�>Y�>z��>�I>��+>"�(>�}��)�}��������D��w۾���6yb��5���G��� ������_Ծi����ӽ,D^�k�(����[-2�Wپۧ�>�4?��<?|.2>}L�=CE>�!����e�OO����U���c_ ��m�4�T���,�01��l�D���½���4�2?��<g�=�ƽ>�H�ذ��`�>{�9>R}�=0d�=��0�c��=gD9='��=P�5>X�=jv=�،>	<�ٍ�1�����1�W�b�r?8���'��"�̾(]���=S��>�:?Կ�>��'�����v}�b�>�������t��H�=�<�>���>u�	�6�C>�/�����cF���>i�ۺQvϼ�𽼠��N�I���[>���>�Ҿ�p>Gt>��(?�Zm?�).?G!d=���>P��>� �>t�= �F>�(G> �>��?�b6?�c'?��>�]�=_i��G�=�<�y9�9ì���0_�c���Q=�ó��-=_T�=.M�@h<rv:=�g�*J�<d�<�(�>d�6?���>���>�@��Jn�7ۂ�=8-�mK�>x��<��>�� ?3~?ء3?m� ?F;�>��N�f����F��>�Ȝ>Hς�ǳw��)@���~=L�?�?&�Y?�*������\>��>6vC?R�?V|c?��?;�<=u�Ⱦ���.kӿx$�*�!������u����;��<���M�r�7��-������S�<��\>��>Mzp>M�D>E�>�?3>|R�>�?G>�Ǆ=%ޥ=%��;Y;��E���M=D���+G<��P�; ��xGƼ򭗽�(����I��>�F��ټa ?=��>&�I>/�>a�_���龅�B��rw>l�>S�N?��2?��:��ftB��RK�Buý� ?�fG?�-�>�2��5>ĺ->�.9>Z�>�Z�>�$��u���O�ƾ!�U]-����<w�?����D���vn��̓�L�KY�>��x=���m�?9Z?Fe�����s��P1L����>s��g�^�赾n�ճ6�T!v��g�Du�=-�>��?7�O�CW�=����v���x�#��G��=�j�=6��> \>'7	��ᴾbx�/�ƾv�>�{i�<�}�>�M��{k? ;I?�b"?T�?�l??�"�"F=?z�>M�7>+�>@��>��&?�%?o��>�t�>�v�Zv�q�F�ݎȾ�>���8�y>�}�>��>{�/>�K�=~>�(K��!>�$����K���������;�48=�MO>��>�\?�O�jM�=`��=���T=Ҟ=��>M�v> ��xAP��c>$RC?R?��9?�8�>����V����эZ>�C?�l? ��>�ē�Vr=�ھ�ݿ�F@<��=�iH��뇾����\�������>1�>V>��g>��_?�d:?��!??��;I}�$y�������Ľ����>�!\>m�!�������`�"uL��V"�Bq��)B��=6�=���=4�)>Z�=DHT�h���b��騽�T,�D��=�ž>cT�>�	?��r>3�a�R�Ⱦn��#�C?/D��}d�������%<�G�>J�<ɲ����'?�C���l��j���<S��ݛ>��?���?��?�G����F�>��ƽ��!�/y�=RvӾ�c=A��>�V�>37�>��=tm����=�b�>Õ���5��֟�(��u	���ʿ7�J��=S��"ھ�\��LH���b��Y=�;ؾ�8��*���K#�������༼�|�����ʴ���!��\�?��?}zo�-1;��勿�1C��
�@(�>��߾�h��d�x��¾��@�w$���� ��"���F5��&�Zl*�w�>�ݢ�4��:�p�Yr�I�<��>��?O�Ⱦ<��Vо_,#>�f�=G���A���B��Pژ�}#�LG?��?�����f��?�<TR?���>���>�p�>P���tOD�?��I?�K�>҃v=���HҊ�<�<�ت?�N�?sy9?�`��S!��N龞0�>H�+?���>e~�>�^>��]�v�Z�g�I?zE?Ɯ��{d�����E�4����>/g�?M���W>��y>|_>(e�V��������9(��m�=3���^����E��4 �;p�>PV{>	I>X �+�;���>�P��`ܾ?���^ξ�T�}n=��>�\̾��&>r��<��;!g3��J��_�R���;�W?�!�?U�2?�Z?�R�RR�;M����=�4y>�F�>�U�=
p4�R��>�?�;�u��j����/?
4�?I @-�?�UO�DGӿ������+��֟�=�%�=�>>K�޽dʭ=��K=�ޘ�YU=���>���>po>N;x>��T>��<>��.>^���v�#��ʤ�ْ�\B�� �����vg��{	�]y�����ȴ�����������ϓ�o�G���T>�T�ɾq��>Z�D?#Z�>��>�2�>�f>��
���to(�C� �f��-�Ѿ�޾]x����/���Խ��A�i�R��P���??���9?h�9�Ɠ(>�
�>��y=_�����f>��>+R�r>o�=!>V��>�m>���>9��>����@�>��k=�ے�ܡp�U�o�lᕾ3ԽXq?fȈ��׌���������R�|=Pt�>���>�o>��B�t݅��Cy�� ?�6��b��������˃�k��>,�?�>^��=^/ؽ�ľs��:->͇�>x�>d��/�#���S��D=!��>�b̾�>o�%>+�'?�t?��7?���=���>��z>[�Q>M@>�g>�d>�Ȏ>�*	?$�6?��(?��>x7~=� Y��mü��=��z�=����H �0�ʼDk�<ț=��`w=�}6=y<��e=Ur=�K�d�=oF=��>]d1?).�>oj>p�]���%�p�T�i~̽̃>�)�=�L�>1��>c�?�?���>��A>ɜ��0��!Ǿ-�>��<>+�z��3��*� ����>X/�>X�?�?�4�v����J=��>[�??�Q'?]Y^>��B��f������ݿ�2��=��#��»0*߼Em���>Ϗ=�*6��H�/��=�R%>p?>��k>1HD>��>�K�=d�?�O>c�0��(>��{��<��=�>�=���3�V=��z=4�%���$�����<��<l��'�����J�?�+C>89>t��=ӡ>���)��	����>���>7�1?pI?6�B��G��2��%[����R��>wqC?7�>��Z�1�>t0Y�^�r:�=z;�>���>!�e���\������C���>�A'?B��;a��/0�ZJ�����>A�T=d��D��?%\Y?r���[���d.��N=�B����=�����1��wо�P���6�-������>,a����=�>�%�?
�?�o�=����uw���‿(���\0 >y�=h��>��S>�n����o��t�þ����ڡ<���>���0?��[?�-�>�B�?	� ?�%?�ܾw=?
�>�%p�"�>E��>�=?I?S�>!�3>eV��C���c��Y�۾�7;�1����=�F�=
�>!�;(E�=�^h>	����ǽ���Sfӽ6T���<���=��J>��>>��p?����DZ>o�w���5�g�9���B>D��Gi��+��>� ?�҂?wa?F�?�,�Y�g��=U�<�=��Tq>Ř;?w�^?�k�><�Ľ,X'=&(���V�������>�k==�B>�Ԃ־�f>��x7��k>2G�>�:<=9�n>D6n?ޒ3?��!?`����+�"F��֎�� =jj���>͵�>�������̉7���c��N�������<2��� I==>>�P>���=z�=���=�4�!�z�u�����<�:���4A>�)�>p��>͉�>�.%>P�ž0� ��D?`�ž��J����=���᤽J�>�=�`ʽ��"?yِ�QΣ��p��\K�Ǣ�>���?T�?���?GLV��dҽ��=���`�<��{k<2+о�yG��� ?�'�=�
U>���=�i����=�2�>�sJ��G�Í��7�w��#�ǿ��<�BT��񫇾3�k1��%�X�齇:����7��G�m�ƾ4��]S�n-9<5�7���;�����澜��?�գ?�� �-��=H]N��3�l�����=����T�����5�M���X|������J.����)�s� ����H+�>n��"!��+ȍ���?�GE�=WԀ>��/?akӾ����پF_���	i>�Ų�XC۾k.���ǜ��0转2>?l�?�v��kC��2�ɺ�>@��>�Ʀ>yj>�ؾ�u����>��?��>v�s������:��O�ݽH�?�)�?��>?xc�oV(�q^��ad� ?7W?KYG?.��b�6�X�H>t/?�?���?�3^��ޯ¾K�?���?C�����e>�n�>�B�>%�I>TZ��Zޫ���P�q�R>�w>���=ߓd=���\dm=�$�=Y�>Cj�=�,��5�U��<�>�:�'2���5�����N���;y	?:����L>�o�>{��= ��w[���r�����t�K?Cگ?�jC?%�4?N"��i���BO�'@=�a�>�&>\�<��u��>˸�>%����e�d��ȿ?���?U�?�xX?%�����ܿ ��7���JW��я�=7��=u��>Ł��y�Y�>B d<�Y��c�=�v�>�1�>�ˆ>c�T>�@>j�B>|�����,�ϒ���	��\�A��.�ߔ����+���#�=����)�*��
�G ��q�H}�Y�뽞4v=&:�z�[>z&8?8?�Ι>�V�<�"�>H�}�C���������&���\I+���ؾ�M��b,�>?b��B��.-��H ��"?�W��p�>t�	?(;��>U��>N�?>�K���]
>���>.q\>v���>zц><��>>���JZ�>ʉ�>nI����_�PPW�������!)m?@��<K!=��0��𰾢���|>�WY?�
>{������_X�Gd	?-�Ͻh�ؾ�����x����>��?x�>����󳾀=�ʃ=�R�m���d><-�����<��=�� >�~�>=G��R��>��>�X1?'V?�f?�h���D�>�O�>���=�8k��˂>4�>�0�>�)?-�h?OA?��>�������L�=4x�<)t������j<T�O<�<��N@=�є=��S��Z$=��<�}#���y��#���E=�5=;�>�b8??]�e?��?�;e�=����}���<e��=<?�Q>Q�?��]?�??}8? j`>((��pO���>zl]>"�|��k��/�>|��>|�H>�?�>�,ؽ�N���[�=�l=!�f>���>rm�>a�>����tż�W��t���Y�)\���>�K����>�^��>^�#?�_����?��j�<o�>��<<���>��>Q�">a�3>O��>�~>8��;7Y���T�j ���gs����<잘=Q��JI$��m>͚>>)�=�����{=c �=SL�K
�UL
?�K$?r,ؽV�O����r4}������G>�?�\�>���>T��>���,y�h�N�d"���:�>��B?2?���V�{=�#	�vb���V�>ז�>xlq><�>���g���� ��'�>�??�?>zh9��F�YOV�b�̾ET?��=Ʃ;�|�?Ɠ?�������N�OU4�z嬾 ��>H�>�������e����^��{���{����=��Q����>Hu�?g���C��>�����裿@���0�U<�=Rg���F�>�>��;�C�Br��<vP������`�X�<�U�;�9�=F�S?r?_lf?�� ?��?�X�����>��>6��=�w>��?K+?��?�z?e�<?C��>��Z��M�p���x��=s�W<�f�<Α�>�6�>@i>A�X=�W!=]�/>�N;�'���%��=��=yU�.�q>�><i�>=?��&�r�;�s%��MN=��1<�B\�^��>�Օ�C�����=.�� S�>��?s�>��=K�Ͼ��о�w��X�=KC'?��>��>B���(��>$�/y�����>�=�O��1V=�q��y�	����>��c>�G�=��>��h?��?���>A���b��HY��,�
(���%ܽ��?a��>��c���2�I�n/��Rl;�	���q=�Kb�G>�R>�!<��>�ص�z��=���+���Lv���� �0���4>ϰ=Ze�>�j>���F��W�˾R�D?㚾-�	�S���Һ�0���9�=��>�﮽=�	?���|��Q��K�2����>6��?Y��?Oyf? kZ�B��I�F>�`>�*>Kt���~P��o���m�Ҙ7>V�=�^��u��֊s<�dT>^P7>�����ľA�+VA��W����3��7t�2ݻ���L�8��>�ž`?����оW	=�5�y����>oFK�!�j�0��=����Z��r)���{�?�v�?���9 �㼝ZԾG��P���PT<̗�,�@���x���P���Ѿ��e=Cž��{���P�R��o��>84�_捿�����A�O�>��7>0{-?ט���?��e���`�*>��*>A�������ޤ��7����;���O?˚4?ϒ�&\���><�t�=]X?�L�>�p�>�Xھ�d]���u>��?N��>}�	��
b�w]��-rV���?�#�?EQ?���<�S��P��H�B�J?R�?p%B?�T�w��3��=�2_?���>��Ӿ�B��헿f��I?ۧ�?�=M��|>��?��?3x7�w 辗�߽�1̾�^F<`�;>��>�⎽�-s�b�>=y�=��;>���>s���Ծ	��>����N��]G��C���#�<>�?�J��l>�Nk>�y>��(�����2���b��:�L?n�?�4S?p8?�6���r����[ۈ=�|�>2��>硩=�7�\��>���>��L�q��T��?Z/�?'x�?��X?_�m���ؿج����4"�����= m�=5�v>X���y)=�5=^� �㢪<J>���>83}>��>��]>�nE>S*>����+(�p������b�;�%���-��E��$��6���������q��B5ٽ�a����/�j2��(�aB��vKz�F1�F��>U\?�ת<�>]�_>�è����TK��XE'���;��{T�bȾΠ^�5۽��ֽ�	���؜������:?����#A>K�?��K>�L�;�cd=�@4><�l��J�>�n>ŭ�>�@A>�;>Mqc=���>>r�<@)��Y�>E����ri���;�4&��Q׾�bp?��>)�����������0�Ի�=�c?�F>=�k�&nԿ���$}?����nž�����������>�E+?�m�>|�o����q���=h��n>��>�	�<�9x������,>,�<�5S�1�?�:�>�(I?�i�?�A\?��_>�����Ċ�o�>�Ž�}�>�o?���>�)?qk?i\?x�3>���࿂����	5=f��3F�D�绩G�Lq��h�<��X���n<`�=�x>fo�<wYn����𢽦$.�>fI?S�?�?�8>e[:�L���� >;�=�G<� _G?��>jQ�>�8?a�?0%?�t�>�
n�(@ ��=�>�j�>�}���}����=�M�=��*��?^r!?9	T��|��!�=lH�>�j�>�*5?�=?�x�> ����R���$�ٿ���'������  ����<�"����Gbz�Q3����<^%�=%�B>"��>���>�<N>�!>Zc!>���>Mo_>���<��=��N=,w��n�����= ��~�-�fZ��4~��X��&��?���2��0)��I�\w���R?5�?T|��>����㽧oо�*��W>���>+��>Nq�>���<Pξf�3��qj�#S����P>F,?�#�>�w���z���=��V�m{�<�[�>΍�>�,)>=H\�B���쨽���>��$>D�>4,F���M���T�)I���M�>eq�=���K֝?Ɗ�?�������������^�@�6>e��=�4Ѿ	L��a���*��(t���o�֢����ӝ>��?^���9���3ž/���]��[o���E>U��=my?_>k=��&��,�&�!����z�ϻ<�>�>|�;�uX�>��#?1�?�v�?��?�-�>�hg=��?v1�� �>LM>�A�>��?�.%?��?��?��U>�}��R�y�F����K�<\8��8�|F�>���>sl�<��z=�ɿ<egJ=0�r<��;�';��o�	����=��y>H�k>���>0�?�׽��<J����C�������{�=�o�<��=g����O$�R�>���>�?���>�>z�̾4���3��+��<�G?�L?�jC?GL�=����E-
�l���S>��>gr�NuǾ,<��K�ð�f?亪> GT>(z>:-r?��?4��>��3����ܸ)�?�A�~z�=�.z>.�>��>fϽ8���@�N�`<V�m�M�?�����=d�����=�u'>4��=�Q>!���3�>P.>r���n�;��=�������>���>V��>�o>L%>fT��b᷾k�H?6|��R<�i(��)fپZ�p���>�E>���n"�>]G򽽿���z��=6����>3J�?ki�?Ma?��C����߮9>��c>"�>�c��|�+�bd��á��3Q$>�9�=��������L<�+m>�ӈ>6��ž�e�A���T��T��J��A��`��z����P;D���9��js��v'��G�*x4>f�I�-�ɽh���2�^���U�޾魱?UӬ?D�˾HW��t�����8�t�G�͵�Z��<�;==�
�$����ֽ�c��8����\E��sX�Kf3����>��ۼ���ݱ��%2�S:>���=���>8~۾��Ƽ8���|W<��E>���)I�,
�����)x&�'�?��1?���+�	�ʆo�a)�=�%?+��>(\�>�b޾�X���;
���9?�=?����o�����i~ܽb�?T%�?��B?��>�}5�ό/�}��6�>�?}�?r���=�~{�g�q?u�,>Mn��1oྫ��3�!��>%�f?��D�r��=�B�>�\�>O#ս.���4'������S>⏆>w�W>=������7�=�>ih�>��>@Rf��k����>V%��N�ϦH����,��И�<Gt?�h�>c	i>�o>�(�Z��vΉ�eR���L?{��?��S?�Z8?QH���E��-ː=�̦>���>%�=�����>��>�Y�lur�k�˗?�E�?���?�NZ?i�m��n�'��� �Wؾ�f.=�A�=�+b>��D�>�`�=I" �;�K�^.>MF�>J�=i�>$�h>vjI>D�9>�ɉ�l�+��0�������.1�i��f��8Q����1bl��$�KϾu�P��*��b���Iۼ����y�M�,)��0̫�6D�=[�+?#�?�߸=����9Y=>W�ĽJ�R�^�M>�˽C�>�IL��� �������$'����# ��^|��5�\�0��h?/E!�R�=��,?tV�=Q�2>9��>gOm��^���u>NY�>`F�>��>��>��$=#E�>a93=N�#>�\�>]d��hXP�0g>���پ7t�_�G?J$=�@*�+��Wn��-i�F =��
?���=��Q�T��Vl��?��ۼ��о<ΐ���G����>�?��>XZ=�:�������<%>��>ai$>��5>T��{����V>�%>Wo�_[�>�O>h!/?��t?��D?������>֝�>��=و
�L��>U��>��>n�:?y��?��K?T^>���;�����Z����#����k;�Q=DHμ�)�8�$>0y1�t$�n�U>�G>���8֮<n׃���[��$>:-�>TNQ?�L4?Y$??�(?x�~�M����
�b��>�&��4�?��>�?��?��0?�2?4�o>.Eݾ��V��>2��>z3=��Hy�
�>`�k>�j����>wG?Ğ$;M��+�J���>���>���>�0?��?a>.ƽ����}���A�����L������=:��v����=p�Y���|��ދ>�H>{3�=,�>|�
=����>���>�A>�_>�:�>}ҽ��E���9=*ː=w�ܼ���;�AH=x>�Jo���3��>�.W��
��/(u��D[=�=?<F'?���\TI�®Ǿ�UԼ��%��.�?!(?��>qΊ>vSF����G<�4о#�?=�+?�r
?��B=�R����1����L=zA�>���>-�>-�Ӿ�򾙼.���,>��>&��>�P��x�`�3�]��"Y�>A�
>�۽�ڛ?�?�YоFMžg���k2�3�M���?>Es8=�S�6�L��վ(ﾂ����2̾�U��x���J�>���?jG����=�`�?��ې��y��(ƴ>�&� $�>�>�Jؾk���l/�{6��}հ���˽�����D<��7>�;?r�?��?�?03�>��k���>Z�ͻ1�?7�=�K�>�
?n�&?��?�-?�r�>Gӫ����(M���x6�]�B�XJ�=?�g>;�{>�U���o�=T~Y=�ݼt#�a���A��<�G�^[��lM>�8�=| �>Mv?�1?K�I>7��>���>�G龢���&�z=7ٷ<��=D&�=�[�b�W>~1?/�O?5�?��>9��g� � 7�5�S<m�
?foZ?c��>���v�=Q����B��J�=��>Sq��^:�	(���*0>�Z�>�<�>�����Z�>8�k?'� ?0l�>a�?��|��
^�_&c�% F>.F>���>V�>;��%q��F��o`���S�E��)�W=W9����=�l�>/�7>��==��=�lZ>�R���_��o�=6��=����>T>V>B��>���=ֵ�=�7�l.ܾ	6?Ӕ�_p�Cp���������/>e>	�:����>�����oi��_���~&� ��>5��?��?�Vz?��3�>x*��\�=��r>��>�C ���
�>�Z�<�0�=W�.>]]���G�oƼ<LeA>[��=eE����ů��ӽ�����6<��b��j!��a��Cy�����oft=:�_���̾5>侱埾�^���5�t3�;(R��ǣ�yS��d{��©?	^�?a�4��J໼���j1�b�.��s�=uJ󽆌߾����a�=2I|�_������p���9-�<VK�ޗG���>�;�<;������� �L��F>�Y�>��3?�8�I��$h���j>K�3�,�	�:��.o�����!tT�$�&?n=?����Q����r�����>; ?z�>��2>�Z���QQ�v��=d�6?��>�������f��ߠ>��?M�?��<?�=D�5��;��v��(�
?7�?	�?n}��aK�"gz���P?頑=OMT<@�>��X����"�?c�>�0�?�\�Z�^>��?\|�>�[<�u��:^~�a�վ���=P��>A2�>��[Z���D�0ݞ>�^�>/ O>U�%��6�WR�>����O��pH�p
�Ѷ߽N��<A�?�G��y�=b�g>��C>�O$�C���넌��a8�1�C?Ѳ�?�ob?�8?+����⾯�ཇ��=���>X��>߁>��C��}�>!��>p�Ͼ��g�����:?N��?��?��J?�n��ؿz����ϧ��@��Z/�=Y�=��v>�< ��Ƨ=�u=��E=l<3��=�X�>�9b>�{>�l>TLc>`\9>�y����'����vz��mI����y�aW��<��[���1�%_���{����!�ཥ���	1r�X�k��G+��R�V�3>�t?���>�={5���?o_o�I�0��ܰ=�	=���G�Im��Wn|��Hi��;��C��򵽐Η�w�!�mr�V�	?Fƿ�D~�=�)?@�;��>�G�>�lP��G6>^�(>��?>��k>��C>+I�>&��='�=
�>-��=K�>��QL�xh�*1����	�U<2?y�D>rf�y���I+���ľ)^?��	?��> 
Q�Oz���錿D|(?v���~Ѿ�����N��`�$?�V?�v�>@���
�F��;�=���="���L�>��>�o+=󽧾q;f=��>��>������>ݻ�>O�?�RC?{�9?�A+=U>�3�>b�>���ߜ>w��>�>dk%?=�T?��0?�>�<(ko�D#!>҂K=@�X��E���g�5mF��ֽP�Ѽ���~J���>��>�y��
Nͽ�#~>�<�<}��<��>�VL?�Q?�?�$o:��X��b���宾�g�>:�=��?�?�?��`>�Zw>�>MJ�='q��ǾǑ�>k[->�"b���J�B>>�͕>!6�>�!3?�d%?�������ᬽ��=>���>t&?�+?� �>M�R�����F	�)�ʿ�!��H!�iWi�M�f����\]��&�j#/<�1O����s�=#�X>g��>�4r>�2>��>�c>��>�LV>��=fp�=��<�����n���=Ūd���=��9��ن�����Ӽ�%�<p��s��j��Ud��b�?��?6�P��௽/cB�kL������RH>�?��?E��>��>᭾��f�>�\�*蜾��>��1?=?������Hf)��+��8y>�(�>+ި>fYn>�'��)��y�͠o>_Q?9s>���<��0��j��9���{��>xUH<w��X$�?�)?����оUg���O�/ F�9��˞>In��}���=�ﾬJ@���������I�u�|�9&�>xk�?�����:%>�x�\J��::��}�����>�)=z?��>�$��n������Ɏ�0�����gXJ>������>&�P?�cX?p�?���>�<�>����>S.�=��?\�?��>�zP>��S?d�@?�0Q?�_<1K��-�	�Z�]�ʽ�����q�=�fE>�54>��8Q*>T�=�k�*�W;<���ƽ���:��h>���>�>�GF>�?��+?=��=�<��������O>@*�=�����B�>f�ǽt�'��i�>?�?M�)?���>XM>U9��s����Ҳ<=��6?�1T?z	>��{�WF>!���?ʾ�gh>�);>�� �B!`��,��=#P���T��۽=��>"�3�5�L>�2|?A+?�?�'^�i�3�[���QF�4�J=*~1>�*�>m��>|��=&����*H���J�}I�<k�����q.���=�0=߇�=��G>W��=�>Z��=FI�=��8�=�p9=�Ž>ҟ�>ơ�>�`>u�f>�߭������I?������O���N�оX ���>3�=>��-�?ą	�[�}��ܥ�G�<�Z��>@�?_�?!�c?B�B�L���[>tbW>Q>j�<l�@�����@��d/>���=#Lv�����ʋ�;�D]>��}>�fʽ��˾�_�CF��&�25�����B����<�<&�64�l[Z��=�1_���������ې�]�Y�?Y������~�����|F�?J��?̛�I󏼆(�w~�C6������3D����ٯ��F��}:�ջǽ�-l��޾%R��R�*P5��>�>�s������|�ޠ,�2�>f^�>'??���=� ��<����l>�ž{���Ӕ�ʩ��e᜿+WT>��e?�Y?��Ծ�$��a�?�޳�>�\�>٧>�+J>f���(��>:w>*�N?]��>�[4��Lu�ZI���7=P�?�6�?�KG?Vi�W^@�@/C����h\?��>�\K?�ӈ�AH��5����>��R>	f�=P��ׅ�Q� ���?1�k?�b�סּ>Y��>$��>y6�5���^"�U���8��<��>�o[<nV�����;�1���.T=���>g�8>ν��f龝<�>�:�'2���5�����N���;y	?:����L>�o�>{��= ��w[���r�����t�K?Cگ?�jC?%�4?N"��i���BO�'@=�a�>�&>\�<��u��>˸�>%����e�d��ȿ?���?U�?�xX?%�����ܿ ��7���JW��я�=7��=u��>Ł��y�Y�>B d<�Y��c�=�v�>�1�>�ˆ>c�T>�@>j�B>|�����,�ϒ���	��\�A��.�ߔ����+���#�=����)�*��
�G ��q�H}�Y�뽞4v=&:�z�[>z&8?8?�Ι>�V�<�"�>H�}�C���������&���\I+���ؾ�M��b,�>?b��B��.-��H ��"?�W��p�>t�	?(;��>U��>N�?>�K���]
>���>.q\>v���>zц><��>>���JZ�>ʉ�>nI����_�PPW�������!)m?@��<K!=��0��𰾢���|>�WY?�
>{������_X�Gd	?-�Ͻh�ؾ�����x����>��?x�>����󳾀=�ʃ=�R�m���d><-�����<��=�� >�~�>=G��R��>��>�X1?'V?�f?�h���D�>�O�>���=�8k��˂>4�>�0�>�)?-�h?OA?��>�������L�=4x�<)t������j<T�O<�<��N@=�є=��S��Z$=��<�}#���y��#���E=�5=;�>�b8??]�e?��?�;e�=����}���<e��=<?�Q>Q�?��]?�??}8? j`>((��pO���>zl]>"�|��k��/�>|��>|�H>�?�>�,ؽ�N���[�=�l=!�f>���>rm�>a�>����tż�W��t���Y�)\���>�K����>�^��>^�#?�_����?��j�<o�>��<<���>��>Q�">a�3>O��>�~>8��;7Y���T�j ���gs����<잘=Q��JI$��m>͚>>)�=�����{=c �=SL�K
�UL
?�K$?r,ؽV�O����r4}������G>�?�\�>���>T��>���,y�h�N�d"���:�>��B?2?���V�{=�#	�vb���V�>ז�>xlq><�>���g���� ��'�>�??�?>zh9��F�YOV�b�̾ET?��=Ʃ;�|�?Ɠ?�������N�OU4�z嬾 ��>H�>�������e����^��{���{����=��Q����>Hu�?g���C��>�����裿@���0�U<�=Rg���F�>�>��;�C�Br��<vP������`�X�<�U�;�9�=F�S?r?_lf?�� ?��?�X�����>��>6��=�w>��?K+?��?�z?e�<?C��>��Z��M�p���x��=s�W<�f�<Α�>�6�>@i>A�X=�W!=]�/>�N;�'���%��=��=yU�.�q>�><i�>=?��&�r�;�s%��MN=��1<�B\�^��>�Օ�C�����=.�� S�>��?s�>��=K�Ͼ��о�w��X�=KC'?��>��>B���(��>$�/y�����>�=�O��1V=�q��y�	����>��c>�G�=��>��h?��?���>A���b��HY��,�
(���%ܽ��?a��>��c���2�I�n/��Rl;�	���q=�Kb�G>�R>�!<��>�ص�z��=���+���Lv���� �0���4>ϰ=Ze�>�j>���F��W�˾R�D?㚾-�	�S���Һ�0���9�=��>�﮽=�	?���|��Q��K�2����>6��?Y��?Oyf? kZ�B��I�F>�`>�*>Kt���~P��o���m�Ҙ7>V�=�^��u��֊s<�dT>^P7>�����ľA�+VA��W����3��7t�2ݻ���L�8��>�ž`?����оW	=�5�y����>oFK�!�j�0��=����Z��r)���{�?�v�?���9 �㼝ZԾG��P���PT<̗�,�@���x���P���Ѿ��e=Cž��{���P�R��o��>84�_捿�����A�O�>��7>0{-?ט���?��e���`�*>��*>A�������ޤ��7����;���O?˚4?ϒ�&\���><�t�=]X?�L�>�p�>�Xھ�d]���u>��?N��>}�	��
b�w]��-rV���?�#�?EQ?���<�S��P��H�B�J?R�?p%B?�T�w��3��=�2_?���>��Ӿ�B��헿f��I?ۧ�?�=M��|>��?��?3x7�w 辗�߽�1̾�^F<`�;>��>�⎽�-s�b�>=y�=��;>���>s���Ծ4�>$ѱ���q�g���i�8��(�>�!�vF
?H��z�=����0?
�E�YĈ������r�<��*?���?�_q?�f$?�ϼ�u&���j#��e�=�ޘ>�.>r�>j������>��?t9��x�
� �Z��>u��?2��?� �?�䌿"ۿ8���U��������!>Vy��_-=���.>�^;�#���]����3>���>λ�>5�u>�#->�>�S�=�:���0�)���Я����8�k�?���5�/_��&%��[� �Ø�����������g^�Í��@�e H�vI0<�+�!���C? -�>��>��>>k��M2������)-��+����Ⱦ���D�=+ľ�尾�k����e�q	�nS���?z_���u�>�\?o=ۡ<x06>�<EP>L�>�A���}�=�RB>(��>�y�>�(>5�4�y;�>舘=u�����y�8�8��9_��\D=�SC?��c��b��+(5��H��^����>��?� d>��$��앿�>}�rK�>��0�_�z����̼�~�>``�>}&�=�m]�%2���R����z�u=��>��=ʝ����|������=�7�>���峗�[��;zk?H3?2.?�z>Px�>ͱC>��>Tk{>S*�n����=��'?3�G?~b1?k��>��=G��D1>@���D�uƱ���8�r�f�?=h�T���=5�)<h� H;+㬻!ۗ=��`=ݮ8���\�>�2?�??s?��l�;�:�Ӿ�ф�/m:>���@j><������?A,�>~� ?GR�>�Y�T8!�".����>I�>�]�t��*��k��n$?�b?�@�>B��8�� g;�h��>₪>��$?�"�><�j�!���=����������ɾ@Y��2Z�����������=��X�Htǽdf�=�;�>J�S>�o>��z>8�#>Ө=9��=i��>��d>�8=�3�=js���5c>=�=5�˽֋��|�W��}�WW=ϋ�ɕv��,��ׂ�	9&���>���f��>��>�3�� ��-��y=��lC��5"?�?68�>L�4?���>��C����P�[nP>�X&?�C?RH>�ņ�����ll�����>&J༉ne>�>a"0��@ν�V��=�}^�a?�G�>���<#\��WK�&��K��>�}&>���ri�?2ف?2�iF��%����	Ml���>ʵ��u��+x����(�|�x�>�����\ޥ�2���[�>\�?�ࡾ- >��d��ժ����🾶;?�G�>-��>T^�=�NP����;�о���Km%���=�|�>��>��>d;�>���>�^r?�Z ?L��>��%��+�>�t����>!>o�>��?�?���>2�&>:�_�8���%��q������<Б�=ed�9��}>��=I=��>5�#��>�;x[н{PK=��������"�<�!8>���=^�=��?��9?��d���G>`�'>{���F�>�=i���@{�1�>ħ���x�>�V?�N@?�
�>�Nj=)�"%��T޾_.�7��>�G?%�&?M8>C4ݾڽ�6G��1�;�*>3=�_�Ӽc���W�@%s��u=���>�> X�>L?G?o�x?J�v?�PP��ZZ�W� ���m�h�q>E�s>~a���0��j�>d���pH���>J��c����X���t����N<)�CӐ>���=��>�
w>2���7?>Z2���`��8'���M��m�p>۬�>Ȇ?�}>ܡ9�6������؞1?��s(�;�������[=ʽ�~�>^k'���>�b?��������z�P��<�=��?@��?��?�S�Y�`�1�_>��>� %>)����)ɾ�d�'t><P�j>��=p������_=���>tf>�ܽ`}��^���C轌�̿�Bo�@?�4�����x�Ϣ����߾Pe�x���2����侪Z���Ju��Lҹ3�Ӎ�_����r�����? j�?���=�׾�}�ZW���<ʾs�>𙾾}�4��о��q�x��q��'��T4�%U�|�'�n����sR=�D�׈��臃��ɾ�z0>��=�t�>��Ⱦ���� �!���#>db�>#���;�&���p����~�?7�?G�y?�L)�$�V��$��a�=\?�|�>�M6>{ga�"��<tm>��W?��0?�]C�����e�E����d�?���?%,5?��z�.Up�-�ܾUb�=�,U?�.?�^�>��]��k�<f�c�J�=�� ?*R?����ه���C��?�s?�i�D�>$��>V^8>H@�����6�>-�`�g璻 �>T$�s��;�dn��f��ų���>���>�^��ď��	<�D��<x��SX�̳��Fc�Oj�=&a?�+7��;�>9Ю=&u�>?K�~
���u�����B8?{@�?H�?*;K?"�оC���6=���>Y��>`��>�<>GⒾ��i>���>�߽jB����-g�>72�?��?��x?v�x���޿Ӭ���Q~�q/��<��=�PB=U��=����=����Y���䘽��&>���>���=*.>.��=�+�=>Z���Z�%��p��1c��V�D���@��L��Cd��Q ��|u��B%�I�ܾ�#�'ϐ������P�	����N�J�=�Z��Gj)>��?��>\�>��f=���=<��,I��l��J8Y�b��8E������gȃ���k�8w����G�툼�����?�� ��c=fr
?����\���y>@J_��N	=E��>A�F>H?�>�1>P�_>��&>��=)�>�>�>tvh������D��� YY���[?�l2��]e�0O����c��&/�>��?pr�>�V�*Q`�Q�E��>`m������Vn���˼uBs>�}�>��<���Ś>�Sg�_�������uo�>̠�>�I>�T4�U����G�=`��>�'4�'��������2?^�}?P)/?$!~>9;���td>�@?���>F���E=�<���>,$?�
D?h�?�k>�=2=���� >�j˽?4'����=uС��>Q`
>mW��zBU>Q?�=n>�3��ה���������<<h;�=r��>M:J?�w�>�Dp>W?H�D/�K8F��C���>RL&��Ԫ=��>?�>4�?��>E�*>x
������������>��J>i�J���T����<m|`>�\�=�?�M.?�ս�r��񀜽��=�U�>$�?��3?��>��=w獾���jӿ7$� �!�t���k�Y�;v�<��N�r`�8Q�-�D\��>�<U;\>���>ٝp>�6E>��>�I3>L�>�=G>	�=3̥=�;�;��E��M=�>E<NQ��ޱ�,�Ƽ����^ы�Z=I�2U>������ؼ��?�{?o8c���Ƚ,�5�X�Ͼ�������>%��>l�>�<�>d�=G��ux^��;��z��?G�c?^	�>�N�c<>��=��]=\q4>��d>���=��؎�Yg�n�E��`�>7� ?��>�,�F`��{�������>���=MĽd��?ˤ�?#P�j��a��,����?���>���<>v<G/>��y�4��-7���/���{E>��>�ޠ?�+<�'N>�wJ��g��}Dx�p	޾���=�_�*%�>C+�>�q�3%���� F=���0����,��>�z>8�>�%�>���>�5?�0?j�?���誵>�n�<�S�>��d>�O�>��>��?�ӓ>��i>�I�=��y������H��=�z�<�">XW.>Trx>�{>�a�=���<[�.>��g=���<�����<TҼe��=��=�P>�_
?f�@?V���#���7,>kLٽ�`>\D>�܀>�.�IK��㴾��}��:�>�7,?��?aM>l�߽c|��r��^������>�ML?1T>�$���Y>e��c������$�h>1��w�$�����#����Ž��/>�!�>�x<Ȏ#>��v?���?�~?�A;����vZ�S7l��W�>k꥽�Â=g��>x�0?:h
�?�M��������ي��7�����El��ڟ=paz��V?�ݧ���=0N�>'14=�3a�����{ �a%a>?w��>��}>q�>;(���*��y+?�~��> ��X�c5'� �z�Z�=�@�>��N���>���+�R����u�����>��?�4�?d�J?�4F���ѽ�5>��B>��=J�u�ٽ(yV<�n�=�Eg>.ww������p� b>S/�>%⣽53���[�E
oſg�M�	�"������8E�cd��AJ��8�<F���u�"=��M�:��m��3X���R���F���f�Իf������sd?o�x?]l�=�Qh�r�B��(�����t�>)O;������?޾�����T�����������iiE�]4�
t�������*X���l{�y�+����ߒ���$?߾fv���j+��|s<� >�]2�/� ��f���v��:r�S��?~vg?)Mo���N�/5��%��=�	?���>��u>�I��E�k=�>��D?�{�>����p'��R����=�W�?X��??-??�V��;A��;�C9	�u�??p'�>����0ɾ��ý`
?w3?ݖ�>������&����>��X?��P�o�l>�(�>�<�>[����0��I�3�����>����?>�
������g_�С:�
D�=3�>ju>2i`�N��4�>$ѱ���q�g���i�8��(�>�!�vF
?H��z�=����0?
�E�YĈ������r�<��*?���?�_q?�f$?�ϼ�u&���j#��e�=�ޘ>�.>r�>j������>��?t9��x�
� �Z��>u��?2��?� �?�䌿"ۿ8���U��������!>Vy��_-=���.>�^;�#���]����3>���>λ�>5�u>�#->�>�S�=�:���0�)���Я����8�k�?���5�/_��&%��[� �Ø�����������g^�Í��@�e H�vI0<�+�!���C? -�>��>��>>k��M2������)-��+����Ⱦ���D�=+ľ�尾�k����e�q	�nS���?z_���u�>�\?o=ۡ<x06>�<EP>L�>�A���}�=�RB>(��>�y�>�(>5�4�y;�>舘=u�����y�8�8��9_��\D=�SC?��c��b��+(5��H��^����>��?� d>��$��앿�>}�rK�>��0�_�z����̼�~�>``�>}&�=�m]�%2���R����z�u=��>��=ʝ����|������=�7�>���峗�[��;zk?H3?2.?�z>Px�>ͱC>��>Tk{>S*�n����=��'?3�G?~b1?k��>��=G��D1>@���D�uƱ���8�r�f�?=h�T���=5�)<h� H;+㬻!ۗ=��`=ݮ8���\�>�2?�??s?��l�;�:�Ӿ�ф�/m:>���@j><������?A,�>~� ?GR�>�Y�T8!�".����>I�>�]�t��*��k��n$?�b?�@�>B��8�� g;�h��>₪>��$?�"�><�j�!���=����������ɾ@Y��2Z�����������=��X�Htǽdf�=�;�>J�S>�o>��z>8�#>Ө=9��=i��>��d>�8=�3�=js���5c>=�=5�˽֋��|�W��}�WW=ϋ�ɕv��,��ׂ�	9&���>���f��>��>�3�� ��-��y=��lC��5"?�?68�>L�4?���>��C����P�[nP>�X&?�C?RH>�ņ�����ll�����>&J༉ne>�>a"0��@ν�V��=�}^�a?�G�>���<#\��WK�&��K��>�}&>���ri�?2ف?2�iF��%����	Ml���>ʵ��u��+x����(�|�x�>�����\ޥ�2���[�>\�?�ࡾ- >��d��ժ����🾶;?�G�>-��>T^�=�NP����;�о���Km%���=�|�>��>��>d;�>���>�^r?�Z ?L��>��%��+�>�t����>!>o�>��?�?���>2�&>:�_�8���%��q������<Б�=ed�9��}>��=I=��>5�#��>�;x[н{PK=��������"�<�!8>���=^�=��?��9?��d���G>`�'>{���F�>�=i���@{�1�>ħ���x�>�V?�N@?�
�>�Nj=)�"%��T޾_.�7��>�G?%�&?M8>C4ݾڽ�6G��1�;�*>3=�_�Ӽc���W�@%s��u=���>�> X�>L?G?o�x?J�v?�PP��ZZ�W� ���m�h�q>E�s>~a���0��j�>d���pH���>J��c����X���t����N<)�CӐ>���=��>�
w>2���7?>Z2���`��8'���M��m�p>۬�>Ȇ?�}>ܡ9�6������؞1?��s(�;�������[=ʽ�~�>^k'���>�b?��������z�P��<�=��?@��?��?�S�Y�`�1�_>��>� %>)����)ɾ�d�'t><P�j>��=p������_=���>tf>�ܽ`}��^���C轌�̿�Bo�@?�4�����x�Ϣ����߾Pe�x���2����侪Z���Ju��Lҹ3�Ӎ�_����r�����? j�?���=�׾�}�ZW���<ʾs�>𙾾}�4��о��q�x��q��'��T4�%U�|�'�n����sR=�D�׈��臃��ɾ�z0>��=�t�>��Ⱦ���� �!���#>db�>#���;�&���p����~�?7�?G�y?�L)�$�V��$��a�=\?�|�>�M6>{ga�"��<tm>��W?��0?�]C�����e�E����d�?���?%,5?��z�.Up�-�ܾUb�=�,U?�.?�^�>��]��k�<f�c�J�=�� ?*R?����ه���C��?�s?�i�D�>$��>V^8>H@�����6�>-�`�g璻 �>T$�s��;�dn��f��ų���>���>�^��ď��dk>�vϾ�QW�G$v�P8��[�=[V���?�Z۾�>c��<�@;>�%E�X����m����a��u]?���?�&?.5{?]V�&bF�:鍾�?j� ?:�>de�;8]Z�a�>7��>�.��/�W�T% �r?�?BN�?=Aj?͉���п����q���af����=�;�=~�Z>�������=&�*��-[=NF�=��!>��>m`>Amb>�8>q�>�Y,>�{��i�)������ؒ�dD�q�V��������۲��>���s�72�������ߴ����u�Z��4�L����N8���>��?@EF>�:\>UJX>�	����<|��Ҟ�"��ҽ���C�8D���u���X��f��4"�P���e���
�x�?�:��w�L=o>>���=�k>o½=4�P=�4i=�>�>�ɉ>����(�<�>��&>'8���L�>��3>��m��}��Dݾ�͚�K�Ͻ�/?Y!��N�5�?�~���ξUp�>��?Eظ>S��g|��[Y�`۪>��W=��?�A@���{�d�N>�Ԯ>��c=���=�)=�Xg��/����<bm�>�4�>�N�=�V��7����\�=.7 ?����"�?�z��=L;?�L?��?Ɓ�=	�B>4��>ڋ�<?软5L�e�i>��>�3)?��I?��?C5�>G >0痾�x���>[d�9���~����$�u��;����\�=�w���A�5}<C��==+�ؼΰ��pd�R�>cw0?���>V�N>�:���Z:���Y�*>��O>3�Y�~=V�>�: ?V�?��r>�S>�&���c��������>�$�>�]���1��(�=6ë�G�>Bf>?o�C?�>��[�+e����=[�>'�3?ҰA?J�>�AZ<zy+<�G��������㑾����7>3h��h���I���P�>�<�=�=+f>�B?=a��=�� >5!�=�z��}~?t�>�I��w_
<����@�����=}lD��0r��PW=7L�<w�6��E���G�R��_=���=	H>��>)�>ߔ�>3��>R�K��~N����>�e�=td8?#H?Z0�> ޼�?��ɔ��KA����G�>��z?��v>�b���Խ8�O>�u��Q2>���>�"`�9t>����Gn�
��>�/�>�1�>���>w����d�鄿���bY>pӘ=�y���̧?s�?Y�
T�=Dܾ&�x��*����=`�j>~�>��1�s�־�#W���B�@#8������>h��>�V�?t�b��N�>�]�&�����l�p���>->3.�>�F>M�
��q��j��O������1��f>	P>�?>��?�C?��>PX�>��U��	?��=!{�>\�)>M��> /?�%?p��>S�=�V��M�-�o����䏾�妽MO=��=�.>��=�7�"|����ꤎ�noW�(�a�����o8<�5�=���=�$>�k>�i	?�D?��ƾ�]|��V�>.�E�4�6��a7>�#�=�;���sܾ�Ӿ�?k�b�>��T?p1#?��~>˲�/�2�����m�==h�?5
�>�y�<St>Y=)A��I?H��u�2s
>�ˀ=�u>�g��@������Je>p�>�Y�!%U>(�C?�y?�t?đξ@"��~�о�!�繯>v�
�KV�>tR??_�<?x�=k�J�T��ؖ�=QI�M�>��v��;Ǽ�[d��+6�}:�>k�̽?gf>+�>������7-���c�׍�>�y�>�Y�>���>Q��=m��S0Ҿ�C7?�����SF�z���#>��Y>'@>�h7<�����U0?$�¾�]T������� ��@?2G�?��?0#G?^��<��:M�<i�`>5�>��%�6;���^�<�w(�q>��Z>������i߽��>l��>B�\>j*��2N��D�>��ƿ�5e�ewD�MCž���nA"�u�վ^&�=瓔�$<þ�-���M��7%��yY��Zj�-���l�u�gP��ܼ>P�?&|?9�=v��`��������	����=��=��Iû�;H�����/���Ͼ���8��F������͇����>�덾i�{���k�r���֩=y�>�G.?��׾�mϾ?����=�.&>��=��ӾD�����1�.�a�S?i�!?�����ϖ!����=�H%?A>�=�J��5YC��4l>�"J?��)?l^t�Cn���씿ᦽ�e
�?φ�?;?;�w�*1�7F����	|
?�(	?�<�>�@���#ؾ(�ɽ� ?S�:?��>���D6����Y�>s\?U�E�_$K>��>jت>/\����j��u�CV���^����8>�6��V�����d�GkB���d=p��>oh>�sZ�s��	<�D��<x��SX�̳��Fc�Oj�=&a?�+7��;�>9Ю=&u�>?K�~
���u�����B8?{@�?H�?*;K?"�оC���6=���>Y��>`��>�<>GⒾ��i>���>�߽jB����-g�>72�?��?��x?v�x���޿Ӭ���Q~�q/��<��=�PB=U��=����=����Y���䘽��&>���>���=*.>.��=�+�=>Z���Z�%��p��1c��V�D���@��L��Cd��Q ��|u��B%�I�ܾ�#�'ϐ������P�	����N�J�=�Z��Gj)>��?��>\�>��f=���=<��,I��l��J8Y�b��8E������gȃ���k�8w����G�툼�����?�� ��c=fr
?����\���y>@J_��N	=E��>A�F>H?�>�1>P�_>��&>��=)�>�>�>tvh������D��� YY���[?�l2��]e�0O����c��&/�>��?pr�>�V�*Q`�Q�E��>`m������Vn���˼uBs>�}�>��<���Ś>�Sg�_�������uo�>̠�>�I>�T4�U����G�=`��>�'4�'��������2?^�}?P)/?$!~>9;���td>�@?���>F���E=�<���>,$?�
D?h�?�k>�=2=���� >�j˽?4'����=uС��>Q`
>mW��zBU>Q?�=n>�3��ה���������<<h;�=r��>M:J?�w�>�Dp>W?H�D/�K8F��C���>RL&��Ԫ=��>?�>4�?��>E�*>x
������������>��J>i�J���T����<m|`>�\�=�?�M.?�ս�r��񀜽��=�U�>$�?��3?��>��=w獾���jӿ7$� �!�t���k�Y�;v�<��N�r`�8Q�-�D\��>�<U;\>���>ٝp>�6E>��>�I3>L�>�=G>	�=3̥=�;�;��E��M=�>E<NQ��ޱ�,�Ƽ����^ы�Z=I�2U>������ؼ��?�{?o8c���Ƚ,�5�X�Ͼ�������>%��>l�>�<�>d�=G��ux^��;��z��?G�c?^	�>�N�c<>��=��]=\q4>��d>���=��؎�Yg�n�E��`�>7� ?��>�,�F`��{�������>���=MĽd��?ˤ�?#P�j��a��,����?���>���<>v<G/>��y�4��-7���/���{E>��>�ޠ?�+<�'N>�wJ��g��}Dx�p	޾���=�_�*%�>C+�>�q�3%���� F=���0����,��>�z>8�>�%�>���>�5?�0?j�?���誵>�n�<�S�>��d>�O�>��>��?�ӓ>��i>�I�=��y������H��=�z�<�">XW.>Trx>�{>�a�=���<[�.>��g=���<�����<TҼe��=��=�P>�_
?f�@?V���#���7,>kLٽ�`>\D>�܀>�.�IK��㴾��}��:�>�7,?��?aM>l�߽c|��r��^������>�ML?1T>�$���Y>e��c������$�h>1��w�$�����#����Ž��/>�!�>�x<Ȏ#>��v?���?�~?�A;����vZ�S7l��W�>k꥽�Â=g��>x�0?:h
�?�M��������ي��7�����El��ڟ=paz��V?�ݧ���=0N�>'14=�3a�����{ �a%a>?w��>��}>q�>;(���*��y+?�~��> ��X�c5'� �z�Z�=�@�>��N���>���+�R����u�����>��?�4�?d�J?�4F���ѽ�5>��B>��=J�u�ٽ(yV<�n�=�Eg>.ww������p� b>S/�>%⣽53���[�E
oſg�M�	�"������8E�cd��AJ��8�<F���u�"=��M�:��m��3X���R���F���f�Իf������sd?o�x?]l�=�Qh�r�B��(�����t�>)O;������?޾�����T�����������iiE�]4�
t�������*X���l{�y�+����ߒ���$?߾fv���j+��|s<� >�]2�/� ��f���v��:r�S��?~vg?)Mo���N�/5��%��=�	?���>��u>�I��E�k=�>��D?�{�>����p'��R����=�W�?X��??-??�V��;A��;�C9	�u�??p'�>����0ɾ��ý`
?w3?ݖ�>������&����>��X?��P�o�l>�(�>�<�>[����0��I�3�����>����?>�
������g_�С:�
D�=3�>ju>2i`�N����>���1*J�(D�(t�ߢ.��Ԙ<�y ?�����^>.,k><?>�q%������������J?���?kmU?��3?u��󝽶�=��>�έ>���=?��d��>&��>�X�B�o��) �EH?��?6��?�V?��l�b�;������i
�6�=n�>H�N>`QӽG�J��<���q���E�	}=�f�>Q��>_�H>^�/>��>->c ���(+�by��Im���oo�8����񍆾ó�[��{�龣�⾂����=�!>4���ȁ��n�&�~��24�=��`>�>L3>�3����m�p��.���c��.U��,�mξe��� ��!��<�w�Ls��Cx�<V�����>��=���>���>A|@�i�>I/�>=7�=�.�>�Wo>�y=j�!>h2�>�T�>Q�>�]�=/�L>�;c��vM���t��_~��B�=	e
?s^M?�QW��³���Z�Y���[ؾZ�;?MQ>f��>�b��v���������>��z=��O���G��#>=G�>�Q�>4	�=^�>����ׇ�|y���'X��ɖ>:ࢽ>�u>���x�[=�Bu={��>�n1��0�>s9_>x�j?�l?6>?"n;=�c,>S�?F�5>�C�>�/?k}6=���>���>��W?C�@?���>��=.7Ծ�<L=�[���o���z7>y�-��(���K ��M���齣��=�<9<yc��U=��<����.a�P��w�?�/@?fr�>��F?y�l��2�Lmf�[춼�'�>=Y꽈~7?���>,h�>�ٳ>��%?QԘ>h��>[�y�F��K��>Z^�>�{� �f������s���>��?�wY?i8�=��ؘ�n�E��&��4�?Bq?��?���>4;_(	���ӿܳ$���"� c���J�7;FH<��~X���n�"�,��o��yq�<�8`>�t�>�m>5-C>L�>]S2>��>x�H>
�=}�=h�r�I��Y�@�F=���N]<�hG����iƼc9��%�����O��F�w�_���e!(?-�=?�ǃ���8<�bG=l])�5�����>[�?D��>�A�>VV�>�Cݾ1_c�����g��=pv
?�ˆ?rD?��]��6�%=��%��]?���>�G�>T��x�ǾG�R��|���?�G>?��>�X���T��?B�ݚ�Ǣ�>��>��/��V�?�H?%H)�(Ʀ������ )�U�>
�>C9�����u�g�O�]���~ھȕȽU��>J2>R�?�r;m>�>����+�~�*Fv�$��K8>�̻��Y�>���=����-�վ`}���v��8>i�Z>j��=/��>�g??ׅ#?��l?�|A?â�>~�ὓ��>���<�G1>Um�>��w?|�>�?�k�>?5ג>R>RBֽ�J�ŷ���4�r�0D>Z/�>b��=�k=�;0>�u>b����>���>���4b����?>F�&�׿=Bi�>f�>^�(��VH���+=WH7���=r	}>G-�>��{����N��j4>͋?�x?\?">PP~����͖
���\>PW3?�).?���>�콵;E�:���6zϾ�C�6��>�ڽ�[�;{c��_捾��Ӿ�	�>q�=�
p>��->&Q�?�u?�R?�S)>�1�^����F���k<�6;�XA?Z�?��z���?�HQ:�Ԃ�GFѾ���܊ļ:����=A��=��+=��[>���=΁�=/SC>��<+����M�voB=���>r�w>�?g%t>�">f����	��\?�i=J�������pc�KM��,V�=ׄ�>%�>��?�釽��(��-����Z�_	?3\�?���?�À?k�׽TZ����=0��=��!=�\>��[���K=%`x�֋���ZZ>�
��+8��$�<�T^>�n>������$"B���=̰ݿ`�~��U��F�eH�J��E��j���B�۾�nѽ~с�_��c�(���u�@�;>�m��ߚ�v��4G����?��c?��q>�=e>B��V��2<�h�>z�˾Ss�<��w���L�=�(*���f�9�Ծ�Z��Mp��&�Ȕl>��A������6q��;�G�=\1�>z�5?9�̾�/;0����=��;u�ֽ3���n|�{���@�(E?/�#?/_��M����G��>�B�>]�>�`�=�Q#�]�o��z�>fW?"8�>q��ك�}�������h�?�7�?�MT?ڜ$�h�M_��[� ?ӷ9?�w�>���������ν.�	?"��>*�$>�#E�:�����+�¾�>�w�?+	���C<<?���>���<��������ݻF�G��>�t��*꾵�0�遮�:׈�9�l>���=�7���
����>���1*J�(D�(t�ߢ.��Ԙ<�y ?�����^>.,k><?>�q%������������J?���?kmU?��3?u��󝽶�=��>�έ>���=?��d��>&��>�X�B�o��) �EH?��?6��?�V?��l�b�;������i
�6�=n�>H�N>`QӽG�J��<���q���E�	}=�f�>Q��>_�H>^�/>��>->c ���(+�by��Im���oo�8����񍆾ó�[��{�龣�⾂����=�!>4���ȁ��n�&�~��24�=��`>�>L3>�3����m�p��.���c��.U��,�mξe��� ��!��<�w�Ls��Cx�<V�����>��=���>���>A|@�i�>I/�>=7�=�.�>�Wo>�y=j�!>h2�>�T�>Q�>�]�=/�L>�;c��vM���t��_~��B�=	e
?s^M?�QW��³���Z�Y���[ؾZ�;?MQ>f��>�b��v���������>��z=��O���G��#>=G�>�Q�>4	�=^�>����ׇ�|y���'X��ɖ>:ࢽ>�u>���x�[=�Bu={��>�n1��0�>s9_>x�j?�l?6>?"n;=�c,>S�?F�5>�C�>�/?k}6=���>���>��W?C�@?���>��=.7Ծ�<L=�[���o���z7>y�-��(���K ��M���齣��=�<9<yc��U=��<����.a�P��w�?�/@?fr�>��F?y�l��2�Lmf�[춼�'�>=Y꽈~7?���>,h�>�ٳ>��%?QԘ>h��>[�y�F��K��>Z^�>�{� �f������s���>��?�wY?i8�=��ؘ�n�E��&��4�?Bq?��?���>4;_(	���ӿܳ$���"� c���J�7;FH<��~X���n�"�,��o��yq�<�8`>�t�>�m>5-C>L�>]S2>��>x�H>
�=}�=h�r�I��Y�@�F=���N]<�hG����iƼc9��%�����O��F�w�_���e!(?-�=?�ǃ���8<�bG=l])�5�����>[�?D��>�A�>VV�>�Cݾ1_c�����g��=pv
?�ˆ?rD?��]��6�%=��%��]?���>�G�>T��x�ǾG�R��|���?�G>?��>�X���T��?B�ݚ�Ǣ�>��>��/��V�?�H?%H)�(Ʀ������ )�U�>
�>C9�����u�g�O�]���~ھȕȽU��>J2>R�?�r;m>�>����+�~�*Fv�$��K8>�̻��Y�>���=����-�վ`}���v��8>i�Z>j��=/��>�g??ׅ#?��l?�|A?â�>~�ὓ��>���<�G1>Um�>��w?|�>�?�k�>?5ג>R>RBֽ�J�ŷ���4�r�0D>Z/�>b��=�k=�;0>�u>b����>���>���4b����?>F�&�׿=Bi�>f�>^�(��VH���+=WH7���=r	}>G-�>��{����N��j4>͋?�x?\?">PP~����͖
���\>PW3?�).?���>�콵;E�:���6zϾ�C�6��>�ڽ�[�;{c��_捾��Ӿ�	�>q�=�
p>��->&Q�?�u?�R?�S)>�1�^����F���k<�6;�XA?Z�?��z���?�HQ:�Ԃ�GFѾ���܊ļ:����=A��=��+=��[>���=΁�=/SC>��<+����M�voB=���>r�w>�?g%t>�">f����	��\?�i=J�������pc�KM��,V�=ׄ�>%�>��?�釽��(��-����Z�_	?3\�?���?�À?k�׽TZ����=0��=��!=�\>��[���K=%`x�֋���ZZ>�
��+8��$�<�T^>�n>������$"B���=̰ݿ`�~��U��F�eH�J��E��j���B�۾�nѽ~с�_��c�(���u�@�;>�m��ߚ�v��4G����?��c?��q>�=e>B��V��2<�h�>z�˾Ss�<��w���L�=�(*���f�9�Ծ�Z��Mp��&�Ȕl>��A������6q��;�G�=\1�>z�5?9�̾�/;0����=��;u�ֽ3���n|�{���@�(E?/�#?/_��M����G��>�B�>]�>�`�=�Q#�]�o��z�>fW?"8�>q��ك�}�������h�?�7�?�MT?ڜ$�h�M_��[� ?ӷ9?�w�>���������ν.�	?"��>*�$>�#E�:�����+�¾�>�w�?+	���C<<?���>���<��������ݻF�G��>�t��*꾵�0�遮�:׈�9�l>���=�7���
����>���1*J�(D�(t�ߢ.��Ԙ<�y ?�����^>.,k><?>�q%������������J?���?kmU?��3?u��󝽶�=��>�έ>���=?��d��>&��>�X�B�o��) �EH?��?6��?�V?��l�b�;������i
�6�=n�>H�N>`QӽG�J��<���q���E�	}=�f�>Q��>_�H>^�/>��>->c ���(+�by��Im���oo�8����񍆾ó�[��{�龣�⾂����=�!>4���ȁ��n�&�~��24�=��`>�>L3>�3����m�p��.���c��.U��,�mξe��� ��!��<�w�Ls��Cx�<V�����>��=���>���>A|@�i�>I/�>=7�=�.�>�Wo>�y=j�!>h2�>�T�>Q�>�]�=/�L>�;c��vM���t��_~��B�=	e
?s^M?�QW��³���Z�Y���[ؾZ�;?MQ>f��>�b��v���������>��z=��O���G��#>=G�>�Q�>4	�=^�>����ׇ�|y���'X��ɖ>:ࢽ>�u>���x�[=�Bu={��>�n1��0�>s9_>x�j?�l?6>?"n;=�c,>S�?F�5>�C�>�/?k}6=���>���>��W?C�@?���>��=.7Ծ�<L=�[���o���z7>y�-��(���K ��M���齣��=�<9<yc��U=��<����.a�P��w�?�/@?fr�>��F?y�l��2�Lmf�[춼�'�>=Y꽈~7?���>,h�>�ٳ>��%?QԘ>h��>[�y�F��K��>Z^�>�{� �f������s���>��?�wY?i8�=��ؘ�n�E��&��4�?Bq?��?���>4;_(	���ӿܳ$���"� c���J�7;FH<��~X���n�"�,��o��yq�<�8`>�t�>�m>5-C>L�>]S2>��>x�H>
�=}�=h�r�I��Y�@�F=���N]<�hG����iƼc9��%�����O��F�w�_���e!(?-�=?�ǃ���8<�bG=l])�5�����>[�?D��>�A�>VV�>�Cݾ1_c�����g��=pv
?�ˆ?rD?��]��6�%=��%��]?���>�G�>T��x�ǾG�R��|���?�G>?��>�X���T��?B�ݚ�Ǣ�>��>��/��V�?�H?%H)�(Ʀ������ )�U�>
�>C9�����u�g�O�]���~ھȕȽU��>J2>R�?�r;m>�>����+�~�*Fv�$��K8>�̻��Y�>���=����-�վ`}���v��8>i�Z>j��=/��>�g??ׅ#?��l?�|A?â�>~�ὓ��>���<�G1>Um�>��w?|�>�?�k�>?5ג>R>RBֽ�J�ŷ���4�r�0D>Z/�>b��=�k=�;0>�u>b����>���>���4b����?>F�&�׿=Bi�>f�>^�(��VH���+=WH7���=r	}>G-�>��{����N��j4>͋?�x?\?">PP~����͖
���\>PW3?�).?���>�콵;E�:���6zϾ�C�6��>�ڽ�[�;{c��_捾��Ӿ�	�>q�=�
p>��->&Q�?�u?�R?�S)>�1�^����F���k<�6;�XA?Z�?��z���?�HQ:�Ԃ�GFѾ���܊ļ:����=A��=��+=��[>���=΁�=/SC>��<+����M�voB=���>r�w>�?g%t>�">f����	��\?�i=J�������pc�KM��,V�=ׄ�>%�>��?�釽��(��-����Z�_	?3\�?���?�À?k�׽TZ����=0��=��!=�\>��[���K=%`x�֋���ZZ>�
��+8��$�<�T^>�n>������$"B���=̰ݿ`�~��U��F�eH�J��E��j���B�۾�nѽ~с�_��c�(���u�@�;>�m��ߚ�v��4G����?��c?��q>�=e>B��V��2<�h�>z�˾Ss�<��w���L�=�(*���f�9�Ծ�Z��Mp��&�Ȕl>��A������6q��;�G�=\1�>z�5?9�̾�/;0����=��;u�ֽ3���n|�{���@�(E?/�#?/_��M����G��>�B�>]�>�`�=�Q#�]�o��z�>fW?"8�>q��ك�}�������h�?�7�?�MT?ڜ$�h�M_��[� ?ӷ9?�w�>���������ν.�	?"��>*�$>�#E�:�����+�¾�>�w�?+	���C<<?���>���<��������ݻF�G��>�t��*꾵�0�遮�:׈�9�l>���=�7���
��-��>%<��M��3G���P2"�|�<��?�A�W�>��h>��
>�'�d錿M����=ｾN?i��?� U?$`7?����W��N���&�=1�>$��>�c�=��[K�>(�>���2�q��=���?��?���?�PX?nfm��ظ��G��ꪾDB���W�= s�=�Y>.���>=&]�=�Ƙ<��%�S_>6]�>� v>�Vb>�[>'�D>�+>�����!��c��T���"Y��U �5��c=7����zv��{O��jݾΟپ�ݼ�(ݼ���{����IK�Y���6=��?v�>\�?A�ʾ�e�>(���� ����>�uH�z�$�/X�u���
��tش���Z��z���0��A4�Pи���?8+=9�j>j�>vE>�%�>���H�->4B�=�A	>a��>��G>Y�><��=��6>�J�=�e��=]#�����#�u�f�nM�>�2��l?$������Qa���<&�F�R����b?�N�>�sV��}��Y�����>^ֽ=�Kν� ��bd�=�T*>�ּ>O�;:��{>����:>v�=���=d��i��<�'	�Wů=d#�>z??j
� ͦ>Ɩ�>�De?�|V?g�X?�
�=�-�>� 3?66�>���2�=��ֽ|9��,?`j?�q?�f,?�x�=;ξ4�����=9+۽���<�N[��U�<&�ͽ�Z�nE�����<�>��=��;yk;<��P�p/żQ��>��[?$�?��?+H����%�LF�e�ɾ���>�3�8-A?	o?C��>L�3?�bM>Г�<Ye�>Gt����a�k��>u�>p?m������J�ʲD>�w>̜n?�4j?�c�<]��J��=�}�=��>�	z?�*C?��>W;>�����п��"�j��d�j�����x~<B2�h�`F:<AQ4�J��-C�<W>b5�>�s>98>�>�>+>f��>|�Z>#�m=ob�=�O�;#���/(�n�/=�������<�_���Ӧ9�-ʼ�F��G��<�a�LR�D�=��ټ",B?7`?�����J���E>1���D�	�1>�Wk?+_7?K��>Kي����k�q�1�:Z0>Y�g?��?�[^?����������9�D��>���>�2b>���������>!ݰ<ѽ�<t�>N��=�౽���y@?�ڦ��FJ>��=���_��?�_�?>9��ھ���e�����澒�Ƽ��&�B#�?bؾ�&���^���e0�@����̂��"�=к�>�ƫ?�=�n��>oƼ�t������L��[�=r����`,?-�>NՂ�L w�?1�Mmо�
;��w�٧�>��>]�>�5?�m;?ure?l�2?{�>(���W�S>�Q>���?M?n/Q?!�?9�>1�,>�=�>�=^A�<���/��۶
>�E�=/��=E��>�
C>��=u���.�=��=��<YE��j=�����Mʽ�9:=�a�>Ix��xd?B?⬜�^��� ב��C���rӽQ�;Y�`>����I�%�U:�=�>���>���>���>�x�=�kݾ����(�h7�=σ!?�YG?��>hƽC	�#���Ⱦ�`���j�>�����S�q��Y��p�b��kN>A>�d>A[6>�?;qM?�8L?�[���F�ӽ���Ld�o *=
K�t�?��>���=+�/8�x2��aA!��#���<K'���>+�=vt7<n_�>��=hW�=��>��6���#�������=Z��>���>e�a?ٓ�=e�f<�.a�m5�iIO?�~�Nn�Ջ���x��H锽vf>�7;>I��*�?����w�����Nb?�g/�>$��?i
�?�k?�ҽҝ
���D>�e�>&F0>�((=�����%<U&��K�=�L>��Z��˞�E�B��A>��>��Խx̾��پ�޽&���0<�O� ������ˠ����z����>��(��P^ֽ稾����/��w��=6�<�������caξ~�ǾƑ�>���>������ݽh����'��3�Kn�= �[�޾ltȾ*�$�����F���IWJ������q��H��s�V��a�>and����k�|��]*����;�HW>�W0?��ʾxo��ƈ�q!X=�>��<��ھ�����]���!��R?|�:?//������ ">��?$W�>�T>�~��SW��c�>S�2?dO?Ģ{������b��oX�#̹?,-�?��U?
�i�_8���)�	U;�Mh�>�_4?��>-v���P��d�۾���>�o�>Ĝ�>ӻ�P_���Z@�֬>��;?�E��<>^�?gAk>�~t�XY��_J�HQʾ��$:'B>�/�;N�T�4N�u��56��>��>��uҾ��>���1*J�(D�(t�ߢ.��Ԙ<�y ?�����^>.,k><?>�q%������������J?���?kmU?��3?u��󝽶�=��>�έ>���=?��d��>&��>�X�B�o��) �EH?��?6��?�V?��l�b�;������i
�6�=n�>H�N>`QӽG�J��<���q���E�	}=�f�>Q��>_�H>^�/>��>->c ���(+�by��Im���oo�8����񍆾ó�[��{�龣�⾂����=�!>4���ȁ��n�&�~��24�=��`>�>L3>�3����m�p��.���c��.U��,�mξe��� ��!��<�w�Ls��Cx�<V�����>��=���>���>A|@�i�>I/�>=7�=�.�>�Wo>�y=j�!>h2�>�T�>Q�>�]�=/�L>�;c��vM���t��_~��B�=	e
?s^M?�QW��³���Z�Y���[ؾZ�;?MQ>f��>�b��v���������>��z=��O���G��#>=G�>�Q�>4	�=^�>����ׇ�|y���'X��ɖ>:ࢽ>�u>���x�[=�Bu={��>�n1��0�>s9_>x�j?�l?6>?"n;=�c,>S�?F�5>�C�>�/?k}6=���>���>��W?C�@?���>��=.7Ծ�<L=�[���o���z7>y�-��(���K ��M���齣��=�<9<yc��U=��<����.a�P��w�?�/@?fr�>��F?y�l��2�Lmf�[춼�'�>=Y꽈~7?���>,h�>�ٳ>��%?QԘ>h��>[�y�F��K��>Z^�>�{� �f������s���>��?�wY?i8�=��ؘ�n�E��&��4�?Bq?��?���>4;_(	���ӿܳ$���"� c���J�7;FH<��~X���n�"�,��o��yq�<�8`>�t�>�m>5-C>L�>]S2>��>x�H>
�=}�=h�r�I��Y�@�F=���N]<�hG����iƼc9��%�����O��F�w�_���e!(?-�=?�ǃ���8<�bG=l])�5�����>[�?D��>�A�>VV�>�Cݾ1_c�����g��=pv
?�ˆ?rD?��]��6�%=��%��]?���>�G�>T��x�ǾG�R��|���?�G>?��>�X���T��?B�ݚ�Ǣ�>��>��/��V�?�H?%H)�(Ʀ������ )�U�>
�>C9�����u�g�O�]���~ھȕȽU��>J2>R�?�r;m>�>����+�~�*Fv�$��K8>�̻��Y�>���=����-�վ`}���v��8>i�Z>j��=/��>�g??ׅ#?��l?�|A?â�>~�ὓ��>���<�G1>Um�>��w?|�>�?�k�>?5ג>R>RBֽ�J�ŷ���4�r�0D>Z/�>b��=�k=�;0>�u>b����>���>���4b����?>F�&�׿=Bi�>f�>^�(��VH���+=WH7���=r	}>G-�>��{����N��j4>͋?�x?\?">PP~����͖
���\>PW3?�).?���>�콵;E�:���6zϾ�C�6��>�ڽ�[�;{c��_捾��Ӿ�	�>q�=�
p>��->&Q�?�u?�R?�S)>�1�^����F���k<�6;�XA?Z�?��z���?�HQ:�Ԃ�GFѾ���܊ļ:����=A��=��+=��[>���=΁�=/SC>��<+����M�voB=���>r�w>�?g%t>�">f����	��\?�i=J�������pc�KM��,V�=ׄ�>%�>��?�釽��(��-����Z�_	?3\�?���?�À?k�׽TZ����=0��=��!=�\>��[���K=%`x�֋���ZZ>�
��+8��$�<�T^>�n>������$"B���=̰ݿ`�~��U��F�eH�J��E��j���B�۾�nѽ~с�_��c�(���u�@�;>�m��ߚ�v��4G����?��c?��q>�=e>B��V��2<�h�>z�˾Ss�<��w���L�=�(*���f�9�Ծ�Z��Mp��&�Ȕl>��A������6q��;�G�=\1�>z�5?9�̾�/;0����=��;u�ֽ3���n|�{���@�(E?/�#?/_��M����G��>�B�>]�>�`�=�Q#�]�o��z�>fW?"8�>q��ك�}�������h�?�7�?�MT?ڜ$�h�M_��[� ?ӷ9?�w�>���������ν.�	?"��>*�$>�#E�:�����+�¾�>�w�?+	���C<<?���>���<��������ݻF�G��>�t��*꾵�0�遮�:׈�9�l>���=�7���
�����>�^�*�N��_H��2���޿�<B�?m���>r�f>�}>��'��ь�����b�SwJ?5/�?�;T?0�8?a�����Y����=���>�@�>5�=$ �B��>���>��5)q�0��?�<�?~��?�AW?�Sm�;Gӿ����������=m$�=��>>��޽8ʭ=חK=yƘ��\=�ي>c��>{o>=;x>��T>�<>H�.>P���i�#��ʤ�0ْ� \B�� ����Gvg�|	�yy�����ȴ��񽾮���a���kѓ�L�G�g���U>�I�v��!>}4$?c��>��>��>��>����C�\�ަ���
��S*���"�1þ��־V���f̽���l%����o� $���)�>����@���T>��л�� ;���>���֐�$,(>�����y�=�5]>S�{���W>~D>�k�<��>t{�<\�p�cFn������<jw9>�g7?a
�m����#�X-���ي��a>�ҿ>Ɩ�=L��H���-��X�>�N�ą��hz^��`��I}>�c?وc�z˛�K��=�CA����1�Q>[�>!Qn>-Jl>�k��D��o�޽�|�>q���+J�e >��)?�`o?{�H?Ѧ�=��>Yj>��=t+�=��>qMw>S/[>��>�?�?���>w��<z.�kv>�:󻒝��?��'6��~�<����ִ=��;��>���rꀼ�D >�~j:H�O�就=�Z`=�E�>uX;?y�4?6�<?�齰HL�˂�[Jj��>��@>Uk/?3��>��?Zn?��>��>�r�>�Q=��B����>�=f釿
Ja�}��=�ǒ>G�>��e?>"?������C�lІ���~�??h��>e,>?��?�>+ր=��HM�rrľ�G/�j��pm�݃8�X�ľ�3���8���=hUI�K�>�t1>�~�>�mo>�>�R>�Y�=� ?W-R>����Б�'��Cկ;J}�=٦F>]=5>��0>��=�V�=�n��{X�5�+��a��Z�罡�B�g�=< ��>��?lFQ=��9|�=��a?�2o?���>���>�?�) ?�N��0U��U�������>V�p?-k�>Y�<i�!����d����>���>�R�=|h��1؟�(���d-뼊��>�eD>�-F>1x����2���*���þޓ�>��<�q��@��?�h?E0������,��hm���ž��[��� ��@p<���-�X#	�d�о�6ھ.��ᐽ�h?�?�"ƽ�٪>�!�Ab��b�s�����/躽�>sr9?��>'�=�5����"�H�(��\�2�ֽD��=��=[?���>C�$?%j�?�c?h��>ӥ־Zs?��f�d��=u�>�7?��>J	
?��?sQ.?7�>�u ;��h�-s��]�>F���@E<>!�X>�/��A>�.�>�:={^��;!����:C��=~D�=�^�G�=��o>�߬>�Y�>��? ��>�?>�H)����V�=�'=�>LS]>�_�=�N���>�wC?&�H?b�?H�?>ŭT����зZ�KM�=�^H?�I?:M�>� ��F���������+=�qP>;�G=�/=�v����������=-"�>�=υp>?u?��)?��?9��<�P%�8Ќ��}��'��t>�$�>8�?���������n�g��:A��dؾ_^�<E��� �=F�>�<�=�=�P<��#�>K���%�����I;=��>���>U�>T�>�``>}����8��I?n
���t��񠾮�;
��`z>0�?>�����R?�	��~|�&���)V:����>[1�?�0�?y\c?�F�r��lY>tFT>K>��4<��:�o|�����1>I��=mTx�V���%<_�Z>}>�;��xvɾ�I�`�T��G���hG�?P��w�B�L���Z��Ć���S=�S��!~}��;����p�Ho��;쩽������y�T���#���s�?/�?Z�����;,�%�{[+�j���-�>�>Ⱦ��s�aľK���=�׾<��OJ����=tu���U������q>��۽�x���[;���Y�e����<�zN?��c�d���)���THJ��&���оd���k���9��+󾰐{?�cR?p:I�����QC�{��=ֲ]?qN�>ے>���M/�<�� >��?��?D�=�>��D:���a���?ȩ�?[~+?H��mKZ�������$�Q?p�"?,)�>:���ҽGLƾ]CL�i�>u�����F�1.]��-G� 6ĽpVo?<ws�zZ->d��>hP,>j��||@��A�=`A��v�=&\>e=;�h�S��=A����0�>G��>b|>�k����޾���>�9�u�N���H�������'`�<��?����>3i>)�>�(�����Ή����S�L?���?�S?a8?a����`���L�=��>��>���=��|��>C��>���Vr����e�?�A�?���?!:Z?O�m�$���������x¨�s�=�0��� �=
ɩ�j鼻	�=�0��*��<�c�=��~>���>�ƈ>�˅>Of>>D����b,��ǡ����@1���!�(b�2՛�.���,�?��A���Jվ�VϽ�]��|6�Z2h������=�M��ī�>w�?���><�&?���>��+>ӑѾh�)�Ou�t�E�Z�#��?���u���`�=i����=�޾ⷋ�K�پ>��~����>�h�>	�6���=�&�>��<��?���a>�\�>��
��c>�=V>�>�3�>�`���C�>?˄=��v���j��u�y׽|G=r�F?_�l������-�1�ƾ$�˾ɂ>F+	?gh9>�%�ž����\���>�#]�V�q�����@����C>;8�>|�=Y����>�ՊB���<U�i>���=��[�t�ó$���E=��>�I����=p->��C?v�h?�;?�^�=��?����>>�ܗ=K �Sk�>���>h+?U�(??EfW>�>�-��a.>+ �<��-j齲�ɼ�����}�F�����=V�����Q�wK�=�_�=�hU�qO�=�Q��?/�;��R>�*H?ϽI?�jf?�x%�l�k�E�'�}׾��I>��V>1h8?L��m|�>j$?"�?n�&?I��>�D\�A@<��g�>���=�h��?Z�|_=�(�>bT�>U�f?�?�������>`$>�����~�>q�?���>� �>8C�>�^=��j�迤u�v��QB��z��3��@�V�o��⵼.�,�S  �o~ؼ�=B>�>��d>��u>u~>5�/>� �>�e=>N{�=��=���������⽁XX=x9���/�Gg/����=����c��C���EM<?���7���?�"?��3���ѼH�nE� ���)�>��>��>���>M(>����'I�G�#�ϔ��rH?��x?��>i����=����5w����>��>���=�n�5�޽����������
?.;?or�>}ܠ� �J�R�d�������>�O�)��Dȯ?�Ru?�������y�ŭ���&������g[�����k�Ч7���.�������<�������?��?@�q<r�>)�N�+����|�f�ؾĊr�F�y>�6?d�>��=�*P�lr�|#;�������t����=�A7=��?t��>�D�>RZ�?���>��K>�B���#?<�=U��=g|�>�`�>D�>~f?FԵ>�&?�co>5-�݇��(7���=��˽���=��>"k3=�7[��>B��=˳����h���O>�^;�E�@�9k�:72�=Pj�=���>���>��=t!=���=��m����Bt�=���[iZ>~.����\]u�u�>�0?��>S�M=G��� �3!
���.>��(?@)O?� �>!�M��_C��+�y��BV�>5q�>j����޽�I�o����g>��~�k�i=vf�<�G>C{?�8?π?���:��/�l6���*��+��|H>�ת>�լ>�L��̽̾Tn#�_CK���J���9�'����J�
9�<\�>�y>�=>���<[��=k�D�;=Q}�����=�=��> ��>;�>��^>\7�=ֻ����᾽�I?;��m���쟾��ξ����,>D�<>�V���?�
��}�"ե��~<�A[�>�f�?���?45d?��D�|���W\>��U>(>W<��<����GW��� 3>f,�=>Yz��9����;�h[>�>y>�ȽC˾�侉�D��,ο�(8�\=���a����ᾳ�&�ny8��':����l:ݾ������\��2"��r��SK�(�0�H���Ծ���?��?�N�=>��=n�/��['� �	��6>����Վ�OA�8�ڋ�����%��[��s�@�.�
�>P�9����Q�T���J�:�e����B?�����ɾfsž>p�=���>
%���� �y��,���7����B?I�d?��1�ҷ��_ľO�)=R�E?Q?p]p>E���'>��>M$-?1�?o�j>�Z���&��4��ؑ�?Cu�?�o9?zzھ�yR�.�=�j		�#S:?�ZF?	K?(s�V�>}"�ZA?n/�>�o�>��e������3���?�U�?{���)J>6gp>9�>�=�����eo
<�����;2�>=�'ʼ���%�!�s�����5> ?�>�?>z�.�������>���%O��H��s����Y�<��?����U�>ҫi>w:>7c(��-��A��I>�a�K?HX�?��S?:�7?j��7���=�����=��>$<�>Uw�=�����>��>�s往5r����q�?c��?d��?p�Y?ݥm�	�ݿ�դ��������w��=>�Z>�"��{�=�༮�*�?U�<-g>�us>�4D>�Z>ƙ>>Lq1>G%T>�'����-� Ҥ�������S��������y��l)��ۼ���������Uz�6�� =��鼹\��#$����z ��D�`>�?���>��?��?9��>��;Ex;��K��.�+�<YP���h�_���¨� .h=�������NK־�
����;��>L1콜��<r�>�Q=�>��>�D�ɴI�~T�>��=	8�=�M�>ۜk>`�W�h#�>zt�=�Z�>V��<t�h��`��D�XZ�zj˽J�.?�Y�����j�.��b����ܾbY�>_t?�*I>s��;����X�A�>�㋾�p��+I����;�e��>�??�H>^�V<�q>}����Ǿ��=b��>&>�۸>l�H�5 D�.��<��> �f�=(S>��C?��y?o�?��<
��>�>��?>���=�M_>��*>�׌>��?*A?��-?�J�>�Ę=��B��ͺ=o=}=�Z���>=R�����B�� ��K�۽}����T�=]��=�`=w}�<UY\���̼��ϻ|ϐ>��M?��1?oBA?����a\��!?�������>$��=7(?wmu=��?(f�>��>ۊ?-|�>E�==O5����>�e�=!щ��r��<�/>z�=oj?M8?;(7��1}��A������>��?��?eҦ>��>�"=���&쿰���I/�����uͭ���H=eV���}E��9���s��%K����>
��>���>��^>jr>�'>�0H>/��>�u->�~�<�1j=���,ν~��w�}�������n��:w3=&��<�
�<8t=4�߽�ʽ>ӑ��-_���>J)?�g�R�;W4>�Ӿ� � ܄>Ɇ&?���>"�?�5>& ���h�ܫ�o!;~*#?A�?�X?���J��=Zvҽ��N0?��?��<����Z$�y������Q �>���>���>$�h�(3@���1�Q$��ԍ>t+�9��N��?��q?��ܾTZ����Si��8J��/8���f������Vg����L,�����I5�T���6P?@4�?1��<��>)�7֯�m艿�8⾰]t�HӺ>��D?SZ>��>T��;�
�Y��*�Ѧ)<�o2��_#=��?!~$?�8=?9LI?���>��>v2��m�>�r�=J�P>=΢=i)??B?u�?���>�E?�d�=�j�H����ڃ<R}h=���=?�>j�(>�J��m9��C�5�4=������+�=���p4�|y�=�¤=C�0>��>W�	?6��=Қ�=Q����M�K�;�ӯ<��>i��f X� ���-k>2?�/?1w?�qG>�>����=��/'�pk�>Yg;?G�C??��>�"���w"��uڽ��=��%>E�<:�O�PG�����G���E˅>�=�|>s�C>8^�?��9?��?�#���Z0��ӈ���+���s<�S>|�>���>��<�
�j]�T[W���M�B�,�ˋ��U�<�@��;d�=C�%>$�>u�P=��>�R�<8r����N��w�;hՅ>�>���>x�@>���=� ����˾XI?M����z�I��<̾D,�^�>:>K�����?����+}�H8����=��}�>��?~��?y�d?"B�����\>E�T>A>&lt<,�8�� �n)���4>_
�=��z��u���չ;�^>5�v>1�˽�ɾG��BD���׿��J�x���j�S���	��5����9sн��4D���'�#ܴ�g9����Z�QD�^\ʾ���1%��U�?��?Ӷ˻��=���=43��0����>O�L�M���$���s�������-L���񾩧h��ւ�g;P��>��
�����){���$�=��/m>��?	\��}>1���=���E�)���
�z� ���`c�?I?�3?E+�Ic��Lxɽ�.�=}^!?0X!?��0<<��/�%>���>��>A�?���[��X��yt��?S��?b�3?����N��#�TǊ�FH>�
�>�=G?����`�>��M>��X?��z=�WE9G�n��v���g���?���?u����jO>���>��>���>zJ�'�O���=��=�v�2:�� =y�߽��i�_��>��{>z��>nB	��\��G��>�꾹�N���H����X��E�<,�?���J>�i>��>o�(����MЉ�#����L?��?,�S?jK8?�)��3�����M�=�>]��>�5�= ��K�>��>`�Rr��$��?e3�?���?�DZ?�m����mw��ѻ��W۾6�=l	C>D�?>.W�L�>-�b=�%'�$S$�s��=j�6>�>�#G>��T>7C>n+5>'�����.����i[��WX������姇��j��E)��g�_�������H=�
�ý.�x�ؽ�UG=��o�[`K>�?Z��>�#?G�>�N>����D�U0�~�~h%���
�!@���P�1Ľ� ���+���}�'=�:����M�>%Hýk�>���>$�=�(>�n�>:����>"��>eB���-�>.��>�T�>V��=u�>�m>>���>�QG;/왿���� y�n�1�}=�8w?��ID��h/�~랾�}�L9�>ً�>N=��:�{P��lh%��S�>(x��h��A��d�>hw�>��>~A��ɯ#>�I�����=UϾ9)U=��>6Si:�`>Z\�4Vr�\{<�?�>V�[��{�<���=q�A?^{?�3?�R�==	?�a�=�G><[>�!���"�>��>�$?h�?~u�>ˠ_>q��=_g��(=�=�l��Q��̞�=#�B�gǁ�J >|!=�g�<b_��;#�<�5�=J�_>ׁ>���=ɩ��疾���>��I?TX<?\?�.j=<�8��-�OҾ�<�>eh!�5�l?���>l��>�?8�?s?hJ?}��>�4���>��=&�w�OF^��>Θ]>��>�Up?V+?����:"־�,�=��W�>2̦>U�6?E�?���>���l7�R>�d���\RA��I3�e�=N� <�կ�el�=�bq���� �s����|�/>�܎>��v>i�>aĊ>�$\>�b�>7��>8�e>�T�=/�n�
O���6���^v=F�½C �r���&<>���>H�<Z�C=�9������N�n��%�<��>��? ~�������=���f;���a�>���>���>K�?��>���ƽf���l󶾘֘>Z�~?��>��ڼ����ʽ|qX�W7|>�*?>��׽-���:�V>��l�>}�?Os�>^Y�F�)��1�_����
?kh���C��x�?�]Y?(fȾ���_2�F݂�K�^���_���ɽ⫔��(�������ݣ��䴾"?��~�<?�Ъ?���<��>qv)��]���y����yFy���>U�?�T�>���> v�wc0�K��1����r�=�y�= J>���>��>Z�!?ըI?d ?	�>91��b
?�h��靜>_}>���>V�?��>��>"�>tg>w��:�4�6�d��I_�<�>%>�wI=���<W�R>��c�(����JD���<r]>�@<��=}�_��ɽs�>�?iE\>�4(>��<���uq⽆��,7�>ABѽ�09��ݾr�L�6?s�Q?Y�3?�Ź>DM��\�W��&�R��=$D?=�L?���>p�E��J��n������*>�jx>h�<�G��T&�i����9��' >xhS>�!P>�i>LWl?B�?�d?�m���:���l��	��Jֽ�z=��>,h�>�'�<$��� ;��8~��C\��n���a=/�9��>=�o�=��+>���>��=��>qD�<��t��a��ְ�=Q#�Ys�>��>'k	? >rwp=#KQ����cYF?�g����C���m�¾M�S;�5>�$>�>���1�>�=�9�~�rK����/����> ��?п�?/2X?��]�����]>�n>�>�%v�w�L���kW��� 5>7u�=����.����=��Q>�xM>���]=ľ�ݾN�������@Z����;m�n�����o��)��yܽ�[��������{�¾2�㾸dS���2=��9���q��X���n��?�S�?�����6�=��+�-�D��7�S��>��!���μ8n�Z�=��3�f��1y���4����޹�� �%��K�>Ib�Z[�������=�Q�a��G+����?�X-�����[$�i�[>��(�\��7�����'H���t �w7?L�.?�����%$��5s��=?��"?��>�@���X���<�U?6t�>��D���L;����=��0�?�ž?;]#?!�"����ھc�ݾ9�=>�;?�	�>�.���>h����|�>�Z`?Bþ:����y�b7��>�3�?�`Q���=��>Krk>5U��6���UO�_�q�s^U�`�'>�B<ko@���.���N�#K}=�{>��=S%��f����>�^�*�N��_H��2���޿�<B�?m���>r�f>�}>��'��ь�����b�SwJ?5/�?�;T?0�8?a�����Y����=���>�@�>5�=$ �B��>���>��5)q�0��?�<�?~��?�AW?�Sm�;Gӿ����������=m$�=��>>��޽8ʭ=חK=yƘ��\=�ي>c��>{o>=;x>��T>�<>H�.>P���i�#��ʤ�0ْ� \B�� ����Gvg�|	�yy�����ȴ��񽾮���a���kѓ�L�G�g���U>�I�v��!>}4$?c��>��>��>��>����C�\�ަ���
��S*���"�1þ��־V���f̽���l%����o� $���)�>����@���T>��л�� ;���>���֐�$,(>�����y�=�5]>S�{���W>~D>�k�<��>t{�<\�p�cFn������<jw9>�g7?a
�m����#�X-���ي��a>�ҿ>Ɩ�=L��H���-��X�>�N�ą��hz^��`��I}>�c?وc�z˛�K��=�CA����1�Q>[�>!Qn>-Jl>�k��D��o�޽�|�>q���+J�e >��)?�`o?{�H?Ѧ�=��>Yj>��=t+�=��>qMw>S/[>��>�?�?���>w��<z.�kv>�:󻒝��?��'6��~�<����ִ=��;��>���rꀼ�D >�~j:H�O�就=�Z`=�E�>uX;?y�4?6�<?�齰HL�˂�[Jj��>��@>Uk/?3��>��?Zn?��>��>�r�>�Q=��B����>�=f釿
Ja�}��=�ǒ>G�>��e?>"?������C�lІ���~�??h��>e,>?��?�>+ր=��HM�rrľ�G/�j��pm�݃8�X�ľ�3���8���=hUI�K�>�t1>�~�>�mo>�>�R>�Y�=� ?W-R>����Б�'��Cկ;J}�=٦F>]=5>��0>��=�V�=�n��{X�5�+��a��Z�罡�B�g�=< ��>��?lFQ=��9|�=��a?�2o?���>���>�?�) ?�N��0U��U�������>V�p?-k�>Y�<i�!����d����>���>�R�=|h��1؟�(���d-뼊��>�eD>�-F>1x����2���*���þޓ�>��<�q��@��?�h?E0������,��hm���ž��[��� ��@p<���-�X#	�d�о�6ھ.��ᐽ�h?�?�"ƽ�٪>�!�Ab��b�s�����/躽�>sr9?��>'�=�5����"�H�(��\�2�ֽD��=��=[?���>C�$?%j�?�c?h��>ӥ־Zs?��f�d��=u�>�7?��>J	
?��?sQ.?7�>�u ;��h�-s��]�>F���@E<>!�X>�/��A>�.�>�:={^��;!����:C��=~D�=�^�G�=��o>�߬>�Y�>��? ��>�?>�H)����V�=�'=�>LS]>�_�=�N���>�wC?&�H?b�?H�?>ŭT����зZ�KM�=�^H?�I?:M�>� ��F���������+=�qP>;�G=�/=�v����������=-"�>�=υp>?u?��)?��?9��<�P%�8Ќ��}��'��t>�$�>8�?���������n�g��:A��dؾ_^�<E��� �=F�>�<�=�=�P<��#�>K���%�����I;=��>���>U�>T�>�``>}����8��I?n
���t��񠾮�;
��`z>0�?>�����R?�	��~|�&���)V:����>[1�?�0�?y\c?�F�r��lY>tFT>K>��4<��:�o|�����1>I��=mTx�V���%<_�Z>}>�;��xvɾ�I�`�T��G���hG�?P��w�B�L���Z��Ć���S=�S��!~}��;����p�Ho��;쩽������y�T���#���s�?/�?Z�����;,�%�{[+�j���-�>�>Ⱦ��s�aľK���=�׾<��OJ����=tu���U������q>��۽�x���[;���Y�e����<�zN?��c�d���)���THJ��&���оd���k���9��+󾰐{?�cR?p:I�����QC�{��=ֲ]?qN�>ے>���M/�<�� >��?��?D�=�>��D:���a���?ȩ�?[~+?H��mKZ�������$�Q?p�"?,)�>:���ҽGLƾ]CL�i�>u�����F�1.]��-G� 6ĽpVo?<ws�zZ->d��>hP,>j��||@��A�=`A��v�=&\>e=;�h�S��=A����0�>G��>b|>�k����޾u��>�ꀾ{2$���?���ھ�V��<L�&��>U�_Vѽ�f?�&�>�:��픿��q���=>C�a?�c�?��?�Y?j�I����c:>�p>"�4?	��>6"��sɾ��H>��[?�d=֒���K$�~�-?�{�?v�@"�b?��@�hp�.����*��n�՜�=鏛=a�4>���G�=5}V="Fz�ٵ�<^�">�]�>i�r>F�u>�3�>��7>�v,>n���Y#�ћ���0���1�,;��i��M˂��l⾁᜾:���>׾�t��y�0���� ]�<�)������3=�-J�1��=�??nx�>��?Aˌ>8�9�,]��4:�;���^�ʾ�?>�*�L��XS�����P�`(���Ѿ���v�����$�p�_?����m�=I�>k�^����>E�=ww�=	O�>��>��>F>�E�=�>�>��>�=�=��->�>�=�|���q��I�v���@L=�>?񺒾�v��!�"Y�����j�>w4?�j>��)�G�����ZE�>C��<^o�?)��岌=0��>��>�|�=
�w;�R��6~������=�S=>+C=�e��y����ʽ �>���>��Ҿ�ͱ=�Cw>Y�#?�Nv?n�7?o�=8>�>p�R>�`�>�p�=|.S>�GO>Y��>Gc?C�7?�<1?���>�Ĺ=��[�G+=S=��8��E�|���"m��h4���,</A��<F=���=��<Y-�=1>)=�<�W��;�E	=�?a�Y?ű�>^��>���g��8����=w"�>0�w�Ϻ=�6X>b?��?��>	�F>y��C�_���>iL>2҆������7�E�k>.	?N�V?��-?_҂��N�<p��=rD8>�>>?�R?O�F?(G�>q����������N��[ �[uM�RDH���Q�;)��ɷ�M\=nZC�~�)�����DL>dz�>!�>ſ�>\��>]OT>-�|>�>�vM>�Q��χ=Ⰴ��%�Ƥ�f��)�P�>�=���;!=��Yc���渽����ĽCz��5fs�����G�>s�E??�j>Y�$R���0�����<{=j�>W�	?�>&�l�s?��N_�óU��y���[�>�L?f�u>|^�_�Z=0ל��	���>�r�=�rB>9�I>^^������񽢝�>��?Cī>��|���f�ex�P{�j+�>���=i��K�?�\W?
��uRg��UZ�_����{o�=�bb��t����??�O�$��4@���7�%u��7�7��>x�?~�o�L�
>Hi��a��Kq����ns�>��Z>.�>54��Wk�CY�;���a�W�W�E=�+>�o�>���]���W?��d?q��?�E�>��=�,c�{|?��h>��_>'�/?	�?$@Z?��4?bA>>o�>��{���y�����?�����������*W>���=6�
�e�����*���û<��ӽn�D�뀘��W���<�T>p��=P\�>�F?�A�:�3*�5�P>�þ����>�>�?��ý`6����>x��>S�@?jT?Nc�>�4�����w>����D-o��31?�	?&�)?l�;'(���_!�SZ�=Ο>/0�>�>�Fx���,�|��!�>��>g>uΆ>�Dz?)_?UCS?FK=Mi�r��{D�'{=�|N>�^��!�=,nƽ�¾.U�t�?���/���L�IS����3�)�d����)�>��v>�>�D>=#>*3=ט��@�D�!��p?D��>��?�>�<,(!�6Zܾ�Ȼ��b?�����gľ��=Փ��RF�>��U���Sܽ�y??P�>^&a�\�ȿ��^�u_<?��?���?U5?T���y�;n��>5��>�>ok&>rZȾ�랽ܭ��C�m=���=�qD�f�,�	�E��;}�=����� �D�*�Z���w��J�Q�uǸ�6����]@��꽳��h�Ѿ{��F?���⵾h�`�1�<���g�A�l���� ���h��ky�?���?��ݼ�
,=dKk��m2���=�,��>�V����G��%����Ҿ1p���Tk�����43��+��d ���j>aۗ��茿��v��J�}ݬ�7��>ەR?��*���˾�����{=��s>�<-��z��m%��3��=G b?kk?���15�`���|�{=�a?�](?>w�=�;S�F�	aq>sU.?�e?Jsk�
������ɢƽ���?H�?��?�ch=߳{�R쾀{6��[ ? L�?U�?�f7���J�)���w>�bD?��=<V:�!���D�Pt?�Ǐ?2�,<>�Q�>k��=V���>p�nI�M]�<nDK>���=��:"�ٽw�1��N佚�>�>��C>��y�3�W����>�	f�`�%���S� ��L��D���
y?(S��}8�<�_?�B�> �,��礿0�d��t$>�Ok?\Œ?r�,?.W8?$����^4'�L�1>��?�ڼNn�<����`>14*?�𠾌���Ӆ)�u�`?<�?n�?4_N?��f����צ��ܼ�����vx�=�`�=Y�2>����+x=bt=���pk�2�>K<�>��w>;�p>�^_>bTJ>��2>����dR!��¥����5m2���%���ᓾ_��<�+E��S���K���<��z��3����*N��U/��]���|��rd>"��><�>b��>��O>F�>A⧾�ƛ�~ʐ��n��"L�zAK�Us5�fS1��̴�T>����d�����}*�������>A�����q>�y�>�:A��P>��>�ɑ��~>+��>`��=Wj�=�O�=&�k=1��<e�5>��x�0�0>:�9>w)���5����U�񭾵9�=��P?G�j�>=��PL��/��mu��s>�?�p$>��3�b^�����Ί?�8Ҽk9��J�]�i�S��y�>��	?�b*>�&���"������(����=;��>&>Mt@�m�ľ�2ؽ�th>��>�Ծ�3�=]v>u(?�hv?h�5?=О=Q�>�d>��>���=`ES>RN>@�>J�?L�6?/+1?#9�>j �=vvg�l=[,X=��@��c�����G���@��0�<�(���V=�`s="��< yo=m�+=	ݼ�ɭ;��=]�?�LQ?�w�>�`�>w1h�z�P�8�+�me>v�a>Lq���>K��>bz�>0�>�1�>���=[ܣ��D�,ȳ�}(�>e�>`����5���(>���>�~>6ZY?-yx?�f���ɾ��>đ�>�y?�?F?�mE?���>qP�=���@|������%�H�,�),�=���qt��,������P;-��7���3�>U��>P�>��^>��7>�v7>&.>.�?�͟>�B=`�˽���R�߻���fsR>΄�<�=��!��8-��x��}��<S�;�L�=��]�u�P��.�>��8?Q�=-���}̽׭�WJ&����={f$>��>oYK>��{�M/g�s!`��n���q
?&�v?��q>�Q����a�|p���>M-�=���>���>�9���Q��:>��<-l�>w1|?}��><�Q�+oA���4��&��{�>�q�=� p���?($j?bʫ����)���W�����u>���z��i����)��+��?�����������ؽ�z�>z�?�qT�^��<S����,h�{�3�&�'�����>�ga<�����&�оt��/�(�z>�&�>)�����T`?
ox?���?��>ī����=�vk?d��<�%?^x.?�h;?+Q?|w ?��[>-��=�=b��+[��z��7��/���#��<�9�DZ=��>o��;�A���<���,�ؽ?��̲ ���Q����z6�;΀0>��>���>�=?_�<�ʅ�!�>9�==�H��=����-?��Ҽ�X�:��>�?��Y?��7? ��>u�%V@�Ϭ(���'�^�9�˭/?~m-?1�?�7�<���z���2,���>U�>�8!=
I��w��v@���Ľ���>뮒>(�,>P�)>gk?�D?7{,?`m��oE�v[d��H�к%��N;>�k>=�=C��<8־��T�U�^�3x9�j�>-';��}��7�<e�3>�>�=C\>��ͻP�=�=R��Cн���W�<#�O��m�>9:O>�>��,>�: �g���Oھ��c?��ɾ��ؾE?5�Xؾ1��>���-���s���??�͢>�퉿����w�Q��IV?Vc�?��?;X,?@���M��2�>���>xn>D�>`6ɾ�`�=��	�+f-> �>����i��²=��>-z=�,�$f�o��ka@��շ�8�5�wN��\\�������-�����#.r���w���R&��m�o�9���QZ��M�BAb��ݾ:E ��δ?���?���=r��� ����*�QȖ��qT>Z�׾�x��&��Yx�܊]�Fg��nݒ��)���CL�P�c��Q$��B�>B�罍a���
��y��/9>/�?�4�?������U�uGO>*� >���=i	�vq���c��;�3���U?.�7?N��s;=<	�^>4�7?��>M�2>�SG�!ێ��>I@?s�?�� >"9��@���Ύ��\�?\��?+�?wq>��f���侱�ɾcc�>���?��>%R�iW���F���?�h?_̲>��_�	֢��D��<?e�?k���c�7>�2�>��>����fa˾ �+������ei<b>��>�����t��]�Y�&����\>c?�>��t��g.�eê>;Pf�	NU�Kkh���/����%�S�?\D�����\�>�x>���X~��.�e�x�;�,?�Ơ?:S?apK?>p��b��:���\xJ>?^?��>�n=ֆ��	��=�I?a��b����A� 3?A�?py�?*ae?_Z��濼T���(��Ȫ��.>]U=�|�=�����
=
K=�B �1��<��6>,�>��>��v>Q/�>85K>��Y>������)�ۢ���"���-@��p��E���O�Z����w����,�ξ�¾�+��JH�<�1|��������P�<]��]P>�K?W�>�<	?��w>�b>hŰ�y�L��#砾�+4�p���P��HnZ�κ(�b7˽�l��B�𾀼����(�.?�v��X=>��>��t��->�W2> ��_{>�L�>;K�<��>�1�<�p>+�=0Aq>�$�	�|>�J�=���ꨀ��<8��_S���;C"D?ͤS�h��5��ݾ���If�>��?��T>�x'��Δ��y�H&�>�G���a�9?�>��gi�>�2�>���= �� v�z�s�T�9�=�a�>7/>Ǜe��ŋ�����=�0�>I𾾘���l>�b?�R|?�U&?�h>�)�>;a=�w�>/�>R�@>��=�>JS?�5?��G?	�??�=w�8��Q�U�#>�ۀ��!F��]������u�F�,~�<�r��O{<@dS=�|�<�=��=<���Z�g�<��>��V?u;�>Db�>����p�g���Q�,!����>�o�=9A�<�g�>���>���>��>U�=�拾c&�x�?��>��>�Ɂ��v��硻=���>__�>*bg?��L?580;NI����*>`�>�'?p�0?S�C?c;�>^d�;��K���l����x��S�����2������������`���}�3=�|>tS�>��q>IsX>�+>h�>g��>�;f>�ő=7�_=�~'�u,<�H���c=~S��}��� Y�`q<�ɚU�K������������Ob1�Ս轱��>=a(?��I;���G��A��E뾋I�>Z��>�_c>gR�>�2>ɭ�Ha��H���ܽkn�>�b@?�i�>S%��(3=�z�%�v��:s≯7>̅�>K��<��ͯ)�$+�;X��>�?�Ƞ>B(F���L�Jmf�j��� �>�,6=D!�����?�b?��ɾ��LA��e�4�%��G>�A�z
��T���t&�Y�8+��9Gq��l���=��W�>L�?�Y�[�=��農�������B���|�>rv�����>��=.0&�3���:�[�Q��0���_a>V<?����P�=b�2?(�?̥?7��>���=�B�<i�w?]y�=�ǐ>w��>Y'8?�IZ?�f?��=>�'$>��z��؇�X0�yR���)>�>��=KQ�=�{�=gw�=\�d=9/�=��N=�e�F�<�Ϙ�B/g=i\�:8��=�>�v>c��>3�<?4f��e��#�>*~�Ң���Ǔ>��
?�=�.�q����>g+J?�m+?4�>n���`9��'����@s�w�?v�?b?��=�;ý���)<�p$
��\�>�CѼ����B���񆙾�z�R͙>N��>`@D>�>�ZS?P�i?�C�?�C��؆��g����nv>z�>�z->mU>`�X������.�t.�Av5��3�H�$���v�u��/�<���>�c'>���<p(�>sꦽ�F����r��7��V����>\��>m��>|̶�C���ٮ����xc?+�׾7Tʾ�b������ݦ>&;�>	���O�0�8?�O?ᡇ�_Zȿ��龬3~?`�?��?�'?�m����0�}E>,��>��~>5��=�(����=���K
�MD�>������ߦ�=�z�=�#={�:�X�达E.�ý�׿�z���%�(����ؒ��k�!%�������i�������������v�W��Hս��&w�ev�����������?���?�v=�:���j�֜)������͂>�4	��1R��9žL��X�Ҿ+��zO��&��=q���W�ڥ����=L���c���p���uU�`�;��_�>�?�_��g���	��@>��n>���u�S���¦��<r<(sZ?��M?�龾�+�-|�\7�=:!\?n ?�i�=�wE�˕�h�|>��@?U�M?.n�=H8���q�b��=r�?j��?پ!?<R��{]� 3 �nМ�IgD?F;W?a�?]����a��6=<\.?lN@?/�>Vz4���}�K ��D?]Y�?��T��@>�R�>���>^��_����M��~��`ގ=i��s��l��A�.��=�=7>AO!>Z�v�S$���V�>����6iC���N�����zW�F̮�˴�>Vy��Ɠ,�m>p>&uN�iG��ީ@�S��=��j?�K�?��?@bI?���<��Z��`y2=yD�>���>���>}/Ѿ�(>9X?*���F��l^���+?X.�?"��?���?�=y���߿ʫ�10���ڹ��)>�˚=��>Y�)���=6��2���\�h��=(�>2�>�	>��Q>ch>�>���u�&��ܚ��s����?�����w3��#���]����� ���>�о��ǽ*����䜼�������>�GG9��:>��?H&�>�?~$O>*������=�3	��d��K���M��VF�x�0�K;3�߼�:/=U��6��� ��*%&��/?�of���v=�_�>�ڽ�5�>�>>�=�/>�
�>m[�=_�1>�;ֽ`��<h��<��A>�۳=��(>�.>"����Nb��'q�5���WKV>N0?�V����[���u��puj�>z!'?�	>�]@��������i�>�g�=��ѽ� ��S����=�Π>ĩ�=�V��L�;�����н��=�S�>�P��V"��O��f,��W �t�>��Ӿ�5�=SLs>�'?ڒw?�6?���=��>��a>��>e��=7P>$T>�+�>Dp?�58?r1?���>ߑ�=��e�j�=5�:=t�8���8�����m� �w��9�@<-�0nM=��p=k��<\�Q=�>=��Ѽ u;�N=o[�>H?���>�>?=���<L�ݙQ��y�����>�ґ��v>K�>;I�>X?�>S�>�d@>�e�8J5��>Ծ�[�>���>|}���೿[#Q=uo�>�ӽ>U�K?F&?�e�K�ܾɺ[���>��?�C!?s�X?L ?��ɼ����;�'���~~�I��u��<������\��վF,4=Ԕ+�(�����S�z]w��ޣ>���>��>y:�>�M@>g>>�>�>��=���=�J⻸��9�M�=�o�����Mz=��齪�=�8�=+�z�i﷽����E����<E�	=_?��5?���>�zK=�i���8�oO2��?��?�N�>� ?V�4>R����q�hLH�P�ƽ� ?L�?�(�>�����ͻ��{-�LƦ>y�f>F�<>W�>�:Լ�@�<��+�����
?��+?�S>K�<SJc���a��Ʃ�?*h>g��=v����?Q�J?��Ծe�����?�|R���2�XZ�p=�ǻ����:�4�;��fz��Ym�I�������y��>*��?����Z�=}V,�3��tC���W�1��>��
� ,?p��=*)����Q�#|о��^��Τ;p��=���>'I�J�ཫ5Q?C�?�U�?W��>(�9��1	��S]?$Z�>���>�w?��1?Y�m?��?���>�w\>4��7����A�kU��{9>�N�=Jb�=��<���=���=��:=t�;&d�<�K=`^��73�K�8=v��<T-5=��=Ku;>�B?x�7?Ǐ���������=Q)�<NA��,�: ~�>���S�uB��>`�?`'?'��>��P==�"����2�Oj��$� ?͠?�?w�=FA�<Ȕ'�� ��8�5>�O�>TOc=�ξDs���-ƾ<AD���>��?�*w��o>i3[?4�[?#u�?�7���j�Sp�������=vľA��>�9�>�� ��-�����.Z��w��#*��g����/�>�=[�>J�T>���>b�-=�r4=�w����ϼ^�J�.�=Zh��]��>%��>v��>�ɇ>+�"�����5设�ma?Y��+"��臾RΒ��3>Q�=l>�e��4�B?��?V���+��T/;�ƓH?r��?]x�?�`2?s̾g���]�>*�>>	!�=~nl�o���,���U�{�9[�>YU�X�2���>�\1>�B�<{R�>����J�����^��i�V��T�?b��R�����Ѿ�T4��߽ܔ�}H���
��'��s�!��~��\�=�:�����;��!0��7�?��?_�Ǿ݇_�7f��YY5���=�G�>*G�̟�f��q0��vm�����#���A�^xO��\��>��}>/�">�:����\�&%q���~���<?���?�O�>B⾒���5<�E>����Ӑ�Gx��\���EN=�K?�\(?�&�������g�+�>��G?�>�>Z,>݌���J^����>Vd.?�}�>ϵ>}�o�1A��─���?Ļ�?X�?��^>�{�"�
���ľ��T?��b?Z�[����\r����NN?�@N?2�W>�����;���'B?R��?ˁ����=�[�>�r> ��;/�q����n�p��(�>��=۴g������a�8�����Oͮ>��n>Q�>����_
?~�ľ�P���]�2ˋ���>@׳=E:�>�����!|>Z��>�?������l	o�4ir=Pu?���?v�=?�_C?�/���㾙�>��>�>�>9�>��|>e����->܋?���=���g��5,?�r�?�N�?��m?��r�F&�L1���𰾻�z�=�U�=��;=�le���=|[
=0w�=��w<��(>O�>�s>�\�>��`>��>�E=>����+�D���䖿��=���%����+����x�����J�K��\`þt���Ϫ�������0���0��o��9�H�ȟr=�'?���>�<�>ө{>.=�6W��C,�m)�BN�ZpR���� 
F��U���{1�x
ӽH�e��*�"p��ȷ�Ҙ8?\������hR�>��;�0�=K0�>*ި<��>��9>�+>�Z>p�h�(�8=�F<��=��A��S!>u]�>%����(��{�P���x�ץ>	w<?.1�́�!�u���ݾ��tT�>��?"b/>��O�M;��k\�*�>�u>���zn�)�6>��>��?��>�v><�U���O���Z�F�1>ʸ1>��>T�=��s���@�L�n>��>��Ѿ��=)>t>�D&?dVv?[;5?�0�=S�>�hV>Yۑ>x�=F�C>PS>ꕊ>�?�5?<.?�8�>{��=�=`�C�!=*�6=�=���f�"����UѼ<{ ���<.�B��E=��u=/B�;�F`=��==�⿼�s�;8Z�<��?��A?̺�>���>�褽��$�}R$��Lk�7��>z�h��]�>��>��>�^�>��>�LE������ �6�}�a;?���>H��������ؒ=�=?]%?��\?�@Y?t�> �8��>�C?9�?�v5?ʢ/?���> N�=�Jн�K��[���~���0��Q�JN8��O ������c���=�H����x<��>^��>�?�>�b>�k.>u~>pbJ=���>�	l>l(����>Rҳ�Rj�M 4>kI`��þqcd=	[��g�O=�O=�;���_Ž������ý���<t5�[]�>�8?Ӻ�>���>�w�-�F���B�/�>��z>�$�>���>4怾��9���x�rY��Nc<�(?��n?�O�>�p3���<&����P�=W�h>�|>�I>�c����/*���p�=��>�Q)?��>5���Pz�R怿\���-+>��=[D9�2,�?̿m?��yu`�̄A���H���&����=�\��6Ӿ�|��D�yB�8w���d���T�t�ǽ��>۫?�m��K�>�� �6^��˾{��!��y2>u(=)�?�>>�p��M_��B�d\ƽ!J>n�>��>��2�U�ֻNB? �?86�?;=�>w[�;�_��E�?�P<���>��C?r�B?��W?%h
?�_z>�d>�U�����_"�6���\<A=j�]=�ӧ���k<Jty=�#�<�e�<=�	>wn,:F��~㪽bv>���L�*4Y�"�G=�>p�P>��?��??� ��h�b2�>:X!>_~��
,�>�@?t1o��!�=�w�>"	�>^a??_�<?0�>�"��)�k��2����[E?d�?��?ίP��]�����U,�'w�=���>L��<�P���˾���M��t2�>���>f�2<%�a>ϣd?"Y?%:f?Z��'N��r���A�����m(:R�>`�8=�������\�4��\���7�G�&����-='�(�=]1"�:l4>�"�>�ͳ=���>�����s�̯��2��=��7>Y�h>8[?n��>"�=]Yq��T;K�l���L?gt��А�g<�=e���ڑo<����%���K����?I���������աp��U�>�$�?"��?'�?��Z�#�����>��>��	>D�Q=�ԾD6�D����}=�>N��F��y��<A����4)>]�/�!��a����ص�jQ��v>F�~���1|��}�F�B��ʅ��\����U�=�+�Ԕ��5s��)_�Ꙁ��߈�Uʯ�����c���a�?0�?��=�90<h�c�2���# ���:>�������{��j���E������y���MѾ�+�B�?�ğ+�5F�>�T
>l֞�R���BKH��Gm�p4B?���?�����I	=��9>l�=����y���5��Y=$�h?��?�a�_���B��>� �=��?.��>�O�=&�پףb���>~L)?ex?L{�=S��t
��
�=�X�?N��?<�?��=�`f�+���F&� r<?+$G?f��>�2���)��&>�o>�-?��e>�t��,��`�#��6�>�N�?��;�k�=oXG>A��=�G'=-ύ��ؗ��ѽ�)I>�?u=/��=��n��u����ݽ�H>X �>�m>����5ݹ�+�>r��j"3�9{�X����%�s�|>��?2hӾ�Է���>i:�>�9¾���i�t�?�N�^�f?�a�?�r>?�G'?�ќ�Y�(��{M���>)��>�>���s5��T[>;��>���g9E�!���g�>���?�O�?��\?T1�����g��ў�|�Ͼ���k0׽�	�=G� ���D>��=JP�=e��P�(=S�>! n>6��>�b�>/>��>O����.�fЕ�ik���Z�Y�F���'�V�0���þ�Yf����G�I��n������½B�6�yA�k�*���a��&��J�=�"�> �>ٗ>�a�>��u>`g���ľ=4G�Cn��A��-����Lf0�+������:r������@��>(�����=T�>��V���`>�}�>.�;�z?>#��>� �=-�=�ޜ>LA>�u�=���>,�I�M�8>�G;q���i�h�ȭA���	��D��D.?��'���<'���J{��O�/���;}�T?h,�>�1G���ÿ������?��ƾ�!��J�N>��+>w��>
	�>bﯽ���Ӝ>�>�����V��-��>�/E��8:+��y�;�>��>.��>
�彐⛼ĽzE?R�F?��a?Ȇ=���>���=��>�!�=n�>�>c��>��?�4@?�W?;z>�=�䟼�">,�<��������l�k�J�I�/0�>�fU=v��V'=g��<����c��=�ŋ>r�߽����Rh���V�>�M6?�L-?�8�>�V���U��<m*�n�t=cf���Ta>�Ok>hm�>#�>���>��:=�C�=#>�.���i�L�>���<Ŷb�T�����%>��?-'?Z??3T�pđ�L�>(Z>Pu��⏚>�7�>���>u��>P7�=� �+;��յ�&7Y��J]�:���H�~�:""���<X�}�����ƽS/�C�u>�.�>���>�I�>�}�=�jY=���>`�+>��=q��=r@>�DR>6�=GI�<C��L4����=�&,�<3�=@��/����L=Z9�=������B?{v?�/�>�$�<������Ҿu�@����>��3?�U�>Ȉ�>�Q�>+���Y�u���*�2*E�E$�>C�?|�>�j½)�<����O���]|�>�-P>��>��������־�7>�=>��?6�?.N��df��/��=�����>9��=m�>�u�?.�t?8O�j-�������*���ֽ+1�>�N|�d�=v䳾
d���ƾ'�n��l4�>��$I�=�I�>Q�y?�߉>LO>�e3����^��8ҽ4�>wn�>[5�>wW>h˽_�߾��X�Ϣ��Ӓ>��d>+��>����֗?#9>G�>��?��?W�>5>O���H?1,^�c�Ǿ;Q����?j5h?�?!�$?�F,?"B>�����"�
�7�V�;�� <O
żMq>��6>3<g���">��a=S���C� ���V���>	�M��|$>��i=@r�=y��=��>ǁ&?h�:>C&,�'�r=-����=^���a�>t�>�y���ߛ>��>� �>3$A?%G.?�Xq>�ؾwD����:>�d>?� ?�)?>���<9JL���u���պ� ���^׾�꯾��C�;��_�3�Ԝ/=9�D=��I�^Tl>r+}?"z?j;W?�ό���+t��� �'ˌ��?�>�`�>�2`>�VS>���F&&��+G��	�[��t�+=��d�n��<�����'
>���=@���2=ߙz����� ��;�}�9v�s���=�S�>9��>��=>�-�<��Ⱦ�v�MPE?��߾]x-��������U<d��<��_=����#A%?�^�=aK��%��,2��4�>ԁ�?S�?�?���x8��Ǫ	>�>��=�J=�.X���U<`��<�R>'C���4��ٮ�����=�W,=��>=�Z�c⮾�-���=��ȿ#SF�������I��������4���*l�P�1�s�̾�F��j��eN��J�F�y�o��/���)Ӿy�;9�?���? Ô���m�v1N��B���e����>D_þM�u�N��	>�����l3�L������8�ge��;s����>a���)W����C��$�dc�;4��=�"?�6�l�b�0�]��������L��\�$���s��X����ؾ^V?0�?����,!��w�p������>���>���>j#������>�>.�C?�?��A�r�}�����s��Nܸ?���?�'?�w�����1��/��ߗ
?˔�>?'?�nҾA{�C��>���>��=�6��?�8��&���`F�Yk?R��?DM���">�o�>k�}>�3������(����=Pj�<=@>ME<=�w<W%��ߙ=�6>��/>EN0>��@�V����>�+���N��H����1�).�<��?j���8>3i>QP>R�(�����Љ�i>���L?���?k�S??b8?�^�����o���蕐=g�>�֬>$]�=���$ݞ>���>�h�Knr�%�Õ?[I�?Y��?UKZ?&�m�����g¿{����߾'�e=r;�=�5>���t5>���<�ñ�}���Yg>=B�>��c>c�>W�>��|>�#>�-~����f���C��«H����sd�`��m�x����쾡m���9�������e#�Fv��m7)��m���� ��>> �>���>d�? :�>�;q>�~����������W�c;�)嗾��\�J���=~�=o�c�Ͼk���B��{���q}�>�@���ج>G��>53*>��?>��>�[B���q=�q&�j��X�J>�.�>P�>lj>����ެ��Ľ������M�@8	�V�=��ھ)?x&��~�����>�\ �I^�<��>Zg�>�9s�ӈy��|��m�?�Ν�-�m���b�弙P>�ݕ>�;>���׆<s�1�O����9����>�#>�ԡ�~��[�0��ѕ>%	w>^���/>� ��Z?��?��4?�Œ<TV�>S�>�M�>S������=�	V>��>`W2?+�1?3�>�y�>�u6<��a�g�f�@���_�]f<�O�;��%=����|]=�O��١�=�>=3g>�=�>nt>��ؽ0�
=���>f�;?Y&?R��>%�z�B�&�5�U5����,>�'8=��6>��>�~ ?���>�M�>[�>�x�=�鸾u�ӾN�>H�&>.Y�= ��(�=vo>���>S`1?���>9���L����w�q�A>{A�>s&?�?W�R>�M>��x��B������mv3�D��y�O<#8=��_��� ��<��,�h^ν��=f-�>��>RÊ>ZC�>%7e>P�
>L1?�>�F-=�=��Z�����9e�����x��c>�b,����=�˽V�＜F�<ù=Hۼ/���Oƽ��(?C�@?���>->���=I�n���b���>|�>�m.?��
?M�>rk˾x꒿�s��۸ھYP?,�?��
?ɾn�pr=̽]� ���U�>9�>e3�=����y���]��~>�$�>�V>�=�����m��ɾ�U��[��=5_=zР?b�?�4��C�p��u���vI��?�~޼�Q�=V�H�{��з�zԢ�9��΃�ƍ�>L?��K? Y�����>8~'�k[��V!��sZ���>�}�>\$?t�>ѭ2��~쾯�#�p@�_%B���>�?���=B��>�_�>�;�<�?l?��P?�H�>�~'�Ƒ�>]=�>�?}�|��L�>l�c>Z?w��>���>c=���6=������������G��.&=+>���=En�=�(f<��#>��==v�W���<��=�@�<֩�<�O*>]��=��=��>G��>>;}>�!l=6Md��ļ��t>�t�u*���L�>ZU���,\�i�w=	".?�8	?���>�\�=�E��礚���"v�;���>��>��?*��΁e>
})��`�����=�g=N��x&�����޾|�f�@��=<\>���n>6@e?��]?��A?�j�">�0MY�C�G�_=�C>�>ř�>@5C=Ҳ�Ɇ�� >��6�1��Jj�;�矾37u�/?>�>"�P>8k�=k�P>�<Դ��f�O������'����>�~�>F�>���>�`">k���<X�,=?�̌�1�� �����o�;`9�>��>�]k��*?�['��k������I����>3q�?�X�?�=:?1`T��w����`>�(�>��=�����9�䝪��J�k>u5J>��������_��5>J��>Z��������ɾe^¼ip߿�ۇ�|j���P�ƃ�!������4it�"����/��_s��=V�$�/"۽~�%=��z=����ԪҾ=]���?%v�?i�ʾ�.��
��m���%���=�9ؽ�O���|�=f�D�)N-��(������g��[�c�>��Ѿ���D�l�e�Q���8�=��3?w@���L����h���V=�ۄ=џ��D���袿��j��=C?�^?yd��Ͼ �=������>7	?�L�>�Y��Ö��w>�Q7?��>y���o��3䨿�d=��I�?,��?��?�Ž��C�5������/>X>�>%�X?N
�==�O�~�=-�>)?�>��m������n��%?�]I?ܓ ��4>ACS>�>��ֽg�1�ǭ���E�l�"���C>�}�<����3��T⼰�=�.�>q">j���P���>#��PK�țB��A"��=�<�4?���e>�7l>oK	>�[)�T���������\�K?�W�?g�T?~�:?pM��<��yý1��==
�>2Z�>���=�L��~�>+"�>x���Ws�
C�o`?n��?���?�
[?2i�=;ӿ���J������T�=�/�=��>>��޽�Э=�:K=9����@�ź>Q��>�o>OFx>{T> �<>��.>������#�����MՒ�=B��
�S���fg�5�	��x� ��@�����b��������ؓ��dG�?��8>�l9���=t<�>�@?֭>��)>5�>�����<ɾ����x�R*��J�[���k�����]����������RH���ɾ6�Ծr�>��ȽB��>љ?ތ`>L�u=�4>���ץ=�ֿ����=�]>9��>��V>sO�>�
>�~���#>7��=�ݒ��q����'R����Ⱦ�G?�Tݾ��V�W ��H>���L��g>[�H?���>W�ɾ�2��������>�R[�|�=��>�G��=�>E�>+I��>�r	l����(>&��=A|�;1����N��ݗ>*��=���l� >{y��2�m?�?�:Q?*�����>�A�>Sk�>X�C��`�=�&?eP�>��?�\F?�M5?燼>��޼�d��g�8��ÿ�����U)>D��=1[�=Ҷ��,�U�̝ý n��fƘ�=�<��<�=�<Ґ�s�ؽQ��=�K�>��<?���>��>���d1�RDQ��.�%�>�����#�>�f�>o_
?���>��>fg>��Z<	���>�ב�>a�&>_�I�ǜo�Z���B�>��p>�15??;2?!�A��H��g=�2�=
ڤ>\?�z5?�:�>*�>O|�A�c������r��
>�#>a���>N�i�3���<�h��@����k>�>Cz >�X�>�"�>w >��B=�b�>�\4=���<���=�h��Y�u�5Y�M�=�=��?��k�	�Я�t�M��:�<�,$�M{�=
:>��T������96?$?�P�=9�=u�N��8���u�F�'?�x�>�?�=?�W�>G��U�x�ηj��!�Co�>Vb�?�G?�����4�>j�'�4�Z��?�{A><ؖ=p��=nI��TI� B>�l��>��J?��>dW��,"���$��0�ic�>��C>y�Z��E�?m?4A�t.��!E��MU�L�Ͼ��?����1=�����9���'���	�Q���>��!?��'?�l>�C>t�*�`B��mr{�!u?��R�>��>1?@?SC��	-����r����O=3,?Ƚ2?���7�>]@?�V�>p��?;
L?�%?l�Ҿ��#?t	>w�>�n�=)T�>��?�F�>Q�>�h�>2y�>U^=g�I��>��+F��B�m��I>0�[>�:=��<h\�=�^�=��!=�P}�'�t=V��=8����.>Ep�=��M�MЌ<�`�>��+?e7Ľ_�>�a����ν�|���=�kM>�7��]��c�ؽ�x>�.?�A
?��>1��;q=žZ�澻H�lߴ=���>Tx�>��w>�i>��+>���N�=���=���=�Z�{?��� |�BX�Ӓ����=�j�>�O>)��>� \?��{?�i_?�֡�V���L�.�@��B���Z�>�>+�?��j>"��DzH���y�D�K��\����m>�����i#=�?���p�>��>Nb>�%>��ˎ���{�vЙ�ƭ�6�j>���>rV�>>��>PU=��d),�A�I?V���Kh������_о�P�M�>�<>�8�Ɨ?V��/�}�b���8=�A��>��?B��?n,d?��C��0�Y�\>,YV>x�>�J/<�>�U	�ϔ��z�3>�N�=�}y�3�����;=]>�Ay>p�ɽ��ʾ*(侮QH���ȿ��V�Un�����缔���Ǿ)��E]V��ɽl ��]��)�1�����ڛ�=E��s��z�=p�>�ľ�)�?�ӹ?2ꐾ��V�"�=���:�z��S12>�s�<�2������Xͽ3z��!<���ZK��%����.vG��8��B�>�V�y6����t�V�+�7�-��*>#�.? ��2\��W��Q/=a�3>j��<�n�Ho����������P?��7?����쾖��}�>N�	?���>1+>o����\�~��>��.?�+?-�����*��z�ü���?Q�?��V?�]������k|׾����k	>� �>�8?ý�j�㲃<���>Q�d?*����%���y��� �/? ZM?��r�T�_>p|�> h�>��N=��׾�Y	��������9�>�w���n�=�Y���ׯ=|=9>�w>ߧE>�Z�(��>����zN���H����q�4+�<\�?���>Hh>��>52(�  ��K�����w�L?"��?y�S?Q'8?�����{�����z��=�Ϧ>���>��=p{��>M�>([辨\r�k��)�?R�?$��?�Z?;�m�P�ݿcզ�~*���ݾfbY>nY>� d>��:��|�=��2�S1���I��n�=�_�>���>.�>��>zP�>�#r>s����(�����/��Vt'�=��h'����	�7����B�b�A=��B�<�+��j,̽P]���� j�����<;I�=�ω>�;�>�a�>�jR>+�>W{�����䄾�� ���C�O?���ʾi�ݾ6\���������|����j佹�G�?3�>A���b��=�Ф>M�=�a�=?�m>�I4>?cy>(�x>l>�om>��a>��b>�<{>�>Vr >�ڠ>�g��%񕿶A3��5�-W�����P?L޾�t���؛�$�j�Y�r�r���<Y?�>��-����3��m��>�?�[M=��=dm޽��	>*o�>�E>�̾�DLg>z�����c��ܼ;)
�>B�s>58&��y��m袼�'�>�D�>�蘽��>���=%?=?�&�?]E?Ѻ���m>L Q>�!�>��=NX�=h�>\M�>�� ?XP?�?[��>�2�:�����x�=���4���W�Y�hĚ�c�����R >��=藮<��8����o��=��+�?�߼�r<�F>�)�>^Q@?fQ�>t%�>�e���=O�u+�;�ŽG��>8� =�EM>�u?�?b��>OU>�9�=�k��E��=U��>�O>�tV���G�m�c>3�?z�?���>(��>W����xC�)�?��8��}�>��?i)a?(?�>��j�IϾ,i��c������^����=D*�>�y?>�������:�TZ1�oUɾ�-ۼ')�>z��>A��>>�?�ώ>�R=K��>�l=>jO�=�=�?%��/�;�O�<�b��;�=E>o)/=��J="L(��"�!�
�4�=��[���K�K��� ?��?"�@>p��=8:������ؾֶ�>��>|�>�y�>\S�>��6�V�M�.���<>���>�Ӂ?�?0?~�M�1��=�?�t����#?�v�>�
�AV>� �=�X��܂���>pRE?���>�����<
��'�[&���5E>���=��>��?���?H��t����5W���v=�@�?��>>୽E�ڿ�d��ZX�����K�2=㎻>
�
?�^?�C�=��X>�mU��ē�X��VN��W��>�!>�p�>Q@�>���=/g�r�k��
6�\ ����>��0?}�<=�(�>i�?�y�>(k�?Q�C?�9?;j����>��=���>A��>e/�>���>�?G?
y>���=:)���V;�x>��8{輟���d�=��>`�e>XK˽�7<<	 >A�U>D�l���=Y�>�p�=J^�=�8�>�V;��>�q�>z?��<�y�=���<A G<D/>�Fk��c>[�>�S�� ���[>/�>�}?tx�>}1�Ĕ��Q��q�������>�c.?�>di��&>��о Dɾ<w]=�,�>��V=�3�������v\�&7?���a>��>��<�x�>��k?ߘC?�2U?��C�Js�N4�  �@$�<�`V>��i>�r�>���=V���{��_�x�@��	l�R>w�u���>w��<���>���>���E�i>�#V=��<,���7x=W���"�>�]�>f��>UU}>�t=�V�����e�G?�͟�x�������CȾOE��8�(>��2>����u?���i}�듦���9�K�>v��?�*�?�?`?�;�C����sR>�pn>܍>��\E���i�qv��#�0>�w�=��j�\��-�QSO>��{>��ٽ9-̾fAܾ�����k8�p�f���
���̾�޾����D�������#(����S��g����;��I�G��z>��о~���?��?oց�#��R�%��r(��8��\ >���qw��AU��%d{=������k�>����ʾ��o@1��2D�@�>������ZL���_�[�=��t>�~G?��Ƚ������
��6>��>%��>$
��3���a���i�)��7?�x+?�ξ�;߾ 7�;K��=�?���>E�>gC�&ξT)<jc+?y�?�=��Ě��r���"K<,�? �?��8?=j����k��]JQ�+��>�;>N�3?v��=N��C$�x�>!��>��>VdJ�������tӷ>�3?��ݽ�sX=���>�e>:��=�Tֽ��lF־��l�o�+>�ԧ��x��Ծ*|Ⱦ�!����>����L˾ӫ�+�>r��j"3�9{�X����%�s�|>��?2hӾ�Է���>i:�>�9¾���i�t�?�N�^�f?�a�?�r>?�G'?�ќ�Y�(��{M���>)��>�>���s5��T[>;��>���g9E�!���g�>���?�O�?��\?T1�����g��ў�|�Ͼ���k0׽�	�=G� ���D>��=JP�=e��P�(=S�>! n>6��>�b�>/>��>O����.�fЕ�ik���Z�Y�F���'�V�0���þ�Yf����G�I��n������½B�6�yA�k�*���a��&��J�=�"�> �>ٗ>�a�>��u>`g���ľ=4G�Cn��A��-����Lf0�+������:r������@��>(�����=T�>��V���`>�}�>.�;�z?>#��>� �=-�=�ޜ>LA>�u�=���>,�I�M�8>�G;q���i�h�ȭA���	��D��D.?��'���<'���J{��O�/���;}�T?h,�>�1G���ÿ������?��ƾ�!��J�N>��+>w��>
	�>bﯽ���Ӝ>�>�����V��-��>�/E��8:+��y�;�>��>.��>
�彐⛼ĽzE?R�F?��a?Ȇ=���>���=��>�!�=n�>�>c��>��?�4@?�W?;z>�=�䟼�">,�<��������l�k�J�I�/0�>�fU=v��V'=g��<����c��=�ŋ>r�߽����Rh���V�>�M6?�L-?�8�>�V���U��<m*�n�t=cf���Ta>�Ok>hm�>#�>���>��:=�C�=#>�.���i�L�>���<Ŷb�T�����%>��?-'?Z??3T�pđ�L�>(Z>Pu��⏚>�7�>���>u��>P7�=� �+;��յ�&7Y��J]�:���H�~�:""���<X�}�����ƽS/�C�u>�.�>���>�I�>�}�=�jY=���>`�+>��=q��=r@>�DR>6�=GI�<C��L4����=�&,�<3�=@��/����L=Z9�=������B?{v?�/�>�$�<������Ҿu�@����>��3?�U�>Ȉ�>�Q�>+���Y�u���*�2*E�E$�>C�?|�>�j½)�<����O���]|�>�-P>��>��������־�7>�=>��?6�?.N��df��/��=�����>9��=m�>�u�?.�t?8O�j-�������*���ֽ+1�>�N|�d�=v䳾
d���ƾ'�n��l4�>��$I�=�I�>Q�y?�߉>LO>�e3����^��8ҽ4�>wn�>[5�>wW>h˽_�߾��X�Ϣ��Ӓ>��d>+��>����֗?#9>G�>��?��?W�>5>O���H?1,^�c�Ǿ;Q����?j5h?�?!�$?�F,?"B>�����"�
�7�V�;�� <O
żMq>��6>3<g���">��a=S���C� ���V���>	�M��|$>��i=@r�=y��=��>ǁ&?h�:>C&,�'�r=-����=^���a�>t�>�y���ߛ>��>� �>3$A?%G.?�Xq>�ؾwD����:>�d>?� ?�)?>���<9JL���u���պ� ���^׾�꯾��C�;��_�3�Ԝ/=9�D=��I�^Tl>r+}?"z?j;W?�ό���+t��� �'ˌ��?�>�`�>�2`>�VS>���F&&��+G��	�[��t�+=��d�n��<�����'
>���=@���2=ߙz����� ��;�}�9v�s���=�S�>9��>��=>�-�<��Ⱦ�v�MPE?��߾]x-��������U<d��<��_=����#A%?�^�=aK��%��,2��4�>ԁ�?S�?�?���x8��Ǫ	>�>��=�J=�.X���U<`��<�R>'C���4��ٮ�����=�W,=��>=�Z�c⮾�-���=��ȿ#SF�������I��������4���*l�P�1�s�̾�F��j��eN��J�F�y�o��/���)Ӿy�;9�?���? Ô���m�v1N��B���e����>D_þM�u�N��	>�����l3�L������8�ge��;s����>a���)W����C��$�dc�;4��=�"?�6�l�b�0�]��������L��\�$���s��X����ؾ^V?0�?����,!��w�p������>���>���>j#������>�>.�C?�?��A�r�}�����s��Nܸ?���?�'?�w�����1��/��ߗ
?˔�>?'?�nҾA{�C��>���>��=�6��?�8��&���`F�Yk?R��?DM���">�o�>k�}>�3������(����=Pj�<=@>ME<=�w<W%��ߙ=�6>��/>EN0>��@�V���۲>쵾2�?��-��վ�����p���?C���Z$�=��k>q�f>���]}�����M���dO?�n�?�cL?M?w���ﺰ�ݙ��=���=1�=>�\<s�=M?V�>C��0A������"?���?)��?AlK?��r���ؿ��������s����ļʆ<�]�>�p<��M>t��<���;�W0<���;G%>EB�>�ܞ>���=�c>�x�>������)��ڍ�*����v�����K�Ǿ�M{�#����p�,��1i�_��<������¾,��6PV��X�w5]>��>�U�>�;>���=C"9>
��� ���Ľ�b����B��Ծ>w����U۾�C(��*Ҿ��ؾ�`�Q\��ֲ>���>!�>,+�>ՙY>��{>��Y>6a�=�3�>������=Ȇq>ㄧ>�>%,>Ǥ>qs�>7��<�������ꉿ�
�DU'>9_��3?0n޾�$���y���/��0K�-F����X����c�a�ꆿW�>�h>�=�<�����4=��;>iq���>�{D>�AϾ<����X>lթ>и5>�pc��85��ɾ[*Ž�7?��Ⱦlɯ>�?G�?�??��S?R�:y?�L?y��>܉=_��>r��>�b�>KlH?b?�7?�'J?�>��;�My��Cf�=�(��^H<G����i�=F�>�g���=�<>t�<�"�#���1����0�� <��=n?�t|?/� ?;?8d��>N�l�P�]о�F(>��>��6?+d�>g"?��8?��?q#�>��!>ޚ[�d�c��_�>�E�=q�I��a:���=k�w>M.%��.?�
�>F�>K@p��H�|�R�U�>��>j(?" �>l�>t1�<AG�֑տZ�#�(i����*qu��D��R��"�:�yZ���)�E��fA���n=ݑ�>,>��)=]C<>B|J>�X�>wSU>�o?=%�=���=��U*�\{�=��Ե�r�ϼ�o=���<RC=��2ԼDw���S���P"��k?��"?{����6=D��|�"�YR�΋�>%�?Q��>?]>�vľ :��`�K#=~�?`Xa?Xy�>�k���<�Q�E���.X>V��>5�o>�|u��j���J��S�=��>t��>�(�>����O�y�m���66_>5�=������?/}n?���3����c�T���ؾ��#�v 	>䤽�V貾�6
�ά@�|�þ����y��M�Y=��>�B�?u��<���<!w
�Ӿ��5����+��б�X�\>���>}��>}��=���)�ھU�ʾi�8��
����nc>�Y�>-|�>�f�>V^?G-?N��>-d@����>)�&>�>]̶>�?��?0��>�M >\_z>FP3>��=����{pF�c1���������=��=S>�`>!f�=e��C+�!b�=�x�=���<" �=��=�ߡ=6��=Ԡ2=��?��;?��мx�����7��}~=)3{<T��=o`�=[˾�+��e�=��>�N�>�^>-��=������n��Se=9�O?7.4?�?�+;��>�B�un���窼�+�>T�	>�J�+�P���&�}4>�m�>+R7>8a>��?�:S?)�%?��*�9�+�>�j�%I�Zƽ�E <��>��>��>������/�Jta���S�?n3�M��/@%�x�>�) >N>�F6>�RD=9)=0�����ɽ_j�K�<�F�����>��?w�?*ab>t�=��¾u��ۨI?S�����&���wʾ[�'��&>?&>���?lR���x�x���9��]�>���?���?T�c?6�/�����E>TGP>lS%>_W���0��D�����d:>�1�=������s[���^>�<w>W(ӽsɾػ�uT�%#ӿHyv��ؠ��e�Omh�^(����^�?>�I��d������k�Z=1��D��%1>�)��&����m�B爾�;�?#�s?�[��E���*��mk���ȶ��/@>�־�㋾y���v����!u��nU��о���þ�o �Τ����a=�^����0섿���Ws�<���="17?��okϾ�`�,s�=J�=#�Y�~��F��-y����$�={(?^�)?�ﾄ��tօ����>ShP?"��>�)�=G��b�e�LE	>�?oU ?ǺU�����U���� �W��?K�?��?���j�:����� =h=?{�>O?{�¾`�3�����P?�q?(C�>����N���>���?d
<?u����>=��>���>I�ő޾k��Yؽ�6�>T�7>Lۆ�����u�c�ڽ�ݯ����>�[�>f��Y�9����>�S�.�L�Q�F����4�:i<xj?�"��>�g>��>�'�U猿rd��]��2M?��?@Q?^]5?�����羊������=W�>�>d�=a] �i4�>���>��[�s�9{�:?{�?��?�W?�k���ۿ����	��>��5��=��6=|y>i�u��7�=2��=Y�}�l㼰�>�
�>b�>H�>��>�5�>���>.��(�*��5���ܤ��v9��;����ԥ��yh�7G�� ��������ۧ>�Ӽҵ$��
s����R�"=�`�,�.>k�?��>]�>�f�=�G?(��@�}k>�`������1 ���
�����#���P"s��0�;���	��2�>qy�=�m�����>)�@����=DJ�>��#>��>�ظ=ugL>Қw>[�/>�>�U>�>�d�>�ɾ>��>B����J`��]��Qt�\���Qv?k�3=+.:��XC���~h��	B��rg0?��=�b�zM��OG����>�����/߾*�Ͻj����>Xd�>{S>�Cs����B�L���r�t��Zd=>%A�=��H:��7�$�6J.>yš>-N�
��>\��>�΍>��?��J?�v@�L��>��>C�?nKL<TM�=03c>m�<k?�??��+?�??eմ=4�m��J�=�k>�0M=�/��^�(&ν�)> KM�xxg����w�N��M>��Լ�F>m�ȼ�н�,<D�>��F?��?�/?sN�;��N��k�R�Ⱦ��=���=���>�X?b*?�?�7?	�>�y;=��¾�Tݾ��><[>سM��U8��ھ��>��>6�`?�2�>	����+�����=R>E�
>��>
?�A�>�4�>�R�����I�Qv����A��<9,7���=H��Q��ƈ=�ˇ�ͧ�ƒ>���>�޿>[��>|��>)�>���>�>�Z>��;��=�$>kE��hx$���6�����v�Ի̽�0�<�gf��$^�C������Ȕ�&^��pܽ���>G5?*�Ͻ{Tӽ_�L<!L��j���D��>�>V'�>C��>�q9>��ʾ3/_���@���C�٨?��i?Ar�>V]齃s<Nߴ��1���>���>vb>	�)��� �<�m�/��=T&?>S�>��>��AC��4�OV�����>�=$z��$Y�?4�y?)6���z�����`a���X'�=˒�<�7� 㓾��۾c&5�J��'�����}�7�F>�E�>4��?����;l@>��h#������\��|<�4��=��?��>N�=غ�l���L}	��Z��<�T��;��=M�>�`?i�d?�z?�S�>� ?��T6�>?b�>=�?8�?S�O?��1?��?��>_��>�(^>���=�^ɽ����s��c���$����2�>��d>�%B>LGZ>���=��㼚���0�c�v;qa*�Q�E�|:?>-Ր>`S�>��5?Z���� ��Xd=�ʾ�e�Ұ>�F8>��������9��7�;XO>}k�>
��>Q��!}��. ����h�=�9?�P?��?�V��T2o>��0�M:�FV�>	,">D�	�O=������nо�\6>��>{!>cڙ���o>�y?�[?YD?�h�<�$:�ӂO���P�U_R���^=���>U��>�W>=!Q��4��x�`�hT���3�6nG��C��+�=jw$>ݣ$>w�>���<�ŋ����o1ýr�I�>uyL>��>��>1!4?W��>^\=�L��܄��I?>]��dQ������;�'��&>��;>�Y��7�?�	��*}�r���ʧ=��`�>��?Ve�?�c?��@�$��?^>HV>��>\�<�MA�k��̂��4>X��=Τz������J^;G�_>R{>_BĽ��˾��DI���ƿYe��&��o�`|(�9��M�����Þ>��;��.����#��3ܾz3 ���;:UW���F�G�}�&;�?��?�c˽�"����6����5��W��>^���b�����������k�뜾�&��Y龓A ���S�.����>F�������|�K�?�<��=�Sg>>7?,Ҿ� ��/W��$���| �&G�=�<��������|��9/?�?���p������Jǆ>g��>n2?��>+2ƾ����5}>f�)?��5?a��=�瘿���U�,>ㆫ?V��?��=?����(���(�N��>��)?���>f�>��־�Ͼd����3?��!?�z�>��X�a��7����-?$\)? �����s>�<?��>��=���Y��F����=�;�>�nJ��f����~ƾ�l> u�>p>E[D��0d����>H��1�M���F�b���R�:�C<�?�󾑵>�k>3�>�r&��f���h��(h��nN?��?A�Q?b�6?�5�zT꾞��&,�=g��>}w�>5ڱ=(��-��># �>w_�k�q����&d?���?��?��Y?\ l�޿~M���r��cv���a�:v'=a��>I�潌��=ӈD>�I:=����e>���>ʙ�>���>��=��>�N�>�#���'�•��֐��Vb���"�$�ɾ����'�Q�u�z�Ⱦ������k3>*W�=�I=M�6�P"�S�-=�_P��]k>��>s�>3�>,�>F�;>��Z��������q������z	�b���۾z�o��ӿ��"a�r���v�����;��>�ؿ=&�>$��>�>�K�=Hi�>(�ý�>��@>{W>���=��M��`l>謥>N'm>��9>�ϵ>��=0���"&|�=�Ͼ�x��L[̾I�W?Y��Y�����G���ƾ{D���>�	�>�A�'�J�pO���9n�N
�>y<Vb־S�&����T�> �>�b�>9¼=@z>R���}���t�=��b>�tf>hM:�g�1��=?e�=��>m����>��?�/?<�?��;?N����R?�W%>>�>o�=;�=��>����fC�>*%?H�Q?-o?V��=K4����=��b>�DW��}�=��O�@�P�6P+>rֻ�h=�xU<O�>��ٽ?�Ƚ`�нЬ��>h=ub>�s�>�>:?�s�>��>����BF�����7��W��=��O�:�>���>�q?ڦ>w�>L>>��<e���Ҡ��v�>���=�E� :M���-��>\K>Q�_?ma?$Hμ&�߾������=�c>��?  ??�4>=qh���7����`��O5��U��;a�U;���w	>Wo ��0i=���>������U2�<z�> ��>7�>���>W��>- �>g �>�2�>��<�I�=���=�z5�BR��N�i��r�<";��U�`-�8l�<��r�f��"�.�Mp���o�v̒��~�>�`"?X�"=dA�qG�ѾSp����q>"�>@�>PR ?5�>��Q�6�i�t r��/Y���H?e?��>;�_�u�Q=���=W)Ľ�py><`>�ȡ>����|���Z�=�C�>
2�>���>���=0�C���]�����\V�>�2=r�����?��h?����+�rݾ&�Z��Ԟ��=�1=��ὤ�l�K|��.��&;�X۾� ��gW>;�>��?	8�&}�=�x������������Ž�c>܎?���>m��B{���Y���0žD�;�m����l�=�8�=fL�>��?`?86x?�-?��?��P����>��O=~�>.]�>}��> �>���>]Os>���>[� >nՋ���#�������6�;�<�>�� >��Y;3l5>�$�=EU:��ٽ�о=`X>�<�;�<F�<H�>�1t>��?�v0?����e�����J������v�AN�>	���wB�͑��
o�5�>>v�)=�^?Ϳ�>�v3���	�l:��.���ἛRD?��)?3+E?��>�==>��-�Ģ˾<E<>NM�>y������I��$��ȔY=-*�>�}�>��q=%a>3?�He?�fY?֬A�� G��iE���l��D��C5�=D��>^�?ͮ�>�\m�����I��$M��e�я/��Y��t�=��=�qT>�C{>��*�y�`=�t�;�o��v`������p=C?O�>�.?i�I>o�7�o%�����J?YF�����j���+IѾ8����>�/=>��iL?����|��S��#5=�]\�>���?���?�
c?rD����]>�5W>��>I�<5�=��u��^��W�6>{��=�M~�n.����<;�n`>F�z>�)ս��˾p��~?�k5¿��I��Ž�����C/��_��_���%%���(�iF>�b���?�Ǿ�N�\�<)���z/�C�I��ɽ]��?��?��H��D��8w�ܺ�	C�@Zu>Sk��7��c����h~��j ��h���=�Pu!��tm�xC�q��>��X������|���'�)QV�{�8>M^0?��žc"��?�NR=�>.�<n��s���]ʚ�ak�$�U?�R9?�R꾼}��ڗ߽�&>e�?b>�>��)>@l�����P��>x�3?u�-?�μn�������Q�G��?��?NT:?7'ν��N��  ������?E�>�[�>qX��	������6�>&�0?[�>�,�<4�������>�S,?�cu���> ?<mv>�"^�S�¾4���q����=�� >����.9��j������Ds�=���>Z�>e�3�A��;�>��¾Ӕ=��+G�w��0�'�Tz�<4��>r�߾ɋ>>�z>~(>� ��᏿B
���3���Q?���?�AM?�(?�wվ*���:S��mL�=(o;>(�>���;L��ux�>�^�>�,����t�$o?ș�?�?c�E?D/޿�&���]��c���f�>�>|X>������7>���q�� ��=��U>�>9H?��?
�w>�ݚ>BR>�Έ�X0�%q��Z��0C��X
�!rپ)\(�(�վ��־Qe���KW��˱=v�=�*�<�vC��|2;D��������,>7�?F�>3i�>*�>-J>����;��r�B��dƾ����<�47�)���������$k�2[��9ͽ����,?/@==�[>�W�>�@�;��=yP�>O��<��=�k�=_�>_E>m%/>��=s��=�x>>>)�=�?�>�{%>����O+��qD�0d�����IvY?�5c��+��坾������<����D�>��i>�6��7vez�*��>�^+������Wм��>�{?x:|�8�Ҿ{��=�N����=�>�e���=�p�>��,�}|�;�<�/�>�#۾E��>�(?�?�m?�[?]8�9�?��?��?8+=n`���N}>qj�>8��>*?+?e�s?>YN?)d�=�P�
t�٭0<Xő�J>^�]5��Y.�=�Ԇ�xf<g�*>
�>#}=w>=:Oz�O~�=��=�Et�z2>h��>0�>?&?i�?{���s���$�����!�>6?�>ݻ�>U*�>H1�>�)-?��>�釽���<�ƛ���㾈��>� ���i�v�R���=���>��>�mZ?
� ?C�O���^�g)�����6=���>�?uj>���>�i�<�p�7���F���	�0��=z�l�jbU>��#[�<,^ҽ���I=�	�<s�>s��>A ?���>M�?F��>�V�>$ek>���@�e�7��
d���G��꼼i��o��=���=��X=�H������U���4>��>�J)=�B�<c�?՛?��=�=֔�S)�։��{�X>v5�>�Z?�>�H�=�4�|S�:<'�!"#���?��O?��>o'.��3^=T>�=\��>b�>�*q>:4>52<��U��gپ�����z>��?��>�qX�`UC���b��p���8>�%�<�����ϔ?= [?���j����~%�
K@�C8����=s$��]��Ï��9^���8��/��g-��.�~=3O�>l��?��z���
=1_��3�����������=��=:��>@6>��-�����~��0�Ⱦ%�T��}H<HX�>���=u>1<<?jV`?�.�?��'?D�S?v�ɾP?���=�Q�>6��>[��>ހ?Gu�>�XK<���>�a�>�j>Б��$:t�ߋ����+��Yt=�V^>s5�>�P
��	>��?��|A��E ���=�V>�?=�X>v�9=�� >�1�=a�?��E?�f
���!���۾�؇�J�>x,=xF����=)+��(��RؽR��=�?�>��>�Ԃ>&�6�}?��e�=�O>g5?��*?ۚ�>_�<�ĖO=����)��o>��9>%G�=���&�������ݷ�x�>ח�>�=�Tr>JBr?��|?dtD?2����V��AD�]h������S\>��H>�z�>�=#X��d���>{�[���$��1#���Y���?<�F>�Va>��>��=�F�������Z��������=����0`�>�
!?�b"?0}��Fx����3���2E?����"�� ����ZϾ��WH
>�">@��7�?=ͽPl������OD�6˶>� �?P�?�_Z?~S��`�#f>ꍈ>rS>��=�ys����� ����:O>�o>/d����k�j�}�q>.F�>������������T���Ļ�T\��
�,�K�$�i��g꾢�H>�ޱ>�7���%��Mt޾�a��Gد��<S��*)��g�܆��$�?�.	�?���?6y>�#= �$��
���N��i>!�C=�U���0���̾Ơ��9㭾��ʾ�4�K��`N�4o1�*��> ˇ�{����m��o���	=��
>��.?��έ���W꾟� >�8�>�y������d{���g����<	F+?��"??���:�%���z�>raA?ܙ�>oE�>V&˾��K�n+a>Χ8?��?���<|����u��R��¹?��?�<%?����u.�Z�;����<�Bo?o>�>Ġ�>B�0[�0t6=�2?l4�?��)>sF9���˾�G?#��?&�!���Q>`9?E>��L���$����⮾��x>�Yh>Ϲ;�UG��࿾��?P==�>ۥm>v�G��d����>�S�.�L�Q�F����4�:i<xj?�"��>�g>��>�'�U猿rd��]��2M?��?@Q?^]5?�����羊������=W�>�>d�=a] �i4�>���>��[�s�9{�:?{�?��?�W?�k���ۿ����	��>��5��=��6=|y>i�u��7�=2��=Y�}�l㼰�>�
�>b�>H�>��>�5�>���>.��(�*��5���ܤ��v9��;����ԥ��yh�7G�� ��������ۧ>�Ӽҵ$��
s����R�"=�`�,�.>k�?��>]�>�f�=�G?(��@�}k>�`������1 ���
�����#���P"s��0�;���	��2�>qy�=�m�����>)�@����=DJ�>��#>��>�ظ=ugL>Қw>[�/>�>�U>�>�d�>�ɾ>��>B����J`��]��Qt�\���Qv?k�3=+.:��XC���~h��	B��rg0?��=�b�zM��OG����>�����/߾*�Ͻj����>Xd�>{S>�Cs����B�L���r�t��Zd=>%A�=��H:��7�$�6J.>yš>-N�
��>\��>�΍>��?��J?�v@�L��>��>C�?nKL<TM�=03c>m�<k?�??��+?�??eմ=4�m��J�=�k>�0M=�/��^�(&ν�)> KM�xxg����w�N��M>��Լ�F>m�ȼ�н�,<D�>��F?��?�/?sN�;��N��k�R�Ⱦ��=���=���>�X?b*?�?�7?	�>�y;=��¾�Tݾ��><[>سM��U8��ھ��>��>6�`?�2�>	����+�����=R>E�
>��>
?�A�>�4�>�R�����I�Qv����A��<9,7���=H��Q��ƈ=�ˇ�ͧ�ƒ>���>�޿>[��>|��>)�>���>�>�Z>��;��=�$>kE��hx$���6�����v�Ի̽�0�<�gf��$^�C������Ȕ�&^��pܽ���>G5?*�Ͻ{Tӽ_�L<!L��j���D��>�>V'�>C��>�q9>��ʾ3/_���@���C�٨?��i?Ar�>V]齃s<Nߴ��1���>���>vb>	�)��� �<�m�/��=T&?>S�>��>��AC��4�OV�����>�=$z��$Y�?4�y?)6���z�����`a���X'�=˒�<�7� 㓾��۾c&5�J��'�����}�7�F>�E�>4��?����;l@>��h#������\��|<�4��=��?��>N�=غ�l���L}	��Z��<�T��;��=M�>�`?i�d?�z?�S�>� ?��T6�>?b�>=�?8�?S�O?��1?��?��>_��>�(^>���=�^ɽ����s��c���$����2�>��d>�%B>LGZ>���=��㼚���0�c�v;qa*�Q�E�|:?>-Ր>`S�>��5?Z���� ��Xd=�ʾ�e�Ұ>�F8>��������9��7�;XO>}k�>
��>Q��!}��. ����h�=�9?�P?��?�V��T2o>��0�M:�FV�>	,">D�	�O=������nо�\6>��>{!>cڙ���o>�y?�[?YD?�h�<�$:�ӂO���P�U_R���^=���>U��>�W>=!Q��4��x�`�hT���3�6nG��C��+�=jw$>ݣ$>w�>���<�ŋ����o1ýr�I�>uyL>��>��>1!4?W��>^\=�L��܄��I?>]��dQ������;�'��&>��;>�Y��7�?�	��*}�r���ʧ=��`�>��?Ve�?�c?��@�$��?^>HV>��>\�<�MA�k��̂��4>X��=Τz������J^;G�_>R{>_BĽ��˾��DI���ƿYe��&��o�`|(�9��M�����Þ>��;��.����#��3ܾz3 ���;:UW���F�G�}�&;�?��?�c˽�"����6����5��W��>^���b�����������k�뜾�&��Y龓A ���S�.����>F�������|�K�?�<��=�Sg>>7?,Ҿ� ��/W��$���| �&G�=�<��������|��9/?�?���p������Jǆ>g��>n2?��>+2ƾ����5}>f�)?��5?a��=�瘿���U�,>ㆫ?V��?��=?����(���(�N��>��)?���>f�>��־�Ͼd����3?��!?�z�>��X�a��7����-?$\)? �����s>�<?��>��=���Y��F����=�;�>�nJ��f����~ƾ�l> u�>p>E[D��0d����>i���G��NC�qZ�W�*����<���>
��g;>�+o>m�->�5'�֟����2=�b�<?^~�?��W?��)?�Ѿ�=վC!��^��="�>�s�>""r=�A��Ȥ>���># ܾ��n�Y���?j7�?��?}�H?m�n���͗���1����e̻�:B��2�=�����Y<A��=�p���C7�<4Sc>l>>\2,>���=>�+<=�0��"	&�V4��Fߍ�-9���5)�m[����Qڄ�CX��6̾�

�ͦ��S罕T���S�����JN���~��N>T�>�B�>ެ�>�Ig>�r�>-/��:m�
J������$˿�@�9�pb��R���-V�.�.���T����l��^��jX�>�%<-�=���>�s��І=�ޜ>�\
�"�B>�Ƽ=��>
�g>�l�=9�~>$S>u�>�s;>�י>/5��G��PLM��/���:�R�����_?c���d2 �g�ݽ�#U��/��R[e>���>J�I>�,�G��tb���)�>��#f/����=Ы�=��=��>��!=$%6q�ܽM{�3 N���nit>cn�==� �r嶾��7�U�W��,�>A����=���>��+?�Vw?�M0?1�/�՜>���>���>�|=c��2���߼���>cP$?2�?��?*�o=�썾)n�=.�K=�D���I,=�ί��J���1�:;U����;\H�w\���]|;V =(�<=���Q{������>'a?745?{K??Ἵp��bZ�ڼ ���w>a�HAT>��>|�=?y؝>��+?�(?m�><���0�%��	?�ޤ=�Di��1�c纾!�d��v�M*�?��>���>�8&<�f9�V2�D҂�d7�>tE4?��?3$��g
�I7�o�ۿƈ�u+��'��c2L�k$������a��'�T>ƾ�nY��ӽ�w�=�Ji>��=��=��/>6>�f ?#+>�ܸ=�*��^���?)=�����=߆Ҽk	�=�Yz����>&��<(�S�)�O=m!���%0������.J�e?��(?�2$�lX��'����@��lV	?��>L��>�O�>ax�=��{�h�2_ľXS��_�4?��/?u?҉��穻mL��6�=�Qg>-X+?��>�:� b��� o�>�	��
�=>�K?"?�M2�XP{��G��Ԯ�)��>�~*=��(��?�dj?�����[��P�UV@���վTL`�W>���Ⱦ��(�<�;��+��v����0�> ܝ>��?��y=��>�@W�렿�퉿	S�S쁾iaս�T�>pH���#S��_����־�]���[p�t��=��>��?��?�Fu?��>'OF?r˷��#�>n��>��>��	?�?�?dQR>�_f>#_�>	5h>�[>R�kQz��$�<�1߼�JJ=|@�>�h>��=�#`=Q��=�(�<$����;'�޼�=�g�=�!={�H>�T�=�{
?��?����p�s]��T����	�h��>��>�Q��8���X�S�+�[>���>��.?�>��=�c=:��D��b9�s�G?�M?I��>����P~>��,����<E6ͽ��>$ȶ={.�J���E���;G.6>g�>Gy�>�=���?�`h?UX?8�>�����%��d����Q���S{=ol?4cp>���+�-�y��5G�ޙt�\�~=�����>��b='�=���>m�i��_�>ޙ/�G�>����3Y>�?�o?�E?���>�z�>KKv���ྡ�I?�y����������Ҿ\�$�pi><�E>y:���:?�#�	�z��ӣ���>����>���? ��?�:a?��<����0Y>E�N>�>{*<8�.�?f޼S��0>pw�=�0}�ʙ���<< �p>
�|>&�Ὦ�Ͼ%�߾!�F���ÿA�V��q_���9�5���iC�E>��W���C���	��I�ھ��.�E���I+�ց9;d�h���ھE��G^���%�?,z?�I��=��K��x��ƹ�'��>!&z������/��!8���������Ũ�F�ξ}����þ�N�s��>T���g��Z�d�Y?�r,�=�4�>��1?uU��F�2B羟qb��1>_�'>�$5��Ƈ��ذ�����:?�@?�о��ɾ��^�`�=�H�>aί>��<� x�->ɼ>��=�3�?�� ?��Ž����{����������?��?��D?_As�A�0�����tx�0�>�@?-��>aH���Vy�H�=��?��?�>��0�37���D$�~##?>v?@w����>\ ?�{>c���y����p�H���-$����>'>ܱ�<;���C��w8R>��>KpF>F�k�{���l�>�˾��9��`>�$j��K�܀F=q��><��T.Y>#�x>�Hz>`�4�1U������:�u�R�8?j6�?��Z?6?����u`���U<)|�=%�c>mr}>Y�����d��>���>��ʁ���#��I"?�F�?3Q�?˘,?�v��ۿ����4���0;e1>�$�����=Q� �R�<=:�j>cK.�>��(:[<;�`>��>�xc>�z/>�7Y=.I�="����"�a�c����'6��(�l��`���j���5c���"�sNξ�ľ���vn���s�/�D���ǽ�����VR>��?�>�?;�d>�>�&�eٸ�?���Ǚ��F��w ���*�#��[����M~��͔��Ժ�T�E�:G;�� ?!Ͳ=)�g=?�hc<s�p=oB?bŇ=�3&�	�>��&>DG�>��>۞>�/*>��=�6>�%�>��]�P��#%P����R���8�4s`?�|��� �n�����B��]��Q@�>& ;?R�>�6�lf�̰��+M�>-:������p�ޢu�`*�>?��>�}>ռ��>���~����<E�=�$>���=9_��D�r�s/>|b	?`P����I����><r�>�?$��>@�>aV=��>�p�>�V�><�R>�9=���>�	?�?�?���=�T�v��=��=Ѧ�oB=�m=Y�X��L6��^�L�Ի��l=􍽽�`��,���YD�m�<���< >p$�>��G?+~#?��@? �;��V���
�>7���?�2ʽus�>���>H�?�'?��?g�>.�>ꦂ��3��q��>�;�=�g�! ���ˑ�;U��=D��?�FE?����Q�|��|<`}�>���>�z=?� �>+I�=g|�������m�;�t&ӽ��~������Ǿ�]p�����]�X�����`�=:��=/<�>hs>m\>>�;y;�>�3�=3�q�=�u@;� #>��Ƽ=�6<�%м��7�fAI=�d�=�<k�z=�<�ݳ<���䡋=�/�`�>E"?�z��2",�{���B���
Ձ��L�>�F$?�>��>�>�>��ƾ�8E�� ����ü��"?��b?	�>3����=�м����)�>� �>���=,ӽt;�� e�U�7���>G?gs�>�dm��d�<1c���-BM����<)�ӽu�?DV?wy�)�x�%��2e�[��~.�=���9ms��)����J�LO��[&����2�;^1=>�(�>��?�je=��z<W�F�4����L���о�n���4�=rۛ>|佋4��Ǿ�_,��D��Q��喽dF�=�!>흞>�W�>V?ОW?Qw?�?NY���X�>Q�>$Ǵ>U�>��?]g"?���>���>��>�U�=tC�=Cн�ɑ�b�MV�=�Q�=к	>�uJ>���2��<��=�;q=�e	�!_ ��>� �=�G�=�	�=c�>��Q>�g�>�*6?#�W�}E �Al����߽�BV=+�>2��>ex�a���� t��r�>��>� ?/	?��>�+��-��v�ھ$}��E��>ME?>,�>�TY>��&>p'��oѾ��>-�,?�,�=ˢ��A��q�佫��'�F>P��>
��=��=��?>��?� ?��>�CE��{�<܄�����>���<>�=��=OH*�qmi� c����R���(��h�=�B����=«=Q�H>R��>��<�^�=��.=���;�T����<��@���?�?é-?��>9�<����{��NIH?B�����hD��{pվ�TD�tR>��>>�F��y ?(��ˀz�R��o>��|�>G��?��?^�d?!�D��4���[>1R>��>��c<A�8���0�{��T�4><C�=��s�����q
<��[>i�w>F&˽z�ȾxC�Rna�����%�h���O�ρ��1��vߓ�Ǿ��P���z��V|�Sܟ�@�S�|f��:[���ڽ+\�g���s���Q��G�?Ԋ�?Б��-_���N�)Yﾓþ֚�>�숾(���������q������젙�56����A�� ��W�>�Z�eg{�BRw�� �]L>6k�>>1T?bbk����q��A8���D>��=  -����������K4?��,?����2�?�ɾ>�L�>��>��=�伾+�/����>��Y?ި)?7=a����ů�T�=�~�?�%�?�C*?�:�S.�M���U�Q� ?֖?��?�*���9���>{�<?��?��K>OV�y��@�ݾ�2?��l?�y���3�>�"?�ƽ>�2�����S{Ҽ4�����=���>�@޼�W�=��-����F�ٺ�>���>�%�/M���{�>0��n[N�(�H������w`�<j-?w~���>cj>�:>�-(�-挿t���ʯ�RL?�-�?�S?��7?�`�����Ŷ��:��=�k�>ҫ>���=!��$�>,��>�t羉s��T�3�?�
�?Y5�?o�Y?�om�U�οt���Lݛ��q��K�i>��=>o�A>�D-��$>6�?=mw��i�=�<A��>}�>�P�>�i�>	�>/W>����(������㋿8�6���	�[�����2g�r���{�����i�>M3��-�=�"<�?8��1�*���_����>=�?u��>En�>�v�>�{�>(���5����:�M��ؘ�t27�>���e�����}e#���I���L�]��P� �J�?9�>m{>��?�����gE?�@>��2>���>��<ko<>�|>߶�>��=>B�>@aĻ�u�>�&��5v����M�ӻ��R��;uN?t����M��3����7�iԋ��%�w3(?�M<x3�%5���垿t&�>��������oI<�',>���>7#�>u�>v���$�=Hn�=�j�%6a=W2�>�h�;j4<�w�*����>���>�~�����=��>�?uv?���>S/�<���>\o�>���>@�>w��=���>��5>2	�>f�#?]��>9J�>(�:>V��&��=�8>0�G����.�-��ո��p���Ai��/ԽڟC�p�<��>D=�$:>���ß��T���d�>UY?�*1?�u�>g{�=D#G��+��X���h�>�g>H>6I'?��6?�?E�>[�>�#�>�䯺^�V����>Z^>:�=��aR�mȾ�	L>d�[>٘t?Sf�>t�r��-׾��P�)�=l�>�A?=H3?�?~��>�$�=!����鿭��'4�l�,�����/	>����O��� T>�ȷ�/3��4��3:>��>���>���>w�>C�2>�#�>n�>�}�T�^��%c���J��gE�ХQ<p�
�_"�;]�c=v� ���*=�7��&�����]�*�����/.���?gS?y-�<�����'��V=��f	˾,��>�?%?�z�>��==Jd���7=����y���Xz?�#s?�!?�JN��R>�߽6X�IM�>�?�]�>�p��w�b��d�����?$�-?!�	>l�z��+�� U��������>�\m=���
O�?9�I?�tþ�m�-����_�8���<<���$"7��,��B�+�(�{����n�񉶾��>�m�>��?�I��A��r|B������$������*�<:]����>(�#>E뮽Z�2�vP�l����^��6�����>>:�=>W�V>;}�>�e�?@i?�>��:�y!�%'?��??�(?�Է<��e>�)?J�?�˒>N��>G�9>�""��)l�ݳ��K�=�L�=���&�=�=�� >��Y;m�>	qW>����DL��L<���<(�=`�N�r*����:���>��@?���=�Sm��c�>�:Y��d�1f|>l� ?�ی������G>�i�>��F>�w ?��?'9?��l>���}��2�`�ٵ>�6a?���>%�b=��?�]	���W�\!>	��>M�
�9샾X-y��>޾����-V�>dЛ>Ɩ >L�W>�:z?7Hi?}�?X>"Z�?�i�B�c��!�|	�=�ʨ>��?�=7���m�m_b��Y[�v8��v�=�k��@[K>�2�=�so>��>�J�=�泽w���k>�(�=�q�=`��=:��>�?�jA?�z�>t�>�L��/#��xM?�Ŧ�\R�55��XP̾�A����6>b�\>�;2����>�Nѽeyn����h[8�O��>[��?5��?�R?R�b��~Խ�$>�	W>-(�==��<LT1���Y�����>9Ŭ<�>�ӧ��}=�=f>��H>'�z�+�*���?(����� 3�ՠr�"6*��1�'���]��� ֻy����I���m���݅�>}/�JE�����2Ap� s�����ޜ�X�?�y?�*������97�1��$�ھǸ�>�%;�o���$p�lu���a1�~Ѿ��!�\��N�u��V�>�؃�� ���Ae��W���n>���>��6?��վ�ؾ�1���aؽ���=��=��̾Y/�������L�i�1?�4?����4!����ҽ顀=�?�L�>�a�=U���������=�q??�J5?D�e��듿q昿� ��u�?ċ�?�:?��y��Ɵ	��(��u?
�??n�>��ӝѾ�g*�ԧ�>�w?g��>�`d�������V��C�=��y?�ݾԽ?3]+?v�^>��D����`0�j���.���=>�^�9�=��c�g��茠��c�=�k�>��о�Z�u��>#$�o�<��Y8�ͥ�ν���=$@�>��lku>�{�>V�:>��.��Q������+N)���S?$<�?�I`?��?{Ǿ&���~NнO�=�A>�)y>i�c<�g3�%�>�%�>���?��Ua�&�?�:�?	�?h%/?9n�)ڿ]���� �����̏�v�㽈C >2'�\�=1�.>V#p�nu<���=l��>�t�=��)> ܣ>��1>2>Q����#������b���T�m�D��j$��(^��꾣��b��yꜾ�Ѿ�Ŋ�����ϒR�ݽ���Eȥ�@퉾7?m>E2?��>/v?^H8>�9�>�a۾��<�}��8����/�����[+��D����i=�5A���ݼ���E�7�
J?�=���=��?�m�e-'>�?!��=�I�=}�k>6��>��>���>�H�>]>>�=>wd�����>p�ऎ���,��9W�4�=�򽩦�??���I\%�[�
�8U��P�ۼB��>� C?�Aa>�\5�����:��Bl�>�l���N�X�:�h�=�T>��>+�=�?&�L�N�l�F�}�"��=��Z=X�=>��<��f��/����=1��>��Ǿ�.�>o�>�SE?�*u?� 0?����?r��>i>�+>\Y>>]��> K>|j?d�9?�:4?i��>ԝ>!sž�xw>�%�=#c���=3l�ӿt�J��;��d�=_�� ��<R�<��
���=��T���W<Chֺ&N�>��T?�?��<?O�ȼ 
f��o�&۫���>{}�=V��l&?�d�>���>0J�>��&?ڔC>1\������k�>��>�|�
h��א/���>�f�=�Y�?�P?;C>/�������=�ǫ>�,?2+?@?�p�<�z=n=	�<�ҿ��ݾZ�3�(���ɾò �/k� ���>Ŷ��@������Z�<�g�=P�>��>}a�=P�M>1Я>ٜ>Y��<�3>��D>��>#9Q�B>4>�������lh�v����&=����=�x�=��'�)��8Ƚ�C�>P1!?ˡ>s����㽑�����T���
>�_�>�j?��_>Sv>!_��Y5� rJ��!!�;{?MHK?/C?����>��;�u��y�&?u �>���=���;SS���)����6��=~F ?�F>���^m��S}��%� �>�=]�,��9�?�Ez?�����gϼ��)��@u�hW�����;u ��Ľ����-�7���\�	G��	�8���~�Y>�ۮ>1R�?�k��h!>�a�kc��O��B+b�#$��O`��>��<�ļ�D>;�(�'X\���ھX�%��o�>�Z�>���>%K�>v#�>��t?�&>��>������>�m>�>^�t>vKV>
��> ]?N.�>^T�>��->�X���� ��}W���p<Y)�T?z=j݇=���=4������D>uB=PA	>�j�=��=I�ֽ ��<:>g�=�1�=���>�.?��Q�$n��L��O�;��r��x�>Mc�>R�B�s��	A�����>���>6�@?��>2�>�����˾Q�վ's�s�?VzC?۪�>?�S���2>����;�;�n?E�>���فn������DH�iVI>�~�>�Q����>��?�
�?��s?�:=�
��F���?�}ా�4"��
�>�$`>��]�O؎��F�G����#��D����M>P5��A�=CK�;���=�>��:���0>q���u�\=�y�:�=�-5>���>35�>
?�Y?#ad=L�
�h%޾r�I?0)�����V��� '׾��sK7>�>�e�M�?�kʽ�}q�ը���"8�-:�>ba�?�U�?k�j?>v���0�z�~>,l>�G>�%=`�j�wN��V欽=�>:U�=�Ŗ�N��������$>�E�>���`¾���o����ط�U�V�m,s������l��ھ�������=��}�p�̾����!e�����Ї�S�d��P�SI��y��-����N�?Lӏ?�� ���˾
�\�$9Ѿ�d��K��>�p������gx��� �a��ҜR��|�f	��;��ᾷ��²>�j�DAk��S�����
�>
��>J�8?~馾\��7H��~>>�?�F-��3���I���U���>F�N?�-S?����_�bz�;�BU�W�?$�?�J�>]�}�V�m����>e)?�F2?�7>v5��Y���HX��2�?\n�?@�C?�?��3"��ڂ��a��Gi?��g?ў�>g�H��ɐ�fڤ>��0?��y?��>��2� P���92��};?Y;�?e$��=jJ�>��>T�e��վ�{�=0���?�=H�?,��=�1��������z����>o?Z$�����@��>�g�[�I��;��p�$X���<�F�>���|s(>�{�>d�>X#�L���S����1�	�Q?�˴?��Z?
�'?�Bƾo)־��A8=	ׅ>l�>V;=u;�+J�>���>�%��:�x���?���?���?��G?�t��t߿j(���ʾ\����l=u�X�[�J>�T��Ee>��>6�������=Z�=>��:>� x>��e>i��=&f�=!��J�#����������T,�:u�R���D_G��2���MY�Ϊ����K��q���4R�����%�/K2�c䜾7,�>��0?�R?���>�%�>9��>>&۾&ݼ�l$G����Z�<�A��/���6��վc�p��G>=v̼��L3��q3?�n���$��/?�����=G��>�}��URh>|X�>g2�>
LW>Z�A>5U�>%��"�=$�)�]?>��元��E^�`�K��D>5����ǉ?4���4�tD�>]�k�̕�@��=�B??��>܈m�)���2A��,|�>7>��ߞ��	�9����<�T�>mq>?R�=�p<�!=�����n��ֽ)�S>Lr<M=B�ix�J">���>�]��$U=�l>D�?e�m?�.?�$>K�>a#9>�ܳ>҂>��>ԴH>�!�>�1?i',?n�?윴>�F=�h��n=��i=5`��zw�2�N�m�	� "� -�;�z;
b=��@���Ƽ�Pi=qG=��3��"���=Z'�>�iJ?�F�>�gT? ���C`��)�<�TW�]��>��D��>�� ?��>R�>���>hX�>W
�=݇��f��v?v�����G�Yr���V��?��>�ϊ>O��?�uD?[���@���꼟��>�,c>5�>��x?�{�>Z��>fzd>^�	��ĭ�����D��n�=��F��^Z��;�B`��9>\��<�D���
&;�D>��A>i�4>Ӹ_>3�3>f�<���>�<�>��=�O!=c�=>�J=��(�l�}<�����ν���=3�=/C�=}v��6�>�S��л ��l ��,�<o�?+�A?�G�=��'=iTc�3��1���Tt>�[?,4?�"c>���=����̳T�R�D�x5νNPK?w~?j�?�����x>c�=�]��.?�;�>��u>��]�X ������xž��2>%�?�%o>�ݮ=��N�F���, ��U�= 4=��9���?\�?������<����kt�����H+=��ؾ�Ӊ��Ἶ�nk�9̀�J{F�	���<��>�6�>���?Y�]�qp��2B5�9���D���ri�4�����>�
H><=�DL���;�|4�T��̪������>��9�ߺ`>^h?>x��?�2?庄?c��_�?
�)?�5����>V�>�2?�v�>���>6m<?��>�B�>��q��r�����=jE�=��<�Q=��!>�����Kl�b'>���<�R��4����f�p�p��d
=`=�<��=3b?���>�yM�ɗ�w�|�~�t=��_�]�s>;� >ķ��x 6��!�<��X<�>�#?��?�ؼ�x�Ľ޾�B����>�d(?��Z?��>�Y�������5�<d���1�={R�>��1>|\����V�z��q���>�s>c�=w/�=7�?�5�?��>?��>��X�����0q���>|�>]�b>���=��&��!U�UǄ��KI�-4�����c{���@�k��6m�>mj�>'}_��F(>�>��	��A�SQ>��9���N>�?ӲL?�t�>�(+>�7���$1���I?8��Z������2Ѿ�'�U>>a=>�� �7�?t����|�䟥��Q=�w�>(�?8��?8�c?1�A�m��
+_>uX>�N>e1<�+?�H���"���1>,��=��|�[���;;h�Z>�x>��Ƚ"ʾH�d�L�5����
4�׳x��LľR���8���#s��d'ǽ�m~�����&���ᘽ��G��5ڽ�y����0��]�yE��ⳡ���?�f?�V�<��㽓@��1¾�2����>Udh�Z��9���k8��{��77������Pjھ��!��#�!��P�>~���'z���i��r�G�Q>pU�=6P?�<��,!�(���|�>f�?9�>N/���~�KS��;2R>^�]?v�Y?���y<�a���һC=�Q�>*��>m>�����|��!��(�,?p�>���=�Q����ϲ�1�?���?BF9?�g��$,=�������c�>��?a_�>����xԾ��4���R?a�?˾?W�;��"���˫�+,X?Ax�?�wV����>�0�>
s"?"侈����=��#�(o">quM?��k>Di��$羕C¾A!�W/U>u�??`��JM¾g_�>龭�N�SH�=��\���<M?�)�V�	>�sg>jC>��'��Č�`�������ϏM?�M�?^hR?p[8?���F��Ԧ�=�>I�>gm�=]a��>5��>A�侗�q�a1�T?.�?���?tY?I<m�L�߿}������/����P�Yչ=UJ[>%Ud�N�3>xc>�$�<J�7�1_P>�5�>�f�>I�C>��;>XQH>�ʝ>����g������ ���|�V�-�>��T\(�4��Ow⽇�������t���-(��ӽ�E��ϼ;�`�=����M��>�:�>I[>3}#>� >[U�>R��?r����`�O�s�}q��9E˾�P;W\�6���g��ͱ�7��YIg�tȾv��>X��=]k%=��>ş?��Z�=��>K�>�8�>�F>�`D>x3>��>��?=z��>��>R9>z�>���=B�J��|}����o��K�y>�?�J��@H��j����<��!>�?^�?��Oq�����ǟ><q�<�����*=S�v=/�h>�P�>�D���Ӽ��/�*B2�ϟ���Z��QY>gF� =���Ⱦ�A��E>`u�>��Ӿ�u>Bw>]~*?~Ɋ?�.�>^1�=a�	?W>��>\U��%Ն>T�>��?+Ⱦ>]u?���>�?ҁ>�����7���5H>�_&=��Oϝ��'>�.�s�=�셾g��>%�޼X�Vd>>	?�=��|���$D�>d`�>'�%?�??�9?���_�
��[����+�>_N�>{��>��>@�?�Q�>{V?`�e>�(}>����6�N��i�>�%��A�₿ˇ�q��=�#�>88e?M?XO�Y��!�">�f!>�8ɺ�4'>�?\?�,�>ʀ�>T��R�.���I���_��J��(�)=|��<"�=f����e>l彑磼9�M>���>p��>��->yw�=��p>#O�>[��>{�a��<�g.>U�=P�=���94</>׉��!�D=�X��3��=!�L�%�J����>�;��=��;
Y��g�?W�>ڜ��z���� t�O8������>�r�>�a�>b=c>׍�>��˾�����)�����+OY?��U?B_>ftὸ3�<`� �B�˽���>1�>℠=��=^?�5۾��=��N1>[R?f?�v#���K���N�6M\��ܿ> �=��?�/�?�K?��AY9=R�B�MS��5���y���A�Q۾{�����)���I���&�������u�>m��>*�?�h>"��;y���㜿�6��fVT�pp�<nR�Ƈ�>�X1��ڹ������Dj�٠C��cݾ̴���ec>'P.>wMo>�?H�+?d�{?��?�4S>�*p���?���>��>N�>Ki�>��'?���>ຊ>�%���>�>!X�>����Ee�� =���=���=�=r�M>��=-�˽���=ן<>�*N= ��&�=wQ>���=��U=�7� >"P?[#?&�.X�=��g�g��� >��!=�EZ>jN9����[X���7=��>���>��c>��X�_�ľ�^o��N�x\�=4�(?ɫ"?_�d>~�$=k?E>@��X��'t>���>@8��a=���������.�H��>N8�>c�`=�(�> ؕ?tu�?�"?W�<>�0\�L����}���/߼��=��:?À���#>3�������U���Fj�H�9��>��0�F�E��T|<#��>�">�>щ=��B����0�=�V�>C@�>�?���>[K"?S�>��}>Y�����Z�G?�9�����=�� l־e7���;>�Q=>�*�5�>��
�d��ס��>�;��>/��?��?�)^?��^�������Q>�>>f��;��7�������$> �v=��F�+�������^>���>vѽU9̾ #۾ή���O���+2�sJ6�"R��_�;��� ������+>roʾt�p=H[�U�g���}º��wF>���� �`[���������?� �?b��>>��Ue8��J\����V����T�������4�����پ�ַ�cbF��+ľ����KWP�--J�;͜>��T��Ƒ��6|��L)�KB��ȲA>,�-?�ƾ��������U=�#>]j�<�Q�W��;����V?o�8?^���t�H�ٽG�>/�?e��>J&!>A*�������>�,4?+j-?�VO��ܫ�������?%��?"?�\�#z.�ɭ���9��Ѫ�>�:�>"j?�C���L�,z���g?��?�e?�����y��S�BZ;?��8?�7���@>=��>#w~>��J����U�F<"#����\=.>�=)=�Qt�W��엾#�,>Ϣ>Kw�������N�_��>*l��<N���F��j�����t�<o�>>��{>)i>�>zg)�+��~	���"���J?˰?��S?p�5?������aࣽoo�=��><Ԭ>uK�=M�����>��>IU�G�q�E��R�?`��?V�?^*X?�k� Gӿ�
��ʶ�����Ѡ�=�'�=��>>!�޽_ͭ=��K=혘�)v=�t�>���>Yo>�;x>|�T>��<>��.>J���i�#�aʤ�ْ��[B�� �����wg��{	��y�����ȴ�W�-���Ǥ��Bғ���G�����X>�N����A>��> �d>���>��
?4#�>����߾n�=��v>�R�%,���c��n����H8H������m�=G��_�#�^?}�n��39>��?���Ci?�x�>�н��m>A�i>�<�>v��>���>�o�>ᕞ>mQ�=P���e��>e�?<g'@���O�4_��/�����>�V)?y�R�)F�=��y�)���|��k#>.߲>�'#�w�c��9�������>>�㽼�������Z@>>o��>�H�=s��<k�ν�C�< ^:�m�i�k��="-�>Q�"�>1F�wEu�g����<Z5�>�}�����<UB>�R%?�O?�4?a3>%�>�Z=�1�>��A>Έc>��>7��>�X)?��:?c3?���>��ҼXǯ��?���S�=�w�ՂA�=����B=�	�<�$�=@�o�2)[=L�=���Tf�b��+�=� >c�J=e�>��-?b?6BF?�
<>#���rX�\���5h�>r��-?Ӎ?�m)?b-]>�T�>)�>1�!>=l4��Y���8�>���,J��y�3���k>P��>Z��>D�?��"?���\p���S>�ݨ=V>3Q�>JLS?��?�Ւ>On>��*���J&�ݮ<�Hj�@ɞ�p�W��s=v6O=á��A3޽ީ6��>!��>&��>*��>Y��>4y>O��>�Q?�x>���=��=Ch�=:�;uA��R>ҿT���ｴcܽ/<>���i\���&�<4~r���G�%���65�=Z�?[�>Θ����5q�y;�2�/�u�>��>��>���>�)�>z�d���4���>(~?щ�?E8�>�!���F<|��=�s`����=z��>�4�=Zi���M���2��Z�<bQ>���>��>�;�=PN�"�0�(V�>ô�<Q%��ޝ?N8O?��o�霽��R��1�`k˾�VM=x�Z�9|�� U�U�6�MP��#7�m��m��ǭ�>|�^>��?M >��=8�\�-���-y��ZC.��kJ=yWD��6>>��.�j}˾�̭����� �(�`����.���4>�8����>��1?k�9?�W�?��a?Z�>F/�"RL?է]��h?[��peZ?uxF?wI?�?�B�>|�p>u��>��m�-څ��KP�Q��������=�/�>zJ콸N���}�=U2@>�8�֯��=.�=^�<�Y����F��X8>�o�<��?�?5ߋ���)���F�Տ����=��=��<�K��������=������>��?�z>�to=޳�m8�~�
�`r
>��
?y��>I�?��^�+��=�Cɾ��B������D�>��=�vĽ3�ƾ��K����>^G�=�{?�����L>�@�?��?��?^�H=�߾���������=4���>Ý����-�������圿?dT��/#����=Bs��=8>	s8>ț>r�	>䊬=p���y�޽s�S=*ٛ>��'>ll�>�N�>��4?ɤ�>L��>B\���
뾸&H?�Q��,��♾N]ʾ�tv�h�>�'>>M��`�?M?�	:r�_ ��@:�$i�>���?,��?�h?�P8�n��]>��^>q=>�"�<�]B��������юA>��=��l����{R<�^>�k>����˳ɾY�Ծ�PC��h���MU��ra�����> ���Ծi!X���>��ᾜ7��_�����=v�T�~B�(�(=X/��lCν���5���֒�?H��?���=<��=����N8��r �=��=�N��J_�?��`j��J;��wK��2Ľ����&���}<���b�h��>=>��Y���?}����jcd�!�>Ҁ3?����-̾!��5�:=�L>/�l=�M���ͅ��������^�B?F50?�پ&�n�����=�?9ݬ>C=>%�<�L�$�D�>�%"?�:?3�w�򐿸3��O�(��M�?Z��?��L?�9-��I����'J@���>�ܣ>���>����H��TTg��Z�>�?�>��A�_R|�+n��~?�-?ᝳ�j�3>V��>�6?����"��S=�Z&��M=T��>ۊ@>������9O��'+�=�>��5���U>���>T���N��H����;!�F��<�?c��>Z�h>��>��(�2������)����L?(��?�oS?�J8?�<��v��������=�˦>d��>.��=�����>���>�]�FLr����?��?ں�?JGZ?9zm���˿�ۧ�@nȾ����O�=�/>�׻>zW��£?�1�>���;6Д��K>�>�>�y6>�X�>��_>��>1e�>u��P�-��`���g��W<��/(��Ҿ3ﴽv*3�v>&>nL�z�����s���0��}�^��=Pb½CA��Z�=���s�e�%>V�>��>+�>��+>��#>q�{�R����^�Yܞ�C��g�C߾&7۾l+j�`z>��G�*���὾���
?3<�<�q�=Ҁ�>m�.�->A*�>��=�dG>�A>x3*>x^>*�p>�9>�XO>!u>�J�=�Ƕ>�~Q>#q`�0����b!�6������p�>��F�J��r߈����;�m9����<`T>��������ez�3���߾>!�߼~eD�����X.�=���>?�>]�����|����Y�-=�YK>��I����=Έ����-=�^��a�>!:�+c�>��>z�?H�s?��=?��>}[0?�v�< '?V6���Д>%3}>���> ��>{}J?��0?�0-?�>��z�.��=�q>�x�	�={*0��)�=-i��V/X>6-=��P:=Q�=F���*%�>�nh>뙇�X	���>�S�>*�-?�?��?�Ģ=3������@۾���>�A��o�?�t->ˎ5?���>�0�>.�X�i>�x��g���Z>o1��2u���0�T��>�b�>��d>��M?�$"?9 ��-�g=�Q1�M�l��r>Ϸ�>�L?�h�>�H�>��<9��F����:�[�Ҿȕ�<X�ɼ+�<�g>Y�&�b%�>���H����<�*��Ζ�>r3�>2wt>l��>F��>O�>lx�>���{��;4��;������ڽ���>NX>E�W�#0����>��I���'��}�>�f����0�ڽN`����>���>�0>&���l�U�2�cx��h?j��>��>�m�>G/�>
��$UQ��_�/Ϳ=��<?w�x?��?��M=�fT��^���f>�!�>n	=g�.�C�꼬�ž���)>>��?4��>+�����R�����u �6$�>Jҽ=B�;`ǚ?�Q?I�꽞��<��@��8�H+���0��h�����������������F뾽���'�M%,>�Y�>�-�?�z�=iI����-��X��1#��Z��ۃ��H�>Iu�=߃��S]P���8��e���Й�����	Z>�ڵ=
�>��?Q�M?k_?,?C:?�����	?޻��-?Z~W>-�-?�?w9�>���>���>Qu�;	�.>X

��đ����=��۽}j#��J>��>�C/>#j��ӛ=S���C�cN7��W�<0�B>F�=(oI��͍=�h�>e� ?'�?[� ��V���V�H
��m�X<Dzc>Z7�GԦ=wID���e>��T����>���>S�?}0��]�e���,��B��=a��>Nf&?{9?N���	r�<�W�������,�&�u>�5�<R(���P���믾�p<��>藁>��d>~i�>&R�?�	�?�`#?�>�6���/���Ĉ�����Y�>$�>��L>���>��0�cOZ�er��kN@�a����̂�R��<b��>��=>$�>� �=���=�{�꼏��7>�i>W�6>Y�?���>���>���<'�>`qd�n+Ծ�;E?�헾\��Y��͜ؾ�Z���>�wb>n��g(?�	�Ywl��x���>���>���?A�?j�f?s8�y��U>�K>��>���<�Q���S�`g���8>MD�=�Dg�?����'C<rqU>�`n>�
��н�`��cz?������,�}�׾Mu޽-(����2���k�=K%]��^G<j�ѾWϽ޾�
��`g&>�zƾk�̽@�D�Ӟ���q�?Q�?��<�??=]��{���< �@9_�%ʽ�N�<,q�󷲾��߾]e���Ⱦr�0M#���l��5�>J-I�����ںy���'�v�8��*>��.?u;�|��F�!���r=�6>G��;J��q���ę���!��II?}�:?�~�f������n >G?'��>z�,>\��<�۽#|�>f2?��(?��T�깏��N��'!Ҽ�'�?�F�?8J\?4��'�E�{�i��n�����>͠?�4J=C���K𾼤P���Z��?�	?�+�|���>���h>ɉ�>H�(��->JK?�9?/�����>$=w"��-�=������=��=]]x�;�P�B�a��H�>;GX>�֦���=z&�>���a�L�R0E�Ǜ��)��b�<�H?����>��`>&_1>,(�~Č��w��7;�g�M?U�?��M?r�6?�U�.�cL���X|=~(�>�ݦ>��=U���܂�>���>��Ul�S����?��?���?@>Y?Cgj���¿|�Y�ž�0��c��H;B�W>(��O������>�B�=�����N�=}�1>8�=2S>�;>�b�>�'V>����* ����Q��!X�2�+�6j	��"~�t�;�uX=�r������������Z�9��.�ظ��E��}��&�b��!w>�?ir�>&ʘ>C�x>���>�o�I���%�A���彴�������ȵ��4���{����Bl������1�C������>�s޼k�]>~��>�О�2&V>�$�>��^=3S�>Z=>���>+�F>��X>@�<>�}>���>復=��>���=9v�(.l��3[��5ɾw��>��?}�$����=nJ�������G.����>>q>�y߽l^��3���R���۷>!�A�	�9��w�F9>��>P�=�c,�ܬ8�ϋ�<��y���v��ZAV>�᭽��>��;�`���9P�[A�>�s����>B�>۳i?��?���>��=���>��)>�,�>�}�=�?#a>J]�>Tr+?��?�x?�D+?pN�=�b��Ǽ�ݷ�����K�߼ň��ED>�=֣%>��־K�=���'�O;���=IJ�=�����<�$=d��>Ю7?��%?h@d?q�n>b
x��8�����s4�>.��G" ?}�>��V?Л�>���>��>GU=䎅��7>��>AJf���s���"�h��>Yɨ>?I�>��b?��?�"�ɯi�]a>����ڸ=j��>0�N?���>$3e>�K>^�
����5�D�7�a���J����A��v$=l����qԽ�/"�F]���`=��>�3�>	[]>Bd�>ַ�>4�>���>��>�|���>�ʷ=��=Q�=(1�>�j�=�?��m��v��<�
����=2P|=@p�;�=�Ӣ� 2n����>��>.]==��=XS��8�)��j�`�>CW?�3?��>{��>�y��*r���#���>�L?��?�3E>4���=@5<<��&��3=$�J=�iN>�����3ǽ�Ԉ���J;���w0�>U,�>4�a���zwO�ǽ�o�>>�=�4μ[n�?HEW?s|?�\�"� �E���5�9����e��"ݽ�c��������>�HvI�� �O_��;Go���o>�l�>|�?y��=H�=x1�Fy���z&[��Th���(�cY?��+N��� ��H�n�����!���Ԋ��E�>ٖ=��>֐5?0:?z
c?��(?��?l]��t?��;�O,?D�>M�A?�?Qd�>���>)�>��>�1�=q ��8��3#�<������H=�&>U>)
�=�pһ�&8���0=b.½����3=�ͥ=3�>ퟛ=�b>��=ko?a?��G������M�+ܻ���X>rf>>�	0>8�����N)>��0��l>��?��Y>�����v��8%����Yn�=�E"?q-�>�ǹ>?M��c���?��4
��Ws=�u�>>�K���������bx�� ��>�t?�%�=K'�>[�?�	�?s?^S.>9����}�� ���gƽ�p�ZL�>������>�@��K[��ꎿU}g� {��he>�q�#E<%�9>	P�>�0�<C�=�O>/
.��*�<�?1>��>���=�3?u�>��9?hּ`_>�M��B����;?�j���t�K�}��Q����R���=��!>е�=r�?��Ͻ[aU�����T�r�T>���?n��?��s?�!O��"ܽ��q>�ޗ=�
C>����:��X�=K���t&>��=
���$�~��A#��Ղ>C2�>��df������>�=����vgR����qP��p�Ⱦ��پTҠ;�Ԉ>�2~�������پ&>>�����Ч=����5�<ݲD��y��#�?���?��N:,	>Heh�O�=�̓��I��b���1��X��j�>�㹾���@ٯ���'|־�ﾹ��0�>�HV�h���!{��(����ęC>G�.?��ž����J�w�p=y�>&s�<�}�+��C-���:�S�U?/:?&�꾭����A�S�>P#?���>�">�2����t��>Ȥ3?`r,?��ռ�܎�}���*��s�?᝾?wC?�����'��<�,�c�j>�>�	?��>������}���CJ?�f�>�I�>P�
�o���1��u�>��?�c��fZ�>/��>���>��{��bm���<<k��r��q$>�i�:C�<�)��sĐ�z�����>
7�>��;���K��>;;꾛�N�#�H���[���4�<�?ڈ��>>^i>�L>U�(�#��;͉��1�T�L?r��?�S?6e8?^��0������Ӑ=��>�Ѭ>��=�����>���>e��pr���3�?�F�?}��?{[Z?��m���ҿ�O��� ��� ��;~=�m=�>�X��#H��:ސ>�8C�U�V>ʙk>��>��>q�p>�">��L>Z��>�w���,�V���4t��
a�G�8�����S�ԐC�ÓX>h�U�f����k]��_�*���=��p���/����=��B�A�$>�%�>�"�>(��>�d=jrG="u��Lƾ�8G�_���1C���;	�����n�ҾX�������H��Iׅ�n<Žt���>��;�hy�>�<�>PA���(>�A�>wga>N�>\��>��<>ق�>9��>(�>0�>���>�O�=N�>+�=�$��@mJ��H��u	��{�}IG?�s��׾&Gi���#��X0��^]���2>Oپ=��M�������:�>:gN�OA��D��7K�>�D>T�=3�g��9�?=��v�8�[���?���>�n��@-��A��.�����.��>j��vrB;�H��ؠ?��?�)a?�9��?�ꮽ��9?��ƾ��>m��>�n�>��-?u�T?�vH?��?���=�1/��%=��0�GWv�P!��0�;~�'>��3=����w���=�.�<��&���=�<�=��;6�m�!<W�>�a8?�?��$?������<�Ҧľ��#>�^<ц ??B�>Y?6:?���>���=c�x�!������C�>xk<���K�N��c>0]	?�D>�mM?�`?���=ָϽH�)>?���>m�?�25?��%?K��>���=�}�ȿ��I�f��+8����'��
:>���={��i?t�G�B�;
��=����sE�>e�n>�>&�>�.>��>�EQ>f%��c>Q�^>��E��#�F�>�5�=�RY��D>�ӽ� �\F�����=��ֽe�NK<l�K=���>�k�>eo?��U��=���G�t�޾��>ZK?��?s�n>�>��$�y��u��>�9��T?��r?�E�>F���(�=*W>&J:���0>�r|>
�5>?	�:	�#����E�<�>�=3�"?�ɰ>MԽ�W9���l�o侃��>Ca�=V �VP�?��C?|��)�-��?��3��;R���پl���+�O6�<�q�:�����2����D�����>�\�>��?"B�=��=(;�n���`��WTY���1>�V꽇�a>>=Q�ч����žm����R�oV���/(>4j�>��M>m��>p_?B�0?��I?�o�>,�T>�콽?H*�>�K�>��>��>�K?�?G��>��>�ú>�E�=2ݽ4,&�El(>^��<i�=�t�>F��=F����3�=�����U?=ə�6��=�4�����Ł9> �J=�5��G�=���>'p�>���T�@�uΫ=���� ����>:�����x��ܣ��>��|��t�>�i�>ڎ�>O�=g0پ8a#��پe0�=�&?H?V�>�h��9�<J�Ѿ��o<���=�^�=�p��q�r�qv辈���h䂽§>���>M��>C�>,9�?DM�?��?�)Y��������������>�67��>���Q��>SO��ۯ�� ����z����=�a�> +H�씜��e[�o4�>Ku>H�X<kW
?{f(=�/۽@~i>B'�>���>pV�>��
?��i?���>J�>�I������%I?�L��KX��С��X;�^&��w>�!=>O���d�?6��%�z�#���y�;��
�>GL�?ب�?��d?o�D�
O�Q�Y>�[>��>$(8<o :���������7>��=��z��B��z�<6�X>�u>��̽f�ʾ�V�`�?�iN¿:�]��I��[Њ���%��(�\r����>�b�>=Z9о*�D�r�4�������>�RD���2�D���8�/��?&�?��Ž��!�?<�O�%��:;��4>�tᾯ�Ͼ�_ʾAFf�J�þ�Y}� 21�����O&�qK���=���>���u�Ww�X�=����<.4>��?|��z� }'��I%�ذ>`+���@��R���w���"��)�5?ʼ?���m2�-�K�ᾁ���>4��>]��b��o�9��ԣ>?�?�LB?8���ڐ�6{��X����?P]�?��>?�>N�ٷ?��^�����F?��?�s�>�ٌ���;����-
?�W6?��>���������IC�>�V?�$L�ql_>���>|��>����Ŕ��z(*�|-��у׻^	6>o�G��w�0�b��G�ml�=���>g?v>,�^��䧾�D�>=;꾐�N�ަH�u ��f��ޒ<��?H���>�<i>ڧ>\�(��$�������� ���L?Nl�?�R?pe8?,�����T����p�=���>�?�>=�=�d�iZ�>��>��@Or��1���?���?{�?0,Z?��l���ԿWz���9�����5j�=깳=#3<>^�ݽ�G�=K!H=묌���Y��]>7!�>��p>�z>�-V>=#>>`?/>��bF#�N\�������C�����o�?�f�|	�(bz�����6��w���¤��y��e���(J�� �KRB�>������>.�?�7�>��
?���>�5�=%��ܾ9K���A����vg�ꊎ����꾞�6����x����l:��0)��s?�ވ�r0>�a�>��_=�g�>��?�ɓ>��~>�>L�!=�ʷ>9�M>�v>ne�>2	�>���=-��=䩥�������d�NJ�� >��>$_?Z��9� (�b�M��R��
Ⱦ��>��?���>,������ꍌ��:�>�Rؽ�7d�����>j�= |�>��]>6"�iF�=����=fEW�7�>��=6�p=�s־�H-�r�=�=�>2Ҿ�)�C���o>�bN?v3?b��>ex>���>�\�>���>X�վHC�<�W�<�4�>f�?�ry?s��>��;t���=ն�=�D&�{�=����;�qO<v���H ���>��<�x�=*pӻ�=d�=�yR=J���oY�|>�b�?7�??�;?��'>�A��x���a@޾E�9=F���Ĭ
?��?��/?Na
?�)?�[i>�J=d��i*�A#>/6����z����=��>�Q>�F?�9?��L>n�g����!g��B�>�.�>�?�?{�	>^#�֝�7п��"�Ų&�򲡽�}��cɚ��-�TڼK��<��I�:��f@5<|JB>{T�>��{>v*@>Ft3>�>��>ӦC>| �=Ћ�=.ĺn��<���;"=%�ἃ�+=��"�m�cZ���k���N��	r��_ƼC����,l����>)�>*ӎ��F���žuG�������!�>�;?���>��,?]����¾$oQ������;�?��R? �>�e,��C=�(��=D �>l�7>z>z=uv5�Eנ�k����\B�*?:>�>���>2�)~J�s�`�<�Ҿ羽> 
!=��h=�|�?��i?Rf��Pp��ԑ�00����F���9�,P�}�'>L?>�Ѿ����? ��^$����[�>�D>ج�?H����?�wھ����n����;�W¾(�ᾎ��>ڐ!=�-�=|Yh�ʰ���Ut��`;�q�q��p�X=�1�>X�?yfE?
OV?5D�>�ד>`������>��>�%�>�r�>٨?��>�,?�,�>LR�>���=w>+Z�۬���yJ�o�<�[�=�(>}��>���m��=�~�<sЄ�{��V�=�)�R9�T��=��6>�	a>�p	>]_�>3}#?�@˼Ǽ:�(���	^���_���m>ƕ�>Рż�Xb�a���}f>$��>2�7?�D�>�jX>%=ľ����L���K��4	�>��?���>�6!>kvz>a�����?�S����=p=䴧��Eݾ�6��2�T���!>��C>J/Y>�yJ>��?��T? �+?�<�Q�1����X�ը}� �ƽv�>��>{p>�M���.�穉�_kz�a�*����<^��[n>��<reE>���>�iv>�=��I�=�˔�����X�>UH��%Q>���>��?=��>�]�>�徸����5?_��F��ĸ��W�V���>z�p>f�R���?�a��wn�4풿=\G�4�>�W�?W@�?[$\?H�d�:q8�7�>]]>�e>t���ei����$���˼�b>X�=_�Ƚ8���$�=Q�>�{�>�B)�do���F��'���Iay��6ľ�]��r����'��b���ؽe���g<��.౾E̾��ݾ�_ܾ���w���������������?�s?y��xf	�[�x�D5ɽ�M��~D>�
 �߬\��ԓ��l�+E�����0������L��������!��?әi�Ft��B��V��V�=|��>�>?�þ�;�Z'��:�=yï<gt�>Ip�(��#̰�%S�li?��?�����ھ�ŽܩT>��>زi>ׇ��=������v%>n1?R�/?L@:��ڹ��������.+�?*��?�z^?�	r��� ú�;�=���>�[+?��8>Gc��$<Ͼ5	��,�.?`�f?�՝>�X�����1O��`�>�˔?�*�����>��J?��q>�Y��@���n���7�����=1�>Q���$r�pֽ�3�
�F>Ǧ^> ,�=>�d�
����>f9�X�N�hPH�4��5W�Ҩ�<�q?����>4
i>��>A�(�{������i�7�L?�^�?�S?-N8?c!��j�������=��>q�>&0�=��'�>0v�>�]�p\r�#��?���?�{�?SGZ?�qm�T�ῷ�����¾Ǫ�[�;>[��=�4�=�����=��q���P�t���y>=s�>Qg>}eC>�Xf>WC?>�1>V����%�d��-����,�!��%��}���X;x��)���Dh̾�,��@ݽ�.۽����Ͻ��r������z>��>ơ�>�"2?K��>��
>sU|�/���,(�pjp���-���婒���!�H˾K\@�����`�=ʾ��������>�1��U�>Q�?PI�=��`>��=�xg�~������><��>��?��>�`U>O�{>��9>?&�9�S�>Y� ��zW�6�e��]��>��>fE?~^��Ƥ�S������o���B�=��:?��
?_O�5u��{�b��!c>��-�1n꼆�u��XW=hf>���>���.b/=�L��R]P�YZh���<�p>N�~>��<�gU�
������~�>�־���`T�p ?:!?��	?�->�h�>J>=���>.->*}��d��c(>���>�BS?zdB?��=Ó4="���->;�=���#s�w�j�b���<�Ү��bw�`Б��F�=��=i|�<�^ܼԧ+�6RѼ1�+=C��>4�F?q,B?\�;?���i���s���Ͼ�t*�^̚>d�>�N<?�S?��?�$?/ß>�vq�־�˾
p{>� '<LI(�53c�/�����>C(3?�+?��?���<���o�=4�>�B5>���>�n?Q�>��>���=+@��-Կ������7=��Ľq
���E�o�4�g�<����2*��p�Ϝ]>R/�>f��>��\>R:>3�>��>kP5>��=Rv�=iƉ<��<��̈́�8�4>�E���Oi=���h�>^3ۼ�����Q��Di�E$�|���GM�(?VZ?�ӥ�������l�'^��--����>�n	?���=�>?�ǻ�S�4�W�he�
���8?IdU?;Cf>d2���=>�Eֽ�;�<Y�>n��>��=̇.=h����ʾ��=.m�>���>7I�>G��.3�<r>��A��gp>�01�
�$=���?��o?�ju��u�_rH��f����:�/��>�����o�=�A�=}��G#K���6�i�ɾRdݽ��U>ɮ�>DÛ?x�=�f�>7����8���"��H�V��o��=}��>eψ=�2��ޒ�;Ծ��<���n�ǾW�ߑ=x��>wk ?���>�D2?G��>�G�>��u���>�أ=�Ѥ>|�?~_$?�@�>��>�ƛ>
1?6
�>n�{�����i��>ҷ����=.�=a��=��E�u�u>%��;���g�#�6��7 �����9��DcO>�S(>{]�>���>5�?]��������	��<m+�>?4�>��)?��	�����C��Q,��ꢂ=q�<?��?J�<>
�W� �j���P��=�h�>��?~�>:�n�W�q��>�/�R��c���4�=/V���i��M��V����N�2�g>�?�>JPa>��M=�/�?��?�Y?Fy�=�܌�5
��c:A�52�  �=��>M��>�ͽ,��#��KD��l�f$*�W�9���n���>�=/�8>2w�>7ڼ��1=�D>˧�<������;>�&�옳=Lf?E�=?P�~>��]=�*׾.����??JĖ�
l��������0�3<��<>U/w>!<��(��>r�����w��V���LC�EM�>�%�?x��?�hN?�j�,�潷�q>�
J>��>�1<�[G�tO���ê�C{f>���=�}I�]@��0I<}B?> MM>;���\��
j�����t���d
�������1���x��ڨ�����[ >�ď���>$���^��1^}��=�g/>��(��WJ�=�����/�ﮤ?¬7?�������=Nu8�#���2Tx���z>����J�ἴQF�"m�s�.��f�a����8s��i���h���3�9B�>u�2�8�o�8O@�)b˾h�>,ʡ>Q=?�́�L+M����δ=���>�>0>Ψ��t��7��p��<b�c?��+?`�0�:վ�tJ���?�o#?l�>�˂��d��am%>r��=�:?��>F-�=�ׅ�(���B��e��?�(�?�3E?��(��ʤ���>��2?H5(?���1��d����`=��?�EQ?�g?��m��:����"�h?쨣?qMi�)�w>N?j��>�ۮ��v��9�������=(��> Y!>ɴX��%��(�ؾ����M�>	��>��]H-��<�>7�E�h��M5��	\�$�=)=��?�����:��>?��>V������L�鸯��8[?�?�?r#8?wSѾ6ή��ט=y�=2Y.>`9�>T]�=+��»>��?#~��^�$��`���>�5�?���?�O?�օ�$�Ww������y%��R�7>��F�n*P>$D����>̌�9������v)>{m�>��0>-
k>��>�L>�^(>�z���o,�8������]f+��N�
��(�k��M�����U�*��D�x�о>��?u�p� �	��$�:�"*�����H�>2�!?�[�>
,?~�q>kf�>C���J��zC���<����_ܴ�����9��o�׾��н+o���;�=ᘳ�?-�ʆ#?v#>����=�?>����RG>�1Ѽj�=g�-��
�>nK�=J��>뇺>�J.>`��>
��=����84�>X����UN��p���j>�N�>n3C?Mc�@u��C��m(�1#C���>0!?z��>��(�+*������	N>/ >;><�Ʌ��|�<C:>9��>� =�Ճ�	���c�O�Y��7 =GN�>��b>g$�m�ؾ���e
>�!�>� ��L���z�<:��>�K?�(�>�_w>���>��?�;>c>)��=�|ڽ��>�3?n�V?��&?3�>f�=�@ŽIM�=��\<��*�(�=h�<��>���要�\ۏ��&>á��^L��o����=Ꝡ<�h����<�I�>,~r?�?]d?\]e>�뒿킑��8վM]{>�1:�k3?,/?4�H?��V?n ?hf�=�,>ca��P���'�>Q_�cL����k���y��>?��>��C?La?���<�%���=/'y�v�>��?�%�>'�?��>f�i<����п^-��:#����W�L<�b�:'s��'���쪽,�����5nx;��>z�>{@>�V6>��r>J>/>o��>�YJ>��=�=�m���d=J���6{u=�:��sؼ��0�;�$�=�ꊽ��[�u�n���Ǔ�::�"�s"?��?��$�i���L�u�l�۾�#��ښ�>�w�>��>���>���=�
���U���9����0?��[?hl�>u2���=��4sͻ�r�>G�>:S>e��	���r��h������>�?ߢ>���$ S��yh�!.�Jn�>����V�=�v�?N�w?�{���j���1��Cx��]4���>_0ؾ�R>04�5�ݾ�n
�P��Z�!˵���>�d�>_S�?�V�rS?��{����;�� ��<�>����Я>Q���8=FԾrq��3��暾��v='�nG�=�_>"�>,�?Q�=?���>�ޕ=:�����>\��>	,�>���>�"
?p��>���>>��>X�?Y�>��S<`���:��tr�1�N��+>�i�>:ҹ=����_w���5>�xS=|��ּ��=��ν��>)8D�Ǥ6>��>�]�>Q��>6���]X��/�����`����=v��>c�?�#$=�`��x��E�>�2?��>Y�|���#�����Й%={�>��(?
d�>�$��|����㊾����[.>'\d>h�b=�~��!޾q*m�Z;���a>׌�>}r�>zc�<�Ē?��r?�CJ?ߊ>tn��lv���y��<~N�=�o�>���>�as>9N���+�Rup�(#I��G���>8����o>./�NM>��>�r��˦b�]�>���mY��ad>���;��>�2�>�x�>���>F>��h.���>?W�ؾ~��
頾�����=��:>Ǧ>���j�>i�N=j1��4��4-f����>�ػ?�@�?��8?�<��Q7W����=���>��&<��D>묐� �ڽ�Fr���'>
�=o���о��d��>�>iC>L#�s.���*��3|� ޿~{�4���%Ǿ7-���&����ξ4������[{���d�����w2Ͼ/��xG�@!J�B*>����r�N���?^�?��J��/��d�>�����z�|��>n��<�88��t0��>�W̾����`B�����b)��V��0U�8��>�7���lz�͒;�i"��!��>��>�i?!�;*����>��s>AT>(�=��ɾՌ��Q����V=��m?�(?�<�������=��>��>o��>�$���R�F���>�:?E.?�f������������=��?-[�?.^:?f�ٽ;����*�;��>��5?a�e=�)�E���*==��2?��m?�'>t�������� ���[?,��?o���yw�>�H8?�),>��R�:������I>y��>j��=c�� a/����#�M�L>5s�>˒Y�ž��>�)�PRR�=/,��i��]=�ڽES?'���*ᔽ��>�q�=j�������J�g��L�$;?9�?��?��@?�c��Bо�pl=�����f>|1�>�>�u��!>uT?a�g��%�U��C�>#�?�0�?�?�����U��_T��M�ɾ֔
�Qj>=K�<k�=d �.a=�P�!U�^A���O>z��>U�=�O	>F�y>�8=�@�>q�����%�h��B6m�c�D��B������-�x!�9�Ǿ�3���ྡྷT�/��R����_0�Rm��=��)����e� >�U&?���>�e"?���=�u]>0ſ�� ��}���(N�s� ����m���{ؾ�ۼ�2�,��\�Q�a��QT<a+��s&?J�n��x�<q�P>��6<[w="��>�>������>�/=U��>���=��=�e>��>c��=�+�>�
>��M�M�K�&�/��w�>�F�>�;=?"�f���hW���������l�>_�k?��>�%���w�7.��m_">s��<�D= ���:�=�D�>���>U���T)a��jl=(��{���7�Q���>���=p��W��5:��s�U>���>��(�2���c|�=%��=�eZ?ݺ�>�\�=����>�(+?�?`<�>HRӾ��cFT?�d?>?��><[�=pآ��4q=���<�WĽ��=���������=�@�,���9�=���;�=�K�=,qu>�XB=r���`3�b�?��??��>�#+?��6>��`�y�s������>_��>.�?0�>	?��(?Ǿ�>W�=ʺ�=���LVؽ��?g���A������=�~�>�Ⱥ>���?�vR?�n>w����T�{0]�c�?��4?@m�>�K>��=��<Ή�Q7���N��⡾�,>j7�	2B>�Ӈ�nѼ��	�e:�IBھ����Tp>>�p���`���q>/���]�>/�C>@o>gzO>��$>/�<,�)�YQ�����Y��=�x�=˺�� �w=��0��_?=+'��vL=$?�=�Լ�g?{l?���;��E���x�02��F���>�,>2[�>��
?�HL>?�����C�jL��[=�%?x�q?j��>�)�N��=82_�����E*�>zM�=&��0��F�L����H>`9>�;�>t��>�%=qR>�'�C�����v>*�a=�6����?epW?%�������ϾOq�����f�>���8�*>���*[ �-'-���7�7���Đ�}$�>�>�`�?b��-� ?1ǈ���3����3��8��\k=;�?!�k>��J>�<��پ�9��#0��>S����6C�=�:�>I(?� ?)+[?'
?�?e�n��>[�=��>�6�>m?�?y��>� �>��>*�h=}���`�O����K<<�.�=�=�'>�W+>p�<�i=|�&=�d=�U�T���;)�<�"�;|�9=��=���=��>��>W�?�Ck����ի�	e����!>���>u��>��5<K���5�Ͼt�;�7�>�O?�� ?�i%������d��O`�<'/�>�?`��>���=6`>,���ͤ��S��rc>��b= �U�����P��T���w�{>��=���>�:>�K�?+y?��A?# >�Pg�����K�y�����$>�>>q?���>\� ���D��{p���J��>T�'�<� U��DT>�S�=va=4�>��x�~�=W�>�z.�쪙�X��>d��5I
?f�?��>tm�>��<��ľUr ��;I?+e��B��>��_�Ҿ����R>ٸ?>TM��?d��V|�͒��r`=���>;2�?ӑ�?�Zc?��J������\>^<V>�>JV'<�;@�u�!�*q�=�4>5��=Sy�n~���S�:D�`>�'~>�ν�ʾ�����J�����~^�c�v����
Yl�ff���/�����6M���r���;�9���yL��{���^t�%=���B���"��W��?��x?�P&��v��Ef��v��� ���J>^�F�M崽�G.�MWp�����׾�� �$EϾ��'�)
���ﾮU�>������a� �L��Q�0� >(j�>��?�!���A����$�#��=e�>��������f°�>���Z,l?aE?�)վ�閾рH�M�K����>��>��}�/�(�Nj�U�v=ؘE?ʽ%?c�+��ƥ��S��BJ���?"��?=S>?�s��"�B��ثL�y��>�%C?�:�>./#����U���c�?ք0?�S�>X��=���=�\�X2�>i�x?�օ�\�>�?
h�>"��<8����ŭ���о����J�>24��D꼩�Y��ϧ4�_��>E�{>c8���˾w�>j�����]���9����4[���<��>���@�@>c>��>�{.��r���Hz�"^:���A?C3�?�9>?KkD?��ʾ�#;����`�����>���>�3�="�:���Q><�>3;��{�+�����>l��??p�?c�?��j��D������_��7��ۧ>��K=��$>ŋM�z��;8���Ʊ����;e��=1q�>FZ>�t>	w�>}Nv>�^>�F��\�!�!v���t��"0=��$����QS�G<�%�����̾��þ�Eɽ�����`c��	e�Ӟ��#�Ž��L�>�T;?C��>��G?���<��>E�����E���O��,���Z�y�R����5վPy-�Hѱ�BA�9(�5.T�?v�>���թ> ?��"��j�=;�r>~0>�U)>�H�>�He��Z>��>�(>�p�>n!�>���>�¼>�m��0���1��L�E��>D�>m?Xþ�����u����� �f>\T?U�>�7��px�@����>��<Zr��W����
>H�i>�֏>q}>'Ip=@[ɽ�r��.#� U�s�>�r=>~�<�[n�ޮ-�B�����?�V����!�.�z�>BX?@
�>�}_��2�>�:?��#?�D�>�ż�V��D��O�5?�?U�?i�?�)5�=m�U�U�66�Z  ����:����'佘D���� �ZhP��b�=�ļ�d]=�^x����M��l�;�F���9�>ycJ?h�?�?��R�~PK�QQb�u�P;�>�s���>��b>�??�"�>���>���<�v�<���F�þ�.�>*w�=��G��X2��Rg=��>���>~;U?�s?�t �W�|��0����<�x�>���>j�?~�>�@I>!���)���ݿ����q �6c�<|���\r���Y���]+��㽨6+���G�_Y����AY%>��>�t�=f�=>���>֮?��>��e;-^>3���A��E>��=3=�k���F����k���;%!9�{U�5r���OJ��8�5��=�Eϼ�?0L ?�閽;ܽM�� ���*���ܫ>��>�z?,��>��=����B�e/�����.?�Tj?���>6�A���=r���x�\w�>�V>�
�=5�Y;�ɓ�ӵ��ɗ~��O�>+��>y��>R[��I}E��9N��]�:��>�sW;zFp=�?H=�?b�J��eԾB�c7��y�-�V4?=����>�>�������z/�Yf��b���3O.>
M�>���?�Ͼ��>����pu�����qF���K��J��>��?\P�>��=-���A;�sP���Ⱦ8n�1!>y"�=�j�>[v?@�?U�_?J�?�Y?���?� �=�W�>7�>��?��	?�O�>L�}>�À>Vv3=���5�������C6<e���=Y�>��'>�<&+=�J=��<U�$�@H����<Z��;=?
=�9�=���=�%>�V	?�((??�=�����,��츽�D�>�y�>�?��X�V*
�9H��S�>
�3? ��>Q��>�ݽ!Kؾy�ݾ�X��Y=�,
?8�>�Ų>�7�K��=2?��D��Lt:��n=��)��v���߾F���//��z�=��0>F�+><�>���?�e�?̡k?�4m>�L��j�y`i��ržxռ]�6?��?ℶ>aw��)�ʎ<��n��T�j�½Oc��8=S<�Wi=�^�>� \>X��=,̘<�j>���>j���+��>"
�����>:;G>��?�V>�>#.��BȾ�}8?Z�l����o��^��H��|<3>^NY>�>�'?M�2�	=`����6�gO�>e¯?p�?�)M?�G����J�A��>`w�>��>���vô�O��;�F9>���>�0�=WX+����N7>��)>��>��=mQ��^M׾b�n=cӻ�i�{�lĖ��&f�g�I�/AȾԞ����X♾�P��%>�������ݾ��*���F'�AS0�E�<�?����?�Mf?ەξV�.�Q�_�ｽ��pa�>�V�<=�=,�]�0q���ľxE�r�T�|Ӿ0*;WTھ����g�>�Q�8Z���z�z�%���k�L)D>k^/?o����l��Y���JU=W�>��<�J�e�����^���=U?��9?ǭ�z{��&���D�>�	?[l�>02>N���˽�҅>��6?�)-?���O���芿�����u�?��?h1;?�|2�����+�������>~}?I��>�+���D׾;]���?ߺ4?�o�>��
�GzM��M)����>LTG?�=���.>)H?�(�>&7���I��`�=�C��2��<�y�>%(8��ѽ// >H�[�6���m�>�Hq>e�)�_Љ�I��>B;꾢�N��H���n����< R?�a�Q�>0Ni>�>U�(�X���Љ��P���L?e��?"�S?U68?�x��w��!Ч��Б=4�>U׬>e�=�P��Ξ>c��>2辉\r����?#C�?f��?&KZ?�zm�Rzտ�ǜ��:��@O��+�->���=�	>����y�=TJ�=!�R=7�<��$><~�>��m>�>��!>�x>�{k>e���=�!�L^��01��bAH��l���$�Ės�L�$�s,x��� ��;��|��½������n�j��!�
�>�<fqL����=�?���>�Z�>%�N>�e=zj���˾�|��H�C���۸��վT?�_f����'�+WԽE���
{����)]?��g=7��>+=?�Sü����b0�>0��=�p>(K`>���=��>X��>ȩ�>{�>u�o>��=%e��&+>t���b*����F�Ԑ�z��>�Hf??�_�����6��V�_%-�l�?��?�V��(ZG�2"���y���W�>�T�;=RL� ����;�=~6y> ��>��#>�����=��ż�l;N��=9#>ph*=Xq�=ԓ�vͦ�Oz�=P��>�{1��u�>�?�@?�6�?$߆=�ԏ���-?�G?h�?Z2�>ѳ>��(>Z�<>��%?B ?�C^?�4?3>�ʡ�i��=��=��Ծh#N>6��>
9*>��C:��L�?1����&>� �=�t�=�۴=s𽿉t>���=?�?�D.?���>s ?9�z������b�����i�>'�>�׿�>��>�?n��>��>W�@>����i򬾆�ξ���>U�
>o![��Yh���"��>[u�>�FV?��#?�0�O5��t����=��>t�?�`4?�!�>�N>����J��N׿�, ��$��Bt�o�Ƽ�hO���H��Sͽq��3���Ӥ����=�Qa>� �>L��>Z�W>�B>�s>�f�>O'L>���=��>����,� {^�!O�=�m�,��Eཡ��qTź�䥽 ��4)�C!�<�;��������>%?�I�R����ʬ�����2���>�C�>A�>���>L�B>@��x�&����.>?�<?	��>�Ð��^ܽ�5��hEY>S��>�k�>�ü�Z��|�J(��x;�D]><��>`�?��=]A��-~���þ&j�>��>��T�Τ�?i�w?t���d�=�G���i�>v��HU>���=��#y��;:�SJa�>#�X���<�=
w�>3ǽ>�t�?00��=���,ȿ�ޒ�G	��z���?�<��?\X�>[���2�従H2���"��ĳ�<{��4�=��m>���>\?D?x�O?�҇?�U3?>|r>%�⾱�?{��>��?�0?�m?�T�>>��>�Ȉ>���>P�>Y=H������Fx=� �=�<k>�3^>���>���<�+�}e�>ecڽT��=�Ć=>��=&=�1�=Yn]>�~ >�>���>N�?2���m��"X@��ܤ�CeJ>k��>ى�=g�ͽ�x���}�.�����>�RD?rX�>HTU>wn����O����e=�o ?�o�>	yh>_m�<�|*=�����ɽ�W���.[>�g�=�ʹ�+�$�4�����<�4�>�X�>��>�]�>D�?��Y?r�3?�襻E���-��r{Q����^��=!$?ޕ�>�ru=g ��H��x�SEW����r���'+�;4�=2�64g=/�>���=<�>)�=�$=�=�͡X=��X=ܶ�>|y�>�,?�x�>�o8>�~Ҿ�� ���?}�ӽ��������I�`z0�䕣>`��>z=�h>����,@��6���\���:>���?/7�?�1?[/#��ԭ��@>�ŋ>�7�=\%e=���.��h/罦�0>��L������=i�TDW=?�
<�8
�wR�h��-���S��j�ܿ�NQ��f]�ďݾ�2��(u	�����_Ӽ�d2���ξ�Y�c���jLV��J<�g=@�$��"���&��p���x��? T�?)�;��.n��3h�i�I���齉m�>�s���ݾ�m�=��QF �v̆�Z_'�e)8��I���a�Αz��f�>ؓ �ӏ��%�l��@-���Z;�om>��$?&�ҾE�̾�%�%�2=�e@>�v=����PQ���ԝ�R�A�G}M?y�*?l�̾l���"�^;O>y�?0/�>f@=>ܓ��5��e�5>Q�?�/?�ᚽ�ܒ�^���E��<6w�?��?�<P?����!��̾���X�>��?��>�|��Ӝ��V���O�>A�X?��>�S`�KO�������>9�M?��a����=�?f�>��q>3ۉ����\6�$�H=��>�>FI�x�ѽ����懽�a>�̂>��J�;��ʶ>��PM�$5��ž���^���>�h���!�>��>by,>���I������|����/?��?X)e?�*?��	���4|
��ח��e?01�>��s>hF����>���>�����i�lG����(?'��?���?��G?o�qXٿ�����ž�מ���=A��=�>�N��a->C�4���;�8���*>�˰>�>>�S�>X�>|/i>�?>���OQ)��㳿zi���cP�$[:��j,�����k�'��b���:Y�4N��US>�ؽ�9�ѐ��)P���>;b[D�^E>���>�6�>}�>�iG>��6>dGs�,*Ѿ|Xt�>^��h��HG���Ҿ��־c��� Y��mW��-O��-���{
����>��y=��=��>_w���=��>��=`��=$f\>53>�>(��=�V:>>�.>�l�>w}�=-u��S>+h���o�1l8��P	�rǽC�6?	�ľ�Jо�$�3�"��(A���>��J?)g�=���PL���ˆ���?e���[˾p�{��5K���>�h�>3��=�S��q�=\�A��g߽�>X��>mF���<���P��Yg��2h~==��>(&�c?ĒB?��7?xF�?"D,>���!c?�x?P�?���>D�w�C�}����: �K?
�7?��p?��&?��J=#2Խ�����Y>��h=�w�=X��<�׎�%��=�G�z`�=�����`=�p�F@&;c��=$�>R�:>��[>\&�>�K8?�>4�>?s&�NN,��C������==j��>���>��>�S�>3��>�'>��=� ��f���#i�>|�>V�M�r�QuH=Ӆ�>��>>|6?ȭ:?.�r��[���K����<A�>��?�)?�S�>�� >��⽯�	�Ơӿ"+$�!�����}��5��C��kj�ݣ;�|$�h�꽘�<��Z>j�>J�h>��=>F�$>� 4>2�>��M>*�=T�=&,���û!�"�=�=6D��Դ�:��I���A;z�%�W����{�}9W��T��/�[�q"�Ĭ?#<?�e�^�����Ͼ�ļ����>���>58	?'�?�8>���VqZ��x)� ��lD?��h?��>~.%���=�;��]����>^�>��c=
(��G~7�oY(����=Z�>��
?���>1vʽ�"U�7�O���S�>݂V>1����?Жx?=��*��;��A��g��_��#ڢ>L�ְ�=�>�*�k���HAо��ξ8�=��>ͫ>���?�<>(1�����sݢ�ɤ�����7־�$�>{�>�~?>�}=���!;�ԇ�)֛��]�zpD=�wL>Ka�>$�?b��>n�I?�?�(�>i۽���>/�<�O�>F�>��f>r�>ۻ�>D�>�)E>�ȃ=ɴ��n�h��v�]<�W�=��c_>M�>�p��k�=�>��ƽX���+R#����=������F�=j*�>��>��>�%N?�S�YЦ�5a=*�b�(;�>�1�>��߼�㦾���L�2��׆���?�m2?.�>Hnq>��
�m32�e��� k'�
�?��?\�>�~������`��3������=.�*>f�����C�̾9	�=[����>��'>aI�>yT?H�a?!I.?�ڟ=
��pA��	9H�-�����>�!�>��?#|>���ײ:�k6[��&G��X�I��<��d�L�<�>��=�U>�_�=kT�=;�>���=V��ؠ�=^�p��D�>f+?�0?L��>�Mo=KE����y�@?��`�k�������N�`z�={6_>������>��^�j�\�g�����9�$��>|T�?�?�T?�l���ν�Vj>
1>E��=x]O=2��#g�����`M	>�2�=�tS�����o =�gj>/6�>��T�ɾ������:]����[���Y��0���˾�b�������Y��M�R��+��9q��ʾ��1�L!�<?J3�bKؾ��վ!ֵ��$�?WY�?@�+>�f����{�U*��6��_!�>�Y������~���笾$�̾࠾@ <�g{��R�;��EdM�GU>�<f����8�Y�]����<�>!@?{�����E�V��'���>�8(>a�ؾ����_փ�$ ?�8?i����ˬ��)ȽL�9>X�?]� ?���>�"Q�ÿ�T�>W{+?e�D?A��=����B��>j�?g�?�@? j���s��d!���0�U+=��q?�=?I�+�N��Ž~��O�=�?�\$?�T��0˞�[(��hm>8C?���U�\>��>�ש>7o�=X���@[1�F�"���
����=�d]�YN��&6��"���G�=��>��>��u�C缾K�>���mOM���F�M ����0�y<�?���>�(k>Ĕ>ŀ'�\.��ǉ�����&M?���?�S?;8?�2��f�V������=g��>Z�>�D�=�>	�
��>���>�f�Xq�c��?�!�?~��?�bZ?x�k�S�ſ�H��K�A�Vm�r:+�r�*>a�>=b3��=u>��Q_�=L`�>l> ?u>�:x>j�9>lp>�G�>�8���.,��w��Ǒ���|����_�&�-���7�������?C��������6>U�&:cH�=5���V���,¤���H�`�=f�#?H��>e�?OV�=��<��	��gݾ����Л�Y���Fڤ��G�A�𕾉V��oo ���%��;���#�C�?�>���>�D�>Mpn>Ybc>L�>�����>��>��>�"�>��>W�>č�>|�?�@>�<=�>�>��+��<
�q)���i>�jS?s�(!��a@���<��&?��9�>��?����=7D�J<���v��	�>JS>�ǐ������+=��B>ި�>w�=�D����<_��=�5��������]>b>
���W<<����ǽ���>;\�X2?5?�y?[(�?W�>���� ?�H,?�Z�>0�>��1?f���D�F=i�<?�F?~�?��;?�%W>*��)h��4�ԧ��{w>2NS���L>�>:=-���[��q����=�0;>>CR=���< �$<x:F>|>�>a�?c��>X?�SP>�y��h������=�R>O7B?;�?xg�>ҕ.>;��>�U?��i>������Æ�>�I�<�P4���H�)p�<�7�>aL�>k*H?m�)?���=�����=�M<>T��=�l>�+I?�3�>���>Y��=u�����C�ɾ�þɧ=h�C�R�4-z�����-��f�^���i��jV��e,>>�>�yg>���>	�>ΐ�>}�>�D�= Լ���=���D�&��.M=��=NE�<��=����ƛ��H�_���>����?��IP��lN����/?ȇ�>��}=)<>Ž��7�o�ץ���d>�?�S2?nV?"��>/������)�;��/�*I?��?&G?NF/�h	A=��`��9|h>{f�>��*>����`b��������h��>�[6?��>��������W�r0���W�>�p�=�� �F�?�6i?Wз���=v�8�-�s�,��V�i>����B�S�v��(�_�*ʾV�ԾG|��Ё�>�>cص?�H��W�>9�����¿F��5��|o�����	?-��>-:��f� ���9�&f(�+㱾�ľ�"�h��=���>cf'?I�*?9�i?�\�>�0�>?���?+�=ֵ�>]��>��?^��>���>穚>�a�>�}�=+���฽]4���-�<\ȼoR>�iy>�1>�!d<C=JA�=9�Y=R�;��3�~=<ų;�ߜ<"/�=%�]>2;�=�?�>�\:?\wi��G�T�_��E����u���>V��>�ڸ�+� >q9J��>��_;�>��_?�{�>�p>lT����H�׍D�_3.> �> q�>d~�>��P<B�C>r֎�;��1��7�Ͻ^'��� M�Em~�+�����Q�<=���>��~>��r?�>?��?�Ru�Ġ�޶|��	R�����O�=mU�>��b>/�=�7��6d�#�t���W��p&�L.<�M������7��>+��>}O�>�VL=p�B���7����X�м��%�K?=��p>��x>��
?[R�>�>v��A�8K?���F�^���R�ƾ�l����>_�7>��нB	?���s�)����C�`��>�%�?o`�?rf?�27�=����D[>O�L>�u>�CD�FD�	����<~��^G>&��=$�t��ь��D��P>�}>&���&��X�޾I'���̿�����4�vZ���3׾/���\Ҿ�p۽�®�%z�MZ��D�=�O��M��.���\��XoW��g�|x�H=|?\Ln?�4m���������p���;T�2>�qӾp�����q��j��p�!���ƾ,��c�⾛���'�o��>,׽���������������>T�4?J�ƾ͵ʾ˄�!�ʼާd=҃�=�{ھv���Қ�)-]��QB?tQ1?C�괾�������=c��>���>��=>v�w��߼)پ>��;?%�9?�=�,����o�%:D<��?�l�?*�%?�=��&��P �_j���f�>�M?ac?�g��/b��i�Žg >�?���>�, �k��mP�*��=f�H?�*˽	.<>���>���=܉E��w��:�������}!���>F&�����G��+����h�>��<�������K�>���mOM���F�M ����0�y<�?���>�(k>Ĕ>ŀ'�\.��ǉ�����&M?���?�S?;8?�2��f�V������=g��>Z�>�D�=�>	�
��>���>�f�Xq�c��?�!�?~��?�bZ?x�k�S�ſ�H��K�A�Vm�r:+�r�*>a�>=b3��=u>��Q_�=L`�>l> ?u>�:x>j�9>lp>�G�>�8���.,��w��Ǒ���|����_�&�-���7�������?C��������6>U�&:cH�=5���V���,¤���H�`�=f�#?H��>e�?OV�=��<��	��gݾ����Л�Y���Fڤ��G�A�𕾉V��oo ���%��;���#�C�?�>���>�D�>Mpn>Ybc>L�>�����>��>��>�"�>��>W�>č�>|�?�@>�<=�>�>��+��<
�q)���i>�jS?s�(!��a@���<��&?��9�>��?����=7D�J<���v��	�>JS>�ǐ������+=��B>ި�>w�=�D����<_��=�5��������]>b>
���W<<����ǽ���>;\�X2?5?�y?[(�?W�>���� ?�H,?�Z�>0�>��1?f���D�F=i�<?�F?~�?��;?�%W>*��)h��4�ԧ��{w>2NS���L>�>:=-���[��q����=�0;>>CR=���< �$<x:F>|>�>a�?c��>X?�SP>�y��h������=�R>O7B?;�?xg�>ҕ.>;��>�U?��i>������Æ�>�I�<�P4���H�)p�<�7�>aL�>k*H?m�)?���=�����=�M<>T��=�l>�+I?�3�>���>Y��=u�����C�ɾ�þɧ=h�C�R�4-z�����-��f�^���i��jV��e,>>�>�yg>���>	�>ΐ�>}�>�D�= Լ���=���D�&��.M=��=NE�<��=����ƛ��H�_���>����?��IP��lN����/?ȇ�>��}=)<>Ž��7�o�ץ���d>�?�S2?nV?"��>/������)�;��/�*I?��?&G?NF/�h	A=��`��9|h>{f�>��*>����`b��������h��>�[6?��>��������W�r0���W�>�p�=�� �F�?�6i?Wз���=v�8�-�s�,��V�i>����B�S�v��(�_�*ʾV�ԾG|��Ё�>�>cص?�H��W�>9�����¿F��5��|o�����	?-��>-:��f� ���9�&f(�+㱾�ľ�"�h��=���>cf'?I�*?9�i?�\�>�0�>?���?+�=ֵ�>]��>��?^��>���>穚>�a�>�}�=+���฽]4���-�<\ȼoR>�iy>�1>�!d<C=JA�=9�Y=R�;��3�~=<ų;�ߜ<"/�=%�]>2;�=�?�>�\:?\wi��G�T�_��E����u���>V��>�ڸ�+� >q9J��>��_;�>��_?�{�>�p>lT����H�׍D�_3.> �> q�>d~�>��P<B�C>r֎�;��1��7�Ͻ^'��� M�Em~�+�����Q�<=���>��~>��r?�>?��?�Ru�Ġ�޶|��	R�����O�=mU�>��b>/�=�7��6d�#�t���W��p&�L.<�M������7��>+��>}O�>�VL=p�B���7����X�м��%�K?=��p>��x>��
?[R�>�>v��A�8K?���F�^���R�ƾ�l����>_�7>��нB	?���s�)����C�`��>�%�?o`�?rf?�27�=����D[>O�L>�u>�CD�FD�	����<~��^G>&��=$�t��ь��D��P>�}>&���&��X�޾I'���̿�����4�vZ���3׾/���\Ҿ�p۽�®�%z�MZ��D�=�O��M��.���\��XoW��g�|x�H=|?\Ln?�4m���������p���;T�2>�qӾp�����q��j��p�!���ƾ,��c�⾛���'�o��>,׽���������������>T�4?J�ƾ͵ʾ˄�!�ʼާd=҃�=�{ھv���Қ�)-]��QB?tQ1?C�괾�������=c��>���>��=>v�w��߼)پ>��;?%�9?�=�,����o�%:D<��?�l�?*�%?�=��&��P �_j���f�>�M?ac?�g��/b��i�Žg >�?���>�, �k��mP�*��=f�H?�*˽	.<>���>���=܉E��w��:�������}!���>F&�����G��+����h�>��<�������K�>���mOM���F�M ����0�y<�?���>�(k>Ĕ>ŀ'�\.��ǉ�����&M?���?�S?;8?�2��f�V������=g��>Z�>�D�=�>	�
��>���>�f�Xq�c��?�!�?~��?�bZ?x�k�S�ſ�H��K�A�Vm�r:+�r�*>a�>=b3��=u>��Q_�=L`�>l> ?u>�:x>j�9>lp>�G�>�8���.,��w��Ǒ���|����_�&�-���7�������?C��������6>U�&:cH�=5���V���,¤���H�`�=f�#?H��>e�?OV�=��<��	��gݾ����Л�Y���Fڤ��G�A�𕾉V��oo ���%��;���#�C�?�>���>�D�>Mpn>Ybc>L�>�����>��>��>�"�>��>W�>č�>|�?�@>�<=�>�>��+��<
�q)���i>�jS?s�(!��a@���<��&?��9�>��?����=7D�J<���v��	�>JS>�ǐ������+=��B>ި�>w�=�D����<_��=�5��������]>b>
���W<<����ǽ���>;\�X2?5?�y?[(�?W�>���� ?�H,?�Z�>0�>��1?f���D�F=i�<?�F?~�?��;?�%W>*��)h��4�ԧ��{w>2NS���L>�>:=-���[��q����=�0;>>CR=���< �$<x:F>|>�>a�?c��>X?�SP>�y��h������=�R>O7B?;�?xg�>ҕ.>;��>�U?��i>������Æ�>�I�<�P4���H�)p�<�7�>aL�>k*H?m�)?���=�����=�M<>T��=�l>�+I?�3�>���>Y��=u�����C�ɾ�þɧ=h�C�R�4-z�����-��f�^���i��jV��e,>>�>�yg>���>	�>ΐ�>}�>�D�= Լ���=���D�&��.M=��=NE�<��=����ƛ��H�_���>����?��IP��lN����/?ȇ�>��}=)<>Ž��7�o�ץ���d>�?�S2?nV?"��>/������)�;��/�*I?��?&G?NF/�h	A=��`��9|h>{f�>��*>����`b��������h��>�[6?��>��������W�r0���W�>�p�=�� �F�?�6i?Wз���=v�8�-�s�,��V�i>����B�S�v��(�_�*ʾV�ԾG|��Ё�>�>cص?�H��W�>9�����¿F��5��|o�����	?-��>-:��f� ���9�&f(�+㱾�ľ�"�h��=���>cf'?I�*?9�i?�\�>�0�>?���?+�=ֵ�>]��>��?^��>���>穚>�a�>�}�=+���฽]4���-�<\ȼoR>�iy>�1>�!d<C=JA�=9�Y=R�;��3�~=<ų;�ߜ<"/�=%�]>2;�=�?�>�\:?\wi��G�T�_��E����u���>V��>�ڸ�+� >q9J��>��_;�>��_?�{�>�p>lT����H�׍D�_3.> �> q�>d~�>��P<B�C>r֎�;��1��7�Ͻ^'��� M�Em~�+�����Q�<=���>��~>��r?�>?��?�Ru�Ġ�޶|��	R�����O�=mU�>��b>/�=�7��6d�#�t���W��p&�L.<�M������7��>+��>}O�>�VL=p�B���7����X�м��%�K?=��p>��x>��
?[R�>�>v��A�8K?���F�^���R�ƾ�l����>_�7>��нB	?���s�)����C�`��>�%�?o`�?rf?�27�=����D[>O�L>�u>�CD�FD�	����<~��^G>&��=$�t��ь��D��P>�}>&���&��X�޾I'���̿�����4�vZ���3׾/���\Ҿ�p۽�®�%z�MZ��D�=�O��M��.���\��XoW��g�|x�H=|?\Ln?�4m���������p���;T�2>�qӾp�����q��j��p�!���ƾ,��c�⾛���'�o��>,׽���������������>T�4?J�ƾ͵ʾ˄�!�ʼާd=҃�=�{ھv���Қ�)-]��QB?tQ1?C�괾�������=c��>���>��=>v�w��߼)پ>��;?%�9?�=�,����o�%:D<��?�l�?*�%?�=��&��P �_j���f�>�M?ac?�g��/b��i�Žg >�?���>�, �k��mP�*��=f�H?�*˽	.<>���>���=܉E��w��:�������}!���>F&�����G��+����h�>��<��������ܵ�GpT��7���>��G���x�����<�>�	��Z%���>�)�>i�d��*���q���X�=xuk?��?�]?!"?7?����վg�|<��d>���>��l�ξi��>���>�@"�'U������?l��?��?"�k?%�w��x��氒�3���5O��>0m=�BH>�q3��Q�=��=��/>:��=u��=ѣ�>C�$=�-=>C�U>�Z>oP�>�t��ls �[��9`��_,��C��$��=I������M����ĩ�k~žo=8�T���eT4���K�ّ����`>a;پ���;K?�>�>D�}>�ќ>��f��-��0h�w�D�Ӿ|Qپ�ݾޞ{������x�t���x��#��>��=�>j2?9�v=y̒=	O�>ơ�=F�=���>�cO>k��=�$�=ν]�I�=ɀ%>
[0>���=<P�>G�^�}`����+�Q"�%l >'fc?��
���1�vo�,����T
���?8�^?�V�<��L��(��2]����>&��<�g���:l�i�_;>4J�=�R�=��N>����о_���c��=/+�>�O�>�G]>�.���ؽ�`�����?���zʓ>�?osH?���?��?Da?�~�>r�>��j��>���>}�R>�K?�`?�=?"O�>׃�=��о���=�{~>�Ѡ�p��^�
<N���w���=��V>,�j>�B��g2<]=s=�e-������5=g�?x'?Ew�>��>��ҽ��2��Ld�0qn���>��5>9@>>">Ӽ�>%��>��?6>pK��/���+C���t ?xS�>�o�;?��=ÿ=�=��^?�SY?��;45ʾ��2��� �I6�>4X?�?,�>�c�>[�6����<�Ϳ�"�)A#��q���n���<��Q�g�������(y �T����&%>��j>L}>��b>n�.>9T1>���>�W>F�=X��=c؄;�I=p~]����<t�̼ ב;�����<P�d<�-ǽ~��$�����3�F闽�<�����>w?�;ż5㚽]�*�����꺾*ޜ>���>��?�%�>۸>�����e�>iC�޽�S�>��V?R��>��ս��{=�Α�&=N*�>6��>.3>���j������G���>ݩ1?�g�>���pj��k��k��PB�>���=��/��O�?%c?��N��A��FG�,���+>ܕ2�z6�Pr�� ���O�о/���a��)<$�?�O�?�$���YA�%������[ ��S%4�$�e>��=�F�>��P��M���ƾ��澃���� P��f>O��>�->7�>um8?��N?]$~?��.?�s�>6T޾�� ?k�->,�>��>�h?��?�t�>�5�>��>�a��r\��ȩ�uþ#(�<��=9�=/[>� o>��b�0��<ȶ�;��=Wڋ:����E�<p>�=�wf=`�'=�X=�>?%�=?���<Qڋ��-���;�vZ��<>�v�>��s=�>����;n+m>���>�??9��>�{=�A��D�*��a�=v鼩�?`E'?؝�>�',>�>՛B�Œ� >8?[�>ղy�8_꾹"�M7׽B[�>�G>�b>[1~>w�?��g?�F?��s���"�5m���uU��ψ�w�=o�>�}�>�Q>>NgV���#�لK��T�Z&,��2����̟=�\�=�>�Z�>0�K=���<�#<�g�w�Q=�p�=x(�;[�e>��>�Z	?�!�>��T=��������?BB��^C/�L���?�R���(���(>�r*><�4�G�?�;�=���B���:3U���>��?���?��?�1A��1N��.�>A÷>֠�=􇼭�^�r����;�U)/>�ܞ=����i�I�=A,x>ǆ>"��1A��b/�կܽYѸ�<��F'�a���X������x��Qh���;��bl��9齝���y�tJS��߂�Q�z������A�l?��g?FO[>��=�x=��c�$�о|>Z�½e��~���1�H=�#>�{���XNľS��D���,�49����V>�!)� �i���e��I<�`����b7>��0?׾������D��>�>�ޅ��	�����FdȽ��]?3�2?�̾g'�,�G��v>=�2?��!?Q?�>�P������Vt�>1� ?�t:?��>-O��-��n��[�?46�?r�4?Iy����	�E���h�����>qj+?KM+?㱷�o��X?=��?�nL?�\�>L��9���.�c�>�#�?�U�^T>-�?� �>��뽲���|��tB��.2�<P7N>P�B���Ү��-½�94<6��>b]>������\Ǜ>&�����m���n��X��D��s�>�?�V"�׷M����k�l?|lg������a��>���LD3??"�?�oq?��?.��3��$>I�%�>}��>�,ǽ�.��G5>�M�>'���z{�p��?��?���?Ŕ3?I�\�'�濾���	A���r��#w�>%>��">��ս+��=M��:��:G���"�=���>�5�>���> �7>��>j�">����|'�OB��4������e4���!�$XԽ����觾d��郾N��{�<ԟ/�T\̽mq��	��f,��!덾��=Ʃ%?+%�>��>w��>��>�M��/�����žU,��٦ ��H����	�1�����e����;�;e��:۽`=��jſ>�`/=XN>�?K�J=,��=Ns�>(^a>)��<,a>]h>/�v<�T>I
l>��=�ɇ��,>��>�~>щr�������:�α��x=�~"?z�#��ֺ�i5<�{��ɾ���>�?���=3�0��a��$�}�q<�>V�y>f��=��h%�=���=Y�Y>�m�>�A�>�H}��s�L�	��˫���v>\�>.W=}�־Mӽ�ݔ<�a�>`���c�>/Z
?j�6?x��?0�-?$�(���>��>Z�>qxo�+��>N[5>�k�>��?�v(?�"�>;��>�	�=$��l��=E>>?�3�s�J�l�}��g�o��ڜ�=X0�=Fq�;\��	�<�h3>QC�<Ý����=�=��?:�4?.>?+?�';)y ���o�~X���(�>���>Ȣ�>�Xa>��"?�&�>�?���>A��=kr��ߞ����>�O>%x����ש�=�[�="�J>#gy?�~o?6�K�ѩ�
��*;� h�>�%?<?o�?Z�2>��u�M��A�ߪ.�P�	�N�>�ؘ�q�+�V��"��V\����<o4�F����>��>��t>)�=�S�=�q�=Ȣ�>�Is> ]C��/>�p���>�aҡ�s�~<�#��PMQ�'��=I�ּ�l��#�e�H�J�'���?����Y��������>��?I̙��U���.l�Q�� ��>�>7�>SM�><�L>���=��-�qi����=�Q�=-�-?T�s?��?�b	��1�<����'>���>�r�>�zn>���=0Tl��l��CF]>ڢ=W�d?-�E?Xd>��.9��p���[��>+��=K#�����?�n?����8��A�Sd�l��h=�u=�
V���H�͏�Z)�~����I�u��"�=�_�>(:�?Y���;�=)�ھ!��ʇ��D���ָ=M)>��>��>6��=�7��/����l��[���$�۵�<��>�d�>�H?aP?w�H?!�6?\-�>L�ʾ���>��|>���>�a�>,�(?�?u �>w�>3eQ>�b�;�������U��u��o&�=A�9>�ن>�=\>�=����h�>��'<�g��=�CW==򼽋#4���=� �=mw�>�?M�1?��>�6�Q�k���s�<*�)SA>(�?+�k>`���jɾU�>���>��B?wq??�=6��A��*���l�*?e�??�j>E�C=��=�e��?�����>w�m>����f���6��a#W�\����>�l>�+�>"�~?L�c?�f??��K�ަ%�7ݍ��H]�Z�<�/>�!�>��>3wo>�к��/���C��BO��<0�-����:���=E,
>|%J=���=�K-=�nO=�۟<��q�*�=��=,�]<G��>x"�>)?�y�>��>r>��ؠ���G?������nw���H��25���H�}L)>G�>��?���nUf��	���SH��Ι>w�?X��?=�`?C��F���">6�c>��>�E<����j3�:�ν��=b E=ȱ��ƎѾ{g�?>T>�~��sž�D���P�#�Ͽ:0�����"z� -�<R����������׾�,ξR�>2�!�zK���>�^(��� �~�T�Z5���?��?vݽ����dN�#��1�����T���H*��GȾ�J���ϕ��π�
��ҷžq����4��4���=u�=�~�|��H-���!����=rJC?����P����4�w=�>E3��_Lk=�[ �w%���v��sv>�IEC?�?g-����wI����>Hǝ>�y�>�f�>հ�{�l����>�c?��?�Z���T���c��#����Z�?���?�??�n�����,Ǿ��ҽSg�>MJS?��]?�̫�ꚞ�kN> ��>=\W?F��>H~��� ���M���?�v�?9c�0�X�n��>b�N>F&��*M��&��Ƞ�����QSj>uT˽W1���=��)��f@=?q�>�H%>��վ����ܵ�GpT��7���>��G���x�����<�>�	��Z%���>�)�>i�d��*���q���X�=xuk?��?�]?!"?7?����վg�|<��d>���>��l�ξi��>���>�@"�'U������?l��?��?"�k?%�w��x��氒�3���5O��>0m=�BH>�q3��Q�=��=��/>:��=u��=ѣ�>C�$=�-=>C�U>�Z>oP�>�t��ls �[��9`��_,��C��$��=I������M����ĩ�k~žo=8�T���eT4���K�ّ����`>a;پ���;K?�>�>D�}>�ќ>��f��-��0h�w�D�Ӿ|Qپ�ݾޞ{������x�t���x��#��>��=�>j2?9�v=y̒=	O�>ơ�=F�=���>�cO>k��=�$�=ν]�I�=ɀ%>
[0>���=<P�>G�^�}`����+�Q"�%l >'fc?��
���1�vo�,����T
���?8�^?�V�<��L��(��2]����>&��<�g���:l�i�_;>4J�=�R�=��N>����о_���c��=/+�>�O�>�G]>�.���ؽ�`�����?���zʓ>�?osH?���?��?Da?�~�>r�>��j��>���>}�R>�K?�`?�=?"O�>׃�=��о���=�{~>�Ѡ�p��^�
<N���w���=��V>,�j>�B��g2<]=s=�e-������5=g�?x'?Ew�>��>��ҽ��2��Ld�0qn���>��5>9@>>">Ӽ�>%��>��?6>pK��/���+C���t ?xS�>�o�;?��=ÿ=�=��^?�SY?��;45ʾ��2��� �I6�>4X?�?,�>�c�>[�6����<�Ϳ�"�)A#��q���n���<��Q�g�������(y �T����&%>��j>L}>��b>n�.>9T1>���>�W>F�=X��=c؄;�I=p~]����<t�̼ ב;�����<P�d<�-ǽ~��$�����3�F闽�<�����>w?�;ż5㚽]�*�����꺾*ޜ>���>��?�%�>۸>�����e�>iC�޽�S�>��V?R��>��ս��{=�Α�&=N*�>6��>.3>���j������G���>ݩ1?�g�>���pj��k��k��PB�>���=��/��O�?%c?��N��A��FG�,���+>ܕ2�z6�Pr�� ���O�о/���a��)<$�?�O�?�$���YA�%������[ ��S%4�$�e>��=�F�>��P��M���ƾ��澃���� P��f>O��>�->7�>um8?��N?]$~?��.?�s�>6T޾�� ?k�->,�>��>�h?��?�t�>�5�>��>�a��r\��ȩ�uþ#(�<��=9�=/[>� o>��b�0��<ȶ�;��=Wڋ:����E�<p>�=�wf=`�'=�X=�>?%�=?���<Qڋ��-���;�vZ��<>�v�>��s=�>����;n+m>���>�??9��>�{=�A��D�*��a�=v鼩�?`E'?؝�>�',>�>՛B�Œ� >8?[�>ղy�8_꾹"�M7׽B[�>�G>�b>[1~>w�?��g?�F?��s���"�5m���uU��ψ�w�=o�>�}�>�Q>>NgV���#�لK��T�Z&,��2����̟=�\�=�>�Z�>0�K=���<�#<�g�w�Q=�p�=x(�;[�e>��>�Z	?�!�>��T=��������?BB��^C/�L���?�R���(���(>�r*><�4�G�?�;�=���B���:3U���>��?���?��?�1A��1N��.�>A÷>֠�=􇼭�^�r����;�U)/>�ܞ=����i�I�=A,x>ǆ>"��1A��b/�կܽYѸ�<��F'�a���X������x��Qh���;��bl��9齝���y�tJS��߂�Q�z������A�l?��g?FO[>��=�x=��c�$�о|>Z�½e��~���1�H=�#>�{���XNľS��D���,�49����V>�!)� �i���e��I<�`����b7>��0?׾������D��>�>�ޅ��	�����FdȽ��]?3�2?�̾g'�,�G��v>=�2?��!?Q?�>�P������Vt�>1� ?�t:?��>-O��-��n��[�?46�?r�4?Iy����	�E���h�����>qj+?KM+?㱷�o��X?=��?�nL?�\�>L��9���.�c�>�#�?�U�^T>-�?� �>��뽲���|��tB��.2�<P7N>P�B���Ү��-½�94<6��>b]>������'�>��羯=M�!H�q��D�6��<*� ?����>9�d>؂	>�N(�n��-剿�����I?0�?��S?�7?������뾙����;�=0��>X�>��=�D��
�>��>��྾�p������?���?wM�?�U?�m���꿷	���Į�׮���Q>��`>J��>LIӽ��X=3T�=ͨ=��ν�S�<q�>^ȇ>��Q>��W><�K>��c>�ً��+/����]���%"�']������g�u��E栾iC�g
���ߺ�PQ</��=~;��_���ܻ��<l�t�� �z�?��#?�N�>�B�>P�>�����xt�|z��i�?��;%���@�����~�C����i�Ǟ!���&������>� :f�a>���>j��="�Z=h�>٬%�
K�<uM�>�A�=�-f=y�=�".>�a�>7�=��R�V(<e<n>+�X���X�-@e�U$��&���F?i��/�ž��$�./�x����>��>�/�>U] �¡��F�m�޴>�D>�b4����R�*�{��=���>]>�q>3q!<;e辺+��= ��>�ڿ<���b�ԿA������>�C���ʹ>���>n?]h�?w�.?�ؾ���>*.?��>���=���=�<ϋ�>K�<?�I�?�U?�?	�T�g�:��~">�!���Ǯ����;�E>��=g��Y%�=C�R=+��׾<�O�<�X/>t���`j[=��=�7�=շ?�:?Y?~E�>^�ݾ0@��Gc�]�r���>�3=! �=3>z�?H��>{��>��>��=����x��Y2�>3׽>Zyi���b��;���3�-<J�?�?v���־̜����?=�a�>��D?��]?J9?er��l�ž�z�T?�w�&�MN�`Ő=)=�)3=lg�A����7l� ����
��	��o�>���>)��>I�*>.�g>(&b>!F�>��{>ݞl��=��=����&��	>_�A=�񺼣��;��~<j^�� ʽ�S���!����]X��L����?T�?��y��= ��2ۼ�_��i�꾰#�>�?��	?��>F��bδ�wf6��C��	B�̰�>+Bg?u�>��d���L�{S=�ko>]��>�/�>T
�>����ݾt�þ<d>���>��>9[#>/�(bV��^������>�1=�����q�?�.p?�ԏ������� �g[�p���a��=�Hj<]oA�����E���=�p��0�龒Ќ��$>�:�>q�?|ĺ� Mݽr}о��]ʬ�	��z�=N�0�UԷ>�&	?�>�/�����;=yM�}ؗ�V@=�I>�&�=�/<?��e?�N?��;?���>��쾢��>�(�>B ?���>���>+Y?���>�˱>�K�>��=r�C<C9*�kn���c���o�<,�=��>N��>�ch=�Kݼm6<>��H=�O2�}%�^��;�!��Z�
�J�>�e>'�<>Cy?ԝ3?+OM<���%⁾6�M�\Y��m��> ��>:�@<�
�����qX�>���>sP3?��?xt�>!�5C�/<��3�p�ۆ�>�$7?Ӽ�>���>kX;�!5��*���H=>-�>���rtD��@���d����<����RM�=�C�>r�>��z?�Ht?@9?�[�%��Q����;}�G9H��Lh>��>�
2?���>=ݾ�J	�}���5�c�'�G*�,��|=�J=�T=���=��X>t�.>C��=^쮽x�/�����F����>!:�>A�?��d>�u�=Tt��Vd ���J?>���w��ha���jѾ�o)�Y�>x�C>.½?�-�&
��%y���<�T��>t��?R��?��b?$�H��%��[>��C>g}>κ�<|�3�|3������Q7>�7�=�]u��Z����c<.]>�j>`-��]žytݾT�?��&ǿ�tl��J)���d�.�ߧ��wo�>㭾��������m���S�43�=�Y��F��
پ�-i�/᯾�q�?9�?^ͼ��ϽQ����$��VǾF��>NF���z;��y�\���T�6�+!��]X��*��q�2�ֺ�?о��}>ZC>�d��)=��+���ϾF�>HLm?؃��0NM��T��t�>�W�>-�>` �Ҹ��Ӭ��4��<[�?9�?�����B���m�?Q?7��>Пc<��t<�t3?hQ?���>�3�����,���қ!��R�?=k�?/#�>}�ۻ�T�������>:�H>.D?x�?��׾�e.>�[?��>�v�=��h��֥��ȝV?�C�?#�*��H�=2L"?9S7>�Yh��F�=�r��4��� i�=�|>Uϫ������_I�wݿ��o�=�>Vt>��"�Z���ܵ�GpT��7���>��G���x�����<�>�	��Z%���>�)�>i�d��*���q���X�=xuk?��?�]?!"?7?����վg�|<��d>���>��l�ξi��>���>�@"�'U������?l��?��?"�k?%�w��x��氒�3���5O��>0m=�BH>�q3��Q�=��=��/>:��=u��=ѣ�>C�$=�-=>C�U>�Z>oP�>�t��ls �[��9`��_,��C��$��=I������M����ĩ�k~žo=8�T���eT4���K�ّ����`>a;پ���;K?�>�>D�}>�ќ>��f��-��0h�w�D�Ӿ|Qپ�ݾޞ{������x�t���x��#��>��=�>j2?9�v=y̒=	O�>ơ�=F�=���>�cO>k��=�$�=ν]�I�=ɀ%>
[0>���=<P�>G�^�}`����+�Q"�%l >'fc?��
���1�vo�,����T
���?8�^?�V�<��L��(��2]����>&��<�g���:l�i�_;>4J�=�R�=��N>����о_���c��=/+�>�O�>�G]>�.���ؽ�`�����?���zʓ>�?osH?���?��?Da?�~�>r�>��j��>���>}�R>�K?�`?�=?"O�>׃�=��о���=�{~>�Ѡ�p��^�
<N���w���=��V>,�j>�B��g2<]=s=�e-������5=g�?x'?Ew�>��>��ҽ��2��Ld�0qn���>��5>9@>>">Ӽ�>%��>��?6>pK��/���+C���t ?xS�>�o�;?��=ÿ=�=��^?�SY?��;45ʾ��2��� �I6�>4X?�?,�>�c�>[�6����<�Ϳ�"�)A#��q���n���<��Q�g�������(y �T����&%>��j>L}>��b>n�.>9T1>���>�W>F�=X��=c؄;�I=p~]����<t�̼ ב;�����<P�d<�-ǽ~��$�����3�F闽�<�����>w?�;ż5㚽]�*�����꺾*ޜ>���>��?�%�>۸>�����e�>iC�޽�S�>��V?R��>��ս��{=�Α�&=N*�>6��>.3>���j������G���>ݩ1?�g�>���pj��k��k��PB�>���=��/��O�?%c?��N��A��FG�,���+>ܕ2�z6�Pr�� ���O�о/���a��)<$�?�O�?�$���YA�%������[ ��S%4�$�e>��=�F�>��P��M���ƾ��澃���� P��f>O��>�->7�>um8?��N?]$~?��.?�s�>6T޾�� ?k�->,�>��>�h?��?�t�>�5�>��>�a��r\��ȩ�uþ#(�<��=9�=/[>� o>��b�0��<ȶ�;��=Wڋ:����E�<p>�=�wf=`�'=�X=�>?%�=?���<Qڋ��-���;�vZ��<>�v�>��s=�>����;n+m>���>�??9��>�{=�A��D�*��a�=v鼩�?`E'?؝�>�',>�>՛B�Œ� >8?[�>ղy�8_꾹"�M7׽B[�>�G>�b>[1~>w�?��g?�F?��s���"�5m���uU��ψ�w�=o�>�}�>�Q>>NgV���#�لK��T�Z&,��2����̟=�\�=�>�Z�>0�K=���<�#<�g�w�Q=�p�=x(�;[�e>��>�Z	?�!�>��T=��������?BB��^C/�L���?�R���(���(>�r*><�4�G�?�;�=���B���:3U���>��?���?��?�1A��1N��.�>A÷>֠�=􇼭�^�r����;�U)/>�ܞ=����i�I�=A,x>ǆ>"��1A��b/�կܽYѸ�<��F'�a���X������x��Qh���;��bl��9齝���y�tJS��߂�Q�z������A�l?��g?FO[>��=�x=��c�$�о|>Z�½e��~���1�H=�#>�{���XNľS��D���,�49����V>�!)� �i���e��I<�`����b7>��0?׾������D��>�>�ޅ��	�����FdȽ��]?3�2?�̾g'�,�G��v>=�2?��!?Q?�>�P������Vt�>1� ?�t:?��>-O��-��n��[�?46�?r�4?Iy����	�E���h�����>qj+?KM+?㱷�o��X?=��?�nL?�\�>L��9���.�c�>�#�?�U�^T>-�?� �>��뽲���|��tB��.2�<P7N>P�B���Ү��-½�94<6��>b]>��������?/�ʾ��tt˾�Yؾ󄎺ȡ�=΃K>������>=/?e��=w}Y��]���¤�B�U�d��?���?&�q?=2?�!�Wr龴+��->e?S��>,���am���E>൬>�	���0f�Ԍ���>���?���?h?A7D��ܿ�J���l���w��f��=�'w���F>`��=��p=�����v����V=K�=r�^>��2>��E>�� >�>�g>⏅��������������W�'���]禽�)��S޾��6��(������Iw��gJ�۪'�񆁾�a�t�ʽ������A>~"?��>��?u�>�[�=�b����3�G*Ծ�VL�hc��@�z>�8����<����:�l���!� �Խbz0�%�S?�n�=׮;%�?��!�Mz�=��<������>w�>	��ʊ>�b�>�;n;��ѽ6>�G=Ex�>]���X����X�0%���=���>�M?;��<>��>������|�>-y?	�(?䝣=�:��(p��q�+��>����E�՗n���	�G�>���>#5����>c���N�ͽ"��=M�B>A�>�m">�� >�c۽-L�~n���>�#ƾ���<G�=y=?/G~?c�:?;(�=�f�>�V>��>#�>яv>ꚜ>�Ǣ>~?��'?%�?6��>��=qY?�6��=0>^� �Jr����4��x?�wcu���[;���,�1=�T�=@�W����=^�=�N��E0<���=���>�]?S�>T�T>�|�\�D�NX�Q;}Q�>�u]�_8�>3��>Tj�>6��>n��>^XW>*D ����5^;F ?��>��x�<܌�D���?_��>�H�?��g?[OY=k��FǇ=�a�=��>�*?.,L?]:�>T	�>���=d�4�˿c��/��o��c����[;��t���n��p����G�u���D=��X>��y>��C>	��=Ll�= z>�n�>v�">7҂=�J�=�_=<��伺н�k��~�G�l>�ɍ=ti2=G��<~]	���V���4<�/Q��$�<����?U�(?��<@xؽ1h���㾸�,�<φ=��5?��$?��?�e�^��	P��#j��m���M�>�_�?S9?�W�x��>����<ƼB>��>�Ys>�'+��l�=��e��t��W?�J?� �>�OŽ˚r��ꐿ��4��*�>�>�;�C�f��?ľ-?FJ��WL.�
M��:Y�>?D�n�i<���y;��G׾��<��8���#�p��;�[<�cI>���>k��?4�۾B�=�qx��*�� ����u��AI>�� =x�>�Ԣ�	'����f�ey���ƾ({�=�8>��?dyB�EZ꽨oG?Q[f?�UV?�?��K?Xnq����>0��:�<��?�[�>��-?��G?��>^S�=�=$6>���1��T�=�3>�:=,��<ɿ�=TI'=}���C�<�����C��
q��(��=CJ=��R<$%�=u�>���>�'?b&��@����<�>}L�=(�>�W�>}�3>̀����-<?w?p�?�^�>�?�<��þ�(�?��N	�>�c�> ?��*?����z���+�|���(<n#t>���D�����X"�Hʾ���=B�>��n>�k�=>6�?��?�?��'>�G{�H������j��^����+?��>�>��3�e}+��y�6s���[Q���!>����=��> f	>ף|>Đ潠a2<j����`��Tٽ�̴=�a�i�}>��?l�?�T�>��^>I����t�-;g?�����羵g���s����=O�=_'��ࢾBm�>�+�<��[�]��������h���b�?|)�?Ki�?�D�=�"��4�>]��>�p�=	��=O��E���m��=��>���>�9��5�����=iy=;Қ>����!�����M���ݿC0E��,P��8��.�Ǿ��� ;;��>���_L�r���8þ%\����7�x�-We�Z����������?|l?퍑��(��I��Q��v�>:�����=SZ��L�s�y�������P�Ͼ*[�i��!����>경f��QDL�>��x<9����<��6?�̾�k����m��=^Z�=Oiѽܸ�񄕿���U�����d?swA?ڞ�(;��b����=�#?�Q?�x	>��fIɼy:�>!%?���>4���ɓ�����=f�?A��?��??7�i�ۗC�M��j�B���?
�?il�>�Wf�y�������?<":?V�>ȩ�Y�{��h���>ڣD?��I��>f>f�>ҁ�>�u���v���T��G�}+>-��;Xj��i��IE�C�=>�f>~�J����X�=?h/���W�G���T�ҽ1m>ˆ�=w��>x���O�>sY�>xe?	�b�S.��%���k�\�?���?�i�?�>0?��+�E1p�1�ʽ�$�g�?�b>a�1>��t� ��>}��>��ƾ�����v����>�W�?m��?���?�R�zѿ=>��i�������>���=/�h>A����_�<���<�=<>���A�=T��>>��>��~>U4>��>Z�>�;��
@!�M���#S���M:��$�r����T����dÏ�����e���� �� �P`�S����i�Rs�,�ɽx����-#�0R?��?K�?���>�� ?J����LY��/O���+>�z��%!� �2�+
�[�1�!>QN�P�O�ҽq*�,�H??�1�����M?��` >g��>R�r=a>5�a>�LN=�3�=>_F>>�[>_ǽW��=˯�o������>k�}��`��ǻd� ����1�s?<1=�H��%?���Ⱦe����F?qg?�΢=��x���C~��߱>��ǽ�Ђ�!}��z�<="Ԃ>q��>�߻=^z�=t<��R���p�:&�=|��>w�����ֻ��&�$Le���<��>#wH��>8>=e>�U1?ȯe?1?C����>yx?|��=���A��>c�>��>e�9?fB?�4?	�>�;Mk��� �=.6>�r�%�<�*�<�^|���i��.��ܤ��J�=��2=Z��=G��=Q�½�K$��b��J>x��>m�=?�?-��>�E�;�3�0B�3�*�>G�>ю>��k>q(�>�+?�x�>�1?>��>BD=�񒾠=ܾr*�>ئ�>��y�����2S�i�:>�6z>87�?y4x?3��=jƾ)�'��ޚ��3�>??�??f-?죙>?=aN��Oܿe^����m��n=�l=I�i� ����잽F���>��2a���<>�4E>sa>8T7>!��=��	>���>�H	>D��=��=@����ٺ��4�)��<�M?;���=%�|=��>%�0>�V��N��X�����V;�f�=��n��r?�a�>i <U>����
��������=�D.><2?��?~#h��.��Bf�Ha�~�;��Q?C�f?��?�Ͼ�9�>b�C=�3
=7�?�x�>�>��9�<F��~��`~���ڇ>V�?t��>���s�v���Y�ITJ���w>��$>�����?��I?�I�"�>���c��f�7��`X�<�Ƃ�m8Ͼ�Q?�	V�7�پ����1����>uc�>If�?~/���ќ��n��io��v���47��r->���q�d>ORB>��L��4|�<�����Z��=�?�?a=���>;IB?�RA?��}?��?]��>4v;��U>=��>$r >��G>g -?���>�j-?ze�>�>���=Mc=��c�=Θ���.>1�c>�n>K�=Z;>m7�j ýdb�=�2�=��;E���^�<3��=3�=�2�=�I�=%~�=��>U�?i�%��k6�Mʼd�J�7�=p�>q�W>���;�vľ� ��	�>v2?#�0?��>�Z���پ_���	n=S�?}!?j?��Z�!^>��	�+����]=�1�>�0�=3��YO�9��� ��zT�='H�>���=�,�>���?�9f?���>�&<����Ә�x�U��b?�������>��>f�?	����j��GR�H�g�A[ �w��>YXd�f�ʼh���k�>-ʇ>eש�
j=;�
>���,��GH���=e'?��>�f?ް�>���=��4L��d?��������$��uڎ��ݤ>��>�*��43?�<V>u^:�%���w�R��K�=�`�?���?�ّ?.�<�6��F�>�g�>���>�$���<�u�>�jp��+�=���>��U�k"��}m>�-�=�-�<�ዽ�O$��0,���4���ӿA?w���Z��m9�m��CV�BIо��;e�x��E��	h���^���֝�9���(g�\a=5uB�H������(x�?���?���P���S�w���R�!>ž!� ?k<�ﾼ[���PT=ʒ��j?���\��/d�y ��o���M���}>����W����\/�u�¾tq��l(>L.�>Z�ھ�멾�9Ͼ�f�>ڙ>��h���	�傱�
ۉ������J?fE?��ʾ�a�Ư<=�F>Xx�>���>���=��DR�ꦖ>��4?�:?\߯����x���=)�?��?��??�O�{�A�7+���y�?
c?K�>D��Yp;oP��$�
?L�9?5��>͵�r0���4����>��Z?h�N��bb>o��>#��>N^�1͓��	 ��ϒ�R����;>SS����f���=�|�=|�>d�x>��[�b��:� ?�R�a�F����<����煽s�&�>��E�&L >���>��Z>���t^��oA�� ܍��r?n[�?�t?�-?�h4���g��#�=�I�=E�>?-��>iV-�P��=C�+>�E�>�^����_��A �>�6�?��@��?�g��ӿϽ��`+���K����=��>�Fo>�4�!]�=�w�<?�<�=�d->�c�>[�V>9!h>"�>>��9>B<'>�l����!��B������N<�<!���߾�J-�.B��င�>���������ý������B�3�>p��=�>�"$��kg0>�=?��?��:?؀ɼ�/\>�jO=���u�,�l��&~F��I$��F��b��'���=��������5*�T�?ߟ����]=*_?�</�ΒX>�?V=�`ټ��>3�>�t>P�K>s��>��={�=B��=6�>e��>�3�&���#@���u��B�<�w��>��0?J,�y(὏���V�������>��?&��>U�z�J(s��ʇ���>��׽�۸�v����q��kxs>�֜>-(��<>k��$�>�¼5�=��>f��/�<Ll����  ���>�ɾ�'�=�LP>��?�Tz?�4?)�=)O�>��=>�>N5�=�\]> �>���>?��1?��?���>�y�=��^��߆=K|�={��z�p���W��x��=����o<n=�?�=�x�;�'y=���<��4��dy�2�Y=z;�>�[?_��>��7>����y��I�a�r;-�a=���=;rp>��#>R�?^�5?C?k�L>1M;�����p���>ӝ�>�9���P��ּ͇^z>E�>&��?��Z?-1$>�����	>Z��U?,��>��O?��>-{=т�=����3߿���(�$�q���ѽ���<�;��b齼�v�0�y���5��ɽ�@>?q>Wuz>l�4>3��=�M0>��>#�>й2=t��=�]���.��A���3��"��Y;%>D��=���=f^=����C������b�~�� ��A�>��?�X=H�W=��ĽZ �,虾���> �>�?�`?y�@�yz�Ӧs��qJ�e����>W�v? g�>���q��>_0�(���$� ?���=�3>�k�=����������4�W>�j?���>� V�0{���~��(?�B`E>�A�< nY��\�?g�4?����� ��2`���B��)G��P½��=$2��J���7F���1���1�A/3�6���_�>=|�>R�?W2о���:)��f������!a>�W>�*�>�P)��J��M5�o�P��-��پ�X=�?�[N�6I<���>�?<0?u�>?ĊD?�]x�r�?�ܾ�9r>f��>�z�>�=?*?��>#7G>��}=Zlk��6��²�9ZX��<�Q�=�t>��>}�>�Z�Qm�=�8>6��=�@=,��<���󐽩)м��h�ڽ�=G��>x�8?�"��c�оp:�<<O>��<䛐>��"?Ƥ�>&&�A(>"��>��?P+?z(?�M>Y��vv�����<}�=�1�>lI?�?�߅�)�\��D侻���d��l
�=�f���)Ͻ���JX���P%�M��=���>I�[>1NO>[0�?��Y?��+?�'[��6�����U�a>�>�X�<�U?���>���>׆d���E�)���]牿"�ƾx�?5A`�`g��u�	>5Fi>Z<=�Xh=9��=��=���|��l9����<�ܶ>@��>��?���>j9�=�}Ӿ��9��4f?�	����3
=�e��Y>}�>��#�.�:��a'?�8>�,B��ƻ�s̊�wC輥��?��?�ʢ?Ţ�<�)��XN�>�[�>�%�=�Q��Jd���Js���:=�45>��>�A\��K����>��>g��>�-R�_�0�����kI��"�Ϳ��K���#�X���}C��Ҙ ���Ⱦ">
��D>�r��\l9�"��WȖ����=���^M��w��8��4��?���?�t%��/:�βk�ja�*�[��>'_¾*A>4�������h������E �6,�"���Ŀ���9|�>c��������J�&����kܽ�2D?,[����A��{b�=��1>	.�5�m���jɞ��Ƚ�Dd?�B.?��ھ$A�e�_q�=�0�>�"�>)�U<ȿ��Y6���>o�?�=3�a��y��Ŗ��M;��?4��?`�??��Y�a�A����R%��E?� ?��>��y��c;���: ?��:?~��>ˌ���ρ���1��>;O?��N�G�c>��>�>_�ʽ�L���P�'�޼ҰD>�hE�r	���M���G�c��=��>�h>V�^��J��R�?D����G���m��<�>�Ś><%�>�$�2�	#??( ?�d-���y�W����rѾ�j?�F�?��?�o'?�.�����"�}��[�+?���>i)U��/V�G�=�f�>hO�$�V�����ۆ>�{�?q��?�|Q?[�h��VӿZz���۸�4V��*	>�q�=�f*>���Pd=yo<||���ټ�>,��>>8�l>��>��B>$wA>8'���y$�%٨��P����:�ts�7$��E���
��l�����%ǾR�־V2d����:'Qq�tP��ؽڛ�;�ž�ݩ=	��>�/?�[3?'�=���>
赽Q��������z&۾4V&�z�S�*������@d��<\@ؼ�r����j�?�X�<[W�=�?@�A���3>�L�>�|>��+=�{>�| >��>!��>�h>��G>�u#>��+�>�h>	�}�e}��<�����;.�=jG7?gJʾ��.�4��A��������>�3�>͟���О��Ă�N�����>#(�FA6���K�<^[��K�>"Ѵ>��,��=6?��5F��IB��}p=�E>������>	?ڽO\O�K;(=��>0l�D�p>���>�!%?9bo?�D4?�,��&�>�$�=��P>�f=Z�X;��>:	�>�-)?��7?(�?Us�>��&=���"��ܤ<��\��Q84����_S�������鼜��'$+=�1!��>%��8��������@?�>�SP?غ�>��|>��WOC�]�]��q�;_�>l~ͻ�1>���=��?qd?��?�i�>w���(���2?c	 >E���{����:�'[�>�u�>�~?�p�?�Ũ=Zm����+>b�>C��>�O?l��?z��>��>�����pؿm�2��4;�z1��:ž�!��vV>���Q���y#�rr���^m>�+�>S��>�U�=a�v>�HE>5�	?6��>c��v4ֽv��G<��:���=A�ݹ@��=u�=���=҇,>�sau��C�;�'~=Ю���d�qS?"?�W=2�j:�(����:���YAE>q�>}�>FC+?6d���(�x}�ij��ľB�x>�{?��)?{9о�Tl>�ZA<�$=��?.�=[�K=��^�;,~=,|羸5�����>ۻ�>a3�=R��=ƌ%�� f���(��5n>?4�=rP��u��?��\?ʪ�����P�������î>������K�=��OpF�Y�*���(��*�������>�m�>��?�����@��Tپ�%���]��[����=�Q	<���>����C���5�e��L7��W��5�>1�D?�|K����7f?�Va?}�w?�!?��@?	k��_ڼ>A�ʾ�Ү=Ӵ�>���>-�?�F?�%?T{�>�`n>�G�<�l���a�<���w}��0">K.M>s�=o#�=wz�=D�;�.¼���<%��<+J�]��i�۩=m�=hG?��(?�a��B[���躻S>!5�=�Y�>��?.X>�$־�9����>��?Z?=�'?V��>�%˾����� �X&">�*?x{A?�G(?|ꐾ�2�ԉ�������<��>�=���ֽ¦���E��Y��*A<,�> �Y>��>��|?=M,?��?�̢=�-E����Npo�v�>��=�=�>,��>2��>�R����;�jv���p����*��>lv�����T�=�>B>fl>ک�����<�y~=ƥ��eq�=�u@�<)�>���>��?8�>��>ř ���@��T?����9���w�	�۾��<�>k��<�5��;�$?W� >�Ov�����!E�|c�=E:�?s��?��?�҃��0���x�>G �>s�9>�
>	�����*��g;=�y�=�B">��o�p��(E<\|y�]��>�ㇽ�R$������������F�+�I���������yY�ǧ�1zd=r�A��r4>�$����O���9���[��-M���4���c���Ϫ��Z�?!��?���c
��i55��8� ����4�=?/��޼6>8) ��2"��u��*�j�f�B�ؾ��,����Ԋ�>�`ߺ����wx.�U9�$�z=(�5?-�޾h�ĽYŴ��A�>�m�>&y��3l��^���B����ʼ4�k?��D?I����Ƹ��؝=n��>J ?���=�炾gg�d��>L
S?>>�ҭ<Π�.׎���=K�?���?��L?����O=����`�Z�t�-?��!?�_�>����y�Y�=��	?�?t��>�r#�*�x����?NR?z\�8j�>,��>�pr>��ǽ�۾��׼AҖ�¢<���>z&m<d(��,"���3�=�<ɟ>�>�1@��j����?/�ʾ��tt˾�Yؾ󄎺ȡ�=΃K>������>=/?e��=w}Y��]���¤�B�U�d��?���?&�q?=2?�!�Wr龴+��->e?S��>,���am���E>൬>�	���0f�Ԍ���>���?���?h?A7D��ܿ�J���l���w��f��=�'w���F>`��=��p=�����v����V=K�=r�^>��2>��E>�� >�>�g>⏅��������������W�'���]禽�)��S޾��6��(������Iw��gJ�۪'�񆁾�a�t�ʽ������A>~"?��>��?u�>�[�=�b����3�G*Ծ�VL�hc��@�z>�8����<����:�l���!� �Խbz0�%�S?�n�=׮;%�?��!�Mz�=��<������>w�>	��ʊ>�b�>�;n;��ѽ6>�G=Ex�>]���X����X�0%���=���>�M?;��<>��>������|�>-y?	�(?䝣=�:��(p��q�+��>����E�՗n���	�G�>���>#5����>c���N�ͽ"��=M�B>A�>�m">�� >�c۽-L�~n���>�#ƾ���<G�=y=?/G~?c�:?;(�=�f�>�V>��>#�>яv>ꚜ>�Ǣ>~?��'?%�?6��>��=qY?�6��=0>^� �Jr����4��x?�wcu���[;���,�1=�T�=@�W����=^�=�N��E0<���=���>�]?S�>T�T>�|�\�D�NX�Q;}Q�>�u]�_8�>3��>Tj�>6��>n��>^XW>*D ����5^;F ?��>��x�<܌�D���?_��>�H�?��g?[OY=k��FǇ=�a�=��>�*?.,L?]:�>T	�>���=d�4�˿c��/��o��c����[;��t���n��p����G�u���D=��X>��y>��C>	��=Ll�= z>�n�>v�">7҂=�J�=�_=<��伺н�k��~�G�l>�ɍ=ti2=G��<~]	���V���4<�/Q��$�<����?U�(?��<@xؽ1h���㾸�,�<φ=��5?��$?��?�e�^��	P��#j��m���M�>�_�?S9?�W�x��>����<ƼB>��>�Ys>�'+��l�=��e��t��W?�J?� �>�OŽ˚r��ꐿ��4��*�>�>�;�C�f��?ľ-?FJ��WL.�
M��:Y�>?D�n�i<���y;��G׾��<��8���#�p��;�[<�cI>���>k��?4�۾B�=�qx��*�� ����u��AI>�� =x�>�Ԣ�	'����f�ey���ƾ({�=�8>��?dyB�EZ꽨oG?Q[f?�UV?�?��K?Xnq����>0��:�<��?�[�>��-?��G?��>^S�=�=$6>���1��T�=�3>�:=,��<ɿ�=TI'=}���C�<�����C��
q��(��=CJ=��R<$%�=u�>���>�'?b&��@����<�>}L�=(�>�W�>}�3>̀����-<?w?p�?�^�>�?�<��þ�(�?��N	�>�c�> ?��*?����z���+�|���(<n#t>���D�����X"�Hʾ���=B�>��n>�k�=>6�?��?�?��'>�G{�H������j��^����+?��>�>��3�e}+��y�6s���[Q���!>����=��> f	>ף|>Đ潠a2<j����`��Tٽ�̴=�a�i�}>��?l�?�T�>��^>I����t�-;g?�����羵g���s����=O�=_'��ࢾBm�>�+�<��[�]��������h���b�?|)�?Ki�?�D�=�"��4�>]��>�p�=	��=O��E���m��=��>���>�9��5�����=iy=;Қ>����!�����M���ݿC0E��,P��8��.�Ǿ��� ;;��>���_L�r���8þ%\����7�x�-We�Z����������?|l?퍑��(��I��Q��v�>:�����=SZ��L�s�y�������P�Ͼ*[�i��!����>경f��QDL�>��x<9����<��6?�̾�k����m��=^Z�=Oiѽܸ�񄕿���U�����d?swA?ڞ�(;��b����=�#?�Q?�x	>��fIɼy:�>!%?���>4���ɓ�����=f�?A��?��??7�i�ۗC�M��j�B���?
�?il�>�Wf�y�������?<":?V�>ȩ�Y�{��h���>ڣD?��I��>f>f�>ҁ�>�u���v���T��G�}+>-��;Xj��i��IE�C�=>�f>~�J�����i�>��]��)�����B���j+���;nm�>��Ӿ�ޒ����>�[���:�����vN|�(��J�?�z�?r�?�&?���U6����9>�	ȾB�<� �>ࢁ�V��ɹ?&A?s�/�p�g.R�WR�>	�?- @F?�n��hH�Eǧ�d���������=�W�<�op>�=��+_	��Y½����a;�"���Z�>�}>��>�/�>	=�=4�=�߈��#�Z;��_ݐ�P�.��������b����eI�ӛ��}�#�6��{��L�ؽx5�S'0��~.���X�u�f�Od\��W�=GSL?67@?��I?XϹ<��.>�{�=ޏܾ=G���M=�~6��(�X�/�焗���l>��.>��w������'�N�?���ݰ]>	�?>/ｪڕ>�s>�j
<��.>���>�s�>WZ�=�,�>w8�>K�>moX>%�>վ�>e:>��j�o�n�=�0��I��R�t>5?�0���Yƾ�5���	�"�����>L)�>�%�>;�jF���i�SP�>�Q�=�s���;3�1_����e>���>��.>CǦ=!ꦽ�0�T0Ƚ4^>R<z>��>-��=>�Խ9=��ʀ�����>�����}>C��>�A??��e?+>?܃�>��->�s�=�ř>���=�G>��D=4�>�>?�,6?�"?�<�>F3>�ߴ�[1�=�y�=I�E���:;ս"�Z��k�=>y��r�<�>/������=��h��]Ľ�	�]��<a�>tG?d�?�? ��>q ���8����ؐ�>,93=n��>E/?�Vy>��?�<?�Ÿ>	�=ns��]�(��>J�q>�z�?\��'�A�;>�0�=G�-?�y?��t�Lz=y"<�5�=h� ?��>��>ь ?��i>k-��b���� �C��ٝr��g���( :iR5��OǾ/1��eW<����$����o=�8>��J>�>�ϔ>rR
>'�>�'>z��=w��������I� ��>w�}>��=�/W=jq,>L	,>��Y��0��A$�Uս2��]@D���>�S�>˞(�kq�{���/�����D�ur�>R�?��'?�;?��<P��Yt�8eE�����=��?�T�>.���)�$�� ��E>p`$>���>�<�>_��=�_�������`�Q{I>��?៞>��L��&%�"�1��l��ɛ>q��=��S�P�?��?a�Y�2�ھ���Z���<��Ża?���S���׾��s�,�߾�Ѿ�۾�4)X�쿕<kޤ>�.�?h'����	�������e�G�����>��<��V>	�>?�x��ȧ�9�>� =?�c��K/�Y��>t�=:N�>��,?�>?P�v?�y�>(�>2?��[	?�qU>,Q�>u�>Z�>#�?l#?�x�>���>:J6��2��%����8�(B�;uj���=��:>�O'>�(<x"@=�0<=���;���<T<p�i>}>���=�0�=D[�=���=���>#��?�W�=ˉƾ�kt��=?5�!����>��k��lȾ/�=�M�>�b�>��t?�^K?�uc>|n�ef(�m����И=H0�>�Ǥ>��>md�}|a�.��"k��¨=��=],>$�X�)�Ǿo{U���N�m��=+�>�T>��k>��f?�`?�{S?v�>ǚr�~E���@8���i>�>s�T>���>�u�=x�3�����p=�z}.��o,�ƣ!� &,���$<_ |=�.�>���>4ʺ=5�=l杽�t���B=�T�=;n�W��>^�?6�	?�/�>j�>e8��[���7?�5����@��=\>���8�޾?�>=�>0��36?q&B>K�̲��RYl�0w/>�ɵ?��?kj?3��2���b,=�k?=g�>Ѽ�>��
���=E >��>k=���E��Ѕ9���B>"��>,#�=ϔ%��?+�PG�<�iÿ�	G��j"�
�꾛bȾ���n.���8n����:6������M�4����A�����,3���|��,��\˾I�?ȟ?
�O��GB��aD���!�#���|>����Z��	��+�2�-��fT��û�w��K~�	S�##���;>�:H�2򢿡�w�=�~��m=���>�=�>��~��IϾ𒆿���=���>�=�cK�*$��xę��ɩ���]?�bK?~���/�?�/=O>!k>��X?���>99�n�S���	>�8�>M�X?��E?��K��z��az�)�D�K��?"^�?�%?����&�Y�_ݾ����5j?C$>��>�-�,I�<���<G�?�`?'w?�$��s�5�H�G��>zZ�?ʥ���u:>�F�>�⌽��{<�f�ѽ���;$Y�<�L> �5>U�Y��Ѿ�4��6>���>@�p>��Z��U;�=?P�i��N.���8�B��ga��t��<{?�ξQd7>��>c�p>�8�&#_�f񋿅��;.�]?X:�?�?�a&?�+��b�����k�6����>(-�>�0��[�����?~i?a&?�?�f�:mS�V ?R�?l
	@��|?2ܜ�ݿ�b��s�������y��=|�=� �=���Tp�=���<_4[=,A�=!#H>̛�>�t�>;�>��B>��
>#��=�ى���)��:������\_I��#�3��:�,�������W����L����̾�νEuȽ��7�T�G�5
B�Š㽱����;�=4�?0��>��?ѳ=�+�<�R=�Oؾ�dҾzϐ��}۾ͺ5���gF��)7�ѫ�2����3M�2Q���?(\�;ߴ>�?�C9�ay>ᗊ=�'>�4<\�~=�X>ii�>?ߦ=���=*�ȼ���=��V>������=����Ö�b1;��ZX�HQ>sW?{���پ��X�:�v�ľPv>���>��=�H+�rڱ���a�s�?Y�¼��۾�	���!�Ӕ�>��?��=��{>�Mz<ɭZ=��>���=��H�� ����D�u
U��b�>�3�>6���,$>���>��1?Z�?%�<?Tv4>���>��%>��>���=;V�>�9�>�ڿ>F&?s-?��?���>�>�~U�j�����R[�*xٽ�I1�x��<ы+;���� =|j=>��=_�u=��	>6;12׼��{=k��=�?�m?���>�q ?���<��S��,~�u�Xn�>��P�ޘ�>�z?V?_�,?oX�>�#>Q��c^���%�V�>�t�>��s��֚����A��>>"e>��\?�4z?����_�����?��=s�>�S�>�?�P�>�_C>Ge_=��mӿ�$�G�!�;8P��;s�<���M�x9�7C�-�@���E��<,�\>!�>7�p>�E>��>�<3>�R�>�HG>,ф=J�=<�;7�;|�E�֘M=N�EG<��P�����1#Ƽ�������U�I���>�:�\7ټ�} ?x ?#��=�r=;��J�����B��>?a�><��>��?]��8G���o����W�G\�>v,W?�L�> ���?>'-�</��=�}*?��>P̙<��<ع#=�S8��f�=/!�>/`�>��>9���m�{�.����R�,��=WA�=Ƭ�,��?_�b?�K��A魾�J�O���bU8������S=�"��C�v�VF��N� ��������:�%]%=���>^��?��ľ9Cp>��*�ݗ��!����@�C�=S,7�⢲>��o>#�I=�"��a��l����4��=ػ�>�B�<In�>0S?�j5?��?*?Y?��?<��>�<�?��[�K�>0?<?"F?�5S?��>�w�>����-�A��A�>}��L�t=( �=z �=Z�=Յ%>�!ʺ�?�r�<W��e�O�(��s7��X�=C�=�D<�w�=�	>;�?��5?t�"�n�.:���;���f<ۯ�=��>)�4��QB�������i>�d?��.?�`�>!�~=ݧ׾�[�{����/�=Sx
?1�?�R
?��=�51>/ھq���+>��0>�޵���u�U��8��p��c��>���>^m�=H6>W?�+?��?����Fc�<���?��v��CU��R�>��>4��=��־ּ��HO�?�B��*(�C�8=$�q�l=���>>XT�>hxQ>��;>��&�&5�=ݘT=/{>�'�;1>$�!?��?��>�	�=�B˾^O�S��?�����羥�#�'#
��[��?�>���>M4ݾ�֍?%w�9���&�Ͽf����>E�?6A�?�i�?����a�r���P>˭�>G��>�i>���.����s=�z�=H��=���z��������.=Wc�>�a^�����7-���<�}��q�\�7����p&��"ݾV��|��������	����G����O���?��:D�x$��m��U����?�b�?c8ݽ���#S/��tؾ$nؾ�C���l�H�|���J��D��,���������+�,�9��l��������@΍�"���]�hܫ�n>�l%<�N���û��&�$E�����=�����+\�MZ������}��ڀ?�O	?���� @�8�c=���=��>�4M>�">�en���+�-�+>�K?X�3?���=����K]����餥?9x�?��?؋Z���[��c��U���?x�?2��;�� ��d��/���RB�>��.?h9�>�M�F���]7���?Ӓ?�8��܀S>{�>��n>�wW=����� ���5�
�=a�����<x�}=�����\н��;(*�> �F>���a��� 7�>&���7S\�k�^�����3>>c���d�>�wl� �<m�=�	�>����x�=Á��RԽ21F?c��?�	S?�|?US��5���?�3=;��=���=��>e .>K� �ċ�>.��>h��2i������>���?���?�]@?\h��G�ܿ-���爮�'Kþ��S=�`�=�P�>�?��^O�!;����˽��~<�ȇ=���>/�>�R>X�=+>�Fp=�-��<��	����s����D����Yf��ɝ��z�旁�'�#�s�;S�ɾ#G���i��w��r�1hE�'�ѽ^���B9�>��V?���> �<?�wY�u8�>Q�J��?�,]�=���>��?����>���ͼ?�=�V�
�iq�z���E:���W?$L
��ğ>T^?��E����>�+> ��:��_>�H>���>cQ>�P�`���o��=���=��=`gn>�8�=�脿i1��-?���L�q�;�=?)�L������5��Iܾ����C �>Q�?��I>�0'��v���v���>?.�"[{���)+��>�>���>�P�=�,'��]��sv�Bgս墧=���>ԍ�=uK�ޑ�������=��>�e����x;�?>�U�>;a?ڋR?��<|�>��#>P'�>��=>SqO>-O�=F�E>׾?6j>?7?K�>L+�=�.o��`�QP>����i�o<��,��}=v��=*�ƽWz�=Ĥ޼SnS�#��=竌>��>b�<��;N�>^�g?P?$�?�=ՓN� f������~)�>��v=�7�>hF/?�x(?�'?�?�Ȭ=�^�w�����Z�>N>��>��s��ݬ�è�>���>@�B?�  ?�����Y%�HF�<\�T��>�
?^�4?Ep�>��>-�0����hyۿw 0�:����;u��<��+>,(������q=����U����E>O�7>\�=��>�ߖ��:�<��=���>��=�TQ�,�>=��="=����I>Z>�^�<�=Q^<�H�	s=e���I�����=S[=���dÿ=�\�>���>�̽�������q�ҾRX�]bd?�D:��Fg?7�f?�վ�ࡾԳ>���T�,���?�|?���=����=�����G��Ϙ�>�,�> *�>�̥�w��nh��Ɲ�>��>�D"?�w?���~R�M�j��6��Ѽ�>8_=���2��?�.h?�$!��)�$���zQ����:�bϼ���6	�}S*�����j�Ⱦ��۾6���҆<���>���?r��*�D>e�ྼ䢿�'������=�7��N>�\W>��=����"�_����8��>Cz�>{>�=��>��*?��?l?���>�R�>�����?��d=��>m�>)�?7?8?�\�>T>U[d����&r���'�\=� S�=FvA>�~u> ��=u�ʹ�h�ꜽV�%���u�Z�a���=k��=�I>��p>ʂ?�b3? ���<Z =�Z�}�f$>��<�w>7.�����S����>'�>Ω&?��>x��=�O��_P���c����=�'?�&?���>�kv�g�7>ܠ�	��
�'>?�a>
r/�����|�����������>��k>=xK<"�=N˄?�c�?gW�?,r>�Y����}�z/׾"���B�=2=�� ?���>Aɿ��Е���f�:g�M�h�,:F��ZN�z�g=�*��L?'>\�>���=�d���~��l>٥�=b)�e��>[�>��"?���>N�#>������A2�[�K?��������|�&��=Z=��>�v���>p��>q�#=?�X�m����:�39Z?�3�?~��?��?p1쾰����4>���>W#>��= G��FT&��m��)X��t�1> m1�{���B�����=��>R���l���������\�Ȼ��j�L�9~d�W�L��2ʵ�����q��>&];�Tҽ����&�V���ꮽ:��	;
��t�%�o��I��?�V�?�A�lӾ�J��8d���Z���`�T*���/�3�Ѿ���͊z����p�����s�!��kf��c����=�N��B�������F��;>����	<Pn�=_(��J]�7c�>::�=��=�7������Α�䣒� ��?(K?���;�!���=|��>�;?��*>V0>C�����A��u>�H?3~?�%���d��\i���ʽP�?�O�?5MG?n¿���1�������w=�nM?f��>\�>��ܾKi;�t@�=��>��'?R�=?��&��g��"��z$?��?�����%>�̃>~F�>������ȼg�R=�X��rD>�w���G�<��#��0����؜9>#�L>���>rcڽ޾��=?P�i��N.���8�B��ga��t��<{?�ξQd7>��>c�p>�8�&#_�f񋿅��;.�]?X:�?�?�a&?�+��b�����k�6����>(-�>�0��[�����?~i?a&?�?�f�:mS�V ?R�?l
	@��|?2ܜ�ݿ�b��s�������y��=|�=� �=���Tp�=���<_4[=,A�=!#H>̛�>�t�>;�>��B>��
>#��=�ى���)��:������\_I��#�3��:�,�������W����L����̾�νEuȽ��7�T�G�5
B�Š㽱����;�=4�?0��>��?ѳ=�+�<�R=�Oؾ�dҾzϐ��}۾ͺ5���gF��)7�ѫ�2����3M�2Q���?(\�;ߴ>�?�C9�ay>ᗊ=�'>�4<\�~=�X>ii�>?ߦ=���=*�ȼ���=��V>������=����Ö�b1;��ZX�HQ>sW?{���پ��X�:�v�ľPv>���>��=�H+�rڱ���a�s�?Y�¼��۾�	���!�Ӕ�>��?��=��{>�Mz<ɭZ=��>���=��H�� ����D�u
U��b�>�3�>6���,$>���>��1?Z�?%�<?Tv4>���>��%>��>���=;V�>�9�>�ڿ>F&?s-?��?���>�>�~U�j�����R[�*xٽ�I1�x��<ы+;���� =|j=>��=_�u=��	>6;12׼��{=k��=�?�m?���>�q ?���<��S��,~�u�Xn�>��P�ޘ�>�z?V?_�,?oX�>�#>Q��c^���%�V�>�t�>��s��֚����A��>>"e>��\?�4z?����_�����?��=s�>�S�>�?�P�>�_C>Ge_=��mӿ�$�G�!�;8P��;s�<���M�x9�7C�-�@���E��<,�\>!�>7�p>�E>��>�<3>�R�>�HG>,ф=J�=<�;7�;|�E�֘M=N�EG<��P�����1#Ƽ�������U�I���>�:�\7ټ�} ?x ?#��=�r=;��J�����B��>?a�><��>��?]��8G���o����W�G\�>v,W?�L�> ���?>'-�</��=�}*?��>P̙<��<ع#=�S8��f�=/!�>/`�>��>9���m�{�.����R�,��=WA�=Ƭ�,��?_�b?�K��A魾�J�O���bU8������S=�"��C�v�VF��N� ��������:�%]%=���>^��?��ľ9Cp>��*�ݗ��!����@�C�=S,7�⢲>��o>#�I=�"��a��l����4��=ػ�>�B�<In�>0S?�j5?��?*?Y?��?<��>�<�?��[�K�>0?<?"F?�5S?��>�w�>����-�A��A�>}��L�t=( �=z �=Z�=Յ%>�!ʺ�?�r�<W��e�O�(��s7��X�=C�=�D<�w�=�	>;�?��5?t�"�n�.:���;���f<ۯ�=��>)�4��QB�������i>�d?��.?�`�>!�~=ݧ׾�[�{����/�=Sx
?1�?�R
?��=�51>/ھq���+>��0>�޵���u�U��8��p��c��>���>^m�=H6>W?�+?��?����Fc�<���?��v��CU��R�>��>4��=��־ּ��HO�?�B��*(�C�8=$�q�l=���>>XT�>hxQ>��;>��&�&5�=ݘT=/{>�'�;1>$�!?��?��>�	�=�B˾^O�S��?�����羥�#�'#
��[��?�>���>M4ݾ�֍?%w�9���&�Ͽf����>E�?6A�?�i�?����a�r���P>˭�>G��>�i>���.����s=�z�=H��=���z��������.=Wc�>�a^�����7-���<�}��q�\�7����p&��"ݾV��|��������	����G����O���?��:D�x$��m��U����?�b�?c8ݽ���#S/��tؾ$nؾ�C���l�H�|���J��D��,���������+�,�9��l��������@΍�"���]�hܫ�n>�l%<�N���û��&�$E�����=�����+\�MZ������}��ڀ?�O	?���� @�8�c=���=��>�4M>�">�en���+�-�+>�K?X�3?���=����K]����餥?9x�?��?؋Z���[��c��U���?x�?2��;�� ��d��/���RB�>��.?h9�>�M�F���]7���?Ӓ?�8��܀S>{�>��n>�wW=����� ���5�
�=a�����<x�}=�����\н��;(*�> �F>���a��� 7�>&���7S\�k�^�����3>>c���d�>�wl� �<m�=�	�>����x�=Á��RԽ21F?c��?�	S?�|?US��5���?�3=;��=���=��>e .>K� �ċ�>.��>h��2i������>���?���?�]@?\h��G�ܿ-���爮�'Kþ��S=�`�=�P�>�?��^O�!;����˽��~<�ȇ=���>/�>�R>X�=+>�Fp=�-��<��	����s����D����Yf��ɝ��z�旁�'�#�s�;S�ɾ#G���i��w��r�1hE�'�ѽ^���B9�>��V?���> �<?�wY�u8�>Q�J��?�,]�=���>��?����>���ͼ?�=�V�
�iq�z���E:���W?$L
��ğ>T^?��E����>�+> ��:��_>�H>���>cQ>�P�`���o��=���=��=`gn>�8�=�脿i1��-?���L�q�;�=?)�L������5��Iܾ����C �>Q�?��I>�0'��v���v���>?.�"[{���)+��>�>���>�P�=�,'��]��sv�Bgս墧=���>ԍ�=uK�ޑ�������=��>�e����x;�?>�U�>;a?ڋR?��<|�>��#>P'�>��=>SqO>-O�=F�E>׾?6j>?7?K�>L+�=�.o��`�QP>����i�o<��,��}=v��=*�ƽWz�=Ĥ޼SnS�#��=竌>��>b�<��;N�>^�g?P?$�?�=ՓN� f������~)�>��v=�7�>hF/?�x(?�'?�?�Ȭ=�^�w�����Z�>N>��>��s��ݬ�è�>���>@�B?�  ?�����Y%�HF�<\�T��>�
?^�4?Ep�>��>-�0����hyۿw 0�:����;u��<��+>,(������q=����U����E>O�7>\�=��>�ߖ��:�<��=���>��=�TQ�,�>=��="=����I>Z>�^�<�=Q^<�H�	s=e���I�����=S[=���dÿ=�\�>���>�̽�������q�ҾRX�]bd?�D:��Fg?7�f?�վ�ࡾԳ>���T�,���?�|?���=����=�����G��Ϙ�>�,�> *�>�̥�w��nh��Ɲ�>��>�D"?�w?���~R�M�j��6��Ѽ�>8_=���2��?�.h?�$!��)�$���zQ����:�bϼ���6	�}S*�����j�Ⱦ��۾6���҆<���>���?r��*�D>e�ྼ䢿�'������=�7��N>�\W>��=����"�_����8��>Cz�>{>�=��>��*?��?l?���>�R�>�����?��d=��>m�>)�?7?8?�\�>T>U[d����&r���'�\=� S�=FvA>�~u> ��=u�ʹ�h�ꜽV�%���u�Z�a���=k��=�I>��p>ʂ?�b3? ���<Z =�Z�}�f$>��<�w>7.�����S����>'�>Ω&?��>x��=�O��_P���c����=�'?�&?���>�kv�g�7>ܠ�	��
�'>?�a>
r/�����|�����������>��k>=xK<"�=N˄?�c�?gW�?,r>�Y����}�z/׾"���B�=2=�� ?���>Aɿ��Е���f�:g�M�h�,:F��ZN�z�g=�*��L?'>\�>���=�d���~��l>٥�=b)�e��>[�>��"?���>N�#>������A2�[�K?��������|�&��=Z=��>�v���>p��>q�#=?�X�m����:�39Z?�3�?~��?��?p1쾰����4>���>W#>��= G��FT&��m��)X��t�1> m1�{���B�����=��>R���l���������\�Ȼ��j�L�9~d�W�L��2ʵ�����q��>&];�Tҽ����&�V���ꮽ:��	;
��t�%�o��I��?�V�?�A�lӾ�J��8d���Z���`�T*���/�3�Ѿ���͊z����p�����s�!��kf��c����=�N��B�������F��;>����	<Pn�=_(��J]�7c�>::�=��=�7������Α�䣒� ��?(K?���;�!���=|��>�;?��*>V0>C�����A��u>�H?3~?�%���d��\i���ʽP�?�O�?5MG?n¿���1�������w=�nM?f��>\�>��ܾKi;�t@�=��>��'?R�=?��&��g��"��z$?��?�����%>�̃>~F�>������ȼg�R=�X��rD>�w���G�<��#��0����؜9>#�L>���>rcڽ޾��
�>]��)g��[d�uk��H���&�#[:?��񾃛�>]��>�>��0��j{�S����м��J?�2�?|�(?xCC?�<o��d*��"�>{��>�+?�I�>�#����y<���=p��>'�8���ξR/�G�?�$�?8��?E�D?�タ���x���c�վ򲉾|�I>�>��J>��� �>�2=�=+������=�^K>:�F>U�^>z.>>�D>>��>]���2 ����~7���6�c���
���P��ؾ�E8��x�Nä�o���`Շ����R#Ͻ�0-�.���d���7�����>�'2?<2?0y�>Ni9���E>zJϾ�^6�I�޾_�!����z��7��h��M����ɾ:�ᾌn�g.��+罾�Y�>8�]���k��"7>�>|w�>k�8>��=���>D�W>n��=��>==۠�<B�B=Y�|=D�=��>�+�<=d�Kmq�^5�Q,#�	��=�d3?Ȕ?��	��$�������T��>��!?�b>b*��h����l��x�>3��=���-�(����9>�4�>b�c>�=�=;|�gG���$����>�(�>>K���œ�<F/�844>���>b� �q
�<,�h>C�,?Ms?9g#?{v���֛>D6~>C�>B7�<���=ܺ>�[�>�$?�=3?��?eZ�>�=�=��3�}r=�3=٨]������� ^W�-�q�z������><n� =:��<��=�:�=�ck�Q�<y��=�>p�Z?�8?Є�>d殾l�6�-C�D2����>h���$=Q0�=,��>���>��?&7�>!<>a�������?�'J>m}�܎��,�[��<�=�h�>��?��?�}t=q`�N��=��V=�>Z�?#D>?���>�)(>Ďv���
�YaϿ�Y��D�:ᓽ �4��ˀ;:�O�b� X����%��@�.��<��U>�[�>�5d>�wC>��>S;>���>��3>ƭ�<ưA=Y�E�)��;i�&�N�s=+pj���0=w�|�v�`�y䪼��������~�)/c��"=�ю��oG�>��<?�`G>�"���ǲ!��s!���?ˮ#?˦H>�V�>�1�����||��D*�i�ϽR�L?��n?��>������ �>�ۥ>�	A>_� >�b$=�.���S(�a�)=Y����>�k?� s>�[q�W������������>kn�����;�G�?��Y?PQ��]��U��j/����j"��zH����ug��9��������2m�fȔ��ş=3�>�h�?Wmn������yҾp���p����P�7�u>�)=��>���=.�7��=���;;����{��=�a�=@~]>������?��?��,?���>�I9>���>z�a�}82?��2�*?�!?�+�>�>z�>!
�=�K=��^���<(�����Y�=Uby��U>tY�=�Ao<�L��}�0��b]>��<�r ���%�� ��l=���;�@Ż��u=|Sy=��>��??%6�=Ŵ˽��;/E��gԅ>��=Y�>�mƾ���F��<>԰�> m?���>�
R>AG���Zľ���<�>�b{>��0?��?	��db�����ђ��~ݽ��>��g�O�˾c� ��K
��4��p�>v׉>`>?�L=	�r?��a?�O? Yw��q9��SJ�o�������;j<��>qj�>]��=ź��#�,��Z�|�K�+.����
���RR����>'P�>�j7>4�k>��:>�b�K�?���R�G%�	����?#��>F��>��>�A��������9�[?�f�XY@���ὒ�>W+�>�U�=O?�����9�?3>��`���z���@���?�3�?M��?��>��$��C�r�>;��>�>¿�<�'.<���<Y���MX->���<Y����Iž�#���ܷ>`��>P�佂���z"�qr��Eſ.'��憾�n�����DSԾv�k]���E�;5�=��;3*Ƚ�>����Ľ�8�ߋ(�cΙ�n����W��{?��l?ŕF��������,�WJ����>�ƾ�^�=:�#*U>�
��&@�*��������7�P�A���ؾ��>�I\�hB�A�n������<b=�+>?|\��N�潚����>���=�ѵ>q����_�0���*�^�,?ViG?�.�ES�Ym=�\�N�d��>ټ�>��=+�a�SI���_G>U=?�R?��\>"��U����嬼�;�?�0�?�S?炼����f�����:��D?=d�>���="X������8�=Wٸ>~��?��O?�(оQ�����E�F�:?�(�?�1��j�>t?�>W^�<͗���P��s�+<���=�~����X=	p���=#/��l]\��C�y˦>�y�>g`��TIH���=|{�q�[���k�O�5����Ii�<�?3������>���<��<>M�W�K�}�΃�d����JI?�S�?Y�H?:�?ɩ/�\�"�Y����=i!?�^�>�f���5�<�8r>��>����6O��<��j'?a�?�T�?��W?ܢ���ݿ�"��O3��
��a1�-�=�T#>��a�Q�<�TT=�O�;Є�=N&�>@�R>Ta1>��=nc�=�E�=����9��G��^����%c�����3��M�����L����򆳾{���.�&����@�����d��Jf��� �������>0p?<!?}r�>f;�<!}�=M�������L�9о̜���2��[۾�3޾�[����6V����h�����G��.�>�V4�Tj�=B�>�W!�W>Ao�=����[˺=���=�>=J>��i>Iv�>5:->Z�=���<�>γ;x�O�O�uA���73�P&�<MQ�>�0A��:xs���=�x���d��>XzZ?+�?���"k�������>��c�]\�
v�xC$��+��|�>��R<)�^>�
�=�l�����
��=m��>��a>6�����,���'�>�?��/������Q>Q�<?t�j?�L?��`�����i�=��>�,�>XSr>\�%�y�|��>�Qp?"�?�R ?td�=�'�*�v���	>g��<�����@���=w��[W�ȥ<��a=(>	>I��=����V�E����=r�=.8�>�PZ?T�>?��>]�7��U9���6���=u,�<L-ξ�!�>�> ?S��>G:�>��=U�,�����i<��?J� >�싿�r���2�����>��e>��Y?��Q?rݾ����.=.�=��>��5?G?�?�>�'��{�e���
�2Z̿)%�(-.����j}������>���)$��*��vｲ_2< �h>Vn>_�U>I�$>��=�>r��>	�>>�*�=F+�=�"�<����b���|�=*����<� ��v��;�.1�K>����K�k��s���W�����K�>G5?l��=('���p�m��A軾���>Vd>��>_A�>��=�� �L�_�BdG�{~�F�?��e?�&>w:���n=,_�>�߷>�>Q�0>1F>r�㽌�ݾ�2�*�<��?�~?�׿>ݷz��)Z�7��x��K��>���x=��?��t?c"���򪾗h���K��
��?��=�?�vbٽحo��)��-�%��<��v�_��=�i�>��?ꗢ�Ր�����ń��%Q��佗�/=���=5R?�/>����6��L^۾�j��&{H�w4���i�>Ot�;��?�A?U�?��0?��>3��>��*��
?tl�=�.�>���>�V�>�p�>Ŭ�>ϐq=G�>c{:<������E��@W�i��=�gB=��c=��=�g�=_���/(<�d�=�x�<ץ��l��d�`o��[Pu<��z=�$>�{�=!��>��,?�Ź���:�iG=DX��I��2T>5��>����q� ���[=��=P�>9^?`ܜ><G�=� پ6?Ͼ���ё�>�c�>�Ϩ>���>��]�.�ֽ�0ֽ�ء����>��Z>��|�����1��{�05�����>�~�>�|/�w�+���{?���?4w?�	���BؾI�:����L�>��\Y�>9�>���= 
Ⱦ���o{p��N���"���x�*̛�+����,�>m��>	̸<�->a�(>�X��<���Ea�q�;̯	=���>c}}>��>d>i=f���3�� ���?���׭����Pv��%��>�`>�t�=�����*?��<> �U�t�����-�Ǵ>��?6H�?�?z��M��<C�<�p>��S>��#>W>��C�I����	�=N�=+�=�vS��c>��=��h>Ƣ̽�������������_ۿ*�.��߀��`)�:�q��������#>�B��C ��Q�Ⱦ�rؽ�=���7:H�P���e�T����
御~����}?��6?�c�=C�6��޾f���L��ʡ
>}8��:��:Ž@����设2Y��{�� '��s�\����i>���� h�LL�o�����<Ud8>��?2|���%'���$��k{>�l�>���}���U�����rkk?ђ2?m����\���;Y;>h�>�B?�ޘ>��ν�5<���k=6,*?I�M?b�,�������aܘ�S��?u?�?�l]?�w��X���/����&?��V?�+�>,Ć��j��8,����	?��?7C+?�K��膿��.�Q�>rm`?p�n��D�>@�>C��=�����a����.�2l��t�;Y�b�du����>4�:��I������{�>��>>�1�o����=|{�q�[���k�O�5����Ii�<�?3������>���<��<>M�W�K�}�΃�d����JI?�S�?Y�H?:�?ɩ/�\�"�Y����=i!?�^�>�f���5�<�8r>��>����6O��<��j'?a�?�T�?��W?ܢ���ݿ�"��O3��
��a1�-�=�T#>��a�Q�<�TT=�O�;Є�=N&�>@�R>Ta1>��=nc�=�E�=����9��G��^����%c�����3��M�����L����򆳾{���.�&����@�����d��Jf��� �������>0p?<!?}r�>f;�<!}�=M�������L�9о̜���2��[۾�3޾�[����6V����h�����G��.�>�V4�Tj�=B�>�W!�W>Ao�=����[˺=���=�>=J>��i>Iv�>5:->Z�=���<�>γ;x�O�O�uA���73�P&�<MQ�>�0A��:xs���=�x���d��>XzZ?+�?���"k�������>��c�]\�
v�xC$��+��|�>��R<)�^>�
�=�l�����
��=m��>��a>6�����,���'�>�?��/������Q>Q�<?t�j?�L?��`�����i�=��>�,�>XSr>\�%�y�|��>�Qp?"�?�R ?td�=�'�*�v���	>g��<�����@���=w��[W�ȥ<��a=(>	>I��=����V�E����=r�=.8�>�PZ?T�>?��>]�7��U9���6���=u,�<L-ξ�!�>�> ?S��>G:�>��=U�,�����i<��?J� >�싿�r���2�����>��e>��Y?��Q?rݾ����.=.�=��>��5?G?�?�>�'��{�e���
�2Z̿)%�(-.����j}������>���)$��*��vｲ_2< �h>Vn>_�U>I�$>��=�>r��>	�>>�*�=F+�=�"�<����b���|�=*����<� ��v��;�.1�K>����K�k��s���W�����K�>G5?l��=('���p�m��A軾���>Vd>��>_A�>��=�� �L�_�BdG�{~�F�?��e?�&>w:���n=,_�>�߷>�>Q�0>1F>r�㽌�ݾ�2�*�<��?�~?�׿>ݷz��)Z�7��x��K��>���x=��?��t?c"���򪾗h���K��
��?��=�?�vbٽحo��)��-�%��<��v�_��=�i�>��?ꗢ�Ր�����ń��%Q��佗�/=���=5R?�/>����6��L^۾�j��&{H�w4���i�>Ot�;��?�A?U�?��0?��>3��>��*��
?tl�=�.�>���>�V�>�p�>Ŭ�>ϐq=G�>c{:<������E��@W�i��=�gB=��c=��=�g�=_���/(<�d�=�x�<ץ��l��d�`o��[Pu<��z=�$>�{�=!��>��,?�Ź���:�iG=DX��I��2T>5��>����q� ���[=��=P�>9^?`ܜ><G�=� پ6?Ͼ���ё�>�c�>�Ϩ>���>��]�.�ֽ�0ֽ�ء����>��Z>��|�����1��{�05�����>�~�>�|/�w�+���{?���?4w?�	���BؾI�:����L�>��\Y�>9�>���= 
Ⱦ���o{p��N���"���x�*̛�+����,�>m��>	̸<�->a�(>�X��<���Ea�q�;̯	=���>c}}>��>d>i=f���3�� ���?���׭����Pv��%��>�`>�t�=�����*?��<> �U�t�����-�Ǵ>��?6H�?�?z��M��<C�<�p>��S>��#>W>��C�I����	�=N�=+�=�vS��c>��=��h>Ƣ̽�������������_ۿ*�.��߀��`)�:�q��������#>�B��C ��Q�Ⱦ�rؽ�=���7:H�P���e�T����
御~����}?��6?�c�=C�6��޾f���L��ʡ
>}8��:��:Ž@����设2Y��{�� '��s�\����i>���� h�LL�o�����<Ud8>��?2|���%'���$��k{>�l�>���}���U�����rkk?ђ2?m����\���;Y;>h�>�B?�ޘ>��ν�5<���k=6,*?I�M?b�,�������aܘ�S��?u?�?�l]?�w��X���/����&?��V?�+�>,Ć��j��8,����	?��?7C+?�K��膿��.�Q�>rm`?p�n��D�>@�>C��=�����a����.�2l��t�;Y�b�du����>4�:��I������{�>��>>�1�o�澒2 �&��AsY��n����˾���F�/���+?+�����>cFo>^��>Y,A�z�喈�'iD�	�6?��?E�=?`(�?O�\�(YO���=�K<>�?)5�>u�=����3�=X6?U���n�(�"���? �?6��?a�c?j
����ҿ�z��^*��BL����=;�=N�>���Һw=�\�=���O�=�/�=JǑ>�:7>pH1>&n>�A>�7>^��%i�����r���g=���&��'�#��H��ܓ@��G�{C��xyԾ�ɽ6*9�����l��K��5=�׾���>fZ%?ۃ�>��>���=�=��#�d��� ��zQ־�������O	��WѾ�S;�s��e�@�ޥ�0˴�@�>��<&0p=�r�>��<��>Z�L>��C=O>���{�=[=f=b>��4>�,>ǣ���I	=���=-˃>T����@�O�������ٽ��p>^��>z̭�o�Q=�����T��Dվ��>=�`?2
?{[�ϩ��ؕG�r��>��J<��X��NP���U�>50>�X_��5>yg�x@�������x>=N�>h�>��'����Gwb�)��>�k�>����*͠�9=K>�o:?�?~�+?3��=}כ>���=�?�p>��C>�A���t7�H��>�:N?�1Y?[��=C�^=�Έ�E�>z�&�2'��S������A�-�1�)=���=��1����=���]�=��/>8s�="ؼ�������@�>�Ho?��?���>�X(�Q+,��M~�%�����>�؉�l;8>h�>���>��q>�S�>*�>Ð�<�#��R��Bڭ>9ן>u>B�a��� |=�>��&>��a?ךM?O$�*�g�f��=��=�0�=���>�(?/�>Z=�2������lӿ�$���!��䂽�6�L��;��<���M�@i8��-�x���P��<��\>G#�>��p>��D>ޞ>]23>�Q�>�SG>�݄=�ݥ=�<�;?�;��E���M=��'$G<w�P�����zƼ�������הI���>��7���ؼ��>��>b��:��FGj�t� ��9~<uU�>�c�>l��>���>��>"���N�mEJ�[Z��[.?|�c?��>�Q�n�=q1�Q>���>g��=!m<���"�H˽����>^�?��>�&��k`T�|�6�^������>zS���"+=?ٜ?~��?���E2����,��N}�����ɣ<k����_2�2ޤ��B�z����	�3�	�ki���(�=��>Ve�?��!�Y�>$Nƾ�ؙ��qw��Wþ���=��w>*p>���=�>�
dо}�߾�z���c���^<DZ&>�)<�O�>S20?�!?e}^?�y-?[�>?5h�{U�>�K1�,��>��>#��>��>2;�>�b0>x�	>6-��
��=6��"n�����޽o��=��1>ua>���=?�G=SR�<?`�=�o�������U�VR������=O�=cYo<���>��?Y߱=�4/�����ཅh�R1�=5@�>[�9��
t���Y���=m��>.�$?���>�d
=�	��י���.>�?�?��q>�}�$�#>ɿ��L���7��>S[>N�ĽSٿ���Ծ��޾�L�h]�>7�>}�>�(>5�{?y�c?�??t�'�p�e�a2��/н��s=�_>�.�>4B=�8�j+�(�m��5[�Z�/�a�ü��Y��l<�B>r>��>��=�s�=/
�1��������#�<<՟>13�>{��>O>aD���a��H(�vF?���G��N��YQ(�1�;=�Q>U��>Jr=��(*?���=��e�7}��/RK�"��>�?�J�?�`C?u7��b��]7�=�V>t�r>VB=��1�L��S����=s��=��w�F�����w�cï>ʋ�>/�� :��p+�����|ȿ�L-����t������ �����Q�<I����x)�qx��煦��6�����?�;�n�c�)ŝ�T����i�� g?�CM?#�J��c��3�`��J\�Ȅ>��j�������ʾ����������1��i��B�8��U#�Z)����e>�	b��`r�ͳ\����7[,����=��?ॾ�z郾|%������j�>�^>��y���� ĝ�U&���X?-?P��&����佝>V��>��>T�3>tTO�\�-�Ca>jjI?i<5?�W/=����	��_������?.��?�^?g�����*����/5���|�>��?��==|��s>;��պ�+?��?G�?4�پ@e�����P?�[o?\K7���>Yn�>bc>��Z��V�v"=��n�,wm=��U��9=���=}�#�YX�]���W?�>$�O>7�%���¾�2 �&��AsY��n����˾���F�/���+?+�����>cFo>^��>Y,A�z�喈�'iD�	�6?��?E�=?`(�?O�\�(YO���=�K<>�?)5�>u�=����3�=X6?U���n�(�"���? �?6��?a�c?j
����ҿ�z��^*��BL����=;�=N�>���Һw=�\�=���O�=�/�=JǑ>�:7>pH1>&n>�A>�7>^��%i�����r���g=���&��'�#��H��ܓ@��G�{C��xyԾ�ɽ6*9�����l��K��5=�׾���>fZ%?ۃ�>��>���=�=��#�d��� ��zQ־�������O	��WѾ�S;�s��e�@�ޥ�0˴�@�>��<&0p=�r�>��<��>Z�L>��C=O>���{�=[=f=b>��4>�,>ǣ���I	=���=-˃>T����@�O�������ٽ��p>^��>z̭�o�Q=�����T��Dվ��>=�`?2
?{[�ϩ��ؕG�r��>��J<��X��NP���U�>50>�X_��5>yg�x@�������x>=N�>h�>��'����Gwb�)��>�k�>����*͠�9=K>�o:?�?~�+?3��=}כ>���=�?�p>��C>�A���t7�H��>�:N?�1Y?[��=C�^=�Έ�E�>z�&�2'��S������A�-�1�)=���=��1����=���]�=��/>8s�="ؼ�������@�>�Ho?��?���>�X(�Q+,��M~�%�����>�؉�l;8>h�>���>��q>�S�>*�>Ð�<�#��R��Bڭ>9ן>u>B�a��� |=�>��&>��a?ךM?O$�*�g�f��=��=�0�=���>�(?/�>Z=�2������lӿ�$���!��䂽�6�L��;��<���M�@i8��-�x���P��<��\>G#�>��p>��D>ޞ>]23>�Q�>�SG>�݄=�ݥ=�<�;?�;��E���M=��'$G<w�P�����zƼ�������הI���>��7���ؼ��>��>b��:��FGj�t� ��9~<uU�>�c�>l��>���>��>"���N�mEJ�[Z��[.?|�c?��>�Q�n�=q1�Q>���>g��=!m<���"�H˽����>^�?��>�&��k`T�|�6�^������>zS���"+=?ٜ?~��?���E2����,��N}�����ɣ<k����_2�2ޤ��B�z����	�3�	�ki���(�=��>Ve�?��!�Y�>$Nƾ�ؙ��qw��Wþ���=��w>*p>���=�>�
dо}�߾�z���c���^<DZ&>�)<�O�>S20?�!?e}^?�y-?[�>?5h�{U�>�K1�,��>��>#��>��>2;�>�b0>x�	>6-��
��=6��"n�����޽o��=��1>ua>���=?�G=SR�<?`�=�o�������U�VR������=O�=cYo<���>��?Y߱=�4/�����ཅh�R1�=5@�>[�9��
t���Y���=m��>.�$?���>�d
=�	��י���.>�?�?��q>�}�$�#>ɿ��L���7��>S[>N�ĽSٿ���Ծ��޾�L�h]�>7�>}�>�(>5�{?y�c?�??t�'�p�e�a2��/н��s=�_>�.�>4B=�8�j+�(�m��5[�Z�/�a�ü��Y��l<�B>r>��>��=�s�=/
�1��������#�<<՟>13�>{��>O>aD���a��H(�vF?���G��N��YQ(�1�;=�Q>U��>Jr=��(*?���=��e�7}��/RK�"��>�?�J�?�`C?u7��b��]7�=�V>t�r>VB=��1�L��S����=s��=��w�F�����w�cï>ʋ�>/�� :��p+�����|ȿ�L-����t������ �����Q�<I����x)�qx��煦��6�����?�;�n�c�)ŝ�T����i�� g?�CM?#�J��c��3�`��J\�Ȅ>��j�������ʾ����������1��i��B�8��U#�Z)����e>�	b��`r�ͳ\����7[,����=��?ॾ�z郾|%������j�>�^>��y���� ĝ�U&���X?-?P��&����佝>V��>��>T�3>tTO�\�-�Ca>jjI?i<5?�W/=����	��_������?.��?�^?g�����*����/5���|�>��?��==|��s>;��պ�+?��?G�?4�پ@e�����P?�[o?\K7���>Yn�>bc>��Z��V�v"=��n�,wm=��U��9=���=}�#�YX�]���W?�>$�O>7�%���¾��>5����P�:�,�{�۾I5����ټ��?]������>#�>W>`> z����Y�w�Ö��=jK?��?Ф8?�] ?�hh�x����=�D�,�=h<�{|>]��<��>\��=��%��/��A+2��0 ?~%�?�6�?Gul?ق����տ^喿T��������@>�\�=u�=>����Z=A�<�_:2�I�F3 >坕>�]�>��u>��N>��.>��7>`v��!&��.��]×�*V8������������d����ƌ!��NǾ�����V���K�� �%��o*�����ո��A���D?Y�b?�K]? (?�m�=G�<���E��S�C�ξ>on�����P����*
Խ�s��N��t���yֽ�*���>�{����=��B>G㽮7u>�H>�>>�tQ>��k>�2�>��=|����	����=��>H�=���>)s�<�Kn�A�v��<�>&���M=j:(?ow=�)s�}6H����,[���ڸ>>�8?���>�(��ꏿ��d��/�>N�\=�?�,�-;�C���ÿ>���>D�`=��^>��^�׾ζ��V�>Dh�>�[>���c1˾m�z5(>�z?�K�e@��Έ���2?��p?��'?��R�� �>��>�E>!��>�^�=Ӑ���<_�>`L?�e]?1<�>:];ܽ$��=p�=o 2�w&��X�ݳ�;�g:�<J�Ȣ:�Y��<{<�<$�ѽ���={��=��=+a=������>U8?�#�>�o�>�rG�5�@��}N�?��q� >����dk�>R��>�?�/�>�]�>�K<>�F ��㻾\f辯��>��7>xL\�y�u�f�"�G�w>�ao>P?s�2?��5��i��vx<'y�=��>�??�,?}��>�%>&]�����kӿ�$�E�!�����%x���;$�<�N������-����я�< �\>J�>�p>�D>��>�73>o]�>�[G>k��=}��=,�;sM;j�E�eON=?����E<l�P��ٱ���ż ���8A����I���>�*A��`ټ'S?��>VY+�@=򽣽ݾ}D��э�?!�>=>r/?_X�>nq�>�^ �0�w���1��g��3?J�k?��> 2E���M�1�.��4�<���>H��>{Vn>��k�7ӳ�-���j�����>�%1?�*�>������c�Y�n����FQ?��ټ�=�8t��?��n?"��g쇾��,���F�ь��2�f+�x����=���5�:!��~۾.��6̖�>��=�Y�>VR�?/��I��=Kǭ��ە�����N��!�=�f�<���>?��=�0U�EI����%���;,�̽ >��>i>}�U=��>�v�>��?�w ?C?l�����?�X�>�+�>c�?pnQ?֧
?�n>T��W�3=�U�=���>����aS�A��=.���=�=E�= ��=��^���g=��=?Y���^<����	�={ۃ=dr�=��=��=��
?��)?��9>,��=,Ȑ����=Nh>���H�>���-h?��{���z!>7L�?�ŏ?�e;?�C��,��[����-�c��>���>��K?���>�$���/�y��E�#�*�5����>G��ʛ��rJ���)+��Kdl>)�>Rt��q!���?NLz?iGC?��E=)A��~��		�w|n�/���D�>�	>�>�����7�T�Z���e�j�?���[��X��@����=*��>&1>�ڼ��>J�=+G�=�U�ؑ�>�5�>Ԕ�>�Ģ>��?��R>���$�K4��"A?�㬾�[�3���g�⾔~(���>Z?s �=r�9?
C�sI$�@���J��?#c�?w��?�:Q?�޾8^����=�(�=%��'��l�7(�r>[����F.>���<Xɮ��֐�w�͛
?��#?��$>}��\�E���>�3ٿ�3�Eo��W��s&�8S2��Ę��&>֒S�/tо�ļL(��ҽ&�=��룽��B���}�!ߦ������?��p?|X�����=
nL���;���ܾm۠> �;����x
.���2=�	��	|Ǿ�9~�����6���N���aA>Kn�����OQ�T�:��偾_t>�7?�������u��*�>���>5'�=� ���&�����/k���S?�Vj?\�=�Ի+����l��>�i?t�*?��N=��Ծr� �O�<�u.?��?�H�=�������#��I�?+�?[�B?�D��U��2$�kc$>E)?R�2?�F>�-T�,�����=w�8?��Y?���>��Oψ�����<	?.�?����<*>��D>��~>�J������d��b���oY=��(>�]=>���D���K�� ��5��>��>���2������u�<���v���j��K �ز>kd����c?cϾ+�e��n�>kH�>��\��s��^�?��"��X�q?&Ǿ?�M�>���>~p��K2�@��=q%���>b"�=#�=>���g�>�$�>>�	���x����Ϧ�>Pm�?"n�?A0?3m`��u��‎�E�ξεľ�$}>�G	>��Z>����a��=Z����U=���=?11>��m>�8�=��>5>)Y>�ȇ>�P|��J1�zy׿�[��w��!�
�I���K�j�6���f��a5�Ғh�xK�������n����f��%>I�=�7#��?��/?�y+?l?�m�2�(x���4�p	�=�0��^���8�#�cs��h>�-�=#����߾0v9	da�A��>�����>�Ɨ<�d9��V7>�>ݨ=���4w7>qkL>�˥�e�J�?>{Lg>�>�g�<4�?
���a��l�yg6�p����a�>��?�a^>����9'U���#��㪾
s
?3${?ke?�2�l_��bG�k�>�l>8����-�þa���>_�>�����X>���b�)���zT�>HN�>KDX>u))�q�ӾV��ፅ>2�>������2�=-�/?��~?�.?.=Y7�>��=5�>��,>!zQ>U��= >#@�>�+?�E<?�]?;)>�>�|�<ф=+���{ݽ��G<3@�#�B���=iF���RO=���=�P>�s
� Պ�6����h�+>�e�>?�E?��?�>E릾~����e��m�<�:�>"ǽ1�?,j�>fF9?��?-��>�ɶ��iž�_�$���>�9>��c��6��Z	x���>��u>�x\?��?�`��Nh\�Wo_�u<;W��>�0+?�P6?I@�>��=	Q������
ӿL�$��="��;������=�_�-��wO�0�;V7&�����.�x<l�O>�ل>t�p>�"M>Vi*>/>�=�>��E>���=7��=�0�;F�;�J�l�H=d3��$��<�G��A����ݼ����~W�A�1>�������&�>V��>gX{��K �W��!S��\���0@�>���>r��>af�>t�;=L	����g���>��[��?�jo?���>���<� 1=J���>���>
��>X%�><d��E��\���֕�=�?^r3?���>L�8��{��O=�[]??v.���=$��?�,�?7�Ⱦ�=���H�^>\����^T>��
��� �d�\�.��L8�V�g�(�̹žm��='"?L��?��z�rZ��.7־᧿$؊�2<����u>%��=_S�>��<������"��t�>k�I�=b�;>�b#=w�>TG?��?��N?���>B�>���?��=�6�>'��>Q�?��?��>��c>K�L>-�;����d�(����˼:8�²�=���=bA>��6�9$
=�O=O�=���HM/="V<��~�.�|��=��=Z�:>��?6�?��=Ӊ�;�KҾ����%7>��<]Ԋ><"-��Qƾ7��aj>�{A?�Z?dJ�>��E�������5��ڕ>H`?=HT? ��>G�ջ��ٽ5������Ş>3�>9�>F��fH���'�t���(Z�>;�P>�x�=]�o���?�D?)X0?Q���?F�G�T�n�[��=>~� &�>=A�>}�>����m���Q� �E�n'%�x:Խ�}�1�
=$��=��>�3>��W>�>)B`�V��yQ�h'>�<�9?��>��>ʹ�<����o�o�Ѿ��n?T�Ӿq���[���"۾|^=�a�><D�>PxV���^?o�m=��Y�����a��G(	?�	�?���?��"?鳮��
>4�<a�>|��=��->x3�;�o>��R����>���>��Ѿb��_=�4?��?�5W>���E��n�<�<���J��`�� ¾�T����;K���]�۽  ����ǘ�+ub��<��q	�paǽ�2��`������H���%�?�f�?���=�T輭�/�z��L뾱�=����3ڮ�h�:����n�Ǿ󪰾�h�r#�3 %��@�G!�>"�\�>��7 }��d(�V�[���>>�=/?��ž:B���t�o�m=؏">��<��@K���ř���^�V?�n:?�뾨���W���>�	?6�>�� >�3���M�@��>4�3?�i.?�Vм�؎��$���8��"��?z��?Uk,?F��S�]���(���=��4?{�6?�>��?�r�㾵�>m�@?T�M?R�>���F���Fy�O`�>���?�����5�>��>���>L���CKI���ν���=����*f>r���C<Jv
��%I�Z	>�1�>�F>k�(�T���M+�>�_ ��K�p 6������F�)z�<�?�3��eb�>�>��>Ҿ�a���Xu�����>?y��?�8?�F?��^4��-.G����=9�>�Ν>Ɣ	><��=3��>ew�>y ؾ�ċ��x ��w?F��?��?ӎH? $����ڿ���v����߾�#�<n��>�$@>{}��}>r�����z��~z�=��v>7�=���=���=H4">z��>o���������	�����b�HS�����h���
������!��BǾ���	�C�Y'߽�}�KB�M��<�33<u㚾pN�>D:
?��?���>Ӹ�>nW=9��!��\���{��%�U���־��N�\ ��oy*��թ�}9�5ؾ5o½e꾑�Q?�&;���=�>`�(�@�e=ĵm>�>�2>�d�>�s>L�=w��=�l�=?'>��>_�>�B>�;�h��Wr�m�H���z>+�$?q�u=��W�H�G��b�)������>9c?�H�>�h,��a��KN����>d�/=������������=�ƣ>���<؎ͼ���Һ�%���7�>1��>��s>2��wv��3$߽[:>�[?~.��JH�ʪA��5X?S3S?UO?R鎽�S�>!rK>Ō�>F� ?��ڼ�L\�Z��6b�>�;:?�m?e��>���=�U�;K�a=���=	���֠4=`�=D���G})=�F��S�<r$=���=A6>S�<66���L��1f��Y�>���>W�B?6�?��>���?�P�BP�=�L#>����>z�> �>hx?tj?0�>���=�I�����$��>Y�A>n�C��Y��4�=���=N9>��G?�m6?���=􃾀YE;�=�;��>̋�>F!?a�>�>y�9�
���&��zR.��xa��f�ŵ�>h�=�eP��;�<��۾x��8��9��k�G>�3�>h��>�rD>E�5>oT�>���>@��>pQ=$�a:���1&������a�<�k���wսMn�9�B=W�N>-B�>�;">0٭=T뽑�ѽ���>�X#?u�>v|���b�<zJݾo�An}>gl?�?�}>�#׽��꾿�@�Ňb�r���6�>��[?�z{>
�-��=�=Tӳ<V�=���>T_�>� 2=�0,��t
�{�}�n[ ><��>�N ?�+�>�X���胿ᓁ�����=�>7G@<ǥ�=�/�?pNS?X�Ͼ3R��e�4�2J���]��aY�ʓ��2 �-����^�6r	��x��~��ً�w,>6�>^��?
���.�=�x������.��S�����?>�Sܼ2�>�I���1�~���;�*�L
���G	>�B�>��T>&!�<��>��/?e�O?Y8[?��?>P?� ��H+�>^>�2?���>!�<?V?%��>��g>r!�=�^�DF"��%w��m�������I=���=dh�>��>8�ռнټ�5>=�K<��!��B�<)�';X볽�&>�3�=���=�]�=�?�< ?�й=w�=��Vm����>jՑ=��I>v'����;1F��1�=�KA?�H?h2�>�������L�	��)�0G�>��>M/?f��>n+6�L��Z������;�ȼ)m�>F�n������=��	D��2��d%�>�>��=$j�=��? 1�?�z?�r�=��V�uK��븾ԧ6>�˙����>�S�>}��>4+D=���TW�T_���V�������ҽbR὚^�<�M�>5�=S�<x��>B�5=�����C�>dI�=�ػ>*��>1"�>���<c��/޾.��� ;?���9+�,�{��>���U>�k>�F?�T>ñZ?��>�b��:9��7:c�|��>�A�?	�?�J?�����B;%��=�K>�7(=�cG=�OŽ�l=�Q���&>��=o���[x���J�=��>Va�>�o�=b�C���*���@����3���z����%�.��~ھ�p�����������������]��ͽ�>�UX>��~�b��t��o�Ͼ���?��T?���=U]>]��X�� �WI>�ͷ�D��kн�,�=����A־@T���Q���d
����!�>qľkh��n��|�!S��D�>���>j2��\7��y�	��>�^�>�� >��j�d���倿ȯ���Yb?/kt?��>�#��qܾHz?��#?�_?�h����뵛=B@�>̚:?�9?�����B��J��;�4֧?�~�?�%F?� ھ�]����'�3>��>�?:�^>�̾eĝ�4��=qPE?��:?�#=Z����g�i2����?��?g{X��k�>!y�>볜>�詾�ڽRnL�#)>L��=�ˌ>�v�=�.��gɾ��\�9:'��>ݨ>�FM�&t�qz�>E��&RS��A6���Ğ&>j��p�?�i �FW�=w�u>O��>J&��T������-�z��hR?b��?7�J?��?I�Y��#{��j�<�<1�xn�>�އ>�N>mT}�yL�>AU�>��`���w��:���>|(�?/��?�C?��w�R�ܿZو�2�Ӿ��������=J�>���<�>�X�:��;��dP>r��>�J9>��(>��C>ϑ>���=�{��ݷ"��=ӿ�c���9��</>�=�̾g����cԾ��#�KY ��7���"澢�j���޽�k\��� �wx�#޽.����3?�P?R�F?��>�t�=Ѳ/�����S����j��8���r�t�о_+~;V�n�A+>W�<=�<Ҿ�v�8и�3ξ��?� ���N>�6>J���:?�=H?��V>�9�<���> �<>p�)�Ol��e��=�L>TX
>X~l<�z�>��A=<']���Y�
 E���i�>p�,?^R�����<�,(����:��L��>3�O?�C�>+��W���n��§>�(=Cx/�uxo��[��S�>�L�>��=p�m>�O�v�������>�s?�C>6��n�ھi�����Z>��?���|4n�}�8��#C?I ]?Jg�>�_�9�g>y��=獭>��>%�1>EE��[l3���>�;?��`?a?3��=AK>��Vr�q9>�R�*�<�ƽܒ�;�8Ȼ��1=�`�����;�X�=J��=��=�BI��:�Ij��'E�=P��>b"A?� ?���>����go��Js�N��>c8�>	���Ѷ>Џ?��^?��>�>����� ����'Ⱦ���>f��=�Eq��������=I#�>���=lq{?�N?�愾2�GKc�� �>�!?+u ?ria?#��>x3��Ⱦ���iӿ$�$�!�ւ�Ad�t��;��<���M���Z�-��������<i\>�>�op>{�D>i�><D3><L�>�>G>-��=*�=�/�;!�;�F�U\M=����G<��P�i8����ż����5��_�I��?��Y��ټ��>��>xj�;{����1�(�׾vk��U�>�G>8P�>G��>�{�=~���On���H��ֻ%�,?��Z?���>���q���������Q��K�>n��> Db>X�S�����ѩ�65/>��>�#?01S>J<˽k�j��f�ON�����>��1��_>���?��?nL������EO��5x�!~Ӿ�F5�0�ƽ�a���`��������;7���ྟҫ�����P�>�Uy?����P��ֹ��D��~`���Ĺ=�*�=��B�t��>(
D>ۡ��p����WĚ���<]σ>��
?J؆>c
!>��>'�>j:h?�&?�[�>�C� h�>���=0��>�[�>�?�З>�n}>�ȩ=�#>�6>��x>�Z���0�~׺��m�=/
=�j�=�om>Xx��)Ľ)��=ޥC<��-���]=�y �r�߼�=q���
P>ؾ?H�)?�z>ן0>��M�׹��mT�=���=�y�>'�Ͻ"��cc����>�e??�@?�,��l�1��(�!�Ӭ�>���>`X?�v�>��m��fʼZ2�<!��6����>�r,��j���W׾\�������>l߬>�N��LJ>�?�zF?�=&?�M���T5��@v����i�<��/��l�>/˪>3b>g�Ⱦ�`$�d�l�E(h�SM7��F���@��W<�!�=å&>�`5>���=�v">���;L��"��h��<�M�;�]�>���>F��>B!H>�1v=2{��^�����;?�$��u��P�q�_ɘ=,9q>��>�1��h�S?6=�>����E�����k�>峬?�ĩ?�;?خ�Ceļ%��=�
o>P��=fӮ��!����>"�k���/>��j>/�<�3*�m�K<A`�>4�#?�c�=�v���a���1��G���E�����H㾪�1�"&�l,��>�}������'�� T@�T$.�|�<�N���ۣ��@��h����>Ⱦ$В?!}?j��=7�d�q�9��)۾3��=����BY)�k׉��;��=��	_��&ݽ=�����7�l�!�P���y�=����m���B��%��ٟ����>�>?�U�3�e�����e>��>N�1>�T��@���/�������E?��m?�N��G�G�B��+�>�Y9?��>㢖����+}E;��l>H['?L�?�mn�e��Iņ��Y˽��?r'�?q�+?���R����vB>��?g��>ENe>?���ꃾu��=�_?� ?l�U�����%b�'\y���(?u��?����e�>o��>Qn�>�~�c]=_?���Ž`h<	)>a#�=WG�����}̾�+>�.?8E?��|=ɾ���>����3(��j��ĸ�� �=�X>/�?�C�����>ˁY>�2�>��E`����������A?�}�?hoF?�?l���'��.o�ª�=��>zy�=��w�T�*�9�?�p�>4!��[��`�(��yD?�&�?���?�V?綎�qٿQ���H���S�Ͼ�(
>���:��%>��ݽ��>�&�=B`R=	0��/>Q�>�3f>F�D>wy+>2P>澜>g�����*�/��~+���,�#�	��z<��\�E���
�S5���֌�H:� =�$=�&����6�s�=p!{�?�#?��?uLL?"�>�F�>2�o�A%�u�Z�ዾ]��	-f�� ���V�r�� ���Oz��d���lþi��t�ھGX?�.��
B>�> Y��͏=��>K�⽷�)>���>i;>m�<�Y�<|G�=T�>���>DR>X�{>�h��j����N������5�>h�o?p�=J�W��a@�oO��N�l����>�=?�S=�3������(Q�͒�>z��=,(�=T�P=�he�B�	=HO�>"I>utw>R���Z���䨽�]�>��>;�>�I��� ޾����@�<F�?�`��,G��P�S?�&[?�*?Z�>=.�>6�?~?/�r>LǾ������i> g/?2�?_m[?#Ř>���=	㎾9�=�k>�un=O��=�4'�����Q=!f=�m�[Q>��>�Iʽ��8�=���7x7��,>'��R��>~vD?2�>��>���{A�g�W�����&>=��*�>���>��?��>��>]j�=^�ܽ��,�ھ�Z�>{� >Vhp�%Uv��Ij���>f!G>��P? HB?�����K�>3=7�=}��>G�>��?B�>RY�=m�ٽ6�:����Y	���r�c���{�1���4ξ=� �8f�=��s�z�⽯�L>L��>%��>��h>�<�=��=�
�>��>G"G>P��<W{o=�q����=�+���=%�~����\hE�]�x���)�폜���|���L=L��<�r��N�?��>	����#��'U=v3u�G1վ�>�6?��>�_�>��>}�Ѿ��x�fzK���T�2��>]�?G�>�%��S>9{"���9�>���>#>�@4���B�����ù<�ݡ>Ŵ(?{��>s�w�%�_�����}���?�%<^Qi>��?�w?*�ܾ�������m8p��R�8<��Bμ�1���䒾;�gm�>%���ھ����*�=侪>\i�?D�ڽ�I#<`�þk���Ǆ��ң���<*���Ԏ>���K�\�������.�Q�=�*�=�Ñ>�-�=f�>�+?l�?��b?h�?�
?�"�D�?�k�=�>��>	�?O;
?���>G+s>^�s>��=�7��K
��Ӎ���]<���kN�=y1 >��3>�1<�0=��=��<�b��{鼮Y�<c �<��=���=��=�>�1?^$?h:>K�>j,��+>�)�>6���r>��<b�@�¾Q��k�>�q?�m?��>hw����7�h��'0���>��>�^?Zi�>����q��N"��"4�8s̼X�I>\����}��,��(.%�e�`��>L�>�>g=7��=D�?Œ?�Bg?]����f��B.��8^���p�=�l�ɘ>���>��#?��;ʆ[��|�������z�i0 �-\J�]':���N=%�>D�E&3�\�S>���=�y�= �=��>��>D�>�>��>�v=@=����߼�mI?Lk���+�W�ϾA`�F;r>�K�>� �>��2���*?C��>u�l�=2������2?5��?��?Ԭ?�uH�3��WKn>x��=��B>��*�`)�����=�ey<�e(>�9��{:3�&h �و�<%�	?��?�d�=������ ���~��۷�m�F��	�����*���ؾ�B����V�J�A�P�d�oT��ɶ&���������*4��^�/��
�t�ˡ�?�Bw?�����'�ke�����q��>��C�-sh������4�=�b��U��פ�T�'�������!��`�>�͘�/�������hg���ao�>�vY?�y"����J��!̘>���>)�=���>������;���b? FT?�~$����Q��T� ?~WR?�&?��_Ͼ��%=�N�>ˡG?��?@���t���nC_�P��H��?�I�?�B?��:�m�%��c�z>>B�?0$�>�k�>����>��S�<��6?�c1?��5=�)K�/N���l�%?Y݌?��=��:�>�:�>e�>,M��n�K�o����=J� > �9=�i+��#g���½�*>QV�>�b�>�;�KE��&��>�߾�WC�'vE�[[����[M�<V��>�(�fm6>ޫ\>a->�#��x������juP��(F?��?!�Z?��'?��Ѿ7Kؾ���H��=�>�>my+=q�!��s�>j��>R6�V�|�����?�?�?�K?�]r���ÿ2x�n����K����<���0Z>%]&<:N ���=������=o�	>ި>" �>�<0>�s�>��w>�v)>���Q��S�¿�3�����5�Z��j��P�S�H�/���nB��U"ʾ��*�k�1=5m����ý5%p�]�׽k�N��>/?z4*?��?K�?1��>}c��T��G�E�0����ҭ�����~��KF���þ���=LO�=]���М���u�>Z9�;G�(=LW�>�����"�>�>���,�>�S�>���>�/>��>��F>�z>��>#c(����=���65z��C��U�O�`*J����>��;?��)�⯛����?FJ�@��j�#?J�6?�|�>?��������=��Z��>�����=�cĽp�u>���>�X ?R6���(->{�aO�=�䓾=�.>�O�=^������=�4����6�=z�?S~Ծ{qJ�.</��F?)�7?�?�-=��C>	�>"s?��O<��޼��>+�;z�*?�z?o��>π�>j�=���<��+>��6>O��ϒ�"-� >���?��=ح��^d>�>�0��I�=�B����=�ϼ	s�=�^�>]Ng?,�'?�<�>��<9�4��������>��>I�f�6|>~P?U'?0�>V�8?�m�>�Y�;��۽'����� ?w��=�$�����2̽E�G>��>�-|?��\?�o���0�����=��@=�>�Ө>�?M�?1��>���=c���bӿQ#$���!�T�������;?�<�EM���7�>-�����R�<��\>f��>O�p>�TE>1J>y�2>�;�>cqG>��=�2�=Ϩ;�;8�F�8�L=8���K<��P�:^���Ƽ}���TȌ���I�p�<��\�w~ռf�?��?��9��j���y�^�������C��>F��>~��>	�>D>,��%bJ�ׇ5�rC%����>��Z?�L�> XB�5��=��C���<Qƙ>���>k�>�.��-iʽ�鲾�95��P�>_�?���>����n�L��~�y���$�>�!���:�=�t�?ni?�R���ֻU%�~O�!@�c�=A�;e韽��%�p�<	L������m�>��>�9�>�?F�;/�,>���ن����v����lkh=�>���>�X��C�氾�.1�q�������X��>3V[>وJ>�v�>RV�>k�U?k��>�H�>��k�yq�>��=�!?���>`��>Gv?oPu>	��>Hp�>�L�g��.ý�/8���3=������=n�C>@_>j�G�[o<�L�=��=;��=�I7�1�>��<h=ڬ>-��=p��=��?��>4\���	�f�I�@�+�-�
>�}=>l�>g���$^���t��$E=$��>!?���>�>!>�&�4Gݾ@����C��]�>�.?fK?�N-=Z�`>l�!����^����>J�!���B����x��Y����@X>���>M-/>zG����?uى?��W?(��>$�����.�g���>Nw7>�se>b��> ��>A7���R�T4W��v�`��=�9�#f$=�,>.�>'�='8.=�B�<US�=I�������!�s��B�>��?�kE?���>��z���׾P���z3?����[��6���p��ؼ3RB>i��>�Р�7(?Nd����I�8a��F����>���?�v�?��?н3�K( ����>I΄>vY�>�1�J��i����N=؇�>yf�=��Ⱦ����`S�N͔>�b�>m۽������7
��WV߿�==�NŃ�cP�����V`E�R��ό�=����=�������U��"����=!����V��4�Ծb����ʅ?u!P?�bi��,4�`�-��z��ξ˜�=K����
ֽ�ͯ�qx���Ǿ��/�&�L�=�򾅟(���|�<� ��?4��&�o���D��'�}��=���>U5�>�H��i�2������;���>���="X۾ŀ�輙��<ٽ�@n?�� ?�پ,�(��I�=yTV>�X+?$]�>� =�fN�D	'�&�>�[?o,Y?q+��!��n��W�ٽ[9�?z�?�IW?NW]�:��S辆1���T#?�K"?6�L>�X@������z���F?�Z?�mM>S�0룿|8��71?~a�?@���>��>�`?��
>C�G�B�ܾ$�����ƾA���M"?���'���,̾����=��@<3��>��b�\졾c ?��s{�+�9��躾�[Ƽ���=��p>N��8.>R��>��e>� �X����|��t㾩Y?���?�{v?ڒ�>�����z��$��_gֽ��>��=q��� u�'�?��)>�������J�*�(?��?���?��,?�H������փ�?☾�G����=ur�=�V[>�����P}>@�=��]�ퟨ��{�=�2�>Ƥ>d�y>1r\>x�>�*�=H~����&���ſ�H�� S��<���ʾ�� ����x��Մ
�=����辩ۨ=��;9�v�0�XT˾�ʛ�$�I)�>d�?oP,?��6?F̜>�G>���~"�	׾-��=��S	������徒�;X*���z<>�<g��Ȼ�p��>�k>��G=x��>+���e�=��>Q�2���>}B�>x}�>e>�N>j�>3_4;P�=���}��z��|@��,s��H�0(���D�>��j?�夾�~<!x���:�$Ӿ��+?��?���>@��&֍��k}�ǟ�>��<\�A���<�8�=g��=�uK>lQǽ�'��8ϼ�A5<��<�F�>܏=�E����=��׽�^�7�>�>,�z���H��=w?|�^?/�(?&�=t^�>��w>�{�>yK!>��>�p�>�,�>��?U�=?�?���>�n�=B��w��=�5�=�I��Ӆ�X% �Ы�]��<��={*�YA�=5.�C��C!=nh���<�N���=�=5��>��R?�?`�?��B���4��߆��*�=���>�^��~/�>���>k�?EN�>-�3?u��>6>G��t��|��g!?�z">��q��W���y��:��<�ޣ>0z?�k?� L;��3���A>}>}g�>�D!?9|:?m�>�8�>�"n<���cп��$��z#�G+��������<�?�\�`�a'�;Y� �͍��<t
^>�`�>�q>:�O>�>̒'>�K�>*�G>��=�η=xn<K�=<��N���=3gҼ�g�;S+��T<)�ܼ���%N���};���Q�`��i�^p?��?��<i"�Y�i���޾�ݐ��7�>���>x�>�z>�@�<����ZM���*���P��B�>�f?�?y�,em>N=�T=>E��>i��>̗�>;�?��������ũѽ!g>x�	?�m�>r�9��/2�P`��QQ��P�>WZ:�r>n~�?��p?"������=Ϥ�|`_�>	������< �a����T���[����	e&�z�!=Q5>ep�>���?V�n�����<������6������A�s�>���>A��=�"��Nپ�9:�]S�Cć�o�G�bO>,��>�x�=�>��&>�+?YQ�=6��>��J�j��>���>�y+?;�?�A�>�5?~_�>L��>v�?WĽO+�����<*g,��Q�<��Q=W{�=��>���=��=�=��>�Ĵ�ದ=�"�:�\y=�:=�M=�">艕=�T>�'?R?w�2���X��?�f�a���=,/I>��>�q�<�H��A��=z�=cA?��*?3�>��2>= ۾D޾�޾!)D>5�?)8?�XC>r������=��w�Ƚ�Y�<Y���u>��F���y���-��<�s=��#>�>����a/�?'4�? �T?�75=Ew�ا��
P��1>�NR>���>\��>���>tS.�
�A�G[���u�!Nƾ�Ľp���恽O�=L�>\��=�X2=@Ԁ��(k>�S���J���$ٚ=E��>���>�W<?��>�>IQ¾2���C?*���������U}ݾ�ݼwk	>�|�=E?,���?��\��fl��(���CG���>���?��?%g?My�J�~�hq�>~��>pDq>`��=5�Q���k�R����6>�O^= ���#�¾�낽�)�>9��>ٱ`< ��ھO~Y��k����N��07�Dt�!i��lоU��5{��OnS����c�Th�VP���Aս�?��(�Bbh�i���I����|?!�X?ja�c���02��x��ľ��>̜���������	�[�{�����Lr�������!���8�v���O? q��d���6��:����=�@�>1�!?qb~��0����>v�>R��=��Ѿ�^���������p}?đ5?�/��פ�����?��3?�>�S��J�s��K2�C0�>�?�?V/�Nc��ݭ��͡n�Z��?W��?�[?�,��f�/�Y�����;6q?LO?�ߚ>����j�����H?��G?�K�>�%�_ٛ��66�JM?��?����a>)��>d5>xe�5'���^��)����f��N�>(��=�J��S��,䐾#^����b>O��>�_Q��l��}��>B�˾c�&��1�<�þ฼�P�= 9:>-�վ��<>�ί>�ڧ>�0�� ��Ό�����~�?=̷?�z�?��?���d��������bo�=�N)>�;�璚�%�
?�H>>�;���&�O�2m(?���?��?g�K?�/�����u���9���I�����=BV�=�>�
i��� >�=�=o���f��=q&>�&~>��B>|��>N>�i>��=>��~[��'˿�����*I���$���۾W@���<=���ξĊ
�{����H���/�:�/��z*�0������V��w�>I�?<j/? "+?�P�>���>�WݾN��}���DZ	��[��nG�.
���d�$�_=�A�<�s�=Ɗ�`���� ����>ѩ;>��: �>(j�buq>#�>�d�=96�>٬>���>"P>݁�=��<=���;{H�=A�&=̍�>����D�r�����2B���2>��4?�:!�rԾ�������w�1�?��5?˯�>���~苿O�~��B�>~^��^`���,�9c%>Ī�>㏚>�%�%$��ӏm�Y�>3�O��~O>$�>�
9�[�E>ck׾��/; O�<]��>ݪ��B�1>> I?o�? �>?��4>�z>|jY>��0>-��=�4�>09�>��<>��?��	?#0�>�>p��=�@ͽ_!Z<L��<��n������� ��=��$*>%�<v>���	>"�Q>���;�D�=#�����Ƽ�r�>#;@?�?%�?m��.�/�9�i��R���(>�j|=U��>o*�>B #?{�>�	?�

>�R����.���B�>ȩ#>��=��p��w���))>ُ(>��d?z�?����z���=I8&>�|�>7�?�?e��>]>2�����E]ӿ�!$���!�Ee��w+��1�;g�<�ǢP��7���-��~���5�<Q�\>�3�>�yp>�.E>��>Z�2>\��>S.G>��=ه�=�q�;#�:3�D���Q=4���I<c�R�(.���wǼ�ᖽ/���K�@2<���x�׼:�>��T?���>RU���v�<E��.��R��a?� ?���>	�O��	��Xq�Z M�Qv����>��?T�?��b���>佋������u�>�>K >�G��HL=@���O�=�H>�?��>�5{�\dS�Sӊ�0���~�>mܣ���>>Ѣ?� }?� ��\4�<�ZA���R�~�ľN}���w�&�-�y�U�[�(�I��J��>���%��=��1>��>��?��<�ȟ�w����ެ�M�?%�>�?>>"��<0,B�!��CT�oӾѶ/����>j��>թ=$��>�n?g?sZ?��?�?� ��@?ʃ�=�.�>�s�>&i?J�?{��>Tr�>�2h>�</{��_��-����
<
���=�}>��,>j
�;d)=�)%=�Z<��[�����G��<��: 5=r��=ES�=x��=��,?\n>?�`�A�����c�F{��k�>N��>ʜy��C7��Gɼ��=�ѫ=��)?�~0?!&?��"��4�>�����>V��>!Q�>e��>��>��>"پK���w<z�=19�=�r;�9	���;�4F��sD>���>���>�ȍ=��?�W�?wHZ?�w>т ��Q���75��4?�C�>Ԝ>X�>s&�>��C�_�P�{XU�HWc���T���<�GO��0D��n`��]�>���=�^=6AS>���>�>���S�Mm?��Ps>#!�>
�>u�0?�I�>x�=����~5?(��+��T��Β�������=����U�?��'*?V	��8�_���\�g�%n�>�.�?���?qO�?#�L��K��>���>aҖ>��G>XN��6C,�@�G���=y����pT������?�>��i>'M�=AH��2��ZV��ؿ��H��'��m�ie$�<x%�����6N!>����Y���s��=$���	�ļ T>���ɦ�=�[t�榦�P��?�^?��:�j<��p�P�R��J���D�>*)��J6>��о��S�刦�0?r�������ĺ�hs>�F�߾lI�>�4d�LZ��Q0i�I���=1}>�?�ͨ��˾�����=&7>$�=^���������I��z�e?�>-?�����;U��Ɯ%>:�?��>G�=DZ��5!� ,�>)L.?w�*?��׽F%��+���F��"�?&��?T�/?_x��S6�i�ྫྷB����3?��?�b�>'����+���ؘ��Q�>�;?*��>c�˾�b��h��؈='�K?5�Խ~�>t1�>5�Z>�By�X!+�6�g=H���%� >��=��ý8�=�����C�\ɝ����=�S�>��	>3{m�1�?L����,���̾,@��r<>�>���>�o`���=)�?�@B>�Rƾ�Ճ�X햿��X�v?�w�? �Y?��?��㾗���Y�?���8�ˢa>���>u&��~���>
��>�����zd��q?�@��?�M?�6i�hFӿ�
��`������7��=�#�=��>>a�޽�ϭ=?�K=y����}=�C�>�>�o>�:x>��T>��<>��.>���4�#�uʤ��ؒ��[B�e ���Eyg�k{	�y����ɴ�u�8�������ʓ�5�G�!��&^>��bѾ���>I=?�r?�J?�<�>| 7>&(�o�'�
���- ���*�=���^���� y�=�ԏ�d�ռ"�>�o�H�}�����?�%����a�f��>J�A�*��<1�x=8�u=,u_>rEl=�*�>-��>O�>	��<,e>C�i�M��<�&j>|�Ⱦ�Z��؉�� �;�B�!��B�=�m?|R�����}'+�=h�f\]��o?�A;? o�<l` ��[����b�q�>w�վힻ��0z�H_�=ټ�>e��>v�½��"=��z�Y&>y\D���>��>!� 5�= ���	���>u�>�2ؾ��=
a>��%?+�q?��3?�A�=f6�>��B>��>ݳ=�I>��]>�|�>r�?�1?c�)?@��>�:�=B�_�
/	=ƋD=�8���E��s����'�=����<226���N=gZW=Ӹ�;KxV=�}T=��x�+�	<��<���>gJ?~�?�6�>2���[<�� p��r���4+=��=�}}>�-�>ȝ5?r`�>��?��>�ݽ�;o���/�>;��=�HM�o?}�/�o��=��=�aT?b:Z?8۽��b��c<�z�=[%?�?0o?�1�>S!>�7�����'iҿ��y$�:�_�*n��J���M�O|��+���.�
=�!6�<��g>�6�>Vo>��:>D�>�:A>YV�>Ui>�$K=�o�=>s�Q���zo����=֎�����<�n�]Q񻐃P��������N����1���e��6��>�K"?"h���<Ii��������v�>c��>��>D�>C�";�l$���\�͒J��ڊ����>K n?k��>�i���C�=g���`=��>v�>��>K'���-��-�����<���>:?	P�>1����Y�⻃���#��a�>v��'f>ޣ�?/��?�h���)ս��F���f�zU����>��C��Q޾KI���J��R��O��=���P�Ҽ���/�>�ў?cV�����=�넾�梿��r���;�>U�>��>��>J-�����f�&������&��"U=;n�>x��>��<�(E>�>ɉ?��>�J�>�ȍ�&[?!&��R�A?K�=��?T�!?�'?��>����9��L�������O=���ʮ<)\s=c�>���=�5Y�##C�m0�=�Ĳ=+e"=eKͽ"S�=g?ȼ*.�=^}�=���=�2+>Z�?k�>��U�M�$��CN��뎽�!*>�n>A>ՕB��qQ�)Q>^pg<z0%?yg?�za>K�J��?�����px���L>7%	?�*#?1̖>)g�� �>$��@����#>[d�f�>���������ܾD�˾)|�>�Ƿ>"��>@�˽'�?k�?Q�O?���=��Ͼ5'��[5"���^=X�>�f�=�V?Ԟ@>ZcM��69��Q/�Y�7��k����]�S}���9��gY>��o��%�<_I0>���>��S>P���]�����9H~=���>��>�)?��>Lհ< )����6?����`��Ѿ�� ���;�G��>����=/>�
V?kEm�g�h�_�����~��Á>6��?���?[��?��J<��g�?��r>�E�=i��=�u���	�c�%���'��}������ܴ�P�j�>�>X�6>�׽�	���5�ｉ���3�6!j�8j��xV��m�\
Ծ3\=K�ؾ�'P>�Kо����OҾݻx<�)>Hd����J���4�����?��?˾�w�=��[��@�3;�="?�ڂ�\>I@���A��Q��ϓY��Tp�E7�/Ϳ�8$C�W�%��V�>^pc���|���I���
��Ǽ�\�>~�>?�iҾt�����M�M��>(6|>m?>6*��Lgy�+��:�z?&D	?��H��[����>���>1�>����6���ڷ�<ѕ>?�?-j4?���Q[�������H�@`�?��?�+?PF��ܕ2�07 �}���C�>D�?�U�>�������5=��?�X?u��>R(ھA�����Ά
>m�l?�i����=�o�>�G8>��@>�HL�����o �Hܤ>�1�=�u2>Akb��T��K��	Jν��>��>gcw>�z��h�>�?ɾ��=��f6�������=�=۾>�ㄾ2�=�_�>e��>]D-�H�r��u����$��?�ͤ?��@?�Y;?91��j䃾����踏;�)>B?�.K�{Sz���>{�>�>����y�
+6�(�>��?���?�W ?� U��O�𠩿>���/����,>� 8=C<>��H���={J�<S�н�W���2�KР>��v>���>K7x>�W>��f>H�|��`!���������19�����k���N����r蔾T�����F课�Z�U೽�_���f���G�ڰ�����^Ϯ>B�?Y�4?�e?>O%->V�����p4 ���#��Z-�,W�rn��jW��*̽<7ڼ4�����E-�:!?�F�>�6ݼ��>k;T`�>\��>
��>m$>�=�=e�>H��=Q��>DZ�=�q=�+>�{<�;m�>k����ֆ��B���C����+�_>HoU?�����A�����=��羾�>�a�>
NO?|Nq>ED��B������#��>[�W��6{�(ڷ=��=; �>3��>(�=~����U=�� �:M	����=���>e5D>>`���Ⱦy���>/��>c�־0�=��m>a�"?��t?�N3?��=� �>{�S>:?�>���=��T>�{\>���>�?��)?w&$?�y�>���=�`�n�<<E=r"H�k ���mBI�����<\j�Ju�=��H=V/<z�<YT=�Լ�YT=�1=��>�$B?��	?���>�����,�$�t���;�"�>׫��}>��?��-?�н>h
?Z;F>ցB��Y�:���>��=
FK��t~��]d;3T8��>�>J?]uB?�2=�e�z
>	�G>"^?�3? �*?�h�>-R�=q<����hٿ%� ����[�����a�9��[{���=�K�����Qg�J悔@�y>�{8>R:�>�nq>�G>]�x>Z?Bɸ>(�*���*l���н��g<��$>ނ��`ƽ�Q��^�Tb�=�F˽RK�e�I���{;	��<)��I�>4�f?�J�>�k����0> �Ҿ�i��.��j�>�N?���=�$@���&��^}��|Y��81�6� ?��?�a?�~�\��=a>8�LM=5��>�>���=�� >%p�� ��W>k,�>	b�>e�>t�ɾh��Ж���N��9>��⼖�=Ұ�?�ߋ?0Pu��׼�>H��Y�-����>��������Ŝ�٬>�v~(��۾�j6��E�=�^>Q��>�Ѧ?/�,��[V� ��6��G��d����=h�>���>����|��ދ�����t���<Ť�>K��>Ʃ>e�/=	�I>!�>��)?�M%? �>���=EA5>1���=?�n��$?v��>��"?
z�=]h��Z����{��t=���1��������=�4�h>ró=rIʻ�j�<D��<nX ��.��Zڽ��2>��*�(�q>+*�=�/%>��/<��?��>B�C��i=����AT�ԅ>r"j>D��>��u=#YD����>�G��x�Q?r?�z)?���`��F�Ͼ��l=l�>�?�H�>�=8މ>�Ͼ��H�	Zr<� �=�姼`�M� '۾��ܾ��x��`>>N|>(X�>ō�=5ڑ?�Ł?o�9?��=Eu� 奿�c�O2f>8��<A��=A��>gk>P :���.��sT�[9\��:���l��f�=��y��b�>����H0q>�->�"�>ߖ����<�/��
o>���>��>ɥK?Y�>wv�����]���2?C�ӽ���]�c��hU/����=j�����`���+?-'w�`�Z�H��ID]��n>���?d��?$��?zH<�բ��U�>���>�G�;3��=9���^)��#�2���=��>�	��^�Ͼ?<��>�sf>��r��ڼ�p7��j��>%ǿ��9�����1�����>�̒d��M|=ۼ	�>���5�÷н�<m��X؂�-M8�e^��G����?p�?>���ށ�j���6���Y�VO�>�Έ�fW�= .S��%=64����q�:d{�D��d��Q��5��ߐ�>fp��邿9�O����Uu=�O�>��?��������	�w�>o�&>���=:�����_�����!B`?I?�}�j-ξ�k��qg)>U�>]r�>z��=0�2�˵j��(>ؾ#?#�I?�,�I���'Q���=<���?g�?�f4?R���s�&�i�˾Q����E?c�+?��>�W�����=�=,��>&�:?���>\Z��o���-���_>2�H?w��+�=G�>L>gh�=*��۽i�ھzB�=->�T>Z��J����Ѵ=f�4>��>�9>��%����>���M�B�G�����S~<9�?J󾕾>��j>3�>Uq(����X���W��L?A,�?ocS?�`8?G���
�����=�2�>��>���=�"��B�>Cp�>����sq�B�??�D�?��?6Z?�m�n<ԿCx���׾�s�zu�=�r�9=���<a_�<%bG��+(�d|�=2�Y>_)�>���>?4i>�*B>�h->���=�+��`�%���׈��ZA�l{���?�7T}���������MԒ��hھ��>�X%9?��=��'��\�v�ս���J.V>Z�?��?�;�>0Vt>y�=�ڱ��о�Q\���m��<!������M��Ty;^�����p�hҠ�i޽�]��C�>��n=6�>��?�j�;�u>���>j"�>�c�>kV�=��r>��=�Q���1�>w�>uЩ>D�=SE��/�*>��m�ovn�Ө�	��/��>�?����Cܸ�����q���������>��.?��{>��7�bP��/U�`%�>2�>6��=)���=Cv�>X�>�VW>2_T�(N�!�>����d����	�>{�b>�X���߾f��m>s��>�KܾG��>#�>��P?ˁy?F�?%J�YS�>���>"�>�V^>�-?��g>;O=>̚?x+?��!?J�>Y�>ѳ޾�f�=H_>r������>��IE=���=t�>	�=ZY3=ЃY>g�t=�"2��v�>��=J5>�`�<�-�>kT?��>au�>�X��X=�9���5��͖�>sk�>�|i>�3�>���>`�?�>)�/>���<�,��U[ھ@�>@��>{�b�����n���?wr>(��>|�?�Q?�U� &M� $�=�7>NWj>e?o�&?�,
?���>=�%;�x��>�RP���F�#���k��]Y�,����&�^_���/��U6#��U}��9�>���>;X�>�ȕ>;6z>�>>�?{�~>mG$<f�ÎO���><fϼ�9����&��eQ���(�u���j�h`�+,�ǤĻk�o=J�:}�,?l9?ΗI>ف���Q��GL�c��(�?cS}?�?R�>꜅>`X��3�_�0����=$*C?bD�?���>��H��^P=���=�x�>j��>+)>��%>
��W&<^l$��Y��J�>ȑ�>A!�>��T�3?1�����a>v�%>�7�ﬤ?T׋?!;�����<�5�i˃�W����!>���� ���� ��+�P ��2/� ����7���>�V�>��?%:ܾQ�������*#��S0����Ͼ�4\��Q>�8?@.��yﱾ8(1���8���W���־+���b�>%o^=@~�>i>��q=l�%?~�>_#?~��=��=�&>$0?	�?��?�v�>Y��>xߦ>gg�>�Ё=��ľ��E�FDC�]x��ߛ=�Y>��1>��s>�)
�8�=�9.�Hf<�6�=襈��E���>ޡ=&�����ݻ�H=s��>l9?yA�\u�7�{� ?X��Lw>��>7Aɼkm��-8�I�����=W�>�?�M�>�x��Ԏ�����p5ξc��=�e�>�"?	��>r��� =E���"�B@,��p>Db>I������/�ς�߆>�5�>�/>f�>]�|?�b?̽M?�1�;@�@��N���8��<$>��)>=a�>v�A>^8��e�G�Ȉ�Bw���hX��@�x9q>�$�	8��cM>���=��=���=���=Q->wD�\���9���^�={�	?��?BA?��>���=7�������I?㞠�o �Q����ѾmK"� �>�	>>[� �\,?�<
��|��ۥ��a=�AA�>��?�t�?�Zd?��D���
]>�<W>��><�<��?�'���^��V�6>@��=	f{�����mi_;ڲ\>P=x>7ɽ(�ɾdY徙�E��Ϳ���r
�~���*��:��DkþӍ2�C	��c�^�'����>׾Mg>ޮD>+'���������X�7��?p��?���=͖�wS�g ���}�Ԃ�=2�+��Y� ɾ�ㆾWR�������+{�i=�/�5��~�nT>���dK���i�o�/���h�l��="?N��V'侵���TZ�7@�=E5u<WGʾ�c�����W����5!?|�%?L|����/���c���>���>gJ>.F>Ȗ���ɼ>\�/? ?
�=𬎿	�q� �<��ư?��?"�7?:��r�+��Z���)��>�@	? �>}���U辉����=�>v�#?�)�>�پ��y��A����>RF7?�vW�L�c>�G�>Lѷ>��X���%���������<��A>�#��R=��d��
�[�9�o<rR�>�tX>��T� AQ����>� 꾦�N�1fH������1��<$V?�a󾲜>:�i>�>��(�����É������L?���?��S?�]8?-E�����k��s��=���> ̬>�ݯ=��7�>s��>�(��Qr����D�?�1�?t��?NSZ?Ӏm�'�п�R��y��������>|p�=���=���h.�9,�;7�=�K��u�=ȳX>��=��r>Y@u>�|>v�X>��� ������;����Z���"�*���k������r¾�i"�������Ҿv��qf�1��Ol���m�����Y�ٽ(t�>�>}X�>��>�5�>�|r>����[Ҿ�kϾ��ھҚ0��޾\����pྶV��{k��HO[�� ���(پv�
?� >��<A�k>����\��7�>b�O>�I�>]�>�6>6�V>[�->?�=�fq>\��>?�#>ٷ���N�\�]��u�-���T����ml>S�4?���H���@C�u�뾇�v��}E>kHQ?�^�>@�9�@叿C���]�>w�<T
i<����V�a>Sw�>��=��>+��Έ�y	�G8�O@�=��(>��&��g�=�]ƽ�pd��=���>Kw�]��>���>;?�U?<v?x���*�>��>,��>ׅ�>곆>��M>�W>�I?�U?��-?� ?�>�˾���=ߴ&>�;s�h�;!�<)h��K�3�`>����>B��.P
�9-�x�V�ґ�=z�F=.�g=	!?�=-?C�>,+�>�
�����R�ZU��5��>���>��? ��>�i)?�;?Q1�>y��>��z>1I���]v�ʳ�>�e�>D�{���R�$=��	>�Q�>�Յ?�a?`%��&\����=�=��~> �?�Xq?��
?��S=�Fh=+��NbӿU$�#�!��D����s��;s�<�9�L��֬�A�-�����O)�<�\>1�>B�p>sE>Ξ>�
3>oX�>�IG>ل�=���=�|�;��;[�E���M=��$G<ߣP������eƼj՗�6W����I��B>�����ؼ��?���>�a��Lތ��-�=B社��
�哨>�Of>�Ll>Y�U?��>�>T�r$���)�ж+�E�?翅?]��>�	$�����L=1>��>wX�>��E��T�խp���.�.�)<'P�=f��>���>s���0��Cf(���My>p>}���-�?���?h_ʾ��+=5��%���~�¾O�>]N <�b<n�6�w�	�.3W��I��w���b�L�>+x�>ȟ?Ⴞ�$^�#׾NF���怿W���l�%>���=ɺ�>���=_q��߳��MJ�\���vC����P>JA�=��>�-y>��Y?�L?y�R?W�?G��>��Ⱦ��>6ʑ>�?�>��>�!$?x��>�ߛ>(=U[|>.]�<�	>~��w����R=�&��"V>��>xE>آ(=龼�<�=S�>z佁5[�/ؒ=@ j�.�=��>�Y>�o ?#�%?�A��)�^N9����:��(>�bP>��>��>Ol�E��47�>�>)?8�
?��<R�Ӿ2AξU���f�@>s �>O��>�Y?�|�=V����ˮ������g�cC>V���P��ôE�q���Kׄ�.��8!�>ۣ�>y��>�n?��g?(�F?N`��Pw��뉿��Y� �<\��=�a�>���>?+`>��̾��>���w��Z:�"��%s�;��U��i1��:�=čJ>�.0>���>4 �>"��=����|ӼnQ�)���>�>:&�>��(?
|�>v��=	z��oҾ��M?SD��X/�����/�ɾ��"�u� >��8>�M	??�ֽ��u��)��\<�Z%�>S��?�`�?�c?y0'��G�n�Y>_�P>>�>��<��7����Fo����#><@�=��w� 嚾I����>>��u>�Bν^�Ⱦ�y�s�U��\ӿ)UZ�9�����:�?�X#5�T*�=W蕼o���b�q)����*��E� �W���=&ȡ�����ٷH����Ecl?�?{?���O/�=�}\�sQ�}E[�yA�W7����=d�޾��׻@���A(��'�=C{�j.���L�>og�Cߜ>�O�m��o{�7&��� ��C>��.?�%ƾu����i��5=V� >(fa<>�^���������U?QE8?,���O��[�뽨w>!?���>�T)>�����3����>��2?PG,?�p��ގ��4���Ĉ� c�?t��?FNM?5Z�=Q���}(=�?O�%?��>�:�P�&��訾�p�=�?n�f>v�)��O���h+�迈>'�H?N��13�>«?d�>��K�'��eD�=̕Ⱦ�j�=�!=�te��V��󧖼v�O@����=W�>An�<����>n羭�L�s�F��6������<(~ ?���}>{@h>H�>��&�)���dŉ�i��6K?ư?�S?4�5?�������8���=8)�>�>��=)^��7�>i6�>X��r��1�qe?���?�?�KV?)�l��ʿX��,f���P���r>Je>m�>X��,��=�2>N��=�$���;��>�w>5+*>���>��`>n@�>["���$�}[���l�!\��|��8��v1��;���*���l龄_�d"=k<��I&�2PL��
���
�=�~�'�%>��?���>��>!�>��->��V���J��ُ���-�#�Ѿ޸ھvJ۾7薾���+�b���7�Ѹ1���]�	? ��(}>�a�>F}�!P;�3
>G�7>�oE>�ƕ=���<��>�O>�;�>�>��=뭹<ߔr�o!>�ꈿ����rH۾��F��.�>�eL?��h=�S�6^e��P�����ܴ�8�Q?Z��>X�q�J��k�����>/�Ӽu����1��6=�M�>�f?��M>�y��H}���nܽc���搽�e�>��>���3	=� =H��<��>����>u�?��>?�\?[�?>���'6=�<�>���>�݁>M��>��>gݽ�_�>��V?u�4?�@?CB>� ���N�=�K>;D�e�l��Ԃ=��>��>��Y>���s�=�;%��Q�+-h>Q�$=�[|=��>xv>��>�=
?%��>j�>�5��G�7�<�=U�6b�>i��>���>�>*P?C� ?$�>|��>���=��?�_�Ӿ ϭ>c��=��t�)�p�`�=���>�>��O?L$�>�ݟ=�h�=�$>)��=3z�>{�>��G?�g?!_�>ޛ�=����nq$�I��>( ��6=�N���a�D�����mU��f1��c]�� �>��w>�&=>�M>YK9>~�n>���>6QN>U��=��=��N7��x�qb�=�;9���\����:,d"��cL;��P�կ��΂�SZ�)2B��?;)?�����2�ɽR��A�۾�9�>KU?��?P�%?�{�>?���?;��K��C��0?�̉?��>Ď����=��
>R	a>L`�=S�"=5��>�Ͻ��=d�a�O�`��='��>ZYE>o4Y=����"�0x澑7[>��>s}�YG�??�������#,k�B ����m>u'꽃�Y��ܲ�XTP���d�s�	ב�`S�9�>N��><�?)��=�aw�i���"������=�M��1	=��8?ͨ�=-�q�5Z��zl�z���������<8R<w>��N>I�&?Q~6?�e?f�?6�>2Ӂ�ͩ�>�L0>�s?ST�>I	?n?��>*M3>��>���=�!=��T�x��s`����)B>#>Z�->���=�
��DG<�L�<	$<t����� �=��Y���>E(>�R>"{�>��?<������M�-��7̽O�><�>�;m>�#�<�����z5=�8�>U��>��?�S�>n��=���r���e���=??h+�>�X?�w�=�m�<���-	ھ�w�=D�K>�
l���L�����Kھ"s��ޝ�=�g>3�=�m�>$�e?fw? �M?h��3�7ˉ���c���G�m��;m��>���=~�Z>@-��w]��1�m�Dt-�'.��* �\���t̤��+=x/�="��=�mK=�ƍ=��;>����3�x�=��=��?��!?�?Š�>��"=O\��l���I?be��&�F���	Ҿ�O<��+>��;>r~��?����z��c���<�\$�>o#�?
z�?%)d?�A�Ne��C^>��T>�(>���;xs@����A���S=>���=c~�/��E�><�lZ>v7x>�R��;Ⱦ����A��ܿlrs�Y:Ӿ�ج�UE��>�L�;�$����B���:���;.���=��;t茶 ��}�־�����Ȑ?�Y�?��Ͻ�����>��\�����Ă=�����8a�z�=#��u� ����v`���j���i�k�_� �>ӄo�W*{�:iu����>-b>1��>�wd?�{��~��#�CM�h�*>O+ƽ�ڔ�4���K����ѽKL?�?�Nľ��B��0�����R�>R�>,>Ƃ������>�L5?k�&?^
u�`���e����E�n�?ל�?�%=?ؒ˼���K��2����?m�?5 ?�dɾ>[������_�>�*?��g> �۾A���p�%�Ŵ
?��T?x�/�>�?�U�>��H�_W��ҽb*��ˈ=��>p=[����9���ֽF&O�T�>��>����m����>��.@��:�� ��̣S�\��>Sw��6i�=zj�>���=�k!�C㌿ʌ��)���E?T�?�wT?#�*?�� ����1�e�A��=\��>�%�>X�=;���I��>�B�>��ٺg�|��W�?1�?bN�?�eX?J'd�O㿧���k�ؾ�m���ؠ=�F�=M�>�a�&��=��ֽ�mx�P������=���>k�>�T�>[ q>vO>#�>#ۇ�%�����������Fv�xt��{� �H�u|��|.���c�=��z���XXy�Eqi��c�����L�mg7�{� >�;�>2\�>�&�>Q�y>�d�<��ɽ�g�զ��O��=+�U�Ҿ�����a���4x0��������(����_	�>��=�y|>���>+S<'\G���>�=>�~>��`>jF>c!�=�@=)��>L�>�y�>jW>-恾ڐP>,9�������þ�z�=c��>�#;?*p��V�&���j����m��:b1���?�>nRh�w_���ޏ��϶>"�=D����½v��<e��>	m�>�/�=��<�o��ڂ�_a���B���T!�=���=�}����B��D>�J
?��5� �>)�?�e?��g?��7?�{=ib�>�?.��>�FF>2c*?Tm?J�T�d<?i�s?�yJ?~�N?E�1>���$���0]�=<����n���t;mB,���E<���=��
��	�>jT�=۵�>4n?>>q>��=�-�=�"@��r�>�{?p��>�=�>�]�H 8���O���hՋ>��>�K�>=��>��?��??
�>��g>��>bi˾Io�>f{b>Ԍe�x�&׻�_Q>JϞ>w~?tj�>�"���~<��j��F�=�p�>�n?��*?�R�>0k>}+�f���Vӿ�"$�G�!��D��r�̲�;(]<��VN�Ano9�D-�+B��v��<��\>E8�>t�p>�0E>! >t�2>.U�>$OG>v��=��=)�;+�;O�F�j�M=��b�B<�(O��ٶ���Ǽ󘽏a��|HI���>�Jv�Ahּ���>%�5?��8�Le^�#�����!���t�>�oY>}��>{&?�E�=X4��M��ؾڑ�ZH�>�N�?X�>>q�����=�y�=?�=�9�='pg>��l>UnW�Y��=���}4�0�>j��>�i'>V]��h��Re!��g�'��>@�=Y[��NM�?כ?),�o�b)�����ǜ�j=�>������=j��J�_2�^�$�����W+4��5>��>���?�㣽mS����gL��1िw�c��7�=��umG?���>y�N��{վ/;B�����(ʾ'�c�2/>��~>�
F>��??��0?5SX?.�? �>�"Ӿ��?,�>Ǐ�>�ʵ>?~/?_!?�6#>L)>q��>�>b�=��gg�������u�ܺ�=D��>~��>;��<��#>�\�W�z��톾o��;�>�?=�ƨ��=�=�Ō>���=�p�>8�?�=�OY�9�"�L C����<��o>��>e�z���.�������<vV�>k�?��>�*=VGs�b߾��¾\2=��?�#?� ?���;f���E־\����,�I�0>�bC�y���*�����c��([<���>G�s>��>DM�?�h?�+0?�5���D�-���E@�B	4��{�.��>8�>�hu=,*��	,��:M���K�/y6�сA>VqQ�n�)����=�>E �>G�)>uS�=$�����X��<���r��<`6�>�6�>���>n>:>�~>⍒�&ھY"I?�R���J�Ռ��K�Ѿ�����>V�6>���N?���68{�����b<����>C�?��?��d?^�B�)����\>�=Z>S�>���;�`@�&c+�2㐽�&6>]��=��y�������:ޡU>��s>�ͽ̈ʾ��v�\��$�h�c���đѾ�Q��	`������d������Wܽ,�Ƒ>�0�� �`�*��=��3�������@ʾ���?�r?�m.>T�����(x!�b���ސ��ag��H�I=,d5����=#s��S���C��վM��<6�,�@�Ql�>�� �ր��di�����=��z>@�1?���N9��!#��M,�q�$>g��<���#��[�����Z�)�K?S$?mG˾jɗ��"�9u�=�S�>��>c	�=*E��-Qt�0a�>f�B?�)?�1���_�����Ԣ<��??��?j3?dЊ�����d����?��?��
?����@�O-K>]�?0;�>f1$�Kݕ��b �b��>p[?��l��E>r�?�W�>������M��+�h�9��>wg>!��=} K��ff��e�Ic>>�>�<�,@)����>��.@��:�� ��̣S�\��>Sw��6i�=zj�>���=�k!�C㌿ʌ��)���E?T�?�wT?#�*?�� ����1�e�A��=\��>�%�>X�=;���I��>�B�>��ٺg�|��W�?1�?bN�?�eX?J'd�O㿧���k�ؾ�m���ؠ=�F�=M�>�a�&��=��ֽ�mx�P������=���>k�>�T�>[ q>vO>#�>#ۇ�%�����������Fv�xt��{� �H�u|��|.���c�=��z���XXy�Eqi��c�����L�mg7�{� >�;�>2\�>�&�>Q�y>�d�<��ɽ�g�զ��O��=+�U�Ҿ�����a���4x0��������(����_	�>��=�y|>���>+S<'\G���>�=>�~>��`>jF>c!�=�@=)��>L�>�y�>jW>-恾ڐP>,9�������þ�z�=c��>�#;?*p��V�&���j����m��:b1���?�>nRh�w_���ޏ��϶>"�=D����½v��<e��>	m�>�/�=��<�o��ڂ�_a���B���T!�=���=�}����B��D>�J
?��5� �>)�?�e?��g?��7?�{=ib�>�?.��>�FF>2c*?Tm?J�T�d<?i�s?�yJ?~�N?E�1>���$���0]�=<����n���t;mB,���E<���=��
��	�>jT�=۵�>4n?>>q>��=�-�=�"@��r�>�{?p��>�=�>�]�H 8���O���hՋ>��>�K�>=��>��?��??
�>��g>��>bi˾Io�>f{b>Ԍe�x�&׻�_Q>JϞ>w~?tj�>�"���~<��j��F�=�p�>�n?��*?�R�>0k>}+�f���Vӿ�"$�G�!��D��r�̲�;(]<��VN�Ano9�D-�+B��v��<��\>E8�>t�p>�0E>! >t�2>.U�>$OG>v��=��=)�;+�;O�F�j�M=��b�B<�(O��ٶ���Ǽ󘽏a��|HI���>�Jv�Ahּ���>%�5?��8�Le^�#�����!���t�>�oY>}��>{&?�E�=X4��M��ؾڑ�ZH�>�N�?X�>>q�����=�y�=?�=�9�='pg>��l>UnW�Y��=���}4�0�>j��>�i'>V]��h��Re!��g�'��>@�=Y[��NM�?כ?),�o�b)�����ǜ�j=�>������=j��J�_2�^�$�����W+4��5>��>���?�㣽mS����gL��1िw�c��7�=��umG?���>y�N��{վ/;B�����(ʾ'�c�2/>��~>�
F>��??��0?5SX?.�? �>�"Ӿ��?,�>Ǐ�>�ʵ>?~/?_!?�6#>L)>q��>�>b�=��gg�������u�ܺ�=D��>~��>;��<��#>�\�W�z��톾o��;�>�?=�ƨ��=�=�Ō>���=�p�>8�?�=�OY�9�"�L C����<��o>��>e�z���.�������<vV�>k�?��>�*=VGs�b߾��¾\2=��?�#?� ?���;f���E־\����,�I�0>�bC�y���*�����c��([<���>G�s>��>DM�?�h?�+0?�5���D�-���E@�B	4��{�.��>8�>�hu=,*��	,��:M���K�/y6�сA>VqQ�n�)����=�>E �>G�)>uS�=$�����X��<���r��<`6�>�6�>���>n>:>�~>⍒�&ھY"I?�R���J�Ռ��K�Ѿ�����>V�6>���N?���68{�����b<����>C�?��?��d?^�B�)����\>�=Z>S�>���;�`@�&c+�2㐽�&6>]��=��y�������:ޡU>��s>�ͽ̈ʾ��v�\��$�h�c���đѾ�Q��	`������d������Wܽ,�Ƒ>�0�� �`�*��=��3�������@ʾ���?�r?�m.>T�����(x!�b���ސ��ag��H�I=,d5����=#s��S���C��վM��<6�,�@�Ql�>�� �ր��di�����=��z>@�1?���N9��!#��M,�q�$>g��<���#��[�����Z�)�K?S$?mG˾jɗ��"�9u�=�S�>��>c	�=*E��-Qt�0a�>f�B?�)?�1���_�����Ԣ<��??��?j3?dЊ�����d����?��?��
?����@�O-K>]�?0;�>f1$�Kݕ��b �b��>p[?��l��E>r�?�W�>������M��+�h�9��>wg>!��=} K��ff��e�Ic>>�>�<�,@)��&�>������W�T��u���m�-.>���>{R�}��>�>�U!>��
����̉��wA�RW5?��?��Z?�6?���x�־�J���>d�>� �>���=-�y��AX>%�>�A��Z�r�_��3?8��?/��?3MW?
�u����D����z��X���Ͽ=�#���/>�9�0*�8I���  K�%;��a(;>�y�>'<�>���>�=>.Y$>WN>�5���q'��(������D6��$;�����_轾��A�:��b�!�^���x��~a:L��b�<|�
��r�;oB8��ھ ��>�J?c�>К8>���<B���R��w+l�Ŋ�B�~�tN4�Ӗ:���n���9��9��Iq־�۾���[���&?�� =�@=E�>��U�} �>�v�>M��=$P�:���>j�>���>� �>��C>u�1>���>Ca�=;�{>Xň=����	���d:��Q�p�;"�C?Ra]�������3�0s߾X���B�>$�?�S>�'�������x����>�G�M�b� ̽!��Y�>̀�>�V�=� ǻ͞�/�w�s_�=(��>QC>�.k����� ~�=^&?C^��⩾K�>�_l?�1?.�	?��>f��~1>�8�l��>�,�>wg�HO�z�?_�f?��?�7�;5��=�L�??>xb>����!�<^���~����=�[=�2ý<���@��x��꺄>��>�C=��*�
�*l�>�;i?�7?�8-?O�Mc{��S0��u��-�>�y��C�?WP+>��-?�:?�6?��=� ���+-���9����><4�>����j3��!6>�Y�>wɽɓ?R?Е}�J7 �b쩾����>yK?A�?���>�c�>�U��� ��ڿ�����	��Cؽ��_���<S����bM�˦'�7�r�i����l�=���>bc�>']�>�#'>��>>j�;>�'�>;>�(���=�h=��\=�t)<��=-؍<��#=B��<
���t�x��T
�6G������E���
߼��K�E	?̅�>r�ýdÄ���+�~���z5���>B|�>�t�>�=?Uf==����A9�T=X�JVP���?�\Z?��z>)#�5;=vb�`W�=�#? �N>��=�l�=D`�U��h>VT�>�B<?�1?]��=����|��Y#��>��ս�k=�٪?�<N?��e�Ѿ�q�	��剾cM>F��� ��'�T�,�� 群-�P����¾��<��>Sr�?@�_��"4>�X�������X�<9���U=9�[����>l�>;~��mޑ���A�%D/�������"���?�#>u4�>�>!2?^�r?��?��?ZlԽܙ�>��=g�>�%�>R�?��>(d�>c��>9n�>�x�=����Q���|��4V;�[�k�y=��>�	>��4�:��<Mz=�lY<}v��q.�����;~�W=
1=���<m��=��>��
?��!?G���d�������7��P�=�wI>R`>!-	��b,����<�;>4D�>-�?n4�>vs�=+8��8��lu�^j0=v�	?��5?=�>X@�d�H=���G~�,�=�>┽e��������2�����Ҧ>'Y�>�2|=����?�F�?ZSY?!y��م���}���(��)?��A���>�
 ?��>�I������;`����������O������<���<t��>���/�2��7?C&��,��hC�$V%>	�ۼ�'?��?���>
^�>
� <t)���"��'?����P���Q���� �BtH>L,�=������X?^�P��.��=ŷ�:�����?{��?��?|�?��慳�v�?��>f˽S�����ž���hl½![�>me����m��Օ��H˾�Ǳ=�+��0��bݝ�J|��׽׽g���e�F�����Mc;��������������惾0)k����<��,���漽�p=^����i����a��췠?r?�ru�����*�Wwо)ѐ��❼��{�>�L��q��r0���ӾP��
��]6!�S�ﾠ���+q>I����喿)��_��L�s=I �>�ה>� 0�gJe>r�\�6L���>�>�;"�$K��P���[��8WN�?I��?w�ž��9�t�U��ؐ=��$?�?d�$>��t����=�:�<��e?�yS?G���s��}���J��+�?��?��%?��y�=8/��iM����>�k;?e�?-v?���
w��z>���>_B!?�W=?A5��#'���%��5?Ϳ�?�́��q^>�>uYH>tˁ��O��(�<w_�����_�=e�=�>�Vu�^7���#�=�!�>5�>r�̒��I��>I��`�N���I�� �"��=��<{�>w���L
>��<>q�>t �Q���-�����J�C?ᘱ?�sV?�x5?B=�8�b�3��g>��>���>�q�= ���+ܡ>��>~��k�J��]?-��?���?��e?{s��kݿ�����Kg���X�<H":17@>�(��l�;"�>;e�=pb=m�>"�>�uk>��>s9)>�s^=~<�=�x��0�*����!z��x�:������ǚ��8�A���X��<�jÓ�b4��}��Ar�����VO�~�>�?���2Eݾ8�>��$?��!?��:>S=���~�=�@��2ož�<�zT��O����djԾ���5v��.=�ד��#��^��x�8��	?F���>��> nξ/(?��<P�.�.�>!����N�>���>�p?}��>��>�	�>��s>d�{>G��=� ��S��M:�[4Q�q�;��C?�]�)g��r�3�}߾}f��:�>��?�S>0�'�������x�^��>8�F�!�b�X�˽���2e�>m��>_��=�Ȼ�����w��f�=�Å>&->uo�f�������=S&!?YP�����ؐ>�Q]?��?x�>��>B�;`wh=g�$>�K���>���=J����>%�O?d�6?��>ӷ<�g������E�9N:�������=�'W�j�>�o��<J!=��ݽ�/1��_� �>���=����t0��Q�>�G?��?���>�^����G��K<��f�m�>6�8�c�>��>�?��?�?�$m>`��a��)����>)�%>�Wj���U����eR>�N`>u.?��?���=�5�m�>�Ϡ�>��><��>��0?��>��>�"�v���GϿ�w�c^�����r��q��Y�����;:����7-�^�h=7IR>Ӯ�>���>���=�~;� �=/1�>�U$>2�.�B�u=��=�A>tsn��R:��O��̖���]V�S6P�X���6d�<�b���!�R͙=������>C ?�	=5��=NI����	���\��>��>���>���> �;>kZ'��w^���7�mVg��)
?AD?�<�>�g���-�=��G<N��<���>�٦>�"�=��}�F<ƾ!�Z<k��>�?Ne�>�W��ch������8a�>���9>���?J�Z?WW)��
���O�ڹ-��U�����N�;�!��0��l�H�����	�����E���5���>q��?����P�e�*�'������r�2x��/&�>�~>ͪ�>���=9����(�0uL�E�0��Iɾ>BG��ά>�f�>\6>�%�>���>�%f?�55?��>��>Jy�>/8�<l|>��>m�?��)?}�>0�=���=힏>�:>���Jt(����:�]�����=�6�>��=֌�=��u����<�ؒ���r���=�kV=^��< ��=����d�=�n�=�?��!?l��=z�������-�*>�O�=~YZ>{�4=���a��=�Q>���>��?���>x�>М���r޾�d�T��=<��>} ??T��>V��
	>TY׾0�@�ׅ >��	>��=��¾�`�����9i����>B�->uV)<.~��`#�?J��?$�>��־]W}�&���l;��)?i0���S3?ü�>	I�9�7�Hp��t�81i�����K1~�ȓ��%�ޙI>ؠ,>��o=�l�>�t�>$��=����W�� +�SpL>���>�i?�S�>L>\\�F�Ҿ�a˾�2"?Wv��@˾`�;u�%���!�n��>1��,?�=�;?�����z������8x�:"�>���?���?��(?���l����{�>�$?k��=�覾?셾[�����Mg�>6f/=-f��0S��+��bH��F�>?������������(����N�h�@��I�]B���;��|s��nd�z�ƾ䃌��#վ�N�� ���M��=�Q{�4Hl�~��pþ&�?ˏw?ԁ���{��Z���׾ q8���O>����A>-���i�s�2���ž�c�(�aK���,���G�>����m䔿N��H����.>�M�>\��>�%�ޭ�>��s��>z��>���=�j�3����ߏ��Z|��Hm?�Aq?�����f���l���3=�� ?n��>��=B��t&_�qfj��B~?�E?��o>��˴����[�φ�?�(�?�T4?n�V�,��t���%>T�E?�>��>݌����G�\����r0>�Z?�w3?&���{Y�� "��M6?4�v?ÇY�Ej^>_{>���>D,>�y���]��K(ҽa�$>� �=E\�>U�E�z�m��TѽQ>z��>���>���>����$�>�
��X��oJ�;�þ��h>u��>��>O�U��*>�{%�>S��>xN���W��Ǜ��SϽ��H?�:�?H_3?H�&?��Iǘ��;�>�k�>�>���K7�=q �=��=���>�𾍑M��5����>`��?�'�?�p>?�-��o�׿�ݓ�Ϲ��ܚ��JQ=�e=��>B����>_��ֽ�����d=���>mP�>�`M>��>���=��>�Q���$��ݩ�Ξ��d>�n� ��&�F��#�!�Ǿ-&�~羏�n��{ͼ����4Wl��.������U<����	�>��?wȷ>�Z >m���j�_��]	�A׾�F�o��<iK����d�׾�d!���?2ʽ��ľ����י�|�>��z?S�D�T���I�?��R�|�>�V>��(>���>~`�=Z��>Ye�>z>�>�u$>�o�<{�M>�Qo>�Mz>5ň=ݣ���Ѐ���:�MVP�qx�;�C?	m\�8�����2���߾����'%�>�
	?&T>l'�˪����x����>3qK��L^�"Ƚ�9$����>Ġ�>Ѽ�=Y����j�#w�&7�4R�=� �>��>��|�惐���Ӓ�=�2+?���y��G�:?6D?8<?i�#?�t3=tㆽ��>�i\� �?c��=7>߽�þM?1j?7G?�.>2@t<���P�<~�h�����a=��}��R�=�}~���=�$�����P<V��h>Pdc>�����YE�!DP�[�*>\��>�%N?JdC?3��>F��(���:�E�M>��>	�-����>SW?�G?3 ?*$?nZ#>k�l���-�RN��>��|=��Z���G��^X�bT~>x�>��H?T�>m�#<K�ȽG���&m!>j�>^<�>�??u�>-�>��	��1�Wѹ��<þT�'��9�-7_�v��\=���<��0�����������<�a�>�F?h8>*�;=>b�>j��>_�0>Y��;�-a=,E�=
��<���=�� =Xη��/->�_=v� ��������(��+�q��$=4�=?~ܼ�i?��?6��� 
�<���(}�����>��>���>���>���=�-���rO��:���1> ?�B_?��>�eK����=�DN�;�'�>짛>�U�=����:�Qܧ���V=���>��?���>�7��g�K�}����v��>&Q��(S>�n�?Σa?r�zF���D���2�`ф�Xx1���<kc�)�W=3�����¾��V|Ҿ���X�>��?�^�/�=�Ӽm����������,>�F���=��=y0߾Z��ۻ`����:��%��rb�>��>�Ϝ>�l�>Sl?��Z?�$!?�m?�N�����>`�>�8�>��>��?=n?f��>��U>(X�>���=�!̼s��;#S��s;L�?����=m��=gY>5�F=J�c=�B=�~-=	��p�޼H<"=r��<�Y�;��_=��=d_>�	�>��?�P�<"�<�����2.��d�;,F_>6�U>������8�k��>XW�>��4?�k�>��%=�徜��A:ؾ��=s�?b	>?�y�>~N���>s��_n����=]X�=�jv�9��j<�Յ���t�;_��>�p�>X?B�f�*=�.�?���?���>Nܾu�����(�7��K&?�e���D�>zs>�
�̬�����]3`�𪀿�ؔ���a=	���[	����='* >���E>��><M>D�ֽ�H.�=ۉ=��>O?�_ ?�a�>�df>]�l�0��E����;?�tO�F�Ǿ�M�����G$���\>�����S:�q"?K'���"!��j���%��E�>\W�?�?M�.?�D������D?�<?�,)=_*N��ǘ������Ⱦ��?�P���f���������>4(T>s+�.�Ⱦ�����
ɺ���G�����`侚v���񹾨��ܤn�0^��}�����Ⱦ ]��+	���q�v���0���u�C��������?�?rO,���*����lZ�A�\%=0�ؾ-V�=FҾZ����ݽO��׾V������^�% þYaa>�V������S��[N�RL�=��?�z�>E�0��W.>@ W���H>g��>��=(�	��M���Ä��T��f�m?���?�_;%.2��^�ox=y�?�?hYb<0�����O�->��Z?�\�>�e��5��H���`ܽ�-�?Tq�?pD4?��μDp9��q�=��>*?h�>9�6?��.�
;:ߪ>���=��P?KeP?<cl��"F�'n?>_�?c���>3��>5+>�	��~��=>TR�lU���>=�QE�#�'�8��C�t��˻��>�;r>ϲ��o�g�v�>X���WT��|>��ı�������];-��>$���X�}=��'>��=:��~c���o����ýpF?�!�?�NC?Ӂ)?���>_׾@<޼v��=�6}>l�>�@%=���yQ>���>q��א{����{��>�+�?���?`�T?~�6�ϿO̒���G�����e����\"�=���o�>�?�=lS��]\�k�>QO�>�\�>vl�>~*�=�>/��=R=��"#+�RZ��v_��k�B�R��Aꤾ`��I�G��.��{1�8'羼n���!��02�+�/=��Vz���j=iʾ��>^	1?/�?�d>���W>��E3;���"6��ϙ� �;�=t�#~���{�=<�:�<���� �4����"����>N���-I>�Y ?i�½��?�s=y=��>�^�>ւ'>	��>t+�>���>�y*>(lK>�>�,{>9.�=(���+���8:�k�P���;nC?s^�J��I�3��߾F+��Y��>��?��R>O�'������x����>�$F���d��"ͽ�T�{m�>��>�޻=�'��Q��cy��5��t�=i�>�O
>�������U�<="�?�Eо������v>]i7?͟>?�?r&�>_���h���>8Wn>���=���=R�#���>a�C?)3?v�>a�=I�����=A�:�$0�1�+=�댼j>ߩP���=�F=f[�=��<�@�<��=G{A=�g�<H�	�%�v=�&�>�Y:??��>��>�cM��E?�'rG��
��[/>
׌��1�>@��>Na�>i;�>m:�>n9;>�m�#uҾ������>O�#>L�Y��1e����]�c>�ru>� O?�/?C��Qx�@�Jؙ=Y�>W ?\%?���>��>��ս'����Կ<R�^����~�uG��e��=\C�8�Ӿ�?>K���� �>�T�>�TJ>}M�>�
>;� <��=�X�> �w>x�s:>I�>�S>=�ح�Fz�=�2��C2�<]4j=�]$�}6�y[߻��.��[ۼO�_:*�?���:��I�>65!?L+w=�|�=�v���F��3��)l>fB�>^�>i��>�>�#�2~c���<�y�ڽ���>�D?k�>.�~�0�=1���7�<�u?&�>��8>�{�<F2��{lľb��=���>�L ?���>VeX�H�n�}���s�����>�̽<E�=D*�?�*e?5z�d����?��:�l���K*L>scW>���s��P��l�l�|Ĝ�i����^4M����>gب? ~߽�>��ɾDՠ����� Ԍ�	 �>�W=��>��A= z�qh�a�L�j�'�l�ھ�� �`��>2�=>t2z>"��>���>^�d?z�2?�{�>=��=���>�e��U?��F>M�?Vb-?L�>�Vn=��=�O>l��=D*�~�:�.�=�Y�;t��=��>��>�P=�B�=V�=GT
=��s�v��<4��=~}$=f�
=
��=㥅=���=u�?)� ?|Щ��Ӥ=�/����h>�B>��->��̽�2����=�P>��>)�?h �>�W>P�þl���I;h���{s?.�8?���>&x��`�=]�;�5t���=!/W=��R�S���� �� �����=���>b�>^��)����J�?��?�?�c�#�x�����=Q�?.?������?��>D�/������޾p)L�)�k�h���o���޽�2�:�6=0�=t_�=��W>�`:>��z<�s�!��PI����>�H?$}>��>�r>i><xl��C�ʾ�0?n&�mf��c�=L;о?�-��H>�鯾�]�6��>��6�B��+���*���k>�<�?���?m6A?��*�k1����>	� ?=+>�E���濾�q��ٌ!��g�>�� >�ѽ��4;ڌغ�R}>v����ྸ��*d�豼�}E��}�����৾�L�����%��.ʾ�J<=$�߾.�f�co��N��;6=L���t�T�>?��u���av�?ؑ�? P��v��`2�l��!��<p%I>[oþu��>%c��u��C����۾X�kC=��=�"����R�>C�l����S^����Ŋ�=R&?\��>{����>g�o�1�t>��>�~>�G ��č�����r��Ya?=�c?
�����Ni�=S.w>�l ?��}>��=)Dӽ���HU>o7?�]?Z�w>�΍��f��Շ��,�?�1�?k�/?�0.�K9��Q ��H�>*�R?��E=a�?�m�=ƾ�+=��=�H?Tp#?�����v�+�?Ès?����̫>Ti>�G#>�T<ڄ��/w½ ��=e���}��=֖��Cs���+J��!�=(��>��>�ѭ=4�ھ�&�>������W�T��u���m�-.>���>{R�}��>�>�U!>��
����̉��wA�RW5?��?��Z?�6?���x�־�J���>d�>� �>���=-�y��AX>%�>�A��Z�r�_��3?8��?/��?3MW?
�u����D����z��X���Ͽ=�#���/>�9�0*�8I���  K�%;��a(;>�y�>'<�>���>�=>.Y$>WN>�5���q'��(������D6��$;�����_轾��A�:��b�!�^���x��~a:L��b�<|�
��r�;oB8��ھ ��>�J?c�>К8>���<B���R��w+l�Ŋ�B�~�tN4�Ӗ:���n���9��9��Iq־�۾���[���&?�� =�@=E�>��U�} �>�v�>M��=$P�:���>j�>���>� �>��C>u�1>���>Ca�=;�{>Xň=����	���d:��Q�p�;"�C?Ra]�������3�0s߾X���B�>$�?�S>�'�������x����>�G�M�b� ̽!��Y�>̀�>�V�=� ǻ͞�/�w�s_�=(��>QC>�.k����� ~�=^&?C^��⩾K�>�_l?�1?.�	?��>f��~1>�8�l��>�,�>wg�HO�z�?_�f?��?�7�;5��=�L�??>xb>����!�<^���~����=�[=�2ý<���@��x��꺄>��>�C=��*�
�*l�>�;i?�7?�8-?O�Mc{��S0��u��-�>�y��C�?WP+>��-?�:?�6?��=� ���+-���9����><4�>����j3��!6>�Y�>wɽɓ?R?Е}�J7 �b쩾����>yK?A�?���>�c�>�U��� ��ڿ�����	��Cؽ��_���<S����bM�˦'�7�r�i����l�=���>bc�>']�>�#'>��>>j�;>�'�>;>�(���=�h=��\=�t)<��=-؍<��#=B��<
���t�x��T
�6G������E���
߼��K�E	?̅�>r�ýdÄ���+�~���z5���>B|�>�t�>�=?Uf==����A9�T=X�JVP���?�\Z?��z>)#�5;=vb�`W�=�#? �N>��=�l�=D`�U��h>VT�>�B<?�1?]��=����|��Y#��>��ս�k=�٪?�<N?��e�Ѿ�q�	��剾cM>F��� ��'�T�,�� 群-�P����¾��<��>Sr�?@�_��"4>�X�������X�<9���U=9�[����>l�>;~��mޑ���A�%D/�������"���?�#>u4�>�>!2?^�r?��?��?ZlԽܙ�>��=g�>�%�>R�?��>(d�>c��>9n�>�x�=����Q���|��4V;�[�k�y=��>�	>��4�:��<Mz=�lY<}v��q.�����;~�W=
1=���<m��=��>��
?��!?G���d�������7��P�=�wI>R`>!-	��b,����<�;>4D�>-�?n4�>vs�=+8��8��lu�^j0=v�	?��5?=�>X@�d�H=���G~�,�=�>┽e��������2�����Ҧ>'Y�>�2|=����?�F�?ZSY?!y��م���}���(��)?��A���>�
 ?��>�I������;`����������O������<���<t��>���/�2��7?C&��,��hC�$V%>	�ۼ�'?��?���>
^�>
� <t)���"��'?����P���Q���� �BtH>L,�=������X?^�P��.��=ŷ�:�����?{��?��?|�?��慳�v�?��>f˽S�����ž���hl½![�>me����m��Օ��H˾�Ǳ=�+��0��bݝ�J|��׽׽g���e�F�����Mc;��������������惾0)k����<��,���漽�p=^����i����a��췠?r?�ru�����*�Wwо)ѐ��❼��{�>�L��q��r0���ӾP��
��]6!�S�ﾠ���+q>I����喿)��_��L�s=I �>�ה>� 0�gJe>r�\�6L���>�>�;"�$K��P���[��8WN�?I��?w�ž��9�t�U��ؐ=��$?�?d�$>��t����=�:�<��e?�yS?G���s��}���J��+�?��?��%?��y�=8/��iM����>�k;?e�?-v?���
w��z>���>_B!?�W=?A5��#'���%��5?Ϳ�?�́��q^>�>uYH>tˁ��O��(�<w_�����_�=e�=�>�Vu�^7���#�=�!�>5�>r�̒��T"�>��q�m�V�y/��Vg����媽6�>.R�eK�>�2?�Ɏ>�20�������)O+��zu?�F�?+�H?V�,?l�#�Ӧ��ݰu��K�>�0?�B�>�����׾p\�>�'C>e�����|�����?�>�?���?�\|?9�s� ߿�ɥ�F��U�����B>H�u;�ĸ=oE9��C�:p$>��_V�;�>B�>��4>�F�>�US>�W->="%>�?��E#�}������S<�w������(R�|�m6����=�'����`���Uz���!��~��O���-�<RS��o��>�� ?D�?�,?cf��P%�b_�_��K�9�U�_%x����jB�9�ɾރ�=eS>;)�� u���;=�5�C(T?��>�hż�H!?[������=V�>ZĈ>�n8�x�>��=���=l| >�W>�8">��|>b�̼��>�.�<�c���m��7���&��=�Ő>�F?��m>�s̾�Kc�f���4ۼN$�>�0?"��=�A"�YF��E^X��?��E�wf���|��l�=dz?���>/��=�mF=)����b�ݙ��3Ӓ>БG>�4>+?���
���ڵ�*Z�=���>B�Ѿd�=vj>�f"?�u?��3?�R�= �>�P>Ձ�>���=��P>��U>RΊ>*�?�2?��,?���>�߶=K/^�?�9=xӟ=s�W�Ny��ݖ��w�����b�<�O��1=�T�=�E���k=pj=SEм�=�J|=[,�>L?+�?;��>������Q���a���E>���>��#�y��>�n?�4?:��>��>��>j��������I�>"�~>�Jh�� ���O�<S"_=�|�>��?Oz`?G������ ɻ����>�},?��7?�_?�R$>�Id�'��9����̿B���n�5�>X�w=T��<d�g�tA�_�;�n���}=,B��J�>tL>ġd>`\k=��=i
&>
	�>��>��4>���>�y�=��.>��U>�$>z�>u`">Ti�=v�V��u����O2A�x��3*(���Ž-s ���>�y5?l�k>:�>A�5:���U�,��W >�NC>;9�>*��>KVH���	x��)GG���B���,?�d?�v>?�/�.d�=ː�&>ܑ�>̱g>c�O>�C�h����LK�͆�>˒ ?��>�*0>�8��2��{�����G�U\�>�q�=���<�Z�?Ouq?�A��-<��JS��/r��Y��Z>�i6�,���S�Gt>��=����������*�=hp�=Y!�>/��?�)��o}=������j����ʾ]�����㽙��>j���i��ı�C���,�����=�$>�K�>	�>���>IK�>�vV>o78?VT?�8�>̆=qn5?@U�<���>��>&��>��	?�M�>ZN<>q�<=����$o�T����v_����=��2>�����|>��g>�Ku�)�=�H�<$�=�8Ľ�9>&T=lQv=�2=	BT>�^�<�P2>*?�75?���=ϰ��IB=�+澕�½�B�>|�?�_^=
?��'����OZ>^%�>Y�l?>�?�%��'���Y�������=�?7j:?��>B����j>��6�XP����>���>'��p῾b�������Gn����>���>fH�>��0>T�{?bh?�Cc?{��=ط:�bߑ��B�Z����A>��#?C�>>>���zq7�@��c|���E��3�mk<��ɽg�t�՚>=�8=훹<6�=kBE>�d">��>����&
=���>�ϭ>��>d/�>.�:=;���[����;ɾ�~'?�>�`_��L� �'#���-��i=-=��_���Q�-?u�Ӄ���檿�p=�\� ?�0�?��?��m?H���}��>�sL>��$>q�=��W�<�ڽ'@:�m	X>H�-��`i�����B>�_�>���=����AʾFt!��E���ڋC������M�"����,�����������Y���/g=���Υܽ�����P<R�k�)��cg��羭)����?�P�?t��3ྈ���`��^t�K�>�Y_���o���;X=�-��e=r�|�7�W��C���/��پ�;�>۟��(����{�S8��z+>\��>۝1?�������ļ��
	>��v>�3�=��߾y����%��`Q<�I�Q?@�'?9����G�f;�M>l�>Λ�>��>�wվ=u꽨.�>T�?d6?�::����������Aƻ��?��?:?���s _�U��b:�:[L?��F?V� ?\��o�\�GŽ�T4?C�b?�e?1"�����|��w>#�?���B^>_VN>+�(>��=4
��R�G�c&���>���a>��a=�7C�@�M�:FK�S�׼�o>�>En�S.���>Gd復!G����*K���Z�
�=��>�㡾l�b>��>O�>�4�����M���%ʽv�?��?��W?�;?����?��d#���6>��>��>�z>�}��d�>7�> ���=ti���ľ}?!I�?���?ШT?�E���ؿ� ����d�9���m��>���=zi>��o���>\SQ>\m�3�=gr>e�>Ch>*B>�5:>ZS?>@7�=��~��*�Z����ل��$(�O��I߾$0���&�����P/H��������� ��4B�(�R�e3��%�c�ʻ7��J��>P&?�Z�>��>�sd>��%>����X� �c0��?�(�V�*�b�
�ھ�V���Q7�Mc?=㒽R꾫@���^:�W`[?N���>>�c
?p���D>`P>��>4���?����N>΀==��[>b��>l\P>�B�=�_>���;Aބ�X(��x�:��``>��>�6?��
���5�b�����l��{|�>9L/?Ӷt=�m6��p���6L�s? �:�h6�ѣ��Ԗ�>��?o"u>�-�=��ν��<���܃��w��;o�>>R\�=·���E��m+�ّ�>Ă���ӏ>�vp>:� ?x�{?�J?.h=s�>�>E�>��*>U�.<�"�>⾧>�?��;?�Y-?	-�>��=w)��(>��>��
P��L0���;�у�MN �����m�i�h?�=N	��J�
>��*>b�M��*>u�>�:�>*�C?�l�>�>���[ZV��]Y����=FB[>n˜� 2�>i�>�>'P�>���=���;����j����B�>}�l>2�L�w���a]>�b�>��>��z?#�??0/��������<l�>ُ?<?�IC?ǉ�>@Km>n���-� �޿g[�'>��&���$��3�=?����e���=�ž~��>���>�Ֆ>_��>��e>��F>�o>I�>+f>$,�����=�6@���'�Pi�=�{�N,:�w�1���i�6|ɼ�(����켡+�����<��ܽU�B��/�=L=�>x� ?��=� >�Ƽ�#���4�9>���>[��>運>�iҽu)E�~4|�:ZI�*/�H,�>��[?A#�>�$���R=�o]��j�= �8>�{�>.��>��������N�zyB>�?O0?�*>�4��E8������B�G�#v�>j6�=h�$�ξ�?�?[����A��0�4�+dl�W&����=�j��Sw�������8,��\=�/L����IhQ��49>^�>{�?�ľm�:>*X���+��(���巊�S��=~�=�c?K�h�R,��4Ͼ�����娽�ԃ>~�>Z�=�m?���>U8�>h�H?��>a ?	�μ��8?��H>�1(?���>/2?�y�>3�
?H��>�N=�S'��Z���K��	<���S>�@�=q��=�+U>�3>����=��=ߥ.=2Fs=@ ׽�v>��~�Re<Y������=уj=sj>�0?�?�wb��^Ľ��L�J'��A>��>��>r��x���i3׽e�>�L?��<?��>�Gs�4�s�sA��ڪ�i��>���>J�H?N`�>��5�2	=\W&�J�微��=��?\V��O���@�?�H9$������ڪ>qY�>[�">@b>g�`?I!*?�/\?�����>���{�-qZ���1�(�=���>��P>u[���+���_�熿�Y�"[9���>�l��_��;*Q�=�j=	lK<���=�� >��>o�E<�ސ�ߏ=TU>�m�>M͹>%�>�-=Õ�<��u��[���19?�uv�|���=���<K��xsK��y��0^���
�>Ƭ��Ԍ������C�>���?3-�?K��?�^���S���K>B�.>�1���(��0]��G��}ِ<�/?����оL���f�ν��>3Ĳ>�o�������V�;�/Ŀ��E��c��WȾWR���򾟤���ֽ�ξ��q7�[P���6�����U˽�(���	���i��w�����ʩ? �?l ���3�]�h�z��{L��s��>
皽4����Ͼ�G�6zS��������ȩ�ǒ#���X����BO�>8ಾ�珿8֓��g�fU>���>�VM?�E���d��%���$C>}NN>�:�=��;t���'�������iI?? -?c���.��oz����>�X?Pg�>�k�=zS����8�7��>��?uX?��=":����x�L�"~�?��?��'?��ݾZ|��"���^���G?�~%?0w?ɾf�������>��?��?X�"�����0t8�A��=QG�?�Z��ͤ>��>�"�>��T�����j�A�t��L8=_+�>0@>����������4�=��a>O>�XA�%�S�_��>�̮���I��
�������D��5�}�>C� 0�>P�>]�>��D�Yw���g��$�����?rm�?�[?:??md�͞��۞p��2>��>�{>5岼�L[��1�>68|>)����b��S�h�?��?Dl�?<�j?j�`�c�ʿ�_��Ꮤ��V���>}J�>��;>��:��7�<�+f=1�+>�3>�>�y>P��=jbM>s�<>`� >�m�=^h~�� ��o�� s��NDF�J������s�+�?�#�]U��{�O�z����]�ώ �py��%�0�ܘ�<3o��ģ>��>��>}/?%�~>�NB>��ȾB����ٽ�?]��c?���Ȕ��Hnu�T�K�i�ԽgY��S�̼AZ6��K?�T%�<p�<e��>¡�_7,>��>\��=%*�=���>�I��3F>��o=c~$>Ko>�u1>I��==j�>�=�c��3��/CA��{">y�/>VW?�7>��^�)���'��� ���>�y�>��k���%�n��4�9���>�^�M����	����=F��>�ط>�>ͨ�=��~� � 1���=�Z�>�PX<�����L*��J��)�$>D��>��ܾT��=�Y>C�*?��j?��/?G#e:ae�>�DU>c
O>���<��Q>�p�>��>Ā?O�?=|0?���>�f�=�.O��G>���=�显�޾�C�>�1�༐K���k5���	>�}>~��<�#�=$'���q=���>'9=;?J=D?e�!??��>%���_�j���O�s�`=tŉ>���=��?髻>���>_.�>���=�`@>JM)�I)���h�^��>�)>��[������>���=��>�c?��9?k����5��=6J>���>e$?4[?��>��=��Ҿ�>���࿪��Y0N��΍�m�=�D%�T�W쑾=�=ӎ�=��_�K�>�=>�h�>�֐>TN��`#>1d>���>��~>|�=ۉ>f�н$sj�b���?CR=5!x=~T����	��	&�y�	�T~�� �<=�o��躞��U=0D�����>Y�)?���=��1>X����������X>��>I�>/��>���� %���^���.�(6�+?�^S?`��>��`�Xٗ=�ɼt�t=�#Z>P6�>��>����ީ�Z����= �??@}*>�vQ��2��sՋ���*��ܳ>�E�=�<<�j�?o�t?a������&Z8��\�m/��&�=����֓�r��V�&�؈�ơɾ;Ⱦ�/:�#�
=v�>��?�zj�w��=z��D䖿��o�S����>W�=���>��+>�ֽ7P���"�U���F �c�1>�i>RO=QM�>,�?~%?��h?n�?g��>��8�(?��;��?�{�>#!?�>���>Z�D>��f>( V=rѼ����r��-dc���4�=P|>���=Ȋ_�����	��
>wH�� �<�jq=�&����W<���=��e>~4&>�3?��!?��^>�]�=�X>T����g>���x�>��=�7���k�����>i�?�/^?:�>��E=����d,���/�S�>(�>��9?��?ghH=�M�
�,��&Ͼ0|>&	t>2Ԏ�;xc�v�=�<7	��~���>�i>�L>%�7>x*{?P�U?8�Q?��l� �� \��*��(��˖=��>^�>���=& ���3��{u���Y�N�3���+��@��.���>>DD=`#>�=��>��>�����<`PE����=P��>̯>���>�"G=���9�� ��#Ͼ9U>?:��t����<�� >/M�؅ƾ��g�\���"b>�TE�'ɘ��C��U��%�?��?Lw�?v&�?p�ԾJ�	���:>�1>�ye>����L �[@��.T�����>�����7����)7>ia
?w9
?�O#����[���F��]��ޱ(��򯽙������'�(��[�^�"��n=�Ŏǽ����� �����d�F�Aɽp�?�jz׾��⾋�����?w��?u�R=�E��DQ��/��vξ�8�> ���{���Dƾ��`=�-��]��7���,$�?u ��\������>q�)�!����r���O�����>I>i�:?��;��cȾ|_��(>递>3��=GE���酿�j��ז��f0,?!k\?0�Z!(��q��)�/>Ȕ_?��?�+�>|���s퇾a�N>�A-?mY?���=	h���w�h��<���?���?��?S����a��կ��澾Fl?�P?�kF?�Eɽ�2��k���m?{|-?,�>+�'�c���"����
�ʇw?��%�e>Y�y>4��>������Trv�m=f�*�R�E��>�̃=�ݷ���i�Y���"��g�=F�>�WK�F'��3�>�.c�V����]���?����k�cj	?�r�e�=��W>����6�Y�Eh��ƼH�(.�=4�l?NĬ?�5'?�IO?�L3�!�8���)=��>�:�>�[>�8*�>D4?=�>D,��\ҁ�÷#��?���?D�?Ii?�g_��ۿ	>���@�����9>Md��.����ֽ��>8�=����;�$�=H��>��3>`;X>�-'>�[�=0�>	̃����3���݉�Շ)�G1�{������+)��{�2W�O֖�����W`��	̽5���P%�ݳ��v�	���P�Z��>��?��?�h?�a>j����Ծ?��`������m��)#׾ŏ��K�̾�e����U�'N$��A���i<][/��Co?��n�.`�=º>) �	ˋ>��`=Y]�=LWm>�l�>��D�%�>ٰ�=�M�=K7�=�A�>E( =J�>DnB�13�ᔸ�,ێ�Bz>>�e�>G�3?+¾���>�*[����̌����>V�?���=�`#�`�˿@�]�?�l���#�QQ;I��>Q�=?�p�;�p>mT���� >�M=���N[(�CD�>i�>�V��2��Y;�� ��g�>C�ؾ?J�=�|>�!)?��v?�I5?���=G�>��U>�&�>�{�=�L[>ԏd>AC�>O?۔6?�2?�N�>���=9�\���Y=�"S=9F��g�l��"��Լ<�
�j<�O���k=-�~=}�0<y#E=�6=�ï��!h<c�	=���>��8?��	?5��>us��p7�ӣ��C�v�_��=�(��= �=mڴ>���>Ȇ3?C�>���>S0��ھk�>��A>\X���n��b=��=�=�
~?S�2?����C��צ=�p<=�>�?@�6?�x�>��ݻ���
�Yп��ѾF�+��qO�Z7
�� �z�\<���`�	
Z�ܿJ=B3>�zZ>�L�>lF�>�	>0��<���>y�=�s(��7�=�!�,��=��k>���=�?>�H�=0S"���=��U<̵u;�䃽aj<x&�UM�čt=zH"?��?R�>�	�&�]���%��5���2?[I?�$?Y�?v�>m/�j)m��"6��I��B�>
ER?٥�>M��EK<7�j��wP��Y�>��>���>�:�<@3s�%����9=�X?2u>?d@�>,�^�:1���	�������>Qә=�eƽ�f�?y�W?��Ⱦ��5�v�)�L�o��/�M�J ���k���߾�������AF˾^�ž���1j����>K�?��J����=�J�������,������=5�D=,4�>��Լ��s��о:���o�9�&��=e�>��2��I?PrU?2�??��Z?�~e>m�>� ���O?g����a�?@�[��-�>�%s>Ys>��=�x >GR�(�����,�情��!�=�����V=AlL>r��=Zk���=C�C����=/��=���0)=�~1=�P�=w�=�(>6�?�\-?�}�=�~�=V�k�0Y�=A�}<��<>^ �C����$=AH�>\�>9(?<ߟ>?`�=�𺾗U�qD:�� ?0,>4�?���>ʳ������*��W�R�!;r>�8�V�ل=�z�Ⱦ�1=?�>"�>�u���i->藂?�N?��!?�02��R/��HO��j���f=>=�r��?�j>�G�=ǫȾ��!�l\T��RP�d0���(�$"�����=>�� >' W>	Eq='8=A����G���m�ʙ�=�j��XH>�i�>F�?�Ga>�c�<Ot��I�ϴ4?0-���j�3`�A�*�hv'=+��jJ=�<�{�K>�;�	���$����#��T?ۦ�?�\�?q\X?���-������=�X�O�>��C��;��=��M�B�>�AD=���,/�����>���>�2>��F����} ��I^������J�`���(��\�?��c���=Ҫ߽�>��Y<�����E<�r��촽r�&�9�ս�6�̬�?��hv�?m/�?~+$�
RJ�я��n2��U�oa�=��p�� ���s#�Ua�K����R׾�{������1����E�X���?��>��ľ�Y��@t�E��\�>%j�>7�??��h��<�t��p@%>��:>��<>-þ��`������a�$u=?��?���6�׾�t/>T�>��>wE(?����qӾ̾�:���F?��d?5:K>򪒿VR��y�K�,�?��?��9?���}�K��^9�ÿ
>sM�>�)4?��>՚ؾZ���a�s�\?*t`?���>��@�V��smP���>ɝ�?7����J�>s�
?���>�U�����S���ͽ�JM>1<;?ˌ<m����jR�"�U���;>�:>��>T}ǽ�7;��e�>���vR�� ?��R�J�U��=�ݽ>1CþA��=��>�)|>a\'�.<��˅���C�0�U?��?�N:?�?�ݠ�w R�̃��ŽZ>0�>QY�>0V�=� �>E�?���De��l��?p��?�i�?��0?��u���п0Y��O�9�����_�=O
�<Q>�Lۻ�/D���&>�L��_-��J�=0��>I7>%��>�>�n�=�]a>1��R��&���g��6Z:����&���ֽ]�%��=ڽ�9��ܕ�R�ƾ�M��o�3������?��� O�9N_���>@j?O�	?��?�b�>	�S�t!���#��<���	��T���������	
|�ݤ��j�XZ�D{�ě��J���Ta?a�'�U�>>�ȩ>����S��=A�>�>~���E>�*5�6�M>�]A<5�J>�zp>m<J>�L�=�>���<�W~���h�<��(Ľ.9�<��8?�	:;N�c�@�#�H���������>զ3?\N�>��%��/���-o�OW�>�|ǽ�9B�,@+�*��=���>ė�>�M�=�k1��ⰽ|����e���e>z0�>�+E>�'սɸ��*���>Dq�>����"Խ����=1�?#��?Ǆ.?�	�|O�>x/
>^�>�mW>}'>���=� ,=��>9B+?L�L?��?��=�0-��`���!s=����h�/�����5���H=k[���ˀ��Z[<�xk=��[=Eѯ=E7�< o>��ʲ<�$2=�>i�=?�%?g+�>Y=�����l��=�N%=���	h>wc0>�X>��>��>�>1�=o�y�8�E�>�K9=\QV��&��:;��`�2>S�?T�x?�X?U&����=nb^>�$�>��>�l?�r3?�-=�a>9��=�n�|�ǿ���Fݥ���<FKj�h`���<��žF��>�T����G���<>�=<>$>ރ��$R��>½
��>��l>O謽f)�>�#<�{=D]�;$!���)�=*��<��=fB�)ػ�����=��l>��+�յ��r��^@	?���>S�K�<-B����*�ܾ'Yb�H�>X~~>_?�
?]�>���ң����0����T� ?Z?�?�q��q��$9b=�B��Q�>���>��>��w}�Ay^�V��<Bs�>��&?���>�=`��0��Tb����h�>���<�x=�?P?�A��q���)d�	H<�1Z�v�=nꊾ3���w�T��$*�����:����s��^���zQ�>�.�?m��#�=&jʾT�����U�wW��ϝ�<��e����>K-�=Y)��:�����lx���.��.<���>P�B��6H?EQ?�h�>$D?@�>���>x��=�?�Ȟ�&BA?	>�/?=��>.��>���<�(���*��m���'=��𖾩Q%��C��6>�"3>]/O=@4�_�����n�G=�"ļ����Xq�<硦�g�=�>J��ۭ�>��>�,?�n9>�ؿ:�s�=	����Ds=�&�< �>S9������r�s=���>y� ?*E?n5�>a�C�Ȏ���<�a� �8S�>�S�>�A?���>lNƽ񁸾D���|��b�>rw�=�&龌������[���H�ų�>f��>�2>�>6ǅ?~�N?��A?�Ș�����x��hT������)�5�>n[=�< =@�Ŭ1��{��z�g��A�����=�.�W$<��>��=1k&>\�=�[�<�C=쒩��b5��s6�w[= �>U�>��>jL=��=#�ľQxɾ-�)?U?��_�n�(���Vy/���*=(�>$U�>��>�����k�����j"��
?l(�?���?��?�����݄�}@I>�x?=%��>�=3>����;�y��>�>&���H���<*�>�s?i�c�����G>�1����H��Æ4�ͬE��lW���������a>���|�����CT=?f
�ɏŽ4O]���������]u��9¾�4�z߭?0��?��`��i_��;|��%�KY��Q�>*�����=~���	�<���$����ɾ�������	��?�a�>o�}�8]��eX�&�Q��!�<�g�>Gk?=	��=ԗ��Z���=|��>F�	>�ʾI-n���g�5�"���c?�X?��;�"��o<{�O2�>x05?6�>��U=g���4Ѿ�2�>	/?�x8?�*�=Ɣ����Y�=%�?�	�?��P?����MZ�j��)�1=D�B?�?��ȼ �轏�Ǿ��n=.�:?�O*?G{N>�����H�"ٲ�(�4?�E?���K.�>ٿ>��A>��R�W�q�� ��Ͼ�<'�ü,�0<8�4=7WC�V���-�=Ρ>9%�>h��� �	���8��8�u�]�=���k��&�&�)>>.?�2�/�����ӽ�t�>��4�lJ���k�e�羹>?���?ZMK?��?U���|��wL*=�Y= ��q$>Ǌ�D���*C?u��>�L�k_��D��?��?GR�?�3?�P�����Ņ�Iʺ��>����= �>l|>jur�P�>!��������� >��s>��!>PX�=�WX>7s�>yP6>S̆��������`��Q�^���ݾ���G�� ̾lS׾x�1�h���}�Ǿ@l�d�8�D���PDG��;��y��|{���PT=	ݹ>�.S>⏾>k=i>�=��~��h�DM�@���5K��h��0��Ic�>2� ������'����߽������>�]��P	>��+?��=�z="��>13�ė�>���=�u>Z�>x�N>�p>�{=�8�>\��>ߐ>5j�=}f���[�p)��Φ�\U;=��,?��q��}����A�j����6�/��=F��>��=c����Dt��Nc�Y �>��o���住�D;[ڽ�:>XՆ>�;�<-�#=�|r��`�<�
��I> ǵ>U�>D��;HȲ��XQ�3�=��>�۲���>=&#>%��>��d??�/?���=�S�=n2���R>�_�=� �>���>��>��(?E��>�q>X��>@_>�9��� �<���=Fx#�9�����`t�=MC<�?�>ΉM�8)>���]�f�A��<�(���ͽ��>\�>��0?�Bp?t]4?�?�;>=J(�G�I�q\��^W�>ڛX<�� ?͵j>&h?�I?�7�>�b>�ھ#3�������o�>�>�~o��ƅ����6U>EW�>e�Q?���?3EO<ho��B��p�&��%>���>?T+>$!2=��I>��ȿ�2����Y�]�e��Y������y���j>9������>5E;��.4=���X�ֽ�6�=���=�7�=q��>���=	m�>y�>+%u=֒>K�8>�>ܡ�;p@���gB��f�<�S��#Į=�OV>N��;����i��:KIO�84D=��(?�8?�}����������	��(�����>��>�?�P�>3�> }��	[�Di"��l��?��H?���>m���:>��b��Q=�]�>+N>��?>6Cؼ�z�"�����Q�>���>��>lk���S�	TO������=�>����˜?:k�?^�r�h�-�M{���k����ž��9>�~z>w��b���F��N�r���������J��0��2��>�9�?�����6W>p� �)*��(���d���v�\o�=��>���=5��=�CS�梿��E���9����M�j0�>��N���=P��>���>��>?>P0?2)?��>JI>tk��� >`��<��>�k8?�|!?�߼>$�?^N]�-�=5���LU�m�=qf�=��$>J�>�Ғ>{�=&�K���!=\�=vOU������a<��=�;=�%=?�<`u�;?�-?�2?���=c5=>5�
�Lէ�4��=�q=��>��޽�~���8߾+`>��?g�	?���>+(
>o%;�q��4��o���?��)?hc�>��>�s�=���҅ʾ���/?^�㼰���Kw��h�0�>?��>�G�>S�1��>��?��y?�N?�>`�@�xM���+�-�k=�8?�?��?�U�<�_���P�h�{��!:�?�ھ(����o#>� h=�e����F>#`>�9=�[�=?<�:LR���(��c3>��>�@�>���>�>~��=/�����,
Q?`k��n��Ǘ�/aվ�h��.	>�E>t���G?����dq�Ҳ��<??�&N�>,��?	�?Y?M�A�	�ٽ��j>\�>>��>�$���d�܏���b���>>�/�=|I��
ɥ��J��@�|>["�>��+���D�
#��Yǿ��P�V׽������������ݾ.���o!���8>3��~&�v�ݾېھ��u�)��Ԩ�A$�:���~?�'?��W>��p��I����<�Ӿ$��>w^)�>yJ"�_!�sD���Ƚ�㼽�'k�"��@�-��
5=���� ���}�b�C���>�w>�q;?�d�-��7,���=���=M_�[s�鳥�w����=W�P?�$�>x	
�`�2�O�k��r�C�?�1�>�x>�������H�^=�7?W; ?~ �)���J政�6�<g�?6	�?��?�fֽt�.����{� �;b?	��>4��>Z���:*վ�%T=�P?o�5?�>��߾=Y����2��>�Zf?ǂн">���>���>�6zw��N8=f���:=u&a�ܰ6���%���ҽh9Z�=E<>0d�>�cO�j7�����>�c��wL��F����j����<~&?h澨�>"V[>�m�=�&�;����;���Hͽ�R?�V�?�R?T�4?�f���T�}��eW�=���>�ʰ>�!�=����>K��>Y�ؾ�]m�~����?��?ګ�?�OZ?��d�-줿/���Jgþ�/��01=�D�=@!u>���.�=�.o�}yL;Y�+=$�@��!�>+�>0��>�Q�>�j>O�}=�υ������ƿ7T���{��[����84<����~;I:�j2��i�=��,��׍���c��ܒ�[�C��Ӿͮ��S� �
��><�>P�>�$>d��=��>�z��#C��$������|���GL��R�����<��:i���Խ8��m꾇ّ>ھ�<u�>��?��>�����>6�	>���>���>'=�KĽ�uW=�-�>�>���>t�=ey�P/Խ��o���h�"�l�#v�g��:��G?.ս�EA���_�3/�,;����=�.?��Ӽ�y4�a�J�v*��f�>N�ٽ�j���)#>aq�v�g<w�>_#=)�f}_���ؽ�G��$od>��&>_�i=L�=�✾�)��B�>�">�������?��y�>kKu?���>��3>�[h>�0>pˊ>r�>��=;1-����VS�>,��>�HA?_0?@m'>Ç�a�D=�p>��h�Ī�����<�᪼�i ��ʣ< ��=�H7:�S�=3�=�ʹ=�{�<=�s=�ؼ�?ND?4�?�?D�.=E�룾
	��-ܓ>!!��'�?�1�>~,?���>_�?�S	?�<>����*n���?��b>;hI���f�K!;/~��p�>]�s?�:?N;�����T�^=���?/>��>�
?�?fU�=���'�Xܵ�g*F�'+6�]�O����=�1ٻw�¼����ڃ��ae�+o�=�b�>f��=�Z�>�8>���>w֟>���>"�O>���=Tt�=h��=J�=��f=}Z�=P�����5��*�;�R�=[Z��]T<a�I�.)���j�4��<7+z=
!?�v&?�X'��?���qj�g���gLr���>�?c��>8y�>q
a=ny�ݘK�.�����2t?J�]?��?2���`>�e���Dɽ��>͔�>n�E>1��<��ý�� ���Ƚ�%�>�?>�>lٽZ[�� W�O
��L�>-q¼y�¾_��?g��?�ƽ��v��R����r��> ��I�>��>(��=��t�&���!������)���y�V=���>�O�?=��$*�=���������YͿ�^V��0����8>?>`�J����Zy���~��ݾ*}_���>xÂ='U�>��?qw?��Y?6?J�	? ��?N<�=v �>�X�>f�	?�?i�>�i>[g>���=~"a:�L�hӃ��1�<Q/(�d�=_�>�'(>&��<z�>=��<=Z?%<ҝk���	�a��;e��;��=��=��=�>��*?�Y�>d�=�I>a�&�2y��h�=�->�Kڼ߸��o-�i��� �>�8)?�4?���>M�V<Nx8�������
�\1F?wH?[Z	?o�8>�t���^�󑲾�Z�=��>/��K~�= �����{O�L~8>r&�>i)i>���>�s�?��?MO?�f�>(� ��D��|����S��W�>a��>���>�Z�>���=��My��ؚ��o��%̽3}�l7>�S�=�/��d>��T>\�=�@�_��	��=�22>�i�=���>���>2Q�>���=+'>��1�����j?��%��n��������żfN�>� J>V >
�
?�Gy��텿�Ą��L"����>T��?E�?N�_?r��پ�D�>��>�s>V��=����8'=4k{�%�J=�v�=S2���䳾���<L�>p�.>a����:�̕���hA�ϯ��h�T���ʾP��J� �U�~�'���{��=Û_�Uo��#���dp�}���7�Xއ�h�==M�"aG�#���kU?~�O?v˻��	��P'�c������@L>?��t[нT�پ�9s�&ja�*��3��,B��*��)��پ�m�>M�[�ڼ��ԝ{�y)�n��c3>�H/?:���-P��p���%Z=�$>�l�:j��v����	��/��	�V?�68?x��v����׽e*>E�?��>�M>y2���\���E�>�5?�*?�'�K;��y���:�n���?��?]m?�� ���$�����zK���[+?T��>���>"wR��_�ֻ����?�?
�U>�1�aLd�i����	?�:W?�_���Q>�/�>؇�>�O�������ǭ{��>�$�=]����Jҽ��\��=o���o=	]�>�ь>��'�����r��>�޾�{H�"�D�H^���I�KU�<6�?���W>W�|>P�=>Y)�������$ķ���??D:�?;�J?O�>?C����!�x>ཧ�=���>&Ϯ>�y>I�F�>c�>u3������^ �[p?���?S�?��Z?��p��о��燿�㡾���Q����2>�-~>DjH���'��e����<=`�<|=�!D><�>��=LH�>.�M>��U>б�����0����������¾�t �p���E�վ�Ⱦsk�8���a��ӏ�AOȽ�s�AL�1ⱽ���6"���Y>E��>�Q#>.x�>��d=703>��+�5ժ�%m=�7��̊��lþ��$�
������B��<ێ;Vl���Ǹ�(��4�>�/>{�ҼS�r><n�=�w����>S��>i�e�&=�>�<8>:�"#�>�QE=vP�>�!�> ��>��+>=�ؾ:p���w�U
X����=m->�z?W*;W�9'
�������l?�q>6t?u_`�8�s�Q}��6ق>+0=�Jڽ�AV=�Y�����=�Ӣ>GOS����8%z�~}���H�:>O@>d�7=qg�<rNv�oa�u�<C��>WV���D>��>5�??ܽt?�2+?j���e3 ?�l�>6H�>~0��ۗ>"��=es>���>Ӡa?�?�D9?+n�=3Ώ��p�=W��=��;��H>m 6=�˽䇂�Z����=��f=$����=3
Z>Y�]�j����HT<�=��?neH?��,?.�?�WX>u4;���U�$}��'c�><��>��?�D�> V?�?x�1��B�>l#E>�P�d<��C�>L�"=R$u��U|�䯾��>h��>�h�?��U?�����!�E%��E�Ś4>�P4>��$?r��>�<�>��<,Z���ҿ[Q$��"�������.�;�8�ewU�P�H9x�,�J���@�<ƒ^>+Ņ>�m>w�D>M�$>�->�5�>�H>��=S�=c��;��yYE���T=Id�&`<��I�/����^ڼ�����j��;�F��D5���	�z樼6?���>{��|L���&��L�hRW�u6�>�ڷ> R�>��>/ܮ=���[�\��ξ��9�3,�>
za?��>7�i�={1�q��=�[�>p�?�XT>����h�2��=��x"=3�>7~�>zW�>��o��\��k�"P��"�>���= UX�F��?c��?�����3q�>q��:�˿�<M�.�ǁ�=)�D��H��Zƾ�P�G���W8�����=o�>XU�?lŽ�\*>�82� ���-�������� �����e�?WS�>�W7��<s��ħ����n��r�=���B����=)�>X�>��?��k?�4?��?�?	�@�>sV=B�?ߛ�>im	?��>m��>K�
>)��>N]>��>S辽K�c���=�0<(��=�>��
>�]�<VRx�S�Z=r3T=�D:�](8^�L=	m����Z���=?��=͓�=��?@�?G�*�0l�����s ��LB>X>��G��jH���߾�G��=^<ky�>�M?>��>������En���)&���f>|K?0??c�8?���������{����=�k�>@�\��~=}H���پ�K!��}>�]>�s}>(�>v��?p��?]j? Q�>UR��c�������e���->O��>k�J?�=?Q�ӽ!��y�f�͞8��T:�����������=-E�=C����q>W\�=�e~���=P����M�>p^=QyT����>u� ?;@/>'��>���="V���̱�
�J?�R���A��.��L�;a�<�wJ>өA>�K,?�o�}�d���}�:��s�>���?"C�?�yd?5�B��$����U>��K>oJ>�<*;/�P�ż���ob*>Cٺ=+l{��������f\>�7�>��ͽ�sžn��Hv����m_�����sE�=�Y�"�¾��S�9^&=1+	98m߾��I��*��Q��D��l�=j�վ�;��]�|����b?z�?�߻=Nx���z��_ؾ$K>�m���G<�Э�9r��
��mOԼ)*� <e���8�VӾ��"� )�>�[�}	����|���(��Ȗ�v�<>�\/?�rƾ&���Cw��o`=cn!>��<���)��CQ��K���'U?)�9?r�꾀^��u��7>�s?��>-�'>�ړ�>���7�>4p3?��+?V�ܼ����� ��I�[�?c�?��?K�*?;Ӫ��q)�%�̾���;��7?� ?�I�>�܄�2���&-$>�Z�>>G?�8�>�)���~����e8?Fix??����M>���>��>��f��g�`�6=�쎾�~3>��a>�B ���Y<~VI�X��cK>M8�>5?*>���������>Y���-O�R�I���
���+�%Z�<��?���p�=Q�i>W>>2�)�����]���k���L?|�?GO?�8?Z���u�=s���5j=(��>Z]�>bĦ=���[�>�S�>,n���o�.t���?V��?ӆ�?iZU?d�j�&I�������������=�=�">�eR>�=��;>�����K�{����Շ=�&�>��>Jdl>��c>-Y(>U�>8-���@+�`���Uj����)���׾�_����呱����b�/�����߾��Խjs�ga�<�\��;�WY��$g�6�=*?���>σ�>f�ǻ���>����G �i�=��J�r�Bg���Ⱦi0��!;��뇾�t�m�������1�/?&�>�n>@��> ��=w�>��>��<��$�=�Ѧ>rGq�{��=�55>C:>�J�>&��>.0%>SJ�>`f�>�Պ���{�Ɍ�89�:�qv�x�t?k^�=�� �������u/u�O/���23?�a�<����X��נ����>�P;��<�=+<~����>N�.>zo>W��{���5T��0L���>��>C�	>�a=<��!���%������>9b���Ѣ>o�>�'Q?�P?�"-?{��|(J>��k=��	?$�>��>oHM>$���B4?9�C?ˍ=?)A?�ٵ=�A�#2�ޫ��P��!���%�L<g�{=Fx;:���=�P=Mz�=�8��9~���k=,E;=Z��<����BF<��? �F?�?]�?�B���,H�%�,ݽh��>ZiG����>!�>X�"?�?���>_.���=��|�f��~��>o=>G	���4��W��JH�>'��>I36?��m?0
v��	�s�]�ݒ>J*�>�;�>�#?Gb?�$>���=b��D���j4�W���2�{�9�A�;v��^��O>�{��[߾ ��pD��k^�<'U?�@�>s�>VQ�>�Z ?��>��=o؃=��=K���C��r�=�m�O�9���=z)��Ľf"�ٍ �6YP���ͼ�%��3�2�|��>�?!#��㯡�C����R��j����>"a?E��>���>�?g;���u/����P$���6?rQ?/A�>5Ɛ�ȁ�<�Y��חn�梎>d��>Cv�>Έ���]�d$���j=���>W�2? b�>_���J,�/S�K4��V�>�j�=�L��͢?�?�ᄾSBܾ��W����7�d��<5��=��=GiF������.�;�!�����9&̽���>=[�?`/>|R>��:�Q݁�TĿ�sQ� (�΁��o3�>���=��B�Eڡ�l$U��5���n�䢇>��=��>�y>i��>y3�>_A\?�S/?���>�A���=.�rs�>z#�>(�?H&?���>~+`>	ժ>/�E>�G�>���H*#�G��i������<}G>��s>��H8��m��\c>zc	��1���`r>�E<��=}�Q<j�<J'�=?�e0?��::<h0B� �u�+��=N��=�ؼ=�S>Ѳ1�a�����>FF�>��?�/�>��e�q��)��k��$g�[Ӏ?ʘn?v�>?O���ۮ�?q����M�>	=�>
����	���c��	�
���>ݺ	?2>�>2�>w�?Bn�?��Z?�-B>a�u��r�b��������>8l�>�X>�A�>'�����7��^He���B�N4���c5�I�O����nW��>�-�=n�@>��>M>�ɗ<��d>ؕ>N1>ڔ>�$?��>�f=�}���ڡ�{DH?X1��I�����D�پ볷��ͯ=O�0>Y ;M?�4���bw�����H�Â�>%�?L:�?�6V?0;���Ľ/�U>g.&>��=��`W����B�lb=��" >q�>m�������!���I�g>�b�>/(���ƾr����)����d�2K�N��m�ξܸѾ�^����n>�"�т� ���W��W���%O��R6��g�����/~��q苾�S�?�̞?ٲ=9`6��}n��[�4/���J�>��1>��۽���Gm=�Ї��5�Ћ�."
�����ed�$��h�>Z�;�C:���ix���0�������:>�d3?�W��Ҽ����CJI=#��=����}0�����*����н}�G?��7?gӾ<2���^�mF>X?�8�>��6>�u�$ ���~>"�&?��,?�|�	ǉ�]>��=~��?�9�?�?���
��*���1=S�S?S��>Ue�>��r�1�۾�!��[?3U�>�;�>;�,��f7��w�Z�>�n?"�o2(>L`�>��|>��J鄾+�`�Y>h��R>!Y>�8��q�%�W�4�/���	>��D>��=ƽ^���_�>�����j3��;�a��V��8�w=�^?6��)e>Ir5>ޤP>�w'�$��Vҁ�!۽�?F?�ة?��4?=0F?�NӾ���������)>��>��a>�M��5�>��>l	־������	�%?L��?�	�?��O?՝r��8ֿf]��%���붾��'>��=C��=˵��[ �=�W�=rH?<�Ea=�>%o]>�f�=Pz�>f-r>��7>�E>EV���*�#¶��윿��;�,������35�z��V����
��6��?þ�N��	
���
=�>@��SW��v]��O����d>8/-?�f?c�?�'<\��>������Ǿv��=M�^��l��?����ݾ�\���}u�`�(�^�l�>J?��'t�+u+���	?��?=t�>���>�j>dʮ;�6�>
pb>^CT=z�>�p>�G�=�0���I�>��>�y>��<U��>f�=��z�o���>�0��8�>��Q>�`?k����ٳ�d;��*
��lQ�Z�?�tX?�
�>�z��� ��8*���.�>��'��Mr=����{�>��'>�����S�����	\g��a����V=�D�>��>�s�{ھ�Ͼh�>I5�>y:���Wg>�͢>6�0?zID?��?�e���>�%>�g�>��>���>w�>�!�]o�>{S7?�:?S*?�+�=m����R=�"�=��̽���<E�>TZk��oe�����)E����=�$���=��>�>�<�J���E����=���>`V6?���>�>(Y�����(4%�Ҹ��> ��寝>�b�>�-?��>���>�_>�=>+|==Ql�Ѹ�>�v>8%Z��l����Ǿ�iU>j�>e�?t?����?�=����|yN�bܠ>d�*>f�?s*?EV>�=���4��)�9�x��_�/�Um���8o�S��7G��?�ɶ=Rپ����=���<�ڋ>�?d�>���>��>G��>.�:>���=jɇ>��	]�P�:��M=����2= Z>m�`= ��<��4�����ý�N�q������=�?br�>�M0����;�S�.O���?����>ٗ ?X�B>b�;?�aI>3�O�[�,�?��7��(�=?��r?;�?���?�$^�r�<��>�u�>T�=��ʽ�����L��P0����>4u�>d�>�(���*��IY��(��ڶ>E��=t\S�f��?��?�G�_޾S2Ͼ R~�u�92�=z3�����;����#�SH�1
.�pu������Q&�o7�>�_�?�1��Pc>����r���0������(^Ž��v�o��>?i9>�d�����Hd	��m������4̽Ԑ=ٌ=�a�>�@?��?Y�h?0|?��?�5,�h?�2>Y@�>�>�?�z�>9<�>qK{>���>'%>h��=C��:��/=����|"�=A��=��r>+�\=����_><�Y����Ѽg!�<F�<r0�=��=̭=�=G�?�k?��z�
GнX��g�<�I���(�>]]�=�b��MHǽe]���=Dz�>���>��u>U����ؾ���\���<=��6?�eF?�?�.B���O��X��S<��H>��>>v�=E@>���o�ᾰ�ƽ��?�?">o�>1q�?\`�?]6P?G��>os_�ñ�%7������e�>�0�dB?���>G㿾�)8�����,�8>�3Qe�4�J�⮮=�Ț9�{����t>AT�>�1�=�[H��G �eU\>��>j�<P1?�c�>9p?N>"f�=q��<=$��tJ?pћ����J1��d�;5�>�b)>,�R>�/	�� ?m��DBt�W���i�<��ӽ>�z�?Z��?(a?MPW��R潤]W>��:>��>�0�<��#��M��K؁�C�>���=K��oT��b#�:�hw>�>ʼ����Ӿ�f���g�H���B�����BǾ{�Ⱦ�S��H�>��]?=����������|�{��w����A�=gB�ǜ��+��� n����w��?���?��"�iǾv�&�XhѾ-|����>*�齸匾���6�H<�VϾ��־����!0������9+-�w3�>?1K�ᮌ�"�t�SC,�&/���d>��.?��վҶ�W����<8�>b��=��꾝���p��	�.���Q?�V0?�ܾHѾ�9t���=�4?t�>(�>ۥ����"��>(�(?\�/?t%+�O���ֳ��+���Ը?=G�?� ?�����f��\̾N��m ?��?�|�> ��)!�Aq�>+4?�&?�2	>���������$?&D�?|l���5x>�'?dP�>��ݽ0?߾��N�ņ�� ��=�G�>ݠ���H��
��[,�\8k<MH�>��*>��b�˾5��>�꾾�N�a�H�*�3��?ʛ<7�?���(
>{h>��>Y�'�_���
k�����L?�4�?��R? �7?���U+��ª��U�=��>~��>�C�=�N��>���>��hr��q�ǿ?5��?��?�^[?�l�6Gӿ����������=�$�=��>>��޽�ɭ=͘K=t̘��Z=�x�>x��>*o>F;x>r�T>ϛ<>��.>n�����#��ʤ�2ْ��[B�� ���wg��{	��y�����ȴ���U�������NГ�l�G�b�� U>�ˇ���-d�h8?�2?DE�>Fa>N>�=`��j1�S��6��![��)����|�����ܾ:����8��9:�c฾ \?����>���>�q�=�p%?������o��e?Xh:>)D?�I)>
�5=��=QX�=��?��<�L�>�ML>@<>��E>m���Y>m��}<��R<���>1p%?�%��Ѽ=�ut��e�cR��`��8=W?��=�;����k������>R���~��F}���޼��>�z?��<�%��I�<E�x��)
�ݏ����5>�X�;^^�=l���2���=�ǿ>ى5�z&>j�>�@?���?[?�0=��?�0�=gٯ>zR�<s-b>��q>�g0>�$"?�X?��,?e*?��+>�:���z�=��<��*��OV�:��=JG=k�B���[=| ��P�A���K==: ��yA>��ֽ^@�=�#;�G>0��>X5$?���>ȱ>��(=�"#�zY�Pۈ�0Hs>ۙN>[��>���>K$?�b?*̣>�~>�t񽃠t���.�]�>">�C^�����L'�=! >�{�>��:?���>	�>>!��+x�����>1�u>���>*�?�?P�@>>�x����+�ҿ�#���!�=����.�;��;�l
I�5����-�"r��ȧ�<3Y>�K�>��p>-�F>B� >Ÿ2>��>�F>Z�=���=�s;�u;$�K�tP=FX�8�P<�rN��G�]���ᏽ�x��\�R��=@�q��e�^J�>F�?{�=(�]��l������_꽛k?A�?�?���>UX";r;S��Y�Qb7��w>f�2?	��?vR?^%��3X<LL[<��>w�>ب8=����u�c=��=<T�.[����=м�>��>��=-�(�\]F�h �s,�>��>���aK�?�Ŋ?3�;���=Q6�g�[��w��3bf�R8�=�u�<��V�*"ھ!�/�X6&���U�>�g���?�>׮�?;��ȨL�aYľ�����i��p��n�?�� &>��?�>@����+��@7�ʐ��Q��t���,�>�U>�i�>� ?��?���?���>8��>�����?F��=>)?��"?��>,&�>��Z>U�>Q��<�vx=��1�g���=����X�<�=>8�6>*l�>X�G>6� =s�6�D(����>�:���CM<U�=ܻ;q�=��=�c�=]�?�J?�qj��7�0zF����T�>�P�> ՠ=
���C.�������~>�=�>*�?�_�>��e=Sq���?����q�;��??��$?dn>p���EɽꜾ����;��t/�>��=7*�����6Mﾥ�ξ~5>@��>N�o>��>L�o?:�g?�?4?�u�>��Gy��3ψ��T�詽x�8?54?�q�>�vC>n�\���K��_�P���+�<��Q��T�=u��=K�R>,��>1�}>4�>Y�V�F��pK~�����K_�5z->��==�>ǩ�>z!+=�������B�:?��O���𾦨�����⠽�O>���>~�<We?���^��Ң�>�A���Q>�?[��?\�?�8���W���2>�J}>�X>��>6��4z����Gd>�i�=��f�x�������(P>�z>����Ǿ���vwW=}���F(���o������ھlY� S�7��=��9�����|̾R��L-��K���-ԽH!�.%>�<{���+�?I��?e]H���2��P���
۾u�z�!x>�ս�@=%J��
�<� =C�b����`���r�?!�4�$͟>> M������t�q�#��X����K>e]0?cD˾H̾��S�+=��'>��=��ﾈǏ��ߙ�t���T?n�,?����پ����bI>�?:�>:�>�Ч�v��ǌ>�x0?��$?�Y�{D��f����R;ĺ�?���?`�??d�N�BtA����@����?:�?�-�>q���9;�"�� �
?ʧ9?Eۼ>���iG��& �C��>��Z?Z�O�A�`>7��>⸗>��ｫ���<�&�l���o�����7>~|�g���h��2>��F�=ٞ�>m*x>��\����o�>A_��bK�.gH� {�SE��o�<N?�&򾄦>,�d>n�
>��-�C���y�l���ԒM?O��?�RR?՜6?')�F�_O��Fs�=W�>���>���=G`�욙>r��>����Lp�Dh��c?���?���?� V?b8l�d�ڿ1���uʪ��Q����>�>�D>bOн�X<�m�=����u��)�>��>�ԁ>'��>�=�>��[>$j>���H|&�����z���PG��J�)>��l�A���J�Y�/K.�'0��cҾ��=�TJ���ֺ�]@�`�`��H'�m؏����=���>��b>��A>�s>%Q3>��нgX����K�߾��Y@��Ҿ����پ������b��;���eA<�(��:���7�A�?,
�=j=��>I���Dw�=|��>�Il>6��=pM�>�e�=Wd=�eo>� 6>�G&>�.�>�ؐ>Xq�l�9>A4��㈿�i��}>�|�>#E?���r�">A�x��kN�m=�b� ��k?&��=����1���dy��>C�ż8ׇ���vQ >�`�>�5�>Z>B_V����<��ҽL���|->��=��=y3���+��M�����=dF�>JL����>��>�2?�`?{?�.�=��>j�=6�g>2�T>�P>�.�=��`>���>wd?�7D?Y�?� >�]��X^�=�LY>e��<md��x���朼������>��Eo>��=�8�Kݼ=�h>ޖy�����w�D=�+?\F�>(n?�?�>O>�8��y��S&���>k���-R?��F?��?�n?�߼k��=Ƞ"=��<|�ݾ�R�>�N=4"=�*� �4�н�>#��>I�I?Z\�>p�!�<57��:��/5>ޑ�>� 6?|�[?MSf>߬�<�������Pӿs�#���!�"i������Ǒ;��;��eI�U�%:X6-��	��H`�<�U\>O��>G�p>AE>v�>�\2>���>��F>�]�=�Х='��;�;�C��:W=���7�[<��L�/�л�Wü����}����fI�6�8�=���ϼ>=�>o�?��=���=L�������<�>���>t�?�&�>�׃���\��I�-�%����=�> ?:�U?ė�>�U�N��=��v���=H��>��U>_�6�t7:��Α=HE
����<��B>���>���>����A����_������K>�p+>>�~����?5F�?���=ZT�N�f���z���f�q�s���=�w�>������nD������3����*�>���>r�?ٿ��ڏ��\�"�,Fo�LЙ�R�7��M,<��\> S?z·>o�����l�8�W�.����>K�=?Z�;pd�>��J>n%?� Q?��n?���>�'+<E=�Rj?�R���]@?��?��?�9F?ó\>�6&?b�>jp�>�]>�t1�˜@�k<($�=E=͔�>!b�>_�H>��l>ֲG��D.������U�%��̯=�O>I�=�l�=�ծ>uY�>�|?�l�+�Z�^���$��D$>�i�>M�H9�>�A�Q�.�[�o>r'�>{)?p��>��j>�T�����I پ��=��?@?I��>�qA���n=�¾x���~�p����>R�=a޷��0ξ~\ξ�=�`2>�x�>Y�F>J!r>
�i?��??D�$?�\E���C�2�K��)���s��h���>B7�>^ =�Z�o�L�o'��1�Y�<��{5>z�a��E`�;�">:��<�ޘ>�]i>�t�=��J��<����ǽ�=Հ��n>O��>��?���>�Ue���˾�+���;?���5�	��������*���8>vi>�K�:?���_t�è�\�E�ɩ>/,�?���?z;f?��6�=����Z> HU>x�>c��<z0�}�$�%���~)K>H@�=Vq�G��	�����W>O�Y>)ϱ�J~���վ��9���΁�%_m�	������u��U7W�.�]=�׾֍�<x���྿�Ծ�׾8�z�)e9��F�R���_�۾��?yR�?5�����d8��[L�>C�����>1�X��n0�M*־<�Ծ����}~۾
}��=!�l�2�-�-��eJ��P�>ާ�=���	7����n�>��>m}+?e��,`3�u��a��E��=���������|�����?����?��?����R������=�_>Z'>!��>�F�>�KǾ�"�<�>�g?�.?�2����X��~�l=���?+��?�=?$1��?#�����Vܽm�>�{?�	�>����(���P�y
?hQ?'S�>M{-�BN���*<���>9��?Iㅾ�>�V.?:H?P�=�(gR����p�����>�r�������OG�Sc$���ʼ�x>���>ڏ����ƾ���v�Y��8W���,�þX�X=�=��>�i*�������1?5�D>��:�>wM�Aư�J}�>�\?~��?چf?�#?���پ��r�<�>�?t��>����u��ݵ�>m�?�b��$mA��� ��~�>*��?�?�7i?' S�[sѿi���{r¾9�j�}Np=�ʽ��=��:�˒U>�����OB=O�=4��=5��>^�>Bt�>�R>`D�>�KX>� ����$�����g|L�3-����O2���Ҿ�.����	���\{�ǲ<kx�>�I>��*����X�<v�n��]P>�!�>铑>.��>�V@=��|><x� �þ�����ھ��)��J�M��'ܗ��Tu�"A�������>t���ž�2)?Oo��_�<��>׻��q��=��>���<�ٓ>Y�>vk\>���>D�:>�n`>�o�=�>��=C�b>�إ>�>X�{fZ��GB�{%��/�=��>h�p����;59^�|�-��?�=���=
�F?J��<���=���0~�#��>��Z�{������7�=˭v>�@�>�V&>�a��ɠ=F����� ��ا=�u�=}�>�Z��ʽ4U����=m�f>6���9>ER�>�\.?��W?��*?�NL�Ti>���>���>�>�"9>��=Hc=E�$?� 2?�M?94?�>�o�x�b>�>!l���|<�w��}�{��9����H>��@�<)�Y��h���ڈ>Mf�<R�Z=>L���J=���>T�(?�(�>���>�O�w*"�B1J��[��Р=��=ZƄ>p��>��?*p?S(�>�E�<�V�䏾�N����>��@���L��qE�����1�>�ߟ>�s]?�F�>S�?>�P\�����=�D>.Sf>���>:�?�9�>$-�=`x�=�	�ܿMM,�O�w ����
ל��PS�C�=��ͽ�V���Ȼ=�ƼT��>]�=]��>��p>�TN>�ٟ>:��>z�>=M�r�����<ޝ>S@=7�>��Y�&Oýdb>��#=�h�l���K6��6 ׼��.>��0:>|7>P@?�-?g>�L�mI���[ѾG�Y�%G?FK?�)�>��>�ù=�(¾J�b�����"����S?J�W?�1�>�K�"p�<� �<]M>Ŧ�>',�>��˽-�#��<3�ܾ������>B��>k��>��	=L;�J�j�(��6�S>���=�#V����?�ř?q�a��C����P�}Sk������w�=L?U�D�C=?�3�	�eK#����n.�ɒ׽n��>Ժ>�}�?�jX���[>e�M�ե���g���c��a��=#Vz����>�O�>?%��F�e������ �����f� ��F�=&�=�{�>�7?��?�`?��?̊?��.?D��=Kw�>>��>H�?�	?I��>��~>���>�<-=q�6��W���T<&Y��R.�=>u>i"&>|v<9�=y�&=��<��@��-�W�r<?�<'<=I�=��=Z>��?g� ?������g�B:(�Ê��[�>b�>A�>�
�>.���ִN�9�q><�>�))?�W�>�Kf>������=���B�='�?��>[%�>tQ�<��>-�J�����������>���� 8�����������s����>�<�>�_�>��x>>R?u�b?�??U�h>@��\]V�yU����>�[���b>9�)?[������+�'q�SWs�o=Ѿx��=ㅾ�޽�=1>���=^W>�V�</�>X���Nl���輾�&=o�����v>;��>�T?Ǵ�>J�=�7��Q���H?.������+����Ѿ�V)�0�!>=�H>6�˗?M+��<{���TU>����>�?�E�?N�d?l�@�^���v\>]7V>M�>@�l<X+8�Ǯ������7>��=��x��s����:�_U>4�x>�;ʽ}uɾ�<��8��ϵ��C�Ɠ �ߝϾ��0�ZBu�oB~�/Ϛ��#þ7co�	a$���i����z���}qE��M�=k�S�eQ��#�����?:�?�K�>�߾���v�E�0����>�#���G���L�7���D�׋ �x����F���,� F_�*�Y�Y��>_�;�
[���A���۾
��>\�\=4�O?��-�ž���|
��(�=Q�$>0����ʗ��,���-P�FRf?��?�8׾?�þ� =H�0>��>�	�>x�=Xv�,}k�}��>��4?�<?�-�������5v��5Z�L/�?���?��L?�*������n�y�Rh?4��>B��>����r�㾺y���u?a�P?��>R"�o����,����>c�?K����(g>�)?���>e��-�ݾE��;��+��>��2=-�=����=�Kv��Z�O���mޝ>Z{5>���q�����>�辣�N�4mH���̾����<�p?���
>m�i>��>��'�3���/w�����>M?�G�?�vR?{k7?@���f��H���ߎ=��>�[�>��=������>�(�>�K�ңq�9 ��.?1�?#��?��Z?��l�P�Ͽ ������������>��=M~,>�Y �p�>ۿ�=�Κ;��6�4r�=��>�nu>7��>���>.Tn>��g>�*��U6&��Х����V8��������u��T���]��D���Ѿ$�Ӿ��ܽ�����M���6`����=������>s^?� ?{� ?��0>��4>�_ɾ6� �G�	�x g�-�þ�� ��U\��Q��%|�W&o��䧽g��@K�7��[J?�eE=d�5>��?�_׽�Z >F�>`t">�$�>��<>���=7�p>6�>`Ԝ>P�+>q�>*(�=��>Q�U=�d���F_��4����>�ԓ>{??/����q�m�D�R!K�%����xw=ު#?�j�(8��g����O�o��>.�>7ؾR�����=�'�>n>�>T^�=��Q���	>�m����]����=���=e}�=�M+��N���>�<>��>,��
�>��>�;%?j!l?Ċ?��̽J�?UH�>+�R>J�w>ݒ�>�a>@I�>0\�>�a?�A?�?��U>����>�W�=v�̾���*Ki�%�=�3�>}�>9��O�2����>4����E�=���<��->��=�d>���>'�S?��!?�?�t>�J����V�X�?s��UZ?.T?�-?Q�G?GN>*2u>�3ӽpm=�D��]�>V�%>74����½��>�w�>8�.?��?4�,�`\M�.���2P�==��>H�>�v)?S�>���=#gC�2��Q�ￄ�����a��>���=��<-RK�qF�=XI ��B_��@� '����=b��>�U�>/�>$��>u��>8R�>�f5>[{�=g�c=�_�s���P=M}>(���'�=]���V�at�=j��H�<{��<�n��w�I����3<�>j�0?+i��G��X#�� p�UAA�R��>5��>���>\q�>��>�d�#x�&�2�՝>��Q?�gM?>N������*e>U �=MT�>�1�>K$L��������H���0M��>���>�.�>g}�=�Z�������վt0�>t�>�1D�4Y�? �?[>̾u��b�Z�2�|������>�b��!�<��2��f$�a(p�I�N����Q�ռ�?�2>F��?��H���k>�����!���z���Ab�>f>c6���>�.�>� �%3��2/�/6ƾ*g��0Gy�O;+>�>��>�a7?��C?Na?-�>��>QΦ�OW"?M��?�j�>w�	?�K?Ǌ�>���>�4>�w�=c�7�v�����܊=�#|=F5�=\�+>o�g>&�=)�;lq1=u׸�lj��ʽ&=�'���2=�J= D�=$D�=xN?L�?$?��.N������s�);-�H>��>��"=�:Q>ҰP��i �҄�>��>3H?��?��<>z`�����L;����=��?*?�|�>��R�C�i���o�<�Q��b>��>��B>q�9��9����վy����A?A�>�=�=�B>��h?��X?�PG?c�2>@`��&���Z\���=]p%��;�>�R?��ݼ˗��jtU���t���>��1�Y�>a����=�h�<4��Y��>��>>�7M�E< �|Kt>ρ}���F>2�=�@�>�)?��
?!��>U��<[Q�(�M�B?P0]�u����D���ʯ���>�v>������!?4����=]������8�zc�>��?�.�?^�[?몆�\j��e>�^>=Y�<
=�;�@u�3F��}�X�du!>��:=��,�&�R�/R�#P8=�A?>9ᴽ���款	!*����p>�����Xھ9Yɾ��ھ�����<w=���:����ؾ4�x����&/��O	�<|�����]���w��ߺ�D�?(�?ȍҼ�����q�c���u��q��>/�?�
��o���(/�~B���/���^���8��/���E��?<�37�>�Y��^�e�G�'����A>�d>	P?��#�N���on�H�潝�>��=®�������Rx�FVJ?a%#?�E�I��^�<>ϒ޺=ѡ>{�?��<>NHݾ��;�G>	�<?��?`�=���� �����>+��?���?�A?Oq8��B��w�{r.�>N?-�?���>`��Rl��t��F��>�]9?BZ�>������D� �cq�>��U?XtQ�IC>�)�>O��>D4�q����9C��s��"�<��?>����ý�K��)S��D\<덕>C�w>cW$�K莾���>��龯�N���H�������:I�<�?���D�>�ii>��>T�(����������_M?g��?�mS?"L8?-���������=)�>��>e�=���
��>���>�$辒Yr��C�gz?�%�?۴�?�VZ?Vam�К�UO������Ɖ����D>��M>d�,>���FF)>]����J�Ə�$p�]L�>)��>	a�>+.!>��>�Mr>yP���f%�R멿Q뚿�k3�kV�X��fh����1��
K��͜�?za��"ȼ����4�5UA�L��fp�*���\�>΁�>ݴ�>
��>�j>�>��e��������9��i>�Y����{f���w�e)I�7
���i�Jy���M�?���I��>�?&��mN>���>�[��ZK>ێ�>l��=��w>iU�>F6�>�I >��C>ZU�=�>�8N>S����a��Z=����=Jn�>3�;?TZ���=����j�9�{n�՘����S?���<�h=�6Ϋ��%��J��>��<��Ⱦ����=�b`>7?�>��\=���=7P6=Q���R������>��>��|:����[
����<�n�>�~ ��؟>$�?�*M?��?�<�>A%��2?���u��>���>��>�T>Z8>���>�y?tI?5h'?J@>$@���}9=v��>R��>��gq(�y���_��[<8>D)��4�H;�ǀ=?^�� �����=�g=V/>��ʈ<�K�>w#&?���>��>р��g�c�F����G�">���<L��>���> !?Z2?�߿>�0>��}������iȾB��>�ϫ=[�T�>��Y�����>��?�_??��?	T�>\X���Y���p>�=�>E�>��(?%�>w�Q>9��=5��|<�M��F���u=A&�=�`U=��4�+S}=åZ;�iƺ��j�{�I[�>!�>��?Zv�>��>���>��>� 	>i���'�>�AL�IE���Ņ��>�$)�Jz	>&���9F<���>�q0�����ۼ��c=BP���3�?�4=?G�5=dL��)پ7�T��;�?vߦ>c��>7��>�)�=� ��0T�2��u6>��N?��M?̵>WV@�Jt�=�A>��v>���>�`�>gB���,��8e=�4پ�>����>A��>]�>a�㽩,�TxT���ܾW��=�2)>M�p����?T��?;x���Ɩ���0��i��4��S�i�����%>�������i����������R=��>A¤>#֞?����ݠ�ax��d���ԧv�K4��/]�1ü���>���>g���:Y���C������p�S-*<�_�=��>h(�>�(1?M�=?M��?c�?��>;����}/?���<>W?�?|�$?>./?�S�>��>!ɝ>Ӕ	>.=�����.��WK�=��,=>�?>*�>m4->�[�=�7��\<X)���U���Q=Y�ƽ��M=2h�=��=<�<�s>��?`�?5մ�e�������+�����>-ʊ>>�<�8V>�܎��E��]����>G0�>%�>[Đ>���	,����+����1?J�>�r>0��{=��:�`&W���=?��Y=J�ݾ�J���&�����E��>]��>���>���>Fe?�7a?DG?�>t!��@���Tv�c�>޾˾�?k??@E��χ����В�4\�uN8�0��=O$g���]�'[`>��=�O >�	>��=)���Ӯ<(D3=:֑>$�6>d�>	�?�;?r�>y^�=�����о�@?ϋ2��V�ݶ�G6�����ܜ>�@�>�)�d�?
3ּ�[d�n���6�5�Ք>޷?q��?��\?����c߽�b>0�d>9��=�O=����q�s��^&�}m	>\��=��K�Ëb�[-��5�}�J>"���dg��/��8�;���a�_��=�z¾�н�����}���_�<�D��x�=d��ξ��1�[iѾ�f#�������O2ȾM_��W��?ӕ�?�!�=�8����w���	�dը�<$�=�ݾ���c�!��m��ۄp��!�	@�����#�A���X���j����>+��RY���U�4�ˋ>�$>�M?�n��8��J�����D��>ُ�M����6��ns����<�n�M??g%?U׾Q羕��=��=���>�?zT>|��	Y!�.-M>��?g5 ?s*ļV87����'��t�?&�?j�@?�f(�� ��˾��2��x ?ܨ
?��>����+*̾��&��;�>,_S?�O�>�������"Z4���>˹m?�^~���S>	�>h?;	`�Z���������g|Z>s)�=+T�='����}��j�2tv�S٩>!�=>=���&b�5��>���2�5��7�	�辣�ͽ_A=wO?y��2{;>�#Q>b�>�6��Ď����M?{`�?XrP?V�)?����Ͼ�秽��=g��>xz�>x}">׫
�R-�>} �>�ھAzg�����?.��?JX�?Qk? ]]��Z�B������M��h�P>N�/>�f�=	R��KJ>VSb>�&+���Z=*U�>0o�>/>#$M>$ҁ>�C_>�͏���)����t:����!��Z �~/��Ծpq��y3&=:r�Ƕ��su��߽���^S��ݾ|���-��t1����>=�?M��>��>Z��=�|>�+ �(Q��e�z��������+ʾ�
��24�	½K-@���g�B_j����<.?Dμ�,<*?�6��W&�=��^>��&>=>=Z�>�) >rB�=�Ϊ=R�~>1q�>� �>��>��>R�?:>+��a����i���2���L2%?��,�c������n�3���Z�m�>̽?����a��i���!�����>h�=����@��y>�%J>=Ψ>��=>I.>�\y��)��hL�t��<9#�>��$=�&�>���B��<�=��>Ґ�B�=i�_?�/}?�bz?"��?��=4\8?��~>�c�>�e�=H�e>�$�>x�ֽu�A?�?�?=?6����Z��z��W��l�⽏K=�k���=$�g=�=x��=���<,k+=��Ž~H�=��<���=<�=U�h>@�>B�!?�q�>J��>]������<~ ����rf*�]��>r-�>�B�>�ὖ�l>s���S��-�Ծ8K��x��>p��=�
]��!f�����"?d~>]�?��|?�uɾŋ㾬��<�����'�>9�	?�)?�(>a�8�`�ѽ��l(￣}���^���A<"T�z/��g�&��>3�>�jL�Uݙ�9���D��>u�>�9�C��=4Z�>��>Fk�>m��>�N>��|=>�����$�Q�=�hA>b�+����������r}��M�彜Q��_5�=�=�5v���Լ��?>7?E�=m+Ƽ����g���{���`�>"+>B��>Ũ?PJ>4��1�g���2�G�@����>~4?l?b�����=(�:�5\����>�P�>i`�<l-׼2eȽ"r���R�=sI}>.6�>ê;>����F6�`X��qо<�>�m#>~쿽�t�?��M?������<N!���+��J�8ޜ>B�>�4>����@��_���e��_��,5�;u�'>`7�>�z�?����7�=�׵�JA����d�fE����I\���>��>\5��*�7�
���� ��C$ӽ_9>�tb>ͱ�>YE?
�?#�o?�=?5.?ޠK���>g�
�?t�$?��?CG?1=�>�?�=���>>&�>��>�P�4���-��z��]�=X�=���>;=UN�`�{=�0��M��p�N�R�;>ް!>%Ư=��(��,>��>��?�'?����^E��.@�^=����j�sr�>4�=�2���Ǽ�ʔ=�͡=@,#>G0?CÞ>��H�~��ʈ��a���ǳ���MI?��b?K��>|����i��n�����˥?]��>=��=[h�=��,;g������>�� ?ټ>rí>��N?��R?�W?����h˾dG_��w%��{��NP�<gY�>���>V	w�N�D��<�f�=�8�&��оቋ=s����I�=���P=��=���<�c�>{8K�
�0��w�'����1����>�9�>Ǚ�>�dt>��>���?����E?�ϩ�Bh�Qwx�����vF<(�T>9�S>����n� ?`a�	���U��\7�'u�>|)�?��?��c?F)����dE>��6>$�
>�ڠ<\�н.hw<-�R�i�6>�>��~������B�����=� z>Μz�v|�����D�.��B���tA�^����þP�þ?�%�!�߾0���������Ŏ��7�ma�������\��i�2��^Ц�T��?j
�?r8�>�]�=�փ�}x�R7��>��+�|G������=��������"7�@6#��U�I|���b��y�>��*�t���e�&�Bq���D�=�8<?�9����ž�����ڤ7 �=%N�7���-,�����_??"Y+?{���;$�[��[>�?�Z>��h=�����wj�e��>��:?B:?[���������uW�q_�?���?qU@?�;�yN0�
���7��w?��>���>�7�� Ͼ~9i�� ?�?8<�>�
�Wi��v !��>N�^?^[F�<;X>g��>6d�>~������]����C����C>W�:��V�X���E��[�=�L�>��>�)I�2���S�>����4��A4�7�w�fO=�� ?y��:�+>G�>��>�a��
���~����Ž�yK?��?��T?��,?�(�����y0��^�q=U��>���>(Z>����"�{>�?�d��Of����'?
C�?�z�?;n_?��c���῝=���`վ��޾�=�ϩ=�b1>p��0�>�H�=@��NI��t��=Q`�>��5>r�>r��>�D�>�>H��1O/��֨��͔��D��Y�{r龘⃾�	ﾉ#�`�N#���'��hqO��:���\ �ț
��
��Oxh�#V�DJ8=�?�<?���>��=�15>:��p�H�8�
=2w��]ž�����|���$������Z�Sb�s�)��Q�$�*�]H?� >�jw=�1?f�#> ��>��=�UR��b�>�꽱Q@>R�D>'q>��T>Z��= �>2$>�5�=��>~�h�4x���U�"7�xTV�<?H_/��9$��Z�N�������^�FI?�҃��Ds�����[������>p>�=�p��)Ň���.>d�>#bs>c��=zX(>���?��oh��\U> �>�->|r�>�w7���0�a6�G��>ų���6?�?c.?׮�?f�D?z��e��>�j>C�1?ӄ?���>S*?�¼%>��I?�1i?�H+?���<�������n �G
���x>��=2����~;d��Ή:>�;ͽ�����>s�l>���<$�[�ϼ	@?=L��>y?Y�>�+? �V���Z��h�S�/F3�́�>X�>�*�>�?��d>�-8=�li=�Ͳ��;� ���.�>�:J>;M��ϔ�/�L���?�t�>��l?�\;?�����׽���>�Pj���M>~��>��:?�:Y>�zh�n����1��L�+���ٽN��=��>�v
���B=��⼔{�����
1�<�>J.{>��>?��>	�>0�>*;�>V�L>�s(>,I�=֢�;�߽���;7:����a<�QF��&��Ss�;5�[�ꢺ=��=s؆���Խ��h=�P?���>�t�=�u>g�aξp�m�uA(>+�{>� ?o�>���>�����I��j:�@)�E�>�pC?6��>����5�&>��$>�J�>�'.>��=�c4���y��)= ���%>`$?�p�>�ν��8��*����`V�>�>n�f��S�?CI�?��L�&�rg��s�S�	�f�wq�>YO�>oD+=v�=+S����y꥾͍���}>�3>fm�>��?$����>�ý¦��`Ae�_A'�	����>N,����>X��=�꾘SE�mN���3�����M��=��>4R�>�G>�:U>� h?P��>�S�>��o�$?�U���&[>�-�=�J?΄?��u>0�>

.>@��=�bc=�rȽ��^����B:����=���=���=�49=�=>L��������h�r�- �v�=9�5=��=B;�=(�#>���>�?��j�� W��3��x���=��>��>\��8�_����4���>=�>�&�>���Xؾ�W{�s���-�2��P0?P�`?�X�>�)����f=ɷ�������>}�=L�=���]�X�&�ɾk¾:c�>"�?|G�=��h>�j?�N?��9?�[�=��A��c�r���T��/R>t2]>�,}=}>�bt�83�̔k���R��S%���Ɔ"����<�Ҏ=Z�>�V>q7�<��=#�<A�L;"/����<9#�u԰>�R�>��?�)>ʮ�韾-��@�I?�_��ɷ�iȟ��yо�2��/>��>>� �ŗ?�/
��]|��㥿~�=���>�?���?jc?]�A����e�[>��W>�>�k�;n�<�\]�<�m�0>�g�=Vwy�&+��U�V;�\>�Oz>��Ƚ41˾x��[�G�����J�D������پ��̾�������ȹ��Y�8�������OQ��4�뾖���7���z�;���R��������?Rg�?eQ>��Ľ�.y�xx�iKa���>a���!�#H�e���䯾D�Y� �5@A���j��iq���=���>��S��J��/�y��#(��~Ӽ��2>^/0?
 Ǿ�ز�:��C9=�o>+r�<�4�oō�����q���R?�Z7?�Q�k���ؽ?�>��?O�>{�)>�镾��꽎{�>��3?�x(?^��玿�u��%%-����?��?TB??P��w�)��_��lI���?/?��&?��,�O� � ޽���>W��>���>�ڰ�e�m����C�>4�T?�H��Z>���>�<>zT�<V�������ݾ�=�@>b�o����؅y�p��N&>b�>�Q>�4�"�}x�>��'�����(Nپ��ܾ���C���W��>�1�k�>a�>�_C>�d��<|��Q��d+
���\?6��?�M?��>'�H�)8�=b�;�E�=�=?�d�>�>�{r�=�<.?�B��Za�E�
��v�>g��?7d�?Q2�?����C|Կ<��������絾��=%]�=K�?>�ݽ�X�=�BW=/���R�޼>tS�>��p>�x>�uS>��=>�J2>�B��+�#����]���JJB��#�#/�Kd��e��v�v3��Ĵ��;��}����1���Ȕ�%}L�+L��`8����q�,�)@&?�?M�=L�H=9��=�v/=ge�%j����8��]�|E �=�����/��;0J����OM�DU�e�?��j<�5a�ݏ1?i�=�n>
>3Gr<��u>�Q��t�=p=� G�F_
>ç<\��>\M>b���a�>
_]�9cj�o&6����=�V@'?;��=�2���Z�* M�D7�D��=Nļ>���<�|������И�ً*>�mm�J���&��)�[>��4>Vn�>�X>�VT=8��ҥ��p�
=�-�=�M>�,>�T>�/x=�4w;~\¼lT�>b����*>�}�>s�<?t?Q?f�9?r
)��C=��W<��?�?�Tl<^]=?�#��?��E?�:?Ȏ�>�c������!��b=B���	����l��Ѧ����9<9�=٥�ɢ=[+>�g�=�dJ�=M�=�\��Jr��'�{>�ӻ>�?휚>/��>�2�O,��E�p�[n�=�2�>t0R�Q�=�?���>1h�>k`��If�L��n������>y�n>�KD��s��&�#�;|�>wR>���>�RT?�i�d�後Z�=�[E���>�4�>�3I?���<�o�=�̮�%|�y[ڿJ>��Q'������$���^�<�[ܽϤb:�6�����½��<��D>~oR>-Y>3SG>ebT>\�b>� ?"+V>�Ь=��>�=��c��N��G�=�ϝ�\[g�Cd/�;�̼�㟽�s��aN��'z��'�D���W�ŕT��P?3�	?φ=����qK������f����>�h�>"3�>�>��U>��(�j_V�0��Tƽ�v�>!m<?��> ">����=٬���%%���+>���>�9>���=����J��m<�=��>���>� �>Ǌ���L�c�3���k�>
�H=d�ѾQ��?w�?��8���=��׾��U�\_?��D><L>��.��n�>����a����Y5��٨�=%�C>��>�1�?ƅ�+=��ɡ� ��(��I	�5�G>�a8>���>GCi=*�����i���0��X��1�*��F8>���>1%�>S�>�*R?L�!?G�2?~�����>�b8>�Y?�o!?u]?�k?��>:@�>�?s<�>�\Ի�X���������	�Q.=�u�;�&�>A���r;>05E>ى�;�޼�m��̼t뵼ڪ�=�Q=�z,>�ʑ>��>�)?&�㽢��� I�� ���m=t>.o�>L�&=������A�ȼn7�>˕&?��X>��ý7����6������qX�@|�>��?۸\>��h��Q>�C��־��H>��>((�=4�½N���!n�)������>�~>�*��k��=��f?h?�*�>�֒�|+6�7|��g�)��Վ>�L[=ʹ��E�8�Ã$>��x�2��⧃���~�"7�^5C��'�	���'�=��]=0�>���=�^=�^�V��=MJ���a��(я��h>���>��>�8�=�C$� bP�0�����I?�S���!�;F��L}ξ���>��@>��-?���VTz�<|���?=�0u�>|��?�z�?+�b?n�?�Ƨ�ކX>�!S>�>Y�m<S�8�c��(Ń���3>,�=�ey��x����<�]>��q>Ž%�Ⱦ�x���>�ɇ�����W��=X��o���8����'�'	���� ��X�,w��w�!�������	�#Ǿ�������=z$�?ߤ�?�=�> �
=�#i�q_�Y�?��l
��'g�:ܽ
����Ѿ;���z�����7�6��gr���������>�V������{�ޜ(������R:>~u/?�ƾD�������\=��#>��<H ��kk��8���U?�8?������$nؽ�b>X?�l�>�h$>YY��o�>��>�K3?p�,?��޼V����(���y��k�?���?�??~C�-�=�ҍ�����?��?�K�>cr���)ʾT��/�?�1?L��>���B���\����>O�W?� O��"c> ��>��>N㽔C��b<�2M���D��}�3>t9���R��<c��<���=���>] x>L�\�-����P�>��ʾ��e�Kמ�}�I=f�w>���>[ݲ�U�'�f>���=ǡ5�e��֐��1�m�d?j`�?��_?*I?�������3���c>)t�>�?HRO>Z��M��>��>K7��Z���N����>�z�?�h�?�{{?� �(�Ὺ婿�t����W3�=�Q>�Y�>>���<&=�>�q>��<�å>�=�>`^>�y�>H�o>jҍ>U��(�)�W���e䙿���cܾXӾi`������6��#M��<���e����<X�=�b��r|�/�½{9����B�0>�?��>�0�>"�>��=���w���:�Q��]�i鷾D���@	�A����=pO��IO��W�7���8���0?`��-F�>lh-?%y?=hr�>�+�>�݃>�=�>�>��=x6�=�*>3��=���>B�>X�>�* >&�?�-�ӿ]�tBi���N�޲���<?^�о�]��Bk��6���žT���䕣>�l��cG�i���UC���b�>�wf=�a���I�h>?h>�k�>ܲ�=��=u�(�s(��}(��v�=^��=��@>rRg>��9���\<�u=���>�y#�7%>=�k>�g? �?���? >_>g�<?M��>�n>���>������:>��)�@?i5�?��|?� �?�8=�DK��D�tA���T�l�3�7���n=j}�BN�=%FC>.�=��=mB(>�Ռ>a�>��<�J�=�	P����>�.?��>��?����M��SK����=�%��>�At>h��=ċ�>0�>�Y
?�����=@�h����G�>�A�>�F��g��X����>Q}�>�F�>��?\
^�ȫ���2*��}6=LL�>]PV>l�!?7��>�r߽���M��C��|2b�e�k�WW����=k�P=��J���=�/�=���=�D�#�S>i��>{�>���>���>�ӑ>�~�>T~>�E>�[=2�>�y��ڴ�������2=B#�����q��W�:��&��!�� �=�U_��_t��}\���?�?�)ͼ��R�}Y8�>�込n����>AH�>���>��>-�=��)�K��6=�n�$��s�>�a?0!�>��>�(�r=��<��>=�t�>Mܠ>�6>�"��[-!��4S��$��'�>�K$?r�>�@���G���b�u}����>"��=��P� O�?W�@?�[���zK�A�.�g���:2�� �>	㽪��=�$\<'��0/�įɾzo�X�ɽ��T=
�>"�?��8��Q�>y���������O�+�;s&�S��ڙ�>�`P>��T�]z��Aࡾ 0�D�����Qn��u�>�,�>��>�F?d?7��>���>�x��8�>J7�=�d?�G?|(?�D]?�p>���=qۖ>���= �=\վ���/��ǽ��Q���=��;>y��>���=N
^=$C滹m��lL�῿�{`�:�G�� �i:R��<%�>�|>>
�>�3?7�	<�㨽7eý���f6�e[�>�I:U�T�{����ľ���N�,>�$?�J>>پ)ˡ��$�K����3�m�?r�G?�|�>~��=���=��ƾ|�h��4>Q�T>>)|>��ֽߕ�3	����T�|>��>N��>Lul>jjb?"�@?B�>?2K����4��j�:~�d�m��%�<�m�>��>��=���MW�Co��yV�=]%����O뽈�=��=[U>^9�=��Ͻ���=��l=�>�����}��=�o�;\N�>��>���>�>���=z��x� �ԠH?䌣����S����ž;a��]5>��@>4~ٽ& ?.����y�����p<�iI�>X�?!��?��e?ru&����fbX>�]H>7�>��<��<�!u-��de��;@>>,�=�`��&����wJ��d>�;>�_�E�ʾ�]۾�L6����g��Ծx�?�g6��Ѿ���o��=�w1=�>�l��&X��"�u�;\��F�k\������������C��-�?j'�?03�>Eb3�ht��M�L�l(�>�ľ�ΐ�@>���==B,����
��a���c� �|�h���Ҿ�.�>��Y��7���}�w)�Q=���n>>�H/?�ž)��Y|�	^e=%d%>�E�<!�<���g��� �
�n'W?��9?~��#���LGὼ�>yt?��>�=&>=���;�� �>t<4?�X-?TT����]Q��?���C=�?���?�G??��K��~?�7����6�?q�?���>�Ї���;OI�h
?N$6?w��>i��n߃��k��z�>��Z?��L���\>���>U��>roའ����>�����g�߻�96>B��k,���n��@�-6�=^.�>&�y>�Y�"�����>Dp�w�N���H������*C�<p�?���]>�Gi>�R>��(�����ω�M����L?J��?��S?:f8?�W�����P�����=��>Ǭ>��=����>`��>�h辞kr�b��?xE�?���?�ZZ?{�m��޿����<̾�ɾ{��=���=�r�>�	�խ�=��F=[t�<[=�� >���>�:>��>���>��R>��>2'��q�*�\w��w|��_H��f���
��0������9�����J������W}��m뽇��u���:kd��l~�]l��2��:�->*��>�i�>)�=8�^���K=�,)Ҿ�l����$˾���������ܽ�4Z����Lu���CO��M��,?��N>d�'?�/�� �׽
;>�F�>Ǯ�>U�>�y�>W��=N=S�[>�h>MƯ>9x�>��l�w��>n�d��3J�@�1�% �\��1;\?�����������3��/��{�~)?�ľ�8A��~o�����3)�>>E��L<h���B>���>��P>9_�>`�S> .���Ia�u�@�2"Q=��<:�>.4T>([,>�D�xl�W��1=�>DN���>J��=%	?�a?�:?E��Ju?'��>i�>�i�>O�?��>�*��|�+?Ehi?�G?�*?)D�=&�-���;'O�t����y%�CX�0	T=�L5��[2>B�=B��r,w>R�=�;�;���=Y��<>�������>D��>yԜ>�g�>��!�������/�x�&����=�>��>�� ?�?f{%?e=�S�g��@���Q�>�+�>��v��Bb�R�q��Kj>��L>�v9?�V\?ؿǾlz6�@�����ݾP�?��>��>A�>�gr>�l �����iӿ
$�(�!��肽cj��;��<�2�M�g)q�,�-�����Vn�<��\>S�>n}p>��D><�>I03>fO�>CG>ڄ=!�=��;ː;;F���M=���G<��P��ۮ�73Ƽ���������I���>��3�T�ټt�?�?��p����p%�d4뾬js�ݵ>��>z �>9N�> 
�=b0����X���8�i@V�TF�>�xj?B?�u?�Z�%=r�	��5�=ta�>�k>�I�=QԼ~�>�%2p�g�<= ?Ē?|pi>����cE��_Y������>��>��ؾ�ԯ?+�n?��ʾ��=:	�@�:�p��n�>3R����&d�=����-.�"Û<��\�Q��?>4��>饴?���ݐ�=&��> ��}$p��� �8H9>�<�M�>���>�2��ʳ�A�c�Ƙ
�滾Po��i�(>��>؎�>�w�>>� ?��D?��??m��|�G?1�T=c��>,�>8�>,�?%�>g>�>&n?���=��><K��|�7�B�=7��I`m=���=�b�>�tx�?�6�WA���m�$z���g(<�O=�"��Kj���=4>ڞk=�%?�1?��:��Y���=��6>Jvw=j�<qw��Wi�	����L�D-�>��>6�5>�j�8�j�w�㾙g��M��a�!?p'?�
?�Tͽ��>���A���Z>s�<=�q�=F&=�@�� �%̸=;�Z>ƕ�=�>�x`>B{??�>?��!?�꽜�,��r��-)�����2w�Wy�>�ˤ>YV�=�ݾc%3�3�o���]���/��;��TB����<�^�=��>9U7>Ԉ�=��>��=m�����t�<��W�	ٲ>me�>�~?+[>gT�=�ꩾEc��I?����H��ˠ�)Nо���`�>��<>G���?����}�^����0=��[�>��?���?�)d?��C�Q���\><�V>�/>�E.<9�>���D���
�3>5�=��y�����Н;M�\>��x>�9ɽ:�ʾ�P�d�I���Ͽ�t=���>�&ξ��&��O��-F�=���<@��3��g�m��;׾LyӾT�p�ЧǾ8Ud�.��-x!��Ν?�J�?��>�I����p���H�n?�{(�>����qZ���r�ӾU��������N��p�)sV��g'��N.�l�>��L�ې�;�q��3%��md��n>�/6?1CϾ)���߄��#=��>槍��lپe����U��a1�ҞK?��4?�_��x�r���m>@M?�e�>b�>�Ҕ�� ���>o35?��,?�HZ�� ��2A��#�#��i�?��?B?Vx���W<�I�i&���>�l?d}�>���<��t�̽���>�?^�>�о��v�� ����>�7?G�>�[�K>���>��`>�'��.�*����R���%Y=$��=.P���$��+�Kd�%l��>��>�Rd�4���.�>+���C� �9��̓���i+=\:�>!�Ͼs$>�xH>�	)>�a,���������/�<u6?�б?�O_?�0?>����̾1"���3=���>���>��A=�sǽغ�>�,�>�v꾂q�f���?	��?�]�?7�V?	�m��1���p��yo��ٖ���˼�hN>XF*��4�t�G�Ȕ�1À��>O[>;�G>��(>]F�=�(_>�I8>�����w+�WȤ�[��&fo��A3������Ǿ��&��.Y��=5�����h���-���s���/��),�,�D��u[���ƽ�T��n�>ٙ�>�ߝ>%i�>�t��6������9�>D�U����iؾ�d���M���]n����/c����g���C�������)?;t�q�=���>����P��>&I=쨟>!�=E�<>J��=E���p>P�=N#9>]�>�7�=H4>B�=�fe�����}����վ����ko=\5&�D��=���JE�<e�2N�>�3�MDG��W���Z��L㊿U�>6\b�- z���޽��=���>\?K>��P;b-4��� >���1&����,>��a.>��r��5�i�ɽ�Ƭ=���>�`>���{<UJ�>��T?��W?�;�>V�)>8ݣ>Md{��{-?��L��M�>��T���<(*�>0�D?��O?u.�>8�?��jW��R#=�L>��=�P�<$�D�4&���]�>N�޽Q����T|�ՠ����<���������NE���>�W�<M{�>�I�?=84?`ܙ>L��������V��g�>r?���=�s&>��?��>6�]? ��?��>d���Yni�By�����>n�>����p��:�a���>�?���>.�>��T��j�9��=�5�>�Z%?5-?,!�>��߽�2M��!� +��u.)��l.���,�����QF��՟�����#Wپ����ѽ��=:FX>�j4>o�>�P�>�5>+��>��>ໜ>n=��j>(�D=��=E���'��=~�	����I$�yt`�1'}����:�*;f�=8j�<C�=&�<+�?�>?�염+M�;��΋ھ�R7�+��>r�>E�>ɕ�>N>�P��^-�����O���a�>#RU?E��>��_�N��=*ݶ=�ق<7��>��>�9�<�D=!Rq���;���KP�>� �>K0�>"���}H�eW�X��W>���=Oď��1�?`?��־W�=х�5kI����8Xļ��.���R>���H��G��0X��]E�O�B=��>	��>��?&;�| �<(7��G�����������Bj�U%�>�0�>�%<>��F�ea�a7i�{��LEF���)>D�s>�	�>�>?��:?2�9?:�s>�HB�S�>6�1=$�,?`?�=7F?��T>� �>W�->}�?���>�Z0>O���Ik�Pz��b�u=zg���NJ=\�=�g�=t<�=��1�ep�;kYY�P�=#��<}�=�F��kJ</D�=�}>��>�W?����X< )�=�l�WjF>K�P>h_)>�>���=��>W=�=�R�>F��>�B?eiE>�0�=����MnоU#<��>�?��>=�>�=>?;�����������>�sw>D��� f��3�_��� �>l��=�R>�gZ>=�Q?��r?Y?3Z����پx��V1��>���� �>�*?����D�:�����F�r�G���w>����w$�-C�>M�Z���>_��=�a{=�v�>B{��騾f:�$�a���m>��"?��I?�z�>��>�WJ�o]��GP?d~L��!��ը�ҟ���,����>��>P>����?���(�x�{����$��l�>^<�?�?�\?��>��O�$0C>%�z=��=`nt>	u��v�.]���^G�Q��OD�	R�����;>�x�=>^D���\�6�Ӿ��'��[ǿC`�AR��@߾ ������/�4�ᾦ�?������:��_��@x����/3����Ѿ�������?�?�{�?O$=/ �E����z�@������o���
>n�Pֽ	���f�<�����yӾ}�'��GN�bW?�91?����mE�?.O�9�ɾcp�=ZS? w�>(��M>A�4����=:�(��k񼯍5��M[���ɼ�!�?v�?�6��ͼ�����=�~=�'?�a?�����(ԽAТ�l�=��-?<�?>U;�Ӡ�ǃ�����9�? �?&nF?*3K���!�����,�8=�(?��?���=��V�g8߽��澗,�>y��>6��� �멏��8�B�>h�6?����*>��?��?A᷾��������)%�><y�����=şͽ�U6�'lN�	$F�Cĝ>�<r�Y2>��F�"J�>5��G��A��B��M��/:$�?'����(�=�C^>a�>D!'�9Ό�aቿJ����M?T�?��Q?��7?��ܠ�tlĽs�[=6��>hb�>�Y�=Ga�\�>`�>�_⾰to�����?���?��?�xV?�j�hB�B��vо�Ӿ��^�JA0=Z��=�WC�k,2>ݥ4�hs�4?@���>!�>��\>�%=>Eli>���>�,>&l��J�$��z�������m��T��-����Ǿ�%�eTQ� �,;��>��H�½l|?�{9�cR�0�d������S�9ik�r�Y?9:5?�.?59�=�v���+��c�d����Aj��d��F�bT�%������#�ٻ���3z�������8�}�>o����>��>#$>��>�`Q>��,�@\E�6!�=�/>��	>�Q>������>��>���7�>��'>��g��g��]:N��e�=%>�!?`���]�'ƾ��p�'M,��7?��=��=��������M�[�?�(�����9N�>��?G@�>_�����>&��>N>z����=���=���>�5�>��N��5�Ϧ|>�>"򾍛#>�.?��P?�m�?�u/?��>n&0?j垾�WW?Lf	>1�	?
>�y4?��V?�j?�׈?GH�><#���4b�=K��\C�1��l_��b��<<�	=;�8�,���%���q>XQC��f���I�E��i��淇>���=��>P�L?[�?l'�>}��?�r�[���?��0��>�p<=�->��>�D"?���>j9�>@:q=G�=n�(���� �)?��3> b���ϗ�v�p�O�>Wֹ>�JP?�a�>;�5>���*=��>u*>?t]	?�	�>HH�=w�<x����gL��LB�$��ծ�y%\��A����G��p���a���l�顙<`f �33>�b�>�L>5��>�W>���>��2>���=h�>1B>����	�����=M�\�i8����=,��>�W�9��X�c�qڇ=�)��`p��;{��?�?�(��A��@�c���Ǿ#/�o�>���>�?H�>.�=>`��G�>�hu��@!�>!P?%�?�IS�{A>FA�=�+�=�<�>-�>�0�=���`x'�|?�������>�D?�_+>�ށ�TT��n�=~p���>��<��:�7h�?D�Q?=�J����M:�"I;�̣.�zh��YX��_������\��J���n��J����j���w>W��>���?��d����v8�&ۑ�x���LMݾ�
 =��>a��>���>��w� ?W�}�����&����P,=}=>E٫>�3 ?*�?��?<?Ģ�>Z���0?��>so?�j�>�p<?A�>�?�.?s�?�T�>[[����-�����=J��=��G>��W>����=�����n6��>ٓ޼RՓ=m ׽�%��}:�}�i>�a�=#u#>�V�>��?)|h�y=<e`<A����"N�->�=`�>�/A>U��=��1(f=�'?$f�>#Ҫ>2t>js������(>w�?�OL?C �>��G�l�U�kQ����=�7,���>*竾�}�<�L���m��Y��?=��*>9�>�O!>޳f?�X<?�R?=,�g�1���_��Q9��7&�X�=�}j=��=h���@k�xr[�����A�t��,�7�>�`��a���>�pT>t�=:
)�W�=�b�=P��t���M=�~=�m�>2�
?�?M��>dr�>|Aľ,�%�dJ?uğ����K$���\Ⱦ.��jk>p�:>�a��?6w��.{��ե���9���>���?���?��`?�gF������a>��Z>�(>�1�;��A��c5���u��I:>J/�=��~��闾P��;��]>�yw>�oͽ�Tɾ��߾=t���Ŀ�7��.;���(�����-���1+�֢ �AT��Ľ�v>��Ɛ<!��Z�C��U$�฼�����۾�ʾu�?D"�?2q����ھ�0O��ϩ�];N��&�=
�t���>�F	�NB=�Y�WQ���&̾QҾ�K6�;Ka���:����>�˾�v��bv��.+����>_�J>Uk�>�žϙ�=�wپ���=�4$�ǽ��!���틿�������Ï�?���>��zⒾ�#&�]���[��>P�>-��>�p��������<�,?�w�>Z�1��j��������M�[��?
ɤ?�6:?�,<�J��"�
�.=k�\>��?a��>ҷ��!��AS���;9>���=fE��̅� ;���D��>��?���w��>�?	�I>U~:;��
�8�ƾ�fd�r�0��-��3@�c>��H�w�i �3ң��!�;��2>�,?���Ǿ.�>+���C� �9��̓���i+=\:�>!�Ͼs$>�xH>�	)>�a,���������/�<u6?�б?�O_?�0?>����̾1"���3=���>���>��A=�sǽغ�>�,�>�v꾂q�f���?	��?�]�?7�V?	�m��1���p��yo��ٖ���˼�hN>XF*��4�t�G�Ȕ�1À��>O[>;�G>��(>]F�=�(_>�I8>�����w+�WȤ�[��&fo��A3������Ǿ��&��.Y��=5�����h���-���s���/��),�,�D��u[���ƽ�T��n�>ٙ�>�ߝ>%i�>�t��6������9�>D�U����iؾ�d���M���]n����/c����g���C�������)?;t�q�=���>����P��>&I=쨟>!�=E�<>J��=E���p>P�=N#9>]�>�7�=H4>B�=�fe�����}����վ����ko=\5&�D��=���JE�<e�2N�>�3�MDG��W���Z��L㊿U�>6\b�- z���޽��=���>\?K>��P;b-4��� >���1&����,>��a.>��r��5�i�ɽ�Ƭ=���>�`>���{<UJ�>��T?��W?�;�>V�)>8ݣ>Md{��{-?��L��M�>��T���<(*�>0�D?��O?u.�>8�?��jW��R#=�L>��=�P�<$�D�4&���]�>N�޽Q����T|�ՠ����<���������NE���>�W�<M{�>�I�?=84?`ܙ>L��������V��g�>r?���=�s&>��?��>6�]? ��?��>d���Yni�By�����>n�>����p��:�a���>�?���>.�>��T��j�9��=�5�>�Z%?5-?,!�>��߽�2M��!� +��u.)��l.���,�����QF��՟�����#Wپ����ѽ��=:FX>�j4>o�>�P�>�5>+��>��>ໜ>n=��j>(�D=��=E���'��=~�	����I$�yt`�1'}����:�*;f�=8j�<C�=&�<+�?�>?�염+M�;��΋ھ�R7�+��>r�>E�>ɕ�>N>�P��^-�����O���a�>#RU?E��>��_�N��=*ݶ=�ق<7��>��>�9�<�D=!Rq���;���KP�>� �>K0�>"���}H�eW�X��W>���=Oď��1�?`?��־W�=х�5kI����8Xļ��.���R>���H��G��0X��]E�O�B=��>	��>��?&;�| �<(7��G�����������Bj�U%�>�0�>�%<>��F�ea�a7i�{��LEF���)>D�s>�	�>�>?��:?2�9?:�s>�HB�S�>6�1=$�,?`?�=7F?��T>� �>W�->}�?���>�Z0>O���Ik�Pz��b�u=zg���NJ=\�=�g�=t<�=��1�ep�;kYY�P�=#��<}�=�F��kJ</D�=�}>��>�W?����X< )�=�l�WjF>K�P>h_)>�>���=��>W=�=�R�>F��>�B?eiE>�0�=����MnоU#<��>�?��>=�>�=>?;�����������>�sw>D��� f��3�_��� �>l��=�R>�gZ>=�Q?��r?Y?3Z����پx��V1��>���� �>�*?����D�:�����F�r�G���w>����w$�-C�>M�Z���>_��=�a{=�v�>B{��騾f:�$�a���m>��"?��I?�z�>��>�WJ�o]��GP?d~L��!��ը�ҟ���,����>��>P>����?���(�x�{����$��l�>^<�?�?�\?��>��O�$0C>%�z=��=`nt>	u��v�.]���^G�Q��OD�	R�����;>�x�=>^D���\�6�Ӿ��'��[ǿC`�AR��@߾ ������/�4�ᾦ�?������:��_��@x����/3����Ѿ�������?�?�{�?O$=/ �E����z�@������o���
>n�Pֽ	���f�<�����yӾ}�'��GN�bW?�91?����mE�?.O�9�ɾcp�=ZS? w�>(��M>A�4����=:�(��k񼯍5��M[���ɼ�!�?v�?�6��ͼ�����=�~=�'?�a?�����(ԽAТ�l�=��-?<�?>U;�Ӡ�ǃ�����9�? �?&nF?*3K���!�����,�8=�(?��?���=��V�g8߽��澗,�>y��>6��� �멏��8�B�>h�6?����*>��?��?A᷾��������)%�><y�����=şͽ�U6�'lN�	$F�Cĝ>�<r�Y2>��F���>å辽O�]H�L,����Mq<�?���w�>S�g>́>/)�.ь��ǉ��F�	L?˰?mS?;�7?k��;����(�=i�>�7�>Z,�=|�����>�k�>J徫�q���
�?��?�f�?��Z?��m��9鿃���?�ǾEƾ<�ҽ/&�=��)>˸_����<�ua'�q"��h~�<h�F>��R>.R^=xZ>��b>��=y���@%���\��ys�N����Ԙ��SG5�����L���m�&O��P�/�{���t���j��8�8��`�=�S��O����e)?��>�2�>Ac�=`�>H���`����ym���8��M������D޾ۢ�:�d��	�y@����B-?%�"= ��>w��>��>Ə<b	�>DU�B����)w<����=-]=C8>
 �=·	>J]�=9d >�`�>u)=�e���]��&�ξ���lM>��:>,�;�� ?��x��߽7M�����6�.>A��>� ��ǔ��a�d����>�bY��5��)�����=��>�?�����Fl>`�==�-9l��u>���9��=�3�>Ư�
L彯��?�E>���uX���!?�	[?2O�?].M?B)�>��7?H�-���?�&>g�?��A>�K<?�x?:4�?㽓?�d?ۭ"�{�1���X��6�i�K��N����<�,�]ǽd~��c Žn>��;6�ܽYw���=��&=5�=���>�D[?Aj?��>���r��c���<�Ȅ>�a0>	P�>��R?���>�H?���>B�O<d1��=����ER�>��>�p��Bv�5,���->�Tx>2Ud?P�?��<ȱ���D��6��=�$?&�A?�	?��=�X�1'R��?�~t��%��W:����MK<�2���71��0�h�*����dž0�
>FX�>v��=���=���>�٭>��h>-�>�'>�N�=)^��m67�v�$I;|7�=u1�=]��<P�=�}@>=��=��="-���3(>��=�Z\��=�<ca/?�])?2)��+��'Y�IŹ�BN���n
?��=�	,?�1?����оU��\A�$�����>|�/?[Q?%���"O�"o���i�9�?�߆>���D>m�ݾvߢ�Z��z/c>���=:�Q>��o�g�w��/+�|Z�zh�>؜�<����?hG?�!���n�"f(��H�iP>�j�(�9
���Ҿ��=��Z��57��׾G9��́>���>�ɑ?�H���$���0�����틿e�y^2���><%?/t?lc>\2~������柾X���\�=���>��>��!?O�?�?�	�>1�>4;c>���=b�?:�Լ�!?C>�L?��>�?�;�>p��>װ4>IWI�<� �����骼E��=�e3=gvD>�<>]�۽lVr���[��.�<;]��)x˽8b�����^�r��߼���=qn>=Ŗ�>W� ?��Z�I^=;hA��׼l]>��=�yD>p�O��;���N��>���>���>,��>�c=��������x  �yw��?V�@?In�>)��>�EC=����ռ��~���>�|�=2U�ǧ����f �����>)?s͢>Y�k>�x?��E?�?�>����3�mx��y�D��$�%�>�7�>B.=?�־�;���l�d�R������G<I/��a�<C��=06,>�c>;��=r�=x�C=��Y�XlH�f	=��<#��>�0�>�?��M>��=��M���AI?�{�����+Ȝ���ξ[b��� >��<>R����Q?0j�{P|�����<�+o�>i�?:'�?A�c?S�@��	�]�Y>9Y>��>�@�<,�;����������1>��=։r��U���6�;�IY>�f>�h���pȾ����29��g��q5S��N%��,��W�I{���q��<Sվ�VW�u�!��y��ƾdꕽ��¾,�`���Ծ�E�x���ף?>��?�JT=�)Ѿ�ľ��`�W{ݾĳ�>
量�v/=���h~=z��c���M�����\�v�@�����V�c >>���И��V�{��o.���2�=�T?Fÿ��Z���"�L��={�=&Ͻ�qܾ�`������GO�z"&?1p?hd��ž��=�\>��S?j	>�q]>O�� r.���O>�Y?�?d���j��#4`���?��?tX?X��<p�O�{J���M�>�L?�	��о>b��P�(�t�p>}�>��>w��=�2��焿v-+��][>�?�>��>kq�>/ՙ>�S��	B��id�=���:8>nG=s*���R;�B���>F�=�D�>�av>���w�̓�>�_�IM��H���������<=�?����ni�=��l>�i>+H#��������Y���K?���?�T?��3?s�ﾕF���~�=�+�>~߫>6$�=��l�>�c�>�
ྍ�d���
�Z?(�?��?�AP?sj��6ֿ�����������J��=D��=�1>�������=O��<��ݻ����f�=v��>T�w>��>�:b>I@>	�%>D��L�(�_;�����,L�mn����Iۄ��������r���#���#ž�|��dK��<5���8�!t��/6��2��Q8�<
�(?[c�>��>��=��Ͻ�R��9��Z�r�n�ܾ��Ҿ������!#���^��ez_�0ԅ��������b��[�>����Ɓ>�'�>�=��^a^>��>�<ٽ'��=��->1�!>��[>\h.>)�~>�2>N�=���<Q�z>i�ᾥ�y������i��;��	N�4�?�\����u>��۾g�	�$��x�E>��>�b����+�緎�F�%G�>���������a�R>�hD>j� =Z�=ߎ =bG�͆m�k�>Poy>K��>�n:>�A�=!���X��h>��q;?>�u�>�zI?�%�?H�8?�"=��>5F�=`i?� �Ah�>��?W�?�/A?�m>?�`$?�+�>���C���4ӽK��R
p�a6�<��<�X =
B"=�E �a��+�G=�[�=Jp�=�,>
�c=��H�B���FU�<�>.�~?CD?��?�e6�ٜF��q�͐�����>z�4>W�(?�rH?�?BX�>�b�>e.�>~P>�R���	�g��>�>p��P�a��!�=��=8�k>�cF?��?9&Ͼ�a���>=�'�=L�>^R�>A�?�kM>��D_�<z��]�⿩��R�*��H�]�k�f%�=��{����V,�x\��e������P>�[>
N�>zn�>5�N>?�X>U��>c�M>�?>>�~=Ѡ�=�*����=>z�= �$�c.=Y�Ͻ�k7=��ڻ8#e�V�Ⱦum1����+���R= �>4i	?��W��U]>��������ܽ=�p>�	�>�O�>ܔ>[�U��¾|vT���H��﻾GU�>�C}?T~"?�{ȽD9L�<�.�9�u�_Y�>E�q>Yw�=�VR=�d���q%�|���$=�=���=�-e�DC����������d�>^<�Oꩼ��?-,h?ɾ���P�&�QJA�������>�0�;��J>C5���[���־K�����l��� �����K��>�(�?@��E[�>�C�bަ�-�t�/v�����>���>eSJ?��>߄��i13�������N��jN<�q�>*�����>\�7?C*?�n�?J�@?�0V>񌆾��L?㹿�i?Vu�>y�??=R?�8V?(4*?\?�=�-����"��Ͼq�����8�3�X.�>&�>�ϫ=x��e�Z<g�=ȳ_=�8[�!LP���=+L <ɻ">�=�iP>3��>X��>��>E2�>S��!)��'8;>Oi�^�?�zX>�£�.#x=�#?>�?5�[?r�:?�`�>o�����]�t�;��	�>U}??�?V?Ls�>��(<Ϟh��V�|� �U�+>o6u>>��8�χ۾���!�'��=��
?q>6E`>��|?L)B?l "?���J�.�a�t���+�����;��Il�>f��>���=�޾� 7��~s��]��j,�z�2���E�Z��<���=�a>[L>���=\g>�q= p ��vI<�'���>Z�>��?\GZ>Ɋo=8䫾w��$�J?a0��v=������˾i���>�4>՞D>�*��?m~��\x��板Ic7�B�>#�?�x�?�(h?q�>�y���g>��u>�6>����^�����:?X>z��=<�}����<u� >s	�>>᳽Ǵž(w�$i�T�Ϳ=:T�g}���#��yѾr�Ծ�~�����k�ܾ;f	��/��<���W�����Nܾ��Ⱦ .���޾
6ǽ�a�?M��?E׆=$�d����#�ס��"�NM����=pA���I��8�1 ���龵^]�#"w��(F�P�־?�=S�c�*6r���V�۱�Go�-	�<H*?����������S>���Aɾ�D�;���`��h���y�m?��E?{iƾ�
�VS����>��?���>,�?�����V����=��&?Q?s��>V�8�U�t������g�?���?w_?7F�MR�����>Ժ�>r�9?��v?�9AǾ�6>��->o��>5��>���KeU�1�����#?���?̲:��C�����>#ɏ>"�F�lS"�+g>ؾ5ю��?��i<���E5H�]�;<�u�>J�?�h?Ij�����>	A�� N���G������R?�<��?���>��i>}�>	)��Ќ�"ĉ��}�ÐL?}h�?�S?��7?�(��779���a�=d��>,�>�=�G	�ڨ�>t�>���?�q�o����?q�?���?�Y?v"m�BGӿ��!��������=%�=��>>��޽�ɭ=��K=Kʘ�
[=�\�>���>o>8;x>��T>ޛ<>��.>o�����#��ʤ�4ْ�\B�� ���wg��{	��y�����ȴ���g���Ȣ��vГ���G�m���T>��0����:?0	?���=�Fe���>��㾈��Ҷ���׼�,�a�;�C��Q�8��������(l;��<�S��/�F��z�>���>
����?�3=�}>=���>�W>m��=2>�>�im>ҰD>���>���>6�>���>�@�=��l>0�>'�b��⋿"H9����������|?a��=�n-�0ƈ��� �A�	��":�>i'?ʒ�g[���^��>���=�W���?)���C>�u�>5�>������>,�*���b��d��$L;s��>�~�; 9.>�~�TP#�p�>�F�>��#�Ce>6��>zaL?7�|?H4?����>3!	?'�>gK)>-�=���>� �>�/?�&S?B�B?��>U��=Y`��mT���t�=�$����4<-�B��������%ͼD���Ql�<*(>�h�=4��<�!�=�Ç;tN�< �==Ѥ�>7O?��>��>�@�a�&��2[��3q����=%�>̟�>��>��?Y��>��>cy>��M>	�L�8	����>�j%>,�l�har���<�~�>C��>W\B?+-)?�j�='�����d>ղ!>�i�>�&?��!?}��>��=>ܬ`=L	���ӿG�#�)z!�
0��_L�S�;��<�l�I��J;iL.�����C��<�^>�%�>�-o>0�F>�!>�%3>���>�YI>��=hR�=�$��X�9�tD�R`\=����P`<��D�e�����'��=Ж�>He��tM��*��ʼ��?��?��?��Rͽ�퇾�߹��|���x�>A�r>�f�>(��>@��>����ȄB�@��4&��?��o?q	�>���"��=j����p����>?m�>��V>��=�3X���žo:��7�>�?"��=�꨽	�8� 5q�ۚ�0(�>�_>�w��ꪞ?#Jc?� �Z�X�]t�����>1�=���l����\˾!�}�s[
�Lu���M��k�>
N>�̫??@�V�=���<s���3���jt�T����M�=?�aU>�;<�h*�X������}���h�=`v���D>�]�=�8?�O?�ƙ?��,?r9?.n���`?f��>F�0?��>��3?�f?�t*?@%B>)�>��Z>T2��|�r����������d��_뼀�W>���>e�R>�젽v,���n=:���pj�����j]+>tI	>�x�=���<f�8=y?�>�A@?��۾����b]=�z���>��?����}Z����>Պ>t�>e�?Qҽ�/�;���e��/Vc��$?��Z?[��>U]뼍~}��@���?���>KV�>����i��Ɂ޾�������Ą�>���>p�>��e>RQn?�bL?d�*?���B?3�73��s�H���v�=Q��>�A�>��!>�Ɗ��o8��p�x�W�����⢽��d���=O�a<3�=��>� K=���=y�@=d�H�bNt��û^�@=�J�>��>��?�*N>�'�=w����Y��F?}���T������dmҾYx�s]>8_>>i���-?hs9���i�ц��#P;�V��>.�?���?��Y?V�g�Y�߽P�Y>V�*>��=��:7�<���
�-����3>/�=�7������*�T=�;>��~>]��(辤�0��D��ea�I˽� ���V�ž2�
�HO�������d��Iپ�-��n��XE��'�'
��c���4��n��?���?�l�>f��i���L,�7"����>]��&��N�b�r7A<[t@�98�3���p�z%��.O�YV$��:�>ta���䀿4Ne�������r�>Z�?�����i��|�_���ٞ)=ΐ=Ј
�q���M����/n�"(Q?l�?�3޾�| �5쬽\v>��>�ƪ>����(ԾІ�<���>:��>�?��˽�����ߛ��S=-�?�2�?m�?��n=%<�5�ξXƽ)?D�>���>����VoнΜP?
%Q?f��=qDH�yI:�����#?U�u?8JZ�;v\=2��>Y�>� �
j��s�=��l����=}�F>�.��j�t���ؾ�|���S����=gf�>+�~�ݾ��>���yJ��E��n��{*���<^' ?x��ȕ><l>C�>�t)��5��L��ļ�jG?��?.KT?@54?p����+�{�c�"��=-`�>�}�>X��=����>��>?�㾿cq��U���?Wl�?#�?i*\?�\o���߿Z���9��Ȭ�uuV=?�-=��K>����V����>5����!�=��<�W>yz>(>U>��_>� >)���=(�Ǎ���К�ZK���!�VJ+�C����)����� '�����(����E=aZE�A� ��_�$�E�X�Z=�xP���1>��+??�͑>᭧=���>7�������nUk�B'�z��т��P.��g���`���.���_���v�[���P�>��=B�	���
?;V��<�=��	?�~>��+>��>oFv>���>ؓ�>���>��>1>F	=5��>�$�>\E���+���f��o�.�@j��і?�Z�=��?��gd���>����BҦ����>�F?s��R��A����t�>L��=,l3�q�Խ,�N���=�t�>���=� ���#�|b����P"�����=2˖<wo�Qd������=���>-Ҿ,�>�?G�B?�	�?�
S?�;P��Ֆ>a��>���>�}���,�>�$�>�v�>�-�>GRa?ד??���>m�>��)����'[�,t���^q=0Sr��eR�EŽ#�1���H����Z+�=�;=��s��.:�d��=t�q>��3>r��>A+B?]�+>��>'��tF�9 U�9���#�>[c�=AL>�K,>s�>x��>� �>>I�=����ξ.!�_��>���>7H��f�|����<���=W�>a0W?p_?�9�h5澢 �=䃕�X�m>C��>�&?]��>\��=<���X��e�l����#��m��<Q�8�S���ɾ�F����b�B�O���_�z�����>M>���>�̖>� �>Ⱦ�>���>Mi3>pv>��+=QL��CJ�=G]c�S�P=���W5=F0�>���/5(������\��<�X=��e<u��I�?��!?Z숾��v��7�e���lž_P�>�#�>���>��|>z�p>���t�A�]&���D�C��>
p}?�?:����D�<^+���;ռx��>��	?��>�Z��u/u��žf�ܻ|T?�E?=t�>l}:�f�D���Y�, ľ���>��=�\��/�?��t?9��I�8�}���Q�%��U��=�t=d��KZ(�����G�k���\�X���Y>�r�>7ѯ?jǋ�'s�=�f���3�������?�ى�=`�=��?���>N��M����(����[þ맡�-�,>��q>F��=ߕ.?��X?sπ?�74?�*?��;� ?#r?�!?��>/�/?��4?2{#?Z
/>�@�>�%�>�)���DV���p,:����Ƹ*>Lb>J�>�uW>��5�il<N�=��3�A�p��(C�O/=+��=/H�=0$;=t�z=���>�?ۋL�_
��0���j�5��������>�Lļhe���Ի�߾ >�W>�>��6?��>9ʻcI�2{6�fL�?=!?c%?F�R?��Լ�r�<�)�����gn>N��>EX��1��V�3�Js���@>��>˝�=�>�>|Ei?Pv[?�;0?�v��)KS���M�8D�^+�n]->�?�^H>D��>����]�L�}��7q���%m�=A拾�P=
��=M/�>v-�>��r>#v�<6�$�f>�"=7��{�@�J@�>��>�??�|�>��*>�_��#0�a�I?yɠ�8?��;���FӾ�J���>z�D>�� �69?g��TA{�R���>�C��>��?K|�?�Ab?�EH��K���[>B�U>$�>ğ�;p<���0����1>���=��x��.�����:��Y>��s>%9���+̾o����I��4����\��E���[W��xr����$���8T�����۽˘����`#�"X[��:۽��Ӿ�ƾB5q�!��?�<�?����mU���I��X�,��#�	?�����T���B�����<r���K��{����'���I�)�,���>03�=�T����i�K'��nݾh��>~�?
�%�Vܼ�4����=���K�@=9C�&����
��zƶ��OT?`��>˲�o�~=��l>��=�A>]�>3�I��H'�M3�=��>�k?L�>U䩾樱�����)���?G�?�
?&r><@@�	W�G�<��?�_�>�n ? ��������ʾĳ3?z�J?��T=��ƾ�<��5��c�)?�O?6Y%����=���>��>ѤE��+��WMp�~���PYݺ�ft>�)>;���fC.<L���LH=a0>�\&>/
�����*8�>��¾i�Y���c���r�
�?ޅ��"?"��h�>�ć>�Q�>>=����v�j�B��<q7f?kٜ?Q�?}:?�s��;� �'�D�cM��	�>��>�F/>0���o3�=7a ?0#y�3�f�?�)�U��>���?�g�?D0a?$tV���Ͽ4���w��}��\T+>��=z�[>]�R�=�A�<j@�<��;��(>Ƥ>O(u>�Z�>�g>b1Y>�4>����@�$�Lz��(��G;��1��E�B�x�Q'�V���X�$�W����x���~N��:��j.�%j.� ��gn���:��O���o?Ev?A^>6��=N�>����x�<�����e��2��-5:����.��w�>-�&�����9ѽ�����,�>4RL>�ȷ�;?��O<ST�FW�>�.�=~}X>��g>P�+>��C>N��=�y�>�x0>;�>��]>h_�>F9�>WƆ�w"|����'���;��]?��%= Ƥ� f��侀?n�!|>,-5?���>:�.�8����������> �s�cڔ��6w�{Ԭ����>�w�>�Y�>6g�[����h5��	�v�>ή�<���i[ܾQ�I�BG�=���>�)�NK�>��>e=F?��?�*T?�x���7�>E��>�ڪ>,�b=+�=9`�>�|>;��>��+?�:?l(�>�ܶ=��y�&�=���<&c����6=ܟ�<F`��x�#{,�-�6� �=&�=%�>���=��>*��=����C<;�1�>[n<?�/0>F��;!����,�PsY�Kc.<O�>Ke�=H!>6e�>�>�>=�>4��>��>��3;��������s?�'�>~똿ɒ�������=�x@>
څ?NB?"#�?c�v\x=��>�[l>w?>�J?���>q�!>m+5����g�%��Fi�E�{�����(h->vL�:A�������+�G����nS��8�>;j�>�ø>��z>��0>I�=���>"T�=�>�F>[��=��=�8m��fc=_E��8�g>�-��,5�<��付0�R����&�;�S��R�<%��<�1�>)�!?�O��OH�}`���T�����>���>Uƥ>W��>�^>0��{�N�$�������>��?��?�KK�N�Y�t�=��=�-n>���>���=��߽~�[-���q�~Q�>��0?�g�>�Z%��@J�C�8��W��%�>#>�`�f�?*�?��#�!�Ž3�� �s��Sᾭ�2��;�=w���7龬����`���Ҿi�������9�>L�>u��?S|$�ao��/������Ӌ����� �=�}�=���>I \>c��:�Ž�����ξg����m7�ߨ�=��=�`f>T�[?��L?-��?}�)?�Q?�>Ҿ(;?n��>bw8?�*�>��F?�\?��?�X%>p��>��x>��<!w��>ݾ�l۽�r=i��>�d�>	�>}�=Q��=�Aٽ&~#��Y����+�b����I�<��=>��>�k�A  >�7�>b?R�V��?�|U��n�>��z2��v�>���=#_>�q��nS=F�|>bО>��?�>�y>4�ܾ����)'/�"�׽�8?�S?
O"?PV۽N3�>�;��ʻ��I��?դ>���>˳侉Y��A㢾�sN��a�>�o�>��X2�>�te?f�h?Q.8?��?��/i��o���c��輈s�;\� ?�՗>��F=8�4�ɩU�p���_�2�9�� �W����:,=���=�� �)�n>G<	>�(>��R>z��=Z�m�5�=E�����>z7?��L?>�>�d�>���)T9��">?�����TE��[��?�,�$Z4>_��=~�?:Iu���>A��j[��F��Zp��.�>��?�$�?yo/?�)޾M����n>��$>��T>|�<I{߽m:0�u����ϊ>�>��ྮ~$�E_>=�t�>z�Z>|W�o�����:�=�q���=�4�.�[ž������\K��E��ƾ}��=�$о����N��!wսܑo���S�
l���4о�ZȾ�.�?vC�?��)=?˾�]P�Kn3�ci��|#>����=��b�)}�3):��ٿ�3CK�ؿ��E���>-�e�u�?]��]��!Xk�L˾��>���>K�2?���0D�R�&��������=��=a��e������Qd���HT?�$?~�׾p���4��=	��=�pG>9��>��(�S>���>�u�>!�6?3+Ǿ>/Ŀ���A��?�?���?z�-?�>O�<��(
��r�=ԯT>`P7>��>u�H�\R��w�&�?�rV?�6�������`y��#��5G?*?�?��x���8>�?��>,��m���;�(���aG=�~�;cm�>�G������T���>�8�={׫=�[˽괾3��>�{;��[�?�X�0��Ͻ��Pj� L?
S��j�=�%>�:>Ax+��
����}�u�p��tM?zZ�?8M?@;?VE��V�M�ҽ��H>vq�>��>q�=pнR(T>�1�>�eg���_�K�'��>ze�?z��?�(T?��`� "ݿ�W���f����¾�2�=�*B>9��>��j��D{=��k�J�E���g�L���!��>�l>yo`>x�]>Cvv>��=}������4��������-�a����3�@���˛�d��3�Ͼ��=�ƽ��:��>ɽ �(�Ԃ>��\H�NRe���3>e?w�>�y>.j�=@�>Δ�����������0���_)���,����(s����?\����c����H
���1A���?�~>�=��6�4?�"1�9Y�<�&?�{O���>��>u⓽r´>0>�W>��2>u�1>n�k>=�~>M��>1֋��W����0��������?[D>�v��Ƃ��������h��V�>�IE?_¾�B���\E�o��>�s;�9U��?���@�Y=>oY?ߑ>� ����[�5+��	U���)�=�>g2�B�=
H��9j��x�u<_��>nϾש�>�
�>ڴ:?��b?*JL?43�=�>b^A>���>1�=,��=6e�>��>-e�>3N?�[2?Ћ�>+��=���'�0Vڽ�N�a�$=��
��i�<��=�ּ���rs���F<��<�X�=(vC>/O%=������<��>��?;��>Z��>~���iC��_�������>�ך=��>k�?��?�7?@H>�.|>�I�G�ľ���Z��>DС>%.[��*}��Tx>�?Y>^~C>Pag?@�?-��k���l�u���
>�0�>Zg?z1?\��>�^��4Q��S�'!�|��Tl�nl'�G�/>'�J>/Qֽ�o{����Ua����޾��e�A~w>K�>of>��<>9�D>��(>���>9a,>���=��=����P֎�ׂ��D�%�)C(�"�>ө�=�X����=
h���	������l9XԿ����=��>P
?-���!B�����;�65���ƾ�?�2,>��=
V�>��><Dƾ8ZJ�nKվ_`����?��?v��>�Ͻ�W1����
S�>�F�>�,$>��>��ȽIYk��!�c��=���>3��>e�>KD���y4�ŀt�gGA�>��>ya>���ǧ?��?>����=���Ux��Va��F��5��=�t"�D�ؾm�7��^� =��Q���i>���>ˑ�?Fs!�2)=?��������V����X��Q��>�LK>�ʰ>)�>��;Q�nb�w'����>n5���Q�=��>'�;?ψO?pZ?e�?w�I?6����e?��>�%?'J�>��&?�*?��?-7�;-	?���>��(>li������x��<�Ď={F^>�c,>4�=%k�9�����<�ݼo)M��ھ�n�=�¸;�9����>�@>���>`@?5޽N���*��!�侮����3�=j�b>��L>�=�P�ý<I�>��?"h
?]3�>���<�1��5�;R��ǵ=�?�/?^��>4����c�=X�ؾ�G�E�&����>2�%�?��W��Sf�=R���&B�>'ĩ=ֽ�=x��>vui?a�L?l.?;4Ľ�3E��(�{9����	y�>��>��=��Y=Ⱦ+V�nyw�˘g�B�/�e�=N�۾��	>�	>� j>C�>��=���>�n\>��>��Y��>@ذ�yG>��>6U<?��>�E>+#V�H�6�&�G?���H������ξ�*���>�L>1���C?9�\w�mؤ�ď?�J:�>ʤ�?� �?�a?��O����TrY>5�P>�n>��<xA<����oy��4>���=iw�y�����<0`>lko>u����eɾ:+�O�"�)ƿ��W�K
%�f*���r徉?��7�۾��=�Ȥ�4�Y�������侤J����7��T�='8���������6C���?�e�?�R3�"T���D�~ �m�-���>�,U���:I����M=C�@�S����U��
���<L�H�f�*�-?�Z�[���-�l�1
�y�9>���>�9?h4�ĭ����J��IQ��Y=�q���*!�����۬��v��	[?�?�5Ǿ�]���>�e�(��>�¸>lٚ� +��1u>x>�>�_�>N�g?��־<�¿������/�?���?H�1?SgO���I������I����=�7�>a��>���X��>ɽ��?��2?:`�<�n�򀆿�Gݾ<�?�i?}����*U>,?7�>^AO�ըx��v��I����=��>���;eQ�.���k��'S�=&\�>���>������4�3��>�{;��[�?�X�0��Ͻ��Pj� L?
S��j�=�%>�:>Ax+��
����}�u�p��tM?zZ�?8M?@;?VE��V�M�ҽ��H>vq�>��>q�=pнR(T>�1�>�eg���_�K�'��>ze�?z��?�(T?��`� "ݿ�W���f����¾�2�=�*B>9��>��j��D{=��k�J�E���g�L���!��>�l>yo`>x�]>Cvv>��=}������4��������-�a����3�@���˛�d��3�Ͼ��=�ƽ��:��>ɽ �(�Ԃ>��\H�NRe���3>e?w�>�y>.j�=@�>Δ�����������0���_)���,����(s����?\����c����H
���1A���?�~>�=��6�4?�"1�9Y�<�&?�{O���>��>u⓽r´>0>�W>��2>u�1>n�k>=�~>M��>1֋��W����0��������?[D>�v��Ƃ��������h��V�>�IE?_¾�B���\E�o��>�s;�9U��?���@�Y=>oY?ߑ>� ����[�5+��	U���)�=�>g2�B�=
H��9j��x�u<_��>nϾש�>�
�>ڴ:?��b?*JL?43�=�>b^A>���>1�=,��=6e�>��>-e�>3N?�[2?Ћ�>+��=���'�0Vڽ�N�a�$=��
��i�<��=�ּ���rs���F<��<�X�=(vC>/O%=������<��>��?;��>Z��>~���iC��_�������>�ך=��>k�?��?�7?@H>�.|>�I�G�ľ���Z��>DС>%.[��*}��Tx>�?Y>^~C>Pag?@�?-��k���l�u���
>�0�>Zg?z1?\��>�^��4Q��S�'!�|��Tl�nl'�G�/>'�J>/Qֽ�o{����Ua����޾��e�A~w>K�>of>��<>9�D>��(>���>9a,>���=��=����P֎�ׂ��D�%�)C(�"�>ө�=�X����=
h���	������l9XԿ����=��>P
?-���!B�����;�65���ƾ�?�2,>��=
V�>��><Dƾ8ZJ�nKվ_`����?��?v��>�Ͻ�W1����
S�>�F�>�,$>��>��ȽIYk��!�c��=���>3��>e�>KD���y4�ŀt�gGA�>��>ya>���ǧ?��?>����=���Ux��Va��F��5��=�t"�D�ؾm�7��^� =��Q���i>���>ˑ�?Fs!�2)=?��������V����X��Q��>�LK>�ʰ>)�>��;Q�nb�w'����>n5���Q�=��>'�;?ψO?pZ?e�?w�I?6����e?��>�%?'J�>��&?�*?��?-7�;-	?���>��(>li������x��<�Ď={F^>�c,>4�=%k�9�����<�ݼo)M��ھ�n�=�¸;�9����>�@>���>`@?5޽N���*��!�侮����3�=j�b>��L>�=�P�ý<I�>��?"h
?]3�>���<�1��5�;R��ǵ=�?�/?^��>4����c�=X�ؾ�G�E�&����>2�%�?��W��Sf�=R���&B�>'ĩ=ֽ�=x��>vui?a�L?l.?;4Ľ�3E��(�{9����	y�>��>��=��Y=Ⱦ+V�nyw�˘g�B�/�e�=N�۾��	>�	>� j>C�>��=���>�n\>��>��Y��>@ذ�yG>��>6U<?��>�E>+#V�H�6�&�G?���H������ξ�*���>�L>1���C?9�\w�mؤ�ď?�J:�>ʤ�?� �?�a?��O����TrY>5�P>�n>��<xA<����oy��4>���=iw�y�����<0`>lko>u����eɾ:+�O�"�)ƿ��W�K
%�f*���r徉?��7�۾��=�Ȥ�4�Y�������侤J����7��T�='8���������6C���?�e�?�R3�"T���D�~ �m�-���>�,U���:I����M=C�@�S����U��
���<L�H�f�*�-?�Z�[���-�l�1
�y�9>���>�9?h4�ĭ����J��IQ��Y=�q���*!�����۬��v��	[?�?�5Ǿ�]���>�e�(��>�¸>lٚ� +��1u>x>�>�_�>N�g?��־<�¿������/�?���?H�1?SgO���I������I����=�7�>a��>���X��>ɽ��?��2?:`�<�n�򀆿�Gݾ<�?�i?}����*U>,?7�>^AO�ըx��v��I����=��>���;eQ�.���k��'S�=&\�>���>������4���>��龺E�I6�S=��)���>5��:?���M1<!W�>�+�>LBҾx⎿T&s����3?��?�M?8:�>V���C��p�<��?q@?� >�->kE<���<��>�rξ!�$�����ҍ�><��?��?��3?67��_+忕������8����=�>��> �K�NU<>��.;�*��pG�;�{>=;�>��U>�:�>StC>ޝx>��X> ���5m �Ҥ��唿�'<�-U��>޾E.�K���h���  ����8&T��7���ܽ{2���q�q�
������/��>�b?��?-�>�i�>��P<x þ�[?�M$��0�i��>�
���򾥝侴W��!
�@dn�P-��A4&������Շ>u�=^�>]X�>.۾=�W�=G��=x�Ǽ�oo>��>�>i����;��7>Ť[>���<w��=�D>�Q�=���<R�J�� ��J�d����H�ϼ���>���HF>��� �ܾ؍��� �>�d>�j�>G�.��W����s��n�>��y=o�Q�J�Y�{G�="�1>��>-Nd>������=�$�GCƽ�8�>X�:>O �>vR�<���Ǌ(����=8��> ${��ʲ���>F�?iԨ?�S�?d�1?�0.?g�O���>�H�yl>>�Q=$�?�?s&�?�CS?ק:?�2���T�6l����И���O��e��:��"�?�=r��=ΜX>��>ކ�>��C>��>�"�=���=X��=���>h�E?AO�>�j�>op�;[���=�}��ʡ^=ɻͽ1�?\�>��3>�|�>��>{t�����Q	�%V�����>@��^Rt�)s]�(ɠ=���>�4?��V?(�?�Z��
�����t��!?�	?���>��>zk����?K�t��α5�a3)���½S"ԻF��=��ܽ�J���Y�	�nX��U.=\�{>��>'4A>�a>�>@>��>+X>]��=a�=馍;��;�'�?%��Ә�=/��@#���r�p&��^�߽^�	�b���1X��1ϯ��"?� ?q� >kO�=�IA�K=��M0�eh>� �>­�>�?+��>)þ�Z��cC��s��ݹ?o^u?��>�**���=rnýq>���>>�
>_������F�����e=⛞>�U�>�4�> ���Q���m�[U
��N�>~#�=���è?c�P?�̔�;4����5��7��O	� �x����>�@>�%;��#[�a.�T����:��F>_�L>�)�>�?��>��>'�d��Z��_���K��)l=��-?��,?��?�Y�<o��Ё��Kt��^�:�>{G>m��=���>)��>�&�>�=*?���>;��>H��?/P<g�>��>�i5?X&�>�G�>�K�>D ">�.��������0J��Ċ��Wཷt=�16>��i>L�*�q�=!�=i>�̋��;�=ԙ̽��2=O�1>�ɽF�>�yE>��>�5+?*�,�¾�Yu�7��v�=$�%>���>/��=&�վz=�z
�= L�>�~!?���>�
[>g�����Ҿ�js=�~?��D?'�>F{��T���!��$ξDE>8�h>�=�?V�����?�a�l�<?�>���=�G>�T?C�%?���>�|�dH� �l��LN�d�w���>�"�>�@�>8.s=��d�
�D���g�!���}��t�U���̽��=G��=(�=.x,>vA�=U��=���=�Ň=�V����;�@g=E�&>�D�=^=?��>>cu��읾�e����;?q������nRw�; 	��|>��>q�>g���L�>��Ὗ.���H��>�W�3	�>ew�?�Y�?*LG?���l�ؽl}y��14=J�">�I=o�̽��D>�Ӑ>R��>1��<Z=��j���h�={��>���><=���~]�����6
>�rҿ/6����y��B�[�
�������C���ɜ<���������2�>�؃�b��=�����Г��M-�?�j?�N�=Q+_���@���ξ����˿��)O�����=m��Y���#�!��a侺������a��'�2��;���>&�7�v2����i��K�v,��ù>'3?8����܉�VU�����=��>h
=�Cľ?�o�����[9ջE�n?+�.?F����'����J�@Ӄ=��?�N�>���>�<��h���%>��!?�1?�*��L{�����xR����?�q�?��G?�DJ�=R�[�������>��?���>�e��ʣ��b�;��?��#?���<Tmɾ�}��R�x��i?w��?��P�>�8>{-?秘>��=s\j�3��I����=E|�=��>��<;���e����Vл	;�=�ͻ>g�������>�\꾇�N��DH��r�jK�u�<׆?���m>�lh>x�>��(����K����:� �L?J��?A�S?a<8?���I�~ݩ��_�=뺦>]Ƭ>7ΰ=�M���>]��>V=�Xr���3�?�3�?$��?�IZ?�lm�8-�H����þ�"����=���=�3E>
BR��V�=���<�P�i+��y�k=F�>î>�	>T�>�,�>i@>����{�*�ɠ��������S�F�����Ѿ)�&�F�������!�u�������G���oZ��p�C0����˽�۽O��p�=@�c?G�.?�L??���=̶V�H2��e�&�����R@�6����(���㾻�����=��=�<j�CX�p$���>6��<�	#?=?a�>�Z|>h��>�Q9��O��R#=��6A=�9=��F>O%�=C�>�U>$��>�f�>��}�6h|���2�a˾�K�ި�>^]v�����&"�w�w� ���?�.�= ��>b�S���6�y=�>�)%��ʾ�湽�ű=w��=d�>�Y�>��:�Ch�+��x���0 >%@f>fWD> G`>?� ���/=Э�> �>���nh�>c��>z�z?,;�?Q�k?U+�>�ga?�����5f�I؉�>��$����>��>,?�S?��#?�_<��¾	�M��pZ�5�U�&��1.�l/ >�L�=XH\>�{G>O\>���=gn>[H�>�(=kņ>A�=��h{�>̑.?��>��J>̺׼�B��`�UxＹ�;6�p=�w?t�?�=�>�>I.�>�/&���<�{'��d��7�>0�u>�;]��"d�?"?�؏>���>�)?	<?�}���Zܾ܀F=/U,>6t�>m?��I?ufH���=��'������,��Z�v���n�>q�>�x>Ld�>j��%n��䦫�N�-�=E�>�y�>	l�>��>�����>�x�> �#;O�z=1>�=���}ｬ�'�J���[-�nR�u_��������g�@O���W=�H�2U5<�4
?�I?\A3>�}z>�@�=�Ø�����{>�`>>��p?wO�>wើd�ݾɴ���K�>�/_?=�	?��<�Γ��Կ�n.1>!˕>�B�>4?�	������{�������O�{�'<�X�=I|*��� �7\E�{y����>�F�=*O��O��?�;?��3�� ���rN��Hþ���0��ɶm<���k�F(�jݾd��1����;t�ֽ���>N��?���\>
r)��b��� ��
$����<��>�(?�$�>G�q���#��@!�Y����=]���P|y>�e~>��>[M}>>�?>�>���>�?�m���%X=x�>�Y�>�>�Rw?���>�B�>���>�%�>;��o<��,���d��=�(׽�5=:.�=zK=`�M�{Z:>]����0>��6<j�O�	;�%T��5�<W��xd><�0>��?�u?�z��'��խH��.�� ��=Gnx<%]��)�)>���ѕ=�m>ݰ?}�>x��>�Q~��X���v��W��DN�=�0E?�)?��z>��,>n�F�ä��D���,<��>L�&�wC�=S�ľ����W���b?V��>����>��[?�0?Y�>�����M��E�mv���xu>;�+>F��>�+7=�o,=eoQ�ؕ0�2����W�l����B�45�=��=� =���=��= G7>��u�
]��J����=���K{>��Q>䒫>�<�>�p�<���۾3�I?���1����F)Ͼ( �:>H�=>����!/?j��~�c祿�=��h�>�Q�?���?�Ad?ԌB��v���Z>�PU>�7>�,<�{>����|�����4>(��=�Sx��
����;��^>�|{>�&Ƚܻɾ�.��I��穿!�ƹ�����!���	��]����j=�x�t�<����+.�Y��� ����(�������:�rm�q,��b��?˷�?.�5>L�c�qh�aPT���о@D�����_>������<�Z������ȣ����k>�\7O�g������>ۜ=����/�}�f�0���x�J�E>�'?|gǾ�ܞ��f�._2=Va@>p"�=�`�Q��������?��N?I�4?�n�T��u��E>�0�>���>��X>	�������P�>o�1?�+?/u��{��=	������+��?;��?�l4?@��p�?���!�-���b>t??��>Ά��.}>(�����?0�4?n��=��n��"0g��[�>�{�?�8���>��?�g�>HG��"��է$��ǽ/�t�mV�=������f��Lj;e�>[�>�J�>{;������>��f�M�5G�&��z�m�<�T?�����>!Ui>&=>C�(��P������;���L?g��?��S?��7?�������᥽��=7��>j�>R�=&���>��>�]��r��^�~�?��?���?�|Z?��l��H⿭5���3�~�l>�b�=Ћ�>�W=m_�=����\�*�H��<�۶>��>K�= ��>@{X>�q>8�>6G���,�`ᦿ:�����7�G�̈þɡ����֤�"~�f�ʾ����������Q�G�p�-��D�s��|�<��^>�+J?	�>?���>o��>��=r,��O�۾�� ��\@�NϾ��4�jT'��	Ҿ��>�T׽>�߽�p��@侧��>� >^$?�"?��>�>ė?��)��<���=���=L��=���=B�>�/�>^��>��\>�6�>R�>, j��?���15�����v�=�rH?
��~4��?��",��#����>��(?� q>��=H��^g�O�>�ׅ��P�z\��f�.
�>=m�>��=FT�>RB3���8��<���<E�Q>�a�>��?>��j����=�"[>�-T����{]?�B�?�%�?
Oq?+B?��?�����E>ax��9�+>H,�<f&D>?�?@�?凞?*�1?��r<kq��ː:����
�P����ս7:��r��:��=�z>S�T>���=�[>Y֤>hIP�w��=�4=g˝�0Y�>�*0?��>��>�#��j�'��P�LA��$D���?�>X$�>��>]�>v�>�G=d+?>�Fz� �����	?+�=�`o���k��H��5>
�>�`\?�/?��l�>\Q����=DC#<~v�>�-?�I
?e{���>c2t���T������|�d��;��=�=z�.>2C :A�������3��������*�>Ư?�3O>-�>�>�>K>G�>��>��f>��=��$>]�ٽ�Խ�&��<�v�D=��>]zF����=+=�<���5��=ܒ��������u:��}n?��?��<�mn=���8-��O�žK�>��> ��>�>?��0>�D
�sqH����[�;�Z��>�=N?��!?ED"�ƕ\�w`����u=�>S^�>ø�>�Y&<���l�ξI�%�;;>jT�>��i> ~�t)O�r7b�L�߾,��>�3�==�U=e>�?�H?����iN�=�B�L#�\��v����=V��<�E���3��%!� 9��
���~K�*���E?Hu�?V[J��|�=�S3�4N��eє�c�����1�ow}>��!?�� ?�:�;�]	��$�f���F���e��>3��=N�>y�?ǰ?o9?1��>a�>���yj�>5[1>.U�>?�>L	?��?���>]�_>:c0>
W����(������a�)�������=��>cb>t�O:���=��3>�j�=��<�	d=�p�=΃L�1Z�:�<�:�>e$X>53�>6�?�ց��˂��b��̕��!�6>��ͽ�� =OE�=�\���A>��~<���>�� ?���>q�����"�ﾫp��~H?��i?�φ>��$����p`�������<��@>�S����7;��ξU��⼏�;�>.ǰ=E}>�>�m?�U?�m?T�D�c��8h�oS��A(�l�?Uޯ><�=�������J�����]��޽\)�եt=�"=ˊs>ȭ�>6^.>c�/>Mnm=���1^�|�T�5���|�>ߦ�>3�>$��<�?>��ľv7پ�I?<o����'��5rϾ�6��B>�=>4���)?�����}�M���>=���>lX�?���?�1d?�2C�v?�M�[>DU>��>�D2<�M>��������4>�8�=Cz��ߕ���;!]]>��y>mɽ�ʾ�"�9H�?c��|�3�mz
�"�+��>[��5۾�
��8`־U=X>o����8�˩ȽC�Tڽ���Y$Ծ}��kY��Κ?��?�H�>��ۼ�7A��R�|��B�ݽz����>��ľ�#2�ӧ��� �*���5��<1��l��V
/���>\vA�FL��U�x���-�ֱu�F�1>)>2?o ž-f�����E��=&0>(E<=�Q˾u%��R�����
�BsX?�>4?� �e����6�	D�=u?��>��Z>��t��:�-Z\>ϱ%?Q�+?�������ì��?�ؼ��?#�?"x5?F���)�<#���F��x�>mF�>L��>��E�@y�g �=��>?�G�>9>m�K��V�t�S�۲
?�j{?۠7���=��?2��>�"}��9����n�gCԾ�n���=\���x$��_G�:tʽ�	ؽ�� >��>�U��)���>����L\�9��H-���`C>&!>c�@?�5���q��{l8>:�=e�A�Pϕ��v�ᓢ�?8G?迲?Mr�??�?n�x��톤�`���З>;�>��g�e��V�>c�>?"	}=�}��zy���K?3/�?���?��~?�GR�]�ڿ����TY׾)�ƾ���=-�=O�">he��tp�����=�*=�E>~�>��>��>?��>q|>A [>e�����.��(������s5�;��Vm�Y��'1�効�˱� <پo���ҽ�#0=n�=����$��z]=��s�<Z>�1?�P?��?@��>B�'=e��=�쓾Hj��}�#��쟱�"�"�������>�<uό<Mj��;r�U5+�[�<t�X����>4�>J�>�?H6?w�(��?μLǝ=���ε�=X�=�9<>��=}γ>��6>��>>���>v[N��=���{b� ��Q�>h;>�����Q�>aw��D��da��2$?�ۥ>p/k>/�b��d���S`�P��>��D=�A�������9���>D��>�tc>e�>9�νI:��i'��K�e��W9=$��>�ؽ1�=_Zȼ��T�~��>]�m�*\��.�>��?�b�?ܴC?6�K?�M�?�<R�ʈ?? D)?�d>�Х���(?De?��?6)�?t�m?A�";�惽P�y:zy����8=Z�p<�	��kF��+��Ϸ_�Z9�=p�3=�@���G�|}�=�ڵ=c�Zѣ�D�F����>^�,?���>�{>+玾uS-��
#�Zΐ��ء�4v�>��v>�|K>�"?Kd?j낼N�7��b��
ƾ����>C�=c�\�f]Z�����H�>7Q?�8�>�-�>�?�=����˙ ����V<�>q�?�+?����.�����.>�t!�_���a�(�Q����������t(=�`1���-���&���h�H����;q�z��=��?�"�>��>�>�>Oa�>*��>��g>�*�=�#W��p�K���'׼���<�!�=($�=�.��Έ��v6=-���}�{�iѽc��1�:�1��_?b�?ugh=�X!>{��<�G�r�����>!R[>I6X>�|�>
>�޽�6Ii���b��D�����>=�M?���>�&��!='\���=�lb>{�>�;�>��=��L�3��3�i=�I>�~{>jđ>n���7Y��@?�۶پ؜�>3�=��<��?H�0?
5P��B�Va�3�F����ox�v�=s��>�r
�a9��LJ�c� �-槾h��F�Ҟ�>��?�DǼ�ߖ>�\�B$��頻�~���~Ƚܲ�>�D>�w�=��=fIv�?�2��V��0��x�Q�k�}>�(1>�L�>�?�Z?H�>�>Y̑>�X��l�>%q=a,�>��=�0�> �?VC?��`>Y�=)F���W;�<_����>�!�Ǽo\+���=�ߒ=z�p=P�>ʇ�=���<$����սL����=�P<�؄:�A�:���=�>�
�>�m?)�� C�؎ɾr
a���>DG�Uj�=?��>V>�:�����=I��>2�?�`>�
a� 2پ�����X��I�¼Y�=?�g?�(�>辒�c�˾I�ƾrw9������>}P=�I�=Ox�n�Wþ"6�>�c{>Z�����)>��^?�dx?D��>e�h����~�J��F=��ѩ�C�=�Bs>tn>�;�>I���n�3�3t��_[��p��lm��2�E����<���=G%>��.>Ϟ�r�o> O>��7�'�k�/��$?нx�?�t>	�>X��>_�G��jg����{I?7�������;���>4A>���7U?�\��}��'���=�n|�>�?/Z�?�Ed?�?�Op�S�Y>�[R>��>��+<��=�y���僽4�5>Vt�=��w��ו��{�;�\>�z>oǽU ʾ9�⾞=��Ͽ-�V��[=
p�1-վ���rK¾�l��,���}w����;s�ϋ��w�4�4�ƾPV����������_�ŏ�?Z��?��>WY=�[�R�_��/1��w��$
�4�>�����=t�u�JА�b
־�徊��'���!A:�$#�>>[`�su��q�p�&-�OB><�cB>%*4?Kt����¾Y��,Z=��=�H�_A���X��~���ӏ��BF[?z�4?�n�������FW>J�?��>r�>����)���a��>�1? /*? ��ꋿRA�����S�?��?�C?ۥ��y5?�������>�C?�k ?���xrξW�G=���>���>���>����"B{����p�>S�A?��8��`�>3�>�ڄ>i�ٽs�����r�����a=���=�+g=4?�G�B��*���>?l�>؂>���z���~��>���|GK��m4�w�׾�N����=2�?Y�Ѿ_z�=f��>�0�=�-/�ճ���׃�Lʾ�0�M?8z�?b�W?�b/?\S���
��?)�:�˻�C�>�ۢ>W3>uǦ�O�>��>�أ�M�M�ͯξ@�?�k�?¿�?B)b?�Yi���p6������¾om�c���Uc�=U]��~�=~(����K���»)�=Y�>v-�=��� �=z��>xy>�ʌ�7+)��̥��i��r�O��������Τ����4������}^ﾢo��"1����Ÿ��/����ҝ��W>�I���u<=yK?��_?�%<?{+	?�h>�n;����!��ٕ�Gn���}(�tY�x*���)�"�e=C��;1�Ľţ|��#�h�>�+��A_?��>?Uu>//>��>��>�,Z>G�=P�<�6L���=�.>T�>�*�>T��>�u>��>�+��&��7OZ�]T�����<~_�>2m���R>EBI�8���MX]�&8�>��?刦>D�(����r��P�>�΃<R>��A$��-��~>P>�ͩ>?�b>�C]>\�� *��/q�1��=��V>p�s>���=\z��f	������U>���O��q�>�
�?ɞ?�??��H?G�r?�p�����>@�=��{>��?�H�>�fT?�S�?�̚?|�?�t�<N��Iļ!p���C�G���]��=xt޽��%=�a<1�J>0LS>Н�>�#>sO^=[F�=��c����U�>��B?���>�@=�=y�2��F,�z�������>|C�>�>tg�>���>�1�=p�	=d�k���վbc����>K�>�|V��SE�H�l=��>��?��\?�?¾ŤY����R5�<�)�>��1?ɭD?�9f��v_�)��"��p�迡�?���A���F��fս��W��P$����<'K,�r����(�K��|C�-ݢ=��=�o�=U�=oË>f�>�W>��P=�+�<��,=D
^=���x�c=��D=Cx�<�Q�>��q>��W�"�ɽ�s>=˼;�M���v��p?4?&����FL=�}����a�u�I>�ҷ>;5?y�?�k_>^v �a�`���!��E~�4r.>ηT?ԛF?�*���Q=�d1��������>5|�>��>9��1d�n�ɾ��{>ӊ�>���=�7{���v��;l�[���z>�>#�N=5�<ǐ?��D?p����n��T�l���,����H=��ǽYm.����Sھ�#�HP�Ad���(�b�.�s�?��?����Za�� M�hVl�怿�W(�Vԥ�d��>k�2?�S�>���N�����@뾙_=���=\uq>A(;>�J
?�6�>�>��>e�=^�>#�����>�Q1>�?�?f�?"��>���>B��>�W<�ɼ��Y�Zɽ�r���ۼ��9=w� ���׽�xe>[ڝ=��T>�|�=�ѽ��6�xt:=���<+\�=�3_�$����;=j8�>��>�?z�s��6g��]m�Y�>�1Z=����P矽�l��ʺ�=,��B��>yB)?��v>�BȽ�]��)���ƾ��<��<'?��]?���>X�"��*(���Q2��਽#\�>Xe#�I��_?Ѿ(�%��V�>���>K�=��a>"�V?�&0?�\�>v`�'M3��w���C����Az>gk�>��>�9V>�r���<��w4�_���1��7R��dk��@0>�ټ	1t=��>%�=$�>?V�=#�(����=�,�=j���F�>�Sc>{v�>{m`>��>#�þ>����C?������vz���Ͳ���#=ӵ6>�T>�̹�u��>�N߽A|�UV���9�p��>�}�?_��?�h?�i�������I>na>���=�`1�K�g�55����P�L>���=�Pk��ra����=���>Ɍ>FF��Ů��Ͼ�w��7�ƿZL����9�6���ܾ�c��پ^7i���u���<��*�x׽ES��{G1���k�Y�׽�H����⾅0���!�?��?�U�>q7���4�"������M��h��XQ>A?�(���z�D����Y+���J�z�p�q�0�荦>�b������߲I�q�$�t����w�>�'�>:姾�>�I��:4�=&h�;�[��� �)���<���k����}?h�5?����#������8>4~*?��>ҭ�=�=��͍���8�=���>�m�>��&��㌿*����<
��?�4�?y8I?E�ڽp����<��ok���>�]?J�>��`=޾*��S��>�-�>|C��7/�.¿�,5���?F(�?�DF�*C�<!�?��>��ֽ�2 ��u���$��TL>7U�=��z=�=��w>	�=��>v�?��>�%�4S���>��(��j��K�#��*��'�>&n^=2�%?v2�����=��=A T>/����O���R��/v�>3�?>A�?�K�?�b?����_��)�w=:f��-�>���>�P>I�5=�n�>�q�>~}ؾS�V�$����K>��?��?�b ?]|վ�z޿����p��KK��,<+�	>�+q>�y��Y�<-=gN���|t��򩹊5�>;�+>���=��=�>�ݜ>8W���#-��k��������?����~]۾.\>�ܷ�GþB�-��V�gT���>H{�;�
�� ������m ���N���9>ɕ??"�>i�V�"ڗ�	^=�樾��
;�'���n��x�-�;������c��q�N���Ͼ�|���þ��/?ӝ�*�����?�a����N=��|>���=��>�Qe=*�V>��>���<��>Ǥ>O��=��=p��=�2>	6���[S�e������=f��k}?����-�3��4��1'�C߆�o�Q>
��>ߋ�>%{S���
�G	��T��>W9�<��[��3���l>0�>�$V>;ƻ=K��v����D�G�;� �=�>z[�>�ڎ<-��A4���==T�>��˽�!>-�w=�Z%?N�J?M?�Y&>O.?�s>����>{��>���>,�h>&�V?�0=?ŹT?$ �<��Z��-��k ���̽��=.c�=|	>Ò�=�¨=m���b��	��<��=�,>��#�S1{�Ƞ�e.+>.�>o,?D�>v�?���2.���N��Y:�3��=�q�<���><Y>�k�>�=�>��=��>��k>�x����ԾD��>dk4>��q���H�?��>��i>a�=�k0?�f>�D�Jl��+��>��>^@>:B�>~��>���=���>q��<^��B��`�u�哿�&��-��=dZi>gQ��P���'=�������Q�==$�>��>C2Y���>���	��=�P�>��p>m#z=܂�>,r�=:6ǽH:��|�n=ٯ��$�=�M���i���;X���s��ջd��?�=�gw=�5����?�0"?d�>X)6=��ɼ{"¾�� ��}W=H� ?k�?�(�=Q#?>��`�F�������+=:l�>o*@?F�p>�r������I��ƥ���Υ>��?kE�=�p�=�Z��u����>���>|Q?R�>�L�=��?�-�~�6Ĳ�k�?>��W>w����?e}?7�[�xR>�rþIx$�p���W^$>­=E-��z��=ܐ�GE����b>g{ʾ����M�D>���>��?��"=5x>����C�����?J�=�er=�q>��c=/�@�l���Ǿr�ҽ�2>*ӹ:���塒>Q,�>��>r��>��>?���>�	?T�a=D�I>z3�=��v>ő>ُ�>C��>���>��|�Ƽ>p��<��>pAؽ.t����ɽ�:@��Z>���>y��>�D�������=,�=
�������km�%L��~G��<>~�> 3�>~
?m�V�Y�~>��]>�dX�7���\>#1l=��M��Ѭ�&×>�Ǽ8]�>�u/?�.�=�$���ξ��羪�������8?\>?�޽�A��]l>*��1|l>m}�>����
��K�5~���$��}~U���>�{>��=�?z>��l?(?��?C��sa&�k�b�z9��u�W���R?<_�>�R>�m��R	�5�d�P8d�?�!���r��@Y+=�S�=�->.�r>��>�F�=��6������'���>���=u�Z>�j�>5�?���=Mm�?˾O��A_D?W7Q���۾�A.�%:ɾ/�1�S>���=�ǀ<��+?cƁ��:}��s���`N����>���?"W�?�T?�8t��ƽ�w<>�)>$�=��Լ�����9QF��!>���=����5�Z��Dɽ>ba>��>!d�;z����O�4\�	 ��·e���˾�l��׾����V��� �ǇԾ6h���?ؾ ��t���=�������Gi3�"L������F�?�I�?��>�8?>�vD�S�'�Ʉ7��B>L7��o����<�);�W*ľ�q־����\��R�+������>�7Ɲ>�y�z�����o���/��J�=��>t|+?;ž�i�����
V�=��D>�9y��l �j�z�e��[�˽QP?}�.?ε�`�V��>�y?�%�>�lc>� ���y*�>�`-?p�0?�P#�1����{�αټؖ�?��?��.?ʎ��g��b��\�=���>�f?1+�>i�f��E��,/>��??&[�>��Q�b�x�_��/��>�3?c��E�>���>�I�>C�ƾO%Ⱦ��(�E�ʾ��x=��>��]=B#��F�a���&9<��>݄>ZV+�'HϾ���>h'��|N�)G��{���#���<�8?�7�`�>��f>0�>�*�!���쉿����N?p�?�dQ?O�8?3��������n�=�>xs�>6��=2\�ik�>$�>-!�JSq����@\?�N�?�c�?"[?�El�(iܿ4��W���O����Ѯ;2==��=�@��m=�P�=e(Y=@.H=�=�v>e5�>8~>e�=b�<}ٕ=����Y(�Z���m⊿5@L��u�����%�������E����@P��t#��\��>S=��0���R����H=��s��$o�^?,�/?/��>�@>��潢�޾��=0p0=�$̾��9ﾃ,
�1�$����a=~�b������ɽ2'��4?��$=:��+i�>f�^���_����>�Iǻ'�<��=ڽ^=1>cx;>8�	�_��=d�X>wS�~Nc=C��={z�N*��_G�!Zx�7��=W�U?}�"��l-���O�0:8�P���`�>ʅ?$��:�6��l���:���>��@�B�g�^��	�>��>e�>OO�џa�vm��=�ah�=��<��Y>(��=n�=��{��)`����;�M?��Ⱦy�\>�!Q;l�(?_��?dZ�>3�a>m��>7�>t��=Y>K�_'�>3+��9�T?�j�>6�?�eY?Gճ=I+��eA����=e���m��=�^
=��J=����6A��/>*�+>�S�M�N>	1�=�Q�����^=w�≯�>�"?r��>�L�>�lF����z��E����?�>�+�=N.A>�>����Ye>�A�>ޟ�=�nW>,-_�K����x?b��>!����O��L��<��=��>c�d?o�>K�A������ߺ=q#�=��>!��>��N?���=���>8�=��ҟ�`�K�*nR�k���:1t��ԁ������뽗��=Ow\��>A�W>k9>Y��>>�6=�iC=�S��h��ѿ>��4>1�(>*�O>��=Ws0=���=��=#A���S�o����	<�`s<)�(��XȽ�C�D�=�F�=<���w��>��?�6��&��������ᾨ�0�;Y�>1�>�:s>1��>{���AN���r9�$b@�!|	?eI?T��>��j�`���
����J��zS&?�?��~=Ȋ�>m�׾h�����=���>�'H?�(>�M���<�6�m�1E>�H��>��=NyQ���?�#|?�;��et�:2��^c���_�0�#>���ޮ��ev�T�ƾ,���}��˛���]	��C�>��>��?j0B���V>Ĝ��+١���l�( ���=��\>���>e�<�h��ԾYv���žAҴ=�[G�v�����g>��>B"?O3?"�H?��?��!?�~�J�>_Yͻ ұ�|d�>'~(?���>}��>�C�=M&>^���b����D�c�\�c~!>J}�<]!= ��<�V�	O��M͌=C��>�Y�=��X��N6u=.p	�y�ȼ�7�;J����=���>��(?��y�&�����>�o�<�nz>%�>�'6��r,�pU���>Y�!>��>�?u�>h/<����)����վa���R�'?��L?�>ն����ͽ���p�=�\J>9=�A���g������ζ���B��>b"�="��>�L>o�j?c�B?c�(?᫥����A'm���7��q[=.M��[��>��>�ڗ=��꾧K7��/m�"NS��18��CV�C4��� =Et>ٕ$>��>/5x=F� >YJ��������ɽ���<()Y����>`��>�?r�E>D��=�$��!+�� Q?���`���	��l߾�.���ѽ��%>� ƺ1R?�ޔ��叿a�������A>5p�?�F�?Or)?ޕ����U�ey�=ZX ?�>�yH���ڻ�d�/�U��5�>�O>ª���ߘ�f3���T���>,s=@a����9�=�̿zj��o��=�]7�'"!�"|o�hs,�%8�A4����;��������*�=q���Ͼ$��"W��q�?a��?^�,>�e���X��pE��a����.>Ok=d�^=l��3�`���A<���+��%����������(�D;>�-��Z���@_��`�ޘS�ȧa>��M?t
���]ᾴ ž�Ի��"�,S�>�Z!�ǩ��^�7��=��?jc0?�о���*���>��?��>@�>���������>_=)?d�O?�<�<wf�y`���~B��p�?��?�p? j�=�A�����N>��>3�>^?��� �
���>{�?��	?�ɧ>듀�,�I��d#�Kl	?�2�>�B��=F��>ߟ�>�Н�2��$��"����">�~�>uV��=��S|���v��cS<�'K>&ր>�m�m���\x�>�	�(� 2#�1�������5<���>�G��$�_>Q�>˱<Q�	�^/���v����J�k!B?B�?RdW?�B-?��e��;$�8�<�ϔ>�Ӧ>c��=��\��>���>U<ξF�g����f?�V�?���?�mR?�R�N�п�.����վ�˾w�*>��=gf\>!a˽V�>�=�mb���;��R>�r�>��>��>��a>�L#>�Q�=c~��� +��ٸ��ҝ���8��?����]�;; ��>]�,��|,Ծ�\��`nC�;n�$N��'��T)�\BF��C�u�=x�&?��*?g�!>LH(>M_>�>n�DB���O~���޾z��A\	�����8��ԕ��v<�"��TǛ��MU��a�ܭ�>�7J=��T>�O?�J>��W>!~�>K�q�|���	>�Fv>ķ1=�Z�S��=u�>O)>>4`>��>��	>ń|�<�`���*�-k�m�}�LY<?'��c+þD��ri��4
��IC>=!?��J>A �GwT�1�k��=�>_彽Cx�,^�'\>�A�>c��>��=WW���A��6���"o��Ҏ>mB�>Ϧn>�><���q#'>��<ύ�>+Ⱦ*��>�i�>��?ǐ�?8>?�*�=Q׿>8.�>�>k�[��>���=2m�=~�?A?��?�e?�O~=����H8�r�޽ `���v�T�ۼh"_=�A�|t�<8��#�B=d�@=)Q��%�g>��>�ۢ����Ơ��7�>a�1?(��>���>���xH�w�$�Ɋ���>7e5>Ϲ>�VE>N:>GFr>�2�>Y�>�\@>�¾P�r?�C�>�\��c�~��U0>��7>�Qw���W?�L�>�����L"=t�t>"ص=��?W�>�J%?��>�ӂ>:P�<�B��ῊA�m�F��ʼ�`d̽�]�p�¾w����v�8D�υd>l��=�H>RE>c/>�>Ǥ9���>څ�>�Fa>��=&��=�쓽�V�<^���a���+�>�;t���꘽P���A���hG;�B����%���ｱh�����>��?�!��<��ټ1�B����@�>{?�p�=ɐ�>ǋ�=�x&��F�X����>�V?�&$?��?�!q=k���pq̾\%^�g�>�?^�B=aӄ>����r>�t�I>;j�>�D?���>�
-=iG������4���>&�:�;ž�l�?��?����E�=*Sp�G��s����?[���D�7�X��� �$�řA���V��Nu�Aᦾ_K;D�>�߶?[.�=�=&�� W��+du�����+>�OK>�?�0>����X���l�F�>]I�=!wt>�r1>=�>�> ?�:�>c�?��>rO�> �Z�8�n><�=(��>a�>��>��>G�>�>��>��c<����<ͽ	��Q���"U��=��H=y�>���=���>=�>��J=���4�N���=D�~�Y��=/>�b����<b�?��?5I����i��41>*���s�+=�Z>�����Q7�#n|>��=rV�<�N�>�?9�,>��~�Fw��
�[�w��
QC���4?O�G?��q��4�'0>�""��H�=��>�����=��b�eP��e5��u����>@��:9>�j>B|?��A?�Q"?�>�j-���s��*�����]d����>̛�>�=�=} Ծ��5��Qp�"�]��b/�:�O���M�f�<��=�W">fC=>f�=�>~�<�����ҽY�)��3��z�>��>�?�\[>n�=eS�����f�@?���V
�����U�ܾ{;��r��=�9>'���E^? �yI}����?<����>%/�?�<�?�^?ױD�h�޽�f>�?>��=�e�;@�/��6��6J<���#>�z�=��T���q���� O>6o>\���Reľ�O�N����޿�M��6.�.�ݾ�ɶ��샾U 9�h�3�w�i�r=�!4��z��A+=�X	>'m�8���1��\+��	��W?CZ?�a6>脑>�R�m�޾����e�=~��<��<D��S=#�� �������½4�߷�����F������>g�_�𙎿�xt��t&�H2�JD>��.?Ҽ¾�
��Wx�!�w=T.>�;= ������
��nS?�6?T��i��C𽨜>�?�w�>!#>���ׁڽ�Ғ>Ѐ,?(,?1n�h��������������?�H�?ǘ1?�-&>���A�Ӓ>���>�J�>��?�!��M0���Р�>���>�n��<8��X�E����"?��&?��}��=*��>�8�<.7]�&������	þ"��;{O>����������/����<I�=��)>�k������>Ď羹*O�2F�*�	��/��X[<-�?+2�Ç>��m>>�)��?��O����[��mM?�9�?*�O?�>:?s�ﾵ��(�����=�%�>�5�>Lm�=k��S�>��>K�侯Gr����H?�9�?�F�?�.Y?��k����9�� ���/[;��;�&�=q	&>����G�F�ի�<��7����4>+��>e�7>�`>St�>�>�Wf=����{.�~���A��
E���ʅ&�U먾G��}Y�NrϾ�4���~��9�Z������>����0��~���#��"�=b��>��>SИ>�=->�GJ>��ľ�[�7{A�2������gh��6��U�t�Hz¾����7��2���*���s�>�25���o�p�>�<o��=��x>�A�=1(�==ǳ>6#�=�G>ݩ�>�ݾ>O�<>C	>#_{>�2>Oc>W��{��������2���`�~?�>�����μ��d�*��յ<�ٞ>E4X>�G�ZL��n�>��>6�;̘��P)���?>L��>�Q>���=%*���]�eq5�����A�=A��>E��=]�|>�W��aUڽ��a>M�>i㲾�?*e�>�;?�c?�h)?3M�(��=��>!�$���l�>��>2cT>���>�fC?��/?��>���=��c�������=��[��~��<�[�<�C �X/�5�I�2�<8n>���=��=�~�=�Zڽ�����<g@�>r"?��>�5�>q�@�7���Z��=Y�>��Q���?_V�>-͝<��>5?��%>���=����O�ؾ��>C�F>ic��[����d��>�/<"LJ?'�6?�炾�㦽f�5>h+>��>���>�]�>Е�>�nJ>V9=i��l��=T�np�����@_�P��X���?6ɾ�W��;x�U&>�~�%o�<)�=ʑ>@�>���>O�>��>�q>�y=�fx>G?y�t����r<;==97W����܎��ii0��#ҽ	�=S�=���ڑ	��K=|M,=j�>h?��ɾϢ8�2�B��׾�����?+%?���>z��>d�>꾥���־��X��/�>��?�6�>6B�(:?=�ޙ�����] ?�(?������>�6�����[�ڣ�>.k1?�B�>� ���$�-Bv�������>}b>��|���?��r?���!��=�$��LZ�=�4���>_��N��	�>U/)��}���%�]����=Y�%>冪>�z�?>a��V����-=�Ԯ��.�hX�=���>�B=�lc?k��>�ˈ�R~C��,��>B�	���HQ�r��=,�>�z�>�+?�?G�q?�L�>JjO?cϽ%�q>��Y=�	�~$>ȅ%?�p?߹�>��"��>��ҽ;X�r����`�G����5�=)ڄ����<^^>��"�#�=�_=��O��=�ų�bR���w-�+7�W=*>��o�>f�?$1����Y>2Y��dt�ẝ>��Y>i��d3�=:b5>����^,>]s?~��>j��xx��+���ł�\"A��=?�Z3?e3�=#菾�J,>Q��0p�>:r9=�*���O�� ��~�K�t����>��>f{�"��>-�|?��a?��"?�DS=���u�*�p.�~
�=ٱ2>*?���>�3X>�ȉ�l�O�����L�W���,>r�5� �<��w���j=�ܥ>��=���=N�Q�0��+����q��v��ͤ>�X?�3?�I�>>2ᔾT;���	@?�c�����K��>3�7���=��Y=@�c�֌����?^�/��G���K��2�2���>t�?J7�?�^?�@���J����|��4??O�q�	���>�	�hu �v3�<�I�=P��K������>C#��k��>b�<��e�7]��u�f>����`�T��8v��.t�#��'�!�����[�M�ɴ���W�wj���H� Ş��Iǽ�V��]G��}T?�?�� ����f�?82�?�ڼ{>�[:�ZP\����>q8g�Āw>�RL��N��¾kR.��ؾ�`߾�j��j�?���$���>�S��[���y�[%���;���A>��-?�x���(���Vnv=2@&>_��<S��e݋�񙿢���U?��6?͂����Io�(�>��?$m�>4r&>V���
D��(�> �0?�+?Ҿ�fÎ������T��J�?�Ϳ?>}'?5X*=��߾��;H,�=�8?:�>`�w>~F&�ڠ�5��1��>}�?��>��4�.�U��4���=�=?��c�=uǚ>�` >����]X�r4r�EXc��EJ�G��=�t�=��A2��V0нgMU=�P>�O;�A�23�����>���YN��pA��@��[$�}u�<M:�>���D	>I{Z>J�>E�(�p���%��n��K?K��?P�N?E4?��U�(����qD=ʕ>�h�>�t�=���g�>���>1#龭�r�����*?T��?���?̌Z?�o��?�p��v;�����=o�=��E>ǹܽf��=d�4=�ӻ�ir<��=��>I=>>rR>T�k>�]�=��=Y}����!����U���)?�>���(L�Mq�s�_�鿔�Ԭ������Z+�/�	��0���E�Q�C�D���m�=�?? {S>��>�>F �=ٚ�����C >�3ؾr1P���f��	���-þ�����۽����=�����P���@?f���V?��)?ahŽ��p>rL�>��ǽ��{��!�>!>c6=QK>�J>sQ�<N��>d��>���>n-�=ȑs��/\���0�;�~��)x>?`wd���ӾW��=
��þxȇ=A�
?�V�>�K��C��q:�>��>]��2TF�ݡZ�w��=��>�)f>�@>�d}���4�}w���5���>�]S>��T�ة�<]���)��p4D>�t�>�0a�y�{>"��=/	?��a?�?G��ߜ�>�>�p��6}�=~Qc>l�=���>O��>J.?e��>��?�u�=��t���!���=���@o�<�t��<��Z��E�����#��<U�*>3�<Q��<���=*x��b铻;7=+7�>V ?w��>��?��z1�5������٘�=Kvh>�=]�=� >�i�>�� ?h=�>Ș�>R��T��L�>|@�>d�5�e�	&�:b>���>DY?�e!?Ġ�<c¾J������)�=*$�>
�2?�_�>b��:L6��������;A����'W��߼Nc�=�rh��I���|�_�=��=��o���f��,�=7׀=*>��ܼK�|=~��>[��=|��=S�;>��{\�?�!<)Xҽ..�H�7��T�����:V=�༔��;���=N��瞒=��=G�?J�?������	0�����!�Ӿ�: ?�'*?�-�> ��>�y�<���=����?�= ?KQ?>-�=b�6����C`F�`��d�?� ?�u�<g�R>>����� ->>,�>�?��<<���])��$r������?�1�=w��Qq�?B�\?��Ӿc�>4q��s�E�P�Q��=�g¾ƕ� �>r��8�y���b�߾*{����>C8�>1��?i�ξNR�=��������-��о^�_���>l�P?���=J����2���.+������5
>b�뽓qC>�i	>�h�>T��>��>�??��?�P?Ӥr�u�>\�=Y�>���>O��>���>Cv?��>j�'>yI�$C9>�;%�"����h%�B��<q=(�z=6BG=��<��>�(Y��3e��E�=�2�L>�(�9=s�=ڹ=;!�<�B==���> �
?-\2��m��F����۽j�=S�=��>�j���&�,ҙ�����gk�=�"?�`?E��=�7��&����Ѿȋ=F;�>I�?qU�>�ra��o��Vd�=���g�>��>f�,��߁�
!¾eP�5rh��I>�X�=��Ƚ�
u>�̋?�y?U��>�{>(ě��ᾤ_�'�O��>�,?�Q�>���>�0�P'y�JՖ�d+2�rg�w�>D=���
��BH>�@=B�>(�/>�'>m"���GD��˽�^r�K�>YzX>�ߞ>:�?�S%>��=%�������UA?P!�����0)>���l����U>�C>(ݔ>�O?ҙ��_�`�Ex��#�$��>밨?+W�?rf?�������=?�>>M����߽E/�:^�;7K->��4>T�p=r���I�#��sm�>kTa>X�=>��Ȇ����q��"ʿQf�Y~�( ־���|&��	�	��a��V�Ҿ���mFB���������|��!a���#��;��g5�������?C|�?�����9�>�Wq�9�L�r/���k�>0���1������+�_�޿���ӽ)-��e	�$���b˾��3���>9��
铿���ʀ����Am�=t=Z?�x��J���@龠VT>/���b��>�6�qS������^U>�?u�e?�������Z��3�>f�'?�p�=N��>�$���'�>u��?:i?T��>[vh���{��eϾ��?�r�?�>�&��97�P���q>"��>�$ʽ���>�\,���O��-�>Z�?�?-?��=?be��
�}��T���f�>n��=f��K?N>��>�i�>����x��\=X���O>(�>h�=�:!��D��1ý�$�=>��=��>��{����9�>c8��N��H�O�������<\�?�h�,�>eoi>�>N
(�_猿Yt)���L?��?�TS?w8?�����������h�=��>�s�>���=(9�q �>A�>gO��tr�by�5O?�?I��?<WZ?Rm��Y�
s��@ܾ!���U�=$G/=��Q>請��=1½����E<v a>�q�>���<�S�>�P> G>�@9>����!�y��6{����B��������5��p���A��	��y�����Az�H���e½�:C��8]�-���_?��� �e�>Q.�>.,�>��=c��=�;��� ���D�<�%��굾������-��K�ȾL�����k��g���0������ ��>4o�/�>�S�>�V�=�	�>�.?�V>+�%>��T��>��>	�>�ǩ>�;�>Tk�>��>��=��=W^����E���$����-۵��D?�'5��s������N�+�����)=$�>P��C8@�5P������2�>�����s��ٜ�a/a=m�� �">�W�=�����9�<�|<��3=H��=gr�>��K�:=�#M��=�<��U�&��>��8�>���>�d�>c�8?��X?�b>�>%?B�q>�P�>>��=��1�z��>LNX>�q�>!?rK?�z?=^8���h�=��=�૾|����U���>�/�`�Q>�i�=m�(�%b>u������= }=9�Z=W2����^�TM�>0B?�?��>�Н<���v;�f��we>\��=�u�>��G>�m�>uE�>�&?;T?�҇>�:��G=���>�->���^r�|�bD��#�y"?H^�>#��{v��4u<��ǽ�y�=c_?d�,?�7?�|�=�)�ſ�`d�y�'�n�9������߽w�>���r��oQ��c׽�nQ��o�;�4> U>o�f=�RR>FL>��>\>��>WJ>o�=�N�=�H��6���N�i�<:'�<�݇=�w<B�^����I���pߢ<U�g��0w��Z��o�ӌ?��)??r>T:�=F���\ؾ�#߾��D>���>�o�>�>���=����Y�4�G����>K�=?�It?F�-?�U�����<�
>�>�?'�K>�0<S^��p0'�qЯ�kn�>oVA?��?�K����^�����/���to>���=�rd��?HB?��m������m[�q���<��>���,%>��G�po���!��_��"�1�(1h���=+��>�(�?OWe����>���.[�����b;������*��!4?59>~8�XQ�ڷ�t��S�ؽ"������>^�X>���>F��>w�>�/�>�~�>���>��=���>�l����>��Y>�K?}
D>2�>W��>-m�>}l<=�$�<�@6�5�O�����l	�a�>R�=�)�= �=���=��o=ת>{������2Y�=��&=���;���=�<`=^L�='�?���>�w=n�!>����I>��>@�f=�]>� ��|��AP>�=:�>A�?a�>9�J=(b��z������3��<iN$?e+�>�X�>��y��>yپY��<p�=�*>��=��׾s+������=;�%>^��>t��=�Km>�y?<?;m!?�W���*�ݼs��%���w�t��C�>�z�>A��=�ܾ/�3��<l�=�\��:/��S�D{D�i�<��=�>��>>��=�">��=�Ɨ�|�ؽ9к�哼�W�>�=�> Y	?�V>��g=de��ڱ����B?�cv��f�s��t����	v����=�w�=�|�93?CT�>m��1��9�G�u��>���?�W�?��k?�k��ɞ
��oE>�I>S�> ��<�P�b��h과��>�a�=�-x��,����;D�>RF'>�Ƚq����۽�_�c���ܿ�����9��,D9�L��U�侢��T���^�?��.��;}���]�t�����R���-X���X��޾/�����?{�?j�&>ણ�������a�4�8>*�־h��E.Ѿ$�
�_վ���D���� ��G�6�:�X,���>f �A���8j�����v�<�~i=�	?�EӾ,޾���.�=xߝ>�E>���t�-��H����9?uE-?�6�V��[)�<k�a>��,?�?�e�<
�����P�[�>��N?��Q?�8>�o���
��D ̽>�?)�?I�0?���U���Ǌ�f"�=��?�{?��>��̾����Kw���"?w|w?ϭ$?���h�4����>�?%�p��j�=���>ȷ�>��l�� 1���9>�5��#=�m7>���b�$>ǽ���U�����U)>IR�>d骾��ؽ��>*e�<6O�ǾH��������<��?���>�i>NZ>@�(�2㌿>ى�ө�uL?�q�?�S?U 8?�%���9�5ݧ�~��=���>��>'�=Z��tޞ>���>����)r�o�W?�?3��?�&Z?u[m�0Gӿ�����������=%�=�>>��޽�ɭ=�K=hɘ��[=���>P��>o>j;x>g�T>�<>��.>l�����#��ʤ�1ْ��[B�� �����vg��{	��y�����ȴ���$���<����Г�w�G�s��ZU>�<���R2�U��>$K�>N]�>��¼�@ս͔P<��������*��R?� ��R�J�,�)�A"Z�����᤾����B�*I�>h�
>��>��>�２x3>7��>[)�>��[=v߸=�b]>��%>6��="�t��H�>̭�=�v�>�'�>Gi��%{k�3/l��T8��Ҿ�/���X?�tE�1S�(㾃I�$�k�eE>5NN��HɽO�c�3�������>����c��Z�PƸ=1�<[��>���>�0�����-�P�"��;�@#>���<H�A>Ϧ����$>H���׆>>�Ŧ���>��x>�>�j�>؊?#�=�?]�F>f�>�wϽ��?63\�'$�=�9c?Q�
?��H?:1?y=ν��|��"�=��޽]�T�Q�=���.��۽��_�.��E�.>pHҽ���>$&<:�ͽ��5���ڽw��>��u?�6�>��>,��=Ag����H�Չ����>�h>?I�>k8�>�c�>�6? dX?_ڿ�P��>R9�=���]�>�ҳ>X�g��G���'��G5>��>��,?r�?�g����V����������k	>���=��8?���>���>t��=���jӿ{$�Q�!� 킽�L��`�;��<�9�M�D���-�`����<�\>T�>Q�p>�E>(�>R3>dJ�>7G>�܄=M�=�Ǥ;L;S�E���M=m����F<�1Q�����ļ ���LꋽP�I�_?�5n�:�ټ���>�r1?$�}=��E�
;+���`��)>��?�d�>���>2^>��t��&�y��Ȓ<+�	?��\?]R?s�|�q,ݽ����G�=��>}-?<�>��X�9���4վ��O=
��>0?�)�>������Y���q��A��Eq>��Լ%����?.u?7�	�K ���*�7�@�����%$>pK����=ӏ��3.������a(�j�H�#��=���>�:�?�2��uWI>%5�����S��lB�	�M<gs���>K��>ՠ�=�֜���D���˾+_ʾw/�=(�l=�d�=湪>g?a�?V1?���>��!?^U�u�>���=�?Ѱ�>T"?���>=�>�Z�>�N>4|>�\4=$/���N�'�U=��4�d�5=�4>� �=6gC<���:Z&=δ�<�ƽ��Z=�S�<�Fy=�O�<E�2=V�2=�	�=��>��>/��=^;1>�"~�vX|��C��$k�=�N>̡g=�?��1ּ�e���f^>�d�>���>��D>��r�������*�7����8?�z,?b��=/R�����g_�������>o�P>���=?���{��Ꮍ�K5=�Ĉ>��Z>��#>ݏB>�{?UpG?�)?�)��n*#��l��|9�� ộ'��t�>r~�>\�E=�R0�h\n�]�T���#�� �:y�B��`=c�>���=�*>i�>���=s�;�����׽���<(g��%b�>�z�>�?&�/>1=v����*��5?y�p�{�޾>�"�cŤ�e�ݼI|Q>�)O>�^�����>���x�c������8�+_�>@�?߉�?��e?�Sɽ�B���>n��>���=�@�<?b�7�>=F��<��/>2>�����r���R>a�!>�������E����!��6���X��:ƾ�����o�D�v��1M��7��oξ����Ɂ���p��mw��!y��8ؾZ8羡"{�ſ�,Y��?�?��?}T��+<�c7�8���"�ōe>�
�����#���,��|��)>%P����,���I�1f��Y��r7>�x��Ϩ����8S�3�+>"OX�Dm?�������U�����\��N��>26�����M��ĕ��a?�F?'����i�z��,�>{�9?$3�>>}>F��_�m�-/�>�W=?���>A�<�3���Z����Fy�?v�?	=?��<6�:�������>�K[?F�>��Y=;Zs��� ���7;�`�>	4�>W:?�߾o�o����@�=�Z$?��X��	=��?�?xAn�SƲ���>��v�(B&�$|�>+����=��k#���P��ȣ�=UC�>t|�>e�a�9�n+�>�}�A�J�#ZF�C��U��{�<.?��V�>_�`>M�>��(�D�W ����
��:K?ձ?��S?�Q8?�F��(`i����=?1�>ᮨ>���=���K��>?��>���P�o���%?��?�@�?��X?�^m��3߿9㣿AH����̾`�>?E<?��=h�c�:�?=/�3�r���u��me=�>[>���=M�e>�b>CC>����1�*��"���ș�?-9���J�1==�:�6����Q���sg.�<�U�ᣫ�dY���Bq\�LVG�-/:����;�<��9�=ғm?H�?Lu�>?��>���>%Gž�r��1�">���Uۃ�n#��T#��������	}��4깡;�����,7?nA�=�"�>��?�ʥ<G�n>t�y>�>�=_��=�>�>S�= 8>��=�\=F�>�Ċ>�x�>��ɽXb����J���C�:d��jϾ��~?��~�+�뼀lþ�V��P���	���=�q�<�G���{�������>��\��&Z���<4&�=dǌ>��	>\h�1�<b+[�A��m-��Mw��~@>��V=��=S\�`��=���:Q�>G���"<)>k�>~JW?��2?�e�?O��� ?�
y�g �>�i>`����-�=My=�eS?I�?~�j?��g?h����-��~���н�q�DS�Rh%=��Q>�#���Kn�����7!]����<>K`=�.��P^=�R�<]k�>�
<?~�>l��>B+)�EWR���7��z�cL.>�����	?L.�=��K?���>�dE>�S�<�5f�]m��z�<�)�>p�>�X�t6�����<��>U�>�9�>�{!?�&:>%_��>돪�0��>�^=�B�>߁�>���>��,���N�ٿ����M-��Hݽ��T�+��#i������T�{���z���
�=*��>��>ǩ�>���==!>LcH>���>��$>�U�=N�=pO����>7݅<W��=Hq<��<>��=ި��Ȅ.��P˽�2N��Aǽz" ��k��P��?ϗ?s#���X�r����HF����>3��>��?N��>d�P=���::�Lc*��Y>��o�>�,Z?g�>�[B���=31=D9T=�\�>g�>Z{�=�����5�3���J�>��>��? >>/%缡�X���k�����Ǉ>u-�<WK;���?��a?��Q��r==�B �:�K��	��8�v>_�TK�<�u�<JQ-�Ә޾���t����D����G>�a??_�%����:,r�M3��잿Z��+� �Y�m��?�v�Z�T>�B�=����[�A�(=",^���=�{�=R?��?A�>t�v?tp1? ��>A#վi�?7�/>l�>���>D�?ذ?��?�M�>���>'l�<���=I��d%���6�<�?N=��;=���>v�S>׾�<З��#�>�-1<y`���4 ��Sv<�H=�zK��=T;2=i�=Tz?��?m��=�!��Ϛ>������y5��7�=��/>d���4e^>�N�>��[>-�?���=�v���?�V[����%!�b�_?��<?�H�=V����!>� �;Ν����=C�>5ܢ==�$�͏���d�s+λ �>��"�#��>�s>�LU?�/?�'?|�����}�v�S��u�{���߼b��>���=�ª>q�ݾ�4Ѿ3�R�dV�m�,������7�	F�<(��=��r>j$!>���=/��=���<p}�;���
<
>� �X0�>�r�>�B�>��>�9�=�%��4��=I?،���z�K���wҾ��q�?->D�E>i�߽�?���x��������&��r�>ެ�?F��?u�a?W�K���1�X>�a>�>�	�<��f��%��\i���I>�^�=\Qa�"H��:B>���\>l�>1 �����;&�K�_��`/��v^ƾ�0��޾ID[�+��9z�;�"@�I���B���3��Bꊾ����^���@g��+�꾑����c�a��?�~�?�)�)i����P�7B���ҾZ�>}�����<�qϾ%���f�<:��������ξ��C�e�&��6F��}�>.X�����|��(��˞��>>�>/?8�ž|c��<���kc= �%>h��<J�rF�������
��U?_�9?�o� ����_��>>�?��>�/$>�e��l��dG�>{�3?��,?�߼�ڎ�������m~�?R�?<S?qN��7�0��N��	�X�%��>Ӝ�>|��>Fe�몾��^�t��>��#?	"?�� �n�c����<?zr?&W�?̼=��?M��>\�(��&���=(p��.�=�T:>�<U��<o����]5�{�+>�\*>w>�♼ԩ��"L�>�Y꾖EN�NH�j�k��l�<e�?O��f>f�h>->bX(�����ى���%"M?Nu�?��S?��7?����"u���B��=�
�>�%�>y��=��a۞>Vq�>'���Dr���kz?��?%g�?�Z?�m�i��#"ÿ2վd� ���'=3��~>>?�v�<h�=㽣=w���6�	��<�R�>���><��>���>��B>{[>;}����N���
��32�"�����G����mԾ:[����25�������h�ǽ߾���=�,��b����~ �\�O�Mi�>�\�>���>SF-�4��=��o��\����$>O������oY�y���Sw���e�Bpt�J{�
�e����X��H5?#%�L:�>�D�>���X�>+��>ۤ	=�'�>v/��&N���>0��>*$}=d�<0�>��g>Qܠ>�v����9;*���L��ϛ�=۩X?r�N�,m���M��H�ξA���<�����=+�?���`���u1�>K�0��»"@B�����UW!�ē�>M�Ƚ;F��5N�<%S���X`>��;�65>7s=�n>��P�==�=�聾+A�=��ѽ3C�>�׻>*C?���?ͱ�?6(>�"f?PH �qka>�\�>�k.>��<��$��k�>�'�?G��?v\{?�u��p��4	�*8��1K��?>��˽�d�>��<i�=ꤔ�Z����<h�=Ԍ	�ê��8�<h��=ʖ<>pxy>7mv?��	?���>�X�>q�L��O���־Gn�=/$�=*�G?�4�>@p@?Y+?g�N?�x�;�E>����M���^�>��>�z#�b�_���!��W6=�JZ>��>�?Cp`�E�h�<
�=)>ӱ�>̗�>�:�>�2�>��>��	�y��Hlӿ�$��!�J`���;_�<���M�O�7r�-�����0��<Ã\>`�>��p>)E>=�>�83>�Q�>�HG>�Є=��=� �;�/;��E���M=���SG<d�P�Ǵ��AƼ)���~���I���>�N:��3ټ8e?��?��M�;�=M�L����M��[й>�N�>�-�>wH�>(��d�ž��O�v*� ���M��>L63?���>��R��X�8�I=߯�=��/>�K�>�V�/]�Ӡ�)D��Pν[~�>���>Gّ>T��=�P`�?q��H%�9+�>�JL���^�5�?��5?�׼1�#����e�i�#������>�O�=:��;���	㙾�ԭ���f���aX��N�>n��> B�?;>ʾ� �=����}R��u�*�ƾ�j.������>��*>u�>�W��_����g�I#D�Kݽ����9�=���>��>DO?��H?ޫ�>��?V/�?��%=iO�>�>�R?�9�>��>(@�>8�>�W�=���� ���^���;�"���q|<�_>���>�w��*�=+��=�]�<��|��|�=b�ȹ�*0���>��=DG�=.>g�?] �>�쮽������6P5�K#�=}nH�z�@>}F�#���m>��u>8]>�,>[�>/[3�l�R�����ݾ8����`?�e?s-i>��,����=u�ﾱ��O4�>���>RK
��|���X���WL�|���>�V�T�>�Z>G�x?�0@?�q$?�dս��,���v���'�2K�5�;`��>��>� �=��ɾ�(�õo�+9[�(T1���+�)C�q �<z >w>��7>��=~O>X�|=;R��I>���W�<Wu6�ʥ�>@;�> ]
?�	L>��=�D��r,���+?��P�����DV�1�Z�y�8��=f�;�� 1'?,�ۼ͊�����#h��+�?��?��?�<y?��0��@�@��=o�>�՞>�$=��$�@�G���=��(=�j����D�<|D��<G>f�x>�݁���;v!�*V�XϿv�;U��]�6��xZӾ�������D��k֘������эȾ�"ܽ���lW&<����L��C��.|�?֫�?��Ǿ���>,�8����� �Ǝ>����p�~N��}��I����K�n����E���i���0��'8�HK�>�@o�E��9Ly���#��[{�zP;>�8+?�ľ�Я��A��d=�D�=�=3�����o��
���Q?+
;?Y��W���s���Q>+�?=�>��(>�����#�x�>67?'�&?���9򏿿���1���YQ�?渼?�v8?�3<���@���
���3�/��>$��>���>����ZqоL���q�>X ?�ɮ>�i �0�h�Y���>=#&?�hR��c>���>��m>yf_�Uܭ���(�����$�;ř">i?�:����YC�6jl���=���>vv>��<��ԙ����>���{
S���A�����#��>���	?��XY�=��r>��>dt1��ڊ��׆�ñ�	,>?�z�?ĊA?]�1?r��$��;n۽L
>�v�>��>719�qֽ�{�>Mp�>�����u����V��>�{�?e��?6�h?
�i�:Gӿ��#��������=%�=��>>��޽�ɭ=b�K=*Ș��Y=�d�>x��>o>L;x>u�T>ۛ<>��.>p�����#��ʤ�1ْ��[B�� ���wg��{	��y�����ȴ���F�������GГ���G�h��U>��M��!����>}��>��=�@�=wE�=m�N�g����.t=��Ҿ���Q퇾qA������ݑ�� ���W��f	�v���aV����	?����~>�v�>�H���>@+�>�]�=�:>�"=N�u=���>�>�a�=��
>���<���>���>vz�`�m��Bk���?�0���·���_?]
4���ļ��3F�� ������>ݭҾ�lb��;��㠿�y�>U�:����{�����=���=��>�H��{���-�=g�i��";���y�r6�>��ѽp�E>!�S�]�4���?='�>��-�Q���.Z>�u?�8?��:?���;�/?hw����>͚�>�ֽl�=&=��5?�.?7?��>�`j������<�'�l�V��Eܽ���=�b1>�@�=�Q���ڽ�!:�>�,<�?k�=[hk<�k|=�m>j���ס�>�/]?�?ur�>G}
>���GP��`��w�\=��>�Q?u?�>/�(?���>X�6?o��;�S�>������,�>O��>�Q��9u�y�G����>�RQ>~�?x)?o��=���<�\'>�]�>�s<5'?S�>k�>��'�l��O�ӿD0$���!��a��W�V;kW<��eK���9mj.��q���<\>/�>C�q>nF>� >�3>�m�>��F>,�=X�=U2�;ם�:��H��K=��BwI<�"L�E⮻B����ʕ���{H�t@�+|��2׼�?Wx?۹�έ�3��������OR���>WH�>�+z>��>���=�������#��mc=쑣>)�Z?���>�t�F(�(j=Q>� E>Sb4>ى�=���5|H�k���8� ��>�r�>�Ȏ>"���S���o��(���>r%r<�/�ba�?�8o?�ж�>�Ǿ�n(�Nu(��.㾾X?"{ȾjVh��Xn>+־`�;��,���Ⱦ��Ⱦ�T�>�@>Rp�?��ƾ>��=g\Q�H����t�':@��k�<|X1?�:�>Wl=�n���.�ʾ�1b>N�9>��>��=�P?���>���>[SY?�X?�d�>�뢾(�&?XY=�"�>�>�6�>��>�q�>�F�>�> ��=��5>���U����<yfм�;Z<Z\�=��~>�9}=���"��=e^�=��b�1���ԗ��|�=V��=tC>���=z��=B��>��?�F=��I=[����$�[:�=-*����}>q��=��9�Ob���;3>��? ̲>�?�� >�𾣝Ľ�����0�tf*?]�-?�>ί�[�������n��c>*�^>��P=\��P�۾��������>�I�>��S>�G[>[G\?� O?��D?��F�<�$�v	k�e�0�<��7K>�>Y=�>�^�>3��Q��j�//F���1��^=�����O=;T>ڝ�<�Ζ>2#�>a=�>fq�:YvĽτ�����]^6��HO>I^�>�%?��1>{B��q��x���I?(A��'Z��C�� XϾ�$���>Q�>>�e�F$?��_{��O���<��2�>O��?o��?��c?g#B�N��NkZ>��W>7#>�X<b�A�e���ٍ�p�6>�C�=~v����|:��Y>�r>E,ǽ#yȾ;�߾�29�D�����K����辑�����)�n(��:����N��`<��Ѿ�q̾�7����;�$�;U��l���E��C��k�?ч�?��q��P���w�n����徽[�>�����r�{���
/��ֱ��~�<��Yӽ�k��3Q�>DN�C�=����>O4`�aK��:!y�)��迼U0>�"1?%˾?C����8\L=��>=A�<u����-���Ҽ���P? 7?>�������ؽ�j!>,
? q�>��>	ԓ�rW��J�>��6?ހ*?2;�����?��� o�<j�?֣�?�U,?�ƽ�n%�V]þ��=��&?Q?��E>�[T�����:���7?��>�"�>`N뾳Us���Y�>�?�I����= b�>���>�޽�q��/�4>+����r=4�<b9������ʂ�������;z#�>*aZ>�~��Y;���>☩�BaD�*C���)�J���<8�?KQ�3�>>���>bR/�A�9�/�����{�!�F���C?Y�?Q2&?W��?N;N�v����ϔ�����{v>�<�>�I�>ni)��>��>�ξ�$��@顾�|'?@�?C��?��?�7Z�(Hӿ���k��������=�%�=��>>��޽�ĭ=��K=�ܘ��6=�݋>���>�o>�8x>e�T>֛<>��.>Ҥ����#��ɤ��ؒ��ZB�� �����yg�V{	��y���6ɴ��ｾ*���ݦ���˓�a�G���R>�
� ���0�p9T?А�>D��>��>��1�Ot��H��������r�DVU��]}�;z���~پ��[>���پ���
/�I	Ӿ`Z�1zP?]��=&ׇ>~�;?���=5϶��N�=�29��	�>�w���Й>�-�>:\{=p�>�z>��Ӻ}���7�k>�*>�׀�Q*y�nn9�Z|��!��5�P?<�ؾml�����5G���֞��IZ��4%?��U>ʣ�`m���J��>z4��h2����i~�=�!�>�u�>fA�=��;\e��8w�������V����>��>���×b�!9-���b=M�>��\����>'��>&�.?��a?\F.?Q����>g�����>9��>��>�z>�e=�_�?Ev`?��?(�?������\�<��;�w�=����ϸ�E-�>8eZ=�I齁F�z��|
=�>�j�==�=��˻�5:�}��!<qa�>�o?C^�>��?�!=>�ܰ�t����Ծl
�>��X�Rٝ>.�>:~�>/��>Tox>�>�,3>_M�U��>��>�W!>S���e���j���H>�����L-???(�>f���r �����/��=��M>20?2x�>��>�ﾋ� �~���Em�%�'����u���4�>�l���ѽ<��=�dؾ��C�e��;9�5>�4X>|�X>�LO�>���>���>6��=���=��>Y>cg㼯Rܼ�+ؽH��'�=��>ս�����ě���'���D�Fgs�*��=�G�*�>�5?�`���d���������$쾜��>����i�>���>��=��]&N�a�[�C��IX�>��/?D�[>V�"�%
Ƽ��A���O�f��>'B�>�R$>���=�紾P8��s����?��>�J?k���1z��.���{���>��A=J�!ַ?)��?,?t����>t��aX�{ձ�\�X�r�F>�.���Z^�|5���7{�N��=]3u=O3�d\��ǫ>\��?�{�@�>�!�;6���MP�C� ��qZ;�&6=J�=��>�?���r���� ���="�g>[�E?l�[>�X�>Q?�"?Qz?h�$?��?�ξ3~�>�Y����O>im�>Z(?,��>�!e>�>��>���=�2�}>=���	=�˽�\�ؽ^�=g8�>�0�=�s���0���|=Mh>U�<E�V=�����\��Z�g��;<T8>.��>[��>�O��C�;䤽��G�c2����(>->^�>�Y��� �<�;���e�#��>��>�sq;_ؐ��j��0v�RCս.�?N�F?r>�>�C��$���T��A�">�	i>�Q==Pꕾ鵾3]z����l;>B�>=^ύ��rz>��W?��>n�>�c��/��f�:���Oo=wL`>�h�=�6�>���=<� �c�3$�d�a�A��eY[>+�[�c��TE�=3�q>�ȉ=�y�=�f>:����=�w���x=>� ��l�=��>Y?ίU>9->F���oQE?Lo������ē�\cþ,�R��="�2>(����F	?)�q�E}��Ȧ�s�A�
��>^��?O�?�SW?RJp����f�@>l\,>��=�ܙ<	� �?~�L��	�=��W=|����<!�l>�<�>�ܺ��:���̾��J��4ο��i��1��4���Q㗾)'�J�����Ľ�w\�b��=�7���Z��/�<��c��s�6`���k��R���=��n�?h`�?�Lv>)��l���+yb��_����>�������P3T�*���A���ϭ���|���}嶾��������I>�o�<XN��������k��c��4�=�^\?|����Ѿ�݄�\��d7�u��>�R��ԣ��Wz�ɰ�>�\?�NQ?����	�=�����=(f?X�>5(�>�����9@>nR?|�3?���>�l��Y���y˾���?y,�?���>�)�=�%#��4������N�=2{1=�i!?�R��;A�/@��d ?��v>���>�z���**8���?=*?`�A�e(�=�m>`�>,��ֺ�]@[�ȧ���L�>γ�>���~2$�-ߡ=t����==�>��=���~�6��P�>��ﾜPP�B� �,[�ɔ.=3<�>�h�=�>!�j>2%>=�!�1ʌ�`����㽺�D?�Ĩ?�@O?8:?AIྒ׾Lս%{9�6�>�A�>�R>�^�Dg�>P�>!�޾�(w������?˒�?^�?�b?�g�"�ut�����x���m�=Q�=�[N>��C���0<��S>�>2�Խ���=��>&U+=8!�>��=�K��ZO>�P��_�%���ÿ7j����R���򾏌پeŶ�X���=���Hݾ�V��s#ž��w���O��"ֽ��������l���5�ͽJ�Z?7��>X��>��>YB��K��g����>��3�����M�h������ׯ���2�+e��UY�8^9��?�	��w>�@<?�#��F�>]d�>2�G� *�>T+7>i�=;�=�0�=Ap�>Ng>�>��=��>�&�=�"t�4lz��z5�k勾l�;�9H?���8c�,+��n��F�����>�V?�=9>R�����_�~��>H�j�)�A�����C��u>F�>�E!>^1���Z�6y���ܽJ}�=ό}>@�=<�1�2O��&K�)�='��>�{�����=-��>kqW?�?ky?�`\�f�P>���/�=-�w>��Z>�T.>@#�=\��>�l�>j��>v��>f!T8r��e��� 0�l�	���#���ϼyU=ox=�.ҽ�K�*�>�U=&�����=q��h{�Rb��j��.��>S9?�'�>��>�ܙ�EF!�"*F�;��~Y�>��m=�̇>|0>d>�Y�=�j�>�;�>ۦ1>��ý���\5�>���>�D+����G���M�<|�E���L?�N?��>�侳a���XB�X�b>p^?��#?a�!>��>ɧ>�0�f�߿�W����P��'�;�<�!�#��nⲽբ>(���j�9͐>0+>�u��2��xf>w���?�>��?i�c>c��=���>1��=B	��tZ�눯;�g�˾�'����=>�5�>�ω>p��4�>)��>7��=�Ln� f�>�&?�b��>��o2
�b ��d۾c�?�-�>]�>aj�>[�a%�no�������=�W?��?��>�թ��9��uύ�K�H�XG�>
��>��2>v�F=@ɾ�ۏ���@Y�>�?'-	?A|\�Y�?���@�Y���Q�>�{�=��U�|ї?�wl?$;���s�=��ݾP/"��_��'��"5�>��,��Ww�p~��G�Y�������c���?[m�?�վ��D>�R�S��4��+8*�D?=���>��>+ψ����a��8┾n�X�ۗ��wn�<z>�,h>ZW�>�6?φW?C�}?�P+?_C?i���ҾP>���<z���D�=E� ?q=?�Dh>x��=���=�r!=��>�?�P����=� �=��M>;M>0޵>O��=/�!��B�=��`>��ѽ*g =��=:�m �դ���D=\��>��?��=���������ƾD�	���>t�>O/4=	~h�1]C�?�p��>���>�l�<�&=Rp��6�[T���諒a?��-?/T�>j��<4>�eؾ!�K��=)'Z>�N߽-V���&.�Mx�n'�;��=̜�Z��
y>;�t?�B?��,?��ڼ����:[�\7-��࿼>벽�Ά>��^>��=$�r����i,d��Q����f1=C�E��>��1�(>�gm>x�">�X�=� >(J�=ꕿ�����cX���盫>2�>\�?{s>�˻���E���?d	����#9��m�#����HN�ݠ>����?��!>q������ DY�H� ?�(�?w��?C;A?�Ə�����c4D>��K>�E�=Ǘ4<!��Q��<j�ƽ��>_1�>+0���>����#=�:>#�'>'��=9��ɡ��Kp|��#ֿ����%��&�ļ��F�.�����Rh��A�Ⱦ����97�܅?>�"�;�f7�-���$ ���U>e������ؖ?~��?ͳ�>�t>��a�����ξTt�>�I��K��	�<?�����j�!�E[��75��z�~����3��8�>$�C�1���3�nQ8�oֽ�mA=��F?uS���Ȉ�،ᾸF'=偱=�v!=�%��V�x����N:�=@K"?h�,?��Ҿ{ϻ��b�^�r>�?r�>[�w>L��U����й>�???^{<��g��Ƀ�EOͽB�?��?��?D���D�I����	���l�>(T?6��>��w�����-]=	�>?�g�>��1=4� �d,�șP���>�Q-?�{Ƚu=Zj�=/$t>̋�������;�T���~>I��>�����)�����D�޻��U>��s>�ʙ�� �����>���'O���I�"8�k���R<k,?���1U>��f>��>>�'�������uV��vVL?��?7Q?��7?p�����쾎:��dg�=�j�>;��>T˲=؆��ʟ>&q�>�����q�����?��?m9�?[?nFl�#�y ��e��hL���s3>��=�)�=����d>�I��^Ⴞ�c�<��>�5�=�9�+{�>�1�>� >EP>~�����,�j���4���yN��|
�Fv&�%������+��<���.��E�Z)W�{������=]���oM���½��~�9<�^2?O+?6 ?��>n�$>�_���V¾����qP��jZ���о�Փ�9{��)޾-*��=d��J�6�3�0��\�>�L>���>h?��=�<dQ<�Y�>����#3=�ܠ=G�>�|K>u
���:>�>I�^>��=8��>o��>��>��{�dc��\��=�.�;9#?�	��o��Ҿ����U��pn>?q�=d*�hrc�rc����>�R��+&�W&h�!��⩬>>�f�>�p>��L=;�ʾ@�:�/`>��>!�:>�
�=����5����;�!�>��%��%+��;D>WS_?�?���?:�=�S�>M�j>���>_C�>m���D�۽�� ?t�>I��>�ӕ?�^�?8;�=;S���(���ӽ6�Y��q��%�$>5`�=���=�1�=�=�2O>�b4��̹��>� =+��*�=c�>A{�>3?n��>	�>��\�?��%�&y���Z�>U���i�#>�>��?��P>��<�d�=�t=�Q�����D��>?wM>�+@�]����sD����>p�>	H?J�>�j�>6茾_<����>�������=��h?��
?9�O>uE������忄�*|�6�O>��������j���=<;1�!�#���=��E>��I�xˣ��?� ?���=��>���>��I>�x�=ۗ'=B��<SH<hؕ�y�<+�*���s>��>ۚ��(��R�U���n<�:q==x3=�����?��?�/��XN��H���5�)����-F?�<���?�>#?OzA��_�;d�EEϾJ���?�R?��{>s�s�:�<��H=���>8��>�gX=\(s=�1�\��
��X
�=Εy>w>��>ߝ�ѹ���3�����>6Ϟ=Z������?R0�?~a�^�<��(��WP�fX�g���������p���==��x�Fc��Q�<�ƾ^D����>�z�?9�w��=/���������_����[ւ=D�Y=�S?�M?�@z��%ܾ�L�� +�����va�=,��>�[�=��>�j/?mn?�x�?�>�	?m���x ?l�g>�ݾ=|ݾ>}Y]?mvf>�>�>���=zӅ>	�=*.�=W��<�F#�=;X�����s�=C�{>K�R>z�#>�P�)۽�(��0�<f⽩�����4�}国���=�@>�?Ҩ�>���>��̽��P���=~����=}I >�g>�+�(���)>>#�>�Y�>AN�>Cf�����s���f�쫫���.?�J?�x?Y[�;�$>��վ�þ����t>7o�}�Ѿ�3�ZEԽ�w�~5����e>���=��/>�^?&* ?V?��=o���f��o�7����.T��F�>L;>�N�<�|W��5��a2d�MB���F�a��bu��x=��>1f> �v>��>��y<�j'=_[C�K=��X�Q:�>��>ICl>��=>A
�=.̵�4�ﾱ\H?� ��������ݾV�J�N�>��>�g��?������x�K,���p9�6r�>��?���?K�f?r�6�[��y]>��\>��:>�Ӡ�MKP�Y~ֽM:>��=�FY�G����ͻ�Q|>4m>��y8��=:�|q� ¿�T����4�߾&_���پ+A��J�M���� >DE��3��4ﾳ���䌆��M�E<�������͝?�[�?`-�>��=�����cb��%߾���|����y��c;c�b�ٍ��6$�;0S7���8���P��;5�k�L��	�>:L)�����X���gb4�$�����=��F?*Zپ����u!��=�)>Ö-��y㾐9������ɽ�7?Ee6?;��b�׾�s �u>q�)?�4�>��E>1������Ɉ>	"=?A�?��o�~<���z���V�)�?�
�?
�5?a\D��68�8��+�J�|� ?t��> ?E���߸��;��f�?]	?�2>����M���we?\FE?{�2��SD>���>��>��ǽc���ט+�m�xeJ<�Ww>n�=�mA��sh�b�/����=�f�>Q7G>2���v��H_>���`��.J�!r���߽ͼ=� ?�V�ߠ�<���=��!>���ֳt����k����DX?�ޱ?r�X?B/?rپ_,��>�#�N�=���>AĞ>���=�?C�ߌ�>���>��پ�>x��Z�u�0?v��?�g�?y!;?�O���Կ����ٞ��-p��/�
>�p>u��>wF�B<>N�.�C�_V�=B(\>YS�>T.�=��>p>�>�]O>��>Ⴭ��,�t�ȿz̙���H���󾼥�':_��JȾ3���B�B���H��4���+>�g��{��>��Dq+��=u��%=��?��?���>�>]P	�~%���'��)�ξ��<�`#�(v[�95ž�~���t��#�<�f4¾G6��t=����)�+�T?�F/>k��>Q�,?5�"=.�$>�1�>�Y���R�����@>���>u{�=a����½-�(S_=�(q>3<�>�m �X��c\�������*J*?NW��o��>�0�s�4����W5�>��p? �d>ݾF��:���u�s#�>IX��P������罇K�>�o`=���>&�:=��o>�VľEM��[�=y<�=�>�>�Fݾ0�Y�#.>��>U.��r>����ǽg8?!�?��?��=P��>n��>�8�>ú=�,оD��ԝ=YF?�i!?O?��n?V�=/�A����=.�7<�V���L�{�0�X1>/�l=���=��>G�\���=YL�������W>���|��>q��=Xk�>��?�k�>�З>��y�r>��(�k��<���~Bp�
��>r�h>X�?I([�:�>�P�>T���ܾ������>��J>e�D�������B	�>���=�D?�u>3>%1b��=�=�g=>��b>W6�>S�?��r>�C�=wЬ�C���S翎��f�8���W=l��=���=��<;��>|���3@� �1>� j>�{�>x$	�����=6?���>���>��>�C�>~ť=�#�5><}�ѽNA���F�<���=#>>��s<^��=�}��{�p����=#��=lJ�<h�Z<���>�0?�X7<,�U��ؾͭ�%q����>9�>��?�E�>Z,��:��"g�\xҾ�=}>#}�>�Xn?sb�>a8�a�=�=Q+f>S��>K�9>h��<L�������*�t�<>��>v��>�%�>w�	�5��)�*�՘?>~s�=F쵾���?�@�?Ü��������`�D錾�����3�^�م��)�l��B��@�љ?��v��<+�=C��>|��?v� �`n7>'龽;���a��X���=>F�>�#�>��?OI��i���w�ž�<�F=4���s==?�>4�i>Fp�>�,?@N?��Z?ȕ�>��1?UHO�Ԫ�>o�N>ī�>�,?��1?K��>y�>�ae>�?:>n�U>ߕ��V���c�V����==��=8/D=_�>�^�>�{>�d�<��}�g$R�*�y��Z��j�ż"8�=E�_>$>\>6	?�(?M:ټ�1�U܏�S��sw�ï[>�r���T>7<}>��}<Q�����>��?��>cPy�ӿ��Ǿ��Ӿ6N2��<�>�}N?�?n�-��n�>�' ��(;��&Q����>X��=	�d�������)����3�>���>~/> Dj>��d? �E?��*?X�������_b�;�W���̼�H���M�>�h�>��=>x������E��bC��S-�*ʷ����=�y�;aE��(�?>��9>O��>(�p��^$���C�:�<خ�=��>�R�>���>\_�>�ø=WР�f���C?�؇����Է���;��;���=5�q>�"۽�??L�����t��;��ܣF����>�~�?�{�?;�f?d���	�|�P>0J>�H>�y�<�`\�:u�3Ҹ�-	[>�պ=�_����*��< )F>*U>AB���e��	�پȉ��S񾿣�?������ȾՒɾ;V��x��h�0=P D=�Sq�����׽�>{����v�Ҿ��F�ߝ���^k����?ʳ�?���>c�
>ɬq�t�����S�]����-v=pl޽P�/1ھxQ޾���=s-k�8�9��J5���S��b��Z������w��W�辕>�>�??��N>OEW�������>Pd?6?c7l�Ǘ��+�����U>O�k?i��>��¾�`ž��۽W��=���>+"�>.d�>�n�����<a�>��>lp�>qӾ=7c�(���|��=���?��j?�q@?�5E���=���=I��v?��	?b��>V���ȾCW��#?�5?��>C{� ӂ����Nt�>^�W?ʆO�F�Z>���>}R�>
?�#3��c���W���
e��9:>�!��~��=o��l<�/6�=(��>6�v>�JO��\�����>S0���N���H�	�����k��<��?Zo��9>��h>E/>ɰ(����qȉ����9�L?9��?��S?{g8?�X��9��������=��>�̬>Cѯ=h��y�>���>7h辡rr�|���?xF�?���?�ZZ?�m�Ti�쮿���dɾ�[�= %�=�~R>�*�H
>ؕx>�'�� �
��d�<X͓>��>	A>
 �>��p>�U�>c����&�ж��k��C7�� �5:�Z��w���2>�
�Q��~¾"����R-�L���總��<;�!���E�L�c��hH?��>?&?�"�>���>����]�-�߾�	>S*n�Z�5���E��� ���þᖮ����-���_��	$?��k>��>�{�>��=��(۾>��>e��;Ĥ�=�>��<��<��>��X>VS8>b]�>�@�>
��>�^h��k���oZ�'\>������	?�m���ӓ�	82�G������<�V�><��>�0L>���3W��L��"E�>��<���F����eJ�L���w�>��>~5D�wx>�<P�X2������=k>��|>A�?�j��������=l��>Ԣ�Xv�=w<�=C�>.2�>��>+U�>W �>���>�*��.�=3�q>$(�!j�>�@1?&)?��o?=/?X��<I�3����<饞=�/\��^�}=��;��C=Xo2��nY�9��=�4�=�H����=8�+=���ϝ=7��Vз>Wz?�N>�ܕ>�[��z���n�s]e�.��<�˾։�>��%?�-?��>���<ݘ>/�=�ݦ�����?(��>3_t�����r�=գ?�,��Wv?�.4?�3�=ݡ��Y�о���>C�=�G�>f?1��>с`>�KF�ɫ�����H�W���Ž֦D���;Ll4����>���>�XV�	Վ�V������<��!�۽I��=r�>�`�>���>7�=ې*<a�A>�e߽�ë�Ocۼp�����<�@>e�_>�C>��:<e��a�V�u�Q�"��۠��U�=�x�>��>�Q������
��)�
�������?~�?6��>_~�=$m?>r��F8��t5�~�>0*?��<?�?uc.��7(�=r=]>�H>,҄>繳>徸Sھ��Ͼ��A=ۛ?��4>,�?)磽Uf�<J�v�9�f>��=D;뾗��?q3�?u����;1�پ�:a��!��⓾}�>y����ʾ񿽽]�F� C���b������=B��>��?3�5��,�>�8��8(s���4���־�>=�Q��Z��>s��>4�̼�37���߾�ݫ�я;>��=�|�=�~�=<��>O::?Ռ'?�|?�>7�>O��`3�>b�>4��=��]>�?p��>P6�>�E�>k6�>��>�Z�>L���θL�k/�Pm��¼�^=��~=<0>�#�=ڳ��_�o�ˁ�2�Z=N����=�J�=��D=!�U>�	>��	?�;?�J���ni��Ǧ���t�����gʧ>ឃ�+Q޽�_=��S���3=K3>�f?6��>���i�󔳾g?ܾ6��}7D?:4?=�>�~2�Z�@��ꋾ���=���PB�>��V��%dz�S�پ�{E����:[�|>~	>��V>�ru?�4?A"?�a��0��Md�1&�D�~��]�ʼ�>0��>�=�<�u��y(,���g��wQ��10��-��&2��)=Ow�=4>"vK>�E�=��
>9�I=�=ؽ��2�<�E��e}�>���>�(�><PY>6��<Ӣ�=��B?䳌��m�i���Ͼ|����=p�o>�\m�?
u��$v�����_~B����>��?6��?B�f?�&��t���C>�$q>�z)>V$��O��w]�	w۽_�2>_�=6���ɍ�������`>?�]>h�#�K#��Ej�y�)ɿ�b��䲾�����;��j�����t���W���i>�9���E2=�p�����(��ڭ��2��s���n_�P��?PY�?�%�=P�޽j�D����;��?tȽ��H�Ȋ�ͱ�;5n۽���}N��u��� ���xe���x����>j=m�ߟ���o�R�:�0i�<4�>�l? ���)J���Y(����<Cz9>=L>
���)���5��������-?�*?��ؾ��ؾ�� ��9�=C6�>���>O�>軔����>�g(?y"?�i�:#ݑ�\˅�"ɟ�蛳?���?�OJ?����?��쾍�8�ɫ?B2?�(�>�d��f�Ǿ�s��j��>v)7?!��>�,��4ty�*$��Ԍ>�{?��X���X>�r�>�8�>�>��菫�d>ּfK���y�:nR=U�=�g�7FҾ-@�P���=K>��>�
������>(�龛�N��OH�F������o�<�U?^��"�>,�i>kA>-�(�)�9���jY�L
M?�q�?�nS?�8?�������馽���=�[�>���>�Q�=Cd
�z��>
\�>��辰�r�����t?�8�?Ѹ�?DaZ?�m��Fӿ�
���������n��=%(�=��>>��޽ĭ=��K=�����Z=���>3��>�o>H:x>{�T>'�<>g�.>3���L�#�oʤ�<ْ�[B�� �9���wg��{	��y����6ȴ��򽾍���Š��wГ�X�G�@��XZ>����;��5�7�^?��I?X��>�s�>�<�>�ѽ~{��L
>+����3ƾWN۾���f���Ͼ>]D�ì7�μ��6��\!?Y]���L�=/�?0]t�ӭd>��>����l�E=�풺3A>�(z>���>к>��ս�4�>[��>t�x>�Y�=bc���$��k�W�����6��M.?��z�ڻ]��䦾�'��[־b�N>��>Q��>�d��N��sю�Q�	?�2���w	��(bi<��>�n�>)6�< u��98�<�	x��ˈ�DJ�=e�R>?�>A�P>���J�6wW=���>��n��Kt�f*=}�?�KS?�?oQ>�;>'�=�x>�`J>�66>\��>u��>(�>�X?)F/?A� ?��N=�,��F������<>��DK�n�ܽ���w��;���C&�=q���.5=.��;��^=����Dy�H�9;���>�8.?���>w-?^���*���X��!L����>#ah�!�(?"�/=��X>�6�>�?E�v>Tǖ>��y�پ��?v�#>�ь�*	����1�m&?8۽�vx?�?��X��ہ�յ=���'��?��>R�r�۶�>�Ou����u����y����$.$<���߻3>6.ƾ_��>u!������[���o`=�V1����Z���t-���>-��>d>>�к����מ=���=�9�p�>�$o��?��H>*�����=<`#����=��=,�b>�b�=��� ?%�N?7�U>�X��b�>KLξ��>o�y�1?,!?]<?擎���5��p��s����>;�C?�_?d[? �F�nw ��%�Q�a��>��>�p>�mY�5��1�`�*�4�=}�>��2?���>��[�E��Ic]�ď���^�>�V =�����?qg?��Ⱦu!>#6,�Wh�c��<�l�<A�Q�Ε�����5��y�>�'���12�m��>�֟>z�?�Ӿ�/>g�R����BO�$F�E4G�|�d>��*?���>���k�쾡��㦼���>c3;>���>�3�=�4p>h�?�?��o?��(?0cK?[Gq���?�⍽��>wU?=��>��?���>@0->K&	>����Ps=9}7��;��D�:x�u��-�<�^�=��9>��:<�R/=�F=��>_=:U����=(c=��=<��=�wD<G��=�h	?��?�~��J׺=�K=
tĽ:�}>X�	��f�=�/"�(�^��?>n]<>�_�>�[�>�
�=⪼s�H�2�5��0 �_Ƚ��%?|�7?;0>��T����a���8�G=�8�<ǜC>c'(��ʻ���ͽ.�Ҿ�v���NK>' ���z�Ɔ>qi?]??��5?CĻa�#���C��#'�X��L���
�~>�D�>4lQ<rC��Q!I���Y�JDI�d�G�#�7�~���"-m�"G�>�Q->�6�=�O�=�47��[=�/��I��:�;A-н���>C��>y��>��'>lb>��ܾ�D	���/?O<��A�-w/�@�P�b\�����<�Dx<�V�=Ж?_�6>��q��ײ���X�K�>���?Q�?a�B?yx%�0oؽ��s>�>s=�Q�=�f>�����\�*��5>̲j>m��Iܽ��ݽ2~K==��>,��m�d��#ɾ��L!ǿy�p�����f!�͸�'��C���:���$A����>����R���ay�
!��d�ʄ9����o?¾ؾ.�?Om�?�=���=w��_��{��]Y>�
C���]�]W�.埾̐n��s����Ew����ؾUW�����>�'"��x����c�@r]���=��=�;?�����ƾ.i��,�<_H�>�͸=Q��UX���}���8e3?��@?"1 ����������>�c$?-��>�>P��Sr��=
LP?��S?��>�I������2eؽ8�?��?�i?�߲=Q�N���J�<����2 ?A{=�i(?p-7�
H&�����1?�I_?!�?=�A�Et���w?��?�i����=z�>�ˁ>�
׽3#��2�*>u=��W�8>0��>.P���u!�C%��p�>�;С�+�T=��X>�o����*�d�>�b��pL�0tD��"��h)�#�0�0�>d����>���>�p�=���|���ƅ�����D?8��?�L?�2?�$�`���aA=�͒>	��>e��=�"��3/�>��>Z��� w��%�'�?'�?�
�?��X?�Xl�����笿�:���$��]��=��̹vOw>*����>!-V<R�ѽo����e3>U{�>(-�>���>�(1>->q)�>J���--�c��ߞy���:�{������h.��6��D���d.��iw�ŀ���\�����Q;n����ͼ$੽�wU�����B?�^:?��>q��>�9�>[���}�׽�|=@z:��D��#�K�Qv0�S�������f���W���E�;����>/P�<�H>9�	?��y<j��>�^�>���=��2>-�m�e�=�n>�;P>��L>c|�>�Vr>���>e��>%"6>�M�x@?�I?��k�eu���?�/�\d���N���,��kT��b��ܙ>��X>�޾�z������e��>d�\�8�>�m,%��?� ��>���>T�<l���=na��*�=��=�A�>tU<��ʽL���gW������@�2>��:�V�^>��>�YR?y~�?ln?��>��??V�=<M>�s=���>d�>�o�=��>�?&g�>�xk?Vj=���24d=$L�����"��P*�e1-=����8R�<��V<2!>¸@>���v��>�����5��~�<N�����>��+?���>I�>����Zo��i�m*Y�� �>�R#����>,>�=�&>��d>*�#?��>2�s>9;���B�Go�>�9}>�Ze��Ӆ�nQ����9��S���h?�>�>�>hE;�8_W�9ŀ���B>��? �>��^>�X�>��Ҿ�� �=���v�B�g���(��*>�e�M7>�S�<������:�lš=���=�E�>���>�B�>^��>�T�>/
�>��2>~��=�{�=�p==G�.=��='_=��;I�=��]>���<l��^Wz�%�f���<GF�=+l�p_�>�S?ǒ>�J��>�;� ���J��f&?w:�>���> �>�v�G�=�{5��=>D�\?�"2?�_?x�����W<`i��V>���>jL?��>�)x��$����9� ��?��!?��>Q��>�p�(8�̻���n�>R�=�9��<A�?s _?�dƾ	=`�׾`�+�O�˾؏?;Q۾c5��ٹ:�K,G�8�#�Yk�<�������uA">>ڵ?�ܾ��9>�� ��q������B��4q=E�6>j??��=2<�Qоjzվ���=<f�=p��>�,�>�٦=��*>}��>� ?,B?���>X3+?����/�>�jH��>�^�><a�>�?d��=Ѭ��	�;�=?W>Ѷ���a�&ҋ=e����F=��=���=%Ы�1�\=���= Ĉ<��5��# ��:��`#9<.�=��=��%>�,a>�A?�?�B,�)�<3Z���@?��kJ=�^=>R�=n���*ͼb�߽���o5c>�>�s?>W��==�������ľߡ<Ts+?��?:�>B����;�����)E=yNO>iUo>�Y�4I��`J�v�j�p�>l�>'	+><�f���l>;�s?�[4?�i?1��B/���t��[�K�?=c�뼊X�>]�6>�
<֌�O�+�(O�T�S���0�����2i.��?�<��>��">�">:=�Wp=�+�=�8n�T^{�u`��Ň�,,�>���>ƶ?gu�>& H��DľK�t�3?1����f�q�>���ޝ޽-~�=��U>��;,�P?򥳾i�p�j��ÀD����>@��?�2�?>� ?eݽ��(�>tL=t�>���;J4v>d�d=��ü4o7>>�>����=R���u�<�N>4{#>��v�NcR��B��c��dϿ؁P�"+c����ξ�[ ��Txh�=8�<�c�G��������R��xc;�Zؽ���JH���E���u����ʈ�?o,�?8�zF��e�w����9%����.�޾��"���{�J;�nȾfG���ܾ�@�l)E���;�Ծq>�X���v����g� ��=V1=��+?\��J;���K�����>��=�䏾��zI���B�<G@	?)�;?��ξ֦���𴽞�!>��>ļ>��>-m���^���E>:�J?�q?#l>���Y�=9��0�?j��?�	�>�C>��h�M�3��Z/���;>��~>x?�>I�?�*j6���M>��?i6R?�G0?�W������/�N�|(?BB=�q1�v��=j�>���>�Ƚ[2s�mS>��@�Cd�>�j>c&>Re���
�����/�~��>�:	>,}��Ӈ�w��>��Z�N��H�u���o ���r<n?�Q�޷>��k>\7>S�(�_����v�����A�L?o�?VR?�G8?������e���@��=F�>e��>W�=�
����>��>f_龴'r��z���?d��?Z��?��Y?��m�̬ؿ�ܣ�S>��:����	>`͌=��i>��ۇ=]6�=�"=�Ė;�Q�<��_>P��=�  >|A?>ze\>n/d>����{/�ꌤ�䕿&�M�+'�KP	���������V�p������5;���h�%\Q��r�f]��;I����h��� �3?[��>�y>ɋ�>���>[��{+��:^=��, N��;"������7���e=X��������վ�m��)<�+�?�-<xf�>,�9?����,m>1f�>k���D>u=�~>�*�=B�+���=S��>�A>rg�>h�B>�G�>�\->�%R���F�G�M���d���/��k?쵾�j��e�W�
����O�1�>|�D>�������������>�|<O�<�K�0��:�
�{>�@�>"P�>'���!w=����4��������>L}l>�ic�$�ξ�;��_+>)Đ>�8�}�,>��>��Z?`��?͇c?m���F�
?Q<h>�L>���=��
=��4>�C�>V?ˁ?҃?��1?��=7u��>��ې��慾�$8�� ��?X=8q:���=,��=�/2>9�u>f�=W��>;@M�K�c9[B=F��<�
�>��&?�ڲ>��>�0��P�\��]m��\��*K>���<���>en>�,6>޾n>w�?��>���>���W1��(?�x�>檁�<��L�d��b>m�m�?�.?��<r�{䰽ۛ��=��VC?�{
?&׽>X�>��x�N?��6���6WE��i����B���7>��Bz�<�h�<�<����eJV<�>f�>ے>�i�>rd�=bV{>`?�>N�h>��>h��=��I=���=�Wg�I�>AKм�A�5m<=����V>�Y=�`	=̇���ܽq��1=Д?��<?�[�=���<�Ҷ=��������4>E&?�?y�8>��=�%�����H��}>�fN?~zW?�?\Q��
̤�C���ح=��>���>�5�> ���S.�q����}����>f?��?:DK��;f�È6�f��a �>��*=@Wy����?�Mp?S����= ���H��a��^|�>� ���X��f潟�]�!��y�@<��*�䕆�⾜=��>H�?�߾��g>���r��|�x���:�q��;�W>�g'?��#>]�_��͉��|��#A���/�>X`�>��?�l�=&j�=
��>�,?�0c?��,?p�E?"3��40�>�jq����>���>�> ?!+r>�
]=p�> z=r�V>x�(����  ��J����\>�O->���>.=�X|9����=�p����=�t(=��>I2^=�oj<�_��R�=h)>i�?�k"?}�ս�j2>�`��g����>���=κ�>�E�Ӡ>!�>;78�-�K>4��>Ĝ>�����`�Y�'��-�/�ʽ�@L?��[?WБ>'����8�b�ᾗ�W�?R>�y�>rȾ��>~��,7�3D�6F�����>M�@=2����\>�d?S�B?B�H?�&)=2�0�9cg��=�{噽��ɽ��>W��>Q�5>X<��$�O�X��0�N"� )�<:�'��=�F�=��(>[!�=&�Ệb>H~=8=Q�L���|�F=e�+=��>���>9�?=>I2�Ū	��(�/�@?`@M���
󆾱I�����̽�<���=۞м�?_0�4�k�h���9A��}�>l�?v��?�oh?�뽆�ڽ��]>�>�P�=�q=��:�[n���,��~E> ��=����l���t]Ӽ��n>�|M>���������ξhk�����E�	���>������	��啾�=�#?�K��:��ž�EѾrr����[��
�����l��	�ľ���=\�?ţ?��=9�V�Z��%�%A!�0�<��s��{�nZ��A���<��%�վ\��,l���Ѿ]�#��M�4v>���M��zΌ���@�7B�<_��l@?[�P��KӾm��:�\�>s�>j��I���e�h��1-=��(?X�<?kʾ��!�T��_L�>L�?mZ?�tj>vc꾈���",S>l�]?��<?��x>I�i���������2t�?Ae�?�?�v�=77d��[%���L����>%��>E��>`�R��U$�&v�=Q�%?1�l?��?!�9����/u+�.ۚ>0Q�=$2�~��=q(�>�4�>��`�ܲ��Ќ*>����G�>��>��m����VE�M����6�bo�>uɬ< :����(�A>�>�h�X�K�PG��
��G;�eV�h� ?��Y�>2�i>���=�I*��C��Ö��3���K?�8�?�lI?�P;?�������:쮽8{=�ƥ>.�>L��==T����>�>��2m�H'��^?C~�?X��?x�_?�k��&��$yſaľ��о�>�c>�Fj>#4���G<�|b=PVg�ġ<E��>.�>8se>��C>!��=z>ʶ[>�����(����HE��:?��X��������t׾�;F��-�����	����ǽ㫛�5�<���<��<#w�T�$��`�r�U?O�>p�C>:��>N��>�ʗ�wy��XA���S-�7$a��������U
�Ϡ�����+�vC��h5|���=�c�?1��=vg>L��>$�H�1I>�>�˙�Wi>B�>�'>?oٽ�+X�{�J>�g�==��>��>�۫>���=?%I���=�$�)�Y�E�[r==q�?8���8ٽ�6������q���^>K��=�Z�>��S���ߺ��,Ӕ>���=�bN<�,��u���u�>8�>�:=;%ƽ�M�<Yk!��r�<IVR>N�L>�P�>m�� %ܾ�n��}�=�Q]>��P�=�`>-w0?�؅?��N?�6���>�?>�Y`>i�=0��>��>G��<,Z�>�w�>��>��!?\��=��V��o�<hW��z�e��0��ca>~z�<<��=�"�� ��=;��=L���5��w�;�zB����7�<���>�?B��>�/?O{P��vp���[��ũ�K4>9�=Q�>;�>2Y�>�l�>V7?/R�>2*�>i�\�����my?W�>�����K��J�=�p�=,�j>���?�?C�����4��=�w;��>�ϳ>R��>w^�>���>F3��f���쿴}�(��'�<��:=��=!|�1�<���b���C@�=�|>�Ak>0a>:W>Z�=7`>R`�>�E�>���=��4<k���<,:b//=|�ʼ�oD>組=5����y�_9�%"�=`	j�`%�O����<��>C�B? W�=�x�<ĺ�>߾�t%���[��mQ?�J?;��>���>�E�\�����Q��>��Y?�4?�T?$/��hL���sý!ü�c�>��?#�>ʛ��о�6�ᚥ�K=	?���>֦>W�q��/�^Ⱦ��h>�9�|���]�?*(�?�|ؾ��˽���<p�C�����>�M往�`�hp>@7�f1*��B�T*����fq>���>�D�?�+���>�4I��#���zu�'��~D=\��>6�:?�,>��������Xʽ�>��>-�?���>�\d>�Q�>]3�=��0>T�?Ǡ�>K�?��k<(�{=��I�A2�>53�>���>]*�>��>�;��G�6>���=$˷;^ɣ����*��=��=�j,<�־=q� >$.>�ة�=��=i�4�����3<e��3�=�>̕=�y��Ϳ>�>��?�BL���	p��;��ح=(,>�.=�/�=i=��	�����<��>/G�>�k�>�DC��Ӿ#�۾z־lG=Jk?|)?Ў�>V�jw������O=mY>�[A>���F����<��#r��z�X�>w�>t�-�ړu>��l?E{9?�ED?k퟽����#=��\1��[=lط����>�~I>��1�I�w��:�c�`��aO��B9���z2g�E�<�;~>��q>�>h%�=�4S=JL�<����Tt��<��;�/�1T�>b�>\�?��^>�c>�P�hN��zF?E�\��Z���3�揇���.(�=!�&>=tּ�l?�(��9z��Y��c�1���/>Ǿ�?���?<�7?��k��<��)4>�OP>i7�=�`>u�!��Z�`{4��Y�=�e�<먲�������l�>Ȅ�=�C��ɂ�����46-�p�п��S�O��G徇�վ8�]��fY��n�%�e殻"���Ͼ�I���.ټ�/�z�J奾�:Ⱦ�v��
;�?2�? ->ls���2��C�`�ăV�޺�=�E�C�G=*�(�[G��!�־�¾x&�%��<����8�n��QY>
x�)*��k򆿥{R��9 �u�p�Ek?�������tf��A��;,��>iQ_�����u�CgT�;%>>�>��=?0޾\@�H����>��'?_`?��>����Y%Q>�&G?��P?ok>����Uh��7ݮ��o�?�N�?2?�=��U�t�� �V��S�>\��>�?�v ���A���>m ?���>@��>N�6�Q�P��&��?4h�>$"��F�=��>�>o᫽��z�C�>�r	��ǣ=)�>\`=Z̈́���	���ʼw���n�>0j>�H׾/�*�V�=���&�:���P����񮉾a���-�>���D[L>�Ӧ>��v>�"��*���u���Yľ�?$�?:Bc?��2?	Ӿ<_־Q&T����=.Ǔ>�R�>v�=	C��ɀ>�ƚ>3����Y�����>���?�A�?�??h,��:�޿b���z�������X>뙚=(�1>W��/�=�˻��M��c�$��=le�>�Uu>�g >:�>��S>T�?>Ȇ����'�����qi���:��@"�Ar�Q�J�E��T	���3 �v��"۾v1콶
��J��N\�9�ʽ���c���_�'GM?�"�>�Z�>A�?��.><'0��1I���V�s0�iL8���˾걉��`���ٻ0"��s�-��E#����0�.�>JS~�hB�>�l?��=F@[>Ի>�P>���� �<������<=���>��
>�;>!��>���>p��>�%>�TN��66�S5'��Ƅ��hF>\�0?Iľ�:�����$�����=���>�9�> ����������>b
�<n�ջ��<��۽
�=>K��>Oヽ��<�2�XB�y-�;2\`=���>��=p�<_F��N��Ch=���> �ľ6�4=X��>�O?�0`?��Q?ou�=�օ>�#�=Q��>��\�v��>.�_>d>�?^:?bj�>�?�n�=3�y�5K��q�H<@�Z�"?�<�c�������t>� �=jz>�w�=DM�=lr>��Z=[UA���ͽQ>ƽ�5�>�:?4I�>œ?඾�YL�DF�r�ݾ���>�>L$>Y��>w�=��B>|�O?m�>�o�>'좽�p�bk%?���>Sk��l������Z >��ż#��?��
?/b=�F>	��������=:?J�?��?M��>m�������>쿌���6�0Z��=\���.=����b�:'����5��C,������c7�J�t=V�H�j���Ax.>C�>���>N�U>��]=ǽt=%��
_=���=E�=�(=TP= B����;4J����f�&[��l����ʎ<k(t=wO?J�??�Б=3�<˳=}�ʾh��*�>�C?�K�>��?���>�P��=��D��+~>�m??��-?Oi�>�0i��ጽ}����u)=Och>�?S�>N ���g�#WC��?2�m�>�3A?�T?�Y澥v����-��樾���>~�=���N��?u?$
���>����#9�Vb��7��>w������?櫾z+�sf��ᑽ��9�<�վ��=xO�>p�?J"��w�J>�v��q�����3�6.V>�,-=M�(?�%�>E��������nr��K�>WA�>��<=Q<>��L>�6�>�e?M�_?�o?��?*!��>\�1�K
�<=\�>��
?�?s�=�ވ�g�=y|�=α�<:b���S����=�Ǽ�r�=H`>�q�=���<��ϽU�>a̤�Z�<�Û=��R�>�A�<�)�S>�<��^>��?�?٢�~�<�o�1v����$>|p�=}��=��3���V<���=�*>Yo�>�BB>���>-dr<��ȾSRǾ@�� `��NP`?�Y?���>Ų��(�ҋ�At��ƻ>i��=�䍽�˝�����	���,���=��ѽ���
j>��s?lI?�	3?Y����=�jUv�+�5�9=��>�I��>U��>�:�=={ƾn�0�g�h�0�H��-�ϛ*�X�?�+<܀">�2N>��J>4h�=e5>�p<퓱���Z�U�"�9�Nq�>��>

?�8D>�}=%y���N �B(G?�/��������{.��?�����/�=>;�U=i%?��<�;�,ò�o�S�M6?:��?��?O}O?�Z��1���4�>�g=Req�[�*>�<������=�$R>0��	��Ub�I�l��29>��>ט����������};	TڿƯ{��yc�j甾��׾�,��CK��־�����6�=��������k�;���g�¾��1���,�:�$�����?��?���=�[>.�B�y� �.hȾoL0��$���>lɈ�w�69�G= ���μ�1��G!����y�d�<�q��c��`����I�$T߼?'=8�0?kǽ�&���mfx���=�J>]�=��ƾ�퐿�a���)=� U?�+?�l���|Ҿ�fe���>P�>Y�?>w��>�3��ܓ��/�>�M?��1?�/>>�){��`��-t��'��?E	�?���>D�>o+]�]�D��@�� ��>�K�>��>?��O���:���=��Y>�Lw?]g+?��x��H�tv]�,��>%?d�/�I�u;/��>�ش>J�#�Q�ž.���$��4��=���>�j5=�۾���x@վ*4����>��!>��)	)�51�>-��9����G��뾈���k� ��V�>
�1����>�;�>�W>�k�����2��N����??4ظ?�?M�?��ξ5 �Ȧ�=8�w=$��>F�>����=�L�>Ā�>S�e�������m�>m��?�n@C�?pM\���ڿW3���L�������n�=o>|D>���%��=���=�*�=�6=F-�'�P>Uc�=���> \�>��=>�Q>�
����(����L��R{/����g��2aV��ݾ�"���a	�rW��k3�����;E�N��*�A�D�]�D�!�����b���$>ț?:n�>
� ?�y�>J��<}�þ�F��ͽ6��e@�]��Y�'{�@S���ӽ!��������H����I�
?4M���j#>c�>�����|=f�>�>�xs>�Y>��>�^�=Þ>&O>�ݼY	>k��=��y>Ǳ�=�-��琿�o����'�p��>j��?~�*��=M�:�y��r0=/�/?��8?w��>�I�s9���늿Ϧ�>��)>��оba��ǽs�>El?��E>�`>x#��nƾ�G`�o�0>]��>�S�#�`�<k��Lm���Gt=Fv�>i칾��>���>]3?�܇?��?�����M ?�Դ>̣�>l�߹�P=
�=?@=�d�>��?DM8?�U?;��=x(���q<9N�=[�N��(��C���ɉ�h�P�8
�=-�Լ>j>CT\�nū=�$>��YҽF�O>�=uz�>l�"?�>��>H��<ww>��=z������>&��6è>y�!?��D?��>{S�>ʀ�>�Y�ݧ���Ծ��>�>НI��a��!Ƶ��'>Vb�>�\?�K?��x�y�Vp>�+I�=t"�>��F?��(?�)b>@�$��7�����ؔ��s����G:=Rc>��[�����ӊ� �=�[�7�ǾƎC�k{`>��&>��2>��>�#t>��L>�>��L>O��[c>ڼ���fG�.��=���=K��	��qp�9�ӽ����t�4�,�+�����<{&�=�r���?�>?�F>�tQ;.����h��{���<;>�X>h�)?��?��
���@��s��c����Ⱦ�?�}?�71?}F���{=�/����c>�g�>���>�~�>r�"�p)>�����)�Up'>�)�>[?'�O=����j�UC�RS>��=�����?ՆU?^���=��<$���kI�����>,(=BRQ��?��-�%���6����]@�q*ڽ3ԭ>���>y�?���{> Z���������eI*��ɽ񐁾���>��#?�H�=D���x��|Ӿ�W��'����'�>�>���>)�]?��y?� �?�R9?s��=��Ri;?X�G>��>���>�\?��>��>#�?��?1vC>b!�<����;R��x��=H��=% �=I �>�ܛ>1�Ǽ�o����>c >S .���{�i=�:a���A�k>��> ��>u	?9)?Go�� ��cZ��}x����?H��>��>�I}���o,��s�=e?�H?�`�>#�1>�������ѾpD�+r?�L�>x~<?cw�>�e�<�=����4�>��>�/v����y�0��|���ｲ�>�>�S�>�x>�Wv?v�L?��:?�%�=��������9�|�=�����>�??K��=���x�;���K�S�Z�#;!�Ď�=g -�rz�=�����=}��>}�Ië<F4�=��=�:�9�<2�"=��>��>�?�t�>�h=ľ} ���I?3P���I��ޠ�P=оa����>�<>/��ާ?�����}�����7=�Jd�>�h�?���?�#d?s�C�/c��g\>�:W>��>�.5<.�=� 5�� ���K3>mi�=>/y��!���Ϟ;��\>�Zx>�[˽��ʾ��㾻xE� d��#q`�����%�K���ؾ�i,�ѓ����$<l�����E�Ʌ��p����޾�����=DY���^;����ȾH�?۰�?�k<�3�[I_��M��Ĭ����>$�v��U��O¾�-�=;��F�
}��ɾ���[�E�J�0�h(�>�,]�;af��w����na=�_D=Rk.?��%�s*?�ِҾ&�7>���>t�:��L��=��q6��9.=>�#e?#�;?j@���d�׼���J�;��>,�*>�҂>�������94?xg?��9?!!�Ǘ�ё��� z�Kh�?��?�C?�u��� 5�����o��a�>���>���>5U��oA��a��Ȋ?��O?C%�>G�QE���=1���?ҕY?NI,�tx>�I�>�j�>�ۉ���h���B��8��7��9/w�>ߙ�={\�8���G���C/н��k>	 �>�f���2D�E��>�׼��D���
�����������;�>·+����>k�&>던>���"D������{��E�3?�X�?So?xe�>d����Xh�{#�=A�>�8�>�D*>C��=�>�j�>i?�[)��8� �ݾ��0?�j�?4��?�l?ʩ���(��d�Y�Y���4r�����=�	�=�0�>�����מ=��;TDü��oz=7�>��~>�6�>�D�>D!>&v
>E��	����e���cq�3�K�@���f����B��=ʾ@�A�fa��<�^�=�@���%��,ֽ��ְ�#gO�=ǒ���=cM?���>ܡ�>��a>cb�=zǎ��H۾�DL��T��/�C������5;�@����4�;�T�s��@����g ?�*#=��5>���>z�y�Τ�=���>WMf=72>��	>KZ�=BT9>*��=��3>��
>��a>�>-㾹�����V�o��@S�,��w��>c�B?�Q#��о�`<�������1?�>*?n�W>��\͊���h�d6�>�*�N���	��<�2.;�oW>3�>�҈>��	>���=����V0����=4�>~*>%��<D�)�=Xu	�L�>���>	��>��V?��?,F�>�ѽyV?�V�>��>����;_>a�<F��=�j?	�L??!(?�u�=Ĺ�����=�1�=�����N`>�P���f(��k��0�����=�Hv��`>p�=�V��wy� 9=���=TY?K�p?�?(?w/�=f�	�o�w�I�þ�d>i	�=u�?D�?��4?瀽>�>Y�M>j�y=�1��TE��R�>c�>N�[�`{x��%��*
>��Z>Td)?+1?Òi�+@���ʼ�ӗ>���>�%?//3?V�>'7,=�C�qk�>ſ'��3�#�n�Ľ�����<�����G=W�d<_RG��_���X�Di�>n��>���>d>�1 =�9�<���>�~:>��0=��=�Ѩ<[@�<F����;�ွ�M���0��8��<��c�80-�"@齂;������p�4��5����?�?�+�f�G�ڤF��;徖�����>���>���>x��>�=&����3X���?��;C�X��>��e?�I�>��#���=E	����u|�>�Ę>ց;>�!��g���	g��2�o=��>�/?��>�a���N��dk�[n�||�>w��=T~�H˞?>�z?�G����=O�A��|^�u�M>Y(R>t/�؆��(���&�#׾�˓�t����:>(��>~#�?�{�%y�;?;þ�᧿ ���b����=ɨ�<�%�>��>6�=�%��ݺ�� �����

�N�TA>9O�>!G�>���>��E?H�>���>�[J�1)?3��=|U�>�؃>X!?�?�>N��>���>$� ?M�ļ��5��핽��e� m=t��Ȉ=��?>�v>(�<���=`<d<BWz�yr�O�T��k��E�=�	>��>>�>�#>���>���>­
�L��V�O�����=�>�K�>2��Q��~	V��O?>���>��.?d�?n�=����_羑"��ۤ���� ?P�/?U,�>��=�0� �.�!举�j��2fa>�>*�~��L�����	E��D>׍�>[�>}l>1�}?&7F?\&?3�ӽ.(���w�Ng,����9�<��>��>��=����-8�p�b�Y�Y>,��Ｓ&U����<�t�=�W)>�j>�v�=�#>,C=�a��2��\/V=c�z��[�>��>�?� �>�ή=#��v����I?�����[��٠��Vо�����>w�<>�����?����}�� ���C=����>q��?0��?0d?��C�B3�ڱ\>�CV>�>�I2<��>�1��[���{�3><��=�4y�#��Z�;A�\>74y>�.ɽP�ʾ�&�}�H�]K���/)��f���Ⱦ�7������W�e�d��z�F��K�Έ���F�yމ��q����<�Ľ<K��ْ��{�̾j\U?��V?�*��o鬾x���&���ZϾ]�>i���'6������4�-�����K�?(���v���D��x��S��%�?5�7<^�o��Iy�&I�4��<�j>:�+?�}�����?�>M}#>9[�k��8��\����$�>
�S?8�6?Ev�Y[ܾ�r�<�ѯ=_s�>��>�\?>z�վR�Q�%�>s:?+-�>��.�͕��|��w<(�$
�?���?�$j?$���^p�����]Dt�c�>E��>ݒ�> �7�2i��T>4�t�F?�P?�]�2n����7�"���@?§�?��-���=�p?��>#���`�K����Dl��%�E��9;?��Y���ս��6�k����R�=�و>^~�>���J�N9�>ѕ��
L�
�E������x�<EH ?�n��>�*h>��>E$&��(���뉿&@��zL?[D�?�T?�6?G���RC�������=���>:{�>�U�=Z���ʟ>(/�>=羦�r�R���9?W��?���?�W?�Jn�Eο�����0��P����=	Y9;O!�=>{ڽ~�y>��=ԧ=mo!����<��>��>��>��>)�>�c�=(^��-/#�q\���i���x�CV�(��)���۾E�2��4�:o������P죽��T=��c<�ƾ*�z�3|�V��#��=��>F��>��)>L��>0>�3���f���Z�i�׾�i3�����z�����xO���>�*�@�L77�N��CG����>E2���>�>���>��<��d>m��>�����̋="�U�w>]�Y>�B�=���>�L�>h�=[����Yڽh�>B���ũ��>\m�X�پ}W�>XV?蝅�5tA���a��<��оD]�>~ ?�@>s�V�͎x���7����>q�=����Uֽ����)�>}�>��Y�5�>�6�=�ꤽEʀ�_M�LH�>�����b���4>�כ>2b�>9~�/P.>(Q�>�W/?��?0#+??��\��>`��>�L{>Z(��"�>,�%>\E>�A?mo8?%�+?K'�>:��=�^���A�=w'>���Z��.�NU(�,��=Z��=��z<��=2�y�N(#<״	>ߪ>w�B=��U�!�P<�d�>��2?���>�H�>֢]��U'���D���!�v��=k��C��>�b�>��?��>'7�>�xJ>��=�s���Y	�>�6>��p�C3R�N&лcyO>��>a9g?�9?���=C)���>ӌ>L��>:�=?�X?�i ?-s�=VdX���	��Կ��!����矽Y���A�L���8�`�Ǽ���<�8 ����Q�Ǻg�T>Ϫ�>��>�.8>vo>�(>���>lA>	>�=��=�e�V4�;�<���E=��P�O�O<}]���We��5)��N�y�x�b�� c����騢��?�4#?���=���(3�d߫�bu���2�>�,h>q��>��>0'>���rm��B��H��4;�>�4x?��?�ԃ�O�8>Fp��7A���>C��>V٠>���=�Ř��T��!P�=���>�p?S
�>j�� �^�|�i����ul�>�>1*��I�?���?%�û;�J>�X�.!x�&�ǽ���>�a7>?�"�eޣ�[*C�S1�4���/�����b!>�[�>l�?S���ƛ�=�놾\1���Έ�8H���pm�r���1S?!�>Br��x������){����ʾ�����+f>��;>H�>*�>���>�j1?ƨ�>�?��d>�=?4�=D_0>�Z=���>�EV?A�!?��?��?[顾�I�ћJ�DbN��ی��U�<hL��*>qZ�=Ts���>V�>e��=*e�b�*�5r��H�w=�P�<TI>W�=Xi�=�>��?΄u�_֭�0�Ͻ�B8��>.�`>Ӝ�>.�`������=�٭>�?_h)?�%�>�Mv>�;�g��C�־���+�2?��?�9?����_E��Y	�]���Z�=r��=^pN�~*j�p������{m�X=���>�>��>ut?&�o?��E?��;>0$ھv׎��`�+�&���$>N�?L��>xt�>���� FS��RR��,��
��W=��b�&i�=]��=��{�d]�>��>��=�4��$2�=�g���O�����>���>'�?0x]>U�=^|Q���$���I?���]_��ʠ��Qо�����>$�<>ym��?���g�}�����3=����>c�?���?d?�,D��(��\>}�V>S>�Z0<S�>�u�Lԅ��4>5��= hy�����Tݝ;%�\>��x>��ɽ��ʾA��S�G�ιݿ�p���`"������7F0�����	�Gm��ɡ���ޱ�<�پK޾��~>^m�=� ��"@׾��ʾb�t?El?�@Y���o��5�b�	���˽͎�>�����ݾ��3��=<7ٽ��m�hpb�	��K*���b���>/���Zy�4_z�U����=dwL>y�"?߆��Ȯ�՚ӾyS)>ى>6��5�쾺�������*�=��c?�8?-�پ�.	�@�#�J�4>))?�"�>b-L>g����D�R��>�.?��?6��=(���T����.�,>�?���?m�U?e�J��m��Q�������>�M?.��>�����2�i6'>�lQ?y?"(�=3U���������BV?H�?��L��8��j
?y�?�*�������K��_����*�fm?BQ��ݽ��]=��ɾ�,�%(x>��>����E�b��v�>{[��A(���/���p����o�>�	⾌�>�&�>�i>=�dŉ����_�T�4?)}�?=�d?M4?�9
�O�˾d�u=.H*>��>"��>^��I��<�x�>Q5�>�{��Q�yu�%��>�s�?��?G�*?;�k�k�������̺��B���=�-�=L�!>>��{�`=�l=��:���ܽ�@�<���>�{>��>��^>��1>ؾ1>�΄���"���������,E����Y����b�O���؃�	��bئ��a��X!F�@����>����!���#]��)�����=���>���>�>��4>��=�f�����ǽ߽������S4�[�������<k��;��Ŋ�U����e��(�3�>j'�=z^>�	?b���y̗;*K�>D�QD'>�h�==t�=�?F>�a���0>��R>�D>�+�=O�<�)�=�璿踇�a�o���%�U/2?�N�?�#��2�>z���c�83>�)$?!S8?�MM>W$�K8��o��媓>��+�������L->�">�c>�����g=�=u���,�i��C��>Z =%��<�Oּ�(�+ս��>"�����>���>ome?��?��>@݌���?�K�>sB�>Ͻ<���>i�>��|�t�?��?�&?���>��>7�`o>�*�<�����7�����K䅽���0;C������g>���Oz=��=e����>��=���>�f$?
�>�y�>.nn��'��=��[��i>�ս_}�>�?�Ӹ>/��>�t�>U<�=���׃Ӿ�	����>'Rd>�]��9����Y���>s"�>��^?�V!?^�������?+����>��>}�&?��:?���>���=��B������߿I��Q[ ��!��5���D&��Q��0�����<�"5�Ŵ>�>� ��z!>@v�>
q|>�II>-{>�+>�w�>��Z>�=L9[=?;J���>�W8�B�=�^��/��]��I�=㉵<}Ӽ�ټ<���c>��p��2 �G�?V�?��H=�ip���%���þ�)����>tT�>8��>	<? �>�qǾ!�_��_�5�־
�>0�r?rl'?�ir�#=�>Y�?�M��>ҭ>$�>>�>�����<����'#���2�>�B(?�^�>����H�M��1�����hU�>�F>ARѼ��?�%^?OF��V(�<U�&�FT�%֢��<�>�!>�H��Eu��~\��H��@�Y
߾i&�<�1�>�?yפ?��Ľ}'�<�������Ӄ���=�����!��=�3>?~��>����.�/�R�L��B�׾�S�P>�r�>;O>�=�>�o^?��H?��?#H?��1>�6̾�H$?���>��> ]�=�~�>�
?�S�>�	?��?�'>��
�	���\� ���C/���>}�>��>��=��=B`d<=5�yE,��&�=L�=;�>ͅ�=N��=p }>��a>7[�>�d�>�E��6/�m4��/�����>a�>�1�>���۾�wk�P�>)��>T8?j�?��>vn�
���G�=��#�1?��T?H�?뒉>Y�n�̿,�@����BI>���>2�`�c����վ���`�H��D�>���>�:h>u	�>	�x?5e?,�h?��=���n,��^X���>;�>�r?��>�^��^���D�J�F��2�������B=q���%g*��@�=�+�=ML�>�1>�ݜ=4-�=]���#�2���E.�?l>�B
?��@?�#�>�M>6	�/<�+�I?4;�����|���Ͼ/��T\>�P<>,L�_�?����}�����x)=�D��>���?���?Ed?�C�?�Ͽ\>�?V>�U>��(<��>�D���4��]>3>Y��=!�y��K����;�\>W�x>��ɽ��ʾ.��	�E��̿�{����W�Ǿ8K��7�<bǾT{m�|����'���"���p�dyc�,]�=�p��P�������"����w�?09�?��i�l��o�U��G0����?[���҅q����=r��x���R3��T$J�E=�cD�?x�>5���ㇿR�s�CY$�C񼽾>��$?Т�ɜ�����z>�'>����������g���eL�3�\?�Z:?O���I7���S�Խ�=T�>��>��q>I���v\�P؄>�}A?8b0?^{=�A��@������?7�?�[?��->.����i⛽>+�>Z��>	��>f�Ѿ�wھ:�>�aq?�9?�W7>�G?������Q��V?x�?Cz{�Ჟ=a�?�>1ӻ��<�b��-1��;��=6�>�@-=��W�u�X��>_��>}�.>~���U�3��>-N���L��/G��d���!���$<
T?���>f0n>ET>�4'��m���Ɋ��B��BJ?l�?Q�T?�>5?(���X��dt�����=�D�>6�>���=7��Ҟ>�q�>��
'q�l8�R�?"�?�&�?enT?�`p��3���4h��@��=e���=]�=Aq[>�[���&>kQ�8c�S���=j�8>A�>��>�jo>y�N>͙7>��>ӄ�������k��y�g�q�U�0��q<�Y��Ծ;�,�E��VR��������a=yBŽUW�U�����8�7���j�P��>،>�l�>��{<�i�$�b��t+��
��c0���	�*)������K���\Q��-�WÒ��7���fؽ@����?H��=y͝>�M?��:����m5�>�AZ>��@>p!N>ܛ=�6�=�½�%>��B>K��>���>7t����=�O��8h�<K��x�1�i�B>���?DJ�1�B��j�Ib�&�ݾ�<�>�I?�UC>hJ�k���W���v�>a�I�l=O׵=�9�=�k>�a>?3�=%����I>�%�=������܉6>4V�=��h<L�=�{q�����@?��о(��>=�?�s<?S�?�v?3�վ�/?� ?��a>l����>��>���=�w5?�aw?}T?'6�>��>�+z<��=n=��\g3���T��E�;+a�<W�ؽ��3�o�=�:k=a�Q=�r#>��>�U��4�����iO?�12?�-?G�?�O<��
��1��e���\>�^=�x�>���>��)?�8?T1�>�9�>r�w=,����ξ&�>Lv}>�0[��̍�������>.��>;�0?��?���W����=S�=�]?��?ϵ#?��>s�>S����,��`ۿÇ(�� ,�9~����`�kwQ��%#=�4L=���	'��?���
>(7G>2�U>��>X��=��>a�>{�'>���=It�=~ƞ���t<��
;�$=�>ۥ=���<-e=`�R>8=O�5��=��.��i�� !�=:p?�I?ª�<��Ӫ���Y���m�> r�=���>\,?��>1L*�Z�r�|�S��e��n#>ã�?L0?��z�.�v>r5O�`��It�>�0�>^7�>�7�=��x�p;��G�K��>�7?���>�h��3�y��7e�C�T��u�>vX�Q�$��*�?��,?�f���[��<�w�YH4��?��P=c4>�᳽$"���'���:�(p����ί��.>�L�>9ר?q~i�i���Δ��j��<��7P�EE)>��}����>W��>����������8�#������>KN?_�^>\4�>��V?��K?�~n?t�*?0�>�� �ɹ�>��>C˰>���>�-L?��?�4�>���>$�>��	=\������v%��0Mu�D>;��=��a>�>��>��g����=��=ɮ��)2@��J����E����={
 >�Q�;(�>��>U	?,����Ϙ<b�����W��2�/�>&-�bs�<x�
��"�E>?A�/?t��>��=;%��P}�a]�(j���?�w9?�I?P`i=𨣽�������->�z�>�ӽ�ޒ^�������4����Wx><ʳ>�J>r8n>�|?�J;?��?�E��.���w���$�����T��<�o�>��>���=�9�)@B���z���Y������;G�X�N�=S�>qm�=�h>�
>���=�����:��˽�{��{ҽ���>Z*�>{X	?��>v�=�7ƾ�I�W�I?육�b��⠾_bоʻ��>�<>��<�?S��L�}�(��&B=�u��>&��?���?�<d?��C�$�%�\>;QV>-
>c/<7�>����{��*�3>j�=�ry�z����;�]>$<y>��ɽW�ʾw,�c�H��6����H��%ʾp���AӾE� �r~ܾV�=佽h��������e����*#1��9=��ӎξ�K�@ٯ���-?*�Y?2���<1��`�pci�y����o�>4����ؾ�i����ӽ�|��"����m=�>��I�j���r�Q�)�x�=e�R����sɀ��� ��U�~V=��'? ���*ܾS<�;y>�6Y<�~9�����٧~��S��o��E�$?��$?MHо��¾��Z��>6#?_K�>������7G�,��>��C?5�?ͰD� Z�����S�>?z�?*�?	/?�`�>ϒ,�.��?��x>�N2?�W�>N.��ה�Vq>��u?<>�>t7��`~�	a����2�n�Q?�?�L9�@K�_��>���>�?����X�~�G;��C�H>���>�m0�9*+��U�d����f=ƞ�>���>^��\�����Z>����&��D�y�6�\ ���M�=��>C�<�ؽ�k�>E�=s��x�Ov��r�U� �0?���?�+?35z?���>���iL���mE�D?8�>7��M� �~j2?��L?Iyվ�o^�����,?���?� @��o?�z^�Gӿ������V�����=&�=��>>�޽�̭=S�K=����|Z=��>b��>4o>�;x>��T>��<>-�.>&���>�#�qʤ��ؒ��[B� �����vg��{	��y����ɴ���ϔ��0����ѓ�o�G����CP>��E���'1>���>t'>�]�>i��>L+>[{��?jȾ�x|��mB�nn��E'��+�q�$�zN����*��k����Q&��8E��5.?� >�}�=��>�㣾4��>:�7>{�=T� � �?�c�>!�>�0>��G����>]��>�Kl��nW>�_>�~��ڲe���Ҿ�/K��{>9I?�򭾞m������YI��q0�>7��>̋�=>�N������u6�?6I>ȧ�<�L�ʘ"�r�(�;�n>��D>}D*>t=>_�r�O�̾(��]��<�`}>��S>~Kj=�hԽ����Z��M�>;.��|N>�[M>)n?�k?Z��>Z�4>���>��>ȁ\>�f>�*>���>Ra�>d?�`C?Gr#?��>0�>?�%�>�>o�b�R>e�o�9��@��p퀼��p=5��/�>��L>�ſ;r�K�ɺt�u��K�-�A=i�? "?0��>�a�>oiD>)��֥<�۹�<Mɓ>:dR>�>%��>�v ?է?ځ�>�J?>�{W>�g��&����>5aG>޺���܌��妾����z�>GK?K_?��j�{�ս2�����8M�=5?;7>?7�>`�y>���7)����7�(��8��9u�����ǧ:L���N.ѽ�����N��GM��R�=�2�>��>2+s>�A>s�=
�>� �>�K> ��H�>�3i=2���z��xc=O���P��=���fl�"Y۽�
���5�@�#Q*=܎��h��I?v�?�ݮ���ýjqo��r��cE���O�>o(�>+�>,�>p'=��A�P�t+�+�
��?�ii?���>�V����='z��=$�ƌ�>��>��=�Q���S)��i���؉<L��>`D?���>����NQ�F?c�Z��ڵ�>��=_�F�'�?A�m?ð��ZȽw�D�(B�s���d->b�1����<2�?�(��%��R������J ��w��"F�>���?��0��|�>Q�_��쥿f�z�-/�d)'=��C����>�=�ԓ��� ��0�&�����j֤�j
�>0�f>�7�>%a9?H\-?�Qf?`?:�#>�\=U�P?,�>

�<�#?W�?�#?�d�>��>Fs�>�>[ാ!Pd�����oW�� =�R;>�3>T�A>�����e�<,b/>�k��>=u�j>Ub�=@+J���.��v�s�$=p�=F�?�;?�מ�m�:��R=�-��� >��?`&?ʝǽ�H��V��&=�ڰ>.>?G�?��U>�\3�>�����5�@���? �?c^�>گ��V}۽�]ؾ�����½!@>٫�>�)���_���c���z
�	~=�ձ>r1>b�|>w-�?a��?�x?�=>G�e�������F>}ҁ=�6�>�M5? �Z=���q�
���E�U�H����Q}�7��RV�@�=��s<�͍>�U>��j>��>y���V��C<�w�=� ?��
?���>�9z=0�=N�S�6Ⱦ�N?�#���ȾLm%��o]����>W�U>HR�����C9?ʘ�>5H�j#���|y���[?���?̓�?���>)�ר���t>���>$��;��=�ȑ��ụ��r��>�Q>R�c�����U����=��K>�Q���׾'t�%��<nH�(���%ﰾlzվ�Ly����F┾�.�.ξ bP��)�o6���mK�6Nc;T;E��j@�J����۾�]��$��?VR�?l���7 �>���Fgk��婾a�>�8Ҿ�w���,]ӾP^�����'34�O7:��nB�B�(�ZW,�{��_������E���	����T�T>�C? ���2������oV���F>�p� A�*j��)���&c�Y�i?�*@?Ynξ{�l��Ò�0[���?�ײ>"v�����b�E>Y��>���>+h ?�����g�،z���=S�?�s�?���>@����E���;��?e�8E8>�CY?u��>�0A�$"<��Oѽ
o��O?���>�1K�{����H�ً?T��?��Z���0>$�r=�Dg>�^>t��	��5��;�z�=�<��+ͽ�,�<�x0�Nѽ�q]>���>.А��/���f����*��(��$�G�!�"�S��>��0?��(�MX%��y�>�گ>�难�Ek������7��"f?�?�a?'�?^vҾ
�;i������>h�t>&�>�t�<����`>��>��z���M�_q���"�>iG�?�!�?�+F?��8�u'��Ox�9����J�/��=�)=L4>tc=���=N��d�=�>��>㪛>{� >��>'�=>��>>Wv#>"��Q�!�F�ѿز��Z�U���/�dq��Nݽd*a��#L�m���M�����dK�*�����p�����ak=*�D=ʚ�Vx>O�>�J>�K�>�K�>ۣ$=��ļ�I1��	��a��2<׾+�%��U�r��z��C�l���|Ⱦ�,?�gn�G�?�ཇu�9�?�
{��>6��<�pݽQ�6=µ�>���>o�>\d>[�j<��>?x�>/�����i>�W=}����G����4�][V��x=��F?Jau�6Q����*�0�Ӿᢾ1r�>j�?��G>L����|�s�e�>p�V���S�ʠνHM��[
�>>FS�=Z��;-}���yr��U���!�=��>��>t@��꠾�6
�|b�=�,�>��������n�!���%?�2?7?�|>RL��L3>J�>��3>��9>����R�e>��(?p%L?��&?���>�]C>�7��>A>H���;�6�w��=�u�*~t����,Y�>D���R��4p�˝�=N�> �S>j������m3�<��>;�8?+V�>���>� 1�)�<��J�}��6>�'(�Ԧ�>7o�>�-?��>"�>��->a�ٲľ�d�g��>�.B>� [�m�q��|���o>2�~>��O?��,?����^Q�7=�j�=꟭>��?��+?�I�>+!>c>ý�����п�*��%�����#��B.=���m���������5���q=�l/> �[>��r>�ww>[DC>�(>�4�>oK> ��=�=�s<��<@�Ԣ+=���U�<����,�B��v��@��B]w�-ؼv���h˼|����>`��>�R �q!6�H�?�l����
���>~�g>�8�>���>wr >��;͈E���A�kpa�s�?o�h?���>WW齳b�=�Ɣ�|�<^Z>\��>��=�i���i���ut��TźҠ�>f�)?4��>�xн2�c�$Ȃ�¤�c��>e�0�A��=vi�?��y?�d+��
��PD��zB��j��̀������K�{� K�ۅ��
�����yؾ�T3�	�>n¯?�w��N�>�ޮ�^}���-h�D,�
�D=˕p;��?�>���E�ɾ�?���t'u��5X����>�H�=���>Ǵ?g?Ǔa?��?��?(��(?�ư=���>{H�>��?4�
?Y��>�w>� x>��%=���h	��`���$<L彼	S�=��>�)>,�<`\#=�4/=��<V�;��:ƼC��<+.*<�|=�ލ=���=�4>�?P!'?K�U��4ȼ���H��UM7=
!'=�ܐ>��=���ԑ��ɟ=x��>b:?�k?W�H=��9ʾ�*�n�/>~n ?i�?(�?�k�=�E�R ��b�G�ϙ�=��>|�ѽ��~�K6���.�b�q��?>�\>n�;Up���x�?��?�Ӂ?�����V*��d����zS�>^�8�V�s>}x?1��< ����=��,V�jG���3���[���<8kw=��>���>8L�=�e>e�R>��<j7 �2��=��>&�?D��>�*�>���=0�g=hA�B�޾�?ϼ���"��\��h���Gi�>��$>F辞dԽo�M?��=RꗿY������=��h?���?l�?;��>jdƾ�߽9I�>Z�5>���>]6�A���Qr=�`�<���>���=�x�ovb���2��H=xk�=�%���&���C��2 >m2����G�q��5Ǿ���wGY���ݾw�6�Ȑ�Ί������u����S����������>����fȋ?]
�?-RJ>Z��=@�1�66��ʾ��;�|�u�q ���r]��)��ľ[¾����L 2�76�
��g>�-��]y��A{��B,�9Ľ���>�/;?�޾E�I�����`.�=mo�>§�<u���K��ԋ�m�O<qSV?}$3?�6辗�־W߻�ڄq="?�+>A�޼��	�,���VS>�c�>-�A?<T%<NXz���� >���c�?��?)?ɛ��!������Ͼ�)�>Vޜ>v�$>1lt�$վ1���(�=&Ik?�m�>�^� ��ԕa�\?��?6#=��I>�u>'�=܂c��'�7X&=ڹ��#����_�P��=�W`��1(�

��,�>�_�>�T�>9�C��]���>�G���_�q�U���%�Z��ൣ>z4�>7d:��;�>���>���;~���R���x����V?*�?�gS?��"?]�Ӿw]ʾ��a��|>�?�>'��>�L�LZ���Y�>��X>�9��^W������?۶�?���?��?@E�]Gӿ
����� ����=�%�=e�>>��޽lɭ=��K='Ș�U=���>{��>o>;x>F�T>��<>6�.>_���}�#��ʤ�5ْ�\B�� �֤��vg��{	��y�����ȴ���C���㢷�Г���G�_���S>��蜾t�>?��>�һ>!}?do�>Y�>ʱ��W�Q�b�þ� �fs�#ľČ��H������s�W��q[m�1���rdA��+?ٓ<{���L�?_ɟ���;�?8�&�X�=��>*�b=>YU>��/=�?�=1�)>A��=M���7�>�aJ�m���2
a�d��>��A+=�Y�>�y|��{<-�4]������:�>��?,�>���u���i����>�9���=���^��׆�}d�>�C�>��>M�C>6��<����7ͽ�Bk>)�>��=W�ǽUA¾��Ͻ�>Mѽ>h�������6��t�>"
?� ?Q��/G�Ѱ�>AZ�>���<��=��Y�������?��e?B�G?1l>>JA�=�A+��a��=Z>��4�t t=����H�<�c���/5���=b�P���=���>7d	<2��$�����=�-4��7�>�qP?L�>DW?��
��ZD���o��R�{��>�����	�>M��>[_> M�>���>dOJ>��#��k�й���F�>$ɓ>��R�/̆��^�=��=�U�>��n?,�?�=�5%��l>>��o�<>DT�>��?�:�>,pX>��p��0�?ӿ��$�B�"��r��Fl��H!<!B�%�c��o<�.�%���LP�<�U>;ރ>��x>)J>�$>M�8>��>4�F>J��=�"�=��z;�,�;? H��.>=����Ax<C>J��w��s�Լ-������C9�^����p�ݼ���>�e&?�Í=�6'��P�����L����?6V�>])>��>�#'>č4�O�2��-���B�Ny?�d?���>��d���=��<�>�=a�x>
4�>z38>?�ͽ��{��<A�O�%=��>��?]x>�$��,�}�C>��p���6>�~�=e��D�?��P?����q��eJ����FX%��֯�b�¾&��e��+����� ��� ����᳾\4�>u�>7̤?�6��{>�y��y������� �׾w���22={�
?�?�=ᵈ�=�m�|���[���=�d�>An�>����#��>�hT?�I?r��?	�'?��>���>�H?�S�=H?� $?�?Z��>���>����1�=���"Ƌ��o^�B��v6���V1>��">F9S>��>�=��D=��k�ϵ
�Mh��n=�{����<d��;+�x=�?�>�d>E�>��?[ϣ��0h��F���U�l�N>!1�=�X�=�?����#��*�B>|s�>$R4?B~�>�얽?��>ơ��>E�yQ�>�A?��%?��'?*��=�yy�1G������8�od�>W�����NP(�s1澧��\�y>q?>v�'���?=���?{�?u�s?SE�@b𾫳��v]����>��޽DZ�>J�)?ҁ��b䷾Ww ��ڏ���Q��d�U������7н>,/>u_$==3G>�B�>�7>���={��=>A> ��=d��=���>�_�>Om�>��
>�s��d�Ⱦ�C��c@)? ���D6�x��������{�>�~��뵾��?g� �o�D�nꂿDY+��د>Q{�?��?D/?�U;�0G�=�5>>�Y>,��<��c=�H'�3�p���y��g�>ZoX>�fO��h���x�����>�^)?�*~=�����I�=;��<�.�������������2��Sl���������?���53���걽v��$��Wi�* ��X4���a����?��%?�ܾaKϽ7_�}@A����پ�>s���>d|�������Hӑ��{��O��@�!�K���!�@���>/]���a���"T�1���]�<o6l>e?·��p�G�s"���\��A�>�>�V���j�����";����f?�9@?]�;C��A���D�m�>�f?`��>9`�Gˆ�g���!kC?>b^?8½d���p/{��g̽�?y�?��R?�%��J�;�H���ZLw�D�?R"?���>eu�Q���1��"7�>5Tu?��?m���)�_����� ?��P?,��9�>��?�Ku=I ��O䇾I�׼�?��/�o���M����%=�`�鹾�?>4�>s/3>�ـ�W/H���Z>����&��D�y�6�\ ���M�=��>C�<�ؽ�k�>E�=s��x�Ov��r�U� �0?���?�+?35z?���>���iL���mE�D?8�>7��M� �~j2?��L?Iyվ�o^�����,?���?� @��o?�z^�Gӿ������V�����=&�=��>>�޽�̭=S�K=����|Z=��>b��>4o>�;x>��T>��<>-�.>&���>�#�qʤ��ؒ��[B� �����vg��{	��y����ɴ���ϔ��0����ѓ�o�G����CP>��E���'1>���>t'>�]�>i��>L+>[{��?jȾ�x|��mB�nn��E'��+�q�$�zN����*��k����Q&��8E��5.?� >�}�=��>�㣾4��>:�7>{�=T� � �?�c�>!�>�0>��G����>]��>�Kl��nW>�_>�~��ڲe���Ҿ�/K��{>9I?�򭾞m������YI��q0�>7��>̋�=>�N������u6�?6I>ȧ�<�L�ʘ"�r�(�;�n>��D>}D*>t=>_�r�O�̾(��]��<�`}>��S>~Kj=�hԽ����Z��M�>;.��|N>�[M>)n?�k?Z��>Z�4>���>��>ȁ\>�f>�*>���>Ra�>d?�`C?Gr#?��>0�>?�%�>�>o�b�R>e�o�9��@��p퀼��p=5��/�>��L>�ſ;r�K�ɺt�u��K�-�A=i�? "?0��>�a�>oiD>)��֥<�۹�<Mɓ>:dR>�>%��>�v ?է?ځ�>�J?>�{W>�g��&����>5aG>޺���܌��妾����z�>GK?K_?��j�{�ս2�����8M�=5?;7>?7�>`�y>���7)����7�(��8��9u�����ǧ:L���N.ѽ�����N��GM��R�=�2�>��>2+s>�A>s�=
�>� �>�K> ��H�>�3i=2���z��xc=O���P��=���fl�"Y۽�
���5�@�#Q*=܎��h��I?v�?�ݮ���ýjqo��r��cE���O�>o(�>+�>,�>p'=��A�P�t+�+�
��?�ii?���>�V����='z��=$�ƌ�>��>��=�Q���S)��i���؉<L��>`D?���>����NQ�F?c�Z��ڵ�>��=_�F�'�?A�m?ð��ZȽw�D�(B�s���d->b�1����<2�?�(��%��R������J ��w��"F�>���?��0��|�>Q�_��쥿f�z�-/�d)'=��C����>�=�ԓ��� ��0�&�����j֤�j
�>0�f>�7�>%a9?H\-?�Qf?`?:�#>�\=U�P?,�>

�<�#?W�?�#?�d�>��>Fs�>�>[ാ!Pd�����oW�� =�R;>�3>T�A>�����e�<,b/>�k��>=u�j>Ub�=@+J���.��v�s�$=p�=F�?�;?�מ�m�:��R=�-��� >��?`&?ʝǽ�H��V��&=�ڰ>.>?G�?��U>�\3�>�����5�@���? �?c^�>گ��V}۽�]ؾ�����½!@>٫�>�)���_���c���z
�	~=�ձ>r1>b�|>w-�?a��?�x?�=>G�e�������F>}ҁ=�6�>�M5? �Z=���q�
���E�U�H����Q}�7��RV�@�=��s<�͍>�U>��j>��>y���V��C<�w�=� ?��
?���>�9z=0�=N�S�6Ⱦ�N?�#���ȾLm%��o]����>W�U>HR�����C9?ʘ�>5H�j#���|y���[?���?̓�?���>)�ר���t>���>$��;��=�ȑ��ụ��r��>�Q>R�c�����U����=��K>�Q���׾'t�%��<nH�(���%ﰾlzվ�Ly����F┾�.�.ξ bP��)�o6���mK�6Nc;T;E��j@�J����۾�]��$��?VR�?l���7 �>���Fgk��婾a�>�8Ҿ�w���,]ӾP^�����'34�O7:��nB�B�(�ZW,�{��_������E���	����T�T>�C? ���2������oV���F>�p� A�*j��)���&c�Y�i?�*@?Ynξ{�l��Ò�0[���?�ײ>"v�����b�E>Y��>���>+h ?�����g�،z���=S�?�s�?���>@����E���;��?e�8E8>�CY?u��>�0A�$"<��Oѽ
o��O?���>�1K�{����H�ً?T��?��Z���0>$�r=�Dg>�^>t��	��5��;�z�=�<��+ͽ�,�<�x0�Nѽ�q]>���>.А��/���f����*��(��$�G�!�"�S��>��0?��(�MX%��y�>�گ>�难�Ek������7��"f?�?�a?'�?^vҾ
�;i������>h�t>&�>�t�<����`>��>��z���M�_q���"�>iG�?�!�?�+F?��8�u'��Ox�9����J�/��=�)=L4>tc=���=N��d�=�>��>㪛>{� >��>'�=>��>>Wv#>"��Q�!�F�ѿز��Z�U���/�dq��Nݽd*a��#L�m���M�����dK�*�����p�����ak=*�D=ʚ�Vx>O�>�J>�K�>�K�>ۣ$=��ļ�I1��	��a��2<׾+�%��U�r��z��C�l���|Ⱦ�,?�gn�G�?�ཇu�9�?�
{��>6��<�pݽQ�6=µ�>���>o�>\d>[�j<��>?x�>/�����i>�W=}����G����4�][V��x=��F?Jau�6Q����*�0�Ӿᢾ1r�>j�?��G>L����|�s�e�>p�V���S�ʠνHM��[
�>>FS�=Z��;-}���yr��U���!�=��>��>t@��꠾�6
�|b�=�,�>��������n�!���%?�2?7?�|>RL��L3>J�>��3>��9>����R�e>��(?p%L?��&?���>�]C>�7��>A>H���;�6�w��=�u�*~t����,Y�>D���R��4p�˝�=N�> �S>j������m3�<��>;�8?+V�>���>� 1�)�<��J�}��6>�'(�Ԧ�>7o�>�-?��>"�>��->a�ٲľ�d�g��>�.B>� [�m�q��|���o>2�~>��O?��,?����^Q�7=�j�=꟭>��?��+?�I�>+!>c>ý�����п�*��%�����#��B.=���m���������5���q=�l/> �[>��r>�ww>[DC>�(>�4�>oK> ��=�=�s<��<@�Ԣ+=���U�<����,�B��v��@��B]w�-ؼv���h˼|����>`��>�R �q!6�H�?�l����
���>~�g>�8�>���>wr >��;͈E���A�kpa�s�?o�h?���>WW齳b�=�Ɣ�|�<^Z>\��>��=�i���i���ut��TźҠ�>f�)?4��>�xн2�c�$Ȃ�¤�c��>e�0�A��=vi�?��y?�d+��
��PD��zB��j��̀������K�{� K�ۅ��
�����yؾ�T3�	�>n¯?�w��N�>�ޮ�^}���-h�D,�
�D=˕p;��?�>���E�ɾ�?���t'u��5X����>�H�=���>Ǵ?g?Ǔa?��?��?(��(?�ư=���>{H�>��?4�
?Y��>�w>� x>��%=���h	��`���$<L彼	S�=��>�)>,�<`\#=�4/=��<V�;��:ƼC��<+.*<�|=�ލ=���=�4>�?P!'?K�U��4ȼ���H��UM7=
!'=�ܐ>��=���ԑ��ɟ=x��>b:?�k?W�H=��9ʾ�*�n�/>~n ?i�?(�?�k�=�E�R ��b�G�ϙ�=��>|�ѽ��~�K6���.�b�q��?>�\>n�;Up���x�?��?�Ӂ?�����V*��d����zS�>^�8�V�s>}x?1��< ����=��,V�jG���3���[���<8kw=��>���>8L�=�e>e�R>��<j7 �2��=��>&�?D��>�*�>���=0�g=hA�B�޾�?ϼ���"��\��h���Gi�>��$>F辞dԽo�M?��=RꗿY������=��h?���?l�?;��>jdƾ�߽9I�>Z�5>���>]6�A���Qr=�`�<���>���=�x�ovb���2��H=xk�=�%���&���C��2 >m2����G�q��5Ǿ���wGY���ݾw�6�Ȑ�Ί������u����S����������>����fȋ?]
�?-RJ>Z��=@�1�66��ʾ��;�|�u�q ���r]��)��ľ[¾����L 2�76�
��g>�-��]y��A{��B,�9Ľ���>�/;?�޾E�I�����`.�=mo�>§�<u���K��ԋ�m�O<qSV?}$3?�6辗�־W߻�ڄq="?�+>A�޼��	�,���VS>�c�>-�A?<T%<NXz���� >���c�?��?)?ɛ��!������Ͼ�)�>Vޜ>v�$>1lt�$վ1���(�=&Ik?�m�>�^� ��ԕa�\?��?6#=��I>�u>'�=܂c��'�7X&=ڹ��#����_�P��=�W`��1(�

��,�>�_�>�T�>9�C��]���
=�%׾Υ^�i�=��3� v�����G��>�o#�U�c�S�>�I
��6�JA~�*~��A޽�?�+�?^?"Za?BG;�sC
��+�y�-> �?�9�>�}2=�.A�tQ�>o��>d|�9b�Zþ�W?���?���?زN?D�y���Կ�N��o���������=��=��;>�Nཝ~�=�GJ=�Ҕ�h_H�|�>�ٚ>�p>��w>��V>�e>>4�0>{+����#�R���㑿>�A�E\���o}f�	�]]v�Q������!�s줽aز�e_��%QG�z��'5�p>����>�Qi?4�>�ܼ��Z��/>������\�7=7�>����/��2,�c���=c�>IS^>`c��xX�[s���}��,?<���!<5�>����4U=�.>� <f�=)M��+=�̼���='�>I1�=�j+>� >�h>w�ֽ4y���Î��W.�n}���HH>�7?�+�<>���i� ��u4�0�[>�X+?�S�>yT��vy��kV���?�_!�u���ͽBY�>9֬>/�>�d>�8>@��;����%�b��>�:?���>��M��������>+�>K�����=>�W�> 1&?��q?7�b?ջǼ�I[>v��>M]�>oI7>7/>7�=��z=�?XT�>�)�>E��>)�=#�+8�=���X���r��*���Z��X�����<���X� >&��=~���>�=>B{��oM��>=�A�>&]?�s�>��?!��H��0u��;�'�:���Z�>&�>5G7>_��>`�?*�>ܱ��b�N�xT��<�>1��<�7��`�_�ac����3?@*H>nFw?��5?�t�=Ծ����YJ����>�*?l��>�B�>���=�K7>���yԿ� ���A���8���=@�i<DnU��᤽���<�
�����}<�PB>�H�>�8Z>1Ff>� m>Xx>�l�>�S1>�^%��i:>b/?�xڤ���=f�!<R��n=����,��j�=��0���۽(�ҽ(���qü�ג<���>�f?���=$�P�ܻ>���^�#��>��B?��/?�p�>cuR�gWM���|�`fX���n:��v?9t`?@>,�����A>Y�>�=�S�>����;�>Aξ�ɽ�yE��|�=s��>�,�>� >�i��KGN�.�S���9�]yU>��=&8=ႝ?�1?���X!���W۾qm��!TN�ц�>F�>栔>wp8��XA�s�����=l���!���)�=ݖ�>��?r�yc�>b澗G���=��骞����@��=�5�>j��>	��=��>�/��J�콼�*��= ��=��>>�`���>y��>��l?�s*?�!?��>��?��&>�D=P��=�>m�=?�H�>N*���w��F+>��>[S��Ž��=5xl�M�ں�g&>��=W�'>؄�$*�����=�)J=A�><�z2�	`+��?0=�*0=A3�=fp�L��>��3?�S=��]>�T�b<��؛#<�:�=��=��.����8����"=s%�>Io?��>uv>k���Pӗ�K 1��6�=ܦ?U_?yD�>������>{��ϼ��>�V>_Q�ʚѾf1��þ��z>���>���=�o�==b>�с?Ħ+?\.?�U��*��ny����8�;��D��>�>(ń>.I�<�����n�.X�����r="mD��Ou=E>���=���=�d�=�6>�a����A�����Y�Z�ݽ��>��>��?&�>&�=��˾acݾ��$?���iE��*�8þ!e	�f�*��Q�>��=�A%?�S�5����p���B���>^��?��?��(?ގ��H��]�8>���a�M;��>����sk�=Ww5�܌�>��>�D��k8�#�k<�>mԀ=m��Y�9�󪬾�Ҿ����P >�w�,��e3�q�������2�������7�m ���߾\9��u�V���6�a�(��뎾>ᾨ���ӱ��0��?��?��-�|�&�Y�t�g#�ޢ��_>�D���E���t8��tk����Ӿ��ﾄM���d��I�4��U�=Ds��F���䋿M����3=p�]>�H?7����˾�КP��j�=��>!����Y���������0?�F/?Tp��t��E��=�Х>��>�b��;>���BX ��S�>� G?�":?��/>bז�����$_�<���?`��?T�(?p����4�P
�"+�>�VK?a��>
�?H�,�!CA��?����?���?~]+?4�ݾ�Jq����?�!+>\@��5=.�>�mb>�&W�佽�vt=^ꄾ���=���>�4=ⷀ�,�v��v����>�">ކu��S����(>�㾽։�~�M�m=����á}�7�?�	�����>%�> ��<�~��-���Nx�{�I���2?�'�?�K?�3?Ճ��\���:��7z���U�>n�h>P5�>����H
>���>���kF��d��c<G?lb�?9��?>S?��a�h��B������-����="ӓ=I,S>�?���_<5�=2^��ۚ��'1�=�ń>�ӈ>N�>�Y>v��=�7>����� +�A:���ƃ�ƣ?���/��W"K����R�����Ѿ��׋�rGK��E=��m��䠽"�G��S<�%�.�K?�{A?
 �>�&?fC��<R�>����Q*���c�2'վds7�2XC�i��u7'�-y���>�����>�2��ܳ��t9?S�5���'>�n>�'��ѽ�:>����=
��=��r>�/�=�&=.�=�m#�����%�{��9_>%]�4	����s���<��;�=�ýC}�>����[��Mg��"�B��ӹ�6��>��>��4׊���7�ex�>����kn�+D�ǁ�=n>���>���{5�ƌ!��f���}=~_<>�@?V�>�)6� ��˙>�C��=�;�>02 �&DW=���>hq�>H?(�?N�!@�=��s>� �>u��>���>�瀺�)����!?s2?�>j\�=���=6;C�N��� SV��`ӽ���=���@�~�-�<�<�>"V �3�">V���[r��/>Z�P>�_c���<�~S>ذ�>���>� �>0�>L�쾒k:��Z���Z�V>>鈘;\�?��>$	�>Y�u>�G�<��w>��~>Z��&���rB�>���<�fI��b5�:��y�?!��>�n.?��?f�(��&;=x�C玼]J�>�>97h>`Q�>�>�C�������Կ���uh!�vZ��_�!��.�<��?�[h,����<��P�(���ۮ<MV>[ו>��z>�
`>� >8�:>�>�>)�=2�3=#f�<dȻ��;�x��=�U�<jǭ:m[N��I]��E��k�a��]�=��A�u�<v�ۼ�?��>���=�F.�����S�w=���H!=- ?�(?�]?�/>�x
�]�(�����V��4�>�Q$?�S�>h����>�6�  ��a�>���>Æ�>.��=C���j����(�z*�>s3�>x�>�1޽2�H���3�=��oy>��~=7��v?�	?q�оS�����K�(`���Ǿ|J>:�z>[�_>����"�l�e*<
�¾N%־�K�= 2�>�:�?�eH�8��>_��g����Wt�V/��a~=>A�H=�h?��>�|>1���5	��b����Խ��<���=�(>��=��?�()?.2�>�6??�O?)j�d��'�<	֔>l9�>B???��?S��>�c��>�M�=o8��L����X���=3��=F�>E� >��=�q>q.�=�c>=���Lb-�t �;�������X<Alk=mI�>9�=NJ�>#�?w�C�I��>��D���P�L[y���>��N>���=s�,��W0��5����>�?\��>��>6���!��N�Tƿ>��	?�v?�S	>��>y���\�2�9>mEG>v >��ۨ�m&[��ןm>eU�>���=7>u�k?BY?R_�>>P��3�h�%@��2PQ�Ps>e��>�?�t�>��H�H�.����a1���[�M�/H+>K��Z�1>E�=�
���#>�(K=�@@=c2>\��U]˾���Ɛ�e��>9��>q*�>��>y�(>+]���mؾJ�5?�i���'�C����� g;C[v=fbO>�`�\�>���Ѫl�6����C��#�>1�?�2�?��R?�e������[>�Ca>�=ς�<��4�э�<���</>�/M��^��K�@c=$:�>���>{':���ɾ�:��fF�T�տ�_D��?�(��W�^�_�������t����b�����¾�q��*���hF㽐�8��N*� ���c^u��s���? J�?�;�M�k�:U��ݾ_~�=<Xq���=�$U�w	U��q�U�վ�E��/�\>��x������e�>�U���n������E��KI>��?j�??:Q#�����|D�
�=���e>�0�>-�s���|��j��_�=��0?w�O?�~4�v�從]�<�l?�@�>�I�> X>�ĺ�9�W�]VZ>gbF?��-?��{>�c���e��饾{m�?�{�?Es;?�*Ҿ��$�d�����>�?:S ?��?�H�o�+�~nҾĦd>��9?��@?����C[�ṋ�t�?j�>� ��q>�4�=ͱ�>w���҅��_��!�ڽb!�u��>�	�>����:6ƾ�Ci��6>�+�>�>q��$	���u>9��J����q�HvI���>1(����H?I(�+E-<�kR>�"�=�2Q��]��ފ�"���B?���?,zd?�WM?��^Q	�H"H�G�@�>7�}>�^>���G�b>��>������ʨ��A?�5�?B�?�D?D�b���Կ&Ř�>v��L켾���=��=��K>N�ǽi��=��T=t�a�^Ѡ��V >�&�>�A~>6Nt>K<W>R�D>�.>΂�z�"�f���)���5@����[>���b�/�u7k�P$��/���ܷ�L��`諾N�u�Ǽ<���F�!�]�A��D?��#?�6?ߒ>�J�=�5T>��^��[�K��� � ��c�T��"��P�T���6�G=�R��Y���ž��?T�
��=\D�>��ʻڶ*>��>�1!����=;L>էc��!�<�㳽Qӄ�hj�<����0����>pb὎�m�FLv��j޾큽��7��Z?�|�'a#��r�����̾�5>�^?�Ui>.�.�;ŀ�z��=C�>�ˁ��=�١8�U�>���>���>�Y޻�:�=`�;�ܔ��6�,��=�fV>\��=ę��x��T̎�&�>%��>�(о����ν�L?��?��	?���<'X=6��<��>���>ԣ`>G; �����1;?��>/�=LԀ>�^�<E"����&��A=i���"���י�m�=�Ͳ�;�p���u���,=���=�Ө>��ה����?>�U>��i��+�>�|?F?��>��e���B��N,��ཚf�>{f�<�5�>)�>��d>��>%��>yX>�#�6�Ͼ�W���+ ?��O=�Ն��Hz�Rv�=}�?^G�>}�)?���>K">�����w��m�=�� =�c�>�(?��'>�_�<�ȝ�W�
��lÿr��MA.����L��<~f=|/���]<�mo< �G�Ȫ�!۾;��r>ᇥ>g�j> pb>��D>��->\��>&>���4,�=�<<�4��̛�Y�.=��6���N=�A �ŀ�<X9���p��Wd���S���<���ϼ�ٓ�l8�>�]�>��=��_�[�=��j���>�ba?�Yx?��>nK��w��&��5�꾰��Hf�>·�?>vs>蘾3�b>�E�<	��T=�(�=�T��*vӽd������㷨=�	?]a?���;��Y=���^$(����B��>�<�=~k�q-�?;�2?<�2�酨��8+��@L��g���pc>a�=�O�=oy<���ZL�!���,׾�r����=)K ?꿆?�r��%h!>�쾾+�{�P���!�оu5�=�{0>V�O?"G�>�?�	��OF��>���������?	�>s1=�q>q?�gD?��z>��>D�i�E�>Yi��N��>�!?=\?��P>�.��=�>�C�>%�x�� �*��$T �*uڽ�o7=?�_=>_�=�2�=�$7>���=�߽a4�/z9��">��=,ĽZ� =�H=;V >��=%=�>B�>����'�=Yz�=/Gk�,��Pa*�����߁=����EM�=�r>���=`;�>c��>�Q�݆��7��=A���>K�>�$?�8s>=[`>72��n��St>�SH�N֜��J�5�i�7ڽ=MR='�>$nB>hQ�=]{>f�g?�,d?�.?y�L�Q��Vy�M)(�X�>>��>�R?Sy�>6[�#����ŧ��E��ui���"���>�0�P�V=)s<]m=�Ĭ>��۹)�>�F�=ǧ�=ו��-�=�S輻:>"�>�?�U$>۸�<�.�����2� ?O���^y���X6⾁
�<����?��Q��>�G�#x��)��7����?j�?7��?�7?$NJ�.R��mɃ���Z>ds�>~.�>2<���>׉=�*�>=})>Uuݾ�Ó���>�?���>�Fӻ+��ÕN�x}�r�߿a�C��;ν�h�y?k�DƟ��GԾ��v<m>��Y��:(��P�=�2i��/ܽ�a��tt�xg9��CP���m�T@�?�ք?kIc�B\���N$��`ӾG\����>t�}������s&�<ݦ9Y���֧�!��\�۠,��eƾz�����>KTԾ����a�c�������d4>E�[?�>���ʾfd��^����=��>�Oʽ�<��ޅ���ʤ��>0?�(J?�m+�� s�X쑽$ӽA*	?��?&�5�j*ھ.������>L2_?}�X? }>w"��[7��ޤ�%�?�h�?շ+?V�þL�����_�>�Ӌ>|0?���>g�������֗�εO>��=?>�?R'ݾ�O��~#�V�>�=<�(�=HL>�ݏ>��T>9���t0H��lp��ѾF�3�>eC��� ���Žը�G�(>kQ>
CF=��;Ԫ9=���>!�.�N���H�s��;��6��<�t?���Y>��h>&>�i(�a��������9}L? _�?pS?�`8?1���2Oﾛ����=�=wŦ>\��>�í=N|�/�>0�>����pr���\�?�%�?%w�?�AZ?�wm�$����و�!
��
�ɾa�>���=�o	>��[w�=5n=�j�<:i��9Lx=h�>�{�>��P>�{,>59>5�2>(�z���,��캿"���LR1����?�Ex��-P*�х@�:��,�"����9J���=�2�<C��>g}�K@F��p)����>�Ȅ>�� ?S��=o >t�U>yϣ��l��s��F���J��̠��<������-���=/��h!��Q���qL��["?�� ��>���>����'>���>�e�=	B>
�*/=��#��� ����A켇�+=��=�i�<�r¾Z���0S�S殾ӱl�����;>�*���/���9�#1[�����v�-�&?��_>�,��)g��ҾA��>��ia0��i˽qx���؄>>�>���;+�<#��=~������u��=��>�n�����߆���=_h5<$��>P6��응=��[�J�8?�ts?�b�>,���}=؃o=�i>C��>a�7=���| >���>�*?�>�Q�>��$>�L�N�v;�*T>$Iͽc���# ��>�%�=?%H�(5���=7��= %>�.=���,a>-����CB?��?C�?%�?(�־�^5�L��8�r=�4�>�S�=Е�>�>�?|�=b�P>�L�>��'��*;�6�K�?�M!>�zq�R�\����>��= �>���>�?�>�(�Z�����<H���2i=�a7?c<?��ɽSNt>���꿶0˿�4�������<������ګ:��2@="�uڣ=�쩽��<UA[>�D�>@�<Zή:1�>n$�>��q>���=2k=��<�K�<y�<��<!S�<�<9ǽ;p���l�P �C���G7��\?�Fs������yB?˭�>��<Jp������o��-�r����>�t?��?G�>��\�F���,� ��@0������m�>w,n?���>����
�=}��:!��� �>�>,��=���*;�����+=���>�o�>��T>�m�@<7�S����0�>Cq=-b׽IƤ?��L?�W�F˾h�#�_��`�[�2�>�9��=�½����D��� �
~��V*���d�1�ӽ4�?:eu?������=T�ھ(����X�����+׽���=�?�0�>Ed5�B������z_>Qԡ�鄍����>U�`>rq�>
��>��>B�L?7��>��>�cP�P��>ت�s(�>�?���>��=,a�>��?���
H���.=\�b�hi����<N���D;=qm
>Ӛd>�y-��m��x�=���X&�;��=�� =R
�S�t=�n)>�K�=�aE>��?��?ٔ��>�߁=)<N��ȶ>�([>�L=�5	�kož�k'�n��>��>��>�D�>�>I0���5�*��W�>k �>\<?x�E>"�=�Q�Pj��9��6%��H*��$��vW���[�0��#�(�S�?Q��=�u���q>�cz?>]C?�!?v����/��.s��I*�I��NZ�����>�>��=��߾3���h�u_�T=1�a�-?E�1*=��=�S>��9>J�=�>M�&=G'Ƚ�j��:7;���S.�>��>e�?VT>�1�=���?��J�I?<Q��&����Kо�� �i>�v<>�g ���?���pE}������<����>���?�a�?�d?�xE��H�)�\>H]U>�>�"<j?�)���5����3>s�=�_y�Q��:�;�.\>�8{>�ʽ�vʾZk�J*M�'����uC��h�q���{��q�E�T��L�����=*_�<68;N᾽j�S�J��>���%������k �"q*?.3�>���=?͗=���q��������>�{�������%��KC>A��΅̾񐫾����־��&��{���1>FG���e����u�{�X�ɽ����vh�>��۽~�=��ƾk�S�;��[>t䌾R��Q����D>;�?�-?L�Ⱦ�$���"*:G����>��?��=hYɽu��7�>bw�>�L?*$�=�鍿�{o�m�>��?Ҧ�?[nk?�:=�v�������g>�?kX?x�V?6ӽY�/˰�8��=T�#?�B?�ؾ����YS��U?���>O��>�u>�n1>V�j�9Ơ�>N<�L�"j	>��>`�x�R� ����c�>I��>��?=�ˆ�D9�>��>�
=�%׾Υ^�i�=��3� v�����G��>�o#�U�c�S�>�I
��6�JA~�*~��A޽�?�+�?^?"Za?BG;�sC
��+�y�-> �?�9�>�}2=�.A�tQ�>o��>d|�9b�Zþ�W?���?���?زN?D�y���Կ�N��o���������=��=��;>�Nཝ~�=�GJ=�Ҕ�h_H�|�>�ٚ>�p>��w>��V>�e>>4�0>{+����#�R���㑿>�A�E\���o}f�	�]]v�Q������!�s줽aز�e_��%QG�z��'5�p>����>�Qi?4�>�ܼ��Z��/>������\�7=7�>����/��2,�c���=c�>IS^>`c��xX�[s���}��,?<���!<5�>����4U=�.>� <f�=)M��+=�̼���='�>I1�=�j+>� >�h>w�ֽ4y���Î��W.�n}���HH>�7?�+�<>���i� ��u4�0�[>�X+?�S�>yT��vy��kV���?�_!�u���ͽBY�>9֬>/�>�d>�8>@��;����%�b��>�:?���>��M��������>+�>K�����=>�W�> 1&?��q?7�b?ջǼ�I[>v��>M]�>oI7>7/>7�=��z=�?XT�>�)�>E��>)�=#�+8�=���X���r��*���Z��X�����<���X� >&��=~���>�=>B{��oM��>=�A�>&]?�s�>��?!��H��0u��;�'�:���Z�>&�>5G7>_��>`�?*�>ܱ��b�N�xT��<�>1��<�7��`�_�ac����3?@*H>nFw?��5?�t�=Ծ����YJ����>�*?l��>�B�>���=�K7>���yԿ� ���A���8���=@�i<DnU��᤽���<�
�����}<�PB>�H�>�8Z>1Ff>� m>Xx>�l�>�S1>�^%��i:>b/?�xڤ���=f�!<R��n=����,��j�=��0���۽(�ҽ(���qü�ג<���>�f?���=$�P�ܻ>���^�#��>��B?��/?�p�>cuR�gWM���|�`fX���n:��v?9t`?@>,�����A>Y�>�=�S�>����;�>Aξ�ɽ�yE��|�=s��>�,�>� >�i��KGN�.�S���9�]yU>��=&8=ႝ?�1?���X!���W۾qm��!TN�ц�>F�>栔>wp8��XA�s�����=l���!���)�=ݖ�>��?r�yc�>b澗G���=��骞����@��=�5�>j��>	��=��>�/��J�콼�*��= ��=��>>�`���>y��>��l?�s*?�!?��>��?��&>�D=P��=�>m�=?�H�>N*���w��F+>��>[S��Ž��=5xl�M�ں�g&>��=W�'>؄�$*�����=�)J=A�><�z2�	`+��?0=�*0=A3�=fp�L��>��3?�S=��]>�T�b<��؛#<�:�=��=��.����8����"=s%�>Io?��>uv>k���Pӗ�K 1��6�=ܦ?U_?yD�>������>{��ϼ��>�V>_Q�ʚѾf1��þ��z>���>���=�o�==b>�с?Ħ+?\.?�U��*��ny����8�;��D��>�>(ń>.I�<�����n�.X�����r="mD��Ou=E>���=���=�d�=�6>�a����A�����Y�Z�ݽ��>��>��?&�>&�=��˾acݾ��$?���iE��*�8þ!e	�f�*��Q�>��=�A%?�S�5����p���B���>^��?��?��(?ގ��H��]�8>���a�M;��>����sk�=Ww5�܌�>��>�D��k8�#�k<�>mԀ=m��Y�9�󪬾�Ҿ����P >�w�,��e3�q�������2�������7�m ���߾\9��u�V���6�a�(��뎾>ᾨ���ӱ��0��?��?��-�|�&�Y�t�g#�ޢ��_>�D���E���t8��tk����Ӿ��ﾄM���d��I�4��U�=Ds��F���䋿M����3=p�]>�H?7����˾�КP��j�=��>!����Y���������0?�F/?Tp��t��E��=�Х>��>�b��;>���BX ��S�>� G?�":?��/>bז�����$_�<���?`��?T�(?p����4�P
�"+�>�VK?a��>
�?H�,�!CA��?����?���?~]+?4�ݾ�Jq����?�!+>\@��5=.�>�mb>�&W�佽�vt=^ꄾ���=���>�4=ⷀ�,�v��v����>�">ކu��S����>T���3Q��4�2�F���C�!�J>S?=Wվ,3E>>}�>��Z>��:������(v��)�r+D?v�?��?
r�>�1ѾÌ�-z:=1��>�t=��K����=��*�>?�?��_�#��0��c�>���?���?��f?����9�&M��颓��g���R�=�=�.>MĎ���.��]=�G�=����<>�Ν>�'b>��&>	�>oP>A2>I���LW��؝�����c[F�m����޾o)����`��B��"@���3�����R�bhY<RB-�v�+�=`l�V�ξ��n>��&?S�?�?w�>���>֘��-���������t.E�AP	�'���#���=B��<���{�A
�'���F?�20�L[�<Ȍ>�^j�Yӥ>��>�M�=��P>�o[>��=$��>3��>J@|<�'S=�ؠ>L&>9'>i��=�@���ܢ��^Z�1�\��>�+?qky�ͬK�9s�P���=�N�T4�>�S?i�\>s�������j���?$?=���jt$� f�����> ��>L�>N�=>��C˾pCҽ�S>���>�-�>�������&Z��0>I� ?6e� z,��=�@?S�o?�S?Պ�=eu}>�uB>��> �=mӫ=b9��<<�0�>�,2?)^_?��>i��=�90��!#=��=)�	��r�<џJ;�yͽ��	�`ڔ<(����=n�I>�}�=��>����w�]*e���=>���>G?�\%?)�K?�w���y�@�Z��
�=❨>�:G����>%?T�?f3?F-l?I��>ƶ����()�|��>���=��m�KYk��~=�I>��h=f��?��Y?�싽��X�h(��6UJ=���<�@�=�U?��>��>�V>z��T_㿾����q���!I�|�F<���:u
�����X��U�u<�2H�>7�>`g�>�&
>Ջ�=c>��>y�P>~66=m��I-U=}f<ʞc��$�=~*�=^�<ؐ��=&�ҽ���k�Ap=e�^<������<���>��?�蚾@~#�*�.�A�#���	;%o?t�z>�r(?3b?}���;ﾽY+��E��ꏾ�G�>
ma?�,�>+P��y)��~��==^��>"?9�">��H�v�`�n��h����X�>��4?&�>k�	�1�jJj����� Q�>��N�+k]��;�? i`?�ྈ�7��G=��0m�!w��h���y�pl�����R
�^� ��pȾь�q�����i����>��?�Mʾ�u�=[���@��X}���9��k>��(�Ҕ�> �ؽ�?�}Ѿ?�2�0��F׾�=\\�>uRl>Ϋ�>W�>���>F�c?�?N��>û=��&?J��=���>76�>hHa?�v>?(��>�G��t�a��=J��>B̛�>1S��S >_7=)Q��y>�
>3�=J=�T�;8���]?�<0 ��t��Xsܽwyq=�O�=i�=}��=�a?ˠ%?��O����;��<���a�<�J�=�>hB �S�b�%�>���>�*,?��>�M�=��mZ���b��=a�>x�8?��?��K=k1�=$?������`��u@>�.���/�G����Ӿd�3�=�D>��^>tь=}}�<��? >�?�4?�<��O8����T�o�
?+7־5�?��>?��=ܣ�>f����)�&b}��p�8�:���;�<�`=t�>"Ν=[���m�>+,�ۀ��D�>��=S�a>A�>�#	? �(?�S�=B�L=���}-���C?fz���)���\�������k<�0>���<�֚�\�G?�ƹ�゙�������Dh�>X��?*��?�&Y?�9�(�Ͻ�$�=��?��H>��>��={����rv�n�?;ck|<�G�P�����?���>��>��q���ξ�{	�\TT�Ƿ��gM�����*�@ld������M_�2��k��n����mK�Ԓ������n陽ȟ�1+^��ɾ鲾Y�?�+�?��2�6����f��m��>ߕ���r�e&��
�3�؈¾��m=��ݽt�ƾPNܾ�����ԃE�Q��%�>vq��运�u���v���k&�Ƒ�>|@?4T��W��_�E
�>�I>���<��>����ދ�yJI�ՙE?'�6?�����-�n>�X�=�&	?���>�	�=�㴾��R�?C�I?��>�rپ����˘���=e��?.0�?S�C?�#��6x=�-{���#>.�M?�,?�="���������l�^�>�ha?8�>Y��qp�;���G?���?�qL���>
R�>�� >�"���ގ��	>��%�<�3�>��;;�@��3.�<���=�Z�= �=ͭP�2�`�8��>������f��y8���n��%��h�[>��"?�̰�V��>H�?�H���e��惿�R���b
�o7?��?��?	�4?Ռ �G� ��(�=�?�B�>*'�>ҽ>��<_h7?�T�>D�u��~o�
�:�M�?�8�?��@\Ay?��m�@<��m���̾D����P=��=ה->5&�]�">���LZ�=�3���@=Qv�>�~�>�N|>��)>�>4>��K�d}�����Fz8����'���������%�[����f���o޾�=���<�'���k\�G���ټu}ھ���>�+?�#?���>V{+>=dh>O~����۾�\�T!�m_�3���u����<f:低�ѾVF���+���0�=<?��=��>(��>�����}=�ӌ>�E����>���>��{=٫�>��>j��=A��=���=F>�yp>m�=����l>��Z�?���n�~E�;�ND?6a_��Z��8+0�;�oR��|�}>�?�I>Ԝ%��]��9Tv��B�>2U���o����^��B�>�˿>,S�==�'���s�������=m��>��=��Ƨ������ǽ=ī*?GeA�qw���>D�=?y|?Pw?��A�2���*6�>W���>�׭�����u�@�2?b�?,��?T��<X�<X:���\l>D솽����=?̖=Ea�B���T<�=�<E���l�=�C�=`�>|�=����k�_=�Ï>�Fd?��.?��?��,���s��\g� ���L??����?�/)?��d?��`?�?��S=(u���쾎�:�+��>�H3>��]�;��<]��.�>�,I>�~D?�9q?:���4�뷒<|o�����>�>XW?� ?��?g-�����otͿ��@�d�����#>+��=��8\̽۸�=U�e�y.��ݴ���l>�>��F>���=���=�9>
�>1d�=�:�=�>JQ��`�(=5Eg=6pJ�H�����=4�;� <�<uQm>�~R���ݽ͊��ݮѽ$�W{����?���>�,���x����/����<�t?/���:+?EXk?{D�=,��s�1���?�{d]��>%O?�߽>�}�EYy�\��`v�=@��>��>[��=����L˽|jo����v��>X��>Qq�>�?=�ZR���u���k�?�p�ϝ��u��?W�`?��J8O��:�V�<���h���ft�=��E�u�����.徘徻����Ⱦ$�:��>�٩?�d�Խj��R������NM�u�>�����h�>}!>����`־�W��O#�.���X��>b�	?M�V=V��>�t ?��?!�N?�;�>2T�>��>��^?~�={��>Z��>T3?!%?�<?_#3>�8L>�|�<c~��ń�r���#<l4�jL|=�$>��k>��=�K<:A$=03�<��l��_�y����3=l�<p�=�->2�/>t2�>�*?��<HV<����{_���<�
>��K>�3S=(bo���gG�<Zc�>�k5?�Y?$z�=��澱����Q.���>�?b�>?4�?���=���=^���f��9��$��>�wf�F�W�A;�3�	��꼾}>D	?>���o��-ԝ?�z�?�&	?��>>35����Q�"�q1?1�,��Y�>e�>粂>(Z>�ƾ;e�aNs�~�L���ν�1'��{��9�=h��>���=/ټ��>�m�����>�mH<�;�=?�>��?���>�i>R{�=�־W|��D?P��#�ǾL�����dM< ݣ>��4><���Xq?�Xo��؉�3p��h$��A?��?���?��?�N���g.�R�$>L��>6.�=h��V���۽�ZK��u>Ǡ���� ,��mZ���>�]�>�t4=�Mʾ:�O�=ψ����+�J��o�5U��ؾp�4��j�^_��u\�b����:C�,��<���j;���0�2F���'澧B�����?�T�?U�<ٳ��~�T�K2@��U���>�z�M���<p�����Lé��:�����C\��q��v����o>V��.����o���b��%B�1$[>0�?�{ᾡ�Ͼ
r���<a�;>�/�8&�[2��6鑿�.�M�A?�F?���-$��ٽ��F=�)?ͺ�>���:ֽ��h��bx�>?H?�?��3}��h�̽*�?���?��D?M٨�	%�e��Y�=�G?�?x��yþ�$��F�*��h?��q?!?0?(��&j��ܥm��m)=>�?Y`��u>>~�?>%[%>[
�jv��R�Cg1=�[�"�7=�w�=�o#�0�i�)�齇��;}�7>*�&>�}��DZ����?Ǵ:���u��F�cϾ�6�=�<�;1<;�l���6��4F���>�c'�Y'���͓��;ѽM�?��?ӦH?��?6	�ȷ��Y0G>�^~>֩�>&">m%s=���=�ך>[3?�����)s�>��~)?
<�?hQ�?�c�?0���dI޿�k����ɾH �����=��=�><N����=�ά=��;�f��q�=w�>���>ǣ]>�m)>��>�V�=-D���P"���Ŀ����w�L�C��YT
����S���#o��9:��$Ѿa꾴�e�Я<�)4u��G�="��1���V�'�>��<?�S*?�Qm>X��>x5>����/*��h���g�x?y�g� �l�!����x��=Q�;Jĉ�-���>�R�����>�<>U�=`r&?��o���	<`�>nþ�?��0>W�f;yщ>�ay>�J�=�AV=6VX>�=X��=���=�񁿿�{��#i��Ҿ	K>�S?(E�Nљ��
L�Ͼ|�'�d�>�S?�:P>� �5Ǘ��x��h?��Fʪ�����wE��j�>���>Z�q>3ze> f%��>���߽���<h�>�M>Y�"�b����M��8�=�w%?�39�e�X�g��>�$?��?��?���0�>�z>k��>�ɠ>f���T���J���?(j?�ɏ?=�'>z�i=�F���>q@��%�f	�=�F>v��=L�Խ��>4����r>lW�=5��=b�+>	<ɒP�����E>�{�>�\O?�|�>��>C@�;��J���_���*�f�>*7F��Y�>�(�>�f\>��>-?┠=z{���`�ݦ��#�>��9>�_n���|��8v>��.>(>�:?��?f]�<�ҽCg�=�̌��>���>n*?�K�>��'>������u�ӿz�&�#��Z��#�,�=qEϽ:V��r�������O�<`|>kr�>�9>�gF>w#�=u��=��	?���>8$>��]<0��>�ؼ�zp=���=8h��';�*V�=�=4��=Tj��(����jk�,[���ŽӁ%����>Cp-?�G ��T���3���
���w��X�>�ي>��?���>�N;>���1�I�U�@�y�����>�j9?���>��1{�=:�p���:��>hܧ>#Un>G��=��F���{�e�,�ŋ�>�?��>�M��?b�zYh�n����޺>̽��
�U��?�C�?sw3�SO>q�7��t��~9��翾3֊>�o�����!/�icؾ�����N	�m@����B��>���?{�.���=⬶�C֨��B���^D��;�>��#�D�Ἤ�w>��Ƚ��p��޾ז���_��Ъ%<��?=#&>�:�>Ȱ�>-/=m�l?d`�>W�?<1V>nn�>���;#��>��>6d'?�:a?u>�>��Y���}��;x��>����k-��h=�<�=�x�=��=t6f>�ٻ<��g>��ѻ���<�ui=$�-���	�M&V;S϶=@��=%�T>Q�?K�&?����#׽20=h�D���==�B> >�>=m�F�|tv=��A>���>Q/?*��>�|?=�����þ0�龍��=��>N�.?���>9d˼F��=YcپA����=�1^>�3�������߾���3�[���>���>)Y�=K��=cT�?��S?x�?{~>:�1뵿�k���m2?��c�>-?�h>Q�>s�=;�f��8�J�[�3�9���n��Z�ࡢ<��e�>�:<[4�=Qx;>��"�0����%B>��7>�=!=��>�3�>���>��>��>H�X�^])�|�F?�˾�CG��`Zx=�4Ľ]Uo�i��>R���J�>z.k?+���S5��3����"���?���?GZ�?#H?���_dJ�ã>p�?�~>H��+�<dP=��_�����/�>�ѷ����o6=)v�<dr=�2=�.��eo���轍���_F;�qW�����\��g�a9��X0�7s��ǹ����� �Q�;�F5��躽^��cH����ؾU	����?���?���������7���<���7�S�����#v�L�������Xӽ�9���o����������4�}6���>��=��d����q��r���d�>�F3?�1ɾ�Ǿ�@K����>,��>D%>�e������b��[r����[?�
I?��3�~�������>��S?�_h>v�y��6�@[�J:>�J?�T?��*�����ǅ���Lb��@�?�
�?�S?H�����p�+�徻=�y>�Y?�)??��1���/�-�0?%�\?��?GRﾫH����/�Z�=��?�X~���w>O�>��<U~����޾�d%��܅�H{=Ȁ>�H-=�.��b؅��L8���=�'>���=��B�0�����>T���3Q��4�2�F���C�!�J>S?=Wվ,3E>>}�>��Z>��:������(v��)�r+D?v�?��?
r�>�1ѾÌ�-z:=1��>�t=��K����=��*�>?�?��_�#��0��c�>���?���?��f?����9�&M��颓��g���R�=�=�.>MĎ���.��]=�G�=����<>�Ν>�'b>��&>	�>oP>A2>I���LW��؝�����c[F�m����޾o)����`��B��"@���3�����R�bhY<RB-�v�+�=`l�V�ξ��n>��&?S�?�?w�>���>֘��-���������t.E�AP	�'���#���=B��<���{�A
�'���F?�20�L[�<Ȍ>�^j�Yӥ>��>�M�=��P>�o[>��=$��>3��>J@|<�'S=�ؠ>L&>9'>i��=�@���ܢ��^Z�1�\��>�+?qky�ͬK�9s�P���=�N�T4�>�S?i�\>s�������j���?$?=���jt$� f�����> ��>L�>N�=>��C˾pCҽ�S>���>�-�>�������&Z��0>I� ?6e� z,��=�@?S�o?�S?Պ�=eu}>�uB>��> �=mӫ=b9��<<�0�>�,2?)^_?��>i��=�90��!#=��=)�	��r�<џJ;�yͽ��	�`ڔ<(����=n�I>�}�=��>����w�]*e���=>���>G?�\%?)�K?�w���y�@�Z��
�=❨>�:G����>%?T�?f3?F-l?I��>ƶ����()�|��>���=��m�KYk��~=�I>��h=f��?��Y?�싽��X�h(��6UJ=���<�@�=�U?��>��>�V>z��T_㿾����q���!I�|�F<���:u
�����X��U�u<�2H�>7�>`g�>�&
>Ջ�=c>��>y�P>~66=m��I-U=}f<ʞc��$�=~*�=^�<ؐ��=&�ҽ���k�Ap=e�^<������<���>��?�蚾@~#�*�.�A�#���	;%o?t�z>�r(?3b?}���;ﾽY+��E��ꏾ�G�>
ma?�,�>+P��y)��~��==^��>"?9�">��H�v�`�n��h����X�>��4?&�>k�	�1�jJj����� Q�>��N�+k]��;�? i`?�ྈ�7��G=��0m�!w��h���y�pl�����R
�^� ��pȾь�q�����i����>��?�Mʾ�u�=[���@��X}���9��k>��(�Ҕ�> �ؽ�?�}Ѿ?�2�0��F׾�=\\�>uRl>Ϋ�>W�>���>F�c?�?N��>û=��&?J��=���>76�>hHa?�v>?(��>�G��t�a��=J��>B̛�>1S��S >_7=)Q��y>�
>3�=J=�T�;8���]?�<0 ��t��Xsܽwyq=�O�=i�=}��=�a?ˠ%?��O����;��<���a�<�J�=�>hB �S�b�%�>���>�*,?��>�M�=��mZ���b��=a�>x�8?��?��K=k1�=$?������`��u@>�.���/�G����Ӿd�3�=�D>��^>tь=}}�<��? >�?�4?�<��O8����T�o�
?+7־5�?��>?��=ܣ�>f����)�&b}��p�8�:���;�<�`=t�>"Ν=[���m�>+,�ۀ��D�>��=S�a>A�>�#	? �(?�S�=B�L=���}-���C?fz���)���\�������k<�0>���<�֚�\�G?�ƹ�゙�������Dh�>X��?*��?�&Y?�9�(�Ͻ�$�=��?��H>��>��={����rv�n�?;ck|<�G�P�����?���>��>��q���ξ�{	�\TT�Ƿ��gM�����*�@ld������M_�2��k��n����mK�Ԓ������n陽ȟ�1+^��ɾ鲾Y�?�+�?��2�6����f��m��>ߕ���r�e&��
�3�؈¾��m=��ݽt�ƾPNܾ�����ԃE�Q��%�>vq��运�u���v���k&�Ƒ�>|@?4T��W��_�E
�>�I>���<��>����ދ�yJI�ՙE?'�6?�����-�n>�X�=�&	?���>�	�=�㴾��R�?C�I?��>�rپ����˘���=e��?.0�?S�C?�#��6x=�-{���#>.�M?�,?�="���������l�^�>�ha?8�>Y��qp�;���G?���?�qL���>
R�>�� >�"���ގ��	>��%�<�3�>��;;�@��3.�<���=�Z�= �=ͭP�2�`�8��>������f��y8���n��%��h�[>��"?�̰�V��>H�?�H���e��惿�R���b
�o7?��?��?	�4?Ռ �G� ��(�=�?�B�>*'�>ҽ>��<_h7?�T�>D�u��~o�
�:�M�?�8�?��@\Ay?��m�@<��m���̾D����P=��=ה->5&�]�">���LZ�=�3���@=Qv�>�~�>�N|>��)>�>4>��K�d}�����Fz8����'���������%�[����f���o޾�=���<�'���k\�G���ټu}ھ���>�+?�#?���>V{+>=dh>O~����۾�\�T!�m_�3���u����<f:低�ѾVF���+���0�=<?��=��>(��>�����}=�ӌ>�E����>���>��{=٫�>��>j��=A��=���=F>�yp>m�=����l>��Z�?���n�~E�;�ND?6a_��Z��8+0�;�oR��|�}>�?�I>Ԝ%��]��9Tv��B�>2U���o����^��B�>�˿>,S�==�'���s�������=m��>��=��Ƨ������ǽ=ī*?GeA�qw���>D�=?y|?Pw?��A�2���*6�>W���>�׭�����u�@�2?b�?,��?T��<X�<X:���\l>D솽����=?̖=Ea�B���T<�=�<E���l�=�C�=`�>|�=����k�_=�Ï>�Fd?��.?��?��,���s��\g� ���L??����?�/)?��d?��`?�?��S=(u���쾎�:�+��>�H3>��]�;��<]��.�>�,I>�~D?�9q?:���4�뷒<|o�����>�>XW?� ?��?g-�����otͿ��@�d�����#>+��=��8\̽۸�=U�e�y.��ݴ���l>�>��F>���=���=�9>
�>1d�=�:�=�>JQ��`�(=5Eg=6pJ�H�����=4�;� <�<uQm>�~R���ݽ͊��ݮѽ$�W{����?���>�,���x����/����<�t?/���:+?EXk?{D�=,��s�1���?�{d]��>%O?�߽>�}�EYy�\��`v�=@��>��>[��=����L˽|jo����v��>X��>Qq�>�?=�ZR���u���k�?�p�ϝ��u��?W�`?��J8O��:�V�<���h���ft�=��E�u�����.徘徻����Ⱦ$�:��>�٩?�d�Խj��R������NM�u�>�����h�>}!>����`־�W��O#�.���X��>b�	?M�V=V��>�t ?��?!�N?�;�>2T�>��>��^?~�={��>Z��>T3?!%?�<?_#3>�8L>�|�<c~��ń�r���#<l4�jL|=�$>��k>��=�K<:A$=03�<��l��_�y����3=l�<p�=�->2�/>t2�>�*?��<HV<����{_���<�
>��K>�3S=(bo���gG�<Zc�>�k5?�Y?$z�=��澱����Q.���>�?b�>?4�?���=���=^���f��9��$��>�wf�F�W�A;�3�	��꼾}>D	?>���o��-ԝ?�z�?�&	?��>>35����Q�"�q1?1�,��Y�>e�>粂>(Z>�ƾ;e�aNs�~�L���ν�1'��{��9�=h��>���=/ټ��>�m�����>�mH<�;�=?�>��?���>�i>R{�=�־W|��D?P��#�ǾL�����dM< ݣ>��4><���Xq?�Xo��؉�3p��h$��A?��?���?��?�N���g.�R�$>L��>6.�=h��V���۽�ZK��u>Ǡ���� ,��mZ���>�]�>�t4=�Mʾ:�O�=ψ����+�J��o�5U��ؾp�4��j�^_��u\�b����:C�,��<���j;���0�2F���'澧B�����?�T�?U�<ٳ��~�T�K2@��U���>�z�M���<p�����Lé��:�����C\��q��v����o>V��.����o���b��%B�1$[>0�?�{ᾡ�Ͼ
r���<a�;>�/�8&�[2��6鑿�.�M�A?�F?���-$��ٽ��F=�)?ͺ�>���:ֽ��h��bx�>?H?�?��3}��h�̽*�?���?��D?M٨�	%�e��Y�=�G?�?x��yþ�$��F�*��h?��q?!?0?(��&j��ܥm��m)=>�?Y`��u>>~�?>%[%>[
�jv��R�Cg1=�[�"�7=�w�=�o#�0�i�)�齇��;}�7>*�&>�}��DZ���5?����`���Z������^�>��]�� >?�	�����]�?�{n>���K�{�è��ur��,q?6��?�Nf?�)? )�1=�����>Y/�>O�>ǚ=[>Qu�����Jp:>K�Ⱦ�?����J�i43?�J�?���?8��?3��kgο%3���aҾkg7���=�޼��>���6�g��h��K���*=W>_=?�l>y���>*m>�l�=��> ��� �'�W¿�Ԑ���.�:N�^�jʆ��y6��(���~¾�����T�>���	��x�@� �Ne��s���d>��?0>?i��>��f>
�T>�-�8���徾 ����(�t�5�]��Wy����v=#�j��{�g��SV�`p�!?�W����޽e/?�6��*W��4�>�o�C[�>4W>�<��>9>�x=�ڬ=��=��>Ȭ>�3;>�_o��vg��l��u4�!��= �I?�잾��˾����KB��X�:���>��.?����8nH������Ք��4�>ᴮ=bz���M>�܆� /=-EV>��=Y�D�^߂=���$�Ë=9�>.��=M�-o���J��==֭�>�3پ�M�=��q>��(?�Hv?j�3?��=g�>��\>U��>�j�=��C>E%>> �}>N?h�<?�w4?��>���=>>]�-�
=r�%=��;���>�j��Hi��L�a�<^�H�Yd0=�i=�U;� X=��H=�OP����:��<��>j?�q�>��>���
R�k�w�Tk��T��>�_l>���>��?}�L?M�*?�J�>/ҏ�q����x��ʾ���>�1:>.�X�桎�	x���>(�<�
?ڕ1?�*>"�����B��>->"?{�?� ?���>� &�x��I�Yw鿧��1ξ'�0>.k�y���ؾ�ԧ���ž��þqwL�ʶ���=�KI>)�=�T��.�=c��>`J�>o`L>�a�>Z%p�v�2<��=�33�ݒ�<ؙ2>V�r>7�û�L���I�=�F��2%>m 9���?=Ɖ��1����?� �>G~�<����8#վ�C� �"��\B>�$=+�
?�%?��=�s��e�R�`�"�/	?pG?Q��>��+��>Y�N�jf���~����n>���>�ui>�>�(�=-*�>1�8?�=j?�7?/~�H[��:񒿥�0����>�
M=�5 =m=�?�j�?D����'��j?�	&�~�M��=����þJ!�u�A��[�kP�w���NҼ�>=�>���?/J��t��=Pʤ�	O���������zD�>g�=S+�>F=�u������.��{��bl�$�>Կ>am�D��>��?�_!?�3�?�?�6K?���&tB?�E?�i���?M9 ?f�*?��?=��>�`=:���옽z7"��Ү��Y&>�6�=�$$���=��4>���<i�L>���=��Sս?�����8������m[=�g=�B�=��>qyN?��<�����e�����N��
&t>ͳ�>��:=��9�j���>V�8?�@<?0x�>�.B�gn���!��B�E�=}�?s8?:�?6N?��%>�޾��j�=5��>���>^#ʾ&��L�� �ͽf'�>d�>���>�C5>��}?�<U?��K?2���;��b�1�/���>U����d>���>`ӏ=mP�;�6���N�/.U��+�~a�=;�?�V��=���]��>hӖ>��_�N޻>�؊>�/޾!w��{
�I�	���a>_i�>.�>sD�<��G�Fn�T����jF?�l��������]�9�р>�g>J\��F��>/:u>đO�(x���Mt�Q��>^��?��?g��?f 羗镾���>�cs>4��=ɗ�m����u>W���u���^>�aܾ�B����a=���=;�<2�,�gԾ%G"�{�y� ��?t9��׺�_�-��^���(&������9�<L f��iL��i	�1���o�x�$q�)p�<>�����f�쿨�ہ����?A��? k����dD�`�4���F��	?�G�r�¾� ����\=4l"� �b�;����������������>aڌ<0���Q[G�[�P�` �����=��K?����񌾞�ͽ'�>��>C�H=�, ������e���6����i?�|H?�2��)߾�ҾS!?�s�?�GU>	5Q>j�޾�e�= M1?. ?��.?�nͼI䗿A,c��l�>���?��?1v8?��|kF���>� ��L�=?�R?0?��W-žz�>|V?��R?ˁ?���������L�>v>�Dk?H�T��n�=�z�>-^>{��=�}��d0����S��(�=j���T�&����3�o��>�A?I�U=�u����[��>|¨��`��E����������9��q{�>���8[�̃�>��<׈E���ً��&��U`?��?A2Y?c�#?R����#�"#>HJ�>k>b߬>E�������=�l=�U6�Td����@�	�?���?�'�?��?
՝����d`��X̪�[8���.�<�7�=�O�>�� �酪=~)&�o���<�wH>F��>q�T>�/�>�>i>�7t>;�g>0���;(�Zΰ�4���5���޾5@���V �Lu����@=��u��;@��{n���:K�׽EBp�o�����s�2>��?U��>o��>z�>�ӊ>Cо�r��������+.��|��窾�
�r!_�M�ž�Q�-P���q���9�$?l��>�慾��?��۽��=߇?��u�8^�>rDT>_6�<ĳz>	���[�=�N�=�H>� �=���>�-v=9@Z�g�_�Nu)���N���U>�"8?��[������_�KF�j���ߪ:?��Y?mt ?6�)�����pg��5�>~���+�=i��������==�?�~�oB�=�2�v��_!��Xu�>%J?��L>���C]پRe��6�>�m�>�׾OM�=8Iz>\�(?a�v?4�5?���=�'�>�^>۝�>K��=�cH>Z�N>�ȇ>n�?9?`�0?e��>��=�2`��=t�8=E�?��|W�fR����J.,�@6�<(Z/��LL=�Fl=O�;�Oj=�@=�üi�;��=���>��P?{m�>�g�>��G�JbI�� C�$���s>�<X9���>u��>p�?&P�>���>��=��$�\���&���غ>��$>��I��p��Һ�|e>�z�>�[I?F�0?���<��"=6#\=~��>~	?/ (?�ǿ>�b�=N�Q�Y}�e��c���8�ܮ!=�I>�Դ=&A��(G���Y�� \���ؼ��&>���>��>�]d>��>���>/�>�(�>|#�>�.�=.'=��=��μ�]�m9=�p���9=�k�<l��=������we�<ﺞ��V�����Ĕj=��?!H?I�$��F��KnѼ�����.��O>� �<���>�H ?��@>�w���x���\��g=���>K�m?;~?�h���o>;[�0r��lK>��>�H=�铽q���5�?��$U>���>�b?ֵ�>�K$�,�u�k?���2+����>�;�=�"<
�?#�?|�_�C�νW����˃�<տ����#2(����Sj����y�*��v�9{�ތw>	��>��?��n�r��=.�ľ�4��/$����{���>z��>I��>�(�=yM�����#�����Bؙ=�>�;�>Dɇ�����_�t?Gjq?_�|?�q?vr?ל&���>}9?�
�>z}#?mF?�	 ?��>�[>�CW�V�~�MΏ��ѽq��_G��W�=���=fc6> >.���	�;���=xó�ܷ?�@G�=i��=g����B:c>�]>�, ?�&-?���>16D��L�=2��L��>W�w�ű�>�)�3bG�֨��:�>=3?��t?�<�>�Q���=������(���>z�?o*=?m�?+�p�Ֆ�����
����I;ܩ�>[X>���T���/�;X!�I�>���>lO�;s�x>��?��7?��>-0{��k�ay��Y��6�>\Ҽ)��>f�?ܐ�>c����X0�����{�z��F��2!�~��>Pe>��w��%>d=�1�>0�L>�&����v{����'
?o�>S?�� >(н�㾽��Z�??s þ:7�I��	��9����j�D?͊�� c�>�A4�%{W�v�����f����>�?}b�?S��?��edǼR11>KH>�w��>-�'�<C<��=�>b�>�D�:�l��>���>���>l�=u�Ӿ6���������R+��˃���3�z>߾mM��#H��![=w�������&�=䮾�_A��o8�9�ϼ�K*���<�����j��桩?s��?->_��̽8�Y��U�FhȾá�>�&�tAK�C�Ӿ�₾��l�~x��G���T	��(W�wO�-�^�H�H>��{;�;���І��<���P�W�f�:Vp?X���,�/M���V=��m>�ف=&���������;��JJ1?J?s� W�(�R���>ܴr?��> �&>�����"���?z\?P)
?���:r���_�����;�v�?ݮ�?gT ?y㥻�]��%+�sU����?K�>�#?"���xx=̪?�u:?�\?�?�>S2J�񄡿�B �4��>�9�?Ѧ/���=b�?���>����T`ƾ�8��֝l�_�>9�F>ңۼv^��	���{����N�>4��>QnC���н[��>|¨��`��E����������9��q{�>���8[�̃�>��<׈E���ً��&��U`?��?A2Y?c�#?R����#�"#>HJ�>k>b߬>E�������=�l=�U6�Td����@�	�?���?�'�?��?
՝����d`��X̪�[8���.�<�7�=�O�>�� �酪=~)&�o���<�wH>F��>q�T>�/�>�>i>�7t>;�g>0���;(�Zΰ�4���5���޾5@���V �Lu����@=��u��;@��{n���:K�׽EBp�o�����s�2>��?U��>o��>z�>�ӊ>Cо�r��������+.��|��窾�
�r!_�M�ž�Q�-P���q���9�$?l��>�慾��?��۽��=߇?��u�8^�>rDT>_6�<ĳz>	���[�=�N�=�H>� �=���>�-v=9@Z�g�_�Nu)���N���U>�"8?��[������_�KF�j���ߪ:?��Y?mt ?6�)�����pg��5�>~���+�=i��������==�?�~�oB�=�2�v��_!��Xu�>%J?��L>���C]پRe��6�>�m�>�׾OM�=8Iz>\�(?a�v?4�5?���=�'�>�^>۝�>K��=�cH>Z�N>�ȇ>n�?9?`�0?e��>��=�2`��=t�8=E�?��|W�fR����J.,�@6�<(Z/��LL=�Fl=O�;�Oj=�@=�üi�;��=���>��P?{m�>�g�>��G�JbI�� C�$���s>�<X9���>u��>p�?&P�>���>��=��$�\���&���غ>��$>��I��p��Һ�|e>�z�>�[I?F�0?���<��"=6#\=~��>~	?/ (?�ǿ>�b�=N�Q�Y}�e��c���8�ܮ!=�I>�Դ=&A��(G���Y�� \���ؼ��&>���>��>�]d>��>���>/�>�(�>|#�>�.�=.'=��=��μ�]�m9=�p���9=�k�<l��=������we�<ﺞ��V�����Ĕj=��?!H?I�$��F��KnѼ�����.��O>� �<���>�H ?��@>�w���x���\��g=���>K�m?;~?�h���o>;[�0r��lK>��>�H=�铽q���5�?��$U>���>�b?ֵ�>�K$�,�u�k?���2+����>�;�=�"<
�?#�?|�_�C�νW����˃�<տ����#2(����Sj����y�*��v�9{�ތw>	��>��?��n�r��=.�ľ�4��/$����{���>z��>I��>�(�=yM�����#�����Bؙ=�>�;�>Dɇ�����_�t?Gjq?_�|?�q?vr?ל&���>}9?�
�>z}#?mF?�	 ?��>�[>�CW�V�~�MΏ��ѽq��_G��W�=���=fc6> >.���	�;���=xó�ܷ?�@G�=i��=g����B:c>�]>�, ?�&-?���>16D��L�=2��L��>W�w�ű�>�)�3bG�֨��:�>=3?��t?�<�>�Q���=������(���>z�?o*=?m�?+�p�Ֆ�����
����I;ܩ�>[X>���T���/�;X!�I�>���>lO�;s�x>��?��7?��>-0{��k�ay��Y��6�>\Ҽ)��>f�?ܐ�>c����X0�����{�z��F��2!�~��>Pe>��w��%>d=�1�>0�L>�&����v{����'
?o�>S?�� >(н�㾽��Z�??s þ:7�I��	��9����j�D?͊�� c�>�A4�%{W�v�����f����>�?}b�?S��?��edǼR11>KH>�w��>-�'�<C<��=�>b�>�D�:�l��>���>���>l�=u�Ӿ6���������R+��˃���3�z>߾mM��#H��![=w�������&�=䮾�_A��o8�9�ϼ�K*���<�����j��桩?s��?->_��̽8�Y��U�FhȾá�>�&�tAK�C�Ӿ�₾��l�~x��G���T	��(W�wO�-�^�H�H>��{;�;���І��<���P�W�f�:Vp?X���,�/M���V=��m>�ف=&���������;��JJ1?J?s� W�(�R���>ܴr?��> �&>�����"���?z\?P)
?���:r���_�����;�v�?ݮ�?gT ?y㥻�]��%+�sU����?K�>�#?"���xx=̪?�u:?�\?�?�>S2J�񄡿�B �4��>�9�?Ѧ/���=b�?���>����T`ƾ�8��֝l�_�>9�F>ңۼv^��	���{����N�>4��>QnC���н(��>X]��d�o�Y41� w5�����^���;r+?�y������ہ>
�R�`3�U�����/���%L?ac�?B�Y?�4?�=�b1��Q����֤>�Z*?
���G�>�9m��S>o�>�9�Y����-���1?���?��?\�p?�a��p'��6���s���|���\<>�ZO=W�B>	p�W�!>brм;T����=��l>���>w�>�>*>f>N$X>��s>�̂�A'��{��O��� ;,�����"��f�}��Z��9�,o���˓��E7�E���Ȅ�վ	�>���-�<�ۉ�q �>3[?��?EZ�>v��>!��>�41��߾	�8���;	:���ؾ�?��R���=�������G����º;:��R�?��<(��f<?,���e��>C�Z>`��=���>���=�->�#>q��=o��>_o>E�>t�>̼>�48�%U��r��L7���M���>x�&?�P��7���R�Rw#�FӘ�4N?��O?��>_��g7��C62�LȨ>������>U`J<l'̾�/9>+�?�u�*�=aJb=�n'��`����>@�>�o�>����ڪ�a����V�=���>��־����dd�=1�~?�e?L+A>���>��<�S�>��1?����i������L=���=?�k?�f?��=��=����D��<�<���2c�2�
<ޙ�� ��@�Y��uF��gA>�cB>����5n��i���lm=��=I��=��>�;K?��'?��> ����d�cQL�w3��ӗ>���*@;0��>�cM? ?���>���֠��s�ﾽ������>��>�fK�����i�����=�O=D1\?���?b������|���I>���>��?��?<��>
�=����1��]��{�*�(�C�=������J�ޘ���)�x! ��O�=��=9v�>�?�>	�=>�))>�K�>P��>F�+>���Q����=�,=�.^<��b>�z�<4Eȼ7h=|6o=��6������6<K��Y=�I�x|f��(?ii ?��/=��{�P�ѽ��{�4��� �>wu?
:? ��>Uq�=��о�Y���B�d�����?M�l?�G�>��	���>��4=��z��
d><z>�r>��u��Ҿ��ٽ��Q>"�?e!?zԛ>�N��׎���P�8����>�c�<[V2�E�?�*�?D����:Y
��D[����-�c�Gd������NZ�W�N��s@Ҿ��p��cQ6>%[�>�)�?j��ͽ����k��%.�����`�<mU�<��=��>��ýI`���cھYv���F�\[[>��>�ԅ�6f?_O?��1?��=?�1�>g�??�{�-?%�O��>��-?et,?��?y��>���=�=�ti�
���s�����(�	> ��<07>�5$>���=�BA�ps��v�=�>>��=�w=ҽ�=�x�;��$����$�W<%q�=�>�,?���>%ã=�����k��Ӂ>����9�>~kF=�RG�U�����>�A?W�n?�
�>H�E����b��R�GL�>e?G�7?��?�׉>��
>b�L�湩�⌠�T`�>��L>�	���I�o���"��0
�>�|?�:>�;>�yf?��]?�pr?M�g���P�c�R�C$���!=��s>~�>�?�>�l�>��B�Mu���wu�F����j�` ���U��3
>�8>��f>!U"����=�#3>X|��=�[�9�x=
��=��?���>���>P�k��U�:!ܾ���r�,?���_�L��+�!��=fR|>�9c�N�?{־`i?��h>�T�������H����>5��?E[�?�~<?�%���Iȼ@
>r{>K�H>ak�= ĩ��f�>�,?�k>�A�>�W��5��ĺ�=�*?���>���=h��d��o��u�ȿ�DO���Y��D�!g���븾Ls-� (�lF��jQ�[پ�,��{E�%ќ=I9½HV��d��ˌ���`E�c�?ֈ�?�O���h��HW���F�H���`��>|��
QO����,I����X鰾E�
�wW8�"8����.����C>���j֕�P�z���;���M�]J�>0}0?�H;��I?��$�=���=��=�k��a���j���9��Ym?#mX?EF���4�4�=��= ֲ>���>:�p>��
��<?��>C(?��2?�'+��嘿nލ����<�+�?��?\N-?~Ă�.d/�۶��O�����> ��>�[>._��r��y�=
??�d%?��>'�h�_���u������>�H�?��=�t��>z�>���>詶����.&�=�����=���<*K��gæ�v����.���?=/�>�N<>�TR�`RU�(��>X]��d�o�Y41� w5�����^���;r+?�y������ہ>
�R�`3�U�����/���%L?ac�?B�Y?�4?�=�b1��Q����֤>�Z*?
���G�>�9m��S>o�>�9�Y����-���1?���?��?\�p?�a��p'��6���s���|���\<>�ZO=W�B>	p�W�!>brм;T����=��l>���>w�>�>*>f>N$X>��s>�̂�A'��{��O��� ;,�����"��f�}��Z��9�,o���˓��E7�E���Ȅ�վ	�>���-�<�ۉ�q �>3[?��?EZ�>v��>!��>�41��߾	�8���;	:���ؾ�?��R���=�������G����º;:��R�?��<(��f<?,���e��>C�Z>`��=���>���=�->�#>q��=o��>_o>E�>t�>̼>�48�%U��r��L7���M���>x�&?�P��7���R�Rw#�FӘ�4N?��O?��>_��g7��C62�LȨ>������>U`J<l'̾�/9>+�?�u�*�=aJb=�n'��`����>@�>�o�>����ڪ�a����V�=���>��־����dd�=1�~?�e?L+A>���>��<�S�>��1?����i������L=���=?�k?�f?��=��=����D��<�<���2c�2�
<ޙ�� ��@�Y��uF��gA>�cB>����5n��i���lm=��=I��=��>�;K?��'?��> ����d�cQL�w3��ӗ>���*@;0��>�cM? ?���>���֠��s�ﾽ������>��>�fK�����i�����=�O=D1\?���?b������|���I>���>��?��?<��>
�=����1��]��{�*�(�C�=������J�ޘ���)�x! ��O�=��=9v�>�?�>	�=>�))>�K�>P��>F�+>���Q����=�,=�.^<��b>�z�<4Eȼ7h=|6o=��6������6<K��Y=�I�x|f��(?ii ?��/=��{�P�ѽ��{�4��� �>wu?
:? ��>Uq�=��о�Y���B�d�����?M�l?�G�>��	���>��4=��z��
d><z>�r>��u��Ҿ��ٽ��Q>"�?e!?zԛ>�N��׎���P�8����>�c�<[V2�E�?�*�?D����:Y
��D[����-�c�Gd������NZ�W�N��s@Ҿ��p��cQ6>%[�>�)�?j��ͽ����k��%.�����`�<mU�<��=��>��ýI`���cھYv���F�\[[>��>�ԅ�6f?_O?��1?��=?�1�>g�??�{�-?%�O��>��-?et,?��?y��>���=�=�ti�
���s�����(�	> ��<07>�5$>���=�BA�ps��v�=�>>��=�w=ҽ�=�x�;��$����$�W<%q�=�>�,?���>%ã=�����k��Ӂ>����9�>~kF=�RG�U�����>�A?W�n?�
�>H�E����b��R�GL�>e?G�7?��?�׉>��
>b�L�湩�⌠�T`�>��L>�	���I�o���"��0
�>�|?�:>�;>�yf?��]?�pr?M�g���P�c�R�C$���!=��s>~�>�?�>�l�>��B�Mu���wu�F����j�` ���U��3
>�8>��f>!U"����=�#3>X|��=�[�9�x=
��=��?���>���>P�k��U�:!ܾ���r�,?���_�L��+�!��=fR|>�9c�N�?{־`i?��h>�T�������H����>5��?E[�?�~<?�%���Iȼ@
>r{>K�H>ak�= ĩ��f�>�,?�k>�A�>�W��5��ĺ�=�*?���>���=h��d��o��u�ȿ�DO���Y��D�!g���븾Ls-� (�lF��jQ�[پ�,��{E�%ќ=I9½HV��d��ˌ���`E�c�?ֈ�?�O���h��HW���F�H���`��>|��
QO����,I����X鰾E�
�wW8�"8����.����C>���j֕�P�z���;���M�]J�>0}0?�H;��I?��$�=���=��=�k��a���j���9��Ym?#mX?EF���4�4�=��= ֲ>���>:�p>��
��<?��>C(?��2?�'+��嘿nލ����<�+�?��?\N-?~Ă�.d/�۶��O�����> ��>�[>._��r��y�=
??�d%?��>'�h�_���u������>�H�?��=�t��>z�>���>詶����.&�=�����=���<*K��gæ�v����.���?=/�>�N<>�TR�`RU��C�>ռ��3�m�	��F=i�z5���l��ך�>pX4��x=>� ?i%�/�̾vꁿO^��0I��g�.?��?'�R?��F?��=5�^�ž�ʺ>̓?� {>q��=ST���>_�?����5�����!�>���?�2�?��N?�2���2�������Լ��Y�>@88>�b!>՛u�[]>�>�8��ǩս��o=O��>{�>���>l>�i�=_�=������.��|��Up��}�`�A���'#��������#��+9����(۾R�K�N'�zz�.Dq���G��j��6��>6]6?��?d��>M���!n>h�����iS�=}��`����O��{龵)�s��=D+[����a�����^�	?W@�^}>�i�>��<��=mCP>�߂��ў>w�>�|�=��=hl'>'��=�w����=�t�>�->��=����2����
#��Z3����<�4?�􄾻B۾��/��`��KؾХ@>m��>�G>�d5����w u����>c"�<��z�����T�_Nj>G�>��ۼH	
��-���L��!x�K��=S�K>-�d=����⪾� �>M>^�>�ž��g�4̫=%$�>y|?�$?�38>4��>ڐL>��>�r<>���>���=�P>h�>��>?�'?�N?��=ݓ{�5��=�&^��v�t��=~���;�Θ=g�ݽ_]9>*�=Z�:=*�E>Y%�=�s;Qo�=�,ڽM�>N?+?3X?�ʦ=�X;�y[������O>%��>AD>�ҍ>�w�>1y�>�I�>�g�=�����d۾绲�"�>�AA��_u��/Z���?�u>�Qq>a�b?7��>�lM<�ס=(��ܩ�>��!>I�>�(?���>�%�>|�;x/�	�7�@�C�*���.�@>�y�s9g��dǽoo[�/�X�n��z�<.��>-B?ҫ�>�Ś=;�ڻ��ۼ~S�>���>�~:��*Ѽ�ܹ=9��=���<odq>0�S�'w��-<(���|5�5��|���]�=�T��/dU=�:�ԟ?�E?��ֽ��轡�G��sԾ���g�>6�>��?���>q�)=�����T�deE���н�?0Tc?V��>��U�in�=�����{@�>� ?��v>Ӡ����1�V���{E���?��?��>Oף�&'H�2pQ���	��Fk>UҼ� >�B�?��W?�f���̺������W����'g=N�n��������J:��"����w�
�+¾&�D��M?:��?kz{�\sI>�y���k���8���?L�-�>S �>���>A�>�be=�>��|�1�mk�$�2����dW5>�J>Ӊ�>� ?Н�>�N?K�>l�	?߫�<U�>2P�>�>���>�0?0;?���>��=9[�<�a,>��=���,�q�����A���S��=��>�vn>�A���C= O�<���:� >2�t=s��=t��=K��<ɾ'=f4>Z�w=���>�o-?�>���>�%=�Ν�J|�BR>�N)>4�(��F����<Q��>L(�>OY?���>����@�2�(�x����6S=��S?��,?x�>�">2�>@����ɾ�n,> ��=����@پ3�btq��Iٽ^Z9>p̢>>>�I>Β?�po?�h-?�^|>��I�/﮿9Sa�c��>.-R>��ѽ.��>�>[����:�"J*�^D��\���@���׽�Z� �=7�=��=�g<0u�=�p>a��=i���W;; �X��q?r��>��?�7D>wg[=�>�����S9?��	�4sz�~=�<����/����I�=@<�;�?�.?�Y��e����w�D�{,�>ϛ�?��?�X�?���+5���Ǧ>��>	��> ��=H�ݾg��=1��Ar�<{�=��NF(�$b����=���=]�(��[��r�ܾ0�;�����\�{?��u��{5����A������&�sAо77����ľ�d�c�ؾ��@������T�K?���ھ��Ѿ(��?��?�v�<Mb�����
��SQ��@���I�or���f����qT����������LZ��L�������=zC<��������N���j��ؚU>n1�>�{�{��%�<�����x弆�J�[�/�l����ޤ��#����??o�9?�,����ƾ��C>8������>Ͽ�>��=t�?�Ec>�>d�H?(d?�Y!=�Q���A���K>�?h��?yr5?����n��#ݾ��߾j.?�1?��=?1���$��r�>��N?�PT?��?J`��}au�>=ƽ���>�m?��=�0 >��z>���>{
�bX�ʍ��#l�������=�D���X=�i�>�pdn==n�=*�g=z��=��u�͸S�b�?���5�>p(�|�پ �ýJB���{?�lؾXW>p�g>���=k�%��4���Z�%M�;�H[?�s�?��??��?\�L��6J�=�����>pۓ>�\=ŵ~�6��>��W>�R���ۏ�8R�)3?/��?H��?ʸ�?�v��hnۿݰ���ث�!�����=u#>=�>?Sʽ�l�=�9z<�)<��;M4
>g�>#^>�ev>��
>c;>��=FI��!��ɎͿB{��i�d��u8�(��
�1����3���a�(1��X���]���+H�, ��e;���؎������r�>��:?Ut4?��$?����|{=����@�
��=@q�Mu!��r����S�
��!ƽ��,��% �ʍ�0��:WܾB��>i���d���>�oG��N>���>v��=^��>�A>W�0>F�>�O�=���=��ν#�I>��=
v=� <=���O{��P_�(���x��=��]?"g��F�˾��0�\�޾W�O�6x�>E�?�>��>������\�n��>.o��j�>>��IȀ>�E�>�,==u���>��ѽ�n߽��L=��=�N`>m�Խ��Z�5V�8?>4 ?�.׾tp;M��=��?�Iw?f�?�)%>Q��>X��=��>�UN>@��>:�>[�*>�F�>Y�"?d)?T!?��=��d�JY�;r~<��P��.��T��"��$?����=H�ν=�j��<�	��h�=X,8>�0�<6�=z���4�>'L7?�&�>��>ph)��B���M��� �F
>"��<|��>��>���>���>�:�>,B> �`����྅��>�8>}�_� �x���޽]�|>�.O>gQ?ϓ0?IG4���1�T�[<A�>'t�>���>�J&?�̱>��#>��h����lӿ$�f�!���Y���;q�<���M����7Ξ-��������<��\>3�>/�p>EE>��>�93>�R�>fHG>�Մ=:�=Q9�;�m;]�E���M=G��AG<��P�E^���&Ƽ���������I�'�>��;�[4ټ�y ?���>b����E��߳�f5��w�ھ!d�>��?j��>��<?���<:���B�=��i�	K�A��>��*?��??����w����#���<�'>���>���>�\^=W�$�L���B����?X�?3�J>�%�<9�M��(.�7��p	>y��U5g>V-�?��g?zU��C岾�H�$R{� ����E>d����p��@t˾P��Q�I��u�������@8��]?bӧ?8>I<�]��CY��lk�[!��[���~8>)~}>�,?R�)>�Ͻ�a���E����T�;\{V����>���;rƹ>cY?>�?�a?�E?a��>9�
�j�>X>�]�>���>W��>M�+?���>1`s>���>�7ƽ4��`�Ͻ�r0�d�:�j߽�l�=]{=B�=._d<+g�=���=P��=xr;��)�ý�^��N>�7�=�>h<>�e?�m)?Å���p-=s-
<����{>2˼�&�;���U�־/��Ą�=��*?B�S?�V?�cO>2nپ�������>.,?��??3$?$ 
>=��=L��}�̾�'�=�#>)E�=R��-\����O����L>��>Y1�<a]'>�:�?b_�?��Q?�G>�& ������m�o��>?��>��]>u1�=I�q<��=�I�9u_���q��Jb�t�S�Q#��w���U=\��>U@>Ӌ��&�>�i�>+�t���D��!;���<쇭=�ѝ>G*?��=DG�<Ю0>�*����R?+:�����a�=�wȾ"M��(n>5�=|+�<8?[����;��dW��˼��Y�e?��?�?�g?k��Ѷ��/		?�;>�>i>�=�!��E:k>���i8½�uR�I�����þ���=�B�>��>�>`1����;C�	�ο�~�)>�e۾����t��,у�k��;�{��BF��+}���u�  �֘B=r䋽�񚽗 ̾o��� ޾4Q�?�h?�Uֻ��3�yB0��E��亾*�>-T��^�i������h�g����վ�־�h�m�T�"�3�����{=�篾����:��X��E���-�>��F?4�ھ���,�{�C6;>F��>N >�V|�0ΐ�g
���ш=V�G?�E? �I�9��BL���>v�:?�;?���=Nyd���<���>0�q?PI ?��>4t�bu���n>
�?⛟?c�?z�/��D��Ya�,u޽��?�t?�A ?`�ۻ�1>����>�kk?�$q?j �G$�u':�þZ�?��S?n⹼��>��>�6>�`A><��֖���^X���=��=�v�=Q'����p�2ǫ���K���>Y�>��:�2����C�>ռ��3�m�	��F=i�z5���l��ך�>pX4��x=>� ?i%�/�̾vꁿO^��0I��g�.?��?'�R?��F?��=5�^�ž�ʺ>̓?� {>q��=ST���>_�?����5�����!�>���?�2�?��N?�2���2�������Լ��Y�>@88>�b!>՛u�[]>�>�8��ǩս��o=O��>{�>���>l>�i�=_�=������.��|��Up��}�`�A���'#��������#��+9����(۾R�K�N'�zz�.Dq���G��j��6��>6]6?��?d��>M���!n>h�����iS�=}��`����O��{龵)�s��=D+[����a�����^�	?W@�^}>�i�>��<��=mCP>�߂��ў>w�>�|�=��=hl'>'��=�w����=�t�>�->��=����2����
#��Z3����<�4?�􄾻B۾��/��`��KؾХ@>m��>�G>�d5����w u����>c"�<��z�����T�_Nj>G�>��ۼH	
��-���L��!x�K��=S�K>-�d=����⪾� �>M>^�>�ž��g�4̫=%$�>y|?�$?�38>4��>ڐL>��>�r<>���>���=�P>h�>��>?�'?�N?��=ݓ{�5��=�&^��v�t��=~���;�Θ=g�ݽ_]9>*�=Z�:=*�E>Y%�=�s;Qo�=�,ڽM�>N?+?3X?�ʦ=�X;�y[������O>%��>AD>�ҍ>�w�>1y�>�I�>�g�=�����d۾绲�"�>�AA��_u��/Z���?�u>�Qq>a�b?7��>�lM<�ס=(��ܩ�>��!>I�>�(?���>�%�>|�;x/�	�7�@�C�*���.�@>�y�s9g��dǽoo[�/�X�n��z�<.��>-B?ҫ�>�Ś=;�ڻ��ۼ~S�>���>�~:��*Ѽ�ܹ=9��=���<odq>0�S�'w��-<(���|5�5��|���]�=�T��/dU=�:�ԟ?�E?��ֽ��轡�G��sԾ���g�>6�>��?���>q�)=�����T�deE���н�?0Tc?V��>��U�in�=�����{@�>� ?��v>Ӡ����1�V���{E���?��?��>Oף�&'H�2pQ���	��Fk>UҼ� >�B�?��W?�f���̺������W����'g=N�n��������J:��"����w�
�+¾&�D��M?:��?kz{�\sI>�y���k���8���?L�-�>S �>���>A�>�be=�>��|�1�mk�$�2����dW5>�J>Ӊ�>� ?Н�>�N?K�>l�	?߫�<U�>2P�>�>���>�0?0;?���>��=9[�<�a,>��=���,�q�����A���S��=��>�vn>�A���C= O�<���:� >2�t=s��=t��=K��<ɾ'=f4>Z�w=���>�o-?�>���>�%=�Ν�J|�BR>�N)>4�(��F����<Q��>L(�>OY?���>����@�2�(�x����6S=��S?��,?x�>�">2�>@����ɾ�n,> ��=����@پ3�btq��Iٽ^Z9>p̢>>>�I>Β?�po?�h-?�^|>��I�/﮿9Sa�c��>.-R>��ѽ.��>�>[����:�"J*�^D��\���@���׽�Z� �=7�=��=�g<0u�=�p>a��=i���W;; �X��q?r��>��?�7D>wg[=�>�����S9?��	�4sz�~=�<����/����I�=@<�;�?�.?�Y��e����w�D�{,�>ϛ�?��?�X�?���+5���Ǧ>��>	��> ��=H�ݾg��=1��Ar�<{�=��NF(�$b����=���=]�(��[��r�ܾ0�;�����\�{?��u��{5����A������&�sAо77����ľ�d�c�ؾ��@������T�K?���ھ��Ѿ(��?��?�v�<Mb�����
��SQ��@���I�or���f����qT����������LZ��L�������=zC<��������N���j��ؚU>n1�>�{�{��%�<�����x弆�J�[�/�l����ޤ��#����??o�9?�,����ƾ��C>8������>Ͽ�>��=t�?�Ec>�>d�H?(d?�Y!=�Q���A���K>�?h��?yr5?����n��#ݾ��߾j.?�1?��=?1���$��r�>��N?�PT?��?J`��}au�>=ƽ���>�m?��=�0 >��z>���>{
�bX�ʍ��#l�������=�D���X=�i�>�pdn==n�=*�g=z��=��u�͸S�b�?���5�>p(�|�پ �ýJB���{?�lؾXW>p�g>���=k�%��4���Z�%M�;�H[?�s�?��??��?\�L��6J�=�����>pۓ>�\=ŵ~�6��>��W>�R���ۏ�8R�)3?/��?H��?ʸ�?�v��hnۿݰ���ث�!�����=u#>=�>?Sʽ�l�=�9z<�)<��;M4
>g�>#^>�ev>��
>c;>��=FI��!��ɎͿB{��i�d��u8�(��
�1����3���a�(1��X���]���+H�, ��e;���؎������r�>��:?Ut4?��$?����|{=����@�
��=@q�Mu!��r����S�
��!ƽ��,��% �ʍ�0��:WܾB��>i���d���>�oG��N>���>v��=^��>�A>W�0>F�>�O�=���=��ν#�I>��=
v=� <=���O{��P_�(���x��=��]?"g��F�˾��0�\�޾W�O�6x�>E�?�>��>������\�n��>.o��j�>>��IȀ>�E�>�,==u���>��ѽ�n߽��L=��=�N`>m�Խ��Z�5V�8?>4 ?�.׾tp;M��=��?�Iw?f�?�)%>Q��>X��=��>�UN>@��>:�>[�*>�F�>Y�"?d)?T!?��=��d�JY�;r~<��P��.��T��"��$?����=H�ν=�j��<�	��h�=X,8>�0�<6�=z���4�>'L7?�&�>��>ph)��B���M��� �F
>"��<|��>��>���>���>�:�>,B> �`����྅��>�8>}�_� �x���޽]�|>�.O>gQ?ϓ0?IG4���1�T�[<A�>'t�>���>�J&?�̱>��#>��h����lӿ$�f�!���Y���;q�<���M����7Ξ-��������<��\>3�>/�p>EE>��>�93>�R�>fHG>�Մ=:�=Q9�;�m;]�E���M=G��AG<��P�E^���&Ƽ���������I�'�>��;�[4ټ�y ?���>b����E��߳�f5��w�ھ!d�>��?j��>��<?���<:���B�=��i�	K�A��>��*?��??����w����#���<�'>���>���>�\^=W�$�L���B����?X�?3�J>�%�<9�M��(.�7��p	>y��U5g>V-�?��g?zU��C岾�H�$R{� ����E>d����p��@t˾P��Q�I��u�������@8��]?bӧ?8>I<�]��CY��lk�[!��[���~8>)~}>�,?R�)>�Ͻ�a���E����T�;\{V����>���;rƹ>cY?>�?�a?�E?a��>9�
�j�>X>�]�>���>W��>M�+?���>1`s>���>�7ƽ4��`�Ͻ�r0�d�:�j߽�l�=]{=B�=._d<+g�=���=P��=xr;��)�ý�^��N>�7�=�>h<>�e?�m)?Å���p-=s-
<����{>2˼�&�;���U�־/��Ą�=��*?B�S?�V?�cO>2nپ�������>.,?��??3$?$ 
>=��=L��}�̾�'�=�#>)E�=R��-\����O����L>��>Y1�<a]'>�:�?b_�?��Q?�G>�& ������m�o��>?��>��]>u1�=I�q<��=�I�9u_���q��Jb�t�S�Q#��w���U=\��>U@>Ӌ��&�>�i�>+�t���D��!;���<쇭=�ѝ>G*?��=DG�<Ю0>�*����R?+:�����a�=�wȾ"M��(n>5�=|+�<8?[����;��dW��˼��Y�e?��?�?�g?k��Ѷ��/		?�;>�>i>�=�!��E:k>���i8½�uR�I�����þ���=�B�>��>�>`1����;C�	�ο�~�)>�e۾����t��,у�k��;�{��BF��+}���u�  �֘B=r䋽�񚽗 ̾o��� ޾4Q�?�h?�Uֻ��3�yB0��E��亾*�>-T��^�i������h�g����վ�־�h�m�T�"�3�����{=�篾����:��X��E���-�>��F?4�ھ���,�{�C6;>F��>N >�V|�0ΐ�g
���ш=V�G?�E? �I�9��BL���>v�:?�;?���=Nyd���<���>0�q?PI ?��>4t�bu���n>
�?⛟?c�?z�/��D��Ya�,u޽��?�t?�A ?`�ۻ�1>����>�kk?�$q?j �G$�u':�þZ�?��S?n⹼��>��>�6>�`A><��֖���^X���=��=�v�=Q'����p�2ǫ���K���>Y�>��:�2���ӯ�_yn��y��ӊ��h@��W�=]B!��>���<ֽ�F+?��=J�Ҿ�}���N������~X?6��?��F?�� ?�"���J#=)97����>4>!q�>��-��S���&>(N�>y�ƾ�P�7����4�>���?��?��>?�qn���¿��U/������h�=1�=�RN>]n���<�=���<�߇��׮��*�=�$�>���>c�U>�(>�� >v�>���y��밿=8��|4j������#��I��~�������!�LϤ�c���b�,|{��l��n���7d����=����>s�3?�D?t(.?8�m�y6q>9TϾ��
�Ur�Qz��������i��3��=�Ҝ���{�Qb&������b��Wל>B˦=���n�>�{=z�8�B�>��2>��=�<7r�=��}>���>���>W�]=79K>#�$<=C9�=�1���@y	�4H���OQ>�B\? %;���޾��8�+��K<꽓N�>h"?/=�>6 ��o��Wd��y�=Y=�O���ϐ<���=s`>]T>�J���N>��*>�Ǿ/=��օ���G�>aޯ>jY>%�͠k�2��<��?�s��>��=�~>�۞>HpS?M�0?�0*>�^�>��>,{�>��>D�>t�>`��>��	?�=?Ģ�>�8�>x,�=�
_�4RH��gn=���
�\wq=E��;��=�s����/�=��<��=X=�o=	�>��n�<LD"���?q�4?��!?�u�>��L�8�Q�X�Ӓg��%�>��=E	?�q.>�9�>�{">�`J>BQ�>S���Ӿiо�?�:r��W��������3�N^�>�ի>'�<?�%R?����*w�c.�>d8�>��?]Z�>`��>)�`=�r5>؁�>�w��)��̇/�V���P>��ĽZ+M��M���b
���A<�2Ҿ�����=�D�>Hy�>�zA>��-���/=�P�>sY�>/�q>�OY>�.;=�y�_�=�����>J�����ի���@*��*y��*=��G�aX=�����d�=D�=$O?�_?�/�x���A(�3��;6���P�>���>u��>���>z=)k��+F��D6���ؽ9}�>m�X?u��>��D����=�ýyo=���>3��>f.>��"���,�ҧ�H�T�Z��>��"?�:�>"��NO�vgj�ݰ��>EUD�dw�>;i�?��e?_��2�̾LN�x��5]2��0�>dl��Z-��Z�����5 ��]��@��Γ��R'��{?ݨ�?�(ͽ:9��D�fQ��s�y��H��eh>���=�1�>ʮ�>tT��d��t�q��$�����P��,_�>�f�>a��>�4�>X�?/��>y�>�>?3� �Q�	?U=�D�>�wd=��>�R?�A?=��>Υ�=�̎���t�I0�}��!�1�;�)���<ۙa=�>�/��9U=X��:%�=FԊ=�UW<#RF>#&�=y�{<�-�����@�=Ζ'?D��>���<? �>1yV�RW"��Y&>���I�>��I>�\�<��<��=�?�o$?�>�@T>^E�LЇ�$�Ͼ�x>�)?��@?��>_K�:�C���N��21r>z.ʼ�ua���˾y������� *����>l�=��U��u�>6΋?�Kd?���>��	>�-���Ţ�W�D�`-�>+�>�?Z,>�p����ƾG�������W�uiR��ٽ�W;��2�ksa>J"h>��>��o����=R>5�þ�齹M�<��\�bJ�="��<K4�>Ē&>�	5=!*�;���<V?�D�Syw�#5�=Օ�n󡾭�=���D�>1H"?�y=lsg�<ڿ�\b���?���?�2�?#~?_��
��[�D>�W�>�k�>��v<�������>�ƽ��=!��=����~���-�ܽ�:_>[�>��z�գ�K����k������Z<�l	��XIx�p��Jڪ�;7:��<n�|>��N ���ֽ. ��@��>�{�\�������}��q�p���'?�g?}Fn>��>ZO����\�1!=wzȾ��T=�0�*��z�����~�ϩ$���Hw�WI�� ����o����]�.�H��l~����ဈ<��c?�g�T��o�۾�[�=�@g>C����!��䘿��Ů>�Z:?�By?�cV�c�w���"�ά>N�R?I�>��?���h���>�a?!�f?���>.>��r���p�>q�?�v�?�4?=,��B�s��&��=lW?�j�>�43?;��"վ����+A�?f�s?��?/��怿����QF?6�? 	�"��>���>�<�>�/�:f���<~;ԓƼ�	Ƽ`u->�]�=��ʉ���#���r>?��>�b�>9E��ʤ��
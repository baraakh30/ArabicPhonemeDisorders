�   �   �?j�����H�H���sH�pn������u<?���v�x�cm�>��7�]�.�4$�~�0�J��>��>��??w�>س�>0��i�=�Ld<�{�%� �{�<���>8|�;9Z<2E�;�h�@AS�7gŽ����)�=�=)��=�=�
>H=U?��?��>9hQ=���=1 ��-����%P��������^p>�"9���E�:�R�iHG�cT�(fL��䩽�x[>�X��.X�=�ǡ=�"�Ӡ>Q�)��=�	?>���=C��=N�>i��>��>�f�=gQ=a񒽣8����޿Ht���s�C!���,>8(�>:D>��:��4�=�%>R���;IY�'�)>pc�>�N�>p��=�+<�n<#Q�|��"�=��l�'T	�sk��M��p־O���Ճ�L�����W������A����# ��h�C�8������\'��Ip>�UD>�#�>L��>Z?��>�l�>�b���;?�1�>�J<ό2?�`�>*�?�)?��>g>�x�=yt��;�3��^��&�<�|@�R��=���>t.>J<��i��=Cb�<6�=�(<JS��]rG����<&!7���=��6>}��>�/?]}���:�E����M��=�8�RH>lA?5�:��b�>��>5�<��aF���?�i����1�>wD�>KC?��>��>"�"<�Q�y=;t��sU�> p�%��=o�k���b��Ǎ=��3��@	=o�x�F�W��=ւ�=g�=��w=�%�<nB?�?��>N#S���"�z|^�?�H�8��S9�a�ž��>w�[=�v�W��!�6�o�O���Q�����.=�ux>�S�=�q�=T�H>�Ĳ�;�A=.`
=��!>BDܼ-�M>��q>�e�;
�P>��=�Q�*,��ۓ�0���ٿ����>G��
���Z=#�m<4-�=�E����=�#ɽڦ���T>�)�>��	?���>>n�=��>>Lu�<UIR=X�þc�������ŽL�����a�5�%��觼�g�m��,�0�Zm��]_�w�)�%㊽n�r������.̽Dі>��>C��>��>cD?ܜ?�p?��=bo5?C��>��n>���>߹�>D�?h�>FsM>��M> {=�J�2�����ٱ�=�)��4&{=ύ=>�$=;뽁�Z>�9+=u�>��?���A=��\=:rI��f=�ٷ=�H=,M�=��0?Z%��*��v��Ao�����o�>uiL?�NU�5�>(��>g�����,�Zž�FR>@S?��.?���>�.�>���]i����G���z>�َ=���>��H��d�.�)>V_E��������ƈ<���=��>x4�>\R>jKS>DSD?vN?��><E���j���G� $�K��=?	׾hz���/ܽBL=l�ཌྷP߾z'��-��!���ྔa3���>C#T>��{=�>+f(�h����2��v	��½et<M�>>|�>���>"��=.p=m�;�ج������e¿�����	������>�^�>��=+l����>��>V,���V>�Z~>Oc�>$)�>O�=Ah�Z��C��=�V�S�@���@P��2�꽥Wf���t���G��1��t�e`T��/%��%�ۉ�
m�Q��^2!��<�,�qk�>�s�>:�>��>]r?��>��>�9�)��>s]ؽo��=��q>vl�>�}�>��>��>#_�=`5��k�ߞƽ	��)��<�ǥ=.��<�D>�N>~�R�N�H>[*�>��O���/>�=p><0q>=~���<�x�=���=3u|>���F�@���!�S�Ե*���>�%?��4�W�?�:J�(�������2�����I�>5�?��?f-1>Ӎ�=��E��Ҽ��~�}ݶ�>��:�w4�n>�4�=Α�=-��=l^�����?��N�= �=��>u�<N�D���k???��k�3�v=�k��j�O�q�'�}��<)d�����=#��=Mm	=�*��UB����3�]5�Z`V�h�@��'뼐-�> �A>�P�=�T>?�����y���B{������P*>&}�>�5�>���>��>G��D� �6�jg}�Ƞ���}��k�jS���~�x%M=`ٹ:%ƽ�@����&��PC�/)���m����=Q= 2�=�֫=/��<��=VҾ��ɽ$�l����5Ͼoų���B�v�ɽ����oM=ծ��	�^��d���|�@~��")}�Z~��4g��U�<���>f�=��>k��>�)?U?�?�>%"���^?%\���D<ˬ�>x�>�&?�?}�=�t����	=Y�Y��� >���y�Y�x�>U]�=��>�Z>��>��~�=�{d�e���r��=ߵZ9_z(=�X=��=���=�4�=�j�=��0?Z%��*��v��Ao�����o�>uiL?�NU�5�>(��>g�����,�Zž�FR>@S?��.?���>�.�>���]i����G���z>�َ=���>��H��d�.�)>V_E��������ƈ<���=��>x4�>\R>jKS>DSD?vN?��><E���j���G� $�K��=?	׾hz���/ܽBL=l�ཌྷP߾z'��-��!���ྔa3���>C#T>��{=�>+f(�h����2��v	��½et<M�>>|�>���>"��=.p=m�;�ج������e¿�����	������>�^�>��=+l����>��>V,���V>�Z~>Oc�>$)�>O�=Ah�Z��C��=�V�S�@���@P��2�꽥Wf���t���G��1��t�e`T��/%��%�ۉ�
m�Q��^2!��<�,�qk�>�s�>:�>��>]r?��>��>�9�)��>s]ؽo��=��q>vl�>�}�>��>��>#_�=`5��k�ߞƽ	��)��<�ǥ=.��<�D>�N>~�R�N�H>[*�>��O���/>�=p><0q>=~���<�x�=���=���>������|�G�:SH��L���>���=aP$�|J�>��,��#,�Fj>͐�=G�	?Ԧ�>Af���>�B�>H��=������Y��)t���=�2�Ӽ^*D<���=�I���D=������X���6т=�W=����:>Bǜ=x[?@4J?:�>�k����� Wj�Sc��8��=g{�<-�D>��>����( �ǒ3�W�A�fK�֧ܾ�^�= �ؽ<_(>ʿ.>���<h��>h�;�θ=m��=�u �)>*�>�z�=��>�h�=�T�=��=>)�;�,7�m�����s$��ߤ�H.���X�.�پ�p3�oLҾ�Oٽ*����S��h����t;ا�=�''>�Y>�%�<�>p~�=�F���P��N7��`;=��ʾ�龮�Ͼ��v�����6!E������S�H�侇���,8������{��~9��n9=?ɋ>�x�=���=�u?�DZ?�D?��	?�M�>�?��K�?�� ?��/?�x$>E�>��սFQ��6)W>���6�I���E����nͻo�D��=�G�=��s=���=d�$�/w�<Qx���=J!�=�T�=zn&=�k=ש9>H���s��>�yk�t�5���������P�y.�=���=���-�o>	jɾ`�޾��Ѿ����3q=
��>���>��>u%�>k��>=�=L��|;��������D>�gt>3��<��0������y���6�Wݢ���z�Vֶ=��+> �*=�t������>1�B?��1?u	?6���,�v��e����8B>��L�+�>�}�>�*5��㦾;s����.�ߓ��x� =�K��3E/>4v�=���=U+=><��=�G�<1g
=id=׼ڽ�X>W�D>>C�>V#>Fc)>1���B�
�0��^����ܷ��>��D�A��_��=h��<Y�D5��"�П��Xu�����QM�=��|>3�.>�uS�`$�� R=�����ھ��j�a>糮=D�ƾM��'��=����px�����&ׄ�!e�s;������[g��A�SĎ�C�b=��>>#2_>��2>��>�.E?F4?���>J�)>���>����D[>~�5>D�?Z�r>t��>P�^=y�*>Q�h���?��݇�㑎�
�;=	���Te�=l$�=Y��=E��=�)>7hI>jR�=�4<>���=���=���=b�ʺ >�9�>)�Y>���>���.�$���+�A��jݦ��%O�Zi�>�w��z�;��%�n�#��M!�c���ddx���?�?�$?�x�<f��>��p>!"7���Z�;-W�d��<��>_i>���=�n�=f�����*�����<�z<�y�=VЬ=t��=�Fͽ%A�>�81?XC?�S�>��þv��H�#�����=N&>9-�>���>����H�'�ي����5�"E���w��"��O�h>B�H����� >�q=��3= �==�=�����{�=�F=���>���=YRp>�J��ýc���I��x,տh���}���.��b��=o�>��!�@j���8]�Y����  ����l=�kg>�5\>Z=wI���Ʊ���=�Xʾ�?��s�D>���.���;�����D���B��ý�\;ͧ��sо��R�/?�������0��ս���=.U>���>��=f�>UG?
7??WJ5?���=�c??أ<D��>H�z>#&?o5>�P?cΙ�Y�Q���� �
o��� y�Z�K=u>�A�=���=Z�>�+*�,>i�PЗ��
k>� �=��Ùۼ�,P=[,���=\BZ>�k>s��>�yk�t�5���������P�y.�=���=���-�o>	jɾ`�޾��Ѿ����3q=
��>���>��>u%�>k��>=�=L��|;��������D>�gt>3��<��0������y���6�Wݢ���z�Vֶ=��+> �*=�t������>1�B?��1?u	?6���,�v��e����8B>��L�+�>�}�>�*5��㦾;s����.�ߓ��x� =�K��3E/>4v�=���=U+=><��=�G�<1g
=id=׼ڽ�X>W�D>>C�>V#>Fc)>1���B�
�0��^����ܷ��>��D�A��_��=h��<Y�D5��"�П��Xu�����QM�=��|>3�.>�uS�`$�� R=�����ھ��j�a>糮=D�ƾM��'��=����px�����&ׄ�!e�s;������[g��A�SĎ�C�b=��>>#2_>��2>��>�.E?F4?���>J�)>���>����D[>~�5>D�?Z�r>t��>P�^=y�*>Q�h���?��݇�㑎�
�;=	���Te�=l$�=Y��=E��=�)>7hI>jR�=�4<>���=���=���=b�ʺ >�9�>)�Y>���>���.�$���+�A��jݦ��%O�Zi�>�w��z�;��%�n�#��M!�c���ddx���?�?�$?�x�<f��>��p>!"7���Z�;-W�d��<��>_i>���=�n�=f�����*�����<�z<�y�=VЬ=t��=�Fͽ%A�>�81?XC?�S�>��þv��H�#�����=N&>9-�>���>����H�'�ي����5�"E���w��"��O�h>B�H����� >�q=��3= �==�=�����{�=�F=���>���=YRp>�J��ýc���I��x,տh���}���.��b��=o�>��!�@j���8]�Y����  ����l=�kg>�5\>Z=wI���Ʊ���=�Xʾ�?��s�D>���.���;�����D���B��ý�\;ͧ��sо��R�/?�������0��ս���=.U>���>��=f�>UG?
7??WJ5?���=�c??أ<D��>H�z>#&?o5>�P?cΙ�Y�Q���� �
o��� y�Z�K=u>�A�=���=Z�>�+*�,>i�PЗ��
k>� �=��Ùۼ�,P=[,���=\BZ>�k>b�C?��D=IX&�n:��۾�D�(00��3	?[���@�|�������=ڕ��[�����>ݾ���6½���>�m\>L�=��]	�=-�����7=�n=�(�=D8��7�<��0�u}�;E��=}�V�^"�NA0=믤��q>�F=f��=�C?�tb?��?�T��Z����Z+�$L@�z���nξV!�;�D>xM<Hf!=��쾚�����]�6�NUо戠����>]0>����*�>L��<(�\���H>j�w=�}�=[��>K7�=r�m='~�>=? Q�=})M>OF���F����ƿρ��uyY������
��;Ŧ�����0PоU
�{�.>�
��vtξ�&��5��=&lt��
�={�a>s]r>��.>�輋�轿�<��o=�t��-���{���z�����|�o���BN�4��߷�ųp����Ď��3\�F��k_>wӴ=���<��>�zG?��5?�?�R�>�+!?9Դ>2�>߃�=�o�><ʚ>�/2?}�>�C?�j�>��d��9�W�
�e�Y'=����U;ݖ}>%n�=h>N�K�հm=GH�=�fe��sҽFk��G�W<��-=bvA>��^>b�C?��D=IX&�n:��۾�D�(00��3	?[���@�|�������=ڕ��[�����>ݾ���6½���>�m\>L�=��]	�=-�����7=�n=�(�=D8��7�<��0�u}�;E��=}�V�^"�NA0=믤��q>�F=f��=�C?�tb?��?�T��Z����Z+�$L@�z���nξV!�;�D>xM<Hf!=��쾚�����]�6�NUо戠����>]0>����*�>L��<(�\���H>j�w=�}�=[��>K7�=r�m='~�>=? Q�=})M>OF���F����ƿρ��uyY������
��;Ŧ�����0PоU
�{�.>�
��vtξ�&��5��=&lt��
�={�a>s]r>��.>�輋�轿�<��o=�t��-���{���z�����|�o���BN�4��߷�ųp����Ď��3\�F��k_>wӴ=���<��>�zG?��5?�?�R�>�+!?9Դ>2�>߃�=�o�><ʚ>�/2?}�>�C?�j�>��d��9�W�
�e�Y'=����U;ݖ}>%n�=h>N�K�հm=GH�=�fe��sҽFk��G�W<��-=bvA>��^>�?hIH��ʾ��Ծ![�-����+���b�>�揽����u�#�h0��l�!���������]���S�Є�>g�>=Rw=����䊼waj�6�P�=y��i�=6����-�%V����uy=��R������׌=ԝ->{�<���=�O.?n�9?W�?{t=��+�N��2f���e��>�z� [꽿F�>��8>�z��f���f��"Z@�w��D�����f>�1P=��<|��>z��<-郾�2�=�#�z�<<��>��>��_>�p>�W�>!p�=�K�=�Uد�
Vѿ�B���%���|�9�Bm�=�Y7>T��D�=.oX�u�M��(x�.���'�=gg�>��>R�6>�=>~>�ل������09�豾��n�%ב�/���qF�\��LQ��&�D�'���dTs��`!�����b:��uI�@e��R>>P�z>�ڲ�E1>d��>p�^?��*?=y�<��>6q>���>"�>	͗>z�>�0"?}?�jJ?h3?z�>ټ��8�\����=c0�=��=I��=�)�>��;�ʣ=�!>�D�=mK�;<I�i��4/���|��Q3<7ʩ<s�>�?hIH��ʾ��Ծ![�-����+���b�>�揽����u�#�h0��l�!���������]���S�Є�>g�>=Rw=����䊼waj�6�P�=y��i�=6����-�%V����uy=��R������׌=ԝ->{�<���=�O.?n�9?W�?{t=��+�N��2f���e��>�z� [꽿F�>��8>�z��f���f��"Z@�w��D�����f>�1P=��<|��>z��<-郾�2�=�#�z�<<��>��>��_>�p>�W�>!p�=�K�=�Uد�
Vѿ�B���%���|�9�Bm�=�Y7>T��D�=.oX�u�M��(x�.���'�=gg�>��>R�6>�=>~>�ل������09�豾��n�%ב�/���qF�\��LQ��&�D�'���dTs��`!�����b:��uI�@e��R>>P�z>�ڲ�E1>d��>p�^?��*?=y�<��>6q>���>"�>	͗>z�>�0"?}?�jJ?h3?z�>ټ��8�\����=c0�=��=I��=�)�>��;�ʣ=�!>�D�=mK�;<I�i��4/���|��Q3<7ʩ<s�>uq?�tR� =�����^�����������>��Ӿ���-|W>�pʽ4)����v�
'�t���h|������>/31>v�4���B��Ⱦ��w�	�������>W3<��{���q������fYe=�����Ƶ(��f&>K��<\ۼ>��R?(�(?�?�x�����o@�Ud9�y�Ѽc��=�ɽ,�>�i5>嵜=�!�<��C����
�O��!��;lL>�=�&>�Y�>�D�>�g�9T�R>��>lҺ�>dy�>H:?�5߽
?ZX�>έ�>�&���~���ͿB5����������C��Fֽ;��=���=�;��>/Aʾ��u�4�+=`�i>O>�6>���>ŭ>;�=>F�_���y���z=�<��+��.7���Wu��a���MY����(�^z����]������U�\sǽK43�?��$�#�?�Q=�a�>�r1>W��>��+?��]?��4?��[>��
?�J�=P3&>	cQ<���>܋�>M�?ĥ�>2�"?Vw	?P��>6
_�V����=��h��S�=h��<�ER>�r\>�:ͽ���=!�=fuȽw��"  >߉�=�3�(��<��G=�2�=�]?��:�J�a��&����D�>\��>�$�=���=�>�K
�65��;���:�?��?�<�>��2�>��=c�+�G��=�7�=�E'=j��O�O>00�=�&�=(Jr��v=ۄ��Ox�٬�<7��=�P9��G�|(��,�콖$?S�?���>w�������Q�
�ξ�f���d=_T��֌�>
#>N�;L����~1�G$������<7>wmm���X>.�w>n�y=�LS=d���=���^����;�r�=@V�=��D>i}=���=�Fo<gk�+z%<5S�=���>�|���v�,!�
�8��<��=��7����0=֋ν�o���r=��`>@�=���=�,X=g3�=���>j����̾Tj��q�� ���^�׾��;���;с��γ;�4��������ؾ��T�i�ӾP�[�Vy��Xd=Wz����<�ٳ>-�>>��>�!?�?B�s>$�N>|��>4 L�D���m�=2��>�k�>\�?�I><W�=*{u����C�;@aԽ�\=�9�=�g-=��$>P�>L��TY=c��=�}�=:+=�<k1�=�r�=���<
�<��RW���>��P���"Ծv*���̬�"��>@�?��p�>yǽ�`>'��2n�A7��ࣉ=�i?�F�>H�w>�Dr��i�>�Z�����>�<l����ɽ4��>�S>�RM<�YμZ>>�ZJ<�zd����< ����>��>͊׽;p=�r=>��(?u�?��?�{�����m������=BM6=�e<�>&�x>��=�[���x=�h��T͈��Ф>����ć>Əp>a�=�q�>C�=lZe��I`��@)=Z�켑s0�q��%=_�]=��1>-󛽑2����~=93����l���i�
�S��1^�=��v>����1p� ����=��žzc��^(<�i�W)<��ҽi	����������
��w�u���==��Ǽ��.�'T5�jb����w��{��ì=�7���vܾ��`�Z����+���&���L��нD�\�f�>�>YX�=�=�P�>��4?� ?��ּ�t�>�b����"=*x>Sb�>a��>���>��H>�\>!�ؼ�$�;h| ��y���>��5�u����=��G>�+=���;�k�2*=���>Ӹ>��>$��=:
#<��=�=��>��>�D�곾��/�w��\1���n�s?�>�۽jE��O������L���ɾEbϾ�Q�>5g�>�Q?9?��>�t�� =��<M�T��3����	=��$>�K=x)�>�o=�Y>��A�/�>�N��A�82>�
���!>�3>z �>�	@?�E?*f�X��Xm���㽑qڽo���ݦ>�(��{u;��Ͼ�:��v�.�7���[���58=۱�-�>6��z����P�>yߡ>��(�7���PN,=����¶H�ξ��q�R>
�<Iw�>���</U��̉=k�0��	���b�O�K��⢾���ߞ=�3μ]"��R]���J=4��Y%��G��1�=���Z=)H�=�|s��4��'���7�K�5�>}<2=�m�����?����:�����>J�;(��]�=O�l�uz����m��d�.$p�?�׽2����Z�!?!*���=X�8?-@?a�4?����,=A>�=X��=�?m��>�C5?p�N?��D>�O�=����O.>q{����2���U>w4;ע����9�04[=sN�-�=k� ;��>�E->�#=o������P�=_��=�9�<׾���?W�����+2��}.%�������>E? ���Iὐ:�>�Ib<��H������A�>	K?Nt7?�F>;�>�`�c��=T�8�Pq�����>��>��m�4�ּoKF>{��=�$ʽ{Q_�Au�ӫ��R���μ�S�=��\>?~1?h�C?�c?����6Ms�dM�c,���a�g�=�☽b๽ ��=/�	� [�5m?�[]C�&}�mUm>��M{�>q�y>%��ek>���=�"����=���=X �����i�<",�<��=�ǈ>䷮<�զ=����0ͼ.o˿d.B���E�k�n��>���>�\����.��	�>�;+�*���Ѿ���=9�=Q	>�D>�K�;ߜ�`E��L��3�*�V�߽��Ѽ�h��y�)\��RP	��t2���佅f�������f�� ���]�n�ͽ|��{�#���,>RU�>:��>�)P>y�?qs:?��+?8A>�J�>�Ԫ<C>s�	?� ?�2?�#?�?�>���>ڜ�=�Se�şZ�J�^�\P�=J����.Rn=��>bh�÷z=�6�>��<n���}>��Z>���<�$>�B�=#A�>���<�w1?uSѾY�ȾJؾ���s�Y���ͬ�=�Z?�� ��%���R>je�O�$&�h^�����>}#?�C?9G��ߑ>4��=^O��Z?o��V��!��=�i>9E>�Խ"q#>�<>
���m�'TB=hg�Y;����>H�=H�8��U�>1@A?��d?��?n��=�qԾr<��츾�=����j�Թ�=��1����E��j�B���6��{��>Be.��9�>�[R>��׽:>���=u<s�3��R5>�o�q���q�=9�>,�=��<��`=7���c�<t��=En࿧쓿T�e��kq�L�0�Ьt��%���N��ے=y�j>�&��C&>���>���>5��=�1p���ɽ+�{� Fٽ_-E�" �7˾�;�<5*�}������� �;b�D����]~������Y��g��`����N�4������<�ѵ>_�4>BR�>CM?r~j?��>q ��ț?(y>>eE`�d�R>%�>���>�t?���>Ս>�yM���=�Q��ۄ���ؽE��=��m<k�=�>,M轪pL=	̸=��=NcR=�=a�=�A4>��2=���=�/�u�=U;&�����v
�%��6�����'��Cu�>��7�����6㾳z-��S�2�����k@5��M������Qj>0L�>E/�>׵����<���<�}���pO>�$�=��n�#��z��.�}��db�d��AUZ���S�-���o=�8�<��e?�,<?ڗ7?�h��� ��z���h��Ρ������w>5�v> �t<����-��0ƾ[�����þ����)�W>�?=�F>Ve�>��[��S�=k�=b�J=�ʲ>m��>ǇV>ݣ�>bʞ>c��>���>���=P����㲿g����Z�]/$�{����9�a��Ș=P�=�N�ủ��:�v�H>�R~>U{|>�C�=�.��0��q�5>���4��j�=�|F=U��)� ���þ��q�Tf �:}c�RM�ݙ��zu&��T�&ӕ��)���E!�ϼ�=	t�>=�=��_<d��>y�.?��?
p�>�]�=E�?c09>�b�>a��>�\�>���=CJ
?'�?B�?6�?[|<�R��Yw3��r��k �o��<w#�=�3�<��;�*==B�=_��������57�8׈=\C�=�S�<С�=$Z�=U;&�����v
�%��6�����'��Cu�>��7�����6㾳z-��S�2�����k@5��M������Qj>0L�>E/�>׵����<���<�}���pO>�$�=��n�#��z��.�}��db�d��AUZ���S�-���o=�8�<��e?�,<?ڗ7?�h��� ��z���h��Ρ������w>5�v> �t<����-��0ƾ[�����þ����)�W>�?=�F>Ve�>��[��S�=k�=b�J=�ʲ>m��>ǇV>ݣ�>bʞ>c��>���>���=P����㲿g����Z�]/$�{����9�a��Ș=P�=�N�ủ��:�v�H>�R~>U{|>�C�=�.��0��q�5>���4��j�=�|F=U��)� ���þ��q�Tf �:}c�RM�ݙ��zu&��T�&ӕ��)���E!�ϼ�=	t�>=�=��_<d��>y�.?��?
p�>�]�=E�?c09>�b�>a��>�\�>���=CJ
?'�?B�?6�?[|<�R��Yw3��r��k �o��<w#�=�3�<��;�*==B�=_��������57�8׈=\C�=�S�<С�=$Z�=�t���|����n=n[#����S9����^>C-��^��v~�>!��hV��n������-̾����Bɩ���>TSD>�m���E��
�Ǽ��=��L>+�L>$���=IU�=�&>�QĻ<?�#C����x�<Ό1=��d�K��=1�G?�'?��T?5ʵ�%l0�����h*�|�о�ٛ���H>���� ������=£Ѿ��_�@�S��ǈ�xZ��[q�>���=c�<�@T>��/�O�'=Ԙ\=��=#�h��u@�p�D>�V>P�>�5�>�F�=Vu%��z�P���o��="���a`��X���!�o�=��貇���:q^���+��J��U�=,�鼊�<ՙ�=��9>N>n_�;R}��į��L=>���=R憾8��!ʾ����]ݮ���n0)�l�����Ⱦ�=� ��W����<���Y�f���s?c�g=�jy��ͦ����>*?4w�>C�9>��)?��X>��=bN ?�'?��>##	?ţ'?p�?�A
?[z�>���<������<��uD���>�^{�^����$>Y^�=b��;�E-����=#ٽӛd�>�=�{>S� >�>���>�1�Hm��>\½;]���4�.��+ �>��8��z�>�Y#>����#����6-���3��A��t>t��> �>�.�>*���Ǣ�f����M<=�%>ͅo��Ԕ<v��=]9J�F<�0=�h��ŻR��]߽��=�6k-<�N>[tp>��M?L
?B��>���;����@žK�����4�;�=�w�=�X̽�>��{%ھgz���������νg�N>���=��ż���=�/=�=V��d#����>@?�=�^�>6�>ߨn>��>�?��>��|='�̽�慾7 ۿTB���]3�8�4���
���*o�=F�=8+�čW�Qm��̮o�1������d�>Jӑ>�;>�;��=�y��	>�����A���u�
�G�DU����v�q�ѽT ��jĽFͽ�8!��`�V=����x��ܹ ���>��>1�>�
�>��A?��:?#[�>H&�b?���5��:9l�>� �>���>���>��?���>���=QT������u������=b+�=��>��S=�i=>�>􊲽߼�H2��A�E���ѽ��+�o��Q�=(ܞ<�m=��=�t���|����n=n[#����S9����^>C-��^��v~�>!��hV��n������-̾����Bɩ���>TSD>�m���E��
�Ǽ��=��L>+�L>$���=IU�=�&>�QĻ<?�#C����x�<Ό1=��d�K��=1�G?�'?��T?5ʵ�%l0�����h*�|�о�ٛ���H>���� ������=£Ѿ��_�@�S��ǈ�xZ��[q�>���=c�<�@T>��/�O�'=Ԙ\=��=#�h��u@�p�D>�V>P�>�5�>�F�=Vu%��z�P���o��="���a`��X���!�o�=��貇���:q^���+��J��U�=,�鼊�<ՙ�=��9>N>n_�;R}��į��L=>���=R憾8��!ʾ����]ݮ���n0)�l�����Ⱦ�=� ��W����<���Y�f���s?c�g=�jy��ͦ����>*?4w�>C�9>��)?��X>��=bN ?�'?��>##	?ţ'?p�?�A
?[z�>���<������<��uD���>�^{�^����$>Y^�=b��;�E-����=#ٽӛd�>�=�{>S� >�>I�>j�(�E0��ﰾ����K�x̡>���>��D��>��żXt�ŕ�^��©^>�q�>Y��>�Z�>>�>&U�>�]_>�Si���:݃�<�jϼ�2n>&*�=��<B>G0�<I}�����HK1��8��G�6��0�9G��;E�d>�P?�2&?�,!?�=�񾊍���۾�0�<O�z=�=f�a>�g/>;u��a���A&�L�� �4�g�or�<�S`=��>��}�=zS3>jU#�pF�=�0�=ǚ�Kg=5��=�"�>T	�>}	>t�=����-����νY�ٿ�ˤ�[�_�,�?�8�� ���~��fO�<������Q����'=z�&�3t�>B>�q>�R>0[�=)�=�∾�2)�Ӗ�*�E�Z���V&\�~��F�ʽ�x���Ľ����M��Ɣ�-���T��'T��<�<��*�ν5~�>yV?�>�6N�<<X?{J?{�>�~>��>=+�w�>�Q�>�%?<�D?F��>5�G=J���9G'��<m��gx�-Ls��[>��h>��S>�@T�i�
>(G�4�սXm�=��=�A>>��a�n�ѽ���_=E�:>{PB>d)>�+?�->���f{�5t���Z�L������>�/g���2>�U�z �FS/�״�G�>]=?N �>���>�;�>��/>OL�>��v�3S�=>��=��z� ˉ>��O>�n�5�s�(�";yH���P4���}���*��=��L=�ӎ=�.=��[>��$?��	?���>�\���Z���ξ�*��Ϝ���>y�>�;=Q�=�븾�'��7��sL�TW���H=�S8=�4>A#�W�8���j<�L(>���g���t	>�0t��`<�qQ>�v�>��o>W &>BTI=�����ߋ�6��M�Կ]_���x��K�	����`�,<�h�`�=j�:����=�q�;n�;퓆<{u>�=�
�HSǽ����N4�=N����]�n��=�쁾��ľI:��̾7��*�{�#=�=��޽�n$��)�-9�E�5����ƩT��9ҽ�b���M�>�D�>W��>)�+?�-b?)��>>�>ڮs=���>}��r=>��?��?���>>�I>������=�F�V8����Yl�u2>}�V>>��8=��D��ʐ�y�=G��=��(=��t��@)����;���<�=+�>�A>�;�=-۰>E�x�,����-��� �3�`��$�= �=����[[�>}v�\ཾ���=/��ý<�>v[�>�4�>h>͵>��V>�0�����؍��:!�X>���>_��=�P�;��f=6gνx?ɽk��; �=&E�;���;E�A=�?Z<:�=Ȗ
?�?�?V�>���v0��w=`����9ȾA�>��<Q��=��Tz�K $�/����	˾,u)��E���ep>�?���>��0>�6R��t �7���lT����r?N>Pm�>ԯ�=��=^B�=�z��{(�0Id�Djֿ'����p���nL��yӼqX8>���m�k��2�<�1���ܽ���=d<��>g�=Ё��H��:̛���h�>��߾m��hݽ�f����ξ�s��apɾ�M��Dg�r�"�ͨ4��Z>�~wW�b�t�>�S�����7�;A�>�?�3�=++�=Bo:?��?P[�>M���e?�?1���#���>�/?j @?��>�6^=Ձ{���d�B�Q���B�3`���Ô>�" ?\�=��c=:��=����k|=Է�:�O>�P�=0)���b=b�����v�R~v>=�>i��=�>?G0>����
�AnB�@���/��ZE�>�`d��/����[��7�l4x������c���_>9>�)�>�P�>ۄh>o|e>����\<9=�֩=-@�>#\�=1�/�!ww��Q�X�y��ߪ=�`>�o?>��=o-Ѽ�A���h>F�/?X��>�0?D��\L������˾��7�aϥ����>�=�8F<;e�1�����=�Ҿ+������d���Z�=�#>���=�6G>��.����ǀ==���>����p�=Z�=�r�>TZ=>*l=()�h�%�L=V�O
#>GvпA튿@6�!Ӣ�r>�5�������n��HW$��&��}@r<A�kL�
�1�ۊ!=�K�=m�#�b;�`�U��]��[I�cp�>ཊ��������]z��q߽�ӽ,�]�=u�0�=.�Ž�\A���'�2���s��Q"q��X����=2D�>')�>��L?�	�>K�>�N{��>>Z�E>9�G=�t>O��>��>�)u>�7ͽ���=��/����O�޽((F��M�=\q=���=XO<�(<�^�7�C=��>��>�-	�~��:r(��Q�潌yL����=�K�=90\=��?�3�Q��-��_�Ⱦ��\=��:��>�"��4�=��?��e��Q��n��G��!!=/�J=b�Z>N�>�'f>*P>����Ht�0>���=U�<dg>n�ͽC+�&�E���u��<���=�R>��<&蜽c��ۺ2���<��/?�"?̑K?fpI�!� �ڔ��i��w���o�9>J�v>ǂ��g��%	������ND־�ۃ��v�f%�ww���=��>>��	=�}8�¢���޼F���,=}���1��=:��=�;F>x��=UwҼڈ��$�~�����O�=M�⿻��dˈ�����d�C"7>���={�4��j½���~��$j���}��S>�O�={)O<w����w�=��F<�A����KT>.NP<ϧ��)	�����ս2 ��@+<����xܽ��;�#�B����_gA<,��+�߽��ڽꖫ=4K]>D]�>u�>��!?�C�=��%=2	�ͧ_>u_��>Պ>-�e>���=
�h>g�>��
=Y�Q���վ��O`1���>��=i�������<�>:�v��=�#^>��>>>��=��.�/����%���z;kK>�VP>�t=�go>���\�ݾ��8�󘞾[�g>��Y�K��>�v���hS>�v侕Q�Q-��N"��v���>B��>;?���>���>g�>j���rc=�;��j�`>iǼ`��<8�>NC��!��=�����~�Apb�#��rT^��r=�~=˦d=W
>�oP?X�?���>#�����n�x?S�MSi�V-��wt�R>�b ���==�<?<���<<�1����E�� �p7ټi�>�E��g��ٽI>��[����ԟ���ּ��>���=�>ی?�V)>*��>���=6��U���m۽Cyֿ[k������-z\�| ��s2��>��#��IO����<͉��6>�~N=M@�=�PY>�MJ=�5�=nJ�=��̼����4a���?=����(���;l����0�����=��־f����L��N-"��)��j�+�c݁�3꓾*�a�D��>)��>Cm�>���>�+?h�+>�<%?�=>���>{�=Bk�>�M�>9�>�>?�3/?H�=���Q6���ƽAQp��������=Aw�=pA�=��>&,�>0�0>��k=����!=���=ι�<o�<��4=$o�=��=�->���=�g>_���Y�
���u����>g���k��eb?<�i�ckݾ�tҾƕ:��P���4�}�Y����</��>�8?[?q��>Z��<���ކ>��=YE/<��[=2>9*�=���;�սj���9�g�k��Be���Ͻ�r�=B_�<��[>V	E<Zl?7?C�?�}t��#Z�v�z������} >}��>B� �ƴ��UE�>�S���8�Ø
�A����i�Š���=��>*���AQ�r̵���
=��9=|�˽4�>�޽�"��=�Ĝ>Y�,>62�>ғ
>G=������b"�q����KǾBy��D��N=�����4�Fp/�����(�T���To�usA>]�=����������rD��S�C����q=������v�t�@_�`C㽩���z�F�B�N�'ˎ<��߉��?�`X&��?���Z�����Ď?��.>W;k>G�>��^<9�>[2?#�Y>��?!��>��>Y}>���>�T?
�/?��>�I>�l�=?�X<�7i<J�ܽ�j:=�D<=�=~�m=��<f�B;)N
��E >�>D*)=�+��ޝ�=+��<љ
<.yn�P�=wj�=�#�>+>�=S2���n�!9���c��#g��%;,?<��5���5!���TV)�,���H])����=�H>�A	?8��>�*�>=j�>V�����=��=��=�=�#� 0̽|,�e�+>f|=���<(�t��q���ؽh=�jI>� A>`�A>��Y?���>��?�i�M,��[��}_��W��i=��?�l[>$ �����iϾ�Ro�����:�曾u�@� }�=0м�L=��	=#N��H�t�f�3<�(��D%�����2x>��o>M�`>c��>��=O%�#�=������߿ͱ��J�H�JJ㾕q�=iuN�@��<����Ǽ��J�2�1����f��w.>!�=-�>�9>=Z�=`a�=�t��*s�����<��{�j@�L��B���g�ʽɡ�����<����b����)�=:�:򽽬۽G�N�&�B��9�>�;��gH>���>y��>B�6?�Y=?K
>��>�Ø>`�>�"�=g?99?ߚ4?k��>�1C>ǳ;=�E,������4��E�=�V:����=ѵ>>��>>jr6=��=���M��<S���3��q���=�p�=Z3�f�]={>C�?��j�-�v��W�����K�d&Z���?ĐX���3�����Qw0<�������Z���>�$>?(4?'�><5�=�3W�ʅ<��=[_>8$>м8>/�>C���@U=�p��+ֽ�����#x�x =�A>�4�>�8>�e>*�<?�?�@�>�#�D��$I��G���=S���ū���\��>����.�=�Z#�6"��,������W�~�>R-���|���_��dS���7��	)��->8_>�k�(
D>��=N���Ɋ>S��=��@��۽��
пE���I�h��_žx�c�Ab=�[>L�5>�Z湂�j�5��w��f��=���>��>�!>��=�p�=0�E>�����D�h�>n�������*��;R����'��Gξ]��<wzu�� ��IȽ�������(�L����Ǿ&ц��Õ>��>�c�>Y�?M? K�>}�0?�Id=$Y?��[>_>?6��>��>(B�>�U�>��d=d~�>�弒vؽ�,H�p�P�6K�=5u�<5O�=��c>�m�=ɲ�;3��<����+>�=aH=#�>?3~=_ջ�)�=zH�=�h�=��>#o޾"�b��Kž��`��_�R�S�#?O�(�ᩧ�l�����8�2	)���b��*�>J�>)8?b?M�Q>�c(> �#�@�=�o>3=���=8�>8�[����O�<0N)�] �67Ǿ��^�!���0�>8��=���=윮=N�>��A?{{?uWn�9�1�z�G�.G�i�==�=��{=|D�>-��>�@����a�g�:��1)��v	��� ��</u>1' =�ϼ$ѼQ~�;I�����n� >��EO���o�=�0�=�Ѩ>1d>�,>�]：� �U*9��̿%W���!G=����޽>yj\<طӽ'�Ǿ�����=Z���:�澬]b�r;�=ݫ+>��<K�'���N�̽�Nv�v����6�=x>>��ִ�E��M*������賫��H>Y"��>'��C��,������4��ߑ�C�Q�����|`�>��?��������g���?MP?���>�n?	0>Ϛ�>�)\���>t�(?�@2?�S�>��>���r6?=$;
�mV�[�.9�ǯ=Ls_=�c�=���=Pܼ/��#ݦ=uJ>R��=���6��=��=3Gd=�=�=�|>>�,?��4���1�8�׻W?�ӷ�����>ȆZ>�O=�Q��>�*�������䇾¦��u�>�I�>�=�>���>�˵>�>����P�u���������'>%w>��s=������=�4�#͋<(%x=&�p�g��|�?&�;��<���>�]-?��>�o�>$R�>���"C��(Ѿ����nžIvW�r0>���>&
>�5N����D�F�����%�r�&gY>�Q>c\�=�t�>n�Ǽ����if��t�;~�=��P�0�=�>��Z>TF�>���>+��;g�ཧ�l�z�ֿ}.��
�*���P��|%�?J�>�؞=o�l���	>Q�	�	a��v�y��>�h>���=o`E�:|�<�l<�F���:�F�=Y�=E���W�L����H���� $���;brs�
.�h?�5:�������IQ�H�������]�=�?�0�>
_u>^?@?�Y�>ݘ�=
M>;�>N�H�֨|>U<�>G�3>~n<�f	>�=�uc>2X�=Np�7�&�d������=z=#>��/�˶0>Ez>v����y�<_7f�շi=�Ij=��iX���(�s�Q���M>�P�>g�8>#�?�ǽu�)������7'���<r��>l�m>����g�>�M��ƃ�L�+*T���>���>B�>�a]>3,�>@&�>�f8�t'��0v}����	>�>̯�>�>�##�sb>>��S�<���=��=�d8>�l�<�����5ֻ}�R>�B(??���>D<>�6E���,���پ�3�G~���`<��>-��>"L9A����z�	?�Fپ�=��v����>��>-�>,�>��n<��/�W]˽�]J���=���0{=-l	=��>]y�>�B�=���a<��?�;k�0���F�R��v���$=�Ģ�@u?�\��فn>t�><�=�J:I�� �=e�<� ��:	�=g�='v>�G�����8�D,�<��-��ξ�r��H"��R���(�iš�y�O�G�g��gн��&�\Tj���6��͆���
��X��>Q[�>�X�>̖�>���>�k�>��>��e>k4>�#���>{z�;��/�ٚG>?ց>���>���>CFּÇ�>ѽ�+7��B>�%>��̼�9�<��<�6�˙��Q*�<�v�=.ۖ>׶�;��#�\"��D�U��F�=�Q�>立=�?i��:nY��O��'��`��Wa�>�]�>9�T=���>j�)�6y����ܪ��;S=H"�>���>j�>Kʛ=ێ�> ���;���5G���߽��=�Q]>�(>�K'>��J=�?A>�B���=�$�<2&ּ���=sv�=A�G=�,==p{=>k�E?" ? �?�og>��ݾ)�/��z��������yCP�ݷ�>.�>
��;`����U)���9����R��n���q>>DBR>A>�t�>�v���hS�	�۽25߽%�=�����;����P,�=+�}>2��=m������]-�z�(����;��jc�/4=h��=˽F����'㸽Gv=�|">,+b>��=`�<
}+���E=��D>�p�=V�GƋ�K�=4�`R���j���.U��s_��_�ϭ� b��<P���2��6�p<�R=#���5��t&�WO��3�>��v<�>GT>���>�?t��>��=_Q�>Al�z(r<�m�c��=;�>d��>���>n�~>M|=F�㽄ӽ�,��"�=��=�+��X�$>���=|螼���=�\��* >�J>�>;1����;��ڽi��<�q>��>>�1�>���+W�>k��_�,��|��a"=��>ew��1��>�ԓ�=̔�� ;�ζ�� h����<\�#>�Q�=[�W>�c�>
�U=9���(x��bƽ�{7>+ž>�C�> J4>���=��g>�.����y����=�`>�>�4�>:�!�oC����>�q?(?3
?�*e>�%���1�N&���f�M���b6]�Չ�>W�>��f=�~��\H���.�\���>p�N���V>�Nd=�a��n>˯����P�w�2�u�%�$��x��'�=�&>^y�>�d�=㨽.%{���U9�ֿ v���	վLS�v�#;D�>�FB=�����]��v�� 6L�LP��k>:>6��=�ӡ���˽$�k���x=p���b����.>���=������Q}���H��ej��(�����F��jG�-$��4;I�-�p��霾!�X��N��{�>��O>�^����=�خ>S�>��>�޼>��>�/�����>�������>�L">}5�>�N�>Ǩu>�1��_&���  ��0�=�<<>$2�=���=$\޼�Ӌ�R�=��.=��>��g>#SY>�4��喾�P�q���z~�>���=���>�u��+����Q�O� �y���ַ>�z>(]� Ǥ>卽@k����Ծ����Y6���^>3 �>o��>���=x��>S"��ж��R�����
��Ё>ΐ�>};>J��@=>�瞽yvü ��<��x==b>��U=	o-��6s���>�C?��?�^�>K�>{8��v��;���� ��z���Y�>���>�R���ʾSv"�|DC�q�8)�=�x̯̽\>�3>u��=s>AIm=C����������=�����^�<�)�=�/>�#�>�g�=���۽=�｀�忽���]�*��C=���j<ə>�`���F���>c�����=��>C�S>G�=d~��������U��R�=�n]�Tã:���=�Ɩ<�ȏ���t���P�L/�'LY�8]��s��l0�˞g�!l�E�7��8�L��I��"�=O��>{�=x�]>w��>#F?Pc�>�Զ>��=�%
>�-y�a�=��#�Mg��\�>�#�>]>?�-�>��=����D����T�/H�=.N�>G!=�M�=[��ϟ��:�3>?c��X&>�VQ>���=�+M����.3���.>^4�>q��=wK�>��>�ܾһ��B�����y��b�/?+�R��m>�y��E
0��������|X��	^I=��	��I��i�>��=W�U����=���d�;�$�>AXT;o�	�7�=(o�C�<�������𐼝\ݼ�]=QM]>��ѽ�d�>0�?/��>�0.?C!D=֝<�!�G�R���ց�G�ݽ��<�0�>2�k>��8>�7Ǿ���P0�Y���/������Ā>r�!=À��Y]>0\�����Y�����>2=�um>�U>D�>F�>��q>��2>y>�=;;��=�o쿍=ÿmT���:����>3��><ٽ}�[��U���<�=���=Խ�g�>�a?k�^>Ee>['>�����*��q>�,$��@���!���ȼ��k�=�㌾eA��,[���f�W~�=G̽���Խ��+��l���9��������><�O>��>��_>Ru2?���>�L
?���"N�>�&N���>"*�>u�!�90>��	>;�=a�?	�?V��>�2ƽ�ヾ%oc=JQ"�=ǀ=1vE>�"W>��<�֧���5��ʢ�Z�ͼ�&�=��=I���\7�.�[=\�Qn>�ڱ>DR+<����$����>��m|���'>.z�>&���|m�==ء��?پ7.�o�;�>��#�8�(q�@T�;qֹ���>��>ŉg�r����P���>ٓ=E�>��: >��=�۾f�׼d8�,��xa��[����:M�o�b�i=|�=�?�"?��H?F
7>�9�L�h�t������e�<�ݏ>�/�>�y�>��!>O���rپ���-�8�~υ���ҽ��<>)pr=��l=��{>�c��3s�=��z�L��d�)��GP>φ�=O�=�Q�=h��=���==h>��&=����c���¿�kz��U�}m!<D�n>��<����
	�9u=�K�=<<��m���L��ߖ��(�=Pȇ=�M�>(��=à`������d�>��=��d���	�?�ľ%�O>ώ۾Y���c��DJ&�oU0>����;H�z�5I�������þ�Ӄ>�p�=���<�i��4�>	l?V�?1� u$?��ؽ����Xg>�{�Ws=r��>�1|>��>)t�>J	�>���N�j����<gR���f=�+���J��z�=�=L��=p�V>���:��=x���<	�>�:�<08����8>,�=X�>E��=�f�_�a!7����/�w=���>��Ծ��=^���D��y��t�h�����=|%ܾɰ��`�����>x�=�􉾻�����{�4���}ʹ<C�%=� �=:.�<���# �MK�lz���齚p༤���0�<��=WĂ>�M*?�	�>�� ?jE�9o?�A�>�����e��C��}�;>&̫>�_�<`����ξD��Vɾ���ׅ�i������=�	>�O��o
�=�l�=��=�5A���>�+�=QB�<ё�<ח>>a�>��=5�5>�ձ>�ѽ������D����%�ӾR��=j�e>�[���<�r��,�>Ғ�� ߇�R��>�����=@@=�\=�Й>�'�<��>L3�>���>�)>����>���k���D(=3�ʾ�}#>oߚ�Y�t�W+=n��7��c0�C|�.�b�wY3�q> .�;�>5	�A?�B5?��>�TϽ{M
?�M���59>pe>UN�@�V>���>oT >�?l&?j1?dہ�5(�����᤹:C͛=űq<#}�<Β=�켙j�����=�;�=No�<T�M����=N��"�=A��=�G>���>?E�=^uƾ����֎'�%�3_9>Tz?�P�=/�	=�s��R�ھ3�3�{^�Ǘٽd�<V�����a��WJ�2�>~7>ip7�X塚&#L�t����>E�x�;�(f����}��J�Oo>�â;�ׂ=��	���q�t�꼙Z>��?B�)?��1?��0>��$��v*��H#�6���G&���>���>�.&>x0=�4���⽻M������6���=&�>, ͼ����u�=-��<e�꽯q&�r5>�A=�V�=�}�>���<��Ҽ�J��*0�/f�=��=�t�;�ܿ}���3G��+���l�:�%>�M�>
�d�)����=Dgz��V�A5�=���<V
���Z>v��>E�?���>jA����/���]=i��=��!�휭��6����O=j ����<A��^�����<;��OP� ��C^�v�V�d�d�v�>��>M|>{t�����>޲?I�c>J�C>��>N���<W�>���r�>�s�>���^mN>�_>Y�r��5��2��,>,y=Q52>���=�>"�B>��X�M�Լ�=oĂ�Fӆ�����j�>����$�m=XK>i>q�> �Q>�ߗ���K���N��
x���D�>�ȽA�>�S���v����^��wP��H�\��%���m+>���}L�>��>��(�q��<��ܽ��������>=+L>j� >w�h<�Hl�)c:E��>�8=hqŽ-�����=g�Y=�"R>*{?4F?��;?����;�m�]�h��xݾ�ܬ�3��=�=>gc�>��=SþG���\���}q�����C;��o5>v��=���c>����r=ÐF<�%��挽|�=m8D>sr�<:�����<Gv�9��=���fb��[V�u���������۾ox<�k�=���<.@˾��0���M�RW<��2���O�������>�>��%>m_����}>+����K�wA)>g��<��N���d�*ڦ�˽�͹��-��!%��=/�B� :�����I�:����h���+��v�O:�>��`=9�G��'���<?D2?��-?���4f�>#�W��;�>7�>�L��7��,�>�C�>�Ӗ>�b?�H�>��,2w��X��ڼ�q�=��=���=�:�ç=�ؼi�r�߃;�5�ݼ~�@=��@=�>O��=�l='��=k�?cU���lھ����������h'�>�e�>n��>�o�H���zӾ^
L���.>u��>�V�>��>X�>su�>��V=2�S���ǽ��̼�E�=��>�\�=�Y>���<2��<u:>�̻=��hC��J�l"�<}|7>�{>�L>�G?@. ?T�?H��>|�ż��0�a@��`�<�/�K�>���>�O�=����iܾ��,�͢��*��zȾ�Z� -^>��>��=���=&�T=�����$ν�1�����=p$�<y>J��=���>*/>��I?n��⧾�˿s3�����K� �d����"�;B�<&<�&��=�DC>�뽇��=��=���=��D�5^�=	o���һ�v>�x׾���)�=�=,ɴ��	ݾY�t��{-<h_��M�=s �����]��A|�����d/�̚j�@�|�7�9������G�>�ݑ>�� ?AI?�z�>��|<8�#����=^o��3�a>�~�>�ѻ>3��>nY>�|>�>{=���:~)ż:;��E�&�ڙ�=f���l>02S=E>)��fGN���<�r�=�n&��6��C��=t.�=�P#=���=�\�=�gT=���>1���Ɛ��R�^���	��c~���H�>m,��^S�=
�)ƾ��޾)�_�+u>=�)>�z�>r�>�޼���>uX��tU�������;��->$x*>p�@��9�;��&��b<9�I>w�p=I߿<�%H������y/�ބ<>NO1>�RS?�?=��>���<v�����g�\1��u����>��>�>>>�7�"���J��B���9�0,��w�q\�=��L>R��>�L�N�N����o�<�}��#���f=%缽mk�=�5x>��>V>��>ڙ.����2˿z���eQ�����\�x1=��"�Y$��>��R�}z�f�O=���=�>��u>f� >:��k��`��=�.�=V8�>R1�>�<d����O���Wɾn��<ڜ��`H���r2���ƾ�;*�yR��?�l�#�=�c��l+2�Z^�=���>BX�=� ?G�?*7�>bA�>��;-�>����M&>1w�=L��>!a>�$>��<>��;�'�<P��9�l�|�;����=�,��G>�`�="'K=���<qIP>q��=���<�E}=��&��p���b=ݯ�=�c>A>�kV=��>�A�8q����7���P��)=X�x>�����g>;�Ӿ�l���~���$�����]I�P7Q>�%�>�J�>��>&/�=ZIp�c�=�/��&��=���<��-=�@>Qc=+�=��=�q�=��B=\꽎Qc=%TS<�hJ<{��=�l�>;%?5��>�D?�솽$���F�7>=�Q=�vp��>��{>]O�>h��>$y<�L/Ѿ�@��;)��#��L�R��:H>��K>�l�=�1>6�׽K��]Cn�g]	�����I�l>`��=�L�><L�>W���?A���zu��n��0 鿛ɿ*Ԝ�ʗ��ߞ�����<�>@z��G=	��>�������^�=�4�>�F_>��N>�:>��E����=�����N�=��[�� ��]̾�ξ�)�Έ��B��!��K����41��/���P;En½�������˘�#�����>P�=-��>v_b?�W�>�%n>G����>5���+_�>{�	>>�<o��>��-?L�>N~�=�d���8ؽ�����@�<&�=����%z>y>� ;>�@t<FT�=���=k�=���N����b;���x�I�g�'(�=�O>��;>��)?�*U�a��Ӌ��꾽����=�{>�bh�r>�+s����}��#�5����=/��>�n�>���>ޭ>w�x>V�=�����/#��u>=���=���=Y9��� �=��=1�J=���=�_J=�����K�n��j��F�K�P6x>L>�i?�U?_�>}�%>�1���G����"�E|a����=P�>��>�8�>걁������\>��=�~��Yܡ�%&e���=#,>�d>ػP>�
�=CZ��&�ٽ�]:�-䛾���r��c`���=@�>��+>×=����	ؿ�I��b�Ծ�9��<x�OI���������P��>[�=B�ӽ��>���>�~9>9cM>7T����<G���e�<J蒽+je�o�(=�캇 ��fM���@��+B?�9�2���=f�׽��Խؾ_�+\˼�:�+W���+��zG���>J�>��>#��>[I"?2��>�z�>B6���½ŵ���U�=�w4��x���{�=g�=��=��=�)=�5N�ɽ0�-�O�\>j�=�x�<lES<x�==��=��>0>J�
>��<�3k=��==�:�<e��=�^>�+�>+�=��>�
��������$��H9��s�>��>�檾胏>Y�h��߾���J��>ؗ=z�>��>� �=oo�>r��>�p�<^ę�s�潽x�=4#�=ηp>�=�"L=ݡ��6ee��	R�O�=A���)н�/�<;�=���>�α=N	^>�pJ?�?��,?�>x�a�V��^ʾW����-<��ɀ>4��>�
 >�H���������-eþ�ɤ��U�I	�=� $>�;�=ұ�=�Yj<� �uc"��h�=������=V;�>�->��d>���>�z�������=�c%��6޿:;���n���$־�j�����Ip��#ʾY
�>V >#��=���>���>��O>�%=����J�{Ѱ=�Ӕ=6�&����<ƈ>�M0��ŕ����������<7+M�90>�>�a'\�;���X%��h���˷�\�:��!K���l<�ѿ>̖�>�o=�l�>
<2?g��>3�#>R�V>�ӕ>����.)��v�~��b>�>B �>���>�m��(��=��|v+�G� �0�=ZP=�?;�"=��:�)���=k;@+�F�~=��۽�������%�p���-=�p(>�f��w����>j����?��2�޽v5,���9��>޸r�zF.<�-ؾ��4��@���鄽�Е>��>g��>P�>J��>V{4=�K4�Y3۽�B�=��+�E)ռ�=�<�G ���<���������H�=�c�>|U�=�
>$l	>x�=��H?L	?v��>����N��������*���4��(���z$=�u��`,>1�����^L6���n�ݾ[d��
���>T>Ǫ�=*|x�S<�<E����!>���=����닻��=�¡>aX�>�<>��k>�6>�?ϻ��^�:����i8t����g)��O�}a[�M�I�굛�O c��� �{�w�|_���k�<���=�>��E�2�Tz��zͽ͑־?���/e=p8���r�2˞�^���(*���K��P��;�}�	�ݽ1����ኾ���c�ž^���䭀�����><r>�}?oB�>��>��'?�*+?�R>�;�>&�r>+�>A�Y>�y�>x+?���>Z��>3Ν>�2�<���j)����b��2B=�Qg>R�;��{>�`�=S�5=|~)>�}�=`V>_���|=T|S={.��sZ���0=�I)>w��=Ŭ ?��=J�th�����_�޾,:U���>���-z���w[�=<�U-� �/�L�G>GT��O���U�>(��>ϲ ==�U��$�=���=�V ���=��d=��G>/�?S�{TM���O��0���	��l��5>`Z�=���>G�f>T�m?^%�>�>?�9�������|�؀�8��>dľ%-��I�=�֘��Z���#�X�q�	��Z�fXھ_�<�u�>�[�=j���
����=Ij�Y������-�:>O�{>�6e>�y>�ӂ>�Ɖ>�>��={$���c��ٿ�Y��7񾊳3�䱳�#�z��ϒ=�(C=�m���0(f����4=p�>OJ�>�=�e>�=B?=*��� ��=�h[=h�D����n���:���$�MO���@����P�f��Ż6J�Ls���%0�M�F�mڽ ��>K��=,�?~�?H�>��D?�x'?s��>�n>�s�>B�(?���=6�?��?Za5?�V�>���>�Y?!$����'h�an�<��)=��<���=�`�=��8<C��������`=@9��m
=R�ļ|D�=,м�Mw���G=Ʊ�=Ŭ ?��=J�th�����_�޾,:U���>���-z���w[�=<�U-� �/�L�G>GT��O���U�>(��>ϲ ==�U��$�=���=�V ���=��d=��G>/�?S�{TM���O��0���	��l��5>`Z�=���>G�f>T�m?^%�>�>?�9�������|�؀�8��>dľ%-��I�=�֘��Z���#�X�q�	��Z�fXھ_�<�u�>�[�=j���
����=Ij�Y������-�:>O�{>�6e>�y>�ӂ>�Ɖ>�>��={$���c��ٿ�Y��7񾊳3�䱳�#�z��ϒ=�(C=�m���0(f����4=p�>OJ�>�=�e>�=B?=*��� ��=�h[=h�D����n���:���$�MO���@����P�f��Ż6J�Ls���%0�M�F�mڽ ��>K��=,�?~�?H�>��D?�x'?s��>�n>�s�>B�(?���=6�?��?Za5?�V�>���>�Y?!$����'h�an�<��)=��<���=�`�=��8<C��������`=@9��m
=R�ļ|D�=,м�Mw���G=Ʊ�=_�?H�˾��%��Ӿ��kbҾjX����>���B�`��t��܍�����1l��ۛ>i7>J�>?i�=���>���=[ي��^���V���ѽ�>��=�C^>��M�<�׽]Lɽw�>�i=�ݮ=�S�;��-={y=��=���=��?\v?/w�>�Y���E��B۾������!C6�	��>�L>�_���i'�٨��������4b,�4�Ͼ���ɱ=�Fp>�/�7�>�<@;�L=� /=w�� �g>Ы_=$U=�嵽�3=�8��M!�==�'�jݦ�/��w��5���*����� >߷��������ſA�}ǼW	e���<�'q����=ЄE>+x>�p��r"�=�(>�þ�Fb�=�ɠ�mR��Yg�_{�
"x�b�Ծ���aJ����,>�#E���?�	��`�n�w��b�m�;�����?��?�m�>�D�>q?q6?���=�z�>�t�=O3�>j�\>�{?�j�>�B�>�U��^h>��!=E�h=>{����D�=�>č{��J>xh���û�f��;g�=cy>���=�rfa�4�E�&�л�x�=DT>���=Ŭ ?��=J�th�����_�޾,:U���>���-z���w[�=<�U-� �/�L�G>GT��O���U�>(��>ϲ ==�U��$�=���=�V ���=��d=��G>/�?S�{TM���O��0���	��l��5>`Z�=���>G�f>T�m?^%�>�>?�9�������|�؀�8��>dľ%-��I�=�֘��Z���#�X�q�	��Z�fXھ_�<�u�>�[�=j���
����=Ij�Y������-�:>O�{>�6e>�y>�ӂ>�Ɖ>�>��={$���c��ٿ�Y��7񾊳3�䱳�#�z��ϒ=�(C=�m���0(f����4=p�>OJ�>�=�e>�=B?=*��� ��=�h[=h�D����n���:���$�MO���@����P�f��Ż6J�Ls���%0�M�F�mڽ ��>K��=,�?~�?H�>��D?�x'?s��>�n>�s�>B�(?���=6�?��?Za5?�V�>���>�Y?!$����'h�an�<��)=��<���=�`�=��8<C��������`=@9��m
=R�ļ|D�=,м�Mw���G=Ʊ�=q�>�P�����K2�.�K�~/��	�����>G%쾩�=�^��D����Ⱦ|����[����v�7�?VH�>߂�>��>6����xļ/�(��Z���M������=�\���X=k�[�����E��h����t�,�Ծ:?O;�&�>��>~�*?�>$�>?����۾Vy
�ϔ�^Uo�'̕�W�>?qq�����1�NV����}<������XX>�
�|��=!��=�V�<�43>M��=zs�<К=]�>��=�8>9� <*��>"��>9��>�O�>|2x>�������տvԳ��e�P@z�:��>e�A>c��>:uZ<��>�)�>&�����z��=?;Iӽu�<t�0?]n�>>�򽱏|�x畾�$<\�I=����wrb�������ν&���G��<~�c�@Ro�H��=����.M�W���6�Ý%����=�>;��>��j>쁦�,?�N?��>Nֽ~~�>}�=�5�=��?H�?�A?�??��N?Z�>xؾ�
�4�t���}[>�o��>Ե�>�`�>O�=��=�8>�)�P9>	_U=\.>n��<���=u�\>h"n>y`>���>���i����6����E��|���<��\d>���Y��=5��.嫾JoȾFb4��#��_оg��;�C�>�\�>J��>U�>O!���É���T��㡽�:D��[�������`h�	��=��1�6���E�����߾�`n�/:ܽ�d">�<>/��>��>?���>�U??��<1˾���𓝾���=���~>[�@������M��f���!�+y-���sMW��9b�l29>B�|=�b6:2��=���=�^v=o.����>���=7j?>���>_�>y	�>4�>
��>��>3	����3q��?X�����|��ߗ���G�>���>X̏� ;�2>�p$=�b۽����W�>׭>Tl�>��>2Y=���<�����1��sd.>�<=֋���4��P�����I�n���A=A�����ֽ�VM�{�[��9����g�-lT�Uv��?	,=Js>ۨ�>��Ͻ�q^�9�[?ʜ?��X�D�>X��>�F~>�i>F�>Nn?_�)?<++?�%&?��>�`��s{��b��r���zA>M�s<��>���=�@>rp�=�w��2��=c���t�����=�,�=�@K>'��=�J�:)59>��>���>U�8~��^���������K���>㚾�@���,���ན��޼�"�e����w	��_/�>�(�=���>/��>�NA�v�P=>�ڽ��ýT̠<�ֳ;fa$>%�s��b��?�<�|:�	��z���?<�j�Y�Y>�Ǖ>E��>b�3?��>?6?#�ƾR���٬�?�n�[����ý{-�>�� �2����)�����\
�]o��&=ϣ�S�=`�]=��<U�5>�h>j�=Z
�����=�z��c>� ����P>�Z�>��>z�H>C*�<����%��=�+���X����6m����c��[4��M�/:��1�i���㽜<��;��>�0v>܈=\H��)3����=��==��=�G=;*����侦�=��ž�㽜�	�f�j�8�t�;K���]o�?h�|k��ݽ�2|�"�=i&��7����
�?[?v-Q?q�?�������>��?T�>�}ɽ��?5RJ?yZ�>��>��D?�ϼ�㽉7?��ؾ�Z�=�����:2>F�=��=[(W>�6t�֦ >�wX��+�=���=�#v��>7��="�>>��w>2�?T[>��5�����|E��c��損��m�>H�پ�C>D�@�����.�������Ծ�K���X�HyE> ��>�W�>vz�>!፾jB�b�y����=�X�������=Y���U����=��4�1kT������ݽ%�q��4>i�>zW�>k�?r�?gX?�:�����|��cT�*f��Y�����fu2�����ǩ�S����r+�=����g�D�8�����Q=*������<Y�x>�i��>�;|!<>
:�>Wë=�[�>vo�>ذ�>�J�>B9�>Ċ�>|�=�̫��a	��ƿ���k�Ҿ�����==�-=��?'�<W�ڻ��=P�>e����
�CW�>��><�t>bo�>�l>����j23�tM0�"��Ь�Dž1����㾻�=���h�=Qe��=�H����oڼ8��	[8�	��u��8�>,�>��=��2=�W?�
�>y�>6'�=u9?���(����K?�?ͨ?�?x�"?�P�=������A��C�{�R�ݹ�>�d�=ҭC>�z�>��>N�����Ji��=��Uj����-=���������>��i>�Q9>sg�>�0�������ǽ���]ڡ�ܠ��j��=�Մ�K�X>J��"���P�I��ȓ
�	�e���[i�>��i>�>%5�>�?��I孽1����7T6�ώ�@�a>Nq>n\>ӖS>Ⱥ����<��R�U*B>�gk��$I=�s�=x>U>�@�>P��>H�?�`��O�о��:����[�����=@gk��KY�wC��zؾ�������������*н[^���22=V�=�n>/��>�:>��>�<>�<ǽpŒ�M��=�:н���>�,>���=2��=JOz>$���	���9ο���)���u̾'@=�!,���>04a�ř����w��SS�����uՓ���=콎>̐�=">o_c=�-Ƽ�{�>�
O�E�+4�f���r�������Կ�����$=t䗾%MV���T�'����I���Ӿ�?Z��4�<PJ��K�v>1?�f�<�)���D?�)?/�?��>j��>Ds�����>?m%?�+?�L?<;?3Q?��P�����մ�&ۄ����>�ě�DW|>�>0�>�S�&����F<���B��;�:�����u�=�^<zt)>۱�=)\�=�|�>���<�O��(�4"2�HS�������\�>��پ�^	��B����Ҽ4E�d��� 	=u!��"��
��k��/I�>��>Ю��gT=d������<�4>q	D=�L>=��>PF�=��5�%F�=�5���U[=g	��K����`�-�e�J��=��>:�?�?�����ʱ�,���{y�V�����W�gx�=J�A�݅a>����l�Ǿ�������žu7辮l��_��>��=��K���6>)�2�d��;�	���S>�W=���<�y�=�Nb>O�a>&i�B*5>S�.>CW/>����׿�#������׾��=��r>�6�=�<�]丽)��$���Դ��v�{7F>���=7C#>�[/>��$>s��>��߾|�z�	�b=`%��F�������ؾ�l���྘���N�{��q��z:c��iF�� �*^k��{��E~������O>)��>x��>�ɫ>O
?wa>x�W>m��=t
?2�>�w=���=���>D�>Խ�=.ի>t*�>��>E�>?΃�d	V���=Z���[��>�\>�)�<�=�=��A=T����'@�-��=��ؽ3�<�~?=��>���=�%$�{�M>�|�>���<�O��(�4"2�HS�������\�>��پ�^	��B����Ҽ4E�d��� 	=u!��"��
��k��/I�>��>Ю��gT=d������<�4>q	D=�L>=��>PF�=��5�%F�=�5���U[=g	��K����`�-�e�J��=��>:�?�?�����ʱ�,���{y�V�����W�gx�=J�A�݅a>����l�Ǿ�������žu7辮l��_��>��=��K���6>)�2�d��;�	���S>�W=���<�y�=�Nb>O�a>&i�B*5>S�.>CW/>����׿�#������׾��=��r>�6�=�<�]丽)��$���Դ��v�{7F>���=7C#>�[/>��$>s��>��߾|�z�	�b=`%��F�������ؾ�l���྘���N�{��q��z:c��iF�� �*^k��{��E~������O>)��>x��>�ɫ>O
?wa>x�W>m��=t
?2�>�w=���=���>D�>Խ�=.ի>t*�>��>E�>?΃�d	V���=Z���[��>�\>�)�<�=�=��A=T����'@�-��=��ؽ3�<�~?=��>���=�%$�{�M>�?�۫>�x����ؾ�h��[ܾ��>+?-�7���y>�D�>�'��2=\<����ܾm��=Z]�=�=e=� �|E�>�.�=�;Žl@��*�ͽ��=�oO>|�>�7/=��4>���l/��,6������8��hp>�<�=��>�چ>r�L>��?�oS?6�%?��d������׾�I����<���^F<5�>4U��2x�P�����Ym��c�����O����>�eT>�H�=Ru>�+��Ǧ>��1�<ν|��W�>G�>?p9>��>3>U>X�	\>e��U"����_<���F�W�-��3=o�q��T����cg">�̮> ��;`��>��l���oK�=>�ýʻ�e]4>DE>�Պ�9�>��;h=bJ�e2��c���W��8�1��>�iy������QY�i��H,1��̲=+����}0�[�f�a���>��>�3->;X�>��-?
?�$>������	?ƌоUN��ғ>r�J�#��>7 �>�>:q�>*7=
L�>?�D��2�:���dt�;�Y�=���<� �=+����|�=b�='��=��:e�S���T=5>O�Yv�j�����<���=}	�>�#>U͡��ʓ���a�Մ�� �O=�?��C��(�ߎ�=�����\>��"����?��>{�$�h����&�K��>���>A��k�ռ�|���O�:9=U�+>�bz��f>ɽ�<����<���[k=={P=�1q���ܽI��M@�=��>?):`?��A?�@�G��{��*��mK=Z4v>��<��uݼ,`
>.p�=���F��p�;���=��n�`>M->��u=�-�>�	��A�m�
��~�λ�W#<$T5>���>�g���(o=�Q>���>>�=s�$=�)ݿJ������u{��/�=��=�%S�ܥ"��n1>$e�=#\f���,��gi���>�ʼ�4Ѽc\>�{�=�#(>�`=[̈́�fW���5���z��3%=/����o+���V����z��(���1N<�ւ="\*>�51����\�I��[>�����s�����I�.?��?�u�=q�q��g�>᪩�Lu�<�
?�e%��k�>&ކ;$J�?��=��>�@W��;��;"߼�N=���=e��=ç=@4Y�� �=����䰽����K	>w�[=��o�Z��%��=�M=�?�۫>�x����ؾ�h��[ܾ��>+?-�7���y>�D�>�'��2=\<����ܾm��=Z]�=�=e=� �|E�>�.�=�;Žl@��*�ͽ��=�oO>|�>�7/=��4>���l/��,6������8��hp>�<�=��>�چ>r�L>��?�oS?6�%?��d������׾�I����<���^F<5�>4U��2x�P�����Ym��c�����O����>�eT>�H�=Ru>�+��Ǧ>��1�<ν|��W�>G�>?p9>��>3>U>X�	\>e��U"����_<���F�W�-��3=o�q��T����cg">�̮> ��;`��>��l���oK�=>�ýʻ�e]4>DE>�Պ�9�>��;h=bJ�e2��c���W��8�1��>�iy������QY�i��H,1��̲=+����}0�[�f�a���>��>�3->;X�>��-?
?�$>������	?ƌоUN��ғ>r�J�#��>7 �>�>:q�>*7=
L�>?�D��2�:���dt�;�Y�=���<� �=+����|�=b�='��=��:e�S���T=5>O�Yv�j�����<���=ˈ>i׌�yR:��gǽ�3�!����v=��?��Ծcu=��߾�>��(`�'���!�$��޽���v�>��>7�B>�N=� >ؽH����m�;>>�x�l�S<�cP=�����&%���4��ie��,���	�Ľ꟧=���>��W?��$?��>�����*�i�H�0M���~��φ����&>)y�>@u�>d�=#���L?������9�ZȾI�(��&?>�!>M/�=�έ��ӽ�1��ȑ��6�>����Qͽ��>�r�=�j�> �?���>�͆>�{9��,ؾ~3�����!{���Q��6�:��%��EI�]gV�
��==��G2�O�B>so@>J��=.��<�.>�nl>^f�>{����e{�(�P�ݾ����a6н-���U�=��H���)<U��� bV<�հ��R��}�/�e\��?��_ż]6$;�Hz>�Lt>#�>ch�>�D?T]1?�[�>����� �>Et>��>e�>SO2�Ё�>�r'?��?9��>���>�]��2p���N�I�d�<G�Z>S�)>�9>w�ĽӘ
<��$=��E=60��}.��ʪ2�ؔ�4��<�_�d�>�>5ל>6'�>��;��CG�	�̾v�>h��>c��ޤe>K��Nd%�V���,��%��'Ѿk�ս���>�7�>I�>1_�=�n��E�'=J֏�p3��vq�<7ԻMԪ����0���x�<r�u�����_���@pC�6eE��KK>��D=+D�>a�6?�#�>M�?b�v�a|�XeK�&�O�>	Y��h�N��>�m?u@��O�=7���aW˾���h��*���N�/����>-�=�*O��k >՗&=ܷ��&��=��G>�]�=�>'-�=���>�ٺ>�� ?�I�>��=��c����������������I����s=��=�=!��GI�}�:��1��*�g�|��(>���==�=җ�=�<���=E��ͷ�,;ν�������sؾ�7׾�����6��R�=q*��Ҋ��Ye�n�u��*�Ls�������s^|���>V�>LW>��K?b:?��O>+�2>�4?&���6�>�Ɨ>��?�@?�'?c�,?"�?ݹ��)e��iH���.D��?�=�>��6>�>�ܔ>һ���o<�r���a�A8=2g-=/�y�,�����Բ�=q��=�l�>c��>I̓��J��}ａ�Z�Õ��������>D��Ƞ(?U@�l�A�P�A��A�YVD���������A�>~�>��>h��=�r��=��
��=[��$.>����K��Z�=�h�������e���/6�Z깽D�=�:���~�>�%B?���>?@?�M�m��;k�k����3�^��A>���>ɜ_>z�{=KY��S���I�W���P�������>�2H��
=<ҙ�=�������"��7b>�U=�,>ŗ>%gv>���>�p?,�>�/+>�`��Y�m��S����u��s�N��?�;��>C�=oU�����}#��Ǿކ-=���=�n!>��>��t>_��=�ԧ=�0�>�F����:�1�<b�#�PQ���ԝ��>������=�v���W����\���v�U��o�K��'z�(�-��K���=b��>�d�>�κ=ewQ?�h?o�>���=�'?c���#�>_��>��>S�?�. ?�� ?�?�[o��OW�����c�!��=�
L<e
>��J>�b>��<��=#��w$��^?6=+@<�.����A{Ḵ��=��=	�?>v�?����Ր�uF侍�H�c�Z�?��Z?� ��C�>��������Q������4�:e�`��o[h�-f�>aO�>�$�=x��~Gὡ�=MN >��<J�*>y�V���t���Ƽ�37��` �Q�=�1N������NQ�|�>�)&>u��>�!5?�[8?w��>��ھ��-�F�m�1�2���_�=&'>Iޠ>j(?��k=��D�N]���m�e����B)��4a�>�u����>�!>��ὒK�������>�f�=��=�đ=5��=�'?�X?�x�>���>�þ2����x���3t���*�p���E��.�=��c�7���u���ü�ҧ����[->���=I\Z=S��<��=6=���ٽ$�!9����{�8�Ҿ6��T�Z�4 N�Q!]>�2���(>�֎<:��R�����d���cm�1$i���=jU�>�w>V,�>~�L?���>���>
�ӽ��?ľ��r�>M#�>�樽l��>��?]?�&?7�C>"�D�ݔнe�+��@�=Qk�=�D�=��=��>���<�=Լ%�潛��;A���!���A��K���s��ؾ�Zq>f��=��>�L� �澬%����@�*VԾ�>B?=&þ��>�载��Ko(�k���#���۝�L[,�	��>�l�>\�>"�=�]��5=ܑ�O�ҽ<�F>���>â��U#=Bh��qD�?���8�q���<�Zz���隽�at>��>��>eT?��J?I?>o��l	�n:��L��ޠ�����S?+�>�">��>ɣ������296��5��qr�(ʙ��>�l >U�7>Y=�<2���{���(�(	>�8s=є4>�~�>N�>iܰ>���>�!=7Q�<Ta��@e�w�ǿ����G��w��%$>���>��+�����R�>><R��I��/�v�h׽���
�нA?�i�>��R>T�������̽;�����;��ć��$6�𤾧�@�3�J�S����1���5N��I��=�e�8.Q��%��齞�?��uv���\>��>ڇ�>y@�>�o9?0�>��>��@�٣�>Q���K���N�>"?q*?Ö/?�&P>�G>���#쪽[᳽�`���=�l5�G�>r}>�Q=jѽ}��=T[���[�n�e=.�=:5!�k�<_�^=��=!��<-� >�;?0sƼ|�7��"I������>�e>��b?��=�Q�>�t�>x��,�&>��'���D��:�>Y��>aT=?-S�>�y�=z��<�(H��o=^�0=͔�<�'&>�4^�ϝW��"�;�����˽
`U�5�����I=�D#>��H>Q >b�˽�*8>ƪM?~~T?[?�R�3���þ��2���u���m�l�=�>��s������H��&����@���'����>���=��^�P}>$c��;�W&�=��8=����=7�=�T>��%> {�=��j��eW�I�Խ��?E���"��I��,������>5ˢ��/����g����7��=�g���y^=�L�=��>E�[>[�=eQb=������=�:< �����%��X�=^�3�����< ���ս�pC�g#�<e�3��'�N����؟��,��N���R�0V�S��$>�>���=3(̻''�>�s�>\v�>|��>��>T�f>e���>=�G|>/�=,��>`��>也>Z��>"�>a�����2$��]�>���=�����}>�= �����b>2Fn��2�=Dl]��W>�Bi����;j��<�n=��X>q��>;�?h����վJ&:��+!���>���>V�?�Ɠ��>�>>�>�����ؽ5+E�*���?��>�{?�??��>�gP>9�i>M�9����K�<���= P;>:'�&�>���/>��w<7����ڵ=��=��+>Z�=��=e���#ސ=+�I?a� ?n�>��C��yþ$7J�!:G���6��_ھ_�H�}DL�e����>d5p�A���,��-��������HS<��=Ɔ>��=ZC>SII�ϾP�)�>��r=�� <p����c>�h!>���<�	P=1���n޼$�۽�P<�$¿m*����<������:���˾�``��W���?�#��rc����?>s�>�x�=�|��U���̾�盾����_x�K�E�˽��wU���Z�n[�|�f�����S־]��W P��7��/���l����I��|1�R���p������>�>�>u,�>r��>��7?*��>�>�>�a>� �>y,�=g��<��>[��>��>q,?��>-�:>�����ɐ��_��I��d�=�氼�����/>[��=X�=v� >$�=�=�<��=U\�=��=�X5=蓝=s��=`� >l>��>�g����쾞aO����ע=F�>�A6?.�Խ&��=���=t� �����E��J���`?>��>��7?���>q�w>�c>Z�/�� =���<x�$=��A>�(�������v@�������׽@:�<�����8�=�:>&[�>��;�'�=I�&?V?��!?�{྄���{������ >�I =ݖ��R��=}�=�<\)������b�@��eJ�>��=��=>!Y��=Y˽�7=�kX��0���=ts�=�~�=��l=h�}>lA�>�Z�>��>h�=m��T�o�ֿ��Wʿ����	%��=��ͱ>)u$>����V��-Z!��6����ؾ$ྎ���B`<�a����ʼ �<)��<A��$C���Ǚ� �=}�f�~޷��⼄�����y��#
���)�eaO�Lf9��FȾ�Y*����R��O�x�zR?��Q�>�@?㬥<ø�>��D?��>y#�>]O1>ق�>�?^>.X ?4?L� ?��?T�?�7>��>t�����+A��A�
��X�=�o�=��,>��>��=�w�=�O<����=�ʮ�~A@�V�;���S"�����=�X(>��f>�21?cr��i�5��� �r�1��YC�B>�1?!�U� ?MM�>�ܼ��B$��'�"s���=6��>��?���>��>^ӏ=�S����y����=<�=ņ=��=b��>'Ӈ<*��='a>�y����=Nތ=�"v>_�>L��>�ʓ=�=x�@?h�K?�[P?c�.�L��ٹ˾�H�w��=�ˤ<�A��q�<ac��n��zھT���#���!���rBj;a��>�2M=�g�=l4�=�Z˽���=�	��;j�C�9>��g�ຉ�]=�?���AW�����C������i�hʿ�H���˟�����$�>��6��Z��N����=p{Ҿ�86��X=G",>wg.?���>��_>A>��[jm>2���1�#���<����	�r��82�N�m�%�ѽ�̈�����tg������׫�уv���P�@$��uz����9?3���>�A�>��3>2>Ȩ?�?o��>$b=@��>�pm��=4�>�ǻ:�>W�>_a>H�'>I*I=�'������.�}�wv>���<�z�3!>���� 	7>��	>-����u>���Q>��l>,X:>3^=�n�:t��=?A�=�Q%?A�ƽ9���5C���6���=S�>��N?��>*Ql>��>wZ��O�I�O�pX�((>�1�>fn0?��>�jB>�&Խe偾�l��p�5=�>��=�5�=���E�o��X*=b��=-�ؽh��=Y�2>�JR>]��>V�1<��>i�8?��\?�8?�4}>}Q˾�-C��2��\��t=��>�(3�=�\9���\��q��"o�}��L�����[*��rJ>���=�u¼�����	�r�LoT��ڿ=�����Y��=1r.>�>�>=~�̼�
������#,��J̿x豿��ؾ��ɾmF��+�=d}g>=.���Gw�Y��U�ѽ %�>���=@?�8�>^�>��_<��J���>�	=HN>�b�=u�;�j`����%������s�p�s�B���)��A�O�ʽ~��fe�>9�J㝾Q��
HO�f��>&��>�ێ=�v�>c13?>�l>�N���>>Ker��"I��7=�b>�(�>�R�>�>Y��>�<܈��`5��Ʌ���=J�<c��=��=�#}�j꽼�f�=��=k�=��ɽ�\=;�N�=@?�=%CǺ�7>��=J�>g�/?(�0��OU��]�P����
>r��=�n�>��=��C�b�\��q���%!�ZG��᧾T�N=Ձ^>��$?r!�>�EE>�7!>�G�'�ٽBt=��T>Q�5>�p���a��w���8�`$B��ٽ.��r৽��>��>9��=%#�<�>�(?8aB?E~�>����,Q�O=�T<�辒�ɽn5G��6����<���~��^y,���F���C��z��7�>�&�>G�ӽb����:=����cK#>��6>&DI;]�2>[z�=�}b>5�>��g>1�!=������0i���տ����iUҾ��"��!��+�/�vi?=�M�L1����>�ػ��r�}Rv���C>�W�>{�8>��=�-{=Q���WIQ��
�͔>�6r�)�m����h��k�/�)� ��
���f����߼a�߽hӐ��M�V:	���&�R�6��0!�ͮ�>��>[�<>~��>��+?���>��>$��>a�?�HE��b�>eJ�>�'?`�?�?���>k�?��C>�A==�&��[վ��!> Q>*1=)�<���>����6��
j={
= W�=!��8>V#e��l��>�<T��=���=G��>�י�@O@��P%��X羮����`�P-?�q>�W��e>dY@�����i�8�o��T�>�>�-�>Xpp>�b�>N�Q>����iX.��)�"�o>���=�A=I��=A��=�z>�����H��0�+En���E=�O<>�j�>���=��=
P?��5?�?Y�<]�վ�LپI �p��?�>:B'��yٽǓ�=}늾9@;��~]�͍����*���!�>����H�=��j>�C�p��gP>�=�l�L&�=2x>Χa>�`>�i{>~hv>da=,�	��\E�i'ȿu)��˼���?K�ĸ ��">��	=��㾼c��'���}2���ߔ����=B >�Jٻښ��2���K�������W��C���+>Ob��O�a��:���=[8=�VX�`߽��c,�Mh6�����u�}�Aױ�~�߾�^��f�=����>��>Y)�=��J>oi!?���>B�>R��=�*�>Zj7>;_>0��>7�>�A�>^?���>.v ?!�V>ڕ�=��������j>4؜>���=��7>���>ޥ����Ͻwa�<k+�;C:T>"��=��\>G*`��H��b�=��պ�;N>?M$?i!N������?V̾��A>]ٽ�yR?$t�=��%���
>�$>����w-b�� ���`��@�>��"?��>��>}�y=�&��DG��*m�?�v>��=��>�mV>��#>�oֽr-���׹�:�޽Xa��^�M>�Ð>˰�>p�==���=�� ?��\?_D+?�ZĽރ��*���%�c��5����>	���ޘ=␄��Or�3���@�R�=�������A=n��>^�/=���=W;�=<gN���
�_f6>��;f� =?��=�9`>�vS>/>�A>N%s���/��
2���=hӿ����+����]�1>�k�=R�>E���\���T2>�>��G9��r�н�@�>�n>
F�>�V>�ۣ���;%I���ǁ�� �m�ͽkM�CC����r�ѽ�uy�WK�����i�����;�S��G�M���>����t3���>���>�=��=ꮾ>DW�>�2�>��I>/�? �=>�/���ӗ>���>��>���>�"�>xI�>m��>EK��5i	��<��at>N\>���=aU>gh�>�p��9��f9��bM=�>�����=dY>�C����Q)�M{>�5?=Q���{7����\���Ľ��=��3?�`�<�[��;y>y �; (�8�
���>��J>C�>��?`��>��/>>N)=ᦾo��9��=�g�>��>]@�=�a�8�񺌨�����eQ���E��n����=�b>g�x>ꗊ=�>=k.?��i?f>�>޿L��F��^�ྃ_������1�䛒�RE�A;$>J�k��At�X^���E�&"@�їݾ�T0=V�>�i"=�&=LD'>���-��ػ>iN>�g��U�H>J�x=��>ĭ:> �<>�3=�{+���E�)!��Cb��1���\=Q"����7�={�>���O��ǟ�>���c*J<��̽���>H<>]>�ڨ>��>H�=�X�8���y�<@����~�\��"��gؽ����%���7�^� ����Ce�����&�/�p�V���c��Z,�V��>x�>O����oK>6�?�� ?�ë=��>��>�ү���=-{>?�I�>%��>j}�>�5�>�Q>�3��煗>[_�>�?��Z�<̇>�-O�X�<�ݶ=�x$=�ĳ=�<�7>i�>���M_o<b�����+>��?s�F�y�F��t��L�b|M��}"�>M?�����H���'>��)��j�������ﳽq+�~���0�>7��	�>o��=x{�m���p�o=��d>�q���8>K�P>�J;=*]��W�=U���Đ���^���;>��>�t�>���>�e>Mq-?&�C?�?Y �=7�;���qJ����$�d���!�1�|���+����=��'-��y��� �+q��bO��7W>�����}>%4*>�;�EW<��	>���=V�Q=�	>�ƚ= ��>��>�ʬ>ݠX>�$=�� ��E��/�ʿW��b!ٽ┥�r�>�
.5���>F�]�%ў=���h�]_��6N=p>�Q>��g< �:>���<�\>S���8��Y>����HL޾�/���u�f��q�Ƚ��i�nv/��>��@*�%�ϽI1��"wþ�ƫ�B�����>�>"�e=�*>�R?>>��U>��>PO2?�ǆ>6��=�#?��?o?k�	?
�5?� ,?&��>��8>�\�f�VB?>?V;>3�=�,e>�c�>蘑�N�Ѽ���=���:��=g >�R�-D��>I��:=�D>��?��Ǿ�/ ��S.޾m�N=��>4��>�1�����>�Rb�x�u�sP�]0پP3q�
-@>�9>#p�>�?Y�h>Y�.><���Ǝ��	M>�JK>��Y>*yj=v������*`��<�8>LZ)�g>;O�=��A�Dᵼ��`��0�����>	?�?1���4�Q����׾Ǿ i����8>���=S}������龲j
�#���F�����M=I�b>��>�&=�N=����鱢=g⼋�=hhN���=��H=	�>[�F=g��;H�C���a�$�ֻ�ד>�=п����gŽ��Ͼ4"��Z�.�B�)�=��烸��[=?�@��<XP=p�5>~�_>�/s=�ս�\+<�5��|J�k��x�M>VS2�"����S��l��l���O��-����(U��^�=��۽��4��kt���o�ߐ�v��>��?�b	>�˝>q�S?���>��A>��%>�.�>�B���(�=	��=l�>��>���>L��=%�p>L3=��]�f�*��]��H�=.�>ׅj<oS4<x�`=#�<��>�.�>�(>>�=���&�-5���#��K�-=N��>:>3�><�>k���ľZ!&���6���-���EMH=���=�>"q�+��,\�+�ξ��}�S�>~L8>�C{>S��>G��> �>�k��=.�e�>��[>�_�=!q�=�Jӽ SX�������Y��欂��ˤ=�ڒ<Zլ�����/�3��=�V9?ъ
?�$?�n��VOɾql
�AȾ�c׾�v�<8�F>�<�n�����N�徤X��a��4���xνC(O�;D> �=�ۛ=��<�>��k!���(>�N�=F"�.B�=�j>�a�>)�>I{<߽�P�2p��K�=J����V�
�.����	>�`���3��v�I�<5�����9JvT<�匼�>�n�>ıF=�!�<�*���#����}lƾY���2��<�������nZ�K.���-��!L��-�<<U��1ߊ�4|��5�𽞸ǽ3;��%걾�Ӳ���n�:9t>�^�>Ϧ�>�>��!?�	�>S�>�|G>'o>Y�'����>�+�>\ ?��>��H>��7�|J=�ф=�Uk��R�BX�>#�=N�I=g�#=�?�=�����=�M>�nM>4L;=��$�~#=�75�x�=�5t>��=>��=�?�Z9����@�(������x�!���o�>��=9���Wɾǣ�f↾eྒྷ�_� ��>Lq�>#�h>b��>DO4>�y�>�����P��u>��Z>���=���=���T�:g���bq=�_���{����#*U=w>�(>#�g�T��ޖ>?��"?�h?�D��[:T�|��c6.�а���c�>+U>|�>u�(>��N�������?I3�4�=�nm��m3>����3m=&�:DW��3��t�=oR>8ͬ>x	����<��=�	>@�>�=8�zjý�tf�����N�=�}ʿM������s�d~��W���a��б)�� ��#7:ck������2�;�!>��,=��d<��=x$ >���;���&�پ��L>TxT�I@׾����u����C�R���[�<"�[�4��W�Ž�=�/�<Ҕ�<�V�?t���%9��>n�>gϬ<�D?��H?�e2?,?r�>W.�>��)���>�� ?��A>u^�>t,�> �����>�9,>�2r��8D��,ѽ��>N'>��J=���S�=�yO����;g<�<�ik>�;�F�=�	�=sg�<�`U����<]_�=�a:>p��>(�������}���Ԛ=�"c>���;W�f��;> �����G=�Ͻ=�!���۾���< ->^�>���>4�|>6�6>X~�����)�?>r��=޲<U��=���q���[����ר���_��}��X>��V=�!�)%���=ԭ�=��?��>6R7?c����ƾ����a���ﺾڗ�<(ˈ=R��~s�\�ٽ�0�t�����������ۿ�oʽ:�=`9W>��.>�+�� � =[�>���=N�<DY$=���>b.�>�>!>+�D>�D�n�� K�	�7�Ez�T�Կ�W����!������)c�3<���J��Tް��Q)�䁒<�����>�A>0�+> �3>�[>���
D��ܬ���ۨ>;y�Muվ:ߜ��Iվ b����z��ʃ�:�<�p>�����&���h=5�
�OB�cb����=�?m;�>7b�><&2?m&V>�H>kA�>p	�>�Fd�R��>�t�=&��=�A�>.��>e;	=�������)h���g�P�N��7�=y>����G㜼K~=*腽�Ź=�o=�&>�.�� �ȼAԷ=�`�9Ud�=l�=d!>W�����>"Ӿ���ƍ������Y=
�>���=���=���>��������[��v����f�eL�=��>��1>�!�>K5�>/��=�a���bA����=��=�e�=��=~�=�j0�
�ҽ���<�E<>�T��2<d}��VP��,�ֽjiq=��ԽLL?��?�&?����S���S�ξi�#�	��=��C=P�|�)h�g���hž`z��fjھT�)��ʊ�;�>?�>ģE=Rs�=p�<���;Y����"�>��=�>�2�=�����=��>� ��8�,�6������տk��ې
�-Y۾�;�K���𮾏$��-0���K�\U{����埽'j4>o�4>+>��׻���;�tٽ~��b���(>�񼀱˾��о���L|K�hG½�r�=K믾����B�<���)ٽ�������:�t��-��>]k?e�B>!�>��3?�V�>C�J>j�>�A�>�[d� �>[��>t��>1��>���>��=y�½�	>!�����f����k�=-<>� <>�=f����a=y�=W(i=迃>�Ņ��O<�Y	�=4�#�ϑ==�:>��5>���=G��>�E7���:���;��
j���=n�>���>���ZY���%>'�&>���:{����������A��0z?���>�!�>.cc>(:��:��M��'>rim=}�d�q=Q���нyx>z��=���=��<����c�	��ͽ!��=�����j/� Z�>@�5?E�%?���j��?�w�)�d���7·��Dv�����u侫���p�&�ԾK(J����FX��PۻA�> ��=
�%15>��ʽx4=7��=`��=z6>X�='<�(���$>�q��u=U-=��5����=̤ҿ�
�� $	��I��r�n��;�oҽ2H�/푾phd����xJ���.=��>Z�>�o�>#a.>��=A���>پtp��wz<U��=	،�����hj�����о"����ļ-&�R+w���%�!�N�q���X��~z����>�>_�E>=!�<�<?�ܧ>r��>-��>��-?�?��~>�Ƥ=7��>A#?�/?�0?��<?s�=s`-��C�H�����(=�?�=��6=">L��=����->��<��꽏��N��=Pt,�M>,X'>��.>�� > %>)�?9&�=�p1��GD�/�U��<{-?+�?#(�=ѿ7�9�=�$�>g�����=��
=���}'�m;?�?y��>��=#»�\5��]��H��=�ԍ>�<�=/�7>3E�&�%���	>�w(����<�D=�K��4 3�of>�>�C�=�X$?=�K?z3?A�E="���D�o�+�bʁ��5ɽ�o併�M���=]��c%�%��8rԾ��&�L箾dT�ٺ�>��q>3�>(�9>��������d>�/��$7�FS>������=�K=GI=�m>}��=6�C��.[���ÿ1/��+ƃ�������4>S̏����,\>��ξ����&���Ԭ�LJ�P��=�>(��=1�@����d��\o�L�M�w<��T�D�^���I��
h�T=�XF��yY�`�0�������<�)(�A�཭H��[b�WK�4���[��>�]�>���=��>�0?�85?Bڢ>���`�?��L>pV�>�Ԓ>�� >r��>�?5$?�p3?Dqk�u��R�=�o�����=?�<�&ʼc>>���;8�J�Q�>�1>n"%>�4�=���<��t���)<~[�=�U�>>/>�Z�G��>�E7���:���;��
j���=n�>���>���ZY���%>'�&>���:{����������A��0z?���>�!�>.cc>(:��:��M��'>rim=}�d�q=Q���нyx>z��=���=��<����c�	��ͽ!��=�����j/� Z�>@�5?E�%?���j��?�w�)�d���7·��Dv�����u侫���p�&�ԾK(J����FX��PۻA�> ��=
�%15>��ʽx4=7��=`��=z6>X�='<�(���$>�q��u=U-=��5����=̤ҿ�
�� $	��I��r�n��;�oҽ2H�/푾phd����xJ���.=��>Z�>�o�>#a.>��=A���>پtp��wz<U��=	،�����hj�����о"����ļ-&�R+w���%�!�N�q���X��~z����>�>_�E>=!�<�<?�ܧ>r��>-��>��-?�?��~>�Ƥ=7��>A#?�/?�0?��<?s�=s`-��C�H�����(=�?�=��6=">L��=����->��<��꽏��N��=Pt,�M>,X'>��.>�� > %>)�?9&�=�p1��GD�/�U��<{-?+�?#(�=ѿ7�9�=�$�>g�����=��
=���}'�m;?�?y��>��=#»�\5��]��H��=�ԍ>�<�=/�7>3E�&�%���	>�w(����<�D=�K��4 3�of>�>�C�=�X$?=�K?z3?A�E="���D�o�+�bʁ��5ɽ�o併�M���=]��c%�%��8rԾ��&�L箾dT�ٺ�>��q>3�>(�9>��������d>�/��$7�FS>������=�K=GI=�m>}��=6�C��.[���ÿ1/��+ƃ�������4>S̏����,\>��ξ����&���Ԭ�LJ�P��=�>(��=1�@����d��\o�L�M�w<��T�D�^���I��
h�T=�XF��yY�`�0�������<�)(�A�཭H��[b�WK�4���[��>�]�>���=��>�0?�85?Bڢ>���`�?��L>pV�>�Ԓ>�� >r��>�?5$?�p3?Dqk�u��R�=�o�����=?�<�&ʼc>>���;8�J�Q�>�1>n"%>�4�=���<��t���)<~[�=�U�>>/>�Z�భ>7x��y����$�P�C��ry��,>Cۥ>`R�1�W>ޥ�=+�u�`����C��*�z������ކv>�u�>�o>���=��R� ����E�=�y>�U=� =�����d�`�=M �=��3���{�R7��[�=7�j>�+�=N%0?W�(?��?��f>NAþ� "�>����!������3����.�6�H���#��¾�%�����FQ�����Sv��h:>�>���=�+�=���K��m'@=��k>�$�>K]A>�%�h�y>J�>V��>Qo�<e�O�h$�������� *������敾Y�>a��;�c<���=huž6`վ�f�>܅�>��j>T��>��=�3�=�%=���n�(��E�����&q����'�g�Ci���v�zy�V#���\��m��=��t��V�"�R�X�����O4�>�>�N�>�e?��<?�-�>�>,�O�bd�>�,��8�j>q��>�s�>^�?+?;?�$?��[�݁��✼����w=�I
>.�}=���>�gZ>�Dk�m����#<�庼�0=���U->��B=7 ����=,�>D3�<�u�>E~ɾ��v�ƾ_���2��W�=[��=q�Ǿ҃�>��Y��1�YŤ��ʘ=Gܻ�k>�Mu>��w>���>.˭>�i���+�����{\=��4>�#�=��<z9b=8���/�=�E�=_)>�0�=z�->7�<:������ރ��a>՝?%�>2�m?�x��UbM��8�����3�5� *$��V>���<T����xt�����������˾��پ=����ξ���>S�`>�}�=z<�LP����|�==ס=�վc�=*�b=��<S�=D��<5��=棎=�	��Sў=I���GϞ���D�^��{���w�#�����y��Ns��_ż����O��D23���#��à�/�B��p<W���{�>�/>S��<;t>la����t��n_�H�����Et��;h�=��ƾa'8�K E�����悽;�'��P��I0�#4���=��?��t>/�=��?dѹ>5Y�<�=J�?�C����>�w�=�L>T*_���>����ҕͽ�Ŭ�L����p��������n>��T=)=�ݼ+�@=�A�����<R��>,+ ��7�4�%�9����i��+����=�}~>qb�=�x�>�ھ�¯�få�#����
/�J^<<�~>����O�^>�����l�� ��=+��>� ��$EV���Q=��>��?R*�>Q�];(�����F� >���=s�I=�ٽ���=���=w�e=���=��(>O��=��f=�N=ElY�������S4D>�m"?8�>F?ͼ2:�^���=��I۾#��������>\�=�?�(�l]���܄��`+�A����A.�"s�>R >Y�=�`�=G-��%6�,]k>J�+>��`���U>D���=�Ó=�v>�O�=�=�=�k�3�н@P�%ن������&��X�!�*�*�=|�>���<S�>�H�W���V�۽���;�z
=��=l����4珽��/�+�v����ۚ�;��I�꾾m�ސ���������JV���_��LὄO<�B�Ž�ɽ���1�����=�?5`>j��>p�<?o��>�o�=<L>c(?mzz�JZ�>'>���d��P�>���=%��=��p�����:%߽�����~~>�\#>�սڡ�=�!>�z=.��2
<��=^EƼ#��ⶽy ½���If�<sdo>�9�=�u�>E~ɾ��v�ƾ_���2��W�=[��=q�Ǿ҃�>��Y��1�YŤ��ʘ=Gܻ�k>�Mu>��w>���>.˭>�i���+�����{\=��4>�#�=��<z9b=8���/�=�E�=_)>�0�=z�->7�<:������ރ��a>՝?%�>2�m?�x��UbM��8�����3�5� *$��V>���<T����xt�����������˾��پ=����ξ���>S�`>�}�=z<�LP����|�==ס=�վc�=*�b=��<S�=D��<5��=棎=�	��Sў=I���GϞ���D�^��{���w�#�����y��Ns��_ż����O��D23���#��à�/�B��p<W���{�>�/>S��<;t>la����t��n_�H�����Et��;h�=��ƾa'8�K E�����悽;�'��P��I0�#4���=��?��t>/�=��?dѹ>5Y�<�=J�?�C����>�w�=�L>T*_���>����ҕͽ�Ŭ�L����p��������n>��T=)=�ݼ+�@=�A�����<R��>,+ ��7�4�%�9����i��+����=�}~>qb�=+�>sЭ�q����7�D��,��Ctx>��>G����>��Ľ~
����<"1�=��Ľr/�=�8�=�J�>?O�>�]�>�x�������&�Kd$>�>6Mq>߂�9H���s��Vm���_=�h>�݆>���=���Ք4�9r#��|=�M>�"?���>��C?���:��%���S��ҽ吾�� >8�=����=�E.��ڭ�dt�����jl��=��v��>z�=1L>��=�t޽��.����=��ּ5���>�f>��Q>,��=@d>�	>!/o>,��>G���V�����ۙ�#&">����μ�@�=Ϧὐ
ƽû��?�<�x�����.N-��	=Q�ܼ�˓<�ֽ��r;�9��e�Y����=���>�0��ds��]�����;��,�̾�C>(��?@E�W�~�����+s��rY�����Sl��2)8>�3>��?�}a>1����?�%�>=�Z�d�>-M#?����6�*>�G>���=�U���C>��<Л=�gڼ�����,��n'��E
>_>�����=��<�'=j��>�Y>>�>����-s��ϛG�rH���(���=J:>�U�#)�>�{���zȾ��V�L����>._b��������>�;��*��7�QΠ<吂�g��=<|���->Y��>Y!�>/]�!˾<'q�*�6>��&>�b�=��F�s7�;��/>����
>�r�>�L�>�=�^��t����IA�6{ûk�U>{�!?&�?�\U?T����v�F�h�ᇳ�g�-�e������Z8<�R��q=�=�޾�ݹ��y��z���|5�����j��>t}`>��H>3�M>�tc��]�W=D=�+��Uw��2�Z>����u":=�۽=pj>��=��]>C�=�������ק���k���?Mܾ�o<�}��('>�w}�II½a�k<���P�k���S>�5�>�J�=qt��?�n=d)�=�O=V�
>U�)>�zռR]��暾C�ȾMr���<;�8�/�B����D�9�������TN�Hн�y������%��d>�?�=1���>�+?�<�><��=-??�����=��:>��S>���H�>���;#?9>���=U���� ����/�,>F�^��H��G�d>�;>F>ix=X��=eu�9�D�\�f�rLf�^^0={�>ӗ>>_��>�X!�,�!�۾D��G-�F$C����>�>�>0�@<vM���!�Df��Z�н�W�=�{�>��[=�d>*�>ֶ�>���>�_�=DgҾL���?�;h��>$>*8N�4m�>��~"V�����H��a��	Q�'>���%>�I>�_�=K�-? �%?S�<?(^����վ�J��P����J�끺<Η>�>���=����u�����: ��W���e��V��/>�:���p�=c濽��ｗ�J>�K>�v^���#>�c>�q->�y%>8Z>.R1;���LG�W��8C˿uw��6J��!��I�V=ס�/���D��!<�^��<M�;M�ٽ j�=��">E��>�s=y$==���I��o5��u=��=>�$���f��V���䭾�A\�� �����*�nr��i�'z���^��k0"�v�,1�e;>�?��>�}>9!?��>)�N��X��+>�����6���=<�"����=�6��I�>Y�>��=�!�	3�˯���F�>�^>Q�c=�z�=��=�T��s><��>_}>�2�>�L_��a������L=6%�>� >k~>�e?lX���#�`[d��£��4����>g�>m[,�7d�]Q�[�ؾdjž�8�<\��>�T��l%=��N>ː>=��>�(>��b�g��=�1�:�Hv>Wxs>��M=�T���=a�i�����L�R�f=��?=2y>�Y+=9�=O�_>�A9>�5?��H?+�?7���C^�#��vxϾ�X���"=�m,>�`=��|"��^��k,�e���ž1־��O<��\>�Z=��ƽM!�=���oE���gb>0�=4���?N>[ώ>�<�3|<�X�=iR��$۳�*���*��\޿�F���*��d�Ѿ9�>޶U>$-$=j<���Tj�٣k���Ѽض½,B>\B7>��>��>�^$>#�>���>O��
 M���:�S�����o>�B���UjZ�-6˾3D��0����*�|���s*ֽ8���}P��bW�V;g�,P�g�>?o�>�D�>��>��x=u��=]>%�>_ۢ>�Z>E0�>���>+�:>+�<>C]�>�ù>�]=�K�EjɽkuW���>9 �= T�=xD>W��=�۽�tv>c>��=q������=C��9D�;��� =�)�=��=��=X��>��S�xY���}����X;;֤�>��`>d����w>y�(��Ͼ�7�
>s�!?P�?�Ȣ>G�>`��>��=gK*>5��iQ=2��=�i>��R�q�9�*���0 > ɗ��I�����]�o=�;��"���[�f�����<_��	�?��?Nx?t�	�w��f���'�<V��7/�bw9=�5����0>�g���+����6���d��2�Ҽ�A>/9>���=�y��I��a��F���ԇ>晆>����5ρ=���>`R7>Nc4>i/>���=z})<�m�*M������TI�B��+�����>/M>����R'��{链�N�=\��W���$�pg�;R�=ƽ�����D(*�3r>�-�W�*>��Q�Ӿ��¾l�h���=���-�m�+惾�#�z���}[���79���'���<��<�+�L1�>���>���>sA�>�d�>�k�>n��<�tP>�g?�}���� ?�
"?�(�>Ay�>63�<��4>$MN>]��=fv�\ӽ;���O|=6�:=�`>�p;>�"�=��#�&�`7=:� >��U�����GO�*Ӵ�H:,���">S�=.w>�c>�G�3 ��M���4�� ���I> F�>�?��(�E>�M�+�@[ܾ0V�=��?��N>o�f=zR�>MB%>���>�>�b���Iݻ?p�=��+>@�l>k���W��`H�:Mz_���c �;��z=W�"�>q>�����x<ꎳ=�{�=�+?�?S&?bN��'�p���N	�<,ɾ �>�KF��R���YF�����U�B�����|�������?ď<
��=sO�=B��;P�=v\6�����>�3�>��뺰�>>���>eU�=��=�b&>Mp�=�5-�z��C|��ڿ􏿆S��۾�S���7=�����6{��{�?=< I� <s������r�=t��=z���!��8^�L�s�������>+���| �2��4��B�9��̾^��<��˾S��7-������'�������@L{��w��;Q�A@�>ӷ	?��!=�҆>��3?o�>`ܧ>�>�(?쩏��??�1'?��>��V>����7a>���>!`>�>>�i𽾈�RA�=�>,>�=��=O�=����"��橼<.>�[��+"<��<�=�Y/�(�=ο�=L�1>_�?�ξ�ľ"�2�?���_YS>���<�Z�>����v��C���E������>��>���>�U�>+5�>M)>���>\�
>�{4���T����=��y>��j=�H2���=B�>�`k�K�,:�=�=o����&=�ȼE)I;��>�W�=��(?��:?�� ?��,>(0����v���̾_�x��>�i><�>�A���'��}8�<��N�"�R`���à=���=�k���댽��K=�� �Do��ym�>��]>6׼��%>��>z�>6�;>�Ry>�b�;|<콿��)_��W��#_�����1�=W0���T�*\3>�Q���w�b�<\e�<�/�=��=lx�p�ξ���m̍������=>���0G�s��;���JS,��抾U�K�<����9�M���۾�����)vs�&'�������G�i�vcݽ�y>�?U�=�Ƥ=:m?�T�>����Ctb>��>&p�>��3>�Ux>w�j>v��=?�F>�Ý>l��>㉑>�9��c㽆1ݽ�Z�>��>:bC�:�b=`<�<��s�M"T�j�9�koy<�R�>���{ɏ�A�R�=<[6�>Щ>�w>^�>pH�\aa��-������q>�G ?2b>goʾp�?������-�r�#��2��<R��"?E@'?u�?M�=&��>�is>�f��5򆾩W=�0p� �;�=���<��!��������m"��h��~��T�>���=�/F>�+O�Uig>>�4?-?~��>@ �u��*SF�/�ξ\|Q��k ���>�S�>&þ\<�>5�x�k�%��W&�^��b����={�6>���I�">�_�������ŽW(�=�1�=7%��l�3>�4D>��>9=�>��,>/�ǻ��= ����9<��������h����x���-/�F5�]��?�\��=b`��5��}��>.Z1�]�4���'<�v��8�������T��n����!��E/�䅾�ւ�$�׽≄�eнUd>�ͽViɾ�@9�ѩӾ�����m��P���SR��g?��w�>���>��>=�=�4!?
��>V�u>��>�@?������$�m	�>_"}>ߦ�>�,�>�ٳ�d��=fdK>��&>d�4��3G��&�> qG>�ڋ>a�4>��=�?����b�z>��M�9Z=N罽r���E�=/�˽� j�$�	C;]	?���`�IY �E�7����>��.?�>Wq2�T"?'4�		�~����(�ڗ����?%�,?��(?<�=��>�y�=��S��:/�n���H����p=��=�\5�z6[�9J��ͼ-���6���\i�=I>�sO>�iF>�r�=�8]>[�#?x�?��#?�u��/_Ѿ�D�l߾4pg>���=I��>J�>Δ?>t�Y>���Z���0�ii4�[��� ���>>Eǻ�Z">���	�սb�p>[e�=q%�<9	�=Q�S=s�1>�J>G�=���=�9=�ጽk���z+���R���m(�}��m!c=QQ�����Ib���;�Xy���5��������
�@���9�m�g�[�f��Qƽ�S_>o���_ͽ��	d���@��Vx�R���7j�q�Q�������:��@��>Y:��Zh�\�V�E�a��厾�Y	��uf>&��>2�>�E>��<??��=2��<Y	�>��?�)�W�k�w��>z�R>�?U�?[�&>�>HM�=�yC��H��wx���>���;�Ҋ>�#�>[W>�x�o٣<��=��k�d=."�o
P��2��Pz1��� ���f<��.�d3�>�X��S&�`���tM���%>�O?��>�%'�/��>>��>��/��)!>�Õ�n��<
{l����HT>�?%�>Q�=������Q������^>	�Q>��1>7_����Uɵ=�ս�MQ�YU<��<�g�׭�~:W>�'L>���=P�?��'?�?�H0>'���C��Ug5���!��>��=���>Y�ȼJae�J���i�������ɾk^a�����!V>�>�_>��=Nm:�$ω��ݔ���>�����	��nQ>L8>���>պ7=�)�>�]k>L��6�����翖�W�cMS���ԾհϽY��D���_��<�B�>�ܽ��;��,�SZ>���#B������M�Z��>ͽOFO�/�Ⱦ�����Z��ִ���s�a?ɾ��E��m����ԽR6��H��[�H��1�e����+���۽�`��Ji��~�����>v�>��=�k�=�"#?�W�>-д�씸>���>��:>,��>�w�b��>Ž�>C�>�Q ?m�H>8�����ѽf�/��V>���=">�|>6 �=�+����;\L>R��=qY-=)�=�<K��>#=���=�;�ƥ>���=�M)?�����������[�a~&��$?��>Fॾ7�"?���=�\�u���-��������T�ܦr>)?]}?vG><=�=�1������=QF�=�OA� ~�>�>�ɖ�l�;,�s>�j�� �q<2;+&\>Y;��,�>;�l>U>�=C5?AQ?XEZ?e=K�g�־\0��}������ђ�>_�>�6=k�Y�� ۾���^�R��U���Ͼ<��Kd#>)�=R|�=�n��NK���r=����<5`�Rn->���ɀ�<m����=ɳ_=n�<a ^�l�½��ҿ������)����ͦ=���<�
7�e���Fd��ES��������=	�>˓<>iK<>6��=��t���?лY\ٽ� �;׽��ɼ�5��F���򗾛���!ꕽ��:�����v�E��{ƽ�ߗ��Y��U�"����<��P`>jf�>#}�>�&?��>�	ٽ���>'�?='����)�R>J���u	?��"?rV?p�>;�D��7���m�r�>ah.>�_�<��h>��>��������j�=��.1��">QY�=y�kS�׭�=Q̔=����?���,H�A`��U��|	�.�?>̰�)_?��/���*���ؾ+O�)�,d>���>ϵ>�ZH�G�x>��=�q�ۇ��
>(ֶ=��8\�=��=��мM;>Y��=H���%��;_�A��Ϯ=t��>��E=; F>��?�I?��)?�z>f���'�B�7�y��e�N���>�>�>H� ?ҙ>�Ծ�BH����ȾA�Ѿ�ռ�>�0= ��=|�2��j���U�:��q>zG/=��/<3�.>�����=�\>z%4>��=���]}��r��*�������n;��� ��>FH,=�
�=W��<$=]N������l>�2s><l�>��>dn��F=�k�>]'5�s�/��ѕ�4 ;����I���
�����.+��e�>>��#t.�7��L>��>ۼ⺂=�#�OP^���(��Ë>9?�N�>K�> >?2�
?M���z�?Y�?�/Ҿ��J<�+�>S���՗?l�@?"�>��:>�߼��>���Iwy�)�>��>�Qm>�>�Р=�����>����<T�A�(�B=�Kl=R�;=Ko�=4�=ӄE>�Ze���=��>j����?��2�޽v5,���9��>޸r�zF.<�-ؾ��4��@���鄽�Е>��>g��>P�>J��>V{4=�K4�Y3۽�B�=��+�E)ռ�=�<�G ���<���������H�=�c�>|U�=�
>$l	>x�=��H?L	?v��>����N��������*���4��(���z$=�u��`,>1�����^L6���n�ݾ[d��
���>T>Ǫ�=*|x�S<�<E����!>���=����닻��=�¡>aX�>�<>��k>�6>�?ϻ��^�:����i8t����g)��O�}a[�M�I�굛�O c��� �{�w�|_���k�<���=�>��E�2�Tz��zͽ͑־?���/e=p8���r�2˞�^���(*���K��P��;�}�	�ݽ1����ኾ���c�ž^���䭀�����><r>�}?oB�>��>��'?�*+?�R>�;�>&�r>+�>A�Y>�y�>x+?���>Z��>3Ν>�2�<���j)����b��2B=�Qg>R�;��{>�`�=S�5=|~)>�}�=`V>_���|=T|S={.��sZ���0=�I)>w��=Ŭ ?��=J�th�����_�޾,:U���>���-z���w[�=<�U-� �/�L�G>GT��O���U�>(��>ϲ ==�U��$�=���=�V ���=��d=��G>/�?S�{TM���O��0���	��l��5>`Z�=���>G�f>T�m?^%�>�>?�9�������|�؀�8��>dľ%-��I�=�֘��Z���#�X�q�	��Z�fXھ_�<�u�>�[�=j���
����=Ij�Y������-�:>O�{>�6e>�y>�ӂ>�Ɖ>�>��={$���c��ٿ�Y��7񾊳3�䱳�#�z��ϒ=�(C=�m���0(f����4=p�>OJ�>�=�e>�=B?=*��� ��=�h[=h�D����n���:���$�MO���@����P�f��Ż6J�Ls���%0�M�F�mڽ ��>K��=,�?~�?H�>��D?�x'?s��>�n>�s�>B�(?���=6�?��?Za5?�V�>���>�Y?!$����'h�an�<��)=��<���=�`�=��8<C��������`=@9��m
=R�ļ|D�=,м�Mw���G=Ʊ�=Ŭ ?��=J�th�����_�޾,:U���>���-z���w[�=<�U-� �/�L�G>GT��O���U�>(��>ϲ ==�U��$�=���=�V ���=��d=��G>/�?S�{TM���O��0���	��l��5>`Z�=���>G�f>T�m?^%�>�>?�9�������|�؀�8��>dľ%-��I�=�֘��Z���#�X�q�	��Z�fXھ_�<�u�>�[�=j���
����=Ij�Y������-�:>O�{>�6e>�y>�ӂ>�Ɖ>�>��={$���c��ٿ�Y��7񾊳3�䱳�#�z��ϒ=�(C=�m���0(f����4=p�>OJ�>�=�e>�=B?=*��� ��=�h[=h�D����n���:���$�MO���@����P�f��Ż6J�Ls���%0�M�F�mڽ ��>K��=,�?~�?H�>��D?�x'?s��>�n>�s�>B�(?���=6�?��?Za5?�V�>���>�Y?!$����'h�an�<��)=��<���=�`�=��8<C��������`=@9��m
=R�ļ|D�=,м�Mw���G=Ʊ�=_�?H�˾��%��Ӿ��kbҾjX����>���B�`��t��܍�����1l��ۛ>i7>J�>?i�=���>���=[ي��^���V���ѽ�>��=�C^>��M�<�׽]Lɽw�>�i=�ݮ=�S�;��-={y=��=���=��?\v?/w�>�Y���E��B۾������!C6�	��>�L>�_���i'�٨��������4b,�4�Ͼ���ɱ=�Fp>�/�7�>�<@;�L=� /=w�� �g>Ы_=$U=�嵽�3=�8��M!�==�'�jݦ�/��w��5���*����� >߷��������ſA�}ǼW	e���<�'q����=ЄE>+x>�p��r"�=�(>�þ�Fb�=�ɠ�mR��Yg�_{�
"x�b�Ծ���aJ����,>�#E���?�	��`�n�w��b�m�;�����?��?�m�>�D�>q?q6?���=�z�>�t�=O3�>j�\>�{?�j�>�B�>�U��^h>��!=E�h=>{����D�=�>č{��J>xh���û�f��;g�=cy>���=�rfa�4�E�&�л�x�=DT>���=Ŭ ?��=J�th�����_�޾,:U���>���-z���w[�=<�U-� �/�L�G>GT��O���U�>(��>ϲ ==�U��$�=���=�V ���=��d=��G>/�?S�{TM���O��0���	��l��5>`Z�=���>G�f>T�m?^%�>�>?�9�������|�؀�8��>dľ%-��I�=�֘��Z���#�X�q�	��Z�fXھ_�<�u�>�[�=j���
����=Ij�Y������-�:>O�{>�6e>�y>�ӂ>�Ɖ>�>��={$���c��ٿ�Y��7񾊳3�䱳�#�z��ϒ=�(C=�m���0(f����4=p�>OJ�>�=�e>�=B?=*��� ��=�h[=h�D����n���:���$�MO���@����P�f��Ż6J�Ls���%0�M�F�mڽ ��>K��=,�?~�?H�>��D?�x'?s��>�n>�s�>B�(?���=6�?��?Za5?�V�>���>�Y?!$����'h�an�<��)=��<���=�`�=��8<C��������`=@9��m
=R�ļ|D�=,м�Mw���G=Ʊ�=���>�%c�b���� 0�F�⾣^@>�,>K�;>���>�;Խ�Ь��-��G ='?��G��yN�Ɏ>*y�>*��>�P=�H����ɽ�X`=��>4=&�*>�>��� �=N�.=}}=�t=>��+>[�=��<G$)=��m��b���>���>��E?�?E>=#��|g>��|4����A���{���6>��>�9=`���9Q�����M�徃|��{mU��'>��S>��k>k~W=N�?�0YX=O�
��;�pw.�B`=��
�#��<���$�=9�=���_=�Pt�;�ݿ�2���?���X 	>/)޾�ּ�����#��=w����>I_���W��8�=���= �μ$���E޽��Ͼ�ߎ�<;E�Z7��K������;�!�=��C��ͽ��H�ˍ����J��"�^@6��;��5]�\�߼L*�}>^�?}=<=m�>���>�>#�>��>�	�=�*�=R��>�^\>$Zi=M5��ܽ'�M>B�>QR�;%V��U1����<�7~>]F=<��<�n=�"a�9�5�}>A�d���;<��+��ֽ�߼h�%�qu�����=�w9<�/�=2��>������Ͼ{]���"���W> �P>���>�E�>~)��7v����,�Ճ��41<:�>�4u<R�Z�9N�=��R>?��>�˧=
U���\���>T4>�
s>@۽ëf=�!��wp<����<�� >(��= =
�J,M������=b�=7?�D#?�:8?�;Z<��k�(��<)�hM����S���<�Q�>���=^<��U�荾�\�i����E��׽���=�&�>��7>��*>ʑp�c�0�!��[0��F����=D=���=i�o�+}�<�{ͼ��>�s^=a���k@��&�\�3w��퇬�nL��D����۽%����<0ō���#�S\"���=Ӊ=���=���=� _>S�<>�������:�=B{��$����e�R�w�֯/�p�Q���9��. ��\5�E�r��S�<t���,��_ཷX_��$?H�>�W�>�C?���=�/>U�>]��;l�>VH�>��=�z�<���9y��!�=t�>~����䷾<'ܽ��%��s�>s�>Ds�=<�=���<�P)�� v>�=[I=qi�=h�;��뀽�.��	�=^3(>�A>�"�=���>�%c�b���� 0�F�⾣^@>�,>K�;>���>�;Խ�Ь��-��G ='?��G��yN�Ɏ>*y�>*��>�P=�H����ɽ�X`=��>4=&�*>�>��� �=N�.=}}=�t=>��+>[�=��<G$)=��m��b���>���>��E?�?E>=#��|g>��|4����A���{���6>��>�9=`���9Q�����M�徃|��{mU��'>��S>��k>k~W=N�?�0YX=O�
��;�pw.�B`=��
�#��<���$�=9�=���_=�Pt�;�ݿ�2���?���X 	>/)޾�ּ�����#��=w����>I_���W��8�=���= �μ$���E޽��Ͼ�ߎ�<;E�Z7��K������;�!�=��C��ͽ��H�ˍ����J��"�^@6��;��5]�\�߼L*�}>^�?}=<=m�>���>�>#�>��>�	�=�*�=R��>�^\>$Zi=M5��ܽ'�M>B�>QR�;%V��U1����<�7~>]F=<��<�n=�"a�9�5�}>A�d���;<��+��ֽ�߼h�%�qu�����=�w9<�/�=2��>������Ͼ{]���"���W> �P>���>�E�>~)��7v����,�Ճ��41<:�>�4u<R�Z�9N�=��R>?��>�˧=
U���\���>T4>�
s>@۽ëf=�!��wp<����<�� >(��= =
�J,M������=b�=7?�D#?�:8?�;Z<��k�(��<)�hM����S���<�Q�>���=^<��U�荾�\�i����E��׽���=�&�>��7>��*>ʑp�c�0�!��[0��F����=D=���=i�o�+}�<�{ͼ��>�s^=a���k@��&�\�3w��퇬�nL��D����۽%����<0ō���#�S\"���=Ӊ=���=���=� _>S�<>�������:�=B{��$����e�R�w�֯/�p�Q���9��. ��\5�E�r��S�<t���,��_ཷX_��$?H�>�W�>�C?���=�/>U�>]��;l�>VH�>��=�z�<���9y��!�=t�>~����䷾<'ܽ��%��s�>s�>Ds�=<�=���<�P)�� v>�=[I=qi�=h�;��뀽�.��	�=^3(>�A>�"�=4~?\p�8���y���)����\>e~�>F>��'>f�O�g���24���T=���=��ջ�ed>w�q=�q�>P>�j�>]$�=գ�[����l=$ƻ=�Q>a�A>҂I��90����=@�=�
�=7�
>���y���Lн���<��=,(>�3?�H�>�)"?jo:�T�����$?��Y྇�J�9��= v=Zk������z��0O��G<��
��X�������ğ0>�h�>��=�;h<��:���� �M�7]5�of�=B�滽v�<��]�0i��>i�>�jz>Pʽh�Ҿb@��&��"����!�7 �^���w?��ɒ���=1����$��8��������ؽ�D�;���������=~{�=�Վ>�_�=r]>�G=����A����[�
�K3����p�Y����,���[�fCv�/^��;�N�����O)a=�{��Ћ���>��>Y8K>��?ה�>RG >��>d�O<2I�>Ԝ�> ؀>���<4R)<�yf=��޻�ze>х8�`X�>A��ʄ���>:h���+�=>/{N�|�<�	3>Mr%���:E&��HP=�롼x�O�H1u=�5޼��˼�#>�*#?�J�澃`�����o�>��>wC?h�V�Y��=��ǽBGd�<f��
ս�>��>�L>T���[��=��G>�xC=>��=���tP>g�=�.�=9�=#y���'��佽;Q�/*��B>�9��Z_�>�=>,[>=�8�
A)���?�UQ?3� ??�a�I8��'A�T���@�Jv=��2>{>t>ˋ�>$����ž�3��p�P3����E�]5������k�>֣�>^i�=��ȼ(;|P>�����՘t<�:u>���=t1�($�=�Q���+���B>S�߿�鄿�D)��'U�E=<��W1��r$=[>�� T��㮱=C��2O3�^��a�t>��=4�<��=�	��S��UT>`l�>L�>lV�=g�	���־1S����m�ђq���R>wI󽻏F={Oý�y����<[�*��:9��<���2��I��=�|?���zn>��5?9�>i��>�􇽉�q>t���{�����b=s]l= ��>+��*1�>c�=M!�>%-���~��A8&�v5�>Բi���߽+�='�:TIٽEM>��=�j>ʥe��	>�Ml=9����^�gԽh�I>��'>�*#?�J�澃`�����o�>��>wC?h�V�Y��=��ǽBGd�<f��
ս�>��>�L>T���[��=��G>�xC=>��=���tP>g�=�.�=9�=#y���'��佽;Q�/*��B>�9��Z_�>�=>,[>=�8�
A)���?�UQ?3� ??�a�I8��'A�T���@�Jv=��2>{>t>ˋ�>$����ž�3��p�P3����E�]5������k�>֣�>^i�=��ȼ(;|P>�����՘t<�:u>���=t1�($�=�Q���+���B>S�߿�鄿�D)��'U�E=<��W1��r$=[>�� T��㮱=C��2O3�^��a�t>��=4�<��=�	��S��UT>`l�>L�>lV�=g�	���־1S����m�ђq���R>wI󽻏F={Oý�y����<[�*��:9��<���2��I��=�|?���zn>��5?9�>i��>�􇽉�q>t���{�����b=s]l= ��>+��*1�>c�=M!�>%-���~��A8&�v5�>Բi���߽+�='�:TIٽEM>��=�j>ʥe��	>�Ml=9����^�gԽh�I>��'>[�?K�
��@�2��q=��r��Y5>{��>��W��r{>Z	��K�ľ�y��8���lcx>�7�=4�&>
l�=�I�=��>�A3>,����t����j>���=��q>�u�=6�=�ܷ=u3ѽ*�%�/i½݇J=�Ǽ��T>{9>R<>��>����;�?LH<?��>�𱾜���l�6ǳ����P~�� K�>-�ֽ��9�����"�5�<��nU�7!�G�پA�=�>�Gf>�>0=н�� ���}��ߺ>mTZ>U���Ѽ��J=~>>(�J�#aN>�""�����T3�7#�x�޿G���&��ﰾ� �=@O�=��VȾ���� �(��J���a�+X＄�f>�޷=$�>f$�=e�=]�=�ž�,����=졽P��[ґ���ؾ|/������Z�t�Tz(�N��;��缨O�
i%�Q�v��q��Z�T׾�O>R��>�=��>�N?���>'�?U�F�bs?�0E=��=�o ?}��>�0?O}.>m�>ƽ�>�ˊ>c74>(�c���D�QU>s![>���=}{�=�->%&b��{r�!�=@%>��G��C�I���A��,!=��=n�q=��>�*#?�J�澃`�����o�>��>wC?h�V�Y��=��ǽBGd�<f��
ս�>��>�L>T���[��=��G>�xC=>��=���tP>g�=�.�=9�=#y���'��佽;Q�/*��B>�9��Z_�>�=>,[>=�8�
A)���?�UQ?3� ??�a�I8��'A�T���@�Jv=��2>{>t>ˋ�>$����ž�3��p�P3����E�]5������k�>֣�>^i�=��ȼ(;|P>�����՘t<�:u>���=t1�($�=�Q���+���B>S�߿�鄿�D)��'U�E=<��W1��r$=[>�� T��㮱=C��2O3�^��a�t>��=4�<��=�	��S��UT>`l�>L�>lV�=g�	���־1S����m�ђq���R>wI󽻏F={Oý�y����<[�*��:9��<���2��I��=�|?���zn>��5?9�>i��>�􇽉�q>t���{�����b=s]l= ��>+��*1�>c�=M!�>%-���~��A8&�v5�>Բi���߽+�='�:TIٽEM>��=�j>ʥe��	>�Ml=9����^�gԽh�I>��'>�*#?�J�澃`�����o�>��>wC?h�V�Y��=��ǽBGd�<f��
ս�>��>�L>T���[��=��G>�xC=>��=���tP>g�=�.�=9�=#y���'��佽;Q�/*��B>�9��Z_�>�=>,[>=�8�
A)���?�UQ?3� ??�a�I8��'A�T���@�Jv=��2>{>t>ˋ�>$����ž�3��p�P3����E�]5������k�>֣�>^i�=��ȼ(;|P>�����՘t<�:u>���=t1�($�=�Q���+���B>S�߿�鄿�D)��'U�E=<��W1��r$=[>�� T��㮱=C��2O3�^��a�t>��=4�<��=�	��S��UT>`l�>L�>lV�=g�	���־1S����m�ђq���R>wI󽻏F={Oý�y����<[�*��:9��<���2��I��=�|?���zn>��5?9�>i��>�􇽉�q>t���{�����b=s]l= ��>+��*1�>c�=M!�>%-���~��A8&�v5�>Բi���߽+�='�:TIٽEM>��=�j>ʥe��	>�Ml=9����^�gԽh�I>��'>ǧ�>
8콺�X�l���G��v���5>n� >���'�u>kI2���߾8>l��_"�琾xA�:���Z��>���>��[>e�k��,*=����C�W�a�;V��;ݍ<q�=�UQ=�N>n�kt������̽��<�䑼;� >�>˛Y?u??��s>G#�.Tw�Α9�d$��t����>K��>�g�}�������Z��Y����þaK��w3����>�9���ǽ,>(����2�n�">2~>_#���۽��ּ��=ou?>=t�>B�0��k>(�w����_ſ����*���(���q�#�裎�j<��>>�,ݽ�`��z�8��ž� q=�[>◗��-<>6=Kr������f��Ή����nӆ���:�΋��O�9�\ԽU�A���$�A�"�0���>O��U�#K�{e�r#��0����>�^{>��>r�>=?�'?a�?���>�%>l~�Iԇ<!�=bt">:|? �/?R8.?��8?l�?#�ڽ��Ss#����=`>7�=�?>֌M>�R�:�:��)>)F>�l����<���<y�m<}�Q>�Aֻ���=���=�~��.��o"�s)��*Q�p,��Q��<���>��־b$�������X�6�8���ɾo�Ⱦy޾8������Y��>�Ӿ>�̑>eo��:�>��!=7tּ�R=i�p����F >=B}>?̍��%��:��< ���PW�i+��������C��'�=�1?j"?��?����E�\[V�%�H�;�C=+�>~��>�`�>u��n
k�D(�[0�y2��X=Խ��<>�м��>
 �;�ꣾF�?���Q_��h�=�q�>��6�hZ>�fF>a��=���>���<#����=�G��K`ѿ�ʝ�ft�%�*��+���:>�">���>/:C=�BӾ�t�bV�=�`�=�C�<ո�����<�߄=�;�=�g>6[/�5����;�hsD�њ������<Ҿ�5�=��V�z����0����>���=W�����_�R�=྾v���$t>�??�G>���=��x>�{/?���>XX�>�o1��-@>�ۚ>������\"=�Ҽ> �?ޚ?��>�{0<����z&�<�pb�u��=�g >Z��}.(><�p>XrB=���j>=���=��$���G<�K�=��:ZL>�{�>\�>��>>;�O>jtF�4����T������N�2>�>�傾	L�=F����;�
>U�<c�A���>Xܽ.������>
P.>�2M��]�<����Ϋ�=��>uk��[�{=��/>DC>7�/<v�໓H�����f��m�H=��>
�>���=0?$��>��>Q����C
���A��=��`�=(��Wԝ>�ǭ>����l/˾W^�%#'��P)�A�����=��y���K>gd�u2��M��=�{޽C:T=�6>�X!�x*�br��t"=�y����[>���>�z>LV=n8���6վ�ۿ�^���M�����×9�n��g���M��b#���먽⟾Ka�����=V_�>0=a�ý�<>^ꮽȖ[���侅榾�*�=�EA�^s��M���~�:��=�ܚ�,���Q����μ�z�<�:V<�]�����T�W��������=(�>=j�<W���`�k>�_[?��1?��?���=x@�>
�I>#��;�h�>�+�<rW>i�?�?=�)?���>);j>}X��xKF�S\B>0->��j>#�@>��9��	 ��B��L�;���=��K�9��5��=k�H9�;�;��I=�G5>k՛>��ҽ�K��и�
k��3W���<�B)?#���ȟ�=�N�� ɾP����i���������W`��)1羰�.�@+�>�D>Ό���=E̽8F��`�=(�<�φ����<j=vjS�Xy�=�a<�[9�G�=h,;���=y��+>�.?��?JL?{����C�-^���%�
��=L�˽��=���85��fX���Hž��̾�4��C���B{=���>sd��j�|z�>�0�;��n�H>�\�>L?"�)�|��>�I˽�{�í�>��=��=������p��3߿X�����Sǜ�~��@�#>��`>5����ªt�h=��P�=	�=��e>-�>�k�>Wi�>��>>cu>����񒡾Hl�=��M���\�
����9���2��o�I"��m��Q�ҽ�P���ؿ��y� �����'8����>͈�>��>��y>��.?�/?%J�>�=S=���>n��=��>�p�>U�q>��>��>1-�>}N?�?���>o�����M�WYC>�ɷ=%q���^>n�(>YR,�+?н�d/> >N>K��=:��=����N��-���C��=\m_>n"u>�P�����h����8������NֽC=�>'M`�w��
��\�\
���4`��(�����_g��䒾ݸ(��>�ڌ>t����ٴ���)�"o#�Hb��
]>v��=lr�=S�����<��>�?���A�� ��=�x�9��<!f�=�|O>�(M?ƹ�>��>j{��2���Y�@�"���=��*��h��Z�ZS_=k �2�T��w���l�"�(�����Ľ�<� �=� T<F�g>~c%>�>�������*����
{=�,<���>>�2�>)�1>X��=a�M<��:����묿h*,�i)�F�վČ*�{P���&��_�׾q+m�_�3�������龛O�3W�n)�=3�>ќ����0�g��쵧�b��g֩��Dd���=�Rc�AN�)�1���_����ƽ1x�Q���W��Ͻ�!��<��?��#>5��>�5�>K�I?�BB?��%?�u3>��>�Ȳ>i�?��?.��>oB>���>�
	?m�?��?���>��ý��.&>ݴ=溾�ɐ�=�/�<1�ٽ`nw<U��="�=��P=������=�g�:��_��Si�<�(=��J>��)���������-�܍����>fM>�ߗ��&�>�&��v������"l���b>�a�>���>"]0>(.
��s>�q<>��s����
�>O�B;�e� ��=�l=QaM��[�=̈�=��t�vA߽����i?=��>��^>���=��P>0z?3�1?Z�;?�C>�>��G\H��3�~�>n����π>a��>N5>@2��&��0��<�l2��>�>�48��s'><�Ἂ=IS$��	����=0�=���N�=�j�=��=�}=��K�=�9&;q��=bȴ<����Hп�(��b��>���#����_�=eQ�>kJ�=0m��_>O���Ǫ�z��>���>�15>���=�ޔ�9�#�lk&�[�������΅��5����9�:Ղ���>�|;��a�%�8999�&�����۽�黽���;����\���	��[�>�r�>��!=#�b>��/?�qR?=�9�_~�> xD�B�?-�y>n��=�{�=ik>eR�$��>RŤ>���[�'�a�����B>��`>)P3=IQ'>:.>��Z���ͼD�E=�q�=�e�F�t>��l>�7'<r7��DgB�'�ؽD1!��A�>���<�8����{�U��k�No>�6(>a7��u�>m�Ǿ���
70�_�Ҿǚw���>A:>�_>���=���>�r�>S怾A�e��Iͼz�X=��>��=��A���q>N�T>����腾�Iս�8�=��=S�8=�S�=]ͽ��>�k$?�!?`�>+��=�Ǿp�W��-�= P;g�����>�*
?楦>��ʾ)�"��K��D����
�>��,�B>��=G?�;B��=���"0L���J>���=J�н��*�=)>�s�=�=B�?��J�:�y���l�=���Eʿ��ܾ4����K��h�>�<�>��i�hb>xO�>F��� s��@�>h�*?��?`Hp>
т�e	�1#���˾镊�[����ѽ�q���v��ڧy���B�����5��:���Ɍ�)K��dO������뤽���,���;b+�>s�>��G>Ei�>H�+?)� ?��_>���w��>N�Ľ��>iS�=S��=:��>^�j>(�R>��>:��>0Ӧ�l�����%>��z>�D�=��A>� >��r��W�<B��xq���P�=pq�>��->�Μ;�B����S���'��$�2a�>��	>r��uN�������]���>X��>o暾N����՗=�����+X�������52��k��玨>G߷>�8�>�o�>��fn=���/>l��2�f�
C*>Q]ݽ=�����=2�i�Y���)���|��N�=���<�՗�S̃> !?Y�T?'��>
���q@���f�F��n��0��>�@�>6w�>Ó>B.G�T+��I��G)��Q�1�:��r9?G>���=O���.��<�=t9�� k=�>����=�>>�>�u���g=5���_m��OJc�կ=�ο̮�;�������i=n��>� {>z%�r���������/��z�0���?��?}�?�@�>��>��i>����4��ݽ�]�g� �X��6�\ ��2�������]�^�]�g��)8�*]�qߟ���&>'����G½A.�0<�>\�X>ύK��L=>eiE?5�8?��>A�>�"? ��=0�=n=��_>J��>,��>Ab(>s��>ڢ8>8 N��������(d$>���>��V>�a�=\I?>�恺�%�;[)
>P\���[�X��7�P>�:�>�q�=0�=�*u�=�!=�*���>Ǿ��%��F�"�F�٤�!u�>���>8���>����p�!���8�A!1�Kz>�Q�>%N�>��>�0��cr=��+>��������#�=����������d>�{�=a��=��:>>Z��l����%��w�
m�=3[=Ax>������#�%?k�?�.�>I�*=mŖ��$B�
F��xL��x�����7��A�>�>%��nV3�'6B�@gH�T2�,��>!Q�<�t">��H>IZM>/2w=�*�����<F]����=���
Z����<�s=>J�>�> �x<4��=`����=�����䒿�F���ư�21�)�V>���=�0�@W4�Y���݌�<r:� �ս���=�`	>�>�/�<I�0��o�>���"���=����־�`��4>߾:eh��Ղ�A=����>s=���Ö�/�Y���1��J��tQR�R�>#?���>�>lA�>fF?�b&?��>�h��0�?�i>%�>��>K��> H�>H܉>��0= �_>���>y	�=g20�=��-��=צ�=�c�<(�>�K�>h��7�\���Ľ#�R=�P�!��=4]Y>��"r��o�QA��p�t�y>���[�#�wns�a�M���(��>�*l>©�m��=���;�����8��0���Ǿ�a�>v?�q?�=�ϧ>kpc>�Vt����Y�>���<%�T=�ߡ>q����f�Y�>�6ݼ��z������E=��>TN>}�4>�Q/�7�>&!?IR2?��>�K<b���ՙH��ǾERt�M���?��F��>4%�>�_��
j¾�[���/��E���f>�O4=�+}>���=�e��ϥ��i��1l4�� >x�/>��3>���<�8<ؗE>�	>�I>	'���Z={�<�0�<�6Կ����o�9.��<"=�냻Qv:>�썾j��=Ԣ�=�l�#������=ʠ�> }�>��R>���t���̟���)�� �^�w5/��o��/��ٝ�����W1��<��� �%>����t��
��M�¾nm���R �/��ͪ����=(��>��>�s=� 轐b)?GB?!�&>�\o>�?�B�=�H�>d2�>��>t��>���>��ƃ�=��>OW�<L���#:����.>MZ>�*G>WUL>J �=�	A�斻�O{� �W=τ>�*�=F[n>l�B=���p��+��*z<Yb?�N⾬
Ⱦ����J�s�<(:�>�mA>Ji��ut�=��+�5�L�Y=C��=� ==J>#9>�m�>ٶ�>Ɩ�>d��=�	ξˎ=�B������* >�]�;�zs=�ч<�� >>y��=��>2��=7^J�N"<�)>� ����7�n�$?�&?�EI?(ǰ<W�߾=��xR�;�M��c[���E=����Jt7�4��;sӾCE1�ƞ0��Z��@��y�=n'�=�M�=��<-��a�퐝���=��}ν��8<���=HC>B@>:Z>5ԓ=�N�g�i���0�@�Ϳ<����C��H�B�_=���(X=,Q��N����=��<,+����R$>x�U���=�V=>:��m�=�վ����jՌ�����U��!n��4̾�#.���X��ظ��H��V>��/|���e�T��,{�;�����b��~J���>��>�,0>���=C�+?��>�*>o|�=Z�y>��)<�jK>_ �=.�W>��n>�B�>)��>:�>+>�@���'(��׽�D�>���=>�y>Ε->��h�@j
>� >�w�=7u�7��SU�"O���=2�>�y(>h,�>�?Ⴂ�1Ǿ�Ⱦ���O��=P#�=%J=b<c��W�> ��2>��L���a=GK����>�LY>�G>�W�>z�>"2>�ҟ���<�<�B;���0=&�=*�>A�u=��4>�I�=~�=溳��l|�!�K�U+�<s�=�]��U��;�"?y��>3=?�����4�\���(�y� ���(����Y>aBx���o�s������TN�Ů2����,E�S)�=oW���X>�|����ͼ��6�$��et�<ā<¡��)!g=��><��(>҆/>^�>��>�y��eb���u	���տ�R��"���&վ4�:��]�=<r6�֏��`S�a����-�E�2��A�<��=��/>�=(��=���<��<>b?������H� >om`�[ܽ���Y�Il��<��i8�2F��gM�Q����G����? ?����� 0�����0>��>OR�>��=p�?�&�>
��>Y�{>���>&.%���%?T���_>��~>�x>�c0>xD>h��=賡�G2�e���,>)ڴ=5D>-�6>qG=� �Gn�!�=��`=��"���ؼ�1���<��h^Z=V�@>0�=w�o>Y?W��F�ݾ�z���*,�n䯽p(�>�;I>ʷʾ,x=�;�y�=҅4>�X>��R���<#�n>'��>߱�>�7R>�+#>Bq˾���ɏ=�3��>ᤶ<������m%�<�R�=���=�l0>�`'>�}�=��1=&��=�Vi�w��<5[?*B/?���>V�ڼx8���v��{����E��:\>[��=B�"\��]	���0��:*���9�(�(�龍���G]�=)C�>�N�GJ�=�=�={�z��ν$��n�=ࢊ> �">�N�=�ol=�O]=7�)��L�𸻥�=��ܿlL���q��6y���Q�i�5='NI��x�3=m����=���������=_`�=���=Rc���Yɽ��=��>�=��=Q��&��~��p�˽�,>�Na���+�C{���T4�U�S�����J��_n�LS�m����j�>P�>��	?���=��e>U$V?�ۭ>�G=fQ3>1z�>�襽���>]>�9g='��=�A�>�^�>��>�QH=��5��Ө�ܒ��-5>G�)>�9=nP>'k��I��;R>��>L�C�M�潵w0��*����=�t�>�8�=���=�w?�'�����f^�����,�Ǽ �>C��=n諾fZ�>$����$>���=Rd2>�b�����=��=>���>�'>஦>\�.=�Iо�������=��:���=�<9��=�3�����<^�>�bD=#�=>Ǟ@>�J=W�A�	�<	�?=�9ڽ{�?�#M?:<�>�Ɂ������y��N����0���I�=���� �P���l���^����$�?m/�/g+����|����&�=Ĩ~>+�p>R/B��'�<���=P��Ք���>��=���<kO>��ػ�[S=�G�=�>���=��>qkտ����*� zh��E��A�=n��z�D8>)����V�i�{���D�B>�D�=va#>ģ/>����&���g�r-d=��=�y;�-�V�b������ʛ��w���'�u���Ǜ_��7y�Ɩ���>���! ���9m��� ��z>ץ?Bټ�>�x]?pD>o\L�E��>,6H>E����>d��<4>�'>���>׃�>}�U>�>$�>�_~�E7���?>W�;>�3���t>�M�ݏ	>�aN>�N>#-E=��v�ٸ��eT���ж#=u��>a~��>��l�)?3�&��Z�\{��'�֡&=y��>��>�A�=O�(>����>�8�=�R�>�!	>��>.%+>���>�κ>��>`ĕ=����S����ڽ>�=�4,> ��=�a<�
�_[�g�s�=>$�*>�w�=>Rk>�͎=�@}=��+�$;>�s'?��9?�CY?���>Y'��8��jL���o��<"��>�\@�Wr���_��	��cJ���+���1�'��� R9=T_�=��f>�EL>���={uN�pq�=?Ք�*Z�=��r>���>��G>v]=�h�=�`�>���pf(�P߻">vݿ�>���񋾁,v��佟��= '�Zn뾼�}�h8=H�>7+�R�%�}|=F�^�b���~�����=8Kz=�G����3p��փ��\>�� н}�'���ս��v����[���.��u)�YN*�$�#�N����XڽPt��dE^�e.�>7�?�)3>�ʱ���?��>�=�F->I>�왾�|�<��D��>��>i1�> �>�x�>̇@>��X�Ku(�9i�^�>z��=غ\>�K>��I�9�k=�w>ߤ7=��M�Zv�n���* ���y��n�hE>l���y�<J47>=�j�s=�J�+�D:�[;*�ɜ	=��2?-"־�yӾ:I:����a�0��߾Z{ѽg��z�C@�<H|d�ׂ�>���>��1��/�k
�K�o=X��=��>%L{>G�1>F�;=��a���y�~������
֔���>��V<� >'sj> �5?�b[?D� ?�='�8��xY�$L�;�)�lM�=-zO=1��>e �>��|>�k��&�4�;��=��r�<P��>��=���=��>� Y=�A��Ie<��">����"H=(>�"�>�Q3>���=po>��=�#V;�L��ͭ�����T��������Ƚ0�>�!\>��~����>h�>\�z�v���]>3C>�mx=C��`Q�8�B����Ĕ�d>�O,��	���*��w����A��!������%��픒>�0����=>��Ƚ���#�pǾ��;(��>� �>���=�>�)?m*?��>��=Oi?���X�H���*���>KS><�μ>}?� ?4�?Qv�>`½�����$<X��=
$>o��>2{�>�W����.��W(>��޼)��㽗S��F͍>%V>iTD>D�>��X>���=������<�"���O�Sվ�z=+�.?U꒾p�������=�*+��ՠ�Z>��F�����Z�P�-R��,{7>��C>�/�R���U�޻�>���=*>���=�?���=�dǾ��R��k��vP��a�<x�=�+=W�1>��x�WA(?CG_?�r(?Չa>�9���e���F��Ԡ�">>U ?=S�>h��>�˾8 �d#$�k�O��yX��!=`�a>�Ք�-e�=6Kp>��:G�ݼR>e"(>��b�>R�>���=5�:�X�=�%�>�=r�=Xi�=U���ϣ�0���`$���k��'��*W#>��w>�8��w>��=V�j�I�罢P���>>,�q=Ъջ�װ=�3�=�C���h�z��=���������w��U�
�Kq����=��b�y:�>K �������Ǿte��.ξiÑ�t?��>�%S���_>�
,?}i3?]��>�꘼��>}�\��	a>q���� ?��>O,�>~43?J?��?��j>�����j�A�$>J�a>�>y�>��>��L�e�ɽ�V>��S��q>�E�>(�1>���=��x>b.�=�[>�
�=��><��>KY�)j-�(p^��������%?�@�<Ff��K�'��z�=���[�˾���Iu��W����[�,�Ƚ���>��>�`���Ǿ�sɽ�B�>��D>oY>�k�>%s=����C���[�O@���;��Z�2M>8;>Д>հ���?�s?=?k�i=�W�OW��^���~v ��Ϗ>���>@6>X��>IJ���x���Q5>�jR��v=�oN>��=�o��ż
�P�$�@�{=�=�D�=�@=>l�>4T�=�B=l	�><s����V�mlϻ�_��$H��c��@���O���\���弄�H�;ڃ�\v�=/�~��@	������=��=�\8=a(Q�!�e������y���\�E��=�>�c������	Ҿ"+���>�����<���4>�?	���=�=��p� $t�B8��5��Vs�>�7��>{��_>D�?�1?8(?��e>9��>w�X>0��>ź���Ո>�\:���>ς?�]?�,#?ӯ�>c��t�a�.��=3M>�0G>���;�p>���pN��x�<���=&x�=-P(=Y`<�e�=�͘�۲���Ĝ=�%<�K�>�)�;Rz6���!�,�V����ѱ�҈ ?�H��)M��"��ئ= �K|��r�;���v���ҁ���R�y�>��t>����������٣�>�>�ߐ>�c>�2����T=�n��b:�<X��3�qq����>���=� !>�9>�5?�$?~28?+O��z���]�0�V�f��_�`>���>\R!>�ן>���>��f��8�b�%� ��~G���۩;<>Q����=![>Qw�=?���f���u6>������{=}����W�>��X>�FR>��B>ۥ�=�"r>�O>��ȿu����=�T��&���)��o�d�����0�����>����]>�0��Uz>�?���V���_J�'\)�8���RRM���A��4V>H�c=��������d��$;�/7���7�������̃>:���M>~���=�����龰���,���>�O:>笈=>��/?]kJ?��#?d�<>��?H�}�=��>����=3�>	]�US->�\?�"<?�q)?��	?�D���<�j8�=�U�=��B>��
=�7N>��ʽJ�;�[,>��=�Ͻ=*�����AJ�<�ܿ��>�<=�=%(�=2�0>휫��x1�� �[�@��+&�oj����??�cr��2��[&2��+]>j�G�m��I�W��7%>U�G��[�������>�A�>TN�����X3@=�q�=ܑM>ڡ3>;q���཰����]:�!���+�8 ��1�=��;���= ��>�zj?V�:?bE�=��9�m����@�đ�9��m
�>kR>�>�=Y�c>A5%�����*^��Y㾑&$�/�-��ޡ����>O:�=Br><��>o�=�x�^��=QP>���q�>�K�=f�>2v��P�>3�>VH >��=�y(�kVǿ.��uuR�H��-C���Mf=���=�b�O�Ⱦ]S��*��=�'>�q�>����!E={晾�q���$������͢��P>잙�����wg�����r�.�[�ƾa"
��{j�W�>�ك�e�>.������������$*��B�>�+��9��=�6?r�N?6?-�?�Bֽ��4?�i>�P?�J���ð>��)��"?��?��4?I�0?�J?T&y�c]��}����=0f�dK>zϒ>Sf���U��M{>H����;q������<~�<=6��;�O�=�YK>�/>���>t���쾯ׁ��W���֙=Z�>�/)��$�����>�}���7��A�n�(	>$j>��>w
�>/��=�l�6c�>�T>�x˾�ݺ��T�=�t>P֤<V��=�Z>��Ѽ�t�=2a�����<���<��=9Y3������m�<`��>�F>K�7?��?30?x���+M��X�*ͭ� F�>�����;?2/�>��0>X����"�G�����^�����G�=l�>��ۗ�>S׊���A��V�=OD�=V����r=�d>��L�/vG>�Av=�6�>n5o>���=����{žn�Ϳ�)V�"�>v�\�U/>L쾀c�=����5O���������<$ý"h�ŋf��u3��[��c�=�h�>T�_���ᾇ�ھ�>��"���d��ܾ���u���������<��砾�ܧ�)RD�^���S�h�2G=���a�
��͇>�ٜ>ޓ��[�����>��>h{v>-Ic>.��>�Ԃ��>���=��>u�z>�g�>�$Z>>#�<��;`j<>�w�rȼ���>����<��<>�~:=i�Y�x�a>����5޽P��>hU=t�H=�=5���t��F�7=�$#=��?��0�r��V��9z��百T��>�<�=LX�a,A��:���%�۷i�~�?>/|d>Θ�>���/�>��?=�x>�?>?��B�����}��&o>����1�>�>�zI��"�E�3�R��M�Fh�=+���R��wJнZ�(>�@=C��>�eB?��2?�9�1��k�ǾU&þ/���Hи���<��E�R��[�Ӿp}+����?-,�5W���f��{�=x��=j�\>D�=���.{���=��ƽ=	=@!�>�(�>/�;/`+>�~>�+ �N�>M8!>��={PJ���ῠ���]��F`�>��==J^�=��J>� ����g�~��>Q�B���˽�f>�h<=����_.�=�ƽ3H޽���;��vۘ��Z�� К<@�f��_���ݽhz?����Gp��Z���3��v����P<�:���U9�@I�'6�<廬>F?%A�=
���>>EI�>�I����>C[?�p�=O�?>8?�=����=��>yNY�j2?�M8��.ɾ]w���Ž�R3>�ǀ<�B>#�=�=�r������}�; @Ҽ��=Z��;h�ۼ`s"<2n����<�_������>�d��]ྀ���O���ioL��>$V>�y�
<�=�e�p�[={uP>� U>?�ܼC��86>J�A����y��>�@&>�u���B�@J��1>o�"=��7>r�-�m�����O^F>�>�>9�{:� ���M�����ԾK�\���2> �)?c�?1�Q?B���
�˾Fj:����������=�?�>�F�7W;�~����!����O�j��c^�_b�;�a�>a�<��ý.>dB���O(�x���ذ�=@��=�V�>3����y>�pa>��u>`���l퐾��6�~`��kڿ��P�ɣ>|���S�>�ɾ�ו<��iϩ�g�L�w������!���_�p�̴Ծ��<��#=�I�>BMX>�g;^�X��c�=�	½K�W\ƾ����?G4����L%/��H���Պ��Z���B5���I�?>��;=�J�=������.>�^?�U���$*����>�H?rJc<,�[>���>��UU�>r>�/��z!�;�l�>�O>�Jf=ۤn>�ψ=�����q��U�>P��=w�#>z�S>[�@>(���>��a=��q=[�O�G���9�������=}_>oԉ��g,>�s�>�{��b����松�?¾ꚃ�k�>^�=��-D�=���}
��S�=Ĵ�:M�ھ����>�gr��H�=��>d9>���	&T={�=� �}�������4�\��_�"����</�=���=�Č=�>>��<a�b��w@�@�����>��?7�?��V?׶=��4�sn5� R뾊E>��W�q3
>��޽3���U}��"��=�)��v�����{N�;�0���>��>�ܼp��>X7��Nf�*(>� �=��V���g>�>Bi罪n����4=ߎ�<�7_��p�=�u���Z��xe��M&þ�޾�ݘ��ѽ�@+>��r�h�z >��x��6.�<5	=2���gH�>���w�=�`>v�Ҿl�p�@#<�ҍ�"�����"�g�M��x���Z<�墾��)�k�A�&�p�^��Ȼ��y�n�$��:;�WY=��	?��>��{<�d?�3?��&�+)>�2?\�̿�>B�=�w��Dy<�Z�>J�w=(���E>�,�<t�x,i� 1>Z��Ƴ�=��>� >�BH�B�=��4>ˤӼc8�HT;�(;=���G����>ʫ2=�6�>���>�w��B8��ِ��.��V��<"��>!x�=��G���Ą�>1=�lD>�����������=>S�޼@�ͼ_�>�LU>�I�����P��.9P�ʏ\<@�=J�\=�R�	�L=�S>��)>rƼ%$N����Uq���,ܽ>�/��uR>�?� ?��"?�[�z�þ>�	�B譾����Q��"r=pI��В1�����zu=�؟�+n꾽	���ƽ�AR콖��>��>t �=l!>?�Q�k����>'U��ν��,=��=�k[=Q� >	r>��>K��=\6b=C�I��M�Q���������[�뺺��6��j��>5�"�j�o=u�?�f��2�<��Y/�({���=+�M>�(��=K��=�v���퍾t�=(牻盍��yn��G���`�ۏd�%�i=�-J��A�]��F�Q�+�@��;�f<k9<���[>�� ?�	;5)K�|�?%�>�o��5#>�>�>�e��'�>���=����Xc>,-�>'ۓ����=�D>��#�����P�hy>y��뱘=K�,>=D�=mb��t�>cS>z�;H����D�;�i�=�G=�,�=��=���>L?#O������	�j�L�U[�=! �⣵>ì̽\�k><޾c�%�����Y��=��>t�>``�>���<zF>�>��1<d�l���)�Xb.=IY>���=s�=�T=���=vN>l��r�;��0ǽ�j$=�?>�@��%�<�j��'>lM;?��C?w�&?�R>��7������KL�s�x����>@^�>夾=�&�97��S���9���ݾ��A����<��>�S�<���=�+ >b(K���̽K�r=.ڳ<T��<o�4�%l	=jj>��>��.<HYB<��S>A/Y=�6?��>п�|��>߾|Uо��<��M>��>3�g��ԧ�����C�!�i��=�z>���>i�=�2E>݋�<џ>���O@����ڽ�"�==U�����|d�[���2���,��	�����T��"�p�Ɉr�?�G�\O^��b�#��V.��B�>���>�ig=�[>.�D?W��>�i?
?T=Ը�>n��>0E
>��>�`q>?��>,��>��>ɣ�>��>�T�h�'�l��^�>+C��Z��<��>��O>�1���\
>�&k�&�=�=f�&>[>g�>l�<!�Ѽ۶�=�x�>L?#O������	�j�L�U[�=! �⣵>ì̽\�k><޾c�%�����Y��=��>t�>``�>���<zF>�>��1<d�l���)�Xb.=IY>���=s�=�T=���=vN>l��r�;��0ǽ�j$=�?>�@��%�<�j��'>lM;?��C?w�&?�R>��7������KL�s�x����>@^�>夾=�&�97��S���9���ݾ��A����<��>�S�<���=�+ >b(K���̽K�r=.ڳ<T��<o�4�%l	=jj>��>��.<HYB<��S>A/Y=�6?��>п�|��>߾|Uо��<��M>��>3�g��ԧ�����C�!�i��=�z>���>i�=�2E>݋�<џ>���O@����ڽ�"�==U�����|d�[���2���,��	�����T��"�p�Ɉr�?�G�\O^��b�#��V.��B�>���>�ig=�[>.�D?W��>�i?
?T=Ը�>n��>0E
>��>�`q>?��>,��>��>ɣ�>��>�T�h�'�l��^�>+C��Z��<��>��O>�1���\
>�&k�&�=�=f�&>[>g�>l�<!�Ѽ۶�=�x�>L?#O������	�j�L�U[�=! �⣵>ì̽\�k><޾c�%�����Y��=��>t�>``�>���<zF>�>��1<d�l���)�Xb.=IY>���=s�=�T=���=vN>l��r�;��0ǽ�j$=�?>�@��%�<�j��'>lM;?��C?w�&?�R>��7������KL�s�x����>@^�>夾=�&�97��S���9���ݾ��A����<��>�S�<���=�+ >b(K���̽K�r=.ڳ<T��<o�4�%l	=jj>��>��.<HYB<��S>A/Y=�6?��>п�|��>߾|Uо��<��M>��>3�g��ԧ�����C�!�i��=�z>���>i�=�2E>݋�<џ>���O@����ڽ�"�==U�����|d�[���2���,��	�����T��"�p�Ɉr�?�G�\O^��b�#��V.��B�>���>�ig=�[>.�D?W��>�i?
?T=Ը�>n��>0E
>��>�`q>?��>,��>��>ɣ�>��>�T�h�'�l��^�>+C��Z��<��>��O>�1���\
>�&k�&�=�=f�&>[>g�>l�<!�Ѽ۶�=�x�>��j>>j�k�������T��@���׳=�>?~�=m��>3.����3�3��Ӿ$�=´�>&
?]�?-�p��؂>�b>�YV���:=�i&=0��=>�4>s��=)<�=&��=��!>i�d=ݶ��C:�׿��X��<��l=R�;>��.�"�a>\>E?�v�>�;(?��>���3�3�����R��=�B����>��>��>�Q?�lGK�͔G��M�P�4���z=�J+=��a>Uo�Z���m>q���������gy=�X�=��X<'�=�>�>9g>`7'>��V=Ȅ�<�O�h�����Կ�$��7��=�~�Ģ�A�j>�-\<3W=>Td�����������e��Ӣ=�-,>`>��ż�e=d<��_>�˾il��]�%>t���4��ҷϽ䋤�xڼ�F\�UW�쬾�{��	3���[l��\{��ȶ�㳒���X�;}��ϸ�>R�>�}���V�>0(?�� ?��?j�R�ŧ��������>œ?��>��	?���>�Ҍ>D��=n�3=�
2�4	���:�~�4>��.=Z=%�A>��<ݠ��40��W����<>O�<m>=�.�=Հ>�>>��=6�?<sT�>��j>>j�k�������T��@���׳=�>?~�=m��>3.����3�3��Ӿ$�=´�>&
?]�?-�p��؂>�b>�YV���:=�i&=0��=>�4>s��=)<�=&��=��!>i�d=ݶ��C:�׿��X��<��l=R�;>��.�"�a>\>E?�v�>�;(?��>���3�3�����R��=�B����>��>��>�Q?�lGK�͔G��M�P�4���z=�J+=��a>Uo�Z���m>q���������gy=�X�=��X<'�=�>�>9g>`7'>��V=Ȅ�<�O�h�����Կ�$��7��=�~�Ģ�A�j>�-\<3W=>Td�����������e��Ӣ=�-,>`>��ż�e=d<��_>�˾il��]�%>t���4��ҷϽ䋤�xڼ�F\�UW�쬾�{��	3���[l��\{��ȶ�㳒���X�;}��ϸ�>R�>�}���V�>0(?�� ?��?j�R�ŧ��������>œ?��>��	?���>�Ҍ>D��=n�3=�
2�4	���:�~�4>��.=Z=%�A>��<ݠ��40��W����<>O�<m>=�.�=Հ>�>>��=6�?<sT�>��I?�m;>Af������� ��G�=H�?f�=9ǽ����>�壾mUA�,�+=�� �
�?�
?r�>��>Ow�>��i>�y�-뼏�O�]k�n��>�4=.�I��)�='�J��$����%=,�w��I��@�=G�B>�R>0���ʔ>d�*?�Y?G<?m�	���ƾN�&��$�Jb��:��%u�>�>|���Ɏ�K���`����ҾFe�m¨��c:��M,>�ީ=#3=���<H�=O-��/�>�4�>8W޾�y\��n�>#=�$�>�\�>�L���%9��˾�6���*��������ؾ�.Y��B�{��=�߮��_���ʀ>�.l��%t��q>10�=m�>>��(�*�������`>����K<�(9���/���0�
[���+���^�h���a��@��M��Y�A�����8ٽ��O�����.�=.���>>���>�=g>�$�>��R?*q�=/͕>u#�>�f�>�)����=��>W�=���>ME?�
=��ɽ�qܽq�k�*��j����`>�N->��>F�>�y�=r���_1�#:�>�}>_)�=hv���,�]�=�Bt<���=���>���>ؚ?����7���j��.�>�G2?�D=���:��'�>1{�K$ �����Ծ�rA>'� ?})?�k ?���>�:v>E��=mB��8���㓼9>IY�=��=��Z�z�~52���޼��e�b����=���=�϶<2��<���<#�3>�S%?�A8?�oJ?Gm��p ��f�/����=8N��8>�k�=�!��UL��D�)Uݾ$��C�o�B���y;>��J>f��==>&�/sO��9�<��#>񥵽5f�=yoa>MY>5%>G�=������`�U�I���׿fU��������3��kW��:�۾�鼇���=�P�=�O�=4�Q�M>�%>�7���ɽ/���S=?t|�J��� �ϻ��罦ʋ�f���|��xFU��)�w5$�y4S��� Y�"b�@^���ؽYu.�$M���a<֬�>%`?���>��h>>�*?<��>�@$>\��>�?͡H��1��B`�>���>Jo�>#&l>�V�*$+�G!>�P����5 �t�I��oɼ�$�=@ϸ=I��=�Y�=I�>�ʻ=[������EB��7�<��2�趼4�=m>�^��L?Q���y��f�<��dK���>��?>C>�5��Zz0?�6��IF�jU����J���>\n0?4�?"-�>s��>F�>�`>E�>��#�Ȗ�=�~�q�p>���9��=2*���l�=c�,�ڻ/�G�>I����
>n	:=�*�;��>�&wu>y'4?��)?,S?V�ʹ�4t��1ڽ���	ؾ�z? �q>�Y���O>:=9�(���D�\��Ͼ�D�=��%>�bT�F�e>E�:�X�s�%�|<R`T>h��=%�/=���;>���>�O:>f�~=�Vu����8�g�L��fӿ����8A,��Ծ>*�>Kڔ�=i���o��๽�ڀ������=��4=!�a>+��>�xӽ�����Y>Ƃ.>�����f�\�!=�>�AJL���l�C����D������� ��t�(�fVѾ�����;R�ǽ�<��x{��zԽ� Y=$h>��?��>A�?�3&?���=�?�>$-Q=�?�R�!��>�?�а>���>�>Ӄt�w�
>�6=r��Z^������S>�<�H�=]Y>�ǫ��w�ͦT> ��<
*=�Q>"k���q����	<�x���-}=��>\��>�?SU��U-��8���?����?�l�>������>��v<E���"��ֶ�p�پ�)�>eO�>�<?��>&Ħ>7_>RH/�GY>GI�UaW��O=@Z>�����*������*�[6ӽaH=�^�=�p>ݏ>`J�<�К>�L?��,?@99?	�Q"��T��}��*9{=��˾�Uo>��=>��<��i>׸����ڦ�8Q:��5��Z�u��8>�5y=���)�C>��μ	�:=,v�=�=�T���=v��>�ڡ>��>�W9>P���'���Y��y鹾7��W���{eҾ@���s��=U�y=V�~�@K�,|:��U�=�t��i<�n>�����J>ZI���󽯭�<_=>9����q���6���㈾�@h\�
9
���I�=>��E�ν.ٚ��-��5l���O��ٽ T3�k�~>-��>���>E��>kx(?R�>	���;>�>��9�`1�����>���=�d>�3�>ĉ�=	zc=�G<F轇�d�����>r"=[8=G:?>��<=Q����=}�%>��=>���ꕽ�?��wŽ�T-=	��=��=�l>a� ?��m����s�1��a9�K����ʸ>R[�>���=��/�K�ľu�|>�/�gT^>��4>#��=�F>�#���g>H04>� Ⱦ�5��ƍ<]P�<b�>��=>y4ƺ���:��E<��e=Dk���*>�[>���=�Ѓ=XK��#��+��=7�M?��?<�B?@�(>������R�A���g��۴?gz�>Y��\�w<�@�^a��x��&��d��`�B�z=�ϙ>��6=D�>����c�π��S�>Uo��>�$>8��>`M>.�>�, =}8��OR���i<�T->���-��-�r�V챾KN���ipD�����#�sY>�ӫ�${(��Uf��5�Un��#e��p7���_�=v|�>ڟ�f^<�#>uM$�ts߾�̾3*��x2@�(� ����<9�ѾK�����F������5��u��S�X=a>�+�=LV">!�>U��>D�?� ?�(�%}w����>O(켜,����>nR	� R\>��=��D>�i>�2>�F4>dTd��qo�V�=٧d>�r!�k>X��<gkͻ�E�2�=P-t=;Ō��֐<�7��9�əg=�n�=�>#h
>�xx<�wT>b1��P�MM�D��Y��>�Y5?<��<��f�<��!Ž�Ww����n_<W�r<�'���Q�����j�>�>vnc�9������=�\>o�,>x��=��=���������k>�-��j������Z�O�H�j=#T;>�@3<��#?wF?kX�>�ȽС��;��4���Бa���"���޽1�>�՘>a����5����G1���þ\�Ľh,d>h��=gV9>�0W>�5�3Cν��r<35�<-Y��N�>�;�=���=g��>p�>A��=	�+>��I>L������#���9<eХ��葼)y8>�wL�^R,�̲��w�'�������������>���=��N���?���Ǿ=u�������Ӵ�<�[j�'G��8Ǿr��.m4��⻽N��<X+پ�ϴ���c���;�V��9�x=�-��=��,�c���?�?ؽ�77>�
?_�9?��?=B�>��a�W,�>�\�>?X֟>�aT=X�=y1>*��>nc'?��?��>6��:1I�2�=�jX>a�>}Ro>I�>�^4��ڛ� %u<露<���<�5���3�N��'̮=+G�=���=�.�=
">m���9�z�Q���g��!����>?n�>�a���ν2ྒྷ~�>pn ������&�B������>0��>S�:���
�b�׽��=��K>��@>;�=Uq�=>@5>�Q� �����!�1�6��5N�χ=t�~<1DF>�e>]W��=?�j?��>��k<������6�<�����"����E=��=���<�cp�#��p��
����:׾�gܽf�>%���p}�W>�%>�������ǃ>�i���>Ƭ[>�;�>���>�x�>#T>��>>D/ �.�����ԿTݰ�a��r�����u���C=�WU�l���PL"��:�mξ)���� >�w�>15,>=�?>�L���c������b޾�;=if1=f�y�N��-7��$
���9�Tb����Ƽ�HZ�������S��jT�n��*d�x��v��GzҾض�><�H>�߇>ZK�>w,?��?�%w>Ss.>� ?qP�>n�>�w�YC�:T��>���>$?��??S��>�b��K	�'N.���<��=���<~ٲ=1>n��=�ջQg���<�p�����kL=�%=��	���=�#0>��2>�xx<�wT>b1��P�MM�D��Y��>�Y5?<��<��f�<��!Ž�Ww����n_<W�r<�'���Q�����j�>�>vnc�9������=�\>o�,>x��=��=���������k>�-��j������Z�O�H�j=#T;>�@3<��#?wF?kX�>�ȽС��;��4���Бa���"���޽1�>�՘>a����5����G1���þ\�Ľh,d>h��=gV9>�0W>�5�3Cν��r<35�<-Y��N�>�;�=���=g��>p�>A��=	�+>��I>L������#���9<eХ��葼)y8>�wL�^R,�̲��w�'�������������>���=��N���?���Ǿ=u�������Ӵ�<�[j�'G��8Ǿr��.m4��⻽N��<X+پ�ϴ���c���;�V��9�x=�-��=��,�c���?�?ؽ�77>�
?_�9?��?=B�>��a�W,�>�\�>?X֟>�aT=X�=y1>*��>nc'?��?��>6��:1I�2�=�jX>a�>}Ro>I�>�^4��ڛ� %u<露<���<�5���3�N��'̮=+G�=���=�.�=��>�Uｏ.O��!F��~�ʾvJ>�3?����&��b`3�����ض�<�)�&,��^�۾s���ֹa>^��>���:��<�Lڽ��2��sֽ�3�!m�����qj����=��#=�� =v9��������M�u���q��`G>�X�=����*?r=?pK�>[����&��H���#�����(��Y >��ս ��E�6�D�U��,���%��M��*Z¾�,߼p��>�>x���O>�=qP�<Y�l>O�1>rx|�Dl>a����a>��>�*:>��=xP>�g��$S�i�����-�@�k։�Ռ�F�>�z�=l���jf�����>6Sžƹ��.]E���w=]0=|	�=a@�=p�=d
E>0ҽ:8�P�=&�=a���G���鈾V���>��E��������;�(��=��>�)Q��ҫ��{þ�k�>�)>�&�>��>FE?�b?u�>ͷ�<��>6I\>(]�>�H�>!��>�D?rڷ>�?�?]�= ����=�툾f���d�a=�� >��s>�Ę>��(�y�=�KR?>T=>6�2>t�=S{���^<�=H�>�9D>dq�>щ�>6o=>�F�V�T�r� �N��eoh>�y?�� �F�M>E+�e��A�?I��n���'��a���E>m
�>�	�>�z
=J�6�;;�-"=��>&��>6P�= \ݽ�6�<��=�b��LK�����Ǿ��L��G\=��6>���>���=:�?p�?6??u<h��Ⱦ(0�jJ9�R�� ���v>��@�Ѥ>w�>���<﷾���7�� .ʾI�0�9��>Q�>n��<� �=7�(�՝�����=�\�>�V�<H�@>�0>�T�>p��=f�>��>%<>�F�e2m��jӿ�����;�H򛾈)���Bo=�8!=�
���r��	�=���<�>A�ս��>h�$>��=�ʻ�Ƈ<2��拧��+=���=��&�"�Ӿ���;���v��D���G���y�޾�;�=fz�������B�i����䭾ާ��w+�>��c>-��>�F�>`�(?�R?���=�"�=fh?8�Ḻ>�CM����>~��> �>��?�!?ʰ�=�B���4��\�T�.<H�u=�b�=��>�d�>I}�<�C:UQ:ܭ<=r�����{�v<���<j��<ݩ�=�u>���=nI$?_��� fG�`D�}�X��I��Ʋ>���>J��<ߧ�=�����.�bM�1ŉ�n=��.?�b?NI�>�q^>n��>KP>ea?�#9���e<&}�=�T�=Q�	�(���.�½�;��8%�:?ѽA��=ܽ�={M��9>���='rٽ���>��D?S��>�h;?���v!�1i(�� �\��>��ʾ
�>���>��>B����B�^	��J.����m�&�Aq�����<X��>��y=�=1�C���>�Î>F=�&>(*�>Sų>.XT>�u�=kj>�{M>!I���Y��쇽p�ܿ�f�@�ӕ.��#>b{> ~��Uȱ�B�Z��s��Q��jɾ�1�=~^ؾ�����������%��SM={&X���<�Խ������ؽU��8:վ��9���fW����� K��
����2��(}��r�)��F�d;ͽ�y7��|
>4wF>�?��=��3?o�?υ?ʐg���$�x�>Zf�>)��>���>�?(Y�>�o�<]
>�W>c�ܽg����d�hw<�e<��Ȼ=�E>m�q=0;���J�=,e�=�
-=�h��ߺ!�t=�g��\=���w=��=l�
>'N�>�'վ���k���X"��-	������>�?�D��=m��~�:�p�
��\���n��w?�}%?�j1?d3q>Z�>�Zt=��=B���}��;�G�@��<CZ>�>2�����xQ=����4�`;$�+�!>lq�=9G=�w�=�E>�8�>��>�?5lu?�5���S�뾽�Y�O�F ��[?j�?�dS�pq����$���ھH����ܾ��}>9νQ$�>)����=���>]��=�O>��=2U�=�8���d%>�i�>���>�l>�p&>$9�=,J��X�=I�@K�z���`<�/���0�>TR=������{���`=?������[q���p��A��d������?w#�����a4˾��C���z��H�("��V�S�ܾ����A������Ţ�Nj���觾�{i��o����M��N������P���M>�
?-�>4�ʾl�?}�H?j�N?] R>���>�X�>��>#��>T�?�AG?��?\az��2�eYx�1�t��¨�W_:��:�=����ֈO=� >G�.=�a!���'�>df
����3m�C��6/���3�7=t��=L�Q=�?OW���mX�M1�S�W�b'���A �2d'?�����?B>����Q��� ���ɶ���>���>W%?#��>��>�3p=��L>)���e���(�==>q�>d`�����.7ܽn�Q��W̽캚���a>[>մ>��&=��U�ھ�=)�'?�8�>�?2��/0���4�B���;��=0 ľ�h>�>��r��v��ѣ۾k������&�J�ھ����I�T>��ἰ�f=��z>;0�[�d��Β�R�x=��>�BD5=Sv��ګ>	=��<Xх�+��7�b=�{�<Z��c��۠��P1��`O���νOV�<�<p=Py!=^
�=1"/�id�)�3���c�ݡ�=d��="=>��=��> ��H����9D�-� ����,��J�ݾX~�w�<�޵�׍�����=�m��E+p�5�����m��Ft�n����9�ҷN>�W>.}�>�V�>�8?;_	?�?X;����*=��>|�O�.��>��?X�
?�a?n�=�E=���=P���:��S�����ː=��P�q�>ܐ�>旄��o>t�)>��s=�2<�����<>V���(<�ǽ=<�.=��=>��?����s4*���!�]�"�~���h;��>,0��Ʋ;<� ��9����7��Ѥ<��
?3�?��>��~>��5>�C�=`]g=:2�����R�n=�y
=9��=E<�;��� >K弘H�8��<� >,R�</��=��>��ҽ���=l�(?"/�>JOq?%�1�'� v%� [�v�>�������>�͌>ť >��۽p�ϾP`$�IV>�G���`����1�%x=�G�=�'!=�>�g��D�=EdR>'T0=�$��TF�>���=�:�>���>�V:>��=
3���E0��ڼ�ڿ�鍿gR%�~���=_>*�v>�UN�+P��o�$��짼þ\�,�½��-�q�ȿR�����9н�ڂ�����NŽ��>ϝ��K�<����*���Už�߉�K�}�lP���Gľ�4�z¾�����V�,q����� B�� ;��M��;��I>���>l��<�q$?��?�?�j���>�Z�>d��>4I&?ð0?(�?���>���;�f1=�7*>�(�>�y��YZ�������U<i��;�a^>0�$=��'�Y��=e��=�29�t��<���=��ݽa6����j=��=�c�==�y>nI$?_��� fG�`D�}�X��I��Ʋ>���>J��<ߧ�=�����.�bM�1ŉ�n=��.?�b?NI�>�q^>n��>KP>ea?�#9���e<&}�=�T�=Q�	�(���.�½�;��8%�:?ѽA��=ܽ�={M��9>���='rٽ���>��D?S��>�h;?���v!�1i(�� �\��>��ʾ
�>���>��>B����B�^	��J.����m�&�Aq�����<X��>��y=�=1�C���>�Î>F=�&>(*�>Sų>.XT>�u�=kj>�{M>!I���Y��쇽p�ܿ�f�@�ӕ.��#>b{> ~��Uȱ�B�Z��s��Q��jɾ�1�=~^ؾ�����������%��SM={&X���<�Խ������ؽU��8:վ��9���fW����� K��
����2��(}��r�)��F�d;ͽ�y7��|
>4wF>�?��=��3?o�?υ?ʐg���$�x�>Zf�>)��>���>�?(Y�>�o�<]
>�W>c�ܽg����d�hw<�e<��Ȼ=�E>m�q=0;���J�=,e�=�
-=�h��ߺ!�t=�g��\=���w=��=l�
>�� ?0��06�i�辽���R�����>��?������=0�>8n���FCܾG����0>��	?��"?�&�>���>L�!>�_��H�1��d�<t� >���=���>��=`D>N�.=�6Q��J��RW>�Y�=��=�t>�:�=�ὃ��=�u?�[?��V?lyW����Wx���dþ�.�=��=l��=H��>�}I>��H�۾*�9������;E�>�_����>7�y>
�b=,M�=�#|�,���;�BY>��I��D���,�=�i�>�0
>��K>K�=�� ��X�μ ���޿2T�������u�����+��~0*�^{����A8���̾�����;�=;{>�Gs�=2�W;�<{�6
��m>d�;��`�O("=ˍ��h$���u��!V����4u�I-��'P��
�K��5ƾ�����a���T��>p��#�Η=^�>��%?'|ý�𙽔zU?��?������=�n�>p]��=�L�Lo�>���>a�?���>a��>A �M�ɾ���wq��1x�0�>�7A>߶=�V=���=C���	� �!��<�n�=�=��	�j0� ��Y��*��=�4>v%>.!?Y"���Q�����ľ�BT=Ŀ�=�F�>��X��D>`?�"���R�ý�1=O~U>�.�>�?�>ke^>b!�>��=+����L�������=(N��Dl>?�8>jp�=��<�w������T=���=4�>��R=ps=�j��^+�=�?x�5?�$A?���� ��D����.�>ԥ��+>��\�i-�>�vY=R����<��8��BU��&��<�C2��!R>��>ٽ<��J�>K�r�8_ѽ]R�=��M`���=�>^|}>��>�ÿ=�"�����4�E��Š���ݿZ���\6�:�/�V���&9ɾ��Ⱦ��P�yd�=����-�?����	뽗���Q�����=�Y���X�<���><��>�F����=���jy��:8�{%\�|l����:�ʊS����E�<���r���n��h��/I���C��D<r�p>�*7?��q����>�A?���>�`}>5JL��->�x��My�>�&�>�`?���>:�>
>N�+ێ���X��ww��F>n�p>Q�=bI;�-J(>;����\=v��=V8<�o�=�������7���a#�=�t>e
�>��?t���WS�5uʾD�޾_�">o�>�;�>�������s��J�ξ����;�{=��>�Ӏ>�E ?��>q��>��=6��	�y�;$�=�M>'(�<�s�>����*<_��=x<�Nk=��>ޘ�=[<�'X�������0��$=ˌX?���>��0?��>󣤾�D��b��k�����C��i>ɲ�>-�=��h�g����3۾�d��y�9�>v��1��$�=I��>�-]>q)�=e��<�#��Wf�W��>1nL�k"��u�R�rM�=d<o=�z6=�	>ü>����� �=mX俐�����`�=��`dh�����ԕ ��M�������=������<�X5����#�=D#
=�����޽귋=*������܈=����͐�����_��ƉA�-��c<��+������Z���2���,����YL��'�$������A�=��>���:�ޟ>+��>��>kđ�~��*�?Ne�=��9>Tq>�(e>Ö>��=v��<
L����#�yK���;�1>��T>����߽�:>�ž��E�:8��=��=R<q=4����]�K���(����H>mSc>j9>uk�>��ھ�����ݾd�ԾC'>��>��!>'��=Н>A�^�aY����ؽ(�(�F�=��=��d>�|�>�p�>Vӡ>9��<Cƾ�N��>��>��(=X��>�d�=�d�=P�>����k�=���=�׭=Bػ�94�y�/�#�0�߼Y?²)>��M?ҕ>�� �d<�_��'�����W��[�>?��>��N=�Rv�2j���0ƾu
��@�K��������>�V�>��z= �=jo��µ
��a�F�\>��Ž����f�=!��<�!0=N��=l@�=�i>q��(�W=9�˿�8p����;����Z�"���1�U�վ&o:�Y|���y��S`��DJ�SSf=���d��"�N=�U =�8�>�@��S��#��>�ӽ�C��f?��>����餾�}��ϩ�����z�ƽq���7���[=h���������<	�ԼT��=���>��e�i?>Bi�>��>>+F�=�4>�H>����b>��5>�B>&X>07>o>��<>M�J�������;�C>J�+>�!=/N��Z�<�މ� ;��$����� >E=!��<-���&���/8��0>�i�=2�Ƽ��?��P��+L��򾁽J�_=2>��>��>F�=(�>�����sd�Զ���(L=ȸ��=^��>���>N�>����𵟾�P���=�k&>�W�:�x`>�k$=}�=��^>ˠ���kN=f��=��">��=y����d��[IͽAl�=�M�?KWv>�ex?1z�>�=���Z,�_W�(��9䄾 ��>��?�5f>v�^��ھ=t��8
�3}=�d�0��r�7P:>�e>ch)>b��=�����ʚ��&��&>neӼ����Y*=e�;�-�=���=?s]=���==�2��Q���ӿ.���i���?k�;S6��V۾���Y쾜�ٽ�r�
|F����>҉��,f��h�<|a�=��<�6���$�O�����s�9c==�Q �"�y�(�O��`+����Ē[�rP�h�������"$�ʌ�	��T:ڽ[`н�?���큽4�>~��>Yc5>Ƨ�=ق*=���>滸>�	�=�i�>���^d����+����<D�[>���>6{Y>T��>?�k>E��X&�����=bw�>�O�>�{{����)>����>$��;������@6>�Z=k8����I���U��=@a>^�l>�G�>�c>#�Ⱦ�p�\g>�CܾN��)�;?z��R��=@u�=�<�A���pD� F��6>�X>J��><���F�j>yu�c�d�R�:�7㽆L�>�jC> �5>Dc�v\^>e��h�m=P+e>��i]�����07=s��M*>��/>C�?��Z?i�K?�+==������(���%��Ӫ�q�#��|��xޥ�#"=e	;�<�Pc��ӊ�"�����>:d=���>���=��=۪�=�v;�M۾(X�q0>_Ƥ�j�>ز��Z󆾃�>�E�>}�>�R>�`N>������@�ƿD���݋��8���g��d�=�-d�!꼓=Й��qi��A��<��>�Vg�h�1�>;LD>��/>ڍ��}۞=9�+>�d=�B�7�ˑ�`���xo&���Q���)�Ϥ;�Ž'`%��wO�����]1�Z�#�[�&�kD�>�_n>J=Ds2>Ͻ!?'L"?Qn�>q��|�">S�ռJL>/�Q>��>��~��>6l�=[�����H=�6e�D�_�r�=z�j=pOf=$
>L�>p� <�#>�l=	:{=k{���=� =CO�fW�"�ͽ��=�-N<s3�<ٿ<7���ƃ���j�*'�Xh-��d?ZԾ5��>jD`=�<� @����������=(��>|"?�F����>|ϧ>wo<U�m�	Ŧ���޽4<=� �=	��<�:F>�!^����=Lh�>}�s|	>�^>U�Y�Z׽��j�`�=��?3A?��N?�td=�:�N�"�כ���&�%B�٧��\>㽎yC���!>���<��c�m���v�/>�/=z�>d"�� ��OP>�M�����rK<��I�ڑ >m��=[�=�=���=!g>o,�=�F�:?ֽ�ܿ�C��α�Y��N�8�=@-�=͵�=)�f����Bw�����9�ǽ_�m���+���:g�=���=fi*>���
ݾ1h��M\+�(tԾ��A�����0�,�m��Z	�+�Q�����w��:�K�>�x���d��??��"�����>zV�;~b��� �=��?͑
?��>f��V�>j�|=W�= �>��>�n>�$�>����Yn�,V���|)>w��F�����=��
>�xz=ITu>�5�=q�=���=�f�<1^}<�Yٽ��<�L��=D���,��B%��&V=O��=s3�<ٿ<7���ƃ���j�*'�Xh-��d?ZԾ5��>jD`=�<� @����������=(��>|"?�F����>|ϧ>wo<U�m�	Ŧ���޽4<=� �=	��<�:F>�!^����=Lh�>}�s|	>�^>U�Y�Z׽��j�`�=��?3A?��N?�td=�:�N�"�כ���&�%B�٧��\>㽎yC���!>���<��c�m���v�/>�/=z�>d"�� ��OP>�M�����rK<��I�ڑ >m��=[�=�=���=!g>o,�=�F�:?ֽ�ܿ�C��α�Y��N�8�=@-�=͵�=)�f����Bw�����9�ǽ_�m���+���:g�=���=fi*>���
ݾ1h��M\+�(tԾ��A�����0�,�m��Z	�+�Q�����w��:�K�>�x���d��??��"�����>zV�;~b��� �=��?͑
?��>f��V�>j�|=W�= �>��>�n>�$�>����Yn�,V���|)>w��F�����=��
>�xz=ITu>�5�=q�=���=�f�<1^}<�Yٽ��<�L��=D���,��B%��&V=O��=�G�>�c>#�Ⱦ�p�\g>�CܾN��)�;?z��R��=@u�=�<�A���pD� F��6>�X>J��><���F�j>yu�c�d�R�:�7㽆L�>�jC> �5>Dc�v\^>e��h�m=P+e>��i]�����07=s��M*>��/>C�?��Z?i�K?�+==������(���%��Ӫ�q�#��|��xޥ�#"=e	;�<�Pc��ӊ�"�����>:d=���>���=��=۪�=�v;�M۾(X�q0>_Ƥ�j�>ز��Z󆾃�>�E�>}�>�R>�`N>������@�ƿD���݋��8���g��d�=�-d�!꼓=Й��qi��A��<��>�Vg�h�1�>;LD>��/>ڍ��}۞=9�+>�d=�B�7�ˑ�`���xo&���Q���)�Ϥ;�Ž'`%��wO�����]1�Z�#�[�&�kD�>�_n>J=Ds2>Ͻ!?'L"?Qn�>q��|�">S�ռJL>/�Q>��>��~��>6l�=[�����H=�6e�D�_�r�=z�j=pOf=$
>L�>p� <�#>�l=	:{=k{���=� =CO�fW�"�ͽ��=�-N<s3�<ٿ<7���ƃ���j�*'�Xh-��d?ZԾ5��>jD`=�<� @����������=(��>|"?�F����>|ϧ>wo<U�m�	Ŧ���޽4<=� �=	��<�:F>�!^����=Lh�>}�s|	>�^>U�Y�Z׽��j�`�=��?3A?��N?�td=�:�N�"�כ���&�%B�٧��\>㽎yC���!>���<��c�m���v�/>�/=z�>d"�� ��OP>�M�����rK<��I�ڑ >m��=[�=�=���=!g>o,�=�F�:?ֽ�ܿ�C��α�Y��N�8�=@-�=͵�=)�f����Bw�����9�ǽ_�m���+���:g�=���=fi*>���
ݾ1h��M\+�(tԾ��A�����0�,�m��Z	�+�Q�����w��:�K�>�x���d��??��"�����>zV�;~b��� �=��?͑
?��>f��V�>j�|=W�= �>��>�n>�$�>����Yn�,V���|)>w��F�����=��
>�xz=ITu>�5�=q�=���=�f�<1^}<�Yٽ��<�L��=D���,��B%��&V=O��=H碾 /̾�	)����a�ྟ�	��!>��=G�f�T>�j���F��ܤ>r�>	i��f�����>���>�x�����>�2�>��-�=��>�W"�n�C��M{�TQнJ�)>sɪ��$=��F��V&<:r�<��U��&>YMJ>EJ�a��>�?F��>�[?vQ|�e����)�'嬽n\��]���a�ӽi�>�i
��a�����=������A��վe8�=�:�>�I�=���I�=[�߼s�ѽ�>;�1>��%�\H��>Qu�<�)>�!�>��u> �=�m��'-���ο9Q��*���1�1�(@�����=N���Aj��[�a�ן�<6�$=��-=I� >o2"������c>>���> EX<� i��� �_��<&����H��θ������"�à��'�����U=F2*=p�H�'I���ud���R���d�~������>��\>��>��a>P�>�d�>�>1��Y ?�r>�w�=�+���.����?�>�O�>
�>Y>�/�>?�#���*����>���=&�=��v>s J>��=�,@=�:=��=l�,�����N����%�������70<�tp>Y�>����r밽��%�
�|�"�8�"��?��V=�f:�@�H>�H�ss��y�����<X�>�崽n[ >�Y�=ѭ�>ނ�>�#�=y�W�i�j-���pNy����(�>`�>�Pf=3�=��2=4��n(^=��K9ohG=��
�1>�5?�?r�2?�~c�74�5i"�T��.+�,mm�R�>��>���>-ZG�Uܒ��`�*� V�_k<�`��=�Q>�b��8�����|>1u�=��T>0�>�ʽB|�����}G>�'�=l�>��_=�/>�������&Lڿ3���l�O���R��q��.���nZ=�>��M�K=�>��ؾ�ľ�޾��)��ɇ��|�����׆>ɳ�>�ž3�k��� ��$ɽ�6B�sm�DsV��e��SA��3�<�$�_��Dֈ�����ҒܽF�:�͡���d�Q��S�?���>�s�=��V�n�<?�o%?'??�>�� ?R���I�_��k����=��>U��>�o>�Q?Lb�>4�>F`ؽ�҅�pw=s�=��h;H#>�a�>�0�<�尿�:��N�罡��=��2�q(�7�=h1�<1��<��<>�>��=\�K�ʾ���|/0��t뾰=�>�PK>/�P�u��>��о֤��;��������[�˥!�u�c��1�č�=>�>��>I�<=��
�2��� +��m>(��>u/�����!���Ѷ=�'�=�U>�O3����a�=6[���k�\�>�~�>�rb?�3?����ݾ�m����O��R�ܽ:��>��=�t��>�~>���@E�.<�8s2��y;���=9h>�H<Pȷ>m('>�G�Z3�?8��h����<�>kC?=��?>�>N�>�m>���=X��d̾@Aֿ	|��}�C���p�P����]9>�:�>�8���Z���Z>���`�=�I�UE>˖�>�<>�M�>�>?ϼm�����Ǿ�w"����
���#�ͽ{�ཚ�;��;�]cN��E��~�~��W����������=5UM�_?��S���-!?g?/r_=�4�>v
H??��>�B��-��>>�?^��d>�=�q=!ӽϜ�>��?��>�S	?��z>:'�w�ٽFOj=PL˽�:>�=f>�9@=U�;=�8>��=}��=�T���콻���v��{����=��K>Tb�>H碾 /̾�	)����a�ྟ�	��!>��=G�f�T>�j���F��ܤ>r�>	i��f�����>���>�x�����>�2�>��-�=��>�W"�n�C��M{�TQнJ�)>sɪ��$=��F��V&<:r�<��U��&>YMJ>EJ�a��>�?F��>�[?vQ|�e����)�'嬽n\��]���a�ӽi�>�i
��a�����=������A��վe8�=�:�>�I�=���I�=[�߼s�ѽ�>;�1>��%�\H��>Qu�<�)>�!�>��u> �=�m��'-���ο9Q��*���1�1�(@�����=N���Aj��[�a�ן�<6�$=��-=I� >o2"������c>>���> EX<� i��� �_��<&����H��θ������"�à��'�����U=F2*=p�H�'I���ud���R���d�~������>��\>��>��a>P�>�d�>�>1��Y ?�r>�w�=�+���.����?�>�O�>
�>Y>�/�>?�#���*����>���=&�=��v>s J>��=�,@=�:=��=l�,�����N����%�������70<�tp>Y�>����r밽��%�
�|�"�8�"��?��V=�f:�@�H>�H�ss��y�����<X�>�崽n[ >�Y�=ѭ�>ނ�>�#�=y�W�i�j-���pNy����(�>`�>�Pf=3�=��2=4��n(^=��K9ohG=��
�1>�5?�?r�2?�~c�74�5i"�T��.+�,mm�R�>��>���>-ZG�Uܒ��`�*� V�_k<�`��=�Q>�b��8�����|>1u�=��T>0�>�ʽB|�����}G>�'�=l�>��_=�/>�������&Lڿ3���l�O���R��q��.���nZ=�>��M�K=�>��ؾ�ľ�޾��)��ɇ��|�����׆>ɳ�>�ž3�k��� ��$ɽ�6B�sm�DsV��e��SA��3�<�$�_��Dֈ�����ҒܽF�:�͡���d�Q��S�?���>�s�=��V�n�<?�o%?'??�>�� ?R���I�_��k����=��>U��>�o>�Q?Lb�>4�>F`ؽ�҅�pw=s�=��h;H#>�a�>�0�<�尿�:��N�罡��=��2�q(�7�=h1�<1��<��<>�>X
�>�����'��().�+Ͼ���<s�>��}=�v����=�����UM=R$*�`��`��t��<�f�>0|�>�4>���>��W=�^��:�>���Y������=���>�p,�y�&>�ۄ=��Q<U�=�p�;�'����Ź7E+>\/|=�.�=H�r>Y�>?/��>�?�;�J�����{�=��о��ݼYC>䀘=���>�]�>>����M05����cͽ���� @u=#�B>��3>D�>D�l=Ö��Lt=0�;���,��A����m>�p>�F�>��>")˽��|��6�^�����O����оk�(�X`7��욾݌����C�9={.�����J)]=�#k>��*>���<C��;z~�=��ڼ�|�a*���9���
�	���^����u���y���ф���)��x��"�"��d+����/u��vN�|�х)>��-> i�>b��>��)?$�?ŭu>������?�2����=d��b�>��>�u�>�>��.>�8������?�����j(>��_�|>ĉo=�p�='m��s2�>����~�=LT$>���·-�L�ӽXi=h��9�d�>�=��?����������U�%WQ>1��>y�>d���y>>m�<�j�EM2���#��\���>Ӡ�>	�/?+�u>q�>'�>����t{=5~��w�����=�Z�=��<�=�=F��=ơ6=��C;7-��{�C �<���=��,>���>6�>��O?P�?5&?����J�����h�[���S>��=��Y>��=�Ǟ>�ͽٲ��"��o��B��i���=s#�=��Z=	$>�d���`�<�iP��VV=��^�����M<�޽�<>.+~>U�o>m��=�t񽃮��~������9;��� ��=/���=��ҽ�����&�Q��똾����4�J��=�-�>�"k>�-�����=?��=D�;�c5���O�����.<�wE ��^������l��ڱS�������_�o�u=��ƽu������V콬�%�𾃾e��RxY>"}�>W5�>}??y2?2�q>�y�>��<��><�ֽ�A>�=�p�>`�?F@�>pr�>0Q>�s��m���%2�� ��!�>/Ŵ�~��>���=x��=>F����>dY�;�S��-ju��b��G��v)<A"����J=p�b>W�>*?���z����a>8��e��6��>��>N�;�Z=*ȇ�L$��<rC��D?�r�G�=Y�>eD,?8:�=/V�>�~n>������=���(����<>�>y[�<�%G>��A>z�b=��=E|B=�be��mԽ�P��n��<E��>0˶>U?���>7~*?�D���ľ��FL�=o��CB�>��H>�a7��^�>���>��_��y��{C���P�N��=�����<~d5>��=�2>I�<�mJ�,*˽��޹g~����,�q�|�;>�6>��	?���>좑=a��	{�֪ۿ>Ϊ��g�A�վ7s>o�=�� �U��{���,��e��d+>��ջK�0=�>�����W<`�<�Q޽~^��i�\�=��N�I8��# =�зj�)ce<�L���䔽�`A��-ϽR9���J�V����2��b8���N�+>�J�>��>/~�>g�_?��>�޼�}�<��$?�����~�>C�>�?P1	?�"?�\�>9܁<�B���n�b(G�8�=�yx�^G>���="��=4>��)�(>j�L=�*��hx^=
��g��pg��4���=b��>���=f�?/�Ӿ< 径0侌��� 0>8Z�>��>��,>bj?*��<p�!�7�^���j>8�>�?L�>j;�>�>8�>�v�SD�=�F��]>�&;�9�>��>��A>� H>���=�J��Q�ݻ��&���<��=��>s��=�{�='�<?��?\��>b�q� u��� ��������!p��S�c>�=��>�]�<��ؾ�H4��gA��v����=�'>�r>�ܭ=!>e>�$Ͻ���'�˔�=�*=T�W=e�T<���=�y7>
�x>c0>w�<婙�!��B�Vņ��ƾ�)-�K��{3y�-S���M��2� �q��.T1��g�>�B�=uL>������<X��z����7�豜�-Yν���VJ������ж����|�\�\Ъ�9�{����@V��dR���	������6V�̓��$�=��y>�c�>�>%�?!D-?|A:>B))>��>�,o>�f�l�>�]m>i�>�>�?->6��=�=�>Jaƽ�&G���@�u�>�>=d>��Q=c�+>�	��!��'��Gg��ɬf�r5|=��%Rh���������r�=R�e>0�>�b��:�&�=v(��0�x�x�,j�>6$>?@�<�u?�x�s#�^�3�;%ؾ���>^�^>�>v!�>9��>�)�>p_>�ま
-�=�F�D���wܭ=�I�==g2>��&>	Գ=I#����<_j�9�޽%���-k��o��= �J>@1>�LU?<7?5�"?�d�@������Ѿ0����t���>��=a�>�K�ҹ�F-���K�ǜ�ϼ��P�<�ƽ��$>I�g=ڝ�>*�>G򽽆I>]~�8^��E�==�@=���=���>n��>k��>��>C#��S߾P�󿯜������&���!<7�\���-�M/��Ru���+�KC��=ƽ�j�<@[�=e��<Y
Q=��=͏�7e
�����}XO<��������־-ݺ��0Ƚ�5��]m���E��G����a�����A���b���[�j��w��.>t�i=��>���>��??��"?h�)<���>�'g>-L��s.�>$b?I�?�?���=�W>�H�>��|=�Ed�=9�����>�l�=�HH>���=���=���,���$R��N �z�=:�;����ʈ ��ꓼ�m=��q=}�>,?�������_������?>��p>�?�4׾^�?�ߖ��'�\�����@N���E�>R�>�	�>��o>�O�>��>v����{)�[�q���=��>h ��v;>\;�=���='~��������r>�ᙼ�Ro>�-u>����FP�c�}��()?���>�?C�1<P42��c)��#��#�S�򽾿?�=��^>Jq�~۽�����r��������������A�d���1n>�k>�ݽ���.�ν��J>��E���x��<>�Y>�\�>ŗ�<
�.<�o(�
4����t���=�5ܿ�|����\���gK�����>�/�[B�v��a���]�ӽ�y�<�W=M7=�|=�Ԕ=��=+x-�B+=��>g��7���C��x ��<��� �ýG��$X���vG��̧�lꎾ�A���(p�?�콊M���w�o��>�Y�>_=�=�+?a
�>̷>�ZϾ�?S����c�>���>�+�>�S0??�$>�[�v*o�E|��Ñ�OW��9=t0M=n}>�.v������B��J�>D�_��Ͻk"�=�ʣ���.��I	>zg;��ٻ=$0c>� �=�%$?9z�ӈ��z_��	��2=Í�>y.?�1���?�С=n�׾"���"��S�;��?�?��?�l�>6!�>t��=%E���N���=�����#>��>�>M��=��>��H=�n�o�<to�;�ü��=��=ܘ'��k�>�
@?PO?G�K?-��>���h
�UM~��A�ar��J>� ��4�����������������@���bdr��X>�O�>2.�=��=3A�=So�-��۽sj,���轏xC���?>(>�9�>�=�=-����Lӽn����Կ������~�D��������]��[��������VӾ����3�>Ug>�>���CW=D3�fOm��|Ծ�*�� ]:�}:���x�(?�;U���!�&���U�؅�CƝ��̍<��:�3ӽ�2	�/��k��ѽƲ��J#���J<� 8>�n?V��>�L>��T?��>�ߘ>�]پ�:?�����[�>Tv�>Ԃ�>O�?��,?���<�.6��wp=�5 �����y�"���#�-{��ى= �=�o=W�=�~;>g4����=��=���=�^�=�<=���<4��=�5�=e�>/�>*i뾛?�D�P�i^@�����7�˽3��>ILa�5��>���o���&��Ȝ������>��?�?�@�=�Y�>>�������
==$�$=��<ﹼ)z>� F=w=L�=^*�=#���f����&U=��R=t>`�]=�`=a_/?.�?8�*?�>m�b��Kݾ���d���P�->��=m��=�L���ѽ��-�,$(��L:�m�3��]⾼.5>_�5>��=��x=�܃;c�5�Q>ܰ9�rM#�3~���/>wW>�>l�4>��;�X��s�	�п=ɘ��e��F�?�
���]�<���Y���@2Ҿ�2��O����=��F=
�H=�	�=�==�K�<n��=���=5�>a�.>l(%���Z���R۽��->�E;UK���R�Q���˾�Y�9����I�a�0�l/�)�o�����}�>��>,�[�T'E?��)?v�>$
L����>�y��H�>�?�J�>�t?�3?�ń<�N����'�@g�v��w�۽�[�=�L����=��n=�P=5�8���<���=2Ă<}�=$>�H>��=H[ڽRh3�������D>�N?��ֽ�����w��A�/(4>_��={j?��ؾ��>i�@�j��F�U徲Q���\>�?�h?���>���>�K>�}B�C�4�u\=���=��=�=&\�=�
>*,>p��`7���s폽R�;Y�4>�5�<Hbe>[�3?�k?C2?禈>��v��>���>咽*�+���;T*�=�б���j�5?���	�h��S��]/���=�a�>� �>lC�=**�=;񕽴�h� ��=��$�����U�q}�>��\>�>�P�=G��<[E^��i7���ٿ=���qؾ���a+޾V˘���Ͻ8춾
f���ѫ���ݽ �\��=�`=��>t >����v?���矾O��쎾d�[��yĽ㓾��f�D����=�^�d'4<.���ㅾ����o��������%�O�����8n�	->ZR�>���>��>�(?���>Z0p>���f]�>�1��ߴ=���>�<?�?-3?�廇�d�V�~�p- ����w�����=���<�x�=~��=� �=ܱ2:��;X:Z�QK~=�� �
�*>鹛=��,>V�>��o=4�<r�=�N?��ֽ�����w��A�/(4>_��={j?��ؾ��>i�@�j��F�U徲Q���\>�?�h?���>���>�K>�}B�C�4�u\=���=��=�=&\�=�
>*,>p��`7���s폽R�;Y�4>�5�<Hbe>[�3?�k?C2?禈>��v��>���>咽*�+���;T*�=�б���j�5?���	�h��S��]/���=�a�>� �>lC�=**�=;񕽴�h� ��=��$�����U�q}�>��\>�>�P�=G��<[E^��i7���ٿ=���qؾ���a+޾V˘���Ͻ8춾
f���ѫ���ݽ �\��=�`=��>t >����v?���矾O��쎾d�[��yĽ㓾��f�D����=�^�d'4<.���ㅾ����o��������%�O�����8n�	->ZR�>���>��>�(?���>Z0p>���f]�>�1��ߴ=���>�<?�?-3?�廇�d�V�~�p- ����w�����=���<�x�=~��=� �=ܱ2:��;X:Z�QK~=�� �
�*>鹛=��,>V�>��o=4�<r�=�?�x�������d\Ľ�
M�.�=�H���w��yi �����)���ھt�=���>��>X��>���>�p�>[#>M:-���]>�T����=��>K7}=�Q���\�z5��&_>���hm��ʽ|����m=e�>�l >4 >��$?Y#?~�?��������������=���=�D�>�>��>a�a>�3���t<�����@߾o��Ao��0b=x>�˗���g>���=`>"�qe>�n>sV>-�R>=�c=b6�=�Ԁ>�F)>?�{���c��P���P.a���h��h���=�lz=��I=c�=�!>�*f>{Y�<�I>��>�2@>����먽5���t�<��<���P,�tZ0=�������������CU�]��T������V����o<?�h���k�O ��v�XC)��M��W�> 
�>wnM>�e�>)��>b(/?آ�>�Z�=8�>�n=�l>�V�>�\h>��+>���>���>�s=6�l=�Jx>8���N��,=7�k��ͼ~c�:�Z�<?�ǽ��c<�V�=
�s�o������<@%�<��<�Z=JR=F	>�*H>%X?Ia��0�E��^�eNн�X��Y���	=��`��!�����R>��ؠ��	>�X�>v{�>5��>�>{�|>�A�=`<��7��>�rs��/P=�`=t��=�� ��'�vU�=Sq��y���ԽP痽B޽�����>��G>cor>�3?Z'?��P?������IY ���4�T�[��񔾈��>�=տy�bUP��
���f�Bh���@��پoD�1��=,�*�/�ͽax>�S���9��0h>�R�>m;>�%h>)"G��[>_5�>i��=*jI>Hy�<�O��qy���޿�^���X�P- � �=�Y����<����-=���>1.�=��(>�^�>�={@>�~>!2=!����ý/[�\W�C3>]ķ����$�p�~Ծf�'�6��b�ŕR������l��t�8��@�-;'�1d�eN�0m�Nּ<S��>$�?V�\>���>�{<?�F?���>�n)?\�>���>�[�>*p%?��>�'>N=J�U�D&x>"DR�>{����ʥ����b3=�=��?>ԭ�><���<�{*��F=��N<݅~�Н�=��l=w=A����=o� ?��ϾKY�},��C��6(�=OC�=��>u�"�K��4��]!�]����F�9����א>[�6? �0?K�>ӆ�>a��<�!ܽ�q>x
��6q��;4�=�569�������h�=�o=q�ӽ�Z����>�潛R�=���=� 8>s9~=�?�?JR?���^���������[۔�hx?��=p���T >T���iJ��� �_k��9�%�Y�u܂=7�=�PO<x��>��i=�-<L�0>�<�=o�r>�$5>�O2=L��>�->�1�>�C>�=������ϕ��#��𻚿�vO�������I���.�k�ks���o�8��#YK��0׽�z�=���>L�H>��7>/TA=N_>�]>b.����N<���=���{*�:����i����_왾\f��s��sf��B�~�����2�5������`��8(�h�>Ԅ�>��p=��E?f/?]]�>�mD>��F?�^?k��>H��>}�?�-?� ?�#�>Uޅ��ҟ��`�>N�ʽ�������_�����k�b=���=[��<��$>��0�����<�_���7�+ڟ=�셻��=:�=2p>�?�x�������d\Ľ�
M�.�=�H���w��yi �����)���ھt�=���>��>X��>���>�p�>[#>M:-���]>�T����=��>K7}=�Q���\�z5��&_>���hm��ʽ|����m=e�>�l >4 >��$?Y#?~�?��������������=���=�D�>�>��>a�a>�3���t<�����@߾o��Ao��0b=x>�˗���g>���=`>"�qe>�n>sV>-�R>=�c=b6�=�Ԁ>�F)>?�{���c��P���P.a���h��h���=�lz=��I=c�=�!>�*f>{Y�<�I>��>�2@>����먽5���t�<��<���P,�tZ0=�������������CU�]��T������V����o<?�h���k�O ��v�XC)��M��W�> 
�>wnM>�e�>)��>b(/?آ�>�Z�=8�>�n=�l>�V�>�\h>��+>���>���>�s=6�l=�Jx>8���N��,=7�k��ͼ~c�:�Z�<?�ǽ��c<�V�=
�s�o������<@%�<��<�Z=JR=F	>�*H>%X?Ia��0�E��^�eNн�X��Y���	=��`��!�����R>��ؠ��	>�X�>v{�>5��>�>{�|>�A�=`<��7��>�rs��/P=�`=t��=�� ��'�vU�=Sq��y���ԽP痽B޽�����>��G>cor>�3?Z'?��P?������IY ���4�T�[��񔾈��>�=տy�bUP��
���f�Bh���@��پoD�1��=,�*�/�ͽax>�S���9��0h>�R�>m;>�%h>)"G��[>_5�>i��=*jI>Hy�<�O��qy���޿�^���X�P- � �=�Y����<����-=���>1.�=��(>�^�>�={@>�~>!2=!����ý/[�\W�C3>]ķ����$�p�~Ծf�'�6��b�ŕR������l��t�8��@�-;'�1d�eN�0m�Nּ<S��>$�?V�\>���>�{<?�F?���>�n)?\�>���>�[�>*p%?��>�'>N=J�U�D&x>"DR�>{����ʥ����b3=�=��?>ԭ�><���<�{*��F=��N<݅~�Н�=��l=w=A����=���>����j��=��1���k=�so>={<�(���=��Ͻ�.�K(@���5�Q1��H�>m�>j�?z��>m�q>i)D>�D
����<��=��)�!�>j�,=74R=��u�4H:�;y�M��n��A:��r1>��B>���<���>��E?��>Z '?��z�=�����w��&!���I�=��̻�_�=���5�v�4�x���/��o���n�>`�>_��<���=�2>�����J|<�=%u=ǒ�������Y>]�>7�?d�>sW��|��{ܾp�t��泯��ߒ�(�ھ��hY�Y���s�[��|�;��=�nH���I>�j1>�Iv>�ް=������	�iG�H�m�4�]���=���j Ⱦq�^� �~���-��c���/���a�t��'.������i
�;���k�N������U+��-�>��>���>dw�>�8?`��>�>��>�-?�2�=2�<�r ?�P	?��?]�E?7r�9s�q�+W��@��-|7��;h�'�Q= Ő=�pe>���=��>h��U�ȻU�=j�0>�S=�]<A�3��B���z=Z3=��o>f�?>ߚh>�A¾*�6��1���6�`�)>���=�=�1��F�>�6>���T���7E�b���e>��{<�}>���>v9�>eȽ>��¾�BO�
�5<O��=ևx>�NI����rs��|Rc�Oiq<S�,�,�P>D�>�<����z���yo�&�����>�E?X�J?q�� ��s���;�O���z��m�x �0K<��g�]���y���ݘ�����\E�������>��=`IZ=f�=K޽ъ;�>'K>�m6>bQ�=o��=ǴQ=��$?~��=�=9�=��U�dUf����=�ɿݗ��R����ؾ�qb=�*�=gg���#k�P櫾;�	�PW	=m���~���0`���3G=�`Z=B��=c�<�7p�������Ԟ<<Ⱦ��!�ǻ3�V8Ծ��м��:����ꌾ�z۾���׾� &�ޖ"� q`�0�m��L�=0��>9�>(��>VK�>�?R�m�{3>,�{>&X�>�9�A̝��d�>���>/�?�}�>L��FZ�=!9��l=��>F�qg[��u>�A&>�C0>����8<n�)�^�;<�*A=��=��>e�����<��R̼I�6<��=�fC>�h�=?�H���D��r�����pr>���>��?F��h�{��h�>@V�^���'��������>*�>��"?��;>�>�'�=_���K8ʻ*;��*�>���=�Ї�sAu�WUs�P>Ľ�����F���E��� �@(>��2>�^<Q���̓>��0?c�>�@!?7��Hv����о�x:���-��p��f�=�{@=O)>��ý��0��ɀ�Ju���Y�=�ia=R�>�/���3��^W=�E'��G�<��<�9>�tH>ŋ�=���=tp�>)��>�SL>y)��nF���w�RL���ѿ���e������K��c����׽��+������=>�H5��e >u�<\�>��`>=�<j6�[u^;�L>�_u���d�.�R<�g��U��*g�*���>��d�3�D��A����󽊼e�Q�`������$����R�+=��>��>�l�>�)�>Q^F?L3>>!k�=߳�=�>y!:>U�����0=i�>H#?�0?��a�@8X=�Ѻ���ؾ�(�p����|>`>�-�=�s=&��=��=�G=�|¹=�y>�Ҭ=�䨻ɢ�:q=�6�=��=�Y�>pc�>���>7��~%��l辔.���>[,g=[��>�⿽K��>��>����P�۾��̾��ʽg$}>��>X2�>��>�;�>�h>���.*5�/=9Hd=$�<>DN>^�齊�ɼ+q#� ���rޒ��_�=���=�Q�=�`�=�0���D��R>u ?�?��/?�=����⪾;0�{b�$���Ϻ6=98�;6�(>�.����������I��tʺ;��D=��V>��=5�<�|��OR=u���2e�l:>��{>�<��>1�>�Q�>Oq�>�����t��zHf>�Cݿ�\��W��«��t6>$� >��k=8��<�v�K���A�_�����r۟=/)=X�P:���7Ɏ=¼��W��>�{�x�9>�>���ƾ��.�Jȿ����Ӗ�w%� <>�J�a�޾,��껾Q���:Qb��ڍ�l.T��5���f�>��?��>p� >%�?���=uۧ=��P<q��>�B��+�e�\a�>��>!�>���>}�c=Ly�=T����"�T�1��r��>";>*L>����-I<�x��ė�<������=[M;=��@�o�������_��<(�)>���>�O�����>a�q�N�״��rV���Q=c~0>Oat>[A�����>k�=����_�ξ�0=�y�>^o�>&� ?�3�>�;�>��O>h@��M~�;e�5=�1�<Z/�=�+�=q��GxW:���E�ƺ����l; �׺�4>��>i�v=����/o>�'	?��>(�5?	 �:����辋yƾ�=�~���܈=��v>�IC>J̢��m�U��ľ�ȩ��>��J=�c3>��=(�	=��\��8y=��<�7�s�;>�@��(kM>�x>�B^>�j>$�/>C~� C���j�3ղ=t�ڿq����1�A`���N�=s��;�e/>�H�=a]ľ�D��&§=L��<]�>E�_>�3�=�(�=?�%=m�>>\k=�/Ծ���!�^=&��T��k &��)j�,A�D Q����:A}�����`���c�e��}��k��;<�@�><���>�+?�>� �=�D?�*)>�t�=�Q�<�@�>���}�z����>�Ԉ>�Z?���><3�=!U;�촾��꾿%��_���=>�)=~�^>�鿼r6�i2�=�)�=]�%>X[<�1>�AA�����l˻ʗ�>;>��>MJ5<��><G��}��h�0��X������>՟?����}��=·�>^�e>��ľC�����~�����>B?m�>�ڧ>_'=�珽��2�
���w޹�s!>�62=G[�m�i<W�t;4a=���$/������">�ݓ>e��>�^��EKe>��?dS?�G?��<R��S�Q�J��p<6�ĽE;~��/>>�2�>	r�>��ݼFg0���E��&�Ѣ�G�Q�Mx>�b޽L�<�>1'7=��6�[�=~��=������=l�]<)V�>�_>RCg>��=�[
�5i�x��s��������=Y7q�э>��>,v4>���l����e���ξI�v���6�c����>���=�� �^��h-=����@�)�W܌��$߼�8��#p��"L��åK������½
3߽ ����t��k��0@b��ޭ�#��������۹���>�H�> �	=5��=u�%?��?�VK>ˑ���?��=�=�=�{��y >ib�>i�>�~1?%]�>e(>o6�cL��}
&�(t�>�:�;��>�Ґ>��F>��ýݝL<�AH>�@e�� ��`9=,��=���=1%+=�ʻ��*>j��>wg�>ߙ
��s�CH���Rc�����k�>O�>-	^��vs��I�>~��=��{�L�T�#��������>-�-?ȵ�>��H>��=>��4������=g`�;�E�=�'�=�O�o��=���=>ֹ���L�������~'.>7�=S3>�۩=�w�>��B?yw,?-�?R���w�Q	l�4O7�?�6>T ��fľya>�j�>e.>Wv)���= �d�V����T�o<�+>��=d��V��<<N�=�ê��h�=�կ=�v��<Ē>��=��>3, >"�>kR>i,�=�J��B[��F��ì���H;��'��H,=�S>ǝ�>�"/>mh*>��/>�!�L�������U��=!�=>^�+>(%�[�=�l�=�Ѳ���Q�nq
>��=O~��*x�H�q��������h=C�����E�� ��V�u�����)7)��8��ݽ���>���>��&>H->c�?��b?��>B>���>R";>��>�{<�Ys�>���>�`?i\?�>5 D>Y�=��O��RE>){�=urj>��<�z|>C_�=�=w<f꘽ĊS�&�>�<���<0�<�,�<z�	�7AB>��>�?�?�=_P�����XO��5վd�ɾ�l?��l���>��	4��we>�+�4�"�P�J�lB�2>w_�>�L?�	d>�58>��9�6ƽ%m�T�ٻ��I=�U����;�_�=�K��Yy:=��>����x#<�b~;��N=�+3�����0>2�Y?���>���>76ֽ�h'�=��x.��M���t�{�B>p�����U>ת0>�f��)�������2����wN��X >��">xș=i��<�k6>\>�����).>:=C��b>ͩ�����
&>�@�>��>xz�=�9�}���,ҿ�n���"�]���9�=4St�Qm�<������?>5��=��U촽Jz
>�=*�4�n.L���F=�W�<�d��W)��VJ=��T=c�����U��вC��U
�����:��
�K{���:��m��b�����2W�<����kV>a?�<���>K&!?,�R?Z<^?�~/?�?q�Ï�>k0]>`5�=BB��Z�>3��>@\?��?+�4>A��=�4���Vz4��<=�{�Ϥ>�=��b=�.>�YQ�+�=U������=i��<��]�������=���=�c>�"�>�>�=����;�Ss_���=�RK۾�V�]�L>3U�[�ݽ���=���LdI�u�=�V|:�|�L�Ӻ�="ߵ>���>~~�>7��>}g�;4�n='Ŗ�Y��&Ͻk�X�nM�V� >*@;ʑK�J�z��sƾ.l�/���U4=_S�� �=�J�>|�M?���>~��>��l=�����?���-�`0N���>�[�>Ô�>���=��5=�����|�
���D�;��k"��%>����e�<H�2>��6>�`�<�=�:<�	ཪ� >��7=��K>�|�=>ǥt>	G=t-�?�j���ٿTt��z�ʾ%�O��\[��r0>sL�>�u�>P�?Ŏf�j.��s�*��1S>�a�>��>�C>o��d^�=��0>�$�����@�;� Ž�W��x��S�Z�<�
%��xؽ"s�k,��~���0>�N��g��o(���E
�4+�#�>�2P>ש>;}&>�?vU?B� ?0K>V&>p}��x�T��ֹ�>@�>�/=?�T"?�&�>T �>��i>�m�S�r��s������=��;AAA=?��=B��=�9=r��Z�=o:�=�΋=��޽y�9�gO�=z9>r�>wg�>ߙ
��s�CH���Rc�����k�>O�>-	^��vs��I�>~��=��{�L�T�#��������>-�-?ȵ�>��H>��=>��4������=g`�;�E�=�'�=�O�o��=���=>ֹ���L�������~'.>7�=S3>�۩=�w�>��B?yw,?-�?R���w�Q	l�4O7�?�6>T ��fľya>�j�>e.>Wv)���= �d�V����T�o<�+>��=d��V��<<N�=�ê��h�=�կ=�v��<Ē>��=��>3, >"�>kR>i,�=�J��B[��F��ì���H;��'��H,=�S>ǝ�>�"/>mh*>��/>�!�L�������U��=!�=>^�+>(%�[�=�l�=�Ѳ���Q�nq
>��=O~��*x�H�q��������h=C�����E�� ��V�u�����)7)��8��ݽ���>���>��&>H->c�?��b?��>B>���>R";>��>�{<�Ys�>���>�`?i\?�>5 D>Y�=��O��RE>){�=urj>��<�z|>C_�=�=w<f꘽ĊS�&�>�<���<0�<�,�<z�	�7AB>��>?h���}G��,��.L��6)>*&�)�
? ���]μ�����������������i��R��>��>�C ?2��>���>�Z�%���+{���s�<��=���={�=p��43����<��$�:�ʔý�:���i>8W>X�->���bZ�<�d?Tp/?9�P?�s>b>��� ��`%��	�=�Y�>���>
��>"�=�&&�%<޾\P+��1�w�<�ՂѼhV�C�=��>s�2>��Q>�CϽ�%Ͻ�yo<��=4�y=[%>un�>��0>)�[>fV>l.6�q~���T���x���ؿ����h\���Ⱦ��<��Y;����~�	�E��P��p���g�,m�=^w,>J�=�=��"�!�j��!�F��q�轼�;��E�fξ�x��+��������\��[<�_8(�R��� ����̤�O��呾��s�x�<���=j ,>AH�>.�&>q�G?�?��)?X�=$ܑ>[H�Z(�=a�]>,�>�D�>A�?"t+>:��=�S<F7��]����ꪼU�^=#�{<,C�Ű�=�k>�2�]?�>mZ���22�<Po���=>o=��]<�>?�=a�o��=?h���}G��,��.L��6)>*&�)�
? ���]μ�����������������i��R��>��>�C ?2��>���>�Z�%���+{���s�<��=���={�=p��43����<��$�:�ʔý�:���i>8W>X�->���bZ�<�d?Tp/?9�P?�s>b>��� ��`%��	�=�Y�>���>
��>"�=�&&�%<޾\P+��1�w�<�ՂѼhV�C�=��>s�2>��Q>�CϽ�%Ͻ�yo<��=4�y=[%>un�>��0>)�[>fV>l.6�q~���T���x���ؿ����h\���Ⱦ��<��Y;����~�	�E��P��p���g�,m�=^w,>J�=�=��"�!�j��!�F��q�轼�;��E�fξ�x��+��������\��[<�_8(�R��� ����̤�O��呾��s�x�<���=j ,>AH�>.�&>q�G?�?��)?X�=$ܑ>[H�Z(�=a�]>,�>�D�>A�?"t+>:��=�S<F7��]����ꪼU�^=#�{<,C�Ű�=�k>�2�]?�>mZ���22�<Po���=>o=��]<�>?�=a�o��=?q��=^fV���h��f��	�=�2}�X�
>�k���ƾ�0��`���!�+b����8����>�<�>���>j��>�{>�=Ҭ/<r�ý�}�=I�=�D�6� >���=�[h<�������UE��S�����$=���=��4>4�t�n�h>nB?�!?�`S?�o��"�h�@)���O��ֶ�
��=g�>};=l�=��Ҿ�.��l���ý��xq!�+��"g�����=��ѻ&�<r62>_o�<>
�jY���Vp>Wg�=�V�<�I>�Z�>�Xt>^	�>3�= e����.�?ƽN��Ͽ�h�?4žHՃ=i��=�9�=�J>�"f���V��xپ��}��`�>^;�=O��=�b��ԣ���9=4M+�U��>J��>`�=��<�������"Ɔ�@�1��M־�]���櫽������I.K��榾��,�vY9���r�]���z�>��=�t�>�7d>�6?s�?��#?1��>��?xƹ>7��>s��>[�m>J?��E?��=���=���>�4��Жi�����[�w����<�	/��F�<�%{>�=�˖���x����<�#=��@��6�=���;����%	K<�g�=f�>� �>�Г�*�/���Q�)�0��V�QG>���>��Ǿ��N��6>���:�Q��`L�����>�D�> �&?�/�> s�>�T�="�ڽZ�7�'l»;6�<���= cu>߹��r ����=�@ǽ��{���C�%jG��=c�>R�6>x]��2R���/J?B{,?o�>?Dw_�u�9���۾�%�QW��W>�X�=�X�>~�m=1���y;���� �����\?���T��9r��|>��>a��=��>Y���3m%�	>@q�=\�:=����,�=�?4�n>N�>�Ȣ=����1fS��3���տ�%���cM�V`��X#h=�=@>��b��ѩ���=$�=��������v�P=T�d>z��>� �=񃚽`����*>����'X[�
���aBt�=J�����Y�ľ.o���Me��<���IFӽ%zȾ01�������J�*�e���E��Ū=#L�>�"�� �=<Kq>21?�?v�@>.pU>��??^��!@���>F��>��?�"?ݐ�="��=��/=Œ8��S��!fL�Q�>}͢=���m�>��S>�J|��;��<�!$�j�=�Q|��
>��?=M�d�;�=a��=~v>?h���}G��,��.L��6)>*&�)�
? ���]μ�����������������i��R��>��>�C ?2��>���>�Z�%���+{���s�<��=���={�=p��43����<��$�:�ʔý�:���i>8W>X�->���bZ�<�d?Tp/?9�P?�s>b>��� ��`%��	�=�Y�>���>
��>"�=�&&�%<޾\P+��1�w�<�ՂѼhV�C�=��>s�2>��Q>�CϽ�%Ͻ�yo<��=4�y=[%>un�>��0>)�[>fV>l.6�q~���T���x���ؿ����h\���Ⱦ��<��Y;����~�	�E��P��p���g�,m�=^w,>J�=�=��"�!�j��!�F��q�轼�;��E�fξ�x��+��������\��[<�_8(�R��� ����̤�O��呾��s�x�<���=j ,>AH�>.�&>q�G?�?��)?X�=$ܑ>[H�Z(�=a�]>,�>�D�>A�?"t+>:��=�S<F7��]����ꪼU�^=#�{<,C�Ű�=�k>�2�]?�>mZ���22�<Po���=>o=��]<�>?�=a�o��=��>�B�����(�g�D�n�>ZW�<(�>�x�=-U=Lg�O0��.�.>���N�ھ�p���'��V=�V��>zc�>��=�L�gh@<�>V�)>�=YD�= %���X���;������=EcǽƐ��0���%�=%�M> 9�>�)�=-(?c'?x��>�D����9꾓�;�}���Yg�*%��*�R�����ǽ�E���3��S����z���Ȅ<��>�>���ڟW��%ν�R��P�Ã_>�>�5>? L>�">=���>�*�>n
U>詔=����¾*�̿�钿4�׾$�_�>1���z�!��,+>�h��f�f�b���P�=*^(�S�F>DՌ>]��>jK>U�>/�o=�s�.���Ex��V%�Z��_]�T��8�5�(㝾��~��:��ff.�MB�xO���|��7ۓ��3	�3B��N9&��-?D�>�@�>��>s?�H�>dw�>��'=���>�d�>��?�a�>�d3>�`?p��>��>M�?�~>n���;�;��:��):=��
>e>;��<;�=�Z�=%>7�>44Q>/a�=d�o�������+>�+>:�>I"�>�-�=��=>6z4���$��*(����%��9�����>��\�Y>
�I�j�=�X>�Q[�N�&C/����Ph>-H?��r>p>�}#��w(<�]h=UR�=u-�=��=eЋ�"A���)=�:�=��=��=Vٞ�yb;��\>-�=6a���v�<�kb?:�b?�)>a%�6�?�
���JI�P`������#>پ��YH��>ž:��G���k�,׾^��<���=��	>��<|W���ʴ�G�Ͻ	w=�y>�ٮ=��>�d'=�(>,Ή>T�`>��>�M;�w�*��B?ܿ�=�����G|����3�Cc`�9���M)�#C��������	��������ƻ;]��fý�������=�P��Ǿ��3rؽ�q�=K����?����_���6�Z�W�
�����Ǯ���w���㜾�� x¾�z �R��5�սD�?�E=�.=�)?��F?�@?�7?��>ui?j	�<_)?/�>+$�>1�>?#7?
2?�>?]�>�ْ�+Q�R2��ͽ��:���=�d>ox>~^�=�z�<�̫=<{}<)��<a-�;�C�����=�Ϫ<4ֻ=�e\>��=��>�B�����(�g�D�n�>ZW�<(�>�x�=-U=Lg�O0��.�.>���N�ھ�p���'��V=�V��>zc�>��=�L�gh@<�>V�)>�=YD�= %���X���;������=EcǽƐ��0���%�=%�M> 9�>�)�=-(?c'?x��>�D����9꾓�;�}���Yg�*%��*�R�����ǽ�E���3��S����z���Ȅ<��>�>���ڟW��%ν�R��P�Ã_>�>�5>? L>�">=���>�*�>n
U>詔=����¾*�̿�钿4�׾$�_�>1���z�!��,+>�h��f�f�b���P�=*^(�S�F>DՌ>]��>jK>U�>/�o=�s�.���Ex��V%�Z��_]�T��8�5�(㝾��~��:��ff.�MB�xO���|��7ۓ��3	�3B��N9&��-?D�>�@�>��>s?�H�>dw�>��'=���>�d�>��?�a�>�d3>�`?p��>��>M�?�~>n���;�;��:��):=��
>e>;��<;�=�Z�=%>7�>44Q>/a�=d�o�������+>�+>:�>I"�>�-�=�k>���=����������lm)��û�*�>�gu���{>;�� �=���.1,�y�*�h��2x��
=t=J ?�D�>�y\��t���qd����=��U�ᘥ�X:+>��߽��=I�ԽlH�>�>��}���<�2��0��;ɧ�= Kr>��=�*<?��A?���>}W��g�/�`�W����mVH��AĽV�;���L��˾o徒��h�>�������-<�0>W�t>hRD>���
k`=�x�>l���_N>����6v=��<�rp>q��> S�r�:=(�����2�d���Ŀ,����2��߾1zd���ս��=ğ�>Cb�>�����I���8���?�=�^=�e�>�ב>)n�=���<-���!���ün���:���E���^�i=���W��뜾i*�%嘾�sn��ޣ��������3ꏼO��PӾ��~���?��;<�o>=���>��E?��8?��?l@>q��>��Խ7�3?�Տ>x><�)?�?_-?Tf9?��?"����J=v� �V<f�z,#��÷=yoh>]�,>��;�v�=��=	W>�:���9Ž*ټ�I>���<a�>�Pv>�B>�k>���=����������lm)��û�*�>�gu���{>;�� �=���.1,�y�*�h��2x��
=t=J ?�D�>�y\��t���qd����=��U�ᘥ�X:+>��߽��=I�ԽlH�>�>��}���<�2��0��;ɧ�= Kr>��=�*<?��A?���>}W��g�/�`�W����mVH��AĽV�;���L��˾o徒��h�>�������-<�0>W�t>hRD>���
k`=�x�>l���_N>����6v=��<�rp>q��> S�r�:=(�����2�d���Ŀ,����2��߾1zd���ս��=ğ�>Cb�>�����I���8���?�=�^=�e�>�ב>)n�=���<-���!���ün���:���E���^�i=���W��뜾i*�%嘾�sn��ޣ��������3ꏼO��PӾ��~���?��;<�o>=���>��E?��8?��?l@>q��>��Խ7�3?�Տ>x><�)?�?_-?Tf9?��?"����J=v� �V<f�z,#��÷=yoh>]�,>��;�v�=��=	W>�:���9Ž*ټ�I>���<a�>�Pv>�B>Ҋ?�"����"����'�1o��,�=�$�>@�t��@�<�7���z˾�=�,��>""\=G��>��>T6�>��>:x>an>����$͎�ͽoi=� �د�==W�>�Ȃ�V��=�t�>���";���������<R�����=�Rx=�u?.@<?sR?*���V�F��Y����Ob���=���=K\���"A��c��N.�?���M�=V�=�0>��=g�	>�J>Adk=.��=?j�<	��e�<��鼅yǽV>�?�=)P> M�>��'>3T=��@����sǫ�����1�����=�JI=�Y�;��l��.]��\f=�U��13-�3�<t?�=V �<�7����=g/v��&���⾻d���N��⡽��������q��~k:������!��L�K��`�½-`��� ��@���0��x��l�c>7	�>,b�=%Iv��L?�?(:i>�G>�=? ��p��>���>�� ?.��=G��>�u>�m���,�>��y�����D9�G�R>u~r;�	> Ā=�=r_ս������=
�=���C��=�=��=��l�����=�_�=`��>�������w��L}*� �����>_��>�����>�;�P2��B��%0��^��=$��>��>HͲ>d����>�g��[ �m����X��^���=� ��?4���Nf�	����$T�}k��S>D+->�Z>2>���=���\�=u{!?�N	?v,G?([5���j���m� �8�4��Ⱦ2�a=�N�=�ܾ=�T1�+Ծ��Yw۾��.��=��J<�$�>]�⽏Y1�-M�=�D�Pʋ��߼v͎>�Mw��P>�!�>sjD>s>����k�5=�����輎~���ɿdZ��u�)����������sf�=��L�CN����=��Y�� j�mJ\=������=�
�<������$�=9��б���>o�f�?�����-=���.>4�����=�\c�zs�vT��᥾dQ��wG���t�;긾8���ɹ;>���>-��=�͜�V�N?
�?�<%=2�-=��1?��j�c>=��>��>e�m>���>a������<�oO>��
�s�uAR���+>,�=L=���=NP>��= \Ҽ2$`>8'ջ^$�4	��l����=��ƽp��;٬�=)K'> ?��7����*�M�C�����:P>8��>Q��o��ҡ���Ѿ+m1�N(�&��">j>��>�W�U�W>:P�>5��=�	���!��R���z; �D\s>-��>
ZڼP�=�Rl>߲���i=�=��=02b>X�=�?y<�.�??'�?�A?!�j�^���뾕B�D�C��̝���;��F��y8>����ݾ��
��vܾ~ƾP(��E＄W�>��>'~L>�%�>)<��H=zp����W��L2\=E��T�=���=&��<5��N�����;|�=i��3��D}���Y���=���?s��%����U�t,�=��	�8���Z�^>�>E�=:��#��<���=�-<=���������z=~���ʗ��|����������z���ƽ&�@�A�>�]H��S��=m�! � �I�M�}������MX>���>��?�v>�D\?pE?�#\>�>,>i�0?�WO>i��>+�?�
?�%;>:0�>ǡ�=� ����g>��=PE�&\���)>X�=��<ԇ>�7�>��[�.Z4�+$>�o!<�νR?<ƅ��h�T񺼇Ɏ��->'��=#�?촾ae'�O�
���Ry�=O��>l�?v�V�X^>-�������h��yz>ب�=�3�>� �>}�^�b��>�>\�@>�x����
���>�u=!�n��=p`>���By%��|�= �b���=�{=�\�=�QZ>�>�v>b�;� ?�>��!?��L?���Ÿ�ڛ��𮾃�<��i>�ˠ::��s<���=:��ǐ�
�%���%��K����"Sq=F��=錪=$��u����!��i��=ѽ�=r�H>9�1=�֊�����<W>�q�=�=�O�;Ƙ������Yڽ�`޿.�~������)�7+��Lh��<�����ԾPWؾ��#�k�޾�J#�L�K<X�����=t��=�n=�)K>���< IǼN>`=�>-7�=�M�����zƾ�`���[�sV�=b��tV��z�����?F�Ϻ���ҽC����������>��>J}6>�q
>��??q?�\H>�[��J?�غ=�m>�j?GH�>E��>>�>����,>|��>��>	)M�������'>Q|�=���=G>�>M�H� ��/B�����=���=�s�=�
�B�ٽ3՜��k}=yi>���=#�?촾ae'�O�
���Ry�=O��>l�?v�V�X^>-�������h��yz>ب�=�3�>� �>}�^�b��>�>\�@>�x����
���>�u=!�n��=p`>���By%��|�= �b���=�{=�\�=�QZ>�>�v>b�;� ?�>��!?��L?���Ÿ�ڛ��𮾃�<��i>�ˠ::��s<���=:��ǐ�
�%���%��K����"Sq=F��=錪=$��u����!��i��=ѽ�=r�H>9�1=�֊�����<W>�q�=�=�O�;Ƙ������Yڽ�`޿.�~������)�7+��Lh��<�����ԾPWؾ��#�k�޾�J#�L�K<X�����=t��=�n=�)K>���< IǼN>`=�>-7�=�M�����zƾ�`���[�sV�=b��tV��z�����?F�Ϻ���ҽC����������>��>J}6>�q
>��??q?�\H>�[��J?�غ=�m>�j?GH�>E��>>�>����,>|��>��>	)M�������'>Q|�=���=G>�>M�H� ��/B�����=���=�s�=�
�B�ٽ3՜��k}=yi>���=
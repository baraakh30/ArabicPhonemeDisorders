�	  �   �gվ#��>���fK���N�Z�d��߻���=u�:���=&���⾴gV���n�R7(>;��������=��M�Z?u Y�𓓾˅�%���;>��C>���>°�=��,�cb��6O���<�f?>��d���ԝ4��,龦(�>�E?uGc?�L�?�a���i�H�J�}u	�
����>��P?��>O|?�:1>�J�=�ݦ������a��CF��m�>w3�>�j��M<����������*���m>�#?�iE>�?�S?eF	?)V?S�-?�~?�Ց>uޫ��:��w�&?�t�?�ʂ=zҽ��V��w8��zD����>߻(?�lA�P�>� ?�D?oo&?+^R?ý?�4	>�� ��?��s�>�>��W�OW��aw`>rK?y�>�Y?���?؜:>$�4�ZJ��g%�����=�>a�1?�Y#?�S?F��>g��>���#�A=��>�Z?Fy?�c?�t>x��>T>��>l�<яV>�}�>6&?
)C?�si?p�W?���>�<e�ֽ���?$���Ώ<hj��>�=�\>\!��Z�e�Hcٽ��컒Cμ�S��}�����f�`�l8O�绋�`=&��>��l>5���{�->�WȾ�9����H>k�ѻC&��"���ˬG���=�x>�K ?��>�B��5�=�^�>/ܼ>� ��*?)�?��?���<�Ud�)PѾ�l=�n��>O�A?< >�+m��Ր��aw�\%v=ʸn?��V?�JB����b?P�]?C`��<��ľ;�b��
�=�O?��
?x�G����>� ?��q?���>��d�{9n����Db��Wj�ğ�=�9�>p`�"�d��?�>��7?)�>�c>qw�=4�۾k�w��#��\�?%��?@��?�?x*>D�n���L�߾m�����_?�2�>�G��o93?$AF���ξ�}��ϭ�+5�b���0n��]W��Y���b.������_��F�=�?�4�?T�q?�c?�|�Al���W����C������9��/T�N:�J�v�]O�W��h����pY��J��c�?t�?���?�-��V)ھ�ƾ3��=�d���-���.>U�_���=�z=������������:?�c�>G�>�fD?�kR��P=��)�ΠK����:58>�f�>�؈>�o�>���<a�R�S+�ذ��)������;v>>Hc?�AL?m�n?-���)60������"���$��|��TB>m�>{�>1�W�.n�{.%��P>�~�r��-�%���	�	�Q�=��2?�;�>�0�>�0�?��?��BN��Us��h0�݃�<D��>��h?d�>{A�>��ν� ���>��u?���>8�>S眾7�5�nX��m�V>�)�>��>��&>[
#���\��K�� ˂��E9��6=��L?�5�8�]���b>�U?m�]���K=�k�>4|[�FSB��ѓ�[N�`�G>2�>�����H>F�վ�]@�r�t�����$&?�q?�����K,��Gu>+?R��>/�>U�?]7�>���N;��?%�_?y�E?��;?-�>��=����f���;.��+=@�>v�a>�E�=-��=�^����a�7��Ar	=�A�=�]&��⽭�;��A�?q�<��D=��G>�+ۿ��K�0�ھ�d��X��d
�
��S�������aq�Z޵�2���n�z�J���M%�}mU��a��;���Im���?ӕ�?}ܓ��_����%^��Y�>��n�/�����a���#��w$߾�'���� ���N��i�^�f���A?.�l��ƻ�ُ������ ?��(?E�W?W ��|�m{$��<�>\�	:o��<�h��6���H�ȿ�F����n?�h�>�*����Ž�h�>��~>9�z>�>%&z�Fn��6�?�?�.!?D��>��)��¿�ϻ�*��<�g�?	5@��@?'��r�`t=���>3n	?R�A>��2�Ϥ����x]�>{]�?޷�?9u=C�W�5Iܼ_�d?�+<�G������={�=}�=s�^�H>���>���$FC��sٽb�;>���>֠����P�]��T�<��W>�x���Y���҄?>p\��f��/��O���)>@�T?=�>�.�=ì,?�5H��wϿ0�\��%a?�$�?���?��(?Fܿ�˚>�ܾ>�M?�=6?6�>(o&�H�t�hN�=���)�������V���=���>n�>�R,�?��F�O����� -�=����e{ɿ��?�&.��頽N�����&���
f�`>ᅼ�/�Ⱦ�q��S���]X>�>��k>A�>j Q>fA[?�vD?�ɞ>�}8=%:���Sս+*��������;�q��cN���yL=�ߴ��,ɾR�4���������)�T���:P�5�T�A8k������20�JF��%��-?���<�dɾ�L�n<�����-5��]�	�}�A��2I���2�M'{����?U�"?�^���C��y��KT>�>�͍E?G�s=S�0�*��ػm>b�-=�{>���=� s>9�U��Q\�Ϙg��#/?�?�n��tU���l">�����0=�+?	z�>���<[�>P� ?�9�;`Ƚ �T>�26>�4�>a�>�U>
~���q��D7?��U?^�����
Q�> �¾�ls��(=yx>iK3�%	��]>{��<�������3N��)��;��W?��>lP)�O����F���/R=�w?Z?�6�> Wj?�C?%��<���1ZQ��b���k=�V?�{i?!�
>�����о$���pS5?-ge?��I>N?f�?��\�.�����?�Dm?�}?P����|�##��E��r6?Ds?�]�w]��$��
9D����>���>H� ?��9�G��>�4?�H�܈��Y\����5���?�@T��?�=�����=q��>�H�>b�Q�b�Ⱦ�x��Y��z4F=��>�!����q����M�0�ր2?���?� ?�2�����BM>[�p�0!�?l�y?�>i�R��=B%�at��QӾ|:3�(G���3��%6=?����;8��Ͼ����ϔ���N'i>�J@�9(=:h�>E�ܽz�߿1Q̿�>��~��]h� �?g �>�z�� ࿾��j�"/K�^�6��wR�r�վ7d�>)+c>h��6���b�&c=��j>N��>�1G����>%�Ⱦ���%/��2&.=*6?��->G��<��y�\q���?z0�㜰�m���F�D�t?��?�pU?�N?��ѽԽ����>����l?:�t?�7?/�)>�)�`mA>�u?�ō��GT�-�*�R��}A>�~8?�p�>:(���3=v�0>��?N�=�8����.�¿f��%�?�?E���6�?e[�?�3?q���9���� �@
ɽ��K?R��=T�ھ%����{D��5���?�?�ν���_?��a���p���-�c�ƽ}ۡ>d�0�_g\��W��ˢ�SXe�����@y���?g^�?3�?��5#��6%?B�>b����9Ǿ���<��>�*�>�%N>]@_�"�u>%	���:��k	>t��?O~�?�i?�������U>�}?F�>��?��=f�>���=�հ��<���">�p�=U�B�jr?��M?�/�>e��=�*9���.�fKF�8R�Q-�ƪC�=B�>C�a?
�L?�b>���\�6��'!�7�̽�0��ἴ�?�]�,�S���H5>��>>��>��D�4LӾ��?Np�1�ؿ j�� p'��54?:��>�?��K�t�)���;_?%z�>�6��+���%��}B�c��?�G�?;�?��׾�R̼�>4�>�I�>��Խ���h�����7>�B?}��D��v�o�f�>���?�@�ծ?\i��	?�#�EI���e~��m���6��*�=��7?r1�D{>
��>�>�={v�ɵ��:�s�X��>.;�?|�?9��>��l?:wo�p�B��[1=�@�>�k?|x?G:S���{�B>g�?6��)��V��f?��
@�m@^?�ޢ�+ǿ>�x���ʾ�W�����Xr���,Z>	Q=��HS>�G�=Z�@��o=�MZ=3Þ>�l�>��=g��>�Y+>a{����п4���k{���>�w�*�=cA7��L=���#�<o�aU�&��<� ���Ѿ��}~E=2��=�T?�T?&r??m�H��>� ���,=��"�2�=�I�>34?4�L? �&?D��=����G&c�n��)������>�>БR>���>��>�L�>W!<ID>�'B>�6�>�|�=P/E=UH4;s�<�iO>���>	I�>��>H�;>�.>J�������Yh�x�{^Ƚ�٢?y���9J��,��E���h���V��=)�.?w�>�V����Ͽ=���^.H?���ֶ�+�-�@�>O1?@NW?d+>�Я�9V��>_���nn��>��βi��(�LDR>��?$�=���=݋F���"�d�Y��Ծ�Б>� /?��7�*�O�ҫt�%D"�!�徆�l>�E�> =�"���:����}�Bc���>Ł3?
�%?�,:������B)���F=K �>Z��=�S�K{�>ѯ���=>k_.�ٴ��)��>�JO>��?Y�=�]�<
i�={�V�K���>@_�>��=��9?�$�>��j	i��v��������>���>��>c=>����P>�4�>$&�>/'㽗�=�/��e��I]>k}#���6���u�>h�9=EK->�s=�q�����*���~?���䈿��Od��mD?%+?; �=��F<��"�4 ��|H��B�?f�@m�?��	�ޢV�<�?�@�?�
����= }�>=׫>�ξ��L�±?ƽǢ���	�K)#�OS�?��?�/�Zʋ�l�x6>�^%?�Ӿ�h�>�v�IZ��E��u�u���#=-��>g8H?~V����O��>�Lw
?�?�^�F�����ȿO|v����>4�?���?d�m�pA���@�Q��>&��?gY?�oi>�f۾^aZ�ȋ�>»@?dR?��>e9���'�{�?�޶?˯�?X�K>!�?�~?7R�>��Q<E��#X��^���U1�=ˤȽ�W{>Tt >O0����:�@Ϗ�]F~���i��M�b�>l`=zx�>�t����?�>�&��N��\v
�!��>А�>��> B�> ��>���>l&�>�>��-��-w�&ۯ�k�K?���?����2n�\N�<P��=m�^��&?vI4?�u[���ϾXը>��\?]?�[?�c�>��<>��2迿;~�����<��K>�4�>UH�>&&���EK>&�Ծ�4D�Up�>5З>����`?ھ-���O��BB�>[e!?j��>�Ю=T� ?u%?@e>W�>��E�cF���|>� �>���>B*?�:z?�a?ڋ��6�5�-}��zx��`._�_p:>$w?�C?���>~���cg����������M<�$=?��d?��۽��?ź�?F�<?��>?���>_���޾�����Y�>�?�&��@��T*���$��?�h?.��>z�d��ϽD K��`
�K����?7*X?��?��ﾸ�[�����	�&=�q߼�"��ކF�poڼ�A.>A�>/˽��=^(	>�>��N��pL�<�A<�bT=��>�Q�=��,F����+?�⭼?�����b=�Qm�HkB�1��>R&d>�D¾:�^?@J��|����;���.\����?o�?r5�?:
����c��,>?�8�?s?���>Ŝ���޾�/�=j���S�|�>
&�>���;��پ���⧿$7���$��40p�&y%?%��>��?7�?ϜC>��>K>��WF�e���ؾJrN���徳Qh�z�+?��Ҿ������=�_ξ��p�K�>��>�e��>W�5?��>`;�>l�>1�x��g�>N�>ɱ�>�k�>���>��>g"�=Q�=�_��S?�����k&�a��7���B?3�d?���>��m��{��!]�SD!?!4�?il�?���>��h��?,���?P?2w��?��-=/]�ë�<���-R�&a��F[ܼ�"�>�'Ľ�Z7�WOL��\�L?چ?��P�"ʾ�ǽ_�����=��?<�)?7�)���R��m���W���T�ɳ��ee�����($���p�����Kڃ�5����(�nB*=Ŀ*?�,�?}7��
����h�?@<���]>>��>ߢ�>��>m�M>v	�[�1�-�[��'�����^g�>�m|?4��>�>?I?d=`?d�]?k��>ռ�>TCž�?�ka<�N�>�p�>��D?��0?�k?�[,?\M'?��?>�6��ﾙ�ξ�� ?�
#?%;?��>$% ?n�#��#��!7����:c؉�dg���2�=N�*�x�����B�j�=1�9>0?�=	���$�1%�f��=Ms'??+�>��m>�c3��X��<.>{�>�kt>���>��¾�t�t�#��>=��?���
�=6�:>��):4j���D伖S�=��=%n�=��B��Z��}D9�ǹ�=10�=_���w\���<O
>/�=h1 ?�?���>P[�>�?������Y�����=4�`>	>[>�'>.�Ծ~A���͗�:h���y>�Ȑ?�1�?h}=�f�=�C�=�Ξ��W��H��O޼��+�<F?�#?-�R?�V�?�=?�="?0�>������G���[����p?�u:?M^�>�	��ƾ[:����&�k�?	��>�U�sA ��Q������콪~;>S�%�w��t���t�.��U>������_{�?D^�?�m���D��AԾؕ��%$;+�I?B��>wQx>M�?R�,��h�4\���>7;�>LH?�U�>�	+?V�?�Ѐ?�� ?a�u]ʿ�����я>���=,|4?e�]?�%�?�]I?>�>,��>Gͽm�о7�(��*<��ý놘�b>TWd>=#�>�|"?�^�>Z�@=��a=N:��������>�I�>L��>Ӂ�>	U�>��`>X&��fA?��>�=��Z�hΓ��r��4����u?���?6i-?�ur<���^�N�-P�>��?�L�?X4?�$��Y�=�f��(���M����>w��>@�>�n>�^�;��'>���>"��>��)����mW7�AD���?��<?�r�=�Ŀ�<���x߾Ǿھ[�+����ϻM��g&>}m��m@8>�G��R��i�Ծbjd��O�H�:V�������s��?6����t�<�G,=�H�=5Qd=����c<�\=�A�<ʳ�L��<BY�� �=�$�˵����=<۝��i�;��˾|�}?!8I?m�+?G�C?�y>�3>p�3����>����A?_V>��P�B���Y�;�������Ƨؾ8r׾��c�0ǟ��F>fvI�_�>�=3>�O�=4҈<m�=�!s=���=ȞP��=��=0`�=�\�=���=��>K[>�&w?.�������NAQ�'��Ї:?�\�>���=��ƾ$@?�>>2��,���)f��~?��?�F�?&�?��h�J]�>ь�������ݑ=�9���i1>Y��=�=3�)��> J>�`�:��F����/�?6y@�w??�ʋ�ҫϿ�.>�(O<�f����[�AU�4�Ⱦ��������?�ɿ�{����=��L>;�&�rס��H��|e�>��>pz���?����=\eC=�H�=8�>f�#>f">���=���-sj=aы<�nS>���=�u��]��o�н�?��0�9��u>j/+>���>y�?�9C?|?��
?����)����߾'
�>?�Q>	g3?f>�D�>�Y�>��?��=?�;P?��?�����a�>���>����>o����nU���:	�F�`?O��?t?�>�Q>��=!>�v^W�(���b�>��??�?@/?�T�ڡ��Y&�b�.������G�s+=}fr�xSU�n����k������=�p�>,��>��>�Qy>��9>G�N>��>i�>�-�<El�=�n��"�<������=턑���<��ż���'���+�m����j�;o)�;f�]<R��;��=��>n��=%��>,�\=ʱԾ��d>��h�A�T����=zȗ�qBC��[�`���������{I>eD>kȤ�a���U�?~x�>fA>K��?�g?�h>������������PW����=5�z=}yc��W+���]�:�F��Aɾ^��>I��>�>�ڬ>��$���N�:Q�=�y�bN��#
?�Ӛ��	��U=�M���Ĝ�1ۨ��|��@�</o?V���ŏ>�;�?N1O?q6�?�{�>ȹi������q><̖�Xw���2�x��;�Ǿ�F? d?d��>�0�n�I̾����ڷ>3HI�!�O�k�����0���η�	��>l�����о�%3��f������u�B�8Ir����>�O?��?UAb��W���TO�O���*��&r?]~g?.�>kK?�<? ;��O{��u���q�=�n?1��?�;�?
>?ܛ=�4=! ?P?z'�?�?"�Y?���j��>��,�om>x�='u>�C>!4��tb�=5[�>��?@K�>�ar��. �i����!�SG2�TY�=r�3>>3�>\#>w�(>��I=�ȃ=E��=[�V>r�>�V�=�-q>�5�>���>����,[׾U^1?؁p����>�lh?>�9>�ZK>3�\���ө!���⽥.>1��Ly&=a�f�^WA���1>G��=8H?��ؿ.�i?�p=-E�^�$?�r�U��T�Q=��x>i?��x>�r^>��>Y��>�׭>��1>?�|>�,>&Ⱦ{>y;�����;C���O��RǾk�o>�͞�q� �H����Խ��H�*h��(���)�i��g��p�=���={��?�����j��!*��^���

?���>�3?����t�#>D��>���>����^���ۓ���'߾X��?k��?�=c>x�>#�W?��?|�1��3�LsZ���u�'A��e���`�$፿����t�
������_?��x? yA?�t�<%9z>y��?��%�nϏ�K'�>�/��%;�N@<=�)�>�(��>�`��Ӿq�þ67�=IF>�o?+$�?YU?�YV��Ke���'>#?;?��2?Cu?�-2?'�:?%����$?��3>�?R�
?&%6?gx/?t	?�=6>���=� w���=����_|ֽ˲ǽQ��t-=�Ą=�*�:y��;N�=8��<H�>�ؼ_�;d=��P�<��==���=���=���>1\?��?Xƭ>��/?�2��\-:��ȱ�oaa?��8>,��=�����)��������k�Q?���?k�\?+�>y�:�����>B;>��e>%ZT>��>A�������U!<�tE=ư$>��=;����-���������.E��ҹ(>�R�>9��>�k �z�+>C�ɾ��ྛ�>}8h�����@�*�=���4�s�c����>��B?�w?�P>�޾}�A��G_��vB?�5?Ӽk?��U?���C'��xV?�ͭf�U�����>�Ƽ�l��"��� א�W���L��6�j>�y��od>����;C�u���m��
��ϻ^>�����=����l��LI��]D>�>D����]�3i��e����x[?̪���ؾ��:��ȃ��BH><�>j��>�T��{P���K�@x��+�=2��>(&,>1�ͼ���pb�����&�>=tE?!�^?��?Y@~��Ss�%�A��s���裾P^��l!?�ȧ>?�U0>Ç�=����|��|b��E��O�>Ҿ�>x�/#E�}`���r�D� �s�>�?��+>��
?�S?��
?�o]?�&)?]J?ʐ�>O'��t��Tp'?�ȁ?Z^=ɋĽZNT���:��/�w�>� ?�]����>~�?�?i�?�GV?	�?r��=�g�P?6��]�>\��>�V[��߰�S�D>�P?��>�%R?��??�>77������b��o:�=�3>��(?��?��?� �>���>땠�)�=8>�>��c?�ق?}�p?��=�H?��2>`�>vТ=��>�7�>��?�O?��t?�RK?T/�>��<���� ���T��l)��&͸�ĚF<���=>��8 Z��I�\4
=E��;�����D��M��".�9f�����;�+�>.Hu>D�'�>�\��1�����;>�I��H������7BH�O��=3es>�?rC�>"����=���>�{�>o�S�(?��?Q�?�����c��ԾB6�&:�>�T@?���={0r�����/+p���e=��j?�jZ?~'N����db?ud]?�j���v<���þ$Ud����/	P?��?��I����>�P|?^�p?x^�>>j���m��Ŝ���a��jo�r�=�ϙ>�B�\f��4�>D�8?���>!e>�=]�۾��v�2X��1�?DG�?Un�?���?��+>�fn�}�߿�oھ�酿?-l?�0�><���/�7?�y�/���������-�������#ݽj�x�,V����,��CP�"Ѹ��>',�>��x?`B}?n�Z?�ũ���f���H��閿p_�_�־�t!���m���K��m@������$���Ⱦ���/w��q�X(3��f�?O#?Q�F���>���h�̾Nþ���=&�z���۽�w>���J;�=��k=O�\��K������X?�Ə>�D�>�??^�O�G�;��� ��?�>���S>�r�>X�:>�k�>mI�V7���̽��ɾ��C���Mt>�Nc?L�J?��n?�I��[2�F���?!���@������NF>ι>$��>�W]�!���%���=�˧q�G,�%=��d-
�Bj=��2?ǁ>%��>�&�?'b?o�
��U��/�v���0�ܰz<)��>Dsg?���><�>�?нR4 �ގ�>��l?���>@��>������$�v�(�����>��>���>� ^>W]�q�_�//��A���7����=�e?,���[h�Ă>�WO?�j#<>��<�v�> ����� �������:>57?�n�=��C>�[��y��Rv��'���V*?��?쓏�$l'����>��!?�?�>��>��?+�>��ľ��u<�?�w[?6P? �E?d��>��=Y3����ٽ�����=̆~>E�p>%��=:.�=e\1���Y�!�.v=B��=��5����SS�����;ӺU<f{=JaG>I�пd{R�P ���m#�#��	-�����6�=t0B���;�|��������HؾJ�������HQ�*썽Zi4�b�#��{�?m$�?�k��l��B�������Ș�'X?jIоϼx=5�\����mWѾ����h̗�.�%�Q�!d���[�{�.?k�R��,����u��q?W\S?mB?�޾����
�G�j>�d���{�[ʞ���aǿn�0�s+q?`��>�� ������>�y&=WVs>�Ҫ<|]Ǿ�4�gG�<;?�j0?!5k>�u����ο*ο��ڼ�J�?K @��:?9�p���Ә��1?�??]��=�iK����ܩ�S�l>�W�?�^?�ū�Q�>��s�=��[?�p��}�G��j-����=�Q>���B��bb�=P��>�4�=*�m�~ࣼ��>Y� >�z��Lt�=z/ �iPP���>KD��ɂ�
Մ?az\��f���/��T��dV>y�T?v*�> 2�=�,?�6H�}ϿR�\�*a?Q0�?ޥ�?��(?#ݿ�Nٚ>��ܾ�M?�C6?���>(e&���t�ʉ�=�V�����㾜'V����=���>b�>!�,�v���O�������=�E���ο�����d��<�v�<���n�-��qp=?��{"��k灾��č�<�z�=���> ��>�hs>D]U>�]?�tp?��R>�9=U�"�|�������<<��A�� @�J���ξ*t׾�Ⱦ�������6��LO6�;��=
�T�J��+�hYj�m�-�`�>?�>�ֻ�ѲD�>QԼ���2���^�3�3�T��β�7)1�y�f���?��B?'���7F�������6���,T?�z��� �� ���+�=�>e<�p >��>��<UM�ȾO��^�'S)?��?�O������m�O>��!��hS<,	)?)9�>�Ŷ<���>��?9��n�N�_>�9>s�>��>�e�=�J���媽��?KtP?�/�����u�>l���3ӊ�aƭ=��/>�Q�I�L���4>��m<#����V�&y���>=Z2W?��>�(�@�������Do��I>b�r?=+�>���>7x\?v�<?�'=ˏ����;���gE9<�kQ?�ve?6M	>yI��AݾM޼�*#?�`l?�-\>B�s��ʾ��7�Q����?�WZ?$0?7�� �������>����8?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?p�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������]�=J�|��ݮ?{��?�����^�=���r�v���������]=�������<��ޙ:��ܾ����͢�!!�We>s�@wC����>�$��3ؿ2�ȿ�ڍ�d���"0�V	�>��>�l*�ݓ��3te��w��@D��A��������>/�u>��0�v⽌S�c�\�[n=>'A�>
L���#�>�����#��� 7��sڽ޿�=�ԋ>���;U������֑?�����Ŀ.ܫ����?L�?An?R]'?��!�$��a0��BX���:p?��~?
�W?M%�I�%���Zd?���SC��^��g���=��;?�|�>�2�
�e>���>���>��s=�Z�������ǿ8�!���?6�?��.�>�p�?L7?���H��>>Ⱦ�2��@/�|�i?=D*>�۾q���/�A��Ծ
?@))?9y̽��־�_?>�a���p�{�-���ƽС>��0��Z\����-��,Ve�: ��@/y���?�\�?�?,���"�M5%?9�>����?AǾ.�<Ww�>T4�>C@N>�D_���u>���:�u	>���?{�?Ej?���B���^>��}?� �>��??v�=b`�>�W�=	����U-��r#>��=��>�à?ŢM?�H�>�H�=m�8��/��WF��ER�#���C���>��a?h�L?|Gb>�5��2��!���ͽ2V1�W�輠O@�+l,���߽�#5>�=>��>c�D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?mQo���i�B>��?"������L��f?�
@u@a�^?*�HӿRҜ��d������> �=�k4>N��� 5�=V�=�*���ٹ���=��x>�[p>��>��a>'�T>�/>�]��B�&�C%��!��7��
�]��)�B�݊
���`�i.��wž�ݾM,�� �ǰx�3:�p5�>��[��=�U?�Q?��o?�� ?q�t��O>�����=�#�y�=�E�>�"2?KlL?6�*?���=}�����d��a��=��3����p�>rI>���>$7�>ͭ>!,깳�I>**?>>��>G)=�R���=�SO>�B�>r��>��>��b>0�a<<C��ô���[�;O������}ĝ?�����_�u��XE��%��昕>z/?S�!>�e���ӿ�����R?[�j��\���>�nN?��?U���Z�>��ME>�f��Ožvߗ�N<��o�dRP�

c=���>�P�>� >k"2�/�P��%�,䉾l�w>"9?d�Ѿ
�-Bb�;F�X���Ku>�t�>������u���8`�⎫��y�>��2?~�?;��p��;�
����<�>�}&>��c�*�Xb�>����u��9�]�So,��\�>��E>4N?ȌN>���=�Y�>���r���[��>�`9>�]M>iF?��*?fQ���#���8��4��|�n>�_�>���>&�>�*�>G�=d~�>�Nk>��/��U����ֽ	�[��>�YǼ��j�2N{��s�=���{��=ۋS=�H���A���X=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��L��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�/)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ%e�>Z�YW��#��t�u���"=��>�/H?0h����O�G>��d
?�?vl򾅬��\�ȿ�}v����>u��?��?w�m�OA�� @����>��?�cY?;i>([۾2yZ�Qe�>ڸ@?+�Q?�@�>?3�[}'���?ն?A��?(h>���?���?��>Դ5>��׾Ǵ��<=���1> /��Q=�>�����
E�#���i-��G��d۾�>f
=���>-��ା �>�w�������nA����>͇�>��<>g/?\'�> ߴ>�>6>㖮�
�/<�?����K?mc�?���On����<��=W�]��?b�3?��v�4�о��>J�[?�i�?	�Z?X�>�{�0���ҿ�b��&�<�2L>&��>![�>�����I>Nվ|RC��%�>o��>4u��U7پ?/���ڻiÝ>;(!?��>���=� ?�#?b�g>·�>54E�k����+E���>%o�>�?�Q}?��?���B4��`���¡���[��gL>��w?fz?0��>s���$ĝ�6�#���,����+U�?G�f?�/�??�ވ?��=?�C?nxf>I����Ծ����s�y>�(/?EaC�#�n�U>K�H��=/K?���>��>��;��U�Ӹ)�F�;���b�P3?P?5��>�\1��E��v��ż��;=u�<T��P�<=�?�>��=��[��s>L�>[">_鋻g�'�&���1>�5=u��=��i�>=5,?TE�Qσ����=��r�O�D��>�~L>����B�^?�f=���{��	��yn���T����?-��?�a�?U*����h�I =?w�?n?�	�>h��]w޾Ҩ��`w�;dx��Y�.�>���>dwq�i得��������?��4�Ž�1!��I?-��>J�?F?��h>��>�{��e����%s���D����.H���B��$��뜾n������<Nž�Yy�? �>ѽhS�>!9? �o>�ߊ>_Q�>�� ����>=Ε>3�l>3��>�ݤ>-�A>��=X.=:�HR?2a���N'�X~�䜯�B?��c?���>ml��X������u?*�?>=�?�w>@
h��a*���?T��>���4
?I@=����X<,���]�Yҁ� 8�\��>��ֽ�;�5�L�){c�,
?�?�!���W̾?�׽K\���r=%7�?7 )?�)�X�Q���o�c�W� S�"q��g��򡾕r$�2�p�'⏿�R��^����(���*=�_*?��?>���H�@+����j�(�>��d>
��>!T�>�ս>%KI>L�	�˔1��]�L#'�ۃ����>#�z?���>��A?/�L?q3t? �W?c
�>�ӓ>��龐�>i�;�8�>�6�>�*B?m5?^�(?�
?��3?�6�>F�&���ﾥ6�$��>�� ?��?�*�>�*1? �.\+�D�V��[=Q��6��d	J=���/w.�J	>L�>�>\�?w.��:�P ��/f>B�7?�S�>�B�>u��P}�hf=���>|?)�>O_���-p��T�¦�>�}�?k����=��$>M��=��ɼ���:3��=�ռS(�=���`1�?�Y<b��=��=?���*�339��$<V �<m{�>?�?�׊>�i�>�c��� ������=�Z>]BT>t>��ؾ�a��$����g��y>Y}�?�|�?�?i=*i�=��=�y��-l��6�����Cv�<��?b#?�OT?-e�?%�=?&#?�>Y$��H��Ee���1��e�?�N?b��>|��4����ˬ�5R�3;7?�I?��m�o����[�����<=qM��(�8��<󭿃P�u@>�!�/�=���?ro�?՛���bn��[羹:W��Ǹ�#c0?v��>��>)�*?Y�(�� ���f�[Y�=V�;?��:?{��>�R?�߉?��e?�CE> ���Ѻ�s����>�Ƿ>��??�ֈ?��?�no?8?��>���=�AP<Է�ԴA��}L�n���)�>��>^��>��?+k^>y�J�rX�HY=���EwM>z�>%�?�	�>�>>GC>��J�g�G?���>cH������=���q���6��&u?�f�?``+?)=���E��@��=��>�B�?]��?��)?vrS���=�,׼f䶾%�r���>�#�>�ޘ>�֑=�H=o>Ʈ�>���>\�]� V8���O�M�?��E?70�=|�ſ��q� �p����$Pf<�.��Xe�ߋ����Z���="�����������"]������ܒ�!E��a����{����>�g�=}�=���=L��<�9ȼ�A�<W�K=�\�<e�=��o���q<�9���s}�����&J<f�H=D.�[�˾]�}?�AI?��+?k�C?��y>F�>/�4�V��>c����8?3V>�P�݋����;�k������8�ؾ.u׾��c�jş��B>�6I�9�>�83>
�=���<�.�=�vs=��=�dH�_=�3�=�i�=��=���=S�>�K>�6w?X�������4Q��Z罥�:?�8�>g{�=��ƾq@?}�>>�2������xb��-?���?�T�?>�?Bti��d�>M���㎽�q�=G����=2>q��=w�2�T��>��J>���K��E����4�?��@��??�ዿТϿ5a/>|�>��>��I�Q�0�H��=�C��
L��u�>��"��޾ۺ�=O�'>HD�����V=ྚ>���<��x�/'a��T�<�Aƽd�=j�A=t�>?�>B��� 4���1=
�=���=$�>5v0=��a����r�={>uU>Vuw>�S�>W�?k�K?
�?���>��M�?篾˸ھ0�>�>G2>?�G�>d�>���>u�C?.`N?^̆?�g?�S<�v�>l��>i�3�� ���2'��վcӾm?�?�Z�>\Ƽ��!�!^$�_����� �>���>=!
?\�	?���.B����F��}B��*d>5�[������̒>M�;;Ӿ�,��~�=n�)=��>F��>D��>-V�>�8&>I��>X��=��=���=B�P��J�<���=WKH>��>1~����!�f����o��I䉼ze�S�i=Rv�<k��YS�<�h�=�|�>�r>���>j��=����_.>����&L�؉�=.����A�O#c���~��/���8�`�A>��X>u����?�?�[>�=>X�?Ԙu?g� >� 
�h�ӾqǞ���d���O��=�>':�a�:���_�#�M�n�Ҿ(¥>T��>�>=�>0�'��MP����<��;�Q:��'?�q<���ս?>$H���aƿ�_����Z��9>��r?Wx����>�?��? n�?�?�MK�g!
����>,�b����5¾�Wֽ�ٜ�ƒ>��?�C&?�
���t�2�˾�����>�E���O�����O0��� ����_�>T��"�Ҿ��2�����M���B���t�E�>��N?ջ�?��d�x���� P���@x��?�Sg?��>�3?�S?�������y����=�n?��?Xb�?R;>�Px=�V <v?V/9?b-�?�[�?n�t?�2��A�>����A�>m>�>95g=dt�<��=9,?` ?�b�>뫃��.���^�ܾ'Z��u��==�>#��>���>R�>�^>�\>��=��|>B�?��>V�>��>��L>������45?h��=��s>4DV?�HS>�	>��=� f����s��<n= ���x��R��q�$�">�$�=0#�>��ѿK(z?�Cc>t���?&����0�=C/>=�ν�X�>��l>�C�>��>|��>� O>�^">�;�=��ϾC�>�}�/!�dC�6�Q�8�˾Q�z>2��P^$�+��"��'{I�E�����i�}O����<�"��<�#�?��󽒂j���(�(���?��>Ri5?�\��*C��<�
>͑�>Տ>g����� ���ᾕ9�?1}�?�-c>�!�>��W?[�?a1���2��wZ�_�u��A��e�׻`��ݍ����
�r7����_?�x?2lA?e��<z&z>(��?�%��я��J�>�/�,;�ߓ;=�K�>����a�o�Ӿ��þ�>��FF>��o?r�?�]?�hV�)�m�'>��:?��1?�[t?�1?E�;?���B�$?^r3>�d?3}?P5?��.?��
?
L2>�#�=5��E�&=#���~犾eҽ�˽�����2=k{=��8�g<��=���<M�j|ټ8;;z`����<gM;=�ߢ=��=}f�>ӺY?�5 ?(^�>��?Ɨ!���E�^����.B?�LR>�K���(_�HǞ�8��>�{?\�?)�a?�I>.~A�#{3����=<W>{g>��B>y��>��$�
v�T�=���=~D>��=胲���M��jӾ-��`�ʼ�U>���>j�>�)p�
Q�=;���է��A<>'E���ʋ��$��.8���3�����>8B?�)?���='��aڽ��l�13#?�;?�j?W6\?������̾��@�#B����F�>�*)=Z�þlܥ��̓�{�,�\�3���k>��K�M�����k>s9��Ɩ��≿�_g���<� >��'�I��(!��w�5�~�d*=>"Cn=ꐲ�C���1������Y�S?��
>�3�B9��J��'�3>�ڳ>�{">	��=Z��L�W'�ka��?D�=�m�T|����ҍ��m�>E�C?��X?��?�}E��,w��6���|���W�����?�A�>�(?$�a>&�>����!w�]�`��D�gX�>���>��R�7�l���g���͛�'�0>�)
?w�>�4�>^LG?�S?Bh?��/?��?FI�>#,.�����U%?��?@�\=X~��vtp�9%=� >����>x#?XB��_�>Y?��?��)?�*W?v[?��=����C����>{�>��\�N%���1>�%O?�޿>�P?"��?Z�5>P�>�Ͻ���Cʽ�X�=�I>br*?�>%?#%?[բ>���>��pɇ>��>>p4?Թz?���>Q=N�?�ؾ�f�>���>.i!?��y��M;?�D�?��?�yK?�?��=�G��r�Ȯ۽�V}�Fü�]�<"`�=������rr���0�=Lu��^���߼hh��E�<�[�<C<��>��l>>7��5�'>�Eþ�䓾4�8>�»t����x��}H����=�vY>I ?W�>�%�ۡ�=gɸ>��>� ��x(?�#?|y?�U�8�\���پb�,����>�QC?W��=��q�5�����n�U�{=�Yn?S�V?x�C�ܭ�U�b?��]?Nf�<=���þ��b�Ȇ���O?Z�
?�G��>��~?p�q?���>�e�z5n����=Fb���j�M�=�p�>�Y��d�2�>Ԟ7?
V�>*�b>})�=�r۾��w��l��*?���?� �?r��?!+*>@�n�3࿅�־���N�a?qX�>^g��ؘ5?��a��������^Am���Ӿ"�ھq��Xi��z��t�[��T��?�G���f=
�?�L�?!Wx?��m?��6�x�+=���z�/ia�B!���%���6��'U�F�V�	@z�V�ob��Ǿ������R�@W�4��?N?��?�}���������l�>ǭ���Jm��]->wc'=.X>K䃼�ڑ�ƢO�����C!?�q�>���>8�F?Rkf���9�H��?�����-�=���>i(Z>f��>9�Խ%�z��6нy�Ⱦ'���7�r�*��>�e?#�M?ة�?i�o=������S@��%u��?��	��>��q>ʮ�>����c��_�"��!M���E���㾥 ������N�GyP?��>&�h>���?�c/?z���x���yM��"S�)*�<C�?6J?8X�>;2,>���<�T�p��>�u?��?g�>Z㲽����&���Jc�z�?��?8.:?�\�>�ٽ�6t������l����Ƃ5>*�w?�B֍�-�>'^?�w�=�L�=��>�� ��?����w���go=�^	?J�>K�>��)�#��T�vu��{�"?�+
?�՝��0*��Ae>�[?��>~~�>u��?<ڣ>�ξ��l�:�>9wZ?G�E?�<?æ�>�:=&:?��ý��~�=��t>��_>�ѭ=�F>���׳n���C���i=�r�=������ݽ+�.��{�ƾ�<���<'�4>��࿡�S�q\ݾ� �%��ES	�d�=�1� ����@'&�D���ճ������Z���T�u�%|D� ���F�����?4P�?z.�U�D�9��� u�tǾx��>�肾�a��=4���{��L��˖��:蹾�d/�q:=�S�n��q��!$?!�����ǿ�ҟ�
޾�i?�� ?��s?p�� �_�7���>wb^<��L�W��5ɚ��[Ϳҗ��@�\?���>��������>EȆ>�.m>o>.��9���jg<2�?�Q-?�S�>[ q��Eǿ�0��
C�<e��?��@��A?I'����M[g=^s�>J?�WB>�t3�~��KQ�����>���?i��?��h=�`W�W?�?^c?�M�q�G�3�H��=��=��=�c
�1K>�S�>���i=����� <>�I�>e�>�����a��R�<6�U>ݑӽ��s�5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=c6�쉤�{���&V�y��=[��>c�>,������O��I��W��=�7	�|�ҿ�>+��)�c�<�P޼��9}�U�@S��s��aCI��*��[�ȫ���;&��N�=9�\>1�<>�3>1�c?Қ?�)�>�q�>���E¾)�h��0=N۳�&�}���B�=�k��&W�������r`	�SM��/�KO�{:��U=��K�Y���Њ#��jf��Q�*O=?,���f ;�uJ�iW��8V��L۳���u�̕���o2��|�J�?4`=?���� W�����q%����"S?��ѽ��������2�>��_����=�;�>��9>��ľ�&'�,�P�i#?	�?-���6Mm�P�7>�4������F?�8�>�G���M�>R<?�N��$X��L>�E�>+v�>��>fÎ==±�*=3�{v?py?�(�����b�Z>����9.�)�j=\q�>Ғ>�#�I>-s>z��=�&����^�Žϑ�<� W?H!�>��)�y���%������7=�Jx?�?���>5�k?d�B?@��<H��U�S�l�
���|=��W?^Yi?�f>����b�Ͼ�M��6? �e?�N>�h��H꾥�.�����?Ȟn?�&?a���~A}�H)���
��F6?�v?9Z^��X�����E�V�A[�>)6�>i��>��9�ڲ>�>?ު"�H'�������-4��ʞ?	�@���?��F<q^��h�=}R?�'�>�O��3ƾ�Ǵ�����\p=TL�>�E���(v�ڶ�96,�!z8?	��?U��>N���ˠ�k�B>y�#����?�?�����=�,�vS�GC��(�b�ޛ���J�N\&=��þ��)��=�?��n��+҄��R>�o@$K�=$^�>󜚽[��Ўп_\����վF��?4[?�W�+�)��Y�J�ȭ,�;-|�+��p��>��>w)������{��<��������>[�v#�>N5W��$��vy��3R�<y@�>O�>.B�>rº�Z&����?9����EͿ|J��&��Y?�)�?*ʄ?Ѓ?>{ <b~���z�(G�!�F?]�p?O/X?:�_��ZE�ҿj?V��gS`�ˊ4��LE��U>@%3?�<�>�-��|=�>j��>3X>�/�8�Ŀ�ض�����=��?��?[n꾱��> ��?<q+?Ij�F6��tS���*��OG�qAA?h2><�����!��+=�}ؒ��
?{�0?*{��-��_?��a���p���-�w�ƽ�١>H�0��d\��P��T��Xe�����>y�k��?5^�?K�?��#��5%?�>	����8Ǿv�<X�>�)�>�+N>;P_���u>�'�:�i	>t��?�~�?�j?��������S>h�}?�G�>j�?��=���>���=����n,�R\#>�n�=i>��?�dM?�7�>��=�y8��/��MF�ZR�w��C�X�>��a?��L?�^b>Y;��QO.��� ��ͽ��0���޼��@��+�v!޽�74>Y>>J�>'�D�.�Ҿ��?:e���ؿsM���{'��&4?��>�?����t�k7�Z�^?Ã�>U����(�����z��?�.�?(�?	�׾79мr�>�֭>AC�>c�ӽ7���B8���7>KB?��WL���o����>���?̭@m��?c�h�]	?���P���`~���� 7�5��=��7?,0�i�z>���>��=�ov�����1�s�M��>|B�?@{�?n��>Ȯl?1�o�-�B�=�1=�L�>�k?�s?�n��%�B>�?G�������K��f?��
@Zu@{�^?c�ٿ^��������l�_�c=v��=�<�=�!��ѐ=P�������~�<� >�`>[�{>�[s>!�)>�z�>��>6���;�'������Ș�3+�(:�u�
�}��"��������WJþ,��Խf���*�z}-���P��&$���=��U?a�R?^,r?��?i�v��>�p�����</���ߒ=�z�>#�2?�M?
�*?jԆ=���c�ʻ���y������K��>�N>2��>�}�>�s�>�I;��F>`�@>/�>.��=��)=\�;�{�<"�T>�,�>���>>��>�(>��'>7������`s��m��X�����??����?C�c�����������=��?ɳ�=Z���Qo̿�^��:�G?���<&�8�ؽ�&>�v-?"�D?��=�w���#6��|">`ǽ&hn��>b`��ԅ��"�FU>ԥ?�-h>I>A�K�S�5��6�d��i�>/�D?�˾􀜽�}��������US�>f�.>�S��&9��ϖ���a��Y��S��=�c+?Z�>=�f��R���|2����$>,P�>�s>hֺ���>d�=Ӓ�==߽�䋾M}.>*+�>n��>�+>�L�<?C�>7����׈��D�>�o>�5>�:?�?�\V��������C��A�v>?��>�Qr>��>J����=���>�it>=5����i���� �vff>����	9� ���r/�=��g�/�>v��=M���F/�I�\=O�}?굧�ˇ�VU�$����E?E�
?9�=��<������ %�����?d�@[��?�	���V���?V�?x���b�=�|�>}U�>x�о��K��s?�����"��K�	��!�(�?�O�? {B�	�����j�!�>�=$?�t־�[�>�v��[��=����u�ͭ#=а�>B1H?�R���O��>�4i
?�?iS�ߤ����ȿZvv����>	�?K�?��m��<���@���>���?�eY?�ni>*_۾�~Z����>�@?��Q? �>�:��'���?�ڶ?���?:�~>RB�?^��?.��>Ԥ�<n<�r�οQ���+K��е�C��>w��>��Z��TL�λ��&T���}�: ����>�c�<0Ө>�IH�7����p>	6;�}��Bl�����>�R�=���>���>�a$?�b�>u�>���=�}i=�vC�p��OL?G��?��oum����<8�=�/]��?@4?f�t���о��>%W\?�ˀ?�vZ?�	�>I��Pk��t��a���0֔<��J>�>���>�����J>�"վm�B�i�>AZ�>�㣼�0۾1���|E�Y �>� ?��>�K�=˙ ?ɜ#?�j>�(�>aE��9��m�E�<��>u��>�H?��~?��?�Թ�|Z3�����桿��[��:N>��x?�U?�ʕ>7���Ӄ��seE�3DI�������?Ctg?T彂?K2�?�??�A?�(f>���ؾԪ����>��?���\%K��Y��C�	��>���>:	?�����;�&�g�3�>��2�	?�@?�g
?z��D�vx����<.S�<z�Z<گq�JF�<Em[>yv>j�=��=>��<:o�=ؠ��63�q��M<_}v>N_�=�+�� C�$<,?ĨG�N݃��=�r�*xD��>NOL>0��ܩ^?�j=���{����Hx���U�X �?-��?8j�?�	����h��#=?��?�	?��>M��~޾����Ow�Bzx�9u���>`��>�tl��	�t���L���1F��ƽt�5�m4�>B�)=pb�>l�>�1_>�X�>U�e�¦� Ⱦr����d�.bK����|� o1��푾��k�=�l�������T>���ϰ�>�?��~>��>��>�4L��O>>D�>�R=PpH>y��=�+d>Hrp>���<�		��)R?�����\'�#�羘���Q6B?�?d?��>X�`��L�����D�?_=�?���?��u>��h� �+�?L��>W
��o
?;Z?=;� �.)�<�V��V��ᆽ^k
��7�>5ӽ��9���L�U�d��i
?6�?����3˾ސѽ�5��Ҥ�=Ѯ�?Yr)?K�(���P�r�q���X���R�w����f��D��m#���o����s��H����(��38=�7)?�9�?����ue���kj��9A�D�U>�4�>f@�>&`�>��S>*��2�z�^���$�#j����>�:{?�[�>�CJ?�lD?r�k?:	Y?Vb�>�"�>�����>��K=��>��>o*@?��0?0?��>T{?��>�a��-��m�Ӿ�?I�$?��?`��>�h?�4�I�
��`�<v��;���pn���s>TU��R
b����;�I'=�>�t?���8�������n>�#1?��>��>����'�y���_<���>M��>zj�>v���d�n����#�>6#�?'���<N#(>?�=n�ܻ�������=H��d}=�� ��_�4<��=g=K�6��^�;:�w<� ���c<%?^�.?d�>
�> 畾
���u�.v�<��>���>�#�>���'|�ٸ����m��ޏ>w��?�h�?���= ��= 3�=��'���쾃���.Z����>'?8U`?��?R;?��?�s=�+�U����_v��}���K%?�E??U�>e%���|��޳���4���/?��>�N8�X�x�"}����1�I��G�>��c�B_��=���=w�=�<>�(�������?��?U�%��h��u��k�����p?q$�>��=���>o���X�m���C�en�>�a�>q;;?I>�>ZV?��?�u�?�F�>���R}��������o�W��=E�[?�Tp?��?�e?�x�>�,!=�5j���þ�B�N�#�OL'�����=_a>ˊ>ȼ�>�h�>`">���m���CcA��D>�S�>��>e�>r��>�[>jZ�O�E?C��>�����	�L㧾�Cz�ƣr��Qn?�(�?��0?D�|=���@��x��Ż>[��?��?�`.?��;�3R�=CVݼ����m��p��>�#�>w��>�И=���=��.>UO�>�*�>5_&������?������?LE?#z�={#����^���;l���w���H�����P�f�K�z�*=r5���/�s5��J�T!���೾z|�^C��ʏ,��&�>�}=���=vZ�=��U<ĽF�<� >w�<�<9}���D<�.�����1�����=,�7=��r^j��N˾_U}?I?.b+?
�C?�_y>��>�32���>Ḱ��%?�V>��Q��k���<;�����X%��|ؾ6C׾s�c�tƟ��>}J��$>w3>�l�=iV�<�W�= cq=䍎=e"`�G|=i��=\̹=B�=�6�==>y\>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>s��=x�2�T��>��J>���K��A����4�?��@��??�ዿТϿ6a/>=�C>��=^�8�y�S��Tl�z��F<�`[?�H�Y�K�˅��$�o>�9��@$�Q����>��_>����>�O��=N�a��>R#|�IN> ���K=|}�=���;�ё=�*e��ID>e�.=�Ty�k�⼗;>u�!>+�=�0=_]�>��4?�N?��?N��>Sb����پ� ��j��>��>w�?�a>;j�>v��>�k;?|K?MC?FF�>IT=☚>���>�7�������*���Z�߽F�,<Q?�B�?Y�?�u�=J�$>iE�N���	�8��&-?�*o?/�,?�>P������!���Z�� ���F=��=�Q���7����v�ҽ�� �:H��! >�׷>Ѡ`>p~�>��4>4�g>�s�>���=�G��<�ؽw���-�=��H=[7��1]�>�6=Os��J�q�ˌ,<�Rּ\��wBp<߈b=�=1��=d��>%`>e��>c��=�W��1�<>�2����I����=�"���:G�e�f��Zz��0-���8�)(>>E*Y>��0������ ?�fU>W�>>w9�?��p?MU->Zd�%!߾'�(iK�w:����=P��=�D���8�˰[�A�L��ھ���>���>�G�>j��>����H�~߲>gm��$1��a?���t4������1������U���`�J�)��3)?���������?�?be�?�\H?�T2��-����>�HJ��.�4.��ٔ���WK?�?��Y=��=�Q>�L̾����j��>��H�5�O�H���z*0���)�ष��4�>���Ѿ�3��4��Zߏ���B���q���>L�O?�Ǯ?]ub�P>��O�U��?惽C|?n�g?�]�>��?��?
x���Z��������=��n?��?i�?c2>x8�=�f��r'?�c�>+ݤ? `�?�?QFq��K+?Ɲ���/'>E��;ْ>�o5=|�[>���=��	>��G?6a?���V�x�����)���~�=f�̼��,>l>$����@����=rQ>���>IV
?)��>�h>���>`ׅ>�􉾂(�oP ?�,�=�c�>wKV?�i�=v�<"@�=�I>i�]��䖾'�5�� >�$#>�^
�җ-�ON{>��5>��>�)ڿ�6�?�)i>$�CC?��I$>j��<��>��;���>U�>TM>�p�>���> F�>�4u>W�/>�ػ�>(>,[4��<	�iJ���N�[[��'�=���Qk��*	�Oj`�5-���U9��8�:�j��]v�G�:�S,F��o�?���~'F�~��\��;;t"?���>{��>����l���b>��>m�=�_Ⱦ#T{��*������u��?���?�7c>��>1�W?�?B�1�D3��rZ�ߩu�,&A��e�Ի`���������=�
�2���8�_?��x?]wA?%��<7z>F��?��%��ӏ�'�>�/��#;��<=U,�>�'��Y�`�u�Ӿ��þ+8��DF>�o?
$�?CW?�OV��
H��>�=?"�,?��r?X6?F3?�h�Lr%?`J>2?��?Y�6?.C#?�U?��W>�o�=a��<#v�=QД����l���J[L�߭=�X�=ύ;/��.�<~�*<x�����Я><��t���<_�e=�@�=��=�>�]a?�$?�&H>�'?
%��=�S�D�ھ+�o?�ô>�->�N<�=��3�z-��e?S4�? 	k??��>R�H���W���2>%�h>�ˮ>jG�>q�0>_�*�:�����=6� >�x�=���=7}�9��>�\������jcн�t%>���>�Nz>�2��w�>���p}��c> XB�+���O�8�G�71��}����>�J?��?R��=����{���-d�H5'?�v;?�M?�?`�=�پn�9�6K��%��^�>.6�<�����'����W:�á���r>�ɝ��0C�BJO>6������]Y�o�`�(�\_m>*�G�tS�=;L� ������>_��X�=������<��vߜ��O?�
>.ݾ"���Q�I�>�j�>��>u�=c�*��H��¢���*���>�n>��<�#�������<T�>O�I?`g?�	�?{Og��X�FF�Ǽ��>��JG���?4I�>��?��>D`>�ƾ�$&���T�?��>��?��	��qP��M�ξ �A��VJ=���>v>�>b!?UgS?]�
?}i?M�/?3�>�?>����Qh˾�&&?���?��[=�`ؽ�?[���8�0E�¡�>:[%?�B�ѡ�>�R?��? 0%?��Q?x?P�>�=��[A���>�a�>��V����L�V>!M?ST�>_]Y?��?Ƥ0>\�4�-Ţ�uֽ����=� >�2?�$?�?=��>G��>L�Ѿl^�>c��>dk?��j?�xO?62N��j?���<���>�~>��>��*=Ȭ�>��w?Əo?qz�?�3?��:=ߘ�;�7U�SZv�=�����;6�>˚*>�x��z[<� ���$�MI�=��s=5F2�(����ǽaVF��o{<Z	�>�r>���4+>'�ľ����?dB>?�>�=Y���4��N=���=djz>�?�Ȗ>>1$�Q��=�*�>�/�>�W���'?�[?i?Gh&:��b��ؾ*�H����>�XA?*��=��m�L���:[t�6�[=��m?�&]?QAU�������b?U�]?�l�=���þ��b�v��;�O?��
?0�G���>��~?��q?v��>,�e��:n�C���Db�{�j���=�s�>_Y���d��6�> �7?�S�>��b>�N�==z۾;�w�9s���?P�?$ �?���?_8*>��n��2࿎�����WM]?�x�>����;{(?`�=����zf\��o���ľ$�������x�=�⭛�4+�Ml��j��¯�=s�?bM�?��r?��_?�2�(�f��T�{�v�JQ���
���)��:��\>�m7�TVS����[������R�;��l���K����?Y�+?9�8��u�>�]�Lپ�����!>��P�5�� �=e/�<��D=B��=�S�8��Uƕ��"?���>���>��@?�N��4?��P(�:�,��S��*"�=_>�:�>�J�>��<���L0�&�ؾ|ĥ�"/�e_z>�zb?(I?�Ko?�{��2�|c��A� ���Z�量f.A>��>�ۆ>��Z��)(�&&��?���q�p������"g�=G�0?�qu>�Ǚ>TG�?��?kO
�2"��8�u�
r1�I4<���>�lf?���>`��>��׽O� ��<�>.e?���>�e�>�rD�r<)���~��i�����>/��>�F?��x>�ҽ�,[������o����0���>�\?�b��Z��i�> =5?n��k�:��f�>����"���;��s{,>���>9	�=J�1>�|�� }��s�놎��)?ƴ?Yy���(+�E�|>M!?��>��>��?�h�>b�¾1>��XJ? k^?�fJ?7@?�
�>��=S��@}Ƚ�j&�<n#=8��>%�Z>˥^=�\�=����Y����:UE=$�=����U��4�<Z�����[<3�<�}6>zI῭aL���� �{��2}�&X^��^��x���&�� 	��Uƀ�A�\�y-x�z��MVD��S��,����?���?����Y��ڊ�$����>|��_? ꏾ�;k�|���XѾ�����7�&vP��Gp��R���:t�O�'?�����ǿ񰡿�:ܾ3! ?�A ?7�y?��7�"���8�� ><C�<-����뾭����οC�����^?���>��/��p��>ܥ�>�X>�Hq>����螾�1�<��?7�-?��>��r�0�ɿb����¤<���?/�@��??ʿ)�<��=�p=���>E�	?�:>v�2�p��G������>��?-��?J.=8�T�n����f?K}�<)B�^��t��=n[�=�3=c��-M>�H�>Ճ�l�H�$A潹�.>��>�x	�93!��e�K��<�~V>O�齉���Ą?j1\�f���/�#H���~>8�T?1�>iX�=��,?
'H�eϿo�\�z#a?��?�m�?J�(?g���/��>��ܾ�kM?6?�9�>M&�l�t�<(�=p��N��9��[�U��x�=�n�>��>Z-��%��-Q�!D��[�=���=�ƿi$��� ��\<�H��"9~�2��w���?Y�׌����g��ѽ��^=z��=�-^>t%�>��Z>۟[>RZ?�vq?]�>�j>���Q�����)�<u�B�'�A��� /D����<�N�����6z��e�[�ɾ�V:���=� u�����r11�y�]� $��[1?��=�!��My�>�(��k&�C�־�ؔ�IEX�e�����M��p����?>?�^����6���	�hi<>;;��e�?fZ��WZ@�p���1�>���7��>��>SΏ����f������Bh0?>h?�ľ>Y���> -�#T=��1?�\�>t�j=�)�>K�?λ;�}eս��`>�>�ؙ>.��>��=�V��X�ͽB�?��X?�A��t��b��>�*��Fp���=_�!>5H��
4�"�a>�/��0ӄ��j�ņ���5f=yW?c��>��)�����4��CY�`<=��x?��?ue�>nsk?��B?�ǧ<�h����S���� u=�W?Di?��>����Ͼ�F���5?��e?Q�N>>mh����"�.�.Q�?��n?�>?-��j}�e��;��hF6?�v?v�^��B��Z���T��g�>���>�>�>W�9�0�>�>?�z"���������3���?ː@��?�Q<����Y�=D}?B�>�gO�"�žD����{�l=���>�v����u�p��Y.�<8?
z�?�f�>e�������6>ׯ���'�?���?�����=�Rܾ,�Z�����{��y=f��8�V=�i�����վ�w�iÒ�sWy�� �>x�@�	�<5�>����_Qҿ��׿A΢���ݾ$W����>TX�>D�l�=H�������Fl��A���p�>	�>������e�z��;�*Ƽ>��>^�X�U��>�A]�e���ق��#��;Z��>���>��>�6ѽ&k¾���?��C̿jx��]H�]?���?o�?�>$?u��W7{���~�P�¼�H?}r?��Y?��ɼ�T��[��j?�^��6U`���4��GE�#U>J"3?B�>��-��|=]>N��>�e>�#/�x�ĿFٶ��������?C��?go���>.��?s+?Fj��7��\Z���*�z.�7<A?V2>/���ɹ!�p/=�Ӓ��
?~0?�{�w.�K�_?�a�I�p���-���ƽ�ڡ>��0��c\�lP��V��}Xe����Ay����?*^�?>�?���� #�56%?��>����8ǾP�<i��>(�>�)N>�H_�M�u>����:�Zf	>���?e~�?j?�������V>�}?�>޳�?$��=*��>69�=/Ⲿ�A��!>�C�=�:� ?�LL?.��>�6�=>�]�.���F���Q���q"C��n�>�Va?��K?�Z>�|��_#(�I�!�|�ӽ:�1���ʼ��@��lC��(ڽ��0>��9>��>��E�-Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��3a~���g7���=��7?^0���z>���>��=�nv�λ���s���>�B�?�{�?]��> �l?��o�:�B���1=&M�>��k?�s?T\o����B>��? ������+L��f?�
@|u@p�^?!T���T���z���=�w�^=���=��C>�"�U?~==o�R<$z���=@u
>*0�>�Q�>,�>�>!ʅ>�����#�6�3ݧ��V`���#�Ah��$C��_Ő�˗�����l��_&�������m��lսw_��q�2=[B�=v�U?(,R?Ӣo?�� ?��r���>�����*=$�#�C��=�u�>jm2?��L?��*?��=���}�d���E��^N��?�>_aG>��>�f�>���>�8)�ܨJ>t�@>~�>O`>��*=v�P:QB=S4M>L��>���>H
�> -;>$�>���%���i���u��½���?{Q���N�)��*i��	8¾�͟=��(?]�=I
����Ͽ��VuG?*�� ,�#�A�e�=�7?V�R?��>���[悽��>��콴�x���>�����9d���@�E>Ⱥ?��>��W>��_���J�Q�m��Y��1�n>�9?*2例#���(���f�y2��&.>,�x>�ƾ�޽$'��
1��+-�>�<??T|	?��v�� �����<n�,�>ƣ�=�L���-�>8+� �S=�o��M�C�*>^�}>L�?��+>$�=W��>����D���ǒ>%LH>#�=��;?Qq?XȽb|�����g�6iP>�7�>pW>>��=,p0����=���>V�n>=�����q���ȽG�m�V >?ս�k2�C*T�yĽ��Ό��@<=k�=�Խ�L�V<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>zx��Z�������u�d�#=Q��>�8H?�V����O�g>��v
?�?�^�੤���ȿ6|v����>W�?���?g�m��A���@����>:��?�gY?poi>�g۾=`Z����>һ@?�R?�>�9���'���?�޶?կ�?�[>�E�?��t?�O�>���;�o'��/������Q�2>���=���>_�z>:|��~�J�[�������6V�I���$�>Yy6=�0�>��དྷ7���Ǩ<ߟȽ~���G�k�#x�>\[[>'JC>8��>a��>�d�>�>��X=���t���0d��
�K?Kx�?���C�n�b°</�=��_���?�|3?�8Q�Tо�.�>A�[?�w�?t	[?�/�>sZ�����3п�8%����<skK>F!�>���>'��*�L>�Ծ�[D�7��>�P�>�����6ھ�P��}�v�wڜ>8!?_(�>ò=(t ?��#?�#m>D�>��C�ϑ�y�F�JE�>���>�?�g?^�?����3�,]��%����PZ�^�Q>	�y?? �>P-��#0���s��S�2���>n�? mg?����?�m�?l/??��@?��e>�#��ؾ[l���؁>�j"?�⽍�=�V=�K�L�O��>]��>$8?&�����S��|������?|^\?�G?�־��R�"�߾+�<`k�go2�Ӑ;=������=}(N>�H <��=�e>�^�=�w�?�L��?{=X��=��>��>�G��>0=G/,?��H�W�X|�=ӧr�ΈD���>`2M>������^?u}=�?�{������Y��9^T����?2��?{Y�?�v��h�h��=?g�?�P?@��>
a��Ԅ޾��ྉKw�x��S��>�x�>�Bz��6�s��)����7����Ž��a�?H�> �?��>��4��F?30^��{3�I�ؾ	}��._j�&�?.�5�n���%u�ý;�=�ڗ?tLp�\�>�O/?
ǃ>*� >�~?H�� �>�V>]/Z>��>�ɥ>��>+��=Sh�<׈_=�"R?���ct'��#�;Ű�dPB?��d?�-�>��e� ����u��8?u�?��?��u>T5h�T�*��`?M�>�z�u}
?d]<=����0H�<�����
��Q���#���>��ٽ�!:��M��e�gz
?_�?Г��#;�=׽&����|z=x*�?�t+?@8&���S���m���T�K�T�T��e��9���#��"p�s|���*��� ����'�vB	=�['?��?�s���\龽���b?h�t:���M>���>� �>G�>m�@>Zm�",���]��w(��c}�7p�>�jt?q�>��=?Y4P?��P?]�a?CG�>��M>�Rվl�?��v>G�>��?�/?,?��%?�?m?�ľ>Bܝ<���D����>Q�?6�?)� ?R.?|.���ʽ%�<t�'��ܴ�,�N�t�潴��&�����="92>�ǭ=ʅ?�����7�DD���qm>'54?S��>��>�򑾧R}�(̶<��>��
?Î�>�8���q�����'�>�6�?1��b�=m'>���=�1h��-�D�=�F漄��=��K<5� �n<��=Ŵ�=ػq��:qJ�;i�;l\�<��>�Z%?��>$�>s���־�.%��<�o�>�r�>C��>���>e��6�u�u-_>l��?[��?qxK>��>Uy5>�g���Ͼ�YT�b!Ͼt;:���>u�??N�M?�e�?d6M?E�?C�i<��*�� ��3:�!���Ѱ'?DR?�Z�>=H)�f@��:���o���?��?��g�+�I��]E�J��Zm$�a���9
���o�8���v�S���%�9�u=��~��?Җ�?F"�>wK,����>�j�5��S-?%B?At�=@V?��1���K���ȾtV��h�>�}J?��>�mu?�֎?6�F?���>*�H��J��S���~�>:��>5[?V��?� �?u��?�?y=1=����Gݽ_
���6M���
�H��ؑ=���>%�>��>�v�>e��=��>�>�ﷺ��d�N�l=-�>��>S&�>Ǣ>lƂ=�GG?��>�������cA���#��t�4�FTu?�\�?��+?>�=�D���E�I���+�>Zۧ?��?~;*?�MN�.�=��׼B����g���>��>6�>���=�D=�L>���>�Z�>X.�:��8��0��r?qSE?�t�=@���k��#t��B����k< ���]xl���=�����2(�=Wᔾ��$�nS���:v���(ş�������o����>�z=��>���=��w<�����D���b=��;�h=
[+���=l<����h�wmb�K���d��;k~g=��л-]˾
v}?�#I?��+?��C?1/y>f>)j2�g�>�L-?7�U>�O�n����{;�߷���_����ؾk׾��c�0̟�(>x�H�V�>�X3>\�=�P�<~^�=Dr=�V�=cL�.r=6��=��=	-�=M�=7�>�=>�6w?X�������4Q��Z罥�:?�8�>g{�=��ƾq@?�>>�2������yb��-?���?�T�?>�??ti��d�>M���㎽�q�=K����=2>s��=v�2�T��>��J>���K��B����4�?��@��??�ዿТϿ6a/>ֽ�>�X>��Z� 9W��f��.���Z��V�:?�9���e����ҽy��C�	����1r����>h!��Q�����>�*�c.�=�Wl�b,�=�>��;dV�0��=�)>[�>J�>pq���)����_�<�~�=�|>M��=���>Z=?� ;?)lg?���>*� ľ/�վ��>��G>r��>6�=Iv{>�Ӭ>�T"?2�I?�P?G��>l�>k��>�K�>�,!��+_��{���㥾�V��s�?Ŋ�?���>F7~=��=�����A��KO����>�1?ߐ?��>Yy�� �hy�4=�#�F��e#���.<`�����潓*�=`㓽�f>��p�=ش>B�>3��>���=��K>�?m>�
�>0$�=	w�<B`K>�ߎ>2�=�f"�[��=��=i�S��:���6�M���d=1����ʭ=YC>�[W=/Sƽ]��=���>�>Ar�>���=졵�Us/>X3��+M����=������B�l�c���}�c:/��6��q>>e'V>'Oؑ�z�?F�[>;?>��?ˡt?�� >00�	�־�	���c�ĘR����=��>[U=�d�:��*`�I�M��Ҿ��>�#�>L��>3!�>��0�HQ�'q�>(IԾ��I�G�>�p���D�V}	�ya�w{���>���N���c��Of?������=�W�?Rf?8p�?F�?��=�f��پ�>�����!�= _�&Z꽱\ɽ��/?�HJ?���>p�������C̾��a۷>�5I��O���ʯ0����з����>[�����о�"3�xg������"�B��Sr�E�>h�O?A�?l5b��V���SO�2���#��q?�xg?��>sI?@A?&���}�9o���j�=��n?���?v;�?C�
>���=dM��x?Ln�>�՘?��?a�Y?U䇾�M?Ѭ;y~�>Ix��N�>�K�=�QA>P�>�>|\#?��8?P��<@��ǂ���j���R�&��mJ��Ln�s�M>f+�=�G��A&�=�y�=��>f�>6��>�>IH�>%0�>Tݣ�y��š4?�/�=��f>UD?�Ҍ>�N̽�y>]�|��� >(���=e�=*9���7=��C=��>U!='��>ڿ�pQ?{��>-`6���?-͡�+�">��D>;�U=�����>�v�=�,�>ޯ>�]>��>�Q�>�)�>@Ӿg>����;!��C��R�Z�ѾC�z>����E	&�����	����H�C����]�Zj��'��%G=�і�<~;�?²��6�k�;)������?�>�6?����#[���>k��>;��>�?��.{������#bᾮ�?���?�<c>��>�W?3�?�1� 3��sZ���u��"A�e���`�xߍ������
�o鿽0�_?,�x?�{A?z�<3z>���?g�%��Џ�3'�>�/�c';��&<=�!�>x+��0�`�+�Ӿ�þ�M��FF>ʘo?&&�?�[?�ZV�Pv���y>�m;?�!6?���?��4?Ӡ*?�f�^�5?mey>}?3�?|-?��?8w?L�>�/�=���=Ȓ>�/��/������o�ѻA>F<���=��>k���4������Q����=���kϼ)ʽ�R.;�N�=!6j=ڤ�=BK�>':U?���>�%�>�F=?�W�r�8�QG��m�0?C�p=�4Z��kr����/9��2��=r�m?Fޫ?=`?��>�R<�iB:�,�,>>��>P>��V>��>�Ľ��G��Sb=��>�=0>��=㘵�ԥ���	�ش���	�;��>F*�>�Vx>;Rս�I>>魪�Dż��vQ>�P��o
þ%(����@�qlM�l]7��մ>�??J)?�\�zMܾ$����PU���?_ ;?]&d?ATw?�d:=���=K�<M[��9&����>�;�d���b��fE���2����	1>Pu��M�����k>s9��Ɩ��≿�_g���<� >��'�I��(!��w�5�~�d*=>"Cn=ꐲ�C���1������Y�S?��
>�3�B9��J��'�3>�ڳ>�{">	��=Z��L�W'�ka��?D�=�m�T|����ҍ��m�>E�C?��X?��?�}E��,w��6���|���W�����?�A�>�(?$�a>&�>����!w�]�`��D�gX�>���>��R�7�l���g���͛�'�0>�)
?w�>�4�>^LG?�S?Bh?��/?��?FI�>#,.�����U%?��?@�\=X~��vtp�9%=� >����>x#?XB��_�>Y?��?��)?�*W?v[?��=����C����>{�>��\�N%���1>�%O?�޿>�P?"��?Z�5>P�>�Ͻ���Cʽ�X�=�I>br*?�>%?#%?[բ>���>��pɇ>��>>p4?Թz?���>Q=N�?�ؾ�f�>���>.i!?��y��M;?�D�?��?�yK?�?��=�G��r�Ȯ۽�V}�Fü�]�<"`�=������rr���0�=Lu��^���߼hh��E�<�[�<C<��>��l>>7��5�'>�Eþ�䓾4�8>�»t����x��}H����=�vY>I ?W�>�%�ۡ�=gɸ>��>� ��x(?�#?|y?�U�8�\���پb�,����>�QC?W��=��q�5�����n�U�{=�Yn?S�V?x�C�ܭ�U�b?��]?Nf�<=���þ��b�Ȇ���O?Z�
?�G��>��~?p�q?���>�e�z5n����=Fb���j�M�=�p�>�Y��d�2�>Ԟ7?
V�>*�b>})�=�r۾��w��l��*?���?� �?r��?!+*>@�n�3࿅�־���N�a?qX�>^g��ؘ5?��a��������^Am���Ӿ"�ھq��Xi��z��t�[��T��?�G���f=
�?�L�?!Wx?��m?��6�x�+=���z�/ia�B!���%���6��'U�F�V�	@z�V�ob��Ǿ������R�@W�4��?N?��?�}���������l�>ǭ���Jm��]->wc'=.X>K䃼�ڑ�ƢO�����C!?�q�>���>8�F?Rkf���9�H��?�����-�=���>i(Z>f��>9�Խ%�z��6нy�Ⱦ'���7�r�*��>�e?#�M?ة�?i�o=������S@��%u��?��	��>��q>ʮ�>����c��_�"��!M���E���㾥 ������N�GyP?��>&�h>���?�c/?z���x���yM��"S�)*�<C�?6J?8X�>;2,>���<�T�p��>�u?��?g�>Z㲽����&���Jc�z�?��?8.:?�\�>�ٽ�6t������l����Ƃ5>*�w?�B֍�-�>'^?�w�=�L�=��>�� ��?����w���go=�^	?J�>K�>��)�#��T�vu��{�"?�+
?�՝��0*��Ae>�[?��>~~�>u��?<ڣ>�ξ��l�:�>9wZ?G�E?�<?æ�>�:=&:?��ý��~�=��t>��_>�ѭ=�F>���׳n���C���i=�r�=������ݽ+�.��{�ƾ�<���<'�4>��࿡�S�q\ݾ� �%��ES	�d�=�1� ����@'&�D���ճ������Z���T�u�%|D� ���F�����?4P�?z.�U�D�9��� u�tǾx��>�肾�a��=4���{��L��˖��:蹾�d/�q:=�S�n��q��!$?!�����ǿ�ҟ�
޾�i?�� ?��s?p�� �_�7���>wb^<��L�W��5ɚ��[Ϳҗ��@�\?���>��������>EȆ>�.m>o>.��9���jg<2�?�Q-?�S�>[ q��Eǿ�0��
C�<e��?��@��A?I'����M[g=^s�>J?�WB>�t3�~��KQ�����>���?i��?��h=�`W�W?�?^c?�M�q�G�3�H��=��=��=�c
�1K>�S�>���i=����� <>�I�>e�>�����a��R�<6�U>ݑӽ��s�5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=c6�쉤�{���&V�y��=[��>c�>,������O��I��W��=�7	�|�ҿ�>+��)�c�<�P޼��9}�U�@S��s��aCI��*��[�ȫ���;&��N�=9�\>1�<>�3>1�c?Қ?�)�>�q�>���E¾)�h��0=N۳�&�}���B�=�k��&W�������r`	�SM��/�KO�{:��U=��K�Y���Њ#��jf��Q�*O=?,���f ;�uJ�iW��8V��L۳���u�̕���o2��|�J�?4`=?���� W�����q%����"S?��ѽ��������2�>��_����=�;�>��9>��ľ�&'�,�P�i#?	�?-���6Mm�P�7>�4������F?�8�>�G���M�>R<?�N��$X��L>�E�>+v�>��>fÎ==±�*=3�{v?py?�(�����b�Z>����9.�)�j=\q�>Ғ>�#�I>-s>z��=�&����^�Žϑ�<� W?H!�>��)�y���%������7=�Jx?�?���>5�k?d�B?@��<H��U�S�l�
���|=��W?^Yi?�f>����b�Ͼ�M��6? �e?�N>�h��H꾥�.�����?Ȟn?�&?a���~A}�H)���
��F6?�v?9Z^��X�����E�V�A[�>)6�>i��>��9�ڲ>�>?ު"�H'�������-4��ʞ?	�@���?��F<q^��h�=}R?�'�>�O��3ƾ�Ǵ�����\p=TL�>�E���(v�ڶ�96,�!z8?	��?U��>N���ˠ�k�B>y�#����?�?�����=�,�vS�GC��(�b�ޛ���J�N\&=��þ��)��=�?��n��+҄��R>�o@$K�=$^�>󜚽[��Ўп_\����վF��?4[?�W�+�)��Y�J�ȭ,�;-|�+��p��>��>w)������{��<��������>[�v#�>N5W��$��vy��3R�<y@�>O�>.B�>rº�Z&����?9����EͿ|J��&��Y?�)�?*ʄ?Ѓ?>{ <b~���z�(G�!�F?]�p?O/X?:�_��ZE�ҿj?V��gS`�ˊ4��LE��U>@%3?�<�>�-��|=�>j��>3X>�/�8�Ŀ�ض�����=��?��?[n꾱��> ��?<q+?Ij�F6��tS���*��OG�qAA?h2><�����!��+=�}ؒ��
?{�0?*{��-��_?��a���p���-�w�ƽ�١>H�0��d\��P��T��Xe�����>y�k��?5^�?K�?��#��5%?�>	����8Ǿv�<X�>�)�>�+N>;P_���u>�'�:�i	>t��?�~�?�j?��������S>h�}?�G�>j�?��=���>���=����n,�R\#>�n�=i>��?�dM?�7�>��=�y8��/��MF�ZR�w��C�X�>��a?��L?�^b>Y;��QO.��� ��ͽ��0���޼��@��+�v!޽�74>Y>>J�>'�D�.�Ҿ��?:e���ؿsM���{'��&4?��>�?����t�k7�Z�^?Ã�>U����(�����z��?�.�?(�?	�׾79мr�>�֭>AC�>c�ӽ7���B8���7>KB?��WL���o����>���?̭@m��?c�h�]	?���P���`~���� 7�5��=��7?,0�i�z>���>��=�ov�����1�s�M��>|B�?@{�?n��>Ȯl?1�o�-�B�=�1=�L�>�k?�s?�n��%�B>�?G�������K��f?��
@Zu@{�^?c�ٿ^��������l�_�c=v��=�<�=�!��ѐ=P�������~�<� >�`>[�{>�[s>!�)>�z�>��>6���;�'������Ș�3+�(:�u�
�}��"��������WJþ,��Խf���*�z}-���P��&$���=��U?a�R?^,r?��?i�v��>�p�����</���ߒ=�z�>#�2?�M?
�*?jԆ=���c�ʻ���y������K��>�N>2��>�}�>�s�>�I;��F>`�@>/�>.��=��)=\�;�{�<"�T>�,�>���>>��>�(>��'>7������`s��m��X�����??����?C�c�����������=��?ɳ�=Z���Qo̿�^��:�G?���<&�8�ؽ�&>�v-?"�D?��=�w���#6��|">`ǽ&hn��>b`��ԅ��"�FU>ԥ?�-h>I>A�K�S�5��6�d��i�>/�D?�˾􀜽�}��������US�>f�.>�S��&9��ϖ���a��Y��S��=�c+?Z�>=�f��R���|2����$>,P�>�s>hֺ���>d�=Ӓ�==߽�䋾M}.>*+�>n��>�+>�L�<?C�>7����׈��D�>�o>�5>�:?�?�\V��������C��A�v>?��>�Qr>��>J����=���>�it>=5����i���� �vff>����	9� ���r/�=��g�/�>v��=M���F/�I�\=O�}?굧�ˇ�VU�$����E?E�
?9�=��<������ %�����?d�@[��?�	���V���?V�?x���b�=�|�>}U�>x�о��K��s?�����"��K�	��!�(�?�O�? {B�	�����j�!�>�=$?�t־�[�>�v��[��=����u�ͭ#=а�>B1H?�R���O��>�4i
?�?iS�ߤ����ȿZvv����>	�?K�?��m��<���@���>���?�eY?�ni>*_۾�~Z����>�@?��Q? �>�:��'���?�ڶ?���?:�~>RB�?^��?.��>Ԥ�<n<�r�οQ���+K��е�C��>w��>��Z��TL�λ��&T���}�: ����>�c�<0Ө>�IH�7����p>	6;�}��Bl�����>�R�=���>���>�a$?�b�>u�>���=�}i=�vC�p��OL?G��?��oum����<8�=�/]��?@4?f�t���о��>%W\?�ˀ?�vZ?�	�>I��Pk��t��a���0֔<��J>�>���>�����J>�"վm�B�i�>AZ�>�㣼�0۾1���|E�Y �>� ?��>�K�=˙ ?ɜ#?�j>�(�>aE��9��m�E�<��>u��>�H?��~?��?�Թ�|Z3�����桿��[��:N>��x?�U?�ʕ>7���Ӄ��seE�3DI�������?Ctg?T彂?K2�?�??�A?�(f>���ؾԪ����>��?���\%K��Y��C�	��>���>:	?�����;�&�g�3�>��2�	?�@?�g
?z��D�vx����<.S�<z�Z<گq�JF�<Em[>yv>j�=��=>��<:o�=ؠ��63�q��M<_}v>N_�=�+�� C�$<,?ĨG�N݃��=�r�*xD��>NOL>0��ܩ^?�j=���{����Hx���U�X �?-��?8j�?�	����h��#=?��?�	?��>M��~޾����Ow�Bzx�9u���>`��>�tl��	�t���L���1F��ƽt�5�m4�>B�)=pb�>l�>�1_>�X�>U�e�¦� Ⱦr����d�.bK����|� o1��푾��k�=�l�������T>���ϰ�>�?��~>��>��>�4L��O>>D�>�R=PpH>y��=�+d>Hrp>���<�		��)R?�����\'�#�羘���Q6B?�?d?��>X�`��L�����D�?_=�?���?��u>��h� �+�?L��>W
��o
?;Z?=;� �.)�<�V��V��ᆽ^k
��7�>5ӽ��9���L�U�d��i
?6�?����3˾ސѽ�5��Ҥ�=Ѯ�?Yr)?K�(���P�r�q���X���R�w����f��D��m#���o����s��H����(��38=�7)?�9�?����ue���kj��9A�D�U>�4�>f@�>&`�>��S>*��2�z�^���$�#j����>�:{?�[�>�CJ?�lD?r�k?:	Y?Vb�>�"�>�����>��K=��>��>o*@?��0?0?��>T{?��>�a��-��m�Ӿ�?I�$?��?`��>�h?�4�I�
��`�<v��;���pn���s>TU��R
b����;�I'=�>�t?���8�������n>�#1?��>��>����'�y���_<���>M��>zj�>v���d�n����#�>6#�?'���<N#(>?�=n�ܻ�������=H��d}=�� ��_�4<��=g=K�6��^�;:�w<� ���c<%?^�.?d�>
�> 畾
���u�.v�<��>���>�#�>���'|�ٸ����m��ޏ>w��?�h�?���= ��= 3�=��'���쾃���.Z����>'?8U`?��?R;?��?�s=�+�U����_v��}���K%?�E??U�>e%���|��޳���4���/?��>�N8�X�x�"}����1�I��G�>��c�B_��=���=w�=�<>�(�������?��?U�%��h��u��k�����p?q$�>��=���>o���X�m���C�en�>�a�>q;;?I>�>ZV?��?�u�?�F�>���R}��������o�W��=E�[?�Tp?��?�e?�x�>�,!=�5j���þ�B�N�#�OL'�����=_a>ˊ>ȼ�>�h�>`">���m���CcA��D>�S�>��>e�>r��>�[>jZ�O�E?C��>�����	�L㧾�Cz�ƣr��Qn?�(�?��0?D�|=���@��x��Ż>[��?��?�`.?��;�3R�=CVݼ����m��p��>�#�>w��>�И=���=��.>UO�>�*�>5_&������?������?LE?#z�={#����^���;l���w���H�����P�f�K�z�*=r5���/�s5��J�T!���೾z|�^C��ʏ,��&�>�}=���=vZ�=��U<ĽF�<� >w�<�<9}���D<�.�����1�����=,�7=��r^j��N˾_U}?I?.b+?
�C?�_y>��>�32���>Ḱ��%?�V>��Q��k���<;�����X%��|ؾ6C׾s�c�tƟ��>}J��$>w3>�l�=iV�<�W�= cq=䍎=e"`�G|=i��=\̹=B�=�6�==>y\>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>s��=x�2�T��>��J>���K��A����4�?��@��??�ዿТϿ6a/>=�C>��=^�8�y�S��Tl�z��F<�`[?�H�Y�K�˅��$�o>�9��@$�Q����>��_>����>�O��=N�a��>R#|�IN> ���K=|}�=���;�ё=�*e��ID>e�.=�Ty�k�⼗;>u�!>+�=�0=_]�>��4?�N?��?N��>Sb����پ� ��j��>��>w�?�a>;j�>v��>�k;?|K?MC?FF�>IT=☚>���>�7�������*���Z�߽F�,<Q?�B�?Y�?�u�=J�$>iE�N���	�8��&-?�*o?/�,?�>P������!���Z�� ���F=��=�Q���7����v�ҽ�� �:H��! >�׷>Ѡ`>p~�>��4>4�g>�s�>���=�G��<�ؽw���-�=��H=[7��1]�>�6=Os��J�q�ˌ,<�Rּ\��wBp<߈b=�=1��=d��>%`>e��>c��=�W��1�<>�2����I����=�"���:G�e�f��Zz��0-���8�)(>>E*Y>��0������ ?�fU>W�>>w9�?��p?MU->Zd�%!߾'�(iK�w:����=P��=�D���8�˰[�A�L��ھ���>���>�G�>j��>����H�~߲>gm��$1��a?���t4������1������U���`�J�)��3)?���������?�?be�?�\H?�T2��-����>�HJ��.�4.��ٔ���WK?�?��Y=��=�Q>�L̾����j��>��H�5�O�H���z*0���)�ष��4�>���Ѿ�3��4��Zߏ���B���q���>L�O?�Ǯ?]ub�P>��O�U��?惽C|?n�g?�]�>��?��?
x���Z��������=��n?��?i�?c2>x8�=�f��r'?�c�>+ݤ? `�?�?QFq��K+?Ɲ���/'>E��;ْ>�o5=|�[>���=��	>��G?6a?���V�x�����)���~�=f�̼��,>l>$����@����=rQ>���>IV
?)��>�h>���>`ׅ>�􉾂(�oP ?�,�=�c�>wKV?�i�=v�<"@�=�I>i�]��䖾'�5�� >�$#>�^
�җ-�ON{>��5>��>�)ڿ�6�?�)i>$�CC?��I$>j��<��>��;���>U�>TM>�p�>���> F�>�4u>W�/>�ػ�>(>,[4��<	�iJ���N�[[��'�=���Qk��*	�Oj`�5-���U9��8�:�j��]v�G�:�S,F��o�?���~'F�~��\��;;t"?���>{��>����l���b>��>m�=�_Ⱦ#T{��*������u��?���?�7c>��>1�W?�?B�1�D3��rZ�ߩu�,&A��e�Ի`���������=�
�2���8�_?��x?]wA?%��<7z>F��?��%��ӏ�'�>�/��#;��<=U,�>�'��Y�`�u�Ӿ��þ+8��DF>�o?
$�?CW?�OV��
H��>�=?"�,?��r?X6?F3?�h�Lr%?`J>2?��?Y�6?.C#?�U?��W>�o�=a��<#v�=QД����l���J[L�߭=�X�=ύ;/��.�<~�*<x�����Я><��t���<_�e=�@�=��=�>�]a?�$?�&H>�'?
%��=�S�D�ھ+�o?�ô>�->�N<�=��3�z-��e?S4�? 	k??��>R�H���W���2>%�h>�ˮ>jG�>q�0>_�*�:�����=6� >�x�=���=7}�9��>�\������jcн�t%>���>�Nz>�2��w�>���p}��c> XB�+���O�8�G�71��}����>�J?��?R��=����{���-d�H5'?�v;?�M?�?`�=�پn�9�6K��%��^�>.6�<�����'����W:�á���r>�ɝ���k���Z>����*�t�3J�_�ܾ��>��W�;����+��I���� �<Wd�=���k~�Q���y�����C?�!�<�v�]��Z`���=ǒ�>-��>��½~��<�+B��׾O5>���>�(X>r�����h][�I��#P�>rLU?��k?h��?��K��/f�a�M�����Q��hS5��?�&�>%�?jL>���==���R0��k���9�
��>UP?���E��?��"r����"����>� �>��=6]?L�g?Y�!?fH?I�,?
�?��k>���`N���,?E܇?,��=�P��v��C�'��"����>�k?���cuL>z�>)= ?�1<?�1U?�d?g&;>�׾�Q0��><��>�5Y�:͹��&>��[?�a�>�O\?Ä?��=��I�*����U��-�=y�(>��!?� ?�h?���>nU?@����K>k��>�p?1܂?�Y?�p���>��>S��>��0���H>�ۀ>5?��]?Om?��=?;��>0�>���*k����z=�|��"r��<N��=cd�=U-̽Y�#��;=�<���p%�{m�=K#ƽ�1�u�=؈�����>c�`>g|��l�=�ޯ��Ӿ|u~>���R	���|�B&v����>#y�=���>ٱ8>�;u�g��>ʨ�>1��>�2��˙3?@�?�?	��<2~�HT�������>�T?t�E>��T�몿����)�t>8�?�Z?�g��ԛ �P�b?�]? h��=���þ_�b����`�O?4�
?�G���>��~?e�q?x��>��e�&:n����Cb���j�2Ѷ=\r�>PX�f�d�n?�>{�7?�N�>V�b>�%�=�u۾%�w��q��p?�?�?���?�**>x�n�O4�������F�]?�p�>�����$?}���)Ҿ�j���S��,߾�u�����R���nգ����>ʰֽx��=?��s?L.r?>�a?_��Uic�g`�	�~�lbT�ئ����@^B��C�[�A�{n�v;�X���8���k5=R�l��FB��˱?,>'?9��F@?{F��(/���"���k>mѐ�t�`���=���Q�=��=��N��*��"��O ?v��>L;�>�1I?�Q��[:�2�=�y�0��I�ۑ�=/׫>"J�>rs�>ob<$6E���4�fb�sS������qv>�zc?q�K?g�n?H��1�������!�al-�f#��~�B>�O>Aˉ>h�W����%�S?>���r����v��
�7�}=Z�2?0K�>�ǜ> o�?T?�	��@��(�x�3�1�w!�<Nh�>��h?��>�m�>�ͽ�� ����>j�l?;��>��>r����W!���{���ʽ�,�>U�>F��>��o>��,�� \� i��؃��v9�g��=a�h?������`��ޅ>�R?�M�:�,G<)u�>�v���!���H�'�p�>�}?'��=X�;>�}ž%�q�{�t:���;?y� ?T�󽪱&�6�>i�X?��5?���>��?���>r�-��Pa��GF?��b?��?��?�v�>d&.>p��=�o��⑊�T=¸z>N:k>c>S=V>H��7���'ʽ�'y=[T>��<0�2������o���<Ŷv>d�ݿ�XL�zbؾ��E ���U�D���������x�#=��:��2��&���#��7�I�mqa��	_��;��LXs��?��?Jl���󒾸�����{� ������>h�r������R���s�噛�I�ݾt���Z�!�C�M�K�g�M�_�1�'?����ǿ)����:ܾ�  ?~? ?`�y?����"���8�;� >���<������������ο����'�^?Y��>i������>���>��X>#Mq>$���ݞ�c��<��?d�-?\��>�qr���ɿ����Τ<{��?��@��A?''��\꾂t]=���>?n?�g@>�W+�x��6����>ݐ�?��?EA>=��W� m����e?��;�H�;�o��>�=�?�=܀=)b��H>gד>�D��J��Խu�3>FI�>�.�֕��p_���<d�Y>��ݽD��5Մ?+{\��f���/��T��U>��T?�*�>P:�=��,?X7H�a}Ͽ�\��*a?�0�?���?%�(?;ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�օ�=�6�щ��y���&V�v��=Z��>g�>��,������O�J��V��=��|>ƿ2#?��P#�sΆ�Ȥw�����@ؼi
J�,�)6��V��P#��"�=�jE���%>�-4>��o>���>�??t?8�>�6�=�
�ht�X^���IP�I����e��w���n;��k�&�G��y����������"��F�e�e����]�G��s��}4��~�x:�3�(?+.�>���,���tm7>dF ��W��d<Z��� �7��&
���l�j5�?���>���.�E�E����d>�|7�q�?��O�I��M*>�nJ=��� ��fT>5�>������G�D���0?$~?����F���"&>�m��3�=��*?�x ?�U<���>�	$?�.��V콷'W>/01>Ƨ�>H��>0�>�}���*ݽ��?sS?���_���/�>U��q�w�Ƙ�=>�K>����/(`>;t�<B���]��t����(�<\V?f׊>k*����0����/"���3=/�x?�i?��>�Hk?�+A?�'�<Y���PT���
���s=��W?��h?>G><U{�d�Ͼp{���5?��d?�,P>��l�_8�͘-��M���?Qn?��?�͝��V}������*�7?��v?�n^��q��m����V�)0�>�V�>��>h�9��l�>y�>?�#��H��ǹ���T4����?�@��?��;<�e��==?|Z�>�O�^@ƾѡ��낵�^�q=,&�>����tev�����_,���8?���?���>����
��ʕ$>�4��`�?�Ə?�qҽE��=��%��v��1���i�=��>M��)݅��9����v0��W�/�VȬ�%�7����>3�@�F>���>��j��(߿��ԿDK��fV���K��Ż?�$?-�R>	����I�)5a�7�{�qW�3&��Jh�>ol,>|N���6���r�Qz8���/�˳�>��l��6�>|]`��ڲ��Ҡ�e	�<��>���>��>�v��rv¾� �?}���ʿ ^����	�B�Z?�?'�?YA?;�%�=u���Do�NCF<'�C?֬i?�3Q?]ۃ�k�Y����Dj?`I���?`��z4�x+E���T>�13?P5�>�X-���z=&B>���>.�>�.��xĿ�궿 4��#�?jl�?�T�*��>Nb�?�Y+?�+��M���{����*�0R�9,A?v1>�����!��+=��˒���
?�t0?S���=�i�_?0ua�}�p�N�-��Yƽ��>'M0�$@\��+���z��be������x�h��?�V�?F�?�v���"��0%?��>�����EǾj7�<Oi�>Ag�>WN>S^���u>��$;�\`	>���?�o�?f[?z���9����A>�}?��>o�?�G�=�X�>�K�=oﰾV1-�kj#>4�=#?��?��M?�H�>�s�=�9�D!/� ZF�*ER����C���>��a?�~L?ZFb>���72��!��yͽ�e1�g�� L@�C�,��߽�35>�=>�>Q�D��
Ӿ��?Ti�>�ؿ�c��$v'�"%4?�̃>Z�?����t�$��0D_?�x�>�%�E(��+������?/=�?��?Q�׾l�˼�>��>�>�Vս�m��k��J�7>j�B?v���H����o��
�>�?��@�Ѯ?�i���?)�UT���a~����7��[�=��7?*L��z>��>��=nv������s�~��>P6�?u�??��>��l?x�o�_�B���2=h8�>��k?�c?�a�����B>��? ������4P�1f?��
@�n@�^?+뢿��ۿQ县T��}�����i;����k�=v����!>N��=�}.�;dX�
�>��b>9̷=,�C>�dA>�X>���=�b���@��砿�����P��@���"��9���ݾb>��:��kzj��	�w<н>�� �,�]�h�a�V����>��=׭U?�R?&p?ė ?�hx�[�>����;�=�*#�QǄ='�>An2?n�L?|�*?�1�={�����d�FX���I�������z�>0;I>̞�>_�>�>�>�v9�I>&:?>>�>�T'=�����	=F�N>�p�>)��>���>H<>L>˴�1+���h�9w�/�̽O�?閝��J����>#���ͷ�7j�=�J.?�>����+п����5H?#���*���+���>��0?�HW?�>�S����T�a�>�����j��<>! ��Ol��)��!Q>M?wɇ>��k>'�,�{d0�b�Z����!�j>��:?i�Ӿ>�<�l�rC���徒�>�n�>#��<�+�=���	��Δ]�tC=WvA?��?��������J��I��JIV>_��>�+�1D��3�>�8�s[�]F�K��ᖁ<���>s�	?R�G>���=j0f>N����J���>��=?�>��??�?b�5�ʽ�����]T��@>�?:�>d�R>Kh��Q>�I�>�%>62�����<ts�3���O�>ڐ<^0���U���=l���x²=eSl=@#���[���`���~?�u��ވ���i/���qD?D5?/�=+�G<�~"����M����?-�@�i�?>�	���V���?�>�?���y��=Zp�>���>SξoSL���?��ŽM����	�eB#��P�?P�?/�0�H̋��l��>qX%?�Ӿ�c�>���Z�������u�y�#=ԣ�>�9H?�S��Z�O�}�=��r
?�?#^�⩤���ȿ{v���>��?���?]�m��@���@����>z��?$gY?�^i>Rd۾^UZ����>Y�@?fR?�$�>�8���'��?�ܶ?b��?�IJ>N��?t?���>Fvp���.�a3���Ռ���=};���>a�>�j��֎E��C�����k�3K�'a>�'=G��>���u���aO�=Fߏ�J����a��~�>�go>�J>�̟>��?N�>5_�>$� =�ݍ���������C�K?���?����2n�iT�<q��=o�^�?&?>I4?JM[�s�Ͼ�Ԩ>�\?<?O[?|d�>.��m>��迿�~��K��<��K>�2�>�I�>����HK>��Ծr5D�@p�>�З>{�k?ھ�,�������B�>f!?5��>ծ=� ?��#?h�j>�'�>�`E��9����E����>Z��>I?|�~?g�?kԹ�MZ3�|���桿�[�X=N>��x?�U?jʕ>4���΃���kE��HI�����.��?�tg?%O彯?�1�?�??��A?(f>͇�Wؾ�����>X��>6QV�*~I�g��f�t��>O�?���>s&v�PZ��w�=~�̾�Ծ�?t�?��$?�LϾS�Q�t�R��l�=N�-�bؼ�Ь=�d>g5b>��>m�{=S�=!'>!�
>M���GZZ���� �<�(�>�B>V���Me��7,?GF�؃�gј=��r�P}D���>#9L>�����^?�b=�V�{����w��?�T����?$��?5e�?u?��R�h��#=?��?�?��>�K��Ɖ޾/���(w�Lcx�Pq�\�>���>vn���ۆ��O����K���\ƽ�n!��J?��>�E�>ݛ?�GP>�x�>(���g}'� ����w��}�Z��i���@/���G�i{��߄��+���Q���ѾGĄ�TP�>��ý���>nB?���>��q>#��>3C�Kf�>�Rq>Q2_>s2�>2_�=��n>"g{> �>b(�R?<h����#�v��5����D?��f?�\�>6�!��n��Ò
�8�?F�?�>�?Tg>B�h��*���?ʞ?�:����?V[@=N�:���<J�����c�����G�>x½;g7��K���a��?bq?I��e̾��ͽ�����n=�M�?��(?�)���Q���o�G�W��S����n5h��j��O�$�Ǜp��쏿�^���$��?�(��q*=��*?U�?܌�l��q!���&k��?��bf>O�>g$�>�߾>OuI>z�	���1�	^�M'������Q�>�[{?e�>�P6?E5I?�	�?_K[?(3�>[�>�$Ӿ2��>!�=A'�>��?Z;?�"?�s?܂?>�.?�l�>=��J��=�����>gP?�H?W�	?�:?"���S���+x�=�$߽�+ݾ|��oƓ>�W3�ﲇ����=�S>��f>xU�>�j%�D�$�����$=��/?`?���> �J�3Ծ���M|�>���>���>	��|���5ȾN��>|?sa���Ƅ<U�>^��=g�a�oGf���>X��m��=�}�=m�E��,�=�;>�1>H$�z��9>�h?>j�>���>U�?z�>(g�>ⅾ�T �bc����=�"Y>ŹS>DW>}پ	Y�����ɋg��x>�r�?�w�?�xo=�B�=o�=ZH���z����Lþ���<�m?̢#?�sT?)4�?A=?�E#?��>� �~*��zK�����+@?P=?:�y>�1�&>G�bW���6R�ʎ�>,?�A_������=����
罢=<=���<����������������s���X�?*�?�5�=�l.�a�ᾼ����t��w?�o�=��=s0&?�8��B0�����:��ԑ>F�t?+��>�`�?��?ґ�?!�>�
�,���4��|�=�>a>@?0m�?��?�#???���>���V��k��d����.��	��f�B>w�'>55_>��>K��>�>��<^�i�G:�����j�~=vt�>��>�(?���>ӂ�<y$F?:��>���N��U���T��w�Q�+s?��?%?�� =�x���J��� ����>�˦?�?��"?KEx��s
>c�(��{��{w���>��>T�>N�=E��;���=V��>X�>�
�,%�t�9�$c/�A�	?m'??(�?=D����j�9��-�������䜀�����>��־�n��=>�Q�� �69�*�`��վyzվ�Z�E)�L�>
��=�s�>/�=l��`�=bW�=s�;g�<>��¹���>���븄�LO+>
�w�c<,>յ�S�˾��}?q;I?��+?P�C?�y>�:>*�3���>U����@?fV>؞P�������;�|���� ���ؾ�w׾;�c��ɟ��I>bI�3�>�83>�G�=H�<H�=�s=���=�	R��=A#�=�P�=rg�=���=��>5U>Bw?	v��C���Q���꽈D:?F�>��=�YǾ'�??��>>+���������m�~?��?�$�?6;?&+l�XZ�>�������'�==����0>տ�=��3��`�>�L>���pf��gi��3&�?�r@�_??���Ͽ��/>�D@�	���-�u���<@ԾL�
 ��W�e?��?��.���?3��������a+;�a>s=Y5�;Wh���>~����L�=_�>�Di>���=���=$u���m�= 
>C|ݼ!:���O�=�6!>��q����X��=`��<��V>�#�>��$?6�8?g�{?��>��j�R�K�荸���->k��>�Ig>�����E>���>t�?5�?EOh?Ʋ�>�b�=G�>MO�>"�!��Q���/�RÝ�->��?ܿ}?�Z(>]�	��ā�~m�R���B>���>g?��>لA>3*	���׿��$��a:��,˽�{�<�#�<�@{���#�P���C�����ཹ�/=e��>�j�>�w>�n[>}�V>zgb>AH�>��>�\�=�C=;��<=�U��m�=5��<]��b���ٟ�<��B�ơ]�.�Y=3���[�]<}=�̐<qi�=`Y�>�f>���>�=����/>�U�� �L��^�=�W���RB�,�c���}��
/�҅4��A>�T>�S���=��h�?�`Z>��;>ׯ�?��u?��">����վ���Cb�X�Q��=��>�`@�&�:��'_�6M��BѾ���>p��>C"�>�l>'�+�� ?��x=-�hR5��V�>�����(�����$q�!/��Fӟ�mi�a0�lvD?�L��p8�=O~?�RI?6��?���>sg��3�ؾH�/>� ����=�����p��)����?U
'?^��>�뾕}D��+ܾ>i齛n�>��e�r�O������62�^�<Y������>��̾�4���������� @��!{�a��>>�I?M�?P�{��H��4�G��(��5�g3�>րk?���>A�?{x?�߽D��)������=�o?���?A��?�>�t�>��=� ?���>�Ϟ?F��?��?wї�K��>�0�>�Cr��\�/��>U[�>�C���{=60?Nl?��&?�Ў���������T0��3'
���>��<n�=��>h�9>��j>M4�Q���}'>շ�>��X>���>��<>�
B>;榾��_�%?�Q�=>?�>-�1?3ۂ>?J:=�����=��@��H��.)�����c��l�	=��;�D=b�����>Gƿ���?�bV>��"�?�)��Q2���Q>3+Q>�ڽ�_�>��;>:X~>��>�>��>Vy�>XI+>TK׾��>�k�O�!��{C�R�R���Ҿ�|>>�����*�Qn�%V�]L�h���l,���i�믁���;�|�<�n�?����p�m��U*�������?��>�{6?�$���Ñ���>���>Gӌ>����Rs��,���>���{�?�e�? Bc>]1�>�W?YM?�:1�F�3��*Z���u�Z�@���d��~`�թ��4���$�
��b���_?�!y?�zA?xg�<�:z>\��?��%�װ��}��>w)/��`;�s�;=ܧ>-i��+�`�Ծ ľ����G>!no?8�?5�?�W��Bi��'>C�:?z2?r�t?i	2?g�;?���]$?��4>��?K?�n5?/?h
?��1>��=�a���*=�������2ѽ��ɽg���4=0�=/��9�B�;��=�T�<,��pܼH�~;\��uȥ<��==*�=�S�=0�>�Z?]��>��U>�67?{��c%�
:���x'?�{�=@&��������_���[u=�:h?�?�-K? tm>��B���S��:>;�>��5>�gW>�ۤ>�uý�"�?��=�*�=��>��=�+�����������]���Up=�c>^�>�_�>Lk=-.>d��<o��?9>훾�(��؈�=�S�x�K�q����*u>��.?U;&?v���s=���$��`��K�3?$�A?�p�>!�?���>+����K�^3�����F� ?d��=!¹�6҄�+Ӫ���n�O>��>A�!��cT���e>�C�!�	��Vm�X�@��?ܾ��><� ��eĽJվ~�����IY6<G���8�a���ᑿPݷ��(A?�=r�u��;���ξ��k;�S�>zyN>�f���==f�b��������)?)s�=�s�7S+����H�پ�bs>��a?RB{?���?Ζ��d�P�N��+�𒰾9w�G�?��>�?��\>��,>V����&�R)|�5tD�>I�>*��>BC�Ձ���y�u��j;\��z>�?i�;>1K#?Mm?q+
?*B? �M?^?֥M>F���ܽ�;A&?���?j�='�ԽԿT�	 9�uF����>�)?մB�'��>.�?��?��&?k�Q?\�?��>�� ��A@�N��>\X�>A�W�b����_>u�J?ߞ�>�<Y?ԃ?��=>��5����䩽X�=�>��2?18#?��?״�>�6?�ѩ��$N=��?)ps?�b�?ȁb?i�Ż��?M6�>w�>�����Ƞ>ӄ�>���>�u ?Mf%?�2?%�'?�t＄5����T���#��=��=��=?I�;����1��ڀ=1%�}��<DS�=��{����%��h�iֲ=�B.>��>�?��lf�=#�۾�QվT5l>�7�<��8�)f�gDc�n�>H2�>}�?N��>�Z��bګ>�4?�y�>_��"]??2�/?��>�4�=��v�Ѡ��\0���
?�[T?@N㼒�9�D��������r��*�?� Y?A��O
ܾO�b?��]?@h��=��þz�b����g�O?=�
?3�G���>��~?f�q?U��>�e�+:n�*��Db���j�&Ѷ=\r�>LX�S�d��?�>o�7?�N�>/�b>'%�=iu۾�w��q��h?��?�?���?+*>��n�Z4��������c_?���>�3��Y7!?o�[<�Ծ�=u�u���9��ب�����l��C˟�w��z���3ֽf�=��?�(t?�(n?��c?�L��׵`���[�mɁ���V�k��A���?��';�$RB�(�m�5���� ��S���uU=2>���}D���?��%?�#��H�>��K����@���`>gҾ����|�=(���\�=L��=�?�\��̖��!?��>ۑ�>j[S?
Y��:7�( *�,^>��u��U.r=�@�>8F�>��>�ڎ�)�H��I"��9�����Օ��7v>�xc?j�K?��n?p� +1�����c�!�{�/��c����B>�j>M��>�W�Z��C:&�yY>�R�r�i��w��8�	�t�~=|�2?m(�>*��>�O�?�?�{	�ek���kx�&�1�㓃<,1�>� i?<A�>�>�н"� ����>��l?���>��>ߖ��aZ!���{�ާʽK&�>(�>��>��o>+�,��#\��j��O����9��u�=+�h?���=�`�Y�>�R?]2�:��G<�|�>��v���!������'�&�>X|?ɖ�=d�;>'�ž�$���{��7��V�,?�W?�k���$��˅>~%?���>��>9�?F�>�ƾ	�⻞�?�Z?�F?�
@?���>o�Y=�_w���ǽ�~!��(6=�9�>�J\>_�z=�f�=x����]��f#��Ib=Ш=�\����q>�:MU�>k<k8�<{�5>-ۿܧK���ھN��O���]�
����xæ�+����}�L_���Ι�� y��D���$�k�W�Ea�
щ��m���?�g�?����냾I����~��������>�Jv����6
��H�����ܾT�����#�G�L�`3g�,�c�@�'?�����ǿ���:ܾ.! ?�A ?7�y?��>�"���8�,� >�C�<,����뾯�����ο9�����^?���>��/��u��>ू>�X>�Hq>����螾�0�<��?1�-?��>��r�*�ɿ]����¤<���?,�@�fA?8T(�(��,J=-�>�	?�E>�3�l�rY��F>�>��?B��?J-=aEW�O����#f?<�{<<�D��Wػ�F�=�q�=Y��<��cQE>]ː>�!���D�_b߽�7>�~�>+���E
�I�W��<N_>�qѽY��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=xg ��LĿ0'�\�!�t��M��欽m'��b��A���a���3^m� -���=|��=+�2>g+�>|%d>��G>)7V?Nk`?��>��J>)�����s�r��1{<ߑ�
H>�w�w�w����H:־�iᾛ��u
�3P�W�j3��@4>�6�ǚ��G��G]�'�T���E?��>���eؾ��.=� ���+�������==E==+�o�Ҁ?�J�>�^��;�}��vR3>���Q�`?3�s�!1��=�q�R}"�R~�W-u�;\n=g"�>�O׾k~��≿Ȉ0?=??d���!���*>������=�+?��?�c<K�>R%?�'+������Z>�3>^��>��>C	>������ڽ�?��T?�� �!ʜ���>+��p-{�	.`=�#>о5�����Z\>���<�����T������n�<HHW?�;�>�)�������|u�R@=g�x?�?=��>Y#k?��B?�å<XB��Z�S���
���v=�W?�
i?w�	>���тоsE��y�5?�e?�M>UGh�Cg龅�.�iA��*?ؕn?
?�����8}�-������n6?#�v?�q^�s�������V��;�>HY�>~��>��9��h�>@�>?�
#��G��S���
Z4�Þ?>�@��?�[;<;�'��=�:?�[�>��O��<ƾq��=���mnq=� �>|���*ev�����O,�6�8?���?���>����r���=�O/�E<�?�8�?�iZ�i�=�쾙X���پ�i<�	;G���~Nt=y�Ǿ><"�A���Z�<��=������>dz@�40=���>���;�+ҿ�ֿ�l���	�C���F;?���>�E<��K�/?�Lo_��T�'2_��Ǿ$��>&(>?�X�TZ��ba��#�X�q=@��>u8Q�Vݛ>|�Z�h鿾���K�m=���>�>翟>'N��D��>��?�'�	#ӿ�h�����p�d?���?�G�?+�#?�)�=.͂���1���ݼl�$?��^?�U?y�')w�ɶ`�2�j?�_��]U`�Ǝ4�HHE�SU>�"3?�B�>/�-�ߴ|=�>T��>Zg>�#/�m�Ŀ}ٶ�F���O��?߉�?�o�%��>k��?hs+?ai��7��k[����*�k�+��<A?�2>)���H�!�)0=�bҒ���
?Z~0?,{�Y.���_?ɗa���p�Z�-���ƽ2�>��0��\\��{���d�We�L���#/y��?�X�?^�?���"�Y7%?��>T���NǾ�:�<�{�>78�>��M>�\_�^�u>}���:�Y�	>��?�q�?�h?"��������5>|�}?�$�>��?Io�==b�>�f�=)�z�,��j#>�#�=g�>��?,�M?L�>�V�=
�8�e/�)[F��GR��#�!�C�\�>t�a?݂L?-Mb>����2�f!��uͽic1�RO�XX@���,�ڜ߽(5>��=>�>��D�xӾ��?Sp�-�ؿ�i��ep'�{54?H��>	�?��C�t�w���;_?mz�>�6��+���%��"B�Y��?�G�?'�??�׾�O̼u>.�>WI�>��ԽR���假�.�7>�B?��D��_�o�^�>���?�@�ծ?Ei��?����:��x�~����~7�r1�=�7?3�o�y>��>���=�Rv�\Ǫ�e�s�'�>�C�?�X�?"��>�l?0bo�A�B�5(1=V �>[�k?$�?�̺=��*?A>h�?����󎿲^���e?��
@D@fr^?d���]��v�m��Ѿ|<㾽�='1|=XK>�;�B���#=�w=CH�A�Ѽ�R�=��>�˃>�__>e�h>/M�=s8��Z��d���\���0`�Ė"�H �E�=��h���_ξ�B��Ow���������tH��.�j�;�T�ғ�����=��U?�R?�p?M� ?́x�T�>����M?=�}#��τ=30�>i2?��L?]�*?lؓ=����i�d�`���A��Vȇ�˃�>�qI>�~�>I�>!$�>\}T9�I>�/?>ހ�>>uk'=B���d=y�N>M�>c��>	|�>�$>>a�>�W�������h�"�x���̽�4�?����@K��U���i��h �����=�O,?�J>�Ց�P�Ͽ5i��a�G?*x��L���s&�Z >~�.?׃W?�L>�n���A���>pZ�m�m��>Z��1�m��'+��WD>{7?�M>~|]>�4�As;���Q��s���e>��7?�㼾��E���o�CK�1~��i�9>��>�;9Z�����^���wi�L�d==�=?G�?~ͽ�H����g�ls��2Jn>L��>AT���ݔ=�=g>:Y(�/���IqK���><�{�=r�s>�?)�>.ő=�7�>e牾��$�+,�>m^2>�9>8(E?wJ ?;)I���n�����w7�[�q>���>�Ń>L#!>��K����=�u�>��e>Nx�;�6�����S6���S>��Z��8X��q����1=���3w�=4u=��ҽ"P@�8�=�~?���'䈿��e���lD?T+?Y �==�F<��"�D ���H��F�?r�@m�?��	��V�?�?�@�?��J��=}�>׫>�ξ�L��?��Ž5Ǣ�ɔ	�-)#�iS�?��?��/�Zʋ�<l�6>�^%?��ӾmW�>����Z�������u��#= ��>�8H?~Z��%P�T�=�{t
?�?
T�?�����ȿLsv�-��>d�?z�?��m��?���	@���>��?�hY?@ki>w۾&eZ����>�@?�R?:!�>�1�d�'�%�?)ٶ?���?�I>퍑?՟s?m�>�"x�}Z/��6��Z����i=b�[;;e�>�\>�����fF�ד��g����j�n����a>��$=�>?��2��-;�=[����L���f�G��>�-q>)�I>SY�>g� ?�`�>��>�=�q���ှ񸖾��K?���?-���2n��N�<Z��=)�^��&?�I4? k[�}�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��H��<��K>*4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��WS��GB�>�e!?���>�Ү=ۙ ?��#?��j>�(�>CaE��9��X�E����>٢�>�H?�~?��?�Թ��Z3�����桿��[�u;N>��x?V?sʕ>b���񃝿�kE�:BI�<���^��?�tg?rS�0?<2�?�??`�A?{)f>؇�)ؾo�����>��!?�����A��#&��'���?�B?}��>-1���ֽ_ϼ���iO��}�?�.\?��%?ӏ�N�`��¾�E�<E��ρ<�b
 <��>�^e>#�>R>���=��>}>�=2m���5�k�k<Ѽ=^�>���=� 7��(��=,?a�G��ۃ���=e�r�xD���>_ML>e����^?9j=���{�����x��{
U��?���?k�?���q�h�D$=?��?E	?q!�>�J��q|޾����Sw�}x��w���>���>eol��򏤿����F��q�Žk����>�C�>O�?�*?mZ>|�>`����0$��B���D^��C�818��>/��������e�ռW�¾4Pt�w!�>�y�q�>��	?l�i>v>���>�/��{��>�ZM>[�x>Ui�>b�[>rE.>�r>�;�;�ɽ3:R?������'���辸����*B?�md?	*�>�pi������N�??��?�r�?>v>�h�+��r?C�>r���s
?4�:=�����<i������f����n��>,e׽�:�M�lf�ba
?S/?i܋�hc̾I)׽-�����n=�M�?��(?�)���Q���o�ƸW�S�O���6h�Lj��Q�$� �p��쏿�^��%����(��r*=��*?g�?ǌ��!���&k��?�bdf>e�>e$�>+�>2uI>��	�i�1�[^�M'�H���aR�>{[{?�Z�>�H?�;?��P?�EM?LV�>�e�>A7����>s�=<���>!y�>��8?�-?�l/?��?�*?�2c>*･�����־�?��?S�?t�?�?����Ž�䩼W'O�Xz�kU���i�=�"�<]�ٽT�j��N=T�S>���>xװ��k;��'���1�=1'?�^�>w6�>+Sо5����� >��>j�?��>�R��|��+^ᾍ]�>��t?�N�>�
>�%U>��>E�=o(�?B1>ö��5Q'>�ܞ�����$�K�>��=ܣ8�i�<�>C� >��_=�s�>l�?��>h:�>oA��� �y�����=�Y>)S>X>�Bپ�}���%���g�hy>qw�?�y�?�kf=:+�=	��=�}���S�����9����:�<��?�B#?{TT?���?Q�=?�d#?p�>�'�gK��_�����H�?�)?E�>��뾚;Ͼ����L�_�k��>a"?9.i�Re�ew�o�.���ԾX�>٥T�0�@�B[������,���������<A�?��?׺�=j4#��t��7o��ٔ��v��?"+Y=�nN>��6?�n���)��A���/>���>@eJ?���>���?�0�?�kf?�O�>;7�76ſ*^���a;>�5;>�mF?�f�?�ޒ?��3?4uH?�>@�ʾ��
�vܭ�aą<���D���G[սA�	>|��>0��>��>g9R>���*�����^�ƽY~?>)�>�y>�?4�?E��>.�E?¶�>G��<W�(x��6C��og���v?���?�&?C�>=���YuE���g��>{H�?��?��*?-�b��*>sr������#o��6�>���>ށ�>Q{�=K�<��>�V�>�D�>/u�U���|6�]t0�<
?-D?�J�=:���/��8|��վiݿ��ز������>~#i�@��k� =�J����{q��_��;���c���*�h1����>gS�;�)9=
�m>�`�=#0> �,>J[=,�$��e=WA>P.�=ȴp>�J%>l�}�m��<>�7=Օ9>f�˾u�}?;I?3�+?��C?��y>�<>�3����>�����@?@V>��P�2���a�;�[���Y ����ؾbv׾L�c�"ɟ��I>V\I���>�83>�I�=�L�<*�=�s=�Î=<R�?=n'�=
O�=�e�=���=��>U>�w?�r��<���hTQ����v:?��>y��=g�ƾA�??{q?>I��a������T�~?h��?��?��?�Uk�쉠>B�Bh�����=1ݝ�Cn1>G��='3��ڸ>eK>̲��^���;���J�?�d@�h??�����Ͽ[)/>�
�����ʻd�?k*��:����L�B��/?�&a����l��>�n%>�޾��m��=�Q �,�=�]�PA7�T�=�_���Ϲ=K��=]2�>�6>�A>:D���}7=٘~��f=wn>!�Q=�Ń=.��=$�$=��8=��>�r>*��>�x"?ƨ6?��h?��>��4�vd�O����mR>�(>Z��>��h��Oa>k��>	9?��;?�5[?���>h�>�S�>mx>��M��{J�!��'H���=^�?m�?�Q�> b�ؐ��%���7�ܢ/�H�?�C?��>
�>���)=ܿ�Z'���7�Wm��^/�<]��1�\�_�ۺ����5��c�㽜|�= ��>��>Tz�>�O>C3>�21>'��>�|>��<V��=;�L���;��g����=�w}<Y+�<���;k�ܻ��=�o�*=`ü��;��=_3K=^��=���>�;>6��>��=�����F/>�����L�z�=�K���-B�u0d��E~��/�1V6���B>�/X>�|��n3����?�Y>5g?>��?�Au?��>@)��վ�M���.e�1QS��ɸ=��>��<�[y;��P`�N�M��wҾ6�>�k�>Au�>?>>��(�+�F��m=�E�e:�WE�>�3ƾ������_�7��g���Չl�Jtӽ�!?4���L>�?��%?Y1�?��?`<h�F��RF>�T0�I�>@^�g���0ܽ�{?
?�5	?�㢾A�3��p̾�"��ʶ�>�I�D�O�����Ǽ0��a�\7���O�>e㪾K�о�3�e�������`B�Bq�{��>N�O?h�?��a�H��XO�����ل��8?�{g?��>B1?8\?i��������A�=M�n?���?��?�	>N��>�<j�m��>��?L��?��?]چ?�%s��3�>Ҍ�>�G<O
o��0�>��V=~�F�)5�=�b�>i�?��(?!q�����R�Ⱦy=�v�r�Cw��U�=�YJ>��>>|0�=�n�<�>�b�=[��~�!>��>��>~\�><>Oǭ�M�����%?��}=1�>��.?|M�>?p;��DC=NE>�s����Vo;���=/[��֡>Ar$=XR=��!����>�ƿ�k?���>�/�3�?�Ծ��c<�/�>�=Fd7����>E�>,�%>�u�>�;�>�I=s��>j�N>/�Ӿ��>��h!��tC���R��Ҿ�6{>�5��k�&��+�+����ZI�S��m;��j�c�����<�dݺ<�:�?R����k�*)�y ����?�~�>6?��������'>���>��>�{��������uy���?��?�8c>�>��W?@�?l�1��3��uZ�V�u�'A��e�L�`���������8�
�	��v�_?h�x?9yA?lX�<:z>F��?'�%��ԏ��)�>/��';�OD<=�+�>T(���`�6�Ӿ�þw9��FF>B�o?�$�?aX?�WV���;	�>�3?79?��x?c�;?`=?�<�E)"?J7b>R� ?���>$0?��-?��?el>'��=�;l��={��d?x�����4�ֽ�1���C=��=��A��B��<6<>�<U���4��B�<kid���A<[V$=d�=w�==(�>��W?���>�l>K�:?����'-�c���N.+?_�u=.���c�҆��[�꾲�=T�m?�W�?�_b?2܂>D�:���?�J^>t/>�>��c>�(�>��GL�Xz=|�
>��>r��=7�����'|�������<;>_��>
g|>׀���w'>����z�+�d>�(R��뺾R^S��H�@�1�Mfv��Q�>�K?{�?���=ɜ龁?��PTf�gG)?Xg<?sM?�	�?o��=��۾h:��J���d�>���<��`���	
����:��
�:ct>�����Ծ�
L���:�|w ������R��m��2�>�fU�4�GԾ`�����5齆&�������%�_��:Խ�1FJ?r�t<����T������tV�=��g>���>ҶZ�P=�=�E]������=�)?(Ţ>��=�[5�2�k�u�ؾOX�>��K?�a?&��?��n��Kk�� H����ȧ���<��?���>��?NjW>+�=`]�����-�c��gD���>S��>���D:�8�����W%�0Ճ>u��>³>��?��Y?�D?u%c?/Y5?,C?��s>��ֽr��Pk&?>�?Z��=�ʹ��O�S8�DC�Eo�>�J)?��?�2Z�>h�?O?�(?gzP?��??�>-����<�W��>8�>_�W�c���Ӻb>NN?��>4�Y?g��?��/>]16�"z��)ʝ��J�=(o>�1?i!? ?�ѵ>T��>�Z�� i�>��>�Cx?9	�?
2@?{��ʇ
?��?��r>�gG��y�>:P�>~� ?uT?��u?��A?��,?ᨋ=C\�<��)���:��=�Qp�<��ս���=Ƚb��<�t=��8�EN]=2�a�u�ҽ�;8)��e��g�Ӗ�>w6�>?6˾���=��ƾ��~�LD�>�v��������
 >ز>{I��E�>�6? G��$Ž�٥>!��>�!���;?S:?)��>�ػ=0�^���;Y-���T�>��i?�`�ݩJ�_Y���X�������]?��[?���� �E�b?�]?�g��=���þO�b�ԉ��O? �
?��G���>��~?]�q?p��>E�e�:n����Cb���j�VѶ=�r�>X�	�d�]?�>T�7?uN�>�b>$�=�u۾��w�jq��a?}�?�?���?(**>{�n�@4࿲���^���W?��>$����#?���@�ݾ�)z��u�����2���G��S���(~���M*�f���d����C�=V�?|?,�x?Q�]?����d�#�[��Mz��YT����C��BE�}�H��58�s h���������~��fu$�S낾��<��ڱ?[4$?׉6�a��>�ڛ�y�ľ�:>������T�=Ry~����<�B=�N��F&�Ū�r�?�>���>xkA?l�\�gQ@�?�-�kE3�H���>+U�>r��>J��>�^�<m��0I����S"��Pؽ�^v>q�c?]�K?'�n?D� ��)1�[���ʫ!��0��)��Y�B>P	>b��>�W�����&��N>�/�r����q���	���}=��2?�K�>�Ɯ>M�?��?v	����*x���1�"�<�#�>i?i��>L�>��ν�� ���>��l?���>i�>#w���D!�H�{�Ra˽�%�>��>��>jp>q=,�D\��k���}��T9���=*�h?`v��\I`�]�>qR?){�:D<ER�>&�v�ָ!����?�'���>�c?u��=+�;>��žZ*�C�{��b��Re)?@_
?`�����+�r��>�"?"��>��>ʉ�?�,�>4ľ�<�V?�M]?��E?$R@?���>~
==���x�̽F ���&=�܈>WKV>���=��=}�QT���`s=�
�=.�������d4<���>�<7�<��->�Lۿ�|>��eξCL
��i��C���p��$Õ�sC%�O�"����ߚ�C���o_�哽qB]���%�Ǔ}��qr���?���?D�þ[���O��H���~&����>?~p�s�C���w��+��˓��zҾ�S��JG$�@E>�o[�՞c�f0B?fΓ�l˧��?��Nܾ8?�H?țQ?
d�W'���g��`�=�>&)�hU��'~�۱̿f����k9?xl�>r�6������� >J��>���>�6��n���ݾtK�= /?`�o?J�>�����,Ͽ�n��f؅=�V�?3A@x#K?o�(�jھ]����>b�>=:>�>c�_]����J7>��?��?�Ke�#5f�1��=ݔD?qA>w�Di����V>�=���<�ɿ� G4>��?>�_�������>>��j>�B=�=[=f��L���>(��F�;Մ?�z\�Df�e�/��T���S>=�T?�+�>;�=a�,?8H�E}Ͽ�\��*a?�0�?Ц�?�(?lܿ��ך>��ܾ�M?LD6?N��>�d&�y�t���=rA������㾺&V����=���>�>��,�A��ƆO�>�����=r��弿�m�&����<�0�GS��\���:��`�6唾*d��V�� E=��=��?>��>�Y>��O>U?��b?i�>��=>Y&(��ʕ�K���[=�R���9��*���)��\��I�Ⱦ���d����
�lZ����1܀�T?ԽV~n��o|�6);�'�s�L�g���b?�n1=�<.�B�ľr�*��R�Ϛ2�d0�������\���U �";���?E"�>�\������/��\��U-=��?����	,�n@�@0=�\��P��/���vÛ>���D�L�w��m�+?a�?���H��vN+>ܯ��E=�k#?Er ?� =�֡>�C(?=p+��V��X>�f,>q-�>�c�>�h>���үŽ�u!?�RO?6�Ž�����9�>_x��A^M�d��=�g�=|}A�����)^>�����e�s<�gv��y;<��&?��=�<� �� �Ⱦ�ʲ�j;�=�S?u
�>��=\�s?�Z2?�R{�^TC���3���J�(>�!X?�S?eL.>?� ��mC����]?��?���>(�%�`���/X��l}�>��3?�?���='j�8�������+?v�v?Ls^��r������V��<�>�Z�>U��>��9�n�>=�>?i #�F��x����Y4�5Þ?f�@ҍ�?�w<<[-����=�:?�[�>7�O�l?ƾ����ف����q=#�>&����cv�����E,���8?��?���>����v���_)>H����?�af? �w�)�z=��jx��u���P=G��<C&�<�g�=A�ȾPK�vTѾ��i֑�� ��8�>>h@�t�=̦?���տ�_˿�z��;��!�����?(��>H�<��h*�E2�wtk�f=F�s�Y�ԥ�Y�n>��=��
��G��ʄ���L�HNؼ�W�>@�#=�>Ͽ���n��������=^�m>�Io>)�>��ʼi����F�?r���+v˿������m`?x6�?��r?,
?. �9n;�/;^�[e<DEK?��k?�1?����?(�j�!��k?}���rx\��
7�?K?�yTZ>Je/?�c�>Ҁ,�v��=�P>�V�>�� >]�/��~ÿ�ٱ�����?��?��?n�羂?��?��*?�o�q���s���w(��7;�;?�E%>�?��v��N�5��i���V?,[/?���ś�c�_?�a�<�p���-��ƽdۡ>)�0�de\��L�����Xe���4Ay����?C^�?e�?���#�@6%?�>n����8Ǿ$�<���>�(�>a*N>XI_�J�u>����:�
i	>���?�~�?Zj?��������7V>��}? �>�˄?���=��>�n�=(v���2��>��=N8��2?��M?H��>5��=�>6�r�.�?�E��P���&C�_�>m�b?��K?��d>�hý{6@��� ���½��+�j��<�A��J$���ܽ�e/>E�;>�n>D{B���Ծ��$?�#�kdҿo1��l ��D4?xt�>��>c�	��7Y�G��(,b?���>.������n��| 1�؞�?5��?�?�I��,�B>�Ծ>h>����Ž>���2W>n8D?�������j��Շ>���?$&@7�?��N�b�?�M�Bm���J~�m���7���=�8?>���:y>C�>Ez�=Ljv�ᪿ�s�끶>�%�?G[�?%��>��l?��o���B�Q�3=�>��k?��?F�D�R��ׁB>��?(v��.��$5�իe?��
@�e@�*^?����0 Ŀ�+��B����_��q=>��=e3(>z����b>AS_<�ٷ�`x��� x<mG�>z{>A��>�>0>��=��=����#�����͕��,y���/��<�z/��Ѿ����=d�el��a���y��۫��b�e���!�K��E�=�X?\XT?h�s?R�?\����>�_��z�<ځ�K��=��>n�3?��L?�9.?��=e����^a��J��`��Y����>�-?>x��>W��>~3�>�3A;2�9>sQ>(~>m��=�a)=����<�7>���>���>��>��l>�#>�����z��<�i��z�� y��|�?I���H�@��x���S�A��+�>>^�
?��>�����3޿�T��&e@?~ ������R���=�6-?Lt?!�&>6狾�W�=$��L#/�󷧽��=Y3>y��fL3�3R>�)?�Q>�+�<F�?� B�5Xk��_��z>H>Wl?bw�5���ݒt�S'b���Yȃ=f�>e�D>pH��樿�)������>�-?Y/�>o���z[P���%�rp����D>? >�.
>'�r>�	�>h~�d�꽯ΐ��\>�Ŕ>"��>�J�>�D8>�+~=�]f>Le�f-8�7��>�̳=k�7>��D?t�?otv={��������J���V>��>6c�>TF>�RR���>?�?��Q>pf<E�Ƚ��7��*C�x��>z����n����Ҧ=�*���[<���<-��7�*� �K��~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�-)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ#�>e�����H/���u��)=���>8�G?ɏ��N�o)@��K
?�?���Ξ��/�ȿ��v���>2��?��?�Vn�M���@�w�>Q`�?�JX?Ɩf>#ܾ�SX�K��>C�A?�iQ?nҵ>�o��Z&�n�?g��?R�?M}^>�6�?c�u?���>�B	���&�§��%Ŏ���=h��;�ڊ> $+>:��_�4�&X��}S���g��u�M[D>�;9=dO�>����"I��� �=:�������2��X'�>V(H>U�w>	�>v?_��>.I�>Nc=r �1���
����K?���?����2n��I�<]��=ѱ^��&?OI4?�i[��Ͼgը>��\?X?�[?2d�>���X>��)迿�}��t��<��K>�3�>PH�>:$���FK>�ԾF5D�\p�>�ϗ>�����>ھR-��]W���A�>�e!?ϓ�>�Ӯ=�� ?��#?5�j>2�>T\E�V9��]�E����>��>�H?��~?
�?�Ϲ��R3�����塿��[�FN>r�x?mV?�ĕ>i���r�����E���H�3�h��?vug?���8?D/�?��??��A?\"f>-���ؾ=���3�>8�?���p@�B��)����>2�?�M�>(ڿ��)��!׻������j	?/�i?�=?��sU^�����t =]�=���<\�~�ֈ����>k,>p�ٽ$��=��R>�9�<�k� 5��ۼ���=Cϒ>�(�=.�7��a��:,?��G��܃�ژ=��r��xD���>�DL>�����^?�i=�d�{�����w���U����?���?�j�?��ٝh��#=?��?!?|'�>H��B�޾���;Bw� sx��y�*�>��>˦l�徽���|����D����Žq='�{c�>���>�^?��>`7?>���>�H��.� �6,�2�u�Y���e�5��,���������0��x�cq��?s�S�>�q���7�>V?
?f�\>��|>�o�>;�B��σ>��9>�A><��>/�>>1�1>6 >Gd��RmɽmdP??��e�'� 2�����jA?�Gc?9��>��x�O���O�W� ?(�?��?S>|>b�i�u�+���?���>� }��3?��[=���y�}<%���v���y������>[�ؽ/v8�lPM�Ğj���
?��?����%w;�7ܽ������n=�J�?��(?��)��Q���o���W��S����)h��k����$�ߚp�(쏿�\��a"���(��1*=��*?��?Z�����"��n$k�;?��Vf>��>` �>W�>\{I>��	�ؼ1���]��M'������V�>-[{?!��>��K?��R?��h?�:R?r~�>5��>�TȾ ��>P5<>>�W>�T�>&�5?�%?!�?��>��,?eܒ>���<�5��������>!�?�.?�P!?�?��J�B@�<A��<\�������x���7
>�t����=��$p�`N>��R>x?����Up,�
�J�s>	�1?�9�>7�/>�W��AJǽ�<>Y�.?[��>�O�>����n_��꾩�>��t?d���{>"M>˅>��Y�m��<�JH;����oڴ=6�ͼRy=/g >!P)>Ud��:�>|d<R�6��
�3 =*t�>�?���>D�>�@��o� �:��ee�=VY>�S>�>�Eپ�}��b$��G�g��[y>�w�?�z�?O�f=e�=}��=<}���T���������:��<�?AJ#?�WT?��?V�=?j#?$�>�*�{M��o^��V����?��,?~j�>�l�w�ʾ���*i3��|?��?�7`�H��e+��ľex׽��>J�,��G|��7���%E�������+���[��?{G�?�99�3�4���������­���B?�f�>��>��>YY*�W�h����5=>���>��Q?��>2��?5I�?Ax?�m�>��%�Z˨��럿́�*">�?8?�u�?b�?Ň~?K�#?V��>8Ӿ������q���i�۽��ӽv��>$x>�@L=�7�>s_�>���=���=??����}�������=�� ?�c�>�c�>��s>~��=��G?2��>�Z��Q���⤾����6�<�(�u?ϖ�?�+?N�=�x�B�E�9G��#<�>�n�?u��?u4*?�S�״�=	9ּ�۶���q��*�>�׹>�(�>���=N�F=�f>��>��>n��V�}p8��fM�j�?�F?A��=�����P����޻�2�ؽ���z��%������E�n�9��D��5��ZQ����Ҿ8uD��H��X�}�� �>��=}�T>9�>��
����[>�8H<[�=�R<��y�y	d=�޷���>�৽��+>�u�=��=��ɾV�}?�:I? �*??�C?�|>a>::�u�>P�u�%�?�R>�#G�����r:�h�������־8Iվ��c�a࠾e~	>-�D�S>��.>���=��A<~��=�l}=ϕ�=�xY8�=�3�=&�=B��=z��=>}>�6w?W�������4Q��Z罤�:?�8�>j{�=��ƾp@?|�>>�2������xb��-?���?�T�?<�?Bti��d�>M���㎽�q�=M����=2>y��=t�2�S��>��J>���K��C����4�?��@��??�ዿТϿ5a/>��ռ J�na�f3�`�ӾH���$?���0? D=���"��>��̺���/�����^��6V>=�=o�k��j�a�z��@>b>���'�>$�>�"�<W�þi�M>�	->�?>"��>O�=5{��I��M=}�>�b�>��>F�>"�<? <J?��v?0O�>�Ϟ�5���ͧ��-#q>��S>b@�>
0=�Kw>�h�>�-?#i?*�J?���>U�9>[�>@��>��!�TV@�4���V�����p�?%��?���=�N���8=�@�)�s���(��U�>ݷ?N�>�ה>�U�����X&�M�.������T4���*=�mr�UU�I���6k�ͮ�
�=�l�>���>��>�Sy>2�9>��N>�>��>3g�<=��=���Q��<�ڔ����=g���$�<;iżh�$�&�E�+������x�;Ey�;��]<J��;I*�=��>��>PK�>D�=�{���,>�����L�d߽=2���eA���c�	�}�&�.��'5�D*C>ܐX>�K��<��J�?
f]>�'=>�}�?�?u?��>]N�?�Ӿ􆝿C�h�X�S��;�=Y1>�b?�%�:�ë_��QM�t?о&��>���>0��>b3h>0+���=�~
s=]m㾒V4�m��>�>��a������p�L��ֆ���\h��7r9�^D?�Ӈ����=X�~?�I?�w�?D(�>����уؾ?�->�j��\=�
�d�s�����V?9�%?p��>̜쾾�E�P�����Z�>ޞ;���R�>�����/����u̝���>%8���t����3��{����\�:�K���Uɷ>C>?zP�?��l�XTv�=f"�x�"��� ���?CG^?K��> S�>L?$�:��𾡕��~�=]�9?C�?F6�?j�%>���>`���'-?��:?HO�?W�?��z?H熾��9?=��>+⟼�䳾��k>~Y>&��=��f���?K.?��?2~Ͻ�5循X�����d�V�(=�4=d�-=�S#>m�>1�����=�O>ا��W��>�?�>��>�;>��>뮥�����$?4�=�>E,?`|>qd.=�C��A��<kT;�d8�d�'�����&A��o<���<v�{=�K�����>��ſ�{�?��w>�)�5E?��辛�5�~:f>tGM>���$��>{8>H�>k��>yғ> >�f�>�+>̾�!>�*��"��rC���O���Ǿi�}>�G���_(���
�)��w�B�Q��K���Pf����r�<�Jg\<��?��!�g�'U-���ԽK�?���> �,?Gߎ���o�"�>�T�>1ؒ>����V떿D*����ܾ���?�?�?�c>P�>��W?��?e1�U*3��qZ��u��A���d���`��ݍ�����V�
������_? �x?�vA?莒<�Az>��?#�%�gӏ���>D/��#;���<=�-�>;���`�|�Ӿ��þ5$�\F>��o?M �?hI?�cV�yf�<��j>b�??ł1?�Tx?��C?&�;?<���5'?��t>��>=�>d2?A�?O��>
��=��<>P�N=���=�C����1,ѽס�ွV��<�=l�۽���<��>-'�<��<�� a�� ��������=�=,W�=��=�ݒ>o[?X��>�8v>CJ5?C8�"20����,3?�!�=4����k|�e���'��z�=LLY?��?}Y?<�i>4~C��E>�@oQ>�.�>��9>W2W>恛>Խʠ��G=��=�ȯ=^(�=8F��ծ���h�:����zۺƌ>A^�>��}>� ���z%>ջ��)�{�j�g>�KQ�jɹ��Q�~�G�e�0�؉w�+G�>�L?�1?�@�=� �し�d�e�9q(?��<?�L?1�?eX�=�Fܾ�>:�ZfI�J��1s�>��<���G]��BN���:�~��;�w>����*n����z<�����J����-�j���!�>~�I���i��A.��3�ɩ�A�C�J�'>ʼ����(����0���??'�8=Eu5��q��h�۾x�v=�:�=�>�F��F)="U5�©���:�=�:-?X�>��<� (���f�)�6'�>�"W?U�l?��{?��D�Mlo��@�����Iľ�<9X?��>�{?���> �=H����h!��L\��;�l>�>��?�~���Z� ����c��bV�>fa�>1��=l�?!�U?�q?�j?{� ?�r�>bm�>ad�������$?}ւ?��=L�	���N�.7���D�z�>��,?0�.���>��?a�?J$"?O?"�?pZ>ez���F;���> �>��U�IL��G]>7�G?��>�&V?0��?�2E>�!/�<����]�����=�>��1?�`$?B�?mȫ>S��>����R>\+?�J|?Wښ?��?�8y?�6�>�`�>n
��X7>�H�>.;&?9�I?3Fn?�E?$k�>�!��vӽ�ὼjԽ��P�)����V��y=6h�=�ν��S�1A<��=���/J=Q��Z�9��y�=��g��L�>��d>w��m��<:þ�
��=B>n��e=�h��걇�p�?e��> ��>���>�2��A�<��>i?�@�w�)?�9,?��e���=��T����-�~��?%|]?�^ɽ,�.��.[��r�J��:ֲP?�,Q?����c�M�b?��]?;h��=��þ|�b����b�O?>�
?&�G���>��~?f�q?Q��>��e�&:n�(�� Db���j�*Ѷ=^r�>LX�T�d��?�>k�7?�N�>(�b>,%�=]u۾�w��q��a?��?�?���?+*>}�n�W4�p~���E���^?�x�>�E���"?�]�O�Ͼ?���$����������7���m���$�l˃�		׽ ��=��?ws?VLq?��_?޼ �� d�D)^����dV�x+���w�E��E���C��n�ef�����
���G=Uil��U1�m{�?k-?�#���?b]e����e��)y�>")m��`=mO'�\�/>�>%������X��"?��>�U�>�P?��k��KI��D�}E$��x�1Ҍ����>���>R��>:~�Lo��!�$ס�EC`���y��7v>�xc?\�K?��n?�o�+1�����T�!�r�/�sc����B>�j>O��>ǯW����Z:&�dY>�1�r�S��w��K�	��~=��2?�(�>c��>�O�?�?�{	�Wk��lx�4�1�g��<21�>� i?-A�>��>.н$� �n��>��l?���>��>i����Z!���{���ʽQ&�>�߭>B��>��o>C�,�a#\��j��_���j9�v�=��h?}���1�`���>�R?��:�G<�|�>Ӧv��!������'�b�>V|?���=ȝ;>��ž�$�1�{�c7��ڻ)?�?���nW+����>�?"?��>8�>Р�?+P�>sK��7;�W?��]?^UI?�NB?�W�>~iL=r���;ͽ,�'��g.=A[�>w-\>�qt=�=����g[���`�"=�ذ=�ո�}%���M2<�]��#֡<�=��3>Ѣ��P�x�Wsܾ�r�H���_���f�F����=���C���_����о�W����¾��m���ڽ���W�?��?��� s�,���?���(��_�?fW����I�����G5.>�?����C"���I�XlT�`&x�U�W�Q�'?�����ǿ񰡿�:ܾ/! ?�A ?3�y?��/�"���8�$� >�C�<-����뾪����οA�����^?���>���/��d��>㥂>�X>�Hq>����螾�1�<��?7�-?��>Îr�.�ɿ]����¤<���?-�@��A?�'�U�쾞�@=��>��?�>>��2������"��>w�?@c�?²M=S�V�u�wce?�z<��D� ۻ�b�=�q�=��=ۡ	�F�O>hA�>�T!�$D�d�ܽ�*1>XM�>A�#��q���[���<Ģa>gH���ʍ�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=u6�剤�{���&V�}��=[��>c�>,������O��I��U��=ڹ�ѿ$�����8*f=z�S<���S������_#�����9_����D�Z��=�V6>tQ�>��>�ì>�hy>�`J?�_k?�6�>+l#>N�B������8;같<����]�����Nf콨���aL	��� ��<!��� �# �1lҾ0�R�{	�f}Y�|����?�O�m��L��[]?`�&>~B����.? �D�۾��A�ƫ;V˩=���n���{�-��?���>�ǖ�$<&�r>���+>�9��a|?����ǹ?�w��=����w�򒮾�k�>�9=����c!���k;?�
?ӧ���U���f�=�:��7(=�6?@��>ST���ۅ>a'?���h9��s�<�(�>�a�>kЙ>�U=�g������L�(?*(M?S@�����A��>	�����7O5>==:�ؽ�9��o��>�R=B��7�r�7�z�==Y<?j>7�)��?�۾;�ƽi-�<J�W?eg�>�$>�M�?��3?�� ;�ņ�q���&P�7�
>"�J?�T?J7:>�	h��X��.��#1?77�?7�>
� ��(���,��}����?d�M?�?�R> g�?꛿�{Ծ��=?uw?�{]��,��y����S���>�K�>��>739�`E�>��>?ސ �����j$����3���?xv@~��?4�j<W$�h�=��?-�>�.M�u�ľ���Z���$m=Y��>.ѩ��uv�;��1�*�A8?L��?�� ?�~�
���">�!���?p̎?�8�!{<���	�y�vs��$�=�r�=E��=9�;����A�lخ��%��I��P��o�>ۚ@���=��>}�G��޿�ǿ𨀿�"��Ї���J?g?�%�=$ĥ�ɉP��Gm��'K��X�����E�>^O>�\��CԐ�F|�y0<�.�ϼ�j�>��߼j��>��G�����A����4<O��>��>���>Lͫ�������?^����Ϳj����W?�?�ф?� ?/�;��i�I=v�PT���E?�p?�T?&�(���U��>��j?m_��aU`���4�cHE��U>�"3?�B�>�-�`�|=�>@��>�g>a#/�3�ĿOٶ�����0��?ʉ�?�o�5��>y��?�r+?mi�8���[����*� i*��<A?�2>+����!�n0=�DҒ���
?j~0?v{�?.�]�_?+�a�M�p���-���ƽ�ۡ> �0� f\�N�����Xe����@y����?N^�?i�?ֵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>cH_���u>����:�
i	>���?�~�?Qj?���� ����U>
�}?oֵ>f{�?���=X��>�=�P��ܬ(��� >�;�=��G�2�?��N?:��>J��=rV6��.�4 E�;�P�_b��C�@��>��b?ǱI?�e>����H
8�PQ!�½~l*�.k��?��])�~e��7>4�>>��>�D��Ҿ�?HZ�ňؿ�k��I:'�b%4?v��>V�?ÿ�Vt����)A_?y|�>[1�����������?�:�?��?�׾��ϼG�>��>%v�>�Nս~���k�����7>�B?�%��>��}�o�r��>2��?-�@��?"�h���	?�L�����~�ǔ��=6����=x�6?����>ڳ�>�}�=�Ku�I��;#s��{�>8��?p@�?j �>��k?W�n��@C�R*=[��>��k?"V
?@���$����A>'�?W���������zKe?	�
@T\@e�`?G��xhֿ����^N��a���v��=��=��2>&�ٽk_�=��7=��8�>��|��=x�>�d>q>U(O>`a;>�)>���D�!�r��A���l�C�������Z�3��/Xv�5z��3������v?��%4ýAy��BQ��1&��>`�?�=9�U?LR?�p?Q� ?�:w���>���|�=�6#�u�=�+�>�d2?��L?F�*?:!�=����>�d�L��KJ��tƇ��f�>8hI>��>�R�>�"�>hс9��I>��>>�l�>�� >7I'=+��&=�O>*[�>G��>���>$�6>�s>h������`6j���y�Yp�����?SO��D3M�����������>^]=�+?�2 >;Ő�'�п+���ӻE?�T��v����'��r>��,?��R?�n>�����+��>@�ܘc��#>�V���j��^)�:�D>f�?��=誥=��B�u�U�ZtB�h�����x�PO?�	;�{�/�"�W-���ھE_�=q>�)3=� 	��U����~�0���1@>�M`?y��>���=O~b���KR��J�>~�>�_�����>o�
>+�:=%�#��_=mM>گ?O�?�%>�\p=թ�>���b^���>5;>�b7>R�7?4u?%t,����V�����G�D�>�.�>��h>3�>��l�:z�=�?�Pd>0;�m�������z�.W>4%�;Xhz��S��1�=�<����>�{=�νѲ>���=�~?���(䈿��e���lD?S+?] �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��L��=}�>׫>�ξ�L��?��Ž5Ǣ�Ȕ	�1)#�jS�?��?��/�Zʋ�<l��6>�^%?��Ӿc]�>,^�$J�����u�;�=j�>�H?�����O���<�Yn
?��?F򾆌��Q�ȿpv�}��>���?0�?{�m�C����?��M�>ד�?�SY?2ai>��۾�}Z��>$�@?"�Q?/�>���E(�K�?ض??�]I>���?��s? m�>�Su��\/�%�������z=�$z;���>>}>,%����E�.���HY��x�j������a>�/%=�>U��㼾�i�=51��Y6����d��v�>T~p>��I>�>�� ?���>���>�$=-������H2����K?A��?d��b3n�)P�<9��= �^�	&?�I4?�[���Ͼ(֨>��\?���?X[?�c�>���=��?翿|��Ҵ�<��K>�1�>H�>�%���BK>��Ծ�4D�`q�>?ԗ>uࣼ�Aھ%-��pף��A�>�e!?Ɣ�>}ή=x;"?C<"?1i>ן>o�@��t��iRB���>��>2U?�:|?��?�@��-0��ӎ����>Y�_�=>
�v?w?�d�>)����Ǜ��|	�?�N�(��4�?5'a?1���4?�E�?k�3?�];?ٷK>^���;Y,n��u>�\!?�)��'B�L%����?&A?�J�>����/ݽ7��4R�+����s?�\?O%?X��rQa���þZ�<��&��L�>��;�N$���>��>.%��m�= >ɨ�=awj�^65���r<d��=�C�>�:�=U�5�z牽��/?�����o���=UCo��H���>�L>�Ӹ�Eq\?ET��cs��N��^���s�Eҋ?�H�?]H�?�_��	�p�(�=?D9�?z�?�9�>�ಾb�ƾ�� ��j���)�s
��>���>=!E<��þ�O��u?����~���u���)-�>h��>��?�9?��Z>��>����,"�|�پ�H���b����1�D�1����vی�N3�����ʾ!儾b��>������>(�?yl>lj>n��>���;���>��0>�Ss>+k�>Ěd>Qj4>���=�ձ<����v�L?����*�3Ҿ*���4AD?8\b?�(�>�m�����x��O� ?��?�I�?Y�>�Bg�y�/� �?w�?텾�$?�bX=�{E��=�<�۲�s�!��b���� �䅖>Մ��0�ŪG���r��3?�}??�i<IȾ�ٽj}��Go=�J�?��(?5�)���Q���o�ײW�"S����/h�)`����$�I�p��揿�Z���"��N�(���*=�*?��?̕���#���&k�g?�mhf>���>�+�>���>֏I>r�	�Y�1�^��I'�|����Q�>�P{?�ڹ>�Bo?_�R?��H?�s~?�9�>�R�>�<����>�,>�]�<�?L
t?��A?/�?���>?���>4.>i	�X��%ɹ>/�?S�9?�!?"�2?Ի���=��g>;H*���پ/�b�s<���=]�E�W��=�U>��?���OK�����n��;�-<??<��>=���!����>ʢ??��>G��>E�i�Zu�EQ�Ԧ�>�߅?��i�=U9">�M���A�=�d�=e�>kcy�Z�=�a�.�I���<��?>�K>H����>�A �4,=�)>���>��?K�>���>񉆾�� ����v��=<�Y>�1R>�U>�Mپ���<����g�4sy>fw�?B�?8vc=��=���=蒠��_�����-˽�@��<��?j�"?;�S?.l�?��=?=�"?�:>�RD���.��n:��yu?b"-?�h�>���ZȾ@���q4�.�?%?� _�^�	��)��_���1���j	>^�0�q�y��G���;E�����%����?$��?$�C���6�3��r����drF?��>�H�>���>�	&�b�o����=>1��>f�R?&`�>I)�?H/�?F�7?*��>��2���1c��)(l��4�=��1?�a�?E#�?J�?&G�>_.�=��r�3[��qg���h�U�"�.�Ҿd�=`B>Ȋ�>G�> ��>�Y>tTE�1�]���&��=�=�>�p�>��z>�r?5��>��>�EO?q��>Y���v9�<����/���]bD?�\�?I7?s�>����0�Z��k=��"̠?��?��?�og���>���(���<Ǜ�>C��>å�>��>���T���C��>�Jy>��� �r��d��=��?�rK?^ ��}�ÿ�eY�7��1$��12�Hc�4���R6������=�����!�ͧ���7��.��4��/��wh��a�-�F�
?5��=��=�e>�"��(I�xc����=��>�l�=t��;ry7=�����8����-���=��{=ᆸ=P����˾Ї}?�2I?Æ+?�C?��y>1$>��3�˙�>(}���;?a�U>��P��{���a;��������ؾ�i׾��c����QO>>�H���>!�2>S�=ݧ�<��=!s=}�=jO��=�F�=�s�=>Z�=89�=�>z>�6w?T�������4Q��Z罖�:?�8�>�{�=��ƾc@?x�>>�2�������b��-?���?�T�?-�?ati��d�>D��.㎽�q�=h����=2>���=��2�9��>��J>����J��W����4�?��@��??�ዿ̢ϿVa/>�+>�	�&�l���7i����|����d?�`v�+�����>�W@���3��ܵq<Gu:>�+�@,�������V	<�@=M\�1�>�=H�?>P8��3��=��'>�J�=Uw�>�X=�=*���i�d<��)>�>0W�>a'�>�?��#?���>r��>�ꋾ�ᾌȾ2��>�mi>��>���=Y��>�\�>��'?�@=?�3?�.c>��=.�>wX�>O*��_�J����2Ǿw
��U�?�n?���>�|M>`z����P�%�� ��� �>�� ?��>��=8H�9}�F&���.��Ǚ��Ն�$�)= �r���T�Nv��E��V��-�=�n�>��>�ş>�0y>0�9>��N>e �>˴>{U�<���=DO���Ү<ɰ����=���o�<s����B\���;��R*�_ܣ���;Tϟ;#Oe<��;�=!��>��>���>�,�=�B��S^�>�䴾�7� �l>�ξ9�A��	5�� b���:��L��o7�>�#�=`�������_7�>Ȏ�>
�G>ql�?|u�?~Ç>�p��bľC����=5��7ʾ@��>3�G>xOi�{%��ZI�f+�u砾0�>2ގ>a��>�s>W�+�T�C�CӦ=9�ܾ)b.���>4ȗ�����<�l��G��7z���	W��<���<?	Y����>*��?�HM?�E�?@��>��K�#��&3>;$H��<���A��O&Q�q�?ך?��>�U��8�*�ʾ9׼��<�>^�L���O�/��� �/�ͧ�����	c�>�餾�w;u�1�!�������@�d)j��`�>��M?V��?�e�l����J�E���Dz��H?�lf?��>��?��?�镽Hc쾂��
ƫ=�j?Q��?���?U6>��Q>�E�=�5?SW3?F�?P��?-��?� Ǿ� ?S,	?������¾�40>"̬>_�>�
�`�>��>}�?3�#�b<�i������i�U�7�*>ͳe��o�>��>��]=�p3=�湽�����>6E�>Z̓>�ok=j0>��=�&���8�_�?��=c�x>��#?��u>a�=Knv���<v�%�'H�3�4����������;+=�<�Ȁ=FS�߉�>�[Ŀ�֊?Sŏ>�J�`�?a��B 2@>��!>/���H��>o�G>�>έ�>Բ�>�>�O�>�K>��Ѿ�=>o3�
y�TOD���S���Ѿ�Lw>����q(���Č��K��񱾕����i�Y>��P;�}��<�^�?����1l��S#�<�S!?�P�>�]5?�����g��%>q&�>��>I�������z���߾���?���?{,c>�:�>�W?cU?��1�r03�~�Z���u�	�@���d�!�`��܍����ߏ
�ف��Y�_?u�x?�YA?#N�<f�z>ፀ?��%�ی���׊>�/��=;�V�>=��>�:���`�<Ծj�þe��lE>ψo?��?�P?��V�,�C���,>C�;?�F4?�Cx?s�6?�=?"��=#?s�>>� ?��	?��6?ae/??8?��8>���=�];:�[=�%��$���̽%���'�����4=~�=�+=��X<%=��<[�Y��R��wD���=�#K=뺬=z��=&q�>� T?#��>�T.>�7?(Z��k�9�89Ⱦ�,?k�=�����}�I����後g�=�tu?X��?�7j?�_�>��g�j\b���I>U�>�>��(>$ʕ>1���ɐ=f��=��">�#>��u��}m�R��m�����%>Q4�>�`�>�X����T>S���M�����>P�d��˪�����N���$��������>/�6?~X?��:>f�ڶ�� |���(?��P?��N? �?��=\��i�H��x?��Մ���>��5�嗾?���64���B.�I h=Z�p>���S�k�a>���3/��s��
=�g�龈0d=cN
���<^��~���n���xu=�P>ЅҾM���+��A���2�I?�"Z=�:���g�._��� >5N�>0�>��`�i��G���MR=X�>��9>�ټ3�ھGJ��L�l}�>37E?��_?��?)$��U�q��B�#c���]��o���M>?�n�>`?3 A>铮=������[?e�B�F�=�>��>�]��DG��0���_���$��;�>%�?�a>X�?��Q?�i
?O�`?i�)?ֱ?'ѐ>L
��8���:�%?ŉ�?;;�=�>ٽQ�V�C�9��FF�Z��>K�*?H�@����> 2?�P?,�$?�<Q?I?�>� ��v@��n�>��>nJX�(����Y>��I?�>@SY?h&�?6=>i�3�놡��ʤ����=��>��3?&�!?�C?�{�>�[ ?8)�����<D�>��s?���?	�p?p?��
?��>��>������>�/?��>Y'8?�0�?��|?"�)?�a8�	ý�E0�5}?��>��,=�^��؃��W(>�~b����;�L�=rD����e��|�29�=��>��=1����f�>ѹ�>��[�)�>Ѩ��������X>�'������"���|�J�&>�z1>Z�?�U�>쀾��=�k�>|7�>���O?cs?@��>�t����_�z�1Fž��?5�b?�>4He�-���)4����>�<]?)sX?���; 3�F�b?��]?@h��=��þr�b����g�O?&�
?b�G���>��~?^�q?`��>��e�&:n�'���Cb���j�Ѷ=Sr�>AX�G�d��?�>k�7?�N�>�b>$%�=Yu۾�w��q��d?}�?�?���?�**>q�n�I4��W��D��"R^?�G�>�/����$?5z��Ӿ%Ȇ�������s���s���'��Ҽ�� %#�/Ђ���ܽ�Բ=ĸ?rr?Q�p?�}a?۳��d��8\�# �V�G�����C�Y�D��jC�L�m�������L!����.=.�c�JWF�k��?F�E?��&���? M�T�:;�k�]>��ʾ؋���t9=~�ʊ<H)d=x�6�m�o�6gž�D?���>s�>Vk?6Qe��f?�B���/,�%��ͭ�<��>�3�>� �>>}������,�ɾ�M�1Se��w>�b?Y�L?�+p?���m�.�7��ak!�V>+�Gݢ�~�>>$�>�h�>�=X�;����%���>��
t�o�G����
�'�f=��2?�X�>(\�>>�? �?TD��g����x�3�2�^�z<"�>(h?��>��>]۽�� ����>k?�7?��>�!!�����8\���ս��>�~�>7u�>J[>78˽zX�؉�Cƅ�:�4��T�=
Ne?Ny�<�����>4oU??�0=@3�=�"�>�ѽ����̾&�9���=�\?�c>q>��3:&�$�����)?��?_ߎ�,(��S�>9�&?\�>�x�>�ۂ?6џ>�nоə��>T?��[?U�B?C�9?0r�>ϡ=-*����ֽX�)��P7==�j>JW>f!=f}�='$���a�tq�5�V=vk�=�#��Hק����9����}��<0Ѿ<=�7>��Ό�R��=��O{��`�7���}���E�Y!�Q��������о��p��� ��C��=����N��*!���6�?�?��f�Q�$֙�0	t������>?�q��-��l�N�������l�������
���F���P���p�ʍ'?8���#�ǿO����Jܾ< ?�G ?r�y?&�{�"��R8�� >���<s����L뾪�����ο(�����^?���>� �p����>ʳ�><QX>��q><ȇ��鞾�p�<N�?*�-?���>��q�L�ɿVz�����<��?~�@Z=?l�%����p�c=,N�>��>,y>7��z ������m�>�?t�?޻�=�^��!_���^?%-<pZH��!��)W�=���=���;c|ེ�t>H�>}�:�n���u���>o>�1��4 �4��Co<!�*>ys��/+�0Մ?�z\�<f�R�/��T��GT>��T?�*�>�;�=ݲ,?�7H�V}Ͽ.�\��*a?�0�?צ�?�(?�ۿ��ؚ>��ܾw�M?�D6?���>ad&���t�_��=�BἼ���I��	'V����=���>Q�>��,������O�)J��F��=9p���ڿ���U4���'=n�u���?7��3g��ɕ�������\���5�B�»k��	�����>�l�>���>��Q?F�w?��>TU>�v���"B�Â�Xq������ڽ� ������#ɾ ��6�򾅢��9���"����<G��)=�l?�� ���nB���a�v)X��i.?��=f�����n󚼎W�~���	�<�OR�������聿E��?�_-?����CD����!���!=4�֒n?{Ӿ���g���GW>c�>���wi�>�ҝ:�ۿ�j�R�<���/?�!?����T�o������'M�s�>=8�?���>C���V�>!?��q��?O.>��\>��y>�Z>sK�=�y�Z8콾'?�NJ?eAv�$����֦>�ʾ]\�6�>خ�=��F����Б>�@�P�;l�s=�鼑��=0T?7S�>p�*��Q��-��Ϯ��`t=��v?�J�>�b�>��p?ʹB?K|�;�u�f�I��]���3=�'P?x�c?d	>���/uϾ ���]�4?�S^?�-`>s�J�'����2�� ��k?��n?Z ?����^x��㒿h��W;?��v?s^�ws�����F�V�h=�>�[�>���>��9��k�>�>?�#��G������zY4�%Þ?��@���?��;<  �S��=�;?j\�>��O��>ƾ�z������?�q=�"�>���}ev����R,�d�8?ܠ�?���>�������p>2�N��#�?C�?�T��j� =�  ��#��\ξ�Tl=7_:�g�=Ao�<�H߾��;��L���������\Xg�8�>�"@+��=Ӓ�>A���N���rҿ��e���
������4?`��>0"�=�䩾�YI��bO�Mn9��E���aq�>x�>�4�������z��;�
�ؼrd�>���hۇ>�O��c���ۜ�
�-<�p�>��>ȁ�>M���˾��r�?�B��xN̿]������Y?;��?#ʃ?G�?���<l�s���|��@G��C?& u?�X?�dE�k�X���"���j?|B���L`��4�%DE���T>'3?�C�><�-���{=>���>w_></�ǇĿ	ն�������?���?Pr���>��?p+?-c��9��/s����*���=DA?�2>]�����!��,=�ؒ�ޭ
?^�0?���(�T�_?
�a�-�p�u�-�M�ƽ|ۡ>��0�&f\�$M������Xe����@y����?A^�?[�?��� #�X6%?��>8����8Ǿ��<��>�(�>*N>J_���u>����:��h	>���?�~�?Dj?땏������U>�}?C�>���?'��=pT�>m��=�0������!'>d��=��`�Q�?�NN?8�>���=��3�]�-���E��R�]��C�$(�>��b?��K?v`>uHŽ1x=�0"����k�*�Ip�_�@�:4��ս��+>�4>��>�;���Ͼ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ua~����7�^��=��7?�0��z>���>��=�nv�ݻ��V�s����>�B�?�{�?��>!�l?��o�O�B�p�1=6M�>̜k?�s?�Qo���o�B>��?"������L��f?�
@~u@_�^?+����l���aȾC)����>���H�=�W�U>��*=2˽��`���>s�]>K�< ��>� �>���>��>RT��}�,��	��	;���� �t<�������-	�{Q���'�h㋾r�־Di��b��4S=�d��ߤŽ@V=��=:dU?޴R?�p?ެ?�wj���!>�����=ǩ��'�=͖�>��2?��K?��)?&�=�ܞ���e��Ȁ�^8���a����>��I>H�>x��>8�>�0���J>�F?>�>>��=!�$=��6;X{=&�K>��>���>�>p{8>N>�P��L���*i�%�x�,ڽ}��?*=����J��w��g拾iD��S��=4�/?�{�=\���Ͽ�����	H?S��'p�e'���>�`/?�aV?'�!>������c��]>w���vh��F>h����yk���'�(	N>Ə?��s>��>�.1�uc2�<kQ��z��_B�>��4?@`����L���j�~�9���ܾ��V>{޾>�";M������aq�"'j�2e�=6�>?_?5��GS��V�c��k���d>y>��.�"�=f�Q>��ɼR����DV��!A=�w�=�)d>�'?L�;>��j=[�>w���򏓾2�>bH>؜m>{7?6
?��v:��Ԣ�)�R�[��>���>�ĩ=�T3<7�F��#>=�C?3a>�Q�����['��V��"^E>��]>���]{(���<���mp7>mx6=,3��W$�����=��~?�}���∿�
�:K���pD?O.?E�=�)G</"�����GM����?V�@�l�?;�	�ԡV���?�?�?�	��D��=Nz�>.ӫ>�ξ��L���?W�ŽŢ�>�	��,#�DR�?@
�?�0�Mȋ��l��?>]%?/�Ӿ�g�>vx�pZ��/��g�u���#=G��>	9H?wW����O�Q>��v
?V?�\�򩤿b�ȿ�{v����>q�?��?��m��@��!@�<��>O��?MgY?�ji>Re۾v\Z����>��@?$R?n�>m7���'���?߶?篅?u*I>���?��s?ݨ�>��u�|9/���}���O�=��y;�D�>)>͛���]F�PΓ��b����j������a>��$=Q�>�����rʶ=����@G����h����>/6q>�I>l�>�� ?"��>ȣ�>�=D΋����	ɖ���K?���?B���n��U�<�ל=�]�35?R4?Mvk���Ͼ�3�>�\?�ǀ?L[?a�>g���B��!���{��P�<}L>'7�>8 �>�,��{	K>�-վy)C����>ϒ�>᣼� ھ�����<ŻZҜ>G[!?"��>+¯=�� ?M�#?D�j>(�>8aE��9��R�E�B��>��>;H?A�~?��?�Թ��Y3�����桿|�[�*:N>�x?�U? ʕ>펏�r����iE��AI�����?tg?�T彦?G2�?5�??H�A?8(f>v��'ؾj�����>? �׽�E�JG��C�6��>i�?:�?�+��s�;�'>�b����˾�a?1��?F�?�~�t~s��U̽SI�<Ӱ>���=���u֬����=�.�>�����!>[�
><ʽ��3�RG�G�Z�l��;��t>��<)ߠ�������.?�)��2a��0�=��|�o�E��>J>">�q��cuk?���J
}�j��ǈ��<L>�x͉?덿?�?�4ս�`i��c7?b;�?��?8?�莾T�ؾe����W���ɽ����$=�j�>U|5�r ��i ���謹�}�Fl��(�4�>f��>�?�?bf>� �>1������Ҿ�i�	�Z�,��$4�ւ(����},����C��}��ݻ�z����5�>.Yx�4Z�>ڿ?�Nc>\lC>�$�>�Æ;lG�>8'>l>���>Ӛb>��>'��=�٧�#d�Q�G?+��X�*�IZݾV|����3?�S?�]?����څ�Ϛ�ʭ$?�,�?�-�?�d�>�\^��|(�c?�p ?�@���� ?�h�=�ͨ���'=�[������7ƽ-����2�><ҽ�7�.H�6z����"?cB?~â:1$����J{��� k=�*�?v�(?�)���Q��o��YW���R�)��rh�S̡��%���p��珿R\���"��1~(�É$=3�*?��?���i�sʭ�[k��(?��fg>g~�>w�>`Y�>�J>ߴ	�O�1���]�E'�	�)�>��z?�C�>A)J?3}B?	�U?.�Q?��>Z��>�­�(��>��N=B��>)��>ؠ9?p�"?�'? �?�&?Z�j>���T���,ݾ9"?��?��?%?�v?\��WRս�~�8�üq�����C�NҨ=�7�;e��x����J��;�0>E�?�N��D8������=��?��	?F�?� ���T��W>��?%p?�o	?7
i�r�]���"�.��>?;z?A-��8t<���=fRB=�w=u9!�
�2=�E�=�8��nj���Ὑ$>AX>P�>{^G=z�>:�=�n�=��g>:��>�V?ى�>�z�>��������R���=��c>�,Q>��>ɶվ
����e���&f�z�>Eȏ?���?�D=�)�=�2�=ڢ����%	�b6����<�i?A ?��Q?�<�?l�<?�A#?�>��r1��WA���̣�ܻ?q�'?�^�>. �S�þS����/�=S?��?�A^�8�9�3R��i����ս��G>�M,��r�t穿��F�X�!=-��k����?�3�?�_@��.;���u����9��C�B?�˺>��>���>X���j�� ���g>h?��J?�~�>�^�?���?ж^?<ȳ>�Z�W��h����ɬ<X�>��?5�?7�?�?��}>
�?Yȭ=&���@߾L$�%��������� ��>Z�>3�y>ZK�>�q�=of+:è2�ە����o��Ր=1�>j+?��>�ߟ>-��>�B?�-�>I=���Jr��:`���˽�	e?���?%l"?�yM=����>���X'�>V��?�}�?��?�k��?B >fO���оe�L��h�>�3�>�u�>��>|��;��= �>�d�>�q˽����7�Q3]����>��)?`(`=]@˿��k�P�F�Pk���ⷼ����K�@��e�=h���8=F�������a澎(��b�þޕ��|	��v���Q��خ ?c>]>f�>'ǌ�'gy������a=y�=�r= ��=Ƣ�=�S׽K�<.ޠ��F<=�Ie<$!���Z���ʾ�e}?�I?L,?aD?��z>�b>a6���>E@|���?)U>�zK�Py���;��ʨ�թ���پ��־Jfc�W����>T�E�f�>��3>.,�=��m<a��=��t=@��=*����,=%v�=崺=��=��=�J>(>�6w?����%���Q3Q�3k罴�:?�8�>1w�=�~ƾ@?k�>>]2��̗���b��,?���?~T�?��?"vi�gb�>T���ӎ�Js�=�����?2>	��=��2����>l�J>�1K���}���3�?a�@̝??�ዿ%�Ͽ�c/>��=S�� �����1���4�ھkp���Z?��c����DZD?�ط��9�͡��:�_=s��ȱ�����HG_��.>��Q��� ~h>��q>*��=�X>�]v���D���̽lB�=��>��=;ٺ>������V=��=y|�=�[>p*�>�n?��*?�E?�k�>~�����ھT�̾Ӷ�>Ͷ�=}֤>�v�=,��=[��>J5?��E?�'K? �>	o=MB�>0D�>B�/���h�b���Ң����J{?L�?2v�>�>=�V3�ծ�x�`�s����;?�M"?�>�5�=�U����Y&�̚.�A���B�8��+=mr��PU�r����l����\�=up�>��>2�>Ty>��9>��N>��> �>�>�<�q�=�܌��ĵ<����x��=����#�<�sż�K����&��+�C������;u�;�]<��;�7�=o^�><7e>�H�>��(=튢���=>�K���F/�"y>�Ǿ��P���J��z�����߽Mg(>Tӷ=�ℽ$���t��>�>���=�j�?�,}?��N>Wa����o���;�
�����P>*�>��w�� �?�N�gC��ү�j�>Ԍ�> 4�>��W>U�*�B<����;P�ƾ�1����>~ꁾ�+�8N����Y��T��9<����b�B�E<��1?1օ����=ѻ�?n�*?T^�?�N�>�*�����dt>YN"��;�;;6�F�q�ao���/<?��?bG�>���	�%�q�ξ+�Ľ��>D!L���O��~����/�v�������>����7�Ҿ��3�f������N�B��r�i�>SN?�?]�Hڀ���N��E�uR�� u?p�g?J��>�8?�{?^����瀾��=L�n?�Y�?8��?g�
>�j�>�����>��?��?^F�?h�?G�¾P ?sz�> ���Rξ���>2��>Xs�<����=��>'_?���>�+L�B����~���Ŕ��o�<�3#=�Y|>C�>��
�e;>�C�=ί�>�C]>�Q�=�I�>�[�>��7>�̢� ��d�*?^�= Φ>��B?5G>�?�,�<l�>��)D�><���	�w5��Q2;O�;�;�R�D�>�︿gK�?R��>��*�7#&?�׾�����>.�=�"$�⹘>I!Ž6pE> ��>�r>>«<Vf:>P{=�6Ӿ�O>���/P!��=C��dR��Ѿ�z>ޜ�*�&��3�,���.�I�遵�&��j�X,��|'=�Ϫ�<�<�?����k�
�)�'r��Cg?�g�>K86?�3���슽��>��>=�>j����j��ծ��On�*��?���?&c>Y�>��W?�w?��1��3�mhZ�K�u��@���d�-�`�KǍ�a�����
�O(���_?�x?ˉA?8�<(:z>苀?:�%�x ���܊>/��U;�c�;=1Y�>���2�`�ԜӾY�þ��cF>��o?��?�?��W��Rk��8'>��:?��1??mt?X2?!�;?p���$?�a4>?�?4?[5?2�.?�
?�\1>%��=�Sû�?)=�������ҽDʽ�� 4=?�y=d	���m
<� =���<�����ټ�e;�#���b�<��8=�\�=�}�='p�>��m?f�"?�T�>.�X?k���6��s��Jg)?lb>Vw�*�R�g�L�w)���/>c8�?R��?#O?��>��)�)���˓�=�ұ>�2 >.��>J)#?1Y�=rS�:R>ܷy={'=�z*=t�q<�\���!K�V�վ%<�=�E>���>���>��ʼ�`1>1����u���h>!+��u��sֽ�O���9��_g��"�>4�I?�?�X�=P���⠓���i�Z�%?x=D?e|??��?�. >�Kʾ�4<��7F�*Z��ݥ>��<&Wݾ�]������	.�*��vm>޴���J��ۻz>:��Z�����q���O�����U�=|������gk���Ͼzm����=~>{�����'�����t%��\�B?�q�=i���:�j�;�����=_��>o?�>�7_��t���B�Dʥ�9�=?��>��e>�?��ྻ�;���c{�>CvE?�Y?r>�?��^�~q��N;���������0<�"?v|�>�=�>�H(>�^>�������K�+?����>'�?~����U���{���hG��H�>��"?'h>:��>
�H?E��>Qso?�nP?fT
?�kR>v]R�׾$�+?���?Gh�=U��(��f�V3r�-��>��U?0���(*�>�P!?O$?]]1?ʅp?f�?̇6>���4��`�>��y>�P�X���8|>��]?�>y�d?�t�?�x>�AM�K�����J>uc�=�!>4�l?�+#?���>-:�>'+�>+Z��t$1>��?�0�?:�?��B?ă4>;<�>禯=��?f���w��>�-?k>�>��? ��?��??+��>yA���{��W�H��	=G�r���<T�=�.=�����(����;[<�T�H�����:� =�ov��*,<{G�=�X�>�t>s'�� 1>	Pľ����E�@>�����5ي��;9��ش=Os>t�?��>K�#���=&�>!'�>ܹ�mf(?��?+�?a�$;heb�Q�ھ�J�)@�>��A?���=�m��d��T�u���e=C�m?rE^?oX�\����_b?m~^?F ��v=�,�þId���ˠO?�?5�J����>�}?��q?�(�>�]b��l�����F�b��k� �=���>6H��Dd��u�>Y7?�2�>.7d>�V�=Uܾ�.x��ќ�o�?4�?q�?N�?��>q�o�T`߿z���8'��?o^?z/�>�\���#?�=ݻ�о>H���F��㾚ાe+������H���&&������ӽB��=
�?�]s?-�p?%�_?�� ��3d���]����!
V��.��/���E��D��C��,n��������o����A= j4���;��7�?A4D?�&�Z{?/J<���	��HȾ�;�>�l��#�꽥��=��P��Y�h�j���� ��AW���?e��>���>A:?�f� !C��"�@2��*�e��=��>�j�>�)�>&z2;#	����y�ھؓ���R���>]^?k�W?��q?v!-��+�~k�H�'��Ӵ<��w���>���=Y��>saC���[��+��-���Z�L��DE��Ta
��K�=~�6?�C�>mK�>�?��?l��d2��D��:`�uq� ~�>��9?UX�>ߟ�>l���O&����>��j?�r�>���>SD���� ��Bp�����O�>�;�>�w�>�>J��#�\�'c����Wj3����=�_f?�:��|[��*�>�GJ?�=1;/�"<浓>g�c��� ����7����>ǿ?���=��5>#����r��x�4���V)?kr?�l���m*��U�>q<"?V��>/�>�q�?���>�����j;�"?B^?%�I??bB?>��>u$=׏��b�ɽ_J'�A�9=���>�\>ay=T��=�\���`�py���R=e�=�bȼ����O��;�ջ�g9d<�p =_�5>��ѿ��g����_���0�����5��*�m�A ׾ve6�1�Ѿ��v�" �ޚ��JD
=��I����y=����!�X;�?�#�?'����iӾ���V9t��l�E�>y��!6 �hJ��"�B��Ӿ3�	�nW¾���Ń��X�~�б����6?����.J��|$��/�Ⱦ�??"'R?�ӎ?)%
����w�*<�>�\v<��	>����Z���=)׿&�!�ֱk?��>���C����>�b�>6�R>�3>qK˾q���~�>	!?`�.?ٲ�>�)��bݿ�g濤\>@Z@z�@?'����9�x=%��>�1?/E>��8��%������>썞?�?�O,=TQX�����If?��<t
D�-�:7�=D;�=2�='��H�<>�k�>	_#�zFB�'�ڽ�|4>o��>�M�����N�+��<)�T>i�ؽIܱ�5Մ?+{\��f���/��T��U>��T? +�>W:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�܅�=q6���{���&V�~��=\��>c�>,������O��I��U��=ZK �
�̿{�$�Y ��_��+;��kν	�����4�Hm�퉣���6�XWܽ�>�'%>%�D>�͕>�Gp>Z"�>D�^?ͳn?�)�>N �=[?*��ד�W.Ǿ�Y=����V=!�ڴ��c-�u`���Ծ~�ݾv��03���z�߾�����L>;�8��v���/@��ru���U���,?R��>.���p�M�>�r�c6�����?7��5z�+���>S��1^�]Ԍ?�I?��W��jt���c�s�;`N?�|�<���SM�)^�>[oA>�A>'��>.�>O��H�@����k�(?��?�ݾQ�����h>�|@�H��zV/?��>/�N���>q'?�����F�7>��>�V�>��?L>�=U����0�M� ?hT?�9��!����>z���g9�/S�=���=��c���*��C+>w�?;������<H��<	�>+W?��>��)����7�������<=S�x?�?�	�>$vk?��B?c�<�v����S�����x=��W?�i?q�>E���l�Ͼ����&�5?΅e?P�N>�2h��龧�.��i�j�?M�n?�J?�b���\}��������]6?Sv?�q]��@���N�
�S� m�>���>@��>�8��.�>��>?��&�qe��Ɇ��A4���?�b@b;�?i C<;~�~c�=��?Y��>�|O�\�ž���~ѳ��L{=Lm�>�y���Nw��u�b�.�@�7?Z�?|�>�����4��R%>ẃ�ĉ�?��?!���&���Ӿ��y��H��ش�=��<�*�:�=bs�� E:�.��"3����t=��>�[@@�+��#�>�v���[�]"��5�m�J�������x��>��>QC�M^����q��dT�f+K�WkҾH��>Y5>�ŏ��)��w?z�W�:�hu꼞��>i6� ��>�P_�����Z՛��@><�Ք>��>$�>'�ǽ"��W֘?����f�̿����K-��#W?�C�?a��?7�?��k;3T��g�h�FO<H?�It?�@\?�	���l�ɵ9�T�k?�&���M?�P9
�ބ9�<��>��/?㔞>p�;�ڭ>}��=��	?-!>W #��ѿJ�����4��?Wo�?���Bؼ>�s�?ta?o�2��˳�؅�EVn��>	>x�? 8�=��ž��@���	��&2?mC?2�������_?|�a���p�O�-���ƽaʡ>��0��H\������]e�����!y���?�W�?I�?C���#��+%?��><���y8Ǿ��<�k�>�'�>1TN>�^��u>�(�:�A�	>��?�z�?Eq?��������>��}?�:�>-�?��=ۄ�>���==9��-@7��v!>8v�=|�;�?׵M?���>�l�=�{9��,/�,$F�NR����9�C�|�>ܑa?�L?usb>p���B�1�Nv ���̽�N1�y�޼i�B��@(�!ݽ5>3>>c�>� D��Ӿ��?Kp�8�ؿ�i��p'��54?-��>�?����t�]���;_?Gz�>�6��+���%���B�`��?�G�?<�?��׾�R̼�><�>�I�>2�Խ����X�����7>.�B?[��D��u�o�w�>���?	�@�ծ?fi��	?���P��Ja~���s7�C��=��7?�0��z>���>��=ov�׻��P�s����>�B�?�{�?��>�l?��o�L�B�3�1=7M�>Ĝk?�s?�Mo�u�j�B>�?������	L��f?�
@yu@^�^?�ῆk��껤������-�=rOY�U�<M}+�R<�<�x���/����>cc�>�'�>a�>6&Y>��(>H�+>�����[(����hA��:%���D��$ž�� H/��p�Ჰ���ξ��
�ش*<�W��~u�{�T�������=�U?a?R?!p?� ?-@{���>J���=t"�8h�=�ن>��2?NLL?=*?z��=�y��=�d���@D�����j,�>g�J>�~�>,�>�K�>S;x�H>�m>>:ހ>-��=�'=��g��=�yN>K[�>���>���>Dx>�3�>BT���$��`�`��J�����<�;�??�
=b�����	D
�uj���WF=&6?��>3����ƿ����[=F?Q��tP��o<��A>M Q?���?��i>�L �(�g�"ְ>�B>?ۉ�>a=6�;�c��Dؾ���>���>�$>�^�>��.��~>�
�^��0ݾ�U>n?>T>�g�F�]�v��] �F������>S�>pK�pÛ��~�cȀ���b>��]?���>(��e־�����[uj>���>C�ѻsF��X�>�&S�>Hn��V� n�=�(;;��><G?�6>><�o8��>��F�Oޢ���>��y>L�p>�"?�',?1��!�E�6���q|a�η#>[?ɜ�>�F>�#�PGv>�: ?�>�Ў�We������" ���>%W��ӣ��EV�J�F=����e�=1N�<_�	�:4�����<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾRh�>wx��Z�������u���#=U��>�8H?�V����O�d>��v
?�?�^�ߩ����ȿ6|v����>X�?���?h�m��A���@����>:��?�gY?foi>�g۾/`Z����>һ@?�R?�>�9���'���? ߶?ׯ�?��>�x?ux�?�?*Ä�(���]�䂖�ģ	=s>�^_;Ki�>����=P�ҡ��S����(�=� �g2�>��=�϶>1��־D�=��/5޾J���U!�>+]>Cl�>��><D�>A�>���>��#>�*�s���rs�u�J?��?��;<o��u<H��=Zr]�h�?"3?#[��	jо���>��Z?O�}? �Z?�;�>�"��Қ��¿�ѯ��נ<�A<>�7�>-��>��T�_SP> �پ
�M�j2�>���>�ӻ'۾}�����q�~M�>��"?���>��=y� ?\�#?��k>鮲>�JE�?��->E��x�>���>$9?��}?��?���i3�5뒿'JA[��<N>\�x?�.?�7�>Wm��w���LR�EM��Y��Mk�?F9g?�d���?m3�?�c??@aA?Spf>L�(�׾;��$R�>�T?cd���+j�~U��������>��R?�,?�u=b�ܾ���ۭ��D��l�>r�c?�()? -M��脿��9�ٕ�<���=	�8=��D<M k<%��=��Z>7J
=��N>�>��E>�H$�GtT��QL=��">�b�>��<ݒ5�S1�=P�&?6d�=.g��991=\�Q��H#��R>w��>��S���D?*�.� '��ݪ���֜�8yi�0�v?ς�?g�?M畽J�V�QP?�Ǎ?3r�>��>p�Ӿ� ��ؾ�wѽ�{��x.�e.�=�p�>�Q�<$e���C�������ً�^��������>��?�'?�x?���=���>T�Ⱦ���l���I�`���.k���!�5�U�Y3@�l<m�(����=I����̾�sN�>���ߐ�>W�>}+>9-S>���>?�:�4A>��>tK'>�t�>ބ>wƆ>M>!�
=�<ӽ�KR?������'�}�������2B?�qd?p1�>i�<������/�?���?�r�?y<v>l~h��,+��m?@;�>����p
?�Q:=���D�<U����s/��Z����>P׽x!:��M��mf�nj
?>/?K/����̾[7׽tq��?��=�r�?_-5?�*���K���W�O�^�WJ�w6F��E������v���l�^O���.���~��M����=L$?+�?-$��q����+k��,�ߟT>��>\��>{��>��@>���[.�/�P��_*��A�����>��k?k\�>��7?�&E?��>?Z�v?!��>8�=)+��p�7>\��=MF$?��?��?v?+c ?Q!?�%U?�z�>����޾Z���?��-?P�!?��>��?rC�N_k��^�-L�Y���9��=��>D���5���> ����<�� =�c?2G��o;��}󾹋>!X8?���>��>����<���pe= ��>~�>��>������l�q���"��>�#~?��
��X�<��*>zr�=L�߼������=M�޼���=m�����4�;��=��q=��
:�A�:�B	<��;���<&�>i
?�?�>�-�>��������R�Ma�=r�b>c�M>�>4�����5.���5g�x]q>N[�?��?�Ij=G��=��>�b���þg������]�<�)?��$?�HR?e֎?sw8?��"?Y >�/� ���ׄ�������?�0?���>l��6¾���i��oj?�?[wg��ͽ� ����+���t,>6����r��?"���=u\�\)۽\��?���?����<<�~��c�����pc?Џ�>W��>���>�+7��Ђ��0�̛�>_	?e�\?젾>*�O?��|?�X?2�5>�>7�'��^���1�<_�.>y�=?���?||�?j�n?Ɉ�>2��=7c%�nܾ���!A�C��­|���=WZ>�ʍ>���>�ص>>�=�tѽQYO�F}��=��{>z��>�_�>�>&�>W��;�F?��>�찾C �������:]*��Ek?ܗ?��,?S�=V���%�L例��>�W�?U��?� ?�d^����=G�D������q��h�>k?8�>��b�h��<�1>�c�>W��>y�-��F���=g?6F?1��=}x��ve����wڞ�1	���5�������ͽ(�V���=�p����q��ͫ�����ԓ¾y��B>ҾC�����o���>�W�=��>���=�=T??�67�<hId<�� ��-=��˼:-j:A���F�t�/���W���v�<;�8<@�W�P�ʾv}?.'I?vy+?�jC?oy>�x>ň6�C��>� ���:?�V>M�N�������;�n㨾yՔ�'kؾ�׾D�c�ķ��t�>UjF��>�!3>���=FĎ<�B�==�r=o��=���� +=�C�=�]�=���=���=�G>,'>�6w??��������4Q�dZ罗�:?�8�>�{�=�ƾV@?@�>>�2�������b��-?m��?�T�?3�?5ti��d�>��n⎽�p�=Q���O=2>���=��2�}��>T�J>����J��
���4�?��@��??�ዿ٢Ͽ�`/>��x>6��>#f_�L�B���I�?��-_�Ƣ?1�1�W�����>���>cJ����[���g;�=]M(>(���z���B�=Z0e�>3ݽ׃�>�+?�x�>���=i����~=�׼=* �>��v=����]b=��ܽrê���>f<�>� >�h�>��?�0?#^d?��>�%f���˾�L¾Cl�>�C�=���>\�=�oK>'F�>Z�5?�PC?�sL?�Ƴ>Vc�=���>෦>��,�Ҳk��(����*$�<�ʇ?��?�8�>� <�:��<���<��U���?w�/?g�?甛>�h�*� ���N�uU'������;,�;Z*���n�=�k�=uY,��"�=��>f|;?��?��>A�\>���>���> �i=��!�-<�<�}7�����q���7��=`�8���G�{�t���=H&l�jx<ʺȻ�����=��=�G>t�>�8�>K�e>�C�>pQL=#?����K>�-���+M�yeT>$��T^N���W�`��g�A����B>�>q>�8	=������>��#>��=K9�?�?ų>�?̽i���^���cx�o����J�<e6�>�5���-8��gO�U�Y�����A~�>%��>�?��>��3��]�n�4=V����"��$q?�#���7��s��}����Ž�7���	�G�,�k>��v?����'>8q?�?|��?��>�h%�a�����=S���l�T�ݣC�W̘���D�/�?��>o0�>��1�&`�)?̾�	����>�I�|�O�
���ޥ0�N���Ʒ�b��>,	����оD3�Xf�������B�"Lr���>��O?�?VBb�HT��`PO��������s?<vg?T�>�H?�=?$ס�%j�rv��l��=��n?��?>:�?{>dd>e���%�?�f?�֛?uA�?�P?<B�Y��>I��=v�>o�u��Cn>l�i>U���%�m=%5#?��?�?���;R����ԲҾrF��'��V�	>Q>�>=>z�>S�='5P>�\�=���=�E}>�:�>�<�>>��>y��><�x�2���H?[��>�f�>ֿ)?���>J�Ž3*����!>��k�� ���WM�ա#�l���(���Qq<z��=�X�=v]�>)~ſ[z�?ͪ�>�f-��,?-�������MGs>��W>��ͽ�u?���>q�>��>���>���=��>�L4>�GӾ�z>���Mi!��1C�τR���ѾЇz>B���-&���3����HI��p���d�9j��/���==��p�<|E�?l|��t�k�w�)�����}�?�Z�>�6?
Ԍ�Rሽ��>��>\ˍ>�R��2����č�&^���?^��?�Hc>$�>A�W?:�?�Z1���2�gZ�.�u��A�P�d��`��鍿렁��
��S��>�_?u�x?�|A?g��<$*z>��?��%���>r/�'%;�7�<=PG�>����`a�>�ӾH�þ7G�IF>E�o?��?s;?VV���=�>rTD?�K?��?�qk?dC#?�wE�x�>q��=�?-�>uS?Rd?}: ?�x2>��2>,�M=�l'=_��.휾b��������X�=WC�=$5�d��=���=b�k�@�����<��+>�)�������ⅼ�p=a��=��>e|Y?6��>>��P?����
��������S?Leg>�꫽���U�z��k���wD>`؉?��?�C?B�C>=�V��>D���>8�>W?>e�>�f�>�b����ݾ3dY=o.�>´�>A�>T�:=jo[��]�Y�a�̋Q=ޡd>Q��>�}>�'��d9&>$����uz�8�d>��P�|����T��G�w1�$mv����>��K?}�?`��=V�� !��c�e�O)?��;?�IM?��?��=H�۾@:���J��L�\��>f��<			�߯��#!����:���;��t>�ߞ��J��ۻz>:��Z�����q���O�����U�=|������gk���Ͼzm����=~>{�����'�����t%��\�B?�q�=i���:�j�;�����=_��>o?�>�7_��t���B�Dʥ�9�=?��>��e>�?��ྻ�;���c{�>CvE?�Y?r>�?��^�~q��N;���������0<�"?v|�>�=�>�H(>�^>�������K�+?����>'�?~����U���{���hG��H�>��"?'h>:��>
�H?E��>Qso?�nP?fT
?�kR>v]R�׾$�+?���?Gh�=U��(��f�V3r�-��>��U?0���(*�>�P!?O$?]]1?ʅp?f�?̇6>���4��`�>��y>�P�X���8|>��]?�>y�d?�t�?�x>�AM�K�����J>uc�=�!>4�l?�+#?���>-:�>'+�>+Z��t$1>��?�0�?:�?��B?ă4>;<�>禯=��?f���w��>�-?k>�>��? ��?��??+��>yA���{��W�H��	=G�r���<T�=�.=�����(����;[<�T�H�����:� =�ov��*,<{G�=�X�>�t>s'�� 1>	Pľ����E�@>�����5ي��;9��ش=Os>t�?��>K�#���=&�>!'�>ܹ�mf(?��?+�?a�$;heb�Q�ھ�J�)@�>��A?���=�m��d��T�u���e=C�m?rE^?oX�\����_b?m~^?F ��v=�,�þId���ˠO?�?5�J����>�}?��q?�(�>�]b��l�����F�b��k� �=���>6H��Dd��u�>Y7?�2�>.7d>�V�=Uܾ�.x��ќ�o�?4�?q�?N�?��>q�o�T`߿z���8'��?o^?z/�>�\���#?�=ݻ�о>H���F��㾚ાe+������H���&&������ӽB��=
�?�]s?-�p?%�_?�� ��3d���]����!
V��.��/���E��D��C��,n��������o����A= j4���;��7�?A4D?�&�Z{?/J<���	��HȾ�;�>�l��#�꽥��=��P��Y�h�j���� ��AW���?e��>���>A:?�f� !C��"�@2��*�e��=��>�j�>�)�>&z2;#	����y�ھؓ���R���>]^?k�W?��q?v!-��+�~k�H�'��Ӵ<��w���>���=Y��>saC���[��+��-���Z�L��DE��Ta
��K�=~�6?�C�>mK�>�?��?l��d2��D��:`�uq� ~�>��9?UX�>ߟ�>l���O&����>��j?�r�>���>SD���� ��Bp�����O�>�;�>�w�>�>J��#�\�'c����Wj3����=�_f?�:��|[��*�>�GJ?�=1;/�"<浓>g�c��� ����7����>ǿ?���=��5>#����r��x�4���V)?kr?�l���m*��U�>q<"?V��>/�>�q�?���>�����j;�"?B^?%�I??bB?>��>u$=׏��b�ɽ_J'�A�9=���>�\>ay=T��=�\���`�py���R=e�=�bȼ����O��;�ջ�g9d<�p =_�5>��ѿ��g����_���0�����5��*�m�A ׾ve6�1�Ѿ��v�" �ޚ��JD
=��I����y=����!�X;�?�#�?'����iӾ���V9t��l�E�>y��!6 �hJ��"�B��Ӿ3�	�nW¾���Ń��X�~�б����6?����.J��|$��/�Ⱦ�??"'R?�ӎ?)%
����w�*<�>�\v<��	>����Z���=)׿&�!�ֱk?��>���C����>�b�>6�R>�3>qK˾q���~�>	!?`�.?ٲ�>�)��bݿ�g濤\>@Z@z�@?'����9�x=%��>�1?/E>��8��%������>썞?�?�O,=TQX�����If?��<t
D�-�:7�=D;�=2�='��H�<>�k�>	_#�zFB�'�ڽ�|4>o��>�M�����N�+��<)�T>i�ؽIܱ�5Մ?+{\��f���/��T��U>��T? +�>W:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�܅�=q6���{���&V�~��=\��>c�>,������O��I��U��=ZK �
�̿{�$�Y ��_��+;��kν	�����4�Hm�퉣���6�XWܽ�>�'%>%�D>�͕>�Gp>Z"�>D�^?ͳn?�)�>N �=[?*��ד�W.Ǿ�Y=����V=!�ڴ��c-�u`���Ծ~�ݾv��03���z�߾�����L>;�8��v���/@��ru���U���,?R��>.���p�M�>�r�c6�����?7��5z�+���>S��1^�]Ԍ?�I?��W��jt���c�s�;`N?�|�<���SM�)^�>[oA>�A>'��>.�>O��H�@����k�(?��?�ݾQ�����h>�|@�H��zV/?��>/�N���>q'?�����F�7>��>�V�>��?L>�=U����0�M� ?hT?�9��!����>z���g9�/S�=���=��c���*��C+>w�?;������<H��<	�>+W?��>��)����7�������<=S�x?�?�	�>$vk?��B?c�<�v����S�����x=��W?�i?q�>E���l�Ͼ����&�5?΅e?P�N>�2h��龧�.��i�j�?M�n?�J?�b���\}��������]6?Sv?�q]��@���N�
�S� m�>���>@��>�8��.�>��>?��&�qe��Ɇ��A4���?�b@b;�?i C<;~�~c�=��?Y��>�|O�\�ž���~ѳ��L{=Lm�>�y���Nw��u�b�.�@�7?Z�?|�>�����4��R%>ẃ�ĉ�?��?!���&���Ӿ��y��H��ش�=��<�*�:�=bs�� E:�.��"3����t=��>�[@@�+��#�>�v���[�]"��5�m�J�������x��>��>QC�M^����q��dT�f+K�WkҾH��>Y5>�ŏ��)��w?z�W�:�hu꼞��>i6� ��>�P_�����Z՛��@><�Ք>��>$�>'�ǽ"��W֘?����f�̿����K-��#W?�C�?a��?7�?��k;3T��g�h�FO<H?�It?�@\?�	���l�ɵ9�T�k?�&���M?�P9
�ބ9�<��>��/?㔞>p�;�ڭ>}��=��	?-!>W #��ѿJ�����4��?Wo�?���Bؼ>�s�?ta?o�2��˳�؅�EVn��>	>x�? 8�=��ž��@���	��&2?mC?2�������_?|�a���p�O�-���ƽaʡ>��0��H\������]e�����!y���?�W�?I�?C���#��+%?��><���y8Ǿ��<�k�>�'�>1TN>�^��u>�(�:�A�	>��?�z�?Eq?��������>��}?�:�>-�?��=ۄ�>���==9��-@7��v!>8v�=|�;�?׵M?���>�l�=�{9��,/�,$F�NR����9�C�|�>ܑa?�L?usb>p���B�1�Nv ���̽�N1�y�޼i�B��@(�!ݽ5>3>>c�>� D��Ӿ��?Kp�8�ؿ�i��p'��54?-��>�?����t�]���;_?Gz�>�6��+���%���B�`��?�G�?<�?��׾�R̼�><�>�I�>2�Խ����X�����7>.�B?[��D��u�o�w�>���?	�@�ծ?fi��	?���P��Ja~���s7�C��=��7?�0��z>���>��=ov�׻��P�s����>�B�?�{�?��>�l?��o�L�B�3�1=7M�>Ĝk?�s?�Mo�u�j�B>�?������	L��f?�
@yu@^�^?�ῆk��껤������-�=rOY�U�<M}+�R<�<�x���/����>cc�>�'�>a�>6&Y>��(>H�+>�����[(����hA��:%���D��$ž�� H/��p�Ჰ���ξ��
�ش*<�W��~u�{�T�������=�U?a?R?!p?� ?-@{���>J���=t"�8h�=�ن>��2?NLL?=*?z��=�y��=�d���@D�����j,�>g�J>�~�>,�>�K�>S;x�H>�m>>:ހ>-��=�'=��g��=�yN>K[�>���>���>Dx>�3�>BT���$��`�`��J�����<�;�??�
=b�����	D
�uj���WF=&6?��>3����ƿ����[=F?Q��tP��o<��A>M Q?���?��i>�L �(�g�"ְ>�B>?ۉ�>a=6�;�c��Dؾ���>���>�$>�^�>��.��~>�
�^��0ݾ�U>n?>T>�g�F�]�v��] �F������>S�>pK�pÛ��~�cȀ���b>��]?���>(��e־�����[uj>���>C�ѻsF��X�>�&S�>Hn��V� n�=�(;;��><G?�6>><�o8��>��F�Oޢ���>��y>L�p>�"?�',?1��!�E�6���q|a�η#>[?ɜ�>�F>�#�PGv>�: ?�>�Ў�We������" ���>%W��ӣ��EV�J�F=����e�=1N�<_�	�:4�����<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾRh�>wx��Z�������u���#=U��>�8H?�V����O�d>��v
?�?�^�ߩ����ȿ6|v����>X�?���?h�m��A���@����>:��?�gY?foi>�g۾/`Z����>һ@?�R?�>�9���'���? ߶?ׯ�?��>�x?ux�?�?*Ä�(���]�䂖�ģ	=s>�^_;Ki�>����=P�ҡ��S����(�=� �g2�>��=�϶>1��־D�=��/5޾J���U!�>+]>Cl�>��><D�>A�>���>��#>�*�s���rs�u�J?��?��;<o��u<H��=Zr]�h�?"3?#[��	jо���>��Z?O�}? �Z?�;�>�"��Қ��¿�ѯ��נ<�A<>�7�>-��>��T�_SP> �پ
�M�j2�>���>�ӻ'۾}�����q�~M�>��"?���>��=y� ?\�#?��k>鮲>�JE�?��->E��x�>���>$9?��}?��?���i3�5뒿'JA[��<N>\�x?�.?�7�>Wm��w���LR�EM��Y��Mk�?F9g?�d���?m3�?�c??@aA?Spf>L�(�׾;��$R�>�T?cd���+j�~U��������>��R?�,?�u=b�ܾ���ۭ��D��l�>r�c?�()? -M��脿��9�ٕ�<���=	�8=��D<M k<%��=��Z>7J
=��N>�>��E>�H$�GtT��QL=��">�b�>��<ݒ5�S1�=P�&?6d�=.g��991=\�Q��H#��R>w��>��S���D?*�.� '��ݪ���֜�8yi�0�v?ς�?g�?M畽J�V�QP?�Ǎ?3r�>��>p�Ӿ� ��ؾ�wѽ�{��x.�e.�=�p�>�Q�<$e���C�������ً�^��������>��?�'?�x?���=���>T�Ⱦ���l���I�`���.k���!�5�U�Y3@�l<m�(����=I����̾�sN�>���ߐ�>W�>}+>9-S>���>?�:�4A>��>tK'>�t�>ބ>wƆ>M>!�
=�<ӽ�KR?������'�}�������2B?�qd?p1�>i�<������/�?���?�r�?y<v>l~h��,+��m?@;�>����p
?�Q:=���D�<U����s/��Z����>P׽x!:��M��mf�nj
?>/?K/����̾[7׽tq��?��=�r�?_-5?�*���K���W�O�^�WJ�w6F��E������v���l�^O���.���~��M����=L$?+�?-$��q����+k��,�ߟT>��>\��>{��>��@>���[.�/�P��_*��A�����>��k?k\�>��7?�&E?��>?Z�v?!��>8�=)+��p�7>\��=MF$?��?��?v?+c ?Q!?�%U?�z�>����޾Z���?��-?P�!?��>��?rC�N_k��^�-L�Y���9��=��>D���5���> ����<�� =�c?2G��o;��}󾹋>!X8?���>��>����<���pe= ��>~�>��>������l�q���"��>�#~?��
��X�<��*>zr�=L�߼������=M�޼���=m�����4�;��=��q=��
:�A�:�B	<��;���<&�>i
?�?�>�-�>��������R�Ma�=r�b>c�M>�>4�����5.���5g�x]q>N[�?��?�Ij=G��=��>�b���þg������]�<�)?��$?�HR?e֎?sw8?��"?Y >�/� ���ׄ�������?�0?���>l��6¾���i��oj?�?[wg��ͽ� ����+���t,>6����r��?"���=u\�\)۽\��?���?����<<�~��c�����pc?Џ�>W��>���>�+7��Ђ��0�̛�>_	?e�\?젾>*�O?��|?�X?2�5>�>7�'��^���1�<_�.>y�=?���?||�?j�n?Ɉ�>2��=7c%�nܾ���!A�C��­|���=WZ>�ʍ>���>�ص>>�=�tѽQYO�F}��=��{>z��>�_�>�>&�>W��;�F?��>�찾C �������:]*��Ek?ܗ?��,?S�=V���%�L例��>�W�?U��?� ?�d^����=G�D������q��h�>k?8�>��b�h��<�1>�c�>W��>y�-��F���=g?6F?1��=}x��ve����wڞ�1	���5�������ͽ(�V���=�p����q��ͫ�����ԓ¾y��B>ҾC�����o���>�W�=��>���=�=T??�67�<hId<�� ��-=��˼:-j:A���F�t�/���W���v�<;�8<@�W�P�ʾv}?.'I?vy+?�jC?oy>�x>ň6�C��>� ���:?�V>M�N�������;�n㨾yՔ�'kؾ�׾D�c�ķ��t�>UjF��>�!3>���=FĎ<�B�==�r=o��=���� +=�C�=�]�=���=���=�G>,'>�6w??��������4Q�dZ罗�:?�8�>�{�=�ƾV@?@�>>�2�������b��-?m��?�T�?3�?5ti��d�>��n⎽�p�=Q���O=2>���=��2�}��>T�J>����J��
���4�?��@��??�ዿ٢Ͽ�`/>��x>6��>#f_�L�B���I�?��-_�Ƣ?1�1�W�����>���>cJ����[���g;�=]M(>(���z���B�=Z0e�>3ݽ׃�>�+?�x�>���=i����~=�׼=* �>��v=����]b=��ܽrê���>f<�>� >�h�>��?�0?#^d?��>�%f���˾�L¾Cl�>�C�=���>\�=�oK>'F�>Z�5?�PC?�sL?�Ƴ>Vc�=���>෦>��,�Ҳk��(����*$�<�ʇ?��?�8�>� <�:��<���<��U���?w�/?g�?甛>�h�*� ���N�uU'������;,�;Z*���n�=�k�=uY,��"�=��>f|;?��?��>A�\>���>���> �i=��!�-<�<�}7�����q���7��=`�8���G�{�t���=H&l�jx<ʺȻ�����=��=�G>t�>�8�>K�e>�C�>pQL=#?����K>�-���+M�yeT>$��T^N���W�`��g�A����B>�>q>�8	=������>��#>��=K9�?�?ų>�?̽i���^���cx�o����J�<e6�>�5���-8��gO�U�Y�����A~�>%��>�?��>��3��]�n�4=V����"��$q?�#���7��s��}����Ž�7���	�G�,�k>��v?����'>8q?�?|��?��>�h%�a�����=S���l�T�ݣC�W̘���D�/�?��>o0�>��1�&`�)?̾�	����>�I�|�O�
���ޥ0�N���Ʒ�b��>,	����оD3�Xf�������B�"Lr���>��O?�?VBb�HT��`PO��������s?<vg?T�>�H?�=?$ס�%j�rv��l��=��n?��?>:�?{>dd>e���%�?�f?�֛?uA�?�P?<B�Y��>I��=v�>o�u��Cn>l�i>U���%�m=%5#?��?�?���;R����ԲҾrF��'��V�	>Q>�>=>z�>S�='5P>�\�=���=�E}>�:�>�<�>>��>y��><�x�2���H?[��>�f�>ֿ)?���>J�Ž3*����!>��k�� ���WM�ա#�l���(���Qq<z��=�X�=v]�>)~ſ[z�?ͪ�>�f-��,?-�������MGs>��W>��ͽ�u?���>q�>��>���>���=��>�L4>�GӾ�z>���Mi!��1C�τR���ѾЇz>B���-&���3����HI��p���d�9j��/���==��p�<|E�?l|��t�k�w�)�����}�?�Z�>�6?
Ԍ�Rሽ��>��>\ˍ>�R��2����č�&^���?^��?�Hc>$�>A�W?:�?�Z1���2�gZ�.�u��A�P�d��`��鍿렁��
��S��>�_?u�x?�|A?g��<$*z>��?��%���>r/�'%;�7�<=PG�>����`a�>�ӾH�þ7G�IF>E�o?��?s;?VV���=�>rTD?�K?��?�qk?dC#?�wE�x�>q��=�?-�>uS?Rd?}: ?�x2>��2>,�M=�l'=_��.휾b��������X�=WC�=$5�d��=���=b�k�@�����<��+>�)�������ⅼ�p=a��=��>e|Y?6��>>��P?����
��������S?Leg>�꫽���U�z��k���wD>`؉?��?�C?B�C>=�V��>D���>8�>W?>e�>�f�>�b����ݾ3dY=o.�>´�>A�>T�:=jo[��]�Y�a�̋Q=ޡd>Q��>�}>�'��d9&>$����uz�8�d>��P�|����T��G�w1�$mv����>��K?}�?`��=V�� !��c�e�O)?��;?�IM?��?��=H�۾@:���J��L�\��>f��<			�߯��#!����:���;��t>�ߞ�d7���o>����ﾁ}o�m�R����4ݫ=+�pq	<W��wQؾ�c��Oǰ=��>� ƾs%�L����j���I?��=�����h�縱��>�j�>���>5���ZIX��;<��°����="��>f8>�������F�{L�] �>ĽE?��^?�Ń?�����r��uB�A���,K����v�?���>�5?�B>���=SO��T���?e�JhG���>��>3���eG��螾AY��1$��\�>�?.>K�?נR?K?��`?i�)?�0?,y�>ﶽ=����#!?<��?�<j��7l��8�\P2�#�?�d4?�����_�>�7	?z-?�)?�SS?\??��=jY�ڱK���>��l>�>Z��ť�S�Z>(C?���>(O?J9|?_!>�#�2��ܒ��3>�dC>��3?�Y?;�?��>}��>y�����=֠�>�c?1�?F�o?�s�=;�?}B2>L��>��=v��>���>h?
XO?��s?g�J?���>Sύ<�$���9��<5s�<�P�st�;��H<�y=����t��Z��C�<�;�m��>�����D�搼��;�^�>�Tu>u�����.>����ˀ�c��>���=gᦾ�׊�<h'�I�=�� >M��>��>��$�n��Z�>��>f���5?�E?T�>C�J�lKg�#ʾ�i"�ew�>��'?�R=��s�������Y�z�>�ւ?�^U?Y����
��<a?�%U?p�p3�+����J��;��P-V?�e�>�J����>�w?��Y?�v�>�+��Rg�x���#;W�ޔj����=ͳ>s��i�i�_��>��'?���>Up>W�>xy�I�q�����?�u�?\��?b;�?�'>�.r���1�����-�q?��?l����(?�������h]�}�I������Ϧ�y���Uʘ����'�0T�n:ѽ���=�?/�v??�j?�N?��پ��^��t\�Rt���^������"���T�a�>��?D�˔j���b��8��þ<ZJ�}dA�>s�?��Y?�yN���?y6��i�&���b�Y)�>$���%:Y�q03���j���?=`,"=��l���
��Ւ�X�?^��>�o�>��.?�[g�@��m*!��@��_�fЖ>�N=��>u��>;�ͽ�G�.)�B� ��t��$��b:v>Oyc?�K?�n?�q��,1�慂�r�!�K�/�5f����B>�r>���>�W�����8&��V>���r�����u����	�i�~=2�2?&�>ǲ�>�N�?^?�y	��i���bx�m�1���<y0�>)i?�?�>a�>rн�� �i��>Jqk?{��>;�>���}���s���5½�>!Xo>�e?�T�>�Cǽ��T��ߗ�"����g&���6>Ref?̮]�A���<�>>�oU?t导Q��]�>��{�l`��,׾9&�}�">�	(?�7=��=KѾ�����P����a�%?�z'?Q�����(��υ>9�
?�b?���>o��?Z۽=�}���z�]<�>>�m?k�Q?%?I?p̂>�ڍ��=��tT׽%$���qa=Qm'>�\>�� �>��</<�����d�=x/�=�Լ��<�2�����[�=�>>�p>~п��I�B���@A�^I��u��om���15=DX������%B�(P�}��������������6"��"�(5=�"�?��?_������(��
����ؾ)]?���q�����Y$#�@Ϯ���r!r��H�3T���$y��fI�ی'?ȵ��۰ǿ����. ܾj ?�  ?p�y?����"�b~8�0� >�C�<O���_��*�����οS���^?F��>�������"�>�݂>�7Y>��q>$I��y���l��<��?�f-?��>s�q���ɿ�p���_�<s��?5�@��A?��)������΄=�.�>�S
?TDI>۪)�*6"��͞��>�a�?���?��c=.)X�Tr���X?�^�<O9�U��+�=u�R=4Dc<p��5�7>��>J�佸�E�8��4�S>��>2Bg�/� @"�[�<��3>����sؽ�Ԅ?�x\�lf�c�/�8T��NR>��T?y.�>�7�=��,?�6H��|Ͽt�\�D)a?�0�?��?(�(?Aܿ�6՚>��ܾ��M?�E6?��>�d&�q�t��w�=gE�{B����㾤&V���=��>�>R�,�ψ��O�������=6���H(Ŀ��Q�������C-�s�E�j�K��
���3Z���������XW�=C6s>��>�V�></>�%O?ya?�Ͳ>?��=ˌ���å��Ⱦ�_%>��Y��Kz�������Ľ��f�4�e�׾���Z-��,�抢��g4�R��=��L�����?*��z���K�Zf@?��=Tp���9���h��g���Ծ��= :'��*�Ov+���_�eU�?fqY?�-��bm�b�!Ľ�	��=?S{*���	�A)�����;7*�����=�/�>��=�� ���B��YS�P0?��"?���Z3s�L�K>.�>�3=$�,?�+?��R�_��>\�,?r�����ܽ��=��=D@�>F(�>��#>Y�����׽�+#?w�X?��2����[�o>������/�=���=4���7<$�='5<1���>=�\�ñ�;CmU?w��>9�"�zv�e9q�/�G��E<��o?��?��>l�m?�D?˕J=EK����\��L�1�j= IX?�Fj?%�>=��H�۾�����-?�\?Oq>�1W�#"��^*�Dz���?Scv?�Q?_-ͼ<�y�z쎿[�����:?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?s�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������{��=����?>��?����F�<O��o�q��-��n/=9�U=s�F��N�V)ﾺm5�!ƾ0��T����(��0��>P�@}-���>�u� ࿇ο�!���۾�w�Q|?�ӕ>�	սP.��ǐi�Ԓs�G��I�����ޣ>~�>�욽��a0{�E�:��ˏ����>A��ω>$�T��)��T���`�=<��>���>'9�>�:��%U��Z�?	)���ο���� r���W?�-�?��??�?U�<�xs�c�x�*o6��F?v*t?�Y?�90��_�fF�$�g?DH���P��T��4��y>�W-?Q�>�L&��õ=]�>V�?��r>�#��f¿垳�^L쾝�?�;�?с߾��>}l�?}y:?�$�'��������0�����L?�J>s���#��-7�F�t��?�3?��E�]�_?(�a�M�p���-���ƽ�ۡ>��0��e\��M�����Xe����@y����?M^�?i�?ֵ�� #�d6%?�>b����8Ǿ��<���>�(�>*N>DH_���u>����:�
i	>���?�~�?Pj?���������U>�}?v�>�ބ?��=�3�>�y�=�d���"��:%>4=�=�&D�V'?܁N?v��>SO�=��=��T/�=FE�ʧP���"2C�[��>�b?&M?��Z>|�Ľ�_3�|� �ѽK,�8W�7>����I�i�7>��?>��>S2F���Ӿ��?Px��ؿ�T���'��A4?��>�?����	t�Ѽ�t,_?[��>����(��21��,�����?�H�?��?�׾�;˼c?>��>�]�>�AԽ��N���Hx8>�uB?���3��q{o��ֆ>���?m�@�ɮ?��h��	?���P��Va~�,���7���=��7?�0�F�z>���>��=�nv�ڻ��?�s����>�B�?�{�?��>�l?��o�B�B���1=RM�>؜k?�s?�Mo�^�ӱB>o�?)�������K��f?��
@vu@x�^?&�տ����j喾���_��s:�=�e�>E~�.b���
\>e?�
���ks�>ļ�>��o>�A�>ρ�>��->*�=�ރ�%|#�E��-���.����{�۾r�]��)3������4.�G4���ޭ��y����q��=T�3�3�ý�C>��=�FV?�P?��m?��>h��>�(��,=�s)�3ņ=H�>|�1?aIL?Ԧ*?U��=D����Te�I}���	��3����>D�G>��>)��>�M�>��;6�N> ;> :�>j]>6�6=z�j;�=#�N>(��>���>KƷ>ep>>��&>c���b����g�����k���Aע?{#��^eM��;���I���!��@�=Ԏ/?��	>4e��BWϿ����LG?�������!,�B	>�0?=fX?�>���O�!�>\�/hm��G>�[��}b\���)���J>iV?�'y>I;�>ɪ(�y<���>��Iվ���>=�J?�	w��H��^�e���R�h���%>��>v=�=[�.��ԓ�;D~�񿜾�?a>/M?���>����¾�׾�ｾ� �>{�=3�=�q�=ݮ�>�W�=Cwd���	�R�>�qh�E��=#
?�v.>0�=a8�>����Y�Y����>�	H>n�)>�+=?ir%?���#�~�"�����6��Qj>dL�>���>Ϧ>BJ�㚴=M��>��i>B@��>���X��_=��WR>T\���^��Bg����=�g��yh>��=����<A���<�~?k��䈿�뾌^��JmD?�+?���=�HF<��"� ���G����?K�@�k�?��	��V�i�?WA�?�	��K��=�|�>�׫>�ξu�L�k�?ƽ�Ƣ��	�+,#�R�?�?�/�"ʋ�!l��8>�^%?կӾ"w�>kh&��y��N�h��0P��=>$+-> rD?�b	� %D�h���U ?��?����ě�J\ѿ��z�F�?S/�?c��?#���������x�	?̰�?Yܐ?�D>�n&�r��;�<>t�?�96?"E?)���M����>A-�?��?�#N>@�?�q?���>^ �2.�����ފ�/��=����ߘ>��>m����E�K6���Ĉ�
g�� �ni>�G0=�կ>b���b���s(�=���� ���r�3�>�l>��D>U��>"�?C>�>�<�>UE�<t܋�l��-��JDF?yA�?E���h����<C��=D����	?{�@?R���$Ĩ���>>NE?��~?��[?ȯ�>������������o��<&�->i�>e��>*����i>������K�A>�w�>JV>�@��i�A��v�B@�>�D?uf�>�Ǜ=B� ?��#?��i>+1�>�v=�T���p�F�ぽ>���>{-?�?��?a@���_2���������=X�4^Z>��y?�?R��>9����ҙ�f�����Q�t�E�!]�?�Ic?��佀?�w�?�C?�@?�Tb>8��!վ���o��>��?���>���oY�ou���?�z+?���>�~�>f}2�2A�=�I)�����?Ǟ}?�2l?�~�ʼ��~%A�M�=HW���r�<��$���7=]��>`=Z�����&=�E�>��>AF�0+2���r=}�=�P�>Ѫ�=A�Nh�;�<,?�G�SӃ���=��r��uD���>3;L>������^?5v=�?�{�0��@x���U�
 �?|��?zj�?�	���h��%=?��?S?&�>vK��	޾7��ZYw�#~x��x�n�>���>�l��ŏ�������F���ƽ�g��C�>9�>}�?� ?�2V>��>7X��!�(��������]���"�5���.����c����O�Hʻ�����Zt�FT�>�؝�ث�>��?d0i>���>��>e/���>PiZ>S�r>K�>�ri>�6>�=�=���9{�D�P?�ݾ4�K��J�����>?�b?���>�䜾U�7�����?/�I?[|?��>J`n�;�@��	?3v?2lm��?���{%���];�9���:�U> 4=�5=��=d�����H�Ѷ��U?�^'?ܑ;�G>���¾8}����o=�H�? �(?j�)���Q�b�o�ʪW��S��;��g�_����$��p��돿�[��� ���(��h*=Q�*?��?ƃ�n�&���k��?��f>���>�,�>Ӿ>��I>ѽ	���1�5^�T'������`�>�b{?=i�>�BI?
I<?H�P?�CM?Z�>4y�>���Y^�>+�<t��>���>m9?��-?o90?8�?�+?Vc>k������ kؾ�?�?�	?K?.�?����p����^��h�h��x�F���Ɂ=�P�<iVؽ�2s��V=��S>��'?l?��'�BJ�kw�>2�*?���>��N>'7ž�b�=��ͽ��>4�.?���>R^�/���� ���??�`�?� ���O���=��>RF�������>gk<�P7=2��=h�
��^3��.(;5p�=���=G8>�(> ������o�>?�?�m�>on�>Y���p �5��5�=$Z>`�N>�!>eo־1��������h��u>�Џ?:޳?*�m=���=w�=�c��Pd����l����i�<�?��!?ZrS?�ϑ?��=?�7%?b��=
�Cn���������7?�,?�o�>�[�R�ɾ}����3��?�Y?�^`����(�����Y_ӽ��>pc/�G�}�U���U|C�kzn�+������l��?�ȝ?QD���6�N�龸ۘ����j�C?W��>Q��>"n�>�A*��h��/���<>��>�Q?��>VO?�Pz?|�Z?zai>��5�z��	՘�������>��@?�ހ?(b�?�v??�>n>�
 ���پW��z�܆��ᅾg�r=�tT>8��>�*�>Ki�>�S�=�|ҽ����D6�;��=>�_>ph�>ᕠ>Pc�>{z>�=7�G?L9�>	����jn��t����@�Usu?|��?RM+?p�=�[�C�E�����a��>�M�?�ϫ?��)?t�S�]�=)�ؼ3����p�Ł�>�z�>讘>)��=��D=�>U��>���>n�7n�%�8�dR���?�;F?�v�=�̿�7~�g�:�&����MJ��ľ�ٞ���,��뫾��Y>�g7��c��\������Kx�H3�����T����1�F��>�g{<���=�PҼzDu=��>?�=Y��<��=��T����+p���u�u�`=��<_����=Tf�>�{м�}˾c�}?A2I?��+?ǴC?-�y>�*>W3����>t���=?�V>aP��x���j;������"����ؾ��׾��c��ğ�s&>8jI��>�33>BW�=)��<�f�= �r=C7�=��K���=/k�=�b�=c�=�=��>�1>�6w?O�������4Q�mZ罝�:?�8�>	|�=��ƾa@?l�>>�2������{b� .?z��?�T�?5�?Pti��d�>���⎽�p�=z����=2>M��=`�2�s��>z�J>���	K������4�?��@��??�ዿТϿ�`/>f�7>�n>��O��2���d�&Nm�=[��+"?a_2���Ծ�g�>&�=S�پ"����\=�=>�6=��-�b�]���=�w��=�R]=��>(%C>��=�t�����=��/=��>��T>8�!<��`��b�I=���=Q�b>��>�r�>�?:2?�;e?��>9�\��JӾ�8že��>���=���>~[�=�AD>ʹ>��8?u�D?-O?FD�>h�{=��>�ۧ>h�+��j�$��D���Q9�<�i�?�?�#�>�c�;v�2��b��v=�4���I�?�.?�N?H�>�P��ݿN}��h��)��½nX�O���h��e���kɵ���=A>��6>m��>I��>�	?�5�>��->��>m~>7�=�	>^�g=9��#4���>���_�	$l>��L>S\<��{x<��)�v`;��=A�<O!��>�=���>�(�>47�>a��==��>Z_����?���>�L;.�H���e��{�Z/*���>��T_>��<>o>��������?�pK>�3>�A�?}[b?c��=�ɽ?�������e�������m=�T�=�O�b�7���W�÷N�T�;��>�>q`�>��>0�D���q�ݟ�;�ھ��'����>9�Že�:>`�)>k�����������=��/=@?g`����>�a�?�%B?��s?	u�>
б�/�	��1R=�P��]<���]��ŧ
��$?
p3?�x?����"H���;��ý��>R�J�yBP�������0���1��{��
R�>X䩾9Jо��2��q��ѣ����A���n�Uw�>�qO?��?f|b��"���cO��f�:��f?��f?=}�>k�?��?\Φ����~���=�n?�w�?�t�?�|
>��=��˽C��>�R?�!�?�\�?9m?�I�w�>q<��>C����=�e$>�g=��=�w?"�
?d�
?��������� ��m�g�o]�<Ҙ=+Ȏ>�6�>M�h>��>> �="�<."O>ߋ�>���>#U[>�o�> 6x>��,��o�[?���>�%�>x�+?�7Y>YSֽ�=*�Hڡ��*2;���G�����<o�2��{!=)�t>tŀ=�c9����>��Ŀ�
�?V�>wJ4���?��޾�����?�f�>6���z"?Ew�}�P>�ț> =�>��>�v�>G�b>�ž�xi>��
���9�AjA�ϼc��&����>Z�e�n�R� ��r�[&l��������xk�c�����4��7Q<J^�?�%���T��^Ͼ�r%�)�;?�^k>=�?fu�	��=�{1=�?P��>��X��%̋��s�� ��?m?�?e�b>	k�>��~?8U8?�_D��7ĽTFZ�� ��3S/��0C�Qu��C��6ń�\��GD���|C?́x?�#?&���
Q>��?����O�����>d%-�k@E�Rw�=�-2>�9����R���:y̾)#��9>��W?�%z?ۈ�>̵��i�;�(>I:?B1?�t?}�1? �;?�x�H7%?��0>Qk?5*?�5?�9/?]?�3>��=�ϥ�@!=Lh���\����н�Q˽����F�1=Hx~=��:~R <�5=��<�<＋}޼Kv^;�(��V	�<Ӝ;=�A�=���=2�>�;J?��?��>�3�?0�R<�W���ѾÚ.?@�6>���ۅ�z���B���V>(Z?�?�F?�[>�����$���>�N�>�z>?�k>=�>N�0�	�-��̩���=)�>6D�=������L�����w=�R>�k�>Fk�>��(���={y~��ek��n3>mƽn�n���gi�!�!�����;�>�k6?��?m{=��߾�Խ-�T�^�?(�J?A�J?�L? cf=�)��V���P�)�l��;�>���=����������X���=��>�<��J��ۻz>:��Z�����q���O�����U�=|������gk���Ͼzm����=~>{�����'�����t%��\�B?�q�=i���:�j�;�����=_��>o?�>�7_��t���B�Dʥ�9�=?��>��e>�?��ྻ�;���c{�>CvE?�Y?r>�?��^�~q��N;���������0<�"?v|�>�=�>�H(>�^>�������K�+?����>'�?~����U���{���hG��H�>��"?'h>:��>
�H?E��>Qso?�nP?fT
?�kR>v]R�׾$�+?���?Gh�=U��(��f�V3r�-��>��U?0���(*�>�P!?O$?]]1?ʅp?f�?̇6>���4��`�>��y>�P�X���8|>��]?�>y�d?�t�?�x>�AM�K�����J>uc�=�!>4�l?�+#?���>-:�>'+�>+Z��t$1>��?�0�?:�?��B?ă4>;<�>禯=��?f���w��>�-?k>�>��? ��?��??+��>yA���{��W�H��	=G�r���<T�=�.=�����(����;[<�T�H�����:� =�ov��*,<{G�=�X�>�t>s'�� 1>	Pľ����E�@>�����5ي��;9��ش=Os>t�?��>K�#���=&�>!'�>ܹ�mf(?��?+�?a�$;heb�Q�ھ�J�)@�>��A?���=�m��d��T�u���e=C�m?rE^?oX�\����_b?m~^?F ��v=�,�þId���ˠO?�?5�J����>�}?��q?�(�>�]b��l�����F�b��k� �=���>6H��Dd��u�>Y7?�2�>.7d>�V�=Uܾ�.x��ќ�o�?4�?q�?N�?��>q�o�T`߿z���8'��?o^?z/�>�\���#?�=ݻ�о>H���F��㾚ાe+������H���&&������ӽB��=
�?�]s?-�p?%�_?�� ��3d���]����!
V��.��/���E��D��C��,n��������o����A= j4���;��7�?A4D?�&�Z{?/J<���	��HȾ�;�>�l��#�꽥��=��P��Y�h�j���� ��AW���?e��>���>A:?�f� !C��"�@2��*�e��=��>�j�>�)�>&z2;#	����y�ھؓ���R���>]^?k�W?��q?v!-��+�~k�H�'��Ӵ<��w���>���=Y��>saC���[��+��-���Z�L��DE��Ta
��K�=~�6?�C�>mK�>�?��?l��d2��D��:`�uq� ~�>��9?UX�>ߟ�>l���O&����>��j?�r�>���>SD���� ��Bp�����O�>�;�>�w�>�>J��#�\�'c����Wj3����=�_f?�:��|[��*�>�GJ?�=1;/�"<浓>g�c��� ����7����>ǿ?���=��5>#����r��x�4���V)?kr?�l���m*��U�>q<"?V��>/�>�q�?���>�����j;�"?B^?%�I??bB?>��>u$=׏��b�ɽ_J'�A�9=���>�\>ay=T��=�\���`�py���R=e�=�bȼ����O��;�ջ�g9d<�p =_�5>��ѿ��g����_���0�����5��*�m�A ׾ve6�1�Ѿ��v�" �ޚ��JD
=��I����y=����!�X;�?�#�?'����iӾ���V9t��l�E�>y��!6 �hJ��"�B��Ӿ3�	�nW¾���Ń��X�~�б����6?����.J��|$��/�Ⱦ�??"'R?�ӎ?)%
����w�*<�>�\v<��	>����Z���=)׿&�!�ֱk?��>���C����>�b�>6�R>�3>qK˾q���~�>	!?`�.?ٲ�>�)��bݿ�g濤\>@Z@z�@?'����9�x=%��>�1?/E>��8��%������>썞?�?�O,=TQX�����If?��<t
D�-�:7�=D;�=2�='��H�<>�k�>	_#�zFB�'�ڽ�|4>o��>�M�����N�+��<)�T>i�ؽIܱ�5Մ?+{\��f���/��T��U>��T? +�>W:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�܅�=q6���{���&V�~��=\��>c�>,������O��I��U��=ZK �
�̿{�$�Y ��_��+;��kν	�����4�Hm�퉣���6�XWܽ�>�'%>%�D>�͕>�Gp>Z"�>D�^?ͳn?�)�>N �=[?*��ד�W.Ǿ�Y=����V=!�ڴ��c-�u`���Ծ~�ݾv��03���z�߾�����L>;�8��v���/@��ru���U���,?R��>.���p�M�>�r�c6�����?7��5z�+���>S��1^�]Ԍ?�I?��W��jt���c�s�;`N?�|�<���SM�)^�>[oA>�A>'��>.�>O��H�@����k�(?��?�ݾQ�����h>�|@�H��zV/?��>/�N���>q'?�����F�7>��>�V�>��?L>�=U����0�M� ?hT?�9��!����>z���g9�/S�=���=��c���*��C+>w�?;������<H��<	�>+W?��>��)����7�������<=S�x?�?�	�>$vk?��B?c�<�v����S�����x=��W?�i?q�>E���l�Ͼ����&�5?΅e?P�N>�2h��龧�.��i�j�?M�n?�J?�b���\}��������]6?Sv?�q]��@���N�
�S� m�>���>@��>�8��.�>��>?��&�qe��Ɇ��A4���?�b@b;�?i C<;~�~c�=��?Y��>�|O�\�ž���~ѳ��L{=Lm�>�y���Nw��u�b�.�@�7?Z�?|�>�����4��R%>ẃ�ĉ�?��?!���&���Ӿ��y��H��ش�=��<�*�:�=bs�� E:�.��"3����t=��>�[@@�+��#�>�v���[�]"��5�m�J�������x��>��>QC�M^����q��dT�f+K�WkҾH��>Y5>�ŏ��)��w?z�W�:�hu꼞��>i6� ��>�P_�����Z՛��@><�Ք>��>$�>'�ǽ"��W֘?����f�̿����K-��#W?�C�?a��?7�?��k;3T��g�h�FO<H?�It?�@\?�	���l�ɵ9�T�k?�&���M?�P9
�ބ9�<��>��/?㔞>p�;�ڭ>}��=��	?-!>W #��ѿJ�����4��?Wo�?���Bؼ>�s�?ta?o�2��˳�؅�EVn��>	>x�? 8�=��ž��@���	��&2?mC?2�������_?|�a���p�O�-���ƽaʡ>��0��H\������]e�����!y���?�W�?I�?C���#��+%?��><���y8Ǿ��<�k�>�'�>1TN>�^��u>�(�:�A�	>��?�z�?Eq?��������>��}?�:�>-�?��=ۄ�>���==9��-@7��v!>8v�=|�;�?׵M?���>�l�=�{9��,/�,$F�NR����9�C�|�>ܑa?�L?usb>p���B�1�Nv ���̽�N1�y�޼i�B��@(�!ݽ5>3>>c�>� D��Ӿ��?Kp�8�ؿ�i��p'��54?-��>�?����t�]���;_?Gz�>�6��+���%���B�`��?�G�?<�?��׾�R̼�><�>�I�>2�Խ����X�����7>.�B?[��D��u�o�w�>���?	�@�ծ?fi��	?���P��Ja~���s7�C��=��7?�0��z>���>��=ov�׻��P�s����>�B�?�{�?��>�l?��o�L�B�3�1=7M�>Ĝk?�s?�Mo�u�j�B>�?������	L��f?�
@yu@^�^?�ῆk��껤������-�=rOY�U�<M}+�R<�<�x���/����>cc�>�'�>a�>6&Y>��(>H�+>�����[(����hA��:%���D��$ž�� H/��p�Ჰ���ξ��
�ش*<�W��~u�{�T�������=�U?a?R?!p?� ?-@{���>J���=t"�8h�=�ن>��2?NLL?=*?z��=�y��=�d���@D�����j,�>g�J>�~�>,�>�K�>S;x�H>�m>>:ހ>-��=�'=��g��=�yN>K[�>���>���>Dx>�3�>BT���$��`�`��J�����<�;�??�
=b�����	D
�uj���WF=&6?��>3����ƿ����[=F?Q��tP��o<��A>M Q?���?��i>�L �(�g�"ְ>�B>?ۉ�>a=6�;�c��Dؾ���>���>�$>�^�>��.��~>�
�^��0ݾ�U>n?>T>�g�F�]�v��] �F������>S�>pK�pÛ��~�cȀ���b>��]?���>(��e־�����[uj>���>C�ѻsF��X�>�&S�>Hn��V� n�=�(;;��><G?�6>><�o8��>��F�Oޢ���>��y>L�p>�"?�',?1��!�E�6���q|a�η#>[?ɜ�>�F>�#�PGv>�: ?�>�Ў�We������" ���>%W��ӣ��EV�J�F=����e�=1N�<_�	�:4�����<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾRh�>wx��Z�������u���#=U��>�8H?�V����O�d>��v
?�?�^�ߩ����ȿ6|v����>X�?���?h�m��A���@����>:��?�gY?foi>�g۾/`Z����>һ@?�R?�>�9���'���? ߶?ׯ�?��>�x?ux�?�?*Ä�(���]�䂖�ģ	=s>�^_;Ki�>����=P�ҡ��S����(�=� �g2�>��=�϶>1��־D�=��/5޾J���U!�>+]>Cl�>��><D�>A�>���>��#>�*�s���rs�u�J?��?��;<o��u<H��=Zr]�h�?"3?#[��	jо���>��Z?O�}? �Z?�;�>�"��Қ��¿�ѯ��נ<�A<>�7�>-��>��T�_SP> �پ
�M�j2�>���>�ӻ'۾}�����q�~M�>��"?���>��=y� ?\�#?��k>鮲>�JE�?��->E��x�>���>$9?��}?��?���i3�5뒿'JA[��<N>\�x?�.?�7�>Wm��w���LR�EM��Y��Mk�?F9g?�d���?m3�?�c??@aA?Spf>L�(�׾;��$R�>�T?cd���+j�~U��������>��R?�,?�u=b�ܾ���ۭ��D��l�>r�c?�()? -M��脿��9�ٕ�<���=	�8=��D<M k<%��=��Z>7J
=��N>�>��E>�H$�GtT��QL=��">�b�>��<ݒ5�S1�=P�&?6d�=.g��991=\�Q��H#��R>w��>��S���D?*�.� '��ݪ���֜�8yi�0�v?ς�?g�?M畽J�V�QP?�Ǎ?3r�>��>p�Ӿ� ��ؾ�wѽ�{��x.�e.�=�p�>�Q�<$e���C�������ً�^��������>��?�'?�x?���=���>T�Ⱦ���l���I�`���.k���!�5�U�Y3@�l<m�(����=I����̾�sN�>���ߐ�>W�>}+>9-S>���>?�:�4A>��>tK'>�t�>ބ>wƆ>M>!�
=�<ӽ�KR?������'�}�������2B?�qd?p1�>i�<������/�?���?�r�?y<v>l~h��,+��m?@;�>����p
?�Q:=���D�<U����s/��Z����>P׽x!:��M��mf�nj
?>/?K/����̾[7׽tq��?��=�r�?_-5?�*���K���W�O�^�WJ�w6F��E������v���l�^O���.���~��M����=L$?+�?-$��q����+k��,�ߟT>��>\��>{��>��@>���[.�/�P��_*��A�����>��k?k\�>��7?�&E?��>?Z�v?!��>8�=)+��p�7>\��=MF$?��?��?v?+c ?Q!?�%U?�z�>����޾Z���?��-?P�!?��>��?rC�N_k��^�-L�Y���9��=��>D���5���> ����<�� =�c?2G��o;��}󾹋>!X8?���>��>����<���pe= ��>~�>��>������l�q���"��>�#~?��
��X�<��*>zr�=L�߼������=M�޼���=m�����4�;��=��q=��
:�A�:�B	<��;���<&�>i
?�?�>�-�>��������R�Ma�=r�b>c�M>�>4�����5.���5g�x]q>N[�?��?�Ij=G��=��>�b���þg������]�<�)?��$?�HR?e֎?sw8?��"?Y >�/� ���ׄ�������?�0?���>l��6¾���i��oj?�?[wg��ͽ� ����+���t,>6����r��?"���=u\�\)۽\��?���?����<<�~��c�����pc?Џ�>W��>���>�+7��Ђ��0�̛�>_	?e�\?젾>*�O?��|?�X?2�5>�>7�'��^���1�<_�.>y�=?���?||�?j�n?Ɉ�>2��=7c%�nܾ���!A�C��­|���=WZ>�ʍ>���>�ص>>�=�tѽQYO�F}��=��{>z��>�_�>�>&�>W��;�F?��>�찾C �������:]*��Ek?ܗ?��,?S�=V���%�L例��>�W�?U��?� ?�d^����=G�D������q��h�>k?8�>��b�h��<�1>�c�>W��>y�-��F���=g?6F?1��=}x��ve����wڞ�1	���5�������ͽ(�V���=�p����q��ͫ�����ԓ¾y��B>ҾC�����o���>�W�=��>���=�=T??�67�<hId<�� ��-=��˼:-j:A���F�t�/���W���v�<;�8<@�W�P�ʾv}?.'I?vy+?�jC?oy>�x>ň6�C��>� ���:?�V>M�N�������;�n㨾yՔ�'kؾ�׾D�c�ķ��t�>UjF��>�!3>���=FĎ<�B�==�r=o��=���� +=�C�=�]�=���=���=�G>,'>�6w??��������4Q�dZ罗�:?�8�>�{�=�ƾV@?@�>>�2�������b��-?m��?�T�?3�?5ti��d�>��n⎽�p�=Q���O=2>���=��2�}��>T�J>����J��
���4�?��@��??�ዿ٢Ͽ�`/>��x>6��>#f_�L�B���I�?��-_�Ƣ?1�1�W�����>���>cJ����[���g;�=]M(>(���z���B�=Z0e�>3ݽ׃�>�+?�x�>���=i����~=�׼=* �>��v=����]b=��ܽrê���>f<�>� >�h�>��?�0?#^d?��>�%f���˾�L¾Cl�>�C�=���>\�=�oK>'F�>Z�5?�PC?�sL?�Ƴ>Vc�=���>෦>��,�Ҳk��(����*$�<�ʇ?��?�8�>� <�:��<���<��U���?w�/?g�?甛>�h�*� ���N�uU'������;,�;Z*���n�=�k�=uY,��"�=��>f|;?��?��>A�\>���>���> �i=��!�-<�<�}7�����q���7��=`�8���G�{�t���=H&l�jx<ʺȻ�����=��=�G>t�>�8�>K�e>�C�>pQL=#?����K>�-���+M�yeT>$��T^N���W�`��g�A����B>�>q>�8	=������>��#>��=K9�?�?ų>�?̽i���^���cx�o����J�<e6�>�5���-8��gO�U�Y�����A~�>%��>�?��>��3��]�n�4=V����"��$q?�#���7��s��}����Ž�7���	�G�,�k>��v?����'>8q?�?|��?��>�h%�a�����=S���l�T�ݣC�W̘���D�/�?��>o0�>��1�&`�)?̾�	����>�I�|�O�
���ޥ0�N���Ʒ�b��>,	����оD3�Xf�������B�"Lr���>��O?�?VBb�HT��`PO��������s?<vg?T�>�H?�=?$ס�%j�rv��l��=��n?��?>:�?{>dd>e���%�?�f?�֛?uA�?�P?<B�Y��>I��=v�>o�u��Cn>l�i>U���%�m=%5#?��?�?���;R����ԲҾrF��'��V�	>Q>�>=>z�>S�='5P>�\�=���=�E}>�:�>�<�>>��>y��><�x�2���H?[��>�f�>ֿ)?���>J�Ž3*����!>��k�� ���WM�ա#�l���(���Qq<z��=�X�=v]�>)~ſ[z�?ͪ�>�f-��,?-�������MGs>��W>��ͽ�u?���>q�>��>���>���=��>�L4>�GӾ�z>���Mi!��1C�τR���ѾЇz>B���-&���3����HI��p���d�9j��/���==��p�<|E�?l|��t�k�w�)�����}�?�Z�>�6?
Ԍ�Rሽ��>��>\ˍ>�R��2����č�&^���?^��?�Hc>$�>A�W?:�?�Z1���2�gZ�.�u��A�P�d��`��鍿렁��
��S��>�_?u�x?�|A?g��<$*z>��?��%���>r/�'%;�7�<=PG�>����`a�>�ӾH�þ7G�IF>E�o?��?s;?VV���=�>rTD?�K?��?�qk?dC#?�wE�x�>q��=�?-�>uS?Rd?}: ?�x2>��2>,�M=�l'=_��.휾b��������X�=WC�=$5�d��=���=b�k�@�����<��+>�)�������ⅼ�p=a��=��>e|Y?6��>>��P?����
��������S?Leg>�꫽���U�z��k���wD>`؉?��?�C?B�C>=�V��>D���>8�>W?>e�>�f�>�b����ݾ3dY=o.�>´�>A�>T�:=jo[��]�Y�a�̋Q=ޡd>Q��>�}>�'��d9&>$����uz�8�d>��P�|����T��G�w1�$mv����>��K?}�?`��=V�� !��c�e�O)?��;?�IM?��?��=H�۾@:���J��L�\��>f��<			�߯��#!����:���;��t>�ߞ�d7���o>����ﾁ}o�m�R����4ݫ=+�pq	<W��wQؾ�c��Oǰ=��>� ƾs%�L����j���I?��=�����h�縱��>�j�>���>5���ZIX��;<��°����="��>f8>�������F�{L�] �>ĽE?��^?�Ń?�����r��uB�A���,K����v�?���>�5?�B>���=SO��T���?e�JhG���>��>3���eG��螾AY��1$��\�>�?.>K�?נR?K?��`?i�)?�0?,y�>ﶽ=����#!?<��?�<j��7l��8�\P2�#�?�d4?�����_�>�7	?z-?�)?�SS?\??��=jY�ڱK���>��l>�>Z��ť�S�Z>(C?���>(O?J9|?_!>�#�2��ܒ��3>�dC>��3?�Y?;�?��>}��>y�����=֠�>�c?1�?F�o?�s�=;�?}B2>L��>��=v��>���>h?
XO?��s?g�J?���>Sύ<�$���9��<5s�<�P�st�;��H<�y=����t��Z��C�<�;�m��>�����D�搼��;�^�>�Tu>u�����.>����ˀ�c��>���=gᦾ�׊�<h'�I�=�� >M��>��>��$�n��Z�>��>f���5?�E?T�>C�J�lKg�#ʾ�i"�ew�>��'?�R=��s�������Y�z�>�ւ?�^U?Y����
��<a?�%U?p�p3�+����J��;��P-V?�e�>�J����>�w?��Y?�v�>�+��Rg�x���#;W�ޔj����=ͳ>s��i�i�_��>��'?���>Up>W�>xy�I�q�����?�u�?\��?b;�?�'>�.r���1�����-�q?��?l����(?�������h]�}�I������Ϧ�y���Uʘ����'�0T�n:ѽ���=�?/�v??�j?�N?��پ��^��t\�Rt���^������"���T�a�>��?D�˔j���b��8��þ<ZJ�}dA�>s�?��Y?�yN���?y6��i�&���b�Y)�>$���%:Y�q03���j���?=`,"=��l���
��Ւ�X�?^��>�o�>��.?�[g�@��m*!��@��_�fЖ>�N=��>u��>;�ͽ�G�.)�B� ��t��$��b:v>Oyc?�K?�n?�q��,1�慂�r�!�K�/�5f����B>�r>���>�W�����8&��V>���r�����u����	�i�~=2�2?&�>ǲ�>�N�?^?�y	��i���bx�m�1���<y0�>)i?�?�>a�>rн�� �i��>Jqk?{��>;�>���}���s���5½�>!Xo>�e?�T�>�Cǽ��T��ߗ�"����g&���6>Ref?̮]�A���<�>>�oU?t导Q��]�>��{�l`��,׾9&�}�">�	(?�7=��=KѾ�����P����a�%?�z'?Q�����(��υ>9�
?�b?���>o��?Z۽=�}���z�]<�>>�m?k�Q?%?I?p̂>�ڍ��=��tT׽%$���qa=Qm'>�\>�� �>��</<�����d�=x/�=�Լ��<�2�����[�=�>>�p>~п��I�B���@A�^I��u��om���15=DX������%B�(P�}��������������6"��"�(5=�"�?��?_������(��
����ؾ)]?���q�����Y$#�@Ϯ���r!r��H�3T���$y��fI�ی'?ȵ��۰ǿ����. ܾj ?�  ?p�y?����"�b~8�0� >�C�<O���_��*�����οS���^?F��>�������"�>�݂>�7Y>��q>$I��y���l��<��?�f-?��>s�q���ɿ�p���_�<s��?5�@��A?��)������΄=�.�>�S
?TDI>۪)�*6"��͞��>�a�?���?��c=.)X�Tr���X?�^�<O9�U��+�=u�R=4Dc<p��5�7>��>J�佸�E�8��4�S>��>2Bg�/� @"�[�<��3>����sؽ�Ԅ?�x\�lf�c�/�8T��NR>��T?y.�>�7�=��,?�6H��|Ͽt�\�D)a?�0�?��?(�(?Aܿ�6՚>��ܾ��M?�E6?��>�d&�q�t��w�=gE�{B����㾤&V���=��>�>R�,�ψ��O�������=6���H(Ŀ��Q�������C-�s�E�j�K��
���3Z���������XW�=C6s>��>�V�></>�%O?ya?�Ͳ>?��=ˌ���å��Ⱦ�_%>��Y��Kz�������Ľ��f�4�e�׾���Z-��,�抢��g4�R��=��L�����?*��z���K�Zf@?��=Tp���9���h��g���Ծ��= :'��*�Ov+���_�eU�?fqY?�-��bm�b�!Ľ�	��=?S{*���	�A)�����;7*�����=�/�>��=�� ���B��YS�P0?��"?���Z3s�L�K>.�>�3=$�,?�+?��R�_��>\�,?r�����ܽ��=��=D@�>F(�>��#>Y�����׽�+#?w�X?��2����[�o>������/�=���=4���7<$�='5<1���>=�\�ñ�;CmU?w��>9�"�zv�e9q�/�G��E<��o?��?��>l�m?�D?˕J=EK����\��L�1�j= IX?�Fj?%�>=��H�۾�����-?�\?Oq>�1W�#"��^*�Dz���?Scv?�Q?_-ͼ<�y�z쎿[�����:?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?s�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������{��=����?>��?����F�<O��o�q��-��n/=9�U=s�F��N�V)ﾺm5�!ƾ0��T����(��0��>P�@}-���>�u� ࿇ο�!���۾�w�Q|?�ӕ>�	սP.��ǐi�Ԓs�G��I�����ޣ>~�>�욽��a0{�E�:��ˏ����>A��ω>$�T��)��T���`�=<��>���>'9�>�:��%U��Z�?	)���ο���� r���W?�-�?��??�?U�<�xs�c�x�*o6��F?v*t?�Y?�90��_�fF�$�g?DH���P��T��4��y>�W-?Q�>�L&��õ=]�>V�?��r>�#��f¿垳�^L쾝�?�;�?с߾��>}l�?}y:?�$�'��������0�����L?�J>s���#��-7�F�t��?�3?��E�]�_?(�a�M�p���-���ƽ�ۡ>��0��e\��M�����Xe����@y����?M^�?i�?ֵ�� #�d6%?�>b����8Ǿ��<���>�(�>*N>DH_���u>����:�
i	>���?�~�?Pj?���������U>�}?v�>�ބ?��=�3�>�y�=�d���"��:%>4=�=�&D�V'?܁N?v��>SO�=��=��T/�=FE�ʧP���"2C�[��>�b?&M?��Z>|�Ľ�_3�|� �ѽK,�8W�7>����I�i�7>��?>��>S2F���Ӿ��?Px��ؿ�T���'��A4?��>�?����	t�Ѽ�t,_?[��>����(��21��,�����?�H�?��?�׾�;˼c?>��>�]�>�AԽ��N���Hx8>�uB?���3��q{o��ֆ>���?m�@�ɮ?��h��	?���P��Va~�,���7���=��7?�0�F�z>���>��=�nv�ڻ��?�s����>�B�?�{�?��>�l?��o�B�B���1=RM�>؜k?�s?�Mo�^�ӱB>o�?)�������K��f?��
@vu@x�^?&�տ����j喾���_��s:�=�e�>E~�.b���
\>e?�
���ks�>ļ�>��o>�A�>ρ�>��->*�=�ރ�%|#�E��-���.����{�۾r�]��)3������4.�G4���ޭ��y����q��=T�3�3�ý�C>��=�FV?�P?��m?��>h��>�(��,=�s)�3ņ=H�>|�1?aIL?Ԧ*?U��=D����Te�I}���	��3����>D�G>��>)��>�M�>��;6�N> ;> :�>j]>6�6=z�j;�=#�N>(��>���>KƷ>ep>>��&>c���b����g�����k���Aע?{#��^eM��;���I���!��@�=Ԏ/?��	>4e��BWϿ����LG?�������!,�B	>�0?=fX?�>���O�!�>\�/hm��G>�[��}b\���)���J>iV?�'y>I;�>ɪ(�y<���>��Iվ���>=�J?�	w��H��^�e���R�h���%>��>v=�=[�.��ԓ�;D~�񿜾�?a>/M?���>����¾�׾�ｾ� �>{�=3�=�q�=ݮ�>�W�=Cwd���	�R�>�qh�E��=#
?�v.>0�=a8�>����Y�Y����>�	H>n�)>�+=?ir%?���#�~�"�����6��Qj>dL�>���>Ϧ>BJ�㚴=M��>��i>B@��>���X��_=��WR>T\���^��Bg����=�g��yh>��=����<A���<�~?k��䈿�뾌^��JmD?�+?���=�HF<��"� ���G����?K�@�k�?��	��V�i�?WA�?�	��K��=�|�>�׫>�ξu�L�k�?ƽ�Ƣ��	�+,#�R�?�?�/�"ʋ�!l��8>�^%?կӾ"w�>kh&��y��N�h��0P��=>$+-> rD?�b	� %D�h���U ?��?����ě�J\ѿ��z�F�?S/�?c��?#���������x�	?̰�?Yܐ?�D>�n&�r��;�<>t�?�96?"E?)���M����>A-�?��?�#N>@�?�q?���>^ �2.�����ފ�/��=����ߘ>��>m����E�K6���Ĉ�
g�� �ni>�G0=�կ>b���b���s(�=���� ���r�3�>�l>��D>U��>"�?C>�>�<�>UE�<t܋�l��-��JDF?yA�?E���h����<C��=D����	?{�@?R���$Ĩ���>>NE?��~?��[?ȯ�>������������o��<&�->i�>e��>*����i>������K�A>�w�>JV>�@��i�A��v�B@�>�D?uf�>�Ǜ=B� ?��#?��i>+1�>�v=�T���p�F�ぽ>���>{-?�?��?a@���_2���������=X�4^Z>��y?�?R��>9����ҙ�f�����Q�t�E�!]�?�Ic?��佀?�w�?�C?�@?�Tb>8��!վ���o��>��?���>���oY�ou���?�z+?���>�~�>f}2�2A�=�I)�����?Ǟ}?�2l?�~�ʼ��~%A�M�=HW���r�<��$���7=]��>`=Z�����&=�E�>��>AF�0+2���r=}�=�P�>Ѫ�=A�Nh�;�<,?�G�SӃ���=��r��uD���>3;L>������^?5v=�?�{�0��@x���U�
 �?|��?zj�?�	���h��%=?��?S?&�>vK��	޾7��ZYw�#~x��x�n�>���>�l��ŏ�������F���ƽ�g��C�>9�>}�?� ?�2V>��>7X��!�(��������]���"�5���.����c����O�Hʻ�����Zt�FT�>�؝�ث�>��?d0i>���>��>e/���>PiZ>S�r>K�>�ri>�6>�=�=���9{�D�P?�ݾ4�K��J�����>?�b?���>�䜾U�7�����?/�I?[|?��>J`n�;�@��	?3v?2lm��?���{%���];�9���:�U> 4=�5=��=d�����H�Ѷ��U?�^'?ܑ;�G>���¾8}����o=�H�? �(?j�)���Q�b�o�ʪW��S��;��g�_����$��p��돿�[��� ���(��h*=Q�*?��?ƃ�n�&���k��?��f>���>�,�>Ӿ>��I>ѽ	���1�5^�T'������`�>�b{?=i�>�BI?
I<?H�P?�CM?Z�>4y�>���Y^�>+�<t��>���>m9?��-?o90?8�?�+?Vc>k������ kؾ�?�?�	?K?.�?����p����^��h�h��x�F���Ɂ=�P�<iVؽ�2s��V=��S>��'?l?��'�BJ�kw�>2�*?���>��N>'7ž�b�=��ͽ��>4�.?���>R^�/���� ���??�`�?� ���O���=��>RF�������>gk<�P7=2��=h�
��^3��.(;5p�=���=G8>�(> ������o�>?�?�m�>on�>Y���p �5��5�=$Z>`�N>�!>eo־1��������h��u>�Џ?:޳?*�m=���=w�=�c��Pd����l����i�<�?��!?ZrS?�ϑ?��=?�7%?b��=
�Cn���������7?�,?�o�>�[�R�ɾ}����3��?�Y?�^`����(�����Y_ӽ��>pc/�G�}�U���U|C�kzn�+������l��?�ȝ?QD���6�N�龸ۘ����j�C?W��>Q��>"n�>�A*��h��/���<>��>�Q?��>VO?�Pz?|�Z?zai>��5�z��	՘�������>��@?�ހ?(b�?�v??�>n>�
 ���پW��z�܆��ᅾg�r=�tT>8��>�*�>Ki�>�S�=�|ҽ����D6�;��=>�_>ph�>ᕠ>Pc�>{z>�=7�G?L9�>	����jn��t����@�Usu?|��?RM+?p�=�[�C�E�����a��>�M�?�ϫ?��)?t�S�]�=)�ؼ3����p�Ł�>�z�>讘>)��=��D=�>U��>���>n�7n�%�8�dR���?�;F?�v�=�̿�7~�g�:�&����MJ��ľ�ٞ���,��뫾��Y>�g7��c��\������Kx�H3�����T����1�F��>�g{<���=�PҼzDu=��>?�=Y��<��=��T����+p���u�u�`=��<_����=Tf�>�{м�}˾c�}?A2I?��+?ǴC?-�y>�*>W3����>t���=?�V>aP��x���j;������"����ؾ��׾��c��ğ�s&>8jI��>�33>BW�=)��<�f�= �r=C7�=��K���=/k�=�b�=c�=�=��>�1>�6w?O�������4Q�mZ罝�:?�8�>	|�=��ƾa@?l�>>�2������{b� .?z��?�T�?5�?Pti��d�>���⎽�p�=z����=2>M��=`�2�s��>z�J>���	K������4�?��@��??�ዿТϿ�`/>f�7>�n>��O��2���d�&Nm�=[��+"?a_2���Ծ�g�>&�=S�پ"����\=�=>�6=��-�b�]���=�w��=�R]=��>(%C>��=�t�����=��/=��>��T>8�!<��`��b�I=���=Q�b>��>�r�>�?:2?�;e?��>9�\��JӾ�8že��>���=���>~[�=�AD>ʹ>��8?u�D?-O?FD�>h�{=��>�ۧ>h�+��j�$��D���Q9�<�i�?�?�#�>�c�;v�2��b��v=�4���I�?�.?�N?H�>�P��ݿN}��h��)��½nX�O���h��e���kɵ���=A>��6>m��>I��>�	?�5�>��->��>m~>7�=�	>^�g=9��#4���>���_�	$l>��L>S\<��{x<��)�v`;��=A�<O!��>�=���>�(�>47�>a��==��>Z_����?���>�L;.�H���e��{�Z/*���>��T_>��<>o>��������?�pK>�3>�A�?}[b?c��=�ɽ?�������e�������m=�T�=�O�b�7���W�÷N�T�;��>�>q`�>��>0�D���q�ݟ�;�ھ��'����>9�Že�:>`�)>k�����������=��/=@?g`����>�a�?�%B?��s?	u�>
б�/�	��1R=�P��]<���]��ŧ
��$?
p3?�x?����"H���;��ý��>R�J�yBP�������0���1��{��
R�>X䩾9Jо��2��q��ѣ����A���n�Uw�>�qO?��?f|b��"���cO��f�:��f?��f?=}�>k�?��?\Φ����~���=�n?�w�?�t�?�|
>��=��˽C��>�R?�!�?�\�?9m?�I�w�>q<��>C����=�e$>�g=��=�w?"�
?d�
?��������� ��m�g�o]�<Ҙ=+Ȏ>�6�>M�h>��>> �="�<."O>ߋ�>���>#U[>�o�> 6x>��,��o�[?���>�%�>x�+?�7Y>YSֽ�=*�Hڡ��*2;���G�����<o�2��{!=)�t>tŀ=�c9����>��Ŀ�
�?V�>wJ4���?��޾�����?�f�>6���z"?Ew�}�P>�ț> =�>��>�v�>G�b>�ž�xi>��
���9�AjA�ϼc��&����>Z�e�n�R� ��r�[&l��������xk�c�����4��7Q<J^�?�%���T��^Ͼ�r%�)�;?�^k>=�?fu�	��=�{1=�?P��>��X��%̋��s�� ��?m?�?e�b>	k�>��~?8U8?�_D��7ĽTFZ�� ��3S/��0C�Qu��C��6ń�\��GD���|C?́x?�#?&���
Q>��?����O�����>d%-�k@E�Rw�=�-2>�9����R���:y̾)#��9>��W?�%z?ۈ�>̵��i�;�(>I:?B1?�t?}�1? �;?�x�H7%?��0>Qk?5*?�5?�9/?]?�3>��=�ϥ�@!=Lh���\����н�Q˽����F�1=Hx~=��:~R <�5=��<�<＋}޼Kv^;�(��V	�<Ӝ;=�A�=���=2�>�;J?��?��>�3�?0�R<�W���ѾÚ.?@�6>���ۅ�z���B���V>(Z?�?�F?�[>�����$���>�N�>�z>?�k>=�>N�0�	�-��̩���=)�>6D�=������L�����w=�R>�k�>Fk�>��(���={y~��ek��n3>mƽn�n���gi�!�!�����;�>�k6?��?m{=��߾�Խ-�T�^�?(�J?A�J?�L? cf=�)��V���P�)�l��;�>���=����������X���=��>�<��ZH����>���u澮�H�������>a��2o��}$�JH��&��I=�<�@�aX ��[-��B���K���N?�zл,߾7v�����#c>wE+?�H�>��?���<vA�Փ�N�}<��G?�Q>�>b��E�3��#5���>�uD?f�\?��?��Is��J��z(��h��5a��G8?��?!�?�;�>{,1=�.B�ţ �	�n�|o=�I��>t??��$�PM�k�V����cC�t�>�|?{X�?�%^?��%?�u%?ڙ?j�?R�2><�e��ڡ��K!? ˄?zY�=��,�&KL�*�-��F_��>�(?����׷>>�G?��F?$U?q)>?+�3?�3�=!���27���|>s\>�oW�%���Cǚ>9^S?4�>�&O?&��?|�;>��N�G������K=&�*>�*?(3 ?��?�K�>��>o����Έ=�@�>*�c?ԏ�?}4p?:V�=��?��5>���>/s�=�>K|�>S�?�N?߹r?6�I?���>��<�|��,���x�������9�J<��b=H���W��.��[�<�<5�������4𼉢;�E�C$�;g�>X*t>;��c�0>m�ľ�F��ϯ@>&���<&��0���bi:��y�=]q�>�?��>%�#�i�=��>T�>����(?��?B?�^;5�b�q�ھ��K�F�>�B?�j�=��l�x}����u�c�f=��m?Ő^?��V��	����a?�F^?a��6�<�(þ01X�����cO?��?�pI��i�>z?��q?f��>ki��#n�������a��,r���=���>i���a��ۘ>��6?H��>��_>�$�=N�پ&w����1�
?&8�?8W�?�ߊ?��*>�m� �߿��׾���O�g?��?g����&?Q�9��ʾ+F��^�6P¾ ۤ��P����[�*�����ԽBe�g���g)>�$?[Wm?��^?��l?uI(�n�d��X�1Ս��Gs����zW���V�"+�#�>�܆��Q������侪_Z<��F��aQ��Բ?�??Jk���?jJ��Kվ�3��ͮT>{�q���e�I�F=�ݹ=���=Mh=��+�$�)�o����?-��>n��>��=?�h���G�<2�\�e�&��L@>3�>%;>��>�dR�{���#ڼ$w���������U�>�]?�mU?[ y?cz�;+��~�N�0�������kۇ>�]9>��a>0 ,�M�	�)c�`�2��p��s�>�����G�
=?�(?`�x>�|�>�?��?�쾠2��ݠv���)�w�\=U��>�kp?�3�>��z>��޽�X���>)�k?���>~�>�Ym��.��o���*���+�>@�F>��>�w>'HH�
{�A���ٍ�p�?�&ȳ=Lnl?J���O��Ѧ>�i??$���$�����>Êڽ�)�JF
�$#��Y��8�>=��=P;>�7̾}-��X��/����m(?�f?���b%*��}>�.&?K��>�΢>"Ԃ?��>�`ž�gW��T?8[?�`H?^y;?�[�>d��<&���9}˽���;=!�>�^Z>��.=���=!�� O����V7�=�=|� ��츽�����Y �,�Z<�k'=�V=>]�Կ��I�������E��O���������ŷ��#��3jپ�q侤I���V �.���q����o�������i�?��?�3@��'[�š��*���[����>}L��� 4�#�_��}��3�)�ˍ���Ⱦ�F �|__�8&Y�"�y��$'?�䉾�ƿ�Ġ���ھ��?8�?רw?��	��]#��6��>�6�<p��������G�Ϳ"����^?��>y��SQ���K�>��{>.?>�.p>qӇ��[��)��<N�?H�,?���>v1p�[(ɿE%����<�_�?Wh@>xA?��(����R/V=���>b�	?ޫ?>�Q1�o7�#���K�>D:�?���?�6M=O�W���*qe?-� <u�F��v߻���=(�=�=�i���J>���>�H��:A�e۽UC4>ʤ�>�\$�·��x^���<r�]>�>ս�-��/Մ?{\�~f�w�/��T���U>��T?�*�>�9�=��,?B7H�_}Ͽ �\��*a?�0�?��?��(?bۿ��ؚ>}�ܾ��M?jD6?���>�d&���t���=�2�nu�����'V����=���>e�>�,���_�O��H�� ��=w��K-ǿ����;�Ÿ��qnD<���;������C��0=��~�Ⱦ#,5�Z�<Q�=A>�z>>�&�>,�\?#8q?�V�>%�p>��=��?Y���ھ�*/��R��#+�<�Y��л��׶��T�n�ྦྷx���v�� �a�ξu=��;�=�R��_� ��~b���F���.?n�#><˾K�M��Z<��ɾ�������{p̾�1�f
n��ş?q�A?�ᅿ�V���=�Zv��a�W?��3�������=�
��X�=�ǜ>D��=��n3���S�%�/?M�?N����8����)>-��f��<��*?W�?<�"<�f�>=#?V*����QZ>�m+>�ՠ>Aw�>$)
>Mԭ��۽k[?v@S?�f�<�����>����X�s�6�T=z>��-��!�1&Z>�3<'����L��|���<��R?�1>>�{S����)��G�m�'1'���?4f�>0��>Ȁ?˷-?==�w-�x�b����7A<�nx?�}?��<f;>�'��wZ����k?c�`?��:���b^�.��#�%��!?U5?U�"?�^=)�z�g ����*��SV?w?�+I�R��������p��� l?��2?Ƕ���?��`?����������R��פ?� @+�?�s5:����r�<���>���>�;��Ѳ�A#�x�Z���=DM�>�/�C��|.�P.����>��?
�?~Ɂ�p�⾕�9>M���i_�?�E�?������ֈ�]p��!q=>��.=�2�<f�u]*��ȾQ;�꺾>R=��e>��@X"M�
�>��q��>ٿ��ÿ�X���f�������?���>Al����ھ�Jx��c�\�'�61M������`�>+�>膕�����>�{�9�:�(��M�>>	�#��>��T�
����➾!�8<Mf�>t��>��>��ld��(��?�[�� )οn\����d�X?��?9E�??G4<nqw�Ph|�f�$�5�G?(�s?�!Z?k/$�m]�K'?���j?�����m�S�1��yJ��:1>��/?P��>n<6�8N�=�}|>��>�:+>�$=�] ĿUԮ���꾢��?�9�?���5;�>w7�?��)?�C�CV���0���1�<�8?��Q>ꕡ����K��w��z?s6?H?�,[ �L�_?�a�7�p�_�-�"�ƽܡ>�0�f\�BQ����sXe����@y����?*^�??�?N��� #�(6%?��>����08Ǿ���<ɀ�>�(�>)N>ND_�ųu>��&�:��h	>���?�~�?j?��������V>
�}?��>��?�^�=M��>��=1���gF��s#>�F�=ED@�5g?�iM?��> e�=�9�x,/��XF��R���y�C�=�>&�a?�L?�Vb>Jj���3��!�P�ͽ�3�s+伅v?�{a2�O��^�4>5�<>6�>�gE�K�Ҿ!�+?aF�R�ۿ�-��W����?A�]>�?�W&�{�-�>&>�?��>g%�����L����`e����?�s�?��?.�Ǿ�:�5	�>�n$>H٠:���=���=�]p�ۘ�>W+v?�e���l�JIs�Eɣ>w��?`�@���?�҅���?ӈǾ�/l�d���rt�-�z>�-?(�����>�-?��=YVf�����v-t�:�>&j�?W��?�i�>��T?��i�����E�=�u9>\�6?[x?�T$>���z�>ik?�@Ҿ�����g	�9MB?6{@$@�)J?� ��mn�i���Ѿr�ﾎ��<~Oq=�4.>��7���}��9x=,�����#m�=>;�>��X>��l>��>3*M>�1<>����@$��䰿�9��B����[)��0;������O���$������߾ɼ��˥�����ϔ��|>
�O?��U?mmq?�?��j;`8+>g��*��=��+��/=밒>~1?tKQ?�3?!�=hΏ���^��6{�*I���ꅾa��>�
2>�A�>��>���>��=�J=>$nB>{?`>[�
>,�F=�VX=��=��>NT�>��>���>i)B>�h$>*�������Sg��ia��7��A��?�.��Z7J������#�����ӽ�=�+?���=0j���ο������F?�������k�ݞ�=Ƅ,?+�^?]>➴�Jo��o>[y�FY}��<>p�ս|�Y���&��BI>Q{?՚>�v�>~�%�b����8��E=[Ej>���>]3оD�o�rpb�_|���q�1>]v�>wV���%�����h����Y�F�	>yD?�L>Vw=�Պ�z��H�>��~�>D�=�g��:>�@�>oͽnn��H��t�=�l"><�>�I?*: >�=Y��>N>���Oc�b,�>��t>>�LB?�T+?��"�+a��Ĭ���5:�_�>Lm�><��>��	>�N��(�=5�>�D]>f�%�Ä��W��3�4��~>�h��e�,�H���S=3i��K(�=\=K��e	@�?�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ|`�>��~��� U���r�ch�=��=[�<?�i�m�����W���>�?����F����տXƌ��$�>���?�?��`��"����,���	?�d�?1�^?"�>��뾺^��_ɂ>��"?��a?��>��[�!�S�!?&��?⦑?6,>m��?��X?�/�>��f�=��/|��Z��}_C=�P;��V�>���=9yþ�X��ꀿ�c��BW�^J�� d>�)$=��>X�R=4Й��§<��<=����4<�R�>�ܝ>�'�>�O�=��?ݣ?�I�>���=KG����b�N#��J?ڟ�?��l�k�q��<f��=4�X�?HG0?�oռ�վl4�>g�Z?�#~?�X?tՌ>T���G�� k�������<�uG>Y�>�"�>E=���-X>Rl־J�?���>���>:]`�E�ྣ0y�^�Ȼ��>��?KL�>t6�=߯?�n)?t�M>%ȟ>�?�����gG��}�>���>�n�>��x?�	?�x���E-�z�o�IvX��SN>e�z?�X?��}>z���5���(���U�|�u?�qd?.ꬽ��?�r�?MC1?b�9?�� >����!��v)=I�>��?���kVE�Eɩ��>����&?b�!?���=���e��lش=�U��"���(�>��N?xj	?{�Ho��rU�%��;��<�7�-~�=5����J'>Ц��)���J�1=�>~eC>�%����u��p���c&>��f>/WI=�� �t#�=�&)?V��=C��;v8���6��Ov�͌�>.S�>8WH���?�5��~R��8ʿ�Wn��ǘ�q��?�F�?⩗?b�ý�Ah��6?Ǖ}?��>(�>�L���`���P����i�a����?�=/�=xW�P->�ՠ�����dw�Vu�<f+�
� ?B*�>o�?W(�>8j>��>\5��yS#������M�P_����!8�>�(����S���4����3n���g��k�>ͭ���>b?��V>)�|>�U�>mjA��ψ>ݝN>�;�>"��>MB>s�>P$>
?�<�>����Q?�;��N%(�|�羶L����B?Fe?�L�>��|�pK�������?��?��?it>+=g�J|+��?\��>�|��P?��=@Z���<󽸾:T��s��px(�΋>��ϽwZ:���N���[��?�?z���̾����5���t)=Αw?�O?��2�	U��^y�:@6��Y�eoս���F��X��u^��'��^
��������)���]�f�8?gp�?(��r��	���:s�Q�?�2�a>Ϧ�>MJm>^��>�D�>����Vm7���l�lC/�%���?��z?�0�>��F?T�1?�=E?���?~\�>L�>����TQ$?�H��E���?JE?�{7?��7?�?�?��Z������������9�>?Ņ?�� ?G�?4�)?�<�-���>��ټ��M½ӈ�>���>����'�h~�>�#=P	?�6ɽP�2��X��i�h>w�=?0S�>3�>v�����ڔw<��>#	?�'�>����_9r�U��_�>ǖ~?�1�x�"=ȳ">��=���K���=%����'�=�/��4��S�+=h�f=	=�=������V�;Q
�<�	C=��>�P ? �>Ӈ>î��|$��
�Uc�=̙a>��[>X�>�׾��V�d���{>W<�?Iճ?�ic=��=,�=�<����������;����	=k�?�&?�
S?|W�?p)??M�#?jw>���!f��dG���@��S?�,?+��>>��إʾ�쨿�|3���?=F?TCa�w���6)�Ż¾*4սq�>�M/��~�"��pD�L'�����e���F��?���?~A�^�6���1����V��;�C?4>�>�l�>j�>`�)���g�G��5;>�|�>�R?1t�>�!I?��?�zu?�=>�R%��񢿫������=@�x��e^?���?]q?�8]?=ٸ>��>����1Ծ����aN�_��ME���s>�E�>��>4?��>��)��p[�3Q��B>��>q-?��>�O�>�0>>��<��G?=I�>Ӫ���s��TO��!p<��s?�F�?�4?70=�����Y�MI��t��>M7�?u۳?��5?1�^�/	�=��P��D�_��>�޺>��>�O=�ߖ=��0>���>�>���:6����"Y?1X=?��=Qƿ�Rr�Ӣq�㚾���;���]b�������]�g�=���_��ݧ��[��ߝ��(���:���М���v�v��>��=��=�"�=t�<�Ю��P�<HY=9	�<��:=�?��5Ʉ;x�M���j�4㛽�b��I<��H=$�%�O*ʾ��}?O�H?��*?&DC?�5~>��>�z4����>�ڄ��k?x�R>D�K�G!���H:�&������
-پ��־��c�f����>�7O�!�>�@/>���=�'�<H�=�p=��=�G:%�
=���={�=���=���=3�>�p>�6w?;���㲝��4Q��Z�H�:?�8�>,|�=f�ƾ�@?��>>�2��×��^b��-?���?U�?k�?0ti�Pd�>���Ꮍ�q�=6����=2>���=��2���>E�J>����J������g4�?��@T�??�ዿ��Ͽ�a/>TC>��>3PQ�y)���g���=�98H��|?��=��ƾAٍ>]�q=��޾
pžT�=�J:>4�</2�c_��.�=V^�Y#=�	u=�v�>�_M>�~=#���;�=�,=���=t�_>�#�אu����6G7=䥹=��\>Z1=>��>�+?=0?�c?���>�l�
wϾ� ���>(��=얱>�φ=��A>x��>��7?��C?�J?bذ>s��=���>Ģ�>��,�0m�p0�W	���!�<ꖈ?�φ?���>�o><��@�e�j_=�*Ľy�?j�0?'�?�%�>^��qAƿ�,7�G��u���Ud�6�Q�<̾���b���x���S>�3�>4� ?8��>�D~>!c�=B�(>���>���=�>>f�> �k�k�<�zk<���=�� d�=�
y��0z����;���6�\�x���8���$z:����=���=)A�>}�>,x�>:��=,��� )>[��c�H���=!���-�;���`�t����.�Y�:��B3>�b>����������?��n>"8>l��?��u?��>Y#�bҾ����es���C�o��=��=nF-���:�!a�S�P�̾V��>�/�>L��=�%�=Hl���+ ����圂�t|�`2�>��`���=��v���J��픿:n�:tU=1�u?����M2>ĳ�?�{?�!�?O�>��4�������<�_ �����5)�U̢�tO��5�?{��>��>"6��vF������[N<ղ�>(�`��VA�����91+���3.O���>H u��(Ͼ�+���p�M狿�vO�mt�٪�>ud\?)�?�!����d��*0�}�	�#����]??�J?iӈ>F &?d?�����پ+)f� ��$wt?��?A��?Z�=�w�=,Ӫ� ��>��?�5�?X��?�Hr?yT=����>l�q;��>�D��_��=��>#գ=���=�%?e�?��	?]���W[	����Lu���^��P�<'m�=Qn�>J�>@�q>u��=��r=�i�=��Z>��>3�>�Dd>U�>ː�>�4��������:?�`>���>f�?���>#CD>d�>��>�O0=4�}<��{���\�ʪ=~=�m�m=f>SB�=l��>۞�:�?c�?�U&��M?������= Y:=ǖ��n�>tH�>�F�>�:l>�}�>)E�=xr	>6��>�ҷ���R>ݾ>k�y�N�z�E���Spx>����^����o@��T���־�����E����*�;5r=�$�?f���\���WC�B%�ۡ�>���>1�?�� �<:N�``>���>��<>���;p������2�ZØ?���?2=c>��>��W?ܙ?�1�3��uZ�ѭu��&A��e�#�`�O፿r���r�
������_?��x?]wA?�_�<�9z>���?��%�Yӏ�5(�>�/�j&;�C<=U-�>D*����`�h�ӾJ�þ�6�BF>S�o?�$�?�Z?�LV��c=��3>Yn?��M?��?u�s?N:l?'�E���B?��>�bk>�R?UR?���? {q?ҏa=�A�=�a�)a��ڽK����}3��.� � �10S=�o>�9����h2>��@�VR{=eGϼ�X=#W�,찼�+�=@_=�8>�s�>�Fp?(H	?��j>I5?ԛ�χ��x�"�MY?�N>�Q2�}B����ޙ��j�e>F�U?*��?ҟ]?��X>�Eh�9]�@<#>�1�>�A�>um�>���>�N
���=�?�<�#>�%�>a��>�%�=�X?�������,�=FN>���>׶|>�Q��V�'>wm��m�w��d>��Q������T�տG��2�v���>��K?5�?"��=��������e�7 )?�P<?O�L?E�?=ߒ=_�۾��9��7J��i�x��>6Ӯ<��'��������:�X�:�	t>�d����þG6�=�6
�_ڃ���V�^0�T�t�#�f�y����;ƭ�D��q�Լ�.>%�����x��|��(�=?mY@=\ɣ�<蚽����V�=���>���>7���0�0��Q�#Kp<U�>���>��>0\��T&�Q����>xK?�d?pI�?�揾�i�� E�6����{�6���?5��>sf�>��>���=u������#pY���D�f��>Դ?����]=���;���:���/>:!?��>s�?�O]?���>,g?�?5l�>l�>��B���ظ,?@�~?C�=Cc1�6U.���>�$�C����>��(?+�V�>�G?��"?!O0?}�T?��?S>֘���b<��2�>)|>�S��Ǩ�5�[>��R?�>�7N?P�?�=>^	-�4����Ƚ��=��/>�0?t"?g?WL�>��?u
�����= ��>�Bf?h&�?��d?�p#��?Qe�>�=�>r�4=�.�>G�?�8?�]?t2f?<�-?���>6k=���"�����N"='w�=1�g���r�61k����<�#���s=qt��c�-�<I�@<}�<�0ּ�[�<�_�>��s>����&�0>��ľ=D��U�@>�]���N���Ԋ��:��3�=���>��?$��>�F#���=0��>� �>���)A(?��?R�?x�;̚b��ھ}K�f3�>p�A?�a�=��l��y��/�u�A:h=��m?|z^?o�W����T�b?��]?h��=���þ��b����a�O?<�
?Z�G���>��~?c�q?v��>��e�:n����Cb���j�IѶ=Pr�>NX�I�d�t?�>s�7?�N�>�b>�%�=[u۾
�w��q��_?w�?�?���?+*>t�n�K4�����#�� 3C?U��>� ���� ?(]���˾!ؗ��:��P�ե�����
׊�1���*b��﫾�aN�_�>rZ?�_i?�Yi?��X?Dl�]�s�Z��~���V�Q��U%��O���A���A�m�_�!�������ŭr=a;�>P�w	�?��,?���=7?5k��s߾�����>�Om��K�4%>s[�9!�=��8>�g$��,"��٨���"?K�>{%�>�%.?2�j���F��X�:�Z��e*�V�S=3~>�E�=��>�ǜ>�)�F���ξ�������v>��c?˵K?{�n?��մ1��Ђ���!��)��B���8B>�>H�>
�R��c���%�=�=���r��*��@����	��nv=��2?�f�>}ߚ>��?��?�e	�붮���y�@�1��#�<
9�>�Ei?���>R�>_�ν�!����>��l?���>��>햌�oZ!���{�ЧʽD&�>�>��>��o>;�,��#\��j��R����9��u�=)�h?���O�`�T�>�R?M�:��G<�|�>�v���!������'�5�>c|?���=u�;>#�ž�$���{��7����.?7	?U��������>��!?�c�>|��>���?~��>�繾�`f��?�/^?�M?��C?� �>��=�2��Zν��C}=?qt>��Q>-8�=�b�=RE!�VZD����,S<�\�=O&�˿�}Y<͊ʻf\<�R@=��7>Nۿ��J�)�پ>	�����	����I벽�b����	�P�����q�x�;F�w�'�3,V�3�c�0.���m�;@�?&�?�ē�)^��u���҂�����$b�>��o�_q��S4��w3�H&�����!��!�[�O�C�h���e�NT'?���ǿ���Jܾ� ?� ?D�y?F�S�"��e8�� >���<)��D��ԝ����ο�_?Y��>����U����>��>reX>�7p>�^��瞾��<ǅ?$-?���>�r��jɿP�����<͓�?��@�A?n�(�Uz쾔/U=�E�>��	?t`@>
�0��1�똰��k�>M0�?a �?�M=�W�C�	�΃e?�<��F�<6ӻA��=�,�=0=���<�I>�|�>��� ?B���ܽT�4>M~�>�Q"�=��;�^���<G�]>��ֽ���SՄ?�x\��f�ʠ/��S���[>��T?�)�>�J�=z�,?�6H�F|Ͽv�\�,*a?0�?r��?��(?bٿ��֚>��ܾ��M?�F6?���>Hc&�O�t����=�7�H�����#'V�Y��=���>~>�,�����O�`2�����=� �%lƿm�>���)��T#��Y= '��m!��ъ'���ֽ�-��_a������='Ҥ�cB< �@=���>��>�k<?N0U?+6�>�<>Xǽ35���Qھ�ܽ�S���������D���7���B��gȩ�o|��4���$�K×���?��#�=»O�.�������1^��MF��~,?�>��Ѿ�LQ�x@�c˾� ���ļ����4о�64��Tj��	�?�.??�u����O��>���/�P<�P?,F�������}��=���l��<�Ҡ>v1�=X�޾�o/�XW�߂0?Q?>�����EI*>� �/�=ƻ+?��?/�`<��>Q'%?��*��\���[>q4>��>v��>1�>v����ڽ�?khT?������l�>�]��z�z�Qeb=��>�5�g�鼞>[>�ؒ<"܌�NV��ޏ�Bļ<�-?���=HB?�\�%�G�2�<��=&&v?Ї�>g��>W�i?��;?�.�+	þX�f��
��~λ|s?��s?���=���j ɾ�?N�WM'?�G?�G=�z��RnǾ�8)�˝��u�>mNp?{� ?��j=��il�����k�A?��v?E^��ܟ� ��iX���>�C�>
�>�g:�_��>)]??���z���W���4���?��@('�?��g<ȑ%�?�=Y�?��>
wO�X�Ǿ˪��bb���v=K+�>� ��_�t��� �oo/��6?�ȃ?���>�Ń�j�0B>�b��.��?�?�!Ҿ�O/=֝��w��\Ҿ�p�~�=�p&=���=����|����l��5U�G\|>�@x�b�u��>|ܱ���ZDƿ����fž\vB�3Y?���>�熾����\K��u��o;��D�d_þ��>:K>�r��򃑾��{��Z;�T.��6e�>�w	�$�>�iS��E������0<���>r��>���>�d���N����?�3��&ο�������әX?4T�?dz�?Pj?O"-<cyv��0{�;��G?��s?,%Z?�%�12]�6�7���?<9��ʚ5�"�@�6�>�8���j�\?c�?_tJ��Ց>h�>D8�>2�>`+�����_C����g=\ߨ?�~�?v޾p�>nV�?6�>R� �������T��������V?cɈ>���G��sC��;۾b??��C?6㐾����_?��a�d�p��-���ƽ(١>��0�Ed\��A��ԣ�<We�����=y����?�]�? �?ϳ�� #�5%?>�>���D9Ǿ��<i��>{&�>0&N>�D_�ɰu>H	���:��h	>���?~�?si?��������.S>(�}?�%�>"�?�z�=�b�>�h�=��,��g#>u+�=/�>�|�?�M?�K�>P_�=��8��/�^ZF��FR��#���C�y�>��a?"�L?�Mb>����!2��!�roͽ�b1��0��Q@�?�,�Ș߽@)5>��=>�>�D��
Ӿ��>8nJ�~�ҿ����{�־D��>���>��?��B���仁� �Z�Q?�z�<������3s��(	>S�?yR�?F�?2S��ʂ<VE�=*��>,�a=�A>Q�|>�멾S*սi]w?/�N>�8o��$辬M=���?r[ @�i{?�3P�=?O������N�����D=��^>�8?sR���u>���>�7�=�ly�듧�A�w�旦>�ڰ?�?���>�j?�>n�ڮ>�c�=���>�c?zO	?�Z=�m���>��?T�����F���*3_?�r
@�@�wU?�W���b���i��4Ѿ���V�u�=^�9>����L�=�7%�����>���>}��>@�5>#6!>M�>>&3y=	>&ۄ�Q�kȿ}���ݮl�5�!�(����_��[�Ɵ����>����+��݇�!A⾉�ξ�J���N�� �\=�z>��@?tSP?g0v?��?oZ�C�U7���i�=k�B�p��=8�4>E2?�6\?�5?�>oa��0IU�3�l�Q͋�bN��\l> 0>n��>���>��>��=�\B>�_>Ok>�0=Ĕ;(J/��̣�%�E>0��>���>�f�>_
3>��>�ճ�LQ��"�f�S�x��ͽ��?�̝��L�" ���+�������=�-?4 >�����Ͽ�����=G?厘�����/���>Е/? �W?��>+$���Zb��J>���_n�O:>�r���(j��)���Q>9!?�6G=#��>�[��F���5��ԓ���>	�?򒾥۾����URs�ji�$��;5ݳ>��k<�� �Bn���炿�]�P��=v5;?�X�>pR��达s;q�|L��=5�>�(=�!�<!��=>	�=6YĽD��xq�*⇽@��=�#�>��?$&�=:I >Y�>Y���|
�
�>7��=��>`&H?k�!?W��O�� %�)p���>Ak�>i�.>M���8�w��=E�?y>`�"�(&�����E��Kq>(T&�˝��W���c�=�j�ƥ>�����78�%�b���=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>���ُ�����`%q�!�<��g>�S=?����>?�=;�E�WE�>�>?�=	��Q��'�ȿټr�64?4��?Tӛ?��o��f���&2����>H��?�x�?�D�>��A�����\>@�S?-�d?��?z�	��곾�n?�W�?6�k?0MJ>���?]�s?��>�8}�y-/��,���������=��k;t��>�>����>�D�M_����wej����_>�/#=��>=�P���
g�=J�������j�g�>vMp>��I>���>�  ?Q��>*��>�=������8Ԗ��K?ɱ�?���3n���<ʹ�=��^��&?�F4?�[���Ͼ^Ҩ>��\?ƀ?N[?���>��B9��忿�r��T�<[�K>(�>�a�>oi��ΉK>��Ծ�7D�8p�>ޗ>����5ھHH��A���/9�>�i!?���>>�=Y� ?��#?^|j>z�>\E��2���F����>ԛ�>-K?7�~?��?ܳ��Bn3����x⡿�[�N>7y?[o?ʗ�>���������H���H�bQ��u��?a=g?�M���?�2�?�??o�A?��e>�D���׾U䫽B�>�?��=�[ாl�=��P ?��6?�&~>�>M���ӽ���=�;,�؆!���>�>O?�76?�Y;�|b�k����=6���E�1=�qW�!�=&�[>i��<�#s���9=f,g>v5�=�M��CO������!���U>C2�=G\׽�V+�� 6?}�����C�����l�[�q��՝>�ݩ>�2޾��e?4�}���C����W����ڨ��9}?zp�?�B�?�	��mnj�1k??އ?�R?��?y��k��{%�V��&?����!���v>�2>{N���QӾ�T���J��9y�bǛ�F4���?T>��=��>�6�>�.?>��O>����:�u�)�l8�&�[�?)
��,1��[#��/>�L3��/a�s�>庾�M<��>�����:�>:��>�>%��>���>���=s\�=H�>�׷>�yG>�ޮ>��>h��>�}�f:l��%R?���c�'� �����)B?�Nd?`�>�j��������b?�s�?f�?.�u>E�h��U+��w??z�>=���m
?;=����-�<O^�����m�����OP�>jWؽn/:�M���f��q
?�?�ď���̾�E׽������=�<�?{7?�\$���I�ٝs��uJ��.9���a�o��?¾�'�s�i����q�rM��ע2�\F�<p$?"�?�������뀘��Th���G��{O>���>��>O4�>F�>'�	�V�?�2o��|,�����P�>���?���>J�R?^5R?��L?��_?^н>1�>a��9m?��>�7z>�n�>�>?��!?��F?i�7?I�"?��)>M��uԾSIA�b6-?i�?�T?Pw'?"?�#���U����=��=�d�Db<�� ���:RC�*����!>�n>]��>aΘ���J���UP>��5?�^�>L�>�-����g�A�>56�>��>�#�>�Q#���i��[޾��?��?���[��=p�6>�GW>��½���2��=t"��SW�=�Q�<'����Q����:>Ma=mR�=$���YN1�{�=��=
u�>,�?���>�C�>�@��B� �Q���f�=zY>bS>�>�Eپ�}���$��y�g��]y>�w�?�z�?>�f=p�=��=�|���U�����U������<�?BJ#?XT?T��?��=?Aj#?��>+�`M���^�������?�+?��>��7�ʾ㨿�k3��v?k;?�Ma���\T)�A�¾<�ս~�>�p/��U~�j����C��\N�b��*�����?���?�u?���6��T辽���:}���SC?P��>4�>���>��)���g�}��;>���>��Q?V9�>��b?2Ղ?�=R?���;��s����s2��c�F>c��=��?�,~?�Ag?Y �?E?��>B~���C�!�S�Ἣ��W���O�=�ֲ>�(8�P�>��?��l<*���ݳ<���˾p/�>�̇=��>A��>g��>�+>X�E���G?���>I)��j��������3�<���u?��?��+?~=�}���E����;{�>�j�?��?4*?��S�^��=1+ռ�����q���>��>xI�>�P�=�G=2�>��>���>�J�!k��]8�vgL���?�F?q�=�����2�<�����¾%>Q�*�w�d�/ړ��䵾�&�M�W���Ծv���6˾*�����پ�a��RG<����>T@>�*>���=K�$�v������=?ܽCW�=���=��r="���>�A�1�iP�=� >LN�=���ۼ��}˾��}?�1I?��+?l�C?g�y><Q>�3�}��>����r=?��U>��P��~��}_;�������r�ؾ�׾��c�c���A:>�TI�9�>�@3>�N�=H)�<vC�=SDs=�ˎ=e[S�.m=�)�=�N�=9��=A��=��>;S>�6w?X�������4Q��Z罥�:?�8�>Q{�=��ƾq@?�>>�2������yb��-?���?�T�?;�?Iti��d�>H��x㎽�q�=P����=2>`��=u�2�X��>��J>���K��7����4�?��@��??�ዿϢϿ5a/>�d�=��佖a�� ���T�+}�蹻�?m�D�נӾ���>��=���r����䒽3fG>R�E>_ֿ��LK���=3�%���=;�<��k>c�>&��<�����b>a��=�o�=^�=�K�=��=)�����=1S�<�g>��K>�I�>8<?�91?'e?�'�>2Su���Ѿ���Ȧ�>���=�ó>4=p=xI>��>�o9?�]D?�~J?M�>k2c=ވ�>�!�> �*��j����O�����<�;�?v#�?�4�>�l<�>?�����;�S��?��-?X�?Mu�>�U����bY&�њ.�#����g-�+=�lr�.TU�M���Ul�v�㽲�=�p�>���>��>Uy> �9>L�N>p�>Ǫ>:�<'q�=���7ŵ< �����=h����#�<wż|���uZ&�7�+�h�����;���;�]<U��;�Q>/��>U�Y>�Uv>��@>k�վom.>6��i?.�e?�=���lT��m�_�e���@-�**�#�7>j�|>E��;�o���%?:(�>։q>5��?o�?���=�I{��`m��R��[��<i��xw6>��D>~44>?	���e�@�-�<h���>b?{>�e�>՛*>���7��Q6=�-ھ5�3�=��>�x��"1����7�	%p������Z���Vo��=LL?ǥ��+:*>6�z?~F?�̒?b��>
n�J�ԾnBQ> 雾�ռ�}���?� ����1?�E?���>�����=��3�̘���A>�f��C�c�D����].��:4�p�Ǿ�M�>��ᾄ;����0����,���ncY�^n�����>k�Y?Op�?���Bv���4�Lw���� ?9�T?h� >5w?�3?z}6�Öھ
����	V?@c�?��?��N=�*=�=_��>t��>/�?��?��j?�)���?��=�q!>s#=��^>h�=j=>�0>:J
?k�?�t?����%C
��]ܾ&i|���\����=M�м Z�>���>�>�!>JQ�=8>��W>��>).�>�T�><R>��>���V�Q�?�*0>P��>�G?�ac>C>e�G>��=&U���M=9��l���м���=TC�<���=�m�=�?�|ֿ^f?�E�>X�S�?ص�QE+��E]<lF[>���`H�>�t>�ɮ>AZ>$��>��=U� >�=_�$�ί�>����@� 1O�-�5�������=�*��8U�q[��p���ל�*S$�z���Le�_�{���?��(s>=�}?|"��J�����M�bb?�2��>��#>��?�J�L'�>�u�=�?���>���U堿~����پW��?��?��]>��>�$S?U�?��4��)$���U�Rv��?��-c��_�s��������
�R�����]?o�t?��8?P��vj>�H�?$y����� r�>�.��<���=���>e}�y��$۾ꙸ�m����R>G�j?B-�?��?�JI���>���>�X?w�R?a��?o<?�,?*|<��^?��>V%*?�|?j�^?m|4?g5??�*�>+��=�+�<�ؼ����R�����g�����"=��=��=�ͺ���=���=T1>H��=v��;��d�����V>>/�=�� >�{=���>4I]?���>U��>־7?��7�������.?gpS=Ad��Z��|��ˍ�c>*�j?kȫ?8OY?ʓ_>T�?�?�D��`>Eъ>0�>�^>Q�>X���C�؏=��>>-�=�qR��p����	��ؐ��	�<(�>	�>[�z>م����+>�-���q��{d>�S��b����S�?G��03�%�v�ю�>՚K?Ul?���=��-���)e�7�*?�P>?q�I?ٽ}?�X�=_�۾|7��G����˜>��<F��1��"���ί9�[�9��p>VI�������G>�O�>��a��uC��ھVR߼E�!�B>=C��WQ��l˾��0=�{�=8H˾�����������X�Q?]�>߱�y���9���eL>	�I>���>�w�<y�ʽ��O�@���
:m=���>��>�1X��H �l�K�KҾ=��>ĢF?}i?��?�p��8���'�H���'���O��e�)?M�>�?��>��=)�i�����w^���H����>��?/UB�f^9�Z�~��e����k�>��>������?�7r?�?�i�?�oA?ӫ�>���>�ܽhr��t�$?+i�?��=1�����>��;��C�F�>w�%?��0�bq�>$U?�?��#?]�T?hC?:C>�%����B�3��>a�>�L�<v���/j>S_G?ⲯ>�b?qm�?��->dp5� ���3/�}��=�[>|�4?�?%�?0�>��>�?,�G��>6?3�?�?�K?;���,o?���>??���݃r>���}�&?p�f?�5S?�C:?\�g>r[r<y>彐��{���å���Ƚ������=ð��ʽ|���U�=y��=3��=`u��f?��lQ����/���=���>�s>W瓾:�0>!�ƾ	d���>>ܡ��Ԛ�������7�.��=G>9� ?Vq�>��&��=4�>�X�> f�%�&?b?��?�4;exa�A;ھ5EJ�~2�>W2@?/*�=ׯj��ϓ��t�V�o=(o?E�]?��^����w�b? �]?Ϛ��=�j�þk�a�W�?P?�
?@{I��>UJ~?"'q?4��>Wrf��/n��ꜿ�&b�
mi��=➜>4��X�d�[R�>&�7?��><�a>���=s�۾�x��
����?
��?u��?N �?�*>�n�@�9`��W����b?@c�>�0��^�&?�zT9gvƾ�>�����o:վ�E��(����ݑ�����ߩ-��ℾ������=>4?.�g?5v?�'d?'5����c���_���~��W���n���_D���G�(�?�D`f�������򦾍i���J��5�?��.?����}Z?���V����W>��{�����h2>5P~�}�=Y?N=�*M�J���,���1?�%�>J�>��N?��:���K�Yr:�yA���#Rs>z��>�K>-��>�I��H|� b,=�d��d�����?v>-�b?��J?)\n?63��0�����%�!��,��֩��ZB>�>�a�>3�U���o�$�y�=�?s�4:��m���i	�9~�=:U2?vV�>5x�>��?��?m?	�����bxw��n1�[C{<G�>qh?���>R�>��ѽ�� �>p�>�a?)�>�V >��]�����y�ׯ��ٝ>��>Y��>��=�[K��*S��[��话�I�R���G>�?������6��x`>_�X?���?��=���>��*��M�s� �Օ�����w0�>���=�M>��i�y5����G[�N<'?��	?�ɍ��&�{��>�w"?Q"�>���>!��?�Г>����$q�<��?3(X?�H?+�A?�_�>�<�<^���i�̽�#�d�!=l~�>5S>=3 =I �=љ��Y������~=T%�=�R�]=���z�<k��9��<;#�<Q9>ӿ�\�z����:վ&k�1��Z\�8z�����vI�r���䠾�о�:
����;����=�=����7�.x�?��?���=}7~�V�V��J��$��>�?$�[�*=������o�=���"����Y�k�T�4�!��)n� �B?�0�뼿}����z�7�>��?���?:��׾V�;��+Q>�}�<���=�ᾌݐ���Կ�����?��>���1��n>�>��'>���=�r>sb��8&���k�>'
?��:?D-J?����2¿t �����<!��?�@زE?�P!�������	�>%?���>�~��0�~j����>�Y�?�k?�c�=T�m���"o�?�0:>D�,�ׅƼ ��={�=7�={Ё�P�]>��M>���p罂��0N�=�x�>NU���a��Q���=e��=W<X�� Z�5Մ?+{\��f���/��T��U>��T?�*�>W:�=��,?X7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?_D6?���>�d&��t����=�6Ἀ���y���&V�q��=Z��>_�>��,������O��I��[��=s��xL˿�	 �p~�Z~�8s�P��������hҽ_���Qp��GV���	>I�>�a>ְ~>5B>��{>Hq_?W�b?ᝫ>�YG>صĽ��}�����L0G<�왾�.�xpk�3U�������־}�!��,�d���Wھ��9�"��=\0T��|���J"���`�cF��-?�m>r;�@L������ؾ1��E��_�ҽA�;�7���i���?�E?���p^���7�Ӽ��۽�]?;�½���J�����=��[��b�<�Ԕ>�ٞ='��]2� 1J��.?��?G ������f(>���x�<^(?_5�>!�:�.�>�#?#�/�=����gY>%_5>Q��>���>F�=�ͮ�� ݽ�q?+S?,�����2��>j����y���\=��>;�0�8�	��aY>*S�<Ä�Q�	�*����]<�QP?�j�>d<�;1;�X������_�=���?\��>�q�>
�B?�zB?�=��߾�`���9���>��x?��j?�S=��0<�T���ES��7?ԫK?����_���.��5�v��tnh>��V?���>�.>�s�GG����ώD?A�v?\�Uk��V���dA�I֭>H~�>���>�w=�W�>�;?��置i�������8��~�?D�@un�?��<�>��-�=�?���>�@�O�ƾ�R��&���*Jw=��>�L��H�l�{�Y�B��j<?{��?���>�j��P� ���	>KӇ�^Q�?���?��Ӿ7�,<�1�'�e��;z=��>]�;�k�<d�ƾ�$�]������n��o,��d>��@<m�� ?�T;-��ǿ�勿8�߃���?�=�>�ѽ��4�G9���8���X�W�ž���>5�>�-�������s��7��L
�>n�=��[�>M.M��hþ�õ�+r��>t�>�g>9��񿾍��?5��ʩ˿?a��C;���S?
֙?�8�?� ?PcB��N���^��z�;��H?�lm?�iO?�:����W��4<�ap?�z�6�m��"I� �	��c�=��>?�#?��M��z�>�A�=�)G?t�i=��o��*ۮ��Qp�p��?�?�����?�!�?E_?�-�������Ѿ<���Vq�>�<�<����c��zf<���� "�=Aq�>;�c�ZW��X�_?�a���p���-��ƽ�ڡ>��0��a\��U����Xe�����Fy���?�]�?��?��G#��5%?
�>𜕾h:Ǿ���<|��>(�>B+N>n_�H�u>����:��m	>W��?�~�?di?�������FW>j�}?BW�>w��?��=:w�>���=�����oA�Wd<>t�=T���a�>�F?gV�>�=�T?�W�/���D��zQ�_���#C�K��>��`?iA?^pc>+���I:�6������D�8�Ay��v5����Λ�D+>kDV>�P>;�Q�y���)?A���$׿k��2�x��?�?�� ?��=�e:漧��=n@^?�$>����'ʿ+1��&�}>�u�?���?���>��������F2>?= ?���>)���{��h<��&>6?�h<d?m��4��̴>���?P��?��?\�O�!	?8��X��3~~�.���7���=��7?`���^{>o��>��=�gv�����1�s��S�>�R�?tw�?:��>=�l?k|o�U�B�3L2=$��>��k?�j?��Y�6�򾋦B>�?y���玿��f?P�
@�s@�^?&ޢ�B�ۿ[+��܅���ٷ���=������=�h�F�O=���;഻�,Y<��=B�>�!~>��>�P>h~1>�>Lv��X�&�eS������k�D���!�����r�����9k�l�QW��	K��/��.���`���C�40���A�� >�4B?��c?16�?�9 >2����7>S�)��-�=�r��J&>�p�>�2?B�~?y�B?�9>-ǽA�L���|����/���~�>�zF>u��>��>慷> ɬ��N�=�[�>+�E>u����G=�9�"��cz>��>恒>�
^>"�<>��>%���G��Xh�´v�F�̽v��?>���d�J�),���W��]����=xC.?�Y>e��j2п�׭�&(H?xǔ��2��M-�˺>��0?�XW?h�> ����T�BA>����i�W@>*� �m���)�ϕQ>w�?Yab>��>��-���6�5'��ǽ�ŭ=O�?�5�����]���]DF��Fھ�J=��M>�nu����D����p���M�;��.�)?��>��ໟ���ϐ��eH��ֳ$>fl>攥�(4=:=b>����nl��q���==OB�=�.�=��?��,>Li=¨>�H��T�D�~��>�>��>�c9?�]!?������{ǆ�,���<|>%��>� Z>�=��E�9��=�R�>$e>�Ϧ����#b*��J(�ǭb>�p���2U�*��2�A=~k�����=؞=3����?�N�}=�~?���(䈿��e���lD?S+?a �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž5Ǣ�Ȕ	�,)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾA�>,Tν_Ü��֖��@������
?�??-"���=�=���>�ͥ>���y����ƿ��9�t?i��?y^�?Jq�=<��ث9�\R?���?�7�?�2�>9��rȽ%?%�X?^K?"�?�+��b�A�a?O�?��n?kI>���?��s?c�>�x��Q/��4��"���VN=?T;UT�>�@>����gF��ԓ�)d��C�j������a>~�$=Q�>z4�,2��nN�=N틽N���f�S��>?!q>s�I>�N�>�� ?�V�>���>�=�t����������K�K?��?"��|�m����<�=*u_��?J4?�_n��'оʸ�>�d\?N��?��Z? ��>���4���տ������i�<��K>���>uT�>������J>��Ծ:�C��>�> 7�>cY��J�پ�.����y���>�C!?���>r<�=� ?�M#?�&h>�z�>U�D��Б�e�E�<Y�>�j�>W�?p~?��?q:��RV3�|��&c��~�[��
J>h�w?�v?�R�>�x���"��.�8��#H������l�?y,g?���j?�7�?M}??�B?��e>���4�ؾ� ��6�>i�?
ٽ��-��A�R]B�8�?���>�|�=��<�>����ɽď�����+�>U�-?�?����Im��o'��2=Fۻ�$�<�&K><]�<�!�=5,�=`|��TZ=�0P>�>�������$>��=Wy>�t�(#��?�s,?!��i��U+=��n�wF��
�>���>8�Ӿ�)`?�,��Be��a���E����p��݃?��?.�?�����
g���>?U�?��?��>p���]��$�پ��N�^�{��y�#�=�`�>O�I�ξ����c�������Y��L� �?��>F��>���>7��>�J>��0�c��K�8���'���W�����J)�^l�F3�[�ھ�(����z;�;ľ�Hs���>t�C�?�v>�?ƪi>ˑ�=S�>�9���tR>8v>�:h>Ǯ�>���>U��>(�5>2ډ����S�Q?B޽�T�&��M������B?�d?�b�>��[��~��o��?Q?n��?�,�? �v>�Nh���+���?t��>$���H	?L:@=�9�<�䶾��큌���&�>-YȽr9��L�f?f�XY	??�?���k�˾�9ҽ����ė&=}�M?��1?ނ��sH�N�Z��Y��f��|0�
k��Sp����U���l������J��{�dD�|�4�i;?��?KB��	�n;����M�dM����>��? �1>V9>��=����:�#�nqR�(S"��ʯ�"?�>��?Pl�>V/L?��V?��r?K�W?�*{>���>MQ���#.?@�>��>�ݟ=5N�>H@�>�YR?�<2?��1?��}>0�ｗP������Z&??��8?�S$?�[?Ճ��������3�V+�=�,�@��=rʽ)�k���O�g;0>�{->C#?Y"��A1A�m�Vp>Z?���>�B�>�;�������l�<��>� ?���>�N�xҀ���%����>�t�?��u�j��<<f>�C,>�#���&�����=�e_�S��=pc��o4�;Mj�;��=�#�=�$`��e;�-3=3�����.</v�>_�?e��>�9�>�@���� �̯�8��=$�X>d'S>�>�7پ}��W#��_�g�Gy>�w�?�z�?��f=��=z��=v���S��������G$�<R�?�K#?3ST?㒒?(�=?Gj#?S�>E%��N���a�����@�?+B$?Ǟ>8��-�߾[��̨.�V.�>��?Xz[��uR��\?�V�Ѿ��<�=��;��΀�T/��S�P�s�D=����N�Dv�?�Č?%( ��*8����Iޘ�����e~G?Q��>�ɭ>9 �>�.�6�^�����4>X�?�I?�R�>|>?6�k?v�i?p�}��O�i��Q䕿6��;s�x�L?�͑?�;�?���?Q�?�`>��ٽg���\��>�����-���V�=�C>*bL>K�>�9�>d�>Ÿ��轈˿�I{y�0�+>py�>T}V>�>�MI>R�x��aG?i��>�m�����碾�,��L@@��t?ݐ?�f,?=z����F�:���EO�>Ll�?�D�?� )?�jT�jH�=A�̼����jh����>l�>��>'.�=moa=P�#>b�>[��>O��a�>�6�x6M�?̐D?���=�ſ'cq���q��藾 Rg<�I��#i�A��+�Z��%�=
��D�%����q]��ҟ����ᅵ�����`h}�'b�>,g�=�)�=q�=��<j�̼7n�<kI=���<Z�=�j���[<��4����(Z��l���Xh<!E=���tľ Fv?U�C?�)?K�B?�I}>���=�=q��Ŕ>�ҹ��	?[�_>6s ��k¾ʡ0�Ā��3L��O���ݾ��f�ed���=>0�8� >�/>l��=H�=��=�=��=/�ӻSiY=�*�=rɸ=��=���=���=��>�6w?V���
����4Q��Z罣�:?�8�>.{�=��ƾn@?��>>�2������zb��-?���?�T�?5�?hti��d�>G���㎽�q�=_����=2>���=��2�J��>��J>���K��u����4�?��@��??�ዿˢϿ4a/>�I>d�=94��� ������O̽�`����>�H��P���d=#�+>0���5!��v�=Cr�>&�x=����~}�>�=�&ӽ�Q���=/�=�
�=(�>Y۽@E�	��=s��=�w�=�aS��w�Qф��ۂ<���=�W6>Q�����>[�?�d>?�?u?��>��Ǿf�Ҿ��˾�[�>L�}>U�>$W�;9-�=�1�>ܝE?TO?c]>?n:> �\��;�>$e�>_L���f��cT�f���Ol�<��?}�?#G`>�z��W��(�H�N�0��:D>��?���>p�?���>8������%��H�2����S����о��� ����]�	N��;�L���>��>h5�>?��>�֜>�Ik>�]f>�T�>�g>~,����N<hN=��=3���g�:<j0�=0�K=�,��:����+>�J=���gׄ�N/��:��<P�"=`�=��>��>�
�>��=���,�.>lk��6|K���=%����A��c���}�\�.��9��=>o�R>p��ԑ�t�?�H\>��9>$��?O�u?k>��]�Ҿ�ŝ�F�l�� S��i�=	�>U�;���8���^��ZM��־���>�-�>,=�>�x�=����a��7Q=
3��3S'�r'H>�I�'�=?
�;��G�2i��Xţ���z��˗=��e?߱��5��>tI�?b6?9U�?0�?i}>9;l�Wi�>��P���q��$���5����0�G?LpP?6��>����[f�h����§<�q6>v1Ⱦ��l����`H�ֻ2<јϾ���>�� ��� �mtE�l�����o�G�������>NCI?��?�~���ih�~�`�W���T���K?��?�N=�>?��(?�k<�ᾟO˽�彝rF?wS�?���?0�&=W=�=��>�;?NJ�>M��?��?�?������"?�~���X>���!s�>��=�ag>�J�=i�>�I?n�?�[̽�a�^>ľx=ž���#�=:���,>���>:��>"]�> _>jbc>��>�!> �*>-�>�׸>A/�> �f�~P��/�$?Jl�=~9�=�@N?��>@�=�k2=�h�;�>O�z�C�>ӧ/�\���CRֽ�"�hD$>�<>�{�>��޿۱?6��>1�b���>�_���=,��(��_:�>��r��>P�z=(L>%.�=��>J��>�>>�]��`g��sE>�'��.��h7�{�/�,%�3��>���;k����$�ڟ�����5F��S2
��0b�[䇿Uo�T�=��?� �=��M�2ސ�tL%��{�>�I>��?��2���?�.ב�*?�P?5��A'����w��F��}{?���?P�c>i��>J�W?�?Q=1��3�IZ�e�u�&"A�s�d�$d`��������
�E��̱_?�~x?A?���<Vlz>ϐ�?S�%������>L/�^;���C=pt�>Z��.a�G�ӾW�þ���>�F>xJo?݃?7:?GT�S$�<bْ=N�P?"b+?a?+g:?r�?����3I?x�>/?m�>��C?��>g|?�f�>�}`>XO >F�����)������l�{�Iз�O��;���fļf݅�%��=�WȻjeR>��<sܭ�j��K�=��=��ؼW�=�ڤ>^[?��?� �>B79?B��#� ��N��>uC?�5>4#�����!�����zl�>E�s?	�?�iH?�|9>s�_�c�>��q>E�>�^[>(��>�p�>#��e�*�}��=�:5>��=��>(�
�W�������[��%=��>>,��>H'z>����O�3> 䢾t�u��m>�Nf��ּ�ԉI��C���3�񶄾$��>RwJ?��?d	�=,q�V���(~b�w3(?'�9?9`M?.*�?~X�=�o���6�,FF�c*�	ڟ>�Z;H	�*������Y9���n�cq>T;������>���}ھjRV�n�3�[�ɾ�ӆ�����(u��	���YO���j�=\����f��A����F?��g���վ��B��1>e;�>��>�K�?º����j��gۃ=x_�>� �>��=,���=>��#��Cڞ>�;?�f?� �?��K��󀿁[<��Y�g�p�Y9s<J�?���>�P�>��r>��v>o>��G+��g('��<3�֑�>)�?\�6�QK�m�|�u����`��e!>��>��C��F?�gX?��>:�?)?-��>�s>�D��Ý���&?2ނ?��=����.�9��h7�VzI��+�>~(?y�:��V�>�o?`?�&?JP?�@?d�>����D�>����>C�>�dV�+ݮ���g>՞L?|��>&�Y?Rn�?A�D>��7�����J����=�)>f�0?��?�?���>��>ݬ����>HV�>�:|?Vۊ?9�)?���=߆X?D�>Fl�>T~>R8�>yV�>�X?�e?��r?��p?��>c�,<�j��7���
����,4�=�Q�:BU�<����Y���;�<�&@;sq�<)�3�����K���}<�k�<�,�y��>7��>m:y��=`lؾ�\o�*P>�_K>���R��6���|>!\x>]�?^�=vPL�����>y��>v�0�c6?�B/?�z�>ۑ�-Q_�1��eQ����>�5P?_��>�U������o��x�=�Bj?xX9?�r������b?S�]?%k�R=�G�þn�b������O?��
?��G���>T�~?I�q?��>�f��9n����HEb���j�wɶ=�t�>eU�"�d��8�>��7?�I�>��b>(�=pt۾^�w��q���?`�?� �?���?�0*>��n�74࿶K�v���-ES?���>8#���?��<����6�~ᦾ���Z��ܯ���2��t�������=����H=V?�g?-l?'Sd?X8��mR�>T�\��L�]�vT�|����Q���A��M1�:�g����G���櫾�;=o����b�$D�?��N?�&��Ь?�W:��V�G����^�>�������=�
�= ��>�[<��$=��ν������_�T�!?�}><�>Y�z?@�[�m�"����)�.,6�t�=9�<Ӕ��#M�>�Jg>۳��%���Sf� ����q��ht>pd?zI?�~k?T����0�1��(�"�*<�E
�� CA>\�
>q��>>�]�b����#�� >�Һr����¼��1�
�[ Y=­2?�p�>J�>;��?}\?�W��3��Z�r�2�.�_ �<�@�>�ei?[�>)\�>�ս�R ����>n�l?S��>���>y���P!�U�{���ʽ��>x�>���>��o>A�,��\�%i��"����9��Q�=�h?�����`��>�R?�ܗ:��G<�~�>*�v��!����7�'�c�>u?=��;>�lž��]�{�?:����(?ei?p���w)�F��>LD"?G��>5�>��?嬜>4�����9j?w�]?YJ?�A?�S�>?�-=A6���nǽ|'�V�0=
��>��Z>wYr=V��=[��*@^�&���\N=�l�=��Ƽ����n$�;�Z���Qm<c�=,�1>� �`�=f��`��,��-�p��|<R��;��4V��ʾ�}���8��"�)�u�=X~��V���/��������?���?��w�H�n�d��Y�Y���}� t�>�l��^�E���4D��-+�kݾ��¾S1(�a0h��W����R���,?Z��lj��q╿5J���?(t#?��b?G�5�X���!��q�c�#���J������rƿl���Xq?��>�:��ob��i�>�Z>~^>I�>�̽����s*K�q�8>��Z?�\+?�b��$Ŀ튴�7|ڽԪ�?��@A?�a(�ȸ�bV=g�>	?��@>x�0�A�R,��?��>�?�?=��?*#F=�W������Me?��;p%G����J��=�u�=h=����1H>��>d���?�)Sܽ�<4>9�>�"�׹���]���<��_>N�ս啽;Մ?�z\�Tf�l�/��T��zV>��T?c*�>J9�=ղ,?#7H�]}Ͽ��\��*a?�0�?���?��(?�ۿ��ؚ>�ܾ:�M?�C6?��>�d&���t�^��=<-�m���d�㾤&V�^��=���>N�>�,�����O�gK��T��=�������
��4����/���ɾ+*���@����!��:�5��@k?�s��w��=C^�>fܫ>}>u?1>i?�`j?��>�)W>��={�X���	�2޽�Z��v����w��ZD���Ѿ?Ͼ�m'��Ǿ��D�p�%�b羋�+�k>�5T�"��M�"�M�M�@A?�w?�h=�޾z?�?uS���Ͼ�ž���t׮���5�B��_����?o0?��x���M�[��m�aH��8�N?�\�\4����in�=j�<�����ף>�Dc>~����?�J�W�?��?9�;܆�}�?>~�M�!<�=T.?\j�>��+��:p>�u=?�1�����Wq�>q��>`�>�`>IXĽ�N��&�	�:)?1�I?͏&���jh'>�뎾��Z�@��=�-�;���H�X>f 0���ž^��;G+���5�=DW?�[�>,�)����@���$��D=Ix???�n�>k?�IB?.��<�g��K�S����~t=N5W?�i?Ծ>
1���;о�`��!U5?dMe?��N>�Qg���龥B/�EK��?vn?Z?����}����Q����6?��v?s^�xs�����J�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�%Þ?��@���?U�;<��U��=�;?k\�>�O��>ƾ�z������?�q=�"�>���~ev����R,�f�8?ݠ�?���>��������3>d���Ȩ�?G�?#?��(s��خ��xv�h���1�Z_=��\=<x��3�B���t�Ⱦ~\`�`9�:��Y>@��i�]>L���r�㿗uп}�E��|����7?���>��/��|�����p���:�wL<�LX���>"�>��̽�S�$�]�B�$���Q=���>�p���>��l����z��K9��>�<�>�~>�y:�E%���?<���b������)Ӿ��^?N��?�"\?_?�>T��4����p
��\Z?��g?y�0?�4佧�$�*��=�P?�#w�{�n�L�1�����a�>֡:?c��>�>�8hb�(��F�>��>e�߾�����)����&��]�?�>�?=���R�>�j�?s۲>�E��X��9� �A콾�����!?��7>��[��*R����t�I�(�+?�_+?���A(Y��_?��a�7�p���-�g�ƽ��>ԁ0���\�ڑ���R��Oe����a�y�h�?�T�? �?=��J#�D-%?V�>9���:Ǿ�0�<on�>�2�>�9N>��^�G�u>&�t�:�"Y	>F��?<z�?�\?��������C>��}?���>K��?�$>K*�>}��=�᝾s���.8#>�#>ݦ<\�>
uM?f��>�o�=�HI�8�%�2E��7A����R�G��r�>��^?��C?	0�>�z漚�{;��'�z᫼s��/u�=�� �O� �w���s><>>�4!>{��w���g}?��U�ؿN��c�&�2�5?��>��?�b�A�s��N!�|�\?���>ؠ��j���Ќ���
�ۢ�?g�?r�?�5־�]����>׬>��>iӽ9٤��^����7>5`A?���u�����m�aň>��?�M@�z�?�#i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*��Կ����Wh���'���8=�Tc=�N!>K/���L�=�m'<*�żū��#>�Ά>xpU>Y��>�H>��:>�#>����i�$��l���J��	O�	J3�B{�Y��N���l�v��A�uX���-ξ ͽ	jӽ
R��-�QI��0{��(�=lTU?\R?Оp?�� ?Q���ה>:�����=<d�˕�=���>��1?�3L?,?��=�@��Hc�1���_��f������>3tI>�?�>���>Sŭ>�y�:5)J>�=C>ɀ>�w�=�6=(����=�R>,!�>N��>�}�>Q�9>AN&>����$���f��{�UϽ�u�?Oz��R�M�ZƔ�
ŉ�ư�9�\=�,?>>f����Ͽ �����F?�O��D��6��
>�r.?3�V?�Q)>���C����>�ؽbEg���=&���>�I��$%���C>��?��%>���>�35��f�<�e�B���6�c=n��>�T��}��z�w�O�I������=�cK=�� ��sL��y6a�J���`>K�S?�b�>�朽t���i]���  �M2�> D=����z�2>�Ֆ>[r���q<,��m�=��J>��ν��?M�5>���=*��>�(t�U�L�4�>(C>�IV>(vA?�L?� �������m��[�>\B�>q�>0 �=�N�#L�=�n�>�O>�=f���]����6C�һ�>Y�m��h�"�����,=3������=��o=:��"A���=Q)�?�ɠ��A��<�~�ý�??��&?���=`�༙c&��o���I��i|�?C�@w�?��X�{�?�^�?8�����=h�>%f�>���&�[�u?��%=^�����pq����?�?^/��܆��O�@R>�1(?�򾾇J�>���몣�;�v�x�=mѦ>r�i?!;)����Fg:���>��'?Rd��e���ܿi���Ƨ?�p�?�w�?�B^����8���U&?c&�?G�]?G��=L��6��=R�2?G�f?� ?l6�BW_�2�?.�?�Z�?��'>�w�?Iz\?o�>B߽��0�J9��?͏��Xr<ꛋ�m�_>�h�=ivžn[D�����g��>�f�|����>|�=��>���>��R�	>ށK�����L�����>�dL>��|>�g�>W�?�>���>�=t����a��X���K?���?����2n��5�<g��=r�^��$?7G4?�+\�O�Ͼ�ը>o�\? ��?�[?�g�>����>���翿|��c�<��K>�7�>7G�>�"��uIK>��Ծi4D��l�>}ї>@���F>ھu/��� ���H�>�e!?���>�ή=�� ?��#?F�j>D(�>�`E�`9����E���>���>=H?��~?5�?mչ��Y3�[���桿�[�X8N>��x?TU?�˕>䎏����udE�nPI����ٛ�?�sg?U�?�1�?:�??�A?�)f>���lؾޱ��z�>��/?f��'�4���ZĽ��?Z�?���>	þ��k�=��+�*L5���0�6@?~�L?��?%[�"=f��߳��@�=�}� �o���t��d��tb`>�D>��H=ی�;��8=�ߢ=�Kb�LQ��z>^d����>+���|B���*>F�+?�E��ȃ���=VZr�"lD�� �>�L>����<^?�i>�~�{�R欿�d�� �T���?���?�-�?B���
qh�;=?�(�?�4?�x�>6�����޾�ྜ-v��+y�H���� >z2�>�l��Q�z�������8���ý7����?�:�>�I ?��>��>>��>'L��)�#�Jw��)�_�X�:����7���+�ǳ�h#��Iz3�$e^�ͻ��]v�g�>�"e�u��>a	?
�n>ןo>�k�>�N�Ej�>[U>k��>kו>�*|>	O>i�=y<ЋڽI�V?e����#�j�k��+??��q?W<?�.������8"��!?��?L�?��#>'f�}N*��?�E?%�����?��>�r���ﻐS¾ЫM�M9�<�s>�f��>�ڽ�%��b1���n�j��>?���<R̾�������o=�G�?E�(?��)�d�Q��o�W�W��S�L���1h�q��G�$��p�"폿�]���$��.�(�"�*=^�*?��?�����+��+,k�?�hjf>z��>#�>۾>�eI>��	���1�,�]�iD'�䱃��9�>=L{?^e�>�)8?s}Z?�\?�f?��9>�>9����#?w��>Dp?���>4�?C�?&HO?�k?N�?�V�>�T"��羉����?��?ϝ?���>�?�u�&��=��
=|�o� ��E�o;i�̼��t�����I�9>U��=V=>�I?�G���r��n�t�>E�<?��>���>�bվ��������T��='7Y?f;>\.P��D���J�fI4?]J�?&��)G=�>�A:>���<�Z0>Zv >r o�gj�=�K<���6��ΐ >�h >\6&���=�v���?�J�4��t�>�?���>�C�>&@��� ����e�=TY>xS>\>0Fپ�}���$����g�c^y>�w�?[z�?�f=�=���=�|���T������������<.�?�I#?�WT?/��?��=?�i#?Y�>�*�DM���^�����^�?�n,?�>h���>˾𓨿k�2��C?=v?V�`�����*�������׽��>��/���}��ӯ�*iC��p����VA���n�?�Y�?�@��6�ڠ�^ܗ�v���DC?2��>�F�>̐�>v)�Osg��)��<>�.�>�QQ?Y��>C�D?Uqo?c��?\R�>A9�3������&�<�x�>i�?�.j?�D?	�N?�V,?��>'�7=.e0��7�@�۽!-�co�$����>w�>�f�>:��>"�=d�>�6��!p��l�_>+��=�%�>$��>%5>Z"�>��c�G?h��>�޾��$�}أ��肾��6�L4u?�y�?�+?M=si��F�|������>^=�?�Ϋ?a�)?�T����=�ּX��U�r�l��>u�>�>h�=��J={R>ѽ�> *�>�r�9�nB8�xM���?K�E?ݽ=�;ſ�`p�O�o������`<�����c�]X��IX���=����{��s����]�z ��^����3���Q���r~����>�3�=G�=7�=Y��<��¼h��<��4=�q3<�=0/e�JgX<�|A����΄������b�;�?=6�&���ʾL~?ҙI?Pa*?��C?��{>s.>A�/�˗�>+�l��p?O�Y>��K��D��~�;����������t־��Ծ��e��N����>c�D��>|q8>D}�=��<J�=-�d=�;�=i�!�pR=��=���=�'�=z�=x�>(b>�6w?Ú��o����2Q�-U�;�:?�:�>�k�=̀ƾv@?��>>�2�����Da�L-?E��?�S�?j�?�vi��f�>m���厽�g�=�����D2>Z��=��2����>�J>���J��ӊ���4�?��@ �??�ዿ��Ͽ�i/>w��=C��=3�P��l��*� �t����.>�$?V0�ӕD��-+>��>S����l�3y�>X�	?f��>_���x��H��}J����=��=nL�>�x=�Q>\˫=���=-&�=�K�=M�>_���)�=����GOo=���>� x>$��=�i�>�?*<?��?��>���2�Ǿ�Q����>b�>���>|U=��C>N��>��D?�#?�6C?+��>����>�e�>d��=S���ξ��E��З=p�h?#w?�;R>-�	���(�y�5�O���[�>`i?���>�ؠ>�������� �-5�r	�g}�~�:w�8�5��`�<�8������b>7��>���>��>��>�_Z>��a>^&�>�Q�=�7�<�B< e]�?��T����e�<�U��/'E=]A<�'<���͵���NǼ4@�<�^k<U��;��|�˰�=���>..>���>M�=�����/>������J���=_���V�A�̦c���}��~.��[3��E>|V>/Z���ӑ��?�;]>#�B>e��?D=u?iV>��h{Ծ�(���Te���Y��̲=�*>�>�l_;��a�ƮM�Pо�V�>��>n̺>�'>�#1���+��[D=����� ��|?Lk��-`=��νk:Q�Qk���ې��f��=n�D?����"�J>y��?�6.?�M�?�r�>�������>�l�)�V>y8��pv���0��U.?�h!?W��>%t��BU<�#G̾����۷>hDI��O�����ӯ0�x��Ϸ�뎱>^�����о$%3�Gg��������B��Or�^�>Y�O?��?F6b��V��3VO�1���6��Vp?
|g?u�>�J?�??q)��z{�Bq��Ix�=�n?/��?�;�? �
>#h�=�Lx���?t�>Ԟ?���?��Y?�
��?>�A>��=*>P3E=�?�=�JW>n
?i�?G�?��ݽ)��Dk�ݾ0���Q�=�`>�f�>��x>�Za>\
>��=lj=��i>��>3�>��>��>���>)u��\����*?F@�=ӽx>�PZ?�6�>�W�;� >0	�=$��=P��=���N~�=�����=���g3>w��=jb�>ݻ࿈�v?nB?�cF�-d ?����P��F��>�jM>��轞(�>��>�H	?�,�>v��>Ս�>ȟk>Ħ�=�i۾��@>��$*2��e�C�O��j'�>�l��_ܽ�T��K�j�j����g���U�`��7�b�Ȼ<���?�:�<>&��;����j�?�3�>ٹK?�E�D��<��>���>�2�>j��Z��ꂧ��5��&�?�+�?�2c>��>��W?v�?��1�$%3�}iZ�
�u��A�+e���`�ލ�����$�
�������_?N�x?EcA?��<X[z>͜�?e�%�����>/�s ;�MY;=��>P�� �`�-�Ӿ��þ��SMF>��o?~�?K?�bV����'�>��P?�j;?㪄?��1?'?����9?�Ȁ>*�?���>l�??.a?f?"
�>�U>�v�=��#<頖�'d���]�*��Lt��>)=_�=E_a=^�B��s�;H�_9��F��ǩX�T�����<�To=u&>D�>�P?Y�?g��>�nB?b���ض*�;:��F?gҹ=O�R�͟���,��3���#>�ig?���?O�W?Bu4>�1D� o7���@>���>�}1>P)k>�X�>a���U��_O�<���=Ѿ�=牻=.�랾�!����sӗ��'">'H�>t3y>D�����#>jꚾ�����h>P>F�}x����]�}DI�IY0��0x����>UH?ȡ?�@�="	��V���c�fY'?��>?"O?�x?�f�=��ܾx+<�
�E�H�+���>ռg�
�=����L���:�����b>A뒾��Ҿ��Q>����'Ҿ Bx�^�L�1���6,=F����h�U�վ,�����Ē��䜲=	�����#����������c=?�r
=;`���vx�����&f=�D�>Q=�>-B�=�O|�WI��+��:�=�n�>O�c>"��=��վ� H��)�Iv�>u�;?��`?�{�?�YY�.�r�KxD�u��h�� J�<��?�{�>T�?A�S>�3�=E2���R�>`\���@�"�>O��>�1�~F�>�&��b���>��?� >�|?WK?���>Y�g?��1?�h?��>�۽Ln��s�%?)��?�O�=�&���,9���6�U�D�n��>e�&?.�#����>��?��?{'?�Z?��?��>X��I7=�l��>��>��M�䇭�g�e>�I? �>v�]?��?�@G>�<�ц���#���Q=?�=ڎ2?��$?w�?��>�m�>bâ����=��>yY?E�{?d�q?Z��=���>n+>�$�>�7�=+�>��>o�?R?,�t?S9?bغ>��D<����>ֽ-�]�o3��of����g=�B�<���� K�>�~<�<
	;���<���<N�{<�{@�������B���>�s>�ރ1>�Rþ8&���@>-������ǖ��D�8�M�=�{>�>���>o^#��q�=��>/{�>P����$?��?f�?��};+`��׾0K��Y�>�A>?#-�=�8j��;��#�r��q^=n?��^?[��t����b?��]?�g�=��þq�b���龽�O?��
?[�G�Y�>��~?j�q?���>��e��9n����]Cb���j�Ҷ=�p�>uX���d��=�>��7?0P�>:�b>�"�=Su۾��w��r���?k�?��?���?-,*>��n�F4��� ��a���T\?r��>j+���*"?��'���Ͼب�����x\߾�_��0>��E>��P]����#��‾naԽ�O�=[?[�s?�mo?P�a?����j�b���\�]�~��$Y�Q����i@E�zE��VD��Dp�����x��8�m�B=Ϗ$���v��ַ?a�K?ń=�|8?�'p��þ=)����>$����4<E�>U�>>�R>��>�MB>�/� 	��߭?��m>��>�go?�AS��@�������n[�~@����>:o�>�m[>(�>��;�
m�y8A���	�+��>>���>�QS?��B?�)g?_K6�K3�Q�u��t#��>̽ymi�pQ�=���=e�>pTӾLJ½˚����BP�(b���|��� �⃍�
�G?�02>j<�>�ė?9??��پ�ޫ��+K�\=��g4>&�?�xO?F�(?���>��!�z&�H��>��h?��>n��>�劾K��ůy��wj�>�c�>�.?���>\I/�y�]�'���P�5��u�=h?9[���-j����>�M?�!�=�;}
�>���dB�E`��w!7�O�>C ?��H=&88>O'��6����x��j����(?�?�Ŏ�p�$�㯀>iF?D�>��>6`�?��>t+���;��	?�0`?�L?ŊA?�0�>��=`ý��˽��"���#=``�>B�Q>�cX=���=�i�&X�eQ��*=�b�=jò�����U��<�)�ңj<E �<<[4>IA迲 g��/�S���q9�{ �nD��g����q྅kþo��d@ӾHǾcY����录�����`�r!��H���o��?��?>_���}��Y��b��i���G\�>��о���c#Q����<�w�y��?d��CV3��q��}�/ h�%i.?��������6���-!��T#?=*?�A�?b%����g80�4�>�w=�ؠ<\(�6���˿��^�h�h?z�>���l���>w�>��n>���>F����b{�=�&�>�^/?�?2N���ǿI2��RK��#��?�@�6A?��(�� 쾚8a=���>%W	?j(B>�(0�� ������>�?Gh�?��H=�!W��b��e?���;t�F����X��=°�=&�"=n��uDI>໔>� ��v@�e.ڽ�6>r�>."*�,Q���^����<OCa>C5ֽמ���҄?t\�j
f��/��R��LB>��T?/*�><A�=5�,?�.H��xϿ?�\��(a?�-�?���?Z�(?Z濾WĚ>�ܾۆM?_B6?�>#c&�M�t�D_�=�)ἅ��J��&V�D�=��>t}>,},�J���|O����� �=���E��B��s�2������a��M���w� ��j����R�r8�&����S��b�<���=Ѳ�>db�>�|>�^�=�
w?�l?�>fP�>���Z�N�iO��4���/d��:�j�L�[7Ծu��{	�5n��@�:���~�\�ɾ�<��>=?��������/>W�^W���!?��=����`'���^�5پ�پ�jH�9
�/m�ms3�;�Y�P��?9�3?�ȁ��xI���;�*���K�$�%�T?�zb�M���#�����T=�^,��*�=eŦ>�)�=�5Ⱦ�n;���O�d*??�U���fh���/>ڶ
��F�<�$?q��>*&���>��"?NO�ɑ�"~>� >	�>,Ž>*� >kş����?w�V?f�
�*(��5��>�=���|�ꨘ=��=rS��ap�o�q>�<�<��?��e�<F���k� X?���>�]*�Vm�穑�@��oJ=�:y?s?Ѥ>�h?��A?{o�<h���%S�����jH=�lY?|k?�<>>ς���Ѿ�x��e6?�d?I,X>.�n�W�
�+����A?�)q?&j?���z3|��(������6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?w�;<��T��=�;?l\�> �O��>ƾ�z������1�q=�"�>���ev����R,�f�8?ݠ�?���>��������	>�쭾?��?z�?/���ٽ�Fܾ�u���^˾n��>Yk8<}��<q�*>�Cξ>K��K<�V���}��� "���\>Bd@	n��C�>������<ȿYB��a��Ɏ��\?4S4>'��J�C)���6����{�D1����u,�>���>8=��N����z��U'�x�����>����i�=D&8�)��`j���䣽��Q>>��>~��=�c!���ľ.E�?���f]ӿ?����O8� �C?B��?ܦr?�o�>zXm�������۾z���\�j?��?��v?N��=������tQ?eH����?]�4�5�Ձ�>�7K?E�? �c���>�D����?�`�>*������7���.�Ⱦ��?�ͼ? ��.��>z�?zF�>[�ž��a�v9���:�o�~=m�G>ro�;�i��ͯ&��+.�����>O��>IIﾳ嬾X�_?'�a�E�p���-���ƽ�ۡ>��0�f\��M�����Xe����@y����?J^�?j�?���� #�]6%?�>_����8Ǿ��<���>�(�>�)N>I_���u>����:�i	>���?�~�?Jj?󕏿�����U>�}?D$�>4�}?hZ�=���>�t�=`ƈ��8�3�=���=�ܽ.�?�R?�H�>��"=�o8��o5��P=�Q�=�Wo����G��dA>o�e?�sA?�?K>�έ��i��
�*�Ҽs���P�Z���SI}���I��0>zU�>5�e>�߈����#?���ݿ�ؘ��z����8?b��>l�?�*)�<�E���_=�qM?0�>�		�o\���,���AZ�W	�?�s�?�c?�k޾�8v�*>�v�>�؉>�e*�M��=�6����R>�z??�Ľ�pQ�g�N�7�>�_�?���?���?>�x��	?���P��Qa~����7����=��7?�0��z>���>��=�nv�ܻ��V�s����>�B�?�{�?��>�l?��o�Q�B���1=8M�>ɜk?�s?�Po���k�B>��?!�������K��f?
�
@~u@]�^?+�zڿ���/%���۾�A�=i�0= �>����aI>#=.=*�����<��#>��q>��t>�>�0r>��8>��$>xC���#�F��ǀ����G���#��x�R6Y�����wq�����0��Ҹ�[㹽SR����K�3��,5�"���޺=�M?�P?z�f?���>i|佖^V>�.��7�=A?$�W%ǻkq�>k�,?��H?��0?aO�>IeZ�,Xl���x��ž��1�Z��>�&�=?�e�>
�>��x=���>RY>�2>	��=3� >� ��G��=�x>��>���>]��>��A>6{8>�ǯ�@䭿p�m�zt�)륽�h�?����fM�}V������ɾ���=4k(?���=nZ��:�οd����E?O��� �E{���=�&?�a?T�+>=����L��p�=8������*>��нwSN�m#��E>%?ʧy>9�=�-�8~���M�hq��h�> %.?`&����þ&4���e�����a�>�Ғ>m��=oS��B�������o���>�;-?�۴>p�\>b���8 ��_����O>��f>�6�=H��>F�J>t�;'<Y��{ �=�]=9u>�w�>S>5I�=��>'K���6��0�?�>��8>�% ?�E?��!{������r����>V�	?��g=�1G��.z�%��=�|�>w�(>V�?�J4���(��������>������*U�<gg->{Q���=� 6>J����]��?0=��~?�y���㈿o�9d���oD?�-?D<�=�zE<�r"������<��s�?S�@�d�?��	��V���?�C�?�����=^l�>�׫>\ξ��L�8�?�-ƽ�Ƣ��	��6#�;R�?��?ʹ/��ˋ�l�vG>[`%?(�Ӿ��>Fv�����F���w��]q�=�Z�>ʱC?��K��PP�0��>vN�>�:Ӿ�ˢ�{Gÿ����w?cR�?�ԛ?ET�=鲿͝-���	?�!�?�Q�?��}>dM��Ȫ=�~>rQ?T��?��"?�\�#�+���?��?8�?��>��?t�a?��>�<�=!%�	´�����k�=��<s!x>K��=�p�C�p�lZ���W�q�C�ˣ
�IM3>
ǜ=X�>-��������=o�[]־X�>���>CQ>�s0>�(�=:�>p�*>�ܖ>-�"��vN<�
_��B`��K?в�?`���/n��K�<䋜=��^��(?H4?[��Ͼ�̨>��\?���?�[?�d�>���=���翿8����<��K>�,�>�K�>\��&<K>E�Ծ'2D�o�>�З>�䣼<@ھ3�����|D�>�b!?���>�ݮ=�y ?�#?dRj>�w�>yNE����F���>=��>�?�~?~�?)���l3�D蒿�ѡ�|�[���M>G�x?�n?6�>W���oV���KY�wG� ɐ�ʄ�?�(g? :���?��?�}??��A?�e>�U�	�׾/���G�>2�?k�,��Q��{��^����>��I?�U>�#�<w>�N��=����*�Rz
?}�@?�SD?��X�kS�����7������ɼ�wS�����1ُ=�ʌ>ŋ]��P�=�i�=;1>��2�2����`�=��>���>O2J>w���-R׽�<,?�G��ڃ���=�r�xD�*�>�HL>k����^?�j=��{�|���w���U�.�?��?j�?���h�M$=?�?�?"�>�K���~޾<�྾Lw�W|x��w�v�>���>N�l�����������`F����Ž-�����?>7r>�D>
�?Z�s>=��i���:�}���<���4���ž<�[�v�7���$�I��B�^��%�=�qžYJ#��L�>��=���>���>�b�<'�<�n
?���<Q8�>��=��>BO(>2XS>iG=>���=��r<U�&���R?߈��(�x��7Y��?;@?��c?���>Hw������9�˲ ?�x�?% �?G�d>L�i�Y�*�j�?w?qp���"?O)a=�(y��ߎ<�W��!�=W��M<��ی>gT��x�9���K��Ok��?�"?��߼ӆϾ�LɽlAɾ�+=�|?�?	�/���S���t���V�w�O�����F0�oD��`(��Ep�3���,~��ņ�֚&��s#��4.?ڈ�?���ҧ�m���GV�k�2�n�U>��>c��>�4�>pm>�A�*04�:tp�Ǐ4�`ū��>���?�co>�=?MV?��^?�q?�Έ>M>��!���I?��=���=�>�g?��$?�g?�(?ZgL?�y+<�W=�O
��d\�h{5?�݁>d6G?��Q?U�>�JK���>1�H<�'��E��4�=�=6�?>�=�J�<h�>Ou�>͹I?�T*�9Vi�'��D�Q;�W?s{!?�u?T�þR<)����?W9?9�>@R8���t�����@_h?�?w�ʽaH���>�1>�б�y���z':���V~��~�=N���Z=����J=Vꉽ��	��$�=?��R�=�n�>[�?��>l:�>h7���� �ȼ��o�=�Y>�S>�>\Dپ1~��?%����g�hYy>]t�?Xt�?��f=� �="��=<x���`���������¦�<��?�J#?TT?]��?C�=?be#?��>u)��N���Z�����ϯ?�,?{~�>����ʾ�㨿6s3�-�? V?�Aa���KS)��b¾�ս7K>�c/��)~�b����C���l����Mɘ�^��?��?X�?�}�6���_���,N��
�C?C�>�	�>{��>˻)�W�g���:>�<�>��Q?��>o+?�Jo?�2x?���>uN_�ถ�"Ӂ��>�V�>m�g?��y?�:,?_֊?��#?]�t>a��:�ı�A��|���Ƒ��T���e��	�>�ր>��>��>X>=�6)�#5ݽtF� ^[=��>�9?tl >��>�A>P�<��G?6��>�龾_�8�������5��ku?�v�?+@+?��=I����E����4��>�]�?��?Ի)?�T�u�=T�ҼK9��#�q��"�>�p�>�!�>��=IM=j�>zo�>��>�w��3�C8��I���?��E?��=�ʿOe�&�v��
��'B	�i Ѿc��f.�k^|�c�����k����Z��f?��>���=���˾O?ҾH^��i��>�x�=���>Ԕ��i"=V�;������;t��=�Tl>p��G���v
���C<�����<W��N>Y�2=wOƾV�x? }G?J�%?��;?�{>͐�=Y�Z����>��Ž��?ʗu>&k��ež5�=�Rɬ��ϑ�-׾Աɾψd�������>��[� �>~9%>Ih�=�D=�?�=r�y=m_G=֙G��<��=Y1�=���=a��=g�>+��=W6w?��������3Q��Z�F�:?�:�>Tv�=q�ƾ�@?R�>>�2�������a��-?U��?�T�?��?�wi� d�>����㎽?n�=����Y=2>/��=@�2�ࢹ>��J>ɂ��J��O���(4�?��@��??cዿ��Ͽ`/>��)>V�@>:(<��/*�l ��WN��K���l?�[-�"�ܾ�>(�=�6���u��vˍ=�>��<g�D�XG��֑=���PA=f�<��>�?>�k=7DI���=��=[>Nq)>X��������^=/c�=`_U>N
'>F�>�[�>�3?��r?���>e����˾j���T�>��K>f�>�.0>>� >�?h�Y?��E?�0A?K{�>Ub���>Z@�>���U\��V�y>�=�܄?��y?��R>�Y����������z)�����>M?.~�>��>S|��J迷�$�f"7��_ӽj$���<�s�|�®�;`�н�m���E�=�[�>!]�>�@�>��>�$>��8>��>�>���<��G=���~��<�/��n=�����{���*3��V*���/�9_R�p�ܻ�ab<W�F��%�m��=���>�>%�>U!�=M����>�ĉ���Q���=������:�J�]��V~���1���P�4	>ڞY>B�$�c����!?��p>��B>��?��o?�3�=~��h�Ѿ�����d�oVu��v�=ER�=jm,��h6�M�`��wJ�fھ�<�>�~�>��E>h��<���y���v=��Ծ�)4���>lZ�E �=�y���W�����=��8El��j�=�~o?A�����>�t�?�5+?�у?:-�>Y�{���羪MJ>#r����g>ҿ
��0|���A�ѧ*?�?6e�>�S��W��@;2!��Q�>חN��mL������3�TDY�/��@[�>
a���Wо�H/�����1���)xC�ɑ��"��>�N?e;�?��]��Q��j(K�#}�h����?�`f?��>�?O^?�˿�:��sq�2i�=�(n?=S�?N�?"�=y�{=������>1N?�?�?5œ?x�j?5l;���?���<��3>u�Ҽ^a.>f8>��=��=>�m?^��>��>�1b�	����e�ͪ�������	}=��Y>F�p>��>)'> +�=S��=��Z>�n�>��>�x>��>�`c>_D�� ����9?��<4��>o}M?|mM>k~7�(	�>��>��>��/=�G>vJ=#�G>���>k�>o�;��b�?c���Հ?�&�>�8*���?Y����;w-̽�:�>?1�|�>�W>�:�>��>�0j>ݰ�>�y>3�
>���C>��־��0���e��rF�����h�>4	��?F|��ܸ��3����	������[��-��5�9�*ZK={��?�{Y�@�x�/�+�k���?���>��$?��V�Y">�i0��e�>�{�>�Q��a���C��� �-��?��?�Hc>d
�>1�W?[�?�{1�b3�Y[Z�ۣu�zA���d�̲`��؍������
����S�_?�x?�dA?<��<� z>���?��%�O�����>�/��
;��K;=_"�>���Ƭ`���ӾQ�þ����(F>K�o?�$�?�K?f�V�t���S>�ri?Pu=?Y��?��?m�?����pg?l�>���>e�?C�L?�C4?�?��>��>��ڼWƅ;�w���<��m�ҽ�8� �(����=�/>��=��=�M=�ب�?�<�=KgI��%̽\&p=��=�g >�=@��>�[?�l�>�P�>e	<?�U5�v�4�Ll��k�2?��C=]�Z���{�����
Ͼd�B>�ed?�g�?k�O?�P>SD�U�5�@]>vU�>6�>�N`>�2�><�kLB���=�� >͡>O��=[Im���b��\�}㉾��<ŀ>��>�Ǟ>�܈�_�$>t<������hI>.�4���	/��j�F�9<3�����~��>��G?	�*?	=���e�)�� ^���&?�B?��?q��?^�#>����fL�:�-�����'�>a�2>�j��<����f��}����KjO>���%����	b>}��큪���d�j�\���j.u�<E�1�>�D���J4���f��=Z�=ۇ��? ��䑿����P?�{>���F�۽�T꾝@>�Z�>Dr>�>�v��;.���@���D�>j�F>���*C���@�D���*��>{C?�<]?ك??y�J�m�&�H�<��q����Nh�7?�m�>��?:�<>r��=ܬ������a�`{D�n �>]U�>�6���@�&Ҥ����$�:�m>��>�[>�?�Q?_X?An`?��)??̄�>l�ս*�ž�T"?�O�?�̂=�x��PB�W4���H��}�>��?��'�Mҗ>�?��?�R&?K.O?�?��=$���_�@����>�ې>��W�:[����3>q�J?� �>
\Q?��?e� >O<�x)��=2����=A(>5#?e�?��?�%�>P{�>�}�;0�>8s�>�[?�#�?[m>?�/F>CT?<BU>ӣ�>l~ʽ�׽>�t�<��?��i?���?�WB?�]?��#��ϩ�!���q��%�3�:��<�*�aؒ9�N�9��T=���<��H�=F.�=�0�=�(���O���=�a�>e�s>���9�0>U�ľxM��'�@>����R��޼��G�:����=�r�>�?f��>e#�]��=���>0�>���h/(?m�??��+;t�b�N�ھ&�K���>m�A?���=��l��x��]�u���g=z�m?�u^?rcW��$��B�b?��]?�5���<�z�þx�b�-�龸�O?u�
?r�G���>�?�	r?��>�*f��n�����4b��j��ȶ=��>wD�h�d���>�7?��>�Gb>b��=��۾�w��P���*?�?���?���?�3*>`�n�4��$��+D���\[?c�>vԣ��?XW�T˾���������߾n����������<6���� �����ѽЁ�=��?�t?^p?��_?� �=�c��c[��]��.?W�[ ����XpB� >��&C���q�t��bV��8����=8{� y-�]�?��'?�R���>�T���l��I��/>�䆾���=��=����O_<U���֗F������H?qк>�	�>�@<?��W��D@�� .��,D��
�.��>���>##�>ǉ�>Փ�a�z�Pem�����{$��.�4�B@v>/wc?1�K?��n?s[�x$1�߈����!�o�/�e����B>n�>q҉>ٙW�%��_0&��V>���r�����v����	���~=�2?K �>u��>rL�?��?}	��p���dx���1�"σ<�.�>�i?�;�>]�>��Ͻ�� ����>�l?�Q�>�
�>�/��h�!�bFt�sNƽ���>7T�>fo�>�f>� 0��S\��ؐ��q��!t=��b�=Ej??��\�1�>qP?�y;�z�<ko�>��c�
J"�U�D\0��+�=b�?�=�U*>fƾp�H�v�Û~���'?��	?:T���1�D0x>Z�?�q�>���>f�?�r�>�Q��'Z��B ?�[?=|E?��=?�n�>JZ=� ��m����/��+�=`��>�J>��J=���=��.�A'Y�8�Eݶ=	�=ߘ;���2��<�1+�{��<k"�<�7>�Nտ0)F���������V��|B��EŽ�d��z�����辨�̾ v���,R�n<���]����]�;�A�-��?���?�bٽ�U��Ҋ��Jw�<�پ�N�=���4��=����C�����������~$`���e����w�8�'?F����Wǿyg��=ܾ��?�� ?�Oy?�X��;"�t�8�D}>�L�<2���;�쾼���mϿyΚ��%_?ת�>���g��m��>N��>��X>�t>K���[���u�<�_?�,?v�> fr�2�ɿ�U��á�<��?f�@�bE?�u:���ݾ�d	>��?�~?f\>�D�e����ľ��>�$�?���?���<��_�c��=��e?i��=�$�F�j����=�o�:,)�=���>�l>.��>�L��+����^�B6`>s��>�#ɹl���|`��B�=�2�>�}�����5Մ?+{\��f���/��T��U>��T?+�>S:�=��,?W7H�`}Ͽ�\��*a?�0�?���?%�(?7ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�܅�=�6�j���{���&V���=_��>Y�>��,�ߋ���O��I��P��=*T�"�ȿ7( ��v&��.s���m�����V���t��~
��~N��@*M����=���=�dt>��>V��>�Ӏ>TS^?�v?B��>��p>a ��v���N���H2�,��|���8Z��vmC��h������x	�G����4�~��HҾ
�9�{��=�%Q�����Fk��b���F��(/?��>�¾D
L��L�:4CϾ�*��A�;��޺��оZ�0��=n�蘞?<`@?ߝ�� IV�U��.��Xq��U?F彜#�
G��h$�=��>�y�<�z�>�!�=��ھp�.���P�co"? w�>r����ž�>�:ؽm=AN3?���>��>Uv�>~^�> %���멽��v>��/>�a�>���> -�=�x���{½��1?�Ks?C���E���(4>
Z���)����W�e*^>мW���>`���@=g�Z����D����:��!W? ��>��)���]W��s���?=V�x?Ho?X$�>�Sk?��B?)8�<�w����S��$�ݕt=<�W?i3i?Ͼ>�H���Ͼ.b���5?�e?=oO>Dh�)��ĺ.��U���?h�n?1I?P���Bk}�_������}6?��v?��^�� ��x���Q��Ш>,��>���>;8�*԰>�+>?��#��Д�w����4����?�O@�<�?�o\<i+%��2�=�?L��>eM�5hž9N���߶�شs=���>"<��>�v�k� ���+���8?U��?��>$��T� �G>U����%�?(�?$Z���c>�+&�K}Z�Wu���=c6i> �@>ˌ >�q���}C�z����ݾ#�!�^U�=q�>�^@s��@˺>�Λ���ٿ� տ����cN�j�]#?�|�>���=�B��'.P���O�J!i��~��E���פ>�q>���	T�<C���#lM�p�_=c7>*B �e?3>����m.��F���yO=̘>�H[=�>��꾦L�/�?�e���˿�?���tZ���s?��?���?�md?l����M�����⽾�f?L�?��D?w5�����v�5=�wj?T����^�P�3���D�O�P>�4?6��>@<.�H�=Y>��>��>��/�(ſ����M� �[L�?~��?���{��>Yf�?c�*?~>�v����ȫ���*��8H @?��/>�*� �I�=��j����	?�t/?�o����]�_?*�a�N�p���-���ƽ�ۡ>��0��e\�#N�����Xe����@y����?N^�?i�?ֵ�� #�f6%?�>d����8Ǿ��<���>�(�>*N>`H_���u>����:�
i	>���?�~�?Qj?���� ����U>
�}?��>���?���=l�>�=�谾��3��[#>p��=gA��?��M?�4�>�x�=�9�!�.��UF��)R�����C����>��a?��L?��a>�ֹ���3�t!�B�ν�:1��!�2|?��#)��^߽ �3>��<>��>8JE�eӾ�?kp� �ؿ�i���o'��54?@��>�?����t����;_?�z�>�6�,���%��EB�R��?�G�?4�?��׾5[̼�>i�>)J�>��Խ���ꁇ�S�7>�B?���D��O�o�h�>���?�@�ծ?Li�;?h&����/=r�Z��D�[��=]x2?[��j+e>��>�_�=��i�U���w����>=u�?���?���>b�h?��x�SGM��1�=�7�>��p?�?]�=2�ؾ��*>�&?4��9������/`?Y4@��@y�]?�ɞ��ܿ���'���X�&ِ<d��:�j>�S%��]�<d�=}�=�YF=��7>j��>�m> K>�D|>Y�u>͑H>P��x9$�0P��{����P�!�3� ��â��N��]~�ײ��
_�|_��j���K]=���@q���ڹ�S��=��U?-qR?gIp?�� ?7�s��>���L=��%�EV�=j�>�T3?I�L?��*?�6�=����c�*Z������J���'�>��I>���>/��>_��>]�;;�I>��=>��}>6�=/X=	�D�@=ūL>�>��>��>_�>�2�>;�ſ��4���#���~>T�?�ho�	�}������s �Y��fe�>-�B?z�9����:A�fw����.?+2B�Z4��yΫ���=%1W?�J?�Q�>вI��B����,\ڽ&�����4>x5�=Hc��*ݾ�6>щ$?�l>^��>��G�N)�4�i������>/hm?l���ԃ4�9O���+I�����? ?^a��~;�|=������S:�k��5f?*!>o�l>hk����־z��Sm��?�?�>d[=�ŋ>��=�E,� ��0�����>�<�>�a?Ҟ>��=M/�>$���7�Q����>�3i>O{�=�A?�w ?�I��ֽ�&���K<�\�>&�>��>Y��=�7���S�=Q�>(K�>P6�=(!����0���f>����gw��-���V�=��%�|b�=u C>��P�l�*��� <�~?���(䈿��e���lD?S+?` �=0�F<��"�E ���H��G�?r�@m�?��	�ߢV�@�?�@�?��O��=}�>	׫>�ξ�L��?��Ž5Ǣ�Ȕ	�*)#�jS�?��?��/�Zʋ�=l�6>�^%?��Ӿ_w�>N>�TG�������u�4#=	��>�#H?�i���O��)>�<^
?v ?t����L�ȿ��v�0��>��?�?�m�/:����?���>*��?�Y?Зi>m^۾08Z�Cb�>�@?�R?S�>�?��6'��?[ն?v��?b%L>\$�?�xs?RP�>��j�N.�Ɂ���Ό�_R�=WL;�o�>AR
>�ݺ���E�;˓�������j����1b>��%=.Ĺ>T+޽Lk��6+�=m�����s�����>��h>m�L>��>"�?���>�t�>�m!=v���}��kך���J?���?���$�g��_x�2��=O�!�d?t-5?�ɣ�������>�NQ?�	�?��_?DU_>q��Q��K��.C���Ա�PXW>9�?lE�>�
�x3*>��ݾ�tF�-�>���>�9��/�о�Kn��I�����>�S?(q�>C���� ?wY#?5�q>�Z�>^C�o��0�F�z��>0�>�?��{?��?铹��_6��z��A����M^���M>v�x?��?���>�$��K@��>�ںz���פ�/'�?e�g?�/�k�?,��?xr>?ίB?Djm>�F��vϾBU��fOy>�� ?Rνf�G���M����\�>l�>�H?�Eٽ�{�=ŽԒ�a�5��?�J?�3�>�2ܾ	Y2��	�����<[�ν>��p�;��%<�c/>*;>i���	cO>��6>�Z>Li?������-M<���+�>#�U>K�$����<S<,?��G�yۃ����=��r�ivD�k�>�NL>J ���^?f=���{�����w���U� �?˞�?4j�?w	����h��"=?��?B
?j#�>�J��$}޾���bPw���x��v�X�>���>�l���b���ۘ��F��eƽj/ݽN ?E��>ض?��>t�>��>zo���F.�T۾_��BE`��a��=��C�բ��׾�#��ނ=���5�w�"��>p�5�)ι>� ?(Xy>�Ob>�Ȱ>/�����a>�G>*��>�Ȋ>_>iB>td�=Sd=�֏�k9R?k����0(�È�ힲ��(B?�d?ۂ�>�b�8������>�?$�?��??Yx>^�h�{�*�8�?��>�*��/�	?�M>=�~Ļ���<����l��9퉽:��u�>Ƥҽ��:��L�ce�n�	?�5?������ʾ���?'�=��V?��?�e�3ai�zGH�t�J��3m���&>3�@������j��J�b�R���ۀ�L���S$�#�ͽ�8F?���?� ��ͭ�����P�V��e���ހ<��=��>�5`>�0�>'$���*M�D�<��Ί��>XF?�M�>RU?��\?��:?{F?f'�>lqP>-ٶ���?�~����>u�>��7?.�?!�F?��3?�'?��>HFf��ʾw�ľ���>N�?��/?(�?�'?�Jڽ�+�Gv�;S��K��8k�a�μ|u� �G�p�μ��o>�9�>lo?���ߗ1�޵�>W^>��-?�C�>��>�w��}�m�_�;��>��?c�>���tns�g�����>�ބ?Z"�]>�<<�5>���=��G��?���\�=\�ټga�=����k�.v%��E�=	�==�B��K�w�b�j����<.0=�s�>&�?���>=F�>=��X� �l��g�=kY>�S>F>�Eپ�|���$���g�ay>w�?�y�?g�f=B�=��=�{��eT��@��b���n��<z�?I#?�WT?ꔒ?��=?pj#?R�>+�6M��|^��z����?�$?օ�>�!�l&f��S����4���:?	�?l�@�<��a=X�ie�`�<���w>0�
�q�������L�\�����Q��٘��T�?X1�?1i�>o�q���fk����澤�L?�m�>	,B>�>�>|;�U]H��"���\��j9? ?i��>�L?��s?��f?���>15پ| Ŀa���O���� 4�	l?j͟?��?�u?fYy>��>;Ƚ8�����4@���_=��Y���=���=U_ >"��>6Fw>M����I�ΰĽ�N��&;��>�%?�@�>2�>l�s>�u�Q�G?m��>X����!���!���T/��w?ln�?�5-?�t=�v��H�
����>��?"�?� *?�BP�r`�=�m��V���n��׶>'ĸ>��>xq�=)�c=1o>��>ӱ�>8	����
�8��)��?��C?lh�=2Hſq��.n�,����ny<߹���Bg��œ��v[�Oy�=����|��Ψ���\��Ҡ��+��"$�������{��&�>3�=��=��=�H�<�缛W�<1?=�/s<#�=�c����<�X1�=�ûR�K���-<;�A=~�%H˾�}?YAI?ok+?��C?�jz>D>�2�X��>_���O?��V>R�L������P;�5E���Δ�TؾP׾Nd��ʟ�)T>��J�)�>/�2>ɀ�=A#�<���=k�u=�=��_��=���=F��=�-�=m��=��>�&>�6w?X�������4Q��Z罥�:?�8�>c{�=��ƾp@?�>>�2������yb��-?���?�T�?>�?>ti��d�>L���㎽�q�=J����=2>s��=w�2�S��>��J>���K��F����4�?��@��??�ዿТϿ8a/>�Q>�G&>Ic>���a���P��ϕ��բ�@�M?��]�,�=��F'>Q���G-��?W���@>=8�����t���OQ����=
W���h�Y�h�dK�>�G�>JL>Q	H���@>�z=�g=J>অ�����pƽ��t=-�Q>��>�i>b3�>O�?B?ǖa?N�>P��<��_̾��>�R�ش?y,>q�>��e>��8?�S?�EW?��>��=Yp�>��>���ׄ�O�Y�оE�A��p�?z?���>K7����X[���4��Y���k ?�h2?e�>��>�%����m-���l����}���;��3¾����dZ��ץ�C�뼧�>���>ױ�>�V ?⤹>y�>{��>��=�==��=����\o�AY���_>7�=2�<���0/��kK��V�=�,/�A��<JE�P�=�[
=u��=<[�>�t>���>qE�=�峾.%->G���C��=����(�C�*w_�r�}��"��W�/0+>��_>ye��������>E�k>�V?>w��?)�j?p�>3���`Ǿ"e��ёx��m;�wе=(@*>�_���2�>Z�l�Q��IѾ�	�>���>5��>��q>��W�@�7�'>��վ��B����>�dƾ�#(��������=���(�����}�<�fZ?Ǚc��7���r?��)?eى?���>M�߾i���k�>+��(�>ږо�hW�d��p�/?�&?��>���k	Q��-v�W��>ڇ��^#��@|�148��pѽ˴�^9�>����5־u�Š���Ô���A���ľ�	�>"gH?N��?U�������� ��V����N>�?4�]?K��>q=�>C�?�?7<�����¯;� >.Ř?�n�?
�?9!�<}�>W�ܾ�B�>�~+?���?�?o??c����+?	g6�Xv�=�4N����=�[l�,F��̹>?�.?PD(?�k7�,��g��b-ھ�����0_=���=-�c>#�u>^|>��=��=��׼E�>���>���=nU>�3�>s��>�ѥ����&?���=H�>A2?�;�>��[=ө�j��<�J��.?�-+�P$���>⽶/�<璻��P=�R̼ٶ�>gǿp��?OU>�F���?���1��mS>��T>�,ܽ=�>��F>�f}>{�>��>�>��>�k'>>)���Z>����P�P-9���V������d>����_�U��%�b��ξ[{#���j�X-��R�7���=���?Hb���T���w���?��?��/?:۴��4�[�u<��>�\>E澰�=ވ�X�R�?���?<c>v�>'�W?�?�1�x3��uZ��u�2(A�e�!�`�{፿����	�
����_?��x?*yA?�T�<�9z>2��?��%�[ӏ��)�>�/�';�@<=�+�>*��L�`�b�Ӿ��þ�7��HF>o�o?/%�?cY?
TV�֞A<���>�K?t'?�{?N+J?��?z����4?��	<R+?ޥ?t
@?�>`�?��>u�;>[/>1�=6��hw��3O��d���iM���3=5&�=M�=���=�Z
>�n�<�j漩څ��]E�&r��)�<M�>C��=��='�>:1[?�C? ��>;�5?7���*��A��2�:?3(=��3����ᛎ�������(>�r?0?�?0�S?��u><)���3��[!>��{>Y�*>�u>�2�>H߉�gD�z}=cF�=�=YΝ=eo���������˧��{�;b�>�5�>{�z>������'>�R��)�|�ɂc>eH��A����X���F���1�Bw��B�>��J?Kv?:��=�a�8����>e���&?o�<?�@M?mT?Q�=��ܾ!�9�K�@����>��<Y��/���&���9�������n>�����_���=�t/����]�wuo�T��K���(���c>��"���������7�>�T�>��<��?�&q���+��H�F?�{�=��׾�Ͼ��p�N>�C�>�?��q={5��9O�`�ɾ����|�?�>�����ۇ�G�'������>�nC?la[?q?�?ѿ}�x�v��@�j����R������HU?N�>#"?�nI>Cƺ=�`�����&d��4H��m�>o��>�Y��5H���������%�Nԓ>���>�m4>j�?l�I?؂
?�~`?��)?V� ?�ӆ>�Q��YƬ�p@#?��~?���<Ҝ"��D���0� s5���?CV?�'��Y>�l�>���>��:?�IQ?C��>Ŷ>����(27���>�Ĕ>�_J�~ձ��5>x�]?��>?YH?�q�?$�>�;!�H`Y���1��R�=Hm�=�@0?��.?�?5V�>|x�>u�R���B>%��>�D�?��?1M?�	�=��D?G>~F�>�S =��?J��>2\?�n?�}?�Zb?Z&�> =Ì8��nt�������S���=��=��h>�S�=`����н9_��h�����@=�!�<7C��C"��"�P��m@��&�>K t>���k�0>�ľ0e%A>����� ��Wߊ�&n:����=��>s�?<Õ>f�#��x�=<�>�q�>���s(?�?H�??�;f}b���ھ��J�
�>��A?�A�=z�l�+����u�T-d=�m?�]?pU�����нa?��^?���Y?���ƾ+:L�վ�SL?#?�^F�;�>�8}?OUj?���>�6d��;j�Xu��tpa�شR�=�=U �>F���de�;�>5�:?!}�>�_>���=��ܾR�y����٦?ʍ?x+�?���?��*>ϖr�f)ؿ�@���Ώ�BR[?aI�>�w����?��4;�c���׉���پ0����{���ۢ�AJ��.�������΢�ƅ�=,�?��r?t�j?��]?�[�	]�0	V���~��U��������^�<�*�C�*�C���l��.@��zj��rF=����v�@��?�C)?Y,A�%e�>���� ��[�^3�>�^��#V���t=6�X�=T�����~��@��ڛ�k�'?d1�>�6�>��??�qY�w[=��,.��n5�����\>�|�>���>��>��B��"Ž�jv�y>Ǿ`���f�)��>v>N\c?�aK?�n?/� �}j1�&f���g!��3�iݧ�ΘB>I>IΉ>eW�݆��%&��t>�7�r�����s�� �	�Q��=�`2?S�>�*�>��?�??s�	��Ԯ��x�ź1����<�>=�h?a��>6��>!yν� �ķ�>ۿl?>��>n �>�c���O!���{��˽��>���>���>T�o>/z,�n+\��u���w��Y9����=�h?�W���K`���>��Q?�J:gF< 7�>�x��!�����'���>��?��=-t;>�pžt$���{�6R���J"?w*?߶��`>��fs>?]b�>���>�W{?{n�>5���h�=�a�>��U?��D?�p6?���>,��=����]ɽ�?�
�/�ȁ�>�L	>�9�� :'=<g��a1���뽔y�=��=t}�=����[�=s̼�ݳ;8U�Nd`>�Oֿ˖G�V��e�۾�����*�}�5�f��	¾��<������ž<q��������������5��]}��&r����?wf�?;޿��?s�롚��q���ڌ#>Vd��5&�=rܔ��{@=�6���r����S��E��{����^� �'?䥑�߷ǿ����y8ܾ�" ?9J ?�y?��x�"�m�8�`� >x��<�?����������ο[���E�^?n��>G� (��@��>0��>f�X>Nfq>���ݞ�.ה<��?��-?���>v~r�ؓɿe����`�<P��?h�@��9?�m>��¥��ڵ=X�?��?J��=z6����ߘQ�f9�>���?�u�?=*���D��_�<�Ia?��=x,%�i�<#��=G~�=9�G=|e�:�'>y�>��ɽ����=|	�x�=�i>��ν����vq��
�K����=�\+�ˠ��*Մ?{\��f���/��T���T>��T?C+�>�:�=��,?17H�G}Ͽ��\��*a?�0�?ۦ�?1�(? ۿ��ؚ>��ܾ��M?bD6?��>�d&�!�t���=�8Ἆ�������&V�3��=Y��>ل>��,�ً�H�O��M��8��=1���Vǿ$>���/�%?��LǼ��=����.=�i�;�|���Ȟ�4����ü�N�=���>��]>�[Q>��>XQ?�l?�m�>���=�Yǽ�����6Ҿ�q��p��m��ľ��F}�����Q�ƾ�
�a��c�=����I:���=�
P����r �m�`�sB��F-?�>~Ⱦ�$M�`J<�]˾5����`�������о?e0�|�j�*��?�B?�r���W�v���]֪�aRV?Ձ�ov�	���>���X�&=�;�>��=:B�D�6���Q�4n?���>p��>׾��=3 ���2<��D?��?j��=,h�>�� ?6X���3��q�>JN9>Z�>�{�>&�G>{����l���?�]?�S��)Ѿn�>�yݾ(�b�����뗦="虾#��=$0=wI�<o�T��2~��9 �(��dV?䣐>�M(�TD�򐾵� ��p=&�v?��?��>Ͼf?݂B?m<�*����Q��
��|D=,nT?�2i?�&>�yg�B8Ҿ�9��˨1?��e?��X>�~f��A侾�-����f1?�k?2X?9U����z�������	��M7?��v?s^�vs�����>�V�g=�>�[�>���>��9��k�>�>?�#��G������xY4�$Þ?��@���?��;<��L��=�;?k\�>�O��>ƾ�z������N�q=�"�>���|ev����R,�b�8?۠�?���>�������">�̛�)��?A��?�:�mU�=JE)���C�FR��,iQ��c>b�+>+M]=��!��E^�d�����;��Y<��=?�>�@����a��>W�����ɿ̱������ॾU�޾f_�>���=�,��Z���s���@��Z���侘��>�K>�cp�t���̓�`�3�nQ=~�Y>f>���ă>6����<6�ɘ˾OX�=�.�>�
->��b>����� ��K�?�-����ƿsE��>�)���o?Y�?�1�?a�Q?<]��+��R|��@�����g?�B?��r?k�=w*ƾ��;��h?�`����U�u92��>C��_l>D?���>X4�|�<n�=��?"��=7�*�ptÿ������Q�?���?���<-�>���?�5?a@�B!���J¾1�+�w	�D�C?�@>>�ʾ�F�ӂK�=$����?A�?� ǽR�'�[�_?(�a�M�p���-�|�ƽ�ۡ> �0��e\�gN�����Xe����@y����?L^�?f�?۵�� #�b6%?�>`����8Ǿ{�<���>�(�>�)N>H_���u>����:��h	>���?�~�?Rj?���� ����U>�}?P�>��?D��=�U�>��=��-W(��^#>��=�@���?d�M?K�>-d�=��8�m/�N\F��=R�  �F�C���>��a?ipL?G�b>� ��R�2��� �B+ν�1����ئ@�ģ+�l�߽�4>)�=>;`>J[D���Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Oz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>D�Խ����\�����7>1�B?Y��D��u�o�y�>���?
�@�ծ?ji��	?���P��Xa~����7�m��=��7?�0��z>���>��=�nv�ܻ��U�s����>�B�?�{�?��>�l?��o�Q�B�{�1=8M�>˜k?�s?cRo���n�B>��?������L��f?
�
@~u@_�^?'6.��9���B��|#����<9c=J�2>��>��̂=]˽�y ���F��{�=�'>a�2>���>�\d>��|>�3a>i��y*%���ڿ��I�J����,B�4�v�mWO���������\ɢ���Ծ�
����<P$�<n���R5���w����=M�U?�Q?��o?�� ?��z�+�>�p���=
�#�j��=�ۆ>�S2?\�L?�*?V�=�ĝ�V�d�;V���C��Ӳ��ؼ�>/&I>���>�>�>�;�>�b�8q�I>�
?>Vw�>�� >�&&=���C�	=��N>��>t�>���>[JD>V;>󌴿���`k��p�"�����?����kL�����(������/3�=
4-?^%�=7���kп�׮���E?
������&E����=r1?��T?�0>���{�f��u>�d�yq����=aB���Vi�u�"�%9M>��?gu�>�y'>�Q����a�s��bx����>�eZ?��.�<ٟ��Є�|a�����&�>G
?�ƃ�r ��m ��4��=(M�Yh�=m�8?S-�>�7��xʗ��j��#T���(->܉>qP>C�>��>w�����}��Wf����=I�q>�5~>�u ?`	(>�am=�A�>����jT����>�MQ>�,>��8?Y~#?��M��Я��^�����Fx>�Q�>�|�>l�>�;�.[�=���>k�b>��-�V�������E��<>�$?��Dd�|FW�	�f=������=gB-=>���Z?�O,i=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾRk�>n`�?W�������u���#=n��>�5H?�S��Q�O��>��w
?�?9a򾿦���ȿ.~v�%��>$�?c��?p�m��@��r@�t�>��?2jY??ki>^Z۾�eZ��z�>��@?�R?�$�>05�Q�'��?׶?ʯ�?�s�>�<�?K֊?���>D��=�u���������=�?�<���>5�V>2�aSA�����2Dh��J���Ⱦo�>���=S�>R�ܼ{�Ƹ{=6���3Ѿ�;a�pҝ>�h�>��h>sfa>��?d��>�e�>�9'>��������g��V�K?q��?����1n�]K�<Y��=�^�K)?�E4?79[���Ͼ�˨>k�\?�À?�[?_X�>_��=���濿�z���ܖ<�K>�&�>C�>�򈽹PK>��Ծ�%D��k�>ї>u���4FھD-���6��XB�>�g!?+��>��=��?��$?}�l>ݩ�>'=�v���f�*����>�h�>ґ?�zg?Y�?�m���<�1@���隿��e�ͅ<>l�u?wf%?C��>HŌ�s�$����=�ԣ�!x?@�Z?*ֽ���>�K�?��8?�IA?�8h>t\%��rо�=q��o>6� ?^FZ��A��/��tt�t�?�?�&?���<)���W�f������ ?3�L?���>��侪�b���;�/H=(�<A,���$��B⾼�J�>���>R $<�8>h��=��=�9۽v1f��e��.v=�8�>��P>���2�=�<,?�G�i݃�C�=��r��wD��>�NL>� ���^?�i=��{����w��� U�@ �?l��?�j�?G��i�h��$=?�?S
?� �>�L��W{޾���nQw�2�x��w���>��>>�l�&�j���-���TF��9ƽ�I�l[�>s�>q��>��?�,>IW�>��|��e1����Y���V�<�ξN��?�8�>�������n����<X̾���OS�>�����><�#?��>��]>�h�>�������>�mI>�P>���>���=���=�>'av=��㽪8R?f7���'����d���3B?e�d?��>@�h�us������?�B�?	K�?<�u>EYh��F+�2
?��>���b
?x�9=�)��u�<IB��W@��Ɔ�*��;��>�Dؽ=�9���L��e��-
?�?�咼�G̾�<Խ�`��$L_=���?տ&?�'�4�Q��h�-�V��PT��̮�md�����}x$�Os�z،��`��j=��̔$�1[=bz-?��?5 �df辤t����e�͘;��+[>,�>��>TԱ>�e>�<�d/�{&X�E�-��O��H��>�~r?x�>�#L?wxC?�E[?�"T?^$�>�6>�y۾kq?�R�=���>� �>��H?�?o1?Q�!?��9?��>m㧽|��IҾki ?y"?�!?�?,�?��"�t-�<�~T=�]�f�JTp�P� =h��<���E<��
>�WP>cl!?���<�f*�3�p >�aI?	�'?���>?�6�;����	�ك?�N�>���>����nS��'�?L�>�>�? )ż�X�<X�>T�H>�k��`Z�'+>JQѽw��=��z�
8j�Od�<��<��`=�B+�qs&=�r��7T.=�k�='�>�q?�-�>I��>���ܘ ���9�=.�S>�I>��>S�ݾ5����2��te�Ģw>�Ջ?س?���=.M>�=	ʚ�V��7y	��c��#�=�?E�?�U?�ߍ?V??�k?K�=����!�������Ө��?�%?�ܦ>:������[���'���(?�>�>U�3��-Z���*�Z�Q�ӏ�Sg=�q#�k3W�0n��E�@��`��i���,���?�Г?kb�>)�g���*��K��Z���]?[�>�E>�Z/?q�5���P��J⾓�»��
?H�!?�l�>8�\?�d�?xY]?I(�>y,�����	���r>>t��>�c?�t?:��?�]??��a>�c>5���Ar�C���������l_���K�='�H>6�>$ ?K�o>�Q>`쑽%���T�� >�FU>�6?N�>��?�G�>�ʸ=MvB?؎�>��ƾ�"�~!���q>�̬�:B��?Y8�?�?�q&<��
��'V�h�Ӿ���>��?r�?�
'?э=�Q��=��B�BþH���I0�>  �>~��>�˜=�l=��>0��>!w�>�龽V#��L<�2s�=�%?�F?�P�=�Mƿ��q���n������8<1Z���&a�Eb����]��I�=�����\ �<^��/�c�-{������v���n���\/n�h��>5	�=�>G�=1C�<8����<֝C=Ƣ;<!�,=�����R�<3(,������B�>/Y<��D=�� ��˾2�}?�<I?�+?��C?�y>A.>��3�~��>�}���A?�V>?�P�R���q�;������ ��+�ؾ�v׾$�c�&ɟ��D>�\I���>	93>tE�=6,�<��=�"s=�ǎ=؊Q�E-=h&�=�\�=�m�=��=��>�Y>�6w?R�������4Q�pZ罡�:?�8�>�{�=w�ƾv@?��>>�2������jb��-?~��?�T�??�?ti��d�>V���㎽�q�=�����=2>��=r�2�R��>��J>����J������~4�?��@��??�ዿɢϿ_a/>��E>�+>�hH��>��P#���@����x2?��"��2��=R>�F=A�;����ԝ=-k>"��=yK��G�A��	�=�����K<%���a�>H.m>�J�=�c��n��=���=f�5>���>O�Z�j`�����j�='�>ͷ�>��>i�>m�?`�0?أc?���>x|f�ڇѾ�\��G�>nW�=	۲>)R�=fF>�O�>6?��C?�hL?�c�>�l�=��>$H�>B+���j����Ң�p~�<�,�?Fǆ?�X�>�<��@�Ut �0B>�~P½f�?��0?��	?�>����d� '���c�za�3J��S=�3J��X~��]h�(�%�	cA��<�=k�_>���>���>�F>qh<>�"�>X��>�>L	�Re����ؽx�ȼ��)<|GC=��м�=�0ۼ��=D��=�Hj;SO=���<�������tw�S��=U��>�=>��>���=$"���C/>✖���L����=���1)B�ld�j:~���.�6��=B>?X>�2��B,����?�OZ>�h?>�|�?.u?�>&��վ�M����d�^{S��=��>_>=��g;�:C`��M�gnҾ���>x�>���>i�n>a�
�S�D��)>X�޾HC���?5�u�H����=f���zj��^�u�iΆ���$�&68?�
�����0�?�C8?�>�?���>o\���8��hH�@�Y���>����={/�=s�>o	?c
?S�j�w>��H̾���޷>:>I�P�O�l��0����Ϸ�F��>	�����о.$3��g�����؍B�Qr���>еO?t�?a6b��W��TO�?��i&���p?Z{g?��>@K?!??���y��q��0w�=|�n?���?�;�?h >L�=%cƽ��>`r�>��?�b�?_*J?��)�@>�>m#f<���>G����]>�">8>/�$�I>��?z?u9?�臽���پ�����Z�\��=#���ob�>fh�><��>��>��>�-=
 >�Җ>�>��>Ip�>g��>B��q����=?%�6>�!�>\4?�f�=-�<$�N��س=���>D�=;"]=~�K�9���>�HF>[C>�=^w�>F�¿D�?>t>v��_F�>���T��<7I>�ڤ>��ݽ?ce>*��=�G�>s��>�F&>���>���>�$Ѿ�<>�Y�����^@���R�m�̾��y>�Y���'���.% ��L�
������o=h���RW:�)�<uh�?=�yh��)��%��5?��>7�4?Iː�H`^���>]��>�q�>���PҔ� ����Y��g�?��?d;c>��>!�W?�?H�1��3��uZ��u�>(A�e��`��፿������
�$���_?��x?2yA?�V�<::z>:��?��%�gӏ��)�>�/��&;�0?<=�*�>�)��W�`��Ӿúþ�8��GF>#�o?%�?jY?�RV���a�[ +>�2;?Q1?+Eu?�E3?Yb:?x5���%?�v4>�z?(?S�6?�.?��
?�9>��=�.�:��3=�/�������ٽ�׽y	��-E=��=���;h<<��=鰌<#���!���%<*3��/�<�~4=���="��=̩�>QM[?��>ɺ�>e�<?�.>9��C���3;?�ƥ=�Q��В�A���M�����=�xl?E��?9�]?�k>O�B��&J�2>���>P�F>n�g>��>#�����>�=�>�B>T��;��{��B��R�����8�|=o�->C#�>��f>T��h�M>>���x��;ޏ>G�����n�������$�BZ+���u����>�3J?j�?j��;][��5V� T���?/<d?��4?A��?)�ݽ[E����?�AfJ�?���K�>*�9`Ͼ�����ț�&o�z}��s�>�轓y���n�=�A��j��	�y��qM��yɾ� P=�I���*����A���n�y>�>y�ž���w���b��3�O?��
>����Yh�U��q"[>�q�>�>0�=�dȽ�5W�@���I�>=���>�`>΍ǼT�׾ǬO�C���W��>�HE?��^?>�?�7�� 5s��A�O��J�~5���)?�d�>�3?�(B>h)�=]������Td�UPF�=4�>ɢ�>�@���F�(���*N�0�#����>{?�,>�i?L^R?*?�2a?�J+?T?���>WýgI���� ?�]x?ڗC:_�u|1�y�&��|?j0?=�ܽ'�E>u^?��?�H5?�Y?�&?�k>�T���F��=�>P�}>zzX������m>�)]?�c�>	~X?�߆?�0�=p�9������Ge�|�=d>��6?ܤ-?Ed?�i�>u�:?ιV��l{>��?[؊?���?��.?�{�=}�;?�q�>Ũ'?)M�=��? 3�>?��q?���?�w[?�>�F�ק���^%���l����0�=v�>��2�fO�=��>V|��`���n=��=�L�x:e�6s�<b�=4]�>b�r>���>,>3Ⱦ�T���UF>��q�03��ʏ�HjD�=�=�z>.�?C��>N	&����=-ݶ>���>D~�j�(?]�?�/?��>xd��$޾	P�.h�>p�A?�h�=_#m��Փ�C6t�Y{=Կm?�i\?F�^�ں��&�b?��]?�h�9=���þ8�b�&�龄�O?H�
?��G�I�>>�~?��q?W��>E�e��9n����Db�G�j�^Ӷ=r�>�W��d�A@�>+�7?�N�>L�b>�+�=�u۾��w��q���?O�?u�?k��?�,*>N�n��3��C��D���T[?&��>�_4�M�?��[��ޫ�qv�������ƾ!ržx���v�ž�t���f��Ix�*�c�G�=U�?��n?E�f?�fW?J�վ��V�TST�&���&0@�1����q��p>�\�m�qJS�z3����?۾�>���_�=z���
B�3T�?��%?h(�-+�>뙾ɓ�a�̾N�F>y霾��N��=밚��<=�`=Z:g�}+'�?���N ?���>�H�>�G<?K�Z��Z<�E�0�Ie6��v��N9>5��>&�>���>!h����+�p���ʾ�<����ƽv6v>�yc?I�K?=�n?�[��)1�����Y�!���/�bV����B>�>o��>��W���9&�(P>���r�0��_o����	��~=@�2?�#�>���>�J�?�?H{	�zP���Yx�3~1����<^@�>� i?�>�>���>~*н�� ����>i�l?�5�>H��>���� ��z�<˽|
�>ܭ>��>�fn>9*.�Ȁ\��`��+ڎ���9��l�=�li?�ǃ�t�`�p��>0R?ޭع��*<���>��|��c!��8�(���
>O�?*��=M�;>��žq�,�z��ى�=�!?�?
\���dJ��2>��?v��>�K�>�t?ѧ�>*�žH�ٽVo�>�l?N�F?}E?��>�Χ=[MW�
���ª�E(�=A��>름>�;�D᪽��� 7���a��=o�=�v�;��M��=@�0�e���3=ܞ>�ֿ�}Y��)��ϑ��t(�[��&w��hf�筇�R�)�6K����D�u��$�"�UU���m�´��$�����?�,�?c@S�m'�s-����`�4GϾpn�>I#�r���S�뾘hs�㨑��m̾$�>�6��w?��k�Q�K��]&?�]��Y0¿���J���(?�S%?�t?����g%���>�zL>�$w;�m���־�љ��'ǿ`�����`?��>�پ��*��ܰ>%�>�̌>*�>�Ql�q��A��<J;�>�/+?��?�H��ÿ����a==��?:t@��A?y�'����[��=�P�>�%
?V�9>��6��j�1ﯾVU�>Z�?޽�?��L=JCV�׼@f?s�j<n�E���R����=�ߤ=�	=V-�<�I>�g�>n��DD��ڽ(�5>��>o ���4�]�e��<%;Z>�Խψ��ӄ?"s\��f�C�/��R��T>G�T?j:�>F�=ҵ,?B5H��{Ͽ��\�m-a?�-�?���?�(?ҿ��ƚ>��ܾ��M?�C6?�>]]&�#�t�;K�=&nἚ줻 ��� V�\��=s��>+�>g,�8���O�.`�����=OL��(�ܿm�]�����@T�8P�d��b���x�|�n皾bb���9���=U�`=Ï�>�]6>iZ=�=R�<?b`�?���>X�>�r�C4����޾����\���@��mLq�u�?$>��[�i���)�
��.���&�V�;�==։S��E����*�r_��?�I�+?�*>�ھ�P��X�8�Ⱦ����5�;1�ʽ*�̾WF;�:Ql�|h�?<D?����K�X����!:�;�v�o}\?� ½_�
�WȾ�,>M���=�>6Q�=��߾�6���;���$?:0?��¾����,��=2��tP;��K?$��>�	>��q>��>1���!�=p�>y�3>�K�>?|�>z3������c�ɽuc?��p?��\��l���?>��¾iʂ�DD����=�e4����=E��=��>���wW��"��'K<�cP?�S�>���l�q
x�	H��+q�=��l?��>\�>�#h?��(?��E����^�T�q@�[s�uT?�f{?2�(>;�Z�!�ݾX`�� ?.?S�f?�R>tKI��c۾09)�U��/�?��i?��?C�<�\�������b׾[??��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������3��=ߕ�[�?O�?�~��Բg<����l��m���נ< Ϋ=P�<@"����h�7���ƾ�
��������s��>�Y@�L�R/�>�A8�;5�pSϿK���Yо+Wq�W�?1y�>d�Ƚ������j��Ou�t�G���H�H�����>3>N���#e��z5~��UM���>��>B(���>Wϐ��n㾧�R�� �=�)�>�:�>DE>�_���پ���?�@꾝�¿�S��r� �ҝ`?��?e�|?_C?J;
>R����˽�(Z��S?���?�/�?���=�䖾�
�S�`?#3�-�5�[q ��|�k��=��.?�֦>7�f�?��=��9>���>�}%=��m�N���ȿ�.K��3�?���?l�¾�U�>7��?�Y?�����;I����%���=��?��g>��.��N־��Z��mB�}C	?�?��ؽV�Z�_?%�a�L�p���-���ƽ�ۡ>��0��e\��M������Xe����@y����?K^�?g�?õ�� #�^6%?�>_����8Ǿb�<���>�(�>�)N>�H_���u>����:�i	>���?�~�?Sj?���������U>�}?P$�>��?�m�=�a�>�a�=���,�#l#>y#�=r�>���?_�M?�K�>�X�=��8��/�[F��GR�m$�R�C�N�>M�a?�L?\Kb>��-#2��!��xͽ0c1��I�7X@�M�,�|�߽�(5>�=>5>��D��Ӿ��?Jp�7�ؿ j��p'��54?1��>�?����t�����;_?Lz�>�6� ,���%���B�`��?�G�?=�?��׾�R̼�>8�>�I�>O�Խ����[�����7>/�B?O��D��w�o�y�>���?	�@�ծ?hi��	?���P��Sa~����7�P��=��7?�0��z>���>��=�nv�ݻ��^�s����>�B�?�{�?��>�l?��o�N�B�d�1=8M�>Μk?�s?<Mo���t�B>��?������L��f?	�
@~u@_�^?)���T���vT�I�����<`�@>��U>ʰ���DJ>2*1><"�=��`=K��=Y"k>�k>ʵ�>W;>4=o>7Ă>�z��(��:пቿ�.e��2������g�U�U�S��+��6¾����k)/���7�{�������F��$EB�T��=��U?�R?=p?� ?��x�T�>w����=�#����=O*�>'h2?r�L?٠*?KƓ=�����d�#`��N@���Ƈ����>�pI>}�>�F�>�'�>�DX9P�I>�9?>���>�� >�v'=M�躒:=-�N>�K�>���>T}�>Q->F�=����>��x6~���Q�dq\����?�At���[�HЗ�I�\�Y����J�=�2?��="����#Կ���+O?�9K��$�*����L�=�oE?|�e?2�J>���կ��e�Y=�P9=��`����=���Dz�Q��xMJ>	y1?|w�=,;�>u32��.��A^��qھ��>��-?���L˾�����+I��������>���># ��8� �-]��ex����>c!?��?)��=�,�[�������\��՗>2u>��Ze>�M	�r�J��.���ʽ��2>?�2>�?�,><X�=ڡ>�(��#�P�\�>�H>�,>�B@?�$?So$��ؠ�����(���v>��>>$�><�>��K���=���>Ʉf>ٲ��1������A�;�T>SS���^��t�ӑ�=H�����=��=k��ɑ?��#=N�~?�}��J㈿��疶�QqD?.?��=@G<��"���~<����?��@�j�?a�	���V�2�?Y@�?���Թ�=��>yΫ>�	ξ5�L�W�?'�Ž���"�	�15#��O�?�?��/�pɋ�
l�>=>�b%?i�Ӿ~��>V!�A��0̆�w�s�9�0=���>YG?M��ߊC�1L9�"?� ?P�������ȿ��w����>�?�}�?�?k�����?����>9�?�-Y?&�k>}�پCcZ��?�>�>?r�Q?��>���"1��?���?�	�?{�F>�[�?'~�?��>��\�1�z������|J�=��<��>ZNT>�"��q�>��̓�ᓃ�R}N�D�	�>l8>�Ur=nX�>�޽fI���pE=�O�ꧦ�Ψ���>�>Q�>M8�>Ƒ?T?�4�>��9=KJ=�f���\��1�K?���?F���2n��$�<��=d$^��5?@D4?�)^��о���>��\?�À?�[?�|�>=���A���߿�iq����<��K>��>�;�>�Ո�%�J>��Ծr"D��5�>֗>�H����ھi@��Q0��S�>�e!?Є�>mi�=��?Op$?`dj>qɮ>ЉC�:z��H�B��c�>���>�X?�{~?)�?f��o4�����ԡ�� ]���N>�%z?�?�G�>�����蜿���M�#����Ga�?��d?9��j�?��?�4??�A?��e>��t�ܾ�矽Z�>��?�8�h�C�d�5��-@��.
?�q?
?j,�{���.{ѽ�������?aeU?+ 1?�^�9^�ZHؾ�,=�<]���7��u�<gg:>P��=���ͬ�=1l�=���=��z��e��g�ۻ�W=ġ�>އ>�ۢ����;,?.jG��ۃ�`Ԙ=3�r�NwD��>�eL>,�����^?ir=���{�Q��*s����T�7��?1��?�h�?�1��,�h�"=?��?�?�"�>�I���w޾,��YXw�"�x��u��>���>A�m����.��������F���ƽ��u��(�>�X�>=�>�=�>y��=�=�>a
������F��ؾ8V=���	��*��1Z�_I�Oȟ���_�89��/�����>��
���>\??�>௃>��>�ӣ=	��>
2�>���>w<�>}�S>�kr>�ҕ>��{=�Y,�iP?'���A&��������Y?{?
�?��=$w��H9�H$?S_�?��?�\n>>�f�m�����>���>�;��	9?�:�<�>R5	���F��n��+Fl�ڄ^>��X�ΙI���:�OO�|�	?~?�e�<3G��g@���i�� >�s?ɜ?�W���J���N��pQ��O��ʽ��E�$ξ��?��1y�����m�@:d�� 
��V#��T/?�t?�V�����q�b�f��(���$>a��>H��>,��>��>���s*�\�^�9H��B¾6��>���?�i�>�F?{;?L�U?L�N?�ݒ>�8�>Z����Z�>ZI�;Ԧ>�,�>h>?U�+?m�.?�?b�-?~�r>���$��/�Ӿ��?T�?ZC?\�?$�?T߁�[��)���#	?�H�l���n�"d{=���<�7˽EP[���]=��R>�?"?��}�'���/a(=�T?7 ?�A�>p��\���S*�B�>�2�>1B�>~���1?��*z�Jŧ>�&�?b�=��=Xv(>(=Z=���=P�<��>����>�� ��.^����;3H>���= %�zOý$�i<SE>V���/s�>��?�>.B�>�?��l� �N��Fc�=�Y>S>�>CFپ~���$����g�FYy>�v�?Rz�?�f=�#�=���=Q}���U��O��������<-�?HH#?XT?X��?��=?j#?D�>l*��M��`_�����g�?��+?�>��ԯʾ�T�� 3�+�?�?�b�F�C�(�ҕ¾0�׽�	>KL/�J� @��K�B�I�:)Z�V���}(�?U?�D�=07�*���u��U�����B?b��>�	�>��>L�*��g�S���8>q��>~CQ?��>\�7?\�?�J�?���>����ƿd��?�=ف�>ٸi?3�?���?3�N?9j�>l>"��=����]~˾/�=��}�<>�}�m>e�t>`d�>��>,~�>�Y�>�7ٽ
n&���z��&�>.��>���>���>��>}j�>c	=�t:?Jj�>����4�u����ʽ���=)�?���?��?sjѽ��5�
1a�ۤ�9��>(��?9i�?�(�>,?���.�=�I�<���Rʬ��>?l�>�A>/f>S\=_�=>-�
?y��>�R��� ���/�.���]?�p?��@=��ÿ`u��mw�I�<D(���li��@����j�
�=E���� �ݎ��uFN�=8������}!��( ���߅�2��>��=`�>7>>��X���ф<��=7�*�Fu=ҍ{�� 	��^�'�����>�����Oy���*<Yڧ�2�˾��}?�;I?ݕ+?��C?�y>+;>Ք3�G��>�����@?cV>�P�������;�L���� ��R�ؾ x׾��c�ʟ��H>�`I��>�83>�G�= L�<%�=#s=�=��Q��=$�=�O�=�g�=��=��>NU>�6w?U�������4Q��Z罤�:?�8�>�{�=��ƾs@?w�>>�2������sb��-?���?�T�?>�?Nti��d�>I��w㎽�q�=8����=2>?��=v�2�R��>��J>���K��6����4�?��@��??�ዿ̢Ͽ0a/>�*7>�#
>ЂR�3�5��d�N�U���C� �%?W7��þ�y>�v�==�辧��H-=q�F>a��=tg���\��(�=d�Z��6`=�H=L5�>x�7>�J�=/����=��=z>~yT>�Y���e����N=�N�=��v>+f>ER?Ў?}+?ᛈ?G
?Ѯ|������$��>��=���>�p>j?;��>�&?��S?�~]?5#�>�R�=�B�> Ƣ>��f�j�����$?
��R>	�?
�l?��>ڒ�a��.�#�y1"��{����>)!?Ff�>���>�)����P'��F.�.���a���]�!=��r��hX��
�}��Lܽ0��=�֪>k��>���>T)w>|l5>�AI>6��>�>U��<_�=tV��7ޫ<����*z=!Φ���<��� ����L�<%�%3��[�Z�:�;i�<f�:Ų�=mQ�>K	>���>���=ߓ��0�.>�Ҕ��lL��S�=X_����B�ӊc�|}���,��4�a+B>��U>�8��0��t�?�Z>�@>ƈ�?�t?�j >�D��]־������a��T���=wr�=mE��Z:�:`�M���о̋�>���>$P�>�s�>���l��νK���O���>�xѽ�І=Ғ6�v͒����A�g����@>�?l?�u���$ּ(�?��?|�?�t�>b������D?��޾ws�=�O����.�&Q�>��&>^�U?TgL?�x�Q d�ؒ̾!X��Ty�>#I��O�(���?�0��C.�����U��>U���о��2�O��88��nB��kr�/>�>�O?y��?1gc�%��/UO��v����8y?�Lg?�>�7?�e?������쾐���r�=G�n?|��?i�?`�	>Md�=?���o��>/�
?�B�?eՏ?�`k?�J�ޙ�>��w�ޣ5>��;�ц>g�>��f=[��=��?�(?O 	?���o
�A^�������U�u�.=�Ѵ=-�>�9�>tk}>2��==�r=�(�=m�Q>Mץ>v��>H'k>���>g��>18�F�RM?�Y= ��>8�?⿯=¬p<�����<:H�=?!>*1	�Y�nK��&|�;.��<��o>[�<���>��¿�t?~�>����i.?Zd߾ =�>�g=���>	"��ƙz>��>���=�K?
s�>���=��>7�>�����^>���3���a3�V�<�սa�8�I>��澩��v߾���๻���U�
���i�@q����,���$>�V�?�os;#�N��)�j����?�?a�6?y
ɾ��=>�V>���>���>�ľ��v�̸��c4'�({?)��?�:c>��>-�W?	�?h�1�3��uZ��u�i(A�>e�?�`��፿����
����"�_?��x?yA?�O�<�9z>F��?��%�`ӏ��)�>�/�';��;<=P+�>*����`�?�Ӿ�þ�8��GF>^�o?0%�?�Y?�SV�Bc���&>�:?A�2?��t?�E2?�H:?��M�%?H�2>G�?��?�/6?lG.?�
?(�5>���=���sL'=!���q:��S�ϽZ�ɽ������1=�7�=����.e�;��=~L�<
YѼ�cϼ#D;�����<��9=(آ=ml�=?�>�VO?E�>@��>9�E?�u��4/?��%ɾ��??�U=$�)�/nE�H&�&辳n>t?�d�?`?EO>�!�\�"��#>�؅>3>�SB>v�>6X���	d�ďt=�7>܆>�>�=�t��:z�9��:K��/�<A,>��>$��>.۽nx�=��@���OU>$s�� ��νs���?�C�K��j���>&r?�{?�ħ=���7P���Ku���'?�%?D�H?�z�?	�x=�}��)�|���\��"ɾ��>M]������������V��6�,�o1>�j��_���=�t/����]�wuo�T��K���(���c>��"���������7�>�T�>��<��?�&q���+��H�F?�{�=��׾�Ͼ��p�N>�C�>�?��q={5��9O�`�ɾ����|�?�>�����ۇ�G�'������>�nC?la[?q?�?ѿ}�x�v��@�j����R������HU?N�>#"?�nI>Cƺ=�`�����&d��4H��m�>o��>�Y��5H���������%�Nԓ>���>�m4>j�?l�I?؂
?�~`?��)?V� ?�ӆ>�Q��YƬ�p@#?��~?���<Ҝ"��D���0� s5���?CV?�'��Y>�l�>���>��:?�IQ?C��>Ŷ>����(27���>�Ĕ>�_J�~ձ��5>x�]?��>?YH?�q�?$�>�;!�H`Y���1��R�=Hm�=�@0?��.?�?5V�>|x�>u�R���B>%��>�D�?��?1M?�	�=��D?G>~F�>�S =��?J��>2\?�n?�}?�Zb?Z&�> =Ì8��nt�������S���=��=��h>�S�=`����н9_��h�����@=�!�<7C��C"��"�P��m@��&�>K t>���k�0>�ľ0e%A>����� ��Wߊ�&n:����=��>s�?<Õ>f�#��x�=<�>�q�>���s(?�?H�??�;f}b���ھ��J�
�>��A?�A�=z�l�+����u�T-d=�m?�]?pU�����нa?��^?���Y?���ƾ+:L�վ�SL?#?�^F�;�>�8}?OUj?���>�6d��;j�Xu��tpa�شR�=�=U �>F���de�;�>5�:?!}�>�_>���=��ܾR�y����٦?ʍ?x+�?���?��*>ϖr�f)ؿ�@���Ώ�BR[?aI�>�w����?��4;�c���׉���پ0����{���ۢ�AJ��.�������΢�ƅ�=,�?��r?t�j?��]?�[�	]�0	V���~��U��������^�<�*�C�*�C���l��.@��zj��rF=����v�@��?�C)?Y,A�%e�>���� ��[�^3�>�^��#V���t=6�X�=T�����~��@��ڛ�k�'?d1�>�6�>��??�qY�w[=��,.��n5�����\>�|�>���>��>��B��"Ž�jv�y>Ǿ`���f�)��>v>N\c?�aK?�n?/� �}j1�&f���g!��3�iݧ�ΘB>I>IΉ>eW�݆��%&��t>�7�r�����s�� �	�Q��=�`2?S�>�*�>��?�??s�	��Ԯ��x�ź1����<�>=�h?a��>6��>!yν� �ķ�>ۿl?>��>n �>�c���O!���{��˽��>���>���>T�o>/z,�n+\��u���w��Y9����=�h?�W���K`���>��Q?�J:gF< 7�>�x��!�����'���>��?��=-t;>�pžt$���{�6R���J"?w*?߶��`>��fs>?]b�>���>�W{?{n�>5���h�=�a�>��U?��D?�p6?���>,��=����]ɽ�?�
�/�ȁ�>�L	>�9�� :'=<g��a1���뽔y�=��=t}�=����[�=s̼�ݳ;8U�Nd`>�Oֿ˖G�V��e�۾�����*�}�5�f��	¾��<������ž<q��������������5��]}��&r����?wf�?;޿��?s�롚��q���ڌ#>Vd��5&�=rܔ��{@=�6���r����S��E��{����^� �'?䥑�߷ǿ����y8ܾ�" ?9J ?�y?��x�"�m�8�`� >x��<�?����������ο[���E�^?n��>G� (��@��>0��>f�X>Nfq>���ݞ�.ה<��?��-?���>v~r�ؓɿe����`�<P��?h�@��9?�m>��¥��ڵ=X�?��?J��=z6����ߘQ�f9�>���?�u�?=*���D��_�<�Ia?��=x,%�i�<#��=G~�=9�G=|e�:�'>y�>��ɽ����=|	�x�=�i>��ν����vq��
�K����=�\+�ˠ��*Մ?{\��f���/��T���T>��T?C+�>�:�=��,?17H�G}Ͽ��\��*a?�0�?ۦ�?1�(? ۿ��ؚ>��ܾ��M?bD6?��>�d&�!�t���=�8Ἆ�������&V�3��=Y��>ل>��,�ً�H�O��M��8��=1���Vǿ$>���/�%?��LǼ��=����.=�i�;�|���Ȟ�4����ü�N�=���>��]>�[Q>��>XQ?�l?�m�>���=�Yǽ�����6Ҿ�q��p��m��ľ��F}�����Q�ƾ�
�a��c�=����I:���=�
P����r �m�`�sB��F-?�>~Ⱦ�$M�`J<�]˾5����`�������о?e0�|�j�*��?�B?�r���W�v���]֪�aRV?Ձ�ov�	���>���X�&=�;�>��=:B�D�6���Q�4n?���>p��>׾��=3 ���2<��D?��?j��=,h�>�� ?6X���3��q�>JN9>Z�>�{�>&�G>{����l���?�]?�S��)Ѿn�>�yݾ(�b�����뗦="虾#��=$0=wI�<o�T��2~��9 �(��dV?䣐>�M(�TD�򐾵� ��p=&�v?��?��>Ͼf?݂B?m<�*����Q��
��|D=,nT?�2i?�&>�yg�B8Ҿ�9��˨1?��e?��X>�~f��A侾�-����f1?�k?2X?9U����z�������	��M7?��v?s^�vs�����>�V�g=�>�[�>���>��9��k�>�>?�#��G������xY4�$Þ?��@���?��;<��L��=�;?k\�>�O��>ƾ�z������N�q=�"�>���|ev����R,�b�8?۠�?���>�������">�̛�)��?A��?�:�mU�=JE)���C�FR��,iQ��c>b�+>+M]=��!��E^�d�����;��Y<��=?�>�@����a��>W�����ɿ̱������ॾU�޾f_�>���=�,��Z���s���@��Z���侘��>�K>�cp�t���̓�`�3�nQ=~�Y>f>���ă>6����<6�ɘ˾OX�=�.�>�
->��b>����� ��K�?�-����ƿsE��>�)���o?Y�?�1�?a�Q?<]��+��R|��@�����g?�B?��r?k�=w*ƾ��;��h?�`����U�u92��>C��_l>D?���>X4�|�<n�=��?"��=7�*�ptÿ������Q�?���?���<-�>���?�5?a@�B!���J¾1�+�w	�D�C?�@>>�ʾ�F�ӂK�=$����?A�?� ǽR�'�[�_?(�a�M�p���-�|�ƽ�ۡ> �0��e\�gN�����Xe����@y����?L^�?f�?۵�� #�b6%?�>`����8Ǿ{�<���>�(�>�)N>H_���u>����:��h	>���?�~�?Rj?���� ����U>�}?P�>��?D��=�U�>��=��-W(��^#>��=�@���?d�M?K�>-d�=��8�m/�N\F��=R�  �F�C���>��a?ipL?G�b>� ��R�2��� �B+ν�1����ئ@�ģ+�l�߽�4>)�=>;`>J[D���Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Oz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>D�Խ����\�����7>1�B?Y��D��u�o�y�>���?
�@�ծ?ji��	?���P��Xa~����7�m��=��7?�0��z>���>��=�nv�ܻ��U�s����>�B�?�{�?��>�l?��o�Q�B�{�1=8M�>˜k?�s?cRo���n�B>��?������L��f?
�
@~u@_�^?'6.��9���B��|#����<9c=J�2>��>��̂=]˽�y ���F��{�=�'>a�2>���>�\d>��|>�3a>i��y*%���ڿ��I�J����,B�4�v�mWO���������\ɢ���Ծ�
����<P$�<n���R5���w����=M�U?�Q?��o?�� ?��z�+�>�p���=
�#�j��=�ۆ>�S2?\�L?�*?V�=�ĝ�V�d�;V���C��Ӳ��ؼ�>/&I>���>�>�>�;�>�b�8q�I>�
?>Vw�>�� >�&&=���C�	=��N>��>t�>���>[JD>V;>󌴿���`k��p�"�����?����kL�����(������/3�=
4-?^%�=7���kп�׮���E?
������&E����=r1?��T?�0>���{�f��u>�d�yq����=aB���Vi�u�"�%9M>��?gu�>�y'>�Q����a�s��bx����>�eZ?��.�<ٟ��Є�|a�����&�>G
?�ƃ�r ��m ��4��=(M�Yh�=m�8?S-�>�7��xʗ��j��#T���(->܉>qP>C�>��>w�����}��Wf����=I�q>�5~>�u ?`	(>�am=�A�>����jT����>�MQ>�,>��8?Y~#?��M��Я��^�����Fx>�Q�>�|�>l�>�;�.[�=���>k�b>��-�V�������E��<>�$?��Dd�|FW�	�f=������=gB-=>���Z?�O,i=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾRk�>n`�?W�������u���#=n��>�5H?�S��Q�O��>��w
?�?9a򾿦���ȿ.~v�%��>$�?c��?p�m��@��r@�t�>��?2jY??ki>^Z۾�eZ��z�>��@?�R?�$�>05�Q�'��?׶?ʯ�?�s�>�<�?K֊?���>D��=�u���������=�?�<���>5�V>2�aSA�����2Dh��J���Ⱦo�>���=S�>R�ܼ{�Ƹ{=6���3Ѿ�;a�pҝ>�h�>��h>sfa>��?d��>�e�>�9'>��������g��V�K?q��?����1n�]K�<Y��=�^�K)?�E4?79[���Ͼ�˨>k�\?�À?�[?_X�>_��=���濿�z���ܖ<�K>�&�>C�>�򈽹PK>��Ծ�%D��k�>ї>u���4FھD-���6��XB�>�g!?+��>��=��?��$?}�l>ݩ�>'=�v���f�*����>�h�>ґ?�zg?Y�?�m���<�1@���隿��e�ͅ<>l�u?wf%?C��>HŌ�s�$����=�ԣ�!x?@�Z?*ֽ���>�K�?��8?�IA?�8h>t\%��rо�=q��o>6� ?^FZ��A��/��tt�t�?�?�&?���<)���W�f������ ?3�L?���>��侪�b���;�/H=(�<A,���$��B⾼�J�>���>R $<�8>h��=��=�9۽v1f��e��.v=�8�>��P>���2�=�<,?�G�i݃�C�=��r��wD��>�NL>� ���^?�i=��{����w��� U�@ �?l��?�j�?G��i�h��$=?�?S
?� �>�L��W{޾���nQw�2�x��w���>��>>�l�&�j���-���TF��9ƽ�I�l[�>s�>q��>��?�,>IW�>��|��e1����Y���V�<�ξN��?�8�>�������n����<X̾���OS�>�����><�#?��>��]>�h�>�������>�mI>�P>���>���=���=�>'av=��㽪8R?f7���'����d���3B?e�d?��>@�h�us������?�B�?	K�?<�u>EYh��F+�2
?��>���b
?x�9=�)��u�<IB��W@��Ɔ�*��;��>�Dؽ=�9���L��e��-
?�?�咼�G̾�<Խ�`��$L_=���?տ&?�'�4�Q��h�-�V��PT��̮�md�����}x$�Os�z،��`��j=��̔$�1[=bz-?��?5 �df辤t����e�͘;��+[>,�>��>TԱ>�e>�<�d/�{&X�E�-��O��H��>�~r?x�>�#L?wxC?�E[?�"T?^$�>�6>�y۾kq?�R�=���>� �>��H?�?o1?Q�!?��9?��>m㧽|��IҾki ?y"?�!?�?,�?��"�t-�<�~T=�]�f�JTp�P� =h��<���E<��
>�WP>cl!?���<�f*�3�p >�aI?	�'?���>?�6�;����	�ك?�N�>���>����nS��'�?L�>�>�? )ż�X�<X�>T�H>�k��`Z�'+>JQѽw��=��z�
8j�Od�<��<��`=�B+�qs&=�r��7T.=�k�='�>�q?�-�>I��>���ܘ ���9�=.�S>�I>��>S�ݾ5����2��te�Ģw>�Ջ?س?���=.M>�=	ʚ�V��7y	��c��#�=�?E�?�U?�ߍ?V??�k?K�=����!�������Ө��?�%?�ܦ>:������[���'���(?�>�>U�3��-Z���*�Z�Q�ӏ�Sg=�q#�k3W�0n��E�@��`��i���,���?�Г?kb�>)�g���*��K��Z���]?[�>�E>�Z/?q�5���P��J⾓�»��
?H�!?�l�>8�\?�d�?xY]?I(�>y,�����	���r>>t��>�c?�t?:��?�]??��a>�c>5���Ar�C���������l_���K�='�H>6�>$ ?K�o>�Q>`쑽%���T�� >�FU>�6?N�>��?�G�>�ʸ=MvB?؎�>��ƾ�"�~!���q>�̬�:B��?Y8�?�?�q&<��
��'V�h�Ӿ���>��?r�?�
'?э=�Q��=��B�BþH���I0�>  �>~��>�˜=�l=��>0��>!w�>�龽V#��L<�2s�=�%?�F?�P�=�Mƿ��q���n������8<1Z���&a�Eb����]��I�=�����\ �<^��/�c�-{������v���n���\/n�h��>5	�=�>G�=1C�<8����<֝C=Ƣ;<!�,=�����R�<3(,������B�>/Y<��D=�� ��˾2�}?�<I?�+?��C?�y>A.>��3�~��>�}���A?�V>?�P�R���q�;������ ��+�ؾ�v׾$�c�&ɟ��D>�\I���>	93>tE�=6,�<��=�"s=�ǎ=؊Q�E-=h&�=�\�=�m�=��=��>�Y>�6w?R�������4Q�pZ罡�:?�8�>�{�=w�ƾv@?��>>�2������jb��-?~��?�T�??�?ti��d�>V���㎽�q�=�����=2>��=r�2�R��>��J>����J������~4�?��@��??�ዿɢϿ_a/>��E>�+>�hH��>��P#���@����x2?��"��2��=R>�F=A�;����ԝ=-k>"��=yK��G�A��	�=�����K<%���a�>H.m>�J�=�c��n��=���=f�5>���>O�Z�j`�����j�='�>ͷ�>��>i�>m�?`�0?أc?���>x|f�ڇѾ�\��G�>nW�=	۲>)R�=fF>�O�>6?��C?�hL?�c�>�l�=��>$H�>B+���j����Ң�p~�<�,�?Fǆ?�X�>�<��@�Ut �0B>�~P½f�?��0?��	?�>����d� '���c�za�3J��S=�3J��X~��]h�(�%�	cA��<�=k�_>���>���>�F>qh<>�"�>X��>�>L	�Re����ؽx�ȼ��)<|GC=��м�=�0ۼ��=D��=�Hj;SO=���<�������tw�S��=U��>�=>��>���=$"���C/>✖���L����=���1)B�ld�j:~���.�6��=B>?X>�2��B,����?�OZ>�h?>�|�?.u?�>&��վ�M����d�^{S��=��>_>=��g;�:C`��M�gnҾ���>x�>���>i�n>a�
�S�D��)>X�޾HC���?5�u�H����=f���zj��^�u�iΆ���$�&68?�
�����0�?�C8?�>�?���>o\���8��hH�@�Y���>����={/�=s�>o	?c
?S�j�w>��H̾���޷>:>I�P�O�l��0����Ϸ�F��>	�����о.$3��g�����؍B�Qr���>еO?t�?a6b��W��TO�?��i&���p?Z{g?��>@K?!??���y��q��0w�=|�n?���?�;�?h >L�=%cƽ��>`r�>��?�b�?_*J?��)�@>�>m#f<���>G����]>�">8>/�$�I>��?z?u9?�臽���پ�����Z�\��=#���ob�>fh�><��>��>��>�-=
 >�Җ>�>��>Ip�>g��>B��q����=?%�6>�!�>\4?�f�=-�<$�N��س=���>D�=;"]=~�K�9���>�HF>[C>�=^w�>F�¿D�?>t>v��_F�>���T��<7I>�ڤ>��ݽ?ce>*��=�G�>s��>�F&>���>���>�$Ѿ�<>�Y�����^@���R�m�̾��y>�Y���'���.% ��L�
������o=h���RW:�)�<uh�?=�yh��)��%��5?��>7�4?Iː�H`^���>]��>�q�>���PҔ� ����Y��g�?��?d;c>��>!�W?�?H�1��3��uZ��u�>(A�e��`��፿������
�$���_?��x?2yA?�V�<::z>:��?��%�gӏ��)�>�/��&;�0?<=�*�>�)��W�`��Ӿúþ�8��GF>#�o?%�?jY?�RV���a�[ +>�2;?Q1?+Eu?�E3?Yb:?x5���%?�v4>�z?(?S�6?�.?��
?�9>��=�.�:��3=�/�������ٽ�׽y	��-E=��=���;h<<��=鰌<#���!���%<*3��/�<�~4=���="��=̩�>QM[?��>ɺ�>e�<?�.>9��C���3;?�ƥ=�Q��В�A���M�����=�xl?E��?9�]?�k>O�B��&J�2>���>P�F>n�g>��>#�����>�=�>�B>T��;��{��B��R�����8�|=o�->C#�>��f>T��h�M>>���x��;ޏ>G�����n�������$�BZ+���u����>�3J?j�?j��;][��5V� T���?/<d?��4?A��?)�ݽ[E����?�AfJ�?���K�>*�9`Ͼ�����ț�&o�z}��s�>�� ue����>!��ʾG7e�~�l���Ѿ
�=LVB��4=M ��b��<���%=���>\_$�h N��\��椧�{E?PW>%���X����ʷ�Dh�>OY�>K?���=2�H�yQ�9��� s=�I�>�+>
ڎ>%�~�h]��~�3��>@?y�b?Ao�?��Y���f���\��D��E���C�=R�(?gZ�>��!?f�4>�=����Xw��:R�S}3����>���>��%VE�㙝�����5��&>�s�>��u>tT?jh?�2 ?��e?��D?��?m,z>>�;�q�Ǿ[w%?�e�?��=���x�[~4���@����>@)?�V��j�>h?A?� +?��Q?��?ʮ>���J+D�?�>�ˎ>�U��Ȱ���g>�M?_��>��^?��?{�->��1��F���ݛ���=4&>�D9?}b%?��?T��>��>U��=��>��>�GF?Ar?� V?c[�>bO?�4>L
?\>h>b?�>��u>b>��C?,+�?\�x?��R?�g=7�'��=���=@��=��=�4�<�>�>��=�!����g���ǽ���=�L��k[�i2�q^-=zj��I�>A�u>�敾��0>�%ľ�D��jB>5⢼ǣ��u1���9�_ư=YO>?�r�>*c%��O�=�E�>"�>����&?��?53?�+�;�b�$پ��J�㨯>kNA?�f�=1�k�z��l]v��I\=�Kn?/�]?E:W����+�b?e�]?�f��=���þ��b�׆��O?�
?K�G��>��~?��q?|��>��e��8n����(Db�6�j�ն=�s�>X���d��<�>N�7?�P�>&�b>+(�=v۾_�w��p���?�?��?���?�'*>��n��3࿔:��|P����]?���>4
��6�"?��;�Ͼ����	*��E#��N���F��yi��n���~$��ƃ��Qֽ%K�=?�As?Oq?�_?r� �jd�Y�]�����V���5�M�E�^E�ԇC��o��n�ܚ��jg����F=PԀ�0@�G1�?��#?s5���>�O����D&о�J>�]��F�|�=�}����,=�N=ey�#v,�uΩ�U ?�O�>-B�>�=?~�Z�x�<���0���5�����%6>�r�>]�>���>�\�;���qa���ƾ������Z>-b?��5?in?gCѽq�C��͇��b&�����B���y+>���=a�7>���G]ǽ�VH�w1L��5_����B��� ����3>��?�]>:�->��?L�	?Y�*�}���6����D��;�=��>\�T?�a�>��$>���� ����>o�l?��>Z$�>����G!�n�{��4˽�>��>u��>Wp>�,�B\��_�������9�D��=X�h?䀄���`��ʅ> �Q?��:E�I<+��>*�u�A�!�����'�<�>c�?���=\�;>�|žW-���{��4��j()?Y�?f_�� �)�|O{>?� ?�}�>�G�>"Ѓ?,��>.þ�+��p�?�_?{�J?�p??4��>�P=䵽ɽ�'�G?=�H�>Х[>k=���=���)�[��h�Y�J=za�=��¼�6��$)	<�e����:<o� =�6>�(޿�>��pǾ$�#�\��#��J4��*��Ӿ���_ھ𖺾����މ����G�`�Ma���l��=����?���?Ik��
�������9醿�ԾId�>@���˼J��V.��E�R���پ&��O)���r���_��<[�U�'?������ǿ𰡿�:ܾ�  ?�A ?��y?����"���8�0� >�=�<�8����^�����ο������^?:��>b�.�����>i��>O�X>4Gq>���`螾�<�<��?C�-?x��>�r���ɿ)����Ϥ<���?�@��??%�#�Y���cQH����>�8?̀u>�<"��:��j;���>1 �?��z?�L� g��>�cO?�Y	�*�-��0(����=a:=>���=���D�>��>ï�&Y���='j�>�>5��=^��<Pg7�G��=�-�>���=��&>5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=s6�񉤻{���&V�}��=[��>c�>,������O��I��U��=2�
��ɿ�w+��L&��`=5 6�nLl�,�	 �����X|��B ���s)�����>y�o>�1[>��L>��t>_�P?�$m?�l�>@��=�<�L���}3���꽃˻�~�<�������9�֠�r�پ2��`)���,�S�Ul農�7��_�=A�J�|����G�f�j���0�o�>"���Ⴞ�L��t��ƾ|e˾���<���1���|�M�e�|&�?p�3?t^��B�.�Ӌ2�.Y�����c=?�T@=�.�+(¾S�+>�z���6>���>n�J�S*��H&8�-��.U/?b�?0���i���k,>���A*=�(?�-�>���<p/�>@�?F*8�R����x>n
>"�>���>���=�h��<޽bt!?�R?<��1���Dߕ>����c]�]��=4�)>z�!���@;_NY>�> =+�{��M%�����`=H'U?��>[�$����:$��T�C��aJ=!�p?��?_��>��k?��E?���<�!��W�Q�,����{=�W?oj?��>˴���G۾$����<7?�yi?V�[>+X��2��<5�����V?�on?|�?࠺�{��l���:���3?N�v?Bq^�;q��w��z�V�Q>�>�^�>���>��9�]b�>#�>?.�"�~E��Z���EV4�o?m�@���?�<<S����=�<?T[�>m�O�+>ƾ�y��*y��
�q=��>���hv����R,���8?���?5��>����0���N->�����?zƌ?0��]|�=I��]�Z�����>MdP>���<DF�=*5��5�v��R���;[�]F�=~A�>O@l�����>�S��Z�忩1⿋���̾jX.�>�E?آG?]]K>�ɾ�qG��Q�@�[���Y��b��T2�>* >4�ܽX̔�����e:��V��1�>�μ>fb>L�u�߷����[IL=��>���>6Sf>����ھg'�?k
վ�=ȿ󣚿����\?u�?��?��)?�l�Z���⃾>�#�0K?0e?E]?�*'<�j��D��!�j?�_��jU`��4�nHE��U>�"3?�B�>G�-�"�|=�>���>g>�#/�y�Ŀ�ٶ�*���X��?��?�o���>q��?ws+?�i�8���[����*��+��<A?�2>���G�!�A0=�OҒ���
?V~0?�z�R.�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?"�>(�?�-�=h�>�P�=x��!B.��U#>s��=�h>�Y�?�M?�.�>��=��8�V-/�ZF��;R�'�Y�C�O�>N�a?7nL?�Wb>b\��;~1�V !���ͽ�C1��	�@^@��,�f�߽C 5>��=>��>��D�J�Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?kQo���i�B>��?"������L��f?�
@u@a�^?*�׿�ɕ�N^�VI��|@�=�(<I��=烽Aa�=S��J�&��JT���=�L>��H>#vl>���>���>�Ɖ> b��'%�Yu��Ʉ��79�wZ+�G�7�f6�ã��˨��$%�q�xû�ZV)�@Տ;��D=gg�f{���=��	>�X?[[>?��j?#��>@;�G*>�O꾙,:=�ɽ��J=)B6>�"?��S?�s:?u��坾�!W��|�N������ֈ�>�0
>���>���>V�>��b���6>�
>>��>S�>v��=�]O�x� =�у>�s�>��>���>�0{>]��>�ٴ�|x��A;������)U�fs�?����@c�����8鳾P��LY�>��3?�+�<ǻ`�j�ؿWȰ�?z6?m�"���
��už�o6>?O>?�E>?��>K.���1��P�=�vR��u\�z��IF\�e�(=1�ݾ��h=4�?5a�>BS�>�FN��L���N�xXѾ�HY>�@G?a������W|��X��2�� >(_�>�f�������֌�3:u�r����=��?Y.?��;�e������D� �{�>�`�>��>��!>�@Q>�W>6u�=RS���w�H#�>�|�>�?:>�X�=ʙ>\ˌ��}W��|�>��J>��S>vy6?�\?�F��刽�?M����bo>���>H �>��>�J�N?@= ?�#H>ί�'���5��������T>dH��M-��#���H=T��)��=���=��;���Y�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ-h�>Ux��Z�������u�ö#=O��>�8H?�V��V�O��>��v
?�?�^�ީ����ȿB|v����>M�?���?[�m��A���@�{��>,��?zgY?ioi>�g۾�_Z��>һ@?�R?�>�9���'�w�?�޶?ѯ�?=`I>#w�?ϡs?d��>�	v�A=/�,Y������	�=��;��>�e>S���X5F��ɓ�/<��Ǟj�{�� b>{�$=E�>k+彰U��ؙ�=������Fcl��>��r>�K>�1�>�??���>4��>s�=V4��i���9 ���K?Ư�?����m����<���=��]�^@?+4?�[�y�Ͼ2��>�\?�ƀ?�3[?b{�>���i)���ȿ�H����<؞L>���>7C�>�l��`�K>�jԾraD�v4�>���>|A��n�پ�悾����ڝ>�#!?FD�>��=�� ?Ɯ#?��j>�0�>}YE�5��/�E���>��>�P?7�~?h?y����X3�9��4᡿H�[��BN>�x?oR?�̕>���䁝�IfE��"I�&�����?�kg?�)�a?�4�?��??s�A?�Nf>�z�Eؾ,ݭ���>*�,?�9?��l �c=���6�K$�>��<?E� ?n2=�5���7�����L��ii�>@�$?�i2? ��zdv����C=� �=7�8�N�.�2Ƴ���5>��>�+����=�!����i�8��2�m���+�>�䄽����x��-=,?d�G�vۃ���=~�r�5xD���>�IL>�����^?]l=��{�����x��)	U�� �?��?[k�?!��7�h��$=?�?P	?Z"�>�J���}޾-�྘Pw��}x��w�;�>���>أl���J���ܙ���F��,�Ž_����>I^�>�`?��>�;>'�>�ԑ�$��������pY�����;�[=/�Y;�jC��4�5�]�E�����Lx���>5�k�E�>�#?��U>�s>\��>�~�<�Ӗ>��a>�>sަ>�9N> :E>'2+>�2�<.Ɗ��JR?������'�k��~����(B?�rd?d/�>=�h�҆��t���w?���?!p�?�Av>*xh�%*+��e?0�>���Ko
?#v:=/��o��<3L�����Y��������>�i׽�:��M��wf��d
?�6?V�����̾�D׽&;��7�q=��?�5(?�"*���Q�`4o�h�W�umS�q���Oi�+¡�"�$���p�y��(L��~M��=b(��p)=��*?	�?e������뭾�3k��7?��9f>���>��> 
�>�I>�	��Q1��]�$'��v��G��>��z?Gȇ>�]G?�7?��Z?upM?K��>)�>EtϾ���>�̖�J!�>V�?`�C?H�?' ?�R?�?+�>Z��U�F�۾���>T&?av+?2�?i?c/(�N����{��5��F���~�m:�k�=5�=�� ���\��~�=Z�>EU?�����8��7���j>37?��>2��>6���s������<V�>fb
? ��>����;|r�BD���>fg�?�J��=Ɲ*>�x�=����[f���|�=��ż^|�=l#|�8�7���%<8��=�=�_�r)�9��:���;<�<j��>��?z�>G9�>Xtz�S1�����U_�=�t>�\C>�>]վJ���0Y��4}f�,ix>���?���?#�=j��=O�=y��Se���'
�#���^="�?%�%?�T?k�?sb5?�5#?���=����ϒ��b��o���^0?&�?C��>X(%��a���b���t%�Η>��>�w)����'�'�ϲ����S��>-������c��8�6��G�y-�����z��?�E�?dk�>�4{���$i���!��b?�Q?o��>�?����`8�J�X�S���20?d�;?��>�[(?�[{?i��?xU�>�ɾ˽�ZQ����e���?ȿ�?�"�?hܭ?%��?��>���>�;��	t��gD���ɽN�R���!��'!>�OY>t��>Ү
?6��>�ͽuĀ�֑�k���ƽSj2>W8�>�iq>���>A�~>���:��G?o��>TI�����K����+��d4�o�t?^`�?�P*?Rp=ҵ�tE�����u�>"e�?_��?Xa)?kVS�0��=[Uռ�0��4bo��F�>pR�>vN�>�Ɠ=�L=��>d��>h��>���fh���7���H���?I�F?�&�=4������:�}>��(M�=�@��]8���_��PX�� �=�E��>xE����<�j��c��+��\'��t���y|Z��"?��7=
��=\N�=C������Ԕ=o~f=;־=`A�Eo8<��=�gr�Q��=;\��o�=��(=6!������|˾��}?�6I?��+?��C? z>�C>4�<��>ق�D?LV>Z�O�����i;�䜨�C���ؾmY׾;�c�6џ��)>JMI�2>'T3>�Q�=�Ԉ<��=�{r=ʛ�=�`���=�8�=
��=w�=��=��>�.>�6w?X�������4Q��Z罤�:?�8�>f{�=��ƾp@?�>>�2������yb��-?���?�T�?=�?@ti��d�>L���㎽�q�=P����=2>x��=v�2�T��>��J>���K��C����4�?��@��??�ዿТϿ4a/>\|>�i>��L��>5��x*�&Y��P۽ɿ>??6���Ծ�mk��埽S}󾧁���'K=A�=M�<Q9��}e���=�y��i��|�`=fW~>W�)>�Ș=��`���E>���=���=��u>L���@�=��1<���Gr>�Ds>�ք>���>��(?�P?Yz?4�>��Ƽ������	�q�;>ȼ�>�a?#چ>Xt�>�v>A@?3�6?��B?F�>�y.>�>��>���5p�q��z9I��l'>��Y?��?���>Ȏ����?���0� �e�6�9�H��>�??6��>�\�> ��%�ῗ6�ׇ3���w�}��;�s$��A��3,�q�o�"&;��<��i=a"~>T��>��>�t>�L?>��t>r�>���=r�>�s�<�I��G�6����|<�����䡻��ǽ�($�GK���W<�3�i�����2�p�ɨ`����=;��>JD>���>���=���[/>ļ��j�L���=�2��KB��%d��B~�Z�.�~U6�D�B>�BX>�N��-��վ?��Y>�?>~��?Au?� >���'�վ�R���he��6S���=��>� =��f;��T`���M�cҾf��>���>J�>�l>�+��/?���u=<!�Fd5���>v��ط��l��q��*������i�A�Ѻ�vD?K<���m�=0~?ܗI?�ݏ?�/�>W���nؾ=k/>�	��6=1�o�p�����e�?��&?�W�>����D���̾#ʽ��r�>�QJ�zP�8����p0�/: ��i��X~�>�;���Ѿ�	3�"h�����"�B���s�0ʺ>*~O?B�?��a�%T��H�N�����|��)?UOg?��>r?-Y?_�������M�=�n?�n�?|�?�>�>V�	�L�?D�?3	�?��?j]L?�(#�[�?�&�=�h�>���=j��>4�=�ρ��)�>t�?t�%?J,?�I��]��6����*���M#>,�6=f&�>�>�3�>�>����eC=9�)>&u�>��;>�D�>v�	?0��>mDa�K[�a?&ƼS��>���>�!�>��='�����=�\׽br��x5F��)I������h�����;��м���>��Կ}��?It">g��f?�㾁����>L�=͕��i��>��W>˹�=	��=)Q�>�>�L6>؂{>2[Ӿf�>,��@r!�Y5C��R���Ѿ�Yz>X̜�0�%�#��h����JI�Y����t� j��5��.=��_�<�E�?����ϻk���)�q(��z{?�"�>�6?�ь��i���>���>?��>�+��Ht������w�U�?���?�;c>��>)�W?��?��1��3��uZ���u�e(A�e�I�`��፿ ����
�{���_?��x? yA?�O�<*:z>:��?��%�mӏ��)�>�/��&;��@<=�+�> *���`�;�Ӿa�þ8��HF>��o?:%�?\Y?�SV�Ҳ=�-2:>�7?�P:?�6{?��M?LH3?��6�F�?�>r=?��?��A?7j ?8=?XA>��=Y��=k��=�R���f��/��.��h��<��>=8&=/51<dX�<&u�=�h�<T�ܽVT���;�5=�=y̹=��=%�=b��>��]?�L�>���>�6?�B�\6��y����.?�`=H�w����N�������W�=5�i?�M�?7FZ?<l>
?���B�v>�0�>�z$>̆h>G�>Ʊ㽔Q?�~|t=)�>��>�d�=dFY�0Z���~	�����a��<��$>���>cf�>6�����>�图�ώ��}z>�|E��d���L7�2�A�Y�5��A�����>�O?0�?.�c=��nP����_��?9E?IY3?ځ?�Ό=?�Ⱦ\�1��^J��P(��7�>��=/�9���ʡ��$�EK�/^>[�'���Q,>+V��� �]�~��EC��;߾p.R>�� �x13=�-��6ž�S�����=�2?>V����������(����J?�=����l��|T�=��c>W��>T��<"&=�A�D�i�>���>��_>�\_�hվ3�R����O>��0?�n?iF�?��l��Mq�V�(�j�	���A���=�m%?��B>.34?���>��O>�o�>��?Qj���;�\��>��>�{V�\KB���e�����'�E�k>��>p���+<6?��? E?t�?(�=?o�?�6�>r�=.׾��?<ǁ?|�=����V<�R�B���B����>��*?3�O��>Y?O�6?_C9?�/\?;'!?�mX>����q4G�j��>��>�yW�/(��mn�>V�@?ỵ>[b?4�~?@��=e]:�9a�����J��=\G>�-?
J?6%?v��>��>�x��F�Y=�N�><�]?RM�?�n?��=�S�>�AJ>���>'Eu=\�>�W�>�6?!M?>fv?��P?L��>|�O<~3��(.���z�W�	;G��;T�L<��B=ŧ��V����/��M�<jY�<'�O��<	#A;��\���a<�L�;���>�W>Pz��E��=��龔Ȉ� e><�ߎ���ȾrP���;�=�l>�A�>�?>{L����<�,�>B �>%#�1I?v+�>�_?�v���{�w���B@��p�>b�C?�jV>6�^�\E���|�����<��V?��2?r\?����p`?�K?� ��vE�и׾� �\x��9}D?��?
��'F�>u�o?�DT?�>�yK�c�m�L^��:Z������$>�9A>-( ���b��F�>W?(�>��N>�b�=㣾T�f�hO����?���?i�?
{�?��+>��s��6ֿ��i�����`?���>�AY��|
?���<�0���_v���#��J��赆�e4Ҿ "ҾEJƾr�޽���Dc~�"�>�?x�|?s|?��m?s�����~��VN��,���T�+v��k&��;�US�)M���b��	��\��ɷ����s=����SA�숵?u�'?��.�N��>@���M�X̾��D>)Ş�I��v�=,Q��z==�^=��f�p�.��֭�c�?Y�>�M�>��<?�N[��G>�0U1���7�����h1>�|�>���>0I�>";Z�,��)轼�Ⱦ3����ӽ9�@>�mm?�xt?`R�?�����sS�|:���7�<�=m �<�o�>S>�>�zž��ɽ�ܶ�{:���u�ꎐ�veܾ��3�3�E>�q!?��	�zC�>���?u��>�����=�_־s�]��ѽ�r�>��o?{�>d��>|�������>sw?n>�>E�>Mzn��H0����]��	��>P*�>�?Ί�>�����Y�����{���.=���=i�`?8�u�V��aކ>oCc?EҊ�OmO=E�>h.���3��پ..���5>d{�>iѤ=`��>�볾�-�C(q��R_��	.?�?p����.(�3�R>��(?I��>��>3�z?�Ҧ>P�ݾY�:|v?%�]?� P?=??��>�����m��
ܽ*�
��[�=��>�U0>�2�=�5>E�����i�^����=��>���9�����<����i��<���=`�x>Q$῞�s�p��B�(� BھV���GZ����>�Eܾ��˾Ҧ��n9ݽ�_�^b=� �=�x��FZ�t{��fd��,@^��?'����Ow��� r���
h??�.��u�n ��>���Ҿ�Ͻ׾�Y��LL�]�9�r���3?����O���]���,�ܾ:�>?6�	?��{?�t:�s�8�4�w�ڸ2>Qr�%�<����i��i.�M]n<��V?��>�>����>J�??Z0>_F�>����ľ�D���!?Oh�>z�>Q�ý5��cҾ�G��=���?c�?�A?s�(� ���U=��>1�	?z�?>��0�Gk��D����>z�?=Պ?kpH=~�W�����e?�<^`F�f,ٻG��=I�=�=^���K>��>� ���@�F�ٽ&}4>Ⓟ>���2��&^����<�I^>�ҽޜ��Մ?Dy\�f���/�ZT��`>��T?�,�>?0�=ǲ,?�8H��|Ͽ��\�M(a?0�?i��?��(?Q߿�<Қ>��ܾs�M?�B6?D��>�c&�L�t�a��=��i:��D��M%V����=J��>�>և,�~����O��� ��=�A��п5��}��T
J=��<=fݺa����q�\�;�l�����N_>�mQ>0�>�*�>�Va>$�.>��k?�da?��u>'=hU:��t7�y"x�l�=>�ϲ�`>u�--I��ݑ��/���Ṿ����{����7�©���𩾄�4��(�o^�ގ���1�IN�c(��Ka?�G���)�U�)�+":>O���䁾S�="���ľ�����m�?�,Q?�M��	E�XqD�`��`OO�=�i? $�ϔ�&j��@*��yü%$켮@�>0P�=k�̾�L�~ᇿ�1?\�?����ԋ����=oo��<�S=wV*?Y��>�o�;��>��?dD�����.]>��=i�>���>�i>�,���/ݽjt?��N?m
�]��?�`>d�ƾT���[�=p/>)QC�Sp���>K3������(,�=�o�����=�V?��>}*����>����X'�WDD=��w?�?���>�Qj?e�B?!(~<����R	T�;`��^=W?�'i?V>P���4qϾ�2����5?��f?hS>��g�҉�Ϟ-�G����?�m?u?��1���z�2ޒ����w�5?pv?�UR�]昿�{��aLO�g��>]a�>�|�>-�;�H��>� 3?�J�q���3���z/�G�?ѫ@�-�?�:�=ӯ]�٧�=��?Ay�>��������ڹ�DG��~��=%J?�j��4�j�v�	�%7v���=?SȆ?��>��d;��.)�=?�A�ue�?��?�8Q�s�)��W��n����ؾ�Z�<�=?�l�2��V'�f�D�����Q�ھ�����'5=)��>�
@4�C�>��$�z����˿o�u�s2?�唶��)�>C��>��:�ǌ��/e��|�MqY���T��K�3�>�!>���H��X�|�D3�p�F<Z��>sG�WE_>��W����:����8<6��>�w�>7S>!^��Ũ��攙?���uƿ����?w����g?|_�?�?��?M��<�0~��)��](�VOE?�~?>`?ϱx��@t��0'���i?I詾�:`�Q4�R7E���T>D�2?���>C�,�4�Y=(�>��>)>��-�!�ÿ�Զ�O���b�?��?/뾰.�>���?ж*?�x�NQ��\f����)��=;xA?;7>���b�!���>�����	?^s.?��ڕ�]�_?)�a�M�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?M^�?h�?ص�� #�b6%?�>b����8Ǿ��<���>�(�>*N>WH_���u>����:�i	>���?�~�?Pj?���������U>
�}?�#�>]�?!��=u�>�c�=���i�3�:F#>Y>�=��>�$�?t�M?IG�>��=��8��/�\F��BR����C���>'�a?�L?�b>a���]�1��	!���ͽ]-1���鼛Y@��,���߽_K5>Y>>�I>[E���Ҿ�V?��`�׿󷖿7g'�Pe4?��>�?\Q��cr��H�M�\?{��>��Bѳ�]���������?̲�?N?*�׾KG��->?�>B��>�Ž����ȅ�:;>�<B?�L��R���m���>c��?�[@П�?Sg�G
?��+E���#z�u!��)���=�6?kT����>���>D~�=fTr�A����ds��x�>IV�?��?���>�j?_Hn��?���=�>,k?ɠ?u�]����I>�0?�:�"V��� ���b?�@4&@�]`?V���hֿ����YN��K���7��=���=І2>%�ٽL_�=��7=��8��>�����=x�>��d>:q>_(O>�a;>�)>���J�!�r��Y���R�C�������Z�A��Xv�Tz��3������?���3ý
y���Q�2&��>`�p�=��P?�CY?Ur?���>�g��U�>pq��/&6=ܽd�=�I?>=z'?	�B?$>)?���=Vo��Cj��z�lK��*Q��"0�>r;H>�T�>���>���>X�o��UR>�|>t�>�>S��=�(Q=Jr
=�}\>��>«�>� �>�gf>�=�=�9��_{��ƀ{�h�.�Db�����?梲�{�;�����yP��襾[z>%�?��Z=RZ��a������ER?)}ξt������C�>��Z?Y|D?~I>�f���i�a���.�����}�A=��/�=���|\��r�>�)?�l�>�>pDB��0��*z��S�%1�=�]?������<(ve�ؼO�奾�zB>I�?b�#=d��D>��;Ơ���r�r:>�4;?w$?��uƾ���ž�.�>�f">�s�<&�P>ə�>��=t'��o���
b	>sh;>ٟ>P�?� >Ш����>�#��[c���t�>;�>�m:�a]?��?�'2���='���XR���Y>��?�	?d�>.�\�=͹=��>I&F>.�=x�ʽ�*�u����>9��=X�>���A��=�*9�O(>i�>�/���}	�<�~?���䈿	�6M��.nD?�-?��=��E<>�"������B���?��@�i�?�	�6�V�<�?�A�?�����=g|�>�ԫ>BξϖL��?2ƽ������	��/#��Q�?f	�?��/�Gȋ��l�>@>�W%?��Ӿ�S�>K� ��ᘿ�9���'u��`�<���>��D?��}�����9�0
?P�>lr�⮢�I�ȿI�y����>�c�?x͓?$�l�02����B����>_��?�\?MK]>tcӾ҈H����>S�9?,3J?L��>9���z���?z�?���?A>䳨?��q?��>Q�>Cㄿ�ſF5��%�)?*�ڽPm�>��@>E8Ͼ��W��U����I�?pL��~�L|�>���=��>��콫�;w=*n�KB��3>���>A�>��l>�T�>4T-?h��>l>� >iY{��`��>���4L?�׎?[��L�m���<��=�[�wf?ő3?���uҾ��>uN\?��?�t[?"[�>d���Қ�����23��_^�<��N>~-�>���>,���/R>�jԾ�>�W�>�ә>@����پ󗀾�V���>�� ?*�>,c�=��?A4"?��G>�,�>�F��G��Z>��R�>�>��?�7x?�g?8����o2�p����ꢿ�5^��N>{�x?��?�J�>���������:*'��!f0���}?��a?�н�?�?��9?J�>?ay�>l�K	޾�����>w�@?�Q�O;B��6��֓��N?0�>���>]�'���>������-��u&��&�>���?��?]#,��{w�t������E����:=���=�!=-�,>qY��^p|=_����>�xս1�����PCV���T>��>�\>9�]���r*?K�<	�^��o�=�\��N+���4>��=�쫾&k�?N��Ƈ�K��1ק���I�~��?��?ͅ�?@��<��y�V|A?R��?	�?��>i|���~پ)���k�����:��#<�� >���=���4���������٥⽰�L�h��>x��>N�?"��>���=�L�>����d��"����˾m'}�F����.� ��̄��[I-��$���{ϼ���6��� ">����Ǩ>�?w�>��>ß�>��s�t�>"��>��>e��>��>���>�X�=��!>z����O?����:�4�y���Ԍ�jK?)|?
��> *������d(�e?���?9�?�v=��������?�"/?�PžCx&?QGe=�9<��پ��yu]�O�ýW>r/�=�t4��  �|6J�w���T��>�>%�9=y���J��E���ׂ= ��? k(?�K(��6S�><n��-X�G�P�C*���g�����ki'�i�p�T���.��O#���[(�
?=�D)?�R�?������l��'�l�a�@�/se>��>78�>���>��E>��	���0���]�`'��o��YW�>Ũy?���=�nR?Y�P?�Fb?D�u?	�;��p>]����v?�=!�wS?��+?Q?9?��8?�dS?�
P?�W;?Jd>����4{	��Tݾ�4?
�)?A+?b�?��>����@(S����=��5�(����M�ah�����O^���O��~���%�>��)?ݰ�2N�p��,e>��;?�C?���>�� ��������K.�>�� ?�f�>Q�#�����a���:?��?��ʼ^/�<MW>Â�=�� >Oow=`�1>�sY�j�.>���<x_�=X�I=@Zw>X>��<���>�"�>�!:<�z�<�v�>��?��>RB�>F��1� ����o�=T�X>�S>>`Dپ
}���$����g�:y>�u�?�w�?� g=��=���=	���M����������<m�?�A#?�YT?���?�=?�i#?�>0��K��zW������?��'?_�>���I&ʾ����"1�zA
?��
?��b���.�"��ɾN½�>�)%���y�DC����B��z���U�B�R����?C��?�YO�Yc6����1"��{����@?HT�>���>a��>2�&���l�|�!�JQH>���>��V?N��>R�S?�[z?a�W?�-]>]}=�~?��D����<[�>�[B?���?	�?��t?��>M�%>�_%��۾�_������_���/��=L�O>�ܓ>���>e�>���=��ҽ��8�ge�=$�Y>1��>�B�>r1�>C8�>��<=
H?U��>R���*!��������l"7���t?��?��+?��=���a�D����4N�>�ç?��?#�*?L�O���=\<��Ƶ�;�r��E�>9U�>X�>��=tdI=k]>�_�>���>c���}�VY7�2.��?@�F?�G�=��ſz�q�H�p�ݳ���Nc<�����d�����Z����=����/���ߩ��\�F���R����鵾������{����>�.�=���=ڳ�=��<ȇɼy&�</K=?͍<�|=��o�e9m<w<9��Fϻx���)T�
\Z<��I=�����Ͼt�x?L>F?'�*?2>?Y�g>�*>�����e�>���?�:0>�J�����=DF��c��C{����־�4Ӿ��r� ��p�>J���\>PM0>��=� =�>ꃔ=�=�
�<�Y5=@��=ി=0��=y��=�G*>��>�6w?X�������4Q��Z罥�:?�8�>g{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?Ati��d�>M���㎽�q�=L����=2>p��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ4a/>��G>��>�Q�Rd,��s��WP�vW��c ?7";�
T���z{>a=�-۾V˾��<N�>���=N�GPR��o�=Pٌ���0=�K=-��>�bH>���=����-��=��=I�=uM>D@<�K%��EH�:�=F�=��z>>=(>Hk�>�?Ϟ/?.�`?�Я>+X���-ԾOgľ�>7�=��>���=W�>���>8�A?�L?�_Q?���>��:<<��>,:�>�7���r��7ž-Τ���p<��?���?Tގ>�p���W!��'�C�0�@{���?�'0?G�?׃>��	��Ov�D(���;����wr��Ɓ�B9<ɡ���*k��-e�B��=z��>b�>�վ>Wk�>��O>m�>��>�f>z��=l�Z=�cT��R9=�&=� �=w�Z��r�z^�%�"��+��=� �<>�<�`V��\�:�
��Aڬ=��>Y>8��> �=C���
5>0�M+���+>���no�h^���z���5��d9����>[�O>��A<�\��c�>Q�=�O>��?��[?*�>� 7�KH�����eJ"���kԙ=�˩>,����37���_�D�`�����;��>�ώ>�Z�>l>�7,��?���x=S���05�`�>�Ɍ�}��X�Wq��3�����x�h��$�y�D?�4��(7�=�}?��I?r��?�o�>�ś�;LؾTs0>�����d=���+r�r���?T�&?R��>r��E�D�)mž;����i�>y�D�� P�LF���~/�����!��w��>�ߨ�i Ҿ7�1�eT��[���OD�F�b��}�>�O?T�?�h��'��MM���5�s�Uo?��c?���>��?�?qު�E�Ug{�W��=<p?y��?��?(�	>c�=�;���v�>��?�6�?H�?��s?_L`��i�>L�F<zzA>\��Z>F,�=}�<�x�=�j?�{?R�?O^Ľ��=�۾D��:H��=Ggc=��>�c�>�c�>0�>���=)��=YL>�?�>M;�>W`_>�b�>�>��žʙ��J�?�j=cȶ>�h?A�>��۽I�)=W0>è?>4.��C#%���#�R�m���w=� >T�&>�F�<+�>��ɿ$ϰ?���<by��p��>���J������=���>�y���>A��<���=f��>ݾ�>�R�=��E>Zz>�'���*�=���S����g�=^K�M����ծ>G/��-�� x
�sE�<�rǽ/Fy��d�g8c�}u�5�.��'���?�L���e�,�8�� ��p�'?���>j-?�mX��&��g�{�?8X?>�!Ѿ�����)�H��?�F�?Gc>�>��W?Ę?��1�
3�DrZ�ۧu��)A� e��`��ߍ����Ӛ
�n"���_?��x?xA?���<\6z>���?��%��Џ�+�>B/��";�<=�$�>���[�`�n�Ӿ��þ�4��0F>��o?�&�?Q\?�LV������X>�zr?݇p?V4�?3?�A?�p��.iG?�V>=O?�I)?	�(?`Q?֮?�Z�>�ñ>�����=E��Uc��@d�_�,�SHA���=D'=L�:�)�:<�0=�=�t�[��<�=�̼F%!� ��<�*>%k\=���>Y�]?bE�>��>�7?���n[8�n���E(/?��9=����⊾�ǡ�
���">��j?�?�HZ?%�c>��A��}B�P.>Z,�>='>A\>�_�>ej�&rE�f?�=�>�>xs�=�UP��]��}	������<�>^?�x>C!佔[�=nɾ��ƽ�֥>�����l�����zJ4���)ԣ����>��H? ��>4Ռ<��ؾ�¼u�Y��?,�?�qG?�P?;(�������J�4�c��84��I�>�a���y7��wګ��kv�.��=G`�>c`-��ߠ��b>a���޾`�n�1_J��|��M=Uc�aU=�k�^�վ�e~��,�=�s
>����?� ��	���ڪ�`�J?�Aj=�S����U��Q��ԉ>���>��>�4�)�x�L�@�p���S�=���>x:> ��sg�nG�N��l>�F?Z�u?Hk�?��\���2^N�L�վd4���x��/F?�%�>�*�>����/�>	}��Db���=�H�k��>���>�M3���R����*���a�+�?��?�/=�?��? 6?���?�R?5?�;�>�n=:����?C��?[y>�Ά=�F)�צG���O�*�?Y:/?�_����>�I?#K?�{?:<]?�D.?��>��־��6�Uǧ>�҉>��k������f�=��D?�
�>��Z?,�?�w)>8�B�h�B��]>��>��=XzZ?p 0?�?_ �>���>�����=���>tc?�0�?�o?���=?�?�82>��>���=���>���>�?�WO?"�s?��J?k��>���<8���7��JCs� �O��ڂ;uH<��y=M��90t��I����<�"�;Nk���M�����R�D�����i��;���>�Es>�<���.>��ľ�W����A>1ٓ�J8��L��r�:��W�=���>�?��>Ʃ"���=h�>^U�>����(?`?��?�+.;5b���۾l�K�m��>�B?1��=tAl�3Y��Kgu�R�f=k�m?�~^?"X����p�b?a�]?�m�2=���þVb�8p���O?��
?Z�G�+ͳ>v�~?x�q?;��>J�e��/n�^���Gb�L�j��ȶ=TZ�>�W���d�.D�>j�7?�U�>!�b>���=(f۾	�w�H���?��?���?���?��)>��n��4�JL�n���k|d?u�>��J�?��F�r7Ծ*猾�,������G¾u����˰��C���Y0���u�S/�� >��?N�q?#?��Z?az��[^d���S�	v��=`Y�����K&��'5���J��F�hTk�V��&?�m����<��}�D�=�tx�?��)?����|�>&O��l�iž�yZ>q�s��I�e�=E,���+9S��<^�Y�R{��y��H$?�>,k�>\e8?�[��=��+���:�y+��T>dك>暠>�R�>pZ���@�gM��=}Ǿ7:��'����f>�w?��o?���?{�:=�>=�@����N4�zi���Pܽ���>bu���(>� �l���2�0|���g�d�����Պ'�N��<s&�?�S�< T�>��?���>v������[��}Z�`Q�<�j�>��?��r>N�?����0	�Ɯ�>`m?.#�>��>���Ds!�!|���ѽѬ�>Ӡ�>���>�h>'�+�|�[�����
*���q8��b�=Nh?�u��	�c�U@�>J�R?Эۺ-�R<�מ>��f�~j ��P�C�"��>jH?�L�=�@>hľMA���z�Nۉ�P�*?�!??_��Ǟ0�~�Z>�.*?S��>�>?׋�>��˾R a=�B?Χ^?��B?�P5?���>s�¼��T��'�HZ���b=\�>ܭ@>�=�m:=�)�c�j���n��<��=��}�e��K���H`�+&�<a�$<  >>�fͿ�,B�f�ƾ<�i����B����r����gx��Dپ�7M�K��s�~� ?�=s(�����ۅ����w�?���??vо��S�G��"����%��+*p>9E����z:���_�Vᔾ���
ҫ�k�;�uK<���|��q�{\.?�e��� Ŀmm����&�E�"?��B?C�u?��龇A3����j>�p���=�ჾ�ꏿ��п�O����C?Fu�>kK��a�;�>w� ?*�D>��T>��A������߃=��*?� ?w��>~e��o������	޺I��?��@��C?��jӾ�c>���>�*?���>&�����������>~Þ?E�?�1>�1\�71(��Ro?eg
>�zо�<�7o��S�=�a<���g�O>�Y�>m��� ľ�ǂ�=�^>�8|><�>Ho��l���Qt<O�>�>J�
=��?=�U���f��b,��2~���>��S?)b�>�=5	+?��F��ϿJZ���]?�4�?D��?�U'?�ʾ�n�>�oھ>N?<z5?�>\�%���t�(��=>U�9S=C�� �T����=���>m >��>�,��B�ѻ��`��=���;i�����.���h=)3��b���唽�!μ��½�(P����t��.9>�@>d�>Vs�>�6>���=|�S?v	o?�%c>1�aڐ��.��V6���{>i㰾��m��)�����;dD���4ɾ����H(��������ͥ�s�:��m�=1Q��ы��6(��l�S�@���+?�h">��ʾ_�U���j<r��v��R+ۻDK˽��ȾQo1�F�q�?��?IV<?�߉��
X��4�q+�o��_?RJ���H�ǉ����=����؁X='�>sN=�d���1�.�S���/?��!?i ¾�����>�9���Y=c�+?D?��r�wǞ>�((?*�%�3t���U>N0>愝>�(�>Ѕ>R���{]ҽ@F?�sQ?��罹�����>�����=x����<��	>�%�{�����e>wu&�󞙾A�+� ��#�=�P?
��>'c��pܾ �x��
�<c>3cv?w�8?߯�<��E?�_?��>�v����P��w��T�=D�F?�@y?r'>V剾|g�{�� UJ?�}v?�&0>Aý�%��@���� ?Gވ?U?��c�H��k�N�9���V?��v?#e^��d��J����V���>�[�>��>u�9�|��>5�>? �"��9��輿�de4�(��?W�@��?~ @<��l��=�O?�C�>��O�'sƾ�6��"�����q=zF�>�����av�����g,� �8?ܗ�?b��>�Â�٫�b=�=�P����?�$�?�M�Q��E!�Ӛp�;/�"qO�x\=��4�c�����KN�i6���L��	;�r;>=�-�>� @�q;�k�>�3���Կ���t�W����B��Ӽk>a�>ϴ��CH���]�L�]�q#8�qm\�S��Ĺ�>��=��&�7�~��`��(�a�N~=�>;O<dB,>�$�`��psC����<��>��>�I>/������E��?�d�� ׿�*��T0/���k?A��?��?Ѹ.?_������Fv<��lҼ�:S?\.T?K�4?�^T�es�ȍ����b?h%��٣�� ��7Q�!OZ>�8?���=�=��T.>
��>�-?��?��A���ÿ﹕��. ���?�u�?Y�����>��?�z�>��'Ʈ���ȉ|�w�;5��?\�=ĳ̾�6m�wM|��Η��g?�Z?Lj;<3�0�n�_?y~a���p���-�/�ƽ��>V�0�A\���˯��Se������4y���?�W�?��?���"#�&%?ݯ>�~��`Ǿ��<Vp�>m��>�[N>�_��0v>����:�q�	>X��?�x�?D>?4��������>��}?���>��?��=|��>ؤ�=������%>�7�=��:�W?��M?���>�(�=^%8�5�.��F�*cR�A��I�C��:�>��a?�CL?7�a>����q:��� �"νu�0���Y�>��1�N�޽�c4>�c<>��>k7E�2Ҿ�?�o���ؿBi��hm'�64?e��>��?#��ĸt����c<_?�>6��+���%���=�m��?�G�?��?��׾�F̼=>p�>ZH�> �Խ	
��+�����7>,�B?��3D��l�o�J�>b��?��@"֮?�i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?wQo���i�B>��?"������L��f?�
@u@a�^?*W�ڿy����G��|N��TZ>_}�=�%�=�c��!
N>j��=��=)z��So;䀘>|�\>fr�>���>�>ߴ�=M������w���y���_2�������v��04Q�"����%������U��w�˽�[j���r�O�����=v�U?zR?�;p?� ?RTy��K>e����m=�_#�_�=r�>dV2?mnL?��*?TP�=�k����d�_���>��~χ�Q��>�I>�z�>S#�>84�><�:�YI>��>>Q��>Sf>��&=m�˺TV=�N>�t�>I
�>�f�>Ρw>�aʼ<B�����
���@�5:�=�6�?�G;���d��3��CL�F��#
Z>u10?W�޼�I��v5ſꭩ��W?0Ծ���G��� >�	?2o?\!�=����=��*L�>^6� "ҾR�9>5\�<���s;L�B,:>��C?��>��>��<�(��8B��;E�]Ǝ>U�8?i��z-���e���I�/m˾��S>��>h��= �
�����Ҡt��Td�saB>r4?�b�>;=޽����z|�����@�>��=귐�32
>b�~>ۨ��P��K��"�=��6>�0�>��?�>+>;I�=���>	����C�)f�>yRL>46>�s??Q�"?��������8}���,���s>��>�y>0`>��L���=Rw�>�1b>�}��v�]��%�A��S>�(h���a�5�K�\�U=nř�Ub�=�܉=Y��+:A�*�5= �~?O��䈿L뾍e���lD?j+?�=;�F<��"�" ���G���?Y�@�l�?k�	���V��?�@�?�
��·�=Z}�>׫>3ξ��L���?.�Ž�Ƣ��	��(#�xS�?��?��/��ʋ�?l��6>H_%?��Ӿ>�>Y��o��<ƃ��q��T=� �>��I?e������7�?�n?s�很ϣ���ǿR�p�Y�>ӯ�?0I�?u�q�a���E=��%�>�$�?�W?;�n>f �~dg��e�>َ;?P�X?���>A�wM3�M�?38�?��?o&>���?9�?
(q>xa�>ȷD��������8>A5�<�e�<p6���f��d�q����zT�)�Y�C:����)>2+�=�u�>7���_��A�= Ո<�3������\�>:l�>��>B�>v��>��>"��>��=e7a�mX��l�����K?�ʎ?�O� um���<�q�=�pU���?�g5?����1ѾW�>��Z?CW�?�&Z?`#�>����
��!ɽ� Q����=��Q>�>&�>k�z�B>�Ծ��:��2�>��>��Lپ�e|��n��b�>�o ?,��>^��=�� ?$�#?F�j>C*�>:`E��8����E�q��>^��>�D?�~?��?ҹ��V3�����塿��[�<N>��x?XU?ƕ>H���c�����D�I4I�������?Gqg?�g�=?�2�?��??.�A?uf>ђ��ؾ
���X��>�*?C�ƻ<H��/�F��f�F?j�>Z�*?���%;�>�|�������^J?�/T?�x?�+)�%&y���8�A��r�=`,���$>�=�h=�	;T���7'�d2V>��=�ٲ�~��n���-�C>B�>7T�=,�Y�3]��A*?!BT�Kz*��j�=�(e�Q�Q�V�s>� $=��ľ+x? 3!���[��X��q��������?��?�$�?F6��<k�R�8?�!�?�?���>:.˾�^���׾3i���kN�t�'�>K^=Kfw>Í�<bk̾/碿/��f�����Ե(���
?���>bn?��?H��=PC�>W3���:���ƾ04����y�?
�@�*��D8��A!���l���	%�<"�ѾW���eT>S?)=C
�>�q?ar>�r�>���>U���(�>��=o׋>Q+�>��|>]�>���=�؟=nM��r�R?�[��� (�9��#۱�m�D?��d?P��>��tՂ��;��?!��?xA�?�xv>�c��r)���>i��>.��M?�)|=�]�����<�ʮ�GD0�S}�������>Z��b�2��[E�>`�K?�?���;�'̾%�ͽ�e��qs={k�?�&)?5[)��R���o���W�\�R��a���h� ꡾�$�h�p������G��[�#D(���,=�c*?M�?mK�����櫾��j��)?���d>�>���>\��>��I>�
�eY1�u�]��@'��]�>r�z?섍>ЋI?��;?(zP?.jL?a��>�]�>�+���z�>Y?�;#�>���>�9?��-?�%0?�j?r+?Lc>������d�ؾk?F�?�I?_?=�?�Ʌ�>�ý�����c�F�y��	����=&��<��׽��t�z[U=�$T>nH3?�)�� "V��7��i�"Y?��G?OG?�da�q��ſ�=?��=oC?P��2ވ���C�_�6>tzy?�F�w��<P�U>H~S=# >Ɂ�=v��<�ͽR��= f=�2ѼBؗ�� �<A�=��,�={j=���=����6�; t�>|�?���>SD�>�>��O� �.��a�=�Y>�S> >�Gپ�}��L$����g�<[y>�w�?�z�?y�f=��=6��=M}��T����?������<��?�J#?�WT?e��?R�=?4j#?[�>�*�M���^�����w�?,?S��>=���ʾ�稿?t3�å?�Z?��`����j9)��m¾q�Խ��>?/��~�]����D�j,�����H7����?x��?U�@�5�6�aO�a���o���^C?��>	Υ>-�>��)��h�w1�,�:>\��>:R?)̺>A�O?|?T�^?q�V>Ř8�Vȭ�⿙��$����">�s@?�S�?�ߍ?�4t?�J�>�>�;!���߾X}��\�#������4��H�j= "Z>�؏>��>���>�ʸ=��ҽh���Q�4��Ԡ=��d>���>�%�>q��>�-}>*�<�}C?\Y ?�)̾����z���c�9R}<y�l?B��?��?��ٻX���37�u�Ӿ)�>7Π?��?0�?ѣF� 4�=�4�;cE���9���>��>4�>�!�=��>-�)=�\�>U;
?B)۽����7b�^Z�, �>��d?�'�>'}ȿ��t�i�`��瑾��<�-��;v�����M6�_B�=q/��Vh������S��+��A���"���x���,l��>�>�Nl=�>UF�={��<"���6�<39B=g3
:-��<�ې����<t�	�����v��'p��,3=<x�=�?ͻՇ˾�}?�)I?'�+?��C?�ry>�>�4�g��>�%���O?0U>SP�go����;�+Ĩ�r��wbؾ�>׾�d������G>�H�{�>�R3>�,�=���<���=!�s=���=�-a�i=1��=�к=�y�=��=��>�W>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>Rv8>c>��R�Yy1���\�J�`�^�Y��!?�8;�[L˾�>>�=6?߾�ž��4=�8> �]=�3�"]\�j�=t�w��:=�-n=��>�C>u��=�d��R<�=ܒF=���=��N>LV��!Y8��,�@�0=y�=�b>|4&>�>�>�-?8�0?f.e?�1�>��p��Ͼ�B���F�>��=�˲>r#�=i8D>d�>�E8?�fD?�lL?�V�>j�=Fe�>��>�'-��*n�^��s����<´�?��?Q۷>Tl=<D<�k��*�<��7Ž_q?��1?Ae?�V�>�I��̿�����"þB�=�	�{�A���Ĕ#>�oi��XüF��\C�n`x>c�>~:�>��>���>5R>W�>!��<�.=��q=ν=!��=ˤ�=I�#<*D�{�����uv=K�j>0==��i9�=�˙���	>�OʼP*�=���>��>�9�>��>>v�����=��S�T��5�>h���L�2���I�6Cw���M�s����>Y��>���=�����`?⿽L��>���?��r?QE�=���=)�v�?l��O�T��T=��>�^A� :;��q�7��iƾ_�>�l�>��>�9m>3?+�d"?���v=r���4��&�>Y�����'�U����p��Q���ڟ�Dwh��p:ŮD?�?��1��=2}?��I?�Ə?F��>W9��Լ׾�r2>|���=��hp����H�?��&?b��>�{��kD��H̾D���޷>s@I��O���Y�0�ۮ�#ͷ�?��>�����о_$3��g��������B��Lr�s��>'�O?��?u:b��W��=UO����v(���q?�|g?�>�J?�@?�%��z�r���v�=�n?���?H=�?c> �=����x��>��	?�g�?`~�?Qq?�J:���>���ӄ*>�󪽿��=t�>��v=��=��?�b?Q?�T�����>
���W�"=kq�=��>�ن>��s>[�=�rK=���=��Q>���>f�>��i>�a�>N�>&�����zB"?�%d>X��>��?	��=HZ�<��R=�'>�/>�پ�+��i�*Bn�v}��\�)=L�t>Ǡ�=!W�>8�̿�,�?W�L>�-�yr?#����X��=��G>
2��W��>��W>��C�PN�>!�>;}�=�c>��>ΗѾ��>X��VJ ���B�U�Q��Ͼ>{>!�� M)���U�콘$H�a&�����)i��́���<��~�<��?|b���/j�i�(��W����?�>��5?����6���}�>��>w�>����QY����\�?�+�?R�`>��>�Y?q7?�,'��=�/[��Gv���@�s�c�w�`�}荿�l����5׽��\?eAw?��@?���<l�y>Q�?L�#�η���ϑ>��.�-�;�l&=#?�>�2���p�W1Ͼ��Ⱦ|��S�?>E9l?u�?�M?��Z���m�( '>��:?�1?Ot?,�1?�;?����$?Yo3>�E?r?�M5?��.?��
?2>N	�=?L����'=�7��~��ѽ�{ʽ��1�3=�]{=�Pָ��
<l�=���<����ټ��;$��Y �<G:=f�=��=��>��\?��>
Y�>�K7?u�)��%8�l��%J$?��M=�4c�>����)���� �|6>�G_?�֪?��S?�O>�$D��xM�0�>�T�>l(>�qK>��>�Ȫ��0X�\�2=�_+>D�2>8��=���gj���
��1~��#Z=�>��>�܏>��ǽ'�*>5I��/A_�5z>�E7����N�]���E��f.��l��{�>TUL?� ?S��=�[H��)�]�ߒ)?[�??Q�J?QQu?���<��ľO�4�4�/�+HN��`�>�p�=�3 ��=�� ��w�<�_Ao�}�>��T��젾�)b>V����޾�n�J�����QN=����U=
�A�վ_����=\�
>D���� ���eت�EJ?	�j=!~���KU�m����>���>�߮>�p9��Hw���@�:���:��=ͯ�>�	;>�̛�
�|G�3��I>bX?��x?ހ�?�Y�������f���0�]@��q;>�@4?�>F�>� �\8�=J���cҾպv�l�W��'�>�{?~��dD�>�p��@	�ׅ9���)>'X?k@+><)'?4vv?ӗ�>��D?�!?�	?S$s>�eͽ�H��}A&?'��?��=[�Խ��T�� 9�sF���>��)?D�B�s��>��?5�?i�&?H�Q?N�?��>t� �ND@�ܓ�>EY�>;�W�:b����_>1�J?���>j=Y?�ԃ?��=>S�5��颾eԩ��[�=>K�2?�6#?�?���>���>b���/��=�k�>l�b?n0�?��o?9�=��?��1>�>qD�=���>Ġ�>C?�@O?��s?��J?�t�>P-�<򑬽hM��Os�$�^��H�;�I<�Cy=>� �Au��1�S��<���;4|��_y��d�^�C��󕼚<�;��>���>\]��f�P>��k����"?>�< �e֎��_���c��;<���>�,�>Ĵ�=�;ǽ]�W>��>(��>IJ%��/?��?��>��)�H�m�'Y� ��\t?�|?���<��p�.'��Q�g���=���?1�?� �5|�
�b?��]?Ge�y=��þ*ib�Kf���O?
�
??�G��ܳ>��~?��q?���>��e��(n�[���!b�'�j�(��=�s�>�P��d�hߝ> 7?�V�>��b>��=��۾w�w�Dl����?��?�?��?�_*>0�n�0�'���{����V^?�)�>L��8�"?�j��]Ͼ�Ή�B,���q����g���l5���Ŧ�`g"����bٽĻ=��?~Yr?��q?�l`?Q �Qd�V_�&Q��q�V�����S�|#E�?�E��.D��ym��
�Z����4��"Y9=�՜� �%��<�?�C0?��Խ��>=t��R��oܱ���>��c��֜�X��=�q��ܻ��=a$3���O��۪��p?A�>�)�>[M?�LF�s�E���T���S�#%��=>�A�>K��>ym>]��}|c������ξ�'����q���:>c$f?,�m?se�?GBn���K��ɗ���J���� ��\��>/��=�r�="v�-��:���np�2恿(�F��k����;_�=�#?��=�i�>�K�?�K�>�����ٳ�|{޾�9f��0�2?�d?[��>J��>��^��5����>&�q?v�>���>ٍ�L,�l$i�l�!��A�>{>�>gM�>U/>՞8�aa�Fy���;��2
A�/�>s�`?�=���J]�
AK>S'T?A�!=��2��>Q�i�'�0�-M����H�S�>|(�>%��<s��=��־��K_�äZ�,�)?�?24���*�Y�{>��"?���>J<�>{�?n3�>��þ�ա�ؚ?��^?��J?��@?g��>��=�ڴ��H̽�!��.*=�>.SR>6 `=�>�=�����V�2 ���D=8��=��ܼ�_���S<�P���)]<�$�<G�1>���V�T�fᾩ	�S��!Z	���o���ؼ$������o`��E�������Kӽ���<X����"���p�.��5��?Σ�?�N�rվT|��d�n������?[����� �LԾ�ɝ��.��|\���*�����_�1;u�1tq�-�?
��˸����+�3��/?05?�"�?*�V��?�;Fj�Yk>��K>k>��z�^�����:���b/4?���>`�#�x�=f��>���>	�>��>�{����V��X8�P�?m_F?���>�d�U5˿	Ŀ:���ͤ�?.v
@�F@?1�)��&����<�>5?wSR>�� �����ڻ�P�>B��?%��?���=��W��돽�\?�L=��.�O1�;�E�=尒=�)ϼ�ý�#>�&�>k	9�\�7��''���?>�ܐ>�Q�����9��ld�<�C>����#�/Ԅ?s\��f�͡/��Q���}>��T?H2�>ʼ�=�,?E5H�&uϿV�\�a(a? -�?���?��(?�׿��Ț>��ܾ��M?<6?6 �>|o&�2�t�W�=jv�L������V����=S��>NU>o},����xO��j��g��=��Q�ƿ��$�'}��Z=wq޺i�[��}�د����T��"���ho���轇�h=w��=�Q>Xm�>�&W>�1Z>fW?^�k?�H�>�v>@佂���	ξ���+J���������������P��߾�	�_������ɾ�BZ��+�?�[��ؙ�Ю9�h|T�Q���J?���;D>ؾV�J�w	�F��V�^�7�T> "<dw��2�1��~�!��?��E?=ю��=R�� O�H�e=�>��c?�����Zb�h>z=)�{=��>Jo~�+2���I�Z�!�0?�z?7￾����P�&>tX뽚*&=�w+?Y�?ˉ"<-)�>�#?��,�޵ؽ\<b>�J1>��>{��>�q>�į��ƽg�?�S?f�����;�>�8���Mo�wV=F�>�6;��{��R>5�<�A��#��q���D��<Y�V?�U�>p�)�JI��-��Ae"�I=�Pw?�E?/�>=5h?Q�B?�.�<�����S���C:o=PW?#Ui?/>=e��E�˾E����5?'xe?oN>��a�y�꾀+�ri�n�?S�o?�p?�@���<|�3����\���6?�v?�n^��q�������V��9�>Y�>���>(�9��m�>)�>?N#�"G�����lY4��?T�@���?K�;<:�u��=�??\V�>�O��Eƾa��{�����q=	$�>&����dv�x��V,�p�8?ݡ�?���>������o�D=��K�浱?9�?�Xi��E
��'���u�����Q>l> >՛�(�����x'�{������u����1��>�@�r߽���>��н.��S�ҿ�>���7ݾ<S�1�?�>�>6�v��7��>�>�]KT�70�v�N�7>þ#�>��>} ��E摾��{�3h;����m
�>�Y�E�>��S��+��u����3<��>:��>���>����j���Ù?�f���(οŝ��ء�T�X?�i�?�l�?.o?�V7<%�w��{���74G?4ts?H�Y?di$�B]�/�7��*j?R���*�_��5��9A�6Y>�H2?	��>z-�S�q=}>�f�>y�>��(�%�Ŀ���5�� �?dJ�?Ǽ��Y�>��?��'?0S�톚��$��?*��-
�9D?v[8>�����!�)K<��4����	?�,?*�뽣w���_?.�a�W�p���-��ƽ�ۡ>h�0��c\� B������Xe�����?y����?F^�?4�?Z��� #��5%?��>����
8Ǿ�<N��>�)�>]*N>�H_���u>���:�;j	>���?�~�?�i?!��������W>�}?}%�>k�?j�=�`�>e�=g��,�k#>�=��>���? �M?N�>`T�=G�8�A/�XZF��DR�x"���C���>H�a?��L?@Gb>���W)2�{!��lͽTe1�gQ�[@���,�^�߽�#5>��=>�>�D�}
Ӿ.�?�p�3�ؿ�i���i'�054?��>��?�����t�����<_?>{�>_2�=,���%���C�7��?FG�?��?��׾�L̼�>;�>UB�>�ս���&�����7>T�B?��D��4�o���>?��?Q�@!֮?�i��	?s��P��a~����7����=��7?L0��z>���>�=�nv�˻��I�s���>�B�?�{�?���>îl?H�o���B�O�1=�L�>3�k?�s?8po�	��B>Q�?)�����L��f?�
@|u@�^?/����LӠ��ɭ�������=�]�<5M%>1C���=-��=|��<���To=���>�[>�q�>�l�>�1i>m��=�;}�s��ỿם��Q�S�k��e��s	=��"�G��Zj��
����̾��D����;�<��r��:N)�]���=��U?��S?�q?� ?����Y$>����Ut=N����=�>�}0?��J?JF,?��=X�I�f��b������ц�x�>�rH>�L�>��>�-�>��;M�L>�>>�E~>4v>�K?=/��;�=�DN>4�> ��>2�>O�=�ʆ=5A��M᱿���R��<�a�?��p���H��g��о��̼���`�=��L?O>>>N����ȿ�󰿻PZ?YΩ��j�����PT�<Z�A?�qY?4�>L&�N��8�ļ��k�6�K�
�>��^�J3���#�#W�>�N-?5�>fI>��7�sOA���P�lڠ���>h%?�Q���'�o�q�L�N�6&��;>�l�>���<�\+�D^���.q�0�}��5>�K/?�s?��LB��u궾���s"^> rI>1!.���Z=��1>V���2�D���2�=B��=�a>�g�>;E^>G5�=�U�>~���n�u��>��>E�<>>�B?��?��������%7I�]u�>%?��>��=e�k��Ը=sJ?S�8>t��՜�c!��~P��nF>�������Kq��~�<\ʽf��=N��=����H�u���<�/~?@���@ň��{�w�����D?�n?ᶔ=�.d<�#��馿�y����?��@0�?]�	��0V�`�?�/�?�&����=���>�/�>(�̾{�L��r?ګɽ΄���%	�ہ ��+�?ba�?`f$�Ƌ�F�k���>�|%?zҾa��>�/���$���a���N���>�_�>2U=?�l�,�j^G����>˔�>��߾E������)[d����>��?�߅?����В���F:�H��>���?��f?���>�E������Z&�=͓F?�fx?n�!?�����&�9? ֧?Mg|?*�@>|��?��w?�p�>�.���5��'���|��O�v=�=H$�>0�>-�Ͼ�J��׎��ށ��aa�L����<>x�J=���>��U����=*���S[��ˌS�Cָ>.�t>ash>���>H� ?���>��>��_=�ڡ���q��>����K?<��?���2n��4�<ų�=��^�V'?�K4?��[�T�ϾXԨ>��\??�[?d�>���-=��*翿P��  �<$�K>b4�>�>�>�0��&BK>��Ծ�)D�o�>�Η><O���?ھ�/���&���@�>�d!?d��>̮=׉ ?�x#?��h>G|�>��D�����E��Q�>#��>��?��}?�?q��K3��Ւ��š�S0[��3O>G�x?^H?r>$���Ꮭ��	#���@�f���R��?�=f?�<ݽ�?T�?h@?*�A?2!d>K��kv־������>�r"?����H��|F�x�x���>�?���>cf�<�9��6���@������	?GIU?�P?�F-�]�X�!ש�Ҏ�<A">�,t����=�O<M����<p�P�,�M=���>4	7�(���J|*�̴��iAs=���>v>f=�,��&	�W!?]=7H�9��=�h���L��@_>��>˜���oe?��M�Вy������m���q�5��?g%�?@&�?$�̽�fh�v�.?í�?(�	?� �>|���X��\@ؾ����J-a���q>���>F����۾蠿����ZU���	&�FE�]'?���>P�?�T�>�/G=���>�{�������۾�����d�س��1��h8���d�eS�%b�=�'���?ɾ�J3>K��)��>b�?(��>Q�>���>��ɽm�t><��>�G�>r9�>�%d=�>���=Ps>՗-��@?���q'�W��o���`?rB_?�?�9>�̀�F+ ��%?ӣI?]y�?��>��R��M)���?ʴ�>�1'���>%l����t�� �̠��4Z̺\���"]=^��>�I��� ��[���a��.�>�*
?Eﲽ@��.%�d���>jo=H�?��(?��)���Q�o�o�u�W��S����[,h�bt��9�$�g�p�鏿!]��%���(�d�*=�*?�?��r���W k�??�Tbf>���>r�>5޾>�I>��	���1��^�-P'�'����Y�>6[{?y;�>��I?<?&~P?�lL?܍�>s0�>�8�����>6�;��>l��>�9?�-?0?��?��+?��b>��������ؗؾ	?_�?�,?!?̨?����	�½�:��Af�~�y�������=0�<�׽یu�9!U=G�S>XH&?@��#�}���P>׺3?�n ?�/?����P���T���v=?~='?�W?Cn�WMz����iU?Ȍv?w�</>�j>?K>��U>0"�=8D$�Ӈ�=o�/=T�>��$>���">�����
>s\>�۽~�>���\k�>��?L��>�C�>�<��� ����}4�=��X>�:S>��>OEپ�{���"����g��ky>y�?As�?g�f=[��=�N�=�Q���W�����.󽾛v�<�?m5#?�TT?m��?%�=?Jk#?��>�'��J���V��y����?�,?���> ���ʾfѨ��e3��j?h?��`��y�)�^�¾�׽�f>$ /�p ~������C���j�v���Ҙ��m�?y��?;��v6�r�)����-���<C?���>���>���>W�)��g��{�u�:>�>�QR?2�w>�l?���?q��?A?�>H@p��Pƿ���p}����>�P�?��{?1�1?Ob�>��>S�?��<��%��z9�17���H�)p���=�~�=��f>��>G�>�����v��M���V[>6	>���>Q�>b�>-/�>O�<��G?��>�[��6���뤾�Ń�=��u?���?^�+?�G=G����E��F���H�>�n�?���?3*?�S�(��=��ּ�ڶ���q���>zչ>C/�>��=�|F=�d>T	�>@��>,��`�7p8�eHM���?2F?��=rƿ��q���p��˗�a�c<������d�*�����Z��j�=���%���̩���[��y���*���ʤ��4�{����>�y�=���=��=���<Wɼ���<�
K=�Í<��=�
p���l<j�8�7л	����1�ޑ\<��I=s��̾��}?oI?F�+?��C?D)y>N�>6�4�?�>r����C? #S>A#H�dR��:s=���%����ؾ"�־�'d�#a��H�	>�5K���>�Z4>��=Q�<���=	y=U�=�|�Y# =#��=k��=��=w��=�S>)6>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>z�7>\d>�R�W1�'�\�[�b�BZ�-a!?�0;��̾�>l�=�i߾W�ƾ��-=�R5>l�\=�G���[�Ӕ�=(-|�H==Ģm=�5�>ɌD>l�=�G��:s�=��H=���=m<P>�$��ǝ6�U�/�ʺ.=���=��c>IS'>�.�>(?O�0?zwd?iQ�>u�n��vϾ�����x�>z��=瑱>k�= �A>�><8?��D?�
L?ʹ�>�W�=#��>���>Bb,��~m��E�ѧ���<:��?`ʆ?٧�>|�L<�eA��m���=���ýp?��1?9?m��>�U����9Y&���.�$���z4��+=�mr��QU�N���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=$�����<�vż�����u&�:�+�1�����;r��;B�]<^��;�K�<-�?(�>>��>��=Q�ھ�W�=����6�S�"�:>��ѾF�:�V�S���p�*�5��]ν9��>W��=3��<�n��_x�>>�=���>5��?K z?�]>P[��_��㧿������o�5 ->�|>鹌�avV�w`�;�A��L����>��>��>��l>��+���>���w=����m5��$�>�g���t��*��#q��6��퟿�h�a>g�d�D??��],�=��}?��I?�Ϗ?]o�>������ؾG�0>�W��%�=���sq��ؓ�6�?z*'?���>2���D�r�˾��]�>үG��O�����<;0�2^�]:��G��>
s���оo	3�^���׏�2�B���r���>��O?�Ʈ?.Xd�p���O�A�Xt��Gi?��g?��>�h?4�?�Ǜ�o,��~��E�=p\n?���?��?p`>0��=�I�����>��>L��?�M�?��m?������>BŞ��O�=&96�W�4>޺C>��=lx�=�r?,�?1)?f�~�[t��f����iG1����<���=��c>���>��y>��=M�=y�=���>筀>�X�>�dn>2p�>zۑ>�����w��`�?�@>Ŭ�>�� ?��Y>S�=j�j<�.�<Ӈ�3b��*�=��	����w=|��=�&�<6�u=a�>.���՟?b��=k��/�?���X>��7)>Q3�>b\����>�\>��'>���>�<�>��w=
h�>6��=������*>�R����Π:�?�H�Z[ž��Y>����S����[��+�����ʾ���y�i�;h����3�U,z=n�?���k�V�QO�=�)��q?Eۢ>�9?d�������$1P>I�?Q��>m��ѓ�l@��
̾�d�?���?|�b>)�>�lV?*�?%/�p�5�
Y�a�t���>�љa�p'_�8��n����
�
=ɽsI`?��z?��@?���<�|r>��?3@ �����u�>�E1��g:��s)=��>٬��.d�f%Ծqʾ���&�F>�q?��?��?��^��m��"'>z�:?��1?�Ot?<�1?��;?h���$?�m3>�F?�o?O5?��.?.�
?&2>!�=�'��=�'=�8����L�ѽ�ʽ���3=�_{=2�¸hV<��=C��<���x�ټ�(;����D�<��9=��=-�=_�A>lb?��'?���>;1?����}I��(߾��7?�<>ٓ�������ۘ�z�羵�>R�?2G�?�� ?�*���^��/���>&]x>b�>�>5I�>]󣼨6�v7�=�O�=�-->qN>���=q���𾏷~��B�<aMp>���>���>$�<�.%�=��Ⱦ�MK�>Tj>�J��=4p/��2�(�=�gϚ��o>�D:?%&�>������!S���c[�s�b?߫?u��?�SQ?�y�}���V��?��$g�DO�>�ֽ��������F��� d��6���>X΢<�ߠ��b>a���޾`�n�1_J��|��M=Uc�aU=�k�^�վ�e~��,�=�s
>����?� ��	���ڪ�`�J?�Aj=�S����U��Q��ԉ>���>��>�4�)�x�L�@�p���S�=���>x:> ��sg�nG�N��l>�F?Z�u?Hk�?��\���2^N�L�վd4���x��/F?�%�>�*�>����/�>	}��Db���=�H�k��>���>�M3���R����*���a�+�?��?�/=�?��? 6?���?�R?5?�;�>�n=:����?C��?[y>�Ά=�F)�צG���O�*�?Y:/?�_����>�I?#K?�{?:<]?�D.?��>��־��6�Uǧ>�҉>��k������f�=��D?�
�>��Z?,�?�w)>8�B�h�B��]>��>��=XzZ?p 0?�?_ �>���>�����=���>tc?�0�?�o?���=?�?�82>��>���=���>���>�?�WO?"�s?��J?k��>���<8���7��JCs� �O��ڂ;uH<��y=M��90t��I����<�"�;Nk���M�����R�D�����i��;���>�Es>�<���.>��ľ�W����A>1ٓ�J8��L��r�:��W�=���>�?��>Ʃ"���=h�>^U�>����(?`?��?�+.;5b���۾l�K�m��>�B?1��=tAl�3Y��Kgu�R�f=k�m?�~^?"X����p�b?a�]?�m�2=���þVb�8p���O?��
?Z�G�+ͳ>v�~?x�q?;��>J�e��/n�^���Gb�L�j��ȶ=TZ�>�W���d�.D�>j�7?�U�>!�b>���=(f۾	�w�H���?��?���?���?��)>��n��4�JL�n���k|d?u�>��J�?��F�r7Ծ*猾�,������G¾u����˰��C���Y0���u�S/�� >��?N�q?#?��Z?az��[^d���S�	v��=`Y�����K&��'5���J��F�hTk�V��&?�m����<��}�D�=�tx�?��)?����|�>&O��l�iž�yZ>q�s��I�e�=E,���+9S��<^�Y�R{��y��H$?�>,k�>\e8?�[��=��+���:�y+��T>dك>暠>�R�>pZ���@�gM��=}Ǿ7:��'����f>�w?��o?���?{�:=�>=�@����N4�zi���Pܽ���>bu���(>� �l���2�0|���g�d�����Պ'�N��<s&�?�S�< T�>��?���>v������[��}Z�`Q�<�j�>��?��r>N�?����0	�Ɯ�>`m?.#�>��>���Ds!�!|���ѽѬ�>Ӡ�>���>�h>'�+�|�[�����
*���q8��b�=Nh?�u��	�c�U@�>J�R?Эۺ-�R<�מ>��f�~j ��P�C�"��>jH?�L�=�@>hľMA���z�Nۉ�P�*?�!??_��Ǟ0�~�Z>�.*?S��>�>?׋�>��˾R a=�B?Χ^?��B?�P5?���>s�¼��T��'�HZ���b=\�>ܭ@>�=�m:=�)�c�j���n��<��=��}�e��K���H`�+&�<a�$<  >>�fͿ�,B�f�ƾ<�i����B����r����gx��Dپ�7M�K��s�~� ?�=s(�����ۅ����w�?���??vо��S�G��"����%��+*p>9E����z:���_�Vᔾ���
ҫ�k�;�uK<���|��q�{\.?�e��� Ŀmm����&�E�"?��B?C�u?��龇A3����j>�p���=�ჾ�ꏿ��п�O����C?Fu�>kK��a�;�>w� ?*�D>��T>��A������߃=��*?� ?w��>~e��o������	޺I��?��@��C?��jӾ�c>���>�*?���>&�����������>~Þ?E�?�1>�1\�71(��Ro?eg
>�zо�<�7o��S�=�a<���g�O>�Y�>m��� ľ�ǂ�=�^>�8|><�>Ho��l���Qt<O�>�>J�
=��?=�U���f��b,��2~���>��S?)b�>�=5	+?��F��ϿJZ���]?�4�?D��?�U'?�ʾ�n�>�oھ>N?<z5?�>\�%���t�(��=>U�9S=C�� �T����=���>m >��>�,��B�ѻ��`��=���;i�����.���h=)3��b���唽�!μ��½�(P����t��.9>�@>d�>Vs�>�6>���=|�S?v	o?�%c>1�aڐ��.��V6���{>i㰾��m��)�����;dD���4ɾ����H(��������ͥ�s�:��m�=1Q��ы��6(��l�S�@���+?�h">��ʾ_�U���j<r��v��R+ۻDK˽��ȾQo1�F�q�?��?IV<?�߉��
X��4�q+�o��_?RJ���H�ǉ����=����؁X='�>sN=�d���1�.�S���/?��!?i ¾�����>�9���Y=c�+?D?��r�wǞ>�((?*�%�3t���U>N0>愝>�(�>Ѕ>R���{]ҽ@F?�sQ?��罹�����>�����=x����<��	>�%�{�����e>wu&�󞙾A�+� ��#�=�P?
��>'c��pܾ �x��
�<c>3cv?w�8?߯�<��E?�_?��>�v����P��w��T�=D�F?�@y?r'>V剾|g�{�� UJ?�}v?�&0>Aý�%��@���� ?Gވ?U?��c�H��k�N�9���V?��v?#e^��d��J����V���>�[�>��>u�9�|��>5�>? �"��9��輿�de4�(��?W�@��?~ @<��l��=�O?�C�>��O�'sƾ�6��"�����q=zF�>�����av�����g,� �8?ܗ�?b��>�Â�٫�b=�=�P����?�$�?�M�Q��E!�Ӛp�;/�"qO�x\=��4�c�����KN�i6���L��	;�r;>=�-�>� @�q;�k�>�3���Կ���t�W����B��Ӽk>a�>ϴ��CH���]�L�]�q#8�qm\�S��Ĺ�>��=��&�7�~��`��(�a�N~=�>;O<dB,>�$�`��psC����<��>��>�I>/������E��?�d�� ׿�*��T0/���k?A��?��?Ѹ.?_������Fv<��lҼ�:S?\.T?K�4?�^T�es�ȍ����b?h%��٣�� ��7Q�!OZ>�8?���=�=��T.>
��>�-?��?��A���ÿ﹕��. ���?�u�?Y�����>��?�z�>��'Ʈ���ȉ|�w�;5��?\�=ĳ̾�6m�wM|��Η��g?�Z?Lj;<3�0�n�_?y~a���p���-�/�ƽ��>V�0�A\���˯��Se������4y���?�W�?��?���"#�&%?ݯ>�~��`Ǿ��<Vp�>m��>�[N>�_��0v>����:�q�	>X��?�x�?D>?4��������>��}?���>��?��=|��>ؤ�=������%>�7�=��:�W?��M?���>�(�=^%8�5�.��F�*cR�A��I�C��:�>��a?�CL?7�a>����q:��� �"νu�0���Y�>��1�N�޽�c4>�c<>��>k7E�2Ҿ�?�o���ؿBi��hm'�64?e��>��?#��ĸt����c<_?�>6��+���%���=�m��?�G�?��?��׾�F̼=>p�>ZH�> �Խ	
��+�����7>,�B?��3D��l�o�J�>b��?��@"֮?�i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?wQo���i�B>��?"������L��f?�
@u@a�^?*W�ڿy����G��|N��TZ>_}�=�%�=�c��!
N>j��=��=)z��So;䀘>|�\>fr�>���>�>ߴ�=M������w���y���_2�������v��04Q�"����%������U��w�˽�[j���r�O�����=v�U?zR?�;p?� ?RTy��K>e����m=�_#�_�=r�>dV2?mnL?��*?TP�=�k����d�_���>��~χ�Q��>�I>�z�>S#�>84�><�:�YI>��>>Q��>Sf>��&=m�˺TV=�N>�t�>I
�>�f�>Ρw>�aʼ<B�����
���@�5:�=�6�?�G;���d��3��CL�F��#
Z>u10?W�޼�I��v5ſꭩ��W?0Ծ���G��� >�	?2o?\!�=����=��*L�>^6� "ҾR�9>5\�<���s;L�B,:>��C?��>��>��<�(��8B��;E�]Ǝ>U�8?i��z-���e���I�/m˾��S>��>h��= �
�����Ҡt��Td�saB>r4?�b�>;=޽����z|�����@�>��=귐�32
>b�~>ۨ��P��K��"�=��6>�0�>��?�>+>;I�=���>	����C�)f�>yRL>46>�s??Q�"?��������8}���,���s>��>�y>0`>��L���=Rw�>�1b>�}��v�]��%�A��S>�(h���a�5�K�\�U=nř�Ub�=�܉=Y��+:A�*�5= �~?O��䈿L뾍e���lD?j+?�=;�F<��"�" ���G���?Y�@�l�?k�	���V��?�@�?�
��·�=Z}�>׫>3ξ��L���?.�Ž�Ƣ��	��(#�xS�?��?��/��ʋ�?l��6>H_%?��Ӿ>�>Y��o��<ƃ��q��T=� �>��I?e������7�?�n?s�很ϣ���ǿR�p�Y�>ӯ�?0I�?u�q�a���E=��%�>�$�?�W?;�n>f �~dg��e�>َ;?P�X?���>A�wM3�M�?38�?��?o&>���?9�?
(q>xa�>ȷD��������8>A5�<�e�<p6���f��d�q����zT�)�Y�C:����)>2+�=�u�>7���_��A�= Ո<�3������\�>:l�>��>B�>v��>��>"��>��=e7a�mX��l�����K?�ʎ?�O� um���<�q�=�pU���?�g5?����1ѾW�>��Z?CW�?�&Z?`#�>����
��!ɽ� Q����=��Q>�>&�>k�z�B>�Ծ��:��2�>��>��Lپ�e|��n��b�>�o ?,��>^��=�� ?$�#?F�j>C*�>:`E��8����E�q��>^��>�D?�~?��?ҹ��V3�����塿��[�<N>��x?XU?ƕ>H���c�����D�I4I�������?Gqg?�g�=?�2�?��??.�A?uf>ђ��ؾ
���X��>�*?C�ƻ<H��/�F��f�F?j�>Z�*?���%;�>�|�������^J?�/T?�x?�+)�%&y���8�A��r�=`,���$>�=�h=�	;T���7'�d2V>��=�ٲ�~��n���-�C>B�>7T�=,�Y�3]��A*?!BT�Kz*��j�=�(e�Q�Q�V�s>� $=��ľ+x? 3!���[��X��q��������?��?�$�?F6��<k�R�8?�!�?�?���>:.˾�^���׾3i���kN�t�'�>K^=Kfw>Í�<bk̾/碿/��f�����Ե(���
?���>bn?��?H��=PC�>W3���:���ƾ04����y�?
�@�*��D8��A!���l���	%�<"�ѾW���eT>S?)=C
�>�q?ar>�r�>���>U���(�>��=o׋>Q+�>��|>]�>���=�؟=nM��r�R?�[��� (�9��#۱�m�D?��d?P��>��tՂ��;��?!��?xA�?�xv>�c��r)���>i��>.��M?�)|=�]�����<�ʮ�GD0�S}�������>Z��b�2��[E�>`�K?�?���;�'̾%�ͽ�e��qs={k�?�&)?5[)��R���o���W�\�R��a���h� ꡾�$�h�p������G��[�#D(���,=�c*?M�?mK�����櫾��j��)?���d>�>���>\��>��I>�
�eY1�u�]��@'��]�>r�z?섍>ЋI?��;?(zP?.jL?a��>�]�>�+���z�>Y?�;#�>���>�9?��-?�%0?�j?r+?Lc>������d�ؾk?F�?�I?_?=�?�Ʌ�>�ý�����c�F�y��	����=&��<��׽��t�z[U=�$T>nH3?�)�� "V��7��i�"Y?��G?OG?�da�q��ſ�=?��=oC?P��2ވ���C�_�6>tzy?�F�w��<P�U>H~S=# >Ɂ�=v��<�ͽR��= f=�2ѼBؗ�� �<A�=��,�={j=���=����6�; t�>|�?���>SD�>�>��O� �.��a�=�Y>�S> >�Gپ�}��L$����g�<[y>�w�?�z�?y�f=��=6��=M}��T����?������<��?�J#?�WT?e��?R�=?4j#?[�>�*�M���^�����w�?,?S��>=���ʾ�稿?t3�å?�Z?��`����j9)��m¾q�Խ��>?/��~�]����D�j,�����H7����?x��?U�@�5�6�aO�a���o���^C?��>	Υ>-�>��)��h�w1�,�:>\��>:R?)̺>A�O?|?T�^?q�V>Ř8�Vȭ�⿙��$����">�s@?�S�?�ߍ?�4t?�J�>�>�;!���߾X}��\�#������4��H�j= "Z>�؏>��>���>�ʸ=��ҽh���Q�4��Ԡ=��d>���>�%�>q��>�-}>*�<�}C?\Y ?�)̾����z���c�9R}<y�l?B��?��?��ٻX���37�u�Ӿ)�>7Π?��?0�?ѣF� 4�=�4�;cE���9���>��>4�>�!�=��>-�)=�\�>U;
?B)۽����7b�^Z�, �>��d?�'�>'}ȿ��t�i�`��瑾��<�-��;v�����M6�_B�=q/��Vh������S��+��A���"���x���,l��>�>�Nl=�>UF�={��<"���6�<39B=g3
:-��<�ې����<t�	�����v��'p��,3=<x�=�?ͻՇ˾�}?�)I?'�+?��C?�ry>�>�4�g��>�%���O?0U>SP�go����;�+Ĩ�r��wbؾ�>׾�d������G>�H�{�>�R3>�,�=���<���=!�s=���=�-a�i=1��=�к=�y�=��=��>�W>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>Rv8>c>��R�Yy1���\�J�`�^�Y��!?�8;�[L˾�>>�=6?߾�ž��4=�8> �]=�3�"]\�j�=t�w��:=�-n=��>�C>u��=�d��R<�=ܒF=���=��N>LV��!Y8��,�@�0=y�=�b>|4&>�>�>�-?8�0?f.e?�1�>��p��Ͼ�B���F�>��=�˲>r#�=i8D>d�>�E8?�fD?�lL?�V�>j�=Fe�>��>�'-��*n�^��s����<´�?��?Q۷>Tl=<D<�k��*�<��7Ž_q?��1?Ae?�V�>�I��̿�����"þB�=�	�{�A���Ĕ#>�oi��XüF��\C�n`x>c�>~:�>��>���>5R>W�>!��<�.=��q=ν=!��=ˤ�=I�#<*D�{�����uv=K�j>0==��i9�=�˙���	>�OʼP*�=���>��>�9�>��>>v�����=��S�T��5�>h���L�2���I�6Cw���M�s����>Y��>���=�����`?⿽L��>���?��r?QE�=���=)�v�?l��O�T��T=��>�^A� :;��q�7��iƾ_�>�l�>��>�9m>3?+�d"?���v=r���4��&�>Y�����'�U����p��Q���ڟ�Dwh��p:ŮD?�?��1��=2}?��I?�Ə?F��>W9��Լ׾�r2>|���=��hp����H�?��&?b��>�{��kD��H̾D���޷>s@I��O���Y�0�ۮ�#ͷ�?��>�����о_$3��g��������B��Lr�s��>'�O?��?u:b��W��=UO����v(���q?�|g?�>�J?�@?�%��z�r���v�=�n?���?H=�?c> �=����x��>��	?�g�?`~�?Qq?�J:���>���ӄ*>�󪽿��=t�>��v=��=��?�b?Q?�T�����>
���W�"=kq�=��>�ن>��s>[�=�rK=���=��Q>���>f�>��i>�a�>N�>&�����zB"?�%d>X��>��?	��=HZ�<��R=�'>�/>�پ�+��i�*Bn�v}��\�)=L�t>Ǡ�=!W�>8�̿�,�?W�L>�-�yr?#����X��=��G>
2��W��>��W>��C�PN�>!�>;}�=�c>��>ΗѾ��>X��VJ ���B�U�Q��Ͼ>{>!�� M)���U�콘$H�a&�����)i��́���<��~�<��?|b���/j�i�(��W����?�>��5?����6���}�>��>w�>����QY����\�?�+�?R�`>��>�Y?q7?�,'��=�/[��Gv���@�s�c�w�`�}荿�l����5׽��\?eAw?��@?���<l�y>Q�?L�#�η���ϑ>��.�-�;�l&=#?�>�2���p�W1Ͼ��Ⱦ|��S�?>E9l?u�?�M?��Z���m�( '>��:?�1?Ot?,�1?�;?����$?Yo3>�E?r?�M5?��.?��
?2>N	�=?L����'=�7��~��ѽ�{ʽ��1�3=�]{=�Pָ��
<l�=���<����ټ��;$��Y �<G:=f�=��=��>��\?��>
Y�>�K7?u�)��%8�l��%J$?��M=�4c�>����)���� �|6>�G_?�֪?��S?�O>�$D��xM�0�>�T�>l(>�qK>��>�Ȫ��0X�\�2=�_+>D�2>8��=���gj���
��1~��#Z=�>��>�܏>��ǽ'�*>5I��/A_�5z>�E7����N�]���E��f.��l��{�>TUL?� ?S��=�[H��)�]�ߒ)?[�??Q�J?QQu?���<��ľO�4�4�/�+HN��`�>�p�=�3 ��=�� ��w�<�_Ao�}�>��T��젾�)b>V����޾�n�J�����QN=����U=
�A�վ_����=\�
>D���� ���eت�EJ?	�j=!~���KU�m����>���>�߮>�p9��Hw���@�:���:��=ͯ�>�	;>�̛�
�|G�3��I>bX?��x?ހ�?�Y�������f���0�]@��q;>�@4?�>F�>� �\8�=J���cҾպv�l�W��'�>�{?~��dD�>�p��@	�ׅ9���)>'X?k@+><)'?4vv?ӗ�>��D?�!?�	?S$s>�eͽ�H��}A&?'��?��=[�Խ��T�� 9�sF���>��)?D�B�s��>��?5�?i�&?H�Q?N�?��>t� �ND@�ܓ�>EY�>;�W�:b����_>1�J?���>j=Y?�ԃ?��=>S�5��颾eԩ��[�=>K�2?�6#?�?���>���>b���/��=�k�>l�b?n0�?��o?9�=��?��1>�>qD�=���>Ġ�>C?�@O?��s?��J?�t�>P-�<򑬽hM��Os�$�^��H�;�I<�Cy=>� �Au��1�S��<���;4|��_y��d�^�C��󕼚<�;��>���>\]��f�P>��k����"?>�< �e֎��_���c��;<���>�,�>Ĵ�=�;ǽ]�W>��>(��>IJ%��/?��?��>��)�H�m�'Y� ��\t?�|?���<��p�.'��Q�g���=���?1�?� �5|�
�b?��]?Ge�y=��þ*ib�Kf���O?
�
??�G��ܳ>��~?��q?���>��e��(n�[���!b�'�j�(��=�s�>�P��d�hߝ> 7?�V�>��b>��=��۾w�w�Dl����?��?�?��?�_*>0�n�0�'���{����V^?�)�>L��8�"?�j��]Ͼ�Ή�B,���q����g���l5���Ŧ�`g"����bٽĻ=��?~Yr?��q?�l`?Q �Qd�V_�&Q��q�V�����S�|#E�?�E��.D��ym��
�Z����4��"Y9=�՜� �%��<�?�C0?��Խ��>=t��R��oܱ���>��c��֜�X��=�q��ܻ��=a$3���O��۪��p?A�>�)�>[M?�LF�s�E���T���S�#%��=>�A�>K��>ym>]��}|c������ξ�'����q���:>c$f?,�m?se�?GBn���K��ɗ���J���� ��\��>/��=�r�="v�-��:���np�2恿(�F��k����;_�=�#?��=�i�>�K�?�K�>�����ٳ�|{޾�9f��0�2?�d?[��>J��>��^��5����>&�q?v�>���>ٍ�L,�l$i�l�!��A�>{>�>gM�>U/>՞8�aa�Fy���;��2
A�/�>s�`?�=���J]�
AK>S'T?A�!=��2��>Q�i�'�0�-M����H�S�>|(�>%��<s��=��־��K_�äZ�,�)?�?24���*�Y�{>��"?���>J<�>{�?n3�>��þ�ա�ؚ?��^?��J?��@?g��>��=�ڴ��H̽�!��.*=�>.SR>6 `=�>�=�����V�2 ���D=8��=��ܼ�_���S<�P���)]<�$�<G�1>���V�T�fᾩ	�S��!Z	���o���ؼ$������o`��E�������Kӽ���<X����"���p�.��5��?Σ�?�N�rվT|��d�n������?[����� �LԾ�ɝ��.��|\���*�����_�1;u�1tq�-�?
��˸����+�3��/?05?�"�?*�V��?�;Fj�Yk>��K>k>��z�^�����:���b/4?���>`�#�x�=f��>���>	�>��>�{����V��X8�P�?m_F?���>�d�U5˿	Ŀ:���ͤ�?.v
@�F@?1�)��&����<�>5?wSR>�� �����ڻ�P�>B��?%��?���=��W��돽�\?�L=��.�O1�;�E�=尒=�)ϼ�ý�#>�&�>k	9�\�7��''���?>�ܐ>�Q�����9��ld�<�C>����#�/Ԅ?s\��f�͡/��Q���}>��T?H2�>ʼ�=�,?E5H�&uϿV�\�a(a? -�?���?��(?�׿��Ț>��ܾ��M?<6?6 �>|o&�2�t�W�=jv�L������V����=S��>NU>o},����xO��j��g��=��Q�ƿ��$�'}��Z=wq޺i�[��}�د����T��"���ho���轇�h=w��=�Q>Xm�>�&W>�1Z>fW?^�k?�H�>�v>@佂���	ξ���+J���������������P��߾�	�_������ɾ�BZ��+�?�[��ؙ�Ю9�h|T�Q���J?���;D>ؾV�J�w	�F��V�^�7�T> "<dw��2�1��~�!��?��E?=ю��=R�� O�H�e=�>��c?�����Zb�h>z=)�{=��>Jo~�+2���I�Z�!�0?�z?7￾����P�&>tX뽚*&=�w+?Y�?ˉ"<-)�>�#?��,�޵ؽ\<b>�J1>��>{��>�q>�į��ƽg�?�S?f�����;�>�8���Mo�wV=F�>�6;��{��R>5�<�A��#��q���D��<Y�V?�U�>p�)�JI��-��Ae"�I=�Pw?�E?/�>=5h?Q�B?�.�<�����S���C:o=PW?#Ui?/>=e��E�˾E����5?'xe?oN>��a�y�꾀+�ri�n�?S�o?�p?�@���<|�3����\���6?�v?�n^��q�������V��9�>Y�>���>(�9��m�>)�>?N#�"G�����lY4��?T�@���?K�;<:�u��=�??\V�>�O��Eƾa��{�����q=	$�>&����dv�x��V,�p�8?ݡ�?���>������o�D=��K�浱?9�?�Xi��E
��'���u�����Q>l> >՛�(�����x'�{������u����1��>�@�r߽���>��н.��S�ҿ�>���7ݾ<S�1�?�>�>6�v��7��>�>�]KT�70�v�N�7>þ#�>��>} ��E摾��{�3h;����m
�>�Y�E�>��S��+��u����3<��>:��>���>����j���Ù?�f���(οŝ��ء�T�X?�i�?�l�?.o?�V7<%�w��{���74G?4ts?H�Y?di$�B]�/�7��*j?R���*�_��5��9A�6Y>�H2?	��>z-�S�q=}>�f�>y�>��(�%�Ŀ���5�� �?dJ�?Ǽ��Y�>��?��'?0S�톚��$��?*��-
�9D?v[8>�����!�)K<��4����	?�,?*�뽣w���_?.�a�W�p���-��ƽ�ۡ>h�0��c\� B������Xe�����?y����?F^�?4�?Z��� #��5%?��>����
8Ǿ�<N��>�)�>]*N>�H_���u>���:�;j	>���?�~�?�i?!��������W>�}?}%�>k�?j�=�`�>e�=g��,�k#>�=��>���? �M?N�>`T�=G�8�A/�XZF��DR�x"���C���>H�a?��L?@Gb>���W)2�{!��lͽTe1�gQ�[@���,�^�߽�#5>��=>�>�D�}
Ӿ.�?�p�3�ؿ�i���i'�054?��>��?�����t�����<_?>{�>_2�=,���%���C�7��?FG�?��?��׾�L̼�>;�>UB�>�ս���&�����7>T�B?��D��4�o���>?��?Q�@!֮?�i��	?s��P��a~����7����=��7?L0��z>���>�=�nv�˻��I�s���>�B�?�{�?���>îl?H�o���B�O�1=�L�>3�k?�s?8po�	��B>Q�?)�����L��f?�
@|u@�^?/����LӠ��ɭ�������=�]�<5M%>1C���=-��=|��<���To=���>�[>�q�>�l�>�1i>m��=�;}�s��ỿם��Q�S�k��e��s	=��"�G��Zj��
����̾��D����;�<��r��:N)�]���=��U?��S?�q?� ?����Y$>����Ut=N����=�>�}0?��J?JF,?��=X�I�f��b������ц�x�>�rH>�L�>��>�-�>��;M�L>�>>�E~>4v>�K?=/��;�=�DN>4�> ��>2�>O�=�ʆ=5A��M᱿���R��<�a�?��p���H��g��о��̼���`�=��L?O>>>N����ȿ�󰿻PZ?YΩ��j�����PT�<Z�A?�qY?4�>L&�N��8�ļ��k�6�K�
�>��^�J3���#�#W�>�N-?5�>fI>��7�sOA���P�lڠ���>h%?�Q���'�o�q�L�N�6&��;>�l�>���<�\+�D^���.q�0�}��5>�K/?�s?��LB��u궾���s"^> rI>1!.���Z=��1>V���2�D���2�=B��=�a>�g�>;E^>G5�=�U�>~���n�u��>��>E�<>>�B?��?��������%7I�]u�>%?��>��=e�k��Ը=sJ?S�8>t��՜�c!��~P��nF>�������Kq��~�<\ʽf��=N��=����H�u���<�/~?@���@ň��{�w�����D?�n?ᶔ=�.d<�#��馿�y����?��@0�?]�	��0V�`�?�/�?�&����=���>�/�>(�̾{�L��r?ګɽ΄���%	�ہ ��+�?ba�?`f$�Ƌ�F�k���>�|%?zҾa��>�/���$���a���N���>�_�>2U=?�l�,�j^G����>˔�>��߾E������)[d����>��?�߅?����В���F:�H��>���?��f?���>�E������Z&�=͓F?�fx?n�!?�����&�9? ֧?Mg|?*�@>|��?��w?�p�>�.���5��'���|��O�v=�=H$�>0�>-�Ͼ�J��׎��ށ��aa�L����<>x�J=���>��U����=*���S[��ˌS�Cָ>.�t>ash>���>H� ?���>��>��_=�ڡ���q��>����K?<��?���2n��4�<ų�=��^�V'?�K4?��[�T�ϾXԨ>��\??�[?d�>���-=��*翿P��  �<$�K>b4�>�>�>�0��&BK>��Ծ�)D�o�>�Η><O���?ھ�/���&���@�>�d!?d��>̮=׉ ?�x#?��h>G|�>��D�����E��Q�>#��>��?��}?�?q��K3��Ւ��š�S0[��3O>G�x?^H?r>$���Ꮭ��	#���@�f���R��?�=f?�<ݽ�?T�?h@?*�A?2!d>K��kv־������>�r"?����H��|F�x�x���>�?���>cf�<�9��6���@������	?GIU?�P?�F-�]�X�!ש�Ҏ�<A">�,t����=�O<M����<p�P�,�M=���>4	7�(���J|*�̴��iAs=���>v>f=�,��&	�W!?]=7H�9��=�h���L��@_>��>˜���oe?��M�Вy������m���q�5��?g%�?@&�?$�̽�fh�v�.?í�?(�	?� �>|���X��\@ؾ����J-a���q>���>F����۾蠿����ZU���	&�FE�]'?���>P�?�T�>�/G=���>�{�������۾�����d�س��1��h8���d�eS�%b�=�'���?ɾ�J3>K��)��>b�?(��>Q�>���>��ɽm�t><��>�G�>r9�>�%d=�>���=Ps>՗-��@?���q'�W��o���`?rB_?�?�9>�̀�F+ ��%?ӣI?]y�?��>��R��M)���?ʴ�>�1'���>%l����t�� �̠��4Z̺\���"]=^��>�I��� ��[���a��.�>�*
?Eﲽ@��.%�d���>jo=H�?��(?��)���Q�o�o�u�W��S����[,h�bt��9�$�g�p�鏿!]��%���(�d�*=�*?�?��r���W k�??�Tbf>���>r�>5޾>�I>��	���1��^�-P'�'����Y�>6[{?y;�>��I?<?&~P?�lL?܍�>s0�>�8�����>6�;��>l��>�9?�-?0?��?��+?��b>��������ؗؾ	?_�?�,?!?̨?����	�½�:��Af�~�y�������=0�<�׽یu�9!U=G�S>XH&?@��#�}���P>׺3?�n ?�/?����P���T���v=?~='?�W?Cn�WMz����iU?Ȍv?w�</>�j>?K>��U>0"�=8D$�Ӈ�=o�/=T�>��$>���">�����
>s\>�۽~�>���\k�>��?L��>�C�>�<��� ����}4�=��X>�:S>��>OEپ�{���"����g��ky>y�?As�?g�f=[��=�N�=�Q���W�����.󽾛v�<�?m5#?�TT?m��?%�=?Jk#?��>�'��J���V��y����?�,?���> ���ʾfѨ��e3��j?h?��`��y�)�^�¾�׽�f>$ /�p ~������C���j�v���Ҙ��m�?y��?;��v6�r�)����-���<C?���>���>���>W�)��g��{�u�:>�>�QR?2�w>�l?���?q��?A?�>H@p��Pƿ���p}����>�P�?��{?1�1?Ob�>��>S�?��<��%��z9�17���H�)p���=�~�=��f>��>G�>�����v��M���V[>6	>���>Q�>b�>-/�>O�<��G?��>�[��6���뤾�Ń�=��u?���?^�+?�G=G����E��F���H�>�n�?���?3*?�S�(��=��ּ�ڶ���q���>zչ>C/�>��=�|F=�d>T	�>@��>,��`�7p8�eHM���?2F?��=rƿ��q���p��˗�a�c<������d�*�����Z��j�=���%���̩���[��y���*���ʤ��4�{����>�y�=���=��=���<Wɼ���<�
K=�Í<��=�
p���l<j�8�7л	����1�ޑ\<��I=s��̾��}?oI?F�+?��C?D)y>N�>6�4�?�>r����C? #S>A#H�dR��:s=���%����ؾ"�־�'d�#a��H�	>�5K���>�Z4>��=Q�<���=	y=U�=�|�Y# =#��=k��=��=w��=�S>)6>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>z�7>\d>�R�W1�'�\�[�b�BZ�-a!?�0;��̾�>l�=�i߾W�ƾ��-=�R5>l�\=�G���[�Ӕ�=(-|�H==Ģm=�5�>ɌD>l�=�G��:s�=��H=���=m<P>�$��ǝ6�U�/�ʺ.=���=��c>IS'>�.�>(?O�0?zwd?iQ�>u�n��vϾ�����x�>z��=瑱>k�= �A>�><8?��D?�
L?ʹ�>�W�=#��>���>Bb,��~m��E�ѧ���<:��?`ʆ?٧�>|�L<�eA��m���=���ýp?��1?9?m��>�U����9Y&���.�$���z4��+=�mr��QU�N���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=$�����<�vż�����u&�:�+�1�����;r��;B�]<^��;�K�<-�?(�>>��>��=Q�ھ�W�=����6�S�"�:>��ѾF�:�V�S���p�*�5��]ν9��>W��=3��<�n��_x�>>�=���>5��?K z?�]>P[��_��㧿������o�5 ->�|>鹌�avV�w`�;�A��L����>��>��>��l>��+���>���w=����m5��$�>�g���t��*��#q��6��퟿�h�a>g�d�D??��],�=��}?��I?�Ϗ?]o�>������ؾG�0>�W��%�=���sq��ؓ�6�?z*'?���>2���D�r�˾��]�>үG��O�����<;0�2^�]:��G��>
s���оo	3�^���׏�2�B���r���>��O?�Ʈ?.Xd�p���O�A�Xt��Gi?��g?��>�h?4�?�Ǜ�o,��~��E�=p\n?���?��?p`>0��=�I�����>��>L��?�M�?��m?������>BŞ��O�=&96�W�4>޺C>��=lx�=�r?,�?1)?f�~�[t��f����iG1����<���=��c>���>��y>��=M�=y�=���>筀>�X�>�dn>2p�>zۑ>�����w��`�?�@>Ŭ�>�� ?��Y>S�=j�j<�.�<Ӈ�3b��*�=��	����w=|��=�&�<6�u=a�>.���՟?b��=k��/�?���X>��7)>Q3�>b\����>�\>��'>���>�<�>��w=
h�>6��=������*>�R����Π:�?�H�Z[ž��Y>����S����[��+�����ʾ���y�i�;h����3�U,z=n�?���k�V�QO�=�)��q?Eۢ>�9?d�������$1P>I�?Q��>m��ѓ�l@��
̾�d�?���?|�b>)�>�lV?*�?%/�p�5�
Y�a�t���>�љa�p'_�8��n����
�
=ɽsI`?��z?��@?���<�|r>��?3@ �����u�>�E1��g:��s)=��>٬��.d�f%Ծqʾ���&�F>�q?��?��?��^��m��"'>z�:?��1?�Ot?<�1?��;?h���$?�m3>�F?�o?O5?��.?.�
?&2>!�=�'��=�'=�8����L�ѽ�ʽ���3=�_{=2�¸hV<��=C��<���x�ټ�(;����D�<��9=��=-�=_�A>lb?��'?���>;1?����}I��(߾��7?�<>ٓ�������ۘ�z�羵�>R�?2G�?�� ?�*���^��/���>&]x>b�>�>5I�>]󣼨6�v7�=�O�=�-->qN>���=q���𾏷~��B�<aMp>���>���>$�<�.%�=��Ⱦ�MK�>Tj>�J��=4p/��2�(�=�gϚ��o>�D:?%&�>������!S���c[�s�b?߫?u��?�SQ?�y�}���V��?��$g�DO�>�ֽ��������F��� d��6���>X΢<�1Ѿ�A>�B"����]���$�W��s��>��u�=�-��zԾ/�8�e�{<�(>�I��&���_���}��eD?�n=�m*���G��e�o=��>�Z	?.H>�=w8��K��z->o��>�8>֔=�U羃UL��j��iqU>��8?N�?���?�J�v�����d������A�_�.?�>|��>��>�s�=�j��+��6o�T�E��j�>�l�>cC%���)�J���*�JM��r>��9?�Mn>-�?	d?>D?.�b?��?��*?U��>��	���#��?�`�?_�>x��;jK����H�����.�>�/?��b�jҭ>{�'?�4?8
"?j�c?�?�]�=��l�=�]}�>�>�>��^��Ϯ��H�>�V?7��>۟N?���?N>a*J��L��q���{�=���>??H�?1?eu�>O��>����N�=���>�c?�/�?I�o?�K�=�?��2>���>8�=8��>f��>]?WO?��s?�J?1~�>�N�<i���=����s��Q���;�I<��y=Jw���s���<(�<��;tt��Gl����̞D�^�����;ٓ�>�}o>����$>뽾P����G>jͥ��k������4�5�� �=y7�>�?\c�>+�(��/�=���>���>^)�--(?@'?��?�ȑ<�c`��4Ӿ�F�c�>�B?�I�=�.h�+Ɠ��s�G=�=|�o?-G^?s[�����$]?AtT?������@�p���40�(v���g;?{V?(�����>|?ij?5�>��Z��%c��ė�i�b�<�+�UЗ=킲>���e�{��><�-?�m�>�FX>���=�٨�5Am�Y������>/Q�?���?�ϑ?�D=>uoq��nݿ���`ɑ��j]?��>w����"?is��-ξ5*���8��)��Up��Æ�����~����#�����ֽd]�=̶?�Zr?Uq?A`?�/���c�b�]��x�8KV��������{E�ЂD�7lC��Bo��g�v���l�����Q=�D~���=��E�?r6(?�a/�_�>pј�t�p�ξ67>>�U�����a�=�ʖ�߀@=p�X=�fh��m-�� ��5�?��>X��>L�<?e�Y�Rf>�151��8������a->q�>��>�y�>�^<"�)���[Aʾ�g���~ƽ�>>#�Y?W`?g��?9��p��]�x��(��K���о�o>�%�=p�L>�y���G��u�'�s�#���S�c�+�����&�leH>s�(?�E�<F��>���?5T�>8�@�,W侨�ܾԨ"�%=���>��{?,%�>��>�f��O����>	l?O��>���>�_��`�"��O|��y���>���>8�?~ul>��-���Z��?��y,���5����=�7]?؀�ve�_�>1AS?[[����h=��>H����&�w����8��>�?iҰ=��D>nɾE����z�ȋ��s?!��>�xо��l�i�.?2I?�h?�R>^��?\�[?iB���=y����>u�l?*�Y?΅D?J��>�9�J�r�:���ͽ��ֽ8�U>\��>1~ؽ�ZԽ���=���~q[��i�~.�B}�=��d��?
=�zp���=�>���<�ݿW�L�fvܾ�������䆾�+������Lt��0��⾔�f�o�������49R�O%a�ȵ��*�o����??��?]㚾����ꔿ��w����
�>�Ql��ne������� ��m����澑����"��J�|Fe�Tec�`7
?�pþ�ݲ�s��������?��?VG�?�3о���}O�b�>�0�>���=�0��Y��
���砾�u?�i�>�����+����>7f->9D�>�D�>��&�E���Z�j�?LHI?iU�>�ĽT
���*��@r�����?�
@'VA?Hl(���쾥�Q=q�>Sj	?��A>q�,����k����D�>-�?�݊?�UT=YfX��u���c?Zn$<N.D�����3a�=ʭ=1h$=յ��I>+	�>+��P�A��<޽��6>eӆ>��4�3�T%\���<�b>AOǽ�����2�?�\���c��+�&�M>U0T?�ع>6�=��,?>�B��!Ͽ� _���[?8��?f��?��.? e���}�>�ܾąL?	�5?|��>�&�rLw�,w�=XԢ�����̦�HV�dv�=r�>>����N=L��|�3��=R������0�S���s�=��1=)��� ���-���P�����]9�3?��c�>��=C+)>�=>P�}=a��=��{?��?�?V=�0%�l+�=�c��� ������4���!=��`�=>��|��g��pP�LE��^�����D��x=x�V��l����ķR���H��1?�=��վ��K���{=l���O��B�R���ž�K.�L�c�
@�?1P;?���e�M�J���"���ƽ��\?K����~뾫c��^ڒ=�%���2<f��>i;�=��Ҿz-��K�C�)??��ʾ�Q���ؓ>�ﱽ)��<�1?(��>�>�¦>	?z��s��>m�G>kÈ>��>u��=�ԓ��U��?��{?|����R��&�T>ޭo�����bթ�V�U>�^=��!%=-a�=����.���m��x>
��=K%W?��>��)�����{��$�'$==h�x?ց?�>\ok?/�B?��<�M����S���ޒu=j�W?�,i?"�>�
����Ͼ�-����5?�ve?gO>�Nh�f��Q�.�E>�K;?��n?J?���3l}���������6?p�?��k�+�u���n�vᠾ���>�|?H�>yȣ�ܶ�>��g?��ѽ���ڐ¿%<�Eұ?�@���?�N|��K��	W�=���>�
�>S	ݾ�"#�7�����]_>=?�zƾV����=��R����D?ud�?�?�b��Pi����=X����I�?�?�����V<A����k�S9����<^­=լ��)�Qs��7���ƾ��
�;D���Aɼ�T�>�A@��彅_�>߶6��⿻AϿ(���Ѿ��r��|?Ba�>8Ƚ���dXj�q$u�"�G�D�H�oE��?�>iY>�Ò�W=����{�H;�uƥ�5/�>���א�>�R������E���)<��>��>��>�ᬽ�R���y�?���J>οu����[��X?���?�c�?�?�a<W�t�?�z�$� ��G?=
s?��Y?/�!��K]�?q4��Qj?���.L`��\4�^UD�%X>�Q3?��>�,���u=>�{�>	*>o-��hĿ���mx��w��?S��?Ր龎��>�5�?<�*?�O�4
��'j���5*�)~����@?��4> ��i�!��y=��Ò�W
?�20?d��:�S�_?�a�I�p���-���ƽ�ۡ>��0��e\��K������Xe����@y����?F^�?c�?ѵ�� #�R6%?	�>c����8Ǿ8�<���>�(�>�)N>�G_�|�u>����:��h	>���?�~�?Aj?󕏿�����U>��}?�>��?@>�=A��>D�=���������>���=�g)��	?�M?���>��=�c8�0@.�h�E�i�Q�	�B�B�-��>*�b?�J?K�j>�f��8)�t � PʽU�)�" �0�<�j�3��ӽ�c;>H>��>[�J�Y\Ծ�p&?*������灿
-�r{?���>�?��ϭ�IS=�E^?{f�>;I�pC��4���m�����?���?}O?. �D�*=�TZ>�#�>`�3>dϴ=D�&�E����->BI?7<�?P��3�z��V�>�²?�.	@�J�?NY�'1$?�+��uf�>��$оZ�k���>�~.?�%���	�=��?n>��a��3��\Um����>_-�?wA�?��>�c?="z��0����=o��>��V?���>v8@��S��4�>�%?����^�� �<�x�s?>w@gn@b�x?����g�|�����������=���=AM>r�C��:�=���=RE=�1f�p�>Ĭ�>��>���> sI>�g>j�G>����N%�8��q呿A'-�A>�ؾ&�D��O��3&��ܬ1����:쑾��%=�M�΅Ҽ�� �e|��9�z=l��=7�W?_�R?�o?��>�������=u�����'=��&���j=��>�3?��J?)�/?�3�=:G����d�H����ť��q��@l�>�+A>��>3��>�o�>��仹,F>�g@>�If>��=(�=�z.<��)=5�?>�&�>�'�>U�>j>&s>�鯿4y��z�g��&s������?����@�d��O���
��N]�=k�)?�P�=C��U�̿e禿��I?Sz���
���N���*>V�-?�l?MGA>� ���l�����=ӽ�q��ci>��7�fw��_Q%�g)D>�,#?�Pe>�Tu>��3���8�n@O�L���Oy>��6?F����4��fu�ZaH�"�۾��L><��>x�7�-���Ֆ��~�c�f� Tx=30:? A?����9V���u�n���K�P>ZYY>d�=,c�=��O>qof���ɽ�[H��!=CM�=0_>.��>��>���=���>����}hl��8�>�}}>�͐>�D?��4?��ҽV�f��o����K��N�>��>�>�^<{�E���1>F��>��>z�<����.�wvh�R��=���/?K�xa���=K�����=�_�<ODP����	�;��}?�7��񈿫�N@���gE?\�?�x�=ѥY<)q"�覿���(��?��@q�??�
�/�V�^�?�Ǝ?�����
�=��>]�>H{˾�1I��?([Ľڠ��3P	�&)��T�?�q�?������k�e�>�N'?5�оzK�>�!�����X����um�B�y=R"�>�JK?�:�W�:�.a��?��	?q(⾙a����ǿ'�t�'��>/�?�(�?�n��ߘ�k7���>t�?�X?=/>��Ҿ�U����>o0C?8�L?s�>A��U`.���?�r�?2��?���=�?�J�?�z?�z�= �l��C���m��l�=T���5`�>�<t����P�P�����Ѫa���T�1�޾=a�`!=�3�=�t�'�����S=�p�����=0��>�z>�,>R
�>f;"?a��>o��<8����Jƺ���v����'K?��?,"��n�=3=_۟=r�Z��b?��4?�a�c�ξ�ʦ>0�[?���?v�[?2��>F���M��M���sܲ��z�<�cM>�e�>�w�>Hm���E>��Ͼ SI�l��>]�>C;��>"־N���/x�H��>��?�k�>���=�� ?%�#?��j>�)�>'aE�G7����E�X��>ޜ�>@?��~?��?�ǹ�
W3��
��6䡿��[��CN>��x?RV?쿕>���~���%E�G{I�Ϫ����?�lg?ju�S?P3�?�??ϟA?�f>'��:�׾iU��*��> z?"���J2�F6�QPp=�W?}o?�s�>$7�=��5>�"��3��3Ѿ0�?��S?/�#?�����o��ʜ��jU<5N���p�≠��*U�
OH>q3>bca����=�ې>��>v@�����$>�?>�v�>�Q">�(��ɉ��:?��|�;)�<���>����Y	R�v�U>�����Ⱦ�d0?�_!�fǩ�{¶��$����>��?�m�?V��?<�I�%�~�<7Q?��?6�?���>��a��כ��*~%�����5��IX�:3�>�����jɾ�ͫ��ܺ��G�۔m��]��:?�^�>Y%?`��>�D�=��~>p�<a7�����׾$[������:�]�r���p��K��:D�������f����>�_{�UǮ>��>
|[>��F>�y�>�Ϻwԏ>��_>z�v>�d�>Y[s>�n1>���="�R��$��q2?�� �_=��'��)o�*�?n	v?���>޼'=?fJ����-? >�?Ҧ?. ���`}�!R4����>k|d?[�#���>��f<z��=���%5~���<76A��O�<�w>4�{<��"�ݑ:��8����>o�>�S%=�/���.d�Ä��n^p=�R�?��(?-�)��Q��o�޸W��S�ft�Q�g�Gs����$���p��揿,W��� ���(�o�)={*?
�?8�� ���$��� k�e?���f>��>�$�>6ž>;}I>��	�I�1��]��D'������C�>�C{?Vm�>��I?i	<?tP?�VL?�L�>-�>�F��&1�>a��;�>"��>�l9?��-?":0?�k?AO+?w�b>���.����^ؾ?~�?dP?��?y�?�1��"�ý<���og��y������A�=�U�<��׽k=v���S=�YT>��	?�n��	�N��^�zAr>G�k?� ?��2>jg��izW�n�H���?��+?�{?�"��ރ���#��U�>���?��c�Z8+>@x>"U=o�c=�E��Yt=�#��n�=��=�>�`=�����P����<^�=�
Y=������9��>�22?!�>a�>�Ŕ����,��_%>xpe>͞9>�hx>����To��el���L��p�>Yq�?��?����&=t�=M�Ծ0ξ�����#��'�>��?�M?�q?�ƒ?��6?Z�?[e�=5��c%q��nd�\V���?�9,?K��>bx���Ⱦ����2�Y�?��? #`������'�������ɽ[�>_1�J}����g\B�1��:�;��cf�?��?�
C���6�!������l묾�@?���>Qd�>"I�>E)���g�r&�A?>Zi�>�JS?r�>�&W?�7v?eW?!\0>߲<���^ό�x��=I4>�g-?m�o? �?NGq?1?(�(>�g5�G���� ���>����M}��q<�mr>Yi�>��>ӕ>�=�)���S���6F=��m>n*�>��u>���>��h>���<R�G?�(�>c���<6�-9���k����<��[u?�g�?+�+?�=�����E��@��@l�>ZB�?~ë?s�)?�T�2��=��ܼ�궾=�o��¶>�]�>��>���=t�J=�>��>�3�>+��sR�=`8�=gM�{?�F?�ֽ=n�ÿB"G��Ծ�~Ӿ]�F>j*�����oL=t	��bh1�f.���� >ł0��|�l�L��)˾�2��mI��.�-�	�?O�>̔;��=+�P�H>�Hh�;7��>*����\�=��b=�1������T��ȼo&2���=<$=�����ɸ�!͑?��j?Ck>?��E?K���EV=����k�M="[#�J�.?�|=��z�|sپ�i%��4���0��?8��hf׾��M�<͵�Ȣt>��f�?yh> e=��!=?�̽�\�=�J=I�=k���D�=펡=3�1���T������=">�~?����ɑ�Nn4���W�v�9?ؾ�>ǅD��;o�.*J?�+�>�W}�2����_�ѱy?y��?���?�?7y�Ǽ�>HE��	���@p�=(	L���>��=�XD��V�>��>s�or�����Q�?}Z @D�>?�����Ŀ��.>��">�>5�T��2��P��w[�fd���#?q�>�!�Ͼ�N�>���=��ؾ4�ľU5=2�&>�IX=�}�iY��İ=�g���.L=b�a=Dw>�9;>Ȑ�=���=�=���=_,3>�c���ގ�;�J�RXd=���=4GW>��>���>8�?��0?Vd?`��>�do�,�Ӿ6尾nF�>�$�=�>���<��
>���>�0?eUA?�JK?t8�>�Y�<<��>���>M�5���j��׾�З�=f�=G`�?춌?�j�>�ڃ=ż&���xw5��b佯�?�1?�~?h�>�T���\&�r�.��0��*@�7Z�*=Mhr��U��= �@��	A��:�=Xq�>���>Tҟ>"6y>��9>#�N>3�>I�>~�<@�=������<qԕ�e�=Uݒ�Fk�<w�ļQ�Y����T�+�vd����;.��;?F^<~��;2��=�?=5�>q?�ط��<޾��0=a3t� �a�C���"EX�׵T���~�������������>>5�>�H��u|��W ?�>a�5>ռ?ÖS?�;+<�#.��ƾ�m��0�%�!�&X >A�/>�G����C�F	X��tQ��έ�X��>�Ҏ>��>�l>.�+��?�V�x=i��tB5��>�^��������/q��9��	쟿Oi�r�ۺ��D?_8��p�=((~?��I?�?�f�>�j���yؾ�,0>�"��m%=
��NXq��c���?,'?��>��?�D�܀Ⱦ1P���1�>l�D�lO�\ ����.�+*�������>`�����;�1�$���0���/�A��,t��>��P?���?��f�S���L��s�[���Ⱥ?re?�>�?[�?@���&������$H�=�Dm?�2�?���?��>~��=8A��j��>N�?��?&��?�s?}�@����>��'<K� >򺕽���=M>>sڟ=���=z�?M$	?}n
?����i	�C���#s[����<{Ƣ=�^�>�E�>�:t>H�=��c=���=��\>�>�>��>�Ne>`O�>[�>������q�%?�n�=c�>��1?�=�>
�i=S⭽��<��F���>�c)(�
��NK��O�<N'��*zL=DͼV.�>�-ǿh̖?x�X>���A?�����'�^R>�Q>�ܽ��>��D>�!y>zǪ>�?�>U�>)Ë>��)>ӚǾ/i�=.N���$��%�@�-�q�þ�%�>:��p�1��V�5y��2�YA������
}X�ms���6���j<Y9�?� [��&U�f ��� �F^?̄�>��?�󙾀]+���I>�?��>S�˾a����l������6�?<P�?ۚa>��>WLX?�r?�94�J�5��Z�'s��]B�Aze�Nt^����U����<���9^?o�w?G�A?v#�;e�p>���?�(�5���=�>��+�.97���\=d��>����i�Q�zDϾ��¾�+��;>��m?���?�w?E�Q���e�� '>��9?%90?�
t?�d2?9�;?�e�m{%?��:>YJ?7?1�4?�t/?�2?�4>" �=v_���#=���䋾0jԽ#�ν�����2=��}=,�0:�<{ =��<������w�;V����(�<T�<=\ݞ=�X�=e:�>�`?�Z�>�.�>F:3?'�$�4�$���v"-?�F?=:lo����Y^���*�����=K�h?o��?�Y?�OP>i�B���B���>,;�>\#>O�P>���>�T �0<�餖=4^>�>+ҭ={�%��~����������< �%>G��>�s}>yu���9#>�����w���a>�J�����xJ��F�ߏ1�<�p��a�>��K?�i?k�=^�龙?�d�;'?�;?	�O?<{?�ϑ=��۾	V7�&�J�<�%��}�>�<�
���� �����:� ���<~>�����Ԡ��db>{&��Tݾ�n�лI�X��XK=J��"U=��~�վ��~�!�=�q	>	���� �U�������J?��h=N褾8�T��纾��>�X�>lӮ>E6���p��@�X���r��=:�>)Z:>#����XG����O��>JD?3�`?sĄ?�|���.r���A��\��`%����g��U?An�>N�?E�<>�D�=�;���-���c�~F� �>���>"L��{G�G0��}����>&�`�>�?��.>�:?�1P?X	?�4]?�&? *?P��>Xv������C&?<��?��=i�Խ;�T���8�D"F�q�>z�)?�cB�З>|�?2�?��&?~sQ?ƪ?h�>$� �!.@�o��>Q�>O�W�^��f�_>��J?���>98Y?kЃ?g�=>̈́5�DѢ�z��G*�=�'>��2?�0#?g�?3��>6#�>U����q�=��>��b?m�?�wo?���=��?��.>�J�>v�=kd�>;i�>o1?�iN?�?s?y�J?`��>�<����I��mQ`��)����;��}<��|=U��opr�'����<�L<J����V���׼��G������<���>4x>�f��H�2>�;����/X->%� ������8t�MK/����=;s�>�y?���>���Us_=�b�>(��>����#?�f?h?���;��c��˾��q�>��=?x�=��i�[ї��Xn�-ע=�o?2Z?C<r�`%�e]?�\Y?��뾙����G�1��'(���`?چI?�6=|Z�>T��?TA�?�B�>z2x�!bR�rʒ�2{.��q��b)=V�*>�X���&�U,'>�ð>��>�U>��9��!�oo��8����>~?@d�?�Bs?mzq>��^���ؿ"z��]�����^?I�>B���f#?.�<X׾*롾�̌�w�پ=Х�zB��B���图���D���COɽ���=�,?�;x?j�i?��_?�$�f�a�|VZ�^��Q�'��A���eG��3?��C�Fp�������v���c\=il�2�,�@�?��7?w!�X��>���&㾪��X	>/+��.'ƽ��M��7�	��=��=�O6���
�$���?k��>&��>�|Q?�i��2�����J��߾�3�>��b>ck,>��>��|z���/��x���������V>��^?�M?�Xp?�d��s�#���z�f;"��k�������S>��=�Cn>�xL�8y/�u&�i�6�!)k�M��˅�n�ȇ�=p2?�1>p(�>"�?\M?�G�������j�fx1�u�h<���>��a?�G�>���>h�,�\����>��l?��>���>	񌾬� ��5|��Ľ7��>z��>�r�>�s>\i'��m[��H���C���L9�
��=��h?$����`�%�>FmQ??*�9�B< |�>ls�e!����fi)�v>1?as�=��<>��ľ ���m{�H���P?��>������N�nh?e?�/?��?�yi?���>)� �/�`�(?��t?@L_?��2?���>$�ʾ������Ͻ��,���:=Q^�>�J!>���<{��=y�=A����@��t�;�����[���~���0>��Y�4?����=���=w�P�N��᪾x�꾛��,�UDϾ�+��5��7�)���)�b�Iqe����U��<���|��0�(ㅾ��?��@Qؾ��ξ?���bh��Z�]�X��>8�I��h���A��\���3��׾�Z6��uj�G�}�*�p��?,����{ʿ�Ь��!5�UbB?�G?=�t?~����"<��N�Y��>,�>>�ˊ=o�噿�9¿�����}?�m�>"u��+���F�>��/>���>�+>.Y&�!�N�n�2�Vϧ>!pS?\��>x�Y�Q�׿����n����4�?4X@�@?ͤ'�U�OL=' �>b�?�B>�,�����Ʊ��K�>��?�-�?�nL=�]X�z&���b?1<sYC����3��=G��=:�=*j���I>>��>�^��@�@C۽8m9>���>�%*�����\�~��<��c>R�ؽI���{ӄ?�l\�ٟe��V/�"���P�>�T?_=�>X�=f-?�9H��Ͽ`]��s`?/�?���?y)?�U���>M�ܾ%�M?�x6?���>��&�u�C��=�(��L�ZV�h��=d��>>�>ʨ+��p��9Q�쑛����=,���ƿ:�$�os��M=�ֺ=�[����r�1�T����xZo��i�v6i=�#�=ܞQ>~k�>�2W>�2Z>8nW?x�k?�%�>C[>�4体����Aξ��N��� �Q������棾�|��߾�	�G�������ɾC���=�\K���������=p���f���)?�>$,ʾ�(7�z��<����5�ɾnk��ij�@V߾�93��Tj��/�?}#A?�(�� /��Ä�}V��m����v?p��R���ÿ��t=�O��wǼ<R�> �=7jݾ#1��c<��L0?��?�>¾����a��=O20���A�.?�?��l=��>��&?���'�^�]�m>Ǽ+>�G�>@v�>��=�
��V���&?�XV?���I��z�>[ѾІ��+w=E�=�H�7佯�>���=�<U�zD��BG潞����V?j&�>X�����׺��n��3Ҽ z?W�?��>9sq?]TO?cU�=�پe�T�9
�}���AT?��l?��>�z��?��4���\)+?�b?ߛ%>�bC���Ҿg�7���L???b�?�y�<�Ej��d��p����-?ѝ�?��o��@������߃���>d�>1��>�]@�:��>� d?F�e��ޟ�Epÿ�K�篡?|�@�� @�+�Q�?�/E>���>�]�>:_�{���7LL��̾">��=?T7ɾ�����J��}ӹ?�e?44�?Z:?Z�������f�=��N����?���?ކž��=��׾p�x��&��a,�+>�i���罤R��G$��c���	�Y���҇��_K>8�@�Z޽�>�E��!տ$�ɿ*fy�9�|�����%�?�e>_�罺���=v�h�n��E�H<���Y��sv>f�>*a0�Ӿ��W�<@��V�P�?>��3>,�S�h���׈��Ƣ���>�J�>�[ >�2"�I:���?m���ܿ����j����u?���?r�?&?@ï��nɾ����tM=;�Z?��o?� 9?�D�#YQ���=Nj?�����`��`5��C��0\>	L2?*��>�a,��h=��>r��>ڸ>k�.��~Ŀ1���R���X�?���?�~�;��>jB�?=�*?f������*��5E+�
�4A?+�1>R���3"�=��k��=�
?�t0?�7�?���_?J�a���p���-�N�ƽ�ۡ>V�0�[\�-\��t��8Xe����*Ay�F��?�]�?��?���Z#�Z5%?��>�����9Ǿ"
�<�~�>�*�>G/N>�L_�r�u>����:�gl	>��?z~�?3h?~��������Y>��}?��>��~?��=��>���<k쾒[�/b >@`>��)=Y��>(�K?|9�>��F>滟�����cA�x�P�W�)�E��D�>?Ʌ?��U?1�f>�(Ž�4�<�l;�P�����~�A�K���T�\(��e&>�8P>3/&>�*k�r��|�?'����˿t����V�׽E?D\�>ӏ�>�x�o8ž�OK��]y?��>���x޳��t���RZ�/�?I[�?��?*���"F�=T�='ʚ>O}>X�Ƚ"y������,>�5?°۽̑��0v�{ix>��?o��?���?�rN�X� ?�v��m���L��v ���Q�H)�>v-?���E��=��?�j�> sb�!յ���o�|��>��?�3�?Ү�>m`j?�����'�e>�\]>5�i?��>;Qs�9���
�>	�:?���T+��[��.�r?��
@��@��?�����������R��ܶ��=�=X��=�s= ������=V�=�6ƽ�;齈,!>���>�>٬�>�`>vwh>�{F>�T��R)��@��vR�����@� �����?��s�B����;��߉�����4��=�ػ�b���� �,=�;1�=�^N?��`?��u?�͐>m�7�G�/>b���W>�u�;�P�=S/�>ΐ?d�=?��?��=8���h�Q�_Rv��&��>X��3?$]�>:��>�D�>���>���3�e>���=�P>��=	X ������5����>ɷ>?2�>M��>o:>�q
>���Ô��z�H�� U�Gμ)h�?0�_fJ�b-��옥��p��=��=��6?1�=஋�~̿wॿE?�K��M��������=�^;?��]?�>�8���XϽj>Z�ڽe�[���V>��=��^�ۼ+�ѳs>m_(?B�f>�dG>�?�?�8��h8�QQ���>�>�V?R��f�X��VX��<b�c������>��>�8=������ew�'vZ�l/=�*?�?����h����R�j���>DM>2�E>�>k�>��6=Oi��SA��Bz�&{>3S�>��?��+>l�=R]�>}�����O�C+�>x�A>�!,>�j??P�$?�������/��Ө-���t>�=�>��~>9*>حH��f�=SH�>#.c>�B�C}���(�1@��>Z>�r��cc���v���x=}���=�/�=b
��e<��4)=��~?���&䈿�뾎b���lD?F+?� �=��F<��"�A ��H��>�?_�@�l�?��	��V�"�?�@�?<
��¶�=�|�>׫>Bξ�L��?a�ŽjƢ�z�	��'#�ZS�?��?Z�/�/ʋ��l�L7>�^%?d�Ӿ�n�>�
�B���z� l�ݛ���j�>��H?���,����D��?{�?t��9�����ſ޽k����>0��?���?w�n�Ɲ���:�� ?O�?��R?�.>�� �����>�B?�k;?�C>�����LC?o�?�Ƅ?��=x5�?'�t?�5�>g  ��?B�='��?���3���b������>.��=�dȾO�^�#t���#x�z�I�"'�T��=}~�<���>����������c>Y�T�-�-'���M?�ȍ>%s8>RJ�>�g?�Ȯ>}>�{��@i=�J���!�!K?���?���fcm�`��<���=�:X���?) 5?h����ξ���>�\?X8�?��Z?��>x}�`���������#.�<r�W>@��>�R�>�;���M>�$Ծd\J��(�>u?�>�ӼJݾ�.~��L�;�h�>�Y ?_�>��=[�?ˊ.?t�>���>�0Q����lOa�B��>7s'?\}?C��?��>-FL����<���T,��͝Y�x,�>q�n?��?�>ۘ��\��yo&>�A>�󽫶y?6�h?Ճ��H?敐?ƴN?9?m�L>gD�,���d=���>�?�å���b�%<X�J}5>���>�B??DL?7��=C���v�@�J�)�>뮾�8?�3R?$?4����s���8�	Jм��=܄�������P�<�4D=�a�=��=¢ʽ*�=y)"=�����lu�)J=e1>^Ϭ>g~�=�:���<���1?�|���/(=R
>G����g���M>-�;���	�iw?ݾ�0��;�����\*�>���?*��?G��?T�ɽ�\���4?z��?�E�>y�?��{(���rپ�.޾k�ľ���o�=�t�>ɒϽ]F���䫿�T���@@���:��a����>t��>5�?�[�>�fW>��>�ǝ���3�D.�M$�c�J�X*���1�j��R��=���O׽��\�������>%Zս��>�v!?e�>���>N�>�:����>��>A�>Uv�>c/Y>a[�=C��=�d==���7<?~���?�^����-��\?�bM?џ�>B��<�v��i�WH'?��?mk�?'�%=�e�4����>��3?�t�4?�>��'������pC�M¾��=k4�<O�>'^�>
@>�� ��D@�����`�?�{?��>6�(����6��E>�ϊ?�,D?0�L�]GB�!�O�)�F�z%����=�-�m;����'F_��ᆿY�b��g��[���m�	"?O\�?���s��Y�y�%�x�a�\����>��	?�v�>p}�>B�	>���W'��}[�J��C���
?C\z?ea�>�#I?�O>?(�Q?$�D?u��>�k�>L$��%> ?���<���>)�>�6?v�-?��/?�9?c'?zCV>f�	�V����ҾP�?�?:>?��?�?�������������u[s������S�=�1�<!Ͻ}�?�Ρ=�U>^X
?U��{a��wB��t?��?>uH>)q�%�q��D�t;��W�>�e�>>>�t:�P�c'�}�.?s��?�/��y=�{c>�S>��=��Ƚ�˂=A�=�wٽA�����U�?fY>6>�~=^���b�Y�zy��s4�oj�>(�?���>@g�>v��i� �B���?�=!3Y>2�S>�*>�Rپ�s�������g��Gy>Ee�?�l�?�f=Qw�=W&�=䪠����&�����A��<q�?SJ#?bcT?U��?׾=?eX#?��>�&��>��lZ��GǢ�J�?Ö?C`]>������<+����5���4?"�A?��M�������ȏ��mܼ�j�>]� ��>e��N��'F�:O�ľ� ����?��?1M���E�����퓿��M�>�?p�4>:9?l�=?��f�1&���&H�{jf>T\?s�h?��>Q�O?�,{?Š[?y�T>
�8��.���Ù�,+'�o�!>41@? ��?�ݎ?��x?��>�q>5�)�8��\�����6v�������W=`%Z>t��>���>�˩>�~�=ɽ�>��ӵ>�}��=� c>}�>]��>���>6tw>�ޫ<M�G?���>�^��q���ꤾ"Ń���<�ʝu?w��?h�+?LM=�����E�F���K�>o�?m��?�2*?M�S����=�ּ�ᶾ��q�$�>�ڹ>�1�>�ȓ=�eF=<`>M�>���>n+��`�~q8�aOM���?�F?���=�Eſ�gp�(Xi����(*<"���c�A����Y�.d�=�E���e��Ԩ�-�Y�꟠��ד����"ӝ�H`~����>e�=��=��=��<���d0�<b�L=秼<F%=������_<�2�]��a���>#��?<l�L=<͞� 齾��c?��[?�fO?Ov�>�ɹ�B�=*þ��V>�[<�z�8?M�b=t.ӽ�����ľ0�þ��
����{�6
�cm��W3)>?Z�=Ц4��>iSx>�n�=ǝo=��= ����ȼPPd=ԇ>��>�o�=`g�=�t�=�ɘ<dz}?�~�3���l1�:LV�rw0?�S�>#�<�c־�\^?28X>fR���cɿj�V��?W�@:��?�S?��O�9�b>K�J�Yt�=8�z<�h�;��=��@=/�����>��>\Q�2��2}̽)��?�� @0�f?����H�׿�3>��7>�>1�R�M�1�#�W�<-`���T�1"?H�:�S�˾T��>v�=�߾�}ľwD>=dH6>#pe=)��j\� �=��~���>=9_s=~K�>��D>»=�^��[�=�A=��=E�M>�����0�hN)��}:=g+�=Yc>��%>�t�>��?��0?�kd?���>��n��-Ͼr,���m�>}6�=�!�>_Ԅ=�SB>+N�>E�7?�D?�K?F�>U�=-+�>J/�>�,�c�m�u0徉��w�<銈?�Ɔ?�f�>r@]<�zA����P>���Ž�l?{1?ۑ?�=�>Ԅ�n���$�Oj2�.���h��=1<Ok��yܽ!�=$��4����I$>Y��>p?~��>��>��^>��r>��>L>�K�o(ϼ��<T>
��=�<v�7�Z�<��>}�c=�"��Dw�TD�5�j=��=��=�ʜ���=B'�>��>m�>�m�=�Nپ��#>i�Ѿ�j_��+>Q����KA�>�y�j����U
�SVսGh>�_w>j�����U��>\l�=!��=�l�?l�?sl;>5��;֦������P�W��5�;̸�=�܀>ơ����_��tt���K�'@����>wَ>�>�l>�,��$?��]x=����^5����>�~����a��?/q�?�����Ni���Ǻ��D?�9���>�=N'~?~�I?ߏ?��>ޘ���ؾF�/>�U����=D���>q�I0����?�'?���>~쾍�D��T˾lQ��K��>!iF��CP�wÕ�v~0��V�������>�z��z�о<�2�ZF��� ���CB���r�9��>^XO?Pɮ?�`�KH��)�O��"�Q䇽X�?�"g?���>��?��?������� ƀ�4�=Q�n?�)�?;�?��>�i�=�k��B��>B8?���?)��?m�r?��=��m�>��e:+�>)ϕ�fv�=+V>���=P��=ژ?�
?T
?S�
��ﾧ�ﾰ�`�M�=Ǫ=&M�>�-�>,�q>��=_[v=�z�=�`>�p�>��>�[e>�@�>���>�-��x$���+?�p>�$�>��1?8�>���=��� 7�J��G�&�_U�~p��됽�m�<鯃<ǎ�=��� ��>�!����?��>�c�/1?��Ӿ�e��� >ZxW>�ӽ� �>CE]>�d>#��>��>� �=jˆ>,�,>	;��>���Y)��8��{M��?ƾ��>-���|�:�W����^�;��~������ui�iڀ�3L=����<���?x��R�m�GR+�ST���?S�>.Z.?B��U����I�=���>��>�+�^T���q���;ݾ�i�?ޖ�?#�b>�R�>��W?b�?�2�
�2�>Z�s�u��FA���d��p`��Ս������
�yL����_?�x?�\A?�ō<K�y>��?��%�����-�>�./�vP;�{I==���>*���QN`�ÜӾ��þ`P��jE>cGo?	�?�???�U�����8�o>�rW?�$P?Q^?!9?YT%?�|�B�>?���=/|?��?�4?2�U?��?�la>�[>E��<W>��oQ������^ٲ�K�����s<)X�=�ڔ=;K<f�#=� J<^��=��^=�~H<H��
���<?=$^�=�Ł=��%>m��>��]?�\�>R��>��7?����y8�9ծ��/?˘8=������9Ѣ������>q�j?��?�SZ?B�c>�A��C�I+>\�>N&&>K\>y}�>]0�P�E�+K�=�>(e>��=!M�V���[�	�U�����<�>2��>ͤ�>��a���5>�����>����S>+zT�(�8�ZNB��N)�dc� �>��L?ѿ?��y=A��]fĽ6Df�:�(?H?H?�:O?Y){?�إ=��;[�?��H�������>�C6<��$w���1��Ȅ7��Y9<�l>:	�������>�������{j��|C��I��F�=��^\>���Fv޾�����S�=@�2>�\��J������覿�H?f�R=_�׾-�Q��D����>j��>�X�>�ˆ��ŽǷQ�Y���%�	=J�>��>9���{���J�E�����>OaC?f?���?�J����h���K�K�D����#ϽJT?�l�>w�?�O<>`Mc=��������[]�ăF����>@��>�[�~�C��2��l���7#�<u�>��	?�>X@?w^L?�?�Y?�*!?��>��>l�ɽ����.@&?Q��?���=o�Խ�T���8��F�x��>P�)?ζB�b��>�?��?��&?z�Q?��?��>&� �BA@�2��>Y�>.�W��`����_>��J?���>$9Y?�ԃ?��=>75��袾�ͩ��m�=s>��2?J7#?:�?���>��>Ĭ���o�=e��>��b?�/�?��o?�_�=��?@j2>@��>Aۖ=4��>ŏ�> ?�NO?��s?x�J?x�>@׍<�Z��D;���|s��O����;χH<�z=G����s�H{�0�<ҷ;�g�������̲D�{f���0�;�/�>qR�>�ॾ��>���������Ob>�^<�����,��c�F�>��=꫃>�-�>I�>����ڮ=y+�>�i�>���.�'?���>��?�����d���ɾ�Z�m|�>�eK?�7>E&p��(����k�OO�=�f?�v`?�K����ʲW?��I?��ھH�_��Q̽+�Y�@�l�:g1?�?��8����=P�}?�P�?cy?_�ƾ��B�#���Se���<R|>Oh5>���c�;��7�=�%?�p�>`��>|��>ÿ]�Y�o���پ.��>�
`?���?�̨?�&�>�(��������Q��`m^?1k�>W7��`;#?�A���о�D1��r������誾ӷ�������@#��߃��Lս��='�?��r?a�p?�_?�$d�-�]�#��IV��b������D�u�D���C��mn�^%��@�����!==�۽��K��Ϻ?�I?����P?�aɾ�{ƾ8���#�?@鏾�!-�䊯=O=P<h>p	W=��*��[�'�����?<��>'�u> n!?�5b�5�8�d�0��N2����ٲ�=��{>��>��c>^�;�ܗ���l�L���l���a��q�u>g%^?��Q?��p?O�(�R�-����0�%�5q�?;����t>7*>Sm�>��#����C��3';��Tv�2���n��-����=6?�Im>�ۮ>&��?Ǳ ?���!m������!4�0������>�8g?��>��>CX��������>�Nl?���>���>ҋ��m��T�w�k7�1��>=�>��>*�n>�&���V�я�׏�4�:�ح>��j?0 ���b�ڊ�>N?�G�z�;;�ݦ>/�
����N�N$� L>�]
?p�=WL:>�5����҅}��#���b,?̣?Ae��Ҩ*�S>�)?���>��>}�?���>�P޾�G���?�^`?�=N?�G?<�>�Ƽ��ZWƽ\�B�Q��;K�>ȄD>%�={��=A��C�&<����;mJc=L䕽�����V'=(������<M=�>"ڿ��F��*ݾߥ�T"�{���z��l��H��{���赾A����)t�¹��"8��qO�$JS����2Mg�y�?�o�?�e��B̏����c��F����}�>�is�
(�*������a��nNܾG��������H�Y�e��Tf�#�?�=z��ֿp�����依��>Pf?��?ʾ:>@�%�p��v>�)�=��=�'���2����ο�k����/?��>��
>O¯>�[>�Q7>�B=2Ƚ}Ǿ�-a��N*?�??kXB?�&n���ʖ��|�=���?��@dt>?���\ﾸ�����>r?E�F>��F1�.,۾���>��?�?""9�P�T�W��ӯ[?:�={)�����>�+>"���S�%�a>��[> ���|w�����z6>��?>NOQ��*b����G
��j�Z>`u���v��]�?�E]��s�h+�i9^�]v�>DG?z��><"�>	?la}�Vӿ]�G�v`X?s��?��?a4>?���B+=ď�g�A?�$?yZ�>���z�����
�=[G���վ\�>���=s(>눓��0��c����s=0b�=|�	�����  �H޾d�<�=G8�=&׎=xt?=gt>
�J��ρ����	Ab>��U>���>��>M�>.?�=+;r?Q�?O�&>u/�x�޼��,��b��4�D=�D\���$��a+��-C=zĄ��\ɾ#Sʾc�:P�i�ƕپ�<����=U�V�+U�����T#[��.���-?��;>����=�I�U�5<��¾����6R���u��R��}l)��f���?@G>?�;��S��7�'_����K���J?/�	A�,R��ePu=Ï���5=S��>���=@�ξ�/��uZ��+?bC?hqܾy�q����=�xƽ+P��sS?��?�S��ݫ�>���>ؠ�,�M�<ӛ>�+�>��N>�	�>�s�<�N������?&�?�R"����GV�>d���}�ѾR�oJ?>c���-��W��>��;������(���ԃ< ��<��V?g��>*�)�����~������*:=d�u?ͨ?֪�>�-j?��B?;�<z3���}T������c=(�X?�/j?,�>��4�Ͼ�M��A8?�$c?�pL>��n��i�,�H��:K?{�l?d�?i_����|��x���N�o�5?��v?�,^��V��ܾ�L�V�>u��>	��>N�9�f/�>��>?�A#��Q���ſ�$4����?2�@��?x�<<$ ����=e7?[�>YP�S6ƾ���ɀ����p=8(�>�O���dv����8/,���8?ٖ�?:��>�T��ʥ�ݫ>�m��)U�?�,�?H���(׌=-*�>kn�����4�<��$>D10=4�K=�I־(l�HX���a���`��)>��@�sl�O��>��mݿ�ǿ�o�&㗾�����"?�x�>��/��ా��e�1r��VE���Z�W��S��>E�N>>�����Ⱦ�6H�R���MS>���>%dG>#��>�խ�4�ξ��%�(r�=���>��?���>?���}�1��?(���Zҿv�e�F�9�\?#�?N�W?Z�(?���\/Ⱦ��%����8?b�?�V?��>�,��ě�';i?�����]���9�Y=�ڥj>�~0?:��>��3�L_/=�>� ?�!!>��2�E�¿e��������?�'�?hS��F�>\|�?W�$?���.ȗ��K��T~/����B?��.>ryǾ�D���<�>��;?�c,?$����L�_?��a� �p���-�D�ƽTԡ>Ћ0�H\�V{��?��_e����jMy�;�?�\�?��?���D#�+%?��>�����GǾ���<��>_"�>E:N>��^���u>l�R�:�=|	>��?�z�?�f?���o����[>�}?G��>�܄?$��=0i�>Ê�=˰��r��/>�3�==�Z�Se?/9N?-�>(��=��:���.���F���Q��A�z<C���>��`?0�J?�g>:?����N�o� ��Uɽ��4�}�0�<�:�5�	�ܽ��1>��<>��>aF��Ѿ3?���M0Ͽ�>��y6ϽqY>?�W�>Y?X�+.ξ��<�i}?#��>g�@��gv����ڽ�Ҥ? /�?N�?�������=IݽoF?Ь�>h�W��!Q��ھ�<v>��E?A�.������t�t�>r-�?ƹ�?]��? N��	?����=��W/~��w���7�e��=��7?��Jkz>m��>��=�hv�Oê��s�ç�>M>�?�n�?��>D�l?�Qo��B��2=�O�>�vk?�W?)jp�����hB>��?��� ���lO�)f?��
@�q@��^?R䢿�/ӿ{�������G�����=�!�=��5>'9��0g={�=Ɲ�<��j��6�=���>uv>S�q>�Ď>�E>�@)>"���8�)�)�������PB=�YK��v
���L����@OP�O��~Qվv@��
c��������9y�1�*�T��=q�8?��j?�Wz?��>��#;1��;y�aá=u�M�X�4>"~�>`�??WO?�8?�>A$���6]����jɘ�Ĵ��L�>�B>���>�?��>fW�=��(>*ؙ>��>�0]��N�=+rY=��=>��=�?�>�>�٧>(�>�Rb>F彿�Ĥ��`�f��ؐ>���?
T!��	5������u��u�˾���=��A?m*>�쌿��ÿ����H?0�¾�5��ϻ��E>��?�-Y?x��>Es���l��ށ��[�f���0<>�"���h��:U��Q>��?��{>7X>w5��7�i�B��2���SG>�A?`W��]��_s���P���辐�>8�>̌�=�m�͘����=3���G�=��7?il?� ݽ���-����P�7+,>�5b>pT>���=�+E>����L;Ͻ� ܽ���R"%>=�>`�? s(>�L�=���>���g��F�>V?>�u>x5E?>N%?�(��md��R��H�:��e>*G�>�s>�	>_&?�S��=�]�>�$V>{��4j~�<��B��^>�m����X�Z�*�'<=8��E�>�=�=���$�!�O=�~?~��䈿��jb���lD?N+?��=#�F<��"�4 ���H��&�?j�@�l�?؂	��V�W�?�@�?�����=�|�>�֫>�ξ��L��?��ŽǢ���	�)#�ZS�?��?&�/�Gʋ�l�16>�^%?�Ӿ,��>Y`(��X��1���pk��J�<:.�>:a?�{ھ����uF\�A?	61?=H�'Ʋ�`����j�̔�>���?��?
X��0N� u�ʽ$?��?p$�>X�=g2
��l�}�>P0D?]7?��,>����@�(D+?mð? ώ?��>>���?W�{?j.�>]7�_�&��[������*5n=v�U�ʿ�>�u�> ��D(��u��\^q���s��v�:��=��<Ѹ�>�3 ����̘>P8�:�Ҿ�޽>��>�+�>�>r��>���>y��>�1�>^w�=�RY�fx�,���K?및?����0n��i�<}��=I�^�D+?�N4?�bZ���Ͼ���>{�\?���?x[? y�>%��S?���濿�~�����<ĻK>�>�>�:�>���9K>:�Ծ�/D��f�>}ח>GW���@ھ�0��aC��GM�>�]!?%��>mή=�%?�&?`�h>'��>P0������L4�-r�>�ϫ>D�?	zf?�-?/�����%�h;��nv����U�sdD>�{{?3�?�=�>�"|�����j�<�D���� � S�?Pl?l�d�}?�?n^+?e<?��>O������g�[�j>��%?��,�F�Z5&�����F7?b?R��>0��<1���ֽs3(��\޾�?O1a?�|6?e�޾�In��T�>C�<�i���f��Y�=#;��a3>�>�=v���==��8=SD��ܗs��U¼ �>��>�]�=��7����*?���=��\>��r�D��r"=�oW>� ��T,?��=�Ѓ�@T��"a�����o-�?:��?�ݓ?D�̽B1d��>�>��?�,?�>��B��Rƾ�Ӵ��kླ�`�q�:��/�=g�>�q>o�ﾤ��M��������#������>ʌ�>B�?7^�>E�Y>n�>Yp���c��;�(N���X�ǐ��-�#�����O(�����y�2��%ξn�P�#8k>�$�U	�>�m"?d�>�Y>@��>2<S��>0��>	֢>uz�>��Z>C�>̽�=�� <���|DM?+��RU� ���
7�16?�^?�4�>X���{�$���F?y��?~��?_y�=��~�#<9��?��?�.��0�>tj�<߸��{/��r�ɾ��O��s�=g�!=�'�>á��t���# �ֽ�����>�/?�%���������s�U
=Hqt?�}+?[�@���k��_h��h?���Y�.�Q>�^��<�׾(�j�ؓ��+���
n�Q�-�"Y�=�>$?��{?Yԍ��_�U���0&R��B/�PK�=OQ�>?τ>H��>"�>$��s>�IyJ�t-��v8�N� ?��|?���>`*G? �=?�Q?�*F?�"�>�0�>[1���|�>��4<��>��>�84?h{,?`�0?4J?i{)?	y\>��)�����پ��?8?Ʌ?Q?��?[3y��R��o^��y��.n����C�=@%�<��^�b����=�dX>h�?NJ�>?��4�u��&�?.fG?�.j>1��:�F����D"��c�>~U�>���=e�b�}����5��~?z¥?�۽�iJ==�=:i4>U�+>y���W>���[�Z>s�_=2j½9Lc�&<�7A�>��t�/�����e�=<�Eb=�w�>��?ɖ�>�J�>YC��� �̺�qb�=pY>sS>=>>sIپ����&����g��cy>�{�?az�?4�f=��=��=Wu��PU���������Su�<@�?VC#?fUT?���?�=?�c#?l�>R%�I��eY���	��U�?#�?;�h>Z���C$������bN����>�?W�o��9���8��5�8{ǽ�	�=���gXO�����aI��:���I��"��%�?���?�|h��bU����ٖ���r��&kn?-��>�ǽ>��D?��AV��ems�ز�>�p�>J�c?1U�>��9?W�?l�h?����ͥ� ��������X)>s�>23R?|x�?��q?��t?���>�Gk>��W�;{�)b'�w1k���o�G�9�>��">�"�>�>
`�>��< ?�=�P��G���8�<=�V�>��>�ʇ>�B�>��>�s��C?{��>�;(L��ߓ�z��Z���?2�?�8#?!�=)g+���F����$C�>gQ�?wq�?*�>�_��`+=��;���d�]�B/_>~�>�M�>��5>X��<��=��?�ܝ>�VL�
�Y�!�I+�=���>+P?��=;��<+J�2z��J?r���R�y�����=�i6>JaO�ƚ�VվkwQ��$:�c���𭾧SC��T����`������?��>�%4�q�m�+=@ Ľ��>S"+=�r�=�<=�X��p�=Һ�<-h]��}b�x��=���=�vK=�n�=�忾V z?;�L?�.?�O4?�d^>lo�=�֮����>>�٦?�H�>�t����z;O�>����r����ھ��پ�d�����d>��m���9>��>�lJ=�.�0R >WAS=�N|==<��=��=�/�=�T�=���=X�=T�>I6w?u�������4Q��T�ѷ:?^<�>�=�vƾ�@?�>>3�������^�-.?���?�T�?x�?�i�~d�>	��h��j��==��E2>��=��2����>�J>_��6K��?���2�?F�@̝??���	�Ͽ_M/>��3>�o>�R��'1���[�^a�G�U���!?k�9�H˾A��>�g�=�ݾRkƾ�c,=K�7>-(e=0���n[�p�=�p��d)=��g=*%�>N@>�K�=����Ѷ=iwY=
��=�PK>������7�"��7=�9�=	\b>�!>�� ?��?)?g?i��>��侵�������Y{>B��Vw�> J3=��v=@�=��.?V�-?cU?��>
U�=#�>�/�>�q��jJ�g@������<�1um?)�?�~�>X>6ꎾOz1�EH:���=�)?�T?��'?�Z>��	��׿����"�羇������=��&>䡼<�cֻS�>=z)轔4)��~ѽq�>!�>���>;�P>M@�=���<ɍ�>r>k�E��?>k����=��>y>�N�=����^��
<���=�������<`���꨽� �=��=��
>��>#-�>6?�����{��U��Θ��^b�)69=mm��R�U��s�,x�o��ʨн��>��`>qy��DB��\��>Vg)>�T�=���?�N�?���>9���A�뽯�����Ǿ$��+@�=���>{y3��3"��xS���S�{����_�>���>�V�>�r>)$-��5B�W�G=��߾�q5�aQ�>�'������Y���q�������'�e����ND?;愿��=��{?�qG?�B�?D�>R���Ѿ��:>����=«�u����?�U'?5��>ǭپ��@�d豾ᓽ��>dA���N�{,��{L4�1��8�ø�>�땾�����*�cC�������D��Y�>��>��L?�i�?��%��v�[�=�E ۾�.���M�>Z�c?�Ю>h��>��	?,������w��<+>w�s?��?a$�?�g�=�P�=�y��0\�>�?��?���?Qp?��K����>S4>;�>�����!�=�|>��=4/�=�s?�y
?��
?�o��=p�h�ﾺ���d�-��<A�=�b�>r�>ow>��=8��=y��=�L]>��>6ڍ>�_a>k��> �>�����
�	>4?wB>CKI>(E?��\>�뻍%���>�ރ<t%=� ʽo`�<���>�=�p�=��=A�P���>U�ѿ�A�?oD�>;&���?1k��JC��H=!Н>J1۽~�>��>}gM>r�>3��>M~�=7&�>$2>�BҾ%�>����_ �cC�Z$S���Ѿ��z>V����& ����R���E�W���{����i������S=��8�<���?j�����i�#*�IV��?Q��>w�4?����L!���>s�>s�>e�������ߍ��ྋ�?��?�Vu>��>L U?�?��1��;h�}j^���k�7@=��Cd��Q�����w*����ׇ��V?3�v?�I@?�v=M�>ݫ�?h$�j��Ğ�>�-�s>�X�c= ײ>��þD�&��nپc Ӿ�V2�Ap>��u?�p�?P�!?sn]���+��>�+J?I�;?�P?�Z6?)"?���{�?[�>` �>�f�>QB-?"�1?�=?�>��>�`�����G�P�.����Ž	P���>���=#W�<��>Au;<��=��(<����|2=��=R 輔ʢ�.H=f�=�;->@��>�vi?Z��>��>!�?����O�J��U3?���Jz�=oT��<����5���>@�\?���?z�m?@�J>�T|��a��qQ>CN0>=�<��>�3�>8�ݽSԛ�4h�=tr�=}k������~��$o!�7�Ծ�������=ᾨ=a�?�^>MGX����=���RB��A2>��V����G��S�dnN�7�ƾ}x�>JyY?X>?�:�=#��v:��/�k�S+? 
A?8�D?�_Z?8�1�f��_?�#zj�!V�;�A�>���=?���	��>#���6��ѽ̶�>`�������a>uv	�V'ھ(�n��H�^��\B=���~aJ=��$ ־�v|�X��=��	>������ ��ؖ�8�����I?I�\=̇��IQS�ᑻ�4}>헗>6F�>��C���k�B�?�T~�����=��>P�:>�z����G[F����� w>�AF?�b?f��?Մ��Dp�M�?�i+��	��r�\�^?�S�>��>!�?>��=9y�� �u�h���I��}�>J��>^��A�-������M�,��>5?P!(>� �>T6K?X?=Z?��?}]?���>{��<����c(?���?ہ�=�׽�xY���7�4$L���>2Z/?��8�ƒ�>kR?�}?�^"?)fO?j.?b�>�s�U}<��̗>�Ò>Q%\�OJ��a�_>ÁL?���>])U?0T�?N>Av6��r��{���
�=�,>2-?Pw#?�?�n�>�>ܼ��A��=y��>o�M?C�v?3Qw?A��=U=?c�F>~��>�;<�>���>�?޻O?�w?,�=?���>-<�#�<o��9���(�<]S���:=-�=9�,�tӼ��<WE=�<4<��=�h��e�ٽI�½���[Sؼ"�?�sT>o�0�4�>�<���E�nBu>z�=
˾���I�<�n�=�J�=��?�H>`U������L�>�f�>�71��-#?�H!?ں??�u'�֌p��{P��͟���?�u-?�M>�y_��=��P�,{�=m"?+=q?o���~�y�^?�WY?��y@������/����J?�Y?.(I����>�3�?�/r?I��>+�Q�P-l�����ΧY���;���=���>���^�-�>��3?s	�>�2W>ذ�=��þ�9c������?��?�m�?"�?�h&>\ji���vB���ρ�W�Y?� ?�����?*I(=�־��w�#��&bվ�O��򫱾r�y�&B��n	�InQ��,��݆��?��x?�?�PR?a�־E�Z�%g�����+4I�c�
�7��F�4�	gC���(�A�_�V�
��:	�|���i����`���(����?ŵK?�Ԯ�4��>��?�����yӾ�>bV�q��z>������7=��]=۳d���~�A>侐�?Xr9>��>o�?��M�|�'��R,�� �j��X�{>ؼ>��V>NS�>���� [��c�'���Ͼ�*�#����CP>T�d?��R?G3m?S*�p�2���y��(���~;q�����P>->��\>�}8�I.����k5���w�T��:Ä����2G�=R�-?J�(>�A�>Dʔ?��
?�`�Ӧ��/z��(//�.�=���>F�T?��>��>�n�����{ �>�Il?��>0U�>������ �-�{��k½��>���>�b�>r>��)���Z�� ���A���29�� >ًh?������e�d�>ׇR?%ł�w�L;�>�!v��#�����()�&E>&�?��=�6>��Ǿ0��ޱ{�k��TD'?�1?�����:*����>u ?�5�>h'�>᳁?
�>��ľ�亻�/?9�U?$�J?�U:?�U�>$:�<k�ν��ý>9���m=��>��^>Nj�<j&�="�ܽ��g�G����=CŊ=t`�#���J�<%"����<�{�<?&>�쿶]a�<꾄�l$پ��ﾥ䊾�A"��,5��>���l�����OO��Wy���H�.H��]y�¬Ҿ�:��$��?�9@�Qþ��ɾ�h��cig������>
�&�b;��K�pwU��|���4��챾`'��]��Ë��Yb���&?�k��8sǿ|����,ݾ[O?�@ ?�y?�#�Q#�'8��">���<N���E�J�����ο������^?we�>~3ﾎ=��{?�>�L�>��X>�Rr>�Ȉ�6���k�<)6?�`-?���>îq�owɿ)Q��L��<��?��@�{A?��(�|���+T=:��>��	?fv?>��0�z4�Oݰ��.�>�2�?��?�'M=�W���
��Fe?��<k�F���ڻt �==�=��=�J��J>*��>��=�A�=�۽�5>2|�>��"�pL�E6^���<ۃ]>��ս�G��!Մ? {\��f�L�/��T��OT>��T?�+�>78�=h�,?7H�J}Ͽ�\��*a?1�?ߦ�?��(?~ۿ��ך>��ܾc�M?hD6?���>�d&�(�t�
��=v<�`����㾓&V�=��=ҫ�>��>	�,����*�O��G�����=R}�EMǿ�$�D����<}"�g�T����~�����d��S���pm�!���t=D��=�!P>��>�}Q>�fW>t�X?:�n?r#�>1�>��ݽ3���,Ͼ#�V�������)�׎������Τ����&��	�a�������ʾ��[��@P=�-T�^-���?�L�X�M�`���,?L l>�����g��	��	�ܾj�L���<k��O�gV��hh�}�?��O?�聿��E��#*��z)�����]?�=�t����a��f>����M;Ŝ�>���F'�cu$���B���@??L����%��b�2>� ��x)!�ք/?�>��f=0ӊ>�!?��)��9�">o˘={�:>� �>[�5>w���|U��?�`?�hs����t�>���V����0伋��=��9�#�ؽ���>�`�l\���@��y�-��ܽY�v?��>���Yg�
�u�K��<hf����i?T�&?��?��q?�� ?�_�=ś��f$�=^��΋=dt�?��f?d7�=���5�!M��???�5E?fR�>@�@�eI�BS���0�r#&?qz?B�?3���7t�� ��~8�:(*?��?����LG�aQܾ�ǐ=�}>de*?8&:�>�W���i?q?(6,��qܾ��߿`,���?��@���?�9��S�¿�����>Ӌ�>͉Ҿ0�ݽk^��n �*��=ݎ"?Up������ZĆ�����7E?� �?j\�>
�F��(뾬��=�L��Pӫ?~:�?�=��UV<UC���k��S��fx�<�Ψ=��%�ޚ)�C�ӈ7�o�ľ�4	�5������ç�>`�@_7ѽ!��>!B4�=1��Ͽ~G���Ͼ^mv��x?�ݪ>��н{栾��i��u�mBH��I�������>��>�ϒ�)���@�{��B;�����d��>� ��N��>S�Q�����䟾0"<R��>k��>0ۆ>���Z������??X��9Bο ����(�X?�4�?�?�?��?O<4�w�Y�{�����F?r_s?��Y?�q ��[�u�0�r�l?����L�[���1��lC�ݤ@>{�-?��>�'0��ދ=�>���>,�>��(��:¿Y����6q�?���?xJ�l��>=t�?�J1?b���#��wܜ��*���g��t=?�^>>��þ��#��F2�M쌾�?:�,?H��a$!�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�!N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>hH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�o�>]x�?4��=6��>/)�=+�����9@�>$>M~,�q?�uI?�8�>�=�r8�@S,���A���O��F�)/C�;�>c!c?E�I?yQi>�>����G��!��F��Rz@��C#��
<���3���ֽ��->He@>Ă>-�O�pѾ��?<���Կ,N�����b??0��>37?G����Kz���'��c?-/�>J�
�t����:�����|�?�?��	?��ؾ�N���">���>(�>ĥ��;���h�,1>��6?��Žp�����x��Y�>�3�?N� @o{�?�D[�܇?q�'f��yl�r搾����wX+>��&?�*���>� ?P�p���>�U���sg��h�>��?�	�?��>N�k?�q��L��W=�ˊ><Ra?&2?�⌾�ؾ1��>k:?�B8�Ew�����;3?��@�?@��e?���� d���KͿ�(����ľ��>�.=�p�=1�*���=ȷ<��m��w-���<`�>/\�>؃>��\>~7H>�!>�Ɔ��(�剦�����Q0�kվ�&��ip��Ȣ��ץ�����̟�ZQ̾�=$<��V=<#�<���������Q�m<�=W?ftj?�Jw?�_X>X�oUW>9A�ŀ)>[?���K=�J>I*�>��5?7�>Ϸ�=yV�(*l��={�n�n�Bѕ�മ>�ӌ>��>U�	?���>�}�=�؉=�(>���=9���&>��ڼ�'�=�~8>䝐>c��>mh�>\y�=��>N�������l�Zf���jI�3�?���p�b��|���D�����в�=Eh/?��=�G����п�����+D?^y��{�z�ϽS=��?{pZ?N�>�MǾ?�~�\I�>"���7����m=���3���%&�Ӧ�>M?��f>�_j>�'C��P$�IV-� ��&V�>܁K?%q��p�h�{;Z���A����db>��?�]=!���͕�ⲁ�M�u����=�{<?��"?���К־za�r���>�Om>ᛍ=�"�=�$>#����$�G_>����<Ob>�׍>�t�>l�\>0r!>&�>(�Ⱦٸ����>�>��y>��8?�."?^f�O�7����;�:�p(Y>��>��O>� H=l��K�>��?Pv>�&=���=<���c\�d��>�;��G��<-�<�	�x��=}�A=���OU��n\��~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��I��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���=4꾽��t�W���l�Q�y�@>w�	?��N?y�� ����-!;?/(?����촿}�¿u\�F=?���?Ywr?u�$���~����p�8?��?�:?�Ց>�W������n>ՐH?�?.K>���g��7�>V|�?l?��>Pv�?��u?,R�>��!�c*�_I��y��8� =a��4d�>F�>�̾�T3�.���R�~�A�`�U6,��>]],=�>�Ž������l=L*��6U���λ�߸>�j>Y�q>�K�>A��>���>j�>K<7��~��p���vJ?Ɏ?s"�Pm��(%=�b�=6U���?�W2?�_���pо�9�>�p]?nF}?��[?" �>%�-���wϽ� ���Ecx<�M>�K�>�q�>ۂ����Q>�ƾ�P��h�>ŝ�>X��8پ�bg�_Y<�G�>� ?��>�`�=u-?��?�>�0�>��>� ���l���>c�?��?��?{??��H�5��'��\⎿�C�.Z�>�_?e"?
��>\������/�==�~�,H�K�?�+�?����F�>y?1?��"?yn>L@ν�'����=���>Ĵ?Je���}�Z+���&>�*�>�? �-?�J��V�p�a=���~����U�>��?��?�����L�'�	�B'�;e���J<��>+Tҽ�ؽL,d>Y=>�p�}k���g]=#�ݾR����E�;���>F��>�m�=3U��+Kľ�R8?�4��)�;��K>�]u�� �a�>��Z�w9��Ƒ?:��ۦ���P�Q����#�Y�?n��?`%�?�L@��o��pN? ��?@$L?�\]��k����8�پ�b�����a� Ƿ>Z;�=���>	蠾�ƥ�\쿿FW������$���>bH�>�?j)�>��N>OǱ>$A������8�`��c�W�?����0��8)��^��A`�]�J�ZϽ�����Lf�%�M>L���l�>��>֡�>?d�>/F�>��<<�p>�kD>��u>���>�{Z>��>[��=��=,����@?����;�%�
��;��O?�O?��><��<X-m���޾��*?r6�? �?H�}>�^a��52��g�>*?�vZ��Q�>�L��ɜ�:�ʹ������H�����%<%�]7�>�׌<#oS��<�cl ���?��?�G�Z�ž��ʾ�Z��}b�T�?��;?v�C�U>�0�a�u�F��a@���$=AMz��-��k�"���[��|��kp��Dp�N����#�c8?-&v?W|�nh�\E�ϕ��i�]�\4�>Y|?�#z>�%?���>d.���4���S���3_H��"?�~�?־�>�$I?o>?��S?l�<?(`u>���>c���{�>A��;�*�>���>�*?HQ-?��'?,?&�(?j�Z>O��%����eվ� ?�?�R?m�?�>��z�gD���@�rGx�?Ti�k�;�yԲ=[�=�%νm"�4x=�5O>�ʴ>LF�B|y�}QW�DQG?�#�?|KúC?N�B=a��<��րt?�WZ?��}=Cɾ��t��q9����>�%�?㘟=�܁=_ǒ����=��6>��޽�b�l�����=I߷������)��Q�>=>�>=h��=̋�=�*v�|	��2����t ?ES?�;�>�p�>�߆�� �f����=�8a>e2T>��!>.�ؾVn���ꗿ��f��y>��?J��?'�j='��=2��=����C��t*�겺���<L�?�#?�T?Ȓ�?y�<?��#?�<>���3������w��A?�w(?���>,.�7¶��f��#�7��?Ν?�c�o�?
���þ�:�-�>���naq����QD�pj�'������?ً�?�Z�_�9��6��9����ج��FC?�[�>�+�>���>Ĉ&�I�o�a����D>ZL�>�T?U
�>OP?_g{?)�[?�1R>õ8�ͭ��ę��
��>~�??�f�?/I�?�x?	+�>c�>h�)��(�7��	�����Hu����X=�?V>{��>w��>���>O}�=��½����{?�qP�=]�b>L0�>Q�>l�>��w>��<*�M?s�>I񭾄��멾�8���;���t?S՗?�0,?m�=L����F�W������>!�?���?��7?��8��>BO�<�ھ١��۔�>�p�> �><YF=��t=��S>�+�>���>'@��S��c%�S˽��?7aF?�p
>+�¿<�m��{S��=��u��R�����Z��a����`��I�=fn��o� ������Y�p�����̭��_��b����0�>��F=���=�[�=��!<����I4�<�:=�.�;�H=,a��(�;�>!��.�p�~�����C;�WR=A�u�ƾ'x?�Ba?LJ?�p?E�k=I�=�m>��y���?��>"���3�½�]v��~Q��z�q$;�ġ�\�%��G��K>��罦��=��=a(;$"���q�=��\�B>C`>{�L=���=k�=6#��烼�a�= ��=�6w?]��� ����4Q�KZ罛�:?�8�>�z�=��ƾ�@?_�>>�2�������b��-?���?�T�?B�?]ti��d�>=��@㎽r�=����=2>��=w�2�6��>��J>���K��k���x4�?��@��??�ዿŢϿa/>Ē=>)h>�`V��t1�.�G��R��iS���!?�4���˾��>~y�==3վ�'ƾ�=0/>�<$=�R�՚Z��ו=|F�"�|=Ob�=cy�>�->��=��~�g��=��*=f�=0<>.�;%�<�P3�~�E=��=��T>K�">D��>��?��4?��]?^�>nт�@���|��6��>3l�=��>�Y9=n��=�g�>�t$?��9?�@?v�>(�	=�o�>���>�7��;����)���;�ي?��?�G�>?�<���Q��<79�0<���D?�.?��?z��>�U����9Y&���.�%���	z4��+=�mr��QU�I���Im�4�㽱�=�p�>���>��>:Ty>�9>��N>��>��>�6�<{p�=ጻ���<� �����=&�����<�vż�����u&�6�+�1�����;Z��;7�]<O��;/��=���>�>�>�O?X�/�o^��:=����Q����=,�þBXO���C���x��D(�u�R<���>X��=�,�:2���5?nR�;FJ�=oĶ?+�d?�>�<�⽾Ӥ�|�B��U>�S{�Q�(>l����|�|�G�I�\�	!龱-�>�y�>�U�>(Fn>/9,�n3E��j=�WӾ��8��>E��A<ܼǠ���c����� ���1�h���<Ϗ@?8$�����=�B}?�R?�Y�?���>�$��gݾ�->}#w���=���Nz��N2�|�?��!?�>X8�WH����4��ԩ>�[�˛1�o�����7�Ƽk=�:վ^��>領�qbǾB!���������-���N���>�,L?'?�?� ��s�f��U\����o�����?�C?Ы[>�-�>���>��۽�����rھ�tȼI�f?���?�e�?I4/>��=�o��q��>��	?���?c�?$�r?iH����>aE�;� >�÷�g*�=$ �=��=Y>>�?�?�z? ښ�|`�Q���S��,F���<(��=U��>;\�>�@�>h�=y>%=[��=J�c>���>R��>��`>��>�|�>�$�����V2?�.P>I@>>��,?��>M]�<�ȶ�gtS<5���.uT�o�=\���ǽ�5=e�]ջ;�������>��ÿU��?��a>̼�p�?4�򾱻����>�\N>�Aؽqf�>ϻZ>��>>���>9�>��={:�>v�*>�'���>|D��&�<CK�9�g�k\��q�>T\_�[	��汾K쩽�j�L�s�A��E?V���b�x2�^j�=y��?*����Qվ��U��:���>E�>A\�>o���>Y�;<�?׸�>�]*�^���)r��A��t��?B��?�;M>
��>��Q?`�?60a�w��I�P�Aw�1x6�bR]��V������tx�Y6��V��r^?Max?�b+?�
%��I>=!y?��6�
���.D�>t�0��?��V�=W��>����>4i�h㹾ҍ����ٽ��L>��^?]��?M?:�4�����+�>:gW?�T?B�?"#�>�iN?˩�?4j?��c>��A?�?��>�_q?De�>�(�=��p>^	>,0�<mD����5�|4��Vp��g���8�=���=�C=�w=�DS>3FP>�h?������`G=t�=�n�<3�>F��=$k�=�n�>3X?A[�>,�>G�.?K���X*�j����-?ѠD=�@��<D��L堾�d�=R�k?8~�?��S?p K>�>��yW�ӳ�= �>k4>x�M>���>Eۡ��)6�U¼=�k
>�>r�=�Ƽƍs�ƌ�Ħ��c��<��!>ސ�>w�>����>��������>��u����R4=����Q)�{\�����>��z?�/?6<���y8�.�P��4?H�t?��%?ps^?�93=~Y,��\:��4.� �-�撁>@��=d��|��E��J�6�@�=�ʔ>-��2���
d>��
���ݾlp���G�Z��w��=�
��sG=���ek۾��c����=n>+����!�a��������L?��i=�A��~�d�������2>͑>�W�>�+��;����A��P��Ԡ�=?��>S�C>���yB��A�A���q>��<?�S?�?�+A��m�����*�T`��oI��x,?���>c?���>�(=�������{X���.�<Э>i��>|`���[�aνn�$��&+�F�e>[V?�� >��?K�R?m'?�=`?�G?P�?�{e>T��<�ۅ��%?�&�?E�=��Ž_oN��8�g�C��k�>�I(?��C�Bؘ>@+?��?;c(?�DP?C?e�>�@ �3�>�o��>响>v�V�����B
i>`�M?���>iyV?�0�?��@>/V3�b����A�����=l�+>;�3?`�!?<�?�M�>k��>E����+�=�^�>��:?�R�?�u?v��=�	?R!>3T�>�=e�>���>��?�K?Ɵn?��F?}��>0��<�׫�t�����j���<���xdL=}B�=KC�a!<YѼ�/Ǽ���<dC/�a!s�o|f��L��.���Y< ��>�Y>a��P4>�	�����*�e>� ��go�0��,v����>nW�>���>bX�>hm�x����P>�ϑ>�:�F?�4$?�xZ?�?t�r�{�<�˾,���V5;\b?�.>2��pk��w�Y���=&6P?�c?/K��i���b?K�]?���?=���¾VXb��X�b�O?(?�H� �>�~?�Xr?���>�4f��Hn�%����a��h� �=���> �6d�YӜ>2=7?���>%�b>�Z�=��ھ�w�'�����?���?E��?���?�s*>8�n�@+�i���do��Do]?��>_)��1�!?�>:<��Ͼ����t����ݾ�����.���꓾�s���#������Ͻ�ۧ=M�?��t?Eeo?��]?h�J�d�/{]���~���W����Cv��C��=D�R C��/l���M���wי��/A=�)V���.��L�?�s5?bc�gK�>���p ���边<>��ƾ?'���Jv=~L��Qȉ<���=��O���9�T᩾9�&?�:�>�Ϩ>�$.?�QQ��*K�
�@��(3��~Ծ�� >ә�>��>.U�>�u�=I{}���������U'��x��F%=>� h?�[Y?�ml?���,�.�+I���;���������W�G>��9<	`�=�vq�m8E��I
��"�"�g�Ӛ%�ɧE����O<�??aj�=F�>���?�C�>w��/��~���O�(���)>��>��G?ݵ�>��>�]����k��>(�l?���>R�>:l���!�?�{���ɽ���>�ԭ>�.�>W�o> 4+�b/\�;\���y��J49���=�h?~^��Ų`�0��>zR?]R>9�F<�x�>+�u��}!�Ģ�='��r>�b?�=�:>��ľ����f{�s���<['?�
?�ӏ�I�&�-�e>Ns"?�[�>���>QY�?��>�}���`99��?Y{^?�G?�@?���>,�(=���4wĽ��&��#=娈>�[>.E2=�x�= ���#^��j���A='ڪ=��Ƽm���0�;�妼q�;<��<��1>��׿\N�����E�x��oS��h����>l��sH��	��dվ�����5�$��<�<%�P^u��(���v�����?���?������>Z���l�����<��>�㉾��ϼtݾ� K�������Uo�~��u�h����𭂿֦?c����S׿�M���o���a?4�?� j?�E����e!>�h��=���>�/U=Bf��X��>z��P��?�U?�O�>B�+�e�'�>�W�>7D?>��j�M>���߾�v�>>�&?�,^?�fq>	�m��?��sּ�����_�?w�	@#x@?r&����9�@=��>��?N>>��(���KI��0��>���?!4�?DY�=�<Z����b?��g�� F�Y"��6O�=rS�= �Q=ߠ �mp=>��>=1��79����U'>���>1p[��|����T��<��l>u�߽�M��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=u6�����{���&V�}��=[��>c�>,������O��I��U��=�F��8ɿ^��������<��༼[���B�����f�~��{޽��=��=�/[>3�>��J>��I>sz^?S�r?ֽ�>5|�='Zܽ�*��p��dIG=ڧq��8��
��2�/�͇�W���澖P	����o ��ܾ��>�֘=��R�9���G:�Ԍd��S���6?ժ�=j����c�����-���4ž�`�=sϏ�|a�ȅE�����Ǧ?�D?�#{�'�a��e�ތd=��q�=	f?�V�'D� ���,6>Q"=9<$=<g�>J�R;�[辢S/�8�W��O)?%�?������>fȗ��=�&?��?cV��Z�L>18?��DK�=ocȺ��$>]r>J�|>.0�=႞���v�>�g?c���Cľ0%�>�R��I2�U�=;
=΃�<��%���>���=ws��/=>����Cnb�wxz?��>of�a��}:�iе�� ��>v?��??��>CT?(;?���>�'�RZ+���F�7�;�2.h?4��?���< d<��	�V�� �U?n�?r�>K+ƾ���75J����Y��>�I�?�~�>�y>�6������������=?���?��p�i���MƾM+����N>Z��>b?�U>��[�=�\o?��"����lɿC5��	�?`H@�@f6�Ú��"u>�|�>�V�>�J��!+���$3��i�f$>fX�>Fm��B�������y�L`?S�?�r?"/h����2�=��[����?�%�?ɼ���h/<�B��i���	���ܽ�>}h��ծ�z�ݾ�\�Z��������,����轑Q>�3@������>��ӛۿ[Ͽj����ɾ����?�>P4F�`��JM��m���B��E�m����>h>|l������{��k:��%��ܾ�>�|���>J�R��H�������_K<�E�>F[�>�ۆ>�j���q��uv�?����� ο��������cX?)H�?Ђ�?��?�?n<Lv�X{�m�����F?@s?��Y?�S��[[��g8�VPl??䣾��\�O2�X<��7F>��1?��>]� �;_=�[,>���>�LQ>*�.��྿�v��,���?���?O��i��>���?�Q2?O�'��K��Q���5&���b��K?+;N>��Ѿ]_&��t,�������?d<4?|�(���*�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?Z�>���?MB�=�j�>
�=����7�[^#>�+�=5�;��[?=�M?�N�>��=�9��/��dF�3R�&��e�C�V�>��a?�yL?%b>����3��� �,�ͽ�0����F�@��:-�q�߽l*4>X�=>�9>wCE�K�Ҿ=�?g\�H�ؿ�u��v�&�c4?��>��?����s�G���K_?}h�>���1���0��M���x�?�>�?g�?|�׾j�ȼ��>��>"�>$�Խ����c����7>�wB?h���<����o���>���? �@�Į?i���(?Y�$���F���H�
�&�-{�v�:>f�?�89��Q=_?2WQ=�*j��IÄ��>�?�?��?��>� Z?KI��6��
�=�5�=j@h?D�>�ʎ;�Ⱦ��$=��,?�����N��АԾ,�S?D�?�@6��?
B��N������i���*Q=Z�=p��=������<_�\<����i=�3)>i��>>��>���>�k>~�>�)>�݇���*�&F���-����;��� ��I
�):����+��j��Q���FҾ��;�$�ջc�c�9�V�0��<���=5�O?_T?��s?���>�A1�:�a>+�H<,J�CɁ=�R,>r�$?'M9?�??l�=�E��(qZ��{{�j[������b�>�(>��>���>�>򆊺��>aoG>KJ>���=�޲=aTͼE�=$Ka>��>E�>AϪ>�a�=�<>l�����\�Z�I�/=���@s�?~���A�䭴�?��@10�Hm=I�6?��?�D؅��
Ŀ�l���W?�z��A[��t⾿h�>�Lt?�ڂ?L�3>9	D�i�ν:�0>��%�@0ֽeo�>W+��à��/�Ⱦ��W>�~:?�zp>�o>�(:�ɓ0��rM�h���q��>�5?}V����<�-�w���/��7߾�Z�>Y�>�U�
���C��CRy���g�N�a=��.?�%?p ��eɾ��R�.Z����:>"�_>r#88�>�>�����W�<!�e���=���=�v^>��?Q�>e�= «>z:����=���>��7>p�,>Z�9?1�!?�ON������t�)�#�$>}>���>x%�>̢�=��G�D��=5��>6k>��~<b&���4�]�<�+S,>���H M���l=�������=Si�=/��n�G�]=�~?���(䈿��e���lD?S+?_ �='�F<��"�E ���H��G�?r�@m�?��	��V�?�?�@�?��I��=}�>
׫>�ξ�L��?��Ž5Ǣ�ɔ	�0)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾSa�>�~�oe����@�u��E&=ă�>>)H?k��G�N�%>��
?�?F�Ӫ����ȿg}v�T��>��?�?��m��2����?����>��?HLY?Si>p۾�
Z��v�>X�@?��Q?�>@>�q�'���?�ض?���?��6>�q�?�}s?+%�>�x���,�����v�����&=���xw�>2�=�Ͼ��A��?���0��-�a�5���>�=S��>=ý�8��E-�=Ԫ���6����k���>DL]>�4>��>Q�>.I�>m��>d��<F@���y��ǽ����K?��?��O
n�@��<y�=|^�a&?~F4?t�Z���Ͼ��>n~\?/ǀ?W�Z?�K�>���5��tѿ�Mm����<8�K>���>3��>ݻ���7K>�վ�	D��_�>V��>2*��Oھ]~���2x��'�>�P!?j��>�e�=�=?�E?��>{D�>��)��{������u��>wp+?��>��l?0T?��Ⱦ�2������z��E�U2�>��x?T);?��V>�[��������=�>|�����CR�?Ÿ�?M�?>Θ+?۾�?��?��?p�>𱒾��ȑ>ܰ�>Ս?���J.D�w&�fB꽛&	?�O�>WI�>��h�'!����!��=�Ң�D�?�"G?��#?����_���ž[�<�����㾼�[$=�'q��
>]@B>VI��h��=&��=���=HM��%P�0ʰ=�O�=�]�>�>�<�貫���%?�l�=��+;JЁ>)�����0��4�����*m۾�ˀ>{ћ�M���f����k��R�=��?�B�?�Ϫ?�'���n�$�$?5 �?��4?��L>��н�䊾ǩR�|�ξ�Q��_�S�� 7>{^ ?�W�>Q�(�e��jEϿlӟ�gm�=� н�?�?��:?�=4>�>~�?�l�@�=��'�l�ʾ��W�<S��G �0��NҾ�U��Yo������c��ő��w1>j ̽�n�>��?薤>o��>GTv>nh����t>�h�>-p�>�t}>�Y>\�=6�>�+�@�潡�V?�ﱾ"$����ͨ����2?��]?u��>Rr�<@����[辎Z'?�	�?���?�=i>Oo���;��l?9�?6��T"�>߮�=>��=\������Gν�Ax�>$�醾>��
��A�P�N���� ?�?=���39i��"R���=��?�%9? �3��X���G��\���O�����؛���ƾ^���R��x��	�d��i��$�I��=�^<?O�o?�O��!�h{�������9h�>|�?��r>.$?��>o���	)�j��R�����?�T�?ű�>�}H?�_9?B�M?�M?$�>�R�>���ݏ?D-\=BF�>z�>6�<?^&??CS0?�
?��?��`>w�����߭���2?��>�$"?��?��>����!����<|�ٻWWh�j#����=��=�>��U�=��=7�O>o��> �>��@&���_?��c?���i�?0�����?W����N?�3??D˽�� ���q�J�\�4GR���y?���t?^=
`�>d{�>:�>=�:���=���;r��=d)��Q891Y,�P_~=0��|�[��]y>3���n/q�)B�}H�>J�?�y�>*'�>r���q ���O��=�qV>GaN>�>T{ھ�}��oė��g�:{>�J�?�^�?��f=,E�=�y�=@@���Y������輾!,�<XR?�#?R�S?�}�?�+>?�|#?l�>�Yؓ�b����N���p?Ӈ+?8�>x�
�����4��h;�)w?��>��^�$��p��^Ⱦ;꽿�9>O�*�N�}��멿6�B��|��#;�7R�s>�?�?��,�'=�f<پ0ݘ��e���3<?H��>M�>�b�>݁&�@Te���]>Y>a	�>�I?�>�O?[{?�[?��T>\�7�]����6L�O>�8@?F<�??8�?"Px?ҟ�>�I>��(���߾_V����8������L=[Z>ɔ�>f�>���>���=`�½[I��\"<����=�eb>�M�>C�>���>��w>�	�<��G?���>dP�����e ��f���:�<��u?��?�z+?k�=u���E�1K��E�>h�?��?�(*?�S�\�=�Rؼr�����q���>䰹>7�>+=�=X�F=Pl>��>�s�>��fb�{r8�C�L� �?�F?��=ZCſ��p�:�q��T��2P�<������g�����u\�=�,�����ܸ��>�]��4���`���q������ғz�KS�>�9�=�q�=���=�γ<�\üe[�<�P="��<=��l��/A<��5�t��q���W����Ec<��L=	�&�D��E|�?Pei?R�-?y6?�p=jB">��'��}�=�&�2C?�㵼������Ѿ"���W7���M�c�ܾ��S�K_�<J`��9J>ӦϽ�f=d��=��S<��r=�aD>�,�=��3�������n�J!>.Ϗ<�K<�[�����=ڋ<>,�y?�t�r/��w2��/�c?fPD>g�?>�%Ǿ|�?��>�q��Iſ�"����?ѻ�?���?,:I?���X.I>�Y�q�=���=��ýT
> ˦=`����y�>��S>4�B�����-�V<:��?��@�\?�B����տ�Ud>b@L>^ >�IU��'3��½���誾�"?�+�wО�v�E>��<r����ž�S⽚|3>��ּ�V��tM�6��=I�s��)��s�=��>Z�F>`^!>`���P�J>>	G���=K7>#�����=O<��| >��>G]>��L=�0�>F%�>t�2?��d?&=7>�G��@�|��޾ q|>�r���y�>5i�=�^ >��>�<?�17?�F?t�>�	��ۍ�>[HD>��7�U�p�;�ϝ���=>Ս?�r�?��?(�<R�Z��k��y,'�̅����?30?j?���>���b]	�c�"��q߭�g�
���ɻW���}��i>ɟ�}�����<��>�|h?:�?4=�>��=���>8��>|�m>iM= �-<�ĳ<�>�a�=���=C_�q�	=��B��|Ľ߸<�W����;`m<�g���;�~���6T�=��>��>F�?B�ܽ|q����i>�>�$�X�l���䱾�oQ�@�a�<N�H�&��~��Q>>~�b>�������g�>�B>��P>�?�k?J�@>{�̽넮�����g��<��/>	�Q=9	�]��j���\�ٮ��4H�>|K�>s8�>�6�>�$I�].l�(�c>'7��c�:�-�?di޽TT?�!FJ�@�66���{��H�A8���?k��%>�ń?Toq?��?^Ҍ>F(�<�оt�=hо��罉������@5��Z��>�;?�	?��Ӿ��&�y�z�$���ǫ>t�(�خ?�ޜ�za$��4�<���:�p>ϩ�r���g+�	ힿ������!���%�A��>/�b? ̬?�@���V�f������L�?HRX?�0�����>f�)?���$�ھ�tI��PA��-?bC�?�=�?��=�D�=�~���8�>݈?>��?Cʐ?g�q?�WS��5�>����0>P�r�oy�=31,>I�=��=Li
?}�?�?�����k	��F񾢶��ފd�� �<���=�j�>dC�>J8�>��>|�=G�=ʾ[>(�>��>��x>�q�>c�}>���$��--?��D>��>>wj#?޹�>S4	�I�3�q�\��}����w��:-�.M��GAݽo�#=��<ձ�;;���F�>kyĿ�I�?J��>��?xh�������>g>��"���>�0�>FZI>�R�>��>�&'>�݁>�*>�Ǿ�4 >)�
��bj>��_V���ؾ��q>�$���Q%��i
������Q�x�Ծ�b �}�_�`~�Ө9�h^m=�N�?v&�<>R���.�j�G� ?��>T6?�ޔ�;�ý�$>���>gd�>K���q��#9����Ҿ�`�?���?=�W>J��>�NV?!?c��rE:��P�%v���A�"l�Y�T�Sy��c�����͙��KoZ?��q?�:?�����h>���?�E!�!:����>��2���C���<̊�>?����S�O�پ3\ҾǬ�_F>�a?$�{?)�?>RJ�A\��,�>LjF?�.?�<P?Q��>U�?Ā#=	��?���>M7;?� 1?�|�>֍N?��?|um>�2>�6�=��y>�t\�8pz�G�F<�$��ܽ ���<�a=ե=+�=�53<-�\=$Y��������;a'�=��|=��4=V�=ᥠ>�_?)��>�*�>�W7?�&�;;7�7���AY(?K��<2i��q���F��rL��Z: >΃f?���?x=S?�T@>��@��E�#�%>��>/�>Zc[>��>�4	��\L�!͒=�]>�y'>�޸=P���%��i=��Ɖ���<" >6��>��m>%L��M>�;��凌����>�m�Tƥ��.1���*�����ń�Pъ>�b;?�D?7�=��о�`߽%@I���9?�9R?�??�Ά?�r��%��!�4���Q������>�����/���鍿�s�T�Іm>��$���!�9>����پ�t�$�N����ɖ?=��^�<��R^��─�I�>��>�����E�w���(H���>O??�u=����=�d�(���L�>���>��>p�K��l��-�1�]k��|L�=lE�>-E>n�S�$�I����7 �>LyE?'_?^w�?@�����r�}�B�wT���o���ϼ�w?�J�>�\?G�@>I��=j>��>���e�/G��y�>���>����}G��/�����m�$��<�>�E?��>|�?��R?�?'�`?9*?�F?�Z�>�S��(I���A&?'��?g�=��Խ�T�� 9�2F�X��>z�)?��B�빗>H�?Ľ?��&?�Q?յ?{�>ѭ ��C@����>MY�>��W��b����_>o�J?���>N=Y?�ԃ?P�=>A�5��颾�֩��U�=">v�2?�5#?/�?�>ֺ�>�"��an�=@ܰ>��c?��?�q?r��=ϟ�>b9>l\�>�Ҷ=;՞>��>�?�M?��w?�gD?�i�>�<���$�������^
��d�:��<b>�=���v�W��׼�$G=�ڃ<>Xɼ�h_�� �sQX��N~�?NZ<q��>+�C>�ƾ�5�=����Ο���=w���0Q_���n�	����>p
5>�K�>ˊ>�$}�U�b�'�>���>�v+��IA?lh?��/?�q#=pf��T��:ߧ�J5�>v�H?L<Ҵ2��r����h��E>ytu?I�n?+�\�{�
�v�b?��]?l���=���þ��b�Y��O?��
?��G��	�>��~?��q?��>��e��Cn�G
��4b�%kj����=���>�-��d����>]Y7?V��>bb>��=r'۾��w�����?	�?� �?��?.�*>��n�"$����8���
2b?b��>%�F�?��<Xdվ򸣾)`p�Q������>��5����Τ�'���
h�~�ֽ~�=�A?�q?�Yu?e�^?>��̞c�uk��e~�";R��#澺��&N�;I���J��yp����:��%򕾇�Z=m���v�3�� �?
�+?���5��>*�m�B��� *���b>	@���?0�� �=�����!=���=O�+�kwE�`����*?���>i>�>w;/?��T�ո8�+�R�'�C��F�>��>��;>�Y�>
�ܽ��^��.W���D@���z�=�u>��c?�K?��n?@� ��Y0�4���X"�*7�`訾��?>�>:I�>1�X� ���%���=�bs�#�w��-	��w=�2?��>,��>!��?]?���x.���z��1��1�<驹>kdi?���>	��>)'׽��!����>2�i?M�>|��>���9
"�4}�pv��O�>���>���>�?>Hk>���e�����ҍ��i.��/>�^j?�A����^�`cg>S?�c=�|=�>��x�����E���w����=��?��=j�?>љ��%��g�p������x)?��	?�>��9)�*�n>q�?���>�A�>�Z�?��>�����h<�+?!�[?��I?�N=?4��>V�=R鰽qŽ�*�+�&=���>�NP>br�=h?�=�W�~�a���%���L=�=�ٞ�Ȣ�5�:���%�<c�<��1>\Cٿ�@��5��:�ܾ���[l7�b���?Ľ�	���uN=Z�꾼e �WǾ,۩�b�:��������Q��U���Z�?�G�?:iT��S�4���V`<���>�Y��N�X�Iz������ �ܾ�z�`,��'K���W�fb�h�*?PΛ���ſ1��-��p�?�,?5�{?��s(;�rF��=��޻��8=���)y���ҿm#��kH_?��>�s�;��F��>�s>a�>��\>cɰ�&9��j��= ?A8?��>r��t�������o<��?��@�A?u5(��:��I=���>p	?�EB>�N/����.��x��>�=�?�0�?.	D=�:X�ϳ��1e?s�8<�E��|�9��=�ϣ=4x=f����J>g �>���ʊA�5�ֽ�6>8�>��]��:Z�f?�<�X^>��ҽі�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=����ֿP��9���<E���D�<x�z�a~�|�?=@c���`<�tݽ�L�=��>�zn>\��>��V>�6>&vw?��Z?��>t>#>�<�ǃԾn�_&������Sͼ˔Ǿ��轐軾��ؾ�T��\�����>��>>þB�)�HZ�2�:��Ra��FY���c�s9}��?�ȼC��x2
�ʂ>w���h:oz�=���=3d���BX�1��tV�?,�'?E�����]���!��Ƚ�H�����i?d�	�;`��,���>��>��>Y�>�j>m#վ�/B�:�]�̍7?�P?@�rm���T�=�ֽ�>�~?�t?O��=E3�>\~I?N�>�Ͻ$oZ=�vG>◨>:{?�R{>[���h*�U�'?�U?�����ȸ��3>RѾ#p쾙5>��]>裂��d����>��=K���D@�۷Խ�y6���_?�2>��$�}6�l�m�m<����<5݁?C�?�=�V?��)?O��S�������
��Ľw?���?�9">
?��F��R�u��>m�l?_�?J�"�����t��*���c�>���?�W?���:�)l��p{��(��Z'?��v?�r^�vs�����I�V�i=�>\�>���>��9��k�>�>?�#��G�������Y4�#Þ?��@���?%�;<# �H��=�;?f\�>��O��>ƾ�z������!�q=�"�>򌧾qev�����Q,�n�8?נ�?���>������>��=4ٕ�0[�?��?ӂ���Cg<$��yl��o��S��<ǫ=� �)H"������7� �ƾ��
�n���)뿼���>�Y@U轐)�>tH8�
6�[TϿ���YоKNq�:�?�~�>�Ƚ�����j��Pu�ڱG��H�������>�fz=�� *a�A��2�7� �-�o��>ﺐ�y >���m�)X����=g�>q`�>ص}>$��&߾v�?�޾�HοȠ����"9?ǋ�?kƈ?�O ?s�n��A+����2�D=��V?��Y?��_?"���l�������N�i?(���a��55�xm9� �B>��)?�;�>R�+�M!o=)�A>��>:�>�5"�lX���j��W��I��?N�?j��9?
��?#E/?�a�8ɕ�̹��;�3���y=GdB?��>�A�����/��=Q�.?@i3?��?��e�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?ֵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>cH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?x2�>�?+��=F��>��=燺���>�� >�:>,	����>�S?=��>a��=���#}$��<�A?H�r����D���>6�\?�H?x48>$�7�)cJ��#��e��:
��{T��8���O���X=>J�f>��:>P4��Ӿ��?�o���ؿj���o'��44?u��>��?���E�t����s;_?�{�>7��+���%���E�G��?>G�?��?�׾
h̼�
>}�>bI�>��Խ���� �����7>v�B?%�C��J�o���>���?c�@Ԯ?i��	?���P��Ga~����7�'��=��7?�0��z>���>u�=�nv�ܻ��Z�s����>�B�?�{�?��>!�l?��o�Y�B���1=&M�>Ük?�s?�Lo���V�B>��?�������K��f?�
@~u@[�^?&{Wֿ�뜿�T�������=B3�=�2>�PڽȄ�=�'9=��6�W������=<ݗ>H�d>>�p>�	O>u^;>�)>	����!�Be��6���sD�.��d�`[���� v�h�'4�������R��7[ýb����5Q�e &�߱_�H\=�?c 7?	�?���>`L==�+g=��4�as<��j�sP� �=�(K?��2?�3?��=RH��`�`���>��-��#��>Ӎ>�?�%�>�Z>��=W˹>��>���>u_b>�= _4>�F�=�/>�#�>��/?���>��>����㓲�ȱ�*z��A	��۽+���?�gξ�n��}A�d���c;�*�?~�=?H�>W�����ݿ�ȿ�?)?��ݽ��\�*���>8�F?=d??��R>_�k�n
���>��ݾM��?��<�j��S���j��T>�m]?:�h>�Bs>�3�W8���P�=���S�{>�$6?�T���<�,t��eH��۾^O>�k�>f�0����t떿o~�ozi��v=0:?k}?	��)Z��[�u�+T��NQ>�[>�=��=�0M>�ci��ͽ3PI�·.=���=pa>��	?r�>�D+�tP�>g��Zf��CK�>��2<_Fk>�I?g=#?��=O��7���46��rX#>bf�>$U>�S>4/�H���筶>F�6>���e�1��y�<�I>���X>�K���D��ܽ(ߏ=9�����=�|N=lM9�Bz=��Qn=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ4s�>Ҍ��W��t��S�u�|&#=���>?H?H��+�O���=�Gv
?5�?0`�)���p�ȿ�v���>>�?p�?��m�J;���@��v�>���?�mY?��i>�۾s�Z��u�>��@?�R?q0�>W:���'���?~۶?-��?�RJ>)�?�qt?��>�Z{�z/����ᕊ��Jm=A��<���>���=3�����H��"���Q���+h���D�h>¯"=S��>���Ǣ�����=����S����4`�?��>Bj>	�L>�8�>9� ?�@�>W�>�0=fr��y'}�uΖ�]�K?Ҭ�?���En��5�<M�=��^��?�B4?��W��Ͼ���>�\?��?`[?�W�>z��[2��yۿ�񑴾"�<��K>G5�>j�>�0��91K>Yվ* D�-y�>(��>Rm���2ھ�8���m��!Q�>�e!?��>U��=��?��?u6�=]�><c9��Ó��X���>�<?�$?�9�?*+?s����G�7��9�����\���>�v?��?�U>Nkp�����]��=C�<���[-�?;�G?�2�Hi?��Y?��(?f�$?ذ�=��j�FF��7x=HaI>^+?��C�@�X��3�Z}��<6�>�:�>�p?��u�����Y>1��Ҥ�?)+?�x=?�|)?�7���w���x��p'<�X׽�L[��T|=�n�<�	>/��=��޽�=��<r>`'�S�p�G�_�=�L�>�����7>�=,?�G��ك�o�=;�r��tD��>�IL>���Ϋ^?�d=���{�;��wu���U����?О�?k�?5���˟h��(=?^�?r?A$�>�H����޾��Njw�N�x�mx���>���>�l��徙�������$H���ƽx��X�?�2�>�4?�<�>�X>�t>Wݶ�BT������  �ndr�) ��B����B2��0X�-F������Yپ�䝾Qel>�,=���>��?->�.�= |�>S�5��ؗ>o�=Q��>�O�>��>;ִ>M��=vʽ;H��[nR?����#(��$꾥D���@?��c?�s�>�.w��h��w��,r?��?�d�?g�p>��h��+�"�?�<�>~`��0?cQ=h��sl�<�R���������0[��,�>2�׽�L9���K���`� F?cl?q�i��?о���4���H-�=Y��?�+?���b�B���h��=J�~Ja���S>����~˾�)�����6��	r�{X����>.`='�9?$��?�����;@s ��x���o���>�I?�;�>?f�>��8=����%L��e~�L�D�$p�N�?}��?,��=�Y�?��>?�_?�k?�߿>��Q>�����?Ϲ=��>��>�U'?�J.?&g3?-�?47?�G�>*|�����G��?���>3�o?�S?r	?M�
�-��1=�üs��uԆ�Fd=�8<~S޽\e�<��=|�~>[�:?-���]�6�C����=}��>[}?��	?���X,����>�_�>>��>IF!>tYؾ����S���?`o{?�*ƽjÎ=�~=C�>��d=[E9=50a=m���]=�$=a�����G=��w>Q�=���;�G7>�/>}-4�ocĽ�?r�?���>��>�w�m� ����Y[�> mm>.�q>�>N���`��'ݖ����s>���?h3�?_�
>}+P>��>" �����W�@�ʾ�e�=^�?��!?
�"?��l?*�N?u?��=y6.�� v�FVg�B�6?H1?D�>�X"�+�о�����4��y�>���>2�A��gX�b!��M��K��{T>n��t�j�m���08�� 1>M�������?� �?��<ce7�.y��V����Q�T9z?;��>�j�>�Y�>��F�b�Q���#���>�?�KK?�#�>��O?({?ԭ[?�GT>��8�\-��!Ǚ���-��4">`@?m��?qߎ?�x?N�>��>��)�g�߾�/��i��y���ւ��$W=��Y>�n�>�>!��>��=�]ȽX���~?�l,�=�[b>�l�>�{�>���>	�w>,�<
=H?���>���*������z���j==���v?�U�?�(?�'=L���&E�������>.��? @�?uf+?�I�;�=��׼�C���w��-��>��>Tl�>���=�D_=�~>f�>F��>�_��I�;�4/���
?��@?�=/�ÿ�>m�Zg�#���q��<�Љ���P�^v��jU��Ӻ=����
�Т���*Y��s��I����Ω�/���r�}�� ?��^=��>
$�=G��;T|ͼǈ=R�{=�H�r=T�A�q��<EP��( �󯃽���N]6;&�A=9��p+�ļy?a�M?�@%?��K?fi�>$�+>�U�[��>Uܪ��?�8q>;�T�Kɿ��U��ȕ�Qc���Ͼ]�ھ�^�R&���>@�Hb�=�+>��=�;�
��=q�=�1X=l����V=��=vp=�C�=_��=�,>�n>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�B>���=
pS�b�0�6�g��j���R��?w7�N,ξ��>:Ϻ=>�ؾ����Q�G=�E5>J�=�� ���W���=q����J>=Z�x=���>�+C>���=ꂮ����=�:=ũ�=�sJ>�7عr�=�C�^�_=T�=��a>F�,>���>[�?d5?�Zj?�m�>�9j���߾�J��!��>-h�=�R�>�����4>��>{�'?-�B?`J?���>�D�=��>VY�>��5��u�����-��?�z=��?lS�?`w�>V��<l��� ���-�H3��	?�8?��?�̜>��&�4���#��a����<6�a>���rD��쭁�U��PYνO��=��>���> �>�m�>oQ�==H>���>�2�=�ň<�>O)�q���՜���=�S��[Y> �<(�'���T�=�����
<������=��-=Ŵ=��?�ύ>��&?҃�=���>#��<��sN>B���>�9��5:m��s�0�4�%'>��=�hh�+���NT?��~>cx�>�W�?mRp?ؿ6> �z�<㾱��R�Ͼu����<��p~>4
Y>��v@b���n�������>��z>y��>g�>��&�:f=�;ן<��Hg���?�};�=�=
h� ���@��&>�؂�;2�D?ۿ��ve�>�ԇ?P�w?�?n�>J�!�q8����L>W���3�����㌾V�����?Q�0?���>��¾p�H�����g����K�>I�'�6�Fi����C�'��=����֕>H���>��Y_*�����������)��3�e�>�E?�z�?��"�����B�c�K��s���?
l?&h�>���>��>|1�=���V˽3�9=j�R?�}�?5�?�~>�;T�:>�l?� �>�'�?�?׽]?�����u?��=�r�������=���>bO ?�z>�	c?a �>zF�=�C
���+��h߾�'g��`��=�e>
�>^��</=�=��=lQA>���<��*>ƻ�>�[>�G�>w��=[�=��Ѿ�x���>?�Y3>�i�>�D?:y�>�Jx�#i�M�@=�����xB���6���[ˉ=ݐ�=��>)��J����>5����0�?��=��ž?Jξ���G*d�{|>}����>Tdd>�g
>�hV>N��>��O>]�F>aX�=,Ӿas>��[]!��)C�ʆR���Ѿ�oz>`���B�%���B2���qI�6r���_�qj��-��n1=����<C�?���k�k��)�t����?�d�>�6?�ٌ�J����>V��>鴍>=@�������Ǎ��g��?���?�Md>eƜ>T�Y?�$?C,�q+1���\�u�q��>���b��M]�����U>��]���ֽ+W_?dw?
IB?):�<�}>�~?��&������>�/��%8��_=ag�>������X���;�bž.����B>kl?�Ƅ? ?]�S�ֈ��QR�>��I?89?Y��?�DU?,Y.?��`��N?RA=_=c>�g	?�?%�	?U	?p�P>�>A�>�
���!穽���@��;�J�%ν��켁E�=��=nǞ=i1�=a�����ڼ��;=*!�������%�<#�,�^B�=v>���>�O?�?���>|�6?l�ͽ@D��y���Q0?���=��c���־�����T	�彌=�;j?�Ȣ?�V?��P>W0�H�d�*f>k��>-� >��3><��>��T�Sg�������T>��=R�=Ƚ/��z��|�4����^=� >R�>K�>k���4�%>^^���v�t�j>��P���WsE��B�y�.��E[�?��>�tE?_#?��=���~���g���,?�@?�Q?='}?|j�=W߾>�>�!:M�n�����>�L��6��*6��L���Ű9�=#7��T>���R���7>9� ���� ��$�a���������5�~�4>7��&����,��M�=�y>Ҽ����R[��o�����k?���=&�Ǿ�x�S�ܾ��W=��>�c�>'���%<�5����]�D>Ч�>&|O>��d&Ծ�':�=���3Đ>>:?Q�W?��{??Rg��|_��c�v��?]��3�w���?ǔl>���>	44>+,=\g���Z��Z���9����>5c�>y�'� �W������D޾��*� ��>�?�2U>rA	?�q?�?�p?D@?�j?ϙ?>��>���¾�&?� �?C+z=�b�ET�U:7���F��}�>��*?5�C��u�>f�?��?��'?B�P?](?��	>E,���@�w�>���>�V�L���8�U>��H?��>�[?�?ո8>�l6�9˟�Wj���T�=�>��2?I�$?�?t+�>���>E����=��>c?�1�?1�o?L��=F�?�@2>���>��=F��>8��>P?�WO?��s?��J?̎�>2��<>A���8���Ts�f�O���;M3H<��y=L���*t��V�"��<E%�;�Y���F��\��#�D� �����;�=�>:l>���*�>>q�ξ;a���H�=ӹO��O[�9>�����B>�>�i�>�yr>m�k�����ɸ>5�>���� ?^�?fX?/���b�2���UM�24�>�+C?�\�=j$L�b8��Կ��z�=��q?�L?<W?���)�^?�H?��>UK����f�߽3�1���:?��?��a��;�>�Wq?X$j?��?�y�J%'�ڨ���r��٠����=N��>8�%�h>s�x>��?�?��>K�>��Ⱦ�~��,B>��6?^
�?�y�?z�?��f>�f���z߿[����Ȓ�mK\?O��>`V���m!?}cZ�48־oy��%%����?K��I����������e)%��:����ܽ�\�=`6?�s?��p?��`?h��ze��]��n���&V����t����B�@�D�S�D��m�$o��v��9��`� =�����?�~P�?v�+?�R�U��>�ߑ��(��߾�G[>��#T��2�=qw���H=��8=��n�3D�O��$g(?*��>y�> �8?�a���A�|-��/�'[�.�@>aW�>��>���>�b�;�����*xľ9�������6v>�vc?.�K?B�n?Nu�{,1�R�����!�5o/�BY��:�B>�x>���>y�W����6&�X>�f�r�W��:v����	���~=ê2?�>���>�L�?�?�v	�Yg���hx�T�1����<6�>�i?�8�>o�>��Ͻ�� �C��>�kj?7&�>���>�ƕ��:#��0v��������> ֱ>j�>�i>��5��!]��C������!�4�V;>�ef?Kρ��n]�f��>-*P?ʢ��EX����>�X5�T�!��Z�)���=G�?��n=y->����#��w��q���m&?V?QJ����)� �p>��?]�?��>Ҭ�?�݊>gi¾�c =��?�j?ݺR?5�H?�&�>��"=�f۽����`�m7�=�9�>�V>4�$=رI=-�5� Gj������=�=��T�0A�@�=vE��+��H�=�,]>{�ݿ��W�����2R��c��Y��1�e���Ͼ�˟��x�;�eӾ= ���S�\N��&X���j���~�D��:☾*�?do�?��W�ԃ׽�I��}c���o����>ւپC��|��-F��DYq���������8�� �L�Z�]���}��/*?�1���Ŀ���w��"Z?m�?Ki?����G��[�
>z��;%�Ϲya��d���п:ׅ���q?��>�B߾����>���>%��>��S>��T���!��s!�4��>�� ?d��>�dV��"ƿ`s���6����?�J@�}A?��(��3�R=�~�>yz	?L,?>G�1��4w���w�>�9�?/�?�L=aZW����ee?4�;%�F�g��10�=���=5=t�sPI>^	�>|����?�ڽ\}4>T_�>�f"���� ]�&$�<��]>��ֽ����5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=v6�����{���&V�}��=[��>c�>,������O��I��U��=��ȿ���X���Â<$��8E|�J�J��Ŀ�1b9 ���5H��Ľ�&�=U��=Z�@>?��>o7>6�M>�:[?m?�`�>N>���iݦ�u5ҾgV���D��**�SY���,Խ� ��1@��޾�G
�����y�VܾL=��ԍ=t R�Dv���� �*�b��vF���.?�v#>�sʾ�M���5<%6ʾɸ�����l���+̾�1�53n�mٟ?��A?f�����V�T���en��ϼW?�������l��F��=լ�l=��>WV�=���3��dS�q'?��?3M���Ô��OO=X�F�j�=�_8?I�?�R�=J��>`X?�y'�����M�=^�>�j�>b3�>�|>dk���]��J�?/�Z?�3�u(���n�>�Z���D���m=�(�=�f��Ǵ���=�;�GK�Gt<�ֆ�7��:vTP?ee�=��2�Ar%�j�����B�i��<q?�1?=H�>]"�?Qp?12<�� �poR�����e	�<B?]�v?m5>l������(˾HS?_�o?/>��b�z��vi�|���?p`y?:�?֮`=�[r������]OF?��v?!r^��p�����Z�V��B�>V�>ҿ�>��9�~d�>�>?�#��I�������W4�Ğ?�@��?��;<�5��=�6?NZ�>�O�FƾJp������~�q=�"�>����&dv����FQ,���8?!��?���>5���������=�ؕ��Y�?"�?����.yg<����l�gk����<Dݫ=/o�PX"������7�L�ƾ#�
�§��S忼3��>Y@il�D �>T;8�3⿍UϿT���Qо'Fq���?҉�>ÄȽ������j��Nu��G�0�H�ɡ��5A�>�F>*��X'��Fu��Y@�Mt�����>����	�>5�N��h��'1����,<R�>DK�>�S�>�Խv\Ⱦ��?�]����ͿJힿ_����T?�՛?�W�?v\?İ�<_H��H��|Һ;�F?�Eo?��T?H.��V�>���Sc?s����a�GH)�5�(�/�=���>�J�>����Ȫ�A_>ؾ>6�<����)���ι����ڤ?��?F�ྜྷ�?"�?�nH?<�"��j��Z�~�u<���<$@l? Z�=m0�^ ��N����*?3�'?!�B��E�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?sV�>�q?�ř<=�>:�=$̼�Or����=�(,>Y  =��?�Gc?m��>�I>�)��`��B��1Q����s�?�vz�>��o?��N?�7>�RU��{ڽ��!�W伹~.�����F M��½������=V�>j'>,�����d�?�h�m�ؿ�c����'�F%4?���>&�?���3�t�����1_?[�>r5��)��N&���c����?`C�?��?I�׾Y�˼��>�ԭ>�2�>ս�����d��:8>n�B?_+��?����o���>���?#�@�̮?fi�t	?��lK���[~�
�1�6�8��=��7?0.�>�z>���>l�=�pv�򺪿\�s�ﺶ>BA�?Fz�?!��>��l?�o���B�4�1=~A�>6�k?.o?�n���򾒪B>��?a������aJ��f?��
@�u@�^?�뢿տ޿'G���I%���">��>(�>I+-�J!��K(>;��d	$>�T�>\*�>��V>՗F>E>	!/>ur�=�>w�a�+��h����y�k�c�S���I��������������E��镓�@��u7���̽�X�M��2׽$O���}?�iT?��}?[?�U=�uO>����7�>�pD�3o��NT�>.�E?��Y?��g?�a>��ʽ�U��}������@��R�>v�d=��>bZ?5��>�"ٽ�+�>C�>��9>�f�<K(ĺ����q��ma�=o��>r¡>�H�>�C<>��>Cϴ��1��j�h�w�s̽+�?����G�J��1���9������i�=Db.?	|>���?пa����2H?���{)��+���>�0?�cW?G�>��
�T�T:>@��æj�D`>�+ �}l���)��%Q>�l?�g>P�t>:�3��\8�@�P�+n����{>]�5?Z����8�zu��QH�jݾ<HM>A��>��G��j�����~�r�i�N�}=��:?>�?v��+����u��|����R>�T\>B=*�=>�L>��`��<ƽ�G�2/=���=�]>�>0�5>.~�7.y>�� �����>�R�>�t>��B?�&? v8��( �+�о$����n >���>[ǒ>M�(>X�/�t�W=���>ex>����Y.� �ռZ��F�>R�޼і9��=�3��=��F�4ԩ=�->� ����M���A��~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>S�)��d��������t��$�<�G�>��??����{̄� p����?���>�>�S3���ǿ��|��>��?K�?�;c������*?�W�>Og�?<M?Ƚ}>́��g٢�g�v>h�6?]f:?	��>!�?pZ�^�?\=�?��?�I>�?s�s?�i�>�wx��U/��8��Ǐ���=,5Y;�m�>�2>����*eF�%֓��c���j������a>/�$=��>Ej�G��2�=j����T���Df�ϴ�>(Oq>�I>!h�>>� ?U^�>l��>��=s����}����H?�
�?Ca�������=*�>SY��'?��O?i�*�о0O?h�w?8��?:Vm?w�?�������Aq��M"���U>�=>=
?s��>Q�&��t�>�
�������>�7>>�'��˾��~�j�M=��s>�v&?��"?Jy>��?��?�[>�v�>�G��ꐿI I��o�>`��>&;?P�~?KD?E���4�d����➿rW� �T>]�t?��?���>[I��1ќ��ņ��_:�CR��߁?�Rg?r㼽oj?�ˆ?�'@?�>?0#h>N9��NԾ�I��.ps>�@"?�u�\eC��6'��J��?k�?H�>o����Fƽ�����<���?�	\?�)"?0!�pa�,���b��<��a�
��;>��<m�}�Cr>=�>�Ҥ��g�=��#>ǭ=�[��c3�� ='��==�>R�=/<�9��3,?^\�����Q�=�gq�6xB�0>� I>���>e[?7�A��}��_��!J��/Y���?�?�?9��[g��\<?���?Y�?b�>Z����&۾�jݾ$�t��yw��A��v�=���>v��A羆������/�����ýQ�s�f2?��>8e&?wg?+k>��>$��[w2��#�n-�q���RO�|�%�J�"񑾻�n�>xC��ֺ��d��2��>(?��L�>W[.?�x>Ut$>2��>S����Z>��c>�F?>���>�B�>��>���="�<��V?R?�����#(�l%�AJ���A?�Jc?f@�>c�d���� ����??*�?��?7�v>�th��)+���?���>z/��z�
?�6C=��k��<z����������}�п�>��׽�8��L�Oc���
?��?_�s̾�oݽo!����q=���?�(?�*�5R�/�o��W��aR�v��ߩf������$��Rp�D����!����m^(�B5(=`*?0�?k�9��@)��Ǖj��p>���j>'��>��>���>�HF>g�	��2���^��3'��������>�R{?g0H>L�l?wI)?O5_?��=?��>���>��E��g?�ŧ�&A>|�>�E?y�@?@2^?*#?bm)?:��=ϙk���
�u���<�)?�-?��?U��>��>�R����νQ�����X$a��A��[�Jh=H�+�L\+��_��=l-?Cg����o�p�L�'!>9(?y��=���>v���e��>�j�>꿺>=i>�
�����UmO�43�>���?߽:�d�=#��=;Q>�%t=�����:�CB�"��=��=�>E���M=�v=u>�#>��p�B�8>0��@���?n��>��>g,�>��}�Jà�%����O=)3�=,�׽8�=ƈN���� @���_� A�>�}�?�?��޼ ��=C&>�þhHҾ{����j����^�m�
?��$?��$?ύ�?|�?��j?�>^�����6��N��� ?!,?��>����ʾ�𨿯�3�Л?Z?�9a�-���8)��¾��Խ��>JZ/�#.~�����D�����]���r��?��?{��?�$A���6��v�R���
Y����C?5�>`W�>��>��)�S�g��!�2;>g��><	R?ۻ>>�O?�6z?C[?��R>��8��!��zș�_ �߼#> �??h��?Ƅ�?�Vx?��>��>�+���߾U���>;"����~|���R=�MU>��>l��>Ӽ�>�U�=�aǽLﯽ�C���=�'\>j9�>W��>��>�Mz>�>�<.�C?�y�>b����1�^c��~���Ƈ��s?EQ�?�,?.H=U����D�x$��k	�>�E�?��?�(?"eA����=��ļOO���4y��v�>l��>my�>4
>��0=�C>���>�b�>�	��G�>�B�F�h��?@F?I�=��ſܪq���p������4[<�
��#�d��є���Z��̥=하�!c��ϩ���[�hˠ�󈓾0̵�����>�{����>_#�=$��=U�=�/�<�(̼(�<m K=n�<<B=4o�Vvk<HN8�ۡػ���T�ũ[<FI=��ʓ˾΍}?>I?9�+?x�C?��y>�m>ŗ3�뙖>�S��y3?�V>�}P�{���n;�'��������ؾ;{׾��c�i՟�,M>��I���>#H3>i=�=���<���=�Ds=���=� O���=g2�=H?�=�J�=Q��=��>g[>�6w?X�������4Q��Z罦�:?�8�>`{�=��ƾo@?y�>>�2������zb��-?���?�T�?@�?Ati��d�>L���㎽�q�=N����=2>u��=u�2�T��>��J>���K��=����4�?��@��??�ዿТϿ5a/>��9>��>R�Z�0���e��/i�>_\�R�"?��7�Wyƾ�O�>ߵ�=��ྫ�ɾSr= 01>S%b=����Y��=�G��,�D=�a=�>\|@>���=!G��!�=نV=���=��J>3�;9�9��n.�;�>=�=�=!C_>�#>�'�>Ď?�?��J?�%�>;���  ��ξ͖�>lT%>s��>�)�=��">fV�>�Y"?7;.?�l,?�+�>Χb=�=�>e�>e���$c��(	�Tr��rH[=z�?��{?_~�>�[�5���|3'��V��2��Q��>�Q6?�'?��> 0����
C���"�A�潝=t��=�h��Li�+(�=��B�~�B�HN->�z�>s��>��>��o>��=V�(>*�>.R>���px>Q&���ļ��N�v$��E�:�;u�=X�f����5�.C��c'Y�䰂���W�O}ؼ��C��ׄ=�R�>�5O>Ą�>ã�<Td���>��C�TK���>B�̾��Z�I�L�,ꏿ��C��O��cnD>�}#>J������	\?�L�>Ƌ�>���?�[o?g�>yڼ�l��ԕ�v	��膾��<��=��=�b,�/�N�ŞQ�i%ȾY��>���>��>`m>�<,�.�?���}=�6�	�4���>�ዾ�1"�����qq�f<��m����`h� �ι�dD?����Q�=��}?O�I?��?4S�>������پj�->с�Ύ=���q�&_��r�?�'?��>^E�x�D�?r������5��>�fB��(X������m.����< X����>����Ἶ�7�*%���|���w>���k�J9�>|@K?6X�?�Wn�:l��zL���.����?S&t?-�>~�?�?�������08���/R<�hd?#��?���?�_�=���=|�����>^�?�D�?(�?XQy?��=����>�E�<9�>���$�=��>�r�=�=$�?�e?+?�����=�$��B���<H�ƃ"=�ڤ=��>4�f>sg|>&�=��=$��=�.^>�(�>�Շ>~E^>���>D��>�ȶ�ʉ���a?bIt>
��>��1?9�>�
��X$��a���k�ٱ���t���m�	pֽc77=�T弸&g=5�vc?
����{�?�=�>Ҿ�-;?'b�(��)4[>R�->v�k=�H�>=N�>B �><y�>5Ǚ> S ?[\�=�fl�;� �-_����>Vf��;t�{����|<�*��1/>̎������<c��3�پ��Z�7�y��cC�aCB;�n�?����m�a�Q��J�=w�?��>��a?��s��ʅ�Y!
?_;>��1=ѥ��ݱ���*�����ˆ?J�@z��>��>>�?]�2?��^�]��>JGO��tn�>�A��Am���z��J������`,��Vn<�ދ?�-�?�O�?�r���?�>�B?�~c��+߽W��������"=�[�>h�ԾU�_��������6��r�=���?���?�.?8��M����>�qL?��?윛?��{?�zr?/\�U?�/�>-�7>���>$�,?$??r�?���>�ba>�����.}�P�۾�Y���@��2�>�*>qx3=o��=P���~�>������r=Q����1�<$�ս)|��/�<D�=�c.>ɦ>(v]?pM�>��>Ex7?�P��a8�H���l/?��8=?ׂ�=���a���5�|>��j?f��?�wZ?��c>��A���B��@>�#�>a�%>"�Z>n��>���|E��r�=W>Q�>�=P�f|��M�	�HP��s6�<�,>aB�>�"�>
����(>i&��~j��DX>lW��1����L�Q
D�H�+��m���>E#M?
?�2�=,��n���5<e��I)?\e>?��M?d\z?P�=�B߾�7��PG�/\���>�B�;.*	�LТ�"��|�8�bj�;��x>f𛾠_����E>a���hپoi��m�����v?=#�&�'�9>L-־����T�u�!>Mi>�K¾�G"�`č�����Wzg?�ʍ=� �K}����=">Y}�>���>�
��nbs��z�Ь��2��=;�>EmP>*�|�?���:��aվm�>%D?-�\?��?��t�g�o��PF�}����������R?Dۧ>��?a�A>/}�='���,`�*t`��^C����>���>O��#�I��ۗ�����I&�'�}>6w?�3>s?VV?I?`f_?k�(?�R?`@�>�ཽ����7&?�}�?|�=��ӽH�T���8�� F�o��>�)?��A��7�>~?u�?z�&?y0Q?(�?��>v� ���?�#��>�N�>�W��]��E�_> �J? ��>�(Y?8Ƀ?l�=>b�5��碾`�����=�O>��2?&#?M�?Y�>��>����GҀ=��>}c?�0�?�o?���=��?�+2>��>z�=X��>2��>?�OO?�s?��J?��>=��<�+���T��1ps�Q����;I|J<v�y=[���t���0�<$��;n��-��z�񼍧D�˚��>��;�I�>�Q�>�>���<>��־�D���B>�"<�8���a����:��=��W>���>�]>�p���=���>%��>!���D"?�?�?�'�<�i�?����H�|�>�"3?q�d=�<m�4n���ـ�e=�*l?��[?��\���QB]?��Q?��;H�K�����+!���ٔ?��2?����7�>9�_?��m?"�?K���`�?�aԊ�h%a����홶=7O�>��.�����A��>׋0? e�>��j=?�;�������V��e?�#�?C8�?7{?5�=������Vl��QY����]?	m�>�Ŧ�*�"?;��(�ξ�ꌾK��d�ᾄ5������p8������ $������ؽE�= Y?�os?�q??_?�� ��{d�ME^����]<V��|��<���E��E�tmC�x�n�Hu�#u��DI��5;=�]����A�bh�?�'?6�/�O_�>:���61�hξ8�C>(p�����i��="d��-B=�p[=QBg���.��P���X ?,�>\B�>y<?#�[�q�>�C�1�ʻ7�������4>���>f��>E��>��_:�..��꽾�ɾ ?���z׽�>v>�Ac?��J?�^n?N���1����/!�'%"���XE>�>-&�>tY��[�B�%�@�=�.	r��`�g揾��	�~f�=G22?H�>�S�>�#�?�?��	�~���5_w�ȷ1��1f<�c�>Õh?���>J��>��нU� �al�>�2i?�8�>6;�>� ����#�I�l��ZV��8�>{��>��
?_�\>��H��R�����Ǟ���P#��Z>2Xe?ܩ�h�G� :y>��F?��<�-���>�Ҽ��.�;%�֘g��=��>r�b��z>�k��>⾪�m��e���+?�2?V����0��I(>��;?l5 ?F��>4��?r�E>?Ծ�W���2?�UM?3�T?�t.?�D�>�tϻ�[���Tؽ����� <ľG>�o�=��S=:?s=�o��)����D���>M�+=qh��ZW�uG<=�X?=ev =�l��L>��Ϳ}�P��$����뾤��Ą��������3 ���B=��Q1w�ꂾ��m�D<��=�Xm#�}ћ������A�?Z/�?�(���8��=֪�PȖ��t�ԝ>:*��?������=������f��^�����K�Q�O/��h���'?N둾J�¿�q��7׾��>�*?���?W��
��D����y>_���#1����CF����ο�-{��Tl?�c�>;�澶����>��>Llu>�rZ>~���A�>|����>��1?���>Qx����ʿ+ù��+T����?0�@PzA?��(�Ӻ��U=F��>��	?e�?>?61��7�����?[�>�7�?���?��M=��W��
�yse? �<�F��1޻�#�=��=�=��	J>RX�>G~��PA�0cܽ�{4>�ԅ>�"�ʼ���^�ꆾ<:�]>��սs��3Մ? {\��f���/��T��'U>��T?�*�>l:�=��,?P7H�\}Ͽ��\��*a?�0�?��?�(?Cۿ��ؚ>��ܾ��M?YD6?���>�d&�&�t�]��=8�����n���&V����=9��>o�>ς,�݋���O��J��Z��=T� �\ƿ=��_:��H=z+�<���U��H�=���%<����ߡU�Q��"k�=�H>�C>Z��>&�>9N>��X?�zb?p��>U# >u�+��줾�:Ӿ�H>=�U���O2��L�r�c���b���Pپ�t���7	��,���þ:�:�YЊ=rO�sE���$�sg��qG�z(,?�>E8��^I��,<p#Ⱦ��R���G���5;li0���q�j��?f�A?���twV�s���R �g楽M�V?/����;�	������=J��F=H�>�G�=_��;�1�znR���*?=	 ?����̍|��>�{'�ӻl<�c ?>?�2=5��>7�)?��2�2W���{F>z"5>�B�>�C�>&�>-'����ͽ�6%?�^?\�ϽY���>�>綾��M��`�=J�#>���>���/>��$��ׂ����;W����=l�O?�{;>�.����������Q;9���?9h�>�T}>R�?]N?TF��w�ǾW�5����t�$��fI?�|?��->|!�菉6
��(�?�Hl?8��>�g�<.���]qM�F�)����>V��?m��>и�r�`�M.m��Ծ۰"?�v?1^�H����L�חU�6�>���>���>�:�il�>o->?p�%������ѿ�[�3�� �?��@
��?	K9<a,�C$�=�?��>�P�<�ƾ����m䴾4�k= ��>r����u��f�,���7?�8�?�a�>�;���d���=�֕�Z�?��?L~��=yg<���jl��e���v�<��=�&�A"�����7�+�ƾW�
�����ȿ�4��>^Y@�n�6 �>?8��4�SϿQ���Uо Dq�o�?���>��Ƚ����j��Ou�޴G� �H����:�>>>�N���ᐾ�v�h�<��"��'��>}l[�n��>- ��j���x��{o3<ݐ>��>��p>����V��~C�?���.�ȿJ؝�i� �l]?��?i?��?��<ьc���o���<bG?Fbu?�"T?hf�8O�ƈ��T�]?<�����J��d7��~S��Ѭ=�u.?J}?��.��`��OC$>]�>�4>�K9�Gƿ����m���WV�?p�?�ƾ���>���?�x?��!�Cg��=P¾�((� �<^�D?�F�>���?�+����I��?�'1?��̽(''�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>dH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?m]�>��?���=V��>���=�;��	��=�'>����s?(mS?���>j��=��4�nM+�=u@��C�����j@� �>{�O?o�O?�>�>��ǽ(M ���-���:�x�ʽ�����:����e��O�g9A>k�l>Sb�=HM�bľ8�?�W�n4ؿ�O��U(�p3?l�>��?����{��+��_?��>�T��A��𗌿�j��m�?��?#�?־�'��c�>�>�&�> |ӽ�Q���S����;>q�B?PZ�QX��d4o�H^�>��?�@s�?�i���?�����F��U�N�۾�J���_�=��?�vԾܣ'>8
�>��7<�'r�*]����^�P$�>W&�?��?��>��{?�<z��L��`�=g$�>��m?b�?]��*����=�M?f�X�������Mu?@@�_@���?�����&�����̷��ɾ��	>ž)>��>�*��.B��}>�@R�A�=�>6[�>��>��c>n�7>-
�=�|>N�}�&B-�E읿�}��Yj�����[���u�'����=��9O��Ǽ��?5��f��/����LK�k`"����<���=|�k?R?���?s�?�¼�>K��,��=�-���f�~f�>.�1?[:_?�C?���=^���h��~��θ�5���ڒ?�=@>%�>���>��>�F^<b>s��>'�S>6�>S�*=Ia�<�Q�;R >kJ�>���>h��>=>��>Q��������h���y��̽�Ԣ?%���l�I�⟕�!�������3��=v>.?(U>���`�Ͽ ���{;H?�������],���>�1?�VW?�>�d����Z���>���Tk� >|}���km�`�)��PQ>��?ork>iz>4�W~9�]�Q��׫��|>��1?�����(8�5�o�ǓE���Ӿ!JU>���>��滌l�}���N�|��
q�j�=�:?�)?M��v��-���$7��CcF>H�^>g�[=L��=�<1>P;���L�F��2B=�]�=�g>Q�?�6;>S{�=��>�#����j�ߋ�>F�L>\hP>:�:?�2-?�)���r���F����[�<)]>�>1m�>�3$>�BI��d�=���>�n>�/��ĩý[6��m�2�m�M>�ω�4�b�Z볽��2=	�LP�=�F�=&f��#k%�h��<�~?���(䈿��e���lD?S+?a �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�/)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>l��R���|܅��yp���<���>dN?�|�ꞽt�-���?T�?���e���mɿ�w��;�>E�?�H�?Ck�	���t;�&-�>D�?D�X?#�k><�Ͼ;ه�d>�:?��W?�4�>- �yO7���?2d�?�ׂ?Q�@>x�?��B?q��>�;o?�]�ſ����:x>*���>ěk>C
��p>�����db���
c��E��f,>�,=z?�>N��7��
�=���?ʾ�՞�gk�>4�>�œ>{N�>�v�>�֕>
��>�[�=��������~���:?パ?����`��.�O>tA�>��/�Z�z>�:?��1>���U�><�^?�@�?-j?�R�>3����w��j����P��W�>]�=M?��s>0�׾���=o���3T��ߋ1>���>��U>����������)>E��>�?n��>�_T>�)?�H?q�>f��>6!�M����Cx��a�>�?n�
?,ʈ?�n?�lʾ�<#������O��K�N���G>�`?Q�?��*>�'~��럿��]<��=�&�=���?�9X?��=r�?>�}?v�.?KD?7��>s$��p�eZǽAۈ>�#?$���HA�U�)����^
?��?g�>$��<���S7��X7��v�� �	?�s_?P�?*�
��T�>�����<�'E<'���!�һ��F���!>��>u�׽m:�=�}>���=k�{�L�؎�<���=V��>k��=��S�.��1^*?R��;�e����}>ɫC�FI��>�f=�r��S2?�._��≿�`��U ���#���?ll�?h�?�ݽ$7Q���-?��_?nE?*(�>�ɾ�þ�����z�A�ϽT���&N�=PH?���=�<��z���w���㍿<��-aQ��5?/^�>�$?` ?f>2ɯ>�gƾ��%�=�!��|�c��p�9��Z1��������*�q�H��k��� ���r�>�/-�Lb�>?D*?��=��>�@�>�⽌(>>��u>�[i>P��>TGg>���=6i�=b�R��B���R?v�����'�+꾨.��	+C?��e?��>:I�����|�G?"В?��?�{> �f�D+���?s��>���z
?�.=5;�C1O<�R���8�l����`)��ݏ>X~˽�S9��_L���c��	?�?�Ņ�Cξ�ؽq���o=�K�?
�(?��)���Q�2�o���W��S�4��&(h��d����$���p��돿�]��Y$����(��g*=��*?��?.��ɗ!���"k��?�`kf>��>�*�>��><mI>Y�	���1� ^��J'�����P�>�Y{?���>�c?�1!?UWU?��\?��#>栥>zɾDP�>���=�5>�� ?�E0?C<?W�G?'^?�v?�0�=����4�&Z���A?C	P?P��>���>@��>����X���=�;����)ɾ�P��=Xi�<��D��K?���=�_>r	$?�7E���@�!����<�G?sr!?�gQ?�G�
�-�l���]�>��6?r�|=W�Wb���3�_9�>=,t?vV/�ӣ�<��>1�<��e�=��I>��ƽ���=��ƞ��:�E�b>:'$��㋽�ڼ��=�:�#��?�?���>�X�>�ջ� ���a����w=Ry0>�t�= �{>�Q/�6"�L��Ju_��t�>3�?8]�?}<=j�=ǖ>{\���6������u���}���?�q?i�(?���?��4?�Q?���>R�,��Ә�1<��1	�M#?�l+?u�>I��jyʾ
6��� 3���?~=?�_��Y�`@&�k^����Ͻ>��,�ț{�����D������%��@���r�?¢�?=�%��R8���꾚ۗ�����CD?6�>��>�K�>a�'���h�\���=>���>�SS?��>�O?�Zv?>�[?PkK>x69�t��	:��=�s<�/4>E?�?���?�Bv?��>B>�Z.�lݾ���U��a��`s�"xo=85I>n0�>-�>�<�>�%>kW��5���E��"�=��M>1��>j~�>�!�>4�>@"=UZG?N0�>���}�	��̣��_|���v�q?��?`$(?Hc"=��i�J������R�>���?���?�W.?ˣM�oZ�=���۩���ls���>zİ>�>�u�=�=��>6j�>ǩ�>G����G8��rZ�A�?�B?.]�=��ÿ]���ύ�V������Y����m����g���_��=ν�WgݽlG��>�"�jS��bT�����
f��+��A��>��<8?�>
q9>"��= v�;Q �<�$�=������3=uѓ�mY�=��𺅪���Z�M�<�m�=:aZ=	꒽EP˾�}?)�H?"�+?��C?/Qx>��>p7����>�׃��4?cW>��O�ً��7�;����qG��&uؾl׾Z�c�a�����>�$I���>L>3>e��=�x�<U��=�x=]]�=�FR�be=��=Mº=r��=B5�=b->1>�6w?W�������4Q�~Z罨�:?�8�>L{�=��ƾk@?x�>>�2������~b��-?���?�T�?G�?>ti��d�>G���㎽�q�=V����=2>���=m�2�K��>��J>���K��G����4�?��@��??�ዿϢϿ7a/>*c8>5�>��R�Q1���^��d�sn[�۟!?Y�:��;��>��=b�޾��ƾjK%=��3>u8_=�����[��@�=Hgx���9=0�o=�щ>QB>M�=������=�(M=���=�cO>�A���3��-'���7=`r�=��a>n9%>���>�A?�+?�c?0N>^�����ɾ�����l�>�g�>�_?M>!��=�[�>}�?�,?�.?!>�>��y>+$�>��>��P
W� ��>����=��?Z�?B`�>�e�����#����Q�)ͪ��k�>��=?��?�L�>�e�����:���"������?>`�<E��a���d�>C�#����)�/>�;�>��>�K�>�1>�ګ��_�> ��>P�$>�k�=p�5>��=�D|�+�8�,�=��E�#�=�h�X�?����<Ŕ4��	���ݼE�'<�;�:��R���a=Ge?���>��+?�چ=�	��>�>LM����F�/�(>;.���:i��mN������E>�uu�]�M>�}8>�G���a����
?��>Z�>���?N]e?�B=*C߾�Y�v��̾����J >5#4>�� ��FF�_�w��I8�����,L�>
-�>��w>��L>BO<�RaQ�O���O���X���p>�A ��T張�!�kw`�G���0��P�Q��=-V3?lՂ�TEn>/�J?�WN?7��?2��> �y��q���h>w�C�[�)����}��5�<�3?�w3?l��>�P쾰�<�Pƾ�?��eF�>�+��9�O,���#+���q��T��Dǖ>�{о�ھn�-�Y��T퉿��7�r�]�s��>�9H?���?�T��i�l�[B�BE�+�<��>��Y?��>�V�>� ?w��j���ǖ�\	>Uφ?f��?��?)?�=tо=����A�>� 	?���?(��?ms?�?�3R�>��~;�� >����( �=>Q��=.��=Z�?��
?��
?��Ǥ	�w �)�,^� d�<���=w�>A)�>3�r>��=Fh=^(�=<�[>Z��>���>��d>w��>�>�h���ϾšV?�g]>A]�>��'?�c>�eq���Ľ�9�,�^�?Ϭ�b�>����0���8�=�!k�<j��`�?�}Ϳ&�?�=�޾e�>?���?ϯ;_��>���=�U,�
"?�.>�S>��>&"�>�S�>
��>��<>;��VJ�=�����YQ��a�n�����>�R�j���K��O.]��(��a���վ	�`��w���f2��x�BR�?��@�t���$��E/=��?�&�>�D?>W-�CUI�t~]>u�?��>NL��Z��f��^�v݆?,`@ΐ>��T>q�?�Q7?{�¼�:�=�,��r��Fp3���s�Kf�
������m$0�a0�=5�?�?\w�?�*���$�>6YU?/�[�M����"d>R��_.����=�^�=a���c���,J-������ߢ>hj�?T��?#B7?��C���m�/T+>�:?��1?�Xt?u2?�;?",��R$?I=6>�?BU?;}5?j/?��?-b2>�?�=�J�A�=���抾�&˽7�νK�7r@={�x=J�9�}�;o�=���<`���Ѽ�.9;�����!�<�v;=[�=��=옴>��L?�p?�Š>��4??y�a��9���M�?+��쀾]\��-� ��I��C>6:�?vm�?Թx?�dR>��8������=>�d>�<�=�p>�"�>�Ч���j���>�/>/� >D�=ܜ��=�����d���*���!>���>��>�J���>�ì��"��Q>��]��װ��SR���7��&��]��"�>��J?(�?��O=�����|���d�?�&?�PC?�Y?jI}?�N�qA�K7��W>�	��W�>�"�=96�!a��?���c3����<$Kz>z�y�J����5c>(��uj���&��A�[�E5	�-/>�P��+<[�>|Ծ��M�X>��P>������a����+���lM?5��<|��������{���>t�>�<�>4�d<M��2����b��=Q�>0�P>�T<���a�>�x����ɇ>59?�b?�q?����"C�Y��B��v}�|��<��?T��>}^�>W�R>��>�������$`�._7���>�P�>�#��i[�d#������ ��%A>B�"?��>B�>7|?�\-??��?��9?�2+?���>x�)�����?���?e��=��%��I����6zT��&�>+�M?�o)��5�>�'?3�%?�^?W[?�y2?">�!�6Q��ϊ>xԶ>�Ł�/���N&�=N�?d#?�B7?\��?��/>Gi5�������K��Y�>��O>e�S?W4S?�R ?�o�=���>������=,��>�c?�0�?��o?:��=d�?i<2>2��>���=x��>~��>?aXO?X�s?u�J?%��>���<�8��H7���Is��O�\΂;�rH<:�y=l��0t��L�7��<��;�m��_J��p����D�����L��; �>2+=>2����=c���U�����=�YѼ��ھq���$��B_>�x>�N�>Rx>�u���
y�u��>���>���$?;��>ƍ%?nA����s����Ğ�>�>�-?�ٻO�qً���Q�c�6>B�j?~>K?{5�������b?#�]? r�4�<�M%þ�b���	|O?�?�9G���>,?��q?��>="d���m�*ޜ�:cb���k��P�=�>����e�Lz�>A7?���>ʕb>}:�=~۾#�w������8?DF�?O�?6�?x,>��n�[9�/���t��/�]?�:�>3y��ʯ!?4�<�TϾ�������K޾�����e��Ζ��P��E%�����8Խ�2�=:�?�3r?:Yp?��_?Cp���va�+�^����[)V���`���F��D��DD��5l�C���K���֚��D=؁}���?��6�?:�(?l-�,�>u�����Q�̾�B>%x��O����≠��G:=�M=��f���/����]?��>5��>ފ;?C�Y�Ԟ;�N�2�8�7�����V5>��>)N�>z.�>P��9('��� �ɾ�K��Jν��u>d?c?X!K?ۛn?�� �P1��q���!�ٟ5�]����RB>c�>���>�V���N&�c#>�m�r���V6��(�	��<�=�2?�+�>I~�>��?�v?P��L ��q�u�@p1��y<��>hqh?�e�>K)�>�Eѽh ��@�>�{i?�\�>��>yv��<��G�|�g%�����>�ά>�z?�@g>��5��Z�i؍�xA���H6���=Ҧe?�\���]�NC�>��P?[k<��<rА>�M��2r!��`��'b0����=[p?�ΐ=�fJ>B�Ǿ�W��0}�6؆�)�?�p$?���N���m>�z?��>4(�>~*�?1�> J̾������?�z??�N?wY?^�?�4=��c������ZU=�p�>��v>�yD��'= ս�����J޽q��<��q=�U��n�)X�<i����X�=�1>풙>���uX�bWȾ�8��㾝L
������6f<(`���J�9Ĥ��!d�$΄��%��/�;���'�`��l|�������?i(�?����������㌿�� ��?�AȾ��Y���� Q��f�m��N��2�\����4fY���[��!s�nh/?�P��iĿ�Y��K۾as?D&?^f?A��ֵO��]�p��=��U=rR��L׾"B���ǿDU��A?�u�>�?���X�<��>�?��+>��c=C6�<�+���K�=E�U?4�J?\S<>hꦽ>�¿���$�j=��?[�@vA?�(�����Q=q��>U�	?��A>��/��Y�,�����>s#�?���?]F=-tX��q���c?f�<�D�eJܻ*��=��=�y=x��-K>�[�>���x�?��ܽU�1>T��>����i]����<>�\>��ֽ޴��5Մ?+{\��f���/��T��U>��T?�*�>Y:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=q6����z���&V�{��=Z��>a�>,������O��I��X��=���ƿ[�$��s�{(=v����[�y��몽�MV�����n�C��o�h=��=zQ>]�>�W>��Y>��W?Hl?x�>)7>�N潠牾Eξ57�m{���������i��ޣ�+'��y߾�}	����t����ɾ.�<�-��=��Y��9��z�M��=u��_��=C?JE	�eƾj2�e���02��C~�W^~=�:[��۾b�6�TYv�cl�?ǻB?�r���a�P�@�<�"��̪���d?���0ݾO�U�G˾<N>r=��=1��>2r>l�p$�JnQ��@/?sQ?�Ǿ�Q����0>��@>�<�J*?|>�>S
[<b��>�&?n�.�-�ԽfxV>k�$>�Ȝ>&<�>�^>���~pϽ�u?��S?�1�"���=9�>��ʾ�{��rg=�;�=R)4��D��fQ>�.�<�6����<��M��	d?<�?S?]�&>�s$�������cϜ�[+�=��_?^��>#��>#�X?-�Z?�=�=��W1l��c'�C7��wJ?̀?Nb(>Ԕ�:+���k��O�,?5��?"��>["�͛0���"�=#�0�? n�?���>�w��H�-�w�y���e�U?��v? s^�ks�����<�V�h=�>	\�>���>��9��k�>�>?�#��G������pY4�*Þ?��@���?��;<�����=�;?7\�>ӫO�?ƾ�z��N���Ԕq=�"�>ˌ��mev�����Q,�H�8?נ�?���>���������=	ѕ��Y�?��?ki��U�h<��Y
l�Mb���s�<U7�=���!�"�R����7�9�ƾ��
�!����ܿ�蝆>BS@�W�0#�>Z�7�#⿟XϿ]�� cоZqq��?n�>QȽ����/�j��Ku���G���H�Ւ��=��>��>ZÙ����P}�(2<����E>�>W��粈>ŒP�X۶�#G����K<��>���>��>����ھ�ϙ?	��V�Ϳ���O��[<W?� �?1Z�?�?H�\<�
r�$�z��
�F?{Ks?ZjZ?L�"�_�Z�b4���f?������Y�0�2�y�1�{�\>ܳ.?���>��-��"<��.>7u�>�7>#;%����a贿����?ޮ�?)C�G��>N=�?�%?�<�A9��������.�d�^��<?0nR>ӝ�?[/��:$����	
?��!?�W����'�[�_?'�a�O�p���-���ƽ�ۡ>�0��e\�$N��"���Xe�	���@y����?K^�?f�?ܵ�� #�\6%? �>e����8Ǿ{�<���>�(�>.*N>�H_���u>����:��h	>���?�~�?Mj?���������U>	�}?G�>/Dq?2x<=7��>��>��Q���=�=˜��a�� S�>��J?��>��=�z��q)�7b@���5�a���Z=����>��U?�Xg?<R,>� ���W����5��N�ۖ��ZN���h�/�Խ耚��$>�Ҁ>kC_>�(~�Wݾ��?Xq�i�ؿ(g���a'��74?ƃ>D�?���L�t��F��1_?膈>�6�G+��L&��\e����?A�?��?O�׾��˼�>��>S�>��Խ�؟�����d�7>�B?����J��P�o�bA�> ��?.�@PԮ?�i��?��)���j }�ٚ���4��a�=t�6?13�0z>)U�>s��=��v�[̪��:s���>�B�?�u�?�	�>%�l?Hdo��jC�mm0=�i�>Jpk?�z?�5�\]��B>_�?������]J�&.f?~@a�@b�_?�������g��<�j�q����7>>v�?>|��>��pD����=fh���˻P�=��>ފ>%4~>�E>U�*>�$>��z��(���������E��;ݾc_�}wX�מ��sE�����"��z�־a����ܽ��x��?0��浽�QM�[�"�@u�?��a?F�?ȣ$?.�� X>>� �X�>$���70���)>q�?A'_?�1N?_:m>�BO���V�1;����Ծڝ����>�|�;�\ ?�u?���>1!>�Ҽ>��#>^�T>C��>S�!<E�<�wӽ�N�=�!E>E��>,;>�Q�>�y�=#i���9����m��	��Waɽt��?��N��F�rlx�ޑt�Ҥ�P�>��??�FW>,a�iNп�<��d�1?z�������X=��D?Ϩu?��ҽ��^���ʽ�T��%L����c�����0��_��v�*��V>w<&?�}}>>mN>�D=�>?�ymY��b���q�>��/?�����p���z�6RG�����lo7>���>�!P��#&�V����x��S�'}H={�.?��>@b��^#��ׂk�)3��S�7>�7>i�==Z�=?�;>�ý]��>g�k�T<� >+�p>{%�>�R�����=�s�>HE��������>�֢��	6>^��?��S?��U�kIҽࢋ��X��`�3>u��>GJ>��o>�u�r)�=���>��f>������=?Yz�|�	��}>n�V='F��m�=�l>��ƾ�����u;=ST���	����=�~?���(䈿��e���lD?S+?_ �=$�F<��"�E ���H��G�?r�@m�?��	��V�?�?�@�?��I��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�/)#�iS�?��?��/�Zʋ�=l�~6>�^%?��Ӿ���>������	����6k�ů�<��>�D?�+��dI�m"�ǫ?��>��2��o}ȿyu����>���?̫�?��g��ҡ9�w��>�d�?ZK]?5�u>�H��XZ����>-�>?d�\?��>��"�bt"��g?���?sL�?�6R>ч?�v?O��>�V�<Ɣ�.���,���'=ϸ�;��>AV(=��;9�I�[��������\�v ��U>�#=���>��
�ɾo �=z� ξ�����>��e>I]>1�>�-?{��>Q��>��X=���g���R���7�C?;�?�z��f���<��=wj#��N�>�N?� =��̾�P�>�yX?0&�?J{^?f�>�׾a�����î�(�.=�5�=;�?���>x�ݽ���>�fȾ��
����>8�x>�/��щ��&漼G�>;?�}�>ગ=�| ?�?ab>�Ǯ>�\B�������E�Y¾>�E�>�?�W?�?k���2�����5G*[�QP>�)y?|?��>����F՛��b �����1n���?(i?�޽�M?�A�?LB?� ??��P>x3���վ�rp�>�N#?-���O��2�ۭn�B�?��?A1�>���rC���%����ƾ��?92V?Մ?����g�ͨƾ�!=�����Ӽ�f�<��,��'>+�>.Rͽ��z=��=���=�y���1��ۗ�2{�<u�O>��=Ȯ�����'�&?2:1:��3�+-�=0�c��(@�>�>F�~>�ؚ��Zo?��S���i��2��[������w�?��?�}�?�VԽ��Y���.?LN�?�-?��>�Ր�����Ǿ���vF��B���=ch�>:4����Ǿ臬�j��6��ѻ�������?ټ?��7?���>��H>��>+��i}-�x ����Լ��D!.��N�g�!�S���Ý�	�X��� �&��ٺ��̡�>K�0���>\��>,��=g�>��>��=�lF>�>T>>(>���>�I>�>�A>��`A��`N?�
ɾ�N%�͙���ɓ�fe4?_<]?0s�>�~�����Oy�d� ?��?�F�?@�!>�n���0���
?��?h�}��?��z=P�<G�v;&�©O�j��� �c�>gU^����^�&h��1?��?��������f`��ើ��h=�)�?�c(?�)��3R�jUo���W���R�GF���a�i���j%��o�?��`񃿥�����'�7�2=aE*?`V�?���T�����i�п=��e>�e�>��>���>��H>����?1��^�{�&��������>۝{?�6>�u?��)?�Ob?,�Q?��>!P�>����W�>wY�=��">�j�>�?�E2?��Z?�5?�M?�DD>�Gx����8�k�
�B?�'1?�?���>���>%���W����N۽E2�����`��<��:<���=fY%�%��_R���H`=&�,?������%��r�J��>a v?7?���>�ʤ�I�쾃坽(�-?��\?|z���p��ʆ� $�k�>WG�?/���c�@=H*>�f=�d��t�ҽ!� �ɂ$���뽍:A�ND=-����Z��r�'=
>�	
����Yٴ= +)�Z�?���>���>���>�BP�+b���1�L��=���>ԡ?�ڛ>�׾u��B����R����>?S��?�\�;�$r=�>9>���X���7پ(m��	�<X�U?��?x�\??�?��8?}�;?7E�>y:@�̔�Ꙉ�{q�#$�>w!,?��>]��9�ʾ�𨿀�3���?�Z?)<a���X:)�]�¾��Խk�>	[/�E/~����kD�������Gz����?j��?A���6�Ay�侘��\����C?�#�>Z�>��>��)�d�g��$�1;>Ƌ�>ER?h�>8�O?P�z?��[?(,T>��8�i!���ř�Xw/��#>�6@?���?t��?��x?��>��>�)���߾q����~�G)����bdV=V.Y>Q��>��>T��>'9�=��ĽmЯ�*;?�XU�=��a>���>��>���>;�v>��<dJG?���>�.��}��Y���}���S/���s?�?c�,?��=S����E�/m�����>,��?�o�?�j*?'�W��=Ь̼���$�m����>q�>Qȗ>�-�=x9=o�>C�>r��>�m�t���7�j~Q���?mF?J��=�\���Uj���t��ѐ��)h<�ؚ�N�x����Qu��ɬ=�˓��+��B����X���������j6���ٚ�Bh�t�>�w'=y��=H��=~&<���}Z�<��=	�=t{
=�OX��x�<�Cp���� Eս>?��"[k<Wi=�Z�;$ʾ�X|?�CG?��+?��B?E�n>�>7/a� ԑ>Y���5�?�X>�ml����ۤ8��+��;����P׾ʠ־�a��ҟ�&�>l.�,>s2>�>�=�B8<ʒ�=`�=Q��=P�E,=q�=yZ�=}��=9��=�l>
�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��#>�X>�/V��P�q����ھX>Z?��=�^Fо���>���=x���j;���>I��>geU�~�I���f���=�3��T�3��=@�>�;>���E|��q>Ҷ���=��>*�=��)��n���@���>E�=���=#��>|�?��-?Qcc?�q�>1�x�q�;aʾ�a�>���=�I�>���=?�*>�>��4?k�B?=�I?���>�X�=3��>���>͉*��jk�U[羄秾��<�P�?Il�?��>�K>=3E�~`��;�� 罐�?yX0?rU??��>�U����9Y&���.�$���u�4��+=�mr��QU�L���Hm�1�㽰�=�p�>���>��>9Ty>�9>��N>��>��>�6�<yp�=%ጻ���<� �����=!�����<�vż�����u&�;�+�6�����;r��;?�]<e��;{�=Di�>�
�>�?$��,<W��G>>�ϼ�eJ'�v>N�W�b�d���F�����X�0��9��O>;I^>��ӻN݆�i�?��>ײ�>|��?G"w?��;���G	��!
���Ǿ[
�Xl��)���>��N�]]l�(�G�𘒾�9�>�W�>$��>�n>H+��L=�Du=�w�M�3��k�>�6���B4�9���cr��o��'����yd����;O�B?���3>�|?�L?�L�?:��>�]v�h�پ�T>l���;���`Hx�&���?�R#?�r�>����D�b�̾?]��^�?u?4��0O�<��Ԧ�(�z��xw�>s�Ͼ܎�ԁ<�Ĉ�*���?8�x,�묺>tP:?zİ?ne��zPm���;����W��<E�>��H?���>V0�>�w?gO=/��i���p�:>D�?�W�?\�?��=�=�ǭ����>�?0S�?�ʑ?s?P�<�6e�>�C<��>:m����=��>�ޣ=���=�?)�?�	?&,��Qf
�w��Y��6�\�FI=���=�>��>�v>S��=l�r=F�=��W>জ>C��>��d>�_�>��>8�����a�W?��P>-h�>�%?S�>g�Y��¦=@>W}L�����.p�'K+����<��=C>'ƽ�*�t��>����Cݒ?c�#���־�?��Ǿ����>X��>� ֽof�>���=%c=�<>מ�>�>��>��+>�����:�=3Z��Y���6���S�Q��W�Y>���
�y$��#+�"��X뵾n[
��Up�y���I/�H��=Ձ�?Q���_��&��U����?��>Ч8?�d7�oٖ�xK0>�>�ݔ>���@����7��پ���?�7�?��>��V>g�}?��G?+�d����<�O�����$K1��C�S�^�v��,2��K�6�Rޙ���p?�5�?}?��{�>)�S?Zjo��<��P�>��'����MN>�/�>o�2�l�<�z���������2>���?��?E�G?�R��G����*>�">?pn-?sjw?�3?�;?����%?c�D>�� ?�R?�23?�X.?��?�79>�1 >I��^ =�0�����=½���������A=�|u=���$97:S
B=J�f<ɋüc�޼��҅ż�Ӟ<<�A=��=�C�=�c�>�gi?�(�>B֑>�j2?��0�Զ*������;;?/>���Љ�[ʚ��^���X>:�w?��?��Q?�	>�D�͂�j�5>�-�>oFa>�.>{
�>ǯ۽hþ�KT���>cE>ٔA=.��1�&�M@��Ζ��}Z=���>Ƶ�>��|>�����(>�I���ez��}d>�@R�U�����R���G�6�1�#Bv�gR�>��K? �?_��=&龬Ԗ��4f��/)?;h<?eM? �?i�=��۾W�9�0�J���ÿ�>w�<6��M���������:�0��:�s>n���J���P�> 9�_ ��������W�5��@j�%"�ig���)��d%i���ڽ�+�=b6f>!dX�(3��x��r���1|?Ϳ���$��I���վ@�(>��>ha�>�瑽���L��
�I@�=��>�/�=[���C���%8��搆>�JE?f�^?:S�?y烾�Os��;C�״��r���VYʼP�?�2�>$D?P�A>�ۮ=�!��/���d�!G�´�>�^�>���skG��M���� �$���>u+?��>b�?�9S?��
?�_`?��)?�?��>�l�����3B&?���?��=vս�T�C�8�=!F���>ߌ)?kmB�#˗>W�?ɸ?q�&?�vQ?��?o�>� �(4@���>i^�>.�W�h����_>6�J?>g#Y?D΃?Ҷ=>L�5�UϢ����-�=/$>��2?#?��?
��>ǿ�>����k�=�|�>+�b?'3�?0�o?��=��?'�1>���>���=���>'�>��?�&O?^�s?2�J?���>�	�<l쬽����tr��O�.�I;��B<zbz=�����r������<���;���������^�<G�kٌ����;5��>J,Y>��IG>����^��K��:�<;@o�]o�iJ��.��=s�=I%�>L�4>�&N�\_�<�R�>,�>�_���
?�I?�*?QӲ�]�#�پH�V����>�@]?Tg>�RO��ܖ��}X�O�=$p?�{k?|{����Z\?m�P?�~���S\��b����o����l%?�&?�~6�]�>�mX?��m?�'?����{.�?Ǐ�G�u��?p� #~=��>'B�j	c��3�=�*>?��>fCνG�=�;	�i[���H��r*?���?�Ӵ?���?�F=ye���Q�L}���H��4^?��>�>����"?����T�Ͼ3K��r%�������u��F���w���$��ۃ�=׽1�=��?�s?�Xq??�_?�� ���c��.^�{
���hV��'��$���E��'E�d�C���n��\�B'��7���G=����?�@�1c�?]'?��.���>|O������˾E>fp��?��.>�=1����H=e�]=`�g��w.�
����?��>���>B�<?�[��>�1�:�7�g}���n3>�]�>���>��>���:��+�|X��ɾz����ѽ�*v>:pc?+�K?��n?�W�2#1�2����!���.��Y��E�B>�R>%a�>��W����(&��>>�W�r���������	��7�=��2?3Հ>ڑ�>�A�?�?�o	�;����9x��1��ށ<r��>��h?�W�>��>�Oн^� �K��>xl?���>�K�>�΋�k\!�0|��bȽ@�>(t�>t��>�p>am.���[�Y���V��3�8���=�h?�̈́��N`�9<�>��Q?ce=���4<��>>�z�aw!�p0���&��>)�? ��=�:>�þ]���{��[����)?�?tj���0�H�f>$?���>���>�t�?���>s�ɾ _���?@q[?�JI?~(;?���>w��<z޳�(IŽC1�� �<��}>�<`>���=��=�+�g�F�C0.�hB =�@�=�@ȼaҽ�:�f��`m�;��5=3�2>�῿$R�Y����� ��p�1v�st��< ��S�	
��aI
����CY<Iݿ�������̧���?��@H��G�!��6��b���Z$��Y�>������l��κe��m��������U�4m��P�S��=�CxL�/?�A꾴�ǿ�ӫ�Ƹ��%?��#?�so?�~��$B�q��U��=�>��mܾp蕿��ɿګH��_V??�>�{�\;��V�?:ߠ>�Y�<�x�=x�f��2�Ne�e?�}?L(�>M�ǾW$ѿ���ƾ����?�@��A?!�(�zA�|�N=j��>f
?]�C>/�+�Y��8���S�>�K�?���?��;=��W����(e?*<|ZE����9��=Kn�=�=����H>�>��\]>�|�ؽ��4>���>N���(��8\��_�<�wZ>�Ͻr��3Մ?({\�uf���/��T���T>��T?�*�>s:�=��,?Z7H�c}Ͽ�\��*a?�0�?���?B�(? ۿ��ؚ>��ܾ��M?QD6?���>�d&�&�t����=�2�'���I���&V�D��=k��>m�>,�,�����O��K��,��=��a�Ϳc& �<��� ;NGX<��d�q/��ȴ�%*�;����S4S�hBg���&=O��=��_>?'v>>�8>(>�Df?�e?���>O:>�]����t�ң����=�%��F��8�(u������׾���w�ﾲr �M�;�Ҿ��=��v�= T����V0��0q�W��?��=�NȾ�;�x <Q�������p<��L��߾U+��.q�բ?_:?Q녿�OE��w���:���ܽ),C?��۽�y��r��1I]>[S�Z�Z=���>�o�=�/վ�-���X��L,?��>ɫ��EJK��+�>d�!��t���=?p�
?@�B���>�8?��M���2��1�<�~� �D>�	?�N�>g�Ⱦ�&�;�?�TF?Y���]��eν���;����E>�>P���.���a�>{?��.�½N�/�����rD��L?��=���[��C�����!���%�t?ȇ�>Bj>��e?1�?�d��/�1�u���"��"�=LU:?ByV?�:;>=VK�EO��*�Ut?�2�?��>�>��-��bN�(���]?���?�>�1w�ҍM���]��0����?,�v?o^��j��!��:�V�G4�>�m�>���>��9��y�> �>?{U#��L������G4��˞?�@ώ�?	�;<TV��~�=�-?�<�>%�O�.[ƾ ��� B��9`r=;�>_~���`v����=,�6i8?y��?���>���̥����=�ٕ��Z�?�?x����Cg<T���l��n����<�Ϋ=��F"������7���ƾ��
����� ῼʥ�>CZ@�U�x*�>�C8�Z6�TϿ(���[оzSq���?N��>e�Ƚ����>�j��Pu�a�G�1�H�¥��I��>��>�4��H��?�{�,g:���a�>�e����> .P�=F������3<B֒>EB�>pă>믽�"���s�?j��1 Ϳ��#{���X?��?���?�o?9�(<Y�z���y�KF��d�D?x�r?s�X?o���U�̦3���d?�)ƾ@(h��/��g,�[�=�1?�#�>(�+�(5<lGo>�}�>�k >(�)��¿�������?���?��c�?%�?��!?B�*���K �,�(�j;��0?�,Q>�1��A8���&���½j�?�%?��"�M�:�]�_?+�a�N�p���-���ƽ�ۡ>��0��e\�'N�����Xe����@y����?M^�?g�?ڵ�� #�f6%?�>e����8Ǿ��<���>�(�>*N>fH_���u>����:�i	>���?�~�?Qj?���������U>�}?^o�>(V�?}N�= ?���=�����ӈ����=K�=��ʽ��>��Q?���>j'>9t�/���B��uY����lL�;C�>l+h?n�b?��S>����C�,������Ͻ'�<�lE;��B�Q9������A>�~>�A>�/ �F���1�?�p�ٖؿ�i���n'�D44?���>��?r���t�H���:_?\z�>�6�%,��$&���G����?�G�?��?۸׾�:̼!>�>OH�>
ս��������V�7>$�B?��VD��=�o���>��?W�@�Ԯ?Zi�~�?)��喂�y�u�}�ȸ#�۫�=Ej,?���H�{>$�>ו�=8�u��ԩ��m�]��>���?c]�?�s�>X�p?��q�f(D���4=vH�>ˬg?ѝ	?�z �O�SE>A
?�4������P��i?��@E@�je?5����hֿ�����M��������=v��=��2>��ٽ]`�=R�7=(�8��9�����=��>@�d>.q>M(O>-a;>Ó)>���,�!�r��1�����C�������Z����Wv�z�
4������5?���2ýEx���Q��1&��>`��g~�-�?��H?���?��?�V	=��^>��k�*>ގ��Æ���>oS?���?�Kp?z�A>�Н��߈��݃�?2��Ӄ��� ?��+=L�?_�>O�>s�<�>�۴>��=�5��L��� g�3�d�*/<�>k��>`�>�SH>L�	>"��������co�s���E�ƽ��?ƃ���2F�͎���ۄ���˴=X"*?���=Xő�Y�̿?���SG?����*��n�L���>�L5?ZZ?�f<>4R��p�=�$3�=԰��X�qD�=�9��X{��$���Q>�h?#�h>��q>l
4�9�$Q�4I��QO>C�6?���?�9��t��UH�e�ھ��M>)ݾ>�c�&������j~�ddh�p�o=yt9?+u?a����R��
-r�#����SW>� Y>��<累=��O>,�o��]����G�;2=U��=^>-�?���=/ZA>V�>!i��Q
����2>�c�>��>��x?�HO?��Y�U�vC���1���io>gm�>%J�>�>c`��v=�%�>��Z>�M&���R��#d�`�j���[>����8��w�-�A�>�����=}7>D ���������~?���>䈿v뾵i��mD?�+?��=ѷF<n�"�. ���H���?!�@�l�?��	��V���?|@�?�
��A��=�{�>�ի>�ξH�L�k�?�ƽ�Ţ��	��*#�1S�?V�?��/�%ʋ��l�?5>_%?M�ӾMO�>W}-�[���N>��܍t��Q�<:�>�I?S��Cs���"���?���>�����2���ƿk���>\t�?�w�?�e�����T>����>{��?��d?!�f>}C�������)J>�<?��b?�$�>����&���?eh�?��?4I>)��?�s?ak�>�.x��\/��7������S�=r^;(q�>g>]���cdF�?֓�Ng����j������a>�$=Q�>���0����=h!���H���}f����>@Fq>*�I>�X�>�� ?l_�>y��>�=�;��~߀�F�����=?��?��&��Ol�Z0�@�>��:�p��>�~>?"�F��:	��ν>�f?��?��o?{��>�����+¿���V�=א�>O�*?��A>ZK����!=�Ӧ�]𶾬��<���>�	O>�Ѿ�[��fN=7��>O�?z��>�岽��?�-?Պc>�M�>��6������a��m�>`?�"?\׎?��? �l�$�@z��l)���C��(R>Gq?�?��B>�A��c���$��#����?��N?Ĩѽ,#?��i?v�"?b(?5q<��K���e=���x�>X�$?K	H��tK��:��tc��a	?I$?�p?j���ϹK���h߸���?%DS?m�
?���X��%��� =�ᑽ/GM�0�r�Q�U=$,�>�3>���GMT>'u�=�bT��e$��	ڽg�8����=Ӄ>v��=�ٽL+��U=,?����㸽w0U>h���eE��d�>�{�>v_�E&y?�9W��l��f\���������*�?<=�?ƙ�?X�!�[�I���?��]?g?� �>����\��R�+��xtd������=�}?-v>'���ᶿ婿W����p���=��?J6�>�?��>��\>4H�>�/�����RA����y/_�7�U{B��01�^^�o���rz(�K���^̾��R��>��=�b��>?w�c>�O>ޭ�>��>�I�>�{>�b�>��>�>��>���=Jq��:w�t2R?x�¾ث(�0��4Z��`�A?6e?!]�>b�g�w����+�O�?�^�?�,�?��v>��g��a+���?Փ�>Y�}���?M�'=��m��͸<�!��4���R�� ������>J���7��KJ��i�� 
?t�?͜��7�Ǿ1�׽XN���m=��?��(?�)�.R�3*p��MW�cMR�})��Ge������?%��Np�]Ï�>��F���oT(��@,=al*?�Ɉ?���H�SZ���Mk��>�=g>{��>/��>Φ�>FLJ>�%
��x1��^��'�-�����>�z?݅�>�I?D<?ZpP?��L?~Ɏ>��>Ys����>�s�;��>���>G�9?_!.?hT0?]]?�G+?��a>����&��q�ؾ*�?z�?�`? �?��?���-v��dَ�զl�?�z�M ����=s��<��ؽ�r�\uW=.%U>�M/?a<۾o�%�u}��- >��u?�9?�7?|��#�.��8>�3?%�'?ǐ^��.��ʊ�����5�>8��?���(��=�l.>Vh\>LX�>������.Po=��>ه	>�s<��.>^F�=1a)=V5B��>�=�������=#@=c�?a��>W[�>G��>�z��>����*�rs=>o?4>2��>R9p>N������~��G�e�>���?`��?5�����=��M>o��U��὾�
��K�彵��>�&>?~�M?Ӎ�?�+m?�>?��s>�	�+9���长8P˾�4?t,?Ϟ�>���7�ʾ�騿��3��?NK?6a�F��-3)��c¾��Խ�>�D/��~�� ���#D��Ő�a��hE�����?�ɝ?!�@���6�d��>����f���}C?��>{Y�>��>��)�T�g�;(�b;>ʚ�>PR?�#�>��O?!;{?�[?�gT>�8��1��)ҙ���2���!>�@?���?F��?�y?�o�>8�>��)����O�����,�݂��W=T�Y>}��>�'�>��>a��=��ǽJ����>��M�=��b>^��>��>��>πw>�:�<��G?Ѝ�>�c����tr�ہ|��V�<�,a?:`�?K�.?���:p*��R^�,��\�>���?��?x�>?>�?�
�=pJ�F�˾����ī>� l>�_�>0��>��=��>�x�>�¢>�B���.
�&�L��G�@�?k�-?e�=:�ſ�;j�yL�/���>>=�Ӎ�-q�K췽�Z�]��=�$���1�e���M�J������U���ş�3{����>�4=a >L�=�ߣ<���w��<��=_X�<�j=Լ���P�<P�!�� �:�+��/�k�t��<�n=�v�g�Ѿ�~?�J?X�+?\�F??�v>4!>C�g�C��>�I���?�P>%�[�x����*�xʥ��ޒ�1�۾]վ"�e�F��S�>��j���>��/>b��=!.�<��=�j=sߠ=�4n;dl%=�w�=��=�^�=��=j�>��	>�6w?V�������4Q�5Z罠�:?�8�><{�=��ƾo@?X�>>�2������}b��-?���?�T�?L�?7ti��d�>K���㎽Uq�=+����=2>`��=��2�d��>��J>���K������4�?��@��??�ዿ̢Ͽ6a/>�aC>;�=g7T��5��$q�;�[�s�@�E\&?��;�Ůɾd�>�Λ=s�Ҿ������<=�
%>��=�j �Y�V��֞=�8��|�(=��$=��>�Mb>���=�`����=�S,=d��=gW>��<@�m�� ȼ�� =&_�=]k>�'>���>\�?\�-?~�a?l��>	���8ؾ����a�>�y�=�ٹ>�oq=ǯ>a�>��-?�@?��J?�C�>^�=��>@�>x#���j��b�~5����=��?�t�?���>��R=%�[����I�=����v�?��3?Dt?~t�>gI�I�7����)��M2�ړ<��F<l,��m���Ȓ<ˊ'�p�$�h� > ]�>Ï�>_O�>�/z>��.>i3,>�u�>(�>�4���=4�8�B��<	�=ʗ�=�ƀ����=PHB=L�½���<ӯ!��b=��k=e�2�
N�͡j��=�?�P�>�?�kǽ(���cgo>�]۾WF�� �=����N��)P�����M	D��-ν�d.>)�w>
�¼���e9?�.>#��><��?�@w? b>���<>޾h��d[�����]��=�_=���&�=��Nh���[�w(��m�>�zq>x{>ɎQ>mR#���=�����?ƾ��4�(�>%#Z�j���R<���g��������
�i�*��<�E?ȷ���6>�*�?�iM?9��?�ڶ>�N6��/�m>�L��W�=(����.!6���)?hI/?c�?bQ����P�i̸�3�ӽ�<�>�PO@�L����&�y������#�>9��r@پ�5�Kf���N���u0��:�(��>_D?dŮ?����I#u�ZE��s��8�����>�T?7ݕ>�v?��?����q �b*��W>��?|j�?M}�?68�=���9��*o?u�>�o�?�H�?�g?a�S�<�?�5>���zf2</�<>�t�>g>� >� ?!��>!�>��	�����������W߾������}>��>1�>	�k>��>���v��=�{�>+i�>���>H?>A��>Ѹ�>y_�q:��cm?[e/> ��>��<?�(m>�q���6�
&=�jždC���l��@����=�'�<�p�<�A��蕞��
?stͿ8 �?=p=��d��?J[���a����o>�x�>)���� �>%�>=��>4f?w�>׵�>���>���=�劾�=��+��-��Bo�s�U�<�̾O	s>#?����̈́���S�T����j�xN龬�V�����r)A��I����?K&���G*���B���=��"?��?�tb?�|��ߨ��У=eb�>�9�>�!��������yҾ�%w?�;�?�3�>��*>��p?:�??�yӼ]��<�v������9�T=�hm��^��'6��~U$�jf;>-�?��?ԏv?ꚼ4'�>SE?�s��̬�b��>w>5��H��I�>��d>@je��P�r�������4�Rta>�N�?��?��>?��RE���O�>̓M?�
1?9&�?3�?<H?�����\O?�A�>U#;>�=�>\-?�:?&�+?�z->]~�=�@<���=�����C���P�5��k����Q��ؿ���.�o9���r=�/>��I<a�C��_����=xv�=����A��)L�=j�>��Y?J��>�>��7?cz"�]�7�*���"�*?�ZW={�~��s��:��y�=�j?Cc�?9�Z?�(X>�A���;��>Ԑ�>�#(>��]>ۨ>����I�el�=y>�t >�v�=��*�ꍁ��2�������<�>.n�>-M�>�����8)>�9���W��i)>�q�Ƚ�b񂾯@���E�>�)q�>��O?�&?�FE=���-�/�am��w'?�'H? @j?��q?�B=�5侗�8�e�I�c\F�Rޘ>���<�����ॿy��5�=��Q��h��>��~��1l�>�� ����S���N�h���]ƽ�����=��<r��e�۽k��=�d>1n���$&��L��u�YU?!�G>(쾇Â�t��~��=#��=m��>x�=~zN���<�?����i���>O��>~.̼
)��^�Z����%�>ag??�v??Ж?�<�H�]��s�^�����;��.?���>R?��>�@
>hkx�'T���4C��AU�$3�>��
?��D�<���:����H���S�>��>����[�>R5F?h��>�{?�I?e��>[K3>���1 ���s#?��?#��=Nh)=C����C��!R����>Fg?�);�䉵>*�?� ?��8?f�_?> ?jy->A���ۭI��=�>Q�>��b�P���:˦>C�O?�J�>	B?y�n?gNY>i+�>����6}��e]=v08>�=?95*?a�>�V�>��>�˾s#�>�x�>@�Y?!#x?w5�?Yԍ<DE�>3�l>���>��:��V�>�? �#?AdM?k&�?�h?��>����A������X���=�54>2h>�\
>��<��� �(=	:>([<���*8>�F���iD�HƲ<2r>�0�>b��>�����>?��~﴾�p�>T輎"徂[N��O�>�e>�9�<�g�>O�>M^����=���>��>Q�#���?w ?��;?޷>Uh��I��W��.��<!CE?�V�=��������P+�1>�w? D?�5;ӎE��b?��]?]h�*=�s�þS�b�f�龑�O?��
?^�G�>�>��~?>�q?��>��e�):n�����Cb�e�j�UӶ=vr�>X�l�d��?�>�7?�N�>��b>A�=u۾��w��q��z?��?��?]��?)*>�n��3������H��t�]?Ik�>05����"?PZ���ϾZ������"�_ ������=5�������u$��܃�X�׽���=��?11s?\Xq?��_?�� ���c�@%^����3pV�.���ԾE�w)E���C�D�n��]�4b��j5���ZG=M10�x�8���?_�B?!0��0�>H�����ھ�������> ���/�����:>��=��<�1>��F��i�=�/��?�<�>Y��>��n?Q�j�,�R��`���_�LN���g6=q�>�1[>ƾ?i�K<�4�<��=�lžO�x������v>�Mc?2�K?�o?�6��1��:����!�D-=��ϧ��F>��
>`�>�DV�m���-&���=��r�����됾��	�,�=�2?迁>��>��?�?�	�$��P�{�:2��̀<=�>yBh?��>���>IvԽ�!�M��>�g?��>�ފ>�݃�<&���t�4�a}�>��>[�?�֙>&%u�G)b�����^"���3��>�Ud?Z�~�s&5���b>=B;?q�<��A��݌>QI��y#�w�;)�颏=n��>\ގ=/!5>�þ�w�e�
��'?l=?������*���s>�*"?Z��>A>�f�?��>	�ľ�+�;^�?�^[?hTH?	�>?`��>&W	=����-ǽ�2#��C=E��>	hU>ҟZ=��=�d�W�T�~N���-=&�=�(b��Iӽ"ig:��ʼV(�<Q�=ق2>-ؿ�DH�hپ�%�����|�������S��̾g9��F�.���MR���]�D�g�t>����n�jw�?�6�?A8���{��;���}w�y����Ǩ>���=(�����Ƚ몦����<���D�A�a�P5k�Y�Z��].?��f�k�¿�ȣ��쾨�3?�t?�7{?y�2��:�8�%�zG>��="�Z�Bϕ�\�ɿ���H�P?��>�I�b�׽h��>LJ�>��>y��>����.�?�?���>ڵD�Gʵ�8ᵿ��7��?�?;v�?�cA?�:(�^�L�X=4��>}u	?5\>>h�2�T��k��/��>��?b�?�sQ=�=W����ee?��;��F��ѻ�V�=`�=Lc=�=�fK>]c�>���e�@��ܽ �1>���>k"����_���< ^>�ѽ�G��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=��#�׿����\��A���_��!�+B�g�<�^�>u�پ:��ly�;�* >ɼ����>��>e�=��>.a?3�?���>f	>O-���%�����X��Ś!������h��[��=U�w��y������6��\�-�D�.���Ӿ�'��P>�Q��ҁ�gp���t�a��	?�g�>ce����m����˰���"M��A">�$����ޒo�ɉ[�(՛?��/?k���G:�����"���*,��Z�?�)=��/�Ա��X��uQ)�+��=�U?�������,�G���N��3?B?>���'�����=��Ó�=і1?�?�%���'�>+q2?��� $��x�=�ہ=~��>~x�>�Q{>r����m�HK ?�mb?Z�!��A��i��>�ľO�l����=�g>������[�>�xV=�$�����=�b��dْ��M?/�>u�&���$���%�,�,>�û�\?��.?�;�=�e<?��k?V/D�׹5�dai���)����E?R<�?��T> a0�8���U����>ݬ@?��>�4w=b�߾�����b?��l?R�%?]Ľ|\��8it��Nܾy�h?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>��������
>����W��?枏?�ד�������,��@o��bھ�?�=�f#>�*��L�L=������*�r/��q���X���̈�>�z@
B�g�	?�P�IK�m�¿�0~�bҾ!a��ז?���>�V���w��N���p�T�T�[��f����>>�>5��R���I{�Ė;��$��ߚ�>y�B(�>�fV����5����8<�C�>�}�>�܄>|d��������?]7���$ο�P�����K�W?���?���?{�?1�<�=x��K� �7�VSG?dt?-
Y?|e9�D`�� ;��e?lG��3�@^�S�=�i�>0�*?OD�>�H澙�2��zJ>�n)?��=&M������<���Ɋ?�O�?]J���?��?Ll?�Kپ���m����N�P~�=��+?1��>}#�@�%�Rez��fT��:�>��=?#N���
�]�_?*�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?ֵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>[H_���u>����:�i	>���?�~�?Rj?���� ����U>	�}?�v�>�M�?���=�O�>���=.m��T�o�-�>t>�Y�)_?�M?7;�>B��=h�?��0�F5E�(�P�pD�\�B��ψ>�h`?uDK?I�c>Lqͽ
�b�i� ���ɽ�D'�(D��׻@��1,�5�ҽ��,>"�:>��>=�?'վ��?=f���ؿf��K�'��:4?Yƃ>�?]����t�����?_?�{�>B�6+���&���\�&��?hH�?��?�׾I:ʼ�>��>#H�>�Խ�ҟ�vm����7>��B?#�]9��k�o�c�>� �?p�@ծ?4i��	?���P��Sa~����7�`��=��7?�0�(�z>���>��=�nv�ܻ��X�s����>�B�?�{�?��>!�l?��o�L�B���1=6M�>̜k?�s?}So���t�B>��?$������L��f?�
@~u@a�^?+�~߿�Ŭ�e���������=�f�=³>J{�����o�>W�<�-����~=�j�>~�}>/Ƀ>6P>��?>{s>>�R��:�*��G��܆��C��/�����Η������=x���])��������+���y(��������6�Y=���=;�U?�R?p&p?Oa?;gy�v�>�����	�<ܒ"����=�>�2?��L?��*?���=?��Ld��U���ᦾ�������>o�E>��>�^�>z\�>���:�7J>r;>>��{>\>�0=��hx=�,M>�ګ>���>�`�>�M|>�I�>Le����hY���F��_���?��C������j�����F�*� �=LFw? >�(��=����<L@?V��7e�v&ʾm({��'g?i��?F�+>��վ����~G�>F̀>�A������e���lY ��f?JT?�7�>t�>~PJ��2U�A�f��ٽU��>/l?���������@�̨��/����=/��>�|�?�2���O� ����;�=7�E?��>�<bV��W��� &�C��>^f�>��<��C<=��>8+��V����S�R/�>�h�=�j>�Z?
8>yIl=���>Ǯ���-C����>CB>!�>>�";?�Y"?���ߠ�$���02�=|Y>��>"�j>[� >͜E�庽=�_�>ˈU>o៼H.��m[���:�RdJ>\>���m���{�i��=��ýa�=2:p=M|�K�4�0V�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ٧�>�޽�H�������q�J�=��>�<E?���\�!�C�tT?Is?�U�^}��Jſ��v�OR�>���?���?q�o����A�/�|�>�9�?czW?�=�>��sh��u�>�R0?�OG?�:�>H/�N�8����>}�?�"�?^-v>�?$1?fi>If��t��oФ�nO��W�=�۽ ��>�Y>ȯ��k(l�����dH��=�X��x���>@lN<h��>�=�#��c(j>`��;ۊ�_�`��V�>[�Y>a��=ׅ>�v�>6�?=�%�>�l�=�=+��?�΁�#�K?[��?���o3n���<��=ȱ^�o?�K4?�s[���Ͼh֨>:�\?���?}[?�]�><��h=��_忿O|���<��K>_0�>`E�>�,��{9K>��Ծ&+D��u�>�ʗ>�ѣ�.1ھG2���U��5<�>�f!?��>Nή=�?�@)?�G>���>Y�1��w��XE����>��>�?M�y?N?�\׾��E��l��i�����Z�KxP>=
|?��?���>�]��)���D	�:�'<$q��U�?�m?Ȇ�����>�x�? s-? �4?&�X>� �۾��]�4�>s ?�F��tD���*�-�-��
?)�?J_�>�0P��Z�� ɼ������HI	?�}Z?��?Dl�	�a��B���G�<� ��c�<xv���%��>	�>�ض���=��4>�=7"`���@;�i�=�A�>�>I3 �� ���<,?�eG��ԃ���=��r��zD���>�@L>��Z�^?-L=���{����>v��^U����?��?�i�?e
��&�h�t"=?#�?�
?R$�>�M���y޾���Zw�)yx��|���>H��>Ôl�L�P���p���)G���ƽ[7����>;�?�?_�>eZ>+:�>����F�w��.Ͼ}aF����p��r�%���ֲ����������D;,4l���>�Rd��?��%?�>���>�7�>O$T�}>�!�>F�>}��>�>U�_>�5>p�>����NR?ك��2�'��5��#��e*B?�d?�f�>�h�x���B�׶?]�?SL�?��u>�h�+�׈?���>�:��$b
?L�;=%��|�<����Ah����[����>\ҽ�:�~;M�Бd��
?�?|���x�̾9�ڽo����o=?�?<�(?q�)�m�Q�0�o��W��S�]H��g�MI����$���p��폿�`��f ���(�9�*=*{*?��?������+�|	k��	?��Of>���>��>���>gI>^�	���1�r�]��6'�T΃��<�>]]{?��>7n,?��J?w�8?�n[?�>1�G>S��ǟ ?[�>gt;ѣ>��9?�(?�,?�|0?�Dh?���>Б}��������?&��>
;�>���>�B?�N�?�lƼ|��=������C��J	�~��=֖!=��V���e>+As>;J3?;�%�2�Ah�S��2�Y?��>a�'?�El��J�G���W"?ݩ�>����s#1��Ћ�������>�֓?f��<d���M�>؜>Ƃ��ӼA�>T�=���=��ͽ��k���.<X�%>��=U���5�<u�>��^>�nнkt�>�?6��>=�>x>��ͦ �����O�=�Y>�S>G>�=پ�}��%����g��My>u�?�x�?��f=�=[��=���W���������/�<f�?�H#?�TT?���?��=?Fh#?�>�)�L��^��r���?�*?&v�>�i����fs���y��?4z?5L��$Q�`p"��\��"cE����=u`�&x��㮿~)G�f�I���X-���?;ܘ?@!�$X,�����o��T{���"O?6��>��>E�?wa'���r�r����>a��>�O?���>��M?-l?Gۀ?I�#?*I�{&�������འ�]>J?x�H?�?)Z�?�"?�j�>���=����7�Bk2�g����ξ�X�M��>Q��>���>��L>4<�<M2���Ǿk�	�ʇP>f�>��>�ff>g��>N�J>P�<_�G?2��>�U�����᤾Խ���F=���u?���??�+?y=^}��E�g?��[M�>�m�?���?�1*?��S�j��=��ּ�ⶾ��q���>[ѹ>�0�>�=fnF=Hk>��>M��>��b�,r8��iM���?�F?Q��=aɿ��%_�[�q��;��
;"=��Ͼ³w���M��I���,�=ھ����>�<�k+�����.��M��m�Ѿ�u�� ?��>Q�	>Ǥ�=����;.�e�9=�4Y����l�=�o˼�1>I��=Z�C<�-<�a����h5 �9T�˾yg}?d�H?2O+?&lC?��y>��>�4�O;�>�ꃽ�7?LV>z|T��d���<���� ���fؾ�׾Pd�h���Y�>��K�D>��2>�<�=��<l�=�w=IB�=�^��=q��=�{�=_��=��=&~>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>W	<>�V>R�3�5�p}�v\:���T��v?֭)��ɾ��>���=#>�f�ɾZT=x>��<v�1�8:S��?�=/�k���=<h8=��>\�2>&�=XTý�!�=���=�R�=C�R>��D=z��t�e=ԍ�=?�o>�G>�[�>�j?W�5?��z? L4?\qw�����m־��J>F2�=��8>|n�=��>2K?H5V?�C`?)`?��>Jv��;h>?�b>�y�$\���ǾE+H�Ѓ���tL?X�l?G_�>� 9�����x�
�b�K��V����?&$G?dZ?4I�>�������� �t���(�`���e>��y�I��=P�>�İ�c����>;_�>æ >�~�>�6�>'M>��O>ج�>��>=M��J�;�?G;�d�τ%��ߍ<�5�%t��pW�x5>,J�>��>j�.��=1��=�Ľ�'S��>G��>�>ǃ	?Zg����9�>�꨾m�v��=��?1>���n�&�R���%��U_��C>)�<>�K��������>�7�>I��=�?=��?��~>�d���׵����d��w-y�2�8>Ë>3���ʹ�3�H��87�����1��>c\�>��>�<�>�Q.��D;�~2�=�ھ�b6��E�>��7�|�[�GK0�8jg��ꟿ3Þ��`����<��C??����G�=��~?"�N?�׌?s<�>�yŽ6�"��=�'a���Q=����E���q���F?�@(?��>m����O�H̾���}޷>UAI���O�`�H�0�z���̷�Տ�>c���8�оd$3��g�������B�EMr�%��>�O?k�?�9b��W��>UO�V���&���q?�|g?`�>�J?�@?�$���y��r���v�=��n?x��?(=�?�>c?�=`���?k?�X?R��?�S�?��{?�B���ߛ>h��;i
>�ϫ�L<>��E>ju-=a�=C?8�?�+�>ǥ�Z������^a��4��<k��<g-�>�>���>�
>�k]=�m�=�8�> E�>�h�>Ɛ�>�:�>a	b>#��> ��u@?��O>��>=[?
m�>�}R>�a/��� >��p=l5���6N6=96G��NO<E_�=�4>+-M�,>�>��ƿ��?�bH>_/־�=�>��J��?ѽ�`�>Ee�>'����.\>0�*>\S�>��>G�?��b>���>Y�~8��)(v>�c��hF�/�E�������s2>�W����ڽb�	�V�NQ��G���k��%+g���s��8����<#�?�����r�I�&������?G��>d�T?�����(N>�>��>���̄��w��^��?\��?�;c>o�>5�W?��?�1�3��uZ��u��%A�e��`���������/�
�������_?��x?�yA?�<:7z>���?n�%�?я��%�>1/��';��<=-�>&��x�`��Ӿٸþ�7��HF>��o?	%�?5Y?n]V�ŋ��BT�=�4J?�p.?�\t?�C??:�U?��m�"?�4R>��?�z ?�
0?{�1?�$?��l>΁Q>V'�=�B�<% ��͚}���������E��	q�=�V.>�=��=Ħ`= {u=}C�<A0����*���	�:�=Sb=ļ�=R�8>-Q�>�8;?��?*��>V)D?5!���6.�+���I?�~o>!?Ǿ����zo�����d>���?���?�fe?�s<����<��| I>ƽ>��@��.�=6�> �1�����&�=�*�>����|�=��_�3�:}=�%y�� ��1>̾�>u�}>ʒ���">Q��TLv�V<f>��R��p��E�V���F���0�!�{�:$�>E�K?γ?�Ǒ=v��¶��d6f���(?�<?�M?��?7�=Z�ݾ�%;�h�I�9��aQ�>���<|���T��(F��@':�a�;Eq>�-��S����c>`���L޾
�m���J�OI��OJ=����>T=9���+׾>{����=�u>�r���>!��E������!�J?o=F�����U�"e��pf>���>��>1���y��@����r��=s��>��?>�ޞ�#��جG����E��>}�2?��h?���?�^Y�d`���_���Q�Dp����ZPQ?���>z�>��>O��=W���ʾ��8� ;@��d�>G�?e�U�lBM�^:�����H����{>�)?t,�=G��>�FU?�?~�f?�ie?r.?�\�>�i��������"?c�?Nu�=|������4���K����>+H(?DN�o��>� ?��?�?+?��U?J�?A�6>5�����C��$�>.I�>
V��#��dv>�F?Jܥ>W?� �?��1>|�6�0ӧ�,������==!>S�4?�&?�;?�?�>�c>T\��N>]�u>_�a?^f�?0�?6>���>���=�t�> 7�ӄ�>��?�+?�F?p�?�X?,�>��<t@������W��j�N3-��-��pBѼ���FHb���½��+���y��ѽK�ȼĶ��u0,�"���ȷ$=�N�>^��>�Lu�-M>��ɾk���8+>�j�ԇ�F�w�z�Խ����Ϗ>���>H�(>^n4��~k=�R�>-��>����?��?�*2?K��<�`�~;�L�����>�N?�6>�`�t����DO����=?h?t�[?�Ɏ��L�	�b?��]?J/���<��þ"c�9��p�O?�
?I�G��$�>�~?��q?��>)�e�sn�����5b��k��ö=�|�>m��d�$�>�}7?=E�>��b>���=�Y۾��w��O���$?s��?��?y�?Z*>}�n��0�����Du��<�[?�T�>ץ�E"?ª���о<���o���Y޾���(��������A`(�R;��_sֽOe�=v ?ZZr?�p?!_?B�+�c��]�~�~�4mU��� \���F��(G�H^B��Kn����s'��J˘��2?=u	���+��h��?�n?��,�_��>��������#�&6�=s��:+z�!u=<�>�R=n&o>�{��*=m��6p�>���>셡>��:?L�}�k�<����G*��M���+>2&>n�l=x��>�1E>l����ʽ�����y@��2�x>U�b?I�K?�2o?($���3����������J������-M>6
>F(�>��I��y��G#��v;��q��������� 	��?p=�4?�р>O?�>��?��?�6�oD��S�|�b�1��+v<�]�>O&i?���>u&�>�ݽv!����>�g?���>�ٓ>#���Ef���Q�b?�0��>��>	�?�`_>#>]��+V�-����"���N2�p�>�]?��p��52�q�>��=?R:�<Fҽ�P�>S)G=����E�ɫ�-=�l?!k>bq�=����[)վ��j��X�.P)?�D?����6|*��>��!?a�>�>�0�?¹�>þ(� 9Ё?�^?AJ?�.A?L�>�'!=�뱽<�Ƚ��&�l�.=��>��Z>�Ol=?��=J�7�[��|��BD=@�=<}ɼ6���<���`�R<�$�<N$4>�~��-�T��%;7����Y޾�W�ɐ���G�(���Yk�&����{�� =/�K�f��~`���?�vw�\����G�?xX@��ZOt�ݤ��>t���>�ݤ>���qA�=����&��Z�ڽ����~x���&�j�>�Y3}�����E'?�����ǿ�����ᾮC ?Q ?ɬy?���dg!��h9���!>���<>ȼ����"��JJο7�����]?u��>�\��ț��-�>�	�>�*[>�p>�%���������<Ɉ?��+?���>9To���ȿ�������<�?�z@)1A?�N*����qXh=\_�>8o	?��A>7�1�Q�������>!��?�W�?��_=*�V������d?�=5<Z�F��û�8�=I��=ż=W���K>;Q�>�l���B�,⽇2>%�>�V�F�mZ��ֳ<��\>�`׽����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=&��Pп���_(� ��o(�PQ��)^������3��Y����ϼ��%<1 �<���=l�p>�؁>!�6>|�<>��a?Bl?�E�>�^>�~��a��j{ƾUm�p���M5�y����t��������Ҿ	���K�1���/������5_�F)m>vY�U�~�<p�J舿l���,�?�?YP��\ڎ��	��c-���p��F>]�սG�̡��ҳ~�ᘦ?�<?ى���u;����� c��t�wc�?4�L=�F���վ��V��P��c=��?�w=�V���B�?�E?I�?#W\�v�w�1�@>��;�">N��>��5?��x�?I�>/� ?�h@����Ľ�����=�d?�H>���Ĺ��?�W?0�y�TsϾZ��=�/�澁��;@�?>
���\6~>�ۓ>���nx!�{t=��*�{��\R?4;�>R����qs��`x��>�NB?a|�>��>�'E?��A?3���ﾱj]�8��bP-�� C?��\?NNO>M�3���Ѿvʾ&�?�_?1�p>��>�j��� ":�t���5?Q2"? ��>�r^>ފ~��|��aI���6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?r�;<��U��=�;?l\�> �O��>ƾ�z������1�q=�"�>���ev����R,�f�8?ݠ�?���>��������>����(�?_ؕ?e�Ѿ��нJ�ND��%2���=a/>�a;�1����X"�c-/�X�a������S�J.D���I>0�@�\��*�`>e�}c�"�ʿ`�'��R2���d�f6+?ꌗ>ظt����z���{�E1�����ż���>"�>�N��ru���~��>�N啼]�>���=%{>�<���ľ�M����<���>s�>��>�æ��F����?����ȿ�˚��S��AZ?���?x�}?��?t�= ,��z-q�$�%:?II?Vx?H@^?=z�]�}�����\?�m��_o�{�E�dH��|�>ƶ*?DO�>Y�)�&�> �@�K�0?���>u�>�����q����9�1ː?�z�?g��?��>�ɕ?[t;?��&���%�����7��@>y<Y?銲>�zF�����ξA��S�8?�Y1?n ��/A�]�_?+�a�M�p���-���ƽ�ۡ> �0��e\�"N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>e����8Ǿ��<���>�(�>*N>jH_���u>����:�
i	>���?�~�?Qj?���� ����U>
�}?�'�>���?PE�=�,�>?	�=�I��v+���=��=�g����>�/M?z�>8T�=�>���/��!G��L�����yA�ۮ�>@�e?+/P?s�R>GUӽ>�i��"����*��K04�ժ4��s����:E2>�pF>FX>��9���־-�?:�7�ؿ�q����(��r4?[σ>��?�9���r���<�8u_?i��>�����;w���X�P�?�?��?83׾��¼1�>�&�>���>�'ҽŸ��w��,:>�cB?��
�ӊ��1n�<.�>���?s�@]��?J�h��	?���P��Ta~����7�b��=��7?�0��z>���>��=�nv�ݻ��X�s����>�B�?�{�?��>!�l?��o�O�B���1=5M�>͜k?�s?kRo���l�B>��?"������L��f?�
@u@_�^?*��ۿ�����r���R���+�=i�=��j>�b���
=�/�<���sp<](>� �>��s>�g|>ΟX>5GD>��$>����$&�����X���=�����(�B.:�s�
�������m���ʦ���罪D��W@O��W;�P6!�8�����=@�J?��T?Yă?$�?}�M��6�=ua��{�h��6����|>��>��>:�[?�+=?S�s>���n}O�����7Ѿ����o~�>Ѝ>��?{?rͿ>t񾽣�z>tk9=5�>I�>�3[����f��<�$Q>���>��?w�>��>f��>���Y��=~������V$�@��?ٵ=S�c�����rVl�"mx�c����p?][>�擿V8��6����D?Γ���N��F��z���h?�Շ?Tm�=�����;I7�>�>�oc����=A�ٽ�۽h�t���>3�?�c>ĥ>K�;��R?���Y�!2��*n|>��3?.ݤ����p�_�=�EѾ�k5>�k�>�Լ1�������pu��v�(��=��9?�O?O���J������0�����5>��>�X�=�0{=�n6>$���{'��8����o=��Q>��>��
?+�>�Hq�5sP>�R����`����>��(�"�c>�y`?�u?zA�� �&<BԴ�h賾�K�=��[>��`>{9>Nc��	�=�.
?猴>D� >�^O�?�M�6H��+܊>�[��8�%�<�޽06�<~˼U`��ǲ$>u >('�K�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>6v��I�s���k�s�t>���>b�?������=��m��>=�?`�G��(���ֿڂ�q�>���?��?�n�m������!~�>���?�XJ?��>��v⑾��8=֪_?l*`?��>����T���??�ɏ?>�?>���?S?nñ>{e���,�-:���"��Ne�=��>,�>�Z�=yѺ�	�F�`����6���J_�#�r�|>xc=w�>8`ҽ?1ѾD��=Ԡ��-���!#�&?�>�(X>�	T>�z�>�r�>�Ѻ>�;_>���;u!���r���X��J?S��?��֯o�d�T:1ɢ=uMS��#?0�3?%c��jhӾ��>V�Z?�K?��\?�j�>)x�b��s����7�����<�`R>Y��>�:�>�ly��oH>��׾��G����>B�>k��)�ؾ�I�������>�>]~!?٪�>�@�=�I ?&�#?)!d>34�>��@�=��'�;�i޶>0�>��?�Cy?^�?f��h'/��ђ��Ý�^X�2hQ>E�t?�:?��>���ܨ��������n����}?�\?t�
��s?)��?S�2?49?��>�[$�-��&��$s>x�!?�~��A��C&�Q�"j?�8?,��>v�?�Խ/�ּ���b���*�?^�[?��%?�����`��h¾�Z�<�����E��<�C���>@>�r��Vp�=Y_>���=�m��6���f<��=.�>�@�= �6������<,?��G��؃�F��=��r�`xD�q�>�PL>����9�^?�e=��{�����w���U����?��?<k�?����h�'#=?9�?�
?�>~M��
|޾4��MWw��~x��u��>��>�l��
得���J����E����Ž`棽��>=�>~�>`�>���>e��>��Ѿ�6׾V�Ǿ 5ξ�@C��'d�ueH��WN���5��3���H����p>�=o�w#���>�����>|
�>q�>4)�>. �>�}7�p	�=��=�"�>Ӳ�>�H�=��">�vY<*&C>��缨JR?Q���9�'����̘���B?8]d?�(�>g�g�����2��h?�s�?�]�?'�u>�mh��+�~w?(2�>���\
?�r;=`��|��<�������G�����>��ֽ�&:��L�of�7a
?�?����̾�׽�h$�=�s?S�?h(%�8�K�~�p�gY���M��]t=t.�X�����ֵj�m���}�G(y���&���=��!?�T�?�����R�X���Yh��6B�lU#>���>Ш�>���>�e>a��@=�"=a�4%%�82���	�>��?zU>uN7?��;?��L?�Bo?�>���=(ｇx�>T��@��>Uّ>x�?�y-?fxJ?�7C?�vR?��_>1��d��:�羿�?d�?�?�?	�?��]�Һ��韽Eӟ��J�� $	�c�f��<���5���Ì>� y>��$?�ޱ=�/6��o"�0#>��4?�?�B3=�{Q����	%���"?��^;��~�ᾄ(��%���>H3u?��=S�=f�,>v��;ovP���]�sc�=z�R�XO>(�H��p�'�4>�ζ=�8>���=q������1�}=����M�>��?�T�>t!�>�-��� �~���&�=IY>�S>љ>�1پ\e������g�V�x>�N�?�P�?�g=���=��=�1���-��������<ј?�/#?IT?��?��=?�7#?e->%��5���P��ĳ����?u�?{��>t�����v������rn?���>�<L�!sy�/�-��̶�ڌ ��+�=�u���q�!@��"�<���l�Y�ء8���?�3�?��%=��4����ȷ��)��XZ? R�>��>K��>V�4��y��x�?k>�2 ?DrK?���>�,N?0x?�"\?��5>:�H�����#��_4�@�>�EJ?k^|?�Y�?o�?�<�>��E>������1�����t˽$g����=OuW>R�w>���>ٗ>��<��½ha
�< M��M�=�o�>���>a'�>h�>;J7>&�'���G?L]�>�����M��j��󱅾J�L�.�s?��?,,?�l=�*�jC�"���
�>c��?��?�@)?�S����=)��C����p��-�>�K�>�D�>⒫=t8E=��	>���>��>���&���8���r���?G?�]�=r:ſ�Fp���s����'�s<Vɐ���d�<���DXY�z�=@��������(�_���������q��c����Vv�.��>��=]\�=o��=��<�[żpB�<��M=~ �<i# =��v���><��>�8��]'�� p4�0�B<�}O=i��{�ʾ��}?��H?�+?�VC?O`w>�">�>7� ��>�4|��R?�vT>K]P�����uC?�����e(��0Eؾ�%־"�b�e����>%�S���>f|3>)�=6��<���=J�k=���=f� �� =/�=᮸=33�=���=u�>>�6w?X���
����4Q��Z罢�:?�8�>j{�=��ƾo@?��>>�2������wb��-?���?�T�?=�?@ti��d�>R��~㎽�q�=P����=2>}��=�2�Q��>��J>���K��:����4�?��@��??�ዿТϿ,a/>�P>K>"�O�Ѷ2���^���W�8���?�8��ž��s>Py>ݤ�KMɾ�t=�;>rN�<����|jQ���=���#=48=�m�>!nH>�^�=�q�����=�$�<���=�o>�t�G�/��7:W�(<R�=�q>ת>
�>�?O6?��h?M4?�c�l����r�є�>X���N?�d>&�o>�?2\Q?Aup?��r?��>B7�߸�>��>[�8����!L9�C�y�j@��o?�5�?���>�=ӻ;Z9�	�ž	�:����~�'?�,8?��>�l�>1���9�s}"�7�,�;��"�S�B=��b��<���<����w2����>��>H��>�F�>�{>�;>�bI>v��>l >�R�<C �=FA<C��<����'P~="�
��[(<��μ�{�:�(;�T}�*2���7�;˖��n1һ��(<��=Ӥ�>���=L�>�f�=*��X>_��!F:���>3ʗ��
1� �n��Y���r*�L�k�ӷ>|)0>>)��'���! ?��j>jeD>�y�?��j?<�>=��M)Ͼ����}s����+.=����=�yf��2<�^�V��rA��0ʾ̛�>���>`j>��=�H#�X�2�]=H���5�kV?_T��>t��!�r����$��L]�
T�3W?�(��UĒ=Dq?�>X?�5�?o�>h�&� �
��>`x���><�#��3 �K��H?��(?b�>][��g�PC̾����ط><AI��O�����ڬ0�a�˷����>������о�&3��f��~�����B�%Qr���>��O?��?�/b�'V��kTO�O��&&��=q?�{g??�>qI???}���n�Lq�����=��n?���?O;�?d>�TH�Q`��ˤ?�>�>7�?ҁ�?�lz?s"2=eb�>��\��U�>?n#���5>ꔰ>�K�>��>�[?J�8?k��>b���i���뾃�����XT�=p~(>>���=i�U>3*0>S�Y>��=��>�iG>ӵ�=�y�=���>�\k>/z�vik��)o?.?����j �>���>�T<+ؾ�s�:��W=H�̾�bA��z�>����jb>���=��=�����t>�ʿ�?��=��Ƚ�>?�]��"5���g�X|�>�I˽��?�qA>��>U��>Q�?��==_�>;ks;G��I�>�z%�Uf3�pcB��6+��A۾o��$f�[^0>,�����6U�A���6��Am��&��`10���->�N�?��u]i�*�T�f|G�>�*?�+�>��,?覕�M�I���V�>�Q�>��5��ㆿ�蟿x���Q�?� �?VDc>8.�>�2X?�?�92�M5��Z���t�|aA�D`d��_��č�g���=�	���ý�y_?K�x?�rA?	��<�?z>r�?;�&����%ȋ>�=/��d;��H=��>Kݱ�\��<Ҿ��þ�&��<F>�n?���?�?�)S���p�c�%>�:?�b1?Gt?�;2?��;?!L���$?��2>�0?�2?\H5?l/?��
?��2>\�=ﳊ�&('=[���m늾/�ҽBOʽ����0=�6y=��K�<�=��<�*�;nټ�;�ូdn�<3X9=l��=��=��>�gF?Е�>\}�>lp?�꽢!G�^�$�E?�䒽rj	�A	��]߽�۱�
�o>���?OK�?#FH?q'�=����w(��$>��4>�W�=�*�>8J�>¾P=�����"@,=x�=��?�)K�$Z����#�9���:B>��>�4�>���> �7���O=-6ɾ�8J�;�_>�D�wM�����9F�v�/���^�"؞>�F?�O?27<Ļ��$���f��q?��;?�nc?9:�?n1<�s�B�i���G��D}=��>�������'���0��456�K�=�>+�ؓ���>6��q�+�p�x;�g���zûO� �z⻼����K¾}&��L<Fy�=� ־�p(���������}J?�:_=������X��%��K�>dˌ>�)�>����M�W�0?��Q9�=*�>��*>�}.:,����`Q�G� �?g�>NB??q?ʻ�?�ƽ�鐿=�v�N�׾�}t� ���"?���>Rl�>�3#>Y��=C~;�A����a��P�9�>�?�A��Cn� ����	�q@g����>q]Y?r��=S��>u�??'K?	cO?͎2?�V(?67e>��I�TϮ�b�?�?�>�_���d���C�8oW���>�Y*?~���>v�?h8?��)?{�W?�!?țI> ��<O���>��>�R�)����D|>��D?��>��>?b�?�,K>Q�.�����0���@�=/L:>��7?Ua#?y�?P�>��>�' ��4�>��2>jxM?�6�?G�?u�,��:�>�?a\�>���['�>84(?���>z{B?�G�?LI?F8>��=%(��8��tC��c�FL�<�TG�shҽ a6�#e�=�۽��p��ft>#>Th
�r<	�K;�Iz*=Q�?x.�>��?��'>X���,g����>P�=��ݾ�μ��I�m>r�ѽ❚>���>Z������'��>���>��
�� ?��?��W?`s�����D)� {
�r?�>,V?��=�of��Y��|���7����?a�W?�J���5�
�b?e�]?�9�2�<�9�þ&%c�%����O?��
?οG���>��~?��q?���>��e��n����YIb��k��׶=�q�>[�a�d����>b�7?<*�>0�b>��=[۾r�w�����d%?�?��?���?�*>8�n��'���������]?zt�>�V��F�"?�����Ͼ�D��E�����ᾟ���{��)P���^����$�����)&׽�>�=ȶ?Cs?�Kq?7�_?� ��d�M^����f�U�j�����ϪE���D�q�C���n�Z�� 1���똾=,E=3]@�� K�팻?�B?�MC�.?�> )o�^�JS�7��>aGl�T׉>5K�<���=�H>0�T���>�$����|	?zR�>�c�>XxK?�����3���1���A�ޑ���.>�L�>G>���>EP��6���7�*x�%�s�3��[�x>��d?�L?��o?>Ž�8��J���G��%���۠�(�D>c��=�8�>�5�����K�>�9�F�v��|�4)���d��g=ر1?�>�f�>�?�K�>Ow��ܫ�V��ʿ8�pG�<
��>�l?�F�>0"�>������$����>&!a?4��=�.i=��̾M����`T�
/���Q?���>��>�-�>x�P��$#��"��΂C�`��;��a?s���&�Y�j>KP?�%�����=�b�>������$�ϳ�Q9�I��<>=1>_U��?��I��}��(?�?�U���G*�̯~><�"?d�>��>���?SН>�pľ�$����?�B_?�;I?ȌA?77�>,l%=^�����ǽ�T&�*=�̆>�YY>��h=�]�=���[�u��W�:=�z�=��ͼß��ah<u��X�o<[��<$�4>�Lٿ��J�������3��a��䎾Y�z=,^~��͝�ἴ��`ݾ�b������;)go�瞊��PP�%�h�J��?K� @%s���D�"�����ܛ)��A�>Ƚ$�����/���#�<`p��� � 齂; �T�D�j�V�3�s�w(?��ʿ�d���'��.?e�	?�?����?��Mo�*�>D�D���vi����@�ſ3`���>?0��>��Ծ*��=_S�>t(�>�ت>��=����<��]S�c+?�0Q?D�>��Ҿ�ſ�����e>�#�?�=@�zA?��(�1��l�T=-��>��	?b@>01�z9��а�})�>13�?pފ?��L=�W����Qe?�<	�F�q?ڻռ�=�+�=S�=8��<rJ>F�>���4tA�RXܽ�\4>�ԅ>��!�Ƞ���]��\�<�c]>U�ս2��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�󉤻{���&V�}��=[��>c�>,������O��I��U��=֕
��Wؿm%&��L�w�/;�`�����ޘ��.��`�9���_F����=0��=��j<�Y>�xE>��">��>>tK?�+T??��>�r4>��Ͻ#��ؗʾ����Uʦ���H�J�-�@�L�ฟ�#I׾B�q��
��D����E׾��9��.#>�NW�qVn�[o$���z�\�X��N?��6>�%�hvY�5Tb=dD��f��V�=D���Jݾ�o[��R��o�?6V?������4�H/��x�@�����R?eD=�>�) ���=^물�B�=��>��>�#���x��\���6?�?����J�{�"m�=ޘN�!J�=�2?�z�>�gk=���>�4?�o��8�ȁ>�~a=��g>�l�>CA>��z�nҽ�?Ig?.�����ݸ�>?�%��¾`�<~c�>}U��9�+���y>��l>,Pj�84�<sC�c%"�/�I?}k�>�j�1��������=��>�=*?�n?���>+�S?v�;?F�
���WbW�9&�ʁv��R?�Om?��U>L*
���ܾE����?��@?���>�}=�)���H����A�>�]?{ON?t�L��j�q��8���DB?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?p�;<��T��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������u>�䗾V��? D�?~������}��][���G��q�=�2G>�+�4�=M柾r
���p�K���LW��4���T>��@r�i�^U�>���=�V�"տy���H�
��.����?=��>��¾����jd��v��c���=�*վ� �>�>����.���sZ{���9�g���P�>�����%�>{qV�����E��7��;���>�j�>�;�>p��7��av�?o����Ϳe���gn�-�W?q �??�?{�?P��;��u�z�v��� � �G?�]t? X?�#�8�]��/�59O?O��|�r,D���B�UG�>���>�'�>��x��l6�zk� y(?(8�=��T�Bs���,�����1n?A��?4 �	�?�҉?�\<?hE��/���ξ!�e�!�$>`�o?�?=Dž����i%��{%���!?��?�qн$��]�_?+�a�M�p���-���ƽ�ۡ>�0��e\�'N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>hH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�8�>�΃?�V�=���>���=!}��+n¼�4 >y�>T�-��2?�ZO?8��>o��=�sL���.���F��oP��d�	sB�>r�>�f?�@K?Sic>��Ž$�3�?�#�D���7��B�:@b=��Tg�[���+<>�:C>�� >�1@�g�پV�?cm�9�ؿ�i��9v'��64?ǹ�>T�?���4�t�Ǿ��;_?v�>�7�i,��z&���J�f��?_G�?��?��׾�%̼S>B�>�C�>��ԽF������i�7>��B?O�C��j�o��>.��?u�@%Ԯ?�i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?pQo���i�B>��?"������L��f?�
@u@a�^?*��V��zD��0�ܾ��<� �=��W>MX<�e�>�=[��A^Q�e�w>�:�>׆=�f�>�d>	aH>|45>�}���(*��崿�W����2��m��?�p�F�E4�j�����ξ�6d���D��Џ�Ĺ	�����۫U�ns��q*�=3DK?�FX?z�?/HJ?sC_����u�=�+��H�>�)�>�	(?�~`?�c?v�>�=��X�&���Ȿ���
��>��x>\f�>g.�>���>�#=>l5=��)<�j�>�4�>~��}��.9=��=\��>�?S�>C�)>�6�>tӲ�aߒ�\%o��۾�z��|�?(�A+{��$��Z�M�R8�=;�=MHN?D�K>Fr���ٿ�c��yS?���p�4�Ω���[�hf?�5�?d�g>���T��=8N�=�U�r ����9>в��.���f�#�}�?�*?Fg>)u>��3�r8���P����&|>%�5?�ζ�FY9�*�u���H�|ݾ} L>X1�>qO��z����3�~�;%i�Nyz=�i:?/^?0�������u�
͝��jR>�\>�y=n �=`N>�&f���ƽ��G���-=�Z�=�_>Q�?9�>�n�=�>Uõ�����޴N>��ؽ���=N8q?�?�6�/E��TѾ6��n��=Q1�>L�>ZA�=I;\�y��=��?�>�ȕ�'�=j)X�z-�%q%> ë=��0�C����n>V��Q��<�=�M,����>=�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>�=�ᕒ�$���<�t�ŭ[>�a�>)�
?z>ݾ���`�R��b�>��x>ԕ�S����6ʿw=l��\�>8�?m�?K4i�����)�� ?��?&C?I�?=K���������0?�e?P3�>����+�J�?�ɇ?�sy?�^>\k�?x�`?��>�qн'��吨�Ǟ��D8>0-�=�`�>6�2>'�����P����p���% _�|t��dO>�y=�̸>�P�l��m�@=� ��\��|�k�UԺ>1�>~:>�p}>KD?�5�>ln�>X` =�"轤����f���K?���?j��Rm����<:i�=�a���?A{4?�a��Ͼ���>̹\?x�?�U[?G�>^��S������En��[�<K>���>��> ���τL>�)վd�E��d�>��>����eھKj��Ɓn���>�]!?L�>���=\�?��%?�q2>�	�>[wB�nmr�j;.���v>�g�>?�og?4�?c�ݾ�B��c�������mW�n�X>r�r?C�?.�d>�p������9�G�f_r�={��?�M8?~Cn�i��>�'w?�x5?MgQ?� y>�ʁ�A�ɾ��K���>�!?���]�A��Q&�>0�K�?9V?���>����uսVJԼ�������?D\?W&?5��3a�|�¾g��<�/"���T�k\<<G��>(N>r!���I�=��>�د=S�m�h6��]<r�=�`�>���=+J7�mՎ�ov+?@pP�����2�=v�p�eaC�-ˀ>YK>7¾��]?�;���z�����f���5�Q���?"��?���?~ҵ�LLh��u;?�Ӈ? ?�m�>/�����پ}޾v�t��7r������>7�>i�r����^q��lE��ę���P˽�0��>�h�>��?9X�>DsD>�s�>�
��[ #���;/<��2Y�����;�Tv/�/��vڠ��&�� ��Ⴛ�s��N-�>����Pv�>�?|�r>Ï�>�>�P��#%v> T>�8�>J?�>�`>��>��=�g^<i|���OR?����j�#�n?�H^��s�@?��f?�0�>.=��#���D��? ?l��?7֛?|rr>��j�%>*��6
?��?/��Xp?".=Z�?<�-��o���#�����(&�&��>7�	���<���L�m����?�?"�M�O�ξ�� �(J���p=>=�?6�(?��)�Y�Q�ȥo�;�W���R�����h����o�$��p��ݏ��O������(��)=Oi*?-�?�m��x�d���k��(?�:�e>)E�> �>lѾ>��I>"�	��1��^�'�ʃ�gC�>@%{?�x�>voH?�>?�V?Ҭ[?ϯw>c�>b��sG�>Y��>:��>)3?�s.?�w:?�"?��1?��t>7j;� ���Pkھ/p?B?@O?��?�?Z�u�f��J�� �;ab�c"��9�<|��<����ռ^e�=�~g>f�7?��̽�)�� :�m����V?	_-?e�B?�t��Bl���=:�8?V5�>w�>�@C�[�8L�{��>��?ԥ)�T=N��>���=��=4J���	=9�=hJ�=7�<����>��=����5.>(��>N��=��?����=�Lc���>�/ ?L��>���>�0�������j�~c=C�f>Kg>eE>n�о����B���	�f�3�p>4�? r�?`j=f�=���=V���$~���t����4=�%?T� ?u�P?�H�?��9?�$?GL�=��f��l���8���5?�-?q�>L�
�Xq���g��i|6�Gs?&g?��b���ӽ�g!�Ož�oȽ���=�6,��bx��T��cCA�"k<�o�������?���?+tG���:��H�6������2�K?��>'6�>l�?V#&���m����N	R>���>��K?���>3Y?R\z?ǿ�?u�(?�c��ÿ��l���^>����63?)?��?BD�?ZU7?#�>�лK�!��	O���$����M����=AC�>qd�>��>�H>l`�<�t2��h��q�2��?$=�0�>�[�>O��>��	?�h�>m	���G?���>(@�����lҤ�����ii=�Cu?|��?�+?�n=Lv���E�I���G�>�j�?H��?O9*?��S����=�w׼�ᶾ�q���>^�>�7�>O�=Q6F=bX>���>ٌ�>��I]��c8��9M�{�?�F?�=9
ƿ��q�t q�'Η�LQ^<j��d�S�����Z���=Z��������G�[�����k���������Y{�/��>���=-��= �=�+�<4�ɼX4�<�\J=�g�<7�={oo���t<r:���ٻ����t��	^<`I=��ʾ�y}?��H?<-+?�C?)�y>}Z>JA��A�>��{��*?�V>Ϩ[��{����<�����%F���ؾ��־#�c��x���>'�H�|.>(�4>���=4E�<��=Y)x=��=5%y���=���=���=��=�%�=�k>�>>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>A�7>wy>g�R�f�1�� ]��a��{Z��6!?x;�2 ̾���>먻=�߾�Ǿ�*=��5>�E_=p��� \�P�==A{��==NFk=��>ED>cS�=�䮽~�=$�I=)!�=c�O>�J��/J:��+�cq3=�y�=��b>`&>�#�>Y�%?&tF?}{n?M7'?|q����	�ҙɾ˝�>����u��>j�8>��v>�o�>T�U?�^?:�b?�;�>>�p�/��>#`�>u���"����ܾ��:���=$�L?1�n?J_�>���c�\�w �m�8�'�7�q
?�aV?u�4?�>������������((W��ὕ��=QJR���� Ʊ<��)�����U>��>�%�>��>��=-��<@>�}�>Ba6>�T>0�P>���Y�x=y��=��=�Ԍ=�FH=\��<Q4�=�\��ƼM��=����j�=��=�Y>=��=���>�>>�o�>OQ�=󄷾=N.>&����N����=}D���qC��*b�G>}���.���4���B>��R>�'��w瑿W� ?We>O8>YB�?9�u?��!>g�
���վe����d�I^Q��f�==B>��;���:�Y�_�MfL�@zҾ�h�>}5�>T[\>2>/�$�U_#�`<�������h�>]�~���<�ff��t�����g����f�ieK�s�D?т�t��=��?OB?e�?�ܤ>f@ٽI+�{�?>1棽�5>��@���1���?��/?�f�>%�̾�rV��:̾l��Ƿ>STI�2�O�����ڪ0�G��ķ�]��>����T�оa)3�Pi������b�B�cr�N�>ҵO?}�?,Eb�qV��RO�t�����o?ig?0�>+A?~/?���tb�m���k�=��n?ѭ�?6�?�>�4=�&��?L0�>�k�?<;�?�|v?]-���>��=�b�=���C�=s�>>}��=lw�>k_7?�Z?��>Lj� ��������R��[>��F>;�>�}�>l߰>��<����!>� A>�{&>��>��-<��^>	ގ>͜#���dS?B�>TT�=�D�>��>U�Q>ab�Cˁ>��}=f̾�hv>�X<Ŝc�l]=D�<�vȼK���1��>_ȿr}�?�M>��ž� G?�q��.=�<w>Ў��i�ؿ�>��>,l�>�Q?�m�>��v=�>!�=|���:� >H}���)�fdI�4��Ǿ|�9>��7���� ٽ;2q�#�޾Ġ�C$p�J����A�\ۜ=���?�=��^�z�)�z�`���?�b�>��@?*́�?����4<���>�ٴ>
��k��|����$׾�?&��?~Lc>�'�>��W?��?�m1��'3��jZ���u��A���d�Ъ`��Ѝ�����\�
�oܿ�H�_?��x?~qA?
�<1z>���?��%�_Ǐ�#�>8"/�,;��0;=M�>� ��	�`���Ӿ��þ	��w�E>��o?d�?V?�/V�M都
 >�:?� +?su?_U:?m[A?�0��J ?��>>�J?|�?�6?�.?}�?"�:>D�>Qx�<	=�</�������t�^���/�[=��=?�ֻL�
=M#D=:�<��ݼغ0��:m<d@��+�<_O=!�=j��=zGy>�j:?S"?0ү>�y?a���������N� ?hp<�boy<쟾樻�������>��?�R�?���?x��< �b�S�žX�=��>!9g���>e?�v\=�ӗ�R�">G�p���=���QN���U1
�r�I���
��B�>y�>�~}>|Nv��k;>*a��\�����b>G�H���þ��6�̔B�M3�np�W%�>~I??:2�=ů�ط���d�ٞ'?�R=?j�N?w�|?�I=��߾�;�y�K�^k���֠>7��:F��1����?��U
4��t�;�d>�?��F� ��$�>���Y�ݾ�{J��	X���>���а����=!4�ȼ��3�M$>
t>O,��ka�0��q��E�N?�V�=M����UԾG��+7>���>�{w=��(���<���%������>�O>��K�*��8du�����a>��=?8t?���?�j2�M̂�S1t�#���X��ZKQ���A?�p�>چ�>�}<��9��kt�~|���Z��%4� ��>�V�>���Iv0�������o3��P�>;=?�Wa>Z�>�{x?h�#?�S5?h;?�T)?�'x>l�-��B���%?���?%s�=7�ӽ��R�{8���E�34�>�)?�U:��z�>Ģ?#�?Vn%?WCO?��?Z�>js �k7?���>o�>^�X�]����]_>�KJ?�E�>�Y?˯�?0�<>w�4�y���U�����=��>H�2?[�!?�w?��>�G�> ڢ�E^�=���>�b?B��?i�o?G4�=xc?�o4>S�>��=�נ>&��>T�?YDO?b�s?�|J?��>�φ<�M��a��v�p��uY��@�:�JE<9Dp=ˎ��7o�����7�<�%�;�����R��2m��`�.������D�;�5�>b[e>���K�>�O���x��>^,�R��̧i���M�x��=L�>�y�>�N>AK����<��>�U�>�t"���3?nh?�U3?ˠQ���p�ա ����%��>]�C?{!>>�O������k����Y?��j?�kT�^��_�b?]�]?g��=�
�þ��b�~���O?��
?!�G���>"�~?��q?���>��e�6n�	���=b�Y�j��Ѷ=�l�>�Q�:�d��;�>y�7?JP�>)�b>��=i۾1�w�Hq���?��?� �?���?]"*>��n�v2�̔����t�d?��>�ޫ�"�?\�<q�Ⱦ�!��
���X�о����HΕ������O���}�Tlr�����I�=[�?��p?@wl?x]?B ��d�8]��q���wV�5�
�c���F�kDE�2@�pr��M���-U����	=��|���X����?;8?��_����>i
��˾o �&An>�+D�
	K��uO>�lp=�4W=���=,#���ؽ�����T?y-�>���>�7?��K�VU?��*� �6�l��;.�=G �>��T>��>�Z:<�~�� :�C��xޠ����Li>Pxe?�}O?�]r?�O��	P8������$�촥�r'���P>��>�ơ>�5L�Jm��*���2�1gu�-��������6� =�
-?���>�W�>N��?� ?�v��1���^{���:��O���>�i?z��>BɎ>}Ƚa��m�>~�j?�l�>���>%�}����m�|���&���>j��>���>0�>^�q�^����>K����'��)�=�a?�a��v�4�#+�>��L?5��;�<�$�>?������.�ξ��ݽ%D">�� ?q#�=�)>{�¾�Sھ��l�x׉��f.?t�?�W����0���k>�h?�i�>Ι�>��g?C��>�.���E<�@%?�g?G�E?kw1?��>>�5<*{.��� J��j�=g;�>գF>��G�^��=匾G���D�	 ��n�=^�H=�ӽ���<�h��a@�=��<�=C��I�^��^�`��6�ɾ��Ac���k��k������þ�d��s�}�*���ń;�����O��RZ�Ң���|�?��?cǨ��ь��<��uCh�\���o�=���fM�������4�#C�>Ӛ��+��'Y��Dc�(�^��a}��"?�^�����>e��N�۾X�3?z#?��x?+h���E�kV�B�>�x�Z����X��jÎ���ÿ���H�J?�ۨ>;9��WHʼ���>(0>�- >M�>M����E��;��?%�A?&u�>"[��y¿�|ȿ���<=�?�@�A?�R(�a��jC=��>3�
?��B>v�*�҅�_��m�>���?		�?��@=�}W�A��3c?|�T<d�C���"��H�=���=�<�����N>Dw�>i�UAL�����/>g�~>�3����b'T��<�<X�Q>GsȽ�p��.Մ?�z\�/f�B�/��T���S>��T?P+�>e6�=��,?�6H�B}Ͽ�\��*a?�0�?���?��(?�ڿ��ؚ>��ܾA�M?�D6?3��>
e&���t����=�7��ڤ���㾔&V����=���>S�>��,����O��<��V��=�	�r@п�� ����x]$=O7ü�\�����1 ����,��O����V�X�׽Ge�;=3�=,^d>ԩ�>��_>�B>zCg?5�u?@�>�_�=�ýq���Z��jc�©O�v��M����.��\��1���2/���F�)�U���YȾ�!U���M>*�Q�e������&��jWg��v?��>�=ľ�|�L�f�q]��u�;��d�=\!�s����Ui��녿�ئ?��"?������-�9�3���޽�=W�n?�hҽ�?)�c���;R>��#�MF��b�>���=�����PP��:9��6?tZ?b���h��L�N=��E[>� ?Nߤ>��>�ر>��>��/�|=d�"'�>F:�=��>��>U?�=�w���Ⱦ��8?�l?V��-5Ծk�>��2�rվw�>�b�>b�$���<�9>=��>�{�xX��V�=u�=;�B?ᥭ>m6�d9�*Ɂ���=TҼV�??�.#??�>�ZP?�G?�ͨ=Y+���q�q_�M%�;q�I?f�?%�m>j⓾U�^�����?d�a?qJ�>��=��0���Q�F$��J�>F�Q?oJ?�C�=K�f��M��������7?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?r�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������ă�=#���b��?�v�?v�þW��/�ݾB�d�*B��u��$Ĥ>D�}�"�u� ��z5��ԟ��C׾�ŗ�����R\>pS
@�����|�>��<»ӿ�������
d�������,?t0�>�᛾�{��Qp�(�Z�Y@?�I�J�����Zk�>� >
����o���ez�|�9������n�>d ��!�>;�U��Ŵ�l��_��;r��>�K�>z|�>h���.���YI�?M���RCͿ�S��v �v�X?[�?a�?��?�'�J�w�J��������F?W�r?u�W?��6���W���2���Q?"����f��9H����_��>��?T�?Ih߾6:�u�<��(�>��/>$U�O��"4��������?]k�?h�'�/?l }?�e?������{����X�d[>�!<?G�G>󧽾y|�F�`�|
þ�f?l�?�+e�����_?h�a���p��-��ƽ�ݡ>�0��^\��9�����We�����Dy����?�]�?��?���;#�35%?d�>�����8Ǿ���<h��>�'�>X-N>�5_��u>5�H�:�ol	>#��?l}�?|j?��������.]>3�}?�>��?JO�=�"�>�O�=�����:��-">���=��:��|?ђM?�>n��=:��/�	F��R�o��!�C��m�>0b?��L?�b>9g���O6�u.!��M̽�-0�+߼�Y?�X?-���߽!|3>�=>�@>O�D�BNӾ?^���LؿNh��Y(�65?���>*�?x��z�c�5�M`?�ȇ>����*���~��`����?�G�?B�?��ؾ�@ּ��> 3�>� �>?�ӽ7B���U���w8>�aA?ޚ�����5n�ȅ�>��?1@��?:�i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?jQo���i�B>��?"������L��f?�
@u@a�^?*�ۿt���O���p��¿�=��=2k>����IS�=��<,y��_<\��=��>��X>�u>��f>�#b>uH4>�����%��8��H��u�J�v���t��K������8���ґ��5þ|0)����Ik���{���t�$2K��k,=�qK?x�`?"*�?�b,?���=i�=���(s���:�KD'>ތ>�%?"68?FK??0�6>#��[��0p�����w7���w�>r(>�s�>ȋ�>F��>^��;��>F >���>��a>�5 ��钽�O
>��$>'��>F�>�0�>�i'>7�=�p���7���y���[�!�?]Џ=K\e��4���"� �S?�*?_k�>�͓�H�ݿ�~��d8P?�b ����1�A� >$�}?	W_?�>-n��v'�����>�`3=������>i��Pw�'Z����>IR2?�yj>10u> �2�5U8���O��®�M�}>`6?���c�5���t��GH��ܾ��P>T2�>��L�e$��@����}���i�6�=�9?�?�(���n��(�s�/i��|�Q>3�`>��=��=@�P>/�[�n�����C�h�7=���=�\>"� ?O�>�G�=��F>�s��
}���>��ɻx�=ve?˄?{�ʽa)��&�3���3�o>c6�>$�
>���<��XwJ=��>�=����Tl�<��޼��}:N>�#����������1�W��R =���=�,`��-^���=�~?���)䈿��>e���lD?V+?	�=��F<��"�@ ���H��2�?q�@m�?��	��V�1�?�@�?�
����=�|�>�֫>oξ(�L��?��Ž>Ǣ�	�:)#�hS�?��?C�/�Qʋ�Ql�p6>	_%?ڰӾ���>O���3�~��s���>���>�L?{��}X��F���/�=?��>b'������ҿ�#h��&?�?D(�?I���o p�˜M��
?�,�?pQ?�)�>۟6�Z�ľ�N'�TYI?��A?��?����<#M��?��?�??\;>��?*M?���>V����"��J��Tƍ�µ�=��/>�J�>Mz>��B��7���܃��-��y�P\o>�"=j��>74�jQ���m�=��x:�n��\��1�>���>��z>M�>Y��>���>0�>cr=�=�X��Ȅ��][L?�z�?���m�׸�<��=��C���?E�.?:�4=�I׾�Ԧ>wd`?���?��Y?�-�>|D�k�����S̷��,�<��V>ڎ�>-p�>���l�<>��߾_.��;�>+��>�C�5Hʾ��~�S�l�`�>� ?ђ�>��Q=V=?��%?o�]>	�>��A��ď��XF��m�>c��>�6?�b~?��?��C4�nb��&����U��F>�(w?�?ȏ>�=������I �l�!��瀽iV�?ie?��V�?��?�<?��<?��l>�1
��߾^���ϊ�>�j0?}��/��)+����?�?kB?L��#[�����g�� ��?�iF?�P?<�ݾ��=�+ϫ�"P���e�=��m=J�ӻ�M��C�=kY>ϱ�����=�s�>B�{=!�����Xx�=+�>�ռ>�Y>r�+ؽ=,?��G��ك�t�=��r�*yD�+�>�KL>�����^?9e=��{�����w��=U����?���?�j�?p���h�_#=?��??t�>�L��<z޾є�4Uw�Tyx�Mw�~�><��>�l�`従���ǘ��DE���ƽz,ν�U�>+l�>!z?,�>�C�=�p�>�Ƌ���5�G�������m����/�:��W	��Տ�~p׽�S�����Q�X�>�̽��>(;+?%�O>㌕>�Q�>���"�w>��<>	M�>�,�>Ss>3~>���=y;	�������T?�H*�Q�1�P�h��V�q?@�H?Y*)?{)G�X���D�R�/?�!g?�{?iO������x1��T??�-?��,��R�>�D�<IvU��*>�˕����B:�<9x#�he�>xb�4�g��k+��M���?(�?īS���վѰ���,��p��=:��?Xx1? $���U���u��P[���W��Q��"
�c���3�%���m�����? ~���|�x�%�冤<P�#?��?���/#ᾥ܁��'l�dRV�`7P>��?{�>(�>큓>���q�>�9�V�l��`�x�բ�>}5{?�[>_I?�C@?3�L?�Ud?�- > �=>��پT
�>K��=��v>�V�> n6?��)?%7?��(?�H??费=��x�FH�;vɾbk?\]?s�?1��>���> ������i�S�ǰ�x��n���2�h =Ir4�&�</�>�c~>�$6?�㜾�c+��9��xP>��G?���>�S?7��}+��3�J��N>�Ub>�x�>nϾ�pk�����>�U?��Ӽn�j=�6e>��=�e~���<bd=˕=ZqQ=��A=��%=$���'A�(Q>��=��=z�=Iz׽�(½<��>�?e1{>:'�> ������a�䣩=�u> �0>n�>��ξQ��F_��Y�i�A�a>�)�?�Ʋ?�L�=x��=f�>���r��ʸ	�����1�<8D ?z�%?:SS?�?�s8?�V"?Bh�=�v�l)��'����|��M�?�`.?a��>1*ھJa�hڦ��]S��/.?h?�e��w} <1q˾!��~rƽ�>e�Ծ��i�B�����kx�=�J�ӽ�N�?�F�?Gv��J�R�z���������75D?g��>L�2>�i?-q��Kh�����[>�@?B>?U��>nZ?��?�(r?q�>[�ظ�K����=�R>��D?3�?Ay�?��7?-Y�>���>����pT��!��+s�Ɔ����,���:�>�>��>	
�>��=��_!n��坾(T/>~�>G ?�'�>6X�>h��=:[ս��G?iW�>�⾾��򤾑���9���t?�X�?5�+?_�=�j�F��%��?�>s�?��?��)?��S���=�d޼
�����p�5n�>B��>�E�>�z�=�D=�<>�(�>t��>������7��%Q� �?ƸE?���=��οc"R�Z1���:���֣<�d�����	�*���%���=�����@�(�BxP��Y��T�t�6+���ː�mV�����>:>P�J>^2>�W=�X����лS�8�D2*=�l�=�[�y�<�J=p>�F���&�<'������齗�Ǿz�}?5OH?0�)?��A?H,r>
�>\o��>m�E�9�?�KV>Ӂu��ټ��h9�襾�����ؾ&׾�B^�>5����=��Z��
>�03>K��=7�<���=.�R=Ҏ�=j+f���=}|�=,�=f�=?�=�><�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��F>� >��O�Ԇ1���Y�@�W���M�e"?��9���Ǿ���>�@�=��㾇^��_=*=�8,>�JZ=|��g�X����=mJ\�y�A=�Jn=�I�>�<>i�=�l��mų=g]]=���=V�L>�R�;qF�����X=���=��U>�`&>�t�>Px?��<?�wm?^�	?f�N�ɾ[���8�>v=�=�"�>z>�+(>U��>��J?I`?V(`?C�>��]<���>��>�W*�2�u��ɍ��-���L"��x?��?_W�>Nȅ�0x�<}��:����-?�4?��?�F�>"V��	U&��.��m���Z�H�)=��r���T��2������㽖��=�i�>���>��>H.y>]�9>4mN>x�>h�>���<K݅=z��܇�<����O~�=���� ��<@/ż(��J>��r*����x�;IL�;�
Z<%��;���={5�>��>a��>�3�=�ض���8>�����N���=����M�C�LLb��L|�7�-��'7��B>�[>�������:^?�d>��;>���?��v?�!>���FaҾE����j��T���=��	>l�=�� 9�'z_��bM�5�ҾZi�>s��>���>Ol�> *��FF���=�:ؾ�C?�@�>�sp� ����ֽuTc�L���!���#[��=']:?'s���!�=b��?HG?�V�?|��>{(����޾�.H>|`i��ˢ<�����a��Z��	 ?�q!?�?��j�E��:̾�㾽Rٷ>uEI���O�����0�0�!i��ķ�T��>������о.%3� f��������B�6Fr���>ίO?��?T;b�W��6MO�a��n���n?�g?�>3@?2B?5��:l��k��Jk�=g�n?���?m8�?V>�=A�����>G�?Gp�?z��?��Z?)��.�>@�&=��+>'hO����=���={=>(��>P6?W�?gJ�>W\���w�d���!��h�s��"F=A��=�}>�_�>���>�Kd<!��w="�w>[�>�j\>X[�>f0�>ȭ�>���]��ޙF?��>�9�=��?���>E��=����H��=��=�P���~3=��h=N��<���=��"�M�	>����휚>g���@��?�K>��ƾ�i?iX��񮁼��X>'�>)�8=���>�a>��>���>e�>��C>��G>�)>l�Ⱦ�>���. ���F�CaE��ξ�in>�z��0N�yA�K ɽ�Y�6�˾ҋ��Ti��u���?0�^=
0�?\�½v�g�/"�2���?e�>M-?}%l�'^A�w�5>1��>��>no��o������{�a��?��?2Pc>n*�>�W?"�?��1�W&3��fZ�+�u�GA���d�L�`��܍�\���,�
��@��7�_?G�x?BfA?a��<�Fz>O��?��%��̏���>�/��;�Wh==�%�>�Q����`��Ӿl�þ:,��F>+�o?, �?(P?�"V��;�d@>��I?��N?��?XU?�c'?X�r��? �=��?oT?+I?ѻ?)?�ރ>�a>b�f�������� w�'^�_A��Z���2}=�d=�<����=��a=��=��=g"<�$�2購ϋ>���=(ip=�F�=j\>�H?7t?�}�>A��?��o�7'�TL��/*?F�>��\���"���h�H��[|�>˲�?+�?�Y?�)5>�ng��pU����=��=Vp=�7>k��>uZ��"�Y�&�=Ԅ<���cU��6��T}��l���i��tv>��l>B��>r!�>��Z�s�#>'���oo��g�e>�t[�C��ƪ���E�>/��TS���>;EG?�!?�o�=��ྟ���*c��$?��??[K?n�p?HuI=��־��=���F����A�>t��;�2��F��!4���7����q�\>�
���~��1l�>�� ����S���N�h���]ƽ�����=��<r��e�۽k��=�d>1n���$&��L��u�YU?!�G>(쾇Â�t��~��=#��=m��>x�=~zN���<�?����i���>O��>~.̼
)��^�Z����%�>ag??�v??Ж?�<�H�]��s�^�����;��.?���>R?��>�@
>hkx�'T���4C��AU�$3�>��
?��D�<���:����H���S�>��>����[�>R5F?h��>�{?�I?e��>[K3>���1 ���s#?��?#��=Nh)=C����C��!R����>Fg?�);�䉵>*�?� ?��8?f�_?> ?jy->A���ۭI��=�>Q�>��b�P���:˦>C�O?�J�>	B?y�n?gNY>i+�>����6}��e]=v08>�=?95*?a�>�V�>��>�˾s#�>�x�>@�Y?!#x?w5�?Yԍ<DE�>3�l>���>��:��V�>�? �#?AdM?k&�?�h?��>����A������X���=�54>2h>�\
>��<��� �(=	:>([<���*8>�F���iD�HƲ<2r>�0�>b��>�����>?��~﴾�p�>T輎"徂[N��O�>�e>�9�<�g�>O�>M^����=���>��>Q�#���?w ?��;?޷>Uh��I��W��.��<!CE?�V�=��������P+�1>�w? D?�5;ӎE��b?��]?]h�*=�s�þS�b�f�龑�O?��
?^�G�>�>��~?>�q?��>��e�):n�����Cb�e�j�UӶ=vr�>X�l�d��?�>�7?�N�>��b>A�=u۾��w��q��z?��?��?]��?)*>�n��3������H��t�]?Ik�>05����"?PZ���ϾZ������"�_ ������=5�������u$��܃�X�׽���=��?11s?\Xq?��_?�� ���c�@%^����3pV�.���ԾE�w)E���C�D�n��]�4b��j5���ZG=M10�x�8���?_�B?!0��0�>H�����ھ�������> ���/�����:>��=��<�1>��F��i�=�/��?�<�>Y��>��n?Q�j�,�R��`���_�LN���g6=q�>�1[>ƾ?i�K<�4�<��=�lžO�x������v>�Mc?2�K?�o?�6��1��:����!�D-=��ϧ��F>��
>`�>�DV�m���-&���=��r�����됾��	�,�=�2?迁>��>��?�?�	�$��P�{�:2��̀<=�>yBh?��>���>IvԽ�!�M��>�g?��>�ފ>�݃�<&���t�4�a}�>��>[�?�֙>&%u�G)b�����^"���3��>�Ud?Z�~�s&5���b>=B;?q�<��A��݌>QI��y#�w�;)�颏=n��>\ގ=/!5>�þ�w�e�
��'?l=?������*���s>�*"?Z��>A>�f�?��>	�ľ�+�;^�?�^[?hTH?	�>?`��>&W	=����-ǽ�2#��C=E��>	hU>ҟZ=��=�d�W�T�~N���-=&�=�(b��Iӽ"ig:��ʼV(�<Q�=ق2>-ؿ�DH�hپ�%�����|�������S��̾g9��F�.���MR���]�D�g�t>����n�jw�?�6�?A8���{��;���}w�y����Ǩ>���=(�����Ƚ몦����<���D�A�a�P5k�Y�Z��].?��f�k�¿�ȣ��쾨�3?�t?�7{?y�2��:�8�%�zG>��="�Z�Bϕ�\�ɿ���H�P?��>�I�b�׽h��>LJ�>��>y��>����.�?�?���>ڵD�Gʵ�8ᵿ��7��?�?;v�?�cA?�:(�^�L�X=4��>}u	?5\>>h�2�T��k��/��>��?b�?�sQ=�=W����ee?��;��F��ѻ�V�=`�=Lc=�=�fK>]c�>���e�@��ܽ �1>���>k"����_���< ^>�ѽ�G��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=��#�׿����\��A���_��!�+B�g�<�^�>u�پ:��ly�;�* >ɼ����>��>e�=��>.a?3�?���>f	>O-���%�����X��Ś!������h��[��=U�w��y������6��\�-�D�.���Ӿ�'��P>�Q��ҁ�gp���t�a��	?�g�>ce����m����˰���"M��A">�$����ޒo�ɉ[�(՛?��/?k���G:�����"���*,��Z�?�)=��/�Ա��X��uQ)�+��=�U?�������,�G���N��3?B?>���'�����=��Ó�=і1?�?�%���'�>+q2?��� $��x�=�ہ=~��>~x�>�Q{>r����m�HK ?�mb?Z�!��A��i��>�ľO�l����=�g>������[�>�xV=�$�����=�b��dْ��M?/�>u�&���$���%�,�,>�û�\?��.?�;�=�e<?��k?V/D�׹5�dai���)����E?R<�?��T> a0�8���U����>ݬ@?��>�4w=b�߾�����b?��l?R�%?]Ľ|\��8it��Nܾy�h?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>��������
>����W��?枏?�ד�������,��@o��bھ�?�=�f#>�*��L�L=������*�r/��q���X���̈�>�z@
B�g�	?�P�IK�m�¿�0~�bҾ!a��ז?���>�V���w��N���p�T�T�[��f����>>�>5��R���I{�Ė;��$��ߚ�>y�B(�>�fV����5����8<�C�>�}�>�܄>|d��������?]7���$ο�P�����K�W?���?���?{�?1�<�=x��K� �7�VSG?dt?-
Y?|e9�D`�� ;��e?lG��3�@^�S�=�i�>0�*?OD�>�H澙�2��zJ>�n)?��=&M������<���Ɋ?�O�?]J���?��?Ll?�Kپ���m����N�P~�=��+?1��>}#�@�%�Rez��fT��:�>��=?#N���
�]�_?*�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?ֵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>[H_���u>����:�i	>���?�~�?Rj?���� ����U>	�}?�v�>�M�?���=�O�>���=.m��T�o�-�>t>�Y�)_?�M?7;�>B��=h�?��0�F5E�(�P�pD�\�B��ψ>�h`?uDK?I�c>Lqͽ
�b�i� ���ɽ�D'�(D��׻@��1,�5�ҽ��,>"�:>��>=�?'վ��?=f���ؿf��K�'��:4?Yƃ>�?]����t�����?_?�{�>B�6+���&���\�&��?hH�?��?�׾I:ʼ�>��>#H�>�Խ�ҟ�vm����7>��B?#�]9��k�o�c�>� �?p�@ծ?4i��	?���P��Sa~����7�`��=��7?�0�(�z>���>��=�nv�ܻ��X�s����>�B�?�{�?��>!�l?��o�L�B���1=6M�>̜k?�s?}So���t�B>��?$������L��f?�
@~u@a�^?+�~߿�Ŭ�e���������=�f�=³>J{�����o�>W�<�-����~=�j�>~�}>/Ƀ>6P>��?>{s>>�R��:�*��G��܆��C��/�����Η������=x���])��������+���y(��������6�Y=���=;�U?�R?p&p?Oa?;gy�v�>�����	�<ܒ"����=�>�2?��L?��*?���=?��Ld��U���ᦾ�������>o�E>��>�^�>z\�>���:�7J>r;>>��{>\>�0=��hx=�,M>�ګ>���>�`�>�M|>�I�>Le����hY���F��_���?��C������j�����F�*� �=LFw? >�(��=����<L@?V��7e�v&ʾm({��'g?i��?F�+>��վ����~G�>F̀>�A������e���lY ��f?JT?�7�>t�>~PJ��2U�A�f��ٽU��>/l?���������@�̨��/����=/��>�|�?�2���O� ����;�=7�E?��>�<bV��W��� &�C��>^f�>��<��C<=��>8+��V����S�R/�>�h�=�j>�Z?
8>yIl=���>Ǯ���-C����>CB>!�>>�";?�Y"?���ߠ�$���02�=|Y>��>"�j>[� >͜E�庽=�_�>ˈU>o៼H.��m[���:�RdJ>\>���m���{�i��=��ýa�=2:p=M|�K�4�0V�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ٧�>�޽�H�������q�J�=��>�<E?���\�!�C�tT?Is?�U�^}��Jſ��v�OR�>���?���?q�o����A�/�|�>�9�?czW?�=�>��sh��u�>�R0?�OG?�:�>H/�N�8����>}�?�"�?^-v>�?$1?fi>If��t��oФ�nO��W�=�۽ ��>�Y>ȯ��k(l�����dH��=�X��x���>@lN<h��>�=�#��c(j>`��;ۊ�_�`��V�>[�Y>a��=ׅ>�v�>6�?=�%�>�l�=�=+��?�΁�#�K?[��?���o3n���<��=ȱ^�o?�K4?�s[���Ͼh֨>:�\?���?}[?�]�><��h=��_忿O|���<��K>_0�>`E�>�,��{9K>��Ծ&+D��u�>�ʗ>�ѣ�.1ھG2���U��5<�>�f!?��>Nή=�?�@)?�G>���>Y�1��w��XE����>��>�?M�y?N?�\׾��E��l��i�����Z�KxP>=
|?��?���>�]��)���D	�:�'<$q��U�?�m?Ȇ�����>�x�? s-? �4?&�X>� �۾��]�4�>s ?�F��tD���*�-�-��
?)�?J_�>�0P��Z�� ɼ������HI	?�}Z?��?Dl�	�a��B���G�<� ��c�<xv���%��>	�>�ض���=��4>�=7"`���@;�i�=�A�>�>I3 �� ���<,?�eG��ԃ���=��r��zD���>�@L>��Z�^?-L=���{����>v��^U����?��?�i�?e
��&�h�t"=?#�?�
?R$�>�M���y޾���Zw�)yx��|���>H��>Ôl�L�P���p���)G���ƽ[7����>;�?�?_�>eZ>+:�>����F�w��.Ͼ}aF����p��r�%���ֲ����������D;,4l���>�Rd��?��%?�>���>�7�>O$T�}>�!�>F�>}��>�>U�_>�5>p�>����NR?ك��2�'��5��#��e*B?�d?�f�>�h�x���B�׶?]�?SL�?��u>�h�+�׈?���>�:��$b
?L�;=%��|�<����Ah����[����>\ҽ�:�~;M�Бd��
?�?|���x�̾9�ڽo����o=?�?<�(?q�)�m�Q�0�o��W��S�]H��g�MI����$���p��폿�`��f ���(�9�*=*{*?��?������+�|	k��	?��Of>���>��>���>gI>^�	���1�r�]��6'�T΃��<�>]]{?��>7n,?��J?w�8?�n[?�>1�G>S��ǟ ?[�>gt;ѣ>��9?�(?�,?�|0?�Dh?���>Б}��������?&��>
;�>���>�B?�N�?�lƼ|��=������C��J	�~��=֖!=��V���e>+As>;J3?;�%�2�Ah�S��2�Y?��>a�'?�El��J�G���W"?ݩ�>����s#1��Ћ�������>�֓?f��<d���M�>؜>Ƃ��ӼA�>T�=���=��ͽ��k���.<X�%>��=U���5�<u�>��^>�nнkt�>�?6��>=�>x>��ͦ �����O�=�Y>�S>G>�=پ�}��%����g��My>u�?�x�?��f=�=[��=���W���������/�<f�?�H#?�TT?���?��=?Fh#?�>�)�L��^��r���?�*?&v�>�i����fs���y��?4z?5L��$Q�`p"��\��"cE����=u`�&x��㮿~)G�f�I���X-���?;ܘ?@!�$X,�����o��T{���"O?6��>��>E�?wa'���r�r����>a��>�O?���>��M?-l?Gۀ?I�#?*I�{&�������འ�]>J?x�H?�?)Z�?�"?�j�>���=����7�Bk2�g����ξ�X�M��>Q��>���>��L>4<�<M2���Ǿk�	�ʇP>f�>��>�ff>g��>N�J>P�<_�G?2��>�U�����᤾Խ���F=���u?���??�+?y=^}��E�g?��[M�>�m�?���?�1*?��S�j��=��ּ�ⶾ��q���>[ѹ>�0�>�=fnF=Hk>��>M��>��b�,r8��iM���?�F?Q��=aɿ��%_�[�q��;��
;"=��Ͼ³w���M��I���,�=ھ����>�<�k+�����.��M��m�Ѿ�u�� ?��>Q�	>Ǥ�=����;.�e�9=�4Y����l�=�o˼�1>I��=Z�C<�-<�a����h5 �9T�˾yg}?d�H?2O+?&lC?��y>��>�4�O;�>�ꃽ�7?LV>z|T��d���<���� ���fؾ�׾Pd�h���Y�>��K�D>��2>�<�=��<l�=�w=IB�=�^��=q��=�{�=_��=��=&~>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>W	<>�V>R�3�5�p}�v\:���T��v?֭)��ɾ��>���=#>�f�ɾZT=x>��<v�1�8:S��?�=/�k���=<h8=��>\�2>&�=XTý�!�=���=�R�=C�R>��D=z��t�e=ԍ�=?�o>�G>�[�>�j?W�5?��z? L4?\qw�����m־��J>F2�=��8>|n�=��>2K?H5V?�C`?)`?��>Jv��;h>?�b>�y�$\���ǾE+H�Ѓ���tL?X�l?G_�>� 9�����x�
�b�K��V����?&$G?dZ?4I�>�������� �t���(�`���e>��y�I��=P�>�İ�c����>;_�>æ >�~�>�6�>'M>��O>ج�>��>=M��J�;�?G;�d�τ%��ߍ<�5�%t��pW�x5>,J�>��>j�.��=1��=�Ľ�'S��>G��>�>ǃ	?Zg����9�>�꨾m�v��=��?1>���n�&�R���%��U_��C>)�<>�K��������>�7�>I��=�?=��?��~>�d���׵����d��w-y�2�8>Ë>3���ʹ�3�H��87�����1��>c\�>��>�<�>�Q.��D;�~2�=�ھ�b6��E�>��7�|�[�GK0�8jg��ꟿ3Þ��`����<��C??����G�=��~?"�N?�׌?s<�>�yŽ6�"��=�'a���Q=����E���q���F?�@(?��>m����O�H̾���}޷>UAI���O�`�H�0�z���̷�Տ�>c���8�оd$3��g�������B�EMr�%��>�O?k�?�9b��W��>UO�V���&���q?�|g?`�>�J?�@?�$���y��r���v�=��n?x��?(=�?�>c?�=`���?k?�X?R��?�S�?��{?�B���ߛ>h��;i
>�ϫ�L<>��E>ju-=a�=C?8�?�+�>ǥ�Z������^a��4��<k��<g-�>�>���>�
>�k]=�m�=�8�> E�>�h�>Ɛ�>�:�>a	b>#��> ��u@?��O>��>=[?
m�>�}R>�a/��� >��p=l5���6N6=96G��NO<E_�=�4>+-M�,>�>��ƿ��?�bH>_/־�=�>��J��?ѽ�`�>Ee�>'����.\>0�*>\S�>��>G�?��b>���>Y�~8��)(v>�c��hF�/�E�������s2>�W����ڽb�	�V�NQ��G���k��%+g���s��8����<#�?�����r�I�&������?G��>d�T?�����(N>�>��>���̄��w��^��?\��?�;c>o�>5�W?��?�1�3��uZ��u��%A�e��`���������/�
�������_?��x?�yA?�<:7z>���?n�%�?я��%�>1/��';��<=-�>&��x�`��Ӿٸþ�7��HF>��o?	%�?5Y?n]V�ŋ��BT�=�4J?�p.?�\t?�C??:�U?��m�"?�4R>��?�z ?�
0?{�1?�$?��l>΁Q>V'�=�B�<% ��͚}���������E��	q�=�V.>�=��=Ħ`= {u=}C�<A0����*���	�:�=Sb=ļ�=R�8>-Q�>�8;?��?*��>V)D?5!���6.�+���I?�~o>!?Ǿ����zo�����d>���?���?�fe?�s<����<��| I>ƽ>��@��.�=6�> �1�����&�=�*�>����|�=��_�3�:}=�%y�� ��1>̾�>u�}>ʒ���">Q��TLv�V<f>��R��p��E�V���F���0�!�{�:$�>E�K?γ?�Ǒ=v��¶��d6f���(?�<?�M?��?7�=Z�ݾ�%;�h�I�9��aQ�>���<|���T��(F��@':�a�;Eq>�-��cg����>�Ҿ���:h�x�N����P)�C���$�:nz!��_�~q���>Ң�>&���>0�����<���wC?d��='�;~��W��kO�=k��>?~�>�*�����h}=�� ��@1>���>��k>}=3�ѾeO����V�>��=?Zu?I�?f�ܾ���&����JV4�8�=���>F0A><�?R1�=��>ԡz�x�&�nw��M��S�>"K?.��&D�r����vA��S��>�(�>7a>5s�>3�?�	?�.^?�?�@?���>�0H�=E����$?��?�B�=pm`���h�L>�U�#�d�>�j?�wk�ɛj>I��>|b#?S�2?IO]?N�?�H�=�S�mlQ�^��>���>vGb�f>��c>b�G?���>z�b?�v?��1>���ʌ��b+��>/
>��)?
�.?�?�ٮ>�D�>�3:��񋼥�>�c?�i?��l?� ;>1F?̿n>�H?���=j�]>�H�>���>ο^?m�?3)J?�!�>��;
�Ž�����ԡ�U';��<�䑼�Y=�$�;�<�M��Xz�<����M���Q����z =8g<�t�>����>e�i>(����>���}�_���Z>��K�m&��R x�;�$���=�`>���>�Oe>
W���=j��>���>�7�1?��?�-�>E�1�Ԗe�/�ؾ�F+���>��=?�e>R�����m�z���=��u?��Q?���^���b?��]?�S�=�
�þ��b��v�j�O?��
?��G�^߳>��~?<�q?��>��e�15n�p��Gb���j����=Um�>^W��d�qE�>{�7?_F�>��b>��=�۾M�w�\v���?��?���?���?h'*>`�n��2�������:#^?���>w����"?p��N]о�W��l1�����z"���~��m����N���E&�#��.3ؽ�8�=��?��r?6q?��_?@� �]�c��^��	��oV����t���E���D�X�C��an�|[� ���������J=����7��d�?��N?/2l�q�>�����9�qǩ��Q>�^㾢-t����=5{���P>%I�b���(������?���>d'>�=?�[����5� �¾G=��#z�IS>��g>�8�>Bi�>�,1���[������6��*�ʽi@߻�T�>s6?v�~?��?nm�R2F��f<�zVA�cN�=g���
"�)�H�d��>px:�(��=:t�Y��� ���=�ʹ�<O���a>V��>�p&?���> /?�
?�L�y��z#���7
�����ǆ�>5yu?k��>�S�>b����3F�p_�>
�\?H�?]?���;�A�,t;�[Xž���>�5?�&�>p�=?�<QH���t��K�S��$���E?�;���9T��.�>�?J?h�˼��<��[>k�&�0�����d菾�">Nv?�J8��wN>ʻ���|E�Q�����轕�(?�m?� ����*��N>_� ?� �>��>���?�!�>l"��\�0<��?$B\?�^H?]@?���>|4=�ڭ���ƽ��)��>'=Cm�>V*U>�{y=���=+����]�����N=Э�=�ِ�����
�!<����*2<D��<�4>�{߿�WW�Z���Xt�ڇܾ�;�ʒ���rĽAY��;�{�C,þ�����O��j���Z瘽�3��%�~�j���u[w��j�?Jj�?���"뾇9��	[������>���M9�������C$�u��z
��C�GY<�N8f��6`�9�8��&?����wǿd���6eپ�S ?ؿ?�Ox?�����!� �8�}a%>�o =2������-��'Ͽ���Fa?�p�>�Q����^6�>�"�>��X>��r>_~��}����<�a?w�-?{��>�m��Pɿ���#��<�x�?Z�@�@?#'�v����;=xI�>�?��r>r���-�zO��~��>�j�?�؉?1�=�W��ؕ�`@e?c��<'4�Y>��x�=t��=�;�<t���/>5;�>h��bO/�y9�s!>��>dp�ɭQ���z����=�m>����L��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�󉤻{���&V�}��=[��>c�>,������O��I��U��=���4�Ϳ���	��7�<��(�"Xս���w���R��u��9m�NL�%>`�=��8>`Ez>�:>�>g�T?,?���>�j'<O��� �d�)n���>m1��`䑾��������ؾ$|��!^�e�Z�%��#�ݳþ�=���=�3R�򗐿�� �o�b�:�F���.?#�$>V�ʾ��M�
7.<�yʾ����0'������F#̾��1��n�]˟?��A?G���6�V�����[��f���W?CH�$�� ᬾ��=�α��s=�>���=*��%3��{S�f�?	G"?�O���ᾓ-�=<�7�Z�>[�@?�#%?З�=zR?=�'?0b;���������>;�	?���>;��<\�l�vʽ/��>�y'?Y��8 :�;>��ɾ0���Y���O_o�EaǾ���=���>"���X�%w�iV��/ȼ=��A?|��=��O���.�S��ƣ�>��;O��?8�v>Ք�>AsL?R�3?�o��m���G�������I>��l?�gZ?��\>����_����U>�� ?9Ih?��f>�v�y�`�2�-m������o>�?�%J?�\d>����H��?���%�N?�)]?6�;��˞��o)�+�ɹ�9�>��]>�/?��0�#�>^p?���=�����¿9�A���?�@:��?] �<���R��=�]?'k�>���s��~������s��=���>C��o}r����f%ݼ�0�>	Z}?Fj&?s��zG.�>�h��O�?Ip�?�ξÐ;���	�x��쾶�=�F��:��6�(������XKپ���0V�`����>I@��.D�>횼����������u���\��~��A?8��>�x��Pľ��D��nY��]6���3�$V���>kL>O�I�E�B�tw�*E�V@�=�8�>%��'8>?T��V޾Q�H���=:��>O��>�<>�xg��9��?�Ӿ��Ͽ�ě��r���M?%�?r �?�5
?��@�*���8��l7���jN?3�`?B�K?��=�MF�Ə��r�_?�7��@n�\�(����@��>�!K?l��>�g_�\r1>�~�=f��>�S,>0�V��?��`<��hV�?��?O�ܾ��?�#�??��>�b$�!���ҳ�����^D>3u?C�0>� -�`?�R�m�:���72?[?Q��
�&�[�_?!�a�E�p���-���ƽ�ۡ>��0�
f\��M������Xe����@y����?G^�?`�?޵�� #�e6%?�>W����8Ǿy�<���>�(�>*N>�H_���u>����:��h	>���?�~�?Hj?���������U>�}?�A�>���?���=?�>a��=^~���A��� >8�=-G�l�?��L?�(�>���=�9��/�!�E� _Q�Y�UkC�$Q�>%�a?�"M?�h>���H�G� q!�aqսpq4�1��Q7D�Z�(���׽�?6>�k;>>T�C�s�о�� ?e���Ͽ)ś�[���A u?��>��>�����ƾ��R�
mn?�">5�jc�������/��ʦ?*��?�?��a���)�:�	�>���>�.���=�ZU���=��5?�@=�����7n�z?P�?yk@���?qq���i?_����bς��]羺r��tX�=�??K��;_^>ޒ�>�PE>*�}������+l����>��?Q��?F��>|e?��\���2��0=�v�>EQ?��>k��='�޾q>e�
?��Ԏ�ȸ��uT?�H@��@�u`?f���D�ݿ�d��T_���u��+>��8�;_=�
�4�&>�ـ� ͽfR��M,>t��>G;�>kFo>.(>��>n��=�܊��2.�fD������g:�"�@��4�ϱ��������vX�,��t����	��Ac������?I�r�P���^;��#>f�>?L=?U;s?��.?�v���g�>��ʾ˹��B���O�>�����Z?���?���?�b>Y��j����w��%⽾3 ˾���>xȟ=��>�Q�>�U��}
��t�>���= a>An�>� >�y<��=�͛=��%>m�>Dr�>"�<>�Z>բ��G����h�Փw��ǽa��?ܭ����J�.���ύ��@��|F�=Y�.?�,>f���IJпj��zH?T����\�N,�ҁ>�0?aW?a?>� ���xT��t>�����k���>n �#�l��)���Q>_?�g>ͧu>6r3�i#8�H�P�����7�}>�.6?+��W�9�`�u���H��ݾ�GN>%�>sY=�oO�����4��Ui��N{=Y::?�t?���������u�	8���Q>� \>��=Ō�=��L>k�c�pǽ,-H�Y!0=U�=��^>�
? Є>���<e�}>�~���@��:��>�@>z�5>�m3?I�8?�K�)傽E�6��'���8>���>Vb�>[�5=�C�e�>��?���>�I�K��[*&�N]��#��>�;ս��� ���?�=�ض���>$���n�����-�<ϖ~?��;䈿2뾕_���mD?�+?�=F<�"�z���4K����?P�@Dl�?��	���V�m�?�@�?�
�����=|�>U׫>ξ|�L���?��Ž�Ȣ���	�#(#�S�?X�?��/�.ʋ�6l�g9>]%?�Ӿg?�>�
���@���$��2J=�b>sĵ>��*?�������팾�5?]B?����Ѭ�؄ѿ ���R�>�+�?���?)P�䠟� �%��n�>j�?�cN?�?m>�Ҿ#&��s'>�hA?J>?/G�>bx+�����??ǵ?��?�M>��?�u?���>ʅ���53�5/���ݍ�.=�=�p=��>y�=�M��ǿG�/^��8��\xj�Y=�/b>��'=�6�>=������ɖ�=i��:|��Vp����>K�k>&(P>�>�6?�z�>pw�>C
=]죽����ύ��kH?E�?T����UD������E�;^�M=c/?�?L�߽3yؾ݂>�ER?_�?Ұn?�h�>hC�"U��ݯǿN���!�<�S�=1��>խ?c�=�3>����$ba��9�>���>�c��!���M}�$�����>B�1?�3?e�=)� ?դ#?'*s>.ߵ>.cH��ђ�I�C���>B	�>n?��{?N�?��44��n��$���[���G>��w?T?�v�>R���rd��ƍ�'/G�K�x�(��?��e?���%o?7�?x�@?j\A?�{Y>+��1۾�����>F�!?��qA��D%����?R�?�A�> ����ڽ�-��������?�z\?�/&?l3�l{a�z�ľ(��<(����ػ*�;�����>{>H���l�=�>9��=+m�q�8��+n<=���>�%�=�3�l���O?�?�9�P��-��!|?��45��@=���>�B���O?��o���E�zி�u���ʐ��R�?���?�%�?�,��z�j��B1?���?�h?{l�>,��I׾�G꾚f	��(2�y)�O�>�>Tv�=U��:^��#��<B����M����|Z�>u��>j�?Y�?2;g>�C>�G��+�#�ҹ�a�G�V��D�����h�$�s�ƾ�^^�4��+ľH��QD�>j��_�>c�?)S>I�T>��>�������>ʝ�>=�D>Կ�>z�w>=N>�w=>�~U�="���Q?����)���1��&�D?Pd?���>;���!=������9?Bܑ?
,�?��m>z�i�G�'��p?�c?s~��x?��==�Ѷ�ǆ<k������H��^���r�>h�ݽm&8�ZK�C�e��O?<?��V�>fξ�GսB\��r=V=� �?K�/?�1�=zP��k��]\���J����-	���ș�S"���s����ݬ��f���yN(��x�<�(?l�?�����*ɾ�av�9���g>7�>���>϶>�/6>7���3���Q�]���y��1�>�wz?u��>XF?�$?5�9?�a?�c�>�->�Ծ��>���b$>���>�< ?[�E?�m?-Q�>f[	?9`>��a<����!⾓�?y�7?\�(?�?6��>d����N��bE�߿��A���C�<!ƽ=�t�=�� �=����q=`�p>�?��-��gP���ѾX�>BIr?�?� �>�)���~��8=�-;�?�O?�^�����>����>p��?�������6 >��>k�=���"ʝ>��<SX��~�=��0�k�>R!>��=��%�v�=Ί4>��Q�M)q<���>��%?��0>n�Q=��K��e�24	��Q$>)Y�>7;�=ȑ>nkR���������1W��U�>`}�?]Z�?��ͼǖ�=�$�=-󻾗;��B��?ۈ�#��<T�	?�L5?�P?zT�?]�@?[�?��#>(9Ѿ�����y���y���?�,?�j�>��;��?Ψ���4��?�>PBZ�����"��ϾM$����">%1��{������_A��*n�F��;���%0�?�P�?��a�/4�c�ﾸq���襾Tc??��>p�>h��>e.�O�a�60��%
>�^�>$<Q?͠�>�?O?"~{?�U\?}�P>s8��ᬿ�̙�i���N!>-Z>?.&�??�Xx?�S�>p>90�������G#�������R=�+[>�̑>+��>��>p��==�ѽ����?��_�=e�c>k��>�ɥ>���>\Ep>&��<f�$?p�>9�¾��4��L���n�@��[?\l�?D�_?e�<S?���Ip��y���>���?��?�1?BC�ήn>��F�e��#����1m>���>���>3sv>D���J�=��
?%l�>ii�����u�A���=^?�~N?�~޼��ÿ��q�?L`�<y�����<s����pt�����yZ�Y�=�m�����
p����V��曾ϑ��F��$!����w�RK�>�eo=�@�=.��=@�<X�*�h�	=C�=܂<��"=,U���<	�,��B
��<����_��|o<�F`=@k!��ʾ
}?��H?�i+?59D?,�|>�
>�?�K�>+⎽B?�T>9L�Ք��H�9�]5��ft����׾�վ��c������>6`C�դ>�o4>z�=��<l��=C�n=�ߓ=q`s�T�=u�=�=��=B��=��>�>q3w?=���k���N6Q��3��:?�)�>"��=<ƾc@?<�>>�.������c��%?���?�U�?��?'xi�8Z�>����NĎ�gq�==ɜ�]2>պ�=D�2����>$�J>ł�9H��S}���3�?��@��??#⋿âϿ�c/>��7>;*>?�H�AN9���=�`i��J)~���?�>��Xľ� �>�T>h��q0վ��d�7�V>CF�=P2��cP���=���kP<��[<T�|>�XA>�t=�����l/>ι�=�q>��i>��Ҽ��⼕��W�=�U=��d>�->I2�>�>�>�g!?��<?&��>�		�{<�( ž��>��>�o�>�s����1=U�>�?�Z?�3?6a�>�	�=A��>���>^���j́��W#�4!��	�<ѐv?�Џ?5k)?X>c޼8�2�VNY�[P���*?�7?�q�>D�@=�n����Y �/���\e��<���|�a�� �<�rj�$����D�=X)�>�~�>˖�>L[�>�E>a��=�L�=!:�>��>hJ���/�=K�+�
&y>��,=���_b��<�n��x�=b_j�rO較��<�ER�i}�<3�g>��p<�X�=�#�>%a>P8�>���=�����,>�K���6K�5�=������@�tc��{�AO.���8�A>mX>+ju�(����?�^>�{G>7��?�0t?qF>X��̜ؾ���� t��%\�qɸ=�&>l�9�b;�]`��mL��6ξi6�>��>A$�>tȎ>!5�_	C�O B=��쾍,��V�>ܛ��杽���\�f�����W؞�u�p�>o1�P<?�
�=��?Wm>?"�?S��>a���9��s�>���I"�)��-oy������ ?��!?���>a���p�A�+̾����Ʒ>��I�n�O�}����0�7��v�����>D��]�о63��a��'񏿙bB�`�q����>�O?��?�a��O��BRO�C���#��K�?+tg?�)�>^Y?/M?q���u�֝����=C�n?~��?�2�?2�
>���=L���C�>�J?���?>x�? Z?�kd��V�>I��z��=��%$>�K>���=9?b=�,�>%�?�w?�ٜ�������.��s����G�/5�=�ߢ>Ԧ>�ժ>�'> �<*�=Y�%>��>iH�>� �>�!�>.qe>ol��:E��Y8?[�%>ZT�>K�-?f@K>(t�<�R߽k��;����<�Z�(������n�F�����S�D�V=&��g�>��Ŀ�n�?�C><Z⾽^ ?مپ,瞽�J%>o�:>����>J�7>��v>5F�>�j�>�75>�>y�	>C�d�=���ƽ.�#5��� ��G��('>U��Pǈ�,A
�fP'��;5�Ϗ˾���޲��l#��=�+����=u�?rg>���گb�$���;?D�>k!!?��<�#�=
��=��)?� �>	�D������c��Ŵ|?��@VLc>T�>K�W?��?B�1�E3�zqZ��u�� A���d���`��֍�����Ӗ
�~d��m�_?��x?�aA?�[�<�Ez>���?��%����)��>0E/�n;��<=͈�>ڕ��M�`�W�Ӿ��þ&���&F>B�o?q �?tM?ZZV��	S�"�*>7?�d0?�w?Kz6?��/?^)��t?�q�=��>��?uc4?�q2?\Q? X>+��=%ܡ�-Rh=o<��h���o�ͽu(���ZI��PQ=Һ�=�D<�<�Z+=Z�,=P����{ ��֩��(�<>�f=��=�x�=�D�>��J?��>���=?n2?JE��,D��a���`)?���=D����(�F��Jv��V�=�e?D�?yFX?�p>��A��d���<>1�A>�4�=��[>�1�>(sa�k�޽��>�>d��=��N=6����X|��� �YA��h��)@>��>�'�>��o��F>Oט�^~��j�>�-�:3Ⱦ8�x��<@��;��@c����>.mS?�� ?L��=�������_��.?&k,?�G?�ȃ?3��=%�꾒�7��H�r�>��>K/=����ݞ�� ��k�6���<u�> ���U��a�e>c�
������i�5-K��z�k`�=�����= ��
վ�)��F�=�t>	���:��8R��{���G?Y߅=V�L�䱹�P>�	�>
�>����H��A�=F���=ݟ�>$C>�*,���lG��R��K�>�H?�`i?�m�?�7����n�(�7��?��[��Ň�t?�0�>;C?��a>%��=	ξߍ �m���/���>���>���]:��B�����+��h>3�?p�=1�>`AF?�?n0b?i�*?�#?ӆ�>���%ػ�@�?��?j%j=�)!���:�q6���<����>E*?���)]>e��>�8?y,?�$L?�7?� 	>���1�e��>C:�>zM�ʑ��k�\>�Q4?j1�>�PX?C��?ռ0>.�>�1�����*+>�4$>ɪ3?qR?qL?M�~>�&?�㮾%����>�bU?��?�,n?�<�=�<�>9�+>] +?��>g�=�>�>�M0?@g@?�@V?�,?SR>Y!=���(dL�O(�����=y��=��=�|�>�Ȥ=;0���_>���=�[5>��zH	�U^��x_���m=9v�=s��>�t>a핾��,>��¾$ԉ�h;>m�U��陾=���Kh;�		�=%9}>HS? ԕ>}x �b}�=���>;��>�����'?.M?��?ua�:�2b�9Iپ�K�^��>��B?���=}�m�����ùs��oo=4�m?�~]?t�Z��t���b?I^?��"<�3�ž��c�ך�C�N?dw?=�H���>�^?[Mr?>B�>�)e��n�*K��$�b�_j����=���>a�zd�S+�>�7?LF�>.yc>���=�
۾��w�*/���L?��?a�?#֊?	�*>��n��C��?۾a����\?�B�>%����5)?	WH=��t�|�BUw�h{޾;���J���V���>�����-�n��m��|b�=d,?}i?�Mt?؎[?�����f�2_�dw�dOT�g������>�`73���G��+k��$�o�c
��_��=�H�m@��;�?�$9?*�N�%C?��0�ZQ�'_���3]>S�|�Q=B���p>�d��m�����卾^�i�a
����?�>���>�)5?;z��-���1?��ľ�*Q>ڂ�>�K�>��>�8��j5��ӂ����¨�>�鼤k$>ȍb?_#x?�r�?�|Ͼ�"��uu��};�4�[>lɃ��=�Y2>�)?5�
�
a��4iZ��p�Gώ����u[������5�=��>OF?dM�>"S�?�I?�Eо�n)�*�Z����ӽ���>�xD?�>`w�>u�ʼ��)�	��>��`?[	?z��>������ ���u�-ك��G�>�Θ>��>#>��b=Ks�=;��̿��p$G�|�;�]?򦾊s�r��>�:9?��0=[�Ƚ��=�==at�_���k]轍k�>�q
?��q>|>�F	�e:�;���5��^6?DE2?�����
&����>2��>I�?�f�>�sg?Ա>� �+�³>�j\??0M?l;?N$�> ͋=����1�<-GK�h���l�>OZV>���=�f�=Q��a<��(�����)>I�d=`jm��s��W�=�=�=�ڣ=ԾL>�bq< aۿOK��Lپ�P�����q
�A4��孽2����X�5浾���rFx�ҟ�+�-���U��/b� ~��
ym���?��?⒓� ;����������% ���:�>�fo��>��Ǭ��Z�qK��G�ݾ\���a�!�cP�,�h��d�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >WC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾s1�<��?7�-?��>Ǝr�1�ɿc���z¤<���?0�@�D?r�)���;��=�?�> �?ʁQ>�(;�- �U�+�>���?'S�?δ.=�M�$U7��Pc?�<�cD��/ں�=�<�=$b=��]>ۊ�>ڱ��8�쎷�4�O> ׄ>	A;�B�2���Z�e;�zL>(��Ժm���?�{U�Ԗ^�\10�Qj���>��P?�w�>J݁<��8?5�*�S���pVa�p%Z?'��?�$�?<�'?���&�>^�t,Y?��0?7�P>�G��~��A�=��нc ?;���A�l�a��<�#�>�q�=4^k�37	���.����~>���ixƿ��$�q��.�=���P[c�-彦����JW�4󟾏n��齴�a=�W�=.R>��>�`X>��W>��V?��k?rݿ>ſ>�罯�����;�a��N3���;�<���8����뾄3߾ţ	�F;������ɾ��7�./�=��F�哒�0���
W�bj^��U9?�[>�m���@���4=��ɾ����i�#���Q�I�q�n���?h�G?%IE�if�~��0���;|߽��^?a]<�����پLz��U�_=��>�d�>�<����Z�2�9���E,?��9??ٶ�4c�,�>X
?��PI>a�9?��>w�;�>R��>�J.����2/�>�O>5�>���>T�0���о��Z��1?wJ?��ƽ�{��hj%>�K.�'M��r���G�<�|����<�f>�L׽l��FV���V��E䊼G'W?Y��>��)��pS�����}==�x?��?y/�>�|k?��B?G�<�^����S�����w=}�W?� i?��>�u��оI����5?�e?��N>Jh�F��?�.��L�<"?��n?�Y?����hs}������l6?�?�#o������l'��>+lF>���>מ"?�4e�f%�=U�?G@j>_P�����d�>�,,�?�P�?g�?��=����l�=~_�>��=��E���j�=P����>�S">�a��B�����4��A:?7�=?e��>��Y�28�.k>��X��q�?|^�?a�jZ9=��о燊���m�`]=&>^I>V�>>
?��%|*�����8�CM ��F�="�>@�k����>���Wֿ�����$����b�8������>
2�>��;F�E�)2,��|�uu�p l�I�J���r>D�=>�M�2�Ӿ�E�>�K��d�� ?�Q�=�r�>peӾ� �zٵ�42>���>��
?�֐>��F��&�����?!��Ah���Ή�&�־��R?�u�?�j9?F)�>.l>�+�HD���h��t�-?Đ?r|?�՚=�*��.x�%�j?�]���S`�$�4��HE�+U>�#3?[>�>�-���|=)>��>�l>�$/�7�Ŀcض�X������?ˈ�?�o����>s��?�s+?�k��7��)Z���*�҅-��=A?�2>f���̶!��1=�bՒ��
?o{0?x���,�>�_?�a���p���-��ƽ��>9y0��b\��/��J��Ce������y���?�\�?��?*w���"��!%?
�>׾���$Ǿ$��<懧>EM�>_/N>��_��pu>�����:�Q�	>���?Ol�?�V?�����樂6e>�}?;7�>5�?D��=H��>���=)^���B� �%>ރ�=�&J��N?�oJ?�]�>`m�=�G9�R�.���E�:�P��F��wD�.w�>�+b?�1K?�qe>C�ǽ��5�#F�)��;4��o
��pF���:��ڽ�`+>"�;>K�>��F��Ӿ�b�>9*#�B�Կ޴���
ཛ�?�[�>�B?���<�=9�yl?�xg>y�)�)<��G
p��N��O�?�*�?@[?<�۾9޽*z�>���>p�>�=d��<�����GW>�� ? ��<�Uk���~��9e>���?�#@y;�?�����=�>���R�����x�CV羮�A��&>��7?N2	�n>���>=�&>h�i�|��M}��ս>A�?."�?���>��d?��k�82��Ly=Y@�>0_?���>��<�����>��>�N[��T\��V?7J@\P	@��Y?��#������a_���򊾥�=��	=1��=���#��<mp�����Lf��=;>���>���=�j>���=�B�=�z>������#�X��@?��QOF���A���J�d�X�̼�Y�r��&�0ܾ������t����	X����HW���<[D�=9T?	�\?Txw??D�>T0����>!�� ��=߆��=$�>kU<?�M?� ?ϙ��N!��ɦl�Oށ��Q��Ha���5�>*}1>$b�>��>�r�>s��<�>"�;>L��>��=�g<xº<>�R=�S>�Z�>��>W�>bD<>ǌ>D̴��0����h�[w��&̽I��?�}��ŬJ��1��,L���֡�=�g.?5�>��}9п�\2H?�	���,��+���>��0?�iW?�a>�-����T�&Z>�����j�	Q>q���Krl��)�Q>_e?Ԏ^>�_x>2���8�,M��J����l>E�7?Ƽ���>��t�߮F��ܾ�ZP>�H�>\�7�Am�V��*|�	qg����=a�9?��?�������,u����%4\>i(Z>���<���=�R>i��$����YE�\=���=��g>���>�7{>jN�<Gu)>�5O�	�;�E��>�3>��{=PoF?��?� ����a0�svڼ�r�>���>L
%>�O[>YF��"�>xS?J~�=G�����O�O��ؠ�>�͗�
��� 3�:S�>񄍼�J)��ׂ��PN��O�ʑ�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�-)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾÞ�>��EZ���"���u���!=�=�>�H?~��I�L���=��r
?��?VZ�@�����ȿ`v���>{4�?�
�?��m�Kl���?����>b��?��Y?d�i>Z[۾y�Y��׌>J�@?��Q?���>����L%��o?���?���?�-N>�H�?z�}?�q�>y7��c1��Ƭ�˔��+>�]㼤a�>l]>�+��Ta3�0݌�����<T{���(���r>�61=.��>���F����=�ͽﹾfr8�>�>��Y>�m�=�w�>Mh
?B��>Yt�>�a=�%���H������]JK??r��E�m��.�<NՕ=��X���?m4?�o�a3Ҿa��>	9[?���?�Z?t�>�j��.���s��>�<(BE>9��>���>2���UK> �վ�iH�맇>�,�>9����۾�Ã��'-�Ϯ�>�� ?��>4Ѥ=�� ?�#?c\k>�n�>��E�0��%�E��"�>���>m-?��~?b%?:l��.53�����*�r�[��DM> y?rK?��>񇏿�f���P��K�D�����?��g?j���?�)�?��??ͧA?�kf>�y�l7ؾ@ծ���>v�7?�о��;���� �*=��I?4 ?�V�>�G��r��=H;�>|�ᾡ:>�� ?1؁?��1?28\�-��޼ʾ3!?=���#�<Z#�x��'܆>Z�>�E1���]<�uX>g��=�^�Խ�� =��x�ީC>���=��7���9=�*?:�M������J�=�Oo�u|?���|>�A>����[?d�;���x�k���������]���?O1�?d��?��Ľ|�f���<?�O�?�?���>[2��7*޾��ݾg�m�b�j���2�=LS�>�*��+澞���%U��Iń�����м+����>��>�?�D�>��&>)��>Xp���l�A�Y����%_��	�n�2��@*���᥾=1��Z��s#����>����Z�>~�?m�I>66>�Ļ>PÕ�en>�Y>��>���>��L>��K><o>�9��`#)�$MR?����^�'���I���~<B?�nd?�5�>&hi�\���_��K}?<~�?�q�?yTv>osh��%+��h?;�>g��6v
?;h:=��̔�<�_��~��@@��t�����>��׽�#:��	M��if��d
?�.?������̾w׽v�ɾo5I<��?�P%?�r(�*�U���w�\�T���R��Kc�uH��Ħ��A �Kbo��������쉄��i)�
B�=*"?�/�?��\������yp�>�D��kz>��>��>~I�>�K>%�
�8�1�/d���,��卾��>h^?�y>�P?�i.?pVM?BE?���=�s�>�pg���?�ڦ��K�>}�>i?aR"?�'?k�? �?�#�>&�G�_:���뾁 ?�<?z��>c��>W��>�x��B�ɽ��<���	��ȫ��`��>� �c
�׽�Ԗ���<T�>�?����8�O�����m>�:7?���>4w�>���#���h�<G��>3�	?$��>�	 �.�p���
���>�)�?1��7=��)>��=[]�>̹���=�������=�Ǜ�C6��<ȇ�=K��=1�˺��S9"�[;��;��<[��>��?ﻊ>l:�>�����.������v�=H|Y>��R>"s>$�پ�ۉ� 8����g���y>|W�?X=�?S�c=!
�=�f�=ݩ���ƽ���k(����<�<?��"?F�T?�!�?p=?��#?� >	��q[���u���ԣ�v�?�$,?)��>6���|ʾ�憎�k3�=�?�??G*a����64)�>�¾ZԽqH>Pb/��~�����D�~
����rv����?~��?��B���6��l辗����^����C?�>�E�>+-�>�)���g��5�V�:>�U�>J
R?�-�>�Y?s�?�r?=����@����F:��?�Y>���=�?tx�?�S�?�[�?d��>��#��h��.� ������e�wEཁb���DW=J�>���>H%�>-�>(��=�LM����C���Ǻ=�>��>E`�>]n�>�u>��:�La<?&ѹ>qǾW��[X��5=��bo���E?�ee?~�?��>���*��M�9F���r?�ۤ?�#�?�?��c���U>J�^��оŊT=b�>]Y ?G��>�r�g���]>s�?&�>4�s���~���u����	?��3?���<5Ŀ5�m��Sn��v����<�y����r��b�� M����=�圾���c��d�R�5n��l����������a�w���>�j�=�� >��="��<����ܶ<;+Y=T��<�|==����f�3�5�E�B<�ch�&�;Y <+�=�<�6ʾ8�{?�8G?�,?1@?�@T>�+%>u�	�f^�>���Sh?B�&>N�[��~��V�4��b�����оi,׾?�g��j��nV>>���M( ><J>'�=�ļ���=��`=C�w=��D��?=<��=���=8��=Ϧ�=��=��6>�1w?���S����3Q�Q'�%�:?&0�>pí=9�ƾ�@?%�>>�0������sP�h1?G��?�M�?�?�hi�.e�>Y��������=}ל��F2>s,�=��2�{�>r�J>�{�&E������)�?��@�??X؋��Ͽ�c/>b�>�;	=��Q���-��7�<�BN��IG��V#?��1�WC徿aW>�>%4 ��n۾&��<p��>��|>D�>�@���=b���ݬ=���<�_>�`)>n�;�� �>I>�<�sm>�<�=yj�;�j=Uw�=,f�<� D=�=��:> �>9�?_9/?�ub?��>�e���о�fþo�>&ح=%�>>Fg=u�B>�x�>��6?�0D?��J?���>B!�=���>�ţ>�+�u�h��;�ɛ��	��<��?[Y�?���>���<�:�����>���ͽ؃?1?��?���>�U����9Y&���.�����/5�g+=�mr��QU�x���Tm�0�㽨�=�p�>���>��><Ty>�9>��N>�>��>�6�<up�=�������<� �����=�����<�vż����v&��+�쏦���;���;�]<��;in�=���>� >[]�>�=6����.>X���@�L����=�0���B�M%d��=~���.��6�]�B>�fX>��D)���?�;Z>��?>z`�?�u?0�>����yվ�H����e�ّS��g�=�<	>p�<� |;��b`���M�2OҾ 7�>��>���>�s>M4-�d3>�@�^=�q�5S4�yq�>�G���8�V?	��Iq�;���2��@�i� �{�C?�2���e�=C�}?4H?L$�?�X�>}♽#jվ��2>�ρ���=q����o��:��z�?�?&?
�>�$�"E�+��YB�X?E>��¾�CI�������R�IO<= ޾���>�V�������"�`8t�f����i����ݵ>}�?6j�?=�T���X�伾HVL>�??�Q?d>�]?�O?m�,>Am�����>
�v?yW�?���?��r>D��= 6����>Է?V-�?H��?8s?�>�I��>a�;f%>ݵ��j	�=iq>6��=���=�g?+
?�n	?�Қ�������I���\��
=9�=x˒>��>*p>}l�=�Co=L�=f�V>~h�>��>r�b>���>;k�>���������:?W�u>� u>� ?BQ[>������;U�_=Xi;�Žû*=y�.��}��������p�ѽ�"�>
�>�����?�	>��پ��"?�禾V��c!B>]1>$�o�Я?��E>�n�>MD�>��>��>��|>K�N>��<��j6��g��w��z>�_�n�ri ���e>$:���2@�]���1�n|�t�ž;�!���u��V��m�<���8>��?^��$z���&[�
�F�-h�>o�`>��B?����K�=���='��>W�;>����?����쒿Ҿ���?��?z�X>\b�>�JM?_�>T/-��&�O�_�\�l�E���6h�;����W��jǾ�����T?fT^?0'?c�m=)��>�)`?�71��'��s�>�ھ4�F�7p����>����.�k�����1���K�#��ZP>��g?�z?�?����5i���'> Z:?�n1?�t?1�1?��;?�~�o�$?n�2>�[?�/?��4?��.?��
?]72>��=���vr$=Mđ������kн�GʽI���3= �}=9�#:��<W�=�	�<�Y�C�ҼwC!;�J��O��<:=���=�<�=(-�>��S?d��>�Ϣ>HV&?#����*��1ؾ~�(?J\��\�Ґ����m����\�=�
c?�{�? Q?��.>ˣ�Rq���=>��>Ql=J�>p��>�	��o��3>�%>��>�9k>�j� yȾ����E_�ۚ�=��6>Q��>�~y>Y��҃>x��rb��Ti>_O�(.��#WI��A��;2�f^��"��>��K?�'?��=�������o_��V!?�7?�M?w
v?�;�=V�ɾ�@;�u�J��#��A�>�<�<5 ������Չ8�j�;�gw>q��cg����>�Ҿ���:h�x�N����P)�C���$�:nz!��_�~q���>Ң�>&���>0�����<���wC?d��='�;~��W��kO�=k��>?~�>�*�����h}=�� ��@1>���>��k>}=3�ѾeO����V�>��=?Zu?I�?f�ܾ���&����JV4�8�=���>F0A><�?R1�=��>ԡz�x�&�nw��M��S�>"K?.��&D�r����vA��S��>�(�>7a>5s�>3�?�	?�.^?�?�@?���>�0H�=E����$?��?�B�=pm`���h�L>�U�#�d�>�j?�wk�ɛj>I��>|b#?S�2?IO]?N�?�H�=�S�mlQ�^��>���>vGb�f>��c>b�G?���>z�b?�v?��1>���ʌ��b+��>/
>��)?
�.?�?�ٮ>�D�>�3:��񋼥�>�c?�i?��l?� ;>1F?̿n>�H?���=j�]>�H�>���>ο^?m�?3)J?�!�>��;
�Ž�����ԡ�U';��<�䑼�Y=�$�;�<�M��Xz�<����M���Q����z =8g<�t�>����>e�i>(����>���}�_���Z>��K�m&��R x�;�$���=�`>���>�Oe>
W���=j��>���>�7�1?��?�-�>E�1�Ԗe�/�ؾ�F+���>��=?�e>R�����m�z���=��u?��Q?���^���b?��]?�S�=�
�þ��b��v�j�O?��
?��G�^߳>��~?<�q?��>��e�15n�p��Gb���j����=Um�>^W��d�qE�>{�7?_F�>��b>��=�۾M�w�\v���?��?���?���?h'*>`�n��2�������:#^?���>w����"?p��N]о�W��l1�����z"���~��m����N���E&�#��.3ؽ�8�=��?��r?6q?��_?@� �]�c��^��	��oV����t���E���D�X�C��an�|[� ���������J=����7��d�?��N?/2l�q�>�����9�qǩ��Q>�^㾢-t����=5{���P>%I�b���(������?���>d'>�=?�[����5� �¾G=��#z�IS>��g>�8�>Bi�>�,1���[������6��*�ʽi@߻�T�>s6?v�~?��?nm�R2F��f<�zVA�cN�=g���
"�)�H�d��>px:�(��=:t�Y��� ���=�ʹ�<O���a>V��>�p&?���> /?�
?�L�y��z#���7
�����ǆ�>5yu?k��>�S�>b����3F�p_�>
�\?H�?]?���;�A�,t;�[Xž���>�5?�&�>p�=?�<QH���t��K�S��$���E?�;���9T��.�>�?J?h�˼��<��[>k�&�0�����d菾�">Nv?�J8��wN>ʻ���|E�Q�����轕�(?�m?� ����*��N>_� ?� �>��>���?�!�>l"��\�0<��?$B\?�^H?]@?���>|4=�ڭ���ƽ��)��>'=Cm�>V*U>�{y=���=+����]�����N=Э�=�ِ�����
�!<����*2<D��<�4>�{߿�WW�Z���Xt�ڇܾ�;�ʒ���rĽAY��;�{�C,þ�����O��j���Z瘽�3��%�~�j���u[w��j�?Jj�?���"뾇9��	[������>���M9�������C$�u��z
��C�GY<�N8f��6`�9�8��&?����wǿd���6eپ�S ?ؿ?�Ox?�����!� �8�}a%>�o =2������-��'Ͽ���Fa?�p�>�Q����^6�>�"�>��X>��r>_~��}����<�a?w�-?{��>�m��Pɿ���#��<�x�?Z�@�@?#'�v����;=xI�>�?��r>r���-�zO��~��>�j�?�؉?1�=�W��ؕ�`@e?c��<'4�Y>��x�=t��=�;�<t���/>5;�>h��bO/�y9�s!>��>dp�ɭQ���z����=�m>����L��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�󉤻{���&V�}��=[��>c�>,������O��I��U��=���4�Ϳ���	��7�<��(�"Xս���w���R��u��9m�NL�%>`�=��8>`Ez>�:>�>g�T?,?���>�j'<O��� �d�)n���>m1��`䑾��������ؾ$|��!^�e�Z�%��#�ݳþ�=���=�3R�򗐿�� �o�b�:�F���.?#�$>V�ʾ��M�
7.<�yʾ����0'������F#̾��1��n�]˟?��A?G���6�V�����[��f���W?CH�$�� ᬾ��=�α��s=�>���=*��%3��{S�f�?	G"?�O���ᾓ-�=<�7�Z�>[�@?�#%?З�=zR?=�'?0b;���������>;�	?���>;��<\�l�vʽ/��>�y'?Y��8 :�;>��ɾ0���Y���O_o�EaǾ���=���>"���X�%w�iV��/ȼ=��A?|��=��O���.�S��ƣ�>��;O��?8�v>Ք�>AsL?R�3?�o��m���G�������I>��l?�gZ?��\>����_����U>�� ?9Ih?��f>�v�y�`�2�-m������o>�?�%J?�\d>����H��?���%�N?�)]?6�;��˞��o)�+�ɹ�9�>��]>�/?��0�#�>^p?���=�����¿9�A���?�@:��?] �<���R��=�]?'k�>���s��~������s��=���>C��o}r����f%ݼ�0�>	Z}?Fj&?s��zG.�>�h��O�?Ip�?�ξÐ;���	�x��쾶�=�F��:��6�(������XKپ���0V�`����>I@��.D�>횼����������u���\��~��A?8��>�x��Pľ��D��nY��]6���3�$V���>kL>O�I�E�B�tw�*E�V@�=�8�>%��'8>?T��V޾Q�H���=:��>O��>�<>�xg��9��?�Ӿ��Ͽ�ě��r���M?%�?r �?�5
?��@�*���8��l7���jN?3�`?B�K?��=�MF�Ə��r�_?�7��@n�\�(����@��>�!K?l��>�g_�\r1>�~�=f��>�S,>0�V��?��`<��hV�?��?O�ܾ��?�#�??��>�b$�!���ҳ�����^D>3u?C�0>� -�`?�R�m�:���72?[?Q��
�&�[�_?!�a�E�p���-���ƽ�ۡ>��0�
f\��M������Xe����@y����?G^�?`�?޵�� #�e6%?�>W����8Ǿy�<���>�(�>*N>�H_���u>����:��h	>���?�~�?Hj?���������U>�}?�A�>���?���=?�>a��=^~���A��� >8�=-G�l�?��L?�(�>���=�9��/�!�E� _Q�Y�UkC�$Q�>%�a?�"M?�h>���H�G� q!�aqսpq4�1��Q7D�Z�(���׽�?6>�k;>>T�C�s�о�� ?e���Ͽ)ś�[���A u?��>��>�����ƾ��R�
mn?�">5�jc�������/��ʦ?*��?�?��a���)�:�	�>���>�.���=�ZU���=��5?�@=�����7n�z?P�?yk@���?qq���i?_����bς��]羺r��tX�=�??K��;_^>ޒ�>�PE>*�}������+l����>��?Q��?F��>|e?��\���2��0=�v�>EQ?��>k��='�޾q>e�
?��Ԏ�ȸ��uT?�H@��@�u`?f���D�ݿ�d��T_���u��+>��8�;_=�
�4�&>�ـ� ͽfR��M,>t��>G;�>kFo>.(>��>n��=�܊��2.�fD������g:�"�@��4�ϱ��������vX�,��t����	��Ac������?I�r�P���^;��#>f�>?L=?U;s?��.?�v���g�>��ʾ˹��B���O�>�����Z?���?���?�b>Y��j����w��%⽾3 ˾���>xȟ=��>�Q�>�U��}
��t�>���= a>An�>� >�y<��=�͛=��%>m�>Dr�>"�<>�Z>բ��G����h�Փw��ǽa��?ܭ����J�.���ύ��@��|F�=Y�.?�,>f���IJпj��zH?T����\�N,�ҁ>�0?aW?a?>� ���xT��t>�����k���>n �#�l��)���Q>_?�g>ͧu>6r3�i#8�H�P�����7�}>�.6?+��W�9�`�u���H��ݾ�GN>%�>sY=�oO�����4��Ui��N{=Y::?�t?���������u�	8���Q>� \>��=Ō�=��L>k�c�pǽ,-H�Y!0=U�=��^>�
? Є>���<e�}>�~���@��:��>�@>z�5>�m3?I�8?�K�)傽E�6��'���8>���>Vb�>[�5=�C�e�>��?���>�I�K��[*&�N]��#��>�;ս��� ���?�=�ض���>$���n�����-�<ϖ~?��;䈿2뾕_���mD?�+?�=F<�"�z���4K����?P�@Dl�?��	���V�m�?�@�?�
�����=|�>U׫>ξ|�L���?��Ž�Ȣ���	�#(#�S�?X�?��/�.ʋ�6l�g9>]%?�Ӿg?�>�
���@���$��2J=�b>sĵ>��*?�������팾�5?]B?����Ѭ�؄ѿ ���R�>�+�?���?)P�䠟� �%��n�>j�?�cN?�?m>�Ҿ#&��s'>�hA?J>?/G�>bx+�����??ǵ?��?�M>��?�u?���>ʅ���53�5/���ݍ�.=�=�p=��>y�=�M��ǿG�/^��8��\xj�Y=�/b>��'=�6�>=������ɖ�=i��:|��Vp����>K�k>&(P>�>�6?�z�>pw�>C
=]죽����ύ��kH?E�?T����UD������E�;^�M=c/?�?L�߽3yؾ݂>�ER?_�?Ұn?�h�>hC�"U��ݯǿN���!�<�S�=1��>խ?c�=�3>����$ba��9�>���>�c��!���M}�$�����>B�1?�3?e�=)� ?դ#?'*s>.ߵ>.cH��ђ�I�C���>B	�>n?��{?N�?��44��n��$���[���G>��w?T?�v�>R���rd��ƍ�'/G�K�x�(��?��e?���%o?7�?x�@?j\A?�{Y>+��1۾�����>F�!?��qA��D%����?R�?�A�> ����ڽ�-��������?�z\?�/&?l3�l{a�z�ľ(��<(����ػ*�;�����>{>H���l�=�>9��=+m�q�8��+n<=���>�%�=�3�l���O?�?�9�P��-��!|?��45��@=���>�B���O?��o���E�zி�u���ʐ��R�?���?�%�?�,��z�j��B1?���?�h?{l�>,��I׾�G꾚f	��(2�y)�O�>�>Tv�=U��:^��#��<B����M����|Z�>u��>j�?Y�?2;g>�C>�G��+�#�ҹ�a�G�V��D�����h�$�s�ƾ�^^�4��+ľH��QD�>j��_�>c�?)S>I�T>��>�������>ʝ�>=�D>Կ�>z�w>=N>�w=>�~U�="���Q?����)���1��&�D?Pd?���>;���!=������9?Bܑ?
,�?��m>z�i�G�'��p?�c?s~��x?��==�Ѷ�ǆ<k������H��^���r�>h�ݽm&8�ZK�C�e��O?<?��V�>fξ�GսB\��r=V=� �?K�/?�1�=zP��k��]\���J����-	���ș�S"���s����ݬ��f���yN(��x�<�(?l�?�����*ɾ�av�9���g>7�>���>϶>�/6>7���3���Q�]���y��1�>�wz?u��>XF?�$?5�9?�a?�c�>�->�Ծ��>���b$>���>�< ?[�E?�m?-Q�>f[	?9`>��a<����!⾓�?y�7?\�(?�?6��>d����N��bE�߿��A���C�<!ƽ=�t�=�� �=����q=`�p>�?��-��gP���ѾX�>BIr?�?� �>�)���~��8=�-;�?�O?�^�����>����>p��?�������6 >��>k�=���"ʝ>��<SX��~�=��0�k�>R!>��=��%�v�=Ί4>��Q�M)q<���>��%?��0>n�Q=��K��e�24	��Q$>)Y�>7;�=ȑ>nkR���������1W��U�>`}�?]Z�?��ͼǖ�=�$�=-󻾗;��B��?ۈ�#��<T�	?�L5?�P?zT�?]�@?[�?��#>(9Ѿ�����y���y���?�,?�j�>��;��?Ψ���4��?�>PBZ�����"��ϾM$����">%1��{������_A��*n�F��;���%0�?�P�?��a�/4�c�ﾸq���襾Tc??��>p�>h��>e.�O�a�60��%
>�^�>$<Q?͠�>�?O?"~{?�U\?}�P>s8��ᬿ�̙�i���N!>-Z>?.&�??�Xx?�S�>p>90�������G#�������R=�+[>�̑>+��>��>p��==�ѽ����?��_�=e�c>k��>�ɥ>���>\Ep>&��<f�$?p�>9�¾��4��L���n�@��[?\l�?D�_?e�<S?���Ip��y���>���?��?�1?BC�ήn>��F�e��#����1m>���>���>3sv>D���J�=��
?%l�>ii�����u�A���=^?�~N?�~޼��ÿ��q�?L`�<y�����<s����pt�����yZ�Y�=�m�����
p����V��曾ϑ��F��$!����w�RK�>�eo=�@�=.��=@�<X�*�h�	=C�=܂<��"=,U���<	�,��B
��<����_��|o<�F`=@k!��ʾ
}?��H?�i+?59D?,�|>�
>�?�K�>+⎽B?�T>9L�Ք��H�9�]5��ft����׾�վ��c������>6`C�դ>�o4>z�=��<l��=C�n=�ߓ=q`s�T�=u�=�=��=B��=��>�>q3w?=���k���N6Q��3��:?�)�>"��=<ƾc@?<�>>�.������c��%?���?�U�?��?'xi�8Z�>����NĎ�gq�==ɜ�]2>պ�=D�2����>$�J>ł�9H��S}���3�?��@��??#⋿âϿ�c/>��7>;*>?�H�AN9���=�`i��J)~���?�>��Xľ� �>�T>h��q0վ��d�7�V>CF�=P2��cP���=���kP<��[<T�|>�XA>�t=�����l/>ι�=�q>��i>��Ҽ��⼕��W�=�U=��d>�->I2�>�>�>�g!?��<?&��>�		�{<�( ž��>��>�o�>�s����1=U�>�?�Z?�3?6a�>�	�=A��>���>^���j́��W#�4!��	�<ѐv?�Џ?5k)?X>c޼8�2�VNY�[P���*?�7?�q�>D�@=�n����Y �/���\e��<���|�a�� �<�rj�$����D�=X)�>�~�>˖�>L[�>�E>a��=�L�=!:�>��>hJ���/�=K�+�
&y>��,=���_b��<�n��x�=b_j�rO較��<�ER�i}�<3�g>��p<�X�=�#�>%a>P8�>���=�����,>�K���6K�5�=������@�tc��{�AO.���8�A>mX>+ju�(����?�^>�{G>7��?�0t?qF>X��̜ؾ���� t��%\�qɸ=�&>l�9�b;�]`��mL��6ξi6�>��>A$�>tȎ>!5�_	C�O B=��쾍,��V�>ܛ��杽���\�f�����W؞�u�p�>o1�P<?�
�=��?Wm>?"�?S��>a���9��s�>���I"�)��-oy������ ?��!?���>a���p�A�+̾����Ʒ>��I�n�O�}����0�7��v�����>D��]�о63��a��'񏿙bB�`�q����>�O?��?�a��O��BRO�C���#��K�?+tg?�)�>^Y?/M?q���u�֝����=C�n?~��?�2�?2�
>���=L���C�>�J?���?>x�? Z?�kd��V�>I��z��=��%$>�K>���=9?b=�,�>%�?�w?�ٜ�������.��s����G�/5�=�ߢ>Ԧ>�ժ>�'> �<*�=Y�%>��>iH�>� �>�!�>.qe>ol��:E��Y8?[�%>ZT�>K�-?f@K>(t�<�R߽k��;����<�Z�(������n�F�����S�D�V=&��g�>��Ŀ�n�?�C><Z⾽^ ?مپ,瞽�J%>o�:>����>J�7>��v>5F�>�j�>�75>�>y�	>C�d�=���ƽ.�#5��� ��G��('>U��Pǈ�,A
�fP'��;5�Ϗ˾���޲��l#��=�+����=u�?rg>���گb�$���;?D�>k!!?��<�#�=
��=��)?� �>	�D������c��Ŵ|?��@VLc>T�>K�W?��?B�1�E3�zqZ��u�� A���d���`��֍�����Ӗ
�~d��m�_?��x?�aA?�[�<�Ez>���?��%����)��>0E/�n;��<=͈�>ڕ��M�`�W�Ӿ��þ&���&F>B�o?q �?tM?ZZV��	S�"�*>7?�d0?�w?Kz6?��/?^)��t?�q�=��>��?uc4?�q2?\Q? X>+��=%ܡ�-Rh=o<��h���o�ͽu(���ZI��PQ=Һ�=�D<�<�Z+=Z�,=P����{ ��֩��(�<>�f=��=�x�=�D�>��J?��>���=?n2?JE��,D��a���`)?���=D����(�F��Jv��V�=�e?D�?yFX?�p>��A��d���<>1�A>�4�=��[>�1�>(sa�k�޽��>�>d��=��N=6����X|��� �YA��h��)@>��>�'�>��o��F>Oט�^~��j�>�-�:3Ⱦ8�x��<@��;��@c����>.mS?�� ?L��=�������_��.?&k,?�G?�ȃ?3��=%�꾒�7��H�r�>��>K/=����ݞ�� ��k�6���<u�> ��<t���b�>��Ć�أc�لS�(��+M=o;���=���8�վv�p�@�>��=*�� o�����ӯ��E?�·='Ϣ�;V5����ϻ>��>��>ӽ%�y����O��6�<��>�2�>3�<���&M�S��s>�X7?e�]?���?o��n�lt�;�¾�	s�4�p��!�>�?�>�5E?�Y�>)�Z�)�澎�9��ol���#��X�>��
?ҿ*�S�7������$���ݾ2�u>���>MW>ǵ�>��>ig@?�E?��J?��?�R>e�b�_�
�ņ#?n��?6C=cb���@�w�6��F����>�)?�=�v��>�	?�?Է&?��M?�?(>0^���j>���>SЋ>T`V��
��P`q>KA?ӻ�>��W?=�?�E>�L0�����2����f�=p�;>�\6?��"?ۼ?ן�>L��>����=�a�>Lg?��?�<g?{/�=��>��e>��>+�2=a��>��>��?,gR?B'u?}ZA?~��>1m�<�7��ؽ~HF��n��tQb;�!�4{/=t
n�e����#�|E�;�o)�ot���A:�w߼^�L��8�����:�A�>�hv>,1����)>-���q���=fN>�pz;I7��������?���=_+z>S4�>��>�- �窰=���><��>~���S%?"  ?��?6�'
`�D�ƾ�U\��q�>��@?�W�=��k�������t���g=�#l?�_?�~E�V�����[?��[?�)ѾU�%�h�̾ʲ���̾T�A?3?��J��g�>4{�?��?o$
?	v���o���� �f���o��@�=)��>���̮^�9H�>�g$?>��>�|x>� �=�=о��u�F캾;�?���?�?��?K >�El��t߿$>�������[?�9�>�X����?�N��˾�	���ڔ�s�ྂ窾�Ω��g��^H��uN*��䃾�tϽ���=n%?�0s?*�o?�L^?�<��oS`��^���~�\IT�;�L��	I��G��B���m�ה�Y�򾂁��˙V=�hf�UO���?H�.?��S�g�?�pk�vL��yپ�_>�W���:�?>�
.�5��3�\����.:��a�4'?Vs�>��>��M?��S���$���.��|G�#yǾ�Hb>p
�>�s�>MF�>w�ͼ_eD�~��.hξ=����D���j>�8P?5�l?<��?&�|�b�
���[�/'���
>柾��y�>3��>m�?���S=���Q���q��u��H�������>�r�Ն�>���>k��>Y��?��?�V)�낾�@`�%�!����o:�=5�+?,�>��>̻<�^.־�=�>=Z?��?���>}�ƾ����h�}��9d�>���>a�?�d>�t�H~f��D��^����83��*>��R?au�����yj�>��0?��=��}=��W>�]b<p�%�D��T0�93=>�?2�1>f�>��羙&�ָ~�@σ���+?RZ$?�Ⱦ� �kX�>*��>蔇>È9>�Xj?�r�>��l�9��.�y>'�a?pGp?��M?
�>��l�^���Yh<���㠽��>�b>1��=��^H��e\����Q���=��2=v����ڽ��e=�g<�37=\Ĝ<f._>y�ۿݾK�sپ����\���
��ވ��*������r*��������'[w�*��-�JRW��#c��ዾe8j��U�?���?'�� .��e\������ ���ȼ>4Sp�.oz�� ��X���ߗ�)w�����Ѡ!�wO�!h��	e�E�'?ẑ�ͽǿᰡ��:ܾF! ?�A ?+�y?��D�"���8��� >�E�<�*����뾮����οJ�����^?���>��.�����>ť�>��X>�Hq>����螾71�<��?S�-?���>Ŏr�,�ɿ^������<���?(�@W<=?��0�1Ͼ���=;�>�?XJ>,G)�!���4w�>a.�?��?D��=2�X������V?%����7�ـ����=�B�=�f�=o����|>*�>�?��{*�&�ƽF7>ϸ�>3P;��V�Ak���$;�DJ>�D�u,1�v�?�)?��Xl��2�ʷN���>h�F?�0�>O�=�-?��D�4Yп��i���Y?���?��?Ӎ?$(���>��羇�@?��7?匇>p'�gO���?��ƅ=���=����+pO����=�H�>4t�=�w)�AW!���4����;�t�<4��X-ʿ�A����夸��'��(�Ľ3�|�@q>�dI��y���o� ���׊Լ]��=FaF>�C`>�=�>ܬ]?��h?:о>a�>(߸�� �-����y���/�Z��wq"��;߾t߾n�����پ�b �-��qPE���9��|�=�'P�C���X���b���F���.?��%>�ʾG�N��	K;3�Ⱦ�����ɞ��<���Ǿ{/���o����?��@?sÄ���T�qX��8,��h��5eU?��S� ��3��:��=�Ӽ�#=�ڠ>9v�=���^�2��P��N+?�a&?��׾�!��%�>�Ef�]�<�n?�w�>�|Z���Z>U��>j�d������0�>�|>B��>*�>���=�ʾ�Z���a"?�.?3h���d����>JHپ."X��ƨ<�>��W��ez=�!�=�%j�l�����[�� $�=�V?�A�>Y)����q���@U�J�?=pux?��?���>B�k?&�B?���<�}����S�rQ�=s=J�W?��h?�
>���о�(����5?�Ce?��M>G�g�E`�f�.�!�NP?��n?�?}Ӝ��=}������uV6?�pm?87S��Ƣ����J�Խ�{�>Qy�>z�>2#A����>�2?���𴓿ۺ¿y-��7�?g�@̠�?��޽{<r7=��>���>	���*������^ž�<�<4/?_֧�m�x�y�@�s�FqF?���?&��>8:��k����q	>Ȣ�� ˴?���?8�ھ&vg>
W�����!��!��=�>���>���=2O���R��h�͓3��=��H��>F��>6s@��H=?��žd濶ếh��|�=ҽ8� ?��o>�Ţ�o����>T��M��B���0������^�>·>����젾W�l��G7�Y{Q�-� ?�}��K�>�[��+ѹ�dR���ҿ<w��>���>ˈ�>s1h�c����ܕ?���ږ̿��;���ID?���?��?=�%?��b=뵀�g�n�ϼ���D:?�u?��a?��b<�YZ����w�j?`���R`�Ɍ4�cHE�JU>b$3?W?�>��-�ٵ|=t>��>�i>�#/��Ŀٶ��������?K��?�n꾊��>��?�u+?�j��6��TZ����*�K?$�>A?<2>����!�n1=��Ғ��
?�|0??y�-���_?�Ha��#q��&.�&࿽t#�>��0��_]�@��+��Tme������|�ն�?=�?hB�?K�p%#��%?\N�>9o��M"ƾ� �<Z�>���>7BO>��[�"�u>����9�l�>s&�?��?��?!���"����
>�~?�>r.�?�<
>(��>�(�=���������7>w2>3o�t�?|�O?���>-�=�A��3�K�q�R�.����D��D�>)Y\?
�D?""�>�ýN�I�Ph�����{+ �n���[D�������#+>�5@>��>�>�?tƾ��?9m���ؿ�l��m'��34?͜�> ?f��͖t�=��9_?�b�>�>�B*��E$���%����?D�?	?<�׾!�ͼ�>{�>�a�>x�Խ�۟�+�����7>}�B?j��%B��N�o���>W �?��@�֮?�i�	��>D�����8$���쎾���=�
��6?Kz��s=>;z�>��P>,��x���Wo�Z��>Z��?��?*!�>J��?D^6��f��=d=&(4?�d�?�?�����l�=��?�2¾^�b�7���Y?�|
@�@(R?�� �ӿ
l���������9�=��=! O>�ꁽ�Q�=�/=���A=�8k=Ƙ>�>��V>��[>%�2>�>�F'>�����'����ӥ��M�E��{����It�� o��;	�q�r�v�þ��̽.´�Ϗ�s�c���=�Ҭ����$>��b?�@?�il?�"�>������>���v�
>���Fo=��R>�`V?'i?ҙ?��;�|��w�7�t��C��	�U�Ε>)�>���>e��>X�>?8u=:4>%*5>Wp>��,�����4gϽh{=��]>��> k�>
�>@�<>Si>8}������-h�tGy�2�ͽ(��?q=��p`J��╿�ɍ�ԍ��&m�=
].?=;>�㑿xп���kH??x���H��N)��>2�0?3W?=�>���^�O��
>0-	�K�l�q�>hA��f�i�;�)��N>��?�cc>Ҭ�>-5(��;�Wz4�[D��Y��=F6?�!����}���u�FCH��l׾�EY>��>�	<�������N܀���o��]V=�u4?��>}�ܽ�ｾ����X��~?U>TF>zM�<�+>I�_>]��uLC���j��k�<;�>��=���>x�7>�m->W�>2��jK���?�>�5<>&r>��D?1?[����� ������A��]>���>r3�>!{
>�׃� E=F�>0�&>A����� ��މ��g��
8>��A<
������F.>�2����=㷆=,0�r�=�F��=�~?���#䈿��e���lD?:+?� �=��F<��"�D ���H��8�?l�@m�?��	�עV�7�?�@�?S����=.}�> ׫>�ξ��L�α?��Ž8Ǣ�Ɣ	�=)#�hS�?��?M�/�eʋ�Jl��6>	_%?!�Ӿ�g�>�x�LZ�����z�u�	�#=���>�8H?\V��P�O��>��v
?�?�^�ȩ����ȿ�{v�A��>=�?���?%�m��A��@�6��>"��?*gY?Roi>h۾�`Z����>G�@?iR?��>�9�!�'���?�޶?���?�\>�?T|?
W�>���i�.��E���P���yA>�wT��ɤ>ԝu>�ߓ�bR1��1��pa��!�v��"���>�Z=�>h��鲾��=뉴�)Ӝ�ȗٻI�>�>��>t�v>��?���>\�>��\=e`���(��V�����E?�S�?B��Ne���=�-�>;b����>�}:?�Yw�v���l4�>]�D?��?�J^?9K�>^���6���]������]B<���=g�?e��>I(T<�`>doʾS�i�>3��>Й.:��.�B�)3�=[�>t�?���>8,>�?-6 ?�~�>rt�>�	J�W���#?��۩>�T�>��?�H�?k(?)����/����ޟ���^��T@>�w?�y?z؛>S�������L�G����a���s?ec?"@�m�	?�j�?��C?tJE?5�h>k��6�ھ��ʽ�Jn>�.?���P����Am>�s�>���>��~>�}@��y!>l�3�s�@��E1�SD?��?�\?������X�����	�K�s=���IF�=��>�|��=��<��<�|�=�o���`>�g���l8��r�<5DH>�8>3��x�[��t0<rW&?�i�;��ؽȽ�>{4����$��e�>��=TS�ۅ|?k콯�n��˗�]ܫ�l{y���y?1�?Q��?��˽�h]��?k�?�?�u�>JU����#�gĺ��s��g}��0¾_:>Mc�>�Vb=޾W4��b����1��w	��པ��>s��>A�?K�>7��>w5�>a�+��J��;Ͼ���J�8��꾓8�\2�8�!�·���h��5ڻ�7���������>M�Q�u�>�Y�>���>��>�Ҁ>5��=3_�>��\>�w>�^�>_�>���=  ==nƑ�%����FR?�����'���������2B?�md?�&�>1i���������?҇�?r�?�v>1�h��1+��c?{<�>>��Io
?�@:=�"�<��<M������G�����S��>�$׽G:�eM��{f��e
?I+?I���P�̾׽���Rkk=�7�?��(?5�)�Z�Q�s�o�GsW���R�O��`h�w[��]�$���p�5珿+`��x���n(��W.=��*?��?ix�[���׬���j�p?��e>u��>�U�>I̽>��G>�*
��1���]�"W'�։����>�<{?��>�J?��7?�M?�K?���>��>�a���K�>³źKD�>���>DZ6?w�,?Ob1?��?u)?�Z>O������(־��?V�?�Z?�h?)1 ?��������ټAӥ���r�f-f��WN=Db<Z�ݽee�O��=�vT>:E?:F�qy8��o��P�j>�j7?e<�>���>���Z��Y��<���>o�
?�S�>-����Yr��h���>^��?�c���=~S)>=��=a���>yۺ���=i�����==�]y>���"<E�=��=p��� ���;Į�;�_�<=�?�?}�>��>PS�Ἶ�P�Nܽ���>-�>�t�=W��X��׮��ob�޴n>���??uA=�^=�<V=D�����%��`D�Ov��b��h�>*~7?�m`?s�?&[.?.�?�����{������tƃ�&d���?,?�i�>@��	�ʾu稿�e3���?6^?:a�E���9)�Ȉ¾��Խd�>AP/��#~����kD�p��K��1ڙ����?���?��A�$�6�ρ����8U���C?>�>4z�>Q �>@�)�h�g�6�j:;>5��>~�Q?[&�>��L?X��?��m?���=��.�����r�V�=��=o�=?�ڇ?��?�B}?���>Uљ<j难�5��f�ؾ�U��τ�r͒�\*�;�|>�t�>���>��>���<5�������9�>U�h>�Y�>Dy�>YZ�>��V>���K�5?�e�>���<�����M���k�=��?1:{?_)#?�D���]�q,�#˾Oխ>�M�?gv�?��'?�`+�Ip>�稽��˾�~�=}͡>���>$?�݊�Ȍc=��>:��>mZ>.��`&��̾��>�0?Q?�_>1ݿ�����笾 ��U�?�ӽe@�j5�����:YK= ��8���	8%�K)���J����d�8𘾨.?,�>="�=w�m<٪E=�d��M��gF>���=�Z	=Fcּ���=���;]{��։��>I���_��&��<C��=�5��2�g?� H?� ?�7?B�>d��=��u����=�䊽�?�HU>��:p^Ͼ 炾����@���O���Ҿ�fe��L����D>��r.�=�,�=�+>��(>Q��=L��=2�;�ٜ���@�O�>)��=ו�=�06>3�>�>"a?��]�֥���V����>�KB?�u;>kB��i��Z?,�C�n�b��b��\����|?���?���?�?�Ò��6�>���o=�[=..����UR�=IQJ�Ep�>(�U>;��:➿Ki����?���?�a?�[���\�Ѣ?-�t>�Fg>;o=�ѭ-��j<�`��ua¾��9?w%�k�澻s���Tֽ8}�޼+��SM=��b>�T>�c��	~�~QL�1P�=���=���;n.:>��=8�=W����&L>�w~=+�=��>`��=4��ϯ���;ņ�=��l>Z�<�1B�>�	?�m-?~�??��>m(O�q����?>�Kv=�w>�=(�&>ї>r?��.?�wH?}��>:�=���>П>g�%���`�lT׾B�Ծ#<s>�Ɋ?:�?�-�>����`,W���$�	l�oO��x�?�HO?8?�ª>�������.��&��PV;���P���>ý���g��f��>��:���=}�x>�B�>�X�>�@>w��=Y]=�^�>��>��A�TC�=<���ڒ�@ۢ=4��4����ǻ/W+=���ęr�
��ýE��W>^�*>���=��>-��>�oz>+��>�����틾�w&>�����0-�>4z��'�5��KN�e����P4��o�Έ!>�Ѓ>J�ƽ'���>��d>G��=���?3Uu?�2y=xJ�Y#ᾖ읿��U����뛵=ǻb>R�M��J�Z�o�DU�{Lɾ�v�>L؉>6B�>Eu>'9/���4��=�
Ӿ'�*��?�>�qt�0;���Oo��o��'9��{�i��TV��A?$5���9�=�8q?K=?���?�u�>�G}���վ��>�Vp�P�}=����X��\��"?b�%?�*�>��ﾫ:�8�
��A���d>qP���iE�Gʉ�p"F���R=����>L^ؾG޾��5�N�)J����N�+��� ?ȋh?\l�?�I.<f>��D���	��ŽQ>�?�>2RD?ݎ�>c7?Q�>���=*l<�����L==�W?Yh�?9��?���=���=5g��,�>�2?O��?)j�?�|r?��,����>gT��M->���	>��>ה=衒=��>�)?��?&֚��������������[���<��=.�>	U~>|�^>�#�=�Q=�8�=Ȍg>I��>��>1/f>�Ş>H�>�����F!�a�E?�N>��>h
 ?3�>�Ъ=��y���8;�]>=��=���=d��<��`�E�d�.N����%I	>F��>+Y̿ꦑ?f�F>����cQ*?�߾�������S$뽹���6?��c>��>��>�>��<�T>��l>ipӾ4>���ZZ!��,C�)�R���ѾC�z>(����G&����C���I��s��8k��
j��(���+=�s׿<ID�?ab��x�k�A�)�k���q�?�;�>�6?ό��󈽊>�><��>aD��P���Oƍ��_�|�?���?,�`>�̔>�+L?�?C�'�����c�vze��q;��<]�~�i��i���}�y���&�佣X?�q?�>?���|�r>e[{?��)��Đ�*f�>�;�.-����=&��>�ꌾ�̇�����3/��A�P4>��s?	'�?�?�W=�"�c���'>T�:?�2?%/r?Rf0?�:?3B�t!#?'�*>HI?�-?�45?��-?#�?R)>�k�=�ml��cN==鑽����佅�ս�_ ��6=�-�=���;�U�;��=�<̕��7y�����;�O��AO�<��B=6��=k��=#L�>]]?��>p��>��3?���z.�.��T(?�!4=�G��!����j������g>i�g?�?�?;;W?r#^>�"O�^�?�!<0>���>�<�=�R>��>�A��7���=�w>�j>���=zu�����E
	�6!��G��<P>E�>R��>�uK���n�����fAD=�2	���
�l��R��}�>��3��	��3Ed>��P?�!?��=?J�����=�h�_M3>�2�?,�>��>�K>���C�;�RG��֙�5f0>փ?>�R.��Q��-������_��=�?U1���U��a�e>c�
������i�5-K��z�k`�=�����= ��
վ�)��F�=�t>	���:��8R��{���G?Y߅=V�L�䱹�P>�	�>
�>����H��A�=F���=ݟ�>$C>�*,���lG��R��K�>�H?�`i?�m�?�7����n�(�7��?��[��Ň�t?�0�>;C?��a>%��=	ξߍ �m���/���>���>���]:��B�����+��h>3�?p�=1�>`AF?�?n0b?i�*?�#?ӆ�>���%ػ�@�?��?j%j=�)!���:�q6���<����>E*?���)]>e��>�8?y,?�$L?�7?� 	>���1�e��>C:�>zM�ʑ��k�\>�Q4?j1�>�PX?C��?ռ0>.�>�1�����*+>�4$>ɪ3?qR?qL?M�~>�&?�㮾%����>�bU?��?�,n?�<�=�<�>9�+>] +?��>g�=�>�>�M0?@g@?�@V?�,?SR>Y!=���(dL�O(�����=y��=��=�|�>�Ȥ=;0���_>���=�[5>��zH	�U^��x_���m=9v�=s��>�t>a핾��,>��¾$ԉ�h;>m�U��陾=���Kh;�		�=%9}>HS? ԕ>}x �b}�=���>;��>�����'?.M?��?ua�:�2b�9Iپ�K�^��>��B?���=}�m�����ùs��oo=4�m?�~]?t�Z��t���b?I^?��"<�3�ž��c�ך�C�N?dw?=�H���>�^?[Mr?>B�>�)e��n�*K��$�b�_j����=���>a�zd�S+�>�7?LF�>.yc>���=�
۾��w�*/���L?��?a�?#֊?	�*>��n��C��?۾a����\?�B�>%����5)?	WH=��t�|�BUw�h{޾;���J���V���>�����-�n��m��|b�=d,?}i?�Mt?؎[?�����f�2_�dw�dOT�g������>�`73���G��+k��$�o�c
��_��=�H�m@��;�?�$9?*�N�%C?��0�ZQ�'_���3]>S�|�Q=B���p>�d��m�����卾^�i�a
����?�>���>�)5?;z��-���1?��ľ�*Q>ڂ�>�K�>��>�8��j5��ӂ����¨�>�鼤k$>ȍb?_#x?�r�?�|Ͼ�"��uu��};�4�[>lɃ��=�Y2>�)?5�
�
a��4iZ��p�Gώ����u[������5�=��>OF?dM�>"S�?�I?�Eо�n)�*�Z����ӽ���>�xD?�>`w�>u�ʼ��)�	��>��`?[	?z��>������ ���u�-ك��G�>�Θ>��>#>��b=Ks�=;��̿��p$G�|�;�]?򦾊s�r��>�:9?��0=[�Ƚ��=�==at�_���k]轍k�>�q
?��q>|>�F	�e:�;���5��^6?DE2?�����
&����>2��>I�?�f�>�sg?Ա>� �+�³>�j\??0M?l;?N$�> ͋=����1�<-GK�h���l�>OZV>���=�f�=Q��a<��(�����)>I�d=`jm��s��W�=�=�=�ڣ=ԾL>�bq< aۿOK��Lپ�P�����q
�A4��孽2����X�5浾���rFx�ҟ�+�-���U��/b� ~��
ym���?��?⒓� ;����������% ���:�>�fo��>��Ǭ��Z�qK��G�ݾ\���a�!�cP�,�h��d�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >WC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾s1�<��?7�-?��>Ǝr�1�ɿc���z¤<���?0�@�D?r�)���;��=�?�> �?ʁQ>�(;�- �U�+�>���?'S�?δ.=�M�$U7��Pc?�<�cD��/ں�=�<�=$b=��]>ۊ�>ڱ��8�쎷�4�O> ׄ>	A;�B�2���Z�e;�zL>(��Ժm���?�{U�Ԗ^�\10�Qj���>��P?�w�>J݁<��8?5�*�S���pVa�p%Z?'��?�$�?<�'?���&�>^�t,Y?��0?7�P>�G��~��A�=��нc ?;���A�l�a��<�#�>�q�=4^k�37	���.����~>���ixƿ��$�q��.�=���P[c�-彦����JW�4󟾏n��齴�a=�W�=.R>��>�`X>��W>��V?��k?rݿ>ſ>�罯�����;�a��N3���;�<���8����뾄3߾ţ	�F;������ɾ��7�./�=��F�哒�0���
W�bj^��U9?�[>�m���@���4=��ɾ����i�#���Q�I�q�n���?h�G?%IE�if�~��0���;|߽��^?a]<�����پLz��U�_=��>�d�>�<����Z�2�9���E,?��9??ٶ�4c�,�>X
?��PI>a�9?��>w�;�>R��>�J.����2/�>�O>5�>���>T�0���о��Z��1?wJ?��ƽ�{��hj%>�K.�'M��r���G�<�|����<�f>�L׽l��FV���V��E䊼G'W?Y��>��)��pS�����}==�x?��?y/�>�|k?��B?G�<�^����S�����w=}�W?� i?��>�u��оI����5?�e?��N>Jh�F��?�.��L�<"?��n?�Y?����hs}������l6?�?�#o������l'��>+lF>���>מ"?�4e�f%�=U�?G@j>_P�����d�>�,,�?�P�?g�?��=����l�=~_�>��=��E���j�=P����>�S">�a��B�����4��A:?7�=?e��>��Y�28�.k>��X��q�?|^�?a�jZ9=��о燊���m�`]=&>^I>V�>>
?��%|*�����8�CM ��F�="�>@�k����>���Wֿ�����$����b�8������>
2�>��;F�E�)2,��|�uu�p l�I�J���r>D�=>�M�2�Ӿ�E�>�K��d�� ?�Q�=�r�>peӾ� �zٵ�42>���>��
?�֐>��F��&�����?!��Ah���Ή�&�־��R?�u�?�j9?F)�>.l>�+�HD���h��t�-?Đ?r|?�՚=�*��.x�%�j?�]���S`�$�4��HE�+U>�#3?[>�>�-���|=)>��>�l>�$/�7�Ŀcض�X������?ˈ�?�o����>s��?�s+?�k��7��)Z���*�҅-��=A?�2>f���̶!��1=�bՒ��
?o{0?x���,�>�_?�a���p���-��ƽ��>9y0��b\��/��J��Ce������y���?�\�?��?*w���"��!%?
�>׾���$Ǿ$��<懧>EM�>_/N>��_��pu>�����:�Q�	>���?Ol�?�V?�����樂6e>�}?;7�>5�?D��=H��>���=)^���B� �%>ރ�=�&J��N?�oJ?�]�>`m�=�G9�R�.���E�:�P��F��wD�.w�>�+b?�1K?�qe>C�ǽ��5�#F�)��;4��o
��pF���:��ڽ�`+>"�;>K�>��F��Ӿ�b�>9*#�B�Կ޴���
ཛ�?�[�>�B?���<�=9�yl?�xg>y�)�)<��G
p��N��O�?�*�?@[?<�۾9޽*z�>���>p�>�=d��<�����GW>�� ? ��<�Uk���~��9e>���?�#@y;�?�����=�>���R�����x�CV羮�A��&>��7?N2	�n>���>=�&>h�i�|��M}��ս>A�?."�?���>��d?��k�82��Ly=Y@�>0_?���>��<�����>��>�N[��T\��V?7J@\P	@��Y?��#������a_���򊾥�=��	=1��=���#��<mp�����Lf��=;>���>���=�j>���=�B�=�z>������#�X��@?��QOF���A���J�d�X�̼�Y�r��&�0ܾ������t����	X����HW���<[D�=9T?	�\?Txw??D�>T0����>!�� ��=߆��=$�>kU<?�M?� ?ϙ��N!��ɦl�Oށ��Q��Ha���5�>*}1>$b�>��>�r�>s��<�>"�;>L��>��=�g<xº<>�R=�S>�Z�>��>W�>bD<>ǌ>D̴��0����h�[w��&̽I��?�}��ŬJ��1��,L���֡�=�g.?5�>��}9п�\2H?�	���,��+���>��0?�iW?�a>�-����T�&Z>�����j�	Q>q���Krl��)�Q>_e?Ԏ^>�_x>2���8�,M��J����l>E�7?Ƽ���>��t�߮F��ܾ�ZP>�H�>\�7�Am�V��*|�	qg����=a�9?��?�������,u����%4\>i(Z>���<���=�R>i��$����YE�\=���=��g>���>�7{>jN�<Gu)>�5O�	�;�E��>�3>��{=PoF?��?� ����a0�svڼ�r�>���>L
%>�O[>YF��"�>xS?J~�=G�����O�O��ؠ�>�͗�
��� 3�:S�>񄍼�J)��ׂ��PN��O�ʑ�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�-)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾÞ�>��EZ���"���u���!=�=�>�H?~��I�L���=��r
?��?VZ�@�����ȿ`v���>{4�?�
�?��m�Kl���?����>b��?��Y?d�i>Z[۾y�Y��׌>J�@?��Q?���>����L%��o?���?���?�-N>�H�?z�}?�q�>y7��c1��Ƭ�˔��+>�]㼤a�>l]>�+��Ta3�0݌�����<T{���(���r>�61=.��>���F����=�ͽﹾfr8�>�>��Y>�m�=�w�>Mh
?B��>Yt�>�a=�%���H������]JK??r��E�m��.�<NՕ=��X���?m4?�o�a3Ҿa��>	9[?���?�Z?t�>�j��.���s��>�<(BE>9��>���>2���UK> �վ�iH�맇>�,�>9����۾�Ã��'-�Ϯ�>�� ?��>4Ѥ=�� ?�#?c\k>�n�>��E�0��%�E��"�>���>m-?��~?b%?:l��.53�����*�r�[��DM> y?rK?��>񇏿�f���P��K�D�����?��g?j���?�)�?��??ͧA?�kf>�y�l7ؾ@ծ���>v�7?�о��;���� �*=��I?4 ?�V�>�G��r��=H;�>|�ᾡ:>�� ?1؁?��1?28\�-��޼ʾ3!?=���#�<Z#�x��'܆>Z�>�E1���]<�uX>g��=�^�Խ�� =��x�ީC>���=��7���9=�*?:�M������J�=�Oo�u|?���|>�A>����[?d�;���x�k���������]���?O1�?d��?��Ľ|�f���<?�O�?�?���>[2��7*޾��ݾg�m�b�j���2�=LS�>�*��+澞���%U��Iń�����м+����>��>�?�D�>��&>)��>Xp���l�A�Y����%_��	�n�2��@*���᥾=1��Z��s#����>����Z�>~�?m�I>66>�Ļ>PÕ�en>�Y>��>���>��L>��K><o>�9��`#)�$MR?����^�'���I���~<B?�nd?�5�>&hi�\���_��K}?<~�?�q�?yTv>osh��%+��h?;�>g��6v
?;h:=��̔�<�_��~��@@��t�����>��׽�#:��	M��if��d
?�.?������̾w׽v�ɾo5I<��?�P%?�r(�*�U���w�\�T���R��Kc�uH��Ħ��A �Kbo��������쉄��i)�
B�=*"?�/�?��\������yp�>�D��kz>��>��>~I�>�K>%�
�8�1�/d���,��卾��>h^?�y>�P?�i.?pVM?BE?���=�s�>�pg���?�ڦ��K�>}�>i?aR"?�'?k�? �?�#�>&�G�_:���뾁 ?�<?z��>c��>W��>�x��B�ɽ��<���	��ȫ��`��>� �c
�׽�Ԗ���<T�>�?����8�O�����m>�:7?���>4w�>���#���h�<G��>3�	?$��>�	 �.�p���
���>�)�?1��7=��)>��=[]�>̹���=�������=�Ǜ�C6��<ȇ�=K��=1�˺��S9"�[;��;��<[��>��?ﻊ>l:�>�����.������v�=H|Y>��R>"s>$�پ�ۉ� 8����g���y>|W�?X=�?S�c=!
�=�f�=ݩ���ƽ���k(����<�<?��"?F�T?�!�?p=?��#?� >	��q[���u���ԣ�v�?�$,?)��>6���|ʾ�憎�k3�=�?�??G*a����64)�>�¾ZԽqH>Pb/��~�����D�~
����rv����?~��?��B���6��l辗����^����C?�>�E�>+-�>�)���g��5�V�:>�U�>J
R?�-�>�Y?s�?�r?=����@����F:��?�Y>���=�?tx�?�S�?�[�?d��>��#��h��.� ������e�wEཁb���DW=J�>���>H%�>-�>(��=�LM����C���Ǻ=�>��>E`�>]n�>�u>��:�La<?&ѹ>qǾW��[X��5=��bo���E?�ee?~�?��>���*��M�9F���r?�ۤ?�#�?�?��c���U>J�^��оŊT=b�>]Y ?G��>�r�g���]>s�?&�>4�s���~���u����	?��3?���<5Ŀ5�m��Sn��v����<�y����r��b�� M����=�圾���c��d�R�5n��l����������a�w���>�j�=�� >��="��<����ܶ<;+Y=T��<�|==����f�3�5�E�B<�ch�&�;Y <+�=�<�6ʾ8�{?�8G?�,?1@?�@T>�+%>u�	�f^�>���Sh?B�&>N�[��~��V�4��b�����оi,׾?�g��j��nV>>���M( ><J>'�=�ļ���=��`=C�w=��D��?=<��=���=8��=Ϧ�=��=��6>�1w?���S����3Q�Q'�%�:?&0�>pí=9�ƾ�@?%�>>�0������sP�h1?G��?�M�?�?�hi�.e�>Y��������=}ל��F2>s,�=��2�{�>r�J>�{�&E������)�?��@�??X؋��Ͽ�c/>b�>�;	=��Q���-��7�<�BN��IG��V#?��1�WC徿aW>�>%4 ��n۾&��<p��>��|>D�>�@���=b���ݬ=���<�_>�`)>n�;�� �>I>�<�sm>�<�=yj�;�j=Uw�=,f�<� D=�=��:> �>9�?_9/?�ub?��>�e���о�fþo�>&ح=%�>>Fg=u�B>�x�>��6?�0D?��J?���>B!�=���>�ţ>�+�u�h��;�ɛ��	��<��?[Y�?���>���<�:�����>���ͽ؃?1?��?���>�U����9Y&���.�����/5�g+=�mr��QU�x���Tm�0�㽨�=�p�>���>��><Ty>�9>��N>�>��>�6�<up�=�������<� �����=�����<�vż����v&��+�쏦���;���;�]<��;in�=���>� >[]�>�=6����.>X���@�L����=�0���B�M%d��=~���.��6�]�B>�fX>��D)���?�;Z>��?>z`�?�u?0�>����yվ�H����e�ّS��g�=�<	>p�<� |;��b`���M�2OҾ 7�>��>���>�s>M4-�d3>�@�^=�q�5S4�yq�>�G���8�V?	��Iq�;���2��@�i� �{�C?�2���e�=C�}?4H?L$�?�X�>}♽#jվ��2>�ρ���=q����o��:��z�?�?&?
�>�$�"E�+��YB�X?E>��¾�CI�������R�IO<= ޾���>�V�������"�`8t�f����i����ݵ>}�?6j�?=�T���X�伾HVL>�??�Q?d>�]?�O?m�,>Am�����>
�v?yW�?���?��r>D��= 6����>Է?V-�?H��?8s?�>�I��>a�;f%>ݵ��j	�=iq>6��=���=�g?+
?�n	?�Қ�������I���\��
=9�=x˒>��>*p>}l�=�Co=L�=f�V>~h�>��>r�b>���>;k�>���������:?W�u>� u>� ?BQ[>������;U�_=Xi;�Žû*=y�.��}��������p�ѽ�"�>
�>�����?�	>��پ��"?�禾V��c!B>]1>$�o�Я?��E>�n�>MD�>��>��>��|>K�N>��<��j6��g��w��z>�_�n�ri ���e>$:���2@�]���1�n|�t�ž;�!���u��V��m�<���8>��?^��$z���&[�
�F�-h�>o�`>��B?����K�=���='��>W�;>����?����쒿Ҿ���?��?z�X>\b�>�JM?_�>T/-��&�O�_�\�l�E���6h�;����W��jǾ�����T?fT^?0'?c�m=)��>�)`?�71��'��s�>�ھ4�F�7p����>����.�k�����1���K�#��ZP>��g?�z?�?����5i���'> Z:?�n1?�t?1�1?��;?�~�o�$?n�2>�[?�/?��4?��.?��
?]72>��=���vr$=Mđ������kн�GʽI���3= �}=9�#:��<W�=�	�<�Y�C�ҼwC!;�J��O��<:=���=�<�=(-�>��S?d��>�Ϣ>HV&?#����*��1ؾ~�(?J\��\�Ґ����m����\�=�
c?�{�? Q?��.>ˣ�Rq���=>��>Ql=J�>p��>�	��o��3>�%>��>�9k>�j� yȾ����E_�ۚ�=��6>Q��>�~y>Y��҃>x��rb��Ti>_O�(.��#WI��A��;2�f^��"��>��K?�'?��=�������o_��V!?�7?�M?w
v?�;�=V�ɾ�@;�u�J��#��A�>�<�<5 ������Չ8�j�;�gw>q���<�ͽ}:��H��R���C8�cy��z\7>p�����=!i� ��%ǽuQ�=���>E֨���3�L����ԩ�*�e?q�=�O9�F�m�}-復$=>�Z?��?����2e�Piy��IW�+�E=Oa?"��<7U4>7���L����jF�>d�D?p�`?߅?gpz���k�S�B��-����������?;ۨ>��?�5K>�R�=� ��$�
��8b��$D�P��>�&�>:�ŗC�[q��sb��2%�iψ>i3?L�&>�?�NS?_�?�_^?�I,?zh?�ޕ>�Z��"տ��B'?�?��=�����R�r�9�"G���>�,?��?����>��?�?��$?��R?Ң?��>�A��a^?�Mڕ>�ȏ>x�Y�����*�a>¿I?Q��>��Y?MǄ?�k<>Q�3����;�Ž�/�=�W>�6?��"?��?Z�>���>��+��a>�xy>�K�?{�?aO~?�K
>;��>�)�>�u�=EV�=0C?v�>q?��=?�;y?�dF?��>����q;�MU?��@+� �f�5��!�p=rC=��\���&�}�"��o���v���=
7~=U����[���;�s������>��r>'���Rm0>�Bžp��Ac@>ߖ��5��l����9� G�=f�>��?Pڔ>�$�:�=|û>���>�����'?z7?�Z?��_;�b���ܾ��K�~�>��A?���=�/l��Z��ӽu�XNi=��m?�3^?��W�����h�b?)�]?xk�=��þ��b�p��u�O?y�
?��G���>��~?��q?���>}f��6n����Ab���j��ܶ=�n�>qU��d��<�>�7?+W�>	�b>�%�=?t۾t�w��l��]?��?T��?���?- *>Z�n��2�<��/~���CW?G�>ǀ��4?)����ȾV�������g ;�j���
������k"���6�g�s����s�=.�?[o?��o?��W?����`��yZ�:�����W�?!
�)G�:>��C��4O�j�Ǫ�d(�h��ZB�=R�n��)F��h�?&$?������?2���l�
�۾��>��w����0�=Z����<[��;R<(��t ��{��0?_�>)=�>y]?k�j��,�*27��U���۾�I�=���>�̱>^�>� ����N�Uiҽ�Ҿ�s���2�=�e>��h?�g?gwz?U�z�t���$����D�>1=#C����>�g�>�)>�@�Uƽ�&������h�{�	�?Cx�n4.���}�G4?�w�=���>{��?ɹ?M���]�ľ�j��Q�W���=1�[>���??@-x>�)"�6
�9��>�l?���>3�>�h��c!���{��˽���>���>���>��o>l�,��\��g��Ӄ��T�8���=�h?}��Ţ`��ۅ>L�Q?d�:|8G<�a�>�	v�в!�����'�O>�`?�<�=��;>�jž����{�5��X(?�?������+�F�l>D�?��>���>ن?�]�>�վ���`�?��d?�@?gG?)��> s]<]H�iٽt	�c�C=���>�~U>ob=��=��=�J��.��g=�=z?�`����_��,�5��<@;=9>����yx�����k0���w��{�ƾK������@Ľ����*�P�g��8���'>}�}�@M��>���m��i�?���?����3 =@������_��j�>-��8>@͓�5�.�Z�=o84��Z���!�7�h�����b��S$�> ¦��:̿�����,?��;?���?.�i�%��+[�*`�=�FB�8Bp�����V���:̿�ɾq�G?�>H?Z��oQ���>k9�>�޺=�Y>�ˣ��&��遾v�?�\�>\߁>?膾���26̿[��=#�?�8�?&yA?{�(�t��m'V=���> �	?|�?>�T1�G��ﰾ�J�>�;�?���?U`M=��W���	��}e?<<��F��4ݻ��=�X�=�z=���Q�J>�V�>Y���6A�\Cܽ&�4>�߅>��"�����^��ξ<�z]>�սB��4Մ?*{\��f���/��T��
U>��T?+�>�:�=��,?[7H�_}Ͽ�\��*a?�0�?���?�(?<ۿ��ؚ>��ܾ��M?]D6?���>�d&��t����=;6�و��{���&V�B��=X��>D�>Ƃ,�ߋ���O��I��h��=N	�Ͽ�L.�� 5�`&���<��u�n�����þ��u����ݓ��-3��>�V8><5>\L{>�gB>�=J>L�P?-�f?�"�>��>q������6��{	�I����R罼�e��C�|���1��(�ɾ�C�d����re߾)?���<2�U��1�'��NZ���A��+?�>��Ͼ��I��K���þ�{��
��Ad����ھ�4�P(n�m��?A�6?k�y��TR�"D�/�J�R���AX?��KS����Ҿ">�i��;�=�>�r>�,�2�1��}T�.74?�$?X�����HI>T��4=)#?	��>��=r��>yJ+?^)�]U��>�Mo>J]�>�?K>������7�}�'?^�^?%����쑾d�x>˰�H��û
=�&(>]�?�F�<�)�>*g	=c6��\��]�X�ǣ(=LW?7{�>�"����~��cu���ˁ=nRl?��>g�>��b?:�L?K%���H�U��$�<o�<�OU?�u?-�4>ӹ���K־�翾'2??+g?�
�>�LN�3�Ӿ''�M3���?զk?�m%?Ho����p� K������j??��v?�r^�is�������V��<�>�[�>���>��9�-l�>�>?�
#��G������ Y4�-Þ?��@���?��;<6!�Ǚ�=�;?�\�>��O��>ƾ{��>���d�q=�"�>����eev�����P,�^�8?���?��>����������=�r���ݪ?���?õO�\�]>Ep*����|?��S�= H�>�o�>��ݽZ��D5���7���{��X=хw>\@�^��T?.ľ�kտ�cʿs���xf�"C��"?��=�U~�u�g�g�+^���S�Ɠ?���v�Y��>�7>��ǽ*F����y�$7�OF��ɂ�>Y-����n>�Z�}p���P���<Ւ�>(z�>f}p>0��󽾔<�?����IʿfN�����x?X?'+�?�X�?��?k�
<Ä����k�[�XL?�5i?F]`?S�x�(�F��C�� ]u?d����6�@�(���$�vSQ>�t@?���>�4���>b�>�Y�>C;��XB,�~9̿Z���%�~ݖ?B�?����>��?�!?�hj���侕�]��=��Z?ua�=ת�V`��a������h�>��?����"�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�!N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?c�>��?�h�=�^�>X�=,�����-�fi#>	$�=�?���?b�M?)I�>�Z�=n�8�`/�#VF�IHR��#��C�Z�>��a?�L?0Ab>cG�� b2��
!�B�ͽ�m1�7�輬N@���,���߽�5>K�=>%>{�D���Ҿ��?Hp�4�ؿ�i�� p'��54?;��>�?����t����;_?Az�>�6��+���%���B�]��?�G�??�?��׾�R̼�>>�>�I�>��Խ����P�����7>(�B?V��D��h�o�u�>���?�@�ծ?]i��	?���P��Ua~����7�d��=��7?�0�#�z>���>��=�nv�޻��X�s����>�B�?�{�?��>!�l?��o�P�B�{�1=:M�>Ϝk?�s?dQo���m�B>��?!������L��f?�
@u@`�^?*3���b��,I�9��+^�=��r>{{D>%Ͻ���Β���ܩ�]�"��_=0[�>|s�>��B>�-+>��>�>�����X)��.���?���p�����J��H�����諭�+�Qi�
��Ӻ=>���Mǅ�P!v�.m�����=i�S?C3S?$er?t- ?�H<�7�>���P&=��0��Ώ=&��>��1?��I?#�)?��=�9��Xc�2��F����e��S��>��J>t�>���>���>��B<͛J>187>&�>U��=�f=���;�j�<�T>�>�>=%�>�4W�0뭾�Y���U��!���ڌ�<	o�>gL�?���E�������	����)���F>��?�dL>B�����ѿ�����B?^t6�e)��=�����>~k5?��Y?Aq2>I�7��5�����<[>�z���@�=�v�������(��>ǔ??�i	>�4�=�h\��A0�Q�îS��϶>̿:?�q��L�;�VT�)�y��߾�>;��=pl*�w�.�Ȫ����2��k�y�s=iU?j� ?2�=��;�D��v����>�L>t�>��!��n>���^�:����J>=�q=!+9>�t?k�->�l�=���>g5��u2a��>F�@>"]*>RY<?J�$?b-D�M��������/�9�t>���>�q>���=݉J�� �=:%�>��^>�P�Sp������.K�GF>���+P��s��]=��ǽ���=�P~=d����E�z�Y=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ~M�>�����G���み�zi��fU=��>o�=?���0��+<!���?'�>���J���ǿ��r��a�>5��?%�?V�i�����hH����>���?��o?J�j>mľWW�@X3>c>?�tQ?|��>�N��$���?e��?�χ?��1>���?� �?׊?w��=}��<i������{2�=Y/%�Y�?��>����%���2���f���{�-x�z�4>���;��?%�u�;�Ǿ�\>-�f�����!�=8zk>,�>�x=�܍>���>���>L[w>/⼊��<��1�K?���?����2n�kD�<��=��^�#'?�J4?υ[�K�Ͼ�Ѩ>`�\?�?B[?�f�>����=��-迿�~��ɵ�<:�K>I5�>�G�>@%���@K>Y�Ծ&5D��n�>4З>,���?ھ�.��O���?�>�e!?Q��>�Ү=f�?� ?�yY>���>W9:�����{B��9�>�e�>"�?�>�?��?��޾�M9��/��̠�8�Y�&�v>�c}?ZL%?_�Q>-���G6��H�G<�e�<�;�=�^w?%�L?�i����><��?9N5?)I?]F->�����ξ�<`-�>?+����E�d�J��p���.�>��a?�?�B&>��^�����Kپ�@4���?�ן>�q?r� �&�;��Z�G^=��_� �<�k=-$�=}ت=���=v���F>���>A��=ci��ܾ��9e=��z>�>\+�>�VC��8�E
/?���<�Ȃ�̛=��^��O�Њm>�J1>�P��-�e?҅1�Uf�F&����)%�s��?��?�h�?y}r��>f��C&?�?x�"?��>�֛���㾑)��q����ٌ��I��d�=��><��<��Ѿ�L���s����c���fK���>�g�>��?v	?��=��>�蒾�,�_G�?���6Z@����h5�4�D��y+�dpw�ͅ�����=�ܶ��v��=>�^ǽ�?7R6?�0>eNa>L��>!	/>���>tc�>�,,>�J�>���>i_>ţ�>z�P��u���FR?|���q�'���;���a/B?�sd?�3�>�h����V���~?z�?�r�?��u>+oh�m3+��h?=-�>����e
?W�:=����ʈ<dI��@��d!��3G�K��> �׽h:�A
M��=f��a
?8?�ߎ�}̾-a׽ۑ����=Mv?�.?Έ"��X�mk��kI���D�6�����q�ƾ��%���p��I����r��z�ӎ.��]+<x�)?J;�?�>��:�ܾ����@oC���9�k&A>~��>_��>��>��> �#��%B��X�+R/�3o̾�?�6�?�è>q�O?�??��M?_\t?�� >
�v>|3�����>�P�=��->��?�zx?a��>�T?�0?ԅM?E? U=�_�F����-?�L?�$?��1?���>�w��Vg�X �0��;ʦ����I>�=ڡ����C�ɽf�,�"�r=��1?�)ɽ]&�B2��=D>B?u�?�]�>ppO�����?�<��?]E�>a/>���!v�
���
�> �?ﾼ<\�<Q=>�=<h�<���<b�,>c���&���c=�`+�1º�m��=�h=��ý@R0=�]w��Ī<%��=�d�>^�?���>�8�>�@���� �����<�=	Y>I�R>�y>�;پ�~��"&���g�Y!y>Pd�?Ul�?\�f=���=�u�=�v��T4����ỽ�-�<B�?�=#?�ZT?���?��=?J#?��>`)�gV��X^��"|��\�?4(?O��>t����̾���d�/�@?�7?�_���!��b'��j;�|߽m�>v�/���~��G��#qC�^�;���۫���E�?�{�?�� ��6����m�������B?���>/b�>F`�>`o(�'Wf�s>���@>��>�sN?�>�~[?�(�?
�m?��>�C"��C��Ö��-�<���<Ы??�Y�?{(l?�:X?_q�>�G�;�,�e�߾!>ݾK����0���E�ȍ=^�>���>�>�>�w�>a�>;���Y��SQ �t]�=�>�p�>~�>�Y�>�P>�r�;x�e?V?�sɾ��ʾC�����~�$�+��?l&�?�?`@2>WI����)�;�B�j[?��?���?%}O?��{��4�=P=Ȭ �I� �3�	?"!>��>�ǳ����}�>�����>�.� ���e�di�⛃>�kU?��;>T	���YZ�����;�x�l�����3����6<��B��r���*�j���W;ܾ{B���忾��þ���V,ʾ[�0����>�/�=�o=nU=u��<��
�W�D�b�52�=�xý��ռ�#>���{R=,ۜ��x�<�և<�w�<7���L˾��|?͖H?�d+?�C?:-y>�>�h2��Ζ>�y��+r?DU>E�R�oF��<�^���#����ؾ��־D�b��1���8>�I� �>wQ3>_��=�_�<�=5 u=�J�=����5=���=�Ϲ=�֭=�]�=>��>�6w?X�������4Q��Z罤�:?�8�>d{�=��ƾq@?�>>�2������yb��-?���?�T�?>�??ti��d�>N���㎽�q�=H����=2>p��=y�2�S��>��J>���K��@����4�?��@��??�ዿТϿ6a/>���=�+�=X����ݟ�t��������{?�&
�!�v�>�Qs�>y��举($Ľ�S�<����������5��r�=hB��w�<��t</jz>7nP>7k%>쇞���)>�j�<�{�=ڳ�>�L"���*=�§�/�%>�)1<�r�>�޷=4t?�"?�5?�`�?�5�>���6���WZ���>�����?��3>���>���>n�^?�e2?N�?�1�>������>\�>��K�/�_�4��/���W�'�W�?̽�?���>��=�5۽@i4�z�L��ѱ=6�S?��V?)�&?�^>"V�
�࿽Y&�ʛ.����P��+=�mr�]U�����6m�E��'�=�r�>#��>��>FSy>�9>�N>~�>�>�5�< r�=�������<)��3��=Y����+�<Jgż�튺�q&���+�͇��m��;Dk�;p�]<:*�;�y�=h��>ir>���>��=Kz����.>x�����L��=M��*B�'�c��0~�&/��^6�,�B>`%X>�ك�r'���?��Y>��?>�m�?�+u?��>�+�=�վ^C���d�iS��ɸ=�W>;�<�ht;��7`���M�x9Ҿ���>l�>�?�}~>f괾񷆿��:7:��$X��h4?��h�=G�6i-�sh�����Ɣ��,c���>�m?��)�w>\�L?��H?M1�?o��=�5'�@p潒G�=;FC����=3�����=m�0=h_?���>)�(?��C�c�!�x̾:n��?Y�>�HH��O�pꕿ�0�T�%��H��4��>�Ȫ���о^�2��k��X���B���r�S6�>��O?���?�'a��j����N��h�/$��H�?	�g?���>�?oV?�ՠ� ��Q�~����=zVn?��?��?�;>KC`=�:���?rp?�ٙ?�U�?�3R?? @��D�>�e>��r>�=
Y>(5�=��R=�=p>?&�?<[?�C#�ɧ �o�����k���6>{��=C?�>�e>���>6e'>�A�< ��=��>ܔ�>��s>�n>�E>�>�o���>���,?~�=��>�Y=?y�N>�\�;�37�v��>8a>%o��A�����H佸���{�=ly=s�C;�>��ÿ�?�MC>���)?�J꾃/L���k=/4 >]����>5�=�;>��>�>��U>��>{x�=I&���L>C�����6��+K��'�AYQ>���˹Q����w?��
��E��	�b\��y���)��&9=)�?B��;�W�/"��oƽ�2?\��>�'?�x��d|<tX>/.?.I>���R[������,����?R�? :c>��>��W?џ?�1��3�dwZ���u�="A��e���`��ލ�=���B�
�X���_?��x?tA?�'�<B5z>Z��?Y�%��ɏ�'!�>�/�= ;�N�<=�+�>�0��(�`�4�Ӿr�þ�8�IF>-�o?�#�?gZ?;DV�ͷ����F>�N?�E?c�^?,`X?�Z?�)�<X(?m,�Td�>�u�>cI?ia?�H?FJ>�z>偍�/�=�Mj��,��x������1�Pyo=�O>�=�<4�=B/>O�;�.O��f>�읽M7*��Q
>�ܺ=Q�=�
�>iLo?|��>�ۛ>�?M?Ֆ�$\�/���v�>�>N����mV�H��=��Ӿ�e�>��m?�s�?��?<��>�:_�=ra���m>{8Y>�{2>;��>I�>����ꊾ,��=�K >m@�=�=U�<�����s�n�S�"�q<��J>�}�>�<\>���$�>b󔾩s��O%>�~����D�{N�m�(���H��놾�i�>��%?�b?V)�=���A>y���g�cd3?�AV?��G?��Z?�A����A�H�+d���X�?њ=磾����K��oGW��?�=�]�=oG���<�ͽ}:��H��R���C8�cy��z\7>p�����=!i� ��%ǽuQ�=���>E֨���3�L����ԩ�*�e?q�=�O9�F�m�}-復$=>�Z?��?����2e�Piy��IW�+�E=Oa?"��<7U4>7���L����jF�>d�D?p�`?߅?gpz���k�S�B��-����������?;ۨ>��?�5K>�R�=� ��$�
��8b��$D�P��>�&�>:�ŗC�[q��sb��2%�iψ>i3?L�&>�?�NS?_�?�_^?�I,?zh?�ޕ>�Z��"տ��B'?�?��=�����R�r�9�"G���>�,?��?����>��?�?��$?��R?Ң?��>�A��a^?�Mڕ>�ȏ>x�Y�����*�a>¿I?Q��>��Y?MǄ?�k<>Q�3����;�Ž�/�=�W>�6?��"?��?Z�>���>��+��a>�xy>�K�?{�?aO~?�K
>;��>�)�>�u�=EV�=0C?v�>q?��=?�;y?�dF?��>����q;�MU?��@+� �f�5��!�p=rC=��\���&�}�"��o���v���=
7~=U����[���;�s������>��r>'���Rm0>�Bžp��Ac@>ߖ��5��l����9� G�=f�>��?Pڔ>�$�:�=|û>���>�����'?z7?�Z?��_;�b���ܾ��K�~�>��A?���=�/l��Z��ӽu�XNi=��m?�3^?��W�����h�b?)�]?xk�=��þ��b�p��u�O?y�
?��G���>��~?��q?���>}f��6n����Ab���j��ܶ=�n�>qU��d��<�>�7?+W�>	�b>�%�=?t۾t�w��l��]?��?T��?���?- *>Z�n��2�<��/~���CW?G�>ǀ��4?)����ȾV�������g ;�j���
������k"���6�g�s����s�=.�?[o?��o?��W?����`��yZ�:�����W�?!
�)G�:>��C��4O�j�Ǫ�d(�h��ZB�=R�n��)F��h�?&$?������?2���l�
�۾��>��w����0�=Z����<[��;R<(��t ��{��0?_�>)=�>y]?k�j��,�*27��U���۾�I�=���>�̱>^�>� ����N�Uiҽ�Ҿ�s���2�=�e>��h?�g?gwz?U�z�t���$����D�>1=#C����>�g�>�)>�@�Uƽ�&������h�{�	�?Cx�n4.���}�G4?�w�=���>{��?ɹ?M���]�ľ�j��Q�W���=1�[>���??@-x>�)"�6
�9��>�l?���>3�>�h��c!���{��˽���>���>���>��o>l�,��\��g��Ӄ��T�8���=�h?}��Ţ`��ۅ>L�Q?d�:|8G<�a�>�	v�в!�����'�O>�`?�<�=��;>�jž����{�5��X(?�?������+�F�l>D�?��>���>ن?�]�>�վ���`�?��d?�@?gG?)��> s]<]H�iٽt	�c�C=���>�~U>ob=��=��=�J��.��g=�=z?�`����_��,�5��<@;=9>����yx�����k0���w��{�ƾK������@Ľ����*�P�g��8���'>}�}�@M��>���m��i�?���?����3 =@������_��j�>-��8>@͓�5�.�Z�=o84��Z���!�7�h�����b��S$�> ¦��:̿�����,?��;?���?.�i�%��+[�*`�=�FB�8Bp�����V���:̿�ɾq�G?�>H?Z��oQ���>k9�>�޺=�Y>�ˣ��&��遾v�?�\�>\߁>?膾���26̿[��=#�?�8�?&yA?{�(�t��m'V=���> �	?|�?>�T1�G��ﰾ�J�>�;�?���?U`M=��W���	��}e?<<��F��4ݻ��=�X�=�z=���Q�J>�V�>Y���6A�\Cܽ&�4>�߅>��"�����^��ξ<�z]>�սB��4Մ?*{\��f���/��T��
U>��T?+�>�:�=��,?[7H�_}Ͽ�\��*a?�0�?���?�(?<ۿ��ؚ>��ܾ��M?]D6?���>�d&��t����=;6�و��{���&V�B��=X��>D�>Ƃ,�ߋ���O��I��h��=N	�Ͽ�L.�� 5�`&���<��u�n�����þ��u����ݓ��-3��>�V8><5>\L{>�gB>�=J>L�P?-�f?�"�>��>q������6��{	�I����R罼�e��C�|���1��(�ɾ�C�d����re߾)?���<2�U��1�'��NZ���A��+?�>��Ͼ��I��K���þ�{��
��Ad����ھ�4�P(n�m��?A�6?k�y��TR�"D�/�J�R���AX?��KS����Ҿ">�i��;�=�>�r>�,�2�1��}T�.74?�$?X�����HI>T��4=)#?	��>��=r��>yJ+?^)�]U��>�Mo>J]�>�?K>������7�}�'?^�^?%����쑾d�x>˰�H��û
=�&(>]�?�F�<�)�>*g	=c6��\��]�X�ǣ(=LW?7{�>�"����~��cu���ˁ=nRl?��>g�>��b?:�L?K%���H�U��$�<o�<�OU?�u?-�4>ӹ���K־�翾'2??+g?�
�>�LN�3�Ӿ''�M3���?զk?�m%?Ho����p� K������j??��v?�r^�is�������V��<�>�[�>���>��9�-l�>�>?�
#��G������ Y4�-Þ?��@���?��;<6!�Ǚ�=�;?�\�>��O��>ƾ{��>���d�q=�"�>����eev�����P,�^�8?���?��>����������=�r���ݪ?���?õO�\�]>Ep*����|?��S�= H�>�o�>��ݽZ��D5���7���{��X=хw>\@�^��T?.ľ�kտ�cʿs���xf�"C��"?��=�U~�u�g�g�+^���S�Ɠ?���v�Y��>�7>��ǽ*F����y�$7�OF��ɂ�>Y-����n>�Z�}p���P���<Ւ�>(z�>f}p>0��󽾔<�?����IʿfN�����x?X?'+�?�X�?��?k�
<Ä����k�[�XL?�5i?F]`?S�x�(�F��C�� ]u?d����6�@�(���$�vSQ>�t@?���>�4���>b�>�Y�>C;��XB,�~9̿Z���%�~ݖ?B�?����>��?�!?�hj���侕�]��=��Z?ua�=ת�V`��a������h�>��?����"�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�!N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?c�>��?�h�=�^�>X�=,�����-�fi#>	$�=�?���?b�M?)I�>�Z�=n�8�`/�#VF�IHR��#��C�Z�>��a?�L?0Ab>cG�� b2��
!�B�ͽ�m1�7�輬N@���,���߽�5>K�=>%>{�D���Ҿ��?Hp�4�ؿ�i�� p'��54?;��>�?����t����;_?Az�>�6��+���%���B�]��?�G�??�?��׾�R̼�>>�>�I�>��Խ����P�����7>(�B?V��D��h�o�u�>���?�@�ծ?]i��	?���P��Ua~����7�d��=��7?�0�#�z>���>��=�nv�޻��X�s����>�B�?�{�?��>!�l?��o�P�B�{�1=:M�>Ϝk?�s?dQo���m�B>��?!������L��f?�
@u@`�^?*3���b��,I�9��+^�=��r>{{D>%Ͻ���Β���ܩ�]�"��_=0[�>|s�>��B>�-+>��>�>�����X)��.���?���p�����J��H�����諭�+�Qi�
��Ӻ=>���Mǅ�P!v�.m�����=i�S?C3S?$er?t- ?�H<�7�>���P&=��0��Ώ=&��>��1?��I?#�)?��=�9��Xc�2��F����e��S��>��J>t�>���>���>��B<͛J>187>&�>U��=�f=���;�j�<�T>�>�>=%�>�4W�0뭾�Y���U��!���ڌ�<	o�>gL�?���E�������	����)���F>��?�dL>B�����ѿ�����B?^t6�e)��=�����>~k5?��Y?Aq2>I�7��5�����<[>�z���@�=�v�������(��>ǔ??�i	>�4�=�h\��A0�Q�îS��϶>̿:?�q��L�;�VT�)�y��߾�>;��=pl*�w�.�Ȫ����2��k�y�s=iU?j� ?2�=��;�D��v����>�L>t�>��!��n>���^�:����J>=�q=!+9>�t?k�->�l�=���>g5��u2a��>F�@>"]*>RY<?J�$?b-D�M��������/�9�t>���>�q>���=݉J�� �=:%�>��^>�P�Sp������.K�GF>���+P��s��]=��ǽ���=�P~=d����E�z�Y=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ~M�>�����G���み�zi��fU=��>o�=?���0��+<!���?'�>���J���ǿ��r��a�>5��?%�?V�i�����hH����>���?��o?J�j>mľWW�@X3>c>?�tQ?|��>�N��$���?e��?�χ?��1>���?� �?׊?w��=}��<i������{2�=Y/%�Y�?��>����%���2���f���{�-x�z�4>���;��?%�u�;�Ǿ�\>-�f�����!�=8zk>,�>�x=�܍>���>���>L[w>/⼊��<��1�K?���?����2n�kD�<��=��^�#'?�J4?υ[�K�Ͼ�Ѩ>`�\?�?B[?�f�>����=��-迿�~��ɵ�<:�K>I5�>�G�>@%���@K>Y�Ծ&5D��n�>4З>,���?ھ�.��O���?�>�e!?Q��>�Ү=f�?� ?�yY>���>W9:�����{B��9�>�e�>"�?�>�?��?��޾�M9��/��̠�8�Y�&�v>�c}?ZL%?_�Q>-���G6��H�G<�e�<�;�=�^w?%�L?�i����><��?9N5?)I?]F->�����ξ�<`-�>?+����E�d�J��p���.�>��a?�?�B&>��^�����Kپ�@4���?�ן>�q?r� �&�;��Z�G^=��_� �<�k=-$�=}ت=���=v���F>���>A��=ci��ܾ��9e=��z>�>\+�>�VC��8�E
/?���<�Ȃ�̛=��^��O�Њm>�J1>�P��-�e?҅1�Uf�F&����)%�s��?��?�h�?y}r��>f��C&?�?x�"?��>�֛���㾑)��q����ٌ��I��d�=��><��<��Ѿ�L���s����c���fK���>�g�>��?v	?��=��>�蒾�,�_G�?���6Z@����h5�4�D��y+�dpw�ͅ�����=�ܶ��v��=>�^ǽ�?7R6?�0>eNa>L��>!	/>���>tc�>�,,>�J�>���>i_>ţ�>z�P��u���FR?|���q�'���;���a/B?�sd?�3�>�h����V���~?z�?�r�?��u>+oh�m3+��h?=-�>����e
?W�:=����ʈ<dI��@��d!��3G�K��> �׽h:�A
M��=f��a
?8?�ߎ�}̾-a׽ۑ����=Mv?�.?Έ"��X�mk��kI���D�6�����q�ƾ��%���p��I����r��z�ӎ.��]+<x�)?J;�?�>��:�ܾ����@oC���9�k&A>~��>_��>��>��> �#��%B��X�+R/�3o̾�?�6�?�è>q�O?�??��M?_\t?�� >
�v>|3�����>�P�=��->��?�zx?a��>�T?�0?ԅM?E? U=�_�F����-?�L?�$?��1?���>�w��Vg�X �0��;ʦ����I>�=ڡ����C�ɽf�,�"�r=��1?�)ɽ]&�B2��=D>B?u�?�]�>ppO�����?�<��?]E�>a/>���!v�
���
�> �?ﾼ<\�<Q=>�=<h�<���<b�,>c���&���c=�`+�1º�m��=�h=��ý@R0=�]w��Ī<%��=�d�>^�?���>�8�>�@���� �����<�=	Y>I�R>�y>�;پ�~��"&���g�Y!y>Pd�?Ul�?\�f=���=�u�=�v��T4����ỽ�-�<B�?�=#?�ZT?���?��=?J#?��>`)�gV��X^��"|��\�?4(?O��>t����̾���d�/�@?�7?�_���!��b'��j;�|߽m�>v�/���~��G��#qC�^�;���۫���E�?�{�?�� ��6����m�������B?���>/b�>F`�>`o(�'Wf�s>���@>��>�sN?�>�~[?�(�?
�m?��>�C"��C��Ö��-�<���<Ы??�Y�?{(l?�:X?_q�>�G�;�,�e�߾!>ݾK����0���E�ȍ=^�>���>�>�>�w�>a�>;���Y��SQ �t]�=�>�p�>~�>�Y�>�P>�r�;x�e?V?�sɾ��ʾC�����~�$�+��?l&�?�?`@2>WI����)�;�B�j[?��?���?%}O?��{��4�=P=Ȭ �I� �3�	?"!>��>�ǳ����}�>�����>�.� ���e�di�⛃>�kU?��;>T	���YZ�����;�x�l�����3����6<��B��r���*�j���W;ܾ{B���忾��þ���V,ʾ[�0����>�/�=�o=nU=u��<��
�W�D�b�52�=�xý��ռ�#>���{R=,ۜ��x�<�և<�w�<7���L˾��|?͖H?�d+?�C?:-y>�>�h2��Ζ>�y��+r?DU>E�R�oF��<�^���#����ؾ��־D�b��1���8>�I� �>wQ3>_��=�_�<�=5 u=�J�=����5=���=�Ϲ=�֭=�]�=>��>�6w?X�������4Q��Z罤�:?�8�>d{�=��ƾq@?�>>�2������yb��-?���?�T�?>�??ti��d�>N���㎽�q�=H����=2>p��=y�2�S��>��J>���K��@����4�?��@��??�ዿТϿ6a/>���=�+�=X����ݟ�t��������{?�&
�!�v�>�Qs�>y��举($Ľ�S�<����������5��r�=hB��w�<��t</jz>7nP>7k%>쇞���)>�j�<�{�=ڳ�>�L"���*=�§�/�%>�)1<�r�>�޷=4t?�"?�5?�`�?�5�>���6���WZ���>�����?��3>���>���>n�^?�e2?N�?�1�>������>\�>��K�/�_�4��/���W�'�W�?̽�?���>��=�5۽@i4�z�L��ѱ=6�S?��V?)�&?�^>"V�
�࿽Y&�ʛ.����P��+=�mr�]U�����6m�E��'�=�r�>#��>��>FSy>�9>�N>~�>�>�5�< r�=�������<)��3��=Y����+�<Jgż�튺�q&���+�͇��m��;Dk�;p�]<:*�;�y�=h��>ir>���>��=Kz����.>x�����L��=M��*B�'�c��0~�&/��^6�,�B>`%X>�ك�r'���?��Y>��?>�m�?�+u?��>�+�=�վ^C���d�iS��ɸ=�W>;�<�ht;��7`���M�x9Ҿ���>l�>�?�}~>f괾񷆿��:7:��$X��h4?��h�=G�6i-�sh�����Ɣ��,c���>�m?��)�w>\�L?��H?M1�?o��=�5'�@p潒G�=;FC����=3�����=m�0=h_?���>)�(?��C�c�!�x̾:n��?Y�>�HH��O�pꕿ�0�T�%��H��4��>�Ȫ���о^�2��k��X���B���r�S6�>��O?���?�'a��j����N��h�/$��H�?	�g?���>�?oV?�ՠ� ��Q�~����=zVn?��?��?�;>KC`=�:���?rp?�ٙ?�U�?�3R?? @��D�>�e>��r>�=
Y>(5�=��R=�=p>?&�?<[?�C#�ɧ �o�����k���6>{��=C?�>�e>���>6e'>�A�< ��=��>ܔ�>��s>�n>�E>�>�o���>���,?~�=��>�Y=?y�N>�\�;�37�v��>8a>%o��A�����H佸���{�=ly=s�C;�>��ÿ�?�MC>���)?�J꾃/L���k=/4 >]����>5�=�;>��>�>��U>��>{x�=I&���L>C�����6��+K��'�AYQ>���˹Q����w?��
��E��	�b\��y���)��&9=)�?B��;�W�/"��oƽ�2?\��>�'?�x��d|<tX>/.?.I>���R[������,����?R�? :c>��>��W?џ?�1��3�dwZ���u�="A��e���`��ލ�=���B�
�X���_?��x?tA?�'�<B5z>Z��?Y�%��ɏ�'!�>�/�= ;�N�<=�+�>�0��(�`�4�Ӿr�þ�8�IF>-�o?�#�?gZ?;DV�ͷ����F>�N?�E?c�^?,`X?�Z?�)�<X(?m,�Td�>�u�>cI?ia?�H?FJ>�z>偍�/�=�Mj��,��x������1�Pyo=�O>�=�<4�=B/>O�;�.O��f>�읽M7*��Q
>�ܺ=Q�=�
�>iLo?|��>�ۛ>�?M?Ֆ�$\�/���v�>�>N����mV�H��=��Ӿ�e�>��m?�s�?��?<��>�:_�=ra���m>{8Y>�{2>;��>I�>����ꊾ,��=�K >m@�=�=U�<�����s�n�S�"�q<��J>�}�>�<\>���$�>b󔾩s��O%>�~����D�{N�m�(���H��놾�i�>��%?�b?V)�=���A>y���g�cd3?�AV?��G?��Z?�A����A�H�+d���X�?њ=磾����K��oGW��?�=�]�=oG���<�ͽ}:��H��R���C8�cy��z\7>p�����=!i� ��%ǽuQ�=���>E֨���3�L����ԩ�*�e?q�=�O9�F�m�}-復$=>�Z?��?����2e�Piy��IW�+�E=Oa?"��<7U4>7���L����jF�>d�D?p�`?߅?gpz���k�S�B��-����������?;ۨ>��?�5K>�R�=� ��$�
��8b��$D�P��>�&�>:�ŗC�[q��sb��2%�iψ>i3?L�&>�?�NS?_�?�_^?�I,?zh?�ޕ>�Z��"տ��B'?�?��=�����R�r�9�"G���>�,?��?����>��?�?��$?��R?Ң?��>�A��a^?�Mڕ>�ȏ>x�Y�����*�a>¿I?Q��>��Y?MǄ?�k<>Q�3����;�Ž�/�=�W>�6?��"?��?Z�>���>��+��a>�xy>�K�?{�?aO~?�K
>;��>�)�>�u�=EV�=0C?v�>q?��=?�;y?�dF?��>����q;�MU?��@+� �f�5��!�p=rC=��\���&�}�"��o���v���=
7~=U����[���;�s������>��r>'���Rm0>�Bžp��Ac@>ߖ��5��l����9� G�=f�>��?Pڔ>�$�:�=|û>���>�����'?z7?�Z?��_;�b���ܾ��K�~�>��A?���=�/l��Z��ӽu�XNi=��m?�3^?��W�����h�b?)�]?xk�=��þ��b�p��u�O?y�
?��G���>��~?��q?���>}f��6n����Ab���j��ܶ=�n�>qU��d��<�>�7?+W�>	�b>�%�=?t۾t�w��l��]?��?T��?���?- *>Z�n��2�<��/~���CW?G�>ǀ��4?)����ȾV�������g ;�j���
������k"���6�g�s����s�=.�?[o?��o?��W?����`��yZ�:�����W�?!
�)G�:>��C��4O�j�Ǫ�d(�h��ZB�=R�n��)F��h�?&$?������?2���l�
�۾��>��w����0�=Z����<[��;R<(��t ��{��0?_�>)=�>y]?k�j��,�*27��U���۾�I�=���>�̱>^�>� ����N�Uiҽ�Ҿ�s���2�=�e>��h?�g?gwz?U�z�t���$����D�>1=#C����>�g�>�)>�@�Uƽ�&������h�{�	�?Cx�n4.���}�G4?�w�=���>{��?ɹ?M���]�ľ�j��Q�W���=1�[>���??@-x>�)"�6
�9��>�l?���>3�>�h��c!���{��˽���>���>���>��o>l�,��\��g��Ӄ��T�8���=�h?}��Ţ`��ۅ>L�Q?d�:|8G<�a�>�	v�в!�����'�O>�`?�<�=��;>�jž����{�5��X(?�?������+�F�l>D�?��>���>ن?�]�>�վ���`�?��d?�@?gG?)��> s]<]H�iٽt	�c�C=���>�~U>ob=��=��=�J��.��g=�=z?�`����_��,�5��<@;=9>����yx�����k0���w��{�ƾK������@Ľ����*�P�g��8���'>}�}�@M��>���m��i�?���?����3 =@������_��j�>-��8>@͓�5�.�Z�=o84��Z���!�7�h�����b��S$�> ¦��:̿�����,?��;?���?.�i�%��+[�*`�=�FB�8Bp�����V���:̿�ɾq�G?�>H?Z��oQ���>k9�>�޺=�Y>�ˣ��&��遾v�?�\�>\߁>?膾���26̿[��=#�?�8�?&yA?{�(�t��m'V=���> �	?|�?>�T1�G��ﰾ�J�>�;�?���?U`M=��W���	��}e?<<��F��4ݻ��=�X�=�z=���Q�J>�V�>Y���6A�\Cܽ&�4>�߅>��"�����^��ξ<�z]>�սB��4Մ?*{\��f���/��T��
U>��T?+�>�:�=��,?[7H�_}Ͽ�\��*a?�0�?���?�(?<ۿ��ؚ>��ܾ��M?]D6?���>�d&��t����=;6�و��{���&V�B��=X��>D�>Ƃ,�ߋ���O��I��h��=N	�Ͽ�L.�� 5�`&���<��u�n�����þ��u����ݓ��-3��>�V8><5>\L{>�gB>�=J>L�P?-�f?�"�>��>q������6��{	�I����R罼�e��C�|���1��(�ɾ�C�d����re߾)?���<2�U��1�'��NZ���A��+?�>��Ͼ��I��K���þ�{��
��Ad����ھ�4�P(n�m��?A�6?k�y��TR�"D�/�J�R���AX?��KS����Ҿ">�i��;�=�>�r>�,�2�1��}T�.74?�$?X�����HI>T��4=)#?	��>��=r��>yJ+?^)�]U��>�Mo>J]�>�?K>������7�}�'?^�^?%����쑾d�x>˰�H��û
=�&(>]�?�F�<�)�>*g	=c6��\��]�X�ǣ(=LW?7{�>�"����~��cu���ˁ=nRl?��>g�>��b?:�L?K%���H�U��$�<o�<�OU?�u?-�4>ӹ���K־�翾'2??+g?�
�>�LN�3�Ӿ''�M3���?զk?�m%?Ho����p� K������j??��v?�r^�is�������V��<�>�[�>���>��9�-l�>�>?�
#��G������ Y4�-Þ?��@���?��;<6!�Ǚ�=�;?�\�>��O��>ƾ{��>���d�q=�"�>����eev�����P,�^�8?���?��>����������=�r���ݪ?���?õO�\�]>Ep*����|?��S�= H�>�o�>��ݽZ��D5���7���{��X=хw>\@�^��T?.ľ�kտ�cʿs���xf�"C��"?��=�U~�u�g�g�+^���S�Ɠ?���v�Y��>�7>��ǽ*F����y�$7�OF��ɂ�>Y-����n>�Z�}p���P���<Ւ�>(z�>f}p>0��󽾔<�?����IʿfN�����x?X?'+�?�X�?��?k�
<Ä����k�[�XL?�5i?F]`?S�x�(�F��C�� ]u?d����6�@�(���$�vSQ>�t@?���>�4���>b�>�Y�>C;��XB,�~9̿Z���%�~ݖ?B�?����>��?�!?�hj���侕�]��=��Z?ua�=ת�V`��a������h�>��?����"�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�!N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?c�>��?�h�=�^�>X�=,�����-�fi#>	$�=�?���?b�M?)I�>�Z�=n�8�`/�#VF�IHR��#��C�Z�>��a?�L?0Ab>cG�� b2��
!�B�ͽ�m1�7�輬N@���,���߽�5>K�=>%>{�D���Ҿ��?Hp�4�ؿ�i�� p'��54?;��>�?����t����;_?Az�>�6��+���%���B�]��?�G�??�?��׾�R̼�>>�>�I�>��Խ����P�����7>(�B?V��D��h�o�u�>���?�@�ծ?]i��	?���P��Ua~����7�d��=��7?�0�#�z>���>��=�nv�޻��X�s����>�B�?�{�?��>!�l?��o�P�B�{�1=:M�>Ϝk?�s?dQo���m�B>��?!������L��f?�
@u@`�^?*3���b��,I�9��+^�=��r>{{D>%Ͻ���Β���ܩ�]�"��_=0[�>|s�>��B>�-+>��>�>�����X)��.���?���p�����J��H�����諭�+�Qi�
��Ӻ=>���Mǅ�P!v�.m�����=i�S?C3S?$er?t- ?�H<�7�>���P&=��0��Ώ=&��>��1?��I?#�)?��=�9��Xc�2��F����e��S��>��J>t�>���>���>��B<͛J>187>&�>U��=�f=���;�j�<�T>�>�>=%�>�4W�0뭾�Y���U��!���ڌ�<	o�>gL�?���E�������	����)���F>��?�dL>B�����ѿ�����B?^t6�e)��=�����>~k5?��Y?Aq2>I�7��5�����<[>�z���@�=�v�������(��>ǔ??�i	>�4�=�h\��A0�Q�îS��϶>̿:?�q��L�;�VT�)�y��߾�>;��=pl*�w�.�Ȫ����2��k�y�s=iU?j� ?2�=��;�D��v����>�L>t�>��!��n>���^�:����J>=�q=!+9>�t?k�->�l�=���>g5��u2a��>F�@>"]*>RY<?J�$?b-D�M��������/�9�t>���>�q>���=݉J�� �=:%�>��^>�P�Sp������.K�GF>���+P��s��]=��ǽ���=�P~=d����E�z�Y=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ~M�>�����G���み�zi��fU=��>o�=?���0��+<!���?'�>���J���ǿ��r��a�>5��?%�?V�i�����hH����>���?��o?J�j>mľWW�@X3>c>?�tQ?|��>�N��$���?e��?�χ?��1>���?� �?׊?w��=}��<i������{2�=Y/%�Y�?��>����%���2���f���{�-x�z�4>���;��?%�u�;�Ǿ�\>-�f�����!�=8zk>,�>�x=�܍>���>���>L[w>/⼊��<��1�K?���?����2n�kD�<��=��^�#'?�J4?υ[�K�Ͼ�Ѩ>`�\?�?B[?�f�>����=��-迿�~��ɵ�<:�K>I5�>�G�>@%���@K>Y�Ծ&5D��n�>4З>,���?ھ�.��O���?�>�e!?Q��>�Ү=f�?� ?�yY>���>W9:�����{B��9�>�e�>"�?�>�?��?��޾�M9��/��̠�8�Y�&�v>�c}?ZL%?_�Q>-���G6��H�G<�e�<�;�=�^w?%�L?�i����><��?9N5?)I?]F->�����ξ�<`-�>?+����E�d�J��p���.�>��a?�?�B&>��^�����Kپ�@4���?�ן>�q?r� �&�;��Z�G^=��_� �<�k=-$�=}ت=���=v���F>���>A��=ci��ܾ��9e=��z>�>\+�>�VC��8�E
/?���<�Ȃ�̛=��^��O�Њm>�J1>�P��-�e?҅1�Uf�F&����)%�s��?��?�h�?y}r��>f��C&?�?x�"?��>�֛���㾑)��q����ٌ��I��d�=��><��<��Ѿ�L���s����c���fK���>�g�>��?v	?��=��>�蒾�,�_G�?���6Z@����h5�4�D��y+�dpw�ͅ�����=�ܶ��v��=>�^ǽ�?7R6?�0>eNa>L��>!	/>���>tc�>�,,>�J�>���>i_>ţ�>z�P��u���FR?|���q�'���;���a/B?�sd?�3�>�h����V���~?z�?�r�?��u>+oh�m3+��h?=-�>����e
?W�:=����ʈ<dI��@��d!��3G�K��> �׽h:�A
M��=f��a
?8?�ߎ�}̾-a׽ۑ����=Mv?�.?Έ"��X�mk��kI���D�6�����q�ƾ��%���p��I����r��z�ӎ.��]+<x�)?J;�?�>��:�ܾ����@oC���9�k&A>~��>_��>��>��> �#��%B��X�+R/�3o̾�?�6�?�è>q�O?�??��M?_\t?�� >
�v>|3�����>�P�=��->��?�zx?a��>�T?�0?ԅM?E? U=�_�F����-?�L?�$?��1?���>�w��Vg�X �0��;ʦ����I>�=ڡ����C�ɽf�,�"�r=��1?�)ɽ]&�B2��=D>B?u�?�]�>ppO�����?�<��?]E�>a/>���!v�
���
�> �?ﾼ<\�<Q=>�=<h�<���<b�,>c���&���c=�`+�1º�m��=�h=��ý@R0=�]w��Ī<%��=�d�>^�?���>�8�>�@���� �����<�=	Y>I�R>�y>�;پ�~��"&���g�Y!y>Pd�?Ul�?\�f=���=�u�=�v��T4����ỽ�-�<B�?�=#?�ZT?���?��=?J#?��>`)�gV��X^��"|��\�?4(?O��>t����̾���d�/�@?�7?�_���!��b'��j;�|߽m�>v�/���~��G��#qC�^�;���۫���E�?�{�?�� ��6����m�������B?���>/b�>F`�>`o(�'Wf�s>���@>��>�sN?�>�~[?�(�?
�m?��>�C"��C��Ö��-�<���<Ы??�Y�?{(l?�:X?_q�>�G�;�,�e�߾!>ݾK����0���E�ȍ=^�>���>�>�>�w�>a�>;���Y��SQ �t]�=�>�p�>~�>�Y�>�P>�r�;x�e?V?�sɾ��ʾC�����~�$�+��?l&�?�?`@2>WI����)�;�B�j[?��?���?%}O?��{��4�=P=Ȭ �I� �3�	?"!>��>�ǳ����}�>�����>�.� ���e�di�⛃>�kU?��;>T	���YZ�����;�x�l�����3����6<��B��r���*�j���W;ܾ{B���忾��þ���V,ʾ[�0����>�/�=�o=nU=u��<��
�W�D�b�52�=�xý��ռ�#>���{R=,ۜ��x�<�և<�w�<7���L˾��|?͖H?�d+?�C?:-y>�>�h2��Ζ>�y��+r?DU>E�R�oF��<�^���#����ؾ��־D�b��1���8>�I� �>wQ3>_��=�_�<�=5 u=�J�=����5=���=�Ϲ=�֭=�]�=>��>�6w?X�������4Q��Z罤�:?�8�>d{�=��ƾq@?�>>�2������yb��-?���?�T�?>�??ti��d�>N���㎽�q�=H����=2>p��=y�2�S��>��J>���K��@����4�?��@��??�ዿТϿ6a/>���=�+�=X����ݟ�t��������{?�&
�!�v�>�Qs�>y��举($Ľ�S�<����������5��r�=hB��w�<��t</jz>7nP>7k%>쇞���)>�j�<�{�=ڳ�>�L"���*=�§�/�%>�)1<�r�>�޷=4t?�"?�5?�`�?�5�>���6���WZ���>�����?��3>���>���>n�^?�e2?N�?�1�>������>\�>��K�/�_�4��/���W�'�W�?̽�?���>��=�5۽@i4�z�L��ѱ=6�S?��V?)�&?�^>"V�
�࿽Y&�ʛ.����P��+=�mr�]U�����6m�E��'�=�r�>#��>��>FSy>�9>�N>~�>�>�5�< r�=�������<)��3��=Y����+�<Jgż�튺�q&���+�͇��m��;Dk�;p�]<:*�;�y�=h��>ir>���>��=Kz����.>x�����L��=M��*B�'�c��0~�&/��^6�,�B>`%X>�ك�r'���?��Y>��?>�m�?�+u?��>�+�=�վ^C���d�iS��ɸ=�W>;�<�ht;��7`���M�x9Ҿ���>l�>�?�}~>f괾񷆿��:7:��$X��h4?��h�=G�6i-�sh�����Ɣ��,c���>�m?��)�w>\�L?��H?M1�?o��=�5'�@p潒G�=;FC����=3�����=m�0=h_?���>)�(?��C�c�!�x̾:n��?Y�>�HH��O�pꕿ�0�T�%��H��4��>�Ȫ���о^�2��k��X���B���r�S6�>��O?���?�'a��j����N��h�/$��H�?	�g?���>�?oV?�ՠ� ��Q�~����=zVn?��?��?�;>KC`=�:���?rp?�ٙ?�U�?�3R?? @��D�>�e>��r>�=
Y>(5�=��R=�=p>?&�?<[?�C#�ɧ �o�����k���6>{��=C?�>�e>���>6e'>�A�< ��=��>ܔ�>��s>�n>�E>�>�o���>���,?~�=��>�Y=?y�N>�\�;�37�v��>8a>%o��A�����H佸���{�=ly=s�C;�>��ÿ�?�MC>���)?�J꾃/L���k=/4 >]����>5�=�;>��>�>��U>��>{x�=I&���L>C�����6��+K��'�AYQ>���˹Q����w?��
��E��	�b\��y���)��&9=)�?B��;�W�/"��oƽ�2?\��>�'?�x��d|<tX>/.?.I>���R[������,����?R�? :c>��>��W?џ?�1��3�dwZ���u�="A��e���`��ލ�=���B�
�X���_?��x?tA?�'�<B5z>Z��?Y�%��ɏ�'!�>�/�= ;�N�<=�+�>�0��(�`�4�Ӿr�þ�8�IF>-�o?�#�?gZ?;DV�ͷ����F>�N?�E?c�^?,`X?�Z?�)�<X(?m,�Td�>�u�>cI?ia?�H?FJ>�z>偍�/�=�Mj��,��x������1�Pyo=�O>�=�<4�=B/>O�;�.O��f>�읽M7*��Q
>�ܺ=Q�=�
�>iLo?|��>�ۛ>�?M?Ֆ�$\�/���v�>�>N����mV�H��=��Ӿ�e�>��m?�s�?��?<��>�:_�=ra���m>{8Y>�{2>;��>I�>����ꊾ,��=�K >m@�=�=U�<�����s�n�S�"�q<��J>�}�>�<\>���$�>b󔾩s��O%>�~����D�{N�m�(���H��놾�i�>��%?�b?V)�=���A>y���g�cd3?�AV?��G?��Z?�A����A�H�+d���X�?њ=磾����K��oGW��?�=�]�=oG��`��� >���fܾ,6l�K�%�,�V->|� �����b �/�ܾ�-���߅�ɛ�>��þR0*�0Z��R.���eF?u�[���ϾV��ʾ��,>ݠ>��>�*�=�V�=��^���ž>ne#?�&>�
��/о�Q+�/h����|>/�K?�^? �?~�p���z���K�2#�^⇾�?P�e! ?�/�>[��>ġi>2=�þ�����Z�!/:�7,�>~��>q#���R����9������D�>��>�
>�]?�aH?9#?�4[?��1?�e?�>Z������G�$??�(�=��ǽʽO�e�8�(�F�.��>�o*?��F�	%�>��?K�?Y�'?L�M?�?�u>����&=���>�Ȇ>�Y��9���z]>ͿM?�'�>�X?؂?��6>�#3��蝾�Z�c��=�>x08?�x%?�m?I�>N?wzd�Ȇ�>�	?���?�I�?@S�?��5>�z�>z�?��>)�"�eYV>)#>��>�D?Z�?�,q?!�?�X�<o���-�h�MxG�ּ��=�/ =�e�5��;�[B�K����B=굂���=���qݽfe��cd�C(H����>As>���'�/>��ľ�@��IZA>JП�>W�����K�;�|��=��>��?je�>�#��i�=�o�>��>O���(?�??�*;�b��@۾��L�4��>��A?"��=��l�oC��:�u��2c=b�m? �^?��W�����b?�]?�g�=���þ��b�.����O?<�
?[�G�I�>��~?#�q?o��>�e�+:n�����Cb���j�
Ѷ=�q�>�X�|�d�U?�>��7?�N�>5�b>�$�=Wu۾��w��q���?s�?�?���?�+*>L�n�94�+���3Ǐ��)f?��>r5��5�?E	�<@��k���V󇾴�ݾ���N���s9v� ���H������Խ
��=7�?�o?T�g?�^t?���f�T�f�`�\���� S�0��/���A5���E��B��r���٠�ӂ����='���ì>����?s�!?���'��>w�H��	���Ǿ��F>����0�y�f=]��<{���#�K}��#�sM��H�"?ߨ�>�)�>Ϣd?������J�5��U���
�m=�{W>"��>>�A�C	]�������"��3�n>Msf?�+K?>�m?���֘5��*��f�(���꼥X��ga>q[>��>�8����(�ͭ5�}m��
��t��V�	��T�<ԟ"?smz>䜲>���?��	?��z��Fgt�M�,�I��=gƽ>��j?�W?~1�>΂Ž` �ӷ�>��l?���>��>Ӑ��lX!���{���ʽ\(�>׭>���>��o>��,��\��i��^���@9��h�=3�h?Â����`��>�R?��:DoG<�|�>��v�޾!����F�'�]�>Ty?Z��=Ұ;>q�ž�(���{�|0���i)?�*?�ݒ��4*�v�>v!?�N�>C��>f��?-b�>�����븺��?��]?H?~QA?�b�>a]/=%g���-Ž!y'�-.=TA�>�	[>�i=R|�=���[]�!�?�A=�=E����ýAa<`K��-9<���<��4>|kۿx9K�ޏپ���v��PG
��ψ�ߖ���Y�����[��1���/x�>}��'��V�O@c�������l��|�?g9�?����+��P�����������e��> Wq�4,�K���X���*������¬��a!��O�{#i�a�e�x�*?m��hrſ��Ae�c&!?7,?�Dt?:��I��&j<�_�>ٜ�:B��$!;����n�˿N���Y?��>�Ծ�μU�>��>�>$8�>����7���cn=���>��*?&��>igV�Vǿ�淿�S ����?,�@hlA?W�(�1��RV=l��>7�	?H5?>[�1�(��!���z�>�?�?��?��N=a�W�ގ�ǂe?=c�;�F���ۻ�X�=�W�=��=���J>�6�>����vA���ܽ�4>G��>t<"����"a^�Iƺ<#Z]>��ս�ꔽ5Մ?,{\��f���/��T��	U>��T? +�>K:�=��,?Y7H�`}Ͽ�\��*a?�0�?���?#�(?:ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=�6ἃ���x���&V����=T��>d�>Ȃ,������O��I��Y��=2���Zƿ\�$�����I=Vm��]U������8"M�����wo�w��Ɍh=k��=;Q>۝�>�UV>�Z>5�V?I�k?B��>Q�>�K�T����[;(���#��^	���S��壾*V�Ԥ߾w	���J��h�ɾ6���8彞7Z�o����O��;H��m��I;?���<��
� �?��p���S�5���>?q���'[�'[����=?>;8~�l�G�F�d�8,��6Ծ��vf?���<��A�����~0>�1!�����w�>$�j�X�=����p�p��33?�;?�ҽ��C��17>����O=I)?M�?}J=��>�C? �"��+����J>b�E> :�>Kg�>��'>K����/��� ?�U?G���❾�ۋ>.���4׉��b-=��>_ +�n�Ӽ�EI>;��<l>��
'������8H<!=W?�H�>��)����������	�==�Px?�?Ġ>cKk?߁B?�j�<�.����S��
���}=KX?�[i?ݰ>p�����Ͼ>h���5?	Je?uN>L�g�����.��@�|�?2�n?��?�c��Q	}�(��ؼ��f6?7�v?�j^��o��b��*�V��2�>�X�>��>c�9��r�>�>?�#��D����-X4�gĞ?��@B��?'�=<]+�N��=*A?�c�>�O�j4ƾ�Z��9z��Yq=�!�>b����av����W,�ƈ8?�?��>���v����=i,��Zu�?���?�:���½�:�������ݾDV�Z >���_���`x�`�z3�bx����<ˈ>�Z@�n�?e?)$E��DͿ��ӿ;���U��o���_H?R�>�=��T���%��dh^�\�e�8��uʽ�s�>�>-���������{�Gi9��Լ&�>����>ƦX��P��pM����;;�>!O�>(�>���][���^�?r���Cο�������X?�<�?�^�?�?81�<6l|��/{�yH��:I?G�r?��X?���&�Z����j�j?q���`���4��E��T>�>3?�n�>th-�7|=gD>��>��>|�.�=Ŀ�����V�����?m6�?���E�>��?r:+?yE��I��f��qc+��	��|FA?C�2>���!���<��)���}
?�0?����O�Y�_?(�a�O�p���-���ƽ�ۡ>��0��e\�
N�����Xe�
���@y����?K^�?d�?��� #�d6%?%�>a����8ǾC�<���>�(�>,*N>�H_���u>����:�i	>���?�~�?Lj?���������U>�}?w#�>/�?y�=�b�>�k�=��e�-�_#>��=F?�K�?�M?FP�>Jd�=��8�</�YF��FR�"�+�C�'�>��a?�L?/Qb>/��p2�!���ͽ�`1�57鼺V@�Ǘ,��߽(5>j�=>>��D�E
Ӿ��?Mp�9�ؿ j�� p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>D�Խ����]�����7>1�B?Y��D��u�o�y�>���?
�@�ծ?ji��	?���P��2a~�߂�&7���=��7?0��z>���>��=�nv�Ի��O�s���>�B�?�{�?���>�l?��o��B���1=IM�>��k?�s?41o��󾿱B>z�?������
L��f?�
@qu@*�^?�X��7������������=�[�=Y�B>ۢ������T=F��<Y�콠��=ng�>��~>bo4>޺M>�.>@8�=����0!������5��s }��:,���0�R^�%{���þ{��w���
�<��u=�]?���ľ��پ�"¾+d�=��T?5�S?o�t?[3?j�
��%�=���pT���]���=wU�>�`@?r.Q?m�'?��
=�O��"�^�o�t������&��!��>=n[>��>+��>T��>��<W�>L>��>�I�=��<ڹ<�|<��$>���>E/�>�}�>/#n�f �+F��&��/k��e^�=k�覢?�ǳ���H� -��(����?̾��>�ew?�ʽ����\?��_&��WaI?�7���U�����o��>ur?$�t?� ��ɐ�!�>�m����>M��H�8=Q$O�Ip>f�ž�r�>�H�>,w;>�t>}r6�E�G�PG�)�Ľ�P>�:6?�R������u������ݣ��	<�a[�>5�2>=52�麊�4>]�=y���<>z�8?�>���о�)ƾ�Bv��߾<�o̼�d>�����9>��w�\f�������ː=�-��C>��?Ò8>8؏=8h�>����7�R�@�>��?>Ǒ>>8*C?��#?�K��d��/b����4���>�*�><j�>ŏ>o!G�W�=%m�>��f>"����|�yk�_.1�3/H>&���<	\�o2r����=S�����=h��=R%�%�@�.=�~?���*䈿��ae���lD?_+?� �=U�F<��"�B ���H��8�?j�@m�?��	��V�+�?�@�?�
��q��=}�>�֫>�ξ;�L��?��ŽJǢ���	�J)#�cS�?��?D�/�[ʋ�:l�/6>�^%?�ӾKh�>�x��Z�������u��#=E��>�8H?�V����O��>��v
?�?�^�ѩ����ȿ3|v����>M�?���?]�m��A���@����>3��?�gY?joi>�g۾`Z����>ͻ@?�R?&�>�9�x�'�|�?�޶?ׯ�?e#>N��?���?�%#?("f��Rc����������>����b��>7�t>y� �����⠿wݘ�tB�4}�50�>$p�<�!?tlC�R���V;>2�:��`վ�	�=��>�7�>��A>���>���>Ϯ>��.?J.�:]��=/�H�ʤ����K?���?-���2n��N�<t��=+�^��&?�I4?�k[�|�Ͼ�ը>�\?h?�[?d�><��O>��E迿5~��ɪ�<��K>*4�>�H�>�$���FK>��Ծ�4D�Yp�>�ϗ>�����?ھ�,��{S��BB�>�e!?���>�Ү=�� ?��#?��j>�l�>pRE��?��3�E��E�>���>z-?�~?�?��h63�����顿!�[��N> �x??G?��>χ������XA��yJ�w���*��?<kg?�(��
?1�?K}??>�A?k�f>��^�׾-����Հ>�?@Bz��G��P8��t� �?��?�*�>߯Խv׽ErG�U����Sо ��>u�S?��A?�c�YxS�y����/=��C>!M!=�i�Bx�<���=>p�=+U��a`5>�.�=��=�L�x�ͽ�:�1T=���>yق=��b�w�=]J,?1�A�����kڙ=�r�glD�!�>(bL>%���+�^?@=��{�M����x���U��	�?3��?�n�?W³�b�h��=?�(�?�?��>�Į��޾nU��w�@�w�bS��W>���>�l����苤����l8��+�ǽ�
q�ʋ�>s�>A,
?�#?U��=�>����U0��ƾ7����_�_����$�~%.�]�)���{+ ��L�;g�&�0�?>�׼�8�>�i?�"�>�4�>���>K�|��>�o*>>��>�U�>�ԡ>"�R>��=�Q8�*�(�.IR?$����(��[�l��//B?��d?���>�m�;?��a�� ?�)�?r�?VJw>�h�tn+��?�"�>[M~��1
?�A=�%��n�<4ͷ����Qύ�2��<�>�-ؽ�9��M�/e�O\	?L�? 8��؝˾f�ս�D����t=�r�?gD+?X)��#R���n�8}Y�NfQ��	��`�ೠ�>�$�};n���d������ (��i5=��)?@Չ?V���1��n��0�k�sQ@�ճb>F��>rt�>K��>��K> �	� 0���]�.'�1F���_�>7�z?s2�>��M?��3?�U?&`G?K�>˖'>���6,�>�K�o��>��?�X?�>.?��?�1?X�'?��>�ɯ����Ȧ׾��?ڟ?�?���>{� ?�_������o9�J���	iB��ſ���=,>��[���Y����=iR^>U�3?���4;�����>�I(?!?�4�>�7��©C��CO����>�؁>Mބ>¾|ht���)�5��>v�n?�௼�n(=�=�>\�=*3=Q���s�;6+�<�M>[��@ǘ��-һ[@�=��c=�n��������<�X>-������>�?�i�>C�>kᅾ~� �}�����=��Z>x�S>H">�iپ�u�������g�L�y>$��?+��?g�j=���=-�=񄠾_e��{���ཾ�8�<��?W+#?<\T?�z�?��=?r#?{J>9��1��dU���ޢ���?.0?�	<>��O���h��d�/��9?��>�U��1��=��þ���J�=��/�ѽ~�Ua��m�3���9��-���R1�?�>�?\��J�`��"�F3��n ʾ��R?J4 ?3�?>�	?^H��脿��p:�>Qh�>��&?�\�>w[?~�X?�R?^$�>���aڧ��ۜ�hR3�U�?cg?)t�?�"�?$~?��f>^�=���=ˊھ�����<=�Ͻ��7�܅�=��g>%��>|ҭ>�D�>�4�rm����������>�@M>���>���>��>t>�un�
�P?�	?�7��H���n�E���yi�T\?;}�?�T%?�~R=���H�Ȥ߾���>	�?���?��=?�a�;��=c�9��ɾ�]��>�Ѧ>���>��f<m�=k>�Ė>=S>LĹ��
��B+���Ѽ�f	?��H?s�B>�g��-�B�'�X�:�@��>޾�	�;��f�5WH���>��
U���5�(;�G��=�f��V��������$�{��>~sI>��">-�$�a(=�)c����=��#���=�d�=�\�>��`=��z��H��|6���������D���'��˾lk}?I?��+?��C?�Gx>��>5��>[ǀ�)p?j�U>=/P�+v��n<��Ũ��$����ؾm׾�ic�2ʟ� 	>2yM���>�23>S�=��}<���=Q�r=,	�=��[�Z|=���=�V�=s~�=�y�=��>L�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?>ti��d�>M���㎽�q�=K����=2>s��=x�2�S��>��J>���K��A����4�?��@��??�ዿТϿ5a/>�%Z���0��zR�$[E��ʾ��>�5Q�~2?��7��������j�>�O��A�?���>���>m�?J���s����=6�>|�(>ԣ�={�{>U8�=��P=S���AJ=A�K=�0>%�=��>�n�<mZE���ӽk�=ā�=�[>��
?Xe2?�6?� |?G��>6U^������u��3�>�Rǹː?�Ғ>��0>O?_�?��?��\?�B?��>8��>S9�>�g<�*�x�����3.���=���?>��?A�>ܧL��;��'b���C���.��,?9�s?=2?�c?�R�Z��PT&�ϑ.�rR��������+=CSr� �U�=���ނ����o.�=^k�>���>��>!9y>��9>�N>r�>z�>�;�<f~�=����hy�<"?�����=y폼���<��ü�E���#�8�+����Ԍ;,��;G|[<�c�;���=[�>��!>�r�>���=vP���+>�����3O��{�=1֥�8?B��a�`kz�c70�g�:��1>>��Y>M�r������?u�H>�VJ>�)�?��s?�,>d����ϾJŜ�n�a�N:X�c�=�W>�#�t�5�v-[��I��ɾf��>�H>���>�:J>����B_��S�<%�ﾉ�G�>��>�����ѽ�y�Q�ద��?���~W�nj*�м0?-i����>z?d?��b?B�?���>n���l���b��=�^�bQ>g+��;��7���f?5�*?�?뢓��(�J̾O��L�>�<I���O�/Õ��0�0���з�h��>5����о#3��f��������B��Lr���>I�O?��?06b�{W��eRO�n��� ��}r?*}g?#�>aI?1@?�,��Qv�o��J��=��n?۲�?f<�?�	>r
>+���U�>��?x�?J��?][{?��2��>��=�?>��ܽ�ڟ=��=@�=&h>8�?��?%	?���������{޾�F���;�:F=4>�
x>�.>��=��<띀=6nk>r>(�y>6Qg>�܌>��>�Ӿ���C�7?�#=�5�>/
�>&��>�ᘽ�N6���>���=<y��	��"����6��:����.=��<�� ?�7¿���?�Z;>*����?�Ǿ~
S��&>�TV=�@��y��>2��=���> ѐ>�yN>�p�=�z>{�=#zҾ�->��(h!��C�/�Q�l�оn�{>����J<&�[���]��ӧG��z��s��?�i�5-���I=�qf�<�(�?�m��JSk�-�)�p����$?:�>��5?�Y��?��$�>(C�>n;�>�T���^������`ᾟ��?���?U<c>��>5�W?�?�1�3��uZ���u�(A��e��`�q፿����
����"�_?7�x?JyA?�Y�<:z>B��?�%��ӏ��)�>�/�';�x=<=�+�>�)����`���ӾS�þ�7��HF>n�o?1%�?tY?7SV��/�Q�$>��<?ý2?��u?�v7?�@@?�K��!?B>�;?�O	?7�4?g%+?�/?77>v�>�M�<�E=�ט��.���̽��ν�,�r�R=�h�= cX�_�<4�*=���<� ���!������gϼW��</�#=0��=D$�=� %?㹂?[�>ݯ>�W?󠾔@������?�?<g1<�\�X�~�kyҾ��4�?"o?�ݵ?4��?�lB?!�	Z��^r�>��>Jfo>��>�%�>Ę_= �ھ�Uy>B>����z�#>U�G�;i�X���ľ��_��wm}�t��>Say>�B���o >����9s�0�c>��L��6���IU�I4H��0�i�s��@�>�bK?ms?��=�y�f���Ue�dk)?�M<?DlL?tj~?�o�=�eݾ^9�� K�<!��Y�>gB�<L������D��G�:��5�:S�o>=G���<�ͽ}:��H��R���C8�cy��z\7>p�����=!i� ��%ǽuQ�=���>E֨���3�L����ԩ�*�e?q�=�O9�F�m�}-復$=>�Z?��?����2e�Piy��IW�+�E=Oa?"��<7U4>7���L����jF�>d�D?p�`?߅?gpz���k�S�B��-����������?;ۨ>��?�5K>�R�=� ��$�
��8b��$D�P��>�&�>:�ŗC�[q��sb��2%�iψ>i3?L�&>�?�NS?_�?�_^?�I,?zh?�ޕ>�Z��"տ��B'?�?��=�����R�r�9�"G���>�,?��?����>��?�?��$?��R?Ң?��>�A��a^?�Mڕ>�ȏ>x�Y�����*�a>¿I?Q��>��Y?MǄ?�k<>Q�3����;�Ž�/�=�W>�6?��"?��?Z�>���>��+��a>�xy>�K�?{�?aO~?�K
>;��>�)�>�u�=EV�=0C?v�>q?��=?�;y?�dF?��>����q;�MU?��@+� �f�5��!�p=rC=��\���&�}�"��o���v���=
7~=U����[���;�s������>��r>'���Rm0>�Bžp��Ac@>ߖ��5��l����9� G�=f�>��?Pڔ>�$�:�=|û>���>�����'?z7?�Z?��_;�b���ܾ��K�~�>��A?���=�/l��Z��ӽu�XNi=��m?�3^?��W�����h�b?)�]?xk�=��þ��b�p��u�O?y�
?��G���>��~?��q?���>}f��6n����Ab���j��ܶ=�n�>qU��d��<�>�7?+W�>	�b>�%�=?t۾t�w��l��]?��?T��?���?- *>Z�n��2�<��/~���CW?G�>ǀ��4?)����ȾV�������g ;�j���
������k"���6�g�s����s�=.�?[o?��o?��W?����`��yZ�:�����W�?!
�)G�:>��C��4O�j�Ǫ�d(�h��ZB�=R�n��)F��h�?&$?������?2���l�
�۾��>��w����0�=Z����<[��;R<(��t ��{��0?_�>)=�>y]?k�j��,�*27��U���۾�I�=���>�̱>^�>� ����N�Uiҽ�Ҿ�s���2�=�e>��h?�g?gwz?U�z�t���$����D�>1=#C����>�g�>�)>�@�Uƽ�&������h�{�	�?Cx�n4.���}�G4?�w�=���>{��?ɹ?M���]�ľ�j��Q�W���=1�[>���??@-x>�)"�6
�9��>�l?���>3�>�h��c!���{��˽���>���>���>��o>l�,��\��g��Ӄ��T�8���=�h?}��Ţ`��ۅ>L�Q?d�:|8G<�a�>�	v�в!�����'�O>�`?�<�=��;>�jž����{�5��X(?�?������+�F�l>D�?��>���>ن?�]�>�վ���`�?��d?�@?gG?)��> s]<]H�iٽt	�c�C=���>�~U>ob=��=��=�J��.��g=�=z?�`����_��,�5��<@;=9>����yx�����k0���w��{�ƾK������@Ľ����*�P�g��8���'>}�}�@M��>���m��i�?���?����3 =@������_��j�>-��8>@͓�5�.�Z�=o84��Z���!�7�h�����b��S$�> ¦��:̿�����,?��;?���?.�i�%��+[�*`�=�FB�8Bp�����V���:̿�ɾq�G?�>H?Z��oQ���>k9�>�޺=�Y>�ˣ��&��遾v�?�\�>\߁>?膾���26̿[��=#�?�8�?&yA?{�(�t��m'V=���> �	?|�?>�T1�G��ﰾ�J�>�;�?���?U`M=��W���	��}e?<<��F��4ݻ��=�X�=�z=���Q�J>�V�>Y���6A�\Cܽ&�4>�߅>��"�����^��ξ<�z]>�սB��4Մ?*{\��f���/��T��
U>��T?+�>�:�=��,?[7H�_}Ͽ�\��*a?�0�?���?�(?<ۿ��ؚ>��ܾ��M?]D6?���>�d&��t����=;6�و��{���&V�B��=X��>D�>Ƃ,�ߋ���O��I��h��=N	�Ͽ�L.�� 5�`&���<��u�n�����þ��u����ݓ��-3��>�V8><5>\L{>�gB>�=J>L�P?-�f?�"�>��>q������6��{	�I����R罼�e��C�|���1��(�ɾ�C�d����re߾)?���<2�U��1�'��NZ���A��+?�>��Ͼ��I��K���þ�{��
��Ad����ھ�4�P(n�m��?A�6?k�y��TR�"D�/�J�R���AX?��KS����Ҿ">�i��;�=�>�r>�,�2�1��}T�.74?�$?X�����HI>T��4=)#?	��>��=r��>yJ+?^)�]U��>�Mo>J]�>�?K>������7�}�'?^�^?%����쑾d�x>˰�H��û
=�&(>]�?�F�<�)�>*g	=c6��\��]�X�ǣ(=LW?7{�>�"����~��cu���ˁ=nRl?��>g�>��b?:�L?K%���H�U��$�<o�<�OU?�u?-�4>ӹ���K־�翾'2??+g?�
�>�LN�3�Ӿ''�M3���?զk?�m%?Ho����p� K������j??��v?�r^�is�������V��<�>�[�>���>��9�-l�>�>?�
#��G������ Y4�-Þ?��@���?��;<6!�Ǚ�=�;?�\�>��O��>ƾ{��>���d�q=�"�>����eev�����P,�^�8?���?��>����������=�r���ݪ?���?õO�\�]>Ep*����|?��S�= H�>�o�>��ݽZ��D5���7���{��X=хw>\@�^��T?.ľ�kտ�cʿs���xf�"C��"?��=�U~�u�g�g�+^���S�Ɠ?���v�Y��>�7>��ǽ*F����y�$7�OF��ɂ�>Y-����n>�Z�}p���P���<Ւ�>(z�>f}p>0��󽾔<�?����IʿfN�����x?X?'+�?�X�?��?k�
<Ä����k�[�XL?�5i?F]`?S�x�(�F��C�� ]u?d����6�@�(���$�vSQ>�t@?���>�4���>b�>�Y�>C;��XB,�~9̿Z���%�~ݖ?B�?����>��?�!?�hj���侕�]��=��Z?ua�=ת�V`��a������h�>��?����"�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�!N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?c�>��?�h�=�^�>X�=,�����-�fi#>	$�=�?���?b�M?)I�>�Z�=n�8�`/�#VF�IHR��#��C�Z�>��a?�L?0Ab>cG�� b2��
!�B�ͽ�m1�7�輬N@���,���߽�5>K�=>%>{�D���Ҿ��?Hp�4�ؿ�i�� p'��54?;��>�?����t����;_?Az�>�6��+���%���B�]��?�G�??�?��׾�R̼�>>�>�I�>��Խ����P�����7>(�B?V��D��h�o�u�>���?�@�ծ?]i��	?���P��Ua~����7�d��=��7?�0�#�z>���>��=�nv�޻��X�s����>�B�?�{�?��>!�l?��o�P�B�{�1=:M�>Ϝk?�s?dQo���m�B>��?!������L��f?�
@u@`�^?*3���b��,I�9��+^�=��r>{{D>%Ͻ���Β���ܩ�]�"��_=0[�>|s�>��B>�-+>��>�>�����X)��.���?���p�����J��H�����諭�+�Qi�
��Ӻ=>���Mǅ�P!v�.m�����=i�S?C3S?$er?t- ?�H<�7�>���P&=��0��Ώ=&��>��1?��I?#�)?��=�9��Xc�2��F����e��S��>��J>t�>���>���>��B<͛J>187>&�>U��=�f=���;�j�<�T>�>�>=%�>�4W�0뭾�Y���U��!���ڌ�<	o�>gL�?���E�������	����)���F>��?�dL>B�����ѿ�����B?^t6�e)��=�����>~k5?��Y?Aq2>I�7��5�����<[>�z���@�=�v�������(��>ǔ??�i	>�4�=�h\��A0�Q�îS��϶>̿:?�q��L�;�VT�)�y��߾�>;��=pl*�w�.�Ȫ����2��k�y�s=iU?j� ?2�=��;�D��v����>�L>t�>��!��n>���^�:����J>=�q=!+9>�t?k�->�l�=���>g5��u2a��>F�@>"]*>RY<?J�$?b-D�M��������/�9�t>���>�q>���=݉J�� �=:%�>��^>�P�Sp������.K�GF>���+P��s��]=��ǽ���=�P~=d����E�z�Y=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ~M�>�����G���み�zi��fU=��>o�=?���0��+<!���?'�>���J���ǿ��r��a�>5��?%�?V�i�����hH����>���?��o?J�j>mľWW�@X3>c>?�tQ?|��>�N��$���?e��?�χ?��1>���?� �?׊?w��=}��<i������{2�=Y/%�Y�?��>����%���2���f���{�-x�z�4>���;��?%�u�;�Ǿ�\>-�f�����!�=8zk>,�>�x=�܍>���>���>L[w>/⼊��<��1�K?���?����2n�kD�<��=��^�#'?�J4?υ[�K�Ͼ�Ѩ>`�\?�?B[?�f�>����=��-迿�~��ɵ�<:�K>I5�>�G�>@%���@K>Y�Ծ&5D��n�>4З>,���?ھ�.��O���?�>�e!?Q��>�Ү=f�?� ?�yY>���>W9:�����{B��9�>�e�>"�?�>�?��?��޾�M9��/��̠�8�Y�&�v>�c}?ZL%?_�Q>-���G6��H�G<�e�<�;�=�^w?%�L?�i����><��?9N5?)I?]F->�����ξ�<`-�>?+����E�d�J��p���.�>��a?�?�B&>��^�����Kپ�@4���?�ן>�q?r� �&�;��Z�G^=��_� �<�k=-$�=}ت=���=v���F>���>A��=ci��ܾ��9e=��z>�>\+�>�VC��8�E
/?���<�Ȃ�̛=��^��O�Њm>�J1>�P��-�e?҅1�Uf�F&����)%�s��?��?�h�?y}r��>f��C&?�?x�"?��>�֛���㾑)��q����ٌ��I��d�=��><��<��Ѿ�L���s����c���fK���>�g�>��?v	?��=��>�蒾�,�_G�?���6Z@����h5�4�D��y+�dpw�ͅ�����=�ܶ��v��=>�^ǽ�?7R6?�0>eNa>L��>!	/>���>tc�>�,,>�J�>���>i_>ţ�>z�P��u���FR?|���q�'���;���a/B?�sd?�3�>�h����V���~?z�?�r�?��u>+oh�m3+��h?=-�>����e
?W�:=����ʈ<dI��@��d!��3G�K��> �׽h:�A
M��=f��a
?8?�ߎ�}̾-a׽ۑ����=Mv?�.?Έ"��X�mk��kI���D�6�����q�ƾ��%���p��I����r��z�ӎ.��]+<x�)?J;�?�>��:�ܾ����@oC���9�k&A>~��>_��>��>��> �#��%B��X�+R/�3o̾�?�6�?�è>q�O?�??��M?_\t?�� >
�v>|3�����>�P�=��->��?�zx?a��>�T?�0?ԅM?E? U=�_�F����-?�L?�$?��1?���>�w��Vg�X �0��;ʦ����I>�=ڡ����C�ɽf�,�"�r=��1?�)ɽ]&�B2��=D>B?u�?�]�>ppO�����?�<��?]E�>a/>���!v�
���
�> �?ﾼ<\�<Q=>�=<h�<���<b�,>c���&���c=�`+�1º�m��=�h=��ý@R0=�]w��Ī<%��=�d�>^�?���>�8�>�@���� �����<�=	Y>I�R>�y>�;پ�~��"&���g�Y!y>Pd�?Ul�?\�f=���=�u�=�v��T4����ỽ�-�<B�?�=#?�ZT?���?��=?J#?��>`)�gV��X^��"|��\�?4(?O��>t����̾���d�/�@?�7?�_���!��b'��j;�|߽m�>v�/���~��G��#qC�^�;���۫���E�?�{�?�� ��6����m�������B?���>/b�>F`�>`o(�'Wf�s>���@>��>�sN?�>�~[?�(�?
�m?��>�C"��C��Ö��-�<���<Ы??�Y�?{(l?�:X?_q�>�G�;�,�e�߾!>ݾK����0���E�ȍ=^�>���>�>�>�w�>a�>;���Y��SQ �t]�=�>�p�>~�>�Y�>�P>�r�;x�e?V?�sɾ��ʾC�����~�$�+��?l&�?�?`@2>WI����)�;�B�j[?��?���?%}O?��{��4�=P=Ȭ �I� �3�	?"!>��>�ǳ����}�>�����>�.� ���e�di�⛃>�kU?��;>T	���YZ�����;�x�l�����3����6<��B��r���*�j���W;ܾ{B���忾��þ���V,ʾ[�0����>�/�=�o=nU=u��<��
�W�D�b�52�=�xý��ռ�#>���{R=,ۜ��x�<�և<�w�<7���L˾��|?͖H?�d+?�C?:-y>�>�h2��Ζ>�y��+r?DU>E�R�oF��<�^���#����ؾ��־D�b��1���8>�I� �>wQ3>_��=�_�<�=5 u=�J�=����5=���=�Ϲ=�֭=�]�=>��>�6w?X�������4Q��Z罤�:?�8�>d{�=��ƾq@?�>>�2������yb��-?���?�T�?>�??ti��d�>N���㎽�q�=H����=2>p��=y�2�S��>��J>���K��@����4�?��@��??�ዿТϿ6a/>���=�+�=X����ݟ�t��������{?�&
�!�v�>�Qs�>y��举($Ľ�S�<����������5��r�=hB��w�<��t</jz>7nP>7k%>쇞���)>�j�<�{�=ڳ�>�L"���*=�§�/�%>�)1<�r�>�޷=4t?�"?�5?�`�?�5�>���6���WZ���>�����?��3>���>���>n�^?�e2?N�?�1�>������>\�>��K�/�_�4��/���W�'�W�?̽�?���>��=�5۽@i4�z�L��ѱ=6�S?��V?)�&?�^>"V�
�࿽Y&�ʛ.����P��+=�mr�]U�����6m�E��'�=�r�>#��>��>FSy>�9>�N>~�>�>�5�< r�=�������<)��3��=Y����+�<Jgż�튺�q&���+�͇��m��;Dk�;p�]<:*�;�y�=h��>ir>���>��=Kz����.>x�����L��=M��*B�'�c��0~�&/��^6�,�B>`%X>�ك�r'���?��Y>��?>�m�?�+u?��>�+�=�վ^C���d�iS��ɸ=�W>;�<�ht;��7`���M�x9Ҿ���>l�>�?�}~>f괾񷆿��:7:��$X��h4?��h�=G�6i-�sh�����Ɣ��,c���>�m?��)�w>\�L?��H?M1�?o��=�5'�@p潒G�=;FC����=3�����=m�0=h_?���>)�(?��C�c�!�x̾:n��?Y�>�HH��O�pꕿ�0�T�%��H��4��>�Ȫ���о^�2��k��X���B���r�S6�>��O?���?�'a��j����N��h�/$��H�?	�g?���>�?oV?�ՠ� ��Q�~����=zVn?��?��?�;>KC`=�:���?rp?�ٙ?�U�?�3R?? @��D�>�e>��r>�=
Y>(5�=��R=�=p>?&�?<[?�C#�ɧ �o�����k���6>{��=C?�>�e>���>6e'>�A�< ��=��>ܔ�>��s>�n>�E>�>�o���>���,?~�=��>�Y=?y�N>�\�;�37�v��>8a>%o��A�����H佸���{�=ly=s�C;�>��ÿ�?�MC>���)?�J꾃/L���k=/4 >]����>5�=�;>��>�>��U>��>{x�=I&���L>C�����6��+K��'�AYQ>���˹Q����w?��
��E��	�b\��y���)��&9=)�?B��;�W�/"��oƽ�2?\��>�'?�x��d|<tX>/.?.I>���R[������,����?R�? :c>��>��W?џ?�1��3�dwZ���u�="A��e���`��ލ�=���B�
�X���_?��x?tA?�'�<B5z>Z��?Y�%��ɏ�'!�>�/�= ;�N�<=�+�>�0��(�`�4�Ӿr�þ�8�IF>-�o?�#�?gZ?;DV�ͷ����F>�N?�E?c�^?,`X?�Z?�)�<X(?m,�Td�>�u�>cI?ia?�H?FJ>�z>偍�/�=�Mj��,��x������1�Pyo=�O>�=�<4�=B/>O�;�.O��f>�읽M7*��Q
>�ܺ=Q�=�
�>iLo?|��>�ۛ>�?M?Ֆ�$\�/���v�>�>N����mV�H��=��Ӿ�e�>��m?�s�?��?<��>�:_�=ra���m>{8Y>�{2>;��>I�>����ꊾ,��=�K >m@�=�=U�<�����s�n�S�"�q<��J>�}�>�<\>���$�>b󔾩s��O%>�~����D�{N�m�(���H��놾�i�>��%?�b?V)�=���A>y���g�cd3?�AV?��G?��Z?�A����A�H�+d���X�?њ=磾����K��oGW��?�=�]�=oG������~#b>��S&߾�cn���I��;�ņS=���GD=,q���վ�+�����=5>��� � �l ��8W����I?�m=#���<P������>�[�>���>�>��z��A@��ǭ��z�=!$�>��:>Q8��9��G����$�>;	G?��{?ř�?����l���C;?�����ƃ��=S0?rA�>4?
�=��=S=H���ؾ�L�wX�1G�>?sQ$�!�2�䶜�������'�
��>Q��>�1>(�'?��F?��?�j�?ZY?�~+?���>)A�^��$?���?��= rw���Z���=�?�B��w�>��$?bx.�A��>��?L�?e�,?�tQ?k?��>�	��#LE�>q�>���>�Y��|��e�k>��D?�ʹ>VnZ?��~?�9:> a5�3��"8��>�1<>/?�?=�?�6�>���>�p��[�=�_�>�c?%�?��o?��=�?}�1>���>w�=,w�>$U�>y�?�EO?ٻs?��J?`x�>tی<�l���̶�a�t��E���;V�<<EDz=��qu���w�<'q�;Qո��9y�����bF����*��;�Y�>��s>/��q�0>dž�����DD>��\���W����=�s��=Z�~>if?���>��$��܋=8Z�>^��> u�y�(?�V?l?�ޭ��b��BܾиK� ��>�t@?���=��j��|���?u�
�t=S]l?�d\?<Q�E���!(X?�,?9���<��4��ZD�J����U?���>պ۾
�N>�Mm?2.?*�>�<����e��<��,�=��w���F?>]��=��'�[45���>�R?3B2?���=eH>����#a�P��?�$�?�|�?"X�?��3>Ѿt�E�Կ(����ݑ���]?�R�>sϦ�A"?V��F�ϾgF��o���W��������(T������$�����{�ؽ2"�=��?Ֆr?�6q?H`?Ξ ���c��]����Q'V�bB��'�j�E�$�D�\�C���m�g���<��*����J=/t��H��t�?z�1?��Up\>��?���4��'N�@�q�([��{���>��>�
t&>+ZT=(��%=��6���2?\��>`P ?�q?����J)K������8������>��?���>�d?�N��L3=���=(n��ܡ�a����pk>�la?Z�M?�Xk?$��0������!�e�ZU��\�8>V% >���>��X���"�H�#�ѡ:���n�������_���j=@�,?rAu>-[�>���?Z?yF	����(>���2�D� <�¹>
�l?Y��>{��>#���k����>/�i?�2�>�_�>���0' �S䀿��k��6�>���>LQ�>ZL�> D�{]��"���Ҏ���4���>��d?"����}�[Qv><I?�p�<5�t<E�>鵂����h�ng!���	>=��>�)�=m�>�Dƾ����;s�����e�)?��
?`����+�o�>�;"?�*�>J��>r�?�N�>}�Ǿ�'0���?�y]?�2H?��??���>�=����Ƚ�'���;=12�>KU>��a=��=�����[��?�~�R=�r�=�mԼ������v<�ָ�la<*��<f�/>�_ԿBwZ�&��n�]��4#��/��)��*6=}���%l7�a�T�g܇��8e��(���ѽ
n��T���|�l�����?�1@�W��;���z���"�� ����?lH���sY�$?��|�&ᾆ�ݾD�R�����z�]�|��s�r�'?T���ǿG���5�,�*?��?��j?Ψ�R��?o=�pM�=k�<�Q���h"��`Xο-���ֵe?���>���W���(�>^��>�Fn>f)f>},��=��Ga=� ?/�"?%� ?�`p�p�ÿ�M����<e��?��@�rA?��(���쾠�T=��>��	?+@>ƽ0�,@����
��>�"�?�܊?+qL=��W��0�6e?�C�;q�F�Ԟֻ6�=�1�=.�=����'K>Ȧ�>�����@�d5ܽ�m4>�Q�>�m!�����]���<q]>wֽ�����!�?�@�dM��kH��Ht��f�>߳W?Eo�>	�">>?f%��ſ�&����?:��?�}�?�?���S=����yA3?	J?�>�$b�l����
>"/��B�;��3:��b��r��>��S>t-Q��	��	��iĽ��;�]��pǿ��#�� �q��<��]��\��������CN��2���sk�<aڽ��l=�b�=�'R>�Y�><<X>z<X>l Y?��k?�
�>��>������*:˾�uֺ����vz����<��C>��U�63�:�	�9I�����R˾u=���=]*R�N���0$�if�D�E��H/?� >�vӾ��N�k2:rо�����橽��̾ap4���o��|�?��H?�H��wiF�3Y	�8�S���_Q?��Ģ��,��:��=����io �8�>�sK=p�����<��+K�ƅ?��?Yp����>ط>白=�4�`�6?YԷ>{�<�T?��q?�誾�F��7��>=��M³<i�<?9�P>:�xmw�X�?��X?�>+�J�Ͼ�3��~�x���Ҿp6_>�Qf>��h=`��rf��j�=������=�9<�Bֽ��E?5�>d������a���_>��GA�kht?�z?i��=�yY?L4K?��HI��F���%��-<�7�P?-�f?��>U�0��8쾭\����1?�0[?�> n}�Yo澅0����Mt�>:]?�� ?�Ký��j�����?�	�\�+?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������Z�=~'��U��?:�?z���><�����l�����"��<���=9����S�Ov7�;7ƾ�g
�.����Ѽ���>\@@)��g	�>��;���Z*Ͽܹ����оA�m���?�ϫ>g��ލ��Ek���s���F��I�붍�ݿ>�E>�`�������P��������?���7��={xJ�ϟ��Қ���q=��8>���>�IM>W�2=8����;�?���^ſ G������@�g?΃�?}�s?�(?Ȥ��	|���ľ�
>��p?5=m?�tn?zT'�M獾<J��d?�^ؾY�v��g,��wC���>��?�Y>�<��`k>R�T>�Y>�'�=̛C���̿�����!�2�?C��?Eq뾪5?^
�?�w?
\�j7��⠋��$�0��=�?��>�3Ӿz�� ������?��(?��"���^�_?(�a�L�p���-�x�ƽ�ۡ>��0��e\��M�����Xe����@y����?M^�?i�?ҵ�� #�_6%?�>c����8Ǿ��<���>�(�>
*N>�H_���u>����:��h	>���?�~�?Oj?���������U>�}?���>D��?�=��>��=���@�Ҽ�)>���=GK!�M#?J�O?�>�=Y�3��</���D���N���\�C���>Tka?�K?�va>�����P�����G̽�+�;1��<��8-��۽�+>T�:>.�>�B���ҾL�?�o��ؿ�h��Gx'�)54?ֹ�>��?w��:�t��3�=8_?�y�>�7��,���%���N�+��?G�?�?ý׾��̼�>P�>�M�>/�ԽN��-|����7>�B?���C����o��>���?ǵ@�Ү?�i��	?���P��Ua~����7�e��=��7?�0��z>���>��=�nv�ݻ��W�s����>�B�?�{�?��>!�l?��o�Q�B���1=7M�>Μk?�s?�Ro���e�B>��?$������L��f?�
@~u@]�^?*hֿ���K��ė�����=���==�2>�ڽ�d�=1�7=P�8��O�����=O�>R�d>�q>�(O>na;>s�)>O����!��q��Q���R�C�-��~�d�Z�J���`v�{��4�������<���&ý ����	Q��+&��8`�J?�=4�N?�ba?��p?]^?�D_��M�=��
�y�=)���	A=�&>Y)5?N]??��?�v>{�k���^��Ղ� �ɾ�%��f�>9�=S��>y�>^>�������>@�/>�h�>�x:>�^�<*�@��
� W�=4�>���>�j�>�>j�0>�Y��0��b%j��%����lP�?�L��h�R��ɕ����� ˾�6<�=!?��=�R���rѿ:ת��?G?�.f��^
��Q��>>�#?j�F?�>׼پ-�.�U�8>'�!�E�r�ج�;ܯ���_��Q�>��>E�.?hh�>e9>S_3�aq���M�3�E���>�SJ?�Sľo���h���t:�l�����>���>�V�:(��䗿L�N��	���>�_>?m��>�<u������q���/����>�G=�y�=��'=��v>k��Ŷ�=G_G������4p>�G>g��>y><>2�>=?|�����\o>�*>���= WI?��2?4�<��A�|�F�A�p�xV�>�>���>�Ҫ=���"��=y�>~8>�Jƽݍ��֛T��d)��u%>%����O��-���=�Y����=��=�,�<
�K��fx<�~?���(䈿��e���lD?S+?` �=�F<��"�E ���H��G�?r�@m�?��	��V�?�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿg��>��l�O���$zV�����7">�ޠ>��W?��b� xD��<��cW�>��P>�w�y`��tHɿ{����/�=W��?��?1���@���}A'�|��>�2�?%AV?+>��3R����fp���Y�>+?u>�>��4�l���`?+)c?2�E?P�K>�+�?Ugm?��>���y�-�
{������WX)=O�=΋�>��<>D�ʾ�J�n䊿����Gd�V�
��gb>�Z�<h�>2�Ͻ�cƾ݅=q?���D��ļ���>?�f>Ӈ4>�>D0 ?�D�>؝�>��<�a�b���5W��L?,��? ���Pn����<�E�=��]�.?�J4?�uW�q�Ͼ�e�>�\?�ʀ?�-[?ܔ>í��8���ܿ�G����<��K>���>"��>`����K>�>վkD�~Ί>���>I:����پ�Ձ��(���m�>
>!?���>���=��?q�?$�N>�rk>�!�&�|�4�s����>���>a�0?�@z?�I?)�.8��և��I���A�v�>�_?$�2?R��=�Ӓ��}��r���	K7>�J�=ta?&I?�N���S�>w�t?�6�>':?�b>{�D�%���hϽ<N>�0?�H�;H�{&�r3˼�=?D�9?k��>���<�W�u�6���	�߳���'?�:'?�
?2�込E\�bΓ�#���1	�J���0B�< Ͻ��>�-�>��{���{=���>s/:<4�㾫����=HM>֑?)8�=�P���C��*=,?F�G�mۃ��=y�r�;xD�u�>�IL>����^?0l=���{�����x���U�� �?���?Vk�?[��=�h��$=?�?H	?i"�>�J��~޾0�ྯPw�)~x��w�p�>���>�l���E���ϙ���F��F�Ž`��z�><�>2f
?܉?�QL>���>j��^2�rƱ�BJ���e�~"־Y�'���+� ��5����B�����*�e��Ak�>��޽e�>{�?�+><2!>3?�[[=5�g>t�">{eM>A�>�xz=t�>�q>Gg'��	���W?�L����#�%F���z��O?p�W?>`?��;R���F �*�?[�y?
�?���>��Q���!��>���>h�\�#�>oI-<\P�L.M=CQ��5��mm����r&�>�a����]��� �uU�
�&?#b;?�[�$���XB�F ���b=$��?W#?+�)���P�4:j�;�R��T������`k�~š�<�|�p��4���v���+���;&��x�=t�(?֞�?m;��Ta��b�e�z0?�]g>���>�H�>���>6f>�����3�kW��)���~����>hx?��2>��\?]bN?�6{? �]?�m&<��=���
�*?׋[=GV�>�#�>+?�O?؝A?�e?�w?v�>�Ѭ��\��*˾b�?d!?(?�(?��>~��e�=d������둾��>��=}~Z=U��E����=^�+>QA!?�g��w&V�xs�K��=��\?��Q?}E8>�d���3�<���ŏ�=E��>��>n�*��;�c��=}<���l?�+V���n<�^�>�mn<���=�x�<��M��=mA=`)O>d�[>�Z2>G�����R�N>����l<B/j>�G=B��>b4?�΍>N��>�Lv�H`�-��
�=
�S>~�i>�->,Dþ����S���Td�w�e>C�?v2�?z�d=��=���=3[��5¾���b�����<t ?�!?�P?�ۑ?�;?�?~�=�B��⑿(��r䜾�k?�?<��>���fKվR+���n���?��?U�i�����6dV����9��=l��=iM�:uv�Xw����9�ڡ>q$�[�!�[x�?��?E��<~�G�o�ɾ���ʟľTX>?r�>���>���>i�K�k�>��� >�?�>5?	��>�HU?O�?q�?�p>�^Q�����b����,<�Us>��[?'1U?}1�?�0�?�E�>��>k����G��t�,�N͏�B�h�Jiþ ��ҏ>1u>��>M��>~�>>J��L���탾��<Ј>�U�>��>F}�>�1�>��r=��E?ʲ�>²���	��'������V91���r?^А?9�*?�-=��B�D��E�����> �?�$�?�,?�Y��+�=2��h���l����>`A�>) �>�\�=�P8=d�>�)�>�.�>�����6�I��?�bC?�t�=��ſiqq���p������a<�-��q�c� ���5[�-�=b���-D�Mǩ��r[�@������µ��	��R�z��q�>�(�=���=��=�^�<%Dм��<�L=��<0=� s��Ko<j�9�p�ܻ�:����R��'\<�$J=�� ��̾"�{?�lK?H�*?e]D??�v>)�
>OBd�D�>�zS���?4�O>Z;9��A��3D��e��k����ؾ*#پ;Xj�Oȡ� �>�$���>��%>{��=?e<���=��=X�=զ�4K*=OL�=�=��=�T�=��>}6>�6w?�������5Q�/S�H�:?�8�>���=�ƾ�@?��>>B2��_����`�.?��?cT�?��?�ui�'d�>a���䎽6q�=f���m>2>��=��2�y��>�J>$��`K���x���3�?��@џ??vዿ�Ͽ]/>dZ8>o�>sQ�o�0�
[��"b�2�\�F�!?�l9�[)ξ종>q�=��ྚVȾ�"=�G->�~N=�Q�Q[Y�c��= 憽��1=V�T=R��>�C>_�=����3�=ec8=� �=L�T>	|	�eN�ފ<�xp=B��=��a>Fj'>G�>�L(?k�R?N�?�š>�V�󊊾���c~�>�j�>L�?��`��u�>��>�K?�!s?撃?p�?N����.�>Dt>Ѵf���o���b�oi9��:>*0�?��h?��T>v�ƽ�'=ÃN��5��{$���?h�K?�1?�
?�!��z�5<Ⱦr[7���z��<l騼�վ����YN�/��=�޻��E>6!>���>�	�>q0�>_�b>�>���>:*>r#4�E�ռ�#���ޜ<��=E@O>��A>i):>�u�=��=�
��"	����!ͤ��}��C�=���= ��>{[5>(�>��=`.���;->z>���]J�{ɼ=\奄��B���X��ny�X�&������.>�:S>����M��{V?�mi>c�J>W��?N�w?��#>w۽g˾�J��_|p��b�A��=VD�=S=p�M53���]���F���ɾ���>�>H>�
>��=P�>��B���=����f�>����>�ڦ��g~�Q��;�g�Y��Q����r��0����^?�։�?�>��?ߘ%?tee?\�>�Q =E�K��4>s���"�W���־��4���=C�?F�1?�?������=�s�ʾi����Z�>�K���O�7&���E/�;�E%���%�>�d��[о��0�/\��}���B�:w��R�>-�P?\S�?�9f�񐁿��N��+�66�$�?&�f?(ؠ>�?�?���X�S#��9I�=�	l?u��?f��?�	>�ɲ=�䥽���>�(?���?m�?Wn?ۭI�QW�>�c�:�">E����5�=��>�W�='��=ǅ?��	? ?ܹ��vJ
���f	���'d�m��<�`�=0/�>~n�>[
Y>F��=�|R=�P�=$�[>#�>@ǉ>��]>&]�>n?�>Wo���|����7?^�=t�>�?��M>��߼"\4;l����C�OA���~罯~��"佚�=���<9Y�=͙�b6�>�����@�?�2>�Y� ��>�����J����1>�4=p�f�z��>�p>��`>��>��]>r��=cϣ>�8>�%þps�>�"��|	�^��x��T��}&�>�F��|���A����X�N�׾`#(�Sپc�q�]"��b�r����="�?X�a��(o��U���1�8?��>b�6?��6���'=d��>~r?�i_>U�ݾC������m�)���t?�b@� b>]�>��W?\?zn0�un3�?\Z��u�b�@��e�!�`�aԍ��Y���x
�)�����_?�x?EPA?��<k�y>HA�?�%�����>f+/��{:��6<=#��>��]�b���Ӿ��þ��C
I>�n?;ڃ?L�?��U��%m�n'>%�:?��1?&Ht?��1?֜;?!����$?�>3>�,?+f?�K5?��.?w�
?[2>���=�窻}(=�(��H����ѽ٠ʽ,�#�3=�;{=R'��S
<u-=C�<׊�ڼ¢;�Q��͘�<sc:=��=�/�=FU>'�c?��>���>�A�?��{�#�R��ؾ�i?e���
;�#;C=OH�i���Y��>��f?擲?��|?�3>�q�����Y��=��T=�>>U(e>vN�=��!�P'���<�+>�����'���G�ھ�PC��0>3��>���>ѧ�>��a=��'>	-Ѿ&A��܆>Ե���v����P
&��1����fP�>�E?V�?��I=%���c�J���$�#?Wrd?!]X?E��?�s��_%�A�2�i[.�5{����>�/r>���1d�����J�E�T���7�?Qi̼�����f>�}
���ܾ(Yl���J�Bv���G=�P�P�R=�(��YԾG)}�Q�=K>t��c_ �����|���YK?�Jx="b���'W�%��0[>7�>� �>YlG�/����>�=\���`�=k��>�5>#Jɼ�'򾋤D����*^m>�o??$�?���?����d����K�ܖ)��5����=<u;?��E>R�?��>�� >�,#�}�߾5+v��\�Y��>Q��>���d$��2��$��9���q�>Α�>�9N>0+?E5?��?�i�?�/?|?{Z�>J
ٽ�۾��?�F�?P�= ���pսt�>�K	h����>n�&?wI
��({>=|?�?��?aB4?I�?c>����=���>6o>�ub��Ʒ���>jY?���>�yZ?�	h?֕=6?��u��m���x>D��=x ?���>Q1?ʝ�>C��>s���0�~=g�>L�b?�-�?H�o?t��=�?��/>�;�>���=�C�>9
�>�A?�8O?8js?ĬJ?���>���<�ȯ��1��c�u��H��s�;n*P<�]{=�4���z��?���<�{Y;q�����c����9A�ҡ��2N�;1d�>J�l>����j'>��žJ���M>����OP��������7�g
�=��x>y� ?�t�>�y&���=��>4��>'���7&?�?t�?��;kb_�&�־�J���>��B?1��=�qp��ے�ks�^W�=h�o?h^?��p����q�b?��\?���X�<�jž�^�t��o�O?hO
?�FH�S��>t8?T8q?	�>��e�Mn�Ȝ��la�5~f�i��=@��>n���Ud�[�>7�7?u��>�Tc>��=+ھ^w������>?@��?cɯ?�;�?q|,>�io���߿�����ӏ�|�e?���>Y~�)r?�{9�V羰;R��;��tr྘>��h:����돾�G �v�R��ģ��)8=8�?xn?I�?F�d?sJ���h�bLT�x��L�\��������	C�FSJ��I?�)�v����,��
���'�<�ϝ���%��
�?��C?��켬��>�=��5�G��z��Y= �w�^�����+���Ŝ>��A>9sl�V�q����)?\��>��+?��j?����z�a�~w#��L��H5��>e?�H>���>�&5=<,���S8�Q����뾠Tg� �u>Ptc?rNK?�En?�>���1��Â���!�n2������*B>��>Nz�>T�W�G��~%�D�=��s����j����	�Π�=�3?"r�>�ڛ>4ɗ?�H?s}�������s�ֶ0���|<N�>�]h?��>��>�ѽ�Y ����>��e?�5�>VR�>:�����Lfr��:���t�>���>nE�>�k>�>��E^��{�������=���>��k?|3���WS��{>f*S?e�̼�z:1�> =k����$n����*Sj>��?zc=��W>�`þk����s�����p)?�F?M`��M*�*��>�p"?A��>���><̃?[�>��¾Ta:u?�R_?l�J?�@?��>�=����ý3*�!�-=��>�Y>l=��=:�/Y[�y#�l[=��=���r1��T.k<X���_�b<п�<�1>�翑�>��[����T����b����fӽ=�w�\ǽ��Ծ�����Q���d��� K?��*A��9Ӿ�����l�?�7 @��x�U�L�B��s�u�`���i�>q�*��{N��I��x潈���C�	�|�l��6��R��}qx�ч��5�)?���fhǿ�"���Zپ��'?4�?�q?���d��8��k>
V=��u�rJ�������>οqJ����c?ܔ�>�P�g��b��>��>�%M>b,^>�9��N����N<�/ ?C�*?�4�>��c��[ƿx�����b<��?Q#@�{A?��(������S=C?�>*�	?��@>��0�4��԰�]1�>�5�?��?��M=��W����a3e?Y�<�F���ػ��=c�=g�=oU���J>�R�>�^��'B��'۽ 4>�!�>*o#��]�	�]�s��<\�]>��׽���Ԅ?jo\�f�`�/�vD��{>��T?k:�>℡=Ί,?�H�zqϿ��\�_Ba?�#�?���?��(?<꿾���>��ܾ\}M?�W6?�&�>�q&���t����==�弅��I{�V��!�=���>g
>Κ,�Vk���O����z8�=E���п���9�[<�yK�����/�c�ܽ"�P녾����	��Ҧ;g˨=��;>��>��>!B>�bY?��w?ĩ�>�n>��Q��L������<��X�1���%2�a~�������ߍ��u�.F+��<Ͼ��E�<�=��C�D�������g��!_� -$?`N>��㾮.A���ļ��}%ݾ� �J�Ͻ�SվG�=���r��b�?�&F?���J�>�]V�����.�w�Q?���/����|��=�6�Q4�=&Ό>sƻ���č!��pQ��//?56?�غ��?����I>3}����7=^.?���>����>��?�){�Y<���u>��=>1;�>�>ߤ�=d������!?Z�N?� !�C��ց�>�~�Pׅ��w>�3>͹W����x>��<�!�'��{˫�O��<ɫU?ᒊ>q3*����_���3�Xv=w?Ù?�6�>�h?t�G?���<���&�T��o��12=	�Y?�gj?O�>u�����̾]�����.?##e?Z�a>�t\�Ď�R/�S-��w?Otk?+U?��b<��v��㏿(�P�3?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=暕�ߑ�?�-�?�j��9Q<]��Ʒl�������<su�=t� �b�$��~���7�4ƾ�b
���̷м�.�>L<@c��Gf�>I5=��%⿄'ϿE����|Ѿ�n�a�?�(�>)��������j�^jt�b�G��7I�*���]�>��[>p�̽���,�8��9�:.(��]�>��H=Ik�>����)�#�!sľ��>�nb>d��>1�3>����p�ҾF��?P�TĿ�Z���e��{?�?��?�?qzϾZ|>�1����bR?�S�?�Z,?u	��ֽ�坼�^?0���b�`6M��L��2�>�DD?ENc>Ie.�_��=�V���Ț>>ګ>�� ��пӲ�����)�?'��?�e�~�*?.��?p�?bE�_�����ľ.��pܻ�t�>�̷>�(����b��'C�w�	����=`��>��:�54�]�_?$�a�J�p���-�`�ƽ�ۡ>��0��e\�'M��9���Xe���Ay����?J^�?f�?ص�� #�]6%?"�>r����8Ǿv�<���>�(�>#*N>H_���u>����:��h	>���?�~�?]j?���������U>�}?Fɶ>��?L��=���>'��=���gf�:X">�#�=W�,�x?hYM?���>�b�=U8�*i.���E�WR��(�p�C����>K�a?J�L?Z#c>�w��Ċ:��F!���ǽ�r/��ȼ[->��/�Y`ڽެ3>^�?>�[>>mE��EҾ	?�h��ؿe���0���4?�L�>\�?�	�Ȅv��a
�?�`?G�>,��갳��y��-���O�?� �?��?��׾f<Ӽ�:>��>Q�>��ӽZf��P��R5>QB?64�ҡ����l��|�>�?�8@���?C�h��	?���P��Va~����7�f��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?YQo���i�B>��?"������L��f?�
@u@`�^?*,b�溿%���7g��UY�=��.�4�= ����)M�+��=a���\�8<���=J�x>갉>�ą>�t�>�	e>�>�5��*�*�-z���ސ��m2���"�.������4�@�)�J}�H��ŵ׾�sܽ0����R�Lp��=��GH�<�=��W?�-s?LÍ?���>�q�Q�.=�K�V(�;�͓=L$�>��Y=R�0?�`?�<?�'�>D/���kZ�W܂��ʴ��}h�Xŏ>a�>C�>�ڽ>/�>���<V�z>�͘=3)�>c">�?k=J"�<���շS>�X�>.�>�r�>C<>��>tδ�1����h�bw�� ̽� �?�~���J�1��8��B���i�=b.?K|>N���=п����3H?���u*�2�+�s�>��0?GcW?��>a����T��?>���M�j��c>�$ ���l��)�#Q>�k?1�>��>!Q�d�'�Js��K��n,�=2)?�\����=�섿7����4y ����>:5�<�b�s܋�ΤY�+%�����=�t/?�?�l=@����(�9wʾ�?s>o#�>̡�=	>��2>����:�e����=m�=�ܩ=t�?��1>���=���>|��f
Q�)i�>��O>��>��??�b?{O�9�����[!��jr>XQ�>�p>HG�=7	K�+��=R�>>_>1Cͼ���p,H�\�P>Ά?��IT�xn��\=#�����= �=m��&�:���<�~?���4䈿f�d��2mD?�+?]��=��F<�"�\ ��BH��\�?<�@_l�?�	���V���?A�?��7��=_}�>�֫>�ξ9�L��?]�Ž�Ƣ�C�	��*#�S�?a�?�/�#ʋ�/l�h7>�^%?��Ӿ��>�k��~��X�����Ł$>���>�R?h�H��$��${�D�?�?��~�DRʿ���rӥ>e��?9��?�M}��&n�}J�iK�>�<�?��?�'�z�¾�>��>�p?q<?h>?D�
�R�,�v��><2Z?4h�?�5A>���?#Qp?��>�W��%�0�JP���_�����=Ѻi=�S�>c	>�Ǿ��A�k@��#����d��5��P>"�=���>��Ͻ�ʭ����=|��/�����o�\*�>Y�i>0KU>���>d0�>3+�>{=�>��=Va���v�^ ����K?N��?8���n�Zb�<�(�=_q_��?a4?�~J���Ͼ�ʨ>4�\?`��?��Z?My�>��_:��Oۿ������t�<�L>�p�>{b�>�Z���J>$2վ�yC����>�H�>����[Hھ-ʁ�Kϫ�^��>po!?�I�>��=#?
�?��9>��>��L�|����R9��,�>�ݽ>��?��q?4y?H1���D7�����ܥ�ϓ_���x>��|?B?*��>�뉿����g�k&�㍬��;�?%�g?��%��?���?�=?�7?( �>PL
�KȾ|(���@>p�,?���(����)��<;?�?^$?ͳ��wWa��`��?ɾ��.�ܞ?,�Q?"��>߈���jS�,蚾_��<t_X��]=�?�V�g;�LQ=�Ց=��Ux!�7��=�=%h������i#=���=U	�>��>�8ѾqI�-=,?'�G�tۃ���=��r�>xD���>�IL>����^?Ql=��{�����x��	U� �?���?Vk�?y��@�h��$=?�?V	?u"�>�J���}޾B�ྼPw�~x��w�T�>���>Ťl���G���ؙ���F��g�Ž�:E�E_?���>��?2�?���>+�>��ʾF{��l���(��{����W;�5�2��
��!��F���=ľop�a&��b@��d>��Iq�>�!?;M>D!g>t�?7�z=Ii2=���=��?�H>'`�=��)>u��>0f�:"��*0L?��þ�N,�P�������S?Dv?N�?u<�<��h����+(Y?��^?$C{?��=�cp�X%���>�V#?B��H��>���;b����d>����P�r�=
�¾7:�>��@X~���A�YJ����?h�R?֦>�Z0�����㠾�Gq=+�?��(?��)���Q��p�Z�W�7�R�}��)h�z���4�$�y�p��ˏ��O������(�u2&=a�*?��?���D�',��T k�??���f>���>d
�>H"�>�$I>�	�b�1���]�+g'�@2���X�>F.{?l�e>�kP?A�N?��j?Ղ<?�+>
%�>�\Ծ�T�>Z։=m9�>�@�>0�=?ϧ<?D?x�%?\�B?��W>B�M��G�?fɾ�u?��?��?@q ?M(�>~����N���.����e��z���Z�=^`��ѽJ�E�9t�<�҄>O�&?���E�C��,�ϝ��C -?I?$?S[������2�1?�-�>�<�>b�@�m�e�z2�i��>�	?#<���4�<�%+>g*�=���=�Q�;��Q�,ov>)4ɽCQ��>;>x�V>��]�6	�y`1=9e<G��>J����t�>��?퐊>�@�>`B��� ���Me�=Y>k S>>TDپ�}���$��%�g��Ry>	v�?jz�?��f=0�=1��=�|���Q�����9������<��?�I#?�UT?w��?U�=?i#?��>)��L���]�������?' -?7N�>�s��Kʾ�X��ur0��>?�?j�\�����O$��Gž�� ��">�(*���w�୿�_C�n�/����3��b{�?�?��|�ߕ:��z�m������0sF?p1�>��>K��>�*.�$�d�^D�I�>Y��>\P?��>�O?`L�?�)�?�Pe=��m���� ��)����^�>�l?f�$?���?�?,�?Tc�>��==wKﾄn0��{��*"n�ӯ���0�=Ħo>z~�>���>��>8_�=�Z�hJ��	7�:m�>��?>�s>��	?q��>c�=��F?�#�>�j���J�mע��f���k@�!�t?O��?I)?��!=���GE��_���&�>�x�?|��?��+?�'V����=�˼���O|�d{�>}��>�(�>2/�=E4P=u�>��>�=�>�X�����B7�X-@�T}?!�E?L8�=�ſ�Yq�I�p��ח�am<?���e�����z�[����=���ݡ�lԩ��V\�^���N��w޵��М�c�{�=��>��=��=���=h��<�7̼d?�<��I=�t�<zm=�Mq��o<��8�2�ݻ@v��v���AX<�.J=�R�až�{?	ED?�"*?�I?K7>�=V��"�>B�k=�t?�Dw>7ȽP�����/�8����U������׾YTX���8�>>y<�0��="��=��=���<�u>�f8=��=�m =4{=��=��L=q`�=��>;>��
>�6w?,���첝��4Q��X�ȶ:?�8�>}�=��ƾ�@?��>>j2�������a��-?I��?�T�?.�?�ti��d�>����䎽Cp�=.���}>2>��=>�2�c��>c�J>���J��f���e4�?��@<�??�ዿ��Ͽ�`/>�d>��0>�=���)��{ؽ0(o������0?C�A�Q����^=`ra=������御�=��>�:�<O�?�(�=�|��ة�=w��<��>�)>*}p��6���0=���={�=��1>�fҼ����0������=��l�k>m�(=���>h�4?�	M?S�?m~>A���U��S�����>�/a��	?lv㽤��>(��>�D?�]e?���?���>�����<�>��>�a{�Ƒ����9��㾽�W�?���?J����-�T�6>e�*�]Zf�	���C��>�W?�[??sƸ>���W��Q�#���(��Z����.����;��V��`o�����F9����0��=� �>��>��>�P�>�n>�P>���>s�=�l=�c�<��L:u��<ʰE�	�=c|��� �;�@��Ș�E9��_�ϼ�C�鎈��S=x�<�=l�=|��>��Z>���>/�>�צ��0>��ž�4=��!�=��>��7O� ���q�Dp��ε�W7�=b�=F��iA��ٚ?c6>�''>�п?��?�)>��˽�����Ֆ�_7�����}�=L�\=�7����>��$L��yO�n�Ѿ��>�>�>� j>�+���>�өm=mᾐ�5��{�>��������;q��������O�h�����MED?7�����=Ɉ}?��I?�q�?�[�>u�����׾�62>����.�$=5�%�q�&ɑ���?O�&?f��>��&D��:̾��q̷>=VI�� P�w�����0��K��ַ���>=�����о-$3��g������@�B�Ymr�Q �>�O?�?�/b��T���GO����C3��Wr?�g?��>@?F?�a��2r��x�����=�n?���?<7�?��
>䠕=Tl��!��>h?e��?�?�}l?�ZP����>�L����>�!�V��=%��=y��=�?>�:	?��?���>@������6�C�羢�A�¨�<��=J�>��>��J>o˫=A�=ٍ�=R>s��>�.�>S.�>���>� }>>ؾ>��bj,?x&>0�?cF?�pM>y���R>��R<�s+��
;4����탾̉_=�a@>�ַ=��Q�W0M��$�>�Ŀ1E�?GT�>ԝ�����>���낼Q��>�ش<,J\���?u�F>V�+>7��>X;_>p;�>��?� �=��ܾ�Q~>���*���UN���z�3����>\J������̼�� 7�茩�uk����Lng��J��X�0�� w����?�{�9ˆ�]��a	����>K(?��M?�p̾�ty<�g!>�?'n�>���%z�����������?k�@�4c>��>�W?��?�x1�]3�$xZ�Ӫu�$$A� �d�y�`�jލ�g�����
��쿽��_?��x?|sA?�Ǒ<-z>���?��%��ɏ�:3�>�/�.*;�U�;=�3�>���}�`���Ӿv�þ�&��>F>�o?H$�?TT?iKV�Rm��7'>(�:?�1?�Nt?��1?N~;?4m���$?&�3>s6?�k?gC5?��.?I�
?�2>� �=S��0�'=Q6��@銾�ѽ�ʽ���q4=��z=.�t�!a
<��=C�<��Lۼ�U";���y��<�9=(��=���=�>��?�K�>�~�>K�?�A�<];�s����?q/���������G	���&��u�>�x?D=�?�p?̷�JQI���22>�ٞ=^��>c�>�8>�|ľ�d=��>#3&�� >ȑu=�9P>�>���N���O��(<�{p>�g�>��;>"=m�H>�hn��!��t,�>�w���W����4��z̾AzD��I���`�>�{P?=�/?�_��&�����@w�^�%?��r?��?7cc?L8��Ͼe��EKC����<ޖ�>X��p>�|ݱ�����^�v V����=�����d�m>���9�۾)�b��E�����7=�	�'@=�}
�X�þ����}:�=��>䍹�
	��_��)��K�L?� �<�Q����i�e7¾�i9>�(�>+l�>h��t]߽��<��칾]h�=�N�>�S>�p�;�:�)�D�?��xs>��D?��{?{��?�p���~�?K����d����ԝ=��8?��z>�z?5�1>���=��?��ھ�S�h&d�&?�>%��>�'�;�A��I���������O�>��h>�$�>�$?�[?��/?�sw??�?�c�>0�J��P�#?��?�݋=9˽�qF�9�C�I����>��&?v�0��՘>�?��?�#?'�O?[�?��>����>�ٙ>p��>�Z�_��r�V>!�H?���>�mY?X)�?�>T�6�1���P�����=_f>�d-?�!?tq?gI�>��>�ڟ�9�}=�y�>�Yb?�ۂ?L�o?Ɛ�=��?{1>%�>U`�=G	�>���>�B?�[N?��r?�8I?rE�>o�</����𵽎�s�L�j����:��-<Pu=k���vz�H�N��<Lː;a˪�/�x��K켦\E�m���H;�x�>��s>����:0>��ľ+�� ^@>���P��pw���,:�Nٹ=�8�>��?���>��#�B	�=���>%G�>����(?��?�?�qe;�Sb��۾h�K�Z�>��A?s_�=d�l�7P��A�u�{j=P�m?�L^?o�W��?����b?�b]?�`�m�<��þ��`�Z<�ɗO?�
?dI�K�>�i~?E�p?u<�>�c�A�m������a�9�j��=u��>'�A@d��Y�>�,8?�
�>��c>\a�=7۾w�����-)?�ʌ?�ܯ?�=�?;�*>&�n���߿�� ����4_?��>�����$?���ѾH}�������羻���|���w�����eN�����ؽx��=�H?n�o?�s?�c?r ��e�$Q^���� S����n����B��*@��B��o��U�C�f��Ј<=櫌�B�/��ܿ?�!<?+D轃G�>r�t� ��H���I��ȅ���a��IP=�}����=��=#�Ƚ�s�wݾm'?��>O�?�g?�p�%y�xK��I��K��v�>J�?�^�>��-?9y��i39��_K�����?�9ґ� u>!�c?�2K?�*n?�����21�݂�V�!��U-�C饾�C>��>��>7�X����<�%���=��r����c���	��9s=^�1?�)�>\!�>��?_�?)y	��3���y�,�0���k<�R�>/h?M��>}�>�MνcD ����>�l?n�>�ݠ>����$E!���{��`ɽ'�>a��>���>�p>n�,��\��X��x|��9���=%�h?r��Q�`���>��Q?��:�iH<�J�>�v��!����6(�t >�n?q��=��;>�ž����{�+Y���4)?շ?����'���q>�.#?�D�>��>
yz?���>�վ�oʻ�Z??�^?7�K?M~<?��>�A�;�x���ܽ����� =���>W�+>�O�;�r�=���>B���%���C=��=����0��ڬϻ]���:{:�o=I�=v"��AT��X��C���%�/���B�����5l�@�����}i��B����R[���PU����E��A�Y���?Y��?O�-�cڠ�=�\��ʅ��4�?i(�^Ժ��uþ(!�Q��
p-��P޾Q8���%ן�������0?F
6��jʿ+����ܾ�M#?@�7?��0?!yg�� =?S�v�����?v ��;�馑��ɿ�@޾��o?�N�>Ɣ��q�;ɇ�>n�>��m>�&T>�轾v�Z�XF*>�T�>�!�>4� ?5꡾��ѿp��/�ڽ�)�? �@_{A?!�(��9�|�Q=U�>��	?Rr@>��.�s>��������>�7�?M��?�(M=q�W�z��%�d?�P <i�E�S��Iz�=��=��=|��ѬI>՚�><�#�=��z�6>lv�>{�'�->���[�ꂫ<�]>T�ͽe%���]�?2J�^Q�v��0u����>�Mf?��>�G3>��?�.�e�Ͽ��?���?`��?b��?}~?Yվy�>����>?�R?��>�9-�(䁿�"_>�3���a:�ݻ�9@�O�&��:?'�j>�G��ҿ����<���<�=����Ϳ�����&�|���-<��.�8�U9�1U��*��(���*T��)���>.>�}=>��>҉|>��r>��V?��w?}�>��>������������t�=�����P�JD���L�������@E�O�{<;�U�A�̾qT�Tc�=Ro.���}�y��ek��r~��%?c�>�,�O>f���6=I	��"{ܾ���<��ݽ	���%ic�0 s�,��?n�J?���d�H��b�������]�j?�Ay�������L���g>?���b>� �>ӊ$<Rɾ��-��XK�,?]�?̱�� ���<�=vm���;Ϻ2?7��>�<=cH�>K�0?�'4����caT>_��=(��>���>�6!>�m��|����	?da<? �`��㌾��#>Ӭ���e8�=��=�w��/����=��j=XO7�mj~���u\�XfH?��>d-<���&�������g->�Pt?yj�>�6�>%@p?e|a?:P��ם�7}���D�T|	�OY?�	�?Vf3>7dݽe����վ��?0{?A��= £�~i־,�����T��>��$?��?_1H���3�h׍����/G?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=��&D�?f��?롭��������r��r�Q-!;�q�=��?�<�ۼ��31�[O���0�l����X�gҎ>VA@��ƽ�a�>�&c��j㿎�Ϳ�������$�H�)?N�>oE�ᙾ�jc��%d��C�*I��E��/��>�@G>Oҽ���~�E��~%��\!��N�>�k�X�>L�s��3W���Ҿ��<��>���>�4>����\ɾzĖ?�����ǿ�R��j��K�j?�;�?)�y?d�?1Q`�@p|�ʓѾ�q�<2�H?�Bs?�0[?��@��9��e����V?���s�u��gA�M�Y�g�S=\'?�# ?i���o>��S>���>K�=\�J��fؿ�뽿��0����?��?.ھά? ��?�M?h������
��m�N�)E>.��>ߙW>�k�<������'����>F�=?^(H�*d!�]�_? �a�G�p���-���ƽ�ۡ>��0��e\�;M��F���Xe����@y����?I^�?d�?յ�� #�T6%?!�>o����8Ǿ8�<���>�(�>;*N>H_���u>����:��h	>���?�~�?Pj?蕏������U>��}?l�>r	�?+�=}��>Ev>zB�������=��P>��:��>�pK?�+�>�Q�k��<!$�jI2�ٖ*�.���>���>9�k?��N?ΐ�>	3��>�"�ܸ(�o���u��=	��=�`���(j�ck��Û=��k>z�3>8�w��V���?-���dؿ#X���p*��4?���>��?Yk���q�����^?'�>�$��c��7��-8�($�?d�?��?�׾��Ƽ|�>!��>¦�>=�ս3�������;>�PA?T}�(ي�$To��ӆ>���?TY@�ӭ?Y�h��	?���P��Va~����7�d��=��7?�0�#�z>���>��=�nv�޻��Y�s����>�B�?�{�?��>!�l?��o�O�B���1=;M�>͜k?�s?�Qo���p�B>��?"������L��f?�
@u@_�^?*�\�g���� ��u��G�=&<>�O>u �cę=�����B��[�<j�_>�/m>B;>�iT>��9>jb0>�eO>eɇ���+�x����˝��	U�����<��n�"�(�}���8z�?���d6�Y�뻙�P����gd�k�,���M�=U�U?�S?ɞr?b��>4��B+>��Y=�"���=���>5�5?��K?��+?�=�㒾�:`�t݀�Y^����R��>SK>é�>�/�>*��>P5��f�L>a>>f	�>�Q>��=xt��KB =BVF>̪>���>@<�>�T>~�=��	��w��4��h�hZ�?�������S��Lq�����ܜ=��?��;<Ց��\dʿg|��˄W?�����6��z!��lq=�%N?�n�?��<dcѾ���=	]j>�������6H>I��������d�+�n>�'?ۄ>�y>�_$���,��<�F����>>x'?���3i�Dxz�2��˾��6>�*�>�j><�T������t����%�=�$?I|�>�(F�_�ʾ��׾�A����Y>�$>u6�=�9�=:�>L�=���m�ȑ��'�P�>g>�?��)>v=P=���>�8��\E�R�>WAj>X�">��>?�?�4;�Ֆ�;��o�'�DU>���>|�{>�.>T3D�o$�=-�>t[>ɲ�<�`�N���N/��%>�vU�v]��&�׽�
�=���=�>G��=t.�1�H���:�~?���!䈿��Re���lD?b+?� �=��F<��"�: ���H��=�?s�@m�?|�	�ϢV�,�?�@�?X��a��=8}�>׫>�ξh�L��?2�Ž.Ǣ���	�()#�XS�?��?��/�aʋ�Dl��6>�^%? �Ӿ�s�>��>P������_�v�o=_�>�H?�����;��y6�y�?�?�������ɿi�v�Q{�>5��?|�?�$m�����΃?�$3�>��?v�V?FZc>ٲ޾մW�q2�>ط<?�7O?q�><���2 ��b?k�?�0�?̯G>s��?)&s?Ed�>��j��~/�Ɓ���m����=�-<�>�u>�{���aF�����ψ���i�����`>�a&=���>���﻾�8�=�]�����C `�!x�>/�n>��G>^��>���>��>�7�>�F=�׋��Q������K?���?���En�J�<H0�=�_��?N54?��_�"�Ͼ�ƨ>�\??�[?ZL�>���0%���Կ�5���\ƚ<F#L>��>�_�>���"=J>2�Ծg�C�ww�>��>>H���)ھp=��(ܓ�;��>B!?��>�y�=|?�&?)�T>�Y�>��J�͖��,:>�X�>7?�>~ ?��?�?���Y6���B����Z�O�d>�"{?5?	{�>���`��;���e3���%~?��m?��Ľ�N?�~�?P�8?��C?So>a���yӾE����}~>32?�罙� ��������%�@?Ζ?�v�>6��;��y�Ѓ���d��Xܾʽ!?��c?�.!?͙̾�aY����
�K<�|��_�=��">^Xн���>f��>kK�<���> 6n>�4>ѱ����<�ޟ>$�i>vp1?�E>ei,��D��0=,?��G�~ۃ���=��r�?xD���>�IL>����^?ll=��{�����x��	U�� �?���?Yk�?f��@�h��$=?�?S	?n"�>�J���}޾6�ྼPw�~x��w�_�>���>N�l���K���ٙ���F��]�Ž/�{��/?�>�U&?\&+?f �>g��>Q�ʾʑ��������S�|��K^�u�8��A�YwϾ5������H(�T׾����-RL>g|�J��>�]�>
�>�ew>ԇ>������>�>x�;�O	�=��>���>:���m""=1�=�@R?r�����'�e��1��B?�0d?>��>ԟj�6��$k���?%)�?o&�?��s>j�h��3+��m?���>���#
?� ;=��"��<����_B�����Ɉ�Z��>}ؽ�H:�G�L��^f�&F
?�8?����A�̾��ؽ ���\o=fM�?��(?��)�"�Q���o��W�S���;7h��g��/�$���p��돿#^���$���(�Pf*=z�*?��?��D��F!���%k��?��hf>��>�!�>/޾>�wI>��	���1��^��L'�亃��Q�>{Y{?��=��Q?``s?G��?з?7�7(�>���ն> /�=��>���=J��?�K?�]G?	�>?�a?��>�����݄��P��>�� ?S?��
?Bi?���j�P�v��:ّ<3��tā�Vs=�u3;����4=q�	���>2�)?����-��O��*l>�K�>n'�>�J?6I�x�s>K�=n�G?�]�=1q#>���eq��xҾ��?��t?�\��=�=ϒN>��=<#�� �$�|!�=6�=���=�D-��Y �0�;6a�=\�=�O>��i=���=��¼��#��t�>)�?~��>�C�>�@��E� �j���f�=�Y>}S>�>]Eپ�}���$��M�g�)]y>�w�?�z�?6�f=��=U��=}���U��t���������<�?OJ#?�WT?D��?��=?j#?*�>�*�SM���^��Q����?"&,?Cq�>	����ʾs먿�Y3�Ե?A[?�a���5')���¾`�Խ�>'>/��}�%��D��_�����&����?7��?i�A�|�6��E辣���CU��Q�C?1�>��>:9�>`�)�b�g��7���;>�u�>;�Q?G��>�cU?��?r�l?[��<�U�@*���O���}����>�_?�U+?���?-��?S�>fV�>��=�z����3����Ӻ������c�=K`>Z�t>M��>jQ�>�><y������!L����<��>^?���>��>��>{Fd>��G?���>矾�k��-����8���C��u?A��?@C+?�=b��fE��r����>솨??�?|�*?A�R�C��=Iм�!��?<u��s�>�n�>v��>��=	�L=�z>�i�>�S�>3"��A��7��L���?�E?:��=��ſٕq�A�p�7ϗ���c<���V1e��۔��[��Z�=�����^�p�����[��������s�@�����{����>oR�=�1�=�m�=w^�<k+ɼR;�<x�J=�@�<9�=тp���l<l�9���ͻ*h��{ �!�Z<�I=���ff��H�?ZA?&%?ͩF?Ec>(/���;�����>Q6�=Ş?L��>I���Ӿ��� A��7)���徳�Ͼ>�G��Š���=c�(�\�=��>�r>&�=�<��,= =P�=�ἅ�>_F�<�=2=���=�{�=�TL>{6w?k���n���4Q�Z�`�:?�6�>R{�=$ƾ@?�>>�1��;����`�0.?!��?cS�?%�?wi�Af�>���Z鎽iq�=%Ŝ�-J2>���=T�2����>��J>����K��nw��(4�??�@5�??����|�Ͽ�[/>~�E>�z>R%K�q-�"�L���e�#o�,�?�&1�3�˾�bS>A��=ܾ��Ǿ�=a�%>�q=����nW���U=~��Β�=Țv=�C�>B�A>�=�˽���=��q=^>5l>����}؁�7��;~�<,�=G�o>Q,>e�>+v2??�S?��?�X�>V:;�-������>��=�(?9��^��>��%>��2?�m?��?�^?�F4=,%�>a�>>gd�_·�X�P�)��͙S��>�?`�?;lr>�9V���Z+��{�D�;;!?��?4?��>����/��"-��9���t`��=�8���u?�vc���[�7�.�	�>O �>���>���>�{3>,�>>��^>��>�P�= ɷ���)=�?��|���R��z&��P��Ҏ�ej�<�=93=��E=ꎚ=�&`�	<��<������=w�>"�H>�7�>���=qg��-�/>�#���$<���F=◣�q�O��re�h,r��,�w�qu[>��>��=|��F��>��T>��Z>r)�?*No?�	>`罞{Ӿ����Q���*��kt��]�<ӆ�XR7�P;k��J�&������>Zf�>�˚>��_>�+�a<���=�pܾ�w7�&J�>Ⱦ��T��n��T�p�9������?�i�:[���E?����N�=U>|?'-I?��?P]�>@b��Vt׾[�+><�k��J�<����m��D���8?�(?���>-��C�6D̾B���ط>eCI�S�O�Õ�-�0����η�X��>����о#3��g������Y�B��Rr����>Q�O?��?�.b�V��jRO����C!��,q?rzg?w%�>�J?$A?���y�k�����=3�n?���?�;�?!>�z*=��X�-��>B?U��?�v�?e�r?�l�@��>A�O���\>�����*5�=:�=w�>���>�7�>$�>\*��A��Feᾭ�������O=�ĭ=��>}j�>��T>|��=:G�=<��='�P>Z�>�X�>�\	>Z �>>х>q�Ծ�/�A	;?���=�i�>U�V?e�>�ӽv��=��L���U��1����̾s����m�=gA7>DI�����"����>Gi����?=�j>��le�>BO޾���;S��>'�=��꾔�>G��>:��>!�.>e>��>�L�>L�=��Ҿ�pT>����.��>�z�z�6�����>EǾ���#���= �����ϾgWȾ(�T���g�$yo��T�?8Tp�*���gB�aZ��#?�?��C?���dJ�=m$>��?߆>$���U���̓���ྨ؅?H��? 5c> �>��W?�?��1��"3�uZ���u��A�he���`�፿ۙ����
�$´�_?�x?+}A?t^�<�8z>顀?�%�\᏾d5�>%/��*;�K5<=&3�>A,��T�`�B�Ӿ��þzC�>VF>i�o?&"�?*Z?�?V����tX>�fA?�QC?�Ag?��%?2�6?�Fi�6�?�@/>h�?���>|=?�K:?��?5pp>��W>)�;�q<�����s�J���L��M�kӭ;�҇<4��<.Iv�n���PBA=��=�K:����<2.�NQ<&f�=��=���=�C@>���?��>�8�>n�?���=Bs�V����?6f(��&����M��}*�F�����>��?PV�?oe�?��>n=(�U����E >)_=ƪ>��?�w>n���DS��`�]ǽ��a>c	>M�>�\���>���+��ٽ
'3>��>�B�>��=m��>�ǻ�f!��� �>f葾x�������L+�t�o��멽�4?��?�h"?�ނ>�C��9���#��11?�Ko?�Ka?bÅ?�5<�P�P�b���:���/��Y>}�;�3�������b�j���<j��=�D+�����#�a>o��޾��n�4�J�%���\=����5S=�z��վ�K�c��=0$>�7��X;!��G��2�����J?��p=������X��Ѻ��`>J0�>��>:@���l���?�H��|��=O�>V�;>�K��a��٬G�lk�l�>D�G?��u?(#�?������t�|1F��C �91���1
��$?FN�>�?�dR>���=���x��&\�e�R�p��>���>�X�l/�����bB���(�o՚>�C�>�
~>�X*?��K?F?e3e?l�"?P�?`[�>�耽�x�h?á�?Cq=*_I�`���
w/��&Q�B��>�h)?��@�	=�>xl!?���>K#?�J?�l?�a�=�����3�R��>��d>�#Z��>��Jq>�YY?���>��c?�dx?�%�=�_J����9�-��3D>��%>ʲ-?�B
?[�?��>��>N̈���=��> �\?��?�o?�>z�?m{>t(�>�;�=.��>��>�o?	�E? �`?�@C?���>y��;xP��
½�𞽰�4�ݪ=�rO�:�[=���<a��z�,	ͼѱn��h�;P�X=32�<h��Z>�	c��,'�>�cu>�ꕾt�/>ټþ����>>�_��w����F����9� ��=�?}>��?=n�>A3"���=�M�>���>M��x�'?�)?U?Aa�;m�b���ܾ�M�N�>��B?�|�=�1k�q����u��o=�Wm?�
^?��U�Ҏ���b?��]?�
��^4=�}ľ�a�����#P?�\
?W�G�2�>>�~?¡q?���>b�e�an�2��<,b��j�^�=܊�>�E�[�d�9�>`�7?+��>��a>�D�=EF۾�+w�C��m�?w��?�֯?��?��*>��n��j����6���8\?q��>A���!? F<�оୀ�A����Kᾛ ��M������E���� ���{��h޽��=�m??�q?�Pr?��\?8L��Pa�{�\�N���U�/&�Q��(�B��uB�:=D��|s��\������Q�<Sօ�>�c��?�"?;��] ?�98���?��	�yE%��∾Έ�)����A��gKO>�$>0���B8y������&?��?�#?F�a?am����Y��W�g���S"�:�>���>�Ӵ>�7?��+�v�Ծ�Q�����^�̽�[����u>I�c?��J?�<n?���Q�0�ʂ�J!�y�#����k�G>7>�W�>lwY�y���%��=��p��`�ą���	��fl=�!1?�N�>9��>���?�4?��Fy��Z�~�ZS0�MP%<�M�>�Zh?P�>��>hLȽX` �?��>��j?��>`��>����.&$�|{��ڤ����>�3�>��>u�~>�A8�`Za�*����@��;�9��R>�7h?C���v�^��d�>7�N?I�A<�d<ۮ�>�P|�G��@�꾚���>��?Qg�=@�C>��ž!�
���r�쥆���&?Mo?󪖾�-#�w:�>��'?"/�>�+�>� �?tUl>�̾�m���w�>�kZ? 
G?R)>?���>��<�a߽.�򽠹���@=a9t>D35>��=�u=��-���O�#��p;=gi.=�]��|��t�o= �-��]<1�c:/��=.ܿ��R�i�}��E׾EѾɳ�_�ݾX�2��������Z�׾��ƾ�YѾS�a�o����Ƃ�(��������}��`�?T1�?ϥ���s=���j����I>��"?i��љh���	�w=S
k��i	��z�b�A���0�������,?pA���̿E��������??O?�?�_���3��@����=֓ٽ�>��@r��	��'þ��T?�ѐ>0G����a;GZ�>���>dx6=�S$>����$��AS�`ۓ>�PD?u�s>R����׿��˿��&�4��?!�?�oA?�z(�t��"9R=t�>C�	?��A><�/�
(������?�>�0�?+׊?�M=ȬW�]~�[�d?3@<cF�kͻ)��=[�=h�=?w���K>�G�>���^B�y�ڽ�2>�^�>a��+���4_��x�<q]>,1۽����ٵ~?#G:��DJ�hG*���i���>�??rfv>��<>�c?p�*޿��E���w?��?s8�?� ?37 ���Z=In�x�<?|�E?�D�>��=�w��� �;>�P�==m."�� k�t,u�%?��(>j����'�E*��=a�;k3>������ۿ���Y"�~ż�
=]��0�U��֋�sW���h��g���O2� �=��6>WW>��>;�>R2e>b�W?܂�?��>^�+>�%w�Ё��񣿾F�'�~݂�,�8�gA��
�L>Ӿ`�о�5���S$�T�Q�IH��ζ���<���W=�%@��y���(��b���Zu���:?�֍=Q�о@TU��㽼x	Ӿ眶� �;=$l���� �O�Fo���?V?p���5_�����W��lO�x~?�b\���������e>F�|=�-�<w��>���<����KE���1��Z?��"?7���mx�+X>�Fؽ�5�t�?�F?�~�;�f�>�&?Ç���Ȋ�[�>c�M>�b~>Hp�>�V���ƾ�R���Q!?�>J?��:�;��b�}e꾰� ��ӎ>q��>�7�=�!��1�=	;�=�@c���<��Y<a����xM?Mz�>C?(�U��t[`��ݽr4�<WNx?���>D�>��h?E�R?9 ����Z�S�(,�O0�Bj]?�p?�9>�
��0���ء���?�0k?���>�Lh��nپ����%	��3	?��?�h#?��S�UxZ�󞅿XO��B?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�*��a�?���?�੾�~<�u�K�n�F���vH<��=�e&��=#�_�� 6�BSľ:`	��Ŝ��������>�@	�ٽ��>3F�a[�ϿR=��k�վx�d���?ƈ�>����堡��nj�rs��WG�xG��H��V��>-�\>>�����e�]� �Z�
�
��C�>�&Y=�	>��:���ݽ�E�}S�=;Ǫ>�Z�>� 2>�6S=�׳��A�?����5��ň���+ؾ��g?,�?_;{?��?���Ǿ����:�$=l�w?��`?���?埦=���pZ彐[?����
�h���;��R9���^=��?�G?�7���缑ǆ=m	?�,�<�\'�bwĿ̧��@�����?�6�?�5���?���?e�??#������ʞվ��1��o����U?+��>,���z��c*c���G�i�>_N*?.��z��\�_?'�a�L�p���-�i�ƽ�ۡ>��0��e\��M�����Xe����@y����?L^�?i�?ϵ�� #�`6%?�>g����8Ǿ��<���>�(�>*N>�H_���u>����:��h	>���?�~�?Oj?���������U>�}?��>}�?���=��>��=�%��Nj@�t#>+��=��;��?2�M?�H�>���=�7���.��$F���Q��y�C���>g�a?��L?�Kc>]��۰8�\!�ޖ̽��/��ؼ��?��3-���95>I�=>�>k$D�F�Ҿ��?�o��ؿ�i��*o'��44?b��>O�?\���t�n��<_?�y�>�7��+��&��PD�!��?pG�?��?8�׾XN̼9>��>�I�>u�Խ@���������7>#�B?��dD��1�o���>s��?Ķ@�ծ?�i��	?���P��Ua~����7�_��=��7?�0��z>���>��=�nv�޻��W�s����>�B�?�{�?��>"�l?��o�P�B�{�1=8M�>Μk?�s?�Po���f�B>��?!������L��f?�
@u@`�^?*$��KĿH��� 쾻k�=X5G>�\6>p�g�>>�Fj=��9���3���=�%/>��>G:>��S>�H>��5>C5���A*�u˝�uG����[�[�����o����^������ݾ�e��^o��]�=��n<�]����ɽ��ý�e�=���=��S?�
Y?��y?� ?��^���
>�M�Ǚ�<n�(�8A�=ej>J"2?��M?�<)?���=Xچ� p]�8��F������f�>I*R>�P�>Y��>�$�>�4�<|CM>Y*>���>��>���<񾫼>�<�g;>��>;6�>`Y�>y�l>��>�ƹ�P<��Q	��[�8��)��뗬?$�ھ
6�����,��}��k�=�?��<Ә���dǿXg��]_G??�˾������'m>��E?��d?�o=�;�����z�>�C��Tc9�	�>����Ǌ]��L��
>���>3�u>�>a�/��4�m�G��ǜ��|>�C,?OH��Gr^��+o��zH���㾵Gq>�}�>�<As�t鑿=�z����e.�=]k;? ��>�,���ž`Ǎ�Z��S�Z>f�u>{ �=U6>C89>}WJ���y�3,W��A�=�@�=�a3>�`?->,Zn=�`�>�P��OI����>��F>�;>��=?$?�w����v��Ƅ��p8��b`>���>��>!�>��K�{R�=n��>�R>>
������DgD�&J>v[��E�]�펽;K=�ԫ�e��=�{=���L�8���<�~?���(䈿��e���lD?S+?a �=�F<��"�E ���H��G�?r�@m�?��	��V�?�?�@�?��K��=}�>	׫>�ξ�L��?��Ž5Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�>�s���ؑ��yz�Hn��AT��U�>n^?����>V�m�/K9?T��>���u��]�ȿ�x�L��>�}�?��?ѩn�@؋�ߡ/��'O>n�?��?k^>�j���w���P�Ӫ?Fx�?��?0�6�j��=��	?�c�?�fx?�H>���?�Nn?���>zPE���1�)ӳ��Y��&T=��<�z�> >��ľ6�J��
��gg��/j��?���g>��%=!ȶ>�nݽtm��U��=H����Ѥ�Ǿ^��v�>lq>#U>�ř>Z�>0��>c�>c<�<�S��I�n������K?y��?�����m�#�<c�=E�^�X�?�?4?��h���Ͼ���>��[?��?[
[?�q�>ћ�Y������������<��L>%"�>�=�>�n���oH>�#վ�SC�6��>�	�>	ډ��ھ�9f����>�P!?c��>�i�=�?>� ?2B>��>��3�X����C����>C�>g�?̡?ܝ?#&̾��@�b����榿��]��T�>��y?�X?(�u>J��'	���>8���e��];y4w?��]?�둽Փ?���?�>C?��B?"]>�C� lѾ�6��Cs�>R=,?		ֽ'�L�v>�����d�I?j��>v�>�=����漲��-��rA?t�Q?�*?�8׾ie��e��f��k�{Y==���E��>� i��c����c=�>��>J�&��`�_�/�23>Y�>X �=�nľ���)=,?��G�tۃ���=t�r�CxD�T�>�IL> ����^?8l=���{�����x���U�� �?���?Uk�?���<�h��$=?�?Y	?s"�>K��~޾H���Pw��}x�uw�J�>���>��l���F���֙���F���Ž��#�U�>���>�?Z?�n�>@\�>���O�|ľm���j�2"�0�F����J��x�}�v}[�]���>�ʾ������]>i�~��a�>67?�P>�h>�ȸ>��<���>cP�>�E�=xo�>��>vOW>=h;=Q�[��R?��Q�(���꾶�XB?��c?_��>�+x��܄�W!��?A��?�!�?��u>��g�.D+�y?��>�}�;S?�5=��_���<�z���t�J �����j�>��ɽ��;�PL�Lhb��x
?T?��t�WϾ�:޽4�����n=mK�?��(?��)��Q��o��W�$S�����@h��g��J�$���p�ꏿ�^��%��D�(��U*=��*?<�?:������%��/&k�W?��yf>���>{(�>(ܾ>�sI>��	�E�1���]��L'�����G�>�Y{?�%7>?�D?�w?:�?�H#?uiW=���=���Ĝ>�p�=��)?��s>J�A? ,\?ax/?J�;?�W?�/�>7�Ͼc8
�c�����>�t.?/�?�?/�>%E��(�Xpk��1>��D�)Ȋ<�fx��������fm����{=��>�)?�%��d�@����<s�<�>�L?
z�>���� ?fҾ^��>| k?`Ҿ`����GH����ъ�=r*�?$����F�U�=���=���=�}b<��0=:3���T'>F�����;"X�����o�=�f3>SL:>�^�<�^9<q2K�Li�>��?g��>�I�>���o� �&���.�=6Y>T1S>�_>�پ	}��]$���g��2y>zm�?�u�?��f=+�=o��=j����T������ӽ����<��?�<#?�AT?���?��=?bZ#?�>b(��K���\��J���L�?��*?X��>_��}ؾM��� 3���?�
?�a��3�G�(������J���	>�>7�����㯿��8��=�@�}�-�R��?�?�(����=����L�����!kG?�&�>��>��>q�1���`�x%���:>�*�>JN?�G�>H�X?0�?]�|?�>�g�c���ۮ���Z�<���>婁?�5?rq?U�p?�O�>��>K�!>3�����G���o����񌚾���=���>E�n>�q�>	��>U+���~�:�6m������I<���>���>o�>��?}�>ܡ!�F?���>Rݺ�*f��ϟ�s���U�@��jt?��?�'?lC2=__� E��\�����>鷨?��?j�/?��V��E�=�����B�����+T�>�w�>�B�>ߠ�=2�=G�>^��>f �>}<�+[��7��2���?�HC?_#�=,ƿŮq���p��З�d<����	�d�ٔ��[����=�������wǩ���[�絠�򊓾�����I�{�'��>�c�=���=��=~�<��ɼ��<b�J=�ɍ<˧=��o�(�m<d�8��Yλ���������\<��I=��;˾�}}?RI?9s+?&�C?��y>�>d�3�z��>2̓�
?��U>�PS�SR��-�:�f�����Ċؾ�}׾�d����y*>�=J�1y>��2>�f�=�j�<���=�Xs=��=�aL��=L��=��=�ǫ=(��=?�>Ҡ>E5w?ꖁ������2Q����ٻ:?y@�>�}�=Qmƾ�@?x�>>x+�������N��-?���?UO�?c�?�{i�4k�>^�������#�=&��N2>���=��2����>K>Rv�L��,M��h/�?D�@O�??�ڋ�ϤϿHB/>��?>��>�&S�01���A�I5����m��Y&?u�<������>�J�=���UJ޾)�<`{�=���;�	�_�G���=nd��U=;i=�K�>��9>���=�&����=�dy=� >QFK>ҫ���G��q̼VT�<�=S��>�z->'�>#?u�Y?E��?�&�>�ž����J����)�>�����D?��=�΀>�^�>�J2?��^?���?�H=? -4�-%�>�Y�>�)u�]����p���6����=%S�?�	�?�K>����N��=��C���*�A)���� ?v�;?�)L?<�>/����YK��
F�|�'�{��=�jT=	��"=�J��F�½��%��ī=��>�K�>��>�ʪ>˦�>�`k>���>C�R>܅>�v�=Ex��]�\kҼ��=�a��屮�=x<�ힻڰ^��L=;��=�E�=f8=4�=~G=u��=���>�>���>��=�ɳ�/>����"�L�[
�=W��%8B�(d�YQ~�2�.�666���B>��W>�Մ��*��+�?jsY>�U?>��?�/u?��>Z1���վ�0��l�d��	S�;϶=�%>�=��_;�AV`���M�*Ҿ1Y�>�&�>�yz>�;>�G �kI����:�M���Z=�'��>��y���e=	�:�ST~� 餿!㥿�k�qe�<v�H?�Ԅ���>%t?�L?���?z��>�� �Z;ܾ*l&>�#���	>E����m�VP�n�#?�M?�?�>�о�<@�}C̾����Zַ>�BI�N�O���8�0�ώ�ҷ�o��>�諭��о�%3��i��J����B�[Yr�E��>U�O?��?P=b��U���QO�T�����r?�xg?��>!K?fA?����v�n���= �n?��?<�?u>o%�<��<���>��>��?j?uNC?lW��2?1}W��P>)��-}���>���>���>2�	?�P�>�(�>ⲻ���1��r־{�/�f฾�]�=�n�>8+|>K��>$D-�V�>P<� >��>3�?Z��>�{�>=]=�d>M����C�+?��=S�>0�6?>ؘ> +-=�c&<����t8ļEJi���n�vm���K��=e�4=�a�Y	�����>�¿va�?��B>�i�?&<վM�+�v�>Y)>E��ɿ>_�>�y>��v>�<�>��=�5a>T"�=
M��YNT>���"��Ji�b%���'J���?H��`h��g(��'�<}LZ�Bg��䚾 m��$��0��F4<���?���q�����f��D���'(?Uc?ȓ??����[p=�v]=��+?��>~fؾ؇������?ؾ�Ӈ?�y @7c>;�>��W?�?�}1��3��tZ��u��#A�Ee���`��፿����
�����c�_?D�x?yuA?��<'2z>���?��%�ҏ��/�>�/��%;��7<=P*�>�%����`���Ӿ��þ:�PKF>Q�o?�#�?�X?IV��7`�S�*>
:?�2?��r?��1?G�:?���DG#?�+->�4?��	?f	4?�/?��	?�6>/8�=�����=�����߈���ӽ��ɽ��弩GA=��u=�"�;�t�<�f�<���<�a��6�@ ;@�Z���<�G=�Q�= �=��s>�g?��>�Q�>�2x?�0n�^�a��ž�?&~��xy2���= ��Gd����>F�t?�6�?�W�?
��<�1J�H$��9�=R��>���>}�>��Q��Ӕ��a=Ⱥ"=�3�<4Iؼ��:>U�ӽE'��Q�!�`�8U��_��>
��>�u�>�@'>5��>�����H�.d>�
��1��:�ݾ��P�jق�(Ȫ�5W�>�W?~&?�Dd>�� `��9M����!?�q?�rb?���?[56>�-���a��F���O=��N>:V>� !�A���Ǉ����H�։Z��@>;3������~#b>��S&߾�cn���I��;�ņS=���GD=,q���վ�+�����=5>��� � �l ��8W����I?�m=#���<P������>�[�>���>�>��z��A@��ǭ��z�=!$�>��:>Q8��9��G����$�>;	G?��{?ř�?����l���C;?�����ƃ��=S0?rA�>4?
�=��=S=H���ؾ�L�wX�1G�>?sQ$�!�2�䶜�������'�
��>Q��>�1>(�'?��F?��?�j�?ZY?�~+?���>)A�^��$?���?��= rw���Z���=�?�B��w�>��$?bx.�A��>��?L�?e�,?�tQ?k?��>�	��#LE�>q�>���>�Y��|��e�k>��D?�ʹ>VnZ?��~?�9:> a5�3��"8��>�1<>/?�?=�?�6�>���>�p��[�=�_�>�c?%�?��o?��=�?}�1>���>w�=,w�>$U�>y�?�EO?ٻs?��J?`x�>tی<�l���̶�a�t��E���;V�<<EDz=��qu���w�<'q�;Qո��9y�����bF����*��;�Y�>��s>/��q�0>dž�����DD>��\���W����=�s��=Z�~>if?���>��$��܋=8Z�>^��> u�y�(?�V?l?�ޭ��b��BܾиK� ��>�t@?���=��j��|���?u�
�t=S]l?�d\?<Q�E���!(X?�,?9���<��4��ZD�J����U?���>պ۾
�N>�Mm?2.?*�>�<����e��<��,�=��w���F?>]��=��'�[45���>�R?3B2?���=eH>����#a�P��?�$�?�|�?"X�?��3>Ѿt�E�Կ(����ݑ���]?�R�>sϦ�A"?V��F�ϾgF��o���W��������(T������$�����{�ؽ2"�=��?Ֆr?�6q?H`?Ξ ���c��]����Q'V�bB��'�j�E�$�D�\�C���m�g���<��*����J=/t��H��t�?z�1?��Up\>��?���4��'N�@�q�([��{���>��>�
t&>+ZT=(��%=��6���2?\��>`P ?�q?����J)K������8������>��?���>�d?�N��L3=���=(n��ܡ�a����pk>�la?Z�M?�Xk?$��0������!�e�ZU��\�8>V% >���>��X���"�H�#�ѡ:���n�������_���j=@�,?rAu>-[�>���?Z?yF	����(>���2�D� <�¹>
�l?Y��>{��>#���k����>/�i?�2�>�_�>���0' �S䀿��k��6�>���>LQ�>ZL�> D�{]��"���Ҏ���4���>��d?"����}�[Qv><I?�p�<5�t<E�>鵂����h�ng!���	>=��>�)�=m�>�Dƾ����;s�����e�)?��
?`����+�o�>�;"?�*�>J��>r�?�N�>}�Ǿ�'0���?�y]?�2H?��??���>�=����Ƚ�'���;=12�>KU>��a=��=�����[��?�~�R=�r�=�mԼ������v<�ָ�la<*��<f�/>�_ԿBwZ�&��n�]��4#��/��)��*6=}���%l7�a�T�g܇��8e��(���ѽ
n��T���|�l�����?�1@�W��;���z���"�� ����?lH���sY�$?��|�&ᾆ�ݾD�R�����z�]�|��s�r�'?T���ǿG���5�,�*?��?��j?Ψ�R��?o=�pM�=k�<�Q���h"��`Xο-���ֵe?���>���W���(�>^��>�Fn>f)f>},��=��Ga=� ?/�"?%� ?�`p�p�ÿ�M����<e��?��@�rA?��(���쾠�T=��>��	?+@>ƽ0�,@����
��>�"�?�܊?+qL=��W��0�6e?�C�;q�F�Ԟֻ6�=�1�=.�=����'K>Ȧ�>�����@�d5ܽ�m4>�Q�>�m!�����]���<q]>wֽ�����!�?�@�dM��kH��Ht��f�>߳W?Eo�>	�">>?f%��ſ�&����?:��?�}�?�?���S=����yA3?	J?�>�$b�l����
>"/��B�;��3:��b��r��>��S>t-Q��	��	��iĽ��;�]��pǿ��#�� �q��<��]��\��������CN��2���sk�<aڽ��l=�b�=�'R>�Y�><<X>z<X>l Y?��k?�
�>��>������*:˾�uֺ����vz����<��C>��U�63�:�	�9I�����R˾u=���=]*R�N���0$�if�D�E��H/?� >�vӾ��N�k2:rо�����橽��̾ap4���o��|�?��H?�H��wiF�3Y	�8�S���_Q?��Ģ��,��:��=����io �8�>�sK=p�����<��+K�ƅ?��?Yp����>ط>白=�4�`�6?YԷ>{�<�T?��q?�誾�F��7��>=��M³<i�<?9�P>:�xmw�X�?��X?�>+�J�Ͼ�3��~�x���Ҿp6_>�Qf>��h=`��rf��j�=������=�9<�Bֽ��E?5�>d������a���_>��GA�kht?�z?i��=�yY?L4K?��HI��F���%��-<�7�P?-�f?��>U�0��8쾭\����1?�0[?�> n}�Yo澅0����Mt�>:]?�� ?�Ký��j�����?�	�\�+?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������Z�=~'��U��?:�?z���><�����l�����"��<���=9����S�Ov7�;7ƾ�g
�.����Ѽ���>\@@)��g	�>��;���Z*Ͽܹ����оA�m���?�ϫ>g��ލ��Ek���s���F��I�붍�ݿ>�E>�`�������P��������?���7��={xJ�ϟ��Қ���q=��8>���>�IM>W�2=8����;�?���^ſ G������@�g?΃�?}�s?�(?Ȥ��	|���ľ�
>��p?5=m?�tn?zT'�M獾<J��d?�^ؾY�v��g,��wC���>��?�Y>�<��`k>R�T>�Y>�'�=̛C���̿�����!�2�?C��?Eq뾪5?^
�?�w?
\�j7��⠋��$�0��=�?��>�3Ӿz�� ������?��(?��"���^�_?(�a�L�p���-�x�ƽ�ۡ>��0��e\��M�����Xe����@y����?M^�?i�?ҵ�� #�_6%?�>c����8Ǿ��<���>�(�>
*N>�H_���u>����:��h	>���?�~�?Oj?���������U>�}?���>D��?�=��>��=���@�Ҽ�)>���=GK!�M#?J�O?�>�=Y�3��</���D���N���\�C���>Tka?�K?�va>�����P�����G̽�+�;1��<��8-��۽�+>T�:>.�>�B���ҾL�?�o��ؿ�h��Gx'�)54?ֹ�>��?w��:�t��3�=8_?�y�>�7��,���%���N�+��?G�?�?ý׾��̼�>P�>�M�>/�ԽN��-|����7>�B?���C����o��>���?ǵ@�Ү?�i��	?���P��Ua~����7�e��=��7?�0��z>���>��=�nv�ݻ��W�s����>�B�?�{�?��>!�l?��o�Q�B���1=7M�>Μk?�s?�Ro���e�B>��?$������L��f?�
@~u@]�^?*hֿ���K��ė�����=���==�2>�ڽ�d�=1�7=P�8��O�����=O�>R�d>�q>�(O>na;>s�)>O����!��q��Q���R�C�-��~�d�Z�J���`v�{��4�������<���&ý ����	Q��+&��8`�J?�=4�N?�ba?��p?]^?�D_��M�=��
�y�=)���	A=�&>Y)5?N]??��?�v>{�k���^��Ղ� �ɾ�%��f�>9�=S��>y�>^>�������>@�/>�h�>�x:>�^�<*�@��
� W�=4�>���>�j�>�>j�0>�Y��0��b%j��%����lP�?�L��h�R��ɕ����� ˾�6<�=!?��=�R���rѿ:ת��?G?�.f��^
��Q��>>�#?j�F?�>׼پ-�.�U�8>'�!�E�r�ج�;ܯ���_��Q�>��>E�.?hh�>e9>S_3�aq���M�3�E���>�SJ?�Sľo���h���t:�l�����>���>�V�:(��䗿L�N��	���>�_>?m��>�<u������q���/����>�G=�y�=��'=��v>k��Ŷ�=G_G������4p>�G>g��>y><>2�>=?|�����\o>�*>���= WI?��2?4�<��A�|�F�A�p�xV�>�>���>�Ҫ=���"��=y�>~8>�Jƽݍ��֛T��d)��u%>%����O��-���=�Y����=��=�,�<
�K��fx<�~?���(䈿��e���lD?S+?` �=�F<��"�E ���H��G�?r�@m�?��	��V�?�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿg��>��l�O���$zV�����7">�ޠ>��W?��b� xD��<��cW�>��P>�w�y`��tHɿ{����/�=W��?��?1���@���}A'�|��>�2�?%AV?+>��3R����fp���Y�>+?u>�>��4�l���`?+)c?2�E?P�K>�+�?Ugm?��>���y�-�
{������WX)=O�=΋�>��<>D�ʾ�J�n䊿����Gd�V�
��gb>�Z�<h�>2�Ͻ�cƾ݅=q?���D��ļ���>?�f>Ӈ4>�>D0 ?�D�>؝�>��<�a�b���5W��L?,��? ���Pn����<�E�=��]�.?�J4?�uW�q�Ͼ�e�>�\?�ʀ?�-[?ܔ>í��8���ܿ�G����<��K>���>"��>`����K>�>վkD�~Ί>���>I:����پ�Ձ��(���m�>
>!?���>���=��?q�?$�N>�rk>�!�&�|�4�s����>���>a�0?�@z?�I?)�.8��և��I���A�v�>�_?$�2?R��=�Ӓ��}��r���	K7>�J�=ta?&I?�N���S�>w�t?�6�>':?�b>{�D�%���hϽ<N>�0?�H�;H�{&�r3˼�=?D�9?k��>���<�W�u�6���	�߳���'?�:'?�
?2�込E\�bΓ�#���1	�J���0B�< Ͻ��>�-�>��{���{=���>s/:<4�㾫����=HM>֑?)8�=�P���C��*=,?F�G�mۃ��=y�r�;xD�u�>�IL>����^?0l=���{�����x���U�� �?���?Vk�?[��=�h��$=?�?H	?i"�>�J��~޾0�ྯPw�)~x��w�p�>���>�l���E���ϙ���F��F�Ž`��z�><�>2f
?܉?�QL>���>j��^2�rƱ�BJ���e�~"־Y�'���+� ��5����B�����*�e��Ak�>��޽e�>{�?�+><2!>3?�[[=5�g>t�">{eM>A�>�xz=t�>�q>Gg'��	���W?�L����#�%F���z��O?p�W?>`?��;R���F �*�?[�y?
�?���>��Q���!��>���>h�\�#�>oI-<\P�L.M=CQ��5��mm����r&�>�a����]��� �uU�
�&?#b;?�[�$���XB�F ���b=$��?W#?+�)���P�4:j�;�R��T������`k�~š�<�|�p��4���v���+���;&��x�=t�(?֞�?m;��Ta��b�e�z0?�]g>���>�H�>���>6f>�����3�kW��)���~����>hx?��2>��\?]bN?�6{? �]?�m&<��=���
�*?׋[=GV�>�#�>+?�O?؝A?�e?�w?v�>�Ѭ��\��*˾b�?d!?(?�(?��>~��e�=d������둾��>��=}~Z=U��E����=^�+>QA!?�g��w&V�xs�K��=��\?��Q?}E8>�d���3�<���ŏ�=E��>��>n�*��;�c��=}<���l?�+V���n<�^�>�mn<���=�x�<��M��=mA=`)O>d�[>�Z2>G�����R�N>����l<B/j>�G=B��>b4?�΍>N��>�Lv�H`�-��
�=
�S>~�i>�->,Dþ����S���Td�w�e>C�?v2�?z�d=��=���=3[��5¾���b�����<t ?�!?�P?�ۑ?�;?�?~�=�B��⑿(��r䜾�k?�?<��>���fKվR+���n���?��?U�i�����6dV����9��=l��=iM�:uv�Xw����9�ڡ>q$�[�!�[x�?��?E��<~�G�o�ɾ���ʟľTX>?r�>���>���>i�K�k�>��� >�?�>5?	��>�HU?O�?q�?�p>�^Q�����b����,<�Us>��[?'1U?}1�?�0�?�E�>��>k����G��t�,�N͏�B�h�Jiþ ��ҏ>1u>��>M��>~�>>J��L���탾��<Ј>�U�>��>F}�>�1�>��r=��E?ʲ�>²���	��'������V91���r?^А?9�*?�-=��B�D��E�����> �?�$�?�,?�Y��+�=2��h���l����>`A�>) �>�\�=�P8=d�>�)�>�.�>�����6�I��?�bC?�t�=��ſiqq���p������a<�-��q�c� ���5[�-�=b���-D�Mǩ��r[�@������µ��	��R�z��q�>�(�=���=��=�^�<%Dм��<�L=��<0=� s��Ko<j�9�p�ܻ�:����R��'\<�$J=�� ��̾"�{?�lK?H�*?e]D??�v>)�
>OBd�D�>�zS���?4�O>Z;9��A��3D��e��k����ؾ*#پ;Xj�Oȡ� �>�$���>��%>{��=?e<���=��=X�=զ�4K*=OL�=�=��=�T�=��>}6>�6w?�������5Q�/S�H�:?�8�>���=�ƾ�@?��>>B2��_����`�.?��?cT�?��?�ui�'d�>a���䎽6q�=f���m>2>��=��2�y��>�J>$��`K���x���3�?��@џ??vዿ�Ͽ]/>dZ8>o�>sQ�o�0�
[��"b�2�\�F�!?�l9�[)ξ종>q�=��ྚVȾ�"=�G->�~N=�Q�Q[Y�c��= 憽��1=V�T=R��>�C>_�=����3�=ec8=� �=L�T>	|	�eN�ފ<�xp=B��=��a>Fj'>G�>�L(?k�R?N�?�š>�V�󊊾���c~�>�j�>L�?��`��u�>��>�K?�!s?撃?p�?N����.�>Dt>Ѵf���o���b�oi9��:>*0�?��h?��T>v�ƽ�'=ÃN��5��{$���?h�K?�1?�
?�!��z�5<Ⱦr[7���z��<l騼�վ����YN�/��=�޻��E>6!>���>�	�>q0�>_�b>�>���>:*>r#4�E�ռ�#���ޜ<��=E@O>��A>i):>�u�=��=�
��"	����!ͤ��}��C�=���= ��>{[5>(�>��=`.���;->z>���]J�{ɼ=\奄��B���X��ny�X�&������.>�:S>����M��{V?�mi>c�J>W��?N�w?��#>w۽g˾�J��_|p��b�A��=VD�=S=p�M53���]���F���ɾ���>�>H>�
>��=P�>��B���=����f�>����>�ڦ��g~�Q��;�g�Y��Q����r��0����^?�։�?�>��?ߘ%?tee?\�>�Q =E�K��4>s���"�W���־��4���=C�?F�1?�?������=�s�ʾi����Z�>�K���O�7&���E/�;�E%���%�>�d��[о��0�/\��}���B�:w��R�>-�P?\S�?�9f�񐁿��N��+�66�$�?&�f?(ؠ>�?�?���X�S#��9I�=�	l?u��?f��?�	>�ɲ=�䥽���>�(?���?m�?Wn?ۭI�QW�>�c�:�">E����5�=��>�W�='��=ǅ?��	? ?ܹ��vJ
���f	���'d�m��<�`�=0/�>~n�>[
Y>F��=�|R=�P�=$�[>#�>@ǉ>��]>&]�>n?�>Wo���|����7?^�=t�>�?��M>��߼"\4;l����C�OA���~罯~��"佚�=���<9Y�=͙�b6�>�����@�?�2>�Y� ��>�����J����1>�4=p�f�z��>�p>��`>��>��]>r��=cϣ>�8>�%þps�>�"��|	�^��x��T��}&�>�F��|���A����X�N�׾`#(�Sپc�q�]"��b�r����="�?X�a��(o��U���1�8?��>b�6?��6���'=d��>~r?�i_>U�ݾC������m�)���t?�b@� b>]�>��W?\?zn0�un3�?\Z��u�b�@��e�!�`�aԍ��Y���x
�)�����_?�x?EPA?��<k�y>HA�?�%�����>f+/��{:��6<=#��>��]�b���Ӿ��þ��C
I>�n?;ڃ?L�?��U��%m�n'>%�:?��1?&Ht?��1?֜;?!����$?�>3>�,?+f?�K5?��.?w�
?[2>���=�窻}(=�(��H����ѽ٠ʽ,�#�3=�;{=R'��S
<u-=C�<׊�ڼ¢;�Q��͘�<sc:=��=�/�=FU>'�c?��>���>�A�?��{�#�R��ؾ�i?e���
;�#;C=OH�i���Y��>��f?擲?��|?�3>�q�����Y��=��T=�>>U(e>vN�=��!�P'���<�+>�����'���G�ھ�PC��0>3��>���>ѧ�>��a=��'>	-Ѿ&A��܆>Ե���v����P
&��1����fP�>�E?V�?��I=%���c�J���$�#?Wrd?!]X?E��?�s��_%�A�2�i[.�5{����>�/r>���1d�����J�E�T���7�?Qi̼="��,�a>�����zXz�ST�3�ƾ�ؔ={x�h#�=h�����[d��o<	>��>	�þ�V�8���m[��Y�M?�m>�}��e�#�%���{�=�<w>�I�>��k��4:���6�:���,=���>��4>y-,����;�?��W��-�>�CP?ub?)e�?�X<��/���M�OKԾ��Y��M=�e�>$m>r�?��>��@=�δ�r�{o�`�J��>X�>Ź/���R�%>۾�{߾�ܾB�>&��>�U�=��?��P?J�#?k�i?ǻZ?o�?��<>�}G�U����&?a%�?�`�=�ڽ �J���C���.�ee?@$1?�Z����Q>o=?�O!?��:?��^?�/?}�E=��4���R���>7��>��d�׺���_>�@?���>��V?`�?��=���k ����ѽ�t�>ْl>H6?��.?J2?Kz>�H�>�����=O(�>�1c?�&�?N�o?A��=W6?H11>&,�>� �=ʚ�>�>�?sO?��s?��J?��>�>�<�᭽w����o�pB�[X�;@�F<��z=��V�|�9��C��<���;�@��غn����F�ȕ���;LU�>u��>m�H���������=ކ�>K�W�� ����
��T��$A�>�"�>P�T>�����㽫-�>���>}Y�@?,$?x��>��=�`�jrN�X���(?�3W?��3>�S��>��(e���r���q?tIJ?�\Q��&�7B`?&c?��ݾC�*�U*��������⾴�S?NO?$M�p��>Șp?Ugo?V?u'��A_��u��A,v�艍��)�=���>�M'�FZv�羂>4:5?-��>���>l�>ii���D`�x[��T?~��?�d�?��?�9B>�fw��]ܿ�r��RI���^?���>�2��]#?#��%�Ͼj^��\&�������"��~T��fw����$��Ճ�L׽�=Y�?Vs?�Xq?��_?�� �d�c4^�����cV�&��!�r�E�8"E�e�C�/�n��\�9�����*2H=y�?�ԥA�W��?;M?\N'���?�l̾�������'�4>�'�������ᅽ�ɀ�-�<� �=�{0���>�����B~?\�>�U�>�J?��|��zG�42C�яN��\��>E��>�}�>c�>�8>��Y�0k̽�X�БD�Ο);��>&�_?�LT?ۨ|?��׽�G�������"��s��K�$�#<����=k	>X�Q�2���"����=(s�e��6&i�����$�בl?��>'$�>��?�@�>i|��gžR���R�v�W>v�>.�a?�ʤ>�=�����������>>�x?|�?W�b>�k��S�K�'I�����>���>�{�>�!�>x݌��<Z�ĕ��wJz�.�!�q�=
�:?��a�D_����*>�Xm?�����,d=X��>[*��<��Tž�}�])>��?R�B>��=�L�J+�'����s�{G)?�N?�Ⓘ@�*� ,~>"?�~�>�o�>�'�?�>	YþO�ǹ"�?A�^?NJ?�/A?��>��=Ф���Ƚ��&�Z�-=!��>�![>�4m=��='��p\���ԙF=a��=3N̼�ǹ�}�<uƵ�E�N<'��<`f4>�#Կ͜T�@��P$��k������ý�N��̓��JЃ� y��l8��.\����%E��zzL�=�T��3��nς��U�?^��?l�Ⱦ�])��.��D[���gm���?�5������'�8�z����zԾT쫾��^��-��~N�>e�g�l�Ӆ'?g���x�ǿX����yܾ� ?OK ?j�y?6�	�"��w8�Ve >��<�(��k������οA/��W_?���>��褽J��>��>	�X>��q>����잾���<��?�N-?���>�Pq�#wɿy���*�<���?��@�wA?ƿ(�4�E`T={o�>j�	?<Z@>T=1�6W�����U�>~6�?���?��K=��W��^��oe?|�<ξF�����[�=6ɥ=it=���N;J>,*�>E�	#A�	�۽Ƒ4>L��>ӊ"���6\^��X�<|^]>��սqQ��a%�?M<Z�)-c�N�*��~��*>k�P?ĭ�>:�=�5?�%B��dϿ�b`�P \?�6�?���?��.?����ܖ>�&߾E$O?9?I�>��(���{���=�6��5�����̾6P^����=�k�>��>��&�h����[����}��=`9�	�ȿy�%�/�#�2�<���˰M��x��̽��͛�| p�J�ѽ;�=��=�6S>pp�>�?\>��I>��^?<cp?7ۥ>(@>�-+��m��j��4��<dk���k �\���A�n⪾���'۾���|���)��j���=��3�=�KR�Y����� ���b� MF�}�.?��#>��ʾ�M�ƙ<�rʾ%l���q���q��/̾�1�s'n��˟?; B?�˅�g�V����$	��{����W?r���������t�=�/��$�=��>ӽ�=-��	3�<�S�$E/? �?�d���:��e�&>Kl �e�=,?���>�I<�9�>j&?B�d��-Y>?�+>Dߠ>�Y�>�t>�����⽠�? DR?h8���J��@��>8r��ʡz�{b=�C>��,�> Ǽ<qQ>�TU<�܊�Ww���w����<��H?n��>��+��w�?C����;.m�=��x?�9�>�d�>l�R?�N$?`@>Z����z_�W9#�aߜ��q^?`�t?˃*>�B��pNо��W�/a1?�oL?���>�hX�� ܾ��!���龗(�>��a?u�@?� F=e$�������_���??���?��i��f���&վk�?��w?��>���>^�4��߭>`a�?��z=�)���5��P"�~ة?�"@tj�?��j<��R;������>S��>����q7�������&Ƽ��?�o��ʀ�JcE���.��^]?E�~?#��>>��� ����=
:����?̚�?bĥ�^t�<���<l�Iu�tǉ<��=���	NQ�#(���6�,n¾��M�����"!�>C;@���+p�>'G�oh��οT�����ɾD�m��[?�͢>"VȽ#ؙ�CPj� �q�WB�G�F�Ӛ��Iڪ>K{F>F�&�T�b���n�L2E���A����>�v�粆>G�������B���K��<��>'��>)8?>�3�g�;���?k�꾒�ѿ�0�_T?���?Eȇ?) ?��c�t�A�U�/,=s�\?d�?a�e?ZQ�W�J����[?�{�Tv���7��J����>�9?���>[:�Q��r7>ԗ?5��>26;�@ڿ��ҫ���Ҿ��?E�?�����>�{�?�D?d��a��@y��6��aPv=��%?�>٣���i��z6�ak���6?�s?���>��]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?���>��?���=0$�>�X�=Go��@�Q�$>�?�=6�>���?�$N?��>�s�=��4��.���E��;R��� �C�$��>�<b?��L?�,d>���6�(� �	�ʽ�0����t?�� �@�߽X�4>��=>B�>@�E�DҾ��!?˩���ڿ:��8ȱ���[?!1�>C�>�4�����l�E��fd?b�>?���]��3ߐ�C�$�6��?�5�?�W�>�˃�(��QS>駴>d�>�Y@���!�ݮ�ɩ=`:?����>���q}�̜N>\��?,��?�+�?jyZ���??��zc���c���վ���n+���3 ?�@�"�*��J?q��>��z�ss��yO]�H�?�?��?|&�>�$�?�"��DMD�5t�>�	�>�̙?lA8?G�M���:���>�h?Wq��* �������?��	@��@ug?���8濳w����������%�=��=I�)>s��b��=(�D=�.���2d<1:>�&�>W�i>{po>�q}>%�6>Ȫ'>�����o!�M��� ���=3��5�����ivz�9�Ԭ���R���־���m�L�#d�g!�<I�'�>�{�=[�=sB?`�Y?; z??�B?��8�>+���ψ����>��V;f�=!��><�5?ћ_?��U?���=
#����l���n�e�̾kɱ��-�>�2�>�T�>0��>w>�>E��>�hG>��K>��=�4�����'uT��>>��>���>Eh�>�@<>�>�δ�w1����h�Aw��̽� �?_���c�J�Z1���;�������n�=�a.?z>����>пa���K2H?K����'���+��>W�0?ybW?Ҟ>&��&�T��6>���f�j��]>!. �ǁl�֎)��&Q>�l?�/>KZv>~O7���2�]��ھ�/�>҆2?�BѾ���8�_�.U��ྦྷ�r>>�>Բ5�.s�c�������P4I�i��=�~N?�V?U`����������.���t�F>�>>���'n�=3�O>["���l�1�f�㼭�=�{X>c�?�$4>xv(=��>j^��{�2���>��H>�>}�;?�-!?`�Ƽb'�4̊��>��V>'2�>4k�>�>�Y�:r�=� �>��M>�K(��ۨ-�;�,�8�T>w�{���y�Q&��*�=|½4l�=���=��|GC��A=�~?���'䈿��&e���lD?U+?� �=ҝF<��"�D ���H��E�?q�@m�?��	��V�>�?�@�?��P��=}�>׫>�ξ�L��?��Ž4Ǣ�ɔ	�%)#�hS�?��?��/�Xʋ�<l��6>�^%?��Ӿ���>�ѽ��6���
���(>#�%?*]?�<:�oTO�����n�>�?e���������пX����*?�?�ȗ?A؀���& [�C �>D�?��W?�N5���@N)�t�c>��+?��o?E�>�V�5[s���?���?+��?]q^>ƥ�?�y?D}?�:�=X�H�x��u�s��">j��=WJ
��$h�!Ȼ��0�qj���q�c]�X�3����=�=XY�>����������=DF����c)>���>�l�>?Jd>귔> �?�b�>�r�>�}�;&m<�a:G�"ř�|xA?~��?DM���h�s��=�G��@#�	*?Q�M?}��C���M�c>	D?1Α?��u?�Ǟ>�ߝ��L�����̾A�� $>=��>�g?��μȤ�<��^T��|�>A6�>PN>����j���~�<�	>�`,?�>?zT�>�� ?��#?B�j>e�>�`E�6��J�E�ݴ�>���>�D?��~?,�?�Ź��Y3����+䡿[�[��KN>��x?�U?���>z����z��"E�*]I��쒽���?qg?�q形?�/�?Xz??͖A?f>�d�K�׾Wn����>��!?���A�&J$�49�jR?�K?��>U5��K�1��>��0s��.?4[?��#?����`��g���T�<���ԡ��ǿ;_�Y���>��>��q����=\>]��=�<j�H�5��h<��=�~�>P��=�}5��ʍ��o8?����<�8��ϋ>>f��(���.>Qⲽ����+�?��7�α��h���G�=Y�?���?�%s?�|���~�\EE?�a�?_w?�~?���ʾ�Z̾b�� ����>�B3C=3y�>t�����*�Ho���t����u�(ۘ�+� ���>TB�>��?��?5=>t$�>l���d�Jy���J�}�s��/���F��=&�w'�o�j�������^��gP�����>ac۽۶�>�?�~'>/��>��>�%�<��>��u>o�>��> JF>�Y@>�
�=M�S;�$��iJ?�䕾Ϫ%�g2ӾȧԾ�2?i�j?	�3?d	�����	���-{?��?`��?w0�>]l�`�1����>��?^���Dd?�|
>{���G=��ɾX����,��һ<���>�F��Z)��6�jEZ����>��?�h���精������yo=M�?M)?��)��Q�߿o��W�.S�c��ph�F{����$�v�p��ꏿuZ���"��u�(�`*=Z�*?�?|�����&k�?�Lf>~�>�&�>��>�oI>��	��1���]��C'�`���O�>hM{?���>��G?G2?�G??)m?���=p,#>�����!?�+�<{�>�-?h�6?�!G?�*[?�?�M?-�x:X�U���������:?޼&?�e%? v�>
n�>Vb���F<(��<b^��vU��s>�a#=YzJ<����[3��d��:>(�?�y�=o7a�iӀ�D�� 8 ?�)}?ߝ ?U���پx&��3�=1'?¦e=��|k��Q��]�>d��?3���5�=��y>�">�'��i	뼩.�=�>�L�=�I��Lņ��Ͻ�-=c�4>\��>�*%;97��Z�;Sa�>�3O?4�?9�C>g�ݭ>��K�%�y�"��>��>�gO>BZ�&��)��)�c�F��>��?�b�?�&����=�^7>7%�����N���H�<��?�{?*!?�aN?�oF?�?;�=�~���XVBu���>C,?8��>���ʾ�쨿Wv3�ޝ?~�?�,a�X(�t,)��¾�SԽ��>VD/�Y.~� ��@D���h����ј���?��?�)@���6���辫���$��!�C?��>�/�>��>ȹ)��g���.;>I��>��Q?{�>��O?�>{?�[??�T>"�8�>/���ϙ�BZ1���!>�@?���?��?gy?[g�> �>ҵ)�D �BW��i��(�]ނ��EW=�Z>%��>�%�>J�>���=QȽ�~���>�f�=�b>ׄ�>Ð�>$��>�iw>`�<u�G?���>NM��R��,��Ӄ�s�=���u?	��?>�+?o�=>����E�^K��S-�>f�?{�?+2*?�S�,�=�I׼��i�q��>ɹ>��>a`�=a|G=k>>��>���>v��{�Pu8���K�Z?OF?�P�=��ſ�Bq��Ur�������:<���c��5���g\����=0��'��੾�Z�4-��߮��)��{Ŝ��}��/�>��="��=p��=���<\�Ҽ(g�<D�K=�Ԋ<��=Y!p���`<us;�'��������F�z�I<��H=����f˾<r}?�KI?ڶ+?C�C?�@y>��>w�4���>^ɂ���?��U>�rP��;��58;�ǐ���&����ؾP�׾��c�����TU>�H�S�>J�2>q�=�=�<W�=��t=t��=�EY��=���=m��=���=���=�>�B>���?X}�*+����'�U��?l�?V�>{�f�����AU?�	?�i�J�˿�/���?�c@+�?�?���f�=>�����z8=��>tG"�Ԓ]�K`�=����(m�>�R�>��~��ѷ����=�/�?Bi�?��D?"|�_@ʿ�>>��7>�j>��R���1�ޅ]��@b�ͣY�ٕ!?�`;��>̾5(�>�Z�=Z�޾��ƾA�*=�5>�a=Ϋ��\�}G�=��y��j>=�wl=O��>��C>���=\��cj�=�`J=te�=rAO>����8�7�=�,�t�1=�=�hb>�.&>��>j�? `1?:Ed?<7�>�/r�P=Ҿi$ľC��>���=�۱>��p=;>ҵ>�p6?�	E?�oL?�۱>��=�=�>���>�F,���m�A��2���\J�<���?�և?���>U�x<0�A���lv=��^Ƚ��?�=0?�`	?�2�>��u��3�݉T����o�<������ľ�bk=�[�g2������>f'�>ԗ�>&Q�>m�>I�b>�a�>G�>�>�C���s=�l�9���� ߼H�V�:���=7�<$ꮼ�IY�������ͽ�?o��?E��G��yp�x>���>c�/>-J�>sR>q7�����=�����>�t{u=y�ܾ�Zq�<⇿�璿/
������F>��v=l��߲��F&�>�K>ш��A�?Nj?Pe$>a~=�c�==����a��_O��Ĺ�X�0��(��5`����"V�|�����>>�>sԢ>�fl>�,��?��
x=%��T^5����>#z���������.q��8��n�i��P��	�D?N@��&r�=�~?ȈI?>ҏ?kH�>je��^�ؾ�j0>?/����=���\q�#\����?�'?~X�>�
�h�D��*��`��>q�>�j��L�"���R�<���:����V�>�ݐ�Ϋܾ��,�Rۃ�⍿H8������_�>�D?z�?L�v� F��Km6�����1��A��>/�G?<B�>H��>�a?TG�=���޾�۫<1ƃ?I��?�}�?Q�=nJ�=���a�>�J	?aÖ?Z��?=Ts?�?�#��>�Ȉ;|V >�z��.��=��> >�=i��=�g?4{
?E�
?�ڜ���	�� ���h�]���<v��=�s�>�,�>��q>i��=�Xi=�֢=eP\>���>�̏>ܻd>�ݣ>�=�>q吾ʅ�y3?��=���>
8?Y�">5,�=0�3�[<�!���z�䍵��a����ǽ���=-�2�əF� �Y��:�>��˿���?o >���?����/=�ô=��>2�}��}+?鍾>��>FU�>���>��F>��>I3$>��ݾ�A>�	����:�M���]��˙�n��>��۾Ճ������@���E�1�����B�j�Rv���.�ǨT����?�Q��C�V� %�IbX���5?m�>h�H?*��*|M��x=�="?$�>�����z���~��?�z	@��u>���>8�w?��)?^��o
W��n{�������8���9���5�?������N~�����Qa?�?(�?O��,>���?T#�JQR�4|�=�aj�d/��M��1?)H꽙�C����q��o�<�ߘ=�e?Qp�??Arv�K��$�B�f?�d?,��?^�>h�J>�8��S�~? �l>���>$E:??/	d?ݐ&?$X>�u>��&�5� ~�����>�Q�`���c�j���>#W=�7������=�����==�� �Q��6`�"䇻��	= -�=Bl�=�Z�>��a?� ?�(�>w�4?i,E��>?�[A���90?��=4�r�a���R������/=�=xj?n��?O4X?	G>��?��k1��J>$	k>H�>�?>i_�>�wŽ��6���=]�=R�,>�P�=P�Q��G���<��Q��� =#�>ŷ�>X�}>���r&>�y���qz�[\c>]YO�������R�hpG�2�|kv����>B�K?�|?�<�=b�辷��hXf�I)?�<?J>L?0
�?�=��ݾ��:��I�=��&��>E~�<�T	�hע��?���{:�m?�9�Gt>�����,����f>Lb�tJ���o�#�K�0���gc=4L�/%J=�P���־�|���=wD>C��k/!�_֗�t��h�L?d9�=
N���\�����'�>6�>�ϰ>G=T��h��GA����q�=)�>l�?>����W��o�G�ϗ��i�>��B?nVg?�x�?�h~���{�F�?��a����Dl<��?g<�>@?W�+>vzC=������v#g�'�?�*�>`%�>���1�P���������>���>m�=�w?ER?!

?C[?��*?<��>�vP>�Q���3���C&? ��?ń=}ս`�T�2�8�dF�%�>��)?�C����>�?$�?��&?��Q?D�?.�>�� ��C@���>?U�>��W��e��:&`>*�J?6��>� Y?�؃?��=>a�5��袾S���!��=�3>}�2?LB#?'�?}l�>*��>S���<�=̣�>�c?0�?��o?ʇ�=��?�62>��>a	�=.��>���>�?tWO?=�s?&�J?���>G��<>���<���Fs��bP����;��H<H�y=`���+t�*����<�;�j��+��j����D�OꐼB/�;�n�>��>��z�̹�=7�ﾾ����n>c)=u����#���]��;FR>��`>ඛ>0�A�K_K�&�C= |�>��>H��Gk	?4
?j��>=VZ�k�C�R��v�?Z�?=�f>*�b�ZD��Io����=�?Cyy?x�]��;b?�s?�о��'����]��L��5+�?Z&?��̾K�U>mk?�8t?�6?���/gG�m������]�Λ�=��>x~K�h������>�ZX?r�>W7">F"�>����q����c���&?r��?��?xۑ?�U�>	�e������lڑ��`?B��>[����?"?��n�\ξ�d�����U޾)P��<����ܙ��%��� ��f��"�� �=�`?r?=�r?-�`?�2��e�O-_��G����Y��L�f����F� SB��@� �n��\��3�v���Ci=�wV��\?�ˀ�?s;?.�ͽ� �>1L��{߾o��l3>�6z�ǟ"��Z��#�:�B��=�A�=?I��nl����P&?J=�>c~?|�<?xni�\>K�Ȯ?�b18�5�1�o�]>D�>�Hc>�n�>�7R=����^������4�[�Oۼ�u>Uc?�K?�4o?'<��i1��n���*"���,�uw��~4A>{r	>�m�>X�-*���%���=���r�S��괐���	�[c�=��2?��>�ٛ>�>�?��?~R	�I®��nx��a1�fA�<��>��h?�W�>v�>2�ӽ�N ��:�>)J^?�*?��?7#r�#9���n���ʾ���>�)?ŏ�>���<w�"��H�� ���Lj��*��.�g<|�)?���2�v�X*�>�_?���<J������>Fq>�ӿ�풑��G� �'=c�?��=�>$�Ӿ
D�k^�� �ѽUJ)?�R?�ג�
�*��x~>N "?a�>��>/�?RD�>OOþ���ʷ?��^?�?J?DA?�=�>N�=cg����Ƚ��&��-=@��>�&[>E�l=/�=����c\��(���D=��=�A˼61��/�<$f��X�L<m��<�g4>�׿�=�����z�����n�8Ո�T(Լr�q��1��#�����]�����'<��.�\B2����˸���I�?r�@7d�����3P��ї��R��]�>~�����#��1��O���:�����ݾ�9��8��qg�����TA{���?<Ol�D���U��{�Z�~]??��l?9��?�p��Lk���i��ɹ>�=��'>=\����i�ʿD�5�y?���>2�����^�>ݻ�>O�>��7>D���}�r����B�?0�*?���>� 	��Q��{)��g-1�+��?,?�?�{A?��(���a�U=8��>�	?�?>QO1�K�S����R�>�:�?j��?�`M=X�W��	��|e?B)<��F��ݻ��=^9�=�^=���l�J>�W�>h���SA�8ܽ��4>�څ>s"�����~^�j��<b�]>P�ս8��Bq�?�6V��V�H��'O��f��>ϫA?��4>l�r=�b?U���Eݿ`�o�x�B?+ @���?>�<?��ɾ?-�>�����[]?��I?�>�>�%�z�����>M����r��E[�e�~��xt=�k�>;H�<:z���	��Қ�!bz�jm>���$ȿ4~*�C!���j=��̻�2g����o��p���︭�[�������&�=�U>��T>=�>�a>�2>��d?9�w?>e�>�>������Q
ѾN?,=Y	P�UIP�9U������F��QO���վӭ�4�QO�k��<��o�=WTR��Ð���-��n��S9��{.?l>�˾��P���ռ�ѻ��u��٦�;�/��2Ծ�B�!�w�/��?cM?������Z��|'���7����;��V?P�/�4��~Ⱦs��=!ر<�3�<T_�>��k=,��G<���I� ]0?�o?���޴����*>H* ���=z+?�W?$�j<%�>�7%?�)�z���Z>33>*��>r��>�3	>t��/�ܽ�r?خT?T9�r���|�>�M����z��:c=�G>��4��J߼*I\>Y��<���YU�偏�	�<v�D?̳>K�6���0��j��u��<6�4=�)f?p!�>8��>-Q?�-?�l�=x�HLc����+<+<�a?'jj?R.>zJ�Z�7�C���(?=�g?�r�>a�9�Ȕ���Y־?�5�?I*(?�$� ,l�o���7꾛�.?ݶw?�^�@�����U\[��>C�>���>S(9�`X�>T�E?�,������<��sf.��#�?��@���?9�<`G���=;4�>dB�>iH��ձ� [ɽ_1��u�B=h�>�|���w���#�#`�3�=?�g�?�� ?hǁ�����=\ڕ�]�?��?5x��3�e<1��bl�����,�</ӫ=ެ��'#�����7���ƾ_�
�!���>F��_��>X@T'轜:�>yc8�14�8PϿ����Xо^4q���?U�>��Ƚh����j�S;u�ÞG���H�h���졣>��>卍��V��ٽ{�g<�O7��A��>_�	����>�{P����1���U(<ET�>�[�>��>�A��*��G֙?��~�ο������X?���?�%�?� ?T��;�x���r�J���G?��t?k1Z?�6���]�	<�ƻG?M���?�]��-��`T��zk>5c?���>X;I��S˽�F�=>?OaN>
[ƾ�º�Q��3�&؞?%5�?~S��?˓�?�4?�Yݾ�<�����>��9>c)?MoX>��������f��<Ҿ|1?��M?�ŧ����]�_?+�a�N�p���-���ƽ�ۡ>�0� f\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?X�>��?��=�i�>���=�9��d�G��>[�=��,��9?��M?P��>ٟ�=O�4��_.��RE��1R�l?�H�C���> b?FM?�Fe>q���8��+ �gɽ�.��L�R�<������ܽ�i8>pt<>`.>
	C��'Ͼ2�?Hj� �ؿj��fu'�#24?���>p�?���w�t�I��d7_?�w�>�6��+���%���L����?�E�?�?;�׾,�̼}>��>DK�>�Խ���������7>�B?���@��;�o���>%��?�@�Ӯ?i��u?Wþ@q��OI��������H��)�1?�����3>}�X?�'�>^||�u྿�#A��?��?y�?��>��|?ꄉ���h�������>֐�?W<�>t޽>��1>�8?,v߾Sm��Fxھ�j�?hg�?�@	�m?�������س�� \���%��l	�=,�=�.'>�p��EY=:��<d����Yt>�ԝ>�.n>��i>\Z>�,I>K�->AM���K�)o��ێ���3����n�����Ap���$��ǩ�n���������&1ʽ,W��c8�U4��ф=�<?��^?E�O?�8<?K� <�؝��Oʾ�%�>�N_��d�=bN�>v�X?�m?k�2?��=�Ch��r�;jq�g�۾��̾��?���>��>�ޱ>`�)>eo=��[>�g.>/��>�}>��_�=��P�@�	%)>�S�>*1�>J|�>uP�=��v>�R��8ⲿ���x���w��=��?/��@�:�U✿s���7����w=��/?R�=s����ҿ����xll?����PW�]�d�#Τ��N?�q?��>}{ʾR�����=�<=!k�S40>v%�?�����=�a��>V�X?�f>�u>��3�ne8���P��{���i|>G36?�趾�C9�q�u�p�H�Gcݾ�HM>ž>�D��k�a������vi�:�{=ex:?Ԅ?h4��sⰾ�u��C���OR>�;\>�X=�k�=SYM>�ac���ƽ�H�#i.=���=�^>p�?��->��=���>� ��T�v��>�Q8>J�,>�9A?��#?�Z �Ş��Ń�B2���u>�w�>/�~>{>�wL�א�==�>K�e>O���(������C�yV>Ozn��ja�5}�}��=�������=^W�=�	��pA���1=�~?���)䈿��he���lD?[+?� �=/�F<��"�E ���H��B�?o�@	m�?��	��V�A�?�@�?+��G��=}�> ׫>�ξ�L�ޱ?�Ž8Ǣ�Ȕ	�)#�fS�?��?�/�Xʋ�?l�{6>_%?�Ӿ���>OV��ϖ�mU���[d���L=&ښ>hO8?���5=ʻ�@��s�>���>����쥿����	j���?=��?&��?�[������*�8��>e;�?��d?�~>3��y��ڠw>I�??yo?��>�h����i�?��?�?i�,>x��?Mi?���> ����5��~��ꈿݲ�<:��<��>!O=��ľpyA����g����c�_����t>�o%=�ĺ>B{��ھ'd�=4�)�ĵ����Y�1�>��g>�#9>��z>�C�>GJ�>�x�>]�W=�;��P)B��Ϝ��C?��? ��j����w�=rT-> ���>s`?�5�^QҾ�3�>��]?�F�?��N?�+�>ð��l���z���u⾇Ǽ���r>�n�>a=?\�V;�8=�M���˾#�?��>�XC=����~q��q齞�>��G?��?���=[�?o&?���>��>a�C�����7�Kb�>�&�>�A�>h5k?��>-t�� �$�����.��6�j����<L�`?��6?�i�>�}��<'���l�-��=��滌�?�_X?�X��3[�>���?w�U?�]L?��>�U��>�����X/~>��!?��1�A��M&�Y�x~?�P?���>9��\�ս�Kּ��������?�(\?=A&?����+a�m�¾�8�<��"���U�C��;ÅD���>��>}�����=�>�װ=jOm�vF6���f<�j�=��>%�=[.7��u����3?[s¼�X�r�>��o�bQ4����>|b�<�־�gؑ?_�^�[����,�� f�<�a�?��?)_?�!ҽCs���}N?)�?�R$?Ԫ?�㾆+���M���/l�j����Y(��`>g_�>GU�R�&�U���낦��/n�Y�~�o� �?5 ?���>�T?�?�G>2?�>�Ӭ�X��M��:���Xl�b�.���C�����������V�3����ϾT����>�d+����>�g?�6>\5�>s��>���*��>��>�3S>�|�>?r>�>Pػ=�<�۽�KP?Y콾�:+���¹���QC?��g??D�>�����������!?��?*��?��\>�l���/�P?�u?����A�?�%=�Ј�7Y=�纾2���`��%pV��*�>�玽�4�c�J���S���?�<	?�׀��W��]k��ə�/�=|�?V�6?�����^���i�D�]��I�~�<�i�Ŗ���?�a�j�+p���������-���=/�&?�g�?\� �Ld��(ľ�ec�m6���>�W�>��U>kd�>X�K><-�{�)�vO�-�-����X��>*�x?���>��E?�X.?�#?��_?~�>;�=>)�羚+?�>���>�?4<T?ZL?D�:?�j�>�?�R�<`�3�P�l�꾅�.?�s7?�B?�9�>A\�>��n�B=r�����Խ�!�6>T�=�|�=Fs4���x�IO̼&Wz>��?L-�=�{g�Ӝ��$x.<��?P�f?H�u>��J�rF'�n�2�J|�>q�?y0�>�;��w��80)��I&?�1�?%%��ϡ�h�;>��y>HgC������S>���?b�C�b�~�����=U��S>�^=�e���켩�ʽ��>{��>�T/?���>�d>и�iw.�)�S��c��pJo>��!>��V=R��T-�������pf�R��>���?@a�?��S�='CB=��m��U8�̍�]x���=d��>|� ?Kia?a��?� !?هN?A/k>X���H���E`�=��?�,?딑>	��1�ʾ�꨿�w3���?fY?�Aa�����3)��Y¾3�Խ�>`m/��=~�:��O�C��^���������?۱�?+�@���6����`����E��v�C?I�>�&�><��>8�)���g�T�;d;>di�>��Q?/��>J�O?Y{?��[?��T>��8����֙���)���">Y�??`��?ߎ?<�x?��>��>�)�c@ྊ=�����a��9�����V=@�Y>?�>��>��>g��=�oȽ�寽(?��U�=8Nb>ki�>�@�>�@�>�w>�Ͳ<8�G?��>�پ��R���������$B��{u?5z�?>+?a�= ����E�İ���.�>�Q�?5ܫ?H�)?!GR����=�+ܼ������q���>�>�S�>gI�=;P=�>���>��>T��,�^D7��O=���?�IF?M��=��ſ��q���p�<嗾�mc<����4e����s/[�x�=����
��?̩�X�[�t֠����k���~s����{����>�͆=@�=�A�=ʗ�<Lȼbܼ<��J=��<�=�up�%�j<R�8�1�ڻ9����D~^<�fJ=�F���|˾Wx}?'I?��+?w�C?��y>�v>/ 5�	>�ك�80?tU>�	U�{Ѽ���:��c���ؔ���ؾ~�׾�7d�[���8>��L�W4>]�3>R��=�Ћ<��=�ir=�Ï=WL"��*=1_�=��=t�=���=�>#>��?n����!���"G�L�^����?������~	��G�?��4?�4d��*ʿ�!�A�?β�?|�?�?�R��w�y>�#���H-=�(=���e�=0�=G����>/��>W�4��ǿD��F��?mI�?hY?R��W�ſmx�=�-5>�>��R�i�3�w�\���a�_���?�;�_
ɾ2D�>y��=a�ܾ=A˾F�<�i->2�N=��
��LX�{��=��o�pP=G<[=i��>�L>��=i���aW�='?e=��=��T>T�e<��S�&�֍P=&N�=�a>+'>G�>��?+�-?��_?T�>at��о/�����>m�=d
�>��=�6>q$�>%q0?y�D?��K?�>NW�=y��>�t�>D-.��j�7�߾�L��(�m�Z �?}��?yŴ>�mY=+:�u�%��0E�~y����?�F8?�S
?��>M���x�$�5�_�*=�K������w��Cr���;���I^���cQ>���>Ǒ�>��>��Q>�A>a�C>���>Q�a>�!�<|w��q�A�<�u<K|D>bU�<U��1�V��e@��#߼�`r<Kq>=|M=���=��b=����0�=��>�>C>���>+��=a;���kk>ޜþ�+/���>���Աg���z��Ň�����XT��!r>P:�=c��-��3e?P�0>�y>?��?�Vi?]��=uU���a�� ���o��%�Tﳽ� �=x6���W���_�h�/��H�Aګ>9ɡ>%\�>��>�y'�eA��7#=�¾�D6����>�i����eq��0a������ad�3�+=�cP?�}�����=�=�?,?"��?Ъ�>-������z%>>�:����=�X:���x7�r�?�*?���>�ž�S���¾�q����>����M�H�G�����4���g�ľL��>[;��LU߾� -����`����|D�0|�@V�>n�K?�A�?�w"��腿6	V�&� ����;�U�>G�W?)�>"?w�>5������5��k�>��r?A9�?�H�?���=r7�=;��1��>��	?�͖?y�?��r?��?�gI�>C��:�� >AB��n��=�u	>�}�=���=�'?�	?�M	?
���V
��	��b\�,��<��=3�>�ш>pr>���=�<r=W_�=h�\>Al�>��>c>���>r��>���_���"?���=���>&G7?�C{>;� =�׻Ԣ޼r=<����派Kfo�zs<*�=ͫ0=�(���A�T�>�ʿAf�?2_J=���fy?=��R*<q"F�ꔎ>��&��?F؄>�y>.V>��|>�'�=�I>SD>ӧξ�G>z��]�&�DVJ��FP��;����>�K��v�,����������C��#��h8 �JRg��.���@�p5�<䰑?��Z�i��&�����3?�հ>�7?�a��µ��"+>���>��>�.��f���܌�z徔��?8��?�/n>���>��y?Φ?>�$�WY��(�x��⃿#>�1#��}5�����򘒿�� �huռDf?a�y?FB?�H��>�Y�?)�(���U����>��=�}�?�2���[
?(���[B����þ'�0� ���=}Nf?u؇? �g?6���מ�K��li?�$�?r�?���>W�>&��=r�h?�#=
�+?!�=?�D?��\?�o%?�)3>޸=��J��`��;�����=>i�������������=8n�< Ȅ�8�:ѽRX�����r=[��p���`��_>��=|��>B�]?�?ݡ�>��.?tp����S��վ�k"?��;=NV���j��)_оx��̙=<�d?�x�?Ckb?2ȸ=�$E���K�{><q�>G �=�H&>U�>!��"�����=O<�=�>�N>�+��I&����������E��_8!>���>�_|>�k����*>�?��ٯz�#Bf>�*U�����4CK�J�G�\�2�ށz��ݿ>�L?�W?�.�=H��.=����g�ԡ)?#<?�M?��?$�=�D۾Щ8���I�P^(�:�>�Ů<8@	��������k�<�'cr�;�q>�v̠�wfb>�e�^ݾknn�.<J�#���I=nT���X=���վ��L��=Ѭ	>i���O� �/���ʪ��J?nk=|U���
V��G����>�W�>��>�:��z��r@�񩬾�b�=8��>�
;>k|��c+ﾳzG�w,�o@c>y9>?�;o? _�?�X��:��#J������;��l�<FK�>!bX>���>���=�O<��׾m03�x�s���K����>��?�=���u��ej�yԯ�L��)��>�i�>dZ�=O+�>��;?�"?�]v?�GL?���>�>��u�����#$?׏�?���= #н����,#>��7��?��3?�Pؽ"i�=G�?V*?O<;?��_?e|?���<�>)���U���>��>Y��~���x>��Y?��>�XY?Vǈ?��'>{	2�h(�����<*��>5c>lzG?s�3?	�?�q>���>�����C�=���>��b?�1�?x�o?c�=��?�1>���>���=#��>f�>N�?ISO?��s?��J?#��>\n�<���tU���\r���R����;QGH<z�y=Ѧ�<t��u��K�<�V�;91�������^�D��T����;7��>��>���.�=ޚ���l����=ס>�ƃ������L�c8=���>5
�>?y�=��O��Q=�'�>���>�u�?�v&?z��>da�=/�s��;)��3��?fe�>�|<�L]�ڥ��Z� �T>�G}?�]P?�����P�\?�Fd?�Ծ!&�c����R�����?L?�g	?O��~n>�n?9�m?�?ĳ�}�d�1���r�x����;�=f�>)�-�w%w����>��C?W�>���>U&>ɢ¾:�|�wq�� #?|k�?H��?o�?��Q>�tm�e�ڿd��	@��Ĝd?6.�>_\��g� ?~1���پ��qYy��+ܾ�S��kI��<�������S�x����f=4?��l?|�o?��_?���#m��d���{�g(Y����P4��M��=�&�=���l����?!ྤb����=�al�/�I�M�?�b%?Ou�����>��������n�|>;���x�j��A��gj�w#�<��==��D���龏"?���>h>�>��=?��s��hY���H�'51���4�Q>1��>"�=Gi�>�(����n�/�Y����h=b������d>�XW?��U?�?�1��O�:�x�'����,=�Z���>Fp>�v>���.�Q�PU�,���i����Y������!�<�a?$�>�%�>k�?�%>��(��7�9����C4�Sb=>tZ?։�>��>Uჽ��7��1�>��h?wO?(5�>����K��넿�����?\v�>p�>���>C�?�%a������e�W��Jj
9!�I?��d�����>�N>��t?��W�����?ؐս�M3�X�����'�h(>.?,�=��J>T�'��Va�X.���}%??!F��x+����>O>?H�>F��>X�?nq�>W�¾ڿ�f�?�e?�H?~�:?�.�>�T<�����߽�{C�{�U=3�>�y>��I=�d�=���T�H��/��=���=)���8Ƚڎ<��㼲�><��=�;Y>���B`�F|;��oi�A��נ�\�������ޟݽ�6���}����f�����߻��>�� ������f�����?�y@`B�����ӻ��L����|��>b��?�]�����.���ʾ����L��B�PT��ل���L�6�&?�����ǿ6���Y+ݾ�?k! ?ڂy?����"��8�n!>'E�<y0��Z��婚�cϿok��K�^?�Y�>RV�q���W�>�>5l[>��s>u%��Y���7�<��?�-?[��>͙r���ɿ�{���I�<��?~@�yA?R�(��I�7pT=sn�>��	?V�?>�0��6�c��g�>�G�?��?-RJ=�W�1���ge?Ǣ<��F�� �05�=g��=a�=xV�\!J>�.�>CG���@�>Aܽ7�4>���>�"�m���E^����<>]>;\ֽF/��=��?�%O�YL����E����Xd>֍A?P̒=�L=�M?6�	��q׿^�����P?i�@�`�?��X?�Ǿ �t>�
޾:RB?$8?>r�>B�(�U�n��;
>��%�*�Խ��I�����G�C=W�?�w}�N����A��L���GD���->��4hܿg������=�=�đ�K�Q�H�̽�����y����)Oz�������=�^2>�%]>��>e�n>�eE>��Z?�+y?��>_�=�6=�L����ݾ�tD=(�����!��S����]�8˨�2m��4辀���5!�>D����V=��ō=�R�˔��s� �-�b��F�b�.?5"#>ȘʾM�M��4(<�oʾ�Ϊ������즽��̾��1�On�)�?�eB?�� W�BK����X�j�W?E��}�5������=����|=l|�>�K�=���d3���R���?d ?~@���r��XD������=G?��>irz�I�>��I?�:��zC��V��;>���>�n�>f��>��Ⱦ>/���E?$�)?����վ]a�>������w��<��>"����U�;w��=������nY'�|?�hς���J?�}�>,�-���-����� 3�=6kh?���>
a>yKf?�B?�t=�� ��U����Z8<A�T?|ah?��'>��彠*ξW��H2?sYh?ˋ�>HR������6^���:?Op?i7?�L
����Տ�c�l�6?��v?�S^�-��/��I�V�;\�>ҏ�>� �>��9���>D�??�D!����xk����2�L�?B�@�{�?'#+<���҇=��?_��>�kN���þ}'��=���o]k=���>Rݣ��vu�PZ �2�(�/�8?K��?ף�>��������=w㗾�?"�?KZ���g<^��HGm��F����<��=��u�=�N�6��KS6�*����H���������>��@�����>Q�H��a��Ͽtz���EʾS�s�\i??S�>M�̽a"��P�f��_p��/A��rC�5~��G�>�!>:���Α�\�{�BY;�����4�>E�����>9!S�x'�������c.<�+�>��>z�>����W��?�k���&οv���F{�4�X?�e�?'�?l?�hE<��t�t`z�E�9���F?��s?NZ?�!���[�Ǖ<�Υg?����Vd��/��(G�]�a>�_/?1[�>�J(��*�<E`#>�1 ?�S>�<0��z¿{>��D����(�?�f�?M)���>eE�?�0(?��^������� )�Y�;�:?��2>�4¾�{��A;�([����?IF'?���X��]�_?+�a�N�p���-���ƽ�ۡ>�0� f\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?W�>�O�?�@�=�Y�>�2�=9=��Բ��3>�^�=GW��?h&M?���>e�="�F��V,�d�C�Q�M�"��ykB����>�9c?V9G?��f>x,н���#�%�N콄(3��z���Q�i<��<佩�/>�/>�' >l~G�׾d#?���rڿL䨿��i��C?��c>E�?8����ɾ��=C�?�w�>�>�g��*a_����?�?�r�?&g?ZӾ����M��>N		?�ݘ>\����>B���?͒�`�Y?u��=Q=���3B��~�>�\�?,	�?[��?�IH��1�>�&��߫_�5�]�4���G��4�=�d)?.���n�=w�>ͷ�2�������0!��;�>cӲ?�/�?Hb�>Ϭ�?Ln�a�P�r�=xV[>�.�?��4?��W�Ԃ�RJ�>��c?�i�����#����?D�@�
@��r?ԑ����鿮:�����������>�=�P�= U�O^�<�9=.�d�!�</>.�>�>/Mp>���>�'J>]�T>rZ��$(��G���슿��A��_�V	��D��@�j�u�j��m:ξ�qž��ļ�<����g������i<�==��0?��R?wxI?�`]?L<���PA�������>$��w5��&�>*>K?�	�?�=?�]�=T=��k���z�֨��G	���p?s�>�d�>:5�>�.�>3��=́�>*��=0�->z�>�X)>!���4��=��>-i�>��>��>yC<>��>Cϴ��1��k�h� w�|̽0�?����N�J��1���9��Ѧ���h�=Fb.?|>���?пd����2H?���z)��+���>|�0?�cW?$�>%��P�T�<:>$����j�*`>�+ ��l���)��%Q>|l?¯f>�"u>+�3�'`8�J�P�X|��nM|>�86?�ݶ�^9�A�u�l�H�VݾIM>���>sOD�-g���������i���{=�}:?4�?�
����e�u�C��hoR>�+\>d=�5�=M>hfc�ϑƽ��G�5�.= ��=h�^>��?��,>�W�=�#�>�d��,]O�]ۨ>��C>t�*><5>?�l$?�_ �-Q��V���U�1�W�s>�q�>� �>�>�L���=<L�>�a>�|��y��@����@�NZW>�儽:}^��F��Vm=�Қ��9�=�r�=�����?��P=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ^q�>�%ż�쓿U(���͂�J�=�~?!#$?|-��N��DT�(?��?* �_���Y@��0!����	?h�?3ԋ?�O[��_����3����>���?q�J?B�">/Wy�԰z��Z>R�E?p�Y?V�>��,�K��(?]�?�/�?% />��?0{?�O	?��[�,D������O���o�=�=[=v>�=~����_D�SX��6��[d�2��'* >QX=��>����о܆=��˽00��e�+=�g�>x�	>]�1>��>4��>~��>��>FZ���
�^��������8?�,�?�Ҿsw�w��>�y�<�_k��3?��_?��+>Zl��mk>E`?L�?�]?B��>_7�����g�¿ԩ�/1���q>��>�?��>h0&=h!�-��`S�>�t�>�
�����9ef���4�OQ>]n(?v�?�&>� ?ќ#?ڊj>�"�>-`E��7����E�$��>Μ�>,B?s�~?.�?�͹��[3����䡿n�[�=N>��x?�U?0>��������E�nI�t�㚂?hng?%<�@?T0�?x�??;�A?+f>l��C
ؾ������>��!?����A��M&�+��}?mP?���>6����ս�Tּ���H|���?='\?@&?����*a�N�¾B2�<p�"��U����;L|D���>�>ӌ����=�>6ذ=Qm�1G6���f<$j�=��>��=c,7�y��(~-?&o�;\��H>�(x��*�H�>Z]�<f�ľ�c�?sW�[�����������:]�U��?�,�?g<�?��Ƚ��k��M8?�ʋ?�8?s�?�?��`먾F�Ⱦ�y����a��$0�.>S��>��&��#�����|��os|�K�j���C�G@�>Y{�>0�?Jl?NjN>M��>b̾����������A�f��$&��P6�t#�j������)�m�c��.Rƾ��_�>�k½W��>��?`�>��>��>/��G��>2۝>KE>g��>��6>�>�,5=�C�<YzϽ�P?S���(�̨�WF��8cA?��f?���>��p�����DZ?�H�?� �?CV>��i��'�U3?�*?X=��=?	?C)C=~;#\{:�4��nP������Jϼ��e>��½Q�5�fIK�ن�ӽ?��?�2Q<)ؾ1������#s=ִ�?�-?Q(���S�m�n��Y��P�%���Gi�롾�#���o��>���ȃ��)�j�
=��(?|[�?�� ��v�n���Rj��F@�b�o>,�>��>���>^�C>����u/�^\�|�&�G������>` y?8��>/F?�H7?��E?' ]??X�>� �>����mt	?��<���>�:�>i�:?�7?��0?�n?��"?�K2>����������?��??5?҄�>��>�jr�����n��qcZ��ļl��=�^O=����q���2��<r@o>\D?��3�=\�NN�T����Fk?�X?��>a+��/;��=�9"?z/%?Ks�>�-�A}��C��	�R?O<�?82"��&�=�z�=f�q>/h#�UЍ�9S`=�;��v���W�=��Ƚ^I*�O��=wVq=$��=��:��ě=z��(��ʓ�>
8?ə�>_��>��[�`�$�]�K�@g���߿>;�#>�	>���K����]9`�M"�>��?�Қ?�V=q��=���=_G��q�ξ�I��Ӿ�ϣ<�g!?�D?p�A?��v?�m_?��?{�=�"��恿&�~��<��7�$?@ ,?Ћ�>A����ʾ��6�3���?T]?�9a����I8)�Ň¾��Խ��>�\/�
-~�*��*D�CT��)��Tw��P��?	��?CA���6��t�����]��R�C?� �>S�>��>��)�!�g�1%��&;>!��>�R?��>v�O?�F{?�\?�NT>��8���)虿}�.��l#>��??+��?pȎ?��x?� �>BK>R *�u0��s������<�s���zW=�(Z>?�>���>�w�>�d�=ߕɽ����?_?�,_�=jb>�K�>3�>�E�>L�v>k��<��G?ǋ�>Z��̃�?�O��uG;�gu?s�?tj+?�=�X��1F�b����>,v�?��?o*?,T����=t�߼6���]q�-�>��>P��>���=:+C=o�>�!�>	�>���^��7��tI��?��E?~��=9�ſMwq�*�o� ���'�f<�M��G�d�'ؖ���Z�T��=����c�������*\�5����������F����|����>�=U��=k�=��<ئ˼}׺<zmJ=�;�<c=eYp��f<W�9�˻tɈ���'��S<�H=�;���sȾ�!u?��K?�]<?��@?I>T�>���9ϐ>�Յ�H�?
�<>�������:�;���������q޾�I⾦af��A����">�5��a>��,>���=�R���2�=��=�8�=e�����<?D�=���=��=�6�=Ĵ>���=��?�|� �����: 7�5SZ?���>�-R�:L���|	?��_?_�g�n�ҿBnо��?m��?-w�?�w*?����V�>�E��IuN�0�=� ��/><�h=�X�)��>�[>����ᨰ��*)���?:��?��;?	�V��ʿ�j4>h�0>��>S�<+0��l��g[���K�F�?�\:�`4پxh�>I��=5�վKMҾ�y�<��+>�r5=��	�`�R�ն�=����K�A=}� =xW�>O�C>�/�=��ؽX��=�l=AC�=�6>!-<Nż���)c�<xT�=/ki>�8>�+�>a�?�x3?�fc?���>�}�=\ܾ�eǾql�>B��=��>v5=��.>�%�>�>4?�D?�L?�:�>�Mz=8\�>��>K,��=n�~�ݾ���+P�;��?��?��>(��;]T��~�TK=�2�'V?^�-?
?���>������ $�O)+�c���ҥ�5R=�c��Mr�,{�Â(�7A���=��>���>vE�>�F>�~=>7'G>�3�>t0>z��<`�d=�n� �<�ћ�{�=of6��Ag<l1м�g��<�:�q�����!+%<R���<��Ѽ ů=n��>NF[>���>9y>����y�>���T.G��U�>>���j���n��v��d�1�ýBo>�/=�g�;��jU?�ِ>'��=� �?�f[?�f'>��_�Aִ��¿j6�_fӽ�=�Bz=꫾4cb�^�s��96�u+�*��>��>�>Zm>,��?��	x=�ᾛB5����>n]����4���q�-��Tݟ���h���׺?D?P:��Yx�=
~?�I?�׏?��>3ؙ���ؾ� 0>�H��!�=����q�v�����?=�&?*G�>�뾏�D��[̾���^�>ceI�7TN��n���0�m�H;�m���#�>�,��0�Ӿ-�2��ʄ�Jݍ��I>���f�e�>��M?��?�
b��u����M�K[�9�q�==?��_?`�>Ѻ?^�?2u����������A$�=�q?y��?���?^��=�x�=����?�>"*	?(��?b��?_s?Ȉ?��s�>�
�;�� >1瘽��=_�>���=�=�m?��
?~�
?�i����	�B����\^��,�<ǡ�=腒>Le�>o�r>}+�=a(h=���=�/\>3Ҟ>W�>��d>��>�K�> ����b�~}2?�&>US�>/�:?��>�mF�� ��<�!���r����$2
�MEl�J��<�55��;�2�,�1�>B�ƿ�;�?X�;>v}���?�
�#�Җ=���>X2���Q�>�j�>w�T>�rP>�r�>��>�>I>����f�6>��� 3�H|X�K�\��.þf��>7A�J%��	��
[ǽ��O��Hƾ����r�����b=���>=�o�?��7=��i���/�e�|�)?��>I�#?`M��&qf;�7O>�n?d8�>���͛���Ih��,��? �?�CA>��>Jw?%*?=C�����!x�E>[A��l0�IY+�n����~���������\P?��r?��?Yu��u3>�l�?dc�����[K>�_D���X�t�G=��+?��Ͼ���H�������A�G�>�Y?q�t?�n6?�B=���[﫽&�E?�2@?�L�?��?�C�>�Z���X?/b�=� ?�4?�@?�-J?<�
?��>p
�=p���A����I����#�fPȽ�����C�=�U�9�Ȁ��
�=-`�=����iP���;��;�p�<��=�|�=X|�=��>'�^?,��>@�>߆5?މ,��<��®�Nf1?9<=�����n��N��Uj���$�=!�i?���?�cW?�Uc>0>�!mB�P�>q��><>וR>5�>�ͽӞ9�H��=M�>�p(>��=�zR�� ���8	�
���8f<t�%>G$�>Iy>�8���/>I=��.�u�$k>P�a�!2��h 5���H�25�UJ�d��>�L?H�?��=�뾤ԣ�Zg�,')?Qm=?�DK?�=�?%�=c׾�c7�V J��T4�0��>g��<~(�򲢿w����K?�WYy��Ym>���7͡��n>f?�.�޾�����Z��6��Ŀ�=���P�=��$�� �ti��NO=1�]>o¾�,���]��� R?�2>I��G�-�n6޾�&�<*�>�Λ>�㋽���HK�}m��n}�=�a�>[;>VN��4��n�N��I#���><[D?1Ul?�S�?��~�TU����N�Q���.��.��?5�>�j�>�)�=�J�=����a�+�Έw�N�.�y��>?�?�])��<g�����_S��?	��۝>{�?�q>f��>4.?�G?�n?��!?�?t�>��o������'?v��?�2�=ص�Z�H���.��>��$?�+6?�x��dS>S�
?[�&?�,?t�V?��?o�=�/$��8B�b�>sv�>��j�����2z>n�\?z�>�.K?�Ts? +>2@7�,���!2�ީ@>��7>�m7?�G.?�	?��>l��>P����A�=���>�c?�,�?��o?���=�?�E2>��>:�=>��>G��>?9RO?�s?u�J?�}�>]{�<H������'s���O�#�;��G<�z=�g�q9t�(1����<*��;�߶��L��a�񼑧D�������;M��>��>2۲�w�x>�)��sA��k3>CK�}����x��7����>ǣ�>>k�>�G�=+ew��0Y=� �>:�>�h��;?�'?��?��>����o4��N��c�>;3?��z=}�M�aD��s|���C>���?|YI?.�6��x7�ug[?ZTc?�Z���H��︾���W4��5�I?tE?3.��u�>�gj?sFo?��>C����O��	��;/��]r����>{D�>�L�!���l�>� X?��?J^�>L�#>�ɾZ���
Zо�<6?�W�?j��?�ݑ?���>��w�y�ؿ�����7���-^?Fr�>�����"?�F��ξ�B��䎾��ᾧr������Nԕ��料�#��y��wDٽg��=��?�Fs?y8q?��_?Wy�A6d�1^�_-��__V�#>���ΥE���D��5C�
�n���_���똾�L=:�@���C��
�?��?����-t�>/���lO���	��[Z>�7����m��ɡ� ]Q������=^�*����K��t�?��>T��>"�=?�ϊ��X��*�JG���	N�=�G�>�\�>I��>� =̓~��>���w������ ���-x>�_?<�M?^x{?�"���8��Ȁ�������Z����3F>�>�Ds>�Xs��F�t_'���@�	9l����&��0����=e�7?!Ґ>��>�}�?Z��>d��c8ƾݛ[��M.��"Ӽ�m�>�rg?���>��A>7T�k�����>�Y?s?�4?F�׾AU��������=L�?>�>���>���>�yj�\x��Uo��y�	��u=NN(?؃��Q���K�= (�?�z>\&�F?�!���J9��� �����P=^v�>��>�2�>t�(<^�tQ�z\k�P�&?�?��OU-��>$?U��>"Bk>�? �>+���p�9=T�?@g?�YM?uG8?ґ�>E�_<e�nx!=��=��>�A^>�5=�
�=q��OJ9����8��<��= �$=�R���P=�C@�{B<�[�<{�M>�~ӿ��I�#�龟���<�z
��н�Q���r�������w��[)�i5ɽf�=��\��u������@�I����?�@F 2����J0���ŋ�������?�.��Mg����w���N�)f�5���h%�\p�������5�?���<r˿<��� �X��>�\�?���?o_�^CE�>u�8u�=�.T=E��k􏾰O��	lݿ�w�=kj{?Rn�>�Cɾ5P��>3�>���>m�;>���	&%��>���><r?)?-⯽|{���z���G> ��?���??uA?Ǖ(�K���S=�?�>�	?d-A>b\2��X��Ȱ�a��>>5�?W�?�@P=�X�'���1e?	�<VFF�'�ͻF��=�=��=J��O�K>��>�����@�޽��4>=��>�!��g�F�^�h�<�\>�ֽ ���`��?�[W���_�ή)��\}�H.$>6.P?�ؾ>�}=l�A?7/7�9�Կ�b�PJ[?_��?E&�?��0?�����.�>����O?�1?;��>n^$��Z�����=�P�J���خ���e�$<�<���>2u>�&!�e ��&|��m��E�=*z�PȿsI����3=�1�mk�9L-��-��g�d�����,r�����j2�=$�=��M>��>�_>=]>ߛ`?��u?�~�>�&>�!!�ȝy��ꔾ\��<�"�����ܗ��A��`�����4�ʾ���������)績��<��= �R�Fb����!��.c�,VE���.?�m!>�%ʾf[N���<f�ɾ�'���!X�����;�2�9Kn����?��B?S���jV�|�� ��`糽�GW?�:��F�12��3�==��t�=2��>��=����3���T��f0?�V?�w��Ȕ����)>� ��#=ٕ+?w?v�b<7�>5G%?�*�j���[>53> ��>���>d#	>q��76۽@�?�~T?-�����ް�>����8z�G�a=O�>��4����d�[>���<&Ȍ��T�������<y;U?�ߏ>_
,�f�����9J�;b��=�j?J�>᧞>`?uFE?#=��徱�[����Z=i�W?�~m?~�>�hŽ/ؾ}��[:7?:k?ׄT>�{��`���1��{��h8?<sf?�&?M���lv��F��\��^]9?|yz?��W��������0�)��r�>��>d��>��.��X>��b?�6�KĞ�l&��(��7��?v@�H�?�m�,�<�ڼ�{?!�>�my�b�q��8��]���yÖ=+��>4I#��l�� �+�	�M�fP<? �?k8?��������=�[����?}��?I�����̻�/��b�����.g<�=��y�����C�����9��ҹ��s�/����F�u��>�@��ڽN|�>��x� �KyͿdꉿ��þ����?9
�>G��;r���da�*�k�-R:�:�A��p��t�>�8>FX������{�ˣ;����pC�>����-��>��T�Rm�������k<�ݒ>Υ�>I'�>�b��	������?�����[ο�=��	(�G�X?�M�?擅?l�?��,<@nv���|������F?S�s?=�Z?"���Z�nE�&MV?~@H��d��69�WfH�R�>��;?���>�B3�\G >�<��]�>#�>�{)��忿���w����?*O�?Q���+�>̡�?+� ?|������������	����=�)?2>����� �[(�A{���?p)?�v�j��]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?XU�>{Ѓ?��=�c?�o�=`幾d옼RC>���=t���}?��L?�x�>3��=��3��/�n�H�ܙP�J���[B��<�>��`?A�L?jon>k���84N�T� ��Hؽg�?������7=�ҲL��ʽ`<7>)�?>b��=�IQ�|�;�d?���y�ֿ�	����V��;?E�>��>5��@�>�{�ʼߺX?s>�>|������搿�T��?�D�?>�?�PӾ�Y���$>.@�>�$�>$�2�⽔|m��_>>0?�`���Lv��v�Z�,>�,�?E�@��?�6d��9?y�þu������e����V��b�<��%?ٯ��o��O�> r5>����������.�~�>	C�?T�?r��>X�w?�s�~�G�x�0���j>><�?��?t8>+���=�#n?��ξ�j��� ��'h?ī@e@�u�?!���6]�{���-���M���O>m��=�,>��'��=�E��͛��%s��)�=:�>�>�y>�AM>�_>� >����`%�R����F��g1A�-��.�1��ބ�����󋾠���I�[�Ҿ��Խ�WJ��ռA���e�1X[�q�>,�H??I?0�Q?a?�2�<n��=6�i>����\r=M��>��??��_?��2?k��=�����[�i,��y{��~��g��>r?�>�>'ض>�\�>�*.=��H>eE>��c>� !>�l5=�T!<��;�SJ>k}�>���>o�>�<>��>�ϴ�=#��V�h�o�w���ʽc��?׼��ؠJ��=���l��C���R��=�s.?c3>����>п�����:H?ת��� ���+�
u>/�0?�YW?!�>T��ӃT���>����j�K=>/ �@zl���)���P>O3?_'>��>��?��2#��/u�h���>�;$?��پq�轘:����\�%¶�h->��>\�&�V1�A����׌�&;���=E�L?Q�?�&��\���K����|��G>�R>�&I=ҹ>*J6>u+=�䅾�\�(�&=6�1>d>�>F?D{,>�1�=l@�>}���7P�ge�>SLB>�i+>�	@?��$?�1�(���Ճ��/��v>��>h[�>`�>^?J��@�= ��>'b>9��s9��Y��--?��X>��|��W_�`�s���v=������=*��=F\ ��=��%=�~?���(䈿��e���lD?S+?] �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾU�>�l���8���y�Ŕr���>ż?�?q���8C=��u�E?%-?�#ξq�����V@_�� ?$�?�Ȋ?�]��斿j�E��>���?��\?*�=�׾�l��g��>@d>?��+?�#?b�!��?�?<?2�?���?fM>ڇ?��~?+*?���K�c��Sc���?�=Sua���>"�>@'��FI�{j���k{��r�8����2>�s=���>}�o��ߦ�� �=�
��(Ǿ�Xy����>�re>��]>J��>��?k��><8l>�[�=��ýJ�@�F���E?	q�?=,�΂�6��=�J>�K�8�>%�<?˭���Ѿ��<>��\?�y�?��O?���>��뾛Q��������\$ս�k>/t�>@ ?��=9?#>e�)�䝾�}�>��>��=)�� =�6a߽?e�=��&?��@?Sfp��� ?x�#?��j><�>�cE�+9���E����>ع�>�:?��~?�?�ҹ�g_3�' ��ա��y[�+�M>��x?�Q?5��>���zl���2E�O�G��:�����?dcg?��{�?{(�?7�??ٛA?�If>#��X�׾C���߀>7�!?��=�A��N&�c��R?�M?{��>���<�ս�$ּ���Ev��[?q(\???&?���)a��þc�<�l#���S�v��;�3D���>
�>�n��=�>�а=@m�S96�@Jg<�{�=�}�>&�=�&7�_c����6?�P4<M1m��I�=��Z�16�y�D>�>���M�?du�ΰ��0������`r>}�?R|�?߃\?�9.���z���M?�]q?��?A�?^��J	����_}��$?����>��M�=z7�>瑾��C�>m���1���(����D��z� � ?�Z�>�5?9?��b>�q�>\�����"�Y���������k���(��}B��E&�]M�"���ZiF�@Q���������>y,��+�>��?q-M>��>44�>����p�>�o�>�$=>��>�[:>g>���=$=H���$R?ξ��(�����İ���B?}d?��>��i�;F���?M�?{-�?�vo> �h��*�1?ē ?p��.�	?7�;=���zi�<7���1��Qˇ�������>+�ֽ��8��<L��l�E
?�Z?x���D̾�Kܽ!v��Y�n=�O�?] )?��)�[�Q�]�o���W��S�/;�uh��u��z�$��p�w鏿;S������(�|�)=�*?�#�?d���v��O���$k��?���e>3�>|��>��>[I>��	�C�1�*�]�I:'�,���JC�>]{?೅>��+?�??+�>?Wme?�Z�>;�N>:���>�?�n">f��>_#
?˹O?|�U?P�7?),?x�?�*�=$�d�����'�Hf5?�:?�?���>��>%5E�'ܽN����-=������н�b	����?s��+4���'�=��>�k?C>��k�!
������s?�LG?�BA��������gة��	?�F8?��>��������|��N2?_�?��M��=��G>CP�=Ν�+ku�Q���-f�!ތ>�;�=ӓ��6 ��v=_ށ��Pm=4��=Ҵ=�n��D�Mc�>��C?a ?5�>��3�/�jLe�ff>{��>���;&�>�~���|���򓿈j���>�ĉ?�Qx?T)
�t*>��p=`�V��M����X,��!�<;�?Ρ]?�6N?d/7?�bg?k#=?�<|�ؾ;����W��8���>�)?D�>��
�ɾ,*�� �5��?{?b��	���,�Ӗľ>ɽ��>�,��)~�lԯ�EC�<;2�~���U�����?��?!H!���3�T�.��V�����B?7�>��>�P�>�%%�nOk��r���@>z;�>�GT?M�>��O?m/{?�[?�+U>�`8�g��$̙���%��!>��??���?i��?y?��>��>$�)� �cq�����u�Ă��V=��Y>?R�>�P�>#�>���=flǽ���_�>�8�=#c>���>:��>���>�v>a9�<��G?)��>R/����m����݃��>���u?���?`}+?/+=�~���E�Y���)�>aj�?���?X(*?��S�S��=��ּ�ض�R�q���>u˹>a'�>Z,�=f�G=sp> �>R��>�� ^�6f8�e�M��?�F?�=�ƿ��q�Z�p�ɗ��}d<7���Ae������[����=����Z�� ©��[�9���Æ���񚜾��{����>���=q��=V�=���<�'ɼ��<,�J=�u�<i�=�Xp�kl<c�8�&�ϻ������!\<�nI=���؀˾m�}?�<I?ݜ+?��C?�y>}>x�3�p��>緂��@?^V>��P������x;������$���ؾM{׾��c�Rʟ�{O>%AI���>Y23>�&�=?j�<n+�=��r=�ώ=� O��=�8�=�Z�=�g�=w��=q�>�X>��?�ko�����O�=����a? �S>��=U���>?�4<?է����ɿ���)�?ŭ@���?��&?Ŗ����>��I�y��=��[>c�M�=&>> %A��4A>|*/?��+�	�ǿ�}v=qQ�?Ǒ�?�QU?⡊���ݿ�n>Z�7>�s>y�R��1���\�t�b�)Z�:�!?�A;�X̾���>[�=��޾�ƾ�,=6>wJa=��f-\��!�=�z�{�;=��l=�щ>�-D>��="���;ݶ=snI=�)�=��O>����5��,���3=��=�b>+*&>8G�>�1?>�.?Ub?���>��x�LcԾB2žT��>ݮ=�>P��=x1->���>�[4?��C?4�J?m��>ۅ=i'�>[��>x�+��
q�{�߾[ۧ�j�?<t�?���?���>;��<�WJ��"���>�;����?��3?��?�f�>E��	���qO�/�(��l�<>н/]E�7#�,=H��M�н�L�=1��>�.�>�Ӣ>]�>�N>�`$>��>��O>��=9�=�v���i0<�C�=�!��.u��˔=�
��':=�9�=�<����Z��m'���-=��T=X>3�>�">{��>)
G>�竾�ا=��_���K����=�̠��9p��o�a�����ڀ~����>��=(oL�瑿��>j�>��&>�i�?!�?Ob�=�z�%(|��ಿ]&���<eڼ�<�=�.����\��U��u2�3s����>�1�>|.�>��o>Ȱ*��<�1�y=f(徳�1�S�>o���~ӼM4���p�i���}(��W�f������E??ч����=�?;'I?�ُ?�A�>�oĽͼ׾��;>�����=�/����N���?�*?���>��|�G�jǾ����=�>�+G���J��o��.1��7��a��C��>'���&4;2�4�缆�ڍ���=�Z*h�4�>�zL?C�?ue�[��:$V�m�n�}��$?W_j?�ܑ>jw??�����P���ڇ�vI�=P�r?��?��?�2�=���=%~��TN�>�7	?���?6��?�Es? 0@�ڏ�>���;� >#���A&�=5y>�͜=P.�=�[?3^
?��
?ȡ����	�C�����)^�?��<�Σ=$͒>���>��r>5i�=��f=t��=p�\>��>g��>��d>�>h�>V����X �/:(?���=��>��3?��>Q�[>
��Uu:=G�晾�����nk����8��=_	|=Tֳ�h�8���>�~ҿ_��?-�>�9�nh�>�x�7��=���<�>�E���� ?-�c>Ar>�4>>V�>Wk=�u>�+>:���K+q>�!���@�p�o�t����(�>���w
�ݿ�7�&=�П���Ӿ�h�������7����;�^�?Zj%<�\l�[8���'�(W,?u�>7 y??��Z΀���>�?@(>�Ѿ�l��|!������s�?�
@i�v>�X�>�TY?�?�&��!���k�m�^���5�7�Z�
�)�R���ċ��#��.5�(vS?r�n?�}?g�a���O>��?~��˄��T
|=w)&�X�W�RB���4�>�9پX,μ���������5�>�n?+ɂ?�Z#?'��%�� ���Eh?�C@??H�?�U�>@>H�M��2b?x��>Ym�>�J?أ.?8ge?��
?_uw>��>��zn��Iܽ"_�� ���.ݽ^��� �.�,�?=;,�=��=��S�=<G� ��7�_��L�=P�I�.А;۠�<���=�Q�>{t^?G �>�؄>b�4?��#���;�7��}W-?�=bEt����%6�������=�Tj?�Y�?Z�V?�\>��@���>��L>��>� !>��W>G�>�9ֽ�d.��ۆ=$�>��!>��=?Q�����������)�<��>��>�|>&���|�'>�xz���c>eQ��'��YR�R�G��w2���w��b�>3�K?z?9{�=Ŭ龽i���kf��5)?�g<?�M?�0�?�8�=�ܾ�9��WJ�Y����>�9�<��9���>R��N;��:�@s>�����ھ�4J>���>ƾ?���No��.��v��}!�b�>g��l_��Ձ�E�>H� >�KʾȦ&�Bё�J=���AC?�Vw>��ڽ��7�����m$>XLS>�q�>�x<>��0�jN��,p�
ri>�Ԋ>���=|�==g��Mip�2�ξ�Y�>�8D?a�a?�4�?ACs�/`x� B��S�Aٙ��ڡ�}}?��>��>~�1>qvg=����(��ѡc��s=�L�>~��>@p$�\�H�V�����ݾ�=�Yե>��?v��=��?��R?]�?,�k?�q1?P��>��K>��ཽ����&?ns�?�k�=��ܽ�<R�Ɉ7��wE���>��)?�8A�ѥ�>��?j?�7&?�P?+�?U4	>T�N2?��"�>��>2�W�iq��M�c>K?���>�W?��?�bF>��4��4��X󘽹=�=kZ>�2?�$?fw?��>���>�����2�=��>gc?�.�?)�o?�v�=i?�:2>���>+�=<��>*��>�?�UO?G�s?O�J?���>��<�7��p9��L(s�w�O�|��;�
I<f�y=��Et�-[���<�z�;�-������y�D� <�����;4�>�fu>��� />�0ƾ�����o@>����ݛ�'���6�*�=d�>�� ?���>��%�/~�=!Һ>���>s��
='?=u?]D?�k<L�b�q�ݾ]�P��8�>{�A?N��=,�j�����#�v�BRU=��l?Ǵ]?8�V�х��Pn^?HF`?��쾪*��#���
��
�x�� d?��?ub���a>�YF?� D?M�?�ԽqaW��T���j�`����ve>L5�>!WO�8������>��}?|�?C��>�d�>���%n�;==�G�??ϛ?{}�?n��?�!->ۑt��}Ͽ�I��|;��c�]?�|�>.@����"?�c���ϾiL��:D��)⾭0��'��C��9��d�$��탾�׽"ļ=�?�	s?
]q?g�_?�� �Zd��E^�l��:XV����
�3�E��E�ƐC���n�8U�����R��DH=�7N���G����?�!?�����h�>��T�Ͼ;��H�O>�ݾ���V��OY�#NM��=�K���]��ݾ((?�:�>j1�>��6?�/~�KB�#xF���?����-<>�I�>69�>���><��=��&�3݌�Z�u�Lw��0v���u>bb?=�L?�q?�G�մ2�����S�"�yP0��1����B>��=m7�>�P^�z9 �o�%�/<���q��;��$�������e=��1?.^�>��>�Ә?� ?��o0��#u��-�:
a<���>�e?ؚ�>+�~>P�㽱���!�>��^?��?A>�>6���6�'���"���GҴ>9x�>��>��=�W^�_��N��D����1��X�=�f??�Ճ�b�9��6>6�B?{�I=�w]=M[�>�j�^d�u�����&�'>�B?3">A9�=�޾��!�X킿^���v�)?�8?_����)�}�z>SA"?{��>���>�}�?���>����I;`#?�U^?өJ?�W??!��>!�=s��=q˽h�&�0�J=��>��U>c�d=%��=���;�[��!"�ғG=�^�=U8��h����T�:�z¼��S<��=�(5>h{ֿ+j\�C��j��f��-��wؽmP��/(龥���P���΅�,�d�b�x�!�=��~�z�}�\�Y������?%�@w��}	B�ԥ��1�{���/�L`�>Z����r=/��x������C���-逾��)��`I��hO������i?�y�=tMƿ�ܙ�b���ix>J�?,�?��&�V�4�g�3�e�=Z�=]�$<ԃ�	ǥ�r8ʿL+��0q?�C�> ���L:=�	&?�T>㊘>��>��|�3���t꽑�?�"?a��>`!��5m��O���v�=w�?��@�zA?#�(�����U=���>��	?��?>1X1�F���mR�>	:�?���?�TM=w�W��7
��xe?>"<l�F���ܻ��=� �=�8=�����J>�J�>�s��WA�"Lܽ$�4>��>�v"����Pv^�zS�<�]>/�ս�6��`ۄ?�i\���e�%^/��J���6>_�T?�2�>�$�=�z-?�3H���ϿS]���`?#*�?'��?d)?��y��>ݾׁM? @6?�#�>!�&�j?u��A�=���b����c>W�i��=gK�>ih>$h,��Z���P�x��x��=��<�ʿ��$���_?�<�@�˸O�4�&�h���J�'�eE���8S���8ω=��=	cO>��>�W>��T>�]?�2p?١�>ò>���.��uL��-<��~���z)�+�����HM�����]ӾQ�	�eb������̾�<�Gd�=GyL�@����3�isj���,��T"?�=���3u_�Ȁ���곾�Q��M�~�k������vF��o����?7�P?�^���Vn��\��nd�=���9�Ia?aِ�x"��k���Y>&�<�������>eg�=���צ4��H0���2?�t?��þ5��a�1>8��!��<>z;?G��>�>�i�>)P%?!����伂��>��>$"x>oD�>$�=���Ǜ��(�*?�J?j=
����F�>����$WT����+�>��E�36=&�->��h�0߈��~�|��(��=�sV?�	�>� *�K��cԑ�����K=vyw?d�?%ڜ>��j?��A?�&�<"~�M?U�Dk�+H^=�iW?nbj?l>��H�о�ܤ�M5?�e?4P>x�a�T�澧�/��� �`�?�rl?	?%�l�^�z� �����c5?aڀ?��a�����+�F�罡1�>g��>��>�M;���>��p?~sH����S��u���}�?�}@���?�r�IN�;�~�Af?=+�>3V����~�,�i�����ύƽ?����ӄ����I��j}=��`?^�?u�?;�������{��=<��{u�?�
�?�Y��4.g<@;��k�A����s�<;g�=C�!���)����8��zƾ�G
����R�ͼ�͆>BG@��齔��>6";�+�j?Ͽ�-����Ͼ��p�6C?��>�˽����?Hj�bgt�;_F���G�����-�>l�>|������F8z�TY;�iΌ�>�>�� ��X�>ϴT�H}���ȝ��$m<�p�>AQ�>�(y>Ioνõ����?,%�v_ϿfX��5���[?��?�o�?eg ?��D<�*��-�o�W�;��G?��u?H�Y?,(5�@�d��}:�5�O?:�w��Yg����b_�1��>E7F?���>=�9��*=@�=ڎ�>9��>�!���˿�%���径�?�#�?��Ѿ�:�>�8�?2G?+ �A��H\��O����=��+?C�+>�ۜ��l�C�O����3�?��-?CQL���	�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?���>P��?d��=�{�>�Y�=(6��#����$>��=�E���?�N?���>�q�=)�-��-���D���Q��9���C�ط�>�c?O�K?�$d>�����XK���NA��n4�	���u�=���(ܽ�3>�>>�/>��F��]Ѿ��?�i�Xο~i��x�X�lK>?X��>�-�>����|��c_�;��`?\,�>��d�������m����?�h�?�?��E(Ľ5��=��>�}�>v�����P�면����=�c4?�6���n|��텿AR^>���?v@���?��c�Q�?�����ꆿn���n����;��>��&?$�۾��s>%W?�+�>/�U��\���lc�d�>G��?c��?���>eHh?���+��S�>۱>�u`?]m�>8��=S�-�ȼ�=O�.?~V��贿 ����k?vX	@@)g?����������G��9Z�U��=-t=�=dPc���=�f�<t�=V<�l!>y�>�{j>,Z�>��[>�>�8>����d7)��ԛ������Z?�(�&�f���M���:�u����>ι�b�ž�ꖽ��Ѽ[����8��9��������=��F?i�U?�E]?\6?�; �=�����]�>��U�N >ژ�>�ZW?Q#h?u%=?]+�=K�|��e������ž�T����>�ʙ>��?��>lz�>	��F>>\>ֹ>^��<{�{�7�w��D>�ߚ>���>>ʝ>���=@̴>b����1ÿ�x�ig��o�Q>��?A��EC �b���d����w�T�w=sE2?���=;���_bҿ�	��>�J?�猽�JQ�T%��ZB�>CO?@�p?���>��������!!>�ʽ�OG��6�=r�,=�ˉ�d���>K�4?��j>�w>��3��6�dcP�.ά���|>�8?�R��dA���r��sG�c ޾}�O>��>�e�-��N��^R|�/�l�mN�=;?M�?�H��i%���i}�v8���N>xX>U=� �=ֻP>6uz��q�p#H���/=&�=�2^>��?u.>��=	ۢ>�N���N����>\�>>�L+>kg>?�#%?���F��#���3���r>���>��}>��	>�{L��i�=�:�>w]>B�ڼ�C���d��D��b[>h�c�if]��c��`z=4���K0�=*��=����m9��+=�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�G�>6lC��瑿kz�Vpc�3��=���>�X(?c�ܾ����eV��G?Ԯ	?�%оZ���:-ſN�]�*�?�?q�?�I`�O ��R�2� 4�>��?�>?��>y=ƾo���F�r>;�E?��Y?+/O>��� Oz�I�'?�D�?&r?'G>5&�?��z?��?��a��?��W���鍿WUf=?`�8�>.7=ǯ־�C�	��7��h�Z�*]�'>}!*=&��>B'��ٔ��E>`���u9p��&�E<�>�=Kml>�E�>|��>���>NO�>H�^�QIf����F����Q?KS�?s��H����d>���>�ƽ���>�Y?�CǼ֜��&�>Lgg?���?[�b?5,�>3'���]��#���<6¾z4���,>Q�>>M?s�.�S�����>Ͼs*�>�?IX>�J��\g?�k)@�~�2>��F??�%?�v4�S�?8u"?ڷx>e �>Ze&��g��c�2�ا|>D�>��>˂u?���> ��8���#������R&^�4��=DOm?��)?>�>1��SҞ�@��<�;�=�� >�ш?��_?~��"�>K$�?yG?EmR?~o�>�����̾�R_�J$�>U�.?�@[=�`�iF龂�s��8?�?��P?9�<�����>
�Ծ'��,� ?�;O?Ab�>�L0��4L���"�a�=�=�l=���ft=��;�悔��x����=)�>4���;���vg�%�D�&ԗ>n�>ȝ.>���Hp���::?��>D=�w�+>�le�����@>;�ϼ"��*��?Up�|�������}���~��=悯?a�?n��?W���s�@n<?���?�5?�j?K���̓��[ޭ��7�� zx�5XI��G3=MX?0�������A���>{�v��������>8��>�?�1?�=@>��>X����&�.�׾<��x-j�r�!��#I��3����󲘾 �?����Dٻ�c��s��>�b ��>��?�A>"�6>pݻ>�}>=��>UQQ>¹�>�Չ>*�=��=���=��J<l�JP?���(,���޾
����G?�f?���>X�T��L���Y�F?�;�?���?�T>��e�sQ1���?}_?1�f��#??��<��B���<�E�����4�Ҽ-����|�>������1��2P��?�?3?I�?�f�CKѾ������u<w=p1�?2�)?�(��Q�ğo���W��R�I���d�os��M)%��p�cϏ�����CÃ� �(�:S%=��)?[�?��0�����K j�N�=���b>��>{�>�c�>H|M>G	�['0��\�x�&��Ƀ����>�{?j�>? D?a�*?��(?f1g?�N>7!>& j�d#?���U�>��%?=�Y?qJ?�N?<��>7?�Y=*�|��z������@?ѱ?Q!?eD�>�ƥ>5���8>4�+�U��[9���=���=T=�E����,6�&.>���>�z<�@�*{�y	���/?ؔ?;I}>]E���D��������>֋?i�<p�r��}������A�>OY�?n���_�Q=�O$>�K=�f�=�z�u���"�<�A&>}��XV�<㬽��>��uM>F\�����:�+����5"��u�>	�?��?"�?鯅��O���n�ɶh>�SD>��>3+�=A\�UӚ�wH���'9�{��>�L�?�ʲ?턍���=��<�lU�Y�.�X� �Uٙ���Z���?@��>�]&?-/w?��>�[<? �>}?����q��Tо���>�*?��>�/�ЯľKg��tU,���?E�?�p[�p,,�O� ��þ�m۽��>��/�6�|��3��Y�@����<�)�쇛��{�?���?�0��-|4��%���ꝿ���zEG?��>�ל>= �>�/�^.o��&���I>jx�>2�M?��>�O?uN{?�\?�>T>��8����ʙ��G)���!>��??�A�?��?Ex?�b�>�>��)�5ྋT��+�����$��|!X=�Z>
G�> ��>�E�>	��=�˽���|�<��a�=��c>w��>S�>@x�>FWv>� �<��G? ��>�D��А��ܤ��Ƀ�=�=��{u?A��?S�+?��=}��E��O��I�>�d�?�?,*?�S����=85׼zⶾLr��/�>�޹>�K�>"��=xlG=R�>/��>���>P��g��a8��?M�%	?�(F?��=�ƿO�q��7q��ԗ�f�[<�d��#�d��p���[��S�=�������Y©�!�[�����蒓�	������W'|�@��>��=���=ϊ�=��<pYͼ���<��K=/��<��=:�q�H~j<�m8��wͻ���`S�I�V<��F=`A ��{˾�z}?;I?3�+?
�C?`�y>�>*B4�JŖ>׈��7@?J'V>:�O�x]��o;�{�������ؾ�׾��c�ڟ��E>��I�L�>QK3>&��= �<��=��s=���=6_��
=�+�=d<�=��=���=��>�>uÀ?&��Zݏ���7��Hͽ�[V?6��>Y�c=�c�֗^?��>�Dx�Uk¿���'�?�� @��?��(?�Q]��|o>Ac�u0�;Sf=�ﵾ~<iԕ='��
p]>��>> d������6����?���?s�H?�N��/eѿ�V>�<>dg>S�Ù0��j]��-]��XW�5#?}�9���;�3�>�?�=̪�^&ľ �D=Q�4>UJ=���.�Z��d�=z�~�m?M=�m=W��>-�A>BԵ=���L,�=��C=��=ؔM>0����8�r2�f1=#��=�gc>T $>Q�>P�?9L0?��c?��>�n�J�Ͼ2¾�m�>�o�=yg�>w��=��?>�6�>}�6?OcD?@�K?/��>�߉=�к>�y�>�k,���m��!�V��"��<�O�?eІ?�Z�>��H<��=�r��}>��0ý�9?��1?��?�R�>H�O� �������8��g���+�ս�s����5�; ����<\�?>�T�>��>�a�>=�U>{d">*��=�>�#'>�>��+7>�Ċ���h�,>��"��K��=��7�	�J=H��= ���)Y������C���=K��;��>���>���>��?ݴ->C9��ʯ}=\ᦾ�\���s>����)]�G�c�a����};��֌>E�:>�-=�����N��>׃�>�`>%��?��a?ꑀ>��ݽ�v��~k����ٽ{�齫�/=�e=Ïվ��\�n�@tP�������>�t�>sb�>0�j>@�+���=��no=ɚ�Ă4�8u�>:���>-%�G��q\p��X��L�����h�>�]���D?�Ї��]�=��}?�G?�ӏ?D�>/��S'ھ֋3>V|��R=8��	�o�a���5�?p�&?C7�>�x�#�C�k;����Rf�>��[���D�#-���@/�X�h�����G��>ֆ��E�ǾM�-��ۃ�Y珿2�>�<m���>�M?4U�?�kf�a��IW�C?�i!Ҽ�?׃^?=��>�f?Cg�>|a<"ڹ�����=m�=�8f?���?��?�F->b��=��8�>d!	?1��?n��?�ks?ۚ?�ȋ�>�
�;�� >����~P�=�>�5�=B�=ce?U�
?y�
?hG����	����	�r�]��0�<�A�=;|�>x{�>��r>U��=ʐh=wƢ=��[>�؞>��>�e>V�>�W�>>��gK��7?L�>~��>7?d�O>>�=��V��:-=$-�������_�̠n�&�2�+h�<�UM��6�<��	����>�[ȿp��?m�%>F;!���?��	���O>��P>OŽǥ�>�J>�_�>��>��>��=�H>���=�8Ӿ_�>�	��!�uC���R��Dо�"{>㱜�#�%�#	�!��lH��3�����~�i��:��ܐ=�7`�<�>�?����f�k��*��i��\�?�B�>VW6?�r���:���>���>�>�H���3�������}ᾭ�?���?���>�n�>ׂ?�]N?A�I��Д�D~�'z�D��'�DCB���������e6�T噾��a?�?��B?^�2��1>�?��m���)>'H��
.������l�>׾j��۔�湆����������H>}i{?��?�R?����{�����a?=!?���?���>�=	;b�y�?��=��>~/Q?}\?��c?��?|/b>q�=�(�!���x���Lz�������z��nL��E���_*<�a=��==]�>&iλ��A�Ľ���ͼ�|��� =H��=hC>G�>��W?F�?NN�>��&?�����O�h뢾Ȱ ?g�=����f��B�߾�>
��Ź=x�q?���?@e?�� >�4�\)<��(>+bd>�S>�?>>E��>����U��n�=�L$>�">7��=�(~�_�K�ć�t����F2�w�->g��>��>^t�":>�鯾\v%�dz%>bƘ�?!��.N��c���.��W��3��>�4'?��?̗�3c����Q��m��?��L?�3*?=sw?������,�u�R=�A�栟>�Q��������x���-��bO=6	K>�U��Q��+a>ص��徢�l�o*G�V ���h�=�
�Z?7=S��Ͼ������=}!>R踾�x�����1��J?'rn=b���^��+���0#>L/�>,i�>�4�H\��@*A�a��v��=V��>�D>cݼs@���H�o��y �>�G?/�i?���?�M��Yd��SG�����ד��M=`E?��>-?��K>D"�=�᫾���"[�BN9�1�>�3�>Y���;7��	���	�R'�w#m>Mz�>784>G:�>��J?t?.�b?j�"?Z�?0�>��l�����$?>�?,®= ���]�ˆ?��/F��>`r#?",��Ց>��?��?��&?�DJ?	w?@3>������=�qʘ>�$�>cX�u	��	�h>�O?V3�>�C[?���?�/>�3�M���Ԥ���=�>��0?Ue!?��?�Ϻ>Q2�>�ˉ��?b=���>��e?��}? �i?U��=��>��U>���>f��<e�>�]?��#?٫J?�yb?�6?�Z�>e�<���a<��/�Ž+���Ι����=�-=������!��J���r�<�1���R��B�=/�J��~��}5���>f;Y>�Pz����=��n�G$m��-r>�~�=gq��􄍾�Ԣ��{->`C�>���>���>�F����=an�>���>:�
��* ?�"?a@#?�� �x�ћ������^u�>1@?ͫ�=�9P��&����n�o� >;�}?�N?	A��s%�Y�b?=�]?�d�S=���þ��b����9�O?^�
?}�G�f�>c�~?��q?ȵ�>��e��7n�
��jAb���j��˶=�r�>X���d�n<�>Ț7?2N�>��b>��=�r۾��w�_q��$?��?u �?���?�2*>�n�G3�bC���4���]?̅�>`ϧ���"?�G�'�;l�� �����=�����+����f��R�%� ����ؽ�-�=�s?*�r?��p?��^?�@�TYc���]�Ƌ���U��f����rzE�E��=C�t�n�M�!���7꙾�vE=X J����+�?�?<?c=R��>�<���z�/2�>kEܾBJ�<�u"=ݮG��c>�>K��������4�?V�>�.?%�G?��p��a�y�`������D�$�>+�>A-�>/��>�ȴ��b��[\�&�<���5���=�h>[$`?�	L?u4s?�p�,���x���4��:4����i��=2 >΍�>	�?���������7��-m��������*��jK<��6?�x�>F��>��?� ?���'�;�[��J��Px�`��>Xg?4�>�+R>�=½L$�"�>#�^?��?˶�>Th���~��&i�-� '�>
��>i)?�9�>h�2��gU���}��`��t��z�>�Z?��p�Q�vG>NI?��=nƊ��tG>�q��6�fX��������;Ei'?1�a>e�P>�O��M վ:����V�1O�>�F'?W2�����~�?��.?�� ?�{F�P��?�K>�*��b��+7?�z?p�#?��/?5�#?�rI>G������gy�J�N=ϑ�>_M'>#o�=�Ա=��B��B���g��"��GH��$ҽ�+�f�<�����}���(>2�忔�M������
��O����Nپ��Kh�W:4�=5���ʪ�2v��*���������bZ����i�v�՘@K�@�9�ϩ��L��^�]�*�a��y�>V���O�T�n���=_Y����7�@��3$��Nb��M�������&?3v�L�ÿ�%��K۳��
?+c?��k?��=�����I�ۛ���X�� ��������ӻʿ:�Ͼ̎l?�|�>�Ⱦ�D�<�!�>��=jd#>NA}>�F��� ���

?n�G?�� ?�D���_=���F�َ�?{B @�C?�����Qξ42����?���>��?��~=�Ʒ����Y�
?��?*8�?%b����/����D˃?��>к�M�z<a�.>t�8�e@��_�=N��>A5�>0ם�{�]���(���>�	;>��4<}������\�=>��>���<�&��2��?��[�$e��</��$��?>�U?J,�>2��=B�,?�!H�9Ͽ�[�ܧ`?���?���?z�(?��Ǳ�>��ܾxeM?M�5?4�>�G'�X�t��"�=�輘�w��@�/V�U��=��>�>�,�����S�iw����=��B�ʿ5)�V�"�r�<��:#"���ұ���rp���� �������-�=j��=��>晌>l�G>{�U>�i^?gx?߰�>)O>_I��^Uh�E#��vk:�≾:A�����j�EX�őھ�4߾���1�#�D!��U��u�>�=>OAW��L����0��#[������2?C��=�'ᾝj.�g{�=�F�� ��x�>�+��V|þ3�I������p�?��j?�����l��o��>=�{��Iv?S�C�e��@�u���\>�Y|��{Q�ɵ?%�z=�����n]�(�z�9�,?�\%?M�u�-E��%ߙ>�!��y��=��O?Ԃ?������>�{d?��3=S��uƏ>���=�0�>��>>�C��D�_=/k0?X�Y?7�i�:5���[=\c���2���?h>ư���L��O�>Կ>BC�<��_=�>��ֽn�S�T?9ǝ>�(�959��g��m�=O��>iVP?�f?�s�=!pY?��S?�>���fD��p����>p�Z?�YV?�^�=ͦý� ��⮨�?��]?g>ҟ����;,���	8?�-=?̼:?]����0��*��]���/@?\�v?�R^��l���DdV��<�>��>r��>z�9�\4�>�>?��"��/��6����R4�ػ�?ғ@)��?ö9<	��o�=G$?|Q�>�]O��ƾ�,��?���[�s=�>x���rMv����@y,�n�8?Χ�?�z�>�v�����=�=�I��?]/�?���Y�������'f�������-=渶=�c�⪄����A6��0ž�(�w薾3ߙ��>��@��Ž��>�;<�n��u!ο$T��svоN~_��?��>h����6��Zg�D�n�>�`FJ�QA��&��>+ ?>��[=f�]�l}s�VV�*�����>�Oý�2�>rzw�����\��+�=�6>���>�G�>���<3���ɔ?"���ǿ���������|?�n�?7��?j+?��\��LB��e^��Ŀ=H�?ȎJ?��=?w[U�����ظ=U`?��߾��_��:�:9��G4>�"?��>�A;�[�N=��q>�D�>�L�=G:C�����Z3��$��8�?h��?mB׾��>	��?^=?�n�qM�����x�S=Ͱ.?�B0>8�u������4�}dh�E�>��?
�	=����1�_?Y�a���p���-��ƽ+ۡ>V�0��c\�K=��+��YXe����.>y���?^�?u�?c��� #�J5%?��>眕�o8Ǿ��<i|�> '�>�(N>GK_�d�u>5���:��j	>خ�?�}�?�i?ƕ��@����W>��}?(�>�
�?�-�=3��>KB�=i���D��">���=��5��;?��M?���>���=�e8�՞.��E���Q����D�C��\�>�a?H�L?��a>2����9�M�!��Jν��/���߈?���+�uq۽0�4>��=>��>�*E��)Ӿw�?��P<ؿ����
a&���3?��>�Y?���Wv�ﻥ`_?��>�>��볿���� ����?��?Y�?8׾���&>˫�>K��>!�н���#R��B�6>��B?�������o�|��>���?�@���?uLi��o
?�p��ȷ���-��:��b�8�#�>�;?���X>��>�#�=>:k�p ���p��8�>Ԛ�?<{�?|�>�Ai?U�f���H�L�<`��>��j?u*?�Ǽ0�U6>x?	������R���^?@�	@�9@�/^?�1��i�������bվ1�J�������=o���>>�<��=ݏ��C==@��>ˡe>���>5�>vi->ڵ>Ҟ����,�EX���.��T�Z�=MG���%�7�$�ê¾�d�����G�b����Ͻܬ˽= =��\I���2��}���1=0�P?$�C?�a]?��?�ʺ�,z>tR��V�=��6�}C��)�<��?��<?��>?{OJ>�m��<J��c��<:���w�h��>c�>���>*�>&��>���=�v�=ꤗ=�]c>#�=>��<�4����=�Ig>z�>(=�>2N�>���=g�~>G$��ed���%��N���D7��_�?�f�����IF��o#�}��M�G�'�|?�b6>�����t�󪰿�R?xl�V��3jO>`�K>��%?�]n?�?�2�� �>�t�>(x��l;�Uk�>��G��ͽ��V�z��=�a?��>z�r>����6=���Q��L��l�>U�&?�>��0:ν�q��3�@���7+>Fm�>��=U3�MW��zv��Ї�:m�=�b7?���>�&�Ɋ��4���r0��_�>���>n����^>�UH>��ڼ"��TQ���v���=�<N>B?�4�=
�@>��>Y`��7(����>�u�>§>e�7?�	?1B����<ٸ��oخ�Iף>ʶ�>���=�<>��)�XS>L�>���=����DL��> �ɬS�P��>��%��,ݾ�[���/ >Cl�q.>ɪ�>.�!�WǾ0���~?���䈿��:d��7mD?V+?�=�F<��"������G�� �?^�@�l�? �	���V���?�@�? ��`��=�|�>!֫>�ξ��L�6�?��Ž�Ƣ�2�	��(#�IS�?�?�/��ɋ�Bl�w7>�^%?�Ӿ���>���#��冿�s��=ú�>��I?���G�v�`�4�I�?�
?�m��m���1ȿfNs�1�>��?�?�k�񶛿�@����>)�?��Y?\�g>ؾ�c��x�>�K@?�mP?���>�\��0/��b?�2�?}��?��I>�_�?�t?k��>1R���~/��@&���=Pi�;��>�A>_z���-F�*����-�� j�z��Igb>��"=S��>�M�~Y�����=o����f����g����>�q>�J>#�>?[V�>�Ǚ>�=�֊�t���-���S+J?�+�?���n�pe�;7��=�)a�D�>y6?b��;{WԾ�Ѱ>��[?Ot}?B�Z?�̜>0�љ�4罿`��%�<��Z>���>m��>b����+>�-��0��ڒ>�a�>��h;&4Ӿ�Ym�m{��4z�>�x ?�D�>W"�=��?xv?1�>�!0>i�.����_���?���>m��>�,Y?�Y?�0���&��א�Q&����,��5>��s?��?E�8>�������b*>j. >\;>?r�?YBe?r�ʾr	9?��?� Q?��
?ˤ�>6����߭�%�p>X�>s?��Ӿ�Qz���w��=���=�>T��=�s>OH��>2Y?ئE��z��&�>O?0#0?���簚����:�>y}���g�YM>%��>�F�=�,>b[4��f>��=G�,=I}¾2�d<|��5ǅ����=p{�>󎒽���=,?��G��ك�7�=��r�xD���>�IL>G����^?l=�"�{�H���x���U�� �?}��?k�?���םh�|$=?��?k?�!�>K���~޾���)Pw�~x�Cw���>	��>��l����������)F����Ž�5�,��>��>�	?�B�>�V>=�>�Q���Ŵྂ��n`��� ���)���#�HD��1̾B�2�Z��yᦾ�ʁ�D>l>C���/�>�T�>�Do>�p�>���> ߼�,�>�N%>q�T>,!�>U֙>�q>"B�=J.\=	,��?G?�㽾���k����� �D]U?�Rq?���>6�,�'�s�k$��YdC?h �?d�?i[�>	5o��~���*?��?�lc�:��>�i�>g��=���=kj����.�>��^�Y��>-��=�(���i��k����:?
�>�=��?)���B�����SpU=�݃?��(?�)�6P�&�n�\U��S�RJ���c��Ţ���%��hp�����m���O�.)��p8=�O)?x��?5� ������2i��>� �h>Xw�>TT�>A�>�JH>+{	���1��+_�2�'�胾�}�>@�z?���=��V?S#?���>C�Y?�
�=�D�>�}����>_/ƽf��!�>):]?�>?�0?B>8?�@?W^6=#�����P���3�9>�3?�5?��?��>���������$���t$��WG���!>��>�����	�Z=S��X�?�/��>��B��=���!#?/�>3*"?:� �D��hb4>1:�=�����?]���W�񰘿,�y�U��>���?Z_�w�&>y�H>��w=�-�]��=*� <�3m="G>^Ȑ�@�:�&�x=lo�=���>U8üYx��2�=Z=)>���<x��>�*?qW??pb�>�����6��5�>A�!?4��>��;>�ǿ�c���6���OS��.�>o�{?��?�N/��=#>"	=Hg����׾�u���7��@�=I�?�S�>"O�>��?��?��#?�FO>��v�����}�����<�?ݑ*?��c>��i}¾{D���.-��.?��?��^���o���W����̽�q�=,n4�lT�,+��x�;���C=MN��c��٭�?�f�?ڼ��;<�Q.�Ĳ������??P�>Vū>2u�>_.�6�a��!�3�>��>U?��>}V_?�p�?Ec�?g~�����z���5���? ���%?��	?<L:?��u?'�?T�7>��=m٨=�v��{���٭���r��zLJ���=A�>>�w�>�W>��}���r�,(��ܽ(>[��1�>��P>bw�>n�T>��|<_�1�S�H?���>�i���a�Ia���v�:̙<�*r??%�?�===��3�r���X��>�_�?���?��/?�6Y�IQ�=�	������`�j��`�>X�>�$�>�	=H��=�Z>]��>�7�>\����`�/�ya;ѹ
?FD?��=BQ����w��쑾�i���yj<�3���Gj�����l�ɞ�=�"��4,������q~��߰����w�վ����U�A��t�>P�2=Ԟ:^�=��<���<���=�r�=�#H=~�<	*���p��`<�1�;�)/=�R��<E���=8���I�˾Sz}?+�H?�_+?-D?�9y>��>R�8��Ė>�̃��?n�T>�L�k����z:�������Mؾ��׾�4d��ϟ�7�>�cF��h>p2>pj�=Q�<���=Op=◌=��3���=���=�@�=�Ĭ=���=��>H$>�6w?W���
����4Q��Z罤�:?�8�>g{�=��ƾr@?��>>�2������xb��-?���?�T�?9�?@ti��d�>L��}㎽�q�=Q����=2>���=z�2�U��>��J>���K��J����4�?��@��??�ዿ΢Ͽ*a/>� F>��= WV�h�'�m�R�U�R�Јc��?s�>�[l��~)�>q-m=���zǾW�<*I3>���<v�:���S�wS�=�ڌ��f�<��9=~&�>�{H>:��=�՝�	<�=��=��=>�?>H�<�I���>�u��<e��=�k>�>�A�>�?\b?�i? �@>�'��6���;���>>:�>L�P>�;>m�=��m>>$?z�9?��G?�%�>T��<�j�>t`�>7⾠�c���"��rᾒ����?�S�?���>W�!>�$F���h�o��묾�E�>�y*? �-?M�>�#��u��B�	���b�.�h������}$�(9D�$�<��������M���=g��>g��>h�>w��>���=I�=��>���=δ�<x�/=���=��Y>}��=��<������3��b#��<���=� :�[��<'
>">�Y+��x�|]�=0��>�8>&I�>m6�=ݤ�	L>&Hھr�3��>>��+D�!2U���l� ���,ҽ�>�%>8��-��3�>��>_54>���?R�u?��>x��Ua� ���������¾cj���=���/�7�a� <?���S��>Yk>�Ó>`#f>�<&�x�5�߫�<�C��k�8���>*v���^�?���h�"������+�m��~�A9M?\��� �9="n?�_H?��?A��>�R��� ۾R4N>�n7��n�=����F��:��^"? 1?&��>3޾�EC��ľ�;�����>��4��P�w����0�2w�7q��Jƹ>�(���	ƾ�x5�����e�����=��m���>�EM?��?:�h�0Q}��L��!�6��T8?Ыg?kO�>-�?3�	?�İ�r�ҏ�劬=jtl?���?�&�?���=57P�g�~=�n>!�?7e�?�#�?�4H?>���WV?�b�K��04��O>��>j�=�H>�i?� ?��>�K��WG�z%��8��%#���(A$>�?u>UИ>��>��4>n�>�Z�>B~>���>��>��k>��q>Rl>!E��[%��)?�>?a�>�(2?��>ֆ��ϳ�����5��[��Zb�!Cý�d<�j�=�N���<F,��.�>E�ԗ?�Yg>����D
?0
��̜��S>J|w>ȡ����?�=M>��h>��>��>rUf>l�>�sX>nDm�u����+����X��ti-�*o޾1TU>i� �g����ϕ�ՖȾyɾKX��'f�B�J���u��g��
=�Gq?�̽ư@�I��>����>H�>�jY?�&��􂯾�<
�=1�>�ݦ>Cc&�-s��������6�B�?�s�?74c>��>��W?��?ߊ1��3��oZ���u��#A��e�=�`�O፿-�����
�Q俽��_?��x?�tA?�ʑ<�4z>���?��%�[ҏ�p%�>�/��#;��w<=1(�>�)����`�k�Ӿ��þ<�^HF>��o?q#�?�W?QV���`�^[�>�P
?�?���?"�#?��.?3ʾ�D?s�=���>�^�>+�.?��:?�(?�f�>�*�>NG<V`�d���@�g�	p���<G7���=N�>mV����A=*M��8�<��c�f<�$>6�<�r1>���<O�=�&�=j�=�=a?���>#AB>ٗg?�i=�QھGH��@?>�<��O�����h��ؼ�*?>��K?"��?[�D?��ӽ#_B�������=F�g>� �=�b�>��T>rN<��M���I>��)>�ޣ=B�S��(��(�Y�Ѿ[č���@=��>��>c%�>��g�>���u x�bSo>�����>�����ngW���#��wN���>�T?(?�>=�]�5�d�c��'#?Α.?`�>?�`s?!�=)UϾY>��48�a�.�p^>�D��W��s���'����-��@�=�g>�e���W��9(�<X�<���Ծ$\G����uc��2>������ۢ�� ��퇾>4>�4�>_ ��u�$�G�������9AI?���p�Z���m�0�h��6%;�p>2��>}e�d
C��S��Vɾ��=3��>l��<�������:�m��?��;#�>�QE?��_?�o�?h��2r��B������m��lsü��?��>�?��A>]	�=�e��� ��d�F
G�!#�>`��>l���G�����%��s�#��e�>��?��>��?/R? �
?��`?��*?{?���>cյ��z��p:&?�?�ʄ=��ӽ@�T���8�@F����>�|)?��B�X��>�p?��?��&?�fQ?͕?ȏ>�� ��$@�aa�>}@�>�W�'Y����_>P�J?��>��X?l��?��>>�b5�����u���9�=+z>7�2?�#?3h?Xȸ>�F�>7X/���=y�>��?c�?U>f?�x�;��%?�}�>�g?Vc���h>I�>��?��d?�-v?��3?���>d��;�`�w�5��+1�;�"�=���=��=�5�������]���Z�b��<�NZ�8E����@��Ӳ�=�퓼���>ˊW>����K9>��̾Tgd��(2>�/=�Ő�T���6�M�u=gTm>>b�>.�>�)K�I�s���>�*�>�_��0?�X?��
?=�|={�R����w@���#�>�^J? >��l�憋���s���b=a�r?c�S?�������e�b?e�]?�r�;
=�~�þu�b��~���O?�
?��G���>��~?��q?���>��e��@n����0b��j�W��=�u�>�S���d��4�>R�7?0F�>,�b>��=zV۾(�w��i���?��?���?D��?0**>2�n��*��j���"�e?��?i��?�>=�������Har������;��=��������´��2�Z_�nýlH�=��?ód?~�a?C�o?�۾l�Y���U���v�)U�E������/�N�cWO� Q�㋂��)(�B`ԾKT���j�=��V�"8�z�?���>v/g<��>���=]���I'�e�>�n��y�p��8��e>,�Y>�2J><ǽ�q�l���ã)?=ʱ>1�"?1G?%���2�>f<�2]t�A�ξ ��>��?��%?�[>��_�� =]RU��/�>l����0=x�o>�|Y?��X?Xt?Z&(��y9��Hn�$�/��RV��sb���=+T>�X�>
?�m�'�����:'��^d���� ��5X�,tf=��!?#�>�S�>[��?���>#h�"�־ �����:��D�=;��>o�U?et?ae�>%D��#����>k.y?��>�]�>�o���V�2⏿��=���>Ƙ�>�L�>Z��>��f��J��������k课�X�>�G?�r��yjJ�<hQ>�X?��$(/�.Ǩ>�?��,�t�nʥ�c���+��>��>Q>MT�bE��"�v������1?q
?�`����0�M �>�(?��>���>�F�?iҧ>o���rn�H?c~V?��J?``E?���>$��<�t����˽9�&���d<��{>�.N>��w=�=L���[K�IA����&=!#�=�z�����4�<ڽ��ب<J�==�6>�����:��(q�DY#�E��K�!�2���;L���$�o-Z���۾p����0��fH���=n.��I�Y��ڀ�Y���p@�$@4���O0�y��U؅�cZ:�*�><���Z�9��Q���9k<�[(�#��о�d���3��L��Ҧ��H�?����������ھU��>$��>�p?�~�[!4�# ��6�=��5��k�<��Ğ�g�Ϳ�d��IJ?T;�>�H��L���~�> >�)�=w�>h���|�:����>�A3?+��>���P:����Ϳh������?�@_gA?t(��B쾅kY=���>�?*V=>��.�Ud�������>��?�݊?�E=�W����|�d?�4<F��o����=d�=�=Ԕ�8�K>zK�>�+��A�9ٽ	 2>��>�$����^����<� ]>F׽�U��1Մ?�z\�@f���/��T��QV>��T?6+�>6�=��,?:7H�}Ͽ*�\�+a?�0�?���?��(?�ۿ��ؚ>��ܾ<�M?�D6?���>�d&�:�t�4��=�:�_����㾐&V����=��>��>��,�����O�H����=�	��ؿ�t�g�)��)��kц<��ټ���H���V���(���T�2'��;��=�A>��p>\՞>��y>yq<>��c?er?���>;v>_���b��
QҾ<��������r;�����񭽕嵾F�ΆV�����������ؾ��d���=�c��I��Z�(��3[��a�I��>�>�}�t�N� q�>�Y�=�����W/>�L�=�	e��Ϫ��ó?�`_?�o:��YϾ�1)>����R?�@���>�%���>���Ԯ齼�C>��3=Ո��w˾T�V��M(?�?U�ھ��H�<���k���A<��1?�l?��:O�>l ?��I�k�P��aK>i������=� ?<�N>Y���a��ſ�>;�A?|���}�Z�b>��ξ�Ia��ߑ=��;$G��S�<�E�=DF�X��.<��ɽ�'n�U?���>WU'��N�⓾�)Q�#��<g�w?�L?���>�h?aEB?��=\����R����X/=T[?
�g?]>��n��ξ�B��)�4?�%c?�H>ām�:Y��$�i��m	?�l?�?�����|u����50�L�-?��v?s^�ws�����H�V�a=�>�[�>���>��9��k�>�>?�#��G�� ���{Y4�$Þ?��@���?��;<��U��=�;?j\�>��O��>ƾ�z������8�q=�"�>���~ev����R,�e�8?ܠ�?���>������ˆ�=�����`�?!8�?l���U6[<����Kl�g�����<��=v��R`&��	���7���ƾ��
��m��?����>�=@N���>�!8�6#��=Ͽ���о�p��?X(�>�ɽ�ࣾ�k�R�u�z_G�[�H�:*��T��>|7>�_>�����y�.�8���(��>$Z�;q�C>4/0��ˈ�J�����l�
Ǐ>��>~;�>1̡������?>!	���Ŀ<Ϗ�F���Ye?���?���?)�?���;���.V��4.���<P?�|?��8?�-�jsĽ�5<��j?_���g`��p4��kE��T>53? ��>�"-�DUv=�>���>n�>��.��VĿ`�:���ݦ?py�?N�}��>m@�?�}+?-a�O�����*����(�@?ע0>4b���,!�r=�����ѯ
?P0?��� C�I�_?�a�.�p���-���ƽ�ۡ>g�0�f\�\R��ߣ��Xe�	��&Ay����?A^�?b�?���� #�O6%?*�>K����8Ǿ^�<`��>�(�>�)N>�J_�^�u>|���:�}i	>���?�~�?Zj?򕏿����U> �}?�>5�?Wj�=<��>Ny�=�'��H�P���+>nQ>o�c�\�?R�L?0��>��=�4���/�\�F�bL��m��B�ݒ�>�k^?�aJ?��_>V���=D��!��Qƽ�<(�m&���?�:��)�o�2>&�>>��>�E�B�Ӿ��?�i���ؿ{c����'��-4?���>�?���|�t�y%��7_?\��>3��)��n'��m�훫?QB�?�?��׾S�˼G>���>4W�>$ս�ӟ�O���/�7>��B?b3��D��4�o���>g��?˲@�ή?:�h��	?���P��Ua~����7�]��=��7?�0�!�z>���>��=�nv�޻��Y�s����>�B�?�{�?��>!�l?��o�P�B��1=9M�>Μk?�s?Ro���j�B>��?"������L��f?�
@u@a�^?*����nÿȉ��)���K!=7��=7�*>�� �|�.>�\�<C����"��92`>4!�>ؚZ>;C�>9+�>95|>��>SP{�@��V��<��% J�����/A������z��}������UƵ�O`�$`6�@���k1���ǽA�����=_�T?liZ?�Zp?�?�/�
d�=_3����=ф���9<m>�v#?��??�n?K�>�~���c�t;���V��.�a��Y�>�>	&�>� �>�^�>;@��=}2>�F>���=�
(=��=L��=�cS>�,�>j�>�J�>8P>HT=���w��Y�T�J���T���?XE���tO�2�La��>����U�=o
$?p��=�ׇ���ƿ��V�I?x��O�վ��
b�=�?CG?�*>�Ģ��$���0>B%�[t���2>���F ��w5<��x>�>7?z{�>�($>�?!��2���;�q1���j>��2?.����	���b�b�:�&A���ì>���>�O�;����8��O�`�n�V��0l<"<`?�h�>$�\��^��܏��E+�=c�>z��=��b=�~2>>�z�����������=%v>��?X4G>c��=@�> �����sZ>��%>��K>t('?R�?��˻�̼�Pt�.O0�\8K>�Ρ>-�p>��>��W���D=}�>�7>K�i<Ȥ�<D�+���r���8>7�<��P��lҽo^=v���Ɵ�=�>�Q���6��=�;�~?���*䈿���e���lD?Q+?� �=�F<��"�@ ��fH��?�?g�@�l�?��	��V�E�?�@�?�
��,��=�|�>?׫>�ξH�L��?��ŽǢ�ٔ	��)#�TS�?��?��/�`ʋ�(l��6>�^%?$�Ӿ�<�>���Gx�����
�v�D�=)��>9H?0�쾬o��ZB�]r?��?���m����gɿ� w��
�>���?ꊓ?tk� ���9���>h�?U/X?e�j>F׾�Rf���>H�<?��T?��>f*���$���?A�?��?k�L>b�?A�s?C��>��a��0�^v���I��3 �=�0<֐>�W>�潾-H�~���$���h����`d>u�=q��>@�佱������=�<������遽D.�>�#r>� B>�_�>� ?<�>
�>��=���&�����a�K?1��?����0n�!9�<���=K�^��&?lH4?�b[���Ͼ�Ԩ>"�\?���?�[?�b�>���|=��	翿]}�����<)�K>�0�>BH�>���UFK>-�Ծ�<D�@s�>�ϗ>�	��:@ھ�+������B�>2e!?��>�֮=��%?�#?�'�>�{?�U,�Ր���b����>���>�r1?#]�?!�?|0�h�P�����Ƽ�����E��>�m�?�Z'?ti�>�����P��b �>�|��uL�oy�?IE�?��㽫_?���?��J?�?=H>%�8�����u!�>� >F�?��U9��$��=Ӽ$?�)�>��?�|���;��-u��"��#��C&2?|�O?���>�ո���P�I�f�@�X<�C�<Wo�=�%���ڽ���=2��>O(ݽ��� C>��p>��>��M��>�'>IRO>��>�Ӂ<��z��=�<,?b�G�A؃����=��r�yD���>�DL>�����^?�m=�=�{�k���x��YU�3 �?���? k�?����h�t#=?��?�	?� �>ZJ���{޾t��YNw�V~x��w���>��>��l�V徒������MF��K�ŽT]�g��>xE�>]�?�2?[�z>��>�m��۽&��jҾ*1�=_��D��{�A����mm�5�����۾�x��e��><�1����>�1?yܛ>�\>�>�>�𚽦X�>�{�=j��=;��>�[�>�F�>��P>�_½��	�bY6?�[��
pB�"��H��|�?>??*)?{:=���#�����?��g?{oz?��>�!���HX�ܣ?��?gB�ȗ�>�?>�r���>E��do�O����(�s*�>��=�3#�
�D�����N?j�5?_H��5���б�����A�=���?X�[?b�!�h{Z���C�_�k��]���t=�現J����>0�w+|�� ���q����[�˸�\��=��*?���?��
�Nl���]����c��B�� �>E��>v�>y_�>v�=J��}5��p�Ni7�� ��\�>x�z?�ZM>��O?��Y?̯1?w/?��%>��>���Z��>^�O=�@r���>v�!?d:?��)?�k5?�?F�=�Lq��6�X���:�>}(L>-?4�#?a�=?¹��S����@-�W���R��\9��Ѵ=��U>=C���b�o!�=AG>�K?WCݽw&�>�t*�����>�VD>"KK?I���R��\>�p >`N'?��1>\Ua���e���C����>�R_?QJp�C��=��=Y��=��;��<hb)<*I*>4R�=���C-��4>� ><>0(S�c���C�;>�B>R�_���>%~??��>�~�>�$�����x����=I�0>��i>���=٘վ�������x�n���a>�C�?Iu�?��=t�>7=�= ����N��e<������BJ<э?��?MiT?���?�N1?Y2?��=7�t���R�|�kh��Xa?Z� ?�#�>��o�$>��������?��>�q��.>y�ƾ��<�zǾ+#W>���Q�A�0袿W�8�5o�=���U�ʽ�	�?Q��?4B˾��v�� �a����Ga?:��>�?Z��>��/�\�f�3-(����=�T'?J�`?	��>��K?b��?Q�a?�,>>�<�%���콛���;��P>w7?�e�?)/�?��r?��>+H$>�c��g۾G��ӗ�Y����|��Z=.d>P^�>�P�>�ͧ>�=�K�8���]�.��=�>f>�y�>�M�>�>��b>�\;�G?%��>]*���������Ń��=��u?#��?��+?/d=yp���E�K����>�b�?���?b3*?ƅS����=+�ռ�ⶾ��q�/�>DԹ>6#�>ah�=,G=��>x��>U��>���e�	]8��.M���?�F?f��=��¿�q�>怾1閾�9_<[苾"/s�y.��Y�MW�=����&�}�����U��`���F������|��冾���>��L=��>�û=��<2���<�jC=w��<�;=�B��tl�;�����񒝽�*���H�;�9=������SI{?��D?~G(?M�??l��>{+>$8����>2L^�� ?�YD>�75�	���3�����9)��
վ��ξh�b�������>gm����>߃:>-x�=���<l��=Jq=� �=����B"=k��=P/�=J$�=5=�=�>��>�6w?V�������4Q��Z罦�:?�8�>q{�=��ƾi@?��>>�2������xb��-?���?�T�??�?ati��d�>X��o㎽�q�=,����=2>^��=k�2�F��>��J>���K��S����4�?��@��??�ዿ̢Ͽ@a/>�c>_��=Qha�*�%�flg�E	����T+?�*�z{⾢�>��W=�Yؾbи�<��=A->(�&;�z��T�e���={ ����=E��=N�>�Y>q�=�If�Y����f=I�>�>�='1�&�R=���<�}O�����\->�=J>1$�>�?�0?�nd?� �>Rn�z�ξ���� �>2��=�I�>���=s~A>�"�>�h7?��D?�L?��>��=���>�'�>�,���m��!徳ꧾr�<�q�?�j�?΁�>k�S<�tA��)���=���½TI?1?<7?��>����6� ��8���׽��<*��=©���#��>�8��ɮٽR�'>8�>"��>���>D=�>��a>K+9>���>�e>��<V�f=�&�`��;�͐��A�<Fýw���\��L�}=<!�O�?;1@�<e2=�o�<��<���L(�=]�>�d>��>�
P>�5���%,>(Ǿ��p��pr>e��
<�#���4�(�:�����lM)>�=*�����Z�>�m�=�{=>�?�?�o}?�Ȼ>�K�=�j������ؾ�K�������[>��s��V���D�j�-��g˾�p�>D��>���>���>��-�:�_����<����`�hP?�w���ER>�'� pP��wވ�i�;�0�<mM7?uŇ�,��X_?�&4?�o?"�>R\�=�fվe�>�F���	��\$��*�<�=� �>�F?D<�>� �@[@�u�����0�>R�> Y�=rI��:��}���M�52׾���>����wݾ<��匿t�����A�1(��p�>�V?ym�?�������$_�C���y�����>��?d��>0�>-=!?*"����ؾ|�t�i�=T�k?w&�?��?Q�;>xP�)�,>Q�	?z,�
��?I(�?�Q|?P�3�?T�5>^	�>5���yf�&����>	�'?��?!h�=m�=>v>5����`���D�&z�8}��H;`E�>,��>�bn>7�>�>�o>k�>շ>�6�>=(?mv�={�r>��������>q��=��g>��2?.�2>9"�=�4��A�E�'�<�pT���D���ӽ1nE���<�49�<��=�����>oĿ⮗?RO>+�׾b�?����Bj��F#>�Ni>�a:��y�>�T+>��>�	�>{�>��=��r>f�.>�Zþ�T�=7��D"�=�=��3L��Dܾ�
�>�ˑ�kvL�F�����(�N�= ��h �_�i�����}�B��<B����?KX뽩�V��"����	 �>M��>6�1?�À��+��9	>���>�~>�������.���2�m �?A��?�ib>��>Q^X?Do?�1�*�5���X��Rv��9A�|�c���`�K|��C������ʽ�^?y�x?��@?Vg�<&Pz>eH�?�%�d���f5�>��.�3�:���@=~�>񨯾��^���Ծ�ľ"��6(@>7^m?��?��?S��so�D�1>8�8?�(?v?�4?Y�:?f����$?5�>>7�?�}?(`1?5�*?��
?y>>�V�=ʹ4:j(=�施KЊ�b�ʽ�߽����`=�C�=��i;nϭ:���<���<���������~���}�<�TE=-�=���=�>�]?c�?8->x�Q?cq��AA����kP?�>l����g_{���(����[E?�?8�h?R>u�U��XQ��i�=�<>��I>�R>w6�>dDW��o?����<�<8_�=�̼^��m��
g��$􈾹DR=�`S��f�>��[>�u$>E�p>���������>N-��\�%���=�+�;-�]Gl�S}�>y?�s?��=t��Pux�V�a�}��>uM?�>f?�K�?Iꊽש��fgi�g��B����g>u�W�����0%������X���T�=�NY>�ɷ�Vt�� �`>j�B��e�l�zI�yJ��wv=�e�}|�<��
���Ѿ�Y���{�=[�>U溾����L�����U�I?aI&=Y�_�P��J��� >���>l.�>��w��_����<��c���=��>��0>�ɋ��'�IAF��1�<,�>�cE?7._?vj�?Yu��Ыr�iC�����T^���Ѽ�h?bJ�>7|?ަA>
5�=
���a_�e�d���F��\�>���>f���G����\󾵳$��x�>�Z?3p >��?ۆR?'�
?*)`?� *?�?u̒>2 ������4&?��?n��=��ӽ�(U��8�(F����>��)?YdC�i2�>�a?��?��&?eQ?��?%&>#� �^8@����>C+�>(�W�I��x._>:�J?,��>�Y?���?p{=>�I5��ᢾ'���:��=�|>��2?/#?_�?%��>"R}>]�Z�O�'=���=��?;]�?�lg?�j����!?&�>�5?�&h�*#�>&?H�(?6�\?,�?�G?���>�&�;�e/��Ž7e��O��=�_>Z�G���=�ރ<���!kٽ�4�<2�} u�؂ռ흓=�h�ս߬����>��n>�t���A>yл��b���%@>����\�����P�G�h,�=�>UL�>���>�1%��N`=a�>3��>� �<�!?�O?I?�HL<q�Z��ݾ��{����>))D?a�=�D_��͏�S?m��ȭ=�s?�ke?�u�������b?� ^?�_�.=�4�þ��b�\��f�O?��
?;�G���>��~?��q?9��>�	f�V?n�)��1b���j�B��=���>FP���d�8�>��7?�G�>)�b>���=2�۾{�w��|��@?��?#��?��?J*>��n�62࿎,򾶊��&Z?��>A����r ?�/�V�ɾ�������@�m���,<������8a��6�*�'����н�ɻ=��?K�q?�=r?�]?>����b���X�� |��>V�|�%j�{�D���C�;pD��Gq��������X��b�_=��a���9��;�?gs?;7��R�>�� ��r��ߔ�0S>����*��F������ר=0��<\�����W�Ȑ�n{,?eo�>P?��6?���2�J���^�OFJ�����j��>���>��	?��>7�����Sc���վ /���=��u>A�c?9(K?@�n?r`��b0�>i��V:!�<;�>I��<�?>�A>��>��V�/`��K%��$=�c�q�RM��v���g
���=Xq1?�>�ٝ>!7�?�?�X�������z���0�W�<�V�>v�g?[q�>o��>�۽��!����>�;e?,��>K�>��g}$�*B|�u����>W*�>5O?@[�>�ˬ�;�X�ۯ���]���6'�҅y>�l?lљ��:���Q�>��f?����Ђ���"�>�뽀E(��
���?�Pړ=� ?�tJ>�%>/埾���۸c�2���u�!?n�	?'%��ل%�~�>ٖ$?I!�>�t�>�ӄ?^�>�4ľ�v���!?S�]?�E?�??o��>� =i����)����.�Ю=%q�>�Q>H<�=��=���a���%�|�=��=Hݼ��Tٽ�du������6�8�=�5>��C�a���뾬T��P�#������m�[�l��c��6���I%�����,������\9�Z#�����9����?�@O��|<��Ѫ��ӗ��-��M�>{C�F0��_پ3��o�/�ɾ��~���>� E|���z���'?�w��(jǿq<��l�ܾ3�?�y?�py?��7�"�L^8���> U�<����v� c����ο�5��U<^?��>�Vﾳ-��dm�>�݁>�W>�{s>u�� �����<�'?�,?���>��s�O�ɿ�^��ok�<Y�?ܴ@v�A?
�%��꾯fJ=�U�>��?@;>��#�������A��>`c�?Gڋ?,7$=pwX��E/�H�d?��<�ZB���@�)d�=�+�=�N$=@+�&�E>�a�>	[!�"�>���ܽ�36>���>O:2�����T�xa�<�n\>o�ѽ�4Մ?+{\��f���/��T��U>��T? +�>@:�=��,?X7H�a}Ͽ�\��*a?�0�?���?$�(?;ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=�6�'���y���&V�v��=X��>e�>,������O�J��Z��=�*��п�" �*��))~=�sg=0��f$����`��X����<���>��ϡ=�=�=^�>t_�>�\B>rM=>�Ge?��k?ԯ�>n>?>�4�����)پ�qa��?k���"�B���b��#=ھK1Ӿ�h۾����v�B����Ѿ��K���a>��~��ڝ�j��bT���o�̠?�̷>' �"�=��L>;��E��7>Ro�=�}�Q�8T�� �?�<Q?򤋿��L�9��Yü����ʌs?>XO��V���^����=\��/�A�B�?}%�=k����*�|3i�wW>?��?7����q����p>7���Լ^Q?7�?O�>�/�>�U?Y� >S��*N<U��Y�>��?J��>p�ž�:����>��U?�0���Ǿ_�;ݯƾ�➾�H��V��>������N�_�>�8w>�ʮ�A~�����=bӍ���k?L�>�?��i����*��T���&>W��?�d�>mަ>i?G<?��>dV�jQ��(4��|7>Qj?�Y�?nĀ=�Zu=&W;����N?��]?>��=]�
�ز��7��\���4?�=�?4O�>.XP�0=�!Wh�����/?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?z�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������K�=�䕾Je�?��?nժ�ׁg<z���#l��?�����<+��=���*�#�;S�0�7��%Ǿ��
�Nq��M>��Ǐ�>oJ@�~K�>D8��"�s>Ͽ��о2lq�]�?.}�>iǽT����j�BFu���G�k�H�䀌�w��>\'>�旽���=�w�Z�9���(��E�>���[$�>@1\��R��vA����<Ë�>6�>Q[�>|k���Q��$֗?R����,οk���7^�@�Z?>4�?UN�?��?���8�p�����/��|G?/�r?"�W?���38Y���9��l?K���P�S.��;���%>2?���>ʎ"�CC�=!�=RS�> iH>�x/�)@���#��~ �2��?^��?�羷��>ʼ�?v�+?���3`���ϟ���0���,���D?8�C>M��@�$��� �J�S��R?�:0?�k��T�_?"�a�H�p���-�T�ƽ�ۡ>��0��e\�O��#���Xe����@y����?H^�?d�?��� #�]6%?�>X����8ǾL�<���>�(�>*N>�H_�{�u>����:��h	>���?�~�?Jj?���������U>�}?Pj�>�&�?Ћ>�W?�R>h������x>���l_ֽ�?sAF?��??v>�@_��-���
c���U��6�a�"E@>Y�R?�Z?�5�>=�=�J=<]\�˪S��{�������z������ͽȿH>G�>��=N
�$��? p��ؿ�i���o'�y54?(��>C�?���ܳt�d���;_?{�>)7�,���%��B�Y��?�G�?�?y�׾�S̼ >(�>�I�>� սJ�������7>4�B?���D���o���>���?��@�ծ?�i��	?���P��Va~����7�c��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?yQo���i�B>��?"������L��f?�
@u@a�^?*~ֿ��	[��出�U��=�њ=2>5�ٽ�f�=y�7=��2�=������=��>�d>��q>|�O>eR;>S)>0���
�!�$\��B���k�C�&�*~���Z����{v�xU��B����������=ý����-�O��!&�M�a�g�=_�U?�'Q?�p?���>s�p��^>6���� =�*&��v=خ�>u@2?�PK?Qo)?o��=e#���c�[��>ŧ��-�����>qE>/�>p �>Eү>}�t���K>��A>X�>��=�34=qq�B_=j�S>�1�>J�>�r�>.��=S�=����ʫ����A��o���g�����?�I������V��uF��d���#�	Y?�'�>��U��Hп�<���P?B�����8��W~
>��>�J?I�`>��'��X!�k��>^���
�K��e'���]���<�D���D�>��>�s>�F5�� ���$�Zu��c�o�9?ǋ�Ĺվ�Jq�S:��_�{��>F�?Կ�=8���q��͚r�D�[����=�`?h@#?�۾'�!�c�u�Vy��G9�>���=�x��1�=��$>�>��!�Q�Ԯ��.Ǉ��5<>1y�>¯?�L*>n,�=^J�>�C��^�P��ͤ>�EB>�m(>
�=?�6#?I���̅�l2��id2�]�n>C��>�/�>	>�fM��5�=Ԛ�>]�a>͗��'��B����E�BTU>�*n�Ql`�L�j��Jv=)��h��=�V�=w�#W=�N
=�~?���$䈿��'f���lD?1+?� �=�F<��"�1 ���H��;�?f�@�l�?��	��V�)�?�@�?�
����=}�>�֫>�ξ(�L�ܱ?��ŽgǢ���	��(#�TS�?��?��/�Iʋ�+l�U6>�^%?̰Ӿ�i�>_s��Y��f����u���#=���>9H?�M����O��	>�xs
?7?�Z򾻨��0�ȿ�|v�*��>��?���?K�m��?���@��~�>ġ�?�fY?�qi>�j۾ZZ�\��>��@?�R?��>�7�Đ'��??޶?��?�5I>kt�?��s?ݤ�>>{�e=/�<#��י����=�%�;�&�>ߚ>R���|F�ۓ�/i����j�[���Nb>j $=5��>^�x滾!ܵ=pr�����=�f�a��>��p>�QI>�<�>�� ?[�>
�>�{=P������I�����K?���?d���m��0�<��=21`��<?�P4?q�t���о�(�>W5\?۵�?��Z?+#�>c��+��k����v���[�<�J>$�>�d�>���J>��Ծ&�A�{��>��>�1��.Yپ�����L�� ��>�� ?��>���=F-?�>?���>t{�>�)E�����h�&�Z��>�?�>�l#?���?�@�>����e>I��`��AH��<�3�P�>�p�?��0?�ٌ>�_��/k��3(>/!½DU���ۓ?&@?EC��Sc?�0�? sH?w�?��i>Zk��l����ć��>PN?��!��A�a�Z3�/;�>���>���>��g� �N��c���&��P��'�?�dJ?�?���^R��j̾۽=��^�#Z=[�n��Ys�=t�.>j5��{�Ƽ��>a%�=�P}�Eo�_�=q�|<jG7>R=�=8����:0=,?��G�tۃ���=��r�>xD���>�IL>����^?[l=��{�����x��"	U�� �?���?Zk�?A��?�h��$=?�?U	?i"�>�J���}޾5�྽Pw�~x��w�W�>���>�l���I���ؙ���F��f�ŽO��K�>���>�$?~��>)��>�W�>Ό��i������m�-��^��v�	^���.�mH���=þ�w��x^��!Ѿ)Z�C*!=�;�v>U�?4S�>�AR>`��>�Y,���F>�hh��.I>��>*{1=�K�=s'�>+�V�����<,O? oϾ�(�����k�_<?
??ɞ�>쵡<4R���j���>��?�a�?�tN>��Q���F���>�0�>��P�R&�>a0�=�#׽�;>�־mC���eĽ��	�!p�>;xQ<t ��d8�S<�[?*?�Q���l�I����->o��?�?^�"?7U���(���L�6/k�)0�5�>6�z�x3�<�E�@�{��d�>��ꂿ6���o��>�1?5�X?�����d����O@��3T����=�u?	z�>�/�>r(�>dS��Q:u�C/����/��L�2(4?�z�?G�>Bg?ӐC?�B9?03<?�n�>�e�>�o�>V�>H��<�+[>�G�>��H?��?�?O�;?�kT?���>Y�9�<ҫ��?k�x>d��>-o?T�9?����*)<��>���<U����UM=2R�=����+���J�>�`�>�&?� ��S�*����Z�=e�?̙�>O�>�����ғ�YZ��K&>>?�D>�y ��h�P�?�3��>t�X?U�����=��>�#�=s-;��l�>���;�����ѻz]���Լ+�[<2XD�RbZ��&
����;ȵ���%�=�u�>:�?않>QE�>�B��,� ���Fd�=�Y>"S>�>�Cپ�}���$����g��Wy>w�?�z�?��f=��=ז�=�|��)V�����������<��?�I#?]VT?╒?7�=?�j#?Z�>�+�EM���]��9��ʮ?U�(?�l�>���	¾�l���-�6�?��>@�c�´��J)��dȾ1��>Z(��Iy�q�����A����;�s�g�����?�ƚ?����;��K�R"��ԋ����M?���>&n�>ڭ�><�-��_�zj�{R->9P�>�pX?�>[~Q?�v?v]?]�e>y1�䭿!y���Cͼ�f�=<~2?�Rz?�܌?.�m?o��>8j4>��&�۾�f���5o�ho���f�,a=��->ʊ�>��>~\�>��>�����駽�v+����=$Q>/��>0��>0��>y\>��,�G?���>�`��-��J�X�0:=�	�u?���?c�+?�=����E�]B���G�>�m�?���?�/*?ɿS�j��=c�ּ�ᶾ��q���>ܹ>�1�>�ȓ=CjF=aY>��>{��>���_��q8��lM���?�F?Y��=��Ŀ��q��nr�*f����5<@g���We��8����Y��"�=P����R����Y��l���}��Wn���ƛ�H{��
�>�=���=Ƌ�=9r�<�L⼜q�<~�L=��Z<^-=)�v��c<<�L���P���l��V�X<"�M=�׷��D̾}?o�H?}P)?�rE?�!�>�t>LJN�	x�>�W���M?��M>��Q�H���<�� ��Wȓ���վ��վ�3d����Ю>c�T�n0>)m;>��=34<Gz�=�%r=��=����|�)=h��=��="ȣ=�='^>�P>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>l-`>���;�nm�P[�8mH��_��yd��)<6?�x����>I/m>4�������b�>Oh�>㺑<����^���7c>Zx=�E>�;g=A��>���=��q=ô��PB�=JÈ>���=��μ��=^gQ>��	����A �=�~�>*�>[ �>�?��/?X�d?���>E�k�H�Ӿ�Y¾�>���=p�>K
�=�^H>�>��4?ָD?�L?�m�><ρ=`B�>�2�>��)��l�)e羉7���\�<���?���?�n�>�T<E�<�� ���<�:����2?��5?� ?ft�>_��jf �w�s�0�=o�'>h꡻iw�"*�����m�g�D����>'��>�d�>D�?�Y�>�Z5>�_�=T?�>,=<�b���O�=�������>t�=)ut�_�컫�m<k�y�)�=R�i<A%�=n�N>�y�<a���e��=舩>��@>�Y�>]u>�t���[>�#���5�"iS>SN�ss6��-6�ٻj�����5�����<E�4>�����x���>�I�fw�=.�?��?��>c�;�;������0d���֨����=:��=�O���P�A�I�4�#��_��/��>Q>|�1?��	?�yL���)�o��=� �w��P6?"
��c�>�W0��a�)��C8���we���>yQ?U��9�K> u!?T�^?Aև?�ҏ>�ՙ�!���;�< .��"�a����U2�����=S�>�\9?��>�پ��J����<J���R�>�Q^>P|Y����5�ž�H��x�V<	?��;��Ծ_y��9i�;§�љ@��27�r��>��[?���?��c��M���{8���������w�>_��?���>5R?��Z?.�ؼ��Dư���>>m:>?I�?��?8�>�����>���>4K>�2�?~�?Ϯ�?)���lT?j��=m^�>EN���n�a�>֖>��='?�#?rN�>�*����e�����	����&��=��=�ʦ>�k[>m�=�#>�*i��&�=/!�>�2Q>�5�>%�c>dA=�i�=�N���A�1X?c�>��&>�0?�s>��=�gs��=N�_P����{�'���p��c���If�;�彮a�<��� ��>��ȿ	�?�w> :����>Q��5��s^>zä>.�<�b�>��>0[K>߃�>�ӊ>�E�=gǚ>E�h>Tp��.>�����
�jO�-=�Z��(2�>��7�hD�����pY,�|c���:��h!��]�~���lb8��I»Ҋ?/3���Y�͇#��@��\
?�;�>��2?�џ�*Ԙ�fSc>��>l�>AS��"��2⊿�Gվ9@�?s��?��b>��>snW?�.?��-�q�2�[��>u�^�@��d�T`����G����
���ýǼ_?,y?�)@?��<�cv>��?�y$��ɏ�<�>�-�Ka:�ԟ%=���>9��|_���Ѿ7�¾1#��J> q?��?U??¯[����X�?>E�6?�,#?��x?��/?�	;?�}(��*?>�:>j�?���>��*?N�2?Y�?w�>>�!>��<=�E=@X��<^�������I����<�Á=G��<�k�-��<��b=���;�(
�DY+��f<�*���=z)�=iRG=}C�=�c�>C�Z?��>�Ah>�jB?���Lz,�2﻾tU3?|\B=CM{��ؓ�U��F ܾ���=�/g?���?��R?��\>�GH�.�>�%� >]��>]5+>	ڐ>���>���V���)=��=�W
>���=�N��F����ω��7�<�+>-��>F�y>�=����)>�ݢ�F�{�vd>�Q�	
��g^Q��H�N�1�u�h��>�EK?�?iR�='k��Ә���f��(?�(;?9�L?A�?�&�=��ھ�9��*I��]��>n�< ����� -��Xt9�ez
:ҡt>�V��"Q���^>�.���ݾ��m�4I���"�n=)���A=r�
���־m�~�]a�=�v>�罾y�!��i������ZI?��X=桾��Q�08��k�>�>���>��*�9Ea�A������=�%�>#�8>�Mڼy�O-E�� s�>�TE?�^?:R�?G���Us��B�r����䡾K���X�?�y�>�3?-A>a�=�ױ��#��gd��F��u�>s�>��4HG��s���$�
`�>�~?��>�?�R?��
?�~`?'�)?/?�:�>A���	��D#?ă?��k=�2�;��{�YE���)����>�>?�Gc�?�v>A?$?c�?�b@?h2�>��=��þ�&���>�.j><&H�?����n	>�e?��>�xL?��v?�=">��=�ծ��^7��>ۤX=D�2?l�'?�j�>4�>UC�>6��wl�=���>��p?�2�?�*q?���=���>�jF>�A?��=^Y|>�r�>��!?
�N?�df?�I?A�>V���1˽f�Խ�cp��(<��~� <��f=�0p���C��(��H-=�Z���߻N�N�O:G���*�ɩc�$�?<
��>�w>Ό���8>
Ҿ�������'>�R!;䗒��{�d�Y���=Փ�>�"�>]Nz>Ψ0����=��>��>p��O{?V�?�f?��<�Ec�D�׾Y�X��s�>5DA?!�>�Jc�����!i��]�=��m?�!U?TN�x� ���b?�]?B��R<��p¾��d�ŉ�� P?�?PE���>�~?V,r?�h�>Mzf��|m��e���f`�]�g����=ZI�>�+���c�zn�>��7?Ƅ�>�_>,<�=:�ھܼv�n����?�Ռ?���?�n�?�z,>ƹn�;�b���O��
m^?B��>�^��[�"?�Y7���Ѿ�������Zjᾣ���hF��C���2���d`$��܀���нB�=��?7pp?�vp?�`?,�����d�0$]���~���V��"�>Q���D��iE���B�`Uo�?��6ז�V=.���a`�?9?��P��?�>	���rLC�6��8�?�/�=y�Y=j+���H�P>���=��A�x�=�}+�3?m�>��2?��M?������J��G`���)�|h)�X�>l$z>.!�>ES?�u�!* �,B���Л��+>#�>�U}>��_?MT?bq?I���.��v�1�#��$�~/���D>&�>�x�>P�Y����`��<5�*_��k��Ӛ�UT�H��<�3?�y�>�}�>�s�?4R�>���8Ľ���s�><��3�:�>�i?��>�"�>��><����>Pii?���>E�>�׍��3�U�f��̽�?�>5�>�$�>���>����4[��n��v�L�)��kJ>%�h?[!s�2e=���x>�/K?��K��;>e�>�4Ҽ�
��2���:�J�=�?b��=��>~x���e�9�]��܆�W?_?n��������.>��?���>쇏>͆?h�>�ܦ����I?�da?JF?�^7?�H�>�B��A���b߽+�V\_<��>��>2*�<��=f7��;�@��F��=u��=�y��N�93�<s,t�E�S=���=��'>��ٿ�I��Ҿ ��� �I���0��2b���E����*��7�����?����N�[������]���G壾��?X�@�v��a{��Jm��r���h*����>�^�DL�[��>I�lN4��O���پ��$��j7��zh�~����&?��h�ƿD��&.�(Q?��?�{?��GQ"��7��*>G�9=��;��澫����Ϳ�ꔾ�\\?B��>�����> J�>X�^>Вp>J�|�P���t�� ?�-?��>L�t��ɿ�m���2�<k��?N@�bC?�*�_���f-�#?�l�>`�a�!�Ta���]��7�>t��?#�?�=��n���"��jx?���=�1��U�[A�=A��=�5������n5>�0}>/S��k�׽J����y<� 7>β<���	�콜�o=�œ>A䗾��!Մ?�z\��f�r�/� U��*T>��T?�*�>;�=��,?�6H�*}Ͽ��\�+a?�0�?Ŧ�?��(?mۿ��ؚ>f�ܾx�M?FD6?���>�d&��t�̅�=�-�!l�����'V����=���>ƅ>d�,�����O��<�����=���0eȿ`��}�$���`<�!=|�#��8��M3�ѱ��oq��bk�Jgؽ��=�P>:�x>�"�>n�@>��?>W]?�>�?	�>�*>� �Jն����Q�޼[�o�o�C�ʻy�^1�W9��A�ξ�K農�����J��f�־��5��"�>��r�"8���+�P�_��Jz�ڱ�>���>	��w�����>�^���Q���8'���(>��}�Y�J��h��e��?�`Q?c���\5)��3־H)�=���52f?���)=�0�M����>�I��Nˆ>�k�>�����I�N�X��(?��+?c{����;�*�=wR��O���?_�?��=�����?�� =�5��=�'���0>U��>q@Y>�����#�˘?���?ς$�9�Q�O>�y��G�:��=Ó�>]Ĉ�6	�ܹ�=	]�>�xo�m
�QOD>c�����Q?[��>�J�����'���S���A��?	J ?�!|>�
J?��O?��E>q���%U���8�=tQ`?�"g?��>�l��o�;�t��ee.?n?%�E>��\��1Ǿ�b"��)�,F?�U?#,	?����l�c��q���b/?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?s�;<��U��=�;?l\�> �O��>ƾ�z������1�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�C��2�?�*�?Pj���1E<�l��Km�+���k#�<d�=82������>(7��Nƾq�
�Z(������Æ>��@�"߽��>��@�<�῝�ο�8����̾��m��)?�V�>��������Vl���t��OF��JF��$����>(>����.���Us��U:���;kG�>s�Ƽ(�z>�\�9���֝���a</%�>Pv�>;w>r٣��#��x�?[v�Gʿ<������o�a?���?h�?��?zL;�f�˃��к���A?]q?�-\?��y�3qs��
3�Vrj?� ��#�]���4��mC�')Q>��0?n��>�-+�U4�=�>'�>��>В.��TĿ^z��e����5�?���?d�龮��>a�?�o-?4�4��'e��K�)�����+A?��4>ڗ�� �!�-�;�H8���?�-?k���>�ɳ_?;�a�=�p���-��Bǽ�ơ>r�0�0X\�#J��^|�He������y� ��?\�?��?�����"�2-%?��>񖕾W,ǾF��<ce�>X�>e&N>	�^���u>����:�@l	>;��?�x�?Z?�������	�>$�}?�ϸ>�q�?�o�=�5?}j�=8�Ӿ=[��`�>�U�=����a��>pJ?���>_1�<��]B2���G�A��W���y>�Y�>�"`?MJ?��`>"���o|�$��e�S��!&=�c!��g�T���}>>��>{ �=a��� ƾ��?Kp�7�ؿ�i��0p'��54?.��>�?����t�����;_?Kz�>�6��+���%���B�_��?�G�?=�?��׾�R̼�>D�>�I�>A�Խ����b�����7>+�B?j��D��v�o�r�>���?�@�ծ?hi��	?���P��Ua~����7�]��=��7?�0� �z>���>��=�nv�޻��W�s����>�B�?�{�?��>!�l?��o�P�B���1=8M�>Μk?�s?�Qo���g�B>��?"������L��f?�
@u@`�^?*	4�蚧�g�¾g��/�I>kNL>1�Y>��8��To=�0u�������p��=�S�>�h�>(z>���>̿>�m>̆�w%'��ǥ�/����(���o�%��֗�6	�ʑ��r���t��P���<JW��|��3ڽZ"�Y��n����	�=��T?��P?[�n?��?�[�q�!>���1=�<��"�QԄ=�ׅ>��2??�L?�^*?� �=Y#���d����Z�������>=�D>U*�>�>X'�>��F�"E>#�?>�j�>��>�)=�Δ;��=�GO>�*�>$Q�>;�>a=>��>W�ǿ(0����>�����F��ȫ?�ؾ_4����"����=����ҾDg?�+?��r�6�߿��ο��C?��i���h9=W\U>���>A\?��>9׾�[6>$Z;<:�ҳ��{��>b,�<����Z�M���->�?G!�>�խ<�B�q��l|A�ܓ��� �A�>?�޾@�
�~U1�	h�W�ݾ3p>�i�>���:_F�n���ǂ������=��4?*�>��Q�J��e�K��
��9V>k�>��<�=�U>T�=�WK����QU�=��a> ,�>:?�d>VD�=���>ʣ�|������>!�=>r�,>�(?S�>˃	=)�Լ�DB�o.���=�I�>�q�>��N>0.d���R=��>5�f>��6=O�"��e���i��wU=�dh��/��}�Q�f=�X�W	�=� �=^W���,��A-<��z?�����i��XR�����7?��?��=�D=i��bk���I���j�?u�@�Ę?��	�gV��0?&v�?*w��Ş�=w�>ʰ>��Ͼ��F��?oEb�Ғ��F��ӢK�~��?���?�S,�`���rp��`>r�-?����~�>���T��@Ά��Jv�~v=LL�>��H?ɮ���U��C>�-�
?Oj?���ms����ȿ�]v��=�>���?�֔?��m�����?���>���?[=Y?o�i>ـ۾\����>P�@?Q=Q?��>N��I�(���??��?A��?�Q>��?�Hk?Ɋ�>z���^@�	��j���b�]=���<uˇ>��">�pþ�Q����������l�:_���u>EO�<���>R��uA����=��޽!矾����>�1>M�@>C�>L�?���>�{>��c:Ջ]�<04��7��8�E?k4�?\"�%�g�3�t����<	i���?�I,?k/y=ƀ���>��S?�?Q!i?��>gn��d���
��.��0>=i7�=̓�>���>S�T�?�.>;O���ǽ��>
��>�z=�;��M}P�X�<J3�>.�?N�>ݹ�=Җ ?e�(?�i�>�X?%�
�T��Z��˞�>P��>�C�>P?�u?I��ˆ]�u���	l��u���� ??��?�{?<�Y>`�y�������z> >� ��v��?�*?����+5>��v?v�r?�<??�s:�%��~����>�f�>�?�/g�u�1�@��\}��N�>��>���>|ޠ�-�>��F>_?-������?v�L?��>�E)�QQ��t����ӕ��6>���=�d=?Q޽:x�=�p>jdA�Eq>��x>�(�=%S��i�)<D%#>�L1>d�>&�<>ӫ�����<)=,?t�G�)ۃ���=e�r�HxD�<�>�IL>,����^?�l=���{�����x��(
U�� �?��?Ik�?z��5�h��$=?
�?_	?�"�>�K���}޾X��rQw��}x�Yw���>���>l�l�d�2�������}F��v�Ž&e=	t�>r�m>���>���>fC>ʥ�>ã�+>�\y�.*�p�g�K�:�X�.(���V��b���-$�<<J��}J�fd>P:�Խ�>
�?���>�z�=|�>��=���>d�6>ֹe>	)�>�B�>2{�>g�>�bi�z���>bI?�1���X7�Z�������)?9p@?�"1?���=-o���Z#�?r Z?�J�?�
=���kE�Mi?��?H����>�.
>x���Ϟ>2q��ƽ4��G�9�>J���d�Y�Q���+w;��>��>U�g������5���z\p=@n�?��*?/�*�ʔQ��Jm��Y��TR��ᦼ�[��%��w�#��p����𫃿T��X�$�.Q=�)?�x�?�����$����k�
?�Ysj>�I�>�$�>{�>m�I>���9�1��O`���'�v���E�>��{?\�>�M<?�lD?��?�ty?"�?<)�>+����#�>��=5�>l�>a�4?�`?)9?�1v?eJ<?Z�F>����
���)���T�>bɦ>?m7?&?�����ȭ�O�����">���� ��k.��D�=�#��6�=��;�H->O�?I4޼�!��'�����=� ? ��>�b?^�A*������;o(>�|�>��f>�U%��`_�*����>V�a?��+�<h�=��->��=�M����1=�ԍ=U}����&>�\=[�o���<�/5>�D�<9
���a8=�><�^+=��=��>�0?w(�>�g�>�f��R�Fiƾ·ֽ~��=�v�>���>O���'��pP���>j�>�>/�?]�?�/�=CpI>h�%>��ʾ�F��0j������t��$%?U�,?=�6?9e�?��:?+?޵�<-�0����L�d��bO�'I?=�+?[�>����Ⱦd�����2���?@(?��_��6��>)������Խ�>t/���}�%����%C�V�f��O��D����?1��?�9�n�7���=%���^���$C?�_�>��>��>�(�mmg��!���<>�d�>��P?���>Q�J?>��?^�]?�>=:�����4_���2H<]'�>7=?�Z�?��?�!Y?zT�>dj >�� �n���(���ϊ��a��0|��>�>&=s>�O�>k�>쇗>��=�� �����ZX��j�=͂>Rt�>���>�`�>nCW>�S��;�G?+��>Z���������Iă�[�<�\�u?���?��+?1�=z�W�E�\,���>�>�e�?>�?�.*?۪S����=׼�ڶ���q�x�>z�>a'�>�ؓ=[tF=~?>���>��>Y�6W�ir8��HM���?nF?]��=w�ſX�q��Vq�-x����_<�ْ��9e�6ݒ���\�y��=a���K������|�[������̓�m���"M���{��\�>�؇=%��='M�=���<anʼ��<2}L=f��<,	=Onm���{<�
6�am�����4���j<��J=սл��ɾ�[}?�H?+H+?��B?2�{>u�>-�5����>�́� )?�T>�xU�hV��^6;�WX�����ϣ־߭Ծ�dc�*b���	>?M�ZQ>�2>O�=-X�<Ef�=�b{=>�=2*$��=7�=�x�=�L�=���=��>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>r�o>1'=�"L�3���7g�<�a���u�,?jF�!������>��P�����ѧ��=1y�=N��6��g�N��l=�H��k��=/�=!�F>C>;`>�"���=�6�=��$>#1�>3H=�=�ȼ�w�<�	>�R�>�)h>���>�?�B5?��j?XW�>�8k�{ҽ��xҾ�tx>
H�=-º>�:=�Y7>�ı>	c0?+�>?�O?���>軄=�+�>�ͧ>_�+��f���v���J�<{&�?r_�?]��>&�#=A�:��q��=�mT���S?+�2?c	?�a�>Ov�f���eo�v�e����=���>1�S>�X����	�W��p$�,Ǿ�8�<��>(��>��>S/	?b�>��F=�c�>�}>�ɦ=lg�=�)�ʿ�<�8=zJI:�!�=ݫ>�k=hhY=֛:5��'�ػ˞�=�]�<�^.�߽`>]8�>Q>��>0�>�����KG>ꢜ��cQ����=AgȾ�	�ݫJ��G���(�|�S��)>�;>���t���&A?Q?�=�ۧ��]�?�,x?�_�>{�¾�ך���ֽ�s��^ ��	�=��(>i��V���S�������>�T>���>���>+y&��+�$�L=I@ܾ*�^�>FM��쑞��*�*�Y�Ș�Ɗ���d�>_�=RQ<?;�p���W<��3?��'?;"�?�,�>Γ�<��u�i�R�$�ڼ:�F�b���ǽ�� ?[t;?�.�>��"�{�z���˾�]��Χ�>� F���O�=���h0�A�P_���9�>"ҩ��5Ѿ03�^������T�B�.�o�K�>��O?�߮?�5a�&^���O���9���E ?w�g?X��>Z�?l??�e���P�瀾]�=< n?��?�%�??�>���<R�=6e?i~>�3�?���?��?�[��O`H>�>�>�{C��5�1e,�2��>���>ZG�>�?��?f���6��Mk߾��:L����=�\�=�2G>�&�>���>�YS>H�<*�=7A�>s��>;�[>"�>�<L>ds>��u�)^׾��&?G�%>ߞ>�):?�\�>�>��υs���=�2=��(J�����<r�K�a�={k�<
�� L�=���>#��E��?n�}>����|�><&�"5�L�<��>sD`=jb
?gJ]=
��=�;�>\�=>s��=pc�>�>����>Z����?�[��Z�a�Ⱦ��>��0��A1�cG�TBd����S5�a 侎�e����x�'�Eip<�6�?H��b[[�������u�?��>\�F? �S�2k�G�a�߄�>鳔>�V�6ԛ�������ľ��?��?��b>���>�X?:�?T�/���0�K�X�,�v���A��Mc���_�_��y���
�d���G_?W/y?`3A?jx<S�y>�+�?�z%��t���=�>�T/�s:��:=�Z�>R}��A[��@ԾN4ž(��U�?>C9m?Ȝ�?8r?*LQ�Ѝ{�jJ3>9?m�$?BJ{?��2?pB<?9���2$?��;>�i?a?��+?��+?�u?x�A>!V�=Ɓe<e=�͎��U��("���ѹ�嵹����<"=h��<=�0�<�x<q���ֻ7O/=�S��mg�<�2�=魓=��={N�>�ZU?^n�>��>z�D?m�ٽ�;�n����:?��Y=�핾I�,-�6龊�<��L?'z�?��J?>�x>��G��*�w%5>���>!n�=��.>YU�>#J�2b�C=B=�"�=E+�=/�_=�=���VA����������� 
>o��>�}>���C�,>m�|�p���o>p�R�2���UM��)F�_�1��?w���>)�I??'��=��羔㐽d��n%?�^=?M�M?\,~?�y=W�ܾ"9��M�^����>�P�<�
��S������;:��<,3r>ۺ��Q��+a>ص��徢�l�o*G�V ���h�=�
�Z?7=S��Ͼ������=}!>R踾�x�����1��J?'rn=b���^��+���0#>L/�>,i�>�4�H\��@*A�a��v��=V��>�D>cݼs@���H�o��y �>�G?/�i?���?�M��Yd��SG�����ד��M=`E?��>-?��K>D"�=�᫾���"[�BN9�1�>�3�>Y���;7��	���	�R'�w#m>Mz�>784>G:�>��J?t?.�b?j�"?Z�?0�>��l�����$?>�?,®= ���]�ˆ?��/F��>`r#?",��Ց>��?��?��&?�DJ?	w?@3>������=�qʘ>�$�>cX�u	��	�h>�O?V3�>�C[?���?�/>�3�M���Ԥ���=�>��0?Ue!?��?�Ϻ>Q2�>�ˉ��?b=���>��e?��}? �i?U��=��>��U>���>f��<e�>�]?��#?٫J?�yb?�6?�Z�>e�<���a<��/�Ž+���Ι����=�-=������!��J���r�<�1���R��B�=/�J��~��}5���>f;Y>�Pz����=��n�G$m��-r>�~�=gq��􄍾�Ԣ��{->`C�>���>���>�F����=an�>���>:�
��* ?�"?a@#?�� �x�ћ������^u�>1@?ͫ�=�9P��&����n�o� >;�}?�N?	A��s%�Y�b?=�]?�d�S=���þ��b����9�O?^�
?}�G�f�>c�~?��q?ȵ�>��e��7n�
��jAb���j��˶=�r�>X���d�n<�>Ț7?2N�>��b>��=�r۾��w�_q��$?��?u �?���?�2*>�n�G3�bC���4���]?̅�>`ϧ���"?�G�'�;l�� �����=�����+����f��R�%� ����ؽ�-�=�s?*�r?��p?��^?�@�TYc���]�Ƌ���U��f����rzE�E��=C�t�n�M�!���7꙾�vE=X J����+�?�?<?c=R��>�<���z�/2�>kEܾBJ�<�u"=ݮG��c>�>K��������4�?V�>�.?%�G?��p��a�y�`������D�$�>+�>A-�>/��>�ȴ��b��[\�&�<���5���=�h>[$`?�	L?u4s?�p�,���x���4��:4����i��=2 >΍�>	�?���������7��-m��������*��jK<��6?�x�>F��>��?� ?���'�;�[��J��Px�`��>Xg?4�>�+R>�=½L$�"�>#�^?��?˶�>Th���~��&i�-� '�>
��>i)?�9�>h�2��gU���}��`��t��z�>�Z?��p�Q�vG>NI?��=nƊ��tG>�q��6�fX��������;Ei'?1�a>e�P>�O��M վ:����V�1O�>�F'?W2�����~�?��.?�� ?�{F�P��?�K>�*��b��+7?�z?p�#?��/?5�#?�rI>G������gy�J�N=ϑ�>_M'>#o�=�Ա=��B��B���g��"��GH��$ҽ�+�f�<�����}���(>2�忔�M������
��O����Nپ��Kh�W:4�=5���ʪ�2v��*���������bZ����i�v�՘@K�@�9�ϩ��L��^�]�*�a��y�>V���O�T�n���=_Y����7�@��3$��Nb��M�������&?3v�L�ÿ�%��K۳��
?+c?��k?��=�����I�ۛ���X�� ��������ӻʿ:�Ͼ̎l?�|�>�Ⱦ�D�<�!�>��=jd#>NA}>�F��� ���

?n�G?�� ?�D���_=���F�َ�?{B @�C?�����Qξ42����?���>��?��~=�Ʒ����Y�
?��?*8�?%b����/����D˃?��>к�M�z<a�.>t�8�e@��_�=N��>A5�>0ם�{�]���(���>�	;>��4<}������\�=>��>���<�&��2��?��[�$e��</��$��?>�U?J,�>2��=B�,?�!H�9Ͽ�[�ܧ`?���?���?z�(?��Ǳ�>��ܾxeM?M�5?4�>�G'�X�t��"�=�輘�w��@�/V�U��=��>�>�,�����S�iw����=��B�ʿ5)�V�"�r�<��:#"���ұ���rp���� �������-�=j��=��>晌>l�G>{�U>�i^?gx?߰�>)O>_I��^Uh�E#��vk:�≾:A�����j�EX�őھ�4߾���1�#�D!��U��u�>�=>OAW��L����0��#[������2?C��=�'ᾝj.�g{�=�F�� ��x�>�+��V|þ3�I������p�?��j?�����l��o��>=�{��Iv?S�C�e��@�u���\>�Y|��{Q�ɵ?%�z=�����n]�(�z�9�,?�\%?M�u�-E��%ߙ>�!��y��=��O?Ԃ?������>�{d?��3=S��uƏ>���=�0�>��>>�C��D�_=/k0?X�Y?7�i�:5���[=\c���2���?h>ư���L��O�>Կ>BC�<��_=�>��ֽn�S�T?9ǝ>�(�959��g��m�=O��>iVP?�f?�s�=!pY?��S?�>���fD��p����>p�Z?�YV?�^�=ͦý� ��⮨�?��]?g>ҟ����;,���	8?�-=?̼:?]����0��*��]���/@?\�v?�R^��l���DdV��<�>��>r��>z�9�\4�>�>?��"��/��6����R4�ػ�?ғ@)��?ö9<	��o�=G$?|Q�>�]O��ƾ�,��?���[�s=�>x���rMv����@y,�n�8?Χ�?�z�>�v�����=�=�I��?]/�?���Y�������'f�������-=渶=�c�⪄����A6��0ž�(�w薾3ߙ��>��@��Ž��>�;<�n��u!ο$T��svоN~_��?��>h����6��Zg�D�n�>�`FJ�QA��&��>+ ?>��[=f�]�l}s�VV�*�����>�Oý�2�>rzw�����\��+�=�6>���>�G�>���<3���ɔ?"���ǿ���������|?�n�?7��?j+?��\��LB��e^��Ŀ=H�?ȎJ?��=?w[U�����ظ=U`?��߾��_��:�:9��G4>�"?��>�A;�[�N=��q>�D�>�L�=G:C�����Z3��$��8�?h��?mB׾��>	��?^=?�n�qM�����x�S=Ͱ.?�B0>8�u������4�}dh�E�>��?
�	=����1�_?Y�a���p���-��ƽ+ۡ>V�0��c\�K=��+��YXe����.>y���?^�?u�?c��� #�J5%?��>眕�o8Ǿ��<i|�> '�>�(N>GK_�d�u>5���:��j	>خ�?�}�?�i?ƕ��@����W>��}?(�>�
�?�-�=3��>KB�=i���D��">���=��5��;?��M?���>���=�e8�՞.��E���Q����D�C��\�>�a?H�L?��a>2����9�M�!��Jν��/���߈?���+�uq۽0�4>��=>��>�*E��)Ӿw�?��P<ؿ����
a&���3?��>�Y?���Wv�ﻥ`_?��>�>��볿���� ����?��?Y�?8׾���&>˫�>K��>!�н���#R��B�6>��B?�������o�|��>���?�@���?uLi��o
?�p��ȷ���-��:��b�8�#�>�;?���X>��>�#�=>:k�p ���p��8�>Ԛ�?<{�?|�>�Ai?U�f���H�L�<`��>��j?u*?�Ǽ0�U6>x?	������R���^?@�	@�9@�/^?�1��i�������bվ1�J�������=o���>>�<��=ݏ��C==@��>ˡe>���>5�>vi->ڵ>Ҟ����,�EX���.��T�Z�=MG���%�7�$�ê¾�d�����G�b����Ͻܬ˽= =��\I���2��}���1=0�P?$�C?�a]?��?�ʺ�,z>tR��V�=��6�}C��)�<��?��<?��>?{OJ>�m��<J��c��<:���w�h��>c�>���>*�>&��>���=�v�=ꤗ=�]c>#�=>��<�4����=�Ig>z�>(=�>2N�>���=g�~>G$��ed���%��N���D7��_�?�f�����IF��o#�}��M�G�'�|?�b6>�����t�󪰿�R?xl�V��3jO>`�K>��%?�]n?�?�2�� �>�t�>(x��l;�Uk�>��G��ͽ��V�z��=�a?��>z�r>����6=���Q��L��l�>U�&?�>��0:ν�q��3�@���7+>Fm�>��=U3�MW��zv��Ї�:m�=�b7?���>�&�Ɋ��4���r0��_�>���>n����^>�UH>��ڼ"��TQ���v���=�<N>B?�4�=
�@>��>Y`��7(����>�u�>§>e�7?�	?1B����<ٸ��oخ�Iף>ʶ�>���=�<>��)�XS>L�>���=����DL��> �ɬS�P��>��%��,ݾ�[���/ >Cl�q.>ɪ�>.�!�WǾ0���~?���䈿��:d��7mD?V+?�=�F<��"������G�� �?^�@�l�? �	���V���?�@�? ��`��=�|�>!֫>�ξ��L�6�?��Ž�Ƣ�2�	��(#�IS�?�?�/��ɋ�Bl�w7>�^%?�Ӿ���>���#��冿�s��=ú�>��I?���G�v�`�4�I�?�
?�m��m���1ȿfNs�1�>��?�?�k�񶛿�@����>)�?��Y?\�g>ؾ�c��x�>�K@?�mP?���>�\��0/��b?�2�?}��?��I>�_�?�t?k��>1R���~/��@&���=Pi�;��>�A>_z���-F�*����-�� j�z��Igb>��"=S��>�M�~Y�����=o����f����g����>�q>�J>#�>?[V�>�Ǚ>�=�֊�t���-���S+J?�+�?���n�pe�;7��=�)a�D�>y6?b��;{WԾ�Ѱ>��[?Ot}?B�Z?�̜>0�љ�4罿`��%�<��Z>���>m��>b����+>�-��0��ڒ>�a�>��h;&4Ӿ�Ym�m{��4z�>�x ?�D�>W"�=��?xv?1�>�!0>i�.����_���?���>m��>�,Y?�Y?�0���&��א�Q&����,��5>��s?��?E�8>�������b*>j. >\;>?r�?YBe?r�ʾr	9?��?� Q?��
?ˤ�>6����߭�%�p>X�>s?��Ӿ�Qz���w��=���=�>T��=�s>OH��>2Y?ئE��z��&�>O?0#0?���簚����:�>y}���g�YM>%��>�F�=�,>b[4��f>��=G�,=I}¾2�d<|��5ǅ����=p{�>󎒽���=,?��G��ك�7�=��r�xD���>�IL>G����^?l=�"�{�H���x���U�� �?}��?k�?���םh�|$=?��?k?�!�>K���~޾���)Pw�~x�Cw���>	��>��l����������)F����Ž�5�,��>��>�	?�B�>�V>=�>�Q���Ŵྂ��n`��� ���)���#�HD��1̾B�2�Z��yᦾ�ʁ�D>l>C���/�>�T�>�Do>�p�>���> ߼�,�>�N%>q�T>,!�>U֙>�q>"B�=J.\=	,��?G?�㽾���k����� �D]U?�Rq?���>6�,�'�s�k$��YdC?h �?d�?i[�>	5o��~���*?��?�lc�:��>�i�>g��=���=kj����.�>��^�Y��>-��=�(���i��k����:?
�>�=��?)���B�����SpU=�݃?��(?�)�6P�&�n�\U��S�RJ���c��Ţ���%��hp�����m���O�.)��p8=�O)?x��?5� ������2i��>� �h>Xw�>TT�>A�>�JH>+{	���1��+_�2�'�胾�}�>@�z?���=��V?S#?���>C�Y?�
�=�D�>�}����>_/ƽf��!�>):]?�>?�0?B>8?�@?W^6=#�����P���3�9>�3?�5?��?��>���������$���t$��WG���!>��>�����	�Z=S��X�?�/��>��B��=���!#?/�>3*"?:� �D��hb4>1:�=�����?]���W�񰘿,�y�U��>���?Z_�w�&>y�H>��w=�-�]��=*� <�3m="G>^Ȑ�@�:�&�x=lo�=���>U8üYx��2�=Z=)>���<x��>�*?qW??pb�>�����6��5�>A�!?4��>��;>�ǿ�c���6���OS��.�>o�{?��?�N/��=#>"	=Hg����׾�u���7��@�=I�?�S�>"O�>��?��?��#?�FO>��v�����}�����<�?ݑ*?��c>��i}¾{D���.-��.?��?��^���o���W����̽�q�=,n4�lT�,+��x�;���C=MN��c��٭�?�f�?ڼ��;<�Q.�Ĳ������??P�>Vū>2u�>_.�6�a��!�3�>��>U?��>}V_?�p�?Ec�?g~�����z���5���? ���%?��	?<L:?��u?'�?T�7>��=m٨=�v��{���٭���r��zLJ���=A�>>�w�>�W>��}���r�,(��ܽ(>[��1�>��P>bw�>n�T>��|<_�1�S�H?���>�i���a�Ia���v�:̙<�*r??%�?�===��3�r���X��>�_�?���?��/?�6Y�IQ�=�	������`�j��`�>X�>�$�>�	=H��=�Z>]��>�7�>\����`�/�ya;ѹ
?FD?��=BQ����w��쑾�i���yj<�3���Gj�����l�ɞ�=�"��4,������q~��߰����w�վ����U�A��t�>P�2=Ԟ:^�=��<���<���=�r�=�#H=~�<	*���p��`<�1�;�)/=�R��<E���=8���I�˾Sz}?+�H?�_+?-D?�9y>��>R�8��Ė>�̃��?n�T>�L�k����z:�������Mؾ��׾�4d��ϟ�7�>�cF��h>p2>pj�=Q�<���=Op=◌=��3���=���=�@�=�Ĭ=���=��>H$>�6w?W���
����4Q��Z罤�:?�8�>g{�=��ƾr@?��>>�2������xb��-?���?�T�?9�?@ti��d�>L��}㎽�q�=Q����=2>���=z�2�U��>��J>���K��J����4�?��@��??�ዿ΢Ͽ*a/>� F>��= WV�h�'�m�R�U�R�Јc��?s�>�[l��~)�>q-m=���zǾW�<*I3>���<v�:���S�wS�=�ڌ��f�<��9=~&�>�{H>:��=�՝�	<�=��=��=>�?>H�<�I���>�u��<e��=�k>�>�A�>�?\b?�i? �@>�'��6���;���>>:�>L�P>�;>m�=��m>>$?z�9?��G?�%�>T��<�j�>t`�>7⾠�c���"��rᾒ����?�S�?���>W�!>�$F���h�o��묾�E�>�y*? �-?M�>�#��u��B�	���b�.�h������}$�(9D�$�<��������M���=g��>g��>h�>w��>���=I�=��>���=δ�<x�/=���=��Y>}��=��<������3��b#��<���=� :�[��<'
>">�Y+��x�|]�=0��>�8>&I�>m6�=ݤ�	L>&Hھr�3��>>��+D�!2U���l� ���,ҽ�>�%>8��-��3�>��>_54>���?R�u?��>x��Ua� ���������¾cj���=���/�7�a� <?���S��>Yk>�Ó>`#f>�<&�x�5�߫�<�C��k�8���>*v���^�?���h�"������+�m��~�A9M?\��� �9="n?�_H?��?A��>�R��� ۾R4N>�n7��n�=����F��:��^"? 1?&��>3޾�EC��ľ�;�����>��4��P�w����0�2w�7q��Jƹ>�(���	ƾ�x5�����e�����=��m���>�EM?��?:�h�0Q}��L��!�6��T8?Ыg?kO�>-�?3�	?�İ�r�ҏ�劬=jtl?���?�&�?���=57P�g�~=�n>!�?7e�?�#�?�4H?>���WV?�b�K��04��O>��>j�=�H>�i?� ?��>�K��WG�z%��8��%#���(A$>�?u>UИ>��>��4>n�>�Z�>B~>���>��>��k>��q>Rl>!E��[%��)?�>?a�>�(2?��>ֆ��ϳ�����5��[��Zb�!Cý�d<�j�=�N���<F,��.�>E�ԗ?�Yg>����D
?0
��̜��S>J|w>ȡ����?�=M>��h>��>��>rUf>l�>�sX>nDm�u����+����X��ti-�*o޾1TU>i� �g����ϕ�ՖȾyɾKX��'f�B�J���u��g��
=�Gq?�̽ư@�I��>����>H�>�jY?�&��􂯾�<
�=1�>�ݦ>Cc&�-s��������6�B�?�s�?74c>��>��W?��?ߊ1��3��oZ���u��#A��e�=�`�O፿-�����
�Q俽��_?��x?�tA?�ʑ<�4z>���?��%�[ҏ�p%�>�/��#;��w<=1(�>�)����`�k�Ӿ��þ<�^HF>��o?q#�?�W?QV���`�^[�>�P
?�?���?"�#?��.?3ʾ�D?s�=���>�^�>+�.?��:?�(?�f�>�*�>NG<V`�d���@�g�	p���<G7���=N�>mV����A=*M��8�<��c�f<�$>6�<�r1>���<O�=�&�=j�=�=a?���>#AB>ٗg?�i=�QھGH��@?>�<��O�����h��ؼ�*?>��K?"��?[�D?��ӽ#_B�������=F�g>� �=�b�>��T>rN<��M���I>��)>�ޣ=B�S��(��(�Y�Ѿ[č���@=��>��>c%�>��g�>���u x�bSo>�����>�����ngW���#��wN���>�T?(?�>=�]�5�d�c��'#?Α.?`�>?�`s?!�=)UϾY>��48�a�.�p^>�D��W��s���'����-��@�=�g>�e�����;�4>����:��.]��)����.�<#v
������~����Ss)�`pƽ�'��ד)��ܙ��b���0?�'�=*�L��$L�w��~��=�A^>c��>�=�;�{�<��Q�jIվ
�}=\�?�0�>��n�"���R�/ʾN�>>OO?�Gr?+_�?x@����j�~/:�F�����=@l�B4$?��>*N?Z�y>�]�=�ɯ���	�9]�%�I����>�	?����:��*������*1��tC>���>��P>Y�?P�E?X�%?q�x?��9?��?K��> '�%"���$?Q̃?��l=��ӽI�T��w>�%�G�S��>�+?ߡ:��}�>=�?C�?��#?1P?>O?�b>�����:=�lÙ>E��>��Y�DO���VZ>w�K?�+�>
�V?3E~?�\6>��0��G������J�=��0>^L-?9�?�?���>� $?0ľ�Y>��?��d?UZZ?���?�L�<G�>�t?֡�>�fR=��	?�j�>S��> �n?%��?f_?��L?� �=ɉ=sdF��P7����w������>j��=�B�>	��r�=�16>g����:�c��������ػ�l�9�%�>���>�֔���4>ұr�� վ3��=�n>]�tu��*�	��&�>F��>i��>P�=��d�4�>i�>���>��?)?H
?��?�G�����G����y�[�?�O�?ת->��o��3����t�F"�<��?J&�?�!��"�>�b?��]?v�=�F�þ
�b�d��
�O?��
?��G����>8�~?y�q?���>ͭe��,n���X/b�%�j�q6�=!`�>�^���d��6�>n�7?�C�>J�b>�Z�=lk۾��w��l��(?R�?���?c�?Z*>S�n�0࿩�ھ>w����^?�?2�⾩�1?�܁=`�ƾ׌Խ����;��o���^b���M&�$��p����z�����p�>P�?�f?Q�t?�V?F���BJ��Q`�"�v���K�D��Gk� ?;���I���<�Ywm�?���^��Kh�֕k=�s�.F��O�?�+?Q��K�>���_7�%����2>�������Ƅ=V@(�{�<�@k=��e�&��"�� ]?���>`�>�:?ۀV��
9�,�2��7��k���>'�>��>�R�>β��YX9����YIӾ��x���ͽ	!v>Wc?T�K?#|n?�$ ���0�'~"��Y6�F���sB>H�>�>��Y����`�&���=���r�����G��w�
���x=xG3?��>���>-��?�?��Y���� w���1���j<"	�>�-i?
��>i��>Z~ʽx��L��>��l?���>��>p���>]!��{���ʽ�)�>B�>ƶ�>��o>�,��"\�*j������l9���=g�h?Z�����`�;ޅ>�R? ��:!�G<�{�>K�v�d�!�A���'���>�z?���=�;>�ž�&���{�7���=,?�?5���
"�`̖><l%?��>���>���?���> ���-��,?[EM?��E?4D?���>��l=�ݗ��麽�0���=��>�B>qS=hp=����U���2���=�<�=�3 �A���d�=u�=HV�;���<��g>Z�ݿ1�P��'޾�M�^��v��ˌ���}��y�rR��Į�-�����l� ��ͻ�i_���q�������a��s�?��?��$��}~�������&�>�7������Sা������y$Ծ�����v �*BG��&h��^`��'?�����ǿ����{۾@D ?p�?7Ty?TW��{"��-8�� >�l�<X���}�뾓���o�ο1]����^?s��>P𾒁����>��>`�[>�3r>*B��b�����<J�?�a-?j��>os��kɿ�.��;��<���?��@�H?��A���=e�>�?���=N���5!��������>��?�r?�S�=F�[�
���5[?BA;��U�.<tO�=3k�=��=c�k��hd>���>No1��U�q���!=�7>Ղ���F��W�p�>�=/�>H(�]=��3Մ?{\�[f�r�/��T��;U>��T?�*�>�;�=��,?G7H�U}Ͽ�\��*a?�0�?���?1�(?ۿ�ٚ>|�ܾt�M?sD6?���>�d&��t����=D7ἤ�����㾽&V����=,��>,�>h�,�ϋ���O��I�����=���ο�{-��m'��=�+ �U�ߺ���=�I
��ྲྀ����̽�1����4�^�>[�Y=
o=���>��[>�XI?� _?�e>ȹ@>&<�h���y����ݽ�"���[V�Ⓘ
##�J�L���׾�Jž������D��Ҿ�mF��l#��cY�5s���WϾ<�O�2�(��F?x_�<v���1���~<Nx��
���="L����B[�͠L�]��?b.?��}�64r����u>�Y���E?Q�������K�{��\=�#n��=A]�>���<qWӾ"\J�}�S���2?J?K��#�����1>~OսH�<տ(?�?�׮<"ȭ>8"?lx,��'ܽ�;X>٦F>Eɧ>K,�>kk >�Ϊ��۽ �?D(Q?#m'�����K�>U���=x��'=���=�+�Dw/���u>���<�+��{���^��ɜ=��R?��>��'�h�D��6�Ľ��f<<.v?��
?��>R�i?�M??���<���k�L�J"��`�=LvX?f�c?��>�_�t�ݾ\E����.?w�f?9zI>�z]����s�,�1���~
?|�f?(�?l�<�%|��)��l�
�o�-?��v?�r^�os�����)�V�=�>�[�>���>��9��k�>�>?�#��G������|Y4�!Þ?��@���?��;<�����=�;?W\�>!�O��>ƾ/{������єq=�"�>񌧾|ev����R,�h�8?۠�?~��>
������� >*���M�?~�?��о�0�=�;��s�z�ž��g��>�ge=.����;�G?�y7����w!P�)�;��l>�b@�>xj�>ߟ<�8ܿl�¿�ڡ���<��� �T�?Sj?=�'>�%���I2���[��u*�0P�����>�&>`�������S�w���A��J1���>�M����>l@�s ��>��c��;�/�>	�>���>�֍�3[���?o���=�Ϳ������-h[?���?kJ�?�L?hY;e#f��y�H _A?��t?��P?�1e���q��ׄ��-h?g
���^�ge2�n�@���M>:�0?�?�>�b+�1�!=k> L�>��'>~+��ÿ�X��L���u�?�t�?�龶��>�ڜ?�E,?������J��+)����<�zG?�^7>�%ľ�P$�  >�UT���-?��7?}�%��V�_?�a��p�B�-�T�ƽ�ۡ>��0��f\��K��v��kXe�����@y����?>^�?g�?'��� #��6%?�>�����8Ǿ��<Ѐ�>)�>�*N>H_�f�u>����:��h	>���?�~�?Mj?��������U>��}?��>E�?�p�=�\�>J�=��AJ-�3Y#> �=��>���?��M?xG�>�9�=� 9��/�iYF�BIR��%���C��>f�a?��L?�Vb>&��=2�F!�̄ͽ�V1���輒O@��,���߽f%5>��=>>��D��Ӿ��?�o��ؿ�i��n'�%54?߸�>g�?���o�t����#<_?�{�>t6��+���%��BC�B��?kG�?��?��׾AG̼e>'�>�G�>ս���o���%�7>��B?� ��D��~�o�K�>���?�@uծ?+i��	?���P��Fa~����7����=��7?�0��z>���>�=�nv�ٻ��@�s����>�B�?�{�?���>�l?��o�J�B���1=KM�>̜k?�s?Xo���W�B>��?������L��f?�
@zu@M�^?.W^ۿ<k������7���r!�)_n;�'�>��<��F>C��<77�� E�;���b>y��>�ٛ>�.�=|�b>�2�>5V��Q�'�~�������k��y	�3����o���ƾ�y������o��I���o���<V�ʽ��ƾ ����r�β�=��U?�R?}p?E� ?2�x�Z�>����X3=�z#��Ä=�&�>|d2?�L?��*?vՓ=�����d�)`��\A��
Ǉ�1��>l|I>&}�>^C�>��>MD9��I>9C?>Ԍ�>�>-}'=��麶h=��N>�K�>M��>p|�>]	k=T��<�5��6-���;��둽���B@�?8J��We�����iȾTz���%�Qo?��>�:��
�׿S���'�E?1[$���jc���`I=�
?x?�;>���J>�/b�>G����j���>R�=��:
$�N��<5��>��6>���>NQ<�L�<��@�'�p���I�>�Κ�dR��$8����w�����
�=�B�=S_�W�/�ɭ�B%�����x�b>��z?���>� о�=���=�U4��L>� ?�p,�]��
�>�~��U�^Ƀ��Թ>�B�=^��=� ?�|H>S!�=NA�>�k��4���>��U>�F�>Z�>?�1!?������V��l���!9��a�>m"�>C�>Ӹ>��0�Q��=�p�>>,B>#��� Ũ����*D�\�V>�(�]�>����`0�<�N��B�!>[��=V��>2:�rH�<�~?���(䈿��e���lD?Q+?j �=��F<��"�D ���H��G�?q�@m�?��	��V�A�?�@�?��P��=}�>	׫>�ξ�L��?��Ž1Ǣ�ʔ	�0)#�iS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>���j��%����s��5=6v�>*�G?R��8Y�mq=��
?*?8��>����ȿzv����>/�?,X�?�Om�K㚿C�?�4��>���?�WY?�^e>�ܾ��\�Ȭ�>�??�VQ? ��>�����&��?ɶ?��?w�G>�f�?�fs?���>;�j`/���[�����y=��;lr�>X�>�Q��W�F�����l	��|j��4�|[_>�A%=��>�I�N�����=7������� Ia��ζ>�or>~	J>��>�?���>�.�>��=Յ��2��w�����K?~��?��k2n�@�<͝�=�^�M&?�H4?�L[���ϾYӨ>b�\?���?�[?�a�>;��>��7迿�}��L��<A�K>2�>mG�>$��aIK>O�Ծ�8D�3p�>�Η>����>ھ�.������@�>Ae!?��>�ʮ=
_ ?t�#?�Ei>��>CE�G����(F�}��>���>f?��~?��?����	3�i����x����Z��P>[�x?J~?gӕ>���w���{T�$�>������c�?yf?�|��?̈?f�>?m*A?��i>U��aپ������>��!?�d���A��*&�V����?2�?���>����[�׽�Yͼ�e������?�_[?�&?�n��`���þ���<�; �\.����;`�u���>3G>Ē��@��=�>6ȩ=��n�8j6��;�<��=k7�>���=k�8�����4=,?�G�?ۃ�N�=\�r�!xD�t�>�IL>�����^?Il=���{�����x��nU�
�?���?Nk�?E��$�h��$=?�?\	?"�>�J��}޾'��LQw��~x�Yw��>���>c�l�y�@���֙���F���ŽwY"��
�>��>+�?g+�>�0E>5}�>��˾�Q!��6ξ�6��� e��)�sB���7�$�(�08���T�soн�Ͼon���p>�<Ә�>N�?�`�>f�>�
�>�&�<qۇ>���="YV>ܭ>۽�>}��>�8 >�=�F���IQ?j�����'�؏��M�� �A?�*b?�e�>"�q�9L��;��x!?��?yU�?�p>��i�k+���?�B�>T�V�
?�+M=Y
����k<�Y�����9����˼�m�>�x׽��9���K�W�f�]?lo?R	��R̾=hѽ����@o=�J�?��(?F�)���Q�t�o���W��S�Q��(4h�r����$�g�p��돿�Z��	#����(�+*=��*?��?��1����""k�k?�kf>���>�,�>��>sI>)�	���1��]��C'�z���+K�>OV{?k�>$@?�;C?��X?��C?X]�>�:�>�ƾ�D�?8��= 9�>>��>�3?"�?^9?�% ?�1?�2�>S��!��ܾ	�?��?Ϸ?���>�?w+w�B�$�~�ֽ�z'�+�&�7`�� >�=1Xh���Խ֔o=q�L>B+�>AZ�C.�����OO�>&xU?��>���>J���9���=��8?��A??��>���Gn�f �ٿ�>N!I?m�<��6="��=�FB>.����k�_�%>:?>o�%>4̏��@���W>�ʒ>^>>(������A=�a#>ӄ�=5�>�T ?)�>�>�����H��9���=JMq>�W>��>8�Ծ�ɕ��G�e�=�>�"�?-4�?qg=ף�=�}�=l���f�ľ�	��l����<Zp?�?hQ?w�?�8?�* ?��>����ߑ�ï��ʒ��!�?��/?B*�>��;�������5.�0�?T��>8�U��P�:J�L>ᾴ��5V�=}�E��7��虿�L��<;�L� ��(u����?@Ӟ?~�d>vB&���Ӿ�e��L�����*?�6? ��>�7�>O|=���e�Z,��P�=j?�SX?���>�'�?88�?۸p?�P�=��?�>ם�0.���H��[,�>��x?_[?�-�?�|�?��%?�}�>le�|����-��cŻ4鍽0,����>��>FX>O�d>K�>UQ?>�s�=�������q�ͽ�:>�q�>��>f+?`?�j�>�nG?y��>�mɾտ	��ו�";���.Ž�t?��?��'?[��=��{>��� �Ѯ�>C2�?��?�%?��g��>OY�iF���q`�ϵ�>���>9
�>���=�隼̦�=���>�d�>6;*�?�h�7��4N�p'?��5?���<T�ο8�u��k��c:y���<����諭�硼vI���`��y��ӱp�䉾!L��[߽
K���Ҿ�䒾�K�~�>b��=$I>�K�=���=4=w=?~k:t��=5�����+n����?=A��<�E;=\y&��Ȃ=o%y=���J���˾�h}?�I?�_+?*�C?�^y>ʐ>ߴ6�K�>�a��z"?�U>��P��μ��<����1��{�ؾϏ׾{�c�@�����>0nH��>�3>&��='ǈ<���=��u=�+�=NVF�u�=(��=@m�=�ѭ=�I�=��>�\>�6w?ݚ�����F4Q�MY罻�:?�6�>�|�=)�ƾ�@?1�>>>2������Ga��,?���?oT�?��?�wi�Xd�>���4ߎ��p�=\Ŝ��<2>��=h�2����>o�J>"��3K��偳��4�?_�@�??�ዿȢϿ�a/>�7�>/�E>^��	�p��;6��/�ξL9?�-@���Ӿ[�>��^>�ܾ|�ھR���l�=K��=#x�ml��>0��ʼlO=3�>!��>��=���l@ʹ�s����=M�|>؀Ͻ�>�1���>���<J| >?8��s�?V�"?9x>?m??�?*�.�d�s��+۾�	�>΢�>h��>p:>L��>�,�>��&?�,#?��a?���>��>*`�>�^>��T����,ɾ1�o�yѽ��?7�?��>���=����f��5PM�љ���E?(M?�)�>%k<=b����]P&�E..��|����}�g(=d�o�"�P�a���}���߽�n�=ؕ�>42�>5>�>�v>�:>�O>��>}�>_��<ί�=�x=�x�<���̏�=,���{�<�\����9ɩ��*������a;���;�@<�p�;:��=���>iH>�C�>ǉ�=緳��:1>������L��{�=�e���(B���c�`~�"0���:���A>W�U>|���6���#?��Y>�F>��?�Wu?��$>���m�Ծ�����_��wU���=bg>��:��<;�/_�5L�=�Ͼ�T�>���>���>I�k>΅���0�h�>j�	�|�8�E��>]t��O�Z� ��t�f櫿\��E�S��LW�J�?�ۉ�e<�3�i?��l?KJ�?{$�>�8�=!�ϾF�,>����h##>���o���.߽1G?V/?��>ܷ���M��G̾����߷>�=I�d�O�T�����0�z���ͷ�ߎ�>������о�$3��g������L�B��Hr���>�O?��?�Bb��W��SO�N������s?�}g?��>�I?>?�<���z�Co���=A�n?ʲ�?�<�?
>���=Tĳ�)��>L�?Ś�?�?K�?P5[��U�>:�=�)�=�B���6�=%��=e�G=91j=.�?� ?[ ?�ѽwB��5�����s�\�|f^=��	>���>O=�>��m>?��<dr��e��=L5�>z!�>��>XZZ>��>?b�>�X��YC�p)%?�(c>�0�=��$?/l�>V�<,-�=�=�oK<5����Ǿ�9~���>J�=�,=jp�(��>r�¿|�?�>dt �'+?�:������b�>��<K�Y=��>��<�>�ý=��x>��M==��>��g>���=���_@���*��^(���پj��>5Y˾��m�m������|u������t�۾�<k�{OY�._1��짼)7z?Ԣ\��pz�!�=��5B>BP?Z�>��?���G�6�	<N��>�V>��������E����վ�y�?���?t;c>�>�W?�?L�1�w3�vZ�Ǯu��'A��e��`�U፿朁��
�����_?+�x?EyA?�R�<:z>>��?��%�eӏ�I)�>�/�';��><=�+�>r)����`���Ӿպþ�7��IF>��o?
%�?TY?�TV��Ud�W�'>��:?T�1?[]t?)�1?�;?�y���$?a�6><�?n�
?�b5?��.?]�
?��2>��=��G�;�0=ĵ����N�ӽ^�ν��2,3=w{=.L�:�d<�=�:�<��J$Ѽ�;񟞼O��<��<=+2�=���=�}�>;�N?�C?`�>vy"?�+��z�m�վw�Q?���>�c���遾��F�s�e��>���?�a�?�WT?���>�������)>l�>6=U�j>��?�6ӽ�hq����ɸ�=E<V>��=���6񜽩��F���"m�L��>Z��>ۏ>|��c%>\�����z�Ċe>��R��麾$Q�,UH���1��[v��H�>�xJ?^�?���==꾠_��2#f��(?J=?*NM?�1�?Γ=K۾�F:���J�'���>��<�d�G�������֒:���1:tu>l������7yq>��"�0$m��E����|��=��#�$<��yt辅���Sܴ=�&>��ľk�%�C�����J?�/C=�t���D�AK��^�">�ɗ>���>��ν���]qF��᧾�|�=��>��;>&�	�o��>�L�?����>ZG?�:r?Ʊ�?�H���Lu�G4(���#�E)޾���<U2?,/�>��?��>�K>'�����wv`�'E4����>χ�>�@���1.���V�s���!F�A=�=?F�>U�4>�Q?�*q?-?R�d?ȊN?���>�+V>������{<!?	�?r�U= ��y[_��A=�%=G��m�>+�,?|�O�^؅>Vr??�?�"?��G?�?^L>�����D�?ܙ>��>��W��ԭ�jF>tjN?ڃ�>}�Z?04?/�>so'�~[���0��e�=
>X)?9U$?��%?��>W~�>�3ʾۊ�>�#?��#?	 �?�y?�/��1��>f��>C2?��!=��>r�	?Jp�>)E?�(q?�%E?��?(k+=���1ӽW�N����=���<F�9=���=���K��v��F� ����:̼V���	�<պ�����<��>b>�>R*��#�#>���u���-eh=<���>���%@���X>ǲ>��|>(%>�
��M�1> 5 ?|�>��y�?�7-?��@?֧��g򁿸���]����
?�zR?�t�=�r��"��h�~���#=��v?Q�o?��h��侁�b?P�]?a�*=�H�þ��b�\��A�O?��
?��G�v޳>�~?��q?a��>��e��.n����K@b��j��=Zu�>�_��d��$�>ޞ7?�L�>��b>h��=#�۾l�w��g��g?B�?9 �?���?|"*>��n�5�s+�*ړ��'[?��>C�����?&�;�_Ҿv���}?��{;޾�I��H>�������2����������޾�'��=�&?Qv?IZn?kL]?t����kc�j�W��"|�d�V��������?���A��qB�)p�h@�(��������lS<�g{�˻B�rش?o�)?��/���>6�������Ⱦ�B>6���g���7�=����=^҆=�9\��(*�x֤���?OM�>���>!�;?HT���>���/��7�@�����1>���>s��>���>�	�::�)���彖�Ⱦ���g��7v>jsc?7�K?~�n?��v(1��n����!�;�0�~(��b�B>NF>6��>��W�O���(&��F>���r��������S�	��~="�2?gA�>~�>W�?r�?v	��s��BZx���1����<��>�i?2�>��>��Ͻ�� ����>��l?���>&�>����+Z!�}�{��ʽ&�>S�>���>��o>5�,��#\��j��y���9��s�=۩h?���S�`����>>R?Z�:_�G<|�>�v���!�����'�I�>�{?0��=a�;>=~ž=%�G�{��6��"N)?<E?Qᒾ>�*��~>�'"?��>�&�>�.�?\$�>�aþM�B��?�^?<J?RA?�I�>��=�䱽<*Ƚ��&���,=;��>�Z>H?m=҉�=���l\���I�D=�X�=��μ'W���<T���J<x�<��3>9ݿNU���ž?����Ҿ�J����?[Խ4�S����[��(p���Ύ���>�P����iQ���������GM����?u�?��x�����!ח��*w�������>e8a����l����b��̤��R�ž� &�*EP�up�8Tn�W"G?E������������,�+?
T&?Z�t?�E�����9�q�����4�P��=�'�>E����ȿ�􆾍#T?@K�>�zܾ���;፿=r��>���=E��>m�W�����%>��>��?�<?=n��}�п�5���	>�^�?97@@;?� ������QS��0??���=�N�Jg!���־;A�>���?�݈?�E�<$�V�ۊ��fbd?���=�+C��ZV;'ʫ=��_=,K=܎��[�o>�2�>�N&���<��'ܽ�.>�f�>hOH�ɍƽ>}Y�8E���c>ލ����5Մ?+{\��f���/��T��U>��T?�*�>Q:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?$�(?:ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=v6�艤�y���&V�y��=X��>f�>,������O��I��X��=����S� c�'���Fh>x��r_�����Y<��<��Ծ�]�ij���=��u>9a�>t��>e��>��>�I?4�m?Ja�>�e�>�\@�,�������Vyr���2�fx[��b�8����ݾ����>���#�I�@�sG2��%�����]>����}�
~0��9e�(fe���?;6?�ލ��O��?��C������Q�S=��>�R����B<b��T�?�??ʠ�f�d����� �=X`N��7�?��|��ho�1��j�o=�G�>T�=���>K�Ľް����Q�f�'�+?|�?����z⁾��D>)� ��H<X&?V?�5�<O�>i,!?V
 �͠-�� =>d$>>�>ě�>���=nW��A�W"?�O?=d�E���u�>�~��0�2��#�=�>�d�e���5>���:�X�7�R<�๽ ��=MLM?պ�>�.����a�:�$�?=�-��T#u?ї�>�+)>��c?�kN?(M�=����R�d��9>��b?-g??��>�pٽܾ>_��d�H?��n?&G>1�B������R*�,�̾$*6?�e?(!?��F�򏃿O�y��gƾ�Y:?��v?�n^�eq��j����V�:�>�U�>���>��9�gj�>��>?�#��E��N���	Y4���?0�@K��?��;<J@����=r=?�Z�>�O��Aƾ�f������m�q=[*�>І��gv����>Y,�ل8?���?�>a�������>��	.�?�ݑ?-�f�=�|��������Q�=�;>�����#����5�D(w�i�Ⱦߋ����=E�n>z�@S��=Ɲ?L�7=���&�տA?��2����yB?N(?��>Y�1�
������S�+hU�6��6p�>ڔ\>R�%���x��6�g]���>���=��L>�h�v븾B���J����>=��>'�t>bv��1оV��?Uo��ѿ�Y���B��b?dǗ?�O�?��>$�,�wR'���:��{	=��%?��i?��O?l-���ܑ��o"�1hr?�G��w�J���?�x�:�
&>�D?�"�>X�*�M/ >|N9b��>�Ȍ=���vѿ����L��);�?��?ۗ����>y�?��4?2KϾ!I��.�¾:=��6�<��B?��j>$���9�^a5���i�3�>+�1?�������^�_?)�a�N�p���-���ƽ�ۡ>��0��e\�*N�����Xe����@y����?M^�?h�?ߵ�� #�e6%?�>d����8Ǿ��<���>�(�>*N>\H_���u>����:�i	>���?�~�?Oj?���� ����U>
�}?�#�>��?Tc�=3X�>��=�()-��c#>��=��>���?i�M?�I�>�<�=c�8��/�~XF��DR�2#���C�/�>��a?��L?	Ob>� ����1��	!�Ymͽ�T1�^��_]@���,��߽K"5>��=>m#>��D��Ӿ��?�o� �ؿ�i��pm'�64?���>��?M��{�t�j���;_?e{�>7��+���%��TB�X��?=G�?��?�׾x?̼2>j�>GH�>��Խ����8�����7>��B?� ��D����o�F�>���?�@zծ?ai��	?���P��Sa~����7�W��=��7?�0��z>���>��=�nv�޻��W�s����>�B�?�{�?��>�l?��o�L�B���1=5M�>ʜk?�s?�Po���v�B>��?$������L��f?�
@~u@^�^?'��޿`ϲ��Z���đ�k��=6Y=Q�n>��m��$�=���=�w��!}�)��>7�>&.�>p1�>ZŪ>���>�f�>�ل�e�(��㗿�����:���9�
��w��������M���m��Ͱ�*�=����k���`��<D)�ŕ= `�={�U?5mQ?�do?7� ?Ĉ�z�>w����W=�R#��A=Ѻ�>�2?b4L?��)?@�=����he��[��Yɦ��%��{,�>Y�G>�z�>	F�>��>?�9XK>Q�?>���>��>x�0=����t=��N>�n�>N��>CS�>�Wz>S�q>���,�� �Z�`�t0ԾF�?LC=�Bd��Z��$���H��V9�7E?`�"��?����������"0?xG��ī��Ґ�f>�:?[�@?.>�ئ�����r�����<�)s���%=1̉��z[�KFF;�
?�qo>��>C�J��9�H�3����Z���sF?m���ɸ��D|��RM�Y޾�*=�=�>Ɣ>lLP������A������=PJZ?�O?U-�=L9���B���
���K>�Ť>%�(=���=<�=>��<�T���!=�N>,�>���=u��>��>��>	��>\)�݆D��s�>��=��>��>?K�*?M�½����ž���>�>\�?TӚ>|�k>�&'�a�=���>D >��꼲3'��pʽ�����>�O8�I$��!6���I�S�r={9>�H5>cW��;����=�~?���'䈿��ee���lD?Y+?� �=*�F<��"�D ���H��<�?o�@m�?��	��V�:�?�@�?!��Q��=}�>�֫>�ξ-�L��?��Ž-Ǣ���	�D)#�fS�?��?V�/�]ʋ�=l��6>�^%?ܰӾ��>6N��R�����3�u��q%=֣�>m=H?�c��naP��&>�HG
?��?��3����ȿ9hv����>)��?�ޔ?��m��#���@�ʹ�>}��?-uY?D�i>r�۾�Z�1��>��@?�R?g�>�`�w(�Q?CѶ?5��?��H>���?_�s?�P�>M�u��k/��&�������<�=�1x;�j�>'�>�����fF�F̓�UF��ʏj�޹�U�a>al%=0�>MM��5���1�=]���|Z��(Pe����>C�p>�I>$3�>O� ?I��> ݙ>R�=C���򀾙ܖ�d�K?���?z+��3n�w۶<
t�=��_��q?*X4?�T~��о<�>VG\?I��?F[?���>e!�f[���ο�����bi�<�M>�U�>x�>��t�K>1�վ�C����>��>b%�� �پ�ꁾ�λHȝ>�B!?�&�>m��=4� ?��#?A�j>[�>[ME�(;��y�E�'��>���>tN?N�~?�?Mڹ�W3�M ��ס�؁[�5N>
�x?Z?"�>�����}���iL��pI�E1��k��?lg?�0�?�)�?\�??�A?�if>�q��ؾr��ӫ�>��,?�Ɏ�E�U��`!��&��8�?�c�>1?����Q�}����#�
���>��Z?�I?�%�T�i��߾�(`=Ny���������L,̻�*�=�A>�Ҽ�׫=3�E>���<fn��@ެ�FL!>34=�#>D�H�Խ���=�<,?R�G��ڃ�y�=��r��wD���>�HL>�����^?�j=���{�~���x��3
U�� �?֠�?$k�?y����h��$=?��?�?T"�>K���}޾���nPw�^}x��w�o�>Y��>y�l���ݏ�������F��*�Ž@�ս5�>�o�>v?��?��a>uf?���c�:�#�k����3�W�� '���3�Y�L�B:0���s��wE�,^�=M���蕍��-O>GFK<��=x ?�١>�>�̬>YV�=��>!T>��>�ĥ>�*>��=[��=� >!�=��Q?Gt���(����)/��b�C?�ub?�:�>�d{�}���\��<� ?�֒?���?i r>�Bi��9*��?���>b4�c�	?��G=�[���m<������/됽!����>�@�v�:���K��[p�8�	?��?o��-�̾ֽ�Ġ��Ym=H�?��(?l�)���Q�]�o�a�W���R����|h�,u����$��p�㏿SW�����נ(�/�)=#�*?��?[�����?���k�z'?��Vf>��>�F�>��>��H>��	�w�1�j�]�.'��_��*D�>:@{?R`�>$�@?xW?�l?7?��M>���>H��\�>�'>q��>S�?�iW?w4?.s6?d�?,B8?���>�����������Y�>��?x�>'D?��?�<;��M;<��=SJ�<`{Ѿ+�K�b<|�Ҽ�Y�����k��=��>)?�v���}G���x�?>�t??l>:�> ���"����>��>?�,?�R�>Ӑ��v��#ڝ��;.?�
??���D�=��[>���=Jn=Y��<b[�=-�J���<���=Q�,����E+X>�a�e��<���<��a��D>΍�>��?���>='�>>��@ ��m�g��=c*]>jU>�`>]پ�3���R���g��Gz>q��?��?h m=���=D�=�K��bڿ��Z��{��>>�<�&?�k#?dHT?T.�?5s<?�)"?}�>�z�rr��sF���
�?��5?!��>Z���Z�����a�%��d?!�?t�[�ܑ̽�4�/CǾ�����U>�J�˹���E��.7�}t�=1g�������?��?�%=��D���׾T���ox��i�@?�6�>�ϳ>YD�>��߼e�*����Z>���>Y�H?$y�>�wO?Q��?��?v��>��@���� ���Y㼾���>z?P��?}�?�I�?��*?Ә�>��q�t_�p'پ_z(���]�8����<�=��+Yi>;D�>;q�>�:>�G,=rhH��*�!��=�&�=�[�>iF�>�s
?>3�>�J�=}�<?gr�>��ξ#l�����]����ս��n?@�?���>9�<L�7W0��� �ކ�>ۿ�?\��?ϙ?����J24>�Ͻ{��=lc��@�>��?K��>[P>0��e8G=�A?��>�̩��J!��2(�e��M?��a?���=��̿xρ���(�<ǈ=��ž�f�#'̽���<����
��V���@��<8��'����X�.X������?��><(>(~(=L���Y�=0�<[�=���=���=ar�=[wZ�0؏�=��<3*�<p!=$�H>*?O��(�(v˾�}?lI?Dp+?��C?�nx>E>�Q3���>�킽R�?h�U>w�P��p����;��>��}:��پK�׾��c�Rݟ�Z>P�I�<>k3>E��=T?�<&��=�s=c�=AD<��U=�k�=B|�=��=���=��>$>�6w?D��������4Q��Y�q�:?�8�>H{�=�ƾx@?��>>�2�������b��-?w��?�T�?3�?�si��d�>���㎽Dq�=���o=2>���=�2�S��>`�J>����J������4�?��@��??�ዿŢϿ�`/>[̉>'�M>ViS�� ������Uؽቀ�:T$?�C �����Q>Ū='/�������S=Y�>o1�=t�p��Zf��m>��1�C����!�<��Z>Vş>��>�ޚ�՚��SB=� >>A�>ER߽N�Լ���}�ɽd�=�]�>.tc>'��>Oe?� 5?�Gh?R:�>y�{�#�ƾ�I̾ꕁ>]t�=5��>��=��`>v�>��8?��C?�M?��>ꒉ=@��>���>��(�h�tO�8���U>=!�?�k�?_=�>�
��.�X�4:�ˑ>��\Ͻ�??�.?�y
?*-�>H������d ���.��雽Mv;�vZ=�r���z��`Y�d�+�L2�Rm#>1F�>`��>�^�>:��>(?j>:7m>I��>r��=
=<7�=D@�<�=�V�\=l��
��<:�0�+��:

1�u=��+��X�ϼ}��<95�;{����
>�e�>h�Z>S�>�`/>�v�����>1�����W���K>D���03��Rj��u�� �
R9��>>_��={���D��X�>m+#>Y��>�L�?@��?�-�>��!�C�۾疿:me�n���F�c:�/�;>A���"�6I�m�C���¾�r�>Q"�>K޻>�s�=�S�d;T�T� >�ξ!�1�h�?M���de�1sA��B�3���`���#I������<J?���\r>q��?S?��?�w�>������)���=
���$>���C���H��WkP?[>K?)�>�9�=�`�H���1�b0�>z���	H�����`3��b	�n�>�p��>"\����;hQ��Z���聿�+�c�
��=�>�V-?j��?��L���u��rj����o��>M�K?���>�G?9] ?�j%�|�ƾw�����=4-z?3��?�p�?�'�=�$�=����V]�>�?��?���?#&z?��L�XL�>~�^=��$>q���˧=���="ñ<瑐=>�?��?Tv?�-��~9��(���쾈%��1�<jը=I�>6��>2��>�r	>�Q=�Y�=9	k>Q��>��>/<N>]S�>�ę>u�y�w<
�.,/?%�<>��<�uI?kj	?�e׽*K�"֌>i��>��<����|'���e����="�+=�O>-ު>�O�> ſ捄?1��>����&?9(�(Q��Q�>H��b1%>��>�7Q>zw�>�a�>��?n�N>[��>��E>�!ƾ؃>�f�͎!���D�L�φ;M��>]O��'�*�U������rZ��'��	����f�]�����9��_<PT�?��L�h�-T,�(C�q�?-V�>l26?0ꑾb�e���>���>��>��j������uپ���?c��?�c>�	�>��W?��?sf1�H3�TjZ�ۜu�t�@���d���`��ݍ�������
�J5��E�_?��x?ugA?	L�<�cz>i��?��%�Nꏾ �>�/�5';���<=G*�>>+��IEa���Ӿ��þ���yF>��o?+�?#B?N�V��U��/�>��Y?��S?T�G?�v.?��C?�(���?,2�>y�?��	?��I?�B?��?��:>�*U>D��=��>W/�����)�]�%�����E�>�=Ts�=4�=��:r����ս��=����K�ͼ9v�� ��=��8>⚛>;�R?�(�>u҆>��9?ne"�dh0�p��"�:?���=��U�=F������h���9p=(c?��?�cW?9u>uM��DG���2>��P>'')>�#>ME�>m���[���>U�!>9(�=��P<�1�wr����@5�������g>�4�>�2>M���g+%>�X����{�M&f>�xQ������(S�ČG�\�1��
z���>K?Z?���=sh��Ϙ�U1f�we(?'<?+,N?��?��=�׾�::��RJ��:��R�>�ו<��[<���-���9�$|,;.�r>�d��Xx�5mq>f�	��-��ha�}N�����D��=u���?�b��ǾɆ��x�=�>F���-�s՘�����J?�Kh;/�ʾ#|N�B���3h%>%�>&��>*,ͽKĽAM7��|�8D{=�ҕ>�o>Y>�G�C�����x�>��E?o[Y?�F}?̴��j�v�ș9��ً�~���?��>�I
?	R->���=�����'��l�Q���8���>}�>��X;��˾#���(���>�?��=^��>6�4?Y?�7T?<C?�?��7>�Z��ݾG]&?W��?.�=�ֽ�����@���>�Yk�>�J%?'O���>�>?�"?bu?�uR?�w?��>ϓ�,=����>��w>��P�枨���>��??Ю�>TV?�Bt?��2><�@{���,]��ʂ=��=>d�6?,�?���>�ǜ>��>OH��v�=�4�>l�b?�E�?�:p?'��=
�?��3>���>᳓=[ٞ>t��>��?QO?�~s?�VK?�J�>���<m*���ڵ�D h��W��8�;�S<z�o=�P[w��u�7�<6��;*ü��������C�����>F<l��>�σ>s����g#>'˾�🀾ӆ>���♾����q$�Oθ=�l�>?�>��>ޗ3��ɳ=6��>7F�>���E,?{R?�?�<�6b�}yվ�}V��D�>5?l��=��i����� \y��z=h:j?c?5bU��:�ٔb?P^?V��=��$ľ�`d�ˣ���O?�}
?m|J���>FE~?��q?Җ�>�-e���m��Ҝ�ab�mGj�G��={ܛ>�p���d�5��>|7?�F�>�+d>Z��=4�۾��w��.s?ȁ�?ү?z�?�I+>��n�'࿓�����4�_?��>���?.?�D�;���a;�����3pɾJ9��nW��D,��̢�)���{�"y�a�>��?�Dd? �n?�	`?8���&K�s4Z�^�z�]AI��A	��4�vI�~TH�(E�Np���=G���4�����=�~h��98�<k�?<|9?9)7���>��O�	�y�����W>ЊL�q������=Z�?���<���=��L�(	ӽc�t�X�?hW�>Е�>�T<?� V�A�E�]7��A������=>�%�>���>�Z�>� �;��������bɾ���f���t>��c?B�J?��m?p��� 1��q��i� ���>�0��%�C>�%>#��>�W��T��=&�O�>�1s��s�� ����	�O�=D3?�܀>�Ҝ>s�?��?v>
����}�҅1��8)<(��>0ye?���>���>�*ֽ~$�E��>�ql?h��>!͠>�勾�"!�v�z���̽���>�d�>�( ?xq>�?*�W�[�SG���6����7�5�=�Ph?�3��ː`�vք>�qQ?ثP��T<I��>�c�� ����:�*��>�{?�=�-B>�ƾ�;���{��j���6)?�+?���Y�*��~>X"?[��>!*�>"-�?�f�>^cþ�����?_? HJ?�JA?�.�>�Z =b
���ǽ**'��'-=���>�Z>�/p=���=�>�=Q\��c��G=�-�=�{Ҽ[߹�ֲ
<����o�N<k0�<�3>�ؿ�A�ң�����I6;A4�?튾�����_�ƤĽCZ޾����s���]\��o�������e�݅��lA�O/�?��?�ľ��[��fX��j�he�>�ľ�)ν���@{������}���%��6��KB��7��x p���'?������ǿ�����۾uM ?]?"�y?l���c"�Q`8��^>���<u揼���·����ο"ۚ�M0^?S��>�U��u�� ��>�>�>C�Y>Zr>?Ɔ��������<��?�;-?��>ep�0ɿVj����<�v�?^�@8�??�g�Ѿ���=�%�>#��>7P�=�]��2��E���i�>���?���?�|G��j��">�ga?�ȼ#�C���=��%�=_�=^S�=l۽Q�~>Ip>tB7��G�ę=o�">�V>�#����%�U��ױ==T��>,�=�F�<8Մ?mz\��f���/�U��U>��T?+�>l8�=��,?�7H� }Ͽ��\�]*a?�0�?���?I�(?ۿ��ؚ>^�ܾg�M?�D6?L��>�d&���t����=41��A�����]'V����=���>R�>΀,����e�O�>����=���	>ȿ` ��������<{`N��6�����->/�>n���b�g�?����=n�1>c>��>�<�>l��>x�U?L7�?��>W�>i%��='���,���c=a0�;����޾�$��Q�c�R��3n߾�!���(��2,�N��Y�!�j��=�7��w��/���UV���K��?H�;�B���j�b(ý����yB����˺hB��8�ľG)S��jT���?� ?ϧ���7y�5о�~�<w�5���W?�Dk�����֙��<>�W����>�1$>K��>%횾�=�,}�4�1?qN?�Թ�WC����>� �%"=t�(?�P�>>��<>�>�u&?~&�����%�K>T2O> ��>���>}� >p櫾��½�?rkI?B��|֚�V��>�K��� a��ɡ=���=#�N�A���Dm>��=� ���� �lI���=)W?���>��)����,�������b?=Sx?�?y՟>�.k?(C?�թ<<�����S��<
���w=VW?�h?ʞ>%}����Ͼ����65?He?��N>lg�=�辛.�����a?�-n?��?���֮}��!��pV��V6?��v?Rr^�2s��A����V�k=�>�Z�>H��>��9�Jk�>�>?�
#�0G�����Z4��?��@B��?��;<d$����=�;?�[�>�O�V?ƾ�x�������q=�!�>���ev�����S,���8?Ƞ�?���>p���^����='����7�?��?�k��6B(=nTѾ����"����|�=�r\>���=z�`=y���]G*�	���V+���N�椧=?��>j�@7%����>��������ο���I��������?�/?%��<+U����H�%a�2$:��-A�p�ʾr�>8�#>��񴌾�,}���=���׼ӫ�>���)zb>��@�����Pю����f�>K�>?E�>�ֽ�s����?���YɿK�����xP?/��?]΄?V�?�~;�<��xHx�j�F�<?K�q?n/[?Y|u����d��Ķj??��~F`�*u4��0E�*<U>��2?�!�>��-�r}=4;>���>�>E*/�.�Ŀ̶�yw��D�?�t�?�r���>ƀ�?!l+?�n��3��VS����*��g��w A?G&2>1���M�!��C=�Mْ�o�
?�0?�r���e�_?��a�)�p���-���ƽ�ۡ>��0��e\��P������Xe�����@y����?.^�?d�?2��� #�N6%?��>,���~8Ǿ} �<^��>�(�>�)N>QG_��u>l��:��g	>��?�~�?^j?�������AV>��}?8��>���?@��=�	�>��=�H��w��#fP>܃>�$��'?�B?yV�>ͷ�=�?����4�Y
J���N�����E��?�>��n?��J?�Ն>=Z��� e���,�@��-%;�q���u�U�GJp����&>z|P>��>��M��JҾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ra~����7�K��=��7?�0��z>���>��=�nv�߻��[�s����>�B�?�{�?��>�l?��o�J�B�g�1=8M�>ɜk?�s?1Qo���\�B>��?������L��f?
�
@~u@a�^?(������ɵ��_���������<tZ�>�⽙��=�^@>�v#=�ƻ�/>ĳ�>�U�>Gν>,��=Y^�>��>L؁��3%�C6��}���(�c�G�#�w�ž�A}�H}�`qs��jʾ�!����|�,>���=N�-=,�>��i*�$:=#��=_�U?�R?;p?/� ?2�x���>����S5=0{#�G��=�/�>Mh2?)�L?�*?�ؓ=�����d��_���B���ȇ� ��>�uI>w��>J�>g'�>��=9��I>�2?>"��>�� >W'=4���]=>�N>P�>���>3{�>�q>�I�=��}樿�&�rXK�p���k�?�볾c)E��K���g�������=�`?c<2F���B��x����6?�$y��< �Y�����=�<?5�?��>s
��|>�<�>�X�i� �>�g.=79��&�<!�>%%?��>��>��'�ҹB�|�p���{��f@>�I?:����k/��|���5�D����?V>T�>}����#=��|��F�y����{K>ml\?`�~>-���u��x�V����(&�>��>zy��NO����9>��=�\^.=֮�� �N�rC>eaM>��?�d>� �=�x�>iM��jm�=>^/>�ʆ=��?x�!?纠=�F%=�8���T���>���>m�>k��=1�;�b	>Z�>^��=u�
x	�t���
����^�>&0�c���P9�'ͼ��}d>�Ƽ�����m	�=�~?���(䈿��e���lD?R+?i �=�F<��"�D ���H��F�?r�@m�?��	��V�?�?�@�?��Q��=}�>׫>�ξ�L��?��Ž5Ǣ�ɔ	�/)#�iS�?��?��/�Yʋ�<l�6>�^%?��Ӿh�>�t�Z��X���u�	�#=̧�>�8H?/W��b�O��
>��u
?�?�_򾡩��[�ȿ|v����>��?���?
�m�OA��J@�r��>���?�gY?Jri>�f۾�bZ����>��@?h	R?�>�9��'��?G޶?3��?��H>���?�s?�R�>�ow�wT/��'��낌�n�|=AL3;f8�>;g>�����]F��ȓ��c��ͺj�C���b>!
&==�>0��u6��7*�=w���
��J�d�W��>d9p>�H>���>�� ?6��>�,�>�A=SU����������g�K?���?O	�ȡn��i�<齖=�aa���?�w3? �k���ξ?�>v�[?�>�?,�[?��>�l�6���ƾ������W�<�2U>'��>��>�B����H> Oؾ�SE���>��>�����nؾ�ă�}���Ւ�>�J ?��>ir�=p�?��#?��j>Dְ>�zD��⑿�6E��N�>�1�>2Y?:�}?N�?cʸ�y3��_��X����Y��_J>��w?��?�>�4��+���G����^�F���i,�?�g?3�M�?Q,�?�]??<P@?�in>���
KؾA.��l�y>��&?�p˽�q�m&+��~���T?��}>(�3?
ק���Ǽܿ=/��<��׈'?�N^?c �>ϗ%��P�1x��sS=S��=����D�8]����=!�{>���=F��=w|>��V>_��샦�f�=J�]>�|�=�qR>���>8=,?��G�,ۃ��=��r��wD���>�IL>9��l�^?�l=���{�h���x��.	U�� �?���?(k�?���h��$=?�?�?�!�>K���}޾���3Ow��|x��w�!�>@��>�l���Z���ۙ��\F��O�Ž��-�?�,�>���>���>�G>3Q�>�ه,�J��bM��op���&�@n7���'��e �ϡ��XKu�&w<�m���H�����>$Ͻ���>S��>:8�>aՔ>�G�>ï�O>�ˆ>��>��N>	��='fR>�CV>T�缁B�d&R?(��`�(����s���F�A?EEc?sf�>H2e�����:�Ә?�?pU�?Nnz>�i��r+��?���>���� �
?{�H=�.�c,�<θ�! �d��r 
���>��ؽ��9�q�K���g�\
?/�?�V��"�˾��ؽ�������=�΃?��&?n'�=�P� "o���T�a�S�S�U��l�1s��Z�&�+�o��펿�=��
��I�*��xA=u�*?�φ?�- ��$�21��L�h�y�:�]�o><�>n�>=T�>�fT>����k3���_��#��%w��|�>A�y?�˃>��B?C?��O?@�S?��>��>˔�����>ty�<�>���>G�#?�?(q,?�)	?��)?�-�>7���|�rp��?��'?�K(?�?�H?�+���n�;{�ս=%`=䈓�^f½��=�XظSЉ��U"���s=�l>�O?�m�̘5����,H�>��??pٔ>aE�>�?��K�b��m�=m)�>�B?D�\>E���W�$�ξ���>#�I?�T(���=�G8>��>�t�\�:H��<�MI<��=E��=�~���Ŕ��C>C�W=R�;�������W�=ʽ�=`g�>�?��>�?�>{0��ݥ �J���,�=�X>2�R>J^>�پ�p���!����g��Jy>�z�?�v�?��f=��=�x�=*s��kK��}���������<��?�F#?�HT?���?÷=?.X#?��>���I��ka�������?��+?鱢>ߌ���׾�ǧ���1�f�?t<?�T� _��p�/��¾YŽ_B>���px�j��d�<����P���������?�	�?��#=�1�%оC?��_���=?
�>ħ�>�S�>kb'��_�+��`>�j�>�YH?z �>��V?V�?�e�?�>��P����;1������{R>m�J?���?��?0�?��>�n'>��J�7þ{N�R����y���c��Y�=u�>8�>��>�y�>��9�(����& L�C�Q>㔪>�?{�>�|�>��C>�R��N�H?}�>.״�!���ž�A�����K2r?���?@m?��<����g2�`=�)�>�\�?���???��i�i.>�I{�rG��Z�J�'�>A��>�i�>=��Ka:>ٯ�>c��>��,�o��"C�G�=�?�^=?��=�ſ{/q��r�W���D|<B���r�f�=����X[�GW�=�
��u��J ���[��������Ub����}�F&�>�K�=�t�=���='�<�����<�JP=T�|<r=>q��z<`�B�M����������<A=<j>G=l�"���˾ƌ}?�:I?M�+?��C?��y>iF>��3����>����$@?�V>èP����5�;�������0�ؾ1w׾�c��˟��F>�BI�J�>�83>�O�=�4�<D7�=Ks=X=5�S�77=�0�=�J�=�h�=���=T�>�]>�6w?W�������4Q��Z罥�:?�8�>h{�=��ƾp@?{�>>�2������yb��-?���?�T�?<�?@ti��d�>J���㎽�q�=T����=2>r��=s�2�V��>��J>���K��I����4�?��@��??�ዿ΢Ͽ9a/>ށ�>�4>�0�3|����=���S���r-?m�d�Ƅ���a>�=�>ǈ��ױ�]�w��1�>Z�J>�裾b�l��h�=9xI�ò��S��=���>��>J�<�y��M�UǤ>j�>.`�>
.�����<�Rr��S�=�(�>�_?\tz<O��>��?Ǚ;?8ww?b��>@�i�lR��2��c�>T>3ֵ>�+�=���>J��>s�;?:�0?^�M?> �>��>vì>���>(���Z��f�����[q�=r��?��?�N�>�Sc����JA!���<�C�Ľo?�0?��?��>���z�Fr#��'�v<r�n���	>OC��"�;�ue>����xT���>�^?F��>[�>��>�a�>��>�T�>�a>Q�l;���=֤�=�w�</>�ږ��|����2�~��'#�<4�6=�,I�᷄����=�v�=z3=��V<V��=���>iI>���>5t�=(���K�2>�����HL����=�!��4B��Fd���}��v.�H�6�M�B>LY>T������?!�Y>�B>���?Hu?�f$>����Ӿ�q���{b�SU�k2�=�+>�=�M�:��l_��sM��bѾ&�>/a�>���>(U>;,�^�<�
�=X�ؾ:�0��;�>���)F��\���k��5���A���f��<I�??���nf�=��}?��P?O��?��>�Ի���S.>N����)�=������a���K�?f/?E�?��Ծ��@��˾�J����>f�I���O�����L�0��J��9���>����\�Ѿ�.3�a��B揿��B�As��v�> �O?�ٮ?[�b��>��\�O����������?'�g?2�>��?�?�ě�_����+Ҷ=��n?=��?���?_ 
>��9=�8����+?s�B?�ԏ?�C�?VȖ?�����O?ob��HU>1�����$�0@s>c�8<I	>4��>��!?�W;?^G������.��e2Ǿ��3����]�_>[�Y>/>�>�->�R�=���=xϲ>��T>��i>�W�>�$>�I>`�>�������;�5?�fe>�}�>�{P?jt�>-XI�<�=_'�=���=��=��C����=:��,��=L��=ns>���=�>s���W��?���>���i�L?ǃ4���}��>ƓS=?�=t��>�����'�=��>�-f>��=�X>	�r>�Ҿ�U>i���� �cqA���Q���Ҿ�az>\�v�,�Ɯ�m�3)P��=��_2��j�26���>�M{�<�?�� ���i�;�)���T�?uF�>:u6?����7ט���>|a�>a�>�����ŕ������ܾ�Ԋ?���?�;c>~�>V�W?�?��1��3��uZ���u�'A��e���`����0�����
��8����_?��x?tA?�Y�<6z>���?�%�;؏�"�>�/�	 ;��|<=/�>�1����`�`�Ӿ�þ�G��>F>L�o?�%�?&V?�MV�Z�m��'>�:?�1?-Tt?/�1?ݜ;?J���$?4a3>�C?�d?jD5?�.?t�
?�2>��=9q���+(=BA��5�W�ѽW�ʽ��ֺ3=�D{=%�B��Z<��=���<?��&�׼�3.;�졼�߫<��9=�Ң=8g�=sC�>�d_?W>�>a�h>j�+?��.��1%�T^���?c����L=W��������"�Q�~|S?��?�af?·;>�?s��W�UGb>N�#>��>�T�=ՠ?�7��X *�uP�;(8z>4%I>�»�1�=�v����#����(=Y��>��>��>�%��n�<ö�����S��=��нiƴ���
�+�� 8�����1�>|�X?U��>(s�Z-���:��Z�_�^C?�t?�ig?5��?}�=��~�Yk[��XU��Px�Y��>��ɽrv1��9���ۣ����3��=�%>r�M�����o>U��Hؾ�i�SJ��)侱�=���*0=������4��մ>`�>#ƾ!�L������`H?��f=�+����q������>>��>d&�>��K�@"M��<�wLʾ�ʏ=���>D{;>��N�����C������>E�H?�~?��?�u.�.����4�8�/�2����>��>�C�>�w?���>���=ɶ���5�a�O���6����>)��>g �p�2���S�龞z#��Z>s�?�!i>�?;�T?6�>�P?�-?�?u�H>��='����!?��?¸(>�*U�"�$�޲\���/����>�7?8���"�>Z�>T��>�M3?/a<?��??��=���<I�ݛ�>�]F>�j��<���E�=ȯM?��>��y?M\?��>>CLa���������x/>ㄉ>�p�>��>X?�>�>g�>����TC>s:?EX{?N�i?-m?�=�+?��>"*?;J�=��@>��?)k?J�,?bl?y�e?�d2?a�<��y0��e�L�K�u��=P��<�\s�{L�t�2��Vg=�� >w;à�;�&���ؽl��<��潎��9���>�-�>u!j���=����	���.6>]:r��������#�c�>oņ>IE�>�>���w�/>Jj�>ݼ�>���u&?�(&?5[ ?�߫<�̀����L���V<�>��^?�>l�Y��Y����e��H@> �g?��g?ԫv�,�2�J�b? �]?h��=���þǶb����^�O?6�
?�G���>��~?S�q?d��>��e�:n�!���Cb�*�j�]Ѷ=Mr�>VX�_�d�l?�>q�7?�N�>m�b>$%�=Tu۾!�w��q��Y?}�?�?���?�**>x�n�M4����9ꌿHWL?E��>��c��>��A��t��=ˢ���>1���^޾xm��_����%L���j�����/�=.S?EK?~�z?,V�?�+����1��R��Dl�.�?����Sm��B�(�9�`�9��偿(e8��v���q��^B�{�{�^�>����?qy(?xH/�i��>���@���˾�H>�*��U;��ܘ=�k��:(=�yH=¦d���0�꬯�� ?�>rX�>H�=?�JW�`=�2�Q�7�J�����.>|�>��>�@�>N�I<߻)���I�ʾ�˄�E�ͽNx>�hb?��R?:hp?>D��5���|�f�+��^�B]���2>>!>T�>v�<�%�"��1)�8���o�ٛ�y>��R�����=	�2?���>zC�>��?�3�>�9��*��2
^�y�.�#=���>��j?|{�>Uv>�n˽KF�b�>�jl?<��>Xܭ>̅��j*�TRw�,+��7I�>�(�>�G�>g>��/�y�T�eE���Ɉ�&�+�;��=*Z?BR��[�T�_�>+�[?Ԍ�<nG�PӚ>'�H�7�'��\��}$��>ht?�{>3�>�ľ2���{��j����*?�A?)A��h(�� `>`�?���>F��>ु?�R�>Kپ�@����?[�^?��G?�[6?��>�;� ���A��nw$�%=���>�2>ܠ='�=6��rP�!d+���Q=�x�=j&��I��J0A<�M���D<E��<��->�$ڿ�@W��eѾ<��H��� �$�e��K=q�ټ��$��7��'ޤ��ؗ�e?ڽ�.ܼ������sI�� v�I�?�D�?f�꽯5꽖���nタr$4�o�>���<���R����f�VoƾP�վ�!��p�A�ψb�Kވ��|t��'?ɓ����ǿ����I7ܾ! ?/( ?�y?����"�]�8�O� >J}�<�꡼������ο1���p�^?���>1�.������>q͂>�Y>]�q>������� ��<`�?w�-?��>r���ɿ�~��	�<l��?��@�>?��� ��m�Ľ�K>���>�?3>ʅ���L��ʹ�Dy�>-T�?�d?��p�P3c����>rJ? �}�U������>P+>��=P��Al��zэ>�H�ͪ3�b�O8��>�2�>O����˼��s�Sn��[N??�tK�q~?�4Մ?{\�yf���/��T��U>��T?+�>Y:�=��,?_7H�a}Ͽ
�\��*a?�0�?��?�(?Dۿ��ؚ>��ܾ��M?dD6?���>�d&��t�a��=�7�ێ��b���&V����=T��>@�>�,�؋���O��I��c��='|�@;ҿ�y�
��x�C=�k`�f=�f��G���I���0ܫ�G����.>
s>"��>���>�H�>Q�>ǁS?��z?��>�0�=����2��kw����=�/+�z���V��&��a��������֘�oM$�SC������3��P�=��0��r�X�<�\�g�x+���X?�>A.�q5����Ѿ|��$����7��������xE�a�k�Z3�?|m?�]��3@�������|��t[��!\?�D{��Q'�������>ΆW>��ս�~�>C�+>;⭾c�<�;Ka�_�-?�
"?�ٽ�$���~�> X�*�=�,!?���>\	=��>��(? 0B����W�I>2�=>��>U��>�_�=FԲ��q��	�!?�T?��ӽ�¦����>-ż���d��x�=��>tp@�Q%���sl>/�~=�*�����'�^�gF��J?U��>�T2�lJ ��|�Ӹ�=��=7�u?�Xt>��>�HR?�PH? �>0!�/'S��5
�A��=r�\?qW?܇>-.��?���T����>?���?�>�-��j��a�(�?��M�?>ُ?�&?�mu�5Z�g���v����q?8�v?�h^��m�����?�V�(/�>U�>մ�>��9�i{�>ԑ>?5�"��E��A����X4����?q�@Y��?��;<�:�(��=(D?ul�>e�O��OƾT�������� r=�+�>����cv����A,���8?���?��>Ϛ�����#��=�Е��Z�?��?���٬e<q���l�h��}��<�ӫ=���V"����}�7��ƾ�
�����/E�����>�W@>@��3�>�38��3⿪QϿ���
bо1fq�	�?+~�>yȽ䋣��j�lNu�)�G�S�H������2�>�w>&G��pf��m�z�`;�x������>��w��>�Q�B"���䟾L�:<FG�>��>D�>̓������3t�?\h���ο�k��Q~�aOY?���?=Ʌ?W�?/��;|�|��%���<��F?�s?f9Y?��$���]��Q<�`"[?�/e���F�-A7��1���>��!?Pi�>�;,�kb=�s!>	��>�ɩ>�7�'�Ŀ�袿�о7-�?��?��۾X�?�H�?%�?x> �!����������l>0f?�?>���E��8L�J'�h�?<�J?x��1�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?	8�>{
�?|��=���>E��=ٱ�	�"��L>�0�=� 7���?|rM?'��>�o�=2�9��4/�4�E�G.R�2>���C��U�>�"b?��L?дe>���Ӊ;�zc!���νԃ0��kҼ�B?�o:(�gٽG�6>��:>��>vD�l�Ѿ��?0p�$�ؿ�i��p'��54?-��>�?$����t�����;_?�z�>�6�,���%���B�X��?�G�?(�?X�׾nO̼�>��>tI�>u�Խ����򁇾e�7>�B?C��D��~�o���>���?�@�ծ?`i��	?���P��Ga~����7�I��=��7?m0���z>���>W�=�nv�⻪�U�s����>�B�?�{�?���>�l?b�o���B���1=CM�>b�k?�s?6o���:�B>��?������K��f?��
@ru@(�^?C	��:쮿����� ���~>W�>�N>Rl����0>���<�����=mZN>}�>�&?�Q?Vs>�Y�>�uM>���C.�w&���,��haD�{F�6�վ`��3�Ծ��վ��z"�U.\�ɜ�=\[p=��<�sK������"<�*��=��T?o;\?�1q?��>s�Խ�'>K5��)<�B���<�>��+??>M?��!?��V<�ʙ�@Xb��^}�����=��A��>ǵS>���>T��>�͐>�����GB>��H>j�>��=�j=�9x=���=��>G>��>�y�>�j�>a�>>G���cC��1Zk�vF�G� �R��?h�$��挿T�q���Dڻ���м�A�>*}i�k맿����?K��NkK?����1�$��.�>f~M?��U?�^v�5xվ��>,�>�=�(����G�=<"�=2����6��Ǻ>D<?���>č�>����p%�\�[�ᩐ�d��>l*'?xx�����P����n�]Qݾ�y=>w��>�FJ<�t����J*~�Q�G�St�=Y2?-@?�R�]h���;�I��&�k=zSQ>y3����="�5>�&A��@l��߽��=r�=tA0>�m ?�Iv>|��=A�>Z������&��>���=�z7>H�M?e+?i��<���s��.�<��Ʉ>_�?ڻa>ˈ=�n]�һ�=�?�չ>&=�p)�c�F� /c�<Z>��׼�84�!�ӽ#Y%�}V�<P�8> DG=����_[�$�ӽ�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ'��>T��j���[�����i�A�={ �>o'H?��	��7D�6(�(�?�R?��]̠���¿�#c�I��>��?d$�?��o�����:��,?�h�?�\?%��>��龆�o���>�XC?��n?UX�>�*��/*����>�x�?���?[�I>P�?��u?�G�>FP_�Rg2�W"������|l=-B<�]�>E,>�!����?�����������e����U>�"=�>��轨���ϯ�=A�����Y�Ϡ�>o�b>
7E>��>��?\��>�>�c	=\;���~�����L?{��?����jm�4\�<4��=^]�9?.�3?�tY�C�Ҿ5�>~�Z?�?�Z?���>}����𝿿<���<˓<��K>���>�;�>b����{N>�RԾ'�D���>�O�>cq��qپl�}���پ�>`� ?>�>�F�=�� ?��#?J�j>�'�>�`E�i9����E����>���>�H?��~?��?�ҹ�][3�����桿��[�=N>�x?�U?wȕ>n��������@E��/I�N�E��?Jsg?�V��?32�?Q�??%�A?�#f>��qؾ������>��2?Z<^���Z�i�<�����>d�L>���>Y�W������}�;'������8>�RS?t?�p\�xg��n�*�=�Ⱥ���=�2�=E�B�<a�=�P�>l"�\q$����=�]=|��빽��e��1�<Q(?m�:>�}���[��G+?�8A��k{��f�=ۊp�ִE�`�x>u�?>?����a?�45��y�����ZN��U��:�?�>�?]D�?yp���g��q;?�È?�B?N��>t,��m�߾q�߾��v��jy��/�g��=�%�>a3�:إ��Ң������j����_��f"�>��>�?1?&;>5E�>����V%����u��}�X�H �as2�5L,�w7��휾��'��w&��þ��~���>��v��
�>9J?�ER>�qi>���>���>��D>ͬ�>��>��h>�>"
�=r; <���FR?����K�'����I����@B?�ed?�!�>�j��������ǀ?ӏ�?�i�?��u>Luh��#+��r?E]�>���0p
?� ;=<�ఈ<�`��3��jC����e��>S׽�$:��M���f��b
?&?�o��px̾L6׽;���u<���?gM,?�+��M�Rvq�D�H���;����d������),�!Ze�+Y��ܻ������R(�Շ�<=�-?�ʈ?���ڗ�������\��mS��5x>���>��>6�>q��=������-(K�.i"��P���g�>�e?OÑ>��>?Z=?��X?RJQ?v�>�ܩ>:����*�>k�R=%��>���>�I,?1)?&'?�??�B,?N�{>Q4�������,Ѿ�8?�$?��?��?ef�>m磾D�hẽ~?�%L�x��I�=�y�����&���:�<Ӿ>O?�*��6�Q�1�`"�>���?�d�>�>�DA��ܾ&�=Gh#?�?�ϒ>zkv��`<����?�%�?�YU��s=�>,��=��F��=E��{�<�EU�kt�=z���sU�|S�f�y���=-?'���<��X�L��t�=Fr�>�?䙊>!C�>�=���� ����?�=\Y>�;S>�>5@پx|���#����g��^y>Ow�?�v�?�lf= �=���=o��q6����N���G��<�?�@#?�KT?��?��=?�m#?��>�,�K���]�������?��,?:��>"�˾pꚾ�(��_�2�!�?�Y�>EZV�҂��PK��ƾZQ��+�=�H/��yl�?A��'yG�H���=�������2�?2��?�,>��@��S���,���ڲ�� B?}��>O��>Oz�>/�xXb�6�%��/3>#��>A�D?��>�0F?���?6ss?�IN>��]��Q���c��U�/;9�>��=?Z�{?ۙx?j��?�c�>H���ͽ�l���˾Ȧ��,@9�Hʫ���>�2�>�х>��>�Z�>8�=�0w�9X>a����+�<�e>�e�> ��>B��>\ �>?h%>��D?W��>ܗ��sr��R慾Q�s�/0r?dt�?��+?`�6=���B�S��z��>�ɢ?���?��&?�ah�ܩ�=��x�?���j��e�>��>İ�>��=/=�>�;�>"��>,��D?�ݖ@������?tP?t�>�zĿ�Rr���D�@�X��t����5}{�?�0��f�����;>5��:�Y��ixm�$��� h�������m��?�u�z�>6}=���=
�=��=��=;�C�_,-=U����X����*����a�E��<`'ֽ�����������<�3��˾}}?M^I?#,?�D?�y>Y>Q%6�ko�>{�����?%kU>��T�c���;�����x���ؾ=׾�qc�k���$�>�J��)>H3>���=���<�L�=��o=�i�=�җ���=���=�3�="��=��=j�>��>�6w?X�������4Q��Z罥�:?�8�>d{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ5a/>J�>�'�>meW�� :��뫾�eq����P��>H�L�ok~��l�>zjE>� ��&�t_>t>�HK=ܳ��k�z�)=b�P��)>�km=��e>+�>`0=PO=�F=t�>r�׼��R<���=�bL�J�>F�<T�1�=�>cq> e�>0Y?�	0?#�g?[B�>��H�w���m���[ �>�$>ݖ�>~J?=6>�/�>�$=?YB?x�H?$�>cm�=)��>��>�],��k�?���,e���V�:ei�?�.�?���>�6�<{Y&�@���|4������?�h0?�L ?�c�>�����v��t�g��=X����lL>=Z��(��<$սL�����;�4�=��>���>|1�>'��>��>޵�>Gh�>J8�=M@�+�#���9���F=�?d���=�Wj,���C=���=xG>���s�[��qڽ�[@>Ӂl>�9>+��=���={[�>�΅>��?A�T>�}��˅�>�{˾��9�'>�*]��]��Ib���p�4F	��+���E�>n�>�+������6�>`�=�XM>��?妅?�]�>_�>�ʾ�tݯ�6 
�$e�ӓ��B���R���-��L��6M��{ھ*C�>�>�A�>@Ä>p�&�HC���=b�����0����>k���V�����ؔd���������X^��Y���3?C�����=�t�?M(K?��?1��>ɷ������8>��e�_��=�3�QW�̮���?{?��>��ھ�A3��K̾����ݷ>u8I�p�O�����β0��K�&ŷ����>;����о�%3�f������F�B�+Wr���>�O?C�?)b�LX���XO�9���+���i?}g?��>�I?�B? ?���x�<n��?��=�n?ð�?�:�?$�
>Z��=oE�>?��R?�}�?"ȍ?���?V���F�>�h>S�[>��ͽTA��>�Җ>4��=i�?�^:?B1$?�]�<|�ܾʹ߾gྲ爼;w����>��>���>KfC>災�r>��[>�>�w�>���=��x>C(�>bD��lj�T�&?V�=�ȍ>�2?݊�>��V=,�����<
K�R?��N+��䷽�B��5�</4���aP=O?ͼ���>�ǿ�2�?�!T>�^���?wy���3��S>�DU>>�ݽ!��>�E>��}>�h�>�ˣ>g>k�>�N(>U�ľz�+>P^�i"���?�`�L��"Ͼ�>����nK����>ܽ?;���Ծr?����c�6�u���1�"J;F_�?w+�=l��"�������?�ҳ>�4?
,��������>���>L��>a���!	�����<�g �?���?<c>��>3�W?V�?͒1�U3�muZ�%�u�'A��e��`�����蜁���
�-
����_?\�x?�xA?H�<28z>�?��%�!Ϗ��*�>�/�:';��3<=',�>8(����`��Ӿr�þ(4�]KF>,�o?�$�?X?B[V�����A��=��I?�X?�
�?��9?�W?�����%%?h]'>��?o?��?�=>?���>�� =��o>�d>>+�j>l?��!݁�P_��=�4�/��;/��=�Ta>�	B�=�=�ɘ�|�S���l��RW<J>���;6I@=P��=��>!�;�%�>�[?�?	�>�=/?�hm�ݨ1�r�¾�F.?��>w�6��r~������+�c�=��_?l	�?�\M?\n5>�?�e.�(�Y><��>�O>r�>)��>�`��T��W{���=ց>5^	>���=�0��@R�i\����b��|�=,=?��>;#��x�5>��þݻ�����>t�^�g᷾AZ!���\���7���}���>��6?
?���=����
��,`��?NfR?iZ?נ�?����Ѿ�yP���H����y��>�E>�����薿�S���~<����;%}w>�׎�����7yq>��"�0$m��E����|��=��#�$<��yt辅���Sܴ=�&>��ľk�%�C�����J?�/C=�t���D�AK��^�">�ɗ>���>��ν���]qF��᧾�|�=��>��;>&�	�o��>�L�?����>ZG?�:r?Ʊ�?�H���Lu�G4(���#�E)޾���<U2?,/�>��?��>�K>'�����wv`�'E4����>χ�>�@���1.���V�s���!F�A=�=?F�>U�4>�Q?�*q?-?R�d?ȊN?���>�+V>������{<!?	�?r�U= ��y[_��A=�%=G��m�>+�,?|�O�^؅>Vr??�?�"?��G?�?^L>�����D�?ܙ>��>��W��ԭ�jF>tjN?ڃ�>}�Z?04?/�>so'�~[���0��e�=
>X)?9U$?��%?��>W~�>�3ʾۊ�>�#?��#?	 �?�y?�/��1��>f��>C2?��!=��>r�	?Jp�>)E?�(q?�%E?��?(k+=���1ӽW�N����=���<F�9=���=���K��v��F� ����:̼V���	�<պ�����<��>b>�>R*��#�#>���u���-eh=<���>���%@���X>ǲ>��|>(%>�
��M�1> 5 ?|�>��y�?�7-?��@?֧��g򁿸���]����
?�zR?�t�=�r��"��h�~���#=��v?Q�o?��h��侁�b?P�]?a�*=�H�þ��b�\��A�O?��
?��G�v޳>�~?��q?a��>��e��.n����K@b��j��=Zu�>�_��d��$�>ޞ7?�L�>��b>h��=#�۾l�w��g��g?B�?9 �?���?|"*>��n�5�s+�*ړ��'[?��>C�����?&�;�_Ҿv���}?��{;޾�I��H>�������2����������޾�'��=�&?Qv?IZn?kL]?t����kc�j�W��"|�d�V��������?���A��qB�)p�h@�(��������lS<�g{�˻B�rش?o�)?��/���>6�������Ⱦ�B>6���g���7�=����=^҆=�9\��(*�x֤���?OM�>���>!�;?HT���>���/��7�@�����1>���>s��>���>�	�::�)���彖�Ⱦ���g��7v>jsc?7�K?~�n?��v(1��n����!�;�0�~(��b�B>NF>6��>��W�O���(&��F>���r��������S�	��~="�2?gA�>~�>W�?r�?v	��s��BZx���1����<��>�i?2�>��>��Ͻ�� ����>��l?���>&�>����+Z!�}�{��ʽ&�>S�>���>��o>5�,��#\��j��y���9��s�=۩h?���S�`����>>R?Z�:_�G<|�>�v���!�����'�I�>�{?0��=a�;>=~ž=%�G�{��6��"N)?<E?Qᒾ>�*��~>�'"?��>�&�>�.�?\$�>�aþM�B��?�^?<J?RA?�I�>��=�䱽<*Ƚ��&���,=;��>�Z>H?m=҉�=���l\���I�D=�X�=��μ'W���<T���J<x�<��3>9ݿNU���ž?����Ҿ�J����?[Խ4�S����[��(p���Ύ���>�P����iQ���������GM����?u�?��x�����!ח��*w�������>e8a����l����b��̤��R�ž� &�*EP�up�8Tn�W"G?E������������,�+?
T&?Z�t?�E�����9�q�����4�P��=�'�>E����ȿ�􆾍#T?@K�>�zܾ���;፿=r��>���=E��>m�W�����%>��>��?�<?=n��}�п�5���	>�^�?97@@;?� ������QS��0??���=�N�Jg!���־;A�>���?�݈?�E�<$�V�ۊ��fbd?���=�+C��ZV;'ʫ=��_=,K=܎��[�o>�2�>�N&���<��'ܽ�.>�f�>hOH�ɍƽ>}Y�8E���c>ލ����5Մ?+{\��f���/��T��U>��T?�*�>Q:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?$�(?:ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=v6�艤�y���&V�y��=X��>f�>,������O��I��X��=����S� c�'���Fh>x��r_�����Y<��<��Ծ�]�ij���=��u>9a�>t��>e��>��>�I?4�m?Ja�>�e�>�\@�,�������Vyr���2�fx[��b�8����ݾ����>���#�I�@�sG2��%�����]>����}�
~0��9e�(fe���?;6?�ލ��O��?��C������Q�S=��>�R����B<b��T�?�??ʠ�f�d����� �=X`N��7�?��|��ho�1��j�o=�G�>T�=���>K�Ľް����Q�f�'�+?|�?����z⁾��D>)� ��H<X&?V?�5�<O�>i,!?V
 �͠-�� =>d$>>�>ě�>���=nW��A�W"?�O?=d�E���u�>�~��0�2��#�=�>�d�e���5>���:�X�7�R<�๽ ��=MLM?պ�>�.����a�:�$�?=�-��T#u?ї�>�+)>��c?�kN?(M�=����R�d��9>��b?-g??��>�pٽܾ>_��d�H?��n?&G>1�B������R*�,�̾$*6?�e?(!?��F�򏃿O�y��gƾ�Y:?��v?�n^�eq��j����V�:�>�U�>���>��9�gj�>��>?�#��E��N���	Y4���?0�@K��?��;<J@����=r=?�Z�>�O��Aƾ�f������m�q=[*�>І��gv����>Y,�ل8?���?�>a�������>��	.�?�ݑ?-�f�=�|��������Q�=�;>�����#����5�D(w�i�Ⱦߋ����=E�n>z�@S��=Ɲ?L�7=���&�տA?��2����yB?N(?��>Y�1�
������S�+hU�6��6p�>ڔ\>R�%���x��6�g]���>���=��L>�h�v븾B���J����>=��>'�t>bv��1оV��?Uo��ѿ�Y���B��b?dǗ?�O�?��>$�,�wR'���:��{	=��%?��i?��O?l-���ܑ��o"�1hr?�G��w�J���?�x�:�
&>�D?�"�>X�*�M/ >|N9b��>�Ȍ=���vѿ����L��);�?��?ۗ����>y�?��4?2KϾ!I��.�¾:=��6�<��B?��j>$���9�^a5���i�3�>+�1?�������^�_?)�a�N�p���-���ƽ�ۡ>��0��e\�*N�����Xe����@y����?M^�?h�?ߵ�� #�e6%?�>d����8Ǿ��<���>�(�>*N>\H_���u>����:�i	>���?�~�?Oj?���� ����U>
�}?�#�>��?Tc�=3X�>��=�()-��c#>��=��>���?i�M?�I�>�<�=c�8��/�~XF��DR�2#���C�/�>��a?��L?	Ob>� ����1��	!�Ymͽ�T1�^��_]@���,��߽K"5>��=>m#>��D��Ӿ��?�o� �ؿ�i��pm'�64?���>��?M��{�t�j���;_?e{�>7��+���%��TB�X��?=G�?��?�׾x?̼2>j�>GH�>��Խ����8�����7>��B?� ��D����o�F�>���?�@zծ?ai��	?���P��Sa~����7�W��=��7?�0��z>���>��=�nv�޻��W�s����>�B�?�{�?��>�l?��o�L�B���1=5M�>ʜk?�s?�Po���v�B>��?$������L��f?�
@~u@^�^?'��޿`ϲ��Z���đ�k��=6Y=Q�n>��m��$�=���=�w��!}�)��>7�>&.�>p1�>ZŪ>���>�f�>�ل�e�(��㗿�����:���9�
��w��������M���m��Ͱ�*�=����k���`��<D)�ŕ= `�={�U?5mQ?�do?7� ?Ĉ�z�>w����W=�R#��A=Ѻ�>�2?b4L?��)?@�=����he��[��Yɦ��%��{,�>Y�G>�z�>	F�>��>?�9XK>Q�?>���>��>x�0=����t=��N>�n�>N��>CS�>�Wz>S�q>���,�� �Z�`�t0ԾF�?LC=�Bd��Z��$���H��V9�7E?`�"��?����������"0?xG��ī��Ґ�f>�:?[�@?.>�ئ�����r�����<�)s���%=1̉��z[�KFF;�
?�qo>��>C�J��9�H�3����Z���sF?m���ɸ��D|��RM�Y޾�*=�=�>Ɣ>lLP������A������=PJZ?�O?U-�=L9���B���
���K>�Ť>%�(=���=<�=>��<�T���!=�N>,�>���=u��>��>��>	��>\)�݆D��s�>��=��>��>?K�*?M�½����ž���>�>\�?TӚ>|�k>�&'�a�=���>D >��꼲3'��pʽ�����>�O8�I$��!6���I�S�r={9>�H5>cW��;����=�~?���'䈿��ee���lD?Y+?� �=*�F<��"�D ���H��<�?o�@m�?��	��V�:�?�@�?!��Q��=}�>�֫>�ξ-�L��?��Ž-Ǣ���	�D)#�fS�?��?V�/�]ʋ�=l��6>�^%?ܰӾ��>6N��R�����3�u��q%=֣�>m=H?�c��naP��&>�HG
?��?��3����ȿ9hv����>)��?�ޔ?��m��#���@�ʹ�>}��?-uY?D�i>r�۾�Z�1��>��@?�R?g�>�`�w(�Q?CѶ?5��?��H>���?_�s?�P�>M�u��k/��&�������<�=�1x;�j�>'�>�����fF�F̓�UF��ʏj�޹�U�a>al%=0�>MM��5���1�=]���|Z��(Pe����>C�p>�I>$3�>O� ?I��> ݙ>R�=C���򀾙ܖ�d�K?���?z+��3n�w۶<
t�=��_��q?*X4?�T~��о<�>VG\?I��?F[?���>e!�f[���ο�����bi�<�M>�U�>x�>��t�K>1�վ�C����>��>b%�� �پ�ꁾ�λHȝ>�B!?�&�>m��=4� ?��#?A�j>[�>[ME�(;��y�E�'��>���>tN?N�~?�?Mڹ�W3�M ��ס�؁[�5N>
�x?Z?"�>�����}���iL��pI�E1��k��?lg?�0�?�)�?\�??�A?�if>�q��ؾr��ӫ�>��,?�Ɏ�E�U��`!��&��8�?�c�>1?����Q�}����#�
���>��Z?�I?�%�T�i��߾�(`=Ny���������L,̻�*�=�A>�Ҽ�׫=3�E>���<fn��@ެ�FL!>34=�#>D�H�Խ���=�<,?R�G��ڃ�y�=��r��wD���>�HL>�����^?�j=���{�~���x��3
U�� �?֠�?$k�?y����h��$=?��?�?T"�>K���}޾���nPw�^}x��w�o�>Y��>y�l���ݏ�������F��*�Ž@�ս5�>�o�>v?��?��a>uf?���c�:�#�k����3�W�� '���3�Y�L�B:0���s��wE�,^�=M���蕍��-O>GFK<��=x ?�١>�>�̬>YV�=��>!T>��>�ĥ>�*>��=[��=� >!�=��Q?Gt���(����)/��b�C?�ub?�:�>�d{�}���\��<� ?�֒?���?i r>�Bi��9*��?���>b4�c�	?��G=�[���m<������/됽!����>�@�v�:���K��[p�8�	?��?o��-�̾ֽ�Ġ��Ym=H�?��(?l�)���Q�]�o�a�W���R����|h�,u����$��p�㏿SW�����נ(�/�)=#�*?��?[�����?���k�z'?��Vf>��>�F�>��>��H>��	�w�1�j�]�.'��_��*D�>:@{?R`�>$�@?xW?�l?7?��M>���>H��\�>�'>q��>S�?�iW?w4?.s6?d�?,B8?���>�����������Y�>��?x�>'D?��?�<;��M;<��=SJ�<`{Ѿ+�K�b<|�Ҽ�Y�����k��=��>)?�v���}G���x�?>�t??l>:�> ���"����>��>?�,?�R�>Ӑ��v��#ڝ��;.?�
??���D�=��[>���=Jn=Y��<b[�=-�J���<���=Q�,����E+X>�a�e��<���<��a��D>΍�>��?���>='�>>��@ ��m�g��=c*]>jU>�`>]پ�3���R���g��Gz>q��?��?h m=���=D�=�K��bڿ��Z��{��>>�<�&?�k#?dHT?T.�?5s<?�)"?}�>�z�rr��sF���
�?��5?!��>Z���Z�����a�%��d?!�?t�[�ܑ̽�4�/CǾ�����U>�J�˹���E��.7�}t�=1g�������?��?�%=��D���׾T���ox��i�@?�6�>�ϳ>YD�>��߼e�*����Z>���>Y�H?$y�>�wO?Q��?��?v��>��@���� ���Y㼾���>z?P��?}�?�I�?��*?Ә�>��q�t_�p'پ_z(���]�8����<�=��+Yi>;D�>;q�>�:>�G,=rhH��*�!��=�&�=�[�>iF�>�s
?>3�>�J�=}�<?gr�>��ξ#l�����]����ս��n?@�?���>9�<L�7W0��� �ކ�>ۿ�?\��?ϙ?����J24>�Ͻ{��=lc��@�>��?K��>[P>0��e8G=�A?��>�̩��J!��2(�e��M?��a?���=��̿xρ���(�<ǈ=��ž�f�#'̽���<����
��V���@��<8��'����X�.X������?��><(>(~(=L���Y�=0�<[�=���=���=ar�=[wZ�0؏�=��<3*�<p!=$�H>*?O��(�(v˾�}?lI?Dp+?��C?�nx>E>�Q3���>�킽R�?h�U>w�P��p����;��>��}:��پK�׾��c�Rݟ�Z>P�I�<>k3>E��=T?�<&��=�s=c�=AD<��U=�k�=B|�=��=���=��>$>�6w?D��������4Q��Y�q�:?�8�>H{�=�ƾx@?��>>�2�������b��-?w��?�T�?3�?�si��d�>���㎽Dq�=���o=2>���=�2�S��>`�J>����J������4�?��@��??�ዿŢϿ�`/>[̉>'�M>ViS�� ������Uؽቀ�:T$?�C �����Q>Ū='/�������S=Y�>o1�=t�p��Zf��m>��1�C����!�<��Z>Vş>��>�ޚ�՚��SB=� >>A�>ER߽N�Լ���}�ɽd�=�]�>.tc>'��>Oe?� 5?�Gh?R:�>y�{�#�ƾ�I̾ꕁ>]t�=5��>��=��`>v�>��8?��C?�M?��>ꒉ=@��>���>��(�h�tO�8���U>=!�?�k�?_=�>�
��.�X�4:�ˑ>��\Ͻ�??�.?�y
?*-�>H������d ���.��雽Mv;�vZ=�r���z��`Y�d�+�L2�Rm#>1F�>`��>�^�>:��>(?j>:7m>I��>r��=
=<7�=D@�<�=�V�\=l��
��<:�0�+��:

1�u=��+��X�ϼ}��<95�;{����
>�e�>h�Z>S�>�`/>�v�����>1�����W���K>D���03��Rj��u�� �
R9��>>_��={���D��X�>m+#>Y��>�L�?@��?�-�>��!�C�۾疿:me�n���F�c:�/�;>A���"�6I�m�C���¾�r�>Q"�>K޻>�s�=�S�d;T�T� >�ξ!�1�h�?M���de�1sA��B�3���`���#I������<J?���\r>q��?S?��?�w�>������)���=
���$>���C���H��WkP?[>K?)�>�9�=�`�H���1�b0�>z���	H�����`3��b	�n�>�p��>"\����;hQ��Z���聿�+�c�
��=�>�V-?j��?��L���u��rj����o��>M�K?���>�G?9] ?�j%�|�ƾw�����=4-z?3��?�p�?�'�=�$�=����V]�>�?��?���?#&z?��L�XL�>~�^=��$>q���˧=���="ñ<瑐=>�?��?Tv?�-��~9��(���쾈%��1�<jը=I�>6��>2��>�r	>�Q=�Y�=9	k>Q��>��>/<N>]S�>�ę>u�y�w<
�.,/?%�<>��<�uI?kj	?�e׽*K�"֌>i��>��<����|'���e����="�+=�O>-ު>�O�> ſ捄?1��>����&?9(�(Q��Q�>H��b1%>��>�7Q>zw�>�a�>��?n�N>[��>��E>�!ƾ؃>�f�͎!���D�L�φ;M��>]O��'�*�U������rZ��'��	����f�]�����9��_<PT�?��L�h�-T,�(C�q�?-V�>l26?0ꑾb�e���>���>��>��j������uپ���?c��?�c>�	�>��W?��?sf1�H3�TjZ�ۜu�t�@���d���`��ݍ�������
�J5��E�_?��x?ugA?	L�<�cz>i��?��%�Nꏾ �>�/�5';���<=G*�>>+��IEa���Ӿ��þ���yF>��o?+�?#B?N�V��U��/�>��Y?��S?T�G?�v.?��C?�(���?,2�>y�?��	?��I?�B?��?��:>�*U>D��=��>W/�����)�]�%�����E�>�=Ts�=4�=��:r����ս��=����K�ͼ9v�� ��=��8>⚛>;�R?�(�>u҆>��9?ne"�dh0�p��"�:?���=��U�=F������h���9p=(c?��?�cW?9u>uM��DG���2>��P>'')>�#>ME�>m���[���>U�!>9(�=��P<�1�wr����@5�������g>�4�>�2>M���g+%>�X����{�M&f>�xQ������(S�ČG�\�1��
z���>K?Z?���=sh��Ϙ�U1f�we(?'<?+,N?��?��=�׾�::��RJ��:��R�>�ו<��[<���-���9�$|,;.�r>�d���k��ा=2y8��[Ǿ�t]�Cq)�1����t>�G��b�>����X6��/"���=2g�=������XW���ܨ�\�<?d�ٽM ���T��@�����<��H>k^�>߼�E�Ľ�A��Ⱦ��=�T�>��>�d���� �����",�j@e>�E?��d?��x?x�*gi�~;G����e��F,佀�?s�>��?��Z>���=]ܧ�Y6��Oj��$1��)�>/��>����z/��&����
��,��>6?'�f>�z�>�
>?%�?��S?�� ?ܗ?'ª>˨���̾�&?��?� �=��׽V`��:��RH�<��>@*?W�:��"�>�?�?D?��R?�M?� >�� �f<�┗>��>�X�����]R>gN?���>��X?1��?H>�v6���E!��2x�=H�>��-?� ?}?�k�>%�>b�	��"!>��>�5~?g��?G	�?�a�@?lL�>8��>��>�0�=��>U�>g[C?�YN?�$?���>���<kX��jC���2���&�<�B�=W/.��B;_i齠�C�(�/��Z��ɣa�+\������+��=c���8�
���>VM\>;1���۴=��㾽�L��jG>�#��1������'#����=� 7>��> 3�>U"��[�;�Z�>�~�>[���"?%\?!�%?9���T�������:;�>�2.?cȮ=�1g��ӊ�)�o�F�%=`�r?�W?i���v��L�b? �]?-h��=��þY�b�Ӊ�g�O?=�
?��G���>��~?b�q?5��>��e�:n����Cb���j�Ѷ=Gr�>HX�?�d�w?�>m�7?�N�>��b>m%�=mu۾�w��q��j?��?�?���?p**>_�n�P4�@Sܾ㤋�dY[?2�?U�E�5�B?��T=������{����0������:������Z��d�i��F � �>0	?�f?a�s?\LW?s��UoO��_���d��=m��S&����iR�<�6��4�7�J���&�v���ꢾ�z���|��?��7�?V(?�6%���>�q���i��ƾ�7>�����Pϖ=�7���K=	v=9�c�H5�Uz����?���>�j�>A�<?r�Z���?�0 1��4�SO�\'>n��>AQ�>l��>3ٶ:��)���ٖɾ������㽐Mu>&�c?ּK?��n?oF � 1��c����!�Ǐ.����iB>��>O�>�1V�[_��.&��8>��+s�?���g��Α	���|=1�2?���>�ћ>�!�?ư?��!��>Lx���0���<���>��h?��>���>�!ν1� ����>��l?���>�>�����Y!�}�{�V�ʽ2%�>*ۭ>���>��o>��,�#\��i�������9��q�=�h?������`�;�>�R?Lǉ:!�G<{�>�v��!�/���'��>�}?͘�=��;>P~ž�"�`�{��5����/?n0)?�U�"@�N��=_?ic�>��>��?�i�>��3�l���&?LyL? j?�93?{�>���=<l�]��_D��8�=�V�>�F�>��<��N>Nv��#\'��3=���/����;;�$=b'=�3��Aл��zŽ��i>U�<<�c�[���˾W>(��������%�q�����J����,���ԾZG���t��;��)��]*n�VA��k�E��q�%��?��?Z���-yﾹ0���E^��mɾ]J?ZB������Վ�������h�m��R>���`���X��8�4�`���O?�aҾB����������
?wN?�g?n\���+��7��<�ϱ=�G+>�D��'�����2���W?A��>�����!�>�A_>Y+>)p>Ĳ�|�0��R8=VQX>vP�?�i?���L�࿋6߿yg~�r��?��@){A?$�(�6�쾄V=ƶ�>f�	?��?>�)1�K�갾X^�>�0�?l��?DSM=ǽW�R
���e?�A<��F�TۻM��=���=x/=��e�J>mZ�>���sA�.#ܽ~�4>iƅ>�x"����e^�Z��<�k]>,�սJ!��4Մ?	{\�tf���/��T��U>��T?+�>�:�=��,?d7H�W}Ͽ�\��*a?�0�?��?&�(?&ۿ��ؚ>��ܾ�M?YD6?���>�d&��t�b��=W8Ἄ�������&V����=a��>��>��,�݋�߇O�$G�����=�u��|ȿ8��#��q<k�7���p��b��㽏8��mԭ�/�Z����YI=u/�=��8>�>u>#�W>�L>�\?V'l?��>�=>��n���j=þyun=�ac��#�[���J��ML����ܾL\׾Q�� ���j	�;�;imM��T��L�|��?�=��%�ڝ"�r�1?�Z�=��従',��;�F�¾�z��	�<0�����A��98b��@�?
C?�h��6X�l���L@;݀���r?�?����Ⱦ?!�5��=���=!�<��]>m���\^��hM�ײ8���$?�.?0X���������=A��ʐ�l�)?�<�>T|����>�?��K��hϽ�y�>M>���>u3�>��>ûƾlㅽn:?��F?�F�Q�����4>��ؾ��0�$���J
!>�K��Cɝ=9�R>z��<a�%bg�d���]��=>�R? ��>����o&�LѾ��=G�3}?QD�>���>7l7?�(?z��=�/�t����>�b4?>Ee?!�/>=Oݽn	�g�ľc�%?:ց?,~�>;8���z�����	�.�>��h?��R?�4�=SȄ�\u�����e�+?��v?s^�xs�����R�V�m=�>�[�>���>��9��k�>�>?�#��G������vY4�!Þ?��@���?,�;<��Q��=�;?i\�>�O��>ƾ�z�������q=�"�>����}ev�����Q,�e�8?ݠ�?���>������.?�=Y�F�@�?�l�?Gq�9�>8��k��C߾Ys���X�;^��)��A0<�����~��L�_� �EUH>KZ@��z=?W�>�����忬�ȿ������{���D��>��>�|>��P�4uJ�|s��U�
Ve��I̾�1�>�Vk≯	���D�N��8�,�)�I���?$u<JP>\dz=�� �	�F%���:�>��?�>nmT�D���`�?rF �z ڿD�v������_?ᚕ?쁃?yQ@>:߇>;%��b��4s#>�?�s?ZL&?�M�=���_"�9�u?�ʾ=oN��b ���N��:1>��F?V7�>�4-��t�=�C�="1?=�>]F ��1ܿ�Nտ��"��?��?�� �.�?��?��?����%���C�G�1��E���A|?j��>�냾X1�_3Q�EGQ��n�>�4+?mX��n�U�_?
�^�1�o���.���Ͻ!�>�4�v?W��ڼp���e�p���1t���?-�?C��?���"��x%?kޮ>hm���Ǿ�l�<p~�>s)�>̱U>*�y�v>�U�0�:���>�0�?K�?�?ޭ��`��?)>�
|?Nܦ>${?�>ߵ�>^V�=���M�-�+>��=��	���?�+F?�c�>�A>�t ���$���=���J���ݾK�A��͉>�*q?=�P?���=#%4�d���#���<:�X��p�J)�R��<��ou!>3f>\�=@q��:���?Ip�7�ؿ�i��4p'��54?'��>�?��u�t�P���;_?Sz�>�6��+���%���B�]��?�G�??�?��׾�S̼�>I�>�I�>3�Խ����f�����7>2�B?e��D��j�o�|�>���?�@�ծ?ai��	?���P��Ta~�'��q7����=��7?�0��z>���>U�=�nv�ܻ��M�s����>�B�?�{�?��>%�l?��o�c�B�6�1=nM�>��k?�s?!Fo��󾡲B>��?"�������K��f?�
@wu@[�^? ����,��ʉ�\���������2�n=�憾msh��K�=�ǈ�� ���<LU>v 1>X<>#S�=�>w�	=�A���x#������5�6����X�(��k��vc�V��V[��0;\�)Ȫ��J���4���֕��8%��KM�0�=��^?.CY?o?��	?�䫽&>Gv�2=Sk>��Z=�1�>f]@?��Y?��!?.BD=����h�Vx������灾ߴ�>+rZ>o#�>��>D�>� ;6�C>*��=�J`>�%/>ߊ>��=ev=�)[>�>�?���>H�>B	�=.H������<r���_��~z���?��þ�A��s�E���b��Y��=.�?�/E>b��Z�ؿbʹ��:?=߲�p����b��">�� ?sMf?.�=�1��� �l<�i��Փ���a>=�[�e���F]��T>�$?^	B>�C>�pF���(�4�R�C���X��=~_1?����b����7�:�S����ޜ�=0��>�|a����rw�ի���ԍ��G>��S?��?r~��xL���ɨ�۾��>(0�=���;Q�=S��=�8�"��(���>��7<��>�`?4�>$	�<%ZQ>�hx��1۽��>k�>�e=\� ?��<?�J��W�8�5]��g���$>���>E&�>^�e>	䒾Q��=8�?]:^>7�6��.s��|��a��Ζ�>kJH��LQ���7<��#>�v׽�>�|�=��|��l��4��=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�_�>;�����F����w�
�L=��>yI?�	��	�Q���4�|�?��?y����o��wȿ�Lp�8�>�,�?��?jm��@����>��A�>���?�6Y?��k>?a�?
D�*=�>�<?�PR?滶>�X��S0��?�?�?Ϡ�?��>��?�ȃ?i�>u=�!�6��^���F��<.��"�>�/>����-��/��+ډ�ӂr��VI�g�$>�»��>�<�Lվ!�>�I8��Sm�LHm�oԱ>�N�>?�=>��>A�*?M?���>���=X�����[�H�K?�?����4n����<���=��^��%?=X4?�Y��ϾB��>��\?ƽ�?`[?�f�>����+���ܿ��������<��K>�S�>�f�>�S��VZK>�վ�C�\j�>}ʗ>�k���-ھN!���L��B�>rX!?ư�>��=0� ?J�#?�mj>�>�pE��+���E�(��>&��>`%?g�~?��?'̹��W3������ۡ��o[��DN>�x?�]?���>瓏��w���D�dG�vr�����?Cg?��N�?��?̧??��A?f>�����׾ṱ���>�a#?��\��Si����=�ƽ�t�>�@x>�?��6�����w8���A:?�[?�4?����Y9����<V�^=�=�F<ջ< R>5�>JqԼ�%�=����L>U��v��Y�U�#5#=U�S>�n>�.ݽ����0,?5�E�烾�ј=��r�uD��>�_L>y��� }^?�H=�v�{�����v����T�1�?O��?�c�?0N��8�h��"=?�*�?u?��>NE����޾+���/w��x�V��U>���>�l����|��򆪿�7��F�Ľ@����>*U�>��?��+?�)�>�A?�Ӿ_�����f����/�v"6���A��:�����h��mՒ���=;˺�N��vKM>
S����>���>�s>i
�>܎�>��e��"�>�6=��F>��>Ί>��N>oI#>�h�=^U���GR?2���+�'����{���3B?3id?�6�>��i������1v?F��?`o�?Mv>�{h��"+�p?�=�>����m
?��:=�r�Ո<sO��*���i��*��s��>?!׽�:��	M�Kff�h
?</?M���&�̾� ׽����Eo=]N�?�(?t�)���Q�s�o���W��S�A��n;h��h���$�טp��돿<^���$���(�nG*=υ*?	�?�9�����)k�?��Kf>%��>�'�>�ؾ>ooI>��	���1�(�]��J'�η��xF�>tU{?���>3�@?¶D?��<?�<>?ᦇ>U'�>c첾#{,?X�[>�g>�*�>I?9�?��?�e?�4?|�>��;Ɩ��u(��(?�>?�`&?Y�>�V?̓׾[��H��=�܌>3��t�ؽ�
=��������&=c]�#�>=f)?�t��HeV�T��<=�>Ab?���>���>L�8�:�S�rr?N�=ֹ�>P��>pi� X(���K��,4?��]?����;�y8>&�w��j~>ks-���X>�qj=�Q=�;<%T'=���=cˡ;SD>��t����=Ǫ�No:=�Ɔ���>��?���>⟇>���
����f����=X�U>of7>d�)>�־�U��r���w�b��nv>�t�?U��?O�^=�n>G��=�����������'��{)=�b?H�?{gV?:�?��8?G�*?>W^�|,������o᣾O�?^�*?�
�>w��Dɾ:p����2��?D�?gj^����H'���žav���1>@-�Fo|�ҭ��0A��:K��K�����x��?Nz�?��v���5��~�o���D���7??]�>W0�>	��>ҽ)���e����B>�U�>TTU?�1>_y�?�D�?��a?���>���ۛi�;b��>3�;�!�mE�>�u�?���?�n�?3��>;��;~!�)U澶Ҳ���m��^��v�
���=RA >ݔ�>cs�>y�>FO�=��1��D'������>��>��>˙�>��>	?G �=RtJ?S�?j���G�43��<y���at�y�?(�?�p>?�[`�{M��a'���?�<	�>ǧ�?���?�?�N�R>5Qx��N־`C�AɊ>G%?.�>x>��}<�fs>^�>LZ�>�k �½辳�1�63M�u�?ިB?�G>��Ͽ);�u����Vݾk�����q� Y�0���|����!<q�̾����ԾEUW����������C־Z=O�7����>�U�=�K�<m��=��=3��/����`<�L�A�=�=+�o�q�����=�_�j/���==ʑ�;9p=H�˾V7�?�D?<r*?�zO?�^>|�J>�'����>��x�D�? J}>��������q�����{���L�羕���]a�՜����=��U��)>61;>m��=��;�f7>�,�=L!�=�_e�2�=@�>�}=��>x��=i	(>f*>H6w?$���+����4Q��Y�$�:?C7�>y~�=��ƾ~@?I�>>�2��T���:b��,?��?jT�?��?�ui��d�>!��⎽u�=F���a:2>T��=��2�⣹>�J>��K��R���b4�?y�@}�??⋿g�Ͽ1^/>�/>pW(�~�oF����\�9�G͝��E?<�#���˾$��>��V�Uy�8���d1�>�=<��x��S>�܃�\��=�̎=k`=�Di>�?4>w�>�=e��E�= ��<���>:��=�0~�i=<I<�c>>��=�0>�f�>ǟ??�to?}�?��>��Z��"��鹾�Ui>^)�D�R>,B�>{��>��>�l?�J}?��n?n�d>n��={��>"B?>��,���0������-塾4��?};U?���>��,>���8dN�w��I>K
:?(2?_?>/>���]�㿐^�:3����������G=s���W9��C5�۷��X�Z���<s�c>�$�>��V>�!>��G>g�0>���>��=�İ=�&<@.���BL=�#��F>\=�	�w��=
�<�>�et=Z����^�=R��V�^<�(������"�=*2�>ش>Э�>x2�=.ĳ�Z�0>n떾݈L�3z�=�O����A��d�nI~��
/�7���B>��V>�؂��'����?�fY>m�?>��? u?� >���w�Ծ\d��g�d�9�S����=?		>&�<��;�p�_��M�9jҾb��>(�>Cݽ>:Yc> ���\7��3>[��4i>�>�5?)�P����>�dF��ց�ly���D��W>y���3�'Dd?�j��?z?��w?��,?.��?�!�>�aM=K�Ř>����P�R�־Aa�p��KY?E�Y?Rj.?��0��PR��˾P���g��>
�K���P�7���]�0��+���o��ֵ�>�訾��Ѿ122��e�������>B�<�o����>��N?;߮?\9c�:灿��N�V��\����?_�g?�Ϝ>a�?��?����������=��m?)�?G��?�
>�*j< G.���	?�
 ?���?Ʌx?yz?��ʾ	�3?�X�>&�=0��=�$�=*�<=�t8���m>�?���>	�?����X��2�Ⱦ�ϙ��`��>�[�=�6>Y��>��P>ӛ=��;:�����2>4��>V>�>���= �>#$->���4�;¯?��>��>g�;?8N�>�=o��+M>���=�4нG2�<�b�(҅������=,��=�&u<�e�=�	�>UJȿ��?�w�>d�0���B?�p	�o�һ]i�=�s�=Gp$��B�>-��=���=���>���>��7=�X�>���=��Ͼ!n>�����$�v�W�:�<�	ܾB��>�ؚ�V8�Y���t)��E8��ƾ����F�^��
m�f�9�@�M�?��	��Y���&��������>R��>��F?Td�� t<�M�=�x�>���>�=��h5���Ԋ��]��\�?Ð�?Ic>��>z�W?��?cX1�r93��zZ��u�KA��e��`�$؍�w����
�i��~�_?�x?�pA?�Β<|3z>���?��%�������>4/��);���<=4��>w0��}S`��ӾV�þl,�{tF>k�o?R�?aF?/V�9���x�$<?6�:?�o?��;?=b?����eM?_��>,8?�&?��%?�>s5�>�҆>�,>��'=�">W���&�������"���伐�=Ў�=�`�<T����==y�=�ϙ�ڐ���FY�1��@L=��)�f�=	�]<df�>��a?���>�S[>l2)?�����4�ʼ���0;?ZS�=����q҄�"�}����m�)>ff?H��?ڎ`?�1]>�oV���e�c�>>��>�e>g7Q>�5�>�m)�~�)�n�=u�,>��)>��=J#��e�����F��KL=�u(>Bx�>c��>&١��i>�����"{�X.W>uI>��k���_��KE�"J2�-��%��>��I?�?�ߤ=�aݾfN��(�f�vQ&?�C?ݬM?=�v?n
�=��ھ�=��ID���$�}�>N�6=W������� �q�3�>;T<|r>�N���䀾�.U>�{���ݾ�-d���8��4�=0����<@��<xݾ�ā��">��0>|��v)#����V��l�D?K=,���N���پq37>Z�>|_�>�������ߊ;��Lƾ�)�=���>hE>x�!<8侰Z[�J���O6�>rE?��^?�&�?����%�q���A�5���G�������8�?Sج>ɓ?��C>0@�=K���S���d�)�F���>a�>���5�G�0���M]�Ǌ$�[��>��?(] >s�?��O?��
?LFa?�+?ف?)��>Aǽ)y��z�$?NS�?���=h����F�Z�E���P����>�A?0l1�)e>�\?1?	�"?�@I?>�?t_>�(߾�~0��6�>�Ώ>dTV�|���ҧW>"�Q?���>��T?Z��?΢I>�K�F���h=�& >{F�=��?�Z?n4	?
Ū>��>�E��]��8��>t&O?�?�xV?X�>B��>��>���>a��=Rr�><��>�?�C?U�i?��=?���>�	=�bͽ�i��$r�����;�jN=5|�=�i�<b�C���߽D�����=�P��b;�<%�Ľ�[���ý��><�=�Ҟ>U/y>h���Ӕ=t�A�>a�����>��>9�\��	�"L����>��>��>¸>��@�EC�=6��>)*�>�|����)?�?�a@?�-���q�Ȱ�[ƾN��>US\?�=�>	�7�	˝�`Έ�MC`>Z|?�6?���]�Z?"�X?�"�Xc-��=���IC���־�
A?�,�> ���H�>m~?Hn?G?�f���j�P����c�4o���>Ϥ>��e�`��n>n�,?s��>E�>%��=xnþ\;o�z�ܾ�8?�,�?+ٲ?�܉?�l�=2_����㿗#��$��|rg?���>�_����?ɿ7=�K�Ç&�$݁��0�dIA��@���㦾�ܯ�4c;�#s����o>��?]�w?4�?��R?|��M�n�jMm��Al�-rg�X�jD �ޚF�;:�Y�D��)o��#����Z����I[<�}�L#B��I�?n�'?�+���>,��$*��a�þH@E>cԢ����Ӱ�=����K�0=pU=�Eg��t1��6����?���>l�>��;?L�[���>��h2���5��"���0>�t�>��>=��>��8�&0�n�K�ƾt��Ozҽ��j>x�f?�R?iq?�Ӛ�T=1�����A%�zj���𞾐">�>���>�4�!���%��5��q�XR�U.���c
���=��1?��v>�;�>$_�?��
?'��tr��;c��e'��)�<���>�Ui?̪�>�؝>��ý�4"����>d�g?,G�>	��>� z�� �9�X�;"��N�>Z6>�F?a��>�A��GR�ŧ������g,�}��=�`_?�~��>m��><�6?\Ti<�Ԁ�^�Z>�"��$'�$�ܾ��2���=�a?r�]>�_W>�ɾT8������ξW�&?��?h%f�{�&���v>?���>��>��?fL�>
9��P����'?�a?RC?߫D?�j?���=������ҽ�6�T6�<���>Ta>n5.>��+>q�0�]��%���>T��=�
t�	�$�r==�HG�^��;!�o=�i>ؒѿlpZ����%#���޾��޾�v�������?���}v�I	���*���^�8�G��]B���5������쌾fah�t��?�5�?7񼾻Ǿ� ��.�b��Bھ�$?�	f��O��䲾�ͽ�w&�1������dJ�+&<�FE�*]*�ѻ??�Ɇ�'𪿍D���O��}�8?>�F?4+{?�Ҧ��$8�$U辰��=;P�<$=�=Z5��\ޏ� V߿jL{��yV?nt�>��پ�|*��թ>���>�V>�>$h��f��Pֻ���?��k?���>x�c���ؿY�ۿYR�=���?��@A?��$�50�Ō=�>�I?�C>�#�?�3*��
��>�ӝ?(�?z%=�(S�^@��d?�;S< �<�=Mb�W�=�8�=��9=3`��DC>���>m�,�S <��#�k7>a&�>�x�����a��1:<$]>��ҽ�(��4Մ?){\��f���/��T��	U>��T?+�>2:�=��,?X7H�`}Ͽ�\��*a?�0�?���?�(?=ۿ��ؚ>��ܾ��M?^D6?���>�d&��t���=X6�܊��|���&V�l��=S��>V�>,�ߋ���O��J��^��=�7���*˿������o+=��A<W���IP.��w�P�ý&G���qe�sV��<���=��>��h>�gL>��$>�_?��l??��> C�=T�T�[�S��ھ�,�=�hJ��j?���r�&���#�������̾���M ������þ6A6�F-	=��N�V��s47���N��(:�.�C?n�=?���T>�a��<��u3��ĉ�:�_���¾co��T����?@AO?�!x�D�F�C�.�+q��LW�;�Z?'C���,��7>F!K<���=���>P�'��(��_��>6�<c-?��?B���]�_��_�=�b ��='� ?���>�����{�>"�/?�w���'�2>F�>+��>���>d�D>*w���|��g0?�D?�_��y෾�~�>�վ<1x�AJ�<��>�j��+ba�Նd>��,;Ҩ���T��*ν��6�,T?��>_K.�U���ҟ�*�}�פ+=��u?�1�>~�>o?��2?zGa=�&���
D��}� �U=��V?\?��&>AfĽ1������j;?X�l?��D>�u{�y����"��2���?��j?}�?0;:�;y�����]���3?��v?�r^�Ys��5��	�V��=�>d\�>���>Y�9��j�>*�>?�	#�xG��ﺿ�"Y4��?e�@G��?��;<x#���=�;?^\�>��O�/?ƾ�y��.���~�q="�>D����dv�����R,�"�8?���?l��>擂�ܩ�(��=`4|�]�?xf�?��8����*�]�v���ھ���<�0���7<1�-��0��.F�\)�����)_Ҿ�=S�X>ʖ@�|L=�F�>x�����ؿԿ��Vp�܂+�ԏ�>�b�=�Sѽ��þ8p�k�x��O��B��:�����>=#>�j+�9������:��'�=�U?���<x[���u�=�ݾ�N[��]¼�s�>��>��>Pϐ��������?���5ؿ����P���at?/<�?4�{?�_�>���=��2�ۊ��%�>ۍB?��R?��?41d� i����?��n?ϭ��B6�T.�Pc!��8�>1�O?���>o
��>H�[>�?F?�I>��x׿P�ͿU�9ٮ?`��?E'��?H��? �?�(:�n��Tｾ(;��y���g}?�=V�����9��ui���q�>�X?�l*�y��t�_?��a��p���-���ƽ�ۡ>�0��b\��G��ۤ��We�*��L@y����?0^�?G�?����#��5%?#�>r����8Ǿ���<���>4)�>�)N>�G_�D�u>?���:��j	>��?�}�?�i?�������Y>��}?1X�>t��?�`�=��>h^�=�����R���#>��=�DH�i�?M�M?�,�>O�=�:9�v�.� �E��Q��x��C����>�db?�$L?F�b>$)���/�g!�H�̽/F2�_���z>��+�s߽n$4>��<>� >h�D��|Ӿu�?p��ؿj���t'�654?���>��?��o�t����<_?�z�>I6��+���%���A�A��?`G�?$�?ٹ׾�K̼Q>�>�G�>��Խ����.���U�7>��B?,��D��%�o���>���?׶@�ծ? i��	?���P��*a~�[��U7�H��=��7?g0�y�z>���>��=ov�߻��
�s����>�B�?�{�?���>�l?m�o�&�B���1=BM�>��k?�s?�ko�<�?�B>��?,������$L��f?�
@lu@>�^?+�ݿHâ������Ѿi��=�g����=�K���!=��f>�!E��_���o�;�Z>�j>`s]>��*> U=o0�=����|*!������r��Ƈ7�'
)�(���y�����%�`��[#�J�;��ƾt΃��r��8�Y�{���L�-�ս���=�$S?^?ǲ�?�-?�g�ה�>x{�����/��Oɜ<шo>��I?�fW?'m=?��,>��t�n�]�!8s��͇��M��C�>��>��>u6�>Q��>�a��`P>��<>�>+��=�4���=ϴ�=��a>�}�>�p�>6�>�-�>�&>!�?���F`�K2��J��?�n���+:���y�.�V���27>��G?�:�>�0����տ~����D?�W����"��:+�F�%>-?��K?�zO>����R�=i#�=X�	��%@���=8*���95��.���>��3?��>p��>y�G�.�2��`��>��<>.�J?��pC����F��Qk��"��ۀ>���>5s�:�3����g���~��*K=>�{[?㽵>H��1���Atc��Ӿ�Ty>�8�=恵>�߬=�8�=?C���4Խ�����\">��o�a�Y>jy?��&>�H�/��>�Ȿ"p�F�>�!k>u�>�?.?8V=Qp������H2��tg>_#�>�o�><4v>�o�_f>t�?"�m>�{y��^̽[�#�>����=^>����g+���)=R�M=�a��۷J=�Ca<�{���r��T <�~?���'䈿��5e���lD?R+?� �=��F<��"�C ���H��F�?q�@m�?��	�ޢV�@�?�@�?
��e��=}�>	׫>�ξ�L��?��Ž5Ǣ�ʔ	�1)#�jS�?��?��/�Xʋ�<l��6>�^%?��Ӿ�W�>ې��T������v��&=�z�>HH?4t���_V���;���	?�C?�A�>��%�ȿ�@v�+B�>��?��?I�m�wg����?�y��>�?gY?g>h>z:ܾvSY��G�>�F@?��Q?	��>D,��)(��f?���?/��??R�=��?��?�0�>n��>8�R�m ��c�����\�+��>�o��ּR(�ŒU�u ��Q�����q��O)�#�b>�w�<���>���2%[�P�=�6��^�����>�{�>�4�>p3i>]3?տ?�F�>H��=뭩�1!�P�����K??��?6���1n��,�<Μ�=��^�F(?F4?�G[�\�Ͼ Ψ>�\?���?�[?�d�>���=��Y迿�{��&��<[�K>4�>;E�>���DK>��Ծ�2D�pq�>�Η>G주�:ھU-���6��\@�>7e!?1��>�߮=�� ?��#?G�j>�(�>�`E�}9����E���>��>�G? �~?9�?�ӹ�Z3�����桿|�[�/:N><�x?V?�ɕ>(���ă���|E�^CI�O���l��?�sg?�Q��?~1�?ԉ??ѥA?S+f>3���ؾư����>8�'?�<�[Gc��)���<�D�>��K>�W?��*���=�HM�<3�|N�M4?a�a?�?��"�?]�v:��?9=�&L=�Q��(�s:��tʞ=��>���=�w�=��=��&�����	�����=�>*Y>N��w2��+�D�*?��<L��V�=ap�=06�a_�>L2A>���m[K?h��#�j��I���䜿�<_����?���?���?�ae�	vk�*�<?ʿ�?Tn?/v�>PqþS�۾�M��'X��$�~��s���>s��>����`��X���l��O�����d�@�b?�Q�>(?�e.?�J@>��>R�;�t$��h־��sr��$���R���?�_�&�*s���GI�o�=H���"���"�>J^;;��>�G?��>mM>e�>�=	��%7>&��>��>W��>�B�>��Y>�l�=1<�x��>`D?�׹���&�[� �/��wW7?Լ`?�u?�"���Ȏ����%?9̏?��?��r>�k�)� �$?�2?�a�sk?�n=u�L=�\-�b�Ҿ҈���{ɽ (;7��>c�x[!��0L��j�b�?h	?��<D"����������=9Ԇ? �(?�#��P�\q�s�Z�:tQ�]���b��丣�m�&��s�ݻ��'Z���8��M +���4=��'?8�?�0��p�w��$�j���@�r�V>�Y�>��>g��>��9>t��B0�z:^�*�$����	�>bv?�6k>�eN?>xU?mk{?�X^?��k>ȭ�>�+Ͼ[�?K
>�Fk>�R�>{o?��
?�.?.>?�[q?�W�>��h|��ɫ�t��>��V?u�?5��>�q#?�?���rϾ�6m>��>;'���rF�0F�=��.>��=�����U�=��>R�5?��^��CP��O3�2�E>���?�͓>E��>z?��U;��=Y$�>M��=���>���� �������>ϭ{?�vƼ7�_=��=��<1t��2�=��>��\=��1>�i�<"�v�L<�,=��%�!���o�"�&�e<b�B;��><t�>�?��>6@�>@���� �й��~�="1Y>9S>n
>�=پ�|��b"����g��ty>1y�?I{�?�f=f �=��=����g��H����I��<��?�K#?uVT?O��?�=?!o#?��>n-��L��\�����&�?�;,?aD�>�����ʾF����!3���?�e?�
a����(�����
ӽ��>2o/���~����"�C�����������?��?�C���6�M%�u���б����C?]��>��>���>Q�)�*eh��G��=>_��>�1R?V�>e�d?���?>�i?'��>7�8�-´��4����=�mB>-� ?d?���?��u?�R�>���<��Z���������a6�������=WWA>��>�%?�6?��A>�<��x����X���>�>�{ ?���>s*?(�h>�����>? !�>��� ��6_��^���g�z�N7x?�4�?OA/?b�k��7�����޾�H�>��?s��?h�"?�2�:->(X���p��F� ���>H?B��>�*=90�<=H�>��h>L�>�u=����V,5�x�:��^'?��4?Q�>�οJ䁿,�m�Zm��,]�<�(��9����o�l�z�#q�=Ҡ���I�热�����	װ��Zv�g#���t��:���E�>���<�I>���=�
=":Y��G��*�B����C����Z��I��<�tO<\Zl<5^a�ޓ�<eI�<IQ�=��:n�˾!�}?U;I?�+?��C?U�y>�Z>R4����>����:?W�U>o�P�������;�δ��t%��˵ؾ�j׾!�c�:՟�H>�%I���>�R3>�X�=:�<Mc�=�s=�=�1G��F=LM�=ބ�=eu�='��=�>�c>�6w?X�������4Q��Z罤�:?�8�>h{�=��ƾq@?��>>�2������xb��-?���?�T�?>�?Eti��d�>K���㎽�q�=<����=2>n��=s�2�V��>��J>���K��F����4�?��@��??�ዿϢϿ0a/>aN�>�%=P�_�4��ʣ�����v6��#�?ў7�BU��0�?��gݾ�P�� j>>z/>�ƾ�I�ٽ�~s�r�>@5�X{M=�x0=k�>�݌=0����<щ�=D�>�F��S>i��jn=��m�z�p>{����s�=I0�<��>�+?t�R?CX�?�U�>E��X�s�x�Ӿ?��>cŻ>G�>9�'>��
?\?4�s?��y?S�>�A�=z�>���>Ӝ9��ݛ�q����P����?煢?N<�=�cn�%����l@���:�̅���?�"L?�r1?Bm�>i4�ۢ�	���wB��F��L�W�k�ʽɾ�+U���������6���=�\>�*T>���>���>�k>��*=���>�B=cԢ��o�=[x�y�$>��<�E�<S��b�ͽ�8�=� �=��<��=�$*=� �=�J��0	�=?ך<"p�=���>��P>�˻>��>�n��_�d>�߸�;OI����=|�KL���u��L���>�3����]>ql>��Ӽ�����p ?J�q>|iG>��?�<h?}�b>X4�-;Ծ�բ�b���'���|>5�>>A׽�v�\�=�O�Ћ��8��>H�>*��>�5>Cj&��Q9�.
�=t�쾁�*�p�?�$
��9�<z?��N�����;���,|T�	�n=NU?�����>��?��G?놔?�J�>Ue���/��3��=�9��ӈ�=k�J��z��VHq�|�;?@	9?���>��"�j(q��I̾6$���ַ>ZI�8 P�����خ0�a���η�P}�>i���o�о�3�3e������
�B�INr�$��>ȴO?x�?�b�V��*SO����;��*t?�g?b�>AC?<?� ��Xq�g��K~�=��n?6��?u<�?�>~#�=����Ѷ�>$�	?�֖?�r�?{�s?F�A�l��>���;b? >៘��J�=
>k��=c��=�?u
?��
?'ϛ�$X
��Bﾚ��_��� ='y�=޽�>��>ʥr>���=�	t=�ɟ=he]>�A�>h"�>�f>i�>�l�>A������k 3?�8F>]N�>��4?�b�>�-�"�>��=�i� -�������W�������rQ�br���=�j�>�qο�V�?,�T>��*�u?�����g�H��>�V[> �w�ZZ?��>�u�>��>�8�>=0g>G;>)c.>r(Ծ��=�j�I�+��I�� G�	Mо��>�����g�{0�w���P�0����i���{Qh�b�}�� 2�ǫ=���?�&y���g���(���U��4 ?!Ѵ>��>?�U��Cf轻��=A��>�%�>aGھ𛎿%*��zX̾�:�?
��?�;c>��>H�W?�?ܒ1�^3�vZ�"�u�^(A�$e�Q�`��፿�����
�q��*�_?�x?/yA?S�<0:z>Q��?��%�nӏ��)�>�/�(';�!@<=t+�>*��?�`���Ӿl�þ�7��HF>��o?7%�?rY?>TV���k��&>B�:?�1?L5t?��1?��;?����$?~:4>X:?�m?�B5?y�.?�
?L2>�T�=y8����(=�Ñ�<���=�ѽ��ɽ���9�4=@"|=������
<��=kW�<����޼-i4;,o��1^�<5�9=�?�=S��=��>�t?��?�'>{�!?X����0�o*�K]�?_Έ=,w���g���<?-~���=�dp?I��?!zV?��>v6�P.!��n�=�+�>�>0�>��?H��������M=(�=�p�=S>�,,���4�\s�_8���А�g�%=Q��>}D}>����7)>G����u�~Ig>��P� m��qzW�n�F�[�0��&u�3#�>�K?#z?��= 辙���hf��*)?dA=?�L?��?>D�=62۾Ә:��xJ��,���>�f�<z��B8���ܡ�a�:��w���q>����>�z��>s����G�z���"�D�C/>A��?�������"`t���Q�O^�>�ᾈ��l�� �����T?L@��ߩ߾�}���������=�B�>I6�>l��"B%��;8�=���w_�=l��>F�R>5`9t?���W��Q��r�>�
C?�^?&�?��b�Rj�FG@�� ��&�� Lv��?kX�>,m
?��>zϣ=�4�����_�`vC����>���>�����?��/�������"��>͂?�/>5�?cJ?�\?J�]?�-2?`�?0�>݌��|�Ǿb$'?ˏ�?"�=�VO��8S� -��B����>��<?���'�>x�?� ?��?,)H?ё'?�>�%˾��"����>�v�>��a�\��� ��>v�]?�ߡ>�^?�Sm?'ˤ=*R:��~U�L�=H�=1H>��=?�?s!?|�>e��>%š��z=���>�c?��?�Sn?��=R?Y;5>u��> ��=�^�>v	�>�?c�N?(hs?@�J?S�>��<�'������`p�&�N��jF;قA<|�}=�V���s��s��<�<{L�;�б�4�o��h�ӂG����V�;��>6r>痗��>#־|����9>�K�u��+����'�4u�=ho�>��>n�>��<��`=WB�>쀽>B[���%?�y
?��?}�R<s\�����y���>fdA?&0�=ga�<4����r���=��n?��W?>o�����V�b?W^?���2t=�{þ�nb�۽� �O?#L?T�E�K��>�~?s
r?8(�>;.e��m�4˜�Sia���h�韵=���>y���%e���>-8?��>�d>%��=��ܾl�w��֞��j?�ό?��?�?��)>��n���߿̆徔ㅿ�Pn?���>����EE5?u =g��e!����s�ߨ �Ay��޷���)��}ؾY���퉾�x�Z�=�p?�w]?U�v?M?��q{��=[���b�I�`�ߨ��!��O\�Q2���]���u�2w�ǅ��(��Z�!<�k{�GD<�$k�?^E'?�>$��p�>&��{��!qǾ��B>����@�h�=����t�<�4B=�bk��.�������?�q�>��>E:?J[]�A�>�t1�sb/���� >���>pN{>$��>�8*��:3�Aaѽ;Sɾ���ҿ���v>lnc?�~K?I�n?�A�_
1��{����!���/�]����B>|x>Ѳ�>W�W�n��4&�S>���r�����Z����	� �~=�2?R�>3��>A�??�p	�/@���Fx�<�1���<�.�>!,i?�H�>���>�(н3� �$��>�l?���>��>�Q��s!���{�W^˽]��>Yح>)��>G(p>�,,��\��^��򂎿#9�5�=\�h?W���ْ`���>-�Q?��:�@<=}�>��u��!������'���>^v?�n�=!X<>�\ž ���{�a���vM'?��>�ʫ�D�����>�?��=���>`q�?8�?��o��V%�;d�>_�g?BR?�B?.O�>�=���!����9�g�U=�Vl>r�V>�=��;= ����g,��[M�K}=��>�{���ɤ�1�=��<=��<m]��y�>0ٿ0�O��N�T�.�Tc ����j^���i��#����d���վ����4na��a,�k�n���wφ��lH�j᡾e�?h�?�'�����c��b�]��(��j?$��U�e������5���1�K0߾����;'�؎?���3���M��Y3?7���ĵ������׷��k;?�+?�p?4U��8$�i�ﾄ|��۞���j=Մƾ�,����ο�㩾^07?w�>����n^�i�>��>���>K"�>��s�����=���>��<?T2?]�d�e�Ŀۏ�����=�?�X@��E?��$��]�+�=~��>�_?�!C>�[½�F%�?���,��>��?oG{?h�<�F� ��<A�g?�����Z>���;FB�=�g�=��1�Ӱܽ��a>f�>ԹF��}�-(z��1R>8��>n��Da�7W��RY=���=���A@�5Մ?,{\��f���/��T��U>��T? +�>f:�=��,?U7H�a}Ͽ�\��*a?�0�?���?#�(?8ۿ��ؚ>��ܾ��M?_D6?���>�d&��t�ޅ�=�6�"���z���&V�~��=Y��>^�>Â,�ދ���O�J��S��=Jf��)ȿ	)��,*��t;ʪ��[�H��j\��R���<'B���
^��'�����=B�>�,h>��g>�<[>!>XR?�n?�m>ݺ�Ũ��\�$���\�=`���D��0���T��j�ְʾ8��-���N�������7(7�YkX=�4D�̍����J�7U5�+<=��_+?��>���������L�� �����=7�������;:}���?��?7���8�z_���<�qý]�h?IH�{>�4���Pz�䩘<��7=��>ә��Z�¾��+�h�^�i�)?��+?�)���~����>�r�S:�=�;?�?j虻��>��$?p>=�(���ǅ>O%/>�&�>b�?r�b>*�ƾa���(?O�u? ]@������a�>Q��������=&im>�Jv�G��w��>Q ��y�ɾ�<v�,<��=�oT?ٛ�>k���
�Q���R��<7C ���g?��?���>f^?Ru+?<b=��쾕bG��z��>��R?�}j?+�=*D	=2��z��P1?	/v?��>�Bw�U����8:�X���'?�Iq?�%?]�ɽ�m�')���g㾛a0?��v?s^�vs�����Q�V�k=�>�[�>���>��9��k�>�>?�#��G������sY4�#Þ?��@��?��;<�����=�;?g\�>�O��>ƾ�z�������q=�"�>����vev�����Q,�[�8?ݠ�?���>������I��=��`��ʵ?H~?J��������R ��v�`9��s;�G��BvH<]̽����8b�ӣ�����D���UC<���>��	@P�3��=�>y�ĽY����(п�q�]���&i�?���>�H�)J��5T��\��;F�H�G�p�{���><�L>Ѕ4�����p�]��^_��?�ڰ��ϱ>�+Y�9���n"�̽:��>��>�{�>�R׼�l���c�?���_�Ͽ�͏�� ﾽ-F?�%�?�?�/�>��)�3?���SE��b���a+?��L?�Uh?tA�<赔�K�ؽ;o?�ė���A���6�xE�#��>:d?4�>�>'��W�=`�&>��>���=���A�ֿXM���!�<�?)��?E���)?K�?��?��#�ބ��ĳ��g�"�۷l��hA?tJ=G3�j���O���>�|3?�Y����Q�_?�a�L�p�4�-���ƽ�ۡ>��0��e\�5H����KXe����@y����?9^�?S�?���� #�N6%?�>�����8Ǿ=	�<���>�(�>Y)N>TH_���u>����:��h	>���?�~�?Oj?ᕏ������U>��}?�u�>�K�?o��=A�>ͺ>斆���绥�=��=Z@%�-�?1�L? ��>�~=h�K�_�3�s;�&�@��5��s�D��!�>�m?b??���>�f�S�g�M�Aӽ��.���m��'+��	���꽹@h>;�->��=6�E��?���?Hp�5�ؿj��Hp'��54?,��>�?����t�F���;_?Yz�>�6��+���%���B�^��?�G�?9�?��׾aQ̼>=�>�I�>c�Խ����E�����7>2�B?6��D��t�o�r�>���?�@�ծ?di��	?���P��a~���� 7�H��=�7?�0�E�z>���>��=�nv�ƻ����s�ƹ�>�B�?_{�?v��>2�l?��o�e�B���1=M�>��k?�s?=>o���O�B>��?�������K�gf?��
@eu@�^?9ѿXh��t(��ݖ�.xZ>q01>c�7>�B+�pv>�/=0�+ʨ=�Z�:���>h{�>kx�>�0�>���>"�R>Gc��4'��B������M,8�I�
�{�
��������}��(����*��B�L���=n�:�?��9������=�U?\�Q?4p?� ?~tx�GW>���j=N#�\�=��>�V2?8�L?R�*?��=M���,�d��\��"/���̇��y�>|tI>�r�>�D�>	�>��9p�I>�;?>1��>C� >޵'=|���X=��N>�R�>���>fs�>E�a>��=-�������bf��rF�6 ��%�?�t��M][�3�����1���<'�9?_HC<�<���~¿e���ZD?�-��vw��a)��7S> n+?��I?�R>��Ծ/2=�=�*����ZL�=��H�Y��������z>��?��x>W>��F���	�XW�	+��a>`/?r���bؾ�[���O�AtԾ�g�=�?vc�4v6��f�������0��Z�=á?B(?VY=赯��GZ�`Os��y>�6�>�]�=�̒==�)>��O=?q;l�l=�"v��W�=�a>��?�d�=6����r�>=��Z>���=��d>�"v>�~\?�/?F�>�8����ͽq��V>n��>~>h��=�<��H`�He�>_��>Z
�<tR��{�X�iKY����>}�<X� �ofb�U]N���<ۻ4>��=K�Z��,P�ES=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��L��=}�>׫>�ξ�L��?��Ž6Ǣ�ɔ	�0)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿh�>�x�jZ��W��r�u���#=ި�>�8H?�V����O�'>��v
?�?p^򾢩��|�ȿ�{v�n��>�?M��?��m� A���@����>���?�gY?�ni>�g۾�`Z����>�@?�R?>�>+:���'�v�?�޶?ܯ�?"�U>'ۋ?�،?z�>J��="=_�`㶿� �� x=�%뺅*�>���>�����|�����1;f�'gp�B�)�!�S>'�b=���>7J9��ۉ��G�>�!�"t��Jq�V��>�^�>舚>6S?�@?��?���>�[�=.�ּiY����K?���?���k,n����<"ǜ=t�^��+?LA4?O�[��ϾV��>.�\?���?.[?Z�>f��:;���濿�m���ؕ<��K>q;�>�W�>����-K>"�Ծ�BD�䓊>�ԗ>�ţ��.ھ�/���᥻�7�>�n!?ͩ�>��=(� ?��#?Dm>q�>�F��n���E�)��>�3�>�C?Z�|?��?
���ھ3��g��n砿��Y��YU>bRy?�?/ٔ>�� !��Qѻ��+�4L�����?Erf?u��-N?�݈?@@?�A?R�e>fz�HLھ�<��淀>�1?�z�ȼ5��������|�>y��>��?r��������W>(������?g�9?2�3?D��＇�*�	��N�=�R'<Zw=w�t����=\5�>��>�Vǽe$>c>��>���b$�5?f>��,�hh$>�����Ž�U.>�<,?M�G��܃���=��r�:rD���>6GL>�����^?aa=���{�l���w��cU����?��?lj�?����b�h�m&=?��?3?R$�>�E��nr޾\��%Tw�;�x�x���>���>Jm���������=D��(�Ž�3���?-��>?�?�Ά>��>A%޾/�;���UھT�H�*fE��#9���6�H9�~����w6�HN�<�þV҈�$��>qV���>$�"?5�X>	>>�,?�R�=���>|�>:�,>�w�>;g�>��>6�*>�żq��L?g7����+�=����̾-=?nb[?.?z�F�J���Ek��?��?���?�<>�n��&2���>x��>*T����?Tt�=�^�Ł��>q¾�F��5�q紼��q>�Y�m�7�@sJ���K�δ	?��?,-�;t@ ����v�����=���?��'?L&�>RR��l�m�Y�1pR���+�&�u�&����#�s�u����Ԃ��W��
*�v`<=9�)?RN�?�p���x���\�s��<E���\>H�>&Ў>eZ�>��Y>����8��3X��^$������;�>x�v?Z k> qd?��O?f�^?6�i?�ټL�>>�ľB:?�#S�{�.>�W?��?v?,U?�c?�a?��?�K�="��sξ�I
?��G?�L? A?��I?I־ȥ��.z>�=�=y6Ͼ/Ž��>�n^�I�
������3t�I�<�V'?�3��3��*���G3>ۊQ?�?��>����&H��ߎ=���>{�?dŗ>��5E���12���>�t�?7&����=ӁT>�	
=�W���� r>����5�=Q!ȼ��� O�=x�>'#M=�}|�Y"#�豐<9��d�">H/?�#?���> ��>������\���=B��>�cx>��>xپ�y����Zx^����>Ѹ�?ꝶ?�"�=LT><��=� ����01��ĭ�� ��}8?g'?\jU?E��?l+3?P>'?F��=P���n���Y��㍾�?�!+?���>@�
�S$ϾG㨿jC0��?j?p�b�����#��5����ǽA� >q6����鮿)�A� s�<sc�/�:�8��?��?�'7���;��i� ���n����C?���>��>���>v)���d���N�J>��>!M?h�>�i?��?�YC?s�>�(h�=����������=ӱ�>��?��?���?P�?r��>��>��s�hҨ�R�ԾO���x��C����]<�F�:f�>�?�x�>�#�K�O�nmt�l��b�>��>�?L^�>|}6?��?��=�??���>�Ϻ�������p�{b�f����Fi?T]�?h3?��]=���q����s��>�"�?��?�?'����=u*���ݾS���N"�>���>bش>��=N���#,=���>7?��=#.$�'�@���C�,?�O9?��@>�w���U[�ہ�)�ξaG�.���Ԝ_��. ��P~�?P���`�&�#����䆾3]��{V��׼��p�=����?�o�=;>�>F{$��W��I���7=��=�	=_t<��J<��l��tl�{	����<�^S;�G�;�ؼP�ž]~?�L?��9?�F?�A>gE>�`����>/�*��?��g>�(��l#����3�:t����s���ƾG�׾΋L����K>
j�9y�=�R#>�V�=�!=b6�=�z�=x��=��
�~C�<��=���=S͢=Qd�=|��=S�>�;w?闁����Y%Q�(\罕�:?^�>�=��ƾ��??�?>�"��ڐ���\��?���?�I�?��?��i�kh�>L������<��=hU��f>2>`�=��2��y�>�2J>>V��G���U���+�?	w@�???�Ͽ#m/>8��=c��=I�L�H7�x�Ѿ³&��"'��;7?o*9�'�����>P�_�n1X�!˾ټ�=��=����כ�:�X�y�=��j��D�=��;>�q�>Fn9>��6<P]L��P>}E>m��>�e�>/Ľ:��T�ѽ�/�=��=�b>^]7>���>K�2?�T?�n?��>���W�`��ϸ�=�>&Me><��>��2>��=��>_s?|�=?��h?��>��=j8�>�vl>�s�����UC�Z���^�;����?k�?<�>xn4��f�����]n0�VD����?ج?D@?N�>u������� �!��R?�����	q?>Vx��jo��>d��E�������|>���>D�>���>���>��M>�ڲ>�>�	K:���<2O޽�3���
�6F����F��l�=$>(���	R=x��Im-��s�����=b5�<��;�� >�:�>ɀ>?)�>MZ=�6|�MW>Q(��^KI����=틾'2�>�Q���v���0�ӛY��W>6lk>�7>�8s���_?@�>�P�=�:�?��j?ųi>y�H�Kо�O��������;S�=̊�=�v)�_u=��%a�B�:��׾#�>Eu�>��>g�>wF���-�q�_>�`�a�O�>�����m���-��|)������B��qb��O^���P?i���^�>�}~?z1?��?��>}Zm��X<�N�>B��1�>���C�-�X���AtU?j�I?���>�=���d�}F̾"
��۷>yDI���O������0��1�@˷����>������о�"3��f��������B��Ir���>�O?�?19b��W���RO��������o?U}g?e�>dL?F@?,��t�Ps��&o�=Q�n?���?�<�?>YP�=nI�dX�>=�?�w�?��?%k?��|��O�>�pM=u�;><мf�=t��=}�=�̉=��?=Y?�?7Z�����ӿ̾��߾�]�[�<��=���>OU�>��n>av�=H��=/V�=^�l>/��>Jӓ>c�`>۩�>��F>�ᅾҋ��� ?2�L>!@�>��R?6�>ګ=��M}=.a^>�Q�=��9=/����6]<�Ą�|�*��b�<#٥�.�=$��>����@,�?�L�>7-�s�?���
�9%�>�	�=�b����>���>l��>�x�>�o�>@�=�>�>%�=y�;~e>/Z�#�~�A���M�q�ʾ�f�>kğ��Y9� ��/��,�A�g~���` �Ͻi�F^���9���;���?�a׽Q<e�"�)�����\
?��> �4?����Nq����>'�>px�>ĳ��Lܓ�̍�u�߾w��?�S�?i<c>��>��W?�?P�1��3�uZ��u�&A��e���`�k፿i���k�
�S����_?��x?�wA?n6�<1=z>Q��?��%��ҏ�d*�> /��&;��Y<=�(�>'%����`��Ӿ��þ�9��EF>��o?i%�?2Z?lRV���}<2��=h�?��P?��r?]g+?��>����1?���>,�?ꜯ>4!?!Y=?��?�C2>X?
>wq(=$dc=�Q�Y����Q*�����WH׼8� =	6z<K=�0���V�<^�=�K�����=�l.�L�+=f/�<N��=���=#٤>�hq?��?��>��??WT��<T��A���6?�:/��S���A=�����ml>q&�?Mү?��p?�ݗ>��Y�ݮK�S8=���>^l>�-
>��
?c0��Y=��'�<\�>�R';�P���x��E���+�o,��6\=�0�=#�> z>����Y&)>1��P@s��_>vO�ȯ���%P���E��[1�Gt��O�>��J?�?��=�!�t��ٸe�V�)?c6<? �J?��~?T��=�׾��9��"K��t��c�>��<�x�|��K��ID;�]j1;%Kw>񜾬��%�B>B�������x�2�<���/� >)e���<y���"�,�`��j>2K>���;��4��a̩�$K?j`ݼD}���P�̐�Lg)>���>#ڪ>Z��0�m���3�a�ž�&�=�&�>��4>���y���HI���;2�>Z#F?k
a?	ą?�(s��+r�+�?�Y������4B��Zp?z��>�m	?
�K>n.�=���S�yc��mE�Q1�>A��>O:�mD�����b����"�T��>�?D�>AZ	?l�R? �
?�6^?Q�(?s?K_�>�
�����<�%?��?�Ϡ=�ཇG��;��RF��<�>%�5?&#�_Ql>��?j?F"?*�Q?,?5�5>���W9����>ϑ�>�2Z��5��'�a>εL?	ä>
~]?��?t�I>��;�I{��]6��X�= �>җ&?��#?��?�>y��>�}{��G=Y״>�{o?R}?�Lo?��_=E�
?M�w>�R�>��s=N��>���>Y�?
�M?S#u?'^K?���>ݿn<�j�9���҈�#=��S�<`̀<O��<��X��ݼ�T�mV�|����;[�
�Â!���_��W��5&=Ж>��>e�;��?>�/'���徚jA>�(8>R�/�0�������=5>r��>���>���>2'��^L->��>�~>���p�
?O�+?�R?͸C�ܗq�O��#��� C?�ge?���=trM��V����P���6>��O?��^?��l�*����b?��]?g��=���þ��b��y�)�O?#�
?��G���>!�~?k�q?��> �e�x;n����>b���j�a�=�l�>[��d��D�>�7?7S�>��b>�'�=1d۾I�w�\r���?��?X �?���?�*>��n�//�Z��/���'�l?a%�>�+���I0?�x<��a��I��kl�?޾��ۢ������ ����ѽS�|�s������=I?�q?V<w?�/Z?h�	�2�d�15g���y���Q��R�$��_B���I��WJ���x�K�����o˜��M'=�zn���H�Q�?W>-?c˽�d	?�I��"F	�����l>�v��Kc�f�=$���<�u�=} I��A�۲��9�?��>��>;�:?�hZ�;�3�67B��E;��z�K�=�x�>Vm>-��>ۺ�m�Q��kɽ���cڃ��T�W|W>m�d?��k?3��?�E ��^7��M��-�E�oͼ�Ϗ�u�9>��>{3>k���\�FJؾܚG���y�7�Ӿh�R�<��c���W?X�>$Y>��? �>b)ž���?��̾NZѽ�D?��?#�?��>q!��P=�R��>��l?t�>���>o`��E!��|�q�˽C��>q��>��>��o>mj-�dw\�Ig�������+9�I��=��h?k}��S`��օ>��Q?'��:�C<	�>�s�3�!���I'��C>��?�U�=�;>�Bž&+���{�G���'r!?-7C?M>���7�YN�>(?�1�>5-�>�/�?6�>��@��=^#/?H�n?�U?!�7?��"?4��=�t�=u|�,�T�������>���>��=&�N>m�2�^��֓h��L�>g �<ނ��5Q1�z�>�z��o=�o�=A��==ڿ�Q�G>۾O��vݾ��
�c���Yod��'���N���ľ����:h���?��6��\!��Go�^f�SPp��H�?���?$q��SEꜿ��t���z�>e�w����"���#Žp�����о�@��[���X�"�T���h���3?�ԑ����A=���款%xX?��>?]�W?��� ������>I >H�S;���皿�zӿW5���|?���>�� �m@f�H]�>P}Q> �>�&T>i)��d���G�����?��`?���>�0��vIҿ4Ἷ���=���?�1 @�ZA?��(��쾧�S=���>��	?vA>�/������K�>=�?��?�Q=��W�����d?��)<�E���ƻ"��=[��=WR!=���I>���>v����@�\�ܽ�5>�H�>����J�a���<�_>Թн?ˏ�/Մ?{\��f���/��T��OU>��T?/+�>9�=d�,?77H�_}Ͽ�\��*a?�0�?٦�?��(?�ۿ�bؚ>x�ܾn�M?]D6?���>�d&��t���=15�����s���&V����=��>"�>��,�̋�E�O�{K�����= ��$ǿ���I�z�y=�̏���ͽ
�ǽ�����ֽ����M[���
���Ѽf=�=I�v>A��>:r>�sD>��Y??�_?˙>��x=��
��#��;�¾@R�=�|���H��å�������~�#/̾���n=��(�fYѾ�=�y�b�7�T����`���-C�4�.�(�F?�ׁ=z9�_�5����=�6�I��:�<�3n�S��7���b�_.�?t�m?���I�F�^-M�*7�<��(�:kg?}V+�~��&u���>G>�i>��[>�4Y�C$�������1���,?Q?j�˾�a��sD>��4�"�><��?��>���7;�>L��>(����.�"�u>��>>;j�>���>��<���j�ླྀ*?^�D?^vF�����5�:>����>�#�p��$+>�簽�%9�K�V>�D?��u��Ҽ9��N	>N�V?o�>�(��o�E�������Hj\= �w?z�?R>�>k?��B?�W=����R����EM=��V?�i?�q>�����Ѿإ�	!5?'f?pV>P�e��?羜l+���_d?t�m??3C���|�V���[�(8?��v?s^�vs�����;�V�c=�>�[�>���>��9��k�>�>?�#��G������wY4�#Þ?��@���?��;< �L��=�;?k\�>��O��>ƾ{������D�q=�"�>���}ev����R,�b�8?۠�?���>������!U�=����*P�?y`�?��^��h�=R�!��b��������,�<~��<��v��g�R\���<�*G�\u�=�B>w@��:�zH�>L#��٠ܿp�ӿ��$��%��#̾�?0Y>>������2��8V��&��z=U�s/+�/K��K�>�B>��2�V� ��v���N7��,"��?��>I��=ێ�e��fsk��X�=�g�>;۸>&��>��F�8���2��?X��i�ܿ,Ő��^��x�?��`?@I�?J��>B'�=��1�|P�Y`><>:?+}?�gH?�$�ZA����d�r?�[��x'���׾��0��{?��|?j�4>�o���>uu?�C<?]�|>�k����߿�K��R������?"	�?Z����>��?��?M�.��D��%i����?�RƽFq?��<�_��xu��^.���9?��?
�~��[�_?�a�G�p���-�h�ƽ�ۡ>�0��e\�yL������Xe�	���@y����?K^�?i�?���� #�g6%?�>b����8Ǿt�<���>�(�>�)N>GH_���u>����:��h	>���?�~�?Mj?���������U>
�}?�>AƄ?��=F&�>N�=�b��b�5���#>%��=jB�:�?�,M?+��>�.�=�`7�ĉ.�\E�4�Q��%���C�î�>�b?�L?��`>���^h3��� �S�ɽس2�sݼ��>��b,�߽�3>~&>>�%>XCD���Ѿ�?3p���ؿ�i���o'�64?&��>��?���E�t�X��3<_?/{�>|6��+���%��[D�f��?�G�?�?��׾]G̼0>]�>I�>1�Խ���7���{�7>	�B?��kD����o���>v��?�@�ծ?�i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?dQo���i�B>��?"������L��f?�
@u@a�^?*�ܿW�����6D��lC�������>�"	�Y��=��*>�ʥ�Ŝ<�5�=��|>��=�#>]��>ȭ0>�s>�����!��������*;V��E�m�"���S�%��$���-�1k���!Ծ\O���)����Y�+��x:��ܼ�w�=m�T?g?�H�?�R?��۽";�>�o,�kOἘ�I��G\�� �> �?��b?�4+?��u>��>��^��6c�����4�,�<a�>��3>�Y�>oy�>�J�>���9���=:pa>qp>��D>4�y>�v�=�K7<,9W>��>��>�T>P#}>
j�=����_��O�t�-���4��L�?�A��D?����4��3���I� >��<?���=l��Qο�{��;G?�g̾%���:��{�>T�?ϪU?���=�Y���8��T��=���A{�sN=|��^Qo�Q�'�6�=>�S�>�ϟ>�!�>��;��%/�;}l�љ��E�=Y�T?�Sﾁ����2�Ca�6*��Q�>O�?��=����ਿe2��9p�H�>��>?���>�.%�j�ʾ~T����#��3d> �6>���#��=qh�=)gc�{��/3�M>.z%>�X�=�?-T>���:9m>�Z����~�x�r>Ç2>.>�C?w8)?�Q)�����W�������u>���>�w>�w�<�^s�̊=��?,�p>����s�K�*�=,���G>�h�4%%��*;d��=ʭ���=�D�<<� �]�R�-D>�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿc�>k���񈿘Lg�ɢl��L>î�>0;W?��澇H�����
?q�*?����ě���ʿM]��|�>��?B�?�V�飿�R5���>|�?ýq?h�>Yɾ�Q�LB>ڔ(?ESS?�̾>Ҙ���$�Ε�>f��?�ڑ?4%>2ޑ?珛?IA? I�=����Y׿Ώ���y�����.�>7�g=yO�����
4��J���mM���Pݾ���>�o��̴>b�޽�B��j��=�������6!�kѠ>3T>��>��>Fd?�W�>ᪿ>K��>)a��Dd�sHn���J?ꖍ?���Ck��e�;ĥ�=p�_���?E�/?�����̾�"�>KoZ?e�y?�=[?�2�>�I	�`��;�������:�^8>�D�>2��>�]���`>��ݾ�?B��J�>P��>Ni<��վ������s�\��>L ?���>��=v ?�d#?�k>-t�>�UE��|���.E��D�> ��>(?��~?��?~v��b73��В�]꡿<�[�u�N>!�x??�?� �>����)���zD�\�:�y��l�?��f?j�	?=��?�@?qCA?��c>d�V�پ����΍�>�T+?�	���{m��1� ��m
�>nħ>��@?�:־��E�3>��� �W�%"?6�\?%�?q�B��&��vK�WB�+�>���=�>��м<d�.><>>����=o˛=�D�<���Y@�#�d<��W���y>j�}����VYE>�;+?j�<��H`�KF�=�Np���:�e�>�'>lDƾNjr?�����g�CM��>���w����?���?�җ?�՝�`�u��BG?�?�?C�?��?�ɾ�����ᾤ��!u|�h�)��_�=Y��>��ҽO���4���A
��}Ϗ�ap��0�sb
?	��>��>U�"?�R>���>�?־��'��_������D��A���C��#X��K�ksg���̽�)�=H����?��yԧ>�W���>�?�X�>��>+��>i`�<�gY>.w>�F�>ah�>4*�>Í7>7�\>g��<�3�g/Q?����u$���Ӿ��W�X?J-n?!?�٩�l9}�8N�V�?#S�?�̐?&�?>�%n��9�p
?��?��8�VD�>v1���m<S�i=n֊�eʉ���|�;�G�>�?��+82��?�m�F�%9?�?����k־( ���C����= ��?"[,?��&�[�N���r�v6X��jQ��z:�w�e�y����)(�ۧv�Ka��K��q���D#�O�N='?�Z�?ڠ�܏�T٧�U>k��D�uz>�7�>L��>^��>��3>L*���6�%CW���)�����a�>e�x?K�>~OX?HQ5?��F?��`?��d>,�>E�վ}�(?P$>G�>v�?0#?_6?c�4?F�0?.�E?�Hh>��l���߾��ܾ��?��?��
?m�?�`%?kg����$��>}�7>�ӽQ{��X>'4��鍽:�C���#>��">�*?z��0�b�ξmh>D�t?}$?ř�>5�n�J���@>���>Z3?w]>T��X�`��i8���>�Ԋ?��B�/���?C�=�<���=��#=���=zKP����=���=�U>�l�=)�����w=҃��(��<��]�I,��P��=�j�>Y�?蔊>mN�>�<��`� ����_O�=��X>x�R>9m>	#پ3q�����G�g��2y>{j�?�n�?T�f=QR�=���=�l��h7��J���Խ����<��?>#??T?划?��=?Vs#? �>�-��Q���d������O�?.�+?$��>a�{�ʾ%����d3��e?�?d'a�4r�G�(�����{ѽ�->'/��?~��˯���C�툻4��z՗�<l�?� �?��G���6�k��[���g���{�C?���>�,�>�\�>�)�Mg��0�7�<>v��>1)R?j��>��O?[,~? [c?��n>-8�����3������6P&>L4?�e�?�F�?m�{?l��>�:>= � ��������Ѣ��s����h=1�`>�k�>�.�>���>�:�=a���ν� ,��b�=֟p>;>�>"ը>��>�k�>k'���E?�� ?D(���"�ǻ���ɋ�܀��{Vq?�֖?�W0?��{���l2�BG쾡��>R��?,ͭ?�"?�8���=�-��I�ɾ���@�>6�>��>X�=z�+=M�>�(�>�ƭ>���;��N4�����	?�.C?�/�=(3ֿҞ��s�u��ξVB߽G���F|�����&[�/>�d����Q	�����}৾��y�6��-o���$��|�>KL=�>�n>��=TXV<W�m��t]<	0=1�F�*��ܽc�����<�^O�gە��[r<��=B����-ʾ��|?	cH?�(+?I�C?b;x>�0>r�1�a�>���Qo?=%T>��T�F⼾�,:�
��o���_b׾k�׾Wd��̟�O}>�II���>t�1>ظ�=�|�<Sb�=Wv=��=�m-�FQ=/6�=4P�=<ɫ=���=��>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>q��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>���>���=�K�|V�#��;g���Q��?�7���������>��@��)��ڢ��a�>G3X>�b=�P�f�b�w1(="���&�;,0��6\q>�eQ=�
>����i�y>=s`J>�O�>����-�e��W��<�->x��>�+�='��>�??��H?�?I��>�
��K��)4򾖥�>w�>��q�ю�>|̺>���>Fh3?J��?i�_?=Ӕ>9�<�V�>U:�>��G��ғ�+R�J���������?Gկ?��>��������!��E�U���<��?w�L?��?w4?�'��ؿP�쾴.6���ɽzs��d���y�����=-�Y����ٲ��P8>�>`>_X>N��>���=�&Y>�à>@�=�A����>�(>S�>0&�<?J4>������R�p�=4��=K0�=�����>��>_��!TļS���Ri�=O=�>�Hv>>�I)>��7��>�G�WyY����>Y
��e;�mu��&�����g�u$����a>3�}>�>>0��l�?y��>/>	��?�W?��>��/�վ����v��D㞾�Л=��]9m;½#\�qSg�Dya�W�8��>�i�>� �>N�m>��+�wS<�A,�=���5�n��>\��a�1��o�OG��&I����`��V�<i�G?����p�>�}?��E?>��?)�>�����ؾ�>A����,����_>���DŽi�?y@$?�@�>������D��H̾ ���޷>�@I�/�O���K�0�Ѫ�4ͷ���>������о]$3��g�������B��Lr�g��>�O?��?G:b��W��'UO�����(���q?�|g?0�>�J?�@?&���y�jr���v�=�n?ʳ�?D=�?�>�	�=���I��>�?�L�?^��?��t?�kH��V�>rx�<~>~x��Z�=Բ>�׋=�O�=:�?��
?-�?�������3e�c�`[\�^\=�*�=-א>�F�>k!|>j��=�Cm=���=%�f>K��>��>4{g>gƢ>^��>a���o@�	�C?��@>�*�>�:;?�D�>U����<�>gr���!�.�0�U�<����1���6>A)">%t�=���>l�ܿ��?�$�>"��yN:?����r&�]��>��;>������>�I�>���>x?��>��W=VQ�>3V=|#���>0�ܾ���V\@�b}������D�>�՗������ͩ���so��a��Z���i�1�w�z���;d=V�?�_��/h�o��ۍ�ʘ?'��>�CZ?��w��ԑ��r=k��>+��>e�޾%珿fb�����t��?p�?�3c>J�>Y�W?͛?�1�*3��sZ���u��"A��e��`��ߍ�����N�
����t�_??�x?�xA?���<�;z>��?�%�$ӏ��&�>�/�E);��U<={*�>$����`��Ӿw�þ�3�jMF>�o?!#�?�Q?CaV�`�Z���.>�:?M�2?ذu?K�-?O�:?�3#�2�!?}�>>G�?�?�2?ƞ0?�@?7�>>2��=�O%�~=���&%��˽}�н~�ż�L'=�'v=J�1:�0к�#1=H��<M!��`���<{�ݼqE�<NT=�|�=��=w��>�N|?2Q�>e+>4oI?�d#��_/��]���l?u�j>ȿ�z��ɝ�d3����Z>�xu?��?	_L?�w�>�q1�"e�j)=�[>bg>���>*
�>�/����|�=|b>E�Y=���=��=�큾a�#�Hi���y�<"8>{��>�gs>	쌽��>H��	�s���M>I>�pz��Ѽ[��8���(��Z_��@�>�F?��?>��=�J�����rf�=�?CXJ?�R?�Dz?���=2�Ѿ�8�%�A���@�Iw�>翐=�� ���\���E�5�-���~��>�C��W�����m>���ּ���\{�at_�r��!�t=@w��n/&<`-��Ӡ��%��D?�=6>�Q¾�j��Q��|@���FA?կK<�Cv��@g��Z����W>�E>�U�>�J�~	��&L��A�Ϗ*>���>:>X�+=����R��g��s>`�N?_�`?۝?	�2�3���2,�5����þ���;~o?���>���>��>N��=�a�� �����S��wO�m��>�x�>���^�'�(����
�|J�����>ٗ?y�2>v?Bz?��>:�R?O�B?ܬ#?���>�Q�`�a�\�#?�`�?ӯ=q���(W���E�V�L���>�y=?��;��d�>/�!?��?� ?��K?6�?P�L>���L5��!�>�z><�O�sF����'>�M?���>k�e?�b�?z�r>�>5�� ����ۼ�h�=IJ�='8?�@ ?i/?�q�>{G�>�b)�6p>h�>�π?�r?;��?�8�k�?7z?Q&>�D>}0:>�f?�>�:?�D�?�O&?�v!?@��h-�����!�;�4"=v=ut=��=��=	AK�-�[�;����{<]����;�]Z������kֻ��7=�A�>�0�>zz�p��=�<,���ᾒ�c>��=�?.�����{��>!��=��>�"�>>񑾁Q�=Z��>���>�����?��'?��U?�� �1V��� ��H𾍣�>1��?�z=�r`���S���>�AT?\	L?^f��[�+��b?b8]?���E<��ľ��`�J8�5_P?*
?��J�O��>�}?3�q?cc�>�Tc��)m����1b��5m�\�=e^�>zP���d��Þ>{�7?��>b�f>#�=Y2ھcIv�x~��H>?���?��?�O�?rd,>e#n���߿*�ou��+Vr?S�>1����0+?I�<C�����]�v����꾲_��}���Lü���Ǿ�XX��t���tO���=�(?-tg?�h?�a?������`���j���{�ZL��۾0*��nA�"�:�@���M�o��{�*��w�/=�1x��@�27�?g�+?�;����>�n���� �É��M�)>s��ϳ�{=��潔�\�d;�<ơh��c�E�����?��>���>�.>?o�X�{=��8�Ź8�����C>(�>-��>D��>7���t�6
���߾ȧ���۽��?>�?�JZ?�g�?$�1>�R�������8�ا�=
UP� �����=K��>�lY���C��!1����3��X*�67Z�k���&��<;M?��>�J=�3�?Ň*?�=��E��*	��u7�7>����
?`l?�`
?�U�>�r��r�O�+2�>�om?���>��>S��s�!���|�_�ҽ���>z��>
�>==p>�d*��\�J[��ㆎ�^�8��=�0h?���hWb���>=�R?:)�;�|><���>��u��� ����{*�->��?zƫ=�<>��ľG���z�^��374?��?T͇�x�4��;�>r�?(��>Uo�>m�?�>�� ���K=�P?�Fq?�C?�
J?�?�>�~Y�oӽ����aH�<O�>�?�>� �=B6�>�֐��룾�M��7W=*��=����=�@�=��u��p&<kM<ڋ>�Jۿ�;J���پ������,�D댾|������6���� ?���p�����e�X�Q�ea�{���AYi�1��?���?�ڗ�r��2ؚ���z�/=� ��>��f��N���������o|����ܾ]�����!�x�K��Qb���_��9?G��}.��F����i���%?WK+?��f?����/��1��.8>Ց�=r�6>Z �*_��?ȿk<T<t?K��>~*��3
����> �>�o�=:%m>��������.�=n�>�.M?�k�>�x4� �ҿ%ٰ�ʲX=#9�?��?+ D?��/�5��q�W=d?�>��?�X>��$��}!�QS���L�>N��?�<�?��=�\�,���6[?*�=��3�Rʻ�|�=*��=��`=�9�C�@>�/�>�-��Z8�"��S�S>SL�>�0��j��\O��|��<C�>�݊�A��+Մ?{\�xf���/��T���U>A�T?x+�>�6�=�,?7H�I}Ͽ�\��*a?�0�?ɦ�?��(?�ۿ�?ؚ>��ܾ��M?MD6?���>�d&��t����=E:Ἅi��i���&V����=«�>؅>_�,�ы�e�O��F��h��=W����Pm �w�A����=6�ν����w���/�w�c<v�H���[�F`C��5>p-�=��>�/�>�Fl>��=�O?�c?�D�>�u2=E-o<�O?��Ͼ�'�AA?����u�+��Bǽ��%��n�������޾��2� �
����3��Cz=�\�槌�&+��a>���]�Y�9?���=�R��(���2>�f�i����IG=~�������$���C����?:�"?z|��;V�z�*�f=^�ܑ}?�嗽QeG��Q���m*>�O�=h-�=��C>����徰��H<��s/?6?sW��ҍ�t	">@��K=��)?�N?�:0<QK�>�a%?/�/�L$���\>��2>���>�>��>����%ؽ��?��T?�!���.��2��>�X��ow��?q=�&>h2��Ѹ��&X>�͍<�	���W���9��$��<��W?K<�>�>�v-$���v�����P��Lt?8G?��>��%?��/?Zp�>ľ��*��Ή�Q(}>ѡ\?��[?&>_^����GB����I?�?u��>xi��� ����7	�f�>�b�?��;?Ҿ}=b��_��\����?��v?s^�xs�����U�V�b=�>�[�>���>��9��k�>�>?�#��G������zY4�#Þ?��@���?��;< �`��=�;?n\�>��O��>ƾ�z������+�q=�"�>���ev����R,�f�8?ݠ�?���>������jo�=f����Ȳ?�t�?�ȯ��?�=D���z��&Ѿڋ<]���3꠽����\�J����������c�d�=<Ju> �@u �W�>J����׿�6Ϳ�j�I$;�ν\>�>�ٍ>�7��0���q�v�_{��9B���<��R7�-X�>�W>c�6��M��끿K���l�A?	��H����t��~X��GA���;�=U��>��>J���0,M������?Ƀ3�"i������Aմ��m?�'�?f��?�k>�_�dQƽ��-KZ>��L?�j?P�S?�$�!K=�d���r?���?1�����mʊ>�_B?K��>n=*���F>�\�>��?���>�v��PWؿtq����u����?�?/�����K?f��?k4?DE�t�y��վ$UC�ʾ&>�Z�?�k�>L$��N(�L�p�#�|��>��?��57�X�_?�a��p�]�-��ƽ�ۡ>r�0��d\��F�����XXe����e?y����?^�?6�?.��� #�p6%?v�>���J9Ǿ���<‧>�(�>l+N>�B_��u>q��:��g	>���?�~�?j? ��� ���6W>$�}?s�>v.�?���=�~�>:ո=���\N���>��>Z�m�8��>��J?�`�>\��="����*�?�H���U�ײ�QB���>��`?�S?3�g>Ys��G��Y~ ���ؽ�A5����<S�.�"ꉼ+=�-�>�k7>e>�sE�G�о.�?�\�N�ؿ;q��*�'��'4?=t�>y?z��:�u�/��\_?a��>\!�����#��R�ڎ�?06�?��?��׾��μo�>��>5ރ>Oӽ���b��<8>ӈB?-���Q��B�o���>s��?H�@�Ǯ?fi��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?�Qo���j�B>��?"������L��f?�
@u@a�^?*����g˾Y��E�<�����|@>,�{>X�=�8�K8��]��<{�7>�&2>�r>O�`>���=�N�=zՅ���!�����r����-��b�o[�q�<���e�}����-�BM�WR������Cn�W��r�-�D�N���=��U?MQ?��p?)* ?>M��i>�A���=2�$�~Q�=j��>e�0?�XK?K*?�C�=,�����d�w-���G���r����>��K>l��>���>�B�>ke%;G�G>-!>>u>�O>:-6=zǺ��
=�O>g!�>���>AM�>�D�>�漩��E��� �����O�X�I��?%y���c��7�{��]���F�*N?�&3>a[����Կ�ƿXSJ?d���n揾׷�>�l8?�|??��>ҾBR�=}�S>l�����^W=��;b�i;��$���r<g�?�?�>:��=g�5�	v7��f���� ��=q�=?Z
��[�3�^�#xC��0�?��>"Z�>c��=��7������^�oش�V��>B3R?�u!?K�۽#����cx���ܾx��>�e�=A2���w�>�˷<5�ҽƨ^���\�TJ�=�"�=��p>�x?�->���=�֤>,H��$Y�y��>1�?>ü,>-S>?�r#?��5ܨ�G��� *�L�s>-��>�S~>��>�+K�4B�=z�>>?d>e��z8��LV��*@��	U>�f�\�Z�G��y5�=��)A�=���=�+��|@�FF=��~?�å��t����p`��R�C?�b?���=8��;�!�ͫ�������N�?_3@\��?V���7W�O#?T�?Փu���]=!
�>(v�>����2K�*/?���^��������V'���?�K�? �P�����4q�O
�=��*?�`���&�>���h����u���&u�5�0=�V�>��H?��O�a���<���
?�.?���;̣��Nȿ��u���>w�?s�?_�n��W���@�x�>e��?�SZ?�)n>��۾0�W�{��>
�>?�:Q?1�>[��-�^�?��?�ԅ?���=�.�?�g�?"l�>ow��s�5��h��"ĝ��r�=���>z�7���S=��L�ʃ��ߪ�ƣ��1�o�䌾��>���<Ł�>Іe���^�n�4>8�~��q޾�Y�����>S6�>��>���>	�>0�>�6?c(2>��;4�o�/?Ծ^�K?_��?%��R2n��F�<]��=!�^��&?_I4?z[���ϾLը>U�\?6?�[?%d�>Z��J>��迿~�����<��K>d4�>�H�>�%��)EK>��Ծ5D�)p�>ї>
���?ھ^-���T���B�>�e!?���>RѮ=,b?�$?Eo>I��>��A�����Z.F��2�>��>^e�>��?�?/���3�F���{��ĖO��TA>�-k?�=#?,�f>x ��;R��0�7<]:�;I*=0ʊ?�l?�×�l�>�]�?�.T?�\?�5n>سD��{� i�=Ƽ>XcB?@�++\��6��p���?��V>��v?�@���.>9?�S�hx����z>��h?�D?�nD�,����A�8I�<1%=��'=�2��qdl�oK>��"� �ˊ�=���=��'e���e��/�<q����=��=@;ּ<L)>\�(?��/=�vb�A'>yNo��>��Gl>^Y�=�J��{�r?X�轶}p��`��\Z�����e^e?!9�?7c�?_��<�F{���O?	�?PI?E�?�\羇S׾d���������b���3�a��=���>ի��m:������Z奿�䍿��Z�SmA���?�J�>�Q?��?C)$>��>s������þ�T�Y~`���C��|R�IrK���%��I��6����w=<9¾�?����>��ٽ؂�>J�2?k��>Ι�>�s?&�D���>J�p>��w>�E�>E�.>Ք~>v�=yҬ��T�I?Tڵ�"�/�HF ������n;?SLN?1
?gҼm͋����d�)?���?�Ϛ?�]>��g���'��y?�.?��,��1�>�U>�~: =�	���%Ҿ\�껮��N���OS�>����.�R�Y�6I�<�>��>�%D��{���
޽L�����=�U�?0�F?,O%�!$%���o�3g��.����&žM���A1#��ށ�U����D��
u��&��&�>�t?��?-�����]ꁾYn��N��y�>9�>�-�>um�>g$>�/Ҿ��0��ń�[�2��9m��'�>��u?�S�>��4?��?��?��_?[+�>��?��ž���>W4�>2���LL�>�~:?�n3?��,?ԭ.?U?D��>i�<�%�ξXK?(T?	0�>���>/��>s)��%��I�_<��];T�x��џ�>��<WS�j�ͽ%�ɽ����i+>�_?���í8�������j>�y7?Ye�>��>�4��K��^��<~��>ڨ
??S�>����Ocr��n�-�>��?����=��)>���=�'��ʵҺ�?�={\üD��=�e��;�;�9- <Je�=c:�=A눻�^ṡ�;+~�;g�<���>�??��>?h�>E��T@��C���ѡ=1U>�GE>@'>��Ӿ�G��K�����e���v>0%�?1I�?�?I=���=L��=s`���̸����×���8�<`?6&?rxT?�?�@?�((?��>������a�����6P?ā+?ݫ�>�/��Ⱦu ���_4�P*?��?��_���(��˿���/�>U.��y}�4��F�C���׻���������?4Ý?Zv6���6��p�˪��8���
D?a��>�>�>���>�&)��f���m�8>"V�>^P?�p�>�nQ?~{?C�]?��V>z�8�ŀ��:������J>">� >?.]�?}9�?��t?	��>B�>_�(�0L߾����2���~��Ƅ�J�=�`>�$�>�t�>���>���=W�ýlܮ�,+2��C�=5Ff>7��>X*�>��>�(}>�~�<}yH?��?}Ɣ����წ����L�w?;@�?�I5?b\��î����/�����e�>��?2��?=d2?����0>�K�������޾�W�>�?;m�>;��=��<Y�t>���>�ga>[�m��f���rB�Mg��ų?c�I?��*>66ʿo�h��ㆾ _���N=�u���^����ʖ��0V�=�bQ�4���Ȥ��&J��m��r�b©�ޱ��_g��p?�|>.>$��=����U"�<Z����>�_�>���o^ڼ:W�=�J�="��U�����;�ʀ��D�=�	G=�Ǿ�Y|?!�D?�n-?1m>?��s>Ә>��5��ؙ>�����?r�Y>	������l�-������`��Y�߾��־��]�󢞾�>R"���>�..>2T�=�9�<��=h.==���=@����F^==*�=@ؙ=�8�=�C�=Sl>��>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>q��=w�2�T��>��J>���K��D����4�?��@��??�ዿТϿ6a/>�p�>��<T�F�}S.��ɀ��w��i��4/?T�L���
�?Ỵ=x�־�_�Yh$>���>���\���]���M=�ؼ�**=!\=S�,>(�>l�B<Tｵ�=�N=g���8�>@r����;�"
�U5��d��=fU>��>���>';3?�2?��?�]�>8r4�3%�����?*��=iڙ>���>,J>x�>��=?=SO?lxb?H�>�4���>H��>1J=�{Č�j8<�������=��(�?Ē�?竧>����'��Ⱦ��s��6��lT�?�Fc?�6/?�??�i���������8�jK=��X���[�� f�(7�=y$��%O���=�{�>d�>ۈ>�ۂ>z"B>�W�=,��>ٳ_>�g#=w��=i`0=a��=�秽�k�<��佸̐�t�=h�=l��;��Xw+=!��=�땽C�?=ڀ�=��=��?}�n>!��>�>�Ӿ;�R>t�ξ�>Y�80t>j!ʾ�^=�^�s�������L�y�����>8��>�d=`ٜ��c?w��>�E>��?u[?p��>غĽ��ľr��v�վ�yz��M#��=���d
������]��p�A]�>N}�>�9�>Cw�>�31��}?��Ճ=��p�.��3�>7v��E,���1�[�n��i��w֠��P���}=g^F?O����(>��?�QG?�ΐ?0%�> Ͻ��@ >��f�k���h��[��M�彋� ?�� ?���>��� �M�=F̾#��J۷> 9I���O�]�����0�in�ʷ����>�����оw#3�1g��;���o�B��Sr���>Q�O?.�?,?b�]W���TO�3��%���r?ag?��>�G?Q@?�.��Br�n���l�=l�n?��?�<�?#�
>��=^�����>_1?-�?��?��|?�Z����>��= ��=_&z����=}�/>T �=(x>��?�Y?�?֨������΢߾��R��!==��=���>��>O�d>y0�=J�<=��=�_>�ݔ>��~>t`>O��>ڷ�>+8���eᾃvD?��d>��>�SE?���>c�ս�@�<��J���,��3������a�Z��ɭ佰� ='d0>�&�=���>9�п$r�?� X>��A�B/?�C�3��ѓ>�]�I�ɼ��>�d�>^E]>�e�>YX�>[�4=Ţ&>�E�;:�ݾ�?�=&���,/�tP>�M�6������q�>I����'��ܤ������'Q����E��ZZ�xdq���*��Y=[љ?v$Ž�����8��Ws�>� ?��>d�T?L}F��;}���\=��?q�>�3۾jU��3瑿0 ׾r��?v��?�;c>��>y�W?y�?��1��3��uZ�:�u�-(A��e�O�`�n፿����
�z	����_?��x?yA?�R�<�9z>P��?��%��ҏ��)�>�/� ';��@<=.+�>N)����`��Ӿ%�þ�7�HF>�o?%�?6Y?�RV��&,����=}D5?FM
?`�?�[A?W$�?����� ?v�
?��V>���>a5?z�A?�7�>$j�>��>L#=?:�>�(���̅��Ԅ�����d���J�J�4
=3��<1/=��Լ��P>�J=��<{�L��)�=Y�`��= x�=��=̧>7�]?��>�Ą>{	5?4��58�Yެ��0?�!?=���ㅾ��������|>�2j?D=�?�<W?&�a>@�H�A�4C>�l�>z�/>y�j>�в>�����?��=��>C>3O�=C�[{����iˑ��S=�(>@P�>���>ci��*�+>�tپB�W��ک=�9�!���u���@)����^��tʌ>�D7?��?���:�*�a�#�c`k�A.3?i�G?�;v?],t?�C�9����Y��7�� ½���>��H>Q��������C�C���=�f�>b�������rp>nȾ
׾
.��Hp�^���=�k�Q��=*���[���˾ ��CK�>�"���E�љ���ڧ��5;?9m4<rK:�:���<ʽgZ[>�_J=B�>�u���c�N��0?���=���>�)>P�S=/v���p���8�e6�>�OE?c__?�h�?�
��~�r�i�B������8���sü	?0(�>q?�BB>q3�=$���O����d��F����>�c�>�����G�A(������$����>�.?�c>�?�R?��
?}u`?�*?=Q?�5�>�������e&?A��?�B�=����B;�+�4�D J����><5?M�=��i�>!?�?'�"?_�P?^?O�9>4��>s/��$�>
ڐ>��P������~>_QR?���>��Z?΃?jv>T~:�J����<���>Bt�=�*?G.?(�?���>��>m���ϐ�=���>��c?�o�?~�E?�">q�?�.d>|�?���0d>�@?³0?*�4?�H?��-?�� ?Wx�=�t���%����;��>=w����TP=��?=)�Y= 3<a�>���L�>y��=�����/��5��3�=м�>��>:�Z�δ�>������Ͼ�*p>�h�=`0�^�O3���>`a�=\j�>�\�>9��3#> \�>0��>�c��n&?�L$?s�>�U���g������.����>,�G?<HM>`Ƀ�xx�9`u�;�=�a?O�I?��A��k8���b?��]?ci�+=���þ�b�=�龯�O?&�
?D�G�o�>Z�~?0�q?͵�>U�e��8n���`Cb�p�j�]Ҷ=�r�>�X�p�d��>�>s�7?�M�>!�b>�!�=yw۾w�w�7t��?�?�?���?�#*>T�n�4�OkϾ.葿�fL?���>2���ZE?�R>�f϶���R�tՐ�r������A�e��*���cx�d���`���:�)�<>�Z�>��?��x?�JE?+�����d���g����4�G���;�X'L���[�UFU������$�O6��j���͖=%����@����?��&?� =�s�>*��4̾s/H>㡾�����=}���YX=�O=1oc�%0��l���"?�-�>Y�>MS;?��X�n=>��`3�K�7�	���Q-7>h��>��>���>
�;�!(�%�ݽ=QɾG4�������>�On?��d?A�{?KL;=1� �����?VR��<�=�Fa��d�>_µ=���>�`�ِ
��5���1�q'a�=�㾏Uy�h[#��u�.$W?��>�(�=Kگ?a�+?0%�����S�����OA>�߸>�t�?�].?ꠎ>:.<�����>��l?B��>��>�����T!���{���ʽb"�>�߭>���>m�o>�,�� \�l��؅���9�Bg�=�h?p�����`��܅>eR?`�:H<z�>?�v��!��򾺵'��>�}?���=W�;>oyž� ��{��8���N&?)&?�G��w�!���>�"?��>�>lA�?4�>���.�w�?`^?%	I?_�<?3=�>��x=l"�������!��=���>ƚ_>�X=B��=��'][�2��V*=��=b5Z�v$����;?uټP	h<�-�<��1>S�Ϳ)dS�%������1#�m�������=k�ϾR?���R��e��� Q�����Q��=�|��2賽 �b� -�Z��?� @w� �Fp�Ї���q���ξ%��>V��;(���x��TDݽ9>����B�����(�����<N�[{j�X�'?r����ǿ밡��:ܾ-! ?�A ?�y?��B�"���8��� >pB�<�+����뾨����ο������^?��>��.�����>���>�X>�Hq>����螾�3�<��?+�-?���>[�r�4�ɿ[���z��<���?0�@OE?���r��3�v�^7�>���>R�>4t�N2�W�����>���?r�?J��euN���=�a?x�)=/�G���<�h�=����ռ��ڽOp>��}>�U,��:z��6��5WS>5�s>�i���X�)���p!=�P=�-��<�5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?$�(?:ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=�6����{���&V�{��=Y��>a�>Ƃ,������O��I��Y��=iX���п�%�0����<�=Y�+<�?>�~�;���'����<,��ͽiO =�>��U>�C�>/;g>�>@`?>ch??߱>�M>m20��G���Ҿh�d���*'ս	4��P��k頾�j��žf�
���p���۾W�&���=
�4�9���s�)�E�d�[9���(?�*3�H�㾇(?����=m�ѾY�ɾ�J=*�<��ľ�V=�< ��%��?{�#?<�~��^��̾i|�=�VO���M?����(�)������(>>b&=j� ��:>j� >D(��A&��pl���?�+�>�琾�S�����>��5�w�<p.?���>Zb��u>R�M?���T��=�ea>4�=�j�>Ҝ
?D�`>4���?�r��>�$K?^��z>���V�>dD�� D��h�x�O��=� ����=}'>F� >B�ܾ�t�=c�p���>�@D?]�u>�9?���p����w2�^�>�ib?Ro�>�}h>�@F?�E?4�<w%��]M��R��N�>�OY?�8?<��=�S}���|��M6?�V]?�{�=�ͽdr��`&@����`��>۸`?�.?����q���*���ݱ�ј<?��v?hr^�[s�������V�K<�>�\�>���>��9�0k�>��>?�#��G��׺��WY4�Þ?e�@��?��;<���=�:?�[�>��O��>ƾr{��]���a�q=G!�>����ev�����P,�{�8?��?^��>Ǔ��թ��$>�����?��z?ew��;!>M�<�I}�
��������;�Z���k�+,�r�V��#�u�#�ɾ�>��p>��@�l>���>�_�02ݿ��ӿ�q���H���X�
�?�j=&�T���d�����{���I�b���:����߼>n�@>��������
n�$�?��0>�H�>��u�=��>�L?���l���O����@�Q>���>+��>�? =�8�|E�?��~�ѿ0���>dԾ�Q?���?�,X?��X>������v��=奦=���>�7'?�{?Io��ş���)��j?�_��tU`��4�jHE��U>�"3?�B�>N�-�ұ|=�>���>g>�#/�t�Ŀ�ٶ�&���\��?܉�?�o���>o��?ls+?�i�8���[����*���+��<A?�2>���=�!�<0=�DҒ���
?9~0?�z�Y.���_?Қa�i�p�:�-���ƽZޡ>(�0��e\�;#�����gWe�<���<y�~��?^�?�?��� #��6%?��>֝��D9Ǿ��<���>�(�>�)N>#J_�g�u>���:��m	>��?Y~�?{j?;��������U>3�}?�$�>9�?x�=at�>sf�=��}*,�%~#>GU�="�?�-�?#�M?`0�>ƌ�=�8�7$/��NF�!6R����C���>��a?܀L?	b>w]��e�1��
!��ͽb1�L�缩�@���+���Z,5>��=>7>��D�w!Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ha~����7�'��=��7?�0�t�z>���>�=�nv�ӻ��N�s�ƹ�>�B�?�{�?���>�l?��o�h�B���1=0M�>Ɯk?�s?Vo����B>��?�������	L��f?	�
@su@A�^?#;J�&G���t��+�3��@��=(�P>,�[�E�,>��^>�0<Q-=�$I>,*�>�"�>��=>R,7>�HG>U��>�>������U��ӥ�w}�ӗ.������:M���ݽ��Ԇ��Z�y�
��-�,�ۈ�8D��D�C�'�=N
�=V?BlR?�|j?2A�>�r���.4>\�"-�<�
�C�>2v`>e6?��P?#`"?CP=|��-;f��'|�썱����J�>P!,>���>��>`��>��<}6j>1>֮�>׳�=�9=u���B=3N>i�>���>���>
B6>Z;>�ԥ�񰿼d��Ѕ����E`�?>�׾��U�q1�� ��,:��:
]��?d�J>�͊�ر˿�Զ�'�I?�Ϛ�!-���c�3*6>��4?<a?��:>(�ƾ������=
�	�!�J��N���Z�?���Hf#��o>^�?Y��>�Φ>!�=��6�W�V"��݄�>�t?$rɾ;����_�I�W� ���>ܽ�>OT�Ґ6��z���h}���i����=�G?7?���~����l��S����a>~N�>��{/'�ϸ@>��>�oK�݄�MIۼ��ݽ�4�>���>9h1>	�=��>Bh��L:����>��W>_[1>�k5?�x$?���u�
�E��3���c>�>/z�>�>g�<��(�= ��>9�P>9�����t��6�vJ'�fN>[Y��g�����WL�<o����I>���=����F<�Uir:�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��L��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�0)#�jS�?��?��/�Zʋ�=l�6>�^%?��ӾMh�>ux��Z�������u��#=Q��>�8H?�V���O��>��v
?�?�^�੤���ȿ |v����>Q�?���?`�m��A���@����>5��?�gY?�oi>�g۾K`Z����>ͻ@?�R?�>�9���'�l�? ߶?կ�?�sd>�c�?e�?s��>/�R>����Lؿ����R*7=-��<dT?�&��Hw�A������S宿�x��#���>X=x��>�4ǽS;�VCM=�6\=vU̾�:��>O��>A�
?�;?��?��>�n�>M��=�z�=1�D�������K?���?����2n��;�<&��=�^��%?bH4?��[���Ͼ�Ҩ>۹\?���?�[?<c�>��v>�� 迿~�����<��K>4�>�F�>�$��IFK>�Ծ(3D��p�>{Η>���f>ھ�)��1���@�>�d!?G��>pݮ=̙ ?Ȝ#?��j>)�>aE��9����E�d��>Ԣ�>I? �~?d�?JԹ�QZ3�����桿�[��<N>I�x?V?�ɕ>b�������tE��AI���9��?�sg?dO彛?+2�? �??�A?S(f>���IؾĪ��(�> 44?���oV���,���7��>p�?�m�>1�,�Ӵ��?Ό<}z�C����>_�Y?n�?�W)��^�]��=ƥ<\iN=-�d�ENs=�$��{{@>�
�=���H�=�=��`<���E)���>zK>�p;=iDӼf߾'1ʼ,2,?�F�?Ճ��ט=��r���D�#�>�PL>e ���^?��=���{���Wx����T����?��?Ed�?�5����h�z=?��?�?�)�>fP��)�޾H��!Lw�o`x�%m��>^��>>Wk����A���Օ��pL��siƽT����?L��>�?Ǌ�>V׊>�,�>�L��#�	����8Ⱦ��b� �t���-�"�"�����5d�D��[f߾+U��3S�>Nzڽ�w�>�U?v�E> �>ˍ�>mZ��ŭ�>I�>r��>�j�>�f>�$>s�g>��=�����Q?�\��bt'�:%�AP���"A?@�c?�&�>�4l������ڐ?+2�?9S�?�^s>2h���*��?���>����	?7=F=3���ê<C���>�H��������>��ѽ�:��`M�Yj���
?�v?˱��̾�wԽ�����2o=O�?f�(?*�)��Q��o���W�.S����8h�as����$�m�p��폿�`��*%��_�(���*=��*?��?L�����%���'k�>?�8Kf>� �>�%�>Z�>�cI>:�	�&�1��^��O'�����+N�>�W{?�>�=?X�D?�l?�aX?`�>�8>�i��"-?��&>���>�a�>�rc?�a-?%4$?��?��!?�l>��=^�뾚���@�>?�?�/?F�+?w�~�sd(���>�'=C␾g�=� >e�d=;�:�}@t����G�`>-X�>\�Խ���A�����>ϊ�>�X�>��?�f�����y��P�>��>Q?�'��tV�b���a?�RV?�oM��TD<oܬ>��̻8�E>��?>�a=��~��ŧ=�܄=�'�="$�T�-������>j�d>�C�� /V<���=S�>�?t �>y�>f�����1��=A.W>�=Q>�>�Pվ&�������g�!�z>ͮ�?���?`?Y=� �=v^�=[��(������^��@W�<Z�?y#?T?���?�&=?� #?��
>�M������������?�;?e��>y~��Eó�����S=���"?��q>=�P�şW�9�/�������is>�!4� po��Ŀ:�|����;4a�6[����?8�?�EK�Za�g�ľ����'����m?���>C��>+��>���eCx����\l4>0�>��n?y��>L	C?�:�?���?k��>��
�
�������[��=�ڬ>�jK?U?�!�?^xh? ��>ާ>d�D��ھ����&��D6��܏��>,��=j�S>Y�?�G�>&_�=z.�0���es4����=��h>�?���>Nb�>�O>��=�>G?��>0���x�
�}��������R��p? ь?e�-?R�=��K	?�]_����>f�?�L�? j+?!�]��>w��Q�Ǿ�ܐ��V�>�ݺ>��>�x�=�.$<}�>���>2��>������6��oo���	?��;?ˀ�=�/˿2y�mf��"l���d0�Y��� g�i����&A��S�=Wϔ�|�#�VM��o�H�,>��j*�������9R����>�f=H^	>�?�=K5<{,)�D���B�9=�]�<�/=�w��+=O'�4L�M�����ֻ^�<26e=ڨ�:�ʾ��|?�I?�:+?D?��y>�<>��+�ʗ�>V|��T?�T>�_�㑻�6�9�>u��>�9�־*F־��b�%D����>�jA�ÿ>��1>��=��<���=��q=a��=~x(���=�u�=O��=��=��=�b>b�>H7w?|���ﲝ��5Q��`�V�:?�?�>�y�=��ƾ�@?@�>>/�������d�++?{��?�P�?��?.�i�e�>��������uq�=G����G2>)��=�2���>"�J>J���K��Ѭ���0�?Ņ@.�??�䋿O�Ͽ`J/>�1�>���<|6:���0�%��Y���p�=ŝ+?�tm�~�0�����W�?��)�݌u�����c/?�Uu=����%�����;=2�/;sB��c>�>4�<BS?>`��9m�>K�]=��>^�=[�ս��I>g�T���
�0�[>�ߵ>���>�B�>w�?
e@?	��?�.�> ����R��=�ܾ�??��>w��>e�&����>L.�>��i?�;C?�'@?�-�>�pN>�G�>�k�>!���=�����������+��͔?h�z?�(�=��3�$��8-�wR0��9F���?҄Q?�8?7Y�>��_���QG�p%e�J�����<y��<b�<��<|&2>�]���P��z�>"E�>�;�>�e>\�>Q�x>��>���>j/���9��_>��=)>��=��K>VԆ��/�<�g�.��=-M�[�8��޷;�ō=�7�=���=9�w��B�=e��>æ>ڳ�>J�=Kﳾ��0>����L����=ݝ����A�d�NO~��.�h4�z�A>X>j��p�����?.aX>�'?>)K�?�2u?�>����վ/v����d��-U�\��=��>UB;�H�;���`��@N�t ӾV]�>�H�>���>��~>�,/�I��ɒ6>�E�]/��6?�\�/��(|�T7�����ˊ���i�J�]�e�6?����y�=�x?#82?�ޒ?j�?Ӏl��i��$70>��Dߞ>(�}��9���;C"?�S?�>?�*��}=�!H̾����ݷ>z?I��O���Ȯ0���ͷ�t��>w����о$3��g��4�����B�kHr�J��>δO?2�?�5b�W���TO�`���.��}q?b{g?	�>MK?@?�#���y��r��]t�=��n?(��?v<�?O >\�=quĽo�>��?zI�?v�?��b?��D�i��>�U=Љu>��#�A�#>�O>�s>�L�=ȯ?1��>-.
?����e��K��*׾A\*�u�=�dJ=^%�>o̎>+Ot>'S�=���=ƷM=N�K>7C�>��>XM>��>D�>Ay�������?Ԇ�=vr�>�&l?{@>Z� �u�=�{u=�^}>־��|K�=�6=�W�=�U�y/�=[D�����=�h�>9׿a�X?kҨ>ͅY��?������>%[">u/>F	پ�X	?�s�=�GD���?�J�>2M�=��>Hħ>�FӾ<>����d!��,C�]�R���Ѿ�}z>4���o
&�����u��lBI��n��Kg�Pj�:.��u<=�<��<*H�?<����k�9�)�{�����?�[�>�6?ی�q�� �>��>4ȍ>_K��v���ȍ�hᾚ�?���?�9c>��>��W?��?��1�'3�'rZ�Ȫu��#A��e�H�`�5���l�����
��x�_?h�x?yA?N5�<�9z>ѡ�?Y�%�uُ�a(�>n/�?%;�n-<=�%�>����`�&�Ӿh�þe6�JAF>��o?$�?U?3eV��.�v�>X%;?m�<?��s?�0?�f2?�c,�$�%?\�t>�E	?�+ ?�8?w,/?�:?� D>���=��$�=���<���oFԽ�l���!<����<(Y�=��<�[ļm|=T	=�ʼ]J��i�<VU�<��<c�<=k!=2O�=E��>�'_?�%	?�y�>�RH?�W"��H�G��=_?��<�Ԯ�^�����	�\����{>�j?*�?��R?���>wJG�8��!>'>��>��>�
�>g��E6�1ߋ=۷�=��b���D><1�=���H}����z�����'>ܻ�>��x>=W����(>�,��y�u���c>��P�I���ZS���G���1�t����>�L?��?q�=��龱H����e��)?�<?^M?��?��=*�۾��9���J�#�����>���<9X	��֢��H���:�hN�g�r>#���������>&X�� ���d���m4z������2>z���S�%P+�O���2��+R.��;^>�澵r����@���R?��J�����!Fc��<��=H�+>�3�>�1��e��uV,���
��wL>l�?F�H=�>���H�Z�K��o��b�>�BF?
�`?S3�?�����nq��"E��� �+�0	ؼO�?��>[�?n]>>fu�=z������d���E�OX�>{:�>�G���D��0��$�g"�
�>��?s�> �?S?��?�e_?(�*?�x?�N�>@}���V��m,!?M�?6�:=},�D�N�S�;�=6��	�>%k?�$W��ݠ>�!?+�?�?�KV?�'?_�=6���G�غ�>�b>q�\�����"T>��N?2ȹ>�`?#w{?LF>W�8���S��Ā�9��<h�>��-?��.?"6 ?�I�>�G�>\
`���&>�.�>d�r?k��?6(c?�T>K�M?���v ,?�u���>��?��?�U?o|?��K?�*?6`2���x�TTG�ǆ�>7;�/�ܽ�Q�<4�&�3�Ⱥ:��<��d=��z��#��xo����0�+����:�R�=�Z;jZ�>�u>����؋4>��ľ{���ry<>�x��컗��E��l�0�ex�=��w>&?�w�>Nl&��;�=@��>�>�����'?L�?�?��Y;�wc�Yپ�P�*��>�5B?*��=6l�����!v�47^=�:p?��[?�zN�B��	�b?:�]?�c�=���þ�b�}龗�O?w�
?d�G�z�>�~?}�q?��>��e�*n����$5b���j��=~`�>`V�T�d��7�>��7?�N�>N�b>�8�=�s۾��w��k��.?��?���?��?|�)>q�n�M4࿳�۾���gS`?K��>��H���+?qü����L�j������׾� �� F�1ڮ���x���J�,K`����Z>L��>A��?)�|?�^?����u�⥄�焈��CF��C���.��-Y���M�r%]�����yK��ᾶ������<ĕj�H�U�3��?5$?uL�4� ?�ǐ��Ҿ�빾pi�>-��t�ս|�>[&�g��=�Y�=��c�� 4�h����!?	W�>�P�>+MC?�{E���G�`X?��))�B�9�?>�^>ؖ>���>�z����F����;2���g��>���L>��o?�c?�	�?�\E=�M����� �=���=���2�>R9<>�P�>So���`L���)�E��}a_���Ⱦ�J��b� �S��ײh?>)�>���>�ǰ?�[?�ː��J;����.��%�>��>�u?�Y?y�>���=�x̾���>6�l?���>��>����V!���{�[˽K3�>�ح>��>��o>f�,��\��j��Q���y9����=h?�}����`�[؅>�Q?Su:�I<�u�>�|v���!����z�'��&>)?k��=E�;>�tžx!�B�{��;����(?2�?Z吾��)���>��"?T-�>X�>S�?ɗ�>��¾��%9lE?k�^?�J?�+A?��>� =�髽X�Ƚ>&�� &=��>H�Y>SXg="+�=���mZ����7�9=�=Fużn;��jq�;I�ȼ��:<
I�<�2>]�ۿ/�U���۾��!�:��*�� F��� >Iy۾�ę��{ϾB�@���H�sS��=�<C����/�"ko���x�|� @7�?2FT�v�%�M���5���o�Z��.�>�d����3=b� ��Yw��ľ�4��ݾ�y����@/n��V��3`5?$i�!+��̃���'Ⱦ��?^6?�w?9�V9���=����=C�>��<����*��V;˿,����]??;��>��̾��|�>� >��>>��9>g���*;��FY����>}@?��?����iƿ�㵿���ѡ�?OS@�A?3(���d>Q=/�>31?�A>�g.�����g�����>?��?��?*y.=��W�M����He?e-_<B�F�����c��=���=��=�y��QI>[�>����>��ٽ�3>V��>j"�C���:_���<G�]>�=ҽ(���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�ޅ�=r6�򉤻{���&V�}��=[��>b�>,������O��I��U��=�X��տ�#���,��*=r�x<���\�;��ڽ)���9����+�����C�˻��>>c�.>�.�>�;b>#̌>�4m?%xk?�N�>�>���x����>�>=Z�{!�����.ݫ�&��~��rK�����/-*��?
�XD��%�0��=�z=�:5����D��']�����3?c_W=�[ƾ8�E���!>_{Ծ��;��<���栾�M�z�h�=��?�<,?¨f���D���'���Ѽ��O���8?U��ھ/X��+�0=E�Q%p=��>l�'=C�޾[�`�kc��&?���>p#�w&����"> ���3��M)?���>e7H>\p�>�K?9��3Aj=��R���>�-"?TM?�Pz>c�ؾr/��?�?Q�]��ƃ���=����Up;����=�ۆ>X����eD����>JU�={����	h=������>p:R?���>��#�35�!Ց��u���H3=R:m?��?A��>x<`?�A?��<�ܾiI�&�/<=SL^?K�Y?G>kƽ8�Ǿ̾�?�e?�D>Р@��` ���3��N�~$?��i?#�?��=��t��1�������!?�v?�^����)����U��?�>��>���>>�9�o��>��=?g�����ÿ�w4���?=q@cf�?A�(<Oc"�̣�=f ?���>?PO��ƾ
����X����u=���>=���j%v�N���(��Z8?�a�?��>s`��&���=�=N�S�1�?'k�?�MC��v=��@�B]k�#��Y>=�U˼ut���μ��\�1�����ҡ�?'�=nzJ>k@��>�>�1�)6ؿ�bѿ����X��[���}��>��=��u��1{��Z��=��|sZ���4�W��$��>��>��� ���� x��;���_�?�>r�@�^Wx>�#C�%2�������0<Ś�>��>%�s>:;P��]���f�?u����Oȿ^'������`]?n%�?|Ճ?��?j+�A	��J�_���H�pz<?��r?gjN?����
��_��j?Vħ���_��3��D��S>��1?��>s�*���k=�;>��>̀>�2.��ſ�Ƕ��� �gB�?���?��쾥)�>��?�.?n��.䙿'����.��b�D?TW:>3޽��h&�U>�B����e
?F�/?�
�7�e�_?	�a�;�p���-�7�ƽ�ۡ>��0�qe\��Q��)���Xe�����@y����?$^�?P�?`��� #�,6%?4�>?����8Ǿ��<逧>�(�>:)N>�F_�t�u>����:�Jh	>���?�~�?j?𕏿����V>	�}?	��>��?��=R��>��=e.��U��� >X��=��H�d�?�RL?���>ת�=I43��z.�hxF�ƛR��	�hD�	�>�Ab?�5K?��g>��x�*�
� ��xȽ��2������8�/�(��*ܽ�5>U�C>\�>��8���Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ua~����7�o��=��7?�0��z>���>��=�nv�޻��V�s����>�B�?�{�?��>!�l?��o�P�B���1=9M�>̜k?�s?�Qo���i�B>��?!������L��f?
�
@~u@b�^?)Zhֿ����$N��,���K��=���=[�2>��ٽ�a�=��7=[�8��F����=|�>�d>Qq>�(O>b;>��)>���9�!��q��<���H�C�����:�Z���XWv�Az��3������0@��\5ý`z���Q�D2&��A`�f��=�PT?Q�E?<`?�:�>���%�,>P  ��:o�F�wm�=�
�>J>?�J?�!/?�=##����a��Ɔ��Z�������g�>I�2>P��>-�>;�>Xj<��E>��+>���>�3m>U�C=>�S7+=:N{>] �>r?7��>�4[>!Ql={����ש���v�Fn��-�= ��?��(�;�#�]��{T�VҲ�vƭ=�7�>��<Q����l̿H����V?�4��� 	�M��/e[>ӳN?Z2]?�%�=V���9x�>���=��)���
|>L����k��$ �$�'>2�?ߎ�>vd>:55�v������	�žf6�>[�?#G��g_>.=~�m/�Uq1���>��>0`���_+�K��a"���:���	&>K�>)�>��=0�ؾ0p�������j�>�ߨ��ď>E��=��>�����x=��ѽ���=�%�=q^�;7�>���>/�V�)�>`4�������zp>�C>��>�#??!1?�b�=�@��`O�Y��>��?^?�&>�c�뻮=��?aO�=	R_�ep���ዽ>tH��+�>K�����q���l���>��ͽ��=Oy�>ec��+Ž?�����~?&y��m∿T�CL���hD?/#?DF�=}rF<+�"�x����E����?�@�d�?�	�Q�V���?79�?w������=�c�>ث>�ξ�L�]�?o�Ž�����	�2#��I�?��?�0�̋��l�<>�`%?y�Ӿ�h�>Bx�|Z�������u�)�#=��>�8H?wV��M�O��>��v
?�?�^�ک����ȿ>|v����>1�?���?>�m��A���@�E��>��?agY?%oi>Bg۾�`Z����>��@?�R?��>�9��'�^�?�޶?ۯ�?�+�=�ڢ?�s�?3�>���=]d�{�ݿ6���>�ƕ�s�=�F1�b���W�4��ۼ�\��b�[�g%�>Џ>��
�t��>�Ľ���]�C�-<"yB� U��yD�$�>�ā>)��>SE�>>�?�\�>���>���=�>x݋������K?��?���%n�!^�<��=��^�0?,4?�I_�O�Ͼf��>��\?i��?�[?KY�>����9���뿿}����Ɩ<��K>P�>'c�>:J��MNK>��Ծ�D�PQ�>��> ���"ھV&������dj�>�F!?��>D��=�� ?��#?�j>I.�>*YE�K6��.�E���>֦�>C?~�~?�?�ǹ�0X3�Z���䡿=�[�,6N>�x?S?��>Q���/}����D��I�᧒����?Wqg?%u��?�1�?�??�A?�Bf>�Q�Iؾۣ����>�q*?�9���A�p�,�j���H�>�b+?���>`%���^>�t��d���c?�,H?X �>%�1��e��# �]=�i
;P�r��#�=S6���Mb>�=	؉�tm�=K �=���=HU���f����=�1�=�s�>}�:>Z�i�)�M=�<,?�G�݃�8�=%�r��xD�|�>iJL>�����^?�i=�l�{����9x���U�� �?A��?�k�?t��ɜh�#=?��??f�>�I��}޾��ྞLw��|x��v���>\��>�;l��	�뎤�ș��)F����Ž88)�� ?�X�>I��>R�?��>w��>\1���-���̾�`��\oq��>�e�!����P��Q���4�u�=�{�S���m�>����;�>��?i�e>�@�>���>�+�����>�zH>*�>���>�s>�+>�:>��]<�= �kS?�̽��2(���+<���A?�a?�b�>��Q�(5�� ��G[?Y��?w��?�rg>/?h�`�,�?
��>����u�	?�H7=�0��n<|�����������f���>�|Խ�8�t�K�.j��,?p?�(��ٵȾI㵽~���ZPp=XY�?S�(?��)���Q���o���W�R S�i��&|h�
���w�$�B�p������n��� ���(�2�+==z*?�-�?�W�~��V"��c&k�;'?���e>t�>��>���>R�H>C�	���1�v)^�eO'�b򃾘>�>1{?�>��(?KGM?fʉ?��w?��>R�>�þ��#?�G+����>%�>t؈?<?��6?N�I?��+?�b~>�>L��eoѾAd�>���>�4�>[�?~k=?ʹ��D@?�<j�=��Ľ����*�@>���>ȟ">���ǭZ��ݘ=ٱ��?7*
��g9�� ���g>P�5?�_�>KO�>�V��p����@K<���>�?�|�>!���o�����>4�~?�m�=S(>���=T%�/��Lj�=C��-��=^W��4
G����:�^�=�Kp=��μ-��v�绹��<l�9=���>M�?gӉ>�=�>����� ��y�y�=	�Y>�7S>�>�ؾ
d�������g��z>�f�?���?�$e=�;�=��=i����+��������<�g?�#?kT?�]�?M�=?�>#?��>%������a���b���?|�9?���>z��8ž�1��������>�'�>�$�D����/�(���m�<�b>�iZ��ڂ����f���b=�9��t���%�?2L�?����T=�ۉ���𬿶�����h?�*�>�!�>�y�=;]0�m�]��{��t>���>�(�?��>�)P?��|?
�\?��X>l�6�D���Z��~���>+'@?lЀ?RK�?��w?��>��>
:'��߾=��n�����骅��e=��Y>7 �>���>��>��=��������	6��z�=�_>���>`�>g��>KFx>*4�<t�G?���>����$I� &��M���,�,�t?���?��*?#�=T���E��.��2C�>M��?�?�?vJ*?��V���=�x뼎����p�ڷ>w��>X�>���=C�H=ip>@�>+6�>0a�9����8�=�G�y�? G?�X�=G�ſ�q���p�
֗�/Ub<� ����d�"���J+[�㸤=�ǘ����ҩ�Z�[����k������-���f�{����>�z�=ˎ�=�"�=+��<�ɼ���<�J=$��<d�=�9p��|l<��8�&�̻����W����[<��I=;��҉˾ƌ}?�:I?V�+?W�C?��y>@@>�3�e��>�����A?�V>K�P�ˆ��e�;�%������۱ؾGt׾�c�G˟��H>EcI���>�93>7E�=�7�<��=3.s=PĎ=0�Q�G="�=�H�=r_�=���=��>�N>�6w?W�������4Q��Z罣�:?�8�>g{�=��ƾq@?�>>�2������yb��-?���?�T�??�??ti��d�>M���㎽�q�=K����=2>k��=x�2�U��>��J>���K��D����4�?��@��??�ዿϢϿ?a/>P��>��=\&Y���M	�����PL>j�?�X)��3���q�=��+?~�����"�
�(=��>t�=s��=3�r��!>��MՒ�Ot�=!��>ZM>)$C�+ք=K3>1�=y3��$V>�%>��	��y���I-=:�>"��>9��><t�>�Q?6^?aC�?r��>H.K�Uu���A��,�>�c>�&?kO>��?���>�I?��i?O[H?)��>N��>b��>e��>����;����<�`�[��&����?�y?�@�>&/�$mv��I�R'<��̽��>��W?���>(7�>�8!������(��>C�3SL��Bs�Q����21���b=<���'˽K0:�'�D>ԯ�>�>��>]�>��>k��>+� ?�D�=q�<}��=���=k��;o�o��u>��3�l����'>�3��ɗA�D=>�:�n���bM<+�>���=��>��>�1�>���=b�;��c>A�ھ�1G�N�j>(�/��:W��CP�Of������5��=;�>�cw=[Ǡ���?��@>-#;47�?�҃?O<>��=� ��B���J쥼�	��\�_>C)�>h�L�d#�17,��^?���̾�l�>�S�>.V�>,̾>������>��P���8�.?�o� iܽ�����n��7���ɏ���u���
��a?'������=��x?��?_��?9W#?Ҿ<=T� ��Jнbx=3��>�1��Ma�W���mD?Յ;?/?�Z�6��/̾?&��*_�>C�H���O�������0���,�Ε��.S�>7����о��2�{_���󏿏�B� �q����>i�O?�خ?w�b�ˊ����N�1��S,����?�g?�a�>�?�W?y�����^��)ҹ=po?~��?�/�?�h>+�=�=:����>X}?�?g�?�o?,��"��>����60�>_J!�q�$>:�u>�h>�`>a�?�?�?9��
�e� �����3�]��4�<E��=_�>��x>R>��]>�m�����?>姓>��>E8u>��>�u�>Z社���w�'?�~ļ��>��g?	�>
(����]����=u��>֜��u|�Z�=$1�=�e=r�:iI���:E>	��>�4㿓F�?v�q>��
����>��#q�>+�W> d}>	�ﾼ�P?��>�%�=HE�>';�>���=[�r>/��=;���P[>A���#��
>�PNL���Ѿq��>}��J�9�N�
��8����3�Qӧ�����f�ɓ���9�� <X��?sh�3�k���#����;?ꖜ>��1?�?m�xɷ���>#L�>^T�>����M��'��@��s_�?},�?�;c>��>a�W?%�?w�1�3�-vZ�,�u�C(A�e�&�`�o፿������
������_?�x?yA?aT�<:z>7��?1�%�ӏ� *�>�/��&;�8B<=�+�>/*����`�@�Ӿ0�þ�7�-IF>��o?6%�?vY?�SV���\�_�*>�>D?�2?d�?�M?��.?���=?6�.>�L�>�~�>�Q?+B?�`?D��>�B>��;��=�{���du��k�v.g�����i!6=:�U>�{ߺ�k��ڻ�N>����k�;:�\��"�=-L��a�f=���= ��>'kX?�1�>�Ց>z�=?����	?��嚾U�8?��M=�a��n��G����־��
>H_r?_q�?�]?�x�>�3D���D���=�1>��6>���>��>n��A���=Rt=s��=�*�=}x�<�~q�k�������ͺ���=~�>|�~>����%>눤�����d>�BR�C廾�,U�CPF���1���{����>BL?|a?-�=�E쾚ǩ���f���(?�n=?6K?�m�?Ƈ=��پU�9���H�$#��.�>��<t���R���٠�'T7�bQ��A�>�ѡ�	�H��œ>P�$�r���mQ^�E,|����hr�=�����9=��+�,��C����=���> ���&����ʘ���L?O�r=S�̾���!�r��8�>Ɛ>d�,>з���'�6V�R�ƾF	&>��?ג��ƽѽ$�*���B���9��˅>��D?��^?���?�〾�p�\�?��m��b❾�k��~?]�>�`?*[>�&�=iT�����d�$/D����>R��>D���<J����,�쾙#�e�>��?ɮ>տ?V�M?F2
?�a?��)?�4?�"�>l����t����?sI�?�uC=��B��PN���@�z6����>f�?��'�b�T>y�?R�>f�?�fA?l+?V�~=�z��D@��d�>�0l>�AN��e���Z>��=?d�>�u{?-�p?��>��2�����=�<=��=�[!?�?p�%?{�>���>
���y�9�>�
[?Wi�?��?� >�8?맬=�d-?���Z�>ҫ�>�!?"lr?�_`?��W?1�%?��=�Ž�ͫ�s�=󜽶e���V"��),��"���>���">�pf��o�<��a=��+=���=I�D��A��I�S>���>�u>"h����5>x�ž"凾@�D>���w|���+���6�㍟=��>�?�6�>�,�[>�=où>Zl�>� �8 '?�0?��?�`�Ta��Qپ��L�'��>CG>?6��=�i�c���u���B=i�n?�[\?mY�X�:�b?��]?@h��=�x�þs�b�j����O?��
?{�G���>w�~?��q?'��>�e�\:n����Cb���j�ն=r�>Y�-�d��@�>��7?\O�>M�b>��=�u۾��w��s���?��?1�?8��?�&*>c�n��4��N⾱��]�[?���>�1��s�3?�������S��5��O꾀]����z�Ο��x󅾇�#�v�q���ȥ�=�(? �?�Pm?�#Z?�8��:�^�2�e�������Q�U����.�G�2�C�̼H�}Ut�<	�QG��b��h!e=�z��<�pV�?w�&?���2�>0j������Ⱦ*>|X��V�4��=/b���".=��1=̓m���?��5��� ?��>vu�>#�:?��Y�]<=��E0�#[;������3>e�>�>��>i<%�3�S��6�Ⱦ��́ս��u>c?�RM?��o?~꽚).�����$�`�� ���I>w�>"��>��S��f��%�J";���q��"��ŏ��
�}�/=�5?��>#�>�3�?I?�f��ѭ��Bk�`�0��B<��>�{g?0��>��>$��{��Q��>�l?���>��>�\���C!�6�{���ʽ2�>*��>W��>5�o>�,��\�\i��{~��9�6{�=Ŧh?䀄���`�_�>iR? ܂:#�H<���>��w�+�!����t�'�u >�?6�=xu;>&{ž� ���{�#2����%?���>~'q��a �p9t>]�0?�>�{�>Hl�?��>����x��e�?��Z?��S?��5?N�>���<�u�����Ld���[=N1�>�Г>L!�=�AQ=i��E�W�U���`<�յ=�����9�,����#�����WDټ
?=>�Ͽ��=�{.��p��ج���)�֦B���^=#W���9�Jԭ��>+�蒺�0叾�M>��Ǿ��6�/���#�y;�?q��?7��׶�jN���ԧ��K��wMT>ael�M 3�r�ھ�����¾����������b(L�GJ��:�'?y���B�ǿ����7ܾ� ?KA ?�y?�ѝ"���8�� >><�<�Ꜽ&��ڙ��8�οb�����^?���>�	�r4��� �>h��>7�X>uJq>h��s垾�B�<��?�-?���>t�r���ɿ�����<@��?��@6oA?(�(�=��#�U=���>v	?��?>�u1�K)�����J*�>�%�?y׊?�M=��W�r�	��Pe?��<��F�\�߻���=.�=s=����hJ>�>\��$A���ܽ��4>�܅>mv#�E�� �^����<�N]>~ֽLF��5Մ?,{\��f���/��T��	U>��T?�*�>Y:�=��,?X7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?_D6?���>�d&��t�م�=|6�
���z���&V�|��=Z��>c�>,������O��I��Y��=��cOڿA�,������==No��2����=�}��k>������6�ܚ��B���E>"��>(+�>��>*_�>�?O?MX?�[>.�Q>�G.�1q�����"h�<�������,���"��!���ݾ��c�7�%��w�X�	�1��?D5���=��V��'����(��U~���C���)?��Q>H��M��jG8���
�¾�/l=����붾P�&��zn��?B�D?�w�T�X�o\���˽,��z�A?8�ʽ^! �>ɾ�>�<�Ἧ'�=^Ћ>���=�H �'C4��9f��?-��>�(d�Cl��Y��pZf��x���|I?B��>�\�=W}�>�7?菜��)�; <J�>���>�!=?h<>�,���׽�i?�j>?��bLd��y>���:N�6_=�I>�1R�_��T>(��=�����U>����&�=�hI?4�>m�,h�(����,󽢳4�) e?��?B�>9Z?*�:?xo�<�����y���>-�2?5�^?8^">*�.�����ھU@.?��d?gb>T���h�RMK�i�����>B7o?��@?�켗���r�����6�?V�v?�n^�)o�������V��5�>#Z�>e��>��9�Dq�>�>?��"��F�����|V4�e��?x�@Ԍ�?GV<<1&����=�:?.^�>��O��DƾS����{���q=�*�>ˊ��Tev�����_,�R�8?���?8��>���������>z�e�?��w?�ػ%�H>d?�Q�Z�cÚ�2���\Rq�b.I��>��侑}�ՍǾ���?���0�<��5>t�@ȗB>�X�>~y�� �޿a�ʿ&b��E�����u!?�dd>�<L��aB��}�}�t��:T�R�V�G����>�">�����ږ��m��e5��s�q��>$���g>��b�Ad��R��mܣ=�~�>T��>��P>d���r�����?z���'пk؝������\?���?_�p?���>�ާ��>��ƾ��:�6�a?�19?c05?�l�?�����j?�V��jT`�σ4��KE��U>h#3?53�>��-�2|=~>�x�>�h>�/��Ŀ�׶�,������?��?k����>���?�r+?+n��5���V����*�y+�V2A?{2>4y����!��+=��蒾�
?�v0?���|"���_?��a���p���-��8ǽ>y�0��R\�A���Z���He�j����'y�"�?�_�?��?ʅ�#�n4%?F�>�����GǾ���<-��>�8�>c9N>��_���u>����:�*	>��?��?�[?��������->N�}?%�>��?Ȗ�=�_�>�u�=�밾�5.�ER#>y�=!g?�!�?ǢM?�K�>�e�=�9��/��[F�RJR�Z"���C���>��a?�L?;=b>&���2��!���ͽ[1�;�輆>@�q�,�r�߽K5>O�=>�>�D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Sa~����7�c��=��7?�0�#�z>���>��=�nv�ݻ��V�s����>�B�?�{�?��>�l?��o�M�B���1=5M�>ʜk?�s??Qo���t�B>��?"������L��f?
�
@~u@^�^?)�yο*���a�ɾ����'�=�>n�>���IZ��J�>k5:���.D>7Q�>�S.>��>{[>v#�>�?�>�7���+�v���g���=��)�hϾ�堽�2�xf(>���w$���mx�R�6��@��=�uѽ󦝽QY��E�=�U?��Q?��n?� ?J�l��,#>����8E=��(�G�=v�|>�]4?�bP?�-(?R�s=晾�zd�N���l��2������>��:>S��>k�> w�>�w�;j�M>��8>CI�>��=Nv$=�ː;�=*�R>��>��>O��>��o>��	>f����3��z�H�A־��n�1��?�Q����4ר�a��y��h��>S;;�e��!�ÿ�|��LL?�J�����,���>��m?�=?Je�=�1E�԰�<A�>��v=i|��Ov�<���*�Y:��A�]Kz>aN>r��>��>�d&��r�?�:� �R�CnY>���>@�;�=7㈿	�`�����>��^=|�{���`���}�������.��B�=Z?�?Z\��܍����C<<���O�W>6j�=G3
>��b=��>h�������3�!��>z�2�� �>�_�>��*>�d>QD�>ה;y�¾�l&>�>:]x>a@?I�?�2�>��f�@!˾'��J܏>��B?O��>xqT>�H"��=O@�>�Xd>#�ܽ|�%��0R���(��7>֓�==��B���=>(#�o)�>��M=I���0۾�L-��~?r��%刿���u��gD?�.?���=��E<�|"�����#}��5��?$�@*b�?1�	���V���?j-�?����[��=��> �>!?ξ/�L���?	ƽO�����	�n#�jI�?��?�60�z���Al�5M>TH%?��Ӿ�h�>�w�sZ�����;�u���#=���>�8H?�V����O�>�bv
?�?�]򾫩����ȿN|v�n��>��?���?�m��A���@����>*��?�gY?Gni>@h۾D`Z�C��>	�@?hR?M�>:���'��?�޶??��?�E>��?$��?��>ː?>$����b���\��L<�=�0���,�>�+�=3� ��Q�h�����a��==��q_>��<�x�>^
8=Aݒ��X�;ǅD�����_���F> ��>�>��?�0?PP�>ƀc>f�]�<�=�R٣�B�K?���?����(n��,�<���=�^�C?	34?�o[���Ͼb��>4�\?q?B�Z?�2�>����6���忿3r��]��<��K>O�>��>�:��Y;K>��Ծ�!D�L[�>ܗ>hZ��{3ھ�7��GȨ��D�>$`!?;w�>�[�=q� ?(�#?��j>n'�>faE�X9����E�/��>Z��>H?|�~?��?�ѹ��X3�4���桿��[� 5N>��x?�U?�ɕ>W������q�D�&I�.3��?�qg?h��? 0�?m�??�A?4!f>ё�rؾ������>��"?���|A�>10�8���?uy?���>���[�������Z:����a?�8I?Wp?� ��Z�6��)*�<��:��һ.�=-48��>>�})>x�� �=O�>i�=�m� ]��(�<#ܩ=B��>mt>�`&�G�z�,?��A�L?��d�=Q�r��D��@~>�|M>�V��k�^?5j<�*0{��䬿q��hS�k�?ՙ�?WD�?˳�;>h�h�<?�χ?�?��>K��z�޾-���v��Oz��O�`>.�> �`�h>侖x��ew���U���Ľ���	�>�<�>\�?� ?��O>�{�>'�����&�ڠ�-+��_����EQ7���.�"�����#�#�=�	�3¾� {��Θ>AЌ�΁�>́
?S�g>�{z>$�>N.��&�>q�Q>��~>RR�>��V>��5>��>"�<��νq�S?����q(��޾%l���v??o]c?r�>+�h�����:��?B��?��?@vj>��k���+�]N?�>XKy�'?I�W=�<u��y���������)��5b�>Xp��`S3�~?K��	v�!?�o?|լ��ξLh���&����o=�1�?�)?��)�Y�Q��o��W���R�e�%h�J���`�$�up�"��\��@&��Z�(��)=�p*?�?�\�pI�ii��ik��>��e>���>�>��>�J>�
�E�1�K-^�A'��у��>wh{?T��>c
8?
�=?A��?�8_?�k�>v�>�4���?�2�V�>���>��L?�?�?�?�&?	'>�8�<�߾�"㾹��>��?i��>� �>�F?�Nɽ�H�<�<��':e:���6�FD�=���=ɣ��3�	��y��
�>��?6u���9�?���^h>K�5?)��>]�>/������,�<H��>F	?Uz�>�� �Rvs����$��>��}?j���=( )>{��=R��H�:3��=���)ߠ=�#j���:���<�=Վ�=��\����Ê<���9$��<ZV�>��?�Չ>E͇>����� �W��X��=N�V>?T>��>
�׾|1�������g��	|>��?�g�?�ug=���=�=���˧���`�Uf���q�<�?,�"?T?WZ�?=?�	#?�>3�-���τ�����E�?_I?��>X���4��I<��)���? �	>�0�����:�
�(��Î��ѐ>Zj�'��kA���6��3ǽI` ���/�-��?)\�?f���V)�\���X��Y���3��>�G�>��>@�M>����\�z�e��1�">�v>�c?��>�pd?��?��\?Lv�>�ϾϽ��T���\=�#��85?�Mr?���?G�Z?��v>rx5�&���N��þBg��l����k�>�*�=��;>�??9Â>N�>Hf��PdK=�׽j2+>�~o=y�>�,�>�t?�|�>�`M=�:?ui�>X᷾���=����虾6wh�r'�?��r?�7?9О=�u�b�B�a��ԉ�>�G�?��?�>?ڕQ��~�=�?��K%���}��"�>�@�>-��>�>�g�=.^<F&�>!��>�.
��_�9O�뗙���)?�3[?0>�Iƿ�r��
r�Ͷ���.|<*��cMd�����:<Z�0�=�����c��ũ�=[��������8�������x��+�>BD�=-]�=$��=���<�kӼĺ<�vU=T��<�Y=�Yv�^�<�r?�D໅���x2s�F[c<5�J=��ݻ˾?�}?=I?��+?F�C?(�y>N2>B�3����>�����@?�V>h�P�����B�;�����z ���ؾ�v׾��c��ɟ��H>TWI�k�>�83>�E�=�2�<$�=�$s=�Î=��P��,=D#�=�Q�=tf�=t��=u�>�R>�4w?!�������2Q�;O罝�:?7K�>#��=�sƾ@?��>>�2�������_��.?���?�S�?r�?hi�f�>Y������q�=pȜ�VC2>���=��2���>G�J>�|��H������3�?]�@r�??Dዿ.�Ͽ�q/>�ڌ>�k>Ŭ:�twy������ؘ�gH����>8�j��q]� H��&��>BI0���֡�N�>X�����n���f�<�y<N>�N�=mh�>f>;H���O<��> ��<��y>�>#��=��:5b글`B>J8�=�a�>�g>�K�>��?B�]?Ǿz?�u
?�����p�'������>��Lz?�>#=���>�O�=��B?��+?+tD?��>&�>1��>��>5c)���}�^J��j�� ���ք?��?�$�>�(��N=�L�,?K��A���>	�A?3�W?+Q�>E����|�:����)���9y<{(�<t}�=W��\��>�׽���0O�=���=\��>��>i�w>�G�>d�>���>d��>�\4�L�C��-=xŹ��֎�mS�>ǵ%>��=�
~��v>MB�� �;n�i>g��T�x���+�=2��=���>�H>���>j�=����/>������L���=
3��B��"d�^>~���.��r6�5�B>hX>�@���*��M�?�Y>?>΀�?@u? �>0-�-�վ!T��(Le���S�z5�=Q!	>�<�؉;��f`���M�U~Ҿ��>$��>���>Z��>��:���+�fA>9��,n�#�>� �l=I����;C��h﬿Ы��xKI�~h��+?+����"�=yq?$�>���?r��>�����/�˃>B;��h�>
#3��TY>��,>WWF? ��>��:?�[���	��B̾����ѷ>EII�\�O�����0���A̷�.��>����M�оI$3�6h������D�B��Lr���>��O?+�?�2b��U��COO�����!�� j?�|g?��>�J?6??�I���o�D}��,h�=��n?��?>�?&>���=CT=���>i�?Ó? W�?��x?9ȗ���
?���?1����M�>Zc�>���=ڼ�x?���>Dc?���.���W亾����|���>��\>ﴬ>W9D>k�>1��=��ڽ�/�=��V>!r�>=��>>�=�\�>�h>%������� ?���=��p>ZAA?P&�>=��=d��=��۽�~�=؟�^7�=V K>2+=�x���1�=9q8<�b�:�`�>�ÿ���?��n>���0?��F�Y>)��>&�>��~U&?�Ί>�}��Q?*��>Os=n�Q>&�>9/Ӿ��>��<d!��(C���R�)�Ѿ��z>W���V &�����h��PI��n���a�"�i��-���;=��K�<�C�?\�����k�_�)�������?�Q�>6?����f���^�>���>�ˍ>\����������\���?��?�;c>��>3�W?�?ے1��3��uZ�Ůu�(A��e�
�`�L፿����$�
�����_?�x?yA?V�<:z>4��?��%��ӏ��)�>�/�I';��B<=}+�>�)����`�S�Ӿ8�þk8��HF>T�o?%�?SY?�SV�s�e���&>�;?�=4?t?��1?��=?dh�,V$?J�*>�~?F9
?9(6?M.?k�
?�6>�q�=L=�wRD=�����n�����]�ӽ%f	�� >=��=QA<�\�;|)=�A�<p\�&z���?;�c[��<-=+7�=-^�=c��>x�N?�8?s?|>�LC?��S���@�5<���?I?���=�S����{�0&��s��e��=H?d�?=uk?T��>��:�fh1� �<3��=�Z�>�ҳ>�,�>����\0�8����	>��=� ]>!8�= ���N��d���{ҽk?�=���>�se>��?��/>/���q6��LW>=8�Ay��Y P��G�;�/��)B�4޻>��N?�z?Mx�=���rJ����_�350?�69?�:K?���?x��=���lm?��G�Dg=��؎>�r��q�����������!4���[�n;>j���-�Y�Tk�>Z�#��T��yk���^f���8��>9x羍����v�3��2ذ���=tً>0F����o�斿b=G?���=�g�,/ԾKj���|@> h�>�&�>r���m6,;�m8�������?onD>H|�<��4�ۚs��o4�gF�>ggE?�_?4{�?Fl��mtr��C�����ġ��Hȼ��?h	�>��?�B>��=	c�����.�d�M�F����>n��>�8�G��垾 ��)4$�`�>��?<>e�?��R?�E?�B`?��)?K�?�ב>�f������&?�K�?���=��Խ�
W��{9��C��*�>�H)?VDH�{��>f�?��?K�&?�R?}�?�
>�� �&V@�I2�>�>�W��^��c>tK?�ֱ>�X?B�?��=>��3��;��4#�=�>�x2?��"?��?��>���>ϊ���M�=�X�>e)r?i�?oTg?��>��?�W>���>��^=3��>��>1t?BP?��p?�7I?M�>;(<�ם�V���6l�}4���J	���[=��[={4�P�(�I�"���~�<Q�l�*$	���9�՜M�3��<�RE����>��`>S��$AL>�DG��>�r>^��<�4��T��vQ�M�X>�S>���>(y�>��|�q�>��>�l�>����)?���>�?ͽ�lc�y�ʾxuc��]�>�;?
i�=��p��Ꮏr�m�9~�=�`?��U?;���
o�\�b?@�]?�M�
=�B�þ�b�P�~�O?r�
?��G�Vܳ>��~?T�q?��>ȝe�u-n�[��� b��j�'0�=%Q�>ja���d�qW�>�7?!)�>ͷb>�y�=�T۾��w�ZL���?��?�?Y�?��)>��n��5��*پDȍ�!q_?�5�>F�o�9N(?�BW�7 ���tM���u���⾛����#L��+�����S���ow���ٽ�>��?L�?*#�?&bc?�rؾ�a��z�F����nJ�B�"�xW�D�S��>���L�pS����)�E�� ���|�"=:�~�}A�Nh�?X�'?z�/���>�d��E��̾g C>�Z����;�=�����C=\GZ=;]h��).��Э�� ?�7�>�Z�>��<?T�[�I,>��|1�Ĳ7�����T*3>Ro�>�Z�>�>+��:@�-����	�ɾU���2Bӽ��v>I�c?\eN?_q?p���+�2���k(�]������FJ>��	>��>��P�5m��K)���<���p�m�
�������
��� =�6?�>@��>4�?��?&��촾�l�w�*���=U��>`�f?��>2U�>���~��	��>��l?}��>��>
m���?!���{��˽��>MЭ>���>�uo>w|,�i\�f��ۉ���9��h�=B�h?
w����`�D�>xR?<Zk:�E<kp�>� w���!�:��ӛ'��>�?h�=��;>��ž��{�u*���(?&S	?z4���6)��c�>��"?�n�>�l�>d��?�B�>��¾�׷;B?tC]?��K?�xA?��>|{=câ�v�½"��J=I%�>��V>�==��=D��OW��� �i.=X��=O&Ƽ�m�����9���C5q<�]�<#2>��ɿ'�I�b�����n�R�	��0���=�0h�l5��x)J�Y���k�Q�=�8ľw����E�)]�;��?H�?�#��/ҭ�<ŧ�aՍ��0˾t-I>%��<s���򲾲�>����:T���$���&��(�j%�(gW�ԕ'?���H�ǿװ���:ܾ6  ?fA ?�y?��˝"�Ó8�Ȯ >��<�*��'��ҙ����ο����^?\��>��������>���>[�X>VGq>w���螾DT�<��?Z�-?��>��r��ɿ5���S��<~��?��@OXA?-}(��C�ͬT=�|�>�	?�>>�/�����}��Y��>�\�?��?��E=o�W�7&��|e?�<'�F�&�ܻ.��=�)�=�=lI���I>:��>��@��mؽ!4>��>ރ�@��s_����<H[^>s�ѽm���5Մ?+{\��f���/��T��U>��T?�*�>W:�=��,?X7H�a}Ͽ�\��*a?�0�?���?$�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=l6�y���{���&V�z��=[��>g�>��,������O��I��U��=Y��S}ʿM�;��O!�d6�<��-=���=Q�/>G�*���X�����L��ڽ�{=�df>~s�=��><>�n>�l?wl?g�>{�>b����㚾-什.�Z�_d�
u����<�#þR��/ξolE�\{ݾ�{�W}��r1���=,�\�M�����8���m���!�t�-?�X5>�ξ��J�
��=�Ѿ䙴����<RG<��Ԙ���%��a�3)�?�E?�)x�|�Q�pi�4J����o�pWD?�	�!b�8��2L<�lo��g�=Ԁ�>^�=���H�F�n{T�a1%?�t?����y�q��I>�Ғ���V�r�.?���>��;\�>��H?���#����T*>n�x>���>L?)L,<Œ��.h��<?�-?C����=�J��CW�M �>)�=�j���nI>W��>�ҽ�7���_�Q�S>8�N=dR?gȜ>"B�\���ϛ�����B�=G�h?Tv	?�i>�b?�a%?�چ��A��0%�����ж��oKK?��e?�M5>³��������þ�B?'h?;�a>�9�����&�����>8$[?��1??�U��Jy�Uܠ��,��0!?Z�v?LS^�!O�����XGV�M�>8��>��>�9�ҧ�>]>?*9"��0��Ի����4��Ğ?[�@]��?dc5<����=s.?,[�>>�O���žb	����s=
�>Fw��:ov����Y,��k8?r��?�a�>m����t���>|��Su�?���?�G���X>0<@���c�[���]�$��u�=<f7����=��ѳS��g�t�����?��=�&I>~�@>�ګ>�'E�������俠S��:�����$K#?9z =؏�����{Ԑ�Y���T��D���#��j�>a�!>�'���0���~z��#A�?2�<���>���(X>�u7�������z�=3��>��>A
H>[����x����?�O��ÿY����}�R^?m��?'z?"T�>���<�傾]����vA��@G?�*b?�
E?l	�cm�k<����j?GY��3Q`�j�4�xGE��U>i"3?3>�>��-���|=>���>'b>�/��Ŀ�׶�$�����?��?p꾈��>݂�?�w+?Xj��6���Q��m�*�@�4��=A?�!2>�����!�>/=�Ғ�a�
?�}0?i���(���_?��`�p��)-���ɽ�W�>.�.�:[�M��jQ!��[d�aΛ�TM{�'�?j,�?l��?���Ds"��R%?�\�>���ƾ�Y�<�:�>sI�>�N>��Z��en>���f�:��Y>��?jj�?)B?�y��k��.>�(}?@\�>8%�?��
>[��>+�=d����<�Y>��{=�Kv����>Y"I?`��>��=k���u*��K�:/Q��e ��sE��9�>��m?^[?�B>�|νHP<�w"�ZJ���˽��H=ՀP�I0=�����H>m;>�1>�\W�v�����?9p�1�ؿ�i��q'�E54?���>�?���մt����-<_?
z�>�6��+���%���A�Q��?G�?Y�?,�׾"W̼>@�>RI�>��Խ����񁇾��7>�B?&��D��K�o�H�>���?��@�ծ?Gi��	?���P��a~�Ԃ�P7���=	�7?J0��z>���>)�=�nv�ۻ��?�s��>�B�?�{�?A��>Ϯl?q�o���B�?�1=OM�>Q�k?_s?�]o���2�B>c�?��������K�Qf?��
@ku@��^?��+ſǬ���Ǿ�����ΰ$�iN>������պ�>;l�=G��jx�=��+>)��=�wM>���=��>��Q>�����c��<���䕿 oY�E�,����t�y;��*a=���~���$ľG̈́�JKL�%45�2���G�L������=S-X? �O?��k?���>��O�np>����=�$���>}�?>5�4?<�N?
@$?�4=���_��n|�&A��A���F�>@��=��>2��>���>�=w�s>}�=���>4Ѻ=�P�=�ޖ;��V=E�I>�E�>�-?I@�>�'�>�<>�ͯ��w��rz�γȾ�>>��?
8"��
�R ��6X�������q>F�?�6����xCѿ�^���]H?H�ھ�f��wk��e�>{l0?[^�>��M=���Z�=�z�<�\�������<������=s�8��M>|�W>U(�>A�s>��>�ӠA��.;�,֠��
�>�'�>Qn���=�L���ݾM�&��G�>�ʐ;,s��]�<��o�{�K�D�S>�B?U�>̴%�ü��xQp���q��v�>�� ��'>}��<�?>y`.�S�K=�H/�ZN!>�Ѵ=@Xv>( ?� P>�D;=���>�������~�f>l�
>�4�>DB?��!?!�=�0���LǾ=�g��>A2?�;�>��!>fZ�=q�=��>!�`>M��+~������� J>�5�
4��CϽԵ�=�ﻼl�>>󼏼���+�(�>�~?���䈿��	e���lD?R+?u �=��F<��"�6 ���H���?n�@m�?��	���V�7�?�@�?�
����=�|�>�֫>�ξx�L�ñ?��Ž;Ǣ���	��)#�`S�?��?��/�]ʋ� l��6>�^%?U�Ӿ�g�>lx�{Z��Z����u��#=Ω�>�8H?WV����O��>�_w
?�?k^򾜩����ȿ�{v���>
�?���?��m�|A��X@���>ܢ�?kgY?;ni>9g۾�_Z�O��>��@?pR?��>�9���'�u�?�޶?���?^�N>���?�5�?���>�}>��b���п�Z���wA=�a� ��>t*��+��Ǖ�m���ݟ��t�o����>S�(=��>����-+�����:��o���7$����>��>�D�>��>f?6�?�?����k��rݽ�7���0I? ��?N����c��XM��	�<��,���>��4?�.���bо�0�>l8L?]~?8^?q'�>���!���^��������<G�<>O��>��>�Y�ȶQ>�Ͼ��B�,�y>SH�>��*�O'ྭˑ��*�;&��>'�#?��>.@�=� ?�#?}�j>f0�>�YE�7��z�E���>��>%=?��~?��?�Ϲ��I3�����[⡿I�[��9N>��x?�T?���>A���V~��k�E�!�H��������?Q`g?Zv�L�?h,�?D�??��A?"f>�v�ؾ����O�>��.?��t�,�&��� �?(�!��>�	?�>ܪ��&������&��}5?PB?�m�>�(7�	a<�dHþ6@�=E1B��T����m�=dc�>kq�=M��!�;o�=붽�����d�apҽ��	�>χ>�Ƅ�Cɍ�r ,?��5�̃�2��=�jr���D�}}>J�K>Zվ�B^?<�;��n{������i��K�S�R�?\t�?�Z�?����Sh���<?�?5~?�h�>Az��5hݾ^�߾F�x�NRz�FB�CE>��><�� �zs���િp���ýS{��?�}�>wt?�b�>YY>���>���&�@�߾���|a_�Hu
��;-�,��s�=	��V�1����~�Ӿ�Tr�ԝ>�ȥ��V�>�x?�i>a�>�b�>:��!q�>��!>'�>�i�>ۍd>�f#>V�.>J�r=�a�{PR?!y���'�)L辊˰��A?Q/d?���>N�n�9��M���?JP�?X��?Sx>�h��K,��X?���>>T|�Jw	?%p(=�0V���<[S��'��l��^@�詎>���k9��K�ddf�I�?IB?�����̾7�潺���҆o=�P�?g�(?�)�Z�Q�?�o���W�S�[9��*h�}����$���p� �G_�� $���(�5�*=5�*? �?������d��k��"?��f>���>�$�>r�>)KI>B�	��1�^��L'�1Ƀ�3A�>0Y{?.ډ>c�A?[O?�}?��i?t��>��>�ھ2��>�ֽ��?�W�>�a?,*?�E&?��?)�$?��>�z>����:�;_�?l`�>b?UY?��?���J�O��$�ğ|=����i�oʄ>�%�=�
};l],<a>�az=e�?l;��5�|� �-c>I�4?�I�>W[�>ꖔ�Z���M�껖\�>U�?�t�>�k �9dm�b�����>�by?���֍0=��0>�q�=����!X;��=��ZJ=����8J��B'=n��=)�.=wr��ߥ;��<]����<���>*�?c!�>��>��o���v��J=&=�>U<�>�1?>S}��B���87����e��q�>h~�?���?In�<�=:� >üоᒉ��;#��K��'�>&��>҈?�h.?&x�?�-?���>��}>����5��l�y�vm���)?
5?�!�>�5��,�;����?_/�>�ic�fO���%������_��1>0NI�t�m��"��%OA�Vvt�<���ͻ��?���?p���+��d��b���4���;�C?\y�>F��>�k
?S|%��hb�9�	�P#W>5��>t\Z?6�>1MU?Y+�?�c�?���>�eվ�+��$5���� >���=�5P?��Y?㷢?j\_?�a�>ؽ �(�����D�-���V�n�aC��+��>�q>!��=�m,?N�>h!\>�@~�0́=�|I=�P�>u� >O��>
_1?��?q�> 2�=�B?>�>�����-	�����P����q?Xs�?�+?�M=���?��
�K�>��?��?��1?Ly����=Te:�����-�f���>�֮>"�t>x��=�S�=M%>s�>���>�rٽ{A�L�9�?���1Q?��G? ��=d���V�n� ��������Im��3��z%�'�"�b�IM�=e���zI ������q�	+���X����݁��jo�d� ?�r�=�g�=�#>峑�(ꖽ:��<�Ü<�{o=���<@����&�<��X��1:{����\��'�G=SW�<H<��˾	�}?�<I?h�+?F�C?t�y>�E>2�3����>p���E?�V>�hP�⁼�J�;��������سؾ�w׾8�c��˟�A>T�I���>�@3>f6�=��<�'�=��r=��=�qQ�=� �=�U�=f�=��=
�>W>�w?􃁿����LQ�I��o�:?���>��=,�ž�2@?J)?>}�����hp���~?���?jW�?��?�`i��X�>bĢ�������=2T����1>���=�2�q��>�J>`D��+���t���%�?P�@�q??�׋�ҪϿ3Y0>��t>��N>�F��L*��%�����b���=�?�����{`>��>ê�B�ǼI>0�>�=��o�[�h���=ཀྵ���>�싽�
�>	ݑ>���ņ!=8好�/
>���=�A�>B���K��H�6��>�a,>�[�>a�>�M�>G2?H�W?�a�?&U?�=�����%��>��P��?C��=<S?p�5>��K?�~?��4?���>_M ?��>/ L>[�>���L�i�];�$��cr�,�?�_r?���>�6_��J�U��>Q���l2!?
�?ٛ�>���>���>�翪|1�~�=�-��A^�;Ӂ�/�a�+̪���ֽ\�����	�=6(�>��>A��>,��>qZ�>W�>⾙>E�=eŽ�>E�=�2�=p�=pU�>Al�=����=���Q㙻H{�:sk�='s�=�*�=�J�=j���b��<���=���>g>r��>h�=����/>ϼ��]�L����=���-B�Id��4~�/��Y6���B>�X>l|��6���?#�Y>�R?>v��?�@u?7�>���վ�K���d�i�S���=��>��<�(w;��>`�O�M�M�Ҿ�R�>Ki�>2��>�e�>71'�@��� i>���S�@�m��>e���l��I���F�ў�`�����`��<���/?� ���t&>���?��N?l�?��>�χ=�O��.�>��Ὢ��>"�,���$>����6�0?^?�#?KI��&�<��H̾�L���J�>
�H��P�����_0���>���R7�>
��X�Ͼ�3�TX���᏿�B���q���>�O?C�?nua�P���O��,��ׇ�Lq?3g?(R�>6?(?󠽂f�hL�����=��n?��?��?�
>I�=���<
G?�?J�?Sx�?�a?z���{�>�pQ�&L�>�H?��z�>ވ>���=?^Z>��?�?+u?H߽p�zN޾�F������*>U�=���>��>�&6>���ț;���=E�>fze>��=bg>n�>My�=3My��F��*�%?��=1M�>
�[?2�>��>��e�g���@�>�M���=6b�:�R=!i<Ab�aUH=��M=���>��׿z�\? >X_����>-$�"�>_�c>씻>���3T?���=<=���>���>�6j<F>!��>'Ӿ�Y>���_!�Y,C�}�R��Ѿ�z>-����&����}����I�~^���T�wj��&���/=� ��<KB�?/.��U�k�	�)�ƙ��!�?+L�>��5?�ǌ�<|��zs>���>��>����������hY���?���?	<c>��>�W?ޚ?��1�h3��uZ���u��'A��e��`�7፿	���T�
�����_?�x?/yA?�M�<�9z>!��?��%��ҏ��)�>�/�';��@<=+�>f)��q�`���ӾP�þr7�|HF>G�o?%�?rY?SV��M5���=�:?N+?��s?��5?jU7?�rɽ�$?�T>� ?v�?��;?u*?�b?~K>�:�=u���=D}�C����ц�������i�,��#='���ϴ<�6�<bRѼ�%��讼�`�<�T�M�o<aoU=�¡=���=Ů>��?.�>Z&F>=\%?�\���K\�䂼��h?ʁ�>љ��^~>4��eQ�����:p�?�\�?y�?PG����f
��ަ=rFn>�X)=_�a>�0�>�a���I"=��=h��=��<�����OR����h���������:o>gt�>�{>eu��q $>�Ѣ���{��Ah>��J�>��3UY�QE�
;0�jFy���>ByL?�?7؈=��羁���c���'?s5;?�I?P?��=٥޾�J8�o1K����֜>�N�<���ݡ�-��q�9����G�x>�k��:=��e>X�ѾU���[���=�����(S>��iZ=�+�����'彾,�m>���=m����s5�`l���7����=?nBo=�ʾX%��!w�3�j<�Э>;�>Ț�` R��QH�0�Ծ��=>�>��z=Kj<��-2��Xd��1��@�>�WE?kM_?g��?�C��P�r�IlB��W��� ��¼� ?9;�>c�?�3D>�I�=���L�nd���F����>o�>^���G��̞��;�>Y$��+�>��?\ >w?��R?��
?��`?�*?I^?�>���(���3&?��?ј�=c|ҽ��S���8�!�E��[�>i)?�RB��^�>П?3�?J('?p�Q?��?\�>�D ���?�;��>�>��W�a@��-�_>(�J?q)�>��Y?�ȃ?J�=>�b5�"آ�ę���U�=�n>k�2?K�#?�|?�v�>S�
?�'���6��'����	?�q�?���?y��=�x?Qr���65?m����A;>=��>o�?V�o?G<{?�`?|y?��#=+�P�,Ԑ����<���������;�,->M=z�^�d�7��1�=x�@���Ӝּj�W=o�M��ǽ�Ԅ=!*�>%r>�+��Z�/>�\ľK�����?>�g���ě�������9�ݸ=�o�>�?{�>��"���=~һ>���>V����'?��?�>?K2;Gb���ھ�eJ��ݱ>�TA?���=��l�eH���v�>�a=+n?�E^?QZ�>0����b?z�]?Vf��=���þF�b�E���O?�
?��G���>R�~?��q?���>��e�@9n�����Cb���j�Զ=r�>X�v�d�?�>O�7?�N�>��b>��=Hw۾ �w�r��L?�?v�?���?
$*>�n�\4࿖��	����c?Xk�>T폾��#?}S������B�;"���վ�!����B�6������AAܽ7{�5d�>�%
?�	{?�k?Y-j?���e���\�݇|�K�0�����'��T�)�J���\�����������=���C$>Fq�$�E�_�?�?ޑ#�j��>0g���dҾ������->t�����c�>�f��p�=��v=�]b�T�^����?�m�>Ӻ�>�A?��P��z;�R�/�2�*�{v̾���=V�>D`>�	�>�}�s�V�;�r��/ľ������~��Ñ>n?�_O?9��?qϭ���/���S�_�ߒ�=i����͠>���=���>j� �Ćo�/fJ�KP���~����f放�"���W��[?k$�>c�1>��?�:?�v	� a����r>�P�037>_��>���?�:5?��i>@�>�$1�Z��>h.m?��>�>8\��'>!�0�|��!ս@}�>i­>J��>c�n>6�*�P�[�n}���ώ�� 9����=kh?*���
�`�ہ�>s�R?)j��(<%�>�Br��~!�|���&�>�>r�?�ժ=�RA>�?ž@�~|�Fˊ���(?���>(���-�^�6>�u$?�J�>���>�N�?�#�>|�^�����y[�>�	V?��C?t@=?��>z� >v��y����
� ��=�Έ>��G>���=��
>�-ǽ�AJ� M��6=�n�=���#ͽy�m=���{Y�;)� <ο>g8ܿS�M�����ھ6&&����R�潵�B>�gh��Bt�����d�3���@��?��G��=����F�<�{졾k'
�=�?ay�?�jx�m��H����G������Z>�J��Pr4������9#�E����Z���������9�Wb���j�[�'?�����ǿʰ��$;ܾ�  ?�A ?�y?����"��8�1� >r@�<k"��ܝ뾞����οJ���&�^?C��>�-�����>Ť�>��X>�Iq>f���螾�7�<\�?��-?��>��r�(�ɿ@������<���?�@�.@?ϙ)�Y���G=���>��	?r�9>('�b������^�>J��?�o�?�|N=��T�X���I}c?�1<��[E�˻��=iկ=6r8={4�{vE>���>,U���2��6�N�)>���>��(���%if���=*�Z>O��bс�Մ?Lz\�Kf�У/�zT��
[>�T?o)�>�?�=~�,?b5H�}Ͽ"�\��*a?20�?���?��(?�ؿ�Wښ>��ܾ҉M?�C6?���>�d&���t���=0�*�����5&V����=)��>�>ȃ,����z�O�7N��^��=���2�߿ !�Y-���28�%��#��=3Z�>8�P���>{Y��v~�Ŗ8�W���.�]><�R>p^>�Ҽ>�aZ>{�4?��@?�Tl=�#>��<�Zu��H����>�����������I3�N��������t����]��E[��q���0�u��=V�I�kr{�;�h��|p�{��}1?��<��Ҿ��F��=<��̾,�����=PP�1�þ%A�
�n�Eթ?�9?l0����g� C۾W30=1C�:L>?�8޾���¾�N�<vc�]"=@j>e��=���
>������?���>#��I�l�0�D>~Md��B�km?�W
?��V>�k+>��?�k��?����(->�@�=���>��?8��<�L��C��'�%?PN4?���ؿe��Lx>�B��X�9���=�>K����=�}]>o�=�C������J��oV=�W?�]�>B�)�*��ސ�R@���C=ʕx?;�?�̟>V�k?��B?J��<�����aS�s�
�nm~=�W?d7i?��>Ƴ���jϾ�-��U5?1We?oP>��e�32�S�.�j��vT?cn?�?�P���I}������v6?C�v?5p^��r��}����V�qA�>\\�>~��> �9�l�>ݑ>?�#�[F�������U4�k?�@`��?�;<��Պ�=�:?�^�>�O��<ƾFx������q=�$�>t����bv�{���[,���8?���?ב�>����8��h,�=��I�.�?O��?�q����A=r�0��KL�ły�c$���\ȽS�?��@>�:�=d����|C�}~��B>w�>Ѯ@���<d��>lg��kҿ-ۿ����8	���Ǿ���>�Ɠ�����¾=֧�@c��r5]� )
�|�޽�>�>z�>�^������9�{��a;����U�>,X�܈>��S��#��~���3<�>���>��>7ѯ��彾	��?�]���0οN���f���X?�L�?f�?�G?L�6<��v��t{���u-G?pps?�	Z?� &�w�]���:�%�j?�_��wU`���4�vHE��U>�"3?�B�>T�-�[�|=�>���>g>�#/�y�Ŀ�ٶ�A���Z��?��?�o���>r��?ts+?�i�8���[����*��+��<A?�2>���H�!�C0=�UҒ�¼
?V~0?{�e.�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�#�>�?�[�=`Z�>6e�=���ʈ-��n#>��=��>�Z�?R�M?Z@�>�b�=<�8��/��WF�YBR��$�t�C���>��a?��L?�Fb>0���+2�!��lͽ�_1�b鼿]@� �,���߽P#5>��=>u>��D�WӾ��?Lp�9�ؿj��p'��54?1��>�?����t����;_?Qz�>�6��+���%���B�`��?�G�?>�?��׾�R̼�>:�>�I�>D�Խ����]�����7>0�B?W��D��u�o�x�>���?
�@�ծ?ji��	?���P��ha~���+7����=��7?�0���z>��>��=�nv�̻��;�s�׹�>�B�?�{�?��> �l?��o�G�B��1=M�>��k?�s?�Lo��󾄲B>��?������L��f?�
@{u@Q�^?Yտ����F�����^�A=!��<ؙ�>�X��}����>��H�:�Q>k�d>��>��>'k>�>ըK>�]�>@<���\*��͓���s�Zb���9����D�H��B���Z>�3V�+���1"�:ݸ�b|/�(��<	kx��n7�!�=p��=m�U?��Q?q�q?D_?`����{ >�Z ��p=�B � �= �>�3?M?n*?r�=xE���Ec�����TЦ�'����>l�B>g��>���>-�>[��=�B>	�G>��|>|�>��?=fi"<�=J�R>��>���>6�>z�[>�>�ĵ�Ϣ����e��ѳ�C��� �?��/��4�Q`��%`��%����ȇ?׫�<�9����οWͿ�V?�t����J�nU���a�>�'?l?� [=AY��r9[=�Rۻew#�I���D��>�n�(L���'��&>W�>���>��w>	�;��5�i�(���V4>��7?�]�����o�j������">U�o>�wc<v#���������X�8�=�&L?���>��2�َ��0�N�о�6>��O>^L�;�˦�|Zp>󉼽�%J�3ъ�nC�����=[�>���>z_�=} �=E�>D	���z��G>	��>mO?C��>n]���n���ؽx�<:e>@�>��>U�B=a��}�=m�?�O�=�(��UY�<~�������=-`�����������>9XS���&=)�=�Q��	��=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?��>�<�?+u�?�]'>��:W��[�ٿ弸�"6�>8�������T�|��<�(�28ؿ����Lx}���uj�>�t�=�b�>��p� ��4�=Ϋt�F䫾��P� �">~.?�G>=� ?ë�>rY�>�� ?���<b;׼���N��u�K?K��?����2n��X�<Ɯ�=X�^��&?nH4?Hs[�%�Ͼ�֨>�\?$?Q[?Dd�>9��;>��q迿A~�����<M�K>b3�>�H�>�&��wFK>P�ԾY4D��o�>6З>x꣼�?ھQ-��KK���B�>�e!?ӓ�>aԮ=�� ?Ŝ#?��j>�'�>�`E��9����E���>"��>dH? �~?�?NԹ��Y3����桿:�[��9N><�x?�U?ʕ>"���T�����E�GI�/�!��?@sg?�Z�{?�1�?��??P�A?O+f>����ؾ䳭���>�"?����8D��$��m���?�*?���>PQ����ҽ���b��]����_?�QX?��$?���S`a���˾_�<��,��~����E<�����G>R>�6t��b�=�n>R�=�b�h5�YJ<���=��>	��=Ҍ4�Tʃ��6,?�H�ۃ��ۘ=d�r��tD��>XL>����v�^?ģ=�\�{����)o��U�%��?���?/m�?�C��:�h�=?a�?
?=�>�9��0d޾_��(w��xx��l��S>��>#k��������%����<��<�ŽTA����>���>(�?�C ?*iM>��>~����&����J��w�]����)8�.�.���us���}$�GF�Ȳ��z�{���>�d�>��	?�|e>�{>(��>+'���܋>�7R>���>���>(�V>��4>�G>�A<'�Ͻ�&R?���?j'�Z��|���<B?V+d?FZ�>#,h��u�����l?���?�f�?1�v>Eh��+��(?X�>���|3
?�};=P�2U�<�H��w��Jm����
���>ٽx :�3�L��.g�*&
?~?x���/6;��ֽ�/���u= _�?��(?��)���Q�hp��W��|R��<$���i�ua��s$���p�
@��ș���$��z�(� t1=az*?�U�?^�T���6����j�ӳ?���a>�>*�>g��>'`G>��	�IF1�ڟ^���'�+�����>	{?�1�>�&6?��H?�F�?1�?��?���>|�Z��4?��y�]��>d�?��"?X/?��N?�Z?��-?�v>:F>U�ԾH�Ӿ�$�>H_�>�?½2?��>.�Ծi����	�wC�<j^2���R>!�,���H�날��K�=�>�<��=א?%��w6���6~c>Ja3?��>X_�>+~���Pr�O=GK�>K�?Ε>�����n��n	����>��?Q���
�=6�*>��=�/2�i|i;XY�=�@���\�=�D9�Q4'< ��=�=�s[9$��:N���W7;�+�<�6�>�u?�(�>��>�X���� ������=�
[>��T>��>�پ���Vӗ�-�g��-x>rs�?v�?�?c=���=.��=(������u��Yӽ���<a?��"?N�S?�i�?��<?��#?R�>ڽ�j��ta��آ���?��,?/�>�����z߾�J����?��i�>zz>Vd������m6�%��7=�´'S�Q��O˿)Q�صҼ����R<p#�?��?������B��\����q��5?g�>�b�>�[3?!�W�Çh��� ��s�=}�
?S�?��>��S?��w?�}?;Q�>��,��t��B@����q�9V>hV?|�g?���? ��?Yc�>~��=�撾��Y���ܾ��ػ]�������'���<>�4�>kg�>���>ɕK=:#��f��ƿ=��5=��>A��>�0�>uM�>*��>�ۻ��F?E|�>��Ǿ=e������W������j?p�?�P&?��=����A�A?����>UF�?�4�?=�0?˿E�f->�@L�1 ��\]�l��>`-�>���>�=�a9=c (>y��>�W�>y����-3�z��r�?�B?v��=D�׿���p���IMC�s���l���9׽*�v<����q�>}[���頽ۤ����s������x�R���;3��>�ɦ�>�i�=)2=�� >s��=
����1��c>���=<õ�W$�=t�y��E����)��y��ܲ�7�"��_�=������ʾM�|?��H?��+?>zC?QIx>F�>�1���>'{��?UQU>��T��Y��j�9�S�������׾��־�uc��7����	>\YK�"L>�2>�V�=���<oa�=��g=���=5쇻A"=;c�=�=���=da�=ݨ>G
>�6w?-��������4Q��Z��:?�9�>@{�=��ƾ?@?\�>>�2��q���.b��-?p��?�T�?t�?�ri�`d�>��bᎽ_t�=�����=2>���=3�2�P��>��J>w���J������G4�?q�@��??�ዿ��ϿXb/>΍�>�j�=p9��-�����?=�]��r���(?��\��iX�BB��n�5?����<�h�!�-�^�m>���=�\�������"��`
��(�>D8�<��y>f�z=�ٽÞ߽��>�A,>t�">ƈ>���/����x<lA=�;�>[w�>@>h��>^N?�&9?&k?9��>�.�����gξ
Ԏ>�=�=
	?��3>��x>J�?��N???"�5?�[�>+2�=(�>d_�>@M�vX��ľ�汽ϯȼUm�?ή�?�3�>}n�܆Q�*�j���Q�FƳ��b?�d?���>�	?P�j��i$$��<(���ֽӎ��n�i=�ZR�~G{��	=P���Ž��=Z�>��>Be�>�:�>�UV>��E>���>Vq�=���;�*�=�V=��<~Q׼{��=�뼻,2;����2^�����
{���Ի�x��sY �>�G<1g�<���=���>a<>��>�y�=�	���//>����L�-��=�E���'B�m4d��C~��/��J6��B>�5X>���0����?��Y>�[?>�~�?�:u?��>���վGQ���Me�_S����=��>� =�{;�^\`�_�M��~Ҿ�6�>���>�]�>�E�>��q�\-���*>r���a�E�>�	���T��=�[����)����}����T	??֕��(�<$ \?�N8?؏�?uf\?=�< �����>`�N����>����A:���u>w�J?D4)?��H?�)ž�H��H̾[���޷>�@I�/�O���T�0���0ͷ�8��>������оp$3��g�������B��Lr�S��>�O?��?Y:b��W��DUO����o(���q?�|g?5�>�J?�@?�%��z�r���v�=�n?ɳ�?R=�?n>�*>h���v�>��>���?�Ȩ?f~�?�ذ��k�>1	�T#�>Qɥ����>�O�>Zy>=�8>`-?�7?�?��9�H�žۺ�҉7���þB#�<��V>�t>y�R>��i>��=�f9�m��=���>+]�>��=��>���>���=5P��%���]??�`=�.�>z�??$�.>�dN<u�c���I=��5>�.���P>>`�=�."=JY-�X�q�b���=K��>ǿrb? �{<W���ҽ�>+�<�O��>�Q >9�>�^���?��>��>A��>���>\�>fy>v̽<zӾL�>����^!�d*C�!�R�Z�Ѿ��z>Կ����&�ͱ�S���	JI��"���i�7
j��:��RS=��%�<�9�?0^���k�j�)������o?'|�>_�5?������~>l��>��>B���M���Cō������?9��?�<c>�>��W?s�?=�1��3��uZ�-�u��%A�[e�z�`�b���Ȝ��:�
�L����_?G�x?ywA?�T�<4:z>8��?Y�%��ԏ�5&�>O/�(%;�E<=r(�>�,���`��Ӿl�þ!0�ABF><�o?F#�?:U?�VV�8��p >̈́.?40(?ߵd?m�?�S ?,��k?*�u>c� ?2�?�`"?��5?�l?��/>)8 >v҈=�]�<Ok��n�v��뒽R8���g;a/�=�!*=s�F��)��\�=�G�<��U��K���9��>��]�=�,E=�sn=vߺ=���>��Q?a��>�v�>�+4?$�-�Ԟ9�����kt0?9�=�C��;�l����g���(>gi`?�H�?R�[?��J>R89���=��N7>���>h>�"b>k=�>q�⽆�)���h=y� >#�=sJ�=��_��F~�a��%���AC!=��>?��>��z>E+��5r'>@:���yy���c>s�P�c��VOT�E�G���1�;�t���>/�K?W�?n��=��龏����f��*)?X<?IlM?��?4ڒ=�۾=�9��EJ�2Y��G�>:�<����Т��.����:�'�k:�Ur>
R��=�˾Wi�<�-���۾�6��VK ����2>>�^c��1f�3�����,���?[;�Zr>���E��e����㨿�&>?���<o�t�e���������ֻ�3�>�m
?�<�<m��<!NS��p����<�.?�Vu>��[���QQ��*�| X>R�h?�;s?�p�?����4���WX�/��Ѯ�-�_���?}B�>Y{6?VM�>�C�=͕���e(��>t�Dy9�7
�>4�?U��ET�b-��(�6�G���>�9?T�W���.?רF?�E�>��T?K�/?� ?�\>��5RȾ�?&?;t�?fC�=oս�FU�o�8���E� t�>��)?9UC�Q �>��?/�?�&?h�Q?��?�/>�v ��9@�Xs�>��>{W�����`>�qJ?Κ�>!Y?N��?�o=>��5���������=��>��2?R�"?��?({�>�<	?�U��p*轰�]>�?y�i?��A?E�P>�1�>�ak>�!?|��>������>�۾>��7?�L?$=z?��?9f�σ<�K�:�-��0�1�߫�ޜ`�v�=���=b�4�JB�=fV�1��=Ͷ(��\���\>���=g���64��N�>S�s>���T�0>>�ľ^.��2�@>Dl���#��Z���':�I·=��>��?ӛ�>��"�v��=a��>G)�>A���>(?�?M?X;¬b�j-۾CyK�{)�>��A?]��=~�l��o��S�u�&i=��m?}^?�W�D��W�b?��]?�g�=���þ%�b���龩�O?��
?��G���>/�~?��q?&��>3�e��8n�x��JCb��j��Ѷ=>q�>�W��d�gA�>��7?<R�>��b> $�=�s۾��w�r���?��?��?I��?4$*>��n�P3࿛p��F��J^?�y�>���#�"?;�����Ͼ/5���뎾�⾷Ѫ����0!���i��s�$�kڃ�׽�=&�?�s?�Pq?��_?�� �,�c�w%^�����V��=�k,�0�E��D� �C��n�U;�.>��$����F=�[w�!>���?�6?I�Ľ���>�׍�����)��伈>��������=x|����9=���,d��,��W���E?���>m�>�c?1�n��:�st)�1�T�K_���=�Zo>�(�>��>{�P�*��z����־$���eb$�/�u>Dyc?ЦK?��n?1� ��)1�����!��G/�=#��U�B>>�߉>��W���r&�K!>�3�r�I��4{��d�	��}=��2?�&�>�՜>X�?O�?Le	�;���y�q1��~�<s�>8�h?�)�>&�>8qϽJ� ����>��l?z��>��>����iZ!���{���ʽT&�>�>��>��o>0�,��#\��j��J����9��u�=�h?���@�`�O�>�R?��:p�G<�|�>�v���!������'��>a|?���=��;>%�ž�$���{��7����?�?�7��&����=ݪ?
��>��>�$�?��>�	w�.�&�)�? �K?�3Y?�6?e��>��<��WL��c*��T<d`�>�^>"3�=4)k>�_���A��Y^�
�5��=�`��n����'�<����ֱ�����`^>=s����j�:���}����_Ҿු�����#�wp�F��Ӄ⾜�������;���TD2�0��
Na���@���?��G�)v�,ά�t�
��Σ��:�>�ʽnD.�!��͆ �{������ھ�z$���;��HJ���h�oeO?����kܥ�E~�Ȅٽ�?4c/?�9R?�� ��3q��4=�%�*>IO��\�H>�*�m8���qٿo\��1�l?q��>Gm�vj����>y��>~Y�=���=�ӾFR��\�<�>��(?��?�U���]w忽�K���?�X@FSA?��(���쾃)R=9��>i�	?��?>91�x��.а�3��>��?R��?��D=�W�����oe?� <l�F���ɻ��=�g�=��=^���K>�>���`B�ѫ۽I3>��>�.����`>_��ذ<�%[>��нp���4Մ?�z\�kf�y�/��T��U>��T?$+�>�;�=g�,?E7H�[}Ͽ�\��*a?�0�?��?�(?Zۿ��ؚ>b�ܾg�M?GD6?���>�d&���t�{��=�8ἂ���T���&V����=,��>ޅ>n�,�ы�l�O��R�� ��=���jɿ�� ��B���<�װ��U��8�ڽ適���v����z��V��K=.g>�f>��>]he>��W>yD[?A�h?�G�>rq�=%�<���k��˾�yw�r�}�,����'�?�i���PX���ྡྷ��8��d�C�ɾ��M�տ��b��1��D�>�/�Z91��Q?�^>���<���{�6q羶���0��u�(����������h����?t�2?!%��h�I�A�|�<�N׼)�d?�<��k�K{��̃�=��_<�9="�>�T�=�䪾~�4��T��5?C�?ǲ��텾���=E���*<��+? �%?���
)�>6�>�
��`�t<�>;�>�6�>F��>C�̹����wF���t ?aq6?����@���M��>�/ٽ�������|�������mX=�{�>Z�7>{C��1(Z�ɗ�n#ֽ؉K?tKH>A�%�`��۹���	�<�_v=��]?R��>.ȇ>�o?�i<?\X�P�gP��ܾ��=�>]?نT?B>�u ��I���u��8�I?�f?��A>����c��C����?�E%?��?���͘}�H!���^���LI?Pv?V<^��/���6�.\W���>t��>�&�>*x9�Z��>�>?�"�v!��cʿ�_4�	��?�u@IU�?ŷ)<� �֎�=a1?���>��P��;ƾ�&��S����q=���>\���;�u�1���l,��8?���?���>�т��A��)�=���W��?��?&�n�g�����7x��7�7��9R�&w�<-�%>J�>s���$����۾�{�[`Ⱦ"��;.>��@j��_M?�z��������ɿa3k�a�-�6��%�?��K>]]>�FZ��@����'�\��Z�Q���$��>�>�����:��X+|���:�W�����>�z����>�+R�O����;���� <�p�>��>�\�>߮��5����?�U��S�Ϳ>`���B�1HX?�F�?�;�?/?$')<}�w��C{��n�G?_s?�Y?(�)�^�]��8��x?Η����;�����2�>�D?�i�>��)���;�w���x?c�>���@�ٿ�E¿W���3�?X��?9����>Jv�?Sl?r�(�P��������5�;�=l�=?�l=T���ʹ
�b�e���$�^��>n�?�5����[`?��^�::o��),�ȝ����>r?"��ZU�v���KL&�'sd��]��%�v���?���?�.�?u�#�%��B#?Kd�>_S���YǾw8�<�R�>A"�>qHM>/�s�!mk>���G:�B�>��?���?��?g��ӧ�2Q
>�y?_$�>��?o�=�a�>d�=O��-��k#>�"�=��>��?��M?L�>NW�=��8��/�A[F��GR�[$�A�C��>��a?�L?xKb>/���2��!��uͽ�c1�MQ鼲W@�L�,���߽F(5>��=>�>h�D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?��GP���a~�����6����=�7?�.��z>U��>��=�nv�󻪿��s�s��>[B�?-{�?پ�>�l?�o�,�B�n�1=AL�>H�k?�t?��o���h�B>:�?���)����L��f?}�
@!u@M�^?�좿�ؿ�������d��`�=�T�=�2/>��ؽ���=��3=��0������n�=zk�>dg>�ss>��P>�L=>1�)>`��G� ��(������unE�����?��%Z�oG��x�Z�����V�¾T@��N�ǽ�α��-T��/$�me���=�[U?n�W?nz?��?YE��˰�=�a���=��]�y=�߇>��4?�\D?Hv,?��=/�����e���y���pĔ�#`�>y�R>���>K��>��>�%��L>/�D>�H>�,�=�#z=�_�[�<�sL>�_�>L�>�+�>��=����Q���9ϡ�_	{��Z!�EJ>�\�?��_��Q+�K�������ھkg>�I,?|->���/b˿:g��"w7?o���v�	�׶߾3��>`9?�eC?�z=VK�i�=�2>��R��2�,�+>�9�@r6�2��/gH=>�>�)F>���= �?�"�L���B�(=��4M�>^�B?lپ='����s���F�O0ݾ��B>	~�>af�=[������R��\�f����=�^:?�9�>pH��Z������rtf��wg>�%,>9S�=
i>e~&>�s��Ӧ�����:4=�Yh>a�h>�G�>Iq>[�<&�I=�Ѿ�����>F��>H`�>K�V?c?7?v����������½wv�>�� ?	��>�m:�ډ��]�>��>��U>�?���{��`���C�>s��Q׻=��z�_�M>1��=vԇ>Q�^�� �������ܻ�~?R}���∿�WM��;kD?8.?��=:�F<��"����$G����?��@�k�?�	�H�V��?�?�?������=y�>Pҫ>�ξ��L�2�?�ƽ3ʢ�̕	��)#��S�?"	�?�/��ʋ��l� >�^%?:�Ӿ�h�>�x�rZ��|��h�u���#=i��>�8H?�V����O�R>��v
?�?�^�멤���ȿ%|v����>K�?���?]�m�oA���@����>��?gY?-ni>�g۾N_Z�z��>޻@?�R?��>�9��'�q�?�޶?ᯅ?�I>���?�s?rn�>�x�D]/��6������==�X;�g�>\\>����>dF��֓�h���j�����a>�$=�>�C佒7��2F�=����DL��k�f���>�(q>��I>)Y�>� ?�b�>��>s�=�e�����R����K?ǭ�?���I n�5��<#��=�Y^�H/?�[4?�J_���Ͼ*��>��\?J��?�[?�r�>���6:���࿿h�����<c�K>&'�>�m�>�舽��K>��Ծ[PD�Ms�>햗>�$��a7ھ���������:�><!?3.�>S�=ۙ ?��#?��j>�(�>BaE��9��W�E����>آ�>�H?�~?��?�Թ��Z3�����桿��[�x;N>��x?V?qʕ>b�������LkE�4BI�:���]��?�tg?pS�/?<2�?�??`�A?{)f>ه�*ؾi�����>�?��-��<�2�!��Hགྷ�>�(?�D	?C{޼弬��U1���6�n�;�L!?��V?��+?n�����t�Ǯ���br=�?���1<$ýɓc>P1>j/->e����\�g��=t�6=4��<�>�ue
=��b=UxJ>�;�%Pq�6 >�"?:�;�{y�U�=��u�k;�5Aj>��e>�(��}g?E�� w�#O������a=���?D��?2��?�8ݽ�h�cv@?9�?q?e��>�;t(��BǾ��E��h�S����_=X[�>��1=8����������C��53���SF�b3?�u�>� ?c9?Z&�>xԨ>#$����8��Ծ��޾��n��l�$�o9E�}�6�4���AV~�@�v=�8��]|�F9�>�c����>�?�(�>��>[��>M�<%�>�[>9a�>#w�>�>�4j>Kq>2�:P�{�zTR?����ѱ'�������5"B?&vd?��>��h�������P{?燒?�m�?d�u>�h��2+�!h?�^�>���h
?�%<=�I���<�R��^s�����������>~�׽b	:���L�Жf�9f
?�%?We�̾6�ֽ#���L�n=N�?��(?��)���Q���o�иW�#S�x��[6h�Jj��5�$��p��쏿�^��%����(�_s*=��*?a�?Ì�4�!���&k��?��df>t�>T$�>A�>^uI>��	�^�1�X^��L'�B���dR�>r[{?v`P>�iL?VS?'�w?j�Z?]�<>�z>��X��>k��=���>Y��>��=?C?u�;?�?�=?��=9���������`��>�?�G?d?_"?�y���.����=z�(����[�=�~<Re���Žl�?�l��=v��>ݓ?�ͅ���/�[j��)(>M4?���>��>��� =���@l>7?�>f�C��	�>q���C�k����qF?�{�?�?Q��;by�=c�=:�B<�N��л�=ܼ=S�=}��<ʻ=��(=T�=�;u>�ڜ=F��<)N��~�<٥�=:?�>0�?rH�>���>*���Y �~�>�=j'Y>d�S>N�>��ؾ�`���%��;�g�r�y>�t�?�g�?�e=���=�T�=�R����������&��.�<�?�0#?�+T?���?�b=?_*#?Њ>���?���B��rߢ�)�?>�<?�[>���EѰ�H����'��$?���>��h��6K���/�H�����9<�f>#�]�~���焱��$�\9>^L
�*Fy�W��?��?�����2�$M��$��]��01V?.��>���>�$?�(��aj�����[>,�>t"]?��>��?;�?�T�?��
?�[����ٿG蟿Pe��ń��!1?��?�Y�?��\?f�?$�n>_�<��(�� �w��h����"��#�>k�J>���>o:�>k�W>��>FH�>�^+��md����\����$�>e��>o�F?���>F�=a�#?U��>�V���������\��N�]Hp?�/�?%- ?�8Y>P��I�}�sz�>%l�?�d�?��?H�l��|W>�r���)�G8����>���>�I�>�+z�V��	���v�>�B?sq��9k%���^�J�h=r��>O:B?_�>W���p�ߛ��E��%���7M�HWW�V<���&��u!=�����n0���-��������v�<P������q���U
?@P�=|��=��z=������`�H=�[ >ƙ�<q�b=���z�<[�N�/*<�I�����[Fj=qYX<�25�|�˾"�}?�FI?��+?x�C?��y>>��4�?��>����+?�V>�yO�����[;�ꓨ��픾��ؾd׾h�c�ן��0>�H�O�>m,3>��=�v�<�-�=os=��=�6O�fo=���=��=E��=rG�=> M>�6w?!���沝��4Q��Z�v�:?�8�>�}�=W�ƾ�@?��>>�2��|���=b��-?X��?�T�?�?�ti��d�>0��㎽<r�=𵜽�=2>��=��2�*��>��J>փ��J��؀��{4�?��@x�??�ዿ�Ͽ2a/>?=�=)�#��xC���l�յ���V$=�-����G?j����۠����U� �O*��*&>���>�ص=!�><t�f���ѼE�ʼ Q�>Ty =E�> =\>Ad=N䓽=�B>�%>69>]bV>eМ��EI��Uh��x���6:>�= ?��>d��>t�?��0?��d?�ĺ>�|n��{Ͼs¾E��>FK�==��>@G�=��C>)ͷ>�7?��D?�.L?iα>;2�=���>�K�>�q,�9&m�_)徱����;�<R�?���?���>��*<CHA��7��'>�;�ƽmK?�\1?�?��>�Q����]W&�.�.�Ũ��C��7��*=tBr�<�T��������U��d��=�`�>a��>3�>&Ly>F :>ϤN> �>x�>���<�q�=]����c�<#���ה�=�����:�<�ż�\���&���+�Z����<�;��;[�^<�q�;�M�=���>�2>���>��=�g����.>����(M�q׿=�E��rB���c�Y~�"D/��9���@>�BV>3��$Q����?�X>��>>R��?^�u?�">C�	��?վ����`�(U���=x>��=�%�:��X_���M�ܛѾ��>�>�>��>���>v�ľ�=����:!$4�}�D����>�U�Q�O=/?�=~.��M����俿��������1LZ?������>L?��4?�{q?[�>���i!ľFrm��?���>;�V��e���xE�T�&?Uj?�u?]q��k��e̾�h��ʴ�>�>I��P�������0�xm�����r�>j���о�)3�gl�����s�B��5r�D�>4�O?4��? b��Z��KO����Ӆ�r?~g?��>SB?q??.᡽�g�T���%v�=4�n?��?�0�?
�
>�:�=�?��Bj�>�?&�?�3�?��q?��?��F�>kV<l%>�藽���=�->꫊=w�=�j?uL
?˩?	ݝ���
�T��.�� �X����<0Ҥ=�C�>聋>n�u>v��=�B�=U��=@�c>9Þ>�Ӎ>0�b>�֥>p�>%P��1�ʾ,??���=��?��,?�t_>*x��f�7<��B>��=�Ը���Ǽ��>h��􂍾|�L�C��c>+I�>^տ�A�?��������w�>پ����m��>p�>$�@��;?���<*�>|/?���>��">�C�>Cy�;��Ҿ�>����I!�C�B��SR�v-Ѿ&�z>�I��(�&�����}��vKI��괾Y)���i��6���\=�T�<�4�?����F�k���)�k���>~?Z�>��5?��Q��Cy>�$�>[W�>�6�������捿5��!�?��?�;c>��>I�W?)�?��1�03��uZ�*�u�Z(A�e�O�`�|፿�����
�Z��*�_?�x?'yA?�R�<:z>F��?��%�Eӏ��)�>�/�';��?<=l+�>*��S�`�n�Ӿ~�þ�7��HF>��o?8%�?|Y?(TV�>m��'>��:?
�1?4Et?��1?h;?t��5�$?=�3>�/?B~?�@5?�.?��
?_*2>��=6����)=^E�������ѽLʽ��񼣤3=+|=�fT���<��=��<q��o�׼�\;� ��O�<p�;=I��=���=Qރ>��V?��?�{�>�
>?��H�D�;�h<ݾ�y-?#t>䓾��j� ]B�{+�f�6>-Db?k԰?�R??%B`>�<E�Ia��E�=Đ>;�>�@> y�>ա��v���$5=�w<�>b��==Y������򾁗A�x"�=�}>�y�>?x|>؛��%'>(؟�׺u�,Yn>��L��N��:�Y��CG�Y21��4u����>�L?��?V�=����Q��b5d��p&?&�9?֡J?�s?���=�$ܾA�9�~+K�|�&��0�>�.=�
�쥡�^���U=�>Ql��u>(w���ET>���#@վ����C�cվ�/>Qp���V�<8��J!޾s��0�<�(>�n��l]�߯��a񥿋�B?
�B=�����V������,@>ɤ�>f�>Ԡ���iɽ�29�'V����=#��>���>�[��� ��I�����>YoZ?$:�?�m�?y����b��og��R��BZ4�T2@=x!?-�?n�>eS<>S����j�Y�3��*g��4��ͭ>p��>�K�������Ш+���#�h�>}3?�ߜ�3?j�$? �L>�Y?��R?xV?�)>W�#��Z���1&?d��?ȣ�=��Խ��T�+�8��F�.��>�})?��B���>s�?g�?n�&?
�Q?��?��>� �26@�Ku�>�_�>�W��Z��2�_>֧J?��>�@Y?�̓?M�=>W�5����jɩ���=}�>ӻ2?�<#?��?�ȸ>��>���c=��>�!a?���?m?9��=�?��#>��>�Ț=���>M��>�M?�%M?o�t?=�L?��>ڒ<�W�����n���1�=�:��1<��i=h���c{w�����<8F<����eB���s���R��`���X�;�'�>�t>w]����/>��ľ�爾�UA>]������L��R�:�;�=�I�>�`?�W�>��"��^�=d�>*�>p���N(?��?��?V��:f^b��J۾�I�e[�>sA?��=tm�kh����u�ޮf=tm?!"^?g�X��:��E�b?��]?Jh�=�.�þE�b���]�O?�
?O�G���>V�~?�q?A��>��e��9n�1��"Db�F�j��ж=]r�>X�#�d�_?�>3�7?�N�>�b>!%�=u۾��w�bq��C?k�?�?���?I+*>Y�n�I4��?���H��\OY?���>������!?w��@�˾s�rK��F<���[߫���������!��+����ڽ�=YX?xZr?�4o?X�]?9&��ia�Yp[��r}�&�U�E���o��IF��RE��D��m�����%���-��%"A=�0��w^4�϶�?^�?���<�5?ᆚ���������_>����FԼ!hE>�:c>Ξ�;�������ƽ̿��e�!?A��>�1�>�-i?����K�|�a���V�W��6�>|Je>o��>h� ?�8�9"��x+����(ؖ�*d��+�p>=�c?/UN?C"p?.���	=4��4���'"�W�{������DB>�m>�8�>[�T�ٸ��X#��?�ƞr�6���U���X�@�x=��0?�W�>�
�>��?��?`b�=p���Ln��/��Ψ;��>iCj?zw�>p��>�2ͽ����>�l?���>��>����X!���{�o�ʽ;'�>]ܭ>̵�>��o>9�,�H#\�4j�������9��s�=��h?����&�`����>IR?��:=�G<�{�>��v�˼!�M��N�'���>�|?���=�;>�ž%���{�A6����?7?�@���)'����=zo?hE?|��> T�?W!>>��"�!��>��=?�i@?�3?QT�>uN"�����Pֽ,̶����;�ܬ>�JF> ,= Ht=?	�6r����n�qt�=]�)>�%�=�<�/ϻPn?����n<�,�M>m�ӿ"�|������̾����`>�Q�����c=U�����=p����SN�`lg�1��S���ݽ ҭ;Y����9�gV�?�ͺ?�0,���K<o����KG��`̾�d�>�aX��7�=�a���h�4�#�q��)*ž�Ҿ/��R�����!?re�������l�����
�T?~�*?.�D?�ķ�� w����W�]>롢>�G>�9��K��b�οA��}?0M�>��+��޴�8P�>��?�E�>l,y>�+�a�x�(�>�ƙ>.�3?�)�>���嵿ӿKA˽\r�?2	@�ZA?�)���.i=���>�0?��C>��3�c�@4���b�>۞?&n�?��}=m�X��zU��zb?+ݳ<��@�&r��5L�=���= =���MDC>= �>��"�y�A��N���6>}W�>-��/��r�Js|<~�a>����h��&;�?�:R��*b���4�y;���.>k�S?z�>�2>W�&?��B��ο#P\���R?A"�?$S�?��%?Z���41�>z�پP?�5?0��>�>'���u�;�I=>�`;4B�=�Ѿ�2V�G`)=���>	>�k"�G�	��5L�&��Y�>д�8GɿΊ'���
��ץ=t���wʽ�*u��dν�.�<�kݾ�b��4����<]��=O�T>���>f�/>�s�>m�^?m�X?T�>�h�=�l �q;{�U�����=�Ӄ�qpڽ79�+JʽF���* �vrʾr뾅��J���'����+����זY�'(��3�(���M�s�5��	6?6޼=�0���@�J�J6۾����f.�W)>;>磾-�-��[��?�R?��m�� F�:��vͽ��<�=4a?�Θ�6&�b����=_�ڼ��T� 2�>_;>�~���Q*���M���-?6�?f���Ry޾��7>O�]��3>�:?��?`B��?D�?;����ͻ>e�>��>F?�ɇ��I����8���?�A?Bsd���@����>�U}����_6�=�_���z����=�}>l�;=1&W�s���Y�9ʲ=��K?�!�>
"��e�1	�����;@��=�m~?9(?F >j6f?��1?��=4Ѿ��C�Q��!Xk=�lA?zJW?`D>�ͽ�оw"���&7?�gT?Es>����r)�y$<�����:?U	y???F��p����ڞ������C?��v?n^� q��,��0�V�v7�>
X�>ۿ�>��9�p[�>V�>?� #�8F��5����T4�Y��?(�@t��?)`:<��c��=�6?7V�>s�O��<ƾ�~��Ă����q=��>�����]v����(D,�Ղ8?���?��>����ئ�j�K=�z�:�?�Ƒ?C����	8='@��B��!�3�gxZ>����	��=�߀>�׶��=8�o���� �m[��ɣӼ�}>��
@7C+�"O	?���G~�5q׿ħZ�$�T�:���%?�^�>V��)����g��-����\��ce�'Ѯ��$�>��~=K��x�t�.?t�Q`9��`�gB�>@��_@�>��K�}$��Z-�����;�Ѕ>I��>��>42ý$�����?����խϿ�����0
��Y?�?��?�?�<��z��m����(�ݵ9?�b?;V?gp��<.P�]�?�\�c?2�z�Y*��Q�Z�ݾ���>��B?��e��e德 Z>]C�>h%?�L�>z����sݿv_ѿ��ྼG�?�E�?�o��f�>nk�?-�?�b9����4ƾ`�=���=b�O?���>
aپ��M-r��׾��&?T:?=O-�o[�2�_?j�a���p���-�L�ƽyۡ>��0��`\��M��֥��Ve����f@y�E��?�]�?3�?f���#�'4%?8�>�����8ǾE��<���>�%�>�&N>�W_���u>w�F�:�Ll	>��?�}�?i?b�������tX>5�}?z$�>��?�n�=;a�>zc�=(���,��k#>g$�=��>��?^�M?�K�>�V�=��8�N/��ZF�pGR�g$�,�C��>��a?ÂL?`Jb>���x2�I!�sͽ5d1��[��X@�C�,�}�߽(5>�=>>:�D�ZӾ��?Jp�4�ؿ�i���o'��54?7��>�?��w�t�����;_?\z�>�6�,���%���B�c��?�G�?:�?��׾fR̼�>(�>�I�>0�Խ����[�����7>2�B?i��D��r�o�W�>���?	�@�ծ?bi�V	?W!�Q���_~����Y7�}��=�7?D0��z>W��>��=nv�l����s�߹�>�B�?�z�?���>�l?��o�-�B���1=�K�>Ɯk??t?��n���y�B>�?7������oL�f?��
@�t@��^?��g俪V��i	ľN���t�*>0�M=U1�=����� �=�r�����ϔ����=n;�>�^>=>�ea>I*>>�;,>�����#������џ�p.����X%�3�r�"_���u�����.��ξ.�q�z��2��u���P���T5�~b�=��T?�#[?�r?��>䮪�&�>�!��h+�:-3��ֲ;O��>o�@?q�K?E�/?-��=tЖ���Z�Կx����x���<�>+#>�g�>N��><�>��<.�C>�|!>C�`>y�=��`=/oF<�ȓ<B�0>�л>��>cC�>]eb>��=������������� �������?W�o���J��Z��6ߵ�{¾C=O�<?�M>.፿� ο�T��Jl<?-|���;��5zq�c�>+5?Khe?q�i=lվ3��jvj>F��p�A�}	w>�[9%��M�C��|�=��>̔�>�[�>�$���@��r��P�X�>O>?-��=d�
���[���m�����������?Z�J>�4⾻=��Vg��H�a8>�w+?�?�UA���޾rT����$�>��K>k�$&
�Fa>7b��T9�Oza�c�5<��k=¿�>�R?�">��)=]5Z>���,�9�~ү>iW>�}�>��?�D?�Ï�7d�򻓾g��N~>-]�>�c�>��I=V4V�v��=��>#WS>�lҽHE��4˽�n��.�>��d����X0�Ս�=��۽N�=��=R$��n���?=j�~?���S�����'����WE?�p?���=�WV<	"�	���"���p��?�@!h�?L���V�$�?ˎ?���	��=O�>ͫ>�^ξ� N�:6?��ͽ�/��i��4!�{��?)��?��%��k��Ϡl���>�&?_dѾ���>�{��$��چ�;.u��^-=t�>JH?,���]b�_>��3
?dy?h}�U���A�ȿ��v���>?��?v֔?*@n�T��?�?�?�>O��?�UY?{�e>,*۾OW����>�@?�FQ?�>��\+��2?�?;�?S\A>���?��v?�>�G�:�6��ƶ�󅋿ӣ�<]��;z��>U>����@B��ݑ�	��^l�_�x	W>ظ$=�>�����}��=�7��m,���E���>� d>�\X>�_�>	e�>._�>���>��<oǊ�se���ݕ��K?%��?����3n���<���=Z�^��&?1F4?Á[���Ͼ<Ѩ>��\?���?0[?Qi�>,���>��翿�|��0��< �K>�-�>�D�>���,OK>��Ծ85D��n�>�Η>�֣�>Aھp-��᡻TE�>�f!?s��>5��=ڙ ?��#?��j>�(�>CaE��9��W�E����>֢�>�H?�~?��?�Թ��Z3�����桿��[�o;N>��x?V?qʕ>a�������7kE�EBI�?���]��?�tg?�S�/?;2�?�??_�A?u)f>܇�.ؾf�����>�6?As��g#0���Y��qѾ�n�>�a2?���>�\���=��>�����ξ�5�>��i?�e<?E�[�Q��bu��T�8 F�q�:S�0��=�=Az0>��>X0��	�=�C�=�Y�=�J�O1'�餶��%H=��> D->>�<c���(5,?��C��Ճ��^�=L�r��XD��>+�L>�����^?�l=���{�����u��M�T����?ܝ�?�a�?4I����h��-=?/�?�?o��>N.��ge޾�b�K�w��x��a���>%��>�g����o���싪��J��b�Ž������?�0�>į?�*?��>�`�>�����~(���Cξ�ǀ�9&.�j�/��DP� j-��X���:!��>�bɾu/���HN>ܰT�Yv?U�6?��>T��>=>a�D�D��>���>9`�>�?'\�>��>0%u>-�S�}���MR?����v�'�n���>��gQB?�pd?��>TIh��y������?���?�z�?�qu>�h��4+���?9��>9��\
?,�:=r��#G�<jf����x@��]�3�>&�ֽ=:���L��#f�i
?��?�����̾�Lֽo���f0q=�[�?�)?C�)���Q��o�o�W��LS�9���h������$�چp��ꏿoT�������(��)=�m*?��?y`�ܔ�𬾚Yk��5?��6g>��>�>w,�>8�I>��	���1���]���&������>{?�`�>+/J?[�C?ΒQ?��D?~�>��>.���=��>��=�ς>�O ?��F?>0?��1?�4?>t,?�+f>��ս�3���ʾ6�	?y ?)~?� �>* ?/���X�������Ú�pBv�	n����}=�����ڽL����B�=k�t>��?� ���6�ځ���`y>��9?Z��>g3�>�H���Y~�8x�<̇�>G�
?䃘>�U���v�u���>�ڃ?gl���	=�*>�=Q��6yJ��{�=�?�t|�=���;����@X;�I�=��=����N��c�<:��<pN=*��>>L?�C�>��>�=��Z��!c�d��=�Gj>_�>>�>0��ʙ��K���[d�s~v>,��?p��?}0H=#��=�|>b����,�����{�ۍ=x�?�q?�@P?���?7:?W�"?<K>��AǑ�����7���A�?%#,?���>���ʾ1稿�w3�ҟ?�P?�3a����l8)��y¾ҸԽ��>ya/��<~���� D���y�������h��?廝?�A���6��q辽���8X��>�C?%�>�M�>o�>y�)���g��)�eU;>o��>�R?e�4>$_?c;�?�]�?�@>����?���Ӓ�m+��f��>�g
?�B�?�ט?��~?��?s�>�2E�K,��'�ؾ�@����J�@4a�1�?�<���>�8O?��g>vσ>I�e=�̾�L����>�>���>�,�>�?cM�>�B>f�.?���>�K�� C��h�����N�=�e?�d�?��>2/»E7��XH�7/��>	��?e�?6?�a��+��=�n��B�ξ`���u?J�>�5u>g��<�פ�M��A�,?� ?�7��"�پT�?�9,׽;�?�9P?��:䛿\š�w*�,��=����y���I�P49>�X��*��>����Ž�¾�k�rj׾���?�oꖾ.�0�1�>��h>3K>���n�@��=˟=����m��Pd�����b��W���`#�<�>�;=ٽ5�o��v�<Ζ�=m�˾��}?`:I?�+?��C?�y>:>c�3�J��>5���B?�V>�P�/�����;�(���g���ؾ�x׾/�c��ȟ�G>�jI�*�>963>�D�=L�<�=As=���=R��= �=wN�=&b�=���=;�>T>	6w?ɚ��ز���3Q��k�x�:?�8�>���=/ƾ@?��>>�2��G���c��-?���?T�?��?�vi��d�>����ݎ��n�=@���A2>��=�2�ɣ�>�J>8���J��'��$4�?t�@��??�ዿi�Ͽ�[/>�ү> ҆=S@�g�M�QŽ׏��>��Q��>�Z��!��x�-?2o�=E5��9��pl=p|>ƕ�>u�,>��c�?)�=ed�RNO<�����F>�>t�=hꄼe�*>p��w-�=��S>����t&=w�=�v��`R�<HAO>���=��>�?6ZF?�c?V˪> ���nBþ��ھ3m>�I>��>�st>�ѿ>���>[�4?�@?p)]?+g�><��=&��>2��>��*�=�Q�K�Ͼ�����\Ѽ>Yj?�@�?ȥ�>��<�9H���/��J@���Y�U=?��=? �?Q
�>L�D߿M�j�.� C�<�>D�X���B��b-��y������a���2=	�>s�>0O�>�*�>��W>���>-��>���=��6=Q��=P9<�	ռM�#�'A.>��һ�}�=�M��]y�=��5��+��.~��P=ϩ%=�em��h	���H={}?{FP>Y��>��>/������=�о�=�2?�=L����O���x��J��	�I�(硾��	>��m>��#=G!��O�?��T>gb1>D��?v0}?p�#>Sl=$�
��R��o�e��ڳ�b=��@>|�P��qT��_�U�����>�}�>��>R�>���Õ=�BP�<Oc,�Nj���?�[:���9�`�_�����d���k ��-"I�P�>>l?�E��D8�>��~?��5?�݋?��>���_����F=������Խ��?���N!!��b?*/?��>4G(���j�z5̾<#��xd�>�I�i�O�𪕿\�0���淾���>O���Z�о#3��o����WB�r�먺>��O?��?�a��?��MO�����ᆽ�g?'�g?[*�>??-?0K���p�����;�=	�n?+��?�?��
>ʍ�=5���<M�>"-	?Cޖ?���?�s?m@��h�>�K�;� !>H���	��=�>�(�=
��=�0?P
?�A?�Q��� 
�3K�&�\���=���=L�>D��>��s>%�=�r=�ͧ=5_>n_�>�9�>�g>僤>bv�>��߾��ؾ
B'?��>�?DT?W"�>Ǩ��L���{�	=�l�Y��������$>{���x��o��=pi�=�z$>��>r<ѿ9�?�^;��ؾ�Z?�ʾ~ ޽�b�=�gm>V�žI0-?��>2\�>�m�>�H>:<*>oD�>1c��VѾ�L>�F��< ���B�*>P���ξ %�>O��VY7����h��s.>��屾��/i��	���f<�T_�<%��?b!�!k�cn(�&��j?���>��2?;(����v>f�>�$�>���gܕ��׎���_��?Z1�?ڤb>��>x�V?~?�3���2�B Z� �t��A�uWd��o`�֍�8����M��.����_?)hx?,�@?��<Q�z>��?.%�3j��6��>�7/�6�:�@I=Cϧ>;5���n`��?Ӿ�yþ=M�OH>d�o?��?�?TW��*o�((>��:?��1?�t?��1?~K;?TU���$?t<4>�?f�?c5?O�.?R�
?�p2>w��=o���+=���������ѽɝɽ�#���2=��y=�&�<�=���<�~�L⼤��:�짼�J�<G�:=�?�=���=�n�>��a?��?h3�>Ņ%?i�A�#�,��ಾp(0?���=�����J5� q�W��~�>VFc?�`�?��S?��|>M�5�������=ף�>�� >�R9>+6�>~7��l���o�L=��>���=�6�;	uԽ!���o���<�s�X�<C;>���>D�|>GW���E&>3��Cy��ae>a�O�k���T�ǩG��2�6�v�ɋ�>��K?��?���=������)�e���(?��;?M?8[?�ʔ=$�۾�c9�΅J�<9�~��>��<��܃��3����:�y:��s>�a�������]>����޾�_n�RI�y羧�V=7��Z�Q=_��5(־Mc���M�=��	>Ș���V �h��������I?]%f=I���W�����J>6̗>窮>)�5�)gy��@�/���H�=4�>�<>՗�����{*G�6Q���=l��?� �?���?3�n��Z}���x:������
��=�>�(�>�?��>*Vz=G䞾P��z|��| �o��>��>3sA��r��<	�)��h�pw>�T?5>�R'?�?O��>�Pj?Ol�>�e�>��>c�:�[蟾6A&?���?��=��Խ��T�i�8��F���>9�)?T�B����>�|?ڸ?M�&?ÄQ?ɸ?��>.� �%B@�t��>]�>L�W��]����_>\�J?S��>>7Y?2˃?B�=>�y5�uӢ��|��7b�={3>�2?'#?H�?���>��>)Н��r=J�>ZvX?�%�?�x^?��>ɍ?{~>���>$�= ��>�e�>2R?lR?��w?|�I?/��>��~<Z����3���o|�����6=w�=Y,�=��Hf���G�PDQ=�,��GR���ȼ]B�8�9��N��V�O<���>�@r>HՖ�2�/>�qƾ�S����@>9ܘ�qX������7��X�=��>!^?V��>r�#�!��=�ʽ>���>�g�<(?%�?-?�O�:�hb��cھuK�C��>� B?�(�=��l�g��5�u��f=VFn?	�^?�-X����F�b?��]?h��=��þ:�b�}��|�O?=�
?{�G���>j�~?C�q?X��>��e��9n����Cb�!�j�OѶ=vr�>IX�C�d��?�>e�7?�N�>,�b>$�=yu۾��w��q���?y�?�?���?�**>n�n�G4����4>���0^?�[�>�̦�#?5���>�Ͼ����q���kO�;���������7��z*%������f׽���=��?j	s?�bq?�`?� ���c��R^�#��sPV�#"��T�q�E�:�D�}C���n��N��L��}���xD=/����*7�㟼?HC?�=��S
?�d�x�4����V>��оr�=b�H=X�?< �<i�\�|zC���?�;U���?��>��>�nz?�w�3�2��eR���L�9!׾8f>_�>ck�>Q�>L�/�0��� ��D�M�}�ji���u>��c?d�K?��n?���M1�j����!� %0�h����B>!�>���>��W�2v��'&��M>��s����_��F�	�x}=��2?^i�>��>E5�?�?UN	�����({w�Mx1���<�7�>��h?�F�>��>�нV� ����>w�l?Ϊ�>�>����cZ!�!�{�l�ʽT%�>[�>:��>7�o>��,�`$\�k��p����9��v�=X�h?���V�`���>MR?�Í:9H<u{�>snv�M�!�F���'��>#|?�=G�;>�zž�#���{�8��>�?;��>u��8+���=���>F��>��>�Ǉ?|��>��Ͼ�� �Ý�>�A?`??��??�>��C=� �y���c
��e<���>��[>)B�=�B>y���cr��񪽭�=F��=hN�<� ���*=��=��x�p<KU�>n�q�h������?���Ҿ�B��:Ԫ�u�_�W;/��Ȅ�춮�(w˾9ݪ�y/m������@��a9�8<4�o:�g"�?'u�?w%�{��7����2P��f��6�?�b=�
���>T�X��=���7�s��q4��Q���&��^H�s�7?Gi��0���i�'�$�??N�A?xND?p���z'��{;�D�e>Ά�=��>�پ�U���6����w}?j�>�&��h�Q��>
?�O�>��>r�P>��&���J�2H�=`��>��8?�d?\t��
޿q[ڿ�A�=��?�"	@^�@?P�3����&=��>a�?d�L>�s�7��`\ž�l	?Yǖ?�?��潲tJ���=�m?�=p�O�g��<�'=���=b
��X|P<nJ�=�n>I�=�ф4� -ȻT_H;z�S>�+'���<��R���=9,9=�U�����Ԅ?�y\�.f�ݤ/��T��`U>��T?�+�>9�=��,?47H�I}Ͽx�\�_*a?�/�?���?��(?�ܿ��Қ>H�ܾV�M?}D6?a��>]d&�%�t�xt�=(ἜQ�����%V����=ԭ�>E�>v�,�b����O�\򘼸��=��� ʿ��%�΍�:��<�4�Ḓ����Ƚ �ٽT|��}p������wJ)=/��=�@K>�,�>��d>\RU>��c?u�p?�K�>�>*���i��¾p'B=:�7�oF ���Q�ԽlY��^��@о��������@,ƾ�DL�� �Y�^�M���Q$�S*L�t@�1\-?dq>>�4�g������ξ1xI<����d����ҵW��?�):?]����\�s�+���Y=)T����S?9��m��>�x�?n0>s'r<x��<�>԰;iUվ�[��@D�/�)?8�	?���������=����|�<��0?ݙ?e��=��w>�?��a�/�D�#�">qK�>�-�>u��>�{�=�ڡ����u� ?�"5?i#0�w唾���>*���QL�p��Sk=��t�b2��kn]>�
�<���[Ô��5��ꗼ�W?���>_*�F��δ��-����==�x?�:?J�>�lk?�B??B�<W���h�S��j
��{=vW?bh?�>4����Ͼ˧�v�5?�e? �M>uh��;龁N.�&��ĺ?��m?��?�S��1}�{4������5?�Ac?�a��Ƞ����.龪ظ>r9�>��?3�$�`9>+�z?\ݽ��[�Ձ˿`y����?kH@�^�?�W���3c=�S���>�\�>��F��۾U]�奰�lʽ��?�Q����M�4I�j�a���?D��?���>S~ӾH�/��f=���ù?v��?�#w��=�T'�4����0��r�=�K�S� >�=_d���C�	`辻$��D��܏I;!>Y>��@����/?����C��@濧��o
'��y~�҇	?�>���=xz���*�>+��I�h0O�Wz��ɣ>m�>堚�������{���:��'���+�>��6�>��Q�}���T�����<���>�G�>��>0�����5s�?g����Ϳ������:�W?dמ?��?�?�>K< �z��t}��ha��TH? 4s?��X?n�9���]��>��i?ڽ^�ʚ=�4�ܾm��X>�U?]�
>+�
�M$A<F�@>rq ?�n�>�������ҿ\���?��?�����>R��?� �>g�/�8렿����<f�ŭ�=��E?��f>�|��R�.Hc��3۾v�>]>?��Խ�K�ŷ_?��a�b�p���-��ƽߡ>ʳ0�1O\��s����8Ve� ��S9y���?�\�?l�?���#��3%?��>����:Ǿ
�<1��>)�>�.N>Vq_�٦u>+���:��q	>Z��?�{�?3h?Õ�� ���Q>��}?�#�>�?u�=�b�>�d�=��t8-��h#>� �=z�>���?��M?vL�>`U�=��8�d/�2[F�HR�#$��C���>�a?b�L?�Lb>�"��.$2�%!�sͽUf1�N<��W@�A�,���߽�&5>��=>V>��D��Ӿ�9?���~vؿ�&���;/�O�4?�[�>�:?���[Rz���Y���^?"f�>���D��ދ�fi �ի?�l�?�	?�r־��ͼ�C>#�>)@�>�&ҽ򽝽U���vs9>"RC?��{I����o�9�>~�?�@>��?
+i��V�>>�������r�`/��ꕽ��=�:?5$���B�=�l?��=
�K��w���P�e0�>;�?�E�?\��>�h?CGX�x�/�w�=��>�5L?H	?�;�<���Sq>+=?{ ��ro�����lF?�
@�@�8?$Ƥ����G����¾��^ '>%Ҽ)*E>Cϩ��q>������k���!>R6�>��'>��d>q�>a�J>��#>�����*�/鱿�w���,�LI�����i`���Q��D+���龉jӾQͽ�<z�_*�>%%�FaC��=Žld�=±U?�R?�0p?� ?Jz��>m����l=��#���=�\�>�m2?R�L?Ҩ*?���=y[����d��P���:���χ��N�>�(I>+��>~l�>BT�>O��9��I>| ?>~n�>j� >��%=����= �N>�U�>���>d��>�=>�>������#1h���t�`�ǽ�?������J��𕿋���b���?�=]t.?ީ>���Bп곭���G?�����%��v+���>ɝ0?�?W?@o>1����DR��[>�)��Bj��[>/ �t&n��*�l?P>H�?�a�>& �=,�	���e���G�HT���>�g,?�5k�6j�>1r�pSz�C*'��D�>��?�b>o��F��*���ԔH��/>|B3?�ʭ>2O����l࿾[��TS?�`�=�k�0���-��>�N^��kU��E7�<��<�³>&5e>�?5�y=2暽RÕ=�����m��>�˖>���>ȑe?i�>��=�4ʽ��þv@E�<D�>�&?X��>�N�=�)��!�=�9�>
v�=��HG�<��B�̵�@YI>Ӳn��q�������0�,d �.�==r*p=���������<!�~?`��䈿��a��mD?�+?���=_�F<��"� ��zG��!�?J�@l�?B�	��V���?A�?�
��۷�=�|�>�׫>>ξ�L��?(ƽNƢ�Y�	�L'#�AS�?��?p�/��ʋ��l��9><_%?K�Ӿ�e�>+~�aZ��u���u�#�#=/��>?7H?^R����O�l>��v
?7?G^򾲨��A�ȿ2{v����>Z�?(��?��m��?���@�%x�>Z��?VgY?�ki>#e۾-`Z�ӎ�> �@?aR?n�>-;��'���?�޶?>��?J>�Ȕ?.�?f��>+�h=7��}������l&=�O���mq>/�+>���`B�����YɃ��e��"�>U>��=��>Z�������|	>��3��~��'�üö�>].>�I�>���>6��>��>�1~>�b�=� �˃�d闾��K?��?����1n�R��<��=�^��+?�M4?s\���Ͼ׾�>�\?}��?[?<i�>8��B:���忿�w�����<F�K>�2�>�D�>�)���JK>Q�Ծ�9D�\p�>9Η>�z��1ھ�.��y���}@�>�]!?��>��=ۙ ?��#?��j>�(�>CaE��9��X�E����>٢�>�H?�~?��?�Թ��Z3�����桿��[�t;N>��x?V?sʕ>b���񃝿vkE�:BI�:���^��?�tg?qS�0?<2�?�??`�A?{)f>؇�)ؾn�����>C)#?ᐠ��*� �4����S�>�u?��*?�4��ӹi�v�m��3�KDA���?��??�`#?����_��Y:������� >=��<ь�?_�=/>ǰ�>?� ���Z�3��=_���fm���ؽ:�5>jX�>���<����9����e=��+?t�M��Ȃ��+�=�yr�JBB��t�>�nQ>Bf���u]?�@��z�����W���zU���?�X�?��?)�����g��<?4=�?h�?�C�>mg�� c޾�޾xOt�������r�=S>�>p�6���������W�����ͽՉ����&?�_�>�?�+?ܧJ>���>ɇ���/�d��Z��Y�d�f��y�)�@�V��&������P�Wc+>�#̾���&�>1S �lO�>Ғ?t��>wo�>R�f>?��P��>��g>��z>QE?���>P�>�"p>��"��ؑ��JR?R�����'�ٷ辛���q3B?�pd?�2�>�
i�z�������~?���?�q�?�>v>n}h�/,+�o?�;�>���mp
?SO:=Y
�R%�<1U������5����ᫎ>�:׽�:��M�of��h
?7/?�����̾�8׽���Plu=gp�?*>)?W�)�7�Q�%p���W�<�R�=v��i�Ⱦ���m$��vp�~����F�������(��S*=MM*?��?"v����8����yk��7?���f>&<�>��>c��>[�H>J�	��1�0�]���&��{�����>��z?U0>j�>?O2H?$΁?e3\?6 f>?�>d���0?J��և�>?�
?�_0?��S?�RC?�$�>�O?]�4>��|��������$�>�e�>f�(?��A?��?"*����ǽ��4=����0��0ri�C'��!(;�Dۗ=~>ν��>��>�S?���n�8����4g>�15?���>���>v㎾�Lr��
=��>c�
?��>u���,�n�7��+��>D`�?�B�>=K�$>5#�=h����ϵ:7��=�Sü*D�=��6���6���<���=�d�=우�t�x:j�[;�%�;5j�<�u�>��?$��>�<�>w@���� �Ѵ��x�=�Y>-S>�>5Aپ�{���#��Q�g��jy>�w�?1x�?I�f=u�==��=	|���R��v�������r�<-�?E#?�QT?4��?8�=?�i#?��>*��J���[��%��ǫ?N,?@b�>���w�ɾ|����2�O�?=�?��`���b�(�D����ͽ2�>A0��~�k篿��B��<�9���Bm��g�?��?ћK�y�6��v羺����q��gC?b��>RZ�>6�>�)�6�h�vg�|�=>o��>�1R?�>�+�?Ntz?ǔ?P_�>�U���ƿpߙ�Jƹ=k4>��T?�F�?;2�?w��?�n�>�\�=�������_��vWT�����<�w�k�>̃��8�>޴�>��?3�3>�
��m��4�<�)�=繜>?(8i>N�?z�>)v�<�Y4?��>���6)����������\?�N�?�W?�]��'���*����-z�>l�?;�?�?:`f���>K���,�!| ��U�>���>��.>�D<{4���A>���>e[�>J�t���Y'9��ķ<��*?�1#?�yQ>�.��%�x�Æ��@H��K�2�6$�C]S��%�<�@ܽT`��I.�	�����������`�P����,����b��#Q���?�}�=���=�]�=5@��F�=���=Eӝ=�Aϼj�|.�<d�&=�''>�w2�F�� �ߴ=�>"'(�.�˾Ȋ}?\-I?X�+?��C?��y>�:>h4�7X�>Q����[?��U>)�O��|����;�����U���}�ؾ�(׾{�c�V🾳Y>L�J���>�3>;&�=�ʈ<���=��t=?��=P7��=��=��=��=7l�= �>/Q>9�u?���ȷ��j�F� %���-?r��>�L�=�ľLc/?w0e>� u�4	���Q�υm?3��? t�?E��>ޓ����>چ���H���Qe��^<K�=�wG=0�1����>c�n>�3�|��=Uc����?hQ�?�%?Az��KLȿ���=-6U> ��:�bS��)��륾ё���~�;�?9��oٖ�
��>���=�k��V�羍�Z=1Q>Nx*>�F(=|N;��{�=��L�F$׼�+/=.�>z�)>�@\=T�^�<T��=�VO>R65>j��=J�R�'cR� ʸ=	">�:>��>�W�>2�?�c0?�d??S�>�xn��Ͼ�-��d��>�	�=Ym�>�G�=�6C>u�>8?��D?,L?�Z�>���=��>��>Nq,�m�m��W������<b��?��?��>(D<�4B�����f>�X�Ľ�P?�_1?Ii?��>�Q����Ya&�v�.�m��?�8D�*=*Fr���T�� �DF�Ĥ����=5S�>e��>�П>zEy>9/:>f�N>/,�>�>wL�<@_�=�f��ʺ�<����Ą=q�����<��ļ/4#�z�+��6���?�;�!�;�_<
�;"[�=���>v�5>l4�>���=������3>,����F���=�s��|�B��x[�{��J�6���g���!>��[>ĝ�G����V?�I:>��4>�I�?ȝz?i>��u��>�����I�����zW�=��3>�4C���$�1R�uqW��?Ѿv��>j(�>F��>��>�: �сP�^�4>�]A���{�?06���=_���V���+k����Ƿj�->`>�3k?�@��Y �>�Ox?�"?���?���>�c��ſ����}=�j%�����I�3�ƾS$���I?��G?��>2c,��*m���̾	����Ƕ>��I�N�O������0�����붾���>,�����о^3��m��Jď�PwB��(r�Gn�>|�O?��?\|a��[��anO�`E��w��N�?ujg?,�>=�?6Z?�䟽����_���H�=In?^q�?O;�?��
>���=�5��Fj�>��?���?DL�?��d?L�S���><n<�*>rǀ��?�=`9>��=�0�=��?�3?�4?+����T���G �`@�ڍ�=��=?��>_�u>Ywt>���=���<���=w3\>�֑>Yz�>�D>�Y�>�ޑ>��nǾ�E?Dxf=s?5n&?��>�����:��b��=`>�^�EZ��y�<��c���&��Uw=њj�V�<>�*�>cm̿��?���<�K���%?:v�OuĽ������>�c�c�5?b��=��>4o�>�6>�}3>-�>fL�{�Ӿ�>�|b!��*C��R���Ѿ�{> ӛ�j�'��T�X���t�J�nѵ�n�;�i�����<��Ŀ<ya�?����T�k���)�:� �w�?�ȩ>E�5?5Ɍ�2��'N>r�>��>���,T������"N�$�?��?1<c>R�>��W?
�?��1�i3�EuZ�.�u��&A��e���`�U፿򜁿ӗ
����(�_?��x?�wA?�L�<I9z>��?k�%��я��)�>�/�';��D<=r*�>�*��1�`��Ӿ�þ4��HF>6�o?H$�?eX?�TV��R��9!>@�:?&�;?��|?]*5?1M#?�3��D"?KW8>tX?J�?�h4?)=?ZV?��d>��+>_�;h��=-O������5�����V����=�=k�+�-��^,=yc5=R!D���:%[�<�����=eO�<V(�=5��=Z��>��[?�X�>�ʃ>z<6?��R8��ū���.?yk=����ɞ�������K����= 6k?4ݫ?��Y?�0c>��@�*�@��@>���>o�#>�#_>��>5*影�B�pq~=�
>3�>!2�=�tV�/��?�吾x
�<�>U��>�J{>[�K�%>�����Q{���d>	�O������Q�9H�c;2�Bw����>��K?3�?$��=���2��r�e��}(?B�;?�}M?Ē?��=O/۾��9��K����mp�>A��<���_�����A:�� N;��r>࿝����v�d>P�
���޾��m��TH�� ���e=�z�~v?=����׾ʣ��u�=�>ؠ��$!�ߢ���W��8I?_a=�줾s�S�SU��} >�A�>�f�>�cQ�-h��y@�`#��l��=�H�>+�:>�@�����I�����Յ>SG?�ob?�4�?R8u���u�t/F��*�����|��?�\�>�<?
�F>f��=��������e��C�p��>���>�����F�>C��;����%�*��>�?�|>f�?zP?*�?A�c?�j%?��?*ƍ>�ͽ�2��xd ?H��?��=�-�P�W��M�~Q���?��G?��D����>ݕ�>���>B�S?<n[?��?� >+���n>֠>� �!����6>�B?ZU�>ec?�߈?O��=�[%�?���w��E�>��>��?�[�>�V�>���>��>;ә���=D�>�'X?�P�?�i?f�=��>i�*>��>?;�=gإ>�W�>J)?�Q?c+u?.hK?�P�>��=<.���M;k�'r�����;��<��=�������&WU��^�=7���.�K)��U;�9;�Qg�;<�<�\�> �s>9�����0>��ľ+9����@>�����F���Њ��{:����=Ct�>��?���>�#�7��=鲼>G.�>���40(?)�?�
?X�;�b�J�ھU�K���>m�A?N��=��l��y��U�u�	h=*�m?R�^?��W������b??�]?e�=�s�þ��b�ŉ��O?��
?��G�1�>��~?T�q?���>X�e�]8n�u��jBb�o�j�ж=q�>1W��d�}?�>��7?�Q�>��b> �=w۾;�w��r��t?8�?~�?$��?U *>��n�3������J���^?!}�>L;����"?H�s�ϾZC���)�� �W��] ���I���r���$��݃�N�ֽ��=��?�s?�Vq?0�_?t� �3�c��-^�����iV��&�����E�Z#E��C���n��_�N%�����ڃG=aCq��WA����?q`?*�\=�>�*m��L���ľɡ�>}ܾP�6�d���o;e�V<�D���UM�����y�
?Q��>s�>o�d?�����/�GeP�D��D�d�X>�AC>"q�>�r�>%�۽ Z��W��D�ѾU^���"��h_v>h|c?��K?�n?Ry��1�Ux��[!�Ľ,����E�B>��
>g]�>�W�����%&��[>��r�����a����	�u*~=�2?�9�>'�>V�?�?��	�����~�x�e~1�zf<G��>V�h?W�>dd�>\�ѽ�� ����>��l?ɚ�>���>����e!��{�Wʽ��>�֭>1��>9�o>�,��
\��d�� u����8�cH�=�h?����`����>m�Q?��:�C<�r�>*tu�ǡ!����=�'��w>�f?XT�=s3<>N|ž^2���{����"#?a�??6~��D6�%>��?'�>���>���?��>�����G�:��>��f?>[?Ru>?M�>I+�=!�5��Rɽ����N�=�U>��C>"k>��R>�n���R��ot�����6�=R'��z�h��9�<�G�<U����W��k�*>z&ۿ-T�٦޾�'�t�Ծ\��_X����漈,�G�U�VD���ܦ��76���J����h�����V���a�S=���?�m�?�`��l��p��:T�i��27�>�i�F�E��=�✽�%Ͼ�2羄W�2�U�0���vP�T�+?��5��Ϊ�|���rl־I�,?�x@?�CX?�Wƾ�4�^w7�,�=��<XY�=�Ƴ��F��t�׿�D��ͼj?���>��3���>�s�=}�=ร>5��1xF�i|<���>T9?B�?q���Wֿ:�ÿQ��F��? �@AL6?���^/��#�A=��>�}?r�>�_ӽ[,���ξU�?}�?6m�?.Nѽ,sM�v�>��g?��>?J��=f�=��8=A��=%���->O4�>d*(��p;�����@>��>��J<F����*E&>J�>>��B��7J��Ԅ?z\��f���/��T���Y>�T?�*�>�5�=�,?(7H�}Ͽ�\�~)a?z0�?���?��(?�ۿ�	֚>��ܾ*�M?�D6?���>�d&���t����=-�����@���%V�B��=ܪ�>��>�,����(�O��`��s��=�*��8ƿ��#�w���-�=ުƼ�c��%�b���D���S��oؖ��c��U�<��=P	>`F�>R�L>`Sf>�xQ?�sd?I_�>��=k�?b��۾�og=��h�12�Z�ء�݃��c(��?߰�H��L�l- ��7ľ��A���#<�=Q�_���_P�3�O�PbK�#k)?;�f>P�ԾZ<��琼u�Ծ����W�<����?�ξ����Z��T�?E�@?߈���9E�����=�佥 K?&%ʽ����}����=?���]>�b@�>l�=�'پ���H��=)?z�?�J�����B#�=A#�����?+��>�1=խ�>-�?���j
��x=!fy>�>��?���=홾Ɍ��{/?�0?*���>����>�wy��Y��R0��!>�^�w��s��>4�>{���A���ȅ���,*=ZW?� �>��)����th����� 28=��x?�r?>��>�Bk?�B?�4�<����YS�^�
�*�y=$�W?"�h?�a>�ぽ>�ϾXP����5?��e?? O>{kh�����.�����?�n?��?�[���|��
��M���5?�o?��X�b��O����V|��H�>Zy�>��>,�2����>�AH?�D�����*����1���?��@5��?���]��V�=���>-��>�~T��2ƾ���6�����/=���>2����e����e9���4?�A�?C�>�蒾4��\��=�=�'��?��?�6нl<7�:�"�X��?����>F\彨�X>}Kʼ�۾r� �*T�����ƭ����<Leh>�;@���?'?�h��zNͿ�lڿZ_���눾Am*?K�>���>ʀ���^�E�A��4�_�b�r��7��>�&%>lY��6�P>\��H�G�"ԃ�-�a>��%>�T#?�ڽ}1������U;>�/�>M�R>��>�*ƽ���<-�?#�8�	��r*m�b��~��?K�?��?��%?��/����^P[����ҺF?�T`?��?�J�=�M0���Ľ��i?�,��R�U��0��D�J>�<?�$�>�%&��%=���='!�>Le>J-���ÿ�����;�s/�?�Z�?+���>�?^�*?7��� ��Į�qu.��/��'�A?�B(>)Y��Qj���@�눙��n?��/?���/ �۲_?VVa���p���-�]�ƽ�I�>��/�?	\�n���  �#:e������[y���?�U�?���?���H#�w-%?�ԯ>���KǾ6��<�$�>��>��N>9�b�g�u>�����:���	>Š�?Z�?~?y���P���Fr>�5~?x$�>��?�n�=�a�>8c�=$�g-��k#>� �=8�>��?l�M?�K�>�U�=}�8�g/��ZF��GR�2$� �C��>_�a?��L?�Kb>|��D!2��!�wͽqc1�9G�mW@���,���߽�'5>��=>>��D�XӾ��?�g�ԂؿV��5�'�B4?P�>�?%��u�v��_?S/�>�U�f��� ����i��?��?�	?�g׾̼�d>A`�>�2�>|�ӽLޞ�}����q7>S�B?�����T�o�g��>��?�@ڳ�?� i��l�>�: ��܄��6g����[s���<^g;?,mþ��=�t	?��q=��U�9����`���>�!�?7��?п>��i?ܗH�{}0�^G�=&�,>�uE?u�?��+=������=\;!?��;s�C�O��b5?��@�-@BZ9?Ȭ��ÿS$���]˾V���Z[>�R<j3�=�4� �<�Db��$������G>��>���=�/>�,u>�=�$�>n�~��$�}в�'�l��F�������}����m�ƾG�3�ȋ�s��Ƀ��]���87���t�%
�������=?�U?�R?�p?� ?��x�R�>*���*;=`�#�̈́=�.�>�g2?�L?��*?�ד=j���8�d��`���A���ȇ���>�qI>��>5J�>#%�>�`M9��I>�1?>���>�� >Tg'=	���^=��N>�M�>q��>�|�>'�>>�>��������L�g�Q*q�+�Ž�?���}K������\��X������=>/?҄>������ϿS��8G?�n������)�:�	>�j2? xX?�:>����Gh�7>�E	�O�k��;�=�����f��+�&B>JQ?G�m>�ޜ>v�բ{��XZ��?ӽ�[�>&;?�F������3]�"�����78>R%?w7�="����ȝ���N`�?H�=TZ*?���>�l��h���wؾ%X�=���>�H�>�Ya��q��R>a>�罽�n���>ta�=E��>��>��}>�Q�=���=҆ľ���=ZcM=�J>^L��xs?��K?=ݩ>�~P>�S�F���
?��;?,�?�C>�!��a�=D�>��`<�O=Ċ�����9�(���R>�8M�BV��:tG��1�=j�>=���<�
>HW<ZQݼ�J��~?���䈿��0e���lD?i+?P �=)�F<��"�> ���H��5�?l�@m�?��	���V��?�@�?����=
}�>
׫>�ξM�L��?��ŽǢ�Ɣ	�g)#�fS�?��?0�/�eʋ�Ql�6>_%?|�Ӿd�>�|�Z�������u�x�#=��>
8H?_O���O�v>��t
?r?�c򾼧����ȿ�yv�?��>��?���?
�m��?���@�x�>x��?gY?zvi>\j۾�`Z�L��>@�@?�	R?��>�;�3�'��?1ݶ?Ǭ�?�4?>�?b�?x�>�]l:�(=�~˷��w��,����=��>H�^>a��� 7��ȑ��E��-b��!���g>5T�<��>{��%W��Z`�=��Ž����.��I��>�">�@�>c�>�?���>7�k>{jL=����v��wԏ��K?��?����=n��ܼ<h��=2r^�]4?@j4?��W�+�Ͼ�`�>�}\?X��?@[?|��>���� ���޿��Z�����<٠K>A@�>77�>e���)eK>��Ծd�C�\�>M��>򂞼^ھ+��7ɥ�b�>�Y!?���>���=)v ?��#?l>��>�QD�h���LF�43�>��>V�?��~?�?c>���2�Yْ������[��N>�y?K�?�ޓ>���:��
�,���H�����0ǂ?��g?��۽q�?r�?��>?=yA?m�e>��^�׾<����k�>�m?��= -��A�`����K?�?��?"@�ѫ߾U��=�@龄����>�
�?��0?����J�3W���gZ=@4>��y�O��=<3�>�:�>HL���Ƚ�1>����WG|�S�G�0�F=�]J=;�?=7�M�x���Q�>>=,?b�G��ڃ��=��r��wD�'�>cKL> ���^?�i=���{����}x���
U�� �?���?k�?]���h�$=?[�?1	?�"�>�I��[޾O���Tw� x�cu�%�>*��>��l�,�͏������E����ŽԴ��7�>̄�>]�?0��>�BQ>���>�
����(�i��� ��\�+[�`�8���-����&��y4�Ӭ�$h���nz���>�����˱>*�? �c>��r>x��>Vn���D�>tdS>XW�>Iާ>]�Q>�6>sn	>�W�<C̽�HR?ޫ��L�'�������&B?}]d?�T�>+�f������cc?�n�?3s�?��v>;mh��*+��^?�#�>K��aZ
?�:=����E�<p���%0��s���w��Q�>ƨ׽y:�%M���f�xW
?�.?�j��?�̾6�׽����Ko=|N�?��(?��)���Q�[�o���W��S��K�"$h�+a���$�0�p�+돿�]��l"��W�(�o�*=��*?K�?l��������#k��?�:zf>��>K8�>�ھ>�oI>!�	�Ի1�� ^��I'�����VW�>\[{?�Ӎ>H�I?'�;?��O?D�K?��>��>�P��F��>�*�;��>��>9?�.?	�0?�?8+?*rc>`���u��1�ؾ7�?(7?*?��?�?gi��1�Ž���������y��䅽��x=�w�<'�ֽ?��(�I=<�Q>0?"�7��7����d>�V7?��>�>�>*s��K��
X=_��>�i
??�>  ��o�~		���>�?��
��B=+>;��=,���V��:�%�=��ͼ�g�=[���w.���<$�=��=��#w�;m)�;�Ѭ;��<���>��?�ĉ>��>�1���z ������=��S>�cS>�>�6׾���C����^g��+y>�:�?�?�.f=��=�?�=a{���ž�+��eL��,�<��?xB!?I�R?x~�?8<?*"?#,>C�����Tτ������W?$/?$�>a�;�7���j���*��jJ?�x�>��+�5����H��oN����>�m4��ˈ�j�ƿ�%H�g�u>]�_�Y�P7�?�͋?����U��<���i��i��5o<?&�V>(�>B�>�C���z�I��*S�=I?� A?�x�>ٟj??�?��g?��>M*a�m�������R���n>y./?�č?�A�?�׆?��c>�x&=OE:�'��Vx̾B.p�~�����\�����6s>��[>7=�>���>		>�hi���=UW���H>ag�>���>*��>AW�>,>Z`J���9?��>�L���(��7þ�4������?�̗?��,?!eѽ�F5�s�2���ӾT��>��?4��?�h?jfS�bY#>k�ҽ7׾F�=�R�>�>�p>�½�p�c.M=�?�9?�� �>���5�xI����<?�>?[�|>��ҿ��������S�=�QT�<{��Rj��ʽ����ؾϕ�H�Ҿ�Ei�i��T���������~������0�>GJ�=�8�=���	���x�!=
E>д=|!b�K">�>�x/��N~�wY¼O�U=�)��Qq=5��=�R��!˾�j}?�
I?D�+?̓C?��y>�e>�<2����>!�Z?��U>�`Q��˼���;���������O,ؾ, ׾��c�ˬ���5>�aL��>�3>L��=�}�< ��=!s=�ӑ=ߪB�I2=d��=]�=㏬=@�=O�>I>/6w?��������2Q�e�A�:?�6�>@��=ˀƾ�@?��>>�1�����c��-?_��?5T�?"�?�zi��d�>���厽ht�=����u=2>i��= �2�`��>1�J>���J������Q4�?��@/�??�ዿP�Ͽ�^/>�ǁ>,�=L�N�V���C�þ5r*���k��#?Ч%���ྐྵn�>��+>�S/�S�q9�=`��>�p>��&=rde�j�= �0���=��
=�I>6�W>��p=����t?=���=:�p=�">"�k(!=4;>,�=h<���=~�T=f��>��-?��F?PȄ?��?�^þ������K�>s�+>��>�a >�b�>��>�w$?��"?&C?Bؒ>��0>�;�>%	�=�d��O��홾#l�����)�?�W�?Lw?�Ѝ<n�M���GW.�z���?�_#?zL ?G��>s �]f濱�>���LOq=5���=$>+1���Ǽ�/��)���𗞾�˒=��>]�=_�$=��>�х=�Ì>��>�	D>&�(>��o�,7>�b<������e����y�fR�&�ý�8
=�*�i�.��U>j�=u�>��9��E�=���>�;>ʗ�>)�=]����/>m��$�L�`�=�1��h$B�z4d�}7~���.�a76�t�B>8(X>f`���"��{�?��Y>/}?>Qw�?CSu?�>L���־�K����d��S�q��=�<>�!=��b;�O`���M�eTҾm�>nW�>�#�>�4~>6���^��ό>��_�(ؗ>��𾚗k=�d����j��s��T����d��xý�kX?`���ȃ>!�z?�B?bn�?��>�N������W��eI��k�>u;/�OTs��.Q�!�?��>�1?\R��V��E̾J��n�>��R���M�n��Lg4�o)<����>�Ɯ�ξ0�5��z��wȈ���D�.�r���>��G?��?�B�Yx�4Z@��f�-�&��l?[�e?h��>];�>Xk?
�����Ҿ��{���/=:rl?��?���?�Ǿ=˶@>�KнG(�>�8-?P��?1�?��c?gv6��?]%;=W>�=	*���<�~^>�B�=�1#=0S?� ?�C?�U�r� ��U�۾�@j���	>��!>�c�>Z+�>���=��g=`�|=����H2a>E�>���>�v>���>�~>�]������O?���=�%?v�>)_�>�I$�-����M>jW仲��nk��]6!�ceW��\�2L�=za0;dkF>���>cϿˢ�?�[��_���H�>!����⽉��>���>WL�A�?�1=���>Qk�>B(->�Ȱ=:8�>KN>.�Ҿ4>���8!���B��vQ�;�о��y>:���cg(��i��P���I�派Ҷ�j��]����<�z�<-/�?�����k�TE)����&?�w�>i5?���������\>�A�>K�>\���/���QՍ����'J�?���?m<c>[�>3�W?��?R�1��3�vZ�ƪu��%A�=e�<�`�������c�
����[�_?��x?�zA?N�<�:z>N��?��%��Ϗ�j'�>1/��%;�S<=�'�>-)����`�حӾ��þ�/��GF>��o?U$�?(X?�RV�z�m��'>��:?��1?�Ot?��1?7�;?L����$?ro3>�F?�q?!N5?t�.?�
?e2>�=p�����'=#7�����ѽMʽ�����3=o_{=qZθ��
<v�=&��<w��ټG�;�&���'�<[:=��=�=J�>X?['�>�Yf>=�"?��	��;�����˸?^��==R6�<�L�v�����o(=��h?mũ?6�^?4!Q>��6��T)���	>�k}>w&8>��>��>���8%��&,=�>-�=99=P�<�F��������=��=Q,�>7��>�N��3>"���F���V>�/�����+�O�&�>���3��ё�ἳ>��I?�? 9�=)�ؾ�}����Q���?�')?�O?�x?�E.>¾���@��b�I�j��S�>��=�
�^���򛿾�+���V�W?>`����}�I�
>@�c�ɾ�E����&��>ž��=��	�*�<���<���j�t�BR��9�I>�}�����~슿�԰��:@?�=
=U����	���e����G>���>��>����f0߽~5=��E���陻�?�m>�9�����;�%����r>KW?J�o?�N�?���O���K[������u��=��?���>rL?p>^�<lך� ���m���=�깻>�>,�,9�}�F��Z���=���>���>��{=��B?<?Ai?��g? �?`]?hr>�S���5���#?%�?�^�=ڠ�*Cj�:�7�Qd?��L?YQ?�-F��o>��>r�?��)?�l\?A��>�>���;�H��>���>v�E�܁��yUb>��I?t�>
�k?�w?���=e�0�Y�þ����1@H>��D>�?o?� ?`Ӧ>�a?fT��=��`�o>��!?e��?J?j�=$(�>e9�>��+?� �>A)>��y>d�(>T_?�X�?|��?_�?R}\�]�}�qN���m��
�<i�=��z����=l��?�����ж��6��h<�����20�)�7�r��<|2=���>p_p>Յ��~J>�WǾ�Y����D>O�������ȁ���H�Pܪ={�v>���>��>�g ��ܘ=�[�>���>�2� �&?r?��?
�J���d��?վ]wM����>�D?��=
Ol��)��D�u�p�[=�fl?Ƽ\?=�T�z*�/�b?�^?�I�=�^�þA�b�Rl�P�O?!�
?��G��ɳ>.�~?9�q?n��>G�e��8n�����5b���j��ɶ=3j�>oS��d�J�>'�7?���>Tc>���=[�۾��w�R���?T�?B�?��?�*>��n�)࿝n���A��� ^?""�>2�����"?b|����Ͼe-�������5-���~��s����%�%������ֽ�#�=��?S�r?T_q?��_?P� �v�c���]���=�V�/��:�tNE��D���C��Pn��I�����@��l�C=&h�T:-����?V�Z?Y�D>&��>�>��U�h�g��=X�U�d�>On=�� ���=-��2����\�����B�)?��$>L}N>�`?�J��+�
a ��H��	�O �>UE>���>��>*�<7�0�wb�����}d���B�{-l>��f?��P?�w?P�Ƚ��4�����<%�Yr������e>�R>G�>��U��S��.$��/9��r���m��׋�$TH=��1?V5�>䟦>q��?�?q�ʰ������2�B�,�.�>�f?���>熐>�H�������>V�l?���>�O�>c���[!���{�s�ʽ��>��>���>%p>Ǖ,�x\�Dg�������9�0��=��h?�k���a����>�R?$�:ƶF<�j�>U�v���!�ݳ�9�'��>�{?�ª=P�;>�~ž]�C�{�%���M#?��,?�`6�y'�Q�.>d4?���>�?(��?_$b=���g���@�?_M�?�ff?�`?�i�>j�p���K����$S����*b:>+�>��B>W�>�T���"��iD�����=��5>=�#�=k�;���>f�ؽ��-�we>��׿,c����оꂼ��;�-���(x����P�����!ӾW,��X�~��m;}G��y_!�������ӽ�1@��?l�%��X��V�����������P?�p��ս[=r����]�,����bl��2c��u$��R��Nw��'?�0���&ǿ҅��d�ھ"�?�x ?;�y?B\�Zt#�89�G�>��<�w��f�E����ο۬����^?oW�>�������g��><�>V�V>�tp>?���������<�}?��-?��>��r�éɿ�h���М<�[�?Y�@%�7?�6(��X��8�=ŭ�>p�?{�C>f	�� !��D���!�>��?��?����H�G=��a?C�<q5>��Ir=Y?�=\&�=4��=�(F�fw->�c�>�&׽/�l,5���=�Ս>��O=�#��&o�=<@>�
+�}yb����?c�[���e�0�/��@��!&>7{T?�V�>_%�=8,?H��cϿ[\�U�`?�
�?p_�?{�(?;W���P�>c�ܾ��M?�6?�~�>7&�'yt��=�=��˼��p���PV����=�,�>>�u)����j(Q�X����+�=�p9˿���%���(=N���2��_��Wٽ�ƽ�2���,����$�����Ý=n�B>ԌX>�C@>�̝>p�S?�cU?^:�>��4> �ٽsی�My־��	���[����^���5�9q���۾[�ܾl����3�5,��nK/�>G�;�Y��f���2*��pG��	>�%�+?�
>�����<�eS��at�]+Ծ��;��
�����~�BB_��Ԡ?�;?��|��O���i<�(@<'�K?4��=�� o���7>�U=x{�:R�>��>��ɾ��6��M�%�-?�I?0���EW���b�=�ˑ����=;r?m�?B�=��e>�&?=�,���ؽ4/4>�~)>��>YN�>t}�=����왽��(?ܴE?�P�-l��=f�>Z`��]�5���>[ǭ=��d�xuY=�N>#$;�BJ��ږ;kQ��Lf=X�U?z�>�)�`j�|���.��f�S=Ϗr?�?V�>�&n?�DD?�)�<�<���`S�����2c�=(s[?N�h?��>����Ծ㈠��l6?*�d?7�I>�m����d�,�v�����?�d?H?;	��C{��摿�m��$8?"�v?�P^�i�����ѯX�r��>$�>���>p�9�[ʳ>�j>?��!�����ÿ��?4���?5q@�?�?7=<̧���=�!?�p�>��P�|ƾzC���
����n=���>�n��	�u���i�-�.38?ֻ�?�f�>B]����!��= 6�(��?�d�?cA��˽]x�C�����+���=qrp��u�>Գ�<4Fƾ_�����D��[�ؾ�!���?>��@����n$?����}�ٿKm�Ϳ��5|�J��=ʥ1?�Ê>�W�=��e�ni��,���p��[�0þ���>���<VK�
j|�T������������>��7�6�>k�I��6��}������8�>`��>�{>C�B�(:�?I��m=¿2R��IX���^?� �?ٴr?�?l1<89����Z��'��pY?H�f?�7?��ν&�@������j?c��o-`��4�A2E���T>�63?�4�>Fa-���{=�->���>OB>��.�ЊĿ���B����ۦ?�}�?�x�~��>'��?�x+?����2��'����*�Y�F��AA?Ml1>����y!��'=�����
?\c0?���7)�?�_?�a�D�p���-�<�ǽG�>�1�m%[�CEܼ���Ce�y���y�׭?,J�?�Ѳ?I��"�x�$?�{�>̔�:�ƾt��<I\�>��>6�M>�RV�)�v>5�*;�F*>Um�?_s�?��?i�����
X>ʣ}?{@�>��?��=��>oz�=�۰�W�"��#>c��=��?��`?­M?9��>���=�Q9��/�0gF��CR�����C�� �>Y�a?6zL?y�a>H���"0�"!��Fͽ#�0�@��?r@�C�)���߽�}4>E�>>8>��D���Ҿ��??s�w�ؿ�d��v�'��74?���>��?����t�ob��4_?4^�>�C��$��4$��y-����?=�?��?ݧ׾��˼�>�ȭ>�E�>iԽ����7�����7>O�B?����2����o�f��>�?G�@]Į?�i�63?���J����q|����6�,����=��6?5���K~>=\�>]Ա=JFu��k��Y&r���>O;�?��?X]�>R�l?�Ll�)@�C�C=���>��h?�O?|��`�5>h�?r?�4���<��Pc?��
@O�@DX?f�-7俹����ް��=��s��=�F=�M>0K�M9k�C+!���>��$9�_�=}~>Q�P>3fm>�}>9&u>Y>Ԃ�����"��ZB����>��-���
�G����0�"����3̾��ƾ=ؽBߏ�_����m���� ȑ���=�V?��R?��p?�?�π��^>n��O�=�q#�\�=u-�>2?b"L?7~*?v��=Y�����d��)������������>b�I>��>E�>��>I�;��J>+>>��~>U:�=M�=rӘ���=��N>"��>Fe�>W�>6[>�x�=Dӵ��!��>�l��L��5�;�?����KK�L����΀�m=վ���=J3?(�>�S���ƿ^k���94?O�����l��e>��?/WR?R8>o���Y���U>����B����w>�F�^�=�7����=XF"?��>��>7M=�;��A5�{Xٽ�˥>�`I?o.��&ĝ�?Ij�ت?������>��>�����{F��a����i�C��X��=@q/?�=�> �ѽM�þ��3���c�蓅>��Y>���� �<�އ>��4����3���=���=�FV>PH?,��=`׽�S=-�ľT�'=V`W>�;u=j�>�Q?�S?�==�K�~�Ǿc��E��>�1?��?v8K=�Lu�zz1> ?Z����\S��c����9��ڹ=��>��׽t8t�0�H�Ms>Y"n����>{G>5z���뱾�,��s�~?�w��E߈���NN��gD?0?;�=��G<�"�� ���9����?\�@f�?�}	��V���?�?�?������=���>Gի>�!ξn�L��?�'ƽ����<�	�<E#��N�?��?�/�`ˋ��l��.>�[%?>�Ӿ]o�> ��u��N����v�n�0="2�>��G? ����?��}<���	?�?����壿��ȿ�=u�y��>�-�?��?!�l�����/@�5��>�"�?OUZ?��f>� ܾ4�Y�6Ջ>�,A?|�R?^�>�Q��
"��?���?��?f�H>
��?��s? |�>k�n���/��i���ǌ��Ip=��;8��>v>�#����E�~���0����j����a>�!='(�>T�佩컾�ո=�������^���>��m>�N>��>�� ?���>���>̿=6V������'W����H?�l�?2��y�i�zҏ<Yt�=V6��?��=?ऍ�h ˾g>�Y?/f�?��b?� �>���j���/���Ũ�^��;�*><;�>3{�>J�/ي>*�ξHt���I>˻�>���<��Ǿ��U��v�	6�>��?Υ�>�V�=�g ?`B#?�8k>G��>�$D��A��CF�Ð�>mH�>(?��~?|?N츾3��Ⓙ�㡿N�Z���N>�Py?l|?6A�>g��������X<���J�ܔ�M�?�(g?���?u)�?�o??�A?g"e>{��,׾�z���a�>��?�&$�O�T�N���f��f)?�p?��<?�d��׾�6;����3w�o�7?�@~?���>a�?���t�����5����<��,=i�� k>�"�=�+�=_���)Jt=���=�+�~�	�v�#� UD=ς1���>��8��0���>�`*?
w�<Z>s�u� =(m�L�B�|fg>D�Y>�+x� T?�Q5���u��ۡ��Ó��8'��0�?P��?4]�?���d�e�lI?8�?_�?��>su��C;ھ�Q��X�½�H��$���
�<��>j=˓��.��X �����~H��JZI��:?��>��?Ɏ$?��>��?�������9�ϡ�A�z�<
龍M
�؅Y��*��$��<R����)�51�����a��>��x�O��>�k;?ƈx>ϸ�>���>��>#�>u�=7H�<�(x>^��>W��>��>۫ =�R}�$R?�ѻ���%�V龻$����@?��d?Z�>�B����@���D?�ϒ?}��?�o>]�e��+���?&|�>�����l	?��Y=�-��)��;�����q�>���E���>n=佫�9�ܱH�2�c�-A?�_?ܛ�X�˾��׽����w��=fs�?�v,?U%��R��Fo�XrW���Q��.�%_�����P#���o��펿L�L��8�&��G=}�*? ˅?au��辱>���'j��K<�}d> ��>���>^C�>�gV>�K��$/���^��~'�[с����>��|?�]�>h�I?X<?��P?i�L?�a�>\��>)���m�>:��;:.�>`��>C�9?6�-?Y30?1S?�X+?��b>��������ؾ�?�?�V?�
?��?]�����Ľq��r�r���x�Y�����=2�<��׽��u�X=;�T>�"?����k���վ�K:>�'?C"�>-�>׾��-g���J<
��>�љ>V{�>��#��=� Xܾ1|�>?KS=� �<j�F>�U>!��n���>`O(��ĩ=�u�=�D�Da9=�/�>Eu�<�<&�t�e��\=<��OK�^}�>��?i�>��>)G���{ ������=!Y>��S>'*>پpu������g��dy>}u�??x�?��f=R��=�o�=�U���[��������Q�<ڏ?><#?HT?���?\�=?�e#?��>��7��~K������?,?0q�>�S��5���v���l/�\:?%��>�e �� �~h����I�>�ԥ>�aW���+������H�C��=��'��~��B�?� �?p&5�w(a��ʾHi����Ծa�4?9I�>���=*�?]�.��`\�-T��->�(�>tO?Ef>=��?=��?�\�?�>�>h��y1пp褿�����=�y�?��w?A�?� b? �> w�=J᡾�����ܾ��]�>�W�i�udl>��)>���>��>�P�>2�>㕾��~�+�6��=�zl���?�Q>�G(?Y'�>O. =r-?O�>m���D /�������+>UTO?��?��i?�\�=�{ʾ�Ҿ~��.�>C��?>�?J ?Rէ��Ú=�ٽww��U�����>���>L�>x�����S�>���>�#�>�n��}�
��H��=v�?0?A�>�ݿ�瑿��b�>�Y���{=E�����0l��	�����<6v�K�C��.���a��$l}���־�ߧ�$����=�!?�t�=���M�>
x;���;�8�m�!=��Ƚ�i�<��2�H! =V5�=�a�=�uh=&����=��>콼}�˾��}?_;I?��+?F�C?#�y>;>P�3�3��>�����@?�V>ޟP�:����;�竨����D�ؾ�w׾��c��ɟ��H>$fI���> 83>ZG�=rH�<�=s=V��=q�Q�`=^$�=$P�=,h�=���=�>:T>/5w?ᚁ�ɲ��\1Q�É�J�:?�9�>[��=�ƾ�@?��>>�/��ʔ��f�p-?��?�R�?�?�i��d�>(��>ꎽ�_�=���<E2>q��=i�2���>��J>���I����5�?5�@S�??�ዿ��Ͽ�G/>��@>H+�=�^Y�d(��E���>%�M�;��2 ?!f;�YN��3@{>l��=��پDR�V=S�@>�S�=U��ۛ[��=�6k�I:_=�]=�GY>��C>>͍��`�=��	;��=NSV>��=����3��0��=��=��+>� �=���>{�?/�8?ѩv?��>�}��7\޾szȾ��>bQe=e
�>vs=�A>���>�94?6k7?ksF?ր�>�k�=*��>iF]>@�<�4*`�z����r���3�=KɆ?�Uy?�o�>�+�f������H3��"�a�?�%?I�?ˉ�>$��{��0��#M7�	U��0������}�rఽRR���w"����td=1fW>�ê>\��>��M>L�>ϭ�>z*�>A��=��=�l�<�מ��A��+�#��=�=a���rb��W<a˒�{����Bý���*J���`\�0^<"z�=�[�>p�>�%�>���=Q_��/3>u�&L�ZЬ=�*��[B��`�'�{�JS0���A���=>]Q>�놽�Ӓ�?��X>�8=>�\�?��v?��!>����LԾ�n��L[��[�#��=e	>�=�a�;��G]�:�L��9Ҿ�m�>%a�>���>�Yz>�j�KDf�5_>>\���-����>�׾�Fν�M!>�9�b���{�����e��t� �%?񭙿�&>ݞZ?�5?��?X �>�ѽ�ؾc=�ݾ�v�>�X#��8꾵�6��[�>�.�>�?Iξ�_@�ZϾOH�ĭ�>��1�K�����u5�^R=�R��l�>�,��;IݾC�B������K��]����>2�B?��?J�B�a����<T���&�J�;��?J�^?�ӊ>��?n?z�ҟ����80�=\`?�@�?��?���=dM�=*����U�>��?��?O�?�}p?0yF��X�>ުN<��$>4���7�=[>]k=��=�t?��
?oz	?�ס��
�����J��#ZX�w>�<F�=ˁ�>�*�>�v>z�=P��=���=_m^>�>{��>�b>�J�>�>�����̾�AB??�S>�?�o?Lj�>h��f,�{��;w�0����t�8�ަּ�e����Q����4x|��>$��>�ؿ=�?h�=���:��>��|�+��G>@#�>0蓽AM?o2�<�ȃ>��?u>py>	µ>i��>3~Ҿ��+>����E���+��[R��^׾�'\>e����,@���-LӽN?�DW��Eh����e�3	z�qm2��\X=���?�R�9;z��N��߯��D?���>��0?3��p�2��S�=?��>�j����ˋ�}�׾2)�?�<�?�<c>'�>��W?
�?�1�f3�>tZ���u��!A�/e�$�`�{���`���)�
�9���7�_?V�x?9xA? .�<�0z>���?��%��ӏ��'�>/��#;�Ё<=2�>�*��Q�`�Q�ӾA�þ�0��VF>�o?T"�?�W?�JV��m�2 '>o�:?��1?�Nt?��1?ڌ;?���_�$?^p3>�E?r?�M5?��.?��
?�2>j�=���c�'=87����ѽe�ʽ��1�3=�Z{=�׸<��=��<��ټL;D!��_)�<�:=.�=i�=$�>�d\?	�>�B�>y$4?�)�[6��⩾�"2?�UV=��~�5݌��N����Z>��h?!�?�Z?�8c>H$B���;�S�>��>2)>�`>�Ȱ>�սV�C�7�t=�$>��>fס=zO��}���	�N����ð</n>��>'�>�H���>�����ֈ���{>.CT��W���S��IN�A�.�I)>�t�>�??�}?cH=����w��+*j�A�%?�F<?D�I?�?#.!=��㾉V?�KTK�Ә(��u�>_~<��
�I͢�������C�,��<��{>����x��i�Q>Q��"ܾ�@p���K�s~;���=ve�v�)�����޾�o���->~�;>?Ŷ�Ȥ$�dc��e۩�UlH?��=+z��Ař�� ����>qA�>���>����M����=�P3���F�=�6�>8�*>u�ܼ?5侳�N��
���>}E?@t_?�m�?Zr����r��lC�ƌ��)����]���:?�0�>�<?��@>f2�=�汾�	��d���F�~��>�m�>�$�M�G��W�����Zs$��ފ> b?�>�?��R?h�
?�v`?{l*?�?��>�a������F&?�~�?Ү�=��Խ��T���8�DF����>r)?�B�ࠗ>�?��?=�&?�qQ?�?�[>� ��9@�׉�>9u�>�W��a��ή_>��J?0��>	=Y?��??]=>5�=Ϣ��l���W�=b�>�2?�#?(�?S��>U9�>�Y�����=E��>v�c?C/�?}�n?U��=�.?��4>��>�Ȝ=V�>	��>64?%O?��s?=�J?��>yH�<�c��&����l��x��1�;0�L<Y�=���ej�p���<��<�ɡ�ghF��Xۼ�F�`X���<�W�>[�t>�Օ�D�0>O�þÈ�tA>d���ۦ��0
��`X;�3�=�w�>�j?���>!h'�T�=�3�>b��>����]'?�P?�E?]�;�b���ݾ�hP�(��>�uB?LE�=�k�� ���u��ih=�m?UP]?JV�2���4�b?w�]?�U�r�<���þR�b�b���O?�
?֏G����>l�~?��q?k�>s`e���m�d	��.b��j��=#��>�o��e��͝> p7?�c�>��b>���=~w۾3�w��;���5?���?�ݯ?��?��)>��n��!࿏��`>��6�b?1�>q��$5?ɹ�2M־3�I�:k|���Ӿ��p���KN��jâ�r��&u�4��|�>-?n�y?_c?-�Y?�.���dc��`O�w��x�O�������6_F�m�C���I�7\u��>�;�������b�=�1B�U�\��ñ?B�.?�4��?�䬾n�!���U>݁��&��"�=�?,��r=T��=�T��R��*���? ߺ>���>��1?0K���0��}�b?��3Ծ�>�,[>2�1>��>4�_<��d��W+�
�־���U���3��>�Gf?r|O?gsp?g���P'�����M*��"��u5��4�v>�pA>�Ĉ>Gs�M"�&3 ���7�&i��G�C&���:����<_%+?.��>J̲>2�?�L?X��f����0���~1�R�V<�-�>C m?PF�>2��>�M��*����>��l?���>��>���Y!���{���ʽN$�>�>��>W�o>ߪ,��#\��j��,��� 9��w�={�h?炄�]�`��܅>�R?�:Z�G<nz�>+�v�W�!����I�'�<�>�|?��=��;>�xž�!�j�{�.;��R`)?i�	?�N��L/'�av>�p?�t�>���>��?*��>����gH
���?8f`?s�I?>�@?�i�>h=�w��*VýH���r	=D�}>�O>�ye=$�=\U�G�a��r#��+=H�=���M���j�;U?��PT<m&�<I�+>�6�O�wӾ��
���8z�Y���e�1��E�����¾�����]����f�&=�/T�c�`��if�`���?��?I�׾�񵾢|���������=?����9��	����ྖ������kkf���T�e�s�씃�22���(?%��Ŀ�'��?X�A?�&!?�u?��M�#�6�:�3�>)J=*�0��,��ޙ�0ο�����\?�T�>��辸ȶ��Y�>��>kf`> o�>XJ������|s�<C��>k_%?.� ?NQv��-ɿ���n
=��?0?@��??j�8���ξ�Z�=h��>L�?�|>HZ>�l���՛����>�y�?怊?�Ö=�=M���ѻ��\?W�f=T�9�]Pi9��=��=[�<L����[>��>���!��t�,� >c�M>>"�-��t������T>)]߽3���0Մ?/{\�jf�N�/��T���T>��T?�*�>�;�=|�,?>7H�>}Ͽ��\�+a?�0�?ߦ�?��(??ۿ��ؚ>Y�ܾ��M?D6?+��>�d&���t����=�5���������&V����=���>�>�,����ևO��P�����=���nʿX� ����dk{<��(��+ͽ�����ӽ�֡�	쉾��Y�������}=S>�ω>��>A.c>V#|>2�Y?S>m?�h�>�CD>�q��`���f��&Қ=��5������OY�l꡾?�߾�;˾s8�t�����y�<�S�a��=�%R�F����:�JFv���*�F	0?Jw>���I�T�߸�E�Җ��T=�=��&���<<�EӁ�Ŧ�?�F?.���p�r������rC���<��c?�n��>x��ľ���=�����*=��>U(�<u�پ�WS��ix��O?��?|G���A��Y����1���=�1/?G3?��]��j�>�{?���I.���>���>��>9#�>��=�]Y�8<�����>Fw?a���;���=;'���	�I��P�L>t����m�>~�+>♄��+��r3�=�=n�S?ѹU>[C�R�������_�kR=�Kk?Ay	?���>�Rb?.�>?������+B�����
=zQ?�&^?#�>���,��|ȁ��Z4?�Y?^:>n�����Ӿ���70�>�5�?-T7?䣽�Ws������a�q�3?��v?wr^�Ls�����!�V��<�>h\�>A��>k�9��j�>�>?N#��G�����9Y4�6Þ?x�@)��?��;<J�r��=�;?/\�>;�O��>ƾ�z��������q=�!�>O���ev�~���S,���8?Π�?e��>��������P>PŦ�8�?��?q.-�?B�>�->�Yǃ��nY�)@>��w>�GK<)���M�:`� � �����0K=n�x>�/^>)7@	G��ae�>�LX��'�kϿk��E�5�7�Z��+?�?z\���g�k�s�ג��9�N�чo��(ľĉ�>�.>�k�������z�T�:�&���"�>�ڼ�>L�R�\a��E��L��<�|�>�>���>���.���/�?V*��a�Ϳ���/���uW?2��?���?�?�Fz<��z�\G~��TM;LrI?!%r?+�X?�p7�NAd��p<�J�j?s茶p_��|3�%�C�ST>�3?�A�>�,��~=��>�d�>��>��,�ſ������?#��?T�ׇ�>4�?B�+?�������~�����+� w�:jB??x<>JT��=� ���<�GI��-�
?y/?�F�O���/^?�(f��g�����,ӽ���>1u0���^� "�<���[�d<���i�Ԫ?��?Dҭ?%�<�Z���S"?���> ����fݾ��<���>"�>�N>-�̽p�{>L����=�u��=ލ�?���?��?g�������3��=_�o?�2�>��?3p�=f[�>؊�=i氾��,�7T#>2�=�x>�ߘ?��M?``�>ϑ�=�V9�W'/��XF��:R�y�#�C����>��a?�L?��b>0���n3��!�"\ͽA1�����L@���,�@�߽�25>v >>�>��D���Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>F�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ta~����7�b��=��7?�0�#�z>���>��=�nv�ݻ��X�s����>�B�?�{�?��> �l?��o�O�B�~�1=:M�>Μk?�s?$Ro���f�B>��? ������L��f?�
@u@`�^?)�Aؿ:���褳��3����>��=�$�=Vi�%�=��=ks:=�#a;P>\I�>�d>U�> >��v>֮f>+�����c�����p�I�g�z�"�Buh���#�\�u���-���
���T���,��`������j/�٘<\,�=I�U?)�Q?}p?� ?�pw�Y>����w7=X�"��*�=�p�>[2?	�L?��*?L?�=&V��+�d��N���1��ݴ����>-I>ў�>*�>��>�	9KEJ>HW?>0��>Z�>x�%=)lݺ��=��N>k�>���>��>@���>���J渿.gk����tV >Ɠ�?U1�Ztg�0'��E#�n�Ҿ��~>kVD?��u�������ؿټ��I?{���c'��\ϖ>��%?:�B?3�Z>2���%�=�i��r�m�F��=��$=:]��[���!����0>,F0?kS�= ��>r)q��.P��B������j?��\?g-V�<�-����{�i���۽��>ot�>�ꕾm�<�
��Ь}�5;����=?���>HL{�B}\���\�G]��t�>�U�>1��>�Y>KE�<���=Er�=al >��V>��=j,X=�F?��">�c=�U�>�b����a�(�>m�U>E�P>F)?�x?�l,������Q���+�b�>N��>��w>���=�0���=��>��a>��$��vw�����a�}	<>�I�Q/j���=�2��=�é�ٶ�=$�=k�*��uK�5�<{~?X\��-������󟸽3�C?�?L(�=�t<�"�Ȭ��D㸾r��?��@w6�? ���V��?eߍ?1���g�=p��>fA�>�ξܡL���?;�ý�`�	�K$���?Р?*�(������ek�)�>�F$?Q`Ծ�p�>�h��W����Y�u��#=K��>�4H?1X��EP�>�1s
?]?�T򾠩���ȿ�~v���>�?�?d�m��?���@�V��>V��?�iY?Kpi>�b۾�HZ�x��>��@?s
R?�>B?���'���?l޶?���?��v>�s�?��?��>~d!<k�%�\�Ŀe^��$�E=���=C"�>�ق>H����aM����ax��$wd�_F�ȇa>;.-=���>��`��d;W�9>�Խ�稾hS���g�>��>e�g>`Z�>��?�Q�>�>�>`w8>��<����� ھ:�K?���?\��#n�%�<S�=��]�XG?3�3?G@Z�ܧϾ]R�>�z\?X̀?�[?]]�>Ͳ��7���濿d��̧�<��K>З�>B^�>�k����J>��Ծ-+C��Q�>��>MF����ھ���;A��e&�>6z!?���>��=�� ?|�#?��j>s/�>v[E�8����E����>���>�I?o�~?� ?�ҹ��[3�����桿֑[��:N>��x?�S?K˕>��������shD��II�����	��?�sg?�e�?1�?<�??��A?�=f>Xn���׾�ɭ�C߀>�W?uw�"�=�A��=�0���>�)?$��>`�D�F˽x�1��U���Ҿ��?�Z?�G!?��Md]��ƾ���<��=N�&��8j�8����>�>��d��љ=.�=�J�=E�K�d���x�=!�=���>���=�T�ܬϽ�+,?��F������"�=��r�GhD���>Z�L>Q���
P^?��<���{�x���~����T���?���?�[�?^"���dh��<?"�?�-?Q�>�+��ko޾ ��h9w���w�y�d�>�'�>
d�@�Mp�������:���wŽ��{��>!��>_�?��?�rc><Z�>ܟ���������T쾶�X�`v��0�B5����xȑ�S8��lO�<�<վN��>Н���>\4?�w>�CK>M��>�R�q��>g�>�<v>�ݢ>}�r>"u>��z>|��<Yཽ�wR?�����h&��F߾����#G=?�Oa?B��>mI%�ac�������?UL�?hq�?t�t>f�a��{+��}?���>T�y�Ln?$�=|���9����z�N�r��v���>׉��3�/I��X_���?_|?^�ؼ�Ѿ6��^���o=�M�?��(?�)���Q��o�s�W��S�����6h�:i����$��p��쏿�^��>%����(��u*=R�*?R�?{������ ��&k�I?��df>
�>t#�>�޾>jtI>R�	���1��^��M'�O����Q�>5[{?��>ÇB?�X?�	t?),x?F�>-x�=�u�"��>��S>H�>Fx.?2W)?� �>��?V�?KM8?%�>00���۾2v����>?�y(?9��>��>�������y>e���A<���=��<>� �=Ō,��O�=��^��t�>�./?.�Z�+�(��ھ�

>n%?"�?mR�>�������V^6��y�>��#?<��>�H:�tP��d�+ë>��r?�9"��S�<1|>~J�=�q>U*�}��=�\�r�>BM*>[�B=Q���e>�>@	W��n�>�9>�`>��z=~��>��?�
�>�"�>s���Ш ���xA�=�[Z>�P>��>�w׾ڒ���S���:g���|>?t�?��?��a=h��=Jo�=U7���~��iA��������<��?��"?�~S?W�?B�<?9I"?�>���t&��A���B͡�Ŏ?=/1?Mϖ>\��FD���띿��(��?�)�>�T�����{&��$�����+�@>�/E��E���l���,8�e�	=N�[*��O �?D;�?d��<ǃ0�i��OǛ�۝��K?Q�>��>��>�B(�9�Y���	��/>j�>��L?��>�pW?�ր?��d?T-�>/��Ʒ�#���,+�=?.>�T?n(�?ր?v�A?�У> >�;�VJ���!��9�q���R~"=Q�}>G��>T"!?h�>2�4>��8�y'�[gs�h}}=��q>�?��>���>I��>�ؼ��/?��>V��������������=��v?e�?�? ?مn=�
���X�Oo(�Ƣ�>�?�Ů?��?v�0���=zd0;��y��L�r}�>�<�>)�>�I=5sn=��t��ň>�\�>y�ƽ>�:���T��x=�?
_)?{�k=��ſD�q�� q��˗�;�c<H��:�d�����j[��}�=ɘ����!���I�[�������������������{����>���=���=���=���< `ɼ��<a�J=���<n�=�/p��On<��8��!ͻj����P���\<�vI=������ʾ�q}?�jI?�+?��C?�z>ȑ>h:���>貁�^c?H�V>u(S�Aü�*6;�+��H_��I�׾�N׾]�c������>�G�q>J4>�o�=��<��=13y=���=��\�D�=���=���=7��=5��=�G>x>5w?���,����,Q�ki��:?25�>n{�=Dwƾ@@?_�>>//��Ֆ���a�#+?���?�P�?��?@mi�e�>`�����V��=ם��<2>-��=��2����>��J>����J��s"��|6�?>�@��??�⋿~�Ͽvh/>��=��>��:��+C��9Qվ���=� B?�󾡰���o�>�=��(��N˾F��>�$�>n{�>MZw���C��=�ʴ�؇>.M=c��= V
>/��<(jɽ�Y>&ͼ(�>�i>خ�2˗�>��W��=-�O>�>�Ѡ>�v�>�G?PO?W�{?��?8z�tU̾f����X�>�#�>���>�O�>��U>��>6?�9?�<d?�>{�k>«>Cš>��
��dw��o� Ε��|,>��?i�u?��>���=�l����.�h<��P�~�>\Z=?n�;?^��>f��!�_%#���0�����i�;0����vz���ǽF�Ƽg�۽���{i>Jک>���>�>�>�π>/�W>m;�>���>�R	>bK7=�q�=��ݽܞû~��o�=q��c��釽��[��F�<��R�=|�;P��<=��=:�����\��=���>o4>���>#k�=`
��$R/>���N�L����=BB��,%B��7d��M~��/��06�~�B>�7X>~���/��i�?��Y>�n?>���?>u?'�>"���վ|P���8e��dS�ꏸ=ھ>	�<�gz;��Z`��M��oҾD��>�b�>AT�>6%�>��Ҿ�6��9������m&?�+��x����=�U?��U��Ě��ee���a=�AM?ׁ���	[��1�?�;G?���?�5�>�-]�(�8�7�?>=��� i>=���.��NH�X�'?�`/?ݏ�>�¥����H̾c���޷>�@I� �O���S�0�W��'ͷ�E��>������оd$3��g�������B��Lr�^��>(�O?��?t:b��W��GUO����(���q?�|g?>�>�J?�@?�%��z�r���v�=�n?ϳ�?O=�?x>l�=O;u�g�?*�?��?5��?�l/?F���3?�c>�-�>�+=�$>Z5>
2��ԭ2>��?�?��$?���M��j̾��ʾ�B���_>�;X=M��>Aݒ>���=0>�D)>,�F>9��>���>���>�Z>�5�>���>M`���N��;@?{z�>��>/�]?3PH�z���q5�=;��>\f>E��<R^�=� ��G"�.=�>윓:�v�>ce�>���>�ſ���?(ά>�����B?��
���E=��>�;b>áͽ�bn>��#>^*N>|�>��c>��b���>���=�X��sb+>E��z6�}�H���<�y娾Fi>�c���q����]���F��r�|����߅X�N+��9�A�e�=�t�?�����W�%�1����y�?4-�>�n5?#S���<���<��>�\�>�I��8�����K1ھn��?��?�:c>��>��W?��?{�1��3��sZ���u��&A�le���`�����j���B�
�}	���_?��x?xA?�S�<I9z>���?\�%��ҏ�**�>�/��&;��;<=+�>�+����`�7�Ӿi�þe;��BF>l�o?�$�?�X?�SV��aF��r,>ԑ<?y5?jx?�~3?��5?@9$��f$?h�D>�>?��??�6?Qr,?��
?<�6>0m >�-����T=�T���։�Kշ�P��9��(�6=�Uz=�d:��<H�D=���<������J�;u�����<תL=g3�=���=�ў>|�Z?�x�>5�S>h ?��-�� �8ԃ�gU'?�r$��Ib��S�E��gp"���B=��w? 	�?T�F?&6>�t)��6�D0>��c>��>>�V>�ǖ>����5����=�d�=�p,>��=</�k����D��ũ�<`��=��?ڷm>
=���s->�絾���%n>\N��ը��g��@�F�!�4M?�*�>��A?��?=0�;�z���ٽ�u�U���1?�w1?dl&?�b?Q��=tS����!�:^�EOc��v>�2=	��;H��L��#�=�l�o�r�>>�s��`�Ѿ�f>E/���m�.MY�J��Ű=l��O���&�T1�,�y���=�u>e���&� q��I���;�N?,=�_Ͼo��������s>ِ�>$H�>$sݽ.햼�"0����\ :>��>^`+>Y$���ھ�";�����>��D?�T_?�σ?F�}��3r�*BD�ʯ��棣������?��>$T?L8>c��=|������t�c�wsF�x�>�u�>-�ٯH����n���#�Ў�>�??kF>��?~�Q?b-
?��a??�+?��?f��>S��޻��?�ۂ?Ȅƻ��>��f,�q�@���,��.?x�?Z��tw>ƅ�>��
?�,?d�[?ʻ�>C�c>B����R��ј>��i>��H�������>ДM?cJ�>ǭ4?(m�?*�>,�����Ψ�=e�>Z�C>�C?��?��?���>1��>vN��@�C>�J�>Ûb?P�?�\?3l);��?##�>ݞ�>
#>؅�>�A�>�m?,�H?�l?��U?X��>J�G<&����
��=�4���<��<�&C=-S�;zn�=c��W���eR�-a�=�嵺��6<�p`=�'(<M.⼡��<���>N�>Qʳ��@>4/۾(�����l>�ә=zò��˕��>���5�:���>�>?R�>ǻ��w(�=��>)I�>?��,�-?$?�?1�=z^�I�޾yK��*�>ѫ4?X�j=6�j��f���te�}5>�c]? 3`?�գ�Z��C�b?��]?��C=��>ľN�b�D����O?i�
?]�G�V��>D�~?5r?���>vSf��Rn���1b���j��g�=>��>d,���d��X�>�7?���>D�b>�6�=��۾��w�:����?�݌?O��?�ڊ?�4+>N�n�g>�����[}��-^?dx�>ޥ�7�#?�g	�;�о_��r����������*���蕾���l"�hb��o�ѽ�6�=/�?Y�r?��p?�_?p��od��]�us�1�V�(���Z��E��MD�v�C��n�yj�(���������F=�<b�G�Z�~3�?�59?���n?"L����
�����S>㖁��B���d=����B��&�>M	?��xd�"W���?J�>�2�>:N7?�}1���J��/�O4��|
��I>�
g>�i>���>��B�
�?����ΰ��^w�Hi�T�w>��b?�PL?h�n?�"��D�0������!��/�j���C>Y)>���>��Z�=��H�%���=�V�q�*��Ӆ���	��y=wS2?�+�>M��>�+�?(?4:�����t��1��|<G��>�yi?�Z�>�v�>��̽M� �A��>/�l?���>��>�z��SO!���{�5>˽1*�>� �>f��>Wp>�,�(\��n������9�u��=��h?#���m�`����>xR?��: �K<@i�>�w� �!�J��'�'���>`v?e��=��;>N[ž���{�}'��l(?�z?�ב��(�k<�>��?���>2;�>_+{?=�>�����pW���?��a?@�G?	9?S��>�\g��
�2���)*"�oL=#w�>x(G>�Ƅ=��=6,��J���F��H�9>ޑ=d�r���JFf����ﳌ�B� =W�K>'u��; Y���Ӿ���1/��� ����ؽ(����(��������ײ�Fɔ�w~R<w�\�蟾�@����z���?�_�?����nվ�n���ņ���о��?����V赾�7��#E��#�侺��Jƴ��ؾ�g�֙��ބ��?����#�ÿkr���J�X��>/?:G~?l���k���[�le�<*7>�=Z@��Ŝ�U�ʿ����A?B��>+�̾�C��S�>��>���>�b�>#���~��j��;��?G�-?/?�!
�Aɳ��6��M�5>^��?@��@?��)���辋k=D��>	�
?��;>��5�Ӄ��Ϯ�s��>)�?�-�?1==ٜW�W���!�d?R�J<�2E��͚�=T��=�%=2�
��1L>>�>ȧ��/?�E�ܽ�k1>��>��!������^���<��]>qZн7̍�&Մ?�z\�df���/��T���T>��T?++�>;:�=��,?7H�Q}Ͽۯ\�+a?�0�?̦�? �(?xۿ�fؚ>C�ܾn�M?>D6?C��>�d&���t�~��=p:�3������'V����=8��>��>?�,�Ë���O��J����=Y���rȿ�O%��8�r=�V�����Y��%U�"ȼ�P���H���ҽlLi='�=K�,>0�e>�[m>@\>�FS?n3i?5"�>۰>.;�Kv��b֭��g�=�K��^G�=����Խ��ľ�t����¾pn�$�'���#�D;�)8x��P=e�D�������5��hy��D��?Y�>[X���Q�5j�ʱ�}��Y�8>"d�����U�S��}�eX�?G9?%\��?Q�����A�#���qM?�p>����[���$ȶ=��;>$ם��j�>��>#�3�7��\�O#?��)?2����9���,>d���2��=�y+?E��>�o�W��>��?a����w2�D�>�T�>���>m8�>vͰ�a;���ݽY?�"M?�1�Nb��<�X>����K#;���}=��<�G��ND=��g>Y�н���!���/����=�W?�Ս>��)����8�����r<=�x?fx?�$�>�k?��B?T,�<EE����S���
���z=l�W?��h?��>�8����Ͼ*�����5?�e?8%O>/?h�)�龶�.�ZC�a�?	�n?�?ؙ�\}��������U6?��v?�r^�[s��^��G�V��=�>�[�>S��>j�9�dl�>\�>?L#��G������ZY4�#Þ?��@���?8�;<N�曎=:;?�[�>��O��>ƾB{��v���1�q=�"�>Ì��Uev�����Q,�-�8?���?e��>򓂾����rH>��湭?8��?̇=2u_>�B�򇀿RX��z��>���=SF�=�M=
�L��xk�+��ľ��4�:>Q��>kq@u��<��=�T*���鿴�˿x;P��aZ�ܳn=z��>�9?CȤ=��˾�?�I���w?��DY�{����>K�>�I���䕾��v��,>�k���Mz�>W�F�C�>��\�=��r]�����<Y�>�`�>��>��۽
XǾ��?n����˿�\���|�%Z?c��?q�?��#?9p4�wE^��i���{���J?n�p?6 _?��Ӽ��T��.f�b�j?�G���H`���4��?E��U>
%3?�?�>\�-��C|=�>�q�>gj>�/�F�Ŀ`Ӷ�����#�?�~�?ed꾞��> ��?��+?�X��1��Q���.�*���~BA?� 2>�P��P�!��5=��璾+�
?r0?�F�#�/�_?�{a�x�p���-�1�ƽ'ҡ>D�0��\�jp���|��;e�?����<y�J�?^]�?Z�?�c��#�I%?��>{����0Ǿ}�<X��>R�>9sN>�_�$�u>���.�:�G�>���?>��?�_? ���=��c%>��}?"$�>�?9D�=�V�>q4�=�򰾄�+�Q~#>���=)?��?��M?�O�>�y�=��8��"/�rZF�DR�� ���C���>��a?#�L? Ob>y��N2��!��UͽEc1�SO��Z@���,��߽�(5>��=>->��D�Ӿ��?Lp�9�ؿ j��&p'��54?1��>�?����t�����;_?Sz�>�6� ,���%���B�_��?�G�?=�?��׾�R̼�><�>�I�>D�Խ����[�����7>0�B?[��D��t�o�y�>���?
�@�ծ?ji��	?�!��F���R~��w���6����=�7?�+{>��>��=@iv�I���%�s�ż�><�?�x�?���>(�l?,�o���B��1=}5�>��k?�z?O�_���qB>9�?������P@��&f?x�
@Ps@��^?�� ܿD[���ƾ5�����=�$�=Ԓ>��&>JVF�Ӱj�#�^�">Д�>�5>G&�>��>h>�I:>B;��Sg'������9����Q��U;���*��,���W'�O�|��?�����᰾���=�b⽜��X����X�ǲ��d"�=Q�U?	�Q?��o?%| ?�Nz���>5��R =$��=Æ>�2?��L?n�*?į�=�r��r�d�>`������Ƈ�2��>��H>��>f�>�>�ڹ��I>�>>D��>A�>��#=���'c
=5O>�"�><�>v5�>��(׮=b����㩿������ƾ9��q�?�پ�,;�gՒ���Ҿ��Q�I��=�/9?_��=���wjп!����c?�d��z�'���8��%�v�,?��f?菇>�۾7�K=,�;K�#�	�]��0>U�����Ӿ�5�5�>�2*?"�>>���>�(�����[;�QB��@n�>�F?4��%%l���u�S�j��R�����>s%�>0惾����~���h�-Zv���=�/N?���>�>m���� ��x=��9}�=ϸ">'؜=��=eA3=� R��߻�Ž�1<$g��פ�<��?-�0>��=���>� ��	7L��>�(E>U�+>Q=?�N#?�eʼn���*�����#���>\�>U��>���=b"E����=���>wee>7��9Ro�����x<��PO>�{�וa�
����~�=N	���o�=�w=(����<�.
5=Z�~?�}��W䈿`�`���AjD?�.?&�=��E<��"� ��^J����?��@�j�?ͅ	���V���?�?�?���ͼ�=�|�>׫>#ξC�L���?4�Ž�Ţ�Z�	�@#��Q�?�?c�/�ȋ��l�D>k_%?�Ӿ���>)���_��*���Iv��E= �>ĈH?����QS�"eB�$v	?c�?b��T���ȿ��v�-��>po�?��?lm�j���!l?����>g�?��Y?�Aj>R�ھ�Z�S�>��@?��R?��>��r�(���?8¶?��?o�l>;�?�{}?0��>��<n�!��	��
v���X	=v� >cE~>d�}>� ��{�Z��j��Y��9�\�K���d>E�=���>������Ҿ_=��𽜾��b���!�>d>hzM>�7�>�z�>�>��>߯=��Žǘ��𣵾�J?�Y�?o����n����<�#�=�R���?�}1?�^ʼ_{ɾ�d�>{KX?l��?7�\?�s�>}
�4�����l밾y�<�_U>�*�>���>+�C�!0N>=�ھ�u<��I�>8
�>�H�m�徇Ⴞ(�ƺ9��>��?��>�ҡ=2� ?e�#?�j>�,�>1[E��7��q�E�H��>$��>M?��~?�?�ι�m^3�����塿U�[�-@N>�x?BT?�͕>G���̃����E�TbI�S���؛�?�sg? O�?�1�?��??��A?�?f>~��ؾ彭�N�>��?�R>�!�������L{�>�D?S�>�Z���y�n���.5������/?PI?�u?�"Ǿ�G\�T����8=�x�P0[=�Ap<�_��[x>`Ց>q�{��(>��8�:��E�a�t�~��M�;�5���� >f��V���Ra�=M<,?8RG��ۃ��ޘ=�r�$wD���>�NL>X����^?�e=���{�����w��1U��?*��?Dj�?��(�h��$=?-�?�?<"�>UH��>޾��ྙTw�]}x�Iv���>6��>��l���吤������F���Žw[��g�>V�>K
?֬�>l�R>U�>���`�"�~P�R����\����u35��/�j2��}��5�!����$��b[��A��>�d��<?�>�7?��i>��z>���>�`ѻfs�>.`O>)�}>5�>,�Q>��6>��>���<%Nɽ?,B?�z��s6�GE���8㾪�!?��f?O�?K�(��h|��u�9��>/�?Y�?�&>��v�4r$�{��>��>����?�ع=�'�=fs�=���#"=�t���o"=1�O>�D��>��M�	�<���?���>�}>KY��X(��������n=N�?�(?�)���Q���o��W��S�ō�7h�Sh����$�S�p�폿�^���$��Ġ(�\y*=A�*?9�?�����!���&k�E?��`f>��>�%�>�>yI>�	�(�1��^��L'�����LQ�>�Z{?䘐>ڒB?7c??��R?d�N?M�>���>��r�>���<�d�>YE�>�7?ѻ+?D�-?K�?<�(?KRq>ك��
��7��^?�?+8?.�?�F?�w��/f���R'������w_��쏖=���<�ν�<���=B`>�(�>��ּ0_��S�����2u>�^i?�� ?��_��fO̽�tD=��d?��?S
�ӎ�6�-���a> �m?�������9�=�m>���Z꾽�������<��M�Ps�<>�y=W}�=G�Z=L�^=oR�6܇��.�:�Ӭ=T�/=�?�?D��>�6�>�Kz�:���H��*P�=CIj>�m>Y�5>O�Ӿ�1��Q���Xd�!N�>���?�õ?��=�6�=	��=$@��%�ɾ/2��̹�u\�<5o?��?)U?��?��:?r�?��>?���ב�؂�|l��P�?�b4?[H�>��ྜ���G�����4�?Z��>*�(�]��E8�����콇�=g�N���o��W��]a����= �j�>�^V�?��?�VT=��9���,��Ķ���j�2�j?�� ?�6?���>�eK�y1o�/F����=��?S?]��>h�!?v��?�d?�4�>����k������:n�;���>%�/?�z�?m��?K&?�H�>�G>���D\����ξ�J����q��%~��J >,-�=�Ы>;�?�7�>k�o>�CM��ѡ��A���ּL,?��?���>W��>���>0���G?I��>����ߎ�N=��ߋs�5@��=k?5��?��0?�q�=���:�G��b����>�ԧ?$�?5^0?j@� ��=~��̏ž�ɉ�y��>��>H��>o0�=�="(/>ˡ�>K��>[��,�6�?�Q��d?�ID? j�=� ƿ��q�2�p��ȗ���c<���We�����[�|Y�=�������Ω�^�[�&��������������q�{����>e�=���=���=���<E�ɼp��<\K={��<�=�*p��:n<�e8�^�ϻ<�����ү\<W�I=����U�žM�}?v�F?��(?��B?0#}>"�">�@.�_�>1���_�?�I>��w������:�wf���闾�:پ��Ծ�sa��u��R>O�E�s>�F0>��=͇{<'J�=�*{=�=P;�c/=��=WZ�=���=���=k�>��>�3w?����ݰ���4Q��M�2�:?g0�>���=&�ƾ@?]�>>�/��ӕ���`��1?���?�T�?}�?S�i��c�>|����䎽�X�=����l=2>h��=��2���>t�J>���WL���K��15�?��@�??�⋿�Ͽ�\/>,2>���>\���XD��B��J�������jX?����������>���>�<B��X���>8��>{�>Mvt�9@��ǅ=Ԙy��*�=e�)=�*8>]b>I�%����<;;�=ߨ=(B�=��>�H�:�))�1ξ;�S�=�	&>�.Z>��>���>�?];?��?7�?�"�<Pb������?�n�>�(�>�e>D)�>G-->��?�"a?/'v?4�?S�r>%?�>�'?�h�o�F�=���8[���a�<|vY?Y1o?*ҿ>@g�>��S�	-"�w�K�u����?�r?��?���>�V����EY&���.�������b�^�*=rr�hU����Wf�)���=Vo�>��>x�>0Ny>��9>P�N>[�>F�>���<rs�=�o�����<m˔��҄=�f�����<�mż�E����)���+��f��䃍;B݄;��\<�G�;q��=���>$<>|��>?��=���kA/>����@�L����=�F��]+B�4d��H~�i/�eT6�2�B>y9X>���3��C�?)�Y>l?>��?/Au?=�>��y�վbQ��|De��YS��ɸ=n�>0�<�vz;�Z`�`�M��{Ҿ�l�>
�C>���>ۿ�>H���g�ӟ)��"�,z�B� ?���,P'>���}�~�#ѳ�(̍�Fbe���=&u]? ���$�i��?�x1?���?�Y?W>�M{���X>�Jw�%�B>
��`R�n�����	?�^6?���>�r��>��(̾�追�_�>�MH���O�-�����0��q6�%��(9�>|r���Zо��2��h�����:UB�}�r�1�>��O?���?��b�`<���UO�ʿ��#��!�?ٗg?�_�>��??�󤽔��v����=Wo?��?k�?�W
>�O�=�2ʾz�)?�[2?I�?5�?��?p~��#?e�_>Q#�>��p=����S��	�u��>�a�>>�/?�T.?=¡�#�U���n��.���O>�	�>���>�m�>��O=����u�9~�=�Ws>A�>|i�>h��>���>I�>*�c���O�>�K?
̥>�M�>X�v?�AE=Gfc�t
�>��>ln�>0.:=2����ڡ���~���_>H3<т>DrB>�>S��ez�?%�>�����
%?�����/�d�O><um=濎��A�>�A�=���=ڵb>�7�>*>�і>v[�>mkؾ�5�=��@�)���Y���V������ܑ>���h|7�w�t�a� /�)��1p��c�\��]OJ������?��)�^��T���
�h@?��>N�@?�ۂ�f��Բ4=��>iϚ>����)+��}U���"վR�?���?Nnc>V�>!�W?|�?�1���2�LfZ���u�F�@�<�d�ֶ`��Í�����Ձ
����K�_?Q�x?c�A?:��<��y>���?�&�h����9�>�/��;�$w<=s�>	g���`���Ӿ�Eþ
���2F>��o?�#�?�9?�V�9�a��">�~;?�k2?�]t?p2?x�:?����$?d#9>�D?��?�G4?�	.?g
?4x2>���=�>���-=�k���3��ƞнŽ'���\>=��=�G����D<�=T�g<����=H���:�k��JX�<d�F=ד�=x��=j�>��\?˒�>�E�>��=?Ɇ��Z�.��h����8?:J>��\���G���@��T�	>:�p?�{�?��l?(��>���pn<��oS<%>e�0>@�`>\	�>J���nh����=ڹ >���=��=8f�Pc��y���zQ<>C&>��>׍>]���u�>P����)w��zq>��7�?��3�c�*C�݈3�Y�v����>�I?��?C�=h��]��?^��0#?=:?�YQ?�Vv?�Ƞ=s�Ѿ	�8��E�{�M��A�>,��<��
����������4��a�W2w>�萾�!���l>P�dn��k��
O����^�=E
��ָ<#6���ܾ٧���+�=#>�¾19#���"��\�J?`j�=�6���g�Է���>1�>�f�>)�b�3-��a�=�+˥�ڤc=T��>W1>Bv��ky澏�G��i��<�>\TE?�&_?�Q�?6#��4s���B�Hk������ɼ?2�><L?SB>�&�=&{�������d�64G���>:��>�����G�h%��E'����$����>xS?I>�?_�R?��
?҄`?#*?`?�&�>�:��p���.%?w�?'��=V�ӽZ�R�WG9�=�B�R�>�(? P�v�>�?��?�a&?I*R?*�?/�>�R���>�k�>�-�>�DU�m��xV`>d/H?��>�ZX?��?�|>
!2��8��K���a��=nS>s�+?b�?d�?���>e��>ں��u!>�n�>q^?{{�?��W?=�%=Q�?���>L�>�,=>�{�>Y�>�?��N?MR|?� _?��?I��<�o���9ƽa@����E��T]=:|��?"<0�<�1Ͻ����~����<}�<��A�Q,<@!��F�L�� =HM�>��x>q]��RF�=�gþ3톾��K>;�<��������A�M=��h>�x�>��>/B��D�����>�L�>���ڕ'?B��>�?�ڂ=�\m����i�p؝>��4?-�<%n�3$��,�q��f�<�a? �Y?�|����P�b?��]?qh�b=��þ�b�/�龏�O?�
?��G��>��~?��q?��>)�e��9n�%��4Cb���j��Ͷ=	t�>�W���d��A�>�7?�J�>��b>��=hu۾7�w��v��U?��?Z�?=��?.&*>��n��3����d�����Z??4�>iL��|.#?ȥ���Ͼ�����ߋ��|�Q�������:$���>������%��˸��$�=��?o?+h?;�Z?����qkb���\��Rz�:�X�/<	�N?�^TE��I���I�n�m�|�����M6����=�Rb�frH�'�?��,?\Y��q?�/��w��������x>5m��� �3>�s;<qC8=���=M,�%���m���?�I�>���>��7?b|]���9���:�9�D�@+�`e&>	x�>�B^> ��>�%e�Æ�����Ѿo���{�0Dv>�wc?��K?�n?'^��)1������!��W/�fk����B>�A>"��>*�W����:6&��R>�B�r�����l��U�	�-�~=��2?F4�>���>�K�?�?�y	� ���]x�@�1��i�<?�>.i?��>Iц>��Ͻ!� �D��>�Vl?�a�>�|�>�~���- ��ry�]5սц�>�,�>U��>��i>r(�|�Z��C��"x��WU9��%�=��g?h���^��$�>b�P?�� ;��	<���>����*!�i4�i�'��(>�3?~͘=N�2>s�ľ�L
�_�z�Uɋ��4 ?��?Lʅ�X!��YF>�X	?i��>#Z�>�`�?-��>@̫����Ip?��c?!N`?^l.?%�></�A;=�+ [�k�ͽ�=ϟ�>%�>��7;��=�.Ž_.s��E�Hi1<��n=�n�=�h��)P�<�+m��X�߻��bLk>�nۿLK���پN�w%�W7
�A툾�����u��#���]��
���]x����&���U�6c����}�l�ky�?�4�?G���%������蓀��������>��q�UL����t��9��ރ�>����`!��O�Bi��e��U?м7�S�ƿ�����̾E�>([G?��v?������3�8��ă=�Oݽ0�g=W�̾�\��R�̿Dl���b??���>Q��B�<˸�>��&>�L>gL�>E $������Һ=S�?��:?�?R�̽�g�������5{=Ռ�?#6�?W�A?�_(���龖�o=B�>l
?�%<>��3����_p�����>/n�?�ߊ?P�3=�CW���６Wf?�@u<�VE�0S��k��=⏜=?H=����M>D�>����B���ٽ�a1>ֲ�>�4�=��	^�!@�<{]>F ս�̑�5Մ?+{\��f���/��T��U>��T?�*�>W:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=t6����{���&V�{��=\��>c�>��,������O��I��V��=���5⿛C��ʾ>���&'�=��a��F�ԗ��H����!�ND����\�z��=��>5`�>�'�>��>iC?͐Z?Ӣ_>|
��}�I=��i��Q�����=e �������:��Y}��a�������оA˾���u����H����=դL�����!��r����I���/?�>+>��I�U�6V˽���6��c��=���)��;�O���{���?��@?�싿[Us�����=�ⅼ'�A?�� �@�
��ȱI>oz��0�:=�a�>�?=AJ����.��,L�&?!D#?�R�����3؁��H^� J9��B?�D?�;�G��>{�?箾F�;bY�>�gl>�S�>5�7>��h���`��0�;3�?j� ?,9N�!搾Wй>�}���V潊>��Ƚ>���~��=um�>F�t=U�Ҿ�G��8�ԇ�=�Ab?X�Z>=��Y_ɾ:Xa��#�=�Dq<2L?�?67�>czj?�^?|�>��(���V��'�Qޙ>�pr?��o?��=D������ST��U,?�l?�T>dG9�G���M)5�C� �;�>�Ƅ?1�.?����@��p���5?��v?�c^��]����fjV�4H�>6�>���>��9����>��>?#�"�g;���ǿ�S4�̞?}�@��?��@<܄�紎=~&?�@�>�P��Lƾo9���o��vks=���>2p��:v����n�,��8?��?)��>�{�������>)����3�?�-�?�b����>�d.���x��yB>ǀ>�'��>�Eɾ��Q�������ݾ����>�>@��%�k0?%)����P�ؿކ���+����5?���>�N3�|���ᤂ�k���W�[��Ȇ��"��SM�>��>�Ô�����`�{��p;��Ԟ��>�j�>a�S��&��`���\6<W�>ݦ�>���>L>��#罾>Ù?S_��F<ο娞���?�X?�f�?�m�?Kn?�9< �v�|�{�Q��+G?Ƅs?�Z?6y%�;]��x7�J�h?i����Y���1�l�;�|�M>�;0?�x�>��$���=9�	>v�>��>��)��ƿ�2�� ���?n�?���[k�>�q�?9�%?�������`=:��J��K?2�'>�r��i���@�D����b?
<.?�(�+��%�_?��a���p�k�-�l�ƽۡ>	�0��e\��=����;Xe����/@y����?;^�?'�?��� #��5%?�>����8Ǿ��<���>W(�>`*N>�G_���u>���:�4h	>���?h~�?Jj?ޕ������T>��}?R��>X��?���=���>�5�=����Ҳ��t>j�=v�<��?6
J?6��>N\�=�J�,�/�t�F�e4P��Z�M�B�v��>�oc? �I?Y�`>g���f�[�$�2Pѽ.y��l�u�A������'>QU9>�>SH�e�Ծ��?Mp�9�ؿ j��!p'��54?0��>�?����t�����;_?Oz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>;�>�I�>?�Խ����\�����7>1�B?W��D��t�o�z�>���?
�@�ծ?ii��	?���P��Sa~����7�V��=��7?�0�#�z>���>��=�nv�޻��X�s����>�B�?�{�?��>!�l?��o�O�B���1=9M�>Μk?�s?�Po���k�B>��?!������L��f?�
@u@b�^?)g�ɿm�D%E�3� ��.I���>d�=��2��g�=+��=�z����=(�>�D?�o>�wx>T�4>9�t>|H�>������(������ѐ��xx��5�b$�F�c�	���T���8��˕���>s���V�=����&`��������=t�U?��Q?��o?�G ?	({�e	 >&��;F
=0�#�!΄=�>gC2?*�L?g�*?��=�7����d�XU��?���BE�����>7�I>ñ�>��>�:�>ڮ+:(�H>�>>�$�>i��=$�+=�غ?;
=`�M>[!�>�*�>�ݺ>��<j�>�p���h��dM��Qʾ^l�=���?����^�l��3��[qξ� '�J>M�:?r{[� )���.п�H��'�U?M�R�Ǚ)��;�N:>m�3?��{?�%>$|ʾnJ>�ň=
/T��ן��g�=�+�;��zF1�n�z>s{?dIn>��>��M��L�,h!��o��>�J?�%��핾IS[�F�k�@��V�>���>b&u�:41������\��9�g�>4,?��?k�ؽOѾ��(�$Y+�Y>�@>ҽ�>2-w=�>bp=��="E�;��>���;�E���?oq=>�
�=��>�嗾��S��>��?>$D>2�9?�� ?���%�y�9Go����l>4��>er>p�=��>��;�=�>�cf>se˼I������I�7�OG>Bw���d��C���)�=�̡���=4
e=���uIQ�W�m=R�~?�|���㈿�뾩����jD?�2?
0�=��E<H�"�b���u<��U�?~�@k�?z�	�-�V�M�?�@�?Z���*��=/��>X߫>|&ξB�L�ݬ?T�Ž�â�ɒ	��0#��Q�?]�?�/��ȋ�tl�>6>�]%?��ӾD�>&b�pv��>��:3u�lC"=`7�>aLH?+w���S�k=���	?�U?.9�<����ȿ�v�	�>�{�?���?�lm��*��?����>�:�?��Y?}[k>��ھ�W�긎>�`A?VOR?e	�>b��'%��?�b�?&�?	I>���?S�s?�c�>jx� W/��0��F����=o�X;6_�>�A>0����aF��ؓ��h��m�j������a>�$=O�>I/�v5���E�=A���wK���=g���>%Dq>�I>�R�>R� ?]X�>Г�>)[= k��݀�����'�K?��?����n��
�<�Y�=�N^�2?�X4?��a��Ͼ���>�\?���?�"[?`7�>y���1���տ��/��>(�<��K>�;�>{?�>�ŉ���J>�bԾb�D����>���>�t���,ھ�>���κ�w�>G� ?(��>��=�� ?5�#?�j>�"�>�ZE�o7����E�ڳ�> ��>H@?��~?�?�й�oT3�:��硿ߐ[��-N>t�x?�T?�ŕ>O��������[D��[I�&䒽�?�qg?�2�l?�0�?&�??}�A?If>���ؾ7��@�>�?T�F��;���!��#��m�>x?��>(���O&��uo�&�*��& �F�?)1Z?�m?� �g}f���۾��<t=���=�ڻr�d:N��=8�>{ ��[=&�=}�$>e���a@8��׾<�>��>��>P�C�����=,?H�G�kڃ���=��r�awD�F�>$HL>� ��6�^?�h=�d�{�X��!y���	U�� �?@��?�k�?N��˝h�U$=?��?�?� �>�I��3}޾8���Qw��~x�mw���>���>v�l��徥���y���XF����Ž	�o�>,g�> 	?��?�5C>�.�>Q~�����)�.��^�Z�]��(N4��{2�3��9��+��%lX�b?��]����7�>8����>�b?�/�>?~>7��>����C~�>Uo>"��>��>�>>%hH>ض>TD�=��z���??5��;!�	\����� �1?��w?��!?
f���i�xʾ��>S��?ϖ?یQ>`gd�41I�k��>�6?�Ua�@�?�2I��N���q>]YҾ,i��������Ɛ>���M�a�Xg�}����<�>�K?��h��愾�����o=�M�?)�(?X�)���Q�8�o��W�-S� ���6h��k����$��p��쏿�^���$����(�}x*=;�*?��?|�� �� ��5&k�E?��`f>X�>�$�>r߾>sI>8�	�*�1�	^�M'�&����Q�> [{?��>�H?w�;?��O?�EK?�ކ>E�>ѯ�z��>�s6<���>���>v7?��,?��1?!?�k*?^aa>��З��*Y־�R?�S?��?2�?�?/.����˽@z��wW��8t�U�Y�;ņ= e�<�ݽ<���\=m�T>θ?%_}=>y&�I�H��=,b�>�/?���>k������3�c�}X>��?�[�>G�'��ہ��"��/k>��y?Z�=�ʟ��3>�F<��T�ļ�S�%�N���<ܤY>�㜽���<%�;>"<�k�9}�=�[2��� >g��  ?��?��>wH�>����+ �5�����=�i[>
4V>^�>=e׾�L���x����g�1�{>ȸ�?ې�?E�l=|�=GM�=Dנ�\5���D�X������<E?P#?��S?#`�?��=?=.#?Y�>������� ���Ѣ��?#])?�ږ>|m�w�Ծ柿)�&�o�?���>΅U�,���h������s ��%�>w�5��q��wt���;��#=pd��[��Oe�?W��?
ƶ���0����
���v1���I?�>���>&��>��&�^#`�b���<E>2q�>��E?�>�J7?;؈?u?a%�>C=:��8�����{1(>Qq�>�MR?v�?�Kg?�[9?x;�>\-�>H�Ǽ?�g���;�^2=xG~�tE�A�+<�u�>��>S��>׿�>K�=7f�=o������CD�=�B>�Q�>��>���>K��>& \�c&I?���>����{3	�����y�~��|R�yCr?�
�?�.?+gB=���v�C�\(��f�>u�?٬?&-?�QH����=nLü�����q���>��>K�>4�=��=�!>}��>3��>��(���4��6��E#?��D?���=�Tǿ�#t�¥q��-��vs�;W����i�qǕ��(Z�ظ�=�ޘ�}��K'��G�`������C�����F����ys��D�>�=�p�=�}�=��<YP�jй<��H=�d�<>l
=�\M���O<�.�O.�9�^n������Xu<�;c=ݰ���˾��}?N<I?`�+?U�C?ʯy>�->��3����>'��	A?5V>ӢP�&�����;����������ؾ�u׾��c�͟�0K>0^I�(�>F@3>ZH�=t\�<\&�=�2s=�=6�P�s=)�=DK�=id�=���=��>�R>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>jJ>P�>(�V�5�+�����<4��yW��bB/?J�@��g��73?.0�U�	��A�����>)z>oL>�V����� ]=b4�;��=�
N=+��=-@>�G�����Z��>���$�>�*?`�c'�Dc==p�d>`�;>�Ɔ>X�*>��?��>��K?��?#?ױѻ(E�����H�>�?��?��>3�>$e>����>$�?V�n?��?�=;D�>/dl>�L2��Ta������<��E>��?�mr?���>��ڽ��V������d� sA���?G'J?�X
?��>�>���`��M���M���a=�t���c��:���7d��~?��h����<$I>��>���>Xa>hIW>��>Uٳ>U�>��=vH�=^�=�f� ,��1=N=X�<te=I��=iu9��=f�=T��=�����";���=G���"��=���>�:>��>ꌖ=���E/>=���(�L����=�G���,B��2d��F~�;/�[6���B>�1X>�y���2���?��Y>0j?>���?;?u?1�>��8�վtQ��Ee�^S�鹸=�>&=�C{;�Z`�i�M��vҾ��>Fڕ>Kt�>'��>�u��W0�N�b�|�W����s?G����Tֽ˒��u���(��$����@I�.K��)�-?c�� �@���?8O�?�?�\�>�\�R��^�=̠>�r��<,/v�Is�����h ?;#7?��?ԀC���&�$ ̾W����z�>9(H��|O�w���)�0�Lv=�ƿ����><����о-�2�`o������zB���q��>��O?F��?�pc��*��Y�N�|D��م�'�?9�g?��>C�?�y?�����]쾐��W[�=�o?��?�R�?%o>u=qن�[�.?P�?8��?���?��\?���Ů>��>>5�<>���=��>��=�����;>���>
�5?��(?�?��G�h�ƾ=�쾪 ��b�>�B�>S�*?{ٛ>w`�>���=)����>���>ā?���>��t=,ش>�_�>��v�A�2?ќ>���>�OT?v��>>��<[�F�vP>���<���,b�;M��<�E��+-=$��S)>b�>��>9���/�?�"�>�8�O�%?9L�/���I�>��3>&�r��!�>�g>Pʳ>�>��>k�n>E
�>��Y>�Ҧ� {i>������o/��B��-�����>A�y� 8��n��Fa�?tK�Ñ���5�T�m�ʱy�N�?�C=��?�߽�if���-�d��? ��>q"?�*��5�ʽ)>uͺ>�Jj>�&侶Ȟ�OU��r���?
��?�;c>��>H�W?�?��1�J3� vZ�)�u�e(A�e�J�`��፿�����
���� �_?�x?%yA?�R�<:z>E��?��%�Eӏ��)�>�/�';�v@<=w+�>#*���`�k�Ӿs�þ�7��HF>��o?:%�?~Y?9TV�z�m��'>ҵ:?d�1?FNt?��1?K�;?���2�$?�{3>;D?Fp?�Q5?��.?�
?�2>��=�.���#(=�!��/늾Q�ѽ�gʽT��4=�{=�?�H<��=q��<���ټڼ;O���P�<9:=zܢ=#"�="��>��9?��?�:�>Y5?������1�����btO?�X�>@��P�<"����(@��%�=A�|?�Z�?ow?+ۚ>4����9�`U:=��O>�� �p> N�>s��p�T($<+>�a^>��=��9�yXg�@G�%��G6=��>�'�>D�>�+z�f*>����ӊ�`�\>۔'����B=w��AA�C.�p�U�`��>ΚM?�
?��g=K_���Ǯ�-HV��%?/?��E?3Rv?E3�=<�̾q�&��K�Kvp��l�>�r.�����Ԟ�ǖ���l@����;>�;W��!���l>P�dn��k��
O����^�=E
��ָ<#6���ܾ٧���+�=#>�¾19#���"��\�J?`j�=�6���g�Է���>1�>�f�>)�b�3-��a�=�+˥�ڤc=T��>W1>Bv��ky澏�G��i��<�>\TE?�&_?�Q�?6#��4s���B�Hk������ɼ?2�><L?SB>�&�=&{�������d�64G���>:��>�����G�h%��E'����$����>xS?I>�?_�R?��
?҄`?#*?`?�&�>�:��p���.%?w�?'��=V�ӽZ�R�WG9�=�B�R�>�(? P�v�>�?��?�a&?I*R?*�?/�>�R���>�k�>�-�>�DU�m��xV`>d/H?��>�ZX?��?�|>
!2��8��K���a��=nS>s�+?b�?d�?���>e��>ں��u!>�n�>q^?{{�?��W?=�%=Q�?���>L�>�,=>�{�>Y�>�?��N?MR|?� _?��?I��<�o���9ƽa@����E��T]=:|��?"<0�<�1Ͻ����~����<}�<��A�Q,<@!��F�L�� =HM�>��x>q]��RF�=�gþ3톾��K>;�<��������A�M=��h>�x�>��>/B��D�����>�L�>���ڕ'?B��>�?�ڂ=�\m����i�p؝>��4?-�<%n�3$��,�q��f�<�a? �Y?�|����P�b?��]?qh�b=��þ�b�/�龏�O?�
?��G��>��~?��q?��>)�e��9n�%��4Cb���j��Ͷ=	t�>�W���d��A�>�7?�J�>��b>��=hu۾7�w��v��U?��?Z�?=��?.&*>��n��3����d�����Z??4�>iL��|.#?ȥ���Ͼ�����ߋ��|�Q�������:$���>������%��˸��$�=��?o?+h?;�Z?����qkb���\��Rz�:�X�/<	�N?�^TE��I���I�n�m�|�����M6����=�Rb�frH�'�?��,?\Y��q?�/��w��������x>5m��� �3>�s;<qC8=���=M,�%���m���?�I�>���>��7?b|]���9���:�9�D�@+�`e&>	x�>�B^> ��>�%e�Æ�����Ѿo���{�0Dv>�wc?��K?�n?'^��)1������!��W/�fk����B>�A>"��>*�W����:6&��R>�B�r�����l��U�	�-�~=��2?F4�>���>�K�?�?�y	� ���]x�@�1��i�<?�>.i?��>Iц>��Ͻ!� �D��>�Vl?�a�>�|�>�~���- ��ry�]5սц�>�,�>U��>��i>r(�|�Z��C��"x��WU9��%�=��g?h���^��$�>b�P?�� ;��	<���>����*!�i4�i�'��(>�3?~͘=N�2>s�ľ�L
�_�z�Uɋ��4 ?��?Lʅ�X!��YF>�X	?i��>#Z�>�`�?-��>@̫����Ip?��c?!N`?^l.?%�></�A;=�+ [�k�ͽ�=ϟ�>%�>��7;��=�.Ž_.s��E�Hi1<��n=�n�=�h��)P�<�+m��X�߻��bLk>�nۿLK���پN�w%�W7
�A툾�����u��#���]��
���]x����&���U�6c����}�l�ky�?�4�?G���%������蓀��������>��q�UL����t��9��ރ�>����`!��O�Bi��e��U?м7�S�ƿ�����̾E�>([G?��v?������3�8��ă=�Oݽ0�g=W�̾�\��R�̿Dl���b??���>Q��B�<˸�>��&>�L>gL�>E $������Һ=S�?��:?�?R�̽�g�������5{=Ռ�?#6�?W�A?�_(���龖�o=B�>l
?�%<>��3����_p�����>/n�?�ߊ?P�3=�CW���６Wf?�@u<�VE�0S��k��=⏜=?H=����M>D�>����B���ٽ�a1>ֲ�>�4�=��	^�!@�<{]>F ս�̑�5Մ?+{\��f���/��T��U>��T?�*�>W:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=t6����{���&V�{��=\��>c�>��,������O��I��V��=���5⿛C��ʾ>���&'�=��a��F�ԗ��H����!�ND����\�z��=��>5`�>�'�>��>iC?͐Z?Ӣ_>|
��}�I=��i��Q�����=e �������:��Y}��a�������оA˾���u����H����=դL�����!��r����I���/?�>+>��I�U�6V˽���6��c��=���)��;�O���{���?��@?�싿[Us�����=�ⅼ'�A?�� �@�
��ȱI>oz��0�:=�a�>�?=AJ����.��,L�&?!D#?�R�����3؁��H^� J9��B?�D?�;�G��>{�?箾F�;bY�>�gl>�S�>5�7>��h���`��0�;3�?j� ?,9N�!搾Wй>�}���V潊>��Ƚ>���~��=um�>F�t=U�Ҿ�G��8�ԇ�=�Ab?X�Z>=��Y_ɾ:Xa��#�=�Dq<2L?�?67�>czj?�^?|�>��(���V��'�Qޙ>�pr?��o?��=D������ST��U,?�l?�T>dG9�G���M)5�C� �;�>�Ƅ?1�.?����@��p���5?��v?�c^��]����fjV�4H�>6�>���>��9����>��>?#�"�g;���ǿ�S4�̞?}�@��?��@<܄�紎=~&?�@�>�P��Lƾo9���o��vks=���>2p��:v����n�,��8?��?)��>�{�������>)����3�?�-�?�b����>�d.���x��yB>ǀ>�'��>�Eɾ��Q�������ݾ����>�>@��%�k0?%)����P�ؿކ���+����5?���>�N3�|���ᤂ�k���W�[��Ȇ��"��SM�>��>�Ô�����`�{��p;��Ԟ��>�j�>a�S��&��`���\6<W�>ݦ�>���>L>��#罾>Ù?S_��F<ο娞���?�X?�f�?�m�?Kn?�9< �v�|�{�Q��+G?Ƅs?�Z?6y%�;]��x7�J�h?i����Y���1�l�;�|�M>�;0?�x�>��$���=9�	>v�>��>��)��ƿ�2�� ���?n�?���[k�>�q�?9�%?�������`=:��J��K?2�'>�r��i���@�D����b?
<.?�(�+��%�_?��a���p�k�-�l�ƽۡ>	�0��e\��=����;Xe����/@y����?;^�?'�?��� #��5%?�>����8Ǿ��<���>W(�>`*N>�G_���u>���:�4h	>���?h~�?Jj?ޕ������T>��}?R��>X��?���=���>�5�=����Ҳ��t>j�=v�<��?6
J?6��>N\�=�J�,�/�t�F�e4P��Z�M�B�v��>�oc? �I?Y�`>g���f�[�$�2Pѽ.y��l�u�A������'>QU9>�>SH�e�Ծ��?Mp�9�ؿ j��!p'��54?0��>�?����t�����;_?Oz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>;�>�I�>?�Խ����\�����7>1�B?W��D��t�o�z�>���?
�@�ծ?ii��	?���P��Sa~����7�V��=��7?�0�#�z>���>��=�nv�޻��X�s����>�B�?�{�?��>!�l?��o�O�B���1=9M�>Μk?�s?�Po���k�B>��?!������L��f?�
@u@b�^?)g�ɿm�D%E�3� ��.I���>d�=��2��g�=+��=�z����=(�>�D?�o>�wx>T�4>9�t>|H�>������(������ѐ��xx��5�b$�F�c�	���T���8��˕���>s���V�=����&`��������=t�U?��Q?��o?�G ?	({�e	 >&��;F
=0�#�!΄=�>gC2?*�L?g�*?��=�7����d�XU��?���BE�����>7�I>ñ�>��>�:�>ڮ+:(�H>�>>�$�>i��=$�+=�غ?;
=`�M>[!�>�*�>�ݺ>��<j�>�p���h��dM��Qʾ^l�=���?����^�l��3��[qξ� '�J>M�:?r{[� )���.п�H��'�U?M�R�Ǚ)��;�N:>m�3?��{?�%>$|ʾnJ>�ň=
/T��ן��g�=�+�;��zF1�n�z>s{?dIn>��>��M��L�,h!��o��>�J?�%��핾IS[�F�k�@��V�>���>b&u�:41������\��9�g�>4,?��?k�ؽOѾ��(�$Y+�Y>�@>ҽ�>2-w=�>bp=��="E�;��>���;�E���?oq=>�
�=��>�嗾��S��>��?>$D>2�9?�� ?���%�y�9Go����l>4��>er>p�=��>��;�=�>�cf>se˼I������I�7�OG>Bw���d��C���)�=�̡���=4
e=���uIQ�W�m=R�~?�|���㈿�뾩����jD?�2?
0�=��E<H�"�b���u<��U�?~�@k�?z�	�-�V�M�?�@�?Z���*��=/��>X߫>|&ξB�L�ݬ?T�Ž�â�ɒ	��0#��Q�?]�?�/��ȋ�tl�>6>�]%?��ӾD�>&b�pv��>��:3u�lC"=`7�>aLH?+w���S�k=���	?�U?.9�<����ȿ�v�	�>�{�?���?�lm��*��?����>�:�?��Y?}[k>��ھ�W�긎>�`A?VOR?e	�>b��'%��?�b�?&�?	I>���?S�s?�c�>jx� W/��0��F����=o�X;6_�>�A>0����aF��ؓ��h��m�j������a>�$=O�>I/�v5���E�=A���wK���=g���>%Dq>�I>�R�>R� ?]X�>Г�>)[= k��݀�����'�K?��?����n��
�<�Y�=�N^�2?�X4?��a��Ͼ���>�\?���?�"[?`7�>y���1���տ��/��>(�<��K>�;�>{?�>�ŉ���J>�bԾb�D����>���>�t���,ھ�>���κ�w�>G� ?(��>��=�� ?5�#?�j>�"�>�ZE�o7����E�ڳ�> ��>H@?��~?�?�й�oT3�:��硿ߐ[��-N>t�x?�T?�ŕ>O��������[D��[I�&䒽�?�qg?�2�l?�0�?&�??}�A?If>���ؾ7��@�>�?T�F��;���!��#��m�>x?��>(���O&��uo�&�*��& �F�?)1Z?�m?� �g}f���۾��<t=���=�ڻr�d:N��=8�>{ ��[=&�=}�$>e���a@8��׾<�>��>��>P�C�����=,?H�G�kڃ���=��r�awD�F�>$HL>� ��6�^?�h=�d�{�X��!y���	U�� �?@��?�k�?N��˝h�U$=?��?�?� �>�I��3}޾8���Qw��~x�mw���>���>v�l��徥���y���XF����Ž	�o�>,g�> 	?��?�5C>�.�>Q~�����)�.��^�Z�]��(N4��{2�3��9��+��%lX�b?��]����7�>8����>�b?�/�>?~>7��>����C~�>Uo>"��>��>�>>%hH>ض>TD�=��z���??5��;!�	\����� �1?��w?��!?
f���i�xʾ��>S��?ϖ?یQ>`gd�41I�k��>�6?�Ua�@�?�2I��N���q>]YҾ,i��������Ɛ>���M�a�Xg�}����<�>�K?��h��愾�����o=�M�?)�(?X�)���Q�8�o��W�-S� ���6h��k����$��p��쏿�^���$����(�}x*=;�*?��?|�� �� ��5&k�E?��`f>X�>�$�>r߾>sI>8�	�*�1�	^�M'�&����Q�> [{?��>�H?w�;?��O?�EK?�ކ>E�>ѯ�z��>�s6<���>���>v7?��,?��1?!?�k*?^aa>��З��*Y־�R?�S?��?2�?�?/.����˽@z��wW��8t�U�Y�;ņ= e�<�ݽ<���\=m�T>θ?%_}=>y&�I�H��=,b�>�/?���>k������3�c�}X>��?�[�>G�'��ہ��"��/k>��y?Z�=�ʟ��3>�F<��T�ļ�S�%�N���<ܤY>�㜽���<%�;>"<�k�9}�=�[2��� >g��  ?��?��>wH�>����+ �5�����=�i[>
4V>^�>=e׾�L���x����g�1�{>ȸ�?ې�?E�l=|�=GM�=Dנ�\5���D�X������<E?P#?��S?#`�?��=?=.#?Y�>������� ���Ѣ��?#])?�ږ>|m�w�Ծ柿)�&�o�?���>΅U�,���h������s ��%�>w�5��q��wt���;��#=pd��[��Oe�?W��?
ƶ���0����
���v1���I?�>���>&��>��&�^#`�b���<E>2q�>��E?�>�J7?;؈?u?a%�>C=:��8�����{1(>Qq�>�MR?v�?�Kg?�[9?x;�>\-�>H�Ǽ?�g���;�^2=xG~�tE�A�+<�u�>��>S��>׿�>K�=7f�=o������CD�=�B>�Q�>��>���>K��>& \�c&I?���>����{3	�����y�~��|R�yCr?�
�?�.?+gB=���v�C�\(��f�>u�?٬?&-?�QH����=nLü�����q���>��>K�>4�=��=�!>}��>3��>��(���4��6��E#?��D?���=�Tǿ�#t�¥q��-��vs�;W����i�qǕ��(Z�ظ�=�ޘ�}��K'��G�`������C�����F����ys��D�>�=�p�=�}�=��<YP�jй<��H=�d�<>l
=�\M���O<�.�O.�9�^n������Xu<�;c=ݰ���˾��}?N<I?`�+?U�C?ʯy>�->��3����>'��	A?5V>ӢP�&�����;����������ؾ�u׾��c�͟�0K>0^I�(�>F@3>ZH�=t\�<\&�=�2s=�=6�P�s=)�=DK�=id�=���=��>�R>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>jJ>P�>(�V�5�+�����<4��yW��bB/?J�@��g��73?.0�U�	��A�����>)z>oL>�V����� ]=b4�;��=�
N=+��=-@>�G�����Z��>���$�>�*?`�c'�Dc==p�d>`�;>�Ɔ>X�*>��?��>��K?��?#?ױѻ(E�����H�>�?��?��>3�>$e>����>$�?V�n?��?�=;D�>/dl>�L2��Ta������<��E>��?�mr?���>��ڽ��V������d� sA���?G'J?�X
?��>�>���`��M���M���a=�t���c��:���7d��~?��h����<$I>��>���>Xa>hIW>��>Uٳ>U�>��=vH�=^�=�f� ,��1=N=X�<te=I��=iu9��=f�=T��=�����";���=G���"��=���>�:>��>ꌖ=���E/>=���(�L����=�G���,B��2d��F~�;/�[6���B>�1X>�y���2���?��Y>0j?>���?;?u?1�>��8�վtQ��Ee�^S�鹸=�>&=�C{;�Z`�i�M��vҾ��>Fڕ>Kt�>'��>�u��W0�N�b�|�W����s?G����Tֽ˒��u���(��$����@I�.K��)�-?c�� �@���?8O�?�?�\�>�\�R��^�=̠>�r��<,/v�Is�����h ?;#7?��?ԀC���&�$ ̾W����z�>9(H��|O�w���)�0�Lv=�ƿ����><����о-�2�`o������zB���q��>��O?F��?�pc��*��Y�N�|D��م�'�?9�g?��>C�?�y?�����]쾐��W[�=�o?��?�R�?%o>u=qن�[�.?P�?8��?���?��\?���Ů>��>>5�<>���=��>��=�����;>���>
�5?��(?�?��G�h�ƾ=�쾪 ��b�>�B�>S�*?{ٛ>w`�>���=)����>���>ā?���>��t=,ش>�_�>��v�A�2?ќ>���>�OT?v��>>��<[�F�vP>���<���,b�;M��<�E��+-=$��S)>b�>��>9���/�?�"�>�8�O�%?9L�/���I�>��3>&�r��!�>�g>Pʳ>�>��>k�n>E
�>��Y>�Ҧ� {i>������o/��B��-�����>A�y� 8��n��Fa�?tK�Ñ���5�T�m�ʱy�N�?�C=��?�߽�if���-�d��? ��>q"?�*��5�ʽ)>uͺ>�Jj>�&侶Ȟ�OU��r���?
��?�;c>��>H�W?�?��1�J3� vZ�)�u�e(A�e�J�`��፿�����
���� �_?�x?%yA?�R�<:z>E��?��%�Eӏ��)�>�/�';�v@<=w+�>#*���`�k�Ӿs�þ�7��HF>��o?:%�?~Y?9TV�z�m��'>ҵ:?d�1?FNt?��1?K�;?���2�$?�{3>;D?Fp?�Q5?��.?�
?�2>��=�.���#(=�!��/늾Q�ѽ�gʽT��4=�{=�?�H<��=q��<���ټڼ;O���P�<9:=zܢ=#"�="��>��9?��?�:�>Y5?������1�����btO?�X�>@��P�<"����(@��%�=A�|?�Z�?ow?+ۚ>4����9�`U:=��O>�� �p> N�>s��p�T($<+>�a^>��=��9�yXg�@G�%��G6=��>�'�>D�>�+z�f*>����ӊ�`�\>۔'����B=w��AA�C.�p�U�`��>ΚM?�
?��g=K_���Ǯ�-HV��%?/?��E?3Rv?E3�=<�̾q�&��K�Kvp��l�>�r.�����Ԟ�ǖ���l@����;>�;W��!���l>P�dn��k��
O����^�=E
��ָ<#6���ܾ٧���+�=#>�¾19#���"��\�J?`j�=�6���g�Է���>1�>�f�>)�b�3-��a�=�+˥�ڤc=T��>W1>Bv��ky澏�G��i��<�>\TE?�&_?�Q�?6#��4s���B�Hk������ɼ?2�><L?SB>�&�=&{�������d�64G���>:��>�����G�h%��E'����$����>xS?I>�?_�R?��
?҄`?#*?`?�&�>�:��p���.%?w�?'��=V�ӽZ�R�WG9�=�B�R�>�(? P�v�>�?��?�a&?I*R?*�?/�>�R���>�k�>�-�>�DU�m��xV`>d/H?��>�ZX?��?�|>
!2��8��K���a��=nS>s�+?b�?d�?���>e��>ں��u!>�n�>q^?{{�?��W?=�%=Q�?���>L�>�,=>�{�>Y�>�?��N?MR|?� _?��?I��<�o���9ƽa@����E��T]=:|��?"<0�<�1Ͻ����~����<}�<��A�Q,<@!��F�L�� =HM�>��x>q]��RF�=�gþ3톾��K>;�<��������A�M=��h>�x�>��>/B��D�����>�L�>���ڕ'?B��>�?�ڂ=�\m����i�p؝>��4?-�<%n�3$��,�q��f�<�a? �Y?�|����P�b?��]?qh�b=��þ�b�/�龏�O?�
?��G��>��~?��q?��>)�e��9n�%��4Cb���j��Ͷ=	t�>�W���d��A�>�7?�J�>��b>��=hu۾7�w��v��U?��?Z�?=��?.&*>��n��3����d�����Z??4�>iL��|.#?ȥ���Ͼ�����ߋ��|�Q�������:$���>������%��˸��$�=��?o?+h?;�Z?����qkb���\��Rz�:�X�/<	�N?�^TE��I���I�n�m�|�����M6����=�Rb�frH�'�?��,?\Y��q?�/��w��������x>5m��� �3>�s;<qC8=���=M,�%���m���?�I�>���>��7?b|]���9���:�9�D�@+�`e&>	x�>�B^> ��>�%e�Æ�����Ѿo���{�0Dv>�wc?��K?�n?'^��)1������!��W/�fk����B>�A>"��>*�W����:6&��R>�B�r�����l��U�	�-�~=��2?F4�>���>�K�?�?�y	� ���]x�@�1��i�<?�>.i?��>Iц>��Ͻ!� �D��>�Vl?�a�>�|�>�~���- ��ry�]5սц�>�,�>U��>��i>r(�|�Z��C��"x��WU9��%�=��g?h���^��$�>b�P?�� ;��	<���>����*!�i4�i�'��(>�3?~͘=N�2>s�ľ�L
�_�z�Uɋ��4 ?��?Lʅ�X!��YF>�X	?i��>#Z�>�`�?-��>@̫����Ip?��c?!N`?^l.?%�></�A;=�+ [�k�ͽ�=ϟ�>%�>��7;��=�.Ž_.s��E�Hi1<��n=�n�=�h��)P�<�+m��X�߻��bLk>�nۿLK���پN�w%�W7
�A툾�����u��#���]��
���]x����&���U�6c����}�l�ky�?�4�?G���%������蓀��������>��q�UL����t��9��ރ�>����`!��O�Bi��e��U?м7�S�ƿ�����̾E�>([G?��v?������3�8��ă=�Oݽ0�g=W�̾�\��R�̿Dl���b??���>Q��B�<˸�>��&>�L>gL�>E $������Һ=S�?��:?�?R�̽�g�������5{=Ռ�?#6�?W�A?�_(���龖�o=B�>l
?�%<>��3����_p�����>/n�?�ߊ?P�3=�CW���６Wf?�@u<�VE�0S��k��=⏜=?H=����M>D�>����B���ٽ�a1>ֲ�>�4�=��	^�!@�<{]>F ս�̑�5Մ?+{\��f���/��T��U>��T?�*�>W:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=t6����{���&V�{��=\��>c�>��,������O��I��V��=���5⿛C��ʾ>���&'�=��a��F�ԗ��H����!�ND����\�z��=��>5`�>�'�>��>iC?͐Z?Ӣ_>|
��}�I=��i��Q�����=e �������:��Y}��a�������оA˾���u����H����=դL�����!��r����I���/?�>+>��I�U�6V˽���6��c��=���)��;�O���{���?��@?�싿[Us�����=�ⅼ'�A?�� �@�
��ȱI>oz��0�:=�a�>�?=AJ����.��,L�&?!D#?�R�����3؁��H^� J9��B?�D?�;�G��>{�?箾F�;bY�>�gl>�S�>5�7>��h���`��0�;3�?j� ?,9N�!搾Wй>�}���V潊>��Ƚ>���~��=um�>F�t=U�Ҿ�G��8�ԇ�=�Ab?X�Z>=��Y_ɾ:Xa��#�=�Dq<2L?�?67�>czj?�^?|�>��(���V��'�Qޙ>�pr?��o?��=D������ST��U,?�l?�T>dG9�G���M)5�C� �;�>�Ƅ?1�.?����@��p���5?��v?�c^��]����fjV�4H�>6�>���>��9����>��>?#�"�g;���ǿ�S4�̞?}�@��?��@<܄�紎=~&?�@�>�P��Lƾo9���o��vks=���>2p��:v����n�,��8?��?)��>�{�������>)����3�?�-�?�b����>�d.���x��yB>ǀ>�'��>�Eɾ��Q�������ݾ����>�>@��%�k0?%)����P�ؿކ���+����5?���>�N3�|���ᤂ�k���W�[��Ȇ��"��SM�>��>�Ô�����`�{��p;��Ԟ��>�j�>a�S��&��`���\6<W�>ݦ�>���>L>��#罾>Ù?S_��F<ο娞���?�X?�f�?�m�?Kn?�9< �v�|�{�Q��+G?Ƅs?�Z?6y%�;]��x7�J�h?i����Y���1�l�;�|�M>�;0?�x�>��$���=9�	>v�>��>��)��ƿ�2�� ���?n�?���[k�>�q�?9�%?�������`=:��J��K?2�'>�r��i���@�D����b?
<.?�(�+��%�_?��a���p�k�-�l�ƽۡ>	�0��e\��=����;Xe����/@y����?;^�?'�?��� #��5%?�>����8Ǿ��<���>W(�>`*N>�G_���u>���:�4h	>���?h~�?Jj?ޕ������T>��}?R��>X��?���=���>�5�=����Ҳ��t>j�=v�<��?6
J?6��>N\�=�J�,�/�t�F�e4P��Z�M�B�v��>�oc? �I?Y�`>g���f�[�$�2Pѽ.y��l�u�A������'>QU9>�>SH�e�Ծ��?Mp�9�ؿ j��!p'��54?0��>�?����t�����;_?Oz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>;�>�I�>?�Խ����\�����7>1�B?W��D��t�o�z�>���?
�@�ծ?ii��	?���P��Sa~����7�V��=��7?�0�#�z>���>��=�nv�޻��X�s����>�B�?�{�?��>!�l?��o�O�B���1=9M�>Μk?�s?�Po���k�B>��?!������L��f?�
@u@b�^?)g�ɿm�D%E�3� ��.I���>d�=��2��g�=+��=�z����=(�>�D?�o>�wx>T�4>9�t>|H�>������(������ѐ��xx��5�b$�F�c�	���T���8��˕���>s���V�=����&`��������=t�U?��Q?��o?�G ?	({�e	 >&��;F
=0�#�!΄=�>gC2?*�L?g�*?��=�7����d�XU��?���BE�����>7�I>ñ�>��>�:�>ڮ+:(�H>�>>�$�>i��=$�+=�غ?;
=`�M>[!�>�*�>�ݺ>��<j�>�p���h��dM��Qʾ^l�=���?����^�l��3��[qξ� '�J>M�:?r{[� )���.п�H��'�U?M�R�Ǚ)��;�N:>m�3?��{?�%>$|ʾnJ>�ň=
/T��ן��g�=�+�;��zF1�n�z>s{?dIn>��>��M��L�,h!��o��>�J?�%��핾IS[�F�k�@��V�>���>b&u�:41������\��9�g�>4,?��?k�ؽOѾ��(�$Y+�Y>�@>ҽ�>2-w=�>bp=��="E�;��>���;�E���?oq=>�
�=��>�嗾��S��>��?>$D>2�9?�� ?���%�y�9Go����l>4��>er>p�=��>��;�=�>�cf>se˼I������I�7�OG>Bw���d��C���)�=�̡���=4
e=���uIQ�W�m=R�~?�|���㈿�뾩����jD?�2?
0�=��E<H�"�b���u<��U�?~�@k�?z�	�-�V�M�?�@�?Z���*��=/��>X߫>|&ξB�L�ݬ?T�Ž�â�ɒ	��0#��Q�?]�?�/��ȋ�tl�>6>�]%?��ӾD�>&b�pv��>��:3u�lC"=`7�>aLH?+w���S�k=���	?�U?.9�<����ȿ�v�	�>�{�?���?�lm��*��?����>�:�?��Y?}[k>��ھ�W�긎>�`A?VOR?e	�>b��'%��?�b�?&�?	I>���?S�s?�c�>jx� W/��0��F����=o�X;6_�>�A>0����aF��ؓ��h��m�j������a>�$=O�>I/�v5���E�=A���wK���=g���>%Dq>�I>�R�>R� ?]X�>Г�>)[= k��݀�����'�K?��?����n��
�<�Y�=�N^�2?�X4?��a��Ͼ���>�\?���?�"[?`7�>y���1���տ��/��>(�<��K>�;�>{?�>�ŉ���J>�bԾb�D����>���>�t���,ھ�>���κ�w�>G� ?(��>��=�� ?5�#?�j>�"�>�ZE�o7����E�ڳ�> ��>H@?��~?�?�й�oT3�:��硿ߐ[��-N>t�x?�T?�ŕ>O��������[D��[I�&䒽�?�qg?�2�l?�0�?&�??}�A?If>���ؾ7��@�>�?T�F��;���!��#��m�>x?��>(���O&��uo�&�*��& �F�?)1Z?�m?� �g}f���۾��<t=���=�ڻr�d:N��=8�>{ ��[=&�=}�$>e���a@8��׾<�>��>��>P�C�����=,?H�G�kڃ���=��r�awD�F�>$HL>� ��6�^?�h=�d�{�X��!y���	U�� �?@��?�k�?N��˝h�U$=?��?�?� �>�I��3}޾8���Qw��~x�mw���>���>v�l��徥���y���XF����Ž	�o�>,g�> 	?��?�5C>�.�>Q~�����)�.��^�Z�]��(N4��{2�3��9��+��%lX�b?��]����7�>8����>�b?�/�>?~>7��>����C~�>Uo>"��>��>�>>%hH>ض>TD�=��z���??5��;!�	\����� �1?��w?��!?
f���i�xʾ��>S��?ϖ?یQ>`gd�41I�k��>�6?�Ua�@�?�2I��N���q>]YҾ,i��������Ɛ>���M�a�Xg�}����<�>�K?��h��愾�����o=�M�?)�(?X�)���Q�8�o��W�-S� ���6h��k����$��p��쏿�^���$����(�}x*=;�*?��?|�� �� ��5&k�E?��`f>X�>�$�>r߾>sI>8�	�*�1�	^�M'�&����Q�> [{?��>�H?w�;?��O?�EK?�ކ>E�>ѯ�z��>�s6<���>���>v7?��,?��1?!?�k*?^aa>��З��*Y־�R?�S?��?2�?�?/.����˽@z��wW��8t�U�Y�;ņ= e�<�ݽ<���\=m�T>θ?%_}=>y&�I�H��=,b�>�/?���>k������3�c�}X>��?�[�>G�'��ہ��"��/k>��y?Z�=�ʟ��3>�F<��T�ļ�S�%�N���<ܤY>�㜽���<%�;>"<�k�9}�=�[2��� >g��  ?��?��>wH�>����+ �5�����=�i[>
4V>^�>=e׾�L���x����g�1�{>ȸ�?ې�?E�l=|�=GM�=Dנ�\5���D�X������<E?P#?��S?#`�?��=?=.#?Y�>������� ���Ѣ��?#])?�ږ>|m�w�Ծ柿)�&�o�?���>΅U�,���h������s ��%�>w�5��q��wt���;��#=pd��[��Oe�?W��?
ƶ���0����
���v1���I?�>���>&��>��&�^#`�b���<E>2q�>��E?�>�J7?;؈?u?a%�>C=:��8�����{1(>Qq�>�MR?v�?�Kg?�[9?x;�>\-�>H�Ǽ?�g���;�^2=xG~�tE�A�+<�u�>��>S��>׿�>K�=7f�=o������CD�=�B>�Q�>��>���>K��>& \�c&I?���>����{3	�����y�~��|R�yCr?�
�?�.?+gB=���v�C�\(��f�>u�?٬?&-?�QH����=nLü�����q���>��>K�>4�=��=�!>}��>3��>��(���4��6��E#?��D?���=�Tǿ�#t�¥q��-��vs�;W����i�qǕ��(Z�ظ�=�ޘ�}��K'��G�`������C�����F����ys��D�>�=�p�=�}�=��<YP�jй<��H=�d�<>l
=�\M���O<�.�O.�9�^n������Xu<�;c=ݰ���˾��}?N<I?`�+?U�C?ʯy>�->��3����>'��	A?5V>ӢP�&�����;����������ؾ�u׾��c�͟�0K>0^I�(�>F@3>ZH�=t\�<\&�=�2s=�=6�P�s=)�=DK�=id�=���=��>�R>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>jJ>P�>(�V�5�+�����<4��yW��bB/?J�@��g��73?.0�U�	��A�����>)z>oL>�V����� ]=b4�;��=�
N=+��=-@>�G�����Z��>���$�>�*?`�c'�Dc==p�d>`�;>�Ɔ>X�*>��?��>��K?��?#?ױѻ(E�����H�>�?��?��>3�>$e>����>$�?V�n?��?�=;D�>/dl>�L2��Ta������<��E>��?�mr?���>��ڽ��V������d� sA���?G'J?�X
?��>�>���`��M���M���a=�t���c��:���7d��~?��h����<$I>��>���>Xa>hIW>��>Uٳ>U�>��=vH�=^�=�f� ,��1=N=X�<te=I��=iu9��=f�=T��=�����";���=G���"��=���>�:>��>ꌖ=���E/>=���(�L����=�G���,B��2d��F~�;/�[6���B>�1X>�y���2���?��Y>0j?>���?;?u?1�>��8�վtQ��Ee�^S�鹸=�>&=�C{;�Z`�i�M��vҾ��>Fڕ>Kt�>'��>�u��W0�N�b�|�W����s?G����Tֽ˒��u���(��$����@I�.K��)�-?c�� �@���?8O�?�?�\�>�\�R��^�=̠>�r��<,/v�Is�����h ?;#7?��?ԀC���&�$ ̾W����z�>9(H��|O�w���)�0�Lv=�ƿ����><����о-�2�`o������zB���q��>��O?F��?�pc��*��Y�N�|D��م�'�?9�g?��>C�?�y?�����]쾐��W[�=�o?��?�R�?%o>u=qن�[�.?P�?8��?���?��\?���Ů>��>>5�<>���=��>��=�����;>���>
�5?��(?�?��G�h�ƾ=�쾪 ��b�>�B�>S�*?{ٛ>w`�>���=)����>���>ā?���>��t=,ش>�_�>��v�A�2?ќ>���>�OT?v��>>��<[�F�vP>���<���,b�;M��<�E��+-=$��S)>b�>��>9���/�?�"�>�8�O�%?9L�/���I�>��3>&�r��!�>�g>Pʳ>�>��>k�n>E
�>��Y>�Ҧ� {i>������o/��B��-�����>A�y� 8��n��Fa�?tK�Ñ���5�T�m�ʱy�N�?�C=��?�߽�if���-�d��? ��>q"?�*��5�ʽ)>uͺ>�Jj>�&侶Ȟ�OU��r���?
��?�;c>��>H�W?�?��1�J3� vZ�)�u�e(A�e�J�`��፿�����
���� �_?�x?%yA?�R�<:z>E��?��%�Eӏ��)�>�/�';�v@<=w+�>#*���`�k�Ӿs�þ�7��HF>��o?:%�?~Y?9TV�z�m��'>ҵ:?d�1?FNt?��1?K�;?���2�$?�{3>;D?Fp?�Q5?��.?�
?�2>��=�.���#(=�!��/늾Q�ѽ�gʽT��4=�{=�?�H<��=q��<���ټڼ;O���P�<9:=zܢ=#"�="��>��9?��?�:�>Y5?������1�����btO?�X�>@��P�<"����(@��%�=A�|?�Z�?ow?+ۚ>4����9�`U:=��O>�� �p> N�>s��p�T($<+>�a^>��=��9�yXg�@G�%��G6=��>�'�>D�>�+z�f*>����ӊ�`�\>۔'����B=w��AA�C.�p�U�`��>ΚM?�
?��g=K_���Ǯ�-HV��%?/?��E?3Rv?E3�=<�̾q�&��K�Kvp��l�>�r.�����Ԟ�ǖ���l@����;>�;W��U��N@e>�����޾):n��xG�q��7`J=����E=�_�˾;m���=��>��ľ;S!��V��v��H?V�r=S[��jZ��D���`>�x�>�]�>�@ѼT�����A�G&����=���>Z@>
���#��$�C�����`z�>�E?�a?Tt�?���1Xq�n�C�*���s��Ħ�o�?ޯ>sK	?1�H>m��=蹰����)d�&OG���>�L�>��:D�����	�����%�О�>��?�D$>n?��Q?�#?�B_?�)?И?W��>�9��}V��/�2?Pp�?)	�=Yw��+�#���7��jR��F�>-<?�Pٽr�w>�W�>]�?�!?ژ\?��?�H>�辠�C�SJ�>���>/}Y�����o>B�G?l�>�1P?��?n�T>�C:�+E���˽��L�=f�>Q�1?�I$?s�?��>x��>p���f$�=ƨ�>�c?�1�?��o?�U�=��?@2>��>��=��>g��>}?nWO?��s?��J?���>S��<�/��a;��OEs��EO�p��;�7H<��y=���,t�MH���<3�;�ⷼ�a�����ӲD��萼F��;���>��Y>X6����D>�2Ѿ2����L>��Y�)���u���2����=��>�?�>U�J��< =��>���>ҡ��2&?�?�~?ǫ�;8f�>��4ё�o��>\�=?�.�=��i�2���l��ר<��s?MjV?!j���C	�(�@?��e?�"���Q���ȾA�T��\k��4^?|?�>�o��V�k>=�t?�Ub?4x?�uZ�_�s��u����S��G$��E>�D�>(@��PX�M܆>�&?#̞>6r�> �:>֖��8zo�P,�P��>���?��?]�?��C>�ы���ῳ��� ,���^?���>w����"?B%�͛Ͼ{Y���u���ᾃ����몾����}���`%�������ֽ���=�y?P�r?L�q?Q�_?'e ��c�4*^��)����U��������E��D��oC���n�C��U���2k���=@=u�ʣ\�	z�?~�1?��S�V?&�R��������J,{> �u��0��>�s	�w�=��K=$@}�r>3�E̕���?��>1��>O#0?kf�t�4��?�%�,�y���\>S~>&h�>H	?��L;��F���ؽA���s}�����&v>�tc?̘K?>�n?^w��1������!���/�CX����B>�r>�ŉ>̀W�j��}2&��T>���r�B��ct����	���~=��2?�D�>~>�H�?��?w	��J��Ex�3t1�⇂<P,�>zi?z/�>��>��Ͻ�� ����>��l?���>��>���rZ!���{���ʽ$&�>�>���>��o>�,��#\��j��O����9��u�=$�h?���(�`���>�R?O �:��G<�|�>��v��!�|����'�!�>Z|?���=�;>�ž�$�|�{��7���v+?�?� ���4&����>�#?M�>�4�>��?_͟>�z¾���?��\?��I?��B?��>m�*=�����˽p�*�* 8=«�>�&c>Mj{=���=�j��'d�$�%��&W=���=��Ӽ���bٝ;�X����^<�c�<��8>��ٿ��<�SGѾe������������ʽ�ˊ����ه��<������8Zl����v;A�Y�/�(l��w�]��8�?��?򧆾�i����m3���+���V�>��$�
�¼���T����3i�D4ؾ������$��0Y�g�P�T�ҷ&?���Ѯ��Ϟ����mw?�_?k#y?5q�x��N�5�,B7>�f=�7B�M!����>˿󂓾��_?k�>�|��&ؽ��>tؐ>�`y>�H�>�|�ӯ��$[���%	?D)-?&"�>@g�6�ƿo����d�<�M�?��@��A?��(����TX=��>�	?
y?>)�1� *��ذ��R�>�4�?���?�#N=��W����tue?to<[�F���޻H��=�y�=��=߉�ClJ>�_�>f_�/�A�g�ܽ��4>U�>�H#���Xe^�j��<�k]>��ս����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�}��=[��>c�>,������O��I��U��=C���؟��:�o(��B	=b)��}�<��u�"B��y@��(_�*�9��A־%ޗ�q��~�>Y��>���>p-C>ø3?�g?No�>z�y>�0]�&�2���ƾ��M��y��򴽅�=�qƌ=罾�BM��� �Y������:.�����F�+>p�A�6]���"�-�q�d�:�_k ?{�>먪�o[5����=A)پ5���A"��L���]����"�A�S�ǰ�?N�<?h}�� N��]�}`��Y{�Y=[?�lc�����|Ⱦ)�7>L{�=�>���>٢���U�js3���,��u0?>Z?_����[��1 *>�� ���=�+?��?ڂZ<%�>K%?��*�C)��][>�3>Lң>���>�F	>;���P۽�?��T?��] ���֐>ch����z��5a=u,>z;5�C��`�[>�I�<�팾>�U��[��\�<�R?Y�>�/(�JW��Q���[��v?=�v?��?L&�>�yh?OE?o��<���X�T�E���W=q�T?Ki?r >pf���Hվ�Ҩ��4?��f?��`>��X����-1�����A?�Ar?�D$?�J8�+���m��E���;8?91?C'a��a��@j$�?���45>�z?
��>�aO�$ޱ><g?q�q�v���ÿ��1�M)�?�q	@a��?$=NW|�J��>�?o�B>ޛ��;Yԕ�������=R�	?(Ý��n�j� �뙵�t�J?��s?��>v9t�KN����=ܕ��Z�?��?����a�g<H���l��m��A��<�ҫ=?��7"����(�7���ƾf�
������ܿ���>�Y@Q轝)�>
E8��5��SϿ����[оeSq�k�?��>6�Ƚ������j�dOu�j�G�]�H������f�>�.>_ؽH��[�t�jS7���=t��>Zd���V>�DT�T����[�<��{>|o�>�p;>����+��k��?3�޾��˿By�����F�]?��?3݅?�?4+������ݿ��AaM=O�h?5��?�??�u���Ml�����e?�¯�4H�����E�Nf>��7?���>��,�e��=v�>���>�Z>�x��������ݻ���?�?_�޾E@�>⚟?��8?�i���=Ӿ#�@��2=2L?��=Aʾi<�n�*�@*��.b?,?��P��,�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�
i	>���?�~�?Qj?���� ����U>
�}?2	�>�}�?���=���>?��=������8">pG�=�)��e?2�J?69�>�9�=��=��^/�3�E�3|P������C��P�>X�d?��M?�zd>6�Ƚ4�K�޹$�=���{.����D���7��5�M�*>,�G>��>�K���׾I�>>kO��+ٿ����Ʃ�?��>R?	f�|Fɾ\+�=�
�?V}>�H(�y��S�n��T��ڤ?��?��?Q���Z���]p��?s>ȫd>-ο�j�8�����
>g�?�b>�Z���q��j�]>�x�?_6�?3��?B{n���>�u0�
���Is�Z�Ծ�C��D��=Z�"?QO��׺=��?�g>���A��[ƅ�ۂ�>p��?3�?�I�>�7a?Fb(���0�=��'�>�rJ?��9?���d!�-�>Q�$?��9� ���f���*i?��@�@��l?����ҍ���+�������S�H�>٩<��6>�^n�e��=�;=>H>��>A��=�Ē>P$.��#+>ժO>��b>�ϴ>�V�d;�ݾ��(���$(�m�B���:�e=s�����)ն��=�$�ӾI�g�ڊžl�,��J�<w��g>��=~�I?f�Q?��b?���>ɧ����>v�m����� ��|�=]�>˝,?	U>?�=?��'=����X6k������J���͢���>d�g>d��>H<�>�(�>�ҋ��'>�-�>9xd>�h:>��=~я�xw�[��=| �>�Q�>HO�>�7;>�>˅���&���!h��lv��nŽ�?#����K�������D���=�/?M�>����/п`}��6~G?�[���"��(��S>�z0?a[U?�F>����sX��4>s���6k�*� >س�� mc�o>(�� F>��?�G>M��>�>���7�<�X����
a�=K�F? $�U�ξyw��~S�L�&�F�>]�6?�9}=�)��ɬ��e���)���'=Ø@?x��>� ���˾�^���æ��&>嚞>/	�;>b="A>�����F��`T��N>1[>M��=R`?-_)>*��=���>ӛ��Q�l��>��B>))>��??�e$?�n��ً�콁��/��iq>���>�W�>�5
>�LL�́�=֘�>~�f>�3�z��ߔ���G�q�Y>�"t�q&a�>�5�w=������=.�=�����?�p;=�~?���&䈿��9e���lD?R+?~ �=U�F<��"�C ���H��E�?p�@m�?��	��V�>�?�@�?��>��=}�>׫>�ξ�L��?��Ž/Ǣ�˔	�)#�hS�?��?��/�Zʋ�=l�|6>�^%?�Ӿ<�>F���6�J0����n�HI���> ??E������n4�oA)?�l�>d��G��~�¿��u�;�>��?5��?�R�`:���C����>[j�?�s?2h�>�p�u����0>��-?��j?�|/?����혵���>�1�?o�{?3I>���?Z�s?H��>:�w�ZP/�4��1����I==_d;�q�>ֻ>����5=F��̓��[�� �j���(va>}%=��>�C佦���02�=�^��gh��S]f�/��>�}q>�I>�]�>h� ?/b�>���>vK=�r��V���(�����B?�Ə?Q�	�4�j�{)�8�=��d��<?�2?iV�������>�GY?�?��b?a�>�$�v𜿨$��:尾tX�<Et^>���>%��>�D��r�G>9U޾�$p�~�>�:�>?{̼�澐�����.��Q�>4S"?���>tz|=��?��#?k�i>?�>�dE��J��$�E����>��>�%?<g~?Zp?Ƒ����3�p��'����e[�Z�M>��x?a�?at�>����}a��}+A��?�J|��њ�?̲f?�E��O?�?k6@?��B?��g>���]ھ�ƭ�^ׁ>m�?]<\C��5���"�/��>i{?q-	?jg�a���ڍ�t���̾ �?Jx?�e?0m�@�P!پM.�<�,�>�X=�(�=��8>��B<��˽�P>�"%>;��;� �A�LJڹ=��=f��>�]>\�������>ޝ#��	þH��LH�N[����>��;>i����yK?J���cu�H���ȟ�?�w?qL�?g��?ƫѽJ�e���6?A�?w[?��>ٿ��ؾ3%㾚Od�$�t�$�Z�>�x�>Ձ<=�պ�:퟿ػ��̇�C׽�~#��0�>
"�>z�?���>SӚ>���>�u̾&&�����	���Z��G�A�"���7��/�����)��~�<.����&����i>ķ���j�>\49?�\�>yE`>���>Tx��s^Y>:�R>�f!>���>=�>��>@�=�S_=��½��N?�a��"(���㲲�O>?k�e?Q��>����\��4��,&?�?Vݛ?��>�h���-�r� ?��>��v�N�	?׽\=�3�
�2<򓴾T
(�go���Z��7ȉ>d-�'�<�HJ��]�@?��?$�y��{ྍ�������_=���?x� ?:q-�ܚO��~l��S���P���<���y�������Ĩj�Y^���T��񀿍�)��Z<TL*?���?������������k�eR=�Y=�>$�>��~>*-�>R�T>����o0(�^yS��*��S���T�>]~?}V�>�p7?��4?2Lc?�_v?���>e�[>��ξG;?�G�<*�>�?�>��3?A�&?Ξ)?)K"?��*?�_X>bY�����9�~?�%?`�?w4�>`�	?.$���:�_'��'�l<����jѽ��=_�.=K���ŵ��1kl<1pz>��?��k��Q��ܾ��g=V�.?�?Vh#?R��yoþc�>�
?C'?AQ�>\H�|d��"��j�>k��?��ѻ/��<3>k�>�g�=.=�4z>#};-+=� ��n�=!U���>&=���=J��eB��$;x =�>)�>��?��>�>K���� ����H(�=��X>:0S>K>_پr}��L2����g��by>Ov�?:o�?�f=���=�=�e���N��k���� <�<��?}]#?�WT?K��?(�=?^|#?f�>o)�dM��&i��"��V�?�~+?�ۑ>�9�P\ʾ5���8]3��/?��?�	a�����(���¾��ҽ�>T�.���}����l|D�D����������dd�?V��?��=�E�5���o��G��A	D?�"�>⁦>Hi�>��)�C+h�U�F�;>�3�>��Q?�6�>]�m?�ϔ?jC�?�˹>�>��4��ಿF�<�=�>k�L?Q�?j�?���?B"�>{�R>��p���f��'��<tU��a�U�->/�>{�>�ߎ>�7Z>W4
>|F$=����Q�1�H$3>y��>r��>�>_�C>Ofѽl�b?f`?6E���t��|4�Asr�%�[�G$e?���?�M?�\���>���7�D�޾�� ?>,�?��?P-?�$���J�=&=���N���L��>0��>r,�>d���5�=V�$>�Ը>��>�	�ڒ�T�D�s*<Cl?Dq<?�D>}��\�^��!�����u恽�Ӕ���b�+"�Q���%>���2���w��Z^q��K��@ؖ�(����L��L���e�>1zj=��%>�>�=y>+=�.�9=�m�=dui=�� =u+�`�=�'7<�,Ӽ��觽F�L�Wo�=�"�=�e̾kax?��I?dT)? ,;?e�t>�>�>����>dh8��?��V>@�0�R(��2%:�3"�������߾.U޾��]��C���u>~d@�o�>��->���=�t�<a�=���=Q�Z=�-<
?4=D3�=��=�k�=F/�=>�>�6w?X�������4Q��Z罤�:?�8�>e{�=��ƾq@?��>>�2������zb��-?���?�T�??�?@ti��d�>K���㎽�q�=M����=2>n��=w�2�T��>��J>���K��B����4�?��@��??�ዿТϿ3a/>��
>�z�=%�Q���3��%Y���}���I��w?9�>�5]ʾ/�>�Q�=*���Ѿ,�=p�E>s��=���!�V��f�=�b��K�=� �='�>"�R>B�=TܽqI�=d =�:�=.QY>_��<��L�����ܹ�<X��=��6>b!->��?���>I=L?��?�`�>G��DY���оY��>��>�j�><����L>�k�>��@?}�<?�t*?�
�>0�ɽ��?�#?oaC��r��-o����3��Q+�?�U�?��>�ii����=�?�VQ��M�=4�?��?7-)?&Z>�U�m��,Y&���.������$E�f+=jnr��XU�E����k�����	�=so�>���>�>VUy>��9>��N>L�>T�>�>�<�r�=
ጻ�ʵ<���j��=������<�pż:��^&���+����l��;���;�]<���;k�=~c�>�N>w��>�#�=�����/>3Ė���L����=x����B���d��V~��.�-�4�ĻC>,cY>�?��|����?��Z>��@>40�? @u?� >�c� �վ�A��nd��WR��κ=�>b�=���;��V`�M)N�6�Ѿ���>��>�ۧ>�z>sQ-�@�>��Ȃ=�RܾhE3���>�\���<���i��z��������f�u",��E?����:��=��?~+M?�?���>8�����(�<>�{�$�<yr�|s��'���h?1�*?���>N��7H�{L̾"���ط>�DI�~�O�4�[�0����η�@��>g�����о�$3�ah�������B��Cr����>{�O?��?0b��V���TO����0���q?�zg?��>|K???�*���z�=t��^u�=��n?h��?<�?� >;�~=�K;���?��?
Ǉ?�I�?T�?�����a�>d���R�q=f��� >Фj>���<j�!<R��>6Y�>۹
?}�]�'�$��R�C4Ѿ��M����=A!<>K|�>*=�>�%�>x�z>�`P=�N<=w�u>j��>�ך>ڕG>剒>�Na>�:��[�(���,?}�e>�v>o�K?~��>/2=�y�3����=�-<��r�S���Ve��g(ǽ-�;Xɚ����<�<��>�zȿƔ�?��V>��(�r��>C���%���0>b��>mqx�6��>.=�>L�;>���>�<�>�'>Q/]>4��=�S��蠷=P���4����[���I�O�߾��>ϸ����۽�� ����<�л)D~�������z�r�z�&+�U�=��?B;��ry��o)���(�n?��>�GD?�2w�Ťͽ@�2>5��>8��>Q����h�;���ə����?"��?zBc>��>o�W?�?f�1�<3��vZ���u��%A�=e�ʺ`��፿h����
�:����_?�x?{xA?�0�<�?z>��?��%�g׏�p*�>9 /��(;��e<=�1�>�'����`�ĲӾ��þ�:�WOF>g�o?�$�?�Z?6WV��ck�B�#>)�:?�2?5t?F3?:T<?���hi$?�0>u}??�
?��4?%/?�^
?_>0>rv�=ns����,=�ᐽ#n��Q�Խ��Ƚi(���4=*�=Ŕ�:�o<�A=���<f��r���N;9��� U�<��9==o�=���=F+*?-U?R��>l��>Q~�?�x>�a��m��؇?�g�>��y�P+��F�^���NL>yJ�?��?�bH?��n=G�J����[>��?�?���>�K�>����V̾�a��%�>$��><�K>��<�ӫ���Ҿ5�t������q>f��>�A�>0,��O�=�M�x���̢;>��A�����z��A;�H�2�G�I����> �F?��?�$9=&V���g�|�a����>)�@?B:R?y�e?Vy
>Vخ���a�k����N��>�9>�l�X7���b��
?�^w=�r>�k�&��K��=Mh8���;J���*�P�����"ͽ�
���F=߾����ྋ�:>���~��_2Ҿ����ڳ���5?�~�>�h��.�㾷���g)��>���>��=u�@=;�������@�;��>1��>-Y��+��9��eվ`�>P�J?�Rw?jU�?j臾Īd���g���1�l�z�	��=�'?�>0�?�>��=�������=(_���E�Z��>�_?(|꾨�2�sA�����ƵD�Ά>�T?E	�>o�?,CQ?�E?BiU??]$?��
?� �>�S޽���Q'?� �?���=��ս�L�S8��jF�Ч�>�F,?e�5���>��?�?��%?)�Q?�E?�>���.�?�㖖>���>vY�yk���Z>��H?�z�>��Z?e��?�O=>5�e�������\�=��>S{1?~Z$?�'?�,�>��>fϾ�@>%��>�_?���?^hl?��<η?��>�?�v=@Z�>b��>A�?�T?{Au?T�B?9�>�<���Vzm���<�;:��<d2<��=l&��Ɠ��3�<Ȑ=D��;r+69X[ =�X{�zĬ�He<O��=���>Yh>y*����%>z۾R���^V>X�;33���$�"�4�	�=��>M�>�>y�6���=��>���>���h&?�?_�?�A=��8\���׾i�h���>��C?&T�=��j�[���%�l��Ѕ=:�r?�)Y?ԓt�H��"V?�fQ?��	���;��T����z�����'\?��>C@��>��N?�pe?MQ
?q���xm�6Ȕ�u`T�K���$�=cؙ>UL��Vy��ߍ>5�(?�IN>��>ر[>�ؾ�a�S���M�>o�?C�?��?�g�"O����꿡��ߴ��[^?���>�����+?U��:kVҾ ����*��UѾak��D:��)���_잾W� ����c"̽�x�=>�?��t?��q?�[?���9�b�h�`�G�~�DY��	�[��A���A�`=���f����4����o���� =�vi�$tH�'��?J�.?d��6?��������䂽��V>��x�J�4��<�=������=.�R=Y�f���P�����?$��>���>�3?�#_��q?��d<�k�8����qz�=��>Dd�>�M�>ߒ�<����O�
��1���+��pv>hc?Q�K?��n?*��X�0��{���!�l.�����G�C>�>���>��V�ɉ���%��>���r�z�U�����	��|=�h2?'�>�n�>2m�?�	?�8	�Q���dZy�5K1��!l<T��>��h?���>ޖ�>>Ͻ�� ���>��l?3��>^�>�����V!�~�{���ʽA"�>�ڭ>ܴ�>
�o>ҟ,�: \��i������\9�Lz�=�h?̆����`�T�>AR?��:�H<���>��v���!�$���'�|�>�w?���=h�;> �ž\%�F�{��5��ӛ(?L�?���	-�a�>��?�3�>cg�> �?���>J;xu��^c?�^?xM?N@?O+�>%<.m߽~ʽ�����b=:��>�GM>5H=B�=����eJ�T���!=��=�W��aѡ���;�����e<��=9'2>�׿�(Z�0	�B�ݾ�ھ6����␾�T�%h��n!`����現�����������S1�.�0���%���\�?���?,���73��O���,�u�7����|�>��i�ܴ��4�پw��m���׾|ྮ_��)��Ko��h��$
?�AG����������9��n�>��?_E~?T����.�.�3�}�^>'�$��i'�vL��П��p˿�q���`?Y}�>M}���ݹ�>Fy�>��0>D>7>�(i�h��n%;�[?w�I?��>����"nܿ.l����<�T�?tx
@�{A?;�(�M��P�U=E��>�	?g�?>eB1�II�)���BK�>�;�?`��?�%M=j�W���	��|e?��<��F���ݻ�=�a�=�u=Q����J>�T�>i���WA�2"ܽ��4>�ͅ>˅"�����r^�4�<|�]>��ս�]��5Մ?){\��f���/��T��U>��T? +�>]:�=��,?Z7H�`}Ͽ�\��*a?�0�?���?#�(?<ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=c6�h���y���&V����=\��>e�>,�ߋ���O��I��V��=^��1Eݿ}4�F���$�>'�ݼ��j���
����u[���6���,��x��>��K>D8@>�@�=:�=�=�ya?y�u?<O�=��>>ho��m�}쾘Q
�,&��%8�x#4�_�������";_	�ʢ��������I�?���[=�UY�������2�4�h�6�&�?�c�=x׾6-F��{��
��)ㆾ�<����������D���x��[�?)�O?�.m���f��m����� �A��^?����:�X%پ���=)��-=�Ӫ>��=ȶ���#��E:��Y0?� ?j���bݑ��k&>߫ �:8=c,?=?T<�>d�$?�m'�KX߽I�[>��/>"Y�>1��>s�
>�䮾MR۽C�?�;T?���l���d�>ɛ��I&{�'i=J�>�4��ܼ�Y>F
�<���TN�����޽<z�O?� �>՘ ��.���9���t�=�с?�F�>��P>��a?�1??���<C'���2��� ��r��u[?I7f?U�7>���ԯ��Ư���/?-"g?��>B�=	پ��!��1ؾ6�>ܥy?�L??��=�l��Ɂ�-���@{0?�2Y?ү/��@�����"�c��T>�)?��>%8M��V�=��>�O�>x��_%Կ=�b����?� @�V�?���=��ͽxվ=c�?�?+W��3q���սX��ui	���> ���X��!S)�н$#?��j?��?���w��%� >Ȕ��~��?��?�Ƙ�a�X>z�~�}������<$IQ>��ý�c/=Z�ɾ����b��u��vq��:,�>K+@�p=���>��r�=����7࿾���X箾:+�Yw�>3o�>�0
>9���WM���A�l(=�2CQ�i}۾���>.�>۞��N��ey�2�:��du:���>�OK���>XQ�����]����<:\��>D^�>���>�h���Ū��B�?����/eп����� ��:U?���?�܅?W�?'@^<��Z� ���Wt=��W?llw?�oJ?&2��sak��N)�C�g?�����P��g-��&M�.j\>ž6?�><)��}z=ą>���>%G>�%��ɻ��G�����K�?5)�?Z��B�>�i�?;�#?��0�\N������"G(�׿���CK?��>f�Ӿ�����1�x�t�t�?V,?��V��m#�]�_?)�a�M�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?ֵ�� #�e6%?�>c����8Ǿ��<���>�(�>*N>[H_���u>����:�i	>���?�~�?Pj?���������U>	�}?�Y�>g��?#>���>S�H=�a���<�y>x��=T���u� ?��D?�l�>?�=�<��K,��@�f�N�����aD�y��>��f?�O?&�l>�?��?q���+��ݬ���P�Tһ���0�j�{�vн��%>�;>n->pX/���ؾ�*�>n�e�̿J���C?��g�>�\�>��?(��R¾rV��ԟ?h�8��f�haͿ��r����jw�?M��?�?죾���<:i1>3��>>Y?���=f	y�G_����=IG�>�P>4��ن��{�>q��?�)�?���?�aT�F�?�_ �鴈�瓀��N����6��>-&4?gO���U>���>�m:>�I{����Fz��a�>�ȭ?��?��>�Xh?Ȥg��i5��}�=9p�>qj?�P
?��ϼ�����5>�t?t#
����dr ��c?�	@��@��Z?�Ϡ��.�I�����������>\�> ]>s�ѽ{�w=I�)����ȭ��Y�=ڌ�>���>^��>j'3>�>��>�[����%������t������R5�]���C���V辈Ħ��{侏l��I	�^��<�}��cڽ�o��� �t˽N>�NQ?j`\?��q?'��>4 ɼ���=(��:_0=)y����=tS�>�p7?�LJ?aL0?8��= p���Ga�X������X2���)�>NWc>���>���>-��>Cm�<��#>��>��|>�>4'�t>�<���<�� >f�>�d�>i��>��7>��>���.��:�i�	C~��Ƚ�e�?s7���VJ��e�������ڹ��=��-?˪>=ꑿ;пk᭿�bG?&��������3�\�>�I/?��V?��&>����RZ�GZ> ]�odg��f >�����o���*�uX>E?��>9��>��R�E��a1�B����le>�A8?�����M�LL��:�G��T�����>�?���<A;"�͜��^M|�S�s����=�B?V��>K8i������2w�@����D>�4o>��<b�>;+8>Z��ý��f�\����)>��n>w=?� >�	>Xa�>�h�������>�f>���=g;?h�?��ƽd!�=n+c�]~3�ȃ&>;��>9�N>)�D>��q��Y�='�?֓>����K�w��	�'j���=>y�����U�t떽�Z�=�6#�%U�=�!4>��㽟�^����~?���(䈿��e���lD?S+?f �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��G��=}�>
׫>�ξ�L��?��Ž6Ǣ�Ȕ	�-)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ<�>e�U���b�����c���
�8B�>?N?����a�&VT�^�?���>���Vk���̿I}��a�>���?[�?�6r�t�����.��� ?���?9�S?�zJ>�����%��9l>�=H?ܳA?��9>܆;��J�E�?Xܱ?�V�?yI>���?a�s?$�>,wz��R/�YU��{���Ci�=n��;���>@>���;F� ����1����j����˨`>;$=*/�>����Q����=q8��?�����g���>Whs>VzJ>	d�>q?���>�ә>�~=�|��/؀�v��K�B?�?6B�Ds�[�F==LV7���?!�7?�X��A��8\>�{H? ��?�h?��>��m���~Ϲ�T��O!=_i�>���>ˤ>a�ѽ�$;>4���T��0�>b�m>���<Ì��ٙY��A�?B�>�M?�3�>x�=;U?$&?X�9>�c>ƺ;��F��j~����>[4�>���>��X?UH?e��~O(��x��銖�LTE���>+hu?9_$?�X>�_�� ����=Wͱ�N>bI�?�+.?hK�r%?0cd?2�c?���?3��>-������c�(����>��?�q=̀6�k~Q�*����>@+�>���>�H��_�;����ʔ:�j�о_�?2�s?MD
?m�;~���5��g�<�q1=h�>ҫ�ń>ߝS>�h�=𕵽@;o>�=�F���M=�n<^��@k=�/>�н>)8�=y2|�S�S�E�?�O<Lϒ����<��_���E��h�>2=>��-�6?)�3��T�j�� ���5,���?�+�?*��?sh���s��*?���?�?�� ?�)�����\���4K�~q�'�����˾�>6�<�x������w���wv�����D�!��>=?F]?��>�H�>zB�>����D�%��>���<�Y�������0� �0��Q	�hP;��V�=���=�(��!���K��>®\��=�>�2?��>�Tx>�z�>���ʘ�=�l8>��>�%�>	Q>HAA>}Υ=č>�v�i�p�P?���\!'��E뾪��� J<?0d?P!�>ꝅ�e`�������?��?-�?�z>��h���*�%� ?j�>�~��?��q=,=�����p���*�����O��~�>�_���>��I��Ya�X;?��?��?߾	�����]�o=.I�?I�(?��)���Q�B�o�R�W��	S����FJh�_W��G�$�`�p������Z���!��i�(��{*=��*?m�?W�������*k�?�u�f>���>��>���>��I>��	�W�1�0 ^�S'��ă��u�>]{?^q�>A
.?UJU?3�r?��S?�=�>G�q>�4�����>v�>��>N�>/6?�:&?�'?($?71?��>��8������%�,?��?X??o?�%?�^���p��U�=���<��J�x=�e�=�t��9�*f�ڲ�=�C�>�n1?�H�A�'�2Ϸ�?��>u��>{C?�dV?�颾�7���y>��>&�;?Q�>�C���O�����Z0?#�?43���6��:>�f+>�-����>j��=�G۽��H����=�	������K>���7�D��Y��=`�ѽ��=�"�>&�?�d�>c�T>F���������~�=H}�=�>��<z�������x���i���>Rz�?��?X>Ua>y�7>U2;�nپ����m�g�=�_1?O"?@�Q?��?�D?$*-?�wa>����\,��r�{��0����?�+?�`�>VZ���ɾ<w��c�2�t�?�E?�`��4�*�(��5þ��ǽ1>�e.��^}��H��X�C��C�������R��?���?)J��@6��辍��$��Z�B?3��>�>��>I)�)g����9>��>�`P?���>��Z?&0�?�oj?7�=���4����ð�̚=
7�>7�`?��h?]~�?� b?=~�>p��>@~������"��ą�\O-�����-���9��>�>�y?[�>twa=��r��J=��f1�<
�=�>� ?rŤ>	g�>,f+>����T?p��>V��*���d�i���v�,Ⓘ�qR?��?��g?b�n�YjB�I�(�\�ھ�!�>�S�?��?V�?�ž*m�=g7�k������b~>s%�>H�>*��=�>�<
?>���>���>Z�s��h�ɀ,��N�<�6�>�0?��>X�׿IW��G�r�����>���t澘�@�p-����нU;K>�[R��x���"��x�E�O��N��+ԾDģ�H�&?��)>�a��H�> Cu�s�黚�>������
��ͽk�>��ǽ%(;l�=���um�<�T�=�<$ߡ�?�ʾ��|?��I?��+?��A?� }>fB>�I>�罕>����V�?�S>u)F�ƺ�L�<����ⴕ��;׾��վD�d������>�M���>o�9>1�=ӥ�<!�=�@^=�=2���|�=�=T�=;1�=���=�>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>Ck9>.	>�R���2�q�Z���_��<X��y!?��9�^�̾�X�>B��=>=޾��þ��M=4[5>wTG=�����[�
�=�u�^�H=Lrf=C��><�F>�Թ=B)��=��A=9G�=��N>��ƻ 0����#qE=�U�=j�]>>�!>�<?G�?�F?��~?r�?W޽�������޿	??^�>/��=
۔�Bh�>�J�>��<?M�W?��Q?+1>�w@�$��>�p�>0�O����||ƾi���4&���y�? ��?���>�P�ρԾ�D(�8+9�Z�>�d3?M;m?���>���'W���� `&�ҋ.�#�����7��)=m}r���U� �`��#�㽬��=4{�>��>��>Iy>6�9>{�N>4�>��>���<Ѕ=Fđ�:��<���聄=`꒼���<�?ü|阺��!�ߜ+�Ш�ϋ;w�;�g\<Z��;N}�='v�>�4>[�>֕=�t����;>H���~J�}��5����8�ʡb�1����3�)<#��	�>��>p���K���L�>X}�>��>t�?�0�?A��=#�t��G��◜���d��͹��3>b];>X���AH�|h�2�>�J������>��>靰>mt>�8�л7���=c޾�*3���>zs���SK��ǽ��h�㦡���a�eƽ��A?w����0�=��?̹L?�?���>l�~�����;>�ꖾ̏=o#�X{�������?�$!?zW�>��ھHMD��Y̾� ��<�>؉H���O�U��� 0�:'�����F�>	[��AdоtT3�#�������H�A��o�I�>ԚO?U��?`�7��8mO�/E�I���?��g?�à>]?��?㥙�C?�ƹ��pn�=��n?�H�?oz�?��>;A�=��D��?s�!?���?Lթ?G�s?[��VU�>���=ο)>�u%��g|>I5�=oQ�<p��=dN ?B�>��?�Ԑ���+��b��k���偽�d�=�w����L>gx�>S7�>/)g>r�=��l�= k�>�o�>��\>�>��>G%����	��.0?�d8>�$�>�MX?���>ZY�/BR��5=�W\�w�c���J�񗽬/�D�4<4�;G����<���>��ĿkƁ?g�k>����?%� �����x>)��>� �D$�>D�=�H>I,�>�>�7&>,�r>�L)>4�þQ]�>���afE���`�ڈ�����[�>�gj��ju�M��PwT�]����,8�p���bf�����G)�$C��sZj?�%����P���$��y&>ORj>��s>5'\?����󽋾���>ݡ$?v�>i�㾵(�� ����̨�?��?N�?>37�>��S?&�?j�B������L��rm��cF���b���]�0H��Aw��F�ӭ���X?w�z?>�F? �C=���>�X|?XX����NoD>I�6��c)�
/�=�7�>�����m�(���̝���^T� �6>�Gq?�\~?k�?/65��$��D�>��N?�rQ?��q?6=?�#?����?���>%?�?
?1�<?4?��?�D>;��=�����я��7h��%��Z ��'���<��/=��.=/!�<C�l<q�=pܛ��ݜ�O�m��������O�R<�\�=��U=��>\� ?�PJ?�@�>��>�.?�W�� �f��ݘ�Z�?E� ?��Ҿ;,�'a��/�پ��>�l�?r��?��8?o���
�_�6
����^>�,
? ��>#w�>�V�>;;?����pH��:�>��>"FƼ�˔�I�w��pھ͌���A�=���>k�>�З>8'�<�+ >�Y辯Ss��:\>4-�h��Ub���D�kq(��
��ۿ>�ZG?�?�T�;�\��w���[���?Id=?F�I?� f?�g�<ƒھD L��G�1A>���>W�>7�����`���J�l缽��>��`��U��N@e>�����޾):n��xG�q��7`J=����E=�_�˾;m���=��>��ľ;S!��V��v��H?V�r=S[��jZ��D���`>�x�>�]�>�@ѼT�����A�G&����=���>Z@>
���#��$�C�����`z�>�E?�a?Tt�?���1Xq�n�C�*���s��Ħ�o�?ޯ>sK	?1�H>m��=蹰����)d�&OG���>�L�>��:D�����	�����%�О�>��?�D$>n?��Q?�#?�B_?�)?И?W��>�9��}V��/�2?Pp�?)	�=Yw��+�#���7��jR��F�>-<?�Pٽr�w>�W�>]�?�!?ژ\?��?�H>�辠�C�SJ�>���>/}Y�����o>B�G?l�>�1P?��?n�T>�C:�+E���˽��L�=f�>Q�1?�I$?s�?��>x��>p���f$�=ƨ�>�c?�1�?��o?�U�=��?@2>��>��=��>g��>}?nWO?��s?��J?���>S��<�/��a;��OEs��EO�p��;�7H<��y=���,t�MH���<3�;�ⷼ�a�����ӲD��萼F��;���>��Y>X6����D>�2Ѿ2����L>��Y�)���u���2����=��>�?�>U�J��< =��>���>ҡ��2&?�?�~?ǫ�;8f�>��4ё�o��>\�=?�.�=��i�2���l��ר<��s?MjV?!j���C	�(�@?��e?�"���Q���ȾA�T��\k��4^?|?�>�o��V�k>=�t?�Ub?4x?�uZ�_�s��u����S��G$��E>�D�>(@��PX�M܆>�&?#̞>6r�> �:>֖��8zo�P,�P��>���?��?]�?��C>�ы���ῳ��� ,���^?���>w����"?B%�͛Ͼ{Y���u���ᾃ����몾����}���`%�������ֽ���=�y?P�r?L�q?Q�_?'e ��c�4*^��)����U��������E��D��oC���n�C��U���2k���=@=u�ʣ\�	z�?~�1?��S�V?&�R��������J,{> �u��0��>�s	�w�=��K=$@}�r>3�E̕���?��>1��>O#0?kf�t�4��?�%�,�y���\>S~>&h�>H	?��L;��F���ؽA���s}�����&v>�tc?̘K?>�n?^w��1������!���/�CX����B>�r>�ŉ>̀W�j��}2&��T>���r�B��ct����	���~=��2?�D�>~>�H�?��?w	��J��Ex�3t1�⇂<P,�>zi?z/�>��>��Ͻ�� ����>��l?���>��>���rZ!���{���ʽ$&�>�>���>��o>�,��#\��j��O����9��u�=$�h?���(�`���>�R?O �:��G<�|�>��v��!�|����'�!�>Z|?���=�;>�ž�$�|�{��7���v+?�?� ���4&����>�#?M�>�4�>��?_͟>�z¾���?��\?��I?��B?��>m�*=�����˽p�*�* 8=«�>�&c>Mj{=���=�j��'d�$�%��&W=���=��Ӽ���bٝ;�X����^<�c�<��8>��ٿ��<�SGѾe������������ʽ�ˊ����ه��<������8Zl����v;A�Y�/�(l��w�]��8�?��?򧆾�i����m3���+���V�>��$�
�¼���T����3i�D4ؾ������$��0Y�g�P�T�ҷ&?���Ѯ��Ϟ����mw?�_?k#y?5q�x��N�5�,B7>�f=�7B�M!����>˿󂓾��_?k�>�|��&ؽ��>tؐ>�`y>�H�>�|�ӯ��$[���%	?D)-?&"�>@g�6�ƿo����d�<�M�?��@��A?��(����TX=��>�	?
y?>)�1� *��ذ��R�>�4�?���?�#N=��W����tue?to<[�F���޻H��=�y�=��=߉�ClJ>�_�>f_�/�A�g�ܽ��4>U�>�H#���Xe^�j��<�k]>��ս����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�}��=[��>c�>,������O��I��U��=C���؟��:�o(��B	=b)��}�<��u�"B��y@��(_�*�9��A־%ޗ�q��~�>Y��>���>p-C>ø3?�g?No�>z�y>�0]�&�2���ƾ��M��y��򴽅�=�qƌ=罾�BM��� �Y������:.�����F�+>p�A�6]���"�-�q�d�:�_k ?{�>먪�o[5����=A)پ5���A"��L���]����"�A�S�ǰ�?N�<?h}�� N��]�}`��Y{�Y=[?�lc�����|Ⱦ)�7>L{�=�>���>٢���U�js3���,��u0?>Z?_����[��1 *>�� ���=�+?��?ڂZ<%�>K%?��*�C)��][>�3>Lң>���>�F	>;���P۽�?��T?��] ���֐>ch����z��5a=u,>z;5�C��`�[>�I�<�팾>�U��[��\�<�R?Y�>�/(�JW��Q���[��v?=�v?��?L&�>�yh?OE?o��<���X�T�E���W=q�T?Ki?r >pf���Hվ�Ҩ��4?��f?��`>��X����-1�����A?�Ar?�D$?�J8�+���m��E���;8?91?C'a��a��@j$�?���45>�z?
��>�aO�$ޱ><g?q�q�v���ÿ��1�M)�?�q	@a��?$=NW|�J��>�?o�B>ޛ��;Yԕ�������=R�	?(Ý��n�j� �뙵�t�J?��s?��>v9t�KN����=ܕ��Z�?��?����a�g<H���l��m��A��<�ҫ=?��7"����(�7���ƾf�
������ܿ���>�Y@Q轝)�>
E8��5��SϿ����[оeSq�k�?��>6�Ƚ������j�dOu�j�G�]�H������f�>�.>_ؽH��[�t�jS7���=t��>Zd���V>�DT�T����[�<��{>|o�>�p;>����+��k��?3�޾��˿By�����F�]?��?3݅?�?4+������ݿ��AaM=O�h?5��?�??�u���Ml�����e?�¯�4H�����E�Nf>��7?���>��,�e��=v�>���>�Z>�x��������ݻ���?�?_�޾E@�>⚟?��8?�i���=Ӿ#�@��2=2L?��=Aʾi<�n�*�@*��.b?,?��P��,�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�
i	>���?�~�?Qj?���� ����U>
�}?2	�>�}�?���=���>?��=������8">pG�=�)��e?2�J?69�>�9�=��=��^/�3�E�3|P������C��P�>X�d?��M?�zd>6�Ƚ4�K�޹$�=���{.����D���7��5�M�*>,�G>��>�K���׾I�>>kO��+ٿ����Ʃ�?��>R?	f�|Fɾ\+�=�
�?V}>�H(�y��S�n��T��ڤ?��?��?Q���Z���]p��?s>ȫd>-ο�j�8�����
>g�?�b>�Z���q��j�]>�x�?_6�?3��?B{n���>�u0�
���Is�Z�Ծ�C��D��=Z�"?QO��׺=��?�g>���A��[ƅ�ۂ�>p��?3�?�I�>�7a?Fb(���0�=��'�>�rJ?��9?���d!�-�>Q�$?��9� ���f���*i?��@�@��l?����ҍ���+�������S�H�>٩<��6>�^n�e��=�;=>H>��>A��=�Ē>P$.��#+>ժO>��b>�ϴ>�V�d;�ݾ��(���$(�m�B���:�e=s�����)ն��=�$�ӾI�g�ڊžl�,��J�<w��g>��=~�I?f�Q?��b?���>ɧ����>v�m����� ��|�=]�>˝,?	U>?�=?��'=����X6k������J���͢���>d�g>d��>H<�>�(�>�ҋ��'>�-�>9xd>�h:>��=~я�xw�[��=| �>�Q�>HO�>�7;>�>˅���&���!h��lv��nŽ�?#����K�������D���=�/?M�>����/п`}��6~G?�[���"��(��S>�z0?a[U?�F>����sX��4>s���6k�*� >س�� mc�o>(�� F>��?�G>M��>�>���7�<�X����
a�=K�F? $�U�ξyw��~S�L�&�F�>]�6?�9}=�)��ɬ��e���)���'=Ø@?x��>� ���˾�^���æ��&>嚞>/	�;>b="A>�����F��`T��N>1[>M��=R`?-_)>*��=���>ӛ��Q�l��>��B>))>��??�e$?�n��ً�콁��/��iq>���>�W�>�5
>�LL�́�=֘�>~�f>�3�z��ߔ���G�q�Y>�"t�q&a�>�5�w=������=.�=�����?�p;=�~?���&䈿��9e���lD?R+?~ �=U�F<��"�C ���H��E�?p�@m�?��	��V�>�?�@�?��>��=}�>׫>�ξ�L��?��Ž/Ǣ�˔	�)#�hS�?��?��/�Zʋ�=l�|6>�^%?�Ӿ<�>F���6�J0����n�HI���> ??E������n4�oA)?�l�>d��G��~�¿��u�;�>��?5��?�R�`:���C����>[j�?�s?2h�>�p�u����0>��-?��j?�|/?����혵���>�1�?o�{?3I>���?Z�s?H��>:�w�ZP/�4��1����I==_d;�q�>ֻ>����5=F��̓��[�� �j���(va>}%=��>�C佦���02�=�^��gh��S]f�/��>�}q>�I>�]�>h� ?/b�>���>vK=�r��V���(�����B?�Ə?Q�	�4�j�{)�8�=��d��<?�2?iV�������>�GY?�?��b?a�>�$�v𜿨$��:尾tX�<Et^>���>%��>�D��r�G>9U޾�$p�~�>�:�>?{̼�澐�����.��Q�>4S"?���>tz|=��?��#?k�i>?�>�dE��J��$�E����>��>�%?<g~?Zp?Ƒ����3�p��'����e[�Z�M>��x?a�?at�>����}a��}+A��?�J|��њ�?̲f?�E��O?�?k6@?��B?��g>���]ھ�ƭ�^ׁ>m�?]<\C��5���"�/��>i{?q-	?jg�a���ڍ�t���̾ �?Jx?�e?0m�@�P!پM.�<�,�>�X=�(�=��8>��B<��˽�P>�"%>;��;� �A�LJڹ=��=f��>�]>\�������>ޝ#��	þH��LH�N[����>��;>i����yK?J���cu�H���ȟ�?�w?qL�?g��?ƫѽJ�e���6?A�?w[?��>ٿ��ؾ3%㾚Od�$�t�$�Z�>�x�>Ձ<=�պ�:퟿ػ��̇�C׽�~#��0�>
"�>z�?���>SӚ>���>�u̾&&�����	���Z��G�A�"���7��/�����)��~�<.����&����i>ķ���j�>\49?�\�>yE`>���>Tx��s^Y>:�R>�f!>���>=�>��>@�=�S_=��½��N?�a��"(���㲲�O>?k�e?Q��>����\��4��,&?�?Vݛ?��>�h���-�r� ?��>��v�N�	?׽\=�3�
�2<򓴾T
(�go���Z��7ȉ>d-�'�<�HJ��]�@?��?$�y��{ྍ�������_=���?x� ?:q-�ܚO��~l��S���P���<���y�������Ĩj�Y^���T��񀿍�)��Z<TL*?���?������������k�eR=�Y=�>$�>��~>*-�>R�T>����o0(�^yS��*��S���T�>]~?}V�>�p7?��4?2Lc?�_v?���>e�[>��ξG;?�G�<*�>�?�>��3?A�&?Ξ)?)K"?��*?�_X>bY�����9�~?�%?`�?w4�>`�	?.$���:�_'��'�l<����jѽ��=_�.=K���ŵ��1kl<1pz>��?��k��Q��ܾ��g=V�.?�?Vh#?R��yoþc�>�
?C'?AQ�>\H�|d��"��j�>k��?��ѻ/��<3>k�>�g�=.=�4z>#};-+=� ��n�=!U���>&=���=J��eB��$;x =�>)�>��?��>�>K���� ����H(�=��X>:0S>K>_پr}��L2����g��by>Ov�?:o�?�f=���=�=�e���N��k���� <�<��?}]#?�WT?K��?(�=?^|#?f�>o)�dM��&i��"��V�?�~+?�ۑ>�9�P\ʾ5���8]3��/?��?�	a�����(���¾��ҽ�>T�.���}����l|D�D����������dd�?V��?��=�E�5���o��G��A	D?�"�>⁦>Hi�>��)�C+h�U�F�;>�3�>��Q?�6�>]�m?�ϔ?jC�?�˹>�>��4��ಿF�<�=�>k�L?Q�?j�?���?B"�>{�R>��p���f��'��<tU��a�U�->/�>{�>�ߎ>�7Z>W4
>|F$=����Q�1�H$3>y��>r��>�>_�C>Ofѽl�b?f`?6E���t��|4�Asr�%�[�G$e?���?�M?�\���>���7�D�޾�� ?>,�?��?P-?�$���J�=&=���N���L��>0��>r,�>d���5�=V�$>�Ը>��>�	�ڒ�T�D�s*<Cl?Dq<?�D>}��\�^��!�����u恽�Ӕ���b�+"�Q���%>���2���w��Z^q��K��@ؖ�(����L��L���e�>1zj=��%>�>�=y>+=�.�9=�m�=dui=�� =u+�`�=�'7<�,Ӽ��觽F�L�Wo�=�"�=�e̾kax?��I?dT)? ,;?e�t>�>�>����>dh8��?��V>@�0�R(��2%:�3"�������߾.U޾��]��C���u>~d@�o�>��->���=�t�<a�=���=Q�Z=�-<
?4=D3�=��=�k�=F/�=>�>�6w?X�������4Q��Z罤�:?�8�>e{�=��ƾq@?��>>�2������zb��-?���?�T�??�?@ti��d�>K���㎽�q�=M����=2>n��=w�2�T��>��J>���K��B����4�?��@��??�ዿТϿ3a/>��
>�z�=%�Q���3��%Y���}���I��w?9�>�5]ʾ/�>�Q�=*���Ѿ,�=p�E>s��=���!�V��f�=�b��K�=� �='�>"�R>B�=TܽqI�=d =�:�=.QY>_��<��L�����ܹ�<X��=��6>b!->��?���>I=L?��?�`�>G��DY���оY��>��>�j�><����L>�k�>��@?}�<?�t*?�
�>0�ɽ��?�#?oaC��r��-o����3��Q+�?�U�?��>�ii����=�?�VQ��M�=4�?��?7-)?&Z>�U�m��,Y&���.������$E�f+=jnr��XU�E����k�����	�=so�>���>�>VUy>��9>��N>L�>T�>�>�<�r�=
ጻ�ʵ<���j��=������<�pż:��^&���+����l��;���;�]<���;k�=~c�>�N>w��>�#�=�����/>3Ė���L����=x����B���d��V~��.�-�4�ĻC>,cY>�?��|����?��Z>��@>40�? @u?� >�c� �վ�A��nd��WR��κ=�>b�=���;��V`�M)N�6�Ѿ���>��>�ۧ>�z>sQ-�@�>��Ȃ=�RܾhE3���>�\���<���i��z��������f�u",��E?����:��=��?~+M?�?���>8�����(�<>�{�$�<yr�|s��'���h?1�*?���>N��7H�{L̾"���ط>�DI�~�O�4�[�0����η�@��>g�����о�$3�ah�������B��Cr����>{�O?��?0b��V���TO����0���q?�zg?��>|K???�*���z�=t��^u�=��n?h��?<�?� >;�~=�K;���?��?
Ǉ?�I�?T�?�����a�>d���R�q=f��� >Фj>���<j�!<R��>6Y�>۹
?}�]�'�$��R�C4Ѿ��M����=A!<>K|�>*=�>�%�>x�z>�`P=�N<=w�u>j��>�ך>ڕG>剒>�Na>�:��[�(���,?}�e>�v>o�K?~��>/2=�y�3����=�-<��r�S���Ve��g(ǽ-�;Xɚ����<�<��>�zȿƔ�?��V>��(�r��>C���%���0>b��>mqx�6��>.=�>L�;>���>�<�>�'>Q/]>4��=�S��蠷=P���4����[���I�O�߾��>ϸ����۽�� ����<�л)D~�������z�r�z�&+�U�=��?B;��ry��o)���(�n?��>�GD?�2w�Ťͽ@�2>5��>8��>Q����h�;���ə����?"��?zBc>��>o�W?�?f�1�<3��vZ���u��%A�=e�ʺ`��፿h����
�:����_?�x?{xA?�0�<�?z>��?��%�g׏�p*�>9 /��(;��e<=�1�>�'����`�ĲӾ��þ�:�WOF>g�o?�$�?�Z?6WV��ck�B�#>)�:?�2?5t?F3?:T<?���hi$?�0>u}??�
?��4?%/?�^
?_>0>rv�=ns����,=�ᐽ#n��Q�Խ��Ƚi(���4=*�=Ŕ�:�o<�A=���<f��r���N;9��� U�<��9==o�=���=F+*?-U?R��>l��>Q~�?�x>�a��m��؇?�g�>��y�P+��F�^���NL>yJ�?��?�bH?��n=G�J����[>��?�?���>�K�>����V̾�a��%�>$��><�K>��<�ӫ���Ҿ5�t������q>f��>�A�>0,��O�=�M�x���̢;>��A�����z��A;�H�2�G�I����> �F?��?�$9=&V���g�|�a����>)�@?B:R?y�e?Vy
>Vخ���a�k����N��>�9>�l�X7���b��
?�^w=�r>�k�c����|>����� �����zQ���˾w`>6"�d���aE$����9F��R>.�=Nɧ��Z��W��֟��>?2R> �a��HD�.������=iK�>%*�>�᤽?F�8BF�(Oʾ]%�>d�>��`>��;.E��t^�$���V�>ŠE?�o?v�?�D`��Eo�:�`�������Vu=��?���>�7?rs��4=t'������a���0�\K�>�?��{�I�����D	�V)<�(xL>B?�KN>4?��]?�:+?%z?�� ?C?�,}>w"��<zž�',?܂?._>��ᓷ���8���H��/?!US?im�S��=��>��?��?�KU?9I?�3?>�R�cSC�0�>�]�>��d�A�����>f�;?6{�>�']?Y��?v��=�KG�9����>���<{���>ʜ?��?7�#?]��>��>r�׸>��>n��>o�?�+�?/k��dK�>��B?S`�>�)<҆0>��B>��?,Yl?��?8l|?�?1��۽���Tq��P��I�V=(�}>��[=kQ���=G�k9r&R;
T�=��\=|E=����*�����=�1=��>>�{>~����/>�Tо����H>�	��Ꟑ�@^���IU���=k�>#=�>7�>}<&��΃=r�>߁�>����#?m?1]?]��zZ��Gо}p�2k�>��C?W��=@%q�>u��Ur��r�<�n?��Y?�4r����ay_?�h`?NU��@���̾s�t���� U?�?��k��a�>Yx?M�n?u�?9B�A�g��H��cSe�S�|�H�=#��>��\�lT�>	e-?���>w��>p��=��۾jn��٧��_	?,��?г?�;�?5bt>YLu����x'��Wݐ��_?n(�>%N��~�$?,�;��Ӿ�+��x;���྾L��|Z��b󟾬w��2!�Qǂ��aݽ��=�R?/o?~r?��^?o���_|d�f!_���|�)�W��, �����pB�J�D�q�F�1�h�zS�־��DE���`=�]h�Z@��*�?:?��pf?�T�f(�G����d>?O���< ��:�<S�d�*"컴xm=	�U���:�����D?��>_y�>�1?��G���O�ѳA��!����x�E>78�>�a�>��>6���km�G�ŉɾ��y�ө����y>��b?c)N?�ro?����T-��u����$��k6��a��L�B>�>-�>��b�HP�=
!��:��_s�[���ӎ��n
��w=J�1?-/�>5��>�B�?́?m�������|���1�Z���`\�>؟h?$R�>�΅>K�ٽ����>�Ki?�H�>��>֊��d��	�w�;�;��>�a�>ײ�>Ԕ=>I�<���U�"~�� �T�;��n>Gpk?���	�`��Ԓ>�U?Y>%�̕�<��>M���!�8�����5�V�=�?�wE=�JE>w�Ǿ	6
��oz�����j�(?/`?z����)���a>�y?���>涬>�?=s�>T�Ͼ$&��?7�]?ٻK?�*>?���>�O�;X8ݽ�R����!�ڶ=·�>o2i>L��=F�=����~]�ei"���K=�	�=콒��(��/����A&���b9e�7=�_<>�࿀Z��]�f�ƻξ^��l��~G��Q����;�;2����������ؽvt_��Q���{������z�p��?j�?�`���������F�y��w�\�>�����
�G�� @�ɮ��վ�����Z"�׬Y�Z�i�o�f�Ц?ƬY=�+���n ���Y�=ZH?���?2����n��KN����><">�O�>��M���'ƿ{�!�epB?΋�>���y���>??��><�>R2���+��o>�If?�s<?��>����Oɿ�@��=]�?-	@�eC?�!�� ���=�T?Ho?���=��T��`����>���?y��?9��<�lR��P;�f?���<l�=��#ɼ��=o�>=,�=d
��\1>���>�<2�����Z+���o>Wf�>f�н=���n0�yst��,L>��������Ԅ?Hx\��f�V�/�zU��'N>��T?�,�>�?�=U�,?�8H��|Ͽ̭\��(a?R0�?U��?l�(? ῾�Ӛ>u�ܾ�M? E6?��>me&��t���=H���k�����9'V���=ȩ�>��>�~,�ϊ��O��B�����=_�$߿X~E��K�tR�>�-K<|!�<ֽ���8�����1R�<r�-�$#��~:N>|�w> �B>�L;t>�k�=Ӂ?�y�?p�.�W�3=Ƽ��#$��m�Ͼ�����]���}��/���$��eyϾ�v�����Ƶ�U5>��],����6�7��I�=�G�1����45�:�u��7 �˽7?~��=�� ���K��6=c+�5���)��/0��8ξ؈���Q�eP�?]G?��R���9�)��>�}��`%��qe?6)�����F��!�=��	>2">���>�Sj>�OӾ��[���]�T�8?�S?9���Ve��^�B>��(���3>�2*?�P�>�_9��'a>�xI?�6c�(f)���>A�����=q�>�>�W��j�׽�Z;?fr@?��ž��q�
�7>�6���]��e�=S����Δ��YW>\�=׾¼A�����d=�2�0ν~~V? E�><B*�q��9��t���F=OVx?��?Z�>��j?=C?_��<h
���U����߬q=M�W?�j?��>�Iw�8-ξ�橾!�4?�e?M�I>�l���".�?��܁??�l?m�?����-}�������W�5?��v?s^�is�����0�V��=�>\�>���>��9��k�>�>?�#��G������mY4�#Þ?��@���?T�;<��a��=�;?f\�>�O��>ƾ�z��������q=�"�>���wev����<R,�T�8?Ѡ�?w��>���������=����C�?6�?�H���@=����0}�~���	>�
&>-r�<R,ƽ�]�P� �O$��b �S)��y�<�F�>�@��<퓰>R����꿼��1����}��i/X� .?�p?w:>�P���(6�Z:���9�V�A��Ս��ė>��>O=��ȾE�{���8���g�?���U�=�<��t����T�_ě>��>��>k�6�hY����?~����̿�����	?��?��?_�.?؝Z�B�N�<�����=Tr?M3�?,��?ZF>&o�gX��#9D?�`�b�Y�R�R��|�ی�>8?M��>L�;�>�r�^=>=��>]>���x̿�.���=�DI�?���?3����W�>:I�?!��>�c�G�}�$��$*N�G��=Z~?�J�=�j��fD����-��@E�>��>+�6��(�з_?'�a�G�p�B�-�"�ƽ�ס>X�0�l]\��)�����Ze����'>y�P��?�]�?��?r��z#��3%?b�>����7ǾM��<i��>Z*�>8,N>�H_�~�u>�	��:��l	>z��?�}�?�h?�������qZ> �}?�P�>[��?W,�=i)�>���= ��|=�-�%> ��=-F��?%M?��>x�=IE5�z�.���E�F�P�9��'7C��ˇ>F c?�YM?YZZ>������0�d�!���ͽ�,�������F����Cm���/>�A>`t>� I� �Ѿc�?:��ؿ^0���l��eQ?f?�>e�?�k�(����@=X]??.�>��R����e��D��ܬ?���?ym ?�s�s�$�E#>�ɽ>r��>��q���s���Ẅ>3yB?9�k�sy���Vm�ł,>*��?��@u�?\T��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?SQo���i�B>��?"������L��f?�
@u@a�^?*�+�պ�:���T��h�>P�S>
a�>�Ͻ��<=��=i��<�ڽO��<�l�>x��>��K>�?S>NK>|x_>ҋ��UX-�����荿�}#��J��$��F]���lş����<���L��l�;�Q�=t�o��g�r�n���<�$�=��P?/jU?��t?�A ?sF`��>,I��=;���ȼ=ˤ�>/�2?�<P?�,?�M�=�O��>�a��A���料|c��-l�>KT>�+�>���>�g�>�gr���<>��N>���>4%�= FK=�|�<z��<�<>"l�>���>��>��	>b�>� �����pt��C�/ur��%�?�l��W�U�+����a��v茾a~q>�* ?���=�3����ǿ>���*�??�3��*����S<>63?n	h?K�>>)Ŵ��$R�	��=�8I;�����>�%��ാ��:��÷>�?��>"�>���H}��Gt�����<�8I?1������Ey�#KS�9ރ�5�>a6?�[�>b:������ڔ����Ξ�<�P(?Z�>�M��u�-�;��r�D�>�L�=� ^�KW�x�A>Y0+=鵰�h�X�(���� >��>_v?�">T��=Y��>%Lq�ڀ���>�>;B>�s;?�[%?r������R
��&$�-g�>u�>z��>��>ŅO�6��=1y?�]g>���k㯽cpŽi�$��cf>��߼5e��۽��<�"��JN�=WM�=�a`��)��sE=�~?���%䈿���d���lD?U+?� �=�F<��"�C ��|H��@�?p�@m�?��	�ޢV�?�?�@�?��
��=�|�>׫>�ξ��L��?-�Ž3Ǣ���	� )#�fS�?��?��/�Zʋ�6l��6>�^%?�Ӿm,�>�<�����o���[o���<4�>J?H�������<4��?�:?�������ɿ�Ix�B��>�g�?���?@um�����68���>���?��S?��W>M6ݾ��8�nĘ>�Y;?�O?�ͩ>�l�@�2�gV??���?��M>*��?�D{?�?�>cr��3�����!���wh�=:B=���>��b>Ab��M����lI��y�d�?>�Ǻ[>nA>=C��>Jֽ1�̾*�[=�d��@ᴾh�?��>���>N>1ۢ>Ģ?���>q��>ɚG=]��x�h�Y	��!�C?��?���֌g��F��i����l?Ti?B��|۾vit>�~??�y? Ll?V0�>����%���ÿ-���tO�<��=�q?�1�>ȁW�Z�8>�UѾ�c;�2_v>#��>Y�7�.v��l���c�<���>]\2?<p�>�����E?�m#?��p>j�>f�C��i����@��|�>�p�>*2??�u?�\?M$���:�8����<]�)�G>�u?=� ?V �>�(���d��8�^�ڽW<��췇?b�i?r����?�Ј?�??��E?���>T׍�o�Ͼ��U�X>�&?3�弻�4��#�(�I��0�>B��>	V�>�4��=��;1v�qE%�"�۾(5
?��h? /&?n Ͼ;�y����<Տ���<�<�O�;�t��,>���=]��[�=��]>�=�]�7��RI�'M>=zU�>���==~3��=� =,?%�G�Sۃ���=t�r�xD�A�>sIL>�����^?jl=���{�����x��	U�� �?��?]k�?e���h��$=?�?D	?k"�>�J���}޾.��uPw�"~x��w�+�>���>-�l���A���љ���F����Žb����>��>��(?���>���>�s�>g��mL$���ʾֆ��li�l?.�}�s�woB�^����վy����=�l����t�?k>�������>(�?�&h>�y>�Q�>�׽u��=�P�>���>	LS>�P>T��>�v>���fX[�U�Q?��'����L��E�??AWd?��>=cl��E��`����!?\��?z��?D
s>�h���*��?>��>}�y�G�?��=R��;��<������H��X�
��4�>����H7�S$J��Qi���?i?�ED��HǾ��������2o=�I�?��(?��)���Q��o��W�	S�^w�.Ih�W_����$�įp�ꏿ�b���$���(���*=��*?W�?�����`1���8k�]?� �f>
�>C��>�Ѿ>j�I>/�	�`�1���]��'����7�>�9{?���>��.?�3?o?W?~�g?�͹>�B=>͙ξ��>_�=�1�>���>��1?��?�?��?K2?k�a>�Iｙ~����ݾ$�.?r�?���>�q�>_{?؞b��Q��[�<X�1=�ي��+�d�=[Y=h�׽�^�<h�"=�t]>��>-�ݽ� k���׾N?u0�>�?�y?5!�5���>���>�l?'��L�w�����
���.A?�d�?΋,�e������>Dx�=� |��X>�.ս����A�=,�&�\k�<K/=����,Q���n�=^|�=y+�=]z@�n�a��t�>��?���>(D�>D@��˩ �!��d�=�Y>�S>_>�Eپ�}���$��Y�g�^y>�w�?�z�?Լf=o�=���=�|��\U�����d������<ף?�I#?XT?T��?n�=?'j#?�>�*�^M���^��~����?L�)?�͔>
j�&=ɾ�����d-�0�?dg?r�Z����ĕ)��ž$`����>�,�9F�|A��~�9�[��;o<�%���g��?��?����0���޾bc����F?aC�>ՙ�>L��>�i(�BKe�
�N�(>��>\�K?$��>��2?��?��?XH=>ytվ���%ީ���<%��>(L?�7�?	�?�v0?�b�>��>'��i����$�y�x�0笾%��[E>q�>���>͟?3�>.r<D�ڽ��<�?�����v1�>}B�>��*>�>�lZ>�v��ZC\?�<?(-���+�
G��yQ���龅�g?�y�?'I?�O���bb�ߥ��I־uQ�>#�? ��?T?q����=����*�=�7?�2?�%>A���5���=6��>zf�>4��<+�ؾ��W���=�f�>�I??��,>�״�s!U�:A��������,⾓|�⤖<�����q���=�����v���=,���b�6��S[���_U�,0?���>Q%>���] ��*�����=�+n>7�]>Rm�=�&��3n�;󾙽P0�z���Z>�o%`>�0(>`<=˾��|?[I?�,?qC?Ed}>�->�p@�b6�>�K���?��T>[R� ��Rf=����r�����ؾ	�־k�c��+���z	>N���>��0>a?�=�)�<c��=t\v=�2�=��Z=V�=�ҽ=��=IS�=��>V�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>+<>�p?>;kM���-�&1��՛����u���!?�p0��/��(v>�F��2$����z~>_>��=�k���o��=ڀ�ܜ�=�=LQU>#@6>uQ=��Tܽ=��>?�=�X+>0c= ��5М��� =~2�=�F>=K(>K1�>&��>]�=?�Gk?�z9>�H1��ܾ�?����>圌>��>�F��4��>d��>@$?@�6?��U?ȹk>�iR�<��>��?���n֚��^C�6<2�͓�`'�?vZ�?׆�>��þkҾD3�ZfA��H�=�T$?4/?j�>G#>�D����#���(��]��ki=���=�g�M��,W.�[Q��.M���S=�־>���>�h�>��n>�s>F�w>���>�w�=�^���=�&e=���s���`�=m4e<r��о�;U��<��ú��F�cT�<)�v=�0 ���x<�v˼O5�=cM�>�F>|�>�ƀ=G����IP>2���!�J�IK�=�4�G��i�� ���/�=L ���>H�1>��B��Z#�>5G>�Lk>
q�?��~?7�3>Z9�m�о^;��Wm�l�Z��X:=�u=�Ku�r�.���Y�Z=J��s�����>:,�>���>0_�=~����8=g���[�C�G��>��^�dՆ��f�s�S�L����ݷ��q��BK>��X?kNu��f�=��?�O?�#h?��>��F=x�Ҿ9��=4�y���e��������G���r"?9%?���>�	�	�C��H̾L��o�>9�I���O�+���$�0����� ����>H��1�о'*3�\���q򏿽�B���r��ٺ>?�O?��?+Ea��=��"bO�H���ĉ��&?��g?jh�>V?�"?<���/�F��o{�=�5o?���?���?b�	>�>9^E���?Y�5?���?K�?�U?�	��1U�>&P>]�)>v�Ž�&=��=�ļ;�f>�~?�M�>`�>{�����ؾavȾ������\�߼P�)>�d�>��g>�n>p&�=���=��=��U>���>_\K>q��>Փ�>q��>'�������0&?�*�=��>~3?ت>�===����<��7��K:���*��)��9��̹�<�T8c�Q=�Xż>t�>�Eƿ���?��W>����g?���^)���Q>�AX>'�Խ��>�u<>�x>G��>�^�><+>�߈>��(>Ǻ���.~>����q0��v?��jP�!����+�>Jx����Vd.�����S���y�?Ծ�\��T���<6�q	��-��?�>���p��2�?	g�ڙ?��>�7'?�Ě��T ���E>��?Q2W>����ٔ�昿=`�����?�v�?�c>�>_�W?�?T�1��2�gZZ�+�u��0A�ce��`��э������
��{��9�_?��x?giA?���<�wz>颀?"�%�C���X�>�F/�4-;�+�?=�Q�>#B����`��WӾ<�þ� �J�F>��o?j�?y?#�V���輋/�=&�F?�Y?d�y?B�C?��.?8.}��0?�r�>y,?�?�O+?��<?y�>.�?>�F�=�����<h_��i���^#����������=Tb�=i�=}ܪ<�01=�j��+;���Ὂ(��.[��oe�l�L>�0�=�m=%�>�RD?V��>�o>8�^?XS=��S�N<���b`?#�>�A��9��hW��(s�n`=��u?�&�?�jM?�+>�`�����x>l��>���>Z��>���>������QM����>M �>
M:ý�x�P���L��z9=&�V>$l�>�>�v�=���>m��q���>��n�,s����4���A�x^3�2�	�{>NE)?��
?sڼ9��=����#g�r��>	�L?�Ɔ?�m�?�J�>,$����q��aV�#�π�>to �	J�Ū�2��T־�y��4QS=�����U��N@e>�����޾):n��xG�q��7`J=����E=�_�˾;m���=��>��ľ;S!��V��v��H?V�r=S[��jZ��D���`>�x�>�]�>�@ѼT�����A�G&����=���>Z@>
���#��$�C�����`z�>�E?�a?Tt�?���1Xq�n�C�*���s��Ħ�o�?ޯ>sK	?1�H>m��=蹰����)d�&OG���>�L�>��:D�����	�����%�О�>��?�D$>n?��Q?�#?�B_?�)?И?W��>�9��}V��/�2?Pp�?)	�=Yw��+�#���7��jR��F�>-<?�Pٽr�w>�W�>]�?�!?ژ\?��?�H>�辠�C�SJ�>���>/}Y�����o>B�G?l�>�1P?��?n�T>�C:�+E���˽��L�=f�>Q�1?�I$?s�?��>x��>p���f$�=ƨ�>�c?�1�?��o?�U�=��?@2>��>��=��>g��>}?nWO?��s?��J?���>S��<�/��a;��OEs��EO�p��;�7H<��y=���,t�MH���<3�;�ⷼ�a�����ӲD��萼F��;���>��Y>X6����D>�2Ѿ2����L>��Y�)���u���2����=��>�?�>U�J��< =��>���>ҡ��2&?�?�~?ǫ�;8f�>��4ё�o��>\�=?�.�=��i�2���l��ר<��s?MjV?!j���C	�(�@?��e?�"���Q���ȾA�T��\k��4^?|?�>�o��V�k>=�t?�Ub?4x?�uZ�_�s��u����S��G$��E>�D�>(@��PX�M܆>�&?#̞>6r�> �:>֖��8zo�P,�P��>���?��?]�?��C>�ы���ῳ��� ,���^?���>w����"?B%�͛Ͼ{Y���u���ᾃ����몾����}���`%�������ֽ���=�y?P�r?L�q?Q�_?'e ��c�4*^��)����U��������E��D��oC���n�C��U���2k���=@=u�ʣ\�	z�?~�1?��S�V?&�R��������J,{> �u��0��>�s	�w�=��K=$@}�r>3�E̕���?��>1��>O#0?kf�t�4��?�%�,�y���\>S~>&h�>H	?��L;��F���ؽA���s}�����&v>�tc?̘K?>�n?^w��1������!���/�CX����B>�r>�ŉ>̀W�j��}2&��T>���r�B��ct����	���~=��2?�D�>~>�H�?��?w	��J��Ex�3t1�⇂<P,�>zi?z/�>��>��Ͻ�� ����>��l?���>��>���rZ!���{���ʽ$&�>�>���>��o>�,��#\��j��O����9��u�=$�h?���(�`���>�R?O �:��G<�|�>��v��!�|����'�!�>Z|?���=�;>�ž�$�|�{��7���v+?�?� ���4&����>�#?M�>�4�>��?_͟>�z¾���?��\?��I?��B?��>m�*=�����˽p�*�* 8=«�>�&c>Mj{=���=�j��'d�$�%��&W=���=��Ӽ���bٝ;�X����^<�c�<��8>��ٿ��<�SGѾe������������ʽ�ˊ����ه��<������8Zl����v;A�Y�/�(l��w�]��8�?��?򧆾�i����m3���+���V�>��$�
�¼���T����3i�D4ؾ������$��0Y�g�P�T�ҷ&?���Ѯ��Ϟ����mw?�_?k#y?5q�x��N�5�,B7>�f=�7B�M!����>˿󂓾��_?k�>�|��&ؽ��>tؐ>�`y>�H�>�|�ӯ��$[���%	?D)-?&"�>@g�6�ƿo����d�<�M�?��@��A?��(����TX=��>�	?
y?>)�1� *��ذ��R�>�4�?���?�#N=��W����tue?to<[�F���޻H��=�y�=��=߉�ClJ>�_�>f_�/�A�g�ܽ��4>U�>�H#���Xe^�j��<�k]>��ս����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�}��=[��>c�>,������O��I��U��=C���؟��:�o(��B	=b)��}�<��u�"B��y@��(_�*�9��A־%ޗ�q��~�>Y��>���>p-C>ø3?�g?No�>z�y>�0]�&�2���ƾ��M��y��򴽅�=�qƌ=罾�BM��� �Y������:.�����F�+>p�A�6]���"�-�q�d�:�_k ?{�>먪�o[5����=A)پ5���A"��L���]����"�A�S�ǰ�?N�<?h}�� N��]�}`��Y{�Y=[?�lc�����|Ⱦ)�7>L{�=�>���>٢���U�js3���,��u0?>Z?_����[��1 *>�� ���=�+?��?ڂZ<%�>K%?��*�C)��][>�3>Lң>���>�F	>;���P۽�?��T?��] ���֐>ch����z��5a=u,>z;5�C��`�[>�I�<�팾>�U��[��\�<�R?Y�>�/(�JW��Q���[��v?=�v?��?L&�>�yh?OE?o��<���X�T�E���W=q�T?Ki?r >pf���Hվ�Ҩ��4?��f?��`>��X����-1�����A?�Ar?�D$?�J8�+���m��E���;8?91?C'a��a��@j$�?���45>�z?
��>�aO�$ޱ><g?q�q�v���ÿ��1�M)�?�q	@a��?$=NW|�J��>�?o�B>ޛ��;Yԕ�������=R�	?(Ý��n�j� �뙵�t�J?��s?��>v9t�KN����=ܕ��Z�?��?����a�g<H���l��m��A��<�ҫ=?��7"����(�7���ƾf�
������ܿ���>�Y@Q轝)�>
E8��5��SϿ����[оeSq�k�?��>6�Ƚ������j�dOu�j�G�]�H������f�>�.>_ؽH��[�t�jS7���=t��>Zd���V>�DT�T����[�<��{>|o�>�p;>����+��k��?3�޾��˿By�����F�]?��?3݅?�?4+������ݿ��AaM=O�h?5��?�??�u���Ml�����e?�¯�4H�����E�Nf>��7?���>��,�e��=v�>���>�Z>�x��������ݻ���?�?_�޾E@�>⚟?��8?�i���=Ӿ#�@��2=2L?��=Aʾi<�n�*�@*��.b?,?��P��,�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�
i	>���?�~�?Qj?���� ����U>
�}?2	�>�}�?���=���>?��=������8">pG�=�)��e?2�J?69�>�9�=��=��^/�3�E�3|P������C��P�>X�d?��M?�zd>6�Ƚ4�K�޹$�=���{.����D���7��5�M�*>,�G>��>�K���׾I�>>kO��+ٿ����Ʃ�?��>R?	f�|Fɾ\+�=�
�?V}>�H(�y��S�n��T��ڤ?��?��?Q���Z���]p��?s>ȫd>-ο�j�8�����
>g�?�b>�Z���q��j�]>�x�?_6�?3��?B{n���>�u0�
���Is�Z�Ծ�C��D��=Z�"?QO��׺=��?�g>���A��[ƅ�ۂ�>p��?3�?�I�>�7a?Fb(���0�=��'�>�rJ?��9?���d!�-�>Q�$?��9� ���f���*i?��@�@��l?����ҍ���+�������S�H�>٩<��6>�^n�e��=�;=>H>��>A��=�Ē>P$.��#+>ժO>��b>�ϴ>�V�d;�ݾ��(���$(�m�B���:�e=s�����)ն��=�$�ӾI�g�ڊžl�,��J�<w��g>��=~�I?f�Q?��b?���>ɧ����>v�m����� ��|�=]�>˝,?	U>?�=?��'=����X6k������J���͢���>d�g>d��>H<�>�(�>�ҋ��'>�-�>9xd>�h:>��=~я�xw�[��=| �>�Q�>HO�>�7;>�>˅���&���!h��lv��nŽ�?#����K�������D���=�/?M�>����/п`}��6~G?�[���"��(��S>�z0?a[U?�F>����sX��4>s���6k�*� >س�� mc�o>(�� F>��?�G>M��>�>���7�<�X����
a�=K�F? $�U�ξyw��~S�L�&�F�>]�6?�9}=�)��ɬ��e���)���'=Ø@?x��>� ���˾�^���æ��&>嚞>/	�;>b="A>�����F��`T��N>1[>M��=R`?-_)>*��=���>ӛ��Q�l��>��B>))>��??�e$?�n��ً�콁��/��iq>���>�W�>�5
>�LL�́�=֘�>~�f>�3�z��ߔ���G�q�Y>�"t�q&a�>�5�w=������=.�=�����?�p;=�~?���&䈿��9e���lD?R+?~ �=U�F<��"�C ���H��E�?p�@m�?��	��V�>�?�@�?��>��=}�>׫>�ξ�L��?��Ž/Ǣ�˔	�)#�hS�?��?��/�Zʋ�=l�|6>�^%?�Ӿ<�>F���6�J0����n�HI���> ??E������n4�oA)?�l�>d��G��~�¿��u�;�>��?5��?�R�`:���C����>[j�?�s?2h�>�p�u����0>��-?��j?�|/?����혵���>�1�?o�{?3I>���?Z�s?H��>:�w�ZP/�4��1����I==_d;�q�>ֻ>����5=F��̓��[�� �j���(va>}%=��>�C佦���02�=�^��gh��S]f�/��>�}q>�I>�]�>h� ?/b�>���>vK=�r��V���(�����B?�Ə?Q�	�4�j�{)�8�=��d��<?�2?iV�������>�GY?�?��b?a�>�$�v𜿨$��:尾tX�<Et^>���>%��>�D��r�G>9U޾�$p�~�>�:�>?{̼�澐�����.��Q�>4S"?���>tz|=��?��#?k�i>?�>�dE��J��$�E����>��>�%?<g~?Zp?Ƒ����3�p��'����e[�Z�M>��x?a�?at�>����}a��}+A��?�J|��њ�?̲f?�E��O?�?k6@?��B?��g>���]ھ�ƭ�^ׁ>m�?]<\C��5���"�/��>i{?q-	?jg�a���ڍ�t���̾ �?Jx?�e?0m�@�P!پM.�<�,�>�X=�(�=��8>��B<��˽�P>�"%>;��;� �A�LJڹ=��=f��>�]>\�������>ޝ#��	þH��LH�N[����>��;>i����yK?J���cu�H���ȟ�?�w?qL�?g��?ƫѽJ�e���6?A�?w[?��>ٿ��ؾ3%㾚Od�$�t�$�Z�>�x�>Ձ<=�պ�:퟿ػ��̇�C׽�~#��0�>
"�>z�?���>SӚ>���>�u̾&&�����	���Z��G�A�"���7��/�����)��~�<.����&����i>ķ���j�>\49?�\�>yE`>���>Tx��s^Y>:�R>�f!>���>=�>��>@�=�S_=��½��N?�a��"(���㲲�O>?k�e?Q��>����\��4��,&?�?Vݛ?��>�h���-�r� ?��>��v�N�	?׽\=�3�
�2<򓴾T
(�go���Z��7ȉ>d-�'�<�HJ��]�@?��?$�y��{ྍ�������_=���?x� ?:q-�ܚO��~l��S���P���<���y�������Ĩj�Y^���T��񀿍�)��Z<TL*?���?������������k�eR=�Y=�>$�>��~>*-�>R�T>����o0(�^yS��*��S���T�>]~?}V�>�p7?��4?2Lc?�_v?���>e�[>��ξG;?�G�<*�>�?�>��3?A�&?Ξ)?)K"?��*?�_X>bY�����9�~?�%?`�?w4�>`�	?.$���:�_'��'�l<����jѽ��=_�.=K���ŵ��1kl<1pz>��?��k��Q��ܾ��g=V�.?�?Vh#?R��yoþc�>�
?C'?AQ�>\H�|d��"��j�>k��?��ѻ/��<3>k�>�g�=.=�4z>#};-+=� ��n�=!U���>&=���=J��eB��$;x =�>)�>��?��>�>K���� ����H(�=��X>:0S>K>_پr}��L2����g��by>Ov�?:o�?�f=���=�=�e���N��k���� <�<��?}]#?�WT?K��?(�=?^|#?f�>o)�dM��&i��"��V�?�~+?�ۑ>�9�P\ʾ5���8]3��/?��?�	a�����(���¾��ҽ�>T�.���}����l|D�D����������dd�?V��?��=�E�5���o��G��A	D?�"�>⁦>Hi�>��)�C+h�U�F�;>�3�>��Q?�6�>]�m?�ϔ?jC�?�˹>�>��4��ಿF�<�=�>k�L?Q�?j�?���?B"�>{�R>��p���f��'��<tU��a�U�->/�>{�>�ߎ>�7Z>W4
>|F$=����Q�1�H$3>y��>r��>�>_�C>Ofѽl�b?f`?6E���t��|4�Asr�%�[�G$e?���?�M?�\���>���7�D�޾�� ?>,�?��?P-?�$���J�=&=���N���L��>0��>r,�>d���5�=V�$>�Ը>��>�	�ڒ�T�D�s*<Cl?Dq<?�D>}��\�^��!�����u恽�Ӕ���b�+"�Q���%>���2���w��Z^q��K��@ؖ�(����L��L���e�>1zj=��%>�>�=y>+=�.�9=�m�=dui=�� =u+�`�=�'7<�,Ӽ��觽F�L�Wo�=�"�=�e̾kax?��I?dT)? ,;?e�t>�>�>����>dh8��?��V>@�0�R(��2%:�3"�������߾.U޾��]��C���u>~d@�o�>��->���=�t�<a�=���=Q�Z=�-<
?4=D3�=��=�k�=F/�=>�>�6w?X�������4Q��Z罤�:?�8�>e{�=��ƾq@?��>>�2������zb��-?���?�T�??�?@ti��d�>K���㎽�q�=M����=2>n��=w�2�T��>��J>���K��B����4�?��@��??�ዿТϿ3a/>��
>�z�=%�Q���3��%Y���}���I��w?9�>�5]ʾ/�>�Q�=*���Ѿ,�=p�E>s��=���!�V��f�=�b��K�=� �='�>"�R>B�=TܽqI�=d =�:�=.QY>_��<��L�����ܹ�<X��=��6>b!->��?���>I=L?��?�`�>G��DY���оY��>��>�j�><����L>�k�>��@?}�<?�t*?�
�>0�ɽ��?�#?oaC��r��-o����3��Q+�?�U�?��>�ii����=�?�VQ��M�=4�?��?7-)?&Z>�U�m��,Y&���.������$E�f+=jnr��XU�E����k�����	�=so�>���>�>VUy>��9>��N>L�>T�>�>�<�r�=
ጻ�ʵ<���j��=������<�pż:��^&���+����l��;���;�]<���;k�=~c�>�N>w��>�#�=�����/>3Ė���L����=x����B���d��V~��.�-�4�ĻC>,cY>�?��|����?��Z>��@>40�? @u?� >�c� �վ�A��nd��WR��κ=�>b�=���;��V`�M)N�6�Ѿ���>��>�ۧ>�z>sQ-�@�>��Ȃ=�RܾhE3���>�\���<���i��z��������f�u",��E?����:��=��?~+M?�?���>8�����(�<>�{�$�<yr�|s��'���h?1�*?���>N��7H�{L̾"���ط>�DI�~�O�4�[�0����η�@��>g�����о�$3�ah�������B��Cr����>{�O?��?0b��V���TO����0���q?�zg?��>|K???�*���z�=t��^u�=��n?h��?<�?� >;�~=�K;���?��?
Ǉ?�I�?T�?�����a�>d���R�q=f��� >Фj>���<j�!<R��>6Y�>۹
?}�]�'�$��R�C4Ѿ��M����=A!<>K|�>*=�>�%�>x�z>�`P=�N<=w�u>j��>�ך>ڕG>剒>�Na>�:��[�(���,?}�e>�v>o�K?~��>/2=�y�3����=�-<��r�S���Ve��g(ǽ-�;Xɚ����<�<��>�zȿƔ�?��V>��(�r��>C���%���0>b��>mqx�6��>.=�>L�;>���>�<�>�'>Q/]>4��=�S��蠷=P���4����[���I�O�߾��>ϸ����۽�� ����<�л)D~�������z�r�z�&+�U�=��?B;��ry��o)���(�n?��>�GD?�2w�Ťͽ@�2>5��>8��>Q����h�;���ə����?"��?zBc>��>o�W?�?f�1�<3��vZ���u��%A�=e�ʺ`��፿h����
�:����_?�x?{xA?�0�<�?z>��?��%�g׏�p*�>9 /��(;��e<=�1�>�'����`�ĲӾ��þ�:�WOF>g�o?�$�?�Z?6WV��ck�B�#>)�:?�2?5t?F3?:T<?���hi$?�0>u}??�
?��4?%/?�^
?_>0>rv�=ns����,=�ᐽ#n��Q�Խ��Ƚi(���4=*�=Ŕ�:�o<�A=���<f��r���N;9��� U�<��9==o�=���=F+*?-U?R��>l��>Q~�?�x>�a��m��؇?�g�>��y�P+��F�^���NL>yJ�?��?�bH?��n=G�J����[>��?�?���>�K�>����V̾�a��%�>$��><�K>��<�ӫ���Ҿ5�t������q>f��>�A�>0,��O�=�M�x���̢;>��A�����z��A;�H�2�G�I����> �F?��?�$9=&V���g�|�a����>)�@?B:R?y�e?Vy
>Vخ���a�k����N��>�9>�l�X7���b��
?�^w=�r>�k��m<��0J>�8��徃�u��2L��f��K4�>?&��Ɖ>�|��K�u@>���8>�]>Ȕھ�����Ƃ����E=P?k����z���ȵ�0���V�>�	�>*�>�]=�"���G��N����>N>�>�o+>M �=���.�����T�0>�bT?2�Y?ws?,:	��:����^��*
��������C6?��>��?%��>�M:=>���_Y��x��P?����>��>M���:`��;��U�����xw>��?�t=&r�>(�]?��?ή<?�w@?ܨ?���>�f�����Ƅ?pߋ?�9T=��t�w�ݽ��'�q�@�V�?��W?����j�P=��(?�\?)/?="N?��?ϾH<^�#�]+"���>
�C>��j�ٜ��w�+>j`�?��>-��?�Ċ?� �>`dl�����I�p����� >�P?fh,?�T?���>���>*���Ή=EW�>��b?	�?K\p?/U�=6?�->$�>Ć�=9N�>(�>E�?UDO? s?'gJ?M��>��<Tǭ��=��	y���9�wڤ;>DT<ht=b����j��g��
�<�?;DϼO僼k|����F�����%�;	[�>��s>���+�0>��ľsN����@>�U��)P��=Պ���:�:��=��>��?)��>za#�٘�=Z��>f?�>���I7(?��?�?u�(;�b�6۾��K���>2B? ��=��l�(�����u��g=1�m?̅^?]�W�%"��kb?�^?�B�<�n�¾�d���꾢
P?t�
?+YH����>M�?2�q?"��>�fh���n��^���b�h&d����=�B�>U��p�c�$.�>��6?|q�>�0`>\K�=��۾�Yv��Ġ�~�?��?�?'؊?x�,>�o��]�tl��eH���^?�{�>�)����"?c����Ͼ����u��a�ᾈת����[j���m���$�0	����ֽ��=��?Gs?�Cq?b�_?7� ��d��?^�����MV�V����E�rE��xC��n��m�#�������jI=�����V��(�?�?G�����?����,W�����!>Vg�l�q=U��2�d��7�<�=��朧����ە��9�+?�'�>J��>�)?Sj�IC��;��_������Ӆ>��a>���=ik?�(>^�j��0F�3�Ծ�c��'�0->/�o?��<?I)d?�~==�R�������$�z��Ⱦ��>��>T>@$#�8J��c,��oK��z��pԾ�����o��{=��B?ϊ�>���=�Ձ?-�>A1���t����Vb��/���?P�P?�?Y��>��N��Q~�h��>l�z?
��>�m>��O�����/{�j�	�n�8?ڽ�>0!?��>d	ֽS9�=&��˯����r��\�>�A�?�̈́���i��>��?F��=ܯ�>Hr>��*>6�A�VR!� K�~��>�3?o0><��=d¾*^+�O��G"a���?3?־=�r��Ss>eL?m�	?���>�yz? o�>b+̾E>�(?;xd?��!?ݣ+?B��>��Խ�������/�ɏ�=r?�>^q>b�R�FZ>����ʾ���2=>D<C�T>�*q<N7�=�%�W���=8;�>+�okH���ž�־Y�����}����K=eo��i�(�BuT�LKᾭ\A�e�����=ŭM���1��R�l���_�?��?v��������ɀ��c�Ӿ�Q?𧋾��Z>K�(��ak��x��ܺ�6	����Y"��O5�I�i��'?8�����ǿ����1ܾV ?73 ?�y?��h�"�4�8�� >:
�<D ����s�����οС����^?���>���� �>*��>k�X>�aq>����➾�~�<{�?3�-?X~�>��r�)�ɿ����7H�<���?��@�|A?9�(�1��~�U="��>s�	?~�?>�L1�F�����N�>�:�?u��?��M=��W�u�	��}e?��<J�F���ݻ��=�<�=XU=���ՔJ>�T�>����OA��>ܽԶ4>jׅ>["�����~^�y�<��]>��ս�2��ț�?�]�-2f���/������>GoV?A��>���=��,?�vH���ο�Y�s7a?�~�?�i�?�'?-n¾4�>hܾU�L?ŋ5?/�>��#���t�n��=!��x�w����o9V�&$�=u��>R>�.�X���M��O�=��=O����ſ��"��d���=��˻��}�pY��Q��9�W�x����Mv�&W���w=��=1�J>�Q�>"�U>v�U>��Y?�_k?r4�>7(>>��܎���Ͼ��<x���
��;��A�%��џ�x6��	ؾ���������g�ɾ��o�L�;cFM��>���F/��u���1�<V?w��=��̾uQ���*�8о)���>��b7�l,Ѿli%��#e���?��+?w]����g�f.��ء:�q̻�*??��ֽ���L߾-U�=���@�𻲴�>y��<�ɾ�B3�� S�.�.?
�!?�¿�{��Dc9>S*꽡�1=ʼ)?�	 ?�sj<Tq�>|�%?���i�Ƚk\>��5>�:�>Δ�>�l>ҥ���
ݽ�'?6Y?Y�i|��;��>�w�������1;=%j>�3��й��Z>�@�<����{��z���̲�<{W?D�>�)�\���0��"��P7=< x?t?�Ѡ>�k?�B?e�<�_��d�S�r��r=��W?�]i?S�>?a���{Ͼ��<5?�e?TgO>�Vg������.�;$�|\?	�n?�[?i���}��1���?���6?��?�$r�����p-�����l�?���>�T�='�C�@�>��A?x��B ���7ɿ��e����?n@��?���>=j@�O�U<Z�>�4�>�{�|Z޾]H�û����=)�>�˾��c��)������2??��?�'�>p�F�ϑ�d��=�������?�?�m����<���8x�L6�)��<�ԩ=�0-��Tp�����`6���о�.�͡����m���>�|@�~�٘�>�Z�O!��4Ϳ�H��?���p�h��'?km>��ӽ8N~��0s��+q�qt7�0�A��u�8o�>c�=Z�-�Hӎ�������F����
P?s.L�Sk�>�o3��4־�`���Y8_߫>0��>P�~>����ھ��?|r�]�ǿ�Ǣ��T�y(Z?���?��p?�:?jQ�<�X������}���W8?��Z?��O?�$���ǈ���$�j?�_��vU`��4�sHE��U>�"3?�B�>R�-�Y�|=�>���>g>�#/�y�Ŀ�ٶ�E���X��?��?�o���>q��?ss+?�i�8���[����*�5�+��<A?�2>���G�!�A0=�OҒ�¼
?V~0?+{�h.�J�_?6�a�e�p���-���ƽ�ۡ>q�0�6e\��G������Xe�����?y����?^�?K�?ص�#��5%?��>W����8Ǿ��<J��>3)�>�*N>�O_��u>��\�:��h	>���?�~�?ej?ȕ������XU>��}?p��>���?���=���>A�>�㰾�7*>���=\<��~�?rU?p��>�%�=�:�,m.�b+J��N�����B�5�t>j�^?;�T?؂�>����kqK�T�%��5���G�K�<��h���������Wme>��^>2�+>x�_��-?����ؿ
���$�'��3?XJ�>rc?N��6q�@W����^?׆>�l��P���^��/���"��?I&�?IU	?=%پ�Iϼ a>!/�>���>~˽k{������^:>�TB?;��A���uo�^,�>^�?!�@h �?w�h��#?#����Lp�� A�����ݡ�4w>�=�>�1��p�>?|$?D�=��x��\�����͏>3��?�A�?�q?!g?f䂿Z�/��G=k{>���?u�?}
�$����%>z�>�G�����Y~�Y�@?]�@?2@7�c?�����&�����Jƾ�~=�e�r1<>��=(L?=޽ht潊)l=3A�=O�A>6>F0>O�=�W�=}��=�2�����!Ԡ�ޟ�n�]��)��V��D�%y�:��F@�0���y���P��@%b��D������x�J3� ��=:{U?��Q?��o?Ѣ ?�]z�߈>\���=��%����=�}�>n62?�L?k}*?rS�=�ҝ�Ikd�����R���&�>��K>���>�'�>T��>����J>W�;>(> G>"n#=�M$��x=��M>tت>d��>=�>BsT>Ȅ�=����+x��x�l�o�e�?�����?F���Rm:��������=(�/?1�=������ɿ=$����F?�෾N���Q6�J�e=��B?�sX?E��=�%����$��� >�����8��0(>z᪽O�9���T] >L�?�0>y�>`�C�+�#�/!F�r�Ҿxʮ=�(?��<���0RY���g������?�>X�>0�7�!��B���p���*���`�N>$Y$?/��>+d~=��ƾ��}�oF��]s>�5>-c2=Ӯ(>��(>�W):��4�1BG��nV=[� =��Y>P`?�w+>}��=��>c���#bO��ĩ>eyB>ǂ,>�@?�%?���a�����GL-�Ww>�*�>��>�>�VJ��F�=�n�>�?b>�6�=��������?�Q'W>��}�2,`��w�|=����;K�=)8�=8� �(�<�8\&=��~?���!䈿��l���lD?	,?�=��F<˂"�$ ��I���?A�@m�?�	���V�7�?@�?u��(��=}�>Z׫>�ξږL��?v�ŽXȢ�:�	�+#�uR�?#�?��/�ʋ�nl�;6>_%?ڰӾ�e�>�� ۘ�0��
�t��=\��>>CH?\H���L�[�8��<
?��?ɀ�Ǥ�5#ɿ4�u��W�>���?K��?��m�m���Z?�R��>�f�?�Z?�$e>��ھ8{T���>� @?��O?��>u���S'�3b?�c�?�҅?-�>]��?�jk?���>�<�N�ҳ���r���,y<�D��`�>0t�=g����%��ی��s���,k��~(��->���<[4�>�1��@ξ���<�l��,ߴ�E���wE�>C�h>L�>!Χ>��
?W'�>�٤>��F=WZ�ڋ}�b���,�K?_ď?>���n����<rn�=�_�B2?rO5?�A6��Ҿ���>,u\?�o�?QHZ? `�>D#�[���nE���a���Σ<�J>��>tx�>k���_�I>T.վ��D��;�>;�>�N���8پ�	���8��r�>��!?<��>ԯ=�m ?O�#?�i>�C�>5�D�6���'F�Ū�>��>`�?w�~?l�?����_h3�g��B��Ͻ[��O>�Oy?�@?2n�>C��R���D��H�K���w�?<�f?+8���?�?��>?�8A?��b>�p�t�׾�b����>\�/?��6an�+YK� �B�L?��C?��>�i�>G�3>�ʔ�RU��꤉=I�H?E�c?s�?�錾�#{��rI��jp=���-g=�v�<יp=��h>5/F>o=�'�>q��<��>�鼽(н�"{>\7 >�j>u<���9*=�4?-�ͽ��*���>M2E���>�cZ>mQ�=���h�m?q�G�p�����PT��M����ɞ?��?���?�@7=����[?a��?���>�/�>�3�������D��H��R�����Wå=�}?Q�<ýѾ,u����������Svu��k�c ?т�>N�	?��
?��*>��>ƿ�N	-�+$��b��\W��3�!]R��;�q��_����8�g]����Ǿ����Aٸ>��-�p:�>�?内>]t�>�ۏ>�dŽ*Ͽ>+��>���=���>���>W>�=M��<+$���ER?ǯ��e�'���0ر��$B?3�d?�W�>�c�'�����?w��?lZ�?2�w>h�|�*�2�?P|�>{��=
?��;=���M%�<�.��$�����8?�.��>PMؽ3b:���L�6g�*
?��?B����˾�X׽!ˑ���=Ar?\�?����LP���39I��]S�A���;�?�8�~��G�G�p��Ј�C���{����	�L��=��?=��?����~���d�_r���G��2r>/T�>��X>�<�>��=i�0���+��v���/��uA�ŉ�>1c�?�],>]?��3?�T>?�zf?u�>`��>��۾�m�>g�(����>���>�iL?d;4?��-?�
'?jH�>d$>�.�<�~ ����r?��_?'��>#��>���>x���#�h=�m���W<�9��j���9=��=����$��Ԭm=X{<={n?G���8�����h>9$8?���>��>�����~�����<,'�>��
?�4�>������p�����>�?k*��p=��+>̝�=N؄�C��4{�=_n��dh�=�w�ӧ<�)�%<���=|ד=0�l��0:r�g:@��;��<4�>ӂ+?�p>���=R��*
ؾ��V�ّX�:�>0��>�/�>��#��V}���^>���?���?>XW>�=->���=V����t������m��Y9>p��>��e?�'~?jr�?�OL?/RK?�t�=��A��`��O����0��Y"?�,?׊�>g����ʾ��z�3��?kZ?�9a�o��!;)�I�¾��Խ�>�Y/��.~�T���D��������_��	��?���?W�@���6�s�辈����_��S�C?�"�>�V�>n�>��)��g�`'�h);>���>yR?k�>��O?�5{?�[?5�T>��8�e2��AЙ�%�4�'�!>Y,@?���?��?(y?X�>Ϛ>3�)��F��S��K}�_���ڂ��U=B�Y>ȓ�>�>I�>t�=q$ȽY߰�A�>�̭�=��b>���>ڨ�>���>6Ow>S��<[F?��?!����]'��lx�pv*����w��?>��?7�+?�z�{(�2Q,��qܾ�>�[�?��?��?dvD��;�=wA�<�対�c����>�a�>NZ�>'ݭ<+��<Aw>�|�>�S�>���n���LTM�1����?9ET?,�=��ҿ��j���w����iFG<H���i[��b����^��;UZ�����h��~�B�uL��b���|�ľ����<���*m�>M�!=�@�=�*�==(�7�dE��K�4�%��;Db>3�=�Ll=��9��==i�k�)?=�è;I�=�W�;YO˾�o}?��F?��*?�{B?:�p>yx>	o9�|�>��z�	�?�M>�?G�$㹾�9�������Rھ"�پ�wa�X����>>�I�0>rb1>��=�L�<W&�=k`t=1"�=�'�*�=c�=�ʵ=5��=���=�8>%>�6w?X�������4Q��Z罤�:?�8�>X{�=��ƾq@?w�>>�2������{b��-?���?�T�??�?:ti��d�>I��y㎽�q�=L����=2>t��=t�2�S��>��J>���K��6����4�?��@��??�ዿ΢Ͽ-a/>}�!> �>�*W��q*�n}���\i�@�?�:;��D��eJ>�{�;�~���S����=߹�=�#=��Z���d�X��=l�t���M=i�!= �>98>�q>羽�B�=S$=��=��_>mt�<�9��{�y`s=�W�=L�.>y#>h��>�?Ua0?QPd?M9�>n�u2ϾC;��yE�>���=�K�>��=nHB>e��>��7?�D?i�K?X��>�ω=\	�>t�>أ,�B�m��Y�Sħ�kT�<��?�҆?s׸>��Q<��A�ԙ�_e>��ŽM{?	S1?(o?��>P���߿�$%��b1�|H����;+=g�|��[���G��$�	wཡ��=+R�>ee�>E9�>��j>�>.>�F>k�>ї>��<1x�= ��Z�<[-꼘xV=�^����H=\�Һ��<���;���:���|�~< (;���<Ɂ(<�۴;��>72_>*ҽ>0�Q>	�־S �=䆫��J���=	Q;�F�8�l��C���V�qԽ��u>z��>FGӼ�j����?-mb>�>��?�mh?=�U>*���m<��ϯ���^���R4�#�="Jl�b�E��U�K�\��Q���>�۟>�u�>=0h>Y�"�	�@����<�Fվ�y1��G�>Ynu�[�<����l�RT������Un�bUǼ�J?}����X�=U�w?z|K?���?#[�>:�����K�>Z���_�=b8�iu���}J��g!?�1)?�L�>����҉T�G%��g2����>�)��:�5�ប���*�6V=�j����>�������,:9��w��������c�Z�r���>��f?���?"'���vc��;��?�G��=�
7?��/?*y>F?S?I����
�o�8���j��W?��?{@�?��]>(��=1ǹ���>�
?U��?4\�?��s?l�?�;��>��)���>Vk��a��=J�>�Ǥ=v��= ?#|
?��
?=\����	�Dw��<��[\��]�<Iv�=��>D��>��s>���=]zc=�֟=��Z>˲�>I+�>�e>_��>lV�>�Iݾc9�-.H?.	)>�Z�>a�=?�(z>"ޥ<ϻ�` )���=��I=�*��ꪾ!#�a)�<�j��]>/��<L��>n�ҿ�֬?z�>����E0? 	���D=Bѻ<dV�>a����?4��>�P�>�� ?n�*>tA�3C�>3�!>��ǾZB>O�	��S���5�[�����K�>�ࣾ�$�i��)�ӽ2�?�ɾ�e�Kbt����K1�4�=i�?<��sZ�w���|���E�>�V�>��1?�戾%c��[>�:�>h�>ƅ�Fљ�ꮋ��9˾V �?�v�?�i>�ۛ>^_g?��?��ӥ?��1���y�{�G��]S��K-��ϙ���o3�̺����(?��m?\+L?V>j��>���?�u��-Ҿ^��>�b/���M�[�>v=?�>��D�����Q2��p��<p���ŀ?5�?�i)?��I��E��f���s��?�<�?�8�?r??n�_?|�v�U��>o����伾P)?�M?�m-?�P?��>���=��.>��>�@������G��q��c< �;���<5��=�y�[Ӛ=�M��kE����i���2�K�=�Jn��+^=��=�e�=�>�>|^?�f�>�>�I8?�$��=8��[���f0?�4J=-���6���.̠�s�ﾽu�=Bk?���?��Y?��c>�_C��>�3�>Z��>��->G\>Ͱ>1F�� �G��(�=c�>�4>�/�=��:�bc���
�n*�����<]I!>�R�>�ȇ=*~��n�Q=X��I ��ǈ>�oa���K����;�jT��T�Ś�=�
�>o{G?8M�>L��U���I���%0f�D�s?�??߾K?��?!�����}���K��i���;�>��!�n���鹵�ը����i��)��WM�>�ϕ�'������>rk
�����t�1��k�̾���>zB�M�s���㠔��`'�V|>O��>�簾��"�9��u3���;?�E�=����)����"�=`�>u�>�=>IS����j�@���8>=?i~�=9(��g�þ�WT��D��xvf>/,7?�r?�=�?v���<b�$=A�YJ��pžb1�=l�?�%�>B�? >ќ	>�S���I���N��@�J9�>�*�>MU�"�Q�]\ɾl8��%O��]�>y?�~v>A��>^�=?���><v?5?�[?fh�>�xǽ�����'$?��?I�.>g��F��p4��;����>8??�4��F'>:��>w�)?��?b\\?s�*?�b>Kؾ�1��ӥ>}o�>Ixn�@��3NB>q�<?^N�>?�~?�F�?�>�:��־K�����=��>�C?fE?�f/?�>NC�>uf����=���>;^c?P'�?w�o?�o�=0�?>!4>�*�>��=�A�>���>��?��O?�s?��J?��>>�<�#��5"��*'l�@O��Z};�wK<�u=��:Zx�OH���<��;�-���.|�4T��C�۲����<�=�>�"t>��Ru0>b�ľ�r���"A>�8L��񺊾�^:�S�=T��>�?�ʕ>[#�~Z�=9w�>�>"���#(?��?�?�=3;ٚb���ھ�L� ��>.B?���=�l�xo��
v�G�f=��m?�l^?��V������d_?�`?1ھ�5��.��*�v�O� �+5??(<?��C�v��>_L~?8�|?���>���,5j�K���k[\�I;T��=�v�>7��pW���>̝0?uZ�>�kY>�,�=]�վ���5|��$.?6y�?�U�?�ŋ?��1>�/l�����о����0y?���>D㣾�iE?�P�;� �*s���wj��ߺ�x���g޸�>���~�ɾ@��z�4Cr��>��!?�3^?�w?��F?���9�O��{�E���W�>�tj0�#�)�6p5�$u�ܢ+� �b�����l$�פ�`>��y��G��P�?�'?�s0����>(����*����ξ��C>J��� ���=�����=�m^=�g�6)�۩�KN!?�z�>B��>zd:?V�]��<��4�b�9�8���6>�2�>/�>���>��;��.����=�ѾÂ�����贇>��S?{X?>�i?��<��/�?���!O#�.�]=r◾o��=+�>a-?�|�����+����C�mb�����������=HC?�]L>�H�>W'�?��?�
L�]Ɖ�c55��0�&.B�z7=9�?m��>��/>���W��V@�>��o?���>�T�>Y�������>~�D��Z�>�>*O?�e>Z���Z�У��s�����?�־�=��v?�~��TbI�$��>�H?i�!��8�;9��>�za����ܾ� ̽�>�4?�>N��=$�¾���+�|�R����!*?��?�af���(����>��?���>[�>/܉?z��>z�Ѿ�� ��?WT?Q@G?�,_?SD�>u��=�Ɇ����-�� }<xN�>�m]>���=�M�=�2���C��B2��h�=���=�-滵 ��0��v�����1�=Ok>�X�=Ow�f�ʾ*7����|r�{5��EØ�8 �hoν��>�����lǏ���fN;�X+�$�#�R$��*l���i�?���?Z���Ծ*��/������:#-?|�R=,i�=fȾ,��<^���]�Ծ�躽�᤾�4�p{@��S��O&?	*��0ǿfU��͟ؾ�?q?,�w?��$
"��	7�!�&>���<�~Ӽ��������&οM�����]?���>Z��ԯ�8;�>{=�>cU>�3q>����U��(Ul<��?��,?�*�>0�}�quʿ�7���#�<�-�?+@�|A?'�(�d��&V=���>?�	?�?>T1��I�����U�><�?���?iM=��W���	��~e?�<v�F�ZOݻ�=�2�=-K=k��)�J>�V�>Ղ�TA�(>ܽ �4>�ۅ>x}"�����^��i�<d�]>��սg(��)Մ?!{\��f���/��T���T>��T?W+�>;�=��,?t7H�X}Ͽ�\��*a?�0�?��?��(?Vۿ��ؚ>��ܾ��M?pD6?���>�d&��t���=j4����Z���&V����=F��>̄>҂,�ۋ���O��F��d��=����ʿA'!��9�>��<���<_^��1���ʽ}\������L���b��Ul=���=��>>6��>��J>�N>"�\?עf?���>T8>l
'�����[ݾĨ<u�`�;����{y��jؽ� �����M�;�E����`)���ɾ�L��O�=�Ya�����a�Q,���5-��lL?�>�r��$�Q��yZ��M����M�=d�9=����Qu��(c���?��S?ъ�T:��nU��k�=>�=<%[?qW��-�����_�>���؛=���>첽N{���JBR�2(?"5?�-ľ�0��Qv,>R��f�x=�"*?s0�>!'�<�ҩ>M�*?�N�r���)q>�\<>�Η><��>-f�=贻�uԽ�?�S?{�ҽ.K���T�>�P̾k������=��,>��������>E�F�x<���C����\���(=%(W?���>��)�*��_�����Z==۱x? �?z-�>;{k?,�B?ؤ<Yi����S�F!�a\w=��W?@*i?.�>u����
о����տ5?c�e?��N>vbh������.��T�%?��n?^?-����v}����R��(p6?F��?����Ē��x�� ����?�>���>�=.�V��>]1l?�D>X���س��V?����?�(@�@��=>>C'��̸=^��>׌ ?����B"��*>D����v�=ѷ0?����CS��R���>�{�>�Y�?y��>N�������r�>`�Ǿ��?��?�i��z
�=i>�Y�v����W�0R�=;�}�d?��.� ��8A���¾ta��?��>?%=!��>�S@\�2��s�>�/G�v�ݿ�Ͽb��ް��t����?�I�>�s��z����Ld�p�O�O�r�7�����2�>��>#����t�{��y;�����(�>{�����>��S��������q6<a��>���>���>DL��.������?uH��37οέ��V����X?ic�?�k�?�`?^-5<B�v��{�,��.1G?�zs?�Z?x^%��.]��m8�=�j?�_��nU`���4�^HE��U>�"3?�B�>E�-�ʵ|=�>���>Df>�#/�t�ĿZٶ�G���r��?ى�?p�;��>i��?ys+?�i�#8��*[����*��+��<A?�2>������!�40=��Ғ���
?�}0?�{�J.�7�_?�a�W�p���-���ƽ�ۡ>��0��d\��H��I���Xe�����@y����?5^�?[�?(��� #�#6%?(�>�����8Ǿ�<���>�(�>7*N>D_���u>e���:��h	>���?�~�?Rj?ؕ������ V>��}?��>ם�?KH�=H�>���=1b��>Ў���&>���=��5���?�7N?9w�>�0�=�/��[,�V,E��pQ��I�^sD�_�>f�a?.�K?��e>+�½�%���!��,㽂"����	�5�9?#������.>��8>�[>I�5���Ͼ�LA?���˿piy�����8?�d�>�a�>q���.R�>yR=<�?�;]=_�B��Ө��t��1�9;��?��?�!?��j��=�<|k�>�?�	s�Ŝ����8�xtR>
�,?zkE�E��J�-�T[�>�Ϳ?"@w�?�\�B'?���߅��dp��_Ծ�q#��d�=��+?	f�"t>E ?ہ>��OA���k��>5��?�1�?��?�%d?"�u�s.���i=扛>2�h?wi�>�<=���q�`>��?<�(���"�Ծd�Y?��@�-@J�f?0�����ӿ	������6C��i&>7:�=j]>�A�G��<�m�<|��:�J���Ӗ=�1�>Νw>"@x>�.>�l>�
>uɅ�99��c��t ��F�;�.������H���|��׌�����E���TC��P��,�q��_|��ٽ��=I�L?n+W?��v?l?��v�[V>���D͌����귎=��>&�9?RB7?nA%?1�=�����F\�I�v�|³�f������>��d>]��> )�>�*�>�Qf���>��|>s�>w3�=-�n<_���W�<��?>�ͨ>E*�>��>4X�=�r�>(H���j���{��v���c��?�8��We����������G��ZV�>#)?�	n=�{�٭������f�>?�������sf��l~>�-)?�-?o&'>�d����?�(/6>`R���m���հ>�A��.����ן�=* �>>�2>t>W>jZP���K�W�[�B��=�iQ?�/W�RҾ�{���6��ן�g�?��>wF�=����d��q�~���7�.-��gL?���>��ɻO
��``��8/���>��>���<2?�=�٨>7۱�f���G�Ƚ��<?5>�ia>EQ?��+>���=-ˣ>�F��#AP�닩>nB>Z,>�@?� %?�c�~��hl���-��-w>4P�>I	�>aN>�zJ�;ɯ=�o�>:�a> ��}Ӄ�D����?�0,W>�}��Q_���t�}zx=,��Q��=n��=� ���<��C&=�~?���(䈿��e���lD?R+?e �=G�F<��"�E ���H��F�?r�@m�?��	��V�>�?�@�?��M��=}�>׫>�ξ�L��?��Ž6Ǣ�Ɣ	�))#�jS�?��?��/�Yʋ�<l��6>�^%?��Ӿږ�>S:���z^�T�F�������>�B*?mF�	��"�l,?���>l �B񧿱<ܿ��f����>�o�?�m�?��]��%���:����>���?�Z?��I>�hɾz�(���w>�[?׈,?�4�>L��M���?0��?�C�? ,�><��?DD�?�k>�ޱ�G'�p��ǎ��q�>�����>�)>����-6�W���}�ex��:;��"?\�@����>�!4��2��T>��&�Z����"%�m��>�o�>7T:>�z�>��L?��?���=��=���<!崾Wp�f1??���?Į���l�h�c<��=�7"��9	?G�,?S�d��J۾bA�>��Q?���?X?��>��	�Q���9&����ʾ�c=�7>��>p1�>���J�>���I������>�E�>�>�A���W��Wh�<�>?�l�>�A�=� ?nr#?�k>��>SD��ᑿxF�ﹾ>��>��?�3~?��?�D���%4��!��� ����[��zP>�y?#?1��>���N=��>$&��6N�x|���
�?7�g?(��K?�?Q??#_@?�b>m���)׾����F��>a�?�X���V�O�:����n7�>s'�>�h?��r��=���ac�C)�'��r�;?P^A?��?&G�@sw���
�c=�<�"�FYP���N=� ��V{�=Z��=Ѥ��Q�=�9>���=��2���,���󼨑h=��>��]=�gؽ2�.�
�7?dZ�)��X�H>Š`�m=M���>e�>{�þ�?�́=�J`�T���Q֜�9������?���?�/�?yN=gꂿ�P?�A�?8e?i*�>��̾(�}�o���ꮾhd����ؽ���>�����|󾴰��񹰿���Y���P����>$�>	�2?5G&?\>`�0?�-���h��ה��V����H��L$�a7O�&lG�J"�Eh�ӱ�|�y=��پ<���w��> �@r�>8A?�DM>�\�>�ļ>P��<�>>g�>e"�>/�f>��+>��t=*�����\KR?)�����'����ղ��T2B?�pd?,2�>�
i�,�������?��?�s�?�>v>�}h��,+��l?G;�>c���p
?�Y:=�B��X�<\V�����/��#�x��>�:׽�:��M�mf�Dj
?�/?���̾�7׽a�P���<���? �"?�&�Φ)��Ss�kc�]cD�̶ʽ=%��畾��#��u��[����x���0��̆D>4?a<�?J+&�^b��+m�I�t���Q�싅>_?��^>�ͨ>��W>1�%�&���H�b(�io����>Ua�?��>��/?�7A?��:?O�k?�T�>h�>6�_f�>�ӭ>��:v�p>DB?]B?��^?��?	�?�ْ>��=�=�T���*?^P?�V!?���>5�	?O�Ⱦ�l��pц��� �?� ��S���==)�d>+��jeX�wfٽ�'�>�F?�
���8����H�j><K7?���>u��>dÏ�o������<�v�>q
?ҏ>L���7r��o��_�> V�?�'�Z�=��)>��=����Jƺ�%�=e0ül�=�
����;��#<�m�=�Δ=�fw�3Է��:�ݍ;��< v�>Q�?ї�>MB�>@��,� �Ҹ�{Q�=�Y>S>�>�Dپ0}���$���g�cUy>Eu�?z�?��f=��=���=F����Y�����������<�?�L#?�VT?ꔒ?��=?k#?c�>�)�$M��@^�����d�?0x+?���>����ʾq����3�=�?�?�a�D���(��U��Jѽg�>1�.���}������C��
�����R���$�?˺�?�'<��6�1�辉ɘ�����n�B?j�>��>)�>+��Gh��T�9>Z��>��Q?���>��S?��{?R�R?U3�>@7��l��O隿�>��>��1?;�?]k�?�p?B��>\�>v$I�Hھ&�@|����Z摾S��=q��> �>\��>�9�>���<��˽��8��(��tw=���>6M?��>[��>D�">����mG?7a�>�����3�^憾����yTb�ֻs?� �?�(@?�����_�3p.����Z&�>_Q�?e�?;�+?�D���=گ���Ѿ�遾5s�>'�>6��>��3=��r=AaO>l�>�>c#�3��.=��O����?=�H?�=DZ��@���Ns�lC����<3�:���3�Xi�~���;69}�&���F���bO��/���"��/򡾸k��H�z���	?u��<�>#�>��ҽi�G����,�<lH/=�ޜ=�P=A>��>/M5=ʚ��TP�<��H=��
>�=;aǾxj?*�R?�8?D6G?_e�>eR�=�Vҽ�R0> �D���?U�3>�1=�ӾQ�\)�������Kξp5ܾ�3k�O���� >�F"���>�>0�=��<��[�=A�/>��=J<�<�
=�.�=��=���=��=S[>�=�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>r��=w�2�T��>��J>���K��B����4�?��@��??�ዿТϿ6a/>"�,<`g>��H��Z��W���n����f���??���:7�02�>�d?��=���^>�?�@>E~="���L����y��wc=�8л%1L=Yr��~>�Î>]L�<< ^���*=�L�f�=�+^>���=:3�;�,��$*)<�@�<���<��=a�>-�?�^:?a�_?(��>�e��I�پ�&ľ^��>��=>��>��w=�	�>K)�>K�<?q�G?�B?t�>�r�<~O�>6�>�9�������䢝�kM>=~G�?,ؑ?<��>M4��k u�����k%��p��G?]�G?�'?1��>o��c��sq$�f�'��̒��Dq<^t9=��x�Vہ�./��`�����0�=Ys�>q4�>CB�>A�v>��0>m�G>��>�*>�
=��= *�aΝ<�##�r;�=�a/���="����<j��<s�� ����N<�:%<zq�<t;�;M)�=N��>ME >�n?z->�T��^��>�Ͼ�&m��RU>0���G=��[�7'��zJ�"�C�M	�>�6�>��<����1)?���>�[d>E��?M�m?�Ύ>�:�D�f,��\L����E���=;��=�[�OS��`J��v���پ���>u�>`�>@�l>
,��"?��w=2��\5���>�s������7q��@��-���qi�9Ӻ��D?hE��ȕ�=�~?K�I?��?���>t)����ؾ:0>�F����=m
�aq��]��;�?�'?n��>�+�D��̾����8�>e�H�.�O�5Ǖ��0�V�鷾�n�>����XLо�3�cr�������B��Zr�,�>�O?��?Ub��U���OO�4���Ǆ�My?]g?6�>�A?+?ZL��[��%�����=c�n?W��?�>�?��>���=����x��>��	?.Ӗ?u�?�Ot?�A�8��>�*�;�k">�ޘ�y��=)K	>?w�=%�=��?Q
?��
?�H���7
�W�����_��=�4�=�ϒ>w+�>��r>���=1�h=ⵟ=9@[>ʪ�>B��>�cc>y(�>'��>����*���7?Xax>3�>%�??�H?䙼�ϋ��zL>j��>�1�@m���ǖ��f���)=�� >�n�=��Z=a��>0տ���?�'=��8�%�6?�HC�	݀����>��=���eǉ>˜<>�n>:�>B��>h}���>NK>r����>�����W�g e��b��`�(>c��� 3�3�վ5k=�<����P��ގ���s������I=?]�?�H�lDn��Ѿ!ٲ����>pH�>��?��y��v��90>�l�>�E>T6������U��q���(��?R; @�<c>��>��W?��?x�1��3�JvZ�E�u��'A�e�l�`�>፿𜁿P�
���j�_?��x?yA?mp�<�9z>ȣ�?��%�tԏ�x*�>./��';��E<=a-�>�)��w�`�îӾ��þ#8��HF>��o?�$�?sY?PV�Hh�(o�=�I?��L?�Z�?&�7?x�<?����?e�d>���>��>B�9?´2?O&?d=�>f��=C�<�3�=G�ν����D��lz�����d�<\�O=���P
��I�z���6=&?F�D9�̀��x��R�v=��=!�=���=�B�>�)_?��>��M>aZ6?[�ν��-�虢���>?��C>�������5n��bѾ��,>)�}?s�?�xY?r-d>�;H� PF�~��={�>'�+>��y>��>!f�H���0�m=�)>��>#�=�2�;��z���T������<D8F>ZR�>y2�>�a�	3 =Cȶ��u���t>٩=�����C��C9����Aٽ���>	�E?�	?�}B��$辅bU��=h���?�#F?�=?n�{?]@�=���n�J�B�L�«��P�?��s=d�����B|��� b�2�<p��>����^���O>��f���b�q�eM�[fо^�8>����=��,��0:��$Z�=s�*>�ϵ������W���}K?y=<p;��k$M�T�¾�%.>���>X��>��M���0�`�+�S�� ^=ܞ�>��>5!�;� ��IO�i�	��[E>"�D?�q?�9x?�6��U�lZ���ho̾�>ǻ��?�P�=�#"?r>�|J>&����D�g�qD�<?DW?
�6�Rx�a����'ķ�R��>�/�>�>�.�>�{6?�q�>J`�?�k$?;F?�@�>��}�K}��� ?Pѐ?�)>����߽M��p�4�5�#?��?������=��>�I?��]?2�[?�e?��k=	L%��J'�D�>���>Rr�	����u>�C?���>�"�?�Η?\��>m�O�L0�bH�&�=�d>��F?��>?��?��>X	�>�����~=Q�>ĭa?�G�?�p?���=,K?�n(>��>���=ꎟ>��>h�?�cN?��q?�hI?���>�<n������s���D�"��;�k<���=k��U�l�ٸ
�c1�<|��;!����~�� ���E��_���q�;�b�>�s>_��p�0>��ľ�F����@>�墼�C���Պ�Q�:�CϷ=疀>� ?��>CY#�O��=Ϝ�>�9�>���9(?��?�?��*;��b��۾͓K�~��>7B?"��=��l��}����u�@�g=�m?�^?D�W�!��A�b?��]?aX�C=��þ]�b�����O?.�
?��G���>O ?��q?ɷ�>Of��<n����*Cb�6�j���=k�>�Q�'�d��@�>g�7?fD�>��b>(��=	v۾T�w��q���?t�?�?��?�.*>�n��4�/����O����m?���>�̒���)?�I����Ⱦ�d��Z�������=��������������;�rX�������H�=)0?�xe?��y?'hV?��z[`�
Oi�̭����Q�����+y��$K�8�,���<�n�o������2{����=5���R��>�?Yk"?����?_)�� Sپ4���&�>L�{���ýBz=�k.��F=dA�<��]�������7|'?�H�>?Y�>,�/?�nx�y�0�"�E�1yN�=����!>l_�>��Y>@�>3�a��D6�;H0�P����)��j���>�dU?́n?z{?^��q�&��$�����4	b�N���Z�a>���>?;�m-,�v�B���O���[��~����Ǿ2"�F�>��>�i�>$�>:(`?y�>U1���j��9���f��3�n�?�E>�s�?�1?�d>w���ᭃ���>�P?2#?։�>EU�nO@�Xꁿ(�� W!?�d�>ϟU?XI�>�GY=�
 �h哿e���g�m�h�=��?Kހ�P�f���>�M?�d2��$ӽ..2>-��=�|��x� �Ž?`?]�?�!T>�2*>.�M��颾����x���ƶ?.f?!�����\��=J�H?і�>��>�ϖ?�>���Ym�=��>~�G?��)?��>?��?0Z�6^C��W$�E{�f��=�e>MP0>xQN=���;A㍾?��oE����>*�>�����������P�����1=&�
>`{�>���U�Q��ɾ��Fپ[7��ǒ�2���봾@<�<6ߒ�@���:���&�<�� R=��*��3L�CՊ��Hx�u"�?I��?s�޾=)���횿�]w�����
?󇢾p�L>�<��p�p���2�޴��(v������/�cP(�y�[��"?1�d��2ÿ���<0þ��>��?��|?������(�+,>��<�F�� +���οԍ�N�e?�&�>����O�����>�4h>�#7>�̌>ݘ��0��gf;'h
?'n?�K�>�!��	�տ����%=�\�?w�
@^zA?��(�[��Q�U=^��>��	?*@>�C1��D�� ���I�>';�?���?�pM=K�W�a_	��ze?�E <�F��޻��=*:�=/K=s���J>eQ�>���}:A��4ܽ�4>�ׅ>�?"����g�^��Ѿ<�]>��ս����ӄ?�w\��f���/�uQ���z>��T?�.�>���=�,?�@H�MvϿ.�\��,a?�+�?ݚ�?��(?�鿾���>��ܾωM?�?6?��>O&�4�t����=�w߼G���X��7V�L�=���>�6>Jr,���ϜO�il���g�=�o�&ɿ�Q �&j��Y	=HU)�;P���Y�ͽ��T��s��9�f��m
�~�b=("�=�Q>�e�>��@>�M>d!Y?.#m?X�>2�*>���˦��o�־y���܆�}�ֽ��m�,G��1������ʾe�����*��Zо�Y@����=%ih�P���*�*^��F�;�-�e?R]���z=��5�9{ýfOƾ��ԾZR'>�X��p��߃�/we�Y�?G�1?Zv��r�d��t,��ɕ=Qxq<�>^?Vѵ������A*>,�C��z�=��H>�M�<�V��uc�3�@��_*?�7'?�M��h��6Q9>�ˀ���;S&?�
?���=�ݦ>|E-?<q�Ng���.^>�S>|)�>=��>��>�]��آֽ�-'?M^?��3ݹ����>��Ǿ{ƚ����<��!>f"�?I�;?�->6�b=��x��ʊ�����<�'W?���>{�)���Bc����v\==γx?�?�/�>hzk?��B?���<�g���S�7��cw=?�W?g(i?y�>q���vо�����5?b�e?s�N>dh���龄�.�+T��$?��n?�_?`����u}����O��*m6?�F�?�M��=���7���Y�w�?`��>_q�=;�5����>��_?�A�,��]�̿��c��ä?:@�@Q�:>c��2��=��?6$�>'S���P������\��?�a>�?w�����_�sZݾ��/?ɹ�?��>�����s�=�达���?5̓?�ϙ��F3=+�#��r��^���꼱��=�4��(�=�	��5��־<������R�=���>�@h��5�>��d��~߿�{ʿ$���!���H�G�?��h>�՞�>$h�ʦw�W���CY��L�+����>#V>�ǽҹ��J�{�r=�r�μ���>�I�g֗>JnV�+%��������:(�>���>�@�>�6������%4�?�|���I˿J1������W?[j�?���?�-?��t��o�G�b��]�w<I?�bk?_�V?�Z���b��>�%�j?�_��xU`��4�uHE��U>�"3?�B�>T�-�g�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*�p�+��<A?�2>���I�!�C0=�VҒ�¼
?V~0?{�f.�[�_? �a�>�p�b�-�)�ƽ�ۡ>
�0��e\��H��/���Xe����?y����?7^�?F�?��� #�6%?��>*����8Ǿ�	�<ڀ�>T(�>~)N>eE_���u>a�=�:�Oi	>���?p~�?Gj?핏�����cU>�}?ٺ�>p7�?�n�=f#�>"�=�x���OE���">���=�2�ye?E$N?>�>��=	U7���-��E���Q�p�r�C�Jy�>'Qb?��M?�td>�����,�T]!�[;ӽ;�3�p��r@�#�����N7>��>>�>�A�NӾ�j#?�@�w�ҿ&匿G9�up?BGq>h��>\��\��<<b�U?H#7>�q�K�;A��0�v��?	T�?�v?����&ȼ)�+>��>0��>&c�����rw�l�B>l9? n ��3���Il�*�p>���?�g	@ l�?�7p��^'?��9���"�5�;,�`|��(=�=���>b�&����>�?P�
>����=ժ��k����P>7}�?�M�?�?Q�]?K���Q��>:��>�Y�?ɜ?��P�Pp��C�=��?Q�ʾ�k�����c?�H@Y@%e|?���L�ֿ��������)|����=O>�c>,}齐�=�sF<{�S;�o�<eB%>���>�M>�fa>�9>�j8>�'">_������\et��x�=��*�P}۾a�!�-����9��������M����ѽ�� �L�½�m<�w�ҽ��^���=S�U?�/R?�p?�� ?�yw�!N>�����=�$�d�=�Ć>��2?F�L?��*?�͒=�㝾��d��T���(������b�>�H>�]�>��>V�>��82I>��?>DE�>��=5�%=��к�A=�NO>0<�>���>�Ĺ><>(>�������O�h���x���ƽ�,�?{����}I��������3��q�=�K.?#c>�s��k�Ͽ6Э�Y�G?zv���A��*��>s�0?�W?V�>�����i��^>���Z�h���>�� �Z�i�]�(��K>�<?T��>�o�=�@��2=�]�u�f������>Z/?*he���z��>g�z�Q�(��U��>L��>�U=1s ������H���8=����=c,?�W�>!=}5��u�ܾ�l$�(�=�AY>o�~��w��=Q:�<��������7���P�=d[>RM?��+>��=�>����4PO���>l
C>ڍ,>��??�$?�x��������k�,��Fw>�(�>K��>JV>NJ� ��=���>�eb>?��iC��J]�d�?��OV>��~���_���t���{=Dg��5i�=$ܓ=�%��!=�%=o�~?Tz���߈����;����mD?p4?4=�=QSI<�z"�����L����?��@�l�?W}	��V�³?T2�?5K����=Fz�>�֫>��;i�L��?tŽIۢ�v�	��#�P�?%	�?�81�H���xl�B>�T%?f|Ӿ�W�>{Ͻ9<���x~���d���w��\�>��I?����G��o�F�?��>�������#Ϳ=�{��J�>*��?�$�?�Pr���	z0�t��>'��?,�f?�V	>�_׾�wV��i�>�4?��%?�0�>CE8��
D���?t��?%F�?-�e>!��?1\f?H�>Z�<?=/� ���D��P9+>i��=���>�4��S���3��ꙿ�f���@����þӬ�>ũ=���>����K����<����(�������?�9�>��)>E�>�h?��>�=�>`~G=xp��"&�I�~��-K?/#�? ���zr�p�<�̱=��`�E?%<8?]��<�ݾ��>�Y?#�?��[?�}�>�	�_-�����s%�����<�	3>���>x��>a�;�L*A>z�־h����>Z��>�@w���־BK��,H��hi�>�.&?Co�>�\�=��?�$?n�o>���>xC�=�����G��3�>��>&?l�~?a/?���� �2��O��w����t\�F�O>Loz?��?*��>�i��I���!c#��W��d��d��?�aj?{�ٽ/o?���?r{??�B?��_>�����վ`���& �>��?<졾��f��'(��F0�� ?�:?� >��>����2�c��Pz�Y�?�[9?:V�>�	��"8`�B�M���<�z/�g,�<�P�=��Z=DK>l�>����N> <�k|<wʆ���Z<؀�=rY�=vK>�2=�aŽ�k<rJ:?w����1�vbt>��G�`����l>��/<��� �?F�6=<]�Sű�����{���?�S�?�F�?��W<Tr��dr\?Bێ?e��>m��>�� ��ݾ1b9�:��1�/���ؾy�C;�]?M��=�ˊ�����.ɿ�ȍ����e���I�>sH�>��?�R(?�s=��>g��6��8���S$�n�f��>�M�F�=4J�k��|�zD�	䳼qKо(������>�@��^��>�?�X>e��>�	�>�� �+$�><��>�M>/��>0�>��7>xg�=�6v<�x��yER?u¾^'�<侂e���bB?�'e?V��>�+F��+����	��c?uג?:#�?Y�>�{f��]*�\a?���>^���~%?�;G=
���7��<C���$�HM]��a9���>�� �5��YH�wis��>	?�?�Lüؔʾ�﷽�{��8�=��?�n?���2�:��Z��?�f�sc��ߧ��GZ�=6ݾB�Eo�4"�����Z����%���>��?ZҮ?�D�s��ӂ�37l�R�2�%uP>�1.?��>u��>CMϼ����\���ln��}@��Rr��p?夅?H��="X?�-U?W�@?��_?�u~>~�^>�$���?�
L�$k>�T?�3?6�(?�=4?��<?{�?,��>�6��������B?�&�?N�9?	G`>2F?�����I{��վ��z2������<�=��1>>�>p�T<U�L��P�>~n�=_�?!}�#4:�h���Q>0�9?>�>��>�������)�#=B��>�T?Cg�>L;ﾯ�k��	�(/�>��v?�����<�4,>�v�=Ӕu������=0���aT�=9;L�� ���;%��=�ě=��;�9=.=;u��;��<u�>�?���>�C�>�@��� �U��e�=�Y>�S>�>�Eپ�}���$����g�4^y>�w�?�z�?d�f=3�=~��=�|���U���������Z��<��?7J#?8XT?Z��?g�=?jj#?��>�*�hM���^�������?N!,?���>���ޭʾ�憎\�3���?@\?�7a�����>)�1�¾��Խ��>zU/�-~�&��ID��������ja����?���?��@�{�6�p��ܻ���c��͓C?��>\�>��>2�)���g�	'�$;>���>�R?�λ><�O?Ak{? �[?g�S>G�8�K��Y���p^'��>�??S�?*�?��x?���>�r>η+��]ྋ�����$�m���まBIU=�]Z>W��>��>ߩ>���=FDȽ+̴�.@�E�=V�b>��>�ϥ>���>^Ov>W��<�.G?�`�>鈻����n9��s�o��M]��[z?Z&�?��0?MJg�Թ���?��q�c�>⢧?�.�?0�"?��N��V�=�޼�a���Qf����>���>���>��<=SC�= >ג�>ws�>p��z��a�9�OV�X?�LH?���=Hƿ��q�� r��T��.Q<����1dd�嘒�Dx[�q��=�����U�z���oO[��!���0��0������R|��#�>�t�=B2�=/�=�X�<݄μװ�<��J=:�<=o�k�35~<ȸ9��9λ�k�� � ��sW<�jD=��	��˾��}?U=I?�+?w�C?ҽy>�>�3�Q��>Χ���<?UV>HP�����iv;�خ��3&����ؾz׾��c�ZƟ��F>II���>�43>�G�=f;�<��=[s=���=��Y���=%�=|o�=�~�=���=n�>�7>�6w?X�������4Q��Z罥�:?�8�>[{�=��ƾr@?��>>�2������zb��-?���?�T�?@�?>ti��d�>K���㎽�q�=R����=2>p��=t�2�T��>��J>���K��9����4�?��@��??�ዿТϿ3a/>�O>�8<S�f��L�w��8���A#c=�F?I�9������[>��>��̾�����+>��N>b�=����)�u��q�=z�����=��=���=Ǌ�>�Ѝ>]�a�@�->�+�P͕=\�<>(�u>e�#���,i>�͐=�]��� �����>n�?�a0?xTd?�5�>n�'Ͼ�:���G�>#�=B�>ׅ=�wB>���>�7?��D?t�K?~�>���=p�>��>��,���m��j德ȧ�s۬<d��?+φ?�Ӹ><Q<�A�����b>�*Ž�x?�S1?j?��>���,O�ګ���/�+�>���F�<=d=�i�B�ӽ����'�a�>/��v��>l�>��>�pf>�>EP>���>w�>>���;�T�=�M������u�y�	�нI�>�F�=�@�=H_4=-� :#F)<Ĝ==��	Sý![ݽ�F�<���>\�a>�Z�>`�o>L��!�">����G��:�=1��>�W���l��*���;E��*��U>
��>>89�N����?C&�=��&>���?�4?q�k>A�_=S��4k�����m���r��^�>aE����R��[�,o����k��>��>�"�>7�l>�,�,)?�h<v=��GT5����>�a��EZ�����%q��<�������i��亯�D?�E���G�=�~?u�I?���?���>k;��Jrؾ��/>�J����=!�t q�2����?Z'?A��>�쾷�D�>����C���u�>`��in;��%���l.�#-$�E2�^Ԩ>Ѐ��F����=�u�������D�^�������>�e?V��?�R���Po�"@5��2 �
�X=8X?,l2?��>� ?�(�>&�����TYt�� ���i?��?���?���=m$�=����(?�>��?�З?�b�?KHt?�?����>�4�>T�f����=1�>�,�=�R�=c
?��
?)?	?�����?�����y�4�R��[= 5�=�>-��>�:n>f��=��=�F�=z?G>�ژ>z�>��Z>�F�>̤�>#3�]b�y*-?q�`>�?��?��i>y1k>��k��1߽��r<�E��⾾f�v�r�=��(���Q==��C>\�M=���>m%п�=�?��<upL��B?��.�0q*��p���x>�c>��?];�>3��=�-?��f>�=��?>z�~>�ո��e>���v���F#��Ug��i����>��ξC.潞�������2�߽B�ž}3����t�/Յ���/����=b�?F����b�g��P�Z�1�>��F>�c#?�H徽t���J�>�4�>�f�<"��Q���3����\�泒?Gy@�;c>��>K�W?�?͒1�43�	vZ�+�u�m(A�*e�N�`��፿�����
����!�_?
�x?/yA?�S�<.:z>T��?��%�dӏ��)�>�/�$';�@<=�+�>*��2�`���Ӿ��þ�7��HF>��o?:%�?yY?8TV����Y���e?� n?��?��A?ٕh?P/N���?+U�����>&<#?��?�;?�Y?��>�#>�)>`��=`���{nѾ������k�<L��GQ>L=^>��=t<����F>��n>�A�=����;�н���n�νo��۽?2=���>�^?>��>���> �7?����28����50?;�H=ڐ��^���졾���:>��j?=�?5aY?ye>hC��^C�<Q>���>�&>�yY>���>�P򽾶H�y�=�>��>���=@DM�TM���>	��Z���q�<� >N�>��i>|���1;>�A��������E><꼂�����w(r�ۋ���c<K��>��Q?$G�>�:��������ޏe�M.F?"?Ԕ"?!�?Y툾��T�;;�1Gu�*8����>�}>��	��e���磿~N��s��«>U��<4{�:��>�1��I�Ԅn�fgJ��GG�>��%������	��e۾`����>�x>��о|��p򍿨4��W�O?r��{���=������>�@�>� [>�*%=l����_D��U��a�g<���>���=��"=c}���F!�B���d9Y>!K?�uj?/	}?���ox��-:T��Y���Ǿ:ٻ_��>h�)>i!?;)a>u�=���"����{��N<�Sm�> ��>׹9�nRV������޾"������>d�+?Al>�>~V%?h!?h`d?��C? 3?'�k>b���Ⱦ�w-?�̄?E��<BEg��j��m$���L��]?�V?@��K�=>Y�>3%?�33?b�Z?��@?�c�=ѫ�H�8����>_9/>�
m��1��2r&>"j?��>H(k?g��?_݅>��8�����t�5�J�>o��=��y?��5?a�L?���>w��>���
�>g�>,fg?�?�n?�����?�`F=u�>:�\��J>��?0[?�ma?F\c?�@4?���>ʟ}����c���ҽ�ػ��M��w�\�������3	=dTr=H
L�&:�x��=���fU�Ͻ����d�>8�s>���#�0>�ľ6<��E�@>^M���C���ي�M:���=(��>M�?���>�D#��ڒ=��>3�>����'(?�??��;g�b��ھt�K��%�>KB?J�=��l�Vs����u��h=]�m?G}^?a�W����>�]?�i?׾/*-��e������	���1?x6?vR%�ӑ�>?L�?:�|?�`�>t���h`h�mR���c�W��O@=�n�>��8�`����>�Q(?ͽS>��>��<�f�v��[~]��?���?���?J}�?}��>�m{�yA�<��}֒���_?�1�>D꥾\#?(gf��mо�e��sЊ�f��,��*L���,��?����&�'����սZ/�=
{?ʍs?�Gq?�]^?�1��/c��l^��5����U��������E���C��B��m��U����������j=K�m��e�ن�?c�4?��ֽ���>��¾����lؾ�Μ>����轊C�=b[G�-#R<���;4������}�$J*?��>B��>+�#?]4r�)���A�A�M����xyG>��P>��Y>CR�>2ݻ�RB�/�Z���~>����X=�WL>��Z?9H?��X?�ǒ=�A�ݮ��}������羡�x�X6�>r�?�S���DZ�Ȩ.�d�!��B��w�Ͼ�}־4x�4�>��&?oӎ>� x><�{?�>�P�
�����s�V�~���g��H�> �n?�u�>�i�>"W��R;���>�\z?��>�ę>�c���%�sRo�V!!�C0E?�|?�A?I
>���,�x��~ɑ���{���>�ȏ?�E��I��=�=/8?�=e��W�:>�:�<|Ǿ$�̾2�齥�?�</?�V�=�:>쎢��ɰ������i�4*?Y0?5���r�2�˅�>)�*?�.�><�>�p�?�f�>6rԾ��\���'?6�Z?dV8?�R?�?.+9�~u���!������=;��>�Ng>L���PH>�k�0��	#���=�&�<�ċ=�����<����:]��r=�E>ӗۿ[�7�$���H�����"�i�����9��j�5�<؅�Ri��9�O�����&�<
2H�)�2���v�Mx�����?HB�?�▾��-�Td�E�¾"�>�uW��)>�ƾ�I �A�t������k��� ����Y� T]� d'?�#���yǿ ���;۾��?�Q?�y?��e~!���7���">���<@Nü��뾑���/�ο����_?�i�>���|��?��>$k�>{W>�s>�Q���\���ӕ<�n?%.?O�>8�q�"�ɿـ����<���?�6@5�A?��(��@���O=�v�>x�
?^xB>"�1�-B���Ν�>T5�?�2�?ϫJ=_�W��
���e?;�)<T�E��ջ=m�=�N�=u9=:�QsJ>mē>���>��#ٽG�2>l �>��߫��j]�]��<�_>��ڽ�敽	Մ?`z\�#f� �/�6U���V>��T?�+�>YC�=&�,?Y7H��|Ͽ~�\��*a?-0�?V��?&�(?�ݿ��֚>	�ܾ7�M?E6?T��>�c&���t�w�==ἎФ�=�㾢&V�f��=.��>C�>0�,�y��F�O��1�����=����J¿��*���.���}�Ľș����G��e�̿W�����H�w�J��/�=-d>� ]>���>�p>�F> \?]Pw?e3�>p��=�;i��c���ľD�C�ߡ�����	~{�e(���'������7���j�*����z�վ��/��vR>��g������;��[d�q�+���3?=�>�=��[�ڰ�Z�Ǿ�|�o=��н�v)�U�(���b���?��8?��s��r�es���P>$�$85?��d���G�����C>�P��]�=r�=t�>=�K���<�zOR���-?��?�k۾4�ʾoC�=��G�=ƀ?���>+��z��>4�.?�����
��=|>��I>�>j{�>~�=���fh5���?ҹ^?8V���5����>�����Ͻ�b�=�C���Y���@>�1>/]u=�x��B��Qd���=;'W?휍>��)�q�Zc�����'_==3�x?��?'�>cyk?h�B?qA�<	c����S���w=k�W?�!i?$�>V}���о삧�1�5?��e?.�N>�^h���k�.��N�;!?f�n?6`?�"��'r}�F�����l6?�t�?2t�$�����̾o��wv?SB?�Ɲ>$�M�&(*>Gg?���q{��ݗ����b���{?�z@�q�?�S->&=Z�݀�= �>7��>�1-���˾��
�2Pľ�5�=�P?�s{�����n��x��	�?4�|?:A?X�]��5��]�=��G��?'�?�У��<T��v�j����F��=6��= @�w,�o���¿4��I̾��������:ۭ�>h�@V�G��>�xV�%�ݿ�f̿�Ä��g̾%-t�(�?��>�`ýD�����d���{�S�L�*T<�R @���>�OM>��v��턾�rk��BA�g뤽�h�>�A���b>N+���Dݾ�9��ɞ�=(x�>5��>S�A>�G�mϾ2��?����ѿQ���-M��Lc?���?Y��?{C?��;|מּA�I�k�W��6?ha?��z?H�z<�x;��(���pv?�#׾cbV����WC����>�P?xe>�b:��b>���>d�>���=��+�7fпc����(;��{�?[��?2����}?��?�?�w��BV��FR���X�B���Hh?�	)>� ������-E��k����?��>�9��l�Y�_?�a�K�p���-��ƽ�ۡ>��0��e\�EL����~Xe�����@y����??^�?`�?���� #�P6%?�>o����8Ǿ�
�<_��>�(�><*N>�G_���u>����:��h	>���?�~�?Lj?問�����QU>��}?��>#�?&�=�l�>9��=���z6��##>�S�=�U@���?P�M?.K�>��=��8��"/��PF��RR�_���C���>O�a?rrL?Sb>�Q��i1��
!���ͽ�1��~缇�@���-���޽�S5>�=>��>0E�?Ӿ֮4?��(���ɿ&�y�W�i���T?�ҽ>s��>c��K��.T>��~?��>ު� ����x��<޻�?���?��?����n:=���=[�8>A?+:<�'h�[ȡ���<�i5?�:>�j焿eXN��x0>�~�?,�	@���?��l��W?��X����Vx���^��>m�2?d���[bd>�?�B�=�Cv��1���x�c3�>�_�?8�?�u�>��j?_
r���=�Զ=��>�p?�/?KE���	��n�1>��?me�����
K �7Wa?p@
@ռ@/�\?ޞ��"Iֿ$W��+[������	��=��=��>bB��iE=��o;�B������>�,�>S�>�	f>`l>�A>�b<>̴���r"���D��L<��|���A�9�K
��%����h�ƾęپMՀ�ċ�EV��kaY�a��yM��m�=��U?�R?p?� ?�Rz��>����Zx =��#��D�=� �>Z2?��L?��*?��=a���&�d�YT���C�����R��>�OI>rt�>��>�<�>a���YI>J|?>k��>�o >X&=�󡺕�=fO>�&�>f��>+:�>Na>�#>����ާ��vu�.�f�-A��{�?���1a:���������'���S�=h)?s.�=�2��YÿLh���G?����-�MT��Pg=��B?Z�^?�z�;���EӔ���w=��������B=EX��L�ս,���)>q/?e�>��!>,V%�
#�׶{�� ��PUZ>B�d?W쎾Nm�P�U�d�r��u�����>���>S}X�Q�+�4:��+ǆ����'�5>.�B?��?=Y)>�
��5��x�=X�ͽ��=�p�=(�[��q�=	�����=��������5>h�9>c?��)>u�f=��>	����B���>&A>w�1>
<?�G#?��Ƽb����6|�;�"�MEz>4��> �p>��="E�Ŕ�=���>b�s>w�e������o���-9���e>��`�(4r�����
�=�M��[��=��=&�	��~Q��tA=�~?���'䈿��8e���lD?T+?l �=�F<��"�D ���H��G�?q�@m�?��	�ޢV�9�?�@�?,��X��=}�>׫>�ξ�L�߱?��Ž8Ǣ�Ŕ	�4)#�fS�?��?��/�Zʋ�>l�p6>�^%?��Ӿ���>0�3�\y����I�)�H��zѽ.�>'6I?����e_=�T(=�9?��>�������!̿�Ax�(Q?��?�A�?䍃�T��.�7{Q>Z��?�N�?3�|=ۭվ̐��	x�>^�C?�I�>J�?%XV�uEv�P?��? �?�uR>��?��y?���>��R��v)�?��X��6��=:�<R��>W�v�FJ˾:0�����u���S�r�L/ž��>�xg=��>��h��1��9�=�:���K�4�����>nܰ>��%>�B>,U�>��>yim>�dk=�豽e�r�0���`,L?���?r���Kn�0��<�̠=c�_�0�?��5?��*�mѾ���>��\?���?��Z?�t�>��ߚ�#����ͳ�� �<GwI>�p�>�z�>�$���&L>�־��A��Ћ>�\�>����]پHw�����|�>W3"?�G�>|�=-�?�*?�L�>�h�>�s6��e��jM��@�> ��>w�?��?�?�$���0�����	룿 �j��f�>��?�A?���>�����F1<ܳ��A��_Zt?%Gh?%���?�ނ?��&?#<?�>R-��þ/�<�%�>�?$?>�#��Tg���=�����?q?ZK�>��̽���O;�?����ؾ��$?J�6?*��>��ɾX*x�'*��Q8=d�����;��P=ҡ۽��=5aa>����>�>��kD�Ǐ�<���=��z=a�>��w=3_���x���M3?�^�N��;�=y�j�:_7�0��>�(�=U���_r?p$从�{�sٞ��j��Cþnz?%�?���?\����{���H?R��?��? �?���VN���
�z��4~�O���k�=�h�>V�i�Hô�pN������'�����=|���>���>$�!?p:?�f�=q�>����Z,$�t�;��έ�i�J��9/���[��rA�<���x��¼A��=����8����>x>ߣ���˹>�/?���>ņ�>9�>��Y=�@>D>�wo>E}?��(>G�V>��N>~�>���RHR?������'����)˰�t0B?�gd?z�>�Eh�^��x��Y�?}�?[i�?�Xv>�]h�	+�L?�
�>���lS
?�:=�]�V��<)U��8X��������>�Xؽ�/:���L�tf�Nd
?�7? @����̾ɪֽ1)[���#=,��?\�-?;���A3��y����B�8�D����=e(��C��P}��}�u�����኿^?��E�辘��>��?r�?y2�"[�g����m��%3�@��>=� ?f5�=]��>~z�=e8%���A1e��^M������(?t��?�!J>�eN?j-?6�F?Ou?��?>���>�ܾh��> ��=�}>Y�>.�L?T?�F?��K?;cD?��>(�����L)�&�W?T�?Yt�>k�>�;�>����}@ν<�.�_�Ƚ?�ν�)L�*��۰>�=<��i��>>���>�%?z
�M�8�)� ��h>�8?���>���>�������� =���>;�?�v�>p����Pp�t 	��S�>K4�?�[�i��<�'>N�=��������X�=�X�<П=�lq�7vC�k�<���=��=�)�����;�p.�ו�;��<�t�><�?���>�C�>�@��� �d���e�=�Y>�S>�>�Eپ�}���$��m�g��\y>�w�?�z�?��f=x�=���="}���U��u�����E��<��?@J#?XT?W��?V�=?Hj#?!�>�*�YM���^�������?ʮ+?�L�>����Lʾ=訿��3�P�?7�?��`�ak��.)��ƾ�(ؽ�>K�-��}�%쯿�XD���tt�m/���`�?���?�@%���7���e���=�����B?kZ�>Q;�>x��>BC)�jf�]
��5>���>�zQ?�7�>CP?2�z?ZG[?�U>�8��g��ܻ��YC��!>�??�3�?��?��x?��>/ >� +�
�����X�#��b�m��2T=T�[>"�>��>�a�>
�=E�ɽ
���9>�jY�=��a>H\�>�>�>l��>:t>8<�<��R?�?�Ҿ9���wV�����Ͻ�l?&�?��D?�7���澌���Z��(��>v�?9�?�?�Ɇ�)�m=yF.=������K�g�>���>\�>*�Q�HY=UЉ>$�>{��>'�m��D��gT��份��>?��D?��=�ȿy�s���u�2��Ͳ <�X����e���{��RZ�`D�=؏���w �����Y�>����G��*˷��9��}�u�#H ?�=�G�=��=s�<��ټ�7�<���=Y��<�~8=f�]�x��<5~߼[���~��;Y�P<?=�e����˾m�}?�<I?�+?��C?��y>�>3�3��g�>�G���5?��U>9�P�푼�ӕ;�)�������ؾ�d׾N d�9���$o>iI� �>m!3>�v�=���<���=1:t=��="�\���=���=6q�=ؘ�=���=l�>m>�6w?V�������4Q��Z罥�:?�8�>d{�=��ƾn@?�>>�2������vb��-?���?�T�?:�?Cti��d�>O���㎽�q�=w����=2>���=q�2�Z��>��J>���K������4�?��@��??�ዿТϿ;a/>�>ZRv>!]�Q>b�7!��>���q�-?!aE��+��4�=���>��G��|��g>C(�<:!>W���m�9ؔ=S�A�:+��S�u��ٛ>1�l>��=��@�u=�rK����>��f>�}�=� j>,�=����L�=���>O��ڏ�> �?�a0?IVd?p7�>an��Ͼ�=��kH�>��=�?�>�Å=�wB>G��>i�7?��D?f�K?z�>߯�=��>P�>�,�=�m��q��ç�̬<���?�І?�Ѹ>�0Q<ݏA����Qc>��Ž�|?�Q1?Hi?�>,7��h忌b1�V<�<���;���2��Fy=�vZ��n��I.�*������`i�>��>�<�>���=�px>�0a>��>߄e>�i����̽��R���R=�z���b>ј�<�S�=���=?t=	�F>�g=�<���=���=�.ɺ��,����=�:�>#�9>�b�>�0>ҹ޾�D>"����L���r��G�Qr3���e�#\��+�:�S��G>��i>o�<N���w;�>�(n>�a>+{�?R?l?X^7>�?ｍH���4���F����0���^�O�C>T	S�X�&���L��P��}��Ɗ�>��>T	�>�i�>��� K�� �=u�˾��E�;C�>�l�f
��>�&�qŐ��ꬿއ��W�^^�=�F?�ߖF>I�?Q0Q?i	�?U�|>��'�dw��A�k>�" �7'��M��v���nz�W�A?p?AB�>��ev0�l?̾㾽��>�3I�Y�O�����0��Z�Ʒ��>�窾��оL%3�>e��"�����B�Ofr�4�>��O?K�?=�a�KZ���\O�u���5��m?�tg?�*�>�D?y??�T��I��)c���*�=�n?��?g<�?�>ep�< �4�-?DG?�0�?��?o~t?=������>�s2�x��=�Lн� �=8�>2>���>�'?��?�.?������Y�����9y���_=b�=��>�b>J��>�>�Y����ŽK��=�9F>i>~�O>1B> �r>����a-�� 3?��>,��>XQ?��>1>����=�=�v���cr��ĕ��؇�V��Da=&/>���=z� ?/ӿ�Z�?q�=>�|?�H�?�S��z���6>);?�?���>T�>@�Q>���>�G>�?�<�#�=R�>D����6s>)m����$��Y�e8�K�>�����x:�hs�:ˑ�SM�=���\��k�l��*��G%�c�=���?y����}��~	��=p����>Z~>��(?�~��������>��?#�>���\v���̒�6�� �?(�@�;c>��>/�W?
�?2�1�,3��uZ��u�[(A�e�U�`��፿����
�d����_?��x?yA?�S�<2:z>J��?
�%��ӏ��)�>�/��&;��=<=�+�>*��!�`�R�Ӿ��þ.8�
HF>��o?3%�?fY?�SV��7���Ϗ�Fo�?�P�?i�?VP2?�ml?�|��f��>¬��i� >�?7�?E�?̫H?}S?ɍ�=�*>���<q̡�UԄ����7Aʽā�d%�=�1>��->l�P=𢏽F�=�?<�<)��;WZ���@s�����=Ѯ>��>��k?F2�>��>@?����2�H���fN?�BA>'����������@y�����=�*|?CS�?M�D?��>���˱�j/>?5�>o$o>�>;ߵ>(��P���?<CgL>r%�=jj�=��'=sud��� �<2|��'=c�7>%��>�K�>,�Z��� >�}��ɆF��[w>���/B���7�P	E�g�-��j����>��:?�c	?z-������W<j���6?�c??�P?Ю�?5ޥ�k��,O�5�h�zԺ�U|�>_�V<u촾R��H:��F�i���&�>�J��m<��0J>�8��徃�u��2L��f��K4�>?&��Ɖ>�|��K�u@>���8>�]>Ȕھ�����Ƃ����E=P?k����z���ȵ�0���V�>�	�>*�>�]=�"���G��N����>N>�>�o+>M �=���.�����T�0>�bT?2�Y?ws?,:	��:����^��*
��������C6?��>��?%��>�M:=>���_Y��x��P?����>��>M���:`��;��U�����xw>��?�t=&r�>(�]?��?ή<?�w@?ܨ?���>�f�����Ƅ?pߋ?�9T=��t�w�ݽ��'�q�@�V�?��W?����j�P=��(?�\?)/?="N?��?ϾH<^�#�]+"���>
�C>��j�ٜ��w�+>j`�?��>-��?�Ċ?� �>`dl�����I�p����� >�P?fh,?�T?���>���>*���Ή=EW�>��b?	�?K\p?/U�=6?�->$�>Ć�=9N�>(�>E�?UDO? s?'gJ?M��>��<Tǭ��=��	y���9�wڤ;>DT<ht=b����j��g��
�<�?;DϼO僼k|����F�����%�;	[�>��s>���+�0>��ľsN����@>�U��)P��=Պ���:�:��=��>��?)��>za#�٘�=Z��>f?�>���I7(?��?�?u�(;�b�6۾��K���>2B? ��=��l�(�����u��g=1�m?̅^?]�W�%"��kb?�^?�B�<�n�¾�d���꾢
P?t�
?+YH����>M�?2�q?"��>�fh���n��^���b�h&d����=�B�>U��p�c�$.�>��6?|q�>�0`>\K�=��۾�Yv��Ġ�~�?��?�?'؊?x�,>�o��]�tl��eH���^?�{�>�)����"?c����Ͼ����u��a�ᾈת����[j���m���$�0	����ֽ��=��?Gs?�Cq?b�_?7� ��d��?^�����MV�V����E�rE��xC��n��m�#�������jI=�����V��(�?�?G�����?����,W�����!>Vg�l�q=U��2�d��7�<�=��朧����ە��9�+?�'�>J��>�)?Sj�IC��;��_������Ӆ>��a>���=ik?�(>^�j��0F�3�Ծ�c��'�0->/�o?��<?I)d?�~==�R�������$�z��Ⱦ��>��>T>@$#�8J��c,��oK��z��pԾ�����o��{=��B?ϊ�>���=�Ձ?-�>A1���t����Vb��/���?P�P?�?Y��>��N��Q~�h��>l�z?
��>�m>��O�����/{�j�	�n�8?ڽ�>0!?��>d	ֽS9�=&��˯����r��\�>�A�?�̈́���i��>��?F��=ܯ�>Hr>��*>6�A�VR!� K�~��>�3?o0><��=d¾*^+�O��G"a���?3?־=�r��Ss>eL?m�	?���>�yz? o�>b+̾E>�(?;xd?��!?ݣ+?B��>��Խ�������/�ɏ�=r?�>^q>b�R�FZ>����ʾ���2=>D<C�T>�*q<N7�=�%�W���=8;�>+�okH���ž�־Y�����}����K=eo��i�(�BuT�LKᾭ\A�e�����=ŭM���1��R�l���_�?��?v��������ɀ��c�Ӿ�Q?𧋾��Z>K�(��ak��x��ܺ�6	����Y"��O5�I�i��'?8�����ǿ����1ܾV ?73 ?�y?��h�"�4�8�� >:
�<D ����s�����οС����^?���>���� �>*��>k�X>�aq>����➾�~�<{�?3�-?X~�>��r�)�ɿ����7H�<���?��@�|A?9�(�1��~�U="��>s�	?~�?>�L1�F�����N�>�:�?u��?��M=��W�u�	��}e?��<J�F���ݻ��=�<�=XU=���ՔJ>�T�>����OA��>ܽԶ4>jׅ>["�����~^�y�<��]>��ս�2��ț�?�]�-2f���/������>GoV?A��>���=��,?�vH���ο�Y�s7a?�~�?�i�?�'?-n¾4�>hܾU�L?ŋ5?/�>��#���t�n��=!��x�w����o9V�&$�=u��>R>�.�X���M��O�=��=O����ſ��"��d���=��˻��}�pY��Q��9�W�x����Mv�&W���w=��=1�J>�Q�>"�U>v�U>��Y?�_k?r4�>7(>>��܎���Ͼ��<x���
��;��A�%��џ�x6��	ؾ���������g�ɾ��o�L�;cFM��>���F/��u���1�<V?w��=��̾uQ���*�8о)���>��b7�l,Ѿli%��#e���?��+?w]����g�f.��ء:�q̻�*??��ֽ���L߾-U�=���@�𻲴�>y��<�ɾ�B3�� S�.�.?
�!?�¿�{��Dc9>S*꽡�1=ʼ)?�	 ?�sj<Tq�>|�%?���i�Ƚk\>��5>�:�>Δ�>�l>ҥ���
ݽ�'?6Y?Y�i|��;��>�w�������1;=%j>�3��й��Z>�@�<����{��z���̲�<{W?D�>�)�\���0��"��P7=< x?t?�Ѡ>�k?�B?e�<�_��d�S�r��r=��W?�]i?S�>?a���{Ͼ��<5?�e?TgO>�Vg������.�;$�|\?	�n?�[?i���}��1���?���6?��?�$r�����p-�����l�?���>�T�='�C�@�>��A?x��B ���7ɿ��e����?n@��?���>=j@�O�U<Z�>�4�>�{�|Z޾]H�û����=)�>�˾��c��)������2??��?�'�>p�F�ϑ�d��=�������?�?�m����<���8x�L6�)��<�ԩ=�0-��Tp�����`6���о�.�͡����m���>�|@�~�٘�>�Z�O!��4Ϳ�H��?���p�h��'?km>��ӽ8N~��0s��+q�qt7�0�A��u�8o�>c�=Z�-�Hӎ�������F����
P?s.L�Sk�>�o3��4־�`���Y8_߫>0��>P�~>����ھ��?|r�]�ǿ�Ǣ��T�y(Z?���?��p?�:?jQ�<�X������}���W8?��Z?��O?�$���ǈ���$�j?�_��vU`��4�sHE��U>�"3?�B�>R�-�Y�|=�>���>g>�#/�y�Ŀ�ٶ�E���X��?��?�o���>q��?ss+?�i�8���[����*�5�+��<A?�2>���G�!�A0=�OҒ�¼
?V~0?+{�h.�J�_?6�a�e�p���-���ƽ�ۡ>q�0�6e\��G������Xe�����?y����?^�?K�?ص�#��5%?��>W����8Ǿ��<J��>3)�>�*N>�O_��u>��\�:��h	>���?�~�?ej?ȕ������XU>��}?p��>���?���=���>A�>�㰾�7*>���=\<��~�?rU?p��>�%�=�:�,m.�b+J��N�����B�5�t>j�^?;�T?؂�>����kqK�T�%��5���G�K�<��h���������Wme>��^>2�+>x�_��-?����ؿ
���$�'��3?XJ�>rc?N��6q�@W����^?׆>�l��P���^��/���"��?I&�?IU	?=%پ�Iϼ a>!/�>���>~˽k{������^:>�TB?;��A���uo�^,�>^�?!�@h �?w�h��#?#����Lp�� A�����ݡ�4w>�=�>�1��p�>?|$?D�=��x��\�����͏>3��?�A�?�q?!g?f䂿Z�/��G=k{>���?u�?}
�$����%>z�>�G�����Y~�Y�@?]�@?2@7�c?�����&�����Jƾ�~=�e�r1<>��=(L?=޽ht潊)l=3A�=O�A>6>F0>O�=�W�=}��=�2�����!Ԡ�ޟ�n�]��)��V��D�%y�:��F@�0���y���P��@%b��D������x�J3� ��=:{U?��Q?��o?Ѣ ?�]z�߈>\���=��%����=�}�>n62?�L?k}*?rS�=�ҝ�Ikd�����R���&�>��K>���>�'�>T��>����J>W�;>(> G>"n#=�M$��x=��M>tت>d��>=�>BsT>Ȅ�=����+x��x�l�o�e�?�����?F���Rm:��������=(�/?1�=������ɿ=$����F?�෾N���Q6�J�e=��B?�sX?E��=�%����$��� >�����8��0(>z᪽O�9���T] >L�?�0>y�>`�C�+�#�/!F�r�Ҿxʮ=�(?��<���0RY���g������?�>X�>0�7�!��B���p���*���`�N>$Y$?/��>+d~=��ƾ��}�oF��]s>�5>-c2=Ӯ(>��(>�W):��4�1BG��nV=[� =��Y>P`?�w+>}��=��>c���#bO��ĩ>eyB>ǂ,>�@?�%?���a�����GL-�Ww>�*�>��>�>�VJ��F�=�n�>�?b>�6�=��������?�Q'W>��}�2,`��w�|=����;K�=)8�=8� �(�<�8\&=��~?���!䈿��l���lD?	,?�=��F<˂"�$ ��I���?A�@m�?�	���V�7�?@�?u��(��=}�>Z׫>�ξږL��?v�ŽXȢ�:�	�+#�uR�?#�?��/�ʋ�nl�;6>_%?ڰӾ�e�>�� ۘ�0��
�t��=\��>>CH?\H���L�[�8��<
?��?ɀ�Ǥ�5#ɿ4�u��W�>���?K��?��m�m���Z?�R��>�f�?�Z?�$e>��ھ8{T���>� @?��O?��>u���S'�3b?�c�?�҅?-�>]��?�jk?���>�<�N�ҳ���r���,y<�D��`�>0t�=g����%��ی��s���,k��~(��->���<[4�>�1��@ξ���<�l��,ߴ�E���wE�>C�h>L�>!Χ>��
?W'�>�٤>��F=WZ�ڋ}�b���,�K?_ď?>���n����<rn�=�_�B2?rO5?�A6��Ҿ���>,u\?�o�?QHZ? `�>D#�[���nE���a���Σ<�J>��>tx�>k���_�I>T.վ��D��;�>;�>�N���8پ�	���8��r�>��!?<��>ԯ=�m ?O�#?�i>�C�>5�D�6���'F�Ū�>��>`�?w�~?l�?����_h3�g��B��Ͻ[��O>�Oy?�@?2n�>C��R���D��H�K���w�?<�f?+8���?�?��>?�8A?��b>�p�t�׾�b����>\�/?��6an�+YK� �B�L?��C?��>�i�>G�3>�ʔ�RU��꤉=I�H?E�c?s�?�錾�#{��rI��jp=���-g=�v�<יp=��h>5/F>o=�'�>q��<��>�鼽(н�"{>\7 >�j>u<���9*=�4?-�ͽ��*���>M2E���>�cZ>mQ�=���h�m?q�G�p�����PT��M����ɞ?��?���?�@7=����[?a��?���>�/�>�3�������D��H��R�����Wå=�}?Q�<ýѾ,u����������Svu��k�c ?т�>N�	?��
?��*>��>ƿ�N	-�+$��b��\W��3�!]R��;�q��_����8�g]����Ǿ����Aٸ>��-�p:�>�?内>]t�>�ۏ>�dŽ*Ͽ>+��>���=���>���>W>�=M��<+$���ER?ǯ��e�'���0ر��$B?3�d?�W�>�c�'�����?w��?lZ�?2�w>h�|�*�2�?P|�>{��=
?��;=���M%�<�.��$�����8?�.��>PMؽ3b:���L�6g�*
?��?B����˾�X׽!ˑ���=Ar?\�?����LP���39I��]S�A���;�?�8�~��G�G�p��Ј�C���{����	�L��=��?=��?����~���d�_r���G��2r>/T�>��X>�<�>��=i�0���+��v���/��uA�ŉ�>1c�?�],>]?��3?�T>?�zf?u�>`��>��۾�m�>g�(����>���>�iL?d;4?��-?�
'?jH�>d$>�.�<�~ ����r?��_?'��>#��>���>x���#�h=�m���W<�9��j���9=��=����$��Ԭm=X{<={n?G���8�����h>9$8?���>��>�����~�����<,'�>��
?�4�>������p�����>�?k*��p=��+>̝�=N؄�C��4{�=_n��dh�=�w�ӧ<�)�%<���=|ד=0�l��0:r�g:@��;��<4�>ӂ+?�p>���=R��*
ؾ��V�ّX�:�>0��>�/�>��#��V}���^>���?���?>XW>�=->���=V����t������m��Y9>p��>��e?�'~?jr�?�OL?/RK?�t�=��A��`��O����0��Y"?�,?׊�>g����ʾ��z�3��?kZ?�9a�o��!;)�I�¾��Խ�>�Y/��.~�T���D��������_��	��?���?W�@���6�s�辈����_��S�C?�"�>�V�>n�>��)��g�`'�h);>���>yR?k�>��O?�5{?�[?5�T>��8�e2��AЙ�%�4�'�!>Y,@?���?��?(y?X�>Ϛ>3�)��F��S��K}�_���ڂ��U=B�Y>ȓ�>�>I�>t�=q$ȽY߰�A�>�̭�=��b>���>ڨ�>���>6Ow>S��<[F?��?!����]'��lx�pv*����w��?>��?7�+?�z�{(�2Q,��qܾ�>�[�?��?��?dvD��;�=wA�<�対�c����>�a�>NZ�>'ݭ<+��<Aw>�|�>�S�>���n���LTM�1����?9ET?,�=��ҿ��j���w����iFG<H���i[��b����^��;UZ�����h��~�B�uL��b���|�ľ����<���*m�>M�!=�@�=�*�==(�7�dE��K�4�%��;Db>3�=�Ll=��9��==i�k�)?=�è;I�=�W�;YO˾�o}?��F?��*?�{B?:�p>yx>	o9�|�>��z�	�?�M>�?G�$㹾�9�������Rھ"�پ�wa�X����>>�I�0>rb1>��=�L�<W&�=k`t=1"�=�'�*�=c�=�ʵ=5��=���=�8>%>�6w?X�������4Q��Z罤�:?�8�>X{�=��ƾq@?w�>>�2������{b��-?���?�T�??�?:ti��d�>I��y㎽�q�=L����=2>t��=t�2�S��>��J>���K��6����4�?��@��??�ዿ΢Ͽ-a/>}�!> �>�*W��q*�n}���\i�@�?�:;��D��eJ>�{�;�~���S����=߹�=�#=��Z���d�X��=l�t���M=i�!= �>98>�q>羽�B�=S$=��=��_>mt�<�9��{�y`s=�W�=L�.>y#>h��>�?Ua0?QPd?M9�>n�u2ϾC;��yE�>���=�K�>��=nHB>e��>��7?�D?i�K?X��>�ω=\	�>t�>أ,�B�m��Y�Sħ�kT�<��?�҆?s׸>��Q<��A�ԙ�_e>��ŽM{?	S1?(o?��>P���߿�$%��b1�|H����;+=g�|��[���G��$�	wཡ��=+R�>ee�>E9�>��j>�>.>�F>k�>ї>��<1x�= ��Z�<[-꼘xV=�^����H=\�Һ��<���;���:���|�~< (;���<Ɂ(<�۴;��>72_>*ҽ>0�Q>	�־S �=䆫��J���=	Q;�F�8�l��C���V�qԽ��u>z��>FGӼ�j����?-mb>�>��?�mh?=�U>*���m<��ϯ���^���R4�#�="Jl�b�E��U�K�\��Q���>�۟>�u�>=0h>Y�"�	�@����<�Fվ�y1��G�>Ynu�[�<����l�RT������Un�bUǼ�J?}����X�=U�w?z|K?���?#[�>:�����K�>Z���_�=b8�iu���}J��g!?�1)?�L�>����҉T�G%��g2����>�)��:�5�ប���*�6V=�j����>�������,:9��w��������c�Z�r���>��f?���?"'���vc��;��?�G��=�
7?��/?*y>F?S?I����
�o�8���j��W?��?{@�?��]>(��=1ǹ���>�
?U��?4\�?��s?l�?�;��>��)���>Vk��a��=J�>�Ǥ=v��= ?#|
?��
?=\����	�Dw��<��[\��]�<Iv�=��>D��>��s>���=]zc=�֟=��Z>˲�>I+�>�e>_��>lV�>�Iݾc9�-.H?.	)>�Z�>a�=?�(z>"ޥ<ϻ�` )���=��I=�*��ꪾ!#�a)�<�j��]>/��<L��>n�ҿ�֬?z�>����E0? 	���D=Bѻ<dV�>a����?4��>�P�>�� ?n�*>tA�3C�>3�!>��ǾZB>O�	��S���5�[�����K�>�ࣾ�$�i��)�ӽ2�?�ɾ�e�Kbt����K1�4�=i�?<��sZ�w���|���E�>�V�>��1?�戾%c��[>�:�>h�>ƅ�Fљ�ꮋ��9˾V �?�v�?�i>�ۛ>^_g?��?��ӥ?��1���y�{�G��]S��K-��ϙ���o3�̺����(?��m?\+L?V>j��>���?�u��-Ҿ^��>�b/���M�[�>v=?�>��D�����Q2��p��<p���ŀ?5�?�i)?��I��E��f���s��?�<�?�8�?r??n�_?|�v�U��>o����伾P)?�M?�m-?�P?��>���=��.>��>�@������G��q��c< �;���<5��=�y�[Ӛ=�M��kE����i���2�K�=�Jn��+^=��=�e�=�>�>|^?�f�>�>�I8?�$��=8��[���f0?�4J=-���6���.̠�s�ﾽu�=Bk?���?��Y?��c>�_C��>�3�>Z��>��->G\>Ͱ>1F�� �G��(�=c�>�4>�/�=��:�bc���
�n*�����<]I!>�R�>�ȇ=*~��n�Q=X��I ��ǈ>�oa���K����;�jT��T�Ś�=�
�>o{G?8M�>L��U���I���%0f�D�s?�??߾K?��?!�����}���K��i���;�>��!�n���鹵�ը����i��)��WM�>�ϕ�4����[b>��� �޾ �n�!J����O�O=MT��S=�]��"־;����=��	>	���� �����Ъ�7RJ?�<k=����U�͹��~>d�>H�>�l<�#Nx�x�@�ì�z��==��>d�9>T���ﾬzG�
��d>��<?z7}?��?��=j�m��D����M[��.)>B�?덪>�`�>��u>�V�>�vO�ؤξ��_��	b��s�>��?�5���|��m���Ӿ:/�V]�=�>x�,>�z?ϥH?�y�>��{?*�?'��>j
�>�=��&��K�$?r�?�]�=�W��A�0� U9�cVE���>ML*?��*����>0Q?�H?�>+?M�V?�U?��#>�f�mbC�nV�>�J�>�fX��>�� KP>��F?�5�>KW?Se�?�'->.D0�S�����C��=��>-/?��%?r?_�>5��>����H�=%��>�c?�/�?l�o?��=��?^42>8��>z��=z��>���>�?�XO?��s?��J?׎�>ọ<H=��k1���as��O�2;�;�&H<��y=˟�W"t��5�P��<	��;�a�����^���D�<���D��;���>?*w>Zl��e�>г���e�=�
>�3˻�E|��D��za����=\Sb>[�>��s>�LB��ŗ=8�>DR�>t���?�F?2�?�g�(�f�P߾�D�ǽ�>ӂA?��>e�v���0�r��u�<~�e?��^?�:�~��>�b?9�]?\f�=���þ;�b����n�O?��
?M�G���>��~?��q?��>w�e�{7n�����Cb���j�|Ͷ=�p�>]W�K�d��>�>��7?]O�>R�b>�,�=hr۾��w�An��7?��?��?���?S4*>��n��2�6F���U��#3^?���>c¦�?�"?h��^Ͼ�Ƌ��!����+�����֥��� ��$ $������ֽ��=�?h+s?�/q?�_? � �2d�f^����a_V�����E��5E���C�|�n���4r��@L��'�H=��R���_�Ϸ�?�;?PM�;Rq�>����p�ۥ	�|
>�����-��b�=7\��>�.>��̽�WٽMľ��$?dÈ>���>�D?�W�[�:��m'�'�E�*��`�J>���>Ӝj>R �>��2-��Հ�"��=ؖ�����Yv>��Y?0a?���?57!>*c�W���4���V=5�
�<�)>	�&>)̟> ������d������k���!� ���N���7>�ha?P��>�֚>	X�?�W?l���eo����2�F���5�n?��?�}$?SŁ>�A����+�`D�>�f^?`ܼ>�/>* ��W�"�8��q`�Tt�>���>&�?R+0>�L���V�JԊ�����j�-��[�>�W??Rf���M�V7r>:C?6�ϼ��<��>��Ѽ�+�_� ��E�ٖ�=���>Z�=�>R���5��+f��Y���?9b;?){<�{-����=4�?z[(?�h>���?�b�=e��q�A;�/?L�g?�4t?�$i?�R	?􄠾+/��E
�0�%��	>�?>;'U>HIɼ{h<��ʽ��4ս/
1<|�='��5m;��w:>?ë�����)z[=ka�=��ݿ@�L�CTþ�������"�����eD���G1�Ɍ�y��j񄾋G��c�潥�R���7��3Q�؉���ċ����?~i�?	�Ⱦ����I������	���S��>�Ͼ�6-ǽ��Sڽ)Yv�[�-�Q���rI*�R1@��1~��3g��X
?����sGͿ\+��K3�Z?�#F?�I?������Cx�\\@> <^>Y���0�;f���W̿�f̾un?�e?����B����?Kȳ>{�>�s>���;�S���\>xZ?z;S?�?���2²��'��6>ǽ���?H�@�AA?��'�C���\W=�`�>�x	?�?>�$2�c��������>Ej�?�o�?��O=�1W��2��d?ȯ4<��E��dK�=���=M� =i�QvI>���>o���EA����-^6>s��>�*'��x��`�|��<�a>�UϽW]���ӄ? n\�`f�8�/�/R���c>��T?�/�>�6�=ժ,?J5H��yϿ��\��)a?r0�?���?��(?�꿾�Ț>��ܾ݆M?�D6?��>�`&���t��_�=��༴�|��K+V�/��={��>�_>͊,�����O�'��D��=r���KͿ���i��R�<�G��=e3�9���B85� �ý��������	=����<),�=��U>��>iOe>J�A>�T?��d?�c�>k<�=N ��1�������=�a�Qٻ����qc��*d�h��߾����K���5	��y��9E�;�=�K�����Q�.��Wi���I��q0?�6p>\\��l�����Tľ�xZ���μ����d�ƾ�e@���q�ّ�?|N?�ړ��b�@�!�
sq��ԓ=�>g?�� �������,��<u==�>u?>��I�c[��A���G�9�#?��?~YǾ3O�����=~��r&ӽ�f"?{?W>���>s?s�Y�39���7�=�-�=@C�>�?۠6>{ï����!?9/?��%�ľq�P>ӣ��%Q���=�s>.'~�N���2$>d��as}�����,��/2��P(?�)>g�_�!�$7��d�P<~���xL?��>ix>z�A?���>Z��Ku��Mb�o�*��:d��_?OcZ?�Tu>p踾,�"�d��=֮	?�[�?�*?6�����0�J�^�P ��Y�> �?�1?M�l���w���@1?�;v?Ad6�����pt���~��k>,>��>7�>��K���V>=�a?��?����u¿[e<��H�?��@�k�?�1?�xv�X��_~?��#?8�ҾP���]�<�Wѽ��F?� e�7�����)��]��.m?���?V ?�h�u�)���>Eq��KԶ?ǔ?�ٽC�����E4�D7��)�;q	>at����@�8�����a��A\Ͼ�����2����A>�&@�0���@�>r蹾nd쿾���}�����8>V�Z3�>ْ�>�v�u]��  s��p��`{i��R���Z��*�>��>C۔������{�m;�?e��J�>���p��>YTT�2
��G����;<�В>/q�>ܚ�>Z���6�*ř?�P���Cο ���|��~�X?�p�?Xp�?2Z?h2<w���{�����G?Is?��Y?Į%��]��r6�<�\?�����Fj�u�4�8�4���>�  ?ְ>zs��3B=�o;>��>��o=��#�U�����{$Ѿ��?T��?��#�>�K�?��	?���hB���]ʾE� �R����9?d�b>~h���?�ho1�7ʡ��:�>��.?�ړ��{/�]�_?*�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>dH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�|�>d�?�S�="��>��=���H����f/>_>�r׼u�?�M?���>�m�=�@���.��nG�G O��&�!3C����>��`?=H?�Y>�ѽ�H�!��Ǵ��R"��kc�-�C�9!e�C��)6>C8>De>W5@��MվYN?���	�ݿ_����$��\j?�<8>>A�>�����폽$-#�O��?KH�>U��������s�[�Ӈ�?@��?�>��C��v(>wU�c��>Ο{>*���q�=�&#��o;=ntZ?:0�\���S�d$�>W�?$�?��?�u��?���k�u�\�R��Ż���*����=�'?��Ѿ�V����?���<�v��>��c)i�@ �>CD�?R��?[�>a?J�m�A�0��>���;_�6?#�?ö[��&����>N�?�ya��Ӌ�\�6��E0?7@,|@#%V?9���������aU�����e�W=e�<f>�0���L���ʽc���A�p�!��N�>ݒt>C�>5�}>�*�=��=0����!"���ί��U0��R ��!��Ǵ��d�H�jw��$s$��m�K����彯W:�.5L��{6��6y���+��_�={C?A�o?�T�?un-?�,5����=� ��$�= 漒�o=ӄ7>Q7?B�&?ڐH?m�i>�bg���V�#�������h@�x<�>gIM>|1�>��>���>�t<��m>��5>��O>�>t�Az�=_my>p��>�>ލ�>���>;�,>/,>�Գ�����Юk� ����ʽ�b�?����N����,����5�����=\)?�)�=�W��{EпD���wL?�	��)<�nv?�l��=Q1?�`?�$>�����k�>>��M�k��=�#�K�x��x*���F>�?ѯ�>/�>F�wp;�z)C�ž�Z��>G�<?�X���þ�+���5��
þ�:�=�8�>s$�=Ӵ
����ɯ~�,��\�m=`z%?b�>�D����ԾL�������'�>�>����q>���>N�>��!��"k�lAC=�I>�s>�K�>V�>�"����<3ǚ�Zу�$��h��>b��>�:|?^G? ��<�E�Z�:���Û�(�9>a��>U�u>K0y��>���>�t�<F��io��A]A��ǽ~�h>_�x=T��foU�6����=z��<�{��7�=�xȽ�~?���(䈿��e���lD?O+?R �=w�F<��"�C ���H��E�?q�@m�?��	��V�@�?�@�?��3��=}�>׫>�ξ	�L��?��Ž:Ǣ�Ȕ	�3)#�hS�?��?��/�Xʋ�=l�x6>�^%?��Ӿ�>��#����;��(�z�jt�= �>��*?�aվ>_���!��-7?��? �ھ0�$�ȿr�}���>L��?�X�?�[�|������R�?�j�?�51?��H>�:����1�>I�I?66M?8��>O��,�,��?�*�?HV�?xhP>Hǆ?�J�?�]
?r�<�@U�k����F��J�^>6�;�>�-{>]H��و~�憂�!@z���Q��p���(>$�F=�"�>1�`�]��qH >�$�ڍؾ蓒���>=1�>��>��>�k?���>ƾ!>v��=��:y]�������"9?�c�?�ྖHh�G� ����=���:
��>��C?����K�x�>��b?g�u?M#[?��>󵶾�0���f���������;��k>+�>���>>k����F>F7�)N���ޏ>���>R�=�6���G��y<>�`�>��:?Z�>{R<�&?\?$?JWp>"T�>�A�ǯ���C���>��>^�?B&{?o?!�y0�=���C����Y�CW>Xw?�? я>@���ɤ���,�.�3��W���d�?�g?���?z��?ʻ<?-1A?�T>�>(��%Ѿ<%��߱�>Oe-?���=F/�S����I���8?-�j?(s�>�������G^����8��夾�"?�J?2?���������Ӿ� 3���>���=�lͽQQ�B�T=B�V>��=�6}>���,�=�"D��X��������>>�?��>�y��V����+?��B�R�(!�>M�k��jw���>3e>���?�|=4t��)���pߠ�3d��Nx�?��?Ӹ�?e���?�y���?AN�?1D?|�-?�Ъ�ڭ��4�����;��#%���5���\>�ʝ>�?�=;{������Ķ�6���������+�>���>�?I�?�=@>,L�>#�|�z>&�q�4s�E}`�3!�h�>�.�&���	��Ň��L���"!ƾyBm���>���s��>�?��H>ĕ�>C��>,E;���>�`u>b~>�-�>h>��I>��>��;���P�Q?�����'��������A?vzb?�{�>Qd�!���� ��?_O�?U֛?��n>A�g�R�+���?m> ?����ag	?v�F=�Nr��x<� ������ς�����-a�>�N̽��8���M�r�i���?�6?⸐���˾	3�#!��B��=c��?�j3?i���a�KDk�OE�MP�l-h�%�b�/���p'�ڕ��:���gၿh�}��f"�G�G=g�?�u�?�J����!0��,�g���=�C�A>1?��>�s�>oam>��ˑ(�[vj�3/,���9��>OYw?j�>��F?��B?�W?�3R?��y>,&�>�<���_�>N^�<Sb�>�}�>�I/?j'$?��4?	 ?�	%?�S>"�������׾}?A�?@}?]N?u??��\�t��-)��Ӝ�Bd�f����=��d=��½�h��t�=xM>�?���M�A�d���C�=	^y?%/�>b�>�߾O�~����=\�?--|?��A?���
�u���X��x�>��?<Z	��	�<@�\>#w���F�<�ɻ�1f>F�7=Bd����>>Q���u��<����,(=S(�=uE>�C��3���;��|�>ص?�nZ>1L*>����������)�5�=�:�>�×>�.>H�Ծۃ���*��Ef��C>3�?�ٷ?+��=�@�=���=$ps��뺾/���������:�?X?��F?���?S1?Ļ?�$�=ZU	�&5���偿�ƚ��,? ,?E��>"����ʾ��)�3�E�?�U?�9a���A9)�3�¾�Խ*�>�V/��*~�����D��=������y��X��?��?��@�_�6��|输���Y`���C?�"�>�Z�>��>��)���g��&�3&;>֏�>�R?C$�>�a?5�u??+<?E��>�8"�G����߭�W�p=��[>��+?{ԇ?��e?�zU?X��>�b>����<žب׾��;�;�����t�=y�<>�>:��>U�>-ub>�Ӏ�)8�V�h�=��=]��>�p>$af=���>;g�>cc�=�G?��>B뾾ؑ�:�������6U@�YUu?�?_+?RO=�Q�r�E��U���7�>}D�?�Ы?*?�7T����=�ؼ@/��[br���>��>_D�>>g�=�&D=��>fJ�>��>g�����I$8��mM��i?��E?ْ�=y\ǿ�t���p�8���v�T<���?]`��E��T�e��"�=�0���)$�l׭�E�Y�옟�2���h ���y���Ox�ޅ�>O�=��=���=�f�<�VټW�<��w=S��<�h=�4L�H�<�.%�E��'m��ѓ���<`,`=�8ʻ��˾�}?e8I?V�+?��C?��y>#>�w3����>%*��_E?�V>�P�a���҉;�ϭ��$$��x�ؾXn׾�c���F>,[I��>y33>YF�=37�<��=K�r=}��=PV���='�=JD�=WK�=��=��>�P>�6w?X�������4Q��Z罥�:?�8�>d{�=��ƾq@?��>>�2������yb��-?���?�T�?>�?Ati��d�>M���㎽�q�=I����=2>s��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�6>�J>�WO���5��|`���m�S#����!?�@-�����R�>1��=�'񾉝־��z<��">j/L=�W��sT�b��=_XZ�V{=�B}=f��>m�:>$�=�ŉ�r��=7�#=���=A`L>��8�<���.�b�p=]͜=�O>�%>mu�>M�'?�*?�+X?�?�lK�<Ͼg3徶Y�>����~�>
��>7��={��>��7?L�?>�9?|��>�c=7��>�Δ>��W��6�/�����4��<��?��V?r�=v7>����G9�C_����2?jY?��?J�x>͞��2h��X�'����w�(l<)ܼ�����ń�i;=��Ծ��#�F�>5�>��z>V�>-�>v">��>�G>���=V��^�ֽ��<����䧀=�JW>Qq�<�_��>m�>�i�;k�<
�
��>���5v�E����=SY�>hZ�>�?�sX>V徒��>^D#���S��Tg=�ؚ��>_�x}��e���o�`u <}#�>q�k>L�\��l�����>Eq�>a�=��?�M�?�>Q��='��0ɶ�0���������=_�	=(/<�����g��CX�������>�֎>C��>�l>�,��?�bKw=���kQ5�R"�>#g��U���)/q��=��%󟿢i�Jĺ�D?�C��]��=~?{�I?gۏ?=m�>�E���yؾ�Q0>�-���d=]
��Jq�������?�'?%��>�
�>�D��B̾� ��Rշ>_NI�h�O�������0����������>�𪾼�оm'3�f��B���ōB�4Cr��>�O?��?5b�S��GUO�����S���k?�|g?��>�K?�=?.���y��y��r�=>�n?��?�:�?`�
>��=?o��g�>�?8a�?���?�jl?�!�X��>��F��[&>e�9�J9k=z��=,�=�@>Y�?P�
??��^�
���YS�>C���B=�7=j�>��>�6W>�>J.�=��=��Z>�(�>�|>��m>x��>�Ɏ>�֕������M?�>��?�n?�0I>�G�>������e=f���gS�Ma���@�</�g>J1I>��=�齾��>�@ٿ�>�?W�>�
�<�"?��~�!=�ȼbS�>M@���>"�>��v>`w�>bh5>�@r=�)�>>f >x�׾M�>#��d2��ze���O�ڧ���ǳ>��i�TM���*N�0B���ڽi�J���z+j���t�U�R�;DA�p�?|
-�����-�#�p�x�3a ?  ?~�?� �����ީ=*��>C?�>����K���1����	��Â?��?
Yb>b��>�+X?]?�7,��r3��iY�w1t��A��|e�fh`�8፿ý�x;��ǽ��7`?�.y?�)A?m�z<2x>�h�?�\%�9K��#�>��-�#6;��-F=��>[���^�D�Ѿþު��G>V�o?�߃? �?�LT��m��6'>��:?�2?�t?r�1?�O;?���z�$?�74>]+?�A?�5? �.?;<?�R3>��=������"=z���F����Mѽ�˽��．G5=�2z=���0
<)7=�}�<`���ܼ'�];̜���O�<�];=&�=��=lV�>Z�R?��?ṣ>�T?�71�3!�Th��0�?$V���9��K��׾]&�ܠ?>�ur?,%�?\TA?΁>�#*�D�I�pJ4>�>2�L>�T�>y�?>p<���.߽1��<�
/>�c�>�N>w�S���a�G�:Ą���>��V>��>���>θ>=�J�����w����#�>�� �3��yֽ�����ɾ��0���>�cy?�7?eh >�!��U�P�:��{�>ɭ#?� /?��{?���?�e�]� �e�f�i�a�>�	>&�JC��ҿ��]�'|���W�>})�=1�����c>��� �m�c�I�-�辱�U=�.���=���w+޾�w����=W�>�ſ�wE!�1���i��+�K?��m=����+W�/����>��>��>�
U���]�@W@�4+���`�=g&�>z�A>b�p�G����F�����E�>�sP?��c?�p�?�����m����k�5�6�����W�,<P)?��>Uq?#^�>J;>T����O��|�T��U��n�>��?�mJ�b	h��|j�A]�t�E����={[)?���=�f?�BQ?�?�xC?�K�>�8�>�K>��z����lW+?NP�?�
�='	��c�ʽ�\1�mP\�ŏ>RB?�!�d+�>�:?��?<H?c�K?�	?���=�Q� �N����>ɻ�>��G��϶�|��=�v?� ?dv}?Bb�?��,>}X#�������
=M1>6/?3h&?vM??Ɠ�>f��>:��+>O�>�d?��?�pm?��W>�e?��=
{�>���=���>�?l�*?��J?�o_?�4?ߙ�>t��=�͔��U%��	���c���f��'�����=���;�Wa��rT=r�%>�<�;�<H�=l耽Рk�]�=�_G����>�O�>�𚾜g>�˾+����G2>Fָ;����+��hB�">Ń�>=�>��i>A�]8=���>ʾ�>`� �!?��?�?� =�wf�w?�815��S�>��9?=��=�LW����wg�R��<7�i?]�_?�{ �U���b?x�]?c^��=���þ@�b�ۓ龤�O?��
?.�G�h��>��~? �q?���>��e��7n����Db��j����=�o�>�R���d��?�>��7?OR�>]�b>��=u۾*�w�2p���?��?���?��?s$*>��n�3�Od��=[���^?���>�_�"?�q��SϾ����q'����ᾙ@��I��}x���A���$�bჾ-'׽6�=�?�s?�/q?f�_?p� �>�c�-^�0���V�>�~���E��D�ōC���n�'w��0�����	�J=V�B�qt�L��?�1?�{��~��>��Ⱦ��L�%��4'	>�D�LI��t�xV�,i�=#�==��u�q,2�R#¾�)"?ߟ>7�>�bB?�%��ۻ4���0�6[���8�ν->SI�>� A>%�.?!���0����F��-�ؾ�ih��>���>k_?�xN?8v?Q���4�O�����4�q� k��uZ�>���=Q\�>����3������I�1�y�v���W��@����>ǖ?���>/�>��?GU�>�4��nN��P}���p�]��<KM?xT?N#?L�>��T��&Q��@�>�l?�Y�>�Š>B6��8� ���z��ný��>a��>��>�xo>�&�1�Z��Ď��	���8�<�=�Eh?x;���\����>�IR?g�<��<�{�>5h�����h�a!�.x>j?�?�=�f7>����1�
���z�����i(?tu?ڂ����%��L�>j4$?z��>�W�>,�?n �>"A��y��;�?�^?��I?m�>?V��>u1=s�Խʋ潌2&��ks=0��>���>vә=�f�=�>�ES��\��Q�f=���=n�'�PH׽0�o;�d�����<�(=��?>�j�؂]���Ҿ?4 �r���K�W�ʾA��D�B��m����Ѿ?���>~�.��st���,]�Ճ�����qx��^�?��@���	���Ⓙ��]�.* �� o>V_%�N$5�7/"��{Ǿ,举�{ؾ�ؾ4,-�=Z�p��lT��?�kr���ȿ���t
��?��$?Dm<?�������4G��=I=��W<r��q������ƿ��־esa?���>�jԾ�*A=���>��g>�->f�=f.��Y��!.��A�>�x+?��>�"���Cҿ֞����b�&�?��@�mA?e�(�D��@YU=�I�>>a	?�?>��0��1��C�����>�8�?R�?fDM=%�W�$G��-e?NE<�F�Ze޻�.�=�̥= ==m���.I>�ג> ���?�Kܽ�5>W�>�[&�����^��h�<�>^>[Խ����Uք?�z\��f�M�/��T���R>�T?w3�>V�=��,?�5H��}Ͽŷ\��"a?�/�?���?��(?aͿ��ؚ>��ܾ�M?�E6?m��>�c&���t��~�=����i��*���#V���=���>W�>c�,�#��?�O��t��G��=�:�,�ѿ� ��$��Y<�+;��2ʽ�ͽ����L��,ߐ�K;�M^޽l+�=���=�N>��v>�<>qz6>�;R?4�?w��>U�=0�����Oپ;�_���h�%I��跾oo�#A���U��;��k��!�
������r��"�=��X�~���F� �4�X�TnS��?wgH>�W�P���7��NԾ�~��J�$��(⽣���[�h�m��Ѧ?¿H?$D��:�W���侸�`���=`�l?w�*���ܾ �	���<�皽���=[��>���=�̾��H��T�C,?�?�uþ��g�=rG�^�<G�.?:��>x����>�|0?˰��+߽���=py�=�<y>{_�>�h>���3��}?2�O?�@����Ѿ�4:>�ԣ��R����=�">E��@w�#��>��g����$%�=\�O��s=��V? ��>�*����B��?�=?=� x?�?�"�>X�j?n�B?���<6���3T���Q�p=��W?M�i?Į	>�䁽�о��X�5?�e?j�O>X[g����{.��)���?��n?ʖ?������|�pΒ�ub��:6?���?/�?�����J�ɾ�k��쮘>�*?�>ֵ:�5r?�;,?ez��x���3�˿���W�?jg@6U�?۷/��iO=�PX�k��>|�!?�gt����G�����L��1���q�>�9�\�i��bV��4���S�?��?��?�п���;�D�%>p��c��?�U�?�_��5���f�'�p/E��"�Ad���7>G�ٽZ^�l���"��ξ�(�d���h��>��@�}�����>�g�����jOĿ��������#��\^�>��>B4Q�zT��qZf�(}��$�T	!��X��K�>��>д�� ���q�{��q;��A���>j�b
�>6�S�M%��/���Jo5<��>A��>��>&��/佾�ę?Bc���?οu������e�X?Wh�?Ho�? p?�w9<R�v���{�h�./G?��s?Z?e%�y6]�w�7�W�i?J��a�_��4�+CF��cW>F2?�X�>!..���W=��>�f�> >(Z-�{ÿ�����6��?�Z�??��6��>0�?�,?����ᙿ�f����%��t<�=?��.>&���lE�w�<�����zj?/!0?���j�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?߃�>|߄?A�=� �>���=ҕ��k���D">���=KF��-?S�L?ܓ�>���=�G8���.��F��R��4�	bC����>��a?��K?be>����t'��} ���ɽN2�#]����<���)�8�ҽߠ4>�B>�>�HG�pԾ�V?_��,�ȿC���<�:�z�?a�7>+@?������9<��p?bB0><����������:�?��?��?�Qʾ���g�����>P>�2Ƚ���6���}6�>%�U?��I���,+`��Fj>u�?Ax@!��?����	?�'��A�m���l�3���쐌����=7�6?��߾��>�� ?p�>�at�����z�	1�>���?G��?��>�rX?��U����|�=�8>e[j?�/?�3�C��.��>�e?��I�&	x�R�G��	V?"@�_@<hv?j��D�߿3��qh����žas�=uD�<� �=I*ܽ���=���<�C=Z�=�t@>�d�>1�>��>�=>%�	>��=�{��į'�2졿�i��7�J��$�/���!�LR�ts}��y��oȜ�QGϾ��۽��ҽ^�U��"P�E�J�����=acY?�`?)�w?HX?>ӭ�R��=���6��=X�����=m `>��&?��V?'()?�`�=�a����_�H���M���݆h�*=�>?0o>U�>���>���>���#�J>e&�>�6>�R>��<���=8��=T�*> ��>~��>�r>h��%�"> ü�6��� @Y������,=,�?Zh��?L�~���+���$nھk<>�?�(@=㜄�ݑ׿�j����P?�4o�h� �J��HV���v,?l�a?ڽ+=t~־�%>��>���<�>˽�]<�n��:I���#�!k>��?�2>o�v>�F��D���U�P��I�>A�(?�.��ǔ$���|�f�H���˾��4>��>W�H�iV � ���Kl���D�S�x=c\.?oG�>�����T��?��/�>䍂>kc�=Ts�=is>뽼�>�G��iH�u3=�X >7�>8X?~->4+�=�͡>n�����L��}�>5D>�{&>h�=?�v#?��wE���t��x�1�!wq>���>?�>;�
>baJ��=#k�>^�i>[#ۼ%���r�T�8��+`>�O��V+^���G��=�����=	�=����=��Z2=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>��B�b��f^������
^���܋>��?eZ��-=�g8����>3B?��̾Ѐ����Ŀ�#j�D�>�1�?0{�?�S��[���?�Ъ�>N4�?5?l?o��>P���[d��'>9�!?�P�?�G?3JӾ&lB�  ?O��?Ud~?�&_>8��?�|e?�Y�>`���(�U�j���끿��,=�d��6A�>\I�=�ͨ���F�Bd���H��F�Y�Zj���h>i�<�|�>���y���T�=
���ݘ�P�ҽ���>���>���>��>�E�>#?��>0��=����F�U���K?�]�?;��?l����<�,�=sx\��*?y�6?3�A�jQ;?�>��[?�?3
[?�3�>	&�%���B������	9�<�1K>"\�>UT�>X�e�P�W>��оE�6�Ɯ�>j�>Y����׾����׻|*�>c�!?*J�>��=QN ?,�#?��e>��>�xD����w�E��x�>v��>��?�$|?��?K���xr1�Cߒ��Y���8Z��YQ>JNy?�?o��>�;���E��N���Ov��m��g�?
Mg?ݽ`?lm�?�J9?F�A?��]>�#�K�Ѿ�ڔ�F�y>��!?��s�A��Q&�5�S�?�U?��>������ս�M׼����m��8�?;\?�0&?B��N%a���¾-�<R�!���N�Y�;E��>�}>i`��X��=;>�ΰ=�5m�N$6�,Jd<I�=���>���=w37��M���T?V��X��(W>�~a��Bg�g	�>�>K��`�?��W�N.��g¿HO����<ڭ?���?�j�??w�u�{��@?���?o��>��?�L��溾��оk5���g�����|��>��!?��^�a���Ո��krſ7����᳾Ϳ%���?\�>MF?]�	?�//>�í>6���)�!���+H�"R�
� �Cw:��Z!�d�◾Ǽ�����bӿ��n����>�[�?��>Z�?[,G>%��>��>�|��я}>hom>L�k>� �>��[>�$%>ܦ�=�6�l�Ͻn�Q?P׾�C�'�5��᭲���A?̮c?�|�>�P{�6F�� ��;�?s�?r��?:�o>
ph�XM+�(??���>�p��I
?�pJ=u���DԠ<$���Z���x�q�m�>)�Խ�x7��L��'g���?9>?@c��e˾�kֽN���Mg=� �?�|'?�(��5Z�w�x�8�U�
LS�N
O�+uQ��L��<��5v��k���z������
= �.Y=#?�5�?��&�߾#D��]cr���A�?;>>���>�X�>��>N�G>�t
�p�%���V�S&���k�!��>Co?�>��w?�??s�.?{�{?4*?5� ?+�b���h?z)n>�{�>�B?��5?��(?�<?�R?��?�>�Mb��]�����l?�,?K�&?~�>t�>��!�8�ݽ����=����_K<
��=��=�ʽ.�ȽCŚ�+�M>X�?(@��]
b�����"�J?�	?׬����)���j�W�q��N>us?�;�>�7A�QT����0�(�?{�?~��< P�=���=oo=n�l�W���=��*=��������J�Z߼�=���XW�[�?=ӵ�=oW:��SϽ��+��v�>�?���>�U�>4C���� �R��.j�=��X>��R>_>�Hپy���$����g�(:y>�r�?v�?��f=I�=��=7����U�����������<֚?xZ#?�QT?"��?3�=?�b#?��>U,�xJ���Z��k����?O�>so�>��������h9�Hn�>_ǀ>҂^� нى8�ᵋ�2����t =�^��E|�����;;���n>s
��^��v�?4C�?��K=�,U�w�������J�?Q��>�_�>�l�>�k2��[�Q��XN>�C?�<?-��>o�O?�-z?6�\?��Q>��:��֮�S>����#��!>�xA?�9�?࿍?"�u?�@�>��>՝,�ٺ�T���P�%�� ｂ���):=`�Y>���>���>C&�>��=�p��>���N�:�)�=�p>YX�>�̨>^��>Wm`>C<��G?�o�>����v�ޔ���n���p<��nu?2��?2}+?��=�x��E�C����x�> [�?"�?�*?�1T���=�lռ魶�9r�Ѷ�>�3�>��>ִ�=˭J=}�>���>x�>u��Zv��X8��"M�\?pWF?ED�=�oſ �o�Ðt���9�<���gk�%����Z��k�=.���̳������b�:�������q���{��Ku�Z��>hǂ=���=���=1�<BL��/�<cfC=�C<��)=�H���K<^�@�¢��ჽ$Zs�i�{<�^=�Իn�˾��}?y�I?V&,?�cE?=ts>�>�����>��X�?%[X>��w�;q���64�8����4���־Y	ܾ�Nd����Se	>�A��P>9>��=�*�<p �=I�e=xʇ=Q ;=6=J�=vc�=b�=��=��>_t>B��?��y��h��pb=��~ �DV8?Tߦ>l��=�oھ�0J?!*>6q��#�ÿ�H(��|?]��?pJ�?%o?{Oj�Mڣ>�C��Ƕ���%>N0����>LFb=���0i�>V�^>S���'����U� ��?�@]�A?����0Dǿ���>�6>v>yS�ٟ1�T3_�� a�G�W�(Z!?*;�d̾��>#=�=p�ݾ�ƾ\?'=��3>r�W=����9[��=�Sw�y�>=.Pp=�>��A>�,�=�&����=_�M=xY�=k�R>��n�T:���8�l�3=���=�c>��(>4��>�x?�/0?��c?�.�>Am���ξq�����>���=8&�>��=��B>���>��7?�vD?�K?f�>�=�k�>��>�I,���m��㾢���|�<�v�?���?Z"�>�WT<7�A��]��k>�>�Ž�6?�`1?�	?��>�U����9Y&���.�$���{4��+=�mr��QU�M���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=$�����<�vż�����u&�:�+�1�����;r��;B�]<_��;!&�=��?D��>>��>��>���-,>����k2�x��<Pm��C=�h�u�L����&�ѽ4�i>'�b>�o�T����>�g>�>g,�?��v?�7�<N\6�F�k�pEƿ��-�����n�<�/�>iϽ�X��#x�@�J�S�����>ϒ�>v�u>�K�=�.���F������4�6�+��~�>{ʬ��/�=���`Qx��T���Q���4o��O��T?�����b�=+�?�%Y?禈?B�h>���?%�M>��?�g�>8���	��lvH�ă?�6?���>��ž�@�w����Ľ���>w��IT�E~���S��������>,^���F����8�
e��<\��y/P����С>�W[?���?��i�E�d��/.�� ���<0�?�v?�ev>�"�>QF?��#����P����=R�A?��?���?�>M��=k*ҽ���>�
?Q}�?�5�?2�s??�5��/�>ߍ;I�>m\��&��=z">�T�=3��=��?��?�B	?�X��ȣ	��:�a��#_�V��<�ї=�`�>���>��p>v[�=��~=lM�=��Y>���>�׍> le>�$�>ߘ�>XԠ�eb	�k�8?}�f>-��>�d?i�4>*��>�񿽖�����=~Q����U�A����<	d`=��<*~=��h���>�ۿ$!�?��>�� �	P-?!�	�v�T=	�=�x�>j�^��p>]�>M�m>a�[>��r>j_�<ߔ!>�M�>��޾4�>M�;�3�I�nlR�9�!�k�9���=�����W7�ʘ%�Y�a�ɉ.�G���S��(�]��|��MW���=U�z?���1�7��i+�X���L�>�qi>t��>�|���6T��h+>\/�>��>�`񾘧����������?�b�?�c>4�>��W?��?��1�J�4��Z�4cu�67A�3e�Yf`��э�x����
�����V_?0�x?O[A?�T�<%z>ƶ�?&��ݏ�0�>e/��:;�ޑ9=�Y�>?��H�a�o?Ӿ׳þS	��5E>�1o?�?)?��U���½Ь̽�b_?�eN?J��?Af?�d$?��\>��o?�iR��7?�*?V?�	Y?��X?���>j+;>*g�T6 ����xm�� ��p��pB+�1Mn=w�=bg���&�N�<���&8�ʾI��+��1`�:�ȡ=3=�{�=4��=>:�>O%^?�>�6�>�9?�����6�tҩ��3.?��<{�y�d=������i�󾃴>G�i?���?�Y?H�U>�B���L�U>J�>��4>:Ub>�I�>dܽ�F���=V�	>��>�j�=/,����X	��$��k
�<�?>���>NG|>4����o'>z���5�y�{�d>d�Q�麾�8T�H�G�5�1�v�I1�>�K?��?�=�6��Q��24f�n+)?,a<?unM?��?��=� ܾ�9�
�J��d�a�>�"�<f��n�������:�wJ�:��s>��
���.b>F���޾�n�;�I��羼�K=�A�?@V=x5���վn�~��C�=B�	>����� �����ɪ�CKJ?�wl=Bҥ��bV�@���<E>̘>�T�>�U:��]x�@�@�����s��=���>�`:>%���)�d�G�m��>��Z?� �?2�?-�=����h���
�˃C�ɂK>��%>h��>(�&?b��>�;>��ؾ.!"�
c��J�G�>E�>�D�>��-�� 5�z� ���D�Q��h.�.�?Yd�=C��>GQ?"�>�`I?�"?W��>g�>N8���ʾ.&?m��?���=>Խf�T�G�8��F�ä�>��)?��B�j��>i�?!�?��&?L�Q?ѡ?��>Ƕ ��J@�$|�>�C�>��W�1P��G�_>��J?��>x6Y?"ǃ?��=>;�5��㢾�
�����=tE>��2?h0#?��?I��>b��>������=���>hc?�.�?R�o?�p�=6�?L42>,��>��=A��>���>�?VO?��s?��J?U��>m̍<�=��G���r��OO�Gi�;>�I<?�y=�M��	t��[�7�<Y��;F���������UD�-󐼸��;w��>_D�>LF��&�J>kO��Ľm�>$���.+�����΂��~�=횃>�B�>^�4>M ��;�I=���>���>o*���/?�a�>W~�>�P�iGR��g��?�{�?��\?�X�>I�N���������}:>�v}?F�?����>��b?��]?eg�i=���þ׷b����Z�O?�
?a�G���>��~?e�q?G��>��e�":n�0��!Db��j��϶=.r�>0X� �d��?�>K�7?�M�>��b>'�=�t۾q�w�vq��B?��?�?���?8+*>|�n�V4�|I��:���[^?���>~���ӷ"?����aϾ����������N����Ы�_Q��� ��XV$�~ۃ���ؽ��=>�?�Cs?V�p?X�_?/� ��4d�	S^�����vV�<d��-�q�E�N�D��C���n��y������)��]xJ=��m���B��i�?�3"?:�i=�O�>u
��Vٵ����G��>�84�0���oZy=�u��>�.�=�1l�Hx��j����P-?��>cĵ>�O?":d��S��NE��d�,'�-<��Q�>I[�=�$? ܵ�x����'��R����x���<��g>�m?� `?׸�?;�O�RNU��m������'׽���#W>�I>��>�,��'��d[4�{NI���r�K��������a���=�&<?w�I>*��>�)�?Y?��辻3�}L �����<}C?O�B?"�>���=�8]��<�`��>�n?5��>��>B���;�)��%z��4�����>��>�A�>yp>k��� a�l���S�����8�O,�=�<b?׃��&Z���>�uT?�aP�m�R<�/�>��Q��;��z������/>��?v��=l[0>��ľ^�A|��)���7)?�l?�쒾nX*�[v|>�"?�>J��>�D�?�>ڙ¾s���K�?(v^?�J?�8A?���>�5 =:.��"�ǽ
�&��%*=:��>m	[>�j=1&�=T��[[������C=p�=c�Ҽ�!���w<�7����e<�P�<��3>�(ۿ�yJ��{ܾ~e���	��'��!��a�̽R�нV� �4�y��^{;��p��p����&�+�H�IZ����f�	�?/��?��������ų��Tq�	��K>ˇ�Bœ�9�ɾ!���]����e^����+/���D�>a��˸]�8Z?���3�ƿWE��e%�[Z$?-�?��+?}α�J%C�7N�!j�>���<ާX��r�
�����ȿ|7��IKx?���>��׾��D���?0I�>��>��=@U�3�l��`{��t�>n�K?&�>�B��@����w���Z::��?�$@v3A?��*����ɸ=[��>R�?�[;>��-�ns�2��}y�>���?��?�h5=��V�����e?o��<�C�J�����=���=(�3=����{?>���>[����6�*2߽>�5>�e�>BO�J�E�e�5=��|>R�ڽ�)½Lц?��<��1����`�{T>
U.?)u�>�`>��>��O�ɿ������F?#	@zZ�?ĕS?EZȾ�>�6׾��J?�['?��>�7&��̙�Q��<�׼*��	��\����C^�>3`�=��������B�v�<k��>�F�� ƿ�#��[���=�c<}'��H]�g���jq�X����[�iI̽�T�<���=,Z>Q�s>*<>Y�L>#fQ?J2m?X��>���=�pl��G���پ��3��� ��r���:������ྒྷ�����w�����s���\D��e=wP�VЕ�N.6���Y�Z�B�G1?�?w>�ڿ���W�k��<�O��;뉾2y�Pb��D�Ǿ��;���g�:�?r�F?]�����n�}���<cug���.?�}޽3	����L�>�`��=��f>��J�\�����C��B�ѡ.?� ?��ҋ��0=>���9�k=w&?�F?�m9<D��>��#?��&�R� �eV>�E3>`��>���>��=+��E%�f�?:T?|��xܟ�ښ>t����a��ʒ=�>a�!�Ҽ�Z?M>��<Gov�x��<�j��H:g<��A?$D�=J�
���>�&�о�G�<ue>AU�?�H���&)?�ǖ?.�T>'�>���h�^P����=;k?��?��>�{���E ���0K?V#�?���>tо��۾��U�����]
1?��V?�:?J{7��R���&���2?�>]?'<��f��YC��#������>Y��>�_�>8���:�>p?]�b����:H��Ī7�*�?@��?�*ɽ�	}���c>-*�>5�
?\M���'�x�C�[ǀ���m�>U붾l���WD\��e��?N?��?��$?|������if�=���
�?{��?8�m��*������(J�v��&���s�=�4�v�<Xy���I$�!㶾s�������m݌>s�@�僾��>�dn�k{�ۣ̿Sq�fM��oq��q�>L��>2<H@���o�9o{���1�����mL�/��>�>�Õ�������{���:�A�����>0���"�>�vR�������V�<���>=�>E��>dӪ��M�����?���5�Ϳ����%	���X?��?f�?�t?#�V<�5w��)}�
P��F?4t?�HZ?��&�ɀ\�J$<�Yj?k���_`�5�p�D���f>�1?���>!�*�+�l=��>#z�>Cx>�.�dÿ��������?���?�����>Qz�?��+?��OS��CŤ���(�D$�;��>?�
3>����K�#���=���B�?O�6?�[	�%!�]�_?+�a�M�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?е�� #�f6%?�>d����8Ǿ��<���>�(�>*N>dH_���u>����:�i	>���?�~�?Qj?���������U>
�}?���>��?P\d>�@?�>9�������\q>���=�D3���?��P?���>rw�=��"���3���S�1\�:���2XB�� S>xoV?`"@?,R`>����8��̱ ��U��hGe�k������x�S�=��;>��[>IU�=���`��
?E� �g�ɿP_���#3���e?��l�9�`>�fJ�����5�S��`q?y�>Ҏ��0���!y��Mm�-�?���?{b?n�����>R��=�-�>�Ϫ>�t<,�<>؄ξ�f�>Q�N?� ��-:�h�:�ʸl>F�?��?���?��k�5	?��&����}����=�*�j�=�r6?˸�N�x>@��>#��=�lt�=����r�
�>�T�?��?���>1�j?�%l�
A�jI=��>��g?rV?�vx����7%B>�x?4��kY�� ��c)c?�@��@Cv\?W��??߿�J���߯���Ǿ�<=�!�=A6~>E2����s�ᐙ��׽�$<tr=$��>�w>�L	>��=��*>V^=%�����a���=F���)F�I��� �Ã���;��r���O$��$;��˾���7�n�{���y��M�S�߽b��=�3q?�1_?{a?}'?�2�4��<�=�w�>2��|�i����>�(?CY?Z�9?���=HG��&�g��Iw��M��u�����>��=<��>)��>�&�>���=\
>���=���=9��<����i�h���<�m>��>��?���>�A<>b�>-ϴ�!2���h��
w��̽� �?B���-�J��1��S9��~���8k�=�a.?#{>���?п7����2H?t���*���+���>��0?�cW?�>����T��9>��J�j� `>�- �W�l��)�$Q>�l?��f>�u>��3�je8�^�P��|��>j|>�36?`鶾D9���u���H��cݾHM>�ľ>�D��k�{�����Tvi�z�{=]x:?ք?�6���ⰾl�u�VC���PR>m:\>U=�i�=�XM>bc��ƽlH��g.=(��=̮^>/W�>H˓>17E<��>Vg辰%�#U�>���=Zp�>�D)?{�5?�#=X��R#��q��j�>��?	��>���<�F����<&�>>��>�z�<#����I<�(H�`g�>R�=�Ci�<�����K���4>�A�>���=!���[0��˖~?r~���㈿)�j]��)mD?n*?&�=�0F<ׅ"�����,E��)�?8�@8k�?σ	�G�V���?2A�?S��U��=~�><ի>Dξ��L���?�ƽ����^�	�� #��Q�?�
�?a�/��ȋ�}l��;>�]%?��Ӿ�D�>�J��?��������n�H:�=�Y�>\�!?�y��M%��4����?>�>����a����ȿ�Uw�;��>���?�/�?��b�QZ����3�,r?��?lM??��>��ؾTo��.�>��@?<�K?P��>wy�=��?��?[��?�]I>�P�?�؀?���>!M:=(fQ���E�q�v �G�_��DF><�=�y���^��d~�]���ϷZ�d��*�?>�{=��>*7�(i����=�"ҽ9(Z�������>��J>[�a>Q?���>�[�> ;�>�`��!"/�B����Y���K?���?3���1n��X�<h��=X�^�&?�I4?i[�P�Ͼ�֨>��\?Z?�[?�c�>��$>��	迿�}�����<��K>�2�>\H�>K"��JK>E�ԾI4D��o�>WΗ>Y���@ھv-��>��$C�>�e!?h��>ծ=8� ?)�#?�j>)*�>_E�2:����E����>d��>�G?��~?��?^ѹ��[3����v桿��[�M9N>9�x?>U?�ʕ>J������mxE��LI�@�R��?�tg?VR�.?�2�?�??��A?H(f>Ό��ؾ߭����>]"?�j��[A��&��'�k�?�G?�l�>T����ӽ��ǼC��������?��\?�&?�����`�uþ��<�-%�����;�M��a>U>f��5L�=�x>��=�o��q7�>
�<ʼ=�t�>@��=P�8�_'��Z+?S\�=T�F���>��r�̪N�(r>%->ߴ��uC?�RC�oц�l���X������}L�?g��?�8�?��a|m�Y�J?�W�?a�>?� �>�Y��9�s{�¯�f<:=M��؎�=D�?4>�=���z���ճ��'���(���K�x?�6�>��?�}?��=aP�>5)��*���4ȾO��ʯb��2�Pq6�T��G������|�X����J��w0�>�贽T�>M�?�� >O��>�	�>�-���b>��>I'p>=�>a�=.�=��>u�=�v���Q?�Ħ��}!� ÷������E?JtX?(��>f>罃��N��J�?�t�?=�?d�>�o�22�h�>7�?[懾�?�U�=��鼽J-��_����V=)�Rr>8�G>G��<��/�\49��ީ���?�?F�=ִ��B@E� G��_(�=Ҋ?�T1?C��`�Y�V�p��\?�G`�%�����\��=ɾW1��q��E��8�}��z�M6!�i�=�7$?��?1���澐����.q�jWB�N�P>L7�>��|>OՒ>s�x>����`<��X��01�is��M�>#s?o�>��I?E�;?=jP?�BL?e��>�r�>:����>�T�;���>��>�9?��-?00?po?k+?�c>��������xؾ@�?�?�??��?U�?����g�½}K��1~j�Xcy����.o�=���<�2ֽ��r���U=�T>�@??��Ӿ8?3�Y�w����>ڻS?(|�>�?>�6��ӽi>$�>̕?M\F?\(���c���*��?M�?��ϼ�\�<	�=��f>,`����=�zĽQM)�Cߓ=�n6��5����=�5컝3�=�U==�����1<�ؽrk6=le�>�?q�>pU�=����2�����Ҍ�>3l�=!��>�r�>N5�=3m�����b!a�g%�>�d�?�<�?0����C�<�5>n�-���پ����&}���O+>�Z'?	��>|@s?`Ԥ?�+�>��*?
[4>_RȾ�钿PM�������b�>w!,?	��>�����ʾ��ԉ3�۝?g[?�<a����;)�ސ¾��Խر>�[/�g/~����<D��셻���=��5��?쿝?_A�U�6��x�ۿ���[��z�C?"�>Y�>��>V�)�|�g�r%��1;>���>gR?�A�>b�s?�k~?�]?S��>~xK������L���/7>'T>}� ?=�?f�?�Ć?a��>�ƺ=�z�� ����"L7��d�cHq�p��32>R��>�?z��>�C�=��4�6���XN�Կz���m>��>���>���>��>��H=`�??���>�@����ྃWξOuh���=,JT?"Q�?I%?��=�� �>9���w�>��?=+�?7,?��x��A>o��������f&���>��>Iќ>:��<�h=-9g>���>��>�_����;~�+�>[d?n�:?��u=�sҿ�&���[���1�������[���M?�����(N'�~�=)Sƾ���쒾ShJ��ޣ���������硾	兾�?P����=��$>�{W= ������<��>��1=��>,\��VH=�@�=��6O%��;�=���<���<�A=�˾�}?ypI?ƪ+?�D?��w>ż>�)1�+o�>Ē��,?�GU>�V�����?:�[]���B��x9پv�׾��d�����Qt	>�zI��>�"4>FK�=p%�<�!�=lt=͝�=-ߺ�4=��=��=0ʪ=;��=�>c!>@w?\6C�n y��W�2�?�ZhA?���>��}���X?���>��W���ſWr$�U0�?"@���?c+?���N]�>�4��ɽ�=����bP�=ۉ}>ɴ�Z]=�]@>dq�=4����i����پD��?jM
@�Z?�nq�um��i�=��7>,,
>�P�$�1�&�c��m��D[���'?_:�<������>3 �=�ܾ�˾#y�<K13>���=�l�Z���=����	N<=t�6=�E�>{�H>-#�=9?���}�=o=�i�=��>>ۗ�;��ռs�I��=�{�=�\>��">ƕ�>��?�Q-?c?��>Xh�Z�þpj¾���>���=mA�>�P�=��@>Ŀ�>Wg5?��B?d�L?zn�>�!o=Ì�>�S�>d�,��th��߾�8����=3�?���?���>��U<S5��7��T>�0���?�K4?�?f�>f��I��|4�������4M=e�M>��	X��DZ=w��h����>�5�>^Z>�j>�Q6=?֙=)�==1�>���=XI2��m�W�=���= Y½6�*>������<��j=����U�qӽ]s)=�5�=Q�=��~=���=�D�=��?3�>Ek�>x�">q�澖��><|޾�S��5o>��}�=`�<]v��)|��`�x.�N	>n��<\�?�����X?i�>��=�'�?V�s?��=H�-�U)z�?	��7)�ʽ\X�<��>�[��lO�a���I������>���>�3�>31m>��+��5?�YYw=��ᾔS5���>���Y���3q�0���🿑i�/���D?�A����=�
~?�I?$؏?V|�>����ؾ��0>���N�=<���&q�	���N ?'?��>m!�$�D��G̾���ܷ>�BI���O������0�{���ɷ�$��>������оz#3�Eg�������B��Mr����>߶O?"�?i:b�JW���TO�����'��5q?�|g? �>�K?�@?�$��sx��r��Fy�=9�n?a��?�=�?V>Ͻ=�紽d�>b"	?鳖?ݵ�?�s?H�?����>�Ԋ;�� >܋���W�=ܚ>�f�=��=�s?�
?�
?�N����	����A��^�ai�<+�=�|�>t�>��r>���=*�g=�K�=i\>�>���>�$e>��>�7�>v�ȾER۾k	R?GN2>�?��
?���>B>~�����*>blA�Gc���b��h����<��g=�
�����E�q��>lۿY�?D�=m!Ӿ�c%?�o�_Y�;��#�;��>v��<c̚>�$�>�p\>[N�>��>��=�u.>*�n>�v >�)� �X��l��*��˾���üx ٽ�����)��q�X :���o�{_�f��L}���]��Ta=���?�劽c_��
�骰�c~%?�Z�>�W�>�C���Ӊ��V�=�B?I:C>���▿�o��B��DB�?Q@@c>�>�zX?�?��.��W6��~Z��et�H�A��d��`����e󀿈�
�����i_??x?N�@?ف�<�?z>}�??�&�ȋ��aP�>^�/�I_;�;�:=���>�|���c���Ѿ�W¾���}BD>��m?�Ӄ?�?�wT�G�l���.>%`;?�?1?��t?�l0?��9?N��
%?�0>�0?)5?�4?�s/?��?�-3>��=�m���=�ɒ������ͽ�̽�a��u9=
��=W& ;�	�;"=�X�<������r��9�s���^�<
�<=Y��=W��=w��>�n]?�t�>�~�>f�6?֪��8�!���)�.?QbK=.���R��}��q��� >�Zj?ݫ?xfZ?��b>X�@���C�t�>I�>50'>.�\>�G�>�j��IG�^؊=�2>X�>��=�4C��ծ	��0����<|�>���>0�>F�#���T>�4��j������>��t�"ȾV���A���;�
%���ǩ>�JR?��%?ʑ�=S�����e�m��3,?
I?�pN?�Y�?h�=ȃ��=B��O�9���:-�>�!�<����C��]ۢ��C����9�">T
��1�����c>��� �m�c�I�-�辱�U=�.���=���w+޾�w����=W�>�ſ�wE!�1���i��+�K?��m=����+W�/����>��>��>�
U���]�@W@�4+���`�=g&�>z�A>b�p�G����F�����E�>�sP?��c?�p�?�����m����k�5�6�����W�,<P)?��>Uq?#^�>J;>T����O��|�T��U��n�>��?�mJ�b	h��|j�A]�t�E����={[)?���=�f?�BQ?�?�xC?�K�>�8�>�K>��z����lW+?NP�?�
�='	��c�ʽ�\1�mP\�ŏ>RB?�!�d+�>�:?��?<H?c�K?�	?���=�Q� �N����>ɻ�>��G��϶�|��=�v?� ?dv}?Bb�?��,>}X#�������
=M1>6/?3h&?vM??Ɠ�>f��>:��+>O�>�d?��?�pm?��W>�e?��=
{�>���=���>�?l�*?��J?�o_?�4?ߙ�>t��=�͔��U%��	���c���f��'�����=���;�Wa��rT=r�%>�<�;�<H�=l耽Рk�]�=�_G����>�O�>�𚾜g>�˾+����G2>Fָ;����+��hB�">Ń�>=�>��i>A�]8=���>ʾ�>`� �!?��?�?� =�wf�w?�815��S�>��9?=��=�LW����wg�R��<7�i?]�_?�{ �U���b?x�]?c^��=���þ@�b�ۓ龤�O?��
?.�G�h��>��~? �q?���>��e��7n����Db��j����=�o�>�R���d��?�>��7?OR�>]�b>��=u۾*�w�2p���?��?���?��?s$*>��n�3�Od��=[���^?���>�_�"?�q��SϾ����q'����ᾙ@��I��}x���A���$�bჾ-'׽6�=�?�s?�/q?f�_?p� �>�c�-^�0���V�>�~���E��D�ōC���n�'w��0�����	�J=V�B�qt�L��?�1?�{��~��>��Ⱦ��L�%��4'	>�D�LI��t�xV�,i�=#�==��u�q,2�R#¾�)"?ߟ>7�>�bB?�%��ۻ4���0�6[���8�ν->SI�>� A>%�.?!���0����F��-�ؾ�ih��>���>k_?�xN?8v?Q���4�O�����4�q� k��uZ�>���=Q\�>����3������I�1�y�v���W��@����>ǖ?���>/�>��?GU�>�4��nN��P}���p�]��<KM?xT?N#?L�>��T��&Q��@�>�l?�Y�>�Š>B6��8� ���z��ný��>a��>��>�xo>�&�1�Z��Ď��	���8�<�=�Eh?x;���\����>�IR?g�<��<�{�>5h�����h�a!�.x>j?�?�=�f7>����1�
���z�����i(?tu?ڂ����%��L�>j4$?z��>�W�>,�?n �>"A��y��;�?�^?��I?m�>?V��>u1=s�Խʋ潌2&��ks=0��>���>vә=�f�=�>�ES��\��Q�f=���=n�'�PH׽0�o;�d�����<�(=��?>�j�؂]���Ҿ?4 �r���K�W�ʾA��D�B��m����Ѿ?���>~�.��st���,]�Ճ�����qx��^�?��@���	���Ⓙ��]�.* �� o>V_%�N$5�7/"��{Ǿ,举�{ؾ�ؾ4,-�=Z�p��lT��?�kr���ȿ���t
��?��$?Dm<?�������4G��=I=��W<r��q������ƿ��־esa?���>�jԾ�*A=���>��g>�->f�=f.��Y��!.��A�>�x+?��>�"���Cҿ֞����b�&�?��@�mA?e�(�D��@YU=�I�>>a	?�?>��0��1��C�����>�8�?R�?fDM=%�W�$G��-e?NE<�F�Ze޻�.�=�̥= ==m���.I>�ג> ���?�Kܽ�5>W�>�[&�����^��h�<�>^>[Խ����Uք?�z\��f�M�/��T���R>�T?w3�>V�=��,?�5H��}Ͽŷ\��"a?�/�?���?��(?aͿ��ؚ>��ܾ�M?�E6?m��>�c&���t��~�=����i��*���#V���=���>W�>c�,�#��?�O��t��G��=�:�,�ѿ� ��$��Y<�+;��2ʽ�ͽ����L��,ߐ�K;�M^޽l+�=���=�N>��v>�<>qz6>�;R?4�?w��>U�=0�����Oپ;�_���h�%I��跾oo�#A���U��;��k��!�
������r��"�=��X�~���F� �4�X�TnS��?wgH>�W�P���7��NԾ�~��J�$��(⽣���[�h�m��Ѧ?¿H?$D��:�W���侸�`���=`�l?w�*���ܾ �	���<�皽���=[��>���=�̾��H��T�C,?�?�uþ��g�=rG�^�<G�.?:��>x����>�|0?˰��+߽���=py�=�<y>{_�>�h>���3��}?2�O?�@����Ѿ�4:>�ԣ��R����=�">E��@w�#��>��g����$%�=\�O��s=��V? ��>�*����B��?�=?=� x?�?�"�>X�j?n�B?���<6���3T���Q�p=��W?M�i?Į	>�䁽�о��X�5?�e?j�O>X[g����{.��)���?��n?ʖ?������|�pΒ�ub��:6?���?/�?�����J�ɾ�k��쮘>�*?�>ֵ:�5r?�;,?ez��x���3�˿���W�?jg@6U�?۷/��iO=�PX�k��>|�!?�gt����G�����L��1���q�>�9�\�i��bV��4���S�?��?��?�п���;�D�%>p��c��?�U�?�_��5���f�'�p/E��"�Ad���7>G�ٽZ^�l���"��ξ�(�d���h��>��@�}�����>�g�����jOĿ��������#��\^�>��>B4Q�zT��qZf�(}��$�T	!��X��K�>��>д�� ���q�{��q;��A���>j�b
�>6�S�M%��/���Jo5<��>A��>��>&��/佾�ę?Bc���?οu������e�X?Wh�?Ho�? p?�w9<R�v���{�h�./G?��s?Z?e%�y6]�w�7�W�i?J��a�_��4�+CF��cW>F2?�X�>!..���W=��>�f�> >(Z-�{ÿ�����6��?�Z�??��6��>0�?�,?����ᙿ�f����%��t<�=?��.>&���lE�w�<�����zj?/!0?���j�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?߃�>|߄?A�=� �>���=ҕ��k���D">���=KF��-?S�L?ܓ�>���=�G8���.��F��R��4�	bC����>��a?��K?be>����t'��} ���ɽN2�#]����<���)�8�ҽߠ4>�B>�>�HG�pԾ�V?_��,�ȿC���<�:�z�?a�7>+@?������9<��p?bB0><����������:�?��?��?�Qʾ���g�����>P>�2Ƚ���6���}6�>%�U?��I���,+`��Fj>u�?Ax@!��?����	?�'��A�m���l�3���쐌����=7�6?��߾��>�� ?p�>�at�����z�	1�>���?G��?��>�rX?��U����|�=�8>e[j?�/?�3�C��.��>�e?��I�&	x�R�G��	V?"@�_@<hv?j��D�߿3��qh����žas�=uD�<� �=I*ܽ���=���<�C=Z�=�t@>�d�>1�>��>�=>%�	>��=�{��į'�2졿�i��7�J��$�/���!�LR�ts}��y��oȜ�QGϾ��۽��ҽ^�U��"P�E�J�����=acY?�`?)�w?HX?>ӭ�R��=���6��=X�����=m `>��&?��V?'()?�`�=�a����_�H���M���݆h�*=�>?0o>U�>���>���>���#�J>e&�>�6>�R>��<���=8��=T�*> ��>~��>�r>h��%�"> ü�6��� @Y������,=,�?Zh��?L�~���+���$nھk<>�?�(@=㜄�ݑ׿�j����P?�4o�h� �J��HV���v,?l�a?ڽ+=t~־�%>��>���<�>˽�]<�n��:I���#�!k>��?�2>o�v>�F��D���U�P��I�>A�(?�.��ǔ$���|�f�H���˾��4>��>W�H�iV � ���Kl���D�S�x=c\.?oG�>�����T��?��/�>䍂>kc�=Ts�=is>뽼�>�G��iH�u3=�X >7�>8X?~->4+�=�͡>n�����L��}�>5D>�{&>h�=?�v#?��wE���t��x�1�!wq>���>?�>;�
>baJ��=#k�>^�i>[#ۼ%���r�T�8��+`>�O��V+^���G��=�����=	�=����=��Z2=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>��B�b��f^������
^���܋>��?eZ��-=�g8����>3B?��̾Ѐ����Ŀ�#j�D�>�1�?0{�?�S��[���?�Ъ�>N4�?5?l?o��>P���[d��'>9�!?�P�?�G?3JӾ&lB�  ?O��?Ud~?�&_>8��?�|e?�Y�>`���(�U�j���끿��,=�d��6A�>\I�=�ͨ���F�Bd���H��F�Y�Zj���h>i�<�|�>���y���T�=
���ݘ�P�ҽ���>���>���>��>�E�>#?��>0��=����F�U���K?�]�?;��?l����<�,�=sx\��*?y�6?3�A�jQ;?�>��[?�?3
[?�3�>	&�%���B������	9�<�1K>"\�>UT�>X�e�P�W>��оE�6�Ɯ�>j�>Y����׾����׻|*�>c�!?*J�>��=QN ?,�#?��e>��>�xD����w�E��x�>v��>��?�$|?��?K���xr1�Cߒ��Y���8Z��YQ>JNy?�?o��>�;���E��N���Ov��m��g�?
Mg?ݽ`?lm�?�J9?F�A?��]>�#�K�Ѿ�ڔ�F�y>��!?��s�A��Q&�5�S�?�U?��>������ս�M׼����m��8�?;\?�0&?B��N%a���¾-�<R�!���N�Y�;E��>�}>i`��X��=;>�ΰ=�5m�N$6�,Jd<I�=���>���=w37��M���T?V��X��(W>�~a��Bg�g	�>�>K��`�?��W�N.��g¿HO����<ڭ?���?�j�??w�u�{��@?���?o��>��?�L��溾��оk5���g�����|��>��!?��^�a���Ո��krſ7����᳾Ϳ%���?\�>MF?]�	?�//>�í>6���)�!���+H�"R�
� �Cw:��Z!�d�◾Ǽ�����bӿ��n����>�[�?��>Z�?[,G>%��>��>�|��я}>hom>L�k>� �>��[>�$%>ܦ�=�6�l�Ͻn�Q?P׾�C�'�5��᭲���A?̮c?�|�>�P{�6F�� ��;�?s�?r��?:�o>
ph�XM+�(??���>�p��I
?�pJ=u���DԠ<$���Z���x�q�m�>)�Խ�x7��L��'g���?9>?@c��e˾�kֽN���Mg=� �?�|'?�(��5Z�w�x�8�U�
LS�N
O�+uQ��L��<��5v��k���z������
= �.Y=#?�5�?��&�߾#D��]cr���A�?;>>���>�X�>��>N�G>�t
�p�%���V�S&���k�!��>Co?�>��w?�??s�.?{�{?4*?5� ?+�b���h?z)n>�{�>�B?��5?��(?�<?�R?��?�>�Mb��]�����l?�,?K�&?~�>t�>��!�8�ݽ����=����_K<
��=��=�ʽ.�ȽCŚ�+�M>X�?(@��]
b�����"�J?�	?׬����)���j�W�q��N>us?�;�>�7A�QT����0�(�?{�?~��< P�=���=oo=n�l�W���=��*=��������J�Z߼�=���XW�[�?=ӵ�=oW:��SϽ��+��v�>�?���>�U�>4C���� �R��.j�=��X>��R>_>�Hپy���$����g�(:y>�r�?v�?��f=I�=��=7����U�����������<֚?xZ#?�QT?"��?3�=?�b#?��>U,�xJ���Z��k����?O�>so�>��������h9�Hn�>_ǀ>҂^� нى8�ᵋ�2����t =�^��E|�����;;���n>s
��^��v�?4C�?��K=�,U�w�������J�?Q��>�_�>�l�>�k2��[�Q��XN>�C?�<?-��>o�O?�-z?6�\?��Q>��:��֮�S>����#��!>�xA?�9�?࿍?"�u?�@�>��>՝,�ٺ�T���P�%�� ｂ���):=`�Y>���>���>C&�>��=�p��>���N�:�)�=�p>YX�>�̨>^��>Wm`>C<��G?�o�>����v�ޔ���n���p<��nu?2��?2}+?��=�x��E�C����x�> [�?"�?�*?�1T���=�lռ魶�9r�Ѷ�>�3�>��>ִ�=˭J=}�>���>x�>u��Zv��X8��"M�\?pWF?ED�=�oſ �o�Ðt���9�<���gk�%����Z��k�=.���̳������b�:�������q���{��Ku�Z��>hǂ=���=���=1�<BL��/�<cfC=�C<��)=�H���K<^�@�¢��ჽ$Zs�i�{<�^=�Իn�˾��}?y�I?V&,?�cE?=ts>�>�����>��X�?%[X>��w�;q���64�8����4���־Y	ܾ�Nd����Se	>�A��P>9>��=�*�<p �=I�e=xʇ=Q ;=6=J�=vc�=b�=��=��>_t>B��?��y��h��pb=��~ �DV8?Tߦ>l��=�oھ�0J?!*>6q��#�ÿ�H(��|?]��?pJ�?%o?{Oj�Mڣ>�C��Ƕ���%>N0����>LFb=���0i�>V�^>S���'����U� ��?�@]�A?����0Dǿ���>�6>v>yS�ٟ1�T3_�� a�G�W�(Z!?*;�d̾��>#=�=p�ݾ�ƾ\?'=��3>r�W=����9[��=�Sw�y�>=.Pp=�>��A>�,�=�&����=_�M=xY�=k�R>��n�T:���8�l�3=���=�c>��(>4��>�x?�/0?��c?�.�>Am���ξq�����>���=8&�>��=��B>���>��7?�vD?�K?f�>�=�k�>��>�I,���m��㾢���|�<�v�?���?Z"�>�WT<7�A��]��k>�>�Ž�6?�`1?�	?��>�U����9Y&���.�$���{4��+=�mr��QU�M���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=$�����<�vż�����u&�:�+�1�����;r��;B�]<_��;!&�=��?D��>>��>��>���-,>����k2�x��<Pm��C=�h�u�L����&�ѽ4�i>'�b>�o�T����>�g>�>g,�?��v?�7�<N\6�F�k�pEƿ��-�����n�<�/�>iϽ�X��#x�@�J�S�����>ϒ�>v�u>�K�=�.���F������4�6�+��~�>{ʬ��/�=���`Qx��T���Q���4o��O��T?�����b�=+�?�%Y?禈?B�h>���?%�M>��?�g�>8���	��lvH�ă?�6?���>��ž�@�w����Ľ���>w��IT�E~���S��������>,^���F����8�
e��<\��y/P����С>�W[?���?��i�E�d��/.�� ���<0�?�v?�ev>�"�>QF?��#����P����=R�A?��?���?�>M��=k*ҽ���>�
?Q}�?�5�?2�s??�5��/�>ߍ;I�>m\��&��=z">�T�=3��=��?��?�B	?�X��ȣ	��:�a��#_�V��<�ї=�`�>���>��p>v[�=��~=lM�=��Y>���>�׍> le>�$�>ߘ�>XԠ�eb	�k�8?}�f>-��>�d?i�4>*��>�񿽖�����=~Q����U�A����<	d`=��<*~=��h���>�ۿ$!�?��>�� �	P-?!�	�v�T=	�=�x�>j�^��p>]�>M�m>a�[>��r>j_�<ߔ!>�M�>��޾4�>M�;�3�I�nlR�9�!�k�9���=�����W7�ʘ%�Y�a�ɉ.�G���S��(�]��|��MW���=U�z?���1�7��i+�X���L�>�qi>t��>�|���6T��h+>\/�>��>�`񾘧����������?�b�?�c>4�>��W?��?��1�J�4��Z�4cu�67A�3e�Yf`��э�x����
�����V_?0�x?O[A?�T�<%z>ƶ�?&��ݏ�0�>e/��:;�ޑ9=�Y�>?��H�a�o?Ӿ׳þS	��5E>�1o?�?)?��U���½Ь̽�b_?�eN?J��?Af?�d$?��\>��o?�iR��7?�*?V?�	Y?��X?���>j+;>*g�T6 ����xm�� ��p��pB+�1Mn=w�=bg���&�N�<���&8�ʾI��+��1`�:�ȡ=3=�{�=4��=>:�>O%^?�>�6�>�9?�����6�tҩ��3.?��<{�y�d=������i�󾃴>G�i?���?�Y?H�U>�B���L�U>J�>��4>:Ub>�I�>dܽ�F���=V�	>��>�j�=/,����X	��$��k
�<�?>���>NG|>4����o'>z���5�y�{�d>d�Q�麾�8T�H�G�5�1�v�I1�>�K?��?�=�6��Q��24f�n+)?,a<?unM?��?��=� ܾ�9�
�J��d�a�>�"�<f��n�������:�wJ�:��s>��
���.b>F���޾�n�;�I��羼�K=�A�?@V=x5���վn�~��C�=B�	>����� �����ɪ�CKJ?�wl=Bҥ��bV�@���<E>̘>�T�>�U:��]x�@�@�����s��=���>�`:>%���)�d�G�m��>��Z?� �?2�?-�=����h���
�˃C�ɂK>��%>h��>(�&?b��>�;>��ؾ.!"�
c��J�G�>E�>�D�>��-�� 5�z� ���D�Q��h.�.�?Yd�=C��>GQ?"�>�`I?�"?W��>g�>N8���ʾ.&?m��?���=>Խf�T�G�8��F�ä�>��)?��B�j��>i�?!�?��&?L�Q?ѡ?��>Ƕ ��J@�$|�>�C�>��W�1P��G�_>��J?��>x6Y?"ǃ?��=>;�5��㢾�
�����=tE>��2?h0#?��?I��>b��>������=���>hc?�.�?R�o?�p�=6�?L42>,��>��=A��>���>�?VO?��s?��J?U��>m̍<�=��G���r��OO�Gi�;>�I<?�y=�M��	t��[�7�<Y��;F���������UD�-󐼸��;w��>_D�>LF��&�J>kO��Ľm�>$���.+�����΂��~�=횃>�B�>^�4>M ��;�I=���>���>o*���/?�a�>W~�>�P�iGR��g��?�{�?��\?�X�>I�N���������}:>�v}?F�?����>��b?��]?eg�i=���þ׷b����Z�O?�
?a�G���>��~?e�q?G��>��e�":n�0��!Db��j��϶=.r�>0X� �d��?�>K�7?�M�>��b>'�=�t۾q�w�vq��B?��?�?���?8+*>|�n�V4�|I��:���[^?���>~���ӷ"?����aϾ����������N����Ы�_Q��� ��XV$�~ۃ���ؽ��=>�?�Cs?V�p?X�_?/� ��4d�	S^�����vV�<d��-�q�E�N�D��C���n��y������)��]xJ=��m���B��i�?�3"?:�i=�O�>u
��Vٵ����G��>�84�0���oZy=�u��>�.�=�1l�Hx��j����P-?��>cĵ>�O?":d��S��NE��d�,'�-<��Q�>I[�=�$? ܵ�x����'��R����x���<��g>�m?� `?׸�?;�O�RNU��m������'׽���#W>�I>��>�,��'��d[4�{NI���r�K��������a���=�&<?w�I>*��>�)�?Y?��辻3�}L �����<}C?O�B?"�>���=�8]��<�`��>�n?5��>��>B���;�)��%z��4�����>��>�A�>yp>k��� a�l���S�����8�O,�=�<b?׃��&Z���>�uT?�aP�m�R<�/�>��Q��;��z������/>��?v��=l[0>��ľ^�A|��)���7)?�l?�쒾nX*�[v|>�"?�>J��>�D�?�>ڙ¾s���K�?(v^?�J?�8A?���>�5 =:.��"�ǽ
�&��%*=:��>m	[>�j=1&�=T��[[������C=p�=c�Ҽ�!���w<�7����e<�P�<��3>�(ۿ�yJ��{ܾ~e���	��'��!��a�̽R�нV� �4�y��^{;��p��p����&�+�H�IZ����f�	�?/��?��������ų��Tq�	��K>ˇ�Bœ�9�ɾ!���]����e^����+/���D�>a��˸]�8Z?���3�ƿWE��e%�[Z$?-�?��+?}α�J%C�7N�!j�>���<ާX��r�
�����ȿ|7��IKx?���>��׾��D���?0I�>��>��=@U�3�l��`{��t�>n�K?&�>�B��@����w���Z::��?�$@v3A?��*����ɸ=[��>R�?�[;>��-�ns�2��}y�>���?��?�h5=��V�����e?o��<�C�J�����=���=(�3=����{?>���>[����6�*2߽>�5>�e�>BO�J�E�e�5=��|>R�ڽ�)½Lц?��<��1����`�{T>
U.?)u�>�`>��>��O�ɿ������F?#	@zZ�?ĕS?EZȾ�>�6׾��J?�['?��>�7&��̙�Q��<�׼*��	��\����C^�>3`�=��������B�v�<k��>�F�� ƿ�#��[���=�c<}'��H]�g���jq�X����[�iI̽�T�<���=,Z>Q�s>*<>Y�L>#fQ?J2m?X��>���=�pl��G���پ��3��� ��r���:������ྒྷ�����w�����s���\D��e=wP�VЕ�N.6���Y�Z�B�G1?�?w>�ڿ���W�k��<�O��;뉾2y�Pb��D�Ǿ��;���g�:�?r�F?]�����n�}���<cug���.?�}޽3	����L�>�`��=��f>��J�\�����C��B�ѡ.?� ?��ҋ��0=>���9�k=w&?�F?�m9<D��>��#?��&�R� �eV>�E3>`��>���>��=+��E%�f�?:T?|��xܟ�ښ>t����a��ʒ=�>a�!�Ҽ�Z?M>��<Gov�x��<�j��H:g<��A?$D�=J�
���>�&�о�G�<ue>AU�?�H���&)?�ǖ?.�T>'�>���h�^P����=;k?��?��>�{���E ���0K?V#�?���>tо��۾��U�����]
1?��V?�:?J{7��R���&���2?�>]?'<��f��YC��#������>Y��>�_�>8���:�>p?]�b����:H��Ī7�*�?@��?�*ɽ�	}���c>-*�>5�
?\M���'�x�C�[ǀ���m�>U붾l���WD\��e��?N?��?��$?|������if�=���
�?{��?8�m��*������(J�v��&���s�=�4�v�<Xy���I$�!㶾s�������m݌>s�@�僾��>�dn�k{�ۣ̿Sq�fM��oq��q�>L��>2<H@���o�9o{���1�����mL�/��>�>�Õ�������{���:�A�����>0���"�>�vR�������V�<���>=�>E��>dӪ��M�����?���5�Ϳ����%	���X?��?f�?�t?#�V<�5w��)}�
P��F?4t?�HZ?��&�ɀ\�J$<�Yj?k���_`�5�p�D���f>�1?���>!�*�+�l=��>#z�>Cx>�.�dÿ��������?���?�����>Qz�?��+?��OS��CŤ���(�D$�;��>?�
3>����K�#���=���B�?O�6?�[	�%!�]�_?+�a�M�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?е�� #�f6%?�>d����8Ǿ��<���>�(�>*N>dH_���u>����:�i	>���?�~�?Qj?���������U>
�}?���>��?P\d>�@?�>9�������\q>���=�D3���?��P?���>rw�=��"���3���S�1\�:���2XB�� S>xoV?`"@?,R`>����8��̱ ��U��hGe�k������x�S�=��;>��[>IU�=���`��
?E� �g�ɿP_���#3���e?��l�9�`>�fJ�����5�S��`q?y�>Ҏ��0���!y��Mm�-�?���?{b?n�����>R��=�-�>�Ϫ>�t<,�<>؄ξ�f�>Q�N?� ��-:�h�:�ʸl>F�?��?���?��k�5	?��&����}����=�*�j�=�r6?˸�N�x>@��>#��=�lt�=����r�
�>�T�?��?���>1�j?�%l�
A�jI=��>��g?rV?�vx����7%B>�x?4��kY�� ��c)c?�@��@Cv\?W��??߿�J���߯���Ǿ�<=�!�=A6~>E2����s�ᐙ��׽�$<tr=$��>�w>�L	>��=��*>V^=%�����a���=F���)F�I��� �Ã���;��r���O$��$;��˾���7�n�{���y��M�S�߽b��=�3q?�1_?{a?}'?�2�4��<�=�w�>2��|�i����>�(?CY?Z�9?���=HG��&�g��Iw��M��u�����>��=<��>)��>�&�>���=\
>���=���=9��<����i�h���<�m>��>��?���>�A<>b�>-ϴ�!2���h��
w��̽� �?B���-�J��1��S9��~���8k�=�a.?#{>���?п7����2H?t���*���+���>��0?�cW?�>����T��9>��J�j� `>�- �W�l��)�$Q>�l?��f>�u>��3�je8�^�P��|��>j|>�36?`鶾D9���u���H��cݾHM>�ľ>�D��k�{�����Tvi�z�{=]x:?ք?�6���ⰾl�u�VC���PR>m:\>U=�i�=�XM>bc��ƽlH��g.=(��=̮^>/W�>H˓>17E<��>Vg辰%�#U�>���=Zp�>�D)?{�5?�#=X��R#��q��j�>��?	��>���<�F����<&�>>��>�z�<#����I<�(H�`g�>R�=�Ci�<�����K���4>�A�>���=!���[0��˖~?r~���㈿)�j]��)mD?n*?&�=�0F<ׅ"�����,E��)�?8�@8k�?σ	�G�V���?2A�?S��U��=~�><ի>Dξ��L���?�ƽ����^�	�� #��Q�?�
�?a�/��ȋ�}l��;>�]%?��Ӿ�D�>�J��?��������n�H:�=�Y�>\�!?�y��M%��4����?>�>����a����ȿ�Uw�;��>���?�/�?��b�QZ����3�,r?��?lM??��>��ؾTo��.�>��@?<�K?P��>wy�=��?��?[��?�]I>�P�?�؀?���>!M:=(fQ���E�q�v �G�_��DF><�=�y���^��d~�]���ϷZ�d��*�?>�{=��>*7�(i����=�"ҽ9(Z�������>��J>[�a>Q?���>�[�> ;�>�`��!"/�B����Y���K?���?3���1n��X�<h��=X�^�&?�I4?i[�P�Ͼ�֨>��\?Z?�[?�c�>��$>��	迿�}�����<��K>�2�>\H�>K"��JK>E�ԾI4D��o�>WΗ>Y���@ھv-��>��$C�>�e!?h��>ծ=8� ?)�#?�j>)*�>_E�2:����E����>d��>�G?��~?��?^ѹ��[3����v桿��[�M9N>9�x?>U?�ʕ>J������mxE��LI�@�R��?�tg?VR�.?�2�?�??��A?H(f>Ό��ؾ߭����>]"?�j��[A��&��'�k�?�G?�l�>T����ӽ��ǼC��������?��\?�&?�����`�uþ��<�-%�����;�M��a>U>f��5L�=�x>��=�o��q7�>
�<ʼ=�t�>@��=P�8�_'��Z+?S\�=T�F���>��r�̪N�(r>%->ߴ��uC?�RC�oц�l���X������}L�?g��?�8�?��a|m�Y�J?�W�?a�>?� �>�Y��9�s{�¯�f<:=M��؎�=D�?4>�=���z���ճ��'���(���K�x?�6�>��?�}?��=aP�>5)��*���4ȾO��ʯb��2�Pq6�T��G������|�X����J��w0�>�贽T�>M�?�� >O��>�	�>�-���b>��>I'p>=�>a�=.�=��>u�=�v���Q?�Ħ��}!� ÷������E?JtX?(��>f>罃��N��J�?�t�?=�?d�>�o�22�h�>7�?[懾�?�U�=��鼽J-��_����V=)�Rr>8�G>G��<��/�\49��ީ���?�?F�=ִ��B@E� G��_(�=Ҋ?�T1?C��`�Y�V�p��\?�G`�%�����\��=ɾW1��q��E��8�}��z�M6!�i�=�7$?��?1���澐����.q�jWB�N�P>L7�>��|>OՒ>s�x>����`<��X��01�is��M�>#s?o�>��I?E�;?=jP?�BL?e��>�r�>:����>�T�;���>��>�9?��-?00?po?k+?�c>��������xؾ@�?�?�??��?U�?����g�½}K��1~j�Xcy����.o�=���<�2ֽ��r���U=�T>�@??��Ӿ8?3�Y�w����>ڻS?(|�>�?>�6��ӽi>$�>̕?M\F?\(���c���*��?M�?��ϼ�\�<	�=��f>,`����=�zĽQM)�Cߓ=�n6��5����=�5컝3�=�U==�����1<�ؽrk6=le�>�?q�>pU�=����2�����Ҍ�>3l�=!��>�r�>N5�=3m�����b!a�g%�>�d�?�<�?0����C�<�5>n�-���پ����&}���O+>�Z'?	��>|@s?`Ԥ?�+�>��*?
[4>_RȾ�钿PM�������b�>w!,?	��>�����ʾ��ԉ3�۝?g[?�<a����;)�ސ¾��Խر>�[/�g/~����<D��셻���=��5��?쿝?_A�U�6��x�ۿ���[��z�C?"�>Y�>��>V�)�|�g�r%��1;>���>gR?�A�>b�s?�k~?�]?S��>~xK������L���/7>'T>}� ?=�?f�?�Ć?a��>�ƺ=�z�� ����"L7��d�cHq�p��32>R��>�?z��>�C�=��4�6���XN�Կz���m>��>���>���>��>��H=`�??���>�@����ྃWξOuh���=,JT?"Q�?I%?��=�� �>9���w�>��?=+�?7,?��x��A>o��������f&���>��>Iќ>:��<�h=-9g>���>��>�_����;~�+�>[d?n�:?��u=�sҿ�&���[���1�������[���M?�����(N'�~�=)Sƾ���쒾ShJ��ޣ���������硾	兾�?P����=��$>�{W= ������<��>��1=��>,\��VH=�@�=��6O%��;�=���<���<�A=�˾�}?ypI?ƪ+?�D?��w>ż>�)1�+o�>Ē��,?�GU>�V�����?:�[]���B��x9پv�׾��d�����Qt	>�zI��>�"4>FK�=p%�<�!�=lt=͝�=-ߺ�4=��=��=0ʪ=;��=�>c!>@w?\6C�n y��W�2�?�ZhA?���>��}���X?���>��W���ſWr$�U0�?"@���?c+?���N]�>�4��ɽ�=����bP�=ۉ}>ɴ�Z]=�]@>dq�=4����i����پD��?jM
@�Z?�nq�um��i�=��7>,,
>�P�$�1�&�c��m��D[���'?_:�<������>3 �=�ܾ�˾#y�<K13>���=�l�Z���=����	N<=t�6=�E�>{�H>-#�=9?���}�=o=�i�=��>>ۗ�;��ռs�I��=�{�=�\>��">ƕ�>��?�Q-?c?��>Xh�Z�þpj¾���>���=mA�>�P�=��@>Ŀ�>Wg5?��B?d�L?zn�>�!o=Ì�>�S�>d�,��th��߾�8����=3�?���?���>��U<S5��7��T>�0���?�K4?�?f�>f��I��|4�������4M=e�M>��	X��DZ=w��h����>�5�>^Z>�j>�Q6=?֙=)�==1�>���=XI2��m�W�=���= Y½6�*>������<��j=����U�qӽ]s)=�5�=Q�=��~=���=�D�=��?3�>Ek�>x�">q�澖��><|޾�S��5o>��}�=`�<]v��)|��`�x.�N	>n��<\�?�����X?i�>��=�'�?V�s?��=H�-�U)z�?	��7)�ʽ\X�<��>�[��lO�a���I������>���>�3�>31m>��+��5?�YYw=��ᾔS5���>���Y���3q�0���🿑i�/���D?�A����=�
~?�I?$؏?V|�>����ؾ��0>���N�=<���&q�	���N ?'?��>m!�$�D��G̾���ܷ>�BI���O������0�{���ɷ�$��>������оz#3�Eg�������B��Mr����>߶O?"�?i:b�JW���TO�����'��5q?�|g? �>�K?�@?�$��sx��r��Fy�=9�n?a��?�=�?V>Ͻ=�紽d�>b"	?鳖?ݵ�?�s?H�?����>�Ԋ;�� >܋���W�=ܚ>�f�=��=�s?�
?�
?�N����	����A��^�ai�<+�=�|�>t�>��r>���=*�g=�K�=i\>�>���>�$e>��>�7�>v�ȾER۾k	R?GN2>�?��
?���>B>~�����*>blA�Gc���b��h����<��g=�
�����E�q��>lۿY�?D�=m!Ӿ�c%?�o�_Y�;��#�;��>v��<c̚>�$�>�p\>[N�>��>��=�u.>*�n>�v >�)� �X��l��*��˾���üx ٽ�����)��q�X :���o�{_�f��L}���]��Ta=���?�劽c_��
�骰�c~%?�Z�>�W�>�C���Ӊ��V�=�B?I:C>���▿�o��B��DB�?Q@@c>�>�zX?�?��.��W6��~Z��et�H�A��d��`����e󀿈�
�����i_??x?N�@?ف�<�?z>}�??�&�ȋ��aP�>^�/�I_;�;�:=���>�|���c���Ѿ�W¾���}BD>��m?�Ӄ?�?�wT�G�l���.>%`;?�?1?��t?�l0?��9?N��
%?�0>�0?)5?�4?�s/?��?�-3>��=�m���=�ɒ������ͽ�̽�a��u9=
��=W& ;�	�;"=�X�<������r��9�s���^�<
�<=Y��=W��=w��>�n]?�t�>�~�>f�6?֪��8�!���)�.?QbK=.���R��}��q��� >�Zj?ݫ?xfZ?��b>X�@���C�t�>I�>50'>.�\>�G�>�j��IG�^؊=�2>X�>��=�4C��ծ	��0����<|�>���>0�>F�#���T>�4��j������>��t�"ȾV���A���;�
%���ǩ>�JR?��%?ʑ�=S�����e�m��3,?
I?�pN?�Y�?h�=ȃ��=B��O�9���:-�>�!�<����C��]ۢ��C����9�">T
���d��<>R>����+m���G�9޾ �=
���̨=�)
�ϨǾ< ���>
>���<D"�����Ʀ�1.J?���=�w��93m��g���Z�=u�>��>�$���h��?��h��U=I��>��C>1�λ��'�F�YY�}32>��A?�in??u�?{/���m���.��ྦ����0�}L�>��>u�?ܞ>u��<�#��,w�(�l�L�B���>�>�>�"��IQ�z�󾶻�T���>�\'?��>�](?TT?^�?��s?��!?��?ya�>-����%?��?�J�=�׽�����f8�9a+����>��0?��&�i�>�?�?�&?ٮR?��?� >j�7�>��Ę>�Ր>h�^��ƭ��r>8|G?�S�>�V?x݀?��->��*��C��Bƺ���=��(>�+0?)&?�'?�`�>���>�С����=7��>> c?�0�?5�o?���=��?�<2>%��>�Q�=�j�>�t�>*?�iO?c�s?\�J?�r�>-p�<�Ȭ�hI���s�T�R��5�;S�J<��y=@��V5t������<���;3ظ�|����p򼢿C�i��|�;K��>�>Fo��b=Dھ2;���Np>��*>�̘��O_��V�z\>-�^>�?��
>Z��N͂=���>���>�����(?���>���>�*�$tk�4���ҽVW�>��V?�j�=8�b�����2����]<t�w?�S`?H�O����>�b?��]?�g��=���þ��b�L��i�O?r�
?q�G���>��~?o�q?i��>S�e��9n����Cb���j��Ѷ=�r�>xX�C�d��?�>W�7?�N�>��b>�$�=du۾��w��q��2?T�?�?���?�+*>�n�4���x)��ϳ^?�>�%����!?
�ѻh�Ͼ�$�����<���?��O����������"&%��H���޽�=U�?�?s?&�q?�}]?y� � 5d�
�_�>~�e�T�_"��\�8(E�W�D��C���l�-=���}���dAQ=.΃��*=�.x�?��(?RJ.����>�_����V�Ѿ�1>U9����g��=�݈�l�:=��:=�n�Z�:�{嬾� ?�ظ>���>7?�[]��>�o@3���3�3��)>�/�>�ے>�@�>Ab��Ҡ'���ͽ�ž���|�D��9Ol>OLc?e$N?w�o? ���`z0�d^��F�!���L��פ�X�3>�>�g�>��`���d�&�گ>��r�(Q����_
����=�v2?�8�>�Q�>���?h�?G��E��[����J/���<@ƹ>��g?m��>��{>�ӽm�����>�xn?ï?i��>ᭃ�p�1����>D��]��>�J�>�Ͽ>�Q>x9@� :h�F���}߆�v_����=i�D?8¥�򂏾bx�>?e?T�<�
>y�>���T�K�}����+ܾR�Z>Ʉ$?�B�=S
 >������P��O��gs3��p&?i?�2���(�s�`>��?��>:&�>�S�?7đ>{G��H�==?'[?�E?�;?U/�>U��<����Ž|�'� �<�~>��k>��S=���=���Q��� ��!7=X�=�YZ�O;���<�+Ѽ��<=l�<Ƕ@>]T�e�A���������������^�9ҏ����Y���Ӥ��摾s3}��_˽<���Fw�j��~���D�F�?���?
���������re�MCپ�]�>���K�=�x��M;+���.����+X��P�����J]e���'?�����ǿ����8ܾ�# ?CE ?��y?I�Ŗ"�dz8�d� >���<#ț�k�����W�ο넚���^?���>	�^����>n��>U"Y>q>P1���ޞ��~�<��?�c-?���>�`r���ɿ����鸢<���?��@ɁA?�(�r�쾫�T=4��>�	?�@>�0������>�>�2�?|��?�O=|�W�'���0e?�<5sF���ݻ�8�=H˥=m�=����lJ>N�>q��3�A���ܽ��4>t.�>�f$����!]^����<	�]>v�ս^L��P�?�k���b�*���j�Ơr>�:@?{�Y>9h��y� ?l�9��Ϳ�vf�&A? ]�?���?9�-?X����d>�־F�U?"�!?��R>��(�=T��T>$�	��|;\�˾��:�2�	>1��>6u=����޳�����=��>�h�-ƿS$�����A�<q�a��nZ���GϬ���V��1����p��w�	g=7��=�rO>�
�>��V>l_[>��W?_>j?3ɺ>��>��n����̾�8ڻk�����#��3p����߆�K߾�|	���������Ⱦ�*K��B=�V�л���5"��q[�3:�$-???�=뤾P�E��\�<�e־�ŏ�:>o��⿽�(Ӿ��@�d�p��?��??����p_��d
�:��rzɽj�]?H*��S��Y���3>�x�����=q�>Z�=U�뾩�:� �X���?�^3?�º�'����N<�⿾G��=v$?�1?a5-<m��>�R^?~%���u����#>縠=71�>;<2>�u7>M~��y�N�%�?��4?��V���#DU>�w��xo���d->�ʙ=�.S�e?�fgP>�؁��LT�3�D���Ѳ��=�X?��R>J-������P�30=�&>�=\?ɺ�>j�>�9n?[�C?nL>s���G[��u�"PҼϺW?\{?��8>�&��J޾��3��03?���?8ϴ=D���ǾX"����\��>0�?��?��=´���f��+!ݾ�h^?ϗq?�͉�w������:_>���>��>�l?MT6�@0�>ݪG?�6���p��n��jy2��l�?0<@�#�?w8߽��ż)�\�ڢ�>�D�>�&�7��;$ún$����W��:?i���T]�R9���>��6Q?ښ~?�֬>6�Ǿ��H���=�ו��Z�?W�?ӄ���(g<��1l��o���I�<Cɫ=f��H"�	���7�o�ƾ~�
����ڿ����>�Y@?L�]'�>�F8��5�lTϿ����Yо�Tq��?��>m�Ƚ𜣾��j�&Nu���G��H�^���ʖ�>Af>Z�=��C��+��t�A����>��>���='ؑ>� G�"���Gɽ��=�$l>�8�>��=d���Ҿ�F�?�迾�T˿!����;C�?5?��?.�y?�Mh?��>��������<��G?3S�?�3d?Cڈ=e����Z�9vg?�(���VN��5��Q7��VV>��<?qa ?�5%��7+=�%>?�� >q6������ꬿ�^�?�W�?!#꾄�?��?5?�3�����R����򾗽ټ��Q?�OT>����s8�|1F�$���6^"?l�6?g����a0��Wd?�'W��:.��L۾��>p�$?�3�@b��d_>��N��I���������?m�@2_�?ַ��n�P�x/�>,��>\F
��ބ�����+B>J��>	�=��ڼ	$�>1�0��r��~�;�,�?9; @O
?�͘�����c��>�u�?X�c>!2y?��p>� ?o�����:R >��?>��H>&μ4�?��K?`�>0"K>_�q���o&��#@���fX�]�i>�	�?�h�?2J�=�Rl�º�%%"�#��]��gv���z�	�X>h���P�=W(>�Y<=��m���3"?YM�*�ؿ�6��;�$�Tj4?x!�>
�?����cu��ۡ���^?Oa�>�����7��������?��?�	?�fھ���ߵ>W�>�x�>]ѽB����l��b�5>��B?���!��D�o�:��>Z"�?��@���?i�i�؏?���`�� 6��<߾Qֽ��=�.>?�ݾ���>��>L|>p{a��:��g	��L�>'^�?�X�?X�>7e?)����=Y�'5�>K\?�;�?�
?�9��3�q�F�]��B?��=��K�gL��b?���??r�?/�K?�١�?g�����)ԾF��o}3>C$�=*�=>� ݽ��>�I=6��<\�<�=$�B>�*:>o8T>a�8>3=>!�>���h(�����2��818����9���?���پR/(�!�$b����w��� ���k���7�Hʽ�g����<��R?\;e??v�?t��>5��zp,>�M�����=<�C�:�>�ב>��7?�;E?�?��v=o��]	h��'�b���vw��q�>�z>!�>�/�>$�>�M۽��U>&!&>��>K��=���=��?���=�X>��>���>Ҡ�>�(<>��>�ô�t,���h��'w���ʽ���?�b����J��*�����B������=�b.?�z>���==пyﭿ�-H?Vܔ�n.���+�~>g�0?�UW?�>�����U��C>��Ҫj�r<>{ �dl��{)�RQ>�k?D�>��g>;[2�V�?��}N�H��Xro>�9?1�ƾ?5�Q�q���8�S��T�[>S	�>c�o�H�!�
���Y#y��+b��t�=��??���>�0���j���T��9Ul��c> B>���;�^>B�P>w�]���zU�)�<�2>A�o>$z?SQL>��Z=�s�>7R��S�x�mݥ>�>$�@>]�<?�%&?�g=�½�~��wT�ۈm>NA�>�a�>�v >"K�[+q=\W�>z�T>�(���z����5���?�,G_>LA�=�]���u�:v��:��8?�=�m�=⹤�^x/���9m�}?�ٗ��T������,>��V?|�?�g���"�=_?B��,������?�k@[��?�����g���?��c?{Ľ�K�=� �>Ʉ�=I>4���о�S.?_P�Q��H�9���ᾘ׷?Nƙ?c>�;��K=_��V>;?��8�.5�>˷�z���dv��=|[�5b�@�>�H?�%���<W���?t�>�ϾZb���h��b�b�
��>i!�?ZZ�?�w�ᤚ�'/���>�\�?�XT?��>��C{��r�>o�*?V�}?f��>���a���A�>�<�?�O�?Q�H>U��?��s?Jq�>�x��X/��1������<=�[;�T�>Oe>����fF�Փ�Jg��m�j�@���a>��$=��>L��4��:�=����<��cf����>�"q>��I>BW�>f� ?;h�>��>8�=�n���怾����J?�(�?����Hk���T�=/�F�?��7?�&���̾V�>�C]?R=?��Z?#��>ָ�|r���߽����k�=�?->Ɂ�>��>_t��r	;>��Ͼ�@G��M�>���>���@�۾>���� �X��>x�"?��>f��=9a ?�Y#?�	j>��>^�D��R��$BE�B�>��>��?�~~?0?�c����2�)������KA[�͚N>��x?��?>�|���j����N�S;�Y����~�?o�g?k��W�?�"�?@?]�A?��d>�����׾�Z���Ɂ>��4?[�۾��?��� �:�����?�\�>�آ=�\c�����(Ǽ�8�Q>#���>�0�?�\^?�~¾ `W�3���+�w<���=�3�<r� ���2�5�0>��>��l�rҿ=��<HӼ�����U�8�=���==G�>�!>>����>V"?�Ž�l����?�U���'W>�<d�n5ξޚB?��	�U�g����#�����p��a�?Rҷ?'�?�:��{�� r?ˤ|?R��>�I�>� 	��໾F����X������M�� �>���>�
B��b$�{Ь��%��]��R�=�ž3�?��?r@?�B?H�>�:�>�۾�M�Z��\�=�D�M���Ǿi�2�Z�����FR�-��I��L����!����>w������>��>tp�>�7�>�w>}-�<��>��X>C�U>���>��=�i=�B���$��LC(�g9S?g/����߾a�Ծ��<?���?j:�>?�A��Z��Z �Gk#?:��?�_�??'E>�Oc��v+��?��$?un����??�Hh>F�g���������Z���~�=z3�7j>�;�����j�]�[�����>g^?]�>�ɾ%f1�����-��=c�?��(?�Y'�8Q���k� �U�R�S��3���o����-�#�3�n��ʎ��X��F����`)��&&=**?v�?~���~��ݱ�ۀk��Z>�[`p>���>��>��>��J>*���k.��[���#��yy��G�>�y?���> �I?��;?�fP?QOL?���>An�>������>�;��>�!�>ƒ9?V�-?�(0?�l?�j+?c>�;�������xؾo�?s�?�L?6	?i�?䅾�oý\|���f��y��偽=$�=	9�<m�׽�u���T=i T>6T=?䉺���+�q���b��>^+{?C`)>����.��'�>�<?j+>�	e?�	?g�ƾH����J��K?���?�}	��M�<V��=Vu<JV
��ɽ�8�=�T�=J��=�fǽpp�d��=K���b�=[ǉ�Hl=R�!=7�=�$�=�b�>��+?�>�ry>k��b���"�K>+��>���=�>>�Tܾd͉�b���`]���n>	��?5�?%�x�m��=���=��0��w�Y 	�p�ӾY�ڮ�>&͹>J3c?��?p!<?Ѿ?So>]��~
��(���.���#?H!,?�>}��i�ʾ�񨿼�3�Н?([?[<a�x��c;)�r�¾��Խ�>�[/�H/~����D�+م�����~����?�?�A�6�6��x辥����[��c�C?�!�>�X�>��>�)�1�g�y%��0;>���>=R?u#�>��O?�;{?#�[?5gT>��8�B1��\ә��3���!>�@?�?��?�y?�t�>��>A�)����S�������Ⴞ	W=�	Z>Α�>�'�>��>���=��ǽ�[����>�c]�=t�b>���>R��>L�>L�w>�C�<Z�>?/�>�a��ٛ	�_W˾��m=��h?�˔?`?!�<H�
�u83���f��>Aۢ?��?�s?��~���=���<��־�yf��n�>�g�>Sd_>̹�=Km=�ݴ=��>��>?��0��!;������?�}M?ə>ſ�=L�Y1v��(��g��<H�̾L�:���\�ac��E�>~���$��;ܾ��F�pv���]��m���ĳѾqR�F�>��=U�>
	=vk��2�eD�<>�>}y|����={��s`>��P�<�=VP̽B_��s��w�=?N=����n?��m?�p�?`��>{�>5�>�/���ݕ><�ح?�fz>���=!C��Hu۽#錾��ƾ�����"�dL���W>υ���Mi>��@>�DJ=��5�7�=)�>�_>@^�<�f����=� >d��=��h<��{=g(�=�5z?9��������㾇��>
L?���>l�ƽI�ؾ��R?,;�>hE^�%h����$�/�f?�L�?Fȥ?�ҟ>k�����>:j{�֎>���>�3�<L�>�9=>4��֝>Y�����w����нٳ?/f @2s?�2����ѿI��'7>I�>:R�K�0��]��Ph�W�yc!?~[7��̾�^�>42�=�Q߾Hľ�*=ד4>�e=�9�n$Y���=ǆ���x<=e�c=���>�P?>+�=S_���C�=܂R=�K�=+*Q>DO���7���+�t-=E0�=`�_>�|%>ڇ�>�b?�b0?<[c?,��>e�q��Ծ]쾾G[�>��=�S�>�l=L�?>��>��8?�HE?�hM?D#�>�e}=�>�ȥ>z�-�t�m��O�Ŗ��r+�<��?~��?X�>��<L(?�p�t\=�)"Ž��?;P1?ny?��>�v�R���%��-.�޴��lpU��*=B$r��V�z� ������b�=��>pm�>�b�>�!y>��9>�LO>���>xX
>�9�<���=p��=��<�ᐼw�=�Ҡ��C�<p.̼�%t��>��^)����t�X;܆];RwO<h��;���<�-�>�L>>��>���=�A��3�=��¾��G��}=Epݾ4�3��V��Tx�R�(�(�"�p�
>��=5|V�tN��j�?s�q>[��>g��?��B?�)>[�ؽ3?�~j���/������_�=&��=P�[�S�H��Oo��M�h2��F��>$�>�8�>~�l>��+�r!?���v=.⾛^5�F�>�����G���Q<q�!9����i�!o�K�D?FD��CO�=8 ~??�I?�ڏ?���>�_��i�ؾ:�/>�A���D=���9�p�S����?��&?�'�>t 쾉�D��%پ-�۽��y>�Ǿ��9����.iH���:>]M�G�>�����U�MBT���q�{���v�C�́���>�Q?�?4���7̇��,;�U�
��B{=�?�B?�$�>C��>R?�xz�c�Ǿ-����;��_?0�?j��?X&>�Ľ=/���0�>)	?㽖?��?)s?.�?��p�>��;ڹ >ؘ��f�=H�>゜=7��=�j?S�
?�
?�a���	�d��
��^�'��<�͡=��>�i�>�r>��=�g=�r�=K)\>�ў>�>��d>E�>�S�>�����S��a+?�>>���>U�+?4�>�.=����H��ZN���x\�{r(������׽��������Y���>H.����?g�">U��j?�����툼��\>��9>M乽y��>s;->��p>JP�>v/�>��;>'-�>�5>>�x��=��쾨�V�$�*�u�� ��?]���=Y=�a�I�>�l��W_D������W�2�v�8�6����=;��?1�&�t�5�7.��QD���>���=�63?I1��\ؼ�ke>c8	?��->cؾ�`��=���.����?��?M�x=��?6�x?��	?Rc�F���f怿��:���'�Sꂿ �X�1ޕ�uF]�5�����=C�M?I�z?�$?�Z�N�>ݻ�?�*-�o\;���>�&�(z�Q� >��?�}W����)�׾�"������>�*�?��?��?��Ⱦ/��@�/>"�:?.3?��p?rW/?��9?�5�2v%?a�->�4?=D?&�4?��-?��	?�0>��=%�<�� '=Ue��S��>�ѽ�Mѽ�z��1�0=�+_=w���< a=��<�Wռ$#�W�;�R����<|0=��=V��=�G;>�?1<�>���Q8!?�U����s���
�;F�?f
ž�뭾�A�פ�2�,��5�>ԯ�?r�?<3?xa����˽F\��^�=��=��i=��=���>�̥=]�%�o"�=*��>�8x>҅��������
����+�]9�>1�
>R��>��>&4=��/>����g�e�>d������X��я`����^�C��?�>!�D?��?��<�ؾg�};;�u�$V?�'�>"�Z?��?��˼�%*�6�!���Q��z>���>N�͋B�����:�����:|�=`0>�H%�����%b>C��5�޾|�n�{J����=$O=����V=^���վ�W����=6�	>����� �����ɪ��(J?F�i=)l���[U��l��M�>-��>�ޮ>X9�,�v��t@����f�=���>�;>�����ﾡuG���6�\>#mO?g�e?��?�1R���s�R	R���	�2���L+4�6��>}q�>��?��>��3>R"r��q��/_�)#�>��>)�?	2�ΩH���`����*�-��%�>�!	?�d���?$/H?�?�]L?�@?��?�vz>�?G��摾��?���?�"�=lNR�W�H�:�<��l���>c?
U��j>
o�>��?+`?�@m?!-?ș�=���	���>-̒>�.^��6���ʑ>C?�!w>g�W?~?��>�!�R:q���[�?㨼�)>f�)?�?��>^&�>���>����a=!��>��c?��?xEp?��=�� ?߆.>��>���=a�>�h�>��?��M?s�t?� M?��>���<������í���,���n�;�2<e�y=����m����m�<x6�9&Ӽ�x���� <�[���:�`:�>J�>;XὡM�>��Ǿ���>��ɾE]M���վ�U���=�i�>4�?��>��P�Jl��V{�>cH�>o�I�* P?��>���>�(>�@M��nݾS&���x>�8c?8�>�덿�������ܨ	���X?�K?���){]�n?��U?�{���f�%�`�K���)�T�s?V~?���|��>eo�?Jh?x?�S�����ƌ��ѵY�M4��y7I>���=��<��Ie���+>��K?_)	?��j>f\�>�*��d��?"f���>Y͏?Ǔ�?p�?=�*>�
D�c��P��������^?��>V��J�"?����Ͼ�#�������/⾩A��:�����O����(%��ۃ�f6ֽƽ=�??�r?�lq?��_? � ���c��^����wV�6���;��{E���D��rC�+�n�Z�s��{a��~H=.򀾴%<�� �?Wl)?�,���>�Λ����(;)�B>�'��#����=n�=U[>=�e���+�E3���f?c"�><��>P�=?�kY���;��u0��7�B���}8>�g�>�s�>��>��];D@&���b�ξ����D�ý�t>Bc?4�K?�n?�>�1�0��[��q!�kg.�/I����B>��>q��>��W��'�K&�[J>�3�r�^�����	���=��2?7��>�ǜ>��?h�?�s	�Zӯ�bx��E1��܍<
��>1�h?;�>]�>Gӽ�� ��<�>��g?��&?�0�>P f���)���u���ս"ʛ>�L�>+��>�dw>�2G�ضp�<��[Z��q$����=�1?�����[w���>s6m?��˼	� =���>FZ���&� :����g��>�?ӢM=�,>����I�H6w�pP��L)?�D?������*��'~>"?Y�>2�>z+�?�>�^þ��B��?�^?AJ?�IA?o/�>z�=�9��hSȽ��&�۩,=o�>[�Z>C�l=�z�=گ�<\��8��XD=:O�=�Ѽ<���6
<D���6�M<U��<��3>�qۿ?K�%�پ�C'�@
�p舾�u��j��c���]�����[x�x{��/'�!"V�FBc�������l�/��?/7�?Cy���,��ҭ�����D������>��q�;^��������,������ì��a!���O��#i���e�O�'?�����ǿ񰡿�:ܾ4! ?�A ?7�y?��4�"���8�� >�C�<�,����뾬����ο@�����^?���>��/��p��>ߥ�>�X>�Hq>����螾�1�<��?7�-?��>��r�1�ɿc���O¤<���?0�@��??��H��W���=��>i,?��>��;�U��x���?`�?��d?]f�:|�G_;��?2��>�v��<�<��.=��۽�z>+�=�6�<�S�>'Xw��;ʾF?�� �2>v �>$[=J\;��v����  �=:T�<(ĳ;��s?��}��rt���1�%)a���=��B?���>�LN>Y�?�S�6�̿�a`��v?L��?ϭ�?�%?3�����>ML��e?�4?��.>�/��|y���>�c>zڧ�QD��G�E��>��X>ScC>�f��	r��Z��U�>9�X=��#�ƿc�$����� =�����[��5��ڪ���T�v%��N`o�����h=8��= �Q>}a�>�
W>�!Z>ycW?��k?>P�>
�> �����ξR��G��#���������=�dQ�g�߾��	���������ɾ�G=�:��=��Q��>�����N^b�[�E�f/?n�>UʾQM��_<�:ʾGϩ�V���J��-cʾk0��m�N�?�_A?�م��SW����H��#��6�W?�.���������/�=����E�=��>��=��3���R��",?)1?T������U!>B��<�K���,?�e?}��=��>
�(?L��dS����=�ό=�C�>�z�>�:Իe�����"�fh(?8Y?t)7��k����>����P����=��=�5���
���u>���׻m�u��;&�<�_�=��V?��>� *�S�Z����¼0nY=�'s?1h?/�>D9k?�B?�
�</���U�m#�6��=\dY?M�g?��>�Ŕ�Ӿuǡ�و6?�d?^�L>��p�"��D-1�OA ���?uDn?��?���g~��ۑ��\��}5?�;k?�,_�I���������^ �>��?uk�>o�E�k9�>*M?�� ���z�Z4���sM��r�?ZF�?��?�9�<���m�T>(��>���=����Q1��~ކ�
����>�Q?�Ӿ�Qe�}[A�ԥ,��!?��?���>y���!����=�֕��Z�?��?e���,g<���2l��o��3f�<ƫ=c��A"�����7���ƾ�
�ݪ��g̿�H��>�Y@Y��(�>&A8��5��SϿH���Zо�Xq�6�?_��>��Ƚ�����j��Mu�^�G��H�H�����>K�>2���R����[�&L$�Ꭻ=��?E�ڽ}�7>P^c���e�.n��ݕ<=�N>sQ�>��>h);c�Ҿ[`�?�g0������v����/��K?��?��5?ߜg?����-R������#�:?���?�0?�k���ؾ@�=�j?o���W`�.�4�6E��=U>�%3?�6�>8�-�T|=V>D��>on>�'/�6�Ŀ_ж����R��?c��?�m�o��>�{�?�W+?�p�13���k��o�*�����;A?��1>����!�a-=�5Ȓ���
?�u0?\��~5���Z?�����u�j��F��=�'�>��`��y̾(��=P8<�(*��t�����c�?��?oʟ?���@�1���?ز�>���%���MJ>�-�>�X>�O�>e���\>�����_�fKս�+�?�s�?���>�r���&���6R>Xc�?B��>���?�O�>�p?�Q �vHT��R��ڼ�>��>����Hd4?�fJ?�ͯ>��>οv���/��C�K�A�f�%���G��(>īx?��z?1�%=�W\=fS?=�W����f¾��P��/����>g���R>�>#������,��G�?�p�ǖؿ�h��=f'��54?��>��?�����t��G�<_?�{�>>7��+��(%���8�嚫?�F�?/�?3�׾J?̼�>M�>BJ�>�ս���������7>T�B?W�eD����o���>Y��?R�@oԮ?gi�.�>���	⎿����%&�
ʋ��+�=�`3?o��F�>��>��="5��@���*g��p�> �?6 �?�x�>�v�?�`��m�W�����*�>y�?��?���C>�����=�g&?Nm4�59s��	�H�z?�#@:@�<?�J���忁d��J�ȾtU��.0�����=FU>����A����°<��B=AXu:��\=)�>D?>�u>9��=~D�=OT=��|�����٧��0��{$f� 3�d/�>�v���� A��g�N��Na���]��m,�I�ƽ��n�P
u���V]�=ՔW?��Y?J�w?mX�>V���>cf ��Oy=] <��@�=Ĕ>��2?�J?�%?U+I=|���r�h��끿��������^��>/nE>��>�b�>3�>F�{5H>*b:>|>:�>�J=���s�=YF>�{�>!��>�5�>�F<>5�>iδ�Q1���h�w��̽] �?p~����J�1���:�������n�=	b.?��>���W=пA����3H?���j)�̶+���>��0?�`W?��>���ضT��;> ���j�Sc>� �k~l�d�)�VQ>�l?WXN>uD>�.�=|;��?�@�ھc��>;tA?�}ӾI�нW$��җI��r���ɂ>I��>�I�=G���㎿��o���a��ڼ=~�5?��>P��v����h�㉄���>>�>�>�3=���=��->1d��+н���lf=�/>�\8>ۼ?0->�_�=��>���
^R��5�>�E>��)>�??�$?�&�D���D��WE0�Vtv><��>���>��>��K��ϰ=D@�>O=d>�/�Ա����xD=��U>�.}���^���p��m=$���}D�=��=� ���;�I�"=�2�?�ٓ���&� ��b�>��=?�LE??��=�P>2�־ث��1���?�J@X܆?��=����	?�!�?���J�>���>`��>b ��1{��q?V�ƽ�I���9�H�U���?��?5`�<�怿˸i��O�=z?�4K�Rh�>tx��Z�������u�c�#=S��>�8H?�V����O�T>��v
?�?�^�ߩ����ȿ4|v����>V�?���?g�m��A���@����>:��?�gY?zoi>�g۾J`Z����>ѻ@?�R?�>�9�}�'���?�޶?ӯ�?�$�=_g�?*�?3?�V�u�.�]2��f���*=�=39>~!f>ַ��
Z�e݋�=����p�����%>�C�<���>���:ī���<kZ���P�x��N�>b�w>�l>~�>��?��>f͆>�{r��m�[����ꂾ�bU?2�?!���Hj�Ct��2��=HK�j�%?�~[?��&�����>v�K?Xa?�>?���=����1瑿lJĿ�Ǿ^o>���=�m�>Ez+?$�"�n @��NǾlp��Fի>$��>�V���g��x)��n���:;�>�A,?�7�>�S>g�?��(?��>c�>��V�]����#�R�>��>��.?��?=$?�Fw��-,�f������=ge�s��=_?6�G?75�>����r�����pҼy�=\h�?ˌW?�8)��E?{Jk?oS?(�x?��x>�<�����ҽ�kU>��?;���B��'���۽o��>� ?���>��ƽL������B]"�����?{a?�{/?҄��w^��Z�����<cj����/;�h*;]D�Mm�=I�7>��!��=�=�1 >
�=�0\��"=�O�<	��=b�>���=:�!�Ȁ��'�!?@�?$��Fڇ;�[���?�J�W> I> �ʾ�Z?��!��{`�檤�儙��/����?���?>�?����m���L?��?tv?�v�>׾�
��A��o���i;��"�Rl6>��>���=��Ӿ}���a����~�ϕ��\���A?ш?b0?���>���=|�>2��rC���ξOi��#T���龦L-��'����:ľ�L�Q(>Mf��������>�xw��\�>t��>w�;76>'�>!2ݼ�1>�?>.e#>��h>�KK>ޒ�>��!>>�����7�"�_?�ꗾJ�������@�W4?��v?�h�>�k>����N��F?J�?���?�0>^{m�7A=�`��>�;�>�����+?�S�;&5ƼuIe=�ۡ��S���)��� �<[8>�Fa�X��[�X�^��l&�>��0?�I�=ᜲ��e�׫�����=��?�??+�%��SN�J�^�ʣZ��
@�0Lm=`���v?��"�4^|���U��UG���#�43�; i0?�Wy?������FϾ�[����� �>��>f�>*?�=0>)(̾��@<X�ұ ��>|�¼>�r?:r�>��I?"�;?�nP?�PL?���>�H�>����r�>:��;�>���>H�9?7�-?!0?�Y?`+?-c>�d��3��fؾ�?\�?1-?�?�?4����wý:	��(�f���y��܁�M��=r��<��׽��u��T=VT>��%?񉣾0Y��&���)�>4K.?K�?ڂ�>q���ț�i�i>l?��?2:�=�0�VMZ�&�&���E?��?�Ǩ��1�=��&>Z�=��ǻ��^=�BM=ԟ�=��>߹����.=��Ӽ:B�=�*�=�+=u�c=�ZH<�?s9k�<\�>" ?ŀ�> @�>6s��=^�-��e^�=�A\>U�L>�r>_nپ5�����>g�~�r>�?|�?��=���=7�=�����Z	����0�=)�>�$?G�V?6�?�@?�!?��>�������߾��&��7S?!!,?C��>���ϲʾ���3�m�?Q[?]<a�*���;)���¾�Խ�>�[/�+/~�z���D�5�����6���7��?��?A��6��x�ѿ��j\����C?� �>�Y�>r�>'�)�:�g��%�[.;>��>pR?�}�>ytP?֔z?�A[?UjW>ں8�ay���d���<�W
>�I??4�?S��?��w?ț�>.�>I�)�d�������]�����6���qD=��[>3�>�}�>z��>���=��Ƚ[+���=��q�= �^>��>1��>6��>�u>�A�<~�*?��H>����ߠ��ھ׷L��Z>8>c?u�q?	�b?��㽒��(�H�͖��@ٓ>�;�?]�?Y'?��.�y>yW��A�Q�xMu>n�3?�o�>-��!�=�$�=��?i$�>��I>�)^���g��M[�g�9?�`?���=Ha���N�2x���u��yL��3۾.p���(>�|��{D�=�׏��0���0��S��������|������߾r��t��>�=�B>v�>��Q>]�(�tL	��>x`���V�=�|����=X<��Um��20�jv��Y��O��<�Fp>&��ۊ~?~�`?t\?�0 ?<�\>I �=�(P��>�H�L*?�.>rG�=���^�)оĒ��ȷӾ0����}�=vV�(�P>^���.>�R>�j��qĽ/�<�S=��!=<r=1�,<%ү;�=��l=��x=:	�=Jʺ<�d=?����ߗ��$�Z��=���?R��<%J�֞g�"�/?? D��S��z���v�?�3�?��?�z>���Ɂ�>TLǾB&z=tA�>�[>e�>� �J�e�2=n>��>`���A���0=��?Ȇ�?�?�茿$�׿���=c��=8�=��A��g$�^D��5K���'�B�0?��]���>K�=���E���n<]ӌ>ws>O�^��=���-��<W�=��2>��T>�>r�ż81">�(�<$>�=1�1>7��(ٟ��v%��̏=e�=��B>c/>���>��?�0-?^�`?�	�>Q���ȣ�;��Da>_,�<R.�>|Qs=%�@>�
�>��<?�tH?��E?�>gѶ=���>MG�>ě0��o���վ�xb�;�Ç?�3�?�˨>��D<j�2�7����=�����H�?<,?3��>�g�>�W����[&�;�.����F����*=BAr�(�U�@���th���
��=�t�>���>�ן>~2y>��9>��N>3�>�>��<�p�=�����^�<� ��s,�=����ym�<�!Ƽj�����*���+�uS�����;r�;lM\<M�;s�=>��>4�=L-�>
� >��;��>�e[��_��!>��������S��|l��A;�����#��>��>�[�F˒���?Ǝ>8�>=[�?o�X?��'>	SV��*�+u����z��l��=�>��>>�5���(���S��"@�K�����>���>�>�	m>,��?��Jx=�3�R5����>����������G%q�{5���5i�)>ƺ�D?@D��Z��=�~?��I?bڏ?�w�>g��HmؾZ0>��^�=��7yq������?�'?��>G��D����g���5��>:E���Y:�G�sF=����=0������>��ľ|����E�o�p�����W>����ަ�> �h?ָ?W��{���C�9�I���&^�n�?nK?۬�>��	?��>$�׽EN�f����=\
�?���?FV�?*D�=,$�=^/����>�,	?�?'��?��r?�;��x�>]`;��>���9#�=�i
>-�=@+�=F�?��?M 
?K���c������rc��U=餦=Fx�>�N�>/�n>�`�=�R=؈�=�oY>�̟>ל�>Ra>^}�>Ã�>k��2���$?7��=7W�>j 0?���>`�M=�ѭ�0»<�1Y�/�A��C+��?����۽k}�<+�廔wO=Zxϼ �>��ǿ�_�?�aR>r��t�?D����a���U>ҭT>C޽E�>�,F>�b�>S��>�$�>��>�5�>��*>��U�=u	� 0�o�8�E[�����>����l�����7�}�͝��F���f�܃��S?�P�=��?����Y����s�����>�d�>U%?��`�7�5���=TS�>[vH>Kv�G��?��Rxƾ}�?��?��>�(�>םl?zR&?|��j�N:a�jj���)M�y�e��X��~���n]�� �6���tV?QS[?n�#?I��=x�>ݥ�?�X-��M���O�>L+0���Q��=�'�>d��ܽ�Ӷ�x��UA�����>�u�?�z?�G�>̇+���x��*>�m:?� 2?�?s?��0?E;?���$?��2>�8?�	?��4?g�-?��	?�->�/�=��0	H=����A�ν+�ʽ�(��%Z0=+�o=��;�<I�"=ܦ<���һ��8�ۺ>t��{��<��6=���=���=��J>�1�?	��>|
�=�bm?���룇��GI��6?����D��P��"z���Q<�S�>�n^?�Ԟ?���>@s�=J��s£�^E�>�5p>���Ѯ�=�9�>Dc����J�>w��=�`=4���z(�h|��1��������>�+U���>n=!>��ٰ�=�⩾��#�>��当���5n��iT�V�:�ۉ����>]�L?�(?�9�=l��k�;�f���<?Y�=?�4?-��?��d�:־(���i���q�i�l>���=j��������,
�rV=3�>�������%b>C��5�޾|�n�{J����=$O=����V=^���վ�W����=6�	>����� �����ɪ��(J?F�i=)l���[U��l��M�>-��>�ޮ>X9�,�v��t@����f�=���>�;>�����ﾡuG���6�\>#mO?g�e?��?�1R���s�R	R���	�2���L+4�6��>}q�>��?��>��3>R"r��q��/_�)#�>��>)�?	2�ΩH���`����*�-��%�>�!	?�d���?$/H?�?�]L?�@?��?�vz>�?G��摾��?���?�"�=lNR�W�H�:�<��l���>c?
U��j>
o�>��?+`?�@m?!-?ș�=���	���>-̒>�.^��6���ʑ>C?�!w>g�W?~?��>�!�R:q���[�?㨼�)>f�)?�?��>^&�>���>����a=!��>��c?��?xEp?��=�� ?߆.>��>���=a�>�h�>��?��M?s�t?� M?��>���<������í���,���n�;�2<e�y=����m����m�<x6�9&Ӽ�x���� <�[���:�`:�>J�>;XὡM�>��Ǿ���>��ɾE]M���վ�U���=�i�>4�?��>��P�Jl��V{�>cH�>o�I�* P?��>���>�(>�@M��nݾS&���x>�8c?8�>�덿�������ܨ	���X?�K?���){]�n?��U?�{���f�%�`�K���)�T�s?V~?���|��>eo�?Jh?x?�S�����ƌ��ѵY�M4��y7I>���=��<��Ie���+>��K?_)	?��j>f\�>�*��d��?"f���>Y͏?Ǔ�?p�?=�*>�
D�c��P��������^?��>V��J�"?����Ͼ�#�������/⾩A��:�����O����(%��ۃ�f6ֽƽ=�??�r?�lq?��_? � ���c��^����wV�6���;��{E���D��rC�+�n�Z�s��{a��~H=.򀾴%<�� �?Wl)?�,���>�Λ����(;)�B>�'��#����=n�=U[>=�e���+�E3���f?c"�><��>P�=?�kY���;��u0��7�B���}8>�g�>�s�>��>��];D@&���b�ξ����D�ý�t>Bc?4�K?�n?�>�1�0��[��q!�kg.�/I����B>��>q��>��W��'�K&�[J>�3�r�^�����	���=��2?7��>�ǜ>��?h�?�s	�Zӯ�bx��E1��܍<
��>1�h?;�>]�>Gӽ�� ��<�>��g?��&?�0�>P f���)���u���ս"ʛ>�L�>+��>�dw>�2G�ضp�<��[Z��q$����=�1?�����[w���>s6m?��˼	� =���>FZ���&� :����g��>�?ӢM=�,>����I�H6w�pP��L)?�D?������*��'~>"?Y�>2�>z+�?�>�^þ��B��?�^?AJ?�IA?o/�>z�=�9��hSȽ��&�۩,=o�>[�Z>C�l=�z�=گ�<\��8��XD=:O�=�Ѽ<���6
<D���6�M<U��<��3>�qۿ?K�%�پ�C'�@
�p舾�u��j��c���]�����[x�x{��/'�!"V�FBc�������l�/��?/7�?Cy���,��ҭ�����D������>��q�;^��������,������ì��a!���O��#i���e�O�'?�����ǿ񰡿�:ܾ4! ?�A ?7�y?��4�"���8�� >�C�<�,����뾬����ο@�����^?���>��/��p��>ߥ�>�X>�Hq>����螾�1�<��?7�-?��>��r�1�ɿc���O¤<���?0�@��??��H��W���=��>i,?��>��;�U��x���?`�?��d?]f�:|�G_;��?2��>�v��<�<��.=��۽�z>+�=�6�<�S�>'Xw��;ʾF?�� �2>v �>$[=J\;��v����  �=:T�<(ĳ;��s?��}��rt���1�%)a���=��B?���>�LN>Y�?�S�6�̿�a`��v?L��?ϭ�?�%?3�����>ML��e?�4?��.>�/��|y���>�c>zڧ�QD��G�E��>��X>ScC>�f��	r��Z��U�>9�X=��#�ƿc�$����� =�����[��5��ڪ���T�v%��N`o�����h=8��= �Q>}a�>�
W>�!Z>ycW?��k?>P�>
�> �����ξR��G��#���������=�dQ�g�߾��	���������ɾ�G=�:��=��Q��>�����N^b�[�E�f/?n�>UʾQM��_<�:ʾGϩ�V���J��-cʾk0��m�N�?�_A?�م��SW����H��#��6�W?�.���������/�=����E�=��>��=��3���R��",?)1?T������U!>B��<�K���,?�e?}��=��>
�(?L��dS����=�ό=�C�>�z�>�:Իe�����"�fh(?8Y?t)7��k����>����P����=��=�5���
���u>���׻m�u��;&�<�_�=��V?��>� *�S�Z����¼0nY=�'s?1h?/�>D9k?�B?�
�</���U�m#�6��=\dY?M�g?��>�Ŕ�Ӿuǡ�و6?�d?^�L>��p�"��D-1�OA ���?uDn?��?���g~��ۑ��\��}5?�;k?�,_�I���������^ �>��?uk�>o�E�k9�>*M?�� ���z�Z4���sM��r�?ZF�?��?�9�<���m�T>(��>���=����Q1��~ކ�
����>�Q?�Ӿ�Qe�}[A�ԥ,��!?��?���>y���!����=�֕��Z�?��?e���,g<���2l��o��3f�<ƫ=c��A"�����7���ƾ�
�ݪ��g̿�H��>�Y@Y��(�>&A8��5��SϿH���Zо�Xq�6�?_��>��Ƚ�����j��Mu�^�G��H�H�����>K�>2���R����[�&L$�Ꭻ=��?E�ڽ}�7>P^c���e�.n��ݕ<=�N>sQ�>��>h);c�Ҿ[`�?�g0������v����/��K?��?��5?ߜg?����-R������#�:?���?�0?�k���ؾ@�=�j?o���W`�.�4�6E��=U>�%3?�6�>8�-�T|=V>D��>on>�'/�6�Ŀ_ж����R��?c��?�m�o��>�{�?�W+?�p�13���k��o�*�����;A?��1>����!�a-=�5Ȓ���
?�u0?\��~5���Z?�����u�j��F��=�'�>��`��y̾(��=P8<�(*��t�����c�?��?oʟ?���@�1���?ز�>���%���MJ>�-�>�X>�O�>e���\>�����_�fKս�+�?�s�?���>�r���&���6R>Xc�?B��>���?�O�>�p?�Q �vHT��R��ڼ�>��>����Hd4?�fJ?�ͯ>��>οv���/��C�K�A�f�%���G��(>īx?��z?1�%=�W\=fS?=�W����f¾��P��/����>g���R>�>#������,��G�?�p�ǖؿ�h��=f'��54?��>��?�����t��G�<_?�{�>>7��+��(%���8�嚫?�F�?/�?3�׾J?̼�>M�>BJ�>�ս���������7>T�B?W�eD����o���>Y��?R�@oԮ?gi�.�>���	⎿����%&�
ʋ��+�=�`3?o��F�>��>��="5��@���*g��p�> �?6 �?�x�>�v�?�`��m�W�����*�>y�?��?���C>�����=�g&?Nm4�59s��	�H�z?�#@:@�<?�J���忁d��J�ȾtU��.0�����=FU>����A����°<��B=AXu:��\=)�>D?>�u>9��=~D�=OT=��|�����٧��0��{$f� 3�d/�>�v���� A��g�N��Na���]��m,�I�ƽ��n�P
u���V]�=ՔW?��Y?J�w?mX�>V���>cf ��Oy=] <��@�=Ĕ>��2?�J?�%?U+I=|���r�h��끿��������^��>/nE>��>�b�>3�>F�{5H>*b:>|>:�>�J=���s�=YF>�{�>!��>�5�>�F<>5�>iδ�Q1���h�w��̽] �?p~����J�1���:�������n�=	b.?��>���W=пA����3H?���j)�̶+���>��0?�`W?��>���ضT��;> ���j�Sc>� �k~l�d�)�VQ>�l?WXN>uD>�.�=|;��?�@�ھc��>;tA?�}ӾI�нW$��җI��r���ɂ>I��>�I�=G���㎿��o���a��ڼ=~�5?��>P��v����h�㉄���>>�>�>�3=���=��->1d��+н���lf=�/>�\8>ۼ?0->�_�=��>���
^R��5�>�E>��)>�??�$?�&�D���D��WE0�Vtv><��>���>��>��K��ϰ=D@�>O=d>�/�Ա����xD=��U>�.}���^���p��m=$���}D�=��=� ���;�I�"=�2�?�ٓ���&� ��b�>��=?�LE??��=�P>2�־ث��1���?�J@X܆?��=����	?�!�?���J�>���>`��>b ��1{��q?V�ƽ�I���9�H�U���?��?5`�<�怿˸i��O�=z?�4K�Rh�>tx��Z�������u�c�#=S��>�8H?�V����O�T>��v
?�?�^�ߩ����ȿ4|v����>V�?���?g�m��A���@����>:��?�gY?zoi>�g۾J`Z����>ѻ@?�R?�>�9�}�'���?�޶?ӯ�?�$�=_g�?*�?3?�V�u�.�]2��f���*=�=39>~!f>ַ��
Z�e݋�=����p�����%>�C�<���>���:ī���<kZ���P�x��N�>b�w>�l>~�>��?��>f͆>�{r��m�[����ꂾ�bU?2�?!���Hj�Ct��2��=HK�j�%?�~[?��&�����>v�K?Xa?�>?���=����1瑿lJĿ�Ǿ^o>���=�m�>Ez+?$�"�n @��NǾlp��Fի>$��>�V���g��x)��n���:;�>�A,?�7�>�S>g�?��(?��>c�>��V�]����#�R�>��>��.?��?=$?�Fw��-,�f������=ge�s��=_?6�G?75�>����r�����pҼy�=\h�?ˌW?�8)��E?{Jk?oS?(�x?��x>�<�����ҽ�kU>��?;���B��'���۽o��>� ?���>��ƽL������B]"�����?{a?�{/?҄��w^��Z�����<cj����/;�h*;]D�Mm�=I�7>��!��=�=�1 >
�=�0\��"=�O�<	��=b�>���=:�!�Ȁ��'�!?@�?$��Fڇ;�[���?�J�W> I> �ʾ�Z?��!��{`�檤�儙��/����?���?>�?����m���L?��?tv?�v�>׾�
��A��o���i;��"�Rl6>��>���=��Ӿ}���a����~�ϕ��\���A?ш?b0?���>���=|�>2��rC���ξOi��#T���龦L-��'����:ľ�L�Q(>Mf��������>�xw��\�>t��>w�;76>'�>!2ݼ�1>�?>.e#>��h>�KK>ޒ�>��!>>�����7�"�_?�ꗾJ�������@�W4?��v?�h�>�k>����N��F?J�?���?�0>^{m�7A=�`��>�;�>�����+?�S�;&5ƼuIe=�ۡ��S���)��� �<[8>�Fa�X��[�X�^��l&�>��0?�I�=ᜲ��e�׫�����=��?�??+�%��SN�J�^�ʣZ��
@�0Lm=`���v?��"�4^|���U��UG���#�43�; i0?�Wy?������FϾ�[����� �>��>f�>*?�=0>)(̾��@<X�ұ ��>|�¼>�r?:r�>��I?"�;?�nP?�PL?���>�H�>����r�>:��;�>���>H�9?7�-?!0?�Y?`+?-c>�d��3��fؾ�?\�?1-?�?�?4����wý:	��(�f���y��܁�M��=r��<��׽��u��T=VT>��%?񉣾0Y��&���)�>4K.?K�?ڂ�>q���ț�i�i>l?��?2:�=�0�VMZ�&�&���E?��?�Ǩ��1�=��&>Z�=��ǻ��^=�BM=ԟ�=��>߹����.=��Ӽ:B�=�*�=�+=u�c=�ZH<�?s9k�<\�>" ?ŀ�> @�>6s��=^�-��e^�=�A\>U�L>�r>_nپ5�����>g�~�r>�?|�?��=���=7�=�����Z	����0�=)�>�$?G�V?6�?�@?�!?��>�������߾��&��7S?!!,?C��>���ϲʾ���3�m�?Q[?]<a�*���;)���¾�Խ�>�[/�+/~�z���D�5�����6���7��?��?A��6��x�ѿ��j\����C?� �>�Y�>r�>'�)�:�g��%�[.;>��>pR?�}�>ytP?֔z?�A[?UjW>ں8�ay���d���<�W
>�I??4�?S��?��w?ț�>.�>I�)�d�������]�����6���qD=��[>3�>�}�>z��>���=��Ƚ[+���=��q�= �^>��>1��>6��>�u>�A�<~�*?��H>����ߠ��ھ׷L��Z>8>c?u�q?	�b?��㽒��(�H�͖��@ٓ>�;�?]�?Y'?��.�y>yW��A�Q�xMu>n�3?�o�>-��!�=�$�=��?i$�>��I>�)^���g��M[�g�9?�`?���=Ha���N�2x���u��yL��3۾.p���(>�|��{D�=�׏��0���0��S��������|������߾r��t��>�=�B>v�>��Q>]�(�tL	��>x`���V�=�|����=X<��Um��20�jv��Y��O��<�Fp>&��ۊ~?~�`?t\?�0 ?<�\>I �=�(P��>�H�L*?�.>rG�=���^�)оĒ��ȷӾ0����}�=vV�(�P>^���.>�R>�j��qĽ/�<�S=��!=<r=1�,<%ү;�=��l=��x=:	�=Jʺ<�d=?����ߗ��$�Z��=���?R��<%J�֞g�"�/?? D��S��z���v�?�3�?��?�z>���Ɂ�>TLǾB&z=tA�>�[>e�>� �J�e�2=n>��>`���A���0=��?Ȇ�?�?�茿$�׿���=c��=8�=��A��g$�^D��5K���'�B�0?��]���>K�=���E���n<]ӌ>ws>O�^��=���-��<W�=��2>��T>�>r�ż81">�(�<$>�=1�1>7��(ٟ��v%��̏=e�=��B>c/>���>��?�0-?^�`?�	�>Q���ȣ�;��Da>_,�<R.�>|Qs=%�@>�
�>��<?�tH?��E?�>gѶ=���>MG�>ě0��o���վ�xb�;�Ç?�3�?�˨>��D<j�2�7����=�����H�?<,?3��>�g�>�W����[&�;�.����F����*=BAr�(�U�@���th���
��=�t�>���>�ן>~2y>��9>��N>3�>�>��<�p�=�����^�<� ��s,�=����ym�<�!Ƽj�����*���+�uS�����;r�;lM\<M�;s�=>��>4�=L-�>
� >��;��>�e[��_��!>��������S��|l��A;�����#��>��>�[�F˒���?Ǝ>8�>=[�?o�X?��'>	SV��*�+u����z��l��=�>��>>�5���(���S��"@�K�����>���>�>�	m>,��?��Jx=�3�R5����>����������G%q�{5���5i�)>ƺ�D?@D��Z��=�~?��I?bڏ?�w�>g��HmؾZ0>��^�=��7yq������?�'?��>G��D����g���5��>:E���Y:�G�sF=����=0������>��ľ|����E�o�p�����W>����ަ�> �h?ָ?W��{���C�9�I���&^�n�?nK?۬�>��	?��>$�׽EN�f����=\
�?���?FV�?*D�=,$�=^/����>�,	?�?'��?��r?�;��x�>]`;��>���9#�=�i
>-�=@+�=F�?��?M 
?K���c������rc��U=餦=Fx�>�N�>/�n>�`�=�R=؈�=�oY>�̟>ל�>Ra>^}�>Ã�>k��2���$?7��=7W�>j 0?���>`�M=�ѭ�0»<�1Y�/�A��C+��?����۽k}�<+�廔wO=Zxϼ �>��ǿ�_�?�aR>r��t�?D����a���U>ҭT>C޽E�>�,F>�b�>S��>�$�>��>�5�>��*>��U�=u	� 0�o�8�E[�����>����l�����7�}�͝��F���f�܃��S?�P�=��?����Y����s�����>�d�>U%?��`�7�5���=TS�>[vH>Kv�G��?��Rxƾ}�?��?��>�(�>םl?zR&?|��j�N:a�jj���)M�y�e��X��~���n]�� �6���tV?QS[?n�#?I��=x�>ݥ�?�X-��M���O�>L+0���Q��=�'�>d��ܽ�Ӷ�x��UA�����>�u�?�z?�G�>̇+���x��*>�m:?� 2?�?s?��0?E;?���$?��2>�8?�	?��4?g�-?��	?�->�/�=��0	H=����A�ν+�ʽ�(��%Z0=+�o=��;�<I�"=ܦ<���һ��8�ۺ>t��{��<��6=���=���=��J>�1�?	��>|
�=�bm?���룇��GI��6?����D��P��"z���Q<�S�>�n^?�Ԟ?���>@s�=J��s£�^E�>�5p>���Ѯ�=�9�>Dc����J�>w��=�`=4���z(�h|��1��������>�+U���>n=!>��ٰ�=�⩾��#�>��当���5n��iT�V�:�ۉ����>]�L?�(?�9�=l��k�;�f���<?Y�=?�4?-��?��d�:־(���i���q�i�l>���=j��������,
�rV=3�>����ՠ��Cb>���N޾�zn���I�,��Y�M=�t��tW=u%�~�վn����=JS
>_c��� �S���Ȫ��)J?��i=}X���-U����l6>���> ��>�_9�~�w�ao@�ˬ�k��=���>'�;>�F���,ﾯ�G��	��&@>d�R?��f?A��?�����Z���]�d�2�M%��IU��!?��g>���>'/>���=���4����T�
,�]��>��?�V�6,S������,�q����>Un?趱�G�>�.7?Ѧ�>�*(?�+?z>4?�=�>&]�	���*�?q�?2	>߆��)iP�_a4��jY���>	2?����cV>7�?5)?�?�I?��#?��	>�t��}0��·>l�>B_K�o��2�u>y0>?�j�>�7[?)��?�Y>�-��錾� ���4=��>D?7?�?���>�W�>!t?wu�� �M=O��>��g?�ć?j?��=���>���=cg?�E->t�>i�>Uu�>نB?�9w?q,\?dٖ>P�<�ټQ�\����n�-�z���7���<s�<�����h����=�z����<�D�<�O�<j:�����%�,��>@$�>����O>D˾n���>kb�����0'ɾ��0���6>89r>J?�j>�#L�ժ5���>�&�>�7B�.�K?��?�[?���>'G�AQ*�k��w�t>��f?]?�=WOj��A��7tr�����$d?�nC?r�\��i�O�b?��]?@h��=��þz�b����g�O?=�
?4�G���>��~?f�q?U��>�e�+:n�*��Db���j�&Ѷ=\r�>LX�S�d��?�>o�7?�N�>/�b>(%�=iu۾�w��q��h?��?�?���?+*>��n�Z4�Q���������^?P��>�����;#?L	8��'Ӿ����E�����}���ܵ���씾�o��C)��>��Ǘ۽.�=��?Z�q?؁p?%�_?��?Hd���]��'���UU����a�/�D�`&D���C��`m��a��9�s���-<=p_��ˏ�����?�S?�}4��S�>Ϥ����%��q�J>�3��P���=�[･%��m�����zr`��*�����>A��>.��>�B?�T�BP9�� �pS�3�����>/��=^�>3y�>z�ѽҩ���ּ��¾�o��$��u>N�c?��K?�n?ܔ�*�0�v��ʝ!�m0���A	B>�>���>�
X�����*&�=>�u�r����������	��=f�2?��>Q��>6.�?��?�	��ᮾ��x�A@1��~�<ڹ>��h?���>�i�>�н�� �ͩ�>�}o?%?ɯ�>�ՠ�*~$��Qh��ԽG=�>�$�>f��>�-�>�t+�c�*?��U���p!%�/��=|�G?�S��	��a��>k�`?��,�)�_=Xu�>�4?�!`7������b����S>��>`��=̖>�4˾�0#�Y�v�O�X�C�(?Nz?f&��}s*���|>U�!?o��>��>DC�?���>_�þ
b˺x5?(c^?X.J?$�A?q�>�X=�б��ǽ��%�V�*=lΆ>r[>Dn=���==���Y�����F=���=�̼�)��� <���w�Z<���<ĸ3>�lۿ�BK��پ���?
��戾:���Jc����b��u���Yx�Ҍ�*�&��V� 7c�K����l�F��?�=�?%����0��8���f���i�����>�q�������N���)��Öྩ���0d!�F�O�&i�2�e�Q�'?�����ǿ񰡿�:ܾ5! ?�A ?5�y?��6�"���8�� >�C�<�,����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾?1�<��?6�-?��>��r�0�ɿc���N¤<���?/�@��E?����Nқ=�K ?)� ?{t�>_�.��_Ѿ�?��?Y�|?�T��n�c��A��hg?�+j>
R@��r��~�.>��}>}=�ӓ�۪K>�*f>� &������d����	>��>IM������a��=�i�>�퐽휚���x?+�[�OLX���%��"m��.:>�}L?�b�> =M>O�'?��9��^˿��[�E�^?��?�T�?�u?��ﾝ�>?����V?�&D?��O>z�C�O��,܋>顣=���<6O˾��V�|^O>fڅ>�>�ŉ�?j �\����=X[�==�H�ƿf�$��|��b=�:ݺ.�[�;}������T��"���go���轁�h={��=ŉQ>[l�>�$W>u2Z>�fW?k�k?|N�>V�>�5����ξm��G��K��X��������Q�O�߾R�	������U�ɾ"6=����=$P��G�����/d��TE���/?>P�ƾJiM�H�<�m̾�>��N����Ĝ�*%žŰ-�g�m�<��?�5A?�τ�v3U��U�e��[���W?������U�����=�ױ���9=���>�=�=��⾹�2��HQ�or.?�� ?ϸ��z���c+>g��er�< �.?�?��;��>�"?)M(��7��^�U>��/>�s�>X-�>���=_����Lｅ�?��V?�x�UP�����>����ׄ�>�=�>��1��k��V[>Ӧ<�O�����k��9��<��N?��%>Y�/���Һ��m;}݊>Ha?'	�>)z�>M�k?@�L?9��<15����e�\5�y�Q>�Ng?�V?UP>f������O�=DU?a	Z?@�>���Ia��LW��/�;��>y?U�/?�1���2��Ј�s��MJd? dS?��z�k���{�G�6���>���>��	?�6�qC�>CW?��@�C!������w*��?b� @��?�b���B;�ܕ��z�>�?�D��ң�M=��(�Z��$��?n����F{��0�$N?��|F?[2i?�Ƕ>܍Ⱦ�r�N0�=?���D�?�_�?�ȩ��ٍ<kz��_m�� ����<�n�=\9���%�����~7���Ǿ��� ��� ��}>�@!y�~��>�:�]\�(�ο������;�l�U�?��>iɽi�����i�L�r��oE�A�G����<�a>7�i>��u$��T�V��k;��wa=h$ ?/��<D�U>~+ǾJPz��qȾ�:�=&hy>�u?���>���F�ھX�?��#����~�t��6��1f?�%�?=y$?��G?:d��!!��9���=�d?7�?ܧ<?�޸�B��&P�=�j?�{��9b`��c4�X�D���U>�3?�:�>�b-�G�x=G�>�o�>#>Z%/��Ŀ�����?�����?#k�?q꾴��>���?�v+?�0�홿6���*��,���@?��1>�����!�g9=��r����
?�0?*��\��c?r?e�=��ED�Q�٠����>l?[�dO��}zF����E����������?I�?L��?ބ���QR��5?c.�>kd����D>���>]�>V�����#�<Q%�#d۾e����$�{��?�u�?�)-?��Ɲ����=��w?M'�>���?�g�=��>���=�e���C�ɡ >���=�.G�ը?�LM?ݎ�>�:�=d�8���/�~�F�x*R��h���C�/d�>_Ka?t>L?�B`>)��0Y4�Cg!�%"ν�0����Y�?��g*��]⽃m4>�O=>��>C�D���Ӿ�M?�%��~׿����ic��+4?��>�o?�� �S�|�JjS<�6]?�ċ>��" ��y���������?eC�?��?\�Ҿu��M> $�>��>~�ӽ�ޙ�ﾅ��0>@??AW�J>��[�o���>�?�@Ik�?>�n�Q#�>q�.֍��ٔ������T��g=��:?7������>]�	?��W>ץx�6읿��q���>�W�?01�?�7�>$��?5ї����-�m>�S�>�g�?��?�����:���5??i)3�Vy:�+<"��f`?&r�?Bl@u@K?�����ֿ����]��n�þ��=���<�`>L���QNS=�*�=-b����<���=	�>u�+>$ (>��>}�>�23>�����A�Pҧ�Ң��u�>��T(��]&�~��1��@H<�WZ�������׾��ؽ�@��v��s��� "��L!=�b�=�W?w9R?��m?�V�>�߁���>������3=�.�K�i=�Ʌ>�0?�fI?�*?W�=TǛ�q�e����~��������>�v<>k��>o��>)�>��!<TS><B>>��=��=m����=��O>�/�>��>�u�>�G<>�>:δ��0��V�h��w�̽���?�}��k�J��1��;;��U����q�= c.?ـ>����>п�����3H? ��|)���+���><�0?``W?Z�>�����T��A>��N�j��e>� ���l�ʏ)��Q>m?���=	�>L�E�/�ɐ������?�<A?�@��S�C�;x�i�O��?�!Ѓ>4��>xI9>sU���,��
\\�%?��s\@>{�(?��>iӒ���ž�=���c�O>A��>��p<�u�=
>��o��e �v�)�+\�=�W`>}:_>�?��><��=h@�>(ゾE����>��3>!F>��0?��/?�h�<5&��:c��ْP��Wz>X�>a$�>x�=��f�Q>�$�>��#>ī-�Co��j*�6�(��;G>�)��W�5��r�;c�K����=���=B�HA��w'=�݊?�(���SJ�gֽ�,�;^]:?�`�>(m�q�����6�� ����ľ4��?.�	@���?|�Y�����É�>���?��Y�o�=� >���>\y׾�'����!?�7��ks{���>��x����?m�?���=�I���/k�6��=�2)?����h�>�y�;Z��P��[�u�F�#=���>z8H?W��ܵO�>�hw
?"?]_�ܩ����ȿ�yv����>b�?c��?��m��A���@���>Ϣ�?sfY?fli>j۾gZ�R��>��@?B	R?Y�>�9��'�x�?P޶?��?�0B>>ё?�0t?�b�>��o�ej+�"�k���͈=�_r�b��>�<>�)��=tC��}��^����g��S���b>��=�)�>���ņ���G�=&冽~˥�e�>�9�>�g>�B>��>\�>�[�>���>��:=g�����ϛ��P�K?���?����2n��N�<i��=��^�h&?�I4?s~[���Ͼpը>��\?8?�[?�d�>��S>��迿~�����<+�K>g3�>�H�>7$���FK>�Ծ�3D��p�>�ϗ>�����?ھ--���V��3B�>�e!?R��>�Ү=ۙ ?��#?��j>�(�>CaE��9��V�E����>ע�>�H?�~?��?�Թ��Z3�����桿��[�w;N>��x?V?sʕ>b�������kE�8BI�>���]��?�tg?�S�0?<2�?�??_�A?y)f>ه�(ؾp�����>�x
?*��4xT�E��^,�<��	?9��>3FZ>�d��ii=�Y=["o�����?�o�?y??��������8
����=��{>��%>�U����^4>�I�=EK��X�>O <��~��Y���"��>�=S�2>>�y�q�.���E>��%?�|<N^f�v!`=�b�I�A�&Kt>"�N>⦾�DV?yp��b�ϱ���G����o�8U�?XE�?���?R��<n��&E?���?�q	?���>�L־{���?Ⱦ�2���?�]�"�\�>�0�>`�;(nܾ�&��e���� ��嗽0�h�=
?��?u=5?Xs
?���>�->��Ѿ&--���־|�پ��2� �ɔ �F��eP�Lپ(�N���o>iW��1DP�
��>�ǽ�?�>!;?
I>gđ>1"�>�.[<�ͪ>�s?>��>R:>��>����81p=ĳX�9��) _?\ڱ� �����W��T!?��q?�:p>=�L����d.$��j;?�`�?��?d��>Ds���eI�>��>s�?޹���~0?21O>>���ݽ�W�I��m��+�C�L,��a`>tQ9�0:�V�y�Tȋ����>��$?aLf<*{ǾjI̽�����r�=}�?�+?�(�ۜN��ho�+:Z��>S��1	��]g��P����#���n�m쎿`���̓�mc(��~-=f/)?ᮈ?�G�	f뾀O��T�l���>�(�a>�$�>V��>Ԯ�>($C>����1��0[��p"�S|�rV�>��w?�>%�I?�@<?u�P?�L? �>��>����5��>Mc�;;�>j6�>]"9?�c-?ӹ/?G? S+?)�b>����j����ؾ��?^?1�?�?��?�E����ƽ6/w���w�Yx�+����=D��<��ؽcCy���S=G�S>�#?�}���\�Q&վ���>>�?�?���>}V������a�>,�>e�?
>��:���r��ݦ��r?%2�?[����<h��=ki|=݋�<��c=�����:cz\>Y����<܃����=�l?���I�=qc-���D=�cƽ�e�>C�?�\�>;��>�4��Cq �b ��V�=h�Y>�8S>�!>�;ؾ�Y��X��3�g��gy>�{�?ce�?+|`=�(�=�1�=�I�����T���������<�8?5�"?CT?�S�?K�=?W#?T#>�(�A4��)��̪���?�,?8��>���'�ʾ��D�3�U�?�Y?,7a�����:)��¾��Խ��>�Z/�x,~����D��{��3������'��?]��?,@A�J�6�1s�k����e���C?d�>_�>�>I�)���g�4$��;>p��>�
R?�˵>X�W?��y?�iU?��F>�6���������=f�=��0?(�y?_g�?�j?I�>��M>̨ ��v�"a���(�����J���C�9��c>Ȥ�>�q�>��>y�>�pȽHۼ��^6���=��@>��>�ݯ>���>�6P>3G
=��?V!�>�a��'����&�X��3t�>q�x?$�?�\M?���w��zF�{K���>�Z�?G�?s.?��<���Z>h��mq�$	���?��>���=ģ��媽��=�� ?��?�q^=zd0��3u�	�M�[�?�T`?�-=��ſ[�p���n��n����}<������d�B'��Y]����=�.�����9���\�"���68������훾&&|�S��>��=���= G�=���<NoǼZ��<-�M=A}�<�=�Ww�G;f<�9������⇽(6���*U<��G=����־h�x?��b?^E??�2?���>C��=��1.'>�71���>�Uk>�}���5����F��@˾����|�������j�ܒ��Ë�=�p���2�=��>aF�=]�,F=�+2=��=��C<�t&=6�s=E��=���<�i=�4�=�:�=H�J?O|������$,�6>V�0?Q��>k�M>K�sZ?fe�>	���ߛ��3�{�o?� �?e�?Z��>��
�i��>�Ҍ��g�=�::>���=$�=)>ǾH֠>t�=4�ܓ���3���?�8@>S1?�,��I(ۿ��=�2�=uGA>��A��'3������OU���.?�E��b���NJ>�>q��!��]렼BzQ>v>�i��Z�L�8=8�	x_=�Ld=�l>�U>q>O�;�V��=8�;��3<&u#>�/��"=O�޻�=ƌ�=�A>�>���>C�?ʙ1?	A_?_@�>�p��޾X�Ⱦ8�>�Փ=[Y�>��z=��5>�)�>�W5?�\G?�H?M/�>���=�3�>\?�>�p*�۸n���ؾe����,�<���?�,�?�w�>�q<��9�}��}�=������?Fv0?4R?�u�>�U����9Y&���.�#����t4��+=�mr��QU�J���Hm�5�㽱�=�p�>���>��>8Ty>�9>��N>��>��>�6�<yp�=ጻ���<� �����=�����<�vżƗ���u&�6�+�2�����;f��;B�]<u��;��=M��>�2>J�>>&>�ݾ|�>hi�pH�q�>g�����'�INb�w�}1�N�&��|>>ф>�@ؽ�����?��Y>�`->D��?��T?B�>�:<�3���@���k����\��"�=��/>A�9�*�)��jM�hGA��ӿ���>���>&Ф>Ƀp>�B,�>��Nw=���,5���>�i��4��d ���o�����	����h����7D?�P���|�=��~?J?L�?p8�>�s��(�ؾ$O->��{�N�=m���<w�������?	�&?��>9쾜�B��59���[h�>���^$7�H��1�L���R>�������>Ndƾ�����?���t��U����A��㝾 >�>J�i?#v�?쵶�
���C9�������8<y?)�J?p�>� ?sj?:��H���=��,C�=�L�?=��?���?���<:K�=�G����>"�	?��?��?C�o?�D����>	
���0>h/�����=zc>W͉=?��=��
?��
?�1	?j���_g��쾡����\�#`�<�,�=&�>��>�p>*��=�&z=̯�=��[>xҝ>-��>P�_>��>h8�>��������,?�z>jY�>n!?�s|>��=�>H���<��+��%>���,�z���-���:Q�<��=��d=��u�\��>�~ſ�|�?yȎ>M\��?q߾� ｽ:>���>�.�O-�>�6>]q>��>3��>�v�=�Y�>�(!>s�=�i�>� ��G�!�7�=fj��,�����>Zo���cd������=��y��
��?��d�v�����I�6��>�[I?�Fa�,z��	X�g-����>���=N�D?Y�����=b=�J	?��
>� ������������#�?89�?�O>ܩ>)Z?~?�(6��R0��_�w�}�;:=�}n_�D.X�1,��#�}����}�P�W?[�o?��7?l�<T߃>G��?˧$��Z��_�~>.�5��l:�1��=�!�>�q���uo�%�Ͼ���q'��=W>�v?̈́?-j?�c^��p���'>V�:?��1?Tt?Kf2?V;?����Z$?Q22>E??�<?0�4?��.?�
?�E0>���=�ʽ��U0=����Xꊾ��ѽ�N˽����5=�qz=Kk$��<HO=���<%I�X�ؼ��:n�����<��8=�ˡ=?�=g�C>}	�?�	?��=�C+?D��y�Q�hq����?eN�EP�޻V�L�q�3��k��=>KR?�3�?���>o�<=���T�'�>��>�/�=F�R=b�>t_>q��M�0>�gr>A�j=F��=�ܽ� ��n���*��3-]>T������>��q>�k�`%>����Dys�wXm>��Q�	���o�P�'�F�1�����.��>%`J?B�?|=ז뾌����g��+?=�??��H?G�u?8@?=�kξ%0���I�����Q�>߉�<���&��y����`4��9�<ɔ~>�w���ՠ��Cb>���N޾�zn���I�,��Y�M=�t��tW=u%�~�վn����=JS
>_c��� �S���Ȫ��)J?��i=}X���-U����l6>���> ��>�_9�~�w�ao@�ˬ�k��=���>'�;>�F���,ﾯ�G��	��&@>d�R?��f?A��?�����Z���]�d�2�M%��IU��!?��g>���>'/>���=���4����T�
,�]��>��?�V�6,S������,�q����>Un?趱�G�>�.7?Ѧ�>�*(?�+?z>4?�=�>&]�	���*�?q�?2	>߆��)iP�_a4��jY���>	2?����cV>7�?5)?�?�I?��#?��	>�t��}0��·>l�>B_K�o��2�u>y0>?�j�>�7[?)��?�Y>�-��錾� ���4=��>D?7?�?���>�W�>!t?wu�� �M=O��>��g?�ć?j?��=���>���=cg?�E->t�>i�>Uu�>نB?�9w?q,\?dٖ>P�<�ټQ�\����n�-�z���7���<s�<�����h����=�z����<�D�<�O�<j:�����%�,��>@$�>����O>D˾n���>kb�����0'ɾ��0���6>89r>J?�j>�#L�ժ5���>�&�>�7B�.�K?��?�[?���>'G�AQ*�k��w�t>��f?]?�=WOj��A��7tr�����$d?�nC?r�\��i�O�b?��]?@h��=��þz�b����g�O?=�
?4�G���>��~?f�q?U��>�e�+:n�*��Db���j�&Ѷ=\r�>LX�S�d��?�>o�7?�N�>/�b>(%�=iu۾�w��q��h?��?�?���?+*>��n�Z4�Q���������^?P��>�����;#?L	8��'Ӿ����E�����}���ܵ���씾�o��C)��>��Ǘ۽.�=��?Z�q?؁p?%�_?��?Hd���]��'���UU����a�/�D�`&D���C��`m��a��9�s���-<=p_��ˏ�����?�S?�}4��S�>Ϥ����%��q�J>�3��P���=�[･%��m�����zr`��*�����>A��>.��>�B?�T�BP9�� �pS�3�����>/��=^�>3y�>z�ѽҩ���ּ��¾�o��$��u>N�c?��K?�n?ܔ�*�0�v��ʝ!�m0���A	B>�>���>�
X�����*&�=>�u�r����������	��=f�2?��>Q��>6.�?��?�	��ᮾ��x�A@1��~�<ڹ>��h?���>�i�>�н�� �ͩ�>�}o?%?ɯ�>�ՠ�*~$��Qh��ԽG=�>�$�>f��>�-�>�t+�c�*?��U���p!%�/��=|�G?�S��	��a��>k�`?��,�)�_=Xu�>�4?�!`7������b����S>��>`��=̖>�4˾�0#�Y�v�O�X�C�(?Nz?f&��}s*���|>U�!?o��>��>DC�?���>_�þ
b˺x5?(c^?X.J?$�A?q�>�X=�б��ǽ��%�V�*=lΆ>r[>Dn=���==���Y�����F=���=�̼�)��� <���w�Z<���<ĸ3>�lۿ�BK��پ���?
��戾:���Jc����b��u���Yx�Ҍ�*�&��V� 7c�K����l�F��?�=�?%����0��8���f���i�����>�q�������N���)��Öྩ���0d!�F�O�&i�2�e�Q�'?�����ǿ񰡿�:ܾ5! ?�A ?5�y?��6�"���8�� >�C�<�,����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾?1�<��?6�-?��>��r�0�ɿc���N¤<���?/�@��E?����Nқ=�K ?)� ?{t�>_�.��_Ѿ�?��?Y�|?�T��n�c��A��hg?�+j>
R@��r��~�.>��}>}=�ӓ�۪K>�*f>� &������d����	>��>IM������a��=�i�>�퐽휚���x?+�[�OLX���%��"m��.:>�}L?�b�> =M>O�'?��9��^˿��[�E�^?��?�T�?�u?��ﾝ�>?����V?�&D?��O>z�C�O��,܋>顣=���<6O˾��V�|^O>fڅ>�>�ŉ�?j �\����=X[�==�H�ƿf�$��|��b=�:ݺ.�[�;}������T��"���go���轁�h={��=ŉQ>[l�>�$W>u2Z>�fW?k�k?|N�>V�>�5����ξm��G��K��X��������Q�O�߾R�	������U�ɾ"6=����=$P��G�����/d��TE���/?>P�ƾJiM�H�<�m̾�>��N����Ĝ�*%žŰ-�g�m�<��?�5A?�τ�v3U��U�e��[���W?������U�����=�ױ���9=���>�=�=��⾹�2��HQ�or.?�� ?ϸ��z���c+>g��er�< �.?�?��;��>�"?)M(��7��^�U>��/>�s�>X-�>���=_����Lｅ�?��V?�x�UP�����>����ׄ�>�=�>��1��k��V[>Ӧ<�O�����k��9��<��N?��%>Y�/���Һ��m;}݊>Ha?'	�>)z�>M�k?@�L?9��<15����e�\5�y�Q>�Ng?�V?UP>f������O�=DU?a	Z?@�>���Ia��LW��/�;��>y?U�/?�1���2��Ј�s��MJd? dS?��z�k���{�G�6���>���>��	?�6�qC�>CW?��@�C!������w*��?b� @��?�b���B;�ܕ��z�>�?�D��ң�M=��(�Z��$��?n����F{��0�$N?��|F?[2i?�Ƕ>܍Ⱦ�r�N0�=?���D�?�_�?�ȩ��ٍ<kz��_m�� ����<�n�=\9���%�����~7���Ǿ��� ��� ��}>�@!y�~��>�:�]\�(�ο������;�l�U�?��>iɽi�����i�L�r��oE�A�G����<�a>7�i>��u$��T�V��k;��wa=h$ ?/��<D�U>~+ǾJPz��qȾ�:�=&hy>�u?���>���F�ھX�?��#����~�t��6��1f?�%�?=y$?��G?:d��!!��9���=�d?7�?ܧ<?�޸�B��&P�=�j?�{��9b`��c4�X�D���U>�3?�:�>�b-�G�x=G�>�o�>#>Z%/��Ŀ�����?�����?#k�?q꾴��>���?�v+?�0�홿6���*��,���@?��1>�����!�g9=��r����
?�0?*��\��c?r?e�=��ED�Q�٠����>l?[�dO��}zF����E����������?I�?L��?ބ���QR��5?c.�>kd����D>���>]�>V�����#�<Q%�#d۾e����$�{��?�u�?�)-?��Ɲ����=��w?M'�>���?�g�=��>���=�e���C�ɡ >���=�.G�ը?�LM?ݎ�>�:�=d�8���/�~�F�x*R��h���C�/d�>_Ka?t>L?�B`>)��0Y4�Cg!�%"ν�0����Y�?��g*��]⽃m4>�O=>��>C�D���Ӿ�M?�%��~׿����ic��+4?��>�o?�� �S�|�JjS<�6]?�ċ>��" ��y���������?eC�?��?\�Ҿu��M> $�>��>~�ӽ�ޙ�ﾅ��0>@??AW�J>��[�o���>�?�@Ik�?>�n�Q#�>q�.֍��ٔ������T��g=��:?7������>]�	?��W>ץx�6읿��q���>�W�?01�?�7�>$��?5ї����-�m>�S�>�g�?��?�����:���5??i)3�Vy:�+<"��f`?&r�?Bl@u@K?�����ֿ����]��n�þ��=���<�`>L���QNS=�*�=-b����<���=	�>u�+>$ (>��>}�>�23>�����A�Pҧ�Ң��u�>��T(��]&�~��1��@H<�WZ�������׾��ؽ�@��v��s��� "��L!=�b�=�W?w9R?��m?�V�>�߁���>������3=�.�K�i=�Ʌ>�0?�fI?�*?W�=TǛ�q�e����~��������>�v<>k��>o��>)�>��!<TS><B>>��=��=m����=��O>�/�>��>�u�>�G<>�>:δ��0��V�h��w�̽���?�}��k�J��1��;;��U����q�= c.?ـ>����>п�����3H? ��|)���+���><�0?``W?Z�>�����T��A>��N�j��e>� ���l�ʏ)��Q>m?���=	�>L�E�/�ɐ������?�<A?�@��S�C�;x�i�O��?�!Ѓ>4��>xI9>sU���,��
\\�%?��s\@>{�(?��>iӒ���ž�=���c�O>A��>��p<�u�=
>��o��e �v�)�+\�=�W`>}:_>�?��><��=h@�>(ゾE����>��3>!F>��0?��/?�h�<5&��:c��ْP��Wz>X�>a$�>x�=��f�Q>�$�>��#>ī-�Co��j*�6�(��;G>�)��W�5��r�;c�K����=���=B�HA��w'=�݊?�(���SJ�gֽ�,�;^]:?�`�>(m�q�����6�� ����ľ4��?.�	@���?|�Y�����É�>���?��Y�o�=� >���>\y׾�'����!?�7��ks{���>��x����?m�?���=�I���/k�6��=�2)?����h�>�y�;Z��P��[�u�F�#=���>z8H?W��ܵO�>�hw
?"?]_�ܩ����ȿ�yv����>b�?c��?��m��A���@���>Ϣ�?sfY?fli>j۾gZ�R��>��@?B	R?Y�>�9��'�x�?P޶?��?�0B>>ё?�0t?�b�>��o�ej+�"�k���͈=�_r�b��>�<>�)��=tC��}��^����g��S���b>��=�)�>���ņ���G�=&冽~˥�e�>�9�>�g>�B>��>\�>�[�>���>��:=g�����ϛ��P�K?���?����2n��N�<i��=��^�h&?�I4?s~[���Ͼpը>��\?8?�[?�d�>��S>��迿~�����<+�K>g3�>�H�>7$���FK>�Ծ�3D��p�>�ϗ>�����?ھ--���V��3B�>�e!?R��>�Ү=ۙ ?��#?��j>�(�>CaE��9��V�E����>ע�>�H?�~?��?�Թ��Z3�����桿��[�w;N>��x?V?sʕ>b�������kE�8BI�>���]��?�tg?�S�0?<2�?�??_�A?y)f>ه�(ؾp�����>�x
?*��4xT�E��^,�<��	?9��>3FZ>�d��ii=�Y=["o�����?�o�?y??��������8
����=��{>��%>�U����^4>�I�=EK��X�>O <��~��Y���"��>�=S�2>>�y�q�.���E>��%?�|<N^f�v!`=�b�I�A�&Kt>"�N>⦾�DV?yp��b�ϱ���G����o�8U�?XE�?���?R��<n��&E?���?�q	?���>�L־{���?Ⱦ�2���?�]�"�\�>�0�>`�;(nܾ�&��e���� ��嗽0�h�=
?��?u=5?Xs
?���>�->��Ѿ&--���־|�پ��2� �ɔ �F��eP�Lپ(�N���o>iW��1DP�
��>�ǽ�?�>!;?
I>gđ>1"�>�.[<�ͪ>�s?>��>R:>��>����81p=ĳX�9��) _?\ڱ� �����W��T!?��q?�:p>=�L����d.$��j;?�`�?��?d��>Ds���eI�>��>s�?޹���~0?21O>>���ݽ�W�I��m��+�C�L,��a`>tQ9�0:�V�y�Tȋ����>��$?aLf<*{ǾjI̽�����r�=}�?�+?�(�ۜN��ho�+:Z��>S��1	��]g��P����#���n�m쎿`���̓�mc(��~-=f/)?ᮈ?�G�	f뾀O��T�l���>�(�a>�$�>V��>Ԯ�>($C>����1��0[��p"�S|�rV�>��w?�>%�I?�@<?u�P?�L? �>��>����5��>Mc�;;�>j6�>]"9?�c-?ӹ/?G? S+?)�b>����j����ؾ��?^?1�?�?��?�E����ƽ6/w���w�Yx�+����=D��<��ؽcCy���S=G�S>�#?�}���\�Q&վ���>>�?�?���>}V������a�>,�>e�?
>��:���r��ݦ��r?%2�?[����<h��=ki|=݋�<��c=�����:cz\>Y����<܃����=�l?���I�=qc-���D=�cƽ�e�>C�?�\�>;��>�4��Cq �b ��V�=h�Y>�8S>�!>�;ؾ�Y��X��3�g��gy>�{�?ce�?+|`=�(�=�1�=�I�����T���������<�8?5�"?CT?�S�?K�=?W#?T#>�(�A4��)��̪���?�,?8��>���'�ʾ��D�3�U�?�Y?,7a�����:)��¾��Խ��>�Z/�x,~����D��{��3������'��?]��?,@A�J�6�1s�k����e���C?d�>_�>�>I�)���g�4$��;>p��>�
R?�˵>X�W?��y?�iU?��F>�6���������=f�=��0?(�y?_g�?�j?I�>��M>̨ ��v�"a���(�����J���C�9��c>Ȥ�>�q�>��>y�>�pȽHۼ��^6���=��@>��>�ݯ>���>�6P>3G
=��?V!�>�a��'����&�X��3t�>q�x?$�?�\M?���w��zF�{K���>�Z�?G�?s.?��<���Z>h��mq�$	���?��>���=ģ��媽��=�� ?��?�q^=zd0��3u�	�M�[�?�T`?�-=��ſ[�p���n��n����}<������d�B'��Y]����=�.�����9���\�"���68������훾&&|�S��>��=���= G�=���<NoǼZ��<-�M=A}�<�=�Ww�G;f<�9������⇽(6���*U<��G=����־h�x?��b?^E??�2?���>C��=��1.'>�71���>�Uk>�}���5����F��@˾����|�������j�ܒ��Ë�=�p���2�=��>aF�=]�,F=�+2=��=��C<�t&=6�s=E��=���<�i=�4�=�:�=H�J?O|������$,�6>V�0?Q��>k�M>K�sZ?fe�>	���ߛ��3�{�o?� �?e�?Z��>��
�i��>�Ҍ��g�=�::>���=$�=)>ǾH֠>t�=4�ܓ���3���?�8@>S1?�,��I(ۿ��=�2�=uGA>��A��'3������OU���.?�E��b���NJ>�>q��!��]렼BzQ>v>�i��Z�L�8=8�	x_=�Ld=�l>�U>q>O�;�V��=8�;��3<&u#>�/��"=O�޻�=ƌ�=�A>�>���>C�?ʙ1?	A_?_@�>�p��޾X�Ⱦ8�>�Փ=[Y�>��z=��5>�)�>�W5?�\G?�H?M/�>���=�3�>\?�>�p*�۸n���ؾe����,�<���?�,�?�w�>�q<��9�}��}�=������?Fv0?4R?�u�>�U����9Y&���.�#����t4��+=�mr��QU�J���Hm�5�㽱�=�p�>���>��>8Ty>�9>��N>��>��>�6�<yp�=ጻ���<� �����=�����<�vżƗ���u&�6�+�2�����;f��;B�]<u��;��=M��>�2>J�>>&>�ݾ|�>hi�pH�q�>g�����'�INb�w�}1�N�&��|>>ф>�@ؽ�����?��Y>�`->D��?��T?B�>�:<�3���@���k����\��"�=��/>A�9�*�)��jM�hGA��ӿ���>���>&Ф>Ƀp>�B,�>��Nw=���,5���>�i��4��d ���o�����	����h����7D?�P���|�=��~?J?L�?p8�>�s��(�ؾ$O->��{�N�=m���<w�������?	�&?��>9쾜�B��59���[h�>���^$7�H��1�L���R>�������>Ndƾ�����?���t��U����A��㝾 >�>J�i?#v�?쵶�
���C9�������8<y?)�J?p�>� ?sj?:��H���=��,C�=�L�?=��?���?���<:K�=�G����>"�	?��?��?C�o?�D����>	
���0>h/�����=zc>W͉=?��=��
?��
?�1	?j���_g��쾡����\�#`�<�,�=&�>��>�p>*��=�&z=̯�=��[>xҝ>-��>P�_>��>h8�>��������,?�z>jY�>n!?�s|>��=�>H���<��+��%>���,�z���-���:Q�<��=��d=��u�\��>�~ſ�|�?yȎ>M\��?q߾� ｽ:>���>�.�O-�>�6>]q>��>3��>�v�=�Y�>�(!>s�=�i�>� ��G�!�7�=fj��,�����>Zo���cd������=��y��
��?��d�v�����I�6��>�[I?�Fa�,z��	X�g-����>���=N�D?Y�����=b=�J	?��
>� ������������#�?89�?�O>ܩ>)Z?~?�(6��R0��_�w�}�;:=�}n_�D.X�1,��#�}����}�P�W?[�o?��7?l�<T߃>G��?˧$��Z��_�~>.�5��l:�1��=�!�>�q���uo�%�Ͼ���q'��=W>�v?̈́?-j?�c^��p���'>V�:?��1?Tt?Kf2?V;?����Z$?Q22>E??�<?0�4?��.?�
?�E0>���=�ʽ��U0=����Xꊾ��ѽ�N˽����5=�qz=Kk$��<HO=���<%I�X�ؼ��:n�����<��8=�ˡ=?�=g�C>}	�?�	?��=�C+?D��y�Q�hq����?eN�EP�޻V�L�q�3��k��=>KR?�3�?���>o�<=���T�'�>��>�/�=F�R=b�>t_>q��M�0>�gr>A�j=F��=�ܽ� ��n���*��3-]>T������>��q>�k�`%>����Dys�wXm>��Q�	���o�P�'�F�1�����.��>%`J?B�?|=ז뾌����g��+?=�??��H?G�u?8@?=�kξ%0���I�����Q�>߉�<���&��y����`4��9�<ɔ~>�w��"<Ҿ�aC>���ڽ�<��-v��1�� >��׾'�"����r ���N����=lv>�"ξ��������C��QR?�Y�<C�k�T�<������-=I~E>�Rk>��=»�f1�s��'�>ce�>�~>s+�� �Zt3��ʾi0c>��G?֞k?�j�?��`�g p�@�hT��-���q{<�B#?��>/�?o�V>�v=�²��@���f�Q�J�x+�>��>:���=�ՙ���I���0%��V�>=?g�\>U}?�@U?�?�^X?ۑ?�t�>���>��5�D���@&?ׇ�?$�=�Խ��T��9�F���>��)?'�B�>��?�?��&?a�Q?��?�>`� ��E@�x��>IR�>k�W��^����_>d�J?y��>�?Y?*Ճ?B
>>?�5�0���G��G�=�:>��2?�9#?-�?��>���>)ʡ�jJ�=�(�>Ac?P-�?��o?͌�=��?]�2>��>�x�=>ȟ>	^�>��?�O?ʬs?��J?���>yd�<�ӫ�Ϊ����q�nl]���v;
�@<�}|=���gw��S���<���;UO��n����%�G�B�Q)�����;���>/�\>󎜾�>��Ͼ���h�=��K>ࠊ���:�����m�5>�Kg>2<�>�2>�@S�j">�ش>���>���I7D?.?n�E?����.���̬6�~W>㧃>;6?	�D=9������Q?��\x>+��?�o?�]�=4�O�b?��]?@h��=��þz�b����g�O?=�
?3�G���>��~?f�q?U��>�e�+:n�*��Db���j�&Ѷ=\r�>LX�S�d��?�>o�7?�N�>/�b>'%�=iu۾�w��q��h?��?�?���?+*>��n�Z4�Y������ӹ_?���>WԠ��?��~��0׾�Y��6����Ṿ�h��1�������^�QG��ι��G�=�_?��v?@Xt?��_?�|��*�g�9]��)|�ӷJ�T���j���I�jLE�Py8�n�N(�
�Ҿ8W����=����	1��ݴ?�k-?���O�>����xC龲 ξr)1>a	��G�#���==au��{O=��Z=q�����S�3����I?� �>%��>ɗ:?��X��B�ى2�T�2���7B>鮧>i1�>ޙ�>ł�;�A�6������;�P��l����g=��o?�h?�R{?��D��XC��?���O�(d������{>��W=��>�^3�2oa�U�!��oP��B}��N�����,����:��;?�p�>�2�>�X�?8��>��0žjrҼ��̾�$}��s�>0�l?�+�>H�B>�4��� ����>^�l?��>k�>����g!�A|�z�ʽ�S�>% �>RP�>�Kn>�,���[��b��rp���$9����=�.h?����b�p��>��Q?��9:z3<� �>_�r��!�m�򾘽%�@
>{S?���=��<>�ažX|�8�{��z���`)?D?�b����*���|>M["?���>D�>�j�?��>�[ľ�s��@�?�`_?��J?�qA?�|�>�y=S���[ɽ�5%���3=�-�>|�Y>j=j��=d��
�]�����VI=5+�=�ͼeU�����;Jg���NV<���<�o3>�^�E�"9Ѿ�M,�\B����t*^��_���ٕ�����8M�凑���*�Pn��m �o<��1z��}|�)և�+�?D �?Y���Qľ夿�4��FҾ3�#?e!��VL���½i����A���ܾ?�ܾ�Ȃ"��[Y�~�g��J'?�g���zǿ����=�ؾr�?9�!?Աx?�����"��6��T*>Y=�\s������ο�̕�nwa?�>tI���=��wq�>]Ն>,�\>�p>3ي��⡾��!=O\?0e+?��>)5m��ɿ T���g�<T�?y@}�A?*)��z��E=.u�>p�	?�6B>�2��\��U�����>m�?�~�?p�@=�~W��(�lKe?7�M<�uE�C �G�=���=5=uD�w�H>�Ǒ>;C�j�?�R~�D�5>ل>C�)�}��I�\�4'�<7�^>�DԽ*���Q�?�8�^�=�X�%�(i�8ƌ>�3Y?F��>]4�>N?
�u�>zɿ��:��?&l@l�?���>=p�Y�>��ھeSa?�FT?�+�>��)��ZR�rk>YH��`���� ߾	�+��f�=.��>w��>#�o��
�0e�:�\���d=�#�,�ƿ6�$����`� =�?-[����%���`V�����Vo�4c轠
j=��=�\Q>'�>O
W>�Y>a�W?�k?a��>��>�����2�;���n	��0���V���l�������߾�h	�)�������ɾ�5X�L�-=h�U��1��9!C�A v�+$4���F?��=�2�����Q==K������'#)�����j��1�+��v|�h��?\u@?<����������>�\����E?i�ټ\hɾ^1m���k>���E�@��x�>��;���V*�Ճ]��z/?�?0ҿ��ᐾH�>�����=K-?m� ?.`�<�*�>��$?e�3����k&T>j8>� �>��>S>Z��I�нϚ?'�S?N	�S򚾇��>���i�}��
w=�� >�[5��Y�[>�L�<�#������N��cq�<-�K?�.>T�$����p����q>!B[=�DK?m�f>y��>1�K?�zN?V(���n�2'C��۾7Z�>;�T?�_??�h>y���W��!��S4`? n?���>��ھz;�yF!�!3ᾫ8	?Sz�?�??�d1�퉿Y����2��/L?��o?�s�l*����,�HH8=��>m��>%��><���^e�>y�?��4>wՄ��Ŀͻ5���?M��?�'�?V��q�&�z��>?#Y�>-֯�ޝξ�ga�x��V�=�(�>�h���,�w
��1���?2�U?��?d�"��/��=ɏ��rV�?��?�u����d<a�Vl�r������<H��=����.#�����7���ƾX�
�9Ȝ�������>US@�A�cB�>*P8��.�6IϿ0���=о�q�e�?�5�>0ɽ�����j��<u�!�G�=�H��y���ۨ>�(>�x�n�S� N��nG=�4���*?�3Q=_�>ߒJ�v�Ǿ��׾EA��I��>�[�>�C�>*<N�ڒ?����ƿ8���E׾N^?��?�?i?��?�>1=[aJ�h;W���齎�L?��?DAb?���݌�N�&��j?#��h`��4���D�iiV>�3?M��> @-�U
=�c>%��>�Z>/��fĿ����>���|�?�g�?�6��7�>yk�?pU+??W�P
��ߪ�L*�֘0�@�@?-^1>�w��+�!�;o=�|c��g?^�0?�A�l���g?	*I�tIA��E>�0����p>�~<�rq����>A���E������w˱��¬?�@�o�?(#q��2� �?�k�>�V��f�X�y�`=�1>g�?�27>�����?c�-�|"���:�p��?S�?�4!?�����I��A}T<P�n?��>��?)��=gl�>�s�=����.�Hn#>H1�=*�>�Z�? �M?nO�>�e�=�8��/�o[F��HR��%�d�C���>}�a?e�L?�:b>�F��H]2�X!�JMͽLO1�g��ID@�e,�l�߽�5>��=>>��D��ӾC@2?y�^��Կy���ip���H7?\��>�s�>��达�=c�=�^?���>�ᾅժ�L��y��6צ?'��?��>˱��9���+�=���>Iޠ>��Y���+�Ib0���c>�W�>��:��5����z��x:>�.�?�5�?܏�?"�[��?�A������Z�m�e��K�a����=�E?��q�>ze�>P�o=[w�\ݪ�P@k���>4��?DE�?���>��d?Y2j�j�5��ZL=��>xb?�?D�'=g־��d>o�>����1�����jp?2U
@��@�gc?�\����ؿ,��0��������=D�=��1>��߽J��<ѾC<���%C���>F6�>93w>mAo>��I>�u->Y�2>��b$�Q۫�������9�����
������������W"�Y�ƾ[���k˽�-����D�]3�������j���[?&�p?��?�f?dH��Fy={Kɾ�/I�y�0��>]�>#�?�:??{�?=�̾8ey�u���z��nO���>��>D>#�z>�\[>k͊=9E�>���>�X�>^�f>g�K>�S��z��{�=�Ɨ>�7
?�A�>65<>c�>�δ��0��.�h��w��!̽ �?�}��@�J��.��6��<���>d�=Ea.?�v>����=п�����3H?>���H'�{�+�J�>2�0?�_W?��>���T��8>θ���j�%^>�  �V�l�ގ)�$Q>�k?�`>�w>��1�6��UP��^���w>�5?������<���t��IH���ܾ��K>��>��,����8ږ�Z}~�t�e���~="�:?��?�Y��ئ���z����-�R>��Z>*�=-_�=z:N>�"c�_�ý9�H��@)=�i�=�c>y� ?�- >=9={x�>
ʾH�9��E�>��>H,>
D?��&?`����Y����l�K�0i�>٘?�t�>j��=-�R�@O�=���>:av>����j;3���M�F��>����y�-�����;s�P����=Z�f=s�k�U�d��=�~?�~��;㈿A뾔m���mD?�+?a�=5fG<�"�� ���J����?��@�m�?e�	��V�p�?6@�?8��n��=��>�٫>zξ�L���?�Ž$ɢ���	��$#��R�?K�?�/�4ʋ��l��7>�]%?��ӾP]�>~������ޞ����[���=J��>�H?����rN���iD�w�&?�h.?F������ϿF���_�>���?�?�؇�eԡ���f��P0?�b�?sZi?GR�=8��v�h=3g�=��1?�$?�M�>��<��z�ɠ�>���?u��?Q�&>'�?�x?� �>������0��浿Fn��ur�<���:ndw>ţ�=`f��f?���Q����^�����L>�%=�o�>R�ս����8v�=��x�ƞ���p��>݂�>�T>��>�?�s�>{��>��l<Ѕ�n#t�����w	L?ވ�?�	�˔m�6��<���=C[��?��5?��Z�Ҿ5��>�\?qU�?��[?4�>~�R2��=t��龴�k�<��O>P��>��>e(��n,K> վ��H�:��>��>�#��́پܑ��X��氜>Aj!?�O�>�5�=ۙ ?��#?��j>�(�>CaE��9��X�E����>٢�>�H?�~?��?�Թ��Z3�����桿��[�t;N>��x?V?sʕ>b���񃝿|kE�9BI�;���^��?�tg?sS�0?<2�?�??`�A?{)f>؇�)ؾo�����>��!?���A��M&�D�`?�Q?b��>,%����ս�kּ���{��L ?Q(\?O@&?����*a���¾�(�<U"��lU����;�E�a�>��>n����=�>;�=EOm��F6��f<�d�=�~�>�=�.7�z���l(?U����������<�p�e�2���>Rk>YG���T?M8��]�Q����ˠ���k����?�1�?C�?�޽�e�w�L?%�?״?z��>ƭ��`����������G3�ͧ�JV=���>1�><�־�����������\��i��F9U?d�)?�E5?v?�9="����U�Y�X�������ы�L2�����/8(�ڋ�����ʙ�Pg<�j\���Þ����>j0��K�>���>_~>�R�>���>����'��>��>�$�>��>��=��ü����!���D�:oQ?j4���&���q奾0B?�d?
X�>��9�z��6)�@"? ��?6��?�h>C�g�E8'�|d?�N?´��?�	=�"r<��ټ.q��yO6���ϼa�A�q�~>ˬ��X4;�e@N�z�O?,C?��;��ʾ�e���ڡ����=1O�?�R*?n�(��Q�j/p��aW��>S���-���l�����O�$�bo�h����K��������(���-=�>)?��?�G��p�j����k��?�&�`>9�>Xp�>V�>��A>l	
��>0���]���&�������>��z?C��>`�I?C<?@xP?�kL?h��>/c�>D4��[l�>�;� �>��>�9?i�-?80?�z?�t+?�2c>]�������ؾ�
?T�?�J?�?�?2ޅ��sý�f���g�D�y��~����=]�<"�׽�Eu�8�T=]
T>>{.?۞վN/�*�[� ?�S?1�L?ez����� �>>�7?on?&��>l����{s�H@���;�>=�?.Գ�}�[;xa>��}�	��<f�佋��=Ge@�>�P>�^��+ć���=q�	=��=�.�=���:��	m��2�;O��>E?���>!�>z���l����p� �=��X>�HW>o�>Ƞ־K���u���gg��{>�֐?�K�?�_=���=���=ǒ���n�����X���Z��<W�?�!?C�S?g�?�=?%�!?��>E3�Q���L���������?h!,?Ƌ�>E��P�ʾ�񨿉�3�B�?�Z?�9a�����<)��¾��Խ��>9Y/�/-~�}���D�������0x��$��?��?A���6��x辻���_��V�C?�"�>�Z�>D�>�)��g��$��3;>Q��>�R?k�>��O?l?{?k�[?�lT>�8�1���љ���2���!>�@?b��?��?Dy?2n�>m�>��)����V�������m݂�;W=�Z>r��>�"�>��>���=��ǽ�@���>�r�==�b>���>���>8 �>!�w>�R�<٧B?	1�>���������O�Ͻ��?��?ޮ4?p<�<V8���L�KW�d��>�%�?���?~�/?rI��8W >d⌽�r��Z퀾��>�`�>o�>t"�=0Ș=F�;>+�>��>�kM�t6
�]R����<e�?�6B?;bp=-Yſ$[n��Fn��$����;����z�i�!q��u�Z��ו=�m��7������[�����{���1���d���Ԁ�Y�>}�=�4>�`�=��<;=�,�l<��:=g�<��=j�q�ڬ�<�Y'�һ~���%�����&<��[=i_�:v� �%�{?h	Z?GQ?�$H?1<R>ľ�<��h�L=Ӟ~��[?��=���:�|����H��rϾ0$!�|���Y9��r���UO>ꑽ#a�=˽Z>�}>UW>���=Ґ�=�~M=jH�=�:�=g��=�=,Q�=�I>��>�&>��q?2�f�䴅�m$?�h0�\�?p�>>�n���!a?<�\>\s�d�ǿL�����?�b�?>�?���>�ĭ�_�>�C羲��kX���=
,!>fk�>� �\_x>/g�=8�"��5����Y����?BN�?ˡR?<���Vr�Ν�>�9>��>�N�t�,��~���Y�57g�J�'?6�4�o���/�>X��=܈�f�ھ���<�G>��=k޽�W�=~�=���dPQ=ZXh=7��>]�R>�t�=�ƽ���=��==�B�=pl_>����>��o��=�=��S>y�:>��>��?��/?iud?�е>�`t�0[Ѿ�y��ѳ�>���=`��>9d|=�0<>jY�>�-7?b�D?��L?\�>>
}=�A�>IX�>��*�!Fl�Ҧ��K���Y�<�ƈ?Q�?��>��;�I�����=�hy��?'(2??�	?2ܚ>�U����2Y&���.�?�����5��+=�mr� RU�����?m�6�㽦�=�p�>���>��>!Ty>�9>��N>��>Ǫ>�4�<�o�=�錻;��<$ ����=����n�< vż�����r&��+�������;<��;��]<,��;�p�=�w�>G�>�D�>�X�=Q���s.>闾y�L�㹾=�����B�FDd��}�_�.�&,6�MA>AV>󇽻/��ʌ?��W>�&?>�a�? u?p�>���վ���m�c�`�T�V�=�n>�X?��;� `�׀M���Ҿ��>�ߎ>�>�l>�,�A#?��w=F� b5��>|�����)��9q��?�������i�KҺ~�D?rF��՞�=S"~?6�I?��?"��>�����ؾ�;0>3H��F�=���,q�)l����?m'?8��>����D��˾�޽�}̷>�H��'P��Ε���0�N��d����>M����	Ѿ�>3��r���Տ�c-B���p�E�>�8O?�Į?/cb�=���O����O���0?3�g?��>I~?�?���0�y|�����=to?|��?�:�?�u	>��=D���o�>ܐ?���?���?	�s?v5@��]�>���;�� >,t��s]�=̜>C�=� �=E'?:�
?.?$֝�9A	�����1�Ħ_�`��<�=�#�>�-�>/p>�H�=��d=�͠=�[>{w�>Ǭ�>(e>���>���>����u�
��P'?Y��=^��>��1??�>��U=����O�<�N��B��,������^ݽ�B�<����k�8=D����>��ƿU�?��R>ƭ�i�?���a�"�>V>�V>u�ݽGq�>�!J>�{>�e�>�ڣ>�%>��>pR+>W��Wo�=,�����6Xb�t������o��>����P���ӻ�����S ���O۾3�w��4���5��׃��ŗ?f���Zb�R�5�>����/?���>;�!?& y�B�i��=�n?~��>2nȾ������S�q�?� @s|�=���>��e?V;A?�H�P�����m� t�t@���{���f�����������P[��G?��N?��?mN=�sE>~�?I2�,u��{�>�w(�ԏ1��><���>	�t냾���Ҥ��;	�m��U�Q?�?�|$?Ef���f��5%>*	:?�0?Ét?)�1?z�;?̀�I�$?��5>uK?7�?1�5?��.?9f
?��/>M��=�U���-1=���0ˊ�˛н��˽aK�|u3=�Fy=S0�l�	<�/=��<��I�ܼ0�;�v���v�<;=K�=��=�	�>6k?��?���>U�:?-�D���J��;ľ�2?�zM=����G���d�澊�l=z_?)&�?�I?��F>�0?�a�<��>�%Q>�MO>,;k>L��>�����a�1��=��!>d>L�=L����$��v�����E�<R>�w�>C��>}�9>�'�>�־q�⽗C�>Ӿ8������v�K�:�� U�;?���?*�@?g ���D)�;g�Ђ��4%?C��>�L?�v?��z��t�!R��ى����<d�>i��L.(�
����٩�:�R��{=�|">�U��_���24m>~S�`Lξ�{a�AA�fM־�u�<�=����=��
�⾊9���g >�h>�S��R"����2���CG?�� =[���\�p��V�����=��>ԩ�>ڏ��",��6�D�.���F��=zi�>�mG>��~:"��B��0��\>ȯJ?�]m?Ĕ�?�a�������W��A���$�wT>�<#?a��>P�,?��>*��Ǭ�H�2�w�c���3���?�+�>�_%��`�+Y��i5��q:��K�>�?H�4�*�3?י!?��>#�e?=2?8J�>`Mx>���Ω�`V%?�?�̡=?�̽�ze�!v:���E��O�>��)?@�^��n�>.�?�h!?��%?��O?��?�6�=P��v5H��P�>���>��U��x��q>e>Z�Q?ۨ�>��T?��?B:>�09�����)�۽V+�=��&>�6?
�#?Ǌ?k �>{��>3�����=`��>�c?
1�?��o?{�=��?`-2>!��>��=���>���>
?7TO?Q�s?��J?P��>���< 3���:���0s�>@O�'Ɂ;��H<i�y=
���"t�NR�J��<䝴;�ɶ�ԏ����D�D��n�����;r�>~�8>�V���w�="X��Ͽ�M->�M>����H��-R��~x>���>Z�>c�f>֜G��5�=8�>���>Q%���$?Z�??$v߽An�J� �=�Q���7>�31?��=�vt��.{�*��=�,�?e�g?	�<���-���[?�G_?�٧�Q�!�����Ǿԑ	��]Q?�C?JΆ��1�>�kf?hׁ?%�?x�B��cm�X#���Rg�~þcs�=q>h�%�T�r����>tUg?`2�>�r�>��=��	��h��	:�����>^�k?���?�i�?��$>|�`��_ۿ���k׃��Z?F��>BƎ��?���<��׾Ů�H��xu���\���ڲ�I,��4����� ��j4���C=_�?)�t?Y�j?da?EY��c�x�i�yr��KR�vO�����U���A�W�@���Z�v���8��7�q���>�Ͼ?H᾿��?!W?�ܿ� ��>�ޑ���D)徏7X>T�e1��2�>	�����=�˼���v?v�>x���a	?u�z>E��>^!F?�G��P�cx¾��I�x����=vY�>�@�>��>���g��"�����ų�e�D��0c>%�d?��J?�%m?�/��M3�V6���(��7��񩫾�=U>H�>Ur�>�$I�;�A`%���=��q�����A��O ��=v�2?���>R�>~�?��>W
����.�{�\[.�n=J߸>)#g?���>#�y>�N�Q�����>Ap?{��>�S�>\v`�=�!�4ꀿ�8ͽ8��>I��>P&�>��\>t���V�Qr��Cȉ�@�.���=�I`?� ��V�J�}�t>�Jb?m���N3�<���>l���Er,�x���,���b>]�?�]�=w��>�۾%l!��U��NTk�'K)?P?�ؒ���*�~>�"?�j�>�5�>�2�?�$�>�Yþ�%���?�^?O>J?QMA?9�>Jt=Z&��	bȽ��&��3,=r��>��Z>��l=���=d���_\�r�
�E=|��=��ͼ�@��ڃ<�յ��CL<�m�<}4>�lۿ�@K���پ����?
�n䈾���� g��f��\d����,Zx�����&�V�:c�4����l�Ά�?�<�?�}��T,������z���i������>?�q����<�P��4*�����V����a!���O��$i���e�P�'?�����ǿ򰡿�:ܾ7! ?�A ?5�y?��8�"���8�� >pC�<I-����뾬����ο9�����^?���>��/��o��>᥂>�X>�Hq>����螾�1�<��?5�-?��>��r�0�ɿb���¤<���?/�@�cA?�)��x�p�L=P �>K
?�@>'71����*������>#�?5�? �H=y�W�8���e?�e<��E�M}�����=?G�=�=���S�I>�'�>����8A��<۽z+4>�ʅ>������^��<a�[>6Yؽ�ᑽ��?��J��M���1�]F��Bn>��c?V�>7�>7��>бe�TQʿ��7��r�?@߅�?���>l�Ҿ�,�>���VYY?�zJ?J��>�7�mb��A�=A��O����/�<�d�
>���>�E>o�m�42�*��*����>i����ƿN6%�s���s�<FM:��_��Z߽e3���1U�4V����m�|���\T=;��=��Q>o�>0[>8�X>��W?�k?e�>�>��ܽHf��f-̾�/A� ���E�L���	��&��Zp�1x߾��	�-������Ⱦ�=�!_�=�KR�ؑ��7� ��b��yF��-/?O�#>��ʾ�M�F�6<�P˾�����އ�������ʾ�0�y�m�`؟?f�A?y˅���V�>�1���󂵽��V?����������N�=H��^9=P��>�=���83�<�R�� 0?5�?�_���搾�r(>ȴ�3	=�+?"?3\<��>��%??�(�o9�F�[>3>���>���>�>b���:ڽ3�?�	T?�G�C����>S྾��y��#^=Г
>4R5�Oؼ][>�8�<� ���C��S��9 �<>�/?[�J�A�D�|�6��*�S2�>Z�=��Y?���>Z��=�f?_�:?^F��{/�]�A�����6�}>sX{?[�Q?	{�>�XQ�[�¾_~����U?o�C?���>��辬ś��}$�̬	�Z�>I��?B(F?�����w�a��������c?G�#?J�p��T����%��������>��>Z'?	,'�؄�=�C?yy��o��Dǿ���-��?��?�Z�?����#���<>�??��>���c��V@��ܤ	���<�C?-���z�X��ΌZ�S)?c)v?D��>|�[�4��&��=ٕ��Z�?��?#����2g<(���l��n���z�<�̫=7�^F"�����7�X�ƾ��
�c���M⿼��>+Z@U轧*�>�D8�:6�	TϿ���[о�Sq�l�?o��>ԡȽo�����j�GPu���G���H����o@�>�5>�W��U���ؚ{���7�/���:�>��P��>�rH��ϲ�Uˤ�(������>��>Ϸ�>gR��#���q �?E���̿"����"�Z?on�?���?z�?S��;�w���u�����F?_q?!�W?�o-��H`�A�!�V�g?�/��h_�s4�B�E�� l>��1?�X�>v	)���E=�"#>.�>j�'>w�-�K+��U��l����?b��?��澎� ?ގ�?��*?*�Oh����+9�C�ռ��<?/,>&����6'�w�@��ތ��N?/y2?8^ܽ��#�O��?��X�{�R�wK&��O-�"0�>��>Ny���>_$>��m��Y��I"�����?�@���?60��(�2��a�>x�>���� e��ս7�>���>��*>�|��F�>�`�����^ۥ=Z7�?�*�?��?n=���ߦ�DD>�h~?���>m�?�V>��>3�K=���� �T��>b��>�4���E)?�U?�Y?��.>6 ��� ��4��F���s�C��f�>k�>?�?>?��e>��/i�=O%�s�
��ov�Ɉ|=����0�>l���$F*>���=k�=�d� �¾���>�?�K�ٿ�*��X!�(�*?�'�>X�>=��z������.�c?Ț>-�%��.��\'��е7�!��?��?���>�R����G�=8\>ׁ�>P휽�%<�n�@��=�;?�������N��j�>O8�?�[@s�?��b�ޅ�>M;�Q����s�fj���[����=��O?i������=���> 5>A�r������iR�&��>V�?Z�?�ױ>�<^?�+V���#�(�=3Xy>�nP?�,�>
*���E�&��>��?��)�6����׾I�b?}$@$x@�qD?py�����mG���Mо�lɾ�gm> W�=�bP>�x����=:L��NN>=�|�=X�)>�Qg>b��=���=�b0>;4X>֑�>Ϸy�p}/��8׿^4��������l!��*q`���L�������g�%�������s���\���?>�$�=�=D�]?�TI?�YL?�>fjq�U��<7\��޹G>�93��U0>��>�)?O<?�m?�r=�4¾��_�dC��QJ����2� �}>3X!>��>�;v>U�>�/�@>��t>׻�>�}�>�B�;J�=�8�9�z=>;��>� ?���>�C<>>?ϴ��1��k�h� w��̽1�?r���W�J��1���9�������h�=Gb.?|>���?пh����2H?%���y)��+���>��0?�cW?�>��`�T�:>0��Ǧj�%`>�+ �Xl���)��%Q>rl?�Ic>*�u>G�2�5�7���O��H����}>9p5?���i�8���u��H�Xݾ�9N>R�>[!>�Ix�F���|��Zg���z=-�:?�[?�洽�B���v��ڝ�TdQ>H�X>��=/�=KL>��f���ĽE�E�2=�h�=k`>�7?�,>�V�=���>�y��SpQ���> �B>=-->��??D%?�4�Ꟗ��"��S|-�	�v>��>vŀ>�> �J���=g��>��a>g��eX��95�aI@�+ZW>̈́~�Q^��v�b{=f�u�=�N�=� �Ol<��(=��~?�=�������R�9����xD?ʐ?F|�=�&�<��"��������?��@���?ԡ���V�j0?F�?�������=�}�>�g�>(�ξ�@M��?|SǽV���q	�1z"�!�?�Ҡ?�-�o����.l�Q>%?�Ӿb�>h���Z�� ��b�u���#=���>�8H?T����O� �=�|w
?z?�f򾔨��;�ȿuv����>��?���?��m��@��@���>z��?�gY?�_i>Dc۾�hZ�B��>�@?R?��>G8���'���?6ݶ?��?�H>B��?L�s?���>1�w�GX/�6.��������~=��`;{b�>�x>����Y^F�]ѓ�]d����j����0�a>�$=���>;�2*��%�=6$���1���g�[��>�9q>��I>�c�>�� ?�P�>Ј�>57=\���1ހ�����mdE?�?����Y��*輀՝<��}���?��6?aq�����̲�>�_? �u?�eS?���>��������Zÿ�y���<й+>���>�f�>��;M�b>�SӾ�m�p��>k�}>].:=�@�����6R�����>�q(?���>��=�� ?�#?�-k>�l�>�ZE�
V���F�z�>D��>�K?��~?�?GB���3�����꡿��[�ҏM>�x?�w?���>􎏿 ����K�cxG�i�����?Zg?�8�m?��?�n??0�A?	�f>n9���׾�í�wQ�>�!?���A��I&��x?�J?9��>w���ֽ12ּ����n����?'\?�<&?ɠ�h-a�þ� �<k�"���V����;��C�B�>G�>ݒ��c��=�>���=>m�S]6���f<�k�=��>�$�=M&7� e���<,?O�G�܃���=��r��wD���>�KL>��G�^?�j=���{�����x��	U�� �? ��?vk�?���h��$=? �?A	?"�>�J���}޾ڔ�MPw��|x�Xw���>���>�l�z��������xF��)�ŽwT���?'y�>�$?��?�-~>W��>8?˾�%@�:]��>&���3o��k�NY�q�����&ⶾ爄�^?ٽ��˾ [�;@r>���^-�>U��>6)�>��>���>ÈػJ�Z>g6O>���>eW�>��<>���=�su=���<���K?6˾4>,����JϪ�ߵR?��g?z|�>$�;�y��*�۾"E2?�Ӗ?��?&/B>��m���%�p��>�i?��s���?R��=��`�"� ����z!��p�=x�½�\�>������"��H��㥾��	?�; ?6�0=;��-9��uܾ�N/>7c�?��V?����{[��F�6q�Ŝb�]� >޹J�;&��?��M�_��э�d���8-0�`�=��2?�eR?+�d ��3̾����P�C��>0�
?���>��>��>��ܾ�:��\`�y_*�7){�ˈ�>3L?踈>�J?Y�:?ctN?��H?'�>��>������>�;���>��>Y�:?�-?O{.?rA?�(?3#Y>h���>���χԾ��?29?@�?a_?��?K����Wͽ5��(̻�����:��(�=�9�<Uq�Y�{�J;4=11M>��?hd�B�_��#�c�>�C?5-?�W�j��1�����F>��?e�?Ğ>�X)�2���)u��{�>��?�n<��=��2>}F�=���ڪ==ճ1>��=4;�=p7=p�<�#>8bd>�A>� =��I�S�8����=mZ�>��?,��>!F�>�#���� ����>s�=�3Y>�;S>��>'Pپ�x��!����g�dby>w�?v�?\�f=���=��=�v��6��j���꽾��<l�?[?#?�PT?��?��=?�e#?��>��,Q��c��9�� �?�",?���>N����ʾd���3�~�?Z?9a���==)�B�¾��Խ	�>�V/��+~�B��9D��������lp��8��?=��?�A��6��x辮���d����C?<"�>$Z�>6�>H�)���g�O&��5;>&��>b
R?��> P?�z?,[?kR>�9��뭿7���K��OL!>$@?�ǁ?n��? �x?�T�>�M>P�*��Zྕ���F&$�AM�i�����U=;�Y>0�>1��>�ߨ>���=�Gƽ�����'<����=Egb>���>�>6d�>F�y>g��<��G?���>�^��U��B�����=���u?:��?_�+?�k=e��,�E��K���G�>yn�?���?k5*?��S���=��ּGᶾo�q��)�>Vݹ>4�>���=�}F=�a>#�>1��>[&�_�,p8�tEM���?�F?���=�¿s�M�$.9�8>d�r�u=�lu����43���(�����=.���%R�pi���'��lr������ݶ�zT��pL����?|��<�j]>��=r�*<~$��	=-�t=u=�<����3H��H�=@�y�36���ѼF*�=oE&=$/
=%}�<�پ�}?�-I?F-3?u@?tb>��>�Y���ҁ>��!�F?\�O>>
мuZ����/�j�������E�߾�tӾ��`��ۣ�,n>�Hr��>V�>�/>�U�:LҾ=�u=��=`��<i�=a�=�Џ=�a�=��=!�>�A>T�?�r�7���BA2��!D��%?\��>�>��޾��?�	�>�d������Ӿ�}?���?c��?��>�z��Ɨ�>
L̾h݅�6ٙ=��=gt�=���>�̉��J�>���>�Y!��W���w��c��?T��?�g?�7��wLݿ�w!>����o���^�}E:���̾�Y ��v����Z?�%�)��[_�>��=8/$�� ��#<�G>���> ><N�4�=>�W��u>��=3n�>�_�>�>w�0�=��=�H�=�;�=�~k>�]5��Vw�S��?:/={�=9�>�>�{�>'�?�e0?Sd?�9�>�5n��-Ͼ�6��2�>!�=K%�>���=�JB>>��7?�D?�K?tr�>s�=h�>��>܋,�|�m��=��ҧ��)�<���?Ά?�׸>q�Q<AVA�<���]>��ŽHu?�X1?#v?�Ԟ>�U����;Y&���.�S����<4�P+=�mr��QU�$���8m�/��z�=�p�>���>��>KTy>/�9>��N>�>��>7�<�p�= ጻ���<� �����=����<�vż���x&�G�+�:���c�;o��;�]<��;�9�=�A�>~?>���>��=�����#>b+����X���=����dxI���c��p�((��K.��'>)�">�u��������?�K>R�F>�
�?pi?YN>{�ܽ��Ⱦ8-����(�Hu�$]�=�!�=V�_�C!@��Z��@D��vվ���>zߎ>#�>P�l>�,��"?�>�w=��eb5�m�>�|��d��)��9q��?������Ki� �Һ D?�F��X��="~?�I?G�?���>q����ؾN:0>�H��,�=V�Y*q�j����?�'?���>�쾥�D��J̾�c��cŷ>�hI���O������0����G̷��y�>o�����оt#3��g��N���^�B��<r�8��>��O?[�?Qbb��Y��hVO���
���o?�xg?��>�D?�=?�!����.���<z�=�n?)��?�?�?p�
>L��=yQ����>.	?���?W��?��s?q�?�pt�>U7�;�� >?}��$�=u�>�H�=���=<j?��
?J�
?�8����	����g���^��R�<��=8��>Ae�>��r> ��=J�g=X��=�:\>�ʞ>��>��d>T�> W�>0U���H
�6"?C#�=�]�>�_1?	��>�j=w8ƽ�f�< �U�ʦC�Cl:��ǽe�ս��<��o�)WS=]5�,,�>�`ĿZs�?�C>� �ۦ?f����R��T>�]8>�������>��M>{�y>���>h��>$N>�F�>69->�HӾo�>|��^a!�"+C�i�R���Ѿsz>����`&�	���o��k;I��n��Mg�j�e.��5<=��ֽ<�G�?������k���)�:���Ғ?\�>r6?!ی����>i��>bɍ>K�������Ǎ��hᾠ�?5��?Uy]<�� ?��]?�+?�,���a���_Y�~�\�y�n���7�bZ|��A���|��0þ��Z���e?1r?�#�>e�a<��>�u?���`�����>��	�k�X����=le�>��|�Ĺ��%쟾7����+�驽��h?���?L�D?V�}��3n���'>)�:?�1?%3t?6�1?�m;?�����$?8s3>�J?��?�N5?)�.?��
?S�1>�t�=�g����'=E���"튾��ѽoDʽ���Ri3=�O|=>�}q	<�v=<��<�4ּ@�;�}��X��<��9=��=��=�V�<|Ix? �7?���>�ɂ?P2��ST���f���?4?�K�>[� �(���UӾ��K���l?Þ�?�>?2z��U�3�x�P�r
>J��>Na~=_Qe>7�f>w�&�'7�<T	�=)�f>=��>V=3>�@�p�%g0�8H⾚��<8�>Y��>c"u>ٲG=� a>��U����H�>��˾�|ܾ�j/�)vd���=�Rfg�fG?Ъj?��!?�1G��'���\�O-�� f7?�g*?V\�?���?
7>c����E�{���4�=v��>�l���E*�����ǻ���R�O�=d��=Uо�8��!\>������q��WG�����e=II
�Z�< �5�־�z��>Ԃ!>	����������7z��ăI?�g}=�U���T�|���CJ�=rg�>�>��I������<=��C���j�=e �>��?>o>Լ|��E�3� ���W>�PI?q�v?p��?�&.��d��&�.�&D��[��i�=��? ׳>�H?���>����IP��:����M�H�q��>>�M>�Xξ�Ci��O����4��	�>{
?̕�=�.�>C�?�;�>uzR?j?�%�>D� >"�=��˾B�$?d��?���=dԹ��Q�=�%E�,{�>�J+?=Q�ϒ�>�r?�� ?�-?�K?�!
?�&�=,@��D�" �>���>��U�����u�b>�+G?>?�>9�W?hy�?��$>�X5�EI���
Ͻ�I�=qn->`�0?��?m�?�T�>��>{��h^v=���>%�c?X�?}o?���=v�?��1>lY�>���=O�>���>�?A�N?hMs?�vK?B�>|�<����m��U�k�(B���;�Z<�qu=DE��>x�������<�[<#w��
�z����O�g߫�^�Q<m�>��>�!����>c�ɾ�Ax��q>
Q>�?��ڍ_�]���Sc>���>�2�>�' >�,*�Zƅ=C��>�!�>�/�u(?�?��?j߽k�X��󾈱��� �>.�X?�n>Wc��ʖ�o{� G�=�w?�H]?������)��a?��]?��[D:�I/¾��m�i��1Q?��?��N��m�>�`}?{r?�?�Od��Fn��G���Xb�Hyv�6�=CX�>9C��td�h��>K6?7�>�-f>��=v~ܾ�w�#��/�	? �?�;�?G+�?�� >�5l���޿2��#ć��uh?B��>�ȓ�j�#?1b�;���l��Ԇ���׾V˱�H����ƃ�����qy��ٌ���x�=QQ?0�n?N�?sVN?��
���U��de�y�t���Z�%$�H*#�S�O�g�J���?��LZ�� �D帾$�n��u�=����?���?4�'?��-���>=������о��A>�Ҟ�'.�N��=�����LG=�V=��j��_2�����o�?+;�>��>�9;?)\�,=�v2���6�����{2->�.�>�v�>x��>l���l)�����þ?���L�Ľ��>��x?��b?��?�g�i����v�4�NS���+ھP��=��>�?�o�e(l���3�	B�B�y����*`�+o���C��
O?S�>���>�ت?�=�>���\��똽�ھ2��=���>2 Q?��>��=ef�����X��>]p�?��?�>8��,���z���Xn���>L��>~X�>Sl�=5�l�){A����Ba��s�)�"�=�5C?����6��>y�~?l�r����=���>��<�t�1��'$���򽻲�>H�9?q�=�D�>�1��x+�$���н*P)?4J?)撾��*�R8~>.""?�}�>	/�>�0�?(�>doþ-�?��?��^?@J?�QA?�E�>��=P���:Ƚw�&�A�,=r��>��Z>'m=F��=��7q\�vt�
�D=�n�=��μL��5�<扵��J<�{�<��3>��׿�;�Q��D��:-�W2�zq��!�BG����n��R��{����0���<ݺ
>ྚ��M�X�z��@��L��?"��?I9���M���Ї�}��\���e�>�쉾��j�Y�@��b-�����<�F����S���H�l�P�Xj]���'?V����ǿ"���� ܾ�?I ?�|y?�<�ާ"�f�8��!>}�<�0����|�����οfy���_?���>x3�&��{��>�ɂ>�CY>d�q>��������<��?��-?Օ�>2�r���ɿ�n��r��<h��?�@';G?]�A������K��r?���>�'>R�A�
� �8��O�>_ʠ?t.^?6���M�P���6=2�i?��d><:8�?��<�"%>K	>ZJ:��ὰH`>�j�>�;����5��»�=Q��>L��;
�Žz�����F9��"`�,GS��7�?(^Q��EV�@J'�^<}��O;>|�h?���>�#Y>+?�h[�Kʿ��H��u?�@Љ�?�c?jk־<��>U)��O?ϟ.?���>�,%��Qi�B�=�Gk�>�������h����='��>ORd>5D�.��U�(�Wh�;(�>��1S��:�#�\�>�������w=�3�<ɮ�]��愾��b?��.���![>���>� �>36�>��->�LG>�LU?F�G?���>�x}>cq���ľ��۾�2������\����U����:!0�猚����>�#�E��Y�����<B�K~=|qQ�:��4)�N`�G<D���*?uV>��վ��N�WH;Yƾ����Q;�<�ͽ�Ǿ��-�Ծk�D��?��>?�����fP�O�	�������ɽ�X?N������������=�6K����<	3�>ڤY=ޜ�:1�޺L���/?�K?�{���:��G�$>Z�G7=��-?�\ ?�m�<BG�>�%?W*����rsT>a,3>a]�>���>&>9��N	߽TT?��R?n���ћ����>�����o�z�=A�
>�8�P"��U>H�<+�������� ~���*<	&[?"<>xY*����wX�����<R8=�R?|7�>?O�>��Y?`]T?�:"�0�
��TQ�h�,n�=)|g?P�S?�9>��<������t)?v�b?Jf>�l|���ξ<�!�sD�w�?�Ye?�#!?�����{�HՓ��^���L?LO\?����䗿�v��~:hT�>�i�>�?1�k�h��>�@?B� >	Ǖ�ސƿ�w�q��?d��?I��?���s����=��>�o�>Z������al��ނ����=�ٛ>k�J�J�:��U��$dڽ	?��.?���>�L�6ླ��=�ؕ��Z�?p�?󃪾[Qg<M��l�<o��z��<pͫ=5��H"�s���7�h�ƾ��
�D����ῼ���>!Z@�Q�;*�>E8��5�TϿ���v\о�Tq���?R��>��Ƚ������j�:Pu���G���H�����aW�>�>���X����z�}3:�������>U����>��J�"���N���+�;�ґ>�@�>��>C���~����?�$��^YͿ�̝�A��J�W?9��?���?� ?�7<<@Kq��y�VrV���G?�s?�Y?���\�b�?n8��f?�+c�a]&��//��}q>׋,? r�>�D5�L��<��M>Q?T�C>�~,�W龿�����b�$�?���?�M��?��?��?N�4�����SpϾ���<2#�D?�a=>Lþ��b�I��*��%&?#?����1��i?�RS��oV����O7��#�>�I�=�X6���8>�P�=�Q�F��2Ԁ��x�?�E@R�?������2���?�(�>�F��������$>�k�>�>^5���ۧ>�:��n��9��<?+�?��?;�1?���$��g�>���?:�>FN�?��>�?�@>Ǵ8�&�׼���>>�CW���?f�B?�x�>��6>h�X��,#�iF?�BuA�P��̌2�5��>�eW?��W?�Z>H̦=�E�=ǵ$�|���D	��jq�<#�`�@?�=�VؽG��=a�i=w4>�%�Pz9�a�*?�yc���ʿ�N��=��=##?u̿>�R>b��9�z�=��?��>2���4��i;z��[��q�?A��?\:�>�D��0P���5o>���>���>AnO��-�;���=�V>�?�ϖ������5��f�$>�7�?o��?�ڨ?�p���	?�f辚�}�4@e��� �����=>�Z?��ľRA�>��?G�=x�p��٪�\ag�A��>V��?x,�?�d�>W(g?5���VE*����<n�>x�]?��?�*���gƾ�>�?��������̾�Ie?V@��@��K?*���gݿI܏�Rr��\�侯�;�{t>s�5>�zt�/�=�1�k�!��ܤ����==�p>0��=e�=�=.!>^�|>���]���E��lɦ�zFd�������F^��
��p��V"���ƾ�j��J����'k��.4J��%�<)�;�T�=Ox^?�}S?q�z?���>Y}k����=�Ѹ��>��X�|T4>S\>�B+?�wM?��>�X6��!��ap�vz�Ja~�"3��G#�>�h>덨>�v�>�^�>���P�=R��>�s�>e�C>ωǽr��������'�>B+�>�;�>Xx�>�2<>��>`δ�A1���h�>w��̽ �?”�ӽJ��1��h:������x�=^d.?Us>���C=п0����2H?2����&�,�+���>��0?�aW?�>|����T��;>���`�j�t\>�+ �<�l���)��!Q>\l?n�N>B�p>�z3�oc:���S��m��a�>ϐ4?p~���G� �w�>rI���ھ�V>���>\ڻd��n���j�{�i�`���}=��9?��?T>���<��Vs�J㞾+F>R(\>� =�r�=��[>��E���Ľ\�J���+=���=OdY>R�?�B'>\^=�s�>�ޚ��rF����>�n>�,>1�C?k)?V���[��х��&�7���~>���>�C�>�>��3���[=>�>�P\>�ə�sP[����H��_>����C�����i�<xHu���>�3�=B�̽q5��<��~?U+��ɗ����꾥w���OD?��?���=:/{<�)"�DB��s깾{��?��@�?y����V���?+	�?�R��[��=M}�>Z4�>�;O�L�x\?��ǽ�A���
�$���?	��?��/����Hdl���>�1%?�Ӿ只>)���D ���/���T<�z�Z����>w�?��;� ެ�e~�K�"?�C:?X���t����տ?�d��=�>��?\N�? ㈿�h��N�K�^,?P��?�r?�$=��¾b��=yI�>�;?0�G?D�>Hj4�4o���Y�>���?*��?�H>މ�?�s?.��>�v��`/�l"��e��;��=�c;9)�>��>D���a�E��Ó��R��G�j�$���`>�c%=t��>��佳��L��=Z���~%��i�d� ��>�{q>��I>�3�>
� ?�B�>��>&9=�ӌ��������F?�?H� $Z�+��<�f�u�F#?�U:?��μL�ž<͢>rrY?}��?�*P?�]y>��
S��V
¿�������<Z�>:,�>���>Խ:�D>�<վ�7��>$�>.$�;\ ��|���C谢>9�?*�>1k�=�� ?��#?�j>�(�>aE��9��J�E�f��>��>�H?��~?��?�ӹ�Z3�����桿��[�:N>�x?�U?ʕ>���򃝿�nE�AI�����^��?�tg?�U��?�1�?T�??Z�A?$*f>h���ؾ@�����>$�!?4$�ƱA��@&�f��y?hY?���>���Oս�BӼ��/�����?,%\?�D&?����'a��
þ6��<s�"�
�T�K��;3SE���>H�>�r����=�6>8��=om�86��rj<��=(��>J=�=w7�������&?��:�)���/Q=�Gu� ^<�sj>9�>���[?ʗ�HEp��b��������F��T�?n��?��?@�����h��IH?$O�?��?��>���"��R���GP��>G�D��僘:�b�>�<��aP��Oݛ��룿�~������5�8�?�:�>�N?��>
��>�4�>�=۾|*��Rؾ,�~�x�\V�����&�dB��������ڽ�Jվ]�L�&LU>4��=aغ>5��>
�->.�k>G��>�=�x�>g�A>��>ݔ>\�F>��=5D=�������9U?$/¾�;.�]�ݾ���#C?�Db?&#�>�ء��\����$?͐�?T��?��*>�,f��\ ���?)�$?���;�?�,3<��X:o�Ľ몸��E���`=?w�dՄ>���{=6��8��$��;��>r�?W=
��:�e]ǽ�����o=�L�?o�(? �)�u�Q�
�o�B�W��S����7h��h��i�$�ɖp�ꏿ�^��A$����(��Q*=܉*?��?!���������(k��?�Ikf>[��>� �>�>�tI>�	���1�u^�:L'�����(O�>�Z{?d��>9pJ?�>?]�R?
aK?/I�>=��>JG��)��>��q:ϴ�>���>We9?v�-?d�-?M?d�'?��Y>hi��<��T־��?��? r?X�?��?Kk����ʽ���-�������[�pݑ=4��<T9߽�����3=?�P>p<1?S���>7���Em�>��:?6�>��1>BC��u�-��=�(?�h�>}>>ێ�ԂX���ؾ�?n�?:�85'>�ﴻ5�/>ioV��&�<�B)>��F<�oݻ��νf͎;�ͨ�ji>�%W>K�k�������
c�͓�>�t�>q�?�_�>�Ј>Z��+� �c�����=�uY>d.S>%>��ؾpd��z����g�)z>Mr�?Ct�?�8b=���=���=����6��û�X������<�b?�E#?�T?oi�?:�=?ba#?W�>�$�j[��u��M좾ڕ?!,?⊑>�����ʾ���3���?\[?v<a�׹��;)���¾t�Խ��>N[/��/~����D����p���~����?˿�?�A���6��x辜���\���C?="�>nY�>��>z�)�w�g��%�m1;>���>kR?��>P�O?�h}?��Z?�gQ>C�;�����2���9f<��>�=?��~?�?x|?�O�>���=`�M�n[�\���]߼f[콢a����=��Y>ݷ�>��>6��>�y�=�ѽ�$ƽ��O��l=;b>�h�>��>]B�>c�v>v8c;?�+?0Qz>�`�L�뾜 ������E��!�?i��?Q\E?��=J��:To�Z�:����>ƨ?�D�?2=G?��G���Z>��W�����vd?��?CY�> 0L�tT�5�>`��>�u�>iӽe�۾�����=��?0="?*1&=��ѿ��j������|ξ/��5��GP(��6��j�F�:_?�؛����J�����Q������,��x^���4v�0�+����>.g�=�!�=�m�=d1��@�_�ݺ/<��ٻ�����P=��#�%�;����HF<�b�<ZG�=4G�=���=J3 ��9ǾG�?�(F?kh2?C�@?u=m>=�>�ޅ�2�>��W��?��0>�UL�*㭾�+C�������������7ݾ�j�Nx���>���Ib>�2>O��=��<R��=���=�Z�=��b;Z��=���=�Ի=��=%��=Vw>��>=k�?;f���W��f.<�O)?qL?O!�=ڃ�kk�?b&?��=��װ�{TξBr?B��?�,�?[�>O���S��>�l��m��;�R=�����w>Ff�>M����r�>���>���Uo���#l<]��?���?� B?�ܜ�I`׿��<��?>��=S���1���L�c�a��~[��?=8�N�Ⱦda�>)��=}�0�˾�=��=>J?�=p��?�[�*e�=��o���V=��V=b�>baC>׋�=�M���F�=͹6=�y�=\�Y>��T�-�u0H��<>Ҝ=0�`>��%>���>�?^`0?�Pd?�!�>Mn��#Ͼ� ���&�>�4�=@�>O��=�NB>�t�>�7?!�D?�K?Ow�>cω=9��>r	�>�,�Ȫm��d��Ƨ�7O�<���?�ˆ?��>��Q<*�A���Sd>��Ž{~?\1?�t?��>Hx��=��d�-�48X�p��Ο�>~d�=�qz�ϛ�<�s���B����$N5����>�3�>���>��|>��B>�h�>.��>�'d>��=�9��92m���Ͻ�:�<�=�=��y=���ٽYL��(d=��K>&�>Z�3>��=�X����T��=�2�>c�>�+�> Q�=<	��s�/>m����RM�@�=�3���B�%"d��'}�O�.�>G6�en?>ƀS>�J��>A���?�\T>v	B>�A�?�u?�5>Z����Ӿ������`�w-W��=!�>QNA�T�;���_���M���Ѿ���>7�>d�>��l>�,��?���w=��wc5�u	�>�e��R���J9q�=>����	i��hκP�D?HD����=r%~?]�I?_֏?�y�>@^���^ؾR0>�%���=W�Nq�AÓ���?�'?�>e ��D���˾���ΐ�>�I�r�O�袕���0��� �Ġ��ձ>�c��}�оz3�[p����~SB�p�q���>��O?�Ϯ?��b�D(���2O���Y{���c?
kg?h�>��?;O?1��*�;������=)�n?Q��?�2�?�x	>:A�=7����w�>4�?Ɩ?ϝ�?�:s?�|@�@�>��;*c!>�j���O�=I�
>�+�=���=8?��
?Z&?�"��6j	�� �A/�{9^��s�<V�=��>e߈>��q>���=�`c=�3�=]�\>
T�>�~�>r;d>���>7�>�ؠ�����ad#?B��>~C�>�,?N�>Z����,x���>��|=۵i��2�������z�׻��}ѽ$ܽ��>c�¿ ӽ?�$,=����a�>�ξ�_��C΋<�>Gbݽ?S�>�M=<�M>ս�>��>�>mș>BQn>����|e�=�C	� ��3�e��m������yo�>�zо�rϾ�����2¼n'F�Ǹh����w
���kg�DJ&��qƼs��?���4vE�/�G��]>�Ш>�s�>��?
⭾��Q�b>9>�,?�C�>���Ԑ����L��m?p?�;�?4Q>y�?�S�?�l?&tύ����Dp���_�jb���EK��q���H�������s�i�ec?I�\?�q�>�ɣ=p�K>�|?�����j�>�@��Rd��`�>;�?%�%־@� �Mb���^�u�+��u?�%�?F�C?c��{���@hF>vF@?�H?�!p?��3?/�;?�	M�	�?\Ln>E[?��?,hG?��,?�
�>x�;>ixQ=kr���=Z�7��ϛ��������6J�����=���=_�:�n٧��5w=~[B;W��DDM�)r����e��_q=7}=��=��=	:p>�1{?�z%?S�[>�eN?��8|����0+A?�}�=�����{�v����O׾��]�_�q?�	�?�F?�q���-N�V��|�*>�qj>�>��>ѧ>ߡ$�1^}=�Op>L�|>Z\>d>"�^�C��}�:��ܾ�x*=�'�=���>���>'蒼��P>į�N��M�?u̫���ؾ�eQ��c�V�B��Dl�� ?'�k?�3
?���`�N��#��6bd?G?}�P?�y?���=u'�BA�g��T�\�)��>0e
�������ſ��K�ȗ�=��>Ifž�﮾�HZ>k��m�޾Z�r��?M�L�,�y=Z�
���c=���hCԾ||��L�=�E
>Ӛþ�����X
��"{L?�>=K���+]\�{$��V>>.�>&0�>��T����]W>�ܥ����=j�>&�E>́��K��~�F�[��vƄ>�}E?�X`?�*�?nς���s���B�� �����[����?:ĭ>Տ?O�;>y$�=J�����.%d���E����>�X�>X��ٗI��5��o���%��
�>�#?�Z>��?��R?�p?��a?�E(?��?	H�>ӕ������5&?z��?�ʅ=T�Խ�OT�+	9�v6F�Nx�>̥)?�C��g�>W�?��?�&?i{Q?��?�>�� �bf@��i�>zH�>T�W��A��`>w�J?N��>�
Y?�ȃ?{�=>��5�h������V�=��>C�2?w+#?j�?�=�>���>�����I=�ܲ>زe?兂?�/j?J �=�#? L!>4��>�=ܞ>_��>f�?�;J?��o?PN?/�>�A�<�豽p�Ƚj�K����:sA�;to�Ov=�)¼��K��5F��8S<�"�<n�v�)���/��e����j��գ<�>�H>ϻ��d�>iX����!�H\>~<A���)�ɾPr���>o>���>�eR>���3>��>h^�>��h4?�?�??i&����G�bx��E�<�ߖ>�E?��=?�V��c��#�n�M�R>!t?��o?�Q����1�.�N?^�]?��\�����n����۾
��h��?CT$?�؈��l�>�׃?��?x��>�U:��b������{q�~���P��=�8~>��>���w����>�:?�}�>`��>�^'>Tq��*]����̾��?}��?n��?^��?@�?>��y�/-�� �����&d?��>��_� ?><9a�ꋾbӖ�'g߾���������y�o��bq�����N�$�1�~=g#?	Wm?�fo?�V?�����f���k���w��T��|�����D�QJJ��L���b�����¾��R��o�="�6�3�?j�?��-?x�'�N�>�r���� ��zɾ<=>�(��_a!��4�=+4Y��mo=�)<=�Sr��nO�ϡ��n#?&��>s��>�?8?[RW�!`@�5�E6����V�>��>4�>���>��(�-�&ώ����Lc�H0u�v>%zc?@�K?�n?�0��21�Ї���w!�B".��d��eqB>ʞ>v�>�W�t[�h2&�zj>���r�i �yt��}�	��}=��2?$%�>g��>9F�?��?�`	��?��nx�Fz1� ׀<?�>)i?.5�>���>�нK� �%��>*�l?9��>��>�����Z!���{���ʽd&�>_�>˳�>��o>ǫ,�a#\�	k��烎�m9�Ku�='�h?���z�`��߅>�R?N��:��G<u~�>��v���!����|�'���>6|?ؒ�=!�;>l�ž�%��{��6���Q)?�E?�����*�k1~>�!"?�z�>�-�>�2�?�"�>�vþnmE��?��^?�AJ?vPA?5�>��=�걽�HȽI�&�V�,=ȑ�>�Z>��l=���=��3�\������D=��=oμs%��a�<�=��{�K<m��<��3>�ܿ�K��X۾��P��ZP��S��d���#�������^Ǚ��w�\��3�&��X��b��Ќ�[2n��)�?���?Az��	���ڙ����u����ȼ>��q�\�|������	�Eo����޾\0���@!�EP�$�h�<Re��� ?�����#����$�>ְ6?J�j?�d�=5E��+#�9��>�� >An=�¾Q8����ʿ�"N���o?5W?D��Ҷ7��u�>���>�>�>��=4�Ⱦ�U |>K�?'L?���>�课d�ӿC���ځ�=���?9�@��>?)l+�]�����=u{�>��?�P*>��q�P%���A�>/3�?�2�?_c<8�W�E����xe?�v�=�8��3�B�>�X�=o�[=�s-�)�s>��>���/#Z�U��B'>D�>����p�B�X�U��=�_>�����潙�??C:�>>�f��SF����O>D�a?h�><��>��0?2tQ��2ɿߝC�Vs�?#�@�m�?W��>$��d�z>�p׾GgO?��8?\��>Y��a�S���&>��. ����ʁ\���*>q#?��>G������~=�*w<�w>���ƿ��$�P|�>M=�6��Z[��;�}�� �T�����bo�ǅ�Y�h=��=wlQ>�h�>ZW>�Z>gW?��k?�K�>r>佝����ξ����G��+���������裾WE�Ԗ߾�	����E��$�ɾ�f��W};M�Z�����A�r���z\+�H�8?Z:G>d�о�1�Q_�<��!<f��d�<"Y#�0�̾� -���k��?p�?:�c�Gm��i���b`���N��}D?Y�V�nd����uQ>��=�i�=���>�PW=��,��}<��e,?&?�����΄�l��=kz���q�<Ft1?"��>�<\=4��>`9 ?P=����$�D�Y>ŦH>�޿>y7�>غ�=�]��I꽌�?�fG?�8�)���dp>� ��.�h�
.>��+>?�P�a��E�v>���=�^\�'";�F �;�G���L?7->�#�'��5B�8��;:��=EO?���>{b:>>o?;�C?F��b�NU�xi���>��_?R?�F>���|���W��ݿR?]s?E�>nZ�����/0����u�?i�}?�$)?����n�o�E����̾ �?�B?��S��������	��d>9?�>�4?RNk��l�>?�'?�o>�C��|��""G�1�?�f�?N�?5K�=/���C�>aP�>
)�>LQ������/>?䇾П�o�>�� ��%	!������/?��U?&�>�ʬ�W��^��=�Օ��Z�?��?σ���Xg<J���l��n���M�<�ɫ=%�=S"������7���ƾɻ
�����aߥ�>�Y@�R轝)�>�C8��5⿜TϿ���y]о0\q��?~�>��Ƚ������j��Nu�}�G���H�w����k�>��>�ꖽw���>|��N;�Zq�����>Ј�I��>t�P�mδ���� <VI�>*��>���>�����b���s�?�6���XͿ���!��P�W?�*�?�5�?��?vw<b/n�r�~���b��G?[t?q�Y?��,��kf���1��j?����	I`�TG4��jD���U>t�2?���>�Y-��r=Lk>	��>��>9/��KĿ=���,����̦?Lg�?�L�)��>pI�?�V+?d��м��_Щ���)��rS�-�@?�1>]1��;*"��I=�Gđ�+?c�0?h�������k?\�?���C���X/w��>��g"�4�4>b&>\!V�E��Ү��N��?rb@��?v$����C�}��>|�>�q�Cm��Ik=H?g>{��>�ɇ>�2n�¿�>0s/��k|��=��?Vn�?��?��z�%H��>>2y�?�¶>��?0��=���>�)�=�E���ۂ�q(>�� >�L?�4�?բM?Z��>E��=��4�p�.���F�&�R�y	��(C�N!�><�a?lLL?��`>_뼽W�(�qo!���̽�c.�w�\�>�Lo?�Zyٽ�6>:;>��>+�A���Ѿ%?�h`���ʿ������=
\(?$�>0��>���Y����`>۞F?OZ�>�	�����!Î��6*��B�?���?o��>����˻��>�נ>�?5�_�Uy�����ҬF>�~$?}���~�8�s�z//>;m�?���?��?/�=�k�?�D��\���E}�.��)'��<�=>7?�c�Nw>��>U=�=�uu��u��hs�	��>YƯ?o^�?Z��>Zoj?��j�ې?���I=/��>{m?|?N �;�����&D>r�?��
��Ȏ��>�mRd?Ɖ
@�g@�_?���}��yՇ�"6⾷�����`�g�n=�>��T=��>7�����'(�W�J>jo�>�i%>�t>_c=>�C>�=�����]տEm���ń��I��T;��?���ǾC��#��ˮ�t�W��ٽS�z��-�%�(�ɔ �����u?>K?���?�8�>��=H�d>�r!��93��Iּ\#>x���v?�dg?\K&?kN�=���a ��\������a���� ?;l>�=�>}p�>��>��c�>⊾=�:>�$�>"����>��D�<d9 >�ȓ>^[i>���>�D9>��>����yL��k�h�J�y��ƽ��?�e���MK���x���d����=�e.?0'>�����Ͽ�����H?�w����V�/��	>�(1?U�W?"�>^ױ��]�+�>����
i����=����	�m�8�)�UAR>��?D�f>�'u>��3�K_8���P��~��%Z|>B46?�ն��A9�5�u�=�H�
WݾF[M>8̾>�C��n�������rvi���{=kx:?��?�;���尾Ԧu��J���DR>95\>�M=�o�=�AM>�:c�ùƽ;H�Ɣ.=���=��^>Z��>��>d=���>���{@E����>��m>*(�=f�6?GY#?
X<�F��C��?8,�H��>%��>3=�>���=�6���=n��>|u>>}�!�؁�$X��SV���l>�ۼJ���u��(�*;7���@>�ϒ=����v���U<<�~?^i��|ψ����b���kD?WD?u1�=�	V<7{"���k��"��?j�@�|�?PQ	��V��?�5�?&���Ջ�=|��>��>�ξ/�L��?��ƽ�'��I�	��#��Q�?��?#�/�Pċ��!l���>"X%?��Ӿ%\�>G���c��~��y�t�ZH=���>
�G?�'���`]�i�=���
?�{?���@��TGɿڳv��5�>���?�˔?:@m�b���O>����>e�?��W?��d>�Iھ�R�Q��>�|??�rQ?��>N��q1(���?.��?Ņ?~G>r��?M�s?��>)Tu�x�/�����Ɍ�n}=��z;��>�>{�����F����y����j�˵��`>~�$=��>F�4�����=
ƍ�f˧��7j�
��>�r>�K>�>�� ?��>���>H�=�[��i����K��6�6?�?�����,G��k�=a�˽qѾ>L7?_�Y?Dｽ��T�>��}?|�p? VR?�r>8�7�x��[9ƿ,0���it=�~">'�?�9�>Ɇ���\i>�� �]1�aw�>hFA>V{�}*��4���=��x>_�?�^�>G�<��?�&+?p�>�/?Sy6��l����T��޽>��?�?�с?Or-?����0&��������x�~�Q��=�l?�-3?KU>n߁����'S�n6dM���?>�A?��w�}W�>E�?k�j?3l?�[>��#�M��@-w�W<�>�9"?j����@�΋%�uy�G�?�Y?���>쒑��+ýCW���1�De����?�]?A'?x���ba�hyľ��<��*��f�F��;(M`�9a>r�>�Љ�m��=g�>(Ϣ=��o�m0�ܞ�<k��= ��>���=��;�xe��,H+?�ll�5���=�5s��B�[�>�yN>��ľ~(^?k�7��0y�{3������QKX�$��?�i�?L�?�창��g�6�<?Ɓ�?%-?���>%3��hݾg���er� T|�Y��+��=�G�>�d�����᩿c���漽�	M��0?�C�>��?l��>�k>z6�>iľ��8���ܾ���v�o�T0�_���$����1����W����$�Ѿ�]O��މ>������>g??q~}>�iq>��>���<ܥ�>��U>dl>���>�N>d4�=��@=&���KR?{�����'�Jj较Я��B?2d?�w�>ſj�'���|�/z?mI�?��?��t>^Jh��*�f?���>�>��ǵ
?�==��UWi<�׶�0����M��A1�>��ֽ6�9�O[M�Чg��
?]?<{s�]˾$2۽U�оʾK>pS�?&�c?�����f�k�W��J��~�'��N�=��-%��1�E�x�Kz��ꍿ����D��н�H$?L�@?�NȾ��ҾE��Z���.��:�>��?���>�?��>��¾����gl��%����8�>��?��>L�I?�<?LyP?�jL?~��>�b�>17��\f�>�3�;o �>j��>��9?9�-?�70?z?s+?=+c>z������ނؾ�	?�?�J?�?خ?"݅��rýwU���wf��y�
�����=N�<�׽�Zu���T=<T>[.<?��ӾXm/����G�&?��!?{�>�Y�����G��R�7>���>uS?(^���]�&���}��'?}]�?�s�7C	>����!b�>Mܠ�I�<H��=��ϼϝ����ҩ��ɿ��`�;Q
�=-4�=�N|��`����Խn��=!W�>��?���>^	�>����� �k���"�=�Y>xX>��>�Fھ{ԉ�������h��y>̺�?|��?,Z=�|�=�D�=�����Һ�Z~��Q���`=B�??J ?VR?�5�?�e??��"?p� >���_������9M���>?}!,?��>����ʾ�񨿴�3��?a[?I<a�&���;)���¾��Խ��>�[/�2/~����ID��녻����~��/��?쿝?�A�T�6��x�ڿ��2\��F�C?�!�>BY�>��>F�)�v�g��%� 2;>���>VR?��>%�O?K;{?M�[?�{T>��8�H1��>���"f-���!>@?���?���?-y?e}�>��>*�7��w�������~ۂ�nzW=h�Y>C��>�&�>˩>��=�ǽ�o����>�fդ=|�b>���>ޖ�>\�>$�w>���<��G?�f�>RK���j�y������L=��xu?�K�?h�+?f�=��WF�[���>�>�B�?(�?�**?�[T�&��=��ݼ􍶾;�q���>�|�>!�>L�=lEG=�>,}�>���> E�c����7��I��?�5E?���=�>׿�i��L��]���?V�Jʾ�����=��]��={�m�h��4�����.S��s���ѩ�3���4���D?��'�΂�=�'�=Ow=eL��H���=!�_�D�~=@�p�Au�=<�7�L�$=��<]B�l���?E8�4�.�˾��}?9;I?>�+?s�C?��y>:>7�4�Ay�>`���>?��U>֞P��q���g;�c���2.����ؾ~�׾�d��ʟ�R>� I���>953>��=I��<�Z�=us=Z	�=��B�)=T�=p.�=�D�=��=��>U:>�+v?�kK�1�s�?��~֔�ͮ?�I�>Rd�=d�����?��>1�g�5Ͽ~sϾ�?.�?�<�?�d�>����P��>����~S=��="^Ż�f>���>�����N�>�n�>�������m��=bX�?��?��G?_���Lۿ���=lM+>'/=��G�^1,�� ���0d�,���,?3�@��ھ%~�>P->R�
�6���C����e>gZ>q��;��*�9>���lM�=�I�����>�n%>�"�=��X��MU>� ���|>���=�� >O�K�R����I�0J�<�ON>E(�=�{�>��?$`0?kRd?��>�m�|Ͼ�8��!0�>���=,&�>���=�B>~z�>��7?��D?��K?�u�>7��=���>B�>~�,�r�m��u得ާ�1m�<��?+Æ?NԸ>IkP<��A�6���c>�\�Ľ�z?�\1?�p?�Þ>�U����?Y&���.�Ɖ�� 7��+=mr�(QU����8m�6�㽧�=�p�>���>��>2Ty>�9>��N>~�>��>@6�<mp�= ጻ���<��~��= ���k�<vżz���mx&���+�T���	�;��;1�]<{��;!]�=8��>��>���>�#�=�O���7.>�5��$O�nԾ=�1��].E�k�b�^/z���,��|1�= ?>�bN>�S���/���?j�T>�UB>��?�t?�>�5
�0%վ|�����R�hX�$�=Q�>aEE���;�4�`���L�k�Ѿ���>�ގ>��>��l>�,�j"?���w=��b5���>�{��˸��(�y9q��?������hi�ɢѺ/�D?WF����="~?��I?H�?u��>�����ؾ�:0>�H��*�=,��.q��n����?b'?���>l��D��G̾���1޷>l@I���O�\���0���ͷ�#��>g���(�о3$3��g������ˍB��Kr����>:�O?I�?~8b�yW���TO���2'���q?�|g?��>�J?�@?&&���z��r��]x�=�n?���?7=�?�>���=�P���V�>َ?���?1��?޽r?��@�Ƒ�>�:�">h����=Y�>���=�'�=PU?�G?g�
?H����`	�.2�L��z�Y�8�=�J�=�ȑ>���>��r>�b�=�c=2��=`�]>|a�>�T�>~y`>�>�d�>yʬ�wb�pG(?�>�>�>S3?��>���<������<&6�-�K���)� ˊ���ͽt�<ϯ=���<�aX���>G�ſ���?�A>�u��U?����սB�O=a>�C4>ss�)��>�_6>��f>��>��>��+>܋�>-�<>r���$���gK���M��Ol��'�p��>6��#pξ�����ՓS�ð:��?��~�n��s���6�M��V��?���͕H�k.V���=ݦ'?�d�>��?��ľ�uH���W=l?Ŝ>�7�#Y|� #��I���E�?��?��+<��?NBy?��>?������N��5a�%Px�ϡE��=}�F6o�l����~�3T���8ݻ��^?ȹ{?���>X_��\�h>:�f?$���Sꗾx�>�4>����]�x>��>��'�^7�t�����jB��X�e��?2/�?�R?P�kfj���&>�w:?�p1?LSt?�1?�i;??��s�$?�s3>y;?	s?AS5?�.?��
?�{1>���=����\_,=�G��@̊�@�ѽ��ɽ�$�C2=F�|=,w��Kv�;ȁ=�3�<ķ���ڼ~)(;������<v�9=�С=���=R�=�o�?w�X?T�>��W?:7����������8?�uk>#FT��+��[��Օ����h�߁?&@�?I�"?�Pp���(�Z�V���,=1��=#Ǯ=.ES>�ћ>��a��b#>��Q>��>�Y>�������1H�;����x=��>Р�>޷�>|
�='��>�޾��Ƚ���>��;"I¾P�y��H_�LL����l1?�}?o"?ȊO���t�}K���h?�y?u?a�v?3j�=B����a�w
��.νj�?������
��3�������D����=&�>[mǾn��t	+>J(-�� о���mUX�������>JN��ʄ������(����c���@>�>`;����4ۈ��f���J?�͒=�7&����C\��Wz��vw>�J�>f��<Ga����4�X�¾�Q0>��>q.>	����)�L�:��f�>>$�o?��?x��?۰=�^��zp�ݷ��8���þ�-�>���>c�:?NM�>���~�N:2�ӎ���>����>z=>Y'7�1�4��?�O�0���辳��>��?�]�>8�
?a{/?���>�2.?2�>��>5�I>2��[��A&?3��?4�=��Խ>�T�� 9�ZF����>u�)?/�B�ӹ�>W�?�?��&?ЅQ?��?��>�� ��C@����>DY�>��W�qb��C�_>��J?�>N=Y?�ԃ?_�=>I�5��颾>ש��U�=>��2?�5#?5�?ȯ�>��
?�ľ!�<���><�y?�}?��Y?/=>�"�>b��>t�?��G>q�=���=��>��E?~!�?�yb?M�>��:�t��2����ڝ���/=; �=ӹ/�o<��=�Я���m(>��>)D�\#?�^$�z`��}�`>����5�>�#u>qQz�֯>����=����=�(,>�6���b�� ���9D>3�t>���>h�.>G%<�Px�=i8�>/��>����T?N2?��?�H/��[�����<=�U�>q�a?��=R\h�Hr��|�n��>>�z?R�[?�tν`�*�l�b?�^?k �[�<��dľ�f���T�O?��
? �G��F�>t�~?%+r?���>�qg��dn���ӎb��n�ߗ�=>�>S+�ڌd��ޝ>�7?֓�>@tb>*e�=�b۾�uw�4ݟ�k�?�?��?���?�")>Fn��2�T�{	���&a?fH�>�y����(?���<;�:|���ܤ��������⢾�0��Iq��Щ�_���J�����=3�?�Wr?��?��O? ���i�D�d�V�o�/V����h���G���B�g�?���l����*]ľ�UT�\>�(~�)�>�H;�?/�(?��+��>�Ö�N�����Ͼ��;>"���W��4�=ѐ���~G=]kV=��k�ج1��q���$?��>��>�;?�l[���>���1��7��S��|*(>g��>���>�F�>u�z���0�/��ƾ���Eb½=�]> 3o?Z	a?8l?� 9�>BW�5��z�3������Q!}>KiL>J�>>��S��R5��IS�����1�<�*�k����|��=�I%?bn>歝>ʒ�?֕�>������w�pP�����<��>�]m?���>��!>��Ľ�8'�M��>+��?�?P'�>��O��u"����y;���>+8V>�R�>�1�=�(���L�6��9�hS4��zm=:O?�b����`����>w(<?1�6<�����>48���&��ؾw�[=V%�>�� ?�>]#>����7�[r���f�0U)?u/?ݒ�x�*��~>p""?��>�_�>w5�?E,�>�Mþ�&���d?��^?WdJ?�^A?A2�>!=,���Ƚ��&���.=§�>�[>��m=���=�9��\��T�I�D=;;�=�ͼ_e����<#߷�6�H<���<^84>�ԿZ�D��ﾦ��ڼ�w���V��Cj����_�ȕX��8��@Ɋ�ʝ��X��� �G6���5��@y���0�I��?��?�5�:3��H��H�[��⃾��>���'�"����=�����;��뤾�9<�a�@���<���V��'?춑�#�ǿ>���F�ܾ��?!J ?G�y?)����"���8�X� >%g�<�i��|뾟�����ο?�����^?���>5���[[�>�%�>�[Y>�q>�8��L��oV�<*�?.~-?3��>7�r�ƗɿX����Ǡ<��?��@͚A?|�(���|HN=���>�	
?��=>uT.��A�U��N/�>��?�)�?Cg+=��W�?S	�N�e?|�<�E�������=��=��=����H>���>����<�NܽC�1>���>��������^��<E.X>(�ɽ8ߗ�[@x?��W��os�aN0�i:q��\�=ܚ+?b��>��ͽ�P,?}\��HϿ�z��6{"?>?�?�?�?�l:?Øv��L>��վ;e?^�.?<�P>���E4���;P�=��'�5�ܾLI/���s=��>Z>u2��Zc�kk>��D�<���=���kƿ�>$��g����<U��� h��1�_ᬽ�Z�J���Sp�c���p=��=K�S>�[�>��T>��\>��W?..k?eǹ>��>#I��e��7T;�����#��Ne�	���X��(���"뾾�޾�]	�d��Ӽ�>`ɾ�"8�Q��<�f�v8���}I���W�P""�?p7?��5>nZ���B���=�*���{~��Y�-P�e��l6 �G|V�� �?~H9?�
����9��R&�ƪ�q�=o�i?���c'뾪�ʾ��H>���q f=?��>����Ѿ"�%���C��]0?U?/[��N���&>N:�
i�<�/?�� ?]��<���>�}$?�2�D����W>�75>D�>���>h�>�ѭ�����?��R?p��	���ɍ>0m��D�r��Ȏ=�>x�7����`	V>���<>��ͻ����ȱW<��U?r��=���� �|"���=\���O?9u+?�>�Y?\�W?��<��*���_�u����=���?��X?�l�=��=�Y��ҾK�?�L?;�>w����,���2��������>�q?�(?K��Z��b@�������d?,o?��r��m���B�T?=u�>m�%?$��>�o��?-�1?�v<Jb��5�¿���z�?L�@���?�,,=��<kZ�<>ڙ>%�?����oľ�2�y6<��j׼;�>؆,�ޱ_�]�3�O��=��??�|{?<	�>��־�����=�����Z�?��?�y��JPh<����#l��{���>�<Ԋ�=�}�v4"������7�0�ƾ��
������㿼Ο�>/W@��罍�>X8��2�LPϿ���nbо�kq���?�t�>j�Ƚՙ�� �j�sFu�ϩG�4�H�'���v��>�><�ɽ!ה�����@5���K��L�>��ڼ�}�>�KF��\���垾:�<D�>Zg�>Q��>Q��������?4���ο������	��W?�>�?I�?��?�R,;M�n�dd��QҼ�D?v�p?�vQ?g7��Yc�ӯ���h?�A���V�.���1�ȁ�>6�&?�%�>Ф"�Ϋ=@�4>�r?�\)>Й/��^¿ͱ����v��?aR�?yk�m
?�ݝ?��&?�*��w������5��7��72C?,�;>�i���x(���=���U��>?pf.?�i���%/�{�b?��:��V4�5�M8ͽ��>���=���1zt>nB�=��n��ꟿ�Fӽ1u�?��@�د?�����L�U�>\��>�^;�ʜ��?�=^�%>�1�>�ܘ>�I&��R�>i\)����l?�>l	�?ӓ�?]�>�;��}\���)���Y?罪>��?#n�>�� ?�(=�$��7Z��T@>��s>X:�����>�B[?�?�c3>*����8�d��Vd�K�X�>@'��[�>N7G?kr`?�JO>7	�����' ��/�^�ؽl=���,T��;����>П0>M
>�uo�(7S�
;?�A,�@�˿�C��d޽�N+?���>�G�>l
��� �2��Y�p?SO�>:�'��&��1Q��@�ƽ���?lx�?Ah?��ؾϵ �:t�=Ơ�>X�>6:ֽ��[�A�r�lƤ>b�1?�4�ĥ���@��WX�>���?�^@��?�р��?#
��&z�1������X���kE>��.?�ξ<۲>�\�>7a1>�l�U豿�,i�AC�>�ë?� �?�A�>9T?V�b��Z.��(�=�@�>Izf?>y�>�rF��\����>t�?t�"�%֟�-����{?��@J�@0�I?l৿#�ۿxT��RP��nwԾ��=Lj@�A�>R�ٽQ�>q͒= �;=#h��i(>L޴>�]>}�>>��&>E>�z�>�U��3�(��ӧ�L���K3.��	$�\���!�������
�ӵ��(E��l�&���<�<Y����CAW�~Lk=��j=�
a?&�:?ٟ�?xm?V_C>�%l>��3�@�{�ⲡ�XA^=�W�=�3?�H@?4�%?��K߾�ee���z�t���ƾuJ?��s=I��>լ>�n�>��ҽ�&T>�b�����=S�]>9�<���H<�=�ʌ>ܴ>1�>���>u�;>��>�д��װ�;�i�=�y��*ȽvK�?*ƛ�N�J�$�� -�������
�=�1.?i��=Gӑ��Ͽ*����/H?*��T'�Β-���	>�0?`-W?�m>�����[�H>�<	�H�f�!��=}�,n�ǯ)��9O>i�?�^>�%e>��;��2���f���ľ�Q�>�sC?[Ι��>B���w�1�9���վPd>qӾ>P�Wn�����?y��QK����=@A?8�?O���=��D~�
����\>�;H>��=�C5=�r>�톽�����b��E�<΍=r�I>q�?M1>*��=Dܕ>������$����>�]�>�7>MXG?^�$?ۮ�9=5ͽ�գ�9�KV{>���>k^�>}д=tH�O*G=�b�>U�V>��	��o��!�S4��1j>~�����[��C����=~J����
>���='ƽ�w#����;��}?�}���ҁ��O޾N�ٽI?�?{=}Ƶ=�������e��J�?r�@��?�  �E�^��J?�'�?>g����>�(�>Gٱ>~uھ��F�a:?;��h�����?�Ks�?���?��oЉ�:yo�I�	>5�"?��ž���>y�r�����=���+q�R��G�?,�W?�2����h��Dq��$?�!?�mʾK-��6cտ�p���>Ti�?m�?`���+n� ы�oX?h��?�%h?��D�����<���>��G?�{4?��=m�O���!�av
?�T�?��?m��=�Ӛ?�_�?0�?j�q;�5A�`���d����=Lg��X�>58>Kg�_�`��������w���.���>(x/=�V>����(ؿ��S�=���b����a=���>x�=Ck�=���>Gh�>�3�>v�W>�^�~��l졾K�Z���K?��?ֵ�Tn����<��=�]��?J4?]L_��Jоn��>��\?��?&*[?�o�>Z��E��>ҿ�ܩ��Xz�<��K>�e�>5��>����J>�1վ
iE��>���>�5���.ھf!���类�ڜ>�d!?���>���=:� ?�#?�j>�0�>�XE�S<��F�E�d��>���>e5?.�~?J�?����Q3����硿{�[���M>N�x?�V?'��>!�������%H��nJ�wܒ����?�pg?��j
?�.�?��??6�A?>f>6��Gؾ2���G̀>i�!?՚��B��X&����A?ۡ?�F�>eۖ�B�ѽ�ü,�������?��\?��&?����_��¾t�<�*޻�e���<
�*���>�7>�������=h�>_F�=�j��^6��et<í�=�m�>��=��5�玌��7,?��b�����Q�=X�r���C�F�~>[�N>;���Lc^?m�;�I<|�*M���@��gyP�x�?n��?[2�?lc��� h���=?��?��?���>�V��Km޾��޾Iu���y����8�>���>/�g��8�eA��T���׃���Ľ�&�<�#?vO�>�1?6�?Z�z><�9>{ܾ�KE� 
̾�{��w�w*���P�$��0��C���Z]�8׽QǾ������>�`��ȸ> %?R�|>j�a>�Q�>W�<}��>..�>ː>#-�>�*>m0=]�9=�\�<A�.���J?,ݿ���1���羝}޾��5?�zh?��?���Ճ���	��'?��?�H�?Ko>U�k���$�?�U�>J�Z�ԋ
?0	�=0�=8v���2׾�(�JFD�7Y�M{�>�d�R�9�"D�I�Z�0�
?S?�m]�*�Ӿf��h���j�=᳅?6)?��(��Q�-5p�F�V�iIR��56��$i�.���&#�Oo�����i���!��g)�b5*=��*?Us�?��i
�pמּ�k�e?��Ki>i��>g��>���>�iJ>�s	�:C1�=�]��'�iv��N-�>8z?���>f�I?�<?�{P?BjL?Ȏ>�f�>�E���V�>��;���>���>�9?=�-?�70?v?)l+?nc>w�������z�ؾ$?G�?E?�?��?0ㅾFqý����<�h�;�y�恁���=k��<	�׽�u��	U=T>z�+?;R*��~$�~��?�&@?=�X>�ov>|½�^|�֝�=2C?f�?/��<H�F�Мw�~��;k?���?}�V�8R7>S,>�mR>)�R�M=G�&>��=d�]��}ǽ!�<,��"��=�,>^*N<s�	=�O�=�nȽ%CO=��?�?A��>! |>��@���羵�����=E�>��h>�i$>깾~ZP���~e�?r>*=�?~��?^�=wv�=vp�=�L��[`Ⱦ���G��Ғ���>v�"?�F?�!�?V9?;0&?V�>�1�=풿�Q��io��-�?,?�Y�>"���ʾ�����3�
�?�?��`�V�xX)��	¾��ԽG_>� /��A~��诿�D��������ᘽ��?���?�%@��6��s�ڎ��>��aC?%��>p�>�M�>��)��g��9�)�:>��>��Q?���>�U?�?ߋc?� >��Q�&ҫ�J���t=�|>�r??�݁?��?�s?��>�m�=Z!r�=������?��`�}�o�
5�=!R<>/�>���>sښ>>��=Q�M�K���j3�%��=� Y>6��>��>ӑ�>�n>��<�ID?�f>�Vɾ#� � ���G��.�H�	��?M�^?��??��>�����O<��c�>�L�?�?��.?�,3���'>=�`��� ������?$��>\��>$�Y���=�<e>��>i�>2�U<e���30����;�?��?�%>�ƿsq��q�o���<<�j���Ie�%ܖ�L9Z��=Wr��u��)�����V�����ԣ��.����ț�[Ax�^��>>Ҋ=���=K��=3��<�Լ ��<z�S=�Ñ<��<Oh�Ph<04���λь�_W���w<C	K=д��D�ɾ�-�?0EG?Q�2?�$B?{̅>j!>�+���zs>�A��?��/>^�2��뱾d�@����Hࡾ��ؾ�d�PQ���>cЄ��p>v|H>8�>A��<�~ >��e=��=r��<��6=Y��=n��=���=��=�&>�Q>��m?��b��E��ޮ��l0=}>?��>�#>�Y���,E?��?)�p�C������)�m?-�?ޑ�?xY�>�6[���Y>��В8�d��=�2�,��<CJ>>�%��ej>��=�w��� =�-�?��?��/?����5ǿ��=�5U>p�=x�S��W1�f�\�W�N���f��O/?�2��὾.��>�ٻ<�M
�Yu˾aD�=wKq>�>>ֽ�R��У=����}��=Z��=���>�|N>��=$̓�c�3>*�Y=�>� �>�%��\DD�p�Ș�<H(�=�Q>b#>`��>~�?�b0?Sd?�!�>J�m��/ϾG ��-�>��=N1�>���=QXB>�s�>��7?�D?��K?���>%��=���>B�>>�,��m��_�oѧ��ʪ<Y��?bʆ?<�>�Q<g�A���Rc>�ŽF{?V1?ci?�Ş>/	��˳�T����n�w�+i�e�F;ܾ�d �֞�=�Th���ս+�x>��>�>+=�>���=^&�=���>�K�>@�&>�<I�d=��s����=$eμ8p�=^;g��K��`�{���r�Q;��x��R�)n�=��_=e������ʚ�=�!�><�>���>�Ԗ=�����.>9ۖ�[�L� 9�=�g���;B�d��7~�g/��L6���B>iX>a����.��[�?��Y>�V?>�v�?�0u?��>�6�~�վ�=��6Qd�(�R�G}�=
�>j/=��;��j`���M�	VҾ��>Zގ>'�>�l>�,�E?���w=���K^5�{
�>#r��c���9q�?��%����i��Lƺ��D?E����=I#~?}�I?�ڏ?��>$B���jؾ�00>Q8��^�=e��Aq������?�'?���>'
��D�zE̾����۷>�AI��O�����2�0�ː�7˷�Ԑ�>{�����оk#3�.g������b�B��Gr����>S�O?��?i<b�[W���RO�����'��#q?�|g?��>�L?�>?�+���}�0r���=G�n?ٲ�?�;�?��
>�u�=�GĽ���>z?�2�?@J�?\�o?Er:�L��>yڋ</�(>:�x��T�=�0�=Zn�=�'�=�?�?�^?�ס�~�����!��b�\�=��<f{=���>���>Ҽj>Q��="�y=	��=.U>�՗>���>�R>��>���>񦥾�
�K�&?��=n��>�]3?���>n�&=U�����<��N���A�j�)������.ԽI��<o�OP8=k�����>S�ƿV×?��O>i��?�A�ѓF�[�Q>�EG>���v�>�C>�!y>F|�>/#�> �>���>�^,>�6ȾA��=a%�L���Ss�HrS�l����V�>[=D�����0��D���N�����w��vr�H2����9�Γ?��*��Y�6�8��s���?���>Pb+?�M���Q �	��=�?��>~G���đ�U�����r}?�I�?p�>p� ?�Ly?R�C? X�D�ѽ�G�$腿��������^��~&���S��l���nu�9�P?55F?��?"�=0�>8�?��澟�x��G`>-X��#b�
J�>;��>J���v�����#ז�EEI���G�[�c?���?BM?J>�ĳm�X#'>�:?��1?�Ot?��1?\�;?N����$?Xq3>ZF?mp?�M5?��.?J�
?^2>��=]s��e�'=5������ѽ��ʽ�����3=�q{=��޸!<�|=��<	}�ޟټe�;}���k9�<:=I�=�=Nx�>�Jt?X?4��>��2?	�>��S��4���Q?������ξ!jԾq'��jX�� =w�c?��?/L?|�&>��W���H�QL>ϯk>bEM>]�<>�M�>k�ٽ�;��PN�=�pO>v[W>m�.>�_ý6���T(��R��W~9=�{*>�N�>���>;\�=Y��>��M�&� ��>h:߾�Ծ���U��.U-�z���b:?+�d?��>�z���2,��}i��Յ��Z?-P�>� z?e�z?7�ߥ9���I�t���҅_�(��><��x�/�*��Y�����@��_I>J��>�ԡ����v�4>_��'�̾�����~��*޾�I'>"�8���>�'��T���m��m�'>X7z>��߾' �Yږ�J`��oE[?r�ƺ#軾Jz���`��I�->�ј>���>��m;�aսX�3�מ޾Y�#<�Y�>�,V>����ͭ�cv�	l��<>�:T?�bv?���?�;���g�M�]��¾��?4�jb?�7�>�?gY�=-`�>HK������J�T9H��^�>V�>bY/��oH��������_��%�>��>��~=a��>SZ?z?�7B?Vo(?Iv�>���>��������?��?F�D>���6}��S7�@we��(?cR??��(�(m7>�7*?(�?��>��f?�)?A~T>�����4����>��c>(#� @ƿ e#>�u>?�U�>.\?[6�?�>>\�>��)�����,;�<�.=�l,?@;=?��<?~��>��?K�������ea>�S?&gk?i�O?��=Q��>�٦>��#?u>=c�%>�3?�(�>�1M?���?��!?��>^�!=�J=L �<[3=|t��c�-=��<	$4>�½p%�<=ල�>)j���o >����x=	���D
o=�%�>��p>���LE.>�ƾ)E����A>�������r���*<�k��=u�~>�?��>��"����=1�>#�>����)?�+?�?^nP���b��(۾�I���>�hB?Yw�=!0l�چ��{#u��pk=*Pm?:^?|�X�����N�b?��]?<h��=��þ{�b����e�O??�
?0�G���>��~?b�q?T��>��e�(:n�)��Db���j�&Ѷ=Wr�>KX�Q�d��?�>o�7?�N�>�b>2%�=nu۾�w��q��e?��?�?���?�**>��n�X4࿡���6P��ka?���><���0?=��5˾����K��'�־�#��Y������ˮ�{ ���������4%�=�1?�r?Nz?F]?�V�1�`���f�z%x��6O���<B	�x�C�O�I���@�Hve�y9�Q��݋��s�;ӵ��om*���?{E4?�&ݽ�?㚾Q8�9�$�=Ǒ��׽��,>�+?�,D�ypS=0c|���ɽ�}����?���>e�>X+<?�5B�z�7��E�d�(�o�����d>�I�>,[[>�?�>�]����t�������j��f1�E,�=�b|?�ct?҂?V��;h^ �Hb����0���=�k&�n��=��,>�^�>�_���$<�1�.�F��?�$S
�DT��z$�
�,=��:?k�|>U�h>U��?��3?z+��u������[�*�q����v>n��?$�?��>�h��Z(����>z�l?.��>G�>h���:Y!�t�{��ʽ�$�>;ޭ>v��>��o>+�,��%\��k��B����9�Y��=�h?ہ���`���>FR?��:�aG<Xu�>�v�ٸ!�l��X�'���>~?���=H�;>~ž&$��{��8����%?�?W����X&��9E>�.?�N�>]��>�?`�>�2Ⱦ8R˼Ճ ?s�]?M�C?�=?[h�>��]�~J½�ʬ��]"�OD6=�Mx>�hz>��=N��=g�0���^�ݘ0����=�J�=���-u��9$�;����p�:�,=�r.>��ۿ�6K�Ӽپ���%��Á
��Ɉ������������E�����x��0�u$��uV�>b����^�l��G�?&�?����o�������������c��> �q�gy}������Ӂ���?�h\���b!�)�O�Fdi�{�e��M?7���6͝�<r��m�up(?^#G?̲.?
Z��v��	�����=�|>5
�=8ݾI!���ÿ|�M�}?9��>K�Ѿ'e9>a�>"t�>�r�>���>񆡾��W��|����>_�^?b�1?gz����ÿ�?��mw�:3�?��@��A?�%(�&O�1@=��>�h	?`%A>׊4�,q��������>�1�?�ŉ?w�n=xFW���ռ?�e?G< D���f.�=ӳ�=�=f���'Q>��>�j�b�?�L!ǽ0>���>�-�����Y�S{<��c>f�ƽ���6��?�o\��	f�i�/��r��cp>c�T?�d�>�g�=Z�,?�VH��?Ͽٹ\���`?g��?�y�?�,)?S�����>��ܾ��M?K6?qt�>�&�M�t��6�=�.׼�oW��㾻?V��L�=��>[�>�D+�[n�c�O�)L��	3�=X��D�ƿ� %����j�<�(��;Z���潬ª��R�=��&�o�g��v i=�y�={�Q>�Ȇ>�cV>��Y>�:W?��k?�{�> >c|归���4�;���+,����V׋���-����\�߾2�	�7��`��ovɾjB����<�S��fEM����60��MB?+}�
s�9�a���~=D��N���>��K������8���`��8�?
?$~��-`�#��>��PT�;=?�������Fz���f�(JĽ�_>,��>�W=8�𾿬`�@a���/?�b?ϊ��U���1�= |��=�3?)m�>�ʙ=?Z|>�S*?��o���Y��ug>�Y>���>Da�>��=�����&ν��?y	D?ح,������$�>�/Ͼ�c��o�o@=	(��)���Z>0O�=�n��|K�*����H,W?Uc�>\�)�%��9t���	�!�?=lx?�?!s�>=k?/�B?�d�<������S�e��u=N{W?S�h?p�>Wa����Ͼ������5?�~e?v�O>��i��C龋�.�����?�n?�!?�����}����5��tV6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?s�;<��V��=�;?l\�>�O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������Q�W=v�B���?,D�?h�m��%�=�w�ܢd��b�zk��Q: >���E�������;�NZʾ���lA�"�<!9�>I@ 	��4�>X(�@)ݿ�3ǿ�Fk����?��y?k�>�Cg�bG���t��t��LD�M�+��yw�Ad�>��>C(���h����|�� <��������>%��O;�>�*]������>��F�<K�>]/�>���>��½�࿾���?S��clͿ�О��	�#Z?u?(g�?�??{;�q�U
��M���vF?�q?��X?��B���^��lR�O�w?���Wg(�u��M=����>�<?�A>�ؾ��E��DD>�:?���>��.�Y��mѿ��v<�?��?����T?��?ʶ�>��%՜�;�j�7���
��ˍ?(e�;����p�C������l���>��D?�eY��X ���_?(�a��p���-��ǽ�ա>��0��[\�2��x��Xe�����Szy�n�?�V�?�	�?����#��%%?�>>���i4Ǿз�<ٟ�>1&�>��N>٥`�z�u>:�	�:��	>���?r�?9g?h���P����0>��}?$�>��?�o�= b�>�d�=�𰾹-�xk#>w!�=��>��?��M??L�>�U�=��8�v/�<[F��GR�2$�"�C�"�>��a?�L?�Kb>W��[#2��!�hvͽc1�5O��W@�A�,�z�߽=(5>��=>�>F�D��Ӿ��?Mp�9�ؿ j��p'��54?0��>�?����t�����;_?Qz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>;�>�I�>E�Խ����\�����7>0�B?W��D��u�o�x�>���?
�@�ծ?ii��	?���P��Va~����7�g��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=9M�>Μk?�s?�Qo���h�B>��?"������L��f?�
@u@a�^?*FNƿ)���B�����N�;2���N�O>��H<q<��L�=��ڄ�=$K>�ҥ>Ͻ�>h2*>��>��v>��$>Y����"�~O¿���	�����[���O���]H� �콒���Â�J�̾�3E��5=��~�ӽ�Fx�C%�YP�=�U?0&R?M*p?l� ?�y�l>����L�=�E#���=�)�>Ka2?��L?z�*?���=ڻ����d��[��6&��*҇�jY�>i�I>Av�>�'�> �>�)�:�I>��>>���>.>Rb'=sK��6&=��N>�[�>���>�O�>;���8H�嫿���I!a��f�����=�?H��0������g��C��XY�>x�B?]=��k�0'ҿ����r^?���0�
��8�%��>k�F?��W?Z�l<3�6��YN�DT�>|���}����7>��O�xn=�I:���f>v�>��O>���=8+7��'��?���X��_a�>ԋ:?Q�����='����-�������>uM�>���=V���핿�zQ�rU�_��>��/?Ơ?��� mϾ?2��+���><\=>F˫�$�(<�,�=�l=�ɟ<&u�?b5���<��i>��?��=rɽ>g&���� á>�|>4��=^YP?r?���=.�C�u?0�� �j�>�6?-f�=���=c?�qp>�> �>�2�˹�M���Z��>pu>i*B�˾!�k��f����H>��<s�t���s�?��"�~?��� 䈿�뾲d���lD?^+? �=_�F<��"�6 ��qH��H�?k�@m�?��	��V�H�?�@�?��d��=!}�>�֫>�ξ�L�۱?�Ž+Ǣ���	�9)#�pS�?��?��/�Zʋ�Nl��6>_%?��ӾNr�>�~�}W�������u�'$=���>�2H?�F��gvP�x�=�x
?U?�X򾐨����ȿ�~v����>��?��?��m��;��@����>0��?�cY?�^i>�b۾#SZ�օ�>��@?�R?��><�!�'�K�?d�?책?r:=髞?��?V�?�n�>�<�;.���b��� >�'�<#��>�k>O�=I`���G���掿��v��Gr����>Zj�=��>�J=I���(a<��r�M�����B�>*ѐ>�E=)͸>�8;?��?A�>f�����\�d�'?��|�K?���?-���2n�wL�<��=�^��&?�I4? l[���Ͼnը>ú\?g?�[?d�>.��N>��;迿~����<e�K>4�>�H�>�$��	GK>��Ծ5D�0p�>,З>�����?ھ�,��kZ��5B�>�e!?���>�Ү=ڙ ?��#?��j>�(�>AaE��9��Y�E����>ڢ�>�H?�~?��?�Թ��Z3�����桿��[�w;N>��x?V?rʕ>a��������kE�;BI�@���]��?�tg?pS�/?<2�?�??a�A?)f>և�)ؾp�����>M�?�1�GV���C�G�����>�?^�>|��=^����"">КX�~UȾB�.?� F?�$?�־K_�8�2�|x�=J}�����;�G=G(�=��I>&ǎ>]���L�=2�Z=|�=�]z��;1۽����J"�=�>���ǲb>w�+?�?_�င��r�=�Ws���C�T%�>��M>�=��H'_?�#@�+C{�L�������#T��׍?2��?Ų�?A���2@h�O�=?$�?T?*�>D3��*�޾F�޾�wr�*�v����@�>�f�>�A�Z>�D2���w��5��+�Ž�M|��	?'��>�)7?�� ?�+�>���>� �;K/��S��)��F�S�$��=��w6�2�؜�v.���"�=�¾����5O>�i���7�>� '?0^�>��>���>F����I�>°�>�P�>Q�?Σk>�=#>�/>z��<ؘ!�XR?l�����'���辰���DB?fyd?X��>.�f���������?���?�c�?�u>}�h��6+�s~?A��>n��}o
?��;=�-�C�<tG��t��O���hM�D܎>"t׽G�9�� M�;�f��K
?��?�p���-̾�nֽ�楾�h�=7�?^F0?�A�҉A�˖p�tUW��4P��M�b=�e��y�"��1y�f������₿�!���s=�&?x��?�F�ؕ�H���p�!<�ɴ8>8�>m��>�o�>�6>)�@�-�|Yh���(�ֆ�����>}�v?���>��I?1�;?)rP?8iL?`��>>U�>n8��}e�><��;i�>� �>N�9?��-?10?W~?Rt+?0c>
�������{ؾ�?�?�G?�?��?�ƅ��ýe����Uf��y� ���	�=-y�<��׽��t�¹T=T>k�?i��29�&�����w>�0?�Q�>��>!���J�z�.x=�Z�>J?�W�>�s��f�bR�w��>�}?b��f=�T&>L��=/��83��צ�=@��ׅ=��:�&!���<���=��=mI���:7��;��H;��<�t�>F�?���>�C�>?@��� �m���d�=`Y>�S>�>�Eپ�}���$����g�_]y>�w�?�z�?�f=��=��=�|���U��u���������<£?7J#?XT?N��?S�=?>j#?��>8+�aM���^�������?1&,?.��>|��&�ʾ�꨿m3���?�T?�-a� ���.)��¾�Խ��>�W/��,~�����D�>l��q��g���n��?Ӽ�?��@��6�vj�!���dV��-�C?�"�>h�>�#�><�)���g�v*��$;>ќ�>zR?N"�>��Z?9�?�)a?�6q>y�6�=s���H��u-�<	�?>�2??��?.ua?(ɯ>�:�=?�t�j>���p�Gl���ӽJn�GUn=��4>S@�>��>�>��=������,I��k<�>H�?���>���>�,>|�ֹX�5?��>��Ǿ]������7H����<��j?D��?��?�:h�3!��62���Ͼ"��>À�?&��?wp?hE�6k&>��5���پh���S?��>>м>	�n�T��s�=�?�9�>v��c���U��]�=ϐ?��Y?G|>#rſ�q�@�r�������O<�����b��'���[��4�=B���P�$���?�X�Q㟾�a���k������S�}����>fÇ=��=ǻ�=s��<�]ȼ�%�<#�N=�<��=��f��lj<q;4�"���F��	׾��R<1[K=Zuܻ��˾x�}?9I?��+?6�C?H�y>e;>�3�y��>����k@?�V>T�P������;�1������z�ؾ�r׾��c�tɟ��J>NhI��>�63>�/�=�z�<��=�s=tю=��P��B=P�=[M�=�l�=o��=L�>�R>P1w?:�������}2Q����f�:?B;�>���={ƾ "@?��>>�/������]�T(?L��?�T�?��?�ni��\�>g碾;������=�𜽠2>(��=��2����>��J>K��vF��b���3�?�@4�??�����ϿD^/>���>����U��#0�����(w�����>�*�Ӆ��}��>�h��lq˾�Y.��M���D�>2XU>D`:�x8<�>��=�pǼ+7J=!Ѕ=�>xNV>W��<�;��=_��=��N>�
�>�t=���=�#��Þ=�w�=�c>3�
>��>��?��;?��f?5��>�����������nfZ>�I�=Kƥ>�>0�v>mә>�DG?LF?�>?FD�>��<<��>�̠>(jE������󃟾 �=Q�?�x�?ʡ�>��\�ު��~��2;�a���?�qA?�?H:�>�U����HY&���.������6�X+=imr�^QU����il�ȯ㽵�=�p�>>��>)�>�Ty>��9>��N>y�>��>�6�<�p�=�Ҍ���<#��³�=-�����<ErżMp���j&���+�������;讆;��]<���;Gy=D� ?D�R>9�>�U>]���Y->0���F�5>b�þ�>��cp�����x�7��QO���=�/�>�%�=����k?`�*>���>���?�N�?���>f��'��짿����_*���L�<�n�>p�I���� _k�4�S��@쾴$�>y��>�`�>��b>&���@4��N5=B�z���/?�⑾#I�<	:������z��r��c�Y���)>p�]?V��r�>��o?X�m?)�?�k�>��&���J=+�8��?���C�UJݾ	8��@?�d?X��>���B�R�zH̾t���޷>�@I�/�O���A�0����ͷ�5��>������оi$3��g������ݍB��Lr�?��>�O?��?�:b��W��DUO����$(���q?�|g?�>�J?�@?.&��z�r��v�=�n?ų�?R=�?�>��4���|�N=�>�?{��?2�?U2m?n}�����>>(�v�=�=;��=��d=��S�k��=,�>�?EQ?pw���
�@Ͼ�8 ����^+P=�鮼�\�>�~>00B>n> �>�=}>Yy�=�G�>�n�>❐><Ǝ>�v�>"��Q~�e(?�2>f�>�H?"�>�;(��!H��Ȗ7�'�ƽ�x��9���1�7_�<�N�>��=RT�=QL�>����E�?}^>'����~?����rR=#D�=P��>hoW�A1�>���>���=$ۣ>L�>�/>Z�c>���=`�Ͼ�a>H��`D!��A���Q���;��x>�"��-�+�������I�g߲�#k�vAi�����O=����<Տ?c���i��(�=���\�?���>G5?Y�����j�>9�>&�>�(��jݕ��v��,�+��?�\�?�:c>��>�W?�?L�1��3��uZ���u�((A�ke��`�N፿霁�ۗ
����_?��x?�xA?�P�<�9z>F��?��%��ҏ�a)�>�/��&;��F<=+�>�)����`��Ӿ̺þt7�`IF>1�o?�$�?Y?TV���U�,�">�8?�/?��s?0?Q�9?8)�|#?�e2>H�?��	?Z!4?O�.?\�?�7>���=�
ܻ�}!=���珉��Iѽ7�ʽ<�����2=��p=�GC�5��;FR=u��<�>���r˼)��;�$��ش<ʖ?=!.�=�l�=Wަ>��]?p�>�W�>۸7?"���h8�����$/?	G;=zc��XԊ�a���&���>k?���?OLZ?Ad>˚A�H�B�->(<�>�p&>rn\>3��>��ZE�l/�=�'>W0>%S�=��L�܌��l�	��B�����<�S>~��>�m>৶�ɵ>����+ׁ��o>5�����<�,M��3��.����>TJ?h�?���=���y7���&\���?�
2?�xB?�R�?�@�=iu���/>��O���/�!�>�'��o�졡�����JQ1�f>e<�%�>}Ė���Xb>wC	�̒ؾ��m��H�t�/Nl=(��c�G=q��*&׾5p{���=�->Z����� ��~��e����H?��]=���IQ���R(>1��>7-�>D'h�h��c*<��M��H�=A��>0%?>������ƘG�+C��0>A�U?�#?|��?xh�a�V�MOw�;�>��	
Ƽ�?r�>��?g�>=�ʅ><��D!�d�S�E�V�?��>A;��a��Ū� +��>�Bz�>�?_m>��?9pS?m�?�f?\J?'P	?S��>���t,��S�+?�!�?� >��q�]�6�>��Y�`?�N?�S"��y�>�?��#?D�?\5k?��?���=�V޾ї;� ��>*[�>Nd^����<yI>Wf/?��>�_?�|�?�J>F�-�;���o7��ly>�w?>�;:?y!?��?�5�>�R?�����ܼN/�>��R?�Zf?�J?@��=��>K~>��?Ί^>�K�>h;�>xM?w�R?fс?�B'?��>h�D=�J��IO�D;��xc��*F�=���-<�=��m�����ν��<�����!�<诌�!/��ia.����;���>Cr>`2����.>M�ľ[)���Q@>Ǽ�?��1��F�:�6�=��z>]�>�>�&�3@�=- �>���>���|d)?�N?��?�V�: b��ݾ�jL��F�>P�A?�g�=u�m�򲔿f\u���~=�o?�]?`V�ԗ��L�b?��]?=h��=��þ��b����l�O?G�
?H�G���>��~?c�q?X��>��e�(:n�'��Db���j�1Ѷ=Zr�>JX�P�d��?�>k�7?�N�>B�b>�$�=uu۾�w��q��q?��?�?���?�**>��n�O4࿳���	��Mmd?���>�j���P;?�E/�&;��gZ�������Ծ��>��u���`���0��7���
��L>!�?E3s?S�q?qK?���A�]�F��`{�y�d��������D�=�$�'�6[�o�}���.���������li<�Ԩ����ҵ?��<?�?ؽ��?���8 �'W���~�=, �����i��=if%��V�<>�,=����R��щ���6?6-�>Z�>�.*? VW�s}��� �R�&�p�m�>�'�>ji]>(��>�Ƚ2�!V�� ˾��(���g��=��z?Ȃj?�Ȇ?���T|�@����@$��~�=/�o�nkl=7>a��>���������J��)J��0�'5���l���>�J<?��1>�e�>A��?Q�?���b���`"r�1@��jg��T�>m��?�G?��J>����*'�N��>��l?��>�>����sY!���{�JIʽ�F�>@έ>o��>��o>�,�\�Nc������,9�zB�=��h?;|���`�م>XR?�`}:�G<�}�>k�u���!���C�'� �>�?���=�{;>g�ž�(�ѣ{����Yj(?�7?����%��GR>�9?���>q��>��?[\�>���m#=Z	?CZ?��B?�=?���>!9<y���ܢ�aC�:�==|A{>ŷ4>�Fp=���=��� b�̇��ٓ<_B�=�hm�����<X;.9F�_<���<�9F>8lۿ�BK���پ����#>
�_刾S����b��!���b�����\x�z��G�&��V��1c�ڣ��n�l����?=�?}���.�������������>n�q��a�'������F+����྄���yd!���O�&i�߾e���V?y?��e˞���x��6d���.?#,?�=?*���#Oc��� ���>Lf�>�	=k��X�����ɿ�/:��_�?�N�>T"�tԀ�i֟>p�?���>�Wr>�������,��Pt?3v?��>����Ŀz~���"��e�?G��?0�A?��(�m��Q=���>�		?�=?>��1�������,c�>K5�?YΊ?�Q=�VW���c�e?�<�;�yF���ûP��=�m�=Sw=���0�L>W��>���TA��ٽ=A4>��>l7"��D��@^�M�<Xw^>��ս����2Մ?+{\��f���/��T��U>��T?+�>�:�=��,?V7H�\}Ͽ�\��*a?�0�?���?#�(?:ۿ��ؚ>��ܾ��M?^D6?���>�d&��t���=�6�/���r���&V����=Q��>Q�>ɂ,�����O��I��|��=���:�ƿ� %�J���L�<�5��עY�9��|㩽��S�.���.o�M齕�i=D�=`�Q>l��>��V>G{Y>VDW?�k?uT�>ǁ>�g彨�����;ͪ��x�����g� �r,���[��߾�	���j��=gɾN�D�탵��U������u%��i��u/�S�2? >�#Ⱦ}�J�7Յ�=k�3D}��T{=H���S���<�<�Ms�C�?ƍ?���_�y������v2��'\?�{N��K��s���A4<�O�y�8>���>y��=Ag��JF�?�h�!�6?x?����Mt�ȶC=3t+�P�X=��"?fG
?��=EJ> �3?��>�םN��Ԕ>��+>E�>���>z�=L����3=��?G�_?�7���ڊ�x߯>�+<�G�����ý�������q���֙h>��+=��;�-2�u)佺�<�U?���>s�&��%�������c��B[=w}?�?��>g�\?Ʀ=?�g*=�㾣�J��J��C=-	L?�+c?��>������ξ�q��bM2?��`?�a>"FR�9���<�1�7����?�3u?,?+�%��q{�Yߑ�=v��">?��v??^�L/����x�V�F8�>}�>���>��9��ų>�U>?3�"��K���Ϳ�Zb4��v�?�@���?�3P<�(&����=:�?��>��O��4ƾ���������Wq=��>���'�v�� �ʣ,���8?
ȃ?i �>:^�����$o=�\���?=��?�ҝ����=���So�	8	��P	���=�!9�T%�;\'�D|D�Fo۾�D�@:f���;�,�>=@5�����>�C��;޿��ɿ�ۂ���޾��>�8�?�g�>U���6���r��{�*�H���@��r��,ء>��I>_�'<h�b��~r�d9��
�v�>L�<���>a�F���dAx�3�F��x�>�"�>��S>�ڗ��Fľ^��?�(�Q�ο����h�>?�?��?��8?M�=t�o��66�
°;O�N?�mw?��_?%ջ��|���z�?�/Ⱦh]1���(�%�EȚ>h�/?��$>";�t<1=:�>��?�
>�;��ɿHȿ˘��?b��?�V徤c?cƢ?�?��)�5n���O̾/�$�4��1�w?�w=����'^��ـ�A���<?zÂ?�R�P9?��_?)�a���p���-���ƽAڡ>��0�aa\�7��ץ��Xe�����?y�n��?�]�?��?��� #��5%?��>p����8Ǿ��<~�>O(�>"+N> ;_�z�u>L	�i�:�sh	>���?~�?gi?ѕ������xS>A�}?�$�>��?�l�=b�>lZ�=��L�,� n#>�-�=��>��?,�M?�J�>nZ�=�8�Y/��ZF��GR�$���C���>��a?��L?pGb>e���2�F!��sͽ�g1�J_鼅Y@���,�U�߽>&5>��=>�>��D��	Ӿ�^*?L�!���пT����޽@�:?e�>n'�>��龰2��ɘ�<um`?�0�>&��=��}b��'66���?U��?��?��Ⱦ ;_����=�6�>�a>8�ͽf��e���>B?:�f����r��=W>�!�?AA@㻬?��f��	?���P��Ma~����7�y��=��7?�0�G�z>���>��=�nv�⻪�[�s����>�B�?�{�?1��>��l?o�o�"�B�T�1=M�>��k?�s?�Yo��󾖲B>h�?2������L��f?�
@xu@T�^?)q{��߃�����K�����=��B=�:Y>D����>�ӹ=������,�:'=x4�>T8�>yk>x^Y>���=�X�=� }�tV&�<Ϳ+���>W�7!C�����-�<e��g��W���d����x� >^��;�#��p=�,&꾗������=��U?�R?mp?ދ ?��x�h{>V����d=�y#��Є=�.�>�e2?��L?��*?��=g�����d�(^��65���ȇ���>;rI>8y�>M�>��>%͓9��I>�(?>���>�� >�'=��ߺY�=��N>�J�>��>C}�><`= k>������ʹ�Է`�̟���$`�?�@��o�?�n~�ʓ���ξtI�>`�3?�O7>�O��4�пM����78?K۝�;������v1>st/?d=;?7�O>��ݾ����>*�l��� ���>��&��rҽ�u ���=l��>Ѡ�=��<�<��>5�i���-��$G�>��??��ƾG��>�����C��\*��d�>�:�>>��=ڭ��^����P�L��<�2>�Y?Ww�>��?�{ �伌�g�]���=|W�>���<���o?�=g0�E�����-F�=����>�?R�>�:��K��>!❾�>u�iH�>�rH>3�b>R�7?#�?\�=�b��#%�V��@q�>r��>��.>�=WP1��>�$�>s��>9��u���ܫ��R����|>Y��85���Ƚ���=������=�F껥�)�Y�L�K�=�~?��� 䈿��f���lD?P+?G�= �F<��"�A ��tH��A�?j�@m�?��	�٢V�%�?�@�?�
��÷�=�|�>�֫>�ξҔL��?�Ž`Ǣ�˔	�)#�dS�?��?��/�Wʋ�=l�86>�^%?��Ӿs��>X��W��4�����u��+#=޼�>��H?���!}��B��?�?���60��t�ȿ�u��P�>�L�??��?DCo��Й���?����>�?�Z?9W>��ܾY�6��>�:@?�yP?���>���\�0�%3?���??�?+'����?]��?�6?�E="���ƿ���P�$>!�u>�j�>a �=�35;�0o��c��Q��s��7����N>�s�="��>��+j���=�T��g��y�<�Ú>I=�=��2=�	?��G?��>$gr>@��<N�=�����nھ[�K?n��?��2n��-�<+��=&�^�G'?7J4?�[�2�Ͼ/ը>��\?V?�[?9c�>��+>���翿x}��嫖<m�K>3�>H�>9$���GK>z�ԾJ7D��n�>�ϗ>p�C=ھ�,�����?A�>�d!?���>�خ=z� ?��#?�~j>�/�>�oE��6��2�E����>6��>�3?1�~?��?\����H3�����8⡿$�[��N>:�x?mS?\Õ>c������NE�UI����y��?Wg?[��??/�?a�??w�A?��e>a��:ؾ�׭�&�>���>��ܾ�W�KY0� [R��?o0?=C?�=NS<��5>)9E�+k����8?e�P?��J?D�����Z�t�"����=�f�=���<����%"���G>ƒH>P��� A>(s>^�=��� >�-��ܾb��I�f�3>�je> �:5>��-?O�P�	�|���=0�p���A���|>{<>oþ�_?�>��*y����4���bc[��4�?���?�-�?���I�j��_@?nM�?�?���>oҮ�/y㾴x�Wt��t��a�3�=%w�>�,��{ھ�ԟ��ҩ�����rս{G���?���>�$?\�F?t�>��>>�پ�E�_V��*$��wH��n-��/:�;;D���]뱾���:7��=Ceݾ��t��J}>��D=�{�>U�>�q\>^�>:�>� �=V�>'J�>�w�>��>��O>�=^>�I>)~��t�&��VR?�����'��v�	Ȱ�kB?g^d?�@�>"f����������?ރ�?+`�?7�u>ٓh�g8+��W?q�>۩��B
?[:=�����<?���L�9���0u���>��ֽ��9�o�L��f�� 
?��?6$���-̾1*ս�u���l>Ge�?�V1?%���a1�?�b�h�]��Z��_����/��D������r�EE��؆��ֆ�?��S.�=͔?���?i�ݾC���.��j�r�0�N��#>~>�>#ճ>��>���=�J�?�*�7 ^���'����]��>�q?ʋ�>��I?�;?�rP?�iL?���>�`�>�2���i�>�p�;a�>�	�>ş9?��-?�50?�{?�v+?[+c>O~��*���ȁؾ�?[�?eG?�?��?]م�ShýfE���=g���y�{u��v�=�!�<��׽�+u��T=%T>m?����'7�q��7p>W�5?�W�>3��>�ǌ�x}�Q�1=�J�>�2
?�c�>V�����n�Z�Y��>���?�OԼ��=ߪ(>�:�=��{���l�=�������=�^����D�'#<X.�=���=���Vl�K�	<�Q�<���< u�>4�?���>�C�>�@��/� �_��1f�=�Y>1S>\>�Eپ�}���$��m�g��]y>�w�?�z�?��f=��=��=}���U�����F���:��<��?:J#?XT?\��?s�=?cj#?ӵ>+�iM���^�������?w!,?튑>�����ʾ�񨿿�3�ڝ?p[?l<a�S���;)���¾v�Խ��>�[/�b/~����1D�E煻������ ��?ؿ�?�A�A�6��x�Ͽ���[��k�C?�!�>Y�>��>L�)�{�g�z%��1;>��>|R?r�>��O?�1{?�[?CwT>�8��.���Й�92�">�@?���?-�?�
y?�a�>A�>��)��ྦྷL��e��#��ۂ��NW=�Z>⟒>z�>�>���=\�ǽSf��n�>�q�=�b>ƒ�>���>��>kjw>�8�<QG?���>��J�� ���x����9��Ru?2�?��+?�=D�b�E�W)��,^�>c�?�?�)?�S�T��=~=ؼ=�����r���>S�>��>�[�=l�D=9�>���>�{�>8���8�678�I�N�|�?�E?µ�=˧���:n�������fÝ:�����XX�������d�L�=I���@���3K�;*����� ����h��[��#��>��=��=f"�=��0=�to��L�<{�<��<v�<r�����<�# ���3;=ɒ�V	:�KZ;�h=��4��˾X�}?�1I?�+?�C?"�y>8=>��3����>����@?�"V>a�P�Z��p�;����*����ؾ;s׾s�c��ş��D>�I���>�C3>y(�=9�<Y0�=B:s=3ێ=�+M�sV=I3�=�J�=��=K��=�>�Y>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?~�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>q��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>���=X�[�j�V�p6A��c-���-�ռ`P�> �&�t��^?+	�_^��3�=��=>&�>�l�>K�־.�D���X>-����60=C{O>ފ�>E��>�.=&�A���>u$�����>R}Y>�M>K�=�;����->QIi=m�>���=�r�>�?��1?�\d?{�>	op���Ծ�c��h�>&�=rb�>�Y�=�H>C'�>m::?=�D?lrI?�D�>�ā=ɷ�>Q�>1.���o�W���X��\��<�/�?��?�5�>��A<��9��[�e;��˵���?zM1?u�	?�I�>eT����Y&���.�������&+=Cir��8U������j���㽦�=�q�>���>��>�Vy>��9>��N>j�>�>�Z�<�q�=
������<� ��嬄=�Ñ��y�<x�ż�:��x(���+�����h+�;���;��]<r��;H�=�m?�j�>Z}�>��S>!0J��?>����J���t=<���qQ�φ�y����
1��/��L4>1��>ߝ>���\)?�l�=q��>�p�?^o?��>���sξ@���P���A��-w=XD�>�q�d���� �P�߾���>T݇>�N�>ɤY>�a(��5��o=�Q��6��`�>퇊��t�W�<��={����xv����P�q�t=�MH?�����/>w��?aM?A�?��>)R���ؾ؜*>y�p��8K����T���r����j$?9�4?���>�I�/KE��H̾����޷>m@I�"�O���Q�0�;��+ͷ�4��>������оd$3��g������ލB��Lr�X��>�O?��?h:b��W��HUO�����(���q?�|g?C�>�J?�@?&���y�wr��w�=�n?���?L=�?r>��=p ���
�>0k
?�b�?w��?�s?C�B����>M�~�;Q>���;!�=0�>�_�=�,�=X?�;?��
?�N��J�	�T�����hpd�a�<��=ȓ>n$�>řw>K��=` w=4�=|�^>Gy�>��>qKd>Uv�>��>��	�������/?Ư�>&��>��%?��>��4�V�;�(���+c�e!ݽ�u*����@:3�;�>�s�����>�m�=m�>Յ���E�?J�7>���ȵ?�47�CG�����>��D>��4=˜>�T>��H>9��>S�W>�9�=<1�>.�1>ɫ��8�.>���H��SX�"�F�V���f�>;�o�������F����q���i���g��iw��9=�o�=��?�SX���X��1����<ޡ?���>v?�S;��Խ��&>Y?9ܶ>2��߭������G��dhz?g��?�;c>��>/�W?	�?�1��3��uZ�
�u�i(A��e�O�`�}፿
�����
����_?�x?yA?<R�<,:z>C��?��%�fӏ��)�>�/�';��><=W+�>?*����`���Ӿd�þ8��HF>}�o?+%�?gY?BTV��r&� �>�b3?�6+?��q?�\-?��6?Er��g ?g?>�s
?j�?�C3?�.?
8?x�A>R�>C�9��A#=�ʂ�1(��lcƽ��Ͻs�1Yv=j}c=(��;�l;o43=�4V<��м���%�:%\���O�<V�U=�̖=�9�=}��>R�]?�8�>ޕ�>߻7? ��Oo8� ���9,/?!�9=����Q���¢����b>+�j?���?JWZ?�Wd>Z�A�/�B�r>2W�>ZN&>�\>+a�>)>｝�E�@��=%;>�F>U�=?WM��ʁ���	�����Z�<,>/��>��{>{���^'>���Нz���d>��P�4+���iS�(�G�^�1���v�td�>2�K?��?[��=�{�1���
f��)?&.<?�M?��?TԒ=��۾P�9�H�J����$�>�Z�<2��ʜ��]����:� �S:"1s>_���Ɛ���A>���d|־``���Ko����M�>W]�tb.>�n�-���������=��q>�MҾ.��Ά�������{U?�ɕ=v���p���N��WJ�=:��>�>�>�4�=(Ƚ��<���Ǿ�>=���>�6>�<�����`�������>T?Ǎz?��?$���M���t�*̽�7�T����=J/?��>�2?+	�=s�>�î��2���K��A��2?��>�ܾ��D��q����W� ��?o��>-E>-?Lz5?[~?��j?��Z?u�>W|�>�W轈T���F&?FX�?��=ӽ�CV��9�d�E�(��>,$)?��B����>0�?��?�'?��Q?�?��>�� ��@@�MP�>Ԝ�>�W��@����_>�mJ?�ֳ>�Y?���?��=>��4��n���y��{��=~R>�[2?`�"?��?}�>$��>4���|=G�>�b?�K�?��o?VO�=^�?�~2> �>7��=&�>Q��> �?2[O?VWs?�aJ?W��>�2�<蓪��l���Ys��g\��oi;�aE< �=a���l�������<��G;�b����\�@��.�>�G���Z�;g��>�1s>	5��x�/>�ľ����A>:���MT��Jn���O:���=덀>/?��>֓$���=��>U�>ڣ���'?��?s�?a}�;1eb��Cھ��M���>�yA?�=��l�\_��:�u�ɠh=��m?�%^?��W����L�b?��]?8h��=���þV�b����g�O?6�
?�G���>��~?g�q?Y��>��e�":n�#��Db���j�6Ѷ=[r�>FX�J�d��?�>c�7?�N�>4�b>%�=Yu۾	�w��q��Z?��?�?���?+*>~�n�T4࿣���b����^?��>Eؤ��w$?�H�4�оuu���я�ᾡ6��_��A%��O���>%�R|����̽��=��?��r?��r?�=^?�� ��"c��`���!U��O��9�kD�L�B�X7E��On���������}(C=���d�2��?>?���;
?����������ʾ��>7'����E�={q����e;.�0=�QJ���߽�y����?�ɻ>*��>�,/?wZ�p4��Q�E�7����م>s̞>�>��>˃潩IC���R����I�=��>#5>^n?�`?͗�?�_4<���䶐�<1"�&c+>9�l���=|�s>�}�>����6X��0��A9��HN��	���g�9O�o�#�M�?zH>B��>��?c��>�'����]��#N�iuM�~�?T0�?���>�RV>ω��%����>ׇ�?\�=?���>��k��z��4��|�\?q$?5%?RQ:>K�=�����,��3:��tR����>DY?vCC��Ѿpw>��?�����e��kͯ>��(>���S!���X���?c�?~|=\�=�gt�J���P~��<׾��)? �?f���l:#�k�@>�d?bt�>��>�jy?j(�>��˾ B"=@�?&�`?�I?Ӯ>?H�>1�<g޽KaŽ�`�fb�<r�h>�.n>���= ��=�!��-Q��R���=���=��;<dݻ��J��9)��&#<e�o=�P>��鿚+I�"
�U���*��$���R��{�=�8 ��������h�׼u ���:T�a^&>放X�=�IG��}y�-�?9[�?�1��H��Tz��>C����ܾj�?��HNT>�~���#�����1��	�ýo�/�����`���;���)?�k��� ���E���R��?"?��%?S
i?E�����(���)�z5>��<=�d,��]��gY��C�ǿ.���r.k?��>����&�����>�+�>ٗl>�aB>�i������k��Q?�*?y��>�O����ȿ\o���S+<m��?�u@&	D?w�������=���>L�?�y�>F�-����>`��\��>�*�?�h�?��=k?P�<~�0�P?;d=<\m���6�s=�=�A=�j���o>�H�>Q爾P�������D>x>�>jAL�U�`����������b>�x =F��=�Ԅ?uv\�)	f�Ț/�zR���E>Q�T?,�>��=	�,?o6H��sϿ��\��)a?�+�?]��?��(?Z翾���>��ܾ �M?C6?���>eh&�^�t����=Q߼����ÿ㾳.V��J�=���>��>�y,�E���dO�	d����=�f�0rÿ~�(�a�!�� \;`���VD��>�����1|��.੾�>�70��ތ=��>�EF>�>4V>"?H>Gc\?x`d?�t�>>��,����V%ľ��^=�j���������8꡾����ȾC��2��7���}��^T���<�R�̈�w�L��䄿g>5��<?��>a��H[�s�w==u�X���>|G��=���_/��2f��]�?NZ.? ����`�����"�����bN?M�J����M����[<|�6���>#�>8ɢ=��ؾܣL�XU�1
3?}�?D����I��m�)>+����p�=�c)?�6�>N��<>��>��*?��z�@��e>�,>k�>��>`,">����,��T�?��M?����Zq��L�>2��E.�Ed�<r�!>��?�P:+�1�	>�u�z���P��r�6�!>e0W?�*�>�E(�s���c��3j���w=�Jv?�?�_�>�ci?W�C?l�<��E%Q�"�
���v=9T?Y i?S�>Y͌�<;X���8?�f?��P>6�}���ྊ�-�o����?1<k?�?u��"�}�<c���P�<?��t?�bN�0f�������VG���>"��>&�>�{7�q��>�7?���D"��p ¿MW4����?1�@i��?���=(0ɽ��&>wn?7a�>��_���m#��f��e�<��	?-��Os��Si2�'���G?B�?�
?žo���aς=�PM�Р�?���?މ����=���rl�_𾒊&���a=�4��&�:����i>��C۾�Z��;=8�	q�;���>z9@*%�;��>9�0�ݿ�9޿@��0�����T�	j?�1�>�����l_e�E�f��G3�,.���W�>���=��Ͻ�F���ℿ��J�����2�>^lh��3�>� ��B��u����w=g�>�@�>:Ӎ>����˾��?&y��̿񣿞�㾮�a?&�?�{?:�?�,��h�[�ԏ����;�K?��b?�,X?e���.���SŽZ�l?M��R^@�C!�����ؚ>^�-?��>��T�0=�\�>�"?\��=�23���¿�滿c?F�y֬?BT�?�Uپg�?�*�?m��>:$��$��>���^s6�Y7�؟b?Ѥ�=�4۾*�V���u����2�<?q?��;	�.�R�_?Ӛa���p���-���ƽ�ڡ>C�0�'c\�AU��G���Xe�~���Ay����?^�?D�?,��� #��5%?]�>y����8Ǿ��<O�>�'�>3+N>_:_���u>_���:�2j	>���?W~�?�i?ە�������X>��}?@�>E�?���=�6�>Ph�=�Ȱ���%��#>��=�x>�G�?��M?�:�>��=��8��#/�^4F��CR�9���C���>��a?�zL?t
c>�����0�*!���̽�1�E 缌�@�� -�,p���4>Ų=>�>S�D�m�Ҿ�-"?��"�п�搿�-����7?)l�>�t�>��뾖U���D�<ֵf?���>�:��Ҵ�r���	�߽��?���?�X?�p˾u����=�;�>��z>�8	�h,��=��E�\>'�B?p�ὕp���qv��Ys>�ٺ?�Y@2�?�Eb��	?�	G���V~��z���6�I��=#�7?P2�{>���>vY�='vv�(����s����>�M�?c{�?H��>��l?_bo���B���1=�2�>�{k?o^?`q���$ C>˓?L������a��)f?��
@xs@��^?G�pi��x���⯾c/��1Y�=��=�.>�f�ŧ>:�q=PU���=�� >�x>�T:>ҿ�>YbI>�h>�Ѩ=����ω���ʿ�О���J�~�%���׾��<�n�;�A���y��d��Iܼ��r��6�Rg2�t%�#ý�y��=�%U?ҌQ?;�o?��>(�c� >�d��K
�<m�#��B=H�>2?E�L?b�*?�=�����d��F�����t�����>�G>�>���>��>�w�:ߧI>{�>>��>�p>�3=䡴�*�=bM>4�>���>/�>��=pu������N����c���h�;fĚ?;�m�<�P���n�������<�>�7?j��=�gp��Lȿů����K?F߾B��MW�b�>�[?WW?3�ѻ&pξm�k���?����U�P9h%>�����`u���O�I�n>�E?T�>_�>���/����S�� ����>�??5N˾�
���u��{��\��~��>��>E �=��J��f`r��Ou���>e�&?Zz�>�i�Zž��9sn��[>AR@>LKϽ�G>r��>�Y��m���!ј��M�=C�|>qq�>�?�K#>�J_=�>;���+1@�!�>UY>+�>��;?�i?��;�����u�\�~l���d>���>�b>m�>%B�X"�=���>�g\>����|P�R���`�}Gc>����v]G�J>|��lU=%������=�l8=�|����2�M��=�~?���䈿�뾽e���lD?[+?~�=t�F<��"�? ��NH��/�?h�@m�?t�	�ĢV��?�@�?����=�|�>�֫>�ξ.�L�ޱ?��Ž(Ǣ���	��(#�\S�?��?c�/�Cʋ�/l��6>�^%?ܰӾ8�>c�����������t���,=�V�>ZG?`����[��<�I�
?�?P�񾇤���	ɿOv��M�>V;�?Ǟ�?8�m��蚿��?����>�B�?0X?��e>��ھ��Y���>0�@?��Q?�I�>3��f*�(*?P�?���?�ɸ= ^�?Կ�?°>�{>���ſ�����>'7�>���>�(�i�}�Cxk�iD��'���/�Y����Ɲ>C+=�E�>Ʉ��;��
�=���h��.0Ͻz�?4\�>s�c>�5>�� ?���>�t>C�Ӽ�K������Y���K?�0�?K��um����<��=
�Y���?y3?�d��HϾ�^�>/m\?[��?��Z?���>;�l����O���m���<��H>�x�>��> ~x��M>��׾dBC����>od�>����پ�炾��GК>�� ?�o�>V;�=י ?��#?��j>�(�>aE��9��J�E����>��>�H?�~?��?qԹ��Z3�����桿��[��;N>��x?V?Fʕ>X���݃��}jE��AI�����L��?�tg?�S�$?<2�?��??@�A?#)f>���ؾs�����>�1?��$�9����{SZ��6
>P�>\e�>�"�������>w���U"�N[6?�xD?a6?�t���a���jY&=�d�<�1=�=3N�B/�=�i=K��כ����>&]D=׾�����Ʒh;�z�=Y�v>���<_=������&?�sN="���&t=�qY�3�<��`>��<r�ľNWz?B���h���������� J��_�?���?ɝ�?��2<��|���`?�ڌ?��?P�?Y��+�پ�ľ�|s�Tv����8��=
��>L=Q���?�|�����Nu��j��}��d�)?��>�*?j�/?L�u>���>�ؾ^L?��h���%�"�N���L�ڋ.��G��־#M#��Pc���D=����qƐ��!>7#�o>��>���>���>��>#k�=���>�8�=#�>��>ɯ'>�.5>t�c=�ya�T���[iQ?��þ�'�7n�-����C?��d?x��>\���tԁ��k���?�N�?���??�s>eb��(�� ?�x�>��w��
?�.=ր1��4t<�n��t���u��9�zL�>(��"4��O��<X��P?)?i����Ͼ��ڽ��/��=H��?� /?o!�~�D��q�`X��,L��;p�t�k��敾#s�t�w�� ���}����Y=�'?���?���:M��E���}o�©O�X�J>PF�>���>�m�>�4>>h��N7���Z�|2 ���w�k��>߇x?bϑ>�iG?	�8?`�M?6%K?���>��>�����>��<�z�><��>#7?��-?7.?8�?��)?��Y>8�޽T�����پ��?��?��?o�?fg?_'��i9����μ�a��y�<\��;�D=�C$;1q�Dzw�\=εw>��?�a���@��S��Kw=.\L?5��>��	?R㵾����,�pE>t6?l��>��ž�HH����	�<��J?����kA=��E>�<~>V�7>n?n=�c�>�!���t>��p�>V����==�C>jX�=�,�oOR=��D>�Z�=;D">���>��-?E.�>d��>69[��ﾲ�ª<�D�>vh>�>���Ģ��:����i��^>�\�?nr�?�Ͱ=�}�=�e	>J��b;޾R1���t����ӻTW�>�6-?ׄ`?��?�V?:�?��+>�X�8���_���v��">?G",?䈑>��9�ʾ��<�3� �?[?�9a����>6)�^�¾��ԽV�>7W/��+~���,D�����@��E���!��?���?Ϝ@��6��n�-���aQ��j�C?�"�>BU�>��>��)�?�g�^'�j.;>���>^R?cҷ>|7Q?_�}?v�_?A�_>�5�����!9��C��<�&>�j<?���?�r�?�o?;��>r�>ch.�׊پث���|�K@��z����a=�V>`��>I��>�`�>z)�=^%½����+�J���=�t>`��>}4�>HZ�>�G]>��<��G?f��>�������R���τ�p9&��@v?!a�?� *?�o =Y��"-D�����D�>�֧?���?B�(?�U���=Z����R��tls�lƹ>c5�>�s�>���=G=�>�b�>H��>�`���XM8��9^��/?^�E?��=a�ſ�q�Z�q�b"����[<�Ӓ�[�d�k����[���=�s��Ǣ�P����`[��n��Z�������毜�6�{����>�]�=���=���=���<aɼ:*�<qL=��<�7=0r�`?o<��7��ۻl����;B�qb<�J=�:��&̾��}?JI?�+?�>D?wy>O>TZ<�h��>#삽�?��S>p�b������f>������꓾�4׾�V־�)d��@����>��J���>�Q1>��=��<j%�=�}=�:�=��t��z=���=L��=��=�Y�=Bm>��>�6w?S�������4Q��Z罜�:?�8�>�z�=��ƾz@?g�>>�2�������b��-?���?�T�?G�?ti��d�>)��㎽�q�=/����=2>0��=k�2�L��>��J>���K��~���~4�?��@��??�ዿʢϿ�`/>�Gq>,�<7?K�]0�9,��d���ʽy�1?�82��߾���>A�X=�����Q����=�0a>�1��*Z�*)U��o�=�[���<x=͓>s:�>���=�.�R=��=>;.>�P>N�=N��<���9ټO�`=���>�>&��>A�?di0?�Td?�>On�%8Ͼ�	��J@�>�!�=��>�M�=��B>tl�>��7?H�D?r�K?x�>�U�=���>�.�>Ӆ,��m�I`�tܧ��I�<Y��?�Ɔ?ո>�kS<b�A��w�eC>�;�Ľ�a? F1?^z?m�>V�ɡ��Y&���.�o���Մn�y+=Akr�yqU�i��cp���;�=�p�>e��>��>�Uy>e�9>��N>	!�>˩>���<2h�=y����<�ᔼ�ф=>���<p�ż�����O'�6�+�X����;	��;�n]<���;za�<�v?8��>�J�>��>��[��!D>z�f$T����<]��")��X��(�����)�*�#=��>;�>�%=�ŗ��}?�%�=l߰>@.�?�<}?�]�>�t׽�������\�3�4��:�=@��>ɐ��sT@��|��_�^���ʾ|��>Gߎ>�>��l>�,�#?�m�w=��$b5�A�>�|������(��9q�@������Hi�.NҺ�D?�F�����=E"~?�I?W�?��>.���ؾd;0>�H�� �=Q�n*q��i����?�'?���>T�]�D��H̾w���> ;I���O������0�V�>˷�_��>������о�#3�7h������X�B��Ir�1��>�O?��?&.b��V��%WO�����2��~n?�zg?��>�K?\@?2��^{��r��Vs�=b�n?Ӳ�?C=�?�>R�	>���?�>}?�ޔ?��?9Jv?�(P�;��>�H\�a�!>�庼��=�
>�hY<��=d� ?Bb?� ?����b��|/��,྽T<�TV=�0=�N>=Z�>��@>���=%�=L�==�>�bU>��H>�,Y>��>!�>�Ծ�2���+?Cߨ>R��>�)9?���>�8��m�����0=FA����X�����M$�t�Q�J}:>y�9=�)>C|=Q��>ο�r�?'ͮ>:�,�;?�b;�_Y`�5w>��=gt�<�q�>��>/��=��>�7>A�=�F�>���=$cѾ��>���� �jB��lQ��\Ͼ Hy>����z'�A�����G��[���`�:�i�Eׁ��<�݁�<ۏ?�0�;�j��)�������?�ר>��4?���נ��E>�E�>=�>P��ӻ���Ǎ���ᾯ^�?��?�)<>��>m�d?��?�	������h��w��-��E[��PX����@y��`!�3�"��CP?,Qq?.�M?�Wf=C�r>a"�?0��]�о���>��3�RL� A�<��>�R���A��Z��־Z��?�.>/�g?i%x?��#?6Y"���m�]'>��:?�1?�Nt?
�1?p�;?9���$?tn3>�E?�q?�M5?��.?O�
?%2>�=�i��
�'=]6���ȩѽ]}ʽ2���3=sf{=���'<��=��<���u�ټ};�)��
3�<�:=��=��=���>��`?��>"�>ʖ8?W�8�:��@���?/?|�G=2���,7��(���Z�����=~g?/P�?A]?/�j>z@��9���>e_~>��)>\5V>��>�-���d2��.�=ާ>}-�=���=���5W��t�
��a����<\+!>-��>�z>@V����>>p����r��q}>�*��켾�L�V@���"�>a�:��>TI?��?��=�徰͖��=]��$%?X4?��F?���?� �=�`ʾ�&D���A�2M��Ѯ>�Z�<t���������<�t(�;|�b>�i����2Ag>X��z5ؾӀn��aL�@�� ^d=\����=�n�6�Ѿ>"{���=�!>A+������,��4U���L?Kb=H^���]�+���a>���>1_�>��E�%�y�O�?�?L��A��=��>�&D>=	����40J�����>�I[?PZ�?D{o?$�A���_���m��.��0�ؾ=L,>E+�>׊�>�#A?S��=%P�>5���8	��eU��r`�*W�>݃�>����T��ݏ��R�*~-�OK�>�5?Sp0>N5	?�a-?f �>:9�?��>?��>i�H>Y������K&?i��?��=a�ԽĤT��9��XF�`�>�h)?��A�R�>�|?��?�&?��Q?5�?�;>�� �/e@��>���>��W�\��
�_>3VJ?�d�>:Y?v�?!�=>}D5��ᢾm2��1�=f�>��2?/�"?��?J��>��>������=�q�>;�b?�(�?��o?_��=�?�1>!�>���=���>Τ�>�?6VO?��s?�J?R�>��< ���w<��B�r���O����;'�I<2sy=-^��t�B�����<���;��L�����D�QW���w�;?i�>�9s>!#���J0>pž���ZkA>Zힼ�-�����<�:����=�R�>�?ˈ�>[�#��L�=�6�>iR�>u��1(?�?>�?#7B;�ob�ֿھG	L�M�>��A?=T�=s�l�|i����u�Z�i=�m?M_^?�WW�����b?��]?�g�q=���þ_�b�����O?��
?��G�,�>��~?��q?q��>{�e��:n�c��fCb���j�[Ӷ=Ji�>W�!�d��H�>К7?�M�>?�b>j=�=�w۾�w�gx���?��?��?#��?�$*>��n��2࿼"���?��T`?�y�>0��'�.?��@�����Ș��ي�98�c㿾Oã�
��;�����F:h�Gܨ��¤=&~?��p?�~?}Vb?���?c��Uh��v�g�D��y�����FB�%�E��DJ�ǜm�X��ՙ�%��n�<:L���#�%�?��+?݉�H/?�흾�I������D>#���L��O�=T����|!=�=G�?�-?�=^����?L�>�h�>�7?�2[�<�3C���&�A;Ҿy�3>��>�߂>&��>�5S�V9'�0�����9���X��U�m=�Ł?{��?�@�?Пc�EIݾ~����	��m!��ν��=�<�>��>\�Ͼťy����s;'���9��+�����O�)yv=M:?y��=#ʎ>[��?��?�)=�)FN�t���KV?���=>���>���?��>]:5>�vQ�+�@�>z��?g?ӷ>��?�Jm��+���D�ǰ�>�>4�>��>��@��n�+���ֽ���17��I>MW?�܉������>�lW?�����=�[�>���<�P���꾕��J�|>��?���=�4>�*����;R�z���ľ%�*?���> ^��Vf(�m�e>x�? ��>��>���?�W>!K��O���?	�_?u�R?/??���>�
��0��ٽr� �:��<y��>�.<>5=v=���=�$���v����_H=���=����*����a��pY���Ǭ<�x<w�D>�S��BA���Ͼ|#����\@����=�������ʻ�=��>�����6k<=�V��z��3w��,Q��R�?��?N���=�
�����; �3\-?���^T�>�	���G�<9���@�'��=�#� �	��:K��[v��&&?�咾+������<Yľ��?A^2?��y?��/h�vP��˸>6M�=�4=����Ɯ���������5u?R��> o���!�.��>�@�>��Y>яw>�Mƾ�ߔ����?�&?��?8����ÿ�K����y�G`�?%#	@1qD?�*'�T ��w�=v�?T�?��>�C������a��>z�?!Њ?�
?=��`���@�6O?�t>(Uܾ�:3Ik=/�=ߦ�=�b���e>��k>7�g�< ֽi&��&G�>0G>O�*��	f�"L���>C��>�)>�;ɽ4Մ?+{\��f���/��T��
U>��T? +�>M:�=��,?W7H�^}Ͽ�\��*a?�0�?���?"�(?<ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=L6�Љ��t���&V����=W��>b�>��,�����O��I��]��=>	��ſ�����%�u�E=E��<h������\C�����I���������tl�=ë>��O>�sq>�hA>��x>��_?��u?o�>�+%>����	���7о
�y=7#t�B���'���o�;������6�ݾ#��2��v�Q�ȾC�b��d=HqM�xh��{K��P��C�H���D?/U������<�|�V=���2�^�5>>Q:����s�0���c��}�?�v&?<����8c�'�)��=�Ym�}�x?j;Ž&��Z����L<��R=�N>4�>�=��о�Hg�L��1?d��>�x��u����0
>�ͽ��>E�(?c�>m�>��D>�??#�H��"m=�Uq>(n�=WK�>�6�>��">5�¾F�1��?t�G?�W�4�����>�h�1S����	>��6�cW>�r�=�{>>�P޽{��p� >�Ӆ=*�Q>��V?g7�>�)����B�����E�^=�y?��?f�>��f?�E?P�<�5𾮹R��#��]=͞U?�pi?�>����о�j��-�4?�d?��U>�e�96�&0����܆?�
o?�?�u�x�}��W�����w�8?mc{?�zN��z�=�W�5"���T�>��?��P>��޾,G�>�7X?x�8�c�E,��#E�[z�?I
@&��?�v>�1��O.>� 7?�t*>��q���=�O���6>4H0?,����~�1Sx������e?���?��;?�X����"�=�d
��M�?�؏?_q����=���0"y�mK��R/p=L�T<�IC��<|�;
�)A�*����^��'U��>��[0p>=�@i�j<���>��!�����5޿Wd�� l�����$?%��>1�۾su��ot�NH�U?/�MN���AU>ۏ�=H�2��(���ۈ�w)T�1�`��+?��ý�ם>T�������N��u�=�9�>uD�>uE�>#oM��龓~�?F%�@ӿ�ڮ������?� �?��k?�!+?�;>�lGS��6�����=V�I?� T?�tV?x����p��PO�<�j?V���}�_���3�ЬC�+�U>� 3?��>@�,�V�w=E	>jC�>��>2�.��jĿ����Ƅ��J�?j��?#^�s�>Q�?��*?wx�����А���+��2�;$NA?�6>G/���!�-^<�N�����
?ώ0?���V�[�_?+�a�O�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?M^�?g�?ٵ�� #�b6%? �>i����8Ǿ��<���>�(�>*N>[H_���u>����:�	i	>���?�~�?Oj?���������U>�}?�>��?���=[�>���=�ⰾ )���#>���=t�?�`^?�M?�
�>(�=��8��5/�UGF��=R�p�"�C�m�>��a?JsL?��b>����p0��� �7�ͽ'(2�h	��	@��D)���Q4>�9=>}h>>>D��Ҿ��/?��7��I?a��"X>K�@?pW�>=8�>r�%� ~G�M!A>(�k?p3�>[�|��8����aN����?�S�?u��>����x���_�>�R�>��>j��z�ƽ(���mM>�;h?�����o�\�b����=y��?\ @E�?����4:?;�I����r��O� ��Y >�
1?L���Tr>�^?m��=mok�a�����w��3�>�H�?zW�?8��>��f?��m�Z>���k=�D�>ջf?X�?�T��F�� 	D>��?��� �����.Xc?!b@;�@R(]?���yhֿ����bN��Z�����=���=��2>�ٽ�_�=��7=��8�>�����=}�>��d>q>(O>Va;>��)>���L�!�	r��W���L�C������Z�=��Xv�Pz��3�������?���3ý�x���Q�2&��?`�t�=�eW?�$U?ٜo?GK�>�b�q>Z<����?<�?��O=w\�>�@4?U�F?L�*?e��=K���?c��́�M��������>�;>���>ݢ�>�8�>GWD;��;>�!?>ƨw>jV�=hWA=G�:&�H=�MK> ث> ��>VL�>�T>���W��������`�!xz�}���<�?�h��;��q�ǌľ=�U�kJ�>kK?+�=岁�H�¿:��W?Pj	�����:��"�>I�=?)vK? @�=�㎾�~l��Z�>�B*��*����>��%�7�6���+��cX>��?(�>�ɮ=Wd4��,�fy�"�6��I�>��??�ƾ��#�]� �������>}��>���;�8ᐿ3J?�N����v�>*�A?�g$?�K��0��'"�ݜX�>��>�>��K�v�>y�?>�u���7���^��>�4a>Gn>�?�} >�w=5~�>�\���G�ካ>�_H>�%>tv>?�� ?Tk��\��L3i��� �0l>{��>��i>�>P�Q�(~�=��>�g>e+�Ԧ����w� �k�D>��
�#���ݨy�l�=����?��=�)=� ɽ�.�tv=��~?Jz��(������m���eD?�/?@I�=��E<w"�j��[��=��?��@�g�?�	�7�V���?k?�?�0����=Lm�>�ܫ>�ξ��L���?��Ž�Ȣ���	�S#��R�?�?"-0��ˋ�rl��/>{g%?��Ӿ�>��)��]����w���]�Z�=�a�>o�E?X���3���ˊ���'?�\
?<�־����Sɿ��h�A��>´�?��?�_x�����-h.�`�?a�?�BF?�Gu=D������S�>��)?�;M?��e>y���qX���> ��?'��?��<껨?�τ?�:?�7�=��4�g*ɿ[����E>~�G>�>H+>Q��2�z�Dr���I\�MP�=���*QJ>�{ƻ�۴>B��1m�u�=L�����`�h�>�� >��C>O�?���>V��>�l�>�����V�p֐� Q��G�K?P��?����1n�S�<���=o�^�S%?7K4?8\���Ͼ:Ҩ>��\?;?�[?�e�>,��=��-濿!}���ɖ<�K>�2�>vF�>F��zJK>>�Ծ�9D��t�>.ɗ>0���E>ھ�(���ģ�J<�>#e!?���>5�=͙ ?��#?�j>�(�>NaE��9����E����>���>�H?��~?��?UԹ�=Z3�����桿l�[��:N>��x?�U?�ɕ>@���񃝿TE��AI�����9��?�tg?-U�)?2�?��??:�A?)f>s���ؾ�����>;r?���AL��X[����_��>�n�>.��>�#5>�+����>�Q�Lɽv�+?�mG?�G�>�1,�e0X��1о���ӡ���ފ=�~
��1,>�2$=���@%�y�r>���=�E��I?��<#a�3�9>�f=('-��>��&?16�=��t�9X�=S�V���R���>�d�fO��W��?%��Z6e��7��d����ꤽ.ƫ?;%�?��?}<�<�&��W�x?��b?��>���>+츾� ��㟾x���q����h7�+Mh=��>ˁE>&Oƾ	2������4����uK���_?a��>z'?��-?\:|>
��>ش����)���þV��Z���1�ru5���E��D����{O'� ��<�	޾ᕚ��گ>�a�b�y>HA?n�)>�>Z]>Z5=kO�>��$>q7?ow�>2��>~�>t�=�ὲ-��7�@?��ž���q�߾)1��@�?�6k?J��>�"�4���@�^�+?Ƣ�?���?W	>�z�J)�oC�>t?��-�{�T>?�<�i����>���-Q�kA���X>Þ�=b�=�%W�g2�`�j�?֩&?���(����D��橾&,>�E�?n�<?���TM�/|�C�]���F��q�;�q�����|!��@x�Ѓ���\y��v�;��U<�8 ?/ω?�-�m�����v�
2U��>���>���>�>�L�>����6��=]���!�aP����>e�u?�y�>�I?G�;?�sP?�kL?(Ɏ>	d�>�;���D�>fH�;��>0��>��9?3�-?_,0?�z?�m+?e+c>Hg��� ���ؾ�?��?�:?[?z�?х���ý�2��xh�D�y����� �=���<�ؽ��t���T=JT>b�?�n����I��"�pN ��9&?���>9�?��i���>Y]~>���>���>�����k�����*>�6\?Qv���0<�p;>�/�=ˉ=��F�N�X>��:��J=T��Sz��RJ2��LI<�]�=h7G�.����'=�+)=Aq�=']�>S�?ì�>�d�>�+���� �����=�Y>�3S>� >�Gپ{���&��o�g��Sy>�q�?�v�?��f=K�=���=���Ih�����P���#�<��?9M#?qST?ؐ�?6�=?�]#?��>�'��G���]���
����?!�*?�z�>���dLž�g��1�1��X?��?�y^� ����*�5c����ཨC>GJ,��=��%���C�g}:���������?��?5�%�Ea6���������W�;?�i�>4ݥ>�=�>A�)���i����aA>r�>�aQ?���>�P?ȗ{?z[?�'T>�8�aH��������4��8#>/�??I��?@�?�x?� �>\>�3*�M�߾����~��ע���肾��Q=9Y>s��>H��>�B�>���=cfǽ�����,?�G��=�`d>]�>��>���>5.w>�<��G?<��>6\������夾]���x�<���u?��?��+?�E=�w���E�3���J�>bj�?���?6**?ܱS�:��=yּZֶ���q�� �>�Թ>�<�>e
�=EF=��>Y��>��>��\�|p8�\�M���?�F?:�=��ſТq��q��闾��^<�Ԓ�6�d�
F��:a[���=񖘾���F���}�[�������������Ŝ�^�{�A��>���=���=j�=ӿ�<6�ɼe�<D�J=a3�<u�=)�p��Uq<6?9���Ȼ����Y�N5_<�I=�����ԾX́?H6W?�d.?��9?='�>=¸=J/K�9�N>|F�����>�Y>呅<�Ͼ`���G���K��ձԾ9�T�^��>���Z> �̽{>W�>Ũ�=1�<?�=h:l=s��<= E���o=�Ϸ=�1#>'�=6�>�4�=+�>�6w?���b����3Q��Z�,�:?B:�>�q�=�~ƾ<@?g�>>�2��՗���c�-?���?~U�?��?�qi��b�>H���؎��f�=�E82>���=��2�ͤ�>��J>����J�������3�?��@��??ዿ��Ͽ�`/>�E>
��=+�T�6�Jfo�@%L�ƯG��3$?�_7���Ӿ`b�> I�=�QҾ�٭��O�=�	&>7R�<��6�cV���=�y�)�X=��r=��>��G>ټ=�5��%��=Hԁ=��=�f]>��3���7�j�V��[=�]�=Ny_>~�=>g��>�?Gc0?sUd?�4�>n�!Ͼ�9���G�>�0�=�?�>��=�{B>��>|�7?��D?!�K?5��>���=�>��>�,�ȳm��k�nΧ����<���?HΆ?�Ѹ>/vQ<��A�ܞ�b>�I%Ž�s?DQ1?�k?��>Z����/R&�a�.��j��78z�*=1�r�3�U������o�[��Y��=w�>���>N�>�By>��9>��N>P2�>R�>p~�<���=�V��� �<ꋕ���=J���F��<��ż#H���g1��,�����E�;X�;N�]<���;e~;=έ?��G>#�?<�>B����v^>ʅ���=��l�=C���T�Ⱥ��Yς��~>���=0ؠ>���>��)�:������>[v߼�.�>:,�?{?�v>(�(��iϾ�ݢ��E3�onT�
��4�B>��꾁`>������gw�A�`��>ڸ�>��>e�l>��+�?��By=���V5����>󎌾T�}���q��8������Di�sɺ'�D?�7�����=�~?b�I?{�?܊�>s`���ؾ�0>=P��X�=��4�p�v����?��&?���>���"�D��H̾7���޷>�@I�.�O���V�0�n��.ͷ�7��>������оj$3��g��������B��Lr�]��>%�O?��?O:b��W��HUO����x(���q?�|g?4�>�J?�@?�%��z�r���v�=�n?ȳ�?Q=�?w>׬�=����>C�	?��?���?�s?2�C�kA�>!m�;^�!>���
P�=��	>>:�=q��=y=?�c?f�?�U��4�	����^K𾝏^��
=f��=��>�>�r>�#�==OV=��=�pW>b�>��>��j>xi�>�چ>���9�׾
y'?�y=>�>�H?�D�>G���j�@\*=J,��X;��"���������>�b0=6�=�F����>W󻿢��?E;>]���x$?�w��
I�%�5>->|ᆽm��>v��>�&>��>��[>��P>A��>ӊ�=�|���~>'��� ��i>�EK�}�� ��>�ϝ��U�J����4�����i���sk�)v�c�9�/�y=���?q����i�"��F���?�~�>,E2?�C���G��ș�=y��>Vv�>#(�埗��э���߾��?��?t�b>_�>��W?��?�;1��m2��tZ�4�u��$A���d�'�`��捿������
����i�_?�x?�tA?�E�<�z>��?\�%�D������>�6/��d;��"==�i�>�6�`�NcӾ�þ���åE>�Lo?��?�G?#TV����>�0?ϟ(?l�n?�0?c�7?�����/?~D>�q?�?<=8?_$1?A?q,E>d»=�֚�߮Y<q헽� ��K�׽���M1����>=��=��ӻ���ø�<���<���Pq*��\�;�Aͼ���<)k2=�^�=���=;�>R�]?�i�>��>&�7?I�ME8��4����.?�@:=���&@�����$?���>[�j?�ԫ?�KZ?�Cd>_FB�4BC���>w �>_�%>�f\>% �>߾��F���=�r>�G>�V�=	|J�[\���	��j���O�<>�&�>��v>�ʚ�4�%>~ޭ�.w��zh>��C�H��3[Q���H�4`,�G}���>ĆJ?�?U��=^i�ʌ��e�� *?��;?=N?i	|?~M}=��վ��7�M�G��(����>}.�<���ǲ��X�����<� �< 2>M��]����">����
�*;j��hA�_ľ84�=�$�L�󺅼��ؾ`����=P�C>���������O�L?�����2���Z"�7���Co\>��>o2�>5�Ӽ���[C=��`̾1��=Y
�>ἐ>
H��}�=�K�\�	�XT>��Z?���?I�~?d@���K���|�� ��%�ohϽe��>�M ?�F4?�y�<1)�>8���$� }^�i�0���>p�>��\(W���U�Q�������>�_?W�T>e�>�_J?��?!��?"8?R�?T)�>�-�𖺾�%?ڰ�?c�=wϽ��M�rr9�J��{�>�2,?3�>�Hΐ>|?�� ?��$?�hS?�!?�>t�'-@��S�>w�>:�V������b>7E?( �>&X?U�?wC>��3������~�����=�O!>zf2?��"?�T?t�>>��>
�����=ܙ�>l	c?�/�?�o?���=x�?�,2>%��>Ζ=���>���>�?�TO?��s?��J?o��>���<�5���@��7:s�v�O�%�;�dH<G�y=����5t�nS�\��<���;� ��6d������D��𐼥g�;ί�>fl>򑓾��$>����������Q>�I�7��
#��gh1���=~�n>T��>ٱ�>��#�Ng�=�	�>�N�>w��H{)?�m
?��?	k2�M	`�(|߾��W�ۯ>>E?���=��l�w����&x��q�=�cm?�Z?��Q�Z�����b?��]?�f��=�7�þͷb�a�龫�O?��
?��G�W�>l�~?�q?��>��e�!7n�����Cb���j�Uζ=to�>�W���d�g=�>��7?4L�>��b>1�=�q۾%�w�n��\?��?� �?t��?�+*>��n��3࿞����:���a?���>V(����$?���drѾ�瑾y���2��KX��4M��|I���.���y�R ��U��=xQ?�iu?spt?�zZ?����
�c���a�&P��#�U��)������G��gC�5�@�M�k����y�:���ZV^=)���M�(��~�?�VO?�̽�?󙯾�����ھ���>z7��d� �z8�=�T ��݊<�i���e�آ��>ɔ���?c��>�J?x�2?Q�E�3�TK�Y^>�����s�=R�>��V>3N�>��<|��jý�������L����>�Y}?�ak?��?h�+:�☿c��l=<�����q�<U>i��>[ɾt[�C��2�B��-Q����H���`��s��;LN+?c^�=&B�>�[�?u[
?�F�۾X���%�	�82�=��>��?���><->��q��j��N�>���?.|'?�>��ܽqb.�ى����I�ز4??�?�C�>!�9>�i�S݀�Fј�D���Mg3���O>��Z?����8���� >�j?���	h{=L�&>�z�>�'��'�r&&��'�>�.
?/@=��>�f�-D
�D��������(?u�>蔾5���)0>��?@��>���>�3�?�U�>��˾��>�w�>�kr?��A?f�X?ҧ�>7ʼ�6T��d齕[���=1y�>B�}>�D=o>E>X����<Y���h���>�C��0J��pWZ���N���8=M��<U��>�Ὲ;G�ɼ��F�V7��+�$�Y���-�EM��H��]iӾ���k��Co��?½wn8��� "n��B6��J�?��?�׼������q���D�U���?8X��$��=;`��s+���p��7���c���NB������l��pY���%?����l�v5��n��?��)?$�n?�a����Y73��oZ>k�"=�Z2=�g �i���Z�ƿ�`����b?��>;m�o���{��>d��>��>�;z><��i=��p����>�+#?�??�ד��Ŀꈺ��)=E�?��@ �A?7�#���Ɠ�=,4 ?t�?WwB>G�A��I����rb�>⾛?.*�?��
=0�Y�Cf��1�[?6z�=�=)���`�-��=��=�.�<����KB>vn�>�G>�i�>��ý�`C>s��>6*��&�2���n�{1=0ƚ>/�ɼ�Z�*Մ?{\��f�m�/��T��%V>��T?7+�>/9�=��,?7H�(}Ͽ�\��*a?�0�?Ԧ�?��(?aۿ��ؚ>��ܾx�M?KD6?���>�d&�!�t����=�4����:��'V����=��>n�>ʃ,�ˋ�&�O��G��n��=�v�MǿM�"�h��ˉ;�q���{��+Y�q�z���/�C��Sb�Y]� ��=~eu=�&�>��>!�f>n>�F]?ޭs?���>9Z�=<���~��~~��\BT=�)������y�4_!��j��{�վ8J޾nB��w��y�՟¾�_T�Ʊ7=aRW�bƔ���v�D��v���`G?�}�O��]C�}�>i,��+�;��=�=�������i��T��6�? g!?&!z���*�9"�n
4�B?;���W?�K�=���֙��eU>I��
��\'�>��>.09�U��|�J�\/?�?�7��e%N��Q>�<���= �+?C		?�kE=F�m>�j6?��X��=c�n>�P�>>bQ�>�W=W�����P��w?l$O?>V-����� ��>����;�����<�	>M�B�.��R>ݼȼ[(������=g���5>��V?��>d)�&��w���X�
�Q=Z�v?��?lU�>�j?��B?���<�V�T����$d=jwV?t�i?~�>����h�ϾB6����5?�le?��J>a�j�D���.��Q��@?�o?�m?	�����}��.��7:��7?��u?'�Z������5U���>�>�l�>�5�痻>��;?X	�n��u׿�l=6�(ŝ?� @�a�?�G =�z����=_�?���>�W���ξn�������h=�4?v'��=Ws��$�J�<���:?��?S8?�������=�䒾nլ?�K�?����-�<���ęk��� ��u=�H�=pC�U%��?�v7���ȾK|����ح��/�>,@�MͽSy�>p�7��Y��Ͽ񨆿�о�Uy���?zx�>:�˽�4��[ci�{Mr�3D��qD�����w]>$ (=�����p�&�����i�:]=K-?>����d)>x�M=��U��?��<���փ>P��>2�>NɽT �v�?$�#��������w��?�ѣ?�#?�8�>GX��GC=�¾O�>H�?_�Q?�}a?J]��������g?�먾�E�z������א>�0?�O5>����<�<m>i�?��=�a<��yÿ�أ�%@5�n�?n��?>b��R+?���?��>��;����4���A�o!��"�S?e�lσ���k�Ȯ\��_�#�G?s�]?콓��_?3�a���p�k�-���ƽUۡ>��0��b\�?N��u��>We�����<y�O��?*^�?%�?c��#�(4%?��>����7Ǿ��<���>�)�>R)N>�=_�ܰu>/���:��e	>��?�~�?�j?ᕏ����tR>��}?
)�>�?�[�=�_�>9l�=���6+�r#>�%�=M�>�̜?��M??�>1��=@�8��/��XF�YFR�8�p�C���>_�a?�xL??ab>����:2��!���ͽ�e1���?v@��k,�^�߽�5>��=>E>��D�m�Ҿ*!?fP���п3T��QmҽH:?ZP�>���>J(۾s�>N=I]?�[�>H�Nm���d���Ų����?���?a?�GӾ����<�=$�>�uc>�lm��������0>߫;?�-������p,r���f>l?�?B�@��?S�]��	?��nN���[~���7����=A�7?����z>��>S�=�lv�������s���>?D�?7x�?!��>w�l??zo�H�B��@1=�@�>�k?Z{?|�y�P
�ʹB>4�?/������>T��f?��
@�r@˕^?"ꢿ���������o��}��=���<��=�rJ�c�=�H�<,��Hݼ��3��ӝ>Qn>�9�>�t>�W>xd>��x�.��jg���͂�J�:��� ��|�@��m޾������_��`���.�q����+�ν��p�M,R�n�����=wT?tO?�o?٦�>H���4�%>����Y�(=�V��_=�t�>��.?��N?�*?o��=q����c�t��2����߂�<��>�?O>p�>%�>l԰>@p�:PYB> =9>E�>���=�"=���v��<o�A>�©>��>��>��T>%U�=vD���'���a�1�Y�8W�C2�?�Ė���H�Ӏ�@즾bmf��y�='A?��%>�����Jɿ���ʕE?�Ѧ���[B���m>�4?�E?� Q>�R��U|,�� >uK�x]O��e>PQo�y��&�5�s��=ڽ?C?�>s:>�3��*��6Y��1n�O��>�9?V˴�Ȩ��j�a�����ܾ��>���>w4=� "�eؑ�Qo���}��&�=<?gT�>��	�~ վ�0���Os���3>c3>b�Ͻ{6>��>S2�<�+M���k�B�=�2>���>h?��&>�h=� �>�Q���K��P�>�+J><�4>�l<?� ?�r��'���h[��d��g�>���>�Fh>tz�=��L��=8��>$j>�pѼn��������8�R>�+{�H�f�OpN�fB]=�䓽�E�=\Ђ=t��1�r�k=3h~?AP��;ʈ���꾺ܻ��=D?Ln?(�=�`-<�;"��禿�巾e��?~�@M�?��	�ןV��N?�*�?2`��P��=�`�>�)�>�U;�YO�\?MƽB���G�	��$���?���?��0�%㋿�Al���>�P%?�;Ҿ���>����<���>����p�mB=ٿ�>QE?_���r��:� 
?m�?.��Tx��*�ȿn?v����>���?���?��l��͙�Y�<����>e4�?%6T?�g>P�Ӿ�W����>�'@?��T?�r�>%����2�oD?���?f�?`�A>?.�?�Cv?���>��p���*�����!J����~=k�����>�'>G��G�Xj��5��{k�]���Y>1�7=�Ѱ>��ؽ9I����=�Ό����0��ǭ�>�Yk>\�E>�>�?�>��>�j!=�I���,��i6��PJ?���?�]�+fd��1���aQ=G�D�I�?"�8?¯H<T�Ծ���>��N?K}�?jBW?�<�>����.��0⿿̱���n=Om>�?��>�g�uqx>���.B�X��>�!u>yz<�O�'"s�����i�>��?�_�>��=�� ?͙#?j>�)�>JZE�{6����E����>���>�D?��~?��?�ȹ�Z3����f硿e�[��DN> �x?IT?cƕ>H�������E�I�I��(��?�ug?�F�?�1�?N�??��A?�%f>͕�T�׾b��G�>�W.?�۾��5�$���H�<h?N!�>G�?F!��v�H�;�+?�9��� >9?��v?��>�f4�A5g����oQϽr�ռ��<"Xr>�&�E�0>T��aܽ�
�=��V>�ޑ�)�="���H&v>����]�>	�<��"=L�
=K&&?ȍ�=�����[�=�XT���8����>�����G���̊?��t�ܲ=������U���F���ۈ?���?Y�?�*�=�N��<?r?�Ȓ?3�?f)�>"=��0־NҾe���8�J ,������g>;Q �J:��k���g�����p��J�%�M��3?�'�>��!?s�?��K>XU�>�Qپ1$,�������a�I��R8��<�@aN��k�C���!+˽�� =H�׾◷�7v>���<�@�>u ?�,@=A�>�%?,B>£<>�9�=�>N"p>;g�>�u1>���μK*���F?0��1,&� �s豾�	?�t~?<?��D��т��G�lz'?�+�?�כ?�i�=Y@~��� �'��>��?�S��J�>')#=��_J�>��	|�ꅊ�珼Dx>).> �P�/7=�b��N�!?�z�>����ξ�`�9����o=9O�?� )?��)���Q�~�o�շW��S�i	�N=h��f����$��p�x돿B^��`!��M�(�ҏ*=��*?p�?W������$k�e?�9Bf>x��>z�>:پ>[I>��	�L�1�\ ^��G'�����=_�>^Y{?���>U�G?�I6?3P?}�H?_{�>�۱>�A���*�>��<<��>��>�0?7�1?�U,? �?
#%?iM>j��u���?Iھ9�?Zg?R5?�< ?�?ޭ���0߽�l𼆖�<�i��
2Q����< ә���
��e���Y=�̈́>�?��A���,��+پd�w><�5?�G�>�+�>�g�������=�2�>n ?�ɋ>�q߾D�v�3����>Eq?	O#�s<��>�v�=8d�=�D=�=>L;���=]Ͻ���hy���.>@+=�:��۩O��b�=��=c\=�[�>A%R?�� ?��l>7�_���ﾩ_<�H�����>鴲>I~�<"v(��z��՜�;�t��>�S�?h�?F�=�$F=���<@�����־�����C����%��?��@?@0r?��?�ER?`�!?��=�@�����-���H��=?�b*?��v>��?7¾����P�h#?SG? �b�ۈҽň(��掾����i>�+�Y�u�.���
�B�X��<���
�l�?z��?nVY���L�	p��V掿Vߥ�e�!?��>1B�>Đ�>^��u��'��EL>u��>�\?���>�6P?��{?r[?ΠT>V8�Om���%�����f!>6�>?B��?%�?vx?Yn�>�>W�+�\��s�����7���EЂ�muL=ޏY>$7�>��>͙�>Ƴ�=7�Ž���v=����=��e>�p�>t��>���>��u>��<��G?d��>�K��ri��㤾Hك�s;���u?ח�?H�+?�=0.�R�E�����L�>�q�?�۫?�*?A,T��h�=3-Ӽ0���`q�|X�>�̹>�k�>	�=56E=''>���>in�>69�qd��c8�zO���?��E?q��=e�ſ�q�W-q��藾 MX<uX����d�}򓽅[�� �=����9q�ө�Z�[�}x��8�������K�����{����>5��=��=yM�=��<��˼�\�<�`L=�ѐ<��=��n���l<:�0׻����cn
�Ϊa<�OJ=$���-pʾ��|?�H?-+?ȣC?��z>��>y0���>�脽�l?�)S>OK�^;���9�Ű��:~��8پ��׾
�c�*���Ȗ>B�H� [>� 4>>�=�G�<���=��p=�5�=�R���2=��=���=tϭ=5�=�#>[q>�2w?X���a����<Q�y罄�:?�=�>o��=πƾ�@?�>>.0�������`��+?���?�R�?��?�i��o�>���ߎ��k�=Kt���`2>���=b�2�4��>��J>���rK��+��2�?�@�??�㋿(�Ͽ/4/>eW>�I�=8�N�a�,���L��@9�9�G�ͽ?w4�>�ξ���>ݡ=�Ǿ�T���Z�=m�7>vF/<��;��}Z���c=�}��N=ː�=6�s>�4>=c�=�첽��=�J^=Sи=��X>�;�0���E�C�=Ff�=HNa>��	>���>��?mY0?NVd?�*�>Sn��Ͼ�%��Y�>=�=Q(�>_d�=�QB>���>@�7?ߺD?��K?�p�>wf�=���>��>Ύ,���m��N徟Ƨ�ܨ�<��?	Ɔ?}¸>&�Q<F�A�3��rc>�IŽ~f?�L1?�g?B�>����俩�$��������T��vV<t񎾆��=A�
��CU���?��(]<�i�>��>��>a��>��M>x:>��>�>�z��)	;�Խ��B�� <I�>�G;S���ㅼ���r�=����B[	�^>½�D�=�Fa=�G��~i=:I?���>lu�>�ȁ>�̌��	�>ld��`����<��ݾ���*���耿0F�;EὋb�>��>���=������>3`��׻> 7�?�sd?�PO>�.���X��h���T{�����Al=���>X�Ⱦ]�6�����3{����8��>;Ύ>\�>p�l>� ,��?�G y=���K_5����>�q��VV�x�q!q�9����.i��7ߺ��D?>���r�=l~?�I?�܏?��>������ؾOM0>�=���=t��q������?�'?��>�����D�C�̾,Ⱦ����>��J���P�s/���w0��J����f�>�
��7�Ͼ�i3���������B�}�n���>O?�
�?�rb�sF����N�Ҩ������?�Hg?�Ƞ>�?.�?��������5��=�o?�t�?A�?��	>�4>���WL�>�l?$Θ?�$�?�)d?\�s�?H���K�K>�/�W;�>앧=
��:�����>r�?a\/?��y���uGؾKm��*,�4'>b�6��T8>u�>�U>(�2>p��=��[>6p=��R>ќ�=<�>V�?<��>Su��sF��7p,?zӽ>Kz�>�a4?g�C>P�_�<f>�\�><Ib��LA��׏�Ϧ{�)�O��S<B�U�>=ā�>@9¿���?4��>��	��,?4�(��o>�g>Jk�>ې�<�>0��>�*/>���>UD>�${>}��>c�=M���aT>��	����4�o�H�����#�f>4���U#-�e��d˽��C�m)��E-	�Bf�9x����9�'��={��?��/���e�T�#�>dŽ�>
?��>��$?�O����ɽia>���>� >°�ꕿ�.��A����?���?Mk>V�>��?7�D?|=�A:��x�[����"���&�4�m�]���=n���$��3���O?���?c8j?���=�B>��?RV
��k��V�>�O/�;�C�H�u����>�����f�3j-���� �+�ɔ�=��?�ۄ?K�;?�b,��1W�Zq#>��8?v0?��s?+�1?jH:?lq��v#?w>.>�H?+Q?/15?T�-?�;?h�.>5��=��)���=�m�� ����ӽWǽ;�ӼG�C={#j=��T;�}�;��=)�<���*�Ӽ�;
����<G=(^�=2��=���>|lm?s�?g,�>@�??��F��F�^]-?J;=vf���;�"��������=�n?��?Gm?s_>W�@��y�q#�=��>�$P>��>�U�>��D��U9��5�=��%>bz�=%­=8K��C蜾��kA��u�<Kv>c?��>|���5�a>�@X��z��ɷ�>^
��<��1�"��4��}�
����>$Y.?͖?��<E0��_�Լ-N����>��?�??2��?%&>�k���O�B�>��=�@��>���ѾF٩��Ȟ��H�$,��w>b����(ʾ��>Q��N�d����D�6����5=C��-���,����(զ���=s3>�=ݾ�d%��吿�$���@?���=p(��Ky#�);�p�=���>��>��:��=�8����YL>��>a�K>D�:�W��[?^�.�4��x>�>?fXT?li}?�����|n��1��;���*����
����>�}�>���>D�W>��3="@���~�>�d��D�̄�>��>��z�M��g�1Eܾ�V����>.k�>
�S>s��>�?G?	?[�t?mf4?���>�č>�( ��Ҿ6�?<�m?���<*��qX��Y5�F�$��
�>��)??Cͽpt�=�5?P?��0?aJE?&m�>��=����r@���>�^j>��o�@������>�%E?��>T�|?�F?���=ӗ�+Z������6�f>��-?[�/?�0?�Q�>E� ?Z߲��_=۠ ?��k?�_�?�m?�͎=͉�>�F�>>��>i>�?Ik�>�6�>L�f?1�h?��;?�8
?dh<H��̧<� U��~cֽ��̽�n6��T\<a��<�Bb=~�i<��C=��>�\=-X���=���6�=UȎ=�M�>��s>���#0>8�ľ�/��rA>˝��@�������P:�r#�=KS�>0�?7>�A#���=P�>O��>'���(?�?�?$�.;�sb�?�ھ3IK�M�>{�A?�6�=L�l��l����u�Q�g=	�m?�^?�V������b?��]?�O�=��þ��b��V�J�O?5�
?��G����>^�~?y�q?���>�e�0n����$Eb��k���=_�>�m�6e��X�>�7?�[�>�9c>��=�E۾Ŀw�JQ���?��?��?3�?�*>q�n�j1��kɾ�Ț���??�f����K?N9;,��Ꙉ�c�k�����n�SB��m��o˾�������\%����>�"?Ja?��h?/�T?(��7N���W��ea���w�}�0�
���h��o�ґH����!�#���ԾA6��z=�=�
q���A��$�?�{*?�q �m(�>)����q�þ�N>N������{7�=Ъz���'=��w=��S�_&�����!9?S>�>\��>W�;?~z[�D!?���0�W:4�7d���M1>98�>�}�>���> ��;�R(�����tǾ�>���佢��>V�a?P,f?���?�=�|X8�ut����E��T<sኾc�>\��=��D>)b���y��G^'���9�Fi���ݾ�ʉ�A���L���]"?$�}>�G�>���?�?���4���A�M�5��6I0>s3�>)�j?���>��>�C����h��>n?��>?8�>򰅾�l"����6�u0�>+`�>?��>[�n>�@�p�_�-~��Վ��m9��@�='Nh?�����d�c��>K9Q?(O���;D)�>(oP�#���*���?����=/�?c$�=j7S>a��5(�5|��h��g&?�R?.���z/��>�#?;��>��>rx?���>�o���c
�Ir?H[S? �E?��=?6K�>z=x��������k5=h�x>F�:>P�R=Iރ=���<�/'�[.�=�k�=�j�;!�ý��;��"����;/G�:5�3>��ڿ��M����\����v�
��s��e����g�t��޾'¾����{���NZ<r��T�m���n�գZ�ñ�?\4�?6��b����{v�)&۾� �>�d'��?�<hþo�o�[i�����©�oN+��M��w��ҁ�YC'?�{�����)<��>�ľl�?l�!?�Uz?����25�` :�	�=�v��hx��3Ծ���X�Ͽ���VZ?���>�*ھ.��Y��>��S>��f>6:\>Y���+���Hw���>k� ?�	�>�\w��ɿ�,���6� ��?��@{'B?f�(���Y��=M��>g?.6>�@5�ak�Y����>�۝?+�?��<="W�sr��?�g?W�4<.jD�P����6�=�o�=_�%=v/��V.>}.�>���9X9�N ս@R4>�#�>�%���G�C�e �<=�X>aQϽ�s��5Մ?*{\��f���/��T��U>��T? +�>Q:�=��,?X7H�`}Ͽ�\��*a?�0�?���?#�(?;ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�܅�=p6�������&V�o��=X��>c�>,�����O��I��`��=��=��!}k���U�~����踾�򼓢ξ*"�c�������~�n�#�?7��>ٜ�>�|�>N��>b҂>V?��m?��x>%� ��԰��{�6;�N�<os��C�������l���j���̾JW�\v��n��¾�S�Kv?�!�a=�tU�|я�M�+�Kf_�� ;��m*?�3>��Ѿ��T���˼)�Ҿ�x��$��;��ٽ� о�"0�4�m���?��>?X�CGQ�5��J�&�
ݛ��P?A����]�Ι����=��ͻ�7B<�(�>>��=Y�۾N�5�-�^��Z ?�g?I'���v��������I��XE>��'?qC?���?�>&?I�������v>:
(>���><�>fc������)��A?P�N?�彔۠���N>�9�D)Z=�L=�>��<��Q�3�>���7r��"�m�o~��m=�W?*��>
�)�:�bY���3 ���C=�x?Ԏ?�m�>�$k?��B?=|�<����S�w�
��Fy=!W?��h?��>S8�4ϾG@���5?��e?�N>]Dh�S`�
d/��H��]?�6n?�Q?����Md}�:A��E@���6?��v?�r^�ps�����_�V�[=�>�[�>���>��9��k�>�>?�#��G������oY4�Þ?��@���?u�;<��s��=�;?t\�>&�O��>ƾ�z������A�q=�"�>���cev����R,�_�8?ؠ�?���>-�������O9>����R��?d��?�v�^h>����7پWr�= �=ۜ�����R�۾�fw�� �H�Ѿ`B|���>?�>Si@Mٮ�O#p>뽺���⿲RȿX�������ռC!U?j>;J��P* ��nl�ӧ���e�FRE�u?���@>�9>��� ��0�p�� *��E=}�>�)��6t>�E>�����`��rv(>շ�>���>���=Ly�:�ʾ�ё?��;缾�G���s��]p?�[�?�u?�"�>�HG>:{�F�F=�X�=��K?�J�?��_?Ñ�>�q�5s��j?_��U`�4�SHE��U>�"3?�B�>5�-���|=�>͉�>f>�#/�X�Ŀ�ٶ�������?���?p꾃��>y��?�s+?ii��7���[����*�FQ+��<A?�2>
����!�H0=��Ғ��
?Q~0?�z�5.�}�_?�wa��p��-�H�Žfǡ>�!0�e\�D����C �S@e�����_y��?�V�?���?����#�%?Fگ>�_����ƾ��<�\�>�M�>e�M>��^��u>QB��:�o>|��?h�?�P?�������o�>+�}?ɶ>��?���=�>�o�=��1�$���">�|�=��@�|p?=�M?��>��=��9��/��F�mQR�����C��ۇ>��a?�nL?�?b>5V��<5��/!��2ͽ]0�~�⼖�?�\4)�3�޽0g3> =>��>��C��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>@�Խ����\�����7>1�B?Y��D��u�o�y�>���?
�@�ծ?ji��	?��dP���`~�t����6����=W�7?}0�}�z>x��>��=�nv�仪�t�s�c��>�B�?W{�?`��>��l?��o�/�B�h�1=�M�>��k?�s?_�n�L���B>��?��������K�if? �
@su@&�^?���ֿi4��#*پ��|�3U�=3���g=2��<��K<7_��7�=�ȿ=k�R>�E�>�~�>:}c>h�=>#m,>��=w���I�#�J���᫈��B��[��(>��Ss��W�3⭾����]����ܾg]>]��d��=OF�� �����=��S?�P?��n?G��>���>q���>=-��UG=g�>b[3?��M?Bw(?�˃=6b����e��-��Τ�Z������>l>>"�>x�>]�>�1\<�A>!�B>}�w>#�=QM=%|P<�
/=�"N>H�>�[�>:�>�VH>�)>�T���q����R�Wb��O&�� �?/b��g�T�r���+���ݲ�ʽ�=_E6?���=!ϐ�,�ο����{f@?�y�q���.�k��=��3?^�I?��5>�T��n�����=:�O�� ���e>�
�/��7�ڦF>�x? z=�a>�;��!/��cm����u��>Rx&?�Aþk?���񆿩�c�Ef���>�-?0X��JM��L���u�RJT��>�O?G?g�k�q+��̾&ߺ�Q=��0>B[>"z�=;&L>M�ڽ��}�(��j9��P�<T�>�?��>Ȝ�=>��>&���F�<�2��>��m>6�>�5?*)*?���ü�������?�z>���>�Ι>�g=��<��y�=�N�>m>�M���"ν����Q�\1R>����a�����0=k�m���=-�i=���_�\�,3=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿf`�>�s�|Y������u��j#= �>�7H?�W��o�O��>�7r
?�?�X�ʨ��2�ȿ�|v�l��>��?���?2�m�2@��@�"��>��?�jY?�xi>�c۾\XZ����>��@?3R?��>�5��u'���?�޶?k��?e�>2��?��z?@??K>/�8�����9����{
>R^u>���>���<5#�'���,���¨��o�d��;�� ��>pc�<�>���<0ᚾ�=�j�CI��%�����>��]=_~�=��>{?[3�>J�>Q!@>�mĽ胾��ɾ��K?Ѡ�?���n��Y�<��=qK^��:?}84?U�Z�Cо��>8�\?˱�?��Z?�K�>.��r(��hԿ�D�����<��J>y~�>���>1����K>�OԾ�E���>&�>�ꦼIOھ樂�8d��VQ�>Q}!?��>8�={� ?�#?{m>��>�,D��&|F�=��>�0�>��?@�~?u�?Di���R4�����Kl���[���L>�Uy?�&?���>R���9����l%���Z�L���S*�?XMg?�4�n?�و?�t??�??�*f>�z���ؾ�����~>e&�>��[<�oD�P�6���{=�$?�1)?/[�>t�8��M����d]��<�վ0��>�g?�hE?���h�����ܾ���;;Җ=�=�=���=f������>YG�>�>���=�^����'��{	��Ҿv">���>>�=H\������k�=_,?9c3��v��8?�=�s�p]D��9�>�DL>^����^?��=��z�	 ��q��6�T��ȍ? e�?�1�?j9���Rh�D�<?��?�8?;;�>4x��i߾L�ᾡ�u�hv����N�>��>�rB��&s���[��!���?�ƽs+ƽX��>x�>��&?��>pTg>y>�ƾ��t+׾8�Ӿ�dO��
;M��7���"�[1ԾDDR���=�+���:���ɐ>O6���>j<#?��G>LKW>	z�>�d>�r�>t0
>���>�H�>�w�=�s}>��>�A�=��߽�2R?Lg����'�D������A?��d?CA�>�+h�(���י�i!?�[�?�F�?��w>JAh�x+���?П�>Ъ�Y�
?�#A=�Y�H�<tp���
������KČ>�0ٽΌ:��M�]�e��
?:�?뾨���̾\Gӽ�����=gσ?)+?�$�z^Q��p��U\�u2O�vJ��۾R��Щ�Bm*�0�r�'���������%(���=�'?�]�?!��<�,q��r-l��A���W>H��>8��>ͭ�>��K>s����2��4[��v,�^�����>�r?��>R!E?:<?��S?U�U?��>�%�>$����>�V���R�>�+�>�<?�,?��/?�?V�&?g>����j���26ᾰ��>/6?ȿ?�%?��	?"[���/���ռ�;��c���G��(=(�=�ߍ������4<��[>��?߻�@�6������h>E�5?�{�>��>[ʒ���j�,=.�>�?%Q�>���	(o��J	�-�>�K}?~��I�=3'>ud�=�����S��|r�=Q�⼹Ȍ=�mļF.��KU<]�=O��=S:׺(�����v�<p�<mt�>F�?|��>p>�>�O��ɩ �ݬ�c��=-'Y>�
S>�>�1پ�|��$����g�\y>&u�?Mx�?1jf=��=Ҕ�=l��?����/�����<\�?�M#?�TT?k��?��=?�f#?��>)��I���Y���(��,�?�^?/�>Lhپ\���U��=����"?v��>ـ@�.K۾�bG������;���"=�F��_�~�|���&�]�(d�=i��U����?���?uC���A�!�����l���HD?���>�/�>���>�/�h���[" �]�=�?x�S?Xz�>dEL?��w?��Z?E�B>4�;� �������<�)>�m2?���?)��?v�w?[�>�Z>�'����ͩ��dI����6��z�=��v>~A�>���>��>o��=�����½(�=��?�=^�>�9�>�>��>�_>��<�\K?r��>kI����	�ϙ��ߜ�Cz�mz?�z�?a�/?#Y�;M����������Ү>[��?p4�?�5? �����=Fs�<��ɾ�Ÿ��<�>�W�>/��>��R>��=���<2	�>�y�>���
�+�<	.��-�o�?\'E?��%>�ſ�)q�Ȉp�oC��ZhX<�n��=�d��k��{�[��=Ba��pY�੾��[��#������p�������|n{�V��>��=��=�Q�=��<{�Ǽ�?�<7EH=�֋<Y�=��k��y<�4�a���2���*���a<*�N=���߽˾h�|?��H?��+?�.B?J0u>^�> (@�,��>"��Y�?�NW>�b�m2��� B��ߨ��ʘ� �پϮվab�Ƕ���L>n�_���>L73>M�=tt<��=�X�=� �=jA��5*=���=��=$��=q��==�>E4>�6w?W�������4Q��Z罤�:?�8�>j{�=��ƾo@?�>>�2������xb��-?���?�T�?<�?Bti��d�>K���㎽�q�=G����=2>y��=y�2�T��>��J>���K��E����4�?��@��??�ዿТϿ9a/>>�o>��2��Z��ܼ��:sTT>~�!?�t9��D���$?�z�>@�=}�ؽ��J><&�>�>�6�=޴x�U/�=�dh��i��+=G��>l�B>A>x��%��=��,�-�>7Q�>��/K��8�=�V�=HX�=���=ߢ=#q?�?D?"f?fO�>� ��
���6��~��>�a�>�^?웇=�n�>�Ν>Y�'?i!@?�[?��>b�=�I�>�, ?F���₿e�$��Z��dӽ�ܗ?��?cm�>`ը����e�Ӿ��"���G�T�?J?!{-?���>��<῿{'��:.�x����8���=�q���Y����&[�g��Q�=婭>�~�>sF�> �{>>;>:JN>C��> v	>��<��=�ub����<m紼�Mt=b����T�<�翼�ƻ8��(�#�0�ʼ�Ś;j�<Q)�<���;���=��>�$>���>�z�=W��Zo/>s�����L�+Y�=�G��B��(d�=~��.��T6���B>��W>�����+����?�Z>�}?>�}�?|4u??�>q9���վ9M��rve��S�Q�=l�>w =��;�.e`���M�bҾ��>�X�>%�>�q>�%� 7���=?�۾�G-�r7�>򠾩�½��4��Mo�U���p��� 	v�����xL?Z/����|=���?��V?o��?a��>R����\���F>8h>�o��<x��C�g�Ľa-?�40?��> z�w�=���ھ-/���̣><M���O�{A���7�o�Y;���4;�>�f��?徴�(���w�g��ӷ@�$ؐ��a�>1C?���?/P�`x���S�pN��7N=��?��i?�ݠ>�q?O?dр<�aھ=6�ח>qn}?���?��?��2>QՄ>�L�g��>��&?�6�?�\�?˯@?yy��zu>a�C>�G�>�����͐>P��9�]���m>��?���>��?S�<�� �_
��ڷ��jｅs^=��+>���>��;>���>wr>��K>o�>�$�>��m>�6?2�>�.�>��'>`n�L��%�!?H�'>���>�f<?�-�>	����GX>�%>�� =���<y�>��>�ә=0�=s��=m�|>�y=��	?AsĿ͂�?��>�q�� ?�x�,/=Ɔ�>S�=>��3�qhr>]�>Ѡ&>��=> Q�=p��>c�>�A��>&(�����IN������0�N>��Ͼ�Z3�K- ������10�	k��c�^u�
%��7�J�X�����?1�*��6�Y��B:�=�?5EX>v7?*�t��{�]f�>G�?���>t:��򝏿��l������?'�?O>c>U�>��W?|�?�1�~3�LvZ�`�u�g'A��e���`�፿r��� �
�C����_?�x?'xA?�k�<�9z>���?��%��ԏ��,�>m/�*%;��V<=�)�>�$���`���Ӿ'�þ�7��FF>[�o?�%�?�Y?�PV�n�p�Lw'>9?��/?p�s?z�1?$@<?r��zf#?�l4>��?�?1�4?��.?=�
?��4>���=���5�=����ع��Reн�Ƚ~��l47=b�u=�:[��<��=���<��ټb�м�*���q�� �<j�3= �=U��=H�?��o??�??.>�?������1�!VQ<�p�?�}�>��!��o������	X�Ra?%�?Q�?���>�cR��5G��Q>g��>Xm�>~t&> �>���n�s��$&=0�=0O=[�B����=�/���a�0�w�MU�<[��}u�>)&�>�����>����d�B��>�+<�F举*au�	�G��,0�2���d�>��N?��?�6=�I�������a�~�&?�A?nM?x�v?�Nv=��� �9��?E�?�=�}��>	K<(��堿Go��aZA��o�Zo>����j��<>݈�b�Ⱦו���������F���)̾���= ��3�k�bM��,L>�K�>[}��Q%��_��������8?�h=�O��ݠ�����>[�>�v>e����2%�\q���>�&?�e�=�<�ڻ�HbD�S���>�C?�2b?֊�?���>jo�jD�e<�Uu�������,?/�>/?C�@>]N�=T�������^��B�_��>F��>�7��I��[�� ���%��`�>6(?oy>-�?��P?�L	?B�a?�+?L�	?�>�`���7���d?SG}?A5J=h~ڽ!�m�&�7�
�7��g�>C�0?��H�
��>}?~�!?<�.?�PT?ħ?t�>���8A��Þ>�o�>7'Y����$<�>C�I?�V�>E�T?��u?�m<>~�-�ճ����ƽEٚ=��=�X*?�R%?�%?w}�>ډ�>Z����=�2�>��b?0�?]�o?���=�?�;2>K��>xږ=��>���>�?1KO?¹s?��J?`7�>�ڐ<Bګ�Z>���u�<�C�Vz�;`A<G<z=-��ot�B/�A^�<��;/���*툼�@�X�C��
��lf�;�W�>�t>u���t�0>��ľ�&��`#A>�H����aǊ���:��v�=���>6?���>o#���=ڙ�>>#�>����,(?j�?��?�Z5;wub���ھlK�t��>U�A?�6�=P�l��w����u�;�f=L�m?rt^?BW�����Okc?ƸS?����0�Y׹�xm*�s��s�:?��?>.�E �>u�i?Z�{?T�?#�Y���h��J����\���\��,�=��>O}�Vb���>I!1?�T�>5��>��=3��t��1�����?��?g��?�:�?p�>Gkp�7ؿ|R쾷�!�c?���>q>��/�(?r�<���Jr�l`����|���秾�1���j���,1�t,S�6᡽L�	>�i?���?�u?��Z?S��܌`��h��#<K����gb�ˣI��J���G�љt�������C��R{=sR�wM�g�?�<9?�t���?�噾�0��L��?,�> k���Ş����=;���*�`+���*��� �x�m�a�?�	�>�>��*?M\^�}�;�O�+�2�8�C�׾04G> m�>(�>���>[ ����O�:������<(���ܽ;'~>N�`?e�W?vw?�T��0�-��;��wA1���y����aN><J9>z#�>j�Y��wA�9�*�a�4�{�k���������A�Y��=JB1?��s>�]�>zќ?8�?y���#���ِ���.��O�<u��>��p?�>�>��>Ң��x����>֑l?;6�>��>�L���� ��s{���Ƚ�]�>Ƙ�>��>Lmo>J$.��\��Z��,|��Š8����=+�h?{X����_�Q6�>D�Q?<T�9�@<}��>�vw��!�`k򾏿'��u>18?�@�=�i;>�qžL����z� ���Q,?��	?���1��@
k>m{'?�B�>S�>�?���>#�ľ�SM��z"?Άs?07H?��J?b�>���
ͽ����m��nV�<�X6>V��>�h=��=7K�tH���Sw����;kW=��� lI�Z���k=�����O��;>�^��]�+�i�"��\0��� �am�<�ֹ�����$����̾4���a���7�qH/�}��h���?_'�| ����?���?�e���#�&B��>k������P�>�R�;�=�����fVZ��\�����@��gG�|������l�'?Vn��p�ǿ򠡿=�۾8 ?UB ?��y?h� �"�D�8��>��<롼<y�Ռ����ο,Ϛ�c�^?���>���8ѣ����>��>��X>�3q>(ׇ�o������<��?�q-?�j�>��r�v�ɿ�������<���?;�@>=?g�M����G,>��>��?��{>�@z������]�"��>���?K
�?+�|=&T���߼��n?y={�+��A<x3�=g>8�X=�
1���V>�+�>&*�=��I���T>t@�>�[��C� �
у�Y����]>��۽v�-�3Մ?�z\�if�~�/��T���U>��T?+�>H;�=Y�,?J7H�I}Ͽ��\�	+a?�0�?��?��(?�ۿ��ؚ>i�ܾ��M?@D6?y��>~d&���t�t��=�1Ἐ�������&V����=���>��>��,������O�FP��f��=C���ƿ��$�@��B=�8�o[��X罭���-�T�g�� Co�F��h=���= �Q>u�>a)W>Z>@cW?��k?�I�>Rl>9�㽒f���ξ�~�e���������f�����Up��߾�	�#�������ɾ�U���%���T�)����,�l|e��1�wx#?2��=�U˾ڮF���=��cB��M,�U�ٽ'ʾ��"��4j����?�	-?�.��o�k��g��,<�e=/JS?'�9����L¾��>գ��}\=Fa�>O��=Xݾo�0��rU��?�!? ���*����a>b"��ѽE"?7��>��??aؾ�@s���=���=��>@�!?xqa>i?T�.�?#)2?�t�r���X>�Ϡ���w�D�\�Z>+R#��:8�8�k>������w�#��뉢��\���]?�Ig>d��7��~k��+0�<Y;���L?`�?��>�n?��,?�i�������C�x���=�=�N?�oD?U�>5�K��������:?;�s?Ba�=�_�%j�g[���!��@�>��?�@?MVC�\hp�,U��\5:��(?��v?�r^�`s�������V�9=�>�[�>���>��9��k�>8�>?a#��G������hY4�Þ?w�@~��?��;<�����=�;?9\�>=�O��>ƾz��i���G�q=y"�>����uev�����Q,�P�8?ʠ�?a��>��������>��˾���?q,�?N������=�	��}��Q߾,�>r��=j�=%3ͼ��Ɯ@�vѾX9��v��F�=Z%�>�d@�ε�4��>��D��ݿ��ο.D��@׭�C���x�?M�>��!�2\����h��o�`�B�=�;�L����>sQ>#+ϽV��_���]>�;�$<���>����z�>�]������ԑ�>�R=�ʘ>��>�X�>�ͽ�о�d�?����̿E���G�Ëb?R(�?�H�?V?��< x���z�~�9�A?6�k?�;^?d_!�e�f��I���j?�n��{�]�+�3���A�~�Z>6�5?2_�>b4+���"=�>}>�>E�>�.�ʦĿȷ�g������?�!�?���
n�>ҋ�?ɴ+?:+�ѱ��Qu��:�,�nC�;	�>?[3#>�l������M:�z6���*?g0?�(�Ҙ�]�_?)�a�L�p���-���ƽ�ۡ>�0�f\��M�����Xe����@y����?L^�?g�?Ե�� #�e6%?�>c����8Ǿ��<���>�(�>*N>}H_���u>����:� i	>���?�~�?Qj?���� ����U>	�}?�)�>��?J��=<[�>(h�=�簾��*��i#>&1�=4�?�ܔ?A�M?�I�>iA�=9��'/��ZF�nDR����C���>7�a?�L?�=b>)��J2�!��hͽqI1���8A@��g,���߽�)5>b�=>�>��D��Ӿ��?Mp�9�ؿ j��p'��54?-��>�?����t�����;_?Nz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>E�Խ����[�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ii��	?���P��Ta~����7�W��=��7?�0��z>���>��=�nv�޻��W�s����>�B�?�{�?��>!�l?��o�N�B�~�1=5M�>̜k?�s?�Po���g�B>��?"������L��f?
�
@~u@`�^?* �ӿ�I��Pg��E����=H�_=��=�ܬ���L��:0�<�����=c�P>J�=��k>�wo>�	}>E*T>8���n��θ��%��j�\�K$�0k�/� �������#�QI��� վ���dZs�7��鰾h���R�����g<�>?M�;?��S?l��> K�!�>�پ9�g>������=�χ>�h@?�C^?1A?�!>;���Bd��ځ����ʾ���ߙ>PR>���>��>�y�>�=m�">��=��[>�b�=���=�@���E���!->��>$	?~r�>��ý�/�����a���:���߽�A>q1�?(6���5N��Y$e��Kl�O�%��e?��>]Q��Ӑʿ�<��ݍ*?����K7���lR�g��>I>?C2�>n�>���l��m����׾)$޾Tw��A��{x��M2O�S׼�i>?|-���)>�(�XY6���'���پqr�>�L?Cݝ������_���n�?�پl[N>���>1&>�`!������r��Ct`��J?>��8?9?�����(��1��j3꾉e?ղ�>��>��>,��>�֔>'7�<���"�>k�>UC齋�?��u>6�r=��>S}����X���a>�e>7[>�?��B?'fg<Eь���U�Z�@�A�>���>���>h�>�����h�;]��>�}>��̽R$��彐󏾭{�><������a���A>��=;��=���=�\$��晾,��~?�}��㈿��e���mD?�*?��=�/G<]�"�4���K����?w�@l�?π	���V�p�?k?�?o�����=*x�>�Ы>(ξl�L���?��ŽDĢ��	�p5#��Q�?
�?A�/��ǋ��l��4>�Z%?��ӾPh�>yx��Z�������u�{�#=R��>�8H?�V����O�g>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?roi>�g۾=`Z����>һ@?�R?�>�9���'���?�޶?֯�?�I>Tz�?rws?o[�>��u��D/��3��|���Z~=�W;U��>)�> ���sF�Y͓�Ia��h�j��~�/ab>�M$=�>a��*����=Zɋ��2���me�﫷>iq>�J>	.�>"� ?*Q�>��>h=[N��8ǀ�����L?͗�?�����m�~�<���=�]��%?DP4?S�e���ϾS!�>
�\?��?��Z?�N�>.���1��E����G����<KK>�M�>:��>�7��B�J>.�ӾeE��N�>�Y�>y���۾A��u����|�>�� ?bj�>�e�=1� ?�"?b�w>Њ�>-%D�����;mF�f�>t4�>??�~?�Y?wƶ���1�+L������{kX�)U>�7x?%�?ց�>����l��hT�T���
���E�?Vh?W9꽂�?�?�?�>? �B?�om>�y ���о����*�p>��$?�A��q4�S��i���?�?�(�>e����>��'	�w�0��&˾w?[P?�s'?��-�g��V����A<��M=ؒ<����ԾS=�Z>��>�.'=�=���<��<��������i&��3=Z9>1��F/����-=,?��G�Tۃ���=��r��wD���>�IL>p��c�^?�i=��{�k���x���	U�� �?��?:k�?T
����h�N$=?��?M	?�"�>OJ��S~޾(�྆Rw��~x��v��>C��>йl�j��������EF���Ž��{�?	׷>A1�>�?밐>)��>?yH�h��"�����cm�T�g�9��8��3�ѧɾO�J��}=/N����,�yԷ>3�μ���>xj�>�}>��>3��>l�W��->q�[>�0�>���>�f�=+L3=g�>5}t=۹��S?�6���X"��(پ&L��n�E?]?���>�:]���{�����?��?(��?*�|>�I\�e2'�x�>���>L0���b
?;�<.L�rDd<�v�� �w��<�+ż��a>�+���1�y�>�U�a���?�� ?�[����ܾ'���W ����k=�{�?�?)?A�)�7Q��o�x4X�6�R��.�f�f��٠�s|$��op�k��.\���惿?(��h0=�|*?��?8����ꀭ��gk�G?���e>J�>���>��>��H>x�	�El1���]���&�'����>�z?N �>#I?�<?��P?5;L?
9�>V5�>ON���c�>*�<��>��>��9?�.?��/?��?X+?��b>���c����aؾƸ?�??6>?{L?��?k����ĽbF�����>�z��By��1�=�$�<��׽�^{�:M=l�T>�r?���=�[��ﾾı�>vF?�<>�X�>[����'Ͼp��=�!a>���=hL�q�kg�����4�>�z?�B��^��=�1W>,�;D�s��P�����=��=@�7>��!���<�Z	<�6,>�5�=z�'�M��Z0=]�=�P�=���>F�?�*�>�p�>�������դ� ��=��O>"FN>�%>�,Ӿ����@���0[h�x�q>���?�a�?H�=-��=X=�=�����=���P�����ؐ�<��?f=!?ncQ?a�?�	<? � ?�>>��C���~��x���
�?�0?1��>ş����@��ٜ�{,?�X�>+PC��E����B��U辣򔽘5�=��D�k����!���:���=4���|{����?���?hB��|u1��h����C����H?c�>��>#~�>���T*N�S���AI>G��>}�E?�>	�0?�r�?�l?�zf>a�� ���ͩ�h,=\��>&�,?	�y?uY�?`�L?۶S><io�ޟ���¾X���k_���1����L�Y`E=Q�]>ܴ�>�!?�>=Ma=�`���S��H���x�=}5S>@�?�>��>��S>�ި=0�7?��>�ľ�'��E���G��������g?3�?�A%?��o=p@��(*�M.ҾG�>���?ٔ�?�>*?V���%>B��;���G��A��>���>*)f>�=�k��:z4>�u�>>R�>�CV�9�%���G�e����@?� J?��>��ſ]q�x"r���N6J<����d�˚���y[�v�=�ژ��W�-��4f[���������p඾sN��C=}�KA�>�]�=-��=�i�=(W�<����j��<�J=5�<Z�
=@f�O�y<m:��I���ɋ���F�5[<�DN=q�޻o׸��o?�]V?H�8?��E?k��>�\�==	ݽ���>�z�I�?׳u>:�q���ž��B�Pָ�b����;�붾E�a��ҧ���>�R��G*>(�j>�1>�
1=��=��=Τ�=��L��(.=]�=���=P�=�2�=��>�)>�6w?W�������4Q��Z罣�:?�8�>i{�=��ƾp@?��>>�2������xb��-?���?�T�??�?Ati��d�>P���㎽�q�=B����=2>_��=��2�T��>��J>���K��#����4�?��@��??�ዿТϿ1a/>��=��=�E�Vh1�3�K��3���:��#?cJ5��޾UO>`=S=���N|Ͼ_K�=ilE>�}����t&�\�==�)�}=ͨ=̯�>9�>E�?�U���$ǽaI��0�>�J>!�3������=���'�-6I=���>C�i>eV?W!?0C?�Ec?AP�>�∾yF$�_�c�>��>Xq
?jop>��>�N�>=��>��Z?��u?�N
?7g#>���>V}�>�Dd�]P�/���й�'S�����?N�j?�T�>6aC>l���i��	���>^�W?L�`?=��>.;�>�U����.Y&���.������;�	+=<mr�*NU�\���,m�����=�p�>���>��>^Ty>��9>>�N>��>ª>�2�<Uo�=�̌�rĵ<a������=���$ �<Buż������&��+������;��;d�]<h��;o��=g��>/>g��>���=|����$/>H�����L����=-��OB�h0d�E~�^/��D6�c�B>�UX>�u���)����?��Y>ҏ?>���?�2u?r�>�)���վ|M��V	e�}3S��=�>7D=�6};�W`���M�gUҾ*?�>���>���>�w>� �ͻ.�[�>�۾u!����>gs��Uc���wн1�f��L��N���&�e������C?M��L	+=���?�!\?���?�L�>�#��+�����=�J���1>̿��;CX��E>��!?�8?j��>��Ѿz%����h�ɽ���>� ��K��T���#3�'���K����>�G��qtľ3�+�CL���͑��B��P^�ဿ>�P?���?8�4������P��z��I��~�>Q9e?��>�?3W?�����Ak��o�=��s?v�?P��?`��=f��=����f.?��?@��??�sT?������>�m�=��A>��Z��U9>��>�� ��0�<z�?�� ?�9?�*�����Z/�p���p1}�"�3=+�O=#6^>!z>�K>D�>��<�X=�a>e�_>sk�>�	}>�ӷ>� �>�|~�&/8�!|=?>�>*i�>�f6?���>f;��3a�ۚ;>���:|����Ƽ�C2������=Yq>�V�=��>��>�(�Q˃?���>�����>����↾,�*>�� ?���g ?tYp>�9>��|>qRm>�^�>�r�>�1%>DӾ�>U��W!�HC��VR���Ѿp�z>s���]P&����~��N@I��z���J���i�n0��?=�Ã�<Z8�?ȶ����k���)��6���?EU�>�6?����q����>*��>���>]��҇���̍��g���?*��?m	d>�Ǟ>�AX?��?�x1�s�1��Z�
@v�X�@���c�:�_�}���K���p
��*Ž�6_?@�x?�A?�^�<{>�΀?�=&�j�����>�/��1;��,D=Rҧ>�$����^�GӾ�þ6U�?pG>�p?�*�?�?B�X��D�.>gO?��@?�at?*A7?
0(?��^���?(]h>�?,$?�.;?�7 ?9,�>��=��=Q�J�n�=�ؙ�~;��������������=�q=�;!@�O�m=��=?((�'�μ��=CR����;�xa=�n�=�>��?ČZ?�"�>���>��)?'��C�႔�e&(?d,�>�g=��ҽaa��S����>@ߐ?4�?A�P?�>b{5�pn�a!�=tԆ>1�u>��G>� �>�tԽ5㍾]��L�=~鹼P������[�`��������ݽ8>�=�p?�b�>�鿽y��=}po�X1���x>���x���u�{��	B�D�9�YA�?"�>6??��'?iN�<�� �b�� pQ���%?93?�9?�~z?Nh�=2�Ҿb�(���Y�W2L��oi>���B_!�0���;��%�H����hT>Ȋb��5ľ�Qi>5�m�ܾ��t���^�t` ��Z�;q5���aF�4�žIc�c�=��
>k���-1�������A?��=�_��jK�\����u5>��z>���>���;~��T8��=����	>��>R?K>t�,�N�߾>�:�m���d>%x<?�M?[W{?���[�{���0�t� �0m��V�;���>��>�n?�Hw>��=؈��h���^�bdT��/�>7>�>����uO�Xo���f޾��%�E�>v��>��c>��?��^?�*?�h[?~0?_�?Zt�>Iܻ;Ͳ�gj?(�x?=h4ٽ��2���"����>�2?f�"�gG>&z?��/?z;?�S?Hb?b��=����3�A����>�aa>�p�!<��[U�>D]?��>�	W?i�d?��=��aԉ���w��->�=+o5?C~%?�`?��>t��>�iϾ�(N>x��>��{?��?^�e?E�$>(�>���>=�?Br>�?�a?^�>�N?�s?��Z?��,?���<��ؽ���#�	l��k=\x�<׻>+,H=�I����]��ѽ�_>�GU<�S�=T��<����`�=�C��~r�>G?t>�ᕾ{�0>M�ľs��� A>�2���l��m�����9��\�=��>�?5��>�#�B:�= ��>m��>����((??-!?�k�:"�b��ھ*TL����>�	B?���=T�l��0��4�u��i=��m?��^?�wY�Z����b?��]?: 󾲾<��sľn�c���L�O?L$?�2G��>3�~?�#r?���>�d���m�{�Y0b���k�O�=˛>����d��u�>��7?&h�>��b>���="�۾��w�M���K?��?YƯ?��?c�)>T�n���߿<��\���u`?���>F����]#?��<ՕӾՉ��o��*1�b�e奄8>������ ��wt�A?���d�=�?�Dp?�q?Į^?� ���a���a��;�"S��������O�@��H���H��nn�ٲ����^�I�p=V[��R���?�6?�N��H�>y'U������Aþ�Ii>�l¾��Žk�=��5�Xj�<��=6S�H`��o�?0?ِ�>g�>�s;?�"U���6�Q@��\8����ʻr>��>â�>4�>�����O���#�`6���I��-q?��>�>��b?a�F?L�h?y�K��;�8o�n�>W?=6������=>�>��>f�G�mн�"�B}7�*Ll����J���U�x��:�$?;Q�>TS�>�A�?��>Ե���¾�<����-��s�=���>�Z?/{�>GxI>��iI�X��>��l?R��>�C�>����d!���{�I�˽��>�٭>e��>>�o>Ca,��\��r���}��H9�F��=��h?�i����`�˅>��Q?�@}:ոF<^�>l�v�o�!���򾍱'��>=�?;��=�;>Xž&���{�g��h)?\)?���%�'��S>��%?`�?~��>S�z?�9o>�پ ~-�'�/?G�q?�L?`mI?�%�>�iM�T������ӗ��1��=�y�>�%>�h�<f��A1þ�)5��N�={��u]�F�o�{7�
��������9�8>�*뿺�n�0~��G��d��r�O���D?�����ꌾ���V���ξ��/=�8=����\<������ԃ�wJ�?D��?�G����N����r��̜��KD�>���y����H��S<��1��q���>���v��󙆿;L���3?����s��t����߽�vA?��&?�:�?d,���4�7�.�d�Ͻ�~=�E�y?��(.����ʿQ����Q?��>��˾��=�'�>�[<&:>C��>ej-�.Sƾծ*�M��>4}&?�)�>$�c��繿WĿK3��i�?�i�?�_@?e>/��屾�:>`T�>�
?CK�=��|�?$�_Ǝ���>\E�?K�?���=u�^�$}��h?<��<�+�%���5m�=x�=����վM�J�%>��>��ɽ�b�^O��*>�-�>'���|A���>�� @�y��>���gx��5Մ?*{\��f���/��T��
U>��T?�*�>R:�=��,?Y7H�`}Ͽ�\��*a?�0�?���?$�(?;ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�ԅ�=Q6����{���&V�n��=W��>X�>��,������O��I��T��=r	��Dݿ�#�f���ſ�=Z,�=;�̽��$��*��=1��bg�#d����l���>X��=���=�Ћ>�Hs>Bv�>��E?�o?�B�>1��=�rc�
�ɾOԺ��m=�uT����������)�5O���շ�$������?�����-)��Ȥb�Q��=U"^��Ʌ��~G�V���I�H��>E֙>x{�Ni�\ӿ=����J��)B�=����$��6P�I�j�m�?�8?�j�j�a�Q�˾wx>ȼ�!AB?�������ԛܾiS�>M��=�(�b��>r�x>���:-��o�hE ?�?(ɽ�yG���6=S���<��?��?)�=o��>'�[?J�ھbRV�D�>}��;�	�>V(?߮�f_�Q���5�&?۪J?r���y˾�%�>���W�=>9��=ŀt�����^ >$8F>�)>?=�1��<謁�����W?�>q�)�g�������"��H>=�gx?S�?Oh�>�%k?�B?���<yp����S���
�=\x=Q�W?��h?\g>#����Ͼ�P���5?K�e?��N>Jh�S�]�.��^�$�?��n?�n?�˝��D}�������TD6?��v?�r^�ms�������V�@=�>�[�>���>��9��k�>�>?"#��G������lY4�Þ?|�@|��?��;<��"��=�;?a\�>ݫO��>ƾ�z��������q=�"�>Ռ��yev�����Q,�^�8?���?Y��>���������/>k��Zݱ?�S�?#S�����=���OI��(M�G�T>�hI=�0�=s����2�_��[׾U䰾ˮm���i>+Ă>S@�hѽ�U�>����`�տ`Y�&|�Kc���z�tY?Sf>�U���R\���U����b��&c�&�$7�>I�>���zY���"���k=��|�=�>Q�z=U��>���c4��ɫ�(�Y>/��>\��>��?>���W%���Z�?�=����ҿ.���lҬ��p?���?�݈?:!�>�������4ҽ�'
<S�N?@�S?�
]?oƵ=�����H=t�j?T����_��3��KE���V>��3?��>�-���k=��>�>�>Ę.��Ŀ�d��Xu���Ŧ?�M�?Gx뾽e�>W��? _,?��	t��,��rz-��Ǫ92�A?��2>�˿��F!�t�<����-2?�>1?�=
����_?ՙa�_�p���-�x�ƽv١>�0�f\�"&��W���Xe�����;y�B��?�]�?��?^��� #�N5%?d�>���I:ǾX��<=��>+�>`*N>.E_���u>"	���:�5g	>h��?�~�?�i?m��������R>U�}?�%�>��?6w�=Ka�>��=���Y�+�c#>Uw�=��>���?��M?N�>�A�=��8�M/��VF�VDR�C%��C��>X�a?��L?XHb>n���#2�>!�x�ͽ.g1�M�7p@�G�+�'~߽�'5>G�=>��>x�D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�c��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?kQo���i�B>��?"������L��f?�
@u@a�^?*XͿ�����Ŷ�aY�s�c><DY>�_�=���'�=�O.>�c�=J�*��*��=�>xu�=��#>�l�>e2`>�a�>�Մ��#���n�k�,���`��5���������!,���'w��}��D=�+L��H-�v�S�-Ð�̤�=r�=��T?��O??�n?c��>Zޔ���">l����=a��P`=�҃>�3?O�L?�|*?u��=�_��"3d�]避�1��`���l��>��>>�A�>�Z�>�ȩ>MҖ;�,:>,.E>��>�2>D=��;�(=�NR>��>���>��>'5ӽ1A	>�޲��ѷ�(���y�+:U=׋�?U����o����c(�ӳ��A��8O?	��>����b�Ŀqʯ��$?�7�������Y�Q_t>�*0?��N?6ۉ>�ξ��8Յ>��ߠپa&4>@��:p���fܾAE>R
�>�ғ�\Q�>�A���/��1E�,e����?��4?!��P(
�v}��$`�ui%��~	>�?C{;P�I������m{�0��J�t=O�B?�(?K�����\c�G5��e�q>m�?A}���r�=.�>��>�'���,��b��>T1>�mt���?8fq>_X�=	 �>�̾Q��X��>�>>dB�>�??	w?ܖ�=���v�������t�i>S��>3�>2�=�*G��a�=n?�ك>�4��o�������J��?>�[S��4���R&�մe>v�5�on>)�=݃Y�������~?���'䈿��0e���lD?X+?] �=��F<��"�D ���H��G�?r�@m�?��	�ۢV�9�?�@�?��C��=�|�>�֫>�ξ��L��?��ŽAǢ�Ȕ	�)#�eS�?��?��/�Xʋ�5l��6>�^%?��ӾOh�>zx��Z�������u�l�#=R��>�8H?�V����O�f>��v
?�?�^�ߩ����ȿ4|v����>V�?���?g�m��A���@����>;��?�gY?xoi>�g۾;`Z����>ӻ@?�R?�>�9�|�'���?�޶?֯�?_G�>&�?y��?�V?�
����)��=��G���&����<���>�]���a��v*��<���w����>����?�G>Vj�=Ko�>@Rٽpg��;��<E��ɝ�%�8��FF>����[>|YH>1?R<?Y;�>�2$>��ڽ�ߌ���C�K?�q�?u�>�m�**�<�`�=�Z���?��3?�h�{Jоϧ>:]?���?��Z?�t�>t��$������:��v�<�VK>���>���>���pfH>�.ӾxwH�JP�>7�>�4��� ۾%(��m2��t�>II ?�:�>@
�=�� ?��#?7�j>�L�>�YE�
5����E�Sj�>Ҋ�>�H?��~?<�?�ӹ��j3�G���衿��[�p
N>K�x?2R?Q�>���K~���F��J�3ᒽ���?�\g?���? �?��??G�A?T�e>,��ؾZ#��P��>��?��Q?<��j+��;>�'?�b?��?����J��Z����5����޶�>OEg?��?)n�ale��QȾ��a=�`<�=dO<7]>ȈO>�F>w>����=���=�J��~�����v��=��)=W"Ƚ�%�;�>4,?�.1�����M��='s��D�fe�>	�K>�վ�`�^?��=��{��ڬ�Z���uS�Fٍ?�?-A�?�g��ch���<?�/�?$?_�>Ap��;�ݾF�� w���w�s��{�>�.�>2pm��J�QF��И��_a��Q�ǽ�s�%*�>���>��?'�
?qߪ>1�>�0Ծw:�
������o��"��;.���1����蘾9�I�Q��<�1Ҿs����l�>�䴽,��>�?H�g>~]f>���>�V�<�l�>�+> �C>���>��e>r5�>}�8>Z4�8F�xBR?�����'�5�� ����5B?v�d?��>�f�4t�����Q?F��?6z�?��v>p
h�7+��?���>z���Y
?�*8=EF���<X���?�������&]�>��ս):��M�Zg��<
?�?eD����̾1oֽJ����o=�M�?G�(?a�)���Q���o���W��S�މ�0/h��f����$�b�p��_��$��P�(�Ջ*=s�*?��?8��-������%k�?�Hbf>���>�>��>7gI>��	�X�1�V^��M'�о���H�>�N{?�J�>��I?g;?�O?��G?���>|��>�4����>�U<�E�>�f�>�\:?�/,?k�0?��?�*?��_>����[9���پ�?>�?� ?fj?�?񔅾��սBϼ��E"���K��#�=�l�<�սG퐽c1,=�)O>M?ƥͽ��5��`����>р.?���>���>>����k�yä=A��>�V�>��K>����p������4�>�u?;����<_>�k�=���y56���=5��;�!m=x�0�ܝ��Y�<i�=ʨ�=���{��(�%�c=y�	=s��>��?u��>6͈>�؅�� �h�����=BY>%U>>�Aؾ*e�����Ĉg��z>���?�q�?)�h=m�=�C�=9Ơ�������,���+j�<��?�7#?��S?T�?�>=?R.#?,>��������������?��-?5W�>)Ծ�6������9+���9?�'?Οd��	��\��rpҾ�,�<���=	^�xS��bK��B%�z�>�X�~d�����? ��?iny� 1*��,��@��{�6��T@?��>Y��>�?�h��v����D�r,�>jy�>��9?���>���>٩�?�?�2#>�>ݧ�p� �*��p>'U?G�q?��?^C�?B��̪�=i��;����|����c���j���X�=s��>���>ʈ�>W�>��T=���=��ϻ��D<V冽rVo>0{?5Â>�n?�O�>D&>W�F?��>k�������������˽(�n?�F�?�(8?�;�=!	�m<��澂S�>���?�ث?�s/?��:����=b��F2˾�爾�\�>��>�~�>-��=�=�>)-�>���>�qӽ��9V;��1ټ��?Z�E?��%>�{ƿ)�i�4���F��ݘ��Ӄ����W۹���E��JC=(���U���ɦ�]u�j˝����U?˾�j��2������>�,�=|�>�B�=Q=ԥq����M�==U�d=�<�l��5=���F�l�cS��� ѯ<R�e=O�0��l˾�}?�I?�t+?��C?E�y>�>=3�7Z�>k'���M?�BV>L�Q�m���As;�ʨ�N����^ؾPc׾��c��ȟ��%>��H���>i13>o��=��<4��=��r=��=E�R��=GF�=?l�=�d�=\q�=�
>�V>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/> ��=�ei>?;O�s�X���=�iH��̅�ݏ ?5�6���ýF��>���>�Y�	�꾑��=4�=�r>3�{>5J��>b��e�.=cD!>w��>�>zxd�xS��F�V=�xCz>�pQ>�q��-��ҽ�f���Ή=
�>���>�?D��>^�O?�`?��>!ؘ���� &ɾ;�A>��>G?{,�=�*�=�J�>�j�>/L?v�g?�{�>ÐR>'��>_��>`�
i�]����̾�G����~?�j�?���>rK�=�����*����=�!G?�?��?�>M>�;�T�㿳l&�9�)��hx���<�j=i{���a�j%�sV
������=ʶ�>�A�>���>L�z>8@>}�]>�p�>��>�f�<I�=�Ri���)<������=����k'7�������v:*K�ҵ���yݻxXȻa�m�o	<$6)<���=y��>�K>
��>ޕ=�'���b/>����H�L�U�=�Z���!B�Md�t@~���.�;D6��B>�X>	Ą��.��Y�?��Y>�c?>N~�?RDu?��>,��վ8N���se�ܐS��w�=A�>?�<��m;�|c`�>�M��{Ҿ!��>Ρ�>X)�>�E�>��c)�� S�=b���A��)�>��w��Z�4/�;fd�J�������2�Y��f98�J?㈋��d<���?��A?�%�?�A?!�$�.F=��QZ=
�l�ȗB=��1������ۼ���>Db?#�?�&��6��H̾���l޷>�@I�:�O���y�0�F���̷����>�����о+$3��g������܍B��Mr���>��O?��?�9b��W��UUO�����%���q?�|g?r�>�J?�@?X#���y�r��	y�= �n?���??=�?�>��>��b��>5/?n��?��?�0b?��I�.�>H��=�Sg>KB����>�P>2����>�?li?1"?E	���W��`羜5㾅?���=(*>���>H�o>��T>�+�=y">���=��l>�`�>~n�>�I>�>��>�-����"���9?���>> �>ä7?���>!�b�� ��\�=��h.����;��=�|I����=� >9�>]x>.*�>�ÿO��?���>��%�(��>����2��V�>^�>����eU?b�=���=v�>(�I>B�u>��>��>Q�ҾN�>���5h!�:�B� R�ACѾP�{>�̜���&���.���3)I�~g���$���i�?1���*=����<Q.�?�����~k�F�)�Q�����? @�>+6?�'������1�>Z��>���>�H��ł��[э�Qo��?��?W>c>4�>��W?��?��1��3��uZ�Ԯu��'A��e��`�����������
� 	����_?J�x?yA?�l�<�:z>d��?*�%��ԏ��&�>/��&;��K<=�-�>'��?�`���Ӿ�þv9�:LF>Q�o?�$�?�Y?<UV���j���%>6�:?��1?8]t?��1?0;?�q�x$?�3>�q?d�?|F5?��.?�
?��1>���=���c+=�I��/ϊ��Tҽhw˽��꼭"3=�|=E':�	<��=�i�<�D��޼��;�}��4��<I7<=@У=20�='&�>�l?��?�>��?F�����K���E�R�]?ަ>8|<=䴏�.1��Wᾼ�<�h�?L�?9�m?�>�N�ce��U	%>�ʌ>���>'�->(~�>�/������#=���Z=�g�;�*>�����dg�����������A�&>�@ ?�x�>�gνR�=�Ӊ�("A�-�>�B�'�����R�IF�Ɠ.�������>rJK?�"?���=�����ʽ�'T��%?=�9?�>?-�?��=����%���U�Y�,�5:�>�IE����j���	����<��n���J>h���9�ȾW�A>aH����s^�"B�B_��{��<̭����<����Q��ew�#��>-Ǒ>�OþB��l���e��,I?�`�=c��a�Ѿ�`^��/�>��u>#X�>iG�q��T�"��Ծ��%=��>��>��=B|Ⱦ�_U�Lp�2�>�D?́^?j��?�ׂ��r�ѽ@������4����̼!?�y�>=�?;TI>[��=n<��ڟ���d��F�)��>g��>�g��I�贛��&�A�"��w�>�O?{>c�
?�"P?��
?�|c?�I*?�?�Y�>�˽Z��� I#?u�?��=�ޯ�d�K�O6��=�L��>r�.?jK4�쮊>��
?�� ?8.?�kM?�K?�>���~�7��h�>���>l�U�ů�<b>y�L?"ײ>�Z?ۻv?p�>�5�gZ�������&>e�*>C�'?I?�-?/��>�%?���J R>��?��?��k?S�J?��>���>���>p�>�T>o�Q?#K?�g>�{?/~?7�B?p�2?/�=CN�����"8� �8=@�<�2G�k�u>�8�=@B��,�_�?�=r{�=b�>쀨��}��d���4�p=!KU=�f�>��s>�ە��1>��ľ<��^�@>�n���L���Ǌ��<:�O��=n��>��?mc�>R�#�i�=c��>�X�>����+(?��?�?��+;äb�b۾ѦK���>�
B?���=q�l��t���u� �g= n?�^?��W�@(��C�b?J�]?����<���þ&�b�T<���O?,�
?ֿG���>E�~?�q?`�>�Ke��&n�*����Jb�?�j�<y�=+Z�>ol�ze� 5�>�7?�I�>�Qc>X�=7e۾s�w�U����
?{��?��?w�?�,*>b�n�����v����]?sR�>̯���)?�Oh=��40���X@��h�ː�"�����{�Ӥ���i�K��p���=�?aj??xs?`�a?����t_�!Lh�hք��S�Ӻ񾦏� �=�yU��dL�$Xr��D�����ܜ�Q��ky[�|W`���?�6?�Z�*a�>av�R��5 �����>>^Ǿ`�q���=W|�;:C=lQ�=N�bR̽�V���_?5&�>	�>$�D?�pQ�_S.��ZA�(R�Y���o1�>�0�>N��>nx>�+���k��xcU��s��.mg�_�e���h>Sva?Z�F?�ia?�p;�?�7��k��L�=t&=k��� �=���=���>B����̽���Z3�HTd�a/��9�����mЬ=�\&?�Գ>��>6É?@��>����Ė�!�v��1�v>&�?sb?4\�>q e>�]�5���F�>Edy?
[?���>�����0*�%����G:�Ɲ�>u��>���>Gɍ>s�ۏh�*����@��o�8��R9=(!d?�����}��'�>%�M?+�=
�={Ն>�"޽���f��2��\>�D?���= >9V���]Ͼ^Xj�Ŕ�D`)?-H?����s"*�@~>R�!?���>Ry�>��?���>j�¾��A�ޙ?��^?ǦI?�-A?T'�>O=Ě��|oȽ�&�b�+=ֆ>�q[>!v=�{�=��h�[�%���bA=��=��ܼ���`��;�侼��6<i�<�r5>;��&$b��0'�����yV��uB���$������ t��	�k	�	aŽq葾�6	��=��Ӿ_ ~�Z8�Q�d����?�?�?�Y�#XR�bɏ��r��VX����Z������=F�j�5�=%L���a	��>�ڥ#��#a���\�!�n��1'?	�x��뼿m˛�-��"�-?G?!?��z?�����6� �5��j�<)3=
A�����ҙ�-zɿ�s��Ԣ\?r�>Bپ���:A�>�0B>�&>[�x>�����ة�J��<��
?�k2?>'�>�[���Ŀ滿?�<�P�?!v@>A?^�*��x辜w=1N�>�E
?/�G>bG7�����k\�>7؞?-ʊ?9�j=�W������!f?�Dd<V1D�ĢN���=���=�D%=���J>���>9%�L�@���̽dg->���>�N5�m�2�]��<�[>-	Խ�I��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�}��=[��>c�>,������O��I��U��=
@���ƿh&�������<A�r���V�+�m���!\�Gˡ��:l�Y0콥�s=4R�= TM>��>�~W>�Y>Q�W?�Al?(�>�J>�������=K̾KQ9�Ձ���y�w��?��;X�����ݾ]�
�
f�j��2�ɾhF^�]�G���g��ڑ�*J.��t�J��z�?쾦<���:D�vlw>�/��5[�7p>�<���þ��5���� ?�?;q,?�������ƛ-�醄>u�*>�Sp?Q8½ho��A����ٞ<q��=��p=�V�>�{�>
Hd�_\�'�f��f?�X:?�ƾ�8��N�����p�d�|=t�?F�2?�Z�<P��>&�?cʴ���S��\>Ƨ>��>�� ?��}�社r���jy-?��D?F���ީ���>u�ƾ�d��=������ >=->>�*>���O�����X��<�(W?ʥ�>��)�� ��[���N�$�<=>�x?a�?�*�>�zk?��B?lx�<�\��u�S����w=��W?�(i?e�>I���7о\���#�5?Ƞe?�N>rh������.�HT�?"�n?0[?����x}�K������r6?��v?�r^�ps�����q�V�N=�>�[�>���>��9��k�>"�>?�#��G�����mY4�Þ?z�@���?0�;<��z��=�;?b\�>1�O��>ƾ�z��������q=�"�>���cev����R,�7�8?ݠ�?���>5������Q@>����K@�?�)�?+���,�b=Y�����n�M6�>b�	>���=���S���BH��f��渾�D6�Mͽ=9}�>m%@͞�;�ޤ>�{����7�<�_�D��O�پ�K?q��>3A�g��	�z�K�|��%z��(v���C�<�f>��=3X�M�����D`>��b�����>ޫ�:��>-�G���H�������=מ>®>&��>Q�ս/��G�?0۾h1׿T@���(뾵5Q?���?��?�p�>��W�_���b$����<�\U?#_�?n_?���=���<>�+~j?�@��B_�4�^�D��U>"�2?�%�>�H.�v�j=oO>���>��>/�.�ߢĿ�3���K�����?�s�?�꾌`�>�q�?��+?a���.���᫾�*��t!�%�A?<�4>�ν�2�!��)=�g��[
?,m0?b����[�_?'�a�J�p���-���ƽ�ۡ>��0��e\��M�����Xe����@y����?L^�?f�?׵�� #�d6%?�>d����8Ǿ@�<���>�(�>*N>EH_���u>����:�i	>���?�~�?Qj?���������U>�}?�H�>�.�?��=�!�>�`�=�ݱ�
�@��&">���=*A�R3?�BM?�_�>&��=݄8���.��;F��
R����/�C�Hd�>�b?hL?�Sb>I3����4�� �hlѽR1���z A�`4�Uཞ�4>#�<>1>�MF�r�Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P���`~����� 7�n��=��7?�0��z>L��>��=�nv�ۻ����s���>�B�?h{�?V��>��l?��o�P�B���1=�M�>ɜk?�s?ejo�s󾓳B>��?������L��f?�
@yu@c�^?��`��ǲ���A޾%��B0g=G>�=�*>��F�_X�=�K�
!������*�=�>'�w>es�>��l>eHO>��>�ۅ�W������Ş�u
|�rS�0��ΰĽ>�s���0��X����ܰ��p��-}��>p�D5�}�
�%��=�ST?ԮP?�m?ԓ�>,���">�`����0=��#��zL=��>�e2?z�K?��*?!W�=���k9d��c��季��؉��2�> Q9>���>&��>LU�>��<�O9>�R>>r�v>]>�=}�H=��=��8=HF>���>�=�>c��>h?���r>ڼ�4�ſQ�ʾ$�;��*>4��?}�o��n��?��B轾�c��Vi��/�?WY?t/��R�׸��(�?%rɽ�r���H��N�<hc??�'?��@>�Dq�iqk�j��~!��l��E�ɻg�;�Cݽ��H���O=�?<��;v"�>@�5��zG�(/_�p�ν�h
?�A?��n��u�� ���q��x-��Z��~�%?��=s�i��ɥ���q���q�,٧=��G?��/?z���_�������1�>��v>mP����z>9]>1��:)w�d촾n>��ɻ�[�>	�?��l> �=-R�>8����n����>��->�C�>�m8?��?��Ҽ��콀���τ�L�z>��>�<�>� �=��W�6��=� ?�Op>y15��t���J���+<��:`>8���=���6�+C�=��Ƚ݄>���= �D����R�<�~?���'䈿��e���lD?T+?g �=ѝF<��"�D ���H��F�?q�@m�?��	��V�?�?�@�?��K��=}�>
׫>�ξ�L��?��Ž7Ǣ�Ȕ	�))#�jS�?��?��/�Zʋ�>l�6>�^%?��ӾPh�>wx��Z�������u���#=R��>�8H?�V����O�h>��v
?�?�^�੤���ȿ5|v����>W�?���?f�m��A���@����>9��?�gY?roi>�g۾9`Z����>һ@?�R?�>�9���'���?�޶?֯�?Ǯ>���?�O�?Wj�>dռ�mB�tJ���m���_�6�{����>�H�>E<����a�����r���y��)����>�<K\�>�S=�T�����=�\���ם�螳���=y3=>Ql�=;��>�?��n>u��>i�<���<��_��L��\�K?���?����0n�� �<�Ҝ=O�^��(?f>4?\�@�Ͼ齨>��\?�À?d[?�^�>y��?��(濿r��`�<��K>�*�>G�>����<K>��ԾLD��c�>�ʗ>�<��X@ھ�<��)����F�>�[!?*��>��=�s$?'�2?\��>���>!60�����=d��5>�)?_Z?]n�?	!??�Ⱦ��4�Z���p%V�ٳ�=��x?�l?���>�ˇ�m[���~N=���Բ_���?�MM?f�����>T�t?�JD?|�'?:k�>ӊ�������{���>z�?@Cu�W(&����kսB�,?�G?��?�(h�����撁���b��5���?��9?ak
?����~x�b����d=J�]����<I�>�~b>�/�=��;��=�	�� >v����n���{_��S�/�h>��v���˽��Q>�#,?��5�"̃����=��r�e�D���>��K>�׿�w�^?J�=��{�%����p���{T�a�?�{�? N�?����h�z�<?�*�?R?K��>�X��Yi޾cྜvw�ۺx����T�>;��>�<v�Z�侜n�������Y��5�ƽn�� ��>���>��?<A?��>��>BF����*�8����پIc��
	��p=��<�.� �:ӗ��)#���<�̾*��f�m>#�ϼ�>f�?�X}>۽B>���>%�w=y�>y1,>OO}>�p�>`/d>@.�>��l>z=��}��ER?����?�'����௰��3B?�nd?G7�>�ci��������|g?�?�v�?�Rv>xh��%+�cV?��> �� j
?o�9=�+���<E-��ּ��ۆ�m�P��>�R׽w):��	M���f�;Y
?�,?����0�̾�M׽^���D5y=�L�?�m%?��(���X���x���\��@���귓������*�i�r��ƅ��x��@��6�/��<!�%?|^w?q����5F��EQ`�x�D�D`\>~E�>���>;�>�b�>"0��b �>�k�K���Yi�>�Pd?.�>M�F?�nE?��9?%�9?#6�>C��>̂��D�?0�>P�>�O�>�?X�+?�D?��
?�*?�c>!�?=����l�۾_�?+�
?>(?�D$?�6?�6���y5��T�=�K��sþ�.w�l30<��=`(��i�Z�=���=�y?"�ӽ�M-�>��Z��>��L?���>�E�>/���
ԾJ&���/>>n�>$�>��	��k��*�/Q�>Őx?c�	��}�=��G>M��=8�������d�=��$�zB	=�߆�k��<Nb8=J��=��=M}�w����~<Z�=W�>Vj�>��?�p�>&�>�Q��ݤ �+�����=��X>S>QE>=0پ�{��'����g�EWy>�p�?Gy�?l�e=�*�=1��=Lv���3��H��S���<v�?�]#?�HT?���?��=?�^#?��>��.@���S��V����??]?�O�>�)��/��o듿�D��E�?�(?�C��=ھ��1�mJ�W����=F�$�w��N`��;�8�E�=dn��w�/��?&N�?r�;�CX�?�$������¾��X?��>��?�7�>�F���|���2�_�s>G?�nA?��>�� ??>�?�t?���>�6�L ���[��pżn`�>�J?�1�?棃?BE??-K�=]��<�f=��Ⱦ�\��
����Qz�Kف=�#o>��>��?�GY>�%p>��K:Ux��b���9>���>V��>CO�>N�?�d�>:"J�{�G?]�>�ľ�O\������郾�)@��u?��?��+?�=V�7�E�T������>�t�?��?�7*?TS�=h�=c�Լ%嶾c�q�� �>S��>8)�>=̔=��H=�S>���>�i�>����D�C8���M���?�E?�׽=P|ʿF�n�?}�������f�F�̾������	�����k�=\Ҙ������ȯ��j�ˌ�0��"4¾�n��ﻎ��l ?#��==�$>���=<��=z"4��ҥ�z�.=`��R�=7���zH=����U�	��u���c<ڎ�: j��z��j˾ԕ}??I?��+?�C?��y>4�>f�3����>X����A?�'V>�
Q�-����;�5����8��,�ؾFZ׾p�c�M���_O>S�I�ض>T'3>d:�=1^�<��=,�r=`��=*�S��J=<��=h�=V�=��=*�>�D>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�1�=�>�Y�a�I��
����,4����(?�d���^���?8 >�(�tb���=>r���]
>���>�M�e��=��=ܲ=-��=::>i82>R܊=��ͽ�-�=��6�=p�=�5ͽ�񇾝4�J��=T�=�>]3>w?a��>L9;?'[?��>�(|��<���»�v��>�$�>_
?��=��>K�>%��>�-\?�c?%�>���=1�>m[
?QD��Ej��Ͼ���D�p��?�C^?P�>��9>G����c<�#��<j�8?���>�j�>h��>�U����:Y&���.�&���֜4��+=�mr��QU�B���Fm�-�㽱�=�p�>���>��>:Ty>�9>��N>��>��>�6�<wp�=�������<� �����=1�����<�vż�����u&�L�+�1�����;q��;��]<���;��=<��>2�>�K�> M�=�����.>'��MK�97�=k�����A���c�j~�$D.�ޭ5���A>1W>�∽5���	?��\>��A>8=�?h�t?H>T��*׾V���Jf�C�T�VW�=|	>�q;�P;�|�`��JN�.Ҿ���>��~>�c�>�ׄ>8�	�]1&�c�ݼ:Ȩ�^hQ�O�>�1�����3c��`��]��b���n�\���<�*P?�G�����мc?�LT?ZN�?ȶ�>��;�� ���g>�/�/� >-`��_�G�2vI�]J?.W>?�?��Ҿ.C�&sྒ躽��>��/�P�>���/fA�����z������>�]�����Ť)��o������l�E�d�v��A�> k4?�A�?�r�,7��Z�\�U��C���>�!l?&�>3�?�!?k<�:��o���@|=ZYh?,�?�H�?ODs=ʥ4>퍫�?,N-?��?} �?�AG?���N��>�j>h��>P9�����>�$>���/��=�:?� ?�*?C��������)���a���"㽼���>ML�>�g>�׫>��G=k�~>WP>?g�>���>��?���>H��>K��>H��J�0�W#?8�g>G�>@�5?���>r�ƻKܽI�=�ռ����l0^��t=� �;��=Q�>��->�->���>!ǿ3��?7J�>�3-���?"[�����{2>؎�>IXž�>/.>z�>e	?v�>A/ >y�O>G�;���Ӿ>���� ��B��R�!Ҿ��w>˺����)���	�vv���9F�쵾�X�a�i�(5��Z�=�P+�<�}�?AS�"'j�܃(������Y?;2�>��4?�|��pNw�g�>���>�׍>�T��A��������4޾��?���?�;c>��>7�W?�?1��3��uZ��u�j(A�e�&�`�~፿�����
����_?�x?9yA?PS�<:z>I��?��%�Jӏ��)�>�/�';�E@<=�+�>�)����`�W�Ӿ\�þ8��HF>��o?6%�?cY?MTV�ƻ5��>��=?#4?>�s?N�2?�8?497�$l%?5C>g?��
?�9?�/?c?ĝ>��>A�8Na= H��@ꍾ��Խ�ͽ�S�6u�=^�=䬜;V^�<d!�<�턼�(k�б���z<(�e��e�;A�?=[K�=9~�=F:�>�_?N?��>��%?��c���?�RIH���S?��=Q@߽�z����_a����l=�{v?ǌ�?��P?�ͨ>�8P���+���=[X+>�>ݽ�> U�>5nD�y_���=+�y=Ua=��e��g8�M�u��d�C����c�5��>�a�>��|>hǍ��&>����n�x�6�d>��O��湾�SU��?H��X2�aPu�H��>E�K?v?e0�=w@�Hx���e�g(?s0<?�)M?��?���=bܾ�x9��sJ�@y�Q�>�5�<k�G������Ɖ:�`h����s>����9�ȾW�A>aH����s^�"B�B_��{��<̭����<����Q��ew�#��>-Ǒ>�OþB��l���e��,I?�`�=c��a�Ѿ�`^��/�>��u>#X�>iG�q��T�"��Ծ��%=��>��>��=B|Ⱦ�_U�Lp�2�>�D?́^?j��?�ׂ��r�ѽ@������4����̼!?�y�>=�?;TI>[��=n<��ڟ���d��F�)��>g��>�g��I�贛��&�A�"��w�>�O?{>c�
?�"P?��
?�|c?�I*?�?�Y�>�˽Z��� I#?u�?��=�ޯ�d�K�O6��=�L��>r�.?jK4�쮊>��
?�� ?8.?�kM?�K?�>���~�7��h�>���>l�U�ů�<b>y�L?"ײ>�Z?ۻv?p�>�5�gZ�������&>e�*>C�'?I?�-?/��>�%?���J R>��?��?��k?S�J?��>���>���>p�>�T>o�Q?#K?�g>�{?/~?7�B?p�2?/�=CN�����"8� �8=@�<�2G�k�u>�8�=@B��,�_�?�=r{�=b�>쀨��}��d���4�p=!KU=�f�>��s>�ە��1>��ľ<��^�@>�n���L���Ǌ��<:�O��=n��>��?mc�>R�#�i�=c��>�X�>����+(?��?�?��+;äb�b۾ѦK���>�
B?���=q�l��t���u� �g= n?�^?��W�@(��C�b?J�]?����<���þ&�b�T<���O?,�
?ֿG���>E�~?�q?`�>�Ke��&n�*����Jb�?�j�<y�=+Z�>ol�ze� 5�>�7?�I�>�Qc>X�=7e۾s�w�U����
?{��?��?w�?�,*>b�n�����v����]?sR�>̯���)?�Oh=��40���X@��h�ː�"�����{�Ӥ���i�K��p���=�?aj??xs?`�a?����t_�!Lh�hք��S�Ӻ񾦏� �=�yU��dL�$Xr��D�����ܜ�Q��ky[�|W`���?�6?�Z�*a�>av�R��5 �����>>^Ǿ`�q���=W|�;:C=lQ�=N�bR̽�V���_?5&�>	�>$�D?�pQ�_S.��ZA�(R�Y���o1�>�0�>N��>nx>�+���k��xcU��s��.mg�_�e���h>Sva?Z�F?�ia?�p;�?�7��k��L�=t&=k��� �=���=���>B����̽���Z3�HTd�a/��9�����mЬ=�\&?�Գ>��>6É?@��>����Ė�!�v��1�v>&�?sb?4\�>q e>�]�5���F�>Edy?
[?���>�����0*�%����G:�Ɲ�>u��>���>Gɍ>s�ۏh�*����@��o�8��R9=(!d?�����}��'�>%�M?+�=
�={Ն>�"޽���f��2��\>�D?���= >9V���]Ͼ^Xj�Ŕ�D`)?-H?����s"*�@~>R�!?���>Ry�>��?���>j�¾��A�ޙ?��^?ǦI?�-A?T'�>O=Ě��|oȽ�&�b�+=ֆ>�q[>!v=�{�=��h�[�%���bA=��=��ܼ���`��;�侼��6<i�<�r5>;��&$b��0'�����yV��uB���$������ t��	�k	�	aŽq葾�6	��=��Ӿ_ ~�Z8�Q�d����?�?�?�Y�#XR�bɏ��r��VX����Z������=F�j�5�=%L���a	��>�ڥ#��#a���\�!�n��1'?	�x��뼿m˛�-��"�-?G?!?��z?�����6� �5��j�<)3=
A�����ҙ�-zɿ�s��Ԣ\?r�>Bپ���:A�>�0B>�&>[�x>�����ة�J��<��
?�k2?>'�>�[���Ŀ滿?�<�P�?!v@>A?^�*��x辜w=1N�>�E
?/�G>bG7�����k\�>7؞?-ʊ?9�j=�W������!f?�Dd<V1D�ĢN���=���=�D%=���J>���>9%�L�@���̽dg->���>�N5�m�2�]��<�[>-	Խ�I��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�}��=[��>c�>,������O��I��U��=
@���ƿh&�������<A�r���V�+�m���!\�Gˡ��:l�Y0콥�s=4R�= TM>��>�~W>�Y>Q�W?�Al?(�>�J>�������=K̾KQ9�Ձ���y�w��?��;X�����ݾ]�
�
f�j��2�ɾhF^�]�G���g��ڑ�*J.��t�J��z�?쾦<���:D�vlw>�/��5[�7p>�<���þ��5���� ?�?;q,?�������ƛ-�醄>u�*>�Sp?Q8½ho��A����ٞ<q��=��p=�V�>�{�>
Hd�_\�'�f��f?�X:?�ƾ�8��N�����p�d�|=t�?F�2?�Z�<P��>&�?cʴ���S��\>Ƨ>��>�� ?��}�社r���jy-?��D?F���ީ���>u�ƾ�d��=������ >=->>�*>���O�����X��<�(W?ʥ�>��)�� ��[���N�$�<=>�x?a�?�*�>�zk?��B?lx�<�\��u�S����w=��W?�(i?e�>I���7о\���#�5?Ƞe?�N>rh������.�HT�?"�n?0[?����x}�K������r6?��v?�r^�ps�����q�V�N=�>�[�>���>��9��k�>"�>?�#��G�����mY4�Þ?z�@���?0�;<��z��=�;?b\�>1�O��>ƾ�z��������q=�"�>���cev����R,�7�8?ݠ�?���>5������Q@>����K@�?�)�?+���,�b=Y�����n�M6�>b�	>���=���S���BH��f��渾�D6�Mͽ=9}�>m%@͞�;�ޤ>�{����7�<�_�D��O�پ�K?q��>3A�g��	�z�K�|��%z��(v���C�<�f>��=3X�M�����D`>��b�����>ޫ�:��>-�G���H�������=מ>®>&��>Q�ս/��G�?0۾h1׿T@���(뾵5Q?���?��?�p�>��W�_���b$����<�\U?#_�?n_?���=���<>�+~j?�@��B_�4�^�D��U>"�2?�%�>�H.�v�j=oO>���>��>/�.�ߢĿ�3���K�����?�s�?�꾌`�>�q�?��+?a���.���᫾�*��t!�%�A?<�4>�ν�2�!��)=�g��[
?,m0?b����[�_?'�a�J�p���-���ƽ�ۡ>��0��e\��M�����Xe����@y����?L^�?f�?׵�� #�d6%?�>d����8Ǿ@�<���>�(�>*N>EH_���u>����:�i	>���?�~�?Qj?���������U>�}?�H�>�.�?��=�!�>�`�=�ݱ�
�@��&">���=*A�R3?�BM?�_�>&��=݄8���.��;F��
R����/�C�Hd�>�b?hL?�Sb>I3����4�� �hlѽR1���z A�`4�Uཞ�4>#�<>1>�MF�r�Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P���`~����� 7�n��=��7?�0��z>L��>��=�nv�ۻ����s���>�B�?h{�?V��>��l?��o�P�B���1=�M�>ɜk?�s?ejo�s󾓳B>��?������L��f?�
@yu@c�^?��`��ǲ���A޾%��B0g=G>�=�*>��F�_X�=�K�
!������*�=�>'�w>es�>��l>eHO>��>�ۅ�W������Ş�u
|�rS�0��ΰĽ>�s���0��X����ܰ��p��-}��>p�D5�}�
�%��=�ST?ԮP?�m?ԓ�>,���">�`����0=��#��zL=��>�e2?z�K?��*?!W�=���k9d��c��季��؉��2�> Q9>���>&��>LU�>��<�O9>�R>>r�v>]>�=}�H=��=��8=HF>���>�=�>c��>h?���r>ڼ�4�ſQ�ʾ$�;��*>4��?}�o��n��?��B轾�c��Vi��/�?WY?t/��R�׸��(�?%rɽ�r���H��N�<hc??�'?��@>�Dq�iqk�j��~!��l��E�ɻg�;�Cݽ��H���O=�?<��;v"�>@�5��zG�(/_�p�ν�h
?�A?��n��u�� ���q��x-��Z��~�%?��=s�i��ɥ���q���q�,٧=��G?��/?z���_�������1�>��v>mP����z>9]>1��:)w�d촾n>��ɻ�[�>	�?��l> �=-R�>8����n����>��->�C�>�m8?��?��Ҽ��콀���τ�L�z>��>�<�>� �=��W�6��=� ?�Op>y15��t���J���+<��:`>8���=���6�+C�=��Ƚ݄>���= �D����R�<�~?���'䈿��e���lD?T+?g �=ѝF<��"�D ���H��F�?q�@m�?��	��V�?�?�@�?��K��=}�>
׫>�ξ�L��?��Ž7Ǣ�Ȕ	�))#�jS�?��?��/�Zʋ�>l�6>�^%?��ӾPh�>wx��Z�������u���#=R��>�8H?�V����O�h>��v
?�?�^�੤���ȿ5|v����>W�?���?f�m��A���@����>9��?�gY?roi>�g۾9`Z����>һ@?�R?�>�9���'���?�޶?֯�?Ǯ>���?�O�?Wj�>dռ�mB�tJ���m���_�6�{����>�H�>E<����a�����r���y��)����>�<K\�>�S=�T�����=�\���ם�螳���=y3=>Ql�=;��>�?��n>u��>i�<���<��_��L��\�K?���?����0n�� �<�Ҝ=O�^��(?f>4?\�@�Ͼ齨>��\?�À?d[?�^�>y��?��(濿r��`�<��K>�*�>G�>����<K>��ԾLD��c�>�ʗ>�<��X@ھ�<��)����F�>�[!?*��>��=�s$?'�2?\��>���>!60�����=d��5>�)?_Z?]n�?	!??�Ⱦ��4�Z���p%V�ٳ�=��x?�l?���>�ˇ�m[���~N=���Բ_���?�MM?f�����>T�t?�JD?|�'?:k�>ӊ�������{���>z�?@Cu�W(&����kսB�,?�G?��?�(h�����撁���b��5���?��9?ak
?����~x�b����d=J�]����<I�>�~b>�/�=��;��=�	�� >v����n���{_��S�/�h>��v���˽��Q>�#,?��5�"̃����=��r�e�D���>��K>�׿�w�^?J�=��{�%����p���{T�a�?�{�? N�?����h�z�<?�*�?R?K��>�X��Yi޾cྜvw�ۺx����T�>;��>�<v�Z�侜n�������Y��5�ƽn�� ��>���>��?<A?��>��>BF����*�8����پIc��
	��p=��<�.� �:ӗ��)#���<�̾*��f�m>#�ϼ�>f�?�X}>۽B>���>%�w=y�>y1,>OO}>�p�>`/d>@.�>��l>z=��}��ER?����?�'����௰��3B?�nd?G7�>�ci��������|g?�?�v�?�Rv>xh��%+�cV?��> �� j
?o�9=�+���<E-��ּ��ۆ�m�P��>�R׽w):��	M���f�;Y
?�,?����0�̾�M׽^���D5y=�L�?�m%?��(���X���x���\��@���귓������*�i�r��ƅ��x��@��6�/��<!�%?|^w?q����5F��EQ`�x�D�D`\>~E�>���>;�>�b�>"0��b �>�k�K���Yi�>�Pd?.�>M�F?�nE?��9?%�9?#6�>C��>̂��D�?0�>P�>�O�>�?X�+?�D?��
?�*?�c>!�?=����l�۾_�?+�
?>(?�D$?�6?�6���y5��T�=�K��sþ�.w�l30<��=`(��i�Z�=���=�y?"�ӽ�M-�>��Z��>��L?���>�E�>/���
ԾJ&���/>>n�>$�>��	��k��*�/Q�>Őx?c�	��}�=��G>M��=8�������d�=��$�zB	=�߆�k��<Nb8=J��=��=M}�w����~<Z�=W�>Vj�>��?�p�>&�>�Q��ݤ �+�����=��X>S>QE>=0پ�{��'����g�EWy>�p�?Gy�?l�e=�*�=1��=Lv���3��H��S���<v�?�]#?�HT?���?��=?�^#?��>��.@���S��V����??]?�O�>�)��/��o듿�D��E�?�(?�C��=ھ��1�mJ�W����=F�$�w��N`��;�8�E�=dn��w�/��?&N�?r�;�CX�?�$������¾��X?��>��?�7�>�F���|���2�_�s>G?�nA?��>�� ??>�?�t?���>�6�L ���[��pżn`�>�J?�1�?棃?BE??-K�=]��<�f=��Ⱦ�\��
����Qz�Kف=�#o>��>��?�GY>�%p>��K:Ux��b���9>���>V��>CO�>N�?�d�>:"J�{�G?]�>�ľ�O\������郾�)@��u?��?��+?�=V�7�E�T������>�t�?��?�7*?TS�=h�=c�Լ%嶾c�q�� �>S��>8)�>=̔=��H=�S>���>�i�>����D�C8���M���?�E?�׽=P|ʿF�n�?}�������f�F�̾������	�����k�=\Ҙ������ȯ��j�ˌ�0��"4¾�n��ﻎ��l ?#��==�$>���=<��=z"4��ҥ�z�.=`��R�=7���zH=����U�	��u���c<ڎ�: j��z��j˾ԕ}??I?��+?�C?��y>4�>f�3����>X����A?�'V>�
Q�-����;�5����8��,�ؾFZ׾p�c�M���_O>S�I�ض>T'3>d:�=1^�<��=,�r=`��=*�S��J=<��=h�=V�=��=*�>�D>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�1�=�>�Y�a�I��
����,4����(?�d���^���?8 >�(�tb���=>r���]
>���>�M�e��=��=ܲ=-��=::>i82>R܊=��ͽ�-�=��6�=p�=�5ͽ�񇾝4�J��=T�=�>]3>w?a��>L9;?'[?��>�(|��<���»�v��>�$�>_
?��=��>K�>%��>�-\?�c?%�>���=1�>m[
?QD��Ej��Ͼ���D�p��?�C^?P�>��9>G����c<�#��<j�8?���>�j�>h��>�U����:Y&���.�&���֜4��+=�mr��QU�B���Fm�-�㽱�=�p�>���>��>:Ty>�9>��N>��>��>�6�<wp�=�������<� �����=1�����<�vż�����u&�L�+�1�����;q��;��]<���;��=<��>2�>�K�> M�=�����.>'��MK�97�=k�����A���c�j~�$D.�ޭ5���A>1W>�∽5���	?��\>��A>8=�?h�t?H>T��*׾V���Jf�C�T�VW�=|	>�q;�P;�|�`��JN�.Ҿ���>��~>�c�>�ׄ>8�	�]1&�c�ݼ:Ȩ�^hQ�O�>�1�����3c��`��]��b���n�\���<�*P?�G�����мc?�LT?ZN�?ȶ�>��;�� ���g>�/�/� >-`��_�G�2vI�]J?.W>?�?��Ҿ.C�&sྒ躽��>��/�P�>���/fA�����z������>�]�����Ť)��o������l�E�d�v��A�> k4?�A�?�r�,7��Z�\�U��C���>�!l?&�>3�?�!?k<�:��o���@|=ZYh?,�?�H�?ODs=ʥ4>퍫�?,N-?��?} �?�AG?���N��>�j>h��>P9�����>�$>���/��=�:?� ?�*?C��������)���a���"㽼���>ML�>�g>�׫>��G=k�~>WP>?g�>���>��?���>H��>K��>H��J�0�W#?8�g>G�>@�5?���>r�ƻKܽI�=�ռ����l0^��t=� �;��=Q�>��->�->���>!ǿ3��?7J�>�3-���?"[�����{2>؎�>IXž�>/.>z�>e	?v�>A/ >y�O>G�;���Ӿ>���� ��B��R�!Ҿ��w>˺����)���	�vv���9F�쵾�X�a�i�(5��Z�=�P+�<�}�?AS�"'j�܃(������Y?;2�>��4?�|��pNw�g�>���>�׍>�T��A��������4޾��?���?�;c>��>7�W?�?1��3��uZ��u�j(A�e�&�`�~፿�����
����_?�x?9yA?PS�<:z>I��?��%�Jӏ��)�>�/�';�E@<=�+�>�)����`�W�Ӿ\�þ8��HF>��o?6%�?cY?MTV�ƻ5��>��=?#4?>�s?N�2?�8?497�$l%?5C>g?��
?�9?�/?c?ĝ>��>A�8Na= H��@ꍾ��Խ�ͽ�S�6u�=^�=䬜;V^�<d!�<�턼�(k�б���z<(�e��e�;A�?=[K�=9~�=F:�>�_?N?��>��%?��c���?�RIH���S?��=Q@߽�z����_a����l=�{v?ǌ�?��P?�ͨ>�8P���+���=[X+>�>ݽ�> U�>5nD�y_���=+�y=Ua=��e��g8�M�u��d�C����c�5��>�a�>��|>hǍ��&>����n�x�6�d>��O��湾�SU��?H��X2�aPu�H��>E�K?v?e0�=w@�Hx���e�g(?s0<?�)M?��?���=bܾ�x9��sJ�@y�Q�>�5�<k�G������Ɖ:�`h����s>�����)���c>��
�m_ܾ��n�v�J�&�f�C=y���R=6��P�վ �}��e�=��>�����,!��2��QЪ�&�I?�g=:8��ԨR������x>9K�>p��>h�<��ir��\@�`��꫙=}8�>_�:>�W���N�߅G��(����=�1a?�_?e��?�:ۓ�f?��/	��a���G�au*?��>{b.?���>6�h>'���m$��S���k����>�C�>%<6�\�p������|;��?�g�>Q3��*?�}�>�[�>ί|?N(?�c�>fh�>9XM=����"v?&�?
<>9�������I��mH��??�N8?N�ž���>�Q�>��'?�B?
g?lp ?�4l��?���[�lڣ>~l�>��q��*ſƒ�>�oe?`�K>Cv�?���?T�=#I�UA˾�'���<弔>@0)?�	?�+"?��> �? �p�d��	�>1�?�HH?L�7?�b>��<>��g>�����>�K�>k��='g>�vS?uӃ?�X,?j��=��Q<�H�Nu�<:UY���˼��{�o	ѽ�4�k���k�;>tܽZ�(�S�7�y���;>�;I>F*L�J;��|�U��>�,�>����)}z�حžU��蔟>/�z>�]���Ԧ�TI�=�c[>��}>08?�[>f�y�jn�=Mb�>rV�>���&+5?���>�]�>[�$=�+��������l��=H�M? ׋<Z��J��KK������p?'?�P��w��K�b?��]?5h��=�	�þ|�b����g�O?@�
?<�G���>��~?e�q?W��>��e�*:n�*��Db���j�!Ѷ=^r�>KX�Q�d��?�>m�7?�N�>8�b>,%�=ku۾�w��q��f?��?�?���?+*>}�n�Y4����v둿�^?�l�>b���^"?`}?�&�ξ�k��q捾n��|֪���
���^��xO%��.����ٽ).�=��?�s?Iq?E�_?I� ��wd���]�����sV��~�Ƒ�$=E�0E��CC� o�/�?���d՘�@.T=xK���Q"�%(�?Bc?��V�>���������V���k>Ѩ���~?�<��[�c>��=@�n������־�?�P�>��?�:;?Z�Y�O��6�'A.�p7�����>_}�>tR�>�o�>��1��x��.茶�R��V�� =��x<}��?̲v?Err?�9ξ��d���t���
��>�*ܾD��>���>Õ>آ��g�=`�&�T�f���r�����-����=��q?7�e=�<�`�?<�,>�!*��ỾP���Q�G�G��=t<�>�K\?�q?��>C)��^F�̗�>��l?���>x�>����g!�J|�u�ʽ�B�>SЭ>L��>�!p>H -�1$\��_������+9�(��=�h?�q���`�	��>��Q?�8�:��G<Gn�>�w���!�����'�4X>6y?z�==a;>��ž�/��{�j��)?��?ϔ��;�)�.4�>��!?��>���>�f�?�W�>"�ľ/g9��?�]?�I?��A?&x�>�2"=�\���ZȽ��%�cC+=QT�>�FW> ^r=���=�5��]�	��QWF=ތ�=,輴f���72<�Q��� B<d�<v�3>Q�޿��M�@Ӿ�9���ھx���)��+���p���#	��ų�F����v�������<��D�l?O���HN�#)�?�:�?llپpC���^���^��|��v��>��~��=6�Ӿ��W�������xpȾ���s?�@|R��G�l�&?%钾ٸǿ�桿+I۾�  ?�� ?�Iw?IZ� ���-:��� >}=�c�����з����ο����`?��>xﾬH�����>#Ɓ>r�[>�Au>/����!���;�<#?�^.?h�>�.q�c#ɿ�H���ք<��?�@�-D?�n>��d�j��=6�?�?܁>��L���#��$0�Ъ�=$\�?*]V?д��)H�"�!>�r?ȕm>CG%��ۻ|��=څ >�>+��!Q>s�">���l��}u1����>�p>G��2as������F>��>�� ��<!�1u?�,���8��p%�2����n>��-?*oB>�֜=Y�L?D++�mTؿ*Ձ�E{?o9�?)b�?4�0?�Ӿ7#�>ba���.s?�=2?k�>��G��`���z==z]���>���P�k�>[Z���}���1=��U=�r�aI��6�T��=0��ƿt�$��Q��=/?�IB`�}���<X����?�r���m�q=^��=�Q>��>�lU>	+Z>�NX?+�k?�F�>��>v���m���˾�?K�����%��p��9��鋣��|�R��Z-	�Z2�h2��ȾO!=���=�6R�H���� �K�b�3�F�[�.?}v$>��ʾn�M���-<�pʾ࿪��Ԅ�Xॽ�-̾�1��!n�o͟?w�A? �����V���R�\����W?�R�@��$묾���=���1�=�$�>���=<��` 3�~S��/?tb?�l���Ð�W\,>>��t�V=��.?�9�>T�<�֯>��$?J+�w�dHM>H�6>�}�>�>/ >�먾(�ｴ?K�T?��н�C��EԊ>����Up�z�= I�=�7�'5��D>��<Ϭ{��(�;Y��f�O<R�M?,�->�%�����'���=`lr>�q?��>���=h��?@�"?�;<�兊�/�l��޾�Z>+X?�/?��>�=2�z�ƾ̜����g?/�-?0��<��G��@������z���=�>�^i?��o?��>l长ޝ�� ���V?��o?`[�M웿�sྜ!&�Q��>�>5��>�s=�록>�#?�����ۑ��"���x:�7Z�?�$@���?�M��P���(�=��>3y�>�y�����,��%d���Y=�e�>�\U��de���6�`�(�@
?�>l?���>@�,���3��=dw���J�?Ux�?d'���F��/��>nc�����D6=��=����H��2�@�/��ɾ7�d����;9�>�@��ӽT��>�&6��8⿙�ʿ����=Ӿ��b��?��>o����g����n�<�{��H���E�m�i�	�>�o>�5�����~|��<����kV�>e��.��>�=L��Z��EƜ����<8*�>hO�>� �>y���o����?
	����οѶ�����=�Y?U�?�Y�?�?��;VHx�����S.B�i�F?��s?uY?]�*�c�W���7���j?�Q���M`�א4�nAE��JU>%3?�Y�>�-�[�{=HY>B��>�v>�/���Ŀ�ն��������?���?jj�t��>�x�?6j+?8g��9��M���*���G��6A?2>�����!��:=�MԒ�׾
?n�0?���1�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>hH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?��>�#�?���=��>`��=S���+�.�>c��=�A��]?W_M?��>V��=��5�O�.�~�F���R�o��MC�A>�>ha?hM?:`>����(�-�!��ν/�P��1�?�g�"�����4>�U?>��>}�F�#Ӿ��?�3���Ϳ"|���5����M?@?b'>>�6�G!�>����xE?���>�2�����v���5S�9u�?g�?4�?2A�J��<�9�>�@�>~@�>i��9o�<����Y)L?R��=G�����S�DV�>9��?M5�?۴�?A}��	?M�iH���Y~��p��6��Q�=�7?M��z>���>�0�=�_v�Y�����s�׫�>6=�?cm�?���>�l?B�o�x�B�
�3=[v�>��k?�Y?��y����H�B>n�?��E󎿇P�jf?&�
@�o@ɕ^?�袿4��ȃ���Ѣ��+��!��<�	X� %>(
��8ڻ���i�a�&�Ľ~�3>�m�>��{>;��>q�8>oP#>��I>4����%�ޥ�T���*�7��<�����:����A�g���"��X�o}��ö��^��o�<e��f�	�L ��`�<��_?�f?�c�?�5s>�|����H>�%�>�>M�%��?k=��>��@?Z�@?_7?��5=(^Ҿ��ڌ��׵��qnz����>�B�>��>wm�>��>z���n>RE*>H!�>��>�>�x==᫒��w>#i�>���>���>�C<>��>Eϴ��1��k�h��
w�w̽1�?}���T�J��1���9��Ҧ���h�=Ib.?|>���?пf����2H?%���z)���+���>~�0?�cW?$�>��|�T�/:>:����j�2`>�+ �|l���)��%Q>vl?}�f>�u>�3��`8���P�@w��'|>�86?!Ҷ��D9��u���H�mfݾ!+M>پ>N~C��f�3�����bi��>{=E�:?��?vu���䰾�u��5���LR>��\>Qg=���=�sM>ǚc�;�ƽ�.H�?.=���=��^>N�?�=۞j=�^�>$}�᩵�@%�>F�[>U,>Tq+?��?�9=B����C���������>+?:�{>Zn$<���%��r�>
S>�����<��@�cc��Ys|>�R&=��~�>GA��2*��M@�R �>��>���;ʌ���Q=�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>�g�/���j���ZV�b��=n��>��?X�#���>vھ�)�>�t?�����1���Ŀ�Bw�{$�>�7�?���?�V�ߘ��yO/���>���?�d?ܤw>�裾S(�(�6>ފ\?�7a?�>)+�䎘�M��>��?�@�?�!A=�u�?3��?��>�C���"K��V̿�.Z��H�>����j�m>�;�>�Ѿ�UE���j������
���P��1�>�`&=9o�>�|H�E"̾���<F.K=S^��⢽�r�>��(>o�>_��>�T2?&�>yA�>I�=�sj��>������w�K?���?$���2n�dN�<^��=��^��&?`I4?|j[�/�Ͼ�ը>ͺ\?_?�[?�c�>"��=>��3迿!~��K��<[�K>14�>�H�>x%��FK>��Ծ 5D��p�>�ϗ>�����?ھ%-���W��|B�>�e!?���>Ү= � ?b�#?�k>�7�>gbE�$<���F����>n��>�<?��~?�?����'^3�����l顿F�[�/�M>��x?zP?_͕>�����~���>D�d6I������?*�g?�'�(�?�8�?�??��A?�e>��
%ؾ�Ȯ�:*�>��"?����<�Hi!���	�:U?%?���>�>�������Ӽ���pC��k(?p'^?�0-?�����\��j¾܂�<�
��M����f�R�7�$>�}>����y��=S�)>�F�=�$��,�U����;�)�=�>���=�C�J�T��?��>:���e�z��!@���=XZ	=G\���b?/���5��|@Ŀ�S��u��=���?�"�?6n?��@��Bv�F�Z?[�?K?ZI?����������{�ɿ���c ���v>z��>'ަ�4.+�\4���!���n}�#���Vzg���?���>�<?���>���=�܌>Ӿ
Q
�)-��徟�f��i5�bP;�F��UB���������P��*�̾�᩾�O�>��`�X^�>��?���>7��>~)�>��܌>c�!>��X>Om�>,3z>�NA>Ш�=B��=�9Q�dsP?�̷���#��Y���F?�c?���>��g������"?�^�?Wӛ?%�n>	�h��'���? `?�����?��3=�In�]�M�g�ľ����*��<6�r�>�D��2r2�b�M�=���4?�?���<P�׾+B �������1>"{�?�	.?T�3�A�_�����}�3���$�d�==ZU���q�S61���k�"4r�M͆���~�2!1�_E=N"?��?B�9Ǽ��8��eml���'�kM�=��>"y >{5�>z4�>Co�s$�r	g�^E�����v{>Ɏ?��>J7I?K�;?ԅP?�bL?X׎>uR�>v����u�>��;mҠ>���>�\9?ig-?L20?N�?�+?�c>����L���Khؾ�?�K?��?�C?ES?�y��[�½����k��{��À=���<"�ԽJv���N=�MT>i�!?��|�$�"���$���?QtA?`�>n�.?�H+��þF�>ˌH>�k?ǺF?�n�շv�|n&��?��?d�G�@�>Ao>�b:y2�#�=FΚ=��}�Kh�<�g�Î���>ŕ�=�������=���;���sGZ�붤=?e��>d+�=�>����?�w��P��eл��g=x|C=yE>ᮾĎ�ic%��F�>9i�?C�?ߘ�2��=Y�X>խ�8���n�ᾃ����,>M]?��?P�1?�ߡ?�(?�?6��>w}�]X���de���f��_?s!,?	��>�����ʾ��։3�֝?i[?�<a����;)�ݐ¾��Խͱ>�[/�g/~����?D�4���T��6��?�?lA�W�6��x�ڿ���[��~�C?"�>Y�>��>T�)�}�g�s%��1;>���>jR?u�>�P?3m{?y�[?�Q>y�8����љ�	��Ր!>��??3��?��?+�x?���>[�>Wd+���ྷ������f��c���^`[=5zY>6Q�>V�>���>�<�=��Ƚy쮽Ү>��s�=šc>`�>��>��>eUw>�s�<e�G?V�>Z¾tq�	E��2m��e$� �j?��?ߜ)?ù�<A�DC���ƾ>��?��?V�)?;�_���==��� �����s�W��>r��>�|�>�X=�H1=�v>D3�>�v�>�09�QW�� 7�O��?	nD?,T�=�ſ�q�Fq�������h<�����d��ʔ�P.[�c��=5Ҙ�\��婩�}�[�����em���׵�!���&�{���>�n�=���=�=�)�<�ɼ��<�J=���<7�=��o��hl<�]9���л�������p\<�mI=
9��=�˾׷}?�=I?��+?�qC?��x>�>�9��>鿅�+?OeT>8�X�ų��,;�`��90��mEپ²׾.Md�'j���>ruI��m>��3>���=�]�<���=b�m=pR�= Wr��5=�l�=��=kg�=U~�=�>ϊ>nYv?��}�o���8J�~�I�<?��>=W�=����M@?8�<>�����Ƕ����4��?9��?�?��?�k���>�k��ɒ�l=����j�<>�¯=8�<�Sߪ>��Y>���ट�p���=g�?�@h�>?�+��.4Ϳ�L?>�M_>�K�=�jO��Y'�����<���+�?Rh>��귾�i>���=s�ƾ�!Ѿ�'����[>_�>�t���oT�܏=􄄽P�@=�ڹ=��>�b<>��=�xӽb�=2&�=F]�=(,->A�J���k��Z!���=��>�{d>�T	>s�>�X?�Y-?4`?J[�>�GO�tW̾�ľ�y�>a��=E��>��-=�D/>��>��;?�qK?�L?,�>Vo=��>?��>��)�hXo������̞�=<m<���?�N�?�.�>�߄<�hk���#�h;��5��ކ?}�+?�0 ?�ߤ>��6&忲������G�DB�'�K=�B���N�����y^�P����?>�1�>�)�>Ѿ�>l2S>Q�T>[S>��>
�=	���ŭ�=96H=�֐=�E=OL?=5��<�YX=/5=iv��9.��Jݽ��T��*������e<�����7=�?��e>ԛ�>8L:=�,Ӿ�EQ;���u�I�<=X}����L�W�x�t퇿�~�{� ���>>EI=�(A�aR��f(?�^>ҍ>�}�?�c?Y5b>U\0��v
�ȳ���.<�����P>i�n>��n K���q�1�i����^��>`ߎ>�>1�l>�,�7#?�r�w=�[b5�r�>�|����3)��9q�@������Ui��RҺ�D?�F�����=\"~?�I?a�?Í�>B��ؾ;0>�H��<�=b��*q�1i����?-'?&��>�쾨�D��H̾���޷>�@I��O���2�0�լ�^ͷ�*��>������оh$3��g������ӍB��Lr�N��>�O?��?�:b��W��,UO�����'���q?�|g?��>�J?�@?&���y�r��v�=�n?���?I=�?}>6��=�ý>��>{�
?L�?ϝ�?f#l?�C�>��>6��<bw>�T��c9�=:��=�=��!>f�?c�??�������A��g���!}�=�.b=�z>t�w>O�{>p�=�J��w9:=�@Q>?��>'��>��P>�4�>�2�>l���3����?�W�=1�S>� ?u\>�xo>(��{g�X��;L����J���3#���Z<d��=��=�9B�b�=����>-�ٿ���?H��>"��*S?Y�2�?TF>�W�>o��>lt��s�	?g@�>�t^=:��>��>���>��>J�;`��Un�<���%�/��n#��5�6`���=����=�� �_(��3)�Djw�������V�#�f��9%���=�ͫ?}󙽎��Cq9��/	���?Cq?�?�پޑ>3���<?�t�>������攖�#����?���?��c>5��>�W?�}?d1�	�1��BZ�	�u���@�n�d�`�`�,ҍ������
�+S��I`?n�x?KA?2\�<B�y>䌀?��%�aO����>��.���:���:=T��>fҰ��A`��DԾ�Wľ6@�P/F>no?~��?�?�mU�|�l�>�&>{�:?ғ1?f^t?��1?�;?p����$?�v3>�"?np?�T5? �.?��
?�:2>Ȅ�=È���'=,6��B抾�ѽDdʽ���W4=*N{=����	<Nb=�3�<���}�ۼp�;v��iѫ<��9=Ԣ=�=D3�>K�[?��>l@�>�7?d	��J7��W��.?��B=�Ɓ�/)��E��s��z�>l?�ë?�Y?Y`>��A� `A�,�>Dy�>�/>	P`>tN�>�����G�	Ռ=�T>�>.��=�K�ǭ}������V��<d�!>��>o�>?�F�0R>;���Ɋ����B>�l��d��c�-��K�x�;��N����>��U?ߡ"?~�=����ǽ��i���0?��@?�tK?��?,�<�m�;���;�׈>�u��>�pN=Yo�C���֥��B��a����V>J����ҡ���k>F���Oھ�Kp�uJ�8D��)=�H	�A*@=y�	�q�Ѿ)F|��R�=�>�ż��>!��m���(��\*I?�Kc=t*��W�T��W��N�>�Ɨ>�+�>`�I���H��j>�1�����=�c�>x�<>��%�Đ�"�E�����4>��T?�/�?6v?�2־Ot��L/�'[��뗽��L�?��>a��>M��>#ڄ>����:�-숿�_����>�b�>�\%��06������޾q��ku\>v5�>�>^v�>b$?�\'?mZ?�$?
�?-׌>�Kǽ�4޾T7&?j��?H}�=K�Խ+U�*9�^F����>�)?L�B����>W�?b�?X�&?K�Q?��?į>�� �+Q@�˗�>�R�>e�W�}Y����_>��J?���>�1Y?�ʃ?%>>{5����M���^�=^
>��2?1#?8�?���>�_?������t�>k�?�O?�<)?��J>x2�>DZ�=��>�$K�
��>9��>�zt>s�.?M~?��R?���>$ ;L�1�����Q���8B���սkܼ|�<��~�c�ν�a���@�j�\�*/��f�����=i0j=�߼��F#����>)�>Si����1>>����߽2i�>>�b���U�D���-=Ԃ�=���>�I?�"f>�!����=���>X"�>������)?3��>�3?Y@�=抈�*pڽK�`�qѱ>=9M?
=<��ۙ�C�n�K7�=D�[?G}�?�k��*��N�b?��]?=h��=��þx�b����f�O?>�
?7�G���>��~?e�q?V��>�e�+:n�*��Db���j�%Ѷ=\r�>KX�R�d��?�>n�7?�N�>/�b>-%�=hu۾�w��q��h?��?�?���?+*>��n�Y4�X��J��5�]?��>y����"?�����ϾrI�������@��7���u-���w����$�̺����ֽ�ļ=�?"	s?�Kq?��_?A� �Ed�+,^�"��L[V�<'��'�O�E�� E�Y�C�&�n��K�����_8����F=ř��+���?��0?�Jj��;�>���i�ɾ��ȾU�@=DL����-�	;�=�����p>�#>��C���E�w���54?٧�>���>'�"?M�d��B�v�=�̹5�cRݾY>�e�>�>�q�>"F��o��8.���۾v��q����=X��?�^�?�ZZ?j�˾CN�Wn����b�>9�ھ�9�>���>�Ƥ�q>ݾ^��=N�:���M��΍����,����"�m>_�@?V�>��>�W�?C��>�^��);8�Ͼ��Ծ��>W?4B?���>^�>�H�	���'�>�m?���>�)�>����f�!��l|�lDȽ��>�+�>���>��o>�r.�-x\���O���)T9���="h?'��(b�nt�>`HR?&ⷺ߂h<}��>(6q�i�!�q��*�%��	>ۘ?��==>�=žT���z�������)?�e?6���ގ'����>�p"?�J�>���>J��?��>1�þ�����?�o]?m-F?%p??��>�X=��j�Ž܃%���=7�>�@V>�A=MG�=n���[�ϳ#�i�*=��=�)ּ��ؽ���:���V��<�ï</�)>Y5ڿ�wL����t�"�P6쾈c��@mk�Yx8��¸���M����Qo��FB�����}�=r��RGJ�ɶ�������?K�?�b��.žAR����[�𬚾��>a�оvt>Q�뾃C� �K�Y&ؾ�"Ͼp�8�rC�Y�g�S-��q"?�ľT��g欿�u羴�/?*C?<�0?o�$�qt���~�Ry�>��;>B��=��$�6����¿-����a�?�?ڣ��B�=��>��>�d>Z�>����Ρ	�O���ǫ>��b?_��>uɹb�ȿ�����)�e��?(� @]�B?�(�p�����;>Ld?/�>�nZ>��^����վ�=�>S�?�b?gR2��jQ����=V��?���=�33�hDs��y>�W�=�TD��E<�i�>9��>F�`�K�,���=�w�>#��>����Z�׼FyC�����ɵ�=_����=5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�j���ÿ�����#�V��<t"�;�n�N�3�@������J����Ck��4�W�r=�)%>>�s>:�{>B"B>@�'>�G_?�Td?�>�!�=M�ý(t��Ʋ�2���W��@)̽�ۘ��� ��E���� Ҿ����G���
��S���F=���=z,R�"���b� �b�b�*vF��.?�#>G�ʾǴM��e)<�tʾ���+~������̾�1��n���?�A?|��W���� �� �����W?���4[�DF�����=rή��=�̜>t��=O��T3�.S���.?��?VE���s�͏,>�[�a�=�+%?�$ ?�G=%�>��'?[��?��G+N>�;>�S�>x��><��=>%����ϽX?fHY?ɋн%���q�>�;��ǿZ��!�=�8�=9@��,���4>MP
;Mm�7^�=��� Q���+W?� �>�)����±��J����==3�x?S'?ߟ>Ok?�B?Je�<�>��b�S�8�
�v�z=*�W?.i?�`>mʀ�9�Ͼ$��I5?9`e?�N>�h�-��:�.�x^���?�un?�+?)��yM}��������G6?�v?�K^�6D��WM���T�v�>��>���>W�9����>��=?qy#��𔿗����v4�H��?�@l9�?̖<�!���=�?���>�P�ͥž./���ڵ�lCo=[��>���͍u����zv.��f8?�m�?n'�>Pp��#��I�<�r9�o��?*�?P�ᾒ��S�)��^�]���jȽqĦ==𭽢��p�w?���l��M����5���A�>�@@����-�>��3�5t�轿X����ms��ޅ�]?\q>&6ɾ���������C���U�:�G��
���>}�>j���T���U{�ذ:�A���#.�>�J���>��U��������+<��>O�>3G�>%r��Q��蒚?h��عο�ݞ��"�o�X?u��?Մ�?O�?G��< }��}��-��nRF?]q?"�W?�?1���`�E&�&j?e���)1`�~�6��E���Z>c4?s��>��-��O�=K��=���>Ȋ>�H*���ſз�ne �ף�?*#�?���j�>q�?�)?w���y���᭾MR)�Y���'�:?J�4>�;ƾ�@!�CH;��C
?\/?Q��_��]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?� �>R�?{��=�a�>�L�=r����f-�4j#>[<�=?�K�?�M?�E�>jL�=2�8��/��[F��IR��$���C�q�>Z�a? �L?Gb>�����1�X!��pͽ.d1�Ru�.S@��,�-�߽�*5>�=>q>��D�_ӾY*?�5��7¿�;���HٽY�6?~ؐ>��>z9��~3��ۼ��D<?��>>���m4��k���Ӄ��Ȥ?��?:��>�)���ep<*U�>��-?M��>t����=y�"�x�F>�:h?S���t�c�|ZM��<?�'�?$9�?�:�?룃��	?���P��*a~�ł�� 7�]��=��7?�0�$�z>���>��=�nv�����<�s����>�B�?�{�?��>��l?t�o�%�B�#�1=}M�>��k?�s?�2o�-�)�B>��?3�������K��f?��
@zu@C�^?0&'࿞���I˲�t���;D�8�J�#�5>���:������>�=΃L=�M>N-�>@c>�.�>}{$>YxY=A��=e6����(�$J��K���I<������� B���A��dV���]K��0���E4��1w����B�V���F�p�J�Q��=[hV?kzS?bqo?�H�>������>L����#=O�#�I�=�~�>d�1?D�L?�(,?oF�=pӞ�!=g��������4���?�>�KH>���>��>��>�:��C>��C>�1�>���=W�M=m��:H=�4S>x��>�)�>�η>�C<>��>Fϴ��1��k�h��
w�n̽1�?����R�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)���+���>}�0?�cW?�>!��l�T�1:>7����j�6`>�+ ��l���)��%Q>xl?��f>�u>��3�Xe8�p�P�{|���i|>�36?E鶾�D9���u���H�^cݾTHM>ž>_D��k�r������ui�u�{=`x:?Є?�7���ⰾx�u��C��{PR>�:\>�U=�i�=�XM>0cc�2�ƽ1H�ag.=U��=��^>�$
?��f>�����?_'�tՈ�H�?���>�Rk>��=?D"?�@X>Mg8�!��������>�L?�{r>f�ڽ��&��[<�ޭ>Ey%>&�'�H��J�����.�= ���#1���M�2@Խ�����o<�!�>�=>wH�m�!��~?;~��J㈿���K��,oD?�(?��=`pF<��"�����F���?��@ll�?0�	��V���?�@�?3
�����=�y�>
ի>�ξ��L��?(�ŽUȢ���	��'#�`P�?�
�?�/��ɋ��l�5>f]%?��Ӿ��>�!��ؙ������q���v=�>�[??O��3#=|~s�V�?cw?,v�e����ȿ�v��x�>�M�?��?{}k��ܕ���7�4��>]�?ٔX?�JY>��Ⱦ�w^�
n>>]L?XU?�a�>��!��qU�\�?��?���?f+=���?���?�z">1����u��ÿVHR���?�C�\ ?:ၼ����1r�ǫ_�}щ�a�m���U��6
>:U�=<��>f�Ľ�Ծ�	=���=������="�>̼!>5�>���>!F?�>u�>�뽽�������`x�k�K?���?���2n��J�<.��=��^��&?�I4?�f[��Ͼ�ը>ݺ\?g?�[?d�>,��>>��4迿~��k��<
�K>M4�>sH�>V&�� GK>��Ծ�4D��p�>�ϗ>�����?ھ-��}S��^B�>�e!?i��>�Ѯ=ߘ ?��#?Q�j>}'�>�`E�::��J�E�ձ�>��>5H?/�~?i�?�ֹ�V[3�L���桿��[��6N>��x?�U?<˕>e���/����#E��=I�����4��?�tg?�T�Y?2�?'�??��A?&'f>v��?ؾ������>:�!? L��SA�4n%�����E	?+?��>!͔���սf�ʼ��g��,`?�"Z?v%?��K�]�"���/�<��	�����E�2<Jqj�[�>�>���h��=�>���=֟k�I�8��F3<}۷=¸�>���=մ8��X��j	?��`>Q���p>$b���9���>�j/�Z�i��U?ZD6��d��yo���F��R?���?DI�?��h?�ɾ��u�'�U?]��?�D?�?>J;�c���A��e >�����þ�vZ=���K*ὂ����搿�^��Mń����@���?�	�>5?7��>�� >%��>���������	�zs��B�T�����6���)�~�����EF��ý$迾�^���>�>J:��3o�>�b	?�
+>pJ�>�t�>F�Q��`�>uL>%�>���>�%�>�Q>��>�O==?�IR?JBҾ�'���𾁺���E?�FZ?r�>M�����t����@x?��?���?2�*>�g�F�%��?֜?��d���>IsX=�E"= �=3����e+��� ��ml;��w>*|#��D�\�E��]��??��?���=�C��!<������xb>.a�?�$?;>2�W4x�{���M����eY����K�J[O�>́��#v�'�y�l�{���.��km��� ?��?)�#���!���⽔st��?��p>�?�H�>�i�>�� >�r��u'�0^p��:��С���>Lނ?f4�>�fI?V�:?�P?t�K?a��>�/�>(������>��B<��>���>��8?;G-?�L/?b?�,?��c>	f��j���*rؾ2�?�?t?U9 ??jM���u����ov��'y�ަ��ڱs=�<L;ͽ~�K�ǍD=�QN>�f ?[���7>�Rd�ұ?Qq?G�2;��??���S�Y��7�����YI?�'?���JV"������.?"ˀ?��a��0�=v�H=�C =W�!�Ş>�Q�<�G8�1��=�-s�c�?=�۽���!>Э%>��;i�+=�ýޞ>�1����>ɸ?�R�>�^�>�Ʌ��� �\���6�=K�X>�^R>��>�Gپ~i�������g���y>�|�?�n�?>�e=� �=9�=Af��@C�����k½�<��<*�?O,#?�HT?��?_�=?�M#?A9>���E��SU���&���?n!,?�>)��]�ʾ-�̆3��?$Y?�<a�Ų�<?)���¾��Խ;�>R_/��1~�����D�N჻��������?;�?�A�H�6��z辳����Y����C?9!�>�T�>w�>^�)��g�S$�1;>!��>�R?N�>i R?t�~?+�Y?3u(>�M:��"��l���1�<�)#>�}>?�`~?�Ѝ?{wy?�+�>��'>�l5�
���2��𼪝ｕB����e=>�I>��>�a�>}�>�p�=~p���E���G����=�Ub>{��>�P�>+��>8gw>�	*< �F?4%�>�������z���L����(��r?�?R�)?9�J=�4�y�C�!���훬>=��?�ή?
2&?K�k����=ޛ����/w�Cz�>+е>]�>�φ=�2�<�J>d޽>�%�>P������v3��xμ��?��??�Ē=�ƿmvr�Oq�����e%<����%�c���o�a��ɦ=��������W��c�Y�E�z��+�� J��m�|�z��>���=���=�-�=Z>�<CO��͹<}�=m�<j�=q�u�5Y<��4������у��໺�Mz<�jT=Rڂ�w�˾m�}?�=I?�+?޿C?]�y>�:>�3��>>���/@?=V>��P�ʇ����;�¬���!���ؾ�x׾ �c�ʟ�OH>_zI���>r83>�L�=DW�<>$�=�s=ｎ=�~R��(=�8�='T�=�n�=0��=�>LN>�6w?Y���
����4Q�Z罠�:?�8�>B{�=��ƾ\@?\�>>�2������zb��-?���?�T�?@�?Iti��d�>?���㎽�q�=����=2>���=S�2�E��>��J>����J��U����4�?��@��??�ዿ͢Ͽ^a/>e�f>�n4=�QQ�����p��gN�V�j�x�?�Q6���V/<>T�X<��ľ�l־����&j>�>Rv��c�W����=�q��D�<�v�=��>u�=>Y��=tS����B="j���>�#y>�ؼg� ����(�=�E�=j�,>f3>�>j�?�.?;be?]v�>Ko�RȾ�]�����>t��=-a�>4�=//>>OԶ>��5?�D?�[M?�>��=sƹ>���>p�+�z3j���V��Ȟ<�K�?��?0��>�Uc<dxA�I���h>�DwϽ�|?g3?�
?��>m=�jgۿr�*������J8�-��;1���UX��s����'���>4x�>I�>���>\&>e�=#;$>�H�>Ҿ�=�t�7�r=X\�=�K>)�E��\+��@�<A���bu4�s�H�<uŽT��"}=����ûi��=��:GS<�)?M6�>�?�V��X�޾Ami>���
�D�="qC��+��"����,'��0Ľ_uX>�*�=9]g�x9��܄�>�^->d�I>���?P�k?b�=�5�b�z����}B�VM����g>�ۣ>�:��X�W�Dw�>,Y�}Y����>�܎>�>:�l>�,��!?���w={�Hb5���>�~�����%��7q��?�������i���Ϻ.�D?�E�����=�!~?.�I?��?!��>���̓ؾ<0>=H��A�=��)q�5h����?�'?��>!�R�D��H̾����޷>�@I�/�O���O�0���'ͷ���>������оp$3��g�������B��Lr�G��>�O?��?�:b��W��EUO����>(���q?�|g?�>�J?�@?K&���y�nr��Dw�=�n?ǳ�?R=�?�>k�=�s�?�>�:?8��?X�?(�k?w�-�fU�>�k���>����t��=��>�&b=QB�=
?��?a?������������X�w0�<�̪=�Z�>�>�q>!��=�,Z=>&�=��H>ea�>���>#>q>��>��>&�۾�޵�eb=?Fښ>G3>���>��.>��K=�ݶ��y�2M���C��gc�Y⌽�"�=@0>�a7=U�B����'��>��Ϳ�Ǡ?��=���?�:�O�Q>cn�=HH>����T8�>91�>�%�>�?��>bK&>�v�> bk>J�ӾS�<=Ǜ$���R�<�4��x-���s�va6>�A���L>��$�ت���3��󧾕*��]��-r�E@�C�k=��?fh���5~�/�꽔�"?�C?�P/?
C���xT>|�ѽ��?D�>@��}��y!�����qh?�
@��c>%��>��W?ؘ?^�0���2�%cZ��u�A���d��`��卿 ��y�
������_?�y?a�A?�Z�<�z>��?z�%������>/��;�=�;=�>z`���a�	jӾ��þ���F>�o?g�?$7?$kV�g#k���&>1s:?�j1?�_t?O12?�-;?K,�y�$?.3>!?�p?Ji5?�/?�?�D1>�\�=��Đ+=l_��t�����ѽ?vʽc����6=��{=��h�<C�=`�<�c�Լ��;����V6�<%$9=�m�=Zr�=P4�>:�Z?���>��>t|6?5#�Cl1��t���q-?J�L=�x�����}g��������=Em?��?��W?��P>�3@��{A�q>s!�>�y>[�\>���>h��P���|=LN>߳>D7�=��b�<����2��-��>��<�C><��>m,|>&��8�'>Mz��0,z���d>D�Q��Ⱥ���S�C�G�&�1���v��S�>@�K?��?x��=UX�<��gGf��/)?d]<?�MM?��?[�=v�۾<�9�@�J��>���>���<=������!��&�:��S�:D�s>A4������"e>B	�A�ܾ��o��"I������e=���޼O=�	�8ZԾq=z��,�=��>�:���� �.'���	�� �I?T�g=������T�̺���>��>��>�=� �k���>�9���Kh�=���>SD;>󘝼6:�_�F�$��Y\>�7K?�qw?�u?8qԾ�[\�}�7����f7�=7�]6#?�b�>Th?��r>]'j>=f��_��eRs���g�"8�>=y�>y�0��A�I������T�4-�>���>��0>�?K	8?b�?�/^?��?���>z$�>	0ԽB-��~�%?���?٤�=�Yӽ76X�>�8���E�2U�>�)?Z�B����>1�??�?�'?��Q?ey?�%>�7�q�@����>N�>�X�	&��+u^>�J?�ʳ>AY?�m�?d>>��4�wآ��������=�'>��2?
�"?-@?i��>��?��վ��O��+?g ?1z�?��c?��>5�>׌�>�PI>KS�>�4->�4>i�= �8?n�y?kCV?8�n>L�R��=_�&���Ľk�><E�r=�GT��z>\��r�3��ӈ<gh��>{;g��=ԣ�}� ��<B��\=�2�>дI>Y���=)>#�����f��l>R��=�ܿ��&J��ýڅ�N�>+�>��>�Wܽ�\>���>�,�>���R��>O%?��.?+��X)^�OZ��Q��Q�d>��0?���E0�VɆ��ޖ���y=��?�I�?ǔҽ�+�&�b?�]?�g��=�?�þ�b�7��:�O?_�
?��G�q�>��~?Y�q?��>��e�):n�-��$Db���j�Ѷ=r�>X� �d�+?�>[�7?�N�>��b>�#�=su۾��w�6q��Q?��?�?���?W+*>[�n�W4��\��OG��R�^?>.�>Dʩ��!?F�<��ξ󁉾ؠ��?Bݾ=歾���b���5+���"��Z��+D߽j�=r?Bpt?�Xr?Ӗ`?�R��VAe�_�]��c��=U�H*�p���E���E�Y�D�[
o����w#��s���4�O=�L���2�}�?z�!?ҁ�a��>o���{оV۰�>�2>R<A��_�>�~H�8F>��=-@s�^\�.޾�o?���>ݧ�>�}H??'K�3�I�Ӎ%�I�'�qp⾺8S>�\�>��e>mV�>+���U>�{���ѾYꅾ����	>�l?�?Q>H?���/�H������;�N�>��T�>���>&�>�����=b��E\�.ԛ�,�셞����� %>��@?`c>Vy�>�ұ?��.?������)�ؾ�(�y�<�
 ?�>i?�?��>����h�E2�>�m?���>TB�>^+��<�!�֑|�,�̽���>`�>�i�>ϡp>��+��Q\�z&���|��R{9����=�h?���h�a�C�>#�Q?�򂺈�U<@.�>.�o���!�1)��3%��>�?z{�=�/=>��ľ���>i{��6���O)?�@?����5�*���~>)"?8n�>*d�>��?��>�¾�ʌ�v�?�^?w$J?�A? �>��=������ǽ�''�� ,=ĭ�>�>[>��k=7�=�X���\�����D=h��=<�ϼOg���<����%�Y<j�<C}3>�ؿ�iH�3\ѾQ$����>@�q2Z��q� ��}�ὑŭ��C��#�9�L���!7��0~P�Q�L����l�]�<m�?���?q_�v�7Y��i�e��+��#��>� ��I^�=�������e�afҾ�Zþ�Y�>�<�N�Q��[F�`\'?륑�%�ǿe����ܾ� ?�� ?�x?���%� �fY9�aq">C\�<�����X�S����ο���Na_?��>�`�:[��}�>���>�Y>�r>�2��p'���,�<$�?�.?�3�>7r�b�ɿ�r���T�<��?��@��L?E�H�?�ai?>?�]�>�#o>������޾fT��擵=Yd�?�K?̌O�b2���>�s�?�ɀ>��C��46<�u#>��
>&#�=�p�+�>#�>�����0=���dz`>���>6�׽b�>5�� w��#�=bd��$0>�6�?��Q�94^���-��
���@>P?w֤>Vܤ=��,?B�;�Y�Ϳ8�g�
P?���?���?��*?�R����>�t��W?AA?��f>RS,��gt�ji�=j+�?F=�>ܾ��S��
�=q�>�+> ��|��6X�	T/��²=���TW¿��G�������S>K� �ؽC[����!�M���i�d�%}���H�=@�>~	J>�e>�+@>E�c>ʦS?/Kj?�>���=c\�w$I��WžI"���ś�Ov�tx�R��t��[��Ģ߾��c\�����0Ѿ�)=��Ǎ=/R����� ���b��F���.?�\$>}�ʾq�M��,<f\ʾ#���$r��Q楽P#̾Ǒ1��n�Fџ?��A?= ����V�����������W?u��s��~𬾘$�=&W��:�=��>�n�=b�⾅3�ZmS�O�0?Q�?]��r{���G6> ����\=��,?3d�>�p<�k�>�� ?�{�YڽW*Y>.�.>ă�>6��>B�>񱫾��l?>U? ���� �����>�޾��}���`=���=033�7����@>\S�<ٔ���a)<�&����;�	V?�-A>��1���������=�8�=�?k?1e�>�4�>fT?]�.?���=5�Ͼ"%=�QI�;�=rbS?Am]?�=t$����޾� ؾ��J?��Y?�(�=A��:|��^���g;���>�_?��@?��=�ы�=㥿\�����S?^�o?o��w��3�׽Ց>5�.>A�?p}�>�~V�9�>���>j��=�lD�����Xi��W�?X��?b��?|�T�]���a�:Y�>�� ?�,i<j �������#��>��?!��l+��K�v2վ��?u��?\?)�)^���U= 	��m�?}9�?�B׾�b��B!��S�);�����I>��g�6�|����{A�ݒ���
�C�ľTνNQ}>��@��</��>V^��y���Pοك�����JKp�%a�>.[�>�ǲ��*��*:��r�u�u�9��C7��罚T�>հ>?Ɣ�0V��6�{�\3;��G���w�>���>�S�$��|���w�=</ߒ>�s�>b��>4��彾;�?����^οϵ����
�X?�}�?�*�?��?Vh<�w�h�y��U��F?�s?��Y?A�&��T\�1�.��j?N`���U`���4��GE��U>N#3?�B�>��-���|=� >���>�f>B#/�k�Ŀ�ض����2��?X��?Ln����>ǀ�?\t+?�g�8��v\����*�ؗ*�s<A?�2>����l�!��0=�Jђ���
?0?�y��.�]�_?*�a�N�p���-�i�ƽ�ۡ>��0��e\�WN�����Xe����@y����?K^�?f�?ӵ�� #�g6%?�>c����8ǾP�<���>�(�>�)N>JH_���u>����:��h	>���?�~�?Rj?��������U>�}?(�>��?�a�=�i�>b��=T���M^.�/�#>���=�	@�b�?��M?=S�>���=E�8��/�S^F��YR�	=�O�C���>��a?TyL?�gb>]���_1��� �`ͽ�>1����@���,���߽�5>*�=>&Q>�ID�+Ӿt�?j5"��sǿ�՞��x{���_?fk?���>��N������=w�x?s�A>]�۾����|�h�뼎��?q��?�C??#��ա<�b�>@��>�l�>�6��TJ�<)����k���t?;-`�̎����j�M>���?:9@Ѿ�?z�:�	?U&��0��m}��/���#���>p+6?2���l>HU�>o'�=51t��I��$�u��f�>�į?���?>��>nk?=eo� �A�y��=R۬>E�f?M�?��;����D>+?D���Ռ�N����d?��
@�@�\?�o��35ڿ������i?¾\�=��0=�e>�h��2��=������ὣ5��L�G=�ɾ>��>t[G>C�=��=tO>���sH"�#���������?��[����D<�/�"��eƾ���� �l�s���Jy���2���6�A����;��=3`_?�
�?�lg?��Q>�Cٽ/ej={�j��y>�R��d�<���>s�$?�??:�C?���=Q¾�5������߅�������j>-
>���>?��>6_�>�v=�z�=[o�>3�>�њ=��I< �e��̜<�X#>�]�>e�*?�w>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?%���z)���+���>}�0?�cW?�>!��k�T�4:>7����j�5`>�+ �~l���)��%Q>wl?EFf>hu>�C3��<8�8�P��O��{�{>�*6?᝶�HC9��Du���H���ܾ{TM><,�>pr>�a�^����
�1i��|=��:?q�?���_1���lu��蝾a�R>�\>o�=\Y�=�\M>Df���ƽ�ZH�,E,=��=�^>s�?j�>'�S=��>+Ή���C�+�>�V?>v>~8??�??Z�Ƽ����_�����2��*�>Z�>e��>3G�=�$D�*P�=_�>�b>��e�J83�����X�&�S>^�b�{}U�]%p���&=?�ֽp�>�v�=��fxD����<�~?���'䈿��e���lD?O+?} �=L�F<��"�A ���H��F�?q�@m�?��	��V�?�?�@�? ��F��=}�>׫>�ξ"�L��?'�Ž4Ǣ�ǔ	�>)#�gS�?��?��/�Xʋ�;l�n6>�^%?��Ӿp@�>���ʙ��4���b�Ei�=(�?�c ?G�2�dτ>پ4?�z$?*����ޢ�����k����>�W�?��?[h�9 ���)����>]>�?ܫ\?t�>\�
�Aॾ�	�>�Z?)�?x�>PYE�z�|�+z�>Su�?��~?;�t=�\�?�a�?>�L>�7Z��]}��ؿҎ��(�?���<��>�������f�G�T�ۛ�������us�+m�>��=�kH>���+_澔=x���=�-��Y-��2�>1��>���>�=0?_l?�1�>���>Cx�3�{�����5�L�K?��?����n����<R6�=�^��6?+U4?7/`���Ͼuۨ>�\?���?[?	b�>���mD�����{��MK�<�K>5*�>�P�>��� gK>��ԾW"D��u�>t��>Wԥ�h<ھ<5��}椻�;�>bl!?	��>��=�� ?$�#?ژj>�'�><aE��9���E�ı�>U��>�H?�~?��?WԹ��Z3�����桿�[�s7N>��x?�U?�ɕ>���������E��>I�����[��?tg?�Q彁?�2�?(�??D�A?^*f>��ؾ֫����>�!?69��A���%��`��?nL?`��>)ƚ�:ӽ��F��J��q��?�Y?��"?]����]�ૼ�Ng�<�������Ӓ<�\s���>J�>������=�>Nb�=o�98���)U�=!�>��=?R9�:��&a?�D>n2���1ݽ�ł�N�#��b>
 ��wý�<X?)D���e���ҿ����7(>�`�?�w�?��f?��v�� |�-i?-�?/%�>�G�>�F��Ӿ0�Ⱦ�~8=C����p*��+�>j(f>���=������Ρ��%��?m\���U��?}�>^�
?&l�>&=G�>F�������
��Ut��(�VE8�K{!�1|�ѭ���q��J>�'�Ⱦ:뭾�N>ٺ�_�>d�#?%(�=�f>�}\>���+�>��=	أ>D��>�A�>�Z>�0>���=+Ȼ�'R?p俾�'�x?���`B?Ιc?�^�>Z@i�$��t��R�?bv�?�e�?�Tu>��h�K_+��b?���>�X���	?�4=,���ʀ�<1�#��v�����ڲ�>��ڽ�9��QL��i���	?�?�S��Vd̾/f׽�L���&>�|�?��0?V2(��3c��X~���N�>r7�n�z�>P�z�ƾ>v2��u�������{��x��/�.��=!"?U�?������(�~�Jg�u8X��O>L�?4�>sՍ>��I>w�/��k���2�����7s�>h�?>��>K�I?�<?�vP?8jL?潎>�a�>�0��Sk�>�
�;c�>� �>�9?��-?-80?z?�s+?b1c>y���:��̆ؾ�?�?J?4?|�?Vۅ��ný�Q���-g���y�rx����=�4�<��׽\>u���T=NT>
�"?�9�:i8����?QML?��>�U7?�0����=8��>�Aq=�:?�W?�;K��ꖿ��K��K?;�?i�U��>��>��������sw�=��=t<A���=����ֆ�<$�Ľ*�E=
��<� C��!=��a;�������<�x�>n�?��>N�>�5��>� �,��M�=YY>�'S>��>}:پ3|��Z$����g��ly>�x�?4z�?��f=9�=��=�{���S��k��L����<a�?[F#?dRT?N��?\�=?j#?l�>�&��K���]����$�?+!,?��>��H�ʾ�񨿢�3�z�?n[?3<a����;)�g�¾��Խ�><[/�/~����ED��
������|��E��?���?A���6��x辫����[��r�C?a!�>�X�>)�>��)�`�g�s%��0;>���>:R?���>W P?�{?_^[?EQ>ܰ8�A(���e������!>�@?��?Վ?%�x?F��>�>@�+�р�0���,�	�������PY=�MY>8�>�t�>��>���=Mgǽ�󯽐 >�*#�=�,c>W��>h��>�5�>�y>�=�<��G?"��>�r���I��������s�0�
�t?ˏ?�~+?�	=)��$"E��1��p*�>M�?J�?>=*?�IU�M�=	�ռ����n��Z�>{��>1=�>��=�E=�o> ��>a��>�z��z�X|7��51��L?<�E?A�=ǭƿ~~q��Ij�۳�����;!��	vb�~z�_~V�hl=і��+��⥾��D���7��:Ѳ�<����Zw���? �=嶼=�G�=�<zΦ�u�o=x�f=�F��/ۙ=�`��C=�Ŗ��U��C��cۻ(�=?z�=�v�I�˾��}?N�I?ʗ+?6C?�y>7q>��.��0�>�g��9?�V>�AP��8����9�w��qO��G,پCyؾ�;c�ٟ���>��K��Z>ȋ3>Sj�=A}�<ZS�=�Bv=:�=\%D��=�!�=�^�=���=g��=C�>��>Eq?��a�-���l�)����*�B?UT�>6����ľ+�>?�wZ>Q�{��"����/�<�y?�V @�$�?���>�쌾�Ua>����>�=����뺾�S�>�9�ӭ����>�F5>�Ծ����l���Y�?�w@$G?'Ń���ѿ^�o>�J8>��>��R��K1�S�[�	�a���Y��!?*;;�>�˾�V�>}��=ض޾�Uƾ��,=�Z6>��c=���l\�n��="�|�OA;=xn=���>6nC>:J�=���(��=�H=|��=yZO>o薻�8<��"+��)7=��=�Lb>(%>��>:�?B0?dXd? U�>~n�?�ξ\.��?�>��=
�>;م=�aB>��>�7?��D?��K?e��>���=��>��>i,�Îm�3�徼q��oS�<Xf�?XĆ?�Ҹ>p�S<�jA�~���>��@Ľ�?mQ1?b??ش�>c�Dſo�оĤ4��0���>��l�󗴺�<��*�yI�4~��l>�=]�?E�?Èq>���=4�3>C�>���>��=�aG:Qʉ=oi=��;��=�٫=E1��}8*>��2=�F�<�(�;�t��iI�k5�=R��=���<&�h=ɼ?Jbm>�R�>c�Z<�6���>#��o��*����Ⱦ\C6�����9���`��U���4>�n�=
@j�o����A�>y�o=o�>��?��Q?�w�=�!�g�%�@[����H�K�˾��>/U%>0R;>�4�f�Y���Q��Ͼ6��>�ߎ>��>v�l>,�3#?�s�w=r�+b5���>||��~��)�}9q��?�������i��}ҺP�D?gF��h��=�!~?�I?:�?O��>'��ІؾB80>�H����=k�n)q�bl��{�?u'?��>쾷�D��H̾����޷>�@I��O���6�0�v��6ͷ���>������оL$3��g������؍B��Lr�>��>	�O?��?�9b��W��NUO�����'���q?�|g?��>K?�@?�$���y�r��3v�=��n?���?C=�?�>��->��&�S�>5!?��?PІ?�wj?�P��s�>�3y=P�=*�x=`�1=%d>����> �?�?1= ?����E���������X��o��=���=�8�>%I%>�9r>=�=�3f���E<�1K>�>�V>Y��=q��>x��>8���7Z��)`+?#��=���=�?c�c=������ͽ��-���I>R����I�fV�HO�=��>�8���%ý*�,�7��>˿B-�?}m#>D@-�7�&?_��V�>��>�>IZ>�>��>	��>�?�Da>¼μ�kT>$�o>_��R��=����6B��w3���/��/H���L>r�Ҿ�7=�
��丽T�!/��|����V���e�	)+�ћ�=��?~ܐ9�A���fE�
7ܽ�?�~?�T?��񾯋H>o�B���?��>�N�@����܌��1���Ɖ?�~�?Hc>�+�>�W?��?I�0���3�7&Z�h�u�SA���d�n�`��Ѝ�����v�
�)ȿ�u�_?H�x?�JA?.v�<Z�y>��?��%�Rҏ�P�>X�.�Z-;��o6={	�>g���_��Ӿ��þUc��;G>��o?��?{?��U��+m��	'>��:?��1?=Ht?��1?M�;?}����$?c�3>u@?|w?�G5?O�.?|�
?m2>�B�=w+����'=U;��0ኾ�ѽ�ʽ��,�3=%M{=rD����<��=��<�Z��ټDC;I꡼��<�:=Nޢ=_�=���>�3]?���>1�>�7?�H�.B8�����.?s]<=F!���������@~��>�k?�	�?VoZ?� c>��A���B�9>gL�>�^&>he\>��>���/E�l��=q>�<>�_�=��K�������	�����+�<6>pt�>�">cC��ɫ'>������}�=�b>Q.T��I����S��G��1�(�y��q�>��K?ӿ?!�=���	ם��'f�8c)?�.<?�eN?��?�g�=}۾�9���J�LV��p�>��<Y���j��Հ���;�V���3o>���-���DJj>����Ҿ��n���J�ړ�ld=8L	���<�|��ݾ5`��!��=��>y���� ��ԗ��:��rfH?'�E=ҥ�
�=�^!���	>k{�>Q��>�u �7���qA�K������=�v�>�:5>O�����$CD�� ��2�>��D?
	`?�8�?Kp����r�cqB��i���_��il���@?J��>}R?(2@>$�=J����;��e���F�خ�>��>�N��8G��1�����&e%�)g�>�?t!>�?hQ?)Z
?�_?@�)? �?�;�>�h��|귾hA&?��?U�=��Խ��T���8� F� �>�)?M�B����>ۍ?ؽ?�&?ʃQ?��?��>!� �@@��>ZV�>E�W��`����_>[�J?[��>�:Y?�у?��=>8~5��㢾�	��6F�=�>��2?�9#?V�?Z��>Z��>l]���=�g�>�Lc?��?{mm?Ȧ>��>K�>[�>p�=aS�>�
�>R�?�)I?�ar?�&J?I��>�<{	������^��L4�	 �<�W<0�=-|�pcW��.��\��<T�<]���m�:z�"�we�D�R#�<-�>5��>����Œ*>r���!o���Y>M8;���{����2����=Qe�>�� ?�M�>_�-�]�=���>���>Xt��� ?yy?$�?"+;O�^�"���KY=��`�>՘6?���=��[�b񕿐*p��Xc=�.m?�d?)��Y�6�b?��]?�b� =�5�þ�lb��V��O?6�
?��G���>��~?��q?���>-�e��;n����*b��vj��=��><?���d��2�>~7?U��>u c>{O�=ew۾ӏw������?-�?M��?��?��*>D�n�/7�f���K����]?`y�>����"?�c�%�Ͼ^T���+���
⾨1�����C��􁦾V�$��ȃ���ֽ(�='�?,s?�Rq?*�_?�� ��d�Q#^�����hV��%��'���E��&E��C���n��K�� �����{F=Г�E�%���?�#?N���>	��mƾxYӾ�e>"�'���e�?Ά�>߻��T�>)>�@�/u��鑽��_?��>���>\B0?m]�V�I���A�,��*���"P>Z��>/�#>:��>��;��Չ[���.е�7+���_�=�.x?�m?�km?�ɔ���C��v�A����>�%۾��h>�j�=.eF>v�e��}!=T}�x�B�o���)�$�7��� ��j@��#Q?Ï>�}>%��?>	?f!��h�� ���l�Q�������>]Z?�}�>���>Ŝ�<��6�ǲ�>��l?���>,�>;����\!���{���ʽ 2�>�߭>!��>K�o>װ,��#\�fi������|9��4�=�h?ـ��s�`� �>�R?̸�:@KH<�z�>��v�=�!�����'��>#�?{��=��;>�|ž&#�Q�{��4��7�(?��?&���
*�`�w>"?j�>�=�>�-�?�̖>w��A�7<?�6^?��H?�>?�R�>��.=����Ľy*�ظ'=��>�4T>[z=rF�=u��f^_�X�%���a=���=��#���ý�s�;�����<:&�<�s)>l�׿T�D������m%��]��ᾋ���}�'쿾\�Ѽ��򝠾F��d���w=0���.��G��T�F�j	�?��?�9�����n���Z�|������>�����>���1��Z�F��K��}Ҿb��� X��to�F{2�U?�]���)��k寿�Ҿ�
??�W?	G?�x�I�|��
g�B��>8iG>��=���ϫ��$eſ�?���o?�?�(�
���`@?f+�>2G�>��=p�u��T�GD���?��?��?�����Ŀh���v�a<K�?_@�{F?�[2�K$
����>�)8?o��>�sh>�׽���8�X4�
ύ>�N�?��:?�#Խ����7_<>��?�s>"5�h<Ĳ>Dm�=����ͪ齬�p>Y��>�伖�:�n��o
J>���>-��O�_���`:K�����=�I��{�>�Ԅ?Ty\��f�)�/��T�� V>!�T?�%�>'9�=s�,?�7H�^}Ͽ�\�A&a?�0�?���?��(?�ؿ�>Ԛ>u�ܾ��M?�F6?���>?g&�^�t����=����W�㾼&V�|��=i��>��>�x,�
���O��]��x��=��$Ŀ�-�����З�!��"����I*������	�i��ͽ'�=ns>��U>$��>0�@>�C>��Y?��g?m#�>��>c����S��7��=������tW��}E1�*봾�|����޾v������dc�-d���#=��=C R������ ��pb�M�E�ʕ.?�A">�
ɾ��M� �'<:1ʾb�������Fa���̾4�1���m�$�?�B?3h����W�x����t��"W?5l�c���)��{�=�ӟ���=�g�>�=���F3��S��'?��$?ʚ��jBp�0=��=ĭ�>��)?\|�>g���T?K{@?S���^Oκ�0'>��=\"�>[y�>�+�=|�f���0�eZ�>��??"�3�#����t>��?����Ӳ�=3yB>S�'�w����=1h����W�>X�b�0�W�/W?��>i*��7��p��̿��E=v/x?o�?Ę�>huj?ۡB?UL�<4���S�
���=��W?�>h?j}>Y�t�dqξ�E����2?�,f?��N>��a���/-��)��N?�Sn?��?�hT�\U}����N;�hX7?B�l?Z[�L���H*���%�=*��>��>eM�>^�7��3 >�>$J����p�݂����_�<آ?�>�?���?XEj��<���F=�%�>���>�c��'���E����"�@O�}�>�����B�KM��g۾h8�>ZS�?v�?r+#��_�&c�<Ov����?)��?.�Ⱦ�&�N
*�~�R�.Lо���=��v>a/H�ݿG���ݾ��־������:�ғ���>��@p�p�|��>��e��&�<�ǿt�z����w�E�S?eFQ>�$���5��B����9��tY���?�w,-�S�>z�>���_��!�w�Q�5���<��>D���5�>ryo�}L���֛���:,��>��>ӧ}>�׽������?n��Կy����iU?�?�R~?U�?�@�=^����nT�� =�%A?K�g?6�H?迼��,v�j��g�j?�r��8V`�̇4� E�m@U>�3?�@�>��-��+|=�>\R�>��>�/���Ŀ~Ͷ��������?�~�?�\���>�y�?{+?�_��6���>���*�z�Q�D,A?��1>�k���!��3=�s�����
?��0?u^��C�]�_?+�a�N�p���-���ƽ�ۡ>��0��e\�"N�����Xe����@y����?N^�?i�?ֵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�
i	>���?�~�?Qj?���� ����U>
�}?1��>���?�n�=���>���=5R��в���X%>���=�W?��@?OGN?o�>�6�=�)6�!�/�4<F�<�O�����:B�8�>1a?�J?��_>�ɻ�k�%���۽k?5�����Y�4��_�Uݽ�`6>��B>?�>�-8�g�ؾ#�&?�0�)ʿ����=�H?3|>��>Ά��r~�Np�� ?g`�>1����b������ �e� �?���?Z��>[p������@>-� ?��>�Y�ʭ�=�'�WR�~ `?�6Ӿe���Fk�	�>px�?�2�?�{�?X���q	?���H���}���P~3�+^�=�l7?|4��Cw>C��>A̞=��t��D����s��ȶ>���?O�?���>x�k?��n�6�A��OE=|�>�si?HE?�!��f2�?8@>>.?����掿����c?%�
@�L@C�]?�8���ҿ䊓�>gJ��t���:��D��y�=����>��=�d����q�a��>�f�>/Q�>���>�0�=	>�K�=��}��f)�����,��ZED����g���R��^`G�� &��#2���澓���C(���6���=���������O=_��<�X?�a?�9�?�8�>�1[�*>o?�R%>e����n��E9>�%?��2?}4?���=����|5m�	��L0��������>h�e>���>�>u��>Y�=�SB>, 7>�a>n�F>QW=�B=�e�=c��>�|�>Q��>*��>lC<>Y�>=ϴ�/2��J�h�?
w��̽� �?����/�J�2��9��H����h�=b.?�z>����>п'���
3H?����)���+���>��0?�cW?��>n��3�T��8>�����j��a>�, �j�l�ˎ)�/&Q>�l?`�f>�&u>�3��Y8���P����� b|>�26?`۶��_9���u���H�`fݾ�EM>�Ҿ>�C��j�h������mi�Wj{=�s:?R�?S9���谾>�u�!9��aWR>�/\>�=M�=�OM>�_c�Q�ƽ�H�{.=]��=̢^>t�
?�mU>�>
=�k�>+V��-(��{�>�֫>�ܵ=>\)?�3?O��=�9̽�0_���/�Ȭ�>�r?#g>.��;�7�,��;��>��>���=�eN���Cz�o�!>E\=�樾�\���<-2B��И=e��>B!C=B`۽v����~?�|���∿�:U��eoD?�$?� �=>�G<�"�����E���?{�@�k�?�	�C�V���?aA�?-
�����=�x�>�֫>�!ξ��L�}�?�+ƽ<���{�	�*5#��P�?�
�?�H0��ȋ�l�->�U%?��Ӿ��>Z����S��:o��Fz=��>�=?s��K�8�Y8u���?n�?��پ�<��K2ɿ�ew���>���?Y;�?Ĺl�?H����.����>)2�?�F?��]>~�Ҿ�K�����>U�3?cYO?�>=���p*���?���?��?�2�;���?F��?兼>�r;It�<�˿}�W��?�>��?ה�>Y����N�M�j��v�\!w�1M~�v3B>-{�=+?�>�,���9��5�c��=Pt��Sx�ִ�>�A�=���=,?H�=?��>�[>ݿ6�������!���K?Q��?.���n�j�<��=9^�6$?�D4?��[���Ͼ��>��\?R��?U�Z?"�>.��%(��7ʿ�Gj����<F�K>'��>5(�>A����K>�Ծw�D��;�>��>�j���ھ ��ۢ���^�>T{!?��>r�=f� ?4�#?��j>'�>)`E��7����E�ñ�>9��>�G?��~?y�?�͹�QW3�r���桿ߒ[��8N>7�x?�T?e͕>���������GE�=iI�֒�훂?pg?uU彏?�2�?�??W�A?�+f>ɂ� ؾt�����>�T!?;� �/�?�Q%��&�0�	?3w?f�><�����j���ǟ�����XH?K�X?�3"?�B��[�"濾{�<�;�����|�3<�ކ�˂>�>�ц���=
>WP�=�&r���L���:D]�=�z�>��>��<�>���O?k8J>U:@�`fk>��>�7���>��R���C�e?n��{n�Zt��vZÿ>��?��?�r?�}뾻{i�5g?��?��	?Ơg=�U/��+о�c/��a>(g��-J�c��>�=��=�_���䥿���݂������MN�W�	?4�>m?Z��>y��=���>侬� �oK��M�GqG���,��^5�� �^������ b�C*���ľ릾��>iB#�69�>'�?�\{>�Ґ>�ݐ>1���v�>�}�>r��>I&�>�֜>1Cy>�O>���=c��<LK?(ב�@~"��۾�Y��3XB?r�V?�f�>�}�<H+t�����?��?m՗?w�f>%�l���0����>I�?��l��?c��=z���ʈ<��ɾU8k�����ӽ�o>����2��#T�N�P���?x[?<ŉ=5��m3h�g��̀�=�ʇ?��-?��+��@Z���t���Q��aF�*�V���4����(s*�.`k��8��Q܁�:���.�c\=��'?�!�?�r�����㹫�Wyh�Z3>�me>���>�y�>���>pUW>����o/���f��,�L/��E��>�z?��>�pI?3q;?IP?3�K?�ǎ>�0�>���H��>b��;�>t��>�$9?S�-?/�/?s1?=�+?�c>�.�����ؾ�?��?iD?ek?br?o��@MĽ4���Yq�,Hx�p�����}=	�<��н�g��KV=�xQ>�(?�3d��U1���4�?r?u���ͳ7?e�<��Ѿ�Q�>��L��!?^h#?3q��jb�1E��#?vK|?��A���Q>�)>�)2��(�m"
>��D<�_���d>�O�<�n���;�sE>�$>�dv=i�~��`�b���Z�=_��>��?���>���>rK��ڋ ����2�=Z�W>!�Q>S�>�ؾ�e������"h���y>�}�?�l�?'e=��=`[�=�f���R��X���y��=�<Z�?�#?�5T?>��?k�=?X#?�>}���G���S��f"��`�?t!,?��>�����ʾ�񨿸�3�ʝ?i[?s<a�����;)�ϐ¾G�Խ�>�[/�n/~����3D��ᅻ����~��)��?忝?$A�N�6��x�ڿ���[��l�C?�!�>Y�>��>Y�)�v�g�g%��1;>݊�>eR?�3�>��P?`�{?�[?8P>��8��P������r��J�">��@?i5�?���?e�w?O��>g�>xZ,�q⾾���� ����� ��&[Y=��Y>v��>�x�>�b�>q��=Rͽ7����TA���=�
f>�$�>��>���>|y>-��<��G?z^�>�����g�К���ۅ����N�t?7�?��*?��=(���'D��*��ce�>�ɨ?Uܭ?�A(??fk�A��=��V����t�k��>�>7v�>��<Z92=7\>	T�>��>Z�.�47�85�U]�N�?�.F?��=�1ο+~��*h���q����Jޮ��pP�w������>w��m/u��u���#�钜��er�/F�����o�y� ��>�}�=���=k��=���=�&<^>�d�<6�I=V�<�
�����l�Ͻ��< 	5;qH���<�h�;�Ĵ���˾��}?�RI?��+?}C?��x>j!>�n2��>|���j?lUU>BQ��h���:�����u+���پz�׾I�c�ٟ�:>+8F�V�>��2>� �=G6�<�a�=�s=T�=^T?�=��=c��=AW�=�N�=B>2>�2w?=����:&Q���2�:?�8�>M�=��ƾ�@?�>>K3��7���w��(?���?�W�?g�?,�i�R�>6⢾�[���,�=Ӄ���U2>���=�*3�@��>��J>3���M���峽#%�?�@��??ދ�L�Ͽ�R/>��K>���=�jO��)���P��D��5�\g?X8��dھ���>���=Ueܾl¾�� <7>\�=~I�� X�ˏ�=`,���D=��=vA�>��'>���=�U��*�=R�=���=��H>�I
��C��9�5DX=]�>NzA>c�>���>F�?AR0?v_d?䨹>�n�Y;�뾾�Q�>]��=�ޱ>Tё= �<>x��>��7?&JE?�eL?6�>OZ=7x�>���>��*�U�l��徼�����<a�?�?��>��G<�lB�Y����>�������?t�0?�?*��>b�����t���1޾Mtf�uq�9��=Q�b��D���>8G����˾D��>�۶>�$�>��>ϋ:>�w=��>�ª>�g,>����s�1>�x�=$j=�7���ڊ=$l��P��;.��=am�_�Ƚ~�<�ن��g��=Q���ּd�=w?X�>�?�b��.#��>a����C>�����X������"����ΎK>�tc=𘚾�󎿩�>˘�<R�(>���?e�z?��b>p��03�E5���,��?WU�3�^>Es�>Ѷ���O��Pv�6S��僾��>�>���>Q�l>%	,�h?�~x=�⾝S5��	�>z���|�����*q�m:��g����i�GҺ"�D?�A��+��=;~?��I?tޏ?q�><���urؾd0>H��g�=&��aWq��E��b�?G'?���>��뾜�D��H̾>���޷>�@I�/�O���R�0�Y��,ͷ�2��>������оj$3��g�������B��Lr�Y��>%�O?��?Z:b��W��IUO����i(���q?�|g?'�>�J?�@?�%��z�r���v�=�n?˳�?S=�?j>O��=�ֽ���>�+	?��?�?��p?H�,�h��>گ}�GX$>�o��4�=�)>CqT=��=(�?�V?I�?�4��%f����^�����n�Ff=Q��=n��>F�>�mt>VG>Gl=�x�=��_>��>�Y�>��K>ğ>��>�Ižf�̾��<?5]J>@t>c�?��w>o��̛�^�<Il�d1�I����&ǽ���=z�C>�\L=�g��
�φ�>#:��o�?�*�=J-�a?���U�>_�	>vС>�h>|,�>��>�Y>t��>u��>y�>TB>��8>������=K���Z��:���4�V-�q�2>ǵ̾p�+>1M/���X���Y���@�꾄Oa�w4���PD�;=M�?�Uͽh%��0�/�UŽM?X�>�5?D1�(�<]���R�?v��>�9��yW���
��H�
���?���?�i>Cȝ>��T?G]?.�0�4�2�q!V���t�SI@�`a`��aa�n�������N�{�Ľ'�e?N,}?_�@?F$O���q>� �?�Y!�Y���lv>/'��:�x-<�\�>����T�l����c�ʾ�o1���[>Zp?��?v�?��T��nm�k.'>ӫ:?,�1?�Gt?��1?��;?���M�$?sU3>�J?Vu?�K5?�.?��
?��1>��=i��K�'=�/��#�ӣѽm�ʽcL�W4=�_{=�O¸�^
<7=㔦<<��{�ڼ"�;�@��X��<i�:=�ݢ=!��=���>�\]?�%�>L׆>K�7?v��J8�����U�.?b[8=x������> ���"��>�k?,��?�@Z?o]c>٘A���B��r>�T�>�)&>��[>u�>�1�V�E�*S�=<�>�>z�=$M������	��f��><�<<>���>S1|>���ȹ'>�{��l/z���d>�Q��ʺ���S�f�G�}�1�=�v�~X�>F�K?,�?R��=&^�x.��AHf��/)?']<?NM?@�?��=��۾:�9�`�J�H>�X�>�[�<n������#����:��9�:�s>M4���)���c>��
�m_ܾ��n�v�J�&�f�C=y���R=6��P�վ �}��e�=��>�����,!��2��QЪ�&�I?�g=:8��ԨR������x>9K�>p��>h�<��ir��\@�`��꫙=}8�>_�:>�W���N�߅G��(����=�1a?�_?e��?�:ۓ�f?��/	��a���G�au*?��>{b.?���>6�h>'���m$��S���k����>�C�>%<6�\�p������|;��?�g�>Q3��*?�}�>�[�>ί|?N(?�c�>fh�>9XM=����"v?&�?
<>9�������I��mH��??�N8?N�ž���>�Q�>��'?�B?
g?lp ?�4l��?���[�lڣ>~l�>��q��*ſƒ�>�oe?`�K>Cv�?���?T�=#I�UA˾�'���<弔>@0)?�	?�+"?��> �? �p�d��	�>1�?�HH?L�7?�b>��<>��g>�����>�K�>k��='g>�vS?uӃ?�X,?j��=��Q<�H�Nu�<:UY���˼��{�o	ѽ�4�k���k�;>tܽZ�(�S�7�y���;>�;I>F*L�J;��|�U��>�,�>����)}z�حžU��蔟>/�z>�]���Ԧ�TI�=�c[>��}>08?�[>f�y�jn�=Mb�>rV�>���&+5?���>�]�>[�$=�+��������l��=H�M? ׋<Z��J��KK������p?'?�P��w��K�b?��]?5h��=�	�þ|�b����g�O?@�
?<�G���>��~?e�q?W��>��e�*:n�*��Db���j�!Ѷ=^r�>KX�Q�d��?�>m�7?�N�>8�b>,%�=ku۾�w��q��f?��?�?���?+*>}�n�Y4����v둿�^?�l�>b���^"?`}?�&�ξ�k��q捾n��|֪���
���^��xO%��.����ٽ).�=��?�s?Iq?E�_?I� ��wd���]�����sV��~�Ƒ�$=E�0E��CC� o�/�?���d՘�@.T=xK���Q"�%(�?Bc?��V�>���������V���k>Ѩ���~?�<��[�c>��=@�n������־�?�P�>��?�:;?Z�Y�O��6�'A.�p7�����>_}�>tR�>�o�>��1��x��.茶�R��V�� =��x<}��?̲v?Err?�9ξ��d���t���
��>�*ܾD��>���>Õ>آ��g�=`�&�T�f���r�����-����=��q?7�e=�<�`�?<�,>�!*��ỾP���Q�G�G��=t<�>�K\?�q?��>C)��^F�̗�>��l?���>x�>����g!�J|�u�ʽ�B�>SЭ>L��>�!p>H -�1$\��_������+9�(��=�h?�q���`�	��>��Q?�8�:��G<Gn�>�w���!�����'�4X>6y?z�==a;>��ž�/��{�j��)?��?ϔ��;�)�.4�>��!?��>���>�f�?�W�>"�ľ/g9��?�]?�I?��A?&x�>�2"=�\���ZȽ��%�cC+=QT�>�FW> ^r=���=�5��]�	��QWF=ތ�=,輴f���72<�Q��� B<d�<v�3>Q�޿��M�@Ӿ�9���ھx���)��+���p���#	��ų�F����v�������<��D�l?O���HN�#)�?�:�?llپpC���^���^��|��v��>��~��=6�Ӿ��W�������xpȾ���s?�@|R��G�l�&?%钾ٸǿ�桿+I۾�  ?�� ?�Iw?IZ� ���-:��� >}=�c�����з����ο����`?��>xﾬH�����>#Ɓ>r�[>�Au>/����!���;�<#?�^.?h�>�.q�c#ɿ�H���ք<��?�@�-D?�n>��d�j��=6�?�?܁>��L���#��$0�Ъ�=$\�?*]V?д��)H�"�!>�r?ȕm>CG%��ۻ|��=څ >�>+��!Q>s�">���l��}u1����>�p>G��2as������F>��>�� ��<!�1u?�,���8��p%�2����n>��-?*oB>�֜=Y�L?D++�mTؿ*Ձ�E{?o9�?)b�?4�0?�Ӿ7#�>ba���.s?�=2?k�>��G��`���z==z]���>���P�k�>[Z���}���1=��U=�r�aI��6�T��=0��ƿt�$��Q��=/?�IB`�}���<X����?�r���m�q=^��=�Q>��>�lU>	+Z>�NX?+�k?�F�>��>v���m���˾�?K�����%��p��9��鋣��|�R��Z-	�Z2�h2��ȾO!=���=�6R�H���� �K�b�3�F�[�.?}v$>��ʾn�M���-<�pʾ࿪��Ԅ�Xॽ�-̾�1��!n�o͟?w�A? �����V���R�\����W?�R�@��$묾���=���1�=�$�>���=<��` 3�~S��/?tb?�l���Ð�W\,>>��t�V=��.?�9�>T�<�֯>��$?J+�w�dHM>H�6>�}�>�>/ >�먾(�ｴ?K�T?��н�C��EԊ>����Up�z�= I�=�7�'5��D>��<Ϭ{��(�;Y��f�O<R�M?,�->�%�����'���=`lr>�q?��>���=h��?@�"?�;<�兊�/�l��޾�Z>+X?�/?��>�=2�z�ƾ̜����g?/�-?0��<��G��@������z���=�>�^i?��o?��>l长ޝ�� ���V?��o?`[�M웿�sྜ!&�Q��>�>5��>�s=�록>�#?�����ۑ��"���x:�7Z�?�$@���?�M��P���(�=��>3y�>�y�����,��%d���Y=�e�>�\U��de���6�`�(�@
?�>l?���>@�,���3��=dw���J�?Ux�?d'���F��/��>nc�����D6=��=����H��2�@�/��ɾ7�d����;9�>�@��ӽT��>�&6��8⿙�ʿ����=Ӿ��b��?��>o����g����n�<�{��H���E�m�i�	�>�o>�5�����~|��<����kV�>e��.��>�=L��Z��EƜ����<8*�>hO�>� �>y���o����?
	����οѶ�����=�Y?U�?�Y�?�?��;VHx�����S.B�i�F?��s?uY?]�*�c�W���7���j?�Q���M`�א4�nAE��JU>%3?�Y�>�-�[�{=HY>B��>�v>�/���Ŀ�ն��������?���?jj�t��>�x�?6j+?8g��9��M���*���G��6A?2>�����!��:=�MԒ�׾
?n�0?���1�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>hH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?��>�#�?���=��>`��=S���+�.�>c��=�A��]?W_M?��>V��=��5�O�.�~�F���R�o��MC�A>�>ha?hM?:`>����(�-�!��ν/�P��1�?�g�"�����4>�U?>��>}�F�#Ӿ��?�3���Ϳ"|���5����M?@?b'>>�6�G!�>����xE?���>�2�����v���5S�9u�?g�?4�?2A�J��<�9�>�@�>~@�>i��9o�<����Y)L?R��=G�����S�DV�>9��?M5�?۴�?A}��	?M�iH���Y~��p��6��Q�=�7?M��z>���>�0�=�_v�Y�����s�׫�>6=�?cm�?���>�l?B�o�x�B�
�3=[v�>��k?�Y?��y����H�B>n�?��E󎿇P�jf?&�
@�o@ɕ^?�袿4��ȃ���Ѣ��+��!��<�	X� %>(
��8ڻ���i�a�&�Ľ~�3>�m�>��{>;��>q�8>oP#>��I>4����%�ޥ�T���*�7��<�����:����A�g���"��X�o}��ö��^��o�<e��f�	�L ��`�<��_?�f?�c�?�5s>�|����H>�%�>�>M�%��?k=��>��@?Z�@?_7?��5=(^Ҿ��ڌ��׵��qnz����>�B�>��>wm�>��>z���n>RE*>H!�>��>�>�x==᫒��w>#i�>���>���>�C<>��>Eϴ��1��k�h��
w�w̽1�?}���T�J��1���9��Ҧ���h�=Ib.?|>���?пf����2H?%���z)���+���>~�0?�cW?$�>��|�T�/:>:����j�2`>�+ �|l���)��%Q>vl?}�f>�u>�3��`8���P�@w��'|>�86?!Ҷ��D9��u���H�mfݾ!+M>پ>N~C��f�3�����bi��>{=E�:?��?vu���䰾�u��5���LR>��\>Qg=���=�sM>ǚc�;�ƽ�.H�?.=���=��^>N�?�=۞j=�^�>$}�᩵�@%�>F�[>U,>Tq+?��?�9=B����C���������>+?:�{>Zn$<���%��r�>
S>�����<��@�cc��Ys|>�R&=��~�>GA��2*��M@�R �>��>���;ʌ���Q=�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>�g�/���j���ZV�b��=n��>��?X�#���>vھ�)�>�t?�����1���Ŀ�Bw�{$�>�7�?���?�V�ߘ��yO/���>���?�d?ܤw>�裾S(�(�6>ފ\?�7a?�>)+�䎘�M��>��?�@�?�!A=�u�?3��?��>�C���"K��V̿�.Z��H�>����j�m>�;�>�Ѿ�UE���j������
���P��1�>�`&=9o�>�|H�E"̾���<F.K=S^��⢽�r�>��(>o�>_��>�T2?&�>yA�>I�=�sj��>������w�K?���?$���2n�dN�<^��=��^��&?`I4?|j[�/�Ͼ�ը>ͺ\?_?�[?�c�>"��=>��3迿!~��K��<[�K>14�>�H�>x%��FK>��Ծ 5D��p�>�ϗ>�����?ھ%-���W��|B�>�e!?���>Ү= � ?b�#?�k>�7�>gbE�$<���F����>n��>�<?��~?�?����'^3�����l顿F�[�/�M>��x?zP?_͕>�����~���>D�d6I������?*�g?�'�(�?�8�?�??��A?�e>��
%ؾ�Ȯ�:*�>��"?����<�Hi!���	�:U?%?���>�>�������Ӽ���pC��k(?p'^?�0-?�����\��j¾܂�<�
��M����f�R�7�$>�}>����y��=S�)>�F�=�$��,�U����;�)�=�>���=�C�J�T��?��>:���e�z��!@���=XZ	=G\���b?/���5��|@Ŀ�S��u��=���?�"�?6n?��@��Bv�F�Z?[�?K?ZI?����������{�ɿ���c ���v>z��>'ަ�4.+�\4���!���n}�#���Vzg���?���>�<?���>���=�܌>Ӿ
Q
�)-��徟�f��i5�bP;�F��UB���������P��*�̾�᩾�O�>��`�X^�>��?���>7��>~)�>��܌>c�!>��X>Om�>,3z>�NA>Ш�=B��=�9Q�dsP?�̷���#��Y���F?�c?���>��g������"?�^�?Wӛ?%�n>	�h��'���? `?�����?��3=�In�]�M�g�ľ����*��<6�r�>�D��2r2�b�M�=���4?�?���<P�׾+B �������1>"{�?�	.?T�3�A�_�����}�3���$�d�==ZU���q�S61���k�"4r�M͆���~�2!1�_E=N"?��?B�9Ǽ��8��eml���'�kM�=��>"y >{5�>z4�>Co�s$�r	g�^E�����v{>Ɏ?��>J7I?K�;?ԅP?�bL?X׎>uR�>v����u�>��;mҠ>���>�\9?ig-?L20?N�?�+?�c>����L���Khؾ�?�K?��?�C?ES?�y��[�½����k��{��À=���<"�ԽJv���N=�MT>i�!?��|�$�"���$���?QtA?`�>n�.?�H+��þF�>ˌH>�k?ǺF?�n�շv�|n&��?��?d�G�@�>Ao>�b:y2�#�=FΚ=��}�Kh�<�g�Î���>ŕ�=�������=���;���sGZ�붤=?e��>d+�=�>����?�w��P��eл��g=x|C=yE>ᮾĎ�ic%��F�>9i�?C�?ߘ�2��=Y�X>խ�8���n�ᾃ����,>M]?��?P�1?�ߡ?�(?�?6��>w}�]X���de���f��_?s!,?	��>�����ʾ��։3�֝?i[?�<a����;)�ݐ¾��Խͱ>�[/�g/~����?D�4���T��6��?�?lA�W�6��x�ڿ���[��~�C?"�>Y�>��>T�)�}�g�s%��1;>���>jR?u�>�P?3m{?y�[?�Q>y�8����љ�	��Ր!>��??3��?��?+�x?���>[�>Wd+���ྷ������f��c���^`[=5zY>6Q�>V�>���>�<�=��Ƚy쮽Ү>��s�=šc>`�>��>��>eUw>�s�<e�G?V�>Z¾tq�	E��2m��e$� �j?��?ߜ)?ù�<A�DC���ƾ>��?��?V�)?;�_���==��� �����s�W��>r��>�|�>�X=�H1=�v>D3�>�v�>�09�QW�� 7�O��?	nD?,T�=�ſ�q�Fq�������h<�����d��ʔ�P.[�c��=5Ҙ�\��婩�}�[�����em���׵�!���&�{���>�n�=���=�=�)�<�ɼ��<�J=���<7�=��o��hl<�]9���л�������p\<�mI=
9��=�˾׷}?�=I?��+?�qC?��x>�>�9��>鿅�+?OeT>8�X�ų��,;�`��90��mEپ²׾.Md�'j���>ruI��m>��3>���=�]�<���=b�m=pR�= Wr��5=�l�=��=kg�=U~�=�>ϊ>nYv?��}�o���8J�~�I�<?��>=W�=����M@?8�<>�����Ƕ����4��?9��?�?��?�k���>�k��ɒ�l=����j�<>�¯=8�<�Sߪ>��Y>���ट�p���=g�?�@h�>?�+��.4Ϳ�L?>�M_>�K�=�jO��Y'�����<���+�?Rh>��귾�i>���=s�ƾ�!Ѿ�'����[>_�>�t���oT�܏=􄄽P�@=�ڹ=��>�b<>��=�xӽb�=2&�=F]�=(,->A�J���k��Z!���=��>�{d>�T	>s�>�X?�Y-?4`?J[�>�GO�tW̾�ľ�y�>a��=E��>��-=�D/>��>��;?�qK?�L?,�>Vo=��>?��>��)�hXo������̞�=<m<���?�N�?�.�>�߄<�hk���#�h;��5��ކ?}�+?�0 ?�ߤ>��6&忲������G�DB�'�K=�B���N�����y^�P����?>�1�>�)�>Ѿ�>l2S>Q�T>[S>��>
�=	���ŭ�=96H=�֐=�E=OL?=5��<�YX=/5=iv��9.��Jݽ��T��*������e<�����7=�?��e>ԛ�>8L:=�,Ӿ�EQ;���u�I�<=X}����L�W�x�t퇿�~�{� ���>>EI=�(A�aR��f(?�^>ҍ>�}�?�c?Y5b>U\0��v
�ȳ���.<�����P>i�n>��n K���q�1�i����^��>`ߎ>�>1�l>�,�7#?�r�w=�[b5�r�>�|����3)��9q�@������Ui��RҺ�D?�F�����=\"~?�I?a�?Í�>B��ؾ;0>�H��<�=b��*q�1i����?-'?&��>�쾨�D��H̾���޷>�@I��O���2�0�լ�^ͷ�*��>������оh$3��g������ӍB��Lr�N��>�O?��?�:b��W��,UO�����'���q?�|g?��>�J?�@?&���y�r��v�=�n?���?I=�?}>6��=�ý>��>{�
?L�?ϝ�?f#l?�C�>��>6��<bw>�T��c9�=:��=�=��!>f�?c�??�������A��g���!}�=�.b=�z>t�w>O�{>p�=�J��w9:=�@Q>?��>'��>��P>�4�>�2�>l���3����?�W�=1�S>� ?u\>�xo>(��{g�X��;L����J���3#���Z<d��=��=�9B�b�=����>-�ٿ���?H��>"��*S?Y�2�?TF>�W�>o��>lt��s�	?g@�>�t^=:��>��>���>��>J�;`��Un�<���%�/��n#��5�6`���=����=�� �_(��3)�Djw�������V�#�f��9%���=�ͫ?}󙽎��Cq9��/	���?Cq?�?�پޑ>3���<?�t�>������攖�#����?���?��c>5��>�W?�}?d1�	�1��BZ�	�u���@�n�d�`�`�,ҍ������
�+S��I`?n�x?KA?2\�<B�y>䌀?��%�aO����>��.���:���:=T��>fҰ��A`��DԾ�Wľ6@�P/F>no?~��?�?�mU�|�l�>�&>{�:?ғ1?f^t?��1?�;?p����$?�v3>�"?np?�T5? �.?��
?�:2>Ȅ�=È���'=,6��B抾�ѽDdʽ���W4=*N{=����	<Nb=�3�<���}�ۼp�;v��iѫ<��9=Ԣ=�=D3�>K�[?��>l@�>�7?d	��J7��W��.?��B=�Ɓ�/)��E��s��z�>l?�ë?�Y?Y`>��A� `A�,�>Dy�>�/>	P`>tN�>�����G�	Ռ=�T>�>.��=�K�ǭ}������V��<d�!>��>o�>?�F�0R>;���Ɋ����B>�l��d��c�-��K�x�;��N����>��U?ߡ"?~�=����ǽ��i���0?��@?�tK?��?,�<�m�;���;�׈>�u��>�pN=Yo�C���֥��B��a����V>J����䟾�,c>^���I�L�r�"QH�.}���s=�`
��VY=��,�о�h{��l�=��>V׾��'��Q���ũ�+6L?�!c=ו���td���y~ >��>���>�&��Y���f?��5���?�=���>�NB>�!�s)���F������>?�E?�e?���?Vp���r��LK�����ݥ����;��?CC�>� ?
�	>�V=��¾\�V9c��N?���>s[�>�����L�]a��e꾫G���>��?b�
>5s?��]?��
?�l?�{(?m?�O\>�澽5þ&�%?G��?�՗=����dO��\:���E���>({*?��F����>e?�?�'?�(R?�K?8P�=�4��A��В>� �>�lX��k��Q�g>��E?�>�/[?rw�?�o3>:�6��{��C8�����='r/>��3?4#?�?�w�>}��>����
��=1��>�	c?�0�?��o?���=;�?�12>1��>1�=$��>��>(?/VO?R�s?N�J?.��>���<�9���5���s��"P�}�;��H<W�y=B��\6t��G���<��;���F�����÷D��֐�[��;`��>A�>ݳ���lw>���ר����8>��=�����B�+^�<�U>� �>郱>ӑD>�����ǉ=���>K�>װ�i�>?�>��?*� >����x9�����,7>�rj?���>�I�S���=���`����*?c�q?F{<�W����T?�Gd?�t��.�v	��;*��;���/n?��?� /�,�>l�?�w?d��>���
�@�������w��V��_�=���>�6+�ve��H��>��?FR?z?2�>���������9?΁�?v�?�+�?#�=>l��ٿ,�����_?S>�>�G��֟#?h����ԾV$���ɇ�afᾌ����㰾�B��cD������M��p�Ž^t�=�n?4�q?�q?"�_?+��Tc���^��B���GU�q��y��	F��E��ID�V�k��7�������n=pts��^=��y�?��-?���~�>C�������\ؾ>�(����!��K"<�ఽR+�=�f�="�W�sK��鵾Z<?7��>Ye�>��<?�R[�/�;�r�4�q�G��a��J->� �>Oy>)��>��*����(����/ž�MD��@6�_3v>�zc?�K?K�n?	S�01�m�����!�C{/��W����B>na>ʶ�>�W����i5&��W>���r����qy����	���~=а2?�!�>0��>�O�?J�?�x	��X��bOx��1����<�+�>!i?%8�>��>!�Ͻu� �v��>f�o?ϛ�>Q��>Q�J�-�$�-9��� 7�b��>���>�U?w�/>.eH�Ϗk��1��8���ג)�Ǭ�=C\?����Ƙe���>��F?�$�<&��;]��>�"���N.��eϾ�4���j >�2?<.�=�{)>ˊﾰ9$�K/��@�3��*?�f�>&����;��?>��3?�V�>|U�>Ք�?UM1>i�M�[=n�
?��Z?4-@?`'?A�>ӭ/�U����8���H:���=���>V%>��m=�>���?G�a�:�4�,=�ޗ=G�I=qTͽ����9 ��qk>=�\�=�~>�ӿ�mC�?9�����b����1�����E��Z�ҼE�Ҿ�]��V����=:���SL��;W������H�G��?/�?� �]�
�@���Po�O���I�>s�;��d ��n�}X�<����߸���d�����7���e��uI��t.?P��𿿼���Ը��U?n?=?��l?_F����a� �5�
��>��U>��->�8�"H��v峿xS��W�^?˿>��F��� ?A]�>�B�=�\2>�(h�C#��U)=<��>�?~N�>�!�De���3���"=��?�F@�sA?�U)�����M=Z��>2o
?
2F>�@.���[�����>R'�?�_�?޿k=��X��5��Nc?�I8<>0A�ۨ� �=
F�=��/=;�y�Q>�8�>����6�b�轺K=>���>������
���W�S�<T�Y>�(��馎�'ށ?�&H���K���� ���>t�G?Pْ>18>�4?ʧ:��<̿�=U��dd?|@���?E�$?7޻��G�>��⾭�F?�{I?�@�>
:0��o�~�`>��R��<<����_�i�y=��>pc>�߽v��ns��O����>M$��ƿ�$��@��	=����Z��)�e����U�����w�l�h�罆p=���=$R>|�>[�U>�VZ>�%W?��k?���>3�>)#߽ϥ���̾���t��Cj����Ӛ����:��z޾+	�Jq�O���`ʾ��0���=lLP�̩���xW��5P�5y�Z;'?�S>L���g����=�X���!Y�xAh=�Dҽ"��=�S���Z�"!�?��??�ډ�j���+�D�\=(���$w?*tz���=RȾ���=~��=(�7=�>�(>�Bھ{�A�!�S�0?u?�þ<򔾦�=�J!�tN�=7�2?u_?���(��>%?��F�nN���Z>H0�=�k~>�=�>���=�Ҧ�5��<8?0d?��j�u���vq�>�;��(+Z� ��=*�>�5�"[�=��=I*�:Zީ�~�;I<3=(�">�%W?�a�>y�)�������/g���>=ءx?�|?8��>�hk?��B?50�<�����S�E7��v=��W?�Ki?��>���B�ϾM@���5?b�e?Z
O>�Eh�ό���.�)��5?M�n?	e?�����h}���w���i6?:�s?�zO����L���L�׽Ř�>y��>b��>�@N��?z�2?��ý���0�ǿ��;K�?C�@8
�?��Z�&�ͼ������>�:�>y���V]���:���ʾ��<_"�> 鲾*뇿�9<�.����0W?�?Z�>������=Vҕ�3W�?��?F����f<i��l��f���ˠ<��=]��A:"�r����7�1�ƾ͹
�ɣ��=x�����>Y@r�0,�>�28��7⿉UϿ���0aо�4q���?Cz�>�Ƚ���r�j�OOu�ӪG���H�ߘ����>QO>:n��{i���p|�e<;��Sf�>� �}��>�V�����F��A�E<�C�>I!�>�<�>)�������ڙ?Ļ��Uο�՞�k����X?�?R��?Jh?	<V�w�a�{�Оۻ�G?�s?�,Z?�,�-k^�+�>��xj?񫾰|`��3� bE��(X>�f3?ŵ�>Ct-�zm=��>���>�>%�,�wzĿL���L��?�?\�?-��P#�>s�?$]+?F\�阿0���r�)��uZ;~??M�6>o�������y;����E�	?�p/?������-�_?��a���p�1�-��ǽ4ߡ>��0�U�\�C��gK�6e�*���y���?�c�?�?MY���"�� %?Я>P����ƾ���<H0�>��>�KN>�^��.v>���;�9�>���?��?�}?t��������>M�}?ʪ�>�<�?�l�=�{�>G��=:���z��'>
K>�7�,�?ZGL?���>��=a�3�#)-��=F��VP��D	��C����>�ib?P�L?�d_>�C�����)#��oҽ�/&��ͧ���=���5�����,>>�<>'>^�?�ްξl�?�	�<�Կ|���c���?M�P>���>�>� l8����=Z?� i>O� ��ֳ��l������"ݥ?`�?�?��־
���=W��>��>�4�=���q؝���K>.c=?s�ڽ!��Zwu��2f>|��?-�@;i�?�d�K%?��]���$�W��n���F[����<�J?(���*��>�o(?x�T>9�o���FEw����>�	�?���?�(�>�tc?2���,��C�ؽ���>�Z�?L�.?��Ľ��$��Ɯ>I��>/\ݾu���#��
f?�@��@�r�?�l��Ģ�?���Bm��;>ž�3>�����=g'7������>^{��z�G::F>��>�A,>]D�>�N>Q,>� >���)u!�Ҟ��Ԛ���=�x��\��G��u�Z����>��8��y�þ�_��.�=�G|�L����
<���=��W?sT?�m?u�?�����o>������|=���
E�=�P�>�0?��I?��)?@��=��L�_�L]��a����q��I+�>�Z>i!�>1�>���>*�༮6E>(�R>�2�>n? >�.=EhĻ�<»J>Q��>
�>���>*"a>٘�=v���f���{���V�<���=g��?���<.�F�����T�K׽klo>d)I?�<>���>GпZM��O?�;�G��t�?��>��Z?T9?�r,=�m�B��@+�>�m��������=2(��6Ӏ��;$���>x?�ah>FIs>��3��9���P�Ȅ��6(~>36?R��<�l@u�ZrG�i۾^�N>g�>#Y��x�9Ֆ�&`~�k�g�i�v=��9?[�?�N��q⯾��t�f���g�Q>;�Z>��=�q�=��M>��d���Ƚ�I�4[1=���=l`>�e?Lk+>/[�=���>�!��i�N�o�>C\D>i�.>m�>?��$?���0����ڂ���,�G�t>$8�>J?�>��>��J��e�=Lc�>m�c>)�Q�� ��@�egV>�Pp�3�\�\r���v=m�����=���=`����9;��g3=*�~?�v���䈿30뾆����D?�:?$r�=�AK<:�"���Y������?v�@�V�?#�	���V���?�>�?��YN�=:y�>��>��;^aL�Ů?L�Ž����R�	�,�"��E�?S��? /�Wċ��l�W>ak%?�QӾ���>�_�ZH���䆿7�u�	�+=�b�>S�G?�x��G�U�*�=�F�
?̅?��𾲫����ȿ�#v����>6�?���?m��~���?��2�>?��?�[Y?�i>��پʑ[����>�A?LUR?�Ʒ>���	(���?�Ҷ?���? �!>ݍ?_��?B ?��=�y7��׼�����IN�)�>��?{t='���Zs�ж���E���AT����p>�z=tn>3�Ҽ����Uq��㉽O�}�H� =��>͓G>�>>�h?��>���>x+o>�ͽ
M��@�{�:l��06?G)�?vk����Z��@/>S���m�\�V?Ygp?�0d��ž$:�>�*`?��p?�N?���>:�>�T̒�&���?��M��<�1>~U�>��>�F�>)��I�Ž�M�>׿�>j�Q�O&��ُ����T>I�;?_c)?�Y�=&(?e�'?ӵ�>��>�41�p���dY�XЗ>���>x�?6�?�j?��%;�
ߎ�$8���/b�(��=+�a?��#?�G�>eۊ��l���ֽM10�Лa<��?��y?�("�΢�>���?,C?Fh?�ֆ>�ت<�
��j�!��=6w#?�6��2A��<�q ���?���>=��>?d=p 9�� �����6^Ծ�?�?L?��?/u���Z���̾�/=���^��:ӷ<=#N6���F>�I�=�1b��!�=�A�=�>�\d�CG�P��<�@�=%{>Ȁ>Co"�7"&�K4,?_CC�
փ���=��r��xD���>��K>l��k�^?�O=���{����Xr��{�T�� �?"��?nd�?�	����h�'==?�?�?�h�>�]���q޾2���w�ǹx��H��w>��>�o��i�Y��������B��x4ƽeF4��#?#��>[5?�w?ؿ�=�?�>Ė���7���ھ�����}��%�u_0�b7��_�����'E��綽j~���	���"�>��x�Ff�>��?�>���>#��>�7
�\�h>1�d>X.�>�#�>�;J>�r>��=�vƺ�8�fE?�龔�/��۴�����K�e?Lw?:D?]Y%=�&��F��{�3?*��?	��?(�.><o�q�#�v��>�k?�W����>��f������}>O)�����L����5�e��>��0��7��c����
�>i�>�)=�������n��3�p=cJ�?� )?�)�&�Q�!�o��W�&S�2p��g�K��B�$�.�p��菿�f��5��֜(���+={*?��?�{��������k�(?��|f>�*�>��>�ξ>R\J>��	���1���]�:;'��׃�O9�>�-{?4{|>�,W?z�O?XI>?i N?�2�<
[_>�U���@?d�>h��>�>l�!?�?��&?.L?�J?Idt>��s�8	�"Ծ�� ?r�-?�F�>�
?y4$?��ݾt-q�_:>w�=�E����`;=�򘽛�����>v��:�ʝ>*+?�ξ�XT����݇)�P�I?n#?���>h�~����߽T?�1?��?E�6�Ɂ�z����W>\.�?3m�#�>���>�B�=�[�͒={�<�H��#>�s�;���=�D�=߲9> 2�=�ו=w��=	�5;S&>��Ὅ��>,w2?�	�>���>�Rӽ��
�t�Q��R�O|�=��x>k��=��	��
|�~ϧ��Ei��&�>��?Qܩ?�<��k9�=g�=c:ľ�<�T�����R�">j��>Ru�>�%=?� �?�S?��>�q=��c���@���k/�}�A?�!,?�|�>���v�ʾ�73�F�?�Z?6a����i5)�~¾�Խ��>�\/�1~����SD��~�����U�����?��?�A���6��i�ӻ��eJ���C?0�>�c�> �>k�)��g�%�.;>���>NR?� �>��O?�={?M�[?�rT>ß8�0���љ��02�'�!>�@?̯�?-�?Ay?�s�>�>1�)���XV��A��T�kڂ��=W=�Z>-��>-�>�>-��=*�ǽ�C����>��j�=�b>w��>=��>��>0zw>;��<��G?���>2[�����褾ʃ�T=�˜u?؛�?�+?�t=(����E��F���I�>9n�?O��?�3*?N�S���=<�ּ�޶� �q��%�>-۹>�2�>���=�bF=�i>�>��>�-��a�7r8�tGM�Z�?)F?���=-	п6nk���dz=U>2F��˽H�������j>��H�2S��䊌�����񊾛�c�BU��mB�������l?�7�<��A<��>�8������S>���B�<='T��=�ɮ���=�_��,�<A����:�=��ƾ\�~?�gQ?7�/?��D?�':>��>w�R����>�;�;�!?SwK>ůo�?���C,!��	������׾/�ܾ+�q�A-��v/>��	��N>��H>�>G_!��K>���=�g�=�o��A�=��=�=!#�=%d>��= �>�)r?�vg�����<�8����+"?�>�q�h�پ�([?� �>z�Ŀ�
��#�?q��?���?��?�Ǉ�p�>��s��ܻ=�C�=�	����]>t�=w�#��?��1���>����=�9�?� @��A?B皿�\ۿ��,>!k?>.�>�R��74�?zW��S�;3U�Z�!?�o5�Uξ@�>/��=;�۾0���_�0=��1>Y:8=b���p[�r�=R�s�-�B=�r=���>I>0��=%���׼=��<=?��=�pH>��ܺ}�(�r�Ao;=��=��]>�!>���>��?ia0?UXd?6�>�n�Ͼ�?���G�>�!�=�F�>4څ=�mB>���>��7?�D?b�K?���>׽�=��>��>��,�۲m�&j�kͧ�M?�<��?W͆?�Ӹ>��Q<O�A�}��jh>�?6Žv?�S1?�k?��>a����ڿ�¾���~C�=v,x=�O�<���zZ��Ii�C��O�j=�<�=���>Ȗ�>�y�>X0�=	>��\>Ӆ�>���>!T(>^ڈ>P�=TWR>wN>r�X>`!�=�E�=��=�F4��Ά��잽u�=5<Ž�ҽ�Q��ͽ6�=&�?�=Q��>��7>Lwྻky>{�ھ�_�`>��	�g�g�X�t���g�˄+�c����}>k80>UM��╿e?��>�DE>�C�?-VJ?���=�R��.4���2���f<�྾Q�=N��=|?ܾ�<O�u�U��lN�����s��>�m�>��>w�m>��+�E�?��Jt=�pᾶ�4��d�>ꊾb�����Nq��2��_��I�h��hź��D?���7��=�^}?iSI?��?C�>P����ؾD.>�&��v�=y���+t��i��3?��&?��>PJ뾻kD�Q�Ⱦ���8A�>�(@�e*N�M�����0�
�t����A�>ü����̾X�2��چ��/���FD���h���>?�P?���?��a�	�����N���
��q�y�>�zd?+Y�>��?q?/��K��*���$�=-�o?&�?�??h>몽=C���8�>�*	??C��?��s?{v?�=|�>��;"� >�����Q�=��>w��=�%�=�q?U�
?F�
?�d��d�	�Z�����^��c�<�ߡ=�>Xk�>x�r>l��=+�g=��=�*\>\؞>P�>��d>��>dT�>����¾a 2?�{V>���>'�?�7z>�Y �$Â�B��=�3W=����������/Z�=�=%�0=�S�AM?@ؿ�V�?~rw>�d��pN?[� "$�;p>���>�Ƥ���3?h�=)	>b��>��>�0�=�{�>�#>W8Ӿ�h>����g!�a0C��rR��ѾK�z>����-&����L���"I��_���a�4
j�-��4<=�-��<E�?�����k���)�������?1Z�><6?�⌾B%���>��>���>�C��c����Ǎ�W`�B�?���?��/>II�>s �?��-?O��;��r��`�e���T��&&�?�M��w���7����=�TxO<,�?�&w?6�y?n���Z>%�?��$�-���}5�>��Y�V�w���=1%�>�'��gf���0���*����=�@Q?XM�?��?Tlz�E�d��+>:?��/?�Ss?�p0?��9?�Q���&?x�4>7L?k�
?'z4?͌.?�O
?;]2>��=����=�1��`4����ͽ����w��ٻB=���=��So><hU=�<����횧��6:;L���<t�<%I= ��=���=�4w>��v?��2?�i�>�b?�?���y���쾃��>x��=�l׾|%�+ϐ��,��dF=U�?���?��?�ʽo���U�)BS>�D�>]�=4F{>�u�<��	=N�Y��Ri>N�=�M>E&�=�z���ջ��9��8R���5�0
�=7��>h]�>��%	A>F�žsu����>ƈ���<���al�ԢD���A�[P��5�>�t?��8?�'>t�������:�}�T�W?�N? �@?�ڍ?�Ľ4;��gs?�S�w��0C���>q?�\
�����������L�f�G=-4u>#ɔ�B=���c>m���ou��aJ��8޾p�=�	��W=`Q��Ͼ��k����=nb>wҿ�߻�>G��(:����M?�Di=O{���^�1���8�(>P��>,�>�O�?q���;>��U���4�=��>��?>ٷؼu��һH�M��(�>d)E?��_?~Ʉ?�8���!s��/C��- �C塾j�ӼF�?�>!$?/?>,#�=,v��3��4'e��F��3�>���>[���G�8�������ٹ$�$�>t�?�� >5?�GR?�
?�_?�)?ƽ?G2�>�U���7���B&?㊃?��=($ս��T�<9�MF��&�>�)?��B�U��>M�?B�?�&?�Q?ծ?#�>® ��G@���>T^�>��W�_���`>r�J?���>�:Y?}Ճ?8�=>\�5���X}����=B>��2?o7#?��?儸>ݩ�>������=���>Dc?�0�?8�o? ��=�?�A2>Q��>��=���>_��>�?WO?=�s?N�J?��>���<�5��6*���"s�3�P�/"�;��H<��y=ni��It��Q�N��<�F�;�W���������;�D�����x�;�b�>��y>z�����@>��Ѿ����<6> :I�����3n�L
�D��=D�d>���>�~>dF�G1=�k�>S^�>Ϳ���)?��?hG?��
=��m��8���x���>�TH?r�$>X�d��E���^}�,��<��^?B`?��0�ZD۾�M?��V?�W���$<����#t����Ⱦ��{?7��>�=ľ�l�>��?�/i?6��>��c�5Gm�Ǘ�~jL��@��>̱�>�V��A��M��>�`Q?S�%?ȥ�>�L�>}j��I�h�`;s�}m"?BV�?�l�?��?<�3>�A����_+��J����]?�i�>Χ�M#?8'���о鋾!����l��k������j���'d#�<����Խ��=��?��r?Fxp?-v`?U& �*�d� �^�
����eV�A��6�Z�E�b4E��D�1Bn���i�q�����\=��i��C���?�='?��*��>�R��Q��Cپ��d>EB����սG��<��r�³t=�Ĭ=��6���������IC?m�>T0�>|�??�Y��<A�|=2�wOA��x��Ţ>���>�f>���>�!��,��U�	ľ5�?��Y����s>�Dc?�L?͑o?�����1�����K#�n
G�,{��=@?>U	>9�>c^���"���&���>�ps��������&�	�O�=W�2?��{>m��>���?��?�(	�����!v���/����<��>��f?U�>&z�>���� �u��>dQe?��>K��>��F�B�*�k�{��|����]>c��>���>g	
>�Ņ�U{�f����Ꮏ;�?�M��<_?cQr�,�N�~�>�V6?Cz:��9�=IA�>���3U4�h�������>#�1?���=���=\ �.q$�@�}��,��ߑ'?�i?yC���G&��{Q>��)?�?�:�>��|?�բ>M�ľ�*=��?keV?<�M?�6:?���>��������������Ux�=���>���=,�<�v�=:5%�w�$�ys7��N=P��=\4��)�� �������i=�p�=�D>��߿��L���޾0���������+��9���1�`�Ľ=�ɾ�:s�{�Ͻ��j��V��EjA���m��/˽1��?���?�"־����ES��jɂ�񌮾1�?��-�g{Ǻz�;]U�6M{���ƾƩ��*���E��倿ԠU�W "?@#ؾp��ٲ�pwľ��>?g_?���?5�!�(3�I�0�n&�>>�=7�<=�оė��쾿��Ӿ
P?_'�>9��H�I��>�O�>Ʌ@>R�d>>0���K���z)�b^?�?�P�>Cb�y�ο'�����<A��?U@�{A?��(������U=��>\�	?=�?>�E1��:�]찾T�>�:�?���?0L=��W��G
�L}e?��<��F�2]ֻ�m�=#�=��=3��W�J>7]�>,s�aA��%ܽ#�4>y�>b�"����^�w�<��]>��Խ픽b��?A�Z�/�1�����F}�0�$>��1?��>�[�>�?47M�3VȿGI[��s�?*�@��?~�$?�蔾؇�>a8ᾐ�@?��;?��~>i�4���n���=d���iM=:��Y�ޗ�R��>�{+>�8���k�����<�b�=����Eƿo� �1]�/��;�����/�X[)�+�½��p��E���p��X{�]3�=���=��Y>{�>�7i>�xp>^�\?;k?�O�>=&>��:��^��;����f=�=��>𽼦������������)���A���������C�/��=�S�[܊�w�^��Ti���.�6?���>����Q��*w=p�h��a��1_�;6������;���R�^k�?X<A?�ׇ�qY������v=����g?*����ߠ�Q�>u�n<��=���>��»����bJ��b�6t/?!�?"�ľ�Ǒ�K�>����9��=��*?�?|�b<��>ܧ%?���s���k�i>�H4>6	�>���>��=f1���r˽F�?BT?�n#�����b{>�ʾos�v�=�P>�(�I ����7>Wx�٩��,F;Rh��9E^=W?d��>�*�5��5���W��'?<=x?�X?_|�>�k?5�B?�4�<���X�S��J���t=a�W?�Pi?��>����о�ʧ���5?�e?/�O>�g����'/��t�F?9�n?:M?Z���]W}�^����a?6?�z??:\�dS��]�Ѿ�����q�>�o�>���>��,���>�=@?'?���䒿� Ŀ�c'�v��??�@?�?�c�=���T��;Ι?��>�Y�W7��\��䎒�t=⼰?P勾\����(=�YG��^?��?��?o���[Z�1��=�ӕ��V�?�?������g<z��Tl�pp��`ڠ<�ث=>���q"����$�7���ƾ	�
�'����~��>X@TC轂5�>�68�\6�1TϿ����_о~Fq���?�x�>��ȽQ���u�j�	Mu�W�G���H�͗�����>��>'w��_8��Z�{��;�␔�W�>�R	�eT�>	�S�|
���ޞ���%<:x�>OH�>f�>�	������x��?�����ο�����@Y?to�?qU�?k\?�|<)�x�)�y����LCG?
�s?�*Z?8j#�]�o�B�R\?z���tXk�J81�P	M�N�>h1?��>�o+����;��$>��>K��=��$����k�������?[��?�I���?�{�?O�;?���������L�2�oV��h??�X>��Ⱦv(��8Q��v���>��"?���+� �^*a?,a��l�~A+���ʽ�,�>`�&�fBT���Y������a�EG��?ք��֭?u��?�S�?�\�	���b#?HD�>Q}��~����x<��>{��>ƀ0>M_��4�>����/?�)}�=v7�?Db�?2?}��������=�|?[��>�E�?�\�=:��>Л�=����]���;">2[�=C>�J?ÅM?Ϧ�>���=4�8�c.�y�E���P�!���oC��T�>0\a?��L?��d>Ku�� >5�נ!��˽X,�#�¼0�?�H�2��/�7<1>8�<>��>�?�
Ͼ� ?���-�ֿ�m�����z�1?���>*� ?����!p��;��%a?��>h��줳������սO̬?��?�v
?-}޾�]��D�>զ�>Vy�>7�½%���A���<>'u>?����Em�E�>�#�?U�@fv�?rie��s?������;`��̾�*���>j�?R�u}>�@�>�[>k�X����t�x��>c��?6f�?ׁ?dm?Fy�9�(�Mm����>Al?��?�=B�N�`>�3�>D�⾸͇�o��V?��@?�@��f?$ې��-ۿFܜ�Khg�F%e~>]~=�>��޺�J>�\M>Q?��/X�=�&k>�'�>P(`>>`<>J�5>2X>>1��=P&|��q�t;��ꮄ�_s)�%���۾+��L&�OR����H�聊��%����� ��m�h�Q��I-���Q����=C3W?��R?Uo?AJ?q����6">�����C=y{!��2�=	��>G.5?s�K?o_*?Ai�=	����b�7ǀ�����!�>��K>��>���>Px�>����JXF>�f:>0.�>���=g�B=�Z���=�GM>_ԫ>1��>Ii�>��>K�o=;Y���G�����"����ּ=P̣?iw^��"/��荿�寽4q��I/V>�~/?͉�<R��lY̿�����B^?���m����U��Y��>:\k?N?}�&>����Լ`� >],��0���Z�=����Bݚ�}$*�v�8>��?�6o>7t>�4�� 7��M�F{���a�>Q�4?����
*���q���@�!bϾ�P>���>�P^��! ��]���m}��je��D�=Ti8?L�?{���J����p��ϝ�2R>�)O><�=&3�=��P>��z�������R��:A=l�==8f>��?�8>��s=w��>*Μ��V��Ƣ>�o">ǰ>�@?_)?]����6��v���$8��nd>D�>�u>i�>�K�r�=s�>�]o>����޹�����D�]�^>&�X�uD����M�P=�mý��=�7�=�+���
�Q*O=�~?���(䈿��e���lD?V+?� �=U�F<��"�B ���H��C�?p�@m�?��	�ߢV�9�?�@�?��G��= }�>׫>�ξ�L��?�Ž0Ǣ�ɔ	�)#�fS�?��?p�/�[ʋ�9l�~6>�^%?�Ӿ�:�>#��1���T����t��s�<k@�>�gB?-�
��HJ���	�� ?'��>���2��^�˿�bz���>�*�?$d�?�i�<���QN�� �>r��?Two?|��>�d��/������=HN?݆X?���>����l"Խ��?��?�_?��>Oڈ?W�v?.?�����*�������e�=�[���a>��=+����8K��̗�F����4c���,�U>(hT=�ǌ>Hq���^�kb��06ӽ�H��a���f�>�>n�k>��>h��>�/�>�4>G��9�[]�������y��RC?��?��þ��b��<n=2���ܜ(�(C?[k?�KU��E;�ZJ�>��}?�Ì?{�N?���>��������,¿{����"S=�>��?Ҍ�>M���	7�>Q��N�ս$s�>��>����p�Y�����$�G��>J.?	?�F>��?P(?z��>��?P�C������`����>K>�>qz?U��?<�?�����hG��ؘ����~�W��G�=���?�?C�>�ˇ�����.�<��<Z��<tI�?y�R?�yf�Ó ?X�?
�.?��F?��>?���X�쾽�\<2�U>�?#ҽ��U���R�-z4=�FT?n�?7x�>mL����r=LG�=�c��<a�]??�s�?e/?K]*�s^y�m 
��	�=&Ì<R��=�6�=C��ȏ>��=��3��;�=~S>�7�=�߁����#��<�>�=���>/��=����H�=,?��G�ۃ�+�=:�r�UxD�s�>,IL>�����^?�l=��{�����x��]	U�� �?��?Ok�?���'�h��$=?��?\	?7"�>�J��@}޾I�ྤQw��}x�0w���>F��>��l���]��������F����Ž�)���?���>�E
?B`	?l'=>|��>tǟ�6�(�����@�ܓm�k���d6�y�$�����ҍ����n��=��������>������>��?� c>\"�>�}�>��&��$�>��~>\~l>��>�i>�V>K'
>dr�*����N?��ɾ5�/��|�4!��7<G?>]e?�_�>���������# �P�?�R�?��?��S>��j��k/��y�>e�?���{	?�0�=?̊<F�U��0Ⱦ��2��5��"���T�>�Ľ�:�6N�o�����
?�x?|��N;�aɽ�u���|�=1�?tKa?Ӆ%��a�p|��q��1/�|?ܼ�] �=�����	�Rw�XØ�h�ro��7�b��=�� ?�e?�a��Y��G�����x�Q�8����>X�>��>� ?=J>hV�Cx-�pKA�G"���Q����>���?�,j>%7q?�+F?�B?.H?�=4<�>JXG���E?�@=O�?9��>��^?�?��?<�?�?v�>����w/��*����#?s@?��?Z�?��>�ֺ�)�K���=���=d2��1�=ţ�=`8=L,�Ԭ�A��;֑>��?y��3�h�]��|0>��k?V5?6�>x���˾s�W=���>�a?��?�d"�ʒs�*� �.Y>Fq�? <��V}=��q<"�9>�)�a�Ը���=��`��d>>A� �F=�"���<]�=��8��Y��������</x�<`{�>E['?���>�4�>���9e&��N��qռ��>��>��X��(��颿"�����i����>�֐?J��?����&-�=��==[���"(�F��5f���	�>>g�>�K�>f<T?/��?�Z?�?�(`��r�c���i�����1%?��#?2܏>:���µ��⦿�c'�d�?�X�>)�\�좝��P��붾|w�"z�=L�-��&~����LE��B�=^�̸�a8�?�N�?��ļ�I����Q*��E긾�O?���>��>q��>W;�Je�[;��I>���>nOS?��>I�O?!{?;�[?KT>��8�#���ҙ��1�`">3@?���?��?��x?XD�>Ɇ>��)��྇"��+��*+�.ڂ��VW=aZ>�f�>��>�>Mo�=�ǽmޯ���>�暥=�<b>_p�>���>�>�>�x>eů<��G?���>0_��ّ�䤾�Ƀ��=�P�u?͚�?r�+?@�=`|���E��R��v<�>�k�? ��?�7*?�S����=2�׼d㶾��q� +�>��>C7�>��=�F=Q^>���>3��>� ��_�Ao8�x#M�d?� F?û�=nƿ'�q�+�p�����e�c<������d���1[�ۮ�=����#��Z�����[�磠�f{���浾����ޜ{����>P��=%E�=��=�m�<Kʼ�'�<K=��<4�=��p���m<��8��	л�ň�i��:v[<�AI=����ƾc��?��G?ћ&?��I?��V>�d)>��T��+�>D����#?寿=��h<vt��z���q��bC�����;y���v��T���=>V<a�,09>4g>k��=�E�<A�=�q�<&x�=k6=�G�=%��=�<w=;qP=m*�=��=�p�=!+}?^��`�����.�49���]1?��>h�=�U��@�d?;�t> �q��w��u�D߃?���?bW�?��?_RH�x�>Đ��T��=��>�5V���j>�?<?��i�>�Y�=��&�9����������?��@�G?6?���ѿ
�>��:>d�>�S���1��[X�IT�t�O�E!?�:�X!Ǿ���>q*�=�9ܾ+�þv,_=u�8>:=� ��\�$M�=KCs��<=��=0�>��=>za�=6��駾=�H=/��=�}S>۪<��2��<���1=22�=l�g>��%>V��>�?:/?F�d?qI�>��p�y�ξS�¾�Q�>�7�=�n�>M��=��?>ӕ�>)�6?vuC?��K?י�>m�=壻>dܤ>{�,��]m��n⾖m���/�<�|�?�݆?LƷ>}%><�1@����%#>�m�ƽ�d?s�2?
?mɞ>ޮ�w9꿗���W��t;� F���=aK���a��=���������=>�2�>��>{;�>ז�>�JL>6't>.��>M�!>�(�<�=O��jn�:0�c=)4��G�9g�W!ͻJ��+����;)i��ތ=�<[�N�V=��=Vt�=
I�>c/>�H�>SP�=�α��y2>.[���xL�L<�=MR���%W�e?\�Eaq��p��.!�~�U>�(v>��½(����?]D>73>��?Gm?�r
>������u;��U����)_��μ=���=;`����<���S��3F�/Z�;��>�n�>H*�>��x>H--��0<��z(=p�C�6���>r�h��1T��#��q��آ�:�����g����:M?ƻ��m>�{?Z�K?���?/�>z� ����>-I��%�=?�-���<����?�??,��>�"پ4�8��n������&~>e9n��(8��X�� ��۽���ț�>�Z�Y����'�(���,��):� 3���>��L?g��?	��ީv��ZP�=������N	?�}h?j�>��>�1�>����Ȭ�w�����8=��b?E0�?H]�?��>P��=O���<�>*	?���?7��?6s?{?�!r�>Ռ;
� >s���v4�=��><��=3�=�r?F�
?��
?Z����	�F����^�2w�<Rʡ=,}�>2j�>��r>���=�g=���=�(\>�؞>��>��d>=�>xO�>�ό���W�J?>]o�>=?��]>l�=R'��@�L<�7��������B�;���M�u=�>>]��=�Im����>QDҿ�~�?__>G���c� ?����$�O->�t�>뙾75?��4��-�>�5�>���>��{>?��>E��>�Ӿ�>���7�!��(C��?R���Ѿ*�z>ľ���%�b��ޟ���I�8Q���F�j��,��-K=�?�<�=�?nh����k���)�����6�?k*�>]6?���8,��!�>F��>W��>I��S�����!V�g	�?���?��M>`\�>�ۃ?�M*?
dO=dX��v�}�O���f�6Ӄ�>�g����7Ԁ���ƾ:�E���?y:�?z��?���� (>��?p�M��݊�eW�>��d��sv��_<���>Z��Z����E��'��;�)�^?Yg?�'?�پ;�w��?B>�@<?"1?�s?�2-?�:?{�	��1,?��8>1F?�y	?�<?)4,?��
?D=0>�)�=��L�� =qʢ�wb�����b��U����^^={}=��׻{�<���<w =#D��j�u�;�q�Z�<jIL=Z��=1
�=�Ӑ>�_?��?�Z�>�;]?�虾�v��󺾥�"?����D���u	�O(����辧����?��?�]t?���;�5�:7&��ؙ=�ۂ>5�>�*;>ⱎ>KԖ�n��Rw^>a��=�U>] ��!��K��:�+�d�d�7�2N�>Z8�>��y>y&�+�0>�㾒�Q���>h�s�3Y�����X�4��j2��7Z�3]�>�H?ԡ?�^�=_i���R���o�@R?;�-?0�V?Us�?`�c�0�ﾯ�B���w�v���?~�{���]������QU��Ù=�`�>5,��n��Yh>�-	�8�۾A�q�XP�"��F�R=�y��;Z=#A��pоMXn��T�=�B
>��¾n�"������쩿D/O?B�=G��lY\��e��C�>�@�>�C�>e�����$�@������=���>��D>���v1��F����lY�>�E?�f?+1�?`.��!?o���E���6��.��;R�?�>�S�>��>@�y=ź�����uj�� B���>���>]��V�G�C���(��=� ���>��?��?>��?<�T?�?S�a?�(?#?[{�>3b���\���A&?��?X��=��Խ��T��9�F�f�>�)?��B�t��><�?�?>�&?3�Q?д?X�>�� �	E@�ϒ�>.X�>�W��a��d `>6�J?ƙ�>g;Y?Kԃ?��=>��5�뢾�ݩ�'U�=8>
�2?i6#?��?T��>_��>�����=��>�c?�0�?�o?���=D�?X:2>���>4��=Û�>\��>�?>XO?/�s?��J?ԑ�>���<8��_9��Ds�e�O��т;�tH<��y=���2t�UI����<��;g���J�����'�D��������;U�>��> ����W>��þ�\��JN�>�[ ;?!���F�t��O�=O�>T��>;�v>BX�W.n=uͱ>��>�`�~!1?��?z�?:/�b��x	��FV����>�OG?���=J^S�Γ������I=cV?�wj?E�"����5Z?$�S? ��TK&��W���Ǿ@塾fd?�b?DȽ��?EL~?�a?�`?�2���LU�O����5Z��kf�l�=�0`>�w"�<u��Z�>�l?]$�>�L>D>m50��i�[���{�>���?5�?�w?>$>; Y������s��c����^?\ �>*9��U�#?+�0��GҾ C���q����ᾪ����E���������� ��Ɓ���Ƚ̺=�3?�q?,�r?^�_?�W��d�c_�qc����T�����\�8:E�D{E�?EC��dl�Þ����a��21@=�D}�h�@���?��&?`Z(���>�J������ ̾"3F>����{|��<�=t����I=��b=��e�r)��έ��& ?p��>؃�>�=?�(]�M>�_G2��8��v����.>���>d�>av�>�v��C*���޽kjȾ�?~�UgԽf�u>9�c?�K?7�n?E6��1��y��Y�!���2�_=��ϢB>�>̓�>5 Y����PO&�)t>���r���� W��e�	���={u2?vԀ>Ƞ�>�)�?9?<	��ޮ�v�x�21���<��>~�h?��>۷�>�%ӽY� �3=�>��n?[k�>%��>yi����p��J���>�E�>���>+�<>�,�ߜn������S3�T�=J�X?򾉾�2M��n�>0�G?h<����<:ױ>�����)�:�����0�f>��?sX���v�= �.$��C��/]Q���(?:�?������7��J>�5?�'�>N�>��?v[>J��B�<�?��\?	�A?�31?���>��I�-Y��"l����7�(�W=	��>0[>�6:=���=��ƽ��]�t�;��隼��=�S�������u!Q�M�<k\�=A3>�)ڿ�:��-��
H��^��v�#�u妾u`,�1n�<@�4.��������ҽ�=���d�:3�����w���������?~g�?V1���a�Z���nO��C
�Ռ�>�������;�[��x3i��H4���ƾ�����2��#M�Ua���c�ei'?�ɒ�O5ǿx����޾(�"?ǟ ?�_{?R����%�"�9��D&>�:	=�}`�����b����Ϳ�Л�S]?{��>��v���>���>��M>.:x>�߂����^�C<�[?k�,?e��>�o�X�ȿT󺿘q�<�?@�7A?:,(���a W="
�>@{	?9jA>��,��B�]į�.x�>-��?��?�I=X�z��?�d?j?�;uE��Żb^�=~̠=	�=�F<J>,=�>���?C�?(ڽ�~6>C8�>��#�;~�Ҹ]�j(�<"�\>�ֽ>����ׄ?�z\�9 f���/��K��vX>��T?�	�>ᗡ=#�,?�9H��uϿ��\��La?�5�?��?O�(?沿��Κ>��ܾ%�M?�S6?��>m&��t��,�=��߼+�����m2V���=���>��>_c,�ؗ���O�*Ɨ�"��=�$��Vſ�p�"���D��e�e熽�!�����X�������v���½9),==�=��W>��k>D�|>��S>��T?�t?>��>,�->c��5^����ξ��j`��~�#���Ȥ�06��'�����>�����"��lԾM�A��X�=p�@��V���$6�>A��\�J��`%?d�0>vB��L�D�=����ͩ���ѻ���7B辴>�G�k��^�?u}B?�/����T����+n���?¼�n?<ߡ�����k���@>3�&�e�|=4��>����,Ѿ� 2��&F�-0?H?)����폾�#(>�% �M=�+?�� ?�j<��>��$?6)��n���T>8o->�P�>ǋ�>�B>�6���Kؽ�U?U�S?@� �����T�>Ԙ���<{��p=�>��4�Z;�%V>B�<����q��U،��G�<8FR?�T�>��-�������1Ź��i�=�z?*c�>�;�>��f?�_C?M�=x���2�[��p�s_p=S�C?�{?>�>�����;�=ľf�:?Mb?M��>�p�r�߾8#4��s����?�d?d$?��Z�zFn�$쐿7���K�*?��y?�eW��Ǚ�b4��0i�'��>���>F��>�=��f�>��9?>u������wĿJ2�@_�?�@W(�?#�=㳚;7<�<���>�&�>R\$�Bݧ�S�|�t'���os=��>�1��,����h0���:�{�[?���?%�?h���v�����=Sٕ��Z�?��?����Cg<.���l��n�����<dΫ=8��D"�&����7���ƾ��
�&���3ؿ�z��>1Z@1U��*�>WC8�26��SϿ��b\оZQq���?[��>>�Ƚ!���;�j��Pu�Q�G�H�H������>ߘ&>ٯ�6U��|N����=��3��A?[�=L�7>S݇���A�¼� �<X��>~�>�>A�a� ���k�?]�̬ڿ]ߤ�H%;��?]A�?�?e ??L��O�����Vټ��F?Q�b?�@?��<"'��	t=��_?���@]b�(���O�?�V>i7?į�>�[%�&#�=��>���>��O>w�#�rN���������˓?Z��?<龓0?�2�?B�@?���������t5"�ńн�^?�>[�G����N�m1��˂�>�<1?�m)���ﾳ�q?�_� ^���?~�;��>����e�����=]�佇TL�$8��6���-��?>\@�s�?����4�?d�>���,�ޚ�=��x>kތ>�5�>��Y��>��-�5N���.>�{�?n��?C ?�ט��m����O>�(l?�I�>��~?rmy>m��>ѫG>�R	���;]J>S�>�	�<��?�=?-��>�p>���we�q0+�,�O��@�U1A��|>"�W?�b?e�V>yB�����~�K�8�Խ./��h#���6����������ݴ=nqN>& �>	��<���M�?J���ؿ�O��b\'�o 4?w��>��?���}�s����n6_?��>!d��$������Y���?69�?:	?��׾�̼A>���>b�>Mս🠽ӏ���7>�jB?w_��:����o���>���?��@�֮?��h��?\��pA���+d���Ծʹ4����=�%?>�����>���>ji>�]|�絹�fz��z�>���?�p�?��	?v,n?�{��p#�V
�����>��k?�+?b^�P� �Gd>��>����ǀ���B���T?eA@fy
@��m?���vͿt���Օ�]���1��=Dx>��1>ٸ8�4��<�YV=�B&>}@.>��>�Ks>#R�=8�G>�M8>G��=�ʶ=~�{����(��H���G�����A�i�i�J:?���:����z��J�E����&�ü��D��Sm8��Y�<��=3�U?�Y?�.k?/(?oY�`>����*��=�t��*�=�o�>�(?j�:?Y!?J.�=4�����_����Q���;mh�V�>K�>�k�>��>(��>`���a.>�:i>�ك>ɧ�=W�=*��� �����V>��>P2�>9S�>/�Z>�L�=����!����t�TF� ������?���J�X�	 ��E�%���|���>&�*?�N=K^����ʿ����O?H�&�q|��D�><e?�sN?>V-&����G>�3�j�g�'�+>�+��b�����8>�?ppi>l�r>g?4�#�8�"�O��d���׀>�N7?����e?���u�f}E��۾��M>܀�>����}������|�Jg���s=��8?o_?PF������s�g|����O>ЀZ>��=>b�=)�J>�|d���Ľ�H��-=p�=�3]>��?'�M>�F�<<
�>���Іl��>�>��>>l�>�\D?�+?���W�ֽ*���D`S��<>þ�>~�v>7�<>i�6���=���>�<>Ǫ�)z���%W��YQ�CK>͋���S�{֕�tÏ�5���=�=&��=������3�=�.�?&=���[h��,ɾ?o����2?ga"?9��;���=�?�����8��Wh�?	@�l�?�iȾ$�L��H.?��}?��>�)>4�?�ԏ>�H�	�E�W^?!��<��s��s������7�?B��?K����u�Krp��B4>~&?x5˾���>�'�d��ot�vjo���=yZ�>UYK?!W�mX/=���>?�k?.������r�ƿ��h�`�>�	�?(�?��l��Ȕ��R�[T?"��?�5c?�':>��ɾ���?�p>\�6?�a>?�W�>h�������>�f�?i�m?4=#>�ȏ?���?�?��l�+�&��̭��쏿=@���<�2{>��=�߶��i^����������Un�!�U#(>�`=�i�>Ғ�r���΢=1%d�܅���g=:��> �>!.3>G�>�/�>��>�x>t����'�G¾�hg�лI?j�?���^i�K�A=���8VNU��-
?Y|;?.5ּ�N�����>�aR?�4�?^�X?��>%���ᚿ$�Ŀ!�����<FPG>˙�>��>���Ę=>C�㾏-5��S�>G�>�2���ܾm����I<֛>}<#?�>��N=U?�;)?���>��>�;���F�D����>�"�>9?� �?��?�!��;�.�d��`���W��k�=m�f?��.?�0�>Y����T������*�t��=�x�?���?�*��m!?�%�?�@?�GQ?K�>�OļB������=��.>�� ?,�
��G���,�<�P�?��
?ZW�>�]�v��:�����u�?{�K?�?xz��c�೯���=o��-�;p<�@�;4">�z
>��]�{Ӽ=��>�;y=*�g��"@�*!<�G�=9!�>X�=ʾ#�����g7,?Y�D�'���8j�=}�r�vD�Ȅ>�L>$��E�^?�d=���{�.��`x��tU�X��?��?�g�?,��қh�=?��?5
?4
�>�>���T޾��?Fw��Lx��j��>���>c�n������Ο��J���Ž��
�?߼�>ݥ?4�?.e6>*��>ȇ¾uJ1�~ܾ�Gﾙ%p���
�Չ2��[����U��Y��žģ��ڝ�>����>É?c3>�>�L�>y�/ǟ>V�u>�<>2-�>�k>�>ͮ�=��~-��A?�6N>����_C�wZ?�ހ?��??4�j>�Z��@42���*?��?���?�U=g�z�y���Ƥ>�`
??Ln���>8=��<>Z��:	�-ʅ�ٲ���t�>�̼v��� ��{}����>�X�>JzF��g���#>>���x�>��?ءE?^W�8G�@�t���V���R��;h=�X<� ϖ���%��z�{���K�����v�d�?��|�<�62?R�r?�|������Uo���f�.�/��8�>j�?���>���>�Ս>���N	�eg�W��{<J�h0�>p�z?���>�J?�@??gR?M?a\�>H�>hi���T�>F��<���>��>aX8?�(?<�+?g�?��*?�JZ>7�<���mӾ�?h3?�?2?}6 ?ᓾQ�ǽ�4G�ٻ:Ɋt�AG��ZV=7o<�n̽�7���=۫j>�?�����LW�sb龵>�<k�1??*?'�,?��P�s��7��:?P�>Td->(���|a�u?�Q�۽;�T?�{����3=sq>��=�2ʻ��9�nE�=i#ͼp$�=\/���}�"&ڼ�QX=���<���1�|�4<f<>&U&��G�>�1? I�>���>��1��I���3���8�R>�=:S�=�a�I��.k���L�g�>~E�?#$�?7ϼ��=�
�=l���QIw�J�� ��{zn>oj>_'?|�\??�?�\R?߳?'�ٻ���7������k��$?��*?/�>̾��5þrH���v0�M�?�v?`����P'��g��©����>F%2�����w��g�D���<�����O����?��?][��To6�Ӕ�{������/J?�z�>/�>y��>o�-�͓g�.��1B>R��>8�T?��>��O?�A{?T�[?>�T>b�8�/+���Ι�@Y-�7�!>'6@?���?��?�y?�e�>��>��)���Z��M��`�C삾�V=�Z>���>]�>�۩>�{�=Ƚ诽y�>��X�=`�b>�}�>���>��>Φw>B��<b�G?m��>�l��q��᤾߃��Y=��u?���?�+?�=�m���E�Jp��F�>�Z�?���?�**?�LS��.�=Hټ۶�r���>�ι>"��>>O�=�)F=��>���><��>�o��r��f8�y�K��?�"F?���=�oƿwNs��-r�2���tOR<�����d�}Ș��`�;�=���H��x����Z�3נ���� µ��|��^y���>� ~=�E�=��=$�<ꆿ���<<�M=���<�=�0o���</��˻L�}�3�":хe<�jD=�@��[9;���?��U?Q7>?�T?�R>9,�=>v��,�>�ѽ�G?`?Y>��-<�֝�<�A��5��K�b������>޾ON�����]�r=��}�6A6>r�>T��=�r�����<==�)#>�^�<Ɍ=�G>s�R=G��=��>j�Y>aX#>r�?��v�>u��e�:�c���M.?�g|>V�y;�ľ�Y?�aY>kR����̿���4�?A��?�b�?đ?�Dn��>�Y��@E�odq=�e����I>���=6�G�Z��>0g�=��;���S�&����?�
@��F?ߥ���̿��=��C>��>!�T���/�F�`�ضE��U1���'?��5���ξ�Qh>�L�=t�Ҿ����f<!�>8^=�0��O�J�=K畽���"��=Mŕ>�MD>n�=|��ˮ:=,��=<>)�9>�����E����%=���=�nB>#Y>b�>�$?C�/?BRd?���>��o�'�ξ9����ċ>w�=!d�>���=�?>���>��6?^�C?)�K?)H�>�؎=��>R�>�7,�L�m���例��c�<|�?Sx�?���>�I<o�>�+4��>���Ľ��?�2?:�?�a�>�l	�M �PC�$�Y��M���>�R��Yj����|%=8�>R�'���<>H(�>8G�>�>1�0����=�>¡�>�g5>��<�o�>�;��|$Q�J��X�=�!n=�;������h)��2�9��%�=!�<~�
��>�n�<R!�=��?Y�>���>JF>>I ���O>�Z¾��T�=i> 흾�X���Q�!as�d���~�e�+>g�>1q��␿�@?z�>��5>5��??�k?�">#����蓮���ݽǭv��u�=�̱=�ꈾ��8�&c��O�q�Ӿb\�>�*�>䳑>�̀>��/�v�:��*�=ZTξ��6�؅�>��R����۽8�q�d*��(���y&b�w3�^�N?hF��j>@Vx?�N? �?+�>y^׽��о��	>R>L�A�=��l�Z��Eҽ�B?�F"?�h�>Q�a�7��O����T���>���rD�����ѱ+�5n�����(P�>J���L��M�;��ꊿ�Z��N�?�S����>��T?]Ҫ?*Y���Uv�L�V�U��/���>��O?f��>�?���>35H<K���7|���q�=%wq?�/�?l��?Fx�=�z�=^���z�>�2	?]Ė?���?xs?��?�BA�>N��;�!>�ҙ��z�=U�>b��=�8�=�]?��
?3�
?�����	����Y�L�]����<�-�=��>�T�>#^r>���=�sh=߫�=�$\>ⓞ>�ɏ>��d>�Σ>�6�>L����}���-#?I�=��?_�9?��]>`���e+����=� <�紾Z���"�;���v)�=)�s<�X�=� ��.:�>A�˿Z1�?�g�=+�g?��/�����[��>=9>r{��#?��Ls>9l�>)y�>�l>�8�>{>YԾ�>hm�r �k�F�p�V��Ҿ�>ZԘ�n7$��������:�
H�����/j�v3��e7?��as<�?����5�o���*����b�?�`�>jb9?U]��&K���	>l�>��>�����?��L���p]ܾ5�?��?�,t>S�>�Ww?E&?W�m=U�n�x���珿�H��7j��~b�~Q��򉐿+��B��=�0�?Nin?���? {b��B>��v?H�����[�>�E���y�C��=%�=4G��d��#��@L��Y��]0>�@�?�=p?�~?�Mɾ�����lH>/�??1�9?��z?(,?U�2?���
.?�=>gL?_	?��5?�	-?�?�&3>��>��p<1�<�@���G���M �Tɽ@�>��&�=��c=}��T'���=c�D=�^��?ů�,?<���˙<��u=n��=Q��=�>W�h?=r+?A��>si?Ʋ������JǾΕ�>ۃ��8����3�ብ�_�����M>�x�?O�?[w�?�Vǽ��-�^���:>��>���Z�]>5�>�"}=��-��[x=VX�=ׇ>��6����C��"'��S-�(7%���y>���> ��>��<��6>YC��BO����>ȍ�������\�:0j�ڤ'����<�>�N�?W?@��=PP;�;���֨~���n?4f�>PfI?��?ہ�:����N��?|�K�]z�>K�ƾ�	�,����Ԯ��Ȁ�K?.>��H�$��X�h>G��' 㾜�����M�
?ϾW=yK�R��=�&��ľ��r�܌�=_��=]῾�g�����P����N?&�}=����Xqu�.Ǧ��^K>�>��>�սV=\��t9�G��C�=�R�>�QT>����5�&�N�M���	�>�nE?��_?i�?L��r�5C�D���h��k�̼1�?+��>��?*�@>��=i���<����d��'G��*�>��>�o�#H���������$����>"?V� >ϧ?�R?��
?5i`?D�)?ZE?�u�>A���R��A@&?���?d�=��Խ��T�9��!F�8��>��)?\�B�F��>�?f�?f�&?ȊQ?�?�>�� �yA@�9��>CW�>D�W�za��& `>2�J?'��>QAY?�Ӄ?��=>@�5��䢾�쩽�7�=�>��2?Y5#?��?���>x��>G�����=ɞ�>�c?�0�? �o?��=>�?�:2>U��>'��=���>a��>�?QXO?<�s?��J?��>N��<�7���8��$Ds�?�O�6ǂ;6uH<��y=��3t��J�`��<s�;�g��JI�������D�S������;X��>�&�>�?`��m>񜻾+�F���>ٝ�<�O�~�����)��5>Ꭷ>�?=�>c�g�t;�=i�>���>Mo6�^�^?θ�>!��>El<��^�&A�퇛���>]�?۟{=J���E��܃���3q>�Ln?4�z?����D�:qb?�%V?-�Ӿ� <����<���H˾�\?�?�2�ߟ�>���?�rq?S��>�
}�{)t�����"]��;�A&=�I�>ܱ���W�yW�>�/?���>�;>J��=��龿�y����V?�G�?s7�?Kp�?3�>vB~��wۿ���J&��n^?m<�>�	����"?w���9о���ѫ��I�Ku������r���襾k[$�E����Xѽ-��="�?��r?�fq?<�_?���d��|^�<��"�U�6���E�fGF�XKE�$�C�kn�bg��^��b��,;M=c�{�=A�kݵ?��&?��'�Te�>�e��bK��Ͼ�X<>N����B�=o\x��G=�Z=^f���#������?�7�>)��>'�<?;^�Z]>�?�2���7�KG��V�3>�s�>7��>5��>
�]��(�zҽ�:þN�|�\�ǽ��u>��c?��K?��n?���&1�����!���-�e���[C>E�
>	��>��W����1(&��S>���r�a��񌐾��	��E=��2?7a�>_Ɯ>4.�?.�?�h	�``��A�w���1��d�<�=�>�h?��>���>~hνt� �U��> �h?���>A��>5^���="��t��Zu�V��>g��>w3?�>v���X�:̎�����;9�)C�=}h?ш�[R�w1�>�DL?/:��Mi<���>?��I�!� ���M}7���>�o?0�=R�K>i�ƾ����1����P)?�J?E钾��*�H3~>�%"?��>@.�>�0�?,�>Hqþc�D�	�?5�^?-BJ?TA?�I�>ݵ=����;Ƚb�&�.�,=Ո�>��Z>b"m=��=?���r\��w�u�D=�t�=�μ�P���<�����J<i��<1�3>��ҿL�R����Eh���2���
���Ѽ{Z���f<�s���T����i��Ԣ�f&��Cj��UV��?v����o��?��?�����A��g��kv���]v�㓰>�_۽�U��$��sν.�����Vc��+��m�5�
#c���+��".?G#;
t���賿��Ǿlhp?^�?r��?$D�,�M�E�3��_>M�Y�u��=�O�C,�M�������G?��>v��w9a�Y�)?�݇>�eż+�>���U>�����d�>�?�e?�q|�C0�� @��]@i� ��?b�@��F?ݤ.���־��>�a�>"~?_w>�{h�&N�H�ƾz��>�v�?/�?<+7>�F�/ ��R?�*\=�K�uz��%>ƤM>��c=��.�M2G>,��>/�ֽ��_�He���>#/�>������T��ݭ:Q\B>:���/�G�;Մ?W{\�Wf��/�ET���Z>��T?b)�>KC�=!�,?c6H�Q}Ͽl�\�J+a?.1�?��?��(?�ڿ��֚>D�ܾ/�M?�C6?K��>d&���t����=rU��F��^��'V���=j��>��>�,�Y��^�O��L�����={�� ǿB%��E�(�<V�|��|,����ʭu�A���˛���Z�5rؽV�=W��==?U>�\�>u�M>�TY>�Y?��j?�d�>C>Vx�&���?<����k���g�[�6k�����.ͥ��T�"V���ͬ���׼��W3��ֳ=�TX��*�����m�|�F޾�c?g��>"_s���i���=���ʨ��R��֛��A1ľzpJ�o�6��A�?B�M?0f���Y�E��hS=m��~�Q?����'BӾ[A����=+�u=��;�A�>�?ۺ="۾*�b�d�^�MO0?k+?ڂ��ݖ���(>�p��H=�,?@?�/v<㧫>?,%?(*���r�X>"�/>qƢ>��>�>�:���X׽FQ?��S?6����ߵ�>���Fz��<`=+>��5�
g���nY>�5�<ڛ���<��㒽ܱ�<ϲ_?���>I��G���t�ܗC����=��?��?���>B�m?��O?�%�=�	�![U��L���<)rR?��V?��=IS�� ����Ͼ�T.?kX?�>�l�mn��B�ܬ��d'?+؀?(�:?
뫽h��C:��V&���D?�\u?�[�s������N�W�>��> �>�t9�y��>8�;?֧'�ؚ��=ÿ�D'����?�@ى�?y �:�&�(Q+<���>�0�>���:��^��������<�?��x�k�CM�T��F:?4��?��?������=�ٕ��Z�?��?x���;Cg<U���l��n���~�<�Ϋ=Y��F"�����7���ƾ��
����⿼���>AZ@�U�n*�>�C8�R6�TϿ$���[оmSq���?J��>G�Ƚ����F�j��Pu�b�G�2�H�ĥ��rc�>�]>5���H���䆿U6�WH�<B�>f8�w�>�8�x���琾��;��>�!�>��p>��(�d\��.ߚ?k2���ſ<G��'�޾i�j?g�?ǡ�?o�?5SC=�v�<���a
�LRE?uO{?{�U?DP�b;|�˖�W�\?���e�r�����K=�]��>J~B?]�?�5��{�=�=�4?#5>�
����3�����F�?�c�?UI��?��?[�E?��!���tPƾ�}��Z>�%?�>���$��;�C�V��D�>46?�'��q��� e?w$d�k����_�L����>��)��Bq��4�=~Ὧ�D������,��ib�?�@�T�?���v��X��>t��>��������.�=6ϙ>vO�>�.Q>G��Ȋ�>];���R�O�>��?� @L�?NO��2��~y�=��Z?�'�>#��?�/�>�;>��V=4���	��= C�>��#>�:�;?F??Ŗ�>U.=Je�p-��C�.�j�w ���]����>��/?ܴ]?�T>�*׽|�;�oKQ�R��%�I�9;�=Ȯ̾ Tν*x&�mN>�L�>$>/�.��| ���?Ap�+�ؿ�i��/o'��54?4��>��?)��˳t�����;_?fz�>�6��+���%���C�?��?�G�?�?��׾%S̼>��>�I�> ս����ԁ����7>�B?���D��H�o�?�>���?�@�ծ?ci�� ?�S��g�g��a��x�T���,�=��0?����kf>y
�>@鬽0���ո��0�N��>P��?)�?hK�>�=m?�݇�Tv6���g`�>��{?,�>�����*�٭�>X��>�4�L8��f��M�U?��	@UT@�>J?5�����ݿ�������g��y��=-K��4D��Sҽz� >c�=	�)�	�S����=~��>>O+>L6R>�z">�J�=�_>������!鏿����>�*���I:��k����(��uy����X��3����z���սw<���M-�t��P&����=R�X?�R?�p? ?�j����>2�����*=ct#����=Gwz>y�0?��G?7$'?��=��M)c�[��᪾M����z�>�DK>��>���>��>F$8�'�G>ơ3>w�>��=$y =bi�;tB�<�nJ>�ŧ>,O�>�}�>@��>k�+�Ť�[�޿j����S>���=��?�r��[��ȕ�uh��ž$�O>��A?ۻ�=^R��7 𿇒���K?�����_�˾�e�>:�k?k�>�9>%޾v�=Mf�>�
�d��1�W>S�Ƚl-��� �6�>>Lw�>��g>��r>,�3�5�9�*�P�sF��k9{>�6?�з���4��mu�wH�޾��N>~޾>�aM��_��O�����
h�s7w=�:?�?�������v��B���=R>޾[>�r!=�߫="M>wjc��p̽�jG��O+=se�=�a>�??o�9>��Y<�)�>���u(e��3�>��d>%�=J�D?G%?vm�.�ֽ�젾8^J���+>N��>�UO>��;>�9F����=vj�>��P>7!w�����9��$�i�R>��E��-���j�K =i:���
>6i=>�����"�|o]<�n�?0*����u�R����|<p_P?-�?���:�=��*�ȑ�������?��@1�?��ɾ��G��?hJ?6KX����=��!?��>TҞ�~H���D$?h8��n�ȝ!�Z�w���??���=�O�������W=�_/?�Tɾ���>����훿�t��%w�~���X�>��[?�[	�x�=J���9%?-7�>[� �֣�5cǿ�Z]�_��>S�?��?e�n��h����E�ް?�P�?	�s?���=��ƾ��(6�=��H?6Y?n]?V_'��9T���>��?#�?[�4>�O�?Z|?��>p�N�'������΄��W|=�L�v��>l��=`�̾~�H��y��l���7�a�{+��� >��==�%�>��9�[���?�=|B��������U�>�>��5>��>��>���>���>���<1�x��H��}�n�K?���?����2n�'M�<���=y�^��&?oI4?�g[�0�Ͼ�ը>̺\?L?�[?�c�>D��Y>��-迿�~��d��<]�K>�4�>vH�>M%���EK>W�Ծ�4D�@p�>З>����?ھ!-���N���B�>�e!?��>�Ϯ=�O?]O!?u�?>�ݵ>O�F��l����B�A�>#�>5�?�(|?z�?S����P;��ڐ�0����S���3>z?x?���>�=��D��W���z>_����?��^?q/ֽ�k?��?��;?Z�;?�R>N4��Y̾i�H��p�>Vu"?����B��2����H\?_�?���>����D��7�	�F������W?jZ?��!?١��oh��ʾ�|	=:n���yຼ�<D����)>��>fJ\����=�`>H#�=iRd��B.�kO<��=���>��=A��_�{�#?�b=�rT���D>��e��qM���">̓.>�¾6D?��V��L��ޣ�������#��Ǎ?�2�?�Ռ?���v7c��N9?�Q�?�%0?N�>���B�����߾��@����>E��/�=uQ�>Z엽��ł��T\��j6���T,���?&?���>��!?M?XuG>ߵB>��Ҿ����;����ѡj�����B��\*�������s;%�&^5��Q��������>���G��>H^?ƬX>��}>�b>��v��=�>�?�>�>L�>Zw�=�1P<�K��E����P���X? `Ѿh���쁾g���=�C?�D{?�%�>N�����%��y^[?-�?@��?B�s>f3U�E�-��??��>����l@)?��8>�ڽ:�ݽ"��4�(�L�<
\z=�ݞ>���nf<��qf�~�j��&?�B?��=��ȾA <(۟�h��=��?��)?��(�ܡP���p�oV��R�C�"��h��A���w%��p�X�����h����(�x3=�8*?K��?F~ �ui�A��&�i�w�>�=Ph>:�>�ɗ>���>�J>k&	��v0��@]��%��怾Ok�>�{?�f�>W�I?�<?�{P?�nL?��>�M�>�&��#��>���;�4�>f��>��9?n�-?�&0?k?�j+?Tc>���I���Àؾ��?�?$Q?�,?�?�	��c`ý:2���k���y�jD���Z�=���<��׽j[u��5U=gRT>��$?�ח���t��Sξ�,�>AH%?L�?YB<>�(�#�>�-J;+3(?��?�c>x e��ێ���V�h��>�ϱ?OB鼃�_=�y:>XoT>׆�Y����\= V1��rS>��D������e>E�=�=N:�=ލh;� M<4,0=�8
?Ԁ?���> �>�������R
�d�>vx�>L�>c~|>�[�|Í��I���.X��R�>� �?c3�?���<j"�>�%=KsӾOվn�������c>��? }/?[�]?p��?�'O?(�7?�|>���5����w������$?� ,?҈�>����ʾ���3�j�?a\?=a�Ӯ�n9)���¾& սڪ>�\/��/~����5D��������j��z��?}��?�.A�o�6�({�� W����C?�%�>uV�>$�>��)��g�w$��8;>���>'	R?g�>�O?:E{?֪[?vT>��8�61���ә��o+���!>0@?
��?��?�	y?�]�>E�>F�)�Z�b������'��ނ�7�V=GZ>ʆ�>��>C�>D�=�ǽ1T��?�2�=(lb>��>ǣ�>���>�w>D �<pG?�>Pܻ�3�Y����X��f|s�1�t?ʏ?�8'?��<��F�Ka����>��?�?�?�C*?2S���=j/׼Έ����h����>���>��>�r�=/7=�z&>	�>�+�>sC�A��9���Q�1�?��D?���=R"ƿ/2r�7qr��`����H<b���+.f��ڗ���Y����=�o��;��������[����������<��PL���rx����>{�=�i�=v��=,��<=�ż�?�<�DM=�Y�<�=It���N�<2`:�ֻ̀�����5%�[�e<#1P=4:��".޾�ז?3�v?�eO?�??N�q�NV�;;�}R:?������?�#�.��=����ؘ5�J�X��)o�b��(m���i����E>�jϼFO>��H>��<JNX�dI>�� ��3>��R=�jǻ�e�=��t=�c�=�Q�=m>wg>E�v?̴{�)���!6�T@�&O??��>#N�=5���a{V?��>�V��Lÿ7�"�4�?�@��?��?�%��Dǰ>�����0����=�3	;$2�>�=�.��J�?�|T=m;�ͫ�����=�|�?=1 @@07?����)ϿûM=G�8>r�>gS�+�/�j�c���d���\���"?K�;������>�%�=jm��]˾�Z=�(>=/c=8!���W���=K���J)=�D=	�>o�=>�n�=�Q��f�=�P=*>�=��S>=�/�)9�#�>��"=B:�=��j>��'>j�>r?��2?Q�^?��>-�v��[�ĵ����>��b=���>��6=h�1>̴�>f=?��H?�N?p��>�Yj=Q�>��>��*��Tk�1�ྠ����8�;���?���?AC�>=jf<c ;��c�ƫ>��ˢ���?+r1?c�?lĜ>Y"��Y׿��m�.4��`>��������J�����LW���`�(��=y�Y>�-�>�,�>Ҙ�>k�>b'=���>��F=��@�z3�=>t�]��=��m>�)�=� >H��=��9u�=F=ɸ�<�����2=�� ��"�<��=`�=L?� >�n?81�=����^m=����&M9��m4<K���%=Z��8b�µ���Z"��	���s>��I> k�}b����?�c>��=>�!�?u�e?���=����ξ@ɑ�H����A����=�A�<F����S���v�&�Q��_��>J�>�Q�>n�m>',���>�2{=HBྂI5��q�>ጋ��'�7d�?q����m蟿��h��=���D?	�����=G�}?��I?�`�?��>�"��?�׾��0>�Ԁ��_=t��z�r����k+?��&?�i�>jq��D�<9���|O=��?������5�x臿yU��շ=�ݤ���>*��L����M�Yo��+�����"��u� �>�?y��?�,���i�a�T�����.}�Y3?�P{?Cx ?�<;?K�?�;���Z�$\���u2>I��?���?Û�?hH�>n��=5��;�>r+	?<��?���?��s?|?��y�>�m�;P� >὘�}J�=�>A��=�&�=�r?w�
?i�
?�h����	�M����^����<͡=���>m�>t�r>S��=��g=Rv�=_.\>�ٞ>�>�d>�>P�>I=��)yϾC,?n:�=�W? �:?eY>�I�[ߓ���-�W���u���.��W��=bu��0���  ɽ��=Z����>�Vӿ���?0��=g��V�?����=��=)�_>H"Q�:��>�	�����>���>�.�>��]>�2�>I@)>�Ҿ��>F7��\!�/OC���Q�\Ѿ�q}>t����!��	�"󽯧J��#���l�]j�W���TL=��x�<o�?�` �rrk�N�)��&���7?�g�>u	6?s���̈����>�C�>�L�>6��Ns�����K9�+�?<��?زv>A��>�?~?�2?h�f���I���0����MA��b����k�fg��Cq��f���'�>�~?۴�?�Pq?Wp
��v0>�l?\6"�gI����=l>��e�UT%>���>���ZӾ����Xa��Q��+�>�0�?u~�?Mk�>JZҼ�Y����=>�r=?[�3?�t?u�0?A8?A6��8*?�}>�?��?W�2?7�)?��?ۿ->��=���K�<�����1��P˽YIʽm8�L�=�Y=m�ӻ~[;d$'=Vf)=�R��	LؼѭA;�����<�=Yf�=[ �=ʞ>f:Z?�?j'Y>z�+?!韾�4���wV� �?3��q־.oӾ�־�R��L�>vϔ??`�?�K?���=c�'�"���&�ʼ��>���<���=�?��;|�O�{��>b�k>���=������5�W���?ㅾM�h�yR0=���>�|�>gnc�l�A>����<L�=*>ђ��e���o�gN���7��4�Ғ�>�hE?n�?b.>Y���ƴ�+q���C?�0?~�B?�΁?]E;k���`�>���B��� ����>�P�h�������ţ���6��%��c>mמ��렾�Lb>}���a޾ �n��	J�a��[�L=|�_jV=����վ�6����=a#
>������ ����Ԫ��3J?��j=�z��fU�o~��w�>���>�ڮ>�y:���v���@�����X:�=˲�>�:>������3|G�v1��>�GG?b?=��?��JMp��MJ��'��%��0��j?PN�>��?�
;>P��=o���Y���kg�BgC�-��>���>|��K<F�X����.��0R"�	�>�$	?[E5>�s?��V?n�?{�_?��'?�?�c�>L��FT���#&?��?Cֆ=]�Խ�HS��B9��AF�tV�>�5)?�D��>T0?��?-�&?8�Q?!??�>� ��Q@���>��>�W��R���	`>z�J?�>;VY?��?��=>"`5�-����M��_Q�=�>��2?T#?$�?�>֪�>⯡���=���>�	c?�0�?�o?�w�=��?�52>���>]�=��>���>�
?�VO?��s?}�J?���>`��<{0���.��GEs��P���;�bH<��y=���B4t��:�!��<"��;̉���/��ˣ񼮥D����H/�;�#�>�>Ƽ����X>�P���E5�s`�= TG�]��[h��{��N>��>o?4��>�����X�=*ؿ>CwM>�D*�a�K?�>m ?�=�Y������>D�??3��<����\v��W|u�7�=�T?N?�+׽}�Q���Y?��T?x3���`��8�40!��c���A�?��;?�����%�>��?�<v?ά?2��{r��*���_��#��h�<Mɑ>:긾��F��@j>��8?�u(?�'=u��� ��x�Q�žD��>b?���?��?��=�<��cUݿ����{��߾^?��>�k���(#?x��A�о̆���T�����.�pW��oO���
��ע$��K��%׽�=�h?��p?$�s?B�^?0� �$�d���^�C��^ U�7�X��G�D��F�wB��Zn�x��������c�`=��}��n@�~��?3'?�w$�l��>�=��Y���̾�dF>�ۢ�kz�5��=�/���/;=xU=�we�C4.�^����?s��>I!�>�;?^[��T?��2���7�[�����/>�7�>�E�>`K�>+�x;�0���׽_�þ�`��	rý�u>�c?�=K?�o?_ ���0������!��Y4� ,���YB>!�	>���>�VW���H8&�=>���r����d~����	� ށ=~2?Fk�>$͜>�(�?J�?�j	�����$tx��E1���<���>l�h?�Z�>�f�>WѽH!�6B�>�q?Λ�>7��>�������"�~��Ƚ?K�>��>�� ?�! >��;�^�]��)�������:���=�G]?�k���D���>�nG?�H< ��<S��>��Ľ���IX޾��Z�=2?y�=L>>���Q`�݉��򘈾�O)?L?�蒾�*��6~>)$"?�}�>�+�>�0�?g)�>mqþ�H�]�?��^?�AJ?GTA?J�>�=O��.AȽ��&�]�,=e��>��Z>�#m=9}�={��Jt\��t���D=�l�=�μjZ����<�����J<���<��3>�H׿S�<�g�ȾZ�������L�/���o�	�˽G�*��qվ�Hd���s�W������3�L����*�-�j��?	��?�'�|G���������-���w��>���5m >�D���k=�)B��Ǿ������]����V�+�	�m�'?����ǿH����;ܾR" ?�C ?�y?;��"�ΐ8�7� >�Q�<�3��J�뾜�����ο������^?��>��f9��%��>���>>�X>Eq>o��|Ꞿ��<r�?��-?J��>Őr�v�ɿ�����Ĥ<���?��@ZHH? {*��w����+>���>�?&�@>�Jƾ���!�ξ�ʰ>o*�?w �?�>��"�{����D?e���x������>A�>@�����g�,QE>C�>f���]�� �^��>V��>�Ch�$���o�¾»=>�	�>Y-����w�5Մ?*{\��f���/��T��U>��T?�*�>�:�=��,?V7H�`}Ͽ�\��*a?�0�?���?#�(?@ۿ��ؚ>��ܾ��M?^D6?���>�d&��t�ȅ�=�6ἰ���|���&V�s��=]��>��>��,�ߋ���O�!J��g��=��{�ƿF}$��]�� ==4V��{\�彆ծ�"�K����Q�n�����i=ԫ�={#Q>+��>aU>\Y>�W?F_k?��>9�>����n��xξdm�Q���.�����0�f������Q߾"z	�Z��|��l;ʾ.=���=_,R��i��>A!�$�b��.F���.?�%>� ʾ �M��1:<{Aʾ0���%������˾s�1���m�h��?�-B?����
W�	f��C������W?���<�] ��3��=��ώ=(��>�'�=x��^3�/�R��/?�?Df¾
Q��f�>.4
��7 =�w)?�� ?��<�h�>=f#?��0�����4V>L)0>z��>��>Y>�{����ѽ\o?վS?���Gҟ�d��>���zo|�]M�=H�>s3�i�p=R>���<Ng���껍���� �<&�Q?�H>��(��*����,f>�<&>2�8?�8�>!��>�b?�4G?7��<�^0��#W�%�Ѿ�7N>��R?�`t?��>c�����Ѿ�Bw�}s]?ZV�?D5�>�B��g��BTC��'�U*?�<s?	�Y?�<N��Qn�������ξ);=?A$d?TA��Ҕ�f�$�����>?cT�>��>�	��'z4>z�I?�mg<� ��6M��Յ:��ن?R��?'��?L}�=�:<�D��>ml?�K�>$�վ�-��e���=&3�>�}"?~k���m�Ⱥ
�w�����X?��q?\�?�,���a��8�=�a��bN�?x)�?7`��ؽc<����k��}��_��<dR�=�.���#�	�7��Ǿп
������2���a�>cL@wo�K��> 8���?Ͽ���Fоj�p�]�??�>��ƽr�����j�W�u���G��I�롌�7�>��>��VՑ�P�{��|;�������>���t�>�yS�N��򶟾�1&<�ڒ>���>���>ZY��Ǧ��ƙ?mi��Uο1����|��X?]_�?]�?In?�@<Θv�z�z�S��0G?&Ws?�Y?��'���]�5���d?-[��*i�7w9�/D���s>��&?�	�>W���67=�aA>���>Kx�=��=����mF��o�ľ�ƫ?���?ǣ��0?$��?��/?9��#@��������ű�<g�L?ګ!>b���	8�2;E�� B���?�1?Ds,����,d?��N���[��X���=���>}�ؽ:��Tl�>i�:ov6�Y	��������?]X@�	�?��^��G��S�>~r�>�L���ю��"p>/�?�O�>���<����oX>4��x�@�sA�<= �?��@J�?���A����Bn>@#u?��>�|�?٣>ݚ�>�n�=P�Ҿ�Z�=h�>{C>q")��?�?���>���=�P�=r
'�($c�Ǵ|�ʻ"���N�v��>%%O?h^?���>��hf_��a,��%���_��A<_�b�~+7���(��^�=O��=�^d>���<o�ܾ�*?V�8�TGؿ����� �d�H?��>Ф�>������4=q4t?W-?>��cA��:녿i�5�X?�?X��?Ĝ�>�]���=�`.>Z�>ճz>q�w�WLX�47N�^��=�!?U�8��ʄ�#�c�a�z>f��?��?[��?o]��
?����ㇿ�N{�#����&����=��1?�r�a<s>���>p��=��t���ZAs�X+�>y�?M.�?[��>:�f?�Jh�f8��M$=�s�>Bqf?��?���<���1�I>��?V���㍿!&���e?n�	@��@��Y?W��|Rӿ�����;��$����=�<5G>�򒻘]`�'#>d�R��C��$�=�̝>
w>{&�>�4>�=�]>�}�1��Q׏��5��d�;�E��+X�cl½W1%��սU�9�H��|�Ⱦ�󓽶u8�)���U���9W���{��b�=Iih?�=`?�`?7?�>����'=>��Ⱦ�=��?��� >XD>H0?�;8?��.?@;v���þ�_^�Q恿�W¾v�7�3ǯ>8�n>!k�>�;�>k�>�j�ʁe>WS>7e�>�2�=R�=�zS�T���<>ץ>�N?�3�>�C<>��>Eϴ��1��k�h��
w�X̽0�?s���M�J��1���9��զ���h�=Kb.?"|>���?пf����2H?)���y)��+���>��0?�cW?�>����T�-:>3����j�Q`>�+ �{l���)��%Q>vl?��f>z�v>��2��8�a�P�ڻ��Zy}>Bv6?�k���n:�� u���H�6�ܾ�M>�ƿ>H�J����8��X#��j���=�i:?	�?8����]��	yx��Ԟ�7�P>�]>�,=�3�=�]L>�g��ƽ�9H�o<3=���=��\>{P�>�
R>�Y�u>۾�C���A�>qf>V�$>�\K?%
$?��?�/+�_����;��dR>l�?K�>~OJ>#�'���p=�?GQ>�F=�zN��p&��Ǧ���O	>�s�=� O�h೼ٽ�=?����>>��d�R����G'=��|?JS���hu�B�(�>�tP?�f�>�M�<(�2>$j�诟�AI۾ 1�?/@ZV�?\$��V�;�>��S?6[��"�= E�>VF�>cW��������>���f������+���?,��?�R�����s|�j�>L�?z��?�>�8��i�����\���Z]="�%?޾-?/�о-�;=�K����!?d�>�߾�ϥ������f>���>��?��?�[���ܙ�9T��@?�4�?�X?gZ�=�� ��p���x�>$>?U!?�M�>8,<�vO;�U�?�I�?�Z? �>��?j�|?��?�\�# �����\����e�Fו�LT�>'������\�A�A����@���Lp�	5-���&>M�X=C��>p>==�=��ф�=&��^+ؾ�������>2Ŕ>ݾ�=�I�>A�>a �>�i�>�喽�����)��ɉJ��kD?�)�?�RԾU�u�Y0Ӽ�8i=\n���?a_2?ly޽.({�>��U?r?��g?k�y>g*�-5��跿��Ǿb��=?��>�n ?�L�>�����=y��_����>�>-��>��Խ�꾧���R]z=���>a?mf�>��(��W?��0?O��>��>�8�����+�X��;?��?��(?��?�@?���	���m�����okN���=��}?1�8?�g�=+�����F�}��2�>-��?<}�?�
�R	-?#�?%�W?��I?��X>��;�b�4B�=s��>��!?���A��M&�W�h~?�P?���>"6����ս�Aּ���~��F�? (\?�@&?2��1+a���¾%1�<��"� �T�z�;-�D���>@�>]���ꉴ==>ذ=�Pm��H6���f<Go�=���>��=�/7�����f&?φ<�!���_�=f2n��^?�	:@>��K>h9þ�lO?x3���x�����((��:W�H$�?���?9�?e&���e�2HE?=�?�2?���>�j���TϾپ%h�ȁ!��V����=���>����(m�Z������{��4�ĽB���?-T�>��/?�
?�x>�[>2�¾Mo0�I�о���qng�.�
��#��y�	��I�����ܽw��N���'��>���� �>p9	?�v>k>C�>Q�=�bY>��Z>/�`>�r>�i9>�0�=��K=L�2��[��dR?��e��\�Ͼ�����8E?_�]?+��>|��j��ʋ��<?���?���?�!o>ִT�/����>��>E����$?���{�j��D=�ƹ���G���k�lP���>��Ľ:�D�:�d�J�z�ħ�>jU?�L@;d樾5�ݼ�ɞ�+N�=��?�:?}/ �K��#��ЕM�b�W�����_<f�qf����%�%h�z`���Њ�æ���2���*=��.?A�~?�_������W���9m�H"8�x�>Q��>�s�>���>2̈>s��
p �)�R�,���:��(�>JՀ?b�>�EK?��6?�S?<L?T&�>�M�>I���u�>�M�;�M�>��>�[7?��-?o.?�f??)?>�c>���9����Ҿts?�?b6?��?`??ゾ9�н�8ݻ�̌������G���6%=v\�<����e����A=PM>S�<?h(߾e�r�M��* �>"�R?(��>`CC����t4�c�=�&?;��>t=y�B��3O��C��6QH?���?�#��=�-n=�/�=ĕ`�����@��[꼵�k>ޠ�}�S������8���Q��A�=��=�}l=)�>���m��>��?�>���>	ۆ�IK ������=��8>H<>Z�>f��|���Z���{a�`>�>9
�?�o�?��[=���=:�>
a��|֤�-Y�7���I=J��>N�?x�V?�D�?��2?�#?銦=��wz���A��v1���?�,?���>����ʾRਿ>�3��?�v?�a���8)�.�¾>�Խ��>m/�H~����KD�������u���ƌ�?)��?��>���6����˼��Mz���C?`�>)�>���>��)�'�g�5��{;>��>`�Q?a�>V�O?�8{?6c[?a�U>��8�����A♿@�X�>;>)U??q�?Ɏ?k,y?���>x>w'�k~߾����-���0���N=}�Z>6G�>v�>JQ�>\P�=��ɽ����
�>�d
�=�Ta>(��>�d�>Ao�>�<w>��<dG?���>"���#�v���yV����H�_t?'��?�b+?ǜ=����@F������m�>��?I/�?9*?PP���=ԧ �To����o���>�Y�>�֚>��=��8=: >N��>���>����+��8���F��Q?RID?���=�� ���j���G	�����=l���f!7�{=�S�`?r�$��<+�]�ʾ/}���9����A����㬾�0�>\7>{��	�>
��:A=�'�=u��i6%>41�9x4=a���"�F�kς�a=��݊T=@1��e �/�?�4t?�)�>Gx/?�">��>ׄ>���>�ؾݢ[?������S>����Ϭ�n���
�ؾ���
Ĭ���t�z���F=�н�r1>��D>*a�<�t1�S/�7ͽ�D�=�,	<)����=���I{�=�O8>�?V�(̊>�*`?��N�>���M1�u���>��>�կ>�H<���W?���>�w���-����d�?��?7O�?sE�>^��ܳ>�(��#Q˽,�=/�=[D�>��=ޒ����>��\>:(�之��$�����?.�@�!?ě�}_ٿ��=��8>sc>
�R���0�%�e��i�w�Y��k ?L�9�clž���>�=Ͽ�bξ�'&=fB6>7|�=P�ODY��̟=J���CZ=�M[=i��>�"H>J��=5�����=�!`=��=�lR>������1��l,�D�K=��=�\>�]&>��>6{?-�6?I|P?��>í������Ծ	3c>l����{q>��Ǻ�
>��>ʺ<?K�d?p�O?��>5߂��֯>lf�>rS*��Tb��oؾ'�����0�7ˋ?�\�?A�>���7S0�G�!��
:�:o��4?߼)?K� ?��>j�A�޿k���w*�J����~���0�<�.����!�=eG��n��4�b=���>��>�ۏ>0�3>���=R>f��>(�=t��;1��=��<�%�<�;\�E0=�,��܃=��ļ�E}<�mԼvf�a��~�����;��93U�i��=b�?#0>a�
?���=�I��$U=����aL��W6=/8��g�U�_�h���{���*��8O�d6>*�+>̶��W��c?O�>�'<>�s�?C�d?7(>�Y��⿾�M���.Խ������K>��=i"���l�D.���b��$ξ���>��>k��>]�l>x,�z#?��w=N��\5�k�>�p�����9�^@q�n=����Vi��ĺ�D?�D�����=�"~?رI?�ݏ?t�>�&���yؾ�*0>�0��]�=*��$q������ ?'?���>� �)�D�vɾ�A��W��>L;%���L��K����7���;����i�>=G���ZӾʤ3�Ʉ�0���fKG��9l�/L�>qN?$&�?�Vi�%���R��L�i=��!?+q?:�>%)
?�c?�-<��-辸�p���=�n? �?��?"-&>k��= ���1�>Y)	?ﾖ?|��?@�s?4�?��t�>$�;� >:���A�=�>�l�=�$�=fr?�
?z�
?\k��\�	�p��q���^����<�ҡ=w��>�o�>�r>z��=w�g=k�=�&\>�ڞ>�>$�d>��>�H�>�č�z�˾"?O@>P�>�<?\p�=`J��[�8����=m�7��U�O'�]��5a���B�rlݼ���<�V\����>r�ǿp�?u����̾�B�>��0A�;�>�O>d���p��>�����>vrY>2�>�׍>��p>mS>�پ��5>�(�p������%p�2z���W>OI��=:* ��q�����=��Q�����]�*!h�ŕ?���3>��?=o�Oo��A7�~�D�
��>���>��I?o�����<��r>��>�~�>�r���쑿�q��RBľGuy?���?(�?>�>Gt{?	9?�#>Aq ��Ⴟ��RX�u�����`��@P���Z��~a��L�?Vg�?�%?q
N�j�S>i�[?���m�w��>��C���
T�=�B>��)�䴽���ԾR`�������>ʕ�?��_?
� ?l�"���q�`)>��:?<M1?�t?�1?H;?�u�%?a2>�?�&?&N5?'�.?��
?�21>��={���;�&=ð������qYҽʽS��2=�bw=i� �o@<8�=�˝<k�켊Bڼ�}!;Qգ��h�<`�<=���=
/�=���>�xQ? �?�a�>�e6?�n��J�b���q��>�IL�0Ѿ.ϴ��v�����m>R��?wX�?�H?�>6���	��W��.?��0��Т>?�>;�=?�u�o�`>��f>�*�=��� 5�d	����+��J�n��;E�`>fz�>C��>�r�wƇ>{q�tL�2��=%�nPɾf�_�)�=��5���R�}��>��??\z?���=	)¾�*Ľ+g�j�1?�d?e�[?Io?�g�=&R�H ��LE�w���>��\W�K|��±���	F�E|o�Q>�TY�c�J����>���P@;��l��gW���ɾ�K�=;����/�=2L���վ�����=D;>��Ҿ.������c��_S@?d�=�œ�n�0�"��zR�=u��>�͑>����Fq	��K�'V���)�=Փ�>7�0>K`a�����GdL��U�i��>�UV?�Ds?b�?��ὀ�u���d�J/�h�����<��6?@��>?�k>�2H�JNžQ)��ms���H�@�>�?�C��BV�c!���=����<�=�&>�"�>�>Y�?DCm?"y?�b?�s?&��>���>$� �r7�A�<?? �?F�>:��KGX��<0�)�@�X��>k?�^��L�>1 �>	u?}4!?�zT?+�?���CW׾�Z���>~��>"zp�����9%>83b?Uڦ>Q~??jw�?,<i>"J'��s����}R>�RT=�p5?̔7?�:�>4݁>l�i>�&ξ�G�='�N>h-V?�?n�c?s��>� �>~�����=OB�)�o>*�H?�.K?>�[?�=�?9C�>S��>W�H���q�=�/= �=��7>1[<��>�=h�ֽIՆ���;����uts:r�Y=���=�\佉S �X�>�[R����>R�s>����E.> �þ������>>�)������̃��j9����=�{>0��>T��>	'�ք�=�]�>O�>����q'?0?@�?b/&���c�9ؾ+C� ��>�HA?��=Ynk�I8��Vt�߸[=��k?�`?
[����b?H�]?�c�=���þ��b�����O?y�
?g�G���>��~?�q?p��>��e��6n�����Ab�R�j�hӶ=�p�>Z�_�d��=�>7�7? M�>��b>`<�=�o۾��w�e|���?u�?y �?1��?�3*>b�n�3࿦b�KH����<?JJ�>��ؾx5?h��<��Ͼ]�����`�vP��S��������^)�֬v���x�>�. ?bGd?xs?6Z?v᝾9*c�Fp�����pl_�������J�dN+�>r8��W\����b���᜾mm<��.��*\�C��?4;?L�%����>#7���������c>��<��P>�9{�=�s�%\ݽL�>�}r���'��Ķ��?Ok7>�ݲ>�Q?��@�/�@�vH�:U������>��t>�m�>~�>�"T=׶X�i�B��̾�{?��vb==�v>�Kc?L7L?�Eo?M����91���16!��I2�L���ۙE>��>U��>��Y�L!� %���<���r�eP����K
���=��1?�W�> ��>6�?�y?+��߱���gs��1�%��</��>~vg?�>5S�>������ٽ�>��l?^��>U�>�����X!�[�{��ʽ%"�>��>���>�o>I�,��#\�Uh������)9�Oj�=��h?�����`���>R?�.�:T�F<Fx�>�v�ɸ!�S����'�,�>gz?d��=��;>�}ž��{�:���n?�p ?��g�D��A�v>-�%?��?D˦>4�p?�E%>�^ʾ��	�u&?�eg?xN?J�S?Z��>Ѽ��j��!I��̈́����I>��G>�H�=���=U5��FL����5��=���=�7�}T���/���w<4�=P�=�/�=ݿ�YK�#پ5(��뾾��Q��ѵ������޽� ���ș��Mz�%�%���J��Z���y��H��y*k����?�s�?;�����!e����pX�����>������:ң��tὤ�����Ǿ�s�����M�L�;Dh�qh���'?���5�ǿ����8:ܾ�! ?A ?�y?���"���8�?� >�C�<@��͛�ϙ��(�ο������^?���>��.��=��>���>j�X>oDq>.���枾^�<��?�-?���>}�r�s�ɿ=���V��<&��?��@vG??�;���ɾ��=ռ�>J?�1�>�u��������2�>�ş?���?�V'=�`�n��Y?�|�;�_B�r:���=�w�=���=M�ýc�>W�>C*D� ae��4��x�$>p׆>T�'�^����h���̼ �Q>�퇽��ɻ2Մ?*{\�f���/��T��U>��T?+�>D:�=��,?Z7H�_}Ͽ	�\��*a?�0�?���? �(?=ۿ��ؚ>��ܾ��M?]D6?���>�d&��t�΅�=�6�y���n���&V�o��=]��>k�>̂,�����O��I��]��=9���DY����4��4)�s�!��Sa��0�����k�v�>E�����g�������4�"�ռ-�=��g>m�>�G3>pr.?@?6�?<��=Tu>n���ֆ�MW�������3>eѿ�h:��A½�����e0ξ`g ��43����_������=V����.�1��n��?1��.??[�=�|7�C$P�u\=�>�O���K&�=��]��,��DO[�H��?[�?ָ���f|��,�F�q�R��ğ�?��5� ���ѽ�F>솦��[�=���>^o/>fኾ�E���C��98?m�?%<��6���qU	>����=��"?�z�>�ز=8��>ħ$?f�@��v'�Q�X>̿>���>�{�>�~>l���c��a�?��N?��벾��>P'����Y�
�=)Ό=��=��3��~�C>���;�����;�ö�����tW?Vq�>m�)����l:��.��3b<=T>x?�1?��>�~k?r�B?NC�<m���jS�^�
� Yu=T�W?zi?��	> ����Ͼ�ꦾFw5?]e?h�M>�Lh��>�{".�6_��?y5n?/�?�����}��������q6?Dw?�~]���������W��k�>sK�>��>#s9�ڤ�>�>? �(&��������3�%�?B�@J��?��N<C�tґ=4=?C��>��P�@yȾ�4������ s=w��>Q ��2Xv��I �Q�)��A8?�F�?�g ?�ƃ��� �7>�]��ے�?F��?޳���2�Y��������	>RN�>/�o�. �=�����_����{$�Z��W���ot>|� @%> =���>�ZF=�Zӿ����>�����������'?fW�=m�K>^v�����p�{�Q�Dh�񇣾��>u	#>s#��S&���y��p<�����>�S;>`I�
-���|��2o&<� �>��>�>p>�蕽����?_�?7��%:ο;\��i���X?Zx�?���?�k$?�N�<x�m��~��:N��-MF?�$m?l�W?�1ּb�j���W�q�j?�W���N`�1�4��CE�mU>Q3?�;�>��-��o}=�>`��>�T> */���Ŀ�ֶ�������?I��?�^����>�z�?}r+?�g�:���U��~�*�Đ&�<A?��1>�����!��-=��Ԓ�g�
?Ć0?����/�6�U?0�^�~�e�g�'��򆽴��>Q��l�5���*��x/���e�����/�k��ɰ?���?%&�?.���$��%?�"�>Jn���-��g�=ʹ�>�>��7>����[R�>�ַ?�>�?�?ƞ�?s?���$��7� >P�y?���>�?�?���=�?Hl=����  �=�	>�2>�������>�C?_
�>�R�=Vx7�/y$��k:��p����FuK���x>ubx?w\?��>���z\��.���:��vb���=��"��4&=A�ܽ��=��~>�
>�3E�qWؾn[i>��#��ܿ�+��VH�D�.?"��>�'	?x�?$뾑τ��t[?HS�=�2�OH���A��ҕ1����?��?���>O"�����<�v>O�>SzK�����������>�
3?,�@�)����z��E��>i��?:��?Dw�?�SI��,?�,�u�����}��s�,7�#3�=�c7?n��v>���>c�=C[v��쪿4?s���>}�?�\�?�V�>*�k?Mtn�s�A���6=���>�Ni?x�	?����u�lI>�?=i�އ��;��v�f?�@"�@]?Ω������Ճ�[о�7���@r</>�t�>m=��&�*>���@G=�5~�j��=W�O>��=ĺ9<E�O>\��>��;>�,��\Q�v�¿���N�p�!tǾ�*߾ÖM=�y��P$��}YA���\��9Ծʊ-�E�i���޾�gC�P��<Hq�<��=p�T?tlR?$Zo?�� ?�x��*>|����4�<��,�)��=��x>"�2?�|I?�%?���=���X�d�s�t���m���y�>�[=>6h�>��>��>�8�;0O>V�>>��>��=��5=�<���u�<MwP>��>�'�>�>MC<>{�>2ϴ��1��W�h��
w��̽"�?����@�J��1��x9��Ŧ��i�=Qb.?�|>����>пP����2H?5���v)�&�+�5�>o�0?wcW?&�>���T��:>տ��j��_>F+ �0l���)�&Q>yl?Z��>o�>�1�����X����;�>�?FB��ȣ�T��3G���V�%>��>�/��ؾȚ�ܷ���v���<>$6?��)?����*�̾N���̹�o	(>����n��=ET�=�$�>���=�!�����<Խ9�#�>��==15?�9R>4� �J>�;��8�+�S*Q>��>�6�=xIn?��?�;M>��;�ԛ���+�� ��=�$�>P�>�'�>r�~=�7>cٍ>T�>�Խ��¾����8���Yw> ��=� ��Vƽ��~��Z8��}�;�P8�J%=`DY�����~?5|��b߈��뾲C���kD?�,?D!�=/aF<��"�+���S��$�?m�@�n�?�~	�ҢV���?�?�?\蝽���=Tw�>�ӫ>
ξܚL���?7!ƽp���6�	��2#��N�?�
�?h0��ɋ��l�:7>5[%?��Ӿ�>�>K��0]�����R�u��e$=i��>�<H?k;����P�2>��u
?:?�b򾳩��� ɿ�sv����>��?9�?��m��C��@�IY�>���?dY?koi>N۾nuZ�!q�>̼@?��Q?2�>�9� �'���?Eڶ?q��?\>k��?8�z?
�>�ûM�2�%S��l��U�=:y�<i��>�/ >�M��{�8��Q���\��,=o��+ �D_4>RZ\=W�>	,�f�о�T�="Ҭ�Y����q�����>6Bg>Tn<>��>R?�(�>ME�>�=%@�%nq�	x��G�K?��?����*n���<F��=B�^�	$?�G4?w\��Ͼ�Ǩ>[�\?j��?�[?�d�>���U?���忿|�����<��K>�4�>yA�>P0���<K>��Ծ�?D��c�>�ݗ>�n��4ھ�.�������K�>�c!?���>���=� ?��#?p�j> �>\RE��/����E�	��>`��>|O?��~?��?�ù��Y3�8��ס��[��vN>Hy?�V?�ߕ>�����~��E�I���I�������?Q�g?V�余�?a�?�a??��A?��e>�����׾CN��PԀ>S��>tV�#����A����.��~"?n?�\�>7�������j��+�Nhc��
B?s��?�`>?PB��(xj���� o�=�t���LD��2��6��ٯ`=�=�=��ýӷ=���=��~���q�5=	]@�p��>�e>��ӽ��{M-?	��C��h�=�r�k�E�n�>e@M>�m���Y_?X@���z������:���fR�>�?��?0h�?�����g���<?^y�?��?��>�対��۾$Dྨ�r��|�7�� #�=���>����
�h;��YM���N��2�ؽVt�̫�>���>�?κ?��N>���>����e[�>��7���g���߶:�PC8�����Y���:�a�0�t�Ͼyw��d�>�p�Q�>t�H?��i>�!�>�?�>WR6=��>�l>�jq>�g>�H>�G>�>J>ǁX��7R?c���d�'����󢰾Q9B?�td?�1�>�i�3���1���s?���?�g�?�Bv>6wh��+�[?�>�>���`
?��9=ψ�ɱ�<�:��î����6��׬�>��׽�:��M�}4f��z
?�F?:���`�̾F�׽[G��X�n=�@�?��(?��)�.�Q�H�o�N�W�{S��y� �g� ��*�$��p�~܏��T��� ��>�(�R%,=��*?��?�y��d�^���*k��?�d�f>O �>�J�>�x�>G�I>g�	���1��^�_'������?�>}I{?&՗>�AH?T'E?�
[?�$U?�Gq>,n�>�m���`?�׼��>�=�>Ng8?[�$?c�5?�~?�u1?���>y�ƽ`d��H$����?d?Ml?7��>V�?yI���}�g;6<`5!�����-��k��;��G=�#��]�<s�=<�t>9�;>�zJ�|�*����'>�o3?�̡>��>���&۾n�>��>�n?�R=��ɾY0j�k(�A��>Wć?�<x	>Bz>��>:ܡ��n�=k��>�V#=���=-���[�=ա_�e�>��z<�sӻ@�ѽ�M�=��ڽJ��Wy�>7�?���>�?�>�?��ե �����\�=�Y>�-S>� >�:پ�{��$��H�g�/[y>�u�?�x�?��f=55�=Q��=Lz��mM�����x���5��<�?rH#?�YT? ��?5�=?mb#?��>-+�8M��\��$���?@�1?�l�>���#0��hc���iD��?�F�>�MT��h��)��i���j˽+�>��)�߃v��C��QDT�Dnt��1�%���"P�?�y�?����m�7����픿�齾��2?WU�>(y�>x@?D1"�Eg�n	�p�+>d�>��E?N� ?rˊ?��?��q?�?�>��̿�SƿLc��C>J�w?��?�%�?37�?�@�����<�>;R�վ�YI�b[<��w$��v�k��]�P>U��>���>��>@��=�m�-�8�����c�=�9q>m�?,�>Ԋ>7��>I��=�}R?_�?/-��i��������½s�伙�S?Xn�?e?���=_Q���-�y����;�>N�?O�?�w?+����=e����ͭ���5����>ç�>��>��w�)�ν$-�=���>ˁ�>�z�9��N2�'.Q��;?/�e?FO�=�>���g��l�	�d�����������\�a>�F����>�+����N���G�s�������c��h�F�=k�]�l��>��L={��=4��=�F->���=�F=Z�O�e]߽�=�W�vy=}�=t��=��>�q.����<�tM��E�=�A˾=;}?�*I?z+?��C?Y{>B�>�"0��d�>�S��$p?�U>��I��ϼ��}<��ۨ�
���<NؾNb׾S�c��<��,�>��I�%5>�d4>�E�=���<��=��s=܎=�z��S=��=F(�=��=���=�>�6>�6w?P�������4Q��Z罔�:?�8�>~{�=��ƾu@?o�>>�2������{b��-?|��?�T�?5�?Ati��d�>@���㎽�q�=m����=2>���=k�2�W��>��J>���K��p����4�?��@��??�ዿ͢Ͽ�`/>+����&��[�{2`��y2�� q�����-?��T���m<�sG<��>�3�ݕ��Wy�ӌ&>�د=m��=��,�s��=�mc�	��<<=�=��q>�?i>7�q=?����e=�彈@�>D۳=���=�'ͻ탠�W|.��ѽ�i\>��>�?B�#?�Q? jm?�?�#s�뻬�^���o�>�=���>��=�W�>���>6�U?�V9?��>3��>r�p>m��>�
�>\�B�׎���(��o���Q�<�U�?���?ޭ�>Ԙ<��A�-U2��V��ƽ=2?F	�>�U�>3�"?"��f��&�~�.�������F�&=��p��Z���RT���]�=m��>��>�k�>�w>6;>*P>��>��>!�<N�=�ā��t�<λ���f�=�z��$Q�<6�����=���9��#��t��)��;-�l;<G<��<jZ�=��>d>��>��=;7���:/>����ȩL�i�=y䦾�@B���c�=?~��/�,�5�#"C>,yW>�;���0����?�Z>�?>g��?��u?&$ >�f��,վ�)��\~d��T��{�=�>Qa=�<b;�| `�G^M�<:ҾU��>�&�>&ۢ>��w>|�,���B�Y�w=[��?{0��5�>�N��D=<�#4�Msp�aӣ�����wvc��uF���;?�������=�g�?��G?�2�?>��>{C��'P־K�'>��q���[=�C�^�\��ɸ���?�;'?ۉ�>\�ھ�B�U�ھ��ڽ߀�>��X��]T��G���M+���;u���vv�>�����BȾ�H3��م�P+��.-H�h�p��/�>��L?qd�?+ h�)聿��O�V���G����?��f?B��>�7?�H?|$������!���4#�=b�j?��?��?�L	>랶=�Z�Y��>�?珋?�ۍ?�h?�m�־�>Q��8X>3C.��VJ>��>�u�=��1>��?��>�^�>���ϻ���K��e>���=�4>��>kۃ>d9�=��0>�/Q��g>t�>���>�Ժ=߆�>�
�>+܀�
���j$?��E>�~>±C?�m�>y@:k��;m"L��M�=�&�\K�/�
�t;,��7>�2=�Jq������>ӇʿO$m?�H>E(��f�>�荾�眾��>���>O��z?��<k��>�ѥ>�y�>��<�V>h�>�x ����=e1��&�A�Q�~4�:˰���>u\e����f��Sƽ�N�j��r��3����_t����Fk=?Qh?�6�F~��A.�9�y��)?�[�>ȝ5?OH�g��E%=P6?I"V>�1��u���A���˾q�?^W�?�=c>��>��W?��?n�1�f3�WuZ�O�u��'A��e�̻`�����͜��"�
�K��Z�_?4�x?�xA?�[�<�:z>��?��%��ҏ��(�>D/�G&;�WG<=$+�>�)��]�`���Ӿ7�þ�7��GF>�o?`%�?�X?_WV�gp�-b#>�8?d�.?�[s?�>2?xR=?N����!?�#>�?��?{4?�0?��?��=>�g>1����f=͘��	E��(kӽ��ͽF;��r�9=�X�=� :�n;:=���<(g��),Ѽ��\�s���w�<��)=�P�=u��=O�>}M_?�f�>קּ>\6?!���d6��孾�4?�A=d��x�������L��4>m?]O�?�xX?&"m>�C�ǚG�e<>�Ɖ>��>�h_>L�>����S�H�j=c>�>���=�FF�`͂��������|3=m�> y ?�ɚ>hf=��>pӛ�V&ݾ��E>�9P�>�/ԁ�Z-�]�+����x��>��&?�?�O�=�������'mk�Y@?7_?fB?��?BC�>I{���3!�y�:�x7#���>��ʽ����4������A��+u�=���>)���{�/�>Ň>�� �Dzо�{e��T��M[��w�=��<> =3��H��5����l=�Ӡ>	�Ծ�Aξ�ē��㥿k>?ў�b����P!�뷾M�=%�>-�>{��:F�^II��a��c�;=�<�>��=�H�O|���V�rM�d�>j�K?]�m?*�?�I�H�v�Fv]�=�멬�2�;�ro?#�>m�?Nt>�?�=^⸾�\(���z�]�G� 4�>�?mu��m�A��7��Z�վ�>;��d�=�X?g��=���>��T?Q� ?"�z?S?>W�>2�^>�H&��+ξ2�)? f�?���= PѽM7W�r�9���@����><�-?��F�r��>B�?�??�0%?�7P?��?��>M���;�A֘>�:�>�X������oa>1zJ?b�>�\?���?Y^P>��6��ܪ�W���Vm�=os>c�+?�0"??�J�><	�>L�����W=S~�>�*`?<�?��l?���=]�?#6>���>.��=Y˜>]E�>��?yN?z�p?=^K?��>C��<��������Hnk��NJ���;�)<�?w=�d�ぽ�޼�  =F<콅�YZ.��6�>�J��/��E5<'D�>�u>e���NN/>�xþ݀��d�>>5��� ���A΋�l3� �=�~>׻�>V��>Gy"�$��=���>���>�e�b�'?��?]k?��_�T�e�2%پ�N�ű>��@?���=��j��䒿��t���y=�
m?ý^?(�Y�,���O�b?��]?=h��=��þ��b����e�O?;�
?1�G���>��~?b�q?P��>��e�*:n�'��Db��j�0Ѷ=Zr�>KX�P�d��?�>l�7?�N�>-�b>%�=ju۾�w��q��f?��?�?���?�**>��n�Y4����n��c^?��>�y���?y]@���־�)���ʁ��bپ$͝�Qu���� ���3*+�Х��;�Ƚ6�=�O?O�t?�Ro?��^?�q���d�,�[�4}x�L�Y�?��W��2�I��6B��bC��k����}��Մ����W=*��w_�WO�?u�4?�d����>� ��~���'�����>�]G�L� =�#�=����)��<��;nV�8�
�������?Î> ��>]>?�`Q���C���dc$�L���p<>��u>u�y>���>x�='4�������E�(�'���v>|Ic?��K?�"o?�S����0��ځ�ǔ!�9�0�����G�G>�
>>��>��S�Ӕ�'�%���=�n�q�	p��ߏ�
�:z=�2?M�>�ɛ>���?S8?A	��$��y�$2��tb<3�>>j?�3�>B|�>)>̽ ����>S�l?��>�>p���LU!��{�N�ʽ�+�>�ѭ>}��>��o>�,�Q*\�ug������9�+��=�h?Z�����`���>R?��y:�B<�}�>Xw�i�!����'���>�}?+��=��;>RqžZ���{�4K��G�I?R}3?X�^��#��V�>T[?{�?nT�>A��?\��>�f�J�7���?#�P?isK?p�@?K ?)�L=�f��������Z3��E>>��>�FT>q-�=W۽��p��]a��?��#�5���=*dd�irF=��g���<=uϳ=z��=f�ڿ��J�%�ܾ��}���S�OW��L����t��M&���D�(��)
�7����T��a��T���3u��Q�?�e�?�u���l��P���H���F�`�>@`��}z�f��R]��z�����⥾����>N��6i��a��'?�����ǿ鰡��:ܾ4! ?�A ?)�y?��R�"���8��� >B�<�/����뾝�����ο�����^?���>���.��t��>㥂>�X>Iq>����螾�,�<��?!�-?���>�r� �ɿX���
��<���?�@�vA?,�(�~���V=G��>��	?��?>-y1�'B��ݰ��^�>�>�?���?�8M=�W�
��ze?Ԅ<��F��ۻ��=�H�=��=|��3rJ>nW�>-f��qA�lFܽ�4>
ƅ>��"���}^�h��<�y]>k�ս���DՄ?z\��f�x�/��T��!M>�T?+�>�8�=�,?�8H��|Ͽ��\��*a?�0�?��?��(?7߿�o՚>��ܾ��M?4E6?���>�d&���t��v�=X�M������%V����=���>��>Ȁ,�Ŋ���O�`u�����=��������k�8��.�j����kC=���1��6�5�Ԥܽ��i��&�)�B����=��=�mM>V��>9�>�[>7dG?M.^?�߲>R�@>�)���`f��p��	�=�3��G�������覽;����#�3����X�*"�y��AÎ� �Y��(���f�n���:�9;�ù0��7?�:�=j9	�Y�H��%���}g�I�:�����W���J�����^?��?x���ߗC�sr�EK�f�m� �O?g� ����-�̾�Я<E���߽Kj�>܅¼ɽ�� �4��A�x�&?�+?����C���9l>A'�����<�%?)b?ٛ�G�>C�?H.���i���A>�>�۫>�'�>��@>Yx��{@u��$?iR?�9�����dD|>"��w<��w==���=b��19�:C�>���=;�Y�l�=��K���T?G#�>ۻ*��F�j2��<L��C2=SUw?g�?�
�>ڽj?AZB?N!�<�q����R���X�=<7W?��i?\�>��w��3Ѿ�^��c5?�\d?�R>7wg��i���.��8�
�?No?@�?;��7 }�G���S���M6?��v?^r^�$s��f��"�V��<�>�[�>���>�9�Xk�>��>?�#�XG������1Y4��?l�@D��?�;<��`��=�;?{\�>��O�d@ƾ�w��򃵾��q=�"�>U����dv����Q,���8?���?��>1�����gݺ=S�þ7��?Aӑ?Ƴ���U�ѳ���}����>u>��=A>�M���&�����,�%�o$���F���>�@���=K	�>:��.ȿY�׿��X����g�־Ql�>���=H|=X����� ��N�Y�y���������c�>d��>�����^y��gf�-L�a��=q�>��	>ȱ>y�<��+��4J��y������>)��>͖�>/;��5��,(�?�ߪ�L���㗿�rྋ�4?*w�?�=�?d�>1�>�D������d�)��GE?�Q}?�0?�S<��Ѿ�N��j?�J��tH`�ͅ4��:E��EU>3?)F�>0�-�+�{= Z> v�>�I>�0/�5�Ŀ�ζ�L�����?w��?�r꾪��>ڀ�?�v+?(m� C��Q]����*�m] �S,A?��1>�|����!��2=�*�����
?�0?@��G*�j�_?��a��p���-�Oǽ|��>�u0�oB\��e�����me�����_Gy��?<]�?�
�?���#��%?Jٯ>^���%�ƾ7`�<yj�>���>��M>��^�nu>c����:�Ta	>���?.{�?_g?����� ��i > �}?$�>[�?;g�=�\�>�c�=X氾K-�Ep#>�*�=�?�8�?��M?F�>a'�=f�8��/��VF��AR�����C��>&�a?�L?�;b><b��(<2��!�"cͽf1��P��S@���,�$�߽�+5> �=>z%>��D�c	Ӿ��?p�̕ؿ�h���q'��64?E��>��?�����t����<_?�r�>�8��*��-$��1I����?�F�?��?8�׾N�˼Z>s�>2P�>[�Խ#�������7>��B?I��D����o�/�>���?_�@Ӯ?�i�.	?���P���`~����� 7�z��=�7?j*��z>t��>-�=�nv������s�L��>YB�?�y�?���>��l?<�o���B�C�1=HN�>��k?�t?��q�P󾓳B>��?C��@����I��f?e�
@�t@"�^?뢿k=������Ⱦ�dɾJ��<�{�=�k>4����<�[��l9��$=��ż���>~�	>9��>���>Z�j> w0=�������ȿ2��������P�|��Re�<��]о�2>��)���E��Ԗ�e���,|�����,mQ����!�=��>?�X?3�w?��?5C���8>����@<�̽i��=�>ģ8?��<?��?��+<%����e�dw��y��sf��b�>9(>rS?}J�>���>=�@���>��.>��>��\>��N<ɸ�::�<s��>�1�>m�>
�>{
5>��>�봿�\��_i�u���˽�ˢ?����^K�k������j���>M�=;J-?�� >P���#�Ͽ/R��U8G?v7���Z��b-��>W�0?i{V?	�>x���iG�	�>���{�j��>/L ���n��*�:P>�N?ү�=�Sc>��/��q%�m�_�� ̾ǩU=�LD?�T.�|��;��v/^�e�	����=<�1?�&����������Q�q�������<&.>?�O$?թ�5�����V��@>*�>̡����w����>����tu+=�+��� :�8�:�!�>� �>�TS>yG�=�
�>sc��D,2����>1�N>^�t>�>?N�?������O�ܾ9��YU>���>+��>?D9>X�<���=zf�>�>\��;tž�����f���_>0�;Qe������_�=�����Si>�=�=O�$<��z�y���~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�d�>z��Z��N����u�#�#=��>~8H?lT��.�O��>��w
?�?�_�f�����ȿ{v�z��>=�?��?��m�&@��
@�$��>��?�gY?Ioi>Ih۾ eZ���>��@?�R?e�>�9�d�'���?'޶?��?��M>���?�pw?���>���n4.��J��2���4=��+<^��>��>�Ǭ�>�9�@��N����?r�>���NY>ա7=z�>A�߽'W���:�=��@��¡�����9�>F��>�}[>2�>���>��>�ϐ>Vh�<�[��Vs��X����K?���?+���2n��N�<:��=�^��&?�I4?;k[���Ͼ�ը>�\?i?�[?d�>8��P>��F迿3~����<}�K>*4�>�H�>�$���FK>��Ծ�4D�Zp�>�ϗ>�����?ھ�,��%T��EB�>�e!?���>�Ү=ڙ ?��#?��j>�(�>BaE��9��U�E����>ܢ�>�H?�~?��?�Թ��Z3�����桿��[�v;N>��x?V?sʕ>a�����kE��BI� ���]��?�tg?VS�-?:2�?�??a�A?�)f>؇�"ؾ������>��#?�#����>���#�9R�:� ?��?���>x��Iڽg�0�T���(����
?�_?~�?
���(b���Ⱦk�=J���X�b��Mv<�H��(>�>�吽]��=H��=���=C�i�J�/����<��=�e�>�	�=��J�j5��.=,?�G�Zۃ� �=S�r�?xD���>.JL>���i�^?�l=���{�����x��U�� �?��?k�?���ŝh��$=?��?(	?�!�>0K���|޾���Pw��~x��w��>���>�l�v���������F��c�Žx42���>��>�d?�.?�<>��>�꘾-�� �ʾ�X�O�j��"��O
-��!�'���ꤾ��Q�V�D��Ҿto�� t>򺟽ݯ�>q\?M��>�@O>���>����d��>.&�>�}W>l�M>K�E>��f>�>=�h뽷KR?]����'�U������3B?�qd?+1�>�i��������?�?=��?�r�?�:v>�~h�h,+��n?|>�>���q
?�S:=�)�Y9�<V������2����ժ�>�?׽� :�PM�qof��j
?�/?b��ȋ̾V:׽n�����n=�M�?I�(?b�)���Q���o�9�W�pS�f��J0h�(h���$���p��쏿�^���$��{�(�xn*=s�*?��?���@��"���&k��?�k^f>��>�$�>3�>�zI>M�	��1��^��L'�<���S�>,[{?���>�I?>�>?�CS?��O?r�>xͮ>����#�>�&߻�Į>&c�>�y:?R�/?��.?A?� )?HXi>���t���,ܾ?y?)?��?�>��?�fz�u�˽���eټi����������=��s=����]�v�tGq=�e[>v��>=����W���{9>b��?��>�v�>�M�4���i�<�?���>�><��X�k8��4���)?Ĺy?�D�=92f=ڃ9>CF�=X�,=���<)ka=A7<\�=	z	<�zw=�@D�8@I=0��<a�<QHn���=��%=v۽t�>��?���>�B�>�@��� �2���f�=�Y>�S>G>3Eپ�}���$��	�g��_y>�w�?�z�?c�f=:�=|��=W}���U��I��'�����<q�?�I#?�WT?��?��=?qj#?F�>�*�M��}^�������?C�8?�r'>(���^�!��/���L}�"r�>p��>�Ky���C���G�F�龊�J=��>mL���/e�ޠ������YV�3�����?��?��;=�����I���6��y�3?�j?;�Z>*T/?+z־�`����,�­=�?�8V?�D�>�cy?�
�?�s?��*?��������¿�堾x��>[fN?�J|?]��?�c�?/J7>����g�@�%���� �<0ٽr|�Aac;���=YL�>�^?�>T��=f�%='1G>�_ĽV~�=�>�i>���>�,?m�>��=C j?K� ?%ɀ�����.yH�e$��d'>JhZ?�*�?oZ$?���s;��m�>ZѾ���>q��?ƒ�?A�9?�f˽� l=��ֽ���������>�~�>�5�>����཯��<ě>s�>3>ս����<��>��=?�;N?�{�=Y���t	��և��$��Aþ��=6N���>>��̆��{�����s].���4��gվt�a����T2��ì�����>�ǅ=�Ef>��=���=�/�=���=�O�=�D/� �=�>�����n����=�zk:|ac<����T�&>�Sy=A�˾͉}?�7I?֒+?��C?��y>�>>M�3�Q��>�����@?�V>ɨP������;�򨨾[$���ؾn׾,�c�!ǟ��K>_I�U�>�:3>Q?�=
�<k�=75s=�Վ=:lO��+=0�=&P�=�}�=���=c�>pQ>�6w?L�������4Q��Z罈�:?�8�>n{�=o�ƾt@?h�>>�2������~b� .?z��?�T�?5�?Hti��d�>;���㎽}q�=l����=2>��=>�2�,��>��J>���K��򁳽�4�?��@��??�ዿѢϿ�`/>��52�:�cX��4�7N�"�J����&?�>��>�,��]W>Er����|3����="Ɠ>�D>�������u�=�l/�C��n#=��>M�{>+��>�Hr��L��R	�Cݐ>�N?�l�=z��xꎾ�9>
�,>�>��>x�?��?��C?[ss?�,�>��ƾޖ�d�ɾ�>�>�*����>���<��>�(�>��N?�?�H?���>��*>� ?�i�>��?�i���9�;��A�����=
�?� �?Ś�>y9-�=���/�ϱ,�7�Z��?x	F?���>�a�>���V)ۿ��+�M�/�������;�S�<2�_���ּ�c��#�fN��G5�=���>�ӻ>�k�>��>��F>�Lv>]F�>�>�k<�ԁ=kB�;��<Y�:ZЁ=E���l�����kn=۸�<	�����ܼ2��$�,E�<k�<���=��>}>���>z�=�	���H/>c�����L�b��=G���;B�d��/~��.�4�6���B>��W>���R3��=�?*�Y>�a?>��?�Ru?C* >�#���վD��#�d�L7S�/��=�->��<�pa;�H`��M��pҾ��>�c>S6�>T��>Q���gD���(=��侰�<�p`�> _����!�t� ��C�|��8����b�uFȽ0�,?�T����=�e?86@?���?Ƙ?��<�T��F�>�#5�Զ�=( ��.c���[��%?O�?d��><񞾏�%�oξ������>�K��P�|;��lB1�A}���c����>����ѾYa3�C��`莿 �@�Q�l��5�>x6O?&>�?�f�YC��{UN�kh���x��%?�e?���>ў?��?�����R쾍ހ���=Ko?`w�?̵�?#�>+��= �d�>�_
?�E�?��?�*r?=�=�U��>®ٻ�Q<>�w��eK�=�L>���=��=sX?��?�<
?7����	�ﾀ>�J�b�Dx�<��=5��>��>S�`>m��=x =�K�=��]>�*�>芚>��_>/��>n�>�'��w�!�'~)?s�x>���>J�?ӞI>f�!��^��:�>��y>M�[=p)��g�h��c�����|�.^#;�*w�Hm�>'�Ϳ}��?�\d>о��L�>1c�]h���On>�x�>7�ӽ�R6?\��=�9k>��>�j>�J$>��>8ie>�TӾ�g>����d!��*C�>wR�l�Ѿ܎z>E����!&�n���L��RFI�|���_���i�y&���-=�x�<A�?����V�k�B�)�w����?�j�>�6?Yጾ̊���>'��>ɬ�>�Q��k���č��jᾟ�?>��?75c>��>�W?��?p�1��.3�7mZ���u�0A���d���`�V܍������
���Q�_?��x?cwA?S�<�Az>&��?��%�s̏�*�>p*/�=;�� <=�"�>���Qa�'�Ӿ\�þy��F>��o?J$�?�K?�V���m���&>�:?��1?�Mt?��1?C�;?�����$?�3>NL?��?>K5?��.?L�
?o�1>��=�d��P�'=���[֌ѽ�<ʽ���?W3=��{=`�7G�<= ~�<2�＞Lڼ�D;�w��sB�<��9=��=(K�=���>\^?D��>b8�>]J7?j3�ڂ5����(0?�-C=.���o�������e񾿁>�Sl?�ݬ?��Z?5(g>��B���E���>jC�>\B(>$�^>b��>�����J��x=�;>UR>�Ȧ=�KW��邾���ƌ�	7�<�� >b��>�\m>�-��>>)/��Q���:xW>�R�:9ɾR�U�vF�53��	Z���>F�F?6?�y=�f��_����g��%?M4<?uLM?���?���=�$׾��@���A�0h���>^��;/0��4���_���:�9n;1��>�h��pC����(>�K������n��	>�1����>�	�^�<Y����ݾ�6��]>���=��+���Z��������??*�<�u���n,������,>��>G�>�e�Q����<��)���g>���>�_> a�=�s⾯�W�]i����>=�R?�p?)�?���a~���U��g��ž8��r
?I� ?j�?=2>�RN>_�վ����b�H�;���>n)?6 ���>���G��1���S�9�\>,��> R>��
?G�Z?[�?�a?��?���>�c|>�Fӽ�贾9A'?ĝ�?P�=7�Ľ�*M���6�}�D�eZ�>�0?�4��)�>�U?�2?�(?�NJ?��?xq>�d��&�:�ን>�V�>5�Y�����_>��K?���>$mX?U��? =>��5�$߬�-����i�=μ%>�?3?z� ?�e?(��>��>�݄���!>;��>�3�?j��?`�l?r�q=Zl??��>�B?2�?����>N{�> �&?�j?|�?(�C?E�?q��e�1bQ�CE�of�=��]=����o="��bE =|�"=J��=T�8�g�7���W,���.0=��J��>$�>l���	>���������5>�
�;�x�"������U�=�DR>|��>i�>�K/�$�=��>�j�>�@"�B-&?��?��?iS1=��f�?;��ჾ ܿ>�j<?^��=y(a�� ��a@|��P�<��l?d%W?��b�3!��2�b?X�]?0g�F=���þٵb������O?��
?�G���>��~?��q?D��>]�e�9n�=��rBb���j� ж=�q�>W���d��=�>՛7?�P�>Q�b>4!�=v۾L�w��o���?��?a�?@��?�)*>%�n��3�f@����RX?��>,��C?�5�9�bѾ�U��w��b��KাI����x��蝾˕(�k���h�ͽ|�=�g?�+l?Pu?%�`?q���vb�G�_�{x���KW�������
qA�A�i>=���i�f�b����j��*�9=��q�02\��Ʋ?[1?�&��N�>U�M��	�!��Gx�>�ɵ���/�>K�=�w#�Ax�<y�6=,H���,�y3��M(?Љ�>�C�>B�9?��V�i/:��-��4�?��[�=8��>�ń>p��>�g=�鋽W4D�_�������O'v>|c?!�K?�n?t?��11�����>�!���/�HO��A�B>ݎ>e܉>^�W����3&��R>���r�����o����	�z�~=p�2?��>���>�K�?�	?qx	�<\��[dx��1�d�<�4�>li?<N�>U҆>:�Ͻ~� �w��>�jl?E�>t�>�Ӄ��R%��x�j�����>�Ѭ>Ju�>�`t>�R��]��� ���_3�b�>��e?����Y[�-؏>y�O?(p<<���i�>�����"�sC�^B*�AY
>$�?��=��>�L��F��D�y��򑾏�.?+�?Ђm�h(��Q�>K`-?�'?�!�>PA�?�|�>����#�ƽ?��a?��Q?0�Q?2$�>��j=,���*�佒�S��jU=�%�>�F�>{ >���=�)��r���`�(��=!�=��"��ʽ�M�=S�=�W��i+=.2>[6�ZR��&�۫��E�� �&∾.�w�rr�p�6��5پ�����f���ZQ�<���>�~�1��ݬv���e�4��?�j�?;����,�����A�{��l���>}�Q�F^��|�����F՞�m"���䟾�!�F�S�T�O��&i�H�'?�����ǿﰡ��:ܾ0! ?�A ?6�y?��:�"���8� � >�B�</,����뾥����οE�����^?���>��/��[��>奂>��X>�Hq>����螾�2�<��?0�-?��>��r�+�ɿe���Ĥ<���?*�@�wA?q�(����
V=���>׍	?9�?>tV1�>��찾3M�>�6�?�?�M=�W��$
�.e?�<��F�lݻT#�=76�=��= ���J>^[�>�q�fPA���ܽ_�4>!Ӆ>�c"��c��r^�},�<�p]>\�ս���[Մ?�y\��f��/��T���Q>T�T?�*�>5�=�,?i8H��|Ͽ��\�6+a?�0�?n��?��(?�ݿ�c֚>��ܾ1�M?�D6?��>�c&�t�t��=<��������8'V�;��=���>6�>s,���>�O�z�����=N�������.��]����7����H!��pʽN����E��׾rg� D�h����V>� �=�X>gb>�<>X�J?�cO?\�>�.&>�H��6h��	۾V;��v���׽u��}�ݽ�E�� ˾Vʾ��+3$��l�DȾX#{��d�<�V��V����X�+26�Xo"�s�A?�j�=�7����e�X��N�#�K���H�=Ffu�sF�nʾ w\��~�?:�?x:���.r��羮u=��3=�mv?'y��0Խ�	����p�iLW�w�I>l�>��*>^㢾ӸǾ	ru�a
;?6?U���[j���=����,>�}?��>������>/�?��`��l�V�>�b�=�B�>�q�> �>es��Y[��T�)?J_L?)	*�Ѭ̾�{�>oؾ�I��=�v=�q�F�=G<>�=c^]����=��B�g�9�� 0?�S5>q+��h�o�;���㼜��<�C?��>5.�>wBb?�A@?�0���n��+�	���W>m(H?��t?�c�=�����߾A6E���@?��z?��8>�*.�هھ�Ia�y����?��G?!�>?�5�~�z��&t����T?��v?�r^�os�����W�V�4=�>�[�>���>��9��k�>�>?�#��G������vY4� Þ?|�@���?��;<��6��=�;?a\�>�O��>ƾ�z�������q=�"�>���~ev�����Q,�Y�8?ˠ�?���>���̩�E!>U�¾��?�K�?��f�gr6��ؾ$䄿k��:�<����B>^_�<q��W|Ӿ���@����¾��e;�ʓ>�@i�����>j8��h�=>��n�M���^��19?z�>�6����ǽ�$������i���e6���~F�>��<>�} ���z���T�Z?X�A������>��<��>�BȽ�S��g�m���9��8>t��>�=�D]=t���̟?4��&ӿڧ�D%���@?�q�?��?[?�3L<�<!��bξ+$Ӿv/?de?cFI?��@�z5��Y�#�j?M?���K`��4�:E�i%U>�#3?q7�>ن-��F|=  >���>vi>7#/�ÄĿ'Զ�۸�����?؈�?ym�t��>W��?dv+?`l��=��V����*�m���9A?1 2>~~���!�/=������
?i�0?�g��1�]�_?*�a�M�p���-���ƽ�ۡ>��0��e\�9N�����Xe����@y����?L^�?i�?޵�� #�b6%?�>`����8Ǿ	�<���>�(�>*N>oH_���u>����:�	i	>���?�~�?Sj?���� ����U>
�}?�8�>�ń?���=�2�>�8�=gM��]��r >���=�;@���?�*M?}�>7Ϲ=~�2�!/�rC��O�$���#D���>xXc?sPM?"�a>��ֽ�OI���"�g�½�+�E�ϼ�A��U�}���`4>��?>�`>UrB�*�׾��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Oz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>;�>�I�>A�Խ����\�����7>0�B?[��D��u�o�y�>���?
�@�ծ?ji�`	?j�'O��'_~�F���7����=C�7?�*��z>���>�
�=�nv�.����s����>:?�?�z�?g��>��l?�o�X�B�}�1=�D�>��k?hs?��j�i�o�B>��?<��U����J�	f?��
@*t@�^?S�ÿ�2���?���O��(��;1>�v> �!�(0���bϽ�k	=;��:=Kx<�K,>h��=Ď�=�a�>��O>�^R>9�����7L���靿i���+¾����`����+Ⱦ��ƾ�5"�//������'ʽ� }�\hW��0��~GĽ��=;�U?�R?1p?�� ?@7y��>������=�R#�!Ä=�T�>�q2?ݨL?r�*?�o�=ʨ��&�d�s[��=;��㾇�1w�>�EI>}�>jM�>� �>B�>9,�I>�f?>^��>� >�'=պCH=q�N>�Y�>d��>�w�>F��=��U9��6Ӵ���k�_�ν�K�T��?����(AN�@���ը�S��ߥ�>o7�>���>�����)��}宿�6?vы��k�9��< ��=�1?	�D??X=�W�����2�>7#��/<�>,0d<��=J{3�7��.X-?a��>i �=g�"��o�=,X�z�f��>u�4?��ľ�L��W�a��9���H�>0*�>��T>�5�j����҇�c���債=��8?��>��;�s����M̪��F�<�A�>┉����<�>$!��ځ���TҾ�o�<,�f;I>��?�/>t#=@��>����bA��5��>��X>]�I>�v2?�?x��e�����z(���b>���>U�>2��= A	���=�`�>3�z>`v:��\�o ��l�[�Y�6>s�콨��?�����<.��IӘ=�Q��n�G�H�Q�4J���~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ>h�>�x�Z�������u���#=;��>�8H?�V����O�>� w
?�?�^�ͩ����ȿ|v����>T�?���?P�m��A���@����>:��?�gY?�oi>�g۾�`Z�ʋ�>ѻ@?�R?=�>�9���'�|�?�޶?د�?�C&>�1�?*�v?��>�,���9�����7����=kܕ<���>d0 >�p�C���������'e��%��Gc>:_=AA�>�|��qξӳs=3Ü��k���);_ע>��r>�3>캓>���>���>Wru>���=b�(�c��S����K?j��?���[2n�PB�<֛�=>�^��&?�H4?�q[�k�ϾtԨ>=�\?s?�[?d�>f���>��4迿�~��J��<��K>-4�>�H�>a*��cDK>��Ծw9D��p�>cΗ>� ��|>ھ�-��l ��)A�>wd!?0��>�֮=� ?�#?��j> 5�>�@E��?��H�E�Qw�>Ñ�>�A?��~?��?>����P3� ��Ρ� �[�eON>"�x?Kk?d��>A���_���ڢN�/=I����8��?�Yg?=彪?V�?&8??^�A?�Gf>c���4ؾ����>� ?�r���-V�1�0��s��wD'?x�	?�*"?7�`��p��˚�=�$�p7���)?("_?='~?��Q��j���� ���A<6*�==�`R>H-���%�=�SY>�F�$�; �;I}>��G�;ａ�=��e>m	_<��R��g켓4,?�^F�܃����=L�r��vD���>OXL>;���x�^?�l=���{����vv�� U���?M��?�h�?'���h��#=?��?{?�)�>_A���t޾(��3Hw�tbx��x�-�>���>��p���v���\����D��/�Žv%�fL�>�k�>4�?-��>z :>uߪ>O�������澝��	�Z����;�	1�o�x�����="��¾~�u���>v�Q��f�>�?l�j>�\\>�y�>�E<�C�>�U>�8�>W�>�.G>Ot:>	�=T*;x����QR?����d�'�P��0���T,B?#wd?�/�>�i����	���u?�~�?�q�?�v>�uh�%+��f?��>E���m
?b�:=�/���<o[�����A=��Gg�o��>��׽�:�;M��Df��m
?�/?�6��u�̾.׽����;ho=�M�?�(?%�)�%�Q�"�o��W�IS�df�D"h�\����$���p�k>X���#��-�(���*=�*?��?G��Ѯ�.���k�c?�K�f>���>i"�>�۾>}XI>0�	��1���]�)<'�Pԃ�zN�>�M{?�R�>|,G?�Z9?�K?��P?�@�>n��>�x��X�?�۴=�v�>��>'J8?�0?PB8?�t$?�4?Lzi>Aށ�7���cI��S?}?t?�p
?�0�>�����Y���@<V�<@=i��I��R=�&�=�_�����!�W=��(>.y�>��S=%'/�s����>��?}��>tT�>y먾{���?�(�>ڇ�>X�,>�b�����߽�r?!��?.�y=�w�=�"\>[�0><Խ���x2>��޺�e�=�M4��M"��Mr=gݽ=۳�a�콷��<\���>|=Jn=�_�>!�?��>[/�>T9��y� �d���^�="Y>�HS>��>�Eپ�x��*(����g��cy> u�?�w�?!�f=�A�=D�=�����E��C��,����]�<��?BE#?�XT?���?��=?Lj#?\�>}��L���V�������?"x4?W�>O��| ��%�����>��?ec�>�)v��-�E�I�v�׾_8ٽ�h>���,to�O,���`�x���9#�A�?�?��?� �=٩+��a������پ5?�W�>;�>�+?Y>��Vb���}�*>`��>�_U?���>.��?���?f��?��?��A������9A�ʺ�>Ǭ?��?�
�?��|?��>����-��l.�\¾�L�V+�5y�����%>}�>��>�ɼ>�b>��>�7�<�̾Ҷ�>�K>�l�=��>3 ?�$Y>��=S�F?(\�>el��9��r���v��	����o?�̎?�-?��b=����B�V��n�>��?,��?��/?DWD��O>�0*���ľXg�c�>���>��>���=�� =ǜ>I�>��>�LA�"N�oY*�2����?��>?D�=��ӿ��j���0���~�T��s�&��k��8؛��B��N��1��&ھ��ƾe>�QE���`Ǿ�@K� �y�.L�>��x�uVy>��>���=�,��̽���	��F��=�Rؽ���=yC�;��=��ǼKi^=���q]]�����Ј˾o�}?;I?��+?��C?,�y>d<>1�3����>2����@?$V>��P�ڈ����;�p���-���ؾ�t׾��c��ȟ�1J>�ZI��>�43>�D�=H�<��=�s=Ǝ=R��=V$�=bP�=�e�=���=3�> T>�6w?Q�������4Q��Z罞�:?�8�>{�=��ƾd@?N�>>�2������ib��-?~��?�T�?5�?tti��d�>E��a㎽�q�=V����=2>���=x�2�?��>��J>����J��ހ���4�?��@��??�ዿբϿ3a/>���=ލa���F��GN�
[��O�d��V,�I7+?Ċ��t���^�=x��P����4��V�<)��=f8�<��)>�
k����=bu4=�=o߈�Ȩ�>�)�=3�=�Խ�$=>��>��=Wv>���&�ĽS.<��h��#�>���>���>L� ?D�?8�N?E}?z�>�A���Ӿ�t��n(?�ݲ>��>Y����>3��>˾w>��<?#8u?�E�>��>�*�>-��>ָ8��䁿$�����!*>}z�?�?�?.��>����x�)N#�D#��;�V�>��F?G��>U�>�U����.Y&���.������<��+=�mr��QU�Q���in��㽐�=;p�>���>��>aSy>��9>��N>��>�><>�<Io�=�ӌ�ĵ<���:��=*����!�<�użk���&���+�x�����;>��;X�]<��;���=���>�2>z��>j�=�ѵ��%>%����F�c�=�����@��b�^�}���/�s�,��TF>�{\>n`��
�����?+_i>��J>�D�?�yr?&�><\�|�Ծ1����k��}M����=٫�=u/M�.65��"]�D`L��˾<��>9�>k-�>D�l>�+��0?��ax=����e5����>���p������,q����ݟ��h�.���lD?�L����=�6~?��I?��?�l�>ph����ؾ@)0>��X�=m��!�o��y���?J'?�|�>��뾢�D�%�žd{�����>7�H��M��G����-�V���j��ѩ�>��5ξ�z0��������<���z��ɿ>)�L?vC�?�i��3��idR����w��B?y�l?Ȉ�>1?�&?�̽HG �&R}����=w�k?5��?)B�?���=���=�k�����>�?�ו?!o�?��n?��;�!��>n�*=��)>�K��=n$>��[=>3(?b�
?3`?h���X���*��F��.I���p=���=�q�>7it>��d>h��=��<Ͼ�=\^>�ή><ؓ>U�P>	�>�J�>3þ���� ?[)d>gp�>wF?�j�>"T��ww;�A��>s����ں�D<Z/;ޫk�.�=�>=5�=f�=���>�w׿�q?{f�>_����>�E���ɑ��%�>Mv�>����'�8?�>�َ=/�?O;�=��>H�>I�>D^Ӿ�`>���8f!�;1C��zR�w�Ѿx�z>����z&�I��cv���UI��x��qe��j�y*���5=���<$B�?>�����k���)������?�X�>�6?�Ɍ����M�>���>߻�>R��q����ƍ��f�
�?���? :c>��>]�W?֙?\�1��3�guZ���u�]'A��e���`�<፿˜����
�[����_?��x?LyA?�H�<�:z>���?��%�ҏ�9(�>f/�?&;��9<=L+�>�(����`�ڭӾm�þk:��KF>D�o?%�?
Y?�PV�ڳI�S�>|>?�#9?f�x?�+?e<:?c��P�)?��J>,@?x�?��6?��+?��?)>>��>�<�?=��p�q�����½N�ƽ�(�#`�</:�<p6�?z<�F=�\=ف/���M��<������<p/=��y=j��=�ؔ>�i]?��>%�O>��7?���F���@����P?&u=>�m�8YϾ%��&����h�g?��?m�K?��{>�F�m�X��>hDv>�E>,��>Ͳ�>�Y�J���O�#>/E�=٨�=��>�$�c��;�����V��<��>���>�>���'�=����_��^�l><��RW ��N��3\� =8���t���>/�9?�>??����T���/��t�B�$?%uO?�Z?��?$>�׾�?�8�9��E��v��>��X=uj���謹4��-��h��=��>�3�?���u�>�����;t�	7�VǾ"��=v׌����=M�%��վ�~꾟�;7��>�������y������37?:ҹ=ș��E��R���V�>&��>ϭ>���G
}�AH�T�o�=X?,�>c�>����R���C��}>�@?�l?[p�?�(��fs�S"�M�B�ž͛d>8'?�op>v ?�/�>���<Dw����� |m�}=����>幟>0�!��.^�<赾�þ���n�Z>=�>��=�,?�P?�F�>��p?��??���>�)j>`�`�(>���K*?�,�?iF�=�}ν%Ś���:�5�*�_��>��Z?���t9b>Ӯ?x�+?�|*?�L2?�Z�>��{>:����
��>Q�>�p�?	����?>V?�>H<F?�я?0o�>��m��"��D">�R>��=��K?�F&?��>K�>��>!d��>&?ˆ?�nG?���?��
�p�>"+t>��$?��6>���>LD�>,��>69k?�:�?�td?�%=?�ԛ=j�2�`~;�T����'B�^m<��=�b<'��Eۀ;��<��>O�����=���=��Ѽ�����-�-}�={}�>��{>Hz��%�$>����e�[;>Z6��ꔊ�p����6� ��=��>��>?��>'���=֟�>"��>�c��$?��?��?���;�;d�?�׾9M�N��>�.C?���=�Rq�t��?�t����=�k?��`?[������e?�]?J����2�N�־Jb�*iþ�1B?R�?��1���*>g?Q�[?�)�>�f�8�c��!���WV�b;�����=_Z�>���J�C���>��H?���>_ۀ>��<ݾAl�>ֈ��F%?ۉ�?R�?�L�?��=�
��V׿g�Ǩ���a?A��>�̕�?��=�Hվ^����`��W�ξ���������\.��j��ߑ���P#�#�=�?4Aj?�{?��k?����6Zb���j�g&���P�(-����y�.��0B�h'I�<r�L���D�p�f��@W=c�u� lE���?�^,?t����>}�x��o󾂪Ծ�dK>&ܓ���񽳢�=0�q�Ȇ=W�U=��h���P��׮���?a�>���>�E?��V��>�u;:�i=�P���i#�=�ܐ>��>��>���aG��x"�R���^Y�fBýn��>{r?v'r?v�z?n2�<a8n�؋�pD���@������if>�ߩ>b��>|S���u���4�m�T��tb�̸�������u=��	1p?���>G#T>�)�?��n?0�[�0I���ƽ�
���/>��~>6�?��?�~>,��=H
оm'�>�Qm?7
�>���>�x���^"��y}����R�>�w�>3��>k�n>�+�a[�����7��W99���=��e?a���m_�X�>1�Q?�����8�:�@�>�.�0��/H���!+�;�>Mc?Ǝ�=0@>�������z�ߌ����'?�$?恾�3�īt>;Q$?���>!Қ>/�?5�>?X	�O@��-?��s?<�H?�N?U%�>R<�<�;)�q���ҊT���=x|�>L��>��=�>	�M����+t��~ž=V���sĽ�Z���n�=���=�$�<=�i>�տ��b�(Mþ˃&� ����^�J��9>��;���`C��\a����־7G�����0}-�dD��h��i�C���?���?�@���q���u�g�#�۾��>�G�=�=����;=�7��Z�"��'r��� ���+�1����R�Y�'?=���ɽǿ̰���:ܾ=! ?�A ?�y?��V�"���8�_� >_E�<$��!��z�����ο̧����^?p��>w�h-��p��>|��>7�X>3Hq>w���螾E6�<y�?��-?���>��r�)�ɿ^������<���?"�@_BA?�m(����;
R=S'�>��	?F>?>G�0��B��Ʋ�ұ�>* �?{׊?N�Y=��W�����d?�z�;�F���»-��=8V�=��=�u��J>yX�>�����?�ߓؽ$U6>_�>Gy&�H��NA`�:�<m�[>�ҽ�5��/Մ?�z\�^f�x�/��T��U>��T?�*�>�;�=��,?o7H�o}Ͽү\��*a?�0�?���?5�(?ۿ��ؚ>��ܾb�M?zD6?��>�d&��t���=�9����K�㾡&V�N��=��>�>��,�ϋ�k�O��E��N��=�D�^�ֿn?#�E��$,�=>���9��z�ԽS>W����$���Ծ%�{��A� ��ｧ>t2�>��T>��h>}W?�6I?RH�>���<�½��c�����vL>#�p�2��۽�3��N!߾�a���Ė�����)���k�Ծ;��c�Y>�?L��t��uYw�x��U���M?�?t�`Bƾ3��^�!�K�u����=aB���j�'�{CO�z��?�?�"��y�,�Z]��A!<О0��{?+��~����k���=8��x�>�@�>)#=�4���G־��7���(?�?(�ɾ�ã�ђ >��*z��/?oo?���=���>�@?,��K%�M->�+>g�>đ�>k�>�*��L ?��H?<��R�¾���>a¾d��;�=��>��`������%>��e=/Ԅ�M�z=@
潎͟�DA?Y��>�)4���(�It��{=��j�n?�Q�>m��>ouN?�7?��r=����4�u �Pg�=ˊB?�de?S��=t+��㞚�Ƚ���-?��l?���>�{�� �����(������.?�?��/?$Ǆ�8k�S������C?��v?Lr^�/s�����z�V�p<�>�Z�>6��>R�9��l�>đ>?�#�nG������
Y4��?V�@��?��;<��D��=3;?�[�>>�O�=@ƾ }��	���z�q=k#�>C���Dev�����Q,���8?T��?���>��������	>V�ܲ?�O�?�l1�o��K���ȍ�f�"������4>U>���<���*�=�_��=��������>C%@Un>n��>��e��ÿ���糮���Ͼ7ꃾ4�?t\4>�^�=_���m$��^\��x*E����(Ἶu͙>��d>ȷ��㏾Hz�~�;���,=�/�>!>�!�>Q��K�ɾ(*�t�<�`z>Si�>�m�>&�⽅̭��%�?Z7�H�Ŀ�ȗ�(�Ǿ��f?z��?��j?�(�>�E@;F(e�󇞾���bR?�p?=Oz?\���/`���C�s�j?d>���I`�Έ4��1E�YZU>+3?�'�>�t-��7}=�E>���>�8>/���Ŀ�ö�5�����?Ą�?�V꾆��>�y�?�l+?dd��=���R��Z�*��>=��=A?}C2>����ޫ!�>9=�妒�&�
?��0?���%,��_?8�a�C�p�5�-���ƽ�ڡ>Ԩ0��T\���������\e�f���e9y���?�_�?��?���(#��#%?p�>(����0Ǿ/��<���>R0�>�AN>��^���u>��+�:��x	>p��?�}�?�k?w���D���Z>7�}?�޶>��?��=�z�>H��=�毾Re8��<#>���=�3?�;Z?��M?���>�r�=�e8��/��)F��R�I���wC�s=�>c
b?goL?��c>\���ۼ)�Z !�[�Ͻ�L2�hK�rQ@�&�0��ܽe3>��<>�> E��}Ӿ��?Hp�6�ؿ�i��p'��54?+��>�?����t�����;_?Kz�>�6��+���%���B�]��?�G�?<�?��׾�R̼�>6�>�I�>K�Խ����Q�����7>/�B?m��D��s�o��>���?�@�ծ?hi��	?��P���a~�r���7�Z��={�7?�*���z>��>?�=ov�4���	�s���>B�?�z�?6��>�l?-�o���B��1=[J�>��k?2r?�to���}�B>��?������LI�^f?��
@<t@[�^?���h��M��� þ�����=>�LI>79�w?>�6���g��j���~E=е�>�w�>Qi>�5\>l`">���=q0��%�'�œ��S����z(��6پVM�@R��L_���2�)�-�� ��ھ��ܽٔ���=v�]��=��W����=O}U?еR?��p?]�?�Ey��>����/Y=� �奌=�Ӆ>�:2?�
L?R+?��=������c�g��N����&��&�>�rF>1��>��>r��>�>�9��G>f�<>Q�>!��= I =�ͼ;�='�O>"i�>]J�>T��>}`>�&->�m��1Ī��Ig�q�a�8����+�?ȓ��mE��-��L�|�P�����=�??G�>:Б��@п�ٰ�1�A?�.��T����խ>v�/?�iV?-`&>إž�r�C4>c^�T}?�Ê >���a�B���1����=+)?䪔>��v>/h��_�R�m��ߏ�"���7|?�w��$��c�t���/���%>�l�>y��;�=���l�����*O��)��=�Z5?(��>�u�=`ݾ<̤�Ͼ���>���>"S�=~6����>aH"�-~�h�@��B�+�>�?[6?&�J>V�p<��i>��tP��?T>�>FZ�>�vN?�?��ɽy罀�Ͼ�'�G~�>���>�ɂ>��T>���2˯==��>�J6>��6�����,K����|�>e�=ⱬ���/�#(Ѽ՛���>���B =/u�y{���~?���(䈿��e���lD?S+?\ �=�F<��"�D ���H��G�?r�@m�?��	�ߢV�?�?�@�?��H��=}�>	׫>�ξ�L��?��Ž5Ǣ�ɔ	�-)#�jS�?��?��/�Zʋ�<l��6>�^%?��Ӿh�>x�~Z�����m�u�o�#=>��>�8H?+V����O�K>��v
?�?S_򾫩����ȿ�{v����>-�?|��?K�m�^A���@�~��>+��?�gY?�ni>�g۾D`Z�i��>��@?	R?n�>�9���'�h�?�޶?ޯ�?ίx>��?��?a�?�m0>�>�8-ɿe�ʿ�.��hs^>���>&�=|("��+��j��jذ��_�e�"��C���=x��>��\�)5)�}b`��s������+�=���>�*�>�CC=��F>詆>X��>�h>��<�C��I���<�K��$L?���?+���m�Li�<q�=gA\�
?�74?)a�/Ѿ��>~R\?壀?��[?�z�>����Q��e������ռ�<`�K>C��>�8�>:���)!M>��Ӿ=0G�<҉>��>aĚ��hؾ_G��`�Z�̞>: ?���>�ɰ=�� ?��#?�	m>���>�ME��3����D�r��>�u�>%�? �~?�?*���7-2�yl���꡿c"Z�hS>_Ly?�'?�,�>����c��\���l9H��\���e�?g�i?����?�k�?h.@?}:@?��^>N���5Ծ穽J��>��/?��ջ�88�Ņ�azk�t	?�b?��>Z��?C��P�v�Ǿ�}��^+?��?��+?�	$������}�hM
=+�<��J<�s�=8�Ǽ�	>
�0>;�K�k��3K�=�O)�/8a�:����={
�;�>w�:�h�ξ�n
>�@,?�!E��ރ����=K�r�|D�4h>O.L>������^?��=���{����jy��	�T���?ǘ�?�[�?;J���~h�]=?�	�?G�?B��>�g��nY޾Et�}pw��jx�G���>Л�> �i���˔������ @��UOȽ$�5��>�j�>P�?�s ?u#9>�B�>�왾��'�?D����*_��.�U�8���2�#��-���O)�H���ƾA�{�4x�>:����6�>��?��k>P�f>���>���<Z�>[�T>�=�>�ì>n�U>��5>s>��q��?Խ7�Q?~�����"�^�"���۽>?3e`?�:�>Z��;�끿.��~?�{�?6��?ދq>��_��2 ��d?޹?�����?f]"=.;���=�-����	�Yʓ�v���W�>�
�\�H�W�E�pM�e�?�%?f,����վ0o�	����Kr=e=�?��(?��)��Q���o�v�W� �R�M���Te�נ���$�Öp�8ݏ�q}����E(��d!=~*?�k�?������_���Fk��y?�H d>��>*9�>:D�>M�H>�u	��#2��]�7'�������>R*z?[�>"�>?�^?q-k?Ӟc?�cb>;��>����Qs?]�=O��>u!>�N?2�
?u�?H?dnN?)>�>�a=)������t? ?\�2?p�?c^�>a���K���Ƚ���=�NU��T��,S=��J=V����+]�d��=ҧ�=ê�>#mt=UO��q���>R��?&�>T�W>oƽ����j�>�Vf?>�>�/?�#�2��=̾M�>�{o?{��=�&�=��>y�=nᑽ��N;4�=SJ�k��=�ٻ�������#��aj�<��*�"��<�)��>H�=z,<=#p�>��?W��>�9�>(D���� �a��~�=�Y>�S>�>�Fپ}���%����g�&Ny>�v�?Ty�?��f=R�=-��=6~��nU������]�<+�?�E#?8UT?F��?��=?�j#?=�>�'��J��z[��^����?�;F?�9�>���
)�ɜ��SZ��6?ݮ�>ǐ���4������^׾$=��w=s���X�y�F��c����@����`d�O��?���?L&=s��f<ξj��?~꾉s?���>r��=��?ݞ4�%S���!�(>�?��@?)��>.�J?vi�?�-u?u'�>
�A�4]���������V�B>��J?��?�?��W?$�>7q+=E�-������Z���j�Ҡ%�Pvi���=�Ɓ>�S�>��>`��>��>nB;���4�������=\P�>*�>[G�> �?:C�>���<��F?���>�������Y��eք�}�s��Zs?kސ?�},?�k=����D�����>Ц?���?¨(?
�P���=��Q׵���q���>�b�>-��>�G�=2s=�R >L��>�F�>���w��(T3��a�\?:B?�H�=
ƿ��q�ׯq�����3f<�����d��7���[�$�=�Ϙ�	��aש�]�^̠��H���>��t3��R{����>�=�
�=[$�=0��<�,Ƽ���<�IL=N��<��=�m��2d<�O=�=o������**�D0V<��D=a��:�˾�}?Z=I?�+?�C?̶y>�4>ݗ3� ��>|p���A?aV>>rP�<���w;�t���m��i�ؾZx׾D�c��ş�{N>�I���>sK3>�M�=�E�<Z�=�s=���=�XW�4�=}U�=+V�=�~�=���=
�>�Y>�6w?M�������4Q��Z罍�:?�8�>P{�=J�ƾ�@?j�>>�2�������b��-?z��?�T�?7�?4ti��d�><���㎽xq�=޸���=2>O��=`�2�7��>��J>����J������|4�?��@��??�ዿȢϿi`/>�s>��>9A��uVw�a�(��M�<5�W�f?������V>��=��{���Ͼk����1>)�<��;�.��Q��=aٽ�2��5��"��>Ƀ�>�e��a�I=:��I�Q=B�Ԕ�>3��<��j=P�������m�=g�~�[��<.n�>�?`hC?
�p?5��>㾬�����8�����>ߊ�[Z�>�֑>�mW>�?�E?��>��4?P^�>�sK>�?�>���>Y'Z�C����h��Ҿ4p�=?[�?mߠ=��B�#��9����3�rn��(��>�A?'6?��?"E�ɛ���08�nJ�G�1�����|	=S��t�s��<+>!���M\��
�<eI�=�K>��?��>�G�>�e�>^��>�ʀ>,=�^�=�O�;�� �0�H��8u=BY;�)�$;�
P=���<V�6=ň'���O�<eI�=��K=+==���=��>�A>��>(��=����F/>�����L�ؿ=�G���+B�/d�&H~��/�V6�k�B>�8X>u���3��_�?��Y>\k?>��?�@u?k�>;*�-�վ}O��5e�]LS�SԸ=��>�<�\y;�'X`���M��|Ҿ���>���>[��>�o�>����on�NW�>�G�O�G�gN ??�;U�Z��!>=i�PL������|�x�s�$�|?�8���F<��s?w�C?'ד?h8?��=�������>���=�Ȕ>Uiﾘh��p�<T�>�!?�-?�e��o�)�Ͼն��w0�>:�O�.CQ������%0��|�Y�$�>1v���LϾt4�S�����KB�/�q��T�>`�L?���?}�P��{��)�L��������s?�e?˝�>�?�!?�����뾺劾���={�k?�a�?�	�?�� >Gt�=d;1��P"?��*?Kբ?L�|?��o?�"��H!�>�q�=�=�>#�j�*�`>��M��@�Rŭ>(�2?xZ9?��?F�ȽW;������羑�j���<�g6>�q�>8Vl>�as>��7>�=�
���\>��9>/�>��>� !>�=����M:��u-?��N>=k�>y??=�>DX��lK���\>��>$�Q��p����;DG����=!R��'�X�����>nտڕ�?S�>(��GR?��Ⱦ��<a�C>Z���<M�>?�Б���'>��>T�>^;r> Y�>"�h>�LӾ��>I���f!�03C��R�ļѾH�z>|z��l&���}n��VcI�8����_��j��)���)=���<?F�?�j����k��)�m�����?]�>�6?j�t����>���>j͍>�E��1����ȍ��I���?���?�>c>��>��W?�?��1��3��uZ���u�	%A��e��`�.፿����
�
�i��t�_?��x?hxA?j`�<�9z>���?U�%�7ӏ��%�> /��&;��A<=�*�>�&��g�`��Ӿg�þ�7��OF>�o?�$�?�W?uaV�V(��O�+>�?B?��@?)>|?L�(?#/?��&���?öU>�?6��>�0?T�+?�/?��)>#=>���<�Y=?�_�|q~���Ͻ����^`�p��=�1m=���X����{;};=}G�>,�H��=���� �<;,�<{R�<߿/>��>��Z?f��>排>�+:?��J�0�Ȑ��01?2�i=i��������M��P����=�4j?Ի�?�7]?���>�9T�.W�97>B�>mK`>�Bi>�&�>j��4 n�6l(=�>��/>�a�=���j��8�����IU=ty>���>��>ıx=|�k>pPe�D�2�_�>�f�M���1E�r�I�#�u�Z�$�@��>�qL?�^H?��>g���j��=�c��z�>��t?{Eq?��o?گl���߾��A�}K��'�h?:AL>y|�g��������15�J��=�8�>���S�~�e|k>������?�g���F��ݼ�_��=�X�Ά)=����Ǿ������=�'>p���>������KZB?!Z=h	��;@-��%��F�>�{�>OZ�>䩡�P(���?�$P���K�=��?y�>K^�<zW���^�bS�"��>�B?H=X?��}?OW��U8n��N�|�������Y�j�?m��>��?�29>�]�=`��\����b�PO�L�>���>*���v>�����2q���	��ـ>I#?<�>�i?=�W?06?&�]?��,?��?ٳ�>~�:�k䶾 �?S�z?��=����Ꜿta$���I�>�>w^Y?	���g�>'��>��$?�< ?��L?�V�>�0<>񠶾��5�oz�>��F>��S�F����=�A?�w?��m?"�?��<k��+�-���)>&[=_N;?�3??��?J��>Xi�>����*T�=�.�>3ud?U'�?��m?���=��?\�4>@�>=O�=l�>:�>0?�O?��s?`�K?�V�>'�<.n��<1����n�r_��T�;7&�<�=�r�O�o�`<*����<��I;_Q���?��}Ƽ!�C��:���^<�>���>�Ig�4>&���+y��PV>�*�]vJ�-��N*��{&>0i�>���>�_O>sJ���=a��>���>j� �E�?�?8#?7)>�8b�5��X#���#�>�b?�z�<�e�����n��0Q=�L~?�WV?c�p���	��b?U�]?�i�=�H�þ��b�V��Q�O?5�
?��G�ݳ>��~?��q?��>��e��-n�]��7Db��k�+�=fk�>`]���d��7�>ŝ7?�S�>'�b>��=ul۾�w�qd���?R��?j�?���?*>��n�+5���c��*3h?!b ?��z��?���=�5��Ws��Y4�:��[q�e�����p�kN��;
C��N�G�ֽ�˷=�E?_e? �n?��o?�s�y�a���_�=녿X)Z�t��\H�E�6�j�\�S�B�D�c�9t%��ZվZ��ޗ����z���G�蘵?�Q+?����:�>�}�����wľ��^>�e��\��`��=/4Z��;=G�/=��W�72,��Ш��L?&i�>�N�>EsA?$NV�f<��a0�7Z=�����>��>=��>v)�>�o�v+�[����п���	]u>�jc?u�K?�Lm?f���2�0�u�����"���&�����#>>�>N�>\�R�g���&�H�=�'�q�+��R��5-	�}�v=M/2?fo~>ጛ>��??�������n�m��.����<�?�>4 i?���>a܈>�#� �}�>�l?�;�>�P�>�>��i
!�Ej{���ͽۜ�>5z�>���>��p>�+��J\��`��99���X8�D�=t�h?8���+a����>��Q?c;@4<Y.�>s,v�K�!��o��*���>�=?o�=��9>�Qľn��?�{������_'? M?<�O��/��֗>��?G��>'o�>�}�?�r�>�پ�����!?or?�=?�D\?&g�>�y�=2=���L�R��a<)�>�P}>�y=3�(>�<���哾{������<��Լ�� ���~�V5�=�p�=R1c=呎<]2>�Կ�?����6������־�c3�|9]�� ����W�澟7���X�sC�;�6p���-���\�Ii�e/�?�Q�?��Q�پ�3��ڂ���۾�I�>S�ʼzS>�
�����=q��=�%�זm��N�a�/�,��k�e�5�'?ȶ��C�ǿ����>ܾ ?�E ?c�y?<��"���8�m� >��<�V�����P�����ο������^?(��>���]�>ʓ�>X�X>�9q>C���Ꞿ=��<e�?H-?���>J�r�1�ɿH����P�<���?�@ǏA?�a(�)�.JP=�	�>8	?�{A>`5.��"��~����>d��?�H�?�,D=j�W�@��Xe?��<��F�����=*�=W)=���w�L>]�>����lC�A߽e�1>o��>�#�T����[�ߏ�<kCY>a��9�0Մ?�z\�}f���/��T��V>��T?0+�>�7�=I�,?$7H�[}Ͽ+�\��*a?�0�?Ϧ�?��(?�ۿ�}ؚ>��ܾo�M?^D6?���>�d&��t�Y��=�2�����i���&V�G��=���>�>��,����O��G�����=���[ڿ~!(�"�㾡ӯ�/�
��ּ���.�K�9>B?彴튾&�|����<w�>�V�>�>NY@>�ڽ>��Q?�^d?�ѥ>�`	>j<ٽŝ��C�Q���=�Z$�ߕ��#���z`��|f�}����MȾ�/%�p������|���-�w�>�M������3�fd��, �4�>?ۑ�>Ljž�2_�}b��a%������=[���ɏ��g?��ߐY�T�?��?�__�ژ[������J���2��$�u?�)���휾ca#��Y=�ܼ��>���>g��>l���]A������U/?i�?�}��;���0	>yq轻e.=��(?�?d T�s��>rn?�'7�S��p�0>+t8>�c�>��>3�>�奄��b�?�P?�>��ُ�p>x><¾;�����=d1>=-�s���m�P>�錼�e���Ƽ
ݰ�\w�=ېC?E�<>V-�@���%|��ǖ=z۽].Q?��?#�>�K�?ڏ6?,�;�#���L���)	�>6�g?A�s?)�=4%"��qž0D��	�.?8\?S�.>Q�_V�g��eӾ��'?��Y?�@	?!Զ=�)e�S���ľ�18?��v?�n^��o��y��J�V��2�>\�>^��>��9��k�>b�>?��"��F��۹��lY4����?�@ϋ�?�;<���Ŕ�=�2?�T�>�O��1ƾ�]���{��=Fq=�>�����av�����E,��8?�?o��>|���ޫ��!�=�챾��?�֡?2�併~�Q�ɾ�䉿)���p�=�����y�=^A8� D��0fB�]8���Ծ����f�ؽ���>��@�����o	?�� ��������i�������+�	?Y�>5�_����`+R���}�3O��tA�n���i��>��>E�f�]$���p��<�,;���>�ͼ��>_�[�������������k>#��>�f�>FL��}ľ���?H���='˿�ĝ���N�L?C��?VЊ?�i?�#��,�W�aha�;�R�e�B?Əl?	n]?�9��M`��$���-Z?�����JI��$���:���x>=?y��>�u�K���$I�>_K
?I>2�)�lS��sV��w�ؾ��?�i�?���w�>t�?]�(?���r��%ݯ�"72��Q�=��C?��>�Ǿg��.���Dr?@E ?h����*�(�_?q�a���p�)�-���ƽ١>��0�lS\���y���Xe���&Jy�`��?RZ�?��?���#�0/%?��>�����2Ǿ$0�<Ku�>'�>F+N>�r_���u>���:�HJ	>��?�|�?�h?6�������9>�}?X��>X܄?��=ن�>%j�=�a���*"��n!>�I�=�=�	�?�M?�Y�>*�=֣:�w�.�֬E���P�G/�ED��s�>�Tb?!�L?�Gi>�����5�%`!�Ԛ˽�*�zj���@�4�(�佻f4>7�A>�>>sF�,�Ӿ��?Lp�8�ؿ�i��#p'��54?1��>�?����t�|���;_?Pz�>�6��+���%���B�`��?�G�?=�?��׾�R̼�>9�>�I�>D�Խ����Y�����7>0�B?[��D��t�o�y�>���?	�@�ծ?ji�h	?ח�oo���z������M����=?9?�����>Z��>>��=��s����Tt��}�>�@�?-��?�*�>�gn?��l��AI�t��<L9�>�f?E�?Q=����?.>�
?0�	�=���S�	f?��@M
@+�Z?����� ٿ�-�����|һ�>h�=�=wA����p=p��=�ҽ;�wI=�!>� W>�d�=�L�>�7m>b�6>�7@>c����(�_s�������=��������7*��]
�$"��\��������ž�9���*ƼK��< �H���_���{�f��=�HS?��X?Q�s?|?���y�'><���g(ּ���O�=��'>�y8?��A?��?+�E=h}����`�ײv�=����I���q�>�n>� ?���>�g�>�$���b>g<m>�+�>�m">4N�=)�w��]W���U>�>�m�>*�>�j�>x��=�=��+.���Q_�����H�z�)�?��ھ�5����R�M�
Ⱦ�>�J?6��>z����ƿ�l���S8?�d��),+�zR��>L,S?�z,?Pl�]0���T��06L>�%��Ꮎ�9M>�����mؽ�Q1�^�=�e?ڰ�>L��>�<1��07���e�D`�Gi9\G.?�쯾#R����I�)�s����>E$?�k���86������fz��;��-no<�d?}�?Kn��Y���/�����>T�=X�ռ@?�=��?�o����4�Ebv� 3>O�>C�;�* ?Q�,>���=ec�>^|��W��&�>�&=>�N>�h1?^�#?�V=n7Ͻ�)����{���>���> �>/0>DX1�U[=j��>�W>�י=p�
J��i�<����=6�=ݳ���g��q�<?s���@�=���=|D⽐�������~?���'䈿��e���lD?U+?g �=U�F<��"�E ���H��D�?r�@m�?��	��V�<�?�@�?��O��=}�>׫>�ξ�L��?��Ž7Ǣ�ɔ	�+)#�gS�?��?��/�Zʋ�@l�v6>�^%?�ӾPh�>{x��Z�������u�w�#=Q��>�8H?�V����O�f>��v
?�?�^�੤���ȿ4|v����>X�?���?h�m��A���@����>;��?�gY?toi>�g۾<`Z����>һ@?�R?�>�9�~�'���?�޶?֯�?{	�>v��?DE�?��'?���>͹n�+�ҿ����F�=�zB>���{��>���PJ��q��'���Xz5����v=�d����>��������>a�!>��ؾ!�q��H�>��?��=\�0>�Y*?�^!??h�>�Ȁ<Z���_�����G�K? ��?����n���<4ߛ=n�`�"?�E4?5�k�+9Ͼ|}�>�\?J��?S[?5)�>����)�������^��=��<�aK>/(�>ם�>=/��T�K>.�Ծ��A��?�>V9�>�嗼u�پ%���r�}��7�>�{!?��>IV�=�� ?8�#?8�j>�%�>yUE��7��I�E�m��>q��>L?��~?Y�?�˹�[3�e
���ࡿ�[��MN>��x?�[?���>����'�����H��I��咽R��?�dg?��}�?�-�?+y??��A? &f>�]���׾ ����Ԁ>q�8?�ֿ��Fa��Ig�"����*j?B?&R?i�|���৺��<���c��7X?�Bm?��9?����O���9��<~*	=�;�<+��=���Ӆ.>��>��/�r����B�<`�C>��Ⱦs<���ѼV>)ܼ�������o\>S',?sD�r���ͭ�=��r�W�D���>4WL>o���)�^?=�=�1�{�����x��zoT���?`��?�d�?3a��/�h��	=?D�?�?@�>���t޾�z��qw�r�x�u��>~��>j�5�*t������>E����Ž� +���> 9�>�B ?h?r>A�>�U���2$��>����վc���Ⱦ�e/�m,����N����6�c!�YԾ�m��٨>��-�h]�>�1	?�ƞ>��:>���>��=wݔ>-�>�ޤ>�c>��ǻ[�S>��>��L<�tϽ�IR?������'��辯����2B?;rd?�.�>��h�Ê��
��ց?ꅒ??p�?�*v>>h�}(+�r?7E�>B��rp
?r�:=з��/�<=]����M�����,��>XL׽� :�M�|if�h
?�2?����̾[Y׽����=:��?��=?բ�`+c��9q�ؒ`�ۮP��=x��,���g��T(�cPy�{9��D���a��%�'���:��'?׻�?�{ �����\���o���W��z�>�p�> d�>�D�>��m>�*ᾠ�8���W��a!�u���>�Zq?c�>�7N?#;?M�9?��M?0P�>�>h���� ?�u�WWN>$��>�"J?�KC?�?
�5?�_3?|-�>8@x<9G����ᾚA ?�w?�u?���>6�
?��c�=��Ja=��/��#��`L~����=��=%��<�2<-L=��G>�?�y�W�*�;f���~s>A'o?���>.�> kE���
���?�<=?5�>������� �h�Jht��D?^\�?3��(B�=�+�>Έ�={����;��>�j�<��X����,��}�B=�L>I�=�yY�5�(��j�ܣ��L}�<vE�>1�?�{>�ʅ>�����F��:���=�
v>��<>�]J>�־C������Li��cv>A�?��?f�=���=���=�v��+�����W���MƟ�~i�>a�?�3Q?���?��=?��!?�o�=l�g��++���ɘ��7?(�>?��>��Ӿ����,�������"?�?��t���A��5��x�"���1�>��'�prr�i7��-Q��Ng=kt��t�<���?)(�?+�Խk	"�ǂ
��.���,��(?��>V�c>��?�1 ���u���8�I�>:v?�`?ኵ>�9f?q�?�c_?d��>l�5�m�������r�>���>��?��?tb?�[�>�EA�� �צ��*� ���s�t���V����">�h>��>�J?9^p>K=U����9>�谽�I>��=��?K��>��>� �>�p��s:?���>�@׾ۡ�����-�`�"<�f?���?�h�>�ǐ>-m
��1�w��vY�>FK�?��?��.?��j��>�z��!Ѿc�Ž,��>��>ҙ�>:�<��5<O>J�?_ڭ>�NP����I_�!?$=��I?��Q?���>��ſ��q�f�p�����0i<����Nd��떽y�Z���=����B��������]�)8��呾 ҳ� 蚾��y����>���=f�=�]�=�ϻ<�.ټ���<2�Q=�&�<9�=Ln���<`�4�Ѧ�?h����ͺ��O<s�B=X�
��/˾��|?��I?�+?�D?r3w>�k>�H�A��>՝a��?k�X>jA����8B�<s��+���q�Ծ�YԾ��b�{���h	>�N�]>��->�%�=J��<���=�:�=��s=ZX���=ƾ�=��=�Ҳ=���=[&	>�
>x�w?m�}�F����EO���%67?�9�>���=w4˾��;?��/>�r���Z���	��$y?fM�? �?`&?i�z�j�>�X�������~�=�s��*�;>�u�=Z66����>��?>�;�P霿�i��xC�?�b@
I=?�%��E�ҿF�.>�	f>P�=UB���-�ub��_x��*�ҳ%?+E2�~뷾��j>k��=�h�FM׾.�<]%^>\Q�=���ܢ]�ͳ�=��j�V4���]=sP�>R�m>N�>[����.=��;Mb=c\$>�;���}�<�q<Wa;=?�*=�g�= ��=]�>ES?�eD?�s?S�?\{�ɤ����V<�>��f>�V�>���>WZ?7�>r�2?��6?hP?b(?ؼ�>S�>�	�>U;4�����1>;�53��Q�<ٶ�?R��?/#h=Rr���v�G35�sH	�T���u�>��?l�>	^>
���_���6�4��aX��i(7�l]��15~�2��u�>
��9�ѽ�w>�p:>���>.?+�>�8�>I�>���>�b�=W�z=b�L>���'L�A�ּ:=�{�;�P�=��@> +�==�,��{��v�ZD����;L�=�F�=e�>)>��>�y=9)��(�(>����<�C����=溲��]@��.d�3��_�%�R�7�j�@>��\>ᰑ������-�>�y>��7>v��?��w?�>D1񽚐ݾB��7�Z��N�e#�=6�	>Uc��/2���[�O���̾.��>�p�>�P�>o��>�S�u�+�� �=�uþ�zI�W��>C�g�k�Z��1���3��`��dv���:t���ӽ}95?���q��=�
�?�U?��?讜>�ҽ��*M>����b�>���D�)��M>�l�?:�*?@?^J��uJ�gc���Z��S��>RKJ�֏@�[Ր�E%��P�<+��9��>c���y~���D)�iф���?(4��!'��&�>!�>?#g�?�Q�������T���$��q�y�>)W{?�7�>�9�>���>�+��Û������>�+l?���?֡�?9=O=<=U=;��?EG?f!�?�n?7�r?]����>b߂>�@J>�����>�QV=b�L�J��=��?�v�>��>�吽�T�I��9�Ys���2^<��(>�X�>蜗>���>����>�כ��ri>~�|>@_�>�U>��k>��I>UU����S�5?A��>}0�>��?���>�#p�!�;_Op>���z��c&��D���p=C���=�	�;�}�;�HU�D%�>)տ���?Q>I��]e?�N�����x2d>_}�=G�����?����(�>�\�>�{>p�&>�W�>>�>>�GӾ�|>��od!��,C�I�R�9�Ѿ�z>�����&����Ez��5CI��l���e�nj�L-���:=�^н<�G�?q�����k�>�)�h����?QY�>�6?�׌�.
��n�>Y��>�>�N���vȍ�f�<�?���?�1c>��>4�W?ޗ?��1��&3�@rZ���u��!A��e�f�`��ލ�I�����
�z����_?s�x?�xA?u7�<-Az>���?�%��ُ�9(�>�/��#;��<=��>�*����`���Ӿкþ3��1F>�o?�"�?HT?	]V���o���'>6�:?5�1?htt?�^1?�I;?���o�$?|K6>@?d�?�45?��-?>�	?ǵ1>���=��e�mn+=j菽���tҽ��̽'-��7+=!�~=�wi;� �;�J=祌<ּ���߼ʜG;:Z��$�<k;=!��=�O�=�ܟ>�=W?���>���>:6?<+
�L\.��Ů�y�6?��=BP������݋�c��-��=� d?IN�?H4[?�<�>��H�^S���!>J��>0sS>�E>`��>ؽ}�k���=�g�=o��=?I�=�B�VL��
 ��e:��kDC�~>*��>��>��3K'>3��sՄ���]>�N��V��c3U���J�B1�R}���>8�N?�H?�6�=A�㾬V��<Ae�T�#?�A?ۺJ?I~�?��=�Pپ��4�q�K��!�%Ԡ>�̰<���䔠��٣�'3�<��e>����Gs��^�g>q=&�q+����n��]5�ꪾ0$�=[��e	>Ӧ�v�Ծ�Cl���-=�M}>y9���u�������7OJ?Ԕ<��޾A�4�l����s2>��>4]y>~N��W>�d;��?��i�q=}��>��4>��μ�.�=wQ�,j��>-:?��g?�a�?.fC�:H^���]�`���'���9ܼ'+?Q�>�x?��>+(�}��W�ӑU��Z���>��>%h�>�s�X�����6�"��_>~e?���>��?��:?a!?K�w?��6?5|?��>�����#?2^�?<�==�P
�h�9���C�O1��?��8?��ؽ:�H>��>؝?��?*�S?	�?]m�=��Ծ�a&�6��>Ox�>�8i�DU��;5Z>��T?���>4 @?�8?OF>A�N��c����Q=�><S~�=l�?�/?p��>NK>>)��>����y�=X��>Hc?�(�?��o?���=�?�V2>���> ֖=L��>�|�>�?uRO?��s?��J?Ǉ�>��<�V��3o����r���N�xc�;��K<�y=p��2]t�������<�|�;�s���v��T��<�D�Ͳ����;n��>Ynq>����#~2>I�þ�����@>���GF���싾�:���= >{�?y��>�%�[�=x�>�D�>��QM'?��?��?��;e�a���۾w�P���>�\B?��=��k�J����u���h=�tn?��]?O!T�����ʝb?z�]?6���e<�Zþifb�O�꾘�N?��
?�SG����>�?��q?���>��g��tn�A�����a�i9h�Sh�=�М>[y�1�e�|��>�6?���>��a>}�=�پJCw�a�����?8$�?�	�?��?�,->u!n�+h࿀jݾ�֦�op_?]�?�?x�xD?|���	Ҿ�
!�2����̾������ϑ�V��؛+��Ӑ����)XK>��?�l?>�n?�MH?�z�f{s���Q�P�~��}b����w �.�$�Q<�|�H�GtU���%�W�
�~���>��i��wa�x(�?CJ6?�0��&"?[=��Y��3�����>�ˎ����� �=)}v�F�6=��L=#�o�.M�)���w!?�ʩ>�?�>(�.?.O�&�D��$��3���ߺJ>�E`>�͜>���>�
y�ăܽ^�D�Ҿ�%���ܼ�Wv>vwc?�K?��n?k� ��1�������!���/��^���BC>�>���>'W�{���*&��N>�J�r�a���x����	�b�}=�2?@i�>���>�D�?%?�Y	��O����x�Vq1�
9�<��>Ri?L7�>��>y<н(� �L��>~�l?���>��>9����Z!��{�8�ʽ�%�>rޭ>���>��o>-�,�� \��j��]���W9��}�=`�h?탄�#�`���>,R?�f�:�H<�|�>9�v�Ļ!����T�'���>�{?1��={�;>�|žB%���{��8���1?��?�ݗ�t� �c�~>|�?���>��>�߀?J�>�]����?J?+�H?3?�-�>#�<�r��+%���pL�,>���՛>f�d>��=��T>�>3�h�?�@cn��$=�%�=L�Ѽ�	.=i!к� ��һQ�����=������D��pȾD��������/�x�û=6�饽���������"�������=��BT�l����p����?���?۾w��Ƞ�l��g2�������>?A弉ּ�b���T��^�.����������˾�9���K��Ti�S�'?�����ǿ氡��:ܾ-! ?�A ?5�y?��K�"���8��� >�D�<�*����뾯����οN�����^?g��>��.�����>٥�>�X>�Hq>����螾�.�<��? �-?��>�r�2�ɿp���@¤<���?-�@�rA?Y�(�	���oV=��>	�	?Q�?>�w1�B��ڰ�?Y�>�6�?D��?N=G�W���	�be?�<��F���޻L$�=��=�;=!����J>�Y�>0o��A�u�۽V�4>ǅ>"����r�^�3��<�]>��Խ�㔽4Մ?({\��f���/��T��U>��T? +�>8:�=��,?Z7H�a}Ͽ�\��*a?�0�?���?"�(?=ۿ��ؚ>��ܾ��M?cD6?���>�d&��t����=g6ἳ���z���&V����=_��>Z�>��,�ދ���O��I��T��=���B�ÿt��&��w<��z�ʼ�܊�{Ľ��N�z������Nfb�B.��t�=z]>`��>�d�>ߓT>#�h?l?�
�>��>ћQ�`+������]�<��J�٢��'�`�����T�ߪ��_�������׆	������h��s>E)C��t����:��_��Q
��g/?�U�>��H�u�4�w������.��E�=<wh��+)�[�꾨~Z�լ?&?:-����C�`^��V
>�;?=��J?�兾����<�侇��=�Y>ђ=I��>���<�0���W��O�OB1?�?�ߢ�7	��cO=F��~9>d]*?�/?2?�<��;>�?�i�����h�>���>P*�>�-�>2�=��ϾW
��Z?x,I?��W���q�1��>�╾F����c��	>T�=�UIԽ��T>|�ѽ��vX�w]�v�>'~V?č>�
)��l�,�;��P8=��x??�Р>��j?��A?*��<~��-R�
��y=_�W?��h?�	>�b{���Ѿr֧���5?�Ee?g!M>�h��Q�[�.����=�?Ruo?��?g̋�	�|���������>4?S�u?J]\�a*���2��[�ĺ�>��>Y��>�^7���>��=?�"�F^��F����~5��?�l@xO�?�"�<�+�Yi�=׋?�t�>��H���ľ䀷�4β���=#9�>Iߦ�#�w�����-'��O7?�V�?6��>Q���7��,@>ٶ��wD�?���?�����0>Gf+��y�~Ѿ��+�'�A>r�=w^��{��R 2�Á�˶U����B��>�A>?@�7��Je4>��z��Nڿ�߿�y���	������@?���>�O3�$'�a^��ϳ�o<�%,�p(P�0�>��=��׽�f��Q�{�a8/�}ډ��i�>x��н�>�o������T��P༇�>���>�@n>�����;�ƒ?��򾘊Ŀ����1���N?9��?eRy?�-?�H>b��-~�8�=�{=?� H?�ge?�?�=
љ��g}=�j?�_��\U`�َ4�fHE��U>�"3?�B�>K�-�ڱ|=�>���>g>�#/�{�Ŀ�ٶ�K���S��?��?�o�1��>i��?Ks+?�i�8���[����*��+��<A?�2>���4�!�&0=�KҒ���
?`~0?�z�k.�U�_?�a�<�p���-�c�ƽXۡ>��0��e\��I�����Xe����@y����?E^�?`�?ʵ�� #�`6%?�>R����8Ǿ	�<���>�(�>�)N>�H_�k�u>����:�i	>���?�~�?Jj?��������sU>��}?$�>��?�m�=�`�>b�=,��-�5l#>�=��>�\�?�M?�L�>�T�=?�8�}/��ZF�aGR��$��C���>.�a?I�L?�Hb>� ��#12��!�kxͽIb1�!H�sN@���,���߽Z%5>z�=>v>��D��	Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ta~����7�|��=��7?�0��z>���>��=�nv�߻��Y�s�ƹ�>�B�?�{�?��>�l?��o�L�B���1=5M�>˜k?�s?�Po���n�B>��?(������ L��f?�
@}u@^�^?$�hֿ����^N��Q�����=���=Ԇ2>��ٽ:_�=�7=��8�o=�� ��=p�>��d>#q>9(O>a;>�)>���O�!�r��[���O�C�������Z�D��Xv�[z��3�������?���3ýy���Q�2&�>?`�i~�=}U?�Q?��o?� ?��w���>Wi��(�=F#����=A�>��2?SBL?e�*?"�=�M���d��-���C���.���N�>	�G>6�>��>�ʭ>ς;�[I>�?>!�>��>� )=�v$�\�
=m]O>�s�>���>���>@�>�a&>桹����t�i���L������̝?A�Ǿ�����Z]���S��ر[<�D@?��=��w��qϿ9��G�E?3W���+�w�� ',>*o)?�#a?�Y=ݾX�8���=a1ʽX�i��>b�#[�g�'/�=�M�>�ƀ>�s�>87n�XI+�Z'F�N2廟�?��?FN,�.E���n~�o�`�Q�ƾ���P�-?ds#�u��M���A���������P?K��>�.L���������$� ���$>(��=�s]>��=�\>�⚽�ʢ�������<��u>k�3>(`�>��\>D��=�D>%����7���w�>��>a�>Ĳ9?�? ������姥� G:�k��>�{?1��>�Zy>��m�@�=�v�>14d>5�=PýVW(����Lp>H����`���RP�=����T�;>0��<��K�Y������;	�~?�~���㈿v��a��ClD?�+?��=��F<C�"�����H����?@�@�l�?V�	���V���?@�?��� ��=�~�> ٫>Sξ=�L���?F�Ž3ʢ���	��)#�DR�?�?K�/�mʋ�Gl�n2>�]%?;�ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾;`Z����>һ@?�R?�>�9�~�'���?�޶?֯�?�OJ>>�?�t?�q�>� l��.����t܌�9y=M2���>�W>�׾�4�D��G��tŉ��k� :�f�h>f=Yw�>�������w�=�E��'C��zo�w��>$x>��L>S֜>M�?�<�>���>8a=��u�A�~�F�����K?H��?���F-n�Ye�<K��=�^�Z(?vG4?�[���Ͼ�ʨ>��\?s��?�[?qb�>���Y;���㿿�z��m,�<z�K>7�>�A�>k��Y[K>��Ծ�3D�Z�>�͗>ƣ��4ھ�������7�>�]!?W��><��=��?~?a�>���>j�:��닿��O��5�>{��>O?\7�?��?~��_%��,���'����a�eEF>�9�?�?�c�>칌�h0���y�l_���ܽry?��c?��4�G�?L�?_]F?��J?v�l>9h�c����!��{�@>>:?��x��f�A)��(U�6� ?�,#?)7�>�ׂ�ԏU���o�;e'������(�>�f?J�?�� �Ħ~����@]=��?��Jf=>�V=A����W.>�B>:KE����=x��=�X�=u��^�b�<�FL=b��>2�>=4��r�T�T�?|	=�^,��M�;��c�{vG�z>��>ա%���_?���gMx�XT���3��千���??�?�<�?Dh�=Gh��R?Q!r?�](?�?�
����6h��� ؽ��;��:	�煕=�k�>�(>�d�!���� ��n5}�'�V��#���>K��>�?��?��A>	߬>�h���&��k��o)���;U������3��".�?S�v:����ԉм��ɾ򴁾�ē>Kbp���>z?]J>��Q>{s�>�2<�ơ>m\[>^e>�!�>�[M>^R>f��=Og'=8����KR?������'�Z�辷����2B?�qd?1�>�i�O�������?���?Zs�?>=v>�~h��,+��m?�=�>B���p
?M`:=��y6�<�U��"���1���!����>5E׽� :�M��lf�Ui
?�-?���p�̾�7׽���� �n=�N�?��(?��)�S�Q��o���W�]S���h�Q����$�I�p��a��'��/�(��?+=�~*?1�?W��=���'��"k��!?��Bf>2�>�2�>��>�uI>��	��1�Y ^��F'�ʪ��TV�>�M{?�>�>�#D?#AE?U?�m?p��>��F>&]��a=�>; 9�c�>��?�#H?�#?�Y!?5{
?�"*?�bJ>�V�� �$�ܾ8�?�`	?,?(��>�n�>6�d^�����rQ����,��y�}��w=�����<����=�|=>Ei?d���8�:���� k>B7?�}�>[�>��������c�<:��>��
?�>6����Hr�IB�S5�>!��?�)�&�=��(>j�=����g��ca�=:Pü�ڐ=��c(=��"<ߦ�=�%�=m�y�pC����:�i;�o�<���>q?��>q=e>�1���д����=eu>Nna>�`&>��־K�����X�m���>?d�?��?���=U��=��=$z��4䮾�<�?��0W�; �?�O&?`�Q?hЊ?c�?� ?��(>w�������}�q^���?=%-?��>j���T�쥕��'���?y�?BD\��3����2�5b̾�!z���Z>�(�3*��R���r�C����<�)*�R0"�#:�?�6�?��� 8�a,�城�# �A�?��>��>W��>4�gww���C�RJi>b��>�`_?GL�>DKK?��?��^?F�/?����u̾�7����l����=B�?!��?���?X�?�謽E���? ����!�������ܜ��pa���>=)q	?`s~>�E�>��>&=�=��,� bq��s���c�f���a��>�u�>�[�>�&>x��M8?"V�>�彾��.�"��4�5�Bs>�lf?U,_?�\?��=ݎ�B���⾮܍>��?���?��9?��F���=�+�=�k^�^�7���>:�>'G�>d=�>.φ��j�>��>% �xq�r�<�2C��!?Hy?��d>�ƿ;>n���q��.��<� ;ڀ����]�]���!Q��l�=6�������H����n�T���횎����Ź��F�z���?�΄=���=�I�=��<p��3��<W�U=��<�1=؞`��@�:�Ӽ-x�;��s�h�"9]<8�I=��
��ʾ�K}?OuI?��+?��D?��y>�Y>�7����>�����9?eZ>U�F��/����:�Gx���w���
ؾ�a־=�d��韾�j>��G�D�>�>3>�=���<| �=�Nj=,��= F޺w�=���=W�=��=�b�=�B>^�>�6w?6���ಝ��4Q�1[�O�:?�8�>�|�=Ԁƾz@?��>>�2������wb��-?j��?�T�?x�?si�Ld�>>���㎽Ls�=(����<2>���=��2����>��J>����J�����4�?��@W�??�ዿ��Ͽ1a/>A�1>�2>��R��0��؂�j�[�.4���?�{B�Gǭ�.�R>^߫=O�ľ�ɾ���=�4>�I�<hnZ��c���=��ν���<�΢��e>��1>���=?ۭ����=�'�=��=I�]>�|�<��޼����}�=��==^>��B>���>��?��/?��b?��>.�h�Ҿv�þ�ǋ>���=��>l��=j�N>k��>�5?�IC?��I?�Ю>�=���>"+�>�+���m�(�۾|���w��<�?�U�?���>Dy��k3=��X�Q`>��e���?�	5?9x?e�>�U����,Y&���.�A����r=��+=Jmr�PU�����Lm�V��*�=Bp�>m��>��>�Ty>l�9>��N>��>R�>73�<�p�=�茻�ĵ<s����=ޞ��� �<Pvż���b"&���+������ҍ;Z��;�]<���;���=���>K>���>|��=*���</>=���ҺL�xο=�;���&B�H3d�d@~���.�hK6�Q�B>�RX><���2����?�Y>=z?>���?�5u?�>�4���վ�J���#e�@@S�ĸ=u�>��<��p;��]`��M��|Ҿ��>?(>iV�>��>˽��=����=>����S�Jʷ=�����>N������B�&���H��a*;��d����;?&i��|#��)�r?�9?wl�?�&�>�Jl�u�=��B.>&ݼű>ʮ���;l�Ҧ/�z.?�E?u�	?��}�1�(��zξ;2����>�fK�[P��ڕ�L0�F��ꐶ�]�>������о��3�󯆿܏�ӯA�Ho��a�>�O?���?�ea�/1��L�N��z��V��_�?'g?&�>?�?�����g�~�/�=n?�B�?E��?�
>غ=W�Ľ,��>�)
?`��?C֑?��q?B��B�>�98��%>=����C�=f(>k�=z5�=�5?(q
?��
?b����
���ﾘ��3�]��4=�џ=���>j�>Ajr>�0�=�`=h�=-�Y>l�>B�>�`>�X�>���>�	��CB^��/?��>���>��f?[#E=b�<�,>==��/��>ԝ�"���n=�M����=)���k>i=>K_�>/�ÿ��[?4��>��_&f?h�Ծ�@<� ?G�>i����=���=��X>Z�>���>��1��ϣ>�>VFӾx>����d!��,C�-�R�<�Ѿ	~z>���3	&�՟��v��AI�qn���f�1j�<.��W<=�%��<�G�?P�����k�C�)������?�[�>�6?�ڌ�Y��̮>���>�Ǎ>}J��`���ȍ�9gᾅ�? ��?�;c>��> �W?��?$�1��3��uZ��u��&A�3e���`�_፿�����
�e��&�_?��x?\yA?�b�<�9z>��?�%�4ӏ�d*�>Z/��&;�{?<=`+�>�)����`���Ӿ��þT6� JF>ٕo?�$�?`X?VV�70F�Mz,>4=?x3?�{?�b0?��1?h�=�#?�m>�9?% ?u�7?��+?��	?͂,>AP�=��g���X=����چ��$�ƽ'g��D�ۼw�>=g�{=)ǅ<#�;��<C��<��f�%��뻬+��|<�"=��=k��=dԥ>�X?�B�>$e>��$?F7�Y;)��d���0?��=��g�{.������[� N�=Jp?!��?D�b?3U�>�UQ��K�zA>m��>��2>acQ>_��>"�ͽ�����=��>��=���=&���<�i��酊���u<�$/>J?&j�>m��gD->����7g���>�$�����,���4G��-��?D��8�>�@G?�/
?CB=.���5���i�R�?�5I?�T?��r?��W=�ѾĆ,��Y�d�p�Xf�>����		��X��Zw����W�{Z����\>��s�p��c\�>*�-����o� �3�b�x�#�9>���`-�=X9&��������hX==je>tY���=��!��Is��F�O?b!3=��'�yY����
��>�A�>�fz>M�g�r��=�7��Gi��E�>��>�޵>�=/���VT�)�O�>�AB?��`?!k�?;pO�lj���D��\�9z��5F���?�>�?�+p>3WU=>����/vT��{<�@n�>�'�>�]��\I�4۷�X2��M��eo�>���>o.>��?m3N?�?Ǌd?`�"?^|�>�Ȗ>���/����%?;(�?�=�н��R�c8��E�]-�>�*?�UH��ٗ>N�?�*?S�'?��P?��?�>�G�d�>�88�>���>��X�����;_>lfK?���>�?X?y8�?�8>� 4��%������`�=�;%>/�1?� ?t�?J0�>�?�����S�=�k�>�j?#��?��I?��a�� D?g�f;2; ?R�>�Ы>�!?%?�v?�k?�U?���>Rh�9�:7�4��O!<4rj�5��<�>�L�=�P>��o�B��
آ=�������<!6;� ����N�3t��=�(�>��s>X���+�0>"žn�����@>�k��F������BD:�%��=���>�?3��>�#�å�=�{�>��>s��(?��?�?��;vvb��ھ= K�F��>� B?��=A�l�&r��"�u�v~e=��m?�^?l�V����w�b?��]?FM�j=���þ	�b��v�H�O?��
?2H�Mֳ>%�~?�q?"��>�e�\n�����Qb�]�j��"�=x^�>*k�{�d��2�>�7?'i�>f�b>��=��۾�w��`���"?��?<�?��?Ԯ)>_�n��&࿸���pu���1^?u��>{z����"?�h���Ͼܰ��㒏�\������ت��v������7�$��J��X�ս��=��?�
s?b�p?�_?L �Ͳc��K^�����?V�p�����VE���D�jTC���n��5�����Rԙ��C=sQ���n� ��?b 3? �ĽU��>�Ӣ�O�D@��w?�=�����"��a>td�V��=�
�<(N�������j���?��>q��>�S?5|D�l25��g0��h=�;��3 q>��>	�>��>��ڽ�$�G�νx˾����A����s>�c?9�J?�gl?���2�0�&U�� ����.����=>�!>
h�>��N����#�1�>���s����Z_��6	��S=�m1?�o�>D��>�i�?i?=��s���"{��/�<��<�a�>�h?���>�f}>���|���D�>��k?u>�>d#�>�H������9u�6���K��>���>��>��[>�2E���R��H���p��\�8�J��=�@e?����a�b��x>Y�S?E�<��X<}��>-���g��O2��FL��C>�Y?s��=�P.>)����/��U�����"(?��?򑾥4*�R|z>_v ?z�>F�>X�?�>����H��}{?�-^?�RJ?-@A?�1�>.}=<���.�Ƚ��&��,.=��>�X>��n=��=���6m[��3�4�I=,�=Ԡȼ�ܺ��2<�����e<T*�<ŷ6>���d�q�,�۾���4l�V+�I=�����Tܸ����y��⾁Ժ����ܟ��j�s�H�;뜾\���f��?S��?�.������4_¿�}���ʼ�M?ǎu���5�Ȥ��*��������Ձ�7)<�(�_��l�Bڄ��e3?c�ɼpy��bG{�� ����N?K`2?�af?�<��_��}���=�0��z��{��됿�S�±���0�?���>�K��i,��k@�>
��>)!m�gT�>	-%�K�оm��=C�>�a?��?�rQ��ʽ�a>̿�m=�[�?_�@��@?r�!��"ݾ=��=���>�e?j=>&LW����Р���j�>��?�?|�q=@?^�VDk���a?U��<��A�7��:v��=�k=���<F��:>�U�>ԗ&���L��f��=�h>��~>m��=���~�)<;�>�}�����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�}��=[��>c�>,������O��I��U��={���ƿ}�$�/{��g=n~��9[�
�U�����S��#����o�t����g=<�=F�Q>(w�>��V>Z>�_W?��k?c+�>�.>U������;����i��)������p�,�p��߾͎	����G����ɾD�a��7b=�qJ��v���)E��tm��C&�[�4?��_=�����	M�k��?��.���:-=#ᇽ�:��q@3��Ou�HȜ?|D?'y��3�w��4�m�{=oT����L? {i�I�־q��SA�=��<�*�=8��>tkQ<_(��MY!��{L�7#?�&?�K�����=c(��=��'? ��>�;=<ʧ>�N?'�X��V׽j�B>Q�N>���>���>r��=���l�ҽ�?rGT?�R��7���/>T�ʾO�>�߱�����=�+�s�����>ar=�|���,��A��0"=h�V?���>��)�
��ː��3 ��(A=~�x?_t?t��>c*k?�B?�v�<	e����S�%�
�H�{=��W?��h?*�>9�����Ͼ0B����5?�Oe?h1N>��h�J�F�.�$�(�?��n?��?ؘ�C:}�X���	�J6?�pv?�^��3�������W���>�g�>[�>�9���>�N>?|�"�.~��G���KP4�L��?�@�|�?x�B<6G��"�=_�?A�>O�7ƾh���k9��hr=���>�7��S�u���A�+�k08?���?$��>J���O���.6>��?�Ƒ?���<�*�=��8�K�|�H�����|�n=H܇>��R>C	�$����4</�P�_�A�=�yS>3q@h��<�>�~=px��UֿV>���{��: +��=?0�>VJžW�y��&��+TZ�*����7�3ξxΘ>>�.���ᖾ�z���9��u��h��>�D���`�>��M�XA��F���Ҡ<��>_�>v��>�N������jU�?��i�ʿq���=�G�W?ڈ�?j|�?�?{��<�b�*��'��;��5?F%h?�:O?r�鼓�D��A'��8i?���Y5Z��B)��?��q>[�2?J��>)�-��=��=AZ�>"+9>^S)��Gſ ���w�D��?~��?E>�ch�>�Ġ?&\4?gq��>���r����0���H���I?��">-��'����1�5J���o?�5?���y��_?|�a���p�S�-���ƽZۡ>�0��e\�D�����:Xe�����@y����?^�?9�?'��f#�26%?��>>���&:Ǿ �<~��>*�>,N>�D_�n�u>��q�:��g	>`��?~�?�j?Ε������U>��}?�
�>�?���=7�>}��=a󰾙{,��k#>h��=� @�p�?P�M?6��>��=i�8��/��QF��:R����C���>��a?��L?��b>E޸���3�|!�/z̽J+2�9��I$@���,���޽R�4>E�=>�>>>�E�g�Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�L	?��H��-^~�����6����=5�7?)�{>���>�=�v������s�)��>A�?�z�?7��>�l?�to���B���1=�M�>;�k?fv?�6l����g�B>p�?6�������C�f?�
@�q@��^?8뢿uo꿜��⧪�#]���}>��=	>�Yǽ댄��_�=ˢ8�5�+���=L�P>��{>�J�>f@�>�%X>p�f>����ɴ�gb��C���{�[���"��cھc���K�Q��K;�n����X7���%ݽk������lH���Ň����=q�Q?�P?��m?Ֆ�>����C>�����@=�P�5�=(��>��1?�L?5�)?��='��Fyb����ܧ�G�����>�rJ>�@�>���>5ί>e�q<�tN>2�C>a[�>��=��6=���=�R>�>�N�>�ؿ>�~�=�-A>�9���%��D�Q�:R7�|�>&��?���Q4�:���)�Ӿ�+\���0=U?�.>=���LԿ����B?:�l�Yt�����C�>�nN?\�Y?��G>��⾎���=��k�u�:������x�==͈�#5�*��=4N?�C<%An>L�p���i�"�&��D7>-��>�88?�����->$|���f��V���t۽�G;?�AK�.����Ε��	���G��D<2`S?�`�>H�B�K�վ�����TN��{�>p�g=ڮ�>�R,>0�8>�m=�$��0
��>7�l>��~>�]�>Ȳ�>Pf.>q!�<�Y��� �>�0�>�R�=T�[?��>������ܺ���ƕ����>~�!?8��>=��=�-����=6��>� >���=' @=O�v�H#q��b�>�	j��:�}�����k�+�=@�&>5�ݼ5��T3����=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾQh�>wx��Z�������u���#=S��>�8H?�V����O�f>��v
?�?�^�ߩ����ȿ6|v����>X�?���?g�m��A���@����>:��?�gY?voi>�g۾;`Z����>ѻ@?�R?�>�9���'���?�޶?֯�?d�q>���?{w?�+�>\}�=~.�Z����i���8>W^��8�>;4�>���+d ������`���R������$l>=�=��>hsR�s-þe��<�� ���̾�]����>���>���>��>M��>�J�>E>�="d]��K�=DK̽����K?���?.���2n��N�<e��=�^��&?�I4?k[���Ͼ�ը>�\?i?�[?d�>;��P>��E迿4~��H��<��K>(4�>�H�>�$���FK>��Ծ�4D�[p�>�ϗ>�����?ھ�,��YR��EB�>�e!?���>�Ү=T� ?T�#?=�z>��>�:�Bg���M�'@�>��>�?_��?��?�x��R�,��o���r��B�U���V>�Vu?݆?'b�>�P��Ey���oͼ�ڀ� δ���}?$�`?/^���w?�ą?��>?�sC?�II>>���þ�EY��Uq>H?;���yS�}�-��I��1?�?��>�T�;MZ�E����'�Gn���B�>AVg?�?����'m�?�ؾ��<��/�|;�O��R��<]u/>t�>�����`>��=�w�=�Z�EFC��#�{]�=�B~>^�>"��&�5��*?p������X�=�Ls���D����>%DP>�����Q_?
^;��z�/���w��a�Y��x�?S<�?`0�?<����g��;?> �?��?�6�>�4��\7��X�Ɔn��es��X�/m>�z�>%�j�*\�!㣿`G��a`��b��������>a��>"1?��>]�B>A��>�V��"��F!�����[�����W3��,����Ti��<)��s��r���z�Վ>?@i����>,?b>�o>���>�Z�P}>��U>D�}>�ݪ>�PW>�7>���=�������KR?+���Y�'�>��񰰾63B?qd?#0�>�i�|���?��{�?I��?Rs�?<v>�~h�-+�ln?_>�>���rp
?�Q:=� ��>�<�T����.��>�;��>CC׽� :��M��of�bj
?�/?h���̾t8׽]D���x=�_�?OT)?=A(�;Q���p�x�X�<�Q��6 ��c��6���$�Ԛo�`>��+m���ƃ�Z�'�5�-=Y*?츈?��L��j?����j�@�?�EEc>�v�>~(�>���>�iH>�	�X�0��_���'��"����>2Gz?��>�,?p�5?�z[?ayV?P��>8��=@�侔$?YL�b.�>Ji�>�w6?��??ε?P�5?�5?)�>Eн�g��mþF��>W$�>�@?(�"?�7#?_b齷G=�c_����?���������,= ͐=�M��.4�=N#�>�V?Ȓ�e�8�������j>�7?��>���>$��N*��U��<N	�>��
?�B�>  ��zr�<a��T�>���?�����=��)>'��=�p��0�Һ?Z�=������=i�����;���<`�=���=��s�p�u�wb�:$�;wn�<��>;?���>NP>�렾�����&>AF>���>��>	ξ1�������e�+1�>o�?��?>	=Nu>� 	>_���h,��Z���	D���HF=iw�>7�?�WB?���?�'?j5*?);>>	�	�~Ɉ�7o{� 㯾�)	?�0?V��>)��Ug�����nLA��A?|�?<']��5��j#��k�ؽ�=���=	�B��]���)���h�$ �>e��%�޽���?��?/�Ľ�yo��*�'��>D����X?u>->dg�>l6?�:��;|�aG�qE�>�|�>��E?;E!?��>�`?+�r?J ?)�5�ܐ���Y����>�u�=or�?З?ac|?#��?C&Ͻ�K=���<�,=�j����<�s%�ʜ�@�=|T�=��`>d� ?���>��=5&��r�m\޾�>>�z>�?:4&?r�>���=�y)�D</?I�>𜯾?�m`о����?$�<xz?\z?�7?_v=q�W�9�S����>͜?�W�?-i?�R��>��
������_��R�>b��>{��>���=S���$o+>�w�>"��>���rM��PF��ũ�yh?T�C?_�=>/ſ!ho�ʜo�XÙ�՜;[��%�`�ӆ��9V��~�=������G~����\�O�y��^Բ�M����|�J��>rl�=Y��=��=Lث<"�����<��y=�D#< �&=�|b�?�<e�3���g녽�kR�6�<�}R=�I����˾�t}?�"I?Bn+?�C?ey>)5>ȧ2����>�5��^2?��U>'wO��c����:��o��������ؾBv׾��c�K����]>�I� e><3>�W�=9��<c�=FCt=<c�=:ub��u=���=���=�q�=K��=��>�>�6w?6���򲝿�4Q��[�x�:?9�>&|�=l�ƾ�@?\�>>�2������|b��-?s��?�T�?A�?ti��d�>���㎽Tq�=B����=2>%��=��2�P��>�J>x��K������4�?��@}�??�ዿ��Ͽ�`/>z�=?�>�8�o6�uѾ|\���D�<�??�:�I命?x,>�a�QǾ�,��@�=z�n>�˄>G�뽬B��=�,���!�=�x�=��Q>�>�>6� �;��<��<A��=CY><O���M��c�T�=��/>���>��">x�>ι?4?!�h?��>��[�ݾ�Ѿ4��>��=��>�>�F>�g�>�+(?}UF?8H?}b�>Z�{=�>���>=�*�*)n��*�[��cG=�P�?�?�z�>�
q<��,�x��U�*����Ӌ?�a(?9	?�ۖ>�S����V&���.�u���*���+=�Zr�U�;����g�8���$�=�m�>T �>^�>PWy>��9>(�N>X�>m�>,U�<�l�=A̎����<����<��=���'��< ż8F���0%�q�+��O�����;Hˉ;�W^<��;���=��>��&>��>��9=6���o�.>Z���?���=Vᙾ9�>�
�c��^p���%����+/>��J>D�i�,3��K��>�h\>dRu><��?am?U5�=-�%��յ�oŢ�Mц���?��,�=0�>&�C�m�5��Jk��4X�`쳾8��>�<�>ܧ�>�S�>�,�)q���=Kپ�D�M֦>�����q�=PZۼ��7�uƤ�B>��x�m��_�35r?�C��y:=��?��?���?Y�?]Ƹ�2<���$>�]��I�&>ۉ��~ǾEt�<a'?M]?Js�>�q�`����>̾�྽�>m=I���O������0�;���ķ����>䪾��о�"3��c�����,�B��r�C��>k�O?��?32b�QR��nNO�������j?�sg?x��>�N?�F?�.��9x�/s����=�n?��?3;�?)�
>(?�=�̟��1�>�)
?>��?@O�?%�h?��B��>\	���D*>XS8���=�4>�l=^U�=2e�>��?2�?\E�������6��de���=�<��>RA�>Q
�>(��=��F=���=&~L>0�><��>�i>���>�>���J�-�rs9?G�S>��>X-6?Y`>�g�<I�=�y��0���-�*M�<���<q�����9*�"H>�3+>�|�>udؿqߑ?�6�>�x
����>���������=�3�>*>A���?J2�>�gѽ�m�>�'�>YsM>/�>sy�>/t̾r�>$!�����'A���J�Bʾrz>�i���M=��r�'3�
EI��Ѵ�cn �ӽf��9���?��=���?�L���$m�B<&��f콓�?5��>�7?,��ֿ���>y��>�>���������l��s��?aW�?�c> �>N�W?��?0�1�3�bZ���u��A�b�d��`�ۍ������
�96����_?�x?��A?�<�,z>/��?�%��͏��+�>i/�;��w<=�*�>�+���`���Ӿ5�þ�(��.F>(�o?��?�J?�OV�If�=ğ�=2�H?�Z?+x�?')?��>�v���
A?���=�/?O�?��(?>C?xڨ>�[�>~iX>6�G=��b<�Ͻu����f�Ze>��C���=M=���=���=o)==�2�ZϽ�L�=Հ��$ͤ��E;�F�?9�=��2>�[>�)�>�dS?���>�X>�X?���d(�#s����#?�>�|�������׾� ����=�*c?:��?Lee?n*q>��;���4���	>�1p>x/>�uX>
ڮ>S���^)��:4=%f�=ƣ!>�|=P$>�ss��?��>�����<r�)>��>�|>Ҡ����%>�C���5{�&3e>ەO�����MR��SG���1���u����>�K?��?k��=�;ɖ�4�e���(?�<?�M?1S?��=B۾)_9���J�J���z�> �<���/��������:�iq�:��s>�s���KS�g��>� ��*��yl� N�J�)��w6>��ľ��f��k3���$�;���=���>��پ�����wʕ��(O?�[���!��Y=�An2�>ǯ>�~>k�>�	��N�L=��5�Y�پD�U>���>I|>`s���TPA�hWþX}>�SE?��I?9[`?���2�|��GI�C� �r���[�kC?ԟ�>m��>l�>j�
>C����f�7R��]K�b�>)��>Fi�y�<��8Ӿ�о�X1��.�>B�>�*�>�0?�E?S	&?�p?�-(?��>���>�~�X�޾�d"?Vv?���<��ֆ��!C��3����>-?�͊�ډe>�%�>��(?e~?"WL?�*?^�>W^���J��>(KT>��X�ِ��� >��9?P��>��I?;-h?��>�="�J��/D�䱫<�ʕ=��6?��>?��?��>��>Bi��/t�= S�>"�b?��?��o?��=��?y�2>>��>���=9�>��>��?PNO?��s?��J?�z�>�ʍ<�������s��9P�b܊;
bD<��y=X����u���9��<'\�;���&�����(�D�����Έ�;Ȓ�>�s>tH����1>�mľ ��w*@>�&��:כ�{���iM:��=c�>�?��>ɫ$���=	ż>���>���6�'?��?
?��;�b��EھŵM�5��>A�A?�8�=vol��x��;�u�i6h=i�m?�e^?	2W�57��^�b?��]?�����<�9�þ*�a�9��Y�O?z�
?M�H�!ҳ>�~?��q?���><e�V7n�����(b��j��>�=V�>"_�|�d����>?�7?���>�d>���=\2۾��w�S���a"?��?B�?:Ɗ?2)>��n���߿1����^����Z?�M�>(���&?�/+���Ծ
T��D*��[�پ����?o���.��;_�����7ʀ�*�н��=:�?Zu?��q?.�Y?9��qye���]���|�`sT�`~�R����G�GE��A�Z=k�}��5������J��<�UK�.�F�`�?��G?�Yg�b?�>`<��1m��`���}>/8���C���w>4�'�A=	��<mhn�(�ӽnzZ�g�?�Ǐ>���>=�R?�A�S�?��;�r�5����̢x>48�>ʄ>���>C��km�I�ȽTǳ�l�x��;罜v>@�b?�eK?h-m?9����)1�('���y!���32���??>�>�	�>�7P����	p&���>�iq�In�w���Β	�c�z=�0?S~>��>�?�`?��	�2���Tvr��i0�tM�<�X�>gTh??0�># �>Q�ɽ�p!����>v,l?'�>r��>�_�����{�Q�ͽ���>�y�>���>7�w>`	/��Z�\Y��o5��qH8���=D g?�����b���>��P?,|�:��<���>�q���"� v�")���	>�?���=��;>��žQ���s{�L��(?+�?)���+���q>�?v_�>��>�e�?�u�>žʖ�<L?X�Z?=�J?Qt>?2�>�q�<D�ͽw����B#�A�3=�I�>��`>�l=��=�@�S�H�&��1;=���=������  <����.~<�<@�9>%�п�:����Ww�ls˾qSʾ���&_T�V��7ɸ�o<c������h��$.��g �н�p�b�Ԫ���m����?Q�?GV�e�	�Ǳ��%g��P-�
x?|�۽����`��Pо��[�����[���:��kP�*Y}�������;?񶀾ਿ�鉿~��O?	��>o��?�,��	�sB-��0�=(��BT�=ƾ0(��ſrc���f?�%�>j�ᾟvq���>���>���=�a�>��p�ʌ��?fZ=R�?�`0?��?�!K��rԿm�������8H�?w@�~A?��(�쾹VW=��>�	?�>>Tu0���!��(�>-�?j��?�P=��W�����6e?jS<�F�(�ϻU��=��=��=n�SpK>q��>�����A���۽�
4>歅>�����jA^�m��<��\>B�ֽT��5Մ?+{\��f���/��T��U>��T?�*�>R:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?:ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=q6�ى��{���&V�y��=Z��>b�>Â,������O��I��V��=����Կ
M5���Ѿ-7D>4Ʈ>�?�=�̩�^��f�#�$��>��9;�޾����ԍ��v�9?���>�l�>�;�>7�4?�wS?+�>�.������t�<F]H��W��*O��U$���0������;R:�3a�jC���������¾Ӣ<����=�qB�t���NE,��%]��B�W
"?�>�Uľ�WC��m��9澔-��Q���5U��V�̾~9��%o�jқ?�K?Lpx��_�ͮ3�쫽�����b?�(�������jǾN��=a��=���=X�>�Ӯ=��̾��'�zfH��B-?f�)?`탾M���襍= sD����=�	7?	Q+?R$�=@��>�2?��7aR���>Sk>u5�>���>/�=N���/'����?�:T?�Xn=0�k��d�=b5�
�-�=�ͽZ>7\��IxJ��6�>�=>f�������»�`;�U?���>"���������0�f�%f<��t?'?P��>�f?2�D?�]�<)��K'I�(���v=\S?��a?2H>!m���VϾ\;����.?�;n?�0>aX;�$0��{�)�F?�a�?�xl?X?��~��?}�L���H��ڋ5?�"g?�Ze�y������G���>|��>$�>�>@���>�?H?z!�d���cּ���<�#�?I�@�w�?T�=m��i�=��>r�>��5�z���ڙ�����Uym=���>���8�q�s��Z�:���=?{�?!��>o؁�m��y�*>'���a�?ݨ�?�nC=,#�A�G��؄��y��l g=��>}m+>��d=?�׾K�$��ݾ�
�BA���>�-U>J�@%$���>/J|��X俎G�(����R��s��S�?k?�:�}6X�N�h�R�}���T�}�N��b̾�>�>@l>XxW�����v�,
1��J���>���[ x>	MQ�_������n+=nj�>��>�j�>�s���+����?������˿QW������{^?h��?���?3?��<(����ֈ�#�;��E?�Fq?:P?�q�B�|�����m?�o���&S���'�2�;��Bo>(?`��>�}-�w,="�>��>w~>>8�"�2~ĿUW���K�|��?R�?:R�~��>�j�?�4?߃��6���餾��4�S{=HC6?3{->�����-�=9�cޞ���?ީ)?6ʽ0�ٸ_?2�a���p��-���ƽ��>1�0��G\��}�����Ue�j���.3y�U��?�[�?�?A��� #�M4%?��>X����?Ǿ,��<��><6�>i+N>��^��u>��q�:�B	>���?z�?�h?��������q5>��}?Eo�>&�?�/�=e��>x��=�����5��U">�D�=�H��Y?�M?��>c`�=��:��{/�}�F���Q�[�<�C����>f�a?�8L?s�b>�z���g.�)�!��Jɽ�3�"����>�Z$5�7�߽`.5>��>>n#>�KD�Q�Ӿ��>��>��ѿ���*t#�x+?�y�>L��>���p����$>�Y\?�~->w��S����f��A�Hϧ?p��?2|?�`ξ�����Q>�U�>�2�>���ܽ5鴾RN>�\?,G>�M����r��>iu�?
��?���?��c�f��>�������F�l�Er���m�L>�(?��&�?>��?���=\�v��ˡ��o��О�>�a�?�?6��>~|d?��`���7�`�=M�>w�r?��?oN������Fp>��
?Gj�kB��V����]?�@C@�(l?%���8ԿTZ����þc�s�f�0=\佉��=��8��N>�.��{+=��=���=>��>Qh>$y�>�N>q��>��S>�ӂ�#�E���7֕�]�M���.���'��Ѿ@�,�j��������{<u`#�p�B>��2��Æ�Z/;{�=4�U?֮Q?�]o?B ?����K:>P����=��"�ǵ�=6�>/72?>�L?�*?:%�=�ʝ�b�d��k��������a��>�H>���>�0�>&߭>�;c}G>�CA>���>1 >U\2=�ԃ��7=_&O>-��>��>�b�>��@>9,A>jj��p���sh��Q��b ��T�?闡���/������V���`�*�%>O�;?��=���L>п�ث��}J?>����+��Vp���%>�,?&;k?ʋ>;����<E��=��ƭm�1>��(�`rT�Z�J>�?�W>Y�>��4�2�1�[�6��U˾��>E�?8�I������߂��k��9��`�����>��t��/��Ҍ�4�p��Vs����=X(;?
��>����C�ξ�LӾ�g���>�)�=e�>ď�>�!�>������E]2�T�z=���>HyK>��?	m�>�>�P�=��־
?l�9��>48�>��=�R?WC"?yWs��y�:��(d9�d�>��O?���>�_�=u��C�=�9�>�|l>GV`��a�<m	��F!��8}>��2�'�_�H��.�<b ��x�=�=\���d�t����=�~?�}���ሿ���Q���oD?(?s �=ؔE<Ȃ"�E����F����?��@/j�?�	�p�V���?�A�?���N��=��>7߫>ξ�L�
�?�ƽe�����	�@#�vT�?��?C�/�̋��l��3>�b%?x�Ӿdh�>ux�zZ�������u�ָ#=;��>�8H?�V���O�e>��v
?�?�^�ک����ȿ5|v����>V�?���?_�m��A���@����>-��?�gY?^oi>�g۾.`Z����>ջ@?�R?�>�9���'�|�?�޶?گ�?�I>�}�?,�s?�D�>�v��f/���⌌��8�=Z ;�#�>4�>���;F�}���r[����j�c��$ja>>#=�̸>�<㽞)���v�=Q_��|����d��L�>|dq>��J>�m�>v� ?���>>ę>=uJ��Tu��o����H?�K�?ۡ��m���<���=�u2�S��>�&?r=$��˄�>hla?fyu?B0^?B�>P��*-��о��:����<32>=��>��>�ܒ�P _>R*˾�9'���v>۰�>��S���ᾛ�|�Ű.<%9�>�/?O��>X"�=� ?r�#?ܻj>l)�>�VE�F.����E���>��>�3?��~?d?�ƹ�H3������䡿��[��8N>.�x?�X?Y��>1����|��Z-F��G��;��)��?�Sg?CC�_�?h'�?�??I�A??f>w���ؾu:��6��>�?�ܱ=�i�Q�'�i�B��q�>�-?��>� o�un>1ݾ�-�Q�����>1�l?^��>��
�-����< �K�[=�N{��ӽ�8�=���=���=�Ϊ>�h<���u=#��=�M�<{���Ǖ��6����=�:�=�RY>�ގ����<�=,?B*C�Z�Rt�=��r�|oD�)�>�L>H����^?�9=�O�{�����y��B�T����?v��?�f�?"���ʎh�=?�?F?�!�>09���{޾Óྋ�v�ݝx�Yq���>���>'k���φ��3���0>����ŽF��ц�>�F�>L?��	?G�3>���>�ƾ<��2�d��3n9�j5%�b%,���1�(�"�, ɾ	��y�:�pо�?m���{>R⳽���>�	?�@\>L�Q>!7�>�5n�&D�>Aj>ͷQ>�$�>=d> "q>Mi�=�=k����S?�}���E �"Q�B��GJ?rzW?P�>@m�����xw��?�y�?67�?h��>]�j���+��~�>><�>��g���?Z=�<dsI���=Z������?5�~,���y�>���>�tN�Yg�n�?��?�)��Ѿҍ�� ��� �n=�M�?=�(?��)���Q�M�o�Y�W��S����b6h�k����$���p��쏿�^���$��ס(��n*=��*?n�?l��A���#���&k�Y?��ff>��>�#�>�޾>osI>�	�_�1��^��L'�=����Q�>�Z{?
��>U�H?�>?ƘC?h�@?��|>n�>𒛾�?E�o�1��>�s�>�g$?N�%?.?	"?z�#?���>O2���P��۾]�?�??�p?ڼ?p�>9��A3+�RDӽ�����B�^G�wP	>� z<�Q2�Hl���<%v:>��?-���7�I���<�k>�8?� �>��>���=��1r�<��>u�	?(��>����r�������>#r�?�D �g��<�-(>Aw�=�<`�fm�m�=6B��;P�=��n�;U3��<&\�=���=4R������:+��;���<���>%?��>k�>�A��V ���j�=�PW>h�T>͙>E�ؾ�'��
���)�g�;�y>:�?�;�?�uf=�X�=\q�=�(���ѽ�-��h��<O�?-#?�*S?ّ?�=?i#?��>�h��㒿�������?�9?!g�>���M������Lz�8��>;�?�xg���&����z٤���~IO>+"8�4��������=-�M�>����q��I�?�S�?�D���E�W�۾�_����;��-?��>#�>��?��9|����)� >�G?K"]?8k�>�HN?C��?<�{?��>��(����~��<>]�伃�F?�Е?�Q�?Te�?]�>0ǚ=����X���K�ξlOP���O�~�N�LwB>@�M>�#�>�{�>?��>�/�=��<H�;\��cY>t~�=T��>��>���>�%a>���=~�@?���>�~���\��<�U���{d/>8�?�_?��n?()�=����T��Pپ��>�Ŏ?�N�? �8?�b~���=�a=���4��È>��>Q��>T��>��=|�>� ?�g�>S�P�5�	�����<T�E?�J?�Ճ>�ƿ#r��9r��2��� Z<
���Ђc�t旽_�\�Ģ=$��������At[�1��������������.<y�CG�>1��=@��=6n�=���<p`��n��<wC=_ׅ<?�=��s���_<��6��l���r��F<�M=�X񻅉˾ӏ}?�;I?��+?K�C?�y>:>��3���>
����@?�V>/�P�k�����;�����~ ����ؾ�w׾/�c�;ʟ��H>e^I���>�:3>ID�=R�<��=Zs=���=�Q�=�&�=1P�=(e�=���=^�>U>�6w?W�������4Q��Z罤�:?�8�>q{�=��ƾq@?�>>�2������{b��-?���?�T�?>�??ti��d�>L���㎽�q�=C����=2>r��=w�2�X��>��J>���K��=����4�?��@��??�ዿϢϿ5a/>w�P>W#>��L��q1�v��d:���1��m?KV7�-d��]�?>:�6=�����趾�i�=|51>&�T=�-��=a�yk�=]~����	�|��<&�c>$<>6�$>0����e�=��=\2�=��H>)�<����c���SK�=3�O>�z>�>>
�>5�?�6.?�Va?9��>֝t�(�̾7���x�>ִ�=yc�>s�=<iI>��>pc7?�>C?� K?T��>�p=��>��>5,�Gm�B��k���2�<��?�х?���>��x<c�?�V)�Ŧ=�L6̽Ŗ?��3?"�?>�>�����B�'�h� �1�*Yd�`���|��8�=L�T�vj
�𗓽��=z�>4�>���>�z>� F>dp>�5�>rj�={���(��@�<�[�="��Q��=�PL�`������<\��<e�!���J��`��ͺ=�h�=�>ٻ\��=�=��>2�>��>.�=-��H/>�ꖾ�L�0Q�=ES��EB� >d�K9~�
/��6��7B>�)X>����1����?�Y>?>���?4+u?E�>d��M�վ=R����d��%S�o�=�>��<�@Y;� V`���M�ݟҾmd�>k��>�O?Z�>L�׾�P�ʟػ����ľUtD= 䉾MV�>�'�4=3�f��9`���|�E�=�)b?����-� >�b??�ك?�M+>�}�=(Y��]�>K�羬젽�W¾���h�	���??/?Ϩ�>k�Ѿ�Ws��H̾/���ط>GI���O�����y�0�s~��̷����>������о�"3�xe�����ǉB�@r�i�>��O?��?-4b�V���TO����V���r?�|g?Q�>�J?�B?�"��Dw��q���c�=��n?���?�<�?`
>\ۨ=Óɽ�{�>�j	?�Y�?��?Djr?��E����>��tQ.>����B�=�j>ѩ{=��=��?��?�|?����fj�*����/9W� �=�~�=�2�>}��>�/x>���=bJX=7�=�&U>G��>�ΐ>wya>�ʢ>�Ɉ>��$��x9B?���>H��>S�?448>���s��=Pe��6s��0���<�%m=����F�Xt��:8>R�>���>�A̿f��?�;�>g|��� ?��߾LC�}�i��3�>
t�g�j>f/i>�=�Z�>�A�>aт>GUj>t7r>���@>�����<��u5���*�(྘(�>�*���}D�:
����
�Z�֊���I�Pr��I����@�v�g=��?��i�E�!��%����?�j�>}2?~Ǣ���@��>|U�>�;e>����(&��㌌�`B�8^�?�K�?k;c>��>2�W?�?b�1�m3��uZ��u�R(A�e�F�`��፿����
�d���_?��x?yA?�O�<@:z>P��?��%�|ӏ�:)�>�/�';��A<=�+�>*��Z�`�D�Ӿ�þ�7�VIF>��o?3%�?rY?TV���m��'>��:?ʛ1?yOt?~�1?e�;?���-�$?m3>pF?r?�M5?��.?	�
?Z2>�	�={˧��'=�3��������ѽ�yʽ2����3=�P{= ~¸;�
<q�=�<���ټx	;�����<�:=��=��=�1�>ea]?��>6|>�0?'���1�3���~G/?�eN=C�r�nׅ�H᡾���_� >}�e?�? IZ?�@^>�>���A���>�ƍ>��%>ڜg>���>�����A�ר6=h�>�!>��=i%4��L{�L�	�	͖�x�A<O>���>�|>��.a'>)F��7�z��'e>��Q������+T���G���1��#w����>}�K?�?�=\l�Lߖ�~?f��)?��<?�M?U�?��=x\ܾF�9��J����q�>���<������r����:����:FGt>�����t�o�j>i��'�ݾ�n\��w��2 ��6>{v��iz�X�������<����.�=n܈>�ḾF���]��9����R?cY�'	��y��93��9�>;(�>���>�H�����=	�Q�!$ �2�4>޹>�~->�Y��\ѾR\�&D��3�>s�E?g�`?o��?�Hs���t�O�F����3	����Ѽ�>?cа>:|?$m?>$��=�ޱ�����a���D����>Q%�> X��H�N������F$����>U}?�)>�5?�T?)}?�}b?�D)?�n?2��>X󓽒z��+6&?�l�?�e�=A�Խa�T�ܐ8���E���>m@)?k6B�Z#�>�?;�?��&?lgQ?2}?o�>�� ��[@��Ǖ>m�>��W�=;����_>��J?�\�>�Y?D��?o!?>x�5����b^��B.�=n�>*�2?tO#?b�?v��>Ӫ�>�������=��>1c?j1�?��o?ƌ�=��?�I2>���>~�=���>-��>~?�WO?��s?s�J?���>P��<W1���G���gs��P��4�;�$I<��y=F���t�[���<���;����5���@�h�D��r��|�;sg�>��s>���X�0>V�ľ� ��"A>�)��P��l�����:�l\�=㏀>��?P��>#�� �=���>��>���1(?��?��?��;T�b�&�ھ�K���>~B?���=G�l��w��m�u���g=��m?�^?[
W�(��.�b?��]?@h�=��þ�b�e��Y�O?��
?��G��>��~?]�q?s��>��e��9n����Db���j�fҶ=r�>DX��d�^?�>��7?�O�>��b>�#�=t۾!�w��q��R?�?��?���?�,*>%�n�*4࿛��h��U`?��>@���E"?6��}�Ҿ_3��[�L��P���)������Y��^'���|�ލ��H��=��?ls?�l?��]?=� �H�f��HZ�Q{�]'Z���������"G�W�E��G�>n��T�3��$O��dI=�+S��s^�u�?D�:?�V��M�>�����.v�e�>W���6i��oC>��K��=zy�<8O=��W��Ѭ*�Q/&?��>Lt�>��4?A0[�DG��G����,����>'By>��>O.�>�6��C����c���i���%��_t>��b?�vK?'�l?c����/��e�� �xk-��쩾l^C>��	>"��>#�T�P����%��>�2q��������
�Z�{=d\3?��>�H�>ND�?#�?E9
��Ƭ���}�Ӳ2�y��<�5�>�i?t��>�>E��t2���>��l?��>��>6x��MO!���{��~ʽ`�>P��>J��>�o>�,��
\��W��!u��!9����=��h?N����a�g�>r#R?H]�:$-L<�B�>�v�ݷ!�����'�e�>�?�
�=J1<>M�ž�F�֠{�,��RJ)?R�?Ņ���2*��y>7�"?��>q�>;4�??��>��ľ����#�?��^??&I?�A?p��>�= ���`ƽfR%��� =8�>WX>B�g=��=�4���[��y��
N=G��=��ۼ�M��0<�~��N�<�l=�5>[ؿ�H��*���
����������k��"��:���y���Wʾ��������j����<O�8���X��Z��l�v��?fQ�?�����ԾY���eB��k���AR�>0�꽚�.�jĺ�s5齡���L׾�r���x���X��v�B���}'?��s�������ɾ�f/?#0?3ԁ?�9)���@�8�X$a=�ݙ= ��<^T��A����������T?�~�>�����Q����>E3>[T>ۭ�>��9�}@Ǿv�m=���>w1?�R�>T\.�g�ѿ\6��kO�=h��?��@�wA?��(������T=~�>�	?ZI@><�0�>������5�>�$�?�?�=M=�W�����e?�(<��F�K�ໞ=�=
�=�U=v��J>hM�>�d�.6A���۽5>���>X�"�����^��T�<��]>h�Խ����5Մ?+{\��f���/��T��U>��T? +�>H:�=��,?Z7H�a}Ͽ�\��*a?�0�?���?#�(?;ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�څ�=a6Ἱ���x���&V����=Z��>^�>��,�ދ���O��I��Z��=�����ѿv������*>��=�|�������'G�<̃���k�в:�/;�Ղ>;�>�L�>�?�>L�>5�U?G�k?�@�>���=-�i�|7���
���Ц=�u��猽I��N:+�L%�����־R2����@��0�ȾJr=��>��7��ȋ��4R��mY�"1&���5?Y�,>+����,�XA:�g���?���
C=�=����<+��օ� p�?z�+?���6�O�"���>�͇���U?�]	�r&��u;�N��j�G=s�=xW>��<Ŝ����J�ܡd�E�?)?𾐾oپ��=I�&�G��{0&?e(�>��	��ݼ>�_?��?��G��Q>:0x>�u�>ѽ�>�JC=E%̾�v=��2?��f?���<�"�ۙ>�����M+���c�>��,��df<˩�>iGC>E���5��O&����<�V?3i�>�;)�����⑾��.���C=�]x?~}?�W�>P�j?6OB?Ɏ�<G���S��'	����=�mW?�
g?e&>�� ξ�𨾐@5?�*e?�E>�Dh���h/��=� ?��m?�?Ɛ��=@}��O�����K6?�v?+.^��^�����QW�$ʥ>ߍ�>#��>I�9����>�>?3�"��7��V���fe4�hƞ?�@gu�?�(3<%�����=e6?��>%?O�a�ž�ﴽ$}���p=,��>����^v����Ɖ-��`8?Iw�?�4�>u������%$>����QH�?8
�?�\B��(����o�If��{;>r�=ƿ[=�~��-����%�>oپ��ݾ8�B���:>��)>��@����o�>�R/=�8޿��ѿ׹��kC��𾎛5?w�>ᗼ�k���v��Mf�ŲS��i�:���Gm�>��>���������{�ǖ9��A��j��>���>lkV�	�������W<ϒ>Y7�>WC�>���!1��/��?���� ο�����i	Y? ��?l�?
�?�^�<L<z�U}�6��>�F?�Nr?�=Y?(��h]�f�5�ĸj?�T��55`��l4�JE��T>f 3?�G�>Ϥ-�H�}=`�>_��>��>6/�x�Ŀ�嶿K���b�?5��?�}����>[}�?�+?�c��B���]��G+��X�C:A?��1>�6���!�43=������
?�t0?Ow���6�_?��a��p��-�C�ƽ�ۡ>��0��e\�zN��j��aXe����3@y����??^�?D�?/��� #�56%?+�>y����8ǾQ�<���>)�>�)N>�E_���u>s��:��g	>���?�~�?fj?���������T>��}?%#�>�?�o�=�]�>^�= k-�[o#>w�=�
?��?�M?FJ�>4U�=��8��/�XZF�@FR�$���C���>l�a?��L?@Nb>����/2�
!�sͽ�`1�VX�]]@��,���߽�)5>R�=>�>��D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�f��=��7?�0� �z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B�~�1=8M�>͜k?�s?UQo���i�B>��?"������L��f?�
@u@a�^?*E�ҿȆ��:t��}����8>�×=�� >����>@k�=�Kʺ���v��=U��>��k>(M�>�\�>�;m>{�b>ﶇ��-$��{���ћ���9����>�	�-i�D�
�$[���RѾ˂־X��"ҭ�5m��#���ͽ� �<�"�=��U?o�R?h�p?a� ?{t���&>���E=W�(�@��=��>�1?�]N?��)?�E�=�W��H�c�U��=া*2�����>gJ>�C�>���>��>��;��H>�F?>S�|>���=�=�W��:=�'N>�Ī>��>���>[��>�.�=�����J��ׇ|��Ԡ</�F��ԗ?����������v�پ�vľ8ȳ=&hB?M�=�ꁿ��ٿ2���O?����~7��O9����>'=6?c�?�X�=o�Ѿ>�>!z��U�ٽ�ξ�=I�����e�0� b�<H�Y?��>�X->C�t�=��v>�����5�>�:?yu�K�胿"4Y�Zꌾ����z?�1=�pD�=3����T�U����=�of?��?�� ��S��S[˾!*�3B�>�	v>�%>Z=>H�M>��=�5��d9��>�T{>�.>�?-h>��V=W�D>�^������z�>0o>��>C?$�?�\0��ܲ��vž/�\��X�>��?�%�>�(�=�[�&��=R�>P� >�iH����k_���=��P>���2Ma�J�ǽ�5=��|�=���<+U�b�:���= �~?f���㈿e�e��mD?Z+?X�=�sF<d�"�) ���H���?O�@�l�?�	���V��?�@�?x
��"��=P}�>�׫>ξC�L��?��Ž�Ǣ�b�	��(#�iS�?��?9�/��ʋ�bl��7>L_%?p�Ӿ�i�>�r�UX����W�u���#=P��>�:H?�]����O��>��q
?N?$Z�֧����ȿ�zv����>�?���?I�m�@���	@��|�>̠�?�iY?�zi>o۾�XZ�7��>��@?�R?��>?�;�'�?�?�޶?f��?!<>�m�?9@�?�?N@>��Q����'Ę�:��=�ڽY��>R܂>lz���A�{S��W����RV�����M�>M�)�z��>ڨŽ�3�b�>�H��<�򾚹.�y5�>$v>/�>���>��?&�?;Kb>��>b9<xҥ��˾L�K?I��?�����m�T��<�7�=�Q]�E0?��3?!WA�Jо�̧>>�\?���?P�Z?�Z�>�r��)���߿�A���<��J>�m�>���>߇��?M>��Ծ;D���>jϗ>M��_ھU�������>��!?=�>��=k� ?�#?{�j>�*�>H_E�:��^�E�$��>ݢ�>�G?X�~?$�?�չ��Z3�����桿K�[��:N>��x?U?q˕>厏�����:=E� DI�����~��?Ltg?T��?72�?�??��A?\'f>���9ؾ������>q�2?���|�^6)�x�a���R?�[6?`o?�Ӿ��ͻJ�����Z��宾�M�>|�>?�;�>��(���������<��������L�ٽ}=���= Є>���V�u=}��=xR�[�z��m�<e4o��=�R�>�>b��=-�����&?7�=������0r�)�G��ԍ>��x>'���q�_?�E�ۆ_�P��� 4��8���cՍ?�1�?Ί�?�����\�\<0?�G�?\�>�i�>�u�����yھ��n��Y�� ���*H=b��>�н<�̾M5��tũ�N�w�0X�7�)��|�>��>�o?�	$?� $>.R�>5)þ���q�(�q&�jw<�6%�y���C���s2��]Ͻ���<�
Ӿ^󍾻��>���k,�>��'?�@>O4�>)��>1(�$�>vF>a��=o�>dP�>�/�>�r >Eb�=����JR?{����'�	�辚���6B?od?�3�>�:i��������wu?�?	r�?�8v>�zh��'+�jf?r*�>f��m
?l:=���)�<NH�����2��YD�/��>�d׽%:��M��^f��f
?�0?C����̾�8׽Ą��8Qo=O�?)?��)���Q�a�o�m�W��S�����h��Z����$�͜p�쏿9^���#����(�7�*=�*?��?���̣�l��$k��$?�T8f>j�>Z�>��>h�I>a�	���1�	^��H'�T����J�>gM{?���>�G?$h;?��=?��B?*�>}3�>w��+�>�{V����>��>�,?��*?!?,?ҭ?�v?�Ev>~�s����B澜�?P�'?�?�?R{�>�Ym��&������1a�����U+�>7�=���=��/��P#�zl�:/�M>?�
��W@�7�ڬU>�7=?&�>j��>߮���}x�#!<��>�?��>��澫�m���F��>��~?w���>=��.>P��=p#�������=U��g��=Z*�����2Å�`�>!ur=*]N;���<V�l�	��<R�x<�)�>]�?�C�>V>�'��? ��z����=��U>VDV>�6>@E׾�����<����g�fz}>�9�?�γ?��U=6�=7�=�4������ҏ�c��P�<�g?H�"?��Q?�v�?�-;?y{"?{�>e���꒿�ԅ�������?U+?�n>�����T��T���D�^l?�m?�\������$���� a>)B>�@j�����/���8����>U������M�?6��?L%#��
|�ɾ,�����B?�é>~�?��>��#�a���Ӿ0��9�>{��>�Ew?Y�>��v?BD�?<�}?���>[Z�,���������?���=��?�?�?2��?a1>��>k\7��	G=E��l�<U���O���>x3�<�Y�>� ?���>���=g:���>�y^��*�=��>j�>=��>�o{>��=��
�e�5?���>��۾��$�CP��������>�c?w�K?�C�?	=G> ���1q���Kʾ+E>���?��?��"?��˾�x	�s;�=b��d����B>����f@>э>��=0 �=�?_�?�[M�+�:��^#��ä=�N<?�F?�'*>Yeƿ��r�Ҟq��O���V�<�/���e�����EZ��c�=��������6��@]�����𰒾�$��W&���uw����>m(�= n�=���=~��<\���g.�<$�R=�/�<a�=	�z�l�R<D<������Z���:O<j�6=����˾�}?�;I?:�+?��C?��y>>>��3����>\ǂ��??�V>�Q�&��;�����!"����ؾ�p׾6 d��Ο�mO>9UI�1�>xK3>�7�=�w�<
+�=�Cs=I�=�@Q�H�=/�=Az�=�|�=���=[�>�P>�6w?X�������4Q��Z罥�:?�8�>g{�=��ƾq@?�>>�2������zb��-?���?�T�?>�?@ti��d�>M���㎽�q�=I����=2>o��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�@>��>��N�j�0�~�j��IQ��W�_"?��6�@þxWv>�Å=<�վ�̾��=^�4>��=l�!�$U[��=EXz�>�;=z;s=��>�cO>�ǵ=/���M�=�%X=���=�T*>�{�;$v^��L�8��<<�=m_>��	>X��>��?k�/?ۭc?�>7�k���;�M�����>��=ᑰ>iς=�?C>S��>H�7?4�D?��K?z:�>CH�=1[�>'�>{,���m����S�uֱ<`�?f��?G׸>6h�<e0>��9��>��Ľ��?��1?� 	?�F�>���]���d��i���v\>���=�ף=~�k�Y"�=�O��U�h���<�������>ɑ?x�>ߝ> �>���>G�>���=��:=ok=�ʽ9�<�^�=� i>�����ު=��z=�n<�,�=W����z�=�5�=�j=��K꽑V�=�7�>/�>ԍ�>Y3z=�,���p!>AC���yF���=�8���<�Aa���|���-��y!���R>�P`>t̓��Z��hK�>��r>׏Y>���?+�s?>�c�֊˾i����OW�w�L�|�=�5>�-�WI<���g��iH�8=ξﶯ>I��>���>��>�6�,l�$��=X�
�Վ�^7�>������5>K+��l�G�|B��G"����G��NW=& n?�ψ���>9]/?�
?bw�?g)�>Xę�b�6��?����OM=�
��A]��g��wh:?Jm?�k>$l;�%`��H̾E���޷>�@I�2�O���R�0����0ͷ�8��>������оj$3��g�������B��Lr�Z��>#�O?��?X:b��W��KUO����p(���q?�|g?.�>�J?�@?�%��z�r���v�=�n?˳�?S=�?{>	�=�n���>~X?��?�?{k?Nn�T�>h���h	7>��>�%��;�8>�<`��=\��>�(?b�	?y���0��AԾbݾ��]��a�=��>=�:�>��>Ɏ�>s�>�F�=�R�=/_>j�>��>��b>���>���>Uܞ�q��:?���>���>6Y1?�l1>2�sew>Y禽�|*=�\H=qd@�|��=w�3��O��s�k�i�\>��=z��>mNտ��?p��>�+.�%t?-Q����>]�>͵k�M��>���>�ͣ<?��>��m>�y>�<�>y��>�����?)>��� ���/�e)���ȾAޢ>����)�L	��^G��)��>8��־6p��|�b�8����<���?����o���q����?���>�CF?`�ӾS� �Q�|=�2�>;a\>�Ծ8��뫕������?��?�;c>��>@�W?�?ْ1�3��uZ�"�u�g(A�$e�R�`��፿�����
����*�_?�x?+yA?)R�<:z>N��?��%�_ӏ��)�>�/�!';��?<=x+�>*���`�z�Ӿ��þ�7��HF>��o?:%�?yY?=TV���i���(>�;?�2?�>t?@1?_�:?����#%?9�0>��?��?w5?ܠ/?u�
?�3>���==b��*!=�Ւ������ϽP!ɽ����a4=�~=^:�C<��=4p�<L�����޼܈6;�榼(+�<�:=f`�=V-�=%��>�"^?���>�\>��,?�v+��2��W���(?1nf=#�t����5
���t�"��=5�i?�<�?�;X?@#L>^�I��@�Ah(>�>�5.>3\f>���>�����:��j*=	M>u��=�z�=V/�g~i�`b��ꦾ�ԁ<D�)>(��>:�{>*����%>f��4w��=c>P{N�T2����S�<�G���1��yt���>'�K?�?I�=~=�`����9f�i�(?Gz<?��M?�R?���=�ݾx9���I��A�Jl�>�B�<���ס����;�:�T��;5�u>~�������J�>�W���]Ih��b)�5K���4>�U �֍�=C/���n��:���B�_>l���<������������O?�>�=w�m�$�\�����>��>8�>x���Wc='�6��;���{I>���>���>�5��Q\Ӿ�]�� ľ��>��A?'�[?��~?4	��(mr�_=E��o������j?�$�>Đ?��J>��=�מּ����
f�CG�Ho�>`D�>.���4H��G��ɫ>�8�>��?O}@>��?��N?O�?�Z?�*?��?�=�>����=���p?8"r?�<[=�m��ٶ�u�P��4�_�?��?�H���[�>'?>�/?�.?P/V?e�?�j>�f�D8@�}��>��>��^�?��X:u<T�??](?��"?il?��>a7�H(�-в�R!">��D�J�3?�4?��(?'��>���>魡�Z
�=���>ac?�0�?��o?Y}�=<�?62>e��>a�=��>���>�?�WO?��s?��J?���>���<�;���5���;s�U�O�&C�;~nH<��y=���?1t�&L����<!�;.���@�����J�D�k��K��;g]�>��s>���=�0>
ž������@>�n��4N��}���ye:�R��=S��>�?���>�6#�X�=f��>�!�>���3$(? �?�?b�!;�b��ھ&�K�P�>��A?���=.�l�ㄔ���u�M8g=��m?ʋ^?KW������b?��]?Ig�=���þ\�b����O?�
?��G��>[�~?8�q?n��>��e��9n�����Cb��j��Ѷ=�q�>$X�E�d��>�>��7?�N�>��b>&#�=Vt۾�w��q���?O�?�?���?n**>}�n��3�pg�)���T`?��>������#?P�q�߾´b�v���@о���������5��3'���x�)�d�����n>��?�+u?�e?R.c?����Gd��S�SS|���V�HU�
-�C�R�9G�;�=��*r���!B�r����6�:�E���W�><�?�E??ᜟ��
?�Cо���˽�0>!q～�>z�T>GS��C<<ǰ=B��xg��"���)?K�>Z�>.�??�X�̽F�ƴ3��R4�~�V�>^��>�g�>G?�>��D��;���$�"�P��Z���<סu>S�^?��M?��d?�����&��w������>�)᭾H�?>��=0�>�5���;��}"��x5���o��r��{�D9�*�4=�$?)�T>T�>�?R�?#���-���/���R8����=02�>k?vG�>	C[>H!;�j�����>,i?#��>���>	e��x�Rxz�g|��r�>�p>
F�>�_>7�/�^�B������\��7�'�F�=�L?�mu������M�>��K?�4�;��=}�j>saɽ�4�+ʾo7C�L�t=²?ɟ�=r>Y�Ӿ�<�<�����tW)?�<?�Ӕ�$�*�ws{>N�!?�~�>r�>D��?�C�>Gž��^��=?�^?�J?s�@?��>��= E��]<ɽr�&��5=��>�W>T�f=8��=�R��\����D}L=d�=0^ܼ(P��U�;kǳ�W]~<�/ =��5>l6ӿD�Q���˾����:��J'޾njl��%N�\GǾ���3ξ�=̾�o�CŦ�8o@��H���<�2Ǫ��W�����?��?�����D��= ��{~���־��>����Mܰ�)��W�v�NÒ����ɰ�����:`��������P-?�u��U������v�־~]=?�*?�A�?+\0�x2�w�8��Q�<�@>�nD���ݾ�6��\�ǿ>��8�]?at�>�z���R*?�"O>	�=[��>��}����I5�Fz�>)?'?�>�D� )ο����㋽K��?8@G\>?o�=�2���>���>x�?�G�=gpt��8��֔�q)�>'�?��?>I���+N��#ټO�e?F>�=�C#�8|=u��=�?I=90
>qF|���>XE�>�_6���p��|ҽ��={ �=xG��;%��݂�P�~<��&>v��P��4Մ?({\��f���/��T��U>��T?�*�>C:�=��,?[7H�`}Ͽ�\��*a?�0�?���?%�(?>ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�̅�=�6�;���{���&V�w��=T��>]�>͂,�ދ���O��I��d��=�V�A�Ϳ���Q�
���1=.==<l���`,ż�@��6�$>���uڧ�
��R��= �<>���>oo�>ƹ�>��>�W?�o=?�+�>��z>�.���M�����m?a>��������x���lѼ~u$�ݾ��!�_�����/�.W�F�9���=�L�����.�K2[�J�6���,?)�=P����Z��:��&���,��/�:�,����˾T,=�x���?�	P?�����f�A��y(ý)嗽K�V?��̽E���Գ����=<��;`�<��>�=Y��4*���V��$?�-?����{N��6��=D�O�6�*=b+?Ϣ
?�+��ڭ>�?-�x��8V3>˛k>Z��>���>Y$�=D7����$��W1?
�V?.)9=�`2���
=��ݾ��4�	{
���>���C{����>����[7Ѿc�����׽�!W?9��>@�)���~v��f��==�x?�?�=�>hk?��B?�G�<�u����S�/��x=�W?i?)�>�?�ϾV^��q�5?�e?�N>k3h�0����.��P�?m�n?�R?7Ü��p}�������Vf6?��v?�^�<O�����W�<e�>ڬ�>��>~�9�`��>J�>? #��Q�������E4�"��?ٓ@|n�?�m=<��=I�=+??MR�>��N��ƾO����'��X�r=��>f����	v�Hb���,��b8?��?�p�>B�������M>bI��'��?Fk�?ݼ��4=�9)����O��5�Ƚ�Ɛ=B�=�ԅ����ژ^��*��B��@J*��y�=��O>�K@�r�Jz>FǽNVͿs��}��뾾f����>�ff>���_&�C9��`��=�d�>q=��>Ծ��>^;>��P��St�u0)�*�p���>�hr�6�>0Y��Ž�5PO���f<'��>��>�0y><�e���xL�?y���˿쨛���
���c?HD�?��?�: ?�т=Y,�� ��&A=+"2?%�{?��B?0}���f��
N<K�j?�y���]���1�ټD�.U>g�2?���>0 .���l=e>j$�>ȴ>� .��eĿj����>e�?y��?�r�,��>ci�?�/?�U��L�����(/��a�<ݰ>? �6>+D���u!�n;�����d�
?]�.?������]�_?)�a�L�p���-���ƽ�ۡ>�0��e\�TN�����Xe����@y����?M^�?g�?ص�� #�f6%?�>d����8Ǿ��<���>�(�>*N>0H_���u>����:�i	>���?�~�?Rj?���� ����U>�}?
�>��?*��=�/�>~�=	���*5�(�#>lC�=ADA���?ڔM?!�>���=
�8��/��6F�-R��)���C���>��a?!qL?5)b>�r���c4��� �
:ν�1�4�鼒%@���)��߽2$5>z=>��>]�E��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��[a~�!���7����=��7?�0�M�z>���>��=ov�ݻ��O�s����>�B�?�{�?��>�l?��o�=�B���1=GM�>k?�s?�Ko�~�U�B>��?������L��f?�
@wu@V�^?�=�����ٱ�G.���%5>:�@>�^">����\">\�����Y��R��@�>IU�>q^�>s{>���>X�m>��o�#����������4��C��4�m�]��}�=��� � P��B\f������z��(P�'RI�� �������=��U?�
R? p?͈ ?�y�ub>���m=��#�0�=8�>�\2?q�L?�*?"ٓ=+���6�d��^���9������ǚ�>D[I>�i�>ND�>#�>�ҕ9��I>:B?>�x�>� >(=���=G�N>�G�>���>y}�>�}>9�A>
�¿
���X�L75� C�=V�?/��)������^�پ��6������g?6�W=~J����ؿ�ѩ�
�C?�򛾠M/�TS{���<>6A?�m?{�8>�#��=G����=LAg����SS�=t5ȼ@�#�P�S���7>@�$?=��>�n�>�eo�E+0��TC�$ǁ�3?"?��i�=_}�U+N����$*>�'�>6�=��(ё��U����w+\<x�[?A��>+���d#�������ݽ��f>{� =��>�ǒ>R�=!�=����B���ff>��>�7>��?NO�>�*�=+�<���#u�1��>���>GA�=�O?�M?<�o�	Z!�^�쾛F�.�>��=?@J�>��>7 5��>�L�>�>4f�=�	u=�\�gm8���>D��p�f��ܼ�
>�@���j>�f�=�f��G��Q[=�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l�6>�^%?��Ӿh�>,x�QZ��w����u�d�#=��>9H?+W����O��>��v
?+?�^򾴩����ȿ0|v�j��>3�?���?B�m�uA��v@�G��>��?�gY?pi>�g۾@`Z�h��>��@?�R?��>�9���'�0�?�޶?�?��>ޗ�?]�?%?��>V'#��>¿<����,>���!?yr�>_��10�Н�����q�<$��~�>r!��x3�>j�=��o����h��3�ϼ̀\>�{>d�?���>Ċ�>U��>)Z?��=����'&�5�V���K?�ߎ?�5�QKm�m�<�ϝ=CQL���?��1?ƧZ��:վVA�>Y�Z?LI�?��Z?�k�>$��7���r���^���}�<->Q>���>Up�>V���J>�2Ѿ@�@�+`�>Qp�>�b����ؾ�뀾�9E��M�>�M$?���>���=� ?��#?�j>�+�>m\E�c8���E�v��>Ǣ�>�C?&�~?w�?Xӹ��W3�0	���桿g�[��=N>0�x?�S?�ɕ>���������dE�;#I���I��?�pg?�Q��?41�?�??8�A?-2f>@��wؾզ����>W�&?����rnp�( �_N��?�,?a.�>��b�+J��ą�h�1�ؔ��>�o?P�?�#�@}��� ����<u$<�=�+p<T4���!y=rE)>q�4��6�=�>��>�@��qD��y�= �A�-ى>�2>���TD����+?͟O�����u�=]r��D�G�>�tP>�꼾�[]?:��z����F
��{�S�,Ӎ?46�?��?=���?�g�B6;?��?e?!�>4O��,.⾓��,o�<����;�i	>i\�>����p�ˀ��io��K����н�@��>�i�>�?f�?�D>F5�>���G��~���B���T�>C��u'�2� ���٧�r�Z�_;��Ⱦlc��!(�>0zʽ���>%�?�Ub>t=�>�>�^���>R#Z>�Z`>J�>���>�Z>Cx>N��<�w���FR?T���3�'���}���-4B?�kd?�,�>��h�w������
y?M��?mq�?1v>�h��/+�!o?iH�>����f
?}4:=A��歊<E@��e���6���c�[��>�N׽N:�lM�q[f��h
?�.?:F��Vq̾�׽�j��V�o= N�?)?v�)��Q�g�o�3�W���R�����h�a6����$�>�p�����c���#��ӊ(�C�*=�w*?�!�?������7!k�
?�bf>���>��>���>��I>l�	���1�I ^�en'�ƃ�;i�>E{?��>�?H?��A?�Y?,�^?��>�J>�����?ڐ�����>b�?��:?��9?�V$?�?v+?�A�> ��'��0�Ӿ��?-~?��?��?=:�>��S�������.W �-e������~;A�=u����|ּ: ]���{>&[?��ԡ8������j>�7?�{�>[��>\0��&��w1�<���>��
?�<�>�����r��f�TG�>q��?	���`=x�)>I<�=<���n�ݺ���=9i���א= ����;�ɵ<�]�=���=a���й�Y�:+�;Jѱ<҂�>�?�P�>�Ç>�����&������=9�W>��T>��>��ؾ4���y2��o�g���z>0��?�W�?�wg=���=���=ԛ���o��3_�f�����<��?}0#?� T?Z?�?�=?��#?4�>���'˒�
���
���p?݊/?���>��[h��й�������?:?��i����(�t�̾Q�=yX�= �8��ȉ�=m��.�yy�=�@� !��-�?e��?���4�U�?<ƾ�բ��"���(?:3�>��>���>x��l�t��'����=�?�]?��>�P?�߅?�Zb?��>Ag!�'���ܩ���48>�S=lRs?6'�?��q?w�?�x�>�2�=>9�fwv�����_���OMľ�k>���>_��>���>�%�>���>�b�=����?���D>�)�>&@ ?�?m�?��Z>!����7?���>���^~8���7K�U�>6�l?�|J?�M?�*>�����m��~����b>�5�?#0�?��?�'�}�=\ڌ<�]w������>�2�>/�>�>��,=�=���>�ˁ>������E��{'�E&+��m?��_?_h>+!ſ�o�=}r���M��;^]��c�"f��`Fa�*ӭ=�ۛ��<�Â��g�f랾ς��	���Ϋ��ʁ��>ʌ=g��=���=���<h ϼx�<�_W=ۖ<�7=�a�tʔ<�(�7���9��e�p�N<f�N=!3	���˾��}?�;I?�+?��C?u�y>�9>G�3�⚖>A����@?�V>o�P�&����;�˫�����͵ؾ�w׾��c�ʟ�vI>%_I�{�>�93>�G�=9L�<��=�s=�=(�Q��=�"�=�O�=Lg�=���=��>�U>�6w?X�������4Q��Z罥�:?�8�>g{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=J����=2>q��=w�2�T��>��J>���K��A����4�?��@��??�ዿТϿ6a/>�b >;� >W�<��)@�C>��t���&=���)?8&@�8����4D>s+i��ؾi���>�=�p'>�v�=�<�-�^����=I�A#�="�	=H��>I>��r������ �=�A�<��>l��>���=��O��=�"�<X��=-�>_�>���>��?��/?�`c?W6�>)�p���ξ�����>��=;A�>�j�=!�D>j��>��7?�}D?T�K?@��>;~�=1ۺ>�[�>b�,���l�xD�EG�����<�X�?G��?��>א><��E�����=��Sɽ�?(�1?�	?��>�����,�!�v�$��=�K,>�6�=f;����̼6b��թ������Ļ6��>q��>�v�>���>%��>��>��>�Q>�I�<w��<�Ԟ�#���2o����=� (�8H=�^��&2������퟼���q	>�,�=2����;]��=S��>Y�>z��>갇=a͵�u8*>�Վ��ND�%�=�ʠ��B>�>�c��z��G,�S7+���I>{*a>ZȆ�F䐿6��>� o>�mP>�r�?��s?���=���ĒѾ�����]�xP�}��=®>�vE��~?�F1a��ZL�:0۾$��>�m�>[��>��>����3��a>��߄��kN>��`��R��+�:=�3�Ií��f���I}��v>�jh?BU��W�K=�Q[?۷>?u�? И>�Q��z�?��?�^��Q6?>�y��I�־�8>�m?�RL?�?w��9��H̾*���޷>�@I�6�O���J�0�Ƭ�0ͷ�C��>������оi$3��g�������B��Lr�R��>�O?��?O:b��W��JUO����t(���q?�|g?+�>�J?�@?"&��z�r���v�=�n?ɳ�?T=�?�>,�a=���V3�>O�?	�?�y�?��a?͢i��X?`W����>�����=zү>E�j=��=�-�>�???6Iƽ\�6�Ҿ9׾��:!��>|�<ͯ�>é>$i>��t=RU->ބ~=���=�h�>Bd�>�G�>`Ş>�B>�g���-�M�*?��m>�Y�>{ZM?��@>9	�|y�=��%W�����.��Cļ�+ڽv�=�üQ>��y=���>n�¿���?�T>p|��u?���Lཇ�9>��>�q=�c?��>��&<�ܝ>X�>蔃>{�b>��d>P��>>dkݾ���f�8�}�QOҾ��>�ھ�M⽖���U����<z����5ʾm1s��|��>���<�y�?a.�K�c�tE�����.?%(�>3�T?��;��h�ڃ=go�>��J>)%���%��������^[�?�)�?�;c>��>G�W?�?ڒ1�>3��uZ�#�u�f(A�*e�L�`��፿�����
����'�_?�x?/yA?�R�<#:z>M��?��%�Vӏ��)�>�/�&';��?<=h+�>*��2�`���Ӿu�þ�7��HF>��o?7%�?lY?@TV���{��O>�sE?�B?@t�?�!3?�?��Y��n1?q�>=�?�?:A?x:?G�?�$W>�< >�v�<:O�=��������C=��g���7�����=.ث=��S����"&�<���<FS<s�;I)Ƽ~�λ�޴<�=;��<�@>qK�><8^?���>`��>/�3?�c%��S5�<��rW.?��>=��|�A߈��碾�0�=�nj?���?�Y?��`>�DB�W\C��">䝍>_W,>Sd>���>�m��}�@��k=Y	>y>���=pB*�
쀾,
����G�z<+�>���>RV}>ޖ��'�%>����mq{��'d>� P��ٻT��TG�Ӟ1���w����>�FK?[�?TO�=��b���S f�^(?]�<?�MM?N�?���=F޾��9��TJ�Ѐ��C�>Ե�<B��
��^�����:�� [���s>r7��_������>�ǉ����r��D͏�q�i��ub>�W�!��l�����'����Z=�
�>k����Z�;��� ȿ°&?��>eG��`���� :�>"Q>�\>���>�ʓ�u`��D�=�J>�?��>q%>�'��&$��<�ތ�>$�8?�{7?�g?������r��h@��D��g��k=v�>�
�>O��>aU��0�=>D۾l��0RX�5G/�i!�>�L�>x+��JF��@��u���og�j�=�(?�>�> 2I?D)?��5?���>p?g��>}!w��` �|?!�h?>�ʽ�z۟��4����>2�/?w��	���s�?���>:�>��)?)�(?
Ћ��R"�����7�>`_�>�@S�紗�
��>y�3?"�>hY3?O�?��y��cC����<��6���R>�C�>:�T?�.�>�E�>!�>w�>�a�J>��T�9?�3o?��c?��?r��=@V?�>)??���4v���?.��>�_Y?	]�?��?0,?	5����V�

�	"�e��=+�<p�x.�=��M���v=�h=ƻ��#��9�=��c;�y���&�Kq�����= �>��n>}D��kA>қ��A���TTQ>g��0���x��i�.�-��=�*�>�[?5�>K��	�=K�>��>���z.#?|?@l?�ZA��bd�N�׾$U@�g5�>8�@?���=uj������:t�暋=��n?(_\?�P�8M�Qb?s�]?W��<<���žH`�ܹ�q�O?F		?< K�l�>�|?Z�m?"I�>�^��k�+V��v�a�gf����=��>C<��2e��-�>#�6?F��>$d>g�=[N�N�x� ���M�
?�?��?�ފ?AN'>Z�m��߿GX�r���΁\?�v�>�r��q�%?�$�ɽ�j������X�Ҿm\��'n���1��ڻ��y���↾��ԽZ=�=�??iq?R&l?4�[?D���'*a�<ia�-}�pFU�3!�&��ܱF�J�E��C�Vs����V��%���Y�=`�f��??��^�?��'?ʚ�G��>p�����^�Ͼ<�m>�3��h�Խ��=�ƽ#a�<J�=g�H��m����J:?<�>�ĺ>��8? W�g�6���'�:�B�Q���K>P�>��>���>��^��n7�:��̾�?��m��qy>	[b?UjI?�l?�T�ZR0�g���,]��O;�@��� 8A>U~>�e�>jv_�w��$�:P=�&\r�����Q��|,��h=�;0?Az>j�><��?[?J��7��x�H�.�^H�<ì�>mKh?y��>>؆>nҽ��@�>'X?���>L��>Sl������W2|�p�<��f�>�@�>O�?�6>{]����t� }���Ј��2<���=��m?��r�k,��p�>�F?�̓�/"m�X3�>ݖ����nо�0�@
�=��?�+ >+-�>)��X���Z�w����ύ(?"H?x1���k(��Z{>6�?�{�>w�>)��?ǔx>:�ξ���<l�	?��T?��H?c�E?!7�>��?<r��G������o�<�{>al>a�f=R�=P%���S�C5.�"0=�ۻ=��ԼFʽ_y�<|�͹�_:�&�<�a->�$տG�A�֤���y�n󾚱,�p7�����V������Fŕ�#5�T$��M��`X��ھ,���	�����T���?�A @���=��ӽ���}v���x3���>��P��w[��:�=t������j�
cD��;s����Y̌�sx(?6��y�¿������㾾�!?�?�v{?�/��,$�Ar/��>�ũ��(�[���O��Z�Ϳ��ܠ^?�y�>����Lt�>E�>�E>80>�n��վ���Z*<�?&&?V��>��z�&˿΀����#�==�?x@�I+?�*�=!
=xm>u?;�1?���=�3��D��C�S�!?U�?u��?DM�:^�~���N>�/�?�_m>���\�׼;"�=r�<�V�=�H\���>�}a>|ea�ӗ�яؽ�ٝ>H;_>\	�K����=�J)�r*9>�� �!�!�5Մ?+{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?_D6?���>�d&��t����=w6Ἤ���|���&V���=Z��>d�>,������O��I��S��=O(�i�ؿ�%]�*C<���<�C���s������=4�X>�m���ž��Ƚ5�6>�Wռ�_=UL�>�`�>��>�OB?X�I?�??hO>�+ͽ@���뽔��{O>�0ξ@8A���ҽ�C�*�r���澑eپ�徶G��B(����Ͼ0�6�Z
�=�D�|��G�)���u���Q�o�+?�<=ɹ���E�J�A�}�ԾJ���E�3=1v?��v�
�<���p����?x�E?�[z�=�O���!�����	�@R?�Oֽ�o�K����%>�J�;e�=�ֳ>�+>�پ��L��W`��-?0@!?i���N��=8��n,��.�=�?��>V��JH�=_��>�3��1����>��x>���= @E=�]Y=�C����P��.?\�S?Fs�_N����>�Tؾ-�����
?�>D�!�<�I>ȱJ>%�G뽾�7�>o,>��ƽ��V?ℊ>KW#��|�w松�����>=i]{?L��>�	�>{*j?ȧ<?�������9�M����t�=}N?4+f?X>;I����ξ9n����5?|}b?`�>��N��C�,�3����?^?M ]?c�?��Z���y��n��%{�	�;?��v?s^�Vr������V�lH�>�k�>��>R�9��m�>֌>?$#��G������X4�Ğ?��@��?�y=<��-��=�6?dX�>�O��/ƾ!W��<���Έq={'�>����cv���s,���8?��?^��>򒂾O���E>�<��z��?b�?��ٽ�u�>]���Ys��[3����>��>'�>�"�>�����k��۽ꓗ����<�}�=Y2�>*�@��g�x�>O��)�q`��.���R��츈�5��>z��>���.�辚cE�?�}��K���2�-w���ھ>;�?>��D;�r���ԁ�lS���=�>j���'�>3�W����<��X: ���>���>��8>�����IK�?<�������l���~��n?���?Ј?��?��z�7r�-ư��Qk�*4:?Eq_?�X]?_yP��o������p�j?ĩ��_���3���D��V>N;1?���>�y-�O�r=l�>>!�>��>X*0�ڬĿ�k��e������?!u�?�����>"�?N]+?ij�L���SQ����*�ր:��@?��2>�����Y!�]�=��"����	?!0?0p��2�\�_?(�a�M�p���-���ƽ�ۡ> �0��e\��M�����Xe����@y����?M^�?i�?ص�� #�f6%?�>a����8Ǿ��<���>�(�>�)N>]H_���u>����:�i	>���?�~�?Rj?���� ����U>	�}?� �>���?���=C�>ss�=�2��Z�2��$>9�=+:<�IV?5lM?:�>��=�$8��/��0F��R���>�C����>+�a?�L?�@a>NƸ�ȿ0��� ���νS�0��@⼇??��/��Q��4>Ig=>n>�ZD�(�Ҿ��?Lp�6�ؿ�i��p'��54?(��>�?����t�%���;_?Ez�>�6� ,���%���B�_��?�G�?<�?��׾�R̼�>@�>�I�>P�Խ����Y�����7>0�B?Z��D��v�o�z�>���?	�@�ծ?gi��	?���P��i`~�l����6���=��7?S/���z>?��>
�=�nv�����<�s����>�B�?|{�?���>ˮl?e�o�J�B�_�1=#M�><�k?#t?)=o�	�سB>8�?��� ����L��f?��
@]u@�^?�����@7��3�/wƾ_�B>��$>ň�=}�U��EJ>Lj>�F����b�A=Z��> ��>�]%>l�B>{4�>��[>8Ѝ��U'�M����E�� $��� � ?,�BSϾѧ���B=�{�t���~w����Q����X�9�(��7��'��=��T?�0P?�n?;��>S����\>����@=Y=���\=���>�1?oPJ?z*?�'�=�/��r�c�EЀ��(��A����=�>ݔX>Fh�>��>���>>-~��1B>O@>�>z>H�<�mQ����<��F>�6�>v��>�ʻ>.y>(�>${��⣷��a��z�Hξt�?-o[�v6��4����z_��,y>;�1?�Ş�����PͿ5��U�%?>�;�����Q��fa>eU?s�]?:>������ǽ��=dX{�X~��G'=����W�b>�h��w�<�	?��6>Dj?��6�q�P�>���4���~�g�3?���������ӎ���b��
,��9�>��?�Cm��A�Ly��a���W{/�r����?j�G?���=6����
�����5b��F>�w>ȍ<>p7i�QÏ���鼮���&͜�ӌ�>ڐ>�n?��G>296>�g�>�{�0X����>�L�>�~��a�,?,m?���=��6��� ����t�=>}�>>p>�>���j�=\�>��g���<O�=��<�L��l-�=0^O��B���z��.����7�~�1>Ɯ>>���_耾��Z=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿdh�>px�rZ�������u�S�#=��>�8H?�V����O��>��v
?�?_�婤���ȿ@|v����>T�?���?S�m�zA���@�ӂ�>'��?SgY?oi>�g۾
`Z����>Ż@?�R?��>�9���'�s�?�޶?ԯ�?��`>���?�x?I��>��&�T�!�3�������/G5;�z!=�	�>uwO>9��BR�_4���₿�^�Q���r>�X=n�>����ķ���=���/Ԝ����ܷ>�8>�_E>5�>E��>��>���>��<ڥF��`��ƛ�gVJ?[�?i����n��O�<�3�=Yd��?t�3?��ͼosؾ���>!�Z?e�|?K�Z?��>BG��K���7����k.�<�[N>��>
��>#����R>�оP�J�Z��>�ɘ>��̼�־�0��Dѻ��>�t ?�n�>���=`�"?��?w>�Z�>@4E�����C<>���>��>��?��|?'f	?�ϾJ:�<N�����k�S�N6>�u?�?&�>���'����Gܼ�����<��?#	^?����>���?^FO?�cB?bߌ>� �|����ĽsJ>��&?[m�=��/���-�.�J����>L��>��?��>��	�8�ݽ�(���!!�!�>~"R?\�8?Bw�8�b����(Q5=%=� ���|��A��<J�>��=������=/�Pb:=��w�h�i��^��f���`>�`=�7E����3=,?.�G�Qۃ���=��r�xD���>OJL>1��z�^?l=���{�����x���U�� �?ܠ�?=k�?���!�h��$=?��?6	?e"�>K���}޾��྇Pw�~x��w��>���>��l�|�0���ʙ��|F����Ž+���%�>���>=?^,�>x*Y>��>)"Y��Q%�1n�x6վ��N�$C,�k�M�3F-���ⳮ����k=�˰�]�Q�̙�>I�J�"��>cj�>���>#�E>~�>�=�U>+$m>��>��>g�>��3>�QC>_μ8D�h9R?a�����'�	V��h��R/B?��d?��>}h�A���ܟ���?|�?�x�?�Xv>iWh�v+��?A�>
���A
?4�:=5�
�aʅ<އ��Z���8���&�g��>4�׽�:�!�L��cf��s
?�??[u���b̾ؽX\����h=OB�?C�?�(�ۅ@��Ko��IA�%VQ��~��y�0��ݡ�32�f4v�����t����څ��)��+�=_�!?Ł?�x�־ZJp��Cb��Q���>��>���>㢾>ܗJ>�%�j�7�]�_�r�(�������>��}?�?�>W_)?J7*?�8M?@�??���>�H�>g��]��>T�=�H��>�k?HTG?^$\?�?)� ?�	&?��>�n�<�����Q�4?�
-?q|?�>,�>����S�>�Fν;F��2Ԕ=�?\>���=%��EƩ�1��=#U�=�J?a���"-�̉��d>\8?԰�>�i�>�x������Xݕ=CJ�>��>��E>7���o���0�>Ʉ?�:�g=C/>�� >I��<qh�<Zg�=�E�4Ϟ=�4�:8�����;z��=�_'=OY�<V�K�V�<|x�;�.(<�x�>D�?ڔ�>�H�>N��y� �ǭ�d��=�X>�S>G>;پ ~��&��
�g�<Ay>Km�?Lp�?g�f=�=��=�i��-G��/���轾��<V�?D#?�PT?֎�?��=??`#?�>�%��F���W��H��Ь?s�?��>aھ3ї�kԓ�"Z/��ԡ>��?g�Tڃ�L�Ѿ�'ɾ|#��O-�=�u۾��j�����
t1��x^�U��K�"��?�m�?�C>e�H�&�����$�þ�J^?�S�> ?5��>��1�14^���-��{>�f%?r`h?���>�G?^/�?��c?Ҳ�>Q��� ��������_�s�='�T?���?���?�H?�0G�O�=>�g >����C��y½����¯�识=�ے>�G�>��>c֜>ou8>�.��an;��B���
>=*�>%��>�
�> ��>��<����wG?��>�n��fQ�k����|�)��^u?^�?ʳ(?]�	=+��F�*����[�>�:�?�]�?�<(?�L��8�=ݼ�����t�=��>�$�>��>�l�=EQ=?�>���>4�>�}����6��oI���?ƙC?�$�=ޔǿ�au��̃�Mk��u�<q뎾(�i�������C��~�=q"��-Y��\���oX�uÜ�����H%��x���"�r��>�y�=���="ش=y�;�f׼���<�)=�`<=Mx*�<��<�}N���o�V^���;\��;<A=��O˾${}?�-I?ۘ+?КC?�Ny>xb>�/2�`A�>�����-?�(V>�Q��¼�ڛ;�����p
��V�ؾ�o׾b�c�����>uxH�X&>�Z3>*�=F��<���=m�s=yy�=��2�t=���=�8�=&�=� �=��>�O>�6w?U���	����4Q��Z罤�:?�8�>�{�=��ƾo@?��>>�2������zb��-?���?�T�?:�?6ti��d�>I���㎽�q�=@����=2>���=]�2�V��>��J>���K��v����4�?��@��??�ዿ΢Ͽ7a/>�cH>��:>�:�
�"�1ま������j��%?2�L�ƾ{!�=K$=��׾39Ծ=C)�=�3�q�e�ONV�$U�=�]�wV�=�V�=A?M>_�A>vd�=���5O�<>�==�=�'�>=9�����Ƚ�DC=���=k�<>p-+>�d�>U�?m�2?Hg?���>_�������y�����>�k=���>Z>B�x>�k�>�(?��7?@-Q?�;�>�kK=�M�>N<�>��#���p���˾����[+�<P(u?Ln?��>w��䁾4���8�M�!�f ?#)#?59�>uF�>���և�/�~�	�Z��{<��ӻ3�*�PC����>>o�>q�Ži=W�V"�hY�>�^�>0��=֫=\��>ᯐ>U�>$)?>���<&t�<L��u�S���<��=����y=۽mE���g�R���=�����h<�S�<J��=��r=zn�=��=��>�l>�w�>�y�=򭳾cN/>�*����L�i}�=�����A��Ad�O~���.��(6�]<B>U�W>{������A�?�6Y>Η>>�`�?F$u?��>l!�F�վR���e���S��=��>q�<�CB;�&l`�Q�M�0Ҿ���>Ko�>밣>n"k>۰*��:�GB=۾~�4��t�>xr��n�(�@&��s��3���ɞ�_�i�z{: F?����@�=��{?�xH?1W�?��>����_�ؾ}�0>[�{��G= S���i��*���?�$?+�>��~�B�6̾���$�>]/I���O�D���.�0��w�=ҷ�·�>@窾�о�*3�pi��D���F�B�}Xr���>i�O?�?�)b��S��COO�����;��Pr?Qsg?��>�H?�8?Q���d�Ck�����=��n?��?�5�?��
>�>�>���+�)>�7X?��?*��?x��?㖾�x'?�(�G.'>�x\��O>f��>8_?��*�>�yN?��L?�4?�����徰���󍾜e��>�?�>c�>_f�>�01>#k�<7}˽&�ܽs�Ǽ?�s>'y�>�
L>��>�o�>���`��`yi?3ZX>� �>`�1?�	W>#�;?I�Չ�>p����r<(>>|��=����.֣>g�E>B1>`�= -;>!=���?��=>kav�_S?��!��>�i�=���>��!=�>iw�>+��=��<�ǫ>�H�>��C?]@�>�	;�9>��
�� ���C�jN���о.�>�o����-�����T���X\�,f�����h��P���N<���<2ݎ?�����h��x'��=�+�?�؛>��2?�����(�>���>���>���}Q��č�;����?Bt�?�Ac>��>��W?��?<�1��3��rZ�O�u��'A��e���`�Pލ�;�����
�m��N�_?}�x?�qA?m:�<39z>\��?��%��Џ��'�>/��!;�z�;=$�>�#����`�НӾ�þ<9�5DF>��o?p#�?�Q?CGV��x��|6>�8?�`6?�v?��8?��8?~d��f?��=#�?� ?{�>?[�:?��>k�">pPN>�U
=+4=�ƀ�?�Y�� ޽�D��(=~�<1w=9`���v]���;=�!�ͣ�����[�<Ǆ��y�!=H�+;q�g=W|�=��>�]?�F�>)8�>��8?�V�|6�����+?{�#=$ru�P�{�tP��]���=J$h?u��?{NY?�5c>r?���<�{I>��>�M%>\>W��>��꽶H@��v=�>�>�6�=��I�%U���
�,Î�Ǉ�<:k">�
�>��>Oف���>䡣��x�T`>-=��{���@L��A��n'�2V`�Z׶>��@?�7?�-�=�쾖̔��]���?��E?�\N?��w?<�=&�Ӿ��/�Q8L�bG���Ƥ>O�:� ��9��񾠿3)<�bm =A��>(��q$��3��>��	�\Ѿ�T}���u���0�q�g>z�B��"p;�a�27��ٖ�@5A�#Ｕ/K���#��������@�C?{�Y>�ξɾ��˾�@>��>�y>�煽Κ�s�]���<�5��>��>hh�>�:�>����������HR�>��??#�<? ,�?��T�|�ڌ8�F�J���q&>�D�>�I>ڔ?��u>���=��Ⱦ�{��)X��!/����>��>�l�5�Q�[�ؾ�gľ ���$|>�+?��=$��>=3V?Q��>�!A?��,?�^?hp>	��!���@�?6}z?OI�e~��v����9��=(����> M?O(�7>���>]w?t**?`�??�� ?�<͔�҂*� �>�D�>iH�	���Q��=��O?+»>��I?p:|? <�r��c<�E���PA�=Nr�=0.K?��?dr�>w2�>���>����(>"?�>_dW?��?��h?/��=�?s">i?��>F^p>�?�?�,?x�?�SW?t��>�.b<:X��W��C[�P`=-����<���c��E��6O<�n7�ap޼�@�<�
>��h�j�9�d���t)��z�>d�s>Wڔ��R4>�t��������?>5
��L���]��h<�i.�=L�~>ǯ?��>s�$��%�=1(�>�K�>�$��M'?N�?�?v��; b�jEھyH�M�>�@?2Y�=z�j�M"��vlv�U�\=-�m?f]?�VW������b?'�]?g�=���þ��b�K���O?��
?�G�:�>�~?��q?t��>��e�4n�����?b�5�j�T϶=�q�>�V���d�6�>��7?�S�>��b>�>�=Zz۾��w�Vb��h?�?&��?|��?{'*>n�n��0���ᾼ.���Z?<�>ı�9�?�EO=l������ma�/���@��DD������s���=�{{�?ܽ\�=d?�eb?{�k?�`?�:�ic�5U�j�����[�v ۾���Q�M��9�~.A� �q��8"��J꾜Fr�PXb=\Q%��Y�۽?>@?ˢb��%?��P��xξ��ؾ��>bJ�<�	��Fh>W��<D���|�2>B��Z&�TP���?�*�>>?�>��9?��O��gC�@���ST��V���k>祝>"��>���>,�j= ���<R�������%��U)�3�u>��b?I�I?�n?s��S2�����U ���L�W����<>3N>�>�OP�����'��=��.r� W�E����.	���=Q2?�π>$�>��?��?�<������w���1���<ە�>�gg?��>`3�>��̽�o��1�>�3f?�>�>�*�>�C��G2�Gfv�%@��j�>Ct�>��>��x>A�&���U��L��ҳ���2�4t>Ģd?�큾��u�Z]�>,�W?L�A=5��9;�> o�P%�IOž^�9���=�?��=&�>Bj�����.w���o�yj?@Q?�۾T�4�G��>��>��L>	�>B�?{>�c��LJ��XJ?\"?�G ?)�F?�>,߽�<�D豽=� ��nq;2�<>�ٕ>���<��;	���Ah��qOO�oH�=���=ÿ	������	�;�?m=��༞��=v)#>m�ؿ��@����*��GB�e��.F���Ir��}.�#}׽ˎ���񠾸����(�役Nv�?y�xa0�t�|�5��?�s@ҥ2��Ր�1��+��9�^�2>�>��{�����S�v~o��v����Q�ih�dR�2�r�c��%��G�'?����߽ǿ䰡��:ܾ! ?�A ??�y?��-�"���8��� >�?�<�+��l�뾵�����οP�����^?��>��=/��e��>���>��X>�Hq>����螾�1�<��?1�-?Ѡ�>ώr�*�ɿa����Ĥ<���?#�@3�3?�i��a����>ǧ�>N�?*�P>������%��`L�?���?�!�?qr�⟂�rI	>�E[?��j>d��¢��Mc>�Y�����T�B�0�>���>��!���}�dg��a�;�U�>��Z�����F����<���>��/���Մ?z\��f�q�/�!U���V>��T?C+�>�:�=ѱ,?�6H��|Ͽ��\��)a?�0�?Ħ�?5�(?:ۿ��ٚ>6�ܾ&�M?ZD6?��>Sd&���t�K��=�9��ä����]&V����=���>(�>[�,����O�O�t<�����=QN
�	ۿ����X���=7�==C��=��B��]��������B�r�a���G;�<8�=PZr>�W�>?�>Ћ�>��M?e`j?��	?��>�J!��挾�Q���=.��ƨI��f;�F;�þ���ش���W�M[��:���1���>��P>h�=��ʇ�x�V�g��kX��!� ?�0=��;K������nǾ�� ��X���������U��Q��?y:?Ͳ|�4 D�ػ�T��ԥ��P�B?�=k�`��l
����>��g�l��=
��>��>*]
��/`��ai�T?Q/?����ԅ�\;>���_J>��?(��>���z�|<���>yk��]��'�t>�-�>�uz=�#==bͪ�@Ou_���H?��l?� �������\>Y[��xN���H�>���~R����q���L>'<���w���9>K� >�P<X!W?ˏ�>��)���iϐ�����r?=K�x?2?�ǟ>^Pk?�B?PΛ<����\~S���
�J!u=(�W?i>i?*�>�:����Ͼ-⧾��5?Οe?t�N>�f��}龿/�.1��	?_Xn?�M?�7���8}����k��L6?��v?s^�ws�����J�V�e=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?��;<��U��=�;?l\�>�O��>ƾ�z������ �q=�"�>���~ev����R,�f�8?ݠ�?���>��������&>�{۾	��?g֙?�г����>�<Ӿ79r��Ua��x>;?��%>	��>͢��8=��Y�{�¾��=�\/=�`q>O�@�_w�㯿> f�<�X�@���y��*���C���!}�<O�0?���*�f�d�0X��=��z6�=焾��>B�>Q,����q��a��&��4W�=F?(F~��2�>:(5��D��� ���?��K�>i"�>V+>�s��'�%�l��?̾���ϩ�b��y?��?گ?A?�E���0�����h���ZK?���?�^v?���¾�ƥ=�j?-[���L`�p�4��FE��U>'3?"-�>�-���|=z(>Ȓ�>�T>O$/��Ŀtֶ� ���
��?��?�k꾣��>Ɓ�?�x+?p^�8��uh����*�l�5�_GA?N�1>ق��=�!�>)=��ݒ�;�
?a�0?�p�Y)�\�_?'�a�J�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?L^�?f�?յ�� #�h6%?�>b����8Ǿ��<���>�(�>�)N>BH_���u>����:�i	>���?�~�?Qj?���������U>�}?�&�>f�?���=�Q�>��=�����,�lt#>���=�,>��v?�~M?*)�>�m�=6�8�e�.��IF�9R�<��C���>��a?Z�L?�8b>yk���C2��� ��ͽ�0�c��3�@���+��$߽�5>��=>)�>H�D���Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ua~����7�d��=��7?�0� �z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�O�B���1=7M�>Μk?�s?�Po���g�B>��?"������L��f?�
@u@a�^?*�/�7��·־]n��t=���=��&>b��á >��X������������=mT�>�/->��>=4�>J��>O��>ӻ���~-�A�������6dE�gG�����:}����n� �~^��إ������'	V����c`'�7���>�������=P�T?�O?�p?��?:�����>������<���nh=S�~>�71?��L?{(?'�=�D����c�v��"⥾_����>�*L>�R�>1��>rg�>&y:e)I>_D>V��>��=�w6="�[:��=CSK>�ç>�a�>�J�>_N=Dɾ>�驿-�����u��=���H�9�{?��|>�������◃�@Ⱦ�O���m?�+<��ȿ&�οn�˿n~+?NE��O&��9��-?>i�H?y�@?�
�=z�O�(�� e�>���jζ�H��>�K���O�ݨ�>H�>��_>��:>�+�>��H��b/�(�3��Lپ��"??Vy�����tB?��5a��վ
��>�&�>¹�o����3���#�8�^G���D?`�6?�=���Z���-6����>�����={�=���=ET��������>��#>�S�>t;?�^7>�>H,�>����!��>�>�S>�I�>��C?=�>��=C�E��M���0�=��=�O�>�`>>[͔>����&�<�!�>�%>Vx����K=7f�y*=���!>��;��J���Nƽ��>n���>��=��K��T��q>�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾTh�>qx�zZ�������u���#=W��>�8H?�V����O�i>��v
?�?�^�ީ����ȿ)|v����>P�?���?[�m��A���@�t��>5��?�gY?�oi>�g۾E`Z����>ͻ@?�R?�>�9�&�'�w�?�޶?د�?�0L>��?��^?��>'Y=��9��嬿\탿�/�;��=�m>�N:٢��`C'�@玿�χ�^�f�N �]X`>��+=���>�y����B�k=�1���_��E�N�Mֺ>&�>�*I>��n>{��>�z�>�M�>�<�<ٙ˽��}�_�r��@?��?gG$�k�|�ڏ�=C�<�J��|��>��7?h�꽟džS��>��`?W�[?�:?@W�>���qٞ�p��A=��LN<��(>o�?�|�>U���w>�~ξM�S���3>Oָ>�Q=�1�nƀ���Ƚ茓>��?a�>0�W=�g?�?�(j>F�>�.P����M:'�c��>�Ϣ>C�8?N�c?CF�>�q��_�.�2f��q9��!kK���T>{�s?V3?���>@L��梿߶���o=r=ʽO��?Y�f?�t7��A?�.�?��-?%/0?�qe>'��<C�ܾj�d��>%�"?� �=�����0�%���̀�>�L�>>DR?���=�{��Ez�	?�g�*�'�[>��N?�?�o�ٗ4���������vM=>��O}��5�A>��=�>�t�E�'>v�½�&�=Ӳܽ�t�E|�='��=�^�>�I�9�Ҥ;����<,?l�G�QӃ���=��r��tD���>�1L>��m�^?Ec=�$�{����w���U����?���?xi�?����ߙh�=?5�?w?�&�>�Q��n�޾3�ྕVw��Ix�Nz���>���>_�k��+��������C����Ž���4
�>�B�>��?|�
?�d�=·�>����/��f�����f��-�H4!���*����w���826�)]�sɵ��Zl�VT�>��G���>��>�9>�#c>��>JB3=�σ>W>8�>��>�oP>�!>��=4;|�R��=R?Q���5�'�W��Z��aSB?��d?��>��d��s��֏�Vw?�V�?�w�?�v>a�h��*��?,k�>����4
?9=����G�<l��������������>�}׽��9�C�L���e�Ih
?q?����$�̾�׽Ҋ���l=`��?�2?i1���R���W�{�U��
Z�HP�=kv��8����q��������	{���L2x=j%?9Y�?�����J����e��B��>�T�>lJ�>���>�>�:پ���E�d�A�%�:���,��>2Lx?䄒>�5?�[;?5�U?�/K?�>���>{^ھF�>O3=���>�?$%?x�;?�0?�>�> ?B��>B�r�s�9S��f�
?A?1�#?�C�>�-�>��u��[;��f��T*������1�����b��;��K��(�%<�2�>XI?�_���a4�����P�m>�3?���>��>��}�0���+�<��>ئ�>p��>���k�a�.��>�n�?�8�A)=	�>��==R<%��(L�=�l4���=�����L�9�P<�ޮ= ��=NU���X���<ƚ<���&��>\H?Th�>7;�>�ʇ��� �Z��"�=g�S>x�X>6>ڍپ4��d��8ig���r>ˏ?>ɳ?��l=���=��=�2���㽾;��<;;<i/?:`"?kU?0�?zA<?��$?&�>��u�����Pq����?kI*?K"�>�;�:���v����x	?v�>�
M�#�꽆N�+���5�V��4�=�����j�k夿�/���B<���Zڽ��?p��?-��=�<�g������!}��\W?4y�>�1�>��?�=�Πs��*��0�>	�?�gA?���>��;?g�?A�q?���>����/�����s	���e�=��3?(8�?1%�?o�I?ݠ�<	y�=k\�<J������F���8ؽ�P�����
ۢ>�>��>j'�>�J>�l-��W�O!���ż�H�>Չ�>;��=c��>�N�=#ܑ=��G?"��>�c����	���Lw�����s?6�?��&?2�=3���`D��� ��%�>D�?���?�$?s�<��U�=#6߼񑳾
���rG�>���>iB�>%��=jV=~�=m��>S��>_T*�h�<5� iռ X?u�A?1G�=�Oſ��p�Wgq�q1����<7���1�e�5���>^��+�=*̘��6�Ղ��H�W��$���l�� ��/✾$�y�l��>l#�=�^�=��=η<�мz�<k�K=�ڞ<
�=x�m�ʬ\<r�4�T-�ۑ��"��U�7<GG=%�ػ�=ɾF�|?�KG?��*?��D?��s>'�>1�,����>xu�K�?AM>��E�ه���:�����Z����ؾi�վnc��a���>�jF�FQ>0>��=�C�<=�=��z=&ʋ=c���"
 =��=�ھ=�B�=�'�=w�>R>�6w?V���
����4Q��Z罥�:?�8�>�{�=��ƾk@?�>>�2������{b��-?���?�T�?:�?(ti��d�>I���㎽�q�=C����=2>{��=T�2�T��>��J>���K��q����4�?��@��??�ዿ͢Ͽ4a/>��m>Lv�>@oN��8'�2ε�H臾cJ��<�-?>H9�������=uM��v����O������m�l>,�J=H�ؾ`�`�KoZ=��߼}�>=��f<��>���=#Q>���T��=�N;r;=�#>3ż@�ཕؠ;(��=q�K=ߧP>k�J>qI�>y�?k),?G,e?9��>Rh�
þLG��?��>�u>�E�>��=@>G\�>�24?�\:?�C?"�>�\�=G�>�Ĥ>%�)�&$f���۾��8�<w��? ��?�k�>�U=�~�E���SC��m��?*?e% ?�>���g��B<��|0��)⽌��=)�>
Z��0A<������꽩鹽���=vH�>���>��>o��>J��>&�>w��>}�v>LW=y�>��=�,:<_�B��&����vRk�F}���r0��VH=x���=5`
>G�G�����퐔=��={��>��>Y��>cڗ=t8��U*/>�:�L�kc�=�a��Q#B��d��~���.��}6�;lB>��W>>-!����?3Z>�!@>dw�?2�t?z>di�=�վ����ve�ڎT�-ֹ=�	>�<��{;��e`�]�M�{�Ѿ���>g�O>�i�>nF�>I��]�.�O��<>���8��`:?`v��jl=��3��,I����\)��A�9��D=H�D?&ez�z�����?��^?���?R@�>tqG=�������0�u�=sg+�`~��f*�=%��>>K+?��>Qmھ^(��'̾������>.�H�P�������0��� �\緾�α>������о3��c��������B�.Br�<�>q�O?��?D1b�@Y���WO�������#Z?�eg?1!�>
M?�A?E��}@�GZ����=��n?��?�1�?SL>�@�>�x=���>%�?e�?���? !�?�^�v
�>=0����>��?'�>�i9?g������6_?F�o?��2?#J�֥ؾ�2�f!���9C�TkY>��`>>bZ�>`>>p�=�m��	���>G��>�"�=t��>c�d>�C�>���b�F��H�?CR�>:E�>o�\?�ӛ>A�>P��OA�>���>6���J��=���<�tȾs|�>�>�?�>;�T>̛r>�̿���?G�*>X���|?~{��uT�>
��>rO=ז�>�H>Q�>�`�>��>C��>/:>�B�>I�%>
)Ӿ��>f���B!�5)C�v�R���Ѿ�hz>���ԝ%�F��,0��*_I�B`��9W��-j�8"��3=�kt�<b;�?����w�k���)����}?�Z�>��5?#܌�����3�>���>���>B��.���vÍ��J�;�?k��?.=c>j�>��W?g�?��1�93�AtZ�D�u��'A��e���`�፿Ӝ���
�m��#�_?��x?ZxA?�_�<|9z>���?�%��я��(�>�/�4';��'<=T*�>�&���`���Ӿ��þ=7�RBF>��o?�$�?�Y?LQV���^��T(>��9?Y1??�t?��1?f�:?�&�8�#?k/2>�?�5?{�4?1�/?˶
?��.>i}�=7�Ժ��;=����I���Aѽ�Rɽ�N���6=��y=�\:x̭;D==��<�$��Ԙ���[���ּN8�<�.1=Cg�=_>�=�̧>�[?_\�>�>��8?��:c5�S����.??!F=�R������m؝���m�=�Dg?sݩ?��Y?�rc>c4@�=h@��	>mW�>LD+>xV>t��>�+۽&�I� Cl=e>�V>[�=��|���}���
ލ���<ˮ>���>�=z>��p��t2>�-����M�?@�>�i9�'���J%�D�-�v����0�>�oC?�I?`�<�Jվh&Ѽ�BS��{?�C?LUW?��n?[��0��KMH�~�D����ʜ>p��<z��8E������ HL�b��=�Q�>{����s����>����K��p�U��Wb���%�k�='����"~=�G*�7.��������oW+>l:'�6�C�7팿襎�P=?H� =Ó���Xu�����>���<L�.>�[>�A�=��h��ѧ���>���>�l�>s��<?�b�'�Q�T�Z�~>�y>?�?S?@�?W�|��Xw��*F�J�ݾp]��h�j=��?_Z�>�?/�>�^�=��վ\	��<f�*1:����>
��>�y�ԽG�>�����ܾ�"��~M>��?��F>�;�>�D?�-?(�W?�s?��?�g>�׽@����?��u?�j=@),��b�eb$�#B�Wլ>�//?蟚�<M�<}2�>�?)l	?(_L?���>�:�����ڕ$���p>��>�	]������8D>E�o?���>�_
?�g�?CӼ��%�4���X9�$�q>��>>Փ3?���>л?P��>/J�>~L��">xt�>&�n?JNn??�\̾���>!�>��0?Z��>t��>��!?�>�E6?��?D�?~,?����P.=>H��U���꽽zbL�=�5�<5E����=���;F^���< A��#����S�����*����=	��>bU>�����ab>h���[���W">�~X<�����G���H��C>�t>-�>�8�>��E�s�=6�>.6�>�h"���?���>��?�̖=��_�NZ���	U�3?,>�WC?�Hg>V�`����{8u�g�J�Z?�Pq?~�u�Vb���b?&�]?�b�=���þԲb��{�O?��
?Z�G��Գ>:�~?��q?��>��e�P2n����@b�b�j�ɶ=hq�>�[���d��>�>Ӣ7?sS�>~�b>qc�=�}۾̼w�Ht��>?��?���?��?�"*>^�n��-�������W?�!�>V!��M�?ZT ���̾.P��W����Hپ����sԶ�~᛾EP��0�.���kĽM��=%?�t?��s?�`?�����d��z^��~�ɞX��������D�3F�C�G���p�������䜾�FD=�b�<OV�[�?3<?���n�?l4}�#$ʾ����c�>5|�i����>.]'�r����2<��0�L�
���?R��>��]>_8?�5��4;��~�k�B�a��&�>/�g>��S>�Y?	N�;ۢm���������n��������\o>��a?g�G?7k?���,�1�+u���'���\Ȥ�!1,>.��=�b�>9�K��
�v�)��?�0s�}��lK������]]=��.?i��>�ˠ>|��?� ?M��䪾�m��.���<�Ż>af?n��>k#�>ƾ���"��>=�l?s��>Z�>l~��CX!���{��P˽�C�>��>Z�>!3p>��,�^�[��a���j���9��7�=�h?F���p�a�T:�>�R?<�:�;<�4�>��u��!�z�򾯮'�ӟ>��?���=(;>edž'�9�{�
����?p�0?����Kt�:=Hj?>� ?@Q���j?�H�>u����3ľA��>��f?�u?��?���>�����rG��􌽙��n��6Ch>J[�>1���E>�5=��E�[%N�߁!>+��>�.��Z�����Z�N�=��#>�����pf=S��[e�����Qo�����J$��6��o����}�� �d�WᅾoT���R�>D�m?�b��l�9�@r�@�V��~�c̷�G���K�'�U�Z>�5������7�$?��Bཆ���&��D$��\e����f�:�'?����ӽǿٰ���:ܾ! ?�A ?=�y?��#�"���8�� >�B�<�,��A�뾮�����οI�����^?i��>��/�����>ۥ�>��X>vHq>����螾�5�<��?)�-?���>юr�$�ɿ`���Ť<���?*�@xz1?�iD�!�� վ><8?�3?J�Y>�%��:=(���;�w?rӍ?��i?��K���^��6�*�d?� �>����_���1>S(F�t�����><(s>��v>�ƽ���7씽>/�<�,S>
CB=w�.�����_>XUr>G~��Y��=1Մ?{\�vf���/��T���T>��T?+�>�:�=��,?[7H�K}Ͽ��\��*a?�0�?��?�(?Eۿ��ؚ>��ܾf�M?bD6?��>�d&��t����=�3��}��m���&V����=V��>]�>Z�,����O�H��*��=%$�˚���|�v0��:�=-ڽ�-�:V�<��㼍�^<;©��:����۱�7vg�;6��=���>Ϭ>z5�> ֈ?��J?Y0�>���>�νfч��Ӿv����־s���x �rT�n3�L��w�¾��"���!��f�K\�"l9��?)>P�M��o���^��@r�;^u����>wn>B<��췀�S���-�׾Ý�^v��I���\K�~h�N�>�ȹ�?�D?������\�v�/�AQ�=�Bھ!}�?���=�#��Ͼ���=�� >�D�>�:(?���>6L����O���u���3?�z?�x����r�=��>"��gc>?	?��>hX��>-�%?~���7c��r~>'�?�Ζ>�Y>-��>�1��(���??.c/?;���*��b���:����Ľ�"$>R���窔=P�aR>E������c�%�/=�QY>:W?��>z�)�n9��	��o����G=�	x?�?�2�>;\j?#C?��<���Z�R���	���=%�V?+Sh?��>��x�(о�Ϩ�16?�.e?Z{K>ȫa��辐L.����e?�n?��?򶴼��z�3
��C����5?�v?�o^��q��q���V��=�>Z�>���>~�9��h�>��>?��"�F�������W4����?#�@)��?JH<<n�&��=S6?�O�>�O�,8ƾ���Ux��4�q= �>p���cv�;��O,��8?ߟ�?o��>C�����x!�=q��Qk�?�5�?z���l �>��žT��\�!�g��=�y�>ٗ���*�>ߊ)�4A|��'��AX��k~�=6t�=F��>��@����x�>�f׼�{��翿��,e���l��Ϋ>���>?cw=��i�.佾8�����[�X���'�
��>��1>g��@=����y�F1�z6����>�1��^�>h։�f㯾�l���Em�	��>���>�>�q�Y������?
̾�t��7Р�S�X�b?�Ҍ?�t?��5?3z��	ڇ�p,��ջ���??0�]?(n?nL�u�3��5)�&�j?m_��EU`���4�@HE��U>�"3?�B�>+�-�Ŵ|=d>���>�f>�#/�m�Ŀjٶ�����D��?ۉ�?�o꾤��>k��?�s+?�i�8���[����*���+��<A?�2>����!�0=�VҒ���
?(~0?%{�C.��l_?�`�h�o���,��Pʽ�ڞ>v�1��yU�~����b ���e��ۚ�JAw����?��?�u�?�� ���"��&%?���>�ė��sþ;�=xТ>uڶ>9@>�(K�]|>����e;��8>k�?&��?V�?`���֦�->!�~?@,�>���?���=�,�>�o�=�ݰ�^�(���#>���=�>�	�?��M?���>��=Yn8���.��$F�BR����
�C��և>�a?�_L?(b>~׹���0�(� �_�νQ�0�,�漼Y@��h,�cr�]�4>b�=>��>+�D�ZӾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��0a~����m7�;��=��7?�0�1�z>���>/�=�nv�ػ��Q�s����>�B�?�{�?��>�l?��o�>�B���1=MM�>לk?�s?�<o�y�'�B>��?������L��f?�
@wu@Y�^?!
�ٿ/���>���8 ��"�=��=)5>Y�սK�=7�Z=-t����~(�=�E�>��i>��p>�iK>�>>�q3>@����� �4��=����C�t���&��<R�ƈ�R�m�</�9(��C�ǾX]��.��<��ќ_�EN%��]N���=�R?�lJ?��h?��>����0�=����jT�=3����=�	w>/�0?I3L?/?w��<�2����d�N�z��c���$���~�>P�3>,W�>c'�>�>���QqP>��F>X�>9e�=�N\=Or�:��<��^>��>�L�>VJ�>}��=���>����r���SVP�����R`޾���?������R�s��'n��%����A>(T?#['>����q�ͿPl���6?E�*����h$����>7�?��Y?>\�>�Lɾ����]�>��p���"�4�=���<w�ܾ�v|>�ml>�Q�����>'����7���6�?�*���꾼?���=R��l�^�X�޶��w<fp�>K�JO����~Ǐ�������ua)?�T�>z#	���U�b�C=@H����=XA>�b�=@�	>į�=y�Ͻ~%�<�7���h>{�i>�ja>h@?8�1>[�=���>�s���_���>W��>��*�ڗ?�r�>8�'>�듾e�ɾ�'��:��=X��>��=�Y>s�%��=ੴ>��=�a\��h=�`�D"�U>9� �\ b���=����?�*�L��]P>��u�#�0�r=�~?{���㈿;뾅f���lD?�*?��=e�F<z�"�J ��;H���?X�@!m�?��	��V��?�@�?������=}�>�׫>�ξ��L���?&�Ž Ǣ�h�	��(#�SS�?��?��/�Iʋ�fl�
7>%_%?u�ӾOh�>zx��Z�������u�n�#=O��>�8H?�V����O�h>��v
?�?�^�ߩ����ȿ4|v����>W�?���?g�m��A���@����>:��?�gY?ooi>�g۾9`Z����>ѻ@?�R?�>�9�|�'���?�޶?֯�?Y�3>�`�?�Di?�Y�>�J̽�0�]��|��l�>���<�DM>>�q=���9Z6��ފ�܋�� s���DzT>�&=%��>NQн��j��=槀�3款(�I����>ڙ_>��*>�'�>���>5<�>T��>H��<ܳ�1Th����/�J?ei�?H���o�)s�<�=L�\��J ?.[5?O�ջ�JҾH`�>�<[?�Ѐ?2OZ?���>ck�@N��^=���1��d��<?cC>���>]
�>�}���@S>�PԾ��E���>���>�7̼�ؾ�+|��+��˚>m�"?�@�>�n�= � ?)�#?o�j>M#�>APE�(��=�E����>k
�>�l?z~?��?>����`3�lג�С��e[��M>?�x??6?�ԕ>�k�������Q��D�;����q�?�g?w�轟�? �?3??��A?��e>����ؾ���ǀ>(?y�3=A'��D��_پH?��)?�*?5�Y=b�ʾ��n=��뾪�&��;�>��)?��,?
ھ�p/��cP��*����ռ?����8	�=�O@>N�f>Ǚｏ<�=��=p>���jc˼u�=�8P=��/>��>Go�e��5=,?ʾG�)ۃ�K�=�r��wD���>RJL>7��	�^?~k=��{�����x���U�� �?���?k�?�
��؝h�m$=?��?�?�!�>7J���}޾���Ow��x�+w���>o��>ԡl�F�׏������IF����Ž����>s"�>�'	?-��>��B>��>���R'�u���k��
�S��*�7��'��f��N��x���F�d����ii��֐>l���a��>��
?T�g>���>���>�I鼷��>�fT>h>�a�>ppQ>�#?>M��=!�L<BM���FR?����s�'�%��D����%B?�^d?��>CYh�À������t?y�?	h�?6Dv>�sh� +�g?K2�>����n
?/�9=��ߊ<5G��������$��Û�>B׽�
:�n M�zf�i
?r,?�t��v�̾�&׽�H��ٹt=8��?	�(?�D)���R�T�o���U���S�l�#��g�=���	�$�^�p�2]�������烿�(� :=\e*?�^�?v�jN�|᭾�j�$�>��9c>Y��>��>fs�>��C>���41��5]�g '����U�>/�{?Eϊ>�R>?ݞ6?�.N?�KL?J��>��>Cyž���>~�<1w�>6��>	�:?��3?�0?�z?Hr3?�b�>��ƽ�����Ӿ��?c ?�6?Vu�>�c
?��t�č��8\�����j�����޽W(h=i�=�������0�=�X>Y�?���;7�����'�m>5�6?X��>���>�����}���<F�>j�?���>j� ���o�wC	��_�>׹�?��	��T
=�M)>l~�=wh���ʃ����=���W�=�#�XD��_+<��="��=�����|��/=;��;��<���>|�?�z�>Pe�>���ƚ �٣�e(�=��X>�S>->"پ�y��e����g�*Dy>ws�?�t�?p�f='�=���=����n`��)��}���Y�<��??#?�MT?䈒?�=?�^#?��>���E��OO��>����?҈(?�L�>�
��ľ<Z��N45��.?*?4`��[	���&��]ľl�ҽ��>��%�!�~��孿�ZC�y�C������d�?��?ƽ�a�5�:{߾6N��GⶾO�E?�v�>�է>4��>@*�4�e��m��,P>��>�R?���>��D?�\{?��_?�Ѐ>�)�+��xH��5�^���8>�A?U��?=��?=�v?g��>���=7��cɾh���F�4��wý�q��%��<�t>�Y�>���>]��>��=��ؽ�h��A����eU=�J>?��>�n�>���>�Jg>�BB<P`F? ��>\Z��\������u��ϼ���q??��?�=!?y�N=�Q�E�������>�~�?��?�&?ۺP�]��=Km�L��5�N� O�>�>3/�>�C�=�6N=ef>��>H�>�%� �:8��J�F�?��<?X�=]�ſ�p�$�r��뗾�j9<�X���ug��	��6�U���=&x������~����Y��|���j��/.��E���@Yz�k��>�Յ=!�=D��=Œ�<��̼1��<��C=^τ<��=IIv���,<�V>��U�������}��T0<�}I=�Ż��Ⱦ��|?yH?au'?b�@?n�~>1#>�I�z<�>�H���6?�QS>;Ch�4����4�\��쏔���վپ��e��잾�`>��H���>�5.>z��=Q|�<`R�=��=�(�=��8Z^%=]�=L
�=L�=V��=�>>!�>�6w?T�������4Q�:Z罣�:?�8�>�{�=��ƾn@?v�>>�2������{b��-?���?�T�?;�?/ti��d�>?���㎽vq�=#����=2>d��=Z�2�S��>��J>���K������4�?��@��??�ዿ΢Ͽ:a/>s>>��c>�O#��A�v�����ݽ���:�U'?Q���:���>��=AM�����+��=���>Nbe<�9�u`� �v��͛�
�k<K��=o�>.u�=׌�=��x�&r=>�>�R�=q��>�0�<�(ҽ�1<���=��=��C>^��=T��>ַ?ǣ)?�e?VB�>�J�9þ��ƾݓ_>�9�=	�>���= N>��>.?p6?rP?��>~�[=��>�`�>o�0��4o�,!¾!j��/�<ڻ�?���?Rë>�j��9�����<���H��?�z0?$,�>�
�>6��i���G'�U�.�����N���u,=�oo��{M��_���W���ὃ&�=m۩>���>Rc�>�Fy>r�;>�]P>�w�>[>���<Q8�=@���<�G��V��=����W��<SJļ���5c���'#�����~}7;�,�;kGR<`;�;��=�g�>J@>���>��=g����0>�L��I�L���=������@��:d�X-~��}.��Y5�@�C>(OX>ˁ���ב�?!*X>�{:>$��?��t?��>I��hvԾ�h����c�R�|�=��>n�:��:�$�_�V�M��oѾ4p�>��=��?��>���g9-�y;s�&��k"8���?�J�a =$�ȼ�R�= ��u2��=�6�)/-��~Q?�,�������?`�Q?8Ā?R�3?�ؽ��m�Iw�<�,����>(��f(P�;i6��<?���>�c?!�����U��D̾����߷>�3I���O������0��8�[ӷ����>�����о�#3�Sg��R����B�nCr��>ǴO?��?w9b�'V���SO�V��7���p?zg?��>�J?�>?'��pw�t���e�=!�n?���?x;�?�>q2A>���c�>Y�&?�d�?�-�?��<?��D)>eΐ=".�>N��>r�>�Z�>�ֽ�̉=L?�P?~��>�K��*��W������V��X�#}W>��/>:��>\"�={�2=��;������>��>1��>�F�>��>���>����QF��w?3��>��z>�/?�=�jx=��(��u>u=6>�<p������������<>PL>�|`>!4�=\�W=�ֿ���?�̉>S븾.^?���z��X�=�T5=C=>��>M�g>��>>�k�<��:>��>�5 ?\<#=��ؾ��>1	�P���=�TW�#Oپ4g�>C_��b�G�����
��$T�i��Y��{l�E�����=�������?+���sg��)��?�gW?뀢>�s/?�Ԕ��"���>{��>��>��������7c��Y���?�p�?<�c>��>��W?^�?S�0�W�2�OZ�͚u�_&A���d���`��Í�\����
�������_?F�x?�zA?Z��<z>ؤ�?a�%����Zf�>�/��%;�D�>=\�>p����`�liӾ�þ�]���F>�to?�?�&?�IV�ٱ8���%>��8?��+?\Lp?#�0?�>?ߡF���?�DL>��?�g?L#;?�8?f�?�%<>)>�>:=Pjq=��������۽5�ݽZ�U�\~%=��=b�ԡ�<BQ�=2r<��G��%���;u@�����<}�=H�=$?	>o��>0j\?���>.1�>C�9?�x��4�G���Gb+?V�U=Rှ_R���^���ﾂ�=M�i?��?vRW?\�f>��C�$�A�[�#>T`�>K>!�V>(��>|����?����=�'	>�>�#�=��:�q�������/����<Nn%>]��>�c>��/:�E`>�������9ã=��8=U��@h����<���՟F����>ql?�{�>�1L�Vm��p�?eo�/��>0�,?L�Y?�Nk?�d����>�����r���=ZI?�<�=5�=��	i���+U��S�> ڰ>��s��H���>�����L�����l�V���>��n�H�>�^����۾�E�>R��>L�w���j�ȕ���$����;?��>~G������=�ž�h>�q>���>[�Fl�A�T�7�����>t� ?m�j>���>��]�Wo��]��>�1?D?g?�?�$��y�,FJ�mWN�@F#��<�?�`*>�q�>���=��>�-
���'���I��t3��`�>պ�>���ǗC�cl���Q��������>ʌ>�	>B2�>wH*?�S?-�U?���>\��>�h>�X�����O#?]N?�,m=&Tٽ��{���1�C�;�o�>o�>d���b>1��>=?�;?[�H?_��>D�<=����8>����>��>�?V����Kh>$#J?2>�>yp6?��{?�l=%��Ga��!��3s=�xI=0�C?��!?��?���>�Z�>ˁξ,\���q>�8w?L�?��?9�->7S?��>�R�>Mu9=��.��H�>iN�>�@?'�?���?�Z?���<7�b�N����OǼ�ep��D׽L�����=w;���EٽΊw�tU�Z�=�#�;���2�3������=�b�>Xt>?ו���0>��ľ?P���@>����A������V~:�	�=/��>��?��>�#�Ӑ�=[m�>���>���a(?��?A�?q?8;�kb�}fھl�K���>g�A?���= �l��w����u��d=��m?R�^?��W����0�b?+�]?[�:=���þ�b���}�O?��
?j�G��γ>�~?��q?T��>p�e��=n�����Jb�M�j�>۶=�v�>Y�k�d�56�>��7?TO�>$�b>���=�s۾��w��q��Y?��?��?���?�4*>��n�#/�1������V?�>UI���(?��㼑�¾Y���a���_޾J���c���Ҩ�i�����@��=�����bC�=]�?z�x?`�v?�_?�����Ik�T�_�\���Y�Pa�hE���?��N�#�A�ũr��t����v���m�<2
U�IN����?n+?2Ů�J��>\���iڪ��Ⱦrw�>����8N	�hY@>Z?���8=��6>��1�j`]�h��CE?k�>���>�B?;�[�<�T�#�A�l�:����A�F>_~�>��>�d?h/<t@����tOξ����R�l�L1t>�a?\I?k�o?����U)3�zၿ�f�ׯ��sb���HC>Z��=ߋ�>��U�������(��A�8q����	���b	�{��=L�7?�΁>|َ>�0�?�?�*�|#���<c�r�+����<�l�>g�c?�,�>[�>1OŽ�����>��l?���>�)�>���C!��{���ɽ���>�f�>Ջ�>:�o>i,��\��?��r_��k9��E�=�Dh?gu���a�-A�>HR?d�d:%jK<�B�>�{���!�����\(�h�>��?թ=�[:>�$žx���{��Ӊ� )?p�?�u����(��S}>�� ?�M�>��>��?׷�>����9s?�^?��I?�>?R��>O�1=�9����ƽ�2(�*�1=Rŋ>�V\>�=p�=MP�G�Z��#�Y�R=P�=�q��\���?><솾�<��;j 	= t6>��ο��a���ԛY�[RS����m�T��=�Zy<K��=]���ɮ�H�h�V��s��ӊ����l��>��I����a�?��?��G`���F���؏��!�e+�>o�����)':��ܒ=A\��O��~���Hy��e��?N��.�O�'?�����ǿ񰡿�:ܾ0! ?�A ?7�y?��9�"���8�� >BC�<.-����뾬����οG�����^?���>��/��n��>᥂>�X>�Hq>����螾P1�<��?5�-?��>Ҏr�0�ɿ`����¤<���?/�@�=?���I�ɾ�_
>�&�>
?_OF>�e��;���<��j��>ȣ�?A�?=7�=��Y�o����.`?\�<A.8�����^�=���<'�m=m�&��3>qZ�>�Y��zX��Ū��\�>��>~��J��m.�Ub�<v�>Sz콁��4Մ?,{\��f���/��T��U>��T? +�>u:�=��,?W7H�_}Ͽ�\��*a?�0�?���?(�(?2ۿ��ؚ>��ܾ��M?^D6?���>�d&��t�ą�=K6�`���w���&V�Y��=Y��>o�>��,�����O��I��M��=�����ʿ�C�#a;��� =�a�</X����'����=�4;=s���� ��1���6<�mb>��>���>-��>�fP>��L?[�??!�>�4�=��$�u������)=��"��䤽gk���d��`E����+�߾O�;���	��KѾ)�;�t��=JO�1&��*(�)�d�� J��#.?��>Xɾ�M���"���ξ����1�$\�EIѾ��3���n�an�?+JB?���/_R�J����;�ҽ���Y?���a
�@M��{y�=�}��w3=�W�>�J�=��⾺	5�Q�T��&?5z#?�Ww�i�PJO>�]�]�?�?|#?��>�J{�ʮ�>�Y�>@ԙ��5U��l�>`�_>�=���>�s�T����
f���3?�Si?N�1=�[>������Ѿ�V�9$>�Q3>½U|�=L�>�W�񃛾Tu�T �E]�=�|T?/�>�*���������2��<�=�	w?L+?���>�Li?��>?cϚ�Y���H�\��>�m�=j�X?��o?{	>����Wʾ8塾%r7?�a?�>m$b�-�Ѿy�)��Q�`A?�xj?�s?P��Zu�8T��a���8?R�u?X^�jM������EO�*֪>�9�>���>Mv6�(ٳ>�x>?���mP��}4��^4��ܞ?�z@��?{��<)��"�=ӛ ?���>��Q�?�ľ
���2���$�=���>݉���Eu�����s$���8?}�?/@�>�w���e�X�M>"ն�R��?2�?=�v�ň>(^��<C���#�9x�>��<0��>���>8����t)��R߽Ů��'�����<���>�@�넾�<�>*'��(k����I蝿!Aƾ�q��R�?Ի�>� ��1˾]�>��׎���:���z�A����>2o>w�����X�{��;�k}��	$�>uN���>�!V���� ���.p<�(�>�,�>骃>�b��松��P�?�u����Ϳ}О�K��+Y?��?Ä?�?8g:<�0{�Cz�u��R�F?̗q?h|Z?~>�^<_�Q�>��j?�_��pU`���4��GE��U>g#3?'C�>n�-��|=q>=��>_d>�#/���Ŀ5ٶ�����I��?���?Ko꾲��>9��?As+?�h��7���\��g�*�x�)��<A?32>t����!�
0=��ђ���
?3~0?�}��-�]�_?+�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?ҵ�� #�g6%?�>c����8Ǿ��<���>�(�>*N>bH_���u>����:�i	>���?�~�?Qj?���� ����U>	�}?�>^��?�P�=П�>5�=H��0;��#>B~�=�1@�Ð?C2M?���>G��=�F7�:/��kF���Q�3���C��v�>�b?��L?�tb>����<�3�� �#�Ͻު/����� ?�C %��Z�J�3>t2=>� >OE�~8Ҿ��?Rp� �ؿ�i��(o'��54?
��>�?���C�t�����;_?�y�>7�,���%��WA�c��?�G�?%�?��׾ V̼l>c�>�I�>ս���������7> �B?5��D��T�o�V�>���?��@�ծ?�i��	?_ �dP��4^~��}�^�6�<��=��7?t+�F�z>i��>��=umv�l���m�s�B��>�B�?�z�?3��>��l?�o���B���1=�H�>}�k?iu?��o��(�B>��?b��x����J�� f?��
@�t@D�^?f��P�6���! �6��$�=�c�=�#�>���Ė
=�e>Xz�=65��p�<���>��>3X>D �>�{n>���>�	���(��E��������q�ݾ�vϾT���Z�u��������֎�h�U<>�=�i̽�o,�� ӽ�Yb�V�>�6S?�S?�?q?� ?�8r�O(	>��!�.=�����T=�,�>��8?�kF?Sf$?El~==�����_��~���ԁ��E.�>�.P>(��>A��>�߱>��{���?>KSI>���>;�=?9�=�޻��=��=>�ت>/��>��>Y�%>8��>o��;A��B��F�����X��?j�z�q�or��(�Ǿ�a��ڹμ��?�N�����|�п���	/ ?��f��I*�c��Q
n>%>?<ib?^��:V3��$��BGz=�����ν�f#��k�>�o�!�ܾy>��?e�W>�|??2�0c*���3���(�`�.�`5-?Pcw�f��������{����2�I�X[�>r9���7D������P��v�.��-���
?�W�>b~>�m��~�k&����>:I>=�C>!i�<���<C*(=��@>�<�SR����>�D�>��?��5>ޏ=�Ʀ>�v����?�xK�>�.>�8$>��:?��%?�̼�����By�=��p�k>͔�>��>�>�bF��6�=���>"s>�Θ�`�t��^��D4��dM>B���U�0HH��3�=�F��w��=�Ӟ=�~����>�
pN=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�z�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?ܵI>Z�?C�s?c0�>��s�],/������9����y=b�p;��>'4>pe��EF��s��k)���Oj�E���)`>��$=��>8������� �=��ɧ��&h�J�>5vn>2J>��>D?W��>7Y�>��=MJ�������-��S)A?r�?����#cf�J�ν��ܼuȈ���?o� ?C%����X��=��K?/�y?�9^?M{f>ѝ1�������������|q�7pL>uɲ>��>�ST<`��>G�Ծ9L.��c>/��>_>^?ؾ�2㾅j~����>7;7?���>R��=�� ?��#?��j>+�>�[E��7��.�E���>%��>�F?��~?��?ɹ�[3�X��4塿�[��6N>��x?ZU?Ε>ݏ��
���4�F��I�"ƒ����?�lg?ta��?�2�?Ʌ??��A?%f>�}�!�׾S���=�>�c?����7��y(�r�+����>>�>�B�>�%��,�Q���8�$����UM??�Q?݇!?DO
�C	_���˾�<�g�Q`�$^,���M<4+>�9>/~��=?�=�h�=�|B���G�� ��j�=T�>�	>���g�K�+=,?��G��ۃ���=b�r�xD���>�IL>�����^?)l=���{�����x���	U�� �?���?Uk�?q��*�h��$=?�?S	?l"�>�J��~޾>��jPw��}x��w�e�>���>��l���9���ə���F����Ž@�
����>\��>>�?!A�>��7>һ�>&���R#���0�\�\��~���9�g%�̱�����Bh(��T�M����}�΍�>l�h���>Z�?��Y>Z�u>~�>%y#�.�>�@u> 8�>S��>J�8>�/><#>�;��ɽbKR?G�����'���辫����2B?�pd?F(�>Zi����������?���?Is�?�:v>E}h��*+�n?j=�>s��p
?�I:=����-�<*V��?��y5����>4׽�:�M��gf�{j
?/?mI����̾�6׽�����"j=}�?)�&?=X+�LR��+p�=;V��SR���~g�v���ʖ%���q��������`��H�'�v^+=ڹ*?Ꮙ?������C���9�l�'�?���\>C�>���>bT�>�eH>L��S�/���]��(�WA�����>��w?��>X�6?��2?-+_?�:??�6�>v��>������>�H=S�>*�?SR?^;+?!I?4��>�?�]>����f�߾��Ҿ�i�>��?�?4�?|�>��E�߽��3��;��j=w�{��r6=. 0=s�7�3¢�sG>��l=J�>��?;�G8�����X�v>ã9?s��>b��>N�����}���=���>��?���>����n����;��>$Ń?q� ��=z�+>���=�墨��޺���=|�伃��=C+M���C� Z<^�=���=�<m�<|�%9�D��ý�<�q�>u�??w�>�>�>�"��?� �������=}0Y>�S>F'>�9پa�� #��W�g�oey>�w�?�z�?�	h=W�=7l�=����Y������齾K�<�?�W#?6LT?䍒?��=?~a#?w�>�$��C��KQ��7��y�?m.?�ן>�����F��lO���=�J�>��?Y`t��������Ծ<�8�Z$>}��P���x��sB�����	��������?�W�?�i���;��]˾���Ԁ;��N?[�>Rٛ>7��>����K��> �5��=~L�>�LY?���>�l8?^
�?7�?)��>�>�-]}�Щ��C<�=$>��,?���?��?/X_?��>��>��L<(fþ��׾d����/�.Iʾ�7=��J>��<>6>�>��=��n>,#轨��=i�t�wǆ��l�>Y��>;>�K�>�=�����"G?�N�>���	L�̍���>��K.�)nt?���?](?�T�<�2�
�D�p����>��?��?��'?U�,I�=�
�S���t�Ǝ�>�{�>V�>R�=6O=�n>��>{�>��=���O:��"���?wGC?th�=8ƿ��q�]q�x�l�e<�����	e��J��ːZ����=w���q��H멾6�[�h����n��Mȵ��X���{{�c��>2o�=�Q�=�$�=���<=Xʼ�W�<�FL=���<%:= Yo�on<�7�C�λ�R����ZvS<{!G=����u˾�w}?�I?=s+?үC?RTy>��>7�1�j��>����l;?��U>&�R�����.o;��T���#��_ؾ>}׾��c��ß�H�>RH��><�2>"��=L �<ǧ�=w s=���=�xJ��S=���=O��=�p�=���=��>/;>1w?[���Ӳ���0Q�
�C�:?,c�>蒭=�^ƾu@?l�>>�)�� ���me�C#?���?�V�?��?�i�Ba�>������,�=�����42>�m�=&�2�=��>��J>����G��C����3�?v�@��??	܋���Ͽ}Z/>�Ey>:M�>�)�t*:��43���¾[YU��O?��辦,>�x&_����@���+d
��m��Z��>;������sS��Չ=H ������ B=.ް>��G>��>��J�\ÿ=�܎=�1N>-��>��7�l����f�(��=O=�=w�>��c>5��>�j?��.?lDd?%�>�h�ü˾S'ž�;�>;V�=�	�>�|�=<�K>/Q�>H'7?�A?�dI?E��>X�=G@�>%(�>'�-���o�<������<���?�7�?�>�C�;.�@�|��<���νY�?��1?��?�:�>T���QV��l�V {�=��=�h�==�V��o�X�&��p�����ȣ�c�>-2�>���>��>r�>DL�>�^�>��Y>�Sg>d�==�nG��f��'�����Z=�m�o�M����=��)P���C���>�[.=մ@=F����=`��>�?>o��>���=����-/>⭖���L�0��=#I���+B�U.d�CI~�9�.��Y6�d�B>.X>�����0����?��Y>�w?>B��?�8u?��>K ���վ�N��3e�/S�,�=s�>�=��t;��N`���M��uҾ�3�>�u�>a�>Ϲ>cB<�PeG�2���zپ��1���>���/�:mm�UI��3��o,��_�q�'��Y5?�ct��WA>���?W�Y?��?�ϓ>�Y�%b�跒=?j��Z�;������)y=��!?��?ö�>_���d��F̾���t߷>.?I�/�O�����J�0����̷����>�����о�#3�\g�������B�VKr���>m�O?��?�<b�W���TO�l�����ir?�|g?��>�I?�??�"��+{��s��am�=u�n?س�?�<�?�>��d>�Q���X�>��? �?��?��?�L�<Z�?�\=3�^>���=$�a�*�d��+��>�b?NR?�]v?����e�rD�7*Ѿ+ww��_!>�|>�>���>��>5�A>dͺ�'8��{�=.��>���>b>{�>P:�>�`��j�Y�r?+��>r�>��6?�%S>!�%�)fϽ��^>�/��߉�=���=�+��)��X�>f~@=���=��U>��&>��տ���?`��=C���s?:�'���M>�yo>04�>x����% ?f��>q�->�Wm>e�>���>J��>?�?-XӾ-B>����y!��LC�K}R��Ѿ?�z>�����%�(������I�瘵��T�k j��&���0=���<�C�?j��A�k� �)�����x?^H�>�6?�����B���>���>�͍>�������ɍ�/u���?s��?�Ec>�(�>r�W??�?�1��.3��iZ�ѝu�A��e���`�/፿�����
�N��C�_?��x?�gA?rI�<�+z>���?��%��ُ��6�>�/�u;��C<=%�>A����`�́Ӿ��þx��E>o�o?�+�?�J?�1V��%�>�j�>���>�@?�3?� ?�!? d��a?8�R>F��?@4=?0�?�n�?\��>}�9=�JS>ث�=�;>V?�����2'��8���?���p=q�X>"K>^�U����&Ƚ&��p+S�9���^��3*�<���;�.>!��=I(�>�]?���>��>�h7?�u�(8��:��:.?�8=�܂�Ϝ��8��C�򾖻>i?���?�X?Ԯ_>��@�T�D�,�>���>��(>B|Z>�;�>�x���J����==c>!>��=��O��~��r�	�����[�<��>���>|E�>�wB�z�*>�X���|�x6>>O�*��ٮ�c�C�B�C�m�5��sm���>sO?�c?��=�޾[�Ž��\���?7?$�Q?�}?3�=��پ0�2�W�J�����>�=�#�����E���v�2�|gp=�zX>�阾�ؾ�r�>p{��<�/�y��6l�ť3��5�>jN��DX=�(�^�^�s!]=G�?\�G���H��O��Cb���:2?H�E>7�վt��+�\��l)>��>ō�>���ȼ	-!���ž�e��?���>�������W�+�da��i�>��B?ݲ[?���?��z�f�q�ݦ=��2���᭾S�k��?�ڱ>Û?N,2>���=\R������`�(zB�޴�>�|�>�h�bG�f���8���e!���>�i?h>�?1wM?b�?�a?��-?�?년>|:��)��=�3?��r?�D�r���׾G�ky.��z����>�*�>g�F�&��>չ?%��>��?��g?.��>�;�ɤ��	�+��>���>VpO�H���U5>�Y?�g�>��R?d�?�ף��F:�6�ܾ�]��4g\>D�=E�#?�/?X0?k�>ņ�>�)F��z�=�4�>-�B?=]N?�r?7�r�3�^?�N >�7)?��I>��>7b=?]=�>�hJ?��?xV4?P�?��=b���,���ڽ�8�#b?�d3>Md=b0��%�b�>���1�;G�N�#������bѽdޖ��=�=��w��h�>��s>�y��2z2>�¾LJ���C>���P؝�/�����2�R�=��|>�� ?�L�>�B%�sC�=n��>_&�>�5��f&?y�?f�?��<�a��Cپ��G�>�>Z�@?��=eYi�ğ��yTu�fA]=�?l?+�]?r�W��b��s�b?��]?vl�[�<�+�þ��b�3N�z�O?��
? �G�Z�>Q�~?��q?��>�e�X'n����W#b���j���=iz�>�c���d���>u�7?�E�>�c>0;�={�۾n�w�<���b�?A��?���?y��?f�)>�n�Y%�������8[?���>j7��3�?�Ι��˾�툾�᏾�߾�L��?|�����=����D'�󲁾���(5�=��?�!n?YRv?��a?�o���|c�%c\��.���U�&s���l���A�sVB��O?�all������a���.=xvR�@B����?W�.?dCӽ"�%?�騾y���CTƾ`1�> ��<6���!k�>{5Y���Ƚ���>����R�<s��I?g��>���>��A?M�r�aKR�l�������]f>���=�
>��\>�5���Q������Rz���㾦v>�pc?K�K?��n?Li�v*1�ς���!��,0�dq����B>+}>:��>�W�]���4&��S>���r�Q��tp��S�	��~=��2?C#�>峜>oM�?��?�y	�{w���Ex��u1���<�*�>i?�J�>��>��Ͻ�� �|$�>jh?��>�r�>�{�v���p�X&Ľj��>��>sk?�~>�*�p_�f���凌���4�mk>�_h?ٱ��nm�m�>�S?�[�<�r(����>�E�.�#��
澴��XA>��
?�x=h7>�(��.���z�0ƀ�q--?r?{ԍ��/��?>�4?��7?O��Ǘ?|�>i����	a>�6?�Ig?�t?�&'?�*?l�?'9&<�b���,�͊���c>\ot>�ι=Pm�=, ?�4T8��4Y��>��`���<~R��=��żgrk��u��r`u>E���FV���ݾ��.����iL��ʙ��!�˽��ɽ����.���v��n ��!���,@[�deϽ�~�'��~��?�R�?wN)�n|��Be�����G�b���>�/���*�F���dx�j ��G�=}��[�зm��`6�4�W��e'?1���T�ǿ����d�۾i�?� ?��y?z���"�Ї8�� >��<?��
���@�ο(���-�^?^�>�m�O{���+�>4ł>�X>x%p>7��䫞���<��?^b-?���>�Er��^ɿdr��N0�<���?�@PK>?�F%���Ӿ:�q=��>��	?d:E>,�S����������>���?���?$��=��S��&l��a?T7���6�^�c�҇�=@�=Ta�<�'���5>+��>���C�~����M>��}>@Ӽ��ս�'U�׆�<:[o>�BŽ�/��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6��{���&V�}��=[��>c�>,������O��I��U��=�����ƿ�$�)���4=?�#�rlb�����LGS��A��s�n�mX�8�g=���=�O>s̅>�W>ec[>aW?d�k?��>˾>ot�鬉�9�;^��ᢂ�����$��<��s��O����޾�	�������=�ʾ]�j�D&(>��@��h���l������z��F?�?>t���G�Y�!u�H���i��bL�E��l㾑��Z�P�?�hU?c�h��.�߆ ��A����\��IY?�<u����B�K�J���i�C.>���>��i���
��^Q���U���H?��?���8���[%>�w�=<�>��?]i�>gq;����>	��>T`a��W�M�(>�>�=�P�>�t�>o:�<�۬���3�t�7?�6_?�	>1K��:�>��þ�y �>~�<CO�=*��<���=&	-���F����V&��N>W?J��>c�)��������}6A=%�x?@?�6�>�k?��B?�f�<#���ǇS���t=��W?i?��>AO���:о�x���|5?�Xe?D�N>cfg��X�"�.��<���?�xn?�[?�於 }����m���>6?��v?s^�xs�����L�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?��;<��S��=�;?l\�>��O��>ƾ�z������.�q=�"�>���~ev����R,�f�8?ݠ�?���>������4�3>d����?���?�"����:>���JJc��0��
��>��$=_��=�,�>.v��_*����Ɠ�}�����ʺ�	`>�r@�{����>i=�ݿ����R����%��X���i_>�
?	tý}���T%�|�z��I���h�cGM�q�>->Lgڽk�I�!�i�[#<��C1=���>�3)���>�(ٽz������z�����>�>9>��	����'�?4�Ӿ�oʿF읿���K?"��?�?��+?�������0���Mq��o�S?��t?�N??cս�2������j?0_��<U`���4�HE��U>#3?�B�>{�-���|=�>F��>�f>�#/�J�Ŀsٶ����Y��?�?�o�i��>U��?�s+?i�8���[��g�*��,��<A?2>d���߸!�}0=��Ғ���
?\~0?�{��-�\�_?*�a�N�p���-���ƽ�ۡ>�0��e\�CN�����Xe����@y����?N^�?g�?ܵ�� #�f6%?�>e����8Ǿ��<���>�(�>�)N>fH_���u>����:�i	>���?�~�?Qj?���� ����U>�}?�_�>���?��=څ�>np�=M���
0�Ha#>���=�~A�R^?�M?W��>�A�=��8�z�.��F��QR��	���C���>R(b?��L?��b>}���w4�!�
ν�<0�=��~�?���*��޽.4>�j>>�8>��E�̥Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�e��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?gQo���i�B>��?"������L��f?�
@u@a�^?*?�ῢॿ�;;EξsQ�=֧�=@y>d���:�=��3=e�p<�L�<���= D�>$|0>�?�>��>dQ>Z��>������(��#���I���I�Tp����L��N��򒾹[�����@ľ� ��P��ꏂ�ktнym�,��W��=��U?�R?Pp?�� ?�8x���>.����<={#����=}-�>�d2?�L?��*?*ݓ=����X�d�M]���?���Ň����>�lI>b{�>VD�>&�>�W9H�I>p#?>���> >�Z'=�=ߺ;\=��N>K�>l��>V�>5T��U�O>�U��ȥ����i�O�뾪�����?x}����:�"t��B����J�� �<c:H?�����ϖ�/�п�k����6? �����gi�=�f�>6?>�j?�8>�k��������x>�/�=4�M���˽2���<�;(����n>���>i�;>kȇ>B*?��b'���0��M��ѽ2>g�.?¿��CH���6]��L�}<�(�>W.�>򂏽��ߊ���z���Z�ldn��d?�V?.%ռ>cp����8y�I C>��>�«<f��=��\>)J@�(��*�F�E;%��L@>;O�>�{?�V)>�n=��>�x���P���>��>����A�5?�35?u�=�7��2��X
 �1>9>��>o��>\C>v�� =��>�7e>\���A1������l��=��p@2�)��=8r�=?�ս�9>��>�*���9��L�<�~?���(䈿��e���lD?S+?\ �=��F<��"�E ���H��F�?r�@m�?��	��V�@�?�@�?��K��=}�>׫>�ξ�L��?��Ž5Ǣ�ɔ	�+)#�iS�?��?��/�Zʋ�<l��6>�^%?��ӾOh�>zx��Z�������u�m�#=Q��>�8H?�V����O�e>��v
?�?�^�ߩ����ȿ5|v����>W�?���?h�m��A���@����>;��?�gY?ooi>�g۾:`Z����>һ@?�R?�>�9�~�'���?�޶?֯�?�I>a��?��s?�l�>��w��T/�/3�������m=ȧ^;,Y�>�p>#���VhF�%ԓ��b��{�j������a>P�$=\�>�p��7���I�=�틽KA��%�f�ܧ�>&q>f�I>�W�>E� ?/b�>ɣ�>8=�^���ހ�t���o�K?���?}��e;n�C�<�N�=�G^��?V4?�[��Ͼ�J�>��\? ��?��Z?�%�>����#��޿�ai��&4�<&�K>�#�>],�>#܈�uUK>��Ծ�1D�T�>�Ɨ>IX���ھ�H���S�� ?�>�U!?͈�>o�=�� ?��"?��h>>�>ΩC�s摿ND���>'��>�Y?�?� ?�
��N�3�<	���+���S[��(P>�qx?l?䛕>=����������]�T��G����?�Qf?�B��|?{�?�>?�B?��n>b�۾w3��o�}>S*?��>�N8��@�w�|�t�>���>��>	�T�����d=���N��s�kJ,?�D?�:�>��Qm�Fz�ڣ<N�<<Q=m+��.a<�̻>��->�e�n�!>ԙԻ�=�=�����i��S�Z����g�>�8�>�:�uc+�4=,?�G�4ۃ�`�=��r��wD��>�IL>��E�^?l=���{�����x��	U�� �?Ġ�?*k�?���&�h�E$=? �?�	?#�>rK��~޾!��.Qw�B|x��w���>+��>��l�
����������F��l�Ž�2"�I��>���>/�	?g��>��,>�N�>�ӄ��S(�t��ެ��VTS�]��,<�}''�$R��ꢾҦ�c%l��Y��.6��¬�>��v�v��>A=?��T>��j>�e�>^��<���>ETh>��>Zl�>:�A>]�@>��>�#<Q�d�UR?(K��.�'��k输����A?\cd?�-�>��l�yc��1~��:?R?�?�O�?��w>�Th��G+�:�?���>
���a
?��7=���c��<8���x~�t���L�I��>��׽�$:��)M�	ne�W
?X?J
���̾:�ֽ����oo=�D�?��(?��)�*�Q�$�o�5�W��S�f���h��b����$���p�9⏿�\���#��#�(�<	)=+�*?�?ؒ�Lz����
k�
�>��e>���>��>��>ݣI>��	���1�
^��6'����#T�>�E{?6h�>`�C?�:?^�K?Y�L?$ܐ>�D�>o���5)?J5�<t��>*��>��7?i�.?;�'?�(?PM/?�SQ>�ݵ�'���a�־��?Ԩ?\?�\�>�?܏�� ��a
��֣���g�<Di�|�=�,�:����W���)=�FZ>OS?^�ý��6���'S>Ȍ5?�K�>�A�>w!��K爾@�<,�>�$�>��>%��;,f����>V�o?m�����<�v9>-H�=��I�(I�<���=&q�A�=}���M�5h�;�|�=��<m��6b<��;=�{����� c�> �?�z�>�w�>҅�}� ��W��F�=�W>�US>	�>��ؾ�d���"��I�g��x>-T�?Br�?��h=	1�=���=�<��鑾����E���<�<��?��"?VT?���?58>?#~#?g>*$��!���1���@����?��+?M��>'��@ľ�פ�p�,���?�?�ic�hT�͘�ͷ˾�����=��(���z�1`����3������g�� ��/�?�Ϟ?�]�;E�:���پJC�����?E?�y�>g��>��>�0�>d��m�?�B>��>b�Y?��>�+?��?V?>?�L�>���㑿Z��{]=f݄>��?��?C�?R#g?�A�>��>������96�䤒��tL�=�����F�'�=��=>�l�>���>�qE>ˡ��X=Q���萼�'�>OW�>�!><T?���>�Po=�G?���>:E�����ۣ�ݱ��c����k?���?��*?��="V�Vd?���-�>g��?�ū?6-?]�S����=���𴾰 ��@�>6�>�R�>�T�=\=t\">:��>���>UI��q�p\8�9�d���?d4H? ��=�H_i�ƹ��ֆ��\��<oȚ��5����X�ҵa��o=���a��}Ь��8\����������������qo�-��>�h�=|�3>ѳ�=j��:Jo�9��<,��<�'׹N%�<�X�+R�<@8����;y�,��"��<���<[�r�7HҾV�z?K�3?��!?�8?VkQ>ٕ�=�.��~ϐ>�w�g�	?�4>�j��4Oƾ=3��������O���羊@\�������>֚���Q>;:A>+_�=�_�<i�>�=LCk='�ܼL�$=���=�@�=���=�|�=��>	�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?��>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>r��=v�2�T��>��J>���K��D����4�?��@��??�ዿТϿ6a/>�HC����>�HU������P�q���+W���?���'�S�m�>�^��8����t��<�q�;IE��r���;��>�=giŽ2)��(�;oh�>{�@>]�>�23="�=	��=���<�={��<�Oi�9@8����=��=�d >9�F>��>u��>��0?K?��>�!D�����7�Q��>~�=���>��N>�c�>t� ?�B"?�O@?̛[?�K�>m>S��>�D�>��@�7S��y־�gܭ<�x?�8�?��>�p���2��@�/S<�>��X'?��1?w�?%$`>�U����9Y&���.�"�����4��+=�mr��QU�S���Gm�5�㽯�=�p�>���>��>6Ty>�9>��N>�>��>�6�<|p�=6ጻ���<� �����=)�����<�vż����u&�7�+�'�����;z��;E�]<&��;v9�=p��>#%>���>o�=r䳾z0>������L���=�Ŧ��B� d�%J~�g�.�>�6�rmB>@�X>H����#��c�?SZ>�s@>���?��t?�o>����վ���R�d��Q�M.�=dq>)d=��B;�J`���M���Ѿ���>o؎>r΢>��n>ѩ*��_>��]�=2E�5�,��>]8��f���^�qq�~�������Sh���>:�TD?p�����=H�}?9UJ?.'�?��>�뚽~v׾;;,>��n=�L�1�k��L����?�'?���>z�쾡�B�ށ̾	�����>ӨH���O��͕���0���
��)���߰>^���_�о�:3��v���֏�?�B���r�o��>�IO?�ܮ?�b�BS��)O�!��sr����?��f?��>��?�O?ZQ��b�f���~T�=��n?D��?�/�?>0
>�`�=Oǂ���?�A�>��?+E�?GuX?�8�����>�L)>l�#>(D>�>�W>�2��J&x>�O?u�>��8?�rȽ�u	�.��L~�����z=m��=�R�>�V>�<X>�G�>���<+B�>��>�ك>�y>�_�>�{�>M�>�g[��QV��fC?���>��??#�5?W�	>���<���c+>�x��t�<�=T ��ٸ� ă>kL�=�
S��;�>�m=<���?Z�=�����J?6ޱ�w/�T�/:~|�>l�>�D�>���>.�">��'>���>vsx>;:�>��>�Ѿ��>^���S��3=��R�S�о��>M���v%1���Vb���O�����CX��oh�h避l�;�d��<9��?����g��'#�9��?X�>=�1?n�������=>���>��>,����㑿�j��>��u��?"��?<c>��>�W?�?Β1�(3��uZ��u�Z(A� e�5�`�x፿���ܗ
�����_?��x?'yA?MR�<:z>E��?��%�uӏ��)�>�/�';��@<=�+�>E*��L�`���Ӿ��þ�7�HF>��o?C%�?XY?HTV�Z���>�2?X�6?�]q?'0?hb=?.�=�u�.?%>�?�7?[�.?H�3?Ah?'yY>�>������=U.��T�~�촶�pD��:Ȱ�p�<�"�=��!<X�t<��=�ʧ<����@V���]�<A)'����;�&�<n)�=�̗=�ɱ>-U?��>�)\>��.?(����ҽ޾�@?�b�=�ǆ�.�"�.�Z��y̾V+�=��e?���?�^?ܢl>3c9��#�[��=O�M>�S�=�^R>,��>���X�@��y=��=�->Ĳ�=���9���y��pd�C�=��!>Y��>��y>o�X��EA>��7�k�k�_>-�K�o⯾��\�p�H�r%*��Ex�Ǽ>�A?y%?�n�=�z������d�?r�F??�S??�?� *=�׾n48�(K��������>�O=Ņ��G����v��m8+����kGI>m���䃾>"�>�,$���� |G��c� �d��^ܾ��"���=V��h|��t�l�	?�)���
m��㺿���S�P?4��WɾsdX���+�>��>�d�>$�'�IP�=$�����A{=��>�e>r'=�Y�v�,�H����q>?�V?�?7Yp?t؛�F�u��l�K�Ҿ�d����p����>�(?��"?�x>./�>�1ɾ����@���(��,�>R�(?�0��bO������+���s�>��?9Q>��?�VJ?pn?
?�?��5?�;?���>L�D����6�!?�3�?蘢=�����X���>�cxC�ϝ?�c)?�g#��q�>}�?p�?�H'?�KV?�@?�s>Ȅ���;�>��>n �>�Y����-�a>P�B?$��>ryM?��{?$W3>l�.�ޜ�4;��eN�=�>��.?�#?L5?1�>�ȶ>(h��PU�j�>�??�m?s`?!��=<@�>�0�<�D?�!�7y?��:>���>>U-?�~?&z]?��>,7���\άL󽣼���V��cmؼ��ƽ�A=�ɣ=����{���ؾݽm�>�����>�=��<K�Ľ�5�='T�=���>P��>�짾c�=�޾�z����>��̽�
i�_�c��ͼ�畼�/j>�n�>%�>F1N�N�=�M�>]>9�2��"1?��?J?���<��q��+�Mܼ=?�>��(?⺫<�E�- ��}D-�~Y<z�@?��C?�t��!���\�b?^?&Q�%=���þ��b�:z�M�O?h�
?�H�]ͳ>��~?C�q?���>/�e�0n���V@b�J�j���=D_�>~H�y�d��=�>��7?5�>@c>���=�s۾��w�3n���?N�?���?s�? �)>j�n�-�0���L��&J^?\��>�y���#?$��ۤϾX���eՎ�3v�̪�v����y���楾��%�!q����ֽ黼=�?�!s?qq?J?_?z� �l�c���]�(��V�������E���D��0C�xln�9;��
��显gD=o�v��j����?��:?w��<�?7���uǾk�����_>%�E����^�y�|��vh>R�佂U���q<\�Ś?v$	?y��>87?z�f�ľ$��
�U�������2>Re>�&R>�d?ֆa=�=�	�=�bW��t%d���;�a)k>��T?�[?q�w?�|�sd(�ς�QC#���<5�̾�h]>�ZL>�
>Mw[������%��'?�4w�~o���m��s��=@�=)�?��>�@�>+��?B�?���2��
D��HC����=n��>[Zz?� ?�9�>'�e���4�� �>J�l?���>��>䌾tO!���z�c�ǽ
�>4��>̑�>a�q>��/�H�[�DЎ�����8����=�!h?{���/y^����>�P?��;��4<f�>�U���!�Rg�0U,�W>l?\��=i�?>}�ž�5���|��W��wq)?�F
?�/��SZ&�鹍>�) ?�=�>���>Y�~?\��>*z���~;��?e�V?�XB?�;?g��>�vj=<���Ž��'��� =t��>`�Q>�>j=14o=n��dI���4�Tw=a��=E���H�˽u�< m�^L�;�=�4>�ڿ(U�W�ɾ���d�~������n ��ڕ��i쁽TӘ�P���b�������D�z�[)ɾ�����ᄾ���? �?D&��z�ž��y�W�N�6��=��G�֭_�#hb����=l�ξU�Ѽt��b�/�R�G�w�ɉ�ËC?B�E�qЖ�Ј�e���Z�?Y��?fYB?���,�)��7�� 	>�cJ�C=w( �G��Ϳ/T��
͆?�q�>�Ͼ�"�;�?�` >;�>^<�>tǾW�%���>~ܽ>��(?�E�>��tPҿ���Jψ����?��@�8?�n��k����_�`�>�U�>iW=>lxI���*�2RR�=��>MF�?�$u?��o<�<L����}vX?W�,�k�?��gT<��^=�S=@��=0�սa^w>1�s>'�t����Ŷ6��Q�>Yd>)@��Խ�I�w�:�o�h>�{.�PQ[�5Մ?+{\��f���/��T��U>��T?�*�>Z:�=��,?X7H�a}Ͽ�\��*a?�0�?���?$�(?7ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=`6��z���&V����=W��>c�>��,������O��I��V��=����տ[�!�
��q��| ��T�{�])H�Ⲿ�ܾ��/����\���f��!w�=1��>@�O>�V�>Rb>w�F?,�R?��>�~@=�J0>�Y�s���-�W��n��W<5�:]��xr�T,��Bʾ	c�8�"����f���.���*><`�-Ɖ�d����_�J�8���]?aR>�9j���K�`5/=M��{[��<,M��ƾ�4��H� ?<]^?�v��ꗿTz���y�?=b2?Gn���F�"Ѿ�>���Kwy>J.�>~=�=Jڽ�O'��8?�P�G?��??� ��V�[R?v2����>�?��=X��l6�>h]�>�U ��{f>��=L�/>
�w>Ă1?6;?U��=�׽V?�S?蕀�b����r=aҾM�[Y>��/<����[U�<H�>�н��˽ܬr����<k��=�%Y?�Е>�&,�m��z{H���S�=�w? T�>l�>��e?D?U�!���澁�M�����=�kS?��`?�3>�V���Qξ�۞�E8>?Ab?Z�>����,���.m0�G�����?k7\?�?ˉI���y�A���N����-?��v?�r^�rs�������V�e=�>\�>���>��9��k�>�>?�#��G��󺿿mY4�!Þ?��@|��?��;<q �<��=�;?k\�>��O��>ƾu{�������q=�"�>匧�lev����R,�]�8?Ԡ�?��>�������7գ=㾐�Cd�?�y�?A恾�D�=�~$�7QN�k��^{�Q �;�\ >)Gռ*�Ѿ����_�5��*�s�g�a<�B�>�N@!q��=��>F����I�ʿ{�r�tbǾS7Z��7�>֚?��>�e�#�)���L��z\����b̴��	�>YG�>��>z�;���w�o���>� ?���>���>���Dφ���:�Q|>�A�>��?Wc>�<z*���+�?Mw����i���^���>��?�e?�7?>!�>?���U੾Y��>�M6?8�?��k?�#����������o?
g������e۾�F"�Ht?Vm�?�#�=!���!�2>��і,?�7�������ؿ�ܿm����?L��?!����^�>f,�?��Y?V�%�)bb����[N+� ��>I�>�0=> ?�����wE���>��d�>F�>d�[>J�]�_?'�a�K�p���-���ƽ�ۡ>��0��e\��M�����Xe����@y����?M^�?i�?ֵ�� #�e6%?#�>a����8ǾW�<���>�(�>*N>3H_���u>����:��h	>���?�~�?Rj?���������U>	�}?n �>H�?���=0�>��=���VF���">6�=�\I��?LM?�e�>���=lA7�1~.�0�E�S�Q���:jC��_�>�"b?cZK?�)b>.���?�f��zѽ��4�$	��>��Y6���ݽ)?7>U/;>Ƚ>��J�F�Ҿ��?Mp�9�ؿ j�� p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>D�Խ����\�����7>1�B?Y��D��u�o�y�>���?
�@�ծ?ji��	?���P��Za~����7����=��7?�0��z>���>�=�nv�׻��G�s����>�B�?�{�?��>�l?��o�P�B���1=OM�>ڜk?�s?^o��󾁲B>��?�������K��f?�
@yu@]�^?"����⮿���E󾢐��R���C>�*(�����K��J��	����>^Cy>??>/|">���=�^>D�3>�o��z�)��}����k�p��.4�}��f?¾\8&�*�V�!�5��7��6����%���0���<*��%4���L��x�Z�=�W?BR?��o?���>�����'>����m,=� �M�=ӡ�>�;3?�L?�S-?>��=�ؙ�O�b�0��襾kV����>*�I>�a�> ��>F2�>���&*H>��@>�Dy>�l�=�r3=�Dp�U��<�+M>-�>��>�G�>�,Z>w��>:����ĵ���:��@��~9��@�?����:�)1��*P��q�߾�Lm>�r!?�A�<������ÿ�N��H�N?q��b]�f �P��>-�3?��<?�̽�л���K>p�=���Kxs���u=N����>��'��r�>X�?�V>E�A>��?�*E��uW���;.c�=%�?�q�����Q�A���+�{��S7>�w@>5�̽�E޾;M��������w���>D�?dp�>����峾AmO�Sב> �;�;�=�`���`�=�)=��)<��F�ߺ��>��>�G�>��>�s���}>���X�=�?�> !%�Ği>���>�5>?�fھ�Ğ>�M)�Җ\��t�>���>�P�>|��=0m��.�>�#?(;�>�B��4�C�j�<p�#��>/��G�!>F�&��R��܋�=1�O>����\.���=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>���˘�v�����t�]	0=���>/G?�k���;��@A���
?:?���錄ɿz�w���>Nt�?/p�?�Nm�ڢ��ff?�B��>�s�?f�X?$f>Zھ8p[��8�>��@?�Q?��>F����*���?=˶?���?HI>=��?��s?Aj�>�?x�DZ/�F5�������=�\;<c�>�X>^����eF�B֓�g��6�j�����a>1�$=D�>/佣7��);�=<����M���uf���>�(q>�I>�Z�>�� ?I^�>ʫ�>Qh=�y��k怾����"�K?`��?����8n�4�<�+�=�^��"?�04?r�Z���Ͼ�٨>�\?7��?��Z?ey�>k���6��T޿��]����<*zK>�3�>nU�>y��@cK>8�Ծ�>D��h�>�>�£�Sھ���F���1D�>Fh!?��>U�=�� ?ۘ#?S�j>�!�>\E�22����E�4��>��>CJ?e�~?A
?�ﹾ�V3�z���f١��[��
N>v�x?�V?Wȕ>����6���-�B��-K�e��£�?�_g?��Z�?;,�?io??ݞA?h�f>��1ؾ�]��]��>G^?�z*��>��b)�V���`
?�+�>]Ի>�x�Y�3� �����W���-�>}C?4�?�|羾�_��Sھ�s�<�59�c�;3J=�8�e>=>�ƛ��M�=�D>��=�z�2I1�膏;<=���>�7�=���Y�<�",?�g+�X����=�pr�;ZD�Ļ�>$:K>	���~^? =�KL{��ܬ��"���T��?'I�?�-�?�ᵽ��h�U�=?�!�?N�?+��>�����޾�W޾�Gw��z����J`>��>���~�㾬l��E���zp��|�ǽt	���>���>/+?��>�Uc>gJ�>�����*$�a��Qz����^�w�#�9�.-,����
��q "��b�ltž�W����>�`���\�>4��>L(>{
o>���>}��چ>.�Z>�Be>�\�>a�@>ۣL>ǣ�=��<�tý�R?B��R�'�UL��۰�ǴA?�^d? :�>͙g��[���'�?L<�?:�?Fu>�g�(�*�F:?��>�q���
?��>=�H�V��<� ��D{�VZ��#����>�XٽP�9�.MM�@d���	?
�?-ʏ��̾
ֽ����p�n=>K�?��(?��)��Q�p�o�)�W�S�b��N3h�wq���$�{�p��쏿�]��%��8�(��H*=��*?Q�?����������#k��?��Tf>��>"�>��>�I>��	���1�^��J'�ƾ��2J�>5R{?�y�=CP?C\?��?�?�i�>���<]��P(�>�H�a?J�.?�J?Q��>PBa?�^K?�R;?ն�>�m�������ؾ�H?��?�4O?/�E?�K?�����<)+�Ry�H�d�3�=BT�=z}���C��3$��"
=�a>��?�Fy�w�.�t;Ծ�{E>lbP?�/>HА>�Bʾ�F�=Rr(>�F=2?�a�=�m���e���:��>�1?���k�<�4>Mw�=�;������q�=,�����=��<<���;E?�{'>��K=��鼌�U�6�<<���=m�G��t�>��?���>�A�>�=���� ����i�=XY>�S>>KDپh}���#����g�%^y>jw�?&z�?��f=��=��=�{��cS�����5�����<��?I#?aWT?蕒?��=?Hj#?Ͷ>+��L��D^������?]V/?�F�>X����ž�����`'�Q�?:��>W*Z���ͽ��.�Ey������=F8�!�����t'@��u�=���R���H�?�?�I�W�+�)Q�8����m��%�9?��>�׫>R��>�_4�$�f�����$>1��>��U?��^>��?��?|�8?R��=cX�����8о�3�>�Π=�|S?��U?��|?`@�?�
�?�?�����M���������ګ��(ƾ�K=
@�=L�>���>Y&�>�)>_Q >��r=N�������&K=\��>��>z/�>��P>�b&��:??�?��Ⱦ��@��
<'S���>쏒?�4?i?/Ӡ��_��y(��Ƅ����>�E�?]��?Ζ�>��c>7oI�(ZA��f?��
u?V$?Ͷ>����8�=Dڽx 7?��>����Zs�\���s�=�PbM?�� ?0�'<l¿��s�y�l��'���)�;�]����t�e���̇k�ؗ�=�̙�����饾�e��؝�Z���&������u���H�>�Ce=^>E�=�Ć<BG����<��r=@N�;
Z=3ts��<�2��^g�V���{�$� ��<#�T=U���+˾�\}?
I?��+?h�C?(,z>�>i3���>�&��pU?�LU>��L����x;�����ɖ��Vؾ�׾$�c�۫����>�[H�!>l�2>62�=5��<1i�=�q=6�=c;T��=��=6]�=Q��=�1�=�>}�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�U�>h}���t���P�(����<m���|a=9uo�2$>�C�=F=
G�=�?վ
u�̑4��j�=m�O�|�GC>!@H�C�=�
>��*>l��>���<>ʼN��ǖ= W>!x�=p�6>�ơ�-Q=�B���&>��>u7V>���>��?"5?�"k?5��>w�6����%!��<��>��=���>)�L=X�/>ԃ�>��-?xv:?f�K?���>�D~=%�>B+�>WG'�N�v���p����W�<��?�V�?��>�r���N8�� ��00��}���I?x�)?F�?�>�v �����P3)�7�B��[�S2G��=Ʋ�^?��R慨h�ɾn�&��'>p3�>gZ�>a{�>oa�>�J+>9�>��>21>6M�=��|>�ݎ���=���8��<D��<�t�=K��=���<��<���2>*t��>1+�=D�`=�����D�=�n�>%w>�u�>�I�=(9��9@>P*��o�A���=CX��GF;�9'b�,qw��y)��a0�ۡ>>��T>A]��fn��� ?8�w>FZ2>��?WRj?8��=�o��:Uؾ����V��� g7����=;�=���x;��@a��MT��yҾ��>���=x 9?�=?A�A�(۾�,	�ӛK��H>�;�=�=���>��B�u졿����ܵ�DF���Ya>{�?�����=oю?G?�p?׋&=\ܾۖ���ν���R��>\ǜ��Ͼ���>�;?X�*?�::?��B�����F̾VS����>qI���O�t�����0�g��cϷ�a��>y��@�о� 3�}b��7����B��Kr���>X�O?j�?.�a��I��^}O����Z���m?xg?]
�>EJ?Y?���R��P2��'��=\�n?̠�?�*�?��
>�Cf�=�����>��a?��?[�?`O?��>nu9?�侾�Ӛ>tqI�>�U>�rؽ��=#�j>�@D?��A?d�$?[�\���־�9��L�F�v�����=X�p>�_�>Z�>�O���L�Ƌ ���=�o�=��!<��=�"�>pԀ>����l�&�|�m?��>q��>\g&?;?�=��>8���2il��.ս72�;���_;���AS�4/�ѭ0��Q>l�F>Vz�����?�'�=��/�F?� �ϰ>ٍC���>�,��E�>x:�=f�=��>*<�=n�T>+$�>��=3���Jr>G����$���7�iK������a}>&��"�����������|��裾9Z�� �h�{낿��H��h�<�?-	 �&Ke���$�ݽX�?|��>U:)?���#Yi��=1>���>1�>Y����=��������ֈ?���?�5c>�>�W?��?��1��3��pZ�.�u��"A�	e��`����q���Օ
������_?>�x?QzA?F�<�Cz>���?��%�ޏ�	�>!/��$;��O<=�-�>���;�`���Ӿ�þ�-��NF>��o?�"�?�V?`V���v<�>��?C�%?n�`?��4?8�?��j4?�M>}:?^}�>�@A?�1?c�?�$�=cW>�=x,�="�����|�T��J�N��޽��;�i"=��=�����Z<7�=К^�B�s=7f��z��=�<;9�<�,�=[�#>1Q�>��W?���>:��>��'?��޽�=2��p��w4?*L�=r��k���Z����Tl�>Co{?��?aF`?�0u>^�2�����g)>n`�>�Z>���>�Z�>1�ѽy��CO�;	V�=ixQ>�2=Y�۽��X����p8��,�R;o>0�>��>=&���#�=�y��3���A�n>+??�����UF�16��W0�#`�ɳ�>jW+?�W?;�`=�&Ͼ�̊�e4l�z?�3C?KSR?�s?0\�<�c����G��~y�>���=����x��Pː�m�=����=�`6>�I_��ߏ��ם>��7	���q�ãY�Yo¾x5>̀$�ЄƽOD�1̾�о�Ty>��=��@ؾ"� �ݝ����;J?�����qƾ��>��E��.|D>�"�>D"�>s���6�M���i��<�J�>d��>Q:�='.۾��)�A���g>�*H?�t?�n?�a�����:���������ǽ~?��>�?�e�<):\=W㍾���`.)��!����>=��>8���AT�t2��;R
�A=�>V?�iX>�tv>*kR?�>�z?C/ ?:5�>�'�>:��=ZI�G?�)�?s��=0�(�!lb�r$e����~:"?Y*?����~�>1x>�#?�DC?N8?Qk�>��)>߾�&T�۩�>�;>�vz�m?����!>��?��>á?�2K?��V>#��Pbh�]^t��Z>aZ>�?7�>���>��:>�1G>���D^�=�,?_�b?�Ǒ?ܙR?xN�>|�?ސ׾g$O?�eK>W�!?��>�^?��j?�Ċ?b�?�9�>e�;ؠ���ͼ��b� ��>��ʵ��=M���]�w���,>���>A4A�&=½Zk��h���hP�!`��� �>�Zs>2��5H>}��C���3+N>�O�<���`�.W'���=�>x>�h?��>eB,���=���>H3�>/���?���>O|?>0'=	"b�"=��To��]�>�!=??�>�=k��q���ar���=kFb?��V?�Df�
���dY?Ή_?�U��1K��aȾBO{����_RZ?���>�)y�8q�>{�o?��T?�P?3��7Bv�xי��m_�҃C� A�=�z>��s`���>g1?�e�>41m>_��=�U�y
_�o��L��>s��?=�?އ�?�T>q�AT޿Bm���ّ��^?/s�>�У�D�"?Z%���ξ�3��G������}ȩ�ᷫ�@Y��K����"&��]����ҽ4��=�"?Z�q?rsp?t'_?����c���]�Bi~��rV�[:����|E� E���C�Ho�R��˰�
S����H=�Lu��<<�œ�?��5?	lb����>����վ�ϕ���;"ƾ#��m�>��L��ī=ο�p������K�x�]s?5^�>A�>q�?q�e�1B�}��A����߾#؃>�>���>T�>��޻[	��8�-��W��W��N�r>�b?�SM?�p?@���>�0��i���K#��*��E��yW=>�k>@<�>��h��"���%�>��o��'��A�������=��0?�>X�>�S�?��?�>������u���0�%�<U�>�i?���>s��>��޽q�!����>��f?O�>�U�>�J���� ��~}�'<��Y�>*L�>�#�>�49>{�.�95{�؉��ￍ��RB���>t?�V���]��ꋦ>L�P?�>���q"����>_�*��N쾯�	�Y��=5 	?��>�!c>V�� <ӾXŃ�7?���-?�z?��m�pq�m�->�%?~�>Hk�>��Q?̽�>`ۿ��F>C@?�]?�/3?�I?�>��:=2�G�%׀�\�:��&�;��{>I�>9Y>C��=w3D���W^��M�=�=y���)�)�nx�k�_�C&r=��+=3�f>�"ۿ��o�ܬ�ތ��������y��	���AϾ�݆��I�N���{;��_�IJֽ4��l��吻��L��\��?��?�b��$�	��C����<������G�>>��fp<82����=�о�=��P>�%�#��q_��rb��:y��[-?��5ǿi���5\�y�v?l(�>��?���A2�1����>]]o�������4Ν��\ؿ�����e�?l�>���"���>���==�^>2��>�ŽlX���s�et>��+?vHT>)�Y�O���m�ʿ��-�$��?���?EC?N�#�U��S=�=?s?Z�+>�)��R���v��>�;�?�ā?W�H=6�[�������`?tpٻ��;��{t��{�=gW�=��=�����<>n�>��i�#�}��y�>曁>��μ���p�c�Hg�<��K>����ڽՄ?�z\�Nf�m�/��T���T>��T?�*�>�8�=�,?�6H�2}ϿT�\��*a?�0�?���?��(?Gۿ�ך>��ܾ�M?�D6?���>�d&���t���=!%ἂL�����v&V�U��=ެ�>'�>.�,�����O��W�����=���v�޿"8&�M 	��@�⃾~��zʳ�oĝ����V`ľ���9�B�v����=M�>:�.>�M>2�'>�LV?UQ@?N�>i�>�TϽ�l�.�������K;�6#�=��ľ�Ͻo ھ_ǥ��ɝ��Զ���(��C�!�达�8���=�O�$�����M��fW��S=����>����������{��@U>��s|�6_?�=����Y��XI��f~�p:�?o$k?tm�:�N��<�y����m��jo?��Q�<�E{c�$h�<�4E���S>0~�>�l<�L��]�C�F<W���E?���>�T־�����?���
���_'?4g�>(�r>9>ML�>a�R�GT�=�0����=P��>�ۅ>2.�=6=Ծ�A=,�2?�H?x���ʽ�|=b鴾�>=�=��k�Je~���>�^T>h*�>�v���I��+~T>��4�)�Y?@o�>[��_k�fC�;(<��^>w�X?U1?A�>`P?\�K?T�X<����-�A���־��q�B�O?�Oy?���=�����@��|n��]�?˚W?�}\>�S�|.���V*�]��?��c?�B�>��۽� ��1���䕾);??��v?s^�xs�����J�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?�;<��U��=�;?l\�>��O��>ƾ�z������5�q=�"�>���ev����R,�f�8?ݠ�?���>������(G�=�3��1)�?�߁?�Y������&����i�����yҝ��B@=$��3�S<%��H����gU��qS���8l<�C�>h@�R�DT�>�r���ڿ|vп�\���ľ�Ω���1?�b?��>�s|���_�gPG�Q�&���:�Wu��My�>@P}>O!ٽԚ��$�H��}��&>m?p� �U�n>/Û�O[���p��d#>4�=>��>��9>_-N���O֫?R\־{���L��	$�r�f??A?�?�?Ÿ��Ꮎg!>P)?
rT?��S?�Г���b19>Y�J?V���fS�K{?��f7�/��>�6k?^(�>z�������]�6��>}(�O�b�lǿ�ƿ�|��~�?�u�?s��.($?���?���>Z� ������hξC��x�>@��!��6]���$6���!�=��9�>�E̽���X�_?4�a�{�p���-�h�ƽ)ܡ>\�0��f\�(P����$Xe����Ay�f��?^�?E�?���=#�?6%?;�>Ş���8Ǿ�<\��>)�>�)N>�K_��u>���:��h	>|��?-~�?;j?͕������?U>��}?��>~�?���=N�>�P�=c᰾�t8��J#>���=Ij<�J�?{hM?�P�>���=Td8���.���E���Q�B(�h�C�F�>��a?�L?w�b>����3��!�E�ʽ��1��a��e@�/=*�1m�0#5>�=>�x>x�C��pҾO�?j���ؿ�j��nu'�=04?���>� ?B��h�t�>��9_?vr�>74��,��'��N����?xE�?��?ػ׾�\̼��>"�>9J�>x�Խ�ꟽ|���7>P�B?Z�KE����o��>\��?��@�Ѯ?Bi�_	?��#P���_~����i�6����=��7?�0�U�z>���>��=�nv�ǻ��l�s� ��>�B�?P{�?���>߮l?ހo�>�B���1=�K�>#�k?st?�1o�L󾘳B>�?�������aL�^f?��
@cu@˝^?����鿅⫿a}Ѿ]�׾0��l�<��=5\A��7+>��w��:y��'F��=��>]:T>G#7>p�d>oi�>�>n����"�4-���╿>=o�>��~���s¾�%��'O�,��&��s���� н�LD��m��L]	���l�����~Ӷ=)Y?�[N?!�k?�)�>��+��>D����@(��n\��%�=g�>ZD%?2t7?�g?�b�=(��4�c�L���wI������/�>�hf>���>��>Y�>�rB�܃�=�B>T�>Ao>l�>�~��}Թ`E>f�>�g�>�l�>��A>] �=t����㦿�{��F��`��!��?�Ҿ� &�r�Ӛ��!�~?>�G?Y��=�Ď���Ͽ�����a?X�����0��ڽ�c�>m�Z?l�O?��_�*�er>�cz>�]��鳽�$Ӽ�:��s���f�"�>?2=�L?��0>�>-��T'��Q�ҙ�تh>e�"?�aþ	�]�6`�Xq>�3�<�7?*�~>���=���T����ؑ��R���ѵ>�\?WM5?�n��7�j���\�J>��ps�>�Jؾ~��>�>����=�T���� =뽗J>�?�#>�<ټ��q>͈����v�p��>�{=D���@?�J"?�c�̍��v����p��4چ>���>�=>�=�E)���]F>տ?T��>�r�������c�1;⽦w�>�m�k���mý���=d��=�J����#���+��)=�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�-)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>э�~)��A����o��o6�U��>s�Q?���_T��:"q�@�?U��>U��X��;�˿��x�=��>���?ƽ�?�6b��l���M>�C(�>���?�a?嵉>�2������M�>i=?;';?d1�>Q���i����%?}ݫ?pqh?�>>=2�?��c?.�>�9��m�0������1�����e-=c�v>�K�=w�Ⱦ<P�j������ p��H����>�"=㋽>�����௾��=�˂�`�� *��׮>4p�>��1>Q�>ʘ�>��>4�>�ک=�X ���a�囤��K?�n�?I����m�8�<`]�=HA\�dM?*B3?c�;��ξŪ�>?\?��?)lZ?X/�>�������hӿ�����>q<חK>A�>�v�>^H~��2L>��Ծ�D���>�ޖ>N�}��5ھҹ��>�ۻiԞ>�
!?CI�>ɻ�=��?B_%?b>x��>�D�⑿�?�'�>-��>%G?_w?��?sd��	2����r䢿�>\���D>�^x?B�?B�>����E���FB��>��Q�Ƃ?�Ch?�d��?>�?�:?}�H?_3]>����Ǿ�٫�(�j>u"?| D��[L���G��E>�A&?N(?���>��a�y>�>�<�=p���H�۫*?��?�v>?G��^�x��Ϲ��؍=g@�d\��5�_>(��=ě�>��=CY�����>|	�>�:O=�q�<>�ϽF���N&>پ�>]��q��=���=!@,?n	H��䃾*ژ=߽r�.vD���>�NL>��F�^?~S=���{����4u��EU����?���?~e�?z㴽�h��=?�?J?�+�>{N��
�޾��z9w��x�$t���>���>�mm��徯���)����D��F�Ž˂��{�>�n/?��?T�? x�=�;#<��ľe�о�R�u��1TJ��?��,�^�����b=�X��:�ǽ
�T>�ґ�NIþ�	�>`� �w&�>�p�>�>#�>� �>�쇾�<�<��>̳�>��>��>���=�?������/S?vB��X(��.������@?׬e?�4�>�_v��������?�ȑ?E��?Iq>ig���'�"�?8q�>�|���?(=���.�=K0��a���Q��z�2�&��>@8���L:�0P���d���?�r?��X�;Ͼȡƽ<���\ o=8O�?��(?��)���Q��o��W�rS�����*h��Z����$�4�p�P珿�Z��'��S�(��*=�*?Z�?+��'���#��*&k��?� of>���>@&�>�׾> �I>��	�ͱ1��^�w>'����&?�>�H{?©J>_�I?�xQ?F�{?�p5?��>ԫ'�qR׾?I?o�=ǜ?!�>��l?Ez�>�oG?VZ�>h`?��? �	��o�Xf���L?vE?�I?v��>n�f>�F���1>)������>h�6�	�O������A��N)N=�X>��>�J?��A�9�<B�� �>0�.?L��>8G�>�񐾈�E���,=ȑ�>���>�Q�>6)	��n��9����>�R�?e��
y9=&�;>�S�=�P��~����=դ��(M�=ea,�z=����<�(�=��=K���?��<�����8=���Um�>E�?'��>�N�>�%��t� ���{�=/�X>S>�>2پez��;$����g�NLy>�v�?�w�?��f=�C�=��=g���(f���������b9�<!�?�H#?�YT?���?��=?h#?�>\%��E��_\������?a7(?��>��
���̾E����h4�m$?�C?�x]�V�!�(�*��Oɾ:�-��=�~5�	���$F��܏>�N��<�d���W��A�?�ƚ?TM�K8������#��X����+@?���>�ݔ>�c�>�/��2d����$@>n��>'oM?,p�>�I?7��?+D? �-I)�垠�_𔿒�>+��>ڦ�>%��?�?��K?M?�D>ք�/�5�pﾂPU=hc��+���-��-�5>��>�,�>�>J����B�=�E�i2"���}>��>'��>+�>̷�>>tS>����3X?�m�>��վ���P�o��>���> �?��?�}D?x:�}��Ș
������>|]�?�ݤ?۵?�]�([>�'Ƚ�侩_]�?�?�Z�>��s>Ņ�=�^��w�c>!?��>�N�r�	��*�8�	�!Z?Ia?��>X�ſ�t�i@`�֑��d<~t����n��m���rU��]q=���\�$�����T0a��C������
���E�����r�wQ�>LA�=g7�=���=�n�<w�&=��`=� �<�L1=F���r��<�\h�!m��n�c��6ͻ�7<��< �r��<˾X�}?)I?�,?.�A?�h>>8�H��w�>JU���V?�$F>L�>轾\�;��y��ܱ����ھ<wپ3/d�
ܟ�N�>��8���>�-0>T^�=��z<T�=d�w=0�=U7�9�{M=���=3m�=?��=���=1J>r1>�6w?M�������4Q�o[罭�:?�8�>1z�=��ƾ�@?��>>�2������Fb��-?a��?�T�?��?�ti��d�>����㎽2r�=����?2>���=��2����>�J>f���J������84�?��@��??�ዿ��Ͽ�b/>�WU>=r�>"�7�)�!�S̔�dy�����?G7�H헾4�>����Ul��VŁ�]�<�p>\S]=��{���h�o�#>aN�<�����<�n�>+��>��4>T���<[�0>��A<���>�=��@�Y�>�>�T�>�,>	��>�W?c�.?+"j?���>��-���Ҿ����>L�=�W�>�'=4[>k��>��,?�1?sN?)��>��{=�>O��>�Z���i�6�P����>{iv?���?���>΂�=q��i��x'5��}D��)'?�f%?��?WQ�>v��������B���4�H�����ǽG��5�����+%���4���n���'�=��5>��>Ge�>�b�>0�}>�>�?�>w�8=]��;ܱ�=�O
>0򾼯���47�=(a��ʢ��M�(>�H�>T��օ��X���=��U�/ņ=H��<ʼ�=���>��>98�>bj�=���L�#>F����J�}��=�s����?�;�b���{��.���:��'F>�aU>�Mw��O�����>Y>zhF>Ds�?��r?��>���Ҿ�Jp���V��*�=�&>ˏG���:��__��^L�cϾ��>��>Xi�>�Y>���6+���>� H���)���>�iԾ�{9�8Z��ߡ�0�������刿z[Z=�a{?�Eo���=B?yP?��f?�>�O��~�׾ߟ"�k���
>�}��Á�NR��.�?�;?)�%?9�(�hE;�9�Ⱦ�,��m��>z�Q���K�O(���.����;�LþԮ>
`���;Y2�����,�����G��'��f�>Y$P?�G�?Z��C{�z�L��������?��h?ѥ>�7�>2*?��f�K�R�b�?��=�o?��?��?m��=�$<xቾ߁?|�E?I�?M�?qX)?y*�=}>4?3�N��:�>�b;�:�>K	��/�>�
�>v+?]M?�4?�񑽗v
�ex��pLվ�]�
z�O8�>6B|>\;�=�AW>�d�z��=쾜=��(>7��>9%b>v=m>ӕ
?�>閾,���1?�x4>N}�>��'?88/>l�;��,���.��ī�6�L��$��8ʽ7R��bw�����m�2=�g����>f�¿1��?��J>�����!?�Dľk��<&'D>]�,>�r�Q�>g��=�\>S��> �>��>��m>�
%>T8Ҿ�h>t��m!�SC�M�Q�,�о�Ny>r䜾j�#����Q���?J��0�����i��-���=��q�<��?7���Yk���)�����t�?���>"�5?�������"�>2��>�>%N��NP��B���o�C�?��?ӱb>���>|�W?f�?�9/���1�/�Z��Ou�D�@��e��`����1��ۂ
����%F_?c�x?�hA?~f�<��y>@p�?��%�)ޏ�C�>X�.�w�:��A=�U�>����Oa���Ӿ��þ�����D>�-o?C+�??�V�pB��K>�4?x�0?��k?�z7?e�3?����9$?��'>�q	?9�?:�8?�(?�~?�K^>r">��'=��<VȆ������ͽ8�뽨� �:N=�=��[:�ԼEٖ<���<��F�����R�*�'�B��i�<�S=��=�_�=��>��U?-�>�Q�>��>?�� >9��۟�6e4?E�=��f�x3������o�㾨l >v�^?���?vX?�;[>�L�V�F��Z>�ш>:� >Y�M>rg�>)߽ۡC�_Z=Y�=�<>j+�=�妽 ����9�EĒ�!`=�4>���>�>?<�Eq�=�W�(
���C�>3��<YnȾF���<\���F�UᖾJ�>�� ?X� ?o<�=�G�PM��Y����>-�7?�U?��y?�νqf��b�#)[��_'�
B�>�D��Vg������>����"��xԽ|��=�5Ͻ�䃾>"�>�,$���� |G��c� �d��^ܾ��"���=V��h|��t�l�	?�)���
m��㺿���S�P?4��WɾsdX���+�>��>�d�>$�'�IP�=$�����A{=��>�e>r'=�Y�v�,�H����q>?�V?�?7Yp?t؛�F�u��l�K�Ҿ�d����p����>�(?��"?�x>./�>�1ɾ����@���(��,�>R�(?�0��bO������+���s�>��?9Q>��?�VJ?pn?
?�?��5?�;?���>L�D����6�!?�3�?蘢=�����X���>�cxC�ϝ?�c)?�g#��q�>}�?p�?�H'?�KV?�@?�s>Ȅ���;�>��>n �>�Y����-�a>P�B?$��>ryM?��{?$W3>l�.�ޜ�4;��eN�=�>��.?�#?L5?1�>�ȶ>(h��PU�j�>�??�m?s`?!��=<@�>�0�<�D?�!�7y?��:>���>>U-?�~?&z]?��>,7���\άL󽣼���V��cmؼ��ƽ�A=�ɣ=����{���ؾݽm�>�����>�=��<K�Ľ�5�='T�=���>P��>�짾c�=�޾�z����>��̽�
i�_�c��ͼ�畼�/j>�n�>%�>F1N�N�=�M�>]>9�2��"1?��?J?���<��q��+�Mܼ=?�>��(?⺫<�E�- ��}D-�~Y<z�@?��C?�t��!���\�b?^?&Q�%=���þ��b�:z�M�O?h�
?�H�]ͳ>��~?C�q?���>/�e�0n���V@b�J�j���=D_�>~H�y�d��=�>��7?5�>@c>���=�s۾��w�3n���?N�?���?s�? �)>j�n�-�0���L��&J^?\��>�y���#?$��ۤϾX���eՎ�3v�̪�v����y���楾��%�!q����ֽ黼=�?�!s?qq?J?_?z� �l�c���]�(��V�������E���D��0C�xln�9;��
��显gD=o�v��j����?��:?w��<�?7���uǾk�����_>%�E����^�y�|��vh>R�佂U���q<\�Ś?v$	?y��>87?z�f�ľ$��
�U�������2>Re>�&R>�d?ֆa=�=�	�=�bW��t%d���;�a)k>��T?�[?q�w?�|�sd(�ς�QC#���<5�̾�h]>�ZL>�
>Mw[������%��'?�4w�~o���m��s��=@�=)�?��>�@�>+��?B�?���2��
D��HC����=n��>[Zz?� ?�9�>'�e���4�� �>J�l?���>��>䌾tO!���z�c�ǽ
�>4��>̑�>a�q>��/�H�[�DЎ�����8����=�!h?{���/y^����>�P?��;��4<f�>�U���!�Rg�0U,�W>l?\��=i�?>}�ž�5���|��W��wq)?�F
?�/��SZ&�鹍>�) ?�=�>���>Y�~?\��>*z���~;��?e�V?�XB?�;?g��>�vj=<���Ž��'��� =t��>`�Q>�>j=14o=n��dI���4�Tw=a��=E���H�˽u�< m�^L�;�=�4>�ڿ(U�W�ɾ���d�~������n ��ڕ��i쁽TӘ�P���b�������D�z�[)ɾ�����ᄾ���? �?D&��z�ž��y�W�N�6��=��G�֭_�#hb����=l�ξU�Ѽt��b�/�R�G�w�ɉ�ËC?B�E�qЖ�Ј�e���Z�?Y��?fYB?���,�)��7�� 	>�cJ�C=w( �G��Ϳ/T��
͆?�q�>�Ͼ�"�;�?�` >;�>^<�>tǾW�%���>~ܽ>��(?�E�>��tPҿ���Jψ����?��@�8?�n��k����_�`�>�U�>iW=>lxI���*�2RR�=��>MF�?�$u?��o<�<L����}vX?W�,�k�?��gT<��^=�S=@��=0�սa^w>1�s>'�t����Ŷ6��Q�>Yd>)@��Խ�I�w�:�o�h>�{.�PQ[�5Մ?+{\��f���/��T��U>��T?�*�>Z:�=��,?X7H�a}Ͽ�\��*a?�0�?���?$�(?7ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=`6��z���&V����=W��>c�>��,������O��I��V��=����տ[�!�
��q��| ��T�{�])H�Ⲿ�ܾ��/����\���f��!w�=1��>@�O>�V�>Rb>w�F?,�R?��>�~@=�J0>�Y�s���-�W��n��W<5�:]��xr�T,��Bʾ	c�8�"����f���.���*><`�-Ɖ�d����_�J�8���]?aR>�9j���K�`5/=M��{[��<,M��ƾ�4��H� ?<]^?�v��ꗿTz���y�?=b2?Gn���F�"Ѿ�>���Kwy>J.�>~=�=Jڽ�O'��8?�P�G?��??� ��V�[R?v2����>�?��=X��l6�>h]�>�U ��{f>��=L�/>
�w>Ă1?6;?U��=�׽V?�S?蕀�b����r=aҾM�[Y>��/<����[U�<H�>�н��˽ܬr����<k��=�%Y?�Е>�&,�m��z{H���S�=�w? T�>l�>��e?D?U�!���澁�M�����=�kS?��`?�3>�V���Qξ�۞�E8>?Ab?Z�>����,���.m0�G�����?k7\?�?ˉI���y�A���N����-?��v?�r^�rs�������V�e=�>\�>���>��9��k�>�>?�#��G��󺿿mY4�!Þ?��@|��?��;<q �<��=�;?k\�>��O��>ƾu{�������q=�"�>匧�lev����R,�]�8?Ԡ�?��>�������7գ=㾐�Cd�?�y�?A恾�D�=�~$�7QN�k��^{�Q �;�\ >)Gռ*�Ѿ����_�5��*�s�g�a<�B�>�N@!q��=��>F����I�ʿ{�r�tbǾS7Z��7�>֚?��>�e�#�)���L��z\����b̴��	�>YG�>��>z�;���w�o���>� ?���>���>���Dφ���:�Q|>�A�>��?Wc>�<z*���+�?Mw����i���^���>��?�e?�7?>!�>?���U੾Y��>�M6?8�?��k?�#����������o?
g������e۾�F"�Ht?Vm�?�#�=!���!�2>��і,?�7�������ؿ�ܿm����?L��?!����^�>f,�?��Y?V�%�)bb����[N+� ��>I�>�0=> ?�����wE���>��d�>F�>d�[>J�]�_?'�a�K�p���-���ƽ�ۡ>��0��e\��M�����Xe����@y����?M^�?i�?ֵ�� #�e6%?#�>a����8ǾW�<���>�(�>*N>3H_���u>����:��h	>���?�~�?Rj?���������U>	�}?n �>H�?���=0�>��=���VF���">6�=�\I��?LM?�e�>���=lA7�1~.�0�E�S�Q���:jC��_�>�"b?cZK?�)b>.���?�f��zѽ��4�$	��>��Y6���ݽ)?7>U/;>Ƚ>��J�F�Ҿ��?Mp�9�ؿ j�� p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>D�Խ����\�����7>1�B?Y��D��u�o�y�>���?
�@�ծ?ji��	?���P��Za~����7����=��7?�0��z>���>�=�nv�׻��G�s����>�B�?�{�?��>�l?��o�P�B���1=OM�>ڜk?�s?^o��󾁲B>��?�������K��f?�
@yu@]�^?"����⮿���E󾢐��R���C>�*(�����K��J��	����>^Cy>??>/|">���=�^>D�3>�o��z�)��}����k�p��.4�}��f?¾\8&�*�V�!�5��7��6����%���0���<*��%4���L��x�Z�=�W?BR?��o?���>�����'>����m,=� �M�=ӡ�>�;3?�L?�S-?>��=�ؙ�O�b�0��襾kV����>*�I>�a�> ��>F2�>���&*H>��@>�Dy>�l�=�r3=�Dp�U��<�+M>-�>��>�G�>�,Z>w��>:����ĵ���:��@��~9��@�?����:�)1��*P��q�߾�Lm>�r!?�A�<������ÿ�N��H�N?q��b]�f �P��>-�3?��<?�̽�л���K>p�=���Kxs���u=N����>��'��r�>X�?�V>E�A>��?�*E��uW���;.c�=%�?�q�����Q�A���+�{��S7>�w@>5�̽�E޾;M��������w���>D�?dp�>����峾AmO�Sב> �;�;�=�`���`�=�)=��)<��F�ߺ��>��>�G�>��>�s���}>���X�=�?�> !%�Ği>���>�5>?�fھ�Ğ>�M)�Җ\��t�>���>�P�>|��=0m��.�>�#?(;�>�B��4�C�j�<p�#��>/��G�!>F�&��R��܋�=1�O>����\.���=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>���˘�v�����t�]	0=���>/G?�k���;��@A���
?:?���錄ɿz�w���>Nt�?/p�?�Nm�ڢ��ff?�B��>�s�?f�X?$f>Zھ8p[��8�>��@?�Q?��>F����*���?=˶?���?HI>=��?��s?Aj�>�?x�DZ/�F5�������=�\;<c�>�X>^����eF�B֓�g��6�j�����a>1�$=D�>/佣7��);�=<����M���uf���>�(q>�I>�Z�>�� ?I^�>ʫ�>Qh=�y��k怾����"�K?`��?����8n�4�<�+�=�^��"?�04?r�Z���Ͼ�٨>�\?7��?��Z?ey�>k���6��T޿��]����<*zK>�3�>nU�>y��@cK>8�Ծ�>D��h�>�>�£�Sھ���F���1D�>Fh!?��>U�=�� ?ۘ#?S�j>�!�>\E�22����E�4��>��>CJ?e�~?A
?�ﹾ�V3�z���f١��[��
N>v�x?�V?Wȕ>����6���-�B��-K�e��£�?�_g?��Z�?;,�?io??ݞA?h�f>��1ؾ�]��]��>G^?�z*��>��b)�V���`
?�+�>]Ի>�x�Y�3� �����W���-�>}C?4�?�|羾�_��Sھ�s�<�59�c�;3J=�8�e>=>�ƛ��M�=�D>��=�z�2I1�膏;<=���>�7�=���Y�<�",?�g+�X����=�pr�;ZD�Ļ�>$:K>	���~^? =�KL{��ܬ��"���T��?'I�?�-�?�ᵽ��h�U�=?�!�?N�?+��>�����޾�W޾�Gw��z����J`>��>���~�㾬l��E���zp��|�ǽt	���>���>/+?��>�Uc>gJ�>�����*$�a��Qz����^�w�#�9�.-,����
��q "��b�ltž�W����>�`���\�>4��>L(>{
o>���>}��چ>.�Z>�Be>�\�>a�@>ۣL>ǣ�=��<�tý�R?B��R�'�UL��۰�ǴA?�^d? :�>͙g��[���'�?L<�?:�?Fu>�g�(�*�F:?��>�q���
?��>=�H�V��<� ��D{�VZ��#����>�XٽP�9�.MM�@d���	?
�?-ʏ��̾
ֽ����p�n=>K�?��(?��)��Q�p�o�)�W�S�b��N3h�wq���$�{�p��쏿�]��%��8�(��H*=��*?Q�?����������#k��?��Tf>��>"�>��>�I>��	���1�^��J'�ƾ��2J�>5R{?�y�=CP?C\?��?�?�i�>���<]��P(�>�H�a?J�.?�J?Q��>PBa?�^K?�R;?ն�>�m�������ؾ�H?��?�4O?/�E?�K?�����<)+�Ry�H�d�3�=BT�=z}���C��3$��"
=�a>��?�Fy�w�.�t;Ծ�{E>lbP?�/>HА>�Bʾ�F�=Rr(>�F=2?�a�=�m���e���:��>�1?���k�<�4>Mw�=�;������q�=,�����=��<<���;E?�{'>��K=��鼌�U�6�<<���=m�G��t�>��?���>�A�>�=���� ����i�=XY>�S>>KDپh}���#����g�%^y>jw�?&z�?��f=��=��=�{��cS�����5�����<��?I#?aWT?蕒?��=?Hj#?Ͷ>+��L��D^������?]V/?�F�>X����ž�����`'�Q�?:��>W*Z���ͽ��.�Ey������=F8�!�����t'@��u�=���R���H�?�?�I�W�+�)Q�8����m��%�9?��>�׫>R��>�_4�$�f�����$>1��>��U?��^>��?��?|�8?R��=cX�����8о�3�>�Π=�|S?��U?��|?`@�?�
�?�?�����M���������ګ��(ƾ�K=
@�=L�>���>Y&�>�)>_Q >��r=N�������&K=\��>��>z/�>��P>�b&��:??�?��Ⱦ��@��
<'S���>쏒?�4?i?/Ӡ��_��y(��Ƅ����>�E�?]��?Ζ�>��c>7oI�(ZA��f?��
u?V$?Ͷ>����8�=Dڽx 7?��>����Zs�\���s�=�PbM?�� ?0�'<l¿��s�y�l��'���)�;�]����t�e���̇k�ؗ�=�̙�����饾�e��؝�Z���&������u���H�>�Ce=^>E�=�Ć<BG����<��r=@N�;
Z=3ts��<�2��^g�V���{�$� ��<#�T=U���+˾�\}?
I?��+?h�C?(,z>�>i3���>�&��pU?�LU>��L����x;�����ɖ��Vؾ�׾$�c�۫����>�[H�!>l�2>62�=5��<1i�=�q=6�=c;T��=��=6]�=Q��=�1�=�>}�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�U�>h}���t���P�(����<m���|a=9uo�2$>�C�=F=
G�=�?վ
u�̑4��j�=m�O�|�GC>!@H�C�=�
>��*>l��>���<>ʼN��ǖ= W>!x�=p�6>�ơ�-Q=�B���&>��>u7V>���>��?"5?�"k?5��>w�6����%!��<��>��=���>)�L=X�/>ԃ�>��-?xv:?f�K?���>�D~=%�>B+�>WG'�N�v���p����W�<��?�V�?��>�r���N8�� ��00��}���I?x�)?F�?�>�v �����P3)�7�B��[�S2G��=Ʋ�^?��R慨h�ɾn�&��'>p3�>gZ�>a{�>oa�>�J+>9�>��>21>6M�=��|>�ݎ���=���8��<D��<�t�=K��=���<��<���2>*t��>1+�=D�`=�����D�=�n�>%w>�u�>�I�=(9��9@>P*��o�A���=CX��GF;�9'b�,qw��y)��a0�ۡ>>��T>A]��fn��� ?8�w>FZ2>��?WRj?8��=�o��:Uؾ����V��� g7����=;�=���x;��@a��MT��yҾ��>���=x 9?�=?A�A�(۾�,	�ӛK��H>�;�=�=���>��B�u졿����ܵ�DF���Ya>{�?�����=oю?G?�p?׋&=\ܾۖ���ν���R��>\ǜ��Ͼ���>�;?X�*?�::?��B�����F̾VS����>qI���O�t�����0�g��cϷ�a��>y��@�о� 3�}b��7����B��Kr���>X�O?j�?.�a��I��^}O����Z���m?xg?]
�>EJ?Y?���R��P2��'��=\�n?̠�?�*�?��
>�Cf�=�����>��a?��?[�?`O?��>nu9?�侾�Ӛ>tqI�>�U>�rؽ��=#�j>�@D?��A?d�$?[�\���־�9��L�F�v�����=X�p>�_�>Z�>�O���L�Ƌ ���=�o�=��!<��=�"�>pԀ>����l�&�|�m?��>q��>\g&?;?�=��>8���2il��.ս72�;���_;���AS�4/�ѭ0��Q>l�F>Vz�����?�'�=��/�F?� �ϰ>ٍC���>�,��E�>x:�=f�=��>*<�=n�T>+$�>��=3���Jr>G����$���7�iK������a}>&��"�����������|��裾9Z�� �h�{낿��H��h�<�?-	 �&Ke���$�ݽX�?|��>U:)?���#Yi��=1>���>1�>Y����=��������ֈ?���?�5c>�>�W?��?��1��3��pZ�.�u��"A�	e��`����q���Օ
������_?>�x?QzA?F�<�Cz>���?��%�ޏ�	�>!/��$;��O<=�-�>���;�`���Ӿ�þ�-��NF>��o?�"�?�V?`V���v<�>��?C�%?n�`?��4?8�?��j4?�M>}:?^}�>�@A?�1?c�?�$�=cW>�=x,�="�����|�T��J�N��޽��;�i"=��=�����Z<7�=К^�B�s=7f��z��=�<;9�<�,�=[�#>1Q�>��W?���>:��>��'?��޽�=2��p��w4?*L�=r��k���Z����Tl�>Co{?��?aF`?�0u>^�2�����g)>n`�>�Z>���>�Z�>1�ѽy��CO�;	V�=ixQ>�2=Y�۽��X����p8��,�R;o>0�>��>=&���#�=�y��3���A�n>+??�����UF�16��W0�#`�ɳ�>jW+?�W?;�`=�&Ͼ�̊�e4l�z?�3C?KSR?�s?0\�<�c����G��~y�>���=����x��Pː�m�=����=�`6>�I_��ۍ���w>�n�����f��;U�>�;�=��I��=��&������5���^6>�Da=�4¾��+�{<������G?*>�+��}H��}=���B�=v�>I��>L2�;��
��*K�(r���> ��>t�V>�{=��n`A�a����l>��:?��n?W�m?���ދ��8V������(�ƈ?��1!?&�?i�>�j�>��׻���������/�Y**� ��>��3?�+"�E�,�����̱!�m>��/�>h?�ţ>J�?�/?��?6�y?�a?�?L�>�����׾SK?i��?�D�=�o��7�q��#R��+2���?�a?�_�U<>	?�-�>\xo?ףT?�Q�>���=�7��RG�Ɗ�>%>�> �S�����xG�>��Q?�g�>��@?_�R?�u�=e�!���Ҿ��½��=��༉�?J[?5 �>�0�>��H>�3 �@m�@�? �d?b��?��q?�q?x�=?�[ӽƐ&?ާ�<
!?y?�{?��\?"�?2��?$	I?ڸ<*�t���;4�8�5�?9���=e��L�����K=��z�<iN	<� ��SF��X�Ǎ�	�=�>��>c%�>ౌ���B>i�Ǿ��c�.�3>���j9��Z���9���=�+>'�>�E�>���Z��=���>�d�>�� �t+$?X�?O
?���<��[���оFW���>�E?_>#�_�)����q��>Bgl?�7[?F��U辟�_?�\?�� �A��jľ3�u�s���j�S?�|�>�Y)���>�s�?��`?V�?Xl��Cm��ܛ�]�a�ԁ��=���>����\f��؟>�A3?$�>T�S>�.	>-�־+h}�����S?��?���?�=�?W�,>.l�(�ۿ?^��l���7a?W��>�J��]L?;�x�~=Ѿ�������a�޾���@���k���D׮��/����U4ڽW��=�Y?�di?�q?8�^?���h[���`��9�#�U�| �$�^G>��K���C�grl����pB�n���:>o=#Wr���H�-ù?�"?��r����>�P\�٤�Ȥ��J�=@柾�;��hl�G~Ž�x����U��%=�+�$�ZK����?6��>Yя>n)?��_��?��8=��k4���վ X>a�>
%�>l�>{��:�(�
��o��x�d��2�yno>l�a?XjP?A6k?5Y�j�2��避G�"�Ȩ��	��$vA>�>�Uo>�)^�h�4��@*��&>���n��a�}���J/�nx�=sN4?ˁ>�۪>��?��?� 	��δ��sn�&q/�,V.�x�>i?,h�>*K�>��������&�>aj?$�>w��>�G)�N��xD��OWj����>��>� ?l'B>l�����^�sg���p���4���=e<x?��}�^C[�O��>\JK?3h<9�=g�>�w����*��*6K�$�>,��>���=��5>Ё��c$���/r�}B��rj?#�&?Vq����(W=#��>
��>��>K�?�a�>��&���%>��*?�@^?��U?�;<?*U�>��=�d��ڭ����U��<F[�>��$>4&G>��L=��@�����ohͽ�Lp<�@�==�|�@I�t�c�6��=���;�[>�(ӿ_LO���Ǿ �5�P|�K40��%S��9&������b���ξ�_��E8���̤<qj�́�����N����6�c��?Qg�?�x��T���9�|�.u��{Lľ���>�q{���=T���	���޾4#�����G7��uљ�8���'?绑�˽ǿ�����5ܾP ?uA ?%�y?����"��8��� >���<�
�����핚��ο������^?Y��>�
�
C���>��>�X>�Gq>���0����V�<8�?��-?���>Γr��ɿ������<!��?	�@�A<?�2޾��8�F*k��;�>'?`!>I!��8��֤�g��>[2�?��_?�k����5��8��bF\?�o@>f�n�k��U��<8)�7��>��:�bi�>հ�=�#p��P����z��>��=���<��j�ϔ+�U��ֳ�>��=�9�4Մ?*{\��f���/��T��U>��T?�*�>8:�=��,?V7H�^}Ͽ�\��*a?�0�?���?�(?Bۿ��ؚ>��ܾ��M?`D6?���>�d&��t�م�=�6�x�������&V�L��=S��>l�>Ղ,������O�rI����=�F
��vѿ���-�)�8�D�\{K����h�h��h��i�s����I��[����>�h={�,>PɅ>�f>�nx>�a?�a?��>X3>=y�0=d��Ͼ�;�ʽ��q��̀�2ݜ��IR�����ջ����i��z�v�!��侲~(���=�'�J蘿�F/��l�������>?�Jo�*sX��~�z�3>z��s���;_S�����(����R�W�z�n!�?�)t?�������^Fƾ#Ǹ�>�_��Cm?�]��Y�D�̾�>c߬�/��>]��>��>����gV��d�"r2?jg?�;��9�p;>h�&�AX<"�!?%�>��"=z�>��>=�5�(2I��/��=|p�>;��>��\=�ľƀ���48?v9?Ჾtkq����>
�����û�h�=�:>(2C�z$�=���>�.�==)�=]B�=˵���jm?���>pk.�l���.��<"��ˋ%�h�?{h$>,`?�3�?Y��>�K��g��E�\�l�`����� ?�>�?I,>�F��@�4�����i?2?E?��*�A�;��"�;+�j3� ��>���>�p�>p�hj���+Q��H�h(?��v?�r^�vs��~��D�V��=�>�[�>H��>��9�{k�>)�>?�#�tG��𺿿rY4��?}�@f��?+�;<� �&��=�;?2\�>�O��>ƾU{��a�����q=r"�>����oev�����Q,�8�8?���?���>������M�=�������?n\i?W�.�饽/>�Y%��Vs}���W����=�j{=��a�gO��ߗJ����Yᾇ B���J=�%�>{"@3`�3��>�i���`Կ��P�79����)D9?M�>c�>w1*��%E��,�F{S�^`�X�Ͼ�X�>^�>|���0��5y���:��Z¼���>�o�I�>��i�����,!���\�;͐>�i�>��e>&�ܽZ]���l�?�F���pο�ݜ�K���[V?��?D�?'�?�@�<��y�j|�9Z�:�A?4�q?ي[?��;��,g�+?��Yk?�Ԧ��:`�_3�\A�;�U><P/?^�>O�.�/��=(8>��>ں>./���Ŀ�]������>U�?���?&\���>��?�+?�V���6;��Bk*�3��;V�@?��.>`Q��(� �[9�g�����?��0?9��r�]�_?+�a�N�p���-���ƽ�ۡ>��0�f\�/N�����Xe����@y����?N^�?i�?ص�� #�g6%?�>c����8Ǿ��<���>�(�>*N>dH_���u>����:�i	>���?�~�?Qj?���������U>	�}?V�>��?��=��>w��=�a����)�O�#>�=�=F1H���?(L?g��>���=pB:��\.�͔E���Q�[���C���>@a?_�K?�`>61����0��� �!1˽ w2�1�߼;iA���$���Z95>�S=>e6>��B��Ѿ.�?7c�:�ؿyd���!'�I24?���>J?2���}t���P._?QO�>,8�L,��s*���D����?�G�?M�?ǵ׾��˼/>�ޭ>mH�>�Խ ���g��j�7>��B?���?��M�o�i�>7��?J�@�Ϯ?�i��	?���P��Ua~����7�Z��=��7?�0�!�z>���>��=�nv�ݻ��X�s����>�B�?�{�?��>!�l?��o�O�B���1=6M�>Μk?�s?�Ro���g�B>��? ������L��f?�
@u@b�^?*��Vq��?ɾ��ʾ�w�?Ω=�>2�]�����*�\-�;����<��@>�6J>I�D=���=��a>ic�=�U���;#�����x&��h�t����6> ��L����4�z����m�^��ڧþ�Ê��� �Y���W��5�X���=c�=��V?T�P?{�l?�h�>���I>_����`0=��"�L��=���>_�2?�CL?Bs)?v'�=oϘ�O�a�E�~������Q��.��>l�J>��>���>�R�>��߻Y%P>�?:>��>���=}( =�,���'=>�N>5S�>[��>�!�>6m>K�I>�����¿��H��gѾ�(�� �?�8���X�����[��o=���<VP?�R>�ݶ��ҿ����y�g?���9'k��T��Ŭ�>�R@?Ө�?-ܾa>k�xV�>`�=�@��,����[��u�=Y��=I<���Һ�;?�^�>3�>���g�U��_C�=>��?��:>����cl��l���X���Ͼ"�=^DC=F��>��L�D��d�w��˖�1l>>GU\?' ?Vk��+���n^���/��с>�V>�$"�@8�=���=�$���Ҋ�� 0����<��<�'�>Ú	?MR�>r:u��2�>O�����y��>��>��5=�G	?��?M�z��$��{�@�����\>e��>/�:>��o�>'����,<�??���>nщ��H=�ż���D��m�>����p[��)��p�>:�ɽ¿�>� 3>T���r�I�
iQ��~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ	��>"M����������t�`o"=���>�yH?ޣ��KG8���8���	?K�?Ҥ�EJ����ȿ�?v��Y�>�8�?�ʔ?��m�w|��@����>��?��W?��m>J�ݾ�Z�Q(�>��??:cP?���>�L��A.��L?_7�?*r�?�6L>���?;Qq?�!�>�� �)�u���NpT=꽙����>���=�Oþ��I�������Q�g�z��؋s>'7=W�>SwｸX��y�=Z;��}=��7>���L�>��}>�B=>�V�>�? ?8�>��>L�B=7/�����*J���J?�-�?����s�I�<L,=t�J��y?�?	6�<�� �*ر>��S?O�y?F?�7�>Rs��R�����
 ��3� ��=W��>('�>�a;�z>/)��5��yI>�e�>̨=�q���֧�a�Vx�>
�-?���>v�=q?�=?���>�N�>ύ#���e�._4����>��>~j@?w�w?q�>�8���Q�����=l��N!N���>�z�?�#R?�z�>`���*������J��]�=A,t?W��>��>�)?nyt?�?��P?���>�
���c�/����>M�,?L����}���P�8��=��>��B?'E_�?þ3o	?�߈�?ܾ7���ݽw=?��L?�0b��拿C������|g=>W*�=�h��E�`>»E>�0����>��.�%�T>*����<ױ�=���� >w��>�=���I+?�>R�������=U�r��BC��˂>&.M>�����;]?�(8�]|�>R������~<W�M�?�S�?�0�?s䶽�h�I�:?��?W�?L��>$���e߾���=�y��\u���"M>���>��Q�%��E'��0`��n7��~����2�����>���>A�$?��"?B]>�>>�9�{��M���'۾��J���0��(2�+$�ݺ2����n�$���>����e������> �'���>}��>�N>��=��>��'=��N>�	>dp>Xpf>Ny>or>��=��<�,ǽ�FR?���h�'���辣4���JB?�Nd?�E�>)g��q�����P�?�j�?�Z�?f�u>�Kh���*��?�h�>���
h
?y�:=;d黖�<�߶�������I��xƎ>~,ս�U:�1�L��Wf�X.
??�>����̾��ս)���R�=O�?�S9?�����&�%�m�g�#��jK�v���7�y��S����(x��{����2��&Ol�����a=w#?Q�^?��оv������)�_�ftY��&�>�C�>�o�>d0�>i̬>���� �Է]���,�1��>Kw?��f>w�O?;�Q?��{?0��>�O�>��;�l��4?�u�=���>u��>�
6?��>��?�?�6?�ܵ>An<5h��t龗��>YF?��N??��>E��>�ý�>��{�n��
�=��s���qkC��a
�-ʔ�=A�Q&V>�"%>/"?�
���z<�F�Q�>�"0?��>���>���n�S����=R�>���>[$>��oH������>�x~?Uq�hI=�*>�e�=������T�=�q�����=�%(��fνؽ%<T��<dC�={�����$=Ȏ@�p;���D��h�>y�?���>�k�>(%���� �!���j�=UY>��R>�>�Lپ	v���'��^�g��y>~o�?�t�?�g=�E�=���=^���ih��&��- ��Ӣ�<�?�P#?jaT?Ð�?��=?�m#?��>�6�7B���X�������?�#?���>���
�˾���F=��?�3�>�L��Dʽ(+��߿�m_ҽ���=j�+�Z�P�i����N���u;���R%Ž���?�'�?�Y�<12&����ؕ��e��>�8?��>�,�>���>�6(�c�i�O	2�E�>�	?�S? �>	H�?���?1;?���b^`�7���S�H���>�j�>c?�g�?���?���?�$?�Pe>}���~Zy�7���+"b��==㕮�T�T���O=!p�>��>�?x\>Ma����S�����|�=p��>M�?R��>3��>�G.>Θ����G?�F�>z�������٣����E?=�n�s?�Տ?��*?���<�U��OD�R?���k�>��?���?�(?5V�͢�=���񛶾1�k����>���>���>��u=�<\=Y�>���>�>�,���T25�3�<�3�?��G?&��=�4տ�녿X�t��]�����������O���j���6B"�������w������B�q�W������[�{��d6�n|�>s��=5��=8ˍ=&��<��?�q���=^�8=s&��Ƅ����=nm�<*��<�����a;��=G�=�d�<�����M~?�T*?��?��=?��>'�g>_����	�>G �n�?�=%]y=���������n�����Ӿ/];�gW��h���6>��ʻ��=��=�HH>-n��%\>��<bP�=ۡa�7��<�>,��=���=��=�s>�w=�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�ؐ>��:>r�N������"�ֽ��5��ڱ>����
�c�>/sP=�^��徧���&==��B>�V۽� b���{�	��<NE�=X�J�/,>�=�x >��� �W>�r�<�]�=�%�<O�=	Ib����<,l>y�˽���>�>S��>L�?}S0?��d?ɕ�>f�I�ӶѾ������>QK�=���>�y~=�F>v��>%o;?��B?2�H?Φ�>�6�=���>Ţ>uX$�nc�qs־s���^�<S��?�?���>_��=IS0�����=��4�\�?Xe/?��?��>_S��濎�'���D�}���x%��,�����Û�f�i��ɓ�5䓾��X>l��>�"c>��>�>=��>��\>:��>� �=��=vzM��/I�<�t�=�Y4>>��=i�>�!>+e�=#��<)7�=w� ��K�=�ͧ<�;+����=Bq�=���>TV>���>j�=Y	���2>pj��/7L��=� ���IB�W�c��'}���.�Á6��IE>�8Z>?�����('?Za>��@>l�?�t?�I>���K2־ђ����k�R�r�=�E>S!;�̇;� S`�h�M��}о��>�m�>ӿ�>��>�p��|0�3vQ�+���A>����>۽T��N��޾m�]����*`����V��s[���O?3�n�I�[�v ?��K?���?�?iU(> 6��f�:>�g���y
����Ġؾk��<"?̮�>F0?��ľ�w2�p̾�J��� �>#�H���O�����|�0�F	�{����]�>�Ҫ���оM,3��e������I�B��{r�̺>/�O?�خ?7�b�r=��4O����XM��@w?7Rg?��>�E?�;?.S�����<S���|�=6�n?��?��?!J>�S�<�'���B�>ЇB?nB�?�í?��?wyk��R?�b��i�>�?��<�=�U�?2f>�Q<Y�%?��=?�&?u;Ž�E���,�T������.:�m�=R��>k��=����1=ۼFH>ia>^Q�=���>)h�>wƫ>o,��9�;�S?$�e>��>�?l9�>\E<+	�����Ͻ$˞���ྱ��h3�Ԁ�tX�:�ù혩==�>e�ǿ�-�?
�l>ϒ���?k䥾��D���S>H69>�I���>0	>s�A>��>�>�(V>�xF>K�m>���v��=
|�S�1���T�i�P�c����cd>x㝾l� ��y-��߽�����=������\�c��聿�8�N��	�p?ӳ���&��c��cȇ��^?1V+<& 0?����g��5�=/�>��P>X�9��1���=�����$P�?7\�?f)c>�>@�W?Q�?�<1�g�2��sZ��u�$A�Ee�9�`��ۍ�����
������_?��x?~nA?��<�9z>>��? �%��돾��>�/�0#;�d;=�]�>㰾��`�i�Ӿ̂þ�}�+�E>M�o?��?S>?i�U��7B�h�B>�p7?Ì1?��p?pj+?b*;?����6'?�>�r?D�?'o9?!)?p?Ǜ:>���=���;2U=5V�������ֽak�����.�]='ca=Ż���J��<���<t�üE�D�� �<��*���;�}6=��=���=Yͣ>��\?�\�>���>�*5?����4������.?�$=q�l����I���o��!>X$g?�"�?ybX?��f>�UE���F�с>�Y�>�4;>d�^>0��>�콛�;�	 =K(>��>�ө=����Ԇ�w'
����J�<
�#>�X�>H�>Eڻ�t�=9���������>�xv�'M���s����I���7��P��XO�>�?�?������2�2�
|c����>a^q?`[w?M`|?��>'#��u��b��K�z��>�\>p�}B��K���#4_���=���>]����ǾuZh>���S����q��qO��N�寮��?�<�2�_�������3ݺh}=�޾��8����.D����P?.�=�X���bs�99¾���=־�>���>6�w������7��Ɲ���r=h��>��->~޻p��%�@�����l�g>��Q?N1u?�Ç?�P���o�بc��(�\�_8>��4?�"�>�?�^k>h��=2����ھ��G���H��n�>��?l;��S��с�8��VH)��֏>8�?)�='�?߲I?���>�7K?W]?��?�|�>@\��Ŵ�S�%?��?�{�=ͲҽyT�t"9��zF����>�)?n�A���>I?�?��&?PfQ?7�?�>9z ��b@�䎕><��>�X��Q���g`>OGJ?���>�&Y?#��?-;>ט5�	ע��˩�Q��=�K >��2?��"?~?��>�s�>/�s��̇=�6�>�E~?���?=�p?[��=@?��D���?_B	�2�?6?6i7?�w?h�w?(*F?�p�>'�@���G�p5.�^���6���`=Y�<�1�<. |=`d��F��8�6�τ=��*�� ��C�;����o�C���M?��W>@T��>�C>��_�f����>%;��N�k�D$��_L��4�ME>�R�>(0�>d*+��I��r�c>�8�>Qy�Ω�>�t?�n0?O� �,�5�����'��>s9?���;G=��~�R
@���B>�2�?��D?v����;A�UCb?�]?v��ܲ=�"���.a�F边�P?ͺ	?�@J���>[E?�yq?v�>�i���n��ܜ�\�`�0�e����=�{�>�q��d�Ag�>$7?��>��a>ĉ�=��ؾ�8v������k?6ƌ?��?�<�?�,>'�n���߿y���}��0�Z?�>S�~5!?�	���Ͼ枊�����ކ��ת�=u��[}��ٳ���%�Y���/�š�=�?ƭr?W�o?8G^?�� �eDd���[�`���zU�������� E��$D�D��0o�����󾫙���wF=�ǁ��h4�x9�?��$?�>d�5?�s��h%��G¾��K=���_`�=fA >M�d%�=�-�<o!���u����!?���>1�->��'? ���gJ��w#�j%���j���>�T�>���>d��><�ͽ,F?���ؼI��9&�̃�=!�t>�6c?LL?��n? }���0��l����!��A1������A>��>P��>��X�n���%��$>�qr����Mɐ�*�	�ïy=l2?��>$�>N!�?�?-T	�&z��E�y�p;2��?H<��>U\h?ry�>ϔ�><\ѽR� ��H�>�Pg?��>:·>������ ���i��uD����>qs�>A��>4�&>g�q�H�d�雎�����d�#��V>�v]?�z�������>yF?x��<m�=<�Ǥ>o����~0���j/�8�1>xr�>���=�">�ھ�1 �)��������)?�?:R����+�bMc>ݛ?I~�>��>�T�?���>Jy���W�"O?bvd?�	L?��C?�w�>���<u�꽗Q̽:�&���O=�N�>��J>�6Y=�=��!�dAi�~���6�<9��=�>D�m5ǽ��;�(����<�̡<��">�Y�|�S�CKо2�qLܾ<b��Z@���[�����}�ؽ����拶��ھIeξ~o��ղ�����ݞ���e�?r��?�՗��¾���C�n�3-)�Vٓ=`���D�=�x��a��
a��\�����LP�}S��������N�/?mƚ��:ÿ�"��wȣ��8%?�?�N�?4���&'��|'�
�P>q�1�����Ԁ���ƿ�WP�̻m?}��>Wkﾪ�����>U|>�>�qi>�����|��+�<6�	?��,?�t�>�����p��\�����=R?�?O@��C?)�>���8=��>�^?gCA>��Y������5'�>{ў?~ֆ?���=H�W�#F��Q�_?Q�R=��7���ɻ��=���=��3=�@��T>�'�>�)��18���ֽc}B>�z>$��I쮽B䀾��<`i}>��F��6��ڥx?�x�y{-��!(��K��[�x�
By?{�>�S�<ې|?�s���;��!ٮ��W�?���?���?{bC?���������־%6]?�z*?E&�>*� ��q�&-۽��Y>B��={۾)b��9�����> ��Y;ɽMz�H���
�=���=�����ݿm��d-����_UI�s��=�}W��}��e��lžn���h�C�^�<��V<�q�>#Τ>���>�n�>�CZ?�[?iN�>k�=���=��u��R��pc���z�����������D����}� ��?�(@J�ZB@�(T�c�z�p	S�~ >�nS��엿UQ6���q�GF�?i��ZGؾ�%j�>�ƽ�����zBx�*<���&��jD�B�0�j�?��#?S-���@Q�?��= �;9� ���W?�*:�?C������p=[��4Z�=O��>���=�aԾK�%��7A��@?��#?|׾q�����E>����]>y�??���>�����>�� ?p��Ž�R@>� $>�Ru>���>u��>㧾���S-?��N?�ɐ�,���k>�, ��Y[���=I�=R3����7��>
�1<N���A=��*��jн�g?�Ҁ>y6������P��ό�	$^>��{?E�><��=��=?�?��<��ھ��N��
��M��>�2?��?`j@>U�S�k0+���Rg?��<?�@�>$7�=ӯ4���L���߾�?�>h|?�/�>�8?�@9��3ۆ�e����~.?Z�v?^�V�Ou��M����F=��>��>9��>&;����>J�=??" ��	������5�G�?a�@���?�_�<'k��y�=��?w��>vZ�6վ	�h�̽�=ԫ�>���5r�x���i�4�=?9��?^��>���/ �݈=E�o���?���?�&����=/�B�r���Ǿ<t'>�iO>�V\>�%�=�*��_��
1��<���H�6�
+�On>�@������?<������j�տ����:�$S�=/�=?.Q�>�9���Gk��#h���9�q��	9<��q�C]�>2(>�:�<=�����"�t}�=2=�>�*J>:L�>�Q���_�����	rؽ��1>���>q�>5%�����:�?��^K￰��������?�ɠ?`A�?V�?u���C�<�-���=Dap?��>?%�0?�=?�J|W��5>0?t?����\�P����[徑F�>��:?��?��>�ʶ��P�>�"�>�c?=f��VYĿ]몿����r�?W�?K3ݾ�R?���?�?�  �C���l����E��'M]?��=Ջ ��L��.�c��VP��D?(?�?e̻18�O�_??�a���p�p�-�M�ƽ�ڡ>��0�%e\�~L�����Ye����,>y����?+^�?H�?��� #�75%?U�>����8Ǿ�<\��>�'�>�'N>w?_�T�u>����:��g	>l��?>~�?(j?ݕ������W>��}?d!�>u�?�	�=#v�>��=o,����%�>S#>@.�=��=�b�?ْM?:�>���=ݶ8���.��8F�;R�[�l�C���>P�a?܌L?�b>W~���3�{!�ԣ̽cT1�5l��p@�~}.��i߽J�4>��=>�I>��D���Ҿ@�?;��"ҿ<Ӗ�t*����1??�>�n?J��mߍ��A:�7e?=a�>i�*氿����^���:�?m�?R�? �߾�4��T�=k�>�ނ>��ӼA��!Mp�Kjc>�D?��<���z��0L��>���?�g@A�?=b��	?���P��aa~����7����=�7?�0���z>���>l�=�nv�̻��X�s�v��>�B�?�{�?4��>�l?��o�F�B�g�1=BM�>��k?�s?)[o����B>��?:�������K��f?�
@vu@*�^?#�(ٿ�c��\*¾�鳾>G�=o��=j%>1"��B��=�y�<U�1���&#�=�3�>�n>�Q�>[�\>q�>>�� >���{�&��竿h�����M��w�֒���}�m3��B��m������V�Ǿ���*a���T�9�A����aV�"��=n?ߡJ?/��?v�>k�����=���~rn>��V�K~_>��>�r7?АU?:�O?I�>�kC��\]����m���~�j�X�?,�x>Fi�>(��>���>I�K��B>�k�>Z��>+xO=��]>#�v�	,Q='�d>���>�Q	?�:�>�=(><>�>��i����i�hk�_���5�?�����I������D�������>=m�?�%�=@S���̿R����:J?����1]�};�$w>]%B?7�I?�#>�%��f˼�5>�` �#�~�lL�=K�����L��N �IC>�_?u�v>%�=�>�>�>��X�!���E�j>y?�ܓ�?��m)j��;�\�
�9>��u>31b��A�_)���W�'���#�.>�4?�?�^/�4,��8��񰾘0z=�pN>>���8"L=NXu>�Z?�/�S�,���%��=��>�!>~�
?��*>0�M=ל�>\����QN�#��>9�3>R�">�8?��?�����f���{U!�&�>�~�>��>��>�$k�Ѣ�=�I�>C3�>%1����!�\�����o�>����%o���*�9><�E���;>��>[�޽%�V�����~?���'䈿���d���lD?R+?� �=O�F<��"�? ���H��@�?p�@m�?��	�ڢV�G�?�@�?��9��=}�>
׫>�ξ�L��?��Ž-Ǣ�Ɣ	�)#�dS�?��?��/�\ʋ�8l��6>_%?��Ӿ��>_���aS��m�x��|@��ذ<v>�z?�������\[��?,|�>)K�k���>�����s��~�>�3�?���?�&m��{��N@��)4"?�W�?�-N?�԰>/U��2R�*c7>��'?|_?�c�>�ˁ�b��"]�>T�?\K?G�H>���?R�s?��>+�x��o/�j8�������=��;���>*>j���kIF�B����Q����j�����^a>�~$=�_�>���(:��:|�=HW���k��Uf�<ķ>O�p>�`J>�j�>\� ?Z*�>�V�>��= �Ҁ�����5�K?���?��8�m�#w�<��=k`^��?�[4?�o[���ϾŨ>Z�\?���?$ [?̨�>"���6��&㿿����~՘<��K>�k�>O�>�ǈ�9�J>i	վ'�C��u�>���>�����پa큾R2��k�>��!?oj�>4H�=[w?N�"?c�b>�ٲ>kSF��됿�kC����>�>�K?�{?�?	����D4�咿&����QY�izT>�=y?>B!?^�>2o��i���o ��\	��C�w�n�?i)]?��j�	?栆?c(>?�[@?�rW>+�@%ܾ����M<�>d7&?x�!�>J��gF��u"�>O)�>��>�ζ�n�?�t�=a���־�?\�?pN�>�յ��b���� �@=��)�Xk�=���<:ژ�S[��f�>�)�� 'Z>u�E>𫽺�����]��&�>$��>���>z��>��L���޾� ?M/�=���?�M>�S��5.��*R>.1�=`�cj?0U`�m,~�1T����������)�F?)��?-�?�R=��z�G�0?�4�?�7?m�d>�)辚�k�5�~i�=�4��d��d���lp��x���`̾�ƺ��}C��ź'�l�C� 2�>z�
?F�?E[
?�>)>Y�>���E�9�����q>�T!���<�Q>$��������$�h���!���H�� ��>�AA���>�?b+>*\�>�>+�=�X:>HQ>��>m�>�>��W>d^�=g����<��H?����v-�����A��-?9r]?9?i����s�B�ܾ�,?(��?%�?Y�>��a�\�$��4�>!i?����>)n=^J=�J��ٷ��ٽ��!��S��n��>`g��`���,�~R�(W ?}�2?�-s=�M��zT�־ž���=Q�r?؆,?v��l'a��p� Q�#�M�^�|=�X2�-���tf3�	�v�cs��U��t�x���|�}=Y�!?�z~?���L�Ⱦ;�����S�ֳ,�� �>#$�>ZX>���>-܄>��꾟�'�9q��c'��U^���?{?.>��]?uai?Y��?T�?R�>M=>�l�3'G?=��=f3?%?9�`?M$? �j?��e?v*N?B�>>R���\l	��2��l?�
�>��?N?���>��`�@����I=��b�+���n�iC׽C��\@��/��B�?��?r�G?��Um[��U���>@��>�?N?pӾT�߾)A�=��~>g��>c�=�־#0Y�Mq"��I�>D2�?�b;��=��.>�7�=V�<�t�=�x>gcp��>� Y=��P���=�F<T	u>O�>�ټ��">M�>�X=y
�>��?d��>�Ɖ>�f��I� �4��)ʬ=�#[>$8T>�/>�پ)r��*����g���w>�l�?ȃ�?�h=ٯ�=��=p����Ͼ�z��G潾þ�<8�?�#?��S?*q�?��=?�"?f>�$��Q���z�������H?��%?Z�>�M���Ҿ�_����6���?$�>m>^���Y1�j\ľ.V���=��0��x}�<}���C�J�'�N���O�B��?5��?ߺ�J>�@N������𹾨k??�Y�>}j�>@��>{-�8�a�E=���5>��?J?��y>r�?�t?l:?/�>m�X��?��I7c���>s�;<nB?n.�?߻x?q�:?R9'?���>푅>6��m�H����M��H'پ�~���sM>O�$>t��>���>O�=
���\L���Ƚ�Z�<��>�'? ڭ>�N�>����򔽫�G?���>�`��Ë�5�d˃��J<��u?��?��+?�e=\{��E��7��s<�>�i�?��?=**?w�S���=�gּb�����q��2�>ӹ>�,�>>�=C�E=�%>Y	�>l��>�4��\��l8�<�M�h�?]F?��=N��yM\�4��b[�-��<F$�ڦ��qiq�����B�=J럾��w����¸���l��pզ�|����*�K��e{�>��k�,˒=� 
>b�=N5�mW��0=�,�<xv�=ݟj���{�ɭ��m��<��>X=�X�=��3��o��ѾU�q?�dX?�2?��P?�e�>�e�=�ʽy��>ݫ2����>�kD>w���M�о��������h���+ξ����WP�(���Խ�=EƸ�?�>��?>;�>q�7=�9>+2=/�:�Qp�6�N<3'=�-�<�PL=��>�}�=�>�6w?W�������4Q��Z罣�:?�8�>c{�=��ƾo@?~�>>�2������wb��-?���?�T�?<�?=ti��d�>P��{㎽�q�=a����=2>a��=��2�X��>��J>���K��H����4�?��@��??�ዿϢϿ!a/>��O>w=��o�y�Y�������<����^�$?�A�G W��H�>���0�3������ümJO=�x�����}���=8�ܽsX�=O��=|�T>@
>�H>f�[��C>X)v=$x<>˩K>C�<IM1=��=b >�J>�H>�Q�=���>�?[�-?Ҝq?8̧>�`��BpǾ��Ծ���>dQ">�L�>b�>�]t>��>*1?��@?��F?8!�>�`�<�{�>XD�>�-�P�^�I�Ծ�?��g#�C��?�?���>E?>? ��p#�)�5��)����>I�#?lC?��>���2��%��O/�"s��3r(��x[=q�x��7���H��S�����j�=�Ĩ>H}�>���>�>P�>>�2R>�"�>�I>#�-=�H�=5��;�M<�uD<{�=5���<���|M;�K��Cr�go��t��ѻw�I<Z%}<l
p=���>O�> ?���=����^T�=�羘�#�W�=霡���(��pc�D�~�w<%��`�g2>���>�ء�W芿���>]�y>�=���?�+h?pF>-M��!��c����w������q�X_�=m[H�6_4��j���K���߾r��>z��>��>r�X>ٮ)�c�T���;#Ⱦ7:����>�"z̽EMF�p�m�⪜�x����V_���<��.?�֓�5�\>�<�?��?�7�?���>%o��aӾ;C�=1ܽ�ك>E���X��>� �߮�>?Z�>�:���'���Ҿm^o����>"�o��^P�b����-��\c;5ܺ�p��>�þ!�̾�u5�:冿6A��@�C�Dk�����>ZN?���?m��h|�UG��L��y
����>�$e?��>�?��	?�l����Ѿ�"O�-��='{g?`9�?0.�?�(>m�e��x�:^��>{?)��?��?[�a?��_��	?e�B�nN�>$��̤>]D�>Y��>��>�?��?�]�>���z	�
�����@.4���<���=f�>�p>�O�=��;��L�o��=�>x	>�8>��8>>���>0���@��pR?ݳ�=��>M�:?	�+>��p�j��Q6P��SԽE�ٽY���k�Ȫ�e^;�~>��.�rU�>]3����?8�=�P����P?��о��U=P��=D�=���ڦ�>)}�>	�>dZ?�p�>ؘy>���=|V;d� ��I�>�<�����D]��k��P־>d���~.>�������6ξ�$�]`;�?�o��A��3��e�y>�?)� ���N��'2�s�ֽ6
?���>��?�����wϾƍ��B�>>??*R�$����}��7�;U�l?���?"�b>��>��W?V�?p60�p2��^Z�֫u�n�@���d���`��Ǎ�����O�
�����η_?�x?�SA?W�<�Mz>���?��%�����<�>g�.�?�:��E==�#�>���Fa��ӾO�þ����8E>2To?��?�=?�U��W��=�@?a)?�8�?�
f?{8?��K��� ?����?S��>\�F?+�:?�]?�k�>��+>\h�<�\�A�νXu����
ZE��`����z=G���}!��t�����=D�=;�K=!ji:8���je�<2�;��@=�b�=�B4>lv�>��`?���>4�>�8?�	���1�Vo��g6?�Ӄ=�>L�1;z�T��� ���$>4Yp?䌫?
IV?]�@>
�B��E�p�>mXw>�b">��m>���>��׽GS�Y�W=��>��!>&[=*m_��l}���D���'��=�X>��>�+�>QI1=r�>�:#� ���>Y>R��y��bP=�X��I�U^0>���>_�G?[*?��=�Ӿ-F˾���ZpZ?�k-?%�?�w?^������<��� ���1?��>,R��5���̎~�b��`
>n`�>23��H��1Kf>�,���ܾ��f��rD��V侬��=����PI=>��Gž�ms�wa�=w�'>�松������FI��b�E?q��=~N��A5�NE�����=��>/�>� ���R��=�������8=SM�>g�P>3͆������U�H��7��>Q;?a�h?Q��?��X�E�r�V}M�!��OꜾq$=�|'?�ɥ>r�?f@�>4<�þd����S�u�@�Y�>�n	?�2&�I6K�E 0�Mt�rQ,��>z>�^?��C>`l?�S?��?T+n?�	7?���>`w�>��,?�bj$?Fe�?�N_=L�ٽ]�Z�gL7��F���>,n(?k�8�KN�>f?z?�=%?��O?�?�>Z�����?����>ẙ>J�X�RX��-i]>KJ?�Զ>��Y?T
�?f@>4�1�V����դ���=YM,>"1? u ?ls?{)�>���>����A[e>�)?A/�?�ĉ?	�q?��=a?��?��1?�K>��}>";?q>?c�-?�S�?9b[?��>�h_��0��3��7��%� =*�^=�=�2>(�#���^�t��w�8�Ц����%=:ѳ;q������\�<���o>�>��s>���m�2>j���}�s��k>�{�<۫�Bo������>��a>�\�>?�>�]��z�=���>
��>7��4�?�J?;Z?�q���j�f�׈:�5��>�/>?���=�Te�I�����i���.=�lT?Фk?�2�=��M�b?��]?Bh��=��þ��b����d�O?6�
?-�G���>��~?_�q?C��>��e�:n�$��
Db��j�7Ѷ=cr�>GX�G�d��?�>c�7?�N�>-�b>�$�=u۾�w��q��^?��?�?���?�**>��n�O4�-V��Rԑ��]??��>�N��� #?x`N���Ͼ�����`��	��7���������Ӌ���$#�
���Q�׽A5�=r?^�q?9�q?�`?��5Md��^�U����W���kF�0�D��pD���B��n��j�������8=�]�i�b�y��?@�2?8YJ��-?��������{���p>C䆾���(]�=��\��݋�[�=��`����[f��?�d�>��>�3?�@���2�o�9���;�&����=�Ħ>���>�o?��=�W��g轒>��r���H��*u>4c?�K?;Yn?p��t�0�p���̄!��P2���ɒB>�)
>���>�W�/+���%�\�=���r�c��i����	�[��=��2?WB�>4��>r-�?)�?��	�n;����w���0�߸�<v�>Ȝh?��>��>�ϽU2!�Of�>��l?zA�>tܠ>{���N1!��$|�U�ʽ���>�ҭ>̀�>�o>u�,��\�;\���a����8����=gh?%����la��B�>�2R?���97<_�>��w��"�%��
Z'�b�>��?���=�:>υž,���|{�����?)?��?@ߔ��+���{>M�!?r�>�/�>�c�?�֚>5�þT�@�x?�^?�vI?%�A?L7�>�=�	���EʽAs%��&#=��>`�[>0�u=+C�=Ȕ��=[���m�H=Dy�=B1Ƽ
9��t<N�Ǽ��><�=�7>>���!�S�{觾��n�����k���J��3��o ۽uT���(۾�:���c۽��.�=]�{Y��5{��K5�d�?�@�?m���o/þ����݄��#����>�0־ �f�[腾}0�`��NQ8��솾��`\�����^o�o
*?_Y��C�ſ�_��{�ھX�?�	#?�w?w��c�#��8�=>�l9<7c���߾����Ͽ�*��D�Z?F�>���X���=q�>j>
 M>�ƃ>:ё�����zO�<Bu?x�#?���>�o���ʿ�N��� �;��?��@[/A?DE(�?�쾥S=s�>4A	?]�>>B#0�����~���S�>Q�? ��?�GJ=��V�s-���e?M�-<Q�F���ֻ�j�=���=��=�'�A�I>n�>����i?��׽�|0>��>�"����X�\�o�<��\>qٽ�㔽5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=r6�����{���&V�|��=[��>c�>,������O��I��U��=���ҿS,�������<���Pj���/ڽ��c�8�L<���KO���F���>و�=��>���>��}>*�\>�
f?2Mp?�9�>vE�<{��˜�T�Ⱦ٠�=�+�����7�@��^��- �:`��&/�ա+�h�����a5���>g�!�菿)�C��l���2�c�L?3L�� ��dS�@��}Uؾb��g�=W�ݼ]S�� ]N�
"��eק?�l"?
熿Tgk�$⪾4�M=��<.P�?D�=V����#�H�d>'\��C��p�>8�>K�}��{��:���(?ֆ?�nȾLYv��w >�D��-�=��#?���>�X����>�&?�D �o��uT>���=�͡>�,?S�">D���;
�O	?�U?,�%�mQ߾{$B>�p��(��Y�=G	6>��t�c�P�.�!>�_�:Zv��D}>���<d$�CFF?G�>r5�%`��ޛ�v�A<�[��_l?�E�>͏�>�
Z?FQ?/E�=��� >�:��@��=�Ke?�e?mu�=MǼB���~����B?�s`?H��>�HϽZ����G���?d[?���>�19��p�Bt����龋	N?��v?Lq^��r�������V�\;�>zX�>���>�9�Nn�>�>?#�G�������W4�j��?x�@^��?�Q;<�"����=�8?U�>��O��;ƾ�~��C����q=2'�>d����cv�F���W,�v�8?#��?��>ș������B>؞꾽w�?��?������=7������۾���=Z�^>ֲz���=��6�S�Wޯ��j��s�@�=�I5>�c@.�����>��=Zq㿭�ֿ�l��y��M�_�� '?�̰>�>�=u����KT������7�1��S��Y�>�>�˽�����z���7�"n�q��>�+�÷�>�^��[������Ҽ[��>W��>^;�>v��o�վ�T�?ɰ�`̿1�������j}U?�+�?+��?�$?���<T����:����ܭ7?{0q?|]Y?Ǎ�n@ �t�<ٱj?K5���J`�y4��0E��fU>.3?	A�>�-�05{=)>R��>m~>�/�sĿ�Ͷ�"������?vy�?�Y���>�v�?�+?�f�^A��}H���*�+����#A?�2>������!�=�g���h�
?��0?���UQ�]�_?#�a�M�p���-���ƽ�ۡ> �0��e\��M��!���Xe�
���@y����?J^�?h�?��� #�_6%?�>\����8Ǿ��<���>�(�>*N>�H_���u>����:��h	>���?�~�?Nj?��������U>�}?�#�>K�?�_�=�^�>#`�=�찾q%-��m#>%�=?�ߟ?��M?mM�>�L�=��8��/��YF�ZDR��!�y�C���>Y�a?,�L?�Ib>m"���2�;!�xͽ�c1�z]� T@�k�,��߽�$5>k�=>�>��D�jӾ��?�o��ؿ�i���o'� 64?չ�>��?k��E�t�F��<_?�z�>�6��+���%��AC�H��?vG�?��?��׾yJ̼\>y�>H�>��Խ��������@�7>[�B?�!��D����o��>��?�@�ծ?�i��	?���P��Ra~����7�V��=��7?�0�"�z>���>��=�nv�ۻ��T�s����>�B�?�{�?
��>�l?��o�P�B��1=1M�>˜k?�s?To��󾉲B>��? ������L��f?
�
@}u@X�^?(�hֿ����_N��O�����=���=Ԇ2>�ٽ+_�=��7=��8�7=�����=s�>��d>q>A(O>�a;>��)>���Q�!�r��\���S�C�������Z�B��Xv�Yz��3�������?���3ý�x���Q�2&�+?`�@2�=R�P?h�S?ufo?�`?������
>s���b�<�5	���=��>8?:�V?��,?���=m
��Cp`��ˀ������7�����>N>��>!�>e��>k.�<�#.>>��>��> �c=��I�.!u=��O>�8�>u��>��>qZ�>FF�>���gզ�IM�����4�ܽ�O�?[)���h�Dm������վ�W��`?)��>m���7�ѿd�&?�X����i���.?>Ŀ?�o2?��7���޽q1	���>�~��*�>�G��>M�L�ߘ;�QYD�~��=��!?	�n>�˶>WkF���A�a=��ׁF=%�$?����]Ƃ� $n���R��N¾�h�=×>��>E<��璿�`��R����=�T?�?4���I��**:��ڼ���=!|�>L�>����e>��n��H�/���x�=�)E>w,t>�� ?��>�\Ӽ�Rx>�l��^=G���e>r�=>~>�D<?�G�>���=BN%��Z���l�4>�L0?��>u��89��5�<i��>���N*˽�$�~)R�����Ϙ>0X!>!������=��8�]�>�s>�����P徊A�9�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>wx��Z�������u���#=P��>�8H?�V����O�e>��v
?�?�^�ߩ����ȿ3|v����>W�?���?f�m��A���@����>:��?�gY?uoi>�g۾>`Z����>һ@?�R?�>�9��'���?�޶?֯�?I>Y��?.�s?���>Uw��`/�\7��R����=W\v;#��>SX>]����1F��ؓ��f��K�j����W�a>G�#=S`�>�X�[T���ķ=�Ɍ�>s����f����>�aq>�I>u�>�� ?ŧ�>��>{�=�Z��Zր�k����"C?��?d/(�m�{�;n.��X�=�]����>a�U?yƽ+��1�)>Q�O?pdk?�|>?׶�>eh�wj��97���{ɾ�K!=�-�=�|�>.5�>Zo�ܼ>��վzG��Ź>���>��;�v*��礋��E�<P�L>�?���>Sn>�� ?g�#?�j>�)�>�`E��9����E�
��>A��>8I?p�~?��?*ӹ��Y3�����桿n�[��;N>�x?�U?̕>x���ო��'E�7KI�������?=tg?�O�?22�?ω??ݥA?(,f>����ؾѨ����>F�!?dFѽ�D��+���h�?E��>�s�>޺뼅}�퓜����8���2?UU?x�.?���Uh��Ⱦh��<.";�����;����D*>�H>:�ؽ)��=�>Bx�=
(e$���a=`U�=���>
�=H'-����;,?dQH�i烾ֺ�=��r��kD���>4QL>	���-�^?��=�v�{����Ht���T�X��?x��?�a�?�c��Z�h��=?��?<�?��>�J���o޾`�MIw��x�N��U�>���>�cm�`�����.R���Ž�v<����>���>�x?���>�G�=$ ?vi���� ��,�þ&lw��@1�t���4���)��㷾�d��[=@�꾊����Y}>lDy��{�>��?=>gŅ>���>�=�{_�>j�>�A�>}up>�߇>f(c>���=������
�Q?�"��;�'���쯾ЯB?`|d?���>.x|��J��{���?�.�?��?%�u>�	h�ղ*�W0?�7�>4�~��S	?F<B=[Z,���s<����5�G��n%�{�>M̽��:��N�D4d���	?3A?Z�:��\Ⱦ�U�(���4�n=P�?�(?��)���Q�
�o���W��S����r�g�6a����$���p�j쏿p^���#����(�� +=-�*?��?r���0��+k�m ?�:f>
�>bC�>�ʾ>�I>\�	�5�1�M�]��='�i����E�>&W{?(�>gXG?�'=?�{P?��L?=��>ef�>�!���;�>S�<��>s��>��;?��2?�1?�?W*?(R_>?�}���5�ؾ�?��?|?��?"X?h��4Pս����^���i�M�m���f=D�=1ν=]j�(�H=��I>�?Q�=8�D�Ȭ��5> :^?�K�>�@�>�� ��A�Y5��ļE?��V?�;j;P^�G!����ZK�>s�?�ɤ��Ec��Q>�ܕ=)v�<�p�=�É>Z���Z"w=\� �aOͽ��Y�i���^mA>;ӽan＾D��5;��<Et�>��?莊>�@�>UA��� �����d�=�Y>�%S>�>K?پ}��>#���g�+Wy>y�?�y�?��f=��=7��=F����Z��_��1�����<o�?�J#?�YT?�?{�=?j#?~�>&(��I��]������?�7D?"��>�(ݾWG��z叿�vO��'8?�c�>��v��$?��3�Kp�a�|��R>��P�����#���-K� I�=(�������?�]�?�^��V`�c�׾���"���O?�L�>:�=.��>X�&��>����V��f{>]?�sW?�6�>s�/?/
?(�`?ȱ�>6')��Ҧ��9���-;6�>�6a?�v?͙?$�?�c�>�Cp=����<��7F"�I��-䚾7z�E�>{ʨ>v/?���>��=�$2�f����8�<n$>L7�> ?�g�>M��>N��=������E?�q�>\�¾N����pZ��?d�#]s?AP�?��+?�}=���u�A�X���%��>�G�?��?)�)?�JV�9��=pƼY�ۣt�'��>ĺ>�z�>���=vXG=�Z>?�>y��>�I��d��G3���G��V?XF?T��=&�ſ�(q��Wq�����/XQ<���Th�u|��x�[�z��=�����l��A���7\�e"����������Ϝ�0}�$M�>�9�=���=��=(Z�<ּ̤�7�<fK=��<��=�4o�;��<��-�>���ň�y��F�<��K=��8�˾��}?�;I?+?9�C?��y>,:>��3�䙖>�����@?sV>ƞP�∼��;�9���M ��5�ؾ1x׾��c�)ʟ��H>Z_I�L�>�73>�G�=�L�< �=�s=�=6�Q�=�#�=zO�=�g�=���=�>�T>t2w?喁�����V/Q��{�y�:?>/�>y��=�lƾ�!@?P�>>/+��}����c��'?K��?�T�?��?��i�le�>����R����i�=ڰ���'2>{��=R�2�0��>��J>���G���0���+�?4�@i�??�拿�ϿO^/>E�=��%>h�N�FV7�����#�o�:�ʾb�.?�������?�; ��=mQ��� �>�2=Qj�>�Ud>�`@�1i��['>�׶��=�#�/=*�L>�S>zoq>>�$��+>�7�=��=V�>?>߭<��C=IL>3ƃ=J�}>�Ȍ>���>T�?o�)?Q,_?��>պk�'nӾ;��-�>��='��>$�=��J>��>75?��B?�O?���>�@X=R�>N'�>l�.��Om��⾋3��'=ݪ�?[��?��>�;<�
,����Iw;��P����?�W-?<�	?��>�U����6Y&���.����4�4��+=�mr�vQU�f���Qm�|��u�=�p�>���>��>JTy>+�9>��N>��>��>�6�<p�=iꌻ*��<� ��޴�=7���.�<�uż�����s&���+�A���ߍ;���;{�]<���;a��=��>dj>��>�t�=p����/>�����L�Չ�=8���5B��7d��5~��/��6� �B>�[X>x?��_6��$�?}�Y>u�?>Jy�?�Eu?_ >��	�վEO���e��aS�A̸= �>�<��e;�O`���M��lҾ;=�>!E�>���>��>�A�z�w�?jW>^��[W����>u�D�^.�����!K�����U���m���`=�C?O�����N�3X�?��y?ڑt?tY�>o�l=d[��%ئ><7��D��=�� �����:b=[�4?�t&?8�?�U�',�P̾���Jַ>�9I��O�����0����1Ϸ��|�>A骾�о=3�d��R���I�B��r��ۺ>6�O?J�?`Mb��V���QO�d����r?x{g?�,�>fL?20?�Q��-X�[t��uո=8�n?���?6�?
>��=���>�?yj�?UW�??�x?��0����>��p=x�[>L�����=�H0>�b>��=�J?z�?V?������n��q��v�K�	˶<�4=��>�ف>��r>�>U�K=a+=*�N>��>5��>2&f>_�>�>�����	K�R{O?g#�>P��=�m?���>E!�kR@=�,>P�=]�+{��ߑ,�bZx��KH�i�ʽ*>��o>d ?i�׿{?e��>����$C?`����t�4�j>�C�>GV���>P�>�f�>y݊>8�>��b>�W:>qn�>4�Ҿ��>!��W!�QC�vR�3iѾ*�z>�����S&�;�����ΊI��L���@���i��:��ZL=�y%�<�;�?�t��k�k�0�)������z?��>1�5?a�;و��G>�r�>U��>A5��y���dэ��z���?p��?];c>e�>C�W?��?��1�o3��uZ���u��&A��e��`��ߍ�y���3�
�X����_?y�x?yA?'�<"5z>���?f�%�7֏��%�>F/�K&;�K.<=�+�>� ����`�īӾv�þ`;��GF>)�o?�$�?�U?�VV�8e<���=TZK?�G?k��?p7L?xX?`/�;�#?�>{?���>*E?��I?�?p�>���>x��=��=5�NŎ��fڽ�@q�I���=<Ϗ=�3�=u�<7f�=���=���d�R�C���^�<���=�8/="�f=�>j��>:q]?t��>}P�>Fj7?��P�8�����.?�z;=���:銾팢�����>d�j?�?|9Z?u�c>x�A�m8C��>�I�>U�%>�k[>F_�>���]TF��
�=�>�->��=ٝN�ͣ��{�	��-��`��<��>9�>9�>U�{�;<�c���֖�F{]��$�~�½C=�u�=��GT���i�ne>��*?�~ ?w�0=sݾ�ü$�p���>Lhc?�s�?�7@?�b������n8��E��69����>�� >YM�{���G����:����=B|�>8ۺ�������e>��
�H�߾Wl�GI���龋�_=�n���W= �
�M!Ѿt�}�Rt�=^> %��l�Р��ᶪ��"I?��=���3�Q��b���>Ř>��>2����v�i�@�ⰾ�9_=�&�>�.3>$)�����LE��w��e�>tH@?p�f?㼃?x}�60r��AB���nu��=�b(?���>��?[��>����∽��p�l\P�#72����>_?���5H��c������I,���J>�� ?M�d>�� ?�uG?��?��f?�)?&�?e~>=�C��";��?v�~?�y�sA�-$H��r4���9�A��>��O?k��Ci>���>�?H.'?�5?�?��;>GQ�#�Q�6�>]f�>r�v�x����lk>�_/?���>og?�?����=�τ�ˡ���
>h��>�v1?��>n��>T��>0��>8����n>&# ?��?�?AY�?�=���\�>C�c>���>�(/<�[�>��>��?<0? ��?��a?��>Q�<�:O���o)r��0�<�W>>}=x۩=�L���[j�"�d�P�Ͻ-ཾ;|�㵈�4X��WJ=|�=���<$��>��u>�n����.>G�þ8a���m>>����3���׈��8����=k��>��?���>w%�*��=0��>o��>����'?v�?u?���:rnb��۾̰M�$l�>�A?���=|m�ȓ��t��^=V�m?7�]?|�[�W�����b?�]?� �B�<���þ�c���e�O?#�
?�nG�Y�>��~?�r?���>�<f�*n����Q2b���j��Ķ=چ�>�]�~�d��V�>G�7?�#�>˰b>c�=�G۾��w�.s���?��?���?=��?1*>?�n�C)�/����D���_?�e�>:ڧ���#?|����Cо�����򍾈��A��\9���������j�#�}ق���ӽT��=\�?A�r?�q?y�_?�G��Pd��Z_����x�U����U�C�D���C��C�	�n�t���\��)6����J=�D�L�F�l�?��5? CG�'s?��d�����?:��&DZ>�c���R ��>	�.<��+=bNc=$:�N.��r��^?Z1�>=��>k�>?�=`��@���E���9����i��=��>g�>���>����fe��'�"H�������[Xv>�rc?��K?��n?�1��|����!�d�,������C>�[>^�>K�U��=��&��T>��r�E��Bl��G�	��s~=l�2?(T�>w��>"F�?V�?*I	������x�l1��?�<G�>�<i?ɍ�>��>��Ͻ�� ����>b�l?�}�>{�>O����U!���{�FpʽM�>�ܭ>���>V�o>�>,��\�`��x~���9�f�=h�h?�v����`��>R?�$x:�CG<�S�>$�w�U�!�.��Л'�D�>��?5�=�p;>Zž���{� i���I)?M@?@ɒ���*�)a~>` "?��>�>�,�?.�>�Xþ�$�
�?�^?BJ?�IA?�F�>�K=ﱽ�8Ƚ��&� �,=؆�>�Z>��m=Ƿ�=���z\��q��DE=)�=JCм&�����<Po���L<���<��3>��տ�U�;�
5�m@��eݾ$�ʾ���]t����UC�0��")����_/�
;A��n���>����T�h��?iR�?N1���䨾�d��_j~�*e��M?�+�q�V�P��R������r��*�����#�j%^���~��zj���'?+菾ަǿ4�����۾R?�� ?uy?�����"�o8��>t��<*؎����N]���4Ͽ㛾B%^?�t�>j��΍��A�>��>�T>�[t>ӻ��h�<`G?�,?\�>�ws�4ʿ����jJ�<�M�?j
@�hA?Ɵ(��0�VP=Ki�>�|	?f�?>��.���WR��%3�>I�?���?�^E=«W��Z �n|e?T�;GG��1ӻ��=�#�=+=���A�J>��>����}A�|M�ڽ4>܅>7�$�`�fA_�>�<�p[>J2ٽ��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=����п�`��J���½�15=�YH�f:J�P����f����Ⱦ��ɾ���<�7�=��>���>�V>��>y�X?cY?���>��!>d��l]��쾨��=�����;ھ�<rJ�����+"ʾ�E��/����׃������.>Z�^�����e`?�@J���_��pV?�>ps��]�K��Ԅ���Ҿ=Z�+� =JY�<�����)A�/:f���?!E?�Q���t����Խ��>��?�ܘ��_�s��S�>a����QA�|R�>2�>����-���>�C ?§?�WԾr<��lU	>�V���=�?���>��a=�|>[�"?~�ּz�I6>�<�s�>��?pG_>�_��p��ث"?�Z?8�h�9&̾�6�=s��P�h�B&>Z!�>�9����	=��>$緼.(H�݋��(��!c���G?���>�F��//���O�����}-��s?M�?($b>��/?�N?X=ӽF�꾯F;�����ˉ$=m�m?�r?q>KXݽx�������t�?�	�?5ݭ>�8�J���4�d�}*?	��?��?���l�i��o����ؾq�M?��v?s^�xs�����N�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?g�;<��U��=�;?l\�> �O��>ƾ�z������1�q=�"�>���ev����R,�f�8?ݠ�?���>������Y5>]�����?���?�q��7�#=$\���r��𾡳�=��^>$�B;B��=K頾;G�]�׾�������w�=>�m>
+@B)�z~�>��ν���4�����n'���%Z���,?���>F��X�����q�	�p���a��K�gQ��j[�>�>�׽{D����{��;��;����>��u��O�>l�h�hs��〣�	��.g�>�G�>RW�>�fý�Cž?�?}���̿����k��U?d�?;�?Y�?�V�����	D�D\�5�>?�,l?�\?u�ٻS�G��C���j?�]��BU`�֎4��GE��U>�"3?�B�>#�-�d�|=>���>�h>#/�ύĿVٶ�����3��?s��?o���>[��?�s+?�i�8���\����*�h�+��<A?2>:����!��.=�cҒ�w�
?L}0?�|�b/�]�_? �a�P�p���-��ƽ�ۡ>��0��e\��L��)���Xe�
���@y����?M^�?f�?ڵ�� #�^6%?"�>Z����8Ǿ&�<���>�(�>"*N>H_���u>����:��h	>���?�~�?Qj?��������U>�}?Pò>���?I;�=܎�>���=�빾����>���=x8���?��D?b�>�C�=3��$.�Q>��D��l
�Cu<���>�}b?O?�;V>��L����#�r�Q�c)����NrY��︼�ɘ��%>C�S>>6>��v�h����?Lp�9�ؿ j��p'��54?/��>�?����t����;_?Qz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>;�>�I�>A�Խ����\�����7>1�B?Z��D��t�o�y�>���?
�@�ծ?ji��	?���P��aa~�.���7����=�7?�0���z>���>g�=�nv�߻��5�s�ѹ�>�B�?�{�?���>"�l?��o�L�B���1=M�>ʜk?�s?38o�r��B>l�?������L��f?�
@{u@M�^?#y;��ିِ���l���=g5�<�\A>�����b�>\�!�bu'�b�<e�P>��q>�>]SP>��^>�	>�����3&�C��I����zL��"�|)����N)�p����'�~6��������+=ء��%�<�'g���M��	>=�D�=�JM?""V?�p?��?JXh���>�2���I=aJ�F�=�e�>(D7?dV?N�1?X�=���P\��{�j��k`�����>\�Q>n8�>�M�>l��>a�==J>>�� >��w>	#�=�_»!��=?sP>[��>���> -�>��>Lw�>޲�㷧��=��e)2��x���?�~~�])�������Ϟ=���e�b��>Y?ߨu��ѿ*F��f�#?wWڽ0�̾D�U��奻��>��C?��=�ﾴx�A�
>'����~#�b�'=D�?����^t�՞�����>�Ӏ>X��>c�@�F)P�,�m�[F��t�2i?S,��U��ء���a߾^���1�O�my�>)3�>�j
�ZƤ��ݏ������<�<?��>�E�>�����t��h �Aa�;%�>#� >���>
_�=d� >�6��5�=�Q�>^ >6�?��>>N߯=u��>�=��a}h�"�>��)>V�*>��??��#?Am-���Ҽ�+h���?�W�P>2�>Hd�>�Y�=>8���=��>t�p> �$��Sl�z."�v�J�0��>.#�!`D�����=���E��=Ղ�=��˽��o��`6��~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿe�>��*]�������u�\c!=`i�>�7H?%����O��J>�r
?��?�b򾯚��?�ȿ�bv���>���?X�?��m��A���@�X�>��?�iY?p~i>�g۾1�Z�;��>S�@?�R?d�>�5�*Q'��?!�?.��?[�S>���?i4w?2R�>Ȅ�U2�a�����7�=���<y	�>W�>�����5��锿Af��L4l�:��/Xb>}�=|_�>����ZǾې�=�{���ղ�J���LN�>�W�>%�C>�=�>�?�P�>��>w�t=�/���2������N�K?��?W���3n�k@�<-v�=��^��1?�B4?j�]�^�Ͼ�֨>[�\?���?N�Z?mu�>���A���翿����v��<d�K>,�>Jl�>{A���K> �Ծ�8D�e��>˗> ����,ھ�������9�>e!?&��>zή=�R ?�#?�yg>/��>BD�ns���F�e��>��>>�?}�}?@�?������2����Ce��J�Z���P>�fx?3�?#��>�����a��>�+G�j���p�?\�f?45�Ի?sy�?I�??�eA?p|d>yD�Klؾ놣�
҂>��!?Ϣ�H\B���&����#?f?d��>�)���뽃0 �$T�<}���?7tZ?4�(?-��+cb���ž���<D��~���<�@��7>�Y>���rl�=Ճ>���=�/o�&�2��{<*<�=)��>�6�=�39�Ϧ��.=,?\�G��ۃ�n�=��r�7xD���>JL>����^?�l=���{�����x��#	U��?���?Pk�?���9�h��$=?�?U	?^"�>�J���}޾4���Pw�8~x��w�c�>���>ۣl���A���ڙ���F��g�Ž	s��\~�>�e�>q!?��>���=c�>G����4�uо���Pkk�!�[�S�F���)�|������ɻ�����K@_��ŀ>�&����F>�*?�g%>��a>�R?���=�}>�͉>�>�>���>R,�>[E�>��h>�u	:V�B� KR?�����'�b�辍����1B?\pd?90�>�i�'���%���?���?Hr�?�9v>�~h�[++��n?x=�>[��yp
?Vf:=���z%�<�V����� :��������>�=׽� :��M��hf�6i
?�/?���̾N׽+f��>�~=䐄?;w'?_o(�,R�Qp�NIV��DR�c��~7j�7����6%�˭o��Ɏ�D�������(�%=߷*?'�?z��(��ừ��lk��B>��h>IR�>���>�b�>ЍA>���)�1��1^�j'��������>v�{?��>��8?��D?�W?�fN?�!�>��>�8Ǿi�>�i�=�¬>^��><�C?wA?�4<?:5?(d?;�_>=5���������0�?E5?>�"?��?�8? ��XԼ��ǖ�NP�a:z�4��bκ:X�<����)����=��?>��?x>O�?���t�>{�8?��>BB?�������N���F'?��*?�Ƌ��XҾ�q�+�����?� �?�j�s�8<�>�YR>i������c�[>�+����S=�h=��=���l�@>�/����<�.6j=�D���}\�+�>�^?v��>j��>���p��]<���=e�\>�R>��>sHؾ����X���6�f�Y�w>O�?OY�?*�k=���=���=����t���7����_��<�?'"?c�R?�&�??�>?��#?�>[��|����� ٞ�P�?��<?��>"k	��⾴���-Lp��m6?���>;��5�]��}���;��,_��#)>d�p�x����@̿�Kf�@�>�Z��'(����?Vƨ?��]��X�1�������D�7���N?���>�+>t��>�X��.���`i�y��=޿�>���?rb�>��M?m�?�Gi?0J�>�J(�~V��អ���R>���>��S?��d?T��?,�?�"�>�~>~���fA޾�Ծ%xؽ>^���k�6B��%��>hB�>�� ?O/�>�݈=�6Z��j�.2\����<���>�(?���>��>赃>ƭ���V@?D�>��ܾ:��N���P��3uؽ+x?��?j� ?CW �O{
�r|R��.�df�>���?���?��&?�|X��5>�b3��оcy���c�>���>vê><A�=EW=�t�=\ �>��>4Z�E����7���!<��?hO?4�(>D~ƿ�r��q�o$���(<�����g�����]����=%ٗ��������\�1���dz�������H��Яw� ��>��=���=M�=���<�ʼ�7�<��S=M
�<k�=z�R���C<6����P3����LOt<b�V=R�û;�ž�z?[�K?�,?>M>?��g>{�)>K�Z��X�>���>�?�&P>i)u�$��d�M�Cn��)Ŕ��a־�,Ҿ�W�6â��>m"9��r>�BK>��=΋Q<p)�=�7�=&Ư=R��<?A=h��=0��=I�='l>C�
>��>�6w?X�������4Q��Z罥�:?�8�>j{�=��ƾp@?}�>>�2������yb��-?���?�T�?=�?Ati��d�>M���㎽�q�=N����=2>s��=w�2�T��>��J>���K��D����4�?��@��??�ዿТϿ6a/>��=��$>��A��;�R�b�v�X�l���Ƀ'?v�J�A���09>��x>y���a便�O>M�G>忸<�y��d�v�ǡZ=pX�;hO�=2.>ɫ�>���=�
.>�`�zh>o^F=�G�=y�=�g5���=�!����<Cj=TO8>	�W>F��>�i?�*?�wV?<��>�|��оok��k�>�>�"�>��;���=��>~p6?۪0?��>?SL�>��ʼ���>�߻>��8�s�`��ݾ�b��	=�7t?;��?μ�>d@��
�a�UN#��_8��#0�_�>�m2?o�'?(�>����쿊�`2-�GT��fF���ƺо
���NC���}�$�����:�>�5�>�m�>G�>>4��>K��>ʹ>� ==<��;�'�s�8=l�*�a�=ͣ���.��,F>D=�9�<��(��s�cU�=��=7�=��=��=���><�>�>�>B�=�����'.>�]����L����=Ms��=�A�Ad�7Q~���.�1)6�͆B>b�W>u���4����?�kZ>��?>���?�$u?��>A!��־W-��L�c�׿R��=�)	>.<��;�;L`�f�M�7zҾ&��>C��>Q��>�ޒ>j��r�a��R>���7u��R��>�Y�M+X��s���u�<���\ݶ�������[�Z�U?Ö����1��x?3u�?�?�i#?s}Խ(t��">,!�����=zpԾ��z�`�A��<@?�a,?�x?��1�z�_�Sʾ����i�>��N�eM���z�1����
,�����>~'��KҾzv5�G�����h9B�|�m�(�>jM?�q�?I�^�J3��P�����ی�*�?��f?��>B4?p?�!��p -���.�=��m?�W�?74�?�y>�@>>���?��>=/?F��?��?�1y?�~��k�>�6>C�>��㼍bb>�>U�>��o=��'?aV*?Lu�>�z�������9���\��!l=��/>w��>ٓS>9ٚ=ȱ���qv=�R�=\9�>��l>-%>_�}>C?�>Ѻ>�i��1��G?��>�<h>�g;?�̶>�<��N�Z#~><� >��@�x�1�Z=K���<5 �=7=��-=�k�>��ǿ�?-�>�;�JZ<?|���ӑ��N(>G%
>���>Z�>K5�>�Ҝ>��>���>�zN>T�>v��>�zɾ�&7>��k$�=8��X��߾3+�>�ۄ��w�7o�q��5j��@�����H"f�A�x�rz1����<���?_��r��-�NE	��v?���>�4?:Ju�t���x�>��>b9�>����H8���4��-پ!j�?�f�?b>-k�>��V?my?n�.��6���Z��`t��@���c�9�`�����΁��a
��Q��r^?�$x?��@?��v<��|>8��?��&��Ԑ����>;~/�܎:��HD=��>�°��qd��:Ծ'ƾ����:B>8�n?��?��?AP�U��=c)�<Nr=?O�S?�L�?M?u3S?՘h���&?l�>�9)?*^?K/?2	3?,d?3>��>a�>�E�T��l|�7��#瀽	䟽8�<�%=�Z$<���<�g�=k�=�o)��/��w��g�O��κ=�4�=����1y<`æ>��]? b�>�̆>��7?���Q8�X뮾�/?;=�g��� ��*�����  >�j?q��?�gZ?Fd>��A�x�B���>�8�>u&&>��[>�p�><��SuE��
�=T>�i>q��=8M�{ځ�e�	��X��L*�<?>�5�>q~>O����e>�=����z���U>�F����'fS���H��/��`s����>�jK?sg?�V�=K��f�����f���&?f�<?�eL?���?$d�=��۾��;��K�/��9p�>/2�<�I��,��\����<�\�::�A~>Q̟����Fme>n�	��F޾Yl��0I���C=G=9��rsd=��x�վ�`z����=aZ>5��iB �L&���%��TdK?�Տ=�G��l�d�%`���r>6��>� �>N����w�`�?��}��z��=q/�>��A>rj
���꾻H�mQ��G�>^�8?6�\?��r? �3��hJ��J����R����0g��?[#�>k��>�Ln>=��=k̾�$��~c���-�=�>U�?2�~]��;Q��}�n�8�)f�>ˎ?5�]>���>��1?��?�{q?@�-?��?Vx�>��B��%P ?"}�?�Pѻ�r1�'�.1�i�H����>#�4?r�'���E>���>��?0b"?�[R?��?l�=ŏ
�a�5��>��>7t��W���=`�+?.g�>7�e?Q߇?�]>��3�\����#��*>�[>v�>?�?��?�%�>W�>�B��d"�>j�?�0�?J�?h�?�@b��.?�b�>M�	?�Bf=��>�?W|?�25?2|?[A?�>�����d�ؽ�H�;��>���=o��=��=A��nr�p�C��4/=H�=�Y�Vt�<��>��������=;�G]�>�s>����0>��ľ�L���@>�_��;J��������:�B �=t��>��?欕>�^#�l��=���>+M�>?��04(?��?�?��";`�b���ھ��K���>�B?���=��l�}�����u�/h=��m?��^?՜W��'���yb?�^?���A�<��/¾��a����1]O?%?lTG�Ҽ�>fV~?�q?e�>2�b���m�:���ϻb��k��Լ=��>[^��'e����>�6?�)�>Y�f>b+�=um۾��w��7��r ?#�?��?�,�?�D(>gWo���߿;��Td��<&`?;j�>�b��>)?���;p^ھQ���0X���+׾�|��h��1���(Ů������rս:��=m?��p?�Br?zy_?��$�`�j�]����jYW� Q�a���tA���A�/>�#/l���	��������G�d=�B��Q�/@�?z�@?�7���j?
�Z��|����u�>4�i�_�D~�0ᓽ�T�D�x=�9s�]�%�Z=�3#?lr�>��>�:?6b�^�2�ă4��;��q�� >�ۥ>��>�W�>��J=�];��D��;Ͼ����Ju����>�ud?�T?��p?�� <�Ѝ���4�
������o�>+%>	;�>s��r?)���!��);��u�K��3?���w��z=�I#?�>O+�>d��?6�?e���*���\*���/�e̲=bջ>|	o?��>��>��j� �q
�> Vl?���>���>C����2 ��U{��˽�8�>�ƫ>��>\/o>K-��\�ܺ���X��#�8��"�=
�h?t!����c��-�>R�Q?�;5��<ݭ�>�͂��"��|+���>�J?!�=�y9>�žQ��C�|��K��W�(?Ĭ?�����8+�k�}>�0 ?X�>��>���?�G�>��ľ�<�?rk\?�`I?�l@?/G�>�O=���+Lǽ�"(��R)=�"�>��W>E�}=�9�={��OZ���%���/=XJ�=�JY�� ��� �;'�ؼd�?<�q=��7> @ӿ@!G�ݽ�������羋�� ~Ѿ���8z�����<阷�����%���6ֽ]�üAdj�����<8���u���r�?���?V��P۾�V��9	��������>��Ӊ=��l�P�_��kc��|;H�}�'�lR�Y�j�)n��A?\$/��¿R��G����.?^!'?�@}?��5�8��E�-�߼4���
��=��;	����1Կʾ�rD?s��>�]�y:�<�O�>�B�>tr>��r> �����=�2#?��>��?���@�0_ο�R�<���?Ш@P2A?�[(��;�ƤC=~{�>��	?��?>�8+�U���������>�}�?Xh�?G!0=�)W�q��Kf?[�
<��G��[���l�=s2�=:�=S
�hL>��>^��>���ܽ��3>L'�>ŏ$�R��&_���<��[>9^ս����ф?�]\��f���/��X��2�>3�T?l�>a"�=h�,?U?H�:zϿ��\��a?��?��?=�(?Nݿ�y��>T�ܾ�M?E6?��>A&���t����=S]Ἱr��2f�ZAV�8�=���>>�>�@,�,��{�O�����?�=oP�6�˿1���1��<^�<�������E��)弹���W	���$��3�=C*�=Q{j>�w>W�J>�<e>��S?�x?P��>Ok�=Y��D������&�r�u��L��U��C�&�������ݾKξڐ��s3����c����(��U2>�-0�刿����s�)�\��?�ď=L�8�4�����gb���Ox�O6>s͔�}X��ݱK��m|��פ?A�G?����S7�������H=l��?����������:>>6=����_�>�>�OȽ4�
��
@��A?}�6?��߾����ȗ�>��/���	��#?�
?BU[����>R "?)t�/ϲ����>�6a=��:>�>?~��>X�������9?��S?8vB�1�BB�>4�ʾ�_A����;�}�>����0b���>x��<������	�j􌽤�L?>y8�F
%�B����B��c'�DQq?�h?7�>?�O?LmH?G��=��󾀺<�V�^��=�3g?@m?#v>ۄǽdӾ]����#?I�`?HY>2�M�|�Ӿ�B4����[^#?^��?-�
?�v�^�s����R�Ӿ��>?Uv?�a]�|�������0`��ק>���>*��>D:����>��>?8��=���K���3�hm�?��@�,�?$;��I�=p?*��>�7P��4ľsi��/����}=#�>x^����w����[�!��=7?�?��>�������RL6>���<�?W�?����J=���+��j�վ�*���f>�L�<� �Q:��] T��z���z� ���>/�m> @�.ڽ��>����-�,�ڿ�6~��v���mT���?{��>��=!/��!T��u��
A��T���̾r��>�1>�A�X�ʾ��w��@��Ū��|?#���Zٙ>�ER��+��nߍ�ب���a�>�'�>{m�>	1��r�X��?!�޾��Ϳ+�����M	_?[��?���?�?��་
/�S���6p��a?~Y?&d?,e>v1��5��e�j?�奄!	`��X4�D�D��iS>�;3?���>�.�3C~=�{>w`�>�t>5k/�f�Ŀ�������Ц?=��?���m�>\��?ʧ+?u�\[�������
+��^��i%A?�.2>�Ϳ��"�jH=�)钾:\
?�Y0?����V�_?��a�b�p���-�Z�ƽ�ۡ>O�0��d\��N��q��}Xe����@y����?#^�?i�?[��� #�6%?�>����8Ǿ�<Ӏ�>�(�>)N>�G_��u>6�-�:��g	>���?�~�?Qj?�������iU>��}?���>��?�8�=e9�>O+�=nf��z[1��#>4��=z�B�5�?G~M?:�>ޛ�=O68��/��9F���Q������C�ׂ�>�b?�mL?�Db>���PL1��!���ν��0��]�#�?���+� �ܽΤ4>D=>'>r�F��Ӿ��?Mp�9�ؿ j��!p'��54?.��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>@�Խ����\�����7>1�B?Y��D��u�o�y�>���?
�@�ծ?ji�؈?_��c���p��o��O7�"C�=�8?J��}�|>H`�>˻=�Eu��	��g�q��i�>l�?�G�?Z!�>�l?�n�`=C�#7.='��>�l?<&?��:MH��;>tw	?������P���c?��
@�C@�Z_?�<����ҿf���=���5��#�>)S=G+P>���ϲc=���<r�<�{�c >�_�>^�k> ��>u�a>�	X>q/>��!�"��&��&����<��:�k@���l�pu��i����%�����3¾��k��Ľ`�-��V7��!�/ �HZ�=KT?amT?}�p?�7�>T��9�>���5y=�<��y�=�g�>�w7?�O?�J)?��=G䚾j�b�����5��A��ǿ>��F>t�>��>cO�>e�|<k�M>QT4>�h{>�Y�=4&=_�;��D=F�P>+`�>n8�>���>4w�>_�>[(������"v*�{ܼ�	A�<���?����R]�5ܧ��ٝ�K㛾��Q>yQ\?Ib�>0���~ѿe��2�M?~ѣ����녾��<>�+?��h?a�>��N��uvD=��R���� =��\�롐�#�P�M�>Q�?���>�ʕ>gB��`E�O\���L���N=�+^?)B��X\>jd��]P^�哾��=Uǽ>�X>L�J�����r�� ��kb�=�*F?��>���==�����WD��]6A>N��>�v��*�=d2�>�=N��8O����=����ca>	?�b,>^��=�,�>����Q�M��d�>}C>�{,>??P�$?}��\���GU���d,�եu>��>'��>4�>R�J�ի=�8�>�b>�����|�b���A���U>��s��b��v�ю~=&����=jG�=�� �(�@�7'=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾNh�>Fx��Z�������u�Ҷ#=2��>�8H?�V��7�O�p>��v
?�?�^�ש����ȿ&|v����>S�?���?b�m��A���@����>4��?�gY?uoi>�g۾M`Z����>ݻ@?�R?�>�9�~�'���? ߶?ٯ�?�:e>�׏?��z?x �>����KD��귿���FM�=��4��	�>��P>Z��7�'�H��aɆ�s�j�%k$� 2]>��<;��>'	�A�쾜I">u����˾��V�7ȯ>r�>�3I>y�>f?U��>�G�>{��<w��������ž��K?5��?���4n�q:�<aw�=]�_��?a4?��(���оOԧ>k�\?��?5�Z?�Ȕ>Kk��@��3���}O�����<|[M>�y�>`��>���@]K>�dվlD�w��>ϊ�>�4��Z�پ%m��Ӡ�ݽ�>��!?��>��=c� ?��#?~k>�L�>�VE��?��NF�!��>���>?��~?4�?Uڹ��3�$��á��~[��OM>��x?&2?	��>������)�>�[P��2���}�?
vg?�㽚�?$�?�??<�A?J�f>��#�׾	�����>�"?i��C�'o'�� ���
?\�?W��>�7���:��G������Ʋ���?��Y?��(?��5_�i�ƾ�T�<��D�p ;���;ۍm�(~>2P	>�D��x�=�#1>��p=U(��ܠ+�z��<�I�=X�>�ҩ=�<<���|��?,?NSD��Ǆ��w�=2s��C�p�~>J�N>F����^?6t=���{�w׬��b��0�T�?�?w�?�#�?���6h�I!=?S��?��?`D�>�*��h߾�.���u���t�Q�k >V�>��J�^L����M����.���ý呹�.��>��>e!?��>qɴ=���>;ȃ���ؾ6j��}쾩Nc��F�i(�Sd+���K����]q��¨=X#ѾR���^2>L>�%�>R?tf>ӳ�=��>}ʷ<:g>�F8>ܶ>9�>ia>���>��>�wS<r�;�JR?q����'����Ʈ��62B?�nd?�0�>�i�鉅�����?���?�q�?�>v>h~h��++��o?A�>����p
?pT:=s%�9q�<�V�����3��r�ƨ�>�1׽�:�yM��mf��j
?�.?/7���̾�?׽D����x=���?��#?!�#���M�W�j�S�T��.V���&��j�iU��f"(�%0q�J���t���񀿶�&�R�<��+?b�?A@��� �Mu����h�3WB�5,w>�>�>L#�>���>�>`��|/��MX��$��H�����>v�|? h�>��<?ȹH?�'Q?~I?���>5�>z�ƾ;;?,yd=���>�,�>�mB?�.:?m�0?��>!M"?��>帮��������fr?z�?yY?��?NH?��b�0�"�V�9��D�s�\�}�ƽ�J�=�#�<�k��B�L�����TS>*O	?zq�=~lO�0h���u>�?W�q==��>"󴽙����m�T�!?�iS?���=9���YK��ľ�8?��?�A��=�G>� >�|�=5- ��_>_M���=�q�QW�=
�ͼA�=�I����=\���QɽH�<�7H<#S�>�?x7�>�Ĉ>����� ������=\Y>�cS>b�>w>پ�s��$��W�g���y>Xa�?}h�?Y�f=���=�6�=�
���������E�����<��?~d#?�FT?�z�?��=?
�#?P�>V���.��BB��@O����?��K?��>s� ���¾z����D��l'?���>"	��!�����!��)�}��x�ƹ���'������s/�mi�>���c��I�?[�?vCսo��\׾wN��LG˾xU?B��>�Ҩ>���>�=a�m���=�A�2>>R�?A�d?K�>�-P?Gj�?/d?�>[�K�W����
��}�=�Y>,�e?iqr?�W�?���? ��>B*�=�L��}������'���-�.�n��=F�I�>�>��?���>�j�=�g2���x��
n�6;>-��>�>?�F�>O�>���>�AD�'�:?f��>@W侠�"������)�׽��u?�z�?�R+?�5�<���c8�~s��*�>��?�+�?�A*?�'`��">)(G����K�c����>�o�>l�>��=o�=���=ϱ�>���>��H�q����*����;��?A�[?{3>{����El��L�����>-o=뱌��U8�8���V����;=����C���˾�p�����x��ȝ���Δ�w������>
g�=���=P̧�i|�<���R�s=��<X�m=�xp��?���a�qȃ�&��J(���-V��W=�Y�<�˾J�}?M;I?��+?�C?{�y>vM>ͼ3�#��>�Â��7?�U>&3Q�w���ˌ;������#����ؾ9_׾�c�՟��@>B�H�\�>�N3>�;�=��<��=�fs= ��=;�L�Ȯ=�i�=":�=��=��=�>�T>.�l?�ab��z����W�Bᚾ�D?]ig>$�>��ξN�-?��K>�b��1��� �ڣ[?���?W�?s��>�ܭ���>�wW��9���=H����&>8!W�W� !�>���>E3<��H������Q�?'!�?1�?�Җ�?a����m>�1>�Ղ=.RZ�<?C�X���ki�������
A?��P�T�ӾA[�>�?Jn�B3��></��>�x�>&ۍ�`�����>����[ �G>�k>E�>h
>鲈�pA�=s�����%>v�=^4ܽs�۽����D>&�=`�q>� M>���>��?�)?�@Q?��>��l�Bm˾= ���f>���=7��>��=u2>a2�>�\.?d??�D?X4�>�� =�%�>a��>eX7��J|����#
��DF=��? ݋?D��>+�9`�������2��ᏽR
?�!?e?�C�>)��5���#�����-���}��VS>�
!��叾����؎὇��q"��q�>�i�>z<�>�s�>�D>}��=)P�>��~�G�=�>�G�=(>���c?�=�^g�jU>	����-1=2`<�Ž&2ǽrF�H�M=�C�=l��<���=K��>�@>O/�>_G�=>���,>k!����J�"��=}���4�@��uc��}�(6-�o}8�jvA>��\>O�z�%鑿�] ?�=c>@�C>��?�u?�">�L�ܴ׾tX��E�j��O�r�=h�>?��Z;�l_�{�O�n�Ѿ�9�>O��>2]�>X߂>0��Pl�V��=�����O����>�F}��~#�Mj��Ww��!������e����Y�7PL?������F=d�x?0K?��6?1f�>X�e�����>7@�����=0˾��n,�=N�P?uh"?�y"?��ݾ �p�F�˾}渽�=�>`M���O�륕���0�t���:���>���Jо��2�k:��N��3uA�-$p�Nٹ>�+N?$ͮ?�6_�轁�C�O�<��F9����?xh?��> ?�?֤����뾥��Un�=�n? p�?�<�?7>��=�휽J�?�?m�?S�?b^�?����?�Ѕ>A�>D�ٽ�?>u2�>?�>"=�?g� ?X[
?.��k�g�[پ����M�=���=�;�>��>���>
����B7=~U�=$ς>�֥>eÑ>�0>;2R>H�Y>���&F��'(?�a�>�9>�0?�R�>Ġ��U�=7d��;t=��)��5�;��[�]�觸��韼Wx�=��=��>'\���Ǔ?y��>�k:�7j=?�Ѿ�p��w*>ͧ\>d�S ?�U+>
��>��q> ��>��>I�.>E�e>�+Ӿ��>B���q!��C��~R���Ѿ*�z>r���"�%�������Z�I��u���V���i����g!=���<9C�?������k�/�)�>v��q?f�>�"6?�g��]3��E�>q��>w��>���mx������T�/�?0��?�Ma>V�>�,V?ק?��-�Ҁ4�$�Y�Avs�L�@��/c��P`����������
������^?�-w?��??��[<p&>�;�?vX(�,r��� �>CR/�o�<��a=���>򇫾A�`�2Aؾ����Mr�"�H>�(n?���?ny?�xH�RM��� >�.U?G7J?�?x^8?�h[?8ꏾ=�6?rm�>fA$?*I�>�C?hxX?}?�g#>�C>���=��k<��Vn��O�6怽-&�=��=�v>�H<�� =�����L�����^����U�0�=��=�.D;��=��>Go]?���>���>�X7?����8�/j���.?(�8=�!���I��:٠�|
򾮭>>[j?㔫?Q[?Qg>#~A��D� �>�"�>�y%>��]>�Y�>����GE��[�=��>�>�9�=�Q��́�+�	�R2�����<�� >��>l�o>�������=�����Y���`�=�Z��SľYt׽�Y�^��F�:�.��>(�3?�8!?���>�2�ty��c|�2o�>�J?]�o?��?���;����t�MY�����7�>��>�:��*��C钿Jl,���g=i��>Qr��BꞾWc>���7�྽zj�H�G�Q1�A8r=��EKR=�.��@о�.{�)��=˧
>r��y��o��r��O�I?��w=�/���cW�j���(>W�>MU�>if�67^��D��ұ�Vo�=ZU�>��9>QB��S��8J���\-�>�-?��f?F/�?�
�����4UG���+��^��Qo!>��?��>�? ��>��5�m�l�ع.�gyF���U����>	?�1�,S]��kýf��S�o��>T�> �[>�o
?]�P?��>;��?�->?}�?��>˓ս|Q���#?O�?�#s=��㽀zQ��]7���G����>��*?j�F�~w�>��?�?#?rLP?˃?Td>Ol���>��n�>���>�W��&��t�\>�OJ?�R�>�Y?}��?�6>U�3��Ş�Χ���F�=h>�1?j�#?��?Qq�>[G�>I ��Ӛ>��*?[�w?�@�?�ل?��@�d��>E>|�
?�ƽ��(=E=?�-?]4(?��l?gGJ?L� ?�5��iQ���+�m<���7�=��=W�ռ�F>�u<��"��J[�Ό@������k:=G =�3/���"���S�>��s>*��Y�0>J�ľ	j���}@>���#E���䊾�g:��۸=�>��?��>��#��~�= ϼ>n[�>����-(?E�?*�?�;w{b�u�ھf�K�&�>DB?H-�=�l��j����u�˟h=��m?��^?�X�- ����b?��]?�I�=�Hľ��b����|�O?e�
?'�G����>��~?�q?���>�2f��$n����p:b��%k�f��=�w�>�\�W�d�*c�>+�7?�>�>�c>"�=Wn۾V�w�ia���?F��?��?���?�F*>��n�a1�l)������0�^?n��>:8���#?&����о��������]*��A��E���Ŕ�����PQ%�B섾Nٽ���=�#?#r?Z�q?��_?���|c�;^�0D����V����s����D��C���C��bn�I���z��<���*�>=?4-�ʾa���?�z7?,�;i9?"^��s���(`����=��X���ؽ�&�������c��+N�<������B�g\K��$?�֨>q��>�$<?p�k��<��1E��N�9����S>5�/>,��>~?� c�լT��ؕ���پ�2��D��=v>W�c?O�K?��n?p���D1�b����+"��M<�ꮥ��WG>��	>e�>�L�����&�R=��r�+-��.��L����= �2?���>e��>�ۘ?y�?y��ʶ���u��o1���<��>�wi?%�>��>_	н1��J��>��l?��>��>�����Z!��{���ʽ]�>�̭>p��>l�o>�,��\�e��邎�M9���=2�h?ق��<�`�Pم>�R?��:s$I<�n�>Βv�+�!�H��O�'�U�>u?ؽ�=�;>�už�&���{��0���$)?�G?X��:�*��L~>"?d��>n?�>R&�?ܫ�>A�þd$;�q�?��^?�I?E_A?��>@�=����ȽLI&���-=Ok�>�Z>l+k={*�=?��1�[��R�#�A=Ɓ�=�μn����<�f���A<*��<�3>^޿�U�����a'�����C����Y��<?͞�6�\�)Gξ���F4���7�VI=�P����k�V����׽���?-( @�ʾ߅��e��bu���1���?�8�xV�<�ܰ���;��Q�I��[m��P�&�g�G��Ub���n�
�7?���^���� ���L���A)?/�*?��x?Ρ�h�0�N_K�v�=�ͽU1�<�%ؾ�B��Wп����U�G?���>X����<'{�>��^>QS>r�>[I��g���>�?�\?��?ꟾ�ؿl�Ŀ}8�^c�?��@��@?,&(�rz���A= k�>U	?S9;>��*�K����ގ�>-D�?���?�==şW�0Ӽ�>e?v��;_�F�zq��*3�=ع�=�==�/�'iJ>Ev�>�N��?���н��.>6�>n? �ip�{�\�T��<��U>3�ڽ�Ջ�5Մ?*{\��f���/��T��U>��T?+�>X:�=��,?Z7H�a}Ͽ�\��*a?�0�?���?$�(?:ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=�6ἤ���{���&V�o��=\��>b�>��,�����O��I��O��=vK�w�ο�����Qx<w�k=]���j?���b�����^��Z-����=]�4>ϰ[>�b�>��X>��f>�\Y?�[o?|��>�\�=��������q8�<�=k��{�9)s���z���P����������:	�{7��x��)�a>�N��ۊ�N	 ���"�Ji�;?TC>b�_KR�Y�m�ϖ�^ݾ�v;>񝽽J����E�H�N����?q�.?����d�y������&�=�7|=�&p?��=��Ǯ	�tTl>A���ː��p�=�g?",:��%��P�|�?l?�o��C���tUK>�!������&?�`�>����i�>i�C?E:C=�ye���>�.��� ?ڥ?u"t>�a��T˽˛)?�HD?&����
�ur&>�G��r��!Q<XI@>�7E�@����>��>7x�����/�b�׺�T?�>y6,���w��z�^�=�Zx?��?�p�>ߘh?ʺE?�Δ<&+��ąN�r!�嬍=Z�X?�"d?��>U<���;���#o4?ݠa?:�G>��d��h澃�.��^��v?�j?�y?n����[z�gC���H�%�5?��v?�r^�zs�����2�V�\=�>�[�>��>��9��k�>�>?k#��G������wY4�)Þ?��@w��?/�;<��V��=�;?i\�>�O��>ƾ{��������q=�"�>���{ev�����Q,�^�8?ڠ�?[��>"������QR>ilǾB5�?�j�?}�'��	f=�q����mQ��{<�I>��&=�C<�aܾ�a��7����*��|p��tW��Å>/,@���>�w$�.7�G����釿xS�}����3�>�>�_&>v�7��|k�$ZB�v;��} �|����>!J>�п��u��&�v�{�6���+����>b���߂>:�b������휾�� �;�>�>o��>6нH�����?�=�s�̿H���k��Y�V?���?3�?m�?���:,ņ��sn�,c�Ű??�bk?`_?�a*�k�m�,E�N�j?�F���5`�z4�QDE���T>�(3?E�>��-�l%~=�>!3�>��>E/�ԟĿ�涿�����?��?�꾉��>���?��+?-X�2C��1j��n�*����GA?˳2>[����!��&=���Ѷ
?Z{0?�� !�[�_?(�a�O�p���-���ƽ�ۡ>�0��e\��M�����Xe����@y����?K^�?k�?յ�� #�e6%?�>a����8Ǿ��<���>�(�>*N>tH_���u>����:��h	>���?�~�?Pj?��������U>
�}?>��>6�?i��=j�>�=����ڨ6�^]#>;��=p?�(�?��M?�T�>��=PC8��%/��F���Q�w��a�C��߇>��a?�qL?��b>�:��\j3��!��{̽��1���z�@���-�{޽#�5>y�=>3>,�E�� Ӿ��?Lp�9�ؿ j�� p'��54?.��>�?����t�����;_?Pz�>�6��+���%���B�`��?�G�?>�?��׾�R̼�>;�>�I�>C�Խ����[�����7>0�B?X��D��t�o�x�>���?
�@�ծ?ii�?�/������'�VO���6���=��8?����y>-��>ۅ�=�Fv�1٪��Vr�|�>H�?ܘ�?.��>Y�l?��n�g�C�)v(=Jا>��j?��
?�� ���O�;>��?Ǧ
��e���#�d�b?L�
@�h@�U^?+w��w�߿Z(��Ѻ�ZtǾ%��=IQ4>s5�>�a�k^=! ������������c�>b�c>Z>\Y>�^u>�Q�=�!������坿b{��L\/������K ���4�?v�f����s��%Ͼ�龨�ԽU+O��ؽC1�G��~f����=�P?��g?h�|?+/�>�}�w�~>>�����������>��~>ƴh?��{?L�/?�qż�;��/)?��_�����$���;�>(+�>_I�>`P�>`�?���=U�>�,ݼT�.>Bl>,�ּ�r���r�=i>j^>֡�>'��>9��>xt>�{��A� �?�3�ּ�`ѽ�?1�ڽ
�y�C����v�LO��A��<�8?��>�����޿֎��"�P?�R��d�����K��r=d ?�*�?f�6>���S����X=����i�>�N��뮾7�<�.5�>a��>�8!>���>?�?�yS��".�$�x�A���K?%o?=�F�=h��Vd��3Z�9J�=y��>w��>:8#������Y��������=��;?I|
?�Խ��Ҿ���]޾d2n>v�I�4��=C����;H>H*��s�=ە�P{�=��l�đ�=�u?�5.>��x==�>�%��<UP�T��>�rB>�t*>~�:?QD$?Q���[���C������Uf>���>�f�>��>�I�]��=�'�>�fb>�݋�od����@$C��C^>�!��6Ec�x�Hg=�}�� >Y|�=��tT���=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾOh�>yx��Z�������u�u�#=P��>�8H?�V����O�g>��v
?�?�^�੤���ȿ4|v����>W�?���?h�m��A���@����>;��?�gY?soi>�g۾=`Z����>һ@?�R?�>�9�}�'���?�޶?֯�?+I>��?��s?�j�>hCx�sZ/�*6��1���r=�f[;�e�>�^>����LdF�Q֓�]g��Ĺj������a>/�$=��>�R��5��'P�=���J����f�]��>�%q>g�I>�V�>�� ?�c�>]��>i�=�v��g瀾�����K?���?���D3n�k��<��=�^�j+?P4?9=Y�G�Ͼ���>��\?�?p�Z?ms�>_���?��㿿⇴����<��K>b>�>�=�>iK��i
K>��ԾD��U�>7ї><5���1ھd3���^���>~d!? z�>U��=� ?��#?`�j>�H�>e�E��8��.�E�[�>x��>�Q?b�~?�?i����G3�W���ڡ�d�[�i;N>Y�x?�K?9��>x���م���LB�/�K��6�����?eZg?�|��?�0�?c�??ӹA?�0f>'#�!�׾�ʭ���>۷?����f�U�T=�xd��?��>��?���%~=�DJ�{�������"�>�1?}�_?�o ��I`�O���=�Y=�cj=oM�<����م�=�2/>�~��u>6%�>P��d�ؾ�F4�j�G>�_�=ŅZ> �ȽIt�Օ^��<,?��G��܃��=��r��wD�=�>3ML>`���^?�m=���{�N���x���	U�X�?���?�j�?�����h�y$=?��?7	?�!�>qJ���}޾ܔ�Ow�Xzx�x���>A��>�gl���ُ������F��7�ŽI���?���>yx	?3��>h�=.�>Q���G�#�Djž9�ھ�yo�2�!�y%;��1:�e
�>";Q*�4�(�!�پ<(��2�/>�m�=[��>R@?�r>bÞ>z�?���h^�>=%c>�v>g��>9�[>��A>'�>���=X��
GR?����N�'�г� ����.B?�hd?S,�>Ui����b��Q�?B��?�p�?�Jv>h�(+�hn?�<�>���Qn
?�@:=Z@��߉<kO��_��0,��������>"p׽O :�@M�cf�9i
?�.?Xݎ���̾�@׽ˇ����n=,N�?�(?��)���Q�ǽo��W�9S����/h�'f����$���p��]���%���(�!a*=~�*?��?��������(k�x?�df><�>�'�>+�>v{I>��	�x�1�_^�}I'�͸���O�>�V{?��>Q�G?J;?YM?��I?��>?��>����-��>�i�<�֯>��>C�=?��2?�{.?̱?_�*?��l>���v���׾{?�?)?��>/�?9�u���zi�O���y:{�ip��S=��Z=����˩���=R"P>?��^�� S�H���x�>#��>HY�> ��>�3��k��$o=��?�O�>�'�=�	ھ�Zh���վ/�(?m�d?$�2�G,O</�->��	=�l���y�=+
-=c��� U>��=�X�~4��wWr>�H�=OQ~:�w�;��>ܐ�1��=V�>[�?��>���>���� ����"��=e�X>RS>Y�>m�ؾ�j��s'����g��cy>!}�?ol�?�xd=�c�=���=������U��e[��PE�<,�?��"?�7T?���?4�=?�d#?�d>��=7���I������?*gP?��~>e󾱣̾$ݑ��Y�kW,?���>�F���ٖ��B���7��H3�wQv����㾿s�I��ش>��� 2����?��?m�0���^���ݾZ����
��j?�?��R>J/?�b�&����e4���>���>�V�?j��>9;?��t?gV?�
w;��P��ˢ�������=�>�DS?�~�?��?ˣ?R�K>��>nĀ�S��;�M�k�4�PU=.G6�L�z��0?Qs�>�[�>d
�>0f=�9��w���ر��s:>&��>��'?Ϊ= b?��>m<L<��4?���>g�ؾI� �Y��t5������v?|��?�?��̼N0�[?�����ٷ>�b�?y�?�d?LǇ��>��V,ؾO6���-�>�z>y
�>l�=�����a4>u�>���>���F�CA+�����?�pq?�c=�!ƿ��q��_q��
����u<�"���e�^���1�Z�P�=�����h�?���v}[�w���ĳ�����k���p{���>嶄=^��=���=���<�ż&�<+~E=L�<E�
=�p��)h<�\4�5E���I���6��^<��B=44ٻ�N˾4>}?�JI?Ʊ+?y�C?��y> >�i7����>�����b?�'V>lKN�<3����:����t����`ؾ'a׾�lc�EL���>��N��>�\4>.�=�<dH�=kis=4�=ͅp���=Wn�=�O�=�b�=�7�=�>�>��u?:����ZBR��e��2:?L�>�=Iiľ��??��7>����o���s��|?�p�?�L�?J?�i��q�>0l���Ί�)F�=L����1>���=��1���>%AT>F������\t���P�?��@��>?�Ō��Ͽ~�5>h�
>m@w> �{�w^���^��P�����TR?����|����=�j�>�"���y)�\ve�ZN�>v�>���=�R���3>D���q��=>�l�>U�>JH�=�Y�<��<Czc�Z �=���>�ב=sx�=���6�*>G������>�>���>R?ߊ:?�%b?�&�>
��Pc��@޾�n�>���=5�>y��=rƅ>\�>��,?�.?�U?�^�>��=�=�>m�>j0&��y|�冕��e�0�����s?r��?��>�	�I�ɽ�Q�q &�]�q���?�X>?	}?cR�>���8��������x�N� @5>�_>f���m�x��]�{��Ⱦ�	�	��>�8 ?�v�>f�_>��W>�|;>Gĳ>ӄ�=���=��=/�N�Eo+�+'E�~���ZL�Õ>|��=�J���G�=�;�ꕟ���Q�s�(=��5����=�Q�=��>�^>�@�>��=�Y��2R/>�}����L����=�o����A�]�c�~�}��.�]�7���A>TAX>ͺ��r��jx?קX>��@>�V�?)�t?�k>���Ӿ�z��SLc��&S��ʵ=�#
>�;��:��4`�$yM���Ҿc��>��>�)�>��}>���XS�Ya=>b����t�o?1`��=e�)[N�}ł�c����ͥ����е!�sc?3u���QI>��f?��=?���?*�>��q��Y�>	j�[�&>K���'dþ�\�=�?H?��C?�	?�Q���Y��=�˾?|��$�> LL�B�O�`��x1���߻e:��+z�>)ϫ��bо�3�T���������A���o�T��>z�N?���?�ra�]��KoO��������??Zg?�D�>c�?Z�?���)��e��=��n?8��?T�?�G	>��=@�߽�| ?JO?�'�?���?ux?R�����>THg=��>�>��Ǩ=EO>%�!>NP{=�B?W�??~���/{
��1 ��k�8�#�U=�z�=�{~>��`>ܘ>��;�s۽�A{<�
`>6�>ճ>e�>�s>�k>��x����7/?3%�>e�S=�/?�G�>�~>�&�,>\%�+�E>S+b��r���W��<Ϭ���Ͻc�9�g$Ǽo�1>g��>+�޿Ꭳ?���>6Vt�M�\?/3*��n��U�>�W�=y[@���?Pgt=2D�>� �>*�>��=��>"J�>�BӾE�>>��Sk!�DC��zR�Ҿ��z>EN��
&���������BI�5���1P���i�e��`Y=����<�;�?�����k�T�)�����C�?�s�>l6?�̌������>�>P��>�k������ؼ�����o�?���?i:c>$�>
�W?��?~�1��3��sZ�r�u��%A��e���`�����Λ��+�
������_?�x?�wA?�M�<j;z>���?��%�6׏�F+�>/��&;��F<=<,�>Z&��M�`�U�Ӿ�þB7�JHF>ҕo?�%�?Z?�OV���<�G> uD?��E?Hid?S�6?*SQ?�Tоu.?���>Q�?|h�>��O?�2?$ ?�����j�>�Ȍ>|�t>���O��R^��t�Oe��m��={>c�<I�����<�m=��ü
C3����;�<c����wG=(
>� >bV�>�p]?!P�>A�>һ7?t��p8�,.��}�.?��6="��Aŉ��<�����>�-j?3ϫ?I>Z?E
d>�YA��7C��c>�U�>�	(>BA\>J��>���0�D���=�>�m>�=V�H��:���	��:���K�<�>���>�O|> 3���'>�{��Yz��Zd>'�Q����� �S�/�G�4�1��jv��K�>��K?��?�v�=�v�\U��)Ff��$)?�\<?�IM?Q�?�?�=��۾��9��J�'T�0�>O9�<���s���e��N�:�a�:�s>�(��BꞾWc>���7�྽zj�H�G�Q1�A8r=��EKR=�.��@о�.{�)��=˧
>r��y��o��r��O�I?��w=�/���cW�j���(>W�>MU�>if�67^��D��ұ�Vo�=ZU�>��9>QB��S��8J���\-�>�-?��f?F/�?�
�����4UG���+��^��Qo!>��?��>�? ��>��5�m�l�ع.�gyF���U����>	?�1�,S]��kýf��S�o��>T�> �[>�o
?]�P?��>;��?�->?}�?��>˓ս|Q���#?O�?�#s=��㽀zQ��]7���G����>��*?j�F�~w�>��?�?#?rLP?˃?Td>Ol���>��n�>���>�W��&��t�\>�OJ?�R�>�Y?}��?�6>U�3��Ş�Χ���F�=h>�1?j�#?��?Qq�>[G�>I ��Ӛ>��*?[�w?�@�?�ل?��@�d��>E>|�
?�ƽ��(=E=?�-?]4(?��l?gGJ?L� ?�5��iQ���+�m<���7�=��=W�ռ�F>�u<��"��J[�Ό@������k:=G =�3/���"���S�>��s>*��Y�0>J�ľ	j���}@>���#E���䊾�g:��۸=�>��?��>��#��~�= ϼ>n[�>����-(?E�?*�?�;w{b�u�ھf�K�&�>DB?H-�=�l��j����u�˟h=��m?��^?�X�- ����b?��]?�I�=�Hľ��b����|�O?e�
?'�G����>��~?�q?���>�2f��$n����p:b��%k�f��=�w�>�\�W�d�*c�>+�7?�>�>�c>"�=Wn۾V�w�ia���?F��?��?���?�F*>��n�a1�l)������0�^?n��>:8���#?&����о��������]*��A��E���Ŕ�����PQ%�B섾Nٽ���=�#?#r?Z�q?��_?���|c�;^�0D����V����s����D��C���C��bn�I���z��<���*�>=?4-�ʾa���?�z7?,�;i9?"^��s���(`����=��X���ؽ�&�������c��+N�<������B�g\K��$?�֨>q��>�$<?p�k��<��1E��N�9����S>5�/>,��>~?� c�լT��ؕ���پ�2��D��=v>W�c?O�K?��n?p���D1�b����+"��M<�ꮥ��WG>��	>e�>�L�����&�R=��r�+-��.��L����= �2?���>e��>�ۘ?y�?y��ʶ���u��o1���<��>�wi?%�>��>_	н1��J��>��l?��>��>�����Z!��{���ʽ]�>�̭>p��>l�o>�,��\�e��邎�M9���=2�h?ق��<�`�Pم>�R?��:s$I<�n�>Βv�+�!�H��O�'�U�>u?ؽ�=�;>�už�&���{��0���$)?�G?X��:�*��L~>"?d��>n?�>R&�?ܫ�>A�þd$;�q�?��^?�I?E_A?��>@�=����ȽLI&���-=Ok�>�Z>l+k={*�=?��1�[��R�#�A=Ɓ�=�μn����<�f���A<*��<�3>^޿�U�����a'�����C����Y��<?͞�6�\�)Gξ���F4���7�VI=�P����k�V����׽���?-( @�ʾ߅��e��bu���1���?�8�xV�<�ܰ���;��Q�I��[m��P�&�g�G��Ub���n�
�7?���^���� ���L���A)?/�*?��x?Ρ�h�0�N_K�v�=�ͽU1�<�%ؾ�B��Wп����U�G?���>X����<'{�>��^>QS>r�>[I��g���>�?�\?��?ꟾ�ؿl�Ŀ}8�^c�?��@��@?,&(�rz���A= k�>U	?S9;>��*�K����ގ�>-D�?���?�==şW�0Ӽ�>e?v��;_�F�zq��*3�=ع�=�==�/�'iJ>Ev�>�N��?���н��.>6�>n? �ip�{�\�T��<��U>3�ڽ�Ջ�5Մ?*{\��f���/��T��U>��T?+�>X:�=��,?Z7H�a}Ͽ�\��*a?�0�?���?$�(?:ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=�6ἤ���{���&V�o��=\��>b�>��,�����O��I��O��=vK�w�ο�����Qx<w�k=]���j?���b�����^��Z-����=]�4>ϰ[>�b�>��X>��f>�\Y?�[o?|��>�\�=��������q8�<�=k��{�9)s���z���P����������:	�{7��x��)�a>�N��ۊ�N	 ���"�Ji�;?TC>b�_KR�Y�m�ϖ�^ݾ�v;>񝽽J����E�H�N����?q�.?����d�y������&�=�7|=�&p?��=��Ǯ	�tTl>A���ː��p�=�g?",:��%��P�|�?l?�o��C���tUK>�!������&?�`�>����i�>i�C?E:C=�ye���>�.��� ?ڥ?u"t>�a��T˽˛)?�HD?&����
�ur&>�G��r��!Q<XI@>�7E�@����>��>7x�����/�b�׺�T?�>y6,���w��z�^�=�Zx?��?�p�>ߘh?ʺE?�Δ<&+��ąN�r!�嬍=Z�X?�"d?��>U<���;���#o4?ݠa?:�G>��d��h澃�.��^��v?�j?�y?n����[z�gC���H�%�5?��v?�r^�zs�����2�V�\=�>�[�>��>��9��k�>�>?k#��G������wY4�)Þ?��@w��?/�;<��V��=�;?i\�>�O��>ƾ{��������q=�"�>���{ev�����Q,�^�8?ڠ�?[��>"������QR>ilǾB5�?�j�?}�'��	f=�q����mQ��{<�I>��&=�C<�aܾ�a��7����*��|p��tW��Å>/,@���>�w$�.7�G����釿xS�}����3�>�>�_&>v�7��|k�$ZB�v;��} �|����>!J>�п��u��&�v�{�6���+����>b���߂>:�b������휾�� �;�>�>o��>6нH�����?�=�s�̿H���k��Y�V?���?3�?m�?���:,ņ��sn�,c�Ű??�bk?`_?�a*�k�m�,E�N�j?�F���5`�z4�QDE���T>�(3?E�>��-�l%~=�>!3�>��>E/�ԟĿ�涿�����?��?�꾉��>���?��+?-X�2C��1j��n�*����GA?˳2>[����!��&=���Ѷ
?Z{0?�� !�[�_?(�a�O�p���-���ƽ�ۡ>�0��e\��M�����Xe����@y����?K^�?k�?յ�� #�e6%?�>a����8Ǿ��<���>�(�>*N>tH_���u>����:��h	>���?�~�?Pj?��������U>
�}?>��>6�?i��=j�>�=����ڨ6�^]#>;��=p?�(�?��M?�T�>��=PC8��%/��F���Q�w��a�C��߇>��a?�qL?��b>�:��\j3��!��{̽��1���z�@���-�{޽#�5>y�=>3>,�E�� Ӿ��?Lp�9�ؿ j�� p'��54?.��>�?����t�����;_?Pz�>�6��+���%���B�`��?�G�?>�?��׾�R̼�>;�>�I�>C�Խ����[�����7>0�B?X��D��t�o�x�>���?
�@�ծ?ii�?�/������'�VO���6���=��8?����y>-��>ۅ�=�Fv�1٪��Vr�|�>H�?ܘ�?.��>Y�l?��n�g�C�)v(=Jا>��j?��
?�� ���O�;>��?Ǧ
��e���#�d�b?L�
@�h@�U^?+w��w�߿Z(��Ѻ�ZtǾ%��=IQ4>s5�>�a�k^=! ������������c�>b�c>Z>\Y>�^u>�Q�=�!������坿b{��L\/������K ���4�?v�f����s��%Ͼ�龨�ԽU+O��ؽC1�G��~f����=�P?��g?h�|?+/�>�}�w�~>>�����������>��~>ƴh?��{?L�/?�qż�;��/)?��_�����$���;�>(+�>_I�>`P�>`�?���=U�>�,ݼT�.>Bl>,�ּ�r���r�=i>j^>֡�>'��>9��>xt>�{��A� �?�3�ּ�`ѽ�?1�ڽ
�y�C����v�LO��A��<�8?��>�����޿֎��"�P?�R��d�����K��r=d ?�*�?f�6>���S����X=����i�>�N��뮾7�<�.5�>a��>�8!>���>?�?�yS��".�$�x�A���K?%o?=�F�=h��Vd��3Z�9J�=y��>w��>:8#������Y��������=��;?I|
?�Խ��Ҿ���]޾d2n>v�I�4��=C����;H>H*��s�=ە�P{�=��l�đ�=�u?�5.>��x==�>�%��<UP�T��>�rB>�t*>~�:?QD$?Q���[���C������Uf>���>�f�>��>�I�]��=�'�>�fb>�݋�od����@$C��C^>�!��6Ec�x�Hg=�}�� >Y|�=��tT���=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾOh�>yx��Z�������u�u�#=P��>�8H?�V����O�g>��v
?�?�^�੤���ȿ4|v����>W�?���?h�m��A���@����>;��?�gY?soi>�g۾=`Z����>һ@?�R?�>�9�}�'���?�޶?֯�?+I>��?��s?�j�>hCx�sZ/�*6��1���r=�f[;�e�>�^>����LdF�Q֓�]g��Ĺj������a>/�$=��>�R��5��'P�=���J����f�]��>�%q>g�I>�V�>�� ?�c�>]��>i�=�v��g瀾�����K?���?���D3n�k��<��=�^�j+?P4?9=Y�G�Ͼ���>��\?�?p�Z?ms�>_���?��㿿⇴����<��K>b>�>�=�>iK��i
K>��ԾD��U�>7ї><5���1ھd3���^���>~d!? z�>U��=� ?��#?`�j>�H�>e�E��8��.�E�[�>x��>�Q?b�~?�?i����G3�W���ڡ�d�[�i;N>Y�x?�K?9��>x���م���LB�/�K��6�����?eZg?�|��?�0�?c�??ӹA?�0f>'#�!�׾�ʭ���>۷?����f�U�T=�xd��?��>��?���%~=�DJ�{�������"�>�1?}�_?�o ��I`�O���=�Y=�cj=oM�<����م�=�2/>�~��u>6%�>P��d�ؾ�F4�j�G>�_�=ŅZ> �ȽIt�Օ^��<,?��G��܃��=��r��wD�=�>3ML>`���^?�m=���{�N���x���	U�X�?���?�j�?�����h�y$=?��?7	?�!�>qJ���}޾ܔ�Ow�Xzx�x���>A��>�gl���ُ������F��7�ŽI���?���>yx	?3��>h�=.�>Q���G�#�Djž9�ھ�yo�2�!�y%;��1:�e
�>";Q*�4�(�!�پ<(��2�/>�m�=[��>R@?�r>bÞ>z�?���h^�>=%c>�v>g��>9�[>��A>'�>���=X��
GR?����N�'�г� ����.B?�hd?S,�>Ui����b��Q�?B��?�p�?�Jv>h�(+�hn?�<�>���Qn
?�@:=Z@��߉<kO��_��0,��������>"p׽O :�@M�cf�9i
?�.?Xݎ���̾�@׽ˇ����n=,N�?�(?��)���Q�ǽo��W�9S����/h�'f����$���p��]���%���(�!a*=~�*?��?��������(k�x?�df><�>�'�>+�>v{I>��	�x�1�_^�}I'�͸���O�>�V{?��>Q�G?J;?YM?��I?��>?��>����-��>�i�<�֯>��>C�=?��2?�{.?̱?_�*?��l>���v���׾{?�?)?��>/�?9�u���zi�O���y:{�ip��S=��Z=����˩���=R"P>?��^�� S�H���x�>#��>HY�> ��>�3��k��$o=��?�O�>�'�=�	ھ�Zh���վ/�(?m�d?$�2�G,O</�->��	=�l���y�=+
-=c��� U>��=�X�~4��wWr>�H�=OQ~:�w�;��>ܐ�1��=V�>[�?��>���>���� ����"��=e�X>RS>Y�>m�ؾ�j��s'����g��cy>!}�?ol�?�xd=�c�=���=������U��e[��PE�<,�?��"?�7T?���?4�=?�d#?�d>��=7���I������?*gP?��~>e󾱣̾$ݑ��Y�kW,?���>�F���ٖ��B���7��H3�wQv����㾿s�I��ش>��� 2����?��?m�0���^���ݾZ����
��j?�?��R>J/?�b�&����e4���>���>�V�?j��>9;?��t?gV?�
w;��P��ˢ�������=�>�DS?�~�?��?ˣ?R�K>��>nĀ�S��;�M�k�4�PU=.G6�L�z��0?Qs�>�[�>d
�>0f=�9��w���ر��s:>&��>��'?Ϊ= b?��>m<L<��4?���>g�ؾI� �Y��t5������v?|��?�?��̼N0�[?�����ٷ>�b�?y�?�d?LǇ��>��V,ؾO6���-�>�z>y
�>l�=�����a4>u�>���>���F�CA+�����?�pq?�c=�!ƿ��q��_q��
����u<�"���e�^���1�Z�P�=�����h�?���v}[�w���ĳ�����k���p{���>嶄=^��=���=���<�ż&�<+~E=L�<E�
=�p��)h<�\4�5E���I���6��^<��B=44ٻ�N˾4>}?�JI?Ʊ+?y�C?��y> >�i7����>�����b?�'V>lKN�<3����:����t����`ؾ'a׾�lc�EL���>��N��>�\4>.�=�<dH�=kis=4�=ͅp���=Wn�=�O�=�b�=�7�=�>�>��u?:����ZBR��e��2:?L�>�=Iiľ��??��7>����o���s��|?�p�?�L�?J?�i��q�>0l���Ί�)F�=L����1>���=��1���>%AT>F������\t���P�?��@��>?�Ō��Ͽ~�5>h�
>m@w> �{�w^���^��P�����TR?����|����=�j�>�"���y)�\ve�ZN�>v�>���=�R���3>D���q��=>�l�>U�>JH�=�Y�<��<Czc�Z �=���>�ב=sx�=���6�*>G������>�>���>R?ߊ:?�%b?�&�>
��Pc��@޾�n�>���=5�>y��=rƅ>\�>��,?�.?�U?�^�>��=�=�>m�>j0&��y|�冕��e�0�����s?r��?��>�	�I�ɽ�Q�q &�]�q���?�X>?	}?cR�>���8��������x�N� @5>�_>f���m�x��]�{��Ⱦ�	�	��>�8 ?�v�>f�_>��W>�|;>Gĳ>ӄ�=���=��=/�N�Eo+�+'E�~���ZL�Õ>|��=�J���G�=�;�ꕟ���Q�s�(=��5����=�Q�=��>�^>�@�>��=�Y��2R/>�}����L����=�o����A�]�c�~�}��.�]�7���A>TAX>ͺ��r��jx?קX>��@>�V�?)�t?�k>���Ӿ�z��SLc��&S��ʵ=�#
>�;��:��4`�$yM���Ҿc��>��>�)�>��}>���XS�Ya=>b����t�o?1`��=e�)[N�}ł�c����ͥ����е!�sc?3u���QI>��f?��=?���?*�>��q��Y�>	j�[�&>K���'dþ�\�=�?H?��C?�	?�Q���Y��=�˾?|��$�> LL�B�O�`��x1���߻e:��+z�>)ϫ��bо�3�T���������A���o�T��>z�N?���?�ra�]��KoO��������??Zg?�D�>c�?Z�?���)��e��=��n?8��?T�?�G	>��=@�߽�| ?JO?�'�?���?ux?R�����>THg=��>�>��Ǩ=EO>%�!>NP{=�B?W�??~���/{
��1 ��k�8�#�U=�z�=�{~>��`>ܘ>��;�s۽�A{<�
`>6�>ճ>e�>�s>�k>��x����7/?3%�>e�S=�/?�G�>�~>�&�,>\%�+�E>S+b��r���W��<Ϭ���Ͻc�9�g$Ǽo�1>g��>+�޿Ꭳ?���>6Vt�M�\?/3*��n��U�>�W�=y[@���?Pgt=2D�>� �>*�>��=��>"J�>�BӾE�>>��Sk!�DC��zR�Ҿ��z>EN��
&���������BI�5���1P���i�e��`Y=����<�;�?�����k�T�)�����C�?�s�>l6?�̌������>�>P��>�k������ؼ�����o�?���?i:c>$�>
�W?��?~�1��3��sZ�r�u��%A��e���`�����Λ��+�
������_?�x?�wA?�M�<j;z>���?��%�6׏�F+�>/��&;��F<=<,�>Z&��M�`�U�Ӿ�þB7�JHF>ҕo?�%�?Z?�OV���<�G> uD?��E?Hid?S�6?*SQ?�Tоu.?���>Q�?|h�>��O?�2?$ ?�����j�>�Ȍ>|�t>���O��R^��t�Oe��m��={>c�<I�����<�m=��ü
C3����;�<c����wG=(
>� >bV�>�p]?!P�>A�>һ7?t��p8�,.��}�.?��6="��Aŉ��<�����>�-j?3ϫ?I>Z?E
d>�YA��7C��c>�U�>�	(>BA\>J��>���0�D���=�>�m>�=V�H��:���	��:���K�<�>���>�O|> 3���'>�{��Yz��Zd>'�Q����� �S�/�G�4�1��jv��K�>��K?��?�v�=�v�\U��)Ff��$)?�\<?�IM?Q�?�?�=��۾��9��J�'T�0�>O9�<���s���e��N�:�a�:�s>�(���+ξ�=Ṋ��!�������M�Ch���f���(�x�>X�O�`R������6;�>�mE�X�ս��5��t�mM>?"�=��þyվ�[���0>�v�>xq�>^� ��2�f'O��5����=���>]�^>֕=�9���\���;��>Q�N?*�g?���?�u[���_�w�O���)(���� =��1?ͥ>�q�>1�
>Ͳ�=��˾�i���)��%�i��>*?yk��n-z��0꾸���)�6�}>?�?��C>��>,�1?��>���?�a(?��>T�>Y�ǽ����?V*?_�=}^��yZ�k{��#�f"�>F�?g0{��2�>�>>yp>4�L?�R?��>�e�=㟻��&E���>��X>�.b�9����O>oS?c?@�<?2)�?����4�(�(J��#E��E�.>���>�-?xq?�>�q�>9_�>7Q�<۽d��>Hge?�{�?���?�n�>d�"?�P>���>�G�;y�>|?3fE?�^g?,�?�PU?��?�;<h{����F��ݨ��d���&��D�;h�=�����Α��i<����=��=���;=,<A�<� B���<.{�<�e�>�s>~���j,1>
_ľ�3���?>�M��E�����d9��i�=��>:�?/1�>G$����=��>���>e��{�'?P?��?�;5db�0۾q�K���>p�A?�,�=&^l��D��i�u��\f=Cn?ȯ^?�V������b?��^?m��ض;��þ}d���/DO?`�	?�G�	�>f
}?�4o?�D ?,H`�Kdo�L!����_�6�n�U>�=X��>���6,f�Ւ�>�X7?߅�>#ne>-��=0"޾k�x�w����	?��?Ϳ�?>܉?�b*>�n� p࿢]��r;���^?#�>G畾9T#?Q�Z��?ɾ�Ɋ�	���wپ����������cR������r����3�=t�?�*u?��x?��b?[����f�~g`��:���nV�K���2��D��zD��v@��i���� ��!����]=�b��7C���?��?��ͼ���>�Ԙ���ʾO�ݾc�g=�%[�V���s�=��N��q��cG=����W������A6?���>q�?��@?7�m�
R���A�fJ�}N�φ�>ċ�>���>y��>�*��g��FN�r�龐�L����� �>��_?�LV?<Ղ?��N���$��������������^�>�jG>�n�>j?��A��u\D�y�"���=�/�پ|ㅾ�������g?�a�>�	�>�+�?}t-?r�������վ5�~�����l�>	�O?�j�>D�7>�d�����)��>�o?�c?�ܻ>\�����"��х��;�n��>S�>)?3�>)�ϽP�_�,W��%S�������N>Oe^?����/�G�j>�8a?ID�;K����>��7(����f(��U�=7P�>���=��w>^�Ѿ���^�s�V�`���!?��?؝���.6�!/5=Mk�>$?��x>�.�?%�A>�n��X�N��.	?G\?��I?�}P?�Q�>�/�ёF��̽��ʽT�>y�s>_Y�=\9%<9��<��i�,	��zý[�<i� �G�=���;����=+�,��O�<�L>g��.�D�s�ľ����:	�_�H�s�\Q�	蕾
q�e'���D��ԬS��C=oBǽ!ݨ��Ͼ��������?E�?����oݽ��y��_����=�f��9>����i��*������nHپS�8��Ts�&�z�`�+?������ȿOC��̜پ�?&Z0?�{?]���[�+���9>`N�=�Ÿ���ھ~㓿!�пTqh�Aq?��>E������÷>E�d>>�g>�~d>r�u�����/T�׻�>o�"? ��>汙����F���$��=��?>�@b)?�DM�v㻾iP��5�+?k$?�G>�rG;t������3?�Ҧ?ڊ?��Z��^\�I�(>O|u?P>T>�(��ˀ��ج�˺K>��x=�
��\�2>�d>��F�W�����n>�!�>U(�j�P��Y��Z0=�qf>F�C�ի�(Մ?{\��f���/��T��.U>��T?+�>�;�=��,?O7H�Q}Ͽί\��*a?�0�?��?#�(?:ۿ��ؚ>��ܾo�M?VD6?���>�d&��t�#��=�6�,���U���&V�N��=;��>�>�,�Ƌ�ǇO��H��k��=�s��'пL�0��L%�=��^8<����?wx�/��^����U����N��'��O�=�X�=��4>A�R>�tI>,�i>�[X?�5k?*3�>�h1>,��D��R�ľ���QD����4<��'A,�����m���D�j>��a� @�y`��6|?�!\�=�M������%��c�/4C�"&?2� >[g���|P�~>�;;�Ծ�����⼊ji��Ծ94��^l�;��?��;?���
W�?F�Ȏ��Y���h�V?��
����=��ޘ�=)`-��C�<EÜ>݇�=Qؾy�/��,S���/?ñ&?�챾�A����>.X���A�<�L?b�?M�E��ƨ>�?�fI�����C��>fD>���>@�>�a�={R��<�˽7"?��N?�½x���҂>�FϾ;�S�O��=�=�'�퟾;cm>����b���#;H�6��8d=�^W?���>FPF����w���C��u|>�dn?�]?��>V�X?B�;?�?+>�Ͼ�.��@پ�y�LEY?N�|?u{6>J�"���پ92оFu?P#P?�.�>��|��hھH�"J�R��>��A?nC?��Z�k6������W����k?Hnu?6&`�+����O�u�J��B�>�|�>�*�>�'8�a|�>�??ص�������R5�T�?�j@P�?��5<�F!�弋=�?�w�>MR��	Ⱦf����_���BQ=��>����l�t�����-�7?�Z�?_�>����R�P2$>��I��4�?ݐ~?)����~�=�6��J�������<���>[��>n>�f5�
2�����_[v�]�=t�=聚>��@��>�6?;r1�8��riϿ�����s�����>-�D?W� ?0�=C�3B3�Xy��D�5I����U�DC�>�>>�"��e�z�g��k3�(7z�"\�>ܻ+�-�i>������t}����a=+�>d��>xv>e�������?ܳ��L̿���K���[?�s�?��?�?�	��`!������*i���N?x�h?��K?��7�n(��h��A�i?�:���Af��1�ab1���:>407?��>�/�/G=k�=>G��>��>�wL����������F����?���?i�ݾ%>�>��?6�)?��ľ�#��� ��*��l�=a�"?�͏>��R��p&�7�;��#���o�>�tG?0fٽ����_?�a�q�J�-�ZFŽ�$�>7�/���[��~��5e������x���?be�?�	�?)��w�"�\J%?ǯ>Ҿ���WǾ-a�<�6�>��>��M>c�_� v>���%�:���	>r��?�t�?�w?Zo���樂D>��}?�9�>Sj�?>x�=H��>�m�=~��������5>��=%����?�oL?�Y�>
��=�`@��/�ПC�xDP��U�	"B�O�>`?! K?�2_>�����;������Ͻ`�5�P���^�8��3,��4�|�3>�7>&�>�V@��Ѿ��?^m�F�ؿ1g���c'��04?_��>q�?h��c�t�|�j?_?�y�>79��(���&��K�I��?�G�?9�?u�׾�˼~
>��>PJ�>UGսV���,s����7>��B?~��?����o���>���?��@�Ү?i��

?���ge��1s���������;��4?9쎾]w)>�?c�6>��O�f���	sj� S�>���?E��?yj�>ÐI?S�t�X6�� �K�?���?�?��u=PJ��y�$=�
�>9����y����%L?�@.�@��H?aL�����!歿/���ᴾH�=��>��>��B�hi5>~����Ƽg	;F@t>|1�>+M>�3�>�>>�w>5HT>�Y��������"�����=��@���ھR�#� ]��@���� �]��Y�ԝ��S�潫2Ͻ�y�����J��%g�=�T?��Q?��l?|3�>A����Q>\���Ɣ�<���g=�)�>AR1?��H?0L'?���=�����c�qZ��PN���Ƈ�[��>uKO>z��>)�>��>ݎ>�h�B>�n4>�v�>��>��F=�It�+>�<#�L>�2�>��>���>Y:=>m�>����3��	�g�A=����ֽ;�?�5���-A�o����@���ش�$�=>�.?x�>����i�пի��D?���&���!E�h�>�x1?�T?g58>�i����%�Ѻ>����\c�$)>jߧ�J�f�����$U>��? ̪=��W>TT��#W��l��5��+_8>���>}��f�>���[� ���S�>	7>2>�i��Re�� n�Q7?���>�y,?�?�ǉ�ٻ��ۦ��h���Mb=z��>�\�>�ai>�W>c�8��5�5)���Pq=쭄>SFV>���>�V>�R3=eϠ>
ے�9lv���>��=8> �7?=�?)��;���[q��.Wb�w�`>�a�>U�n>E�=�=,�`��=�*�>�;> {����	�ֽ���}b3>f�`��o� ��7=*ۃ��=~!t=4��&�����o=�~?���)䈿��e���lD?U+?n �=ɞF<��"�D ���H��G�?r�@m�?��	�ݢV�@�?�@�?��D��=}�>׫>�ξ�L��?��Ž1Ǣ�Ȕ	�/)#�iS�?��?��/�Zʋ�;l��6>�^%?��Ӿ���>�c��^��F���u�<#=���>9;H?
"���7O���=�y
?�?�?򾫖����ȿ�v����>A�?{�?m�m�U8��@��Q�>'��?AhY?��i>�h۾�iZ��[�>Q�@?�Q?���>[,���'���?�۶?���?�i1>�h�?_1S?|o�>���A?������z��������>��>K-`>�V���c�T��AE����%��f�#xn=�;]v�>�]	�����i=�Wd�Hh��v?;���>��=[�8>�6�>���>�Z\>i�>u�	<�~��:a�MLx�kK?���?c��n�n��Q�<�t�=�MZ�g	?k3?��㻝RӾ襦>[?P]�?�[?4e�>��j����i���w��<V~O>���>�e�>����H>Z3ӾG�B��!�>�p�>������ؾ{���3��q�> P!?n��>2v�=� ?�$?��m>�&�>W�D�P����PF����>�>�/?�f?��?p���X�2��L�����m[��"Q>GKx?<,?� �>�{�����ÒZ�=���:�?�;g?��2g?���?*�=?pTC?�g>�`�$X־o	���y>�?ќ�;��7�]�<�j�J���>u>�>�b?���t9D�	p�m�����N?��x?F'?v����8`�_���vW=�	�=�z=�ud�ʊ�<�%�>�Q>��@�v5q>�^ >Q�>�g�L3���@���%�=P��> �l>!�׽��)=,?C�G�Wۃ���=r�r�)xD���>�IL>����^?Ml=��{�����x��:	U�� �?���?Tk�?o��9�h��$=?�?a	?}"�>�J���}޾N��"Qw��}x�ww�G�>���>��l���A���ՙ���F�� �Ž	@��ö�>�A�>��H?��#?Ju�>6�>��5���G���O��em��{i���2�2<'��B��f#�|�Q�X�X��<Yn����m�.3�>]����>��?�ˌ>N-1>�}4>��@<H �>�>O>� �=g�1>���>iF:��Q��Kx�ZPR?|���f�'����寰��B?7�d?�_�>܁h�uv��ʭ�E|?t��?(Y�?�/v>Vhh�v\+���?`��>���nJ
?or:=�K�G0�<T��q�� ��ps��s�>Tg׽�:��M�}Gg��L
?��?4ܖ��S̾aսF���2n=�s�?+'?��*��qR�2
o�B�W���S��ü�|h�����8G#��m����������(���=gz)?9͈?z ����A����i�Dj?�#Gc>1�> z�>���>�U>��	�9�/�rS\�1'�^;}����>{�x?$7�>@pL?�M:?�J?h�F?���>�ܟ>�ΰ�0a	?�ż�B�>��>�l,?�Q)?x�-?�?0�'?'�e>0��Ą �v־$�?�!?e_?d?<�>�Z��f�������X���u~��i#�EBw<3;�.�����<���B=��Y>�N?k첼��A��¿�L*E>�?[4�>Z�>�E�ظ��=��<j��>��:?�! >I
���G��o�;l�>��x?ڣֻ���<��=��C�s�ݼN�!=��=3��*!=.��ܓ=L��<ޥl=�݈�ގ�=�P=��=���=i�>v�?â�>8��>����܌ �/�����=pX>�qR>x>RپUy��_����g���x>k�?�t�?��g=�*�=�u�=�>��Y��m ��*��@7�<��?�G#?�}T?�?��=?*t#?�O>��I:��F]���墾�?4�+?���>����̾�H����1��S?��?��^��z���&�������½���=_!.��2|�ऱ��?�X�<�>�..�����?[�?���i5����TE��	��$y@?���>���>��>T�*�� e����{U>>�>h�O?~��>�&\?�)�?!wm??=>�F6��߳�4З�
J.�,p7>3d_?� �?/�?�H,?�8�>F��A�3��1.�����g(��)ʽ�ɾ�V>�h�>�	�>���>G��>䉲=�6c��&�>¾B�5=3��>��?¤�>0)�=i+=#1�=��F?�#�>��������!���Dt�
G�)�u?�%�?6$?�M9=T!�W�@��5 ���>�~�?���?2�+?e5S��\�=�8��U���8w��>Rc�>�O�>�ɣ=�#=e.>�m�>f��>�)
�"���7�g
�;1?�xC?+7�=�ӷ�6�L����ﴥ�I����ƾ:;���KM�5꒾c,_>Ç����ڽJ��^���i;��z�a�Ⱦ�2¾`T����?��=���=��<��g<%��<��<�Ȉ=Ph�<����z�i�=ڏ ��LP���"�"J�:_�=��H=(�v��!����n?��D?��?��?���=e0j=�c��)>�¼���>�Jy>���Zp��_e��ƾ��~��{Ͼp<�>�G�B���BH�=@�*����=I<>�z�=5^	;ʌ�=`��Ν=���<�9d=��y<�3�=�x�=ێ=� �=N�>*5w?m���J����/Q��=�y�:?�9�>5h�=E�ƾ9@?E�>>�2�������d��,?���?�S�?��?Jni�%c�>g��:���dw�=����dA2>(��=�2�ȡ�>�J>����I��y��33�?^�@��??����ڡϿNd/>H>q�$>�$I�R�8�A����&6=��?�T3�򒾑S�=��=�Բ�Gp��i�> �o>��<�ى�W�R�;f�=�)��?�<Vn��kF�>��_>�>��_�p�=��=%�>�/>[��W̑�`i=�J=0>'>��>pH>&��>�?%�.?�Wc?��>�Tf�}';���Ƙ�>֒�=[��>�=0]=>���>|�6?F�D?{�H?�S�>x��=��>�>��,���l�:#��P��~s=�v�?$�?-�>q�;R�C�0��n[:������)?��/?��?�s�>�����俬�+�Ъ0�������<��}=�(Y��cT�אl�|�
��Fν�=T$�>��>ڗ>��f>^C7>�KR>N�>�>�t'=��=�S��v��<j���TxH=�i��ё
=�x�Mz	�vN�7��0�ǲ
���<z�點FZ��KP<E�	>X��>u�>4{?�92>��L�x��=ɔ����@��� ��O��#F���a�Kww���(���B��f[>�Dd>��/�����G�>�\>{�>���?b҄?6T_>@��ۥ��3���s��;��
mU�ͼ�p�M��żK��V_�L����
�>�?v>0�>Z@>� �(5/����䴾�9���>�.����=;��E!s����2��ǿ_���
>�g?}�|���=�O�?��7?!��?CC�>ґ��n¾���>nh����=�۾��(�;���>�qD?��E?�4���ԁ��H̾k��7ݷ>�BI���O�u�ԯ0��!��η����>t�����оy"3��e������m�B��Qr��>;�O?^�?K4b��U���SO����i%��4o?{g?1�>:I?�A?����z�So���u�=Q�n?=��?Y<�?��
>�}>������:�YU?���?��?�4�?���>��?��m�\D>�P���<�e�����>Px>b�\?7�?ߒE?�U��E�b�6���ɾKs3�Ή���>8#?�3�>5�>������=��>!�?Yw�>4`>���>���>���>;S��s ��&?���=⑏>�2?�-�>�V=<���Z�<3?�)B?��C+�|��sr�7��<v�X�/kT=�iʼE�>�AǿBh�?&S>����?�b�0�&��Q>F�S>@߽�M�>6DE>k�{>�>���>�>�Ŋ> .)>��Ѿ��>Z��2!���B�8R�6pϾ�.{>to���X$�g��U���E��´�o��$i��0���4<��.�<��?�� �N�k��*����J]?cߪ>�i6?X����M��vF>C��>q�>I���	���΍��>�V6�?D�?<pc>Td�>�"X?#9?�-��?-��Z��Ev��A�c�d��K_�|ٍ��΁�k��{½%`?�dx?��@?D@�<�wy>O�?a&�8��� �>%�-���9���:=<U�>����N�_�R�Ӿ�aľ�c���H>��o?B��?�?o�S��l�I�'>>[:?��1?�t?-�1?M?;?����$?�2>�"?,t?ڌ5?
�.?I�
?�2>���=�E����(=���Ê��6ӽ�&˽�0�<�5=�|=	���,<�0=lƧ<�H�Ӽ(�:� �v��<�6=@n�=)k�="��>[�[?�W�>Rf�>�8?}��q5����g(?�6=��e�Ƒ��t��e�����=��i?�\�?�R?�X>�A�$N��[>j�>/M>��w>Fl�>��:�d�|��=��>��>��y=�m��[w�E��Ǽ��E����K*>Z��>�6�>d_>��5p=ެ��i����=ꍌ���K�w�ʹ�o;�*R �<�V0�>��?��?�FR=�����J��I���>�F:?���?-m?��z���nO�R��w!=��>�&f>��پ%*�����]�I�
qż3�>��m�05E����>�Eʾ�پ.0���j��������.�Y�>x�"���Ƚ+Pb��?jߵ��z��-���2���Ŝ��c&?7�2:޼Ҿ�Y1�p%����8>y_�>�.>��5=zQm�ɭ	��v��*�>V�@?���<��
>����(�
�ܾd.�>QD@?H�T?�
s?����/u�w@����ޫ���J=��?���>���>�Ԇ>=�6������Z��pD��E�>oo�>X�� kB�-2��O۾V&#�2SX>���>>�~?��F?�7�>�iM??Ng�>�k�>��½�}Ǿ�R)?`0�?��<`
J��2!�W�)��I��&?7B"?AuR���>i�?��>�C$?I�W?g�
?�L�=��Z�8�w�>#Ӈ>��[�����3a>E�:?�$�>�	]?�$�?$1�=�=��ށ�(t��>B�Q>��H?x>�>l�?p��>�H�>�\��9Z=P6�>BI`?�Ʌ?J�n?�U>��?�">��>��5=�D�>�o�>��?�CL?
�x?:�H?~�>,��<6�ɽ���jB���+�4Ҏ<�����=HN8���M��JT��";=��~<Ƽ'l�;��Y��zD�<l�;
_�;���>:�r>:�����4>�8оi��͞:>�C�����\���=� 
�=���>�?2��>V���"=Ѫ>M�>���l�)?N�?�J?pլ;kX�V	�;om���>aS7?���=+�d�gs���~d����<"]?if?�fG�F����b?�d]?5���<�k¾f?b���_�N?�
?�d@���>�v~?�oq?Y��>��_���k�݋��XY`���]��%�=��>���e�7�>*�7?Y��>X[f>��=FR۾�ay�m���)[?��?@��?t�?��'>��n�.}߿7����WwI?��>��ɾ[-?Eż5궾��_��^�*	�������ž5@˾B���M��s������G�=��?�n?6jx?��`?+t�$�W�"ua�l���M�jP������3�PQ�6=�6i�ep&�H4�!�۾OwἋzM��C��S�?(G�>]x=C�?�Y���a��M7L�9��=�l��3L4<��9� 罀|<>J�#�b��ޖм�8���L?�?&�q>rzE?�=~�lb�i���T����
5>>�P�>���>��>[�������g�)�K�t���c[�=M}>�Z?K:?ݶZ?I;���� �*ĉ�����)���UV�>�1}>�6x>ɏ��/�8���,����U��/������k�����<nC6?�>���>���?�?bW8���`�Y�-Xc�x�s-L>&>E?��>U>�BҾ�����>@�g?3�?-�>������z�o�ٽÛ�>+2>�~?qH�=H��1Y��R��!������v!>aW?�=���U����>��G?)��;΃0>�>�Xx�3#6�:]ؾ{<��2�=d��>�k)<ݩ��ht�������o�����A�)?��?�n��4�)�l_~>{T?Y�>�ª>�~?�Ŕ>� ����Q;6�?͔Z?�F?ŒE?	�>ԃ=�z��Ƚ̜%��WF=��>x�G>:�?=M,�=~P$���R�W8��j�='�=m�Ļ�}��ց⻃,r��x</e1=�2>�5˿�<�5�	�A>��?�+���"I����=ifN��������劾�gG�UH� ��#��������+��G�? ]@�@O�+������`����ƾ�>E�&��П>�7��*uλ�Z����������ݾ"XX�3�W��6�<�&?�?����ǿr���t޾��?� ?$�v?�?��� �jA8�� >3p�<W�u��1�R[���PϿo򜾝�^?]M�>*�𾠠����>E��>z3S>5St>�t��������<��?_�-?;��>A�y��Yǿ������n<Ŷ�?��@a�??�h�E���q�=���>1L?�7>�H����Y�����>r�?ˍ�?�4)=1�P�ѭ
� �Z?٨�<2�3�����=�=A&x=������3>�̍>V("���N��6���W>d��>��C���5�?�H��Ǻ<=�1>������O��Ԅ?vv\��f���/�R���Q>��T?�(�>`*�=`�,?�3H�gyϿZ�\�$a?@0�?��?��(?ֿ���>�ܾ�M?0C6?Q��>/e&���t�AB�=s�q���d��1$V���=Դ�>>~>+�,����rO��5��"��=���{�Կ~{&��7��a9=y�=m���K(�K�=��Yȱ�����,}c��&ԻYi>�,p>���>�l>�d#>��]?��m?�ܐ>�d�=���W���u6��	uսݭž�����l��\��!"��K���_1Ⱦ��	���� '���%E,�v��==Q�.���ҍ��:W�IMG��d7?+�+>v�ɾ�I����<$J�)=����<B��;�վsC&�#If���?�9?>i���uY����@2�`���BT?����P�����b�>�|����=闣>&>m5	��	%���L�Ͷ4?�?�۾14���V>�@�����=�)?��>�*�=h�>8?�Y�4(���>T��>M,�1<�>X�><ͭ��Խ�%.?��j?�?�)ޠ�Rk�=Pc߾�g���=+�/>a���4 >2F =g]�<҇ʾ|�=��<�-��TR?���>J�%��b쾜���?��4�/>�0?	r�>�?��?�a[?��>�l��x�%w���[X���]?���?i�">"K׽��⾪MԾ�� ?�wU?}L�>觽��޾���Q�;��B�>�#%?`	�>YH�=!�F��W��0��{ ,?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������%>2���ɸ?�p?rW-�pM=��=���>��̈́�����3�=��_>q�߽2'��j�뾼��#��1~����ǽL��>��@�to��?��Ҿ>I��6⿍�g�L����ݔ���L?/�>�?�8q�s���M��q�� ����I�;���>0�U>B'�T"���LP�B������i�>+�����d>�1��ʸ��������<��>=�>�Ib>�������C�?����5Iɿ;q���7ﾲ4?L�?��?�n,?5�=aɾ�����=yXN?4؅?�w?ͯ��L�c������j?�[��gV`��4��JE���T>k"3?59�>Q�-��K}=�>Q��>�z>�/���Ŀ�Ӷ������?T��?�m꾎��>#��?z+?g��6��ed��J�*��.��:A?02>q}����!��#=�tϒ���
?a�0?�i�W4�e�_?֘a�G�p�[�-�O�ƽ�ۡ>��0�Z\��7������We����Hy���?�]�?��?���J�"�%5%?��>ޝ���:Ǿ���<���>;'�>�+N>�-_�3�u>J
���:��j	>U��?�}�?j?֓������Y>��}?ʱ>U[�?��=��>m��=óľ��o�>L��=�ڙ:���>��O?{��>��>Pd@���(�3�G���Q�!�{k?��"�>�)g?��G?�Z>ߓ��+�����$�<��2�2�����&2��w����N>+T">�dF>38�����?Mp�9�ؿ j��"p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>A�Խ����]�����7>1�B?Y��D��u�o�z�>���?
�@�ծ?ii��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?hQo���i�B>��?"������L��f?�
@u@a�^?*�俿��Gž����(�<l��=��:>�w0�E��=d��<l}�ur����N=��>Y�>|>���>���>��>S9��/)�V��?����KU�	����Xξ$��W���u��������d���\�4�m�6���.���ܽ��齩�>�FO?ͪ8?D_d?���>��⽋s$>�m �4j�U��t��<��t>X42?uH?Cq?���=���)�i���~�,g��8m����>("G>p��>�o�>�A�>LۼH�>��8>� �>aM>z�=D[G�6<��6>xM�>�i�>�^�>^�<>� >@���|*���Hh��y�y=˽١?�͜��@I�t��������>���+�=t�+?�#>	w���rϿ�լ�GeG?����Mc�p�.�K�>Y�.?QW?�.$>�Ȱ��-T��>�!��g�<��=��f��G+�I8U>?P�j>&ݎ>��*� #�'f��Y�H>|�>%�����"�L���x� �凵�w'	?�(B>�� ������{w��c>���=�?u��>�SN;낔�;⍾�ˈ��?=�1g>�J�=�
)>Tl>����^\ ��Z�		�=K�= $�>� ?��>���]�>
����`��i�>���O���Q?��?|H>5?����L7�h*�>"�>�_t��?>�o6��q�=u�>��)=���=�>J�� ��L��5a>�d��=_j>���=_�횾=߾༇�����=n=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ!`�>�c��\��R����u�w�"=g��>�#H?#Y��^6O�0>�p
?�?O<�-���O�ȿ��v�l��>���?=�?��m�A��[@�Ǎ�>���?gY?S�i>�z۾�&Z���>]�@?q�Q?E�>e��'���?�ض?���?�v=>���?3�g?X��>7s�86�//��N��A��n	�=*j�>��@>'����S#�_ᐿ�^��+�U��k���>��j=��>Z н�þ� �=ĳ �����Zj����>�XA>e>���>M�>��>"(�>`9L=�d����R��XK?E�?����l�?�<Ķ�=�J^�-?��2?uD2��Ҿ�>L[?�~�?�Y?��>r��/�������泾uؚ<pXL>���>k��>�Ƈ� VG>�
վ�lF�);�>�Ę>�q���^ؾc܃����oq�>�7!?JE�>���=�r?tD?ʏh>H��>�9��|��WZ��}�>���>�-�>&s�?�Q�>B���:��Q�� ���4,���,>�d?W�(?��>O����M���م�܄��)��Xr?!�i?���=A�>O�?h�;?��Q?�$�>+Y�:6�ྜb����>�0?>Ni=jQ�:�;��Bt<��>cn?H�	?���~=�<�-ֺ�ݵ����r��>
1Z?�Q?k\������=�5=/:ѽ/0��� =+�K�|�=�Cq>�Z�=׳9<�v>�; <�[��*ː�!%!>L=�\�>JG9=[7J��n&��+?Q�9���� ��=��r�O�D�� >#�L>�V���^?w?�	�{�8��k�����U��ۍ?=O�?�%�?�����-h��'=?.�?�,?r��>�:����޾� �y+w��x�|p�+&>�%�>�~��徚���ƍ��U���P9ɽ�6����>.�.?��]?[�
?��
?��>�;5�	 !�_�P�A�T��U��׹E���Y��E�U�X�<sj�~Bּ��z�/^��dV��?!>�A���	?-�(?�(�>ֈ�>�ļ>b���+�ؽFj�=�<μ C=KT> py>��=���K.
�b>R?n����'�}��`���	B?f^d?0�>�{i�)p������y?��?�c�?�Ev>�Wh�?+��X?�=�>)���T
?m�;=�����<�2���������r��m�>_�׽�:�~
M��zf�Tt
?}?;鍼eX̾��׽敾��=D��?"f-?v����B��)w�S!@��Y�����pR#���Ҿ2�8�ކw�􎿩X���s��4#�$ql<g�)?l�?����, �������i�t�C�ri>���>iV�>b��>΂u>��@72�Y���vP|����>�q�?���>�G?#.?˨N?�??���>��>rB��v��>�=%k�>D+�>DD?�"? )?z�?�p*?�,>��ֽ�e��h ̾��?R?yU?���>�/�>w(|���z��3c�5���0p��9��͔M=��!<�9��
֣�3�/=�M]>�h?~N�-4���M�X>&2,?3��>7��>?Џ���@�f>="��>f,?}�>q3���JX����d��>���?tμ#�=�Y'>Vף=��ۼ�ϯ���=��Y�`}=��&<T�żH=(�=5��=�|<H� ;�'ٺ��=Ӕ`<�H�>	%?�>]��>�4N���B��}�>)E>=��=�\W>�p ����/횿	Gh�X>L�?���?@�-=�>b�>@ݶ�E�ھ�L��ľ��Z�16?�$?�(a?��?�I?�/?�& >�u	����R.|�z"��i!?-L?,��>�s��<���˗�-]7���?,6�>$�S��X�)�$ݐ�ܧo��>K�$�:� ���x1��A>��¼ ��?���?)�9��J(�ӎ�H���Ím�ݙ1?���>� �>5�?��߱?�3�9��%�>�b�>��?+��> ZJ?WKo?ߗ8?��z>��0�� ��Kn�ٽ�=�Sp>��m?��?�Vc?��4?�(�>��A���R<�����;����=霾g�k=���>}�l>��y>ٔg>!/��sP��5=�SD�Ya<57a����>C\�>+[>�\<���;�G?r��>�X��~�Τ�t���d+<��au?��?"�+?�=E�6�E�����P3�>Db�?֫?�*?�RS����=_ּ����pq�!I�>���>N�>1�=:G=.�>�I�>��>����N��:8��%M�T�?d+F?��=}�Ŀ~Tp�r|t������"<������b�µ���`�}�=ڱ��1����"�W��ס�a���#��2C�{�č�>���=���=���=�Z�<��弌��<�T=B�K<j)=��n��U�<)=6�d��]}���:���O<�.P=*
L�q�ƾlx|?>}F?�*?�A?$�t>�>�6I��B�>��t��?ҩT>���t���k<� ����X��m{۾��Ӿ�b��7����>+^�p
>�3>���=���<%��=��l=:6�=�3�O�=~��=[�=o��=��=�*>��>�6w?W�������4Q��Z罤�:?�8�>b{�=��ƾr@?��>>�2������zb��-?���?�T�?>�?5ti��d�>M���㎽�q�=O����=2>~��=r�2�T��>��J>���K��J����4�?��@��??�ዿТϿ4a/>uv~>��v>�_G��~Ҿhߕ��}Ҿ�pd��ʝ>'eJ�������=��=D 5���!�����!�>�k<�� [���=>��_��j���=�`s>!�<>�J=>�V���#-��&�>�Q6>� q>�Q�=����)����>��=69�>G�>+|�>�?P-?��`?���>Pul��˾]oľ���>h�=�6�>�2�=��R>��>!�3?�(C?AG?C�>��=:�>0v�>k*�cg���ؾ9���͘<At�?��?��>tx=
'����<��妽�a?+0*?Ì? �>PK�����.�DEW�n" �S�>�8>�H�=C�>o�|���������Q��<	>n>#��>�֝>��>@��>-�<�f�>��)>��Y�.��=΍>W���U!ҽ.�#=�u�=xp��1(�&[����
��}Q�{tT��m�=�>��ݼ�d˻�P>���>l?�>2�?� >��8��V=��D�ЮY�f��٢���F��4k��T{�/&)���Ǿ8I�>U�`>�{��g����>>RG>M|�>:�?Q�x?#8�>[:������$���S������ņ�5>�x`�W�G��@�-�X��>���>�f�>a��>�\v>R�2���J�:�y=�;뾃U6�w��>������<)3��*�Q��V���ܕ�J�j�b�7��~<?3�����>|]�?��??k�?ю�>�5�U��i!J>�����!=1�	��Y���Dc<�|?��?I�?*�վ��^�?�˾������>�G�?gO��|��y�0�F���K���L�>J۩��Ѿ�3��~��[��B��p�r��>�mO?`�?�$a��f���O����(?���2?%Dg?ql�>"�?{"?�*���*�E���ɹ=K�n?�v�?���?�u>+��<�P�W�?W35?dT�?E��?�U�?��>ܱ�?�[�����u����|-�%�=m��=&=?�8L?��?�$�� 8�B��E6�?�����<X�=���>��>ǹ>��l>��=�>�#�>�
?M��>�M�>\G�>YH]>P�����r?����� ?��9?��>�|>Uy�=&2�����$���D0ٽ��_�><[��o$�LΦ>����*Z>��ɿT�?��4>s�o���V?����9l�=o�>Z�������>O�=;��r>���=��=l��=L��>�_>O��e�+>�%���/��R��RU��+����=j���@�����wM��{���8)(�eJ(��=����þI�G=�W�?hX;�0Ux���#�0�<��>��>�x>?���Ie�<c
�=�$ ?���>_���&Z���v���X`�?E�?�6c>��>��W?��?w 1�¶2��~Z�Uzu�-5A�4#e���`�5񍿵����
�����x_?��x?�cA?�l�<�Az>���?:�%����r"�>/�);��<=1:�>����`���Ӿ��þ�p�	F>��o?��?<?��U��&�<wi>m�?fX/?�k=?e?]�2?�+�s��>�7>���>���>�{\?�,?�9�>���>�c>�@�TX=ba��{s����D��ĺ���ڽ�g�=Jl�<ʋ�&Kn=j�<O=�*��k�(�`J�<���������Gt=�C�=�L^=���>��\?���>.�>��4?t��F�Թ����,?T��<'�2�R�Y�}��u���%��=c�U?�?��Y?US>FAG��'?��><��>�3>9;�>�>KL�gȆ�	��<�>��=_�K=1S˽����[�����'���6�&>�`�>i��>�Հ<w�=7���d����=���߄��U,�;�,����3"3��|�>ָF?Ί�>�����ݢ�m�ٽ<PN��r?8��?}�C?n.k?-=r>�3߾9�,�P��勉�8�K>�_�#!�����-��s�_�/�e>Yɛ>������%�>[k��������k��Y�v��p:�h��>�?��(
�R���a�:>�a��$˾�9�����xO��ՑD?�|�=�Ѿ�;���T��2�N>S�>��>� "<�h#�ۼJ�=����U�=�?w�>!�S�dn���C�*L��E>�T:?�S?E�F?Zt��Hqq���,���4����+�a>�n�>��>�Z?��.>;9=��}
�q��NI�-�.�a?U��>c%�X\�	����$ξQ4�*��>~�>=%�>O�*?�*a?��?J�6?�?c�>\�>� 0>�վs�?��u?O�S�a]�ޑh�M3@�����w�>�ܵ>��+=y��=��>7?�)?�D?۩?o��<jz���I��"�>ڲ�>�p�!L���$Y>1�:?��?��I?`z?ǽ��d7��獾{�>���?=��>�R?~?�n�>�م>���>:�� ��Á ??۔?&��?�?�_�>�
{?G��5�>�=E��l�>��l>*��>�5F?E=�?���?��4?S1T=50B�����ې�����y�q��"=$�@��bS�s��<�7=(��=_�=Z���X|>��=��S��R��+�1�%��>��U>c,��W�=
��v��~'�=�/�<�掾7�7�^bY�Z�z>=(�>fh?�k�>����h��`�>1�>���T&?�^? N$?�3p=�?k�n�Ҿ�:��puI>�E?ͅ�=��[�����r~���L=�um?`/9?+{���⾁�a?�N]?�L��
>�̰ľ�i��M��TO?�o?�,>�/��>+6~?cXp?�]�>!L[���k������a�>v�[m�=
��>����d���>��8?z��>�;i>z��=��ݾK	x��A��˰
?鵌?J��?CӉ?-,,>^m���߿��޾�p��]f]?�s�>*ϛ�*f?ro���ڱ�mj��3��]Ѿ����1���u{�n?��&�I��̋�k᪽/j�=NC?��m?�8�?�e?J%��>Y��(_��8����^��R�e'��K���=�*IN��"y��f�Uw¾_ݫ�F�Ѽ��[��GC���?�e?�;L����>�2z���ʾL����H�=Q��1x���G=�,��>�=Q��<�A���ͽ����d?�>�`�>��3?��c���@��5G�X�G��/��bd#>���>;q�>��>K��ֺ?�f0w�Ǻ������z���l�>KC`?M@X?�y?V�җ��X��!���=���dݾa��>N��0~�=ɚD�A�x�A��i�;�G������K��m���=D4?��>.h�>D��?J&�>�0ھ���1B���Z�!W��J�>1[C?�v,>yߧ>�i��� �E��>�l?���>�֮>
�����\����ͽXG�>�f�>��?I��>�_$��Y�񰇿��N�)��C>��Z?���{o_���t>XoQ?��=�:=}9�>莠�@���/����?�5%�<�,�>H>^Q1>��;���<���Њ�)$)?�R?��þ̘'�\�>��?�?�F�>���?l��>S@���n1=�?��G?[aT?gZ?�	�>ě��f�G�?Mٽ���R�=#�>�C%>�~=�#=�L̽���ݝG�O �=�)'>����,/���Q�<�󹒚�;��a=�>Z�ٿ�uG�w|־*����i��\��$��'쓾�=q=@Fľ>����X8��-@�R�&=>bG�����8|��W1H�v��?��@��=�ѫ�=M��W!���^��&S>���>�����R�(�
�4�ep��)SL���Y�Z��>쓿ߓ'?y���y�ǿ���IAܾ ?�? ?��y?��O�"�2�8��� >���<�М�S��_���Y�ο����\�^?��>=��8�����>���>!�X>�Fq>����ើ��<��?q�-?0��>Ҏr�ړɿ����<���?��@<&>?g�Bھ�;j=���>�F?�a%>�K����Wq���R�>�,�?iU�?$�H=��Y��%����`?���;z4��<��=�l=�y=w�|�:>Iہ>�����>f����>�Γ>�W��)J�!?�꘧=ٞ�=�{��An�=	Մ?�y\��f���/��T���R>��T?�)�>�>�=��,?98H��|Ͽ��\��)a?�0�?���?��(?Zݿ�֚>��ܾ��M?�C6?��>e&�h�t�[��=h3������㾀&V����=ҧ�>&�>�,�x��@�O�a4�����=�g�_�ʿ�70�TM �KAx;�r-<���&	�7�g���)�^)���P�mj;��>C�>=�m>��v>0�u>h�>�*a?΀?�Q�>���=xd�����ľ��+��Z���l軪Ƀ��Q��t��U*޾ �ξ����Œ�6>�|x��8�7�
��=�TL�<���&�t�e��K���-?��>l���O���<Pvž���A{�3����־��4�d�l��ܝ?.l;?�����W�Y��uႼ}����u]?R������믾���=��4<�T�=��>U��=�Dھ��%�O�O=?��?3�վ����-�>iGM��׊=�G'?�?�I��k��>a�?s<�jU����>�6>`����~�>r��>�m��H>��QO?3�a?&͐�)-���/>�弾��N��$½ ��<P�����>KG�>M�@�קȾ��B>��x<�r���R?���>�,� � ��M�o�r��pB>��h?u��>��?���?Y�_?��(�*��$���p�D'��qT?(��?��>uee�M쾰� ���?T�n?�s�>���cʾxEH�V�'�˼�>,]�>$��>�Յ=�;y�����qw���#?��v?�s^�Ws��$��@�V��A�>�]�>���>��9��i�>��>?##��F��J���	Z4�Þ?|�@=��?g;<<�����=);?i[�>ӬO�<ƾ�u�����=�q=G$�>Ƌ��-cv�B��V,��8?���?d��>�������e�N>�V\����?�Di?�p%p=�.�	J�dI�R�3��G�>;�E>S�.���N���}��#���ږ�;����.�>y�@)o�]��>0�����m���������m3N?��?�է=6�!�N�}���5�a&���7������h�>2�T>e�j��E����t�Z#8�
GA��f?I����Q>�Y����������=�GI>��I>�r�=��2�"���"��?�z־�ʿq�����xCI??��?��?�)+?D1ҽ�搾��q��z�=ɨY?gv?��D?����j����r�o�i?�����iU�C�7���3���b>[�%?ڈ�>؟%�U�=P ?>�j?0n�=�7������"�� ����?qa�?���#�>墜?z2*?nX�GF��O^Ѿ��0�HT�x5?��>�]ž�^�-�)�7z��6�>xqI?b$��==�[�_?�a�K�p���-�f�ƽ�ۡ>�0��e\��M��,���Xe�
��Ay����?J^�?e�?��� #�c6%?�>`����8Ǿm�<���>�(�>	*N>�H_���u>����:��h	>���?�~�?Qj?���� ����U>�}?�>Ƅ�? ��=���>{�=�	���M�p�>9F�=�?%�ki?C�M?�>�>���=�b6���-�Q;F��
R�j8���C�z�>�gb?1zM?*�c>Zs���3��!���Խ��2���7�C��N/���\�0>��=>��>��G�ǍѾ��?Jp�5�ؿ�i��p'��54?-��>�?��q�t�����;_?Bz�>�6��+���%���B�`��?�G�?:�?��׾�Q̼�>5�>�I�>��Խ����[�����7>+�B?^��D��n�o�l�>���?
�@�ծ?qi��	?���P��Ra~����7�i��=��7?�0��z>���>��=�nv�޻��Y�s����>�B�?�{�?��> �l?��o�O�B���1=;M�>Μk?�s?UOo���k�B>��?"������L��f?�
@~u@a�^?) ��������=�ˏ>|M�=>�|>e�`=vr�=�~��A����<<?�>��>��=,��>{�S>�
p>��>�����G*�뎦��n���69�#���׿��@���V����4�h�ʾ�S���w����d�.�5�?M
��+0��>(@?Ӻ$?'�\?ܹ�>�c�UK�=-/'��G���X=����=��'?j�D?\?
P�=y���O��dm���|��@�+c�>8t�=��>Eg�>�In>��g�>�>N4�>4Q}>�9�=�}>L}�=|2ػA6�=��>��?���>�Y,><{>�#���겿�Y~�����H��ѥ?ݘ����8�������m��O_��C\>m�?)�߼}㏿ʎǿJ���d�;?u!���t��t�v��=� G?(�Y?',U>�h�
J׽W�f>q����i�ˊ�=����e��#��/�s>�?hJ�>�5�>��2�0o7��R����D�>�3?Wq��xf<  t��G�������>��>/��=�\�UY���?��'R����8<M�+?H�/?�ű��EȾ��X<Ѿ�{�=�dh>�`	>��=�o|>�����p��޸�:=�@�=2f�>�� ?��>T�6=��>O���{'a��$X> n�LL)���L?a?�>�΄����;��,�A���d;�=��>��=@���P�d=B�>�>�<=����)J=�\L���<�8]=i�����~��=�1���<Ob�<��<�5���[I>�~?���'䈿��[e���lD?M+?� �=��F<��"�D ���H��F�?q�@m�?��	��V�:�?�@�?��8��=}�>׫>�ξ	�L��?��Ž,Ǣ�Ô	�)#�jS�?��?��/�Wʋ�2l�~6>�^%?�Ӿ�;�>�N�-G��U$��[v�l�=�=�>�cH?(1��J�O�0K?�se
?�??]i�������ȿn{v�VP�>6��?�ڔ?
�m�&<��F @��.�>��?TmY?c�i>v�ھ��Z�2�>h�@?R?��>C���&�?�ȶ?��?DSB>wd�?<?fE�>����51���=���Go<O\r�YB�>h�1>h��.@Q�C���}��Y�>���A+>�y=�>rn����+��=��۽�䠾Κ�E�>��>��>�Bx>`~?L��>x��>,D�=�9�T�b�M����`E?~�?�X���m����"jO��Vƽ(��>0?Q�=����n�>�%F?�*~?�m?>U�>�J�8���Xſ�����W�;��C>�? �>�����>������X�̅�>��>��żn���}��s����Y�>w� ?h�>=��=,"?�2?lv�>�|�>bo ��Y\��G����>|�>�9�>pP�?���>�B�K�8��Y��q���;��)>��^?l&?n�>�����p��%琽*C��������?�NO?9[�<��?"o~?�?l�=?�[�>^$P>M�,��s񽋭�>��+?��#>ϢW���*�{"&�`l�>�O?a��>�=U=N׽�rs���ܾ�6뾂*�>��t?b|O?_<˾cb��
 ��_&=�cɼ<���oۼ����a>�Ib>�Wk�R�>�r��0Y��Ľ>ъ�
�C<md5>lFZ>��m=`�K��p��*=,?��G�Eۃ���=x�r�+xD�p�>�IL>��t�^?Sl=���{�����x��O	U�� �?��?Fk�?���8�h��$=?�?g	?o"�>�J��~޾f��CQw�~x�uw���>���>��l���B��������F����Ž&��:,��>��)?�lL?�?
�>JJ�<����()���)���=g��7�)Tu�فQ��-G���Q=2�,��M�<�h��a�M��ˡ>2�=Q?.�+?�.?��>2�>�?x�8t�=A�Z>�5�<Ǥ>���=xS>M_�>.�>�<z<mL?SG����(�������¾�D7?��Y?��>7�&�|}����e'?���?'}�?zq>^�e�9�,�D4�>�>z�~��?�Y=$�<6=�j���r���ý�L��I�>�����,�4nO���x�!
?�s?F#>��;Ǿo{��?nվ��=kp?���>�U�;�j�b׃��r�-�|��T>>�Iƾ��#�����n��������������f�E۩�X":?��^?�8߾�[��&����u��E�6��>z�>]�Z>�s>�z�>}���y�d�A�Hb�s����N>{*e?�v�>(�4?]�0?�T?E�&?��E>�Ȟ>X'�z�>��p�� �>iK�>�)?��?}?5�?y�?n>A�n�B�����Y?�R!?�,?���>A�>�����Y"�a�E�X��������㽨�Q>�^	�I��yL� �>�q>�[?�d ��19��.�UG5>��*?_>�>1&�>�⇾l�7�)��=�P�>z��>dEo>h�̾E�e��6"���>�̈? �ۼ�l�;�9N>�d5=1��<���<�"��p��/Ĕ=�ߘ��Jý͔=^�=,�H=g4��<�L��p=̝=y1:���>��?�<�>D[�>.#������X���ԧ=k�R>��8>��'>��پ�	��Y��,g���S>i�?�b�?�'l=��>��>{����ľp��-���=5�?d�!?�.R?���?X�>?]�?��>���g����l��T+��-�?�?CZ�>J$���ݾW���99��5�>�?xN�������%���Y�o˅���:>?��>Xk������=�	�
;'��Ҝ��I�?3��?r,<S]?�h�J)���⾍lD?S�>���>9�>��:�8�[�C-����=ە�>��@?���>S�Q?��j?�Y\?�} >�!�妿�)���H����>�`d?1�~?p.?�6?ڀ�>\>i�	�net���Ӿ��7��Wk��>��2�[=6U<>k�>$��>���>c�E=��a���<����c ��h�>'M�>��G>ԣ�>��>n��<�G?l�>����{�e��Vg����;�1iu?�S�?d�*?*�=4/��F�vW���C�>�>�?P��?	�)?��S��f�=c�Ӽu����r�;L�>-v�>��>w=��N=��>���>Z��>����{�7�I[D��?k�E?���=�Ŀ?6n� Lg�������;N ����i��5���,f�4�=������C|���x]�͗���ǖ�uո�W���d��a��>ڌ=_W�=A6�=z��<��Ѽq֩<�Z>=o�o<�R=C�{�tt<�1�H��)������S4<y�+=m{.��Xƾk|?mH?��)?�xA?�Yq>Ę>e0��J�>I�z��_?{�Q>/7J�T0��4�3��槾���P�پ]vؾ��`�I����	>�c�w�>2�3>�T�= \�<�>�&r=�i�=��	<s�=���=�e�=�p�=Í�=�%>1)>�6w?L���	����4Q�gZ罣�:?�8�>�{�=�ƾX@?��>>�2����ob��-?}��?�T�?4�?;ti��d�>D��䎽.q�=Է���=2>���=t�2�d��>��J>����J�����4�?��@��??�ዿȢϿLa/>1G>>:�>�?K��/A��������J�s�1?��C���+�>R'>E���+�"�NA�<YL�=��;
#Q���L����=�� ��9��<A_�>y�A>aћ=�Tʽj*(>�>1�H>���>+6��0�&�F%��]�>��=fg}>�f^>���>�1?s�'?��X?�y�>j�U��_Ҿ+�ξ� H>(�Q>��>�	>>A>>q>��?ƥ5?d�6??f�>D�=>���>D$�>V�-�;�U��|�c���D�j=�1�?��|?�1�>�>�R���W��j6���'<�?s��>Vz?k_�>��Ut ��:�k�\�ʽWǿ=��D>����ݴ����������|�>:�?l�>�J>��.>��Z>.�>�
�>��B>=ڮ=�>,�潁Q��k��i��L�m=��>H}�Ԗ�=�2=0N��"�>j����ٽ���J�<s��=��>��M>H��>��}=������=�x��ClI��>a=b�����A�R_�g�w�j,��:`���,>�&.>;��r����M�>ښ�>yqt>�9�?�7z?�P>>�f ��оˍ��( ������Xr=�~z=�nl�$�5�S�D���J�@�оR�>�2�>�Q�>W�>vN�����􍽾TҾ\/�k
t>���,���W�ㅿ����ǒ���P�bŀ�'"?�y���>LD�?Yk?x��?܏ ?G��<���|�;͜���$%����5��ƾƏx>i?}N?�1羑$���˾�`��ĸ>c%G���O��e����0���#��Ϸ�{&�>4&��w
Ѿ��3�����=쏿�'C�ap�w��>�fO?yҮ?�`�~K��j�O��=�����~�?fvg?�9�>�'?�I?�Ǟ���/��0*�=_�n?�d�?O��?ά
>�4|=�Eվ�?��[?Ls�?۲?y��?K��>�%|?�l߾{�B<�$��ټx=޽�ҽ��>!�\?Kci??~�9�q�4�]��L1�45��ğ<�N=>[�>��	?H��>�>t|�=�Z^=I�>�M�>hD>���>�e�>A]�=�ed��� r6?d>��>�0?�p�>�+>Z�g<<J���k��u����4彘�ӽ���a�x=2V{�uV>�-���>&�ƿ���?�f^>7"1��)?�<���>H��>�&�=K�нh��>'�r>�h>���>�,�>�?�=���>�Oh>,�Ҿ�h>�g�Y�!��(D��'S�ReӾ�|>n����#���	������E�� ��Ǌ���j�rJ����=���<U�?���:�k�,*�-����&	?�Ѫ>K�6?w���E��՗>���>e��>�h��׸��^���R߾��?��?��c>��>*�X?'s?�m.��7.��Z��t���@���e���^�廍��:��y
�P�Ž��[?j}y?��@?�7�<CA|>�{�?�&����,І>�o.��P9�>�G=�f�>���2]��dо��ž��$3C>-�o?̧�?�}?,<U�	Vj��}(> &:?P�1?�rs?l�0?:�:?�0��#?��4>q�?��
?!5?�.?i�
?��1>�=�����"=H]���/��D�ҽών.0���5=c}=�WN�1�<~?*=�ò<a�ڼʼ�;�L��\�<L9=�!�=���=���>:2]?�S�>ދ�>�<6?�����8�*���+?�M2=u�{��y��X�����D��=8�f?,�?&=X?	�_>qKB��A���>�ۊ>��*>H_>E�>.�7�F�ׇ=��>�7>�=�Q�ʳ��ur	���t��<Y�">'��>tz�>q���(�S>S,���򖾳�S>�\-�dD�� ew���0��ѾJ�:���>��-?�<$?�e�:�V���+��.a����>;Qu?�&x?�a_?�%=�	���d� ���9�>"�>h;ٽZb��k響
�����6��%�=��>�ܠ�1���p
�>I��z5�HKx��[��iM�Ǿ��N��F?����롾�`�<t3�>]��;�����.\����}6��C�>?~&6=���ׁ�������%>��>/A�>���=��<Tc.�����|�=ߓ>(K�>��>�]پ[�5��;q>�P=?�FM?+-??�%����p�HOA�B5Ѿ뱑� �=Q�>>v�=��?�Ӷ>� �J����TR�qJG��>K��>?���{<��̽V�������N��{>>G�>�Y�>�m?zE#?1�?���>|�>`�>���,���'?(�~?He�<�H��}e�nl.���;�)ã>��?�D���>	?��%?%&?^�-?�)�>V�=JP���+��>�2l>gW�E+����=	zT?P�?��7?c�y?�D->�=-����3����=YTv>�SA?L?X��>)c�>Pב>K�(���g�> ��?k��?�?��T?H��?VӼUmS?��>@��=���>��h?U}?/��?���?�}?Wv�;�)��=�wH�I�<Mv�XE/=Lh�=QH߽�;������u�V�ڻ��|���Ҽg2���4+���0��X�<]?�>��t>����C?>�Lž�����6>����hj������W-,�Cҩ=L��>��?|	�>����t=�a�>�¾>��b�(?�E?�?��k�e^_��ؾU�@��ˮ>c�8?��=Akj��ؐ��+u��J=R�h?�Bb?g�o��;��J'd?�[?�
����<���ǾfjQ�'�Ͼ7�1?�?�b��W�>�tt?`�s?�K? �h�E{X�����aH^��`Q����=�c�>e��eOl��]>��A?a?��v>�A>��߾��k�<���.?|u�?�?5�?&��=�}i�<�տ�A������]?h{�>4���m�"?,�*�Ͼ�z������_v�m��)ȫ�6ꕾ���p[$�Y���k^ս�8�=G�?�s?��q?"�_?�� �B�c��U^������V�g����&{E���D�H�C��n���7��Bh���G=3����-�XQ�?�v?��8�M��>=z��tL��Wؾ
�.>���y��7��=i����M9;k\;��g�ͨD���Ǿ��!?D��>�»>֊7?u_���K�ӗ2�1�:����:�>*j�>���>���>J	<�)�yb �R��3��!� �8�>\$^?Y�S?h�q?![��X�#I����'�a�(\��xXD>��>X�>^���d�Y�hh'�-�Ll^�%���I'��V��'�=G�6?Lӟ>�˲>�.�?O9?�_�vH˾zp��g�;�ց��ۯ>�^a?���>Я{>�㰽]���+�>ǖj?ϸ ?��?2Խs¾�/\R��2<>���=��?��>Y11�����&��+���o�%f9>�Zw?A�����]���>f�Y?Fyy=�$>�Ӓ>w<�_G���ѾJۋ��� C?bdb=�=$���ˬ���M�Ng���6?�?�Aվ�>2�zZ�=��?�0?�#'>:`w?��>���A=~�?�&??�|V?�V?��k>x���%��n��.*�,N�=��>s�I>~ Լ�s=�_���-��ܽv�S�	>�ų�j�b���=�Ju�y���=r��>8���M�N�x�>/�Qn���t�Jxe���޾��a���Ҿ�n��ޠ���8�C���KbؽPÔ��(��^����?�1�?|̊=0��E��ž��p�9�`}=�˸�{->Ό}�Vc=����jڨ��\���	%�,���i���iN��Z�'?3���ڽǿװ���:ܾ! ?�A ?�y?���"�s�8�� >;A�<�/��c�뾀�����ο9�����^?G��>��-�����>���>��X>�Gq>����螾�0�<r�?E�-?S��>��r�/�ɿ_���kŤ<���?#�@��/?��.������#{=�8*??�ʺ�8�� �����E��>���?*?q��XJD��\=��m?O=>y}$�^�%Xu>�7�=nؔ<��*����>���=�}��G�����	�ڄ>}'x>�U��o8���y�	���'@>�����Q�3Մ?�z\��f���/��T��U>��T?�*�>�:�=��,?A7H�A}Ͽ��\��*a?�0�?��?��(?Kۿ��ؚ>��ܾi�M?]D6? ��>�d&�#�t�w��=@7ἁ���B���&V����=\��>��>��,�����O�H�����==|��uۿ�8>�:1����;�$4��}���ĽI�E���Z��~��qU��^푾;���]D>�D�>	P�>3K�>��>:nO?w�W?s��>G��Nrh�0h���ʾd%��j����I(>�>� �V�2��e������9��]�' ��aM�o�1��=}�N��~���-�l�a� �>��E
?�x�=<.B��u���z�����]�<���RIe�S1�I�S�5�m�V�?q/9?�����b�#:�LX�=�����\?@�H�[��jg�l��= �Pkj<�A�>'��<�>���D���V��9?��?_l۾�i���ܖ=Bw��!>�]�>���>�� > 7�>@%?˳����&��֦>J�>���=��>�`}>u����u���*?��_?�ɒ=�w��'�i<˲���F�� q= :>E?��>�2����?r��=�k<��1=W?r]�>��)�\��L���Bg�^8=�x??kǟ>��k?��B?�J�<Uz󾐏S�S�
��w=P�W?Œh?,�>�~��uо߮���'5?9�d?4�O>�i���.�/��ɐ?��m?xk?p��Y�|�풿)��5M6?��t?�_����La��7H����>���>W6�>�5�J�>&t??.���n��E���;0�V��?3�@���?W�<._� �=�n�>0��>؈L�N�¾�����ӵ���=M �>gc���,q�}��%�C;:?΅�?_?�~�#���@)>��q����?��d?р��m>�G��rf�󗰾���0�S>���>��.>?�#�{�+��7��F[�� ��^��Ly�>�@h�I�I�>����~׿q5׿L&��%����<���>�!�=�-Q=����[���n��	S��c;��~�-�z>,�2>�i���M���4y��7O�K½��5>3d���"?a�Ӿ�����a�^BP>B��=���>�y�����̺��H�?�˾��ɿ�x����m"o?��?!wr?b�;?���<���0�ξQ}���UW?�|?`�P?7�=O!��}�����j?�]��jT`���4��GE�U>�!3?iA�>`�-���|=�>���>;e>}$/���Ŀeٶ������?ŉ�?�o�@��>ށ�?`t+?�h�V7��D]����*�C/�<A?+2>����˸!��0=��Ԓ���
?�~0?�x�|-�Y�_?+�a�S�p���-�a�ƽ�ۡ>��0��e\��L�����Xe����@y����?L^�?k�?���� #�l6%?�>b����8Ǿ��<���>�(�>�)N>H_���u>����:��h	>���?�~�?Qj?���������U>�}?Ƿ�>�݀?���=M�>��=NK���9�����=���=�׿�4,?��J?4\�>I�=iF��� ���=�oKI������IB�C�u>��g?k�P?HI�>��3V���?��~��k�n���<'�I�߅��I���|>t>N>��B��9ﾻ�?�s���ؿ�e���P'��94?���>�?���@�t�G��6_?jp�>�8�B)��"���-���?�G�?b�?��׾M�̼��>��>�K�>I�Խ���������7>��B?\���:��`�o��&�> �?E�@n֮?�i����>\������3�]�6��6��G<>��M?���G�>u�?�h >w�d�5����]���>�b�?���?��?w/T?��d�eRC���(;�U~>�g?l�?��(��z�j>R�)?��i���R�����%9�?^@�@\i?-)��h�޿����c۾=�̾���=��=�h>�������5ѽ�;����<d��=�8�>�J�>�Լ>D�>u~>�Z>�܌�%>,��j���a����5��V�]Q��V}��M.����Z�Pvھ���>���"=A��<U����U���J=H��=B<9?XLS?�C?��>������u<���U�c==����J=G����r4?I�G?�<?�*������jD�ۖ|�թO�?�ÂT>O�>�[�>�d�>_BG>$nD;E��=��>y��>
Sü�$D=~! =ˑ�5�=x�D>\$?���>�|8>2h>%��.���Si���}��׽TO�?�����B�����%��z;��_��=2�*?D*>Fx���п|����#G?�b�������2�t�>��-?�KU?'�->����A�o��K>b��\lm���=c�罭�l�}H&�JZ>Gw?M�0>�O�>u��f�q��Jq�^�lֽ>@��>'龀��>�M����,�Ⱦz �>7�>X%��U��㗿�����|�+M�=�M:?��?;F��O��1>@���� u>[m�=%{�=B�=�k�<ۈ��X<<��ɾ�Ed>jA�>�XM�n��>u�A>��>^��>�-��`�p�T�;>g�=J��=$�?<>?[.S�H#���I=��!�5*>f[M>�/>�J���k����=�H ?Q��>mw"=
K� Xw�Z��>�N>�9u�N ��!�μF	�=%���OZ�=#ذ=4ѯ�������m<�~?���(䈿��e���lD?R+?^ �="�F<��"�E ���H��F�?r�@m�?��	��V�@�?�@�?��N��=}�>	׫>�ξ�L��?��Ž5Ǣ�ɔ	�*)#�iS�?��?��/�Zʋ�<l��6>�^%?��Ӿ�g�>�{�XZ�������u���#=���>m9H?;Q����O��>��u
??�`򾌩����ȿ�zv�a��>S�?���?;�m�XA���@�~�>J��?ogY?Bki>�h۾"ZZ�Ǐ�>z�@?u
R?@�>>7���'���?�޶?��?�:>�-�?N�{?hT�>�Ǽ�ӱ0�A�u��'��;*P=�k�>0�	>���� F=�'J������/^����w�.><3P=���>,����&���6�=Avýb̞��3��B�>��>t8>�B�>G�?Tż>,wz>3c=-�G��H|��Λ��4K?Z�?��JBn�-�<1��==LY��J?�T3?�(�RuѾ�.�>�L\?�Q�?S[?�P�>q�����[�������K�< �M>$.�>C#�>n����F>Xվp�@��>�;�>��&/ؾ/���ѯ	�ޗ�>�� ?��>bĥ=E�(?�,?d�C>�c�>���c�n��G9����>���>� �>�%r?���>��)^�/ɒ��;��S�0�7��>'1U?�6?��>@�������p�p�~��'>��\?�7?��#��
,?l�l?��>��~?�q�>�������En��I�">�j+?+yC>�OF��������Ȋ>P�D??�>�8B��Ɋ����=�D+�#���/?L�??e$?���"�">���==���<�I���M��^=�&y�>_��=M*��/�P>���=��Q��|����̽�.A�D|>o�>*��=8�F�==,?a�G�Uۃ���=��r�xD���>IL>2��~�^?l=��{����sx��B	U�� �?��?k�?���8�h��$=?�?�	?�"�>zK���~޾���wPw�6x�w���>���>��l��*��������F��G�Ž=�����>�#?'0\?��)?�6�>Ic)>ϔ� �,�TL0�{�Ҿ�_D�G�վ��P��a�'�\����ۇ<o�=桱�S����
>��N���>i��>���>�y�>A=�>-輽ř�=���<�7ʽ�}�>��V>Z >>-�=��=~�>�JR?	�����'�-������)B?�id?%:�>�i�������wv??w�?�q�?E6v>�uh�;%+��m?3�>���6n
?��9=I~��w�<QQ����F;���7�J��>��ֽ�:�<M��5f�<m
?.?����߄̾�Q׽������i=`��?�?��-�x X��`s�#]���Y��um��u����60%�zXi�L��t��2����m.�I5<�v0?���?�t����޾�i��j�v��l@��_E>p'�>�ɩ><�>g�n>�����$��
Y� � ������>��c?y}�>ӈB?�;=?��P?E�9?�gy>b˃>0����>����v�>*W�>A�3?�e?��(?�?e ?F�A>�3	��&���оG�?��?R.!?�*�> �>�?@��n+�f(���oS�r��m����r�=�d�<s��J��;���D�>y�?6��)�5�g���\>��.?k�>Փ�>����Q�e��n<���>��?�ę>�羼�h�Q����>ynz?���c�<'v*>�d�=����x%�;aק=b%x�KB�=QM��M��ꩌ<�=*�=)4'�[S�<�[����<�J=�S?�x?�3�>��> �=Z��R��Y�+>d�>q�>A�>��Ͼ��#唿1l���6�=NG�?-�?`-�=�7>i-$>����b��*�U�ھ ��<7��>�	-?�Z?nR�?d�.?1�>�>o �V���),u�����.�	?@�?xԶ>��ľ�(龳����).�m�>}t�>�Ja��r�_�(�v����Y��%�#>.�m��UA��tqF�]��"��8Ie�$��?��?���<}$���־����PϾU?�1?���>s��>�$�-�w��T;�s�}>�?2�G?ut�>$�L?�*u?�E?暒>C��&[¿t����\���=}�*?��?v��??
'?v\ >�|�=���l�a�H�h�;�ʽP
����=��>~�>�F�>�>oQ��hѐ���]��]H��ϼbQ_>���>��>c�p>+K�=�~C=�G?,�>���p�\����]��:�:��u?��?`+?"�=mb�%�E����q�>]�?��?�8*?'�R���=��׼������q�ݷ>y��>��>A��=�C=l�>F��>���>�=�Jg��k8��UM���?]F?�|�=ێ¿?�l��h�w��j��;�v����b��>��J7^��T�=�o��Bj��V���O�A-�����I���5����䀾���>T^l=�p�=Q�=h�<�ɼN��<|WX=��T<ܱ=���e�<�GJ����+�u�V8�;`Ԟ;E�b=�����ƾ�.y?]�J?�h?u,?l�$>d>޺	�>q��#;?&>9������J�J���?��׆ؾ�����Y�>����E�=8K��v�=��%>R{>���<��<$1~=A;>�Q˼i*<��==�=3So<�2$>�0�=��>�5w?��������O3Q�M��:?/:�>���=D{ƾ�@?��>>h1������oa��.?���?+U�?��?�hi��c�>���c⎽bp�=c����:2>��=��2�[��>��J>H��?K���|��Z4�?.�@��??�ዿ0�Ͽ	a/>��T>w)'>LD���%�@�f�Amx��04�Q$?�Z3��ͮ�R��>TJ.=w.�\����9�=�>C��q4��fT��[�=�{�$��BMU=�S}>�?>m��=������=���<`��=Q5>>��ۼ�4� x�;П�=n�V=�N>k�.>�E�>��?��/?��i?�O�>�?��wѾ�����s>*,^=��>��=�� >C��>�9?�/?|"E?��>���=OM�>�Y�>�/��Cn��������:Z��?��?�c�>kx�;��9���"��9���޽�?�)?��?�>v�ɛ���aO���T��]��e��<误=lf�ͽ<�ɽ-I:�4&v�b���>b�?$Ϯ>އw>7�g>;ז>�x�>�A^>$��=?�=^�ݽ�ɛ�{_�<<6�<oy=�PC��i��kg;4�>P��=�CH������ۺ=9ױ�?�P�
q	>��>«;>��>[�
>���}�=D�}���G�]|<�Y���6��
J�,����6��9W�:D>0�]>8�ob��%q�>V�_>��>ߢ�?<�r?�hb>}1y��ؾV�����f�bE����<��=,KU�HK�@�I�>�>����q[�>0I�>aЯ>&�>�P"���4�Ȓ2=��ᾐ�0���>�򄾐��"��c�t��������a��<�;�YC?}r����=p z?2L?=ԑ?9�>'\�S�þ C>�?��K�;���e{�� a���e?�;"?�2�>:|߾r�C���˾�E��*��>�F�!O��L��,�0�t����෾�w�>z����о'-3�c���%����B���p��>�>LyO?�î?�a��R����O��#������?�Fg?9�>ah?�?�ġ�����{��D�=V�n?`�?f��?v>'(�=%Cվ���=��E?��?�ǣ?�O?@��>T�V?�A�Lٯ=�&=^D����nA���h>r_.?��H?_?�z�&~.�u,:�!�6��(��F�=��o=� z>�*�>7�>�:�>ᙕ>_�1>p�>n��>?8�>a�>�?Uo�>G�E���
�!;5?�:>�H�>�	#?�c>�D=/V�=����;3����p̽Fh���o��<��w=!��=�cּ�Ԕ>��ܿ�F�?�Y>QD��^=?S�����>eM�>�]����Ԃ�>�ip>h��>��s>8��>�[�>���>[4>e�Ҿ�T>+���!��B��sR�m^ҾΕy>�p����$�}Z��G����G�匴�ra��j����l=�6L�<r5�?�����k�=�)�R���s�?��>!>5?`錾Ɂ��/B>ݞ�>�Í>-3��z�� ����D���?f��?Gd>�>kX?k�?��&��*��Y�ar�
@�f�1�_�gf���F��f���`ѽ��\?�w? A?N1�<w�x>]�}?�t'����40�>_.��:��ve=��>�԰�G�d�WҾq�Ǿ6e��1D>[o?�(�?�s?7�O�
7�&;->��9?��2?>�i?��(?p1?�!򽔀#?%>��?��>�,?�+0?�T?o+.>�	�=XQK����<�7���Ä�+J�-ܽY�^�Y	�<�;=�Q�<�H�<��A=�i<�j��[!����<�-�;}�:=�:�=�!�=� �>)�\?�L�>�Z�>�G7?9��w�:������+?�� =����G����!��˘�=�h?%G�?�wX?g�\>"#C�H�F��r>#	�>T�*>�d>v�>��ܽ˖L��p=mr>��>:��=-�d�1:��d�
��Ő��M�<)�+>i��>�_�>�_̽�(>0!���P��C�>��t�;���n�T�	������V��x�>��?��>,ə;�ľ2@��>$W�#)�>�/c?'�?Ǡj?ru�=:�1��O-�8�t���5s�>���=�w���/��6d��3�<�O�9>�s�>6����`<�%v�>y?_� \@��퇿��F�X
���'k�g�p��F?l1+���q�,N���>�X=t����-��֠�@֢�7�<?-i�=�짾��Ӿ��ƾ�BR>���>��>[伆6<��3�a�ɾ��=>Q��>LV�>{>>ڛѾ��6���$>W@?��V?{�V?竓�1�m��N�n� �����#�=|K?�X�>|?�[>8�<������U�W�9�S�>���>;r�a�/�6�ɾ�d�VQ�+ �=R�h>N �>#�?u
1?j,?��,?k�?i��>ES�> �#�������#?ݍ�?M��;��~���'�Q$�Z7�a�>�r�>��۽.��>��>�+�>�#?�F8? i?ùR=u� �������>�o�>��l�ە���i>�s:?x��>�X?^��?�ll�i]�o�J��Xֽ�	>O�>�+B?��p>h��>qV>�5�>D�X�?&�H��>�F�?��?N�i?�K?�3h?s�_�?�>�B�=�3�>��??-8?}?S��?�ښ?�� ?�;*�F�?�=�e��@A�{��vs��{�F���t��BU>��t�=�(=�<<���;gg��Μ"�gzýS~��l�>�U>��o��o>� ���⫾��.> ۼ�HI�c���or��U>֏�>x��>�۲>��@�w=H`�>Py�>7��Y�?:8?�U?�%>��K�
�Ӿ~_�Ί�>��&?d�%>�~\�q䒿%�b�v
>�}?�Nb?��4���%���b?}�]?�����<��þDUc��D�%_O?�
?ȬE��ڲ>�N~?�q?���>Dc��#m�����i�a��#j���={ߛ>F?���d�$��>�"7?k��>��d>��=?�ܾ~�v�B����m?+ƌ?��?��?'>"n�:�߿~����㏿��]?�k�>B��sR!?� R�X�;�����3����ݾ�g��PԮ�?"�������!��B��D�׽:f�=�?pp?<�r?�a?B���.`��^������U���{-F� �A�*E���p����n��]Ք��`C=>Z�e�G��.�?[�(?�>���>����8n��h�:�.A�<�B�Be��<�0>��/>�Y>x��=y?o�9�I<�J��x*?��3?��>��!?�b��+��O�N��F��N;�,��>t;�>�R> �>q鈾���m�����
���;�8�2�>��[?Q�>?(E�?M�=���5����ξ��;\�㾿�>c��V�>D�������k�����>�B��E\���x��n�o^-?���>u�?'�?M`&?�������"��`�Y�e���А>7�B?~��>�q�>�bj���&��>�2l?��>-Ǥ>ъ���ό{���ҽ��>.�>��>Pc>Cb0��r\�<��y���]/8���=-Pg?k߄�``�6��>-�R?S�;�8R<���>�z�> ���ک)�b�>b?�/�=��5>K�ž��	�j�y�v����[$?��?0���2���J>�g?z?���>��\?��>�W̾�
��p?W�=?4�Q?\7?�J�>�RX��!�b\������:��>l�3>�ܕ=�bI=��3���qV���=��=�0�gQս��=�"�T#�;u�<�,L>9�῞&I��ʾ�!7����fc��/�������}�i��.�ھ�K�򀑾𡓾O�0��K۽���C�1�T�+Z�?J@�`?>�)���̜��Ǉ�=ÿ���>����E�>�L�Īp���Ӿ��򽨜��þ�l�x^������'?ݍ��ĭǿv���CGܾ ?I ?ky?����p"�Ig8��!>uF�<����r������οQ}���_?B��>d�+���9��>4��>�&Y>L�q>����؞�!�<F�?�n-?�S�>J�r�Ɋɿ�������<r��?��@��??Z=%�]�Mk=?�>iB?��<>Ә>�y������YS�>J�?��?Z�4=%�X�+*�*d?�,�:{�D�K����=P�=�6=
,�rF>�>�$�P�P��Ƚ��<>��>�������a���<�tV>��ɽ���5Մ?+{\��f���/��T��U>��T? +�>R:�=��,?X7H�`}Ͽ�\��*a?�0�?���?$�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�ޅ�=�6�≤�z���&V�x��=Z��>d�>Â,������O��I��T��=���ֿ�2=�>:���½f��������x=�N	���n�${��X �����,�Q$> �7>H9>/Q�>,O?�T?i�>]�=	sֽO*S��ƾ��ｫ�4��0�ů��[Y6=�뇽b���Ҿ!�˾V�������Ǿo,?��h�=S�H�k�����%�e�d��RF�b�*?��>W,���Q����<�Hξ3.���?�����	־z�7��}m�5�?n,G?�|��VS�n���U��ⴽ!LW?�3��T��*��=��� d�=���>e_�=�澇�8���W�B|'?b}.?�^�B_����=�֗�s"�<��?�l�>#WH��'?%'?2ղ�n㌽�?�E�>��=�6L>�`> ��2����=?�$s?�E�C�����=��꾆����!�=Seh>гb�i
��s�>�ӂ����UV&=��Y=7�.=��L?�ڧ>�6&���[^��+!��r�>�R?���>���>y�c?�,E?�W���M&��U)�,����g�N?;�?��Z>�1����n����m2?uA�?��>�`L������X��4���o>E��>��[>�Yj�)q���υ�p���|�@?��v?s^�xs������V��=�>�[�> ��>��9��k�>�>?�#��G��󺿿kY4�#Þ?��@���?f�;< ����=�;?_\�>��O��>ƾ{������~�q=�"�>���|ev����R,�^�8?ؠ�?���>��������>�dx����?��?|�B�Ka�<kD��U�1���tp:�]>�ؑ=�;c����y 
�t�Ҿ@ о���1�)��>�^@?(����>fD���ѿ�9ۿa���­Ծ��G�D@?�u�>��]����qd�"M��%3'���5�ߋ���[�>�0>m0���Z�� �u��3�~�Y��#�>��罳�>hXP�F���¼u����<�6v>���>K|x>V;�����8?�0�Xzſ����D���a�W?���?��?�&?q�V�a����b�����)A?Pz�?:]^?~�ܽ��Y�G����k?#�m��L������.��2�>��|?�@�>wEҾ���� V�LĀ>������c�q�ſ�I�P	����?b$�?WO����>���?�)?U��6����5׾��ž܅>��?�^���[���ʽ�<��	n�H�?Y�C?t��KYT�X�_?ܚa�A�p���-��ƽ�ۡ>�0�e\�6K�����JXe�����Ay����?>^�?a�?@��� #�c6%?�>@���79Ǿ��<���>�(�>�)N>�G_���u>����:�%i	>���?�~�?]j?Ε������U>��}?2��>���?&��=��>���=cr��8ȝ���>"��=yS��Z?�nL?���>W�=6:��-���B���O���w0B��h�>��_?N�J?uf>yѽ�5<����ʽ�)��oټ��C�{����?�$>��9>6P>ɖD��uʾ.�?�o��ؿki��4p'��54?b��>7�?L����t�l
��:_?�v�>8�,���&���F�(��?�G�?�?��׾�?̼Q>E�>SI�>��Խ���΁����7>�B?m"��C��J�o�t�>���?��@nծ?i��	?���P��a~����6����=��7?&0��z>��>��=�nv�ƻ��&�s�>�B�?�{�?F��> �l?��o���B���1=�L�>i�k?�s?o��c�B>��?��������K��f?�
@xu@e�^?!�#�Ke����꾼3ʾ�\��lݽi��=�Y`���=��af�����A�=}�>���=k�����=�̅>�i}>�{��]�&�����
���hgN�r ��!����tl��D���3X�ǧ�$�^�0���i ��������Ȓ
>K��=rT?�Q?�]l?���>>�����>�G����<?2�W��=/,�>��-?M�L?�(?���=揟�/�c�=���񂦾�e��V�>�lL>x_�>5S�>-�>BY�;>J>�?>籁>l$ >\IO=dm��!�<\MI>�h�>7��>�>C<>l�>�´��2��F�h�tw��̽2��?������J�1���;��̉���ݟ=�^.?=�>����<п����*H?픾�$���+�D�>��0?�[W?]�>�갾�U�V >r���j�@d>"	 �Tl�(�)�6Q>�\?
4>W݌>����gh�mAh��x�����=�� ?	K�p>�ۆ���
�)������>t�>b�=�2������҈��P�~K<ʥ ?�a:?�T>�%���������;�>lC.��Re=�I>`���0f��3���͐=�m�>�*�>�W�> ��>�;�=��>�ٮ��FǾ�3i>H�A��Qd=�{5?�5?��]>���=y\2�bjZ�U��>d�>���=\�+>>2��h�=~��>3Z7>Rd���(�%m�UT�Е">4��=�3`��`�=�n*�� =ɋ�=�Vy�J�����>�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾhO�>3r�#4���,{�[�k��ڕ=���>��4?u�ܾ2����L��?���>�s��q����п������>���?d�?��g�i퓿ޛ@�f.�>���?�Z?͠�>�:ξ�����
>�_!?�\??�Ϭ>�#� \���?�u�?�Jm?��B>ً�?sd?�k�>8����2�����u��I�����	>[`�>Tao>�yq�:�+����Ow��>�?�
���=/0=���>�Y���V��h�=끽�v���r���~�>���>-�[>��|>a<?���>��g>P֫=7�ּ @��6��"�D?&R�?{��X�~��N�g[U=� �K��>�S�>���=�����>~�Z?#�?&�P?d�>���y����׹�������Z��[h>�;?Y�>İ��Y?,>������ �W�I>�t�>�=�=�(ﾹC~�q&���Q>�#?.��>b >�� ?�1?�t>�l�>�%�)�}�n�F�Г�>\W�>*��>�?���>.����0�q��(����A���?>Gl?J ?B��>�$������嚽����u�<�ds?e�j??�����?Ϭ�?��?��c?�7�>�{�<�-'�������>�@ ?�Q>�|T�L�@�����>{�>n�>�/s���3� 솽��㾔nq��2�>tpo?L�%?�;�mM��HѾ�g={�����>
�=!#K��:�=I̅=�d޼�X>bY��>��=r"��6i����m�A>��F>"�<G�A�$<�<"=,?r�G�Qۃ���=|�r�5xD�R�>�HL>f����^?Bl=���{�����x���	U�� �?��?Bk�?H��6�h��$=?�?H	?�"�>K��~޾5��Qw��}x�sw���>��>�l���<�������{F��I�Ž+�����>�8"?��r?��&?Vj�>%C>������y�?�����hd���V@���n�|�a�t<�I��l�׽��5=+����'���U�>��=?�N=?;�>(ʾ>ߞ>h@=�J�>��J>�:�|9>���=�:?>��<�Eͼ�(R?�|��һ&���徫ⰾ@?��c?V��>r\T�7��ט���?���?Bڛ?�.y>�vh�@4+���?��>g׀�4/	? L=�l�oι<<����A	�����͍>%�ͽ9��>M�Z�`�?��?I`�i�˾n�ư�5`�=��p?��>�,=�qZ���c�!�x�n�m�!�>��螾=H��/A��P�������텿7�G��:@���:?�'`?������"��!]!�u+�g˽�>��|>�'?��j>�r��-��-`���0��8��UX?Ϧ:?�G�>�A?��/?ƨS?0F?�	�>Gb�>;���7Z�>_�*�7��>;��>i�'?IB,?!*?N?B�%?�v[>.���� �R5�5F?��?�#?Y��>��?fV[���m�|�n��}��O ��P?��I�P=�t�$�뽭WѼ�=��H>3!?�_��`9��d����h>66?#��>G=�>��AB���ɿ<�>�,?	�>�~���p���
���>�݀?���:=#�(>�O�=���r�l�Ci�=?ׯ�(=�=+�q�Ǜ;��=.<�&�=�I�=��9�#��#;˴;4�<�8�>�?�ɘ>=ҳ>P1���;s!���.>Yx> >LT> 
�{k��t����a���>#Ώ?�s�?+�Z=gNA>��>C0��2� ���-�x�:8�>�.?�r?Y�?j)K?�^?S�=������.䎿����Z~1?L+?�>C������礿UG/��{	? v�>v�]�?#�u� �)�ʾ#�W�
>��-�<�t�ͭ���A����x��+@�����?�ʠ?Ot����.�@���՚��*���^�=?�-�>
U�>���>(�,�2|q�>���/Q>���>L?#ʲ>��S?P^?�$7?�ռ<W�5��:���5��U	)����>��I?�k?^̍?�?b�=_�L=��������μ���+=+5�<�x¾�9=~MO>�
>��>\^�>B�>9�x�F��F����C>�w�>tV�>�y�>~B�=������>a�G?/6�>����;��U��\��7�<�0�u?v��?R�*?�I=2���E����F��>�_�?F��?&�)?/�R���=ۖռ3v���Iq�\�>�k�>��>���=��M=j>��>s��>����i��8���H�g?[�E?x�=)Xٿ�%������� ��8���e���V ��9�p���4�羱=�����F���ξY��,���u��.�Ͼ���߀�mh�>��/<���=�n�=:�D=��=�fr��l4��be<�++<S�н ˓��J������96��zd�����<�n�t���h}?�IF? �*?��;?^>�>8�q���>�MQ��?1]t>+{�?��μ.�U��If���Nվ�;s;\���|�=w�P�Ъ>�8%>�{�=/�<W�=_�q=q�x=����o=-P�=��=�	�=��=�S>J!>�6w?Y�������4Q��Y罾�:?�8�>5|�=K�ƾ\@?��>>�2������\b��-?���?�T�?M�?�si��d�>1���䎽�p�=渜�d=2>)��=%�2�[��>��J>����J��W����4�?��@��??�ዿ¢Ͽ�`/>h�m>�Z�>�\�iMD�RA�U�1�Z�����>uT+��=���7�=:�u=;t�������0>�3>�'�=K6��,�`�!�n=�/)�}�<���=9�x>f��=h.�=s,R���%>�n<���=kld>�
t�g*���=t�����=�P�>�\�=�E�>k�?x0?rud?�˸>��k�]Ѿ�{��m*�>q�=מ�>��~=H�C>�N�>��4?u�@?�J?��>(��=�E�>?n�>��*��im�f8龆���3L�<V��?/l�?�1�>� �<��9�����P?���Ľ,�?�,?�f?���>CN�0��02�@�9���������Q�Bw�I
��tM���3R�+��2�=\�Q>F4�>�[k>:>�T>��T>���>�>'��=�N�;2�=�9�<-:=�^>���<vK>�6>� �=r׻< S���K=���=M5=�>-i=���=!��>��>�o�>��="����F%>i0����K��p�= ʣ��QC�E�b���{���.��9��LB>?�U>F��^z�����>7^>^eI>���?Htu?�A%>a���־�%���5l�P�]����=���=ȍE���:�CZ��-L�
'Ҿn��>K�g>鲦>U�>"�$��
H�e`>�D���gݾ(�>�o�=�Mj=wdo�)���������`�o��=\D?A�~���>:̜�?��<?�S�?�X�=����񾷾�ۍ>m�8��\
>�L���!�K��=� R?Z]?��>ƱѾ���8#ʾ�����c�>�S�R�'S��01�٤��l;���>K�����̾n�1�.탿ƙ��Y~G��T}����>�_@?j[�?G�a�ҭ���R�#���� ?��a?6b�>Ce�>�L?V x�z�7'��>.�h?B�?�_�?d >�W=�.���>��9?5�?�y�?�m?�Y`>�!-?�*����>F.�����2L�Je$�m�>�4?A�@?6=?�RֽK�%��A��J2��q�'=�i���>��>�f�>D�>�)�>�v�>��<?^��>Ծ�>Į>���>P}>3#����)��qc?��~>���>G?��>Rl�=I w>�K�宩�ˊ������S�_V�]O�=|m�==��>kH��K>�N˿�?��>ꐯ��c?c��r��<߇n>f�.>��>���>��2>���>!�=&$�>��>2�>��>;�ƾT�#>��2����C���S������W>𙕾fl߽����)٥�L�6�J������	dc����=5�6�=�q�?�U
��gk�
P"��xٽ��?�~�>D*+?@=����6��>���>tJv>�K�+Ғ�R����E�u�?C��?��b>켞>�W?�y?�j-�(0��dZ��t�x�@�hpe��8`��1�����b�
�{�½a�^?*y?�@?�ǈ<�Oz>Β�?�)%��|�����>�/�^�:���3=�{�>���j�_���Ҿ��þ�a��ED>-�n?l˃?��?�Q�E��<Iޚ>S]'?�*?�|3?6��>=0"?ӥg��
?�f>�J)?<}'?Z^*?˓?��?zS�>e�E�R�λ� �=T�%�P��
�س���?��)�Ԕ>�p��J�=�5�=�b�G���λ|�W=��<��<1۽���=���=d�>2X?�*�>f>�>�d;?c��7�����/!(?f��;/({����Z����𾶔�=}]a?���?#�R?ÚP>�>��q7�;N&>�߀>+
>4V>�?�>D���6\��6�=W�>�>T�=���������n�	(�<��2>�]�>J�>��W=L]>��7����>����Dľ�A/��A��P��Š����>4Z?S��>O��a�ݾ4�M���W���>7>x?m�t??��?Vϰ=���c�U�ʫK���۽�!�>�
�n�þ�|���8���0��(�>��?1$��fV��Dwu>���Χ��h�t�O�K��� ޼�+����5�=��۾����ٗ�=�>���k�uڕ�*$���F?��U=�����M�ʊ��>�kU>Ѫ�>)��둅��6�bn��S��=���>�>xs=��꾃�9�q���A>��.?�a>?�Es?e����g�@�D���e��M�>�?������/>��f>�xƼHQ��_�=.z��D���?G�>�_A��<!�(j�<���H�:�{>��>���=�3�>&�"?H� ?�JU?�{?��!?���=S�=�3=��"?�4�?ȩ_=����K�P�9�~XI���>�2"?��7��:�>P�?��?��%?��J?-%?�d>]���2=�tH�>�>9�Z��p��W{>^G?,G�>$�V?�x?)K>�1�lU��3�����=v@%>�z+?�v?��?Kʶ>�f�>~����u=��>u�P?Q�w?@m?o�>�}?�b�=���>�G-=2�>Ր�>>�?=�5?"]?�AK?)�?�{(��ν�뽴�s�h�>�͡=-V%=��>�=;������-����E�;�� �$E���ː;����4!&<�sv=0��>�,�>`-��ܑ>,\f��R��x	>rա���ƾz�i�0�S>�e=����@?��>�p���4+���=]&�=����>�CG?\sF?���+u�?-�ȏ��[O?ɣ}?�BžYH��+r���򉿦�n�Q?�?��3�TQپ��b?�]?� �=�s þ}�a��M���O?�I
?
�H�η�>]?��q?m��>�c�6n��,��b���j��׶=�%�>G>�\�d�3�>Dt7?���>��`>�L�=�۾�*w�x���w�?N	�?'�?v��?�M)>�n�[�& ��t���d�\?"�>$��� ?�z�9c׾W�����������t���V�����m4����0���u�0�	��϶=�?Dbn?�r?5`?�U�4�f�nY��z�^jP��������I��D�q/D�!�p�+���;�4O���F�<'!�p�\�xN�?S�+?+�ɾ��@?�]:�b'��e*w�^
�=V��TQ6�I�>�[u��W���)�>/��I�3��m��v?G?�>���>��\?�'i�23P��?����+� P��䣓>�/�>8�>���>!������\�)=�se���q���˽�"s>�a?)/I?]n?���?1�'����;!�߇9������F>�j>F�>��W���ݯ$��2<���r��������o���
�=�-3? qv>��>��?�X?�%�[�|���0�J�1<�X�>	d?���>��>�н�� �y��>v�l?+��>��>Ӊ���X!��{�X�ʽ�	�>lޭ>��>'�o>�,��\��a��m{��9���=��h?*z����`�Bօ>��Q?6;�:ٗI<*w�>�v���!�:��}'���>�n?�ժ=)�;>әž-���{�I��:+(?z�?E �?;��֨>��"?�L"?aJ
?O]�?�L�>���.�=�|%?�OO?fC?��$?�v�>���)n�%�ֽ0�޽xU�=;9�>ӷ�>���g4=��d��8p��͗���)=2�">��=���=A�<�~!�Ō�j�/�р=�h׿DP��������Q��_U���H�����d��(�|�����Q���i�ƾS�T���9���eF���������G�?7�?�[S�Ah���T��1?��$b5����>����ý�=Ὠ����"پĒ�ဈ��I�V�Z�sA�PE��O�'?�����ǿ𰡿�:ܾ4! ?�A ?9�y?��8�"���8�� >�C�<�,����뾫����ο@�����^?���>��/��l��>ܥ�>�X>�Hq>����螾o1�<��?4�-?��>��r�/�ɿb���d¤<���?/�@�6?ASH�_e��41�<J�Y>4-e?$�>��<,Q���窾�>��?���?c���kp�SX�>��?���=^����F�%�:�;����je=u��?��>��>ߨ(>��R<�nT��nF>��=X)��g�f.�����>Rg�>F)���>2Մ?{\�Zf�q�/��T���T>��T?�*�>�:�=��,?T7H�b}Ͽ �\��*a?�0�?��?�(?4ۿ��ؚ>y�ܾv�M?bD6?���>�d&��t�̅�=v8�Ҁ��)��'V���=��>2�>(�,�ċ���O�OJ�����=�	� rݿG?_��v���/=���<!�=�V���p���	��],־�{������1>)8[=11B�^~h>[x>�u�>.4J?yR?h�>�|�>�T��9���MYӾ������Nt����<,�x>A$�%���33�U�DXѾeվ+���6���=�Fd�4m�?-F���~���b�z�8?(�=H�����\½I�ﾒFm��[j���V���߾a���Ȃ�8��?6L?苌��
L������Xg����r?��'��B�#~	��_�>�)>��T>�Q�>�Y�>���쾤��mF�p�?��?������]�iC>�s�����<o��>?��>������G>�D?k�x��H��7�>Ò<��2>B��>C�>݀�-ĕ�jI? yG?�|]�ptM�R��>F �����S?�=��>��o�t��<���>�i�=DX�:L��`�;�=�sM?$F�>l$��>+�����;ˊ=�9n?�.?7X>�cG?~�`?�T<x��t����޾/|= !I?�cO?��>
�e�%��;�����$?�O?��m>���LcA���D��Y���W?��[?hH?���>`��Ԗ�L���?��v?�k^��n��/��~�V�17�>fe�>(��>��9��}�>��>?��"�l@������\4�޾�?�@Ç�?A�><:�]��=1?^G�>>�O�s5ƾ�c��х���q=6�>�����Rv����nA,�|�8?���?���>����I��nD>����
L�?��?����M>�P꾇C5�Y��]�_=�� >������>��t���U�s>>ľ)!ݾe��>�1q>��@<`I=�?=kf>2X�bݿ�W��3L�ё�j�
?⧋>�N��bL{;e��(}�&�Ҿ�#=����!�>��E>��=(�q��,L���L��=�?D��=:ʳ><����ɾ���Ĵ���H>�2�>׬�>��1�0T��%Ċ?�'���,Ŀ�x��*����X?���?���?�v?��/�����rMO���KX?�M�?_�P?�O�4�:	-�j�h?T���-l]�mk5�+C��R>>�4?Bn�>��"�E�=ZZ>��>�l >��.�Ϣÿ������?�y�?#b徛��>�^�?"�$?yg�+���������'��'<�CA?��0>W��� ��W>�2ב�AP?á3?,p ��n�<�_?`�a�o�p�-�-���ƽ-ܡ>��0��a\��>��8��!Ye�����>y�Q��?�]�?>�?X���#�6%?��>����8Ǿ>�<���>�(�>#*N>>H_�u�u>����:��j	>-��?�~�?�j?˕��'���!Q>�}?��>w	�?�;�=���> �
>\�������&>�Ϩ=��Ž3~?2xT?4$�>�5>z��/�&�E���M����)A�
��>�d?��Q?�#A>���n�j��P'���!�0�S�>��sF�-�7���
�u,>��1>�5>,Y�&����?/�'�׿�a��n)��u3?�>{�?
� ��p���"�߇_?�ω>4�����������pB�?���?X�?0�־n�ϼ�n>G��>��>�bսm���P$����9>�A?r�5��!�o��/�>��?o�@�K�?XYh��	?K��3��>q~�%����6�j�=��7?���Y�{>,_�>6X�=��u�P�����s���>�E�?VU�?/%�>~ul?�4o�V�B�)6.=�Σ>�Qk?WS?ڃ}�*���B>�|?�'�����>�f?�
@Dq@cn^?Ţ�u�̓��y�����p�����=-�f>�mw�6�<�d	=����"z�ۀ��*�>#>��=ڂ�=��>��>����S+�.!��or���XA�#����׾��3���"¾�6.���Ď�-<>�ҹ��������E����>��Q?�|H?�,e?o?�g�x�*>Cf۾!��ʠ>�lQ�=Û>�,?�H[?�%?��;Vѡ�]qj�$�t��鞾��z�S#�>L 8>&�>��>��>5_+��T>�y.>ov>i* >��=�����<P�=���>��?%@�>�4<>n�>�̴�\)��D�h�r*w���̽���?�����J��$��+!��P������=�Y.?ǜ>���63п��c.H?x�Q5���+��;>P�0?�WW?��>j��~�U��=>��J�j�XY>9 ��l�T�)��@Q>�b?�E>�݁>��9�q!��Q@��ܾ�l�=��3?l�Ⱦ.�G���A�D�<��뾌��=b�>H��=�z%�N/���ހ�k~l���<76U?U^%?1�K�4�Ҿ��c;¾̬�>� �>X��R��=E�={FܼP/�|/9�W'">W�=Y�u>:�>�?�>%k> �>٠��#�ǾF��>��-���>��S?���>��ؽi4[��������G�=�>���>��9=ڹ�^�G=z��>8�=&᤽����=�Yu>���=O�X�ߕI;��=o[D���'<L9">H�<G'��:����~?���'䈿��e���lD?S+?c �=*�F<��"�E ���H��G�?r�@m�?��	�ߢV�>�?�@�?��H��=}�>׫>�ξ�L��?��Ž7Ǣ�Ȕ	�))#�iS�?��?��/�Zʋ�=l��6>�^%?��ӾSh�>�x�zZ�������u��#=k��>�8H?qV����O�g>��v
?�?�^�ܩ����ȿ|v����>T�?���?\�m��A���@�p��>+��?�gY?�oi>�g۾"`Z����>ջ@?�R?��>�9�8�'���?�޶?ϯ�?�G>XD�?�7s?���>
���+/��س������=U�;�*�>��>u�����E��K��~���j�����_>��&=���>��ݽ�o����=�w��㨾�_d��ķ>��q>3K>��>� ?�
�>n��>T�=^��	���-�����H?Bی?>��W
X�ck�=��=��$�?�4?�x�P���-�>��i?4��?	�O?���>��tţ�f����?���G<��L>�Y�>���>��ʽgH>���b��v>��>bM����;�R]��!P�"Q>K0?�e?c��=V� ?M�#?��j>��>^\E�k6����E���>W��>iI?��~?��?#Ź�~U3�{��0⡿�[��BN>�x?R?#ȕ>'���{���?�F�-_I�������?�jg?C�v?4�???x�A?�(f>Tt�i�׾���c��>�K!?߯���R4��{܀�'?.�>*�>��9�Yo����=��� �!z ?�_?0�?�C��^�'YǾ�P�<M�3�j�(�jA6=�l><�>�6>������=�=4>�:�!�?�!��=0a>/K[>��-=�!�k5ԽЍ-?>h��v&i����=�Dy��wD��!�>�*>P���=j?��d���|�7������Y��r�?���?�G�?�����d���5?�x�?.�?��>�듾���������@q�0<�{g'>Kr�>��yn�~'��	���	]�|�ƽ0-$����>D��>ߓ?�1�>">+F�>�M��.���Uپ����صP������.�?�"���X���;��ɋ�6���3\�V;�>k��nZ�>��?�"h>�5>b��>�ʛ<�G�>�c>l�a>�΢>!]E>�3�=s�=!#��7����Q?�L��>�ލ羹����$@?Q�]?l��>�P"������-��FT"?A��?���?���>^k���=��x�>���>adq�{��>�b�=�3f=ܨ>��S������9������U�>To����G���H���/��I ?q�?�{����̾|�#�ʚ���bp=5�?~)?�_*���Q���n�sX�RSR���
��Ph�Ȣ�r%���p���������⃿��(�� =�-*?Iƈ?z�����(2����j���>��#e>�g�>[x�>�!�>��H>+
��1��R^��W&�S7(�>o0z?��>H?hX:?��N?��I?4�>e0�>�������>g��;�l�>#'�>7?0�,?2�-?/�?7A)?UQX>[�򽍑���,־��?g=?��?�� ?��?�щ�:Ž;�,��k��x}��E���d=b-�<S����h���s=C�X>��?hy���S#�?�o��>��2?�c�>���>P�3����J4<���>��>c��>a��\e^�GH׾�=�>Z�u?�輙\F<�H�>�>jj����<���<�,�Aa�=����FVs�%U�=W}�=�*;=��a=CX=~k(��Fw��=ı�>�;?⚊>ns�>ǅ������`�=q4_>%�[>T�>?�ؾx���S��>e�|�y>{m�?ó?
[=4u�=]�=����5þ���7���z�<��?%�!?%�Q?�j�?B�=?W�!?�	>� �����Z��6�����?nr)?���>�"��=��畧�;�7�X?U��>�0Z�R����!�Tʾ�,��(�=��$��Vl��;���@<��c���wt����?���?DN��^�-��ھt+�� b��pJC?T��>�ǯ>B��>�U � �g����81O>���>.�I?�ۿ>� O?X�s?�^?�f>&�6��]������0u��^>7�>?��t?��?��x?Lͳ>�E>(����ھ3�侮�꼷ᘽ끾�=<X��>�x�>7��> �>x,�=�m��/�����S��= 5>��>�I�>���>�\�>WL&==3B?Uw�>����������I}����<�<r?0<�?�9:?%3;^ھK"5����^^�>�.�?��?g�%?^��f�=��9�Hi������R#�>���>���>�=�1&=m >�p�>6��>1GM������u��<�?�o3?[�=��ҿi��_8��Ǳ���d�yRn�&�'�[!��r���=l�c�i]#���A�A{�����J��jP����Ⱦ
퐾��>ZS�=�>�q�=d�L�?�<<~>�9>���=a�\�/ڡ�Ŀ�#v���&���&�=6�=��:=ǽ�㞽J{ƾ�sy?��G?(?�<;?�q>�V >|ʊ����>RQA��?ٔD>��r��#��4[1�L�������Q׾+�Ҿs_����ȱ>m_p��
�=n�?>���=-D�;��=mQ�=ǣ=�6_��ȱ<|��=T�=��=}�={v�=� >e4w?=���N����.Q�+�@�:?�H�>���=Mmƾ�@?X�>>�1��L���c��&?��?�S�?f�?�ii�Eb�>U��	���L�=�眽,Q2>���=��2�`��>ɿJ>���D��*����4�?s�@�??�䋿��Ͽ�4/>m��=��>bG�����J�g>fn۾[4V�Z�E?��u���H�9+?6H�>-k��y��<�\>�8l>�M
��L>�{x��'�=f�<Q��;�G�t=�>�~�>F��=	���齵�"��sq>��Z>�t���b�_�h>�"#������<�p�=qk�>�!?!??9�x?�/�>�Е��l�f���> ���Vg>�&A>��W>~�>�?�r7?DQ?�2�>�="Ζ>�ɦ>t��"GU�Ѥ���H��b*>k/_?��?�x�>zJ���3��z� ��
f���޽)e	?W?��(?���>�M��`￶~U�Tsm�h}���?n=�8j>u��x�y5;ۧ=��(u�� R<�_�>�m�>�>�V>�5�����="��>/%><�޼G^=>{�E=䀽���<��='Ǽ�:=>^f��&���@̽04=��=��j<��=L�>�q�=���=n��>�p*>���>��ż�`Ӿ@>x���<�>��44>�׿�X�5��^m�?�j���&�Q���p(>��R>�m�F���`�>���>YM�=�?�ӆ?��.>��Q�s�ܾհ��S�Y�W�!�$�F>)�0>�oQ��RI�mKY��=�/ٶ����>x`�>���>9��>i�@��&�#8=���L3���?HQ���Vf�zI*�X�^�h�}��ufo��2=�� ?'���ޣ<:���?��/?8�?-�?6�%�p-����=��þ*x�=��ܾ�Ԇ=m$k�У	?��?��>�ɾ��"��;̾F�����>��H��P�������0����f��>a�>.ͪ�oѾ:%3��a�����|B���q�>��>'hO?q�?%a�7D��S'O�E��
~��p ?<ug?;8�>�=?vP?O٠�/C��'���θ=��n?Ή�?v-�?W�	>۶�>P��Ͽ>�B�>/�?�H�?�A�?�M�=?��>н�$�Oܙ>��6����҈2���?g��>�\Q?4��OO	�1S!�ft+��x��ԛ=g��=�q?�>�%#>�_�;X}��T��=Zہ>�!	>d�	>�5>O�o>,-�>g�h�D�� pG?��>( �=ZK?��8>{�����,�=]9ֽV� ��޴��鯽��1��QH=�\����=��II�>t�Ϳ��?�P�=�о��H?����ߙ6>N�K>�s�X-Իl��>���>��>���>/��>hR>��>��>$.Ӿ��>m���P!�}C�YR���Ѿ4Kz>!���j&����?���4I��;��\�/�i�U'���4=��h�<_>�?����L�k���)�����w�?u4�>�6?����މ��>��>�ԍ>#1��Ӏ������e�ᾚ�?���?,:a>�D�>��W?��?��:��n8���X�>�u��=�0sa�~�^������j���g��Ľa�]?4Jx?��=?=�!<�|>|�?��$�:��܇>��/�c�;��7E=K�>z��
Z\��7վgRþ�Q�)�B>�~p?�-�?�?�U]�>�~f>�m<?K?�5C?K�?�&c?>�{�-��>/�>b��>'p�>�l(?Z?h�>#�k�k>��q��S>Ů���-����]���X��o�<�>>����u�6��%&>e~�=�쑽�������5����>=��.�jQ�=gIc>��>d?^�?�?h%?�-���о�U ���Q?�X�>C���4���>~�_�N�Ny�<��:?�c�?�c?Y)>�-˽��wg���D��c#>��>{8�>�y�;/㧽��9>t>٤_=��J�}߽�&1��Gھ�롾z ý*FM>�*�>��|>u�~��2>�੾Sh���o`>��b��R���3>��fF�wG1�`������>`�H?��?���=]7�Mr��U#d��J%?�??U�K?y?�=��Ծa�9�SF����=C�>1��<�/Ǡ����ɹ8�ܒ/<�|o>�C��^k��	�Y>����ݾ}o�ZfJ�����C=����,^=[	�t�Ӿ�����=<�>�������b��V:���I?b@�=�2���X\������l>7~�>���>zjK��(p��7=��<����=e��>�e:>p��>_��E�.��2]>�X,?ǯV?��?,�a��P���(�sb/��ؽZ�b����>v�>�P�>!�=cuy=(����׾$�f�s�D��?�?S?:�fQP�󛌾��ؾ���>���>�q*>yl?��@?���>3�K?��>?�?f;�>�V�=y��|h?_uy?�|"=�2��Qa���!�T`D�	�>�P!?�HE���R>�1?|�?)G?�aL?�?+��=r4о�j3�0?�>�-�>�V��;���@�>e:?��>�Lp?9�d?u��=m�O�j4�C�O=mD=���=��
?���>>9?��>���>�6��J-o=
��>��c?��?�;o?�N�=��?t5>���>~�=��>���>�?�M?�s?N�H?},�>��<M���%ҽ�qt��p\��������=����&������ =9�
<���|>��G}Ѽ��(�+D����z;4�>lݚ>�㑾��>0߄��hҾ5x�=�p�=(8þ=��b��=H�����:WTP?�>�%S6���Y=���>xy/>�_����>��B?�c?�x��
]�Z<?�P'a�S�B? ~�?���s����H��w�����]��\5?��?�[���¾��b?��]?Fc�}=�_�þެb�a}���O?v�
?$�G���>b�~?��q?m��>�e�L7n�9���Cb���j�w׶=�o�>[�}�d��:�>~�7?�Y�>��b>f!�=x۾��w��t��x?��?�?��?6**>}�n�4�LB��wя�mY\?���>ֵ���"?��]���Ծ-en��t�����X���3���Ѧ��u��c,!������=��?RDh?�s?n�b?)�����^��8]�����aK��u������E��u?�M:�n�0����쾂����IP<2�2\����?�=?����"?�̲��J���;�e�D>�v��Li�U��=�jg�����T�=Wi���4��z�-<*�?���>�~>�0?'(H���.����^�Q���Ǿ �=MՆ>y��>d8�>4!>J�������Ѕ����du>��b?T�K?Ԧn?� �N�0��U��vQ"���#��%����@>�
>�ŉ><�Y�B��&���=�U@s����������	�ѣ�=[B2?L<�>��>��?�k?�;	�Ɇ��}�w�A�0��v�<��>'�g?7��>X��>|dԽ� !���>�/l?���>К�>zp��ۻ �w�{���Ͻ�b�>y�>2��>�*o>�@,�Pe\�O���C����8����=�`h?S����$b�n��>]6R?M;���A<ؽ�>v܀�� ����yg)�i>%?:�=��9>9vƾ�{��M{�m;���;.?��"?m7�����>�8?�x?^�>Q�j?��5>�S4��DD��T?�.?U�R?9g8?��?1L�ֱ��S���>�d�d=q��>%Ն=�>����=;����W�ԒE����=�?>j�N�Es}=L��=iɿ��A=�=X >)߿�<[�Y�`>�c�p�!��hH�f����O�8貽K���	���8���+(]��f=EI���ާ�!Tپ�0���K�?���?˸$�~�Z�������˾�`�>���;Q	�=�|��dh�C� ������~�p7�o���3[���p�T�'?������ǿy���77ܾ� ?MA ?M�y?����"��8�?� >�>�<A՜�}�������οl���a�^?���>�	�M ����>>��X>�Lq>3������:��<��?E�-?���>A�r�k�ɿ#�����<��?�@�,T?K���w���^�1� ?ԯ�>�=��ͽR��~ހ�"y>��?�4�?�UZ�u�|��78>�8w?�֚���=K��=L$�~p��%�n�|d>��>;_�k�G�,��D\5>��/>�|<ҁa�&^���=T�>Ek��[��1Մ?G{\�Wf�y�/��T���U>��T?+�>�:�=��,?C7H�Y}Ͽ�\��*a?�0�?���?	�(?�ڿ�Uٚ>��ܾ��M?<D6?���>�d&��t����=�:�<���o���&V�2��=Q��>_�>��,������O��J����=�\�)̿�s.�.e&�	�>;�2���/m�����~нe�;��۔�^';�D��F+]<q*>�>�"a>>q>>-�)>PU?�,h?���>\��=���R̄������C�;�s����E��,� ����*`��Ծ�q���'��r��ȼ�N�K�+�2<gI����.�;�}It��_3��?Q�O>�����@��+I����۸���ɑ<����?d��8�p�t��ܞ?ݱE?
�x��K��,"�k���
p�U�O?����vk���kl�n>ְ���>$�P>i��=J[���t�MeO��p+?��)?�4���®�[Ѷ>���<��=��	?!Lg>#����>h�?Ƨ��Z�S�J��>ƈ�=#>	��>(,">-l�����M?m�<?�]����<��ؔ>�T�M3���D��v�>�Kؾ�J��T�>bBg�5��㐳�R"%�vI�=P?v<x>�rF�]o��Mپ~a��
�=[��?ǖ=�~��"K�? �?0k��D��n;�a�#��X�;,,m?/K?8.�=�B����Ax��̀?�Oe?�qn=�����I���T�Ǒ�;$?D��?�d>gr>��S��;�������>?��v?s^�ws�����8�V�d=�>�[�>���>��9��k�>�>?�#��G������|Y4�#Þ?��@���?��;<  �L��=�;?k\�>��O��>ƾ�z������N�q=�"�>���ev����R,�f�8?٠�?���>��������K>o���X�?��?�oN����>v#��������N�!>Q�G>��E��=!V��]���B�("�}�N�8ݬ>Nj>�0@�l6<�y�>�P7��M�]�����G��s1��-?�EE>.0��Q��{iq�5M��
��<H��o�Km�=A6>�ݙ��]�P���v"R�R��=ݺ�>k*=>h̭=���d�߾E0J�j��>% >)O=��?-�>dD�/��?�0O�>���ƚ�Τ��1(?�~�?�s�?t,�<�N���7>^�Ƚ0��=�zS?��?��^?�-V�/D=�tݼ�j?�^��^U`���4��GE��U>�"3?&C�>�-�p�|=b>!��>:f>�"/�N�ĿSٶ�/���8��?~��?�o�x��>\��?�s+?li�8�� \��i�*��)�J=A?�2>Ӎ��;�!��/=��Ғ�q�
?�~0?mz�-.���_?�a�;�p���-���ƽ��>��0��a\�K/��s���Ve�����<y�V��?3]�?��?���[�"�Y9%?��>>����:Ǿ��<4�>'�>�.N>�a_�%�u>%���:�_o	>��?�}�?�j?3���&���7U>��}?QK�>���?�u�=���>�>���#Z��: >��>C������>��H?���>V,�=.
*�i"(���A�Q�C� ��d?��>�?d?q�M?��*>�ܲ�����e~&��s�ő��E��v�_1�)��i��=��[>��9>	�y�s}���?"p�"�ؿ�i��o'�}54?(��>$�?���O�t�����;_?bz�>7��+���%���A�9��?�G�?8�?��׾�[̼�>��>�I�>ս��������7>�B?M�yD��M�o���>���?��@�ծ?Ri��	?���P��Wa~����7�j��=��7?�0��z>���>U�=�nv�ۻ��\�s����>�B�?�{�?��>�l?��o�Y�B�S�1=(M�>��k?�s?�^o���<�B>��?������ L��f?�
@{u@P�^?%�J߿=k��#���U���>�k��<�0�=4�>��UO=��=��A=C1=gp�=\$p>���>]�	>H�=_�<�=����t0&�6?��$�����M�zl �ѝ������D���C���������U�����=Y�<C�8�a�Z�S�$�1E���>w�V?��\?p?
?:_���ۄ>I��bg<K]佅�����>Y�=?��G?n�)?��S=�ۚ��t�Q�n��(���+���7�>�=>x�>h�>�~Q>%�U��jC>``�>ͩ^>�^Y=�^<��ṿs��?>8Y�>蹿>=n�>�;>m�>�˴�m2���h��(w�8�˽�?J ���J����9��6V���ޟ=�c.?��>|���$п٭�sH?�ٔ����+��z>�0?A8W?S�>d)��O�U��>�+�Ώj��� >�����k��)��P>�m?� e> �u>O�3��N8�?O�zx��f~>�5?j���SA�ӓs���F�a[ܾboO>U�>�d��M����~�Fwi�s�w=��:?��?*d��Y���g�r�Kn��9�W>_>��=덨=L�G>I/U��BνNG�J�?=D��=�_>�m?.��>�^�>��>�P���Ws�G�k=�S=i�>Ӓp?.�?PԖ��jJ��6�����;��>Tv?@��=���=�&���۹���?b�>����\&>�ý�Ӆ��ـ>Cx&�Z!���Z��f�>��M�ts�=�m�=8�b�k���K>�~?̀��<ሿF�g���pD?�(?��=E#G<��"�u���FJ���?��@l�?,}	���V�Q�?"C�?������=�u�>A٫>�ξ�L�l�?*%ƽ�Ģ�Ǔ	� 1#�S�?�
�?��/�lȋ�l��2>3\%?3�Ӿ\�>kr�#[�������u��R#=ۦ�>�@H?�k����P�~�=��r
?�?MD�(���=�ȿizv�l��>���?1�?��m�N=��@����>��?$^Y?Ri>]z۾�}Z�ʉ�>J�@?�	R?}��>!*�r'��?�Ҷ?y��?�)G>�ѐ??�s?�J�>7�o���.�.����̌�n(�=/0;�K�>��>�{����F�[ۓ�L���j����H�`>�i(=���>A�ཡ�����=g���f��%Rp���>��o>�GJ>-Ӝ>�" ?ZB�>ә>( =YL��=_��S򙾩�K?۱�?���{n�"�<��=!^��?:4?WZ���Ͼ�ը>J�\?��?�[?W�>L��A���ٿ��y���	�<o�K>=6�>_7�>�P����J>(վI!D����>־�>2���M;ھ�������0�>�]!?_t�>�+�=(� ?�#?�xj>&"�>cHE��.���E�]��>��>;?��~?[ ?9���/W3�	���ݡ��[��UN>��x?CT?�>����b����?�{I�N	�����?x`g?!��@�?<6�?�??��A?ef>���ؾ«���>�!?����@���&�<����?��	?���>HᠽR��2����������?��[?�2%?)|�Lg`��������<GXD��u���3<߾r�U�>��">�U��Z)�=/F>쵩=ܓl���9��m�<�i�=Ƒ> �=�m8������6,?�G��Ã����=��r�;xD�9{>�FL>���l�^?b=���{�����m���%U����?��?jd�?  ����h�4=?"�?B	?���>W%����޾���w��Rx��z�N�>���>�q���ފ��&����B����Ž`J���>���>i3?B0�>m�>;`1>���m_��F���c�	��R�i��$�8�\�(�ź7�WF�rE
�|�P�����������>��i.O>���>X�>1��=!��>o/�hHT>�>4D1>���>��W>m� =;�=���գ�M�N?�4��>�)��x��+��}�=? `b?5\�>���\H��� ��?�3�?�?`w>��i�w,��?J��>v~�ط	?#A=�S����<M��������HT��J�>}Cս�:4�JI��y���?�c?�&��$׾��������	�n=�M�?")?��)�W�Q���o���W�}�R���'ih��U����$���p�/ꏿ"W��t����(���)=y�*?2�?Ȅ���1���k���>�Rf>���>��>ܾ>�wI>��	�V�1�z�]��4'�Џ���]�>#-{?�|�>6L?4ON?s�R?�g/?AW�>�?�վm��>�W}�8�y�Z��>�'C?p?0�+?sy�>,�&?��q=��������0ƾ!?��? ?��>��Z>�+����Խ�U{>)�=D����C���H=�Ի�y�=�Iq�22��,�#>&?[DM�G94�OJ�k�>H?l��>#+�>̑U�/z��~.�^5?�5?M��=�_Ǿ��Y��+���?j�W?�L�oVw<`J4>e�(=ʨ_�h�=�#>�{$=��l=CA�)��j�Z�l�	=�2>h3��}Gܽ�n<|��<�Q<ۙ�>�V?�x�>��>�}��D� ����\��=�}[>-S>>?>ٴؾ�"�������,h���{>2��?��?Ēu=�(�=��=|=���r��6�����[R�<�<?��"?�S?�Ց?jL=?�K#?��>���h��j`¡�vy?^�'?c�>	���˾�\���W2��?��?�d�#.��p ��������'>��,��u}��z���?���߻=x��朽i�?¶�?X_���8���很+�����/�I?{ɳ>�>j�>��%��g����[>= �>1�P?��>$.N?�d{?�y[?l�V>�N7�	��9W������^�'>	>?�ր?�?�?ܫu?zO�>/P>�_'�5���g��U��1e�S�����B=.�X>|��>��>���>�=,:ѽ���z�8��h�=D0b>���>��>^��>[�|>�9�<P�F?���>�"���x
�7�����xӼ �l?<%�?��)?���<���A��`��q�>�Ԧ?崪?�'"?�I>��f�=� �=/����v��m�>��>n.�>��=�K=]��=��>�~�>`�ܽ����8����}?t~??i��=�A޿h�^�Ҿ�����������Q���q�R�[��F>Y� �z�>��\�x�B���-=Fj���從� �d�ݾ�B�>`��=;�Y>�_>^�<�#	��Z>1��<���=���=֎a�mQ = ̼]�#=:H�Tkc�=�0>�Z>y��^�ľq?�vK?��+?��A?:�m>�J>��𽝐�>F��f�	?Q�H>�O���Ⱦ�Q���� Ћ�T���#�Ծ�]\�������>��U��>�N>�V>7I<�=�T�<@b�=��=��S<���=m�R=��="V�=Z��=�w�=�6w?U���	����4Q��Z罢�:?�8�>q{�=��ƾs@?u�>>�2������wb��-?���?�T�?:�?Cti��d�>N��o㎽�q�=n����=2>z��=�2�W��>��J>���K��O����4�?��@��??�ዿТϿ9a/>��=��>Y1^��OW���=����\o���R?�r���3T��?��>�<���8q�|��>gdν�1��J�%���u.<6N/<��=̐:!X�>�q�>p��=$fw��v(>�=�&�B��>���_�{�6�s=e=�s�<�#T=�ħ=V��>�Z?G�)?��L?���>e4��i�����5`�>0�o>��w>�{=ymӻ!B>?ۍ6?IP?K�e>/d���v�>r��>�?E���b���ʾ����\�=_�?�"K?�SL>!����;.�&�I>���ν�&?��+?�`%?Kj�>R���.翽5�G�4���Žv�ּv��;3L��x���]�h�Ƚ+Q�1�>	i�>���>�s>rIp>�7G>>�>���>�;>�I8=#��=�ܻ<y��=gY=���=Ǘ̼�'n�����A9�|<������k�<cǻG��<Ol�<���=Z��>�%>��>�?�=8X���n)>̓��J2E���=��>���b��р��.���,��39>�0E>$�J�������>�ai>��K>1�?Ȣr?�_>���!Oʾ䚿x|��_Y��!�=SR>��Q��>���]�G�J��-Ӿ�<�>9}�>8΢>Qs>W))��=��Wn=��ᾡq1�cT�>ق��W�����3r������ޞ�g���q�D?}ׇ� ��=�b?5�K?�U�?���>�檽�y۾{
=>��y��Ɠ<���8op�F��(�?�!?Hl�>cu�EE���Ѿ�w���h�>�>�àU�����u�-��8R����o��>�󰾜ؾ��:��C��P���B��Y�9��>�.E?�:�?\�L�3(���
K���I����m?��f?ݢ>l'�>�?n��o���Ef�u|=��h?bQ�?���?ܸ�=�4>�F����?u��>}^�?=�?�)?�GU����>iO> �K>�ҍ���[>�L>����|�>�Q�>�:?�4R?/T���Z����`ž���қ�<L�=H��>�]�>�}>=z�=N7n>'���J9�>}6�>]�o>NOU>Zǥ>�D�>�� ������e?4��>��b>�za?u���.�ϼ=y�=E�>����^6�X�=$E�袐�;W�>(��s->}��>$L@>E�ƿK8z?,��=h���Z?�>��� �==�>}��; �߉_>��>A#>EY>7�R>�a׽-׾>t�>&3Ѿ�><`��Q ��A�qQ�Z�Ҿ4wt>j ����&������꽙�D�X�������h�P���]F;��?�<Rُ?�����Pk�� +��C��?��>�7?��������&>��>�"�>�$��v�������=w�ߩ�?���?/b>ߞ>FaW?�$?�~1���3���Y�}�u��D?�8�c�$�_��d������\
��齽�X^?W�x?Vv@?�w<�|>gp�?Y&�[?���։>�W.��3:�P�B=ꧥ>�|���W]�T�Ҿs<þY���ZI>o?���?n?y�T�]�U��,>��;?N2?es?*�1?.>?�O��`#?u�/>��?��?�6?'#.?�?�0>��=�1B��#,=���ވ���gȽ+�ǽ,ݼ{ '=�:Q=4[T�#�;�D=��<��"�Լ�s;?�ɼ�G�<�8$=��=��='�>u8a?eR�>A%�>@�?�OB����D�����9?Ƨ�=m������:��̡׾���~<c?,|�?��8?�Į>%e��]C���_=V>�?*>Os�>�+L>��-=�����ɻ,��=�(>ձ
>U�G&�$ 0��턾�=�>�O�>$9|>�}�� �*>�/���rv�pb>d[S��趾E�Q�dG��0��3w�z¼>��I?�
?�j�=��������f��%?�=?R"M?��~?y!�=�z۾xB:�DbG����_M�>|y<69�)á����9�:�N ���Ot>*7��ɀ¾�(
>ŉ�qN׾O�k�Ȥ>��������h�Y{�=T�����J�d�_>ZH�=��߾�5�.���Nߧ��\H?��t=b���K��Xe��p>>�y�>�Ǭ>�<W�"e�*9>�	�Ǿ8�߻��>aJ`>�#=��D�)�6�f��RĈ>t�@?��f?��}?�k��lm��$6���T��~�n=xK?|�>uq�>��=�=I���������h��2O� ��>�J?�]*�bKL�ä���1���k0��A�>2��>�� >?�?DlH?�t�>%,i?A�)?U�?91�>B災�_���A(?ٌ�?,N=���]��I7��D����>
t"?�u/��[�>V	?�R?��$?�H?�?�>�6�|c@�Yĝ>�n�>6	b�h!���>�G?���>e�Y?2	r?��>f�*�Ʉ����Yf>�a�=��&?�?��?�N�>c�>����|ĵ=���>d1b?c��?1�l?���=}�?AJ+>)��>�ؕ=!��>���><6?T�L?N�n?h�B?y�>�Ε<������|PV��2�<׳<�+<rn�=t���X�4�n�Hל<h
 �'z�@X��6�%��e�V����<:���>���>�瓾�`">vRվ����ץ<>������_Qw���L��=|�D>'K�>�&�>��?��l~=���>J��>���-k?ܨ?bS?��2��5_�Y8���s����>�P?�In���J��0����v��4;<hb??9g?V���(�b?��]?^�s=�4�þZ�b�d���O?�
?n�G����>2�~?F�q?��>#�e�\1n�$��V5b���j����=l�>�V��d��K�>$�7?9>�>y�b>u!�={۾]�w��a���?a�?� �?��?U!*>��n��/�WI��:{��Ow\?ˮ�>l���"?*�.�5ӾJ��������� ����g���ҥ�x�)�"D���Hٽ�9�=�?�Ws?)�q?+3`?�� ��8d���]�	�}�n�T����e��4RF��"F�)D�Rm�������P���X<=t�2�_�e���?g�.?�O��=*?*�.�����!�����>- Ҿ����h�>�N`�+ѽ�U�>�~�������Z"��?l��>^��>c�?h�9��R��Ѿ^�/�R��v�T>��>RQ�>�T�>G˼c=��v�C�Ǵ��$澁SB�}_v>�\c?W�K?��n?h��1����o�!��x/�����zB>~=>7�>�:W����T'&�V8>���r�$��7���{
���='�2?:�>��>�C�?��?#W	�e����y��[1��ۉ<��>�i?��>��>4�н� �s9�>kUk?\��>��>����Yb�̀w�NϽ�?�>{��>��>c�l>6�&��C`�%c��fێ�;e6�?� >��i?����)X[�V�>%�P?�ﰻOX<�>����i"�yO�;,�V>d�?�r�=n�0>:�ľ����|����F)?�Y?�Ӓ���(����>�"!?Y��>�-�>w��?�o�>@����@���?M�]?\uI?��??���>p�0=�r��f�ƽ2&��B=�>!c>�zp=~��=7c���c�. �dB=
��=�fȼ����$�R<���<��<�.>��ڿ�7\���)	ھ���������k��ݗ��+��}��rL	�������彰 `������>�Rɖ��6ϾD�?��?r�ӽ$� ������������?����A����r�}���^��+m��U�u�-��2P���R�M�'?<���ɽǿﰡ�:ܾ-! ?�A ?;�y?��T�"�^�8�;� >�A�<@)����뾢�����ο榚���^?Q��>��t.�����>���>��X>Iq>����螾�2�<��?�-?���>��r��ɿC����¤<���?#�@m�=?k}$�����ɱ>.P�>}z?=�>�74����f���"����؂?�œ?d�V��o���%I��V?��%���'�hȽ�ר���=l1r�,_��a@�>�m?�����i �\���]p>�E�>�B<�e�����}�Pj>n0��g7�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��=l��RJֿ�dM��U4��ú��퉽��F�ن�vX�;%U��'ӯ<��$=,�>!U�)�9=�r>��u<>=�L?��E? 8�>�k>`0�љϽ�X��~FD�^�4��g�����w����x���ʾ���9���$�}�־�9��u>ȍK�����pN�'ie�Xxc��$?T/�>	���-B�?ݤ=�5$���ھ��;�.=k�̽X�+��Z�;��?Z+?�|��ilK�/0׾3 >>0篽VUC?N����#��]޽�f�>���=��=5:�>'F0<D.'�TK�r�=��u?ԁ&?f
��N��o��>c�[�r��=�E
?��Լ6;~��+�>w�?Cd�Kk8=��>vF�=�,����>M�I>�鶾(�Y���3?j`u?6֪�w��a��>m�R���:�>�7>��<�
*��C$>���d�b�>�8>�t���@�>��6?�Է>������Ks����W���>��[?���>8�q��}K?�@?����Ƃ��,���Ș�;r]H?z,?^\>f������"��M�`?h�]?�Ʈ=��<:P��lB���ľ�=�>�)�?�2?Z>cmm�����O<J���?��v?�r^�as�����t�V��=�>%\�>���>��9�Ik�>��>?�#��G�����Y4��?|�@��?H�;<��	��=�;?�\�>��O��>ƾ�{������K�q="�>^���cev�����R,�0�8?���?Г�>C�����k)>ַ����?t�?lxk��G>��A�C�G�xӾ��>К�<�'����=q��`�E�
7����E߾����a{>��@�S>� ?yZ=���%)Ϳ�􁿁�ľi{i���%?�W�>��1�t�����x���b��w�5�19��)$Z>ڏ_>-,��N���k�iM[��59�D
�>ɑ�>V��>o$�A�Ծ�p�n]�<��>:?�� ?)x�i�̾V��?i���Ͽһ��-����??gg?���?Ω>b���!=)�%>� �XA? �(?�\?�\��f3���=`�m?�2����Q�B�#��
!�Py>X#7?���>Z	�B��dK���q�>Y�,>XN��ս�N6��;¾ñ�?�=�?��Ѿ���>:t�?z6?�������%�9�d��V�?�Ғ=�浾E�'���@�z����.�>�?ܥL�v�@�Q�_?a��p�a�-���ƽ@ۡ>��0��e\�K�����$Xe����EAy����?^�?k�?N��� #�E6%?\�>4����9Ǿ]��<q��>�(�>�(N>|D_��u>����:��i	>���?�~�?*j?ܕ�������V>��}?�>6p�?��=O��>�&�=�?����:�Y>���=?vm���?ML?�s�>���=�w��-�M�=�ݕM����|�D���u>��e?��P?ΞT>����� � �$�#�����2�e	(��($����>l�:>ܿ7>��Z�Dʾ
�?�l���ؿjj��b'��44?*ƃ>S�?���%�t���%9_?煈>�>�;*��'��-!�b��?�J�?��?��׾2�̼� >��>NB�>/սeɟ�Tr����7>=�B?�3��B����o��>}��?�@�Ӯ?��h��	?���P��Ia~� ���7���=��7?�0�/�z>���>��=�nv�ۻ��N�s����>�B�?�{�?��> �l?��o�N�B���1=-M�>Ȝk?�s?�Fo���6�B>��?������L��f?
�
@{u@X�^?!o�ӿJ���n׾\Ѿ��>�9s=��P>��ƽ��>þ=�{��&U���I>�>F>i>L�\>�$">�(�=���	�(�)������{n:�0I����9DQ�b����Z�$}�Q�Ӿ ��v����xs� %�i�0��b2�A=N�{��=NDU?�8R?�=p?�G ?�v�4 >,a����=�!�)�=`Ȇ>=2?�kL?;�)?q�=�;���	e��>��`��`����>��I>�-�>�:�>���>��:��K>�;>>�4>�� >��'=2*�eA=�TN>���>��>_"�>��7>A>�b������i��;x�$��j�?Cq��t�J��J������;,��Z[�=�-?�F>CK���Ͽ�g��b�G?H���u�t�)���>�90?P�W?�c>m����}r�N>��1b�f
>��IFo���,�+�Y>��?c�f>�6u>Ő3�Q`8��P��p��W|>�*6?�� E9��u�ܜH�3aݾ0LM>�ɾ>e�D�;j��햿�~�q{i�m({=|:?��?󇳽�ా-{u�!I���?R>uN\>v�=�g�=�NM>Sc�)ǽH���.=��=T�^>V[�>ǌ�>��S>���>OȾtY���'�>��Q���>��E?��?�N!��d���f��!$����>��'?"�;tM:>�&�i�<촎>�:>�R���o����C�}��>��{��(�`[Ƚ�.�<گ�<1F���0>ʸ���&��A�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿth�>dx�tZ�����w�u�;�#=���>�8H?�V����O��>��v
??(_�֩����ȿ�{v���>h�?���?H�m�~A���@�b��>��?fgY?�oi>�g۾�_Z�Y��>��@?�R?��>�9���'���?�޶?ݯ�?�I>Ɍ�?(�s?�j�>Bx��Z/��3��1����~=�\;�^�>�Y>U���CgF��֓�)g����j�9����a>T�$=��>�E�64���-�=�����G��+�f�
��>�(q>G�I>
U�>�� ?L_�>#��>��=�d���߀�������K?ݙ�?C��b�n��E�<ƽ�=DG]���?��2?���x�;?˨>�3\?<V�?��[?>��>���ѧ��c������{��<u�L>���>���>�`���bJ>Svվ_C��ŉ>�O�>?���Lھ������ݻs�>M!?�9�>�-�=� ?�#?z�j>�%�>�bE�1:��a�E�Ԯ�>]��>�C?��~?�?ڹ�TW3�����ޡ���[��HN>J�x?�T?Õ>U��������D�EI�2����?@gg?V��?.�?r�??�A?if>�g�6ؾi���|��>8#$?80�5�3��)3��<��?��
?a"?[���R(c�"Q�=�����ݾ�n�>��w?Ϭ
?�e�J�=�5n���:;���;?���+%˽�u=N�$>���=*�.����=_I�=���==t.����"���L:>9�i>賽=ת ��w�=,?��G�kۃ���=^�r�/xD���>�IL>���=�^?�l=���{�����x���	U�� �?��?Jk�?	����h��$=?��?S	?I"�>�J���}޾���*Qw�qx�qw�{�>���>��l������ϙ��F��p�Ž� �����>�b�>��	?�F ?�V>e}�>f��F�%�(���>�
�,�W�-��;�@�Z�.�����+��#�$���T����s�J��>y����g�>3?�ez>L9^>A�>�;p@�>�$a>:�w>Ƞ�>Ar@>�K2>J�>� ⼊��k{P?�績��&�`��\b��L;>?\�a?�Y�>ٚ����ԩ�B?���?	��?�|>�_e�U�,���?�� ?sb}�2�?~�L=���<�j���"�=����6��9�>��Ͻ_�7�A�J�%sh�O�?�?��ͼǾ���z��8]=���?�,,?o1*�DsP��|p���[��F���μ�h��3����'�FCm�ˋ�;ņ����k�'�/6�=,?��?Iy�z�߾I��u�$]A���>T~�>���>�E�>�0>D�o�5���U���j�j�W4�>�y?6��>��E?p<?ڬN?�J?�>�%�>*+�����>�<jZ�>���>�W5?Q�*?2j(?��?�(?6�N>�3���J���־��?�?� ?��>4��>􅾔����=<��u<l�z������=��:@������<)�8>U�?])a='M�1��,��>R?���>�x?�@�Fl�1n�=��>�3?^8�=�,��M��	�s�?"u?��L���	=	^�=f�Z��^�=�H=;�6�.F�=��)�:(�='k�� ���$���P齲�k>%v̽�q�<��:=�e<J��>��?�/�>
�>�����z�8��`�=�\>W+R>k�>�%ؾ�]���闿�kg��mz>[��?�!�?z2n=p�=�<�=p����	������U�����<�?��"?��Q?�t�?�Y=?L@#?\X>pN��h��M7��)m��v�?r�9?�1�>�¾ѡ�HǍ���G.�>3?м{�6$ܼl`��qؾf�޽
��>��9�B>d�ͧ��e��^&�j��� ��!�?譥?n޾o�.��ξc���U�>�/I?!)}>1�>Z�?!�ts��<�C��>5��>�A;?( �>��O?7{?��[?LET>��8�t���ř�J�/��">�@?Ϥ�?��?/y?�J�>��>�R)����(�����z��ꂾ��V=u�Y>Y��>��>]�>�Z�=_Ƚ��	?�3 �=Üb>�b�>���>��>�bw>u$�<P�:?��>5l��t4�kF��h����nR��Bl?�ɏ?�b?��=e��F��p����>i��?h�?ib"?�!��>/��T׾��y�l'�>O�>oH�>��2>F��������>Cw�>E�����<��n$=���>�E8?�%�=<b�
Ν�U��H���s(Z�&�_������v�����=���w�>-6;8P��S�q��Ͼ�ȡ�}�2�E.��*	?��>PI�=��j>�n���<D�X��=g�P�=0�$>?U���X� u7��(=�.�=v�J�`i>�lX=ڑ�T��^~s?7�E?i�*?n2?�F><�)>Tе��a�>���;�?��Z>"���SƾI�$�+ٌ���R�d�Ծ��žmCi���� >ʖӼ\>��>N��=5�.=vB>*��=��=��T�o�<_�>�^=�1�=9�/><Q�=ͺ�=�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=J����=2>p��=v�2�T��>��J>���K��B����4�?��@��??�ዿТϿ6a/>(^5>�>�D���8�dϸ�8�۽Sா� :?��;���)�PR�>B�->�vо`¯��"?��_;��	����>J3��l=/����>�'�2�Ӝ>	A;>F��=NS�"!)�B�漱a
>���=+02>}�
=l�t=LZ����Ƚi
�><5	>:<�>��?�,?(VV?Nd�>���J屾:=��'�>�(>�2�>�%�=�.�=��>�'?wV6?��W?��>�w�=nd�>���>4�/�b���YQ��XL���?<�?��`>�.�=�M�&}���*�?�ɽ�?W�?�y?>��>�,�	X�X�)��3�)���Kl9��,�<�Ղ��N>�Z��Hb��[���Q�=:��>���>I�>�q>y�7>O�L>�=�>ր>_	=�Y�=�� �3�<���s�I=�v��~��<���@:ۻ����6�#��'.�Ǝ�;�\���$��n����={%�>n�>j��>0�=�����^,>M$����K��<�=������A�y�a��;|��e/���5��CD>��S>ҍ��4��G< ?�:[>A�D>�B�?-/u?U�">8*	�� Ծ׆��\�k���M����=E>�=�T`;��_�N���Ѿ���>B�>��>*��>1��<2��#�<8��)��?K�~���ͽ�X���:��n������3O��H�ܥ?����D�-�^R�?�ka?>;{?@�>	+�&����>}Jz��B��?�r
��՟6��9
?N�?i�?v���8������轼i�>w;:�g�����S��ώ�9v�����>����ݫ4��N��1x��#j���G�8�'�4$�>�)?�y�?A#8=�9E�߇F��*�g��8�>?�Q�>�? ?�g,?e�=q����wA�="D�?��?V��?���>jVM>:{����B?��E?ʮ�?�?��?>�
�5�	?
!�>�-���� ����>5O�=�z�� �=�P?���>Kf
?�i���� �w�����Q��h\>���;�z>�%�>�J�>_�ƽ��ƽ{�<�L{�@�>g�"?Yp>���>�Tu>��j����D?�D�>�QG>҈??m><�0�� >�
��Ps����<;�^�O��K �
�<ױ����~���>��ʿK=�?��m>.�龿C%?���!�Ǹ�Đ>��L>J�Q��9�>Ρ�>���=r�>��>h	>���>�4j>�GӾ$v>g���a!��,C���R��Ѿ�xz>k����&�����c���@I�^i���f�^	j��,��0<=�3��<�F�?������k���)�O���̕?ja�>�6?Gތ����}�>I��>�ɍ>�B�������Ǎ��n���?��?�Aa>�b�>�W?kj?�[4��8���Y���t���>��b��%`�씍�������缽�_?�\y?��@?���<��|>�?HA&�����D�>��.�>;��\R=�¦>�w����[���Ѿ>�þ�q���E>!p?飃??��S�W���~�&>��@?��1?�Lr?D�1?�c9?�]�C1&?Yi+>���>t{
?ը<?��0?)��>�5>G��=�O;�Ɍ�=ؐ�������t�����r��{gg=��=-�<m3=�)�=��=$Fl���ٽ��^<��\���<@�{=n�=g��={�>��[?���>|�>G�.?d�/�A�1����!9/?�n=τ�� u��R���"�8��=r�h?�i�?��T?�mk>d�9��?�h�>q�>q� >�oM>�t�>C�Ƚ�!7���O=[�
>�>I��=R�-�#��8�������=k8>��>?�z> F��U`->������y���b>�R�� ���>P�?JG��1��q�3�>x(J?�?s��=~0��$����f��&?/�<?�N?�M?=��=��پ�%9�LI��Z�:S�>��<����9��bˡ�H:�P �;�mn>PM������z+T>R����6t�{Z�{�_O�=;���%�=�Hξ��޾	ᶾF��<��;>26��:Y�̦��0���??���<,py�6Nн)�𾹺�=��>@�>��H�l���:��P��s�<��>Jr>U/�<-l��/�A����9}�>�D?a�]?GM�?O���5r��?����%i���ɼ|�?���>�?hC>�a�=K���g���jd�KG�0��>���>����F���]C���#����>��?�4>>W?7R?U	?�_?�)?�c?��>����
���
� ?�?2��<�罽����8��mH���?��5?�JY�Ġ>G�?�?�?!T?��?ZQN>5E��:��>�b�>�.\�,��2_�>�<Q?��>��T?T	{?͐>B1��%����h��u>�B�=Ҝ?�_?�?��>w��>[B�����=�@�>�f?�~?��s?��d=���>)�=��>T��=]1�>�, ?��?	vD?�z?�O?��>A\;<z�۽�B⽿���;������<`L�=S˪;)��+M�M��3����2��㟺�3��|1�7�r9P|?4�l>����<��>-���Ec��ʅ>	x��콰�����������<Y�hN?�IŽ���M��;���>�oս�i��M�>�(?�!!?�+��c��	2��Jܽ0�>�u?b�-=�q��O��#�h��l�LG[?��u?Y����	��VX?ɁG?X����D�,ľ���8b˾s8L?�=?��6��>�=}?��`?���>�#!��v�aӘ�>�`�Ik�c��=e��>���g�q��L�>n�6?��>�Z>ZO[>2̡�u5]�r����d?[��?���?���?"�>��s�p̿���������]?'��>맦���"?		Ȼ��Ͼ�����ԏ����`{��hM���s��@���'�0a��"�׽��=,�?,�r?R�p?l�_?�� ��c��]������V��O�b���E� E���C�x�n�0G���������K=���e9�?_9?±��H??D����3�%2���>A�)��������>���,z=g��>8l�9&��>&-�V�>:�>���=��,?�>�ݰ+�}����)�"���D������<a0�>��4?�{<ü�<�V�< ����s���ͼ8`>�']?B�A?�j?.���(7�P��.���\�������:j>��=��Z>~Oe��u�� �aw5��Ym�~�����K�
��c�=1c4?�B=>1=�>��?:�?m��Iా푎�]Z)��i�<«�>r�a?��>��>�\�����>�p?�2?X"�>�Z�:��3l\��T��p��>|��>�� ?�d�><�ܽ;xL�Ր���ӗ�&�6��>��_?�̀��J���$>>?2!>�]:=��m>��5�q1$�X���'���<[�?��W>�Hy>�.y��h��x�g��4k���"?7V�>Nx��d39�}�>��.?��>ǉ>|t~?f�>6A��ƊW�K?q?`?IdF?ʸ*?|[�>V	��N��=����콰RT=�Z�>��>*9=o�>�9x��x��C4�O�=�)��=wm�j�������d�<f�<�u�=_>�T׿��P�&�ݾ��޾��#�
[(��Z�L/�2���'�H)���㾳Q��qCݽ<���>��O�L������j��!��?	��?J7���]⽗{�������J?TG��20I>/����$�HԸ�(�,���ؾ���Q�N�|�իp�}'?'����Yǿ�\��E�۾M ?0} ?�*y?�����"�,�8��!>�9�<�}��xa��՚�4�ο���ʋ^?�G�>|)�u�����>|��>�Y>�Eq>xY�������<�?��,?��>��s�8�ɿTF���Q�<#��?��@��=?Pl��%ξ���=�c�>f��>���>B�F��(�/c¾aŷ>L��?��v?��>_=>���(�^�5?��M���6�޻�H=Ȏ=̰E=;�>���K>��>�U��!(�#�+�)>L�Q>��p�lm��G<��pF�����=��ȽZU��Ԅ?�z\��f��/�`T���X>��T?�)�>]>�=�,?6H�0}ϿC�\��+a?�0�?U��??�(?ܿ�ۚ>��ܾ'�M?�C6?��>�b&�`�t����=W��J��	��B'V����=���>��>�,�����O��>��}��=5�	�;?ؿ����J�]:V�M�ͽ��X�q`}�����;��$Qݾ��� ٽ$��K��=Y�>���>ޫ�>"�J>��G?g3J?o��>�݉>����혩�	0������y@�E6����5�;ua���X��Ô�4ӳ��2����Fְ���(�Eq>�e��w�?X.���}���O�1�;?��>H]�����ۜ����Ѿ&�<�����\}���'��h���?�d7?�p����g��p���=�P���_W?)IͽO� L���4>���H�=�4s>�A>�C�sr��h4�c?�@&?!|�l�k�Q��>@us�H����?po?�F0�h�>[�-?|����Dξhٻ>��>��<�=�q>�w��|yJ��?8?��_?�IӾ��羆��>aľ�=��&=n> �A>!	�^�w�ͮ=Ti>�
��=!��)5�0�9?�½>�>C�x��fw��֎ټ4:x�Kw�?v@?��.>{#(?{0?v��;i���o� ����>bf>em?��O?�X0>�H�<!_�G�;���G?<�?&>ʽ�[�:�q¾q�;��$����>��?���>�1��/X��f����
�F?��v?�r^�s��}��O�V�'<�>�[�>���>f�9��m�>đ>?�#��G�������Y4��?p�@2��?��;<�$����=t<?�[�>>�O�<ƾI|��܄���q=d#�>����fv�����W,��8?ɠ�?;��>𓂾?���(>����ҵ?�p�?�ۦ�ne>��޾Ɠz�۫�?�>����x�<���>ҵ����ΛE�PI�kڽ�n0<��r>=c@�-��{x>	$=�"ֿЧ��ڗ$�����*����?�d�>Yy�\_s��?��R_��>b5��g��q�TQ]>��(>��N��-���Ӑ�;�q�g(��1
?�y_>Ȇ>R�=쵅�H!��DI��� ?:�>&��>,�B�P"���?�m���ÿ�o������p�a?3�[?5�x?im!?�s\�Ȣν�%���'`;{N?
�M?A?b6=����<�=��j?T\��?`��y4��1E��9U>,3?�(�>��-�
�{=��>+p�>q>�/���Ŀ�ݶ�����5�?���?8b�?��>x�?�g+?�\�n)���Q����*������=A?�j2>F���L�!��/=�Ԓ���
?If0?�|��&�ѵ_?;�a���p���-���ƽ��>�0�v\\����q��7Me����N2y�P��?^�?*�?����#��:%?��>a���P8Ǿf�<���>�%�>�N>��_�̇u>��0�:�AD	>X��?�}�?�f?��������
a>��}?\޷>�?���=���>��=�Ͱ�������)>c�=X@9�J ?�7M?���>���=(T8��/��	E�!�O��j���A�X�>�`?&}I?�^>�ĽhYD��G��~ʽ�e1��z
���>�pg0���Ra/>��:>��>Z9���Ѿ��?Ip�8�ؿ j��p'��54?$��>�?����t�V���;_?Qz�>�6��+���%���B�^��?�G�?<�?��׾�R̼�>F�>�I�>`�Խ����X�����7>/�B?\��D��u�o�w�>���?�@�ծ?ki��	?���P��Ra~����7�d��=��7?�0�%�z>���>��=�nv�ݻ��S�s����>�B�?�{�?��>!�l?��o�Q�B�{�1=:M�>͜k?�s?Ro���Z�B>��?������L��f?
�
@~u@]�^?)X:��ͣ������Ѿ�qY�3�=��>س���b���p<w4��@q�8�->N��>�s/>�Z>��>�>U)T=������,��6�����PoF����q�$�!���O	��4W�|�о-:�y܁�9�1�fQ��n���8����8��T����>�K?�T?�Om?
� ?=��>���\;�����X�<r�c>9�9?uL?t�?4�v��|��1o���u��+����>��>��1>��>��>R�>��1�[:>7�3>�m3>��>>�g*=��;�.�;$v�=FY�>i��>�>ec<>�i>�ϴ��@���f�>0v���׽v �?���@�J������h�����{ؗ=��-?��>����5�ϿOk��G?�]������+��}	>��0? �V?��>q���xa�a_>��Q�h��f>�����h� �)�h�P>��?*d>�u>(�1��5���O��P��Ԙn>_�4?M����6�%�p��E��{߾��=>�տ>_�U�5f��T��]B~��Mh�)Iw=� ;?�W?M黽cڱ�l}b�:*��twR>b>/��<�T�=p�C>g�`�͝Ľ�I��k=o��=J�P>h?�>��-=���>йf��;��C��>�'>Jv>��B?�g�>��qǥ�@���\`==f�=D�^>���>'E�=�|콨��<ij>3o8>���VR���S��l���r�=�����2����Խy���=��=L{j�b<� =�؎ڽ�~?{���㈿�뾏b���lD?w+?��=��F<I�"� ���H��
�?e�@�l�?��	�̢V���?�@�?�
��+��=�|�>H׫>�ξ˔L�ı?� ƽ�Ǣ�	�*#�;S�?w�?&�/�Zʋ��l��5>�^%?v�Ӿzh�>�u��Y�������u���#=���>G8H?�R��W�O��>�Mv
?�?�\�詤���ȿ�{v�F��>F�?���?�m��@��\@����>^��?�eY?Mli>2j۾<`Z���>|�@?DR?��>�:���'���?�ݶ?D��?�,\>���?�|?���>�΅�x�"�ƫ���c��v�=�җ=w��>" j>�]��E�u����m���we�rB�G�=>e�=W��>�0�B���V?>�"��?���9����>��T>R>ú�>��>7��>�@�>m�3<�"D�_Ge��h��_K?Am�?B���8o���<��=��g�],?�{5?F���gо[ש>\?��~?\�Y?���>X�H{��K���(ĳ�d��<V�H>6��>��>������F>h�Ҿ��@��>i��>�3����ؾ����i�J���>Z ?e��>^�=Î?�d)?���>�>� =�|��l�3��>�&�>�?M�?�H)?�-���(/�N��~���_cZ�=0T>ڕb?o�?q
�>#Ҍ�����F�˻����w;1��? ap?iݢ��u/?�̈?@�?��4?9z�=��������W�]�5>��?��&�s-���=��
���?��?�O�>��C>�R��\�>���bG���z?a-j?X��>X��]j��<;�=�=v��昽��;�>�2>��>E�)�S��,�]>�PP��aľ'��j��>&�=��>�~�=��m$>T2?��v�d���{r�>�4��
%�܈E>��q�zUt��j�?0;������Y��%��� ^(�G*�?�?�?\n�?Kۤ�*Wk����>7X�?-.�>�e�>|Wk>0Ǿ:� ��B4�t%�� ��j���+�>Θ��]��̈́t��h����M�CH�=e*��y�>>{�>B�?�?�<�>?i|��ZP�	1�H达�B���A���]U��P�$�����vg�#&��k����ր>Me����>�?:��=78�;��>� .>���>�mV>���<7' >r �>̇�>�a��!��֓=�K?����"��S���U��E�6?-!g?��>�v�������ﾫ�"?T&�?�|�?8!6>}�i�BY7�74�>2t�>�jn���>9�;���s���,��}O3����;��\<�u>ۼ��5��2?�,�d��`�>U#�>��9�Ǡ��$er�q����W�=�ˇ?�*?��'�-�K��\l��U��N�FMV�'Q�b;�����ưn��e��8@��Z����%��<=Ba)?.ŋ?JR �Uc������
j��(:����>��>�!�>��>�=g>i/���,���f��2�	}���>z(r?V1�>��M?T�X?IB?5[f?��>���>�0��z;G>�N\��
>��=��<?��J?�"?��?� 7?Nus=�RȻ�sǾ̾#�>g?�~!??��>t��>�_B�i�*��14=�Ju�8(�WQN�`&����6c���:����h��?�9>�0��+&�a��>�c>?8�w>��>�\`�S6��9`��)��>�B(?׫�>�x�8|6���վ�M<���?tL����e=�f>��>Ķ�<�����S>���rǽ��N��w;�+ >�/�=,��=�Q�=1���v����&>���]��>k ?�:T>C�]>�^��N�x���b3<�a�>�ha>.=�=	��T����4���r]�܃>HA�?���?2��<�e>=�=u�ľ�ƾ.# ��.�ǼV�?&?�EB?&>�?�r;?�:?v�6>=&�Y:��V��x���{�?�,?I�>�&�,迾�'��?�2��?
&?&/]����M(&�q׾���_>��0��v�筿�?D��i\����c��O��?�j�?�&����4��!�͗�⌯���F?���>���>��>`,���a�"��1wM>BO�>�yL?x��>8�U?g<�?�0T?6z�>s��8�����xY$��->@U<?�ro?�֌?�y?''d>Wl�=D�D��ɽ���i��[�j���Ђ�wdI��H>��>���>���>/�}<�+Y�D+���M���>�4�>���>\�?��>��:>�{�=q�5?
��>3���n��Iʜ�L����rս}FV?}Y�?sf?aZ7=b���N��,�l��>E۠?e�?���>�`����>��<��Ͼ��~�=л>B��>��>?N�݈ >&�>�Ҙ>c�>��Ar��,�i?�\?��R?Rn�=��ɿ?�y�{�Ap��~�m������`����2�`�䟎=r��x�����!l����vœ�`���C���7�. ?�B�=F_�=3�=1��<�ּ1�=<5=�؆:6-�<D��5����b�\�����袴;��<���=�n�&¾��{?[JJ?}�+?�}I?0�>��0>�U����>�@J�@a?�FL>����WF��wwA�L���/���޾3wؾ]�a�כ��K�>�\�u>*�.>��>�S<��=Q�=�%i=g��;�<$=�^�=��=Ql�=C?�=�>ԭ>�6w?V�������4Q��Z罤�:?�8�>2{�=��ƾx@?�>>�2������|b��-?���?�T�?>�?Rti��d�>T��F㎽�q�=T���>2>p��=~�2�S��>��J>���K��,����4�?��@��??�ዿ̢ϿBa/>��=���>N���R�b�B=3Ƴ���8��jw?&k򾝧ܾ �?��>�-�kl���=�t>��E���=7E�w��=wF�;���=���=�%�>�w>O̼Ï�6 >��G=#�^=�X>�c缫ض��$<�eW>2\=Q	>���<e��>c? �.?	x\?v��>�d��þ�����6�>Z�=O�>y{=�?>ӵ>��2?�gC?�VA?3�>N��=ݝ�>���>�'��e�^��F���<�7=~��?rk�?ծ�>��<U�>��3�n�5�
�>���
?Wq6?�=?�>���;�� � QZ�v�X���-���E�`Υ�0�������l�����>�c=��\>�q>��p>���>m�y>�x7>%��>J�/>_>��@>
N���J��~�<�:k=�	��>���%�s���/�iGJ=�9�=f%�=#��~�=�0�=*��=���>r�>���>7�=/��1/>�Ȗ�՝L�t��=�,��8 B�>9d�^9~�T�.��66���B>.�X>2������?�?��Y>��>>Um�?GSu?OK >2���վ5K��@e��}R��Ǹ=��>.=��U;�?7`���M�ScҾ���>i8w>��>���>y`�,[(�q>F���;��8�>Q��� -��=���S�J��nH��bkf����o�$?�>y�Q��=�*{?{5?%w?�=�>dN˽���T�*=f��/�> �[���i@Z�%c)?�)?5��>�!���.��k־+Ʒ�;�>��&�y�^�]��_',�M�<���Di�>�M���c侾�5�&膿U"9A�>|M��.�>Y=?���?j���AÃ��D��o�¥콫Q�>��o?�β>��?�[	?ذy��Y��k%��w��=y�t?�t�?L �?>[�=�U`>)T8<?�?��?�r?'�?U���ߟ'>��U�����z��Z��>�	�>���=��Rb�>�8�>��,?�zl�w�ؾ�G۾HǾ���������";�q�>�A�>�?��O]_=T�!���>Z܎>�T�>��z>�h>�>�ȃ>��F� �/���Z?�}>=�=Za?�-[>�������>�V��D�u��ޏ�½. U>�7�=Һ�>k!��9��>S�ֿ�[�?�ߗ=�U~��j"?����ʤ�=y+z�B��F���77?�0?�>�>Z�L>ߗK>�'�>^�>�R�>L&о��>-��� ���@�qP�J�;^�z>|ɗ�ڎ+����^n�uE�M���cX�l�k�;����<�)+�<���?0���j��L)�I3����?,��><�4?�h������>�u�>?(�>ƃ��򸕿I� ���?x��?bc>X��>��V?W�?�0���2�~Z��zu��@�Q�c�|1`�����c���c-�۬��ɳ_?�By?3M@?���<dKz>uV�?#&������:�>�H.���9��T1=�>�ܯ�D2b��;ԾCd¾c��LC>';n?k�?��?βU�f��<?%>>f>?�M8?��?~6-?�7]?B��� ?�>6��>�4�>e[;?0S9?b��>\�[���P=��Q���?1|�^u�A���|�8����:=��#=�j��C=�<�5j�n+>�o
��"�T�̽����A��=O�=���=N�>�W?�c�>=O>r1?���Z0�l���[/?�ޒ=�y�E4����`��~%>�Td?¡�?�(<?F>��a&�dV�=���>�*%>�g>�a�>n�$��]�]��=OϢ=B��=�r>���;2Җ�~ ��q��!P=�>��>�t�>��H�˙+>�t����h�m>=8L������e�)E�%'2�+�k����>,�K?[�?��=v�����e?a��#?n+6?�H?N��?lؼ=�߾|�9��CB�F� ����>X�<�������V���u=��ʡ<&�l>	���^Ƞ�T_b>���a޾ϋn�6�I���羁M=�r� �U=1���վ�<�{L�=�S
>����� �e���̪��(J?�yj=�j��1tU�6^���>���>�ۮ>#�:��Aw�:u@�ޡ��pv�=���>h�:>�����~vG�+�E�>�bE?i_?]M�?�U��|r��RB�����rڢ��hż	?E��>��?3�B>���=/ձ�˼���d�Z�F����>��>���G�񀞾��󾮃$�i�>q7?�� >c?��R?wT
?rN`?�)?n�?QM�>ذ��蜹���#?X2?��<��PP��F#��C;���>��'?}>r��g�>#?]?�D?o�J?\?"?�[�=����,�+*�>�_�>�-S������-�>�?L?	Cr>K�^?`dz?��>�'��/����<7�>���=R(?!$?�K?G�>�z�>�����=�f�>��b?���?�o?���=��?��1>�D�>�q�=4�>��>�D?�IO?C�s?v�J?D��>]+�<���JJ��j�r�\�J�QB�;�N<,*z=�����t��Y��<���;�F���%��H�VE��\���_�;���>;5>$>߾��@?_���J���������;½z1ǽa����B>48g<�?y�n>Mw�>3�Ԡ?"�g���%��7?�,?9�A?���c墿>	������sA?/Ǥ?&V��/�S�����R�뽀>�1s?q˭?�t��I�L���b?�]?5g�z=���þ�b�{�龏�O?��
?��G���>R�~?��q?޸�>U�e��:n���0Cb�q�j��ж=�q�>�W�?�d��=�>�7?(O�>�b>�'�=�q۾��w�:o�� ?	�?��?���?z+*>��n��3����o��8-`?� �>�I��rC&?�һ�ξ冾��{��잤�0�����2'�S��+�Ƚ���=1N?,�s?�p?fb?�� �Pc��cW��?��JXV���uy��C�s@�C�A��o� ,�a(��8��P�*=\*O��+`��̾?�w?��>��/?K^���׾�h���lO>�6�d06�8*Q>O��&���4;qk��U����K���?�z�>�N�>�-\?��K�I�0��Ѿk$Y��C ��8>��>��>ו?�Hc�+����翽��Ǿ(�Ͼ'���<v>�wc?(�K?Šn?�� ��1��r����!�d�0��/����B>K�>�Љ>�W�����J&��I>�
�r����L|��6�	���=�2?�#�>͵�>�;�?��?��	����#y���1���<&��>'i?�m�>��>�Ͻ�� ��m�>�I�?�M$?L	h>-9;�.Ⱦ�f!��2����>oq?Y�A?���>/أ<o�`�\Қ��a���q8��6�=��v?�Z���ؚ��>�?��=X2�=��>����g	�>]���t�IG�>r�>�Bֽ~}>كþ% �F�^��y?�a�!?KG?Ao_�ں1�2��>̏?��?cʬ>�W]?��>5����[��?LFM?$�]?��e?�~�>��y?�:6�ٽ�[����"�UA>k��>�'�=T",��jw�񽎘G�Ώ/=�b�<`@7�a�c���=��t�q�$��_s��e+>��߿QbW���׾wJ��q�:��M{��0���о���V�F��xվ�ӭ���F��Fl�2KO����~܋�M@�w�?@����>>F��tZ��&���IE�>�˼�;F��h$����i����σ�t�y�<]�a�6�9D�إ��8�'?в��T�ǿ3����$ܾu  ?4 ?Y�y?G�B�"�Q�8�P� >J��<����y�������οD�����^?��>3�G���>���>,�X>P<q>����瞾�R�<��?N|-?��>ͅr�	�ɿ����ㅤ<���?��@��@?	&���辇`=;��>�t	?ߑ:>Z�4���f��A�>Zy�?�׊?Q�X=��X�#5�U@b?�&<9�C�`�ݻ��=���=)=�/	���H>�>�$��e?��ͽ��<>�]�>ֈF��z�Y{[�LK<�
`>��׽�����τ?�X\�|�e�d�/�BH��Bi>��T? �>�Ġ=ҕ,?8OH��ϿP�\�u1a?�1�?b��?��(?�޿���>O�ܾH�M?�16?x�>�J&���t�f��='�A�����?V�W��=��>\�>2!,�����O��̚�@�=����˿>&��X=�������q�*Z��ն�Fy�k��� Tj��>h��Ž�һz5�=O�x>���>6�=��~>g#a?��q?���>�BN>���&!��)ᗾ���:����g�彸�]�-2��ꪮ�����j
�j �=��x��F�Ӿ]?�ƪo=�,R�����и&��<g�2t?�Ο-?$4>��ž�IH���.�?OҾ9J��n���uq��i0ƾ3-5���n���?ǯ@?f䉿�J��\�8|��ƽT�Y?�ǽ����=��N�>!m�~�=ߚ�>zS�=��׾�	"�m_L���?�d�>پ�z���r�=+H���N���A?w\?�XM�U�>�>�)��D`׾��^>���>47=>{�=>������r�
?u�.?��ѽ7�F�(��>o@�����3��=e�>�	���~W�hF�=J>�<w���j佯�A�����1?.��=p�.�l�;��;95��L�v��?FT�>#�=w�4?��<?%���Fؕ�}B*�@������Qi?=g?��>>��G�0�y�� �m�y?'r~?��4=�9׽@SR���V��w��5?�z�?�V�>;�<Zs]������`�?��v?yr^�Hs�����2�V��;�>\�>���>��9��l�>.�>??#��G��Ⱥ��=Y4��?x�@s��?m�;<1#�Û�=�;?8\�>a�O��?ƾ�z�������q=#�>���aev����cQ,�I�8?ՠ�?R��>e������>{3��޻?���?����RB>Qv̾��c�����<=b�!�M�X*�>�x��Yq�Y�����]⎾��>r>ެ@Nn���;�>���<"Oڿ�U���%Z���Y����w?ђS>,��9�����h���/�e���^$�^yνҪG>4�>]zL�	.�����8�V�j,�<,%�>�=r��>n��T���xQ�m#>���> �?���>\�H={!;�,�?��־a��1������F?L�?���?��>weݾ�?���=�C�=�l?b5?y_H?3����>�Z�>(�j?�V��M`���4�L=E�1U>�3?|?�>ݎ-�u�|=_(>?U�>|j>%/�!�Ŀ�Զ�����{��?e�?�o�h��>���?�z+?�k�b3���M���*��'J��BA?��1>����9�!��=�/咾:�
?7z0?���{3���_?�ra���p���-��vƽ=ߡ>��/��L\�65�����qe��	����x��?�^�?C�?M�C�"�g8%?ί>㈕�b7Ǿ�s�<;��>��>��M>�`���u>�
���:�10	>	��?Xn�?�{?����樂^>��}?�5�>��?�0�=4P�>h��=���\�7�b'#>��=p�A�μ?��M?AE�>O��=�9�o1/���F��R�l�4�C���>�a?��L?Fra>ù��/�.!!���̽�g0������?�_/�ߌ޽�05>��=>��>�>E���Ҿ��?0p�+�ؿ�i��go'��54?���>	�?�����t�n���;_?vz�>�6��+���%��=C�a��?�G�?A�?��׾"U̼5>-�>�I�>Z�ԽZ���T�����7>;�B?���D��[�o�G�>���?��@�ծ?Xi��	?���P��Oa~����7�l��=��7?�0�*�z>���>��=�nv�ݻ��V�s����>�B�?�{�?��>�l?��o�M�B���1=5M�>ɜk?�s?.Oo���o�B>��?"������L��f?
�
@u@a�^?*�2�������ξ����4t=CĊ=b�9>Lؽ�f=v9"=+pO���<u�=#!�>��4>6OK>cXf>��=�Q�=c
��,��0J��.U����@�"G�<��<J@�h�I�p�I��T3���e�� �����0��j�Nu9���N��c��q�=CT?�}Q?[n?��?`6���5>������<� "����=)1�>�2?��N?\�)?�'F=�>��%�f��������և��u�>��;>�C�>A��>��>��0��RX>�TK>ćx>�>u�=��C�;V+=��Y>��>	��>��>�H<>0�>˴�	+����h��w�L+̽L��?�p���J�T*��)������GZ�=d`.?Ⱥ>Z��`9п@ﭿ�,H?F���� �r�+�T>�0?�XW?�>�����U�pU>ӫ�+Tj��Y>G �Yl���)��Q>Gt?�Yg>�Ou>�`3��8�vP����a�{>��5?�*���G9��u��[H�t[ݾ�KK>���>��.�v)��ؖ���~��i��{=�|:?gV?�ಽJT���u�b:��iWQ>��[>y�=Ը�=�AM>��`�1kǽ�G�P�,=ȿ�=�^>��?��a>�|%=E�>�`���f�b��>�<.>Uvb>~�&??zV�%pB��U��4ܭ��Z�>�F�>��=�R�=�-n� ɺ=^�>T>�]E�O-x�����G�B+>�9ȼ��d�W�G��=3=��p����=GVj=d3ǽ\��{=�~?���(䈿��+e���lD?O+?� �=P�F<��"�B ���H��E�?r�@m�?��	��V�D�?�@�?��=��=}�>�֫>�ξ�L��?��ŽDǢ�˔	�!)#�iS�?��?��/�Wʋ�>l�e6>�^%?�Ӿ�=�>.	!��|��^���#}��n:<>��>��L?����(���4�;��M?�y�>h۾Of��*�Ŀʆs�8��>k�?k�?�+n�@����@�y ?���?�oO?�Kv>۷�wM~���>D-H?��Y?�?�>�)���6�Ȏ?�^�??��?A�Q>�n�?�y?�)�>�O`��* �*����$����<m�f=Uһ>[�=,M��xh:��~�� \��xlT�����j�>��<�D�>A��'�����=Z2j������z�_b�>�V�>N{i>5��>���>]��>�p�>ŧ��ἽO�k�������K?L��?[��2n�}�<���=_�^�H"?�G4?��\���Ͼ�֨>��\?���?��Z?�^�>���38���㿿�r���g�<9�K>�2�>wL�>�1��- K>��Ծg0D�u�>�Η>���c?ھ�(��r���&.�>�_!?���>��=�� ?��#?�Sk>?.�>4*E����S�E��D�>:�>�M?��~?[�?5M��h:3�y!���ҡ�oV[��!N>�y?"9?*�>���w��6;�8�H�e�����?%bg?����8?""�?w0??R�A?u�e>m����׾�I��Au�>+m?T���/�'��*A���>�4?��>�]<ɤG�)�Թ�ԾD�݇�>\�f?^-8?��վ�^�[���M�<�����`?��e�E�)=�'>�Y�=��~��R�=�~=�}}=y�b�($���0�<��=�V�>�@g=U$'���L��D,?�E�7���=ʩr��hD��w>$L>`���w�^?�L=�Q|�l���h��/�U���?���?�I�?�ﵽݫh�=?�7�?�?O��>.7��܀޾י�X^w��x�Tx��>ԝ�>;wg���侘x��m|��{M���Ž#���z�?�z�>oj?�*?@~>^u�>����&�p̾��ھ�e\�r�����"�:�7�+)�O!��A�5���<�a���Ag�02�>}�����>G�?��j>�R~>���>��<Z�>�!n>�0L>�(�>�n>|e�=iЅ=Ef�:n:���z5?]����0�f̾Q���>R"?3a2?`(?�e��p8������o8?I(�?�T�?�3a>�Ol�+�[��?�p�>�zU����>�ܚ=�9���.>�<����*��g-�6�#n�>
�W������3���o���
?i��>�Щ�{N���6Z��m����p={T�?�(?��)�n�Q��o�ʸW�S����m�g��{��i�$���p�]���5P�����(���,=8x*?�!�?��;�٬�[k�=
?�.+f>f��>�>�>�D�>`TI>6�	���1���]��]'��}���L�>�5{?=s�>�NF?$<H?�G<?��f?��>�:�> �>�>:�<h�_>Q�>=?�z?�i7?�B	?��?�:V>��>�M�]4�PQ�>�?,?�z�>��?���]<�{�N�=�)�F�ν��<#܌��94�6W���=��/>�?!��J�,�����=�>��+?h��>$��>fͿ��-� )�=	��>��?Kq�>�9ƾ��k��<�庵>��5?uU��ȁ�<��	>�,7>zb<�Q�l�}<�4ν�)�=�@=��A=�� �q��=Q�=���<����?P��Yq<�Z��~�>5�?��>dm�>�I���� �������=�wY>|rS>ٿ>5Fپ�|��1����g��ay>6z�?�z�?�:e=���=�K�=ep���Y��k��EｾjI�<%�?�9#?KT?ƒ�?�=?�^#?A�>��P@��7S�����	�?�f,? Z�>2���Ⱦ���2��T?�0?Ϟ`�a����'��ZȾF}ս�,>�0��|����`D����h���1���K�?���?�ZV�e�5��6辏}���7��=C? T�>G-�>p�>$�'�~�f�]#��p<>/X�><�Q?�>n]Q?P�?�P?��>;!�##��v]��i6���U;>��0?�bj?���?�jj?���>V7>����7��>%��D@b�D'���㤾MK=�6Z>\��>�J�>#\�>Y�>������h=;�C�v<��^>-v�>�u�>�>	3G>���ZCB?G��>�ƹ�5?^��]��AC)��#i��
b?銥?,g?
J۽�����j���|����>���?؄�?w�_?>d���">� �l�i������>�]?
?=�>�I�XD���>��>;�
=q�����*�F*��$��>��>t��>���(��{���� ���x���s��/4��;��T���/=T��Y':�
��I��K�徳���b���#<׾qă�B�>��v<���=}�=��4��e�;&�=377=�ޞ=��=�d�<`�O=K1x���ٽ(���Ỽ�d���j`>i��=�Y˾�x}?�I?�}+?֌C?&�y>�>��2�P��>;���{Q?8�V>�R�>�����:��_�������ؾ�׾�d�����@>/ I���>b�2>Q��=��<np�=s=�W�=�N�Az=wl�=(Q�=�ƫ=���=]�>>�6w?8���첝��4Q�'Z罙�:?V9�>�{�=��ƾF@?_�>>�2������Gb�
.?���?�T�?%�?�si��d�>%��䎽�p�=淜��=2>���=y�2�[��>��J>���K������s4�?��@��??�ዿ��Ͽ'a/>�e>��=�hG�� ���*�İ�|�о4�!?UQ��\S5�릖>���>�<���H����>d��>�C��0@���2R�=|��N׽��#<#��>*�{>ތ��ᵸ;���=���;>C�A���k=$=���N�0d�,��9�?3>n�=�C�>W�?��?��g?+�>�;��R�پ�j��c(>ܘ�>��'>�"��6��=І�>�j&?�gC?�,a?���>˘x���><��>D�Z��e�/��ځ����>E@�?��p?�>2��PXҾx��l���DϽ�4? %?�;�>~��=�d������7�:�u�桁���/�F� >���Z��D톽�N���d;�k�<F�=���>:6E>�3>�8>��=oU�>Z�=ˣ]=��?���ؽT������۽e�I��Y�%Խ"!���W=Y9�=L��=T�>���<Ey���<���=i��>C� >���>N�=�A����(>� �K�9��=�T���IE��c��t|�ܨ/���5�mwC>iH>`��0��:� ?�to>��<>!��?��t?�>n�
�}Ѿ�r���wj� `D����=��>E�4��n;�*^��L��tǾ���>	F�>Z_�>�-l>�X̾9j�6��=N����4�W�?���V-�"���0)Y��2���a����5������(?撈�	�<�_�?�10?sX?d�>�>�������v*���8������|$>�h�r>'�%?�+?|�?[�׾vR��R�׾ ׽
��>mU"���Y�嘿Li%���;�����~�>؜����ܾN�7�<ԁ�=s��C<;�=_`�y�>��??�Ӹ?z�N�i����E<���"����s��>��j?ӳ>���>f��>֎ּ&��a0����=�}p?SP�?���?Ԏ#>O~	>S� =t�?c%>f�?�ʚ?�s�?^۾��=��(>SF�<F�<��S�>u;�>�)=bʾb�}>;��9v�?�����.��x��۾>\��NMJ�
�X(m>D��>XB>l�e�L*�>Z���e=Ľ�5�>+?�>��1>nTl>H��>�4W����`?��<L�$>YN? 4<=�=�J��'�2>jL������0�c1G�f�I��x�w^�;F��=�C>m��<�7ֿq��?=��:|����%O?���|`�=hߚ>�Og���ȾL�?S��>G3#>z^�>�}�>�e<$h?K3�>�4Ѿ�>��
������C�p{Q��CҾk�y>т���!�']�x� �q/L�j⳾mP���h����ϳ<�I��<�M�? �	��7h� �*�i��8d
?�G�>��6?�c�������
>�:�>��>����c��7[��O���?v��?�c>�G�>�W?�?ϻ0��G3��MZ���u�`A��ud�̯`�մ��.a��-E
��Ӿ���_?��x?]lA?�%�<��y>�z�?��%�����b��>Y/���:�C>=�K�>�ɰ���`�.�Ӿ��þCR��F>��o?)�?	?{�V�Ld�R�> �9?'�.?0qt?a3?d=?����#?D�4>�?�"?=�3?�-?�	?�0&>�_�=����F4=���E���vؽ@��	�3(=��n=w�s����;ܿ=7E�<������eP�m���ݣ<�)D=���=�D�=�L�>�hW?uG�>��>�??�����d꿾b*3?[]]>�P��摋���oT־!{)>��S?�!�?�qa?�>XJ�nD���='�O>�>fp*>`؝>��r�!z'����=Z�d>P�>I��<��;�\���3;��E��0:<FBr=���>Eξ>�z="H�=��佀��;��>	��w4����_�5[���W�����Д�>�8d?�&?��\>����b�=;�_�Dp�>�c#?�R?vہ?n�p=��3�O��#�!��<�W�>�T,>!��T���
��D�f�>���V�M>)���k2�`%+>� ����ߡb�B!!�c��vp>�=�s
=m���'y�I>~�D{=,��>[�
�M�$�mc���e��q�:?PI<�2AݾMR�ZI:�'�=+��>4�6>���%����4R�6�+�I��=���>�Q�<�&�������,����K��>A�B?�Z?���?���]q�oKC��|����$t��?`��> �?.kH>%�=r��oA��;b���E���>�M�>����C�&����.���0����>��?��>_�?D{U?l�?�\?'?�,?��>kY��B𺾬:&?|��?�{�=���FE���:��J����>(?X{@��Ǘ>G�?�?�#?�-T?a?�=#>v+��(�9���>�j�> l[��1����o>�M?nt�>KX? ��?Yu>˾4�����5'e��y�=��'>�5.?�o?��?8��>|��>�V��8�=�L�>#^^?��?{�n?���=��?׶>�G�>�Đ=��>i�>Q�?��N?��m?�N?j`�>�a�<|��yƽ\�l�*!�E�߻#7�;��=������Y���\��<v[;nD����A�p�m�9������=��z�>�ԍ>/���>��E�4��=��>t� ����Q����c��y�>�M�>�)?/��>9�b���>Z*r>�L�>��8��~?�2*?p�$?�5q���T�KsN�y<��{�$?p�?:<>u�h������凿!����?��O?�}���в���b?��]?�'�%�<��Gľ�b�x����O?��
?��G�I�>�~?t�q?��>�{d��n�g���Yb���j����=*�>�J�}�d��6�>�7?�B�>��b>�r�=:K۾kx�d!��a�?>�?���?�Ԋ?��(>��n��࿿��[W����^?H�>�㥾�#?� λ��Ͼ1���D���B⾖K���R��kH���=���k#��m���Tս��=�?�Mt?3�p?�:`?��r�c�r�^��9����V�ւ�Q(��E�A$D��ZC��o�A:�$���(���jG=��j�D�_�-׸?�(�>��<��>�#	�� Ѿ9�:����>�Eþ���<ke=.�I����=5��=%���������d��H!?�o?���>dL?N�f�>O%�T:�AB��#)�l�>�g�>08�>` ?�t�����'�������M�tܽ��v>�+c?�XK?*�n?����0������*!��,�64��.wC>i�	>xɉ>!eW���� �%��K>���r�ѧ��:��8�	���}=�12?�2�>w}�>��?D�?�q	��6����z�u+1�c̆<�|�>�Hi?���>ӱ�>Hս�� ���>��l?C��>��>�����W!�"�{�\|ʽ,#�>�ޭ>���>��o>��,�\�qf������9�(o�=i�h?���t�`�ޅ>�R?�Ê:S^H<�q�>W�v�W�!�����'���>�}?k��=��;>�yž�&�l�{�?1��.(?Q?1���+)�sbo>J�?$G�>{��>ή�?t)�>N{��w?�z�?'B_?oIG?�s??���>�Y=jo��Io˽�i#�d�=ĸ�>�`>�Q=���=���|P�h�$�i�$=+��=(���F���d�;_�Ƽ�o�;�h=$/>Q��^�ߤ�g
9���m?�{���K��ph��lڽ�Zо殓���R��:������|=���b������艾��?%W@z���7ō�p�����R��l���?Bp��\���^��5��n�9W �ε���95�Tc��♿Ϗ�	�'?������ǿ�����:ܾo  ?�@ ?K�y?�m�"�f�8�ө >�D�<������6�����οR�����^?W��>�
�]6�����>���>W�X>vKq>t��K螾a�<x�?ڇ-?X��>�r��ɿ�����ˤ<���?��@�MA?4�!�s���x=?��>Q]?�QB>=�2�~4��m��D��>*��?�E�?6.�=�N�Z���)�\?+��;�kB���<�o�=��= y=Ԃ�:�c>��>�7�ȵK�it��! #>��>���f��e�����\>�����Ny�4Մ?{\�tf���/��T��+U>��T?�*�>�:�=��,?`7H�V}Ͽ	�\��*a?�0�?��?��(?Vۿ��ؚ>��ܾ|�M?UD6?���>�d&��t�p��=�8Ἑ�������&V�Y��=%��>؄>�,�Ӌ�y�O�H��U��=�����_�0��:D�~���f�{��cd�D��;�GI���p��P�=�J>�%>r)^���>�'�>EbG>P>%>��a?%@W?��>Jr�=$�<���	�	���
竽��W��wk��e-��0�#m���n������n˾.�Eپ0����C��m�=I�#�����(���5��>��e?�������H?��Ee�f۾J��`�V7o�-�˾w4U���r�G�?��>?�6��h�� !��ӽ$��d�I?�\���������=E<O�>��>�5;<����ƍ
��8���!?�r?������3����w��q��=�8?���>�]="�?��>V�2����<�z�=�5�=$�>�_�>Eh�=����A�뽮��>��*?��X��Ǣ�A��>�����>�-�>�D">O)(�u5��s�>��g=�o��1Ͱ=^�=w�;b3U?eD�>k��X�^�W�QJ����tYo?���>p�k>KRb?:b=?v;�=&@׾*+7�H�9~�=��R?�1b?�+>����Fs⾄0��R??�3w?궁>�Mn�Fn��;�;�q. ���?/
�?p�+?YN�>[��e��������"?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������1�q=�"�>���ev����R,�f�8?ݠ�?���>��������=�ˍ����?>�t?��&���=�1��cs�
���}>-N�=�Y>���=��ݾ9�*��n��E���苾���=�>�v"@0E��Ә�>_�n���п��Ϳ�璿ߗ��g�پ��)?sX&>�e�H���,�=���M������?���4��>`��=�Rs�Ml��(a��A1����;��>FUL<P��>*א�P��������<W��>�5�>9�[>k����c�?�� ��ȿ�b�������R?�E�?*��?n�2?��Y��X��.���=��G?OKs?��\?%ǼC�0��b�"�j?�_��tU`��4�uHE��U>�"3?�B�>M�-���|=�>z��>g>�#/�t�Ŀ�ٶ�5���[��?߉�?�o���>n��?ts+?�i�8���[����*�T�+��<A?�2>���=�!�B0=�OҒ���
?V~0?{�g.���[?��.��?S�#�1�r�A=�ט>S����.���$��C��{+K�!��������?I?�?И�?^��u���T ?�ҩ>5��^��;.�=���>!H?[�>����p��=7���/�iO�>��?+�?��>Kծ�M���h�>U|I?=%�>� �?��=��>_��=ݰ�1%��r#>e�=��@���?ʀM?���>���=��9���.� 4F���Q�J%��C�U�>��a?�;L?1Wb>�踽1=3�t!��̽A�1����i&@�.�-���K�4>��=>O>�sE���Ҿ�?t�F�ؿki��Rl'�V04?E��>��?J����t�~���=_?A��>�4��,���$��o;����?bE�?0�?��׾�e̼n>-�>1Q�>��ԽP��������7>��B?��C����o��
�>h��?)�@�ծ?i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*�V��ぺ�	�޾V�}46=��<�)H>`���5��=aսc��}�<�.]>Z�>�+@<��~>�K>�E>�l4>���A2�,珿�6���<D������L�����Vu<��$
��$t��<���:���淽��ӽc�K��8i�Z=
�=��=l�U?pR?�p?� ?��w�w�>S���:j=Ʌ#�,ل=�)�>xd2?n�L?��*?�ϓ=ؚ��?�d��Z��SA���Ň�iy�>CgI>�y�>�:�>k1�>�G9��I>#3?>iy�>k� >��&=�C�?@=�N>PO�>H��>�r�>�a:>^�>״��=���g����a̽�Ȣ?^���IK������`��(޺��=�Q/?(O�=J}��s�ο�j��SG?��������%��K>KE+?�T?�>뒲�7s���>�	��Li���>>I���p���(���M>�?v�s>���=�b5�`c&�������"�OcC?�� ��-w=>�c��w��� �"=>M>�;�nI�'������r�j �-�=?k3�>c������̋�("� �G>Lb�>��2�W)�<�[>(6�:݌����=nz�=�>�p�>�	?��P>Iؽ`�>��"��'��%�>��	?o�=# +?�oW?%D���6���=��Ž4f�=G��>��>���=�(�ԼB"�>�P7>��G�����J�W��r]���=����]�����

>v��/I�>�	�=����JS�I>�z?�����P|���׾8�=|�S?X5?�Qe=��A��,J�"Ҙ���t�)�?<!@��?����L���?�?�Ȇ�.��:���>��>�ᐾ[�仨�?3�?�6�¾�����J�m�?�5�?���=a\���ό�8�=v ?�Ͼ=f�>�y��W������u��j#=��>�:H?a_���N�O>��f
?�?H� ���[�ȿ�yv�L��>S��?]�?��m�@B��S@��k�>?��?VmY?nIi>�_۾�Z�8��>��@?
R?-�>�:��s'��?��?ڦ�?yI>J��?��s?5h�>�)x��W/�e5��<���v=c�\;ka�>�Q>����neF�\֓�'f��h�j�H����a>?�$=.�>�I�2���8�=;�I��)�f�_��>g,q>��I>R�>�� ?Ma�>ꪙ>��=PN��#߀�'����K?���?���{'n��ѿ<1Ϝ=��^�z%?dH4?�\��Ͼ�è>��\?��?
[?o]�>=���=��㿿Cw���y�<?�K>��>vF�>k��biK>&�Ծ�"D��X�>�>Č���Jھ*=���&��r=�>9b!?���>�i�=�@ ?��"?v g>4��>�E�$쑿�F�@��>���><�?t�}?NA?������1��)����� W[��M>�cw?u�?�{�><���镜�Ub{���T�����T��?v�f?���E?���?`!A?�8@?��b>��Y־������}>�:#?�����.��e	�:΁� 	?Q�>݊�>�)��ws��ڽ��$�q��?`y^?Ҵ?����k�0���}(=�3�t�������<<K�=��|>(����=dw{=x�Z���꽅�|��Q׼��߻�-�>}�=͙ڽKJ.�(=,?=�G��ڃ�d�=��r��wD���>JL>���I�^?)i=� �{�A��\x��U�� �?���?,k�?�	��Ɲh�$$=?��?S	?�!�>J���~޾g�ྌPw�$�x��w��>���>ͩl���ˏ��晪��F����ŽT��>��>��?j� ?cN>Y��>����g$��v��K�[�&�$N7��(.����Ǣ��� �D���_ľ �&s�>v�����>]d
?��n>�x�>@2�>��ۻ�,�>/�H>�F�>ğ�>��\>�.;>@�>�\X<WEý)�Q?����k���i��:ܒ�
io?��^?�[�>+�5��������0]E?��?R��?�g�>�e�����f�>X��>[Ú��	�>�07>���=�
���e�H���W)��kѼ�>Ѫ0��i�L�_��͎����>Jz
?���=W��;=�?����q=`;�?��%?�*��eP��)n�k!W�uS� �*� �k��ץ�e^%��Xq�0
�������ǃ��*��=��,?�?�<���ғ���"h���?�"i>���>��>-��>8D>�	�w�/�`/Z�N�&�fv���z�>�h{?�J�>��J?��N? s?��P?���>[?��ѾK)?�u&��x�>��?sS?6�#?x�*?�?�)?���>#�X=VW�ľ�/?�?u�?X4�>�?�X=���=���=f*ľ�T����9k��z =��T���<�N�=��	?���:s�,�n�Ͼ�m�;���>Y:�>���>��]�X���(cJ>E��>܈?��>��������/d�>g1/?�V�O�I;��=By
=ST=�H�=��_��J�u~>*�׽oͽ=�H=�1=��o����:֏7���y=A����B�u�>��?���>�C�>:A��� �ܵ��j�=Y>�S>>MEپD}��X$���g��\y>�w�?\z�?�f=Q�=T��=�|���T������������<��?VI#?�WT?ꕒ?��=?j#?r�>*�M��F^�����Ǯ?�b-?OPU>1%;Q����䚿�X'��~�>hc�>�~T�i�Ͻ��T���T��@5�����OQ��Pr��b��mHB����:+��$���?A�?dq>�>�l1�g���'��p�d?���>���>vQ�>���b����&�Y6�=��>��U?��>�Q?w�{?��Y?Rvd>�4��7�����:�b<�>ɵ<?6ƀ?�e�?�~s?@P�>��'>�|%�Ztܾ<��j},�I���������9=��\>|�>&�>}̝>/�=ܰ��fȲ���D�ox}=��X>
��>�g�>/��>�A�>��#=�\B?��>V��TR
�Pי�r�����S�p?'�?�82?Ԭ=y���I9���j��>���?7��?s ?��H��� >�_^��ھ�sh���>8��>�֤>8IS=�-=1�1=��>'��>���
��E/���-�E� ?��K?�=-=�@ȿ�y�4��&����<�������`���g��K�=.5��!�Ƚx���B��¾%x��y[�����k�{��?�=��=��=P�F<���<�c�=�vI�Fܼ�S=Ε��K##=h��d���	�f�<{�<��=j�麜�����y?R�B?)?�s<?u3x>$>��ɼ���>�v�ʟ?W}L>���I����T@��U��oË�t�׾
վ�we�6���x> �B���>��+>f
�=�#7<�X�=��f=B/�=;���\��<�,�=}5�=.Ӥ=Pc�=�(>��>�6w?K�������4Q�=Z罎�:?�8�>l{�={�ƾf@?��>>�2������vb� .?���?�T�?:�?ti��d�>D��,䎽5q�=÷��+>2>��=O�2�G��>?�J>����J������|4�?��@��??�ዿƢϿa/>�{:>^	>�Vr����P�ؾ7sþ���~�?�;�ϳ;��>S��Oֽ��ʾI*�h& �����=�nvu����=��ͽ�������;�k>�4
����=C�̼R$�<zJH�ʍJ>;>|�ܽPou;��I>��۽�"=<�=�鶽ޓ�>�E?`�a?Y�F?��?���+[㾡<�8��>zB>:��>ܭ>��>;]�>�G^?�D�?�ft?���>o�>��>j%�>+Hj�_�}�q����	�6���,k`?�
M?.�>���<��L.8��*�C�?>�w??�n?)�>��(>>)�&���&�v_4�����ܺh�1=�Vl�S:2��W�9f(��ǽ��=a��>��>�|�>9u>�31>��H>o�>�<	>��8=0��=\�(����;�5�U9�=߿�;kt=I]���+;V�����'m�;�v���]���ی�.~�����=���>�L>y��>�|�=���s4/>;���7�L�kͿ=�D���'B��/d��C~���.��U6���B>95X>�i��l2��}�?|�Y>�Q?>��?ZAu?��>��Y�վ�N���[e�tTS�8޸=��>��<�@s;�
Z`���M�oҾz׾>�4�=V�?ߗ�>��̾��-�KR��0���$��R?
���5w>p���VLm�򹖿����i�{�HS6�\�!? ���%~�{/�?��@?���?�1�>(�=�C����>!�[�,Û����F��.w�=&?b?��?�Q�>���VI��{m��>"Р�RR��؀��C2�EL����̾7��>u��s��<��r���Պ�E-J� ��(�>+?+$�?��(������>�E'��ݰ:J/�>��o?&��>�}?��?�k[��̾��6�M�^>��a?I��?qZ�?��p>,L�=�E�	�)?��,?:u�?�I�?M�?Ѩ]�8�d?����SPH�n~�=��
�E�4=(�>��>��?�X?X�!?��%�����Ѿ��.������5>M��=�?�O�>��>"��>=0�̻>NE>=��W>I�>Xՙ>*<�>4�w>2��� �9?���=���>Pm+?��>��<�7�=vt�=��'�E>Ž�WQ���Djq�<�=����:�=x�<�3�>��¿Z�?'q�=�b���?%վA_=�@[>�t>y;���>��v>O_}>��>�>t�>u>�7>�߾g>��
�<e(�g�C���H�"
ξ�ye>����(3�q!	��2��ae���Ǿ�S
��m�����D����呓?@3����h��$��`���
?��>�6?�쉾~ �<�5>V�>�c�>���̉��)��׬վ�1�?�?�ec>���>|�W?�v?h&0�tS3�!xZ���u�-�@�x�d�Y]`�x���k���l
��;����_?}�x?�3A?�-�<'z>���?S&����^J�>n�.��9;��9=l�>B)����`�n�Ӿ��þ����uH>��o?�>�?XQ?LU��Hk�|�%>��:?671?��s?7�1?�Q;?W�A�$? ?4>r�?GG?u5?I.?�
?[�2>a��=�9��o�/=����1+��^нK�̽�����P.=�Q|=���9$i�;$!=+�<l���
׼|I;����=�<Ȍ9=C =1��=m7�>(�x?�R5?%߼>T�[?��3�94,���+�=y@?��=�C\��S뼄�x���'�D�>챚??�?�h�?�r@?���u?�cg�>[�>1�=%�D>l޼>]d�<�ʾdo0�� d=��>�e>��">�T���b	�ǵ�>��'>�?�W>5G�pd�=;���kYQ��_�>A�5������I��8�[�P~�ԓ���>�M?rK?�홼[���$� ��`�_�?�XL?�6?�G�?r ��j�	E�QkT��b۽��;>�P=>�l��>�w]����5�^g�>,�������y�>K�վ�s��jg�1�N�"�As�>��]�w�x�`f�8����|��벽;6' �P�Rr��Zɋ�]fs?�7Ľ�{���ĺ�(���:}Ħ=���>i���
���P�R�?">�>#?;>v~�=N3�l�6�6�#�tGk>�J?� `?,�?�>%�z�d� iF�N�h�p���R�^F
?���><?Ԯ9>"�E>#�;�R	��_@��8� �>3/?�]$��P�F����-����QT>�?���=���>�<?�z"?_Sl?�N/?ߎ�>�J�>�;����þ�P?,҈?�w�=]6�$��;�+���G��6�>|-?H���TS�>�o?��? �?��a?���>tcj>����%�4�>n�>pp��@����>aR?�3�>l�9?�~?�\�=�:�=ْ���.�9B�=~�;'�3? Y?p�?-��>kȥ>޸;��=�)�>�2L?�$w?�-�?U>��
?
ٔ=��>�6��jֻ>�2�>V�?[Z?S�~?0P?��?�.�;��� �k���cCz���;;�C{=�(�<��5�f����D��A�<��>>Ec=} <'���ߚ��۟���ռ��>!w�>�E�Iު> ����O=��>��O��8D�_a�N��WoI>O�=;�'?�K�>q���E`>^+>�B�>�3���>��(?
5?M��;�����"������>�P?��>F��J{h�����+>�E�?λW?l�5�o��O�b?��]?�g�=�p�þ�b�[��t�O?��
?��G�4�>>�~?��q?L��>��e�P9n�,��+Db���j�&ն=�q�>_X�r�d�m?�>��7?�N�>p�b>�%�=�u۾��w��q���?\�?��?���?�(*>A�n�W4�w�������
^?�)�>}�����"?�_�ξi���T���.ᾐ�4��;����b�$��e��\iٽD׽=�?��r?��p?ˍ_?B� ��\c�>�]�=���V�C5�+����D���D��@C�̐n��;�����$򙾏uB=;,����X����?�o)?Jj<L�?�d��2���"����>�O��o�����<�s��^d=��n�������R{����?Q��>�(�>?�3?V.X�F�.���8���H�Ҭ!�F��=�L�>˳>��>�>׽�Y2<T%2���	���E�n?��v>
nc?B�K?'�n?�l��1��|����!�'0�;u��=�B>��>[��>��W�,��71&�rM>�)�r���"t��S�	��7~=�2?�!�>.��>�G�?'�?�	��p��?�x��n1� �<g.�>a i?3�>Jˆ>�н�� ��L�>&�l?ls�>yԠ>β���R!���{��ɽ��>nޭ>о�>*p>Ŵ,�3\�.^��~��m�8��`�=�kh?M���K�`�0�>9�Q?v�7:#PE<á>�t�w�!�̮�Z>(�c�>؞?��=#<>_�ž�>��{�|쉾�?#��>����9�2��
W>�V?b?�P�>�o�?=ۇ>:2ž ��%?�f?5N?�:?93�>��=�U�<�'���Q1���<�f>�M>%]�=8>���"M��^Z�s0x�6%;=�U�����ܠ�<��!<��;<���<�U�=�)��~���D�����&��꫾�pb��X���ZV��B��D}���"�nf���5�=���Lƾ�Ka������,��~�@�$�?$<�b�����҆�{����>AT��)�(����~��G�4������`�1lW��Q��b#c��a'?yH��޷ǿM���}�پ7U!?Uz?)�x?���C�"�m�7�g~!>���<�&t�+�뾈����ο�#���^?��>��J᣽��>���>�[>b�r>�È�L��Ѡ�<I?1�-?���>�q�āɿ�`����<�2�?��@|�D?dJ�;�����X�-�?WSJ?)XD>Ņ�����ᾦ}�>nr�?�l�?�CL>��E����HN?��|�m�>���x�=We�=S�>���v��>;�>�����i�`0뽦�B>���>�����z(��5�ӽ6�I>U �xm�=5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�ޅ�=l6�����{���&V�}��=Z��>c�>��,������O��I��V��=3"���ƿ�$�,����=˙�%IY���56��U�T�N��J�o�$>�z�g=�|�=`�Q>䓆>�cW>UaZ>�W?L�k?��>��>��彵P���;*H��H��������A��Sv�����ྛ�	���^����ɾ�L=��ϔ=_�O�@ބ���*�$SX��@��&?��)=~����E��C���þ�:��jɓ�Aa!���׾�UH�oQk��&�?c�6?.Q����R�K������^�@(W?�J�����1��6�T=��9�ʻ>1[�>�A�=����J#���M��,?�??奾+����3�=�
��F7=��?���>�8�=@ء>�?�'��?�.�N>>0
P>@��>r��>���=�%�������?NDT?! ��CΝ��n>�b�x�˺���>>F}��r��sS>���=c���%����뽌��=�$W?��?�5&�wO�Z��<�Ո>�U��jA?7�? �>QJ?Q�I?O��<@!���u�yҾ?T�=�G<?!`?�>������w�U��Z?�+�?뼜>�ٿ��	�?[�����$?W�h?�tC?T}��:����� X3�l�0?��v?s^�ws�����O�V�e=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?��;< �T��=�;?j\�>��O��>ƾ�z������;�q=�"�>���~ev����R,�e�8?ܠ�?���>������rj�=�z����?���?j:����2=�]%�+q�OiƾP�=C��=5Q1>����K������f?�[��S�u�3m�>D@�7��V�>xYľsB߿��¿�,���֢��=྿�?��?N��=�������\� BO��a'�f����o�>���=R�ϼ�o��n���2�1A�5^�>S�w�=��>�q�����:����|����>#��>��s>�H�~S�����?w'���˿H������)W?⨛?A߁?��'?��D=ܫx�01��_=:��EN?Ա[?�zO?�љ��'�m־j?_^��]U`���4�_GE�pU>�"3?�A�>(�-�$�|=;>i��>�e>�"/��Ŀٶ�\������?N��?�o�P��>P��?�s+?�i��7���Z����*��+�=A?02>�����!�!0=��ђ�!�
?_~0?�{��-�U�_?��a��p�}�-�m�ƽ��>S�0�0h\�^���	���Te�����<y�!�?�\�??�?Я���"��6%?��>�����AǾ�F�<��>A�>�4N>�_��u>���:��w	>��?�~�?�`?v�������6>2�}?�*�>V�?���=�F�>�G�=�氾��.��]#>F��=?�?��?^�M?��>b��=��8��/��WF��>R�]$���C�e��>��a?��L?�Kb>�%��D�2�� !��ͽ>1�"~꼂�?��,�S�߽I75>c�=>/>�E�u�Ҿi�?%p�}�ؿ�j��Fp'�x44?u��>4�?9��*�t��o�4_?[l�>�1��,��`%���S�+��?�B�?p�?\�׾�F̼��>���>5H�>��Խ$��������7>&�B?��LD����o���>��?��@�֮?�i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?oQo���i�B>��?"������L��f?�
@u@a�^?*�hֿ����YN��Q������=���=�2>�ٽ<_�=��7=��8�v=����=i�>��d>-q>=(O>�a;>��)>���O�!�	r��[���P�C�������Z�C��Xv�Wz��3�������?���3ýy���Q�2&�H?`�#�=��U?b�Q?2	p?�| ?��y�6P>�}����=�#�_��=��>�g2?��L?�*?oS�=0����d�MX���:��͟���v�>�hI>rY�>!:�>�>|S�9�I>ۊ?>�t�>�>�'=��ֺ:?=��N>�u�>���>q~�>�P�>�Z<����<a���u�TK��ĵ����?Of���>����֪��%e����=��>j�=�D��ŰοO����HL?4Ⱦ�v#�P#Q����=��?�|?��z��%߽��{�~�>jG�c�����=��%��x�����i�>���>��>�&=h�.���(�5�.�Z"����=?�.?�����B���L?��y)�Gھ�0�=���=.q¼'��s��q��54����>�<N?u	�>��ݼ����Z����ΤJ>7Ҳ>��뽣'�>sYk>A[�˪<�^��]^>Q�ѼV�q>�E?��=��i=W�Q>�������>�>�A>��>��o?<��>�����c?�_��YP�Ӊ?��>""�>s�=�������=^��>s�r=�K�8{j������L�9=�>:��<��]�"(ƽ�g	��ѕ>�:�<��b<n�d�mdt��~?~��䈿��aO���oD?�*?��=��F<�"�����D����?S�@�l�?^�	��V���?�@�?��}��=s|�>v٫>rξ�L�g�?�
ƽ�Ȣ���	��'#�BS�?�
�?��/��ʋ��l��6>�\%?��Ӿ|��>�������d��k�u���$=���>�H?����01N���=���	?#r?�D�R���g�ȿ��v��7�>d��?��?��m�� ���c@�k*�>u��?:$Y?��i>A+۾��Z�s{�>'�@?lDQ?0a�>|B�D&��?$�?㍅?��H>#��?��s?���>�w��P/�7/��0���{�=�zX;+p�>��>����pLF�B���;f����j�۶���a>�$=GB�>ǂ�RK��(�=}���mB��.'g���>,q>E�I>�3�>�� ?��>��>|K={V߀�T�����K?}��?����1n�C�<���=�^��&?�G4?p[���ϾLӨ>ȹ\?���?#[?<c�>����=���翿�}����<��K>*3�>�G�>�(��.EK>%�Ծ�4D��r�>�Η>�ޣ�Aھ`,��t����A�>f!?��>Ѯ=�� ?c�#?�j>�(�>IaE��9��v�E�ʳ�>+��>�I?]�~?��?�ҹ��Y3�U���桿r�[��:N>��x?�U?pʕ>>���ო��fE��8I�H�؛�?�sg?XW当?2�?މ??�A?6%f>��0ؾ{�����>NP"?u7V�-�6�k�����>��>�a�>�˽���s7���['��ݳ��?p�??w ?�1�h!`�l�ݾ}�<$��<Y8��Ϝ;�Q�<歬=%�>��k����=��>"=7���R�W%=�8y=y׉>Ew>�1��rx�s�'?�dD����� �=y�q��D�~�v>�S>{Ǿu^]?�4�\�w��A���b����_��m�?sJ�?���?p�˽��i��c=?@�?>�?�D�>�q��n8�Νݾ�5|���s�@a���>���>�ٿ���ھ5���B�����������9�Q��>y��>�x?l��>�N>
H�>�쉾� ����6���F�_�XO?��'���������E��?��ԻǾ�^����>6�[��Ž>g�?�b>e5v>��>1�6<fi>x�V>�}�>�>R>l�>-�=�O�D@����X?��(���$Ҿ:،� �?�kW?Ƿw>�O:1������&D?��m?��?��A>v�k�������>��!?��w��
�>�g>;/>Ŷͽ�����6s� l���竽��>���,�5�O�M���1�2�?�/?�i/<�L��M*�����סn=�N�?��(?��)���Q��o���W�z
S�z����h�U<��c�$�@�p�菿W�����ǡ(��A*=5r*?��?׈�އꬾ�k�L?�b�f>_�>�C�>Ż�>y&I>��	�]�1�v�]�P'�i���F�>�d{?7/>/EE?<{K?`�m?E�J?묇>Tb�>�J���?��>=r-?g�>�,�>�(-?��F?�?�l,?�̂>�>v�kҾ�`?��?��>�� ?��>�(m�����a��	�=>ۗ�~j,>�,�=�~�=S����O������=3O$?��e��+(����PX><J=?'�?>M>�Bx�_��'>���>�N+?��l>�����H�:O��"�>�`t?e�Y����;���>�+b> m½iμ��">ݴ���F=(=��;}�
���=�A�X"�;��j=fF�<!�5�^H>�U�>��?��>}�>U"��� �ё��7�=|lY>��R>�Z>�8پ���V%����g���y>�{�?w�?h+g=��=�@�=X��y\�����t���G��<��?�A#?�dT?I��?/�=?�:#?��>�>�~R��\P��1آ��?�+?�7i>=�ƾ�&����8:���>�J�>i�V����I���B���?��,�<.)�țM�|;��OP:�3=��<+�P�ѽ�[�?� �?�@�{�:�����)Y����??AyY>�Q ?��>��;�_H����S>\�>`]?]B�>6�_?�+v?��Z?Uu�>/� �yR��$���	T�=Z>>�h.?��?�"�?)��?n?�_#=������>�̾𢤼�Q��*]��D1ǽ��0>'6�>�ͫ>��>+5�=��޼^�Y��Z��W��=�m�>(��>&r�>8?4�>`��=A9?�V�>Rޥ��\����9����9���s?>Ps?^aJ?���/p�����⺾ֆ>�ʐ?"��?��?�l��ȯ>1��9Q۾jľ�>�l�>�3�>���*��<��-��Ԑ>�w�>���o��Fq��.�=� �>E+D?�h�=�_��äl�cľo�˾��7<�B���o~�RWڼ�����	=��V��T��*׾q�'�{x˾���e`۾{{��F��P�>`�=j�>��=��<�C����=���=C�9�=�<"Q�8�U=��@�q5+�c����(;_�<��=����˾�}?	AI?Y�+?�BC?�z>\�>�>1���>\`���M?McW>B�P��k����:��V�������`پِ־��c��ɟ���>��F��n> f4>
��=F�<���=yTm=A1�={/���=���=Վ�=�ƫ=܈�=
>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>ە>Bȉ��恿2�G�6���������_�W�?+Sb����g�>��������8�����:���bE	�/Q~��4��V���V�=e��=���>�A";� p=����k�>��=��=ML>���;DH/����=�z=|D>c�>0��=�p�>�Z?�>?�>?e^�>-i�����u�M}�>F�W=���>��o>ǂ�=y�	?�6�?��?��o?��>;?�>8֕>q�>�����z��f���Ҿ�f��˚?�>^?~�>�G�= v��*M��V�Y��c�-?a�7?��?��>U�+��V&�D�.�����ݷ>S+=Ugr�$6U�
2��v�"�㽦#�=�r�>���>�>�^y>��9>>�N>��>n�>�3�<Mj�=����ݪ�<�͔�r��=�
�����<#�ż󋉺��"���+�������;�`�;�Z]<�4�;i.S=��>� 4>ڒ�>���;b���e!>��G���9�~�!=��O�o�(�Y#U����,����(��`>{�>��]��E���J�>'O�>_A�>]m�?�k?�>	��g��ߚ��1�BEZ=K��=?�=�GQ��4�2�F�W6c�Q\���u�>��>>ƚ?�*�>7�
�o6��ٯ��Ծ;��o�>���Ą>H�K��z������YN~���o��H���?!�������B�y?��U?��?���>��f�o���o��>�@���'���c�#��-۽,�>��?Z�?<���Q˧���Ҿٞ�9)�>f�"�P4B�q��Q�/�!���:��n��>�ҾzZ���i1����)Վ���<�0�q�ӭ�>�M?��?����~���c�M�TM�����_C?Ӿf?c�>Z%?��?x� ���Q�D���=;}b?��?�4�?�L0>�޽�8��?? �!?�8�?��?�~?b��{a.?E'ؽy}�=:TȽ�ѩ��ĝ=�,�=��>�b4?8+#?�'@?�P��h�'�Ҿ�����#��
�=/��=aa>�8^=h'�>n>aE���l>x��><�>�#,>e>ۃ>�fz>i�̾'�+�ڭ6?��b>!,�>S1?n�Q>��=�*�=�n&>!¹������:��$½�FB�3^�L�=�Gv=���=ٽ>�Aſ��i?��=R���� ?�p���,�<>���>��>��>��>EL�>ʸ�>�%>�iq>.޲>�>���C�=rK���ۼ?�G�:�����&l>r���ʽ�y	�"U��R������u)��y��E��oM��ƽ�W�?�bX��s�(�B��=H� ?rB8>Л7?}���.���"1�>w
�>�S=��⾃Ў�$�P�,7澆��?i��?f;c>t�>�W?S�?��1�3��uZ���u�@'A�\e�f�`�፿Ɯ��[�
�e���_?��x?$yA?c�<D8z>Ϣ�?"�%�ӏ��(�>�/��&;�K<=+�>�*����`�׮ӾٻþB9��HF>{�o?�$�?UY?2RV�]wp���'>��:?��1?�Lt?[�1?�N;?N��[�$?�@3>|�?�\?%�4?�D/?�@?B1>���=ˤ���q-=�ґ�J��ۆн�I̽8���n�7=�ou=��ڞ�;pt=��<�4��~vȼ�z;�ᘼeҥ<��8=\{�=]z�=+h>�a?	d?=��>�1?q������N�ľ �F?����qا�'3���������	�>��w?j�?� q?�S�>6�hĠ�7�>ᦅ>�hn>
�>g�>|�=W?&��)�=�\>�b1>pEI��,ƽ>ʔ����Ǿ�%C<�O?=�*�>��y>4��uI#>c��Q{����M>/,.�	����R���;���/��Sq��v�>�XK?�?���=D�㾇��=�n��?|�<?ͥ\?�π?�G�=`S;��0��P���N�@��>�r�=����9��������8�r�b<^6->ծ���A>�q�6>�J�����&q���D��E�'�f>ݘ��`�=U��h��;�)�s�>`�>8�徸O*�����$՗��;A?տ�b���e�T�u�ؾL>���>Y��>�]��ȽI�9�'���:>�[�>�8=�� >�\���(��#�J�><�6?kF?���?����Q�:��D?�����#�-o۽4ZS?l��=�L?9�>�T<nͤ�����~Q���7�>��?� >��^`��o���񈾨���ʰ>G�>��m=��>�iT?�Z�>�?�Y?��>S�>׻Ž������(?3�t?,�<��|�爾�����<����>��?Э2�v�>��>�#?g?:�?
]�>' >������>/�i>�bH�bW���e>�Y)?�!�>J)6?E��?O,�>Nk�L�d�����ʻ>?^�<3�?C��>��9?C5�>�>Y>bU�����WB>�.R?�<?��?㗚>c�?����7�>�D�=t�6�Wv�>�G+?Txq?�o�?��]?�hD?DӚ<]wN�腽}�򽹛��*<�Q�=s_�>Q5�=�Z/��߽�=��=A��=ek���=�[�X{��G��#,�>IZ�>�W�Q@�>2����-{>O���aCq��������"I>9�>v`?6W>��:�E�>Q��>��>7�&��P?Z�$?4?�w��~IO�߭��J�w�~�>H0?3&�>��k�}ŋ�l q��v�:qXv?zMw?�a�9U����b?>�]?q���<�|ľ�c��o���O?5�
?��G��;�>�I~?��q?V��>
lf��n�����b�u�j����=ě>�h�� e��;�>� 7?	��>gc>�;�=�۾|�w�z2����?�?k��?��?��(>�m�=�Zm��{E��"^?ǁ�>*;���"?Oa��<�Ͼ�3��{	���%�8�������H��Sm����$��惾ֽ̅��=��?ss?�Rq?��_?W� ���c��:^��
��CoV��)�����E��E�	�C�ԭn��X����t+���dG=�a!�����?f�?�~A�q��>Fnx��ʤ���9�>�����^>s>�����N�>�T��`�����L❾7Q?結>B��>m�0?W�T����-�ԹC�r`߾1�>@*m>��>��?���.�N�<��=n����W����I�q>YoS?�P?�Dp?�L0�d����۟!����l��3G�>�@\=���>u5��䧽;����@��5f���7����� �P'�;��8?J��>7�e>o��?���>`�Ӿ�㵾<���X�T�ļ�?��\?{��>k(H>����$����>��l?Jr�>9֠>w���!���{�y�˽��>�ح>Y%�>�p>C�,�k�[�!\���u����8�W��=��h?�t��Αa���>YAR?�[:�F<�}�>��s��!��4���'���>�S?bv�=��;>�ž�={�ꉾ�R+?�"n?x'��pV�Z�?�"h?�q�>T���Nj?�j�>���u%>Τ	?��m?
��>*F?�=�>�>��B=p��A��؁]��Ô>N�I>f�=�k>�����9��Z��K���3�g>9���9��<�u</�NRҼ�g�=	I�=s�㿸\����P(�����5�����2}��Q����ß��H��������O�7��WƽG����q����^�4��?�� @>���]^T��X��JÊ���:�8?�:��Z�ۼ��mL=��'�C:�����m�5�a�]�l�Y����K�'?�����ǿﰡ��:ܾ ! ?�A ?5�y?��2�"���8�� >�A�<�,����뾠����ο3�����^?���>���/��m��> ��>�X>�Hq>����螾20�<��?3�-?Ҡ�>��r�&�ɿ[����ä<���?&�@��>?Q<Ҿj.ɾ�ғ<U?-!?>1E>6؝�{I��z{�A��>�9�?��?Pϡ=�-O�6����W?�"=<4��
��{��=l��=rh�=LT�	`a>�æ>RK��!����Ͱ�>��S>�ڽ����*r��eD=�j>a�W�M51�Մ?Oz\��f�z�/��T��Q>��T?�*�>.<�=F�,?�6H�Q}Ͽ֯\�2+a?Z0�?C��?)�(?@ڿ��ך>q�ܾ�M?�D6?���>d&�^�t�J�=!N��ޤ���H'V���=W��>2�>l},���x�O�c�����=]	�CпM��q3/�p��^�佛��`�E��5�����T�~�t��Q��l>�>>�B>8x>n>�^>'�X?G�e?%=�>��>��s�����<��<+x=^	��mj�9����<��JT��׾����B�"������'�H����<�uZ�b��8�=�Ȅ��u�C�ru??\\=M�����I��Ͻ��m�ٞ��A��hL�ړ��>��s�ѩ?�,K?�����N����{��bd=�ir?"ǰ�k���?���!>��k=�9~=���>��g>F����D.��]���O:?'T?��������=p-߽�>t�?У?0�=��f>���>�rD��>"p�=:��=�A�>Ǝ�>&�v=�F��J���5?�M?"!�-�����>+�Ӿ��E�g׻=$@�=� �n2��\a�=��>�α��^�=����6]�='W?���>G�)�� �,N��Y��==W�x?o�?I�>�8k?��B?I�<z�����S����9w=�W?��h?Ч>�����Ͼ�6����5?�xe?��N>1Yh����4�.��o�>R?�n?�#?���b}����n��s66?��v?�r^�s�����?�V�A=�>�\�>���>�9�Ck�>~�>?�
#��G��ﺿ�QY4�!Þ?��@~��?� <<� ����=�;?�[�>)�O��>ƾx�����:�q=�!�>ˌ��>ev�����P,��8?���?L��>���������=nc9���?"�?�Y#�L�=���0m��+��[Z^=Uw=�
"=�y�<����3�O��~޾u�(��,�<k-�>7�@�kҾ�͓>p��=Z�޿��ݿ�^��-�N�޾�<?���>�#�=V:ɽd�\��+(�I����~���Ⱦ9��>�X>Ч��/
��� }��/�������>:AA�â�>�"K�'i���K��Ϸ=p(�>!:�>d'�>��b���x��?�B����ſ�����T���I?�?۰{?�:%?���=����1|�����V?C�V?
�V?S��c�{4/��j?�]��=T`�C�4��FE��U>#3?�@�>_�-��|=d>ߋ�>Ic>S"/��Ŀٶ�{������?���?�p����>���?�t+?j�v7��jY��l�*���)��;A?�2>+���	�!�0=��Ғ�j�
?�0??{�4-�#�_?*�a���p���-��Vƽ���>�0���[��.��� �SLe�����.y���?�T�?��?�^��"��@%?%ޯ>a}���Ǿ���< \�>��>̨M>f(_��v>����:��	>c��?�f�?�t?�~��+��&>�}?6�>O�?
��=�P�>���=����:$3���#>���=�Z@��?|�M?�F�>R��=�e8�  /��PF��1R���]�C�K��>-�a?��L?^�a>���1�F� �{Rͽ�[1�_?�MD@�N�+��'ཅ55>�=>�>�E���Ҿ��?Lp�9�ؿ j��p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>;�>�I�>>�Խ����\�����7>1�B?Z��D��t�o�y�>���?
�@�ծ?ii��	?���P��Ua~����7�h��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>!�l?��o�P�B���1=7M�>͜k?�s?�Qo���g�B>��?"������L��f?�
@u@a�^?*���A�����̾>
�A��=r[��˿=����<�$����e��b������c�>�f5=
�ɼ-e>e>�.N>�b��j�$�Β�����8���c�˜K���&��оu���6�0���&���[�D��GOs�L΄��?l�*��<�:�=��Q?ZR?|�r?m	�>(X�bG>�����+=a��ݐ�=o6k>�A3?�P?+k*?��w=�⣾h�c��-~�5�������Ĳ�>�$O>�v�>���>Lٮ><�Y;�AP>��->��>zF�=ꔶ<��O<BQ�<�@S>䣪>r�>F��>&>%��=������;Mx�<���^E���?���{� �4Ɂ��%ž���=V
?��.>$����S̿������P?=���P���<��A�>/�G?|yN?��>n��xT���k>���<[��d�=S�l�� �=��U.�>ܿf>Q�>d>"lR�k�5�k^=�������rL?�l.��a�<��A���A���¾����P��>�W��A3�K ������[�3�=��=?��?�.���v��'��u!��+f>��>�=M������>��"=�{�:���J��)�����>��?�68>�Q=XF�=����P���Jѻ>��J>�D>�p]?@�?�����$.�
鷼
�l��ns>P�>Fޝ><'�<��W�7R�=˺�>�q�>3�I�֎)���'�;�Q�Y�8>�6����J��ؼ`u�={�ݽ�D�>�ʽo[��ȷV��y!<F�~?�I���Ո�� 뾦u���D?~?zz�=�X<�g"��q��m��?��@%�?�|	���V���?�	�?�O��L~�=�>GU�>��;z�K���?f�ƽ�ˡ�8	��.#�v&�?7�?ۿ+�Z����k��o>��%?�HԾpl�>st��Y�������u��#=T��>�8H?OP����O�3>�6t
?�?�S�<���L�ȿ�{v���>�?���?��m��@���@�]��>��?�hY?Eni>$^۾n`Z�>ƹ@?�R? �>�9�E�'���?�?���?�I>o��?yIs?D��>b^��.��������?I�=z�!;�>�>G��	�E�/{���	��(�i�:)��|a><S'=b��>b8콆������=5q}������j�R �>=�o>�F>�r�>��?G �>kM�>�
=:����F�y��L?h��?���; n�y�<�[�=&�^��*?CK4?Bs]���Ͼ���>O�\?3Ȁ?�Z?�=�>8���)���ۿ�.i��'ܕ<�K>��>�0�>�Ɉ��K>�վU�C��j�>��>&����.ھ;������0�>�Q!?��>~�=�� ?�#?�Oh>蚲>�E��s��d�E���>�8�>�:?=�~?b�?�����1�K���\��=&[�z�H>w�w?.�?��>�p�����W�lT��(��Ԃ?��f?�gݽF?nň?�>?�~A?�c>qT�H�׾������~>��?$�Z���?�����2����>8|�>p?�[���=�藡����{�پ?��.?8�I?������F��O���2�<�~*=��y<T�ɼ�U��#�=��S=�=���?>�z�=Pm>,�<����>4���7$>&�|>2o�;,aӽ�x9���+?���*���W��=��q�E^E�BN�>zJ>iC���_?�@��z�z���J����J��Ë?J�?��?�����1g��:?7��?D`?+��>�*���⾎羅ڀ�?G����5U$>�1�>��]�پ)���*���'���"ӽ&�_�[��>�J?��?�D?M�>c^�>3}���F׾�������SC��	/��7J�9�C�(�����=U׽��:=$��$�d����>����	?�w�>yM~>�n�>�?�>ρ:q�\>I^�>�>@ɪ>�z8>�/b=��<�;�=Kև��fW?3���'��T�$����{7?Ne]?���>�@�;{߀��Y�Ǡ?"ԏ?=�?�iO>��b�]�.���	?��>�Fz��� ?if�=w5=�h��;����>�ƽ��ܽ��4<��>��ҽ�'��5I�:V�J�?�{?@���^9��@��+���Oo=�M�?��(?.�)��Q�r�o���W�S��}�f8h��c����$��p��ꏿ�]���$��?�(�-o*=�*?9�?���L��q!���"k�@?��cf>��>K$�>	ݾ>(xI>I�	���1�j^��I'�+����P�>�Y{?��L>l.e?��U?t�4?q?���>v�i>?g#�n�>�WN��	�=��-?r�9?]?�	_?-�?W1U?2&=;]/>S���3'�C�B?��^?K8>�y>�M?R��Ͼ�h$>A�>��z��󓾸�ܼ�zR>I��������"����S>ѫ$?9���8�ʗ���	!>26(?�H�>?��>��A�R낾��˻�y�>V�?��>���h��g��Z�>K`k?S���.z<�p/>50�=���hZ/=R`*>΅���H>��.�<U���=���=}��=�ǟ<�*>�(��>��=�#4�QU�>��?Ŀ�>���>�텾� ��m�mf�=*�Y>zS>��>d�ؾ����(��l�g�|!z>���?�~�?�2j=-��=���=X��iI��b��>�h�<n�?�6#?�,T?���?3�=?Q@#?]}>+�,O���I��J�����?�0?X��>#Ҿ�������Y�(���?]�>�;�d�ļ �=�Z�H�����X>�`��d������>Y��rJ�8(ƽ�?G�?+J ���#�����`f��&�ľˢM?��l>|u�>��>�SH��C�f]��4>>$�>'U?�J�>�b0?��{?�NB?��=�ǾY����_��Q��=i�>��?d�G?��?��*?�>�>���=a͖������V���u����N�'���)A>�8>_�>x�|>o�>i�]>��a���r>�d羫T�=E��>. �>��><��>Y�=��P>!�H?���>�ľ�'�b)��%�^���N��j?�?��8?�S<�� ��B��ܢ�c�_>쨢?�'�?��?��l�˖�=Aк��~��3���,�>�5r>�'�>@֐���3>�H|>�y�>��r>-Np�{B޾=�:�Ai��k'?�m?fҘ=�i�H����$���x�<x���˾V��  �T�L��������o��~fO����,ݾ<��h��� ����>��)>#�>c�=%�h�H�#�M���i�?����<�o>ʬ��˼佊9�<�&=,>��=�x��ٞ�6t�v˾ȇ}?t*I?��+?��C?5�y>�>��2�$w�>z��VS?��U>�&O�^���n;�ڡ������ؾp�׾9�c����R>�$I���>E3>��=6��<i��=5#s=L̎=J�I��$=8�=��=�y�=�?�=S�>�l>W6w?c��������4Q��X�G�:?�9�>P}�=,�ƾ�@?��>>�2������b��-?y��?�T�?A�?�ri��d�>����⎽�p�=?���=2>_��=��2����>��J>f���J�����O4�?��@��??�ዿ��Ͽ�a/>`ȟ>9=M�q�����=��/d��D����V?r݄���⾲��>��m��t^����|�<G�>�6��1��q�����=���<���=�>�=�\>0?>��=
��f�&>?E=�G�=T�->��<�C佉9�<�何	�>�x�=��D>K��>Z�+?(D5?�j]?Xc�>H>�<7���6���q>��v>eȜ>��&>��>R�|>��)?P&?k�@?MF>\g>�z�>2�?�c�ލ��ƅ��B�^�����v.H?�Ҋ?+��>��/����,r��d ����uN�>�)?�#?S�p>��;�⿸o$��N3�sŽ}��J�ټ�@��]����ƽ�R.��,����>0'�>q�>�:�>�~Q>��1>��b>��>���=	��=�G�=�0���ێ=R!d< �={�L�c�=��<Ϗm���%��=:�UZ�<�V�md�G�ƹfz�2+�=�4�>�-t>��>�t�=�㤾�F>�q��s@2�B�.>���tY5���c�. z��)�B|U��P6>uNJ>�k\��X��C��>w��>7sy>��?�=}?�I$>��$�ϗ��zp����s��>����=<�1��@'��Z+��b���?�������>�>`6�>*��>��(��c/�(��=����
�/d?�.����=j�Z���Z�p���㜿h|R�^ņ<�-1?�����D�=A�?e1Y?긶?)'
?cI���Z�5�s=�i:�8��=v'�㊻�o��Ó�>�{)?&/�>������%T̾�1���
�>8 I���O�����$�0�L��������>����оP'3�e������z�B�5ar��>T�O?��?�ib��Q��KPO����؅��b?�vg?\��>I?4?����^�s���=��n?���?X>�?��
> 6�?k+�"?T�d?\��?��y?��?(e;���/?x���
�>�	>[C��I}�ŭs�� �>��p?�n?�h^?������}����Z�[�4�뽹,����>�u�)�>YD<��/(>G��=��>�r�=k��Q�>ζ>>A��(���+F?�j>>��>Cs5?��>����=�j>40��C2� 6l��\�}���/*��с�*@>��=s9�>����ć?;�L><��[Q?"#���!��&�=L�<>��
���>��m>m�5>�_�>���>�#'>ic�>Z�>!Ӿݒ>����W!�+1C��xR�+�Ѿ�z>�����&�ܔ����SI�R���_��j�`+��==��ܽ<�E�?P���$�k�k�)�������?[�>�6?P����È�#>���>�>���+���5�-lᾫ�?G��?�;c>��>��W?��?|�1�u3��tZ�;�u��&A��e���`��ߍ�W���p�
�H����_?��x?�wA?�p�<;z>ƣ�?I�%�܏�o0�>�/�L';�`*<=~-�>(����`���Ӿ~�þ~/��GF>��o?$�?�X?�PV���i�.o)>�F:?{�0?�pt?"O2?��;?�C���$?ލ4>bI?�8?�5??/?��
?�2>�w�=ME��to,=��wŊ���ѽ�	˽���A�4=N-x=S�v���<��=T��<Q �!j輈�b;����Ռ�<BI9=�Ѣ=�=#ޕ>��M?�?��>�6B?1���<O ��Ԩ�Ӣ7?5�r=�K�������d;
���=b�u?j�?��b?r��>�6�>e�R�#>Qy>�V?>��O>���>�|�=�U4�^=�4>��=�j�<�w���;S�i��!r�)`�=ׄ�=�A�>	�>!���
>�#��1镾��d>�T�)��Io����F��"�I�j���>c�K?��?,v�=�ؾ9�ཱུ�`�Vm?fHM?Z�J?��s?�v�=���P�L��S�@�E�kR>�+G>d羲լ��`����8��$��
�->�1��%��1u�=�� ��+=��pl���&�{��Z-�>�z�Uր=���澃������3�>�0ھʨ�����
)��͂K?��N�9�V�ZzY������>d��>�uE>ot�� ����^�=��<��?,ub>�{=�?9�_�.�;�t>9Q?��Z? �w?�+��p"I�ʉL��g�����:\<*n?A��>"#?*��=��=���)
��<u?���I��>�*/?<|,��-e��������;���>eO?���l�>��x?R7?��3?}�+?�?���>֤"��վ� ?���? ��=rĊ����:&���@�߅�>��,?_Ζ�T��>��A?h�P??��K?��?�:�=�˟��Q�yR�>��>ŤM�*����*�=��?�M�>��'?���?F��=��S��l��z`�<t>�7���+?z6??��?O��=N�>%Y��Dc�=��>`�b?;a�?�:p?4��=s?�2>��>�.�=R)�>�W�>�?�O?	�s?HbK?h!�>�k�<ȼ��W+���Rs�PPK�c��;�
S<u~=�C�g�r�����<�Ր;�㽼X�������F�����.��;�H�>͇�>F(�M��>����z$����>��½����	���f��h>�>��>a��>S>-�&��FR>�Ώ>�!�>|0/��~?h=?�/?l_��l�:�F�3��A�>W�"?`�>^���ץ���p��:�p=8��?�R? ���栾1�b?�^?���=�Aiþȍb����*�O?z�
??:H�{�>�?r?�u�>�e��n�����b��Aj��-�=���>�R�>@e�?�>�67?	�>��b>)�=��۾��w�埾1?��?aޯ?��?�T*>�fn��1�)^���)���.^?�2�>����-�"?���[Uо�뉾�m���h�DW����������5�%�����C�׽A��=�S?ڵr?� q?Iv_?V �f�c�j^�}��9)V�%���;�mjE��D�=�C�6fn����um��f���bS=�G����.�x��?+ 2?�Y7>��>Ḩ��f�֛�!��>�5׽������P��I�>�K�>}��T/�A��0�ýBf?�ڬ>���>��/?7'G�u�C%� ���!���P����>�V�>2~?��J���3��|ƽ3�����뎾 +v>@rc?P�K?=�n?�R��%1�Q���~�!��/��W����B>b>��>��W��o��5&��N>��r����Lp����	�+9=
�2?	�>���>dH�?�?�~	��r��
^x�'{1�Uσ<["�>�i?)�>GȆ>�Sн�� �ߣ�>ܡl?�W�> 	�>̦���c!���{��Ƚ��>���>R��>h/o>@�,��\��R���k��h�8�hH�=�zh?gh��|�`���>�Q?Bq;9�lU<� �>��s�ۭ!������(�`g>T?{�=��<>��ž�N�ً{��*��&�/?�&?�$�w%�z�>�k?���>{R>�U�?ٗ�>#Q�	~>�"?a??��+?s1?wK�>�� =w��㸝���S��d�=E�>2�>���=��>�e��pzͽĔ�}'	�^�)>U���g�	V��|�W��
	=%���>���P/|�� ��>�,��i3�n`�an��Gý;��%���-
����5׾o���/��l=��w���Ҿ�rX���@R�?��m>�1�����:���>��Ծ����M������,s���������hf����g�Ís�.�'?Ϻ���ǿⰡ�;ܾ,! ?�A ?"�y?��D�"���8��� >#:�<*��	�뾉�����οp�����^?���>���/�����>P��>�X>�Hq>����螾54�<��?��-?���>��r�-�ɿ����¤<���?�@��@?���y߾l�<��>�?��;>��:�ֿ����̋�>�A�?�<�?��X=�[S��3�H�c?�c`<M_?�8Ԅ�	��=��=��=�O�ta>e��>��6�LK�e��"y>r��>�����qv��bb<��r>0��m�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=u6�퉤�{���&V�}��=[��>c�>,������O��I��U��=�d��ƿ�$�f� ���<j�Ȼ �Z���潜3��VRa��㡾aHr��	�j2j=Q��=�V>+׆>Q�T>V Y>}�X?�{k?��>,>O<轳���KϾ�~+��������9��k��ܚ���3��߾��	����;��H�ʾ��<�b�<hv_�dJ����9�q�R��
C�k�'?.֕=����p�3�e�1��ľb���#琽B"�l����E�e�o��y�?��I?cG��dN�ò��|=��>��_?���Ξ��m�]|!>�h��'v�=>��>���=�\Ҿ�� ��2e���)?��?��۾0���,>4ք�KY�=�?�b�>�=Cdn>�>:�sSz�3��=D�>K�>�ƾ>���=�����uؽҔ?�vE?*J�d#��N
�>�P���yJ���">���=L E�KC=��'>��N������l=h�С�=

W?�؍>��)�����3��X����;=��x?F�?�ß>�Ak?��B?1}�<=S����S�K�
�)�x=K�W?��h?׿>9���C�Ͼ���k5?o�e?.�N>��g������.�j��;,?Gyn?�[?~���p}�Z
��_��zI6?��v?s^�xs�����L�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?��;<  �R��=�;?l\�> �O��>ƾ�z������/�q=�"�>���ev����R,�f�8?ݠ�?���>�������j�=�iq�?��b?&�|IX�e���~�=�Ӿ��e>N&>�$O;_�C� �þ �#�G����
���� ��=�>K�@Tl��n��>w����UͿ�&Ͽ�#�����	�����>4�>�8�>�Ӿ\�1Q�6���9I�n����>'>3�����S|�09�!gļ�J�>Zj����>��]�NK���J��<��;k��>3��>Q��>�ɽ�뼾���?�}��d˿�4���y�R�W?b�?ǃ?�)?�@:<@�g��瀼 ?H?ffq?��X?�L?�D�R�pTn� �j?z_��bU`�ю4�cHE��U>�"3?�B�>J�-� �|=w>���>=g>�#/�u�Ŀ�ٶ����N��?���?�o����>{��?�s+?�i�8��X[����*���+��<A?�2>(���O�!�K0=�UҒ�Ǽ
?S~0?{�K.�\�_?*�a�L�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?M^�?h�?յ�� #�f6%?�>e����8Ǿ��<���>�(�>*N>hH_���u>����:�i	>���?�~�?Rj?���� ����U>�}?�)�>#�?��=�`�>\��=Z簾+�.�l/#>JO�=B>���?�M?m<�>�&�=�8�/�aUF��BR���I�C��>�a?|}L?��b>�B��Μ2��!�A�ͽ1�漻Y@��L-��߽5>�=>u%>k�D���Ҿ��?Mp�9�ؿ j��"p'��54?/��>�?����t�����;_?Oz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?X��D��u�o�x�>���?
�@�ծ?ji��	?���P��Va~����7�l��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>!�l?��o�P�B��1=8M�>Μk?�s?�Po���g�B>��?"������L��f?�
@u@`�^?*�1���ÿ^־���^��<tT�L~3>>�m�
��=j�=������<��R<��>e.�>W��>;;�>M�A>+�V>�{��*������څ�Ŧ3�˽���o����Ӿ�&��n��	��l%��ˉ��R�ѽ��� ��U�������=��T?�dR?�{p?�� ?ˤp�=�>Z��� g�<): �P4�=�M�>��1?M?�+?��=������d�!ր�奾�T��k�>�}H>���>ei�>��>=;��I>�C>>ڭ�>Љ�=�.=�lػ��<2LL>��>�
�>it�>�.>~ދ=h ���X���+v��K�Ԕ$�c��?"l���L�����꾾2Ѵ�?��=vm?Z��=0፿�ǿW����n\?�z����!�{���h>x�/?��]?P�=d�⾬��G��=�  >�k��]� >�a��8�A=��٠>u^�>��>L��=U�.�T�%��RE�ef���=[�3?�I���7J�I�>��u.��2�����=��L>*
x��9'�V'i��*u��D����>�04?q��>���<f�X̾1Rҽ��>�/�>>�{<2�3���>�����>���(��<��=��><� ?��.>@���)/�>�I��R����*X>�!x>�>g�$?ƨ ??7|��~>��@햾� ?a��>( �<�]U=��u�w����?�	�>$���7.>�L�)C7<;a\>qB=�a�YF��Ɛ�/9��.m�>g"�m'�cy��m�U>�~?���(䈿��e���lD?S+?^ �=#�F<��"�E ���H��G�?r�@m�?��	��V�?�?�@�?��J��=}�>׫>�ξ�L��?��Ž4Ǣ�Ȕ	�2)#�jS�?��?��/�Zʋ�<l�~6>�^%?��Ӿ�g�>&y��Z��g����u��#=���>�8H?�W��=�O��>�(v
?+?�]�ʩ��M�ȿ-|v�F��>��?���?&�m��A���@����>��?igY?�oi>�h۾|^Z�8��>��@?�R?��>=:�ҋ'���?�޶?p��?K�H>\��?e�s?~D�>;u��</�g,����1�=��{;F:�>�>�A���\F�ϻ���U����j����5�a>��#=��>��0:��SK�=�"���-��=$f�7�>Joo>�cI>���>�I?�,�>��>4E=�ڇ�kЀ�)��=�K?$��?J���*n�_��<Ir�=��^��?H4?�\���ϾNڨ>N�\?���?(�Z?�T�>����/���ܿ��u���<g�K>�*�>�G�>�?���K> վ�D��a�>)��>���~5ھH:���(���-�>'_!?lr�>Z�=�?�&?��u>���>߰;��䍿AG�H��>��>�?�?P}?����0�0�v���|8��Y�CK>v�x?��?W��>�������&���ַ�Xli��	�?��k?�Z�"6?#ۍ?��@?=~;?��l>��:�ܾ�i�]�t>�$?eZ�,�:�-���|���6�>���>���>~r���
�/��(��!���Av?�
+?&�!?Bi��fF�X�)p;�>�<O�G��tCH=�q�=n�^>�K�c�G>S>��=Eo���*�yݽ=�`=*a>*W�=�c��NR���9,?FdG�~ރ�)��=�r��xD��>�]L>L����^?�D=���{����Ww���U�
 �?���?Jb�?c��a�h��=?��?�	?\	�>c3��h�޾�w�-w��nx��v���>Y��>��k�\������i���E���Ž\��d��>�y�>�p?�{�>TA>�G�>#Ǚ����H�پ���(�J����0�6��%��u
�����%���<lվ��h���>V֣�䝺>�?�D}>=Ԙ>ۣ�>r�����>��>SQ>n�>��>|Y>o�=��I=�H���;R?���V�'�z��P�����A?$Wd?��>�h��n�����O;?5U�?�m�?6�u>�Yh�t%+�N?��>�:��X
?�;=j�É�<n���[@��t��#����>�X׽(:���L�T�f��k
?��?8���73̾�׽P����on=�O�?o�(?Y�)���Q�6�o���W��S�����&h��L����$�3�p��⏿a��"����(� +=�*?�?|��.�����.k��?��0f>���>M!�>o�>NxI>��	���1�Y^��N'�㪃�5O�>�[{?+��>kW?}�*?�5D?bM?^��>�/�>�о��?��T�=�S8?��D?��?�>r�>�d5?p�>ڗ�y���*�
�*�!?ǋQ?L�>�?�/?���-U��|Y�=��V�ao\��1�;<<:[�W��:�8���\�s�>$�?w:��&8��0���`>�+0?Df�>ʓ�>󒌾Y���+i<E$�>4�?�d�>5����l�%���^�>�|?��A=x�%>y��=���d�J��=����C�=�i���:�L�;;i�=&�s=p2h;X ���A;��;ZZ�<�s�>�?6��>B�>�?���� �����t�=�	Y>)S>d>pHپi|��?$��^�g�xby>�v�?�x�?H�f=��=f��=Bw���Q��|������>��<*�?{J#?�VT?���?.�=?g#?-�>�%��L���]�������?�W-?"�r>��߾�C��:B���%�lA�>.�>)�=�
.��A�����B����=���k�n�U���1D��P<>�ځ�����?$V�?�S�2�����ՙ�Py���G?�?��>���>�e(��/Y��c,���M>��>q(h?b0�>�j?=p?�@?ql�>�u�韢�������<��@>;C?�v?*�?ԝn?kB?�ч=GZ�9�	����ž|O9�gJ:�慾��0<@�p>��>
��>�i�>���=�C��ݢ	>�x�C1t=
b�>�?&kd>I5?��w>�==�G?3�>2h��k��ō��j���|;�pVu?3��?�Z+?��=-U�VzE��l�����>^_�?~ϫ?*?�S�;��=>2ؼ�w���p�	��>\�><<�>T!�=�G= >���>�n�>����1��]8��>J�V?��E?ܳ�=�Ŀ_�q��So��	��Ұ�<n|���c�>��\�
f�=6��cX����xZ����㤕��x���}��$�|����>�օ=��=���=�<~�ټN��<0�I=>y<�
=M�o��`<~�0��	�䋽�	廇O�<8Q=X^ĻP˾��}?(I?Q�+?�C?�:y>�>�&3����>Y���� ?�U>MP��ʼ���;��C���ߔ��ؾF׾��c����J3>�vI��p>�{3>�;�=g�< q�=�s=`��=��\��=��=b"�=�Y�=*��=m�>Nu>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>p��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>ࡵ>����q���/��e\������?� [�,A�k�>��1�C;�gþm�ξ���>��ϾX�i�嫄���K;Z}=���=�+��G�>���`=��X�o.�=�Q�=V�&>�x�=���=放_2�q�/>!�U>Q��=q��=�ʡ>?6G?�ڈ?��?�;o���F��Nr�=\I>�WI?oሼZ��>&�>�Y?7U�>4�)?v�(>��E>�4�>���>A�1���i�"���b��ӫ��?Z�w?�1�=�h��%�r�X�b��+ʾ�M�>�7?�?gb�>�U����9Y&���.�$����|4��+=�mr��QU�M���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=$�����<�vż�����u&�:�+�1�����;r��;B�]<^��;���=��>_�>���>��=}2����.>Z���[qL�7�=t���@�A��d�-~���.�,6�>�B>bmW>�w���&����?��Z>�?>�U�?�u?k>��O�Ծ%��ʸd��S� n�=OE	>Ir:��P;�LC`�(�M�		Ҿ��>��=F?��>���Zq�w���:�jj־��M?(���K>����\�Z���m��먿�O^�%�ֽ��J?�����Ƽy�v?�F?�+�?j��>�p�=���x�>�P���~>�k �����=��(?%�>��>�fo�m��E̾����з>�>I�L�O�㾕�"�0��2�bҷ�V��>��<�оg!3�d��(����B��Ur�Y�>��O?�?�b�Y��hSO�m����nn?�xg?��>C?�:?�ɡ�i�	t���_�=�n?|��?h9�?��
>-d�I�=�Y3?�r?��_?���?�=�?l���el?#O���y>�d�>�>=^-=n;��;=U�s?Yh�?:N�?��^�2�#�6IܾUC��"b�5&>m�?�;X�>��=;A>m��=�K:��ýy�>ƸA>J��>���>��>������(�=?d>���>?�?�xt>q�[���<�if>�p����ƽ����v�%�=tR���E��v=l�<�)�>8=��BA�?��=��žJ��>�o��6��=�X>�ۥ=QR��)�>)��=4ݲ>���>o�u>l��=Y�>s��=�FӾ�J>���~_!��$C��yR��Ѿqz>�����&�ɔ������uI�xX��a`�j�a.���8=��l�<�F�?������k�<�)������?�U�>!6?������׶>l��> ��>�>�����������K�e�?���?�j`>$5�>
�W?�?�p)�oE5�7�Z��v�+�?���a��_�4%��+���\
�y�½��\?��v?4�@?H1�<X>x><��?�}'�����a�>��+�Y�:���==u�>RϷ���d�IIξ
��A�V�J>hr?���?7l?Kc�R�m�� '>ű:?�1?+Ot?��1?�;?����$?�n3>�E?2q?�M5?r�.?n�
?.2>K
�=�����'=�6��W��ѽ�}ʽ����3=�h{=�xݸ5<n�=���<b���ټ�v;�(���4�<�:=X�=��=��V>P7k?��>���>��[?!��n�>�ƍ�]k?U��>54<xf��5޾}A><��>`?l��?��?���>%��}�ѾLj>HK ?ϳ?>t C>P�q>2��g�t��=�N�:q��=�e���˱=~�T���ɾg�ݾ��?�?4>���>#[>2��*6>þ��h�z�;>����&���N�M^X�Yk��\��k�>�F?��?{�<h�lo���h���?��B?��J?˷y?x#=�����GB� iF����9��>[=7;�� ����)E�	��<��R>��A�=ֽ�T>��ھ0�J�U��H+ ��'��� 5>�l��`�z=�/���lھGq)��Za>�W>�!�=���������3�T?G ���D˾�ѕ��$���>x=t¾>F,>�IŽ9μʬT��
������X>?N�-=�'�=]F�H�O�?���b>��N?p[?�Ow?���4�]�$eT�,o	�GS���k==��?;L�>��?��>��=�1ľg�޾x�]�~m$����>�*?��+��S�3�_��������O��=r?�rF>Ɓ�>
P?�?�H?+* ??�?���>� �ү�� $?��?'~�=�!޽�B�	/2�4HG�m��>J�'?f/��И>��?�b?�&?X�P?�9?�!>M�����;�ؾ�>K�>P$Y��ɯ�"�c>��H?��>��U?���?m<>��9��������^3�=�J>�y3?Vn#?V�?��>@�>������u<�ʬ>�N?J�x?s?��>Ee$?F�=��>kA =�G�>
��>� �>��U?��i?9�U?a^�>5�I<��������"v�\�ݼ�&<�pR=�9�=�y[�Q�r:F\ĽK�P<i��<�ꜽ[ļ�h�����L��2��8��>��y>p��a�@>�g���wy�dqZ> �:+��{���sE���=�|>��?��>�k-�!�=.��>Q�>A�J�#?*!?�]?!�8��)d�	�Ͼ��6�
ط>"*=?}j�=�dm�8哿�s�ƅ=�n?�:^?�cQ������b?*�]?�g�6=�5�þ�b������O?q�
?��G�a�>��~?�q?���>��e��9n����}Db�(�j��Զ=r�>eX���d��>�>]�7?�O�> �b>��=�t۾��w��o��?�?��?i��?,*>��n��3࿨���F��^?�}�>f1����"?O���f�Ͼ�R��|���%�@�������I��$q��(�$�F%׽��=@�?cs?�@q?��_?b� �� d��=^�� ��jV�K1���u�E��E��{C�ݲn��]�������"�G=b����%��5�?H�?s����I�>w����� �*꽾U�>�������<>�C���}�=k�<�
Q�.fO��.L�x�?=�>�>�>�T:?�%4�P���<���2��&"M<���>w�>�>2�=�½��#�����9F�zYڽ�=v>6`c?stK?��n?
��1�?����p!���/��U���C>��
>���>~�W�Go�9.&��K>��r����Y����	�	�}=��2?v�>�ݜ>XF�?�	?�s	��T���x��s1���<�&�>(i?K�>~�>iн�� �;��>��l?��>*�>B����H!���{��_ʽ��>�ҭ>���>��o>Л,�\��b���|���9�+�=̠h?T����`��؅>R?y�o:�K<�b�>!?v���!������'���>:�?Ԫ=��;>ޘž4�r�{�M��>�?
�(?��a�f[/�{��>NS#?��>�|K>In�?&��>ͧ��q��<�l?�O?�\,?)?D?��>���=`"��� ����8�咻�Ir>xc>"P�=QV]>:-�nO�g����;��=G���Juٽ��-:�<7.����<��>�P���v�ê��R��(��a�*پt�Nr��UE��e���C;m�O�X,�������>��E�5���b��^�	@�D�?�K��v���:T����3������>?������ѽ۩1��і��m�
���'��ZA���`��z��%��˔'?3�����ǿ߰��;ܾ#  ?�@ ?1�y?U�G�"�P�8�Ҫ >�(�<g>����뾲�����ο������^?���>��0�����>b��>f�X>�Fq>���I螾�;�<L�?v�-?��>��r�Εɿ����fƤ<7��?��@�??���JC�0�v=%� ?i�?9(R>|�R����ȑ�����>Wl�?���?$~�=ގQ������Z?hbn<�F;�{��M��=���=��=[۽��D>��>��;�1}O���1�l>�J�>�4�S����gh�^y��6>�R�@er�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?$�(?;ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�܅�=t6�؉��y���&V�|��=[��>c�>Â,�ߋ���O��I��W��=�O�F�;3��l3�av��ۉ��|3��e�a����6��ܾy꥾�׽��>�\>�&�>4��>�>�y�>��`?<�T?���>�?0>��u�%gE�&^���0������y �mǽ6�3��� �2M����[�(��(�����	����4<�@G=�;T�5N��H�0���j�!�P��0A?�k�=��ݾ��@�L-��MӾ_e��s�~<^:?�Ra�2[@���v��Ũ?*�C?'����W�������z���hf?�����x����3>�g����<���>��=�u�7�X||��8$?�8�>r�����"/�=@	m�]C>�?��>8���?P��>1,���0*�ΐ�����>�8>ng#?7�|=�����p��v�>ߣ?8�j�(����N>6��v���x���"�=E���Z���-�=W�<7Ԁ���'��=%���*QN?�6�>P����E���R�2>��=S@?�?�	�>l�=?�O?�Cc=�~��Ѱ<������=ƌU?PP]?>�ӑ�ET׾n�体�@?.�n?靝>2q�����vse�c'�+�5?�P?�0&?r���g���ۡ����ҕ+?��v?�r^�gs�����5�V��<�>�[�>���>r�9�6j�>�>?�#��G��غ��gY4�Þ?8�@W��?½;<_!�X��=j;?\�>��O��?ƾ/z��������q=� �>����ev�j��SS,��8?��?>��>蔂�����=����$�?�{?e)� �����~?X�j�����'>�㨼������=	c˾�3%���쾼���S��ã�=Gț>H�@������>��=��ο)�Կ���t���wԾ�~D?�u�>�����4>D�C�W���Ӿ��+����ų�>	>wϓ�.���(�}��a7���d����>C��8�>fU������h����<0 �>C7�>O3�>�+ֽ����<*�?`��p,̿������o�S?6˞?>X�?CW?M{Q<W��r�q���Ƽ�L?�&k?��[?� n�2e���d�#�j?�_��uU`��4�rHE��U>�"3?�B�>O�-�Q�|=�>{��>g>�#/�v�Ŀ�ٶ�8���X��?���?�o���>p��?ss+?�i�8���[����*���+��<A?�2>���C�!�A0=�RҒ���
?T~0?{�_.�]�_?*�a�M�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?M^�?h�?յ�� #�g6%?�>e����8Ǿ��<���>�(�>*N>pH_���u>����:�i	>���?�~�?Pj?���� ����U>	�}?�$�>��?Ck�=$a�>��=^ⰾ{�,��U#>��=<?��?��M?�F�><t�=��8�j/�tWF��ER�U��C���>��a?J�L?`@b>�
���2�!�!IͽlQ1�)Y鼴_@�Nt,�vy߽%(5>��=>�">��D�S�Ҿ��?Np�0�ؿ�i��/p'��54?���>&�?.��մt�;���;_?�y�>�6��+���%���B�P��?�G�?2�?v�׾HT̼�>��>�I�>t�ԽO���)���C�7>)�B?*��D��;�o���>���?��@�ծ?ai��	?���P��1`~�߂���6�>��=��7?�2�Z�z>���>��=Kov�����q�s���>�A�?yz�?	��>T�l?M�o���B��1=�O�>֛k?Gu?!fq����B>x�?-�����EJ�&f?+�
@�t@�^?���hֿ����_N��N�����=���=׆2>��ٽ-_�=��7=��8�@=�����=q�>��d>#q><(O>�a;>��)>���P�!�r��[���T�C�������Z�C��Xv�Wz��3�������?���3ýy���Q�2&�>?`�	��=��U?�Q?�wo?=� ?�fh��Y>ub���.	=��!��=,��>9�2?�FL?LW*?=C��y�d�(���4?��ĭ��l�>��F>� �>��>���>
�ź%�I>�0?>
�>��>��)=���R=��Q>���>{!�>�#�>��>�=���6]��vSl�����e^�DH�?H��Y�/�����
����<F?\������Hǿ�M��6hT?�꘾E�#��
|��i�>�#?�R?���=���>�!�!>8B�<^V��6Ex=�+H�j�Խ�����>7��>�0t>���<ѯ/�WW3�ܯI�l�վZ{)>�1?�����X��M�jz[�4���bX�=:c�>��U���I���r�^G���>���ͨ���"?�&?�n���U�܊��7�ڽVs>vx�>ۮ =;;� X>b���aGm�j.��;��=�Ƚ�|%?��>�X
>o)C�YŘ>����rj�����>��>�[�>G��>�<?�Ծ{�D�%�T������u�>^|>�̝>J��>�K�����=uj�>ޅ�>�]L����= ���	�$�d�I>��=&7�������>㭽^�u>�-��3�<=���t�>K�~?n}���∿y��C��spD?�+?��=��F<��"� ��1=����?�@�k�?^�	���V�F�?_@�?���R��=z�>�ܫ>}ξ=�L��?�ƽ�Ȣ��	�-,#��S�?p
�?k�/��ɋ�tl��->hZ%?U�Ӿof�>��-Z�������u�e�#=��>=H?�\��f�O�|�=��p
?Y?7e�ƥ����ȿ�wv�j��>��?���?��m�d@���@�c��>ʟ�?�hY? ]i>�j۾FvZ����>�@?��Q?��>;��b'�a�?߶?�? �D>��?�r?9��>\V>�x~-��r��Ư��2Ӄ=�MD<��>҅>&���E�x3��3���<�e�k��f>x=��>�8��¾�=�=��W������w��>��x>v�C>H�>��?�v�>Ө�>��X=��`�����u���l�K?\��?��%2n� G�<Ѣ�=��^��&?�H4?jn[���Ͼը>��\?4?�[?�c�>���;>���翿�}��Χ�<^�K>�2�>�H�>�%���HK>�Ծ�4D��o�>Yϗ>�磼.@ھ�,��,x��C�>qe!?���>�Ю=Ƙ ?��#?��j>.-�>vaE��7����E����>���>TG?�~?H�?,Ϲ��Y3�.���塿)�[��-N>b�x?�V?�Ǖ>����Ɂ���xF�!3I�����뚂?�pg?Z\��?�0�?}�??L�A?d1f> ���	ؾ�����>/�'?���){4������x����>S�
?Հ�>g-������r��|0��D龌�%?J�B?C?�-�?_n�^z�� �=�}��7�9����Ks�W!�=p#%>�ī���=�C>$�����I���.�粗=�t<^r�>�9�=��p��9��$,?��E������=��r��DD��`�>�YL>����^?Dy<���{��ڬ��r���hU���?���?�F�?�l���h�g�<?�*�?�!?���>�����޾��߾��w�MKx�V����>��>�W�^�{����Z��bQ����Ž�K�n��>j�?�J?��> |�>VM�>ae���{��D~�x�6��BW�����5�C
�l�!�R�Ҿ��S�A��<��ݾa������>��E�#��>8?��)>�ҧ>q��>��O�)�>/�->ؑ%>�y�>�)}>6�)>�5E=�%�<��&�9�J?�k��C9�J��B����_?�Xq?X�>�N;+Ȁ�A���C?��?�n�?�F>�t�m#�u��>!�?�X��0�>|B0=A)�=�B�t�پN�?�|��� �<�'f>ẽߏ?��%H���@�j�?V$?G�`=�־�������Gj=��?�(?w�'�4�P�HFo�s�V�neR��#���sk�=u���"�$%o��(���>�����<C(��<=�#*?o��?FW���§��j���@���_>���>��>�f�>��J>C	��r0�4�\�:P&��{�?��>Xky?3�t>f�c?4p<?��(?tl?�?,Dk>�"��?@��=4wT>�W?�{B?P�-?��$?3	?c�1?�{>���;[��{���Q?q?�?P�>5�?
@�����:M	�/1�<�5��cս^>gG�=��录[t�/�< [V>�j?c���GA�Ź�%Cs>�x3?IQ�> @�>�zY�����=)0�>d�>*�Y>ʓ�K�>��X���O
?=q^?�$��<=qo,>s�=�����9�<�=jb��%�=`�L<"�߼�;�<В>��-=\�t=����<X� =�$��Lw�>V�?�v�>R7�>�=��8� ����ނ�=�Y>'�R>�G>8پ�|�������g��y>)l�?�u�?��f=��=��=Cn���P�����D��AT�<��?�J#?�GT?ې�?$�=?V#?��>� �	G��1Z������Q�?�9?�K�=RÏ�8���Gԯ�F�c�Ψ�>Q��>"+(��9>�Dd��[پȉ>P�>�K��:�Ҕ��ꃿ��N=��/�H����?%��?� =.�9���-�[b���Y���m�?qx�>�6�>/^?��j�Ne��;��|�>�� ?�fc?u�>+�X?��?;�N?���>S�*��B���*�������N>��E?F��?�.�?��f?��?��!>Wc���#̾(Ͼ�"��ɫ���삾˼�;��+>��>+�>�0�>�e�=�ӼO`ؼhF�^m�=��c>�1�>b�>�ȷ>Q�q>�q��t5F?���>Qa���n ������c�����}�s?M��?m�?��c=����K>��D�S-�>�F�?B��?/�"?tB����=�������v�����>y�><�>x����=�O�=���>p3�>wa�nB
�k?��g�<e?s�Y?�G�=�����:m�������������i���E��!m|�x�d�L�=�ZF�ۛ���{�.��pz��r���Ϊ��v}l�eu ?��J=㋧=1�=�F<Ė��7/�:��=�����o;nP*�"	�=bqR�Z��M�>��u=�=о:��V˾?r}?xI?��+?<�C?j�y>=�>F�1�ш�>j���dK?uU>[�O��p��|R;����������ؾiH׾��c������>҇I���>�x3>'��=t�<�Z�=�s=�0�=�`B�=8�=Zܺ=�M�=.l�=��>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��n>�@�Xm�H�A�ʛ��V��o�0�GW8?[�X�U�-��Y�>��=�'�s�&��j����ǽA�˾F �=����(�=�?o���k=XҺ�-kb>��y=஋>զ�x��=��=׻�=�e>yL8�.�1=����Ȉ>r{�=��>�3=P��>�I?�QF?i; ?#�?H;;;2��Z� ��)h>�(�>��>n$�>��>���>��]?�U?[�i?j,�>F�>��>T��>�:��]��&۝��M���=>�XKZ?�?��>;��Q��}ȑ�������6p�>B[.?}��>y@>�U����9Y&���.�"���\5��+=�mr��QU�_���Jm�.�㽹�=�p�>���>��>8Ty>�9>��N>��>��>�6�<yp�=�ጻ,��<� ����=4�����<�vżW����v&�I�+�[�����;���;��]<���;J��=H-�>��,>��>`��=]<��p�5>�G����K�1�=�J���A���]�J��)M.�[�>�ā9>�M>3q�����3��>�Gl>v�#>r��?��u?�-2>�����Ѿ}���My���[��<�=a>KM �3:�Qc���K���Ծ��>]0>��?�?Km7��2�U)�����&�+��IT?L��#w`��7�>/e��<q��:���B~<�Շ	�<jK?�����ɟ=�'�?��>^�?��'?5Z>�@ھ��i=�����
�������پ�m���>?���>��W>����b4�Z�˾�&��w��>9�H�R�O�@h���1�nEݻb��fް>�q���7ѾE3�5i��Q�����B��-r��ӹ>9O?=ή?+Kb��O���O��X�M~����?R�f?[�>Kw?�.?A���6�����ӵ=�%o?�h�?3+�?4�>�m�=�PZ=h�>��a?	q�?#��?��?�5�(�Y?�雾�s��Ƣ>���Ÿ>W�>-�i>�-D?+a�>q�5?\�P������������_����p��ԭ���? �>75>�0�=��k���=ǂn��n�>u�>|��>m�>��r>6E���
�|�0?V��=��>nq2?�e�>�/=R���f>�=��Խ$�C�{e�Jҽ2�ƽ뎒;D�ۼ�=P�%�L�>��Ŀ䠖?��5>e����$?p5��񘼂�L>�V>>���=��>A8/>c~�>���>��>%��=Ň�>o6*>�2Ӿ2�>���J!�9C��MR�J*Ҿ��{>q���%��x�����zI������M�c%j��/��]/=��J�</�?f����k��u)�����?p�>w6?Č��刽�E>���>��>W��Cf������Wv�%ŋ?���?�A\>Aң>��W?#?ڿ�fV5�']��u��J?�3�^�G�\�����f�|������Q.X?k5w?�<?���<M�w>���?.�,�Y����>�*�M\;����<�-�>Q���!�X��ʾ�����v�W�G>�n?�S�?��?!�R�!�j���'>Hl:?WZ1?7t?C�1?*�;?����$?�#3>�f?1?�5?<�.?T�
?�2>�B�=ᜏ��"*=bё�+���ҽIɽ���Q�3=>�=#�j9���;�}=�:�<���͂ۼq!;�]����<=�<=$��=Q4�=�>��?�&?L��=��b?l�=+O��~5��[?Iso>�ɽ#n=�R�!I���>��g?�g�?�?.;�>/�[��f����1>���>�&�=:t*=��>k�\�_%��D���h|�>8�>�G����ȼ�t�<���D}��T>�!�=*��>C�{>)���
(>ծ��k�y���d>ȷP�AȺ��S�P�G�y�1��Rv�$��>��K?��?;��=f!��약=#f��(?4?<?� M?8�?y�=܍۾_�9�(cJ������>|��<-��G������wi:��
�:A�t>c����Ҡ�cWb>R���r޾��n��J�n��l�M=s~�avV=w�(�վ�F��z�=;
>ճ���� ����LҪ��*J?-�j=(v���nU�oc��I�>μ�>Y�>��:�!'w���@�U����G�=ε�>��:>
�����wG�h3�,�>�Z@?�a?jf�?* N��d��'�L�	�֑�\� ���?5n�> �?^[>J�=�땾����|j���J�Xc�>m��>t+�]FQ�����I��.y-�Q\�>�'?�\%>��?��U?�?qOT?��?K0�>��>Ί�o=��R&?�2�?j��=PUϽ��O�ԕ7��%F�px�>�1*?m�B��1�>��?h^?�6&?:#P?v�?nD>�1 ���@�\ە>��>�W��u���^>��I?�Y�>�UY?���?��@>��5�i��z�����=<>̱1?�}#?58?��>P�>L���ZZW=c��>,�`?+��?�uo?>O�=w��>�%>��>2y�=W��>���>?_�I?�zt?
wH?BZ�>kٯ<+���4��������W<�߉<�p=n�
��)z�X�#���<\S8<���{߼�g
��S:��H���5<�5�>!�>Eɽ�"�ǼH�HI��PsM=�u>����I�۽�r���	>?�(>?j>E�>wb��������>��>�D��S�>�9�>� ?(=�=��H�
Eξ�LJ�,5�>O	Z?2�>?B�6l������6�=���?�rV?̩�a���b?��]?�g�=��þ��b����+�O?��
?��G�y�>��~?��q?��>O�e��;n���\Ab���j��̶=�o�>�W���d�c@�>��7?ZQ�>^�b>"�=Mo۾��w�Pl���?�?u�?���?8-*>�n�3��o��jO��<^?ڇ�>�5��N#?�t���Ͼ).������ᾕ4�����d/������.Y$�mۃ�c�׽8�=�?g	s?QVq?x�_?>� ���c�-^�o	��aWV��'�o�|�E��,E��C�Y�n��d����*����G=!VJ�!���y�?FYF?O�R��O@?�������&�ѽ�����м����=�v=�J> ���}�>�Hx=��]	�d��>@�?f�u=sAM?��-��p1�4���0Z��1��J 8=��E>F	�>��>�Z�=�ˑ�Y�����1<�W-���p>�hv>b?�H?��l?p,
��0�����d��a�ԥ����4>�

>��>�[�ʵ�%)���>��)p�_�
����A	�vOt=��1?�R�>�G�>i�?��?�y�0Y��6:p��J.�|��;�>�>Cpk?z4�>�>�M׽,� ��d�>��h?���>1P�>�%����!��~��(�����>j�>�.�>��m>���Q��5��1���L�<��&�=m?�����`�9؃>IeT?�*����;M>�>}\��B��l��mU�I��=��?�5k=�o>˾��Jr���{��L)?�?6�t'����>~$"?��>��>�C�?_7�>�������;x?7�Z?�kF?w�@?���>=�*=,�ǽO9ҽ^�#���)=K�>��T>.x=pl�=IW��g���O�E=�==�������\<y���H�; $�<��6>�'�l�Y��I߾����!K�ڐ(�ߙ�����s��e%_�ؖƾH�C��[M��"1�����tže�Ǿ�qt�F� @�@o9�����_��=������X?z?�R1��ٖ�d�T�����l��ϕ��W�ID�_�=��bl���%?a򌾣�ſ�ġ�.+پ/�?��?�dy?)T�����9��->)	<�d�㾰���zͿ�&���x]?��>��ݎ���e�>fNx>|�^>0ۂ>ጾޛ���x3<hZ ?4^,?l�>�tM�Pʿ컿Ce":ē�?Ũ@'�@?^�'�i4�fvq= �>/�
?�C>�n8�Y��DԳ���>j��?�Ŋ?�[=ϥX��M߼q�e?�t< �D�m���b�=�&�=��=J��H>���>����9?�b�߽dH0>t��>%M ����^�)��<�d]>�Uս�"��4Մ?){\��f���/��T��U>��T?�*�>S:�=��,?Q7H�`}Ͽ�\��*a?�0�?���?'�(?6ۿ��ؚ>��ܾ��M?ZD6?���>�d&��t���=�5�j�������&V����=_��>o�>��,�����O��I��a��=��`࿱�G��4�~�=��C�֪&>`O��������پ|����tq�HyF�1�2>-�>]�;���=��>�U?�ZI?�ޑ>�%>飛�a�C����DU�����^��t>S��
������L��R������P^��r�<�bØ=-�Q�H��w�"���e�hzE�LT/?��">�5Ⱦ�K����:�t;�g��J�v����aɾ��/��#n�b�?B�C?�녿��X��%��s�3��(�Z?�����@�����=���T�6=���>'<�=&ݾ��-�6R��U?���>B��ƣ���Q=НR������V#?d�>��%>E�A>��&?C8���w����>��F�>�L>�!>�j���������>�>?ʪܽ�M��x>���0'�=��
>�>30b���&�8�>f�콁Ρ��PP=�m=�P���� .?hȰ>��4��I�_��)��ꑽ���?)\�=:��<�7b?�%?24���-�����a&�n_潨��?��8?�Y>W(>�E4־w_����(?�%�?C">�J�Q�=��V:����GX1?�kp?n�?�K�=Q~���Þ�L�´9?��v?s^�xs�����O�V�d=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�%Þ?��@���?D�;<  �T��=�;?l\�>��O��>ƾ�z������+�q=�"�>���ev����R,�f�8?ݠ�?���>���������=0��0�?�Q�?����[>���>v�����&n�i�*>l���J1(�� ����P�y1L�mi��@¾������>�@Yr�����>�1��<�Կ쾿&Շ��p׾���?��>���>O"�=''��o8U�O�b�2�4��&�-m���?p>Ɉ�>f���0Ⱦ�r��Ov�x}��a? \x��iO>�q�����iV �_�=��{>�x�>ǰ�>Y�0>�tѾge�?��Ծ�Rɿ%1��a�����?h�?�B�?�f�>�Ȑ���-���w�U=o�h?��L?ד<?�f��t�=�.�=�~j?]ꩾ
-`�	�4�ME���T>��2?Hd�>�]-��+{=u�>u��>�>�6.��rĿJ඿�����٦?[V�?�f꾁��>�A�?C<+?/I���}��>�*�2�:B�@?'y0>����6� �~2=������
?��0?�T�C��X�_?�a�I�p���-�j�ƽ�ۡ>�0��e\��N�����Xe���Ay����?I^�?`�?���� #�Z6%?�>`����8Ǿ��<���>�(�>*N>�G_�j�u>����:�'i	>���?�~�?Gj?���������U>�}?��>�5�?ג�=��>�B�=�ʵ�CɼGP4>���=�&�5Y?��N?�|�>Uב=^#��1/�eG�%�N�;U�A|B��>�Q_?1�K?dQ\>����F�7��<!�$8���2*�l����>��x��9׽�;3>��3>�+>�US���Ѿ��?Lp�9�ؿ j��#p'��54?.��>�?����t�����;_?Oz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>E�Խ����[�����7>0�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Fa~����7���=��7?�0�I�z>��>��=�nv�޻��G�s����>�B�?�{�?���>�l?��o�N�B�i�1='M�>ɜk?�s?W[o���|�B>��?/������L��f?	�
@zu@_�^?,�nֿ�����U��b����=X��=H�2>�ڽrG�=޲7=�*9�͓�`��=��>��d>	q>:O>�`;>��)>����!��n��ݟ���C�E�q}�C[����Cev��}��5����������Hý{_��I+Q�C&�~.`���=^�T?�P?��n?H�?��=���">�� �@�=0�&��-�=-�>�L3?�K?��(?.��=����7/d�D逿Zl���������>��P>���>���>��>�Э:7IA>��8>�x>�>��=�� ;���<hL>�M�>4h�>��>)C<>t�>@ϴ��1��Q�h��
w��̽(�?���� �J��1���9��֦��dh�=Ob.?�{>����>пM����2H?!���b)���+���>|�0?�cW?�>���r�T��9>տ���j��`>, � �l���)��%Q>ql?毃>BAp>��$�x�/�=P�����6G>�1?���4�׽�j���G���q:>��>�u=N4!�:���~ي��n�<ŖM?�?�Wh��ǵ�d����L���#�>�q>0�8uMQ=|}>й�r����?6�xm�;L�=KI>��?�nK>ݜ��H>ƛ��Uc��!>���><�m>�!4?t+?e�¼�g���o��ӂ�D1>j�>
��=�d���P���<��>K��=x"���$�n��PHf��]�>C�=r���%'M��Q{��C鬼,q�>�c�Z�,�|}m��~?���(䈿��e���lD?R+?d �=��F<��"�E ���H��F�?r�@m�?��	��V�@�?�@�?��H��=}�>	׫>�ξ�L��?��Ž3Ǣ�ɔ	�1)#�iS�?��?��/�Zʋ�=l�}6>�^%?��Ӿ���>���D��?���v�J�=�>
�H?5���j^��U:�u�	?]?��vl����ȿ�Fv�}��>�x�?^��?��m�;/���1@�w��>4��?=�X?cj>�N޾<B^�=�>�6A?ҠR?;�>z��"z)�H4?g��?ì�?�!I>jU�?��r?"W�>�N~��K/� ������`�=O	�;u�>@h>�o��!�E��u��+����j�4B�޽d>g�"=\c�>Lt�g���w%�=
���ݧ���g���>�Kr>�hJ>?��>�~ ?Ɉ�>ju�>�u=�1���{���ϕ�l�K?㲏?����1n��G�<��=�^��%?wI4?�C[�w�Ͼ:Ө>��\?���?j[?�e�>����=���翿%�����<u�K>�7�>)G�>P,��FK>X�Ծ/D�nq�>�̗>h裼GBھ;-��s����B�>qc!?Ǐ�>�̮=� ?�#?��j>��>z`E�8����E�{��>���>=J?��~?>�?@й��X3�� ��桿��[�"CN>�x?XQ?:Õ>��������FE�GVI�<񒽳��?�kg?:彈?~0�?��??��A?�/f>�l��	ؾ������>��?�6�k;������]�>�W�>�f�>��0�	�ѥ}; ������>�i^?�"?����C�Z�J�Y،<ƨ��_��eR���޻C�>5>e����b�=��>��	>;�m�0&S�qmS�*q�=:�>V�>[�4��f��<,?��G�vۃ���=J�r�_wD���>NJL>���T�^?ih=�=�{����cx���U�} �?9��?�j�?1��N�h�W#=?t�?U? #�>�H��}޾��ྍTw���x�!x���>��>�`l����������E����Ž�����>y��>�?Q��>��M>�P�>vk���<&�*X�ܣ���]�1+��98�8k-�P��9����#�a����
¾L�{���>�
�����>=
?zTh>3%z>=A�>�A���b�>��Q>�M}>���>�Y>��5>��>A.	<��ҽ��I?؍��Wl.�[���ھ�]4?��S?�?��;��ъ�N�ཱྀ�?���?��?D�>+ai�G�:���?�F�>�i��q�>�{�<�1C;n��<�������Π���2i�>�m�.���>�|=��&?%?�m����E[�신�Q�n=�M�?��(?��)�{�Q���o���W��S�ݘ�'7h�j���$�ϛp��쏿�^��%����(��u*=��*?\�?ǌ���!���&k��?�|df>B�>~$�>�߾>uI>o�	���1�0^��L'�����XR�>}[{?%|�>N!?V�5?vt?�y?�?��-?��3�o@?���=�<�t?�
Y?�G$?���=�w$?_2?z~!>�.�<l9$� ���?��b?�+?P&>��%?o,��=������np �2렽`�>iiT>cW�|4��x��`J�>�-�>���=	�,y�7�<6(�>y�W=�7?� �����<�(��D�?QSP>��>�Z�=珿���A��>B�a?'-��{z���>ǠR>3V���8c��S���$��)�>�4`=�ü�k��%w>]���x2�������0��P>{u�>��?���>T?�>m8��&� �^��Pv�=WY>�S>~>�Dپ�|��d"����g�<Yy>w�?w�?wf=|�=��=�~���_������������<Ѩ?�A#?
OT?���?��=?Bl#?�>+��L��^\�����?��+?x��>��x˾�ި�~Y3��?�x?4&a�f���)�D4¾�Qֽ"8>~�.�S�}�A��� �C�������e���'r�?	��?0�?���6��+辚���|5���C?aG�>Z��>ތ�>�)�sg���/�:>���>|rQ?��>��O?�-{?��[?�V>��6�����7h��)� >0�>?�F�?��?%Ex?��>U#>U�$�W�޾����� ����1���6K=Q�Z>��>���> ��>U"�=Aǽq���"�9����=J^>!�>L(�>#�>�y>���<q5A?w��>2X��3` �2ƒ�a�y��G����e?�]�?�G)?]�>�L���Q�����e�>���?=��??<���k;�=��1��[ľ����D�>A��>�s�>��=�����O=�w�>=~�>��������Ԑ �򝏽��	?}??�=�t�餚���
�໸��*H=�椾�*u=X���0��u>� �m\�ܑ�?�;�YP����q����ţ����dL�>bb6=:l5>�^2>��=������;H6��/����>K�+> �ֽ�29�LM�=�iS����&��<L�z>�Z�<�8˾�s}?I?fk+?%�C??@y>��>J�1��t�>�z���2?)rV>�8O�b����;�䫨��@����ؾ�@׾Md�#���&A>� I��h>�3>c �=��<w��=pr=�֎=�F� �=J��=}%�=E�=D&�=Y�>�<>�6w?S�������4Q��Z罞�:?�8�>^{�=�ƾr@?��>>�2������~b��-?���?�T�?9�?^ti��d�>O���㎽�q�=,����=2>w��=[�2�-��>o�J>���K������4�?��@��??�ዿǢϿ9a/>,gv>I��>Y1G�q�5� 伾�;�$־�@J?���bc)��a�>�ͽ��̾6�1��[?}�{=��:;�7>�/��W�꿽��ӻ�$��G�>�p2>���=��=/����D�=D%��|K>�1L��>Z��T����=�Y�=��	>��>��?|)?..w?�?	}=78=��$!�� ?:��gt>�$>=�>2/�>y�>~�Q?
WS?7b�=�ye�r�>Y��>^�w�����ʾ;df�����oh?�Ȅ?�W�>��������� ���2�3%R�>y@$?��.?���=��W�~h1���5��rν7�<�6b>5�v��c�����{��ܸ���`�=t�>W��>�6�>��?>�@9>0��>A�>�3�=sK><<�j=��<��>���<�����T�ԏ�ī'�����w�=�+=����e-/<��1�_�_�2H,=a��=1:�>�&>�\�>�=�ӳ�",>�	��,�K�%�="����A�\d��~��c.�QN4��xA>��V>����H+��I�?n�]>�m>>C[�?�$u?0�>����վA0����d�&�S����=�
>��=��	;��_��M�p^Ҿ�i�>%[�>�j�>�ft>��*�U�;�P��<��վ$2#��J�>������f�����sn��I��A��MRi�O�\�]�9?���@b�=���?��A?��?m^�>�JU��\ݾ��)>m�m��9�=�F��^�;�ɽ�Y?W�,?�$�>�a���D�5��[6żmq�>6>[���e��꯿N ���=�¨����>>�F�ed�vc<�(��t���<I�?wQ�h?�>?��?ѣ�=��r�pKq��Tf��U��#?�Ӕ?#��>�>�?�Ž�����Ž�?�>^�y?`O�?q��?�ؗ=f^�=�g*=?%?��R?֞�?[��?A΍?��^{�>�L�����<y)>{��>�*�>Q� ���~>��?�R�>�+A?G�ֽ����ľ�Z��^7f��8��,�F>�m�>��M>cw@>8L�=4�=�wl;�>�ݔ>PA�>G�>a�>Hw�8We��H=��;x?h�9>�s>��3?({�=������>�(>YU>Zr��{=��<�-��l�>&�A��������=]Rڿ���?��M>�ᠾL"f?�j�ڋ?��i�=�W��Q>A�>r��>L��>A�T>���>�˂>^�;=���= �ҾK�>+��<�!��C��IR�l�Ѿ%�{>�S��`<%���4��GqJ�Ҵ��
�*j����ʏ<�Z��<��?����`k�3�)����C�?#��>8�5?#�������>�"�>���>����њ���፿���?��?��b>XB�>Y?bZ?d�+�H�)��KZ�r�v���=��Hd�^��^������D�(�ؽ9�`?�Cz???�2�<�
{>:�?XT(��˓��ˎ>	=.�[q:�=RX�>߽��jAl�k�Ѿ���/�!�˒A>ىl?��?A?4A�
}��Hs.>�A?�IT?�3�?�@?; Y?w玾7�?���ż>=y?�:>?�4?�,�>��L>_�>	%�mn>g�Ƚ��x�����k��c��"�v=�ݚ=��k<2.�@�;=?=�)/=K���Fj8���<�u�;d�E=��)<�7>yi�>�T?���>��>[F?��a>y���('�9�F?ڢd=���қ���U=�o���$Z�'bf?0��?�<?'S�>�M��-V��<w=� >v��>��>�	�E������W�>�9�>��=>���o5$�>�վ�����L >��+>R� ?�GP>�S=�pH>���6��X��=�l&��IO�'@��:�<��Y:�� �����>#&+?]%?XW�����I�{��Dz�˴�>'/w?y;U?]Ă?���=+[�!�C���*���#����>�`����� 6�����������.h>��ľ����!�b>��ׁ޾�n��J�j��X�O=J-�lbX=-�ܢվ�\�N�= �
>Ģ��+� ��������J?��j=oc��}U�TT��i>�՘>��>�	;�;Ww��|@�zy��v�=t��>�!:>F�����G�y�}�>e�7?�Hd??D�?�%��D�F[(���f�nϽt~?ģ�>R�#?4�>��3�[���A���i��e"�%��>Q�?�A6��|j��Rž�
�Ļg�q"�=���>�%>ƙ�>��'?���>a�)?�7?W�
?d7�>��=�|ľ��(?|�w?)6�={&���c�1�'�{N����>�XC?~���ܚ>hv?��>~a�>�]?%&?t>����R�/��֗>3�>��J������>r?j��>`�]?N�t?Q�'>�AL��ʏ��ʾ��2�=��=o
/??���>���>`��>�ܠ��y=E)�>��b?B�?O�p?���=Oh?2>�m�>�ɛ=Y�>o��>��?a�M?xCr?�0K?� �>v��<k���TJ��n\n��Gܻ��;#�m<�,z=Y������B�(�(F�<E�<e���)S��$���=�7���>;w��>
��>�;��|M�s�.�����D���>�o��ɓ�f�=�7�������>�	?�מּ�)�>Na�>a��>9��	a?-l�>�??X�<x��̯������6?qG9?U	�<������@�m��Zo=�.v?���?�0
���۾D�b?B�]? g��=�G�þT�b���L�O?��
?�G���>��~?)�q?q��>N�e�a8n�:��$Cb���j��ж=3p�>�U���d�@�>ޙ7?uK�>��b>��=�w۾N�w�Kn��T?e�?� �?���?�"*>-�n��2�D
��	p���M^?�>C���y�#?% ��ξ�Պ���u�߾k���p�����.^��?#�w��ysٽ	��=��?^s?:�p?�D`?ݰ � =d�h�]��1����U�-.�\��^�E�sE�T�B���n��t�����"���=I=�i���K��)�?��"?�!�0�?���{ؾ ⽾���= �7��0����=��(� �üZ��=��x�YJO��d��?��>�؛>��;?E�[�9�<���&�Yq:��z侪�>-�>۲�>}r�>�p�<B�U���߽��|���- ��G�v>Cc?uL?��o?
��x@/�7Á�=�"�,�;�&����L<>Ns>	6�>�J��[�f%��">�~vq�G��C����
�C�=�m3?�d�>���>p��?��?�	�n�����}���/�}��<t�>�vh?���>���>^7׽�d!�!��>:�l?*��>Y�>���HL!�x�{�rʽ|3�>b�>�i�>�o>��,��\��\��z����8�D�=1�h?�s����`�Bڅ>��Q?W�:9I<̀�>��v���!�(��@�'��>Ir?�ժ=k�;>��ž����{��6���m(??ڍ���S%���J>�a?��>?c�>��?s��>�V޾�[5;#??�I?W::?e+?y��>b�<��Y��5������ =uNR>K^�>�΂=X��=�۽'�s�avO�m�?=d�=�.!��l�f�n��}��5�#�<0�>�F׿��N�ƃ �k�n��eپ�:��.'�޶�����
��;�Q�D/;��J�����J���<N��p��C��?�	@')=�s��OJ������$}�g
?��+�dy�=�祽��k��R��U�D.'�G�&�F�N���c��⃿+z ?*����rſ๓�Xz��_�?��!?�6[?2�Ҿr�lG9���m>�r;>��Ƚg'���߃�\7ҿ�I�Q�c?���>�پ6�o��{�>�ǐ>��1>:S >BdY��֔����<�-?�#?P��>�]¾CϿ�u���l�=�[�?�@��2?%�R�_�Ü`<���>�$?'��>�Ͻ�s޾�A:�M�>��?=�w?y&�Mg�k�>�?�憽4�پ��K=�-�=�j�<��"��8���Kw>�r�><�7��y���f#�4}>�d�>�E����M��X���<珷>r{>��4Մ?*{\��f���/��T���T>��T? +�>K:�=��,?W7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�ޅ�=a6�����{���&V����=Z��>i�>,������O��I��`��=�,
�N�ѿ�����%��!a�6=h=�$������c����fT1���=���>��y>�(=���>��&?�<=�5�<�S?��=?(�>�>HS��Σ��TȾ�-5�4��(߾��½�e>)�½�0����	��=�����$v��x�
��u<��[�=��N��o����*�bc��GG�S(-?-0
>�˾+�C����<��Ҿ�C��_��4��v\��T-+��~�h��?�<M?n�v���Y�"3��!̽eUнK�f?x��s���<��/�b=����%р=���>FG�=6!쾸�$��N���?�?�v.������)���wjk<�1?��	?H�&>'�6��?��8?3����>��k�i>�>���=�-�����<)�>��0?3��[s��d��> �k�.�O�oԋ=�k{>����2*W��-�>��{�=&��M����&�¼<q6?xo�>d��8������6�/��I�?*n�>)��>��\?o�?Q9� Ž�������Lu=?�x?�o/?IS> i��7\�������xM?xe?�>I����6��D��z־2�?�QY?d,6?��=^ׁ�<0���t����D?V�v?kj^�Ip��i��u�V��!�>�O�>���>��9�=l�>��>?r#��H�������M4���?��@���?ܓ;<)4�y��=�9?�a�>�O��@ƾk~��"���ɠq=�%�> ���igv�3���\,���8?��? ��>و�����8�>ͳȾ�ɰ?�E�?�c���}>���*�G�p����%��&8�>�����ר<H6�$0i�-E�����q��Y8)����>, @�0��t8?�Y�����¿0��exľ���yN>�`�=Si�=��9���=�B}^�=����:�"�'��5>-(�>`��_޾ǚ��5�e��Y��e?����
�>V����Ǿ���7��FY�>Z̨>�]�>>h�=X�W��*�?z������Eа�oE���*?3m?��?�M�>�o�=�4�4'����Ae?*H�?�/I?7�����>`�|>�h?�2��[2c�&�.��s=��EZ>?B?�g�>���A�>0>�d?m$>�C��ĿI*�����\�?�]�?oAܾ&y ?I]�?I4!?��������������=wi@?G�7>��-/-�Y�>�����S�>ݕ!?(׀����4�_?ƚa�"�p���-��ƽ�ڡ>T�0� e\��T�����#Xe����Ay����?+^�?X�?7��� #�\6%?�>p����8ǾN��<倧>A)�>�)N>�F_�9�u>����:��i	>s��?�~�?*j?��������V>�}?>��>�C�?j��=r�>S��=���	�:JH>��=�c!����>�GJ?Y7�>{��=B�*�pi0�oD�/T��g��A��{>ZLh?'�O?w>Y>����o\�a�$�p`��C�x�����W��z��t|�g�&>�A8>���=�x;�iEؾ)�?��!�5׿ �����J1?��>�>���|BZ�8nԻ��\?�m�>��#���U��o��� �?C��?�	?�lҾ��0��F>�Ș>�!�>�/��x3}�đ��>)>�_C?�H��̌�n�k��E{>�:�?��@[Ұ?q�a��	?�!��P��t\~�����6�V�=��7?^%��z>���>HL�=�nv�ɺ����s���>?�?Zz�?���>�l?U�o���B�H�1=(X�>ۙk?�r?K4r��	�{�B>Ԭ?Ѱ�����NE��f?��
@�s@��^?HT��T:��m���S����my=�=��C>\iA�H�;i�O>U^�=0�߽J�=��>(.	=��>��=HDO�|�J>c����#�d�ÿ�<���S�����q�վ����\��μw�I�޾�؝�x�Ǿ�4~�c�=0�䇤�e�����4��=��N?��Z?m�?�?�}�}�?>5���f���{��h���w>C�9?�ZX?O�$?���=����]8Z���e��٨����Y��>X>�B�>�>w_�>�?w=��i>�;<>�r>��V>���<��s�;�7;>Y
�>Q��>�+�>�D<>�~>ϴ�0����h�w���˽[��?�z���J�N1��x-�������n�=a.?��>?���?п���0H?+���1(�~�+���>Ѽ0?^W?f�>���ږT��,>*����j��@>IP ��xl���)�$Q>ml?�@�>��>D`���1��F��Ѿ!m�>��D??����0�Rx�^�+��۾ձR>]ƺ>?���3w�ʖ�l�s���i��&=��L?�c?n�������`t������)�=��>�rV=��<��>�V��b��8�C���Z����=��#>�[�>Z�v>���=C¢>Ů�dM��Z��>�i&>��?|�T?E��>rI�;J�
�H���K>qm�=R=>�Z�>xף��hͽ6YY=J�>��=�����\=��K��?���z>u�\����/�vs�=Ne����>�)">_q�=���������~?C�� 䈿T뾖[��2lD?�,?I��=��F<L�"�Z���A����?��@�l�?��	��V��??@�?�����=�z�>�֫>eξԙL�K�?p�ŽJ����	��2#�Q�?o
�?�0�>ˋ��l��2>�\%?�Ӿ}��>����\���ㆿ]Iu���#=���>��G?����MZJ���=��i
?v?��%�����ȿj�v����>v�?t��?X�m�:���v�?�g�>���?��Y?��i>��۾��Z����>у@?B1Q?���>9���&��O?��?R��?I>̋�?��s?\i�>�)x�;T/� 2�����U�=�];M[�>
:>]���vaF��ғ��c��f�j����u�a>��$=��>5佃1���G�=9܋��?���f����>~q>��I> Y�>$� ?�^�>���>bN=f���݀�������K?䫏?O���&n��l�<rP�=U^��G?�F4?�^���Ͼ��>��\?̸�?f�Z?��>h��9���ӿ��c���~�<,YL>�=�>:�>�k���K>D�Ծ�D�!T�>߮�>c��  ھC'��'՚�+	�>�L!?�>�>�+�=�� ?��#?��j>��>�`E��8����E�f��>U��>K?��~?-�?�Թ�Y3����㡿��[�-5N>:�x?�T?�ɕ>Ǎ�������XE�J�I�������?�ng?}S彺?�.�?��??�A?>�e>��� ؾL٭�g�>o�?���'O����؏��8�>��?���>ؼ��i;P���zա�Ң2��<?�]?��?��0�@���`ǃ���/=��F�� ��T�<����Y�=[N	>�}�<{�^>\��>(�l��3���v&��$���0�(��>��=p�D�� �	),?�U?�~؃�p)�=��r��D�7>4�L>���ޣ^?ͱ<�N�{����km��UpT�6�?a��?�Z�?����xh��=?��??�?-�>z﮾{5޾u�p�w���x�]c�e�>���>��b��徍|������9��s�Ľ ��	�>YZ�>�'?V
 ?��V>���>}���4 ���뾎��b�Z��)�n2���)�v��m��96�Q�A�������z����>��Є�>t	?�*h>��w>r9�>·ͼ�n�>RBh>�*n>.��>�^>�>�~�=��<^��%�;?o���W:���Ӿy���Z??�c?9��>���䢃���۾itV?	؜?���? ڿ>0=��KV���>:p?�e�LB�>���ή��ߑ���ؾ��=�+F�>�[���?v�K�yG�h����o���?k�?�Z������J��&���1�n=oM�?��(?�)���Q���o�|�W�KS����4h�h��e�$�Ϛp�폿y]���$��Ǣ(��~*=��*?G�?׌�����"��&k�?��`f>��>P%�>s�>%rI>l�	���1��^��J'�ɶ��T�>-Z{?��>��E?�VS?7'~?V;v?%��>���>�D(�/��>i�ܾ��&>�ē���9?�x_?�Z>���>�߲>��>���><�ݾ��%?��*?�6?�?��?�k��w/���(@��29�V@�=퍴=zȗ>��޺u���ؿ�Cj,� Ud<4I?rJ��(	N��ؾ��G>��?��)?�ɵ>߳�<� � ����&?��>�@��������[�d#�i�?��a?�+\���<��U=wژ=2.�=��<���=�=5S>,v�����/~ <���=i����]=o�:�`�=+n���L���N�>��?o^�>�ֈ>������ ����Zı=�Y>t�S>->��پ3s��M���jg�� z>+u�?�C�?�f=��=�&�=����*���d��LV�<�?>�"?T?R�?��=?�#?'�>?�4��jS�����q�?׍.?Ȝ�>�p�����-z����5�`�?��
?N7^���ֽ�+��I���Ѭ�k�>3�#�(R|�ɬ��}F�a@&�K�Gqѽ���?���?�JY��u!��n�Μ�Aʾj�A?��>M�r>�	?���n:j����?�=o�>��9?I;�>{�S?TS{?c?]o�>���]J��+�����ݼ�9�=�^.?_�J?���?�P�?٭�>eD#>�t����C;¾��W�;���\<}��} =W�>�&�>�6�>�Ջ>�{�=?�A�P3C�@�r�ls�=G�/>��>���>)��>yw�>!�>Z�?�^?��� V�ޙ�?�,�1����d?�_l?�A6?�O�>o�C���l�c�%��?ά�?��?�:
?q!����#>	��b�������)�>e�>�d�>��b=%�8P>{��>c)�=��=;���6.*��i�Lt�>�?$�;>���� �����)�����Ž�4��U�D�A伾�@Ľ�?�߮�1�S��/W�����-���.�&��Δ㾐�x�w4�>j��=���=d�?>0�ĺ�J����r��_Z=>ڽ�þ��<��=�11>	�B��'�_>���=^�a�H-ʾ;(}?�H?t�*?VDB?=w>�>�v(����>�?��s?$�R>��`�vL��=�:���������$ؾ��־��b����*S	>N���>�q4>*��=�m�<���=�f`=���=��9<�=�U�=F8�=W�=F��=�<>o�>�6w?N�������4Q��Z罉�:?�8�>�{�=��ƾr@?��>>�2������{b��-?���?�T�?<�?Gti��d�>G���㎽Zq�=���>2>���=p�2�<��>��J>��� K������4�?��@��??�ዿɢϿ[a/>�+4>�ϰ>�	���m�Z(�����O5%�
{u?�E��LA���ƣ>��?�{K�ZI��D��>Ri(����=�}�>�?�ح'=Ƞ�^�=��!>�>v?�>x] ��ݼ
�2=�*����4(>s�5>8�B�S��<;���I��tF�=��>��>��?��(?�{Z?U��>�N�j�ܾT�>���=�S�> �<ѱn>k�X>a�?��N?��,?��>���;��>B9�><e,�Cz�)���W��p����j?��k?|Գ>`��}֏�_��_*��b�=J?�s?�q?���>���k࿓M-��E/��d��?����k�<Wt���K���k���6������x>�d�>9�>MΤ>�k�>��6>D0T>��>4�>���<�P�=��<y�;1���/�=������x���+�<%u�<�u��٨�e��<O��<ǵ�<N��ƚ�=a��>�>�5�>�<�=����.>nE���xL�ue�=�/���B� d�~��.���5���B>2�W>3������j�?_cZ>Ŕ>>Gs�?�:u?Ek>�i�	�վ�@����d��CR�o�=��	>Tl<�؀;��;`�m�M�PhҾ��>	!�>���>a4�>L�2v1�'#=�;���F��}�>k�`��'�F}���>@�I����s����r�ʽ[g�>u����#��{�?��Q?m�?�)?U�7��ٶ>a<��#�u>c�5�j���o�|=&͇>ț5?�b�>����c�g�ʾ�н�¢>�UD�PN��̒���+�|�F�m�����>X���c���}h.�l���'����A�2sW�g�>�<?|�?�����k��M��Y!�˺�*�?�^s?h/�>�?�}?����6�?�k���>�`n?���?D��?�^�=�,C>����?�?�g?�,�?�w�?٠�?U�	�Ҥ7=����p��G >��>��>م^=Ö�=[�>�46>�h?�}���"���)(��꾺�[� "L�#"5=M�K>�p>�F>��f>F}>'!�=�\ӽ�">K�}>}1�*�"<��.>]�=���<�S�?	U>�ȸ>��M?����>�, ��أ�w�>ǿ��>�`�='Rܾ�1>�Q��0�;����^>	Ͽ���?�3�~���qva?�A���K>�S�>�׼b_>1q�>�u?>	4>���>���>6<�=���>���>��Ҿ�>���t�!��C�9~R��!Ҿ�}>[ל�i�$�l4������KJ������i�W���k�;�.>�<t �?���D#k�*�����/�?�g�>7)6?���������8>]��>42�>;����/���ƍ�n$�*:�?���?Pb>�1�>`W?*�?��5��f:���Z�w<t�e@�&d�n(_�"����偿�����_?͈y?I�@?��<��x>�F�?Ď$�)}���P�>i/���:��C3=y��>���~�\�)�վ��þ7�'G>фp?�Ӄ?�,?E�W��c��a>��@?��A?UŁ?U�9??oH?@G���%
?���=��>h��>��6?�a;?T��>���=f��=��c�>U����g���շ�ۄD�4�<�b�=�\�=��H�����P���4�]=�6;=A���9=��2<v��;�U�<+��<+g�=w˻>-�c?B��>�`�>��
?%g1������؟;?��=-�i�]�����`�����t�=�6�?Ү�?�!?�ȡ>�����=>-2">`6>�,�>���>�����Q��%��4�=���=�:X=�Ƞ=��%�� �����p����>���>��>NV�O�(>�ã��W��ڡd>�Q>�Y>��a�C��F�!�.��*g�!F�>+H?��?��X=��c���3 f�yO!?HsB?��P?**�?�I�=KG��?���L�������>{������$A��c�����4��fs���w>}騾������>[B���ؾՋ��@z����Ѿ������]�9�d�	��������i�� �^>2�E>��v,2��L����¿'[<?C�=>������&z���o8>^J>!?��ۼh�(���3�O)��Ҁ�=�T>?>,>�U>$����9��(���?�>�	9?��a?��?Y�C��1M��D7�X�"��c���f!��G�>��>��?�k|>[6｟��6U龡�W�ǳ��b�>M�?=u&�Im�V��MUq��"+���=Ht?�z�>t_�>e8??# *?:m?
��>��H?+�>�`����վeB?��a?ɽ=�%F��XȾ����7��??n��>2�U�_|?>�0�>�I?���>�?�>�q�=&���� �sc�>!�M>�XB�_گ�g$��(>?3u�>e�k?@?>��>���H���א�8�U��uB>��;?n?*�?wB�>���>8��`Q=��>Y$e?�?�?̛u?���=X��>�*>�v�>1ѿ=���>2��>�S?�rM?�q?��O?$��>�ף<~����c��bYn�*��k��;[D<��n=����]��.k��I�<�PV:H����Q�D����RA�Z�Q�A�;���>eWt>2;��\A->��ž�o���f=>"y�q������q�:�ӈ�=��>� ?Cg�>7!�'Ð=�M�>f�> ����'?S�?�?��';;Vc�xfپ_N���>�B?u2�=��l��f���u��xp=�*m?�q^?�G\�����V�b?��]?�/��;��þ�#_��D�FEN?h�?�EL����>E�~?^3r?��>!�h�7l��n����a�o1l�@�=Ϝ>���C�e��Ü>��7?��>�ac>1�=پ��v������	?�M�?��?\j�?�(>Q o���߿���UZ����^?/�>D��O�#?��Q�Ͼ^����܏�f�ᾉ���a���U���ç�a&'�����Dܽ���=I=?�&r?�q?F6`?�, ���b�*]������T��e�H ��YD��E��HC�X�o��L����w��4'G=��@�gMV�)��?QB?���Z�?1���u�儾�����θ�Ld���D�=�>!p����Pv����m�ľ�~�>�`�>w�>�eM?BH=�~O���~r1��({��뛽
^>�c�>��>�廽mvϾp&D��3	��uP�#
C���v>R`?�9I?�sk?�%	��Q2�I����Q�b�B��`�F>�|�=���>YtG��
�1k$�8>��?t���sF��*	�k�=�{0?p��>ߐ�>k��?_?gJ����Ӑz��D1��4�<�Q�>j2b?�>J��>�"˽2�����>�Tl?���>�8�>�Y����!��#{��{½4��>Ϧ�>�1 ?˰n>B.��[�W鎿����o7����=�tg?�턾pa��H�>I7R?�֟;�L<�#�>���,!�����t�'���>]�?�Q�=��=>�Bž�A���{�g��9&.?+�?I���w:�O>��-?)[�>��>��?�#�>����A�<���>`[6?)�L?!FK?:�>B�o<B���̜��=� ��:(.>��{>d��<�.>��ǽ����$ ���=�4>K��O�M���<���<�GG;��>يd>v�ο�3/�V�
�����վ<�)������*:��|:��\�}�r�y��|�>� ��x"��Y��bD��I4�jt��C�?��@�e>>+7�w�ȿ�l���	��L�=�Pվ�R��Ū��hka�2���{'���;?0�z.��?ӆ��s��7�'?���νǿ��:ܾ! ?�A ?`�y?���"���8�� >�?�<`4��[�뾂�����οg�����^?���>��5/�����>���>ãX>(Hq>���2鞾*/�<��?k�-?���>Q�r��ɿ!�����<���?�@�A?�i��UݾA�:=H��>˯?%�>B��+
��й���>��?@��?�g=��]�@J<i_?dUμ��E�w�;�a�=��\=~��3���6�M>n��>�	�ћe���ƽ�;>��i>���(�*�E�sώ= H>���s��3Մ?�z\�Mf���/��T��WV>��T?+�>�7�=��,?-7H�<}Ͽ��\�+a?�0�?���?��(?_ۿ��ך>[�ܾ+�M?�D6?K��>�d&���t�/��=::��y�����&V�*��=l��>|�>݁,���%�O�X����=L��[>ܿ`[���U$��P�>O�
�����!7����8�zv�=�����ͼD�=c>ž�¾V�>
?ݱG>�I>:?a�.?Aq>��>"��j}�ﳒ��_�=��Ծ>�.>��j>�
U��@���P���C��|�I����Zِ���R��|�H>��R��1����?�n���?�>�H?Kc�<2 ʾ$d<�7��<�k����¾���=u"��{���-���n�5�?�?�Ug��MV������=�`�K{?*���;�Ǿ��׾�d>�>�y��%�>�NF>�l��wþǒN�c&?��?�Yz�H���a�U8����<F�Q?��>;� >���> ��>\Ⱦ�5��	�f>���>���>&�>���=�&��%������>�_j?׶<�ൾ���>H�"��0��n�ʻF�o>��{��.��и�>^�=e��~��	]��V^�=��V?~3�>�2)��������nL*�]�7=�x?6D?��>��k?N�A?��<*���S��
��]�=ZlW?;ig?�h>X����ξs����5?��d?�I>{dk����7W1���i?2Fm?�?N���e|�1E�������4?6�v?�q^��r��\����V��<�>�[�>,��>��9�Fn�>-�>?�
#�MG��\����W4�|?�@��?�<<x���=;?{]�>��O��>ƾ�s��!���+�q=@$�>�����dv�h��FN,�m�8?2��?���>����1��?>b-��#��?쐘?H!��E>i�(�xo��"���־TP=Oˀ�1���u;Ѹf� �F����mWǾp����:�>�@t澣��>{量��忒�ֈ� wǾV����6?�,?��^��,���A�r�J����� m�f͡><i >�M��_ƙ��n}��g?�����_�>�0M���>��S�첾����!�i)�>N��>���>�wȽ�^¾�{�?˴���p˿���!��εW?�3�?[��??2?��<bz�n�i�y���=?��m?DlY?����]8�b��"�j?�_��tU`���4�wHE��U>�"3?C�>X�-�ײ|=�>���>g>�#/�r�Ŀ�ٶ�5���Y��?݉�?�o���>n��?{s+?�i�8���[����*�(�+��<A?�2>���H�!�80=�FҒ���
?V~0?J{�[.�b�_?��a�3�p���-�J�ƽ�ۡ>��0��e\�}R�����xXe���7Ay����?7^�?J�?\��� #�6%?��>d���M8Ǿ��<l��>�(�>�)N>I_���u>����:�+h	>���?�~�?Qj?���������T>��}?�Դ>�L�?4��=��>~f�=�4��&��%>
0�=�9�T\?�NF?��>��=��*-���E���T�[ ���A��q�>4�^?XL?D�q>�l����z��."�i���)�8�R�ʼb�G�6�3��᝽�f)>�#>!)>�QJ�&DԾ��?Kp�8�ؿj��*p'��54?)��>�?����t�'���;_?Oz�>�6��+���%���B�_��?�G�?>�?��׾�R̼�>=�>�I�>R�Խ����`�����7>1�B?M��D��t�o�s�>���?�@�ծ?hi��	?���P��ua~�A��7����=D�7?�0�X�z>���>�=�nv�ϻ���s����>�B�?{�?���>�l?��o�
�B���1=%M�>�k?�s?5o���ֲB>��?ޱ������K�^f?��
@Zu@��^?��*Ƨ�?B����#>KŊ=�P�=��X�]>à��ʼ���K�<MX >:�=�C�Ty�>�ؼ>��>ƊK>E���.+��>��ґ�����Rj��$�����Q���侜�<�l�-��%�W�]�5$��Z̺=����U�l5ѽ5��=�O?�D?|~f?�>�>2u�̤t=�B⾌5����3�b��=.Wr>�.?�\D?Y�!?!�*<iÕ�=
h��{�~/�������>��>>���>w��>�i�>���<��b>�g>� b>->��=}�z<u�2��8<>3�>+_�>>U�>�Q0>ʣB>�O���+��dm�Af���q޽1U�?`���L�YL���ɋ�ڎ���'�=�%2?,�=� ���ο�=���I?ڑ���$�J?F�c��=�(?[yK?�r>�����-׼�o�=���pQ���j=ӭ��رD�����,r>( ?Kw�>�L�>����0��+hW�<s���>�
?�����<^�Y��7��S��\O�>Y��>Ȃ��4P�(N���|�R���8�?�ȖY?�s$?-Ԕ��H�<����޾O�>n>�AT<���=�.�>�X3>�/�������꽶�Ľ�>�U?xh�>P�]=3��=B���7��1Q�>��>oe�=ayp?"S?`�K�zX5�H������>GG$?���>���=��h��B=Ⱦ>�7�>L�=�m��tQ�(�����?>�%¾�h2�:�B=��a=�Z|��l=�29��?"��{���΢��~?����㈿!��b���lD?+?���==�F<��"�) ��)J���?x�@�l�?��	�#�V���?�@�?7�����=J}�>k׫>�ξ�L��?��ŽxƢ�M�	��)#�TS�?k�?*�/��ʋ�	l��8>�^%?��Ӿ�h�>ki��Y�����G�u��h#=ߚ�>m@H?u[��K�O��>��w
?�?�d�������ȿZuv����>���?��?��m��<���@�c��>��?]Y?�xi>4q۾�]Z�ֈ�>�@?�R?��>�=�Az'���?9�?���?ϭI>j��?a�r?t��>�~���/�����9��0�|=������>�o>�׾�2ZC�����뚉�>i�D���^>�(=@�>I��j὾V�=T���������p��>�8w>ʞC>Z�>N�?<J�>}�>��C=voz����������K?��?�i���m���<r��=��^�Z�?*4?0IX�F�Ͼ���>��\?��?�~Z?��>N���:��^����H�����<�JL>���>���>�#��� L>~7Ծ�D�C�>���>(F���ھ�y���܌����>�$!?�R�>��=Uo ?��#?��l>��>ضD��摿��E��~�>��>4{?<+~?J?������2��sѡ��[�E�L>�x?3n?@��>n}�������h���B�6��t�?�g?|⽩�?��?�??�(A?�'d>&�VU־3��u�~>�+?::�<�#�E�6��Ӈ�E9?�:�>���>h�C��D�W�&=��徨V��2�>�+L?�?�#��b'��ž��=�k�<����'��`н�o�>@�X>������=��X>�s-��]ƾ����>7�M>�O >�z�;�O���cO�+,?�{&�i���}�=W�r���D���}> P>�B����^?� 9��h{�׺��e��Q�T�x�?'d�?��?����Ah��a<?��?V�?{V�>�+���޾;c⾉.w��~����w~>T�>�ZS����
 ��0L�������\Ž:`��F��>a �>c?{�?��>��>N
��G���r㾄��\�l�k��S��t�� ](��.��S���`;�@ʾ<���?�>�2�<I�>�?6xP>T�+>���>Ϗ�<��k>��=�v�>�P�>��>C͌=5[C>]٥<X) �gER?���0�'���辙���2B?��d?2/�>o�h�	���~���?�{�?�i�?�v>�nh�i,+� |?gn�>4��	m
?�:=���TՈ<!c��k������:��Բ�>b׽�:��M��Sf�i
?S+?@S����̾�4׽gڟ�&n=�c�?.�)?lw)���Q���o���W��{R��)��1e��ܠ��$��Do��򏿒Մ�p
��J(��*=�m*?!o�?���w���ͭ�!�k��,>��c>�R�>���>}��>�MN>��	��2���\��b&�_,��q�>�N{?���>,k9?�SG?|�s?��Z?=C>�$�>=��/?fM*>��>O{�>��4??�?��?��>��O?���>��)=�������>{�`?�MS?g��>R�?ֻ�e�¾�eỘ��:*���mɼF�
��>�a������46<���Dw?�d�z�6�dA��)�l>��5?���>W��>4S��$��7�7=�[�>�?䨃>�X���j������>���?�:��.=6�">|��=*ת�����=�f���5�=G�g�,�AE�:�ȹ=l)�=���ʎ�;|.@�TJ1�H`�<�x�>��?���>��>�T��ʦ ���(5�=��X>�NS>�%>�Aپ�y��|"��1�g�qey> s�?�w�?��f=�
�=Ջ�=uo���8��b�����`r�<��?�B#?J\T?���?O�=?hX#?��>�!��D���S��N��ڭ?N.?7L�>�Q۾�Ȼ��Ѥ�\�$����>vY�>K[�@�+�������-��tf�>F��m�E�����N�7����R��_�Q��?� �?��-<k!7�X^�����3���]@?�u?�gQ>���>{X	���Z�v�uS>a��>�=]?߸�>�DS?Ɓg?:?��s>����_��^X��óz>Q�{=|�?U�q?,�?��D?��>Zю>^Dֽ�����˾������@��i���;ƽg�d>�e{>ƻ?��>U�`=E��U�ؽ��s�"�)>�=d��>F�>Ow?�p>�~=bCA?3�>�����2����z
���۲�8��?�[?�*?��<=���_0���V��>�ے?�H�?'Y'?�&)��>�����ȕ��}��!ߠ>u�>��>3>�O��܌>���>��>�/����1��W)=%q�>I�b?|� >��ǿ��u����b疾��<������h�pҡ�2�J�U�=c^������֟�Zhe��ߨ�tT�����������r����>c�=^��=a�=���<�:����<]{c=��<�V�<�-
��B<L�Y�$�;������;��<=4k=����ƾV�z?9CF?��*?Z�=?��\>y >���:�>|6���?��U>s�(��̶��5=�?���;ڍ�,�ܾMiھ��[��b���'
>Q�c���>{{>>�6�=<��<�<�=�!o=��t=�Q���*=Y�=t��=��=/V�=�>yF>�6w?(���󲝿�4Q��[罫�:?�8�>.|�=�ƾf@?��>>~2������Tb��-?]��?�T�?*�?�ti��d�>����㎽Ur�=�����=2>���=��2�h��>y�J>}��K�������4�?��@$�??�ዿɢϿ`/>{��>��z>ܫ���A��}���s����P�[?gR���ǾlU=>T��>���<��.=��.>��m�=��B�6��=��н��=��};R4g>�Ϝ>�\��S������G��=�=�=ܗ8=
��y���%��
$>T�M���k>,
>���>?�0?t�V?"��>����M��;����?�;9�>9�^>�/�>q�b>�O�>��2?�-@?��D>���=&t�> ��>Q#�߶`�NF�%?e���G< d�?��?��}>�fؽ��Q�:�����}���?{�U?��?��4>{=�uX�u�C������^=7R��x�9<i6���ߙ=A���.ռ���Ӹ�=}Ɂ>c�E>	?�>>�>�ݑ>hz�>F<>ħu=d��~�=���=
 D�s�B�,�˽%o�<���<q��X���f=�h=>)pM==��=D>{�>�62>?��>��=����OY`>�$��j�@��"�=�%|�]�;�he�!�o����D��_0>�^>���m#�����>^�n>C�>��?�m?m�=YE_��n����f�1�޾g�n�=��=>���'K�
v\�R�;�
)˾��>�x>�?mz�>}��-��V&��	־�] �j�?������c9<,���:#���a��쌐��\�V�?�`���"�
�?3C?��?+�?c\������E>�a��uȔ�^�s��M5�ƴ�=*^	?���>�{�>��˾�.�̾��z�>w�I�\P�ƕ���0�&��x㷾�k�>����о5�2�hd��A؏�nkB���q�̺>qO?0�?ėb�A���fO�b���у�AG?�g?ß>�P?�?Y��}E�}���~�=!�n?���?TE�?��
>TO�<����d�=��?���?�ۘ?A�?w>d���>Ո�=�A�>ʪ=�]þ$Л�?�$����\>���?�f�?�2{�T��R�ž�ھ��_�1X���N^>���>�h�>�N>R��=�jy>Yd=��R=qu�>�y>,�<��}>�*�>	���œ�co.?�>8�>u4?#8y>��9=�$���(�<��h��n��v"�®A�_�%	<q2�	c =�.���>��ſ��?rd>���Y}?}�龭�X�;�c>w�*>b!�
��>��5>;n>-L�>�>�4>��>��>>�Ҿ"�>�����!��eC�s�R�m�Ѿeg{>mS��'�7r�OD���I�ZO������i�����X=��C�<�6�?�����k�+�)����x�?���>`�6?r)��������>���>���>q���I9��+n�����0�?���?�;c>��>0�W?�?�1��3�vZ��u�W(A�e�4�`�o፿윁�ݗ
������_?��x?�xA?:O�<@:z>;��?��%�xӏ��)�>�/�';�wB<=�+�>�)��W�`�Z�Ӿ?�þj8��HF>��o?3%�?uY?TV��1��e>7F?��y?��?���>�K?pξn�*?�>s�X>#<0?6p?1
�>��	?)�>ۅ�=t'�=�>��K�^^=�;: �8H7��V�=`�=�؀=ᮆ>M�>��k�һ�F��Ӗb����������:40ݽ��@=ނ>>E&]?�j�>�4�>j_1?x �Y	$�;@Ⱦ8�Q?v�>h��*�D�M�����ɾL+���0j?���?�P?4Ə>6�I��I7�'iM>��>I>��">���>���9~y��|>���=1�=�]���DN�{����D���K �H�>ȿN>��>�7>�/�=�D>�(���]&��G>�L��%��6�B�e>��W�L�Z����>\�D?��	?��V�4i��{<ǽ�ia�vW?�B?=5N?�܈?8>3(��X�5��m<�Yǉ�3�w>�<#���͙�IU���7�)�=���>.l��D=��j�>G����߶�<=m�`u��F��NV>43��L>B�˾?�$���̾��>2.�>[�+�߾�*����板��J?�-�=��r��h����ʒ>��>?�?�U彇�>�8�Ӕ�|@���	?���>��B>��4���H� �p�'`�>x�/?��I?��?6�W�q�V�^[?���~
��/��t?I-�>�	?a�=�0h=�qs����$O��$����>�V?X�1��(i���¾F����u�E�>�7Q>�,7>���>��I?19?�?�
?�(?]<)>��'��-����?�]l?M��<�������}1�<0A�:�?mל>/VZ���>mg�>V�;?�
{>�?�[2?�?�=���:�Ƶ>݁X>�LF�n��t@�=�mG?0�_>|�]?��U?q�>�l%�fÆ�V<ʽi��=y�<��$?ȱ??�v?#��>_P�>��*��=�q	?�qn?�8p?tv�?��̻;\?��>��>)<�<�">�l>?��D?�i?u�I?�9?�B =>�)�����ٽn�Y���߼��=�;C>3�m^W�2"�P�7=����g�f���^8������|F=@Wp;��>˶~>NS���zD>p弾�0o�X(C>�"�����tQ��1����_�<4�`>4 ?~Ŗ>�;���m=��>��>�d��r?Z}�>?�(?�Q�=Y�O��B���Lz����>�,5?:����l�1����[{�Jr�<��f?SO^?2;��%�վS=c?T?]? ��;:�F þ�^��a�9>N?e
?��N��X�>�}?R�r?~7�> �f���i��v���$a�.<g��}�=n��>�4�аg���>�7?���>�Ng>tz�=ʮ׾kVv�
����?}ߋ?׭?,��?_ &>6�n��߿��澈���io?;v�>u�g�_^.?H'��꼾�𖾝'����Ծ�,ݾ���E�d������=�݁���d���\�=?�6[?��u?пd?��о.Z�PMJ����a�=�a����J��nF�O|C�j�2�A�p��Y�J��

�����=�(>���I�$2�?��9?fǼ��?����\�����ڮ=2(��jj��z�p=�.<-�;(�׻wv��V�5�������?���>nD�>�Q>?�VN�x@��{.���H��"����#>K0�>��>��>�=B�P���o��P¾�+���&��c>+[?�H?�h?��ʽ%�/�=삿�q������������>��>�e{>9�L�:�����<�B��/s�����㕾�� {>';7?� �>wX�>��?�i?{����OǾg�i�jp;�+E=̕�>__?�U�>�d�>i���8$��n�>9ll?�w�>k��>U/��/!��{��zȽ�_�>�C�>���>�n>��+�c\�E��$���_8�%��=��g?C����`�%�>O�Q?bE;I�L<:��>T6��x"�Y4���&�*
>�"?�C�=	�;>wƾo��O|��U���)?��?]���/�*���y>!?´�>��>�҂?!�>�¾�w�;Q?l�[?�:H?�!A?z�>U�=ꮽOzŽ�	'�ċ%=N>�EZ>ܞt=]i�=&���[�����I=LF�=
 ޼�ӵ�cj�;�Ҷ���<��=N�2>�տ7��[��A��:
���0��Y��K���I��,�Soվ��}��[�����O�����)�w���̽=,\�D��?Z�@ll=�CV�(u��h޴�ײ7�Q�n<��ž�vX=��@�����h޾��پ5<�N���Fa��z��Џ�|�'?G�����ǿð��6;ܾ�  ?�@ ?��y?��;�"���8��� >�;�<='����3���=�ο����I�^?���>*�-+����>���>3�X>mGq>+��"鞾X7�<
�?��-?���> �r�!�ɿ􊻿_Ϥ<g��?:�@�lC?�L"�ި���J=�A�>-�?��.>�U#��/!�������>1p�?�)�?��b=��V�TWC�bT^?W��;snE���޻��=��=e�</��n�H>~�>^����c�V4��<N>���>��k��򽷝P��[�lc>S���x��5Մ?+{\��f���/��T��U>��T? +�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?$�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�݅�=�6�����{���&V�}��=[��>a�>,������O��I��P��=`��Uf�.���M�_T�=y�N>�6j>yz>�
? �5���x��Ȉ>㛻>w!?�I6��b�G�\? �?a�?:�*?2�:?C��>���=v�׽���T0x���>ٍ&�D0>0�<��^��-���������p��LоlŎ�Ҙ�H:����=�3D�'|��,.�  z��~Q���$?c~>d�ƾ�@�[���%ξ?���Ἷܲ���;�1��u��ߟ?�*O?d����Q��,�7��:.���1R?�os��澑ޑ�i�>�c���"=Z�>-/�=
̾�b6�R>[�§?��?M���iؾ|-˽�׼U��Qo?�9O>�G�>I�>��>���]ƾ��;o�>��>Ɲ-?��>���Ľ��?�*?��r<G�^��z�>3�����ɾt_��,L�>9. ���
�f`h>��>�z�hܽ��7��:½��V?͍>۷)���1���tg��;=�x?E�?�O�>�%k?R�B?Gߛ<f����S�:�
�|{=��W?�h?�H>5�J�Ͼ{+����5?Eme?>O>��h���:�.�
�	�?Q2n???����}����R���6?��v?�k^�9p�������V��9�>�U�>W��>R�9�z{�>q�>?�#�G��\���V4��?%�@y��?�<<p(�*��=:?�_�>�O��@ƾ�������U�q="�>���Qcv�T��wU,�ׄ8?۞�?���>N���y��B�>�;R�?�`�?!�T����=��c��O6���Լ��=��������2i��e���*�:�财������O>��@N�ɾ���>E����׿n���֝��,Ov�{;;?��9?PU��oƺ������f��l��9!��XB�&_�>��>j����Đ�Nv{��<��1��Y�>��*��_�>�TP�\+���֛�TY@;+��>���>�U�>ο�������?F�����̿#Ҟ�CK���W?�ʝ?�p�?=�?,
�<Rix�.w��H+�*sE?7�q?eUX?��,���V�i���j?k_��`U`���4�_HE��U>�"3?�B�>A�-�-�|=�>{��>�f>�#/�p�Ŀsٶ����Z��?؉�?�o����>n��?ls+?�i�8��e[����*���+��<A?�2>���;�!�@0=�$Ғ�¼
?1~0?�z�Z.�Z�_?�a�@�p���-���ƽ�ۡ>�0��e\�:O������Xe����@y����?J^�?c�?$��� #�P6%?�>k����8Ǿ��<���>�(�>�)N> H_���u>����:��h	>���?�~�?Nj?򕏿�����U>��}?89�>�Y�?,��=�1�>��>����K<�ak>˖�=Q�ƻ[�?G�S?���>VO�=7�.�%L$���N�DjU�d�����B�Yn>Vk?��R?.D�>�唽4�(�:+�����L�b�I=�L��>ܼŶɽBF>`k)>�&.>Y�$�� þ#�>�5�H�ۿ1���o�`�2?�O�>��?u�վϤ�o����*b?G�>������易��6���?7W�?�H?�ɾj��! >m�>2�e>[\�I�A��ג��#R>B�>?���Hu��<s�ے>��?W�@�0�?J�^��	?���P��Wa~����7�]��=��7?�0�B�z>���>��=�nv�ݻ��T�s�ù�>�B�?�{�?��>�l?��o�G�B���1=*M�>ɜk?�s?JRo���v�B>��?������L��f?�
@zu@_�^?$[��M{�����(�Ⱦ���=|�>{��>����>OE����&t8> �>�V�>h�P=��<\��>i,R> O�>����I'���ʿ���T�D�<�۾l�
�5�q��@!���&Q�u�,�����|�>�H�)�׾�H��1��Q[<(��=�FU?��Q?%�o?�� ?r�i�ez#>H�����<��"�$Ў=��>s�3?z+L?Q~*?��=�����"b����`���*���&Y�>#�C>ђ�>]��>?'�>�;�;�*I>�3=>Rdz>�0>LI"=���:!�=m'M>c.�>��>�F�>"�6>0�*>�����,����k���gT����?蔾];��䖿l4���qžx�=�5?@�>����ѿ��?5F?�Б�����9��]>�z1?*�M?�*>]֧�T]��g>nK��Nc����=���[T�H9"�xMG>�\?ڽ�>'��>�:��s>���b�և˾8"���3?kE��b�N>����vU�-<�l�P>O�6?O�=r�W��թ��(p���!���޼O(?�l�>��0�j*��CeI��>þ��d=Y��=I�p>k��>R�
>����1�bu1�/�3>7%>�i�>9J?㨇>6�=Y�~=��˾+��K>�<�>F�=JA?J�?����j���־GA��T�>U�>R��>�a�=�)R���;
�>���>���<�ݽ����<��e�>"��||�U&J�HfG=����y4)>��^�􄸽�fK�e,P��~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾOh�>{x��Z�������u�v�#=R��>�8H?�V����O�g>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾;`Z����>һ@?�R?�>�9��'���?�޶?֯�?��H>j-�?�hs?`S�>��r���.��س�7�����=;�;�Y�>J�>c׿��E�M����u�i������_>S�%=��>��� 
��@!�=W���X��H�q�a�>�Zo>�G>ҝ>�?���>��>��+=��.%������WL?ڎ?2��m����<[�=@�c�� ?W02?���veѾ�%�>� \?�?��[?�5�>��V��pq��dĳ��J�<t�M>��>A2�>*<���FE>ьվTEG��}�>�k�>s�>��Jݾ�3���j)�˚>*j ?���>��=b�!?I# ?�Bu>K�>�J:��6��(�4�P��>,�>2��>��}?��?#���2.��㋿+}��]`U�tV>�w?ZY&?�O�>j[��d������`	��6F�@Y�?�Y?�$�T�?@��?�`I?BY@?�}I>��ҽ?%�&���>`+?-�O��3-��q4��.���?��>�h�>�G�D������"��\Ǿ��?SGc?�-?9(��k�X��|��=��h�`���Y�<�k�v�8>P�:��)�Y�%>�</>r��^n��^����2����R>�8i>������Z���R�(?P�;߁�N�=ls���C�_>��]>=.���_?Y%��uy�ɢ��
���$�_��3�?5��?a%�?Gį��jf���7?h�?+�?H��>�p����־��,������5���>K�>�\:<�)׾֤��㤿s&���ʽ5}�����>P��>�N:?�R'?�>Y>@��>nԒ���'��8�־��I���辮�=�Xw+�����7� �M��l�#�ھ2j����>�ռ���>�?Y�W>�^~>}�>*�#�=<�>͙�>&/�>�$�>˺=�w����z���LR?�����'����䪰��/B?�kd?2�>�\j��������v?��?�o�?�Lv>"zh�r(+��t?+�>Y���b
?�:=:��|��<�D��1���P��������>��׽k$:�,M���f�Z]
?�&?
��i�̾��ֽb����o=�K�?�(?��)���Q�m�o���W��S�?��+h��m��c�$���p��珿uZ���#����(�/�)=��*?c�?C����])��m!k��?�d.f>E��>�,�>�޾>;�I>��	�V�1���]��B'������R�>S{?4`�>&C8?�3B?O
o?1FW?`�>@7�>���"�>�X>�]�>�� ?L�[?��?�.?(�?A�%?��b>�e��������X?��G?��?�ޓ>Y�?Ǧ�<���=g=���=	�侩��8k���>�!]�<�/L=9v/>m�?�)1�w�9��v ���>\A?�U?bܼ>u�b��1_�)�=�>�>'��>bv>~y��7c�
����a�>?֋?�
��k=��+>���=��=<����*��=��)9�h�=*'޻�Z�59����=iǠ=���;z{�;���5� <��1<���>�#?�֑>c�>[KX��%��0�����=�1u>�S8>�r>��ʾ����q���f[�=�>� �?2�?/v=U�>)-�=���������S�����m�
?4 ?+�4?�#�?Ek>?��#?�2>K��~폿2����0��j�?�X4?�̆>���&�ξ;y��t?)����>��>��c�nUV<����M�~�.���!>��.tO��]��.�[�%.y<���c��?��?Re�?`>x�@�:�Ծ>��^�����-?`�7?wO�>���>9��s��_��>�)�>~�z?BB�>��F?F�~?ʿi?�ĸ>aaɾ��y�D�̿�s��h�>ܓ;?�?���?8�\?H�>%%~=�g������5o�Q���^��Ǿ|���>�*�>h�>?��>��q�%H+���ƽBޠ=Jg:>q�x>?��>���>��>>��>��7�d"8?��>;1����"�/��$���#8���?l�w?�:?���9 :���4����Mۍ>Hޞ?��?_1'?ݥ%��m�=1Uk������#��R#�>$�?�7�>�I��,>gu9>��>?0�>��Ⱦq�*��x�@K?�I?6`�>�Ŀ�jp��u�j��hC�<UO��i	r��g�w�>���=��3J������Y��ꣾ�����T��l���'Uy����>��=��=�L�=D��<r�׼�:<�uk=k��<]=��f����;=+�� %�k������;��;�=)=v�l�d��5�s?@?@�#?��.?�}7>s��=50���]>��۽s3?��K>����	�������ї�i܈��پr�;*:V�X���]T
>o�m���>�`7>}��=߻1�5��=Eו;tb=�y�:�s:=��=M�Y=2�=.��=��=��X=�6w?W�������4Q��Z罤�:?�8�>i{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?=ti��d�>L���㎽�q�=N����=2>t��=x�2�S��>��J>���K��I����4�?��@��??�ዿϢϿ7a/>4Ts>�w�>��J�-�d@��8���G��2?s/��������>5�>����o��v�<�;�>���>�(Z�;�>�GH�=C	���Wu�����5�>J�>e�M=񝢼5k>�@�=3? �o|�=)��<f`;E.X�3na=7I>:�T>w�=�y�>`�?��-?"�f?'�>��a�)���>���3�>m�=n�>�e�=�}N>8�>�D2?��B?pB?h��>�c�=Gj�>Ht�>+ -���p�QU�F!���n���?�Ѐ?���>Y'<��A� ��9�7��?׽�?�E&?`��>BԔ>!W�ڼ��	'��.����z8�:4�0=��n�M�D-�?M���߽$;�=���>��>T�>�|z>�9>�R>	B�>+m>�}�<�G�=`$�!$�<�������=�K�G��<���tV���q^�2�5��1�����;�dI;�0<٬;"�;>�]�>�.>@��>��>D"��P�;>j���<�)��<�2=�qG��YT�1�m�p�u/�2�h>q�D>�!�:����p�>�l�>�4�>�q�?��i?Mg�>�_��t�������žH�p�3�=��.�ۺq�I-�J�+�I�_�+Mx�"J�>qcw>i]�>薃>ڂ
��#+������ؾ-i9�g��>�������f�#���P�Ւ����� �u�4&s���:?����L˽�_�?�Z?";�?�k?�~�L����c>+�;eϬ��.<�����G�S�?�'?xL�>KYվ��Q���˾���ɕ�>ʋI�~P���۸0�m�	���� ��>Kު���о��2��m��0돿$8B�U�q���>�aO?�ܮ?�Nb�DB��}O���������m?-pg?Ѥ�>�j?? C�����a0���=�n?��?H7�?�>���=. ����>�y?�7�?O��?_ٯ?����e��>�ڨ=��>�Bս�>��D�>}�>�h�=��>�?E�~?�qu�7�վ���0�SW��hB��䬽/˨>t<�>���>��_>7��<���=b�>_�s=���>��>�#?��>ЩQ�׶�öI?�O>�8�>.�5?���=��=��:��X���x=�{��]�ƽ��<(��E>T=>5Z�y���GP��>�ԿK�?-Ί>;���ntO?����?=�S>��˼.۰��<7�H>� �>�
u>��>	�>h!w>�n=#=Ӿ:�>���MZ!��+C�׊R���ѾB�z>���+#&�Ԗ����gI��~��2c�d�i�T-���@=�H*�<�E�?�t��!�k���)����=�?mo�>�6?K��D���j�>d��>Lݍ>�V�����������jᾊ�?���?�1c>�>o�W?��?|�1��*3��uZ�ӥu��"A��e�2�`� ߍ�R���ݗ
������_?�x?oA?Ė�<�4z>ڞ�?��%��Џ�*�>P/��';��t<=�8�>�)����`�1�Ӿl�þW8��?F>�o?y!�?*N?0WV���=3��>�W3?��1?��k?)�)?+�E?�3��:?&�\>�w�>:�Y?��[?�E?��?��>R"�=,�=�`��J�-��S�53��(��E�kA<Cn9���Y>�C!>h�=�8άq��U��JSu<#����>s�s>`��;�`t>��>�-Y?�6�>@nh>�/?�D���1�eK����*?�@{=!Cr��m��ݟ�����G��=z�g?�f�?[�Y?��[>�/A���C�j�>I��>%�<>�JQ>���>o�2hT�Q7Y=�=>q�>wt�=i�����m�?v��y�O;s�>���>mԠ>�����)>�����ҾW�=�.��-)᾵��QS%��1"�a���X�D>
XT?��?㩶=�$��C.��W���	?,$?�h?}?���ZɅ�-�H�jQ���ȾT��>gc&>���Ϙ�������2�>���>2�޾M;����X>xS�����Y���_�7F��S��<�%��[3<$b��9ľޭؽ��>���>[C��6�6��Փ�����dB?���sǾaΛ����i@
>��Z>ww�>j*���=�u�������=���>p>�>[���1��*�J��_��>��?�pi?���?���4L�������|��z�n��;?�Q?�?��>F�~��$�=�j�M�:/=�J��>�?ȧ=�j=M�rP���ܾv$$��ۇ>��>�cu>á?�'8?� ?��X?�^�>�|,?���>�����c����?��u?z��R1m��՜�g0�9BO�#�?�.?�����	>��?-�	?��?��?x�
?�}>
\���."�ɽ�>妇>[H�P���o�=�WB?ѓ[>��?ͨ�?��E>������ü\�'ڽA>h�??=3?��1?x��>c �>:䇾9
�=n
�>ƭ`?U�m?2f?�#�=��?�dD>>�>�;�=�U�>��>�?˰N?��m?rhW?���>�_<T-�����גJ��A��¥2<��<D]�=bFU�-��񤼼���<[��<1X'��v�;5D4������O�Ni�\�>�-t>���o�0>��ľ�9��#B@>>'�����͊�D:�uø=���>`�?JΕ>��"�f��=˶�>�@�>v���(?j�?��?�;��b�m�ھx�J���>��A?�P�=X�l�do���u���e=n�m?_^?9zV����X_?�R?�m�:�C2;�<�;,@̾zI9?�5�>��g���>��d?�/r?r�>��!��^Q��+��w}`��%���y> �>ŀ ���x����>��K?|�u>��>X@�=&𜾺^���Я�?p �?�ٵ?�?6b==PO`�\+տd��s]���M\?G��>�<���!"?�aػ��оʏ���ތ����˩�뒯��̗��-��0/'��j���R׽P�=T�?W�t?�q?j�_?}� �Vd���]����^�V��'�����^E�$E�n�C��/n��7��*���2����*=Ϩ\��DN���?��B?�c<�/?	a�����ܷ�N��=S�a��o�p3�<�����Kf'��LѾ�=b���c�?0?J��>8��>��)?��e���7��p�:��
�^=��>�A�>���>e�;�B�R���b�e苾�=���w>TLc?�K?dxn?�P ���0�P��I[!�T�2�j;����C>s�>�>\yW�E���)&��9>�1�r�$��u~��d�	��= �2?!�>pg�>Y�?,�?�	�n%��M�x��m1��	G<w��>toh?�V�>݇�>��н� ���> �l?Θ�>7��>d���2]!���{��gʽ��>@խ>��>�=p>9�,��\��U���y����8���=&�h?�~��e�`�Eυ>�R?��:uQJ<~�>�,x�m�!����p'��>�o?���=�_;>��ž�6�B�{�R���w&?��?ר��۟)���r>��?�_�>��>wY{?��>c����+=]H?{�9?T�K?B�D? ��>���=$i��=ө�����=��>G>��Y=�=�c�9�V���
���|=�R�=rz��$����qN=�����Ԣ�T��=��!>�Wܿ�P�Ì�@�����|l��C���Dk��u+�F��<{ ���l;�B��Fl̾X)���j��0�������>�њ�?G�@��<��x��z���������f>�+ؾl���{�뾙B���3�q鼾�L$��V��?:�҂���t����'?ʻ����ǿ�����@ܾw! ?)F ?��y?I�	�"��8�)� >Zo�<`|��-��ɚ����ο������^?���>�	�,��3�>���>͒X>jQq>���m瞾Q�<P�?D�-?=��>r�!�ɿk���HҤ<R��?��@��=?�j׾�!־�C�=��>�U?.1>�q�������Sy?���?E��?��:�}F��8��>>?��˽y}V��� >�d>ͺ���i<�b���>��=8���yN�H<���m�>�/=?t=��Ỻ�7�{��>l/��3��%�C�5Մ?,{\��f���/��T��U>��T?�*�>R:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?$�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=6�뉤�z���&V�}��=Z��>c�>,������O��I��T��=�����'�G��J�Ȓ��G�����;��I��b<>?��>��f�����%<���E �,��������n>>�z�>@@H?��\?(ڔ>��=>�-���z��ƾ���K��;ƽ������=��݁<{޾���`�&@оK��<���ƾ�<��c>��U�*����R��C���zK�4<�>�E�=��辘qX���>�O���:��
��`�����X����r�?�	s?	x�
b}�a"��P�=w-*��߈?Șx���A�r������=�7>;��>)��>d<�>׌.�d J��_Y�9;?I?bM��rNӾ���\F�6�f�@�\?�?h}L>^ O=X^�>�s��A�M��>��?�ɭ>*H?$��>*�� _&��h?5&?8�u
���I�>4��co��nn�pN�=�W ;��ӾFz�>��ؽ��˾�\�=����46���V?�͍>�E)�����k��W �V?=�Hx?�Q?�-�>�Lj?O"C?�ơ<����fR�!
����=�)W?��h?��>���9�Ͼ;����5?r@e?{�P>��k������.�8W�.J?�gm?��?����"*}�j����H��k5?��v?�r^�bs�����d�V�'=�>�[�>H��>��9��k�>�>?�#��G������AY4�)Þ?s�@���?P�;<> ����=�;?L\�>@�O��>ƾ{��˃����q=�"�>񌧾lev����~R,�9�8?Ҡ�?:��>������ .�=��پ2��?`-�?rF�	0�=i뾥Fy���炾��Z>=2���&���+E���f*���ӾQ�����>�@m*L�qx�>�Ⱦ��N�����iC��ܳ��� ?��&?���=��R��H��f��sȾ�g�e����@�>��">���VǍ���{��� ��M=6Ī>��w��	>�uƽFv���<��E�`=z>���>^\>t&������?�Ծ�ſE����T߾�F�?u�t?���?�f&?fv=� ��]�����>a_-?��z?��Y?�ѯ���d��U��%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�_�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.��_?�a�s�p��-��	ǽ�_�>�0��A\��4��a���Ye�z���w�x�#�?�W�?d�?+�'#�� %?���>럕��VǾ�I�<(��>F�>��M>{�]��)u>7��$;�P_	>���?�q�?�?��������P�>��}?� �>�?X�=�V�>�^�=��jp.�uk#>��=oE?��?Z�M?tA�>�^�=	�8�/��RF��CR�/��C�N
�>��a?�}L?�Ib>����1��!���ͽx�1����{P@��,��e߽�	5>f�=>G�>��D��
Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�_��=��7?�0��z>���>��=�nv�޻��W�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?Qo���i�B>��?"������L��f?�
@u@a�^?*�����Z����;���=���=�H>��뽑q>8�t>�	���q�	�<���>N͔>�:>*��>I�o>�%~>u2��H�$�bj��O=����8�����j
����!*���>�
��4wľ<���A2�� ���ȽoF<�%>����=�U? �Q?��o?u ?<�z���>�E��mp=��#�[7�=���>�G2?#�L?v�*?��=�e����d��?��
��/���y]�>�I>�:�>J�>��>u�":نI>�K>>��>x� >N�(=�s����=WO>�>
��>�U�>9�>��
>*?��iѮ��P_�zZ��Q���ؕ?g7̾˶2��Ѧ�釾	����B>��L?��=�{����Ͽcµ�DD?���o�
��˵��������>7�j?�(Y=)⾾^�<W��=rRѽf:d��^>hj��$w����!���=��?�!�>�
Z>*A1�t52��R`�5՜�S:�>=V%?AXϾ,���8u�rD��BɾM�>���>ok���0!��@��������d����=%1?��?C����RǾG>f�O	��Ah=>�h>>S��=�Д=�q>س��	.��M�׈�<&P>2jy>ؕ ?%�9>9�>=�sf>k���)j�99�>���>��N>�N2?p�?`輲Ŵ�v��tӽ�ɯ>�h�>ܩ�>q�I>\�>��u�=���>�P>���|�S�L����ŢN>@�����;�ݡ��=S=��߽;�=��=�� �~�]���b�rb?�Ŧ�
��DP��ڽ6D?��?$5�=�'v�7���ۦ�oܹ����?.A@m�?�t�8W��?SO�?3������=�]�>�8�>�0о9�X�	?(�̽���ʡ	�a��#t�? ��?��Y����k�U.>8%?�,;Qh�>ux��Z�������u���#=P��>�8H?�V����O�`>��v
?�?�^�ߩ����ȿ0|v����>S�?���?c�m��A���@����>;��?�gY?toi>�g۾B`Z����>л@?�R?�>�9�p�'���?�޶?ӯ�?�
I>x��?ɘs?(n�>�"x��\/��0��:����~=ݺQ;pu�>!�>9����UF�-ғ�~e���j������a>��$=��>�e�.��K�=9��_@���\f����>N-q>��I>�T�> � ?|a�>h��>L�=wc��LԀ�����]GL?���?�_��m�-�<e¤=!�`�M�?(u3?����;�:�>E�]?�%�?`[?�$�>�/����Z˿��?���l�<�(L>�m�>�I�>�����L>��Ӿ�BE���>�
�>�<��uݾ�e��ᾯ�%��>�!?1��>�2�=� ?��#?��j>1A�>�FE�� ��5�E����>���>�(?��~?=?]e��#_3�H��~䡿�m[�75N>��x?7i?�ٕ>G���K���D�I��>G��[�����?�Zg?���/&?'�?�??�A?}[e>���f�׾M���ŀ>��+?�{��XJ�p���U��e�?q��>���>9w��CS>�e��=*�
��!w��:�>��[?�'?�X�
�Y��\�1=�.�'f��4҈<�
=9�>�>I� �N>�<�=EU�=mb���Y������5>�c(>M쟻KJ�\U@��",?�A�/����͗=�r�D��~>p�L>X��0�^?#�=�ܺ{�����q���pT����?��?�W�?����h���<?��??k�>9I���e޾���w��y��w�[>O��>��`����P����\��
h���{Ž�#K��C>��=?W%_?8�4?A/?*8?P�ԾO);�m�u�M�= ��Y�4��j�e�[�֦M��j��q����=�i�4u��c�>E.�=���>�X�>-I�>�-e=(�>��S>�ޘ=��>z�>eH>�=���>�>!�*<�=T=P�R?�v��*�'��%�v��N�B?Ϭe?[<�>�j��񏄿���?B�?E �?)}>0�h��1,��8?~5�>��~�Ï	?s�<=Qj��N��<���_t�3����3�>��ν��8��QM�Y�a��-?Sp?�z���1˾��ѽ�����n=�O�?~)?U�)���Q� �o���W�S�\P��h�$P����$�<�p�?쏿/`���#��Ϡ(��4*=�*?��?я����L*���(k��?�}Pf>��>�&�>�>�I>��	�ʹ1���]�E'�K����N�>S{?�>%;=?/�H?�
T?�e?�>�P�>���5��>�ȝ=u@>ч�>VP6?�w?�#?�%&?f�9?8Q�>t+�<Щ��ƾk$�>�0?���>�A?C4�>h�l�_�뽎7��13<�[V������Ƽ��>[�ð��8=��>5c?f!���f8����~Cl>��+?���>�G�>���}#��4�����>� ?\<>�����yV�?���k��>��?����\=�� >\�=�v��G&<]V�=�7����>�]C���V�+�j=�2">��<�1o=�e=�[��� �=h�=Xq�>�?���>�!�>�>��ڪ �,��z.�=�?Y>zS>�>�Oپut���"��g�g���y>eq�?�y�?�g=W�=a�=�r���H����彾�T�<�?B6#?�OT?X��?a�=?~Y#?��>C ��A���X�������?�M?կ�=C�ξ.�O��r��2>����p?��S>����`�Խ]��) ��M�G+/?�i��쏿ee��^�m��ھ��������?�$�?==�H��߸�"mo�9�о��?��A?в>Y�f>��Ӿ�E��9���k�=�1�>rE?bٷ>5.H?��}?��b?��r>$�9�y��d�����;���=��E?}3�?���?�}?�²>Ѥ>j-�� پD��z�������Rm�:;�x>�Ń>�\�>���>9�>w���0����[�mh�=6XI>��> �>&@�>+ϖ>l�G=��6?R�>�)�����:D���)��G,d�ze�?��?��?"��'$����k��\�>A\�?�2�?�;A?�1�&�>�鑽�|���炾њ�>g�>"�>��(>󒼼866>/�>A{�>��=�S���� ���=��>:�F?�� >�pҿ���^?��H��������y�`��딽�-�eb>Wf���-���ɾ
�n�[�¾����Ū�F,��ź?�� ?^"&=T�=�s">��
=�hH�u�<�[�=m��<��=�W�<߯�=��׼ъ�<`�A����;,�����<a�*=��ž��x?�E?L&?-@?g�^>CC�=I꼯��>�Q���1?��v>�:<�k����F.�[��=�����Ծ��;��X������>�sl�ܟ>B�4>أ�=Ӓ=;"�=�Z'=oo�=+�qlC=	��=��=���=۰�=��>�F>�6w?X�������4Q��Z罦�:?�8�>d{�=��ƾp@?�>>�2������xb��-?���?�T�?=�?Ati��d�>M���㎽�q�=F����=2>l��=s�2�T��>��J>���K��>����4�?��@��??�ዿТϿ4a/>��=z�
?�e`�"�_�{�¢;U��r�2?�ǚ��䨾?�&>
D��N��Ȣ��b6�̌�>��>	���`���=M.�ag=K�;���>k6>Q`=��=rRĽO�>��<��=N��\r<�_��=��X�޼��>}��>B��>�?�B8?��_?���>���G���8�;7s>���<��>56q>E��>�>�>���>�a/?�'?�)�>m��=���>܌�>�8&�_��A#f��@�h����gh?Ή�?���>)B��q˹�H����mM������?�LT?�bC?*�|>������4��$�����Eܽ��<�HU���=��V>�ɝ��H�4�T�EDl>͐7>.�>��>��l>���>р�>�!�=����=w�佋ʔ��.0=U� =_�H�U*>Rު=�Ʉ=�n�=�q��о� �ӻk���3=�a>^��=ZN�>�s>�T�>uτ=���)d@>�h���`L��/�=>j����9�^)c���x��L+���9�^�I>�BP>S0���c��:��>\�N>�F>� �?��t?]�(>�L$�e���u��_L��T��R�=_L>��J�l�:��d��P�L�پ�|�>T~�<c?�N�>˹��$�V���N ��P����>�= ���L�d��e޾�L��iF��T薿��D�g�?����l4����?�U�?b�?]�7?��!����O;?��þ�nW=�'G�Hξ��_�@��>�& ?��v>~�־�A.�.H̾����޷>AI���O���u�0���^̷����>����i�о$3��g��������B��Kr�V��>	�O?o�?�9b��W��GUO�����'��tq?}g?c�>�J?�@?�(���y�s���v�=�n?���?D=�?�>�1�=s����D?+[?�۠?�r?�6�?�r���s�>��g=q�@>]�M�	_+>{>��<�|��G9?��??%���Ѿ�߾1"��7 �� ��=�T�;C�>E��>}A>U,Z�I�'>`#>]>J>�N�>r�>U�>i]�>��>�ܢ�,C�"�&?Oy�=�^�>Ĥ3?�u�>6�/=����h<6��]?���0�煥�V�彯��<��L��&-=|&��k�>�zſ�8�?�7F>K���	?����A��i[>۶U>�e�5�>�
O>��r>���>��>�w>^K�>A">nFӾ�>����d!��,C�@�R�v�Ѿ�}z>˜���	&�����w��\BI�Kn��Dg�rj�9.��M<=��Ƚ<H�?������k��)�6���O�?�[�>�6?rڌ�]����>~��>�Ǎ>�J��R���Dȍ��gᾗ�?��?�;c>(�>��W?��?��1�>3�qtZ���u�x%A��e���`�O���������
����G�_?��x?�yA?w�<k8z>���?��%��֏�M*�>a/�&&;�7<=�,�>M&����`���Ӿ�þi>��NF>��o?)%�?�Z?gNV��Z$�a�7>b;? �1?kt?���>�h!?��O�̹?�C�=�d�>.�?��;?u.?U�	?�h>�ۻ=J��=M��=mp���kw��#���5�{B�U.[=�=��>�\�<.jd��o���=�.�="�½M�9�^�(=q�ۼ���=��<Mu�>OTA?�P?RA�>�<8?����=^��{���N#?�v\>:����)��_$%�"E��6,!>�nq?o�?�K\?Y�>?2X��Vz��!>e��>R�=,�2>_��>����o�ϽG�>�H>0�ʼ[�ؼ�i�38+��?��%�!��x�={1?lu>�]��/�@>�@��QE����>\}?���Ӿ����h�<�9�0��꛾ky�>��C?��?�:�<���5���e���?3M?��Q?�gw?��*=�軾��4�v�Q�g �-~�>ؖ�����嘿�>��̴=�И^�lQ�>�J��l����>n���(_��U����T�2��>��־ٰ	=��|�}W"��ѫ�WG�="�=LY�հؾ�o��(��`cc?x^t<&��R���R\���u>C�:>g�n>bC�����C_��)���Ɲ�߻�>+�i>bO/=gW�E2����P�>��A?��f?�Ë?+��l�r���C����NI��<�I��r?Ԭ>�?�;^>���=*A�����b/^���@�K��>��>S�(�dP�*b����־S"�>^�>��>x8�=$~?ԎS?Fp?��R?�:0?���>E4>�K��Sɾ��)?�Ƅ?�&,=�=���<+�DS���>��7?@�J�R6�>��?�e?	�
?1�h?�(?�1>����97�z��>s�>�d�ED���{>�M?� �>�wI?g~?�Bc>&C�B���A��k)C��Y>��2?.�?�7?���>���>�Z��\="�>��b?x�?�o?zF�=�?�q1>ױ�>��=�N�>.��>��?�SO?x�s?[�J?��>�1�<񺭽q����9r��CT��p;��P<$�v=p����t�7����<�̟;}����C��V4켿H��$�����;_��>0ޑ>Ɯ��j>�=Nb ��'v��>�p��K�W��������9۽���>���>{�<>��S��>��O>�K?�.@�W�?��&?\�?? �'�mVQ��h#�ᕀ�ӌF?N��>���>Y��������"����-a?��\?ɥ�
�B�b?��]?Ph��=���þ˵b����N�O?(�
?��G���>��~?k�q?`��>E�e��9n����Cb�-�j��ж=er�>4X�<�d��?�>-�7?�N�>�b>j$�=�t۾*�w��q���?g�?�?���?-+*>a�n�D4�d���@��^?-��>I/���#?���޻Ͼ"���'����!������1���v���h$�����L׽��=�?&s?(Gq?'�_?�� ���c� ^����J\V���N�R�E�
0E�,�C���n��Y������ڟG=^b�u�C�Õ�?%?�/��A??�����ힾ+�ֽ��="���&����)>#D�����=�m�>�$����?�FH����>+�>C�w>=�4?�7�"4��w:���f��Ꜿ)>�>]Z�>zå>c�N���aj+=t�ν�U޽8&P>�v>c?-�K?�Jo?���1�Ĳ���� �&7$�rݨ��8D>7l
>(��>�@S��~ �C�%�w=���r����k䐾>�	��U�=�*2?Z@�>��>�W�??��4a��t�t���1�L�Y<�1�>��g?���>9c�>�ؽ�C!���>08s?3��>ܟ>��d���(�lon��9+��}�>���>�U?��>j�J���_�����-����Q"�'�9>x!l?����ؠ���c�>Skd?s�;������>ⲽ��&��J�Ӕ� 3�=gh?Z�!>K!2>�;���龫ov�r/����)?�?���+�+�u�>��?O��>wu�>�-�?�ߌ>�P��L�<3D?�PI?��P?
*???M�>���=s�]�H�ƽ,("�=�<Ս�>��o>�;=D��=F��?�b�e��t��;���=����W��`�㚫�P� �a��;`�@>�οbN�N�վD�/�n���b	���}�-
�<2�������꽽xb����e5.���ڽKk
�����m�X���ܨ
@F�
@�i��8��P㻿�x�9Q�&i�>�`��E�G ־}S�T�����Bm��@�}��ԕ.�g[��1�&?ޔ��;yǿ}.��a�� ?�b?F3z?�����"��09���">!I1=�M���龹j��/�Ϳ쥘���]?3#�>��ﾏ˪�h��>!�>��[>zoi>�%�������[<A�?{�.?���>��e���ɿf��'W<���?�#@7zB?$���^Ѿ�>"C?`�>j\s>黚�_.)���5��fs>��?!�=?����z�x�ڟ#<�}3?Ǣ��[�z��퟽M�>��>>�ɼ�*�{Y�>6��=ʠ�V���s��;,�C��Z�>9�%> ��؉}�����^1>�k����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�ꉤ�{���&V�}��=[��>c�>,������O��I��U��=����ʿ!$��� ��� =k�ʼ�96�|��?<��)lr�����+H]�7c�q4K=a��=@�5>�z>ݏ4>�b>\?�bn?�P�>l��=����P}��T־��]<���L��W�d���A��-���,о ���4�����%Ͼ];�`��=�aP�sގ�!Q'��Ce�vD�R/?�P>��Ǿ��H��q�Ⱦ����j࿼VH���D����/�$q�3i�?�E?�y��}pL���X?�ld����Q?�N������թ����=L�󼁙:=��>V��=�ݾ��3��P��u.?^I#?M��{������>0QY���N>��>
<�>䋎���򻸪H?��3=WS�=|�>��=1&=a?WD�>�[���Ix�%��>?�T?��m�{?��ޠ(?qǾ����8��=֗�=$S�C�ǽ@s�>%0��g?��������!�[�E?��>i�)��5���̾� �>�%�dcI?��?42��:�i?r'?�>���h��V��m���"�=��T?\�Y?{�M>�)�����4���tB?�4d?���>�a)��2'�9`+?]��?��?U�f�Z�D��I����YX`?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?x�;<��T��=�;?l\�> �O��>ƾ�z������1�q=�"�>���ev����R,�f�8?ݠ�?���>������q��='9��'�?���?Ry���� >6�b�b����O<�?�=�h����<��[4��+�L��)��oW�=4Rs>Q@�c/�W�>�I���쿄ɼ�$<����ھ��&�<)?���>�p�o﷾ʡk��<u�e&���+�Ubp�4�>���=lӘ=T��r�l�[���ɰ�|?�.<���>z��0��Ȣ�%Q��d{>��>�- >�b��# ��4�?�?�����홿����|t?I�?[_�?��&?t<�������,s��>�D?m7j?o?-���:�<ݼj���j?�B���L`� 4��7E��U>7.3?I,�>V�-�|=��>0��>˂>f
/�0�ĿӶ�}�����?P��?��꾌��>v��?�+?e�5���F����*�7d��3A?E2>������!��=���
?�~0?����&��_?�a���p�;�-���ƽ�ܡ>��0�d\�H@��
��AXe����@y�s��?#^�?d�?q��� #��5%?��>����9ǾK��<���>�)�>�(N>�K_�Բu>����:�j	>y��?o~�?j?���������V>t�}?<�>��?��&>y2?��*>�ո�}��=��>ss%>��нT�>�S?���>�/>�*��e,��@���G������J���L>�Is?9qL?�G>ڍ����Ľ��
��ь���2���6=�s��R���F�+�=y�2>Cq>"}��^�Ծ��?1p�0�ؿj���p'��54?ָ�><�?S���t�����;_?�z�>�6��+���%���B�V��?�G�?%�?q�׾R̼*>��>�I�>� ս����3���!�7>�B?���D���o�U�>���?��@�ծ?Ti��	?���P��Va~����7�c��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?�Qo���h�B>��?"������L��f?�
@u@a�^?*rhֿ����qN��h������=D��=��2>n�ٽZ^�=�7=��8�+=����=g�>)�d>�q>7(O>�a;>��)>���G�!�r��]���0�C�������Z�A���Wv�Sz��3�����S?���3ý�x���Q��1&��?`����=LK?�=]?�+{?�?�_�PHT>���?ہ=�[=�~&t=~��>,'?��P?��?�M<~"���b���w�A/���z��>��5>���>tS�>v�>�I� �1>�R8>�Dc>*�=zЈ<y}s�OF=X�!>�>��>n&�>�<>�>���������h��Pw���̽��?�����J��������Z��yR�=z.?�\>���,п�魿�eH?�9��{Z�=@,���>R�0?�DW?�_>῱���W�#Z>����h�{>>(w ��Bm��m)���Q>��?>�h>,Yt>FD3��%7�,�O��ʰ�9�~>$�5?�+��˄6�SQt���H��޾�hL>�
�>ܟ#����ݖ�>��P�i��%z=��9?�?N)��ð��/u�AC��-�P>��]>4�
=�-�=��L>��_���Ľ��H�}0=V��=��^>�f ?�b>�P�=̃�>D���3������>˼">�F5>�1?�3?��.���ý��c�z�6��N\>�F�>��0>o�>��K��f0=���>��>�n~������=�F��!�@>'ˣ��C�ې��\�=�fq��B�=�q�=⺽�)��������~?�s���刿� ���kD?�?;��=?<&�"�_����(����?��@�`�?�	�[�V���?Z;�?����ݍ�=�d�>���>��;�yL���?țŽ�ܢ���	��_#��Q�?`�?џ.�Z̋�y	l��>�o%?כӾ���>'���T���タ�����=>"�>��P?X��(zֽ�ax���?�i$? !¾d���&ÿ�0c�D��>a�?�k�?��d�6���
Q��)?��?��;?���>�C�"߀�a&>kN?��W?t��>7�2�՘4�.��>���?{�?�I>/��?�s?jm�>�+x�YZ/�&5��2���=v=�'\;�f�>�P>����LfF�\ד��g��w�j�S����a>��$=t�>i>��1���2�=����J��[�f�K��>J,q>u�I>aS�>!� ?�]�>���>�{=.r��䀾����r�K?~��?6���2n��L�<"��=��^��&?9I4?�p[���Ͼ�ը>�\?N?�[?�c�>/��>��迿A~��&��<��K>+4�>*H�>t%��EGK>��Ծ�4D�lp�>�ϗ>�����?ھ�,���h���A�>�e!?C��>iҮ=ř ?��#?�j>�(�>;aE��9��0�E���>���>�H?�~?s�?8Թ�AZ3�����桿<�[��:N>w�x? V?ʕ>Y���߃��beE��>I�����d��?tg?�S�?%2�?��??�A?�(f>���;ؾb���a�>�{!?F���v@�y�"�����?�?���>�J��(�ֽ�I�������8�?��T?�%?I8�er\��Ǿ���<� �����y�";��v;r�>v@>�,����=$>��=p[d�F?��t�<X�=
�>���=Ѫ1��C���%,?��2��₾���=qGr���D��,>>�I>ל��ӷ^?�1;�;	|�����kZ���/U���? ��?OY�?�ֳ���h���<?��?�z?���>nO����޾��0w��z�ō�6">U��>nS�6��iC��nB���Q���;Ƚ�q��>�w�>�?n?��g>���>+��ʷ�!���^Q����P��!���.�C*:�iX��v���+A���T�h�ξ�������>����"־>�q?�~>mAc>�m�>/�\<�r>��@>�7[>Ę�>�F>Tu.>���=I�/�6�d��D?[Ӡ���2��%���۾��O?��*?���>*�S�Ղ�
��@?v�?1ȑ?�-�>,�L�dq*��f?'��>{-��{?�>��={�¼��½qA�����AnO��3U= ��>��۽�L7��2�Ԓ�c��>!�?�.�<Nپ��<����� o=�L�?��(?��)�g�Q���o�4�W�aS�m��Dh��d��K�$���p��쏿r]��<$��N�(��*=Ɇ*?��?u���&���$k��?�fbf>F �>�)�>lؾ>�kI>��	���1���]��L'�����kN�>�V{?���>p,?�df?��|?�P?^\>s�>e����>Z�a���>�0�>�?> >?���>���>�6&?s�=�2��Խ�׵�79?�-?�??�f?S ?=���S��鄼-'ս�]�k��� ~��HEs>҆Y��m6�6|j<z�#>=�?�݃=Q�޹H����q?�c=��A?��9���J���B?��P?8-?�|	��8V�+����&?��&?cl���F=�!>��=H=	Q���S>\�:����=i}A>^y��2B=��<=0��ؓ=A�ʽ�L=fB.�9�<���>	85?<�>ҘS>ȶ����31�����ǐ�>��>A[>n�ľ�����'��&\��)�>TX�?�8�?6>M">1g�=���N����
��٭�ѦD=&n?��>��9?Գ�?�G?�k.?��f>���L���p����_���?B/?��>���>qv��Ȅ������
?tq�>4[�A�b=�AT�U>����Jڽ}@���^���B�o��>��C���.Ľ�\�?���?����d3�uR�
���]����LT?I'f>D�S>��?ܤ)�"�;�3F"�~�>�b�>�+4?nG�>H_N?�a�?Lk?���>Z�=�垬����9?<7-%>5>?-"w?,��?thr?��>��6>��ý�Zھ*���2�t�*����K�&=��[>�E�>���>U{�>'��=��.�FV����߽20�=�Kx>�}�>��>W��>rBV>)����A?�\�>����;>߾�E���+�`��6_?yz�?}�?/#:>� .�T�����0�>",�?�>�?�r?���F(>����Ѿ:钾H��>TI�>4�~>#�P=Ȑ����>`�>l)�>3�9��+�#����~��>�HE?��<�g��)���H���Y9ȾH�]��i��}��m����e���?�����F)�����r�'����� �O�|��OC=]��>&���#�<��>�x�=uI=x�>��?>��h=O_#<Tl^�u�;{+�=�̭<gSs��Ky���>��->�Ύ=�^˾/�}?�LI?k�+?�C?ciy>3n>�H3��Ö>~G���6? /V>-�P����gO<�&���i딾�ؾ�y׾B&d�����>v�I�6�>�3>>��=Ɖ�<n��=��s=!L�=�2a��3=���=Sk�=��=+��=��>�@>�6w?W�������4Q��Z罤�:?�8�>a{�=��ƾo@?��>>�2������xb��-?���?�T�?>�?Bti��d�>M���㎽�q�=J����=2>k��=u�2�R��>��J>���K��E����4�?��@��??�ዿϢϿ8a/>%ݒ>ĝ>��M�x�+�B���]��/��(4>?E�[��e��W�>�=��b߉��'�^؎>?��<�h>	Ѯ=�/�*K�=�~$��j���%���?�A�=Ú�<�@�Y^��$�<�
�;���>�T7�?��=�-P=(��׷��|�>=�T<v��>��?��<?G/h?֦�>�<޾e��m�����>�)�<��?�V�;�!��&�>�B?TJ?��[?���>m��k?�?6V��Q���d�վN~��_(�� �?�r?�Ѿ>�h�=� 1��-�f�h>c)�>�?K�7?IZ>{�}+�K�*�ڐ+�6�<B���O>��J���3��u�=��'�1z׽E��=r(>K�N>?��=��=2�=)@{>>�>�So>�2=�õ��_7��v"=k���s� >Ǩ�$�a���l>%�ܽWFC<[�ۼ� �=�A>>�$���&�<�_8>h�>F6>e�	?c>.v���A>'�辤�8��aX>,"���3I�io�]T�v`B��:���Ó>���=�3�+׌����>��>��>O[�?�?R?>'��n���͵������־ zK=�0>��_>�"���W��1(���j���Ⱦ�8�>�>&��>ˤ�>��ھ�!���>�c���'�v�?F��ˮ�=��,��po� ����я��Kd�@����
�>AB��X"޽��?�L?��??v�>�X佌��;���>�6���T>d�U�I
�a�%>��?'S?��>GG������ A̾����۷>/I��O�������0���Jȷ�⊱>
��о�&3� f������k�B��Fr���>��O?��?�Db�X���SO�Z�����Ep?zg?��>�J?�??6��r�!v��YH�==�n?���?�;�?��
>��P==aV�m?>/$?{Q�?Bգ?���?� R����>n����<��b��={/V>�������>\�>�q?/����%�;~��c2���S��q�=Ǒ1>�~>I�>��|>[7>�>�"9>�ѓ>No�>-�>�C>T�!>�zI>�����϶`?F�H>��W>�X?]Xi>ɂ�>�BG=�	z=�}J�����aPֽ��ɽ�)��ZnA>�5L�.�j�s��d��>윿����?̯�=�*�,#8?�%�U-����>J?w��E9=�X�>�F>�@�>�"�>�?!>���>䇶>�
��Sz>���i��ۏt���?��;��>�ϼ���1�����ҐH��돽�����d��̡X�	b�E�<��Y�`ؕ?��\��y�L6��n�=.?*?䟣>�wD?�s��oK7�!����?�w�>�fľ�c��
���Ͼ��?9�?�`G>o�>��q?��(?��*��/��V���g�Q���K�{y+�Sy���|����������?�E�?��5?���=֩j>��?l^2�2Wk�H��>�%l�^�%��EW��^>^`P���ڼ��������o���Se>��;?K[�?�?�|��m֑���=�38?D�3?��}?@E?5e?�\�a�*?Ѐ	>q��>�a?��/?�S3???�>�,3>?�`=*���,�=г��{8�����)�k�%�^N<���=p��;3�+=�Ի<+�=�'�<��ٻ&B�<�⮼ �o=��=�
`=�>�=
��>�^z?�( ?&O�>�U?<־��6��d�:6j?*�?j�>��G��!'�X�n�TGL>s�?_�?��N?�T�>0��8��T�ڼ��+=h?>�Ԍ>z��>.ǘ�b T�WM>����=:>���>���<&�}��^�^)̾J 9=�,>y��>�<|>o���WJ)>�Ϣ��`y���f>�Q�`K��h�S�d]G��U1��9v��d�>p�J?�N?���=9&龞�m:f�Ǐ(?O<?):M?t}?r�=��ھ��9��@J��/��h�>;��<		�Eg���䡿Ix:�XՔ:�q><����	����>���*6��~2S���2���:�=9� �*&�=+޾�P	�)�O�̽��==������ȡ�mۭ��$=?�A=�����h�8t�>!Ӛ>.��>G3x����=r]������-=���>El�=�z�Y�ݾh��D�b*�>E?i�_?%?�?������o���H�Ϳ�t�u��zܽ�]?k��>���>>'h>��&>�����}����U�\u'��]�>*#�>q%���`�Kl���u�0%�Z �>��>!>,�>˒G?��?)d`?�>9?{��>��(>���پ!w.?�҃?���<G�*�72潬ZW�R�P����>��2?FH#�R�i>��?���>l�?/
g?O?١2>(�¾�4�yD�>Y��>��d�
���r>E7?Ԙ�>�;M?��}?��k>�?6��#s�I�W���8=��=J�/?0-?=U?��>X�>������=+e�>?l?��?�̀?�P>{�?�n>��>��;���>�i�>#?�@I?�f?[�B?�<?�ڗ= b<Y�<=�s/�$L���=ף���>�<o�`����f�G�=Q�"<2�w��n�=0JX��o_�l�-���F�je�><��>�!���V>~����{�{KO>���M�n�M좾w=��G����>��>�m>�.�������<p>&�m>���>��>�Z?��=?9�Ծ�|t��?��bֻK;E?��I?��>V���<��=O�mý�E�?�*�?y$���׾5�b?��]?�h��=���þ�b����O�O?��
?��G��>��~?Z�q?V��>,�e�6:n�*���Cb�r�j��ж=@r�>0X�#�d��?�>>�7?O�>��b>F$�=pu۾��w�yq��h?p�?��?���?'**>g�n�34࿉���H����Z?7��>�@4��;?g@�=�����	C��-��i�oa��aY��>�����t�\7�[���*��I>v_�>m�g?i�^?LU?7c���(\�,�L�M5��v#9�&q�33�a�1�J�2���U�^zi�&�!�*��������.;��:m��k�?�&?mD��B?�Y�=� ��S��1��>|���qX��ɾ<ky6�׋w=�J>��^�+r��j������>���>k��>�G?w�1��B�� ���x����C>i��>�>/�>�4<�dJ׾sn��Ѿ]���>ъ��w>�b?��K?Q�n?U_ ��C1�P���RE!���'�e�����<>Ӣ>P��>]MZ�L��"$��>���s�h#�����
���=W2?�y~>��>�,�?(s?���W��"y��U1���\<�W�>R�i?i.�>爇>ɢʽl�����>�bm?�$�>s��>���ȅ ��{������>��>���>$�s>�3�j]�'�������&�3��=U�i?�}��r
h�l �>N�V?�O�::�Z<X8�>Qu��d �Y
 �\�"�1^>��?d��=��3>������	�J|�(���r)?�u?�<���+�jV>l� ?}��>ʴ�>8ʃ? %�>�¾�;;Y�?'_?��I?�@?���>��/=$Ѭ�w]Ƚ�%��s,=H&�>ԧ[>;�s="P�=�+�_�X�::#��=I=έ�=$6ռ�7���&<�D���>O<� =&�4>�r��KM��0ھ)�-������-���>�C�v���o�"����+������pٽ�������"�s�w�h�0�ľ��?�'@�����澁'���s�e�(���P>�6���낾��;�ܾ"���(��&��L���d��у�9��%$?n'��jjƿ�@��t��Mr?&G?\v?M��� �f�8�!�>":Y=ê���P�qL���Qο����}{Z?40�>���M��tb�>|n>��W>�z[>2����@���O�<rI	?Q�+?���>��j���ȿ跿28=�u�?��@B�G?� ����0�;1�?ct?��>��^��+�u0u��o�>��?02P?�Ȓ�p�F�!]=�jQ?��b��w�})<m�=�p�=�ɽ������>�I�>X����_�̭2�Qf���>�EU=Qņ��^���>I_�;�e��Uɾ1Մ?6{\�cf���/��T��^U>��T?%+�>�:�=��,?e7H�_}Ͽ�\��*a?�0�?���?!�(?Nۿ��ؚ>��ܾ}�M?`D6?���>�d&��t�
��=�6ἕ���t���&V����=a��>H�>�,�����O��H��U��=(�R�ʿF� �}!�Ku#=��<��Ĺ3dR�1Ғ�~���sP�O:�E䠽)��=H�=7})>tQ�>3Ȅ>Q$Y>�\?��v?��>#��=I�O�ϛ¾��O��ל���1��_�.��f��w�ξ�����D����2���� ��8�_~�=�VM�k����H�ךU�C�W��J$?$��=&u���>.��E3�7�h��S��,�$=� �(��[� ��dq��Ħ?�K@?le���O����D=�X�:�M?[MC����c�����=j�\=|.a=Ma�>H�<=��澳|�
4�K�!?��?�Ͼ^|���
>�K�}��=��$?f�>�'��}�>#��>�c��.$�=�	��ǁ=���>$��>�N�=����o(���J?��K?b�4�G,t��f>U˓��X����=ǳz>�����Il�w^��V��;'\�����<�$}��∽�<?��>�,=��*�N֊�X������b>?�f\>��O<� ?�,?�r"�t1��s������<v�#?���>=�>j�6���*9�0?Z?�[�?�_W?�벾��K�`
\����� f?#o?�hS?Lt�y���X���ݎ־��?��v?s^�xs�����S�V�c=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�$Þ?��@���?F�;<��W��=�;?j\�> �O��>ƾ�z������@�q=�"�>���ev����R,�f�8?ݠ�?���>������r�=I��_޹?lU�?o���l�=��y�h����|�n>�M���4/���H�/3�k�;�>�U��B��\H���(����>� @�����A�>Pk���y�Y�Ͽ�[��/����#���?�"�>Lô<���ƈA���-�������������>w��=�$�u�a����(��*E�a��>+	��?E�>i�o��������Ɔ���>��>Mm�>޼;���ʾ�O�?	3��?��畿z��Ym?��?x��?��?�2�����0�nqh���@?�+x?G:?9o+�T����Y=��j?)_��dU`��4�VHE�9U>�"3?�B�>1�-���|=>G��>�g>l#/�`�Ŀqٶ�����?��?���?�o����>\��?�s+?�i��7���[����*�5�*��<A?c2>A���e�!�B0=�^Ғ�ż
?Q~0?�{�].�l__?�b�4�n��u-�#pƽ���>Jf/��-V���ґ��!f����z�ロ?�8�?"�?!N���#�w�$?��>�ɗ��4ž�O�<�Ĩ>�o�>��O> BW��s>S��x�9��s>�Z�?Y��?!�
?p�������w;>��}?� �>bB�?J{�=���>�w�=�۬��tV<M�>�� >}�s�\��>f�H?��>��=�9>��/��F��UK�V��	WA�:��>;�f?D�L?�F>\�P�M�Ms�����L�����L���>������>�R>�b">?k?�NNҾ��?ck��ؿ�h���'�^.4?t��>p�?���L�t��N��+_?���>�3��+��"��N���?L@�?��?پ׾��˼�J>zܭ>qA�>uEս���󆇾��7>کB?*�C����o���>5��?Ͷ@Ю?��h��	?���P��;a~�@��7�1��=��7?�0��z>0��>��=�nv�Ի��$�s����>�B�?�{�?���>�l?q�o�G�B���1=M�>��k?�s?^8o�8�ղB>��?7������L��f?��
@wu@V�^?0���ܵ�������������=E�Y��l>)�j:�Q�=֯<ϰݽJ) ��4,>�l�>�ޟ>���>ߐ,>E>)�>���X+�����1y��"<��x��&���#��佾f[��Ӷ.��\v�=:���w����1��Kkټ0c��a��L �=��T?�T? :t?��>����&X1>Yl��>W=+)��/p=�[�>��/?�|K?�4#?Fޅ= ��u�`������!��Kۉ�h��>�M>�|�>��>�ͫ>؄<p?>cA>���>��=�3�<��!� ��<�@Z>U�>��>/v�>�<>��>g������h�h���v��Ͻkܢ?�ʝ�edJ�F�K��H����M�=1-.?>'>q���4�Ͽ�ϭ�%LH?<������*���>��0?�V?�D>a6���P��>s��m�i� �>�� ��Ml��)�k�P>ˑ?�K>��l>��1���9���c�>���� 1>�*?��ѾE�,�6�l�Q�L�s���#;:>�י>�↼o,��.����u��LS��s=�6?��?�����������0ܕ�v�1>�p>J��=��_=�7%>.kZ����n<%�[�=V��=L�}>�/�>Ey>�L=��>����#]����>�Ȇ>׳�>�?,=M?7����=s��q���AQ�-Z�>�&�>���=���<�(�P��=�� ?�Iu>��_��A��_����y�u>�ǒ<u� "J�.%����v��4�>+��>a}�Ꝣ�3��<e|~?𿦿�ӈ�J]�Z����oD?��?a6�=��S<�#�즿G����~�?f�@Aj�?�D
�ӷV�&1?�֍?����0,�=ɳ�>��>t�;�dE�+�?��̽�6���4
���!�%կ?�J�?%"'��t����l�g�>��#?رҾ���>���qC�����vw���0=4)�>P�H?�f��BYX�}X;�=O	?l?3`�˲���ȿZu�q��>;��?�?; m��
���i@�/��>�?�3Y?��k>�oܾN^�ą�>�B?�AQ?˹>�{�y�'�8?
�?�T�?kNI>7l�?#Ns?��>xx�P�/�� ���(����=��<;rq�>�, >�k��cqF�8���X鈿t�j������`>�'=Qĸ>�f��h�=Jg��+���G;_��>y�q>�:H>�U�>�� ?��>71�>�=����Ё��N���K?ñ�?r��]2n���<���=ħ^��%?�?4?�#\�n�Ͼר>}�\?���?k[?�T�>��L:��w濿|��>��<�K>&2�>lA�>,���?K>��ԾP$D��p�>�͗>�O���<ھ�,��nj��-C�>�e!?���>�ۮ=G� ?�#?͏j>z%�>vbE��8����E����>��>(G?X�~?��?Jй��X3����c桿/�[�a?N>�x?V?�ɕ>�������uE�=:I�풽)��?1rg?L]�e?�2�?�??<�A?X$f>��9	ؾ	����>�� ?�e��@�{-$�rB�\�?��?�Z�>�6����ڽ��@�\{�+x���?<�Y?d$?�U���_���þg��<���ݨ�c�;��r�ӛ>�	>d�v��ǯ=��>�h�=$-p��,6�X<�6�=u�>s��=Rq?�4A���9,?��E���	��=��r���D�ڜ> !L>�����^?z^=�;�{�g���x��,�T���?O��?zj�?[ش��h�c$=?��?��?{A�>�6��9�޾��w�*�x��_��&>��>�gm�|�d���׎��OA���ƽ�F佱'�>
�?GX?�E�>��>�c?y ھO�Ⱦ�
�k�"��+R�#�4�U�1��+a���+�;TǾE,�.���p��]Z��`f >2�N�tb�>]�1?�އ>��">���>�������=���<�&�=G~S>:���g���=E沽3�h=G3J?��|�3�3�0༾�T��S?� m?���>A��(�������F?�g�?�"�?��>�N��݆O�,��>(��>9���)��>�S>�W7>ϑ߽�z�5(4��%��=#���>��ܼ��=��s$��ߙ�Lo�>�??�)��`+ɾ����򌠾o=MB�?��(?k�)�B�Q�*�o��W�!S�;c�Mh�	�����$���p�}쏿�W��A"���(�{.*={�*?u�?5~�N�S4��Wk��!?��_f>e��>�/�>b�>�PI>��	�>�1���]��9'��~��0G�>�`{?� �>=�G?��>?��U?��I?��>e,�>�\�����>Ǯ;�֞�>Y��>�4?e7+?NC*?)6?�(?4�`>Ʋ���:��2�پ�
?�|?��?Of?�w�>��OʽCD���1���	~�dK��E�m="Ԅ<V�Ὓۀ��DI==XJ>��>��9>|�V�{�H�P��=��b>	�J>x@?�"�Z8����>[q�>*!?��0?�H�R�q��� �%?�<�>w?s��2�=��B>��q=iJ�=��ܽ`bl>�邽��>޹��q)�l낽E>\8������~�=K��<�O�G%0=��>m�?M��>�ч>'݁������MX�=��_>W�]>H@>�Ծb�������Q�f��;�>�A�?�?�=� �=���=Ot��������}��m��<�?&Z#?�2R?�?��=?6�!?)�>���1l���w���ѡ��W?).?�>�
׾����s%���q�G��>scQ>au~�ʞ=V�^�kS��8X̽D�p=w�]�o�%��ت�o%��Id̾�'��2
����?�?�;��,�q���{�.�+�1~�?��G>�&i>��>��,��+�о}�J>��>�,v?ݏ�>U�O?�{?�(b?m�u>%C7�F̬�1=���<�>��<?��?k�?b&u?7��>ե>�*�?�پ�C�1�5,�J���es�<cG`>0��>Ң�>���>�J�=Gdؽ��ý��3����=��}>�:�>r�>���>�|i>��-��@?h5�>�����̾�I�žb�H��O?�
l?
�B?�=)*�sp�͙!�f�>��?8\�?�$�>�@�7\>�ŷ<'0ܾ�3��"7(?%��>l��>^{*�������=1�>}�*?���(?�O�'��:���"?�?��G�9GĿ�ap�c�k�/����^<�����nb��_���yY�D�=����H���n��?�c������G���N��^p����t���>%�=��=�x�= ��<~OҼVQ�<�$.=>�<�=�S�"��;&�N����.���a�����<bsO=��3�ߴ��szl?��Z?�K?�-?�v9>��>rĽ�0�>ǽ��>xp^>8�������|��az��+����J����Ҿ�6a�g_��z7>R�q��6�=8�4>0��=�{�<��=O5�=U�=�~���#�����;�y�=T,�=�Z�=v��=��>�6w?X�������4Q��Z罥�:?�8�>k{�=��ƾq@?z�>>�2������yb��-?���?�T�?<�?Ati��d�>O���㎽�q�=L����=2>v��=q�2�U��>��J>���K��A����4�?��@��??�ዿϢϿ7a/>�&E>�JT>�b�L"8����.����=�;'?��^�<�ʾR��>�)��%��⊽��>�.�cm���K>��H���>��<c�ڽQ���7��>Wm6>3UH>U���傉��Ǵ<Ә�< ~o>p����Ő���=Ҁ役������=A�g��	�>�?�0?�bS?ib�>?����/����U�>)7O>�Og>�Ǟ=���=�>�Q?SX?$|J?��>�}3>���>�g�>Z1U�����=Ӿ2������P�?ie?��>�Y�=���V�z]��<#��>�!?�T'?bR~:��$��� �0~�����歽'ﺽ��A>j�ͽ��5>�4K;����EV�D�>��B>!�>͹>�o�>���>?��>�C�>/��=��f=Vc�=�
6=E�l=.��=��=�O�<le>T1u>S�=�����)�9~ɽ�����h=]�=vrڽ#��=�5�>8vA>�Q�>ř=<���%P>h���J@�&��=Ԍ��/�>��f�Pz��2� �E���+>)�H>���������>�YM>I�H>]`�?�~?V*#>G'�n�Ѿ���ꌃ�
�k�19�=��=хm��dB��[�_�J�Ĕʾ���>Ox�>Jͮ>?�v>Z:%�#'@��.=)n��N5�l ?Qʱ�����#�!q�[A��NV��e�e�bQ��\?4?e���.��=�[�?��F?+��?��>A��������>�&Z��7�<�1�	h}���ɽ/x/?6(?�?+�˾�U*�$̾/ɾ�ڡ�>�MI�XAP�뮕���0���!��/��ű>L���&9Ѿ%�2�vS���돿tEB��/r��]�>1bO?���?j~b�&����N�������?�|g?
\�>�J?An?�c��N��o���5�=%�n?ϳ�?n�?:�>_����
�F��>�#O?��?i>�?���?3
����?��Z�
7=	{��^	>(��>ᾤ>=c�o>��*>r�e??3ҽ�K�������=L^�mlڽ�ռ�B�>_�h>N��>|�>xnQ>Nڛ>��??�?�^�>��>�$?!�D�&f �̲i?���=r�I>y9? �i>���>��)==��>�j���� ����D+�N��=A0�>(=񺘾Aݖ�"�>�iԿ[ɦ?*>HƸ���`?`Ls�K�>�n�>��=,3<��R>]�_>�E�> [�>�\Y>��N>~�>,�>VھA{)>g��:�=�`Ue���D��/�#�b>�J��j/�nq�/[h�sTC<�������9�^�*���-���q���?>��X�- �'�����?�>�p ?¸Ͼ���z�(>;�>�V�>1:Ͼ�����5o������?�g�?,�q>~i�>�&p?�$?3Z����N��˅�V�����b��e����O�(�-��a��V��?�x?�r+?��->͢r>H��?i�E��k���}M>�U���9���`;���>�}��3n�о8�޾�뽞n�>6s?��?��7?8�ླྀ�T��l>y^@?7�;?�hp?��-?�G?�'�ŧ'? �>Ef�>�?d0(?)?�j�>]>�t=�L��ɍ=y���;��$���t���V�����<5�=�5�B��h4=�<!�7�P-��3��������<�1�<� �=���=x:�>@��?56-?M]�>��D?pԞ��vK�Iwu�y
n?�w�>�c=*F�>��L���A��aɽ�Pk?�\�?��J?�?��0�%���l�=���>�AK>�~>��`>BFC����`�-= �>��>��V>��d���њ��a�\>�(�>O~>�u����(>�8��)o�W�Y>��A������=��@��2�RZ��Dn�>��G??���=\����ְ��Ma�(�$?�$7?�uF?J�?s̬=�hѾ�+?�&8M��{���>�j�=V�ֹ��:���9':��Wu<�x>�������Zp>���D̃�u
g�h8��-˾���=z*�>j>j������U��SaH���g<?�I��r�P���4����F?*��=�3��\�k��_ľ8�K>��f>+��>_��� ��=?K��L�5G�;�w�>u�>�=�ھ�Z�M'����>�A?"�a?z�?��J��Uv��3A� 
��j���{��li?,ؼ>U�?y�>v��=�ϵ�=V�!a��8�l�>){�>~��wL�O��N���>%�M�>�+ ?\�$>))?�UJ?Y�>/{L?M�6?n�?I	�>����Ͼ#4?���?�|�=0�K����35��2n�� ?<�B?��r�ES>�A?MB�>e(�>��y?M�?�>Y���I�(�讠>5�>-�i��_���4N>��I?*�>7~V?�V�?NbK=���,�;�C_�r4彃	>�0?��>A� ?��>���>�X̾Q��=��>�-z?��?ת}?C�+=�?V�>a{�>|)�=��a>��>r�,?)A?)�_?g�J?��?��<�5}��ꦽ������ΕͽXC����U=M4ݼ�v1=�dM<r&f=G�.=��z�\��=�Փ����U֤�%��<8��>�o�>�ƫ��Og>���������>G�;�6K�/Z��ob>۬�=�>Zy�>y^>R.|���ܽ�,�>v��>Y�$��N�>��U?�U`?N�>�I�|�Ĝ1���"�E�(?xY?f��>�聿:����1��s<��<X?���?^�� �%��b?��]?�h�:=���þc�b�ˉ�O�O?]�
?B�G���>r�~?��q?k��>�e�:n���\Cb���j��Ѷ=kr�>#X���d��?�>ӛ7?2O�>��b>�"�=�s۾'�w�]q��/?]�?�?w��?�(*>@�n�4�&w��B��v^?L��>�D���"?������Ͼf0�����d�� ��(��DL��r����$��׃��"׽��=�?ns?�[q?��_?î �_d��7^�U��n[V���O�u�E�lE��C���n�xU�S ��[-��<�F=�Y�E]���?n�+?��/�=;?�vs�>����M{��վ>7���t��\>P晾R}>\�>�I�r�{�Kaþ~�?��?|�>�~L?��'�.1>�!�:�Z��W۾oPR>�
?�)�>��>k���5���������ݽ�<3=^ v>�Xc?�K?.o?0.��0$1�u�����!���1�����@�B>#�>#+�>�OU���^%&�7>��r����l��b�	��R=�2?l!�>�\�>8E�?��?+�	�C���?x��1�56�<n�>�3i?���>�%�>6Խ�� ���>�dj?o��>�G�>�t��� �̢}�R�����>/��>���> Fr>���uO�}����l0�#>��i?B���]$b���>i�T?��<-Xj<Qw�>����)����--��&$>H�?�(�=8�D>�uѾ?��l����⇾@�)?Ƨ?xߒ��+���>�� ?�r�>�ޥ>N��?�u�>�+¾\<P<��?�\?F�K?pyA?���>y�+=E���|ƽ��#��=|q�>��W>np=B�=9�� aY�H�#�-�R=2�=V��2>����;-l��VJ <�\�<�V;>.wٿ�oI��1Ⱦ��$�L�����Rg�ǡ�=�4��|on��]Ⱦ�����:��`�[�b�]��0J��؊�Cw��v���C�?�@�\t�9�����������f ����>����lm����������$о�
��|�׾B</��Ar�$܋���'?���˽ǿK���$;ܾ� ?�@ ?L�y?9���"�y�8�ϲ >�s�<������Ś��J�ο����~�^?3��>�	�+�����>@��>ԡX>�Kq>���瞾+E�<��?��-?���>��r�I�ɿx���N|�<s��?o�@�,K?֦����rշ= �?�#;?�۾=SK���Y���Ѿ���>��?~�e?�੾3ۋ�5��[a?~���8������u�>��.>=b������Yx=N��>hpW�Ev����o�k�"�^>��=�DξUع��#>����M��b��5Մ?,{\��f���/��T��U>��T?�*�>R:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?:ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=p6�݉��{���&V�{��=[��>d�>��,������O��I��V��=nF���ӿ���V�����</�q<���;lɀ����������t�z�x��=@_P>�4:>l�>t�M>焣>`?�ԁ?���>�K>�~#������?�ʖ�����j��A�<�����gM��4�s�-��9���/�����ZSr��7����=�>�'��^\<���i� �T�eK?��X>���%�����}۾�Ȯ���m��$��O��TF'� hq�Q�?i�9? �����H��/	�r�=*?q�_dT?A�3� | ���C��a=�_�*�w=���>w��=Q8��q��]B�_�G?�x@?�Tվn�����>.L=Ƕ">zs&?��??9�����>&�p?Xg��k���&�>��U>_�:='�>3�>ң��Ӯ`�.�?�\x?�h�\����%?�3ľ�0���v>=ލ�>�fþ 7E�P�_>$qd��Ӳ��1�<���q�=
6?N/�>l ;��(,�0 �1��<�O����?IÒ>��ӼLcj?��>6,�=6&g������+��B0>��B?�K ?�A>ʞ���P����ھ��]?�Bh?��?u��c�4�)uK�����L?��?�K(?����B������O�5'?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?p�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=����Q��?N��?�.�����=��kk��R����=j��<���d�$��s���#�"b��ׯ�$���.A�Ɇ>ֱ@�/����>W6�Ӕ�Mhȿ�u��snҾ@}/�̀%?��>K�������vX���a�����/�_���t>ΏM>�m2��ҩ�e���6H8�����S�>��!<%>���=������5�5��/>[t�>���>(���@H�n�?�ા�ɿU����ξ_�X?[��?Ѽ�?�!j>��S�F�N�@P!��#>�oS?԰r?^&?�5���x<ƣ�=ϴj?nL��rU`���4��GE�)�T>m!3?�<�>��-�^m|=�>���>�>/�܀ĿNӶ�����k�?��?�t����>���?��+?�n�54��hc��#�*��6��->A?S2>-����!�a.=�.ܒ�q�
?cz0?Mt��&�9�_?�a�Q�p���-��ƽ�ۡ>��0�7e\�)Q��Ҥ�aXe���&@y����?3^�?C�?%��� #�I6%?F�>\���,9Ǿ~��<��>)�>�*N>bF_���u>����:�j	>���?�~�?6j?������	W>��}?m�>�˃?
o�=���>#��=�S��H-غ�7$>��=u\C�[�?�6M?r��>�2�=�,3�V8/��G��O�� ��?C���>_�b?2]O?c!S>8Dɽ�L�#�!� ,��ۣ'�b�f��H��XO�f齝�$>@�O>m�>hG@�%�о��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Qz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>;�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��@a~����7����=��7?^0���z>��>,�=�nv�λ��b�s����>�B�?�{�?���>�l?y�o�]�B�d�1=�L�>��k?�s?�=o���R�B>��?3�������K��f? �
@xu@4�^?'�xۿ���}�������_��=��a=)�^>g����r=nr�=p�
=V������<*bY>d�\=��>qQ:>ZQ[>ne_>'��h�-�[;������K(O�)(�g��u�n��.0T�ԧ��&��ݼϾ1��4 �ߟn�Z�����6��Z��=IwU?�1R?yp?� ?'�x�� >����n�=��#�>��= �>U,2?��L?�.*?Բ�=�ɜ�޸d����$���B0���7�>H�G>�!�>s��>Q�>X|#�YH>�N?>��>s>�M)=Sꥺ�#=�LN>܈�>9s�>V>�>�H<>�>δ��0��p�h��w�y�˽���?a���d�J�L*��i&��u�����=Sd.?k+>���85п{�z)H?����R�ۦ+���>��0?~aW?�n>����f�T�{.>L���j��;>�[ �8l�F�)��Q>	j?pq�=NYc>X���9�1*o��@�A:N>& &?Rѯ�� �\�e� �R�,�ƾ�W
><�h>g����*�?r����}�C�N�f��=�^@?�?'�	�	��������۾4�>�.7>�	?>�Q�<�a�=����>�;�>��`>Y[�=�=QZ�>	�R>p�=#��>1<��y|��F��>mN>H��>�#?q�<?��V7z��/y��A��ίI>1�>�kl><o*=�@�!1x=�{�>2�Q>��2��3꽱"�����.�~>#����l�y�f�Z0�j4�,^=�$>>~=c��!P��~?���,䈿��e���lD?C+?� �='�F<��"�: ��fH��F�?n�@m�?��	�ݢV�G�?�@�?��2��=�|�>׫>�ξ9�L��?��Ž?Ǣ���	�m)#�cS�?��?��/�Mʋ�@l��6>�^%?�Ӿ*��>)2��B��������v�G�'=�̹>��H?�E����v�=�9��	?�?��X��6fȿG�s�-@�><��?���?�l�mx��*A�I+�>u.�?n�Z?�\l>�v޾�g�=ъ>љB?�R?�)�>�x��/�kJ?%[�?�9�?��H>h�?dcs?�-�>�z��p/���� U�����=
-X;4ߐ>�w>�Y��o.F���e6��=Ej�U���`>[
$=��>}Y佀���m�=WҌ�����a�ز�>!�p>gbJ>�]�>Ɇ ?�=�>l��>��=}���D����)����K?첏?���2n�R6�<3��=��^��&?�F4?�[�V�Ͼ�֨>��\?
?P[?�^�>8���<���濿�}��W��<�K>|5�>&D�>x2���GK>��Ծ4-D�
q�>�З>��	Bھ4.������5D�>e!?`��>�Ӯ=� ?.�#?(�j>�$�>�aE�e9����E�"��>���>�D?9�~?O�?Q޹��U3�"	��=㡿��[�W>N>��x?/W?'̕>���������F�FI�����?dkg?�T��
?�+�?��??�A?+If>����׾�֭�O��>�a!?5��\VB���&��4��1?�?0l�>�����ӽ�S׼2�5����?�\?W\#??K�`��������<|U/��L���<��Z�x�>�N>�*���	�=��>2?�=1l��16��6=<�֯=6�>Ս�=-8�����-<,?uDG��҃���=��r�xD���>�:L>����_�^?i=�.�{����u���
U����?ߠ�?�j�?[�����h�� =?��?|?n&�>G��'{޾���N^w�Ғx��r�|�>���>��j�K�[��������F����Ž�����>���>F�?=C?�,`>��>
��?�!�G��W����^��<�,8�L�3���Ǟ��)-�,G�����(턾ec�>�%��Cƺ>>V?d^d>)t�>w�>�<j��^}>j�I>�e>��> �<>g�4>�>�<�u��Md5?�0x�:U��J)�9;����!?ȵ!?9?(Y��A܁�&ھF�9?�?��?�9�> ��Gd2��$?{��>�d<��2�>R�u<�FE==��=\?޾�#=ez����D�?�}�������6�����?~��>ӟ6=<x��><����o=jD�?�(?(*�z�Q���o�>�W���R�I[�
�g�𝡾1�$�O�p��叿 S�����!�(��q(=�*?x�?*��pm����U�j�I?��f>��>��>"�>\8I>U�	�ؽ1��]��<'�#]���V�>38{?�G�>Fx/?7�S?PO�?�]C?�\/>��>3�!��?Ӹ���"�>@�>�t?��M?��>]��>2?�R�=/��_K�������>S�>��9?*�?\��>���e�^�;�ϥ��·��؆=-(<>��ڽ��	��E0����C�$>(�?�~>�T���!�p��=�;�>���>??��2�z��X�>q�>�dU?��"?�}~��������1�>��>������5>o�'>��C��8���>��[��>����a���gS;DE�=^��<MS)�S��=/޽�q��]�=!U�>.�?>�B�>����� �����=��Y>�S>�	>MKپ�{����Q�g��Gz>l~�?,q�?��g=�D�=�8�=ٽ���t��ݱ�V⽾M��<��?�E#?:T?�}�?V�=?�#? �>b���J���3���ߢ�}?fM)?�(�><Nþ�eξh<�����~?���>��V�����t|�B�Sc%��:�=���xB��L���Ќ�v߬��%���9����?U�?���LG��?ɾ-�e�#���-.?F+�=�a><��>�)־*E�������=��>>�b?x!�>�E?嬂?:t�?�.�><�;�Vۦ�n��1����<-@&?�$�?|`�?�ő?�ؾ>A�=���ھ-t��f��)��F�^��#�==>�9>W
�>kI�>�c��ހ��5/C�қ��l>�+r>��?T>-^�>��"=�1m�G?�^�>�����	����c������Es?�u�?��"?���=K��I�+d��^��>��?g�?@{"?��^��x
>�]C�v�Ǿy�{�Ĥ�>�"�>~�>�@�=%��<h[�=���>���>�g	����.��\���a?8o9?�<�=ſ�(o�S�o�;���ߴ�W���.g�D���ؒW�gQ�=�����'�V��!�[��	������沾�N���Ҁ�[�>	��= n�=���=�B�<B4���O><�M5=�ɸ<t�=s%I�Mb<.�G��m��Uo��ψ����<��C=T��mx˾�w}?�)I?�+?�C?y>��>��2���>�|���M?��U>S�.y��`<�����&��dؾ�y׾��c����'#>��I�%d>��2>��=��<�t�=�r=�]�=��v���=*D�=S��=9��=��=�*>��>7w?7���ک��S.Q���罖�:?eG�>�,�=�ƾ�@?w>>�1�������~�?���?3>�?g�?�j��Q�>dᢾ���/6�=�ҝ�P�1>5�=R2�4��>�*K>���V��*���x<�?��@�??l䋿K�Ͽdm/>$,]>Y�Q>��_��-�ދ�+�y��p�Z57?M�;���W���>�g��׫�f�W�^L>�Pӽ���=�ă�6�D��<8>�~2�G����m��P�>�o�>���>Q�O�����
B=�����>�-,=�������i�D�1��W>>�>��>(�?]�P?�q?T��>������L�u�2>��Z>�9j>j�F>k7�>���>(^S?�n_?d�N?",�>"UM>�w�>��>7�`��F��`|ؾ/fǾ#W��]�?o��?#��>��J�?I��կ[���S��5#��$?��5?��O?bIP=�P �?�E#���N�mQ̽����|?>_a��A�;�����C����m '=d�>�^�>b��>��>oI>�]l>?t�>T.>ڊ�=j�=,�J=�B�=�X�-�>��j�Ղ��r0=�u����>'�=c�1>�K=Y\���8ݽ
]Y<��>>�l�>(  >9K�>V\>�(��š=(K��2�J�r >��^��~B��:]�� e���?�v��͕o>x��=���3냿�@�>�19>��*>F�?��z?�>!O���N��Φ�ڝk���=` #>�^2>Iݓ�u�D��T�@�M��B��o��>+�>�4�>z�l>i�+�3<�>q�=v߾�3����>�2���`����p�u���A�����j�/ֿ��>?�v����=!C�?��I?bՎ?k��>�g���aѾ��4>��z��=k'��Sn����$?�'?�P�>�xᾲ8?��"ᾛ���H��>"�S��`�Nm����:��F"��Y�����>�Č�'��g7/�[��[퉿F
8�l�;�;��>��/?H:�?��9������C�+�
��?�;���>XY?((�>:�>��?gzͽ�K�Ҡ��S�9>�Kb?͈�?�Խ?�(�=q�,�C�����>�//?I$�?�w�?V��?�����?�V����\��,�;��F�e�M��uO�`*�=�U�>��>�3?���#��x���Wھ�}"�F��=��9>]��>���>W�L>Od��2��=�\�=sͱ=���>�,V>��>=�>��>P�2 �^�p?�>U��=P�P?���>��k>i�r�)�`>9���!�JRj�jr��?�����f>����݃�:�M�/a>�ҿm>�?��h>jɵ���G?���Pr=>o}�>�>;<�=���>^ݺ>-�=+?�>�?�I$>�?�9�>��Ҿ�s>"��`!��FC��AR���Ѿ��z>������%�������,SI�&`���K��i�4��J=��u�<��?����Yk���)�������?��>:'6?����=���{U>�>l��>�����z�������s��+�??��?p\[>F�>�	u?�-?�8.��)��O�����0#$����XWP�8���%�\���(���W<ƪ�?�d?��4?/�>c��>�P�?gK@��r���[�>�~^��48��$<���>����z<
�{X��/�þܤ꽭r>�?"��?��8?�c�J���3Ǽ�;1?6�0?49�?#fX?�=o?�G����3?�� >�w�>�%?��?�L?(��>�W>'�=׼=x�j>y�b�?S������нF=�+O=�=�U�<J�ǻd�=)%=+˻G�n	V=5�=/s�<HX�<��=�U�=���>��p?ZS%?<`�>�e?}{���(���l?�^%?Ě�X�.���re��$�=F_�?���?c��?LQ?�>�n�I�x�=T�>��l>3&a>�u<>5&��`��p��H�=��= W>˄�>@�����-��_O�}нK��=��>�X|>�慽��.>v��-�t���f>�P��ָ�sQ��F���2���|�<'�>E�H?��?iA�=�_��,����e�8�%?�=?7M?B�?���=/�ܾ�9��cI�����6�>d�<�}��f���
���R9�
j<��q>���� ;/��q>�>�Rh��Ԯ]��1�����=x������=ߘ�	��{���>kX"�_-r�PN�x��������3?�`�=L�N�����YVؾ�l>��>�+�>���$��=u�c�8ɾ��T=���>Z"�>�}����gFH���꾬��>��<?Ttd?0x�?J80�{�g��RL�s8��J��������=?G�>�?�'M>��*>�7��D��*W��=�d��>��>e�'���W�������ω��v�>���>K�=�~�>y�M?��
?�9v?��5?�'�>�>Z>�|�j�¾.)?�K�?E�G=%a̽�&�%C�)>����>N
+?P��f��>0�?���>��)?��R?b�?��I>�iվ�65����>eU�>��d�1���	�>��H?[��>��P?���?��/>�5�-���O!�?hE=��3=6x=?�!?��?���>}n�>�զ��M�=�>�(d?�?g�p?�;�=վ?3,>��>|�=��>�G�>c?�cM?��q?:�I?_��>�D�<0ˮ��Y��d�x�l�P�X?�;_�<'�j=?�VNb�x}
��=��(<�~ļ#�"�ټ��6��u�|�:y��>��o>��ľ33�=�A��;h��"�5>R߇=�[��B#���S=��2�|WC>+��>��3>��i�l�����>Ϸ>�x�8Y?�m?��E?��ֽ��a��#��.`���>� ,?�2�>����ӄw���g�'>�a?�W?z��<�
���b?��]?o6���<��þ�b�"��O?�
?~�G��8�>�~?��q?��>vg��m����{�b�([l�R�=���>x�� e����>��7?Ws�>˅b>TI�=�7۾#x��$��"?2��?��?T�?AL)>i�n�=��}���J���^?���>!���#?������Ͼq<�������a������]1��y����$��[׽���=��?Y	s?�Uq?{�_?Ȱ ���c��*^����bV���� ���E�$E�ۉC��n�K]�&$��&��QOH=
���k�e�W��?}>?�"��t)?H=���(��nY���>6�$��-�`d�>�]u�T;F�$>�U��T���r��D�?M�?��<>��W?�2�N�S�j2�]q�IY���!�>��>� �>WL?�Kֽ��>��%>>�����/>�4 > �v>�c?�?K?=Vo?h����0�e����|!��=(�#��	�D>�>��>�
U�$�	�%�j�=�(�r����򏾢�	�v��=��2?9�>�4�>��?o?U5	�	����x��1�<�u<H�>"�h?:;�>7��>Z�ؽ|%!����>��l?��>�>򘌾SV!�-�{���ʽ�'�>�ݭ>#��>��o>�,��\��g�����I9�d\�=l�h?t���!�`���>�R?�{z:.�F<�k�>�+v�n�!�����'�(�>�t?��=��;> |ž����{�=���)?�?����]|)���v>t!?���>_��>+��?#L�>򥿾�컟P?pl]?�vI?@?�H�>�}=�g���ƽ_b&�cm)="��> \>��d=�2�=����Z�bv ��'D=�=_�Ҽ�O�� <�w����K<8�=)*0>o��CP��z���}�xk����iUq�H����_��Vz���оWܾ ៾��O4E�>=���ʓ�ߗ��@I��n3�?�!@��F�3��X���&��B�H���>@kֽ�ּ=v6�m���پtW��J�`��쾇�,��X�� ��S�'?(���T�ǿܬ��nܾ`& ?D ?S�y?s���"���8� � >�/�<}L�����G���q�ο����:�^?U��>��G��U�>Q��>w�X>��q>���r����.�<8�?}{-?��>4'r���ɿ���6t�<��?��@%8E?���־�M�=e�>���>t8q>��p����Ґ�i>S��?�q?�Ѕ= ���=w<C?��`���o����fH>V-I>R�ٽq9^��[>j��>�Dx��)�����4�6��>Jmg=�S(��.��F�c=���=�7���'�5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?X7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=o6�򉤻{���&V�}��=[��>c�>��,������O��I��T��=�`�D/Ͽ�����p=�{#=D�;'�˽v���s|���H���γ�p��=J�>&^7> #i>)=+>d.�>M�\?��~?���>�0�=�Kh�ǰ����Ͼw�0���������&�J�T;�}Ī�kݾ��Ǿ0%�[n&�� ��¾I����=�h5�����^E��∿��b�w� ?�j[>�;��%�*�C�����}_��:��=my��'���z��S�����? {:?���1E�l}�&ޤ����9a^?4J���T�-н'	>���=~�"�Q�>�q>T�����}E���/?��?�S⾀z{�!-Y>X1=�AN>�}?�N?��S�Px�>oM'?4����s�=Z�G=5P;;��\>��>�az>T����BV?�ch?p�*�-ˋ����>�O�I�����0<��>Ǡ���4=�=�>�'�4G��x��;?���7;�j�:?p7�>�::�������*o=l�;�v?jw�>����B?ɇ??σB�6���|�������#���/?;�K?I�3>�V����Q����,R?�E�?k�'?]z �s��]u��M¾1�?��I??�?"���lA��'���KtɾvK?��v?s^�xs�����N�V�e=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?m�;<��U��=�;?l\�> �O��>ƾ�z������7�q=�"�>���ev����R,�f�8?ݠ�?���>������&=�=�7����?��?�죾uE�<J����y��{�B��=i)W<�=���/l=>��y�/�o������h`����<a��>-�@�]��R�>Z�����ǿ	���׾�,�[/*?cX�>��I�$X����Q�unK��H���"��;���H>��2>�4�.*��3m��aDP��＾�?bF�l2A>QB��ﾙ���0�Ͱ�>p��>��>�k;=O
����?�&޾.�ƿ���9�ɾ�6�?�?Zƒ?��#>��s��\�t�X<��k>�,0?|fR?L"�>]OX�K�<n��>%i?���*�]�x�&���4��ct>p�=?���>�@!�?
��m-/>���>���=i��QHƿ�쵿�&���j�?���?^��2�>��?C:?����M��X���U2��^�W�>?ߗJ>ݷӾK ��N2��.��ɉ?�+?�e<��p�V�_?"�a�H�p���-���ƽ�ۡ>&�0��e\��N�����Xe����@y����?K^�?b�?���� #�`6%?"�>g����8Ǿ��<���>�(�>*N>�G_�X�u>����:�/i	>���?�~�?Oj?���� ����U>	�}?�ڶ>���?J�	>��?��>���펆=^�=S�>/K���?d�=?v|�>�H@>o�i��10���@�
>S�����D���~>s?#JU?)�S>-����n��N�#�I�Ž6ڽ��q�EE��\�ռv����J>�aJ>��,>~����#���?Mp�9�ؿ j��"p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>;�>�I�>D�Խ����\�����7>1�B?[��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�c��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?NQo���i�B>��?"������L��f?�
@u@a�^?*�:���ʿ�
Ǿ*Y۾��=�/>Ta>�"��v�;	Q=b~{��g���>!��>��Y>9A>��=�e>R_\>}i��֥$��n������8c@��y��j���ƾ�&=������ƾA����^ ���A�<�Tݽ�h�I���e�=��O?}�W?�[�?�	?�)v�gu>���I�=Z�!S>��,>p?"]]?2Z	?+|<�o���yl�/�q�$⳾W̓���>Y�=>���>��>�&�>b\���>�u>=}Z>Y��=�6=�g̽n](<8W>�j�>��>"5�>0;<>	�>�Ǵ�"#���h�	w���̽(��?Ԏ����J�d���C������i�=�l.?�g>����*пT쭿�3H?�����*�N�+�@�>g�0?0pW?#�>�M����T�7>
%�S~j��J>m���l��)��P>�?�Ow>��>}�&���2��bM�w���`�>��+?|"��>����G�H� �Ӿ�2T>�!�>I��<0�#�顜��փ���}�D�f="�B?�9�>Y�ҽ�K��.�z�5ɜ�j�S>��t>��X��r�<I=Q>֏l�y6�C�a�;<<<^��=�._>e�
?��H>(�R�pk�>�*߾��\�>�A>o@>�:?)$?�b;�"D��׽&;k��||>�Ҕ>C�=񾝼xJ潓�;�z�>��>��S�F -��z��e��<f|e>MUk;���MTf�į��W����<�c	>CUd<Te�X�P��~?���(䈿��e���lD?S+?] �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�Y�>�i�Z��f����u�PW#=�e�>:LH?�h��bQ�e�=�$m
??�U򾄙�� �ȿ�ev����>d��?��?%�m�a>���@�I��>՜�?�mY?؈i>�~۾m�Z��{�>��@?bR?�;�>�@��'���?I߶?{��?�I>d��?X�s?�l�>�9x��Z/�B6������=r=��[;�e�>�T>����fF��ד�"h����j�w����a>��$=��>ED�;3���5�=�����I��Z�f���>k-q>g�I>�U�>�� ?�a�>���>�u=%j��f‾G�����K?{��?:���,n��U�<���=�u^��?�<4?5�U��о�>(�\?���?��Z?�k�>����J���뿿(���~��<�9L>q)�>�0�>�c��%K> �Ծ�D���>R��>�� ھ�7��-����>�Q!?��>�;�=�� ?��#?�j>}(�>eaE��9��M�E���>&��>�H?�~?e�?{Թ�6Z3�4���桿�[�Q;N>	�x?V?�ɕ>D���̃���`E�\4I���R��?�sg?�T彾?32�?��??�A?�)f>��zؾ������>:�?��ǽ,�;�q��L��`?ͺ?�q�>ܱٽ(ռ�c<�� &��Q?�iM?K"?ݴ�%R�)�����=��A�2�<�<�Y=���VE>�+�=>Ss�0�>�,'>|��=@���7R��b
=�=�#�>�� >ڌ��sȽ�,?�`>��悾Gy�=�Ir�cD��~>�J>*h����^?�<�_i{�G���r���xT�a��?��?�J�?:���zh��<?��?�J?
.�>����޾&m��y�8�{�TW��o>���>�Q3��E�y���`v���I���ǽA���1�>H^�>:>?ֺ?�m>��>����,�������5_�$o��'��8�����梾�l\���*<�V;g���7כ>����"ڱ>�"?/k>�r>�K�>H��"IV>Q'4>�o~>q`>.�@>RSN>�F>���<��v��sQ?z+���4(�S�̧���yA?Ne?w��>Ia������ ��< ?�r�?�Ν?��]>ZYh�|�*�C�?�,�>h����?�G�=8W�<�v<{&���r��a�����=�>�!ǽ��:�:�H�+'b���?5�?)$z��վ۽8�����n=/N�?��(?��)��Q��o���W�qS����8h��j����$���p��쏿[^��%��ڡ(�-m*=��*?8�?������v!���&k�?�df>�>C$�>'�>�tI>.�	���1��^�L'�����mS�>,[{?�$�>aI?��<?��R?7�L?��>�>$j�����>���:l��>��>�O7?��.?�2.?��?��*?��[>$����o����׾t�?I|?��?[�?d�?�х�%wʽz���LUi��$|�D�v��#=@>�<�hٽK�p��D=|�N>	+�>��=��8��� ��'��n'�>5�>��>�6@�]������>�1�>p8�>t�[>�%n>Y0x��7ɾ4��>�#�>�L�77y=W6>�^�=�����˼�_q>�O���ST>�m0>��������� �=�>�� R>e:<�La =�m�>~�?���>�:�>���%� �-�����=�ZY>�:S>>>�2پV}���(����g�r�y>Lz�?�v�?T;g=M*�=A��=)|��([������佾)!�<��?�B#?�QT?���?;�=?$g#?��>%��K��EX�������?�)?�4�>`��+̾����;T��?oȻ>�OJ���<hnp��Lվ�L��7�.>j,�>Q����0��>r�V��Q�����?�#�?.��q��ܾ�#��iĉ��&>?@yr>��A=e��>��$���#�4�%�Q��=,k�>�RV?)�>ČI?ő�?ԟo?���>��3��y���g���ˆ�D��=��8?{1�?B��?�i?�_�>xn>�ai�6�ӾiZ�(����<D��ٝ]<�x[>D�>���>U��>�����f�w��]�����4>��>p5�>K�->_ۦ>��Y>������I?W�>�]������<��]Lr���&���t?�#�?k�1?�<H=w�%��fH�3�>�>sI�?٦?<?��_��>b��i����	o�F��>4G�>Z�>f��=f��<m�:>���>��>�-������>�4���?B?e�=��ſ�>q�ոp�h���N<�撾��d��A��$yZ�LU�=����<�t��D[�i����$��e����眾y�{���>
\�=~��=s�=my�<�>¼�<�]N=pϏ<�=�Cq��Sa<�;�p���@��[�޳o<��G=��)S˾{}?�I?֌+?>�C?��y>��>i�4���>�q��2B?ȵU>�MQ�bL���m;�Z�������ؾ�Y׾��c�����p>�_H�U�>�3>0��=I��<jE�=L�s=���=�a�!�=G��=��=r��=r
�=�>�>>�6w?X�������4Q��Z罥�:?�8�>b{�=��ƾq@?{�>>�2������yb��-?���?�T�?=�?Dti��d�>L���㎽�q�=Q����=2>s��=v�2�T��>��J>���K��A����4�?��@��??�ዿТϿ6a/>��T>w>��Z��I��� ����yо��P?*_/�e
�Ӻ�>�+�=�T�=��IR(>��B�;��C�>l�I����=~~�� ;�<��>x
>Q��>,`��E$��0�=�Ͻ&��>1�=�E�=%��b�5�̩A���>$��=聿>�G?ҀB?��?���>����v��ݾ�͇>f�>�9>�6>��>��A>�=?��Z?�Zp?� ?�φ>D�>�n
?w������9]E��&���=�R�?�1�?m~�>�4>��%�FՋ�����<Gy���?�C?�Z,?�t>|�������"��GI���V=p�=��)���<A��2������^j�=���>�L�>[�>�t�>��=G�`>��>J	B>+	�<�L�<w�<Z�h=TJ=�=pл�1>�mx=b����8$=�?:1> r�<�ϗ��{�f�F=�V>��>2[�=���>X>�=Yݳ��gB>�kn�v@�eL>՞���DW�efd��zM�ݶ[������>�+M=I�f��l���D�>�,j>pn�=���?  Y?%>H���Oq�Ġ�>��i�=6�2>�i�=�rc� �Q�;�h����j��> ��>g�>���>���-�-�Ժ>��R#�t�>.i��F׼S\D���K�b{���ݝ�]�d�zͼZG?V\��32�=^��?<�Y?qX�?L��>��ʽO�t~*>��K�W=e�!�x�N���ý$�?�@&?+��>���+>I��QѾV���s��>ܿD�3R�q����2�>�u��ޯ���>O���gzվ^�2�E��꜌��C=�Fln����>JF?�&�?E~O�U��u9L��+�������>��f?C��>�o?t?u%���s�
d���_�=vcp?�R�?~�?A>ͣ���߾��>�?:��?w��?e_�?um侅��>h�ƽvo�=�;-+�>'ݡ>?s��<RT�>��>�Q?�R\�J����Q�� T��w�{Ã=ǁ<���>D�$>!�U>Ȥ��P�=�dG>�i:�-#>B�H>��>�>�>]��>ځ�����v�?�|�=v�P>�Y??h�>@�<얽 �>�� ��4w���ѽqL���-�=&+Ⱦ��¾�/�_�D>��ӿ��?��>����b?,����>vq>wʄ��8>�j�>�h>��=v)c=���>CB�=���>�>�Ҿ�>:��3�!�eD��JR�p>Ծ�>�	��R�'����_����G�����N����i�xM��[�;�D/�<.�?� �K�k�uG*����U�	?*c�>�6?�Տ�4����5>tU�>��>����p'��R捿x����?���?ۋ_>��>��Y?T_?O;)���D��Y��w�5�<��/]�9~_�%���G�|�.L��򹽭d?Atx?��A?R�=�sy>�g�?8>)��|��Gʓ>Z2���:��V=�ԩ>Jذ��0M��iо��̾���[�H>�#o?���?D�?�CO��h��{��=A�2?��+?Z�z?ӳC?�;D?z�-���$?(: >cr�>�?�???$?���>�>c��=����=	�k�񰄾ꀼ�1d��\a#��'�=��U=^���X'���Y�<��+<䑻ȟ�����M�Ż���<�K�=r�=Nw�=���>��?�e?wÒ>�ֈ?>�ɾ˚���(3�&˚?�?������P>��!�'���p!<V��?�W�?A�E?k�>���u�d��S\>�r�>�2=�1�>� �=�٫�G=���~��A�>�/�>�+>Ѳ�=n2�2b/����w��Ʃd�P��>��w>Yψ�N0>�6���u�әi>�J��2����<�lH���6�Pa|����>�.C?��?�ׄ=L.�un����d���$?(R<?��I?��?��=�پ�<��J�$I'�߃�>5�=l��J��T��
8�?Oջs�c>@��Z��h �>��پY�+�d�.cb��H���,G�ۻ!�"�>@3��'E˾S��P��=1�=���J�]r���{ȿ��=?f�3>�9��A�/�	��};=-�q>�>I��=p����.��-O�ۡ�=*7?��>�#>�,��%=�]n�?��>��B?�vZ?�|�?!]����t�?A�����c��R�N��U?�K�>ߊ?0�:>!��=���F_�08`�0)H�^k�>��>K��egD��<���?�ô$����>;?7�>��
?�XJ?pX?�_?�+?��?���>���������#?�'�?]�e=�)ҽ��b�N;��C� �>z
+?ʂ:��B�>��?�S?�%?RS?��?��>���bB�[p�>l|�>��X��᯿)DM>l�J?�ȹ>�Z?��?��%>60�{���泽Y��=�>=�-?!"?6Z?���>t��>�������=h��>��b?f0�?��o?���=
�?�:2>^��>���=|ğ>y�>
�?;O?��s?�J?<��>�Ɏ<"1��Wn��Hus��	J�֔�;��H<[�z=���Ys��^�%��<��;���_\���:�B�D��!�����;Xe�>k~o>f0ξ��n�2��؊��C�>$5�=�3��㰾T=�)v��?���>O��<�Aʽ0�=� �>^<�>Gl�=��> �<?8L?�x�a�u��j�rY���o?��c?''�>��O��h��8�q��E��!��?�A/?ҹQ��-.�d�b?��]?8h�]=�v�þ#�b�3��d�O?(�
?�G���>��~?��q?��>��e�y9n����Db���j��Ҷ=r�>AX���d�FA�>�7?$N�>�b>� �=�t۾��w�up���?��?�?R��?�**>��n�[4࿣[���>��.^?���>V���
#?�����Ͼ�<������ᾆ����:��Ԕ��n�$������׽�ͻ=�?��r?<q?N�_?uw ���c��$^�X���zV�$)���_�E��E���C�ͮn�rd�nM��O"���(H=��\�Z�n��&�?[�?n�����<?%
f�ۖ��N���!��>�x��Z��@���%����'>��_>{� ������o���
?3�?6�>Sd_?Z�F�&�B���$�S�Y���ﾪE>��>�p�>�H�>�-���[��t8�����Z+�-C˽�w>��b?�1L?co?j����/�A(��{"��.������B><8>�F�>0�V��f�ك%���<�Ir����;���-
�v҅=�73?5�>,��>���?�?zL	������{�:J1��-�<�8�>��h?+n�>t�>c׽D���w�>׈j?��>&��>����*k�[d}��|��:�>E�>���>j��>i*=��d]����h�"w-�R��=-�j?5*��e����d�>�]^?�a�<;g=c��>�ҽq�!��o��E����=&�
?�:>�p:>��ξ�%�P���Ѐ�cJ)?�7?���L�*�j�~>�!?�[�>�c�>+�?��>þ���"?�]^?�J?�FA?��>|� =D:����ƽ�#&��B%=y��>��Z>��r=��=K���]� M!�X�F=��=�YǼ�鵽�m�;������6<p�<ۮ3>�:ٿ�d@��\ž7#����*%��_��Wmm��i��d��0h�������w��^8��+�V3������]�r���f��?Xx�?Im�����K��ۊ�
گ����>q���	ւ�����\蜽�rս�4���"V��+i;���[���{�ʓ'?B�����ǿ밡��<ܾ�  ?�@ ?#�y?����"��8�#� >�m�<�ܜ�ߚ�e���s�ο���o�^?���>m�3��4��>���>i�X>�Fq>���G��<g�?�-?ߢ�>Ӂr�֔ɿ6���i��<���?3�@��B?�3$��c�N�a=��>>�?�Z>�����!�����>x��??�=�T��g𼥋`?��ͻw|D�e̹��=^�==ʭϽf�A>n��>[��}�L��|ͽ)�)>�X�>e�D�����f�z�<�^>8�ν3�ܽ5Մ?,{\��f���/��T��U>��T? +�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?$�(?:ۿ��ؚ>��ܾ��M?_D6?���>�d&��t���=w6�8���z���&V����=[��>a�>,������O��I��Y��=��-���g#��U��*<C	����=��0����4�2�(�¾�o��g��zG�ג"��H�)���iv>���>^�Y?�Qa?��>-�>L㛾[��TǾ�=4��Q"�GP1>S:5���l���q���?��K�����������r�v��8<�?��=sO�h����3#��f��3D��X'?�Q">�þ�G�B<��Ⱦ�>�����:���K���~�,���p���?P�D?����g�R����q=��?����V? s�`��v��S��=!�����i=<ا>`.�=��پX>.�15R���;?�� ?��������{�>�I<f	�=_"'?�'?|�(�I��>�?P�̾1fm=�>�=
S:>��>E�?0�n=S�Ⱦ�C��/?�(i?�l(���Y�#%�>�о��^���z���n>I��Y�=� �>EDþ��Ѿ�h6��i�N,���*?=�>�3���!�Ց��
��<�z8>܉r?��]>��5�_�J?���>���=awս��[�쾩�(>��/?�� ?��L>n[�&����Ѿl��?��X?	��>k�=����JU��A;��T?7��?��5?��H��P������e턾pO?��v?�r^�us�����O�V�r=�>\�>���>��9��k�>�>?�#��G������yY4� Þ?��@y��?*�;<��U��=�;?i\�>��O��>ƾQ{������	�q=�"�>����ev����$R,�X�8?ڠ�?���>(���̩��^�=tԸ���?m��?LɎ�qb#>M��yp^�J��Mt1>}���'���>������g�"���t�/-���̾k�K�>��@��½a��>��k�~���ʿ(ʖ����F�^�t2/? C�>�켺ʫ��f�y^�Zﾱ%�oT��!xI>��>�W{�2{�GӘ�I�?��9���i�>�J��@>�gK��?��!�T�� >��>L�>BU�>U�=�j�p��?�������zQ��$ ����?Ed?Ib�?�ӳ>�m�1�X=ģ߾9�f<��$?�t6?g�?Ţ,=����>eJj?/g���7`��4�E���T>�G3?��>&�-�v�o=��>�0�>�>��-��iĿ慶�ٴ��_��?W7�?K�$��>�c�?��+?���2��<P��hk*�ē�:a�@?�U4>��þ�(!�1+=�ؓ���?,�0?��s��_?|�a�&�p���-�r�ƽ�:�>��0���[������+�,se��	���Yy�k�?_U�?��?A�#�,%?�į>�ƕ�YEǾ ��<P��>^D�>�N>�_�Asu>A��R�:���	>��?�b�?�c?]����2O>��}?��>��q?$�3>�?Sd�>cG���{����=+�>`Z���?/t??�>+wk>8���1� ��R�b%5���"��mG�UYY>ݸ�?��e?��3>H�$v�'����ӽ�����'���M�O�=�SJ��>o�>�>I���U	D? ��tA׿�T���*,�Z1?�p�>8� ?_D ���m��D�q�_?�4�>b�򀴿�*���I�T�?���?��?�4־I�ּ9�>?�>Je�>ӋϽ󢤽[��ބ3>�@?d(�ؒ����n�o܄>4��?R�@�r�?�k��	?���P��Va~����7�^��=��7?�0�!�z>���>��=�nv�޻��Y�s����>�B�?�{�?��>!�l?��o�O�B���1=7M�>͜k?�s?�Qo���g�B>��?"������L��f?�
@u@`�^?*ݚ��2�������¾�:�=��}=,�&>�+콒0{=j$,���e�X
����=�-�>�Tl>�>��>��R><�:>�(��~�%��^��n9��hz;�V;#����oh?��V�ZԘ�l� �T���+�ݾA��8E��MR�S�d���۽��$��>`�G?�OZ?=�?�W?�ӣ�7a%>q@�8��=�25��o=̹�>$#?�VB?��?�@<=�P���_��I������$���<�>@M=>��>�>p�>m;��^	>X�7>r�G>���= ��<��i���7=!|'><x>�K�>���>�B<>h�>-δ�P0����h���v��!̽�?����b�J�-���>�������~�=/c.?�~>����8пh�H2H?���o+���+��>��0?�^W?w�>�!��FWU�M>����j�i>�4 � �l�/�)�U0Q>�o?�r}>-K~>�!,��1��TL�����h��>4[1?�˼����!�y��0L�u�Ӿ�;:>�S�>^P�<f�"�0���J����w��~�=%@?�>�2㽕u����s��橾�%d>r�D>����b�=~�6>��yyý>�0�.�Լ,AN=�nd>]��>��B>Q� =!N�>x�྆jH�+.�>1P>=��<�/%?+�C?�_ƾ@��=�;��nL�{��>hk�>I�x=�V��������>\��>H�=>y���p�=�(��n�O��qq>�B>v��2#�s�B�܎����U>�-��E	��~J���~?���*䈿��'e���lD?\+?g�=!�F<��"�1 ��BH��6�?n�@�l�?��	�ѢV�:�?�@�?
�����=�|�>׫>7ξ��L�߱?��Ž�Ǣ�̔	�O)#�oS�?��?�/�Qʋ�Gl�6>�^%?�Ӿh�>h�mY��B��y�u��$=���><<H?_����O�~�=��o
??QP򾲣��-�ȿ�rv�+��>A�?O�?��m�@��|@� ��>$��?�bY?�i>�~۾tZ�2��>C�@?[R?p�>�7��'��?3ܶ?\��?V�H>��?��s?�k�>�x��^/��0�������=&�_;sc�>�]>)���`F��Г��`���j�����a>��$=��>��9)��xJ�=�勽P��C�f�!��>�5q>��I>O�>�� ?Lb�>���>l�=�A��r܀��Ζ���K?�?A��8/n�W�<���=Ś^�N)?B4?��Z�^�Ͼ�Ϩ>L�\?���?��Z?�c�>���<���濿�y��K��<�K>T0�>RS�>�5���3K>o�Ծ�7D�4s�>�˗>nU���Eھ03��Z����A�>�e!?V��>��=H� ?K�#?�j>�&�>�`E�t8����E����>K��>5F?�~? �?�й�VW3�����塿_�[��;N>��x?�U?�ɕ>A���6���N�D�O,I��㒽���?fmg?�X彊?J2�?�??x�A?%f>u��8ؾ����]�> �'?�ｓ}=��o�h�"���?*�?do�>����(T��3�< ����ƾD��>��H?�{ ?[�����\��˾��=�-û�z����L<��=.��=b��=U'&�$f=gB2>�=v�~��gd��q�ȽU=�ǐ>m�=ykI�.�7��=,?�F��Ѓ���=)�r��qD�P�>:=L>����M�^?�Y=���{�����x��KU� ��?���?�f�?����h�a=?�??�$�>	@���~޾��$Qw�Ґx��{���>���>Vj��
徦���镪�eI���ƽA�Ž���>�5�>��-?�/%?�>�/�>�+¾I�������O��hB�� ���&���2���ՓѾ5;]��}ͽ̽ľ�a��B�e>4뽉9�>� ?��>oP>��>���R�#>�&�=�8V>��`>�[�=�(�=���=�o=�dR=�)O?`D���)��,�׺���z??��b?N��>8��������e?CA�?��?ʐk>(g�?5)���?	� ?�R~�w�?j�g=�r�;�:�*�����>���r<ۼ�K�>�Mƽ�?���G�%t�c�?B�?��&��ʾ��˽�2ܾw��I�w?U�?�1�ΖN��g��*T�>7=����:@c���.���{"�6�l�麏��@��D��i����>�*?�#�?o�����;�����n�=F�׿o>*��>�>�R�>˒�>������M^��:���m�GR�>M�w?V��>��2?9�Y?�*z?=�O?८>��I>[���5?�yFx>��
?Қ?^?g?�~�>��#?���=���H`�~ ��?#�3?Ld%?�n?��>G۬�"}�T����Г<�s=��>u�=��9�b̽5�󽙡Q>���>��@>�$X�\5L���>=z�>�u�>�L2?�-�9�"FĽxy�>��G?K?р��#�]�ս��?'�2?wX$�ɪ �� ->v{@=k�P�C���ŇX=��}?�=���=��Խp�>�������2>����HQ3�M��>�d�>��?�>�2�>�:���� �������=VY>S>�/>?Rپ�z��}����g��y>v�?4k�?�f=�`�=���=Ƒ��eY��,�� ����:�<L�?��"?�T?Vp�?�=?ā#?X�>P'��S��R�����?�
0?K�>�v��Y���������b�?�>��Q�.+S�{Q~��<뾶�ؽ/��=�7�Mh(����*㜿u���&�6�L��}�?�݉?ri��2��(�$��ǈ���L�
�?�,>�c�>04�>���� !D����勼�t�>��^?>p�>iA? х?��}?��>A��N����J��J4=���=��?c5�?���?R�h?�V�>�R�=������R���?�#�(N�㨇��^�=��`>vhp>�n�>J1�>���<F.>���ݽ�{��u�=��]>B��>�ߣ>�ʮ>��?>�s���iE?4?,UȾ���(Xw�� ���l��:�U?���?Y<?�6�=�����{� ���?^��?:m�?��?��I��'>�(�=���'�پ	b�>)�>UA�>��A>�'Z=��P���>�f�>sһ�����#4��:��G�>v=?��(>g�޿������y�%����)��sܾ����4Q���"�ŉs>���7f/�3Y������Q�u-����]H��%=��?	�>�� >Rk�<�)������/�����<�=4>JJ�<����]�<�¼��=��<!�=��.>'��=L�!� б��*q?I�Q?�(=?��L?/��>�9=><���)�>��w�ڰ?�[B>W;d������a�|���;���b�پ=��XQW�4��.>J���3>վ]>>3��;ֱ�<(L�=~i=��;=�=v�'=���=�ȥ=���<f��=��>�6w?���ײ��14Q�VY罏�:?*9�>~�=R�ƾ�@?��>>�2��g����b�;-?A��?�T�?U�?!wi�?d�>����ߎ��r�=����<2>@��=��2�m��>c�J>���J��t���{4�?b�@��??�ዿ�Ͽ3_/>��5>�?9>�ac�[L�[O�����s���K�A?�g��8	���><���%4�S"	�j$>��=|�=��=i$(�A?x=�_#�0@���Լߖ�>�
>�l�=�������HѼ=�=dj>�$�<�0�8��<;���s-���5>�n>:��>P�?5 ??��o?-x�>/:��T.�C��	*�>ю�>�,�>t��>�J]�x���;0z?**Y?��h?�Q�>$��;���>!��>.��}\���s'��R����o�?pge?B�?�	�>:<��c刿s�>���i>Kj4?��R?�+?�L����8.��_%���-���x�{W���4=�kl��_�7'��kH�:��Q��=��>d2�>��w>J�U>l
J>��Y>��>0��=��<Lw�=)=��� �9�%c=�Ǧ=���I��<$�tAe=Zy�ű��ӗ�i?����a�<�/=��=dW�>�&>L��>�˘=����7q">s�����F�|@�=И��M�<�j�a��Mz�*,��1��~N>TVQ>�j�o㏿)��>i�W>0�R>��?6�t?�>թ���ݾ5���)xx�ւJ����=�� >��9��Z=���[�f=P�n)˾-r�>���>�>�z>��'�37��J=���2�S��>�貾\�P�ؒ��i�ǻ��擘�
�q��Eý 7?���"v#=܁?FG?�
�?�/�>�%��4¾�_>>|�}��k=�z���m�d-����?�l?�2�>.�¾j�:����'����>#�s�{�P��ϕ�X2��)�@~�����>����`��,��"���I���W�3����z�>.�V?��?��M��1w�r�C��*
�̃��L�>i�X?Ϩ�>�>g��>��s�q���y��:w=up?�
�?�Ϲ?�!J=WǤ=K������>/K+?F��?�?���?�ţ����>�eA��,�����c�E>���=�<��]��dN>�l�>��?�D�R� ��h!�	��Y`��P��>���>�ku>��>�j>>K>�>i>N�>C��>��>o�s>�F�>���>��E�ۖ8��Ut?��=�h>��k?@q}=��>����fl>�� ���H r�D����$�;pc">s��(�ʾN�+�<m>�5ؿ��y?�S9=�W��7S?y˝�4�}>���>��>(��:�7>�j�=	_>��?�n�>\�>�?���>�پ��>tp�38"��6D��QQ�c>Ѿ��u>H����I!��l�[l򽘡I�ۡ������k�M�����:���=ޱ�?I]�e$i�ֺ)��2��s?���>�%6?�������{>|n�>]͎>�������y���ia߾ǹ�?W��?�g>�i�>�*o?��+?����9	���U�/A��B��'�C}K��L|��9h�!����Ϡk?��Z?��&?e'��Ҏ>�8�?��6����r�>�X���P��i��n��>����Ȼ��ɖ�&q侢�-�܂�>�b?�?��T?����%�����;�N+?��<?G/�?�^E?�k?�V���!?T�+>z��>�?��1?9c)? ��>#��=��<5ݥ����=ϐ=�Qч�E����
��� ����=�p�==9$=Π`�H�>V���J6*�F�]��.�����<k,�ә[<a�=�n?>���>��v?T�&?IT>=>?��Ⱦ�.��ʘž!|�?��?�q>���>�A���u�*��>�Sx?e��?�a@?I��>���}���S>��k>g��� �>.��>�09�L��p�e�I� �>e�>)˿=�|�����:��,��>wW�>&|>�ۉ�r�(>�b���Uv���f>�4Q���(jQ��G��1�u�s��%�><�I?pl?�}�=���ś�הe��'?{z<?+�L?��?�C�=��ݾ'*8�nJ��I_�>]��<�������R��é:�Y�);�	v>�㟾���(�I>���ٵ��X^�,�S�{��o��=�{��| �= ��]������"��=L?_>9ߠ�7k���������D?81>ŕ��O�����S��=���>��>�_�=Ԯ-���S��6����=A��>:3�>7C�<���bS�$���x>�2?Q�I?�X�?��5�mn���V�r���ײ����;�n?���>}?(>�v�=���E���^�.p7�G�>?�>��K<���˾�%���>�(?�\�=r&�>�7M?�?��\?�4?�"�>:�_>N/`���׾@?�C{?u��<{�"��s=��D���>Gr(?��=�z�D>��?�c(?"�?@�[?S;?P��=o�0SE��ߚ>,T�>�;R�6F���^�=��??��>�Y?J|z?|��=4O9�ᗬ���p[�=�R>�2?�?A�?Kp�>��>����he�>��?D�v?7�?6G?����ؠ?oP�>�Y�>W�=)&�>��>@?�GX?�$�?
V?~��>l��;e�,���T�����;x�-=���<Х�=��2&=�Z�<�u�<ʢ+�����L����<�26=5U=�V�>�Ht>�����0>�nž[����B>
M��!雾F��O�;�C��=�ހ>�F?Z�>�#��=���>"��>��	�'?�?�?'�o;�bb��Q۾�L��P�>oB?�v�=U�l�~���*v��i=s�m?�H^?6�W�����a?(�]?��@�9������e�`Nﾾ�L?σ?��L��m�>��?��r?�0�>�e�A�i�|����a�ǫg�R��=7"�>�"�I�e����>T�5?���>>`g>��=a�ܾ�Cz�a����?��?�9�?�Ǌ?ۼ)>zn��D῅0��$/����]?���>q����#?��S�ϾA?������ ������q��;\��#���l%��ꃾ�*ֽB�=P�?��r?�]q?ǿ_?ɠ �B�c��S^�6���}V��+�X��w[E���D��zC�~�n��k��&��c���h�J=e�h���;�Ge�?x�&?��:��>�Y��e���
���nw>Cl��!��s@�<bI���C<c~�<g~�������^W?���>�'�>~f>?�[��D�@5��,���$N�=%��>���>�#�>�:�<I���e ��ľ�앾6I��Ȱ�>�gb??�J?U�k?�D��3.��#����!�F��<6帾P�C>
P>���>�[�c�����2>��~q�'*�$i���O�vP�=d�%?��U>�E�>�˕?���>�8 ������X��?l;���L��>&k?�S�>B��>�l�0��9�>�2g?���>�%�>�҃��֗w�����v�>���>�L?�Qr>��H��>[�1����荿�`9�,:>{�j?�u}�X{T����>
�S?�90�p2:����> �|�T%&�������+�ߌ+>��?�Ҵ=�D>O�þ�
��{��낾�Q*?�?�Ϥ�C�"��j>���>�?|<�>D�{?"�C>�R ��8���?�JY?H�Q?��8?�h�>$���;�"�����'�&�8�@�2�>,�^>��=��:>P&%���]������<{��=��� �<B<d1ؼ��E=
r=ү	>�MԿF�`�Lg澞�޾��	���+P� �G�n�k���Z�H�d�ξ\�������P�<�F�2~��ܹ��Kx�Dn�?��?�,|���-�Y]��д��n!����>�V�KkI<pH�ܼ��V�����nGH����v'�KY�d��-?��d�����&���ھ��?��
?��v?ؗ#�L7�l��Uk>3�=N��`]��+��P�ֿ����Hg?��>��ܾw����>7lr>]�@>�H>�1~�N��˟P=��?�f4?�>٘x���̿�?���p���E�?��@|A?}�(���FV=E��>Ό	?��?>�A1��D������K�>�:�?��?Q�M=��W�=�	�Gze?+�<j�F�xMݻj1�=bA�=�X=���ڗJ>�T�>:���MA��-ܽ�4>�څ>�"�����}^�
G�<ǌ]>��ս,��5Մ?'{\��f���/��T���T>��T?+�>\:�=��,?[7H�_}Ͽ�\��*a?�0�?���?$�(?<ۿ��ؚ>��ܾ��M?^D6?���>�d&��t�݅�=�6�#���w���&V�n��=W��>^�>,�ދ���O��I��`��=�� ��e˿)�"��'��2=ܻm���P������V��肾J���7uW��ߤ=��=��>>�C�>��|>��O>.tZ?V�q?ɏ�>Ww>��9�	x���|��q,�=��O���׽��<��5��,��m
׾/&���x�v��zm�v�־�4��K��A?I�L����A�������#w@?�^��"���/�h	���Ǿ��2��U%>��Խ�TȾ��-���q��͛?�V@?tҐ��ш�n�����<2>џ�?��:�ˮ'�[�5>aB�=Cr�>��>�M�=;��bq�_w[���0?��?�Z��������$>��j	/=�@,?b_?FM<�)�>�$?�].�u��.`>�+5>�u�>��>�>/����rֽ�E?S?�C��]0�����>+���~�_�k=վ
>4H8�p��#Z>���<<鋾fA��׉�S��<h�W??�>{�'�9f�:���m�v=M=x?���>(0�>r#l?ͰD?gH�<Vm���S����D�=�P[?9�j?��>E�y��Iξ�ߩ��4?|&c?��H>�f�)�꾝�+�o��_>?fm?�2?���b��� �v\8?��v?Jr^��r�����,�V��=�>�Z�>��>!�9�Zm�>g�>?#��G��)���NZ4��?��@r��?�	<<i&�K��=�;?k]�>��O�i=ƾ�v��������q=�!�>�����ev�4��O,��8?䠃?���>_���ĩ�m�>�l�bC�?lk�?�:J���	>���dBu�
6;{��<��X>�9K>�L�f �v=�R�Ҿ�/�?q���<>��o>�$@��ɽ[� ?�睽iT�e�ԿS�e�XǾ���=^?۟?�һ=.΁���F��n4���/�/`��l��¨�>��>L���h��-x|��c=��q��h��>\�����>�kW�0ݳ�����3v�<�~�>���>'\�>½V���Ֆ�?ֆ��oCοʉ��S��k�V?�Ɵ?(i�?!�?K���k����v���H?ds??*Z?5 O���k�zT_�bt?ժ��,���B��� ���s>��>o��>ץ{��z�>(?�>��?'�)>�u�bҿ,�ݿp	��6�?�y�?�n�ū�>�$�?�+?�ݾҫm�<����$F���>maL?��M>]��	V�:�D�y���'?� �?`���-�[�_?(�a�P�p���-���ƽ�ۡ>��0��e\� N��(���Xe����@y����?L^�?g�?��� #�a6%?�>`����8Ǿf�<���>�(�>�)N>cH_���u>����:�i	>���?�~�?Mj?���������U>	�}?�&�>8�?{��=Yb�>A��=c𰾆/��W#>Yk�=�m?�ݜ?�M?
O�>�F�=��8��/��YF�<HR�%���C���>��a?m}L?n2b>8總0�1��!��oͽ�`1����Hu@���,��߽05>�=>�$>)�D�#Ӿ��?Mp�9�ؿ j��!p'��54?.��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�x�>���?
�@�ծ?ji�4	?���O���`~�˂���6���=�7?3���z>E��>g�=ov�t�����s����>�B�?�{�?���>]�l?��o��B���1=�L�>��k? t?R�p�󾲱B>��?������/K�Df?�
@uu@�^?���ݿ��������̷ ����=��a>�:>�{����=�J�=.��=W =Q����J>�S�=��>��>��<>`�L>_���s'�X:�����n�0�������K�Iyܾs���1
�Fڹ�9���@�Ӻ�6���.�w�L��L��ߒ���>�<U?8pR?�Tj?��	?r�U��N3=�
�K�>��k�ng=,`�>�y*?�X:?� ?��>����<Xb�<�z�Ǧ���������>�z]>[��>� ?t��>�>����>R�m>�|�>+"(=~�7<�D�<���<on:>b{�>��>� �>I3>y��=˷��PƿH���~��/�>i�?n�ݾ:2���j���
�'<����>��=?��>�O����˿=:����5?L
?�_�5�Z�K���#>i�$?[�A?�|=>�:�|��Lb��1�{�򽌃t>�'{�����}� |a>���>nH�>i�>T�X���6��}o�ĉ� !�>��X?�C�;�ᾱ����&�����>�/�>f��<�
��Ռ�u������	L>[�!?S�!?1��6\7�*3�ӯ�����>��>���=��=�ͳ>@�->����T��!^�>B�O>G�>��?�%>k2�=o�>�Y��`MG�'�>�6>Qg)>��@?�%?*��Α��o��D1��p>�C�>���>l	>)�D��W�=$y�>��d>n� �����9]�ə:��UQ>��~�q�`��8��ӆ=[U����=ߝ�=����FA�z�1=Ն~?[p��숿V�V����<D?i@?��=��J<��"����YH����?�@�a�?�~	�ʖV�i�?�$�?*ڝ�dH�=��>��>D*ξPXL�۫?��Ž�i��!x	���"�/F�?��?f�-������l�H�>bY%?KiӾ�Z�>,��K٘����Uyu��&=��>�:H?����9sG�D�:��?h�?Z��h��Cɿ��w��d�>6��?�Ҕ?m�=���Jf@��j�>r��?�bX?��i>U�۾>�X�xю>r[A?��Q?3�>���M,��?��?�܅?%�X>,�?Kv?=W�>8l4=,6#�.Y��e����N�=
����>��>^˦�e�A�'���..{�:�i�� ��U�>Vh-=��>��P��tþ�69>5 1���þ���ti�>��@>�&W>?�>R>?}��>��>�c>/�����������T:?��?�D1�u;W��v��/k�r��=��&?�W-?��+����'�>�\?���?F_?�Yc>��پCҢ�����|9I��w�=<��>4�?��I`6>wϾ�����:�>G�>��b��؈־"�=?ҍ>A*�>��>��=w�%?�u$?��v>޵�>�e9�攀��]D����>p(f>� ?q?��?Kd��,�B��Ê��*���wo�N��>'\~?Uo&?��>�p��r��*ͽ!��#�'���?��B?1�����2?��?%�L?�? W�=�敾���q#>>��>d�%?�?w�d�>�o_��?{��η>��!?vY?}��<$�M�����Z�J���	?rCf?R?Kb̾�d���1,L=�M�<�]��IT=�����B�=2=>��+���=�v�=Gߘ=��M��
��Ok���3�=��h>v@�=�����@,?�=�F�����=��r�|:D�(�~>��K>�c���^?�6<�
�{��"��������V�Jȍ?���?�t�?�n��#�h�d=?��?n>?aE�>������ݾ���a�u��0y�ך�]�>�K�>4V����YZ��iv��y;��N�ƽ�罣�?.�>�?��?�,�>��>�������о`Q���Mu��t&� �F��hI��#��v���m#�N��=c˾{͍��RS>>�%�֧>(q�>�O>P&L>P�>޻ǽ���>�]>7i�>���>��>�g�>jw�;э���<�x\I?�Y����:��Cپ�z�?Hw?bv?�-F=O��������?=��? @�?�`�> �^�A~��)�>�5�>��`�	s?خ=�@�;C�<ՠ��_���=��ŝ>c�
��b#�<4M��쐾.5?M�?��?<��Ծ�}���ѐ����=9*�?�� ?ˈ!�FIB���h�7dN��YZ���#��m��e��p� �4�p�z_���9��oā��L�:��=�e,?E�?Q�������2%��{9k��gH��F�>]��>�,�>+t�>���>sF��N?��`�8�-�����	?z��?U�>�9?�2L?�D`?[na?���> ��=[x���?��l���>֌�>�Y=?1�	?��?!�0?&�+?��>�:νpr�����#?��?n�?�h?��?�]���Z���0>h�=m����Z=��= ��;v����נ=�pr>h@�>�X?���g�8������j>�v7?x��>���>���,�����<��>n�
?HP�>����Xr��d��W�>w��?�����=r�)>X�=����?�κ'S�=[A¼��=�j���;��P <#u�=�۔=[�z��O��'�:�$�;�c�<K�>��?��>L�>,l������g�RȮ=��V>��S> �>rLھS\������g�Nw>�/�?A<�?�l=��=��=��������	��۽�%f�<s�?��"?�#T?�}�?�O>?�q#?�� >�{�����W�����_,?��+?'�>����P̾Oᨿ5�3���?J ?]�`�R��E�)������.ɽwH>~.���}��򯿁QC���d����C��?��?��L�*�5�G���������)uC?���>���>�k�>	�'�y�g�/���@>~L�>JbR?�x�>s�O?8q?*[?��>t�)�Ț��� ����S>���e�@?,��?3j�?�zF?���>�ׇ>$�����������o�7ܽ�@��aJ½(j�=�}|>�C�>k$�>��A>Bw�����{ʻ�k�=8Ci>�?�A�>Re�>���= $���G?4m�>7���KL��T��3���X1�4�u?�g�?��*??�=WY���E�������>�9�?�̫?�y)?_�T�8�=�Ҽ:ൾ{tq�Ը>D��>8͘>�ԍ=Z;=.�>��>�L�>�q����;8��fK�c�?�
F?
�=%^��Yqj�$��0�?��gm���ܾ!͂��V�������	>�>�4>�"#���o�vp��hU��uL���f�6b��'��>4�>��Z>�G9=��Y��]�$���.�=1�˽��F�m�ǽv��=�MR=�+J<wZ�ƚ���Z��Ӽ��5�
�Ⱦ}�|?B�I?�_*?J�C?�Ҁ>�>WU����>C��.�?��G>�Eh�)E��!�D��5��.s��D�Ӿ�Ѿ�5d����L�>�Sj���>+�4>i��=1�;<�L�=��=@ܘ=�@X�/\.=�V�=N�=̞�=��=�>�i>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>^�9>0�
>d�Q��/�DJi���o�0O�ϐ"?�6��V;J�v>b��=ܞݾ�P����x=��=>&�i=�
&��?\��p�=��N��L=��X=�>3�@>��=8��؟=F�%=�?�=\-O>&칻q#��h7�*�%=��=��]>��(>ԍ�>)�?�]0?S[d?G�>��m�11Ͼ�B���U�>�S�=_;�>7�=ۼB>��>��7?�D?��K?h�>�{�=�>��>Õ,��m�f��	ç��Э<(��?�ˆ?h��>��K<�A����M>�O�Ľ�n?�@1??U?и�>�Z�ӂ���G���+�EM=%3>�m4�Q���+�=����B#���Ζ>��>m>c�>ďu>�/a>O��>F9>q֙�?W>�@:�Y���~�=�]�==Y��=�7Ś�z�ֽp�~����U�Ti�MƖ=]��=�Z�9>?H�>���>aj�>x��=y�B�^(�=����&�E��m>�PX�$}?���|�R�����`�3R�����>�O�>g0�=����5��>/k->���>	��?��?8�>#�%�2�b���\$������X>	�>��Q��o�<�m�J�L�(��Zy�>ޮ�>�o�>y�S>�!�z�'���2�8��{\@��?<i#�/in��L��M���~V��>h��5�5��V�=��T?	���R��=��{?�jX?SM�?�E�>%�<<ȱ���>����4X���D��4o[=�?�`-?���>��i�A��H̾����޷>�@I�2�O���O�0�W��(ͷ�?��>������оq$3��g�������B��Lr�a��>�O?��?":b��W��AUO���� )���q?�|g?"�>�J?�@?�%��z�r���v�=�n?ĳ�?M=�?M>K�=G�7�P�?z�>��?��?��F?�
��s?��)>��>ͱ_���9�	-���yP�h�=q/�>��?L9&?�9�<�%��ʾ3����7L�]{�=W��=G�,>E�>�,�>��>�/�>�kQ��a�>���>B�%>�ї=��d> ��>����mp	���?->�R�>��/?��]>TN�;(��j�n=ˑ�d[�;�8�5�-��q��<6���'�s=j�r�A
�>f���ǖ�?HZ>�x��	? ���m��!?>r�y>u֔��Q�>�E>�	]>-�>�:�>7��=�ې>�xJ>�ᶾm�0>���R���.���3��P¾��d>�}Ⱦ�Lڽ��ǋN�baW�E㽾��p�1�u��b*��H�=���?W�
��
R���+�K�:����>`�>>��A? ��V�;���J>g�?�ڤ>�6��V���T��1���?ri�?�;c>��>I�W?+�?ѐ1��3��uZ��u�(A��e���`��፿���(�
������_?��x?8yA?�^�<�8z>��?��%��ӏ��)�>�/��&;��@<=,�>�*��N�`���ӾR�þ�7��JF>��o?�$�?�X?pUV�J�=��5>��_?��p?J,�?.4G?<�?�i���q1?C��>���>���>b3?�?���>��>8ݷ>u�$>< �=�ļI�Y����(W��uh%��a<\< >1R;.��;Vy�=�
#=�c�;�� �z��<��:] �;��=Z{u>�#>Y��>YP]?Ow�>�9�>�8?�P�m8����w@/?OJ;=F���iǋ�7΢����&�=�zj?��?IZ?f	f>��A�Z8F��>��>�L&>��\>�>]���C��=�>k�>�1�=w�M�����	��̐����<Uc>.?�>�M�>O��0f>rdm�Z�u��̨>�m#���Q
�(>1�B=�h���!�>��H?�	?�>����l^�b�[��>�?g�#?茣?j��>$�A��5b���~���>�_?��E��i;󢠿���<#��[b���>�	J>;�Ҿ�2>R��a���O7a�ݫM�`ž��=Ca��-B8�q�����^���o>��+>��������$���"��T�I?�h�<�����4|�j+��H�c>ī�>3�>�-=��,��$<�h>޾1�*<`�?W�>���ƴ����*�rIǾ�ډ>��I?�.c?���?z�`�QJl��rI����S霾�ԋ�#M ?���>w�?(�D>#ƨ=Eh�����_���B��2�>��?4��ʐE��ơ�^o��'��>:3?*�>�?U?�?��_?��)?�?���>���kþNB&?b��?��=��Խ��T�%�8�PF����>�)?�B���>�?�?��&?�Q?´?p�>1� �]B@�2��>�Y�>"�W��b��_�_>#�J?���>�=Y?�Ӄ?M�=>��5�@碾�ө��Z�=L>�2?R3#?ű?��>h\�>�A��kl�<$�>8�U?J�x?��q?{�->��?/>�o�>�P<��>�L�>,�?�P?P�p?m�=?���>6��<"���vE��<�:������K�;�N�<_Oq=��;:�d��>����*=�#�;��`���;�Hܻj����@����<�X�>l�s>@��H�0>��ľ�N����@>�ᢼ�E���Ԋ���:�ݥ�=���>?���>�S#��=<��>OA�>��� 1(?��?�?�� ;��b���ھ��K�p�>kB?���=D�l����T�u��1h=W�m?ъ^?}�W��#��M�b?��]?6h��=� �þg�b����c�O?8�
?>�G���>��~?b�q?C��>�e�%:n�+���Cb���j�|Ѷ=kr�>TX�^�d�t?�>c�7?�N�>e�b>�$�=vu۾�w��q��n?��?�?���?�**>s�n�T4���t&��g\P?%S�>��]��(?�w;��!德�s�ۑ��^ݾ�Q���J��*��������Ƚd�G��`�$�=��
?��k?��o? 'R?Q0ʾ�R3�[�K��)m���N���о���7���O���C��~�7�R����P���&>��^�h�M���?�8?ڟ���n$?����i�lʰ���g>��P���%���s<1\ǽ��&;sJQ=U����ؚg���?��>�K�>�#?˲U�i<�z�8��0'��	�\�)>�Ȼ>�*�>���>@V=����	Q��ᾁ=$�c#� Gv>+Tc?V�K?So?����D�0��x����!��)�qɦ��)E>#
>C8�>��Y�s�z�%���=��hr�^e�tِ�x�	�حy=ò2?Ee�>(�>�c�?
?�m�%7��z�u�_�1��m�<K4�>��h?PZ�>���>z�н�� �~��>��l?���>�4�>h���F!���{���ʽ|6�>K�>���>�o>�u,��,\��j��|��9���=m�h?l�����`��ȅ>CR?���:X{I<e��>�)v���!�����g'�U�>�z?�9�=!�;>UFž��֟{��?����?��>�ä�c/"�HC>w@?8^	?C<�>��?���>�/־�x��^�>/�C?XL?uxI?˒�>�:���&������/��g�=�8�>��#>'�=���;DXy����DFH�w��;��?>#����[C�1�q<���p'��!=_�_>n�ѿ�TB��[Ǿa����ྗW���Չ���ʽ
�{�
F�鎻�����μ��5;4�m���.P�1[x��v��yM��?���?�G���[��±��m}���X��>Ues�<���
Ѩ��c�ݪf���Ⱦ����!#��^��Y��#]���N?�2�=����������?��?3�h?�H'�y�O�R���s�>cE�<!�'�K��k���v�L.->m�`?�P�>���t���e?�FI>3�=Q,�>�|Q���ξy�>���?�3?c�>Cټ���ڿU�ȿ�1x=F��?8� @y|A?��(�T��tKV=E��>.�	?*�?>;W1��F������Y�>�:�?+��?�=M=��W��	�`~e?�A<C�F�O>޻p
�=�5�='g=���&�J>X�>��JA�ABܽ
�4>�Յ>jy"������^�*��<�]>�ս4��$Մ?!{\�vf���/��T���T>��T?"+�>�;�=}�,?W7H�N}Ͽ��\��*a?�0�?��?�(?3ۿ��ؚ>x�ܾf�M?WD6?���>�d&� �t�e��=�<Ἤ�������&V����=U��>Ȅ>ɂ,�Ћ�чO�I����=���ƿ��"����(&=�"�;��d����Y���W�����K�l�����A�I=\��=�R>*��>nW>'�Y>��V?�l?�g�>��>B��o!��A�˾X�������������4�����ˑ�S-
�nn�����ľ�II��t�=��X�@���=�(���f�s_���,?��=�D��Z���輇�澜>i����<P"p�X�־(
0�>�a���t?:?{J����q�o�,�����t&��KW?rf�Ĉ�O�Ⱦ�Q�=Q����?>0@�>�	�P��XA�~SM��U0?�?P���:]���)>���=��+?��?$.W<���>�%?m+�׎� \>�4>�ۣ>_�>y�>]��5�۽Њ?yT?���Vݜ���>�����z�]�]=�>�3�l��t�Z>��<���u]�k���N~�<�`W?pؐ>�V)����菾����;=�4x?~*?0e�>�i?ȦB?3��<���)�R���
�F;J='�W?�Ch?��>s{�GJҾ]��IM4?0�c?^�P>�`�a�뾭�/�ΐ���?i�m??pa����}�gY����I6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������n�>��w�'?�?a:�?�����O><�9�y �����|�>펿>Z��=�Td<śƾkD&��j������F=��Z=p��>l�@i��E�>F�d��\�F�˿�������n[�Er?
?'�>\�2�oA6�x�E��3���B�����X�>��=�F���枾"mq���9���ϼo��>�7���>�hz���Ⱦ�N���
�=���>J�>��>��Խ1��_&�?ȿ����ǿ�v����y�X?�ա?��? �"?�&�<Ѝ��o��U���6O?�(l?
Q?>�D�[K/����Kބ?#&־�:(�E���7��$>��?�N�>#���"�=e%1>��5?N#>z9[�/wۿ
&׿���>�?�]�?�¼�@�>���?�y4?{�'���m��e��|2I�W�F�V�?--��pV��u��4�=�4Yw�G{�>��J?�4⾅���]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>jH_���u>����:�
i	>���?�~�?Qj?���� ����U>
�}?^$�>��?o�=�a�>d�=P񰾓-��k#>�"�=��>��?��M?L�>RW�=��8��/�E[F��GR�\$�C�C��>��a?�L?�Kb>(���2��!��uͽ�c1�Q鼬W@�_�,���߽=(5>��=>�>c�D��Ӿ��?Ip�3�ؿ�i��p'��54?/��>�?����t�����;_?Oz�>�6�,���%���B�e��?�G�?:�?��׾[R̼>/�>�I�>�Խ����e�����7>/�B?B��D��t�o�W�>���?
�@�ծ?Ui��	?���P��Pa~����7�V��=��7?�0�,�z>���>��=�nv�޻��X�s����>�B�?�{�?��>�l?��o�P�B���1=>M�>͜k?�s?BPo���\�B>��?$������ L��f?�
@~u@^�^?)8J����V���������=E�=�>1�����=�@��v.���5��+=	�>��y>$�>�z�>t�>Z��=x��������ɥ����w�mQ�kf��{-�<�����ϾI�F��$��|)��4��=���0g	���˾p���.e�M��=�U?�R?�p?�� ?x�x�U�>ܥ���F='�#��Ƅ=R-�>�g2?�L?m�*?hۓ=l�����d��`���@��tȇ�N��>�qI>��>�J�>&�>�`N9g�I>"0?>N��>4� >a'=YH�-_=��N>N�>u��>,|�>ھ3�}?>+���Ǖ����}�����7M[=v��?+���@�[�V���U���U�	���L>-�/?A��=Ј����Ͽzn����9?� ���D����0�;��=t�3?��N?x�=51�����w>�[����KG�=��T���?�I!���=�9
?T𝾟g�=�2S��2�v�r�j����?yD=?��?��ߛ���]���#��xԾ�% ?G� ?pk�=?6�����I�����A]D��X$?�x?��=K?��6��h�@��K>0 �>4hw���=���>R�����.񽐘�=��>*�< ?�T)>�=D�>�י�+�O�L8�>OBD>�0>Av??�($?Z�i꘽�{����*�̨y>�x�>�<�>fA>�I���=�!�>>�b>��������Y�B�Z_W>���M�^��>i� �{=�ʛ����=��=�9�Q�;�0-=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ3��>��P�������u� �#=��>6H?�`��W9Q���=�s|
?�?\d���� �ȿ��v�	�>k��?��?O�m��<��l@�b�>V��?]cY?b�i>~۾�{Z�[��>�@? �Q?��>�@���'���?ݶ?!��?�I>���?4�s?�v�>��w��W/�>8�������=�^;Kr�>�q>����ubF��Փ��e����j������a>Ƨ$=�"�>:Y�_9��u$�=���HK����f����>,q>�I>�X�>�� ?�a�>���>��=-b��逾������K?���?-���2n��N�<Y��=(�^��&?�I4?"k[�}�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��F��<��K>*4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��^S��GB�>�e!?���>�Ү=j�?�'?X7h>#��>p8�{��s<�_�>��>v� ?�1c?��?gb��`I3��N������d��Cp>�n?y+?�޽>�!���쥿�͠��bĽ�ϯ����?��I?�y9��}	?�r�?�J?Q4F?�>�>�����i�xRb>�W�>�͠���3�ʮ*�����t�>$�
?{�?�<>�`8�#���xR����	�?`�R?�j#?����;5@����I��=�S��,���=.�Bb>��u>�o
�^��=���=��>�#�Y�r�8YM���
>���>���=wM��-��,=,?��G�~ۃ���=��r�;xD���>�IL>����^?ul=�
�{�����x��	U� �?���?Vk�?n��<�h��$=?�?S	?l"�>�J���}޾D���Pw�~x��w�o�>���>e�l���I���ؙ���F��-�Ž��*�>�*�>��?�X?�qb>�P�>D���'�νԾ�6��]�x����=�Ol1� �����@u�@�K�GǾ-L���ϋ>OAH�j�>�
?���>y�>hT�>u&��>�$>�ǁ>,�>;�W>7�`>́>,V��D�hKR?����'� �辍����2B?�qd?2�>�i�ꉅ�A���?]��?xs�?�=v>�~h�b,+�n?�=�>Y���p
?�Q:=k?��4�<U��O���.��E���>�C׽� :��M�3nf��j
?�/?;��ˊ̾�;׽���D^=:ׄ?��(?�"'�Q�M�pn��qW�.�P���Rj������%�%q�w���v?��Dr��P&�ˡ<==o+?��?s����P���W�i�Z�<���q>r�>��>��>�OF>Dh�#�/���[�C�'�nZ��6q�>�z?1`�>��H?-0=?VR?t�M?�9�>�1�>�G�����>p�<�ڥ>�,�>1:?�*? F-?
?�^,?�d>>D�S���پ�
?U�?:�?��?�?�����ଽ[5ۼ2�����}�<��=��<�(½<�]�� G=:;Q>dT?ƪ�ޫ8�i����j>�y7?���>!��>����'����<���>L�
?qH�>p����mr�DY�4J�>F��?�����=S�)>?��=����^hκ���=ω����=�����;�M <χ�=�ʔ=,�q�'�O���:�ψ;���<��>�?|Ċ>�\�>����N) �B���w�=�Y>��R>�K>)پ9����$��Y�g�^)y>�>�?�V�?�ei=���=���=\q��b���V�~����V�<�?�#?�T?�W�?��=?�l#?��>.���D����������e�?]�,?B/�>G���ʾf����03�Cq?qj?��a�b��5�(�3�����ӽ��>]�/�/�~��,��-]B�����������D�?���?��D���6�94羜���0鬾 �C?�Q�>���>���>j�)���h�����>>$��>��R?,��>��?���?��m?���>A� �A�ȿ�1���,>��J>
�{?K�?�,�?A�T?2��>��>X�R>�ƾ-J޾��z��q:�U���������=	�n>͍�>�E>e3�=M�$�H(*��'����>���==8�>��>��>� '>Mm���G?���>g����E夾&ă�r;��u?���?�z+?D,=܅�"�E��*��c�>�i�?��?�*?h�S����=��׼/���Ջq�b�>,й>(�>^�=�?F=o!>`��>'��>t���d�(c8��MM�N�?�F?H�=~���i�_��������
�¾�zU�(�<�,����<@����O��v����F��W7�4	����������?��=�>�j��>��=�ؼ��=�V�꤆=�#�/��6W��ș<�tb�4%���#�`xB=p>��˾)�}?�:I??�+?�C?^�y>�<>��3����>m���V@?�V>۠P�8���˄;�$������%�ؾzx׾��c��ɟ�JH>`I�$�>O93>KK�=CS�<0�=�s=n=:�Q��=	"�=XP�=�h�=��=��>_U>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>lv>�=@oM���/�oSd�9N{�
��rd*?�a�e���>->�n����ܿ���s�=�g>�u==c�A�NZ�5�=�����K<Q~=�$}>�R>�?P>>9��^�=��#=�8�=�$b>K�<ʹ�>���o�=&>�s>�>�0�>�?_C1?�?e?�ϼ>di�+�Ͼ������>$O�=�L�>
=��E>�r�>�6?D?�?L?�̲>�=R��>��>��,�N�k���F��=�<�O�?k�?��>���<�|G�s|���;���½�?t�1?Mk?-�>����>࿪&�ۚ.�Z���
κ.�,=��m��K�)����Z��� ��=�2�>���>�q�>�x>Q�6>��J>m�>��>���<W��=ٌ��Ј�<���0��=ņ�����<n�Ǽ[�/9�<D��35�ı����;���:B}Y<��;���=���>��>���>�m�=�ò�s->
��D�K��b�=�=��#B�+Qc�u�~�=:/�x�5�D�D>��X>1(�����F?�W>р@>��?�u?�">���"Ӿ�Z���a��V�.�=��>:<� .:��h_���M�~�Ҿ�??*J�>c�?�̾>d���������
�&�`�NGR?i=s�2t.>w7=<����$���~s���S4�4�>i?)̈́�$�~>�D?ZHb?�w�?���>��2����z�$?�	3�u)�>��X��v��_®�u)>?A�?PT?3<��u�H̾����޷>@I���O�*�(�0�E���̷�Տ�>�����оd$3��g��������B��Mr�r��>��O?��?n6b��W���UO�����)���q?f}g?��>vJ?`@?	&��{x�q���x�=F�n?��?=�?I>V��=C3�7�?EE?�1�?�[�?J�2?�(���{?� f>ͩ�>�l3�+S�>r@��:���XaV>��0?6^�>c?Wy��9�&�\�þmI����_�>s�=��8>j�D>���<���<��<��׽[w�>��>�|�>��H>Q�W>�V�>t᡾��)?9>�9�>�;?ŵt>�F=��q�%=~�0L���������+뽪�=�n�<NI=*_��s��>�fſ�1�?��M>VW�R�?Se����J�ς1>�G>@�н�r�>�>+�>?��>P:�>��>�7�>z%>�Z��0*S>����&�ٻ:�[QC�o�ǾS�>���7P�v�������}�����!���b�4���� (��k=���?[ҽ�o�>f5�p\�in�>Ks�>AT;?h-���M�,>&��>�>�>J#�f��4���Ā��j_�?�4�?�2c>��>��W?"�?+{1���2�|rZ���u��!A��e���`��ݍ�����U�
��)����_?��x?`wA?�Β<cPz>E��?��%��ۏ���>I/�-;���<=�&�>�$����`�ԬӾ��þ1.�oHF>#�o?��?�X?VEV��\l��&>�7:?4/1?Q�s?v�1?��;?{����$?�X3>��?��
?��4?��.?<�
?�3>���=-]����#=x��Bˊ���н��ɽ���4=}='985<��=���<
���{ؼ���:g���<A�<��;=�9�=���=���>�@]?�!�>U�>͗8?)���m8�O[��ˎ/?цQ=8�}��ы��I��"��*�= aj?��?XZ?�Mf>�C��E�!>���>��+>�]>D��>ky���=��z{=�X>��>>�=�P3��ɀ����H����<�.>ћ�>�3�=����v�>o��q�q�^P>8D�L�a�r���9A�Zq�qA��>`�D?UK%?7I�=��;��ýEY��?ZG?�I?�i�?ç6>���1^�\�W�w\2����>P
>%����/1����9�e� ��֢>CP����a>����޾�n�� J����;�Y=ao�Ǧ==f��Y�־U�{��e�=��>�t���� �^Ֆ�ao��UJ?~Ax=����W�������>�w�>Uǲ>,~5���x�w�?�����q��=\�>��;>5�O�c��[F������>��B?GF\?=��?�ׁ�'�o�A[?�2����̢��F��p?�Ϟ>��?,4>v��=V�������b���E��b�>���>>,�-vG�sN��0������䆜>u�?c�>��?�mT?�`?Ib?��(?cp
?�>���R׺��&?1q�?�p�=X�ս:�T�V�8���E��c�>9G)?n&C��I�>}l?��?��&?�}Q?Y�?�D>� �oB@����>7�>I�W��2��U	`>iyJ?:³>�tY?�ǃ?g>>&a5��d���t���t�=&� >�*3?�K#?�l?�0�>��>꠾y�s=���>r;b?⤂?�ro?���=�E?j2>���>�[�=|�>�Y�>�?i�O?P�t?�I?���>Ȏ<<���%����0q�u*v�a��;m�D<�s=B��%�s�V�����<��;뼼�B}�����5S;�T���a<���> ��>萚�c>nҾጾ�K>�_���	��6��U�?�,,�=�nx>a��>Y8�>qz,��j.=4�>E	�>���w(?]a?�8?t�><6]�]G߾)e��ޚ>dB@?c��=l�g�?񔿈�y�q�=/�f?��\?�i�S�����b?��]?~h��=���þ��b�-�龵�O?x�
?s�G�k�>��~?��q?N��>��e��8n����Cb� �j��Զ=_q�>Y���d��?�>�7?JO�>#�b>d(�=�s۾��w�)p���?��?G�?1��?�-*>A�n��3�����e��� ]?+�>W���� ?4|ʼ�"Ӿ��u�	ȉ��@�㬫��_��q���������!� >���GʽKT�=}�?�p?�r?d�Z?4N���$_��~]��@��X������/��A��D���I��:q�����*���鋾Sc�=�qJ�_�h�;��?��L?�dȼt�-?���|s�L_C���>��f�I���NB=Z?2�E	��Ԟ=�g�ii	�W��c?�
�>?��>}CT?��Q���M���Z��H-�C�Ѿ~�=��>L�><�F>C�s�n�"���6��,�����_�/�u>�rc?�aK?.�n?s�w 1��l���!��1��A��ȄB>\>���>z�W�K��5&�w\>�u�r���������
�%N�=
�2?TC�>鸜>-�?y�?��	�{E���fx�?~1��{<ﱹ>*i?��>{�>m�нw� �6��>��l?��>��>Lu��MB!�'�{�H�ʽ���>�í>��>?%p>u�,�\��i������9��o�=Ŵh?}���a�[݅>!R?|"�:	iG<9{�>�!w�Y�!�߫��'��>�u?ǿ�=�T;>�zžQ���{��	��-?|r�>�Sվ���9j>��>��>Uy�>�kt?hz>A����SV�K��>���?�W?4]?<�1?I=v��;�aQ�I�&��>�/j>��>
==��<a�E���]<Bf��EU=��	��v���_G�:�l���=`�=8�>4Q⿎Cd�H�˾_L	����,��ט���[��x���0-�^������̗��t4��ԋ<���Kwv�E=��j)�����?���?n%پ��Ⱦ����zw����Ѝ?q_������$���DT<�wG��㲾����Pu(��dH�`"u���j�A0?�\�Լ��ߟ�٘����!?;�?�^o?���{�!��t���S>��_��$$�_j��������˿��5��Ag?J�>�Z��U����g�>���>�hH> B�>�x��Tp��
�<LX?V*?R7�>��.� ɿN¹��Cs=���?t
@�SB?1`'����>M=j�>��	?�lB>��/�T���n��*j�>c�?�?�fM=�xX�U�5��kc?L��<�kC����w�=�٤=�SD=%��2aH>9��>T�Z@�T�н��4>)��>���[2�7�d��<3�d>ҽ3v���ӄ?�v\��f�o�/�WR���P>��T?m,�>Bq�=��,?�3H��{Ͽ�\��,a?<.�?��?�(?�࿾�Ț>z�ܾ��M?G6?L��>�_&���t�sf�=�m�C|��i���#V����=z��>Zw>�,�M����O�ʞ����=���&iͿ�D[�����3���Eཌྷ��jyG��Q��⍾H����4�Ę�<Up(>�ǀ>15h>�X">�>7>:�R?d?���>�:�=}N�([j�B����v'=�����_��J8��)W�6���5ھ�J�m��w��%�+;k�S��xؼ��I�&��ǝ+�>�t���*���6?�=�v�sRS�}�����vg���Ə=޲�Va׾-�A��m���?EW?K���#Eb���0ս�>�2�?�0�7��ެ���Yg>�b>8�>���>���=Ɋվ.�*�ƴO�,d/??���������>9��D=į)?"�>�J�;;l�>��"?��(��'н67T>�">�Λ>a�>M�>}٭�1U�4r?�"U?�Y������Kϊ>����)�~���=[y>��+�-����J>�ƕ<���7U[�͈��	�<�8b?lF�>ԓ���&�E�2��T�==�<f?�ʟ>ܭw>�dj?h�H?�9=]I��RF�B}%��ؽ�
w?��v?��V>��ڽ��������i�4?dV?w�>�������:3��ƾ�n?�:?<b(?���	���D��۝��@?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?r�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>��������@>�Q����?��?/빽j�+>�=I�rֆ�Oյ�z�K>���>��;S�ҹ	���7��B�������6��a���ؐ>V`@L���߫�>X����濻Uȿ^x�T�Ⱦ͸R?��>�f��ۋ8�[4M��gC�/m��{C�.󂾸��>��>cv�������d�9b8��
=M ?�.����>$9���'��Q����<�ח>9q�>혍>�"�luʾok�?�R���ѿ�=���4��J1?���?���?v�?|)�=��^��y��;�=�oq?%F�?�&�?���=R���Q�����?%c��˨%�K��L��t�>R"?�>,pN���/>h7�>�I?E�P>[H&�dп��ſ����tt�?���?�׾�Ee>If�?�_e?5#F�����l辗�%��ؽy�?R���|���6���a��a��?P�G?���p���]�_?*�a�N�p���-���ƽ�ۡ>��0��e\��M�����Xe����@y����?M^�?i�?ϵ�� #�e6%?�>d����8Ǿ��<���>�(�> *N>jH_���u>����:�	i	>���?�~�?Pj?���� ����U>	�}?N��>�9�?��l=ɖ�>w�W<�����=x�>.Y�=��f���>�+>?���>���=R>���+�JL�]�D������>���<>�a?��G?t)a>(mս����(�'C>�R��a��7:����{�M����>i=)>w],>S�j�g㾈�?/h�O�ؿjg��:O'��54?(��>��?��q�t�����?_?�l�>�2��+���)��zT����?�G�?&�?-�׾]K̼K>�>�B�>e�Խ<���}��Y�7>��B?����>���o�#��>��?/�@;Ү?E�h��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?kQo���i�B>��?"������L��f?�
@u@a�^?*�
ڿ ���p���̡��x5�<��Ὕ�E<|Ľ%-�>���=��]=j|��6��Y�u>�˟>G	�>3;e>B��>��=�ρ�3J��磿����ⶀ�
�]�3��ӽ?�վ��齦������������ƽ~��=�Mg<�4쾿���V޽t#�=�U?��Q?\�o?)� ?D7y���>-C��!P=�f#�DB�=���>�N2?��L?X�*?��=TL����d��d��k"������J�>vjI>%a�>yF�>o�>�7�8f�I>&w?>m��>�� >��&=�pۺ�=p�N>gV�>"��>vV�>�����4>7���8W����x�6W�f�\>'ѥ?��ƾ�4��B埿��j��v�����>J)>?3n/>�L���7�����B?
������玎��$�9B<?��\?��0��,}����<q�2>9�H�PKվ=>���;���e#��>�z8?�>v��>A&A��gR��Sl�]z��EZ�>ox ?_���⪾��n����f�#��>	5�>z�_�7dC�:�����M�ں(�L�A=3{*?�! ?s���{HC�����5�¾-n�>��n>�4�=(	�;L>q��U&A��Dl�r
�=��J>G�>\?�	,>���=ꚢ>���|KP�ҩ>�C>=�0>l�>?�#?��#�o�����w�'�vhy>���>L`|>eH >�=K�p?�=K��>b>j?�>܄�����vB�)Y>��}�,�_��r�Y�w=�졽f'�=� �=%��˗7�k�,=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ8�>�����p��Au���(=@��>vH?���~zP��-<���
?��?n���{��@�ȿʏv�Q��>���?��?ɇm�:��
@�tJ�>Rj�?%�Y?�Ij>��۾�M[�Ȍ>r�@?��Q?J��>&��m*���?�ն?���?�_m>�?���??��>�<q=�% ��\���Ȕ���M=x�= ��>�K'>`��`@�V���_9y��|_�=H��Hc>2�8=^��>Sʽăľ��>�Ӷ�	��9���&�>��=�U>�x�>�C?��>��>X��9sνf�F�-���w�K?V��?��e�m�{�<p=�=L�]��Q?:4?�W���ϾyG�>�]\?�Ӏ?; [?�3�>�1��5���ڿ����u��<�}J>���>N��>S���nQK>g�ԾxlC�:��>Y�>琥�Iھ�ǁ�w���R�>�\!?jO�>���=ݎ!?ە.?%�y>/Ι>�I4��܆�w?��>6�>�3?b�|?�?������>�#���2�����[�(�>��x?6�'?;�>T.���%������]�<�?=�׈?&�8?�?%��?�,�?Z�9?�8B?�e>2s��*�=��<I��>�?��c���C�_��U���Ř>�,?�r?횞=�����)&��䔾]�G?|\?�
J?O���e���c�=hUp�H�K�M�w=�8T��1>���=����V(>�1]>>�=�����l��ۂ=ְ�=���>�M>��_+Ͻ,=,?�G�vۃ���={�r�9xD���>�IL>�����^?ql=��{�����x��	U�� �?���?Sk�?���;�h��$=?�?M	?y"�>�J���}޾?�ྵPw�~x��w�b�>���>��l���J���ۙ���F����Ž�^�F'�>�r�>���>.~�>�Wt>���>�5��0�.�Ki�ބ��Tb�lK��R>��{��d����4��H�uн��8��P��>b��n�>!?��X>�ޏ>���>! �ft0>/$޼���>��>lȔ=p�>s�a>��m:�l��<R?W���K�'����Ӱ�MB?0pd?�'�>	3i�p������St?$��?�j�?%2v>"xh�-5+�	i?�;�>����Z
?�	;=���b+�<]����U����x����>L׽v:�,M�}�f�t
?�#?e��ˎ̾��׽A��E�n=��?3�'?i�%��O��Cp���W�_DN�7��Zih��ޡ�P$�)r����lu��J��2�%���(=��*?�I�?�f�}����?Yh�  <�Ǒk>��>/�>C�>�N>�	��e3� �^�p�(��߉��:�>�_~?O��>NLI?é;?�8P?3,L?Hf�>�N�>Х��oQ�>}#�;祠>��>�L9?�.?�>0?h�?1�+?�b>�������=Rؾ l?��?��?�?�?�E��nG��Z���r�{�x��J~�"}=kķ<��ٽ��|�)�]=�T>@p?~;�=�v;�]��v%�:G2?��?�ι>�M�����.7k����>~8�>��>�s�[�i��f*�G:�>�ow?�PY��7�<b77>>ّ�;JQ��A�=NE<��ټ��=~���#��*W>�S<Kx��$���=���=���=XM�>�??��>22�>�J{����Ћ��=�
f>8}X>�U>�,پx>������Ctf�c�s>wU�?�J�?7d=���=5F>?�����¾k�	��ù�"�=׀?$^?J�R?D��?8�=?b� ?	U�=�������;��8���\�?,?:ȑ>�����ʾ�⨿�g3�Ī?@?(a�P��)��2¾�cս��>�8/�})~�������C�-d�z����8{�?`��?	0A��6��q�&��������C?	�>�@�>Z��>��)���g���;>U5�>��Q?(��>!�]?K*�?��z?
~�>��8�ſ8{���w�<	,�=Hz?
H�?�J�?3UO?XKQ>d)>�繽x���\��-����w��3<�n>>y��>�s�>z |>Y��>niQ����퐽���<.'>C=?�Հ> ?�>��#��G?���>�q���P���������T.:�Iiu?���?lX+?��=���@�E�q���l��>m[�?7�?��)?�SU��p�=�}׼�m��(q�pp�>�V�>�5�>�Ǒ=�mM=~�>�u�>�{�>�$�p��k8���P�9e?'IF?�ҽ=�ʿ��#�a�4���*2��c���M�4A��}u�tF�=:늾�2���̾��l��X]��=]��븾�𚾻$����>Mr=G�>I:�=�=f\��=���=e.�����<<��ٻ�;��?<��k�����'<`��;O�^��L��˾��}?�4I?�+? �C?��y>iF>L3��>ę��N<?OV>�P�W����;�,����&���ؾ�p׾��c�!ǟ�P>�<I���>�*3>�;�=?I�<���=?;s=���=J�S��7=��=)^�=�c�=z��=��>IO>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>x<>>!�U���9�_T��h!`��6ν��?��&�4�?0>/��=������'Q�=�6>�갼�8���L��z�=[�4���D=�=g >s]>�?s=g���>b�=7�	>��>Y��<�U��>�����<[;�=�y>0->d��>p�?�b0?|Ud?�>�>�n�B'Ͼ
G��P�>s�=%E�>��=�pB>䀸>��7?a�D?��K?��>Ǩ�=�	�>s�>"�,�̲m��m�vŧ�� �<`��?�Ɇ?Oո>�{R<��A�̝�h>��!ŽTr?_M1?�n?M�>�X����6M&���.��$����>�s�)=Tr��S������(�5����=FT�>#�>��>	y>��9>��N>~��>ώ>���<�=�4����<w����=(ߔ��'�<�
Ƽqс�QI!�V,�V���u�;�2�;�bQ<ȶ�;+��=yT�>8>.��>)�b=?e��YV/>1���-�N�ǀ�=�C����>��c���}�4�)��=���5>o,O>� ���q�����>�dh>�2C>S �?�u?��>�*ӾL��l��e�;��=B��=14�f�7�^�X�/M�3MԾ�J�>�*�>\v�>�ڭ>�6�^ �� <���~rf�^�1?����OD�=<>>h��h2��ir��b	1�Lm\>"oP?�W���>�g?�]�>��? L%?�(��^ �i��>�t���|>�@�d�$��^;��7?�.>?hk�>Mc�)�f�.b̾����i��>��I���O������n0�[��ͷ��߰>�&��GoѾ5�2��Z��R؏�gB�zr�v��>UO?�ܮ?�8a�Ff��eOO�ސ��ʈ�z?��g?��>,?�/?j���/쾱7��ո=�%o?���?1��? 1
>̜�=ר��, ?I�?;[�?r	�?k(d?����ɷ>��=;��=LQB���>��l=�V���)=��?��?�?Էὼ���ʾ�Ⱦ���>��>�~>3��>��}>>�����f=���>�b�>��>Xy>�B�>r�>M���}B��0?)4>Z�>)�O?��w>���EC�3>�9�$s����������%A�<7"�<2��=���<�Q�>�ȿ�?>l�>�����?����e���>d�v>T�G�+�>o =��G>���>�+�>��`>ف.>�=Ӛ����6>-ZܾJ�c��V<�)C꾯�*>�U�\_��[��h�'xB��	���}[���v�[��LO=6��?�~<�*c��6��?��=�?��>�dG?f��}��UE�>��?�Ɖ>� ��r��������
��K�?���?��b>/	�>_�W? �?��1�O3�?]Z�ڙu��A�~e���`��䍿;�����
���Y�_?C�x?�]A?��<�nz>��?��%��菾�3�>�(/��;���?=V*�>�����`��jӾ�Vþ���@=F>��o?�"�?�F?}wV��Zl�L9'>�i:?"v1?48t?*�1?i;?�����$?BQ3>^?�??�45?%/?��
?��2>dk�=_���$=�命�Њ���ѽzʽ����4=*_{=�N��k�<��=�<��\ܼ� ;����	L�<�;=�͢=��=P�>D�U?���>��>J�;?���7a;������7?�_=�^���l��P���(��#i�=Z[e?h��?��V?u�S>��@�z�2���5>3:�>_(>�j^>���>��	�T�f��j�=97>w>��=���[��K��]����w�=RI>�(�>}<_>�)���4'>6go��]v��]5>f$��H����(��6�u63�F]�~T�>دE?h�?yF\>�޾��%� R]��?3\?�:?O~�?hɖ=m���G�F#�0����_Z>�V�=~Ӿ�F��t�����F��4L����>����8��`S>u� �뾄jx�s�S�S�ƾ���=J�.b�;����վ��I��C>�(9>�A��n%��-���"O?�d=+������?��x>1N�>��>$�ǽDN��rD��鴾���=BH�>?`I>�Vu�XV�OP��=	��:�>�IE?@M_?�c�?�-��xs�b�B������\���ȼ��?���>gX?��A>���=Ң����c�d��G�t�>���>���G��=�������$����>�4?�d>5�?��R?��
?O�`?%*?�I?�%�>-��x����@&?��?�=��Խ��T���8��F����>R�)?��B�B��>Њ?��?8�&?�Q?״?��>n� �?A@����>�Y�>g�W��a���_>��J?x��>>Y?�ԃ?�=>��5�e����q�=`>)�2?�5#?�?J��>x)�>x���F>K��>�9m?X��?}�\?�-==�?]>���>�?<ؖ>�z�>�q?I�U?��}?JVI?t��>�#�<N��D��+B���2���'�<�j>=��W=�b���B��\����̻^�:����JvD;/.
���X�Bބ<�~<�O�>��s>����0>V�ľ�S��H+A>)G��NF��M���վ:�(߷=���>"?%��>E;#��t�=y�>u�>;��^(?B�?�?�6;~�b�� ۾:�K��/�>�B?i��=b�l�6y����u�k_g=��m?i�^?;~W�4���pL?~1J?���z�J���`=�hu����J?͞�>3���O��>c�?ˋS?��>�ƽ]FU��疿ld�&�1��K�=���>�����c�@��>�b1?��?"��>K�F>q�pO����ʾk(?|��?H]�?�\�?l�r>��c�2�࿡�𾮾���l\?"�>����s&?@._���Ծ3��S͆�еپȢ��%:����Ӎ��V���>{�'뺽E��=rC?�&p?�?s?�qZ?���9a��P[�8�|�n�Y��{�� ���>���B�,�F�Nzs���x��{a����x=W�)��8>��=�?z�-?⛛�\�?��������t�X�b>4�w�K�� ,�=I�<W<�
T�=������ƽ�xb�ҥ!?|��>��>|�7?X�o���5���'��s2��U����>ڷ>F�>��>���^�|�@��=QK��q�q�>�X?@X`?���?U�=Q��S͚�SqA�n=��ѽl��>}��>	l�=ָ~���G�%��p���6V��j��Ӿ��&��o<�T�>+�>��>���?k��>�p
���ľfPþ��2��}=���>ф�?T4?�ʶ>zs��qS��z�>3�q?f	?�S�>ۧQ�=�������c�C��>��>�?��>U<n�|�j��W���o����/�.:$>�7e?)c��%�}���y>w]D?w-�=y��tQ>��7�������P~��->IS�>}I>>ޒ�>뉾�7���䱾`� ?��?�7�(���W>Ŝ?�<?(�>x�?d�O>���rr潣> ?RJ]?�SG?ZE?<��>ܳ���������Q'����=�H�>? `>��=�ђ=/*
�߯c����?��=N^�=���9z����X"�;��<M`q=�fs>�����h�A`Ⱦ������D�'�>�^e2�{n|�L�½[	���V�����t;e�{�+=I��+�`��^�h�J��i�?$��?S'��V'p��������I����p?�Q����ҽ�b���������`���R�O��q�Y���q��d�m�'?����u�ǿ>����=ܾ[ ?�@ ?N�y?i�ў"�[�8��� >) �<뜼�뾫�����οC�����^?+��>+	�D��	��>۞�>��X> 6q>��Mݞ��O�<N�?�-?t��>�r�1�ɿ�����X�<��?��@NHA?f)���&d\={F�>�h
?kh?>%3��?�iD���*�>��?�?�\X=�X��	�)�e?�)<��E�UE����=3-�=}�=m�9/K>�!�>��~�A��ڽ	�3>S��>L-#�""�{]�3"�<��Z>ڶֽ%\��4Մ?*{\��f���/��T��U>��T?+�>d:�=��,?Z7H�a}Ͽ�\��*a?�0�?���?$�(?;ۿ��ؚ>��ܾ��M?bD6?���>�d&��t�ޅ�=`6Ἐ���{���&V����=[��>[�>,�ދ���O��I��g��=���".п�������:ǽ���� �������҆�q���s����y���>��n>���>�F[>�~R>�Md?z��?�c�>q�A>/1�k׾ִ�Ҝ�=�>R�/�6%8�D7�����������ľ["��$&����Lо%�F���=<vJ��鈿 <��Is�d�#��s>?F�=�&�Gj?�b��<�Ⱦ��Ɉ�(��=U�������8�f`����?�&A?�E���ur�A*5��´���>��~? ז���$�sg�� �M=d�9>qO�=W��>��9>a��<a��^�|B/?�p?�2���8��׶&>����`:A=6W,?��?T?���>�>M� ?6$��Zٽ�a>�A>ֽ�>6�>�[>���~ὰ ?��U?+t� N�����>�žU�w��Ox=>�e$�F�����R>ϱ�<1v������FG��h=�T[?���>e�"��������Qm�	I)=�Tp?m�>�4]>.qk?�RV?:�=������a�v�,�N2�E(f?rv?y�>��м1�߾�3��95?�![?�3|>���W���2��|
��?��s?��+?�'��X}�����UO۾�7?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������Rb>�#�z��?��?	�v�˘>��!�y��j��Y�j>ՕY>O:�=dF�=��"��fQ�@ž<߾�4�n�>�D�>�{@f=�'
?(_���B�տ�qv���޾�x��!vJ?�F�>sd�Q����a�\�s��3f�����w���>�>������K|�� :��¼���>T��>pfK�Vդ��:��Sd*�-��>���>>br>'�Ž�)���o�?���9�̿�������EoV?�S�?���?��?���?���|�p�W�<��G?x�v?n�Z?x��_a��LH�zcs?A?���?��7���&���N>�)?��>��5�.s=�>s�+?u%->&**��8��Ŀy'���?a�?	���2�>Λ�?�=?�X�� ��Uɾ�G;�H�<�fm?�us>���4%�h\6�M�<� w&?)$?
�~�^��\�_?+�a�N�p���-���ƽ�ۡ>��0��e\�*N�����Xe����@y����?N^�?i�?ֵ�� #�f6%?�>c����8Ǿ��<���>�(�>*N>fH_���u>����:�
i	>���?�~�?Pj?���� ����U>
�}?�#�>��?<i�=�`�>9`�=��D�,��k#>\�=��>�a�?��M?hJ�>5V�=�8��/��ZF��GR�j$���C���>d�a?S�L?�Mb>���9,2�!	!��nͽ�a1�64�/Y@�ə,� �߽�(5>y�=>�>`�D��Ӿ��?Dp�5�ؿ�i��p'��54?1��>�?����t�����;_?Tz�>�6� ,���%���B�b��?�G�?:�?��׾�Q̼�>9�>�I�>D�Խ����]�����7>0�B?W��D��s�o�~�>���?�@�ծ?ei��	?���P��Va~����7�c��=��7?�0� �z>���>��=�nv�޻��X�s����>�B�?�{�?��>!�l?��o�P�B���1=9M�>Μk?�s?�Qo���g�B>��?"������L��f?�
@u@a�^?*>������9[����¾�m�='H�=��>Q����@=a�Y=�U���<_�~>�Lr>�Ɖ>��Y>i�0>1�,>+O���o �Ǖ���J����F�k��D����V���������/ ��������b��G��^��V*������м���=mSP?6_T?��q?�w?�a���=�;���4=�4�z�=�]~>�")?.G?B�&?@�=�~���`��_�����c������>��7>z��>�j�>��>��<�|R>��5>�{>���=��c=�,�;?�4=?�Z>�X�>3h�>�z�>���<���=���昭�2�������8�>���?FF/�FhW�T̢�<�žYx��}t>��B?�m>�i��vV˿xc��o3?M�M��'�hRl�S�>�o$? /?�W�:������m�z=A�������,s"<�Y�ŕ���E��,�=˿�>K�=zE>��j��oD�?�N�l��H?�*O?.���Mkξ�܇�#l,���Ͻ���>E�?�1^=���퍿�F��������GW?I�?J �=�C��}�Ⱦ���Φ�>���>5N>�2;�H#=� @��>������->�[�>�-4>�?��%>1��=�/�>�u��GHC���>ɕ;>�2> ??�Q$?g��1��'K����0��Ax>���>`��>�	>�F���=d��>��c>�8$��Bz��Z�&"C���Q>��i��w[�-�t���q=&����=̿�=UO���:���(=�~?���*䈿��Se���lD?Z+?� �=0�F<��"�G ���H��I�?r�@m�?��	�ݢV�7�?�@�?��Z��=	}�>
׫>�ξ�L�ݱ?��Ž4Ǣ���	�<)#�hS�?��?�/�Zʋ�;l��6>�^%?��Ӿ���>���2��!���u��6#=v]�>�H?�����(T�`w<�N�
?�?��'���Zɿ�v����>��?�۔?�km��D���)@���>m�?%eY?f�j>��ھ�[���>��@?:5R?K�>�0�:)���?�˶?䨅?�Nh>kڑ?Jlx?��>��6�'�xȷ�zH���<�=��=��>�><��,�U�(���Ն�g�e��n���~>~"�<���>_P��h֢��B�=^���Ǿ:�c����>M5`>45s>O?�>��>,R�>�b�>66F=!X���"���XK?|E�?���n�2��<���=}�X�t�?Tn4?�'��yѾ�o�>�-\?mÀ?��Z?�K�>~{�)�������f��ok�<�wJ>~i�> ��>����/fI>"�Ծ-@�L��>\'�>T:żθپv���ػP�>�.!?Q��>���=p$?��!?�^>U�d>�6���x��c6��ɠ>p�4>�6�>m�?�g6?+��� �d�K����i��v�o���>�?�&?/��>��������,�ǽ���-vG=�?��?=�ľR��>��?��A?�m>?���<�=�5�پH=G��>�K
?�ʂ���J��5�H8S����>�B$?=�?�C�=����@�l��%���;�,.?f�X?Qg'?�v�V
_������}9<d�Z��2��=�5�=t�o=$��=��O�s48>�j>D�;�����#8�"��<r�#=Ǚ�>�y>x����=,?��G�>ۃ���=G�r��wD�G�>>IL>�����^?'l=��{�����x���U�� �?��?Nk�?o���h��$=?�?:	?"�>�J���}޾F�ྌQw�/}x�:w�D�>���>�l��O���ޙ��mF����ŽR�>�>¾�>v�?��?��S>�k�>���{%��u�o��$^����(�7�D�/��Y�����!��~��þ����yѕ>�w��տ�>.?�j>
�y>�^�>�1��5�>�aO>l��>��>B�U>O]7>��>0"�;ѓսF�Q?Mg����'��1��8���A?��d?���>��k������ ��K?C��?f�?J�v>	h�h+�X�?��>0���I
?�V8=���R/�<�<���H���Iy��Q�>"�ؽ4:�tM��e��
?�1?����z̾y�ٽ�܎�`�<i�w?��?�n#��;��ii�J~M��_C��䊻4!�`m���D/�[x�%�&u~��́�n����=��2?೅?%��~�	�A�ھ�<k�2����>��>o�X>�]�>�s�>_����?��k���@��?��Չ�>"#�?���>L�&?��*?VsF?�D?���>�^Z>������?�W�=�q>L'�>U?Ζ
?G$?RW/?&~2?��U>�B���Z�>����?��?"6#?^?]�>������%�&>}e*>�����H��dV��<X4����켢��>u�l>�+?��=nY)��D
��]>Tz#?�.�>��>ӈ�� ������=�� ?�}?��k>�_"��1����!�	C ?Q��?�����iL<�n:>q �=��&=H��<�.>sT)���S=�m=��G�Y�<� p=�w�=�R=��ջ�'̽�zE=�#�=���>l�?�j�>fG�>�k���ᾎ��0N=X�T>X�l>)0>���Pۄ�����_��n~>)ˈ?�]�?�he=�c>�n>�8����Ͼ�����Ӿ�Y�<�A?�'?��O?g
�?XH?N4?Ӄ=��,��d��V���탾�@"?,?T��>���9�ʾ�憎��3�(�?.`?�>a����?)��¾E�Խ|�>#P/��)~����dD�[y��������/��?0��?��@��6�)~辮����P���C?&�>�V�>�>ȹ)�>�g�L �a5;>���>�R?Od�>pN?%>|?�?]?di^> 5�r��$癿a����(>:�@?,��?���?��v?���>��>�6!�b�޾�A��p�;�58 �^����;6=�Y>�p�>:�>3Ū>6��=��̽������F��Ǯ=i�f>n��>��>aB�>�v>鮇<,�G?���>�0���z�	ä������<��u?R��?l+?�=z����E� ��"W�>m�?��?�"*?
�S�st�=�:׼���rq�v�>���>�>�=;�E=Zn>�>=��><�pY�a\8��?M���?i"F?���=vʿc�t���j�g���^���J ��|u�՘����S�4��=6���@���9̾s�~�%f��������䥑�:bu�)?qE�=�3�=*2�=�N<b���cω=���=�[+�I_��Ϗ�ɞ�=%+_�"k�<��¼s�'j)�[�U��TE��_���]r?��P?��3?�vH?��>�#�=�����~�>5���?��<>LD���F.�E荾}Ry�pqѾ��޾h�t�x��:~>�蜽�->-	K>��">f�'=">1�=�=+�)����=���=�=��=�m�=�t">�_'>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�5>�>4?T�z�2�< c��?l�!}I��#?|�:���;t?v>%��=iAھ�ͼ���K=j 7>qCI=*"�%]�")�="[z�0�C=�n=��>-�F>G�=ٷ����=�T=�=�O>����7�]����57=!z�=`�Z>}�*>*�>H2?�!N?k�o?�w?b���A�Ҿ�fؾ��>�P9>���>�<�|>��>-?�[?�]o?DG�>��ּϻ>0�>���_������ͭ��~?�]e?5��>H�ɽ���l�6�E;��(b�%�?a<?�H&?���>|������%�GE1�4��]e =MW�<�D���#��(���3��3��w�<�U�>��>h+�>�D�>��:>�U>�p�>΢>b�;f��<�>_�J����]�漝=���^к�)<>g�<�hg<$n��Y(m�q�<��0=	�=zo�<�=`��>'x>)��>�x�=ǳ�� />�֖���L����=?���B��d��3~�f/�P�6��C>UX>���s7���?�7Y>�u?>w��?^Eu?w >�E��lվYN��9�e�`�S�V�='�>�=��U;��`�+�M�ȚҾV�>�D�>�=�>���>����_�
܎�\-���O-?��d���;>�a�K�f�G��������K�zO>�o?E�����R�Z?d�n?3�??�)�1�5��>��ռ#O��;�I��e��Ff�ݛ�>Fr@?��T?��$�GI�jE̾[%��
ٷ>EI���O�p���#�0���ʷ���>���о�)3��h������B�`r���>u�O?a�?b��U��/YO�����,��$t?\g?
�>0B?�=?�ڡ�[j�'t����=3�n?��?�9�?]>�>9K7����>��?��?p��?�-?�ܼ�J?#�L>�i>{"��i��>	�>���
�s<��X?l?1� ?^�
�B�2�?=��������S��jR>j��=�?>L`�>R_��٣;��=��<~��>'��>�2�>�-h>��H>x�>N�|���?���=�>5/?��w>.��<]⨽�q�<�+9���U�F75�0�o�/p˽��<��b<�e�<���j�>�%ſ@�?X�^>��.(?�����a���k>� I>i����>W�>�vj>U�>`��>.�=!�>#7I>�mξ�?=E��V����?�I�?�w�ݾ<*=>v����I!��X�o�۽S<��Z����\��a��_|���?�e��<��?6q����B�EA*�=�]��z�>Wу>�5?k�@�yzཹ;>t�#?T�c>zw�gT���ɉ�u��N�?���?�>c>�>��W?��?Ȋ1��3�*uZ�m�u�J%A�e�9�`�4፿f���+�
������_?/�x?�yA?�F�<�8z>z��?`�%��ԏ��&�>
/��$;�PB<=�'�>�&���`�
�Ӿ.�þe:�0EF>\�o?%$�?Z?�KV���N<�2">��W?�fG?�Z�?�P?��?l`��7�4?�5�>�|?e�>gX?*Q2?�J�>DΣ>]9x>{��<�U��\0i� �S��x�����ձ=ï>u�D>�e7=B�=$��<_��6���>`?�=@�:=��1=a_�=�x>�Z�=�l�>��[?�	?	�>�=?�=��ɿ,����2?�=y�t�~��l�����ھS�(>s�v?*��?~�a?DS>�B�c�B�ZO>�`E>�� >ԍa>M��>��ٽQe�G�=:�Z=�@J=N��;�0J���`������އ=�CW>v�>�yk>䭵��T>���1s��c>��L�˅���}T�,B�W3�.)y�|Z�>)�L?�]?��=���&�ȽH�c�J?jvB?N?]z?�M�=@)龫v?�W,>�������>���;V��=���e���o7�A9A�v�>ϲ���Ȱ���W>������r�p�N�KܾE��=���5�a�;���Ѿ֑�T-�=��7>������(�����������B?�}�=@՜��IK��깾�s�=\��>��>��W�x���3lD�sN��F8=%!�>�E>�r�:a�꾁ZD�V�
�G:�>��D?J�_?���?���mjq��B� #������t���?�>�s	?��C>���=L��� ���0d��F����>��>����6I�������E$�:�>��?�>�s?+�R?��
? b?89*?�?���>渶��U��:q&?�\�?�R�=�ͽ�lO��7��eE�<�>פ)?[@�D�>�?�?�|'?�Q?(�?�N>�6 ���?��e�>9�>7�W��ɰ��N^>�rJ?���>�SX?�u�?��7>��5�睡��1���:�=�">�2?��"??^?��>SVQ?��ھ��>���>�??w��?+�E?m[���k;?��>��>צ����>��>���>�NS?���?�46?��>���=���=�����p�����1�;���7�O=�J���6 ����X�<��f=GSս�A=ؔ�5m����'�r��X�>��s>��1�0>��ľ^O����@>:���dZ��7ʊ��j:���=�~�>��?���>�b#�ܳ�=n��>�G�>��0(?��?�?p�';%�b��۾��K���>TB?��=#�l�ׁ���u�q�g=��m?̈^?��W�
!��2�b?��]?�g��=���þ��b���%�O?�
?��G�	�>��~?8�q?���>r�e�G:n���~Cb���j��϶=Qr�> X�U�d��?�>��7?�M�>5�b>J(�=Ru۾�w��r��)?u�?�?���?I+*>��n�[4࿒����-����]?Q�>_ۦ��R#?#�뻄'о���3#��4!�������&���Q��c"��ނ��6Խ�r�=>�?D�r?o]q?�`?� �ƙc���]� ����U����rY��E�,E��C��	o���ߗ��)����WL=T�s�	!;�Ƕ?z�,?�N���� ?㹗�l���6���:�>�܂�y�νZU-;ڭ����><Ks_=��1��? ��W��1�?�=�>,��>"�D?�DW�_�7���0��5��uݾ�->�Z�>x�>a��>jk�=�$������$ܦ��Ә��|S��;v>eyc?�K?-�n?�`��%1���� �!���/�eZ����B>�o>�Ɖ>�W����5&��S>���r����;r����	���~=S�2?�&�>s��>P�?�?�}	�\c��u`x��1���<b-�>|i?�A�>��>#н^� ���>��l?
q�>�ڠ>����W!��{�6ʽ���>��>*��>��p>��,��7\�'|��5���:9���=0�h?Z�����`���>�Q?T�:�K<� �>5�x��t!�ш�K�'�I>l?b��=7�;>��ľ1���{��r����,?g�?��w��"���>��(?c�>�C�>���?9�>6T۾���?bj?��L?DE??��>j�<=L�����3?���M<��q>��>>=Y��=���QP�v�!�#7O=B2�=�ǘ�������l=4�뼷t<���<�02>�ֿ��P�'���@������	�zD���Y����K����-���Kp�"l[�O����/#6��cx��[��:�c�K�?��?hӔ�*�����L쇿1��w�>�����*D�⡋��걽�ᖾ/��@q8��Q
�	�[���|��c��T'?�̑�c�ǿౡ�h1ܾ��?� ?o�y?%#��"��8��� >�B�</���sX�z�����οP���'�^?#��>m�ﾓ������>��>U2Y>~�p>|k���랾��<?��-?�H�>}�r���ɿ�y���v�<���?8�@مA?ќ(����T]=ly�>`�	?��?>��1�z��m��Q��>��?��?�1P=W����3�e?5<<�F�NԻZ�=|�=]�	=u����J>PW�>
t�:�@�1��I3>32�>zF ����Zp]�rw�<�:]>�Jսg���5Մ?,{\��f���/��T��U>��T?�*�>U:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=x6����{���&V�|��=Z��>c�>Â,������O��I��V��=5: �B�ȿh�$���!���<�~�$����u������̼T���{�X�k�ʽk#�<��=sO>�*v>��1>`xM>œW?E�t?7�>Γ>4�2�/���;�ʾ�G�<\���R>�y/�����̐���־�P��������&��nľ4�W���<v�� ���C��is�A|,���I?�A>���9B`�3C�=Ip|��h���}d>��.����+I�A~c��/?Gt?뉿FCN�9���2$�y�?�W���,�u+�^E��� &��!q=w�?���=w�8�4-k���~��x0?oZ?�\���'*>�� �h�=��+?,�?JeZ<#$�>%H%?M�*�#9�L\[>b�3>�ܣ>��>2D	>v��b9۽q�?�T?p��g���Yې>�b��{�z�Ja=42>*:5��H�Ȥ[>-'�<����>V�&C���~�<�zI?D�>�v��<�G���W)����+>�t?���>O->4�q?++j?�q��D��i'o��bB��h���x?4!�?�:>����Q��I���x�D?��J?�6�>@���þ'*�=��w\?Ł{?��?�.K�+Oq��[��җ־DI7?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?~�;<��U��=�;?l\�> �O��>ƾ�z������1�q=�"�>���ev����R,�f�8?ݠ�?���>������ߞ�=$ڕ��Z�?s�?Z���FKg<���l�nn�����<Bԫ=��F"�	���7���ƾ��
������俼���>�Y@VR�(�>�B8�Z5⿟SϿ���Yо�Uq���?P��>�Ƚ.���
�j�OPu�ڲG���H�����S�>��>�b��y䑾m�{�f;�����>v��j�>��S�'��F���j]7<��>=��>^��>�%���㽾���?rP���<ο���T��M�X?�e�?�j�?Lm?#6<w�#y{�9G�	:G?��s?�Z?%m%��5]���7�˒Y?'�;�L��%�z�:��=�
>?f�>+�7���=cMz>n�9?��>�D�1 ѿkdǿ����I�?v��?��۾�x�>e�?#�?�	�;�����>}"�l(,>XS?:�>��˾�N�S���<��S(?b>?��N���.�]�_?)�a�K�p���-�u�ƽ�ۡ>��0�f\��M�����Xe����@y����?M^�?i�?ϵ�� #�f6%?�>a����8Ǿc�<���>�(�>*N>jH_���u>����:�i	>���?�~�?Rj?���������U>	�}?]$�>��?o�=�a�>"d�=L�I-��k#>�"�=��>��?��M?�K�>4W�=��8��/�C[F��GR�V$�@�C��>��a?�L?|Kb>&�� 2��!��uͽ�c1��P鼩W@�e�,���߽D(5>��=>�>j�D��Ӿ�?�V��ؿ�e��$t'�;(4?"ڃ>	�?n���t�Oc�K_?�r�>j?��0��x-��/j�4��?�I�?\�?+�׾�]˼ >�֭>�8�>+ս퟽k���8>?�B?��":��c�o�M�>���?�@C̮?��h��	?���P��Pa~����7�]��=��7?�0�.�z>���>��=�nv�ݻ��Y�s����>�B�?�{�?��> �l?��o�H�B���1=2M�>ʜk?�s?aRo���q�B>��?������L��f?
�
@~u@Z�^?+O�����i�����OL�����=��=�qP>9�R��=>⋉��l�p=�1>�G�>�{>�i>}�I>��6>Z>Vu���&�6s��s<���Ni�@�V�L����<�
��Ӿ�`-�e����䋾����yM=HԽג��ڧ��s@����={\S?~R?�Yp?�b ?YNt�m�>������<���K]�=�߃>��2?��L?��)?Э�=�9����c�ހ��k��筊��>C�R>D�>��>��>X����E>�&E>.v�>Y��=a�=����<�Q>{��>���>�7�>vX@�O�r�����_?��5�{�o\����$��*�?ݢ��.f�s���@���𺾚ŭ��[?�>���ǿFW���?������	H��:�>m<=?�?>���6徹�=���>h&r��\پ�����Bh��7��<8�� g�>vk�>�߽v�q>G�/�G��2Kx�o�)���>�4v?:	�Z���NX�(�Z�����:��>�w?l�,=c��z>���!��N����佭7?/	?��>6(�D=������-2�D��>���>�jڻ�:>*7=�8۽��K���\>��?>���=�5
?�%>���=�n�>�f��ui'��>��%>�T/>72??��'?�f��~���=w��6��!�>$��>��>��>�T9���=\��>w�>O""� ����4�פD���T>E��0DZ��1f��(�=�1v���=��=����(��d=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>��D����Ԇ�tgu���=���>MH?-u���_]��7�]?u�?�8��HΤ��Pɿ��v�� �>��?z��?�Ol�5j����?�p$�>���?R�Y?@Ci>2,ھ'�Y����>�"@?��R?��>I-��*��?�E�?���?�I>���?�s?�k�>9/x�nZ/�o6��ؖ���n=�[;3e�>3Y>�����gF�ؓ��h��c�j����a>��$=��>F��3��#:�=��H����f�7��>-q>��I>W�>q� ?�a�>L��>�y=�m��kှ������K?���?���2n�4P�<���=�^��&?�I4?ak[���Ͼ�ը>�\?p?�[? d�>.��J>��A迿/~��Ҫ�<e�K>4�>�H�>�$���FK>��Ծ�4D�^p�>�ϗ>>����?ھ�,���M��>B�>�e!?���>�Ү=�?�DB?Oǉ>Mj�>K\L�$���:B��.�>�PL>2�>q��?�;?x�
���Q�����Ī�n�d�ɹ�>`��?+%??��>�ل��񎿑�_������>Ϸ�?o�?�:8��x?q7�?/�L?�+?��>x�о�����6>���>��!?����A��?&����A4?�]?�-�>�Ó��-׽O�ټ�������%?^'\?9(&?i���Ha��3þ���<!'�A�P��+<�uA�>�?>s\��1U�=R>D��=�Am�V6�"�m<��= B�>v]�=m�6��p��2=,?��G�|ۃ���=��r�:xD���>�IL>����^?nl=��{�����x��	U�� �? ��?Yk�?Y��>�h��$=?�?Q	?k"�>�J���}޾5���Pw�~x��w�Z�>���> �l���J���ٙ���F��Y�Ž ��+G�>���>�?{� ?�.O>0[�>jN��SD'�%��J�t�^�wt�B%8�ڞ.���Ĩ���J#�t��� ¾��{��}�>q��(P�>7�
?H�f> z>z��>�Ż�t�>��R>j�~>��>`�V>>�4>��>o�+<Ͻ�KR?����	�'�g�辍���o3B?�qd?1�>9i�1������q�?���?Qs�?.=v>�~h��,+��n?�>�>9��Zq
?�S:=�=�0:�<V��F��#3��\���>/E׽� :��M�#nf�|j
?�/?�����̾�;׽麯�"��w<]?#� ?�⾤�4�35���kA�<���J��b�='~5��SE��w`�����g�l�A_��d�i{�=�#?�8�?�t�R1�V�㾎\*�.��G�h>��?���='Ѭ>��>�$�Mt��5T�8�h��v��I_"?���?K�>��E?e�X?�>p?b�Q?���>E��>!,�6�>p9>`ǯ>�U�>[EO?��(?'?�;?F�>?��*>m/<���ҾЏ�U�>ܓ3?��?ڐ?R$?b�����9�>r_���{Ͼ�����&E���3�j=��='�=(%_>0N?�{>�7�}3��]K>��?�p?���>�ܾ����>X�"?l��> #M=x;��|����$�c?���?����������=\�>�ż�h��
>T4��bb�=���=��O���U=)r,>z~v=����;����=�3+�{p�=�p�>s�?r��>E?�>�D���� �����a�=9�X>�S>.>�5پ����%��=�g��@y>�s�?�y�?�g=�6�=g��=�y���S��V��������<�?^@#?]RT?u��?��=?4h#??�>d(��P��F_��6����?�,?KZ�>���}�ʾ�娿�3�?�Z?�Pa����")�f�¾�ս�>%=/��~�����@D��+��t���白���?���?��>�U�6����WĘ�tL����C?�O�>َ�>U��>��)���g���_6;>��>JR?z�>Y?��?�j?��>��A��ﻤ�E�<B�}>hY6?Rx?7ߗ?�ap?���>��O>�#A��˾w���U�<A,�����i�7>�VI>�U�>m�	?���>a�{�:�q(_:�pо��=�cM>�>��>q\�>��>_=��G?��>�E���}�FǤ����Q�<��uu?ğ�?	�+?̮=�����E�i3���<�>�g�?R��?	6*?��S���=9wӼ�ﶾ@�q�'�>m̹>�+�>3��=bF=q>���>�n�>d��:`�=h8�9�M�S�?�	F?ꧻ=p~ȿ�J���٫��ξ'��=w��)/����ܽ�x�����<=P��i]ҽF�0��O^��*ǁ��ֱ�"���<�����>Yy����L>gj>�'�=Rw#>��=m
F�|�>��U>O����ܽr=i3 > N@��5��=�=<�>�w7>!�˾�}?�;I?�+?��C?9�y>;>b�3�V��><����@?dV>��P�����i�;�7���� ��L�ؾ"x׾��c�ʟ��H>_`I�2�>�83>�G�=~L�<%�=�s=�=R��=$�=�O�=qg�=���=��>YU>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�=��=ɹR�=0��PR�g��V����d?�C��Ͼ]j�>D	�=@�>ƾ�Ҋ=Z},>6Y�<��@��2^��'�=���$'�=ڗ=���>��>�(=oW7�K��=]��=T�*>Pn>^�`���e�*��tA<{I!>vx�>t'd>#r�>g?BW7?2�k?��>��:�<�þ<�ξ���>�	>H�>�})=�x>½>�1?�EF?2P?��>��j=�Ϸ>��>�/+�=m�HYؾJĘ�m�=�y�?���?���>�y��oO@�	���/��8��\7?xa,?L�?��>�	�R�心u)��5�[|���M�4�	4|��o�<�7S<�}q��_�<Y�=��>X;�>~ג>1ZR>>+5>���>�;>��=Ӊ�=hA��M_�<h`1<�M�=�y�=7!�=��F=#�-=��/>��=�9e�-]�=bگ��|�����=���=|��>]<>���>���=���XB/>ظ��B�L����=8G��F,B��4d�I~�/�sV6�<�B>�:X>R~��&4����?��Y>�l?>���?fAu?��>�!���վ�Q��Ce��TS��ɸ=�>��<��z;��Z`��M��{Ҿ���>$��>f��>'KI>�5'��g>�lԻIpϾt�.�2��>O�M�K4�=N����y�݊��Я���\�Bq�=7�O?˃���=V�z?41?��?Oo�>��7�%C�5��>gb�Q��Ĥ-���~�>dI��,?��G?��>=�
�R�\��O̾�)���ַ>�KI�a�O�����ϳ0�����з�{��>������о�&3�h�������B��Or�I�>ͰO?C�?N;b��T���QO�<�����up?Bvg?\�>�K?�??
��b{�p���J�=��n?#��?�<�?�>i�>�/B�Y,3?8�R?[D�?^�?�H?���q\�>��>O��<��J�ٖ�>�J�>7�=4��>:�.?��>���>{�ػ$t������3��)�� �=6{�=��s>ę�>�ͽ�)!�n�=e�>S��>�P�>~��>�C>��>}w>�Ъ�����+?��>�4�>g�1?�2A>qF��dܻ���=���`���z�����R"���<oN�<f�;=Xݻ��>����GЗ?���>@����a?B!�������>:��>;���nz�>�\>�z�>M��>J�>�UB>0SW>uܗ=E ܾ	�>n����"�h,?�s�Q���޾�u>^���/������ؽ3�[��򾾪{���e����Д;��>�;���?����b�Y@&�kҽ��?!�>�H,?�_��T�s�?n%>˨�>a*>�����Ɩ��A����ӾЌ?�t�?g;c> �>F�W?C�?ِ1��3�vZ�#�u��'A�[e���`�J፿省���
�D����_?��x?�xA?tR�<:z>)��?q�%�=ӏ��)�>g/�';��;<=,�>)*���`���Ӿ��þC8��HF>=�o?%�?HY?2TV�kl`�]&>:�;?IU3?��t?@2?F4:?M����$?ԡ;>�?@m
?�6?�.?��
?�	6>���=�啻.�=)	�� ����н�Ƚi�޼ �9=x$=��3;O�<�S=��<u�����Fo);���@o�<��/=Ѡ=���=|�>T�\?���>�8�>� 8?"����7��{���d/?�B=��O���j���G�\�>��j?���?��Y?+�c>��@��,?��8>���>��&>�j[>�n�>���F�p�=9�>C>x�=�8F��u����	�ґ����<�>�H�>�;>�Җ��PF>����֒��/�=��6��#������~#���/�0o�#��>g�E?��?�LF=U��-��Z�[�,�?2�8?҅C?F��?��%>��zO��,,����?��>�>��B����N��5C-�/ K<b�>5Z�'����c>	���޾*3n�'�I���澙P=����Q=P��#^־�A�P�=��	>����H!�=4��������I?��k=&����U�#!���>�/�>�߮>Ѓ7���{�I�@���먖=��>>t;>}k��Ti�KuG��w��_�>�{E?6�_?��?�%����r�A�C�p;�����������?�Ȭ>]C?�Z@>�.�=���������d��G�D)�>���>���H�G� ��������$�?��>8�?��>]^?UfR?�
?Y`?-�)?��?���>࠶�����
A&?h��?�˅=��ӽ��S���8�X F�r �>{�)?P�A�<t�>i�?N�?��&?�pQ?�?Z>� ��U@����>BC�>��W��g����^>�hJ?=r�>�"Y?�?��=>'�5�a7��u������='�>B�2?0>#?k�? ��>���>&z�����=�Z�>yWW?=y??�b? g>?a!+>�[�>��V=���>��>��?b�Q?��q?�L?���>�(;����ýHH��"� �{�<�3=��3=�@��9����c����<�v�< w������_�u?��/!��i8@��>�r>������.>��þ�J��C�C>����
�����:�=�0ѵ=匁>��?�B�>��$����=ʺ>���>���'?��?��?�;{'b���ھ�H���>�eA?5��=)�l�+q��nu��e=�Qn?LJ^?��Z��5���b?2�]?ɜ�=��þ��b��"���O?Y�
?=H��ѳ>7�~?��q?X��>�f�H0n�����Mb��j�G��=Q`�>�Z���d�p?�>ʍ7?�%�>�c>�z�=�f۾��w�������?`�?Q�?���?�A*>��n��/࿘��Y��1d?}��>�z���+/?ů��oƷ�ach��><����ۀ��୾�ي�ᆟ�^���$W;�N���&=b�?���?Tem?Eq?6}���Zk���N������H�_	��1��5I�ME�2�P���������]ͷ�Ż�=��f��r_��t�?�*?�M�Z�?�j��Hƽ��)��艈>�e���;V�oJ=%����=|��=�����53ž��?�
�>�C�>k?? ^�W�9�1�.�5�:�̯;�9>߯�>��z>�2�>��*�F���"��4�۾u𔾲ٕ�F�m>Y-k?Ly?�=�?N�=mB��џ�#��N��=��w�>���>Qj�>jC�to���"���5�I�W��y��S����	���=	?E<>�K�>�Ԡ?��>'���/9��R捾�������=�?6oB?���>~t�>Ǔܽ���@M�>88n?&O�>���>�>��ݔ#����+�Ƚ�[�>�I�>�K?� �>U�)�ױ\����L���
�9�Ǳ�=��d?+���v�b���>��M?Є
;Mɳ<���><t`��!�X�G�$��+>R�?1��=I�?>��ž
,
��x�����;�?���>r5��vY�Jk>_&?��>���>�ӓ?G��>\��� ����>�N?#�R?��B?��>�:A>�[H�� ��?8����=`�g>�`>N�K>��t=�IX��֥��&]�-r�=X��>RT>t��-̻Uؘ�^���r�z>!����ҁ�E
�s�M?˾�<��>i��N'�C�ƾRI�)_澺���  \�@ ���ڽ�xP�ȈM�P��c�x�-?@!��?"�̾3i,=�Q���%����о.T?	�� 9�3���'������!�xF�ۄO�L�]��ad�/���'?8�����ǿ,����:ܾ~ ?A ?��y?B���"�8�� >t[�<�'��מ�;���^�ο�����^?%��>�
�B��2��>Ǡ�>[�X>�?q>���3鞾�,�<��?χ-?���>�r�q�ɿ1�����<[��?��@�uA?��(������V=���>��	?��?>>1�:��ڰ�KB�>�;�?\��?ȞN=��W��
�ue?h�<��F���ܻ���=_��=x1=���|J>Y>�>fw��LA��3ܽ[{4>ʅ>�v"�\��[^�x=�<ӕ]>:�ս�=��8h�?@w_��U������=���<�>x�=?<ۇ=#�@=`�?AR �᾿�����:?Ţ�?���?f�B?������>a)��^;?�)?::�>�3�_a��3:P>����>Ǟݾ�J�=���!�>V*�=�ǡ���Ⱦ��M�k_��->n���YԿb)���-��R+=n�<�B��m.�9��N�����5	G��v����=N��=��Z>�v>F,>.�7>,�d?�d?�ו>��c>hʙ�����2��|�,<H���2��G@����z�*и����� ��1������
�%5Ǿ�=��=�8R�V���L� ���b�R�F���.?Kj$>��ʾ*�M���,<mʾ����w���饽@3̾��1�fn��˟?��A?Q�����V�]���f�����d�W?�J����PI��=?���*�=�!�>���=���� 3�~S��0?hH&?�ᚾ�Đ��1>K�����*=�C8?��?.v=2D�>�z
?ձB��ݽ'Ҙ>��z>h�>��>?]^=��~� �˓?��N?������2>�Tž�UU����<��=]E��x;�w>W����C��-rb�:��ox��eS?~ �>��+�����r�����?�=��r?P��>�J�> xh?w<?�J=���SpU��x��"<=��[?��l?f>j�[�T6Ͼd���5?E�_?��@>}f�g���B4�`��G?�1j?�?�押��y�Ǥ��.�KX;?~�v?b^�cZ�����8�W�vd�>.7�>`�>��9�v&�>�>?�"��A��Yѿ��4��Ş?��@�k�?��6<Ʉ�G�=�?q|�>�^O�7mžW���赾-�l=���>�x��Wv�� ���,��9?��?���>�낾�W��� >�<v�a>�?��?"Hþ@$$=�@3��s�9ͽ����=��<��=��B�̛�Մ2����V6��|��d*��>:h>��@���C(?P��Z濇*���5��u+���ޕ�y%?;�}>K�i���U�c�����B�m��Z>�9�1��;�>��>�ۖ�ؒ��|�^�9����%U�>����>�I�����eР�-�:^m�>v�>�K�>�z��߽��ԙ?������ο�������|sY?�?�*�?&M?�D�<�,v�_�}��􉼋cE?D"v?�[?��e�`��_&��)j?Se��xt`���4��!E�|^U>B^3?�`�>N�-��1z=��>#h�>��>�.�2hĿv��������?6��?-���>d��?��+?�{���������P*��+�9 S??�/>�¾�]!��=�%	��4x
?�/?'�����]�_?*�a�K�p���-���ƽ�ۡ> �0�f\��M�����Xe����@y����?N^�?i�?˵�� #�e6%?�>d����8ǾC�<���>�(�>*N>tH_���u>����:�i	>���?�~�?Nj?���������U>�}?)��>���?	�=��>��=)��Ol�P !>]�=m:�Ɯ?iN?:Q�>\��=�9���.�ZAF��R����CC�7��>�a?��K?��b>R^��v)�Kc ��mν~I0��J� @���"���׽�5>P�=>m�>s�C�N�Ҿq�?�t���ؿAm��x(���3?N�>c�?����s�����^?���>_��6���1����>��?,'�?	?�׾�μ�/>ʭ>p��>��ӽ�.�����4`8>!B?l�����
�o�b�>���?x�@Uɮ?��h�}� ?B�?b���s�z�#�H��ޛ
>��>*���|=�]3?F&>�i�9��k:T�"��>�7�?�]�?P��>MD�?|j��vo�aAG<�ف>7�?9{�>��a�o�4��	�>��*?r+�kE��zG)��^�?�@K�@��4?m;��egֿ'���7L������J��=Q��=!�2>��ٽ�m�=,�7=n9��?�����=��>�d>�q>�(O>�a;>�)>����!�Tq��ۢ����C���M���Z�2���Tv��y��3��(���,3��1ý~���Q�23&��*`�^>D�I?lof?�7�?-s.?�K�=�]�=�H��<��=�#B����=��>�BC?r�[?-K	?�~� �~�%V�{~x�ԛ�vϔ�6�(>�G'>��	?G�>���> L�=�
h>E3.>�m;> &>S�>��=<7��p��>��>5v�>�
�>}C<>��>ϴ�1���h�	w��̽� �?���0�J��0��!>��%���x�=P`.?�z>���w?п���%0H?����&�ɻ+��>��0?�`W?m�>�
����T��)>���e�j��b>�& ��yl�ы)��!Q>�h?"�6>Cv�>�6?��:�������#�>xW?h���"�L���O�86���,�>L��>�_��3N/�Oã��f�u�о����`?�b�>��+�b(Ѿ~��G�)�%��> 푽-�+���>&�W>��#�?`½�uh��&�=dQ�>ޗ>[	?a�d>䓰=�m�>/�����j�oT�>��>�#{>OD??�M?|q��]躽�����潵>�>Gz�>J/�>8Y�=
�Z�J�=���>`N>��3���������<�w>�B�����嚽F �=$�g�)��=�-�=M��DI,�p3�=�~?���(䈿��e���lD?U+?W �=F�F<��"�C ���H��F�?q�@m�?��	��V�C�?�@�?��V��=
}�>׫>�ξ�L��?��Ž3Ǣ�Δ	�4)#�jS�?��?��/�Xʋ�;l�n6>�^%?�Ӿ���>M�TG���X��=��w'��)h�>� ?}���Ǘ=�FZ���>p)�>�Ϳ�����Emɿ�QY���?���?��?ׁg�<f��?�H��b�>x��?VW?et,>�׾�j��ұ�>��+?A^Z?�N�>��ͽ�`h?�:�?�tT?9vt>�ۖ?�\�?]�$?�'�=۸E��ѿ��~��6>: �=F!�>���>1�ܾ�z�����U�m��eb�����s =l��s|�>�c���ݾ�ԅ>��3�6 ��I$>���>0[=�ւ>ro�>p�+?���>���>�cĽn�+��z9���D�W�K?���?���1n�J��<���=d�^��(?jC4?�4]���Ͼ�Ĩ>j�\?p?' [?�a�>��� @���忿
������<#�K>L+�>�C�>����>K>o�Ծ�D��_�>X��>Q���=7ھ�'��h���G@�>Ne!?���>���=Ǚ ?Ü#?'�j>)�>aE��9����E�7��>���>�H?�~?��?�Թ��Z3�����桿��[��:N>��x?�U?�ʕ>?���σ��w]E�lDI����K��?\tg?WT�+?,2�?�??-�A?�)f>1��Dؾ������>�?�4Ӻ�	a�jh�8w��
b�>��"?�=�>�q��ҋ��2o=�'��žf�?|�?�:�>kA7�A���y0Z��%H��O�=�B�<��m��O�s�<>��<�P�18>W�w=l���������}�rR�=W�F>q��>��!>V%������-?9+����p����=J����"��H�>@:߽Jn��-U?�JW�����,���a����d�"��?Z`�?��r?�=<ᆿ2�T?1��?�k>?�_G�-|ξ�Ѿ?E=��#˽LhȾG7>��>rm�(��%��.��ʅ��%������>��>$�	?O- ?T�K>N�>}
��J�'��J��`���u^�����_6��.����p�����-���ż���B�v��o�>�N�����>� 	?�f>��y>6��>5���O��>�P>�Bx>Ĩ>[!X>�B7>z� >`�<�� �/?厸�Q�?�����t����#?a�r?8��>jh��x�aX�&��>�y�?Y��?,�p=6�z���I��^�>3O?i ���f�>Z���3 �=�E�= ���(�0�`R=��=��=�j�����8��Ę�v��>��?YV��Q�)�5z�����2�s=�C�?
�)?�)���Q���o���W�k�R�]��WKg�A>���%�G�p�я�q6������L�(�^�)=�)*?t5�?y�#��o���uek�{�?��8e>���>��>ְ�>5�H>��	���1���]�R\'�
h��q(�>��z?�s�>�,.?�1;?Q�4?F�F?J[�>0 c>��E��� ?�,=Jw>�~�>�q(?̆+?p�5?��?�x?B�>�+n�K8��	�龽��>�?��?���>�g�>Y���M^�O���[=�qܼ���=�&>�]~���D����<��;>�F�>^���u�E5�+)���D�>7�>?˝y>�`9�S
[�T/:u�$�r�2?b��>:�G�່�F+��f?U�?X�jܐ=0��<_ �=Z[>#+a=dC�=C�=�=�,��� �^��=x�<���=�;> .>�\$�w�����S=�u�>��?���>�C�>A@��;� ����7n�=Y>�S>�>Fپ�}���$��*�g�O_y>�w�?�z�?�f=��=��=�{���T�����M���*�<�?0K#?�WT?Ǖ�?��=?j#?��>�*��L��r^������?L�?=��>�7���ʾ�9��U;��,?�?��D�l�ݾ��K�|����e��=&�X�j�����?��?� ���_�77�?(��?�T���.��|��٠�g���K�1?�}�>���>~��>��1�<�n�d���q>�(?��S?$߶>ʷO?�(�?d�k?Sˁ>��%��)���;��I�*<W >�~9?[�?��?ѱu?��>!��=n"*��.޾�V �buO�h]�Ot��S�e=���>�˥>D��>;̣>�k=^q�����)� �y��=�Ȏ>�7�>���>�4�>�w]>$7r�PVN?,l'?mX�Tr���c��Â�����=.�?�@�?#	3?�
;6��[28�֓��6�?<��?&�?˚A?���:���=��W��[��V�k>py>#�>;A=�5D>/k>�>,w>������
���@=��>��#?�m>��Ŀ�_q���v�5ɚ�.��;���{�\�΢���b�ޮ=�����v������W�@I��/��?a���_����u�[^�>�{=~��=?a�=���<�c���D�<��E=I,|<Mu=?q���l<'�#�;����·�ݗ�vO<�U=Ɉ�G3���wt?��`?�O?n[7?�AJ>L�"�b��Z�>�@�<7?��>��'=*~��38?�q,���J��h�پ�Ӿ�u�G0��`�'>�wH=d�7>��A>��w>0���_=��=oG�<��.�X�>�S>�ޕ=X}�=�9>�(>(�>��y?.Ow�U���I�1��^��-,W?��z>ҁ�2��".4?/b�>9�S���ſ��=���?)o�?�k�?Yz�>���+�>V����l/��[k>��A��>$��=�.����>H\�>�E�zt��gd׾-�?P�@7�]?�{�g2���>�&6>�@>�'T�Ms1��4X�M�e���I�>'!??�;�m;���>U~�=��۾ǌ��R�=�</>�� =9$�QX�g�=��d�q>=�T=��>R�D>r��=�[�����=�K=�	�=�/J>���@�d���@=΄�=H�[>�>A ?�? �&?�:?��?Y����A侸��P�>;c�>H�=V�7>�E�>�t�>9�)?*�(?�X]?�>������>o��>d0w��:����9���w��=��?s�X?�>-H�=
�8�j�qtI���>��,?/2?�x?�P0>�X�h]꿗�(�5=��$��k�;�=��$���kp��i"�\�o�YA
>���>g�>t�>3hS>ž	>dX/>G�>��	>۬���=5=�:�<u��;Zy=j�
��E�=l������]�m���ޫ����<�Gf=��'<+hӼ�u�=; ?!Q6>Ggl>:d�����O)>۽��^�+��+>QZ���?�V��3ߒ�����+D��g>�qP=�ƹ�u��f#?J-�>��<�X�?�g}?�*=����>��	ʖ��n��>�;z,�=՗:>�l���X��Xc��m6��C����>E��>���>��g>��*��E>�Q��=�����5����>�����9��{�o�}򤿠����i��뺺��F?�̇�b�=��{?5=I?D��?h`�>��
�վ3=1>�������<NC��p�����ie?%�'?�g�>Bd�_D��^��r�_H>1���HK����Y����߼����*�=���7?��
���j��9���%V�p����=�>V[^?3J�?٨��y�:�n�k��WV�0~U>!�?(g�>|���JK?D S?�X1�����ť���ɾ;�9?27�?\��?���N	�=m��\Y�>n?�ϙ?�ב?��l?c�1����>M��<>�>Y�(�D�>z�$>���=��=��
?�H?B�?�����և������9p�=�<�7l=�+�>#w�>�Y�>mr�=K,0= ��=�:X>�4�>���>�o>��>� }>�m���6	��S-?�4=igu>��X?��=�޼��5�ճ�=���<SE���ʾ^��>�U#>ҫ&>2����WK���>L���?��>_��jK�>�zA��^�>��>T�>�F���"1?P* ?[�?��X>���=�ٷ>?��>I�3=��,���=�H&�u8��i��`���2H�>���Nm�����<�{�{?ٽ1���� 3���l����j)H�8�h>�<�?+L}���.�3��ޯ��L�>"��>�!?�'�����W#>���>��>qn�`���^ҏ������?*&�?�;c>��>@�W?�?��1�3� vZ��u�V(A�e�U�`�}፿����
���'�_?�x?,yA?�P�<2:z>N��? �%�lӏ��)�>�/�';��@<=s+�>(*����`���Ӿ��þ:8�(IF>��o?7%�?yY?<TV��T=�=>��D?n�E?wҍ?f~C?
?��E���=?�K^>QȺ>i�'?G>N?˵L?~0�>��>>��>3P�<ps��a��w���W�^�����=JI6�T�=3��=���>J�ż80 ��_�<��n=��	�6����<�� >�0�=�Ų>�\?Rj�>�j>@-+?��#�>�&�a�n�j�A?�w�=�z��p���՚�ZL�i�E> �m?�̨?��]?�'>�\��V�>F+q>a�">��h>臛>�3�	{Y���5=���=�7>�B�=nܼpz�������jn9&�>���>�#>�����#>�Σ���x���e>��M����%�Q�1�F��1���y���>�5L?��?�=5��}�f��'?�4<?:L?f�?@��=�?߾��9�_�I��=�ؠ>��<� ��衿ܜ���];�|�/�e�q>-�� ����-b> �� n޾�n�{�I����/�L=�{��}W=t�#�վ�B��>�=m
>������ ��
���Ҫ��,J?!j=@c���U��p����>��>���>��:�_(v��y@��׬���=O��>��:>�z����mG�,4� �t>�pK?�Bd?��?j�\��t��.E��M��������Fl?�G�>�?�D>�=�R������k��&J���>g��>����l9���������-��К�>,�?m�=d	?s�M?L�?�a?�!?� ?߼�>�/?�:��^B&?І�?/��=��ԽV�T���8��F�� �>{)?��B����>��?�?��&?Z�Q?,�?��>�� ��@@����>AX�>��W��_��
`>��J?��>�5Y?�у?M>>�5�(⢾���=2�=<9>c�2?�5#?:�?�>���>u���C{=�{�>��a?��?�6o?˓�=)�?�J->fF�>]8�=G�>z��>L�?a�O?�s?�hJ?��>~�<Ƣ���Я��>}��Q9����;��&<[<T=�H�9�?��y"���<rJW��ͼ��C�b��h�K�N���^G<��>?j>f{����>�ʾ���,J>�PV�ˡ�&m��r2�4�=�p�>9��>v�>�h:�ⅅ=Ɗ�>p}�>�3���%?�C�>�D
?���<�X�8!��{���Ř>ـ0?>o�\��}��C�q�|ũ=� v?;�h?,�^�4m�s�b?��]?)_�`=���þ�b��c�!�O?A�
?��G��۳>��~?D�q?g��>!f��;n�����"b��j����=�x�>_O���d��U�>�7?2u�>�@c>�M�=�۾�w��<��Y�?b�?���?� �?��*>$�n��2�#l���뇿��j?&>�>O�þf�.?Y���kǽ���:�.���#��{��Ć������&���p��솾��	�"��<��?W�?,>n?->z?����N�v���J�N*��~F�c��/��!J�	<I���D�Xpt�p�,"��Ҿ��=�肾��=�S�?Ft?S�m�!
?�,���پ����F>hKԾu̽A��<���
��=�2�=�x_���6�l����*?�v�>{s�>�F?�Y���A�{;&��g:�H��/>dA�>Z�j>���>�G����I�`��4�ؾ�w���u���bc>�ul?3�R?��u?�4+�C{��G�#�reS<vv���?>@�/>g�p>*�o��{%��$��g?�&�z��2#��X�	��4�=D�-?V��>Z�>�Ò?n+?�� �6����Lw��('��=�Ƹ>�Ye?�M�>|>Ԟ�������>Y�l?���>�a�>a���D!��|���˽�k�>8w�>B��>�Sp>?�,�g'\�Na��0z���9���=��h?���za���>,�Q?^��:�tN<�Z�>��u�c�!�%�^�'��">s�?���=�;>�lžk���{�O@��B�)?{�?3)��	�*�n/~>��"?�	�>���>Ϡ�?|ҝ>C�����Q���?�_?\	K?N�A?�1�>��=#��RŽ��'��M-=�+�>�Z>��q=���=.L�I�[����<5I=�J�=�u�d䮽{0<���D�X<�3�<�H0>�eۿ?K�j�پ���C
������񱽣z��֋�F��E����.x������'��6V��c������l�4��?�0�?*m���8����������B���\��>Mq�!�~� �����핾n��R����i!�2
P�*i��e��Y'?�����ǿ����2oܾ��?�G ?�y?;��("��e8��6 >a��<����z�����7�οf���0_?��>� �9]����>En�>��X>z�n>�܈���3�<Rn?A-?���>�q�]ɿ�w�����<��?��@f�@?�Z!����Y:�<f��>!C?*BQ>r����S,��y�>�×?��?��J=��T��e���^?V��<�1A��'�;80�=���=s�<��½r�V>���>�ӽ`_���A�n>u�>ί��d)��x+����=���>��2,�'��?	�A�	b(�ՅҾG�Z���e>��6?l���J��==kN?	f���ڿ�񁿍��?���?���?;+?��Ⱦ��=՗ž
�L?8Z"?���>�()��/��cʚ>y�>>��>�뾝'���t�>I+�>�I�h�s�s琾C ���2k��[�>����ƿ�|%����-�=-G��ՒK��L�5���`5T�������k�����T=C��=��R>f��>��Z>'_X>��V?=Jk?���>2v>��eA����̾��5��L���F��@���أ���쾖�޾����+�����Ⱦ�=���=�"R������� ���b��DF���.?��#>1�ʾ��M�x+<� ʾ�ª��Ԉ�������˾�]1�5�m����?U�A?߅���V����F�丽ݪW?�����Zm��"�=$j����=��>���=up⾲�2�
mS�]1?=A?���^����*>b#ٽk4=Q�(?���>WyK<���>��"?�� �{���c>F�G>�%�>h;�>�_
>����Z!׽G�?�N?� ��:���FՋ>Oeʾ?�l���=�=��.�R.r��9V>���=mu��(Ƽ�v���>=��,?�|>a�%�I`)�)����i��2@>�Ht?L��>g��>
]M?�"$?��L>�ʾI*M�:� ��r��ee?��m?T>��ب�'Bf���
?��S?����辧SU��T�' ��;�>U�{?��?w�3�?�{��^���Y��(a?1/K?L�h�闟�}h������->*<?�>��=�kd�>2�0?.W��ݵ������<�/�?��@ŵ�?Y��}:�~>H�?r�>����Nþ Y��������;�?�T��E {��S#�˥D���(?�*q?L��>��X� S���E=g��ɰ?��?�ݾ����n�)�:%f����"�z���Ľ"�~�f�0�p���(��x��~���>Ӿ�ɽ�^�>��@����S$?B4I�� 뿸����Ĉ��žĶ��v.?�>cS�7�¾��{��-n�[V=�!^��(>��t�>�/>
 ��������{���:��Ӑ��>�\��c�>1�R�o뵾v����4<��>�T�>|�>{���RG�����?�o��G�Ϳ1s��d��ZX?9�?zH�?4�?�"<(�s�g�y�͉(��zF?Pss?S[Z?����]�Z�>�B�j?�]���Q`�4�4��IE��U> 3?�;�>^�-��|=|>|�>�>�/��Ŀ�ض�(������?���?�e�4��>x}�?Aj+?�b�5���H��\�*��E�|2A?].2>G����!��-=�˒��
?��0?({�34��_?�a�c�p�.�-���ƽޡ>�0��k\�Pa�����Ve�~���Cy�$��?M^�?H�?��� #��4%?#�>U����8Ǿn#�<��>W'�>k*N>�P_�e�u>����:�pd	>m��?n~�?j?{���<����T>�}?��>��?���=��>|6�=����N4���#>�A�=p>���?^�M?�H�>�n�=H�8��/��UF�YaR�j4�ĠC���>%�a?b�L?�b>�˹��z0��� ��ZͽJ�1�F-鼘5@��H+�c�޽�4>��=>=->�HD�"Ӿ{t?k�&�� ׿��͞�A;?�Y�>��?ȋ�+$�����=�Y?��>���}��Pw��x����G�?I~�?�� ?:�Ѿ��`�ƥ�=r�>�h{>��X���p������>��9?�穽 ����d�a|>Q�?!�@�?�_��?pW�hS���H~����7�j�=��7?���x>n�>v;�=��u�ꍪ�O�s��{�>4�?pI�?��>Cwl?�o��qB���-=<]�>Q/k?�2?^֍�i��$C>we?��Fێ�lh�@�e?�
@�M@ `^?����������{��}Ҿ\�r�=a��B$I>�b�=��;~�m�W>�C�=�ř>%�>ǽ�=L��=M>/P>��(>��{������ֿ2����@L��5����[���xi�ԹP�kB���k�]+Ǿo�0��K��,5y����<]��=�-F=��j=x�a?�^?�X�?��?X����=��ܾ��>7vٽ���=��>;2.?;A?�"?��p=���5Ku�����y��s�l�>h�>�Q�>#�>��>��v=:PA>�J�=���>�O�=���= �=K�;�4D>Z~�>� ?g��>�C<>��>Eϴ��1��j�h��
w�U̽1�?����P�J��1���9��Ц���h�=Eb.?	|>���?пd����2H?%���x)���+���>|�0?�cW?�>��T�T�1:>;����j�5`>�+ ��l���)��%Q>xl?��f>�u>�3�@e8���P��w��'j|>�46?�趾r;9�K�u���H��`ݾ�GM>�¾>D�Ai�.������li���{=�x:?��?�N���ా�u��E���VR>x?\>5>=XY�=�`M>�^c���ƽH��.=��=��^>��?��&>�J=��l>b|������#�>&�G>���=n/5?�Q%? ���,�	h���1����>H��>�L�>�L>��gn�=���>"�1>�>8�r��>��^A��B~p>qa�=#�m��.[�6�m�(&���^�>}�>]�4���E��~�=�~?���&䈿��4e���lD?Q+?P �=ɝF<��"�D ���H��F�?p�@m�?��	��V�A�?�@�?	��Y��=
}�>�֫>�ξ�L��?��Ž<Ǣ�ɔ	�)#�gS�?��?��/�Wʋ�6l��6>�^%?�Ӿ���>´��혿������u���=���>n�H?���@;��];��	?��?��n?����ȿ��u�@��>�_�?/��?�l��E��S?�ڢ�>���?�iV?�[a>��׾4X���>�z>?��R?rͶ>�4���*��?�k�? �?i>>0s�?��?܀2?����V7�A]��/�����>#�ݽ�->��m>M-�DfP��%���f��(`��H�k�=��v=Oѳ>"��(��'0�>F:�=�оYsu����>?4�=[�>��>��?>�>��>=墽҂ѽE���p-p���K?���?$���2n��N�<Ġ�=��^��&?tI4?�k[�S�Ͼ�ը>ۺ\?e?�[?d�>.��D>��?迿!~��ɩ�<z�K>4�>�H�>o$���FK>��Ծ�4D�Sp�>З>�����?ھ�,���J��bB�>�e!?���>Ү=̙ ?��#?Tnj>���>"eE�P-��*�E�X��>��>>;?�~?��?0���sE3���桿׋[��gN>��x?�Q?Xӕ>�������5�A��GI�`��R��?8Jg?�潯?n/�?�j??͎A?�9f>��2�׾6̭����>"�I?ݎ1�mZ
��%����N?e�>�b=5"R���G>��m>-�;�#�
*<?��?B?�堾}�6��	����=[	������:>V�=��X>	g�<m6�����<mY>�>S�txԾ}��>�G>�dE>�[>��l�勛�W>,?��F�(Ѓ���=_�r��zD���>�,L>`���|�^?��=���{�A���s��8�T���?o��?�`�?�̴�z�h�r,=?V�?��?�"�>;A��{޾�t��w��Xx��|��>���>�p�R!�Ύ�������J��z�Ž�SV��?Iy�>�1?� ?|�s>���>3,���T����� �5`���#���A��!!��	��˦�i�j���}��[ܾ�r���>\�T3�>��?L�>:y�>>m�>�R�B��>��Y>K��>�W�>
 >���=G�=�>��Q��3P?���RQ#��B�r�����:?�^?�g�>d����΀�˕�3?���?�=�?�L>��j��(���?&!�>��c���	?3=b},�B�A=.z��_���t�һC����tT>|yռt�(�11M��rm���	?�M?=Q�ʾ��1��⟾D�=ދ�?�0?$�.�)T���r��X�D�J���?���r�����_Y)�#p�ӄ��΃���"����,�Q!=	�)?���?���u���P�k��>��-[>���>�n�>���>�U>c���0�C�_���'�@߁����>��x?��>>�I?=<?GuP?�jL?0��>�c�>�4���i�>���;��>P�>��9?�-?-90?�{?yt+?u3c>��O ���ؾ�
?��?RJ?l?I�?�ᅾ�qý�7����f�A�y�O��� �=Kz�<`�׽kGu���T=9T>.k�>q[��d�"��S���z��?�]d>
��=;�N�����yѝ�k�Q=��K?+��>��󰐿9im�\?uפ?��=�f�=�>�d=������=�a�=�uJ��΀<�߃�7�㼐���ñ=�Vl=�-�<�8=�r�=KTj�*U��k�>��?Z��>
:�>�;��Ϋ ����데=��X>� S>=>?پA{��'#��&�g�kVy>�w�?�y�?)�f=;#�=G��=�w���R���������<��<�?	I#?�VT?��?Z�=?�l#?	�>�'�dM���_��u��S�?�,?肑>���s�ʾ�𨿺�3���?C^?�;a�b���6)�f�¾��Խ�>�[/�p/~���D�T	�����#�����?$��?dEA���6�t�������L��p�C?K�>K�>T#�>��)���g�'��;>ӏ�>�R?6�>�ZP?�{?n\?�uV>|�8��"���X�� ���{�">�D@?/Ɓ?ο�?��x?D�>�,>��*�Ĝ���q��4��n��:�`=�%[>�6�>��>���>Ռ�=�cͽ�ί��@>��k�=�=d>��>�G�>���>K�y>��<��G?3��>y4��(��G��.؂��}9��Pu?�7�?"+?��=�;�CtE��{��.T�>�\�?�ث?�*?�PS����=��ռ.��v%r����>?�>Ę>6-�=�=H=�,><��>�j�>UH��C��17�QLA�e�?D�E?�q�=a����Az���ɾZu���">4�ɾ� w��=������4�\�����o�6z���jϾ?���Jo�w��-=T�d�>�yB=ׯ�=<4�<�r>�n;�=���;�u&=HD=Z�Ƚ��J=;����?�uYS��t�=�ǰ=���=�n�y����:�?�Og?�IL?�%Z?��#>��|2H�"�>�W���>���>�=��˾��(�����7	������R��"<��F���ؗ=6����>�g�=�B_>*A>8��;z�y>�F�=��=�	>t.�=`->��=��>SJ>?{�=�z?�d����FW���ýќA?׼�>���:��;��I?�e>h�h��㩿��ݎ�?���?�޽?�m�>~>���>�o���C1<u�=���Qk>��O=H٠����>�!�>����Ք���~�e��?8@# 4?���Ko¿`Ѩ=����*��rb���D���N>[�Ҿ.U�>wJP?�ya�T/߾AP�>���>���U�lH����	>f+?4!\>Y��Ö>!�<��>��= �.>�=�>E�>8p=,�E=h��=�
�=�`>CQ�=��<�P>��=ir��c>�>���>`�?t-0?}�c?m�>�,m���ξ����eҋ>���=Lv�>��=l�B> �>v�7?��D?V�K?O��>w��=�
�>u��>n],�Ǚm���Qy���3�<t]�?#��?P�>'`P<A����[>��9��Z�?�-1?�1?���>T����]&�l�.��B������i+=�Nr�0�U������R��n�Y�=Nf�>���>r�>Tmy>�9>��N> �>G�>)t�<�^�=�A��+��<�(��
��=�c���h�<+�żܣ��ɱ&���+�G~��f5�;`�;|^<%��;���=,E�>\�!>Br�>��=J����@(>�Ǚ�c�>���	>$G��M�C��g��I��'����"u5>�t+>�h��m���W?�IH>$�>���?dy?V�=�ݽ�MҾ�f��'�7�ȆX���=��=�ua�	A��_�-�B�;�8�>��>�t�>w�j>�%,���>� fz=ԗ�|K5��N�>�g��@� �T����p�����響n�h�z���bD?4.�=ڑ}?,�H?͏?u>�>�ѓ���־+�->�u��d=�X�[r��Ք���?>�'?�:�>쾋.E�ۡϾ��ͽ�D�>�K�_/P�>ݕ�q�-�����Y�����>�%���Ͼ�`0�����@) C�mZl���>�N?KL�?Q�j��v��£P�S1������?��f?��>p�?��?!���]	�W쀾Ͱ�=�m?Jp�?Я�??n
>5��=�ٱ�'��>ì?��?�n�?W�r?�O;�C#�>���8F�%>-��<C�=�b><��=[��=��?!}
?�	?G���[�����]��Qh[�ۂ=��=ƌ>�>�~>���=�`i=a�=�EW>n��>�u�>��`>K��>�Z�>�-�	����$%?�x#=q��>�J?:�=�8>���= ��4��	��Ɣ��'���2�<r��=u;bf��U�;�>}�ʿ�?nl�=��A�iZ ?���ZY�<�^=��=�X���\?��>>�>�D�>��>h�A>q?a��=�(Ծ�w>uS��!�p�B���R���ɾ��>����Yh����P,�;�A����)��]�i�������9����<���?b� ��di���)��/���?�7�>3?	懾�p�>�?�>]ޓ>Y���Y0��c���-��:�?aH�?�<c>��>��W?j�?W�1��3�MuZ�x�u�<(A��e���`�0፿�����
������_?��x?�xA?�Q�<�:z>��?e�%�;ӏ��)�>_/��&;��:<=�*�>�(����`�H�Ӿ��þ�8��KF>�o?	%�?�X?�SV�F�m��'>��:?ћ1?�Ot?��1?a�;?�����$?^o3>�F?�q?7N5?��.?$�
?B2>�	�=y
����'=�6���O�ѽc~ʽ���!�3=@_{=͸� <��=���<H���ټ��;�%��6%�<3:=��=�=>�w]?���>�2�>9�7?�C��18�vx����.?��:=s�������Z5�L�>5�j?j�?.dZ?�d>��A���B��<>�s�>;&>�/\>I��>�F���E��އ=��>�n>���=��J�����4�	�����v��<�>4l�>���>�=�<��v>pΠ��ۓ�e�}>�6����Ͻ.��<��f���0��˾��>�W?��<?��T=�����/=�1��ڋF?��?/,?�
�?(T>t	�]���J�&Ut�$7�>,Wp<��ξY��l!��e�U��i�%H�=p���x��~�4>[x���Ӿ�Us�dL�|�ݾ`�<��/�9�=�7����I��f��==k�=�����:��˓� ;��|�B?�ʉ<$X��QĀ�]�;̀>�ƅ>�7�>�*�<�ю��X.�c��#�=r>�>�G>�JJ�����@��x
��}>WE?�@d?'�?�ɛ�d[��Z?��.޾�&c�4�R�z?���>�L�>�P,>}��=S�;c`�u�m� rG�O��>I	�>���)O��ѡ�*���9��	�>�Q�>�Z2>�9?@,V? �?v�Z?�K?��>�I|>yW�`G��)9&?���?C?�=σԽ�T��9��(F���>�)?C�ج�>�z?ɑ?��&?��Q?��?��>� �3@��~�>�Y�>��W��j���`>O�J?���>�EY?�Ƀ?� >>)w5�٫��������=��>]�2?�/#?a�?��>p��>�9��+h��3ۚ>ҶY?��n?]P?S���~�>�TQ>X��>֝�=���>���>);�>(S?rxw?LaH?�k�>��<�L_�M���<�I:�}�<ød����=�/ʽI�O��Z!=ZX=�Oq<�6���nD����������=����#�>Y�t>(_��۟3>fƾ�����:>~�f���kz����@�%��=�~>�B?���>W"�uh�=ą�>-�>���F�)?�>?�p?���;�c��۾�2J�c��>��@?wF�=��l�ڗ����t��h=�n?9_?��O��x��8�b?��]?�g��=�7�þֵb����i�O?^�
?h�G���>��~?D�q?2��> �e�9:n�'��Db�,�j��ж=Gr�>=X�l�d�R?�>V�7?�N�>[�b>�$�=Bu۾��w�|q��{?|�?�?���?�**>|�n�C4���޾:��ʇc?fW�>`����4?����z�Ǿ<5�1i̾_�
��5����1[�����O?��N�����r:>3D?��q?k5j?B�]?��%Ut��]�+]��_M�+������VA���?��1���i�vtӾ�إ�����/>��n��l;�5�?�D!?ҰQ�49�>������xO��e>�X�������=��[�SX=�k	=@����+U����`�?7�>f��>.H5?D�]��I�
6�op<�[����b>F��>�ϒ>���>Zd�<�>���������N�!���6n*>1iq?s�n?�M�?g�˾��Q������D�=Y���(��>i��>�u>E�6�;h���=���?�-�~��R0�"6��������<$��>�t�>��?"�?Ph&?4���튾&o���r �	�=��>2?f?��>�>����h4�>@�~?i�?���>������!�sR��ߍ�b��>��>��>}w�>�2��k�G�MƂ�W7���h���=XTC?@���!���|�>�5p?ȃT�z��=[�_>�=*�_J�n󀾬)��Kz�<�'?�@�;->�I�`��a���)��R')?(w?9����*���{>P!?%��>o�>��?� �>&Y¾�J��%�?��]?�4J?5�A?�T�>��=0-����Ƚ$}&�ٲ/=>��[>&]v=�T�=�-�\�#��'�E=�k�=(+˼Վ����-<�����[<�	�<�,3>k���&*�a����.�����ɭ���Ӿj��ԧ���+5�K���6�#����lږ��A�b�K� e���̔�p���@��?;��?[Q"�Ě�W%���>���}�k�>�Iξ'�">�(��1�������WҾ�@�d�E��6)���֔'?���ܽǿް���;ܾ�  ?�A ?�y?��"�w�8�:� >�J�<�+���뾐�����ο�����^?y��>��*3��I��>6��>��X>�Jq>����螾�:�<��?��-?��>D�r�3�ɿX���q̤<���?�@�4?�.�*��saJ=`��>��>nA�>��/���$�rE��(�?�'�?�*s?���W�r��b(�n?ܓ�>�Q���B;�N�=g��<D���,��f�=>4i�>mU���q"��;��g>�5R>��m��3b�� ���ƛ�n�^>e���qvҽ�҄?dv\��f���/�yK��]>\�T?e��>��=�,? H�OtϿ��\��a?,�?���?�(?ɿ��ʚ>��ܾ�pM?s<6?��>�I&��t�n�=�6֥�P�㾙V����=��>/�>]h,�-��AtO���� ��=]�����ÿ,���&�3��<���oK<��*�T	
�<�#=�3���$v�'�ս�"�;�ܬ=4�>�a�>R�<>���>��S?^�a?��>��">���\p��&�Ѿ�����m��x�R�p��J��ɮ��tʾ�4������.)�w��i	Ծ^�=��=LR�)���rs �܂b��F�n.?��#>vʾsM��8<[�ɾ{��6΄��Q��!̾o�1�� n���?:�A?�����V��0�RL�����mW?Ua�qB��~����=�	��=�˜>Ă�=
㾆�2�2*S�� *?g� ?$쩾�Ճ�'N&>Ș�S�f<y$?���>t�H�VŔ>��?�Q������ w>��:>��>k��>&�>�
������
�?��e?�O���Qx� �v>'�Ѿ|E��e�=;�>ȉ:��S;���>=�=.<��;������u*����S?Ӭz>�.+�QX�B����g>�=*+y?Q�>HK�>ggp?�>?@��<���;Y�v�	�u*�=}�`?�bY?�[
>P/}��M۾5���kP2?�a?|�T>hPX��6�X5�ce �e?��f?m ?}P �/=��5<������.?��T?�@R����1�WD���H>���>��>s[L��W�>i�)?S���w��е���H��f�?�y�?>��?�{ ��=���=�L�>��'>�5�T�������A��P>��?v?��n�j�_!��\��_'z?b��?�%�>���e�1���=������?�u�?�о�TŻ%����?��겾��=�wt�=��=���T~�Q	2�*����D�2��o����O>��@�W=;���>���B�rο�熿����W�8B*?K�>���t���L�n�IY�r�8���9��������>�s�=N���ۉ��I�w���<��d����>�(J��;�>exW��W��r��������L�>��>1��>������jȗ?�F��p̿�ٜ��#���Y?R��?�ʀ?}!?�j=Cm|�w�t�
N���^D?�Cs?-�\?�^a��lq���!�j?�_��yU`��4�lHE��U>�"3?�B�>V�-�?�|=�>���>g>�#/�y�Ŀ�ٶ����[��?ډ�?�o���>l��?gs+?�i�8���[����*��+��<A?�2>���I�!�F0=�=Ғ�˼
?M~0?"{�\.�"�{?�cg��qm�.�k|G>���>��˽�I��sHG�j����b!������I��J�?m��?�U�?PW��z���>F[�>�f���*���i�#��>���>��>�=�/�>����"I����U�?ω�?��>C��������)=Z&i?}��>9>�?]r>CF?8�U=��������J>�>>�낽�g�>�S?��>��^=�i]��
B�9�G��3\�(��"�<�R,�>v�\?kI?t�{>�c&��	�|v(��1�C���Cw=>�ٽǝ#<�~Ž�T�=�W>��==IO��Dھ���>Q�#�5�ѿ�]��
�����>���>b#	?گ�B���r�=:?xg�>���U���e놿N�ս��?�U�?�]	?�亾ۧ����p=c��>M#9>�p[;\QZ�pT��m�>��9?���^�2t�d%A>�T�?��	@�ԡ?�6c����>�g�ԇ�%􀿓�
�絾	D�>��1?n=��ߛ>���>�<�^\�q���dI��ô>Y۱?7%�?���>�Y?dd`��/��n3��S�>�;\?-�>{{.���վ�q>v8�>����$����F�c�f?�@Gr@�-'?0��-�ֿ�霿�5��h���Q��=U~�=|2>��ڽ9�=��6=,K8�U���)�=��>,�d>)�p>'O>7;>�=)>'����!��v�������D��Xn��Z�D��;�u��n�G:�����K9��JhýV���;Q��7&�U�_�L9�=�-V?K5W?/�q?x�?�P�΃>~%��h=jo�� �=x�>M�1?U�G?��$?�D=q����f�i����`��:��~�>'�G>�>�>ER�>7(�>0=�5P>?>�Mw>��=J|J=>s�e4Z=��N>�ƫ>���>��>�C<>��>Fϴ��1��j�h��
w�o̽1�?���S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?'���y)��+���>}�0?�cW?�>��y�T�4:>8����j�5`>�+ �~l���)��%Q>vl?y�f>�s>�f3�[K8��P�����|>��4?(����6��u��H�cNݾg�K>P�>���=��͖�Js~��h��{=B:?��?�N��4:��V�v�H�����R>n][>��=h�=��L>�[]��Žd�H�_(=\��=��Z>�`�>g�>���N��~�S����?�����>�é��!�K�v?�)?VD��߲4�Zj����[�.?��?,�.>A,|>C�Q����=8��>���>��B=�tP=�2s�A&�9�=Aa���ǽXNQ�=|`���9{=�l]���h�"�z���`ڌ?*;��U(z��Ӿn1Ľ�6T?u�?%�'>��>:lξ�A���(���?��@�_�?)����v��+�>��?~�O���J>��?(.H=�<�s!]�~*?n8l<������$��o��O�?�8�?,�6��Z�'�G�鰁:ѳ�>�iнV	�>�I�^W��
���v��}=Kq�>6�G?���5�M�ܸ<��v	?�^?�u�Φ��}ȿ,v�F��>��?.A�?�5m��h���]?�cm�>Q�?KZ?0l>�ܾc�U����>�??csQ?;�>���*���?���?Z]�?|�>��?�}�?�?����}%�����m�m���3>Ӭϻ�L�>2��>��3�8�1���ŏ���l���5����<u�<W\�>)�U�*굾	�=i�M����"���+�>�'�>F�l>T��>��>�%�>��x>�=����P�{�����w�K?���?���2n��L�<���=-�^��&?�I4?�l[�{�Ͼ�ը>ܺ\?c?�[?�c�>D��S>��B迿9~�����<��K>4�>�H�>�%���FK>��ԾB5D�zp�>З>����?ھ�,���W��?B�>�e!?���>xҮ=9� ?Y�#?�j>>4�>bE��3����E����>��>YB?�~?��?�ٹ�AY3�1��/硿^�[��N>��x?KS?��>��������HG���H�YȒ�ڛ�?�tg?�R�?X2�?��??o�A?&f>���?	ؾ�խ���>(�?R s�K�K�@~(���]��/�>�a?��*>.�
��ۢ=��E<���������>ΘV?��@?�F˾�eC��$��	_O=��P�͐�<n�<!G�< <r>�>����h�=<M�=���='L���X=�D; >��N>��S>Q�=_�3�S�ؽ@,?��S�����[�=/�r��ID��R�>�QJ>P%���^?2�<���{�V����[����T�b�?|k�?�*�?�����eh���<?w�?b�?=��>�׮���޾�^�Ow��pw��!��c>���>eUp���侈d���\��O���ƽ��D���(?r�>q�?Y�?M��>��>�q,��m��S��.R���^��/��4�[N�N� �����X���j�Y�ھ�P��QP�>�\j��9�>��?�>�`>r�?%�Q�d�>��H>Ql1>֎>^*>�c�=��<S3��F���"U?I�ž�;%����w�¾`OB?$g?=�>�1V�)Ƃ�����^?���?)�?�?�>vWe�F4/��?eQ?�6����?�V�=�������9�<���d�ٮ��ժ�y�x>����1��#P��'����?�#?T��;��������p=�P�?�(?�)�L�Q�V�o�$�W���R�x���/h��=����$�ϐp�o珿Aa���%���(�s�)=r{*?�?w�0y����5k�/!?�lf>���>�<�>��>֢I>q�	���1�^��='�����E�>E{?'�>�jI?�)<?��P? �L?v�>]�>�G�����>��;�B�>dl�>
�9?м-?m0?"?�5+?>�b>d������#qؾ�?e�?�8?��?�h?�.���~ý�ߨ�XIj�2y�WV���C�=1�<M3ؽ2�u��?Y=�S>��?��6�c<�"��7�p>�0?��>t2�>�%��$@�����=&�>�L?�>�Q��m���ܾJ?f?0�ȼ�%=��>��=Z�����<2�<T[{���p=��a�YS���� =�2�=�Ln=Z���v�<�;�\?���<Nr�>�?Mz�>O��>�������`�
���=��G>y�T>��+>�Ӿ����[嗿;�g�)�~>���?跴?(�A=ٻ�=a�=d���Ϲ�>�P���n`Q=�,	?��"?�rQ?]�?Q�:?^�!?Q@>��G����݁��_���?�,?���>h��#�ʾ�N�3���?�^?R!a� ��\0)��\¾2�Խj�>�X/��5~����g'D��$������☽ɘ�?���?�B@�W�6�{�辒���$���G�C?NB�>�r�>��>�)�&�g�4�� ;>�u�>��Q?G��>dT?���?�+`?�aS>�4:�	h���c��`V�;�M)>T�C?☆?�Ջ?��r?9�>ز�=F[@�����u�@��z
��ڀ�%�$=�	r>Ĥ>Z�>#W�>�"�=P�ʽ����9�/���=�p>�-�>횪>B��>넂>��<2�C?<b�>�9ľS�����5�������b?�ׇ?8�,?N�=u�,�C�?���g��>�k�?OȨ?E*?�gT���=�_��k{��6���8��>���>«>��=!�A=+>q�>!��>X-�%��2�5�z�����?�LE?U"�=m3ǿ��n��;v�3���Y �<}�����k����@�b����=�鑾/���w��)�X�+A��@|��$ۯ��������h?�=Rr�=��=F�<7���]&�<��:=y��<�`Z=ƳK�'(�<�.d��崺a{��{_������/=�.@�l�վ�
g?��{?�c?�;o?�z�>��<���>۶?�����B!?V��>�>a/�����'������2�q�_��Ǿ�El<5r�=�:7>�> i>��w=��!>�#-��Һ;��,�dh�= Д��x�='#@=TCt=�r^>!�>�j?Va�W蕿��C��8Ͻ"� ?.��>��C�,�˾�,?/2>.gt��
���@�/d{?�0�?#�?H�?/������>�>�����6�&>�[��'T8>�ݒ=9��%�>o��>��ʃ���/��"�?T�@.2%?"���ƿ�>IhZ>��L��]P�~L �Sg8�wy\�'=��F��>�iD�8��h�>��>�'���z޾�����}>�>���=�(L�XU�=����=���nϷ<ߍJ>�B>B�=ѩ<��-�=�5�a�>�G>C��9�1;jӽl5��;�=ߖ�>�_�=�_�>�3(?��/?9<m?�2�>G������ƕ�32�>,Ľє�>D�ǻR%;�1�>�o6?�:?�>?i�>��>�
�>��>L_,���~��ߙ���ʾ|)p=�r�?�Ku?��>�>�ܽ��.�Y�@��n��l+?��2?�?��>�G�+��zi&��.�nV���䣹.�,=<�r��W�l���~� ��73�=��>���>f8�>w�y>�9>8O>4�>ä>��<^��=�Q��W�<�����=�������<O�ļA5���0�j�*�"M����;�`;�X<���;�H�=��>h�>�7�>U�=	��2a,>�����J�/��=`�����A�H�c��)|�K�,��&;�+�;>��S>�x�U���2?�Y>qH>z��?-"t?��>�h�!оʾ��J-]��eW��$�=��>��=��;��;`��N�w�վ/��>��>��>��l>v�+��?�;rw=����N5����>���%���:��*q�4��:����i��p�c�D?�F�����=r~?��I?ߏ?w�>|���ؾ�>0>�*��Q�=��)q�������?��&?rm�>?*�<�D���۾���(�>��a��Y�5��Î!�&��;WGξt�>Hɟ��Ծ��"�(K���E��>v>�R�~�[G�>GnU?㉲?�+d�n ���E�?�g�ὶ�?�i?�v�>qA?L�?�����߾����dO�<��Y?"&�?�f�?ƣ>�X�=񟽽J`�>��?@�?�?�lq?��9�P��>7�<��(>m\��`s�=�>s��=���=��?"�
?
&?�k��7l	����t���Z��B�<D�={Z�>?��>�ce>}��=��[=��=l�c>���>_��>��a>�Ц>��>�d��zѾ'?&�>1E�>--]?S�0>�^�=�|�=��%��˂��Ic�Ah	��t<��c=��ƽ���aL�{D���,�>�;ٿ�y�?{2>�"�eg?��4��/�2��>I>ͻ��1��	?�W>��>��`>��>�@u>��>2�X>��
��C=���	�&���L��sY��?��DE_>�8ξ�7�P�߻�G:��@��\�Y�T�`&y���c�=i=�?b�I��5��S�ć���d�>�?��E?�Iɾg��<y&>��>���>�����������5����?I�?�Jz>E��>�[?~&?�匾i��<�s���i�������5s�o����nt�����
���G?»O?�U+?U�g>��D>%׏?#�4��� �w.�>3�[�g 2�ڑ�=�u�>b얾�,J;��޾@�����V>,�x?�n�?j<?ho��{���0>�n>?o�3?�z?a3?�W4?� ҽ��0?S ><k?y~?��6?�,?�?%`>_��=7�;���;du������[��6�������r�==��z=�.<k:c<��\<,�7<;ͻ4lI�:�C��o߼��=0h=�+�=���=�!�>w�w?�Z?�_>��*?\��� �D��~�C <?axi������,��B��̾H��=eH?��?�|R?a@>�N�R�J���J>�s�=�b�=�@R>̻�>(����Ċ�-�=��=�q�>[hu=T6��v!ž^��jG�f �D|~=���>B��>X3\����=����V���9�>�1ܽ�Zƾ��i�Q���>
+�+�d<]�>��e?E��>�������d�=>����z?�3$?�IF?��?�ՠ=��y;��i3�򐻾�?\��=�^�瀰�N���9n*���n��Z�=��ʾ'����c>	���޾*3n�'�I���澙P=����Q=P��#^־�A�P�=��	>����H!�=4��������I?��k=&����U�#!���>�/�>�߮>Ѓ7���{�I�@���먖=��>>t;>}k��Ti�KuG��w��_�>�{E?6�_?��?�%����r�A�C�p;�����������?�Ȭ>]C?�Z@>�.�=���������d��G�D)�>���>���H�G� ��������$�?��>8�?��>]^?UfR?�
?Y`?-�)?��?���>࠶�����
A&?h��?�˅=��ӽ��S���8�X F�r �>{�)?P�A�<t�>i�?N�?��&?�pQ?�?Z>� ��U@����>BC�>��W��g����^>�hJ?=r�>�"Y?�?��=>'�5�a7��u������='�>B�2?0>#?k�? ��>���>&z�����=�Z�>yWW?=y??�b? g>?a!+>�[�>��V=���>��>��?b�Q?��q?�L?���>�(;����ýHH��"� �{�<�3=��3=�@��9����c����<�v�< w������_�u?��/!��i8@��>�r>������.>��þ�J��C�C>����
�����:�=�0ѵ=匁>��?�B�>��$����=ʺ>���>���'?��?��?�;{'b���ھ�H���>�eA?5��=)�l�+q��nu��e=�Qn?LJ^?��Z��5���b?2�]?ɜ�=��þ��b��"���O?Y�
?=H��ѳ>7�~?��q?X��>�f�H0n�����Mb��j�G��=Q`�>�Z���d�p?�>ʍ7?�%�>�c>�z�=�f۾��w�������?`�?Q�?���?�A*>��n��/࿘��Y��1d?}��>�z���+/?ů��oƷ�ach��><����ۀ��୾�ي�ᆟ�^���$W;�N���&=b�?���?Tem?Eq?6}���Zk���N������H�_	��1��5I�ME�2�P���������]ͷ�Ż�=��f��r_��t�?�*?�M�Z�?�j��Hƽ��)��艈>�e���;V�oJ=%����=|��=�����53ž��?�
�>�C�>k?? ^�W�9�1�.�5�:�̯;�9>߯�>��z>�2�>��*�F���"��4�۾u𔾲ٕ�F�m>Y-k?Ly?�=�?N�=mB��џ�#��N��=��w�>���>Qj�>jC�to���"���5�I�W��y��S����	���=	?E<>�K�>�Ԡ?��>'���/9��R捾�������=�?6oB?���>~t�>Ǔܽ���@M�>88n?&O�>���>�>��ݔ#����+�Ƚ�[�>�I�>�K?� �>U�)�ױ\����L���
�9�Ǳ�=��d?+���v�b���>��M?Є
;Mɳ<���><t`��!�X�G�$��+>R�?1��=I�?>��ž
,
��x�����;�?���>r5��vY�Jk>_&?��>���>�ӓ?G��>\��� ����>�N?#�R?��B?��>�:A>�[H�� ��?8����=`�g>�`>N�K>��t=�IX��֥��&]�-r�=X��>RT>t��-̻Uؘ�^���r�z>!����ҁ�E
�s�M?˾�<��>i��N'�C�ƾRI�)_澺���  \�@ ���ڽ�xP�ȈM�P��c�x�-?@!��?"�̾3i,=�Q���%����о.T?	�� 9�3���'������!�xF�ۄO�L�]��ad�/���'?8�����ǿ,����:ܾ~ ?A ?��y?B���"�8�� >t[�<�'��מ�;���^�ο�����^?%��>�
�B��2��>Ǡ�>[�X>�?q>���3鞾�,�<��?χ-?���>�r�q�ɿ1�����<[��?��@�uA?��(������V=���>��	?��?>>1�:��ڰ�KB�>�;�?\��?ȞN=��W��
�ue?h�<��F���ܻ���=_��=x1=���|J>Y>�>fw��LA��3ܽ[{4>ʅ>�v"�\��[^�x=�<ӕ]>:�ս�=��8h�?@w_��U������=���<�>x�=?<ۇ=#�@=`�?AR �᾿�����:?Ţ�?���?f�B?������>a)��^;?�)?::�>�3�_a��3:P>����>Ǟݾ�J�=���!�>V*�=�ǡ���Ⱦ��M�k_��->n���YԿb)���-��R+=n�<�B��m.�9��N�����5	G��v����=N��=��Z>�v>F,>.�7>,�d?�d?�ו>��c>hʙ�����2��|�,<H���2��G@����z�*и����� ��1������
�%5Ǿ�=��=�8R�V���L� ���b�R�F���.?Kj$>��ʾ*�M���,<mʾ����w���饽@3̾��1�fn��˟?��A?Q�����V�]���f�����d�W?�J����PI��=?���*�=�!�>���=���� 3�~S��0?hH&?�ᚾ�Đ��1>K�����*=�C8?��?.v=2D�>�z
?ձB��ݽ'Ҙ>��z>h�>��>?]^=��~� �˓?��N?������2>�Tž�UU����<��=]E��x;�w>W����C��-rb�:��ox��eS?~ �>��+�����r�����?�=��r?P��>�J�> xh?w<?�J=���SpU��x��"<=��[?��l?f>j�[�T6Ͼd���5?E�_?��@>}f�g���B4�`��G?�1j?�?�押��y�Ǥ��.�KX;?~�v?b^�cZ�����8�W�vd�>.7�>`�>��9�v&�>�>?�"��A��Yѿ��4��Ş?��@�k�?��6<Ʉ�G�=�?q|�>�^O�7mžW���赾-�l=���>�x��Wv�� ���,��9?��?���>�낾�W��� >�<v�a>�?��?"Hþ@$$=�@3��s�9ͽ����=��<��=��B�̛�Մ2����V6��|��d*��>:h>��@���C(?P��Z濇*���5��u+���ޕ�y%?;�}>K�i���U�c�����B�m��Z>�9�1��;�>��>�ۖ�ؒ��|�^�9����%U�>����>�I�����eР�-�:^m�>v�>�K�>�z��߽��ԙ?������ο�������|sY?�?�*�?&M?�D�<�,v�_�}��􉼋cE?D"v?�[?��e�`��_&��)j?Se��xt`���4��!E�|^U>B^3?�`�>N�-��1z=��>#h�>��>�.�2hĿv��������?6��?-���>d��?��+?�{���������P*��+�9 S??�/>�¾�]!��=�%	��4x
?�/?'�����]�_?*�a�K�p���-���ƽ�ۡ> �0�f\��M�����Xe����@y����?N^�?i�?˵�� #�e6%?�>d����8ǾC�<���>�(�>*N>tH_���u>����:�i	>���?�~�?Nj?���������U>�}?)��>���?	�=��>��=)��Ol�P !>]�=m:�Ɯ?iN?:Q�>\��=�9���.�ZAF��R����CC�7��>�a?��K?��b>R^��v)�Kc ��mν~I0��J� @���"���׽�5>P�=>m�>s�C�N�Ҿq�?�t���ؿAm��x(���3?N�>c�?����s�����^?���>_��6���1����>��?,'�?	?�׾�μ�/>ʭ>p��>��ӽ�.�����4`8>!B?l�����
�o�b�>���?x�@Uɮ?��h�}� ?B�?b���s�z�#�H��ޛ
>��>*���|=�]3?F&>�i�9��k:T�"��>�7�?�]�?P��>MD�?|j��vo�aAG<�ف>7�?9{�>��a�o�4��	�>��*?r+�kE��zG)��^�?�@K�@��4?m;��egֿ'���7L������J��=Q��=!�2>��ٽ�m�=,�7=n9��?�����=��>�d>�q>�(O>�a;>�)>����!�Tq��ۢ����C���M���Z�2���Tv��y��3��(���,3��1ý~���Q�23&��*`�^>D�I?lof?�7�?-s.?�K�=�]�=�H��<��=�#B����=��>�BC?r�[?-K	?�~� �~�%V�{~x�ԛ�vϔ�6�(>�G'>��	?G�>���> L�=�
h>E3.>�m;> &>S�>��=<7��p��>��>5v�>�
�>}C<>��>ϴ�1���h�	w��̽� �?���0�J��0��!>��%���x�=P`.?�z>���w?п���%0H?����&�ɻ+��>��0?�`W?m�>�
����T��)>���e�j��b>�& ��yl�ы)��!Q>�h?"�6>Cv�>�6?��:�������#�>xW?h���"�L���O�86���,�>L��>�_��3N/�Oã��f�u�о����`?�b�>��+�b(Ѿ~��G�)�%��> 푽-�+���>&�W>��#�?`½�uh��&�=dQ�>ޗ>[	?a�d>䓰=�m�>/�����j�oT�>��>�#{>OD??�M?|q��]躽�����潵>�>Gz�>J/�>8Y�=
�Z�J�=���>`N>��3���������<�w>�B�����嚽F �=$�g�)��=�-�=M��DI,�p3�=�~?���(䈿��e���lD?U+?W �=F�F<��"�C ���H��F�?q�@m�?��	��V�C�?�@�?��V��=
}�>׫>�ξ�L��?��Ž3Ǣ�Δ	�4)#�jS�?��?��/�Xʋ�;l�n6>�^%?�Ӿ���>M�TG���X��=��w'��)h�>� ?}���Ǘ=�FZ���>p)�>�Ϳ�����Emɿ�QY���?���?��?ׁg�<f��?�H��b�>x��?VW?et,>�׾�j��ұ�>��+?A^Z?�N�>��ͽ�`h?�:�?�tT?9vt>�ۖ?�\�?]�$?�'�=۸E��ѿ��~��6>: �=F!�>���>1�ܾ�z�����U�m��eb�����s =l��s|�>�c���ݾ�ԅ>��3�6 ��I$>���>0[=�ւ>ro�>p�+?���>���>�cĽn�+��z9���D�W�K?���?���1n�J��<���=d�^��(?jC4?�4]���Ͼ�Ĩ>j�\?p?' [?�a�>��� @���忿
������<#�K>L+�>�C�>����>K>o�Ծ�D��_�>X��>Q���=7ھ�'��h���G@�>Ne!?���>���=Ǚ ?Ü#?'�j>)�>aE��9����E�7��>���>�H?�~?��?�Թ��Z3�����桿��[��:N>��x?�U?�ʕ>?���σ��w]E�lDI����K��?\tg?WT�+?,2�?�??-�A?�)f>1��Dؾ������>�?�4Ӻ�	a�jh�8w��
b�>��"?�=�>�q��ҋ��2o=�'��žf�?|�?�:�>kA7�A���y0Z��%H��O�=�B�<��m��O�s�<>��<�P�18>W�w=l���������}�rR�=W�F>q��>��!>V%������-?9+����p����=J����"��H�>@:߽Jn��-U?�JW�����,���a����d�"��?Z`�?��r?�=<ᆿ2�T?1��?�k>?�_G�-|ξ�Ѿ?E=��#˽LhȾG7>��>rm�(��%��.��ʅ��%������>��>$�	?O- ?T�K>N�>}
��J�'��J��`���u^�����_6��.����p�����-���ż���B�v��o�>�N�����>� 	?�f>��y>6��>5���O��>�P>�Bx>Ĩ>[!X>�B7>z� >`�<�� �/?厸�Q�?�����t����#?a�r?8��>jh��x�aX�&��>�y�?Y��?,�p=6�z���I��^�>3O?i ���f�>Z���3 �=�E�= ���(�0�`R=��=��=�j�����8��Ę�v��>��?YV��Q�)�5z�����2�s=�C�?
�)?�)���Q���o���W�k�R�]��WKg�A>���%�G�p�я�q6������L�(�^�)=�)*?t5�?y�#��o���uek�{�?��8e>���>��>ְ�>5�H>��	���1���]�R\'�
h��q(�>��z?�s�>�,.?�1;?Q�4?F�F?J[�>0 c>��E��� ?�,=Jw>�~�>�q(?̆+?p�5?��?�x?B�>�+n�K8��	�龽��>�?��?���>�g�>Y���M^�O���[=�qܼ���=�&>�]~���D����<��;>�F�>^���u�E5�+)���D�>7�>?˝y>�`9�S
[�T/:u�$�r�2?b��>:�G�່�F+��f?U�?X�jܐ=0��<_ �=Z[>#+a=dC�=C�=�=�,��� �^��=x�<���=�;> .>�\$�w�����S=�u�>��?���>�C�>A@��;� ����7n�=Y>�S>�>Fپ�}���$��*�g�O_y>�w�?�z�?�f=��=��=�{���T�����M���*�<�?0K#?�WT?Ǖ�?��=?j#?��>�*��L��r^������?L�?=��>�7���ʾ�9��U;��,?�?��D�l�ݾ��K�|����e��=&�X�j�����?��?� ���_�77�?(��?�T���.��|��٠�g���K�1?�}�>���>~��>��1�<�n�d���q>�(?��S?$߶>ʷO?�(�?d�k?Sˁ>��%��)���;��I�*<W >�~9?[�?��?ѱu?��>!��=n"*��.޾�V �buO�h]�Ot��S�e=���>�˥>D��>;̣>�k=^q�����)� �y��=�Ȏ>�7�>���>�4�>�w]>$7r�PVN?,l'?mX�Tr���c��Â�����=.�?�@�?#	3?�
;6��[28�֓��6�?<��?&�?˚A?���:���=��W��[��V�k>py>#�>;A=�5D>/k>�>,w>������
���@=��>��#?�m>��Ŀ�_q���v�5ɚ�.��;���{�\�΢���b�ޮ=�����v������W�@I��/��?a���_����u�[^�>�{=~��=?a�=���<�c���D�<��E=I,|<Mu=?q���l<'�#�;����·�ݗ�vO<�U=Ɉ�G3���wt?��`?�O?n[7?�AJ>L�"�b��Z�>�@�<7?��>��'=*~��38?�q,���J��h�پ�Ӿ�u�G0��`�'>�wH=d�7>��A>��w>0���_=��=oG�<��.�X�>�S>�ޕ=X}�=�9>�(>(�>��y?.Ow�U���I�1��^��-,W?��z>ҁ�2��".4?/b�>9�S���ſ��=���?)o�?�k�?Yz�>���+�>V����l/��[k>��A��>$��=�.����>H\�>�E�zt��gd׾-�?P�@7�]?�{�g2���>�&6>�@>�'T�Ms1��4X�M�e���I�>'!??�;�m;���>U~�=��۾ǌ��R�=�</>�� =9$�QX�g�=��d�q>=�T=��>R�D>r��=�[�����=�K=�	�=�/J>���@�d���@=΄�=H�[>�>A ?�? �&?�:?��?Y����A侸��P�>;c�>H�=V�7>�E�>�t�>9�)?*�(?�X]?�>������>o��>d0w��:����9���w��=��?s�X?�>-H�=
�8�j�qtI���>��,?/2?�x?�P0>�X�h]꿗�(�5=��$��k�;�=��$���kp��i"�\�o�YA
>���>g�>t�>3hS>ž	>dX/>G�>��	>۬���=5=�:�<u��;Zy=j�
��E�=l������]�m���ޫ����<�Gf=��'<+hӼ�u�=; ?!Q6>Ggl>:d�����O)>۽��^�+��+>QZ���?�V��3ߒ�����+D��g>�qP=�ƹ�u��f#?J-�>��<�X�?�g}?�*=����>��	ʖ��n��>�;z,�=՗:>�l���X��Xc��m6��C����>E��>���>��g>��*��E>�Q��=�����5����>�����9��{�o�}򤿠����i��뺺��F?�̇�b�=��{?5=I?D��?h`�>��
�վ3=1>�������<NC��p�����ie?%�'?�g�>Bd�_D��^��r�_H>1���HK����Y����߼����*�=���7?��
���j��9���%V�p����=�>V[^?3J�?٨��y�:�n�k��WV�0~U>!�?(g�>|���JK?D S?�X1�����ť���ɾ;�9?27�?\��?���N	�=m��\Y�>n?�ϙ?�ב?��l?c�1����>M��<>�>Y�(�D�>z�$>���=��=��
?�H?B�?�����և������9p�=�<�7l=�+�>#w�>�Y�>mr�=K,0= ��=�:X>�4�>���>�o>��>� }>�m���6	��S-?�4=igu>��X?��=�޼��5�ճ�=���<SE���ʾ^��>�U#>ҫ&>2����WK���>L���?��>_��jK�>�zA��^�>��>T�>�F���"1?P* ?[�?��X>���=�ٷ>?��>I�3=��,���=�H&�u8��i��`���2H�>���Nm�����<�{�{?ٽ1���� 3���l����j)H�8�h>�<�?+L}���.�3��ޯ��L�>"��>�!?�'�����W#>���>��>qn�`���^ҏ������?*&�?�;c>��>@�W?�?��1�3� vZ��u�V(A�e�U�`�}፿����
���'�_?�x?,yA?�P�<2:z>N��? �%�lӏ��)�>�/�';��@<=s+�>(*����`���Ӿ��þ:8�(IF>��o?7%�?yY?<TV��T=�=>��D?n�E?wҍ?f~C?
?��E���=?�K^>QȺ>i�'?G>N?˵L?~0�>��>>��>3P�<ps��a��w���W�^�����=JI6�T�=3��=���>J�ż80 ��_�<��n=��	�6����<�� >�0�=�Ų>�\?Rj�>�j>@-+?��#�>�&�a�n�j�A?�w�=�z��p���՚�ZL�i�E> �m?�̨?��]?�'>�\��V�>F+q>a�">��h>臛>�3�	{Y���5=���=�7>�B�=nܼpz�������jn9&�>���>�#>�����#>�Σ���x���e>��M����%�Q�1�F��1���y���>�5L?��?�=5��}�f��'?�4<?:L?f�?@��=�?߾��9�_�I��=�ؠ>��<� ��衿ܜ���];�|�/�e�q>-�� ����-b> �� n޾�n�{�I����/�L=�{��}W=t�#�վ�B��>�=m
>������ ��
���Ҫ��,J?!j=@c���U��p����>��>���>��:�_(v��y@��׬���=O��>��:>�z����mG�,4� �t>�pK?�Bd?��?j�\��t��.E��M��������Fl?�G�>�?�D>�=�R������k��&J���>g��>����l9���������-��К�>,�?m�=d	?s�M?L�?�a?�!?� ?߼�>�/?�:��^B&?І�?/��=��ԽV�T���8��F�� �>{)?��B����>��?�?��&?Z�Q?,�?��>�� ��@@����>AX�>��W��_��
`>��J?��>�5Y?�у?M>>�5�(⢾���=2�=<9>c�2?�5#?:�?�>���>u���C{=�{�>��a?��?�6o?˓�=)�?�J->fF�>]8�=G�>z��>L�?a�O?�s?�hJ?��>~�<Ƣ���Я��>}��Q9����;��&<[<T=�H�9�?��y"���<rJW��ͼ��C�b��h�K�N���^G<��>?j>f{����>�ʾ���,J>�PV�ˡ�&m��r2�4�=�p�>9��>v�>�h:�ⅅ=Ɗ�>p}�>�3���%?�C�>�D
?���<�X�8!��{���Ř>ـ0?>o�\��}��C�q�|ũ=� v?;�h?,�^�4m�s�b?��]?)_�`=���þ�b��c�!�O?A�
?��G��۳>��~?D�q?g��>!f��;n�����"b��j����=�x�>_O���d��U�>�7?2u�>�@c>�M�=�۾�w��<��Y�?b�?���?� �?��*>$�n��2�#l���뇿��j?&>�>O�þf�.?Y���kǽ���:�.���#��{��Ć������&���p��솾��	�"��<��?W�?,>n?->z?����N�v���J�N*��~F�c��/��!J�	<I���D�Xpt�p�,"��Ҿ��=�肾��=�S�?Ft?S�m�!
?�,���پ����F>hKԾu̽A��<���
��=�2�=�x_���6�l����*?�v�>{s�>�F?�Y���A�{;&��g:�H��/>dA�>Z�j>���>�G����I�`��4�ؾ�w���u���bc>�ul?3�R?��u?�4+�C{��G�#�reS<vv���?>@�/>g�p>*�o��{%��$��g?�&�z��2#��X�	��4�=D�-?V��>Z�>�Ò?n+?�� �6����Lw��('��=�Ƹ>�Ye?�M�>|>Ԟ�������>Y�l?���>�a�>a���D!��|���˽�k�>8w�>B��>�Sp>?�,�g'\�Na��0z���9���=��h?���za���>,�Q?^��:�tN<�Z�>��u�c�!�%�^�'��">s�?���=�;>�lžk���{�O@��B�)?{�?3)��	�*�n/~>��"?�	�>���>Ϡ�?|ҝ>C�����Q���?�_?\	K?N�A?�1�>��=#��RŽ��'��M-=�+�>�Z>��q=���=.L�I�[����<5I=�J�=�u�d䮽{0<���D�X<�3�<�H0>�eۿ?K�j�پ���C
������񱽣z��֋�F��E����.x������'��6V��c������l�4��?�0�?*m���8����������B���\��>Mq�!�~� �����핾n��R����i!�2
P�*i��e��Y'?�����ǿ����2oܾ��?�G ?�y?;��("��e8��6 >a��<����z�����7�οf���0_?��>� �9]����>En�>��X>z�n>�܈���3�<Rn?A-?���>�q�]ɿ�w�����<��?��@f�@?�Z!����Y:�<f��>!C?*BQ>r����S,��y�>�×?��?��J=��T��e���^?V��<�1A��'�;80�=���=s�<��½r�V>���>�ӽ`_���A�n>u�>ί��d)��x+����=���>��2,�'��?	�A�	b(�ՅҾG�Z���e>��6?l���J��==kN?	f���ڿ�񁿍��?���?���?;+?��Ⱦ��=՗ž
�L?8Z"?���>�()��/��cʚ>y�>>��>�뾝'���t�>I+�>�I�h�s�s琾C ���2k��[�>����ƿ�|%����-�=-G��ՒK��L�5���`5T�������k�����T=C��=��R>f��>��Z>'_X>��V?=Jk?���>2v>��eA����̾��5��L���F��@���أ���쾖�޾����+�����Ⱦ�=���=�"R������� ���b��DF���.?��#>1�ʾ��M�x+<� ʾ�ª��Ԉ�������˾�]1�5�m����?U�A?߅���V����F�丽ݪW?�����Zm��"�=$j����=��>���=up⾲�2�
mS�]1?=A?���^����*>b#ٽk4=Q�(?���>WyK<���>��"?�� �{���c>F�G>�%�>h;�>�_
>����Z!׽G�?�N?� ��:���FՋ>Oeʾ?�l���=�=��.�R.r��9V>���=mu��(Ƽ�v���>=��,?�|>a�%�I`)�)����i��2@>�Ht?L��>g��>
]M?�"$?��L>�ʾI*M�:� ��r��ee?��m?T>��ب�'Bf���
?��S?����辧SU��T�' ��;�>U�{?��?w�3�?�{��^���Y��(a?1/K?L�h�闟�}h������->*<?�>��=�kd�>2�0?.W��ݵ������<�/�?��@ŵ�?Y��}:�~>H�?r�>����Nþ Y��������;�?�T��E {��S#�˥D���(?�*q?L��>��X� S���E=g��ɰ?��?�ݾ����n�)�:%f����"�z���Ľ"�~�f�0�p���(��x��~���>Ӿ�ɽ�^�>��@����S$?B4I�� 뿸����Ĉ��žĶ��v.?�>cS�7�¾��{��-n�[V=�!^��(>��t�>�/>
 ��������{���:��Ӑ��>�\��c�>1�R�o뵾v����4<��>�T�>|�>{���RG�����?�o��G�Ϳ1s��d��ZX?9�?zH�?4�?�"<(�s�g�y�͉(��zF?Pss?S[Z?����]�Z�>�B�j?�]���Q`�4�4��IE��U> 3?�;�>^�-��|=|>|�>�>�/��Ŀ�ض�(������?���?�e�4��>x}�?Aj+?�b�5���H��\�*��E�|2A?].2>G����!��-=�˒��
?��0?({�34��_?�a�c�p�.�-���ƽޡ>�0��k\�Pa�����Ve�~���Cy�$��?M^�?H�?��� #��4%?#�>U����8Ǿn#�<��>W'�>k*N>�P_�e�u>����:�pd	>m��?n~�?j?{���<����T>�}?��>��?���=��>|6�=����N4���#>�A�=p>���?^�M?�H�>�n�=H�8��/��UF�YaR�j4�ĠC���>%�a?b�L?�b>�˹��z0��� ��ZͽJ�1�F-鼘5@��H+�c�޽�4>��=>=->�HD�"Ӿ{t?k�&�� ׿��͞�A;?�Y�>��?ȋ�+$�����=�Y?��>���}��Pw��x����G�?I~�?�� ?:�Ѿ��`�ƥ�=r�>�h{>��X���p������>��9?�穽 ����d�a|>Q�?!�@�?�_��?pW�hS���H~����7�j�=��7?���x>n�>v;�=��u�ꍪ�O�s��{�>4�?pI�?��>Cwl?�o��qB���-=<]�>Q/k?�2?^֍�i��$C>we?��Fێ�lh�@�e?�
@�M@ `^?����������{��}Ҿ\�r�=a��B$I>�b�=��;~�m�W>�C�=�ř>%�>ǽ�=L��=M>/P>��(>��{������ֿ2����@L��5����[���xi�ԹP�kB���k�]+Ǿo�0��K��,5y����<]��=�-F=��j=x�a?�^?�X�?��?X����=��ܾ��>7vٽ���=��>;2.?;A?�"?��p=���5Ku�����y��s�l�>h�>�Q�>#�>��>��v=:PA>�J�=���>�O�=���= �=K�;�4D>Z~�>� ?g��>�C<>��>Eϴ��1��j�h��
w�U̽1�?����P�J��1���9��Ц���h�=Eb.?	|>���?пd����2H?%���x)���+���>|�0?�cW?�>��T�T�1:>;����j�5`>�+ ��l���)��%Q>xl?��f>�u>�3�@e8���P��w��'j|>�46?�趾r;9�K�u���H��`ݾ�GM>�¾>D�Ai�.������li���{=�x:?��?�N���ా�u��E���VR>x?\>5>=XY�=�`M>�^c���ƽH��.=��=��^>��?��&>�J=��l>b|������#�>&�G>���=n/5?�Q%? ���,�	h���1����>H��>�L�>�L>��gn�=���>"�1>�>8�r��>��^A��B~p>qa�=#�m��.[�6�m�(&���^�>}�>]�4���E��~�=�~?���&䈿��4e���lD?Q+?P �=ɝF<��"�D ���H��F�?p�@m�?��	��V�A�?�@�?	��Y��=
}�>�֫>�ξ�L��?��Ž<Ǣ�ɔ	�)#�gS�?��?��/�Wʋ�6l��6>�^%?�Ӿ���>´��혿������u���=���>n�H?���@;��];��	?��?��n?����ȿ��u�@��>�_�?/��?�l��E��S?�ڢ�>���?�iV?�[a>��׾4X���>�z>?��R?rͶ>�4���*��?�k�? �?i>>0s�?��?܀2?����V7�A]��/�����>#�ݽ�->��m>M-�DfP��%���f��(`��H�k�=��v=Oѳ>"��(��'0�>F:�=�оYsu����>?4�=[�>��>��?>�>��>=墽҂ѽE���p-p���K?���?$���2n��N�<Ġ�=��^��&?tI4?�k[�S�Ͼ�ը>ۺ\?e?�[?d�>.��D>��?迿!~��ɩ�<z�K>4�>�H�>o$���FK>��Ծ�4D�Sp�>З>�����?ھ�,���J��bB�>�e!?���>Ү=̙ ?��#?Tnj>���>"eE�P-��*�E�X��>��>>;?�~?��?0���sE3���桿׋[��gN>��x?�Q?Xӕ>�������5�A��GI�`��R��?8Jg?�潯?n/�?�j??͎A?�9f>��2�׾6̭����>"�I?ݎ1�mZ
��%����N?e�>�b=5"R���G>��m>-�;�#�
*<?��?B?�堾}�6��	����=[	������:>V�=��X>	g�<m6�����<mY>�>S�txԾ}��>�G>�dE>�[>��l�勛�W>,?��F�(Ѓ���=_�r��zD���>�,L>`���|�^?��=���{�A���s��8�T���?o��?�`�?�̴�z�h�r,=?V�?��?�"�>;A��{޾�t��w��Xx��|��>���>�p�R!�Ύ�������J��z�Ž�SV��?Iy�>�1?� ?|�s>���>3,���T����� �5`���#���A��!!��	��˦�i�j���}��[ܾ�r���>\�T3�>��?L�>:y�>>m�>�R�B��>��Y>K��>�W�>
 >���=G�=�>��Q��3P?���RQ#��B�r�����:?�^?�g�>d����΀�˕�3?���?�=�?�L>��j��(���?&!�>��c���	?3=b},�B�A=.z��_���t�һC����tT>|yռt�(�11M��rm���	?�M?=Q�ʾ��1��⟾D�=ދ�?�0?$�.�)T���r��X�D�J���?���r�����_Y)�#p�ӄ��΃���"����,�Q!=	�)?���?���u���P�k��>��-[>���>�n�>���>�U>c���0�C�_���'�@߁����>��x?��>>�I?=<?GuP?�jL?0��>�c�>�4���i�>���;��>P�>��9?�-?-90?�{?yt+?u3c>��O ���ؾ�
?��?RJ?l?I�?�ᅾ�qý�7����f�A�y�O��� �=Kz�<`�׽kGu���T=9T>.k�>q[��d�"��S���z��?�]d>
��=;�N�����yѝ�k�Q=��K?+��>��󰐿9im�\?uפ?��=�f�=�>�d=������=�a�=�uJ��΀<�߃�7�㼐���ñ=�Vl=�-�<�8=�r�=KTj�*U��k�>��?Z��>
:�>�;��Ϋ ����데=��X>� S>=>?پA{��'#��&�g�kVy>�w�?�y�?)�f=;#�=G��=�w���R���������<��<�?	I#?�VT?��?Z�=?�l#?	�>�'�dM���_��u��S�?�,?肑>���s�ʾ�𨿺�3���?C^?�;a�b���6)�f�¾��Խ�>�[/�p/~���D�T	�����#�����?$��?dEA���6�t�������L��p�C?K�>K�>T#�>��)���g�'��;>ӏ�>�R?6�>�ZP?�{?n\?�uV>|�8��"���X�� ���{�">�D@?/Ɓ?ο�?��x?D�>�,>��*�Ĝ���q��4��n��:�`=�%[>�6�>��>���>Ռ�=�cͽ�ί��@>��k�=�=d>��>�G�>���>K�y>��<��G?3��>y4��(��G��.؂��}9��Pu?�7�?"+?��=�;�CtE��{��.T�>�\�?�ث?�*?�PS����=��ռ.��v%r����>?�>Ę>6-�=�=H=�,><��>�j�>UH��C��17�QLA�e�?D�E?�q�=a����Az���ɾZu���">4�ɾ� w��=������4�\�����o�6z���jϾ?���Jo�w��-=T�d�>�yB=ׯ�=<4�<�r>�n;�=���;�u&=HD=Z�Ƚ��J=;����?�uYS��t�=�ǰ=���=�n�y����:�?�Og?�IL?�%Z?��#>��|2H�"�>�W���>���>�=��˾��(�����7	������R��"<��F���ؗ=6����>�g�=�B_>*A>8��;z�y>�F�=��=�	>t.�=`->��=��>SJ>?{�=�z?�d����FW���ýќA?׼�>���:��;��I?�e>h�h��㩿��ݎ�?���?�޽?�m�>~>���>�o���C1<u�=���Qk>��O=H٠����>�!�>����Ք���~�e��?8@# 4?���Ko¿`Ѩ=����*��rb���D���N>[�Ҿ.U�>wJP?�ya�T/߾AP�>���>���U�lH����	>f+?4!\>Y��Ö>!�<��>��= �.>�=�>E�>8p=,�E=h��=�
�=�`>CQ�=��<�P>��=ir��c>�>���>`�?t-0?}�c?m�>�,m���ξ����eҋ>���=Lv�>��=l�B> �>v�7?��D?V�K?O��>w��=�
�>u��>n],�Ǚm���Qy���3�<t]�?#��?P�>'`P<A����[>��9��Z�?�-1?�1?���>T����]&�l�.��B������i+=�Nr�0�U������R��n�Y�=Nf�>���>r�>Tmy>�9>��N> �>G�>)t�<�^�=�A��+��<�(��
��=�c���h�<+�żܣ��ɱ&���+�G~��f5�;`�;|^<%��;���=,E�>\�!>Br�>��=J����@(>�Ǚ�c�>���	>$G��M�C��g��I��'����"u5>�t+>�h��m���W?�IH>$�>���?dy?V�=�ݽ�MҾ�f��'�7�ȆX���=��=�ua�	A��_�-�B�;�8�>��>�t�>w�j>�%,���>� fz=ԗ�|K5��N�>�g��@� �T����p�����響n�h�z���bD?4.�=ڑ}?,�H?͏?u>�>�ѓ���־+�->�u��d=�X�[r��Ք���?>�'?�:�>쾋.E�ۡϾ��ͽ�D�>�K�_/P�>ݕ�q�-�����Y�����>�%���Ͼ�`0�����@) C�mZl���>�N?KL�?Q�j��v��£P�S1������?��f?��>p�?��?!���]	�W쀾Ͱ�=�m?Jp�?Я�??n
>5��=�ٱ�'��>ì?��?�n�?W�r?�O;�C#�>���8F�%>-��<C�=�b><��=[��=��?!}
?�	?G���[�����]��Qh[�ۂ=��=ƌ>�>�~>���=�`i=a�=�EW>n��>�u�>��`>K��>�Z�>�-�	����$%?�x#=q��>�J?:�=�8>���= ��4��	��Ɣ��'���2�<r��=u;bf��U�;�>}�ʿ�?nl�=��A�iZ ?���ZY�<�^=��=�X���\?��>>�>�D�>��>h�A>q?a��=�(Ծ�w>uS��!�p�B���R���ɾ��>����Yh����P,�;�A����)��]�i�������9����<���?b� ��di���)��/���?�7�>3?	懾�p�>�?�>]ޓ>Y���Y0��c���-��:�?aH�?�<c>��>��W?j�?W�1��3�MuZ�x�u�<(A��e���`�0፿�����
������_?��x?�xA?�Q�<�:z>��?e�%�;ӏ��)�>_/��&;��:<=�*�>�(����`�H�Ӿ��þ�8��KF>�o?	%�?�X?�SV�F�m��'>��:?ћ1?�Ot?��1?a�;?�����$?^o3>�F?�q?7N5?��.?$�
?B2>�	�=y
����'=�6���O�ѽc~ʽ���!�3=@_{=͸� <��=���<H���ټ��;�%��6%�<3:=��=�=>�w]?���>�2�>9�7?�C��18�vx����.?��:=s�������Z5�L�>5�j?j�?.dZ?�d>��A���B��<>�s�>;&>�/\>I��>�F���E��އ=��>�n>���=��J�����4�	�����v��<�>4l�>���>�=�<��v>pΠ��ۓ�e�}>�6����Ͻ.��<��f���0��˾��>�W?��<?��T=�����/=�1��ڋF?��?/,?�
�?(T>t	�]���J�&Ut�$7�>,Wp<��ξY��l!��e�U��i�%H�=p��&����s>�K���%־M�n���O�In�֔n=nv���)=FK�T�ݾ����;�=rP>����������%���;FJ?�lN=,(��:�I��0¾n>�G�>���>��E����A������u�=:a�>�u<>hX��a����G�(��5)�>�SC?��e?���?�?��kz�� J��D)�܈�N�=�.?���>�?�>�*�=����0b�we���-����>�A�>�3?�$������G羁>���>�Է>�'==g�?lJ?��>%��?��.?@�>�$1>%��<v���\?�Æ?�6W<-��=�E��=��}V����>b�>�M���g�>�g?j�?�C??3/W?Ő�>|?�:�ס��F�*�y>P�>�{n��h���m?>��\?�s�>zX�?�a�?9ԉ>��5��	������3">��>OG?�� ?(u?���>F��>�ǡ�đ�=���>�c?.�?��o?
Z�=s�?�2>���>t��=���>���>�?8O?D�s?��J?���>g��<���+d���s�8nS�2Ɋ;�I<��z=0B�iWu�h���Z�<l��;�᷼�����&�{�D�v��ق�;�T�>T~?�u����>�����j��-�=��:=/� �c��
D��ݬ<�;?�W?�M�޾A<3�J>�?�Q�C�?ߦ=?�>�t�<g�����	Q���O�>i�'?�*x���Y�i�o�T3���bƻ�'|?/�G?��'�Ys¾f�b?��]?Kb�-�<�T�þa�b���|�O?>�
?�G�Xճ>Q�~?��q?���>��e�':n�,���/b���j�@ʶ=m�>�B�T�d� �>.�7?�L�>K�b>��=1t۾u�w�(v���&?�?��?���?�B*>p�n��(࿁���>���^?q��>\���$�"?X
�W)о�㋾V��g��]���2���z��ah��7n#�U���<?ؽԴ�=�?f�r?uq?�_?  �f�c��^����s,V�W��/�B/F��E�mC���n�G)��f���Ø�"?G=Í���޾�M�?�.�>�ɡ���>n�ھO9�k�ᾧ�>�ob��2��L���c�#X>���>�����4�����c?���>ѻ�>^M?2wI�#cF�z<1�|V�Ur�� ��<��>)�>&?�J�>�����~��?׾�c���T���u>��d?�I?sho?^C�Q�0�
���ƫ��w(�=��t�7>W�>���>�^E��8
��&���=�ѧo�/1������w	�Th�=�.?�1v>���>�#�?�?e��w����U�2����<',�>D�f?3�>�U�> E�m%�}��>��l?��>���>^Q���g!���{�!˽>O�>	�>��>j�o>��,�8/\��l��/~��Q�8��/�=ƌh?W�����`�g�>X�Q?�:m�F<њ�>P2x���!���H�'�7>+w?�[�=�m;>+�ž�.�͘{�B$��-6)?�?����)�q�~>f�!?���>���>��?ٝ�>�wþ����!?�_?�aJ?Z9@?U��>��#=Y����Ƚ�&�6+/=��>!|Y>ƶm=�0�=L�M�[����im?=P.�=Aeȼn���P^<�����T<���<�3>f���[�E�?��T@�l ׾u���
]_�qT���T�ݩӽ�+������Q��$�CȽ��n7���a��K-g�70@q_@_������+��uK��	�Ѿ�v�>�^��n�/ݰ�xց��P��7s���]s,�5l{�f�����}�z�$?�+���Cʿk������0
"?�v?�Zu?2 ��f�X2>�1>"��<���<;�/���<˿_)��\?�B�>����-���@�>(Ԏ>�
[>�A>`�m�p����5�9	�>�;4?��?��:�V�ʿFɿ��Ε;���?�Z@�8?:44�����դ>���>��%?A�$?�dоL89�m���p*?,�?ˑ�?��轿J��%�F=�)?�v�)����]���{὇�>�=�=�RQ��\>�i�>�^������B>�r
?�o�>]qý���<h���>��>����".�5Մ?+{\��f���/��T��U>��T?�*�>U:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=z6����z���&V�|��=[��>`�>,�ߋ���O��I��S��=�����ǿ���R^%���K=�s�<��s��������"�����qYi���ͽ?�j=�m>��E>v:�>su>,Kv>S�b?�q?���>͡#>_ڽ����k��A����i�#	�!|��"���2���o����"��N�#�?�r�ľ_OG�;��=��P�����c!'�|�_��F?��B)?��#>��Ͼ��K�H8�Kɾ�,��1s�H�ӽ�_޾�6��p��8�?|�F?�<���UQ��0��N�� ��+�V?ç	��������2i�=��n��<{W�>�q�=�k����.��K���)?��$?�#��xm��j'>J}�[�λ��-?�?/v�מ�>}?\ G�bDw���>-r>|g�>׉�>)~0>b���h�Ľc�?m�I?� ��×�(�>V;����T��pE=/~�=��V�SD��nK>�
=ןx�:�?;ThȽ��=�W?�7�>��)�S��7Ə�.��.<=2 y?i?��>x�j?}�B?��<�Y��g�S��L���p=x�W?ui?�k>����WϾT�����5?��d?�)N>��h����!�.�L�Ur?uZo?��?�-����|��̒����:�5?��v?�r^�cs�������V�*=�>�[�>���>t�9�l�>��>?G#��G�������Y4�Þ?��@m��?��;<�!�>��=�;?�\�>��O�-?ƾ�|��������q=�"�>����Zev����4R,�=�8?���?P��>Γ��ǩ��	>���lά?�x?.����:ǽtE񾷨���!���,>﹉>a8>e�;�Q�!'����㾀1�8�ʺ���>L@�n���?��{����ɿ(�g�{��D(����?�2�>���=���=��!�ʠ����P�?���3t�zE1>��u>���=��T�
Ό���8�@�8��m�>?�:9xA>}�������wȽ��>8�?,7�>�xC=:U羸�?[�!��Vֿi�����⾙/�?4}�?VqP?	��>?k�>B��B1���lU��N#?�x?|E?�->���H�;��j?�Y��iI`�_�4��0E��BU>E3?to�>��-��Z{=��>�~�>��>M/���ĿKԶ�_���
��?}~�?�d꾓��>�~�?H+?^�[8���I��{�*������(A?`2>`;��4�!��2=�]咾��
?C|0?|��E��!??��a�W ����I����r_�>A��<�D��G>�����=e�	(��H���q�?G7�?��?�� ��"��e?l/�>��ƾ�����=�r?�>�_�=H>�|>+���~i��'�>*+�?�]�?�e�>]���䧿m>)rx?[ζ>y3�?���=���>>��=F4���q�=�%>3��=�H�f�?SL?��>?�=��1��f/�3F�E�P�_c���B����>��a?BvK?"�^>,ж��1��!��>ʽ=�2����x#D�� �0R߽:�5>�BA>I�>6�I��sѾ �?#k�@�ؿ�h��{�'�,%4?S��>��?����t��H�$._?eg�>�6�B+��W#��;X��?�@�?��?C�׾�iͼH?>H��>M�>�uսD���Z��3�7>$�B?�2�C��i�o���>L�?{�@\ٮ?�i��>����i���g�%(�\o�_����?7Ϛ�t�
>�] ?ʀG� �w�x����wj���>���?w�?��>MX|?@��aAC�H�]=Zޟ><f|?4�/?��<�����9>w� ?M��늿.:�㟈?��@�/@*6P?������׿>��#����S��A��=���=k$/>Vn۽ ��=�|6=<"6�_�m�=1�>��f>�p>RYQ>�S=>~T+>�����R!�������qC�g������Y�H�Mps�����������X2��+���j�����P�i?$���U���=��U?�8R?uoo?f��>BRz�&z>�>��B��<�E#���=�_�>��1?�L?�c*?��=�Ϝ���d�A-��lէ�m���=�>�JH>�D�>���>�̭>�CZ��,J>w�=>V�>V��=Z�%=�=�&O>��>N��>��>�k;>ǎ>�Ĵ�`7��'�h� %w�˵˽T�?�i����J�7)���M������v��=zA.?�>���H7пe�[>H?��\�.�+�n/>��0?XW?��>���6�V�r�>P��S�j�4>^E �S�l���)�``Q>�~?@f>��u>�T3��d8��P�K`����{>+�5?�1��a^9�h�u��{H��lݾ��L>ӱ�>){9��<�g��~��i�`
y=�:?}[?�O��Jﰾ�Su�A��vXR>�[>��=/��=R2M>�?d�t�ƽ��G���1=[��=�y^>�p?Z�=vd>n��>�g`�j��H��>2-I�����V�<?�`Z?6)>�qe���Ѿuh����>1>�>>�	�I1�=z�[��<�=2_ ?`�>�d��X﮼4)��o�C�N:>��=]�y�d\o��=w>J�YI>E�D>
G>�ӷ4��J>>b?٥�)���"���~u>��J?�	�>5.>�&>�"�"��J�c����?e @��?�(���G���?�wq?bw���<f?�+�>0]�����Ż>RÉ�	{վv?6��䀽��?�|�?|�3�ά����Y�U�X>�w?�_��}g�>cx��Y�����6�u���#=���>k9H?�V����O�O>��v
?N?�X�稤��ȿY|v�J��>��?B��?U�m�@���@�A��>��?�eY?�ji>:a۾�UZ����>�@?�R?�>�7���'�D�?�ݶ?J��?"�H>l��?^�s?�7�>��u��o/�\��&���Y�=w��;�:�>��>z��%\F������S���bj�Ih���a>~#=��>�W��?���ص=~(���է�A�i��>�
q>E�H>KH�>�� ?4�>D��>�X=A����
���m��{�K?���?#���2n��L�<��=8�^��&?�I4? n[���Ͼyը>غ\?l?�[?�c�>8��J>��1迿>~�����<��K>4�>xH�>�%���FK>��Ծ�4D�mp�>�ϗ><����?ھ-��&U��`B�>�e!?���>gҮ=m� ?Ϝ#?�j>�.�>�_E�9��V�E���>��>�H?��~?� ?ι�W3�6���⡿��[��+N>��x?�P?�ɕ>����;����NF�/I���k��?Fqg?�I�<?�.�?�??j�A?=f>���#ؾŎ����>�-!?���A�v�"��<��?Y�?���>'f��"�ڽ��8��ի����?�U]?�"?C"��]��������<J�8�:ޢ�;QO���>ǒ>�� �=e\>���={�r��B1�w*W<���=t[�>���=<�>��臽t&,?��=��̓�R#�=�xr�KqD�_9>RrL>N�����^?�L=��{����x���|U����?���?Ze�?Ct��\�h�:=?-#�?�!?�>�v�޾���"w��ox�'h���>i��>k o�4�侾���,����,��F~ƽ:�Q�|?��>�U?M��>��'�7�>�5�����A�ǾE��9~U��C$��\5�sW	��kᾞ�n��d�B�=6߾X�����>�)��ݞ>%&?n >�}}>L�>�Ƽ;�r�>�oD=c)O>^�`>ai0>�8q>�63>���=ehɽS;?Ѐ�R.*�v@��n�ν�W?��'?);C?�E��s��l� ���?��?� �?�'i=Ao�2,>� ,"?ә�>�I�Sk�>T�I=�H9=�4H�z������L�=�^�=3��>kl½�S�^rK�����S?y3�>�EN��=
� �>����Go= >�?d�(?� *��Q�ۧo�p�W�	
S���>h��f����$��p��ꏿ
^��,-��|�(��*=[�*?��?���l������k��.?��-f>Z�>�'�>-�>N�I>��	���1��^��B'�����.��>�c{?dG�>H�I?��;?bjP?�!L?g$�>!�>l%���6�>8��;\��>���>CM9?��-?F0?�e?�Q+?�,c>���5��דؾ�?�c?�?�?.�?����N½�O���h���z�d�9�=�<��ֽH�r�/U=�*T>E'?O_侇�W��<�o?uqB?G.�>�DC?x�w>!%�uk�^����:~>��4?�p>�4v�P��� ?�\�?�p��V�=�>�):��+����r=u����g�=�E�+N0�y,�<WX�=!`!>a�j�\1����<���<�SG;D,>��l�>Xb0?�Y�>�n�>;�"��t�>���,w=�k�>c�>0�>0�ݾ�苿���O�l���]>x��?ó?Y�/<���=�>��m�<�ľ�F������$�=F�>6�?�O?"�?��F?�c?Ԩ�=���ߒ�������? ,?���>���%�ʾ2�T�3���?�[?�7a�����=)��¾��Խ}�>U/�-~�����D�P�������~����?|��?�,A���6��k�!���
c��#�C?��>�Y�>��>��)�&�g���;;>ҁ�>;R?״�>�V?�t?�[n?�c<>��C�ɪ��k���ɛ�S�=��;?��?V�?j{?�f�>lI�=4o8�}�ƾ�����s׻�������=��q>�'�>�>�%�>���=�$��Φ���u�,��<W�>~��>��>��>|:�>l�s=.W(?d}?̪���')�����WS��7��w9|?�[�?�"]?�l6�qK�io�v��_��>:�?m��?�j�>�ɏ�8�U�A�=��	�,~���A?���>>��>h�=�1�>�w=���>���>�K�g��©p�w/%�vn'?��G?+�=F	ƿNp�̝o��}�����;�����:d�؉��6�Z�9�=����91�o���b]�S���Qb��]w���r��_/}�xo�>܇=�X�=���=�ͥ<�Ӽp�<��M=f��<�=�d��Cx<��7��ϻJ���>����5<�uT=�|e���˾wq}?ɛI?ч*?��B?~y>�>R�A�v��>����)?2�V>��T��8����;��Ԧ��h����ؾB׾�Ad�㬠�3	>�I�J>D|1>��=�K�<���=%l=��=9%��(�=��=�:�=Ҫ=01�=g>1�>U�W?'�~�>T����k��B��3?���>C�?=�l��fk/?�;>3�dB��/;�x}�?���?� �?���>$�����>����w����<���=3�O>�{+>M�2����>��W>3�?�����/6;�!�?�Q@	�/?(ȋ�Yqֿ���>W_7>��>�qR�^?1��<]���a���Z��w!?);� �̾I�>�W�=Ţ޾��žF&/=�5>�b=pr��[����=��{�kg==a�l=�׉>hmC>5�=ꌯ��L�=[�H=)��=0�M>�ј�V5��(��2=Sq�=g�b>�K'>�I�>s?��'?�Uf?�o�>����AվO󵾫��>ߢ=?=�>�l=	�(>�&�>�<?M76?�>?�B�>���=�ΰ>q_�>��+��k���p1���=&�?\��?"��>׏����u�B$�5q6�*�t��?e ,?L?���>�I���߿"��ɬI�]��V�=���<[�{������|�BF�A�F��=y�> ��>�0�>���>w�p>��~>��>���=q�d�>S����༜��=B�=i"�=������3��L�=�?�;��2-�Yj���2�<�a>=�a�=J�>Ec>lj�>s�&�U͘��`ļj{�R�f�>n��hN��,�?�w<{��Q�m��<�%>g�{�zvƽ����d�0?!�&>Ӧ!����?�r?�r�={�nϹ�������D>��3;F���l>�������{�������ճ�h��>H
�>��>��P>i�8��Z8����;Þ�
�G�	?{��8Y�=l���s�a���E���y�Z�z��*6?�����>H>��_?{6?��?���>���Y̾�>a��6�{��b��x�!��<�p?uF?�i�>�þ�D��O��q��7U4>gl����o��g���gF��e��Y�_�-�=>|{A�o�Ͼ#`.���x�Y��WG�����;�> �G?�z�?P�׾,Ey�����;����!����=D2?s?`t�>�V
?;���ث���"k��x�=>��?R�?��?�u�=z��=�������>}�	?���?�P�?�ms?�7����>�;Y�>WY��v�=��>�i�=5��=8	?��	?�s?˽���������0�]�o�=��=���>��>�p>�=(�]=�`�=��W>u�>���>P)c>^�>��>�½�Ȃ���G?�َ=�Y�=�P�>9F>A,���  ����=	T������6ߐ��G��� ;$�E>��=p�=�J�<[��>O������?G�=^���8�?m��[�=�Z >K'M=O�!���K>m~p>	�-><ǘ>' �>N�?>>6�>�(�<�8��y >X����M��Ex��2K����E(m>nӌ��㕾�E���8�V�o�þ��.k�fj���<�!����ĉ?m\��M�M�d��@�P��>��X>�?���޽k��>+n�>g6N>O��፿O׀�Y�;�w�?���?�&>>�y�>�Jd?��?��K�k1x��^]�$|g��8�zY�G�Z�����IF��J�9LA��?c?*�q?�~??�ۡ<Y�z>�,m?Z?�{���2o>�&��u>��P�=6ݘ>�Ⱦ+�j��1ʾإ�"I�BbC>��g?:(|?O	?A�{��@�V�>�,7?Q�0?�)t?�M2?ġ;?r���$?��2>(�?k�?��2?��/?i}
?�G">���=��:ƀ]=�[��y�����ӽ�)ýE��J�F=�m�=v�<�r_;P��<k�<n�ۼBSļ�fֹ,P����<�$8=�f�=�o�=�e>�?��>����b?���~!>�|%>�;�X?WL�>-�	��ؾ5�$�/�<������J>?<4�?|O?�;):S���������>z��>(�+>K���{�=����g=���L=�b�=ͩj>?�>i�ɽ�i�����þ{">�4;=��>+��>�J�P�G>����0=��Xg>��E�W\���FT��N�:o3��z�m�>$RQ?ږ?i�=P=�ؠ�Y%m�5&?8"B?��J?��{?�聼"����7�V[D�N�轩�>b(<�#��d��񾜿�W*��B�<��{>`���[���I�Y>=�
���ܾ�5m���B��5��tR=+���w]=�(���Ǿ�c����=gI>ң���������벪�I�G?5/=2F��OQ�.���¤>�v�>���>��!��B����B�Up�����=Lt�>�:9>��?�&㾉�=�ߵ��p>;?u�p?.(o?�躾;��D�c������\�8>�4?�r�>ҳ�>��='��=zh�e���C�>���ˣ>���>g�+��8@�h���ל��R�_��>�|�>��<ã$?��0?��?"�E?t?�>�?aY�>����l���%?=V�?!��=�hԽ�2W�}9��vF����>�_)?NB��,�>(1?��? �&?	�P?BC?��>���M@�_Օ>���>��W������^>��J?b�>��X?���?��;>��5�f��ot���\�=��>��1?#?�?jz�>���>�P���=���>F b?7�?�p?��=��?+�.>LM�>��=s�>Q��>��?��N?1t?t"J?c@�>y�<�|��s��3*g�8�6��Т;��,<"��=>���l���%���<hm�;i��K�k�����@>�``��g��;�)�>�n�>����.�=�~��Tf����=��j>�h��b���ڟ���˽4 t>?r(�>	n ����=��>1�>�L���=?t��>	�>?�k_���C�#kо����l>>�N?є*>��C��W����v�it<�Jo?QR]?�˾[��:�b?��]?1h��=��þX�b����Q�O?�
?��G��>��~?b�q?��>��e�:n���Db�:�j�Ѷ=]r�>AX�E�d�m?�>x�7?�N�>a�b>%�=ru۾�w��q��l?��?�?���?C+*>P�n�[4࿘w��y=���^?��>7U��#?�����Ͼ�Y��(:���z���뫾S#��^u����$�2���t�ֽx�=u�?0s?yVq?��_?ձ �� d�>^����uDV�x&���B�E��E���C�:�n�I\��?����|vH=b��/��8��?���>R�`� I.>�f�m@�h�8���>�ɀ��	��Z�=`T�<�z,>M��=�(��j����
>'?dT�>��Z>�GX?�xn�Üa��#Q���5��@I��>J?F�?[6?�	�N꿾�f��梾�&R���!���t>r
c?#K?7m?�8���1������!�G.�!��u�F>��>I��>$vX�����%���=��Vr�5N��!����	�ƭz=f1?O��>A�>��?�?J:	�+T���{�s�1�곋<�@�>�5h?`~�>I*�>,�ͽ,G!�7o�>��k?��>�(�>����8�#��+|�bG��e�>�˷>]N?zCq>�7��	\�DЌ��[��@�9�1��=�h?~Ĉ��\� V�>�,P?� b���$�cw�>�Z�l�$�2���K��đ>�0?���=�H4>����	���z�iu���@)?�*?ْ�]}*�S�}>�0"?�L�>,�>#�?�>�Qþ�=��?f�^?f	J?�A?\z�>�4=Q!���Ƚͺ&�x�+=N��>�Z>�tk=��=C���T\�>*��E=�M�=o�Ѽw$����< ��F�M<���<��3>k��˙M���k��:ľ��e���憽T3B�޽-⫾�Z������Z5������4F�.5W�^ZX��=T�oF�?.��?�F���P��3ht�<���y�>^�[��L�=<Ӂ�Oz��鍾���MD��_�?�`c�8�]���>�O_'?2����$ȿ�B����ھ��?�$#?Lz?�1
���!�:�:���>���<�c@8r�ྒ���S�Ϳ����E�^?7��>������@t�>��>�NR>��u>(W����)�<�?|w/?!{?��a��˿�컿_2�;�w�?8�@dF?�\��zҾ�?>��v=@R?�_7>%�����b�[S��n��>~E�?�nm?kv�{�9���>�?�����#A�g�(�c+\>�W>7�?�����o>`	E��4-���B���<qF8>ʔ>0�<y����৽�R>��=�J��@��yф?�\\��f�g�/�HG��HY>��T?is�>G��=ݠ,?�AH��Ͽ�\��,a?�2�?ڟ�?u�(?�ѿ���>g�ܾf�M?06?"*�>�t&�խt�9��=���腦�u��
V�I�=j��>x>��,��r�s/O��C���t�=�h���ſ�D"��C�%�L=�\</�����彸r����b�,����q�iO�|=pf�=�iS>}؅>��[>�rV>�s^?�@q?H��>�>�]
��А� sӾ���;dq�{���
���8'�S~��[�쾟���F��G�����;8�;�ݢ�=ČS�������#�o_��8J���-?�@>|�þ��H�٣;<y�Ǿ�*���;��#��Reþ��-�&�i��Y�?�KB?˶���U�6�-��� ݦ�c�Y?yn������N�=6zU��iL=�> �=�#ھD�1���T��+/?��?X����?����>����{�<?�'?���>V��<\��>�%$?�N �"�߽�oV>��(>բ�>���>��>yA����Խ�?��T?'��㢾�>JD����o�ǩ�=6�>�3�w�>��2[>>
�<f����Ļ墽@��<�X?���>���i.�3@��*�=^�*>ƅl?�L?|5!>L%D?lL:?c��=�%¾�Q�"%���="�Z?էH?�3>��wj;\�ʾFa?�n?�}�>ݦݽ8j��xQ�wB�ip#?��P?�S"?^}K���q���������D?��t?E�]��������ɤ_�x��>�1�>m�>�8����>�1=?�i&��Δ�y���3��C�?�X@?8�?+lM<�N�ܒ=Fq?��>�+Q�0ľ}���uͰ�r=i=+��>�X��"uv�����(�g;?EP�?M ?�y��@"�Io�=����]�?��?Z�����T<<�.l�����H�<���=��.�"�����7��ƾò
������P��h��>A@�H齓q�>n9��6�HHϿ��cо1Eq��?R��>�Ž\�����j��u�\lG�E�H�����D`h>��s>�Ԡ�E;Ͼ�ۏ�:���O����>R[>s>>>d����7F��a�<�p�>�.�>5�>p.>@`����? ����⁣��Ti�J�n?~��?<��?�a�>�������	�$Æ��Z<?6�N?$�5?E4<Cץ��ӝ�[�j?�}��?Z`���4��=E��U>u%3?aJ�>Y�-��b|=&�>O��>�>Z/��Ŀ�ֶ�9�����?���?�d꾳��>���?w+?�d�0���f����*�����P:A?Q2>�g��J�!��8=�&ݒ��
?�0?h��lH��=?��U��ъ���N�p����o�>h���-�=��^�u�<��x��ҕ���J����? P @.�? ��t��?B;?+H��������=v�?��c>)�>V�Ƚ �>�y��)I�=O>2��?�d@�w�>Uꗿ�����[=�Qv?%��>��?���=���>���=퍯�����F#>���=��;�?|mM?���>��=i9���.�M E���Q��c�YD��ڈ>W=a?�/K?&n`>aḽis+��B!�G�ӽ��3��i��A��&�V�ڽ��4>u�=>U�>��D�.�Ѿf�	?����6ݿP���@�~���0?�%>f�?��:"(��V˼SkL?��o>���-���?���ĉ�gl�?�~�?Y!?١˾����$�=a�>>��>��k�m��i{��+>�3?�m9���o�J�>���?�(	@ω�?4g��E�>������]|�t���n���_�;?z�ھ�͒>V��>��<uj������c�'�>��?���?�m�>��^?�lR���%��%<JLs>�a]?D?���=T�z:=/k�>����������e��?1@�@԰B?/��\>�����9��׹�����<DCs=��H>��<��T�;�ș=����Ñ�k��=���>_��>R�>�T>���=%3>w���4)��򞿩����A�"��e� �@�H���=�r��X���N��O�e�M"�<���������h���;�h�=��S?P?q�p?���> CB�,b->sd����M<�&���w=m�>R+2?E+L?��%?���=E��2�a�Ⓛ�c9��m2���]�>�8>J.�>E��>��>#Q;�^|J>�->�;�>���=9>[=½I<Y�=�L>���>��>�"�>B<>��>gδ��0��J�h�ww��)̽- �?Մ��v�J��/���5������id�=b.?�z>����=п!���H2H?/ ��I)�Ƿ+�-�>��0?0gW?�>�����T��*>X��ʘj�^p>�' ��l�܌)�(Q>�h?�uf>�t>Wq3��8�Y�P�AU��{>6�5?5X����9�fdu��0H�Iܾ�M>7,�>~$W�i��dϖ���Fi��z=&:?{�?6ų��s����v��Z�� 	R>e\>��=��=�>L>�oa��ƽ�G�=#0=���=S(_>X�?�^�=NCf>6�>�.=��L���h>�s���3�>��?$*V?�>=G��)��V��Z<�>ْ��Dނ�N��>K9���@>:��>C�=��ٽ�
�I���M����>׾�>S^ý/1������%i�E�>$w�~����5;>8>�q?������3�ݾ�"t��J-?@42?��_>6)�=[o�U�������n��?��@��?���5[�G&?a��?穌<'����>�?x�:�h��}D�>�1r�B�˾�9�t��;Tϴ?�&�?8����a��!f�Y�>L47?�#��N�>hI�{L��� ��"�u�rl(=���>�H?������R���>��T
??/��T����ȿ�=v��+�>���?��?�m��1��G$@�/�>���?�xY?�Sj>��۾�^[�/(�>�@?��Q?��>J��V'���?5Ѷ?f��?��H>���?|�s?|D�>��x�h/��1��������=��y;��>�H>�����aF�bē��[��r�j����	b>Z�#=�*�>F4�8`���>�=�~���$��[Af�B��>�p>`I>2<�>0� ?j�>]��>��=�c��gˀ�7����K?6��?9��2n�`B�<a��=6�^�'?�H4?4�[���ϾԨ>��\?:?n[?�b�>���=���翿&~�����<7�K>6�>�F�>�)��|CK>��Ծ�4D��p�>�З>�����@ھH-��ev���B�>�e!?���>�Ӯ=v
 ?�u#?�\q>e��>ƝE��䒿�F�9B�>��>|�?:?~Q?ra��*i3������Р���Z��$M>�Qx?D0?���>�s������`�l��h�D���#l�?Md?�-�c?婈?�@?�r@?j�^>���Ծ���#L~>�"?�����8�2�!����#	?���>��>8M���!���nI=@������8�>�N?d[5?3)�Y�a�(鞾�5=���r�";�5���t��M	>�>�e���=�Z>�>�b��Jx�Qn<c��=�K�>��x=A���w>�~:,?��F��σ�I;�=��r��sD��>aDL>o���ӫ^?Eh=��{����su��r�T����?��?�h�?1���h�{%=?��?�?F�>H��|u޾��ྮww��~x��s���>��>��m�a���������A����Ž���WU�?{)?�?�'X?�̛�G��>����.�ğǾ_�$��;���t���C�f�>+6� �Ń��
m�>����a�b�f6?,��g�X>���>`�.>����j>��u<�g�>)g�>�C�>�>��ϻ�Ā��!�󋡾b�S��9h?[oM�,�
��>���?d#?>hX?�	^?ޖ�>�륿��E�?�=�5?`ܹ?���>�Al��XE�G	t?�c?�A�1c�>[Un��=Q>+� >�澁=��RsZ>,�;6ط>�'�[�s���M�_���9?sU?����]��NM�>wW��u�q=*b�?��(?b�)�l6R��o���W�ەR����g�����[�$�mmp��Ə��&�������r(�]*=��*?��?_��@��0}���^k���>�p�f>���>J�>��>�J>Ѝ	���1�?^���&���?��>�z?v��>�E?X�5?f�[?9?�=�>���>A����4�>����>�t�>�w4?H,)?�_?��?�97?�b^>8�7�����m���?=G ?�y?[��>�u�>���H8�����l<1W��|
��8��=g�=�ɽ�(���+I=�;k>i�?}Cj����)��uǂ=��J?׮?��>����4k�5TP;UA�>��(?�l�>�־�X~�9���J�>0�$?�����<0M>�h%>��=�;����=���=j�=�I�<�x��������=^�<���;8V�-틼͇>2=c<t�>�?Q��>E�>UA���� ���/V�=�Y>�&S>�>�Cپ�}��B$����g�J^y>v�?�y�?��f==�=��=7|��8U��V���������<��?LG#?�UT?ݕ�??�=?�j#?��>�*�%L��{]�����q�?�!,?M��>�����ʾ�憎h�3�T�?{P?@-a�����2)�D�¾'=սϠ>�Q/�c,~�����D�s���@���f��\��?þ�?jQA���6�S��Լ��Y���C?�!�>V[�>`�>Y�)�S�g�y"�u=;>p��>�R?H�>d�?�]?��0?�<�yg�Xd��[�|���T-+>
2^?��|?"�j?�5?=�
>�
�>3m�=���{�
��9���&ξ��=�-5>8�?ԟ?���>yP�='܍�"@��ڻ���w=��?w�B>;~�=�^?&D�>�3���F?��>$���O�d����SB��9q?�6�?�'?�UG=R7���C�=����>.l�?c�?=�&?��]����=l�ؼ@���JUf����>F>�>�n�>�%�=�=I=��>"'�>떿>��������:�'m^���?)�D?{X�=+iſN�p���i����Vv<�����^d�𾕽\�Z�c��=xܘ��E��I���Y�F�<����״�#L��z}{���>�(�=8w�=���=���<k ּ�<a�?=o�<0n=ֲr�;�<�$��ݘ������hY���^<�
N=��6�ԫ��-�?%,s?�x ?\�i?�E�=�rh>W�����>v���o�>q<����h����EV��ݾT���l����-Y�ʨ����#>Jɼ�>x�F>��=B��=��>��On>���=M��=�">�P	>�p->a� >�W8=�G,<�v?�N����tQ��j�y�:?�?�>x��=�%ƾ�??5�<>4,���1��Ǎ�oR?���?�3�?��?�<h�z5�>�񢾞2��f�=,��
�2>k�=N�.�d#�>�SE>�V�����v���W�?̧@+�??Vߋ�)�Ͽ&/>7#3>e�o=��@�����A������վA�?�R��¾��>*x>u  �㕐���Z�$==��>���k�g�z��=��4Y����	>���>M�m=�q>�N���NH<jλ8,*>&
F>|�ȽbC�<X���?~=�1�=q��=� �=�9�>V%?�O7?�sV?9�K>�p�N���z��K(�>�<L<�!�>Β(=Cǉ>~��>]D%?��$?o�:?]��>��;ɷ�>1��>H/��,_�=�U��٬�<�?Ҕ?��>� ��Vx�4+�d1-�糡����>�� ?mo
?�O�>����:�C��%{-�K������)�Y=�8r��q3�!m�A;:��U	����=n��>��>ٙ�>ꪈ>�L9>��T>1L�>[`�=�䃻�R�<3.g<T�O<򆎼;�=Ra
=)�~<u�ͼ�����N;����;ч;�B�<|�=$B�;��=�
 ? �>�>�_=�na�Ȳ�<x`���#�h\�>C��ux��9W�D�`�ĉ�����#[$>ui>S��Z����?�
>�ެ�ya�?�<x?)@�>K��)d��ۥ���ľsLz�4�=UJ>Ҵ�w���<��6'�����ua�>��>�*�>V{>�b.�ޣD��u�<�t���#����>~l���ۼ��4�4Mp�����Y���i��A<�bE?m������=	�x?��D?$!�?��>���Ⱦ��=1���u'n=�R��/�x��-�?n*?���>b��{*@��tؾ��۽�_>�	n��X������45�J<�������>�6��5>ƾ�+�����/؎��5H�����ڞ�>��P?	ͭ?{:i�7邿��D��W�!|��H�>�!e?��>h�?5��>�i��ެ޾B���ɕ�=>En?hd�?���?b�>��>�q����>��)?c��?�ԉ?�n?x�
�&��>,1����&>�Z����=�f>�]��*>��!?���>)��>L�U��<�����¾�I8�j�_=ѧ��⾠>|�j>%��>��<@}a=��=Bm>��>%ou>`�n>z�>�Z>�ξa*���O?��v���y>[��>��>ǖ��(2����<����fk�r���^^���
>#�>�f����=t`=�y�>㻿^Ģ?;e�=%Q�Z��>l�پ�t��z)�>�*���D��#24>�ǰ>h!�>�f�>���>��>��>Θ�;���~R�=4/��#���J�K;��
��o~>Е��>�ٽ�o��|U��Z�����	u��q�����/�)��&�=р�?�t��Z���u�&��7���w	?jH�>V�/?�}��U�=��=��>d*�>�$���)������:ݾ{�?���?Q(b>Do�>��W?G�?8�2���1��Z��mu�u�@�oe�wt`�ѷ���>���
�#���|Z_?l�x?�A?��<'Kz>��?�^%�M��^��>Y/�t�;���:=ȥ�>@M��9�`��ԾX�¾!��pG>�o?]��?-�?�%U�&�X��(>Zb9?Q�1?>�o?[3?��=?p[�[v?��0>#V?��?�7?�9.?Y4	?e(">���=r!��m~�<�����~����Ž�Ͻ��;��?�(=��x=���;��R<��=AԀ<K3��}ȼ�ߑ:d����<p:=�Ƶ=[G�=C�Y>��v?���>;�>`gI?bI���]3=���+?iϗ�����#�P���zҾ��=R?Y�? W?m�>�k�R���B�>#R>��r>��>�@�>�D��]���D�=�ݐ=��=Il�`"��(d�����D��l��=�=>r��>�4?*�v��J�>٠*�N�i���6>i]>�K⽥����a��yu���޾d�>"Kt?�4?�լ=t��Q">��i���A?;N;?M�;?��T?���Ʒ��-p�t�)��xN���>	�y=
�*��¡��[������TV>��>{~.��⠾=-a>*��A�۾߮l�rYJ�����M=V*�(�_=�L���ҾMQ{��3�=��>Qd��x��^��,+���L?4W=���]@c�D%���>�>���>}�-���_��?�鬾��=֯�>�5>N7��p뾭_E��!��9�>2WC?��e?���?[_����x�>E���~��O��2�?ޕ�>�M�>z�4>���=N�������`�/�3�� �>&��>Ll�O�D�9U��D�羪�a�>f�?:Z�=�[?^L?k ?$V?_�&?�?�O�>�"ս����;�%?�ڂ?wě=hW���M�8:�PF�Я�>B�,?�VC�i�>�?��?	D#? T?"d?�+�=Hs���<���>uT�>�4Y�F����n>��M?ꭷ>��V?~��?�(>��5�ș��Z6���i�=�>�3?��!??��>�Q�>G4���vb=�K�>�
h?���?(�r?�G>�e?��>���>d�=�0�>�>�?�M?�v?��@?F��>�qD<b�����Ƚ&�b�q��a-ѻ�Ρ;ѓ�=z�ڼԛ���j�Y@E<���<��5 ��p ��8�m��Q~�cy�>b��>j禾���>\Dʾ�2���_>���;��ϾY�dn�n6D����> �B?��>3�F��s�=vl?R?B�a�ӡY?�
m>��?	�=(L?�<>��\>��,�n>wi??&=�W��Ć���Q��f�<K�j?�j?Z��
�i�b?��]?sV��=�$�þ��b�����O?�
?��G�h��>!�~?��q?���>�e�4n����&Bb���j��׶=�n�>�\�p�d��O�>�7?�P�>��b>�#�=Ǆ۾j�w�f���?��?���?���?�+*>��n��4�����P��j�]?9�>�����!?����pϾ%��`������n���`���P7��Hͥ��n!�?�����н���=�E?�s?1,q?��^?$� �toc��,]�l���T��i�ic��)E� E��ZC���m�T��H��ӗ�NNB=v�g�C+��Q�?@?�m�����>��þ�A���ے>�DM��)3<�=��
����=A	�=n�a��!�������1?��>�P>�qY?dT�ۈ/���,��:��6پ+�>�?��>v7U>6d�5�C���=�'����
�m�=B �>�Z?0N?��f?����g�7��bu�!!�=�'>�֡�߈�>C>X>��<1z�p.�=2��G�Z�k���پ9�Q�&"���ĽI1?06�>���>~��?��>�4���Ծ���������9>��R>�?1?�?��>4U8���#���>�\k?tx�>sq�>����}�"��|�o�Ͻh�>Y�>�<�>��f>op0�$�Y�����N���8�(�>�Wg?�k��l�^�҄>��P?����<�͟>�ӌ�H'"����&�'�d�>�0?�x�=X�E>w�������{�g����*?�?�7��7?��٨>��#?��?�-�>oqz?��r>�PȾ^�;=^�?��J?�+8?0�=?C��>H⪼����qֽ�j1�/N�<���>|�n>�#�<~��=�R��0�?��8B�'v�<1K�=��M<7䁽砼��D=�5=�J>�'����P�mh�K"��{˾���:����������D+�`���;��	�������ʼ�O7���K��S��<��0@|��?^��q���є�U�a�(�����>5�`��%����v���w�o�eѾ��G�8��fc���7�B/���'?������ǿ/y��BMھ��?_ ?ARy?8�T�!�%X8���>��<���,��W�����οp
����^?� �>����������>��>8X>H�r>;'��l���fi�<]&?"0-?6f�>c4r��gɿ$\��d�<��?j�@o�,?�>�_������Q�>�}>x�A>-���������#^�>���?%s?L����y}���>��*?�Xо��[�!J�;�h>��>��r=xݭ��F"�ւ�������X���=?1>�B>��ǻ�-��F�W}�=�>�=�=ٽ�M=5Մ?,{\��f���/��T��U>��T? +�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=r6Ἶ���{���&V�}��=\��>d�>��,������O��I��T��=��	��ƿ����"��k=�<Fs�?Q���6ս�M���J��1\z�"��W^=�z>��^>�/�>&W>��Q>y�h?��n?���>xc�=��U���	侴f)=�ۜ�Y�(�"P`�b���Z��݄�*��J.	������
������=��ˍ=�4R�I���.� ���b���F��.?��$>�ʾ��M�1�*<��ʾ����)������D̾{1���m�ԟ?)�A?w���V�������v��[�W? (�B�����=�,���=N�>3�=��J�2��XS�ڐ2?���>�)��s���>�%��c3>�?W~.?�>�/>r��>�X��ʩ=MD>��=>x+�>�7>/p����!�ī?S%p?��޽@㱾���>o���s�w��]��0�X�T���_}p=��>�t��X����F>5�9>�ћ���V?ز�>�x&�r)�5���,�<�ؐ=roq?^v?�1�>�9d?YM9?9'_<�򾯶L��'�ׂ4=�N?a'd?�@ >����־����m7?0�g?�Z>C傾�!�3��S���	?��j?FO?�  ��Lv����� �ʰ6?��p?h�\�][���	�Ԃ|����>�)�>�2�>L�>�`�>ߐ;?�,�K��콿�.�x��?��@2�?U�<kE��"~=g�>ҿ�>�7-��Y;,���R��Ja�=3��>{a���]y�z@�����H@?j��?��?���f�����=8����? (�?<I��hi<���Ql�����{��<$��=� �kz�*���7��LľL�	�֢���r��*`�>n�@	��O"�>t;�*Cῳoοj�Ͼ�Bj���?Ъ>K۽ 3��ni��cr�L�G��wJ�+���v��>|z!>}j>����xe�,�a����?��=�&�>$�f�Ɇ�H�(��GC<�yS>�b�>�Z�>�������0�?� �Xܿr���8�о��?IҖ?��h?��?r~_��Ƚ�A��Щ�E��>��C?DIY?���C�!��E�=�j?�_��9U`���4�HE�|U>�"3?�B�>~�-���|=r>w��>�e>9#/�=�Ŀ�ٶ����_��?���?�o꾃��>N��?ts+?�i��7��[����*��Z+��<A?2>����!�0=��ђ���
?S~0?;z�Q.��-H?�Od� ���'���=G� >r�k�M .>0̧�IK��O^�QВ�"����;�?U@Vz�?7�!�W�(�Wx?f:�>[*�v���qe>k��>ͮ>�)�>�/�u��>��%�j�<��x�>��?l�?:?�J���+��h�e>V?=?n�>��?���=v.�>���=~����� >\��=H�8��?rVM?j�>%�=��7��-�ēE��$R� ��L6D��d�>�ha?�<L?��`>����93��� �c�ͽv�1��b󼡽?��q*���ܽ`�4>��<>�G>pC���Ҿi�?��hۿ�+����s��x:?�2>�'?���\�~�CHл)KT?��Q>�!�\䵿S�����7\�?�-�?��?����v�](>tDv>H��>�5׽=�e�AN��D>�??`�ő��Op��W�>�q�?[Y@�+�?Lh��u�>;h��蘿�����H7���;����9Y?�%��>���>�@=<t��b9��n<j� ��>�^�?��?��?ED`?�i��+?�}$=�e{>��O?���>���Q���$>p��>��#���������&�?	@��@�iG?	-��g׿���&ܴ��������=���=�q7>m[ѽ���=\�;=�3p�󍬼"��=��>Ѵj>��o>d=P>b>>�<)>:l���]!�+���V��e&C��K�~\�4bY�#{��)q����k��[���$d�������Q����L��H"���U��H�="1V?��R?�St?ld�>ț���j!>���{=^
���i=�J�>��(?�.>?(?�U�=�+��Z�a�w�fe��X���2�>��E>���>���>,1�>��;x_N>2�>�]�>Y>�X=�bF<ve�<�;>%>�><7�>�G�>6M<>K�>�̴�W1���h���v��̽A �?{����J�H0���9��)���Y�=�`.?9�>���0=п�����0H?_ ���.���+���>w�0?�dW?��>��HU��G>����j��Q>8. �pl�B�)�� Q>�n?0i>#Hq>'�3��\8�@HM�J ���y>-5?�C��S-��;t�^�H��� MQ>���>rf��*����l�|�	c��T�=�:?��?������xNn��E���U>�Y>�D�<��=��S>o�e�֓н��I��w)=|�=��]>���>D�P�$�>T)�>��J�r� ����=+�?��ϖ>�@O?��?��Q��x��0)v���!��[�=��(<���=5�[>���;�=���>�=dJ���cb:�Z��M����=���>�#��M�r��=9���`��=��5=E������1�=&�l?F°�b��	�ھ?ĝ��?�� ?Ob�>�6K�0�4�-���`��6��?�C@?��*���d��!?.�W?�{ �xc�a�?�iv>͖��݉���(?�M�����* �:��=���?��?���k��H���U��>��*?�,��'�>���oV��m퇿@v���M=✷>�K?4���\�uk<��9	?i?.F�N`��"ȿ�v����>|�?���?��l��\����=�;��>���?��V?��t>�߾��Y��D�>�h??g6M?q?�>]������I?�/�?�v�?I�W>8��?\n�?�C�>B�e��D�%���酿��&>�=*p�>�d>�����	4��e��w�XSp�?��#c�>{�<e�>d��?Ἶ�7>X�z����K*�+2�>c��==�>��v>5��>���>w��>q椻�Ľ�SZ�"���x�K?5��?���2n�gx�<���=j�^��&?�H4?��[���Ͼ�֨>U�\?���?�[?qd�>���=>���翿�}��Ȩ�<��K>�5�>_I�>�)���GK>	�ԾD2D��n�>�͗>����\>ھ�+��Kg���A�>�e!?���>gή=�=?3�!?�Uw>��>D�I�O�����E�9|�>ή�>̬?�_~?B�?e�����-��e���B��	/Z��Y>��w?y?G1�>�⍿�c��{��P�p�,��� ?pqf?G��8t?>ч?��9?�S<?޸t>�(��ؾϨ���>?�
?.���;�����X�<��?�@�=��I>&]����*>�b�>~
��B�	��2>�gP?E?^	.���Q�V<FH-=�-M��م�S���&1�=x�=掙>�����}�>�Ct>/��� ��_��:�V>�_�;��=�D�=��*�)j���	,?�E�'v��xŘ=�s� �D�q�~>��J>����_?��<��{�F���D��x]S����?�W�?�x�?b���\�h��S=?�?<?X��>=Z��f�ݾYNྕz�Fax����H�>�)�>�T|��<供A��[T���G��M�Ž�e�5�?n?rX?��
? �K>�3	?�=�P�����9��?�����t��L��K���J&��TQ�&�.>���ل�K�Y���?�DB�5ތ>�s�>;�F>��P>9A�>ȷ�=�Cn>D��=feٽ];�M:�F��y��4{�n &��6J?946�i���w�o���ϩ/?|�?��F?�4�����q�%�QP�>c�?��?ɴs>��h���qS-?:5�>TL��6�&?��K����=��%�)�|�9Ӿ�����޽`6�>?�ܾ�b'��)���k�E?���>�����>
���>����P�=�o�?5r.?M4�]R��"p�(|Z��G��n;N8>��ቾ�{!�ʾn�7w���^y�M����'��r�=JK+?�D�?[x��ᾣ�����f��);���W>��>�w�>��>g�>�����)�RK�<!��.�����>3��?&y�>��H?B0:?H�O?UzK?�C�>�ѫ>�� u�>VY�;�ל>���>g�5?̦)?.?��?�*?�bV>�� �84��е׾wz?��?�&?� ?g? �{��rƽ���>t�pt�݋?�W��=]q_<�ɽ]�_���R=��N>m�?��&�,i-�����O��>;�5?tȾ>}>�>*=H���w�=�I�>�w�>�mN>�Wؾ�Y�̜�u�>w?�n���= �>gC>0�=�ł����=�o��\�= ����	��k�=���=M��=�ݼ�����^=�^�=��c;sn�>(�?B��>kJ�>=i���� �����H�=��Y>@T>�>әپgz�������g�Wx>rh�?*��?�-e=��=$t�=xb��d���W2�,��O��<��?�M#?�aT?���?��=?�M#?�y>V�x;��}V���	��u�?/,?�c�>8��~�ʾ� ��;�3�a?*2?h�`�&L��)���¾e�ս�>�@/�k@~����3�C�c�����#,��4{�?��?��B�a�6�J�辚Ř�qo���yC?���>��>��>I�)��xg����C�:>#�>�
R?�*�>�9?��|?�X?p0=SA�P*������@>�yP>^wR?l q?voF?,@?2�>��4>}Ύ����_�a�d����[��w��T��;z��>G��>Q�>�*�>C�#>�MZ��s�SG�(���/�a>�<�>��>��>�2>
a����H?J��>R󵾴d��{���,!���;�n?��?�� ?�^=�n�#E9������%�>"��?x��?��?`�I��O�=#��޲ؾ�D���q�>s	�>Ў�>-vz��Š�bا=��>���>��T&���6�?sܼ��?K<?�x>K�ſS�F����H�پ P�=���������0���O>������9�r���\Z��^�Z���ߗ��@V���:�xT�>��%���r���=�=I۽�j��߄=���=׈�=�h�Υh=�6*=�r�ダ�U*>=WӉ=��=e��<�~��?�0L?k�1?M|9?._g>�r5>�h���/�>�ۢ��C?�9?>��m�$g��J�?�@���ҙ��{�پ]�ؾuw���43)>��Rm!>Ƀ3>f%�=Jp�<�>�j�<��=!��;V�=���=-�=�H�="�=r�
>���=�Q?3q�H���cem�׉���6?<�;=:Ӽ>v#�.�?�3>%���'ǿ[P����?O��?O��?��?=����>����	^����>�Ѝ>�#���!>�m ���
?-�>�-�/���R�>P�?�?KJP?|p��I�w�>�Gb>�{���YC��*�MT��o��❾���>=)�
���hx�>_�U>>��3��%	�.�m>��2=
{�D�A���J=9�ؼ5��<��=���>7<;>�Z�=C����'>TH�<� I=@�>�<!���U�ʼ�]"=�#�={nO>T.>��>�?�n1?>�c?��>W䂾�ž1W�����>r�>e�>��=�*&>%��>4�1?��5?;[E?�}�>?�b=)��>���>�M&�O�q��q��Ld��(��[��?<r�?��>ct?=��G�>���78�H�н��?�f)?��?�e�>Ua�0�߿�%��/�?˔�H�;�3=�Gp��J�~���2��ѣ彽��=fȪ>;�>⮟>7nz>mj;>�|N>��>��	>}F�<.��=I���U�<x��깃=؝��:e�<B���v"P����9.�&h�����;`Դ;F�a<:��;��<��>[�y>�6�>���������> ����["��x�>B��/�3��nB���Q��%��r���g>���>(F���ŗ�u#?P,�>>�:>��?W�X?@0�=��<�p�Cp���W`��/��M4>�'w>�cl��� �N�!�_,���ؾ�>�cw>�ާ>u�=>�;c���h��k��	X��ᚾ��4?�I/���?���k��_A���w������V�7�r>��)?MÃ��'w>��`?2d@?A��?���>Q���Pv�+�-�qq��x��!�V���н�Ms�̦7?]�.?�t�>����#�/iӾ��Ž;e|>5ߊ�#�R�֍��"�9��ʮ=����/-�> ��C�ľ �0�����[���D�!A���>��Z?�/�?Ѳk�����D��� �cR0�^�>�n?��p>���>r�?���1b���ԍ���=w�n?5�?t�?�S>�33>t㤽f��>�ͨ>T�?EM�?��K?;e�ä�>�z �Z�>�A�9<I޹��a=�N>�F�=���>Z-�>��>�p߽�0�
��L��fG�������<��>>�{�>g�w>��_>OX���?��s�>9>�y:��A>:m�>��>4B޾Ol����Y?z>��<�ܸ>i�=ը�����;��F>«��d�@(�}�<�=e�F��R=>dM�#��>S�˿�5�?��'ξ�B?���/��=�5>>�ֽ4����?糉>��0>�MB>���>J�=�	>eB=�
��{�=��%���=�h�7��.��A ���>8`����7�/���6��p~�ڨ�d���h�g��p��xO>��?8��<�2��Lb&��}���y?�B_>�_V?�Ui��i�f>�� ?�5j>���替�܈�e^־@t�?W�?�;c>��>N�W?"�?X�1��3��uZ��u�2(A��e�#�`�u፿����
�����_?��x?yA?�U�<�9z>C��?��%�Xӏ��)�>�/�';��@<=a+�>#*���`�U�Ӿ��þ�7��HF>e�o?)%�?\Y?LTV�_q����>t�(?ɠ6?��p?�?Y!6?]+)�3,)?��=��>�?�8?Oo$?�L�>�\E>-�>%��"����e�t�ow�umսr8��%=u�s=��=Q�;'eu<���<�S��
��>�<l�w�<>?=oҔ=���=]`�>o�\?���>��>��7?�z���5�o����.?�+4=5��ެ��訠��M�!��=��h?_M�?&�X?�]>�xC��B�^�>�1�>t#>�g\>��>�6���E�#-�=��>�>QA�=��?�1ꂾD������[�<��>���>�ۤ>�Y=f�>Q¾Ȉ��	Ć>,y��/ƾ� �=�J��
"�d����>�>?�&?���=�@ྞ�Ƽ=_���QA?�+?��G?D�\?�=�ɴ�� '���C�K�.�ծC>�Ѽ�6������T̐�B�0�(��=�,�>V����\���aI>��D��ǚl�,�K�b��)�<n������=����4޾O'��R�>X�>ϴ;�� ������ߩ���D?^$Q=�ߛ�O>G������3>�d�>�Ȥ>IĆ��(���B@�bt��� �=B��>F�>H��9@ྱ>�Ԕ����>�i6?��c?&��?����8���D���[��� \��v?�R�>ӹ?~>q=q<�=?�G�%i�1ij�H�z�>���>&J3�1�lW��|��&� �L��>l�>�ҹ=`/?��*?��>�??��<?{?/5
>����ު�+c*?��y?��=Ƿ�1�'�	;:�U]C���>�?��K�O�>�U?B�?��?#�N?��?j�=�
���+��֘>��>��X�Hp���ڬ>)Y?�ڵ>�E?��m?_c�=�%�{�崽��=��>q�5?W&?X?�|�>k��>�K��;�=2G�>?�d?�(�?�n?	K�=�� ?N�'>�@�>QF�=���>�=�>^]?�DO?'�s?4�D?�F�>t��<EŽ��ǽs�K�F�3��v�XJ�<��=������0����<�G�<l�M�������j<!��㍼���e��>3��>��#q�>;����!��t�>sVG>�7��p�뾞��D_��۷>i�)?@θ>�b^���\>��>��>F`k���T?���>�Y?S�b�08R��U���p�w�<"��>�-��D�\�g�u�Z�f��&���}[?qc?��v��!���b?:�]?���ך<��þo�c���2�O?��
?ֹG��#�>u�~?�q?I��>?e���m����Ob�9j����=�w�>.����d��4�>?�7?�Q�>2�b>�E�=[�۾Rpw�VN��(�?�ʌ?;�?���?6�)> yn�=��2��"鑿'y^?���>���3*"?���(о�������59�HĪ��L��)U��<��Z;%��-��=Խ��=�3?){r?Vq?�_?�Q ��c��G^�F��V��8�nj�*�D�P�D��C�y�n��[��&�� К���A=w ���^���5�?�]?�Z*�J^2=��پ�<׾ �>h�c>yi���x�
M�> �<����?���ڨ��..�gDϾ�	7?ʌ�>H+6>�
?��*�e��I���žfO���/e=�T�>��?c��>4��o�����>�ݢ����'�<��~>^/a?�L?o�n?Z��2�G�����@�l��� F>��>E�>�jb�$V�lv���=�q&s��*
��匾V���CQ=NG1?�*�>�Ɲ>8 �?1?��	�Wf���Pu���1��;SH�>+�h?��>U�>��Ƚ�>!�i��>=�l?���>��>�����[!���{�h�ʽ�/�>��>��>��o>M�,�>\��h��ڀ���9�]��=L�h?с����`�d܅>0R?g��:��F<bv�>��v�^�!�����'�>�u?�m�=��;>už&���{�x2��^�*?�/?H���>�,�oN�>P4%?���>u��>�~�?�7�>�<��]�<��?��U?֪F?|YA?��>Z'�<����"꺽�,���=m-�>)�^>uG9=r��=�v��V���!�|�="��=́�'ǰ�岅;n���8�<�	�<�y,>-Pڿ��J���پ�����o��F6��&������Y�	�(7��7��Y{����]�
�$)U�g�b�U����|h�)�?J��?�ҕ�-�������?�������I�>`wc�Fp���ݨ�RU��i���]ݾ����RY"�
�O���f�ne���'?`Ƒ���ǿ/����+ܾG ?�. ?{�y?��7�"��s8�Q� >�`�<�]��[c������ο6����^?˿�>Z ����C��>��>�X>�)q>+��➾��<��?�q-?���>0,r��ɿ̈́���I�<���?��@3�x?r^��P�������~P?�q1?.o?�w>���	���	,:a�{?\��?�Y�<:ue�[w	<�!�?/M�C����>P=>AЇ=��>=� .��>2�>�->CHҽ :L�H.���9���=:>w6�>�v�����Ҿ�>��u>�?�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��=����ÿԹ%��M �<v=��m<zq��^� ���ڽP�R�����m'S�|����=�x>bQ>Av>�	F>{�k>S?�d?>p�>��>���m�_�þm<�<��P��$� ~�9�/��r��dܾlѾ`�k���
��.ʾ��>��ap�q�=��L��O�7��-v��MI����>�^�>����%�Wbf��Ͼ�?M�}�>��1��n̾����n��u?��&?@�r���C�j�
�~��r�н�
*? �I�T������͜=��>��>�'>S��=��������@�"�7?�f?^&��u����Nl>����%1�<�?�K�>����ZV�>Ms.?�½ȕz�� >&��>�g>�v>��W>�C���U��I?��I?�� ��R��s��>�_��(I��v�)>�:�m0�<�ʼ|Á>��J+���s�=�t���ͻ<�|Z?�[�>^�!�Q��(qy��i<�6�=A�o?��>vכ>��`?�|9?6}=a^����K��s�u�=<uCM?)�_?Q(�=�>���4Ҿ�����D?��u?v�%>R���
��4��྄�?��O?\�?m�>L{�rN��E��8A.?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?s�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������z��=�ϕ�]�?i�?ã���c<6���l�UT�����<v�=�F�ǃ!�����7��ƾB�
�u���߻��A��>bT@H��=2�>c08�{1��FϿ	��*[оWq���?�z�>�Ƚn���"�j��9u��G���H�Vy��^�>)�=]Z�<�J�Ko��(��%����>��z>k�?C�,��L��2f�,��=@SL>7�>Ь��]��=�����u�?�Uо׭��Î�L���⬸>+��?Y�?ݹ�>�ݽ=m���7�
	�=N^�>9N?U�1?)1���;�/�&�j?�_��bU`��4�eHE��U>�"3?�B�>W�-�d�|=�>���>g>�#/�r�Ŀٶ�<���L��?���?�o���>n��?vs+?�i�8���[����*���+��<A?�2>���K�!�+0=�KҒ���
?]~0?{�i.�[�_?*�a�M�p���-���ƽ�ۡ>�0��e\�4N�����Xe����@y����?M^�?g�?ֵ�� #�g6%?�>c����8Ǿ��<���>�(�>*N>;H_���u>����:��h	>���?�~�?Qj?���������U>�}?�M�>��?c��=�y�>#�=6ް���+�0�">�+�=xb>�W�?��M?�!�>��=�9�0�.��%F�|GR�W���C�n	�>Y�a?�L?��`>�y��v�1�3� ���ͽ��0�NF뼰A�gF,��iݽi�4>6=> >��D�NSӾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>A�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?vQo���i�B>��?"������L��f?�
@u@a�^?*<H��|̈��Jƾ8��G�>�њ=��=����e=�p=^��=��X��I;�q�>إ�>��G>���=E#�=ט2>)�s���0��Zÿ\.���-��-(���S��'���:��3y	=� r��N���9n����=��=�;���{�����;T��=�R?�Q?+�r?'0�>f/�de>kN�<�&�F��=�+�>$�/?�@?, ?[��=�"���d�.�}�&F��i�����>�O;>���>_m�> _�>�d�<��Z>��>`z>��=���=�벺�Ϫ;�+U>�.�>gW�>��>M<>��>�˴��/���h��w�̽���?s�����J�#.��\8������k?�=r`.?�>����;пc�,2H?�����,��+�[>��0?�_W?z>�����T��@>�����j�1Y> ��vl�ߍ)��-Q>�f?�7f>��t>sc3��g8���P��l��9�{>a�5?3�����8��pu�wH��#ݾ�M>�Ҿ>nF�0&�͖�Y�~�o�i��t|=yT:?�h?��������}u��
���+R>*d[>�=N��=�M>�{`�,�ǽ,H���/=��=��^>L��>:í=}��>1�>��d��͖�M��>�]>���>�+Q?���>|6��ޔ�T��=�ܢ�X�����>�5�>(�8����>>{�?�ά><aҾ&=ۼ�=߼bR=8%2>���;3�^����Z=޺D�!�*=�@�<he�=B_����8��~?���!䈿���d���lD?O+? �=d�F<a�"�5 ���H��&�?o�@�l�?��	�ϢV�a�?�@�?�
��l��=H}�>`׫>�ξ��L��?��Ž1Ǣ��	�M)#�LS�?��?I�/�Pʋ� l�E7>�^%?߰ӾNg�>�{�VZ������u�m�#=��>@7H?NQ����O�A>��t
?#?!Z�K�����ȿ�{v����>��?~��?��m�8@���@�_��>S��?�iY?�ni>f۾hZ�b��>!�@?�
R?5�>�9�[�'���?޶?+��?�!I>*��?n�s?n�>�1x�vZ/�4��#���Kn=�?Z;�h�>�j>^����hF�bԓ��a��F�j������a>��$=-�>_\佾1���Y�=�ދ�:>��d�f�ݛ�>x)q>V�I>Q�>�� ?t[�>ख़>��=Cu��U݀������K?���? ��1n�ԉ�<>��=Ѱ^��%?6G4?8�[�c�Ͼ�֨>W�\?ؿ�?[?i�>���=��R濿|��\��<��K>�,�>K�>	���CK>�Ծw5D�ak�>�ϗ>�����>ھ�,���Σ�pA�>Te!?��>Ү=JM ?�"?Ow{>�U�>�hG��ג�#F���>1�>*:?�}?�<?�	��`�3�����A���Y���<>ly?��?$��>V��-6����<��T�it� ��?�c?,�ս/?Gƅ?�8?��=?�2z>����޾�=����>�?�}�M�7���.��H ?�w�>�f�>թ���Z�}��=fE���)��>��W?~?���`mK�T����=�D;�0����)������>>�[�=Xѕ��ۣ=>@[>*��=��d�j�I���=Ҿ�=�L>� �=�(�/o_�e:,?�H��ȃ�W�=��r�Z{D�t�>^=L>�����^?^j=��{����os��0�T���?��?@l�?�;����h��=?�?� ?^�>IQ��`�޾L��=_w��|x�js��>��>R�n���C������F����Ž�@�/��?F��>��D?u�>��=��?2y=	����N�'O{�#%��}���xľ`�V�8��㰺�vK> m�ur��䀾"?XD�Dr�>2Ǜ>�-�=ڙ�=,�
?vv>���>�yS>�F�<X�r�����߽�6�����q��?�?���Av�����N4�;$U?��?p�`?��<&։�q�1�+�>5T�?5��?h|1>��{�����w,?~��>K����?&?V���f>
m�ZՑ��B�����=�X>>]���D�w`L�-���M?�3.?C$��.K�7�>;���Ss=�?�8)?i�+���R�=p���V���P�M1�O�b����gC!�Jlp�����Q��e��<�)��M;=�D+?S�?���P��9٨�k�Ca;�\�h>���>P9�>h��>�<C>��*�1�ЌZ�̍$��v��v��>i1}?�B�>��H?Ɍ<? �Q?ӎH?p'�>l��>�����i�>���;m%�>�j�>9?�,?-?�C?�+?��Y>�� ��x��Wؾ��?�^?�D?D?�W ?p�mH���ؾ�v�K�,����T���=d�<��Խ��k��C=��T>�
?v4�0��x�b�>om@?���>�l�>�����h��=�=٢�>L(�>V:_>��˾�w[��4�K��>��?(���r^=��4> �=��<�'�</�>=)���o9=�ؚ=����q�<�|Y=w��=��[<���gv=�<P
>=mt�>��?���>%E�>{B��6� �f��Jf�=�Y>$ S>l>Gپ�}��v#����g�Wy>w�?�z�?�f=��=ʑ�=�|���S��z��z������<z�?/K#?�VT?���?�=?�h#?c�>�'�WL��#_�����ϭ?y�+?޷�>����ʾ����4�3�gM?��?�F`�:��b�(�oOþ��׽��>�1/��c~��꯿�2C����a�'������?Gݝ?��?�	�6��.������ѫ��B?��>���>�~�>S^)��g�8���)=>!�>��Q?`q�>z�I?�}?i�]?��!>Y�>�� �����3�c� >�=?�T�?�D�?��d?��>�m=>��9�}\�=�پ����ӽ(��Ǆ=���>���>�>"�>t��=N,��<m^��S��=�O>�l�>p�>���>3�j>��7=9"J?���>l>�����S���>r��a��sr?U��?)U)?N� =Ŝ���>����_��>�M�?�?O$&?�O�D|�=��
������:��\�>վ�>���>�
%=EP"=�>���>��>��4�/a�hA3���s��?�C?8\�=��Yd��a�8�t��B$=�8���$�?F�������>���>?�>��4��&��=���>���E���	�>K��>nM>��e>�0p=�o�<Z�2>���=�쵼/9�<%%M��(=��56=c��=䋏<�&��3=���=iҡ=�A�<i����z?�}F?y)?�;C?�u>�V>��6�繓>�����?��c>x�8��þy:4�6`��b�����ܾN�Ҿ�\��`��h�>�Ձ��F>�D=>��=j'��8�=q�_=v��=u�;��M=�}�=�A�=<ܾ=+k�=��>/>�6w?X�������4Q��Z罥�:?�8�>d{�=��ƾq@?�>>�2������yb��-?���?�T�?>�??ti��d�>M���㎽�q�=J����=2>r��=v�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>2`>2�]��0F�5�#�2���]�s������>���ͽ��<��>�+G>^n��Zξ�g>ˬ$>T��Y�A��7�����=]Y������7��<�HR>R|�=d�F=a׼(�>\�>��=�V�9ˏ���!>�QF=�!H� �b=C��>�U?>�b�>�?f�0?�ab?���>�p�:
Ѿ����>�X�=�:�>�=ZTE>���>2�2?��B? UF?C]�>�]�=���>�5�>�..��d�H�׾����=UI�?`�?��>���<;^O�;��:�l듽�Q?�w&?�H?� �>�>�4��\&� �.�l��;M�9J%)='s�ΧW��v��8����ὔ>�=4�>��>��>e�x>�K9>�O>w�>n�>/B�<��=�Ӎ��0�<~������=�;��
�< ļ~o���#�G+��������;���;1�`<�4�;ܛ�=���>=)>��>3,W=�ݦ� g1>�����L�7w�=�ࢾ��;���[���x�ۻ,����<J>fiB>r���z����>pDZ>MY?>@h�?�)~?�>Y? �jƾ���7^I���\���=�C>p�D�.�9���S��"I��-Ӿ��>%x>��>��r>�.���B���o=h�\k����>Bw������[����^�q�������
d�w�V=j3?.��B>&q{?׶H?&��?��>i��^fѾ�>ؓ�'�=�_���"�h���+�?$?��?���&?��<̾n��c�>�I��P�Ÿ��K�0�������ʉ�>3𪾣�о�3�'c������i{B�p:r�Vغ>ĳO?��?b2b��V���UO����H���6?5rg?��>�J?q6?	K��<g�X������=b�n?���?8�?�>d�>3d��>���>��?��?%+E?qC>��#�>�(R=�7>��	�%"6�9:�=I24>~�=���>8��>
� ?̀��
���྆̾�F	�����:R��> �>���>�׽�Tv�;R�<$��>��o>O�*>�b>���> E<=,뾋���~p?�����=���>ru�<�Ľ��?��m�=�S6=�!�(��� =�f=׺ ��Je���=�*�=ɡ�>�����?]�>�%����?���܇=ț�>�9#>S2�u��>� O>�}�=�]r>u�>B[<�=��^>����!>U6��(�!���R��a��i־�.3>n��LW�#'��
�0��L������j]h�Pq��c$�C�̼���?�	⽉�O��+�l�b��<?n��>�)?���9��B��=�.�>���>_�\����'��uS߾h�?���?'.c>�	�>ӿW?��?�1���2�WrZ�«u��'A�Ne�a�`��ڍ�3���H�
�������_?��x?drA?��<L=z>ٞ�?5�%�����=(�>"&/�$;�!K==\C�>q0����`�]�Ӿ��þ{��aF>Ǆo?�?�[?�bV����j�/>Ƕ6?�~,?�r?�Z,?��1?b-���?C�>8W?��?<2?�c ?�{?ʋY>Î�=�X ��1=����������Ƚ�{�u��A�h=jG�=Mo	�p�@�>K=t�)<����8��'��f6�>=-�u=D��=��=��>1�\?!�>+�>|�7?����7�����7-?��-=Ѣ����=*��zW��� >��j?�?(�W?4�e>3�?��!D�a>[�>��%>�W>�!�>��':E�-�=V	>9>�5�=��G�H߁�����
���ǵ<xB>A�>��>�F����A>yT����1��Ԙ>��	��̾n(���hL��g/�Sn%��^�>z5=?�?R��=N̾C�����s��*?��!?�5?_o?=�>����6��H��y�Z��>��<��3F������q.�;��=@�Q>"I��&����s>�K���%־M�n���O�In�֔n=nv���)=FK�T�ݾ����;�=rP>����������%���;FJ?�lN=,(��:�I��0¾n>�G�>���>��E����A������u�=:a�>�u<>hX��a����G�(��5)�>�SC?��e?���?�?��kz�� J��D)�܈�N�=�.?���>�?�>�*�=����0b�we���-����>�A�>�3?�$������G羁>���>�Է>�'==g�?lJ?��>%��?��.?@�>�$1>%��<v���\?�Æ?�6W<-��=�E��=��}V����>b�>�M���g�>�g?j�?�C??3/W?Ő�>|?�:�ס��F�*�y>P�>�{n��h���m?>��\?�s�>zX�?�a�?9ԉ>��5��	������3">��>OG?�� ?(u?���>F��>�ǡ�đ�=���>�c?.�?��o?
Z�=s�?�2>���>t��=���>���>�?8O?D�s?��J?���>g��<���+d���s�8nS�2Ɋ;�I<��z=0B�iWu�h���Z�<l��;�᷼�����&�{�D�v��ق�;�T�>T~?�u����>�����j��-�=��:=/� �c��
D��ݬ<�;?�W?�M�޾A<3�J>�?�Q�C�?ߦ=?�>�t�<g�����	Q���O�>i�'?�*x���Y�i�o�T3���bƻ�'|?/�G?��'�Ys¾f�b?��]?Kb�-�<�T�þa�b���|�O?>�
?�G�Xճ>Q�~?��q?���>��e�':n�,���/b���j�@ʶ=m�>�B�T�d� �>.�7?�L�>K�b>��=1t۾u�w�(v���&?�?��?���?�B*>p�n��(࿁���>���^?q��>\���$�"?X
�W)о�㋾V��g��]���2���z��ah��7n#�U���<?ؽԴ�=�?f�r?uq?�_?  �f�c��^����s,V�W��/�B/F��E�mC���n�G)��f���Ø�"?G=Í���޾�M�?�.�>�ɡ���>n�ھO9�k�ᾧ�>�ob��2��L���c�#X>���>�����4�����c?���>ѻ�>^M?2wI�#cF�z<1�|V�Ur�� ��<��>)�>&?�J�>�����~��?׾�c���T���u>��d?�I?sho?^C�Q�0�
���ƫ��w(�=��t�7>W�>���>�^E��8
��&���=�ѧo�/1������w	�Th�=�.?�1v>���>�#�?�?e��w����U�2����<',�>D�f?3�>�U�> E�m%�}��>��l?��>���>^Q���g!���{�!˽>O�>	�>��>j�o>��,�8/\��l��/~��Q�8��/�=ƌh?W�����`�g�>X�Q?�:m�F<њ�>P2x���!���H�'�7>+w?�[�=�m;>+�ž�.�͘{�B$��-6)?�?����)�q�~>f�!?���>���>��?ٝ�>�wþ����!?�_?�aJ?Z9@?U��>��#=Y����Ƚ�&�6+/=��>!|Y>ƶm=�0�=L�M�[����im?=P.�=Aeȼn���P^<�����T<���<�3>f���[�E�?��T@�l ׾u���
]_�qT���T�ݩӽ�+������Q��$�CȽ��n7���a��K-g�70@q_@_������+��uK��	�Ѿ�v�>�^��n�/ݰ�xց��P��7s���]s,�5l{�f�����}�z�$?�+���Cʿk������0
"?�v?�Zu?2 ��f�X2>�1>"��<���<;�/���<˿_)��\?�B�>����-���@�>(Ԏ>�
[>�A>`�m�p����5�9	�>�;4?��?��:�V�ʿFɿ��Ε;���?�Z@�8?:44�����դ>���>��%?A�$?�dоL89�m���p*?,�?ˑ�?��轿J��%�F=�)?�v�)����]���{὇�>�=�=�RQ��\>�i�>�^������B>�r
?�o�>]qý���<h���>��>����".�5Մ?+{\��f���/��T��U>��T?�*�>U:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=z6����z���&V�|��=[��>`�>,�ߋ���O��I��S��=�����ǿ���R^%���K=�s�<��s��������"�����qYi���ͽ?�j=�m>��E>v:�>su>,Kv>S�b?�q?���>͡#>_ڽ����k��A����i�#	�!|��"���2���o����"��N�#�?�r�ľ_OG�;��=��P�����c!'�|�_��F?��B)?��#>��Ͼ��K�H8�Kɾ�,��1s�H�ӽ�_޾�6��p��8�?|�F?�<���UQ��0��N�� ��+�V?ç	��������2i�=��n��<{W�>�q�=�k����.��K���)?��$?�#��xm��j'>J}�[�λ��-?�?/v�מ�>}?\ G�bDw���>-r>|g�>׉�>)~0>b���h�Ľc�?m�I?� ��×�(�>V;����T��pE=/~�=��V�SD��nK>�
=ןx�:�?;ThȽ��=�W?�7�>��)�S��7Ə�.��.<=2 y?i?��>x�j?}�B?��<�Y��g�S��L���p=x�W?ui?�k>����WϾT�����5?��d?�)N>��h����!�.�L�Ur?uZo?��?�-����|��̒����:�5?��v?�r^�cs�������V�*=�>�[�>���>t�9�l�>��>?G#��G�������Y4�Þ?��@m��?��;<�!�>��=�;?�\�>��O�-?ƾ�|��������q=�"�>����Zev����4R,�=�8?���?P��>Γ��ǩ��	>���lά?�x?.����:ǽtE񾷨���!���,>﹉>a8>e�;�Q�!'����㾀1�8�ʺ���>L@�n���?��{����ɿ(�g�{��D(����?�2�>���=���=��!�ʠ����P�?���3t�zE1>��u>���=��T�
Ό���8�@�8��m�>?�:9xA>}�������wȽ��>8�?,7�>�xC=:U羸�?[�!��Vֿi�����⾙/�?4}�?VqP?	��>?k�>B��B1���lU��N#?�x?|E?�->���H�;��j?�Y��iI`�_�4��0E��BU>E3?to�>��-��Z{=��>�~�>��>M/���ĿKԶ�_���
��?}~�?�d꾓��>�~�?H+?^�[8���I��{�*������(A?`2>`;��4�!��2=�]咾��
?C|0?|��E��!??��a�W ����I����r_�>A��<�D��G>�����=e�	(��H���q�?G7�?��?�� ��"��e?l/�>��ƾ�����=�r?�>�_�=H>�|>+���~i��'�>*+�?�]�?�e�>]���䧿m>)rx?[ζ>y3�?���=���>>��=F4���q�=�%>3��=�H�f�?SL?��>?�=��1��f/�3F�E�P�_c���B����>��a?BvK?"�^>,ж��1��!��>ʽ=�2����x#D�� �0R߽:�5>�BA>I�>6�I��sѾ �?#k�@�ؿ�h��{�'�,%4?S��>��?����t��H�$._?eg�>�6�B+��W#��;X��?�@�?��?C�׾�iͼH?>H��>M�>�uսD���Z��3�7>$�B?�2�C��i�o���>L�?{�@\ٮ?�i��>����i���g�%(�\o�_����?7Ϛ�t�
>�] ?ʀG� �w�x����wj���>���?w�?��>MX|?@��aAC�H�]=Zޟ><f|?4�/?��<�����9>w� ?M��늿.:�㟈?��@�/@*6P?������׿>��#����S��A��=���=k$/>Vn۽ ��=�|6=<"6�_�m�=1�>��f>�p>RYQ>�S=>~T+>�����R!�������qC�g������Y�H�Mps�����������X2��+���j�����P�i?$���U���=��U?�8R?uoo?f��>BRz�&z>�>��B��<�E#���=�_�>��1?�L?�c*?��=�Ϝ���d�A-��lէ�m���=�>�JH>�D�>���>�̭>�CZ��,J>w�=>V�>V��=Z�%=�=�&O>��>N��>��>�k;>ǎ>�Ĵ�`7��'�h� %w�˵˽T�?�i����J�7)���M������v��=zA.?�>���H7пe�[>H?��\�.�+�n/>��0?XW?��>���6�V�r�>P��S�j�4>^E �S�l���)�``Q>�~?@f>��u>�T3��d8��P�K`����{>+�5?�1��a^9�h�u��{H��lݾ��L>ӱ�>){9��<�g��~��i�`
y=�:?}[?�O��Jﰾ�Su�A��vXR>�[>��=/��=R2M>�?d�t�ƽ��G���1=[��=�y^>�p?Z�=vd>n��>�g`�j��H��>2-I�����V�<?�`Z?6)>�qe���Ѿuh����>1>�>>�	�I1�=z�[��<�=2_ ?`�>�d��X﮼4)��o�C�N:>��=]�y�d\o��=w>J�YI>E�D>
G>�ӷ4��J>>b?٥�)���"���~u>��J?�	�>5.>�&>�"�"��J�c����?e @��?�(���G���?�wq?bw���<f?�+�>0]�����Ż>RÉ�	{վv?6��䀽��?�|�?|�3�ά����Y�U�X>�w?�_��}g�>cx��Y�����6�u���#=���>k9H?�V����O�O>��v
?N?�X�稤��ȿY|v�J��>��?B��?U�m�@���@�A��>��?�eY?�ji>:a۾�UZ����>�@?�R?�>�7���'�D�?�ݶ?J��?"�H>l��?^�s?�7�>��u��o/�\��&���Y�=w��;�:�>��>z��%\F������S���bj�Ih���a>~#=��>�W��?���ص=~(���է�A�i��>�
q>E�H>KH�>�� ?4�>D��>�X=A����
���m��{�K?���?#���2n��L�<��=8�^��&?�I4? n[���Ͼyը>غ\?l?�[?�c�>8��J>��1迿>~�����<��K>4�>xH�>�%���FK>��Ծ�4D�mp�>�ϗ><����?ھ-��&U��`B�>�e!?���>gҮ=m� ?Ϝ#?�j>�.�>�_E�9��V�E���>��>�H?��~?� ?ι�W3�6���⡿��[��+N>��x?�P?�ɕ>����;����NF�/I���k��?Fqg?�I�<?�.�?�??j�A?=f>���#ؾŎ����>�-!?���A�v�"��<��?Y�?���>'f��"�ڽ��8��ի����?�U]?�"?C"��]��������<J�8�:ޢ�;QO���>ǒ>�� �=e\>���={�r��B1�w*W<���=t[�>���=<�>��臽t&,?��=��̓�R#�=�xr�KqD�_9>RrL>N�����^?�L=��{����x���|U����?���?Ze�?Ct��\�h�:=?-#�?�!?�>�v�޾���"w��ox�'h���>i��>k o�4�侾���,����,��F~ƽ:�Q�|?��>�U?M��>��'�7�>�5�����A�ǾE��9~U��C$��\5�sW	��kᾞ�n��d�B�=6߾X�����>�)��ݞ>%&?n >�}}>L�>�Ƽ;�r�>�oD=c)O>^�`>ai0>�8q>�63>���=ehɽS;?Ѐ�R.*�v@��n�ν�W?��'?);C?�E��s��l� ���?��?� �?�'i=Ao�2,>� ,"?ә�>�I�Sk�>T�I=�H9=�4H�z������L�=�^�=3��>kl½�S�^rK�����S?y3�>�EN��=
� �>����Go= >�?d�(?� *��Q�ۧo�p�W�	
S���>h��f����$��p��ꏿ
^��,-��|�(��*=[�*?��?���l������k��.?��-f>Z�>�'�>-�>N�I>��	���1��^��B'�����.��>�c{?dG�>H�I?��;?bjP?�!L?g$�>!�>l%���6�>8��;\��>���>CM9?��-?F0?�e?�Q+?�,c>���5��דؾ�?�c?�?�?.�?����N½�O���h���z�d�9�=�<��ֽH�r�/U=�*T>E'?O_侇�W��<�o?uqB?G.�>�DC?x�w>!%�uk�^����:~>��4?�p>�4v�P��� ?�\�?�p��V�=�>�):��+����r=u����g�=�E�+N0�y,�<WX�=!`!>a�j�\1����<���<�SG;D,>��l�>Xb0?�Y�>�n�>;�"��t�>���,w=�k�>c�>0�>0�ݾ�苿���O�l���]>x��?ó?Y�/<���=�>��m�<�ľ�F������$�=F�>6�?�O?"�?��F?�c?Ԩ�=���ߒ�������? ,?���>���%�ʾ2�T�3���?�[?�7a�����=)��¾��Խ}�>U/�-~�����D�P�������~����?|��?�,A���6��k�!���
c��#�C?��>�Y�>��>��)�&�g���;;>ҁ�>;R?״�>�V?�t?�[n?�c<>��C�ɪ��k���ɛ�S�=��;?��?V�?j{?�f�>lI�=4o8�}�ƾ�����s׻�������=��q>�'�>�>�%�>���=�$��Φ���u�,��<W�>~��>��>��>|:�>l�s=.W(?d}?̪���')�����WS��7��w9|?�[�?�"]?�l6�qK�io�v��_��>:�?m��?�j�>�ɏ�8�U�A�=��	�,~���A?���>>��>h�=�1�>�w=���>���>�K�g��©p�w/%�vn'?��G?+�=F	ƿNp�̝o��}�����;�����:d�؉��6�Z�9�=����91�o���b]�S���Qb��]w���r��_/}�xo�>܇=�X�=���=�ͥ<�Ӽp�<��M=f��<�=�d��Cx<��7��ϻJ���>����5<�uT=�|e���˾wq}?ɛI?ч*?��B?~y>�>R�A�v��>����)?2�V>��T��8����;��Ԧ��h����ؾB׾�Ad�㬠�3	>�I�J>D|1>��=�K�<���=%l=��=9%��(�=��=�:�=Ҫ=01�=g>1�>U�W?'�~�>T����k��B��3?���>C�?=�l��fk/?�;>3�dB��/;�x}�?���?� �?���>$�����>����w����<���=3�O>�{+>M�2����>��W>3�?�����/6;�!�?�Q@	�/?(ȋ�Yqֿ���>W_7>��>�qR�^?1��<]���a���Z��w!?);� �̾I�>�W�=Ţ޾��žF&/=�5>�b=pr��[����=��{�kg==a�l=�׉>hmC>5�=ꌯ��L�=[�H=)��=0�M>�ј�V5��(��2=Sq�=g�b>�K'>�I�>s?��'?�Uf?�o�>����AվO󵾫��>ߢ=?=�>�l=	�(>�&�>�<?M76?�>?�B�>���=�ΰ>q_�>��+��k���p1���=&�?\��?"��>׏����u�B$�5q6�*�t��?e ,?L?���>�I���߿"��ɬI�]��V�=���<[�{������|�BF�A�F��=y�> ��>�0�>���>w�p>��~>��>���=q�d�>S����༜��=B�=i"�=������3��L�=�?�;��2-�Yj���2�<�a>=�a�=J�>Ec>lj�>s�&�U͘��`ļj{�R�f�>n��hN��,�?�w<{��Q�m��<�%>g�{�zvƽ����d�0?!�&>Ӧ!����?�r?�r�={�nϹ�������D>��3;F���l>�������{�������ճ�h��>H
�>��>��P>i�8��Z8����;Þ�
�G�	?{��8Y�=l���s�a���E���y�Z�z��*6?�����>H>��_?{6?��?���>���Y̾�>a��6�{��b��x�!��<�p?uF?�i�>�þ�D��O��q��7U4>gl����o��g���gF��e��Y�_�-�=>|{A�o�Ͼ#`.���x�Y��WG�����;�> �G?�z�?P�׾,Ey�����;����!����=D2?s?`t�>�V
?;���ث���"k��x�=>��?R�?��?�u�=z��=�������>}�	?���?�P�?�ms?�7����>�;Y�>WY��v�=��>�i�=5��=8	?��	?�s?˽���������0�]�o�=��=���>��>�p>�=(�]=�`�=��W>u�>���>P)c>^�>��>�½�Ȃ���G?�َ=�Y�=�P�>9F>A,���  ����=	T������6ߐ��G��� ;$�E>��=p�=�J�<[��>O������?G�=^���8�?m��[�=�Z >K'M=O�!���K>m~p>	�-><ǘ>' �>N�?>>6�>�(�<�8��y >X����M��Ex��2K����E(m>nӌ��㕾�E���8�V�o�þ��.k�fj���<�!����ĉ?m\��M�M�d��@�P��>��X>�?���޽k��>+n�>g6N>O��፿O׀�Y�;�w�?���?�&>>�y�>�Jd?��?��K�k1x��^]�$|g��8�zY�G�Z�����IF��J�9LA��?c?*�q?�~??�ۡ<Y�z>�,m?Z?�{���2o>�&��u>��P�=6ݘ>�Ⱦ+�j��1ʾإ�"I�BbC>��g?:(|?O	?A�{��@�V�>�,7?Q�0?�)t?�M2?ġ;?r���$?��2>(�?k�?��2?��/?i}
?�G">���=��:ƀ]=�[��y�����ӽ�)ýE��J�F=�m�=v�<�r_;P��<k�<n�ۼBSļ�fֹ,P����<�$8=�f�=�o�=�e>�?��>����b?���~!>�|%>�;�X?WL�>-�	��ؾ5�$�/�<������J>?<4�?|O?�;):S���������>z��>(�+>K���{�=����g=���L=�b�=ͩj>?�>i�ɽ�i�����þ{">�4;=��>+��>�J�P�G>����0=��Xg>��E�W\���FT��N�:o3��z�m�>$RQ?ږ?i�=P=�ؠ�Y%m�5&?8"B?��J?��{?�聼"����7�V[D�N�轩�>b(<�#��d��񾜿�W*��B�<��{>`���vΡ�v�g>����v���t��B��l��*�?=>u���=-�&�����I�I���=�@>����Iz��?���9���;T?�>�=uw���A}�?$��>�Ԥ>�>�_;=T5 ��N��=�����=��>/މ>�
T�"��H�L�́�M�~>��J?��b?�K�?{���x�q�5-O�����s��9�?D?t�>��?34`>Z�=c���z��[j�x=H����>+4�>��!�[�/�ۃ���g��,`.��r�>�}?�|�=*o?]�R?Da?�]?��1?׷?�֛>l<���ž��>��}?d�>am>�=��UDi���]���E?�a?�K��̏�>�-?� %?�&9?W��?,?�U>&����E�q��>�O�=~Xp���#�W>��6?]K5>��u?h��?�C>�!�Rþ����俽�X �"�?_-?9y ?P�?��>�ܡ��4=�T�>��b?+�?.�o?��=��?�J2>���>���=�Y�>�#�>��?�>O?q�s?�K?�}�>�Q�<*���|����r���N�r��;�H<��x=9���is�T��t�<n�;3���S;z��f��~�G�ȗ���t�;��>έ�>`q��9��=q���E��	��>�Yf>y�R��Z�=�v =��>�>��>A��<��0�= 	�>���>B�:�S�j? ��=��>���<�ձ�"+�"6>���>-��?�r?�掿Xض��酿�E�=�V?}�?�"�w�T�U�b?��]?�d�I=���þ��b�ٌ�?�O?��
?j�G���>��~?��q?��>�e��9n�:���Db���j�yѶ=$q�>^Y�{�d��>�>�7?*J�>
�b>�*�=�u۾��w��o���?_�?,�?���?�-*>��n�K4�G��q��u7p?Z��>����p$?�6[�T�ྉ����y��=�žƘ��x�ɾa捾j3���-��Hl������<�l?��u?��c?Wwe?O	��X��bc�L��U����K	��A��A���M����+�����ٱ��<=�Y����C���?�%?�:�/��>�D��8:޾mDž�NL>cC���v���I�<|=X�hv�=�7�=��K���4��b����"?^��>ث�>��4?T�L�/�':�KiK��n��R�=�c�>@�>Q��>����Qh��(,�]־�<���N��-�>�q?�<c?᠂?I�S�a O�Ap��s�8���>(C���>���>_l�>�>�< >�T��GI�������1���z�P� �o��=m�a?1)1>�B>��?;�>Խ8��Ҕ��ѽre���5;��>�C�?�Y�>���>��i�J5&�<��>1m?���>2��>�狾��!��{���Ž��>�ծ>a ?g�l>G.��`[�G���Q���8��)�=:h?&[��x|_��W�>aQ?��:��:<���>�w��z!����%�s�>J�?��=&�:>�ž�es{�W��Ŷ(?�,?�萾�p)��>`� ?���>y�>N�?뛛>�H¾8ho:?k|^?�EJ?�A?l�>��=�����ƽ��'��G-=>�>�Y> �o=�=|M�4Y�M��MD=�t�=��ļ@��Og�;��ż��T<��<��3>�׿6�J���ݾSO-�ݮξ�����L*�,ܽ���F��n�龟���K�p��7
�S�g���
���M�;$��;�u�r��?�?� ��T��%���i��٫��Ȉ>�����@���ԋ<S��ݦ�(;t_��=���w��^a�.?"-,�$󽿗�����V�!�>[�,?ζ?쾶��=�z����>hD�=�f�<]FѾ�U����������vI?��>=Ҿc���?��>q�V>D,3>��d�����;�2?�C?��>����3ٿȿ�a�=~� @Ȫ@��A?3�)��	��YR=i�>��?��K>�C1�|3��.����>zr�?�V�?�V=
wW�F��3�c?�<LC�y*��.�=D�=���<�a�/I>:��>\���:��vϽ��>>#z�>PH1����ÌZ�gD�<�d>�uϽY��Ԅ?�s\���e�^�/�#J���m>��T?��>6١=(�,?�>H�p�Ͽ �\�v�`?�+�?;��?��(?������>t�ܾy�M?�e6?��>#{&�U�t����=�lݼ����~㾡V����=���>z�>��+�,��*�O������=5��lǿ��{9����=��]9����Rӽ��ƽ�qټQ���	}��=��υ=��>�b]>��>�8?>�(I>��`?mn?�٧>[�=��'�����qx��y4����~��d�E��~�yژ�Z�����7���K���ܿ�܄;��ˎ=oT��&���E)��mY�pu)�m�?���=�赾\C^�`�_=9���ی���9��Ja��¾�/;���i�Q�?��K?�`����j��i#�\a��؟�Z�P?�̽Ŗ��վ��=u=|��=�̼>�==0�[lG��K�&s0?kZ?͊���[��d**>�Ӽ=��+?2�?��\<�2�>OD%?�*�66�E[>Đ3>֣>#��>�F	>��B۽b�?��T?�������ې>U]��!�z��a=O">�;5����c�[>#��<��{�V�!L��诼<�=?��^>��G�׆���3�ҙ�U}t>�d?� �>�k�>*��?�B?ֿ=ʾ�T�AK���=`?ӂG?���>�F���|��E�.u?}�?0��=g����ǭL���)�Y�?Pޅ?7?)<�=ݣX��앿��o�X?({n?>
V�U0��&_ʾWD㼽�>A�>��>��5��>�A�>��ƾʼ����ɿ�f9�z�?�@��?a�9�kR�=գ#���?�P�>� N>M��� �����2��=0��>�f�/�O���ؾ�(��.1? i?ϱ�>�3��QNԾ���=\����0�?I܇?5ģ�>�=&���L}�����v>�b{�=<�=��c��D��W2������U�^0��/P�����>�@�(�Z��>a:w�W�ۿ��ο�뉿����s����Y?�kK>߹����ɾ�2x�jr�E�N�lT;���I���>>�Õ�������{�q;�y��� �>��6&�>)xT�6���w��`v4<��>s��>ī�>+R��� ��ř?5���3ο袞������X?Z�?`i�?�w?A�<<��w��{����)G?�s?!Z?*�%�R�]��7�+j?L���fb^���2�2:F��Or>��6?B �>��-��{%=g">Y��>o>'<*���¿�Ѵ�����!��?��?��� ?Pl�?��%?���扚�tg��%��#<�!F?�BL>p$ľ��#�D :������?3[1?�� �]�_?+�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?ֵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>_H_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�"�>��?b��=�a�>�c�=$��-��d#>�.�=�>���?t�M?oK�>}g�=��8�V/�\F�)HR�/#���C�,�>(�a?m�L?aEb>G��Q2��!��zͽ�\1��G��T@���,�N�߽@&5>��=>>y�D�jӾ�/ ?���ο�x��b����>?*$�>��>��L졾�=%��?�^�=�<�����)��M�X�M��?'u�?�#?�,�=Ȱ���>�n?"��>�^V�,���MҾ|�g<��L?6Nx�Ai��q�x�qt:>2�?�?@�K�?`\���>�ڸ��怿ϭe�c4��ӧ��%>��L?����<��>z?L�u�:~�1�����]���>�2�?z:�?�#�>r�O?��`���K�:9�=~n�>~bE?�i�>ȇ*�+7��o>s��>�z9�A���!�ʈ+?��@��@�(X?!ݢ���忕������9�����=�Y=7$>����v�J�ߓL=��=��ټD�>3Ú>d�Y>�� >K>�gO>�R�=�:��b��e���������G��3۾5������:��ޚ��Ĥ������D��7�gA�;�B5��4�����4�[=g�V?	�k?�?M�>�+Z�D�>=.�(���w�A^��>��>�[7?�j?Q�g?{V=m����v��w������'	f����>_R>b��>s�>>�>��=�U>ָU>j�6>�<�=Q�=��мm#�=d�z>+��>p��>��>6"(>g�%>���������{�(n�^�Ƽ���?U����5�G�����u�l4���M�=!m2?�>g���7�ѿ�n��>H?���#5��U ���-���(?�L?�Ii>v�g��-�`Y�=� ߽��e��*>��^���.�^av>�@&?�f>�u>s�3�p8���P��y���z|>�36?ⶾ�69�W�u�U�H��Yݾ�QM>�ʾ>�C��k�,���>��ai���{=�s:?Ǆ?򈳽�ܰ�2�u��2���kR>8\>�=�o�=�PM>�c�_�ƽ�+H��.=��=~�^>g�>��h>됎<-�>����7`���u�>�ˊ>�`*>#X?�Z=?��ŽF��I���>[��P>(i�>�6�>�t>T�K��8�=���>r�O>��=�ɽ<{ؽ�(��G>@�����E��f��Ca�==ͽ�p�=��=2d� �>��
>=�~?���䈿�뾂d���lD?Y+? �=W�F<��"�= ��@H��=�?d�@�l�?��	��V��?�@�?���s��=�|�>�֫>)ξ��L�ܱ?{�Ž8Ǣ���	��)#�SS�?r�?s�/�Gʋ�l��6>_%?�Ӿl��>�52���މ��S���^=	6�>�G?������@5\���?�q�>4��8��zȿxo��4�>0��?eœ?s�r�IᖿL�$�� ?�*�?Y@J?&{0>�v���y��!�>��A?�1?cVX>�!�F�%�_j?��?T��?Bk�=�}�?�'�?M�>� v<ǘ�e\ǿQ�j�@?=ꌾ�̪>����Łݾjy־yy�� c�rg��(�ˠc>���<y��>�}R��վ:�R=�'��L�r�].�1r�>7v�>ۆ|>v��>�5?v�?�?>R�Y���]���Ӿ����+�K?u��?���92n�_T�<|��=x�^�w'?sJ4?n[���Ͼ�ը>�\?L?�[?5d�>���*>��迿�}�����<G�K>[3�>+H�>�#��zEK>x�Ծ�3D��p�>�ϗ>���#?ھE-���x���A�>xe!?C��>�Ү=� ?�#?<�j>�$�>�]E��;��j�E���> ��>�L?��~?��?�ٹ�UX3����\䡿1�[��DN>��x?�Q?�Ε>_���V���W�C��lI��������?rg?�`录?[.�?3�??�A?B(f>:���ؾ��� ��>�!?W�m�A�:L&����?�O?���>�+����ս$(ּ���r��� ?&$\?<&?)���(a��¾<8�<G�"���T�Yb�;�D�N�>M�>���w��=>�ʰ=�Jm�,B6�+(g<�l�=}�>{��=�-7��n���X/?H82�TDԽ0��<yd\�1���b�>�?:>R���?O��d䅿�vJ���@�=,��?���?��?>�M��w�twV?�ܒ?@�?�>�#������喾"i���R��派�9�>3�p>��>h�ʾ����U�������ý�U�E??~�>�=?OA?���>dv�>=E׾NJ��߾ b�x�m�EE�(�F��9�D��=o���j��s1�w%׾7^��7S�>T�!�R4u>��>�P^>���>��>���=1v�>�q�=-B�>W;�>ڸs>t�>�=BH�=Yɦ�:-Q?�JϾLN���վ�?Ⱦ�_?*�s?��>V���冿�����/?E̊?���?��	>E\�L����?��?������?�3�=����[�ӽ~	�ܶ���2<�<���>|n,=�=4�(�X�3g��>�>���>$��=���k|{�O��}+�=dL�?��7?�&���E��"|� bs��8H�*_I��H�n�ɾ�9�~:n��\���r��~x�z$�܎��d%?႔?7�X��w��� f��`�U�>=?��,>v��>U q=pZ��1o-��$S���Q���E�>�`�?^]�>�uI?o<?{tP?�UL?p�>%j�>����6��>���;��>�>�9?��-?�F0?�v?#`+?T�b>ML������ؾ$�?�O?�?o?h?׶������`'���f��y������c�=�ƹ<�ؽK�s��pT=�	T>�%8?Ln���:��}��HT?��Y?d��>�N`=mo�Q|�����U>8sk?���>+���Bi��"$���>c:�?@{�\B@=?�>�@*>X���y�=�ߨ>}�������Z��*���>ع>�Op>��P<��%;�o�?r����=�>��?N��>$��>rՅ�/� �w��K�=z�X>�S>�>�Zپdo�����zh���x>�l�?���?�9g=�}�=
��=����j��$��񧽾7@�<�f?�G#?�T?P�?�~=?h^#?��>����8��f�����u�?k!,?
��>����ʾ��Ɖ3��?s[?s<a����;)���¾��Խ��>�[/�`/~����CD�녻���4��!��??�A�H�6��x�ʿ���[��m�C?"�>/Y�>i�>^�)���g��%��1;>N��>�R?4�>|�T?���?�Z�?�1>_L��壿B ��������=��???Ƅ?&ه?��?'_4?%��=����/��J�.�5�{���ֽ��?�u�>{�i>b�D>Z��>ϛ�>G�<�*м���"���=��9>��>���>B��>sr>����M	9?)V�>��Ͼ�Z����A¾��<A�u?��? 	L?EԵ;��7�m�Q�@
��>Lj�?d	�?�1?���46>����氾"q��p�>���>w�>ꀸ�m�=�� >��=>ܫ�>&p3���6�=/�}#->u-?WD6?�� ��&ƿ?�q���p�䗾|e�</���[<d��e��
?[���=�>��20��֩��+[����J���ۧ���̏{�~��>�R�=H��=?6�=.	�<7�ʼEw�<�NI=���<x=\�o�.Xz<&V8�����I������)\<�H=$��ɾ�|?"kI?E�+?C?�l>��>�頼�O�>���pg?<lX>�Z(����5�1�w����ޑ�D�ؾ"�׾��`�������>��]���>u�3>���=cĂ<���=��= �=s�����'=�E�=٨=�8�=u~�=��>O4>6�y?�A}��ц���2�)��<�:?��>o�i������v6?���<W-���x����9���k?��@e[�?��?[���z�>�%u���!>*�����=�j�	>^�|>���0]�>^��>����ݎ�h�`�,۹?S��?d^9?3���(���e�f>b�B>��=|�T���1���P�bX��[�S�!?� 9�l�žĔ�>��=����̾��<05>��=g�～tX�^�=[h���=�Cn=���>�&D>PƲ=������=tg=vg�=LH>���;��0"���7=.r�=��]>{3)>̔�>K�?1�2?��h?�^�>�\��R�ؾZ���^ؙ>�6�=���>=$�=77Q>�ƿ>F�??�^C?[G?��>��&=
��>B��>�1�!�n�OپY���ƈ;�?ㄈ?�_�>��;�IF����E>�B;��<a?��0?�w
?��>aC��������%�F�����޼�!�<ŋ��"��6B��h�W��O-9=���>�@�>@ū>��3>�u�=�'>�R�>d�>��=����#�=v��<�Wb��>�=R��=c��<]ý���<@ӿ�l�:=��2=<��=P�U=��%���/=ۿ�=��>�_{>���>2"<>�P��<h>�#׾�b��p>vB��"�7���u�v9���L��?�<Wh�>,��<V�g�5��\?-wY=��>���?�5m?W�>Լ�=8��1���@E��Mz�ĝ>z�+=�J���N���p���P�k����>�a�>qC�>} l>�,�c�?��\{=���%5����>J����T ������p��4���ݟ���h�T$繗hD?�>�����=�q}?=�I?��?@3�>@ܚ�˓׾t�0>@��^'=Fq��r�����Z�?��&?+h�>�˧D��A̾ľ��ҷ>�BI��O��ŕ��0�������r��>bા��о'3��d�������B��*r����>\�O?��?�-b�Y���PO�C��ZY��l?{g?��>rN?C?޵��{����j�=*�n?ĸ�?�:�?(�
>ν=���"�>�%	?T��?��?�{s?�x?��W�>���;-� >�����Z�=��>+�=/!�=�l?]�
?v�
?=���t�	������6:^����<�ơ=���>�|�>��r>=��=>Zg=7\�=�6\>4ݞ>Fӏ>��d>K�>
P�>ʧ̾����B?(�>e��>?'?_��>��>��@�4>������j���G�ґf=ʼ3>�,�=����dT����>��ʿ�D�?�G=�"��8�>F4����=pu�>��;>d�R��d?o	��j�>�>�^>�h�=���>�%~>��Ҿ��>�S"�=2D�)R��rо�|>�~��Z
%���	�&>�98H�f��k��H�i���,�=���<�#�?�����gk���(�ۮ�V?R�><6?����|���PU>t_�>�7�>ڑ�������qUιf�?��?�b>X
�>�$X?��?��1�4�*9[�w<v�� @�Y�e��_�
��k� ���}Ľ�&_?��w?3X@?��x<��z>���?/�%�B���a�>�.�]�<�^�N=[y�>�U���*b���Ӿ�¾
�IPF>�n?R��?s�?MYL��<K��H-><C9?-0?q?&]'?��+?�Ǒ��C4??/>�7?Ay
?�)9?�[.?�?��0>�>�=?
��Q(=�L��_�������ֽ:G���C=KA=�E��� �<�AH=�K<��á���v���3��;�9C=W�=�=3��>wL[?�y�>�ߋ>h6?Y�1��=�`\����;?� /=�Oy�O�������qR�r�>ңh?7�?$S?��S>��9���I�s><A>� >�^]>�#�>���P0���=�6>@F>匱=c���l���
�'��h�<X >�M�>AB}>5���g(>i�����x�e>^�Q�ِ���hO��hG�ڟ1�=M{��+�>��K?�|?��=��������g�&�)?�N;?}#N?SV�?~�=�|ھ��:�n�L�d#!���>�C�<�U[���w��%�;�_����'m>[ٟ�Ue��ņg>D�	� ��HUs�U\M��R�ܡp=�
��:=t_�4վB@o���=�L>[�� ��w������J?ە�=򋨾̕I��X��K��=�>�]�> c��s��GD>�^���*�\=;��>�>(����PF�.D �#>�&W?fS�?qB�?8��5����J����/��A	½y�?D"�>!N?�"�>o�>�Ӷ�?�Vd{�!�d��`�>3��>��g}M��M���ؾ��1��?�={L)?�I`>Բ?�y|?��6?�2b?�e?�+?x��>Xa�<s��� ?P��?S�>u�4�])��M�U�Y����>b��?zw��+�>i4?8~L?��k?�Z?�>�!*>hm��Xe�'qn>b�>>3}Z�w��α�=u#I?��?�?�?�=]C�,� h�����|�>�f?Bd!?�E^?�z�>�W	?iоW&����>��f?}�x?�aY?܍g=��>h�>Ew�>fe>��:>��>���>ÂZ?��?m�\?<��>6�<'o��Y ����aƽ)v�=N�?=cB̺�����������o�藮<~��<"�=��G�CDƽ�K:�7�V=[E�>Mc�>^B�����=!��>���֥><��>E�͔��7�=�U)>{g�=��>
rD>�a�I�=o��>�q�>m5���-?�6�>�Q-?*9�=��y��������>,� ?h�?� �>*.l�g���N�l��=��?��?�v~��`;���a?��^?�?��=��$¾�`��Z�ϻP?1�?�K�C��>��~?�7r?��><�i��Vn����/�b�_h�u��=d��>� ��=a�k��>�t6?٤�>}O^>[�=z�ݾ�tw��p��f�?B��?�I�?~z�?�*.>n��u࿹^����9(_?�k�>�J��f#?0;��Lо�*��Ğ��G�߾ʞ��Ϲ��dҔ��E����#��̃��|ݽ���=f?��r?<q?�_?m�z�c���^��e�jV�1�A��w�D���D�KC�:go�s���<��=����Q=Ņ�wu<��|�?��/?��|�>����l����ž��>3e�H���jѼRs���>ϼ�=��_��Nk�4_���a#?3�>H0�>�-?��]��5�;�e�/�������O=��>�T�>�V�>&"?��O��nL���}�L����9C����=�~?�LU?1�w?E��=ۍ4��O��p�����>Ku&��;>�	�>�R�>qU=���)i+��G�1H���A��c��ß����=ʬ�?Y�|>�m=�k�?J�>5�6��󛾜���B�,�s��Ю�>�֋?0�>kN�>�ؽ�LI����>�u?֎�>��>|�;X�����`Լ^��>��>�(
?���>�����L�{���፿�E?��a=#=b?� ���h���O>�~[?c ���|<���>�����&������-���>$�?�p�=��1>X������
�w��ٱ�H�#?k?a����(��p>8_?#}�>T�>S6�?�/�>�E��Zq�<�J?Z9d?��L?��;?,��>,@[=<��fdнl)��M=��~>�M>b��=�l	>��� _�	=�2�7=��=f�>��#н�<ο¼yp|<i�Y=Y�G>lIпxT7�FK�������"�R�򾺊����3 8��@�{�ž幁��䘼˼��\?�C?��V\�f��k�����?S��?��Z�)ϖ�y՛�\���mL�{�>��#��:t�>k��w<�E|��Q��oq�:�K�/��Y�1�W�D�'?巑�$�ǿZ����Dܾl ?A ?,�y?4��"��8��� >?[�<pN���뾅���G�οǧ����^?���>�
��R�����>���>�X>TMq>k��瞾&g�<��?b�-?���>�r�Жɿ]���Ǥ<���?�@��E?B�7�,[�|'A;n�>�{6?��>��I����zjO���M> Q�?�O?P�Y��Y����==��?���>ޅ)��[���h>�!�=��X�7
��ǙT>�3�>���;t����c<0�>"�>����t��G���>>����<��-��JȺ��w?�D;��F*�� ��J�� k=�J?�+�=g�k>+�Y?��g����-�^�l?F@|��?
�?`$ѾX�Y>@W���I?gTQ?5/q>�d=��	e��\=�>>�_>,���(�B?�=6�D>�p�>4u�����v��e�;O>�����ƿ� �����F�;8(�<�쥼�#+�5���z�"�-��w�l��f}�<K=8�>A\K>#�s>��4>�#M>F�_?�qo?,`�>���=W"�C���ľۣ:=_�c��I]�C;o���ƽ������gپ���b������Vоc=�0	�=�O��J����&��He�|�B���-?�9(>`^ξ��N�OM�;	P�������ߟ�iD����ʾ��2���l��'�?`�B?�����nQ��`�Q�u��Sɽ#W?p�������A�=���gNL=���>�vz=���2���N��L0?O?�ٿ�ۀ���}(>qt���=,?� ?��m<钬>�%?+�+�E�sZ>ˀ3>$��>��>�>@����ڽ=?�T?�H�񮝾ȁ>?뽾��y��^=�D>v�7����\>���<8���j�Uِ�h��<a�M?-n�=4b5��}� uܾ�<� �>Y�T?�kg>(��>��f?\.?�8:��⻾6�7�0m�H��<�N?��^?Qc�>vun�����e�)�b?��?7�> Z�{׾��4��{W�;U?�a�?��8?lM>��f�	����B���|?�t?�����l��1�J�r�>��?R��>�'c>�<��n�>�b>J��>�i��\��&L���?���?���?�
����<AZ� v�>��?�)>�����A��踄��H�=3��>)�ľ{1	�d�����<���>|/>?�O�>�r����C޲=cb��鲵?ۆ?�|���7=dH���j�����\���>��Ǽ�>� �ᾗ�����N'	��S¾�u�1�>�@�>*�o��>� g�� ޿�п.u��Ǿꮾ��?
��>���Ǻ�0������ŏK�Ί4��$3��R�>��>e���?����%|��;�f`����>���Eԉ>6�O��ȶ�l)��oK.<��>��>?��>U۬�/������?t���O�Ϳ�f���g���X?>�?�,�?�?P<I�w�4!{������F?�Ts?ƊY?�%�'�[�>�1�U�j?g���6�_�U�4��D�R�W>%3?/,�>��.��l=�>��>H�>).�ĿEz������d�?:1�?�����>��?+?�;��������')��<t���@?�O5>����8"�K�=�i�����
?T�0?������,�_?�a���p���-��ƽ�ڡ> �0��o\�>F��g��/Ye�Y��mFy���?�^�?�?H��) #��3%?J�>6����3ǾB��<�{�>s#�>4N>e_�)�u>y�P�:�ec	>?��?9|�?k?ܒ�������J>k�}? �>Ln�?L��=fW�>h��=����穴��(>�=>K:P�X?A�M?\3�>r��=C<�rw/�e�F�a�R���R'C��>�_?7N?p�b>�3��	�'�/�!��%ʽ�K7��ݵ?��]���׽�%7> �>>3<>�E��׾ V?���\ֿ�n��'Ⓘlh$?`��>���>$����v�	i=m�J?<��>�I��v������T�V��?�V�?/�?Q��!������=5�>��>��E����X�W�>H�K?���><����}��,�>�.�?#�@H÷?�e�hI?SS��t܍�����cE�D��\[8>�f	?�9��(i�>��?No@�Zl�p��愄�:��>�ۧ?ƞ�?G7�>+jw?���m�0��)>$*0?[?v?���>`����0��>�8�><�R��w��Ds)�Q�h?�@��@n?�4�����Y3����;}*��s=Yޠ=�(#>~����> �����=�zŽ,&=}j�>�:�>uIv>��$>d�>�y/>�����z��2���[����9�%������qy��(�V�Y�f����n��W�
�XR2<�E���hd�,-�u	�������_?!�w?�Q�?�?����C=D�Ծ���<_΋���==;>��.?	m?DZ8?��W�fFʾ��}�u��4���y�e����>h�1>^q�>%?�>C�>Iw�=���=��>��>�o�=J+i>���=��>��1>��>���>��^>*<>ٜ>!˴��/����h��6w�z̽���?�}��e�J�1��&;��͝��LI�=Z.?�l>j��=п��`3H?9���n.�F�+�	�>��0?q]W?Λ>z��0U��=>�����j��i>Aj ���l��)�D&Q>�p?�f>�"u>��3��f8���P�h����f|>�26?�඾�R9�\�u�k�H�-Vݾ�+M>x��>,mD�jh�����]�Ri��{=;m:?�?�t��4���[�u��3��1?R>t \>^,=l9�=�4M>��b�Zǽ%H���-=��=��^>v�?w0*>�A�b'�>X�k������E�>X��>���<��h?��5?`���nO�z����1��İ>Y�?���>�k<�ƽ��@����>�"�>�=M-�=�gy��貾�u5>�EV�e���(�C��9�<vd����p>3z>?���M@����<��~?@~��㈿��V���pD?�,?J�=(�E<D�"�{���$=��4�?9�@=j�?;�	���V���?+B�?���H��=fy�>Fӫ>�ξ��L�
�? ƽq����	��0#�xO�?��?��/��ȋ�l��$>�X%?��Ӿ�k�>����Q��T���9z�bX�<��>^(F?���G�c�ŀ8���?�?���|���dȿ�v��Q�>I��?� �?P�l�z�����?����>��?��X?4�`>^o־v�L�?��>��=?/1N?6m�>�j���BJ?:ɸ?G�?n��=rܩ?J'�?��e;�|u>m��N�Y��9�?E�����>G�	>�1���R���Cp��������I1�����>��<��>`)1��nݾ�;_=��=������=���>��>|�g>x�>Y
'??�N<\����Q;�4߾��*�I�K?���?����1n�V8�<S��=��^��)?�M4?һ[�+�Ͼ?ר>޺\?5À?�[?Db�>#��U<���翿�}��Ԗ�<��K>�0�>YE�>����RK>g�Ծ�5D�o�>OΗ>���Aھ:.���򢻏@�>�d!?��>~�=ā ?|�#?_�i>@�>}vE��G����E�X�>sL�>??�	?8�?|���I3�'����Ρ�!_[�|qN>��x?�P?�r�>�~��1e����B�H�wT����?��g?�}�4�?z�?bu??9�A?�-f>����׾���@�>��!?��� oA�E&����o?�C?���>�ꔽ�^ѽ,7��>�Y���=�?�m\?��&?���`���¾^C�<_"�9.��m�;�]W���>�&>������=��>;��=�
n��m6�n�Y<�T�=��>�m�=��7�����WC"?�?�;PF�� ���
y��1��!�>�o�> �	�ńo?Ë�=,�@�2'������jբ���~?ᓹ?S֌?0��Ek��wR?>�D?�?.�>��#����c������-W�s�F��W�d�>��=D~ξQ������Ŋ���\���Q�6i?���>��?�?	?��C>P=�>�����X(����$�ﾥrs��#��S@���}���_���b�'�gξ�����'�>'o����>f�?M��> f�>*)�>��R�'?�>|�1>7��>�C�>�h>�8>���=�:�Sֽ�R?�LľN� ��?��Z���	�E?e]?�4�>i}e�}Ճ��r��t?ٍ�?.��?.f>��h�(�2����>w??��v�PJ?�[^=�<�2�6��+gԽ:��<K.��Z�}>_�Լ��9P�*ͬ�b<	?;~	?���=���SB���c��?a1>���?�#-?9��S�J�����I�+�=����9ӽ���߀6�'{_��v�*�w�C�u��&�7�<�?�?��B��~
�<�B��q�{�x�M��>ɛ ?��=5��>���=�|��U.:�m�o��)����51?�_�?�b�>�rJ?��<?�M?�J?��>��>_Ц�^< ?�}�:~.�><�>r�9?y'0?N1?�?��*?��f>}�������׾�%?��?d?��?��?�T��"8ǽ���~p���z�mv����o=B��<Sx׽�n�2gs=�RZ>�s0?Qf��Z�)�+o߾6�>׳X?���>�z�4oY���_�ؓ�R��>��q?��-?W����9[n�lb��R�?Q�*�8W�;��=1�<����<ѽ|虻�?9=�n�3�� �3K̽�`[�05={�Ƚ�y<Ա��4z��3Vs����>?�rt>i�l>Ց�"���i!�i��=�9(>��g>��@>��ǾD�������h��Ux>�T�?��?�zF=�l�=ܮ>�������`K��\Ҿ�L6<�?)�?�S?
��?��-?	�?��>����������7��G'?m!,?��>�����ʾ��ۉ3�ܝ?s[?�<a���c;)�Đ¾|�Խ��>�[/�U/~����"D�0ꅻ�������?濝?�A�c�6�y������[��Z�C?�!�>�X�>G�>=�)�U�g�s%�\1;>��>TR?gv�>BT?�~?�P^?�)W>E?�dR��5ɘ���<��>��A?��?�y�?� �?g!�>��>��$���辡w�#�ϼ�T��V��_�\�Z%?>a�>�>���>�B#>F�Խm���B�>�'G=G�q>��>�>���>�i�>�;�<KtD?���>-�ƾA$��(��#g��R�
=V<�?��?5&H?�( >��?�E�l��y4�>*F�?�@�?Q(?n~�w�>K�����x�����^�>���>��>�Z���$�<��@>��>��>7��� ����~=>�?��,?6}<��ſ?oq�(tq��뗾=UH<�����[d�!����#[��X�=�;�� p�
����\������u��p����z��k�{���>h��=i��=
b�=���<h̼NV�<GbL=i�<j=�vr��Re<��7���˻K��Q�D��T<I=X<�Kپ_ �?�F?�{3?��G?�	l>k5?>������>�����?iݚ=��Aվ� ������@���y꾣��X�n�	믾_�>˧6��C%>?�'>pG�={��=�K>^�<=Ԥ�=5��<I0Q=˥�=���=�}�=�M�=NI>�%>5�t?g�GȀ�kp��u=S5?��z>B4=�{��xc?x��=u�������-
	�E܎?[ �?H��?�(�>&6��A�^>s���fE����-����=ov>�{��v&�>�d>��"��6����o��А?�v@8�D?$���:���'7r>�:>��>r�W�k�*�;���M!��#2�BS1?��A�qg���9�>7q�<4F��*Ǿ:0ȼa�>���=0Uֽ�~K�%��=$Z���߀<B�=w$Z>m�>V_W=��a�l�a>��=���=��=������<;x��RP��m�=���>FSU>��>�}?�0?4�c?���>]�p�\о�'���3�>���=ڱ>C�=F>���>_%8?�D?��K?]̱><z�==��>�y�>��,�a(n�>~�e���6�<��?�ц?��>DK<XTC�P$�+%>���ý6+?�51?kY	?qk�>����Iֿ�r�ZjJ��%Ƚ�\4>f>? �Iǽ�H!=�H�K���=o��>q��>��}>Y�=`�>��>��> �q=C�S=��>5N^�zps=�x�=P�[�:�����=��/�9p< �r>1�%��\��aG<���� ���s�@<��l=�3?��a>���>��=H(���o5>V2��Z`R���
>򯟾S�R�i�l�|"w�O���>�xY5>vr�=���5���(?~,�=/�>ޟ�?��s?�|�>�'@�a)��꛿y��~6��̎�=�Ч���u��D�~�_�/�G�����>�ߎ>��>k�l>3,�`"?�eDx=��� n5��>�V����t<��3q��=��p��i�
�̺|�D?D��`��="~?�I?�ُ?�f�>�Y���jؾC0>C���y=u�iIq�N����?x'?��>C�;D��þ�2���K�>�w�gp�+����^ �����\���\H�>1���z۾��%�T1����1�E�� ��C��>��K?>˭?�r�*兿.eM��U���<��?��O?x�>�7?�r?GVݽ@= ��򹾠U=��o?)��?���?
� >��=D=׽wu�>�]	?�ו?D��?Zqq?��D����>ч<�C>z���=���=��p=�'�=�x?��?x�?�����q>辀7��J�m��@D=&I�=�؏>s@�>�c>�j�=�bS=�Ǭ=�)\>;Р>���>]�T>{K�>(I�>�Qƾ/\���1C?��>�>�>p ?K|>�K��>��B�=K�<����|䰾AV"����=�=>"r=����B�<�ҙ�>�xп�d�?T�>;��vo?x�'��N�o�=L �=d\�<`L?G��=8��>�]�>�G�>w�=�3F>�Nx>��ݾ�I>�l��L#�柄��o|����z֊>����]���|I��&4��*�Ϥ��R���Xd���w���?��]����?: ��O������������>�>(7?���������ޖ>
�>�]'>�d��հ�S@��_����?w&�?z�b>)n�>��W?��?�!1�_�3���Z�Lxu���@��7e�jr`��э�񚁿�
�|#��o|_?]�x?pNA?�B�<`5z>���?2/&�u=�����>\/��o;�]�?=_��>bm��Ca�ӒӾ�4þzq�e�E>bWo?d��?��?��T��As��/>`D;?ؔ/?��q?��/?��9?8c�*�(?�->vj?d�?��5?|�0?�%?��/>���=�U���(=����犾�*ս=�ν�����>=���=P6�;�%�;��=���<�Q�n��iӺ������<��<=�D�=w��=�Ȧ>�]?��>��>m�7?c����7�!?��j�/?� ;=����ĉ�������->*�j?u�? vZ?V]a>��A�"�B�r�>�(�>OD$>�]>Sv�>e�(F����=�$>��>�Z�=� M��ـ�!t	��W��W��<_� >N�>���>C�=|6/>)��|^��DD>b��C�F��Q���?�h#N��	о��>C]?�4?@��=����Sq���4���oM?:sB?�{W?2�~?��=�Ӿ�9��v��m�D��>A>�^���'���T��]U��	g��~�#>v��¾̚`>ZW������O��ti�3����P�3%��{<Y�%�sNžӠ��ü�=
kj>$�����o������W?v��=��*E�����n2�=���>u��>:SM>���rL�e��^]<�7
?���> �ӽ��羾�F������>N�F?ca?�L�?��|��qq���F�?���Y����-#?�t�>��?�@>��=aٰ�ʽ��Dc�E_C��r�>N��>��ckI�s ��F��c�&�dڎ>0?	�!>� ?��Q?M 
?d"^?��(?TJ?�ϐ>tð�bH��i ?|��?��{=��߽�D��?��`B��[�>��#?����9�>��?w�?�i?�oO?i�
?�/�=���:��>Wt�>L�V�oi����o>�gK?��>K(M?:�~?�G>c�-��L���Hཚ��=`�B>�=6?ץ)?��?C��>C� ?�亾���<*	�>
*]?���?Li?���=���>MQ&>p�>�#	>��>G��>��?HI?��o?,�Z?U^�>��<\�r��p���.��\�\�� <���=�=�=�����;H�߳P�`��=��=�Sr<��;�W��#j��>����z=v�>'��>�������<�׷��ξ�%?>Mg>��̾a�
�y������>.P�>��>':�=�O��g���>�>��?�1� 7P?�|`>�C?B����ň�#�"�Aq����>�7k?a�>z�]������G|�?wp=��:?��&?y 2��ŏb?8>]?Hs󾼌=�Q¾rOb�3�羚P?�
?H�Je�>��~?qr?�v�>��e��n�	�� b�Ug�nj�=75�>dm�`De�T^�>+7?���>e>���=�_۾Ջv�*>��96?^Ԍ?��?܊?�*>Otn���߿UI���.���^?�@�>q��n�#?�����о/���W���ғ߾
ꪾdɬ��ڔ��ڥ���#��6��d�׽��=��?��r?]dq?>�_?Ӽ �݆d��z^����+�U�]�����E�gID�m�B�n�n���Q��H���w�R=����@��>�?�"a?Ƙ���/?����e�(��牾X�K�Y��<D���XD�0����=�=�G��3�R����4'?���>�?��T?2GQ�V�Q���S��8�P[���a�����=���>`�>��=�jw��/��{���e��,�=]�>>Z�o?'�V?�q?ݑ��v�������[ �,jn>ǾpV�>���=ܧ�>��(=�+ǽ��DY9�<qw���$���������%=>�R?��=>f�?>t(�?
4�>�3E�c�p鈾M,0���⽱ �>X��?iY�>�m> ��������>�4o?�r�>��>;ڑ�;�&�ìu��2�����>���>�<?¿p>ū,�	-\��D���ʌ���6�KS�=*�e?}6���TQ�
�t>�AM?��<�+;5צ>3�/��V���Z�B��>í?@�=�_.>+�˾E��uu��(���?)??E?�Ւ�?�*�E�~>��!? ��>M��>��?���>b#þ$$%�Z�?�_?�,J?a�@?b��>��=�ð�� Ƚ.�&�/�,=�|�>��Z>�l=FQ�=���P\�E��5sE=�i�=�ͼ`��Ò<��M�P<��<�4>˟ܿ�@���Ͼl������`�u���{���������о�>����0��/��% ��s���f�筵��^�t��?��?�v��,��xq������ှD/>�T���*���X��]:�t�¾�d��y�+�@��c��S��x?滋�~�¿Z&���k��:	?�;%? $?�����+��$O�HI^>]��=zN6=������Z�¿�&���\?�N?V����!���>4�>0��>��4>����?�x�]<� ?*�F?���>v���ݿ@����<�v�?�@�tJ?� 9��I��9D=�0�>��,?7�a>��6��^������>�^�?h�i?����>�*5�;{�\?+Y>O�(��_N��=>ߦ=�i��j�m�>�U�>=3B���N�����&>���>-;�<�mŽ�r�TYٽ�u@=�Kh����<�+�?ߺZ�RX�')#�(�w�2C�=��S?�Ԙ>��=&@6?�RO��tҿga�C�S?�z�?���?#�6?W�����>m�ھ��I?�}>?�х>D5���m��s>Aү�N�V�S����bR����=���>�>�\&��
�%�^��������=�n�+ſk$!�7��~I��Q���|<���0����h�2m̾��o�XF���I=�	>�80>7�~>��>�	.>��j?0fq?W"�>��c=l{�#Z��2���O���X��V:*��VR���ԽK�*������V徠��O���3���==��8�=Z�Q��@��-\#��)d���B���,?" >�3ʾ��N���%<�ľK���]��,���D̾{�2�k�m�.��?��@?���G�U�
�A�PӮ�b�V?�����*���D�=]�Ƽ+0=�z�>ߕ=���(w2�?�Q��,?�*!?�#���H��FTG>F����=j+?�>T�w=>��&?cJ@�$��+ă>��'>[n�>���>��
>�.�����s�?�P?�	Ͻۻ�����>񜼾��S��Q�=><%>X�2���:�9�T>��<.�e�b�[=}/e��x<�#A?嫌>�A.��t�{���w�;d�=��S??��>�>��=?&DY?~�=*b�u�B�#�}�㺾�K?�^?i3>
������-���|?c�`?��>��b�w���/�C ���-?8�k?ޱF?\_Ǽ���������$K?��z?�����]����]}>��>1�>��=d�Ӿ��X>n�)?�^�E���*w��LyK�qG�?P�?� �?j#���4?<G?�+<?�?ײ����Ľ`�?=u�E�	�v�ڗ?��s�v�B��S��m뽜� ?�d?�S?��4��C���=8[���.�?��?�H˾r�=��"�{�<޾G֗���>���1�����ܾ�z.�@ȹ��g������-����>S @��o�>��;�㿽ҿ�sy�.��o�t��t�>k��>�jd�������X���p�y�@��)>�c+!�UȢ>(>%��a3��k�{���;�>����>)��nv�>73U��<��P���Le1<���>���>\2�>E����螙?nB���ο"}��mF���X?�,�?�=�?�a?�4<�cv���z���+�u�F?�ks?��Y?tA���[�2�6�j?���_�{X4�'7D�J�S>a�2?��>s�-�G�~=��>���>�P>��-�h�ÿLh��$���q�?}5�?2��;��>][�?�t*?���s��B_��9*�4�>�m�A?�3>������!��=�鎓��E	?n/?W	����W�_?&�a�N�p���-���ƽ�ۡ>��0�f\��M�����Xe����@y����?M^�?f�?ص�� #�_6%?%�>e����8Ǿ{�<���>�(�>�)N>�G_���u>����:�i	>���?�~�?Oj?���������U>
�}?1�>@�?� �==k�>܄�=�Һ�Ɯڻ��1>[��=�����?�K?O��>#r�=u�D�T�/�pIE��N�+} ��B����>M'[?��J?�\>���A�P��q��������m�'H���k���*�,>�7>ܭ>�69��Ѿ*�+?
�D�ELӿ˕��`�C���6?F�i>��=����(پ�i����X?~'>]�4�I(��$mq�R�8�n�?P��?X��>�!�)��w�'>���>Qӏ>����C����ĵ����=fU<?�l�(��.��� N�>�*�?i�?��?l~���?������n�w�K����p�=[?�H徳5>�v�>1��=ʃy�^檿�q�>���?1��?���>�Da?�l��0�-�>2��>�]?WA?�pM=1�˾� c>��?�K��d����o�V?+*@r@m�`?=�����<���9˾���ns=��v=�'�=+|��zw�=��=6�N�Z���=.H�>p�>�HW>fx$>r�>پ�=I���f �+�Ŀ�t��\�M�	��Rl�V���h��d:�����j�о ������AQ�fi���P�ϯ�UD��z"�=!�U?�0R?u-p?� ?E u��k>������<d{#���=��>Y62?�>L?v*?�Ɣ=�X���d�lw��ZN��0퇾�g�>�I>l'�> ��>�(�>����}I>�2>>v�>YO>[ (=�֊�ը=��N>Q7�>]��>�T�>��>~
>@����뭿�h��< ���=�N��?�́���J�����e��Qە���=ߔ9?l��=����[EϿ��t.N?����!h�i�>����=:�:?��F?/ӌ>%图v����=q�m���f�v�->&C)�����-�#��f^>+Y(?�f>�2u>
�3�]c8���P�P����h|>~16?g鶾�*9�c�u�@�H�YݾN=M>���>\GE��j�9����Fui���{=n:?��?�&���簾�u�6��YR>I\>T�=�[�=�LM>-c���ƽ�H�r7.=���=�^>���>`9^>vٹ<ƍ�>-��������d�>h�C>��	>�C?�V%?�'���Ľ���^�:�e�Q>"��>ۄ~>��>KyS�z� >/��>�f_>���������&��Ga>��0;��l�ή�,�=�yy����=�_�=� �I67�(�<�~?���#䈿�뾺d���lD?U+?� �=��F<��"�A ���H��F�?p�@m�?��	��V�4�?�@�?��H��=}�>׫>�ξ,�L�ޱ?��Ž-Ǣ�Ŕ	�M)#�hS�?��?��/�Xʋ�7l�z6>�^%?�Ӿ�^�>���J��\|�{.w��l�<���>�dA?�����1��ϔ��%?�o?�����@��2.Ŀ�m�R��>���?�X�?��}�[W��J�)�@?��?�C:?�	�<����䎾5d.>��/?�@?��>��.��*���>?��?��?P7>��?��?pU�>&�S>M,���տ��4���?{���i8�>w�=���A���s��[��)w��/�y��>�U�<BҚ>z�̷�-�=�[V=}]d�3%�=��>�?o�>N��>��]?��?˂r<�S������Ȳݾ��K?���?��R4n�;��<���=��^��(?SG4?��[���Ͼ�Ө>Ӻ\?|À?�[?5^�>/��>���忿$}��r��< �K>�2�>
G�>x ���GK>��Ծ2D��o�>�ϗ>����=ھ�*��F@���B�>{d!?���>mҮ=�A ?��#?Ժh>Y��>�HE�qA���E����>��>�?̒~?�?�����G3�6����Ρ��r[�b�M>��x?&@?�8�>Y]��gP��8<�@�C�h��F��?��f?���?�A�?�|??��A?�%e>��4ؾ�7��XT�>�v!?*��ϵ@���'�@��Ơ?�L?*�>hۖ��	ٽ�;̼�z�����?Fm[?�M#?4=�a��������<ޏ ���`f�;�<"�ͩ>">�^����=S>�u�=��o���6��v<J��=���>�4�=�7������,?��q��½;�>�z��A8�;�>A1�����P�?�ɾ�0��t譿����DtD<��?h�?kMu?��h���p�;Q?$��?��?riJ>�u���ܾ�춾�獾M��gھ؊}>M�>�5����N�����q���Ӏ�����$?��>'	?�i�>x�u>�>O���n6�EDӾ��!�~�����@�����B����|���;�'�P�E�˾-ԃ�%<�>=C*����> `?&��>wE>tu�>�����>\�`>s�t>[k�>��a>�>|>J,N=���	�Q?�þg�$�n��u[��%D?�b?!��>I6������5���a)?��?�J�?%�g>�e���&�R�?Zj?%���R}?�=uD���ż�3˾� #���3�^2�a΍>)V��e+6�Z>E��&l����>��?)��x���:ڽGt��	@n=7:�?(�9?��0���D��r��a��D�������I��s��$�og� ���	K�Y���7)��,=Mu)?���?�	�����^���t��L��x>Џ�>&��>���>*5A>9/���1��P�5�$���y���>.z�?���>��I?��;?0qP?�lL?���>�_�>�*��pf�>%��;���>�>֙9?�-?�<0?�v?�s+?�@c>�x������#�ؾ�?ѣ?�K??ܱ?7߅�wUý@��5�e��y� ����
�=���<h�׽^�t���T=�T>p7?���=< 󾳊V���	?���>}?�N?�ؾ�%�?Vk��L�>�GU?%l?~������	>��)+��e�?�.{��cj<�
�>��@<4{�=�\ �Q�>��=vE=��4=r���m��ߡ�=XEd=gO�=D+j<�f�<q|f=�'0=P��>J�?�p�>�C�>��� �3����=�X>y�R>�3>*
پ�v��W$��^�g��oy>~q�?X{�?pf= ��=* �=�j���_��C���ٽ�g��<��?>A#?OT?���?;�=?�b#?[�>���yM��h�����U�?,?���>���\�ʾI�����3���?j�?�;a�mX�OB)�L.¾jҽFz>�b/�I>~�������C��~:�z�����y�?�?��B���6�r�������Q����C?���>��>t��>-�)�j�g�����:>���>��Q?}�>Ha?y�?a�K?N-�>��D��+����*�>�1�=U`\? |o?�.�?��?�o�>`1�=��^�u"�����Qt��g�� ���fL>XT>列>�͠>M�->�ʱ=T?ҽ���<�&��V;>�@�>��>
r�>�g�>�.Q>�}��N<?`"�>�:��	���(`|�־����<��[?Ԉ?��J?�|�=)wȾ5Y�k���-N?�?r�?'�8?�q��T1>�z�������;��Ƿ>P��>���>�9N�E�X>tR�=�z�>s2>�=S���ؾ�;;�s�>��L?f�0?�_���ſkp��r�����qMJ<^��Fvd�D��Ni[����=�������F����]]����o����ݵ�1_��soz��2�>+�=U��=S��=:�<�K׼�(�<Z�L=�ґ<��=S�u��j<��8�f���׈�\�?��7M<*�H=����y?@'R?>9?V�=?�ȋ>��%>�b�ʳ >�����%?J�<N*���Z־��4����A�q���Ӿ�~��\x�fȤ�S?
>b5�׃>��r>�(/>Q0�Z6�=,�e��$>#�=�|=.q	>�)�=�ń=��=e�>��>�rv?c0v�̓��,���/=��
?�U�>����u��׊U?�RY<�V��"b������k�?g� @���?�T?$Pо���>	��\�>�
���h��?u>H��>lb���7>9�[>~<��~��S���6��?��?�JI?�|�8Ź�)�s>(�>9F�>��8�z$�k�>�ƾ<�P��3$?�-$����� >�QZ>����پE">p��=��<P���7�Q��=i��k7����"��\�>�d�>j�K>(��#��=��=
H>�?9>ϟ���뽣�>�O0>N��>�K�>b�=���>��?��D?Y�n?g�> O�UQ�NA;[��>;�`����>Mϔ<m}=�>��F?0?��(?C�>���=Y�>���>0�K�����	���Ѿ-
�\�?Ӆ?�>�~�;J�޽�!��4�����2?��$?I�>1�>(:�C��B�)�u�%���콑VW�ʱ�=��8�U:!����|�t�Ĵ��X�=�>�$?,��>J?v>b�>T2(>���>�� >;LW=�B=ڿ���7�;�Sb=�J�=��׻k��<�	�M��=�� =M�3�R~�z���I��<�67���<Q�8<R��>��>��?Ֆ*�֬��t�3>�I����F�K�>qX���hk��[��m�������;&Jv>�Y�=���������?rL�>��>	��?�*v?D��=�>����P��Ӂ�;����:H>�6�<]�z�R�ơq���0������>5��>��>�j>�F+���?��0v=�޾�	5��>MX��Η��M��:p�H����̟�:�h���k���D?���m��=�*|?�ZI? 
�?i�>+|���lؾ&�2>-'}��7=�u��7y�����=�?��&?�N�>cm龄=E���˾�ִ�X9�>tH��O�����S0�L������a�>ɫ�\ξ�3�I����T����B�X�s�~�>��N?�8�?�a�<���.O�>�������?.�e?g��>�k?d�?����������=j"o?�w�?5�?%�>R��=2Z��6��>��?`�?�͐?q?(=�~��>�g<̀ >��t��o�=
�=���=���=B�?А?�M	?YR��������ﾚ[�
3=���=&X�>A �>�r>qh�=�s�=�[�=ؔ`>7G�>�a�>)rd>��>�E�>���6[־�\E?k��>IN0>Lna?C��>�2޽3�F�:���V3R>?�ԾwUi��&�m�=��>�V=h�����j�k]�>�ȿ�W�?r��>S�/��x4?���9�J� ��>X. <�3>[��>a����>}��>��>.�=�r>��a>_ ̾q�>h����%��X�IU�cϲ�t��>%Z����E�����ܽ��K���/�羕lf�bi�бC�K?<�Y�?�5���h���&�d[�/?.��>5�@?yC����Ž��=��?�3�>�������Д�Hھ���?��?KF>�ĩ>�l?��1?W�l���qh�����T�v�s�3�N�����%�|��M�?-� SR?�#]?D-?�yH=iF�>a��?�<�cp¾��>q?��X�z�>H6�>ƴ���a��ej��+�ľ��C��"w>�`??]}?��?����k��_'>}:?�1?Rt?��1?��;?Tb�x�$?`�2>�@?�L?�P5?�7/?�
?�1>���=��ǻ3*=&a���Ȋ�q4ѽ;ʽP��~�2=@}=h��|�<f�=a��<+i�\Fּ��;�$��;/�<f:=�Ѣ=���=���>>�]?Qz�>@Ʌ>%&8?jm�`8��P��I�.?��G=La��t���LH��K��R>�j?�~�?�&Z?e|c>�X?�2CD�z�>�s�>�(>e�\>�C�>���{>C�� �=��>��>�Ģ=��L�혀��'�q���ķ�<�>���>�3|>�=��"�'>D����?z�$�d>�sR�t����S�1�G�k�1�4�v���>`�K?��?4p�=�]龟햽"`f��F)?�f<?vUM?��?%��=��۾��9���J�̏��<�>Z�<	��3���� ��D�:�N�9�>s>�D��vΡ�v�g>����v���t��B��l��*�?=>u���=-�&�����I�I���=�@>����Iz��?���9���;T?�>�=uw���A}�?$��>�Ԥ>�>�_;=T5 ��N��=�����=��>/މ>�
T�"��H�L�́�M�~>��J?��b?�K�?{���x�q�5-O�����s��9�?D?t�>��?34`>Z�=c���z��[j�x=H����>+4�>��!�[�/�ۃ���g��,`.��r�>�}?�|�=*o?]�R?Da?�]?��1?׷?�֛>l<���ž��>��}?d�>am>�=��UDi���]���E?�a?�K��̏�>�-?� %?�&9?W��?,?�U>&����E�q��>�O�=~Xp���#�W>��6?]K5>��u?h��?�C>�!�Rþ����俽�X �"�?_-?9y ?P�?��>�ܡ��4=�T�>��b?+�?.�o?��=��?�J2>���>���=�Y�>�#�>��?�>O?q�s?�K?�}�>�Q�<*���|����r���N�r��;�H<��x=9���is�T��t�<n�;3���S;z��f��~�G�ȗ���t�;��>έ�>`q��9��=q���E��	��>�Yf>y�R��Z�=�v =��>�>��>A��<��0�= 	�>���>B�:�S�j? ��=��>���<�ձ�"+�"6>���>-��?�r?�掿Xض��酿�E�=�V?}�?�"�w�T�U�b?��]?�d�I=���þ��b�ٌ�?�O?��
?j�G���>��~?��q?��>�e��9n�:���Db���j�yѶ=$q�>^Y�{�d��>�>�7?*J�>
�b>�*�=�u۾��w��o���?_�?,�?���?�-*>��n�K4�G��q��u7p?Z��>����p$?�6[�T�ྉ����y��=�žƘ��x�ɾa捾j3���-��Hl������<�l?��u?��c?Wwe?O	��X��bc�L��U����K	��A��A���M����+�����ٱ��<=�Y����C���?�%?�:�/��>�D��8:޾mDž�NL>cC���v���I�<|=X�hv�=�7�=��K���4��b����"?^��>ث�>��4?T�L�/�':�KiK��n��R�=�c�>@�>Q��>����Qh��(,�]־�<���N��-�>�q?�<c?᠂?I�S�a O�Ap��s�8���>(C���>���>_l�>�>�< >�T��GI�������1���z�P� �o��=m�a?1)1>�B>��?;�>Խ8��Ҕ��ѽre���5;��>�C�?�Y�>���>��i�J5&�<��>1m?���>2��>�狾��!��{���Ž��>�ծ>a ?g�l>G.��`[�G���Q���8��)�=:h?&[��x|_��W�>aQ?��:��:<���>�w��z!����%�s�>J�?��=&�:>�ž�es{�W��Ŷ(?�,?�萾�p)��>`� ?���>y�>N�?뛛>�H¾8ho:?k|^?�EJ?�A?l�>��=�����ƽ��'��G-=>�>�Y> �o=�=|M�4Y�M��MD=�t�=��ļ@��Og�;��ż��T<��<��3>�׿6�J���ݾSO-�ݮξ�����L*�,ܽ���F��n�龟���K�p��7
�S�g���
���M�;$��;�u�r��?�?� ��T��%���i��٫��Ȉ>�����@���ԋ<S��ݦ�(;t_��=���w��^a�.?"-,�$󽿗�����V�!�>[�,?ζ?쾶��=�z����>hD�=�f�<]FѾ�U����������vI?��>=Ҿc���?��>q�V>D,3>��d�����;�2?�C?��>����3ٿȿ�a�=~� @Ȫ@��A?3�)��	��YR=i�>��?��K>�C1�|3��.����>zr�?�V�?�V=
wW�F��3�c?�<LC�y*��.�=D�=���<�a�/I>:��>\���:��vϽ��>>#z�>PH1����ÌZ�gD�<�d>�uϽY��Ԅ?�s\���e�^�/�#J���m>��T?��>6١=(�,?�>H�p�Ͽ �\�v�`?�+�?;��?��(?������>t�ܾy�M?�e6?��>#{&�U�t����=�lݼ����~㾡V����=���>z�>��+�,��*�O������=5��lǿ��{9����=��]9����Rӽ��ƽ�qټQ���	}��=��υ=��>�b]>��>�8?>�(I>��`?mn?�٧>[�=��'�����qx��y4����~��d�E��~�yژ�Z�����7���K���ܿ�܄;��ˎ=oT��&���E)��mY�pu)�m�?���=�赾\C^�`�_=9���ی���9��Ja��¾�/;���i�Q�?��K?�`����j��i#�\a��؟�Z�P?�̽Ŗ��վ��=u=|��=�̼>�==0�[lG��K�&s0?kZ?͊���[��d**>�Ӽ=��+?2�?��\<�2�>OD%?�*�66�E[>Đ3>֣>#��>�F	>��B۽b�?��T?�������ې>U]��!�z��a=O">�;5����c�[>#��<��{�V�!L��诼<�=?��^>��G�׆���3�ҙ�U}t>�d?� �>�k�>*��?�B?ֿ=ʾ�T�AK���=`?ӂG?���>�F���|��E�.u?}�?0��=g����ǭL���)�Y�?Pޅ?7?)<�=ݣX��앿��o�X?({n?>
V�U0��&_ʾWD㼽�>A�>��>��5��>�A�>��ƾʼ����ɿ�f9�z�?�@��?a�9�kR�=գ#���?�P�>� N>M��� �����2��=0��>�f�/�O���ؾ�(��.1? i?ϱ�>�3��QNԾ���=\����0�?I܇?5ģ�>�=&���L}�����v>�b{�=<�=��c��D��W2������U�^0��/P�����>�@�(�Z��>a:w�W�ۿ��ο�뉿����s����Y?�kK>߹����ɾ�2x�jr�E�N�lT;���I���>>�Õ�������{�q;�y��� �>��6&�>)xT�6���w��`v4<��>s��>ī�>+R��� ��ř?5���3ο袞������X?Z�?`i�?�w?A�<<��w��{����)G?�s?!Z?*�%�R�]��7�+j?L���fb^���2�2:F��Or>��6?B �>��-��{%=g">Y��>o>'<*���¿�Ѵ�����!��?��?��� ?Pl�?��%?���扚�tg��%��#<�!F?�BL>p$ľ��#�D :������?3[1?�� �]�_?+�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?ֵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>_H_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�"�>��?b��=�a�>�c�=$��-��d#>�.�=�>���?t�M?oK�>}g�=��8�V/�\F�)HR�/#���C�,�>(�a?m�L?aEb>G��Q2��!��zͽ�\1��G��T@���,�N�߽@&5>��=>>y�D�jӾ�/ ?���ο�x��b����>?*$�>��>��L졾�=%��?�^�=�<�����)��M�X�M��?'u�?�#?�,�=Ȱ���>�n?"��>�^V�,���MҾ|�g<��L?6Nx�Ai��q�x�qt:>2�?�?@�K�?`\���>�ڸ��怿ϭe�c4��ӧ��%>��L?����<��>z?L�u�:~�1�����]���>�2�?z:�?�#�>r�O?��`���K�:9�=~n�>~bE?�i�>ȇ*�+7��o>s��>�z9�A���!�ʈ+?��@��@�(X?!ݢ���忕������9�����=�Y=7$>����v�J�ߓL=��=��ټD�>3Ú>d�Y>�� >K>�gO>�R�=�:��b��e���������G��3۾5������:��ޚ��Ĥ������D��7�gA�;�B5��4�����4�[=g�V?	�k?�?M�>�+Z�D�>=.�(���w�A^��>��>�[7?�j?Q�g?{V=m����v��w������'	f����>_R>b��>s�>>�>��=�U>ָU>j�6>�<�=Q�=��мm#�=d�z>+��>p��>��>6"(>g�%>���������{�(n�^�Ƽ���?U����5�G�����u�l4���M�=!m2?�>g���7�ѿ�n��>H?���#5��U ���-���(?�L?�Ii>v�g��-�`Y�=� ߽��e��*>��^���.�^av>�@&?�f>�u>s�3�p8���P��y���z|>�36?ⶾ�69�W�u�U�H��Yݾ�QM>�ʾ>�C��k�,���>��ai���{=�s:?Ǆ?򈳽�ܰ�2�u��2���kR>8\>�=�o�=�PM>�c�_�ƽ�+H��.=��=~�^>g�>��h>됎<-�>����7`���u�>�ˊ>�`*>#X?�Z=?��ŽF��I���>[��P>(i�>�6�>�t>T�K��8�=���>r�O>��=�ɽ<{ؽ�(��G>@�����E��f��Ca�==ͽ�p�=��=2d� �>��
>=�~?���䈿�뾂d���lD?Y+? �=W�F<��"�= ��@H��=�?d�@�l�?��	��V��?�@�?���s��=�|�>�֫>)ξ��L�ܱ?{�Ž8Ǣ���	��)#�SS�?r�?s�/�Gʋ�l��6>_%?�Ӿl��>�52���މ��S���^=	6�>�G?������@5\���?�q�>4��8��zȿxo��4�>0��?eœ?s�r�IᖿL�$�� ?�*�?Y@J?&{0>�v���y��!�>��A?�1?cVX>�!�F�%�_j?��?T��?Bk�=�}�?�'�?M�>� v<ǘ�e\ǿQ�j�@?=ꌾ�̪>����Łݾjy־yy�� c�rg��(�ˠc>���<y��>�}R��վ:�R=�'��L�r�].�1r�>7v�>ۆ|>v��>�5?v�?�?>R�Y���]���Ӿ����+�K?u��?���92n�_T�<|��=x�^�w'?sJ4?n[���Ͼ�ը>�\?L?�[?5d�>���*>��迿�}�����<G�K>[3�>+H�>�#��zEK>x�Ծ�3D��p�>�ϗ>���#?ھE-���x���A�>xe!?C��>�Ү=� ?�#?<�j>�$�>�]E��;��j�E���> ��>�L?��~?��?�ٹ�UX3����\䡿1�[��DN>��x?�Q?�Ε>_���V���W�C��lI��������?rg?�`录?[.�?3�??�A?B(f>:���ؾ��� ��>�!?W�m�A�:L&����?�O?���>�+����ս$(ּ���r��� ?&$\?<&?)���(a��¾<8�<G�"���T�Yb�;�D�N�>M�>���w��=>�ʰ=�Jm�,B6�+(g<�l�=}�>{��=�-7��n���X/?H82�TDԽ0��<yd\�1���b�>�?:>R���?O��d䅿�vJ���@�=,��?���?��?>�M��w�twV?�ܒ?@�?�>�#������喾"i���R��派�9�>3�p>��>h�ʾ����U�������ý�U�E??~�>�=?OA?���>dv�>=E׾NJ��߾ b�x�m�EE�(�F��9�D��=o���j��s1�w%׾7^��7S�>T�!�R4u>��>�P^>���>��>���=1v�>�q�=-B�>W;�>ڸs>t�>�=BH�=Yɦ�:-Q?�JϾLN���վ�?Ⱦ�_?*�s?��>V���冿�����/?E̊?���?��	>E\�L����?��?������?�3�=����[�ӽ~	�ܶ���2<�<���>|n,=�=4�(�X�3g��>�>���>$��=���k|{�O��}+�=dL�?��7?�&���E��"|� bs��8H�*_I��H�n�ɾ�9�~:n��\���r��~x�z$�܎��d%?႔?7�X��w��� f��`�U�>=?��,>v��>U q=pZ��1o-��$S���Q���E�>�`�?^]�>�uI?o<?{tP?�UL?p�>%j�>����6��>���;��>�>�9?��-?�F0?�v?#`+?T�b>ML������ؾ$�?�O?�?o?h?׶������`'���f��y������c�=�ƹ<�ؽK�s��pT=�	T>�%8?Ln���:��}��HT?��Y?d��>�N`=mo�Q|�����U>8sk?���>+���Bi��"$���>c:�?@{�\B@=?�>�@*>X���y�=�ߨ>}�������Z��*���>ع>�Op>��P<��%;�o�?r����=�>��?N��>$��>rՅ�/� �w��K�=z�X>�S>�>�Zپdo�����zh���x>�l�?���?�9g=�}�=
��=����j��$��񧽾7@�<�f?�G#?�T?P�?�~=?h^#?��>����8��f�����u�?k!,?
��>����ʾ��Ɖ3��?s[?s<a����;)���¾��Խ��>�[/�`/~����CD�녻���4��!��??�A�H�6��x�ʿ���[��m�C?"�>/Y�>i�>^�)���g��%��1;>N��>�R?4�>|�T?���?�Z�?�1>_L��壿B ��������=��???Ƅ?&ه?��?'_4?%��=����/��J�.�5�{���ֽ��?�u�>{�i>b�D>Z��>ϛ�>G�<�*м���"���=��9>��>���>B��>sr>����M	9?)V�>��Ͼ�Z����A¾��<A�u?��? 	L?EԵ;��7�m�Q�@
��>Lj�?d	�?�1?���46>����氾"q��p�>���>w�>ꀸ�m�=�� >��=>ܫ�>&p3���6�=/�}#->u-?WD6?�� ��&ƿ?�q���p�䗾|e�</���[<d��e��
?[���=�>��20��֩��+[����J���ۧ���̏{�~��>�R�=H��=?6�=.	�<7�ʼEw�<�NI=���<x=\�o�.Xz<&V8�����I������)\<�H=$��ɾ�|?"kI?E�+?C?�l>��>�頼�O�>���pg?<lX>�Z(����5�1�w����ޑ�D�ؾ"�׾��`�������>��]���>u�3>���=cĂ<���=��= �=s�����'=�E�=٨=�8�=u~�=��>O4>6�y?�A}��ц���2�)��<�:?��>o�i������v6?���<W-���x����9���k?��@e[�?��?[���z�>�%u���!>*�����=�j�	>^�|>���0]�>^��>����ݎ�h�`�,۹?S��?d^9?3���(���e�f>b�B>��=|�T���1���P�bX��[�S�!?� 9�l�žĔ�>��=����̾��<05>��=g�～tX�^�=[h���=�Cn=���>�&D>PƲ=������=tg=vg�=LH>���;��0"���7=.r�=��]>{3)>̔�>K�?1�2?��h?�^�>�\��R�ؾZ���^ؙ>�6�=���>=$�=77Q>�ƿ>F�??�^C?[G?��>��&=
��>B��>�1�!�n�OپY���ƈ;�?ㄈ?�_�>��;�IF����E>�B;��<a?��0?�w
?��>aC��������%�F�����޼�!�<ŋ��"��6B��h�W��O-9=���>�@�>@ū>��3>�u�=�'>�R�>d�>��=����#�=v��<�Wb��>�=R��=c��<]ý���<@ӿ�l�:=��2=<��=P�U=��%���/=ۿ�=��>�_{>���>2"<>�P��<h>�#׾�b��p>vB��"�7���u�v9���L��?�<Wh�>,��<V�g�5��\?-wY=��>���?�5m?W�>Լ�=8��1���@E��Mz�ĝ>z�+=�J���N���p���P�k����>�a�>qC�>} l>�,�c�?��\{=���%5����>J����T ������p��4���ݟ���h�T$繗hD?�>�����=�q}?=�I?��?@3�>@ܚ�˓׾t�0>@��^'=Fq��r�����Z�?��&?+h�>�˧D��A̾ľ��ҷ>�BI��O��ŕ��0�������r��>bા��о'3��d�������B��*r����>\�O?��?�-b�Y���PO�C��ZY��l?{g?��>rN?C?޵��{����j�=*�n?ĸ�?�:�?(�
>ν=���"�>�%	?T��?��?�{s?�x?��W�>���;-� >�����Z�=��>+�=/!�=�l?]�
?v�
?=���t�	������6:^����<�ơ=���>�|�>��r>=��=>Zg=7\�=�6\>4ݞ>Fӏ>��d>K�>
P�>ʧ̾����B?(�>e��>?'?_��>��>��@�4>������j���G�ґf=ʼ3>�,�=����dT����>��ʿ�D�?�G=�"��8�>F4����=pu�>��;>d�R��d?o	��j�>�>�^>�h�=���>�%~>��Ҿ��>�S"�=2D�)R��rо�|>�~��Z
%���	�&>�98H�f��k��H�i���,�=���<�#�?�����gk���(�ۮ�V?R�><6?����|���PU>t_�>�7�>ڑ�������qUιf�?��?�b>X
�>�$X?��?��1�4�*9[�w<v�� @�Y�e��_�
��k� ���}Ľ�&_?��w?3X@?��x<��z>���?/�%�B���a�>�.�]�<�^�N=[y�>�U���*b���Ӿ�¾
�IPF>�n?R��?s�?MYL��<K��H-><C9?-0?q?&]'?��+?�Ǒ��C4??/>�7?Ay
?�)9?�[.?�?��0>�>�=?
��Q(=�L��_�������ֽ:G���C=KA=�E��� �<�AH=�K<��á���v���3��;�9C=W�=�=3��>wL[?�y�>�ߋ>h6?Y�1��=�`\����;?� /=�Oy�O�������qR�r�>ңh?7�?$S?��S>��9���I�s><A>� >�^]>�#�>���P0���=�6>@F>匱=c���l���
�'��h�<X >�M�>AB}>5���g(>i�����x�e>^�Q�ِ���hO��hG�ڟ1�=M{��+�>��K?�|?��=��������g�&�)?�N;?}#N?SV�?~�=�|ھ��:�n�L�d#!���>�C�<�U[���w��%�;�_����'m>[ٟ�Ue��ņg>D�	� ��HUs�U\M��R�ܡp=�
��:=t_�4վB@o���=�L>[�� ��w������J?ە�=򋨾̕I��X��K��=�>�]�> c��s��GD>�^���*�\=;��>�>(����PF�.D �#>�&W?fS�?qB�?8��5����J����/��A	½y�?D"�>!N?�"�>o�>�Ӷ�?�Vd{�!�d��`�>3��>��g}M��M���ؾ��1��?�={L)?�I`>Բ?�y|?��6?�2b?�e?�+?x��>Xa�<s��� ?P��?S�>u�4�])��M�U�Y����>b��?zw��+�>i4?8~L?��k?�Z?�>�!*>hm��Xe�'qn>b�>>3}Z�w��α�=u#I?��?�?�?�=]C�,� h�����|�>�f?Bd!?�E^?�z�>�W	?iоW&����>��f?}�x?�aY?܍g=��>h�>Ew�>fe>��:>��>���>ÂZ?��?m�\?<��>6�<'o��Y ����aƽ)v�=N�?=cB̺�����������o�藮<~��<"�=��G�CDƽ�K:�7�V=[E�>Mc�>^B�����=!��>���֥><��>E�͔��7�=�U)>{g�=��>
rD>�a�I�=o��>�q�>m5���-?�6�>�Q-?*9�=��y��������>,� ?h�?� �>*.l�g���N�l��=��?��?�v~��`;���a?��^?�?��=��$¾�`��Z�ϻP?1�?�K�C��>��~?�7r?��><�i��Vn����/�b�_h�u��=d��>� ��=a�k��>�t6?٤�>}O^>[�=z�ݾ�tw��p��f�?B��?�I�?~z�?�*.>n��u࿹^����9(_?�k�>�J��f#?0;��Lо�*��Ğ��G�߾ʞ��Ϲ��dҔ��E����#��̃��|ݽ���=f?��r?<q?�_?m�z�c���^��e�jV�1�A��w�D���D�KC�:go�s���<��=����Q=Ņ�wu<��|�?��/?��|�>����l����ž��>3e�H���jѼRs���>ϼ�=��_��Nk�4_���a#?3�>H0�>�-?��]��5�;�e�/�������O=��>�T�>�V�>&"?��O��nL���}�L����9C����=�~?�LU?1�w?E��=ۍ4��O��p�����>Ku&��;>�	�>�R�>qU=���)i+��G�1H���A��c��ß����=ʬ�?Y�|>�m=�k�?J�>5�6��󛾜���B�,�s��Ю�>�֋?0�>kN�>�ؽ�LI����>�u?֎�>��>|�;X�����`Լ^��>��>�(
?���>�����L�{���፿�E?��a=#=b?� ���h���O>�~[?c ���|<���>�����&������-���>$�?�p�=��1>X������
�w��ٱ�H�#?k?a����(��p>8_?#}�>T�>S6�?�/�>�E��Zq�<�J?Z9d?��L?��;?,��>,@[=<��fdнl)��M=��~>�M>b��=�l	>��� _�	=�2�7=��=f�>��#н�<ο¼yp|<i�Y=Y�G>lIпxT7�FK�������"�R�򾺊����3 8��@�{�ž幁��䘼˼��\?�C?��V\�f��k�����?S��?��Z�)ϖ�y՛�\���mL�{�>��#��:t�>k��w<�E|��Q��oq�:�K�/��Y�1�W�D�'?巑�$�ǿZ����Dܾl ?A ?,�y?4��"��8��� >?[�<pN���뾅���G�οǧ����^?���>�
��R�����>���>�X>TMq>k��瞾&g�<��?b�-?���>�r�Жɿ]���Ǥ<���?�@��E?B�7�,[�|'A;n�>�{6?��>��I����zjO���M> Q�?�O?P�Y��Y����==��?���>ޅ)��[���h>�!�=��X�7
��ǙT>�3�>���;t����c<0�>"�>����t��G���>>����<��-��JȺ��w?�D;��F*�� ��J�� k=�J?�+�=g�k>+�Y?��g����-�^�l?F@|��?
�?`$ѾX�Y>@W���I?gTQ?5/q>�d=��	e��\=�>>�_>,���(�B?�=6�D>�p�>4u�����v��e�;O>�����ƿ� �����F�;8(�<�쥼�#+�5���z�"�-��w�l��f}�<K=8�>A\K>#�s>��4>�#M>F�_?�qo?,`�>���=W"�C���ľۣ:=_�c��I]�C;o���ƽ������gپ���b������Vоc=�0	�=�O��J����&��He�|�B���-?�9(>`^ξ��N�OM�;	P�������ߟ�iD����ʾ��2���l��'�?`�B?�����nQ��`�Q�u��Sɽ#W?p�������A�=���gNL=���>�vz=���2���N��L0?O?�ٿ�ۀ���}(>qt���=,?� ?��m<钬>�%?+�+�E�sZ>ˀ3>$��>��>�>@����ڽ=?�T?�H�񮝾ȁ>?뽾��y��^=�D>v�7����\>���<8���j�Uِ�h��<a�M?-n�=4b5��}� uܾ�<� �>Y�T?�kg>(��>��f?\.?�8:��⻾6�7�0m�H��<�N?��^?Qc�>vun�����e�)�b?��?7�> Z�{׾��4��{W�;U?�a�?��8?lM>��f�	����B���|?�t?�����l��1�J�r�>��?R��>�'c>�<��n�>�b>J��>�i��\��&L���?���?���?�
����<AZ� v�>��?�)>�����A��踄��H�=3��>)�ľ{1	�d�����<���>|/>?�O�>�r����C޲=cb��鲵?ۆ?�|���7=dH���j�����\���>��Ǽ�>� �ᾗ�����N'	��S¾�u�1�>�@�>*�o��>� g�� ޿�п.u��Ǿꮾ��?
��>���Ǻ�0������ŏK�Ί4��$3��R�>��>e���?����%|��;�f`����>���Eԉ>6�O��ȶ�l)��oK.<��>��>?��>U۬�/������?t���O�Ϳ�f���g���X?>�?�,�?�?P<I�w�4!{������F?�Ts?ƊY?�%�'�[�>�1�U�j?g���6�_�U�4��D�R�W>%3?/,�>��.��l=�>��>H�>).�ĿEz������d�?:1�?�����>��?+?�;��������')��<t���@?�O5>����8"�K�=�i�����
?T�0?������,�_?�a���p���-��ƽ�ڡ> �0��o\�>F��g��/Ye�Y��mFy���?�^�?�?H��) #��3%?J�>6����3ǾB��<�{�>s#�>4N>e_�)�u>y�P�:�ec	>?��?9|�?k?ܒ�������J>k�}? �>Ln�?L��=fW�>h��=����穴��(>�=>K:P�X?A�M?\3�>r��=C<�rw/�e�F�a�R���R'C��>�_?7N?p�b>�3��	�'�/�!��%ʽ�K7��ݵ?��]���׽�%7> �>>3<>�E��׾ V?���\ֿ�n��'Ⓘlh$?`��>���>$����v�	i=m�J?<��>�I��v������T�V��?�V�?/�?Q��!������=5�>��>��E����X�W�>H�K?���><����}��,�>�.�?#�@H÷?�e�hI?SS��t܍�����cE�D��\[8>�f	?�9��(i�>��?No@�Zl�p��愄�:��>�ۧ?ƞ�?G7�>+jw?���m�0��)>$*0?[?v?���>`����0��>�8�><�R��w��Ds)�Q�h?�@��@n?�4�����Y3����;}*��s=Yޠ=�(#>~����> �����=�zŽ,&=}j�>�:�>uIv>��$>d�>�y/>�����z��2���[����9�%������qy��(�V�Y�f����n��W�
�XR2<�E���hd�,-�u	�������_?!�w?�Q�?�?����C=D�Ծ���<_΋���==;>��.?	m?DZ8?��W�fFʾ��}�u��4���y�e����>h�1>^q�>%?�>C�>Iw�=���=��>��>�o�=J+i>���=��>��1>��>���>��^>*<>ٜ>!˴��/����h��6w�z̽���?�}��e�J�1��&;��͝��LI�=Z.?�l>j��=п��`3H?9���n.�F�+�	�>��0?q]W?Λ>z��0U��=>�����j��i>Aj ���l��)�D&Q>�p?�f>�"u>��3��f8���P�h����f|>�26?�඾�R9�\�u�k�H�-Vݾ�+M>x��>,mD�jh�����]�Ri��{=;m:?�?�t��4���[�u��3��1?R>t \>^,=l9�=�4M>��b�Zǽ%H���-=��=��^>v�?w0*>�A�b'�>X�k������E�>X��>���<��h?��5?`���nO�z����1��İ>Y�?���>�k<�ƽ��@����>�"�>�=M-�=�gy��貾�u5>�EV�e���(�C��9�<vd����p>3z>?���M@����<��~?@~��㈿��V���pD?�,?J�=(�E<D�"�{���$=��4�?9�@=j�?;�	���V���?+B�?���H��=fy�>Fӫ>�ξ��L�
�? ƽq����	��0#�xO�?��?��/��ȋ�l��$>�X%?��Ӿ�k�>����Q��T���9z�bX�<��>^(F?���G�c�ŀ8���?�?���|���dȿ�v��Q�>I��?� �?P�l�z�����?����>��?��X?4�`>^o־v�L�?��>��=?/1N?6m�>�j���BJ?:ɸ?G�?n��=rܩ?J'�?��e;�|u>m��N�Y��9�?E�����>G�	>�1���R���Cp��������I1�����>��<��>`)1��nݾ�;_=��=������=���>��>|�g>x�>Y
'??�N<\����Q;�4߾��*�I�K?���?����1n�V8�<S��=��^��)?�M4?һ[�+�Ͼ?ר>޺\?5À?�[?Db�>#��U<���翿�}��Ԗ�<��K>�0�>YE�>����RK>g�Ծ�5D�o�>OΗ>���Aھ:.���򢻏@�>�d!?��>~�=ā ?|�#?_�i>@�>}vE��G����E�X�>sL�>??�	?8�?|���I3�'����Ρ�!_[�|qN>��x?�P?�r�>�~��1e����B�H�wT����?��g?�}�4�?z�?bu??9�A?�-f>����׾���@�>��!?��� oA�E&����o?�C?���>�ꔽ�^ѽ,7��>�Y���=�?�m\?��&?���`���¾^C�<_"�9.��m�;�]W���>�&>������=��>;��=�
n��m6�n�Y<�T�=��>�m�=��7�����WC"?�?�;PF�� ���
y��1��!�>�o�> �	�ńo?Ë�=,�@�2'������jբ���~?ᓹ?S֌?0��Ek��wR?>�D?�?.�>��#����c������-W�s�F��W�d�>��=D~ξQ������Ŋ���\���Q�6i?���>��?�?	?��C>P=�>�����X(����$�ﾥrs��#��S@���}���_���b�'�gξ�����'�>'o����>f�?M��> f�>*)�>��R�'?�>|�1>7��>�C�>�h>�8>���=�:�Sֽ�R?�LľN� ��?��Z���	�E?e]?�4�>i}e�}Ճ��r��t?ٍ�?.��?.f>��h�(�2����>w??��v�PJ?�[^=�<�2�6��+gԽ:��<K.��Z�}>_�Լ��9P�*ͬ�b<	?;~	?���=���SB���c��?a1>���?�#-?9��S�J�����I�+�=����9ӽ���߀6�'{_��v�*�w�C�u��&�7�<�?�?��B��~
�<�B��q�{�x�M��>ɛ ?��=5��>���=�|��U.:�m�o��)����51?�_�?�b�>�rJ?��<?�M?�J?��>��>_Ц�^< ?�}�:~.�><�>r�9?y'0?N1?�?��*?��f>}�������׾�%?��?d?��?��?�T��"8ǽ���~p���z�mv����o=B��<Sx׽�n�2gs=�RZ>�s0?Qf��Z�)�+o߾6�>׳X?���>�z�4oY���_�ؓ�R��>��q?��-?W����9[n�lb��R�?Q�*�8W�;��=1�<����<ѽ|虻�?9=�n�3�� �3K̽�`[�05={�Ƚ�y<Ա��4z��3Vs����>?�rt>i�l>Ց�"���i!�i��=�9(>��g>��@>��ǾD�������h��Ux>�T�?��?�zF=�l�=ܮ>�������`K��\Ҿ�L6<�?)�?�S?
��?��-?	�?��>����������7��G'?m!,?��>�����ʾ��ۉ3�ܝ?s[?�<a���c;)�Đ¾|�Խ��>�[/�U/~����"D�0ꅻ�������?濝?�A�c�6�y������[��Z�C?�!�>�X�>G�>=�)�U�g�s%�\1;>��>TR?gv�>BT?�~?�P^?�)W>E?�dR��5ɘ���<��>��A?��?�y�?� �?g!�>��>��$���辡w�#�ϼ�T��V��_�\�Z%?>a�>�>���>�B#>F�Խm���B�>�'G=G�q>��>�>���>�i�>�;�<KtD?���>-�ƾA$��(��#g��R�
=V<�?��?5&H?�( >��?�E�l��y4�>*F�?�@�?Q(?n~�w�>K�����x�����^�>���>��>�Z���$�<��@>��>��>7��� ����~=>�?��,?6}<��ſ?oq�(tq��뗾=UH<�����[d�!����#[��X�=�;�� p�
����\������u��p����z��k�{���>h��=i��=
b�=���<h̼NV�<GbL=i�<j=�vr��Re<��7���˻K��Q�D��T<I=X<�Kپ_ �?�F?�{3?��G?�	l>k5?>������>�����?iݚ=��Aվ� ������@���y꾣��X�n�	믾_�>˧6��C%>?�'>pG�={��=�K>^�<=Ԥ�=5��<I0Q=˥�=���=�}�=�M�=NI>�%>5�t?g�GȀ�kp��u=S5?��z>B4=�{��xc?x��=u�������-
	�E܎?[ �?H��?�(�>&6��A�^>s���fE����-����=ov>�{��v&�>�d>��"��6����o��А?�v@8�D?$���:���'7r>�:>��>r�W�k�*�;���M!��#2�BS1?��A�qg���9�>7q�<4F��*Ǿ:0ȼa�>���=0Uֽ�~K�%��=$Z���߀<B�=w$Z>m�>V_W=��a�l�a>��=���=��=������<;x��RP��m�=���>FSU>��>�}?�0?4�c?���>]�p�\о�'���3�>���=ڱ>C�=F>���>_%8?�D?��K?]̱><z�==��>�y�>��,�a(n�>~�e���6�<��?�ц?��>DK<XTC�P$�+%>���ý6+?�51?kY	?qk�>����Iֿ�r�ZjJ��%Ƚ�\4>f>? �Iǽ�H!=�H�K���=o��>q��>��}>Y�=`�>��>��> �q=C�S=��>5N^�zps=�x�=P�[�:�����=��/�9p< �r>1�%��\��aG<���� ���s�@<��l=�3?��a>���>��=H(���o5>V2��Z`R���
>򯟾S�R�i�l�|"w�O���>�xY5>vr�=���5���(?~,�=/�>ޟ�?��s?�|�>�'@�a)��꛿y��~6��̎�=�Ч���u��D�~�_�/�G�����>�ߎ>��>k�l>3,�`"?�eDx=��� n5��>�V����t<��3q��=��p��i�
�̺|�D?D��`��="~?�I?�ُ?�f�>�Y���jؾC0>C���y=u�iIq�N����?x'?��>C�;D��þ�2���K�>�w�gp�+����^ �����\���\H�>1���z۾��%�T1����1�E�� ��C��>��K?>˭?�r�*兿.eM��U���<��?��O?x�>�7?�r?GVݽ@= ��򹾠U=��o?)��?���?
� >��=D=׽wu�>�]	?�ו?D��?Zqq?��D����>ч<�C>z���=���=��p=�'�=�x?��?x�?�����q>辀7��J�m��@D=&I�=�؏>s@�>�c>�j�=�bS=�Ǭ=�)\>;Р>���>]�T>{K�>(I�>�Qƾ/\���1C?��>�>�>p ?K|>�K��>��B�=K�<����|䰾AV"����=�=>"r=����B�<�ҙ�>�xп�d�?T�>;��vo?x�'��N�o�=L �=d\�<`L?G��=8��>�]�>�G�>w�=�3F>�Nx>��ݾ�I>�l��L#�柄��o|����z֊>����]���|I��&4��*�Ϥ��R���Xd���w���?��]����?: ��O������������>�>(7?���������ޖ>
�>�]'>�d��հ�S@��_����?w&�?z�b>)n�>��W?��?�!1�_�3���Z�Lxu���@��7e�jr`��э�񚁿�
�|#��o|_?]�x?pNA?�B�<`5z>���?2/&�u=�����>\/��o;�]�?=_��>bm��Ca�ӒӾ�4þzq�e�E>bWo?d��?��?��T��As��/>`D;?ؔ/?��q?��/?��9?8c�*�(?�->vj?d�?��5?|�0?�%?��/>���=�U���(=����犾�*ս=�ν�����>=���=P6�;�%�;��=���<�Q�n��iӺ������<��<=�D�=w��=�Ȧ>�]?��>��>m�7?c����7�!?��j�/?� ;=����ĉ�������->*�j?u�? vZ?V]a>��A�"�B�r�>�(�>OD$>�]>Sv�>e�(F����=�$>��>�Z�=� M��ـ�!t	��W��W��<_� >N�>���>C�=|6/>)��|^��DD>b��C�F��Q���?�h#N��	о��>C]?�4?@��=����Sq���4���oM?:sB?�{W?2�~?��=�Ӿ�9��v��m�D��>A>�^���'���T��]U��	g��~�#>v�+̜���r>9U����%�z��X���־$z�=>~�A(<�x�=3̾��g���>�'>��ϾI!��Ɣ�$M��q�Q?(��=PQ��-����/ؾ�~�=E	�>L��>]��W�71<�O���od�=���>�2>�;F�S���L\A��~����r>��N?Xg?�ܒ?��v�����8����c���95߽X�?�'�>I��>A�=��(=�}̾�����]���'���>P$�>��i@��a��w� �4����>��?��>�%-?�2O?�#?~�^?��"?���>n>[����H���L&?y��?a_�=��׽2�T���8�pF�5 �>*?��?��_�>��?ѓ?��'?��Q?�_?��	>=M�J#A��.�>��>H�V���*_>�FJ?B?�>��X?���?�w=>]�5��H��>��$��==�!>d%3?F#?Kz?
��>�|�>����_�=C��>Qc?�-�?��o?��=� ?��2>)��>�1�=���>�{�>8?�UO?��s?��J?sv�>,ߍ<C쬽����/:r�C�M����;�H<��x=�{�ruu��p�\��<n@�;����S����q� �C�î��g��;�`�>��s>�����0>o�ľ�:��_�@>�*���Q��Oۊ�ς:��ѷ=���>}�?y��>7]#���=|��>H�>����3(?��?�?�;ٟb��۾�K���>�B?ա�=L�l������u�h=��m?��^?�lW��#��s�R?&1q?����ty3��>Ǿ@����>'��&?��?�Js=�ˋ>��?x�?�*? A�w�\�������e�4�}���+>���>q3��t��>\�%?�5�>�*�<���=nv��������O!%?E=�?ᜱ?��?�
�=��u�����y������}`?���>�E���S+?!+޼�?߾��%������]}��_Բ�wN��� ���F�
օ���ҽ O�=�?B�r?'�q?uA^? M�m�f��:c�wNz�]�H��� ����E���@��zF��&j��I�h���炾L �=�#k�>�2�dn�?l[/?cR�8�?����V?��|���^�=�z�����;�m���amB=�ԑ=��k��U.�-�����?���>�X�>MV.?/�m�-�7�,CN���$��m��z6>��>zz>��>P���TL*����о���|��<I�V>�d?'#S?�P?�97��V2�)�s��P)�(�p=�x��/>?C>9nW>���c��e�z�:��In��{�U���@�*Ƌ=&lF?W��>^�a>�'�?�?�9�hlھ���Ay5�.=��t�>��[?7��>@>�� �y�K:�>Z=l?�`?'�>⾃�%�=Ă�����-?��>���>h<�>jJ���b��&��ظt���2�TC�=��e? ����C��n�=D;c?ծ�<�iS��]?o��<��/�&������m�=�9�>��n>��=Hs��1�-����Td�!�(?��?^����?*��R{>p�?��>�4�>��?[ӟ>��ƾ��v;S2?��]?~�I?�.B?�`�>�=�z��K�ҽ<�(�ƅ2=!��>fe>�iy=���=�z�+�f���&��-c=n��=����Ƚ��f:9мY��<J�$=;@>s�ڿJL� G�~1�2]�)��`��v�P��V����t��ɾ������׽��P<ni��G�9�-��k��z�?��?"`5��˾0���酿(��\T%?U��3���o����}<t��ǲ������D2��18���P�WtV�"�&?�<��w�ǿ&����ᾄ>?��?��y?����"�q8���!>���<�?��\F�֚��dο4�����]?V��>@��ڎ�����>f΃>GQ`>F�j>�Ɔ�Mx��)��<K	?��,?���>�t�}�ɿW��M
�<���?�@|�A?� )�%x��XQ=���>�	?2�?>5�.��s�p������>��?Z��?�\?=(<X�.��	f?9	B<Z;F��*ۻ���=�6�=��	=��@�K>�*�>��2�C�P�ڽ/2>A�>Q�!��5�J_����<�]>�pٽ����]��?��R� �W�d� ��By���=��j?'�>��=�A2?��8�E<ҿm�`�QBX?���?b�?�<?����m:Z>�羇R?�@??M�>��0�"�n��	7>�}M���)����-g�0�=?��>ށ>�U0�}��O��������>J)��wȿ�N"���k=6���u������<̽yF�����Hӄ��s�9��=���=�aH>C�u>YI>q	i>�T?6�i?�;�>��>��ǽ}��r,̾�錼�f�(�ܦ���t&�{������H�L������O��u˾*9�� �=�*l��:���],�	0}� T+��5:?��Q>���ѢI��t<'����y��Xp=��5�Hž�+�	f�tK�?n`?q���D� �!6��M��0=μk?n�#��u���C���6>F��=`��=�e�>�6�h� �y�.��L\�}F0?��?'o������@*>X�!
=lr+?{�?ـ<�j�>ځ%?�(����:Y\>k6>?t�>_	�>�W>y���
ܽ،?L�T?^�������p�>�}���#���R=q�>�V/��R�K�Z>Њ<�2����U��e�����<TG?�Z>�=��6�����Ƈh>>-+>u�?ؓ��?��?tS?q�A>�.��2��`0`�oR�=�r#?`�z?oM�=�j
��Ӳ����T�-?��*?��>�wt<5�b��.E��Շ��63?L_?�U?Ri >@Kn��ﰿ���%T-?�5o?��{�4���F
¾g�)>P��>�V�=zh5?w�)�r����~?L߹:C8����ƿ��C���?�f@���?���2����>���>n�>���A���]Q�=d��ҏ��[�>n�Y���7�=�̾+0:�!?�,?xq�>�z������m�=����wZ�?��?'ª���<���Ml����! �<s��=����w%�����7�5�ƾ;�
�����������>OF@=U潃;�>�O9��+�RYϿ(�sϾx	q� �?O�>=^ȽP	��n�j�nu�Z�G�nQH�I鋾�M�>�>㳔�J���A�{��q;�|#����>��
�>M�S�U&������8�5<@�>\��>O��>~*��f罾,ř?�c���?οF���ڝ�{�X?,h�?�n�?�p?�9<��v�A�{��{�U.G?�s?Z?r%��=]���7��j?�_��U`�q�4�rFE��U>�!3?�C�>�-�&�|=� >��>qg>�#/�2�Ŀ�ض� �����?]��? n�s��>À�?�s+?i��6��n]���*��Y-�<A?2>Ս��+�!��0=��Β���
?�}0?Bx�.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?<�>��?ۄ�=�d�>�=��9C-��u#>,�=�B?���?2�M?KA�>mc�=��8�b/��ZF��DR����C�)	�>��a?��L?��b>5ܸ��:2��!�q�ͽ�61��B��@�9�,�6�[�4>]�=>0�>CxD��Ҿ�;+?]�,���
��.�=bVV?��>_"?�^��=˽7?�>ȤO?[��>G�����Ǉ��%~=���?���?��?""%���<!V>>I*�>hp}>����DX��7�r�ׇ>=�>_�@��䟿����F�>���?(@q�?��W��[?�����(�w��7����n�ż�YJ?����Yu�=�H??J�=Ƿs��"���/y��Q�>��?C\�?�?��U?��l�I�ފ>�r�>է??�X�>G��=6/þ�+�� ��>Z��Nu������}z?�]@�Q@�j�?�&��t�п�\�Ӿ�9@����=3� �Қ�>���f���zR����=�=��C=��f>��$���=��>�u�=u��><R�� B&�¿������/��/�����ȁ���5��#��v¾$� ��n
�d$�����dd(�3�n�cj�=�nS?4V?��n?p�?v�<��y9>�����a=]��2=� �>�H1?A�L?�(,?�=咚�G�b�d�}�����*��.3�>J\>��>ɝ�>�=�>SO�K�(>�:>��>��>S=�������<�J>J��>FA�>�%�>��4>��+>V���1����u����Z���!�?bI��\gM�pt��O���'���%�=��/?x�=2J��.n̿�R����L?P��D��ɽ�G�=z&?"�P?�!>eo��@3�_O>�O����T�!7�=F��^����^)�M
M>�&?ɦ�>F�>��'�B�%�&�p��&��B[�>w	A?yTվ��[��J�g$d��"\�J�>T��>�*]��G/�S��J*��Q;t���>4/?��?�M)�������d�y�#���H>B�=�=g��Kh>��=Ik���6��49�7~�=_ >�>�Y?��+>�`�=�ͣ>�i��zP�x�>�B>^�+>�@?E(%?���~�K����.��v>�g�>"�>0i>YJ��h�=Vc�>��a>������{���?�9AW>��|��z_��%u�.�y=�ї����=�|�=�� ��'=�HS&=�~?���(䈿��#e���lD?S+?i �=�F<��"�E ���H��F�?r�@m�?��	��V�=�?�@�?!��Q��=}�>
׫>�ξ �L��?��Ž4Ǣ�ʔ	�/)#�jS�?��?��/�Zʋ�<l�6>�^%?��Ӿ���>UԼ`Ԏ�SWm��_��=x��>.[?��ᾇ��aq>%(?�o?Ƌ���-��͓ʿ�>X���>H�?ӻ�?h��8Y���zo�)J?)��?��!?0P�>���� ����>��?N�O?j��>��R��9��B?p$�?��?�HF>2z�?lFt?6��>9O����0��²�Ѧ���X�= Q ��L�>Z]>�[��<+F��-�����j�j�� �[Sc>��5=�8�>��dN��{��=��������(W�>�r>BeU>���>4� ?/��>�S�>���<V���L�z�8����^B?Ov�?$�q�]��O��X���&��>���?�y>�(�/�=�V�?�@�?�}?�|�>�$�EU���ĿPv��\�?��s->9)�>���>[a�p��>�S(��V=R":>![~>ۭ�=�G���ﾊgc�0|�>1T3?<U?kr>�V?U]7?�T�>��>��;�:G��MR��K�>8y�>��?F(�?��*?-������sK�����)�\��	>~�x?0�'?��z>�ߘ��%�����\�=k�g�p)p?�sa?d0>�?���?��n?a�W?v�>Zl� o��+G�M��>��#?�G��.�ڻ?������?�?08?
B���l���)�=��g�|K��4&?�k?�=�>}�K��)�������=e��=uG�=�>H�^�.��������=o|:>�������@
����=���=9��>aa>^d��=���s)?y�*�����(=e�Q��e%�2�>�]=��r�Z?.c3�4�|�wޟ�A���lv�[��?s��?k�?D���^f�l?f?'?���>躌��l�X�ᾟ�F1����@� >/��>�߽ )��̮�z������@��:�S"�:# ?�k�>i�$?�?%�%>��>�-Ӿ�/��k��u�R��` �ls:�}�&�����&���.��?����1:��\��>=�h��/�>�E)?z�H>�A�=)��>�T��u��>�2i>�V>1��>��Z>��$>�>����3��K�L?ʳ����4�V����V�a�K?��{?�?�n�����B𖾵�$?S7�?�W�?�q>�5��^�L���> �"?�Yg���?1m=�Y\�LV<����r��	b��d峼j�>WMM��?k�߼(�����/?6�1?
n$��p��P��b\��Th�=�U�?q�+?�K)��R�v�m�8V��P�r�?�	�g������_$�ʧo��(���郿���(���3=��)?�d�?���N�9۩���j��a?�hNq>�u�>�ߗ>Γ�>b&K><��K(0��6[�C�'�����u��>b�z?.��>� _?O�:?).?u\?��b>�D�>JE��@�"?H'-=HJ�=S�?:�??��7?�+5?
�"?�?��	>6���N�����j�6?�	0?��<?x��>s�-?�!������f�;G ͽ(Ug��F>{I=���5y>�!<�!Dd>X?`~�� :����Es>U:?#E�>���>bO��i����ę=�l�>�?��>���íz������>��?�!߼8>;=�� >z��=��p<r��:*�=���=yN���ە��U����=��=8i�=��(=[U%����/鯻+��>�7!?��?��>A��S-׾`�v�*4���>�@$>���=]a�i��ҙ��B����>��r?��?0�6=#��==�>����_׾���}�!.����?n�9?�ja?�3�?,�{?Z�g?|�>0�c̓�����}���^?y�#?�ǭ>�<�����|��2M�\y?�5?SjT�l�O�$�F�������a>�x�i�o�����	O���"������̂�?��?�@=��L�+Y��}[���s���H0?�6�>5��>�Ƕ>T�D�b�{�����>��?żU?kW�>�P?�{?;[?��S>&�8�=-��󴙿����">��??'��?��??sy?D��>w>z�*�c��~A��2�"��p���V=��Y>���>���>�é>��=��ǽ褲��A�2O�=ćc>W�>��>���>��v>i�<��G?�`�>X澾���ʤ��׃�aB�eu?�ː?N�+?e='A�v\E�@����v�>qf�?ë?��)?Z�T�Y��=U)ۼ���ޓp�ۉ�>�ɹ>�љ>_-�=��A=qe>�U�>���>v����ɗ8�'hM��
?&IF?�}�=�wο�A����}�25}�.�Y=�v���h��.�������ݻIV���'=�x���UY�A�������1��������i]�
��>�=ۗ&>�t=��O=�һĐ�;t�=���<��<u��Ij<3����a��Ʌ��m���̥���=���ˇ˾��}?5FI?�+?�C?��y>e>$\4����>1ǁ�60?P#V>{2P�j��o[;��������G�ؾ7o׾��c�R˟�J>dI�ۭ>L3>&+�=��<`��=��r=`��=�S�m�=D�=�L�=�^�=���=|�>�M>�{w?6dm��	��@y� r�<�)?dK�>��'>����+|-?Y�>>���wߵ�/�f2�?���?�n�?�R+?G�־^fm>v5L����<F��뵖�s۽x��>�d��W�>��>���y����"����?5*�?�BL?' k��пwd�=�a:>)!>5R��G1�;�a�М`�uyX�I�!?�p;�܇̾v��>	ã=��ܾ�¾��?=�H4>�}I=D� ���]���=Qnp�[�6=�Qs=⃈>K�B>"��=�=��3��=(�X=��=<HP>&���),-��,� n6=L�=qp_>0:&>���>��?yl0?qZd?��>�m�-Ͼcm���J�>ؤ�=�#�>�t�=�B>3g�>��7?4�D?l�K?��>�o�=}�>^�>�,�t�m����{ӧ���<���?>ӆ?4ϸ>f�R<�{A����xl>�<Ž�g?�A1?�u?��>zc�S��g���m��!�>A����t�g�Ҿ�}���ֶ��
6(�7�#�I(<>��>��>��D=���=��><��>P">��J>%n�X��	C�=�#�)��=��<>|��>�<ײ����=�	@=�jV>NU�=գ�=�f��lb<���=!��>��:>̟?=m>��־X�>��Ͼ�P�?<�=Z����G��-f�Ed���%��)�|�7>��L>O{q��%���?��w>�
�>�T�?q�d?��;C㐾(���u��-r��BI���<=�f>��F�F��h�xV����C��>5�>��>0�l>,�R$?�j�w=�x`5���>�{����!)��8q��?��m���'i�)KԺE�D?F��ݜ�=� ~?p�I?��?���>m��$�ؾ�30>�H����=;�h,q�qp��@�?'?e��>�쾴�D�-H̾p���޷>?I�
�O���.�0�_���̷�叱>������о2$3��g��������B��Mr���>'�O?y�?�:b��W��
UO�+���#���q?�|g?��>
K?%A?5$��y�r��nu�=a�n?���?d=�?�>�Ž=����9�>{(	?��?���?��s?u?��g�>�A�;�� >�|����=��>�M�=���=�m?+�
?��
?w-����	�������]�H��<̟�=<z�>�Y�>}�r>���=�Bg=sV�=��[>z˞>��>`5e>^�>F�>6D������,?Z!�>��>2'L?�>�P�ʲ?��<��>2�;W������(�ߧ����=XE�<�#%;;�D�b>�>�˿���?�z�=7�8��(L?HW� �(���>�v>D�=3��>9&>#zy>L�>aPZ>|��=�>�A�>�~��:��>B��O�F�j��a�������>Wu�˔j���ݾt�= (�N��(�ᾒ�s�x2|�d#0�b�=&��?ncK�=�7�4V��q=՚-?h�5>^O?����w��=�O�>� ?V��>ʝ�n���Bŉ����G͛?�h�?�D>T�>���?1K^?]��Y꿽,m�=���G�W�m�$���R��ڽ���g:��q���k?��\?ۻS?�M[=9x>c�T?�8̾�2q�PX�>sG\��v<��(>��>Z��xQ���������K�M�<>�_?�P�?�G2?J+#�Z4���^>`�?pU,?�?��%?:�b?sM�@�O?IU?�Ɯ<��?�i/?�j8?V�
?Q��>��K�D�����ɼ.ڽ�����kw=��@;nʹ�&�;=��= W@����<<�G>�yp=H����ʬ�9�S��;����<2h=呍=0��>��]?I��>TȆ>2n7?���}8�X���/?��:=5��vV��n㢾���D�>fk?���?uZ?��a>j>B�~�B�Nq>��>Ӄ(>hC\>�#�>b!��VF�D݄=�|>:>l��=��P�+���	�$���?�<j�>���>�,�>����->#Ķ��[��s>��-�C~��OgX�S�G�]W-�2Oh�G��>�G?��? �W=���>�ý�@i�zP)?��>?�P?vt�?�!`;@$���;��>���3�)��>%u�=�l�a����p���<�b漌M�>�%��_᰾�5�>H���R��-���In���ھ��'>PG�.����@�����;�S���>w�>?�þ"&��ߗ�u���#FQ?ך>l��K����پ�i	=��/>��>]J��"���=;�
4�����=���>в�=�ý�0�:��4�C��>�QF?�h^?R?L��7�v��A�_��ڗ��HE׼^�?���>m ?��:>ᮝ=: ������b�pD�,��>�(�>����I��#������"�ƌ>p?Z2>�
?0�S?;�
?��_?�(?X� ?�h�>S��f˷�S8&?���?�=l�սX�T���8�*F���>ˌ)?e�B�ic�>~?��?��&?��Q?��?�@>�� ��Y@� ��>O?�>��W��L���`>�J?�ó>m:Y?�҃?�>>6�5�񢾝Ѫ�|t�=oO>F�2?�<#?��?Z��>�j�>���&�=��>57c?0�?Z�o?��=��?��2>���>zі=���>_��>��?*1O?`�s?��J?�p�>$��<�,��Q���:s�7�F���;��J<��z=���lv��,����<�\�;󂸼�|�?U�liE�G��0��;O<�>�Am>���f�>U!�)W�� ,=�E�=�����Z�W�M��xy>tg>E��>ê#>�����=�"�>��?X5��?�9?E�D?]��].Z�79�tc�����>+�1?_��񁄿�A���{v���
>g�~?�Ay?"���/׾ :D?Z�w?�D?�h�]�o��n<��q�4�Y�?�A�>��ŽQW�>�5�?I΋?<?����hx���)�]�On־��>=^��>x r�V_M��XK>At:?�Ο>�s >��*=���È�����V.?jVn?�x�?[��?���=p9{�>�տn�վ����oe?��?v�;�L>?È =�4�6�4�K������
ľ��;9��X��{���E;���6��\��=��	?�$|?�9�?�Z?�y'���v��J^�4\���P�߄��6@��T��M�V Y�4�a�"��qw��Y�½��\>Зv��A�M�?,�,?��:�� ?艍������8����=~n���� ��?i=��J�7�X=���=�3�S�V�����ſ?(��>hs�>/<?H`��^>�{/�	@@�h���,�5>��>�B�>
��>�����<�i�޽���On������s>��d?�SJ?9Vp?���5��^���!�����V��_
Q>F@>�L�>��a���&��'��>���p����M��Ï��O=e	/?�D�>�j�>��?�#?���Z6���m���/��)�<�+�>Ye?uU�>�w>-#ν� �iľ>x�~?#��>��?>Ͼ<@C�Y�����y�]z?~5�=?��>^�y�8�j�����ڀ�>,��%�= �`?�E��%9y�K?�Q�(?�y�=@9��\?��>4�M��R־��'�">��?R�,>٤	>���:A!��${�_f���B)?p?"���*�*��'~>��!?C^�>.�>S5�?�,�>|�þ:�.���?��^?�AJ?�<A?8��>��=|��o:Ƚ��&�F�,=\��>z
[>/�l=�H�=_���
\�o-���D=�s�=1�Ӽ�W����	<6/��92U<�"�<	4>n�ٿ�15����)F�-x�&�^�����;�NսA��~��
g��C�Y�V��3�.;6�<�d 
�������J���?���?E��wȞ��`��5����۾� ?�bƼ���"���8gE��[����������%���w��6���ZG?Zm�J˿렿<
���,?m>?p#�?r� ��{>�ǻ�X.a>�O�=�}=Q��������cȿ0y^��q?l�>I�� �>��>���>��>]�F>�o��.X����=��?��*?��>=�-�6�ÿK"��)o�<��?��@EuA?�(����ԽT=���>k�	?�?>ͦ0�Rs�|������>"�?�Ê?�UH=�W�vw��e?��<��F��ۻw��=�#�=�C=���K>�6�>���XB��ܽ"m5>�	�>M`��<��?_�8Y�<�\>^�սKj���}�?��R�<�H��$��bo�1�`>%�}?��>�_5>�?��x���ʿ�5�V��?Q�@2�?$��>����>Q,߾��7?��R?^U�>?�;��l�LgV>���2���Qľ��b��u?><�?��`=8�ɽ��'����t�<v�=C��>ƿ]9��&��;=$C<��	����&���鎽�B��@u�
���"�=r��=�i[>Ԙ>�=j>���>v]?�y?�J�>�=�=�r'�������dr=^@�Y�o��ᨾ��0�=��JU���7澅l�Cx�;���U־?�@��M�=c�R�>ɒ��.��p���9�)�4?\X4>�E׾� N�gJ3����-����~&;g�ƽ9�Ӿe�5�ܾx�=�?%WN?�e��s�=������L����b?'�5��9�������o=��<��=��>EHL=ߓ��i8�� b��J0?f5?�c��������(>�� �T�=m�+?�?��d<v��>@�%?lo)���{�Y>�r1>ѡ�>�2�>x
>>���bڽ	�?9�T?�T��L���9�>�h���kx��y^=�A>��4�����-�Z>��<�c��xF��H���A�<�O?���>ϯ/�`��
�����=�B�UV?��?>m�>��h?r�*?��E��7Dd��J���=Ѵf?�^?s��=U�=�yľ'QξY
?R�D?��$>ҁ��*��,�w��f&�>���?��?b��Ӧ��K���Uy(�*�=?7�f?DmP��A���վ��<�|>�`G>6%?QK��">�\'?�'C��٩�qOÿ�>��?�� @��?6�$��MV��ִ���>�>nMj�y�ʾϺ��+�)<��μ��%?�ھ��*�n��H�-hk?OG?:6?A�������=�\���Q�?5�?᫾.�<����l����8ˁ<g��=om&���,�]x7��ž�
��v��:$��yن>�>@t��7>�>w;��*�9Ͽ�����Ͼ�l�h?.y�>h+̽ाǍj�C�t���F�mKG�3����w�>.Z>�۔�	����{�F;�(4�����>Iw	��Ո>2�S��Z�����,�!<���>��>/>�>���Q-����?ۇ���4οĭ���:�H�X?�L�?�k�?;F?�,<�v���{�*��?)G?��s?F(Z?�'��\�۩<�u%W?���"�X�B�VZ�n�T>�p*?z9�>�+@�jJk>�>�>0�?���>�����������.ܾN��?�}�?��DS�>B�?7?�c�|]��M��F������=4S�>4K�<èW� )���O��}3�@N?6�+?��L�u�xm?-K�U$S�����c���I�> �< ]�\6=�`��7q��ҩ�����5��?��@���?� ]��^:���?�/�>�k��P��5�W�_3>H��>u��>����2�>��������'>���?�+ @�"?ބ��ۨ���ἇ��?s�>��?��=�D�>�f�=�᰾A:&���!>Q��=~4�`�?4N?���>�'�=?�9�ψ.�0#E�F�Q���eEC�A��>��b?*�M?�_>�V���,�j`!��(Ƚ��3�nJ��=��6/��S�X�8>��?>b?>QAD���о��?ڷ����<��__ƽ��.?���<��?�m�ʾ��+��>��O?Ui>��ؾ�`��W���1�1��o�?E��?G�?�lپ	�8=�Mm>�~�>��6>�'Ͻ�������g>�s?�F���'����r����=���?A6@#�?�;M��?8�ھ �t��1������&Mi���?Ԙ��Q>��>CX��t��2���-�n��T�><�?�h�?ޱ�>��_?��n����z)�=��!?[�P?��?x�=�q�
4M�[.�>E�0�������&��ES?$}@��@<�?�/��H���%��A#���ܮ�y�;��=4|>��8ҋ=��6�7�˽HN&;�0A>k��>�.L>�,�>�d>�.s>� c>�ć��k&������榿�m6�����q�㨠�	����P��Ǡ�ڿ��橾����5��R5��G�罳T���T��=�RZ?fT[?o�W?=[?�$��� G>�����> ;���ө<X�>��0?��:?x�?��=Z��a������c��L.�����>P2�>)q�>�c�>���>��Ͻ`*>
/>Ra�>շ/>u�>=UN*�}^����G>u�>��>5+�>��6>$.>E1��X��a�j�e:����нJ"�?�����(K��H���Z��������=g-?��=�ޑ���Ͽd���wH?�^��r4�M(�+�>�)/?|�S?�>i:����_��V>����e�>(�=/j�z,t� �(���R>z�?��S>%�>�|3�=�:��Y���̾ώm>VH:?`��� M�7�w���L���Ӿ�4Y>�O�>�Ǽ� �}D���@����N���=R:?ޙ?�4ѽ���#N���X��wg7>�yM>��=�2�=n�V>�;��2���Qb�Wu!=���=��i>&B?d+>3��=�p�>�˚��uR��{�>;�G>��)>�??/$?ax�tX��"H��$�,�Z�u>9p�>���>j�>$�J�Hy�=IJ�>�$d><�
�aۇ�����c<�A[>��`Ma�X6x���t=!*��2��=�=����fh=�:%+=P�~?O��Ǎ�����u����kD?*$?���=��a<.y"��\��������?@�?5����V�3�?�!�?�x��?0�=���>^��>�Ͼ��M��?��ɽ�p���$	�)�$��2�?,�?u�;��s���_l�s�>^>%?��Ӿ'�>�_��{ޝ������j�C��<:��>e?�6���v�����?��>Y�Ҿ즛�`v˿�u�Eu�>�)�?��?X�m�3���Z+��T&?A��?5zQ?�q>܈���m�$��>��Q?r=?`��>A"��oV�;��>l�?
��?!-E>Ш�?&�k?��>�Ƹ�+VK������򅿔U�=���@�>{�>�mƾ��D�T����抿�j������q>�� =h�>�5Ҿ|��=��0J���A�<��>�>�`>p��>�z�>��>��>�T;�g���|[=��`��5i*?*�?���u�w9=�N����Y�l0�>F�W?���=Ν�X�>��x?<Pm?�(X?�S>d� �"���fE��5����<何t�=$�?V��>GA��1��>/�z����<�m�>�s>��:!��ۀ�u;����>��M?"��>���=� ?p�F?T��>+:�>H�>��ѳ��4���>|'?/m#?��?�H?������!��؊�eۭ�=�b�VfN>��X?�?��Z>��^�ߝƿ�xA=�12>�=s���_?��9?��9>=ı>⨐?y�d?Υ9?��=s���\ھ=BȽ!>(>��!?i���A��L&�*���{?�N?���>�*��6�սN�ּ��(t����?�(\?p?&?.���.a�Eþ�0�<1q#�*XU��<�;g�D�x�>s�>�s��K��=�>�Ұ=�Mm��P6��(g<�b�=�>@�=P27��l��g�(?�L�׍�����=�Y��L��m%= �>�O�SU?\4����f�����z���Fף�g�?�n�?�)�?2�Ƚ�[��H?2|�?Z5%?]b�>� ��s�����^N�|/��QG�pJ���<�>�Ǧ=9ᅾ%̖�h8���U|�y�=�J�:�?�>��?��?{AW>c��>�ȴ�ߚ(�xH�/���]�k�B3�ګ� Z��踾�z�[�D������ύ����>�'�;.*�>
?s�R>x�>���>�k����>�H>��l>�D�>��>�> �=I1'���JR?Y���%�'����䳰��1B?Bmd?�6�>�Ji�m���f����?��?�q�?-&v>Q�h�R,+��m?WG�>���@n
?y:=[H�Y��<PW��Q��KG����w��>?׽W:�2M��sf�:f
?�/?�����̾!)׽�.���$v=�m�?x)*?�%+���P��2o���X�ySQ�L�)���i��Ƥ�`�%��Yp��Z���{��y烿�E(��7=Zb*?�B�?�g�ƻ쾢3����k�u�?�Pcf>@"�>�>���>ɽC>͕	���1�\�]�<�&��G����>��z?�nl>�~O?�V? q??spF?n*>e��>��ƾo<?�@�=��w>a?��5?��?	�?�?�I?��=����-������3?��B?��?[��>���>E�Ҿ?aa���z����=<ٽ*�;=�'�=�*�=�r��k*��
�<)X>�/?��v=��T��� �c�>1�H?��>,��>t�5�B�=q� ?94�>��=?��>�b-��>��>���z�>Q�?�2��j��Wx=Eg��"���|V�q��>�>c}>ۗ>f��=��>�w�>6��>!.3�������=��g��H;=�?`?jW�>��>mま�$ؾ�_=�Eo/���>��>j`>��ɾ]�������#j��F�>��|?�e�?	&>t�=eˮ>��ľ��ھ�����<��(:��T�>r
�>is-?�v�?�q?�?��<SM��ˍ��|����;�?a,?>����ʾ��$y3���?d?�>a�mk�c)�;J¾�8ԽB�>�b/��7~�����D��0t����r�����?���?�#A�a�6��辵���S%���ZC?6��>m�>V��>O�)���g���DP;>�_�>��Q?9Ȼ>�R?0j{?9�W?�qP>68�����mӘ�*졻�� >��<?��?}�?�[x?C��>ܦ> Y3��[�߅�� "���꽈����a=X0Z>�@�>��>B.�>���=����OŽitB��̞=�b>��>��>��>>dn>��</�7?-��>���_������(�þ)ڔ��?��^?��7?�g%�ӓ�S�r�G�"�*��>U��?���?,EV?� ��>-y��b��y������>?f?RI�>���m���+5?=#,7?i�>�զ��r
�p����=�.u>��J?��0��ƿI�q�}�p��ė���d<�����e�g۔�"[����=������[˩�=�[�崠�����.���U�����{����>q{�=o��=$�=�a�<�pɼ�ݽ<c�J=��<�=�p�8;m<R�8�ıϻɫ�����t�\<��I=����ƾ�v?��S?I.?<E?ZWp>/�1>G�ǽvL�>��z&?��>t��;
��\!�ۣ��d#��MT�U�� �d�o����>p+���
>��#>S.�=#�,��)�=�a�=� �=B�����Q="�=���=ѹ=E��=ˣ >��>ֻu?E�a�v/��Or(��W">�X.?G�>Q�1>	'־�O?��T>!���J���J�e	�?�?{�?.
?�I�ή�>�7�"н���Or(��A�>�=>L��Cp�>L�o>=
��s����
>��?!"@�8>?|���+�ؿ��">q:8>k+>�R�{H1�j%\�{�b�S�[���!?W;�=�˾!��>g0�=<�߾NǾ�3.=�m6>�Pk=I���[�Yq�=֫y���;=��k=	G�>��C>���=�٭���=�L=�U�=fO>B�`���4��<,�]�0=V��=�b>�&>6��>l�?2�0?�{d?.K�>�Rn��TϾ%�����>���=S߰>�,�=�yA>n$�>��7?��D?��K?��>���=  �>��>��,�h�m����< �����<:��?
ކ?��>��_<#�?�Yr�Qb>�XEƽZ0?�L1?/�?���>w3�T���O"��p>����<0�/>i��=I��\���z�k��M��S���^>���>�Q�>�݊>ء�>G�>�ʝ>���>l5I>uۏ=��d=4d�=��,<�ֽ�b�<RI�UѼ=�I�=�޹=A0�^tZ<���=���v�\<�	;�=��=S��>�D>-�>@/�=F��-1>�I��-�L�,��=���*MB���c�3�}��o-�� 3���>>��R>����!����?4	Z>�B>
�?-5u?�t>���x�Ӿ	3���?a�S�Q����=��>CkA��+;�r`�>�M��~Ҿ���>iu�>�[�>��V>H�.��;;�; l=��Ҿ2�6�F�>p�v����R����[l����lO���d�'>�j�F?�����=\�?�OO? ǌ?�t�>S�轸־�*G>L����7<S���Sý"�?g(?$n�>�쾠h?�p�ƾH����>Ʊ=��T����2��Y�I
����>����`�ɾd�2���������h_C� oa����>�0S?Q0�?M~^�;�~�P�D��� ӂ�:��>g$^?�q�>h�?{� ?�> �˩���s��� �=��t?�\�?r��?C��=�=>̷�`x�>�}	?��?ᶑ?�s?��@�B}�>E(�;�
!>�a��x��=q*>�%�={6�=�?qB
?��
?�|��ş	��K������\���<~��=��>�m�>mDq>��=p!j=�C�=��[>�,�>1��>( d>���>�+�>�ގ����ؘ&?�p>���>��P?.�>*��v�;��o���,�,����=A�3���<Q��=I;�}En��Dݽ���>�mҿ/S�?x�>4A;��+8?9���Ǖ<B��>mđ��R�<A��>���=��>J>��o> �>�{>�?>WҾ�-�>d(��=4�>st�[H��ڞ�����>Cm���������P�U���ݽy`�� ��A�w�WV}��=����*�?�U9�X׀�b�����=|�F?�oo>v93?�ƾ�;�s�>��"?�'u>w�� ���6�������u�?���?�}>&p�>W�n?��M?FQ�\�C�N�f���mq���p�1Z�DϪ�誆����m���X?s9?�?�>N��>��?'��Fo��ǖA>�WQ�swL��`<>ɂ?8Hc��g���˾�Փ�u�'��BT���=?�~?� R?��-�� ��n�|At?�р?S��?�H2?���?�A!��>�K?�:�>Tl%?m�(?�Z? �>�=R�$�j��H�!��}��~��P�,�6Ca=o�=��=�ƞ=#����jt� �.=�ڽU�ڽT~=���<3�K����=��%>�O>\P�>[�[?�>�>��>?M5?�R&�$�9�W ��-?�T=�h��K䍾:���N���}�>��i?�a�?O�Z?�e>�2A�@���>�>k� >sZ>L��>g߽�8�3ӏ=��>U�>Z~�=;��`��T���|��E
�<|�>�9�>�Br>�Q�=���=Z;=���.���>�Э��/���$x�z����lH�d���
?J��?�n.?���Q����M�;슿z�U?�!?�t:?�1�?�<8@q$� cF�ڏL�"�{��Z�>Sw�<�>+���ſ�n��H/��*�����=!R��_᰾�5�>H���R��-���In���ھ��'>PG�.����@�����;�S���>w�>?�þ"&��ߗ�u���#FQ?ך>l��K����پ�i	=��/>��>]J��"���=;�
4�����=���>в�=�ý�0�:��4�C��>�QF?�h^?R?L��7�v��A�_��ڗ��HE׼^�?���>m ?��:>ᮝ=: ������b�pD�,��>�(�>����I��#������"�ƌ>p?Z2>�
?0�S?;�
?��_?�(?X� ?�h�>S��f˷�S8&?���?�=l�սX�T���8�*F���>ˌ)?e�B�ic�>~?��?��&?��Q?��?�@>�� ��Y@� ��>O?�>��W��L���`>�J?�ó>m:Y?�҃?�>>6�5�񢾝Ѫ�|t�=oO>F�2?�<#?��?Z��>�j�>���&�=��>57c?0�?Z�o?��=��?��2>���>zі=���>_��>��?*1O?`�s?��J?�p�>$��<�,��Q���:s�7�F���;��J<��z=���lv��,����<�\�;󂸼�|�?U�liE�G��0��;O<�>�Am>���f�>U!�)W�� ,=�E�=�����Z�W�M��xy>tg>E��>ê#>�����=�"�>��?X5��?�9?E�D?]��].Z�79�tc�����>+�1?_��񁄿�A���{v���
>g�~?�Ay?"���/׾ :D?Z�w?�D?�h�]�o��n<��q�4�Y�?�A�>��ŽQW�>�5�?I΋?<?����hx���)�]�On־��>=^��>x r�V_M��XK>At:?�Ο>�s >��*=���È�����V.?jVn?�x�?[��?���=p9{�>�տn�վ����oe?��?v�;�L>?È =�4�6�4�K������
ľ��;9��X��{���E;���6��\��=��	?�$|?�9�?�Z?�y'���v��J^�4\���P�߄��6@��T��M�V Y�4�a�"��qw��Y�½��\>Зv��A�M�?,�,?��:�� ?艍������8����=~n���� ��?i=��J�7�X=���=�3�S�V�����ſ?(��>hs�>/<?H`��^>�{/�	@@�h���,�5>��>�B�>
��>�����<�i�޽���On������s>��d?�SJ?9Vp?���5��^���!�����V��_
Q>F@>�L�>��a���&��'��>���p����M��Ï��O=e	/?�D�>�j�>��?�#?���Z6���m���/��)�<�+�>Ye?uU�>�w>-#ν� �iľ>x�~?#��>��?>Ͼ<@C�Y�����y�]z?~5�=?��>^�y�8�j�����ڀ�>,��%�= �`?�E��%9y�K?�Q�(?�y�=@9��\?��>4�M��R־��'�">��?R�,>٤	>���:A!��${�_f���B)?p?"���*�*��'~>��!?C^�>.�>S5�?�,�>|�þ:�.���?��^?�AJ?�<A?8��>��=|��o:Ƚ��&�F�,=\��>z
[>/�l=�H�=_���
\�o-���D=�s�=1�Ӽ�W����	<6/��92U<�"�<	4>n�ٿ�15����)F�-x�&�^�����;�NսA��~��
g��C�Y�V��3�.;6�<�d 
�������J���?���?E��wȞ��`��5����۾� ?�bƼ���"���8gE��[����������%���w��6���ZG?Zm�J˿렿<
���,?m>?p#�?r� ��{>�ǻ�X.a>�O�=�}=Q��������cȿ0y^��q?l�>I�� �>��>���>��>]�F>�o��.X����=��?��*?��>=�-�6�ÿK"��)o�<��?��@EuA?�(����ԽT=���>k�	?�?>ͦ0�Rs�|������>"�?�Ê?�UH=�W�vw��e?��<��F��ۻw��=�#�=�C=���K>�6�>���XB��ܽ"m5>�	�>M`��<��?_�8Y�<�\>^�սKj���}�?��R�<�H��$��bo�1�`>%�}?��>�_5>�?��x���ʿ�5�V��?Q�@2�?$��>����>Q,߾��7?��R?^U�>?�;��l�LgV>���2���Qľ��b��u?><�?��`=8�ɽ��'����t�<v�=C��>ƿ]9��&��;=$C<��	����&���鎽�B��@u�
���"�=r��=�i[>Ԙ>�=j>���>v]?�y?�J�>�=�=�r'�������dr=^@�Y�o��ᨾ��0�=��JU���7澅l�Cx�;���U־?�@��M�=c�R�>ɒ��.��p���9�)�4?\X4>�E׾� N�gJ3����-����~&;g�ƽ9�Ӿe�5�ܾx�=�?%WN?�e��s�=������L����b?'�5��9�������o=��<��=��>EHL=ߓ��i8�� b��J0?f5?�c��������(>�� �T�=m�+?�?��d<v��>@�%?lo)���{�Y>�r1>ѡ�>�2�>x
>>���bڽ	�?9�T?�T��L���9�>�h���kx��y^=�A>��4�����-�Z>��<�c��xF��H���A�<�O?���>ϯ/�`��
�����=�B�UV?��?>m�>��h?r�*?��E��7Dd��J���=Ѵf?�^?s��=U�=�yľ'QξY
?R�D?��$>ҁ��*��,�w��f&�>���?��?b��Ӧ��K���Uy(�*�=?7�f?DmP��A���վ��<�|>�`G>6%?QK��">�\'?�'C��٩�qOÿ�>��?�� @��?6�$��MV��ִ���>�>nMj�y�ʾϺ��+�)<��μ��%?�ھ��*�n��H�-hk?OG?:6?A�������=�\���Q�?5�?᫾.�<����l����8ˁ<g��=om&���,�]x7��ž�
��v��:$��yن>�>@t��7>�>w;��*�9Ͽ�����Ͼ�l�h?.y�>h+̽ाǍj�C�t���F�mKG�3����w�>.Z>�۔�	����{�F;�(4�����>Iw	��Ո>2�S��Z�����,�!<���>��>/>�>���Q-����?ۇ���4οĭ���:�H�X?�L�?�k�?;F?�,<�v���{�*��?)G?��s?F(Z?�'��\�۩<�u%W?���"�X�B�VZ�n�T>�p*?z9�>�+@�jJk>�>�>0�?���>�����������.ܾN��?�}�?��DS�>B�?7?�c�|]��M��F������=4S�>4K�<èW� )���O��}3�@N?6�+?��L�u�xm?-K�U$S�����c���I�> �< ]�\6=�`��7q��ҩ�����5��?��@���?� ]��^:���?�/�>�k��P��5�W�_3>H��>u��>����2�>��������'>���?�+ @�"?ބ��ۨ���ἇ��?s�>��?��=�D�>�f�=�᰾A:&���!>Q��=~4�`�?4N?���>�'�=?�9�ψ.�0#E�F�Q���eEC�A��>��b?*�M?�_>�V���,�j`!��(Ƚ��3�nJ��=��6/��S�X�8>��?>b?>QAD���о��?ڷ����<��__ƽ��.?���<��?�m�ʾ��+��>��O?Ui>��ؾ�`��W���1�1��o�?E��?G�?�lپ	�8=�Mm>�~�>��6>�'Ͻ�������g>�s?�F���'����r����=���?A6@#�?�;M��?8�ھ �t��1������&Mi���?Ԙ��Q>��>CX��t��2���-�n��T�><�?�h�?ޱ�>��_?��n����z)�=��!?[�P?��?x�=�q�
4M�[.�>E�0�������&��ES?$}@��@<�?�/��H���%��A#���ܮ�y�;��=4|>��8ҋ=��6�7�˽HN&;�0A>k��>�.L>�,�>�d>�.s>� c>�ć��k&������榿�m6�����q�㨠�	����P��Ǡ�ڿ��橾����5��R5��G�罳T���T��=�RZ?fT[?o�W?=[?�$��� G>�����> ;���ө<X�>��0?��:?x�?��=Z��a������c��L.�����>P2�>)q�>�c�>���>��Ͻ`*>
/>Ra�>շ/>u�>=UN*�}^����G>u�>��>5+�>��6>$.>E1��X��a�j�e:����нJ"�?�����(K��H���Z��������=g-?��=�ޑ���Ͽd���wH?�^��r4�M(�+�>�)/?|�S?�>i:����_��V>����e�>(�=/j�z,t� �(���R>z�?��S>%�>�|3�=�:��Y���̾ώm>VH:?`��� M�7�w���L���Ӿ�4Y>�O�>�Ǽ� �}D���@����N���=R:?ޙ?�4ѽ���#N���X��wg7>�yM>��=�2�=n�V>�;��2���Qb�Wu!=���=��i>&B?d+>3��=�p�>�˚��uR��{�>;�G>��)>�??/$?ax�tX��"H��$�,�Z�u>9p�>���>j�>$�J�Hy�=IJ�>�$d><�
�aۇ�����c<�A[>��`Ma�X6x���t=!*��2��=�=����fh=�:%+=P�~?O��Ǎ�����u����kD?*$?���=��a<.y"��\��������?@�?5����V�3�?�!�?�x��?0�=���>^��>�Ͼ��M��?��ɽ�p���$	�)�$��2�?,�?u�;��s���_l�s�>^>%?��Ӿ'�>�_��{ޝ������j�C��<:��>e?�6���v�����?��>Y�Ҿ즛�`v˿�u�Eu�>�)�?��?X�m�3���Z+��T&?A��?5zQ?�q>܈���m�$��>��Q?r=?`��>A"��oV�;��>l�?
��?!-E>Ш�?&�k?��>�Ƹ�+VK������򅿔U�=���@�>{�>�mƾ��D�T����抿�j������q>�� =h�>�5Ҿ|��=��0J���A�<��>�>�`>p��>�z�>��>��>�T;�g���|[=��`��5i*?*�?���u�w9=�N����Y�l0�>F�W?���=Ν�X�>��x?<Pm?�(X?�S>d� �"���fE��5����<何t�=$�?V��>GA��1��>/�z����<�m�>�s>��:!��ۀ�u;����>��M?"��>���=� ?p�F?T��>+:�>H�>��ѳ��4���>|'?/m#?��?�H?������!��؊�eۭ�=�b�VfN>��X?�?��Z>��^�ߝƿ�xA=�12>�=s���_?��9?��9>=ı>⨐?y�d?Υ9?��=s���\ھ=BȽ!>(>��!?i���A��L&�*���{?�N?���>�*��6�սN�ּ��(t����?�(\?p?&?.���.a�Eþ�0�<1q#�*XU��<�;g�D�x�>s�>�s��K��=�>�Ұ=�Mm��P6��(g<�b�=�>@�=P27��l��g�(?�L�׍�����=�Y��L��m%= �>�O�SU?\4����f�����z���Fף�g�?�n�?�)�?2�Ƚ�[��H?2|�?Z5%?]b�>� ��s�����^N�|/��QG�pJ���<�>�Ǧ=9ᅾ%̖�h8���U|�y�=�J�:�?�>��?��?{AW>c��>�ȴ�ߚ(�xH�/���]�k�B3�ګ� Z��踾�z�[�D������ύ����>�'�;.*�>
?s�R>x�>���>�k����>�H>��l>�D�>��>�> �=I1'���JR?Y���%�'����䳰��1B?Bmd?�6�>�Ji�m���f����?��?�q�?-&v>Q�h�R,+��m?WG�>���@n
?y:=[H�Y��<PW��Q��KG����w��>?׽W:�2M��sf�:f
?�/?�����̾!)׽�.���$v=�m�?x)*?�%+���P��2o���X�ySQ�L�)���i��Ƥ�`�%��Yp��Z���{��y烿�E(��7=Zb*?�B�?�g�ƻ쾢3����k�u�?�Pcf>@"�>�>���>ɽC>͕	���1�\�]�<�&��G����>��z?�nl>�~O?�V? q??spF?n*>e��>��ƾo<?�@�=��w>a?��5?��?	�?�?�I?��=����-������3?��B?��?[��>���>E�Ҿ?aa���z����=<ٽ*�;=�'�=�*�=�r��k*��
�<)X>�/?��v=��T��� �c�>1�H?��>,��>t�5�B�=q� ?94�>��=?��>�b-��>��>���z�>Q�?�2��j��Wx=Eg��"���|V�q��>�>c}>ۗ>f��=��>�w�>6��>!.3�������=��g��H;=�?`?jW�>��>mま�$ؾ�_=�Eo/���>��>j`>��ɾ]�������#j��F�>��|?�e�?	&>t�=eˮ>��ľ��ھ�����<��(:��T�>r
�>is-?�v�?�q?�?��<SM��ˍ��|����;�?a,?>����ʾ��$y3���?d?�>a�mk�c)�;J¾�8ԽB�>�b/��7~�����D��0t����r�����?���?�#A�a�6��辵���S%���ZC?6��>m�>V��>O�)���g���DP;>�_�>��Q?9Ȼ>�R?0j{?9�W?�qP>68�����mӘ�*졻�� >��<?��?}�?�[x?C��>ܦ> Y3��[�߅�� "���꽈����a=X0Z>�@�>��>B.�>���=����OŽitB��̞=�b>��>��>��>>dn>��</�7?-��>���_������(�þ)ڔ��?��^?��7?�g%�ӓ�S�r�G�"�*��>U��?���?,EV?� ��>-y��b��y������>?f?RI�>���m���+5?=#,7?i�>�զ��r
�p����=�.u>��J?��0��ƿI�q�}�p��ė���d<�����e�g۔�"[����=������[˩�=�[�崠�����.���U�����{����>q{�=o��=$�=�a�<�pɼ�ݽ<c�J=��<�=�p�8;m<R�8�ıϻɫ�����t�\<��I=����ƾ�v?��S?I.?<E?ZWp>/�1>G�ǽvL�>��z&?��>t��;
��\!�ۣ��d#��MT�U�� �d�o����>p+���
>��#>S.�=#�,��)�=�a�=� �=B�����Q="�=���=ѹ=E��=ˣ >��>ֻu?E�a�v/��Or(��W">�X.?G�>Q�1>	'־�O?��T>!���J���J�e	�?�?{�?.
?�I�ή�>�7�"н���Or(��A�>�=>L��Cp�>L�o>=
��s����
>��?!"@�8>?|���+�ؿ��">q:8>k+>�R�{H1�j%\�{�b�S�[���!?W;�=�˾!��>g0�=<�߾NǾ�3.=�m6>�Pk=I���[�Yq�=֫y���;=��k=	G�>��C>���=�٭���=�L=�U�=fO>B�`���4��<,�]�0=V��=�b>�&>6��>l�?2�0?�{d?.K�>�Rn��TϾ%�����>���=S߰>�,�=�yA>n$�>��7?��D?��K?��>���=  �>��>��,�h�m����< �����<:��?
ކ?��>��_<#�?�Yr�Qb>�XEƽZ0?�L1?/�?���>w3�T���O"��p>����<0�/>i��=I��\���z�k��M��S���^>���>�Q�>�݊>ء�>G�>�ʝ>���>l5I>uۏ=��d=4d�=��,<�ֽ�b�<RI�UѼ=�I�=�޹=A0�^tZ<���=���v�\<�	;�=��=S��>�D>-�>@/�=F��-1>�I��-�L�,��=���*MB���c�3�}��o-�� 3���>>��R>����!����?4	Z>�B>
�?-5u?�t>���x�Ӿ	3���?a�S�Q����=��>CkA��+;�r`�>�M��~Ҿ���>iu�>�[�>��V>H�.��;;�; l=��Ҿ2�6�F�>p�v����R����[l����lO���d�'>�j�F?�����=\�?�OO? ǌ?�t�>S�轸־�*G>L����7<S���Sý"�?g(?$n�>�쾠h?�p�ƾH����>Ʊ=��T����2��Y�I
����>����`�ɾd�2���������h_C� oa����>�0S?Q0�?M~^�;�~�P�D��� ӂ�:��>g$^?�q�>h�?{� ?�> �˩���s��� �=��t?�\�?r��?C��=�=>̷�`x�>�}	?��?ᶑ?�s?��@�B}�>E(�;�
!>�a��x��=q*>�%�={6�=�?qB
?��
?�|��ş	��K������\���<~��=��>�m�>mDq>��=p!j=�C�=��[>�,�>1��>( d>���>�+�>�ގ����ؘ&?�p>���>��P?.�>*��v�;��o���,�,����=A�3���<Q��=I;�}En��Dݽ���>�mҿ/S�?x�>4A;��+8?9���Ǖ<B��>mđ��R�<A��>���=��>J>��o> �>�{>�?>WҾ�-�>d(��=4�>st�[H��ڞ�����>Cm���������P�U���ݽy`�� ��A�w�WV}��=����*�?�U9�X׀�b�����=|�F?�oo>v93?�ƾ�;�s�>��"?�'u>w�� ���6�������u�?���?�}>&p�>W�n?��M?FQ�\�C�N�f���mq���p�1Z�DϪ�誆����m���X?s9?�?�>N��>��?'��Fo��ǖA>�WQ�swL��`<>ɂ?8Hc��g���˾�Փ�u�'��BT���=?�~?� R?��-�� ��n�|At?�р?S��?�H2?���?�A!��>�K?�:�>Tl%?m�(?�Z? �>�=R�$�j��H�!��}��~��P�,�6Ca=o�=��=�ƞ=#����jt� �.=�ڽU�ڽT~=���<3�K����=��%>�O>\P�>[�[?�>�>��>?M5?�R&�$�9�W ��-?�T=�h��K䍾:���N���}�>��i?�a�?O�Z?�e>�2A�@���>�>k� >sZ>L��>g߽�8�3ӏ=��>U�>Z~�=;��`��T���|��E
�<|�>�9�>�Br>�Q�=���=Z;=���.���>�Э��/���$x�z����lH�d���
?J��?�n.?���Q����M�;슿z�U?�!?�t:?�1�?�<8@q$� cF�ڏL�"�{��Z�>Sw�<�>+���ſ�n��H/��*�����=!R��hڠ��[b>���t޾"�n��J����NM=�~�%]V=@�<�վu,�Ĩ�=�(
>ܷ���� �_���֪�	/J?W�j=z���bU�jn��<�>�Ø>�ݮ>ķ:��v�&�@�����*�=ɸ�>;>[1����xG��7��Mw>pw>?�Vl?�E�?Ð�������?��\龂߬�4g�=�+ ?�Q�>�}?.��=��<���V�*���Z��2����>�T?�4���h��������6���W�>�.�>:YA=���>qa?vl$?van?S?F��>�T>��W��^���#?�؁?��=e����t���:�1PG����>wv6?BNS��v>R�	?�,?��?�nO?R�?S�>�A��?�1&�>`��>Y�S������_>ɈI?{1�>�TY?���?g�q>��3�芦�o쥽L��=?5>��.?�� ?��?��>r#�>Ќ��L>�|��>�H}?vt�?M�<?*7�>-g�>쁇>�m?m�R<��=H�[>ͱ�>n�[?�w?�gY?�>&�P<�B��nS��Y���)�;�n�u�<�Z�={X�=�\ѽ������=s�='����el���| =�K=�*=���>���>����;>��Ҿ�����ET>��h�����m䚾[�v��=<l>��>�m@>�K�2ɧ=�ۮ>�o�>�=��~?�
?x
?���<U?S�Q��L/�V�>�e$?�{�=�n�;���s�t��A=0y?��a?f�������L?�	v?�c%�9�����ᾐ"�*�0?�X�>��f�O�T>���?9��? �-?�}���<'��PC��r ƾ4��=$)�>�!��{�V��>iE!?���>�Ł>�|�>�/���a����ʾo�>��?į?���?#>�bb�����E���6��d�a?�>�>�G���<2?�������jZ��,揾�z־5�������Č��)��|������R���h��=*?��p?�q?'V?� �Eo��b���t���T�Q��:+��)G���?��E�0Ve�x���bܾ4�l�`�=`�|��+2��O�?z!6?��K�e�'?�����N���B��=������K���=Р伨K�=�i=I0~���o�����1!?'�>���>�)?��_�ЧD�qF�8��H����f�>
��>�OJ>]��>�\���7dӼ�X��r���f=D{c>��\?�`Q?;�?8��d5��#z�	1)��߶��j�ͲS>!�!>ऍ>�x���7!�	�,���A�L�e�r��^Ƒ�<'���=�+>?���>�އ>�>�?��?�c�\§��;���'���=m��>�XX?b��>�%e>	�� �"� E�>��g?X�?��?)'¾n�'���j��'��T�?��?hm�>;�>T��%m�W|y�񈃿/�1�/^>ϔ1?�������t&t>J6|?\��=2��y��>������c��5�>�<�eH>��?���= 
>��
���6��灿�>���=)?��??��v�*�^>�+"?K��>5��>��?꽜>*�¾X��5?m^?�J?��A?���>�!=�M����ǽ��%��-=ȷ�>�[>��m=_^�=����[��@�~XF=)��=�
ʼ�%���<�
��)�P<Yc�<=�3>l�޿g�J��پ���i�� ��T,�
�v�`�6d6�/Ϻ��^x��d��4d;n���0Z���h�"����-��k�?��?���У�@������JԹ���?3\����������e��� ���Ѿ#���sD��X��QW��JD��$?�����ǿ����ྪ	?T�!?[>y?nY�a#�}v5��%>���<�����t�,����/ο[���3Ab?�Y�>HP�u���	�>M�>�'L>�Lj>+���h韾"=��?��+?H�>��|��!ɿ�����=[��?��@=6A?��'� >쾃7O=7D�>x�	?1�;>�e*����Ř��"2�>q�?�5�?�'=��W��-鼂�e?���<�|E�ؖ����=P��=���<�8�iI>`?�>{/���@�R:ƽ�5>�>���+���bP�T��<c�Z>~~׽z���� �?y�S���;�#�*�L`����=C�?x��>���=Y%E?��z�̲Ͽ�]8�:��?�@>e�?�?w��q�>�O˾�8&?2}`?�յ>�/L�,J��>�l��կ��@��m"�.��=��?�n>���;�V�%]�#�5|�<N��kǿ���(!�-�-=�|=���f�(�e駽ww���p��5�;�����I�=o�=�P>�~>�fB>�Qk>�;c?�Bx?�b�>�!�=��*�Z����z˾~	>=nf�Q�"�Uӕ��U���Ͼ��־>���������/�ž�=�]�=�6R�I����� �e�b�/�F���.?t$>��ʾ(�M���-<�pʾV����݄��ޥ��+̾Ζ1�{!n�͟?�A?C�����V���2e��y����W?�O�s���鬾���=+���ް=]&�>���=���8!3�X}S��/?/?? �þ����MB>�$�e�<VR-?�^�>�<U�> 9"?�\4�v��L>�)>>kj�>VP�>&��=�[��~�Ͻ�r?�AP?�����w��>h?¾U��u�:=D�=��:��X���t\>H�=װ��Rxɻm��P��<o�O?Nc^>6p)���ͽǰ#=sPѻ\l?��>Q̘>ȡt?ͯ9?Q�<�!��� e�;* ��g&>-LY?�si?�	>��<�r�ՉѾ�&?�"M?��;>��f�#q�P��M���O�>��?��,?�M��P��!P������@F?2�_?�V����y���
�<� �>8bR>�?��.�z�[>��N?mh��1g��1M���`"���?6 @Y�?	�Q���Z�
�=H}�>�O�>q���諕��@��H뾬���w��>�����A�Zp� ��	?�f?��>i��m�۾9��=zÕ��Z�?A#�?���Ԅb<���jl�=m��{Ƣ<EM�=���S!������7�Ǿ��
�����Mj��䬆>T@�9�O��>�s8��/��HϿw���kоVjq���?ѥ�>�Ƚ�s����j��Lu�a�G��H��j���>؁>%�� ��M{�});�=;���@�>���K�>0�R�_���굟��)<�ג>���>��>ŕ�����~��?YJ��u"οb����{��aX?�\�?�M�?�f?��L<�w���|�2��!XG?��s?�
Z?J�(��q^�D�8�� g?L���u�]���,�5�E��O>�r2?u�>��*�I>�=4�#>'�>�{>��'��WĿ6�����bӟ?�X�?���| ?�R�?�.+?�t��=����*��%�<0�0?��->5
ľY"��x>�Ą����
?;4?����`�K?_?/�V��`��0�2�ֽj/�>]M�;.�5�w΂�0�޽�d��_���S|�Z�?�E�?��?�4��&4���$?�I�>����5�h���T="��=1��>��>�r׽��>����j��h�"m�?�-�?��+?���	
��ǹ���u?�>q1�?�O�=/1�>�@=���Z�+=f8�=���=6{]�u�?�'N?'�>�η=�����6�Qn9�H�H�fj��ў;�_��>"�\?�nD?�,C>5��I������������q��p�n�[Y׽��1���9>�q>��Y>yr���&?�
�Y(ֿ�Ɇ�Ǚ�����>V{�>-e	?��mP�A�=T^N?5�{>W�究�5=���m��v�?b,�?l?k�Ӿ���<a>s�>�x>iK���.��<m��>s$?�M���Ǉ�u�v�L��>���?]�@I�?x�g����>������bs�pl"���Q������<Z?����-=�u�>�
� 0��Js��-Sn���>2�?�E�?$��>�[?�܏���+�ŭo� t?�,�?3����::>� �2�|����>f�7�:J��ژ ���?(�@A@��v?������&	��%ʪ�l���->�-=0�8> Jn�˽>%C���[�=<�e>�	�>�~>�7$>�V>�/W>�No>b~���B%�O-��橋���-����V �.\�D�Ԭ�N��̭�:/��<�Q�4�����ق�*F����l<nU=�!j?j�g?L3g?#�>��½�P�>�	:���p>G��^ #� ��>s*?]�)?�E#?��9��-�myX���v��x�������>NO�>i`�>�D?x~�>����	�Z>�g=��>C�>��=-�������)>�E�>��>?��>�C<>��>Fϴ��1��k�h��
w�r̽1�?���S�J��1���9��Ҧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�> ��v�T�3:>;����j�5`>�+ �}l���)��%Q>wl?��f>u>��3�d8���P��z����|>06?�涾.9���u��H�=^ݾLhM>QԾ>WnC�2k�Q�����zi��{=�z:?2�?rF��(ܰ��u�LD��`?R>L5\>E=���=zoM>�_c���ƽ5H�8e.=���=��^>�?3`">J#=<��>�υ���9�"��>T*X>:"$>��8?�@'?~����B���qD�DB~>���>(̌>�w>mB?�7�=@��>�X^>������w�n��C��?>�-��#;]�iۀ��a\=Wꩽ�	>�g�=�Fý�r���<��~?�|���݈���<涽eD?�;?���=�vF<�q"�����Y����?q�@s�?�x	�U�V���?=�?D4�����=0��>$�>	ξ�xL���?{ƽUآ�H�	�A8#��Q�?m�?&0�kǋ��l�79>_%?	�Ӿ�"�>�Q�p ���;���y�������>(�H?����i��0�"�J?	�>�)ᾥ���˿�0w��.�>F�?Z��?�:a�^���E�$�3��>r��?�K?b�p>h�ܾc�戢> �7?A�S?��>�"�>�.�P�?�~�?���?�?>X��?Ӣv?�|�>�~{���3���� '���Hb=�Y=G��>��>�����H��T��9ʊ�f�j����}�6>�\4=1o�>�޺�z���e�=-7������������>E�`>�'_>n�>/?���>�`�>��:�C��&I��B���8?�?�����_��T��ЈT�{�Y�&��>�*0?|�X ����>�"~?��?��j?�8�=~J�TM����п�b�����7&>}�?��>��<B��>����R~��N�>�٨><Ž ���׾���8���>�/?�u
?.M>��?,�'?�ި>�m�>Q@G��j���]D��G�>G.�>�@?6�{?�"-?�CJ��L)�����٩���p�&�=�j?�?��>^��L𱿇2�S�c�z0���r?&�S?��I��Q�>�:�?��[?3�[?�Nf>��'�ث�8Z���>U�?�ˆ��Q�Eq:�43����?���>N��>��3���=���=��9�G�,����>�1S?��K?}����8����2��<��T;��m<g��=�b=$v7>�C>�ὸx�=��H>�=p7�~2����=���=��f>�L=�><�o;��<,?�G�4݃���=��r��uD� �>�LL>���^?,d=�j�{�!���x���U�� �?Ƞ�?xk�?�����h��#=?��?�?� �>.J���{޾���1Qw��zx�9v�t�>=��> kl�������7���9F��$�Ž�K&�\�?0�>	?y4?%S>��>������ �$������D����1t$�,� �9��橾&K��B�н�֪�����.�>C�
��x�>8k!?�0>Uf>ί�>�R��6�>m�]>.�j>�&�>��>,�L>��>��l=-���FR?_����'���{���&(B?�ld?d�>�gi�.�������?���?�j�?��u>��h��%+�g`?�u�>����t
?��:=���C߇<Re��~��|u���\�q�>/5׽�:�M�x�f�i
?�/?=拼�{̾B�׽x�����t=��?�,?H�(���R��'o��V�74R��߼�)_�d>���"���p��7���΄�<��m�'���=F�)?���?UJ���ﾋ����k�8>�qk>�y�>x�>MV�>��R>�.���.���\�J�'�������>#�{?�}>APQ?��I?L�T?�??�ȁ>Vd�>HѾ��?,k���>Xw
?�>? b)?��,?4<?�?eyA>�{��d��Ӿ ?��?�1?֮?�L?����(�½�����=��$��O0�A�=3�;״ƽ�����A= �[>�?k�b�I�)�G���>jv6?�be>J�> �	�hK�v<]>���>K�?�;i>`;b�0)��wݾHu�>�ٜ?(�F�]	>�	Z=�3>�֟���|�}�q>�����=�ΰ������=��=r�>�0%�5��]�7��X;�/@+>���>�V?o�]>|��>K(����c$�}	�=>s)�>7B>�ť�_�u�t����Z�៞>���?|�?�N:�Ӧ=>��=��p�{��9DԾ�	��8�=�N�>��>ŽH?��?��[?� ?f�>e4�����݇�5�E2'?�!,?���>���0�ʾ�򨿶�3�G�?QY?:a����B)���¾X�Խ��>qP/��)~����[D��������ug�����?���?SA�7�6�S{�t����b����C?��>�]�>�>>�)���g�#��4;>ƌ�>R?���>-P?�C{?25[?��R>9�]EU���p"�Z
!>�-??��?�!�?6�x?���>�>g8.�Ox�w���@���򽍩��45Y=��Z>衑>>�>CJ�>���=�Ƚ�a��2�?��s�=Xb>P��>�K�>���>e�u>�k�<7?�y�>�8��g_վ�Ua�~D��NC��Jt?}Β?�0?��<�(�M�@�q1�+ �>
Ӡ?�u�?r�<?�s��<�=�G=�P��=9��1�>�B�>Ҧ~>X��<.!�=%�M>�W�>|�>E^����f/���r�f
?��@?
>�ƿ8�q�~�p�����e<L����e�W͔�%	[����=h�������ʩ���[�ճ������5�ء����{����>x�=>��=L
�=w��<��ɼ�Ž<.K=n��<0�=��o��m<��8��cϻѬ��\v���\<)�I=L��5�ʾ1�}?.
P?�?/?��??�|s>�|E>�ཱུ��>p_���!?���>�-_�]����q#��Ѫ�?	��"ݾ8�ھ�:n�-��)�>�6�w�>'^)>��=x����==��==���:��1=d~�=��=�O�=R�=��=�>@�Z?�Bf�Qu���Yi���>"V#?N��=�ݾ>%����8?��>��z��f���߾1�]?���?�*�?ч�>���O�>��}��jn=�yF=a���5�=��?;D����>6��>���"����g��$�?��?�[??�Ո���ӿ��J>�{>t��6o`��w)�2P�=�l�;A����-?��;��S�3��>W���
l�w7ھy��={p�>O�_>�{�<	�a�g&�=��<��;)j!>4��>��1>$
>L�����=�I�<¿%>yc�>sl�=�O��c	ٽ���&�='i�>z'>[l�>Fp?�d;?!�d?�e3>�����澧����(�>}�F��2>��t�7oI>zL�>A�3?�<?�*F?)%�>�T;�>��>q6&�WMZ��ʾqQ��7��� ێ?���??��>���S�O���r]3��lǽ/��>��(?FA?�F>�m�
����L �Ď2��=���1肻��s�y��盆��	� g�=p�#>�7�>��>�6>71>�=>��>"�>Ψ�=O�B�0쁽r��=��G=�=z�m>	��<y}O��Ԟ=�}=
�$�S�����G=�\<��=��<�D<�=���>�>�l�>L"�=۲��2>�$��JNL�"��=]��'-B�A�c�Lt}�o�-�y5�3�?>VRS>�3��8+��L?bX>�A>��?(Ht?J�!>/C�f�Ծ����0�b��N����= �>ĘA�$�;�{k`�<�M��xӾ���>�@�>Pg�>;�m>Yj,��p>�i��=����!4��Q�>�F��>�����p��a���k��D`f�����E?���>�=��}?s�G?��?d'�>N䦽Hվ9+>C�����<��/M|��f���T?�^)?�P�>a1�+oF���Ⱦ@�����>~E�$P��,����-���L��Տ�>����];�N2�����с��D�A��Vk�F��>l�P?��?P�i�uU}�i�M��3���c����>��g?ҏ�>�(?�l?}@��/8�X��C��=�q?ށ�?6��??��=�|>�µ�^��>N��>L��?�w�?Q]?̅��'0�>}�<�tO>�]�6�=z�g=YA ={�>�7?jq?��>�|L��;�����C�˃�kٱ<u��=�w�>Zք>�s�>;f>���=ڲ�=]e>(C�>T��>�(I>�j�>��+>ol��e[Ծ�?E9�>M8x>P)^?CY�>C�*������5f��P���6�z�u�	�� ��<L���������^��>�����j�?�>�a�,�I?%!%�ݩC>��<>���>5^>3H�>b�C>�b>�4�>���>�vy>�<�>؋r>���&>���}35��UR�K0a��p��"�>:���$�������%��L�p���v�^+��wx��ہ�k92��&�=Z|�?4=X�����"K�9�>z��>:HE?q���ԗ1��[�>���>��>;#�U ���ٚ��辫؁?4��?�gS>$n�>F2g?n@)? ��#���@�F�z*v��d ���j���c����p![�ު�P�E<8X?>Z?j�$?8�=�j�>�:g?�) ��圾�;�=����C�z��>��?
�ؾ7	��Zc��ܣ���;��X>��T?��?H�>?�,��������T>��E?Zt5?��k?
�*?9D?��a���+?�� >]�?��?��:?ݳ.?�
?�>�H{=K�����<ʟ½���m���y���<���=�=H3+�Gb�nJ�=2'%=�ݢ�wK��7ș<$-�h�#<��g�S5a=��=@��>@�T?l?k�>��
?m���G�DӁ�ֿe?���=����
��r����� ��F'>��d?�f�?Zej?��>������l>!?@>��>Gr>���>6^�.�k���->�]>�u>a���ؽչ��*����0N���z=H
">���>��i>�d�=)Vi>e��bɽ�j?G���ɅԾ����ܐ���DE�����U�?���?�{?-��4,�Mʿ�|���]?�(?�W?]�?�1>���\*r�GT$�ٳ��5�>B�6><Q*��j���S���90��jƽ�}j>��Ҿhڠ��[b>���t޾"�n��J����NM=�~�%]V=@�<�վu,�Ĩ�=�(
>ܷ���� �_���֪�	/J?W�j=z���bU�jn��<�>�Ø>�ݮ>ķ:��v�&�@�����*�=ɸ�>;>[1����xG��7��Mw>pw>?�Vl?�E�?Ð�������?��\龂߬�4g�=�+ ?�Q�>�}?.��=��<���V�*���Z��2����>�T?�4���h��������6���W�>�.�>:YA=���>qa?vl$?van?S?F��>�T>��W��^���#?�؁?��=e����t���:�1PG����>wv6?BNS��v>R�	?�,?��?�nO?R�?S�>�A��?�1&�>`��>Y�S������_>ɈI?{1�>�TY?���?g�q>��3�芦�o쥽L��=?5>��.?�� ?��?��>r#�>Ќ��L>�|��>�H}?vt�?M�<?*7�>-g�>쁇>�m?m�R<��=H�[>ͱ�>n�[?�w?�gY?�>&�P<�B��nS��Y���)�;�n�u�<�Z�={X�=�\ѽ������=s�='����el���| =�K=�*=���>���>����;>��Ҿ�����ET>��h�����m䚾[�v��=<l>��>�m@>�K�2ɧ=�ۮ>�o�>�=��~?�
?x
?���<U?S�Q��L/�V�>�e$?�{�=�n�;���s�t��A=0y?��a?f�������L?�	v?�c%�9�����ᾐ"�*�0?�X�>��f�O�T>���?9��? �-?�}���<'��PC��r ƾ4��=$)�>�!��{�V��>iE!?���>�Ł>�|�>�/���a����ʾo�>��?į?���?#>�bb�����E���6��d�a?�>�>�G���<2?�������jZ��,揾�z־5�������Č��)��|������R���h��=*?��p?�q?'V?� �Eo��b���t���T�Q��:+��)G���?��E�0Ve�x���bܾ4�l�`�=`�|��+2��O�?z!6?��K�e�'?�����N���B��=������K���=Р伨K�=�i=I0~���o�����1!?'�>���>�)?��_�ЧD�qF�8��H����f�>
��>�OJ>]��>�\���7dӼ�X��r���f=D{c>��\?�`Q?;�?8��d5��#z�	1)��߶��j�ͲS>!�!>ऍ>�x���7!�	�,���A�L�e�r��^Ƒ�<'���=�+>?���>�އ>�>�?��?�c�\§��;���'���=m��>�XX?b��>�%e>	�� �"� E�>��g?X�?��?)'¾n�'���j��'��T�?��?hm�>;�>T��%m�W|y�񈃿/�1�/^>ϔ1?�������t&t>J6|?\��=2��y��>������c��5�>�<�eH>��?���= 
>��
���6��灿�>���=)?��??��v�*�^>�+"?K��>5��>��?꽜>*�¾X��5?m^?�J?��A?���>�!=�M����ǽ��%��-=ȷ�>�[>��m=_^�=����[��@�~XF=)��=�
ʼ�%���<�
��)�P<Yc�<=�3>l�޿g�J��پ���i�� ��T,�
�v�`�6d6�/Ϻ��^x��d��4d;n���0Z���h�"����-��k�?��?���У�@������JԹ���?3\����������e��� ���Ѿ#���sD��X��QW��JD��$?�����ǿ����ྪ	?T�!?[>y?nY�a#�}v5��%>���<�����t�,����/ο[���3Ab?�Y�>HP�u���	�>M�>�'L>�Lj>+���h韾"=��?��+?H�>��|��!ɿ�����=[��?��@=6A?��'� >쾃7O=7D�>x�	?1�;>�e*����Ř��"2�>q�?�5�?�'=��W��-鼂�e?���<�|E�ؖ����=P��=���<�8�iI>`?�>{/���@�R:ƽ�5>�>���+���bP�T��<c�Z>~~׽z���� �?y�S���;�#�*�L`����=C�?x��>���=Y%E?��z�̲Ͽ�]8�:��?�@>e�?�?w��q�>�O˾�8&?2}`?�յ>�/L�,J��>�l��կ��@��m"�.��=��?�n>���;�V�%]�#�5|�<N��kǿ���(!�-�-=�|=���f�(�e駽ww���p��5�;�����I�=o�=�P>�~>�fB>�Qk>�;c?�Bx?�b�>�!�=��*�Z����z˾~	>=nf�Q�"�Uӕ��U���Ͼ��־>���������/�ž�=�]�=�6R�I����� �e�b�/�F���.?t$>��ʾ(�M���-<�pʾV����݄��ޥ��+̾Ζ1�{!n�͟?�A?C�����V���2e��y����W?�O�s���鬾���=+���ް=]&�>���=���8!3�X}S��/?/?? �þ����MB>�$�e�<VR-?�^�>�<U�> 9"?�\4�v��L>�)>>kj�>VP�>&��=�[��~�Ͻ�r?�AP?�����w��>h?¾U��u�:=D�=��:��X���t\>H�=װ��Rxɻm��P��<o�O?Nc^>6p)���ͽǰ#=sPѻ\l?��>Q̘>ȡt?ͯ9?Q�<�!��� e�;* ��g&>-LY?�si?�	>��<�r�ՉѾ�&?�"M?��;>��f�#q�P��M���O�>��?��,?�M��P��!P������@F?2�_?�V����y���
�<� �>8bR>�?��.�z�[>��N?mh��1g��1M���`"���?6 @Y�?	�Q���Z�
�=H}�>�O�>q���諕��@��H뾬���w��>�����A�Zp� ��	?�f?��>i��m�۾9��=zÕ��Z�?A#�?���Ԅb<���jl�=m��{Ƣ<EM�=���S!������7�Ǿ��
�����Mj��䬆>T@�9�O��>�s8��/��HϿw���kоVjq���?ѥ�>�Ƚ�s����j��Lu�a�G��H��j���>؁>%�� ��M{�});�=;���@�>���K�>0�R�_���굟��)<�ג>���>��>ŕ�����~��?YJ��u"οb����{��aX?�\�?�M�?�f?��L<�w���|�2��!XG?��s?�
Z?J�(��q^�D�8�� g?L���u�]���,�5�E��O>�r2?u�>��*�I>�=4�#>'�>�{>��'��WĿ6�����bӟ?�X�?���| ?�R�?�.+?�t��=����*��%�<0�0?��->5
ľY"��x>�Ą����
?;4?����`�K?_?/�V��`��0�2�ֽj/�>]M�;.�5�w΂�0�޽�d��_���S|�Z�?�E�?��?�4��&4���$?�I�>����5�h���T="��=1��>��>�r׽��>����j��h�"m�?�-�?��+?���	
��ǹ���u?�>q1�?�O�=/1�>�@=���Z�+=f8�=���=6{]�u�?�'N?'�>�η=�����6�Qn9�H�H�fj��ў;�_��>"�\?�nD?�,C>5��I������������q��p�n�[Y׽��1���9>�q>��Y>yr���&?�
�Y(ֿ�Ɇ�Ǚ�����>V{�>-e	?��mP�A�=T^N?5�{>W�究�5=���m��v�?b,�?l?k�Ӿ���<a>s�>�x>iK���.��<m��>s$?�M���Ǉ�u�v�L��>���?]�@I�?x�g����>������bs�pl"���Q������<Z?����-=�u�>�
� 0��Js��-Sn���>2�?�E�?$��>�[?�܏���+�ŭo� t?�,�?3����::>� �2�|����>f�7�:J��ژ ���?(�@A@��v?������&	��%ʪ�l���->�-=0�8> Jn�˽>%C���[�=<�e>�	�>�~>�7$>�V>�/W>�No>b~���B%�O-��橋���-����V �.\�D�Ԭ�N��̭�:/��<�Q�4�����ق�*F����l<nU=�!j?j�g?L3g?#�>��½�P�>�	:���p>G��^ #� ��>s*?]�)?�E#?��9��-�myX���v��x�������>NO�>i`�>�D?x~�>����	�Z>�g=��>C�>��=-�������)>�E�>��>?��>�C<>��>Fϴ��1��k�h��
w�r̽1�?���S�J��1���9��Ҧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�> ��v�T�3:>;����j�5`>�+ �}l���)��%Q>wl?��f>u>��3�d8���P��z����|>06?�涾.9���u��H�=^ݾLhM>QԾ>WnC�2k�Q�����zi��{=�z:?2�?rF��(ܰ��u�LD��`?R>L5\>E=���=zoM>�_c���ƽ5H�8e.=���=��^>�?3`">J#=<��>�υ���9�"��>T*X>:"$>��8?�@'?~����B���qD�DB~>���>(̌>�w>mB?�7�=@��>�X^>������w�n��C��?>�-��#;]�iۀ��a\=Wꩽ�	>�g�=�Fý�r���<��~?�|���݈���<涽eD?�;?���=�vF<�q"�����Y����?q�@s�?�x	�U�V���?=�?D4�����=0��>$�>	ξ�xL���?{ƽUآ�H�	�A8#��Q�?m�?&0�kǋ��l�79>_%?	�Ӿ�"�>�Q�p ���;���y�������>(�H?����i��0�"�J?	�>�)ᾥ���˿�0w��.�>F�?Z��?�:a�^���E�$�3��>r��?�K?b�p>h�ܾc�戢> �7?A�S?��>�"�>�.�P�?�~�?���?�?>X��?Ӣv?�|�>�~{���3���� '���Hb=�Y=G��>��>�����H��T��9ʊ�f�j����}�6>�\4=1o�>�޺�z���e�=-7������������>E�`>�'_>n�>/?���>�`�>��:�C��&I��B���8?�?�����_��T��ЈT�{�Y�&��>�*0?|�X ����>�"~?��?��j?�8�=~J�TM����п�b�����7&>}�?��>��<B��>����R~��N�>�٨><Ž ���׾���8���>�/?�u
?.M>��?,�'?�ި>�m�>Q@G��j���]D��G�>G.�>�@?6�{?�"-?�CJ��L)�����٩���p�&�=�j?�?��>^��L𱿇2�S�c�z0���r?&�S?��I��Q�>�:�?��[?3�[?�Nf>��'�ث�8Z���>U�?�ˆ��Q�Eq:�43����?���>N��>��3���=���=��9�G�,����>�1S?��K?}����8����2��<��T;��m<g��=�b=$v7>�C>�ὸx�=��H>�=p7�~2����=���=��f>�L=�><�o;��<,?�G�4݃���=��r��uD� �>�LL>���^?,d=�j�{�!���x���U�� �?Ƞ�?xk�?�����h��#=?��?�?� �>.J���{޾���1Qw��zx�9v�t�>=��> kl�������7���9F��$�Ž�K&�\�?0�>	?y4?%S>��>������ �$������D����1t$�,� �9��橾&K��B�н�֪�����.�>C�
��x�>8k!?�0>Uf>ί�>�R��6�>m�]>.�j>�&�>��>,�L>��>��l=-���FR?_����'���{���&(B?�ld?d�>�gi�.�������?���?�j�?��u>��h��%+�g`?�u�>����t
?��:=���C߇<Re��~��|u���\�q�>/5׽�:�M�x�f�i
?�/?=拼�{̾B�׽x�����t=��?�,?H�(���R��'o��V�74R��߼�)_�d>���"���p��7���΄�<��m�'���=F�)?���?UJ���ﾋ����k�8>�qk>�y�>x�>MV�>��R>�.���.���\�J�'�������>#�{?�}>APQ?��I?L�T?�??�ȁ>Vd�>HѾ��?,k���>Xw
?�>? b)?��,?4<?�?eyA>�{��d��Ӿ ?��?�1?֮?�L?����(�½�����=��$��O0�A�=3�;״ƽ�����A= �[>�?k�b�I�)�G���>jv6?�be>J�> �	�hK�v<]>���>K�?�;i>`;b�0)��wݾHu�>�ٜ?(�F�]	>�	Z=�3>�֟���|�}�q>�����=�ΰ������=��=r�>�0%�5��]�7��X;�/@+>���>�V?o�]>|��>K(����c$�}	�=>s)�>7B>�ť�_�u�t����Z�៞>���?|�?�N:�Ӧ=>��=��p�{��9DԾ�	��8�=�N�>��>ŽH?��?��[?� ?f�>e4�����݇�5�E2'?�!,?���>���0�ʾ�򨿶�3�G�?QY?:a����B)���¾X�Խ��>qP/��)~����[D��������ug�����?���?SA�7�6�S{�t����b����C?��>�]�>�>>�)���g�#��4;>ƌ�>R?���>-P?�C{?25[?��R>9�]EU���p"�Z
!>�-??��?�!�?6�x?���>�>g8.�Ox�w���@���򽍩��45Y=��Z>衑>>�>CJ�>���=�Ƚ�a��2�?��s�=Xb>P��>�K�>���>e�u>�k�<7?�y�>�8��g_վ�Ua�~D��NC��Jt?}Β?�0?��<�(�M�@�q1�+ �>
Ӡ?�u�?r�<?�s��<�=�G=�P��=9��1�>�B�>Ҧ~>X��<.!�=%�M>�W�>|�>E^����f/���r�f
?��@?
>�ƿ8�q�~�p�����e<L����e�W͔�%	[����=h�������ʩ���[�ճ������5�ء����{����>x�=>��=L
�=w��<��ɼ�Ž<.K=n��<0�=��o��m<��8��cϻѬ��\v���\<)�I=L��5�ʾ1�}?.
P?�?/?��??�|s>�|E>�ཱུ��>p_���!?���>�-_�]����q#��Ѫ�?	��"ݾ8�ھ�:n�-��)�>�6�w�>'^)>��=x����==��==���:��1=d~�=��=�O�=R�=��=�>@�Z?�Bf�Qu���Yi���>"V#?N��=�ݾ>%����8?��>��z��f���߾1�]?���?�*�?ч�>���O�>��}��jn=�yF=a���5�=��?;D����>6��>���"����g��$�?��?�[??�Ո���ӿ��J>�{>t��6o`��w)�2P�=�l�;A����-?��;��S�3��>W���
l�w7ھy��={p�>O�_>�{�<	�a�g&�=��<��;)j!>4��>��1>$
>L�����=�I�<¿%>yc�>sl�=�O��c	ٽ���&�='i�>z'>[l�>Fp?�d;?!�d?�e3>�����澧����(�>}�F��2>��t�7oI>zL�>A�3?�<?�*F?)%�>�T;�>��>q6&�WMZ��ʾqQ��7��� ێ?���??��>���S�O���r]3��lǽ/��>��(?FA?�F>�m�
����L �Ď2��=���1肻��s�y��盆��	� g�=p�#>�7�>��>�6>71>�=>��>"�>Ψ�=O�B�0쁽r��=��G=�=z�m>	��<y}O��Ԟ=�}=
�$�S�����G=�\<��=��<�D<�=���>�>�l�>L"�=۲��2>�$��JNL�"��=]��'-B�A�c�Lt}�o�-�y5�3�?>VRS>�3��8+��L?bX>�A>��?(Ht?J�!>/C�f�Ծ����0�b��N����= �>ĘA�$�;�{k`�<�M��xӾ���>�@�>Pg�>;�m>Yj,��p>�i��=����!4��Q�>�F��>�����p��a���k��D`f�����E?���>�=��}?s�G?��?d'�>N䦽Hվ9+>C�����<��/M|��f���T?�^)?�P�>a1�+oF���Ⱦ@�����>~E�$P��,����-���L��Տ�>����];�N2�����с��D�A��Vk�F��>l�P?��?P�i�uU}�i�M��3���c����>��g?ҏ�>�(?�l?}@��/8�X��C��=�q?ށ�?6��??��=�|>�µ�^��>N��>L��?�w�?Q]?̅��'0�>}�<�tO>�]�6�=z�g=YA ={�>�7?jq?��>�|L��;�����C�˃�kٱ<u��=�w�>Zք>�s�>;f>���=ڲ�=]e>(C�>T��>�(I>�j�>��+>ol��e[Ծ�?E9�>M8x>P)^?CY�>C�*������5f��P���6�z�u�	�� ��<L���������^��>�����j�?�>�a�,�I?%!%�ݩC>��<>���>5^>3H�>b�C>�b>�4�>���>�vy>�<�>؋r>���&>���}35��UR�K0a��p��"�>:���$�������%��L�p���v�^+��wx��ہ�k92��&�=Z|�?4=X�����"K�9�>z��>:HE?q���ԗ1��[�>���>��>;#�U ���ٚ��辫؁?4��?�gS>$n�>F2g?n@)? ��#���@�F�z*v��d ���j���c����p![�ު�P�E<8X?>Z?j�$?8�=�j�>�:g?�) ��圾�;�=����C�z��>��?
�ؾ7	��Zc��ܣ���;��X>��T?��?H�>?�,��������T>��E?Zt5?��k?
�*?9D?��a���+?�� >]�?��?��:?ݳ.?�
?�>�H{=K�����<ʟ½���m���y���<���=�=H3+�Gb�nJ�=2'%=�ݢ�wK��7ș<$-�h�#<��g�S5a=��=@��>@�T?l?k�>��
?m���G�DӁ�ֿe?���=����
��r����� ��F'>��d?�f�?Zej?��>������l>!?@>��>Gr>���>6^�.�k���->�]>�u>a���ؽչ��*����0N���z=H
">���>��i>�d�=)Vi>e��bɽ�j?G���ɅԾ����ܐ���DE�����U�?���?�{?-��4,�Mʿ�|���]?�(?�W?]�?�1>���\*r�GT$�ٳ��5�>B�6><Q*��j���S���90��jƽ�}j>��Ҿl�����\>�B�D]�K�k�C�G�����HM=\����=����ܾ�����f�=Á>�E���:"��5���z����J?���=s���=W��Ѹ��>��>PZ�>6�>�A�|��	@��ծ��/�=�~�>2>�9ȼ$m󾛿G�x=��u�>�eG?�g?a�?Yhb��Zq���>���k`���l#��8?�F�>~x?��=>� �=M���C��?d�DwD����>��>i� ��*G��������7%�s�>��?�O3>@�?�L?�3
?�
]?N�?2�>3��>���*��)�&?t@�?%��=RxŽpSG��5���A�GI�>L ?���л�>��?WW?$�#?$�J?��?���=����#7���>�V�>ĚW��
��'E`>ݠJ?'[�>��U?]��?��G>�[2�0S��v^,�R�=3?>�5?�_%?�d?�3�>l��>����_f�=�L�>W�b?w9�?!�o?c��=Z�?�!2>��>7�=[��>T�>��?T=O?1�s?��J?���>�<N6��O����s���N��g�;�H<��y=��5Lt��?���<Ҁ�;�[���I��U�OD�������;���>~��>_����f�>��E���={#>�M���[���Ͻ�ۈ=8�^>��?K�`>����{�!=�:�>�u�>B����p?��>#�?��=P%��z�����{Y�>��k?`�8==�o�����Hq��K���?j��?�ԅ��~���b?�]?�^�R=���þz�b�h����O?d�
?D�G���>�~?�q?���>��e��8n�M��<b�!�j�ʶ=Oo�>nW�^�d��<�>��7?SP�>��b>5$�=�p۾��w�g��L?�?���?���?�,*>��n��1�d�������Z?�[�>���x="?p��ξ1j��+���{��鳾���ᘾX<��1z��W���B�V��=�T?�Bs?��n?��\?����e�b���\��3��Z�S�] �yi�Q�D���E�'PE��o��F�� ���s���3B=ݬ��U�-��z�?(�%?�ѽ�b�>'g���y��jrȾ��@>����U3�k�[�\���&�=s�=��M���7�GM����?� �>F��>C^;?+�G��f6�#3B�3@1����r|�=Ⱥ�>c��>���>Kö�R������־�\��7��^�g>&�s?^SZ?��s?���=�Xa��E��C��ԯb>�?u�Ǽ=��4>e�>���a==��׾oB�q�����F�]֛�JI-�n+�=Z�G?a=NԦ>��?�8?�P�K^⾙�~��%%� >i��N>Z�?R�>���<zd�=x�^��>��l?ܹ�>��>�a���W!���{���ɽ���>��>���>��o>�G,�V
\�Va���~���(9���=��h?n{���`�_��>y�Q?�/�:́J<���>�dv���!���
(��4>�?i��=��;> ržf�.w{�A+��im)?{^?�L���*�$�>�`!?-f�>�>�o�?��>��þо~:5a?��^?�I?*a@?���>�#-=5�����Ƚ��&�&W)=p��>�oZ>�l='~�=S(�_�[���� ;= e�=�����?<���]+S<�� =-'1>vۿ7�K���ܾ����E����4������͊��p$��д�ܤ�����`g���/��PP���l�37��֠t���?��?��+ꊾt���G�2����D�>�k��O���*���J �ǣ��6M��-��c{"���S�#�j�ݞc��?ֲ��G1Ŀ�֡�O�˾�0?�<?�AL?f����7���F��N�<�����νc��d�����Ͽx���ҞW?b��>kbǾi��ձ ?��d=��#>�N> ��1g����=�Z�>̃8?X?/f;���¿�����=O��?S	@4D?�)����VE��"�>ϔ/?��s>A�߽�j��FT�>|r�?&Յ?����g�J�a���W	f?ބ�=dn��˻��=���=�#�=����&>�}>I&��E��(�?�Wt>��">j�_��ȴ=��\�_�+��~>�O%�W��3Մ?"{\�sf���/��T���T>��T?�*�>d;�=��,?K7H�_}Ͽ�\��*a?�0�?���?=�(?�ڿ��ؚ>��ܾ��M?fD6?���>�d&�%�t�܅�=�:����y���&V�=��=4��>�>ڂ,�Ӌ���O��H����=!(���&Ŀ�x1�Ϗ?��
T>ϲL>�9����)0����ؾ 䋾��澑^[�;�S=3�>F�>a;�=\Q�=K:<��\?
�? ��=3��=�I��#����3�g2}�����"����P��Kھ�_�*x���6��#�ub1��/��c˾�J?�^�n=lR�}����(�73]��B��,?W�>�ݾO#L�YἿ�վld��r���y��Ӿa	4�	n��ş?�"D?ᢄ�H�U��7��O$�/���
6N?L��L�G���b��=�x#�"�<A��>�j�=��=W4�=N���0?�*?��������>���3A=��,?��>_f�<g0�>܋"?&���O��n2G>[>v�>���>�>b<����P�?=LU?n��#���g�>�g���s�r�D=�[>k�:�@pǼd<> F�<Dh��	�4�H�����~<��S?�'�=m�L�
7M�F�����r>"�=dTO?j��>�ى>o1{?� ?�{>4o$�h}j�ӫþ��h>uog?�?�f>]��Ry/����`E?��?_-�>�G��c���&.��5��m?X?�#�>�/a>��?���_�]Ѿ�|�>S�v?��]�@�������U�=ݤ>{`�>&��>��7�v�>�V>?�M&�w>��We��7�3�G�?�@/r�?<v<���f�=�l?�6�>�M�xpǾճ���U���v=�>L����u��& ��1.��7?�y�?�E�>��S���X{=đ����?%<�?�1���)ν�)/�5��3��X5�<�e=��e��+�[^7����[� �
���>�h�>@@sjs���>Q��ѿ&��@4��i��F�ԽoV�> Y�>�p�=�U���B���p��hM���t��&��h��>��>0璽c���?={��*;�A��>@|	�~/�>�BQ�AI�������R)<�>�>�g�>���>��nj��M��?2����ο�ʞ�
x���X?�ў?23�?��?$aZ<�t�7^|�n�!QF?�r?�.Z?E���Y�v�+��h??����^�$ 9�YXB�~>&�2?��>
�-�JD�=��t>t^�>�&>7l�����p���V˾�r�?�w�?k�w��>܄�?�D5?ܓ�^!���̛�!�$�N�&;��.?O�;>�ZѾcg��rH�E���,��>0&?S�4�`��]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�1�> �?�+�=LT�>���=R찾 +���$>o5�=��=��d?w�M?��>�
�=$�7�T/���F�C�Q�F��C�v�>�a?�CL?KYa>�z����1�!�}-ν��/�1��?�0����[�4>�=>E�>�D���Ҿs?�����׿}p���h���'?djw>���>��[��_u=��G?��>/��|���׭��i㷽��?#��?�?��Ҿ�|��q=���>o®>��i<��u-����J>�.9?����"ag�� d>ڞ�?��@�k�?#�N���	?I����Uv�����7�[F�=w20?y[羑��>�`?
^�<%h�B��'�y�B�>�Ӭ?��?H��>Іi?,�g�6�:�/sx�U�>y?q?mkx��g�=Q>�� ?m��+W!��czU?DK@%�	@�T?ۓ����,}���Ჾb����>3+>��>��s����=�V >k�������R=oy�>�8�>���>v[g>�R�=��=�B��P'-�|1���B���a����:Y!�������⦾P������Q�ݾ|�8�@r,��VC�!��;_y��Jd���`=*�`?�q�?��?���>���v�G�����q�<5<}���f>xf�>0� ?J�a?Z"E>2��7m�kX���Uu�.�U�1�?��=�ޭ>�`�>"s2?�%�:o�=���>�q�=��=�&?�Sx=�҆<��^=OSY>[0�>8)?D�%>�s>tƳ������a�r9k��\�����?�m���RR����`ڞ���þ�`�={�)?`>⭒�N�Ͽ�����I?��������0�h>�,?/�T?�� >g%��ӏ_�F>]3�tXv�Q��=���j#w���-���?>�?�}f>a#u>ѕ3��[8�ۻP��u���t|>�6?j���+r9�\�u��H�Ԁݾ!M>U��>�hD�0m������� Oi�~�{=&t:?˂?�ͳ�밾��u�C��LR>rj\>H�=�p�=scM>�Pc�]�ƽ�	H��a.=���=��^>��
?��=Ls漰�>�.��Xq��m�>��>�w�=Ln5?�NA?����5�<�U;��z�~�=�?��@>�}S>��8���R<� �>^E�>GS<��A�0����=�@�>k��6��ah��ɩ=����G*>�U�>�	���Y��g3<�~?���%䈿��0e���lD?X+?� �=J�F<��"�@ ���H��F�?q�@m�?��	��V�@�?�@�?%��l��=}�>׫>�ξ�L��?��Ž4Ǣ�Ȕ	�4)#�eS�?��?��/�Uʋ�3l�u6>�^%?��Ӿϝ�>)��j��,|�T|��e �7O�>��A?�Ծ��8�X�����>�?����eF���ƿT�c����>���?�?��d�����V[I�vM?��?�sK?�8>vz�<2/����>1P,?�K?s�>QQ����?("�?�e�?<�3>�-�?�τ?�*�>�<f>�Y9��ԿC�����>�70>�_����^>=���%U�����)b���M�k[Y��X ��B�=���>ʌ��Y¾���=��Ͻ����|�B��8"? ,�>�W�=�/w>ߗ@?��?�{>H�<	/=k���ѹ�m�K?���?����2n��Q�<Ꞝ=�^��&?pI4?Aj[���Ͼ�ը>�\?V?�[?d�>R��H>��F迿C~��r��<9�K>M4�>YH�>�#���GK>��Ծ�5D�bp�>�ϗ>����?ھ3-��_E��:B�>�e!?���>�Ү=�#?��$?|�>3��>o�/��ҏ��,=��M�>7�>I�?J�u?v�
?�§��+��ʌ��k����b�� `>�(s?�s?Tք>k�������s�e�::����d�c�?��X?������ ?��?�ZP?��??�+>�6���ɾ�{�	�>��!?,��$�A���%����?�?��>����ҽ)ͼ��1����? �[?��%?�%�.�`��¾<��<os�NP����;�6�A�> I>ш�u��=٭>PZ�=�n��6�7�\<ִ�=[֓>��=��6�hk����(?�(=���V�a>��O���n��e>}~��2U>n�]?��R�{�h��b���w��Q��{B�?�;�?���?1�����k�g,o?�h�?��B?<K�>b�ɾ������)���Ⱦ�y*> ��O�>�]x>}n6<,�ľ ���}���C����ν�YM���?S�>2�?��
?�=Y}�>,�;��"�2�������V�?�9�EV.�ۭ�9���?c�9�Xu8�b�Gƈ���>J���ԑ>��?��5>VZ>�ï>��xu�>�43>@>%�>��u>V�T>�P"=�^�<�=_D?���i���M77��WݾXp$?�R�?6\D?�x"�ʀ��rԾ/]:?��?��?�1�>��]���6��j�>��%?�ܗ�ն? eŽ��=嘽�?���r��vsK��� =�>Yר���E� oY�9�/��T�>�7�>)���B���;�N$����w=�̄?�B(?m�(�oBQ��Hn���W���R����X�k��n���$�R�o�eh��!��._��Tm(�(�/=<�*?6f�?��]�����y�j��?��3k><!�>�H�>��>��I>v��0�=�]�z�'� ΁����>�}{?� �>#�I?X/<?��P?m]L?��>�٨>L^��<��>^9�;Rw�>ua�>m'9?��-?Z^0?^�?+?q+b>`�������Q�ؾ�?�d?�?"?6�?3ᅾ��ý[���՝h��&y�P$����=��<Q�׽5�u���U=	�T>��-?O.h����������,?Wu?ju ?�a��V�^�|��>�jH?��H?���>�Iž8�n��M/��j�>��m?��ǽ8o�<�>>�j->�����m<FZ�=��<�Y���z=�?�����=�E�=�	�>�q�=��bm���^-<�����z�>D�?T��>}E�> 3��F� ����(�=�yY>S>��>�\پ����$����g���y>#|�?�~�?��e=+��=<��=fS���/�����/��^��<{~?�C#?�`T?���?�=?�`#?�>M)�eI���^��4��J�?�m?�@�>	���4Ҿ$����*�?���>hpg�rZ�+8�p�޾�\޽���=j�?�+(���X�A�J7=d����\��?�e�?��@���<�����"�������eJ?���>>E�>��?σ�5�X�4'�Js|>��?��S?B0�>��d? ��?+%W?���>��F�>��ƞ���h>6<h>=�?��z?s.�?�q?q�>W">a�'�����ɼhY1��.����}=Wx>��/>)��>3�>M�=Vc"� ��<�)I���=?+o>�?���>��>�~�>W/e<�0E?⃰>��$|����|���䲉�xFk?�?'?��7>2�&�p�D�g�����>�̹?v��?9)L?}Ɓ���=fT^�0Ɏ�A���fO�>�$}�u�>��佽�>�t���C>$�C>�T�?����ﾏ�>��'?~�a?g�Ҿ��ſ�q��/q�\K����s<��|d�����T�[�*B�='Ę��%�I���1\�Y���
���a��2���|�H'�>P�=#3�=]A�=Ә�<Kg̼���<�E=V-�<��=��p�-g<��:�PL�����f�K��<<%E=�ֻ��־.̀?��E?Z�,?�HB?iW >M�9>�f<��L>�*=�M�>0?�=��i��|��T��HI��Z���ѾY����|_�er��~}q>ßཱིF�=�":>�~�=�<��=��=��/>w�޼+�V=?��=X>�N>�q�=�� >\!�>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?Ati��d�>M���㎽�q�=K����=2>r��=y�2�T��>��J>���K��E����4�?��@��??�ዿТϿ5a/>�A:>�>�DR�M�0�*p]�@�b�]<V��#"?g;�̾��>��=�'ܾfXž_� =]�1>��o=���rZ�旙=q�w��\==�Xf=���>n�F>m��=;'��?��=�<H=���=�DP>�{���$�ij)���3=�8�=aod>�n%>��>JV?b�+?&�e?J�>
0H�z�ľ:���u
�>i�:>�׭>�;=Cu.>�ܭ>�!3?�@?�B?�ޥ>�˺==�>q��>��)��bl�ݺ��,ؑ��ƪ<�f�?��?ǲ>Ǽ�=�O�s����>�0���t"?�7?��?z>!�����Y�uC���{>/����!��� ~�0F�kZM�4�ͽ�њ=���>u�G?���>�.>�3<j}
=I��>�>�ɋ��9�~�*=M�=���s>�ֽU�O�=���5���O=A8�����=�4>�Z'���>>=���=6�?XPd>�N?:-$>۠�u�S>z<�ۀ5���>J-��9�N򃿇r�����G鼢,�>�>�ڗ��雿��>ۼf=ز�=5��?!��?��N>��8�m%����ꑠ�T$����Z=�57>��T��EQ��`���o�+-�/��>���>��>��l>�,��?���w=����a5���>w��W��� ��)q��;������i���κM�D?�?����=�~?�I?7ݏ?��>�G��h�ؾ�N0>m!����=���'q�������?;'?��>���D�6"��x@̽��<Zކ�࢒������h	�3�y;e�V��x'>��O����.|��$�I��f5c��P��;P�>�/G?3��?∾Q�n�Z+����4����>�y?u1?�y'?��b?�&=��m�f�O���.>�D?,�?�p�?�|�=�O�=g�����>��?`�?�(�?޲o?6,+�Lv�>m��<έ>tQ����=�>���=���=�O?ko?��
?������3��
����
^��6$=��=��>��>Γv>�9�=�j�=���=�e>;�>g�>��g>�G�>��>
S��Qﾐ�-?+c>��>u�!?��>��*�b-ɽ�ؙ=��]���e��v�罙�L��ӵ=��<�J(=�h�D��>ÿ5p�?�.G>��<�?������[��<`>�o�=,t�����>�T>��>9��>��>V��=��]>U��=�����L=>37��*�����3��v�����=#��3�c�i��㮾B����hѾ
Z־��C��Ē� 6�-�<n��?D�ؼ�a��67�R�3�r�>YMg>8_
?�@ž�>���=i�>��?q�־�J��.���\Ҿ'L�?��?>c>L,�>ܧW?�?W�1��2��VZ�Tu��A�(�d��`�F؍������
��Կ�e�_?M�x?<_A?h��<3z>��?'�%�׏��I�> �.�W;��=;=[�>i��9w`�ŮӾМþ���*=F>��o?'�?C?�tV��!f�9@(> �:? �0?�Rt?�V1?c;?͝�*�#?[�6>ٛ?4�?v�5?��.?��
?�0>p��=l��s*=���ո���'ҽ��˽��o�2=�~=1�A��	<�=��<��ۼC2Ѽb�;�����'�<��:=rˣ=}��=P٣>v]Y?��>	T�>��6??/�<G2��Z��z�0?|�P=�끾�����඾����n�>7q?��?H[?�A=>�s@�#�C��<>�]�>�>]�D>6I�>N���z4�rs=��>Y�>p�=г��;�k&�n���:$�<��&>�z�>Y�|>�=���i(>P��Hz�H'd>�3R�m�����S���G���1�Ww�w��>�K?�?�8�=�g����f�U)?\�<?�<M?Y�?�'�=q�۾)�9�h�J�x��ҟ>|ձ<�������� ��b�:�fS:@�r>�=��{B����a>�����߾�Ro��J�X����~=.��	%=ښ�A־x�u�l��=Ht>�[��{c"��Օ��_��dK?�To=x��+�A�{����v>'��>�Ү>=�N�CM��(>�?��F0�=��>R�?>GӼF���F�; �$Ky>�F?=΀?&��?�E���w��HG�S�
�I���H�>��
?�AU>4ؙ>�K>�w�=��پc2,��>�@A7��?��f>!�"�5(O��7��c���]�L��>~�?*�|>Y\ ?��'?��?V:?Ow?Z�>�p\>�0<��g��A&?��?��=l�Խ��T�� 9�[F����>�)?��B���>~�?��?��&?��Q?%�?^�>`� �`C@�U��>�X�>��W�gb��S�_>U�J?���>n=Y?�ԃ?1�=>��5�1ꢾ�Щ�hT�=�>i�2?�5#?��?��>��>�@����o=͓�>�^a?���?��k?��=��?h#/>�>�T�=���>N�>�?�`K?ktr?΀E?l��>]X�<!���(%ǽa������)�ڻ 	b;�Dy=Ze&�e�J�_���v<�ߞ���2��i��p�����x�����-#�>��=�(������4���۞�=���;Kٽ�þ�V�=��=��R>୼>l�%=�@ʼ.V�=�>�>��?*�E�-?���>�)4?��-�>�l�����㽨¨>x�C?��=*u�.!��Mo���<7�j?]X?O�T�`���J�b?��]?Lh��=���þD�b����b�O?A�
?p�G��>��~?^�q?3��>3�e�#:n� ���Cb���j�1Ѷ=Br�>>X�M�d��?�>��7?�N�>�b>Y%�=�u۾�w��q��t?{�?�?���?�**>g�n�O4��}���l��f_?=��>+?%�i�?�$�<�B����s�����D��{��g����:��+с���p��@��WN�p�?y?�߀?4�V?�H���W��y�Iu�� I2��������;9�ed5���Q�e����0������پ@V��@��@ �]�?�d*?��ý�q�>�T��J9�pǾ�vt>�ެ���0���O=�<>�8M=���=�_�"g�c�ľ�'?m��>���>��3?$=M��44�Y:��1���Ǿ�u�=ڊ>��>Fi�>�����k����2�ܾ]����۽d�b>��{?I��?븆?K�='�)��V����7����=�{��9>$s�<��*>	`������n�,���S��!q�l~�3���_&��x�tG6?=��>P��=3��?��?<X�����<��}��1\��a��> 6�?�m�>E�<>@A�>�;��D�>Z3l?+M�>}��>z���� �4�|��U̽Q&�>��>��>�yl>�+�ƹ[�v����⍿�_8����=jRh?o��Nuc��<�> �Q?+1��W&<>\�$0!�5g�I�(�Tn>�?46�=ɤ=>rƾ�f�5Az��C��.v)?8�?�Ғ�4x*�r`~>�"?�!�>�c�>��?��>��¾�蚹�}?��^?��I?�A?���>��=�Ů�F�ǽ��&���)=�&�>AZ><i=���=�����\�����dE=�I�=}�Լ;/����<�ǣ� �T<���<�3>1Mݿy�H���޾ѡ�&���r�n��7$�����&�h*���Ř��ek����r�-�.�S���u�=ڊ���q�a4�?�J�?�����񑛿��~��S�@^�>�z��2��#��[�dD���^ܾ"i���	!��uR��)g�J�]�^@'?h�����ǿ񍡿��ܾ%�?gI ?��y?n�y"�HW8�}o >��<џ��<�ؒ����οE�����^?���>Q]���� �>֠�>5�X>�q>@^��.�����<�:?��-?�C�>�r��uɿ������<���?��@�.?�}M�M��rm����>xZC?���>{�X��}��W����:?=�?/0�?��g�Y�5�u���9�9?+eq>�e&��$>=��>uA>�>�����=��>��!>�Ӌ�1"�<N૽ki�>��A\4�ٛ�=¶��۝�=o �>���<��`K~?�B0�9I���>>w�Й�M�Q?}�>��3=1*?��a���ؿP�j���v?�� @��?
+G?����x<>�y�{�Y?��*?�ڄ>��꾫ja�`5�>E��0E�f�ɾS�l����=��?�q�>n�S��⾪��6��,=�[�ƿ��$�xj�y�=s����[�j�+��G�T�m6��;�o��}�q�i=��=S�Q>~Y�>P�V>Y�Y>x^W?�k?�\�>ܱ>(,��y���ξ�?�y.��C��ʪ����ޣ��ƭ߾�	�s��C����ɾ�P}�T�<?�Y�R����7��rf�E~"�Z�@?�[	>9L�,�A�Š6�*뇾���� �?����`�9�5�^� )�?9�,?����CI���4�Ol��u�=l
�?d����&j־j�<�x�==:3=���>+쐻�v�>+��;�J
,?4?x�ľ����I>D���Q���(?��?�t�<-0�>�#?��)����#�>��H>�:�>�5�>�0J>0����
��8I?N�Y?��d�ۏ��'�|>?���v��G,>���=� R�a��C�@>��=Z"���'<�܆��*ֻ>�??���=X�6�������2�����\? �? �v>L�q?�&?�R�=����b�!�����="�?��}?��'>A1A�߈��K�ƾ�X4?���?!�>KH�=��̀j�w��O�M?G4e?���>x�>�T��#���jܾ-�>��~?^G\�o]����¾Sf���}>���>���>�����>�($?�B�:v���н����Tߛ?*@��?{���v'�^ =X-�>I,?Er�\����j=票��W>�j�>��Tb�cAC�ὺ�R=?@v|?oS*?���-�>���V=xK�UΫ?T��?�rb�z��}�o�s�ߞ�����<�}�������p�������7�fӺ��
��ݿ�K�ֽ��>nb@
�5��>�����ֿ�}ҿ�>��X��\�7���?���>̽�ڢ�c��炿L�N���W�P����X�>��>�K��������{�\~;��ߞ����>g����>�S�J��X퟾Wu5<U�>u��>�݆>�?������ұ�?}-���.ο���G��K�X?X�?�b�?EV?C+<<]"w��
|����&$G?�ws?\#Z?�$��Q]��5�P:j?4���K`���4�W�C��]U>�1?*r�>��+��bh=��>�C�>FZ>	�.��Ŀ����cm��/��?h�?{�hR�>��?�,?D���������SK)�u�:��A?�|2>������!��<�����S
?�`0?9�������_?ŕa���p���-���ƽAϡ>�0�6c\�Y��Ș�[e�
��sQy����?�^�?��?&����"��1%?t�>p���J4Ǿ���<u��>b#�>�=N>d�_�a�u>!���:��e	>��?�~�?�l?m���@����=>��}?v$�>��?�n�=�a�>Bd�=�
-��k#>�"�=��>��?��M?�K�>�W�=��8��/�'[F��GR�*$�+�C�0�>s�a?�L?WKb>���� 2��!�duͽ%c1�#P��W@���,���߽:(5>��=>:>f�D��Ӿ��?<3�e{Կ�蘿@qR���=?V�>7L
?��
��ۙ�-c���s?ܙ�>�������ȇ���ec�?���?��?��Ծ�V�p�=���>m��>Y�1Xܽ�~Y���4>�]2?�Ӓ�$Tu�f܃��ԁ>��?p��?I��?�_�?�X���v��na��M�;h�1=��3?5h߾:�>���>1I=��i�D���SO�
��>9�?#_�?�>�T?�#p�g_�{6->�|Y>��6?���>�ɑ��9ɾo��>��>Gt�i蝿0�\y?��@b�@���?�v���6޿:����B�����td�=��=9�>�Ž���=m�3<X�;
����>T��>�U>�
p>e�>��9>�	�=_����|@Ϳ�K���f��p9����l� F������ �ݬ��S릾���PM���q�Ѿ���Ᵹ��z��2^?�OL?��z?�,?����F6>�c��n��z�<�lm��Η;�w�>M+g?��;?���>d:��l�\v����:J�#��>|D�<I�>(�u>I�x>��<���>zT>���>E! >xÆ=�J�<\6�=n
�>�%�>��>k��>~�>��>w\���ݯ�
�o�����(A�����?}䣾pO�����I5���>����=4�*?�
�=�^���Q˿�z��ܵJ?y��՘��ֽ���=�7-?"�S?��>����?1">�7� ,e����=�X��9�z�;Z#�whC>o+?��C=��P>��8�+.���w���о�-�>��M?�׾A�k�hCe��$?��ڜ��%>�Y�>����q4��m��(^�V?��-=�Q6?.u2?����pƙ���'��;oH<>H��> �l>(��=���=[K-��֍������G�=��>��>/d?���=��-;&r�>k���ӄ��H>nZ>�k�>�6?��1?��&�r�u�}��M-��/�>��?('�>O�>��T��,7>��>|>��5���(���������=�B�=��������O=��b��2>)�;R8ͽ޵t�V�<�~?���(䈿��8e���lD?W+? �=a�F<��"�B ���H��F�?q�@m�?��	�ߢV�B�?�@�?��"��=}�>�֫>�ξ��L��?��Ž8Ǣ�ʔ	�=)#�iS�?��?��/�Zʋ�7l��6>�^%?��Ӿ�l>�mʾ�$��6~f��I�����=ٲ(?��X?;Q�v�d�
�<�1?��?4�����z��sĿ�?j��?�ݼ?� �?K"��+ȏ��g�?jJ�?�??v�\>��վ(���8	=�cm?{�g?�;p>Sg&���k���"?�ՙ?�AL?m��=/�?E@�?���>}��=u�%�辿�\���]>$�u>B)j>�;=���ϫ7�v ��z��n��-O��Z�=�k>v��>���=#Ȯ��Z}�6�R<�4˾�����?@�H>�>���>?E��>a�r>4�<`ҽF�5�v����K?���?-���2n��N�<Z��=)�^��&?�I4? k[�}�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��G��<��K>*4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��VS��GB�>�e!?���>�Ү=� ?�#?�k>NQ�>\6E��,��O�E�6`�>>��>X�?��~?r�?R乾= 3��Ⓙ�ʡ��[��AN>�x?�\?L9�>R���q���MX��G�=X�����?�Cg?ο㽒�?��?u�??�WA?��e>9@�޽׾ ������>Q_#?�6��@��\%�ـ�*�?��?���>�����Ͻ>:k�����S���(?EX?�$?����_��L����<}Nt�p�%�]��;�	����>��>� ����=��>�C�=�w�ջ?��b�^�=���>X��=s�'�c䧽d�6?n�*��^h���
>@�d���I����>�tP>�����T?w.*�Ks�&۳����T����0�?�j�?�[�?f3?��>]���H?��~?`�?��>�����ƾs�c=~������*
�X�=�`�>�D�<�Z¾u��������J������GKj��?+��>�1?��?7�6>�4�>П���l=���Ҿ��\�0���]�î��;�����{y�R#��0���z� ��>�ӎ���>�\
?_,>:k�>h��>�?��}�>wR>�yd>AG�>��;>� >���<�^�����cI?�#��k+�j!�h�Z��9P?� ^?8��>�؉<\߆�*����^"?��?�k�?Z��=�J����e?���>
&W�Y%?va�=�6;��)>���G����;�!�$=�RI>�>�uqZ���g�o��D=�>��%?�'<H��7>�D���=�>Zp�?�<4?Δ��J�����hO���"%�hd/>)1���cľ���RbZ�*�"�s�g�{�6�e��a�Q�/?{�?%�����0Ⱦ}�1��O��-�=sg?2��>c?��^>\Ժ���$]��D)��w����>�|?*m�>�I?�<?�wP?�mL?���>�b�>�9���X�> ��;�>���>�9?b�-?`:0?�?s+?%c>e������}ؾ�?��?�H?�?%�?�ᅾ�:ý�=��5uh�_�y�eu��²�=�	�<_�׽��u�ˣT=��S>��-?9u�ّ#�j!�!̃=�u�?�w�>�?��
;��>�@C?O?}�d=�g��C7]�Dó����>�S�?�M=}�=�GD>T�=6��=���<�>}<�<�$�;���=�U�������N�4b�;-/�=�a>���>js��Lnn�N[�>AY?�>�G�>fֆ�Y���_���k�={:a>��R>q�(>,Nپ脉�#u���i��{>���?䖳?Ӑ�=�z�=@�=筠�w@��K3�C$��j5�<es?1�!?4�W?��?;?:�"?	�>*F�I$�������Ӹ?:\+?F�>��U�ʾ���I�3��?��?KAa��2��)���¾h�ҽo
>n�.��~�����C��y�\w�r�� g�?*�?2�B��}6���羋Ƙ�����Y�C?rZ�>!|�>3�>��)��Xg�jF���;>��>=R?(�>ѝR?v@?6�[?o�U>%l7�r����������<��,>��<?l=?�ߍ?�Hs?X>�>�>:�3��'��~����D5����� �=�oR>��>��>���>��=E�ֽ�О���:��\�=�S[>���>��>e��>=s�>�<^�L?��>n���G4�������ܑ���p�m?�a�?1�,?,�=���OCU�5������>k�?ְ?��5?He���5�=T�<�M����T�J^�>�ٗ>���>:�8=>��=��=�x�>�>v�*�@0 �٨)��$��C�?T�8?Ll,=��ſ@om�MVu�����������GZ�?�i��c��=yW��܇�����S�r��c���W���ޟ��B�{�% ?�߂=<�>���=���<ğ�����<j�+=j̆<'�F=B�@�g@�<3�E��S��y���R�cW<;DJ=��@;��Ⱦi�}?W�V?ni8?�Q?��1>Z��=q����q>���y�?ܼ6>R�ֽO����m&��1��ߪ���^Ҿ�\ھY�����Lj�=����B��=��>��>�Q=o�=��$=]��=��;D��A~�=��=���=uU�=��>>W�>(qr?y�_�q���7$�S=���?�%�>J�=�����!1?盌=ԏ������|���̉?!.�?S)�?��?�@��&sc>��G����J�ս�>C,>=� ��>z>��r>��>�38����=&��?0��?�]a?|�z��W̿�B>�Y5>UR>v�R��P1��P`�@oa��5W���!?�;���˾n�>(u�=��ܾ�ZǾ>_0=v�4>�DY=0��[�9��=.c}���==.,u=�^�>)D>�D�=㵽�;�=�BS=~
�=1�O>��ͻ�+D�)�&���2=�_�=��c>.T%>��>�;?b?/?�Bd?4��>!lz��b̾�ֿ����>���=\��>f�[=R�%>
��>�:?�E?Y�M?;"�>��Z=�>[%�>�2,��k��羣���i �<��?�e�?���>�ZB��W�Sq�}=<��15?� 0?��?���>�U����8Y&���.�&�����4��+=�mr��QU�N���Km�6�㽱�=�p�>���>��>6Ty>�9>��N>��>��>�6�<�p�=Dጻ���<� �����=�����<�vżm����u&�T�+�6���_�;��;0�]<���;�y=M��>��,>���>�z>r��z�W>�窾1~e��� >�x޾��B��S^�[�d�����`����e>rK	>�"�5����M�>$�~>Q$F>V�?D�}?�!�=uW��۫���ܗ��Q@������={��=�ǅ�h�G��p�%�S���ݾ_��>Qߎ>�>n�l>�,�5#?�d�w=��3b5�p�>u|��9��.)��9q�@������Zi��eҺ�D?�F��G��=I"~?�I?D�?���>	����ؾ�:0>�H����=g��*q�i����?'?��>�쾝�D��U̾�����ַ>�H��P�S�����0�F��r������>rΪ�<�о�3�
`���폿эB���r�JȺ>v�O?��?��b��H���-O��������o?�cg?�/�>A?([?"-���j�V��&d�=v�n?��?e;�?�@>YD�=�x��Z��>��?z#�?&]�?��q?��9�i��>iQ�;�%>ҿ��˸�=�>J�=��=��?�?�
?��Y	��2�!��B7_���<��=���>i��>��t>#��=6zP=�O�=�$Q>�Ν>���>�g>0x�>���>*����u	��	(?�P�=�j�>�30?��z>��3=���� =M�I��@�Y�)��๽��۔�<%�R�/=��Ἲx�>2@ǿ���?�T>d���`?�i���&���Z>�kQ>�ֽ�W�>�FH>6ay>�$�>_g�>��>ce�>�*>2	��O��=���V���=d�7�S����pϝ>�!��e���Ӿ�s��ѳ�wz־�=j�<����%���o=���?���^X��q� ����t?*�>|?�N�u1�Җ>;?��g>G����-��-���nv��o��?�l�?��r>|a�>�S?��?��7���I�QU�!q�Y:���`�]�儍��Ԅ��}�C�o��b?�}?��C?�黤�g>2��?��$��T����>,�+��-7��7=G��>���G�z��徎׻�m �>O>ds?i`�?��?W�;���v�Xj)>L�9?�1?�=t?��0?)�:?[����"?��5>?"
?u�3?��/?��
?�p3>��=����v%=�␽����jDҽ0�ϽѰ���)=5p=�.:K�><��=L��<�ۼ��ּ�n��0�����<��8=��=���=3�>�\?�A�>ߔ�>�*7?�k%���4�[���&A+?c=�,��퍾�1����辙>3l?�	�?�aW?*�N> %@���7�m� >g{�>9�$>$�R>b��> ����<�xZ=�� >��>Ѣ=1h���w����a閾���<ݾ>��>Է>�oػ���>N;���ξ�*�>�ϾO���ح�׏����P�����s�$?W�|?TU?��>Pv�ݢw��%����?��;?#]?�߉?�E�>�ƾ�8e3�d{h�̔���P>��>;��˘�f���{���V�&�:����l�����\>�B�D]�K�k�C�G�����HM=\����=����ܾ�����f�=Á>�E���:"��5���z����J?���=s���=W��Ѹ��>��>PZ�>6�>�A�|��	@��ծ��/�=�~�>2>�9ȼ$m󾛿G�x=��u�>�eG?�g?a�?Yhb��Zq���>���k`���l#��8?�F�>~x?��=>� �=M���C��?d�DwD����>��>i� ��*G��������7%�s�>��?�O3>@�?�L?�3
?�
]?N�?2�>3��>���*��)�&?t@�?%��=RxŽpSG��5���A�GI�>L ?���л�>��?WW?$�#?$�J?��?���=����#7���>�V�>ĚW��
��'E`>ݠJ?'[�>��U?]��?��G>�[2�0S��v^,�R�=3?>�5?�_%?�d?�3�>l��>����_f�=�L�>W�b?w9�?!�o?c��=Z�?�!2>��>7�=[��>T�>��?T=O?1�s?��J?���>�<N6��O����s���N��g�;�H<��y=��5Lt��?���<Ҁ�;�[���I��U�OD�������;���>~��>_����f�>��E���={#>�M���[���Ͻ�ۈ=8�^>��?K�`>����{�!=�:�>�u�>B����p?��>#�?��=P%��z�����{Y�>��k?`�8==�o�����Hq��K���?j��?�ԅ��~���b?�]?�^�R=���þz�b�h����O?d�
?D�G���>�~?�q?���>��e��8n�M��<b�!�j�ʶ=Oo�>nW�^�d��<�>��7?SP�>��b>5$�=�p۾��w�g��L?�?���?���?�,*>��n��1�d�������Z?�[�>���x="?p��ξ1j��+���{��鳾���ᘾX<��1z��W���B�V��=�T?�Bs?��n?��\?����e�b���\��3��Z�S�] �yi�Q�D���E�'PE��o��F�� ���s���3B=ݬ��U�-��z�?(�%?�ѽ�b�>'g���y��jrȾ��@>����U3�k�[�\���&�=s�=��M���7�GM����?� �>F��>C^;?+�G��f6�#3B�3@1����r|�=Ⱥ�>c��>���>Kö�R������־�\��7��^�g>&�s?^SZ?��s?���=�Xa��E��C��ԯb>�?u�Ǽ=��4>e�>���a==��׾oB�q�����F�]֛�JI-�n+�=Z�G?a=NԦ>��?�8?�P�K^⾙�~��%%� >i��N>Z�?R�>���<zd�=x�^��>��l?ܹ�>��>�a���W!���{���ɽ���>��>���>��o>�G,�V
\�Va���~���(9���=��h?n{���`�_��>y�Q?�/�:́J<���>�dv���!���
(��4>�?i��=��;> ržf�.w{�A+��im)?{^?�L���*�$�>�`!?-f�>�>�o�?��>��þо~:5a?��^?�I?*a@?���>�#-=5�����Ƚ��&�&W)=p��>�oZ>�l='~�=S(�_�[���� ;= e�=�����?<���]+S<�� =-'1>vۿ7�K���ܾ����E����4������͊��p$��д�ܤ�����`g���/��PP���l�37��֠t���?��?��+ꊾt���G�2����D�>�k��O���*���J �ǣ��6M��-��c{"���S�#�j�ݞc��?ֲ��G1Ŀ�֡�O�˾�0?�<?�AL?f����7���F��N�<�����νc��d�����Ͽx���ҞW?b��>kbǾi��ձ ?��d=��#>�N> ��1g����=�Z�>̃8?X?/f;���¿�����=O��?S	@4D?�)����VE��"�>ϔ/?��s>A�߽�j��FT�>|r�?&Յ?����g�J�a���W	f?ބ�=dn��˻��=���=�#�=����&>�}>I&��E��(�?�Wt>��">j�_��ȴ=��\�_�+��~>�O%�W��3Մ?"{\�sf���/��T���T>��T?�*�>d;�=��,?K7H�_}Ͽ�\��*a?�0�?���?=�(?�ڿ��ؚ>��ܾ��M?fD6?���>�d&�%�t�܅�=�:����y���&V�=��=4��>�>ڂ,�Ӌ���O��H����=!(���&Ŀ�x1�Ϗ?��
T>ϲL>�9����)0����ؾ 䋾��澑^[�;�S=3�>F�>a;�=\Q�=K:<��\?
�? ��=3��=�I��#����3�g2}�����"����P��Kھ�_�*x���6��#�ub1��/��c˾�J?�^�n=lR�}����(�73]��B��,?W�>�ݾO#L�YἿ�վld��r���y��Ӿa	4�	n��ş?�"D?ᢄ�H�U��7��O$�/���
6N?L��L�G���b��=�x#�"�<A��>�j�=��=W4�=N���0?�*?��������>���3A=��,?��>_f�<g0�>܋"?&���O��n2G>[>v�>���>�>b<����P�?=LU?n��#���g�>�g���s�r�D=�[>k�:�@pǼd<> F�<Dh��	�4�H�����~<��S?�'�=m�L�
7M�F�����r>"�=dTO?j��>�ى>o1{?� ?�{>4o$�h}j�ӫþ��h>uog?�?�f>]��Ry/����`E?��?_-�>�G��c���&.��5��m?X?�#�>�/a>��?���_�]Ѿ�|�>S�v?��]�@�������U�=ݤ>{`�>&��>��7�v�>�V>?�M&�w>��We��7�3�G�?�@/r�?<v<���f�=�l?�6�>�M�xpǾճ���U���v=�>L����u��& ��1.��7?�y�?�E�>��S���X{=đ����?%<�?�1���)ν�)/�5��3��X5�<�e=��e��+�[^7����[� �
���>�h�>@@sjs���>Q��ѿ&��@4��i��F�ԽoV�> Y�>�p�=�U���B���p��hM���t��&��h��>��>0璽c���?={��*;�A��>@|	�~/�>�BQ�AI�������R)<�>�>�g�>���>��nj��M��?2����ο�ʞ�
x���X?�ў?23�?��?$aZ<�t�7^|�n�!QF?�r?�.Z?E���Y�v�+��h??����^�$ 9�YXB�~>&�2?��>
�-�JD�=��t>t^�>�&>7l�����p���V˾�r�?�w�?k�w��>܄�?�D5?ܓ�^!���̛�!�$�N�&;��.?O�;>�ZѾcg��rH�E���,��>0&?S�4�`��]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�1�> �?�+�=LT�>���=R찾 +���$>o5�=��=��d?w�M?��>�
�=$�7�T/���F�C�Q�F��C�v�>�a?�CL?KYa>�z����1�!�}-ν��/�1��?�0����[�4>�=>E�>�D���Ҿs?�����׿}p���h���'?djw>���>��[��_u=��G?��>/��|���׭��i㷽��?#��?�?��Ҿ�|��q=���>o®>��i<��u-����J>�.9?����"ag�� d>ڞ�?��@�k�?#�N���	?I����Uv�����7�[F�=w20?y[羑��>�`?
^�<%h�B��'�y�B�>�Ӭ?��?H��>Іi?,�g�6�:�/sx�U�>y?q?mkx��g�=Q>�� ?m��+W!��czU?DK@%�	@�T?ۓ����,}���Ჾb����>3+>��>��s����=�V >k�������R=oy�>�8�>���>v[g>�R�=��=�B��P'-�|1���B���a����:Y!�������⦾P������Q�ݾ|�8�@r,��VC�!��;_y��Jd���`=*�`?�q�?��?���>���v�G�����q�<5<}���f>xf�>0� ?J�a?Z"E>2��7m�kX���Uu�.�U�1�?��=�ޭ>�`�>"s2?�%�:o�=���>�q�=��=�&?�Sx=�҆<��^=OSY>[0�>8)?D�%>�s>tƳ������a�r9k��\�����?�m���RR����`ڞ���þ�`�={�)?`>⭒�N�Ͽ�����I?��������0�h>�,?/�T?�� >g%��ӏ_�F>]3�tXv�Q��=���j#w���-���?>�?�}f>a#u>ѕ3��[8�ۻP��u���t|>�6?j���+r9�\�u��H�Ԁݾ!M>U��>�hD�0m������� Oi�~�{=&t:?˂?�ͳ�밾��u�C��LR>rj\>H�=�p�=scM>�Pc�]�ƽ�	H��a.=���=��^>��
?��=Ls漰�>�.��Xq��m�>��>�w�=Ln5?�NA?����5�<�U;��z�~�=�?��@>�}S>��8���R<� �>^E�>GS<��A�0����=�@�>k��6��ah��ɩ=����G*>�U�>�	���Y��g3<�~?���%䈿��0e���lD?X+?� �=J�F<��"�@ ���H��F�?q�@m�?��	��V�@�?�@�?%��l��=}�>׫>�ξ�L��?��Ž4Ǣ�Ȕ	�4)#�eS�?��?��/�Uʋ�3l�u6>�^%?��Ӿϝ�>)��j��,|�T|��e �7O�>��A?�Ծ��8�X�����>�?����eF���ƿT�c����>���?�?��d�����V[I�vM?��?�sK?�8>vz�<2/����>1P,?�K?s�>QQ����?("�?�e�?<�3>�-�?�τ?�*�>�<f>�Y9��ԿC�����>�70>�_����^>=���%U�����)b���M�k[Y��X ��B�=���>ʌ��Y¾���=��Ͻ����|�B��8"? ,�>�W�=�/w>ߗ@?��?�{>H�<	/=k���ѹ�m�K?���?����2n��Q�<Ꞝ=�^��&?pI4?Aj[���Ͼ�ը>�\?V?�[?d�>R��H>��F迿C~��r��<9�K>M4�>YH�>�#���GK>��Ծ�5D�bp�>�ϗ>����?ھ3-��_E��:B�>�e!?���>�Ү=�#?��$?|�>3��>o�/��ҏ��,=��M�>7�>I�?J�u?v�
?�§��+��ʌ��k����b�� `>�(s?�s?Tք>k�������s�e�::����d�c�?��X?������ ?��?�ZP?��??�+>�6���ɾ�{�	�>��!?,��$�A���%����?�?��>����ҽ)ͼ��1����? �[?��%?�%�.�`��¾<��<os�NP����;�6�A�> I>ш�u��=٭>PZ�=�n��6�7�\<ִ�=[֓>��=��6�hk����(?�(=���V�a>��O���n��e>}~��2U>n�]?��R�{�h��b���w��Q��{B�?�;�?���?1�����k�g,o?�h�?��B?<K�>b�ɾ������)���Ⱦ�y*> ��O�>�]x>}n6<,�ľ ���}���C����ν�YM���?S�>2�?��
?�=Y}�>,�;��"�2�������V�?�9�EV.�ۭ�9���?c�9�Xu8�b�Gƈ���>J���ԑ>��?��5>VZ>�ï>��xu�>�43>@>%�>��u>V�T>�P"=�^�<�=_D?���i���M77��WݾXp$?�R�?6\D?�x"�ʀ��rԾ/]:?��?��?�1�>��]���6��j�>��%?�ܗ�ն? eŽ��=嘽�?���r��vsK��� =�>Yר���E� oY�9�/��T�>�7�>)���B���;�N$����w=�̄?�B(?m�(�oBQ��Hn���W���R����X�k��n���$�R�o�eh��!��._��Tm(�(�/=<�*?6f�?��]�����y�j��?��3k><!�>�H�>��>��I>v��0�=�]�z�'� ΁����>�}{?� �>#�I?X/<?��P?m]L?��>�٨>L^��<��>^9�;Rw�>ua�>m'9?��-?Z^0?^�?+?q+b>`�������Q�ؾ�?�d?�?"?6�?3ᅾ��ý[���՝h��&y�P$����=��<Q�׽5�u���U=	�T>��-?O.h����������,?Wu?ju ?�a��V�^�|��>�jH?��H?���>�Iž8�n��M/��j�>��m?��ǽ8o�<�>>�j->�����m<FZ�=��<�Y���z=�?�����=�E�=�	�>�q�=��bm���^-<�����z�>D�?T��>}E�> 3��F� ����(�=�yY>S>��>�\پ����$����g���y>#|�?�~�?��e=+��=<��=fS���/�����/��^��<{~?�C#?�`T?���?�=?�`#?�>M)�eI���^��4��J�?�m?�@�>	���4Ҿ$����*�?���>hpg�rZ�+8�p�޾�\޽���=j�?�+(���X�A�J7=d����\��?�e�?��@���<�����"�������eJ?���>>E�>��?σ�5�X�4'�Js|>��?��S?B0�>��d? ��?+%W?���>��F�>��ƞ���h>6<h>=�?��z?s.�?�q?q�>W">a�'�����ɼhY1��.����}=Wx>��/>)��>3�>M�=Vc"� ��<�)I���=?+o>�?���>��>�~�>W/e<�0E?⃰>��$|����|���䲉�xFk?�?'?��7>2�&�p�D�g�����>�̹?v��?9)L?}Ɓ���=fT^�0Ɏ�A���fO�>�$}�u�>��佽�>�t���C>$�C>�T�?����ﾏ�>��'?~�a?g�Ҿ��ſ�q��/q�\K����s<��|d�����T�[�*B�='Ę��%�I���1\�Y���
���a��2���|�H'�>P�=#3�=]A�=Ә�<Kg̼���<�E=V-�<��=��p�-g<��:�PL�����f�K��<<%E=�ֻ��־.̀?��E?Z�,?�HB?iW >M�9>�f<��L>�*=�M�>0?�=��i��|��T��HI��Z���ѾY����|_�er��~}q>ßཱིF�=�":>�~�=�<��=��=��/>w�޼+�V=?��=X>�N>�q�=�� >\!�>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?Ati��d�>M���㎽�q�=K����=2>r��=y�2�T��>��J>���K��E����4�?��@��??�ዿТϿ5a/>�A:>�>�DR�M�0�*p]�@�b�]<V��#"?g;�̾��>��=�'ܾfXž_� =]�1>��o=���rZ�旙=q�w��\==�Xf=���>n�F>m��=;'��?��=�<H=���=�DP>�{���$�ij)���3=�8�=aod>�n%>��>JV?b�+?&�e?J�>
0H�z�ľ:���u
�>i�:>�׭>�;=Cu.>�ܭ>�!3?�@?�B?�ޥ>�˺==�>q��>��)��bl�ݺ��,ؑ��ƪ<�f�?��?ǲ>Ǽ�=�O�s����>�0���t"?�7?��?z>!�����Y�uC���{>/����!��� ~�0F�kZM�4�ͽ�њ=���>u�G?���>�.>�3<j}
=I��>�>�ɋ��9�~�*=M�=���s>�ֽU�O�=���5���O=A8�����=�4>�Z'���>>=���=6�?XPd>�N?:-$>۠�u�S>z<�ۀ5���>J-��9�N򃿇r�����G鼢,�>�>�ڗ��雿��>ۼf=ز�=5��?!��?��N>��8�m%����ꑠ�T$����Z=�57>��T��EQ��`���o�+-�/��>���>��>��l>�,��?���w=����a5���>w��W��� ��)q��;������i���κM�D?�?����=�~?�I?7ݏ?��>�G��h�ؾ�N0>m!����=���'q�������?;'?��>���D�6"��x@̽��<Zކ�࢒������h	�3�y;e�V��x'>��O����.|��$�I��f5c��P��;P�>�/G?3��?∾Q�n�Z+����4����>�y?u1?�y'?��b?�&=��m�f�O���.>�D?,�?�p�?�|�=�O�=g�����>��?`�?�(�?޲o?6,+�Lv�>m��<έ>tQ����=�>���=���=�O?ko?��
?������3��
����
^��6$=��=��>��>Γv>�9�=�j�=���=�e>;�>g�>��g>�G�>��>
S��Qﾐ�-?+c>��>u�!?��>��*�b-ɽ�ؙ=��]���e��v�罙�L��ӵ=��<�J(=�h�D��>ÿ5p�?�.G>��<�?������[��<`>�o�=,t�����>�T>��>9��>��>V��=��]>U��=�����L=>37��*�����3��v�����=#��3�c�i��㮾B����hѾ
Z־��C��Ē� 6�-�<n��?D�ؼ�a��67�R�3�r�>YMg>8_
?�@ž�>���=i�>��?q�־�J��.���\Ҿ'L�?��?>c>L,�>ܧW?�?W�1��2��VZ�Tu��A�(�d��`�F؍������
��Կ�e�_?M�x?<_A?h��<3z>��?'�%�׏��I�> �.�W;��=;=[�>i��9w`�ŮӾМþ���*=F>��o?'�?C?�tV��!f�9@(> �:? �0?�Rt?�V1?c;?͝�*�#?[�6>ٛ?4�?v�5?��.?��
?�0>p��=l��s*=���ո���'ҽ��˽��o�2=�~=1�A��	<�=��<��ۼC2Ѽb�;�����'�<��:=rˣ=}��=P٣>v]Y?��>	T�>��6??/�<G2��Z��z�0?|�P=�끾�����඾����n�>7q?��?H[?�A=>�s@�#�C��<>�]�>�>]�D>6I�>N���z4�rs=��>Y�>p�=г��;�k&�n���:$�<��&>�z�>Y�|>�=���i(>P��Hz�H'd>�3R�m�����S���G���1�Ww�w��>�K?�?�8�=�g����f�U)?\�<?�<M?Y�?�'�=q�۾)�9�h�J�x��ҟ>|ձ<�������� ��b�:�fS:@�r>�=��{B����a>�����߾�Ro��J�X����~=.��	%=ښ�A־x�u�l��=Ht>�[��{c"��Օ��_��dK?�To=x��+�A�{����v>'��>�Ү>=�N�CM��(>�?��F0�=��>R�?>GӼF���F�; �$Ky>�F?=΀?&��?�E���w��HG�S�
�I���H�>��
?�AU>4ؙ>�K>�w�=��پc2,��>�@A7��?��f>!�"�5(O��7��c���]�L��>~�?*�|>Y\ ?��'?��?V:?Ow?Z�>�p\>�0<��g��A&?��?��=l�Խ��T�� 9�[F����>�)?��B���>~�?��?��&?��Q?%�?^�>`� �`C@�U��>�X�>��W�gb��S�_>U�J?���>n=Y?�ԃ?1�=>��5�1ꢾ�Щ�hT�=�>i�2?�5#?��?��>��>�@����o=͓�>�^a?���?��k?��=��?h#/>�>�T�=���>N�>�?�`K?ktr?΀E?l��>]X�<!���(%ǽa������)�ڻ 	b;�Dy=Ze&�e�J�_���v<�ߞ���2��i��p�����x�����-#�>��=�(������4���۞�=���;Kٽ�þ�V�=��=��R>୼>l�%=�@ʼ.V�=�>�>��?*�E�-?���>�)4?��-�>�l�����㽨¨>x�C?��=*u�.!��Mo���<7�j?]X?O�T�`���J�b?��]?Lh��=���þD�b����b�O?A�
?p�G��>��~?^�q?3��>3�e�#:n� ���Cb���j�1Ѷ=Br�>>X�M�d��?�>��7?�N�>�b>Y%�=�u۾�w��q��t?{�?�?���?�**>g�n�O4��}���l��f_?=��>+?%�i�?�$�<�B����s�����D��{��g����:��+с���p��@��WN�p�?y?�߀?4�V?�H���W��y�Iu�� I2��������;9�ed5���Q�e����0������پ@V��@��@ �]�?�d*?��ý�q�>�T��J9�pǾ�vt>�ެ���0���O=�<>�8M=���=�_�"g�c�ľ�'?m��>���>��3?$=M��44�Y:��1���Ǿ�u�=ڊ>��>Fi�>�����k����2�ܾ]����۽d�b>��{?I��?븆?K�='�)��V����7����=�{��9>$s�<��*>	`������n�,���S��!q�l~�3���_&��x�tG6?=��>P��=3��?��?<X�����<��}��1\��a��> 6�?�m�>E�<>@A�>�;��D�>Z3l?+M�>}��>z���� �4�|��U̽Q&�>��>��>�yl>�+�ƹ[�v����⍿�_8����=jRh?o��Nuc��<�> �Q?+1��W&<>\�$0!�5g�I�(�Tn>�?46�=ɤ=>rƾ�f�5Az��C��.v)?8�?�Ғ�4x*�r`~>�"?�!�>�c�>��?��>��¾�蚹�}?��^?��I?�A?���>��=�Ů�F�ǽ��&���)=�&�>AZ><i=���=�����\�����dE=�I�=}�Լ;/����<�ǣ� �T<���<�3>1Mݿy�H���޾ѡ�&���r�n��7$�����&�h*���Ř��ek����r�-�.�S���u�=ڊ���q�a4�?�J�?�����񑛿��~��S�@^�>�z��2��#��[�dD���^ܾ"i���	!��uR��)g�J�]�^@'?h�����ǿ񍡿��ܾ%�?gI ?��y?n�y"�HW8�}o >��<џ��<�ؒ����οE�����^?���>Q]���� �>֠�>5�X>�q>@^��.�����<�:?��-?�C�>�r��uɿ������<���?��@�.?�}M�M��rm����>xZC?���>{�X��}��W����:?=�?/0�?��g�Y�5�u���9�9?+eq>�e&��$>=��>uA>�>�����=��>��!>�Ӌ�1"�<N૽ki�>��A\4�ٛ�=¶��۝�=o �>���<��`K~?�B0�9I���>>w�Й�M�Q?}�>��3=1*?��a���ؿP�j���v?�� @��?
+G?����x<>�y�{�Y?��*?�ڄ>��꾫ja�`5�>E��0E�f�ɾS�l����=��?�q�>n�S��⾪��6��,=�[�ƿ��$�xj�y�=s����[�j�+��G�T�m6��;�o��}�q�i=��=S�Q>~Y�>P�V>Y�Y>x^W?�k?�\�>ܱ>(,��y���ξ�?�y.��C��ʪ����ޣ��ƭ߾�	�s��C����ɾ�P}�T�<?�Y�R����7��rf�E~"�Z�@?�[	>9L�,�A�Š6�*뇾���� �?����`�9�5�^� )�?9�,?����CI���4�Ol��u�=l
�?d����&j־j�<�x�==:3=���>+쐻�v�>+��;�J
,?4?x�ľ����I>D���Q���(?��?�t�<-0�>�#?��)����#�>��H>�:�>�5�>�0J>0����
��8I?N�Y?��d�ۏ��'�|>?���v��G,>���=� R�a��C�@>��=Z"���'<�܆��*ֻ>�??���=X�6�������2�����\? �? �v>L�q?�&?�R�=����b�!�����="�?��}?��'>A1A�߈��K�ƾ�X4?���?!�>KH�=��̀j�w��O�M?G4e?���>x�>�T��#���jܾ-�>��~?^G\�o]����¾Sf���}>���>���>�����>�($?�B�:v���н����Tߛ?*@��?{���v'�^ =X-�>I,?Er�\����j=票��W>�j�>��Tb�cAC�ὺ�R=?@v|?oS*?���-�>���V=xK�UΫ?T��?�rb�z��}�o�s�ߞ�����<�}�������p�������7�fӺ��
��ݿ�K�ֽ��>nb@
�5��>�����ֿ�}ҿ�>��X��\�7���?���>̽�ڢ�c��炿L�N���W�P����X�>��>�K��������{�\~;��ߞ����>g����>�S�J��X퟾Wu5<U�>u��>�݆>�?������ұ�?}-���.ο���G��K�X?X�?�b�?EV?C+<<]"w��
|����&$G?�ws?\#Z?�$��Q]��5�P:j?4���K`���4�W�C��]U>�1?*r�>��+��bh=��>�C�>FZ>	�.��Ŀ����cm��/��?h�?{�hR�>��?�,?D���������SK)�u�:��A?�|2>������!��<�����S
?�`0?9�������_?ŕa���p���-���ƽAϡ>�0�6c\�Y��Ș�[e�
��sQy����?�^�?��?&����"��1%?t�>p���J4Ǿ���<u��>b#�>�=N>d�_�a�u>!���:��e	>��?�~�?�l?m���@����=>��}?v$�>��?�n�=�a�>Bd�=�
-��k#>�"�=��>��?��M?�K�>�W�=��8��/�'[F��GR�*$�+�C�0�>s�a?�L?WKb>���� 2��!�duͽ%c1�#P��W@���,���߽:(5>��=>:>f�D��Ӿ��?<3�e{Կ�蘿@qR���=?V�>7L
?��
��ۙ�-c���s?ܙ�>�������ȇ���ec�?���?��?��Ծ�V�p�=���>m��>Y�1Xܽ�~Y���4>�]2?�Ӓ�$Tu�f܃��ԁ>��?p��?I��?�_�?�X���v��na��M�;h�1=��3?5h߾:�>���>1I=��i�D���SO�
��>9�?#_�?�>�T?�#p�g_�{6->�|Y>��6?���>�ɑ��9ɾo��>��>Gt�i蝿0�\y?��@b�@���?�v���6޿:����B�����td�=��=9�>�Ž���=m�3<X�;
����>T��>�U>�
p>e�>��9>�	�=_����|@Ϳ�K���f��p9����l� F������ �ݬ��S릾���PM���q�Ѿ���Ᵹ��z��2^?�OL?��z?�,?����F6>�c��n��z�<�lm��Η;�w�>M+g?��;?���>d:��l�\v����:J�#��>|D�<I�>(�u>I�x>��<���>zT>���>E! >xÆ=�J�<\6�=n
�>�%�>��>k��>~�>��>w\���ݯ�
�o�����(A�����?}䣾pO�����I5���>����=4�*?�
�=�^���Q˿�z��ܵJ?y��՘��ֽ���=�7-?"�S?��>����?1">�7� ,e����=�X��9�z�;Z#�whC>o+?��C=��P>��8�+.���w���о�-�>��M?�׾A�k�hCe��$?��ڜ��%>�Y�>����q4��m��(^�V?��-=�Q6?.u2?����pƙ���'��;oH<>H��> �l>(��=���=[K-��֍������G�=��>��>/d?���=��-;&r�>k���ӄ��H>nZ>�k�>�6?��1?��&�r�u�}��M-��/�>��?('�>O�>��T��,7>��>|>��5���(���������=�B�=��������O=��b��2>)�;R8ͽ޵t�V�<�~?���(䈿��8e���lD?W+? �=a�F<��"�B ���H��F�?q�@m�?��	�ߢV�B�?�@�?��"��=}�>�֫>�ξ��L��?��Ž8Ǣ�ʔ	�=)#�iS�?��?��/�Zʋ�7l��6>�^%?��Ӿ�l>�mʾ�$��6~f��I�����=ٲ(?��X?;Q�v�d�
�<�1?��?4�����z��sĿ�?j��?�ݼ?� �?K"��+ȏ��g�?jJ�?�??v�\>��վ(���8	=�cm?{�g?�;p>Sg&���k���"?�ՙ?�AL?m��=/�?E@�?���>}��=u�%�辿�\���]>$�u>B)j>�;=���ϫ7�v ��z��n��-O��Z�=�k>v��>���=#Ȯ��Z}�6�R<�4˾�����?@�H>�>���>?E��>a�r>4�<`ҽF�5�v����K?���?-���2n��N�<Z��=)�^��&?�I4? k[�}�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��G��<��K>*4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��VS��GB�>�e!?���>�Ү=� ?�#?�k>NQ�>\6E��,��O�E�6`�>>��>X�?��~?r�?R乾= 3��Ⓙ�ʡ��[��AN>�x?�\?L9�>R���q���MX��G�=X�����?�Cg?ο㽒�?��?u�??�WA?��e>9@�޽׾ ������>Q_#?�6��@��\%�ـ�*�?��?���>�����Ͻ>:k�����S���(?EX?�$?����_��L����<}Nt�p�%�]��;�	����>��>� ����=��>�C�=�w�ջ?��b�^�=���>X��=s�'�c䧽d�6?n�*��^h���
>@�d���I����>�tP>�����T?w.*�Ks�&۳����T����0�?�j�?�[�?f3?��>]���H?��~?`�?��>�����ƾs�c=~������*
�X�=�`�>�D�<�Z¾u��������J������GKj��?+��>�1?��?7�6>�4�>П���l=���Ҿ��\�0���]�î��;�����{y�R#��0���z� ��>�ӎ���>�\
?_,>:k�>h��>�?��}�>wR>�yd>AG�>��;>� >���<�^�����cI?�#��k+�j!�h�Z��9P?� ^?8��>�؉<\߆�*����^"?��?�k�?Z��=�J����e?���>
&W�Y%?va�=�6;��)>���G����;�!�$=�RI>�>�uqZ���g�o��D=�>��%?�'<H��7>�D���=�>Zp�?�<4?Δ��J�����hO���"%�hd/>)1���cľ���RbZ�*�"�s�g�{�6�e��a�Q�/?{�?%�����0Ⱦ}�1��O��-�=sg?2��>c?��^>\Ժ���$]��D)��w����>�|?*m�>�I?�<?�wP?�mL?���>�b�>�9���X�> ��;�>���>�9?b�-?`:0?�?s+?%c>e������}ؾ�?��?�H?�?%�?�ᅾ�:ý�=��5uh�_�y�eu��²�=�	�<_�׽��u�ˣT=��S>��-?9u�ّ#�j!�!̃=�u�?�w�>�?��
;��>�@C?O?}�d=�g��C7]�Dó����>�S�?�M=}�=�GD>T�=6��=���<�>}<�<�$�;���=�U�������N�4b�;-/�=�a>���>js��Lnn�N[�>AY?�>�G�>fֆ�Y���_���k�={:a>��R>q�(>,Nپ脉�#u���i��{>���?䖳?Ӑ�=�z�=@�=筠�w@��K3�C$��j5�<es?1�!?4�W?��?;?:�"?	�>*F�I$�������Ӹ?:\+?F�>��U�ʾ���I�3��?��?KAa��2��)���¾h�ҽo
>n�.��~�����C��y�\w�r�� g�?*�?2�B��}6���羋Ƙ�����Y�C?rZ�>!|�>3�>��)��Xg�jF���;>��>=R?(�>ѝR?v@?6�[?o�U>%l7�r����������<��,>��<?l=?�ߍ?�Hs?X>�>�>:�3��'��~����D5����� �=�oR>��>��>���>��=E�ֽ�О���:��\�=�S[>���>��>e��>=s�>�<^�L?��>n���G4�������ܑ���p�m?�a�?1�,?,�=���OCU�5������>k�?ְ?��5?He���5�=T�<�M����T�J^�>�ٗ>���>:�8=>��=��=�x�>�>v�*�@0 �٨)��$��C�?T�8?Ll,=��ſ@om�MVu�����������GZ�?�i��c��=yW��܇�����S�r��c���W���ޟ��B�{�% ?�߂=<�>���=���<ğ�����<j�+=j̆<'�F=B�@�g@�<3�E��S��y���R�cW<;DJ=��@;��Ⱦi�}?W�V?ni8?�Q?��1>Z��=q����q>���y�?ܼ6>R�ֽO����m&��1��ߪ���^Ҿ�\ھY�����Lj�=����B��=��>��>�Q=o�=��$=]��=��;D��A~�=��=���=uU�=��>>W�>(qr?y�_�q���7$�S=���?�%�>J�=�����!1?盌=ԏ������|���̉?!.�?S)�?��?�@��&sc>��G����J�ս�>C,>=� ��>z>��r>��>�38����=&��?0��?�]a?|�z��W̿�B>�Y5>UR>v�R��P1��P`�@oa��5W���!?�;���˾n�>(u�=��ܾ�ZǾ>_0=v�4>�DY=0��[�9��=.c}���==.,u=�^�>)D>�D�=㵽�;�=�BS=~
�=1�O>��ͻ�+D�)�&���2=�_�=��c>.T%>��>�;?b?/?�Bd?4��>!lz��b̾�ֿ����>���=\��>f�[=R�%>
��>�:?�E?Y�M?;"�>��Z=�>[%�>�2,��k��羣���i �<��?�e�?���>�ZB��W�Sq�}=<��15?� 0?��?���>�U����8Y&���.�&�����4��+=�mr��QU�N���Km�6�㽱�=�p�>���>��>6Ty>�9>��N>��>��>�6�<�p�=Dጻ���<� �����=�����<�vżm����u&�T�+�6���_�;��;0�]<���;�y=M��>��,>���>�z>r��z�W>�窾1~e��� >�x޾��B��S^�[�d�����`����e>rK	>�"�5����M�>$�~>Q$F>V�?D�}?�!�=uW��۫���ܗ��Q@������={��=�ǅ�h�G��p�%�S���ݾ_��>Qߎ>�>n�l>�,�5#?�d�w=��3b5�p�>u|��9��.)��9q�@������Zi��eҺ�D?�F��G��=I"~?�I?D�?���>	����ؾ�:0>�H����=g��*q�i����?'?��>�쾝�D��U̾�����ַ>�H��P�S�����0�F��r������>rΪ�<�о�3�
`���폿эB���r�JȺ>v�O?��?��b��H���-O��������o?�cg?�/�>A?([?"-���j�V��&d�=v�n?��?e;�?�@>YD�=�x��Z��>��?z#�?&]�?��q?��9�i��>iQ�;�%>ҿ��˸�=�>J�=��=��?�?�
?��Y	��2�!��B7_���<��=���>i��>��t>#��=6zP=�O�=�$Q>�Ν>���>�g>0x�>���>*����u	��	(?�P�=�j�>�30?��z>��3=���� =M�I��@�Y�)��๽��۔�<%�R�/=��Ἲx�>2@ǿ���?�T>d���`?�i���&���Z>�kQ>�ֽ�W�>�FH>6ay>�$�>_g�>��>ce�>�*>2	��O��=���V���=d�7�S����pϝ>�!��e���Ӿ�s��ѳ�wz־�=j�<����%���o=���?���^X��q� ����t?*�>|?�N�u1�Җ>;?��g>G����-��-���nv��o��?�l�?��r>|a�>�S?��?��7���I�QU�!q�Y:���`�]�儍��Ԅ��}�C�o��b?�}?��C?�黤�g>2��?��$��T����>,�+��-7��7=G��>���G�z��徎׻�m �>O>ds?i`�?��?W�;���v�Xj)>L�9?�1?�=t?��0?)�:?[����"?��5>?"
?u�3?��/?��
?�p3>��=����v%=�␽����jDҽ0�ϽѰ���)=5p=�.:K�><��=L��<�ۼ��ּ�n��0�����<��8=��=���=3�>�\?�A�>ߔ�>�*7?�k%���4�[���&A+?c=�,��퍾�1����辙>3l?�	�?�aW?*�N> %@���7�m� >g{�>9�$>$�R>b��> ����<�xZ=�� >��>Ѣ=1h���w����a閾���<ݾ>��>Է>�oػ���>N;���ξ�*�>�ϾO���ح�׏����P�����s�$?W�|?TU?��>Pv�ݢw��%����?��;?#]?�߉?�E�>�ƾ�8e3�d{h�̔���P>��>;��˘�f���{���V�&�:��������tGb>��
��ܾ��l�8TI��[�!�C=+��$�V=���վ
(����=z\>=G����Z�N���qJ?L�k=���V������R>Wޗ>�0�>��:��|��?��ӫ����=���>��<>���e��F��k��څ>�aE?Ŏc?�0�?�7m�:�t�e�E�C,�E��M�_�1d?2G�>�?f)>R��=���R*��a��J��`�>�	�>ߴ���I�*����Ą���>�K?�i>�"?d�S?6�?6)_?$�&?܈?���>ƪ��3鬾rE&?چ�?�-�=��Խ�T�d�8�*F�\��>�)?�ZB��̗>C~?%�?�&?�Q?��?�>s� ��5@����>HJ�>��W��\��_�_>եJ?���>g3Y?Nу?0�=>�s5��ۢ��ѩ�vd�=K>%�2?j##?��?���>m? �ƾ2��=�0�><�,?��x?y�? T�=~� ?�>���>Kyg=�>(�?�,?[wP?��m?�z ?���>�E�����Ȯν�g�RЅ����;�җ<.=�[�\���>���M8]=PPq����=��:VX��G��ć;�ϼ=c�>jo>�����?>�;ɾ��ͽt��>xg0>*�t���ս~r)�ʏ>�!�>�'?�E�>rP���I>}Lq>Fi�>Y����?�q�>�v+?���=��I���#���p�n9�>EIs?�1�=�uu�\��`�I1�>Qq�?t!�?�{8�u�
�6�b?��]?�g��=���þX�b�9�龙�O?��
?]�G���>��~?F�q?���>{�e��8n����m@b���j�Hն=Fq�>�X���d�!B�>�7?�L�>��b>�#�=u۾��w�8o���?^�?� �? ��?Q)*>�n�u2�}$�x��W9T?@��>R�o?	(x�_bž���e卾�[�Qy����������� ����lMǽ�J�=�B?�Yo?בr?2_?3����lf��2^������U��~�����uD��B��EC�#�q�?N��������DE=�y��m��l��?K�;?�	<���>!��&%��Ĥ�W�>�þ�����<��I�)>���=%m9������Ѿ�}
?Y�>��>V�4?��J�c Q�UL�Y�,�=4��}Ͱ>���>���>�:e> =��L����>��ק��f��<`���p>u?��p?ζ>?�>`��<���Q�4��=�������>�	_�0ݓ<����Yx]��䬾�(?��Tg������Hn�i�>a~!?ɡ�>P� =P�h?�&�>�"�����!�-�;�M����<�]3?Ft�>�Ar>hy>]�=�N �>��n?Q'�>Λ>a���,�C�����E��>��>oP?��p>��'�֦U�@ύ�� ���;:���=;zg?0݀�
�r�(�>X�T?�)=si�<"m�>�r�Aa'��S�v�6���>3�	?��=�u:>��ƾ�q	�6w�C���o�=?���><�u�}�q?`=�a?ha(?�E�>�p?�u�>
׏��7�<��	?�ec?��U?G[%?�I�>(�m�j����:X�����l�U>�:'>�0<_�=���*
��z2�EG=7\�=$v�dk��>�<�h���諽Dn��>	mۿ�$K���پ�����Z>
��ވ��S��L���������Jڙ���w��.�1�%��U�Kc�����#�l��e�?�!�?�>��S��\�������e���hA�>�pq��t}�v���n��g��t�ྒྷ����v!�5�O��h���e�QD'?u���ȼǿ������ܾ��?`�?�y?u:�N�"�/�8�� >�\�<躣�!�뾷���$�ο������^?���>c}�S⤽���>A�>�QX>��p>vЇ�y.�����<4�?=-?a��>�r�#�ɿ����$��<ȼ�?V�@�B?st(�$��R=#��>��
?R�>>SO(�E�	t�����>U=�?2��?s�^=�W�ZN�R<c?K�<�;D��p:��F�=J�=�V=_���H> ��>w��4�=�nڽp4>���>������^�#�<C�^>��཰����Մ?�y\��f��/��T��T>`�T?�(�>�N�=A�,?F3H�yϿ׫\�,a?�/�?���?`�(?�ؿ�	Ϛ>��ܾ��M?�B6?!��>Wb&�L�t�yi�=�Ἁm����G"V�n��=���>t>d~,����O�=\�����=4� �����hR-�z�����=qؼG"��ԝ�I6}�Ru�^K��c�Q���{���>�>�P>o3O>/+8>;{>tA? �^?�J�>��>
�۽�Y��9Eоt�ӽJ&��Ma��/.z���o�6����׾����$���w��q
�����==�j��=g*R�ɓ��~ ���b�V�E���.?TT#>#j˾�}M���9<0�ɾXb��G���Zh��~H̾�0�8 n����?�A?����@�V����x��_1��YeW?ΰ �&!�f
���C�=���}�=lR�>f]�=?�$ 3��US��6?@�?����땾`Y(>T��\7=�?�,?�꽋��>r�!?���φ��+��=�>S>�>�>_P>ͫľ����
c(?�A[?�����ǾJ�u>Ƌ۾�4���@>J�=z|d�5�Ƚ�(�=j�ﺙ���R>��]�W���7?l�.<��4�`�+��T>�-�=�`*>��[?��>(�>�V?�$H?�g^>�m�h�Z���V8ϽǙc?��j?��v>�ֽ��������`?Xa�?:٩<'$1��Ծ�	P�"��\F?2N?p6?��(�5s�ҽt��>"�.G?o�c?w�]�Kӑ�u� �A�r�=��>�)�>���>z��뫏>��Q?��ȽAח�����Sn�]֜?�2@�n�??�;{�����<�?}��>�]������HM�����|�M=7h�>����B^��8-�w�3��Z
?6�v?P �>�?���7�]��=v�߽�̰?�@�?��V�R<t���a���0��� >�a���3�F*w�Z徖��.�O����k�޾�U+�~�>�4@����>�*>- 5��˿��ȿ��o�YW`��K��B�?���>���= O�3'��P���JY���Y�{N4�2l�>�.&=�2>'o\�k3���H� V��j�>Ȗ=#��>Q�=Ȉᾑ+r��g���_>���>&q>��B<�����?�'�m�ſT啿��6Z?!�?WcX?'�G?�ɔ�T����!'>�J�>��r?.�-?��'?E0����f�>B�R?�%��[f�x`A�>M�4��>��?�k�>�;��{-=��>�9�>�TY>t�3�1��^d��"p���ܙ?/�?�0�D��>��?��.?ב���)߂�Y������@?��>�e��"��E��ތ�م�>L� ?8�+��	A�k�_?5�a���p�@�-�jǽ�ݡ>0���[�@�����V1e��⛿��x�A�?J�?��?y���"��
%?'	�>����'Ǿ@'�<���>G�>��O>(\b���u>��r;��i	>��?�{�?zQ?�q������^�>��}?�k�>㐃?�;:>���>^I>񃠾��p��=�_'>tRս��?"4I?� �>��=��N�`���F��Z�����V\=��:~>tf?U�H?��;>�7���ǽ����j���2�9��=�����Ŋq��W,>$$>K�.>�����PC>\�����ؿ�������zW?�2���0 ?hR&��#���ߜ>6-D?DN>gFN�����P̒�L�+>	��?�$�?��?9x���K<�6��@��>���>�\�$�W�����?�=��J?7\�=�nj��=�kρ>�4�?5�?76�?XJ�G�?��Ծ�%l��GF���׾}Y9�f��=a�?�K����>��>�ܝ;!�}��5��F
C�#��>a��?�v�?[#�>��m?Ģ��)���y�i�>�I?���>-Z�= �ھ�h(>��	?��������+�
q?�[@(<@,w�?sf��u�ſ�↿آ��j�����=5x�=oSC>Дw�_��=`�<�+��Z�5����=��>U*�>��O>��#>�p�=��>�E��C��[���H���k�t����!�<}1�����"�!��J��򠩾+�i�h��"=��)���W�� ih=U+��E?F6g?(��?�s?���=bt>��
��g ��Ŀ��%9��h�>
a;?maT?3&�>k`m�c�d�܈� ^���W����#>AB�=#_^>:o�>��}>���ݤ>j�>*ʫ>�f�<�P�=��&>峋>\�F>,��>���>�PH>�C<>��>Eϴ��1��e�h��
w�I̽0�?z���Q�J��1���9��˦��	i�=Jb.?|>���?пc����2H?!���x)��+���>x�0?�cW?�>��=�T�+:>;����j�5`>�+ �{l���)��%Q>vl? Sf=Y�z>��F�1�6�=&����ǎ>��<?����Mj[��M~��9���
��>��>!��=���趇�f�f��������=9�5?2�?	hZ��־Z�Ӿd�׾Vj>�¹>�bT<뗀=��>u���q7^��r����V�k�=��>k�:?ب�=�*>���>X��4�R7>���>e�=�)r?�d?}x���D>�T���!�>Ӽ2>��2?���<s4�<]J���'>�n�>ZQ�=�+s<���bh��\�}�-��>^���m'潃r�3�u��Z4�A��=(ٓ=o�r��Fe�/"=��~?�{���ሿ`��a���qD?=&?8D�=ݴC<qy"���0+����?��@he�?r�	�y�V���?5@�?�杽 _�=��>ϫ>Z'ξ��L�x�?Gƽٷ����	��#��J�?��?�/0��Ƌ�"l�%J>.M%?��Ӿ�F>㕙��H���`�H���<_���>0�w?Nt*�}=�A<��y�>w�	?����$��'Wſ�x�$�0?y�?�>�?w>��84���$?8��?>M?�(b>,���cg�n�>Ff?�3r?@?`6ھ�j�7�?�u�?v(�?�sc>�
�?��?:ʹ>�t���%��P���{��>��>�FN>�o�>ѯ�=����l8��C��?�K�u3S��xV��7>Cߣ=#��>5�w��C-��/��c�i���Qn>ܾ�>�j�>��>�|�>$�?���>�U�> =&<T��%�=��LK?�F�?2w���g���<��=)�3��x?s4?T�üm�Ǿ�+�>�fX?q8�?�5\?�А>,���ܙ�����	��T��</ O>Ŗ�>N�>N���";>3�޾;�5�IT�>[Џ>�54�=�ھ���=��ɢ�>�V$?`m�>���=�$?�?�y>h�>2�5�����>�[!�>���>9+�>lvz?�_?��� �,�jy��񱗿�TZ�|�V>�bt?C�$?8�>��������|�0��G<>^�1}?Hq?�1�.W?��?[�E?��I?M�><V����cW����>U�-?Ě<"t-����U>�!.?�O?=�>�ع=�ev�u�<�P��o㚾m�)?�h?5?����][�w����>�q�>Y#޽�E���	����=EU>���ge�=���=��=�/��J��=�$�=$�B>g��<	s/��^�!�4?5�&;����;�>]T��3d��>�1�?��6�`?��%�5t�=Aٿ����������?���?�=�?�躾p�y��@?��k?��+?&D�>1�I�xr쾡��!엾L�ѽ5$B�3k���>��=�'��G���>���[e���i+�� r�6�$??�� ?��$?�>�G�>-?w��G8���)���:� oZ�x����� &���;���I%����<��о�/Q�ʁ> C	�u�N>��.?po�>��>���>�	�n8>��^�n|v>�_�>̠�>�Q�>�a�=\��=�=�pH"?}���"�9����<�M�Q?�cN?�)?卾�y���!���p?�ޚ?[<�?=xm=�e�N�3�3%?�?�E��KD�>��)=��<:��\�{̾;Ů=�[f=���>i>N#U=!`�"���7�ؙ	?�s?��>Z{��謾��׾Ao>�c�?�_#?/�(��wt��<���^���9��
�=�i� �|���+��e���i���l�ԃ�\�L�GCK��%J?��?	�ɾ��>߾��r���5��a�>�7�>.�>a��>��J>D�)��wY�b���5��ɜ�Y:?�d?�H�>�'F?��;?VJW?�VI?���>�V�>z�¾�8�>Q�E=uU�>���>�#?��&?*�7?�"?bS/?�0F>��"�����%�ҾD(?`K?��?���>M�>����ě�;<	����j��d~�8�= ��<�S޽1��(6�<�S>,�?o���?{B��:�|R�>��`?J��>ȋ�>\�����۾�+��S�Y?�D?�V?
�f*q��$��U�>���?rr�<�5�=��q>��=������`��<�6�;Kl�=���O�'��$�=?�/>�_��.�<�g�=�Z8=A�>�~�=nb�>��?��>�M�>��I� �����ϯ=��X>?S>�r>_|پ�~�� '����g���y>ce�?�m�?��c=n��=��=㔠�s�����콾�2�<:�?�L#?�T?��?��=?��#?��>��A��JP����j�?W�+?��>��Oʾ𴨿c<3�e�?��?�f`������(�؈���BԽ-�>��.�y�}�2���5�C�9*b���������^�?Sҝ?�@���6��?龫혿���`�C?\�>2��>���>�)��#h�;C���=>�$�>q�Q?�5�>6�b?j�{?jy??�/0>,�&�a���қ�4-1>�<�>��N?�Zj?Uy?�'h?�4�>+�F>��i��I�� gϾXӃ���;��p���/i=�>jQ�>a&�>N��>G�=� A�Y�e�5^�~��=�> �>�Y�>��>��>��=��J?���>|����8��"���υ��c/�yn?%��?�Z-?.\N=Hl�Q�I����:��>�v�?'�?�h/?D�^�т�=��[�З��r�F��>T�>�z�>�W�=�i=g�>���>���>A�?��{�f�1�1���q2?�}C?�#�=
�ο�|���ľ���˪�>�V�����Q󑾀���DK~�f�޾6��}c�`�=A����C��u��`���͵���&�>���=�Ē>'�=l������<$�=�����;�����j��_w��d�㻔H�<,��������Л=Z��=	�̾��|?� J?C�,?�wC?�v>u�>��K����>��v���?}K>^�r�&ͺ���3�|������۾^Wھ�b�󖟾�>�fW�!g>nv1>��=BGz<�&�=���=�j�=D�ʻ�=��=n��=AY�=���=\t>��>�6w?��������3Q��Y�ŵ:?9�>
y�=�ƾW@?[�>>t2������b�.?���?FU�?�?vi��c�>J��	Ꮍjq�=ܽ��;2>Y��=��2����>��J>͂��J������%4�?G�@v�??�ዿ��Ͽ�^/>S�3>�0�=Q�R���2�(�_���W�#�Z���!?�*;���̾+��>0�=^ݾh3ȾD�=Z�2>͸=����Y�P0�=I�o�j:=���=���>�$B>'��=�ΰ�P�=�E=I$�='`L>2�����/�ˡ6���;=gȽ=��^>�F%>��>�s??�&?��f? _�>��u��¾ot۾��>�*>t��>�R=o�>�Z�>�1?U�??�Q?�g�>F�=���>�w>e(��$d�ײ���j��dq�B�?��~?��>O+=�9e�M�"���T��h���,?��E? &?�#y>�#���ӿx�+� X,��^(����ㄹ<I����@�@Ŧ�6�2�c襽��>��>�7�>-M�>%�V>5l5>\�e>��>>]�=�^=��=��,=�a��.��T �GZ�<F�(��� V���9��.�?E���X5�7�|�>=s;c�>�U�>M�> ��>H���d>>���\!U�goϼ�Y���\D�f�R�NZt�P4�����i]>=�>%̌�rD��>mG?���>�Q
?$��?�`?0��>>��&F	�"���&��|��B3�;�X`>��U���֦F�}�=�������>
�=�}z>��P=��
�2�P�CT�<W���B�R&w>O�=������ս?Z��#֨�������8��2I=�?z)���Lx>�+�?u�~?�n�?3��=ֲ>�.���(�Y���P�Q�<���������j?E�>�W�>@�վi�p�i�����U�7I�>
i��<G��o��T�����q�����>4�7�7��¤)��㋿�F��GJ*�S5��ޭ?�2?A��?�z|�(�b��l\�0@�-���@��>0Lr?pG?UC6?�?|}�=i؏�z���f>(N?G��?au�?n{�>��=�Y�����>�?�ٕ?+��?�On?�wU��n�>�):�b>S]ݽĹ�=Np>M��=ʂ>�-?�?�n�>�㡽py	����)�PP�C�<v�k=~�>_6�>�w>Xb>�o�=�<�=#�h>�>9s�>�o^>��>N�>�}��wi��(?��>/�>�*1?Ņ>7=9"��y��<빊���U�\� ����TH���R*=���<º�<�Hd����>+�ſ%�?�CJ>�D���?��LD����g>zW>��ҽ��>YxE>��>뵳>�t�>ذ
>"��>(�>e)���>_���X�	�5[{�<�n��{����>f4ʾ���X�&�)Mi���P�m��q�<X��Ŋ�t.�r
�=�0v?���k2������E���^�>ׁ]>��?#/�JB-���U�y��>�Z�>B�j5��������_�?�+�?�d>bԟ>7TW?X?�!0�Í3���Y�v���?��tc���_�Ϫ��ˤ��jc
�{ ����_?�y?�A?S��<�m|>�?�w$�񹏾?}�>K�.��C;���?=��>�\��Fi^�w<Ծ�tľΐ���F>-�p?�d�?s�?��X��k�=̩G>�?�w&?�fD?�t*?E]?�t��%?K�=~�>C7�>R61?��8?4�?@�,>*a<]��fs�<nD��?�,��A)��ֽ��
<#U=�qk=��F=2��;��޼��1=[K`��Չ�FB\=�<�;=�<Y��<a��=��>�oH?{?7?�k4?���˷�j�� 0?�Us>�� �¾D��\aƾv�>W�?JW�?��?��*�YA��M%����>y�W>6�3>~�@>�w�> l�ǋ��H�=�O>�>��>�>=������,��KMݽ>�*>ڲ�>w�>@�u��>Z>����_"l�[�>x{��쑾4�-��5>��/&�^Ã��[�>�^M?u�?���=����q����X�*�'?�q>?�tR?�Ss?��6=�]�F���5����8�>7�T�
��Z�����\9�"w1=j3Z>����
�   �   ���>0�ؾ=W)� �Ⱦ6X��ֽ�=޽?j���>�ܜ<������?
��[�̾��;>��>"̩>��B>2X>�¥>I���-�>��=}��X�[�[�^>=t=�
=V�=�R=Z�]��/����6�>[�=���>s)�>q[���|=?N�4?���>͐&>���DI�_�xK>֓�����;O
�*��=@ڞ��-޾	��}�t��lҼͼ<�u[���l>k?>�����Jн@SD��Ű��}�=�9F=��b�	贽7'�>��=n.�>Zz�=u+^��V���MC�k��G孿�������kZX=�n�=Č=�5;��%=�ǉü1�<q�,�P��a-�>��>{1O>�� ��ײ1��7�=����v��.Ψ�9��R_���)�=�\�=��X�����i��;Q��T溾=��O1m�����4�����(�)}�;o(�>���>� 	>��>�*?hE?ݗ�>E�)=���>v$�P°>qK�>��	?p�>Ń6?��>I�E>�>��B��z۽Nۦ�7�=SqN>"3�>�>J�>��H�M,���
�?y^=�6�=�� >�ɂ>��J= f��<*��?7<�^>��>O��u61���.3A�1���΂k=�?yL����%>�r���g0����p�Ǿ1u��GX�>�-�>Hg�>���=�~{>��v>���Yb�O��>�8�=��&���<��ý8�$>R�<��ռo�x;�dO��G�U��<'sd=�Ob>@��k�P>�1?,�*?�W=?���=@��p` ���"���۽�z���P�Y��>�X��	���&꾵�	��ξ�K��=R��&�&�ؕ�>�]>��H����%M�<xk(�n�"<��B��=wb��Bʸ=ϭ=V��=���=/%伮�O��̅���Έ먿�D徦�Ӿ'��L��=��9>,�Ƚ�A�F��H�o��ȡ�Z����m�>o�:>a�=լ����/��m#������t�H ��^��&�������h���tj<�UN������/�n��=?��� J �����d�4���ں2��f>�J�>��><�>�>�,?h�?�ߏ>��8<��>{��=&<�>�P�=p�?���>�Q�>�	��;5ٽ�����+�%�|d�2�	��م=�`�<�9>��z>	G���L3>.��=}O>)&<��}=�!T>�=Q���ޤ==7�;�$>'ȍ=�������
��x,�[V��8>�8�>�-�U"�>��T����<l�~�c�B�����߇>�T?�j>��>�p�>��¾���>�s�I�7�`��>�Y>�v��q�=N��$'���=���@��Q�D=u_�v!>�5%=@>��?h�?��>��>�Ⱦ�oA���g�>%a��꒾���>bT>��c����V��D�;
�G�>��2��򽽛!�>�*�>pOT�t>�="�>4w��N�#�:�R>G�=�k=F4>&V>�B�>e����A>�;��XG��ÿ1r���t$��񠾜m>���=���=Q�6����=���C���<I��U��D=T;�=�O�=�3ܽ�#_���߻t`�����,���?��&��"��j����:�4AĽ��վ��>4����˽��	����Պ�Q���$L�=�?��?�}>nA�>���>�p?'ؑ>�0f�74�>�_��F��>WU�=977?�>�"#?���>5��<�a"��V����a�
�[�G>��g>�=er�=�4b>%Y�󟙽w�F=���=�	����=��%>o3�=_Y=!��=e�X=!K���NP>.	G���U��{A�o�|�F�¾�����96?/��ņ��;%�A9�0J���  ���r���=U�>r�>���>߽�>#������m>��ȼW	��,>f�B�QS�^��UJ�=�5��y��B��U�=���=�Zu>40�=��V>�5?�?	?9�d>t�ξWh*�*A��N��:� �r&���\=���'T���:��E�¾��2�ؾ_
=ᅡ�B�=�>�e>����rv�Bc������H=Un<|�>�.;��Z>H�>',�>:�|=$�,�U6�����῅�ÿ�<���d���@��@;�=
��=�(��N�ω8>�R)��B��=��>=�u>��>nlT==����������}\���&�T¾��5Ͼ��m�Un�~w,��%ƾ�d
;��J�3�xݾ8����r�� x��d���Ƅ�9��=1��>C��>�Ѩ>!ѿ>ҥ?_�	?�>���H�>�>i%�>��>��?���>J)?�q�>��>�>�d��a��R���=����mP<Æ>��=��`�>G��=Z��<,��=�W�=�6>e�\;�~=\��=�U=�=���>0�ؾ=W)� �Ⱦ6X��ֽ�=޽?j���>�ܜ<������?
��[�̾��;>��>"̩>��B>2X>�¥>I���-�>��=}��X�[�[�^>=t=�
=V�=�R=Z�]��/����6�>[�=���>s)�>q[���|=?N�4?���>͐&>���DI�_�xK>֓�����;O
�*��=@ڞ��-޾	��}�t��lҼͼ<�u[���l>k?>�����Jн@SD��Ű��}�=�9F=��b�	贽7'�>��=n.�>Zz�=u+^��V���MC�k��G孿�������kZX=�n�=Č=�5;��%=�ǉü1�<q�,�P��a-�>��>{1O>�� ��ײ1��7�=����v��.Ψ�9��R_���)�=�\�=��X�����i��;Q��T溾=��O1m�����4�����(�)}�;o(�>���>� 	>��>�*?hE?ݗ�>E�)=���>v$�P°>qK�>��	?p�>Ń6?��>I�E>�>��B��z۽Nۦ�7�=SqN>"3�>�>J�>��H�M,���
�?y^=�6�=�� >�ɂ>��J= f��<*��?7<�^>.?fI�������H���b:>���>T.f>0� >��>�e���� >�,þ,P�=j�r�]輦�=:+>ߤ�>�S�>rL+>!�]�l\R�;�W>D�>���	X)>*iO�y7�H�����/F��'�;w��=�C�=� >�=$��;��U>|�T?X�?Ha?j��>m��S������m��9����>�Z���=���r۾����ržٱؾ�����;\r=����Y>Ȭ���0��Wn=��V=$�==Q?<�	�>���=-��>b��<��=P�)�g$c��`�vI�=�ѿf���oB��Z�辻t�_2�����/㓾�G�:D�=RԽ�LD<#�">r�>n�>g�> $=��U�F�=X����"2�؄p�ýq0ž�=T�I��	���
Q<���@B��~�=`:��Ǵ����JL��D��s���^塽�=�>�R�>K��>〼��?���>k�{��>�X�1��e�=�[S<��u>Qr�=�K�>"�o>v>��V>!o��,t
�޽�ܯ>�{>���=���=��=F���!�7>r�>>P(轔Ė=hA�=�����^O�v�=�=�y=V��.p�>��=I�.�C،���!��C1���?�Tw>B�y=�<�>͖��+x>�U�<73�u�%/���½�R�<���=���>b�`=s���C�<�b>���=⏏��B��/�z�ܘ�;�̇����=�|�<C�/9��_=c��<ah=��%>�͓>JN/?�s@?�R?utQ>��ᾤ¾!���y�����>_%l>��.�:��=����9��Ӿ�>��������i�<�L*>��=���[=Rw����I���>�x8>�Ž�0i>y�T>;�u>��;>���=�#D�� &��D���{���Ϳ�?��L�վ�׾�cP=�l0<xҖ����P=6����Bs��M^���Ҽ�{=��> :�=΂M>�y�A��=��L���Wֆ��Vͽ�h����L���D���<H�=n�;;�E������J��[��o�ʼ����'d��1)��K���}�>��>t�?�嚽)��>���>̼Խ��
>}=cӾ�7.�-"�=E��=[E�>Y��>���>��>,B>��;�pt����0��Ԉ>�B>�물&�3=5�r=}r����=h��=Ǖ�~�Q�-�
������}��)e=��>�Ƽ�d�.?fI�������H���b:>���>T.f>0� >��>�e���� >�,þ,P�=j�r�]輦�=:+>ߤ�>�S�>rL+>!�]�l\R�;�W>D�>���	X)>*iO�y7�H�����/F��'�;w��=�C�=� >�=$��;��U>|�T?X�?Ha?j��>m��S������m��9����>�Z���=���r۾����ržٱؾ�����;\r=����Y>Ȭ���0��Wn=��V=$�==Q?<�	�>���=-��>b��<��=P�)�g$c��`�vI�=�ѿf���oB��Z�辻t�_2�����/㓾�G�:D�=RԽ�LD<#�">r�>n�>g�> $=��U�F�=X����"2�؄p�ýq0ž�=T�I��	���
Q<���@B��~�=`:��Ǵ����JL��D��s���^塽�=�>�R�>K��>〼��?���>k�{��>�X�1��e�=�[S<��u>Qr�=�K�>"�o>v>��V>!o��,t
�޽�ܯ>�{>���=���=��=F���!�7>r�>>P(轔Ė=hA�=�����^O�v�=�=�y=V���?��齐���᜾z�����>�݁>��>�����*��?��==Z��=����=�3?>��/>���>�Ԇ>��C>VG"�OZнJ��=��8���6���9>�aȽ�F��Ċ=H�Ҽ�YG>��=d.>��J=YÑ��+>�?>0�>��B?��O?�@Q?0'�=W�
�����E_���������7>
��<���<�l�wl��z6����~�%�r����$�h=��o>���>�Y	��%�Ε�=��}�"W�=4D>��X>�H=��>�b"=���<��ǽ��4>S���3��ſe��a���L�?=m��b����@���Ž5�>�{���j��ɻ�ǁ=��u�@�">�[�=��=s;T��y��B�B�F�۽*y0��?z��� �D����½.n�<G<y���1��L悾���!���ED��<��c�X����0׉>c�?�X�>��
>_�8??Z>h�=�W�=j{�=ю�'S:>���=�M�>|�Y>���>��>Q;=ֿd>u�h�U=����N��=��ǻ�4>��E>�;=���=��<�^<�����:��c���'�#�=(ӻ�����H�%�
?�6پ8������BϨ=vp�>Uh?�l@>&�%>�?�<p�֞-�6�5��}_�]�[=QGS>���=T\>>��>&-�@�c�0Eľ�>�2>��/���<�+��\a��
��=l4,>T�=��/<��,�o�Ž2ZF��D�>/y�=�w>��?�a?^#?F=����(ͽ��y��1���(�b(�=�hZ>>��=��<&k���
�.Q��D~��y�bz>�=��?=�L���=�u���%>�]�=C1�#)���=@`m<�e>��=�C�=W�����⽟���������ݪ"������rM=�I(=�D��Uת��"弸���۵k���E��y*>��>�h\>2�׼,�:���= �+>ǰB>��=��7�����2��~Ƚ��=i�꽞%������֩��{����O睽CE�y�e�Ww�s���Y&��(?���>z(�>_�<?6|�>CPm=K��<���>�m����>R����R>�X&��|�=��7>@�>�j>�H	��T���^�0�>	�=_�G��Ǫ=�$>��5�֦�;�_)��r_=�P����`�Ũ^=�O+=W	d=�@�=�Y,�	(x>���LՐ��/�|$��c�a�Y���w�>���>CJm��pѽy?�����6�&T��7)>����8��˻�*N��-�� �B>p���P����=��a���U�פ>Ac)�\����Ő��0f�z�������b1�l�����d���o�q5+>n�m=u�$?`.?���>�Ɔ>��վCN��.)�1x��JW���i=��R�o��ҾdM;��Y*��Z���wI��L�<v�3>�͑<`+�;�rA>�L�=��Q<��:>���=���;��=5Y%����>�W�>}:>U��>�QR>��ǽhۻ�����;��1���\��ۡw��lu>����:����>҈�=�5J�[�=ׅ�=�A�=1#�>�¿=���=��#>\F�>���Ͱ��tx�!�����ϾL����0���򧽽鐼~��:R>>/���ž�ݠ<Sۻ�*u��&N�����J�)?��>�F9��5�>"�?TD&?��?Gu>ᦶ>azt==�?}��>�L�>�X3?��>�� ?�+.?� ?��>BNh=^S�����<�Q=3��8��=N�g>�9��
�=���=8Q>��Y>��8<�D�J�;��>z�>��>�,X>&�=�`>?-ž�?Z�$2}�b��J%�=�i*?nk¾�쾸4.��e�&�@�˼M�{��"��m5&��F�����>[%�>�s�=�>�>�ғ;M�d�%��?��m��)1�=+K=��<j���T8���_���w���QEQ>k�>�v>8�;?��s?�&?8sf>9�F�̕T��P������8b>�K=߻Y>���;��o�Ҿ4� �tG��|7��
ƾjE�c�r>������ʨ�=�S�<�K�J �;bΦ>Cs&�e��>]'e>�v>��?஗>֋�>�߄>�������,߿�ش����ʪ���U�<�y�<P��>�2n�g�1����5Z齿�ὡ;��� �=�u>��^>~�=�١=�5�=���:��w;$9
�S�S�1����@=��(���=�c��ͥ��'�ƾF�o�3�&�)V��^����ݽ����rµ�l�Y�7�?���P������>?�8?�1�>V�=�� ?��>>��?g��>��(>%'?*?��#?I�"?8@?�jɽئ?�6���"���*���e�c=�@+>`i>K��<$�|�Qy|=;9��ɂ�]�F��$EE=)��=d�ػn��<��T>�S���<�AJ��D�s�t���ϱ�>�׮>�:�����/�z�������y=�S����ݨ6���
�A��>��>�0>If
>c�Y>?ٮ��P��#�=� �n�M�iY�=�3)�l�]�fg�<����x5���E�pż��\�<z��=��[>��C?�UZ?�-�>���M1��ym�O�-��J���>wa}��H^�*ý�n��v���iH�s^���~��� 㾹x�ZT�>���sz��W>�I<1���{�<�?<�ù��=c5�>�">g��>�*m>X��>��=>��<G�U��0ӿ���f�}�IF�s�F����<`��=��>	����p+=�%2��)n�Y[��:.��>ʯ>�O>y�">)z=f���H���ܒE<j,�i����v��n����#���辕�A��{��J�S�-�9��z�<OK�4!�����º�^�?7��<�+(>���>�\?XK?V$u>�b���2?$�r>1m)?�,?NQ�>��D?S�>'�?��0?��?O)U=�吽шE������s=��/=��>>�v>��>��2����<w�>L$��{���kU�=�	ݼ?v���*�=m��=5 �=YT��L��6L��;�O�a�����l�>��?����*
۾�� �:<��.u˽Ҡ�����­��[����������>$,=v����W��н̖��g����쬾	xȽz�>=�Ҽ�c��TG��꾇ؾ�}�e8n���>G>��?��;?h��>���=�-ؾ��e�;�5��������=:�>3ɤ��h��"V��z�� ��\ɾ$&;��h�=�S�=r��>�+�0Ț=\�A=Gc��)�M��=C��>{�=<2�T�>kԙ>�x�>�)�>b�>���=�6�E������������ؾ
]�2L�<����n�\>U�
>G��i��=K����.�<��>b�>?0�=S��=7D,>q�t=G�+>��ʾ�LI��(�=�
�9�位n��Q8���h��0��&ܼ1E���E��},=j��*9<q9�<�\�?
���$�;��>//}>���>���>�?�{-?��>_���<�>��B>���>a�>Ta�>S)?��?��?� ?q��>VB轀8���,�{j=W���*|�=���>���>���=>��Q=�08>	þ����E����Ӵ=#�,=,>5	[>M�h>���=FH���=�g9O���B��)�e(>YfN?u���f9־�1B������f�Ѿ閽_��"H�F����-=�&�>�{O>��>9��=��>��=�v�>��a�l�ݾ_K�<6p>�:�=Z��!���$��h'��V�V���1>��>���>atB?6�C?�e)?���=n�1��E���/����a>B�B>�u�����k�����lZѾ����!����<�G>w�<i߈=&g)>W��<R۔��" �jT>do?=�w>��>��\>�a�>�&�>>R~>ۃ{>Kё<*���{��7;��]�����о��o�G��=��<l�B�~�����`>���;�<w�wE�>��<���<��m>��b>=�<�Ҿc�Y�&f��$��� ���e�9� �H=�>"�U��ؽ�^�=T��"�J�jľq�ս&����E��RTӾ]bi��v�>d�=�^>�4�>ӅI?o�?�u?i轗:�>xKK=�?���>�Ȁ>ȸ"?�4?��?�?2?�n?�0n=}����k�n��;v��]YI=yA�>�q�>&�=�e>{��tǹX���;<���>>�Y1=��=q4>ޙ�=	��=�?���<椾v%�� V��c>�`�>d�=߶�>�x>��4�R>b�>�><>�Py>G�|>��:;I>>�i.>��>����������=�X�=޽�M=�>I=*����= ��=N���L@=��=
Z=��$��r<vx�={��=Ǽ�=��?4#,?�c^?�B>�z��YR���:���'G��F�����������~�ľ����ؾtE���t�2Ek����SqW>g^�>r>�U:>���1l��=�)�R�ʽ���9�%��i>=�=�a�=��6==�=/������8m�7�������C���U0����>���=1�!�كn�jvɽY3��X>�si�<����6&���/=v�=/?N��`�;�{-�P�=�;����q���@�V�}`9���=���;n�m��fɾ"�½�������vC�ԓ��W���ɖ�����6�Ǽ���>.���Yx>n�"?�8��do>c��>�#=��=��>�\�=P>Ի�=I�>0�;��%�r.ѽ�Y&�v������=��������=>�� =	�>H�<4��=P,�=H�=R#��fϼ9�����=�o-=g��=s�?=+TK?�NV�މ��f��!�`�RI�>8g�=�v6>��3>[�>��7�	's�*�7���p啼�>^Q�>�#>��<y�I>v=B=�c���N�=�=������h\=���=~���o>͓�<���입<� =�NP�ܓ}�GJ��RMc�<N=Ct=h�:?� -?�F?��=������ھ�:����(y��߅��f�f�����=���1j�9��X���5�<��=�-�3>+{4>N�o>�n>�ڮ=�:�;7�����)������V�/K��ZJ��ݼ�y�=U��=�a�=���'���ɿ�D��VG���v� Խ|�<�4�T��Ӓ=�q��[Ծ�$��I�;6��>���>6B�>D�w>{��2�>����=�<j>�S���a�qw���%�|��K枾�(��������p��u�={;�b�*���]���ټ���s��[�d���*�?��+> "�>��A?u$=ns�>�_�>��>�$�>��>�͵>��>��x>�o#>�/��G\>�v�>����ME����8�==������E�n��=Ɠ�=��ڻ��='*=��=��=~[�=
�=��c=#�{�V�&�s=	!�=�?���<椾v%�� V��c>�`�>d�=߶�>�x>��4�R>b�>�><>�Py>G�|>��:;I>>�i.>��>����������=�X�=޽�M=�>I=*����= ��=N���L@=��=
Z=��$��r<vx�={��=Ǽ�=��?4#,?�c^?�B>�z��YR���:���'G��F�����������~�ľ����ؾtE���t�2Ek����SqW>g^�>r>�U:>���1l��=�)�R�ʽ���9�%��i>=�=�a�=��6==�=/������8m�7�������C���U0����>���=1�!�كn�jvɽY3��X>�si�<����6&���/=v�=/?N��`�;�{-�P�=�;����q���@�V�}`9���=���;n�m��fɾ"�½�������vC�ԓ��W���ɖ�����6�Ǽ���>.���Yx>n�"?�8��do>c��>�#=��=��>�\�=P>Ի�=I�>0�;��%�r.ѽ�Y&�v������=��������=>�� =	�>H�<4��=P,�=H�=R#��fϼ9�����=�o-=g��=s�?=��0?���o�\���$�G�G�؂�>��>��=j�X=Y��:@&����,=n"�=O�>#x�>#}�>Q�>=��<%=B>���>�Y{<�8M<NZ�AH=�
X<Db?=<���g��=�Ɯ=�.��î��++=�q�R6ɽ�E�<t;���=���=kIv>��&?�:?��?�W�>�����]�:�ڥ�������a��N�߾�S��$����'��Z(��:q�����;��6�=O��=��>2��=��=>��q{�=�a�h�7�N����=r��<��=�qu>F��=���=�R��������� ����X�������'��s��ӂ���9�
z%=�w�>��>|��>�F�>��>{�b�E�����A>->�J*��D��X'�<W�|�<1��]����@���g �=�fN������>���Ѽ-H�������c�]�N��7U�����=�-?M�g>�
�>�F?��y�9|�>+��>;zi>ʊT�ro>i�=�(�=�����SG>�#c>�1>�X��5�=��"����=�~��3�<c�S�J=�=�򭽰�=���=�&>5�<��<��=n6h�V�;�U=�>��N<v�4?�=>����p1�O�f�m�=R->�5m>=<�>�ؠ=`]��M����=�>w>Y`�>�+>��>�=>I�>��>#���|���*��������(>�⍼˸<jg��|�꼩��e
�����=��r��v㼹�˼Z1>�F�= >Y?�w3?8�3?n��>ƭ�Ѻ!�а5�� ��ӟ����˽v��F�����.�9�5������/r��e`��TK�=,��>M^i>�>Y
_>���ؚ��^��������^��'�a>c�2><kc=/>�0>Pj�=�׋�����ٿ��k�|1�r�f������>���=�(=�x�=(� ���>=�>i��;�g�<�}m�����w=P�;�y��>�Њ>�Lྱ�E�rMY�2�������"d~>� �m�6�Hy�/%��Ľ�WR�vx �RVG�r􂾬<���ŽAL2��?}�r>�ש>Z�+?�.>SP>�]q>��K>�*>Q<�>�Oh>�Ȩ;�*>�O>ݷ�>(w>:��ɽ�Y�F�$���{=q?��j�c<�(�=-�o=D���u�=�1�=�k1>.m�<�V
�<�J�zHV������wf= >�5�<٪?�-m�U+N��w�O� ����>��>1�>
���>7��'��M���j����W��e>T~E>|X�>$�=^Y�>T��7+�6�署�>��>쮽4O�j
�=W4>���M��'�4��	>�qp>�L>�{f>�M�=ԅ/>�u7?Hi5?�?bA�>��ؾ�U���3��K�xGͽ[�����E���c־�n3�I"S���O��&1�ȋ>\t�< ��>���{=O�s��;B���̽qM >ۼH>�.>=��#��>@��>vjF>}�f>���=�G!�y�����ӿ�a���І�����Y|&�8��ܒ=�k�b���N�׾RR�sㆾ��1>���>�.�>��>wp=���Ε��cT�{�q=�d�	%���ؾ"�����1�=���?xe��pY�����ՠ}���G��;�i�J�1�H�Z%콧=N�i�>�>	��>|$�Ĝg>�`>�Ď>I�><?Ȓ>P�?0�>��>���>��>Y�>�%?\�T>��K�ƣP�e��]/�>�H�>X4>�-�=�/>kX׽R���ϣD��y+>�.�2�<�<�'�='ՠ��.'�}�"���>F��>�v���Rc�"뾁2:��C>b_?%�?O�־��H��jS��dU�2��b��0>�`0>�@>���>��k=`��>mk�=�؂��NO<��>�ف=�CR��9�<R��
�ͼ3�<  �g���H�	��{�^rd;�f�=7�>�P�=?�>tB2?�r+?��	?�-�>�3���C���5��b#��<����ϽX����d� �۔7���D�.�J�.�����E=��%>rMM�R􎽠��<�D�G�n?2=E�>U��=�e�=��p>��>�p�>MI*>�*9>G]=5�#��$!�rR���z���(��X���q����="�<
sǽ`6,������wj�tB�)��;��>U��>V��=�T�=hl�=���=|��Hi���н�l�qzʾ�����i��p&������������V�1Q������ء���+�(�K��~�>0��>��>o�H���>׫�>@�<e�=o�I?�?���>��>s�9?���>�v>԰?�?�>M�ν���QF���Bh>�U�>Ě>w>���>�jw=�'r��Qɽ��=%����#!�������L=ѓ����n=�h>6�@>� �>����k�'HӾ~l��Ӳ=���>�O#?������������õ�y���P�mG��K=;�5=y�>E�>�7�>���>(�#��.�5��=� �u�%���ϼ٥���; ���g���@��{C��5Z��G�z�=�T9=��<��x>ph?v�A?m��>v�;��N�{�V���<��D�.�vz�>��=a�O��Q���5�,�K�(T��������)J>��=L�����ȼ4���缏i�<u�s>K�,>{���q�=ap>� ,>��b>�.>�>���<*��h:ֿ���v9�56̾nY�=͝>��(�F����'��B��"����ҥ�k=˂�>��>c��>���>ʊ[>_�4>�j{�jǋ�(�%=����HTݾ�H��O�q����=���F	���н ���S$���c�q-�b}&�h'���V�4�2�C��>��?=�m�>O�>3�<?#��>W�f>J

=r� ?��>bȉ>J��>`��>�?sL�>� �>	i�>ͱ1>�O�<MH���5d�
S�=a�>��8>=�>�}1>�D�����<�����6�=_��=@λ�C>��>R�$<�}=��-=��->eY ?&�*%'��e����I�{+!>�ǿ<�(�>�쾗��=�I���1��Ϗ@�� ����t����`g�>�f=�K�>P��=�@L=�9l<5�=4o7=�@���@�ܺ,���<v�`���=���=+�)��s���w~׽l�>�b.>>&�>�k?�j,?��>�T�>�L��M����>�<P�KH�>/Pƽ�ۀ�3b��z��{Y��dL�q�,�E�ٽ�����Q�=h>ٽ�g<�j�=W@'��=���i>���>�
�<�>/$N>��`>���>�:�>�ρ>B�>Re�9���t6࿔.��xbž���o=T޻�R賽<"Ⱦ�m��i�P�`:���󾦭q�
��>��>U�>�>�=�>!S��[���s��^�����"!⽇D�� �k=ݙ��������(�3����J�9U��'��S�#���SH򽟁^�r��>��[>���>o�>i�?�u�>��?�#P>��?���=���>�8�>�?Z�!?�7?���>�; ?@J��3���@���k0�o"	>��=��=W��=3[ >��2��'y�[�:J=+{"=k���Vn<#V�=cn<�0���G�<V�$>�T?���G��Œ�K�[� ��=��>N;?���������G������������H�Y>�K>.��>L�=W�V>�@{>m��
��=�=���VW�=�����<���=��½'�	��������K*!�_��=,����>��X>әT?�;O?�?±?'98��M�k*��wͼҦ��ړm>��h3ʽ�fž�O�ēU�Z���M�5U��dȼ�
a>�O�E�����=��?MN�K:=�V�>�z]=X��<��c>�_�>1Ȣ>F�z>r!>��=�Z ��yD��̿�̭�<�����Qڽ��G�,�k��{Q���=�xt�s������>�D�>fM;>0� >��=���=1(��A\���ԽpYI�����s�<2S���#>U<6�lq�����y��Kؽ��F��N�<����S�x��)��r�>'��>-g>��b>qY ?rp+?SK�>�=�4"?"��>X$Q>ZA�>��4?I"?��>�1�>���>��V>>�1��	�\͕��>�0�>���=���=�C>J�Խ�SF�8�����Q>��V=O����;C=���=��ۼ�I�����=��
>hN?����]��G�7pM����f��=O1�>q��'�>$�F�R���΅�-���\�Ռr>�Xi=���>�l>Rs>��x>�D��ӽ4>�Qp>͌������5�R[����<�pI=�tȽ{��זx�X�"�cD���y=}�X>E�>�`=>ht?H$8?;?"� "�Gx����Z�����e�T>lk>�7>�{{���;�?���'��@k���������}r>LE�:�5s<Zc��6��7
�$=*�a>9q���Z�;zɴ�^��>���>�i�>a">t&�=<�:��a�qgڿ��h�޾��੅� ��>rT���a�f�D��Ɛ�����G�h�g�,�<��><�AM>�\�<��c��p~��q>�5��%�=�IȾ_�d�#�ϫ��R��=L��=��Ļ�Ye��>��(�"'0��Vk���<��7���X�:^O��[�>d�&>:��>!P?���>�V'?`?p��>���>Y�m�/�?�T>��>�?q?�$>:8�>�3n>a�?>�@�}�|��8=�y�=��F=�@M>�:H>z�<�r�������=�S1;��ɼ��F�Ǚw�h�&��=I=��>�;�>�����D���K�QMX������l>:zG>_��;+�����ʋ������4�V�����B
�%�>�Te>�'>`7�>��I�$�fy5>8��={�<�Q�{7�<���=A����R���i���S��b���o���Z�=�T�>��0>1<�&_?�BI?��?0Rk�i����
v���=���J�1ȼ�(D>g8�>;�>𖞾W*.�C}�����2��z��e�U;OQ�>:`-�ɪ�<�b�<�����E��#�<��=�>�=.�r>;'�e�|>���>" f>���<K�~<(t8�9V�,Ѻ�����H�����ܽ;ra�.(��c��<c�Y��ؾ���,V���-�nԛ��܂>�>rp�=Q�=���j߽r�X�9C��5~;�M~��վ��!�+?��r��=���6����5�1OZ�i�½{����$�=@὜~��R��J��>
�C>�,�>��?�C�>�6?�|�>���>���>]%�>W�?�k>B�K>@��>o�?;x�>EK�>�=er=�|��\�n+�=Nv:>���=_�S>��x>[X�<�u��-� �xmM<�V�>��>~��<d�A=o��;&����$|��9@>'�����ž�Of��Q�2͠����-W�<��>d�>"/>3���pP���,��?���پJ�x>�%>�[?�N���̈́>YiB>R��<���=��=�[{;��=)�=}�<�7�=�����ɽ)zѽ�ޠ��1n��<=���=�o>�O<y�$�"�?�N.?��>U~�!���#u��[��՜�����a)?-�G>���>{��W)�:�V�d�!��bY���t����	>�נ=�.=�q�<`	޽���3d=�~S>�J�=ў�>���=��>u�>[�?�ˏ>���=/���y�7����c���?h������4Ag�i�=��ýJ$��f�g'���FĽa��� �r=2�.=zOr>�=�i8��w�=�x�<�6�<����$��!�ōK�+y���	>H�����'8˾x5	��O�J�g��?������(ĥ���׾(�Y����>h��>U0�>t7?�ҕ>kn?���>�h>�/G=1P��_u>��=ND�>G�>I�
?>��=cL>U�V��_>�F�(�E�	M>}w
>�">[4�=��=�	�jKн��E�G=T=-_�=�:�q��=Ȕ=��$��&U��ǜ<��>8�>(3[<f~Z��h?����0�ξĶ���#�� ��"�>�1�1jɾ��3�VwB�����M�M�Q�>�V�>J*>k�>�	�=���=j��=̮I=W-1�O�'�_߽���=�y;=�W"����g��Qaž�},�T��=\�>�H>,.>E?��8?OP)?��p�W����w�O�+�=U��blѾ�\>��B>Q�>�н�H�Ѐ:�����E-��y���̿<�4>Sψ=*V=U��e�8���W��>2�>�D��2�->�>���>4�>ʺ�>��>/��=6��t��Rʿ�릿�,��O�v�]]9��v>&Ds>���>`|�=����d�jɼ�[U�C�>/��=��W>
��<�`⽟�Ͻ�/ҽ�O�5Ǐ�j䧾UR�.�_�O��ix.������%���]�:&��6��LQ<4��^)��2+��3|9�I��>�$�>���>���>�n>��?�?|�>3�o>��#=�?,~d>q�>2R?W�?�>?��?*�>v��=�|ڽ}����'�=��>�(�=ā�>9 �>�0�=�y��ǜ=~4�=�ߌ<� �<��1>w��V��.l=t���O�>8�>(3[<f~Z��h?����0�ξĶ���#�� ��"�>�1�1jɾ��3�VwB�����M�M�Q�>�V�>J*>k�>�	�=���=j��=̮I=W-1�O�'�_߽���=�y;=�W"����g��Qaž�},�T��=\�>�H>,.>E?��8?OP)?��p�W����w�O�+�=U��blѾ�\>��B>Q�>�н�H�Ѐ:�����E-��y���̿<�4>Sψ=*V=U��e�8���W��>2�>�D��2�->�>���>4�>ʺ�>��>/��=6��t��Rʿ�릿�,��O�v�]]9��v>&Ds>���>`|�=����d�jɼ�[U�C�>/��=��W>
��<�`⽟�Ͻ�/ҽ�O�5Ǐ�j䧾UR�.�_�O��ix.������%���]�:&��6��LQ<4��^)��2+��3|9�I��>�$�>���>���>�n>��?�?|�>3�o>��#=�?,~d>q�>2R?W�?�>?��?*�>v��=�|ڽ}����'�=��>�(�=ā�>9 �>�0�=�y��ǜ=~4�=�ߌ<� �<��1>w��V��.l=t���O�>e�#?��5=���Oھv׾�ȋ����=�q2?3Z�[��<�_3�q��=3����L��,�? �, 	��3�> ��>+>*�=�f6>��>�<߻�Ԍ=x(�{�	�1LO���=���=��<E�=�v������e��?F�;�J�<߽�=y�>b�>?�r@?q�A?ڪ����/�����VC���ռ�;=9�=���=�� ?M����ݾy��pPG��Mr������~üї�>�a �r�;��a�=1��<�U�uD4=5l�>HD=��<�v���>3�?�4?�1;>��������t��04ѿ�����Ⱦ�r'��*��P�.�#���ӻ3]9=L����5�#Nc�k������=S)t>�ə>N�=��=B�\>�t�E/Y<@����k��Ď�U�}��v�����=(1������K�I=�=T�Α��<��JǽZc&���k��_��@>wh�>^��>���>9�-?m�G?�2?�5��4?<���v�)?�	��܀>DN?+�.?��"?��?��>�j��@ɽ�t��D���>���=ҵ�=�H}>ẙ;,_����o"�=$�=��ڽSO�����;�;y7�=t�L>K�=��?*��`�$��=���Ĕ�N"�>:�?�����c>���4H���#��� �Lh�=^�E>߅�>���>�>��>�����>=�Ҽx(>/4�=� ��,��/��.j�;�~$=ss$��J�1p�W� ��'�<
��=�9�}��=��x=�?.9H?f6a?{������:P��e?�O4��d>s�>��e>3K>)�+�^H��B�!G��4�)}���\<֌l>P�(�PI��⧼�w�ԧ2�l��=��6>�ͯ�`��=/�D>ܥ�>���>S#�>ᮬ=6&��1&�k���vؿ��������-�	�v=���>Ŀ4>'t<��&��u��Ʒ��H��(潙Cd=z*X=�w;=��J=��=�,�=6�����Z������������-���	�T��F C���"<�tf�[y��䳭��-��yOr��.V�m滾sÐ��q��g>��?oT<>6��=�/.?��0?l�I>���=(� ?浖���>�8�>Dz?�0?���>�0�>o�T>�z��F�����=���=w��=�*>}>�ԉ>��C<���:K�z=�|��pfH<�jd��1W�����<%L2>�>�� >�G?GN���oZ�x���:�ۓ���b>��?�料>�6>�:�X�#���΍Ⱦ�[7>��>)�?��>�>�=ջr>�q=���<m��;���=t�ڼ�_�=�c�;�x߼�/��_	�<[C��r׽:��B���_ٽ< ��=쓇= A�=�>�F7?v�J?�@9?��H>�Vj�x�q����c�>�7����>��*^�=�@߾��<`!��*���˾��u>�a�<N�k>�#�}��v=ɜA>SE���4?����=���=�+9:"#-<�D�>*m>�b�=�<�S���܁�� �&�ɿ�ו�`r���d��p �s����D�>��>ӳ�̑�=��ɾWu�>z x��>|I�=��
>R� �<$>c��=!!!���޽c�}�Md[������q"��.m�(�>�XP���'������Q��vQ��*���\��K ���A�K���"�>��?�Õ>�\R�Z8/?�V?gc�>X�����>B�����>v2��^?5�P?B��>�6�=��e>��]�(���P�$�4~o���>L��>��=�S�����>g�����=͵뽶iP>�8�>��A��c=0�����<��>���=x2>9�?���<�Q�e�Ѿ�������iؗ��*�=�m�?��I�ۅɾ��/�0� �������=Ht�>���>X�>��0>��<>��=����'x=�̽�����=*�	��
>G��=%�.��ʼ`(;��.�w���<:.�=l�>���>E'?�?�4�> >�J���R�j��������>{�\����>�/��`��^��@9�V�
��I� �:����;���=�4�=j��=��|��ߒ�s(��@+�需�X��=�M�>x�Q>�w>�'�>�YV>r[�=�9�����տ�һ������8�A<��YOA=�~�=݈h>R?��h��X���T�=����+!=��=\�9>��=��=�)=�P0� ��]�V�sNO�2����"������\=&�I��������2�< 7��A�M����o��!����͇��SJ����>���>�+�>c�?Ј'?�3?��?��d���>�;��?k`�>��>��R?PU8?;�d>��[<�]A��9��(
���׽��M�ܷ�=b��=[�J>�ѕ>��B��P=t},���Q�z�½]���ܽ�|��o[���7�=�*>�>��2?߲~��������+�]�V2νy	&?K����>�X/�������ھm�����1�[>��>#�>�:>�>A،>��<ؖ�=���3�/r=��Ͻ�>S3=�?<˃v�(��UEs�Yb��G0�<yC��Y�S>)��=q�><?��>��?�C�=�x��I�ړ�
v�=U=ߑ�=��Y�*�=!M־�N��!��s�6�þ��Q��"��`�y=ۊ
>jߵ=	��=��L>U+R�������~=���1�=��]>C�?�B�>Pj�>F�"�a�=�3���"���~ҿ�o��u���C�����x���)m��#��|=f�p��:&���X���ý�qS<�G>d1>���<��=,��=��˼d(������U�T�O��=i�m憾��'>��p��������\�r=sIϻ%������'zz��K ��jf�H4��]?i=��?4�&?�{)?��C?\1?�L?�����R�>�C��kxV?�߹>�?�-?�>_=�=L7�>`Њ=��������n��b�=9N���=��>$_>�]�<�"�pbļIK�=~��<�u1�gL���Z���=��>!�$>�|?LR��7����;�y'�j�Ǿξ�>���>����.�ξԽ�⠾y��+���aQ���|�G��࢜<(�Ҿء>���=�t[=�Z�Ϧ���>.֥��s-<@��=ʢȽ#�ͽ��W������A������Q���������ī�ɫ�=@�>>�4?�-?]��ˊ��#��I>����h?%>_ݽ��H>}fu>K[��?�ӽZl��T�����S�<�DI4>+��=��=�h�>\Q��|�����Z>�6=�P�5v>��#> l>L�>�B�=�	��j>%U}=y��΀�U��%�پ�����{��/dt>��ҽu���_,=��'�L1��ﺛ�V>���<��4<�`�=+��=y�=�~����F�����x�=�s��w�[	��>v1��Z^�rJ =2q'�y�(�.��=����2~�"��\|��L��JO��~�=�s�>��>�1S�=�"?���>���u�<���>&B<��V>u�a>��>�>�v�>�2�>,̤>f�l>��>L��c�㽾��<�?��k��<��>��=!����3�=� ��Y�<B��= W��ӽ�=��=�+=���=�z�>1��>��<i��w�H�uB�ʹ��=ȶ��܍>��G8�<5ޥ=������ؾ_+��j=T���(D���O>����\�>�y.>��4�="�j=�r�=E��<���=b-��i�L���ƽL"=)>Nie>��(�|ح�����#�+=�]<=���>Ի�>�l?�Q?�~H�L����6>����}~�����]�=L�>�����>M�������E�� -��;ݾ�z���~>:>�պ�(�k=l��<��� H���5=����>�d>����>	�=�-�>�� ;��6>�^>�ֽ7�h�����h,�ن�<P��=V>���ڣ�췕�tF����<��>~'x=�V�̪��#н��<�;�=P�޾��e��v���
�'�Ǿ�Z��{��!���a��3`=~I=<�y�	�������H��)���u�z�@�u���L�>���>o�>�$1��?j�>�?�>@ф>���>[�<�!����9�>�F�:+�V>ZX�>�p?���>�Q�>;�i��==�	�>��1���=��%>�>f�;F�=��\>p��l�*�)r�=�%R���I�>|=4���>27?q��>[K����~>��%��7�������>�=�w�)>�[���9
:7�־d<�vw���8�=wڄ�;��-'�\�a>[�c>�#>͵��� ���K">;��+<,�n�=chw�j���;̭��M�	���3���>�=�����u�<:��>(�?��Z?��D?n��'����;E��\T�9����P>�ba>�:�>0?M>Lk���_	�'0��K�#���T����)]%��#>�%ԽK����v�>�`�<╾�fG>h�> ʵ�3$�>C�>.<>~M�>���>Ry�=*J`>v<��5ƽ�_��t��Ō�K�B��%	�D>�{�='Y־�ZX����I*�#����i���7>��>g��>8,3=�R��G��>����P��ۣ�s�h������佁�׽yO=6W���:�D�ӽ"$��sP���G����н���=�	p@�+�/���Z>��I>��>'j�<��?��>fr?l!��xP�>����V�='�Q=���>���>I&>��.�ߺ�>|!�>��>C�ɼR��5��tv>���K��DfY>�߽D�½Dz7=R�F<���;��9�8=#Q�<{Kr�r�<$C>���=ْ?�f�>�=���!������+�~�t�[I?���JE	>p��>.W>_c�!���`�|�1�n���0=�>��]�[v�>x�5>�2$���\���w�2>��;��N>[�>�����
�$9>J�=l�{���S��|ѽv�g�8?���.��d��>��>�ku?�r?�뾀��Z�M�����c����Խ��$<�b>>��o���s�x�!�E�}���-��$���:��~)>1|=�L=��>�E��6���HU�2�)>yk�e�n>/t}>J>�rR>�԰>o��>p��=�S�;\�=|ٿ����+���F�=��>�-��о6`P��������B^��0}!�b��I��.8>>�	>��x�.>;E}��?��s-���=��$䂾��씽�m�\��=�}��TD�������̽^d=�o�8�&��Gڽ&[��o��>Ǝ>s7�>|��XU.?�0?< ?�X���>������=/�c=!?�b%?ߡ�>E�J>T?E�h>���>@��0O���/=nA>,K�C2�=@w�>�ν�V��F>:��������̽Bh$>	�ɽ;����=���=�U�<PD?� �>�[��=��lE�c�F��'?"�H>���>�ַ>��o=��!�[�������^\=22 >K�>�_����>�F>�&�D_��:`��s�_.�@��=P^�<ؠ����B�uq�+o<���= �V��v�<�@���ힽ��ȽN�>4�>�D?�;?�� ��嘾�p[���%�u���nh���%����5<赊�HM̾�]��{w�]W�n��L�����E>��u=w�>D����NϽ�'9>\2�=#|��o>��l=�&a=Eg�=8�>5X=��
>@w><NK>���,�����f$����|�=ĊP>By��@����UAH�"�4�˔����ʀ�7G��UB���=�%z>R���	�d��VN�"'���� �M�I м����?q=�+˽�5=��?��0b�Za�<��'��<Q��퇽�RY�q��>��1>�B�>��P>��)?B?���>C�g��$<�8��S}j�e�=�!?�&?f̸>m�>3{�>��h>sf_>�﮽�_����=�B=6�<I�F>y62>�f6��qI�-�+=2�̼,�%�p�i=�r<S��Wa\=³=����B�N=�*X>�q�=����~",�<��*e��8j��Z1?1�?>�(�>N�"����~>��k�F��)���d�>O�?� վ��>��=�t(>��h=Q�p��
�<�6;{�V=r��J�=:�м��=��<;��=�8>s��<��q����=W�C=|�>�R?�=?��7?���D����sѾh�"��6�xb��{�n>�B�>j(��Ee�=�2 >����b��J�о
�g>%���،>J'���H�4:�>	��=��j�Q @��x�>V�A��&�#����1>��:>��/>�r>�`>.?����,>�7��%̿�����4��2�<4�>�E�>
�*���`j&>�<>��������v�v�r>fd�=����O�/L<{SB��u�����=�%�Bn��_��pX���'����8��@���G�� �Y�x��Ó��9������)�R5��A�>���>Gv;>T��>�?���>Ȥ�>l'F���e>H�P���>[�d>XY���q>�^�>��>��=��U�6W>�5��9��� �3��=>@�=Q9�<?,�>֯>�X����h= �]>�m=R�*��b���+4�y�s��AZ>�O"�e޲>*$�=l��=m���)�3`̾1&��Ŭ?�T�>���>o�x�t���ھnǾ⚧��ڼ=`>E�?�"����>�h�����= E>3�S���=-
���=��Y�u���F��֢F>ϻ.�aN��T=���=pq��'��@K=ϋ>+��>u8E?�??3kA�4�M�����!������߽��B>w�6>�&�>/�>�/��#�H��F�b�*��
���ɽ_s�>Ĉ���fM�Z�x>7|%�v$ ���޽�3=�b��>?:���=tg�=ͷ);�U@>V�V>� �.� >��𹿟)8�.Z9�(4�>6��>���>��ϼ��J��B����>z5_����;�;'����нe�7�:�P=��>>����<�����]"c�"X��A�ʾ?���QC�m��=A@�jpa�Ȃ���b׽��(�)AԼ���+�G��}ؽ!��>���>bH><s�>t��>�Sj>���>�w�R����Ќ�G<>�^>EZ�>�M�=us�>7߷=r77>�5Ľ��X>�F��a:����w9E=>��={+>�V�>�r�y<�<�},>:U�=6��0[ ���,׼�2q����<E>{���r=��Ҽ	(侚��S2��:ξn/~�}�?H��<}��>S�ľ����;����ϙ���E�=o`i��D�>ʑ��G�>��C>NՐ>�@�>ǹ�|%��6�3�<�a�"F���%
���=���<>o@>(�x=�&=H*�=M
 <����FL�>�2?�dt?\o?��F������O�Z��ƾ����*_�>�>zخ>�6�>��=~�'��������� ҾϹ��S��>x���k������>`��O<�<`����A�= p��ʮ�=2-�>/�>_�=�j=5��=��D=�ۧ�y\�=oJ׿*Ǩ��nM��F��Z�=:_�=B�M> �� ����>�>���kiȾ��>��,¼K�.>�`I�����=ޕ=�ξnk�D(��s��ξIp6�u�W��^��؏+�FW�=,�K��Tj�f����s3���z���M�6�澍�o���{�F��>�^�=��=��8>g�?^�'?��?����:�>m���:��=A�>�->*��=v}}>�z���ұ>�V>Z��>6�ŽL���S4��ͷM�/�=S�=>%0>:f�=��=t/>~l>
�����N��Jཻ5;=;�F����=��=	4>(j0=�=�?���@)����F7��H6��w�?�~�>1�>����;K�Rh˾ǖ��nn��'~~:��>��?I�&c�>��=L>�F=p�ݽU�0>;(���;>yK��>->vI>�j�X=��:=�*��2ct>w�t>�D�=%Ã=�=/=���>��?��F?dQ?��V�UH��4��md>������|�i2�<���>��>���>���=oy�fP���<�����2��f�=�튽��x� �@>|�Ƚq�������Ľ�d���(�>�P���=.��>u���>[=�v�:�1��J�%[鿾����q �&{���1�����;�4���ky�v�t���=���i��Za���վ��'���ս�{ >���>�ڊ��N�|'ֻP��9���r#���e���2=��h��7��dr]�0U�<͑��\�9���m����p%D�ȗ��������>�m=~�"��Z<>�-?e�?>F�>i؇=*I�=�Eü��>�a�=�{�>��>��+>��B>-. >r2ʺiW�=�_ ��#�����3 �<�=�}=�cP>U����"=��Լ���t����+��|�oZǽ���i�ٲ=#E;>��2>s/g:����NԾW�!�?1���]�]?�E�=�̩>#����eDb�km��Y��<�>�Q�>^(�<�J�Ƈ�>w�>�G!>���=W��,M�_�l�3��W�2�\)�>������"�=�.�:����աX>W">�7i=`�A�]�>"T7?qh_?�O]?�����#���g�,���*�u����=�#?#�>$>�&�>��8�S��t��l���)��{v>�M�~���
�> "�1�ݽ��>N�*>�s��1{�=�6>xk>�I�>q@E<	����U>�$ ��;=;��ʻ�j/(���"��>�_>~C>��3���ؽ�~">"C�;�;��@qG�2��=�%�=�EP��S�[�ٽj>fվ;�p����=�������D
���]��gu�b�۽��T�==����X�:����&K�����A�iu:�>K��<�<��!�>�5�=ߞ���ㄼ�o?p�??��6>�P>4�T��1>r��+�<��½�$�=�ɡ���=ˁ
?�~�>����O�{�
=�=~�{<�[=>rHa>#Y~���f=T)>��7;~l�z�t��.�>O3>n�r��l5�r��=�<�==v>������ldѾ<cҾa�J�1�t �>X���^>rdҾ�w�=�=���ɾtw���ͽ�e<(�i>�f#����>N^�=<ꆾj�>o=��>r~�=k
�I"���u�2���c=�ه>n��=e$���1(�|�C�vϚ��T��1�>/�?�"�>~�>jB�������ڞ"��� ���6�^[=���(�w>"U]��f2���|�D�v��Y|{�d
>�Z�>���=��v=���f��:ei�a3>jŞ=�kf>�o&>�K �_���޾>5��>��=�nB9pI�#��b�����G(��{����k��j>������r���v��)�ڽа�=��(��{=�A>$��=��=�(g>_�*Ӱ��4���;X��%���oH����׼_��x*<��.����O�A��j�b�<���m���ν��d�c	��z�>�{�>;��=���>�!B?��#?��>jĆ=M�<?�����%?�R��N��"y>!X�>�?S�>�?�>q?8ut���i����<��i��=��=��S>w%>��=,�b=��½���� �xo����=m���>=�(>��>�y>H�=�P�=˾As��d1w�
�����>��޾"G�52��W=���x�Y�6����Ǧ��n)��:�=�����R�>z�g>�ץ=�����`u=�r�>��>cLݽ]��(;ƽ��޽�Qo>��=6�>�a�޽"\ʽ�$4���=�Ň<Hե>�9(?���>���>3|�=�?��������J���U�>>��=���>�;�>#�O���r��� �q�A=�C�̾���<r�7>C��=
�E>�}��N��l��^΢=�S>g�۽��%>�M�=¬�>�#�>�]>�~=&�(>И��O����T㵿���BMY��]���๾�׼6筽3���/��a��&վ����6�:�>�:�>�?{>��=��=����] �� � ��vD��g�i���Q�M�����%���>~F[�ɗ��g��G���2���۽?�6�s"!���U��#�>�� >8W�>Ű�>R±>���>9w'?'�*>M�1?u������>T�=�VQ>�@>1V⼚�>W�?8�>�?C�׽l�y�Rmg�A�����>��Q=�i;>�=��:#}=�b=鶼���k���ν(m&=A�=Q �=^�R=�c->���>��r=z���_��|���Ͻ> ��T,�>��d��4t=�_Ͼ馽�S���q��M��[�������u�����>~�=$( ��q�<�Lh>Àf=���=�:|���*�h�=sd=�t`>ʻ?��*p>R*���/˽�y�Bzx=2Ͻ4>�?.�>{�?�췽����_���
������ü�o�=��I>�(>�Y�2��������!()�d���'L=^�=>H��=ZG>�G���TB�O���>9�f>b�i���?=�Q���5Q>�m�=ֺ�>�~�<��J>H���Ƚ���/�����=���9���t�n��m\=�G��-|ѽ��=�ն��"���l`�$wi�g�d>f�>��C>�9�>�~
>4���]���6�!��d=��Q���h��dN��J!(��4ƾQ �=qNK��W
�D���Yx����Ӿ�w���Ҙ���C�z �s`y>)����v���@>�o�>�><�>?���>�1?I����a�>��=V>�b>��]>%�?zZ?i��>ڡ�> ˚��N�Kj�=g	�5�<=��> �&>X%>�^�=���=����#H9>`m:���j��=�d�=t��=�>s�K>y��>Ҳ���	�}Ӿ��Q��ھ 8"�_o?��=��>=��+� ��T��ܔ�<�
��jn�����]���Ѿ)�>�Bݽȵ>yD����:���=�
����=�U�=�>�Cn�p>-ȑ=:Y<�����c�<�j����=��X<H>�z?؈?��?s�#>�#'����%������Q����>7��>���>���=�r<�ɾ
þ}�����<�d��;y�>�Y����]>���,�iL�<�e>�B�=L�8�v�>���D>�9�>��}>3V�=\��=�d���g�'�ʿ}��J1;����z�/~^<�7>���<~d��4�`>�c�U@J��q�Bf��`��<r��=ʉ5�*��=�:�9f�=L�o>�.����ۼ����Ȯ�a������������W=P�l=����	>'&I�����'	�ޝ���w������>k:�>g�>��e>�(?�Z�>�^7>�\n��[�>����|-�>Wo�>��>q5��$ӆ=TϺ>��*?cg�>�B�>�?�|�L�|�-<��=��>˲�=��>7�.���>z�r��zC�ǹ���放<��w�ֽ����>�;=3Be>B��>�  =E�r�U�#�Џ��YaԽ$�>wĵ�]ƽc���@���H
ľa��z���\��Qxؾ�M�=���9��>rib>j�H�B��l
Q���H>&��<.A��|i�yc	��^�ts>��=5��=����c�%>� >����<Ⱦ��i>S?<�?"�?Ӈp=�74��:��?��?Ͼr->�Vh�k�q>:��>&嘼�ǽWH���$�B|G��^�)�c�I�>JƳ=��=+�>�3��Uu��)	=x��>����>ԉc=#z	���=>��a>���=�� =H�R�<��=����ʿ�w�-gF��̕�x�>���>wc
>�8��w��T苼�3��dE���"���>��E>��>�p�>o`�>�پ�疾5�Y��ѽE�@� �, ���-��&����1�;~�Խ*g���On�����]5��-�+���Ͻ7{���>���>�S�>'�>"F�>!?g�>Gf*=%"?MT>^��>g��=���:5�>�3S>p��>9�?}1�>�֗>P>�EC�����=�jc= �=���<8�B>��>()=~s>�1�=5>�q�\=���')h��(��u��G>)�>��?���/�>��j�����$���%P>�y ?��˼��J�"��>���&�oP�����H�=��?u��>O�#>m�=�g/=���=E:c<��ں�ۄ��W����ɽ&(�={��;v9�h]Q�.���2��=j�=P �:-mg=��X=��6?��2?�q?1�t==���9�<�$J�,���M�8�e>�̾��-<Fs��2���6����D�}>��\�>vc<oe�;�Q�<� �~s��<�Ł>�r>�&>��>>���>�x�>b�>�Kf>[�<�����2/�c���R��X^��w��UDa��4�G�>�a"��F��н�A��������=fڕ>��>̘�>��=>�<���>af�=|��Ӓ����T	��һ�"ܗ>�-�������ǳ���	>�΃��3�{�9�=���s��2��_	��1>��>ZJ>9>�c�>��>�Ĳ>����?{�^>��v>⠇>���>>E*?Ђ?���>`��>��-=����'��L暾��t>�r=Qy�=��>�O�>1Nս)��rڊ�M��<�ν��l�B�5�j���ޅ��e�<��=�>��?����&�7C�-�޾��軨>y:!?K�;�gr�2;�<�½�6¾M���/���6��V�<�?�#>@Ay>�l�=N2�<b�e=VB0��y�=T=�=�Q�=�6����=
��=^q-�˸[���&�E����e�=���=
:�=�\;>�R>�ND?R/?���>�p�z^�,*/���14۾�˾,k�=6gY�N�N�yV��m�Q�W��@��.)��:��==��E>�=���M`=�����X�x~7���=��`>u�=��j=��>^3O>V��>��>��=L >���>�/�����[����o�V�ޞl��rt��=**��F��=��>L�Ѿ�T���U���{�>yQ�>)1�>1�=����������#�7�d=v�e�-O���$��� 0�v����=YW�=��(��Ӑ�q��=�PK��P3�*������<�2��d�$�)�n>�i�>��>�+�>�6?�*�>Eݭ>�@���!?���>^>!5�>�f?X\?�;?���>�$?��=�!�=��?��h���6>���=�L�=JA>yAU>��M�0=�ʁ��e�<*��{����4�I�-���Ľw#,=�S����=�k*?���m�5����nIȾ�:������>��=6�=m��<��%������hv�xd|>^�:>i��>�K�=�E>���=p��x*�*�>��h>��U��*����K��	>���<�D��o�C<B:�;�����}�=|�}>]h�=D�'O�<�%?Y0??gcv���H�9[�;Ϡ������j�+�+>=k����a!��J��|�?�
e����[�=9�@��(2>�j�=�K>�h=�6����q�y�B=kpm>�)�<�K�<�� >��j>w�W>�:>�P�=�=��=�|ҿ9Ԕ��˨�_��6��;K���	��0l��>(`=k�i�x�پ��=m�<���<f�>o�=>�F=f:�<����a�H�������ǖ�ֺ𾗅Ѿ�!��S�%>���艀�����O�<�˾C{�����u���ž��7�����Q�ӼU�>���>:4>�#?���>�%?�{�����>��>mA�<�>� ?lU)?�?�d�>���>���=���"1+���3���'>��'>R4I=�`g=�l6>�Ϡ��I�^����A>�B��>u��2W��3۽��"��=�Q�=J�?�a_���0�f&�w����y�P�<��>R�����>Rĺ��@�$���#��;u={ZH>
�>I��>��>	'=���=B���CȰ��C>2O�>�a�=�ܷ��E¾���= ?>�x5��G(���c�&�ٽ[�=���>��1>�L�������1?�5?�+?*�;��ľ����*;vվTt�37Y=�Ț�H5.��M��:�2�)��8�_s3�'\�����r�<p{/>r��=M�\<lU���J��X6�T3�>�3=O��=��p=%n�>;��>�M3>K�=O����Z��Gʻ��ϿGw��������h�v��=��>�7��_zz�Җ�;3/���n=MW*>B+7>�ݞ=-j3>�+�<��[>G�d=�?�༱+�d��]̾�W����>��oi>X9�kaL��Yþh0�=z���,=kֽ��.���q��tʼx���>7��=�)�=C��>2\?�*?�(?�;��?�oR>>��>�(�>�s�>�.?�X�>���>%	�>[�>�j��ƾ��fi�>b �=��]=2ॽ���=߄�+ �<��?c��v =�m���B��V��!6��VĽ�s����>�k*?���m�5����nIȾ�:������>��=6�=m��<��%������hv�xd|>^�:>i��>�K�=�E>���=p��x*�*�>��h>��U��*����K��	>���<�D��o�C<B:�;�����}�=|�}>]h�=D�'O�<�%?Y0??gcv���H�9[�;Ϡ������j�+�+>=k����a!��J��|�?�
e����[�=9�@��(2>�j�=�K>�h=�6����q�y�B=kpm>�)�<�K�<�� >��j>w�W>�:>�P�=�=��=�|ҿ9Ԕ��˨�_��6��;K���	��0l��>(`=k�i�x�پ��=m�<���<f�>o�=>�F=f:�<����a�H�������ǖ�ֺ𾗅Ѿ�!��S�%>���艀�����O�<�˾C{�����u���ž��7�����Q�ӼU�>���>:4>�#?���>�%?�{�����>��>mA�<�>� ?lU)?�?�d�>���>���=���"1+���3���'>��'>R4I=�`g=�l6>�Ϡ��I�^����A>�B��>u��2W��3۽��"��=�Q�=`ϖ=�e�=A��.�m��� ��t�w�ؠ?%�Q>��=YO�\�<^f6���Ƽ�>P��������Rq=�j����>��>�k%>�7ֽ�*��%��T����>=�t>Bb�dSu=6N����=�*T�K*O���5=�_4>��M�5[�>+
?vU?�f?ݗ���ʾ8*�6�������	>���=Z﫽�C->�*1��}��Y�<�� �(�Ⱦa�;���)=��S>���=��R��X�=B���n��4q�>�G���ٌ=�M�v�q>��K>��>�g=��|=�^a���4>b��������*�����h�����id=r K����<W[�P�w�l* >xI=�I���q���=k������0A�>� Ӿ�����m�+���˽��E42�{d�6�]��㼆Ʀ��4�0eA�x]�@>#>��_��Vh�4�z���I�%<�>�H>��z>��>U�>�c�>Ru�>/s��zH�E�k;<Q�=:p~� Q�>V�>��<�4>�W�>��=>x>�ͽNT���ƽ��=�>�=�]�>ڥ��.|��ؖ��h�=}�=��ܼ����I��e�i<�P�<O�_�w���h�>�A >����RJ���.�����h�پe,�>r�&��9� ߾��W=�)��� �����-qa>Q��٣�:�!��љ>ȅ>C/>�6=���6�<,ս-M�=M����/!��rF>'?�;tн�=hc��0r>��0��S���+�؉�>��!?�?��-?\��-,��[�ﾏ���Pս���/߲>-��>P�>̺>z�?��I�1�оJ�㾱�&���<8�>B�7�T#���|?=�<d݉��������@v=��(��s�>4��>檉>��1>v�=��>7>R=v���ճ�w���G0�A9���U޾Ľ=�C������nRn>_P��<������+��=dy%=�����/ԾP�0>0�e>�~�;)�^�e�s�Sؼ^�x��E��	a�!��j�J�">��ڽb�������a��� ����.�м����dǽ�?�>!�M>�ϗ>~��>}1>?1� ?"P�>c����<>�>�`Q>�͛���9>�s >I �>��,>�l�>yH?u��>����|��/�E�+�=p�9>+�0=��J>���=*�>Z	�����}>��SC�߰���{|<���1�����>��E>圀>�G,>�ۻ��7#���/��ȍ��d�r��>���U0�K��R�o�ھI����T��
�>D���)���Y��1�>�#>��>(">�{C��X��n���S�0>��>4��<��<ď!�1���n7>��	�"���hԪ�)�Ž�rȽ�ѧ>��+?�a,?.��>Gco��Y4�~%��#�ԛ�� U�-?낮>J��=�3>�d>{���d��Zؾ�n�?@�=++�>�~�l�5�<$=p�f�F+��j8��4�ܐ5>l)�<XE�=���>Y�+>p�T>Oj">�ּK��=o�=z��;��=J��&�F���g��=�y>���<]w2>��@�����g�=�c�=a���A�Mk�
I�>���>eҍ>y����}���1�d&���˽zt-��s����< .�K>���"��T�=��-�$�Ҿ��'��7�����&�g�<4k�Ņ�>.Y�=�>U��>&@(?��?�?h6ͽ>��>�ж>og>����p�;>�Ԗ>��_>�x<���>!'�>�'�>S�������Z�Ap�=��=��<>��>ᑈ�q���M���-1=��;�{6���y�S�X=ƕ���V�=yU�=E��=#��>�h�=� �������t��M���4?�:��5g��4�	�3�=������w���:�9y����Ǿ���Y��>��=p�%>ɉ;����U�����в�=*VZ=(E�A(F>�1��&U=�<>����j�=+C����<튼'<�>W#?���>��?3�Y�����R��eپq2>���J�f>�p�>�D�>D�]>��
�	:�g¾8ƭ�p�i3'=a3�>��c���_�K�*��v�=:���ٽb�Ľ�΀=�,�S�>��>�L=�#V>�l=R�>_�����=z￡�	�C�_����P>��>(kc>ø�����Ҏ�>�}->�ƾ���,Vپ��>�	?�½X����>E�M�C^e;��=�ռN�,�!���Q�q��<b����3��m��������V�r�ܽd44���|� S��'\U��`��Я�>^�?>f��>-��>�]?7��>�	?ʻ����>��a>��e>��$�5>�i>�]>̿N>'?82?���>%��������$�|�>��S>f��;ʵe>p �2�=޻�=MX��xb5��T��Ł�t�=8�;�R>��>�@�=�.?>�E���E���;��+]��Ꞿ;��>c߇���������1�=i���ӷ�H��}	�=��
����%ɫ�r�>��<>�:h>A�=�%��e� ��Sܽ��>����T�R|�=�뙽*��<��/>I��=X���K\��E.T�B��<z�>��3?"�C?u��>kϽ�E��L��>�m��2��%q?�ݟ>�/�>���>���.	��ھ}�ƾd�9�������>��=�����9>$��=t�=x��rX>x�O=+��C��<{uk>�u�>��>��<6s�>���=�D;��ݿ�ծ���/��&�<��}���3p>U�(�нO���<��-���PX,����4��}�q<�X�= �:M�">�񤾰����T��O߽\�c�H$����q�����
����ս��}=������������=>���ʿ.�kt��;��>dr�>o�>ꛝ>E'?Q�?���>�D���?E2>O�q>Z⽼!�= �>��>�J,>��?�	?p��>W䄽�uv�% ���-�=�%�=3x�=�>,J�< �>R�=�%�K��:�P��^���սjʼB��=��3>�z�=�g>u�������Ƚ���U���%������?�᡾�s�>�F"��o<��O���A�� ̾����{��>b��>5�(>_��>v�>�a��Ȃ/��5(�}�P�=�<���=��J>��7>���<�t�=�A����|��)�`�$�0��,���T�M�>16?O?v	?]���뾭�P�Q��=ٹ�>�˾"�>�7�=]0�>���Nt5�Y��H�E�ʔ�'��=��޽sG��5�*=��
=rMO>��B>�Z��j�,�t�B���佖L�����>:�@>���>�/�<#�9�7������e��㽿ӑ�bz�3�y>v��=�������s��)^<%' >�P�����=�?v>��]>t�P>A�>��<���='�^����g:k�JR������� ��q��{hm�����M=(��rܽ������"*>�;Z���=�
)׽����ʯ>�66>�+>��;>�A?E�3?�F?��վ��=�����!�h$��?�>��+?�$?Y�?���<rS��c|�.���s�E�=�1>��=BT�=���=�V� ���1=B<��=C��孝�Y�G;b-��.�(==�Z>-i�>5q�>��u>������k��?�>�'�3lľ^�>I)�>z�v>���>���s��ľ�ȟ�M�c>g�>�(?��3>)q>X�9>���EQE� t����1;<R>����>�5{>���=n�S=q  �TX�<n��<|u>���)�¼�k��<>�%?��>N�?�`.�MF׾���f=������;�6�J>D�d���`>6þ�Q�DT�0�5��ڲ��6f>�z����ɼȠ=� `>�w�>-�*=��>p�<��h�sj��)�=#�=C�i>��P>u�&>�b2�K��n]��G4��6�99��!�����#���Ž�gM�t۰=�?��V]���E=����T����P�K��>�p�>T4>C�>�����=��G��L=='>R�~�\��&��ڙ�{U�l��=�E��	\�nX�h܇��_��6����?��=�X�d��5 4�mS
=�#�>D��>��<:�=Q�o?aF@?�3>�Ծڷ�>Sоƕs<��?��'?��?�g?dז>I��������r�{d��=S�">���=���=S.s�*�d��2<#��= �=��;`|���>�������=%��>NnR>��=|^�>�l>�]�@v��õ-��3����G$@?*�=3��=^ߠ>����/�����!ʾ����� ?n�>�_>Ԇ>�c���)����=V<��$��;Cu�E>T�7>������=dc�;s~�<(�<H�<���V�p��p"����>��<?>M-?�*?v���-^����۾�l׾*V�������.=l��ob�>�*:=�(��n�,��V����!�n�M�Ԗ�O��>x�>8PB>��'>��X�2b��r׾f��oR>�X�q�X>�S�>�>ůE�t!ս��5�h� ��%�Ѥ��5��I���+��C�=�(�>��Ѿ��#��"W=Ō�G[>NF2>���E�h>�!h<h0��z�����W=	�<�q=Ur������վk`t��G:�y���|���>Ɓ�����
���I�D�<�m�2����½	˙��`�=)�>P��>�{�>��>�o?��=?0M?
�;��>�.<}af��">�1�>�_ ?I�>t��>�>�P׾ڑ��b�A��֠��� ��!�<��2=W��=B>��=+��=���NM=?�.=(ۄ:��:�wJ��X�>��>0�@>x�5>���>噼Z�����=�:?�����I�<˛>�y����>~}+<0����$c�`@��oþ���>6�?;.?��
>�j�>��>�o>n�$<��3=}e��ձ=��>�0=�I[>��[��c== �=<� �x	�ɱ�N/$����ٺźC��>��-?��<?Vn�>*ښ��ā�˫��ox�=���.<�=�׏>�	��"�>i=�����X��7&��y��5�B> s��[�=%��GF����]>���=#�j��=����*5\����=<��=[hB>hd>��M>�PI������%��?:�D0ٿ���jAZ�K�E��]�>��2>V酾��,����>�������>X�t>�q�>���>12�>�Y?>�λ�i�=Art�͖�vw��A޽l �������ľ�^z�����a����,��;�'|��0�U�������&d�<���>ҽ�>��>�L�=��4?�n?2�7?l����">HJ���A�=^dK>�.�>g�?D��>�w=Z����Vq��G۾澞�L|i�[�=H�H>��3\/>2�f>���g
>	�r=`R�=4�C�&����G�f=� >���>� �>�H�=���>p���� Q�=�H#�A7�x'>@�>����>�w��)L����n��p���TP>�c�>`��>h�>:~�>>+(>����I꽰����F/:*䩼\ S>x�>���>��=�Q=4�=���=�x�<K��=�ܴ=z�>�-\�.k�>,�3?�?���>�hW��P޾Cp���$���	��`/��n>2D�=��>�\����⾛�'��������Ź�2d�<$�	>�,�@'ν^�s>������;]5�=�Z#�d�u�r�KOf>-`�>]2r>���>�����lǽ�1��,���2пzL��o��r��_�=�B>p5ƽa���,���>����=��=�C,��g�>僩>�矽�뽱<h��>�ʓ��)�t��3���M�l:��ԁ�.�W�d?��q0�;<��������}�����~g:�,X̽q��o!ּj�1=��>;�?�H�>Gp=��8?YE�>3�>*�׻��>҉Z��Q;�:n=Ǝ?���>�c�>���>nV=��/�$���8�FF$��+�>b��>��l=��>�M>���łʽ��7*=��s}���F��q�����r�������=$�>V��;+C��c�w 0����xY>�G?��E=��>�q�zh��=,�?O �U	)��,���{Q���|>�U.>�`G>*k���CV�Vŋ<uÁ>��H>���=���= ��u5j�hyo��2ۼy0=���\v����]��fh>AZ�=�ٽ;@�=��>�?ب?͔�=����s�澻n�g.ž�Ij�Oܢ=�:�>dR~>
����*�@���1޾���,����q�t>�N>(��5Q'>{�K>A��]�㽔��=��3;�C8>�̐>��>N��>�	=/�t>�JW�ۆ:�o�k���߿E���B��p-��+G��m��Q�=�t����=N+�=��m�)c�����ҹ�=���=�>��}>}4�>J�>-�ν�:�=Ii)��� �Z��p/���������ˏ�����ag�G����o����S����&�BS"���44p����>?�>/�>��>5?�(?f=҉��0�=��ػp#�>�3�>���>R��>�>:�F>�H�>Ѐx�ϝ&=���� d�"�>�I+>m6���ȼ��%>�;u=&>	M>�}�=?4��h�gv��O�:=�8�=ϳP>�a>��l>���>��=1����n`�_��=����ᕶ>�3o>�=��c�ž���������R���QP�X���OEf� 5�>+��=%�$:��H>��=��o<ĳ���&=�yS�����{��=�]c>�Y���T:���Z��@y�G<��,!ѽ��k=5R�>�$?f��>�*?��J�8z��	�c����پ�Uƽ[P�=��=�j>�뒾����*!�ܾ����Iž8�u�_^6>���=�}=(�=��<<��<y�j=`+>�]�=6v=�dS>��W>K��>,Xf=�m>o[�;I� �����[��F���A��s���ӽO��=�����<�����&��Wx����"���%>�[>>��^>e�h��>D��>{#�f��=���l���U��)N��T��7X*�a(�Cf��O�(]��� �Jᙽ�)A�44�pi!��؃�ؤ���~�>��<�5�>�J>��*?|��>EI?�fC>l:>���>���>N��>�k�>$x ?�@�>/��>���>���>�q�>�٢���B�����N�>�7>�O> jJ=la�=s���G�������\Ԩ�[=��=�e���rC>w�t>N?>�)g�2�
��d�>J��ھG�>�l�|���b�R���
�<-� �6���F<
4ҾO�l�쾚��>�> F�=��>T+2<"Y�����&��i��=���,2�Q�7�b�w������p1�F��U���IԻ�oI>�?N?���>
�|>���_�(�Y�7�����j>KV�>d;�Nc=V󎽙�0���.���V���d�>t
<��p>$�˼\�P���I>�/�>��h��\f�G/>�t˽�d��:S>f �>�>��/>u����=�z�=W�=���-�����Xc���z��P=b�`>d@>AՂ>�c�97�]��#�=B��=�>t�c>i��>{Q�>VF�>O��>ɪ���Q�p�I�0��/װ�D�����[U����7���	=V:M��1��+H_�C�����Y���W6��1���)�>6_8>{�>�`�>�A?�
?>m'?s.�=�#>����V>�W=IC�>K��>
?��>���>nՓ>"���=ƽ�d��ܤ=�w>�)=,�����>�>��j=��@��.����:×=zZ�=V(�= �Y>�'5>0�4>�H�=�U?�D>��J�[@�`����z=����h�>��q>)Ӽ&���x/;a��{��iV@<��$3��C�=T���*>m����<&�>��W�2gb=�4�=CR>�ݑ��g��ŃD�G$̼��I�z@U�Eaɾ�wE�4=��(�!���)�=�/�>��
?�?\O(>���w����~���þM�N��7C>tHh> J>a�=�<��Z��n�����Μ�K�H�v2�=<&)>�yݽ�2P>Jn=�<o��;�> ^ɽA�l>��6<��>	�>��=W�>P=2揼KL�<��ҿ�HV���Y����|�ѽ�B��5��(���@��1y/��c����ֽ�'>e�7>ΧB>�^c����;�T=��>;��>�sM��95<�1�%�����^9�;�ռ<w2�(`��U���/���F����+>�������;�4�������=�o�>�K�>��>2G�>�?G?}̛>��>���>��>r�<>R
�>%>zH�>�>GT=?�4�>��>bu��H�������(���<��>�eN>�_�X���o>�P��T=����'�u�y(E>?�N=P �=�5�>&zh>�$�>���>�@�0ɾ2�j�|}�!
��f과���>��j�E������CS���������J����E��h~�:���6�>٦�>�u��:>�Kx���@��m½�&�<���j0I��M�=[��=�z̼��������Ez�����N�
���[�U��>-�0?��?��7?�v;�U���5�&u�����e�>I�O>tNv>ɑ=�3��Dz3��3��5������-H�=�a>��u=�� >. ���,A;3c7��H>!�,>Y��=H�=H�f>6��>�G>�b��=�*>$/�����ؿe���z�Y�X��]^>J3�>�47>�$�> ��>6u�=��ྵ`���=O��<�>��>�q�>>��>��>z�N�]����R����W��H+��\�/��ٓ���H,��V�W��l���`?�u@M��tX�� ��.t���Z��ׅ���m�>�P�����>�0>ϲ�>�&?QMO?W��>=��=�I ?}��>��Z>��>W`$?�Y?���>�Q ?�U?��>ϊ��~���Fu�#�?�ܸ>N|�>�e>�Y>��=��=/}�;��Ľ���/r���6=؎b>�k<ͬ�>+.�>h�>O��emL���3�N�i��&��&�g��$�>�{���q���L��kǾg��y���վ!� �f[�L�B>>�f>�S�>�U->�v���\<\u�=��:=�4R;iε���4=V1=����3޼Ub�`�:��Z����̛�@S�=E9>���=�4E?�7K?c�9?枼����Sw)��B/�{�ֽ���<#=?���*�+��������E�	���о�L>Y��<�>=m���;�<Q���+?-�W���f>�=��"�b�u>̜�>�0>�}�=��>\�C>��>�K`��2���[����̿Z���Y���<�r8>0�C>z�R�G�@��D�1���N�����x�=<�:>�_>�D>��d>��!>	>���8]�^Gܽ��/��*�"Ȝ����RG=#Ǒ�iS�����Ga���Z�WvV�]ߠ�p���z��ӫ���{\�Ā�>H�h>�4>o�6>k;!?�9.>
��>�C�>2?]��>��>3�?C?؅;?��+?�9?��<?�=��� �ƽ1 �d|%>	0=�k->�tT>��>�݂��Jf=7>�(���G��ܷ�<�!���	<_#=NfA>��w>��>ha�<<�9����|^�f=��վ�N�>*�=�Eľ��C�钎=������x�����������L?�	?�ܛ>Z�>��=�\k=�R�<��U��=
��hR$�&%d��Jz�x�x�����������B�=�-<ٌ'>M)p= m�>Z^b?�/1?�vi?gc��$ ��7�)mC��J�a���D�%> ��^W���뾔���3��BH��O#�y
,���u�\��=����>B��{�=�J���8����>�n�="C�:��?'�h>:eU>T��>���>��=�M�<H�2�b��Í��r��������'���뽛��^�����<�J�>�D?>�վK��9�B>#�C>�6#>�>�,�=V�T��M�=�Pa��2+�x��l���	���<i�mI���=v34�?�	�3�3��)�UF�������~�%�XJ��X��g �>K0�=���>���>=U?A��>�+?g�=؅->�D�>�Ζ>� �>�>?)/?7,?к?�?)?x݅=�Ⱦ]&έ�5�RC=��	�@*�=�PJ>J�>��ʽ�<�=�]�=�P;��0�s7���O<����������6==�?>h�>O��emL���3�N�i��&��&�g��$�>�{���q���L��kǾg��y���վ!� �f[�L�B>>�f>�S�>�U->�v���\<\u�=��:=�4R;iε���4=V1=����3޼Ub�`�:��Z����̛�@S�=E9>���=�4E?�7K?c�9?枼����Sw)��B/�{�ֽ���<#=?���*�+��������E�	���о�L>Y��<�>=m���;�<Q���+?-�W���f>�=��"�b�u>̜�>�0>�}�=��>\�C>��>�K`��2���[����̿Z���Y���<�r8>0�C>z�R�G�@��D�1���N�����x�=<�:>�_>�D>��d>��!>	>���8]�^Gܽ��/��*�"Ȝ����RG=#Ǒ�iS�����Ga���Z�WvV�]ߠ�p���z��ӫ���{\�Ā�>H�h>�4>o�6>k;!?�9.>
��>�C�>2?]��>��>3�?C?؅;?��+?�9?��<?�=��� �ƽ1 �d|%>	0=�k->�tT>��>�݂��Jf=7>�(���G��ܷ�<�!���	<_#=NfA>��w>��>ha�<<�9����|^�f=��վ�N�>*�=�Eľ��C�钎=������x�����������L?�	?�ܛ>Z�>��=�\k=�R�<��U��=
��hR$�&%d��Jz�x�x�����������B�=�-<ٌ'>M)p= m�>Z^b?�/1?�vi?gc��$ ��7�)mC��J�a���D�%> ��^W���뾔���3��BH��O#�y
,���u�\��=����>B��{�=�J���8����>�n�="C�:��?'�h>:eU>T��>���>��=�M�<H�2�b��Í��r��������'���뽛��^�����<�J�>�D?>�վK��9�B>#�C>�6#>�>�,�=V�T��M�=�Pa��2+�x��l���	���<i�mI���=v34�?�	�3�3��)�UF�������~�%�XJ��X��g �>K0�=���>���>=U?A��>�+?g�=؅->�D�>�Ζ>� �>�>?)/?7,?к?�?)?x݅=�Ⱦ]&έ�5�RC=��	�@*�=�PJ>J�>��ʽ�<�=�]�=�P;��0�s7���O<����������6==�?>��>�����|Y�3��WkV��=�s���UE?�B��gz��tT>�ýKKp�&.P��:�������Qd�=k��=�8�>�:?>��/��@۽B\�=1���q�c=J�.=��>c�=HY�,��T��J�z�(N����>=F!	>�>��u>&ֈ>� ?}�:?�P?���=放��I���)�����6��_߼)���; �<$������ ����E��ݷt���<�h>���_5>'��<;ͦ<���IQ�=�X��m;���p>��Z>�bj>K��>*��>8]>�@�=M�/�������ܿ`I������ʑ9�����ap>��>ϩ�����h?���I���:?_>7�{>z>�ϲ>}�O>і/>��>����R���*�0����ľ�y��P#��[�=ɹ-�SHp��)D��c���C�l��Yַ;k=��c��[M6����m�>�3�>�H>�z>E'9?{�*=��?PPC>jU5?���=�ׅ>�X.?��?��>A?Wj8?�l5?��>bc������E	�TJ�>��?;z>��C>��>�`���V�$�>W����Q]/��Ԅ�K�$���'���,�k=^�>���>�>>/7߾B�>����kѾ�ZS��2�>�R�Q�=�|�|>\ ��o��s𞾤�ԾF����>w#�>��6>P�>IQr>sު���3����<Y$�=3xO=5��=u	}�B3d�6��=3Un>��>�����װ�����	�<pW!=��=yŘ> ?��.?�UB?+(������5#<&}+�y�=<���<9^9���&>g|����w�ؾ�ƾ�p��a���Z=^r��0�g=�e<>I�V>�@u>65��gh�<D9C��4e>��*�JD�=�2�G�ӼhR(��ڼE�>b^8�]#�=�(��wտ�w��o�澠�p�q�>p��>a�۽�Ir���}=�L=oq���f��p/=��< ��>���>	L!�y��a����9�:>�b�=�R�C�����Ӭ���;=X豼_^��E�:�rD�p���g�ܽ����/b���I�!��yn<���>��>^��>��j>�>ɬ�>ѽ�>O��c�>Tg>��Ǽ�e>ώ�>鸪>�??�>��=�n�o2��-��x)���\>�3>u�4<�)�����=�;y߽vz}>�'�]u���d̽�y�=��>[��=�t>0�Y��������>�>>/7߾B�>����kѾ�ZS��2�>�R�Q�=�|�|>\ ��o��s𞾤�ԾF����>w#�>��6>P�>IQr>sު���3����<Y$�=3xO=5��=u	}�B3d�6��=3Un>��>�����װ�����	�<pW!=��=yŘ> ?��.?�UB?+(������5#<&}+�y�=<���<9^9���&>g|����w�ؾ�ƾ�p��a���Z=^r��0�g=�e<>I�V>�@u>65��gh�<D9C��4e>��*�JD�=�2�G�ӼhR(��ڼE�>b^8�]#�=�(��wտ�w��o�澠�p�q�>p��>a�۽�Ir���}=�L=oq���f��p/=��< ��>���>	L!�y��a����9�:>�b�=�R�C�����Ӭ���;=X豼_^��E�:�rD�p���g�ܽ����/b���I�!��yn<���>��>^��>��j>�>ɬ�>ѽ�>O��c�>Tg>��Ǽ�e>ώ�>鸪>�??�>��=�n�o2��-��x)���\>�3>u�4<�)�����=�;y߽vz}>�'�]u���d̽�y�=��>[��=�t>0�Y������>�=)D�=�G3�_.2���K�>lӾ�C�����>x�<L� ;�Y]���������3���n�=R�=�ǭ>�ю>J��>��>YK�>�8O������=r�>�� ><'(�q��=V��=!B��ZZ>��;<u�q���4	�WU�q�t<-�m=ޭ�>?�?�?��W?��˾3�ʾ����9/��i8�U��<�=�I�>�W==��0=!-����	V��⩾$#=G�㽌2&=/��>o��>2�=o`A�l5��Z=��m�����c�2>�ǀ�~����=�<P�F>�yG>��G>���X����?࿒O��������s����p�<x�f��o>VǤ�������v�9��:н�A$��$%>|%�=-y��LD�BP���1��k���E� Sо����l0�!N��yiJ=-7>1�N��V7�]i�<_\J��de��þ[�̾jʾ�8L<�z=��>���<��>��>�(?�]"?2��>hϽ_pV��3>wL�>�pA>�"?��
?�EU>->�iJ�����g~��ٽ}��=u��=^r�<aIF�S�>�A�=ȐǼ%��E�=:J����P=���=ѱ�=~;�=�=֡==��f=�4r�߱G�$���@��b������5�!��>�㨽���>$���'�Ҿ�^�����F�(�(8w>ĩ?yH->��>U0�>�(�V �=�C>���<L>޺>=Qo��`�=w]p=��/>��=�>�ػ��{��s<�Ъ=%�X>hC�>|�?�??H?��f�s{/�.��y �Q���6>�^�<�jc>�gݺ�|>�E����������6�==u�7�C��=�8�>Cď>��=�K1>��ƽ|�T����=^�a��"ܻ�������I��8�7>vǛ>�#X=1����y��������� _-��о�Qؽ�!�=�Sq� ���C=����N��������j�c�Te�#d�l�>�@>P2�=�b����ɾ ��C6\�Bo��T¾f-�W�پ�;�=�o>��Ͻͽ���R����z(�e����ˋ�!���^� ?��?��Y>A��>�6?R*?��"?9�=*r�>W�(>&�ἄ��>�?��?y�?^L�>�lb�Uꟾ��<����?;�t� >��8��桽N Խ� ->��8=�<!��
�<�����c��\��H�=��Q=V�=�4�=T92���k����>�>>/7߾B�>����kѾ�ZS��2�>�R�Q�=�|�|>\ ��o��s𞾤�ԾF����>w#�>��6>P�>IQr>sު���3����<Y$�=3xO=5��=u	}�B3d�6��=3Un>��>�����װ�����	�<pW!=��=yŘ> ?��.?�UB?+(������5#<&}+�y�=<���<9^9���&>g|����w�ؾ�ƾ�p��a���Z=^r��0�g=�e<>I�V>�@u>65��gh�<D9C��4e>��*�JD�=�2�G�ӼhR(��ڼE�>b^8�]#�=�(��wտ�w��o�澠�p�q�>p��>a�۽�Ir���}=�L=oq���f��p/=��< ��>���>	L!�y��a����9�:>�b�=�R�C�����Ӭ���;=X豼_^��E�:�rD�p���g�ܽ����/b���I�!��yn<���>��>^��>��j>�>ɬ�>ѽ�>O��c�>Tg>��Ǽ�e>ώ�>鸪>�??�>��=�n�o2��-��x)���\>�3>u�4<�)�����=�;y߽vz}>�'�]u���d̽�y�=��>[��=�t>0�Y�����j�"?���վ�;��LE���=c�=��>�,a>m���xF���ɾ�%~���Ž���<V��>�!�>K��>u�>���=4>�>J����=���=�@,��,��{�=N=��5=��$>łͽ
����;!�;��쿽.T�=��>�Z_>rw>L?q�? '?O�>�I@�5A?��*����������>K��>A!��r���L,��|��;2	����i/s��� >Ho�Iۻ[�=��=P�u���+��?�=��N��C���;L<��>��&>N�.>٧�=�����&�1¿W P��o˾����g�� ��ʹF��Ò����=���<���<�w=6X
=Y�<�� .=���;���=(=L4=8�D����'r��l#j��3��|��3�yH��^pټ�<l�6�ؼm[e�,�"����
���ٽ[r���۽lB�>�-�>4��>!�Tt�>_3?7#?I�h��V<  �>�*�>��B>�P�>{h
?'�>dT���9�ˌ�`.����-�����Y->>� S��P�=�g�>*�6sƽ�F�:K��=�!>�Թ=���O�<�M6=Gg��ם>��l>վ*?ѭ�����C�@� ��6��=�AN>]�%>�u��Qs>�n$�g���ܪ�������m͜>YG?>���>]Y�>ڒ�>�x>�q��
N�=/�=��a�{�E��<��!>s��O��;T8����ѕ�Z�-�s<=��a=�4�={��=)�>�S:?��*?�%&?�̐>��4���N��� >İC>�1�A�=�1X>{b�>�4����ؾ��<�J++�Ҥ	��k�<�z���h>�S��������=�1ݽ̼�=������=P�8>�I�=�M�=eh�>2X�>�u6>Wc�=���=�5)��X���!���<����!����Ӿ�j>L�c>��ҾU���>#�->�H4�����j�>��;>��F>ƀ=V<���=�fu�R�����=�kw��޳�b��l������ֽ�"��
'���U��۽����$�5�DE+�������Xǽ$o>�k?j�>+��=�-6?�*�>>�B<��?W�P>�+�>��
>��>�??�t�>��U>,�>A�= ��+S��cžT�/>�`>zj�=�:�>�F�>	u����[�_�����>�u=������<��-=�qP=��3���:>vΊ>&b"?�����O������q2����;��>g�/??;ܾ6�>���|���!�8t �D��=�?S?¥a>ښ�=i�>+�=+�=�?��2��;��>�}�<�>�43�A��=N 4�~}K�
����cmp���Ѽ�s�=�g>(ԝ<\	>ܐ5?��?�P&?�s?~$��p�,H�ϡ�>$�����=l��>ݑ�>좇������0��cE��1�A�_�|ͻ�T>�c̽�)��.y�=��	c½q=#I>�̼�8(=��=k��>��U>*��=�L(>U�Y=�W�^j�E�׿J���i���\��DX��z����K>�p����g�=�Lý��ڽ~i�<�^[>+�L>���=��=�4`��A=�m����;����_��[P̾���U�k����į��1R�=�ݾ��C���轍��M�K��`p�!���R"���YL���">#& ?V��> ~�F�>�?��>�><j��>���>�k?��C���>O*8?�>���=B�X>���>�L�Ǽ)�暾��f>���>��>�!Y>�M>�����;w�j����>��=-�u�X�>�D�=924<��<��=$�>a;1?{����T-���=�3;�iz(�.>�>
��=")z�;;�>�����f+�|'�c��=��>z��>r7�=�c�>S�p=Y�>�G>��=haȼ�#�H�`�y3>�� <�/ٽ*���F���S�T�8���:��I���F��>ω=͏:>��j?��F?ꕸ>�s�>�Z��n�4��]v�=; �̎#><��>�?�>[f�<<��>�m�7�W�#�L��@<��!e�=�K����a�'�;���=W	>���y8�=���=l�->�ܜ=�ɣ>�Ny>'��>Y�'>w��=O����D�1Ѻ�����5dԾă ��;;�z=lɎ>Z�;T�྿V�=�ǽ#�Խ��ǰ�<y�=��= 8w���s=p�=���=�̽�e���v���V�2E����)�*���M���Xw=���!!l=�������;lֽ�����O�v�t�����~�{>�*�>���>x��>xO?n�?���>C֥�y�$?�U�V�"?Fu>���>!<C?L��>�9�=g��>}-?Q¬�����	þ�1(>���>ŷ4>a�>G$u>��V�$�~��w�6>�g�<�;��E�={��<�`Z=�e=�G>�C>?vv�����e��Ee0���E=��>&��>��>���>�����-�׾�Z۾�9F�Vxa>(i>u�s>e�>�S5>�6=漄i=̡0��B�=/'A���x>�.�=�q�<���=S�޻�6X��/T�׶�<e��=�=):�<���=���=x�B?U�H?��!?�ð���:�4(�{J#�z5۽��Ѿ�<�=G-�>�B�>���rD#�n�D���D��M���1 �����R�>�O��n���>DM�,���PA��h)>;�+��2&
����O�>9�>�'>�8�<j�v����<�쇾Fj̿�D��!����M|��<�=DW��D�>��B�,���Pw=4jq��.���.�� ;�ܴ=�b>%�>�
d�\�<=�=|�����N����!�� ��1M��H���) ��#����S�3a��IM�;m)5�w�0�{<��@���[W��2�> ��=2�}=.>;�?9G?��J>��*>��Q>`��,�?߲>%d�<���>�k*?�-�>�:�>&�=�i+�N�5�.뉾i-C>_-�>/@k=���=S_�>T�;K����<���=iN=겋�祊����H �;?�">Q�>dɉ>-W?������=����6%��W�4<#<��(?������޾��2��⬾�d���>���>7M���=M��>���>ʜ�>0�=���ڙ�=l�=��<��\;����8��{�׼�d��誽��*�ŉ8��2C=��!<���p�?>�^�=%x�>}�/?F�>d�>Ϳ��ǲ�
3�ͷm����4F=�˿>|I��=I0׾R�������/d|��D=�N���7 2>J��;����S�>�3�=�"#<m1J=s~V=ߢ�<F{�=̌�>�j�>�k�>7	>/B=��	�!�}��w��"���k<�G
��*���>����׾.�=��>O=݊6>;�C<3%�>��=���=D_>.O=%~>� �;v^=r�=IJ�����M��2 �����=����w>���{��U ���;��)��U#C���R�����d�����6>U��>1�?@�>�!?���> ��>!��Q��>��>���>�hn>��>1�C�]!��0��>��J>B������w�1���x�� �={�b>���=1��=�>T
��r��=^�=^
�=ɹI���#��O���e�=�UL>.��=E$�=D��>n#꾸������%�D����uʽ�!#?�M�,p��n��9*�񒑾����}O��oD=���>�\�>�Ni>��>&>@p��56�HM>��Q�uH�=8,>�R��ja9�I>���=�t@>'�==h�!�?���L�I!��*�=�&�>P�Z?�q�>a^>TG�=//��a��'о:�3��B���%>E�	?���==0��PN�	G"��sR���Z�M��;���s�>��>���>�2>�`>�>��<��K�>�#ǽb1�<�%>4�'>4D�>�t�>���>���=����Ͼ�,��-Ib������]��/��:�j���b���.ɾ�8v�,�� �$��H<�Z>=f��o[��|D>��X�'��w@��H��=�x8�����ڂ�U��d%	>;�>��n=`y��k����Ծ�2ξ��%�o���Y>���=�S�=�q�=v��>ݙ�> �?A�?&��>�`?�4�����>���>XE�>���>�S>ږ=+-<C�>9`�>�V���b\��������+m=�����0�<��r=]f�uEe��|<<r�n�f����o��2k̽2S뽞B���=��B=��k=�7�>�E����ƾ��ξ�D���)��&��\,?��=>��>�e��
ؾ]׾�1P���n��x�>h��>�A�>��>�}>>+>=3sK�8��=wI;=�)����=��=�'����=u:��y� �ͽ�$������8�=(��=��>�$�<�ߦ>
y:?�
?N{=?�a�=�qD�w�
�1�/�.���"���
�>�+�>>�}>?�v�s�񾤘<��Kݾ:����@�o���=�>NKl��,x�[��=!;>�@���P �<�ב���� d�=��>�L�>�_�>R�R�q��F��� >��7п�c�����+�վ�I<J�.>��9���,�Ƶ��`����R���<.Ӡ�`�5>��2>4F�=�7�]�����S!`���+=���C��vՊ��Q���e�>��=x7��Z�������/���t��fX�rc�bv �Z���� h>?V�>��>_6?m�>+?��+���>���=���=[�>���>��>�h�>;��=~](�Ϛc�����k�lS��Q6>���>�s=�L>��=����rt�=L? >J�H>y��=���`�:�7���ir�=��>�l�=TA>�  ?e����Ǿ\־��,�Kx���l�R�1?E5���G>��9��b�E����xl��oM>�ϭ>8�>��>�ڝ>B]�>��=�N�6�,�[_�=���=�|�=�f=k��*=#ʻ��̷=B�=2�*�J���~;�z9<��=�m�=T�>=i?p��>�
�>-�5=���s�j���Eսg�վ�E>p=�>���>q�r���>�-�s���d��� ��d(��V2>#NK>r>�>��ټ�R���sV����=-ý�:����=%�=M�5>55&>��5>wyǻqO�."<�[S�^
��T������ѽ׸���D>^j���7��:��������(}��;�<���>��>Ȃ>�� �SV�<Ę�]}��k��=��">P)���=8վF�Y�=Rk��1>f�쨅�v|���d��hZ�^%���-��q�0S���ë�=O��>��	?�c?ʟP?�1?A
?mL�sP�>�D>d�>��>@�>�υ>ɚg�ʎ ���;u�Q�o�p�n�%�LӒ���˼l��px�;��">o�+>�k�<?;�ٽ<�Ɋ=+����s��]mJ=�m�=CE�<�L=)��=���=�7�>�E����ƾ��ξ�D���)��&��\,?��=>��>�e��
ؾ]׾�1P���n��x�>h��>�A�>��>�}>>+>=3sK�8��=wI;=�)����=��=�'����=u:��y� �ͽ�$������8�=(��=��>�$�<�ߦ>
y:?�
?N{=?�a�=�qD�w�
�1�/�.���"���
�>�+�>>�}>?�v�s�񾤘<��Kݾ:����@�o���=�>NKl��,x�[��=!;>�@���P �<�ב���� d�=��>�L�>�_�>R�R�q��F��� >��7п�c�����+�վ�I<J�.>��9���,�Ƶ��`����R���<.Ӡ�`�5>��2>4F�=�7�]�����S!`���+=���C��vՊ��Q���e�>��=x7��Z�������/���t��fX�rc�bv �Z���� h>?V�>��>_6?m�>+?��+���>���=���=[�>���>��>�h�>;��=~](�Ϛc�����k�lS��Q6>���>�s=�L>��=����rt�=L? >J�H>y��=���`�:�7���ir�=��>�l�=TA>��>Ѫþ�l��D���2�]M���F��4?���t�Ҿ����7�����"��=�Ӎ>�u�=�w�=" �<���>�(�>�J:>��1<��.�5/����=���<u�a�����=���<������>:��a�̽�������T�=Ms�=�J!>ÕA?��>W�?@��b��7�W��y�=��=�����n��*�����y3�!0�	��Z�<�>z;- ~�M�X>�$<Nt����=V52�AV��j^>OqL>�����7<�V:=�E�>�e>K�>��A=}�����EY���|��z����ʿ���C���r���e�����枷�����(�h�a��b���V2>�iZ>,>^�=>���=+T><�2T�P���8�� q�����i��������H�>���=�tN���ξ���5x1�7��|ك�N;C�7kC�����&{��J"'>>�G?���>�&$?�0�> �?)!0�*@�>y��>{N�>0��>C/�>�w>,�<>�K]>X�=�|;=.���Չ��O8��\PS>3��=��=lo�=m�=�D⽤ýU�
=~��=k]�=��ӽrV�17��L��=�>ԇ�=%�O>���>-���n�Gg�2����Q������m�>�Ŏ�l;2=t���1�󾫽վ*���&<�KM>/�>	,�>�f�>��>x�<�צ=9P�<�"�F�n��ah<f�e��;�<�G>\J�=Ә=��b=��;�Y���B=60�=��">�N>��s>�#?�?>�?Y�f��͎�q��3s�-ܲ�l>���>�$���j=Q�ܾh����)��ݫ�O���^!x�����͔=��>� ����<�%�=Ǟս�SN=sT�=T�{� �#�&!�=Tq>�6>wӂ>�k>=|��"�ɽ�NE�ٖ�e��i�������>�0Q=��[>�{��2�9�b��^ʾ}:ܽ�x`�x�\>to>ߓ�=	�;��=��� z����>oE�5)=C������HB��=>�䃾j#���}��K��%���,��cl�v��3ډ����G��Oh�����>��> ��>|�J?%x�>J�?�ș�O��>�����O�>k�-?}��>9ξ>0��=D�w>w���p��gEQ�_�D��W6�E0�<��=��>�>�=�����6�<�r�<Z���q�P�����	���<�=B�=@�=t$?9X��$%��`�Xͧ�T(.>��(��n
?y�����\�Z^��*ᦾr��8���+�N=-5P>�G�>)�=���>)")>��>�>l�X��n)>T�_��*2=��5<����w��<[��� :����6qܽ~�=$1G>�u<H�>���<�2�>�0?��:?��!?vw��u�%��Q2�n>齁������=�?�&>	�>XG��{��F�,�%��v���'�7$�< �> ̅�(�R��}�=�i��=�:�='�=���=�B�A�>�"�>�0�>"	�=�6=\�(���_����Jӿ(��-��lUŽ��M>���=����4����>��=&�+�(��SJ	>8��>K��>�ϴ=^��=?K>�i>�T��E$x< ɾ�V��00���∾��s��A9>����B=����#���bT�� 㼤腽x�7�{����9����A�|>�g	?@� ?{h�=�^�>6�*>� ?+@d���?Kű=�ܡ�S$�>f�z>G�=��=�Z�>��=sٲ�?ҥ���A��1��L.o>Ƀ�>U�;mu>�F2=�ks�:��<{};>X8y>5_=�������g,��7����7>��=ǔ$>t$?9X��$%��`�Xͧ�T(.>��(��n
?y�����\�Z^��*ᦾr��8���+�N=-5P>�G�>)�=���>)")>��>�>l�X��n)>T�_��*2=��5<����w��<[��� :����6qܽ~�=$1G>�u<H�>���<�2�>�0?��:?��!?vw��u�%��Q2�n>齁������=�?�&>	�>XG��{��F�,�%��v���'�7$�< �> ̅�(�R��}�=�i��=�:�='�=���=�B�A�>�"�>�0�>"	�=�6=\�(���_����Jӿ(��-��lUŽ��M>���=����4����>��=&�+�(��SJ	>8��>K��>�ϴ=^��=?K>�i>�T��E$x< ɾ�V��00���∾��s��A9>����B=����#���bT�� 㼤腽x�7�{����9����A�|>�g	?@� ?{h�=�^�>6�*>� ?+@d���?Kű=�ܡ�S$�>f�z>G�=��=�Z�>��=sٲ�?ҥ���A��1��L.o>Ƀ�>U�;mu>�F2=�ks�:��<{};>X8y>5_=�������g,��7����7>��=ǔ$>t$?9X��$%��`�Xͧ�T(.>��(��n
?y�����\�Z^��*ᦾr��8���+�N=-5P>�G�>)�=���>)")>��>�>l�X��n)>T�_��*2=��5<����w��<[��� :����6qܽ~�=$1G>�u<H�>���<�2�>�0?��:?��!?vw��u�%��Q2�n>齁������=�?�&>	�>XG��{��F�,�%��v���'�7$�< �> ̅�(�R��}�=�i��=�:�='�=���=�B�A�>�"�>�0�>"	�=�6=\�(���_����Jӿ(��-��lUŽ��M>���=����4����>��=&�+�(��SJ	>8��>K��>�ϴ=^��=?K>�i>�T��E$x< ɾ�V��00���∾��s��A9>����B=����#���bT�� 㼤腽x�7�{����9����A�|>�g	?@� ?{h�=�^�>6�*>� ?+@d���?Kű=�ܡ�S$�>f�z>G�=��=�Z�>��=sٲ�?ҥ���A��1��L.o>Ƀ�>U�;mu>�F2=�ks�:��<{};>X8y>5_=�������g,��7����7>��=ǔ$>P��>�+>!�M�|Y��oL���F�F�?�0?z:�D�>���P����������F��=|"�>q�>���>̩>�|1>]���8�o�>=�?k>�1��[>3B��ʧ������tD��Kk�������w=i��=�>o��=�潱p�>�qO?��S?�% ?u��*S���A��1�4~�z|D�jB��5���=�������c�=�>�4�/�/�ZoW�;jɼ[އ>�t�H ���~_�[�G����=j��D"�>͢�=%�=Z�=p��>k��>��>>�e=�=����:�aM�myܿK���ݐؾ����P������o!�%��d�1�!F��<[4���H�<�4{>ܓ�>Z�>��>�>O c�`�I���3����<Ӻ}�_q��2����������j�;"���\���>�F�D���O�~R{�9���=A�t�\���Q���>���=�ߓ>/q�>�g?jV>?�:>��}>��[?�͗�h�?h"?�W+?��=?�?>��>��D>��6�x�Z�̖��栾���=��e>�R><!�=V�.=-�ӽ��&�ʋC;M��=�=��&�n��_ ���l�C��=h�7>;)P>�o?繾> ̾+�о�y:��7�;�W>�q>��¾�\�>�E�y�̾ӗ��@���$=��>Q>6��>L��> np>,�}>|w;����<�y=?��=���Ո,�2��=��ջ���=mI���G�#`;�`���_->΢�=�tg=�=ν�v�>��?H?H�??'��
�߾�#+�d�$�M������$�`��y���(Y=J{Ѿ-H��S�Dk��Q����?���#��G�j�?>.�2="2�>#� �I?�����>(����b.�>k�>�T0>^D>��{>:����B���q���&��o˿���ag�UD����ļp��iЍ��S�<�%��GQ��7�=���=�t'>H�>�B>Zj
<k�=���=��$>%M���E):�Zg�Ÿ@�yѷ��:;��q*=�I=��M�@U{�<����G�׽�+���w�C罞&B�v)=�����>� e>ϔ�>�=>��V?�Q�>�O>��>��`?Y� ��*>w��>�2?ε?פ�>�\�<!�=��\����U"'��l|�O��=�7�=���<��=:
>2m��i��=�b3>��=�EC=k�<�D���6M�#g�=�P3>-=p>H_I>��>��=T/:����g.�Se�<��>��F>�KҾ��� ���,X=�h¾d?㾕/=����=[��=���>���><�g>\�> F�v�ں�n>(�j>�U7=?�=�J�=��h���ox:��n����ܽ�ҁ��8">��>�/�>{�<CU_>�E�>��I?�
A?�u�<7�.�d���W�T���6�$ց>s�����<�m����Y(�Kw��r����)>�'<8�>U1¼��
���">�q���vC;�M>�)�=�\}���>��>т>�;l>(��>��=93�G�&�����w�ȿ=]������.ͣ�p��c��f�=v�R>Q>P���=#�����y���ҽꆑ=��>t`=�>a��Fg�~^�Gc�p`��醾|1f�
&�_O��a��x-�+�����[����"8��b��y�����Ɩ�x�R�J���V�N���>���>�7�>���=��O?s�?�!%��}T�s�(?Zc>�-�=�$.>��>��?[� ?�>y݂>����Vž}��1���?�{>�օ>�02=�,绨��
�нq�r=���>�YT>�L7>��v��
������ɽ���u�=m)>Ļ�>�>����&����=�Eýs6�>2+׾I�������j�,�����镾��s=2~>51�>��=���=���=9�'���>��>C	=�K�SMC=�J�2[c��䌽�Žr���(���U�-F�<�i�=������=׼s>Jy?��6?�FG?���М4�ʒ����徢��_H��S:>�c��C�;�7�r��C���L���Y'ɾ��P�w��V>�>�.f;Ҟ�p�'�<����K�=�)>�B;;m�>q�W>�q�=�H�>���=����$���8@Q=�Ŏ�X��Я�s��h�����>6�>t��<`��N`+<<L�=����D��!�=���>�K�>��>+u>�==��$>����B�<�=6������������o���o˽�gZ��t�=�P;���R>�<���[�⽶j�erB����J+�ѣ>_�H�q�>�m�>�&?�в>�v�>��q=��?0]�>
+�>S�?��?�?��?w=�Ži���P3�����M�x�����Fp�=ͽ�=�#>��=3љ��ɔ=$+��&"k���]=V\߽�;��q��=��=f�=�>��7��>�xB>6��о��ݶ7=���<B��>oU��Rɨ=Bg�=Rȷ�/�r�E݊�Ǚ	>vlH>n��>};�>9�L>��W>4� �מ���ײ=��=>�=#�����$>��I>)���D�=,'=<䩽1�y���=�,=$ڛ=_�-<��>-}?�!?��N?�"���>���8�'f�_p��=�:���=�ۆ��?v�cu߾�<��T=����� ��q�"�J9 =G>�R>1�=)Kr�b�@<��>���X���;�=�j�;�1>n1�>�L>NȽk2��E��w7��kؿ�K��H�۾P�#���%>��<�!%��|4� �i�� ��{�8�@(��,>W�>K�=�ψ=����"���2D���ͻ��1�p���1�ý�dŽ��m�z�N�{YҼ 
�3�Z�ֽ�'-� ͻ�q�����1�>͎>[�=�^>˛�>�)B?a�x>	�>���;�r%?vD=�S:�u
?��)?��7?�#?�bT>w����W۾�۩�^�'�;��TH$>��>$m*>�0��>�������6=�=��=ަ��V�d�UO��6�V)�<�e�=H�;>�I�=O��>~#.>��1������W���Ӿq��>��?���2�>�+��K�b����Dھ�S9�CyG���K��>R�?|C|>�o>2AP=f����f�=2��i���oD>�����?�ӋW=��>���=fsq��u������ޠ�w>Ԩ�<�Լ>�03?�I?[L?��?�y_*�L�X���=�ii��ohһvƎ>_x>�(i��￾pԾ ����#��"��Ҿ\Ek�� H>M�-�RI>�q	>�A#=���=,	�<Y�>۹��[U*�\���.��<�A�=���>�{>�W�;�3[�����~�!��9C7�x	%���l�>:��O���l�rF��9�� !Ӿt�j�+B��r>>)iG>�@�>�=��٫�=�IK��Ց��R��y�=BӾe6����ҴN�t������<��"������x��m��~�^�)�`�Gխ�{䛾p�˽[8�>`�=+��>�9>pV?W�`?�ժ> �N>��]?1f6��F<ñ�>��Z>h�?�G?Db&?��&?��H=���F�x+����<��4�<=?��==Y�3��z�=���=��==Ӎ=�e)=��/>�D�;�=!hP>��>��=�>�Y�=���I?�\�q�����l>a��>��B&>�h�������=�p�l,�B5˾?���M�,>a�>���>�FO>u/�J܅=3t�=7@x���>{�;>Ƞn�'����\<N�6>!i��:���\��k^��x��Y�>8��>��>M?B�:??-?����aUF�Ey�n1S����Vn!>���>@��>����Ĩ>�^��T�7�`(����ؾ���=�
�>��4�E�)�2�e������̽���:�B>��ؽ�D-��7�<�tj<w�>�~�>�l.��S��l�K��"�J��l����ɤ���
��=ٲ	>�Њ��B���>�<6>�������M	>"��^��>�M�>'-a>�>ǵM��M���c~������+���e�	^��摪��Be��GϾ��=❴�����N�->ڡZ�p���e<pb���ƾ�-���J�>$�>U3�>8��>�#?��>�g�>}�>R��>�	ܾz"���6>za*����>�v�>p�=TA?�@��e8a��߽�镾E^�>�&�>G�>d��>'o%<Q�{=?�f>t�>��>IV�=�軽^��<T�y>U�E>vή>3�>��7=�i⼩�j�+��"E��\O�\l��Ϟ��\�s>�u���!��P��X� ��ϰ����p�3���-ǾA��>�?V.�>��=z�X>Rs>���=3��dR�`�^=2� =���<$2��i��<�<�sG�H�E�P݇��є�=xl=?&8=��>:?8P?��i?�����P�t"D�6;)�䳾x	=%�=@^E>zÒ�,���-ξ�й�^?'�(�3��ݒ���g���B>���O�$=�Ə>��=��~=��>���>�_��}�Ee�<�{ >Þ�=�2�>m;�=xӘ=���c����鿣�՞	����f�=0&=QR�%���↾�'>�u����*��C����</^>�v，C�=!Tg=�6߽y)��sF�z�>����n ��a��@p��Q�S�{bܾ��a����6���>�Ⱦ���H���}�Y��g;c�˾�{��)�>�Y�>Є=�`�&X?��E?ӀU?��>6�?�����f�>NE�>Ay?$?�OA?�	 ?��6?0c>�,2�?=üT���ƒ�;��b��=�mA>�>�{B��X���>_1>��=`x;=���=��%��s=�k,>5�T>@�>��E���=�=��aҾh�F��F��*LU<���> �=�z$��B��st�e"��_M�q�F��FJ�"ش<� ��|�>#=�>�5�=�/>½�l_�<>	==iS>t��e��<��>AÌ=/�<�4>��?<�qi��� �מ�O�8>oK�=�`>*]�>|/'?I[w?xe8���L��sM���9�e
�� ?^�G�N>߹�<I�9��ͦ�qhG�����)��X�8����S'�=�ق>����ӟ=p;�>�� ��J=k1>�gz=�X&�S�_������6�m==2~�>�Q�=���<8,	��<��"�E�Ͽ=�����0�X��q_�;������^qr����9����<󒚽�kJ������>g�>{��>i�>+����	�a]W>ɻ߾��e�.C����}�h����1���*����������վK!����Ľ�ſ�]I��E��>.�L>>+v>�����!D?~�;?��?4�j>�jS?�?�y/�!�>���>r�#?N�1?��0?149>8��>�^�=6�ƽˏ�g��<C
�a�G���F=C(p�Q|<��'�=�`�=��>3��=�81<)і=���<�?&>��^=3?�=/�=�3Q��6��0%��m�-qc�o������	�>�����\�/�O�����1���*���uĽRլ>��?�ʂ>�#k>��#>)�Q�ɓ����h�=�C4>݆�=eZ>f�C=�2���_��R�7�����q:O<��a>��\>C�>'m?��?J�[?%<-�2�f�N�ao��3Ƚ-��ͫ>�(>I)��)�~�񮄾���]����#��o��BP-;��|>�c�I~�)��>�=�(��ҩ�9_�>�����
;R��=@Z>���=z�>�CF>z˽�s������׿����k޾�{����=��=>�:<�p������
E>x�{��Y`��L=�[>�t�=\�=w>�>��=v-�=�>���p��k���')>U�ܾ	��Rf��g��
�����c��6�
o��wWa������׾"A��@��|޾�Y�>��y>27�>��;��7?5gQ?��9?G˻>��?hC2>�>4R�>!�E?ݰ?}QI?�G?m$�> �K>m�S���S������<����'��tI�=G�(>`B=t��5l�=ݕS=���=Z�=D>
t��#W?>D�U>�]�=���<��>�m����"���]J'��P���>9�>�������>?þ�_X�̷��_Mξ֚�����rR��>�0X>4?N>js=��>�f6��F�=�bh> K�I����X�=S�=����Y���9�)ߕ��h6�Z�n�~��=�f�>$r�=:A?4�U?�
,?�^���8美%*���8����)T�~�/�C�����w��i���^�ݾg(�e�I�ԑH�.;>�B ��U=`��=�A��,�<�6>�G�>}�>���>+l�=:;�>�ň>���>�u�>�Z�=9�N�ib����ӿH��� ���`9������ϒ<a��>�2O��X	��콼��>X�6�φ�>}+$>V-�=�F���>��*>�����'�2��Uo�=��Ǿa�������5%>�FD�;^�sn �P�>>H���医���Jad�x�F��!��>��>P��>�`J>>P?��3?���>�A�<iP?��=D�>z<	��4? n<?K�?��9?��J?K�>0�$�O���#�+�C>�/=��<�
W>X�>�tD�yƎ��4����=>��=.�)=�!=�����'��=Y)>C�
>�F"?}�D>�"�����D0��bz��/���&?8�1�G>��"��֢���.�Q�-����0�
�irξ�]>92>S>q<>�Q>[	��O��={&
>W�½6좽�=�uҽ;e�kn�}�`�*�'�)�|�j�`��ƭ=H��=�L%>��]>�f?�l?��L?�����2�ʍ,�#�d�������	�*[p>�[\�v*$>w��r���������-�Mj�����=<s�=cd>�Ǌ=j�-��Oz�ð=4&�>4}x>n��>C��>f`�>GĮ>�o?�=�>UMJ><��L��n�ֿ�+��D��H�*���ý�ν�m���=����E>)e�B#P�ךϽȠ�>�0K>^w�=���<�Au=m�>��/� ���s�B�d=���7W��n~����=�]��G�=� ]�+�9�y����=��������� ~�l__��p��ן>��8>��>'+�>m�;?-??��?;�i�Q?��=�W?W˾>�!?1-?�~?|C?q�,?ly=>��I�������L�N���*���b���+�>�ۏ>�r�*|���-�b({�c;����Z=�V�=$能�����Z�[�>o/�=�?��=�I!�R��}���~о(l���I�>�(Ⱦ��>�)���<�����}(��C߾N������T�=�r>2J�=�*O>��=W�u��2>	�>K3s����l�=�qݼ�uѽ�5�����[֐��j�������=p4�=�hJ>�fx>��d?j��?��3?ͺ$�^*ԾK4(�Ϧ�������V{�=_E�I�ȾD�׾O���Z"�/�F���G��䃾�<��N��=o\ż�D>L�>5�\�b{g��e�>ֱ`>bʂ>�;�>!�q>�8>���>\Z?�i�>6ַ=1{F��
��Jѿ�調E$����p��a���n�=��t>�O�~Ɯ��2m�-�K>YՇ�tKS>�#>_����=n��<�d">Cl"=�h�z�m�����͠��B��d��G�=�;��Ƙ���;��=br���#�����R�vڽ[��«���ɠ>��>瞝>���>�L?�c ?��?��,��jE?�M�>�!?��T>��3?��-?��?�q1?G�/?���>���U�O�M����=ʹ�=R���g�&>LY�>@�+�k+���ؽ��r=�L�:���=��6;^t��z�"�l`ٽ�!=��=z�?q�=�"����	(�\�����/��>tZ	��h�>hg¾_��=�h�/��ɾ�+�M[⾯�?���=�u>N�A>�ɼ�劾�>���=�����=���>=�l�Ο��3�v%�;F�Y�,>�Qx=F.�<�'�=n,t>-̑>%]X?�V}?�1D?j\*���	����}�!����N�E�������4��n���޾��2�L(������&d�'@�=ٱ�=��>Q�!=�_E��̽��y=w���\��>yR�>]	�>x�>Ϳ{>My�>6/�>
>OX���쥾��ܿ�͵�����
���R��ty�EZ�=��{��
�<���=k��(��=߶�=^w,>�ܾ=-���z�O>/�W>� R>�=�I=^�{��s=����񌻾��'�~�>=���0u(���աb=n�G��h�����Q���G���#�N[ý�!�>a��>�c�>��d>�@?-�:?�K�>%$�>kmB?lɾxt�>Rg>�?�)?�!?m,$?�9?%@�>��>�Ic�ƍ��=">eoY<mw�3�>�/�>Yy,����:�:�����k�0�x���>���r�(��z��<g�<��>�m����"���]J'��P���>9�>�������>?þ�_X�̷��_Mξ֚�����rR��>�0X>4?N>js=��>�f6��F�=�bh> K�I����X�=S�=����Y���9�)ߕ��h6�Z�n�~��=�f�>$r�=:A?4�U?�
,?�^���8美%*���8����)T�~�/�C�����w��i���^�ݾg(�e�I�ԑH�.;>�B ��U=`��=�A��,�<�6>�G�>}�>���>+l�=:;�>�ň>���>�u�>�Z�=9�N�ib����ӿH��� ���`9������ϒ<a��>�2O��X	��콼��>X�6�φ�>}+$>V-�=�F���>��*>�����'�2��Uo�=��Ǿa�������5%>�FD�;^�sn �P�>>H���医���Jad�x�F��!��>��>P��>�`J>>P?��3?���>�A�<iP?��=D�>z<	��4? n<?K�?��9?��J?K�>0�$�O���#�+�C>�/=��<�
W>X�>�tD�yƎ��4����=>��=.�)=�!=�����'��=Y)>C�
>�B?.l���t�����~j��)��x$�>>�'?k5G��[�>�����P��{YP�@�K�o{���T>�;?�}?�4?в�>��l>�>;v�d���=Ǭ�=䔖����=B"�P��=cH���Ͻ����x�������ތ���6<���<�O��Dd�>�30?��?GOw>��E��̾x(u�_���Y�0"���\E�}ө��Q<e��CV��+B�zn&����n�`���:&�>R�=X��=�����9���W�ګE=Q!>a���t">&�>�&�>.��>�>��=ҡ��η����X�翦�¿�A��
�D��Lؽ�ɽN1><�,�%$��5ľټ��-���7J(=q�>NM�>J�j>3�=s��==>w@�����[h�.�.�?��9��5���I�F��A���c"���ҽ�b���S�(��ƾ�� ��׸����/�J>Q?�>l��>�?#?VT>?�E�>��>-r��05?��e>@7?�;�>�C?�D?4��>�";>U��T�	�7���>l��F��ղ=VS=���=���=��>��4���>�l�=B�׼�P��Wtg��"�<�1��+��-�=u�=���=m��>V���I?;���SH�X�& �>�x�>��ʂF>��ߐ��0�/��G����B��>|`�>���>Ih�>^��>&�=�Ĳ�\�D=�ɳ=��>Fy���#潖�!�C�=�-�2����IJ��(r0�Zl-���������K�)>V�>�� ?���>�?@A���a��K<��$ɽL��
���鼁�z�&a�91d���ﾄd��S<���"����3�!��]n>f�<>�W4����< �;6F�=X�+>w)>E��V>`��=�>���>nܐ>�%�=��=Rk)�����e]�ߝ���޾��/��Uӽ4����+D>и!������������X�<�Z�>�]�>J��=&��<،=>�l>�t���b��h6��9�}��.'�9U���+�<�X>*�ɾ��A������!ӽ�iT�悇������h�0��5'�xgv�]�>N �>�?���>��6?ab�>��g=W���=b)??b��M��>�p�>��?}?��>�[�=U�V>b�\�^���F�9W�m�>Mj�=�3S>w��=�C>,��vP>�)3�w=�7<l���+�<��f� �<��u=�yj>g->m��>V���I?;���SH�X�& �>�x�>��ʂF>��ߐ��0�/��G����B��>|`�>���>Ih�>^��>&�=�Ĳ�\�D=�ɳ=��>Fy���#潖�!�C�=�-�2����IJ��(r0�Zl-���������K�)>V�>�� ?���>�?@A���a��K<��$ɽL��
���鼁�z�&a�91d���ﾄd��S<���"����3�!��]n>f�<>�W4����< �;6F�=X�+>w)>E��V>`��=�>���>nܐ>�%�=��=Rk)�����e]�ߝ���޾��/��Uӽ4����+D>и!������������X�<�Z�>�]�>J��=&��<،=>�l>�t���b��h6��9�}��.'�9U���+�<�X>*�ɾ��A������!ӽ�iT�悇������h�0��5'�xgv�]�>N �>�?���>��6?ab�>��g=W���=b)??b��M��>�p�>��?}?��>�[�=U�V>b�\�^���F�9W�m�>Mj�=�3S>w��=�C>,��vP>�)3�w=�7<l���+�<��f� �<��u=�yj>g->��?��սѷZ���:���K�U�U�P%�>:m�>Q(�fs?��f��D�C���E�k�6���>P?;�?��>>-�>O�
>�ͼ���=��=��+>��X�9>n�W���O���g=�h4��t�=�������o�.��Ij���ý��^���>%T:?�^$?i�?{�p��m��n�H�Q`�"�����r[]��B��h">(迾������7��r�}�"�̻s�(��]�E>5��C�=�m��=�w�O]N��g���]�=E�?�j8�;�z>�܍>�>��>IՏ=��<ʽO6}�%��2���ž	� ��}����V��=w�r>'ɹ�!wI�����r^==��ռ;�Z>GO�>��;>}F�=�x>�>�m>���转��߀��ɾ�t���D"��軽!s���>�\��u�
��k9���0�����a� �4�ݽ����`<�9>�֦>B3�>���>��,?F��>��P>P�Ͼ��F?���o�?X�>t��>Nx<?��??�=
�������޾�����1��$>��=���=[}�=|�x>[2��n#>��="��=�@��Y�ǽ�
ầ4�<��G=�b�=66>��	>��>���;&E�����$�,�1S��I6�>��?����Oɻ>E̾W��G���: ߾�^Z�q�w>f{>B�>��D>.�>D�=�Q����Q�e�=i>��=|��=iU�rX�<��2�D߽��Խ���9߲�iW=�v�=ll�;�/=��<�??��D?%|a�t�X�3���!���&����2 >1)`�c=����ž�s�X ��'�,��PR�s;�=)&�>_�><$p������:���}`c=L�>j� =>>�>_3>��+>`�>c��=�|���A���s���&���Z���,�a�u�X�7�,!��T�=_�H�B���>�2�l1��?�ٽ%�2�8->��^=���=�/�lN5��2��nξ5[��W�B�7�;���s����k�<h�ƾ��1��C�5׺������+��_c�������=�7�=U"�=]� ?�'�>�}\�֘??�9�>[�۽ ��0z$?G��9ڇ>2��>R�?��"?�>��2>��{>�i>z�8�r���K��?>WE>�CU>+�<�A>��	���>a0 =��>�.l�����/C=���ln��40=��j>� >�?���ҫ��������o�
��	_��?�X1<5�b�W�ǽH�ѽB����o��V��q���*�޾� >�_�=��>���=�f�����p>�S"=�#�J�=�v�>��=���=:�>�ؽQ��Ǽҽ�DU=�,<�D��>O{�>shf>Vp?��?�~*?���>쾝���ھ��/��fQ8>�QJ=�0=n�m��^����Խ���>�W�7Y���K?=�>� �=-9�;�ee=ď�=�g�d)�=�L<�E��*#M�*�>e�">��R>�{-=��$>=J޽o����cԿ����j<������|:WJ����>�JT�Ih��hY�>��ڽRA��{�<����F6d>x��8<B?���>4�,>"�;��`��N�+�5i�<s����Ⱦ�ƚ� �->�����H �=�7�{�zo���W�����z�$�x0���@�ɖ��>�� ?�:6>��-��Vl?6=?��>�p�?��ݽ�T���!=>'�>7/�>[w�>@��>�q>�$F<�D�<+�D�����|1>����I: >�A>�TP>��O�ʭ����=`󥼹r$��Z@���Ž�����y�<0�J> ;���z>��>d�/���Z���?0��9Ѿ�|����2?#�Ҿf�n�?�V=�Ar�3���vs�������l#��+��>��l>1��>⹴������O"��~=6��=�~�;,�-�+O�=�}�=?�&�g�=1e��u�#��E�����]H��;>š�=�,>�x?}�?�0?�2���@ݾ'R
���-�бp=a_=sA>��<.jW��^���1ڽ׌�}�_U���"A� 3>��=�O>;׼	>��=�;>�>-��Gn��-��;m#�>5Y>υ�>�.>���;�C�������ݿV.��C�̾_�����<HF�U���/5p�%nh��=�������̱�=Z������=$_>&=�>�n<>NX=^�B<bK>Ը����!7ݾ����ξ�D>O=�������G�D���/&�2���!�˽l�O<�������a%�p�#>	/�>T�c>���_?��=?m�?W?<?�>��>��B��P>{��>n�>v��>Po�>���>x�=so���Q���N��H��::���D>f@8=Y��=�8�|�½U'S>���=�F/��h<�;|�߼�þ�9�>��:>�IF>�Y? ���/��JQ����3P��BF|�0Ě>2!ɽ#�=��Y>�+>�1��b/5�؉]�v�2���ܾ�/!=��+>��J>hi��ƽ��޼�������<�	>��Y����=�fὈ�!�O./���k��.��_R��믽>�ѼOV=;5>7�>R�?�>��4?N���<쾨��+� ���������W5>�0��A;��-t�vٳ��s����ƾ{�%�uQX��n`=��=���=�.�=��;1�=g��=y�=�V�5ż�E�=���>�q^>^�o>'��=����ں;vU]�{��A使۩�Pr��zͫ�1�y=Ƣ�<�>=�(�<Q�D�RW���V��B����U=ũ�>�\m>F2&>�|�>�N�<L�>DH�>k_��/=�����+ξ�f�ֽ��_Y��q]���3<�����9�*�=�zo�]<ν#b��6m��wL�&M>���>�mk>ٚ2�h�u?!>? ?��=9�>;bY>�A���c�=f��>Qs�>$��> ��>K=#??_1:�k��g���愾8��=�m�4.>�l>><X�=�Y�ǝh��p�>�T�<w�p�럽$=v>�C=��>V̒=>�>H�!?�fq�
þ'�Ѿ�$�F�Q��b*��ܒ>�bq��G�Ⱃ>�/X=��T��e2� 8 ��8;�־	�>�Q�>]%S> Î=w;4V���䮽X->O�#>��P��~�<,%=���H����f� 4-�z'���B���;k�X=�>��8>�c?�j>%�*?�����W �D����9��bt���C?=�D�~Qҽb���%����5�ܾ���2��»Ck>�[=Ǧ2>��>^� =�d�=lW=I#�=���=~��<Î�>`Vr==��=&�=5�9=b��j*���忆��,�پ*��,]�L��n^%�*��>�GG=X���o���}��gY��T�>��>��>U�=B=A>�v�!'��l��f�	XV;�@�4�����+S=[����ə�x���*����)�y���8�\�U��+�A!���$��(�n�_�>��>|�=�Ki?H*5?Ҁ?��Y�>�>wj���߆>��>�
>��>/��>��D?��-�� =�+����l��=Rν��Y>�:;��=�M!>�T�=���=H�>p�]=�Ju=u�<�)�=��u=�xf>�H>�5>6(�>X�s��c�Y�g����E����+`�O��>T]�������>�I̼���Z�ʾ�c���n���߾4>�^�>��/>���<ʆ=T�4�b�=����==�m~=���=��=��=��=�~u��f<pm���=�v�<S�=�>���=UF�>}N�>�A@?�\����*��X�ά��'��>����+>f���R�������p�q�u%��)�g��1�U��j�=l"ȼ��=�SE>�=��=nS�����S��<Ԕ=\�>��S=��=r�v='��<�>%���Q�o��8u��	���+��%�ἡ���(�>+_>����Q.��&�2h[��(ܽ�ON>�y�>��>RC�=�>a֬=�C�>�R�>TM�dr����W�پ�o��>.;���2����z��U,�'����*E<,ة��G߾s�U�o؍�\ؠ>��?֐��):�wZ@?<-?���>'<����>��.>/a�~�>�7�>�o�><c�>�#�>�?@��P�z�b駾�C\�,��_=iO�=>��=z�l>)��_t�#y">.��<x�����<�h＜(�<#�Q��2=>C\>�!>`<�>��A>��J���`�b�̳�=����$;?Fҽp����~ƾ^���M�����c~��B�>@�H>����ꕾ�/>� I�y4�={Ԝ>�g�="���Hr�=a�+>p7��r��<�y�����1���ϼh���!=�@���%�>y�? �2?"sM?-��>A��>�2�'�
��ZѾ����>x4��i�6>˯�>!�C�004�~��u�&���9y̽�9u>ڟ�����F���S�=	��^?���h>ϟ�=�X�=��
>��><��=�z�;�n\>�>��:;�`=:����������]���8���;>)1>Ƶ���I>q=l}���ֽjo�2A�zr�=N��=n���"�>n��>?��<�]!>~sν�X�����&�zj����6���x�=�l���c���m���*��YT��k}��
�ҧX���ξB�<>��˼�e�>��F��I�>�L�>F?H��6;�>,w�>x�>��?X-%>�^c>���>S�x>"Π>�9�>��f>��Ž�d���sȺro�*��=�$/>B�>N�=[��V)�%��<I�i=tӻ�҉=�Z>�[��i�<�6=�S>���>(	@>��E��þ��g�2ہ=�=���>W��=^��=��R=G����A����i���ѻ�};>��9da�6��Nv>� � S�=7��>	B=x\^<�n"�)3[�;i���SK�����hV�Hؓ��>���T��3��*��fF��|�>c�+?p�R?�f?ъ�>]TV���P��3����꾳����e�<	�>g�?b\�>Uj�������;�*�X�,��d����q>�
)={��=
}~>,���Dl�l�.�>-������=	>��=��Z�K�H��9�=9��>p�F�\�}L�m�Ŀ}yؾ��u��;��X>��=(C���L������Xvt��k��zc�B;�����t�>bl�>�G?�q?D�N��,="�,��@d���¾];�@u��FŜ<ގ<�x�<*�+�S��n��	Ą���[�;M�d��n^���T�r��>���=�a�>����?d��>�(?�������>�>�.[=��6>-AѼY87=���>�5=��r>��c>\�y>s�F�E�T�R$<��A����75`=.>*�y=<��<���=���=�#�=��=�ߎ=�|>��<;����>��g>��>�]>S�7���پ$=�����{�,I�>d��=�Y�>�þd3���ؾ����;S�e�>e��=Q:���~�ϗa>N�c=.����E�>��@=�����z$>���=��׽VjM�j�/�"�2ZF���	��ά=X�=Y�f�xn���.W���>Ho?�UQ?��H?��W=�I=�H��ɫ������ӻ���)�>9��=�>�Q(>E/K>�\�o+�����,��Ҏ���L>��=vu�?.=^
>)���g�J�x�4>�����>ށ=[]V��=>���jˎ=W�=KW�>��������ƿ�$�.=%�~��=�Q�>�Z>�T!�&8=pA�<���%%*>�N�m��~�	w�>%�>S)?b�>�tr����<E�8�94��������d����;��r=��)>�^+�d���;E��P�����9�}��F�v��.V���>l"�=g�>79	=��?��?-F?����o�>j�a<�d��Ha�>$�a<.m|>���==����>
z�=K ~>嶹�����b*=�"��f�=�:>tjI=*6�=�E��{�="Z]��bN>U�>*������=��aCo>�\#>�{>H�?���>�x�����_�=�ڙ>R3i�^d�>�g�>�Zh�((þdm�����RM���澴ᔽ�~7�}j������iE>0�z="�x>��=l��;]+�<ih�=?� >[L���1�#����p�1Nk<G >�'���`��d��>BH���0�-��>�?KL?��H?�/>��:��+�{�˾{۹���ľ�D�>m��>��>ΉF=AJ�=T���a�]��P'�Ð��QW>jJ7=RS�<�*>v����0�<NW���=�H���>u*l>�1=s/@=% >��޼��F=�Q>o$=8tο�����8��#߾����ٱ<�ʸ>^3F>��ɾUb�>ї?��-=|
�}W�=���>��>8s�>d?-��>yL��XF<��x��������"�t9��I���t�~�Xݖ=q �m��6��>K��z��f�i���L/D�sQ���>7�>27�>�e�=��!?��>�?�难���>�/q>��>�<>��==�&>��H�߼�ަ>��d>�>��������K7����Ӽ���=�&�=ǡ$>��5=O�p��Y�<H�=>>
g\;/��~��=���>u�\=C� >�O
?��>2�8��V+���Y����>m d���>��=��a<@+��0^�D$ݾ�����3�҈��F/=Q��E0���S>X|#��@�¸)>�=����vp>��=��^��jԽ��ͽ��4=�ǈ���&����5Dk���O�j*�z]ɽ��>��?��\?[W?���>��5�$�#�B�
�/��i��o�?}ȸ>dt?s�]=��=!P!�������eK��[����4>9�0>
鵽Ō�=�p�=E��<-F���=~f^>:2P>Y>w'I=9l>=q>qɟ<%,B>Q��=	��*#Կٹ������߾�H�_`;
�>x��=��
>yb'��|޾�!�=�y�i�=�b�#�6>"�t>D.�>��>�����<C�ݽ�&������L��<���q�����@�˼z����c��=*
�14��v������WҼ2�>��\�>��O>B�>M)�>&�5?�� ?ZQ.?U�<��>K�>VQ>�a>�$>L�#=�)w>���>_�>���>?��=�Q����T��;M�@��;G߷=y��=ί��:>�5�>�[��#��<�=k���=���=��}��f�='T�>ע?����y\���,���,�9b>�<�<��?*rJ���u�GM=񋁾|�>��<5㍾�����{�T��P׽d��>��M�	��=���@|�=��)m>>�O>�_�<�c>�QX�;�!>�B> D����Ҿ��<�sн}d�>�>�g>�j�>/�E?@[?|�R�5�*�Z}��l��^F'��N����>�jG>��꟔=5)���ݾ>�����<��M�������a>�"�<�L>�:>�Q�=Ԫ��x�<��>��@R=v���}b��Ȓ>�~�> ׽*�I=�K���O�޿�뤿="e�Xlپ��-W�=-9�=�;����>��'=�Da��Y�Zl=Xt>B^�>hn>'?>28?�2��r���ٽ�ŽV��R�0�A*��?������Z���>J���%���+��u�J���,�AX׾�斾���R�;�.�>��2>��;�2?��>.�>�ӱ��p�>�>���İ�=�Z�=�1y��+�>�I�>2�?V�`>�/G>	Q�\���-<?�{��#_=���=O��={!��
�وD�l)A>���<����;��;�I9>��>��>��)=Ai��+?��E=�e���*�w����P0>�?�A5��}�i���l��1�>&/�������4>O�#�3/�=QH��s��>��߼:������@��=�fH��r�=iE�=s.Q���L>������S=�w<�>��\�m�g��G� ���]>��o>�=�?�(?��2?to�}s��@���,�y��a��݂>I�A>�x��@�]G���#���	������K=��i�γ>�3s<]�>m>���e���x�</x�=�Q���>�i���"d(>�=M>�E>�iV>n*���6�mֿ�Р�8vy���޾�͓�ى�=S�=�z��(��*�E����Խ�>?��b�>��~>,�=꒠=�(`�����B�\=.�&>�K�S����(��B�ƾ��h��K���֮�ԪV�T�<,(�5�����:���ľ�M�?��\;�2 �>��>�ph=SN5?f,?rs?�`����?�qj>C�l�oR>�><�=�'?��>��?n�I>���>�:��4[�_J�=�/�=HG@=$�>[�>����h���><M����i=��
>->=R�=d��V/z=!&L�\�=�?�����n;���#���5�I�ɻ~�i=L��>��l��T?��eO�3�l� =8P��b�^�����/�3��$�����|�>��k��R�=��1�N�<��o�B��=��Z>]�佽aS>))�=
G�;��=
"�馄���(�y���jl>��e>��}>4��>��)?[^Y?8=׽�?��kC���=X�����>&C�>ȼ�=7���
z��F��'�)�x�׼O�,�=.�!���w>�J�mH2>4J�>�n	=�!��m����=I�D���-׸�U׽��=��{>�=>�Cp>�/.��k�b%鿄����wY�O�ﾡ]c��L�<�Y�=�`��n�+�0� M���<�u[>� ?�:�>zZ=�qn��(l��欽ꍔ��b���g׼|����,�CS�����肐��������=�'���tӽ�`W�ʜ��V���Q��JXh��۲�F�G���񽇴�>��>��=�S?Z?B�?�K޾[ȷ> >��|=O�>e��=�ך>s?��?>"?���>�n=�ڽ|u&���[=��<�H��9>$��=у�;�^+>^V��ux<N��=>��>��l=0򤽔RJ�g�A=��>�h���;�C��V#��=>t�Z>�Y><���9<���׽�ߥ��'�p,��dw���>���=��=�q�پ>0f
���>9"`>�����⽴�f>�9+>[߶=cW�>~>�=绨=�0�����`B���	^>��>�@u>�O$>u�%>��>q�&?;?����(*�����Ϧ=�ط=�f�;�-�>7�a><s���BW���������K�t���>�7���=�W�5KL���w>��+=^rP���:�f�>���-h�q�ֽ�>=ڻ�3M$>��<M�=`�����G��ο/���#����� �? ����9��I�=����Rh��ij^�����V���Ñ=�o�>�?��꽍P���r	��!�;M�/>���>vJ��q)��<��&L0�G�����.|~�Π��Ym��EFR�?���<��M������㬾�����ľ/��ɷ�>��|> =��<?"��>��>px��8�>@/=8,���o>��%>h
O>{?�j�>Jp�>�7>��)���k�������=j{������X=r>�������v���p�=��=2�>�P>C�*>����2����
�,>���>�L���oE��f��z� �(
�Ba�>gyg����=��������ͳ>'"��Ot����C>��=��=������K>���;�f��]>�
7>3_=��1>���=Ox�m,������~�K	N���r������=?ټ�#�9=?�=j��>�B�>5�?ݜ?]6�`����͔I�6 ���#��Y��>%qr>?o����=�wǾ���8�l����f3>�h�Lً>�k
=��5�/!A>��f=�����`k=�L�<F���I�=���v!�=8��=)��=�̓���q=�\�W��ݿʮ����𦾛�mmZ=�q�=�|���U�BϽ���C���ܽt�>"@b>��>9�3��?���*�U�=���=��f��2-��&.�V݂�Kj���z��#���u���� ���U�;���<��ϽTꕽ��O�]^u�^�V�2����:�>�>�8�>��?���>���>�෾."�>�S�P�����d��OF>wa�>�H>���>�2h>MN�܈�b$��2	h=N��=�*����I<H�=�H$����=U�=��`=5ɵ=mR��,�=�Ć>RǄ��nF=@�=���=��?���:�"���<�H!*�̡C=���=O�>���=!�N�vz_��2�g�����#�U>�h>}E�>L�=���>ޑ ���[�#�;B��׾�<���� OY>C<c��8���1>OI={w���½�K���T��l2>V:;<�V<��L>b�+?�(*?�j?�w�=�/����M�[M佗�$�FEO=��>TQ�>��>C�D��N	��)�c�8�1�&��`�����"�>y�[>��>g-=>Ԑ�=~6��f��}�+=�|�;'%����=?R>m�=�^>��==�-������՞�����R��􊟾{�3�3��h��f�߆����=�	�<PJ����B����=b:�>w��>�P�>���=�A�<�_z>��g�?��</���C��,s��{�˾��4|�'k|�Q�P���j�+�#���#���>����-�d�%�W�̽���<2˥>x��>a�>E�9?0Z?�Y�>K�>��q>+����>pk�==�=�9y>�_>���=~S>@&�=%S;��̽3
��>�.=��<&7>'��=H��=�6ʽd� >�T�=shQ�ߵ�W��=X��=��:�=L~�����=y>�@ ?Pt��%[2����,yL��%��C}%�tg<��<�=��]H��y�f�l�޾lį�a(��+=�\L=R��=Zi>%��>A�g=����Ί�~�1��E�=�
>��h>�XB�I	��Ȧ>��u��H��@���2������=Z�G=�{>��'>8�w>�"?�?�L�>�G>�e�L�vA���Ⱦ�4�=��>�K�>��>,�N�R��
,�L%�w�ᾑ ��k�d��$#>��>�v_>��)>'�q=������ýJr�ߛ�x3����<>��>S/�>���>B��=��(�#(���ѽ����������9X�������>H+��I���E�>�~�<��˾%}�=U5">�S>H^>յ2<���/~�1Ŭ=��Q�^c���\6�ǩ>��T�ݾ�.˾����5�)(=�徺�˽�N��X��I�6-4���a�yM�Y�k���^����>��>��W>>?���>[�>��i>$w�<t����Ύ>�ﭽ��=1kh><]�>�{�> ��>A�Y>�RC�R!�G����Ѿ=8�p<C�=���<3Pm=��
=���>�2Z;�8�B)�=�&���r�������ʽap=�(b�×���>^r������7徆��U��=ד
�MdT>���=�]�>&����&��Z����;�===kV>�� >-�>j�>1g�>���=�|_������=l���7>TZ>�3��έ���ѽe}&>J�>�ǋ���#��!�^��b�=ۦC>~gw>3c.?`��>�#�>�E>��%��;�J����R�I��^>ʛ�>��>)Ej���^�������t澇����>\\�=��>��>L��=�i-������g��o�r�:��|��s6=���=�9�>F >7ك<���o��#q�I��� "�;ə��K���׍>�6[��-��EVA>���=�����;h��X(>�k�=L=Gf����*��3���,
?�7�=�R�=���%.�6��<j�+�S�4���_<�8�X�<�����~�m�^�`!�k�m�\(������~5�xg�>��>�ڦ>4�-?�5@>��>��=��&>6���_�>�;I>[OX>���=S>˰6>LZY>��=��P�n�l�p���=�R�<	(���h$>1h�=&�;�<> E>f�#>�e��$K���׃=�/=��>���=p��<Y�=���>n�Ծ��ܾ
3/��
L�W����2�=��>7�>�9`>s�
�32��xl�Q >�`�>��>�o(��[��.A>7��>���q���Z�搢=��9=��=$��=�ɵ=���=���q�P>Ḟ���]��ED:5��=i*c>6�>��C>��0>��?ߚ?e<!?�_�>��v�ك)��d�7���>=Y=�>�L�>*�=�w��6f�������H:���d��h����>!B>�	>kc�=�(>�=��𬐽Fh,���ҽ@_=�t;�p@=�{{>�җ>Bݩ=g�!�(���iD�Av����cir��^'���A���v���a��;�.Ͻs�C� 
�<fI�=��_��W���=2 �����<4��<,�	�yY>Jhk>��@qӾ� 
�'����7���nU9=�)�y��K6���to� ���*>�D����,پ7$ھ]L���6�=�M�>Ř�=��p>��:?Cz?!��>%>�]�{�q�g�>��>=|�=L4��ݭ�%�\;�f�>��>��X=�G�i��s=ց�;XgL��l>=+�>3���X���$�[�=�B�=��>���=r�*�Qqm���B����=�τ=���>2���_��I���G�9�=�<�>"َ>?*�=�PI>�Ѳ�p���o	�+�j�o�?=�>F_�>rNs>��X>�ȹ>EJ����y x��ݽ׾*>룯="[�=I۸;'��=��o=��/��U�5�
P<���ަ=��>1�(>�Vz9kI?]�6?`�?��k>2���v(��祾�ȭ�\�=P7o=VO�>2-�>=Zf�]`���7�0��\�1��ݐr�X�|=é.>Չ�=�>k�<����井��f��E���%W����=���>]W�>�>��|<���e�0,����ŏ�Y�ɾr�߾��6<}U��_���7�����>���<m;�S�y>�h�=ͻ�=J�<�@ �N�w�`�z�N>�C���Yl>�Q=R������K���E¾�|�0�<���;o��k���g�_"�S1e����nw�4�������>.l=�_��0��>*�? d�>���>.\h>7���ö�,x�=�bc�D��>m7�>6�
?y�?2�>��>ܦ�=��;�U�ǽ*>%_5>�h�=е�-�7>���S�0=J�M>G?�=�=�Q��m����F�/�=x^>����T�<���>��2��YV�\>F�<��,�>�Ӕ>�h�>�W����{�r"��ʾ����a~J����j�`Ⱦ�?v?H�>�jH�x[�=���=�7T�7��:�8|>Ii�=X�\�!�>g#;>�"�=�a:< TѼ����=eL�$i�=�ה>�D>	d�>��?P?pKF?��<',�L�����^����k�=%��>���=o�W�=���ȭ�>��
嬾�#����(�����+>3�c=�@���?>�!��(VI�N�=$��>���=t|U>M�=����G>k�>L�z>$�r<�/ҽK�0��ݿ�Q��`H��8�pB��<���+���΋}>=&P�5H�牾��=Q>hi�>�	�>s��>,�%ˆ�!�/�m=�{o��h��䠾��s���˾j|ά�o���#P��?Z���п�-�i�J���MX�H}�����K�h��?�>̲�>iI
?0�M>��?eSZ>#ko>~�����Y>#U>�ֵ>(��>�ZE>��>�� ?�` ?��>�\�=)<��+7��e9���3=u�7<��:>��e>�Ej>ɵ߼w�D0��-� �T�:a�,>����%�
�lؽn�=*�1=�Z>��>Ǽ���o�TP�d}�'�J>�y��>�����̠�ՠ}�؇ݽ�*-�q��x�о]-K�,�̽���>ү�>9��>���=�=bx=X���+m�=�Q�=)v����J��K5=�y�=�����ὶ������E�н/� <6T=�u>�،>+�?@�>�*3?�:�|� �k�������9���>u՛>Z��=E����l���ʾo��ċ��]��v��Y�ʣ�=�!P>�ސ=��#>%��s���E��;\`>A2��Ұ����<)0<�|V�=2>�U>��n����>�7����¿��߾��������$�kr>�D)�{�F��I
��)C�i���cX>+��>�$>()>��>A�=V�E�m;0>\�2>�9�.���1-����
���ݾ���>.o�=�H޼���Q3�=�^�=Pt�<���=MΎ�ZbW��$�0BC�Up�=y��<��?s,g>�-?��>p�#?"�>�m?%I�>Nۘ>$�>��?y5?��??�K?6?��U>���-��9���/.���!��<�Ƣ>��j>6�ҽM G���=+j���i��Ib=��t>���<.�뼭G�=�{>v��=��>~�x=F��=4��[��!�>���=�<�>�o��,���<����>W[>�4]�	���X��J����>=<��>,H�>���=�&�=�Y�=5����J��0>�e
>|o�=6�3����=�k�<�qO�q��=&�	��/c�ܲ�R�>��T>՚u>?��>!/?�v=?l�������a����C��6���5<UMj�|)4>�����������:˾��F%��6��� ���F>�襽5?<��>aM�=֛����;�1>b ҽ//;;��4>��%=F����=s=S=v~=11��{���5��|ٸ�a�2��5�����<����O�=�O�=����f�>�ԫ���@�\d�>^]>?���>�>��:?����Cƾ�ま]]�i�1�jD������I�箾v��<�y�抺��9o����F۽�U������g��ÔA�DI���	�^n�>�0�>���>�;A�Cs?�=Ч�=e�>10?�L;>Fȅ>�=Ek��C� >�c ?
�%?�b�>1�?o�:��F�������>P��<_�H> >[=�> ��p�e��q>��=K�#�:�=w.�=�
>�=��=����ޜR���>�|�=9�b�!5��j�ϔ>ٴ�����>\Cؼ%),�w�Ǿ��-��:�>��>�Ұ�c,��T�z��=��>t�>L)>�4�<+��<Uco�7Z���H\>�L�>Wc�a��
ߌ���8�Թ�^��ʇ�L����I��>A��>�__>���>~$?�v?Z� �<8��a��ľ훵�z�Ƚ��><B���Ǫ��_��R����3� n��r��=�f����>�Oz��H����o>Lo/=��"�=�ą>�H
�.�c:�,���J�<œ=U>h>�!>)���lμ�v����ӳ�~�þ�-�!�<�`�=�P/>b�� t�&�v�3��:Y ���M> �=��f>';�>��>W�x�B���za��G��>� ���t=������ھ����y�]�!����=LDF���&��K�*y��V���߳�Fxy��.����t>�iP>; �>.�����>�X�>N٪>
>>Vs	?��>�O�=q��>��5���'>��?l�?XT%?� �>�/���UF��z��= �S�r��=s9<>%">�J7�^UX��3>��>��>����I?>��=k\�<g�>�R"�������>��=�]N��!�!m��ŉ�=�]<�޿>n=��1��]Ѿ���)=�;�>����"��H`����m<~j�>�!�=_�����=CW�P�=c�3>��N>����y���Mw��3:<3V=4������s�J�m�b=,�R>�g�>�ނ>��>�P?E�^?�����������h�7�;�=O�>�.>�������+���A��n����>�fj��0>R� >�{��]��>�QJ=Y��uȸ��a:>j�F=%�=�֢<7�Խ��1>�>�%$>�}�^s������L��;�����]����>��%>���=/�⾯8��=�ܾ��l��>_/�>�V�>�}~>��a>��#�Ѕ�묑�$����+��
�{�4�;��$����e�0��7�F��H�|��)�rp�=7>U���>���v�[�I���uN~>�.�>�u>tlw�ц;?镎>��S> ��>�R?\��=ݨ>���=mPo�-�w��%�>��?�.5?Hz?����@L�~�n��mP>B�>�ZT=m��=�}X>���Ψ@�3��=�z=���=�O@�!�9v��=Ո�=���=�)����x��L�>�������OB�՗�P!=_������>�C��q=��"˾[25>	�
>jW��'˾]���Y�/X9>�"�>�,�>�Z"=���m'��0;X�l`��Ͷ=*A��s�=	#�=��;>F�=�ٽ�C�;���o�v�< �CH�1Qq;3 �>�)?㐸>�\;?�%/>�̾4�þᔿ�
�o�,=י�>ї�=��=�R
�/鰽�����T��/ξ]U���>t��>1/���>�	�=�fV>+�>���`�׻�6ŽJ|>u5>X%:�xS>�V>�;�K�ѻ���T��a����0þ$������Z�E>�B�=��؄g>�콍���?~�>"��>�ݰ>3�?ò?�>v�;\�>wd\��Mս���=�P���6��پg>�l���� ���R<��߽	�=����MXS���Ì;��%��g�>�0�>�}>�v>$��>�բ>?h{>��m��;o>wļ��%>�^H�|<@���= P>�S�=��l>�[߽�M�=�m;�����Ѹ=Wb�=�c�=���=x V�����c�	>L%>� ռ�D�=�d��v��ﱍ=�n�=),�=�� >'�=��>�B��	m׾g9�����_��<�Y¼t�>:e�}����W�a\>/�=i���.Ǿ�濾T�Ͼ���>�O>�>�����y)�ƴ߼yߋ�Cf/�=�?>��>֗>FK><>��3<e<�=d������7'��D	>��=�Mk>�?[��>�4?,~�=񥅾�4�[&⾡C�۵�<�?�=y�%�r���ﺆ��ӫ0�
b�dþJ�D��k���n}>V�=:o�=��>��=]Wv=q��<5�z=m�q��oI<�ჽ�=�%�>M6\>��>$�(>�-�FP(�;<��ؗ��茶;-!��P<=��<>�.���N<gU��8F>������!�m��;��=B��=��[>�J�>�jm��<w=�[�>���k!�=�D,<m���7�	�ؾО�ۑS��ju� ��GP7�ʢ.��Μ���L�ƛt<�4��%��0 ,��r�=�*�>��>�P8>���>�5>�YU>-z��͚>�P�<�8�=O���Q=Y �>���>���>��>�_>��
����8+�H_=�\��1.�<gb>�.=͓���۽�$�;O����^���L�ظ���^��Òb>�*p��-����=�|�>S9h��p�оM\��'>�I>\<w>�᪾�o^��ĭ����=�|*��ξ���9�'�վLD���^>��s>a�=��m��#�=�ZŽ�2�����<�F>�Ｏ����>>��=����=��;��hq7��5��z�>��=:�>�#?\�@>�jQ?���<LG���
�gS�o�ϽH:`>�<�=1;L�^M���,�>޸='�o�ۦ�m!���M}��OuU>�A��I���h�>�<����)���%0>`�;M��<�!$=V�}>��`>Xƹ>;�&>�8/>ΆA���G���ڿs�al��j\/�������O;�����u@���c>��=Ƅ���U�=H=���=��>p�C>���D2ĽM$��rս����a<���Aӽ��`�3d>�!h�2Bj��W�%�
�a�UN��&=��-��c�F�_��t���=���>h?��s>I\0?�b�>�=�> 8�=y��>Qƌ��JG>�4�=�>N* >N��>��>	�>r��>��6>0:��c���)�=����O���*�=�o�=/iw�Q�<p#>�̽�j�D���6�M=�9<7ε=ً�=%3��U��=�7?��u����|N�xF���|�=:[̽i�?��Ž�F9�I�<ԣ����ʾՀȾ<��e����>�J�>C'p>��b>W�̼vʗ=�[��<R<��O=6��=&ռ�t������~�=h6=����Q�%�Hu����y�W��=܋d=�{�=].�>�R�>m�>q�-?k�v���l��A���Q='���R�7��ù������=��%���+��	����j}K��\���.�>6u%�F�>{�>��d<���<�Dz<c�a<��S>˽>�F�tOF>C��>G5�>@I<!.>d:N=.��RBͿ0������蟾7X��]ܽ���>�pӽϗ����	?m�=E�ýH�>�s#>ص>Of?���<����1z��=�U�j, �>����ޤ�����͜��T0��F;8��|���a���_��>ռ�X�g��z?��F/���@�R����>�%?���>f>�?�,�>ʫ�>�:=�B�>�!w��<�=yL>_�j>�dk>�˨>鹢>�{�>{>�wJ>j�9�A�-�	�=������=�h,���=�F�=M��=�+ѽ~E����x=[��=z�3�����(N1>�=E�"<fE�=Yl?�������]JL�̼�~H�=?��>Oi���<���@>D+�<8���E�@��h��`�U>]�>}�M>6iϼ`�1V��G�==��(�^o<XG<�݌�������<"G�=^Z���̻ސ*��X���Z�=��0���3ZM>Un?b�>Z&?`^8=��$��8U��i>�h��������\#���c�W��=�3�� i����牾ߤT�DdQ�4'q>���<jp��)�=o(=\j
�@��=P�=bq�R=��W>��>W.!�~Ӥ>���=cT;�O���썽�bѿ~*����Ž�Cݾ�T6=��=�NA���н�UM�3�=`�B�ؤ^��>��5>���>�Kq>�g=x�������X/>�s�<�!L����"��L���� 	��ý��߰ >�=�8�#�@�0����N��z�6��B[���+��3�G��|�>��>ae>'?�%>���=�=�ŭ>c��<_�5>O�><�\=IN�=��?�-?���>z��41���X�Et���=���=��>�v�=��=>Z�6��_��W%�=�դ;��@��I1=�Q�=�Ua�c<(=T�߻���>O3-=�'?��=˝�=�!�����ؾ��>�Jξ�˾�W���؝�wH��{Ͼ?��,Խ��$>��>�^:>b~{>iY�>�
�S}I<&�̼��"�u�pa'=w�>s
v����=�=S:=�uG>�r$=T:=}��p����D���l>��B?��>^�?oH�|��;�"�Et�����;:G<�ɨ=��1>�y2>v�U��:x����+2����҈���>���>�?�>h��>�> ��>�����=�ཊτ<$�Q;�,�=%<5�t�Z�yql='��=��=�{���aҿ����ݾ�H"�<�+>/R>�%�>�ɕ��8~�'��>�y����#���.>�X�=YL�>q�*>T���CV�X�����ֽuo
��7�x�o<�� �쳅�����,���:��h�ͮ���!����B�񂐾2����L��^��tW���ʽ��L=	;�>��?�<X�)=?�s�>�0?#��b��>	��>��>9x�>U)�>�E
?�n$>��>�u>i�����>䜄� �������1x���_>���=p+�=�!�=c��~�>̆н��v���Ͻ��<�<=�\�=���=�c>%��=?iU��~򠾨J⾳�����w�1�
�>Ⱀ��q�c�#��ξK�	��
þY���j�>;�>�-�>G� >s��>:P">����%���<>&-���׽��=W�>�Bp�G,�=��=N��=�f =� ���F�=HI|��qܼ$Y.�7e>�SC?e;�>�\?r��?߾8'��oV�N1�=��=�(�<S�=���>�F>*y2����"?���/�yY	�e6����m>��>R��>�k}>q�>>0H�=&| �d-��
�� f�=��">Bf�=��P>�
�>2��=�\�=���)	|�xIͿc﬿k��z%��g�ڽ�>> ��>�"�XIY�]{>���jf�z�>|�:>4�]>��$�c+���ƽ�]	>�F���� �p�`��<�'��Y�-G��� �N�;���;l����\ؾu���`J��5�ҽ�5W�������\�9���+��w�>���>�U>��Z?��#?*î>����;�>�vD���/>d��>�{>�W>���=�� >i��>��=I�9>�l˽^�\�Z0��h�y��f��.=�.<>-�<5�L�3��=�*мG�0=*T��e��'��2^��<;�=�I>
�>ZW�>�> >6t����Y� ��#$����<�Ͻ>�O�<��>l�<(%������
�b�վ20��v}>|�~>�E>zI�>|M.>=ε�}G&��B���� ���ּ��>̈>��/>�N<6X��1�=g�<����S;��=q&~�꿑<W�l>��A?�P?��'?J@|=��I�A����7�В��i�E��5��������3+������B澖�þ!?��n��.xսf�;4�>�ş>�Ձ>��>'=z:��YI��]x��_5>I[ >�,=-�'>�y�=U��;f��=��<�t:�Z�ʿ����޽վׁ���<�T;���.>.f=��{>	�+�8|��ݪ>�?�=�>g�>��q�-iþ5ۋ�;A�>ѪH�ʿS���'�f%� ��(R���_��z��Zr��9O׼`܍��&7��U����p��%-��,�&g[�|ֽc%7�]��>W�>v� �R%�;���>=7?�|<<��e�c�S�wm:�Rn>)߽�� ��ф>�?
�*?��?sr:>jXe������<�p��Ih���>}��<�>V׺�<��a'�G�=z�>�Y���?�jZ�ג�<y��=G#=�Q�=&?U�ƾv�	�[㩾�����h��t=�(��=�p���ȋ�x���k�����u9��N<�5l>È�>���>ײ½�B><?�=%���l���=��	��AȽ�n���:>-���qy�=�>-n1��D�R�(w��я$�����`��Um�=d#\?��?��?���=mþPg�&M��=��[�X�����'>&,�=��������%1��bL��SD���н�f־�U>;'�>���>JE�>�?>} �<�L��4�=e~=�9�=���XȂ>��z>�	�>�ZD>��ؼ����ҽ*�ѿ�󛿄��ߦ�G>�Y+Y�eAe��e1=�4	��	w=i�E�]�*�P>�c�=i>RSq������*����I�>M� >{�b���>Tn���d��ׁ�|��=�찾փH=f����B��J�M��'s�틾�&�U9>�y���r5����>�?Br�>u?:?B?]���>���>�'�>'��>*�
?�;�>��j>�^A>�=&c>'�`>��{谾�rZ�&�_�����\��=�E>�:<�0	��Ռ��v�=%�>B��<K��� �=%�)=�
>K!>Ʉ�=,�!?�M����ᾈ�ʾ;b�Y������<w	K>b�7�1;ѽY��=&Zľ�t8��}#ֽ��>��?�{�>a^>Ő>-/�=����73/��8μgdB�� =�t�<Yj>d�=On�<Eg>g5&>�S�=+�U��#>�틻"⋺��V>dOy>�6?o?��?�>>�i����	�k����:[�g	s�� =��`>��G>q�0��ھ�,!��2���&���ν_�=���v>���>_�E>�8D>�j�=�/=�"�z �锾��=w�޽����;�=��$=�����=e�żVd��Z�ſ�������
�����=Q%�=��>x��=Qkn��A�>������=rT+>�� =�q>P��<�*����D�޷���TjJ���(� gG<���s9v��/����=��򍾞M8>�.^�!!-�����h�� ����8��/���Q� K#���>��?!Q?\�>ʹ-?�v?R�6>��8��X�>ɠ�=�?>�W>��>�
	?n��>�!>)�{>̦�=\#C=�>̽gtJ�\�{=��}�k�=��->��>���<��=&��C{�=�?6�|D���x<���=�E>�>�mb>ٸ>Z�>|��'%�]W׾�?���нV���>�.��u��=��3��J��B�3���*�IK(�v����dѾ\�N�k���"�>x&C>�M�����=J�;[g��<8�=j!>6�={�=7!����� ��=RS\<���=�>6>o��\>�[5>�1>Z"?�0?B�;?��x�?�(��&��_����Tj�	+
�N��>�(^>�΁>6@<6Y���G۾?��Dݤ��5����<\a>g���k٧�<B;�Ԭ߽51c��*�[�ɽ�����>!2R>?�<>�><�R���>A�>m~c�y�w�����%�ֿ$�辠[���;
/��]�8>Z�U�O�ཽ��=�9��n��H�ܖ,>���&1>5v�=z�>w�>,Ӿ��˾�PG�jɃ� u�����G��Y���*�>�I���T[h��3нSG�5��/���D�M�6�LĿ�ec)��|�=tc>��u>�4\��]/?|{"?HT�>���=}�f>'҄��Ƚ��x>��e�=���>�0�>�6/?�Ε>��>f8��˽���=l�>�>��0>-��=�i�<�=h������n�������д� �=`�q�6�D�=$��=&A?����4WD���ΈO�
�r���q����>�m���-/��ǻ� �ӽ  ��>���=���&쾟�߾�8�>�Tf����^4>���F�0�AQ�=������6<��=�!:��rü�q��T(��)^v������F$�W��+g=���>��?��?WA?9~�����s�Ѿz��*J�=>�>,�>4�>y�ϾM��qϵ�����oh����þV ���ݨ>X��=/����sn>�]>�B�S=�i�=�pͼ�Y&>��<�[[>���>;�=��\>�8?>/G�<#4n��ۿ�q����ƾ3����v=���=��x�djD�ė�=��L�vq����&���<�>�>8h��r#>:�=>T��>���>	���bŽ@%�<�6��7|���l�*-���}=�&��b#��:#罆0&<W�slK� Hd�2�6�>w��(�n�O���k>���>���>�
�=�5?�A?�M�>>��={��>��	>�ڽ��$�*�z�Ǳ>Vؼ=�:_=�R?�8�>�˞>��'4"����=�{�H��=->��j=��7��ݯ=[��;�R<=��޵�ȵ�=8�"�� ;�Ib=��=
��=ؓ?�=9>������L���;��4<�k(>�?�E�u(��L~��2S%��;񽎖	����:�>s�J�ڞ����}���`>7��=���=�}U>w>��i��*�<;�f���5�=,�����)��	>����ڧ�@�����9�]��h���>2-.?6�.?K�.?��н�)g���A������'�4N=�#?���>�>����?Խ���i6����x��aC�����=Q�۽�^]��4>�>����,>��GnϽ�P>D��>5�=w�=W�>2u�>��=Oӊ=v�T��pտ�����������}�=�h=];>�M����>�0�>X��_��v�=�w6>�K?>ѵ>wm�>DG?��>�ʛ�n�<�pQ���sB�aMӾ.m	�F�v�<o��8�%�z����`���[��
D��C!���=�<h�������iWx>-P�>{��>�9��1M?0?�K|>����D�>�h��).j�P.�>OY��O��>[[�>�a<���>���>��>��`-�&k�<pP�=I&�=�L>#j3>��ͽg�8>��<�+�yTc����h�O>�~��A��Se>b�w=��`>�6�>�9�=����A۾J�4=(Qҽ"�W>^��'M��I.{���۾�wǾ=�*�Xح���=̬)>'�P=��=�@>�y�j����
>8i=qoͽ Ez>&��;�
��V*�\=	��}��^�=vu�����=�ǃN;�c� oa>��>x�:?b,T?�Ǿ=��$�8[̾w侶����=���>z	�>���>I��=ok���r�͟�������оb��9>�G��k׽��=�� >�S-���>[Ű=��X��T�>�=*>g��=t�+>hn>:��=O�w= i�<lH=Ë𿵂��8I��2���,�L*L�ϴ�ocb�E>�{�=^E���7����" ̽���=oM���/�<���>nz�>��>�T�>^�`���1��1��J(�`Uܾ�н3 �� M���Z�CP��Փ�>pW��̲�2�1��Sr�	 @��@��Q�d>\�}>*��=�մ��?C=?џ�>RD�>/�>69�;��'�^�m>!X�=�>��>E/?�(�>��gmx=oT�����-�=� 7=���=.�<�Z�=,s�^��=Q�=�k\�w�<�O�;����?��ѽy0>��<E�=��>s*���%�����+�";���C�Z>�>9��=ӑ�>ī~���Ҿ<�8����2@�d秽a���.X���넾��>�j�=ҍD=L4	>��<�����(�=p�]=�ӽ�+>5��=EH���7={y�>�-��	����?p�|-��dE����>�U�>�2?��H?g����=�0�;���f1���@=c)?��>��?��N>)~�7>꾾�W�&������'h�>r��q�2���	>��p> ��}-4>inN>Eh$���_=��>,�Y�G2��M>�˹<2nJ>a��=d�=���¿�о4��%='��=�$>�UD����:��<�>����M�cZ���<>:�=�싽�,�<��>��>�2���LW�:?��u��)�	�-�����]�O�����2=��˾��1�X�p�)���Fڞ<�����ž��An��q�>*�>��>Ư���?8�?�s�>OĘ=d�>�
��l�<�ް:>��v�eg�=�>@R�>N3?��M>���>�����G��9�= �=1��=�@#>�_>�P���^�v�/�;���<ˮP������b��B�={6V>n��=4��=M�>������aϾ:��ϩy�k쩽M0~� ]f��v<>,U���<�聾��(q�����6�<��>�\�=UF�>!e���R=:��=��	�ZO�Ƥ�=�z>eyѽ�;ٽ0X�<'E�:�`��׶��*r�y*����<��=`>�+>���>2?[��>��K<U�*�""��+��[����۾ڀx�!���q&���=��Y��ԡ��A�	�������%潳�z=t1��
�YT[��{�IC�������2>�	�=���<y>Y�>�Պ>�
�>p�s=�0�#�	�L��=q�R���H�ݾ.a��𷽕) >}V'=jϷ���
���\>�w�v?�����=��>�d>���>8Ɯ>�d>,n`=�MH�O��=��I�C߅����-;�	��r�p�ܙ��r�<�}��І���x�&��#$���н�6��������y)>D�>BW�>Yx�>�;(?fu�>)��>'\�>���>�I;=a�}>xaN>��>�>�J�>,�>�7k>�mS>�(�:��W�JXA��$->=�<>�@=>��0>8�����=%}<�O�9h�<��`�܏���NB=��4>�/�=��=�7>�?X/O=�Ӿ~��|~�(���͙=�.�>h!��n>Vb�$���ߐ��kӾ,ƾ�E��
ܱ�F. �V:>ٴG>j�~�*~�;���=5(�=m��=̌>���>�~n��ē��B�ra��Qx=��PW������;�d�,<&�G=,�_>� �>�m?��C?2(<?�4�޲�_O�\���齇��� 라�}>gSH=rb�Nv��ʧ���ﾅO��ľ�)ϼ�������{�<��ս�VT�4�=y��>�>���=,�U>��}>E��>ڛ�>��>��6>v6�=��$������ҿ鋗�����@�t��>l�y>��<�4�ߢ�,�<���ӆľV>��?e��>4�"?��?+;�>"�=8P��r :=G5����Q��J��g����s�$��ķ=2��֢�T���6�]���"�-�w�E� �f�Ľ��>�>��v>ذ�>��>hm�=�^?l
>��> c>��>�!\>281=�?&>�$~>#�2���>wH�>N�3>��C��;==q~>�g>2��>�{y>�a�<�H�����=ZK>����A�|8&���Y=���=Yk>>�I�=�B�>��=�\�>���������w �����H���2x)> ?\<w�>4[�<52�`=Ϟ��������wq���<=F҇>�`��꘽�Z��ڋ%�����&*��z�>�j��Aψ�6M��s�V���&��x���,T��n�zW��3�=�O7>��=P�>�d?g�?�y�=�"4���|���~e�N���'��R<=&/���.�7�X�,N������X�����(���,���>�ˎ;��/�����G�����<�jA���4>�1���<|Q>���=̰3>���=L��=ڗ=f�S���$�b�>�r��6��1�� �=�k@><�=0����c��F�=��ym�������$ >)�b>�F�>I��>��u>��">��i=g"(>�I ����Ѿ�nP��a̾˝��gP���=`)�<
��몋���K��fB�E�>��r�������|�8�>���>��>�`�>�?���>��>P �=�Ο>�м=&`(>��>�=��>c�>0&>�ٮ>�,�>sTl<�c��<��@>�v>X��>�nE>n��>��=
!���,>��_=������c=Vv+=���>=Q>�vV>AN�=͝�=���>QVþ�\1��o��/0���ĽǄ�$h�>�M��b? �&����� {����̾�پ`V�z.>�@�=�9�>�k�ܚ��k(R�,�ܽ� ֽg��=��>~��=K�\�]��=z >� <�A���0�@��NT����=���> �;=�O?�&? ?DfI>����|q2�)���[���G�/wϽ��;��s<�ֽ��>�V볽�:0���־����o�2��9f>G̿<��1>-E�=tˉ=V�=�C4��l�=�O��8����?�=��>��C>��3>��!>�>���8�������&�����~�<�b->Q�4=jJ�I��v�*�����F��B6F��Q>œq>v��>C��>�=��（ו<E�>Q':�� ��2ϛ�	>��0�\W�� �l��f�=���Y6�������:���ؽ�Ž������,��� ���v>Z��>���>�_�>uG?�j�>&+?!��=�b�>��`>Һ>�oV>����I>���>��>bZ�>�w>�Xn>�Y�0{0��L/>�=��?>[��=I>���<?��j[�=U�h�a�G�/]�<��;�'Q=��=�~>��=kS';6��>O���@�/�u��,t*�l�̾|�;=��>�>Y>�x!>^�/>��-��񠽭}1�HY���= l5>pw>s�;>/��J�c������=��=���=)s>u��Iv�YvZ��==�(ƽ�l�V�^�WͽyԽ����<��>��S>��?�(?�;�>@��=��&����'%�֌9�����Hb��9�=G�0�����р�����E���JӾ�l���b�½<�=���=�d<������=Qw�,�2>�R��3X�=�L�=���=���=�a2>�q�=�J�=�9����R�9��󖿴/��!�#�	��>��	>h�><߮��9�5�20C>&������<��a>@�>�6?U�>��0>�ؽ��I�>1�>��ؽ���`��?K.��ƾJU �����۳=d���z�˽���C
��r��Wa��8����C���ɽHT>�[�>Ut�>e$�>�*?~(�>�4?h>�<9���$��������>*Ҥ=ܡp>�J>�l�>7��=��<H���t�C�2��>&5&>� �=�N=gR�8��=W�>�u>��j>S���n�=g�>��>ջX>�>�;>���=j?�pS�L�3�v��l�F���i>��?��?Β���Y�
�>��4�����%��@��@��Cվ5�>�et=��5>�i#=�DH>���<Γ�;B#�n��=���%܁���>A�Q=�s+=�U�Q�S�'8�c%"�Q�?�;(����ѼVa>��>?V?�8?ZZ�=�X,��C����֬����>cԅ>I��>�ܚ>�<�=�y3�!H��������*��t ������>��7��;�*�$�v�[�����= 
9>�,��>(H�=B?���>���>+��>�<=����	��tC߿ޤ��&���p6!�Y� =zE佋Ia�����ӥ��&O���г��z�����<�j=�ϗ>B��>N�>�T�=T��>4g>yM�}���I�3%���U�;�$�+>�z���[��9?b�����Z��:ud�>�Y����#
���9���>y3?EI�>�u�>�??��>1�c>�ڙ>�?XC�����(�#�P��>�`�>Ӻ ?<�?��?Nu!>��M>�d��ئ�Zן���= �Z>��7>W��=��ؽ�|>�^5<�?����.ӽ׉�6lJ9� �_��=yT�=p�j>��?��ؾ�A��a��;��X����>m��>�:���V��=�۾e4�uu��� ��2��8�K�P>NZ��	�=Z�>�r�>���O�>*�ս�Z�=b��M��ߢ��s�.���=�s&=�4�*�Y���~f���B�=in�=��{=֜8?,Q=?�/?zs.>#��1���-�o0��v[>���>�$�>,�>J����2��Ӏ�F��$�R#ﾍM���g>�R���=f>gve�9S����>]�=7
�:|d[>v�=�N>B~�>���>o��>yU>�¥����:ÿG������o���T�6$5>���=wYE=<�^;&�x���	��<���כ<>\>��(>�\8����<��:>�+*=i0+=9�������ᔽ^��`���G�?��=�p��*~�=�`�`�%=�8���"�����G����Cw�����k����>3\?�غ>F?b6?�a�>�����T>�?1?Í�<8�>������Q>nw�>�(?D�/?L�=?��>�²>Y*��s@�I)K��P�=-�>�D�>���>�G7��f>��ͼ���������`��[��!�j��x���:=�?=%�_=�#?ń���;��,��,5�x�<>y˒>��/?ܷӽI��d�=�<f��r־�gҾ3 �M��tv��͝�>�%>�@��l~3>�yG>a�Z�^�a>��A��Б=�A��R�G�1��<�L�<�v���?
�b�����a'���g����+=@�4>�H=`�C?��/?�b?��=�	"��I�ő�nz^{=v?�>7Ȏ>&&�>fCe<��GƩ�
��i3��ݾD#��^>��$>�Y>���a���6�ɾ������=D����<K�>�P�>�>bH�>Z~>(O>�t��T����ÿ�������%W����yO>û����ʽݮۼZ4i��l���A���M���,�=E~�=��u���>�{Y>���=��>^�ٽF=��(m�:��d:���t�f�>�ϽZs}�Q�y�c�>Zoǽڛ0�@�k�V��Ƣ��!�3�ON���@_>� ?�o�>���>�+?4j,>�]�>z.�uM?�k�>������=�*�>H��>�?$�=?��6?"�>)�7>�7��)[�����k�O�>���>�J�>�`�=2 >�H�<7	
�*�M��K�5R;Z�Ľ���=���=��=��>j?�pS�L�3�v��l�F���i>��?��?Β���Y�
�>��4�����%��@��@��Cվ5�>�et=��5>�i#=�DH>���<Γ�;B#�n��=���%܁���>A�Q=�s+=�U�Q�S�'8�c%"�Q�?�;(����ѼVa>��>?V?�8?ZZ�=�X,��C����֬����>cԅ>I��>�ܚ>�<�=�y3�!H��������*��t ������>��7��;�*�$�v�[�����= 
9>�,��>(H�=B?���>���>+��>�<=����	��tC߿ޤ��&���p6!�Y� =zE佋Ia�����ӥ��&O���г��z�����<�j=�ϗ>B��>N�>�T�=T��>4g>yM�}���I�3%���U�;�$�+>�z���[��9?b�����Z��:ud�>�Y����#
���9���>y3?EI�>�u�>�??��>1�c>�ڙ>�?XC�����(�#�P��>�`�>Ӻ ?<�?��?Nu!>��M>�d��ئ�Zן���= �Z>��7>W��=��ؽ�|>�^5<�?����.ӽ׉�6lJ9� �_��=yT�=p�j>��?��ؾ�A��a��;��X����>m��>�:���V��=�۾e4�uu��� ��2��8�K�P>NZ��	�=Z�>�r�>���O�>*�ս�Z�=b��M��ߢ��s�.���=�s&=�4�*�Y���~f���B�=in�=��{=֜8?,Q=?�/?zs.>#��1���-�o0��v[>���>�$�>,�>J����2��Ӏ�F��$�R#ﾍM���g>�R���=f>gve�9S����>]�=7
�:|d[>v�=�N>B~�>���>o��>yU>�¥����:ÿG������o���T�6$5>���=wYE=<�^;&�x���	��<���כ<>\>��(>�\8����<��:>�+*=i0+=9�������ᔽ^��`���G�?��=�p��*~�=�`�`�%=�8���"�����G����Cw�����k����>3\?�غ>F?b6?�a�>�����T>�?1?Í�<8�>������Q>nw�>�(?D�/?L�=?��>�²>Y*��s@�I)K��P�=-�>�D�>���>�G7��f>��ͼ���������`��[��!�j��x���:=�?=%�_=Ry"?�V���s�'��
$�9�=��]�?�U�>� ����=���hD���%����g�>#?[2%?#9�=�;�=��&��~p;Ҫ �. �=x�8>'�=N�2>���a<���0����;�	�p���?]'���=��>�Ҵ=�,>���>��Y?
�>Hm$?X�g>)	�š��"%��哾�=�r�E=��>��>�k4>Mܴ�](,�u(-��{���_=5�o�L�<���=�5�����j����f�<�/��T)�=j7b=��=�t>&�>��>�v>�b�=�2ݼ���=e��JԿ 咿h�����FA>�X�>�p>�b5��T<���>� ������Ρm>]�z>�uS>7�>���=���<Q�1=Ơ�>�F.>{��]|�fE������X��Y��>����>���o���3���(������%!��	q�%�-C���Y�>���>�Z#?��>s��>�>}w?���<���#2>��8�g&|>�/�>8��>��?���>�30>i�8�ę��[�(�𖝾�MZ>�E�>
�\=C�:=��=e�wn7=��C>)��=ʂĽ���l��jٻ^̅���=�&>$(>�J	?������о܂��F��DR�<�l�S��>a�T>YA��:
{��v�Yk.�}��_�3�Ѡ�>3e�>�q�>cv���.>r��<�5�����U!>.P>o�S�Z�<�=u��{'1=ܓA���v���$�ŗ����E=�cG>�[#>46r=��s>��0?�ڙ>�d?�T�;�8$�O�⾱a��H۠��1�=q�>3��>� �>��i=���
=�տL�*a���">Kʜ�*�Y�H��>^=�=S�N�&�ƽ<w�<�\d�����2������HM=��)>��%>��>��K>bс�:ۃ�+k���ݿ>ߗ�n!
�E����=)��=Hǻ��H����D
'>Ҽ��¬ػ�)T>d>}�>j��=�܁�_����=�z�>�1�>Q���a�Ͻ�����
�ྺ�?	>�3��=�~5��P�_��>�$�c��T�G�O�L��4$��2����=5W�>��?��>���>R�?��7?�>�d$�>HT%>?(>^^�=o>�>�?M��>%o�>���>X�=��+�Zך��7o�߃�=���=�pb=`�=��>�!>/L=&}=�E�=��>>]>�_'=<Q����|ln�&>Ԥ�>AC?#[�����3�����G��!���{?p�����Ǿ<C���9��B>��c.={�=K>\>�>	�>���>�e�>�����4�y���S`?>]ȳ>�>��5=��D�=G��=��m2����gn=�>�{>u��>_��=��%>�D??wE?�?g][=?����M�J��և���k>P-=�_>��k>EC���%���3��,4���*���h���/���=>�K�>��)�T���燈��V>G.X=��νrN�QyT=�6>��4>���=pN�=l��T���6j��ߌ��xٿ�'��,�<�����0�>-?e�@>0�(�,ڔ��)�<o�<���>�&ܽTC=���>۵�>��νjB��4E&<��y�c�;=�)��Mj<<�ۇ��%���ƾ�:�
�c ;yXg���̽ �@�>���f�������*B�̿�L��>(��>Z�g>��W>�?�A�>u�>֫9>F�>��>O�m>�4�=�9=ET���ؽi��=�?@��>�"���Ľ�D���<�=Z�=#X�=X:>�@���ȉ�o�{>W�=am>>ƪ�=�	==� =Q�I� ٽ��p=��V>��?�.�X��H�i?���I����ك�>yn�=�k���r�����Ǿw#� �<�V\>l�>>o��>�(�>Re�5g0<"Zﺚ��ů2;p%ٽ*�=��绚��'����ʯ��T�����<�]D=�/�O�l�C��<���=}9v>1�D?Ig#?;��>��=>���)������6ʇ�aP>���>�PV>�;r>����7Ҹ�:AB��E ��?��zW�K���̄>�r>��P>:�=Ò��� >��u��}K�}�׼���=��/>*�Q>9u>PR�>SK�>�/�=	��_Ͼ �ڿF覿����� VT>x,'>�ѽ@~�.-���a>�\=4�>YH�=�->b<A>�f=��'��pU���2>ޫO��A�=E����z�f-Ǿ;�ľ��_��ͽ��D�+
�=������q���ɽ#G���"�����LĽ�K,�q��L[>�B?T	?��2?QC$?>$�>=O�>�(w�!� =�f�<^�>��>�-<>��I;c=QZO>���>}��>��Ҿ�`�z��.��=z;f��Ӷ>�Q�>տ>8V=q��<������?>*0!>�=�[߽^TJ�m ߽ą���?+>B�f>��?�.�X��H�i?���I����ك�>yn�=�k���r�����Ǿw#� �<�V\>l�>>o��>�(�>Re�5g0<"Zﺚ��ů2;p%ٽ*�=��绚��'����ʯ��T�����<�]D=�/�O�l�C��<���=}9v>1�D?Ig#?;��>��=>���)������6ʇ�aP>���>�PV>�;r>����7Ҹ�:AB��E ��?��zW�K���̄>�r>��P>:�=Ò��� >��u��}K�}�׼���=��/>*�Q>9u>PR�>SK�>�/�=	��_Ͼ �ڿF覿����� VT>x,'>�ѽ@~�.-���a>�\=4�>YH�=�->b<A>�f=��'��pU���2>ޫO��A�=E����z�f-Ǿ;�ľ��_��ͽ��D�+
�=������q���ɽ#G���"�����LĽ�K,�q��L[>�B?T	?��2?QC$?>$�>=O�>�(w�!� =�f�<^�>��>�-<>��I;c=QZO>���>}��>��Ҿ�`�z��.��=z;f��Ӷ>�Q�>տ>8V=q��<������?>*0!>�=�[߽^TJ�m ߽ą���?+>B�f>��.?e�&�e����$�ɛ�|��=�X|>�?�F���h��?>��"߾�j>��g��$�>]9�>����rǾ�~��O�R>����q3�( �y)/=U��<��M>��J�^J���J�>�=:�Rw��!>ZHs;T������.����ve>As��7�\>A�	?K�+?��?�u�����^O�=���1��S=��>��>p:X�6;�����0<?���侜'`�%b��zg"=��Z>�'�~w�=���<�]�=���W4>��; t���ʏ>�5��\(�<&�>�`.>#�>g�Y=�;��N��߿�����F�.X�;��=<@��t�=tA���=�K!>�K���00=�6y���^=�Щ��3L>�2>'Q0=�Q�>����~�i"�3�=32������|嵾I7=J����X�_s��@d��_�6b�D�ս"�2��K��
F��u��j�=l��>O�>��T��H[?��A?{�?�!>���>��=�T:�l��=�L�>�
?��>`��>qX9?��?��>�G�taW�
��=�� �})>�Q�=4�3=��=h5�<�&T>X�<E�5=��r�C4z��Lƽ�:>=�M>k���ߝ�>��>��N�͗/�߆���1��'=Q�@>�a�>`J��+�ּNԇ�#ŏ�Q2����<7Qx����=�#�&{J�UM ���>����Db���9�{�c�	>�j+>W}��٘�>��Z��Pw��<=�n1=d�b=ҹ<�M�r>,�AF�=y��=�IK>r�O?a>?�?瞽>L	�ILA�,3�7���t'�9�>���>�5ǽ���M��',	��盾���=ŕ�jf��k>��c�Ղɽ��
>�ǽ<���ͻ!>�x|=�gX��>�:����=��>�	X>��ٻ�>Z�!�=E|�?�ʿѾ����侦�Ӿ\�������=أ	�"c�����>�$�<a�S�N�ݽ1��=г��z��r�>o��>��`>�x��93y= !>'��=+|���L录�2�1��=鵪�%i=Ww¼(1�My޽�О�1�z����p��[���׹��>�e>�zL�f?���@?��3?�?d�{>�?�2���pZ��>;�>gS�>I�#?�G?��@>��4�u�=�L}����<&��=!�K>�P>�����_׽E�,��?9���J>��>n��=+&�qԚ��r
�m�i�ٜ,>�j=N>Z?�ܽ2p��8��Κ)��[Ƚ��=�* ?�?���芼���p��d�S�oU�����=/d>�*�n`��%h-����>T��<���Fֽp���`�#���̼����`�< P۽4r!���`>�_+��7!�
�ͽ�s >6h���E�sB�=tM�>��>��#?�TU?��<���j�O��U(��:L��!+�K�>��=��=8�쾠v@�ܟ^��}%��kb��6��Д���>�ז=-�={o�=�d�=��=(v>�l���Vͽy����=���/e>�8=�>���<���>���������ؿ����5靾@�ʒ�l�@�@��B�A�r�P�SC>W���4=W�f��ŵ���D>_�>3�J�Y7�-^>���=<Ѐ��~�=�@��ȾqH�����=+�/�(�ѽw�`�=�m�dj�������$4<��f��^�5���6M�����=�1?'��=S�C�v�5?&AG?( &?RoS=���>g"ɽ����T-	>�D>�$#?ڹ'?4i�>�<?b��>�̑>����p�X)=��]��&>
>��K>OU� �=��>��=m�$�ˀ��Y��_9��:�]�=\>��f>�W�>�H���d�W,�&8코6A>n�>.�����;�&e,�9Ծ�>;=�r�Q4��*���8�����j)�=�>`GL;�@½�k�`����)���>e���v_>���=-���� {=��=^Y�Nʏ��<c�zg���~�=N�>A�T>P�>E�;?<�!?ط����3��ʾ�5[=�����s�>�_�=L���+
��!sl�����Ӿ$=�=��<�U�'�>x�=�>�=A��=lм�4S����>Cy@='Ko�
 �=������<PO'>���>b��>�ר=sAY��Տ�E��ꓭ�����D��>�sB=��=S�Y��S\��`������>hq>w����E�Z6>�?Y_&=���<B������+���鼽�:��О�zi��C���j���)���[���<91��K�+KY����,Q���;K�1�D��۫>�$	?V��h�ǽz�?4&?�:�>����?�@�>�C"���輦�>l�?f�?�A�>��>B�>"w;�Z%%�܅,<��->�(p>���=[�>�nռЖ����)=���=���<�ڋ�%���-�@�[�]R�>��>(b�=B1"?-���Ǿy����,2�WB_�;	=�1?1@c�h��j��g۾h�"=_�>��A��	��ڈ�Ի����K��>��J=c�Z٪�c����7�<DA>5Y%��s=`Xy�l�|�;@�=�J�=�%<y�D���<�İ�&�l=$��:�v�>�
�>x�[?��P?��O���2��;�uV��tx�£.��)0=)�z=g���#��\��>�1!�ҍ����i����}�>#ft=:�
<B�d>ͥ<�b'�8[>�%�=e$�M�>�+%��v�;�����f>�C=���=��y^̺;Jڿ�0��������݅�J̭�Z8��о�@_��>�_Ľ��:�t�˽��h>vB+>C���n��\iq>!>r�=���<��=��=��������� ���A�;p�߽.˺`1^��k�w9�;4-z<��#��X�k{,�<Qf��j��?7�=�?r><�8w�i-O?Ms-?�A?�r߽n��>2�e=��>�>��>�d=���>ǜ'?�D?�H?�+�>�?��2�����=u���=��o<�@=��r�p������=���bd�<][7o���ܼ�/=�X�= ��=�j$>�?gýH��R龴�a� оV�\>;p%?��Y�i=�g�&A���Sd�7h���գ�K�<�40����<_Q><�T>,�G>ҙ�=���=-�'���=�6e>����sL��M>�����\��'�C)?���U��1�0{F=Z*�>u��>4ƃ>���> �?�!?��Zu���'�X��"���>߽p�>u�>��:����;����2P���Ƭ��u��
>�+C>�e��ƽ�;�JX>^�@۾���6��QW>K𓽢�i=��>�X�>�ߢ>W?��o>���<f������cJ׿�f����
��q
�Zw�>�;ſ	��r���XO=6�>�L��V�x:�����>����
�=�ϊ>�ѓ>Rcg=9����S�xЃ��	�����۟��m��.�'=�2����52�����Kv�S"�;M����D�O��?�x�G釾�Lr=M?���>t��>[P?�oO?� �>a���1�>m����Ԃ�#>n��>�&=�?�y�>��>k���y���$(E�� ���#q;|��I�=d�>03�<�<z<�\���߅=!߆=o��<Y���:-���=�8�=���5>��?��:�f���#"�q�8�RI���l>?�>�>��Mֽ�Д��e��G���N�z��8�ܽ_�>��>5�;J��=_w?�1$\>�=��=���=��>�E>+����<�
�<���6ؽ�zͽ8����n��=|w>�O>8v�>k8,?�&?MB*?�R"�?��V��j-ܽud�hl���>��>-)7>�!=ǖ��mW��2rھP�ξ���q_=�=>l���Ů6=M�_>��+��}��?f񽑋�=G����O�Ղ�=�Z�=���=FD]>��Q<��q=��u�]%���zܿ�y���u(�oZ��Ԓ	?��>��2>D�ߌ���8>�.�V�vϩ��8�=��"?�Z(?]�!>onG=McG�+�7��u��l�1����[ݾ�~d�����@�;f�ս'�<�]�j�}���jT �\�6<�V�@ +��`m�_��o�>�>���=Fψ<�I
?��>���>�"H>WF?U��:�w�=�sj>٣>�␽���=mp�=�>V�=m��>[?��m~w�pKȽ��\~`�,>�=f�>p���NG�=��>���=�}�=�!@;�W>��}��=�쭽&Y�>��d=J�?��9��Ҿ��n-��u��>�;�l�>/���Ė�=O�='aO=����7�����#����%�),�>9P>V@>��k=)d6>v��=rq�=g�Ǽݿ�=1����ӽD��_��\�ཛz��e��?��S����<��>��6>��l>d�?�'?��+?|U��yN���E�ȗ��8��Q�i�U4�:��ݽ�a��d#1>JS�iҾ� 1	� i���*��׾��I�>J��%k>�FB>�V�=�������*��=��H= {>�,->�*>�H�=�>�>Z�%>�׽]-�Iv���7���5-�բ$�t�="���"f��D�8���M���)�+�L<��=�근���>�� ?�==����58�9;�?N�b���}qq�k���ߐ����2-%>0=�yq��"8��6ͽXb���C���p�QB�C%l�\�<� #)�k^;�&�>�Ɯ>m��>��??��?9?��G���>��K=/N��Z<�(�>�,�>�m?���>���>�8�=��ʽ��V�4����BC�/��il=��]>��>��;���=Ԑu=�� =3�>�&!=��M=x��=��->��U=	'���|�>u龥�/��/%�����(��:c��7Y>�޽��,>��=B	�<��=�3ս��pف�k57�h>��S=�Ĵ>�}��G���́�l��<V��<�nW>�}ݽ���<�ր=����Q��6L��j��ю�z�����>��>MI>���=}�?P��>��4?Z�=E�Ͼ�
��n־G�o��]ɾ���-A���i,����������LǾ�!���=?���;�oY}>�;��s9>�}g>E�������	=��！�,����<1��<���Ft$���V>gOr=L�<�}�K�1�T�Ŀ~���($��A��+��ˡ=��9Y������8e>����䩾O=ֽ�b!>��>�s�=8mM=Ё�=�v������>)�~��0����3����p��9S1�����
}�>���b}=�Ͻ>#�:�ǽ>��Z-Ѿ�&���=�Ϫ�>�]�>�F�>� ?\�>��>��>�O�>R[I=�ʳ=@�H>�='>�S+>z?�>
3"?�$?�<>d >�J���[�/�>�½=?�->�W<G�=[e�=��= �H=�o�=|�=Ǝ>g>6��<uH��˩�=]|�=�� ?;s�����~2�k����������>Q=��W�н�V�>)����E������۽s���G�=:>�s�>Ǆ�;Ι��I���*=�!v�;��=�9�;Sؗ���=��=��<`޽�����^{�WM�)�=ci�=�[�=j�D>�b>?��8?=�E?�>,��̣'�]�۾7Jþ�8־zr����{�<I�D������C��S���/�{M��.��|�>�L>�0_>� �>�l�=���Q��
y�=�$�Y�2���%;��=��d>�1Q>�t>^��=M����C,�6�������h!��B�PN��o��F������$���Y�Tg���B�=Oh >l��>Z�=G;��3�=fr��R�>��=_�g=Ad�<Z;;B���v)X���_=�塺`��=���O��ń���5�\�Ӽ_�7������\R��W�=���>��>Y��=�O?{��>���>e�g�� ?%A�>�ђ>@፾/Rq>�V ?nA�>�C�>O�>S��>��<F@O�'��a����7����n=��>~R�<[���.��V�=Ke.=���={��=��=2�F=�l�H�=�-j=E�?��K徾*�о
W�����=�L>U�>~1S�0ze=
�=&飾ukپ����,��;7��>�8%>&�g>���>���>��=*�;J)�=/?۽�����;>ɭ�=+�B=�K�="���$o��,����j�=h����p+>&�*>�q�=�c�t�>Ҿi?O+X?��f?���B<��`�H����e����js�=��2>`Ŗ>��D\]���=���8�@�H( �N���K>�^v>���=�Q>� E>�*���v�
4==	� ��_�=d��>͢k>��2�=i���%̽B*Ƚjx?����Fۛ�شJ��5�@�=n��:ܱ=.Hɽ��<��޼v�B<.�>�t�>֑s>�����0�zR,>�8�=�C��i�u�!���;�˾����4~\���f��2�4<������=0�)-��?�����r��J�8�rr2�=�̽��{�>��>*ҝ>iJI>Cr�>Z$1>���>��&>˧�>y���[_�M�>�!�<כ>�k�>�?г�>o�>$�|<�ߡ���j�_��=;��
��=(q�=���=�E�=P䠼1��e��-a=�
=}�=�C�<��;?U����=z�7>���>�I�Û��2�T��>L�=+�=��;�����!;�=�ȽÒ������]�0�}�=���>>r7�=L�>u�置�9�h��6k�6���H>���=8!ӽE҈=�.e=��	�FF�<];�=���=Y�x=�"�<;����f<}u�>��,?�NC?�9?85>�Y��)tӾM(־�Mx��p���ꐮ��D���N�A:��Nb߾�+ھ~�Z�k��͵̽,�>�+>��>*ǋ>�a�=��������>��m<>��t>g2��#��O�i��{�hi�=e�)=�6��i���:���
�;oG�[��X�׾}���7�=fCb�Fv�>�;�>���>~�%?c�_>�@#=$��\����ؽ�����>���&�,�-�i~ؽڏ��ՙ���԰�=3{J����z1�c���5��*K\��JL�3�,�9�2�؆@���\�M��>�L�>�ԋ>[�"=���>���>�!?�b[>Q(�>���=��ͽ(5��8Á=�r?=�?E ?��\>�����hu�k
��j�*:켵;8�ϼɍQ=2-�=% ];��|�2��Oٽ�Q�G�>��(=p�>�d~=jB�<�=�-=�Z�>h���C?��B۾sW�t?���=4�>Q��=/�>?�*�Aݶ����nϾ�de��p>���>cC�>+@�=��>�?���3�-�^�ߎt�:<>=��>-r{>���=X�=n��=��b<���<�\>� =w/+>�Q
>2��=�AO>2Ͻ�hJ?=�Q?�pI?���=g�B�6���*�
6ľ�
��!k>�L�>˯�=�R=ukP��`��v�ž��������y>��=>�2;>sx>I��0慽j��
K��Y�� H=��
>�k�=�3v=��=���<�D>�Iĺ*��0l���Zq��������ڝ����0��%��Ro��	\���<�"~����=��>�=�����ц��(E��F9���?=�}>����6>^N�����AA�����'X��l�;��x��X5B���IP��M���Hc��Rtܽ8^��U�>$��=�AO=�L%��B�>�W�>���>
I>'��>�\!>��=��;�͑�(�>0g�>��>��}>+���<͆C�u<�Z�=�6�l&<�A=�'�&����t�����<�H"�d���Z�^Z=R�|=��I(��~��U�=]�?��Mp����� �u"b���+>���>�+<��J>�("��(���	�Q�ξYV>��?>�?~�$>*�{>�SF�?��w��p��
���"N>��/>x>Ʋ>W�'>�2:�oK���*�=m���>�=nM�=��x;��/<���z�:?�(?_�[?�YŻ
��N����UѾ�K���a>V��=��1>>]=<�Z����?*��A��H���Ftf����>� �>�n=�JJ>*�D=Ȫ{�ϓ����=x�5�b�<��C>���=���=�A>O��<��0=����i��#������f���i8���>��L�ˁC�ϓ�	��3�1=Bj�J6����3>o�j=5e0=��I�wA]������<�=��&=4������=��G��}<x�8���F:�=>Pʽ5���1�p����:���"��+�E� t�3�~��v�g�==���=3��>���>�e=#�>?`�>f]�>=�J=CH�>Zǽ7����0�<�>(?��:?���>�K���ξj��=�A�p]�n�V�b}=��
>��>��>��=���ݝ�������V='�X=��&��8=�B
�Q��E9&=���>��#?oS���G�%Ӿ�a��l���<��>�,�[$8�A<<����������� ����>���>��>M�>�ʓ>�<�=Xq�vX��=Sf�=��=(Џ=(�=&K�=��f����O����=n����<>��=)d�<I�B=�W<>��[?�PD?z�?%�_�SFG��;���"�|�����KA��!��^�<��<ytN�`�����!�{u��������>S�w>Y��=�m=^0=F�"�)��@�W=<Ҽ���>4��=�ܡ=�$�=��=q���2�<�Pܽ{ꆾ9��;����ˌ �n���Y4��S�:=����έ<�Y.>���Q�]>\Xx>P�=�?�_{���$�H��<˘ؽrȽ봨�F��U��=����NG����c�j<�(
�:b�)�k�a9$�h�ｺ�8�Bᗽ�}��[k����%����kN=r�>��>�7�=��V?��>]� ?o�9>�w�>-�\>��d>.2>��>�%?�p�>��=����	����>�½M����y��1=��=4Ԇ�ŗ4>��+>K���T₽I���R.=�~�;�{��h�)=�� �_�~;;`>|�A>��?<乽��Db�M��
Y=1�>y��>�y��3��T������;����a=�/1>���>�~>�ls>�Z >��_>�&
>��U��B���6>�݄>� ~>&b���K�=W�r�Ҩ5���<��<w�2<j���VM=���
<2�H>(]>�D>�N?]?2�"?��N�~�¾�"���FY3�\�>s'�>m�>�=�=���9�b"
�ܫ����k�9�p9ν�a��ú�>���>�i��m�YQ#�L[=?�'=���=a0�>�ԣ=�h>V�>UaW>7lb>>���Qǀ�����ݿ�Ƈ�O���[��jXX>����m<= >���
�9>+>%[>,���������;��<hS[=V	c=F���6�LgԽ�(e�Nk��?9Ͼ�Ѿ�������u��,6��ʾ�}!��ۗ�t-,�5���xM�����W����Ť�6�>r��>���=i��==�?Ǧ�>��>��=|u�>%��O�Ƽb�=�#�>��>�#�>_}9>��>�
>C��=�#�{�ý�>2=#��=�c�=��h=�f����<�x*>��)=�%:�h�e��*6�0\Y������<7�0=t�>��?�m���+����Ry�$�=�7�>?�K��q���žS�����ҽP��=�2�>.Ӯ>Z��>ǜ>�N=��,>R�y=�|>��HY����=_I$>�1>��=�Qm;�Ż�˟���=���=��7<�N����,�|<�>s�|==�~�6N??<�O?b?�80��-Q�k�6��4�?�>eI�>���>Ɓ�>�BJ���Ͼu����,�h%�����jU��9�<<>7B>��=�� >hAN��������q�;=�S�p(�=t�t�Y:=ək>FЃ>��9>�Z=>�;��sa����Q��y����g��vh�=�0k���`�E�+�gӱ����h�45[��ޠ=!�=~��=e�ٻ�=��]!>`Y�=+m�>����iA�=$H>�$�hG��|Ǿw�-�)��ޠb���1��r_������8�W��rM�����`ok;�(*=�6|>ۙ�=~�{>� �>�?|\�>���>>��nb=Ǽ
>��>���=T�>{,�>�v�>�p�>��>tu,>\C�;�� ���ݖD�G�d�RvA>���=3�D>�m>}[�<�id=R�>Us�T�2����t=H�=Mg�=�����= :?b��ў(�����!
�I��`���ۄ�>��^�m�ھ�ݾ'� �]r�;�j>���>�\?�A�>OU�>@u�>��[>���=wk�2!��`x����=k�<>���t��;"���N��]0�U��﬽�l�;{��T(�<ᓎ��]��Ӟ=A3T? �U?@C)?�i���ھ�8�����S+�[I>�Ε>%�>��2�/���]o3���:������h����w��������h>���=�߳=�e#��j/��ލ�	DL=��>)L�>sʑ>,�o>���>ek>>Y��=���=*�����;�ο�쒿_���t$�=�1����=l2��*����+2>Ѓܾ]C��� �h��=��Q>J�˽�c�e��>xd���k>��t>.�=��<�
A�_���T���oG=<�m�˿=�ވ������"���~��Is�V*l�=�������<��q�B�>Nٸ>��4>�m?�?Ϲ
?��>���>pf>�0
?m:�>X�>g�>�3n==�<|�U>e�P>틝�4����X�z���Vؽ.��=��=�AP=�^>vj�=KuX�g��=Z��9&�	����/�"|g=�<>R?x>�w�>{�?W��<�־������FFH��r�>�]?�H���:¾����/j/��}*��D�=Áv>r�=>MΖ=y�>pYj>"E>>�m�=� 8�)���B}��l��=��Z>��=�C:�������LQ=���<�F={8&=ɉ���ؚ�S�5>��S>���>��?�o?4Q'?	�D�+�����Q�4�����J��=�-b=�p�=HŰ=��M��> �����j������U�'�$�~\1<T<�>���>'�@=B]%�%"�N1¼�9=ِ�>���=�C<=� >�|G>�>{@�=Q�!뒾-
x���Ϳ֋��������d�>��> =R���-=�@�>y|>��\>�%��B^��J>��Aw�n��a�$>�X�����ږ�/ ��Җ<MIz�\��?2w�����5������5M��`��P�@�)�����
N��~ܽ.7g����!��>���>�cM=��K=���>ы?!N�>4�a>0�>�ct��G>��?�<�߼dQ�>���>��"?
�>X�߽Z�|�W�Խ/<¼İ=e��<<y>�(�>��=�/+���+=�\�>�0k>���<���#�-��=���(=��y>P!�=4F����?��I��
�ʾ��ٴ�A��>���>��Ǽݩ�
�(��r�����F��>� �=��,>�@�>��=7�>���<A�3��(0�ӝ����=/�1>��=��<�/>J:c����]�;�1=���=��A>�J>P�h=�H=���>�)1?��]?'CP?�l^;���H�B������1C<b�=��>�e�=AA���? �ѕ����^�߾���XE,=��V>�s*>��=�* >�3�{�.�!>ʚ>��C>���>L�>�qb>��;0�D��cнY2>�woM�Rɿ8�w�����U�����>�t��+���Hm����r�=EI>�J^=�������7���^��Ѻ=��)��=��G������fB�<HJR�^j����p���W�B`q��Z�"!�31��xm7�8�F�V������:�|��!�?��>�l>����ぽ��>�&!?X��>v8>��>�˽� ��5���oX�>s�?|�?��>��=J>O��>�Nѽ9S��u�1=���<`f=�iν��=F��f-=��=�`v<�i����I����lp�Q��=�c�<Mʻ=f�9>��n>�_g��d�~�5�(-��B��IX�>� ?;���>վ��(���<���^�{��#��`��.��(�<>[��>�$Z>��=�@�=�����T���[��_:�U���=� >���=� �=��F��U��\�5��]��Ӭ=��:<�>a�R?��#?�U6?���<w���F_�d�4�~?޾r	.=N�>'�=�	&=����_�ྡ�پč��*������о�a�<z&�<�>���>���<��ɽ���=a��=mp<<H#�=����ٜ�b�	?b�?+W�>�A�>����;���ç���'��Qͧ�����P�=Ue>��ڽ<Y=�o3�=���=d$�XZ���y��Y�>S�>&��>n/:>��>ݓo>Mͼ=F���ќ��S�#@���n�������R>y��<G���������彯���d\޽�4m�
���=��j�u��>CNO>��>ϸ�>mH?��#?��>"�:�V� ?,�>?��>O�=pt�>&|�>&P&?�Y ?J�H?�o�>�2�
�)��QY�ŋ��/�
�N=cC>I�g> ���!��=�td�䲽�08��W�Kc��E_��8�=]�=�/E>�4�>]�`>���:̳.�r%$�{w7�Җƾd"�>��?��ｐ*ھ��3=l����0f<W�F��H�sb���4ؽ��#�Y��>r>b����eD�aD3��JM���k�6����k<���>����z>f7�=����� ƾ�M�=cFн��=�[1>0-�>5?��*?r~T?o����&!���f�t�0�x���:>״�>�l?�4�>,]߾3�̾?����2�ڀ��E��Z��A5>�����q�Q%�>��b���2�=�=q�!>�6���>V�>.^��>w�>	\e>U9�>��b������X���/��l�I�7���K>sI�>�� >Qh�qꝾ	
=�e��?֎����=�x> �z<
R�<��<&B�=��X>r3$�͢f�b�>>�O=(=����T8��� �<Y�9=��I�ѫ%�~�E�>@��r����2>O��1�B?�l+t��H�>��G>�_v>��w>9�?�!?���>_;���?��f>���>2bj��P�=��p>���>{�$?�z'?��>��=q�O��oW���`=3SK=r-�=��>� �>Y��+�Z��è���2��8�>��=r�8�b���g<��P����s>'�t>誽>nP>����5C�n�2�s� ��%�>Ǖ?�d��y��^T�k��=��3�i2��<����2��#�>[.��l*�>�͏>N�(>w�<β�V(��h������o�5=�%�>�>B7'=�/[�:\K����B+�j�|��h>х�=|�>� X?i?l?��[?O豾�s쾸���E'�3�$��ֱ>'2?��M>	�*�X4>��!��/�46�	#X��Sn��A�=e/��n=�?f>j7u�B�T=>2K>��(>��T�G�<�]ν���=�{�>��?c��>��/>����x�ӾT	ڿ.O���;(�F�ƾ�18<�����޽w������e��=�_&���Ҽ_�>
:�>OC>UG�>.�6>�5{>w��>�)]��;m�T&;]�\�A4�� �t�x�]���>}
��v=��lL��@'=G��S�S����uD����O��+��O�>��>��>o>���>��m?�5U?���>��=� ?R[`>\��<B n���?�?6$?��?�� ?��B��*���˽�M�ۿ,�,-�=D>w�X>W�=�뽿�ʽ��F<v���������{=p�3<&dμdA=$m�:̺=�+>Է�>�IܽF���Pо�=����k��>���>���7��J�e�>[%�������Z��*��W�>��>@��>��=7��='+m>�w����/�>-�K��߰=��>g��J�g>ϵ�=cmC�9���E��������޼�5>�t�>�[??�C4?�|??t���UX�tS?��W3�3mL=��r>��>.�>R�f�X�b ˾)���	/��L@�W�$xнl�=>8f�TY����>��>b���>��<�}�&�9>O�y�4>���>T�>n�'>�)�=8����ھ5�ÿd�����*�h�<]�>(�>i���(㼽�V>��c��o�k�<�?�ݭ>�>�?�Xz>��Y=�Ė�u�"E+�Z�|�jxs���8����*��Q��V��!f�zٿ�tj�����d�<�V�UY��ң�Q�*�ˏ�>���>$ �>��>q�/?�C�>���=㫁>*W?��>7W�>$𽯽�>D=�>�9?�??��=R�龱�N�E�;���=䷯=��=�9>Co>�W�=(Lt����=���=L7��X+�h�����=@|=��Q>,C�>�>�>#�+>v�=0���� ��=F���
�&�`�2!?7쯽H�Ӿ]���r >u+�{K���Q���&���z-�<�	I=bd�>a	�>�w5=H��;�h��#�������v=�� =��>YV�F�B>�Ĭ�Sܘ�ڇ����|���)�w�H��=�,�>�D?��	?��s>�	c�wU��OB�h�پ���6�<��ּ���>���ZL��\�������	��7z������L!��W9<�|Ἲ����>辛> �ż�}�=�νjS=���>2��M>?"�>*c�>��>~���D���ΰH��yVʾ����J{�=��K>j�����E��9>U+�=�C��E;���=�p[>��q>|��>yU>�ҥ>��f>k����Tz��YD��PĽ�%���?B�*����g�;UoӽS�o�5�����齥�i�ɂ�(��<��ｅ�����<���=�c�>0K�=�R߼�s(?]4<?$�1?]��>��:�ʂ>�ȑ>��?�
q��?�?E?�?��*?�|�>'��<�����Z?����=k�k=�\�=��%>٧�>����/z�=�L׼�9=�;>m�=��=h7��&K�<�r<���=H$>��>�a���8ҾBMݾ���"Up��K�>�?A�ʾ�b��ぢ=����~a�����=Ф�F����,>�T>cSd>a��<����z�=�V>h_>W�K>������������V�>��\���_E�<��XqL>o�=��=Q\%��iL?^!I?g4�>�b��j���3f��@7�Oܓ�Tr�>�4�m�>
�>#�uٯ�������q�	�󤥾=��=-��>'�G>��> K�s9�7��9�<.�=��>��)>֩m=��3=ބr>��>{��<gǽN�b����q����C��\��#�������y=���=��[�=�;���W�<�ӽ� ~��]>��۽�h�>|�n>���ʽ����2��su���-쾀���������>^�e��y���#U��Ҽ;��4��bp��ml�<!�U��ʾ�E�o
�>�˓>���>H��>�}<?��>y�F;XG��~%?-� >�W]����=g�\>�,�>���=���>�x�>���>���=���eT��
t>�V>i�E<�R�=�E>��Һ�+>`T�>�J9�����9���vu=���=��༌�ռδZ>�L�>+^#?Y ּ.ھu*����̿=|6�>�+?1=�%彋�� %�>Z�Y<�D/�e�>�����U�=�=�E�=kX�;d�=�fH�rq�S�>q��=8�ļ���f!ݻ6�=^�>�}ƽ;�)�0�=�m�K�k�_<���>>�P?=M-6?�^4?=B?k��=�%�V���J5�С+��B>Y�=��"�4M^>�]�=����������ɾ�������d`�]7�=�~?>3?=��=-m��w�<���=��]��~����ڼ�>�)�= ���W>�>��h�xP���T���¿ZǤ��F*�ۍ��Q~�=b�߼�Bq�6"=wJ$��v����>[u��iE�"'I��B�=��a>M�w>L�.>�F����>�P>괅�卟��`Ⱦ�����4���߱����������lF��tԽ��8�f�<ғ����Ĥ��J>=�>�I�>J+�>��>��?���>�_;�̂v>mg>�*�>��4�M�1>AϪ>H	?=|bf>�_?G\�=��=~�D�]����ɜ=�=��<�x>Y+�="ǟ���>>��=k캽�M=ј�=�����B���2>�n>z�/=��&>��>�a���8ҾBMݾ���"Up��K�>�?A�ʾ�b��ぢ=����~a�����=Ф�F����,>�T>cSd>a��<����z�=�V>h_>W�K>������������V�>��\���_E�<��XqL>o�=��=Q\%��iL?^!I?g4�>�b��j���3f��@7�Oܓ�Tr�>�4�m�>
�>#�uٯ�������q�	�󤥾=��=-��>'�G>��> K�s9�7��9�<.�=��>��)>֩m=��3=ބr>��>{��<gǽN�b����q����C��\��#�������y=���=��[�=�;���W�<�ӽ� ~��]>��۽�h�>|�n>���ʽ����2��su���-쾀���������>^�e��y���#U��Ҽ;��4��bp��ml�<!�U��ʾ�E�o
�>�˓>���>H��>�}<?��>y�F;XG��~%?-� >�W]����=g�\>�,�>���=���>�x�>���>���=���eT��
t>�V>i�E<�R�=�E>��Һ�+>`T�>�J9�����9���vu=���=��༌�ռδZ>�L�>+^#?Y ּ.ھu*����̿=|6�>�+?1=�%彋�� %�>Z�Y<�D/�e�>�����U�=�=�E�=kX�;d�=�fH�rq�S�>q��=8�ļ���f!ݻ6�=^�>�}ƽ;�)�0�=�m�K�k�_<���>>�P?=M-6?�^4?=B?k��=�%�V���J5�С+��B>Y�=��"�4M^>�]�=����������ɾ�������d`�]7�=�~?>3?=��=-m��w�<���=��]��~����ڼ�>�)�= ���W>�>��h�xP���T���¿ZǤ��F*�ۍ��Q~�=b�߼�Bq�6"=wJ$��v����>[u��iE�"'I��B�=��a>M�w>L�.>�F����>�P>괅�卟��`Ⱦ�����4���߱����������lF��tԽ��8�f�<ғ����Ĥ��J>=�>�I�>J+�>��>��?���>�_;�̂v>mg>�*�>��4�M�1>AϪ>H	?=|bf>�_?G\�=��=~�D�]����ɜ=�=��<�x>Y+�="ǟ���>>��=k캽�M=ј�=�����B���2>�n>z�/=��&>��>�a���8ҾBMݾ���"Up��K�>�?A�ʾ�b��ぢ=����~a�����=Ф�F����,>�T>cSd>a��<����z�=�V>h_>W�K>������������V�>��\���_E�<��XqL>o�=��=Q\%��iL?^!I?g4�>�b��j���3f��@7�Oܓ�Tr�>�4�m�>
�>#�uٯ�������q�	�󤥾=��=-��>'�G>��> K�s9�7��9�<.�=��>��)>֩m=��3=ބr>��>{��<gǽN�b����q����C��\��#�������y=���=��[�=�;���W�<�ӽ� ~��]>��۽�h�>|�n>���ʽ����2��su���-쾀���������>^�e��y���#U��Ҽ;��4��bp��ml�<!�U��ʾ�E�o
�>�˓>���>H��>�}<?��>y�F;XG��~%?-� >�W]����=g�\>�,�>���=���>�x�>���>���=���eT��
t>�V>i�E<�R�=�E>��Һ�+>`T�>�J9�����9���vu=���=��༌�ռδZ>�L�>�*�>�v��>O�?���N�G�Wa����w�4�?l�m��h�%��)�>�]3��̑�0a��E-ھ,꫾�B>/��>^��>�t�=W^n�������=�5>j��=��<�n���Y�=�Z�=��=st�������������E�S>Z�r>>=�?��??���>��+>n�� �F�ȩ ��ս�����>*�=Զ�=�ƴ���征K�����yV���2@u��1>b��"�<v��=V!e���	�;ӫ=��>�̻	�)=��&�+�=�B�>l��>I<v>�]>Z���j���eҿ����9۾���h�1�����G>�.>��A�=�P����b��\]��K�<�!|>�">X%#>��2<�� �(��������ƽ:m��%��A���0��(���RSL�D^�=5p�����>��z�u��g���ݽ�\��-8���g߽� �>&��>��
>���=�c:?��(?��?fg|��&�>���>??j���7�+\m>Ni+?��?�'?RA?M�>��3���q�w���>�^�>;�x>����x>������ɽ cA��Hh=�Ƚ<�.X>�"��]�=��x��,|=�>�B%>�/�>�j���)���ܾL�&����=�����>�="�sV]=� G�#Ƚk�˾���VYݾ��ؾ��:'>tG�>J�>���>�)�����&�=H���h�l��=������>x�>c�<����۾n����5�]��Y>��>2�=�b>y�4?�~�>���>���>��<��k4����u�V��#�JQ?�WW>�	�Hm����ξ0;��R�� ׺�
q����>��������a_@>�b=�ܼ�=>\�j>�i��Vp��0�<.1�>l��>���><N�>By��0��s���vɿ?"��9�Ծ)z��g������7�>��n=E:�������߾������=�^�>���>?�p=�ĉ�0M/>8g>Ym���T������:��wV��]ս��羋Tr��f���r;Y$�i������U��j��|
��h�8��g�>E�>���>n��>�$?��>�a�>x�=	0�>��>o�*=�sr�v�>ks�>?�?w�6?rN??@���[ ��:���U���u>�>|�=D$�=^��>&Pl��!���,=�Ԝ=�� <�i��7w��oվ;��	��C>칄>3i">�/�>�j���)���ܾL�&����=�����>�="�sV]=� G�#Ƚk�˾���VYݾ��ؾ��:'>tG�>J�>���>�)�����&�=H���h�l��=������>x�>c�<����۾n����5�]��Y>��>2�=�b>y�4?�~�>���>���>��<��k4����u�V��#�JQ?�WW>�	�Hm����ξ0;��R�� ׺�
q����>��������a_@>�b=�ܼ�=>\�j>�i��Vp��0�<.1�>l��>���><N�>By��0��s���vɿ?"��9�Ծ)z��g������7�>��n=E:�������߾������=�^�>���>?�p=�ĉ�0M/>8g>Ym���T������:��wV��]ս��羋Tr��f���r;Y$�i������U��j��|
��h�8��g�>E�>���>n��>�$?��>�a�>x�=	0�>��>o�*=�sr�v�>ks�>?�?w�6?rN??@���[ ��:���U���u>�>|�=D$�=^��>&Pl��!���,=�Ԝ=�� <�i��7w��oվ;��	��C>칄>3i">��?kcU���������%��?(��	��~�>0�<�$��</e��AҤ�͎���s��iY������7Jʼ	t�>���=K&>Y��>�g[�k�=� 8�=�,�=�X=G�X�5"">��`>2�o��Q��|�c��?�R��\B=<��=��&>��f;��v=�d/?�r�>��?d��=M�<�	�徉 T��=��xWR�"/?� ��G�E�lR������!0I���,��(���c>���ݻ�=D��=�>"R�=����c�+>��>�Ȏ�:}��a�>>�>u<�>]��>}0�>b!�=q�)���ھ0�����ҿ�������c�ȥ[���G�/Zؽ<?>���a�+��%f=V~������<��+Si=��=�9{�vOu=d�>e�?>�����!��$������s��~y*>��ـ��ܜ�"L<R!�������qm�����҈	:f0�=�m�>�A?�V�>
M?�)?�g3?�T���s�>�V>�v�`�>
��>�y*?Nc"?m�?�{�>�� �,8z�C>��&�J>&�U>'§=	Fg�g�>�3A�ms9��xY���">h��=Q��k�E�_x�����J�<�4	>!>�?Bkv���������0�ӑ2�n���1��>�c����k=�ﰾg���{d�;g���Ć�VP�g�м@	�>0!�=��S>ce>��1�&�<a��P߽�f�=�O� %T>�Ip>�L��鶎�뇯�Sd���ջ,>W2>�~�=��7�6g�=�<?�#�>.�?)�=<H�9����ﾞ	3��2F�n
�>[���J��Ly��>���^'�>�"�`��T�|=us���>>��9=���>�k=��=. >਷��P�v;���>�N�>_u�>�k�>��r�5i���a��}s	��?ֿؘ�ŀF�L��Zd�'v�=RS�O!]>@u����q��!��まp- �������=�+|��7���Ӈ�	M�=�i��*'��H4�<��G������̇⾇�.>�2���wU��Y���������&�����22O��X������j����=���>��>L9�>E�D?Dq ?E�7?����>k]Y>���>
	?Yc�>Z�?�w�>��>���>���.XQ���콧�>�Q~�=�9h=Б@=�&�=�_�=�[���Q
�b�r=�G=>�T�<v��ݡ,��5��A���ë6>�� >��=R�>�ξ5�ž_���wNm�Z	�t�D=z>4-"�@�\=p���+=�b�=�JܼSK��^��i>���>K��=1�>�k�=�佽�`
����=���<
Z�<��=��ѻ��z�=D	�=��j>���=�N.��9�������+>H�n=����RAI?s
?I�7?���ܾ���c�#�&��P=am><����I,�daU=�Hؼ�WY��S'����p���D���ԫ>]Z>�{>p�2>�>>ŝ3�����J=�Z=��=]l<�˅=M�ȼ�1>�؞�$�;-}˼xh�;�@���u:���ѽ^2����
�7&
����k�g�A�z��i<���K�,#F���R�^����-a�=g�C=~>Ss�����������{��3q�j]��� ⽂Ρ���~;�"�=�R�����O�i���Y��c"=��>��D=� M��Wz�Ckܻ���>W>N6=P�Z=j��>ǎ?���>�X�>=G�>f޽�;>z��=}]�=�o>�	>�׊>XA>	����������9�r�-DB>�n���<G�����Y>>������ruE>����=i�z�λ���g�c�j>,�>ر��A��t�>I��/��M"�C�����=ҹ�<�H�>��=�8���
���7>��>�8��w����Ͻ%.>kT�>QCv=8��>�ӟ<�*���׽�~�<ү#<G�>���1m��S���>E=\�>�Y6>X�~=fX�<]l=4Y
=�	�t_���(�7#h?
�i?}kg?�X��ۥ��)�:���C��W>͔�>euֻ.Tz�;�NJ�O�����.�1��͖���S��@�=�~�USV>]f�=�=��F��M������>ܽ9+�=Ц��}�=�I>�$9>�]v�߯����Zv=+ 俁�v��ݨ�F�<��4�������@���>���=5є�4�����ٽ�
�3R��~Y=^)<�yv>�=zt,�����K����i[��Ǥ���g���j&�=���CS��=���w����~�B�2���N����xj�c����=mK�>��F>���t>�.�>��>R��=�ᶽJ�`����9<>�>���X���,>|�>o=�>� �=!ޕ=�-F>ͫ˽J���W�>�s�=�F�P��=7G>58>���>�L>d)�QrмU�X�3> �����yU�=�!�=�Z�=�?�<t�>I��/��M"�C�����=ҹ�<�H�>��=�8���
���7>��>�8��w����Ͻ%.>kT�>QCv=8��>�ӟ<�*���׽�~�<ү#<G�>���1m��S���>E=\�>�Y6>X�~=fX�<]l=4Y
=�	�t_���(�7#h?
�i?}kg?�X��ۥ��)�:���C��W>͔�>euֻ.Tz�;�NJ�O�����.�1��͖���S��@�=�~�USV>]f�=�=��F��M������>ܽ9+�=Ц��}�=�I>�$9>�]v�߯����Zv=+ 俁�v��ݨ�F�<��4�������@���>���=5є�4�����ٽ�
�3R��~Y=^)<�yv>�=zt,�����K����i[��Ǥ���g���j&�=���CS��=���w����~�B�2���N����xj�c����=mK�>��F>���t>�.�>��>R��=�ᶽJ�`����9<>�>���X���,>|�>o=�>� �=!ޕ=�-F>ͫ˽J���W�>�s�=�F�P��=7G>58>���>�L>d)�QrмU�X�3> �����yU�=�!�=�Z�=�?�<��>�g���K������� G��^.��C
�7�?]^w����>��ͽ����1aW�����ap����< �L>�[�>�N>(ӈ>m�߽�뙽��=5פ:�UX>�>���u	[>�4���Y��<�=/C>�3��1�+���^�;��f'�>әe=�ǔ=�;?
Z@?�67?e_��|���3͹�_�V�j����]j4>-�>3��<�><~�9������W��RV��u�^��_>u�->��=�.�>�䌽���W�<����w��� >׾��F#>2�>v�>ے=؜��Q�v=��)9��ˈ����쀽5��=+mh>��s=w&���\I>����"���������(X!=��1>PM�=T�;>U[��$V���ǉ=������������Q��!�.���&>`^�����=�V��Z���u�fK'��ν7ۙ�m���Bp����p��>���>�f<=� G=��>�Z�>aw>��b�}�>������Б<���>}@�> N�>
j�='b=����<Ԥ潣���>V
�=p[��h/����>� ̽5ݣ�p�>�=��&�0c��BV�P'��_hr>;>�Ho�H�T���>�"�V#����׾&)׾U�>��#>��>\���$>�FI�����B=l�e=�A��
޽�,�:	�>(�2>M��>=��<A�⽷?�;��9<�t�=�ȼ� �H>�Ľ�3����=@�>��o=�7�=mg=B�(2ܼ0�="���}�/?�PI?* P?Z��� �%s��Z����kR�JN�=�5׻i"�>۔�=�U���տ��鶾	-��]N�䐾�ة>�q�>?Z�>�a�=� 
��zA�����>�Џ��!z=ـ	���F>޼T=��>>J�=�D�#BE��	i�vŲ�+�?�w�Ծ\�� � �ܡ��>j@>�=h6���T<�VP�iD��~��;`Z�>F��=���=��=q�>��o��I��I�н���ؾ\J��J��'����>;>\0� �X����Z�엒��ݞ�ו/��%ʽm.l�ew�)�l�sg��V�>���>���>��)?\Lx>K�F�s��I�>@����>��^�����a�>�}�>@��>D�콜��<|/���o6��]>��=��>60�<ZV2>�x>�Y����>4>�[��v7�va��]��ͽ�2�>=�>�6�=�?S8��������&�R@��d �>X?�6����T>����.z=g2ս��B>�j(>������һo���jF�$_=ں�<�[P�xC�9l >eG>v�>�i��>�Nw��^�27$�G�==pU�x|�=�zZ>�\�;-�)=�� <���=�jA?b?Wv�>�c�>Y>����O��h¾��$��=� d�>=�۽�
���Fa��*�n��{`�`�=�z@��B�=�ӂ>�o�>Eގ=5�@�
��>�'>h�"��Խ�>�{b>���=	ࣼ�ŀ;>����=�[V�Or�=`���ǌ��� ����|����MI�--ý^M����*4��������ܯ �4��>���=���=��`>%g�=��>���>��=��վ�詽���3}����ա>�n�Aޖ<R0���5@=Y�M�E���.G�L]��)$��Mt�>����>U?�|�>�\?e�?(q�>��>�'�����>�o��`$>��>�1�>o��=��=�{�>�U�=l)6�x�%�%�����P���'>�w�ɲ�<�`>�n�œ��٣�=	�!>�G>d���47<���=H�<^A�:�`�;x�>+�=7�?������O��)˾�4�;�(�=S��>�җ�h��>'k��Kؾ�5޾�޽��:�=̕1>�F�>}->?9X��f>@*	�M�/�d�w�Zu$>�֎>�>=�ך��I�=��HW�����8JI����0�[=�x>�7o�:��=�`����,>>_=?t�h?��>�垽�ﺾ�FF�򁗾!�ս��>j?&{�<��>����?'�6�/��c���c���=�:m���> :�>��E>�̋;�(�����4>��B�B�=e�=*?<x�Z>=�>r���t�ۭ�=�≾���U@��M����P��g��?�]��*�:�\j�H�?��ծ��^���oP������2�>�N�>X�.>}H=U��d�>O�>�m>�E��L��7����N;��T��,�>S�_�4��=`��7��E�t�j��9��X��hͽn����x�k�r>���>���=+w>�JZ?^e�>�"?!�`"?��h������>v9L>(��>�W�>�ן>{x�=��;�����#���ڔ�?*�=��r=�[���=�\�=8ýQ��A#ݼ���>��^=�aY<hY�=��<?)�;�O+=K_'>O�>ӓ?#σ��J���^���=`�c>]��>SC.�r�:>b}�<����#�=a*'<�ol=Ӄ��귻K�P>O��=W��=;6��_G<2���?�p>$�<9�Z=��'�iz>�N;�L�F>�ѵ�=:����=B�>W\�< ˡ=�>5<^�>�jD? iD?]`<?��>�K����*�FQԾ��<��:��b��>޼�<��7�"�����{���}2���%��u��r4���>�7>���>�y���1�� w���u>i����kZ����=��s>%0=@��=V��<)����ֽ�����<ԫڿ4슿l�1�v �ϭ|�P1�������g8��{�o��/�&�駨�Ք�>1m�=z >�}�=-���u�>�T>8L�{뾮f�㣾N�Ž�-�ɬ>��w�b4:����i�=�[�� ���	5���F��pĽ�����Y��wO>wu�>��>�e>��;?�n�>�x�>�h\� �>���5=�w�=�0>��W>�E�>���>8D�;;�'�Ae���}X��
ܽ�U�>k�W<xOn��<x=)�=-J�aH�=]�Q>v>ӕ������ͨ��1@���o=��=���<��=�?S8��������&�R@��d �>X?�6����T>����.z=g2ս��B>�j(>������һo���jF�$_=ں�<�[P�xC�9l >eG>v�>�i��>�Nw��^�27$�G�==pU�x|�=�zZ>�\�;-�)=�� <���=�jA?b?Wv�>�c�>Y>����O��h¾��$��=� d�>=�۽�
���Fa��*�n��{`�`�=�z@��B�=�ӂ>�o�>Eގ=5�@�
��>�'>h�"��Խ�>�{b>���=	ࣼ�ŀ;>����=�[V�Or�=`���ǌ��� ����|����MI�--ý^M����*4��������ܯ �4��>���=���=��`>%g�=��>���>��=��վ�詽���3}����ա>�n�Aޖ<R0���5@=Y�M�E���.G�L]��)$��Mt�>����>U?�|�>�\?e�?(q�>��>�'�����>�o��`$>��>�1�>o��=��=�{�>�U�=l)6�x�%�%�����P���'>�w�ɲ�<�`>�n�œ��٣�=	�!>�G>d���47<���=H�<^A�:�`�;x�>+�=7�?������O��)˾�4�;�(�=S��>�җ�h��>'k��Kؾ�5޾�޽��:�=̕1>�F�>}->?9X��f>@*	�M�/�d�w�Zu$>�֎>�>=�ך��I�=��HW�����8JI����0�[=�x>�7o�:��=�`����,>>_=?t�h?��>�垽�ﺾ�FF�򁗾!�ս��>j?&{�<��>����?'�6�/��c���c���=�:m���> :�>��E>�̋;�(�����4>��B�B�=e�=*?<x�Z>=�>r���t�ۭ�=�≾���U@��M����P��g��?�]��*�:�\j�H�?��ծ��^���oP������2�>�N�>X�.>}H=U��d�>O�>�m>�E��L��7����N;��T��,�>S�_�4��=`��7��E�t�j��9��X��hͽn����x�k�r>���>���=+w>�JZ?^e�>�"?!�`"?��h������>v9L>(��>�W�>�ן>{x�=��;�����#���ڔ�?*�=��r=�[���=�\�=8ýQ��A#ݼ���>��^=�aY<hY�=��<?)�;�O+=K_'>O�>��>c�徵���2D���¾SC+>렢>%*?]
��Lս�v�`��>�g��x�������j=ß�>�?Õ�>^�>�R=�W1>t�=��h<X�X=k��=A^ѽ������=���=�z:�u��[P��(�ou>�Ԣ=��=�2-��
�>hx9?��0?�==?l����M[5���0����=M1.>R��>��L�;%>B����|�#ʾG�l��Z���Y@1<rc>�B��S�4>�^QŽc��=R�>.�;�U�VN���=4I�>M��>yRW<\~:��$��7�'�޿�*������Qξ����]��={�e>V`&>T�=,4V�{蕾��z/(�?t>P��>+x> '�=�}&�]�<Q�Ӿ��o��Za��4��'��c�b��ѾaZ�=k`Z�r�<��tY� gw<`x>��O�����nk����f��c=調>�W�>�k>�F�>�(?�A�>ZYk>��G���>iz�=�L��5Ͻ�C�>g��>�~?���>�U�=�oc������X�#V��7>Z�W>L��=�J>#�p>d�K�%���q�fL,>7<4��=��(��뽽�K�<�{(>��,>W�=e�H>%�3��U8�4CK�,Kо|R�Î�=�#(?dd�<F����}=	P�>=4&�E�	�Ճ��֬=8��>`d?F]>>D$>���4M>-�t���u<�q=�%�%���҈�� �=�:�>�3Ͻ���������d�=�UM>��>���=��p><?�?�D?�-#�0\#�'�;���+��Q�=�5f>'%�<����P]=�Ą�K
���:�<X���Ӿ0�%� �'�;�L>�Uн�H꽗e8>/��>�\�lc��g�D>��=�U��Ei,�>��>��>�b0�b=B�RK�����k ��=��ٙ	���˾�3�����Q�C��5��J�=�����-�K"<<ld<��m>���>lh���O��MμF�=�B�>���>�|��6�Ɛ�,�þ~���b >���=,\��7������=�jȾ�v�����8(����Ҿi���\섾���>�<�=-Y�>#��>>�?�%?�#?��9�'�>�e�>{n~> 
�U�?�+?��;?=��>K��=y}~���K�ģ��͢�]�^=�s>%�9={�=�5>�V=��_��XI��O�<(8E>5`�ki���M�ܓ=��1>4J>���=:�>�S齡�"�f� �yѾz��=�����=?�l���o%��}>�{�>!C!�mQ�����<>Xe�>"�%?�=�=�>�F�=/�=�>[�<>�E�<��r�����	����>^}�<�e�����D���x66>U��=��=��<��>�R:?x�.?�B.?iS�;.�$�p����)�9zֽ0D��k.���=��&>'����F�C�þ'U����blн!�B9�<a>��!�����՘p>���~JȽZ�ǽL,>%;=�zɽ96H��ۅ>���>b��>��Ѽ�0��m#��s"������¿�^��MӾ@��=�6>��t>p��=r�i�@ �a���:N=��>uV>RӢ�d�ݼ-{Ǽ�ڭ>(+���ս7���2;��i��ߢ���������%�=(�b�c����V��+��o>�M�X�yݳ��j���콖�I�>�>4ko>2�>߫R>��>fͼ>/U
?wM~�V��>'?U�>���\m�>�?�{'?��/>M	�=�¿��>����
�+{�����>9!=��t�=��>:>B>|S@=c�>�zD�A�ݼ�f��쏽Yɂ��Î=��?>�F>/�q>:�>�S齡�"�f� �yѾz��=�����=?�l���o%��}>�{�>!C!�mQ�����<>Xe�>"�%?�=�=�>�F�=/�=�>[�<>�E�<��r�����	����>^}�<�e�����D���x66>U��=��=��<��>�R:?x�.?�B.?iS�;.�$�p����)�9zֽ0D��k.���=��&>'����F�C�þ'U����blн!�B9�<a>��!�����՘p>���~JȽZ�ǽL,>%;=�zɽ96H��ۅ>���>b��>��Ѽ�0��m#��s"������¿�^��MӾ@��=�6>��t>p��=r�i�@ �a���:N=��>uV>RӢ�d�ݼ-{Ǽ�ڭ>(+���ս7���2;��i��ߢ���������%�=(�b�c����V��+��o>�M�X�yݳ��j���콖�I�>�>4ko>2�>߫R>��>fͼ>/U
?wM~�V��>'?U�>���\m�>�?�{'?��/>M	�=�¿��>����
�+{�����>9!=��t�=��>:>B>|S@=c�>�zD�A�ݼ�f��쏽Yɂ��Î=��?>�F>/�q>e�H>%�3��U8�4CK�,Kо|R�Î�=�#(?dd�<F����}=	P�>=4&�E�	�Ճ��֬=8��>`d?F]>>D$>���4M>-�t���u<�q=�%�%���҈�� �=�:�>�3Ͻ���������d�=�UM>��>���=��p><?�?�D?�-#�0\#�'�;���+��Q�=�5f>'%�<����P]=�Ą�K
���:�<X���Ӿ0�%� �'�;�L>�Uн�H꽗e8>/��>�\�lc��g�D>��=�U��Ei,�>��>��>�b0�b=B�RK�����k ��=��ٙ	���˾�3�����Q�C��5��J�=�����-�K"<<ld<��m>���>lh���O��MμF�=�B�>���>�|��6�Ɛ�,�þ~���b >���=,\��7������=�jȾ�v�����8(����Ҿi���\섾���>�<�=-Y�>#��>>�?�%?�#?��9�'�>�e�>{n~> 
�U�?�+?��;?=��>K��=y}~���K�ģ��͢�]�^=�s>%�9={�=�5>�V=��_��XI��O�<(8E>5`�ki���M�ܓ=��1>4J>���=
�	  �   �۠�<]b>K���r޾Лn��J���羇OM=��/OV=��S�վa/����=�$
>����� �����֪��.J?��j=u�� eU�n��M�>���>�ۮ>�:�'�v�i�@�I����<�=���>q�:>ya����~G��:��Q�>sVE?UD_?�b�?�=���s���B�׋���m��^�ȼO�?���>�c?�ZB>��=N�����ue�2$G����>[��>����G��%���[��X�$��X�>%?� >>�?�R?��
?��`?�*?<<?4T�>!���*K��/A&?x��?}��=@�Խ��T� 9�?F����>&�)?P�B�䶗>&�?��?��&?��Q?<�?��>o� ��D@���>MW�>��W�
b����_>
�J?>0<Y?�ԃ?��=>�5�j좾�թ��J�=�>��2?5#?��?t��>8��>A�����=[[�>]�e?@��?!Xo?h��=��?#T6>��>�ҋ=�N�>�}�>�?�L?Q�p?�I?���>��<�W���[���S��"�ƞ�u�;/*b=����L C�����v=�h<�N������̼|7��%g� i�����>�Su>'���	.>��¾J���{sB>�^��r��'o����8�C��=T�~>�T?�W�>�3#�'��=��>�w�>6����'?5�?�?% ^;�,b��ܾ)HO��>��B?ְ�=��k��퓿��t�#�n=w�m?�^?��Y�����ji?��P?���R(Ͼq�ཱྀȞ���Ϳ�?！>��ؾ���>�6�?�@?�_?��*�ȓz�e���N�#C|=���;\�>��˾�X��T&>q?��@>��9���8>��X�~?��8��?�Wv?"�?�˓?��E>�����cH����o7�?�Z>�Ҧ�?�Ž#����X����T���UӪ�]���v���ģ߾�u��E��|�%�''�<-�O?f?��?cs.?�n-��ds�zU�4���H{��Oξ9O���W�^`p��s�y��L�J������.w=5)�:�A�Ԍ�?ظ'?�/�W��>���������̾�nC>Br�����z�=����@=�Z=c[h�x.��9�� ?+*�>S�>.�<?˶[�G,>���1���7�����8�3>o΢>D��>2^�>Un�:�-�t��ɾL݄��	Խxv>d?�J?��n?�
���B1�C<����!�mC��צ��p?>��>��>M�S����N&���=�-Ms��H��M��hx	��}=�1?�ց>i&�>���?e�?M���z��4�x�2s2�P�s<л�>��g?���>D�>�e�������>�^?���>�t?4��v�6�Yŏ���l=Q��>���>��?��S>�Jm�y��?S��ۉ�x����=��O?�����>a�X?b�k<�q�;.>��m�*A-�\�����R=Ƕ>�w�=,�%>���a@���E4F��F?č?VD���2��$�>RF?MG�>*��>RW|?�P�>~f��D0��� ?`�`?�X?96?J�>L�K=�0�e�ؽ���[#�=���>b�X>TF<M�X=x~O���ۀ���D=[V>V�@=)ݾ��>��`��2�<��üg��=ۿ�~K���־Vi�J��H�	���W���O߅�1��E���x��a�r�?���+�.US�w�b�����hn�mS�?�P�?��|�������A�����%�>:�s��z�������8��� �"���X� ��P�i��2e�O�'?�����ǿ񰡿�:ܾ4! ?�A ?8�y?��8�"���8�� >YC�<�,����뾭����ο?�����^?���>��/��n��>᥂>�X>�Hq>����螾r1�<��?5�-?��>��r�/�ɿb����¤<���?0�@'}A?��(����ZV=0��>�	?P�?>�P1��I�����S�>�<�?���?W�M=��W���	��~e?�2<��F���ݻ��=l=�=V>=E����J>�S�>���UA��6ܽ�4>�م>at"�����^�9��<0�]>�ս=G��LՄ?�z\�1f���/��T��^T>\�T?�*�>�<�=��,?-7H��}ϿҰ\�*a?�0�?'��?��(?_ٿ��ך>�ܾÉM?�C6?:��>�e&���t����=��������A%V�|��=W��>�>v�,����	�O�;0�����=�p����ʿJ�	�	�:����>�3���@1�'$�h�R<Ԥ~��g�%�=׮�=։>��r>�[r>�y�=�>0>T?�^?|��>j�G�2k����!�7�Ⱦ��ݼ�W>��:ｘ���0�F�5�����\��n�����b�ؾ_ =�H�=�6R����p� �\�b�"�F���.?�u$>��ʾ~�M��-<�oʾ���	ڄ�⥽�.̾��1�*"n��̟?��A?���� �V�
��d�6���f�W?�Q�Ϻ�@묾���=Y�����=�$�>8��=���+!3�lS��f$?H-?�0�������f>���Og=�!?���>୙=Ӡ�>n7?^(7�:Am�Պ�>ՙ0>Κ>��>�>>�[���	ѽTF ?ˤU?A��z���4x>5;�2�~*�=�P >���9�<�F>!��������ֺ�t�Rŉ�I�Z?l��>�Q+�����'��;���_=���?�o�> sU>4�s?#H?�%��Mݾ�oH�>�$���FU?o�~?��>�^k�:�˾3%��m0?�%\?��>���vᾩ�+���
�Z�?�iu?�_.?d&@��&f����H�2?�9x?��]�f���vQ��,p�wŠ>A��>@;�>��2�\
�>F??ND7���������UG4�9k�?n�@���?��-<�x�=!�?FT�>�zU�n�˾�
���g���L~=���>H���j����V8��R.?�}?�"�>�*s�\���a��=ٕ��Z�?��?䄪��$g<����l�en�� ��<Gѫ=�
��H"�P��w�7���ƾU�
�}����ݿ�$��>Z@�U�+�>xC8�6�TϿ1���\о�Uq�0�?��>�Ƚ���� �j��Pu�׳G�x�H�����4r�>&m�=i6!�Dۆ��v�r�*�M�m� ��>��-����>�s��g��#�׾2-żT"�>��?B��>��ݨҾ�B�?����[yϿPx��j���6?9�?K��?��3?�P=�����ٜ������=??�;n?��^?)ټ,��W��6�j?�^��wU`�(�4�XHE�!U>�"3?rD�>w�-��|=�>~��>�f>"#/�/�Ŀ�ٶ�W�����?��?�o�j��>1��?�r+?vi��7���[����*��*��<A?p2>Y�����!��/=��ђ�4�
?�}0?�}��.�Z�_?'�a�N�p���-�j�ƽ�ۡ>��0��e\�<N�����Xe����@y����?N^�?g�?յ�� #�i6%?�>c����8Ǿ��<���>�(�>�)N>�H_���u>����:�i	>���?�~�?Rj?���������U>�}?��>�Ć?�U�=S�>+��<<'ݾ�sɽ�Q9>tbs�����4�>��`?���>�A`>w4�+��K�Au��)���B��I�>�-W?�]8?��>'�,��m���-��0�'��i���T����?<՚ٽ30>>��.>��>�]�x		���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�~�?#��{���4{�IR�)<4�?5�=,+?�����{>C��>�I�=1x�|a����s��	�>�S�?�{�?���>IGn?E,h�d�L�G�==s�>u�q?�7?5~:�㾐�1>�H	?��ƾ��[���k?ǘ@s�@]!b?	衿�<ӿ�֧�a�����Ǚ��ig�>T��>\�	�RlY>A}�=�e���L=H��>��>���>��>iq>�@>!�J>�o{���.�_���X�Y��5q���	�)��b1���e�~��	��A�d��^�"N����R0<���j�������=�8o?>g/?�wa?���>���c�=)2��;�5g�������Q>^&'?L=?K'*?0S�����}�d��,���:ľ����׆>��=���>��?�u?�<�l�>�B
�B)>pY��
v<�*�f��oL>�u�>� ?�� ?�C<>��>Cϴ��1��c�h��
w�̽.�?����V�J��1���9��˦���h�=Db.?|>���?пc����2H?+���z)��+���>v�0?�cW?8�>����T�<:>A����j�/`>�+ �rl���)��%Q>zl?|f> �u>�3�48���P��o��UU}>�6?�<��0�9�e�u��bH�K�ܾ�M>H��>�2L�]��▿ ���i�gmy=�$:?�`?u8��:��u����`�Q>4\>�=K�=ÛL>'�c�bǽ�G�jk1=Y	�=�b^>'?~.>���=���>w��'�N���>�@>��->�A?(�$?���+���4��l�#��v>N�>B]�>Ⱥ>�J����=[l�>�uh>�$�q���_k��
C��[>�Pn��^��Vl�Hk�=)ޝ�(��={Г=�l���A��Y=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�v�>5e�AX��t	��G�u��#=��>WGH?�l����P��=��{
?�?�O�>���W�ȿp�v�9��>�
�?F�?��m��<���@�@�>���?qY?1�i>�e۾�lZ�=s�>��@?�R?P?�>B.��s'���?ض?̭�?�J>�e�?#s?�Q�>9J���/�Dn��6��j�{=��:I0�>^�>&U��'G�m5���r��w�j�Ϟ�+b>$=���>�K��2���3�=���������o�m�>�sn>EMK>��> ?��>�>}=d}��*���f����F?�D�?��B]���|���[���L�>w��>���=��ᾟ�>�W?��?6�K?Y�N>����樿��ʿ�˾4��=�^>���>�?߻���=�O������>P�>�B��I��QMj�W�5=�j�> �-?�]�>_�I�0?��?�պ=0�?)ZD��񏿰�V�U�>k C>�1�>��?��?����.�>�����m���lt�4�C>y&�?"?�L>�h��3����A�<1��
��>���?�E?'NZ�r?��?��0?'��?��>eF������'�<���>S�?}���B��)������?��
?[.�>�����Խ��*�������$?/Cb?}^?3���7S�L���w��<_�1��.�<AL���F<t>��=|�ڽ��>z�c>'��=��Z�3U7�%�+=�o>���>k��=H�=��p4�l�N?\n��~���O>+����M�I>�n�>�1 ���y?&>h�@�۪�ʩ��� �D�w?���?M٫?�=IHL���S?6�?�1?5�?5N��N0�t���'Ծ�t����׾��>�[)?n�׽���Jr��y1��Rq��o�Ǽ�g!�M�>�>��?�?��C>XY�>p�>�)����?����[��v�]�+�\�"�̈��o��a���@ҼJ���Q;�;R�>D�����>��?)�M>�ׅ>%�>�Z<oΙ>�w)>RU9>�y�>}ax>�-;>��>CN5=��r��|R?���#a(�|x�l0���??z}c?f��>�끽�υ�����R!?`E�?>>�?b�u>�h���-�^�?� ?LN���?��D=�Lk�f�M<\ٵ����xM��0��O�>�[�%8�%�J�޷a�=�	?�D?�끼��ѾCC��"��H=m��?�!?W@,��R�?�p�!Z�?�U��ܼ�����᤾A�$��Cr��l��R������w*���%=e1?{?uw�\���{��f4k��2@��W>���>�Õ>�
�>q�@>�V��S6��\��i%�߲z���>�x?��V>2�@?�;?%H?��[?MΑ>Z�>"e��ž
?�'E=w�>��>(�6?f *?��,?I�?~t ?��_>%ѽ��߾w��v?��*?�:"?�E?=��>G�?�̽͡)�-ν��֗�~�b������W!n��d4<za>��?t���W9�w��ުi>��1?��>kv�>���#:=Ɓ�>�+?���>������s���� ��>��?Ib��=y�$>�й=�ܻ�ߞ;P�=P:ɼ$��=��� S�{�<���=ց�=�;�S�<^,D�4���<��>`�?�f�>4�>�g��Z� �ڨ�e��=Z9Y>eMS>>@>�Uپ^����'����g�ޠy>|�?ƀ�?D�f=�	�=���=]���0��������� �<̠?4A#?�PT?M��?5�=?�n#?�>z8��Q���Z�����Ұ?�!,?���>���I�ʾ�𨿠�3�ʖ?�Z?%=a����;)�y|¾Q�Խ��>�W/��,~�����D��������_��0��?}��?x�@�u�6�|�=����f����C?��>O�>��>��)���g��#�\J;>ހ�>��Q?Z�>P?	{?��[?WYT>��8��#������Z'M�i�">R�??��?7��?�y?��>��>u�)�o��~?��x�!��|򽅏��T�Z=��Z>vB�>���>�5�>���=�ʽ	����@��G�=m�`>�l�>���>q��>��x>F��<�n^?�-�>��#��x��2����y=�#h?�ڌ?D5?ʒ:=̲S������Ɓ�>�;�?��?�=W?��i�x��=�ӽ����������=s��=���>�>�Tb>g�>Q�'?dU�>``�h�&���W�~� �X�>��_?��V>�qǿ"�����b�㫾��x�W#�STa�A!ƽ^B)�N�=�0���0���ᆾG\9�Y.�����b���,���(�����>;�=:� >��
=q4�=�I���º r=o8�=e<;=z�_�贂�H�Ž����m��$��g�:(�!=B㷼M��*�s?��*?�1?�:?�ɇ>�s�>"���A>~rG�B��>�G�=Sm�<>쓾!��͖��Ъ��(�Ⱦ	�޾%�a������L`=��ܽ���=��*>��[>i�>���=:~��>�=ƀ(���J�3dZ=&�<��=&.�=�9>�V>͐w?.��s���� P�د��:?���>���=Jwƾ�_??�8>1����㹿b����~?� �?���?�"?�m��d�>z�����%l�=''���h.>���=�(�-ռ>ɯK>"|��f���$�����?�J@?j@?�����cο0I/>+�">D�>:OR�E((��m1�p[��=뽗�$? S=�8���]>�wd=1�ӾT�����+=�o>�==����*�R�F��=@���i�<׻E=C�> �4>��=@�4����=�U=!U>�t(>|gu���$0���d=}��=�n~>��h>���>��?U0?�Ud?:.�>o�m� #ϾO���=�>��=u)�>�r�=�4B>̀�>x�7?��D?%�K?>[z�=��>��>��,�c�m��n�9̧�;�<]��?�ц?и>ET<,�A�ͣ�7[>���Ľh?V1?�m?9��>,}�w�ӿ�M��ۨ0�O��/������r����S=�>Q�]����O'>��>9�>X�>��>|
N>%��<�f�=|��>��=�9�<`�[=�2E;c�=�⽉A�=�Y���4�=
�=`~=�X�<�%=p�k�'�_�,��+<<ӊ<Z�=���>W�>�*�>	�=-����,>�b����L�vl�=e]��S�A��
d�{�~�r�/�X�6���B>�X>\�������?W�Y>��@>�J�? �t?Z�>=�jX־Kj��O�e��T�o��=��>��=���;���`�P5N�:sҾD��>��>��>��l>,�&%?�!�w=4���`5��
�>�u���o�Z)�H8q��?��S���Ni���غћD?\E��ս�=�~?F�I?�ߏ?y��>SJ����ؾ�!0>eH���=��Aq�Pi����?u
'?*��>"�h�D��|�7��*� ?ޭ�e`�Kh���bP�∾����>O��^�;�fJ������V>/�Ă��pm>f�)?�V�?�|�������4]߾���=C�>z�0?��f>�g�>��>yn�(��+��-`U>�=~?YW�?	��?�q=�o<�q=H��>�^L>Z��?�?)5�?��a�?1c"��O%=��u��->�5P>s>&]�=Z��>��>q�?�oS�h�ܾ��;���d����=*��U�
>��>�T�>O�t>l�#>��>���>	� ?ظ�>�Q>t��>Y��>�L��d��\%?�P�=K̏>G�1?r�> da={���V.�<w�B�uB�&�,��f���Qӽܰ�<���vEX=7흼���>�ƿbٖ?��O>�i��s?p�����C���W>��\>��ֽά�>"D>�>���>mH�>��>X߈>\?)>\FӾo>:���d!��,C�(�R�۽ѾN|z>����
&�O��py��BI��n���g�Yj�;.��?<=�ƽ<'H�?O�����k���)�������?p[�>�6?ی����>���>�ƍ>JK��/���ȍ�0gᾉ�?���?P��>�Ƈ>p9?ۜ?�*;�MϽffd�'膿O�A���O���v������ъ����8�� s?Wg�?�AC?�╽��> �o?�V� �E�*��>t�����[8>t�>n)�������vW�13��W�>b3�?�͓?�,#?��l�mV�pz�>�.?f]�>b?��'?922?�r��>6G?�p�>~�>��m>ʋ'?O�?��?��D>�E>��;��a�1�f�z�-9�� ��¸�^�=Up=rᎺ���=d�'����"��3�=����ؽ���<��!=o�>]�<T�>+]?r��>�G�>$�8?{����6������.?�V=O܀�PH��}]���w�A�	>��i?�%�?&FY?��g>^�A��MA��l>�t�>�,&>hY>Į�>����@�Ur�=��>�>���=L�Y�S_���	��7��DН<�r>`��>�O|>����Ko'>f���z���d>FR�����&/S�ؿG���1��nv��v�>�K?��?���=K�=q���2f��!)?B^<?�iM?0�?���=�۾��9���J��!����>��<��G���, ��N�:����:\4s>$j�������rb>�8
�P�ݾ`n�o�I���羢�6=P����N=�����ԾG7}��-�=zi>}v���j!�������� �J?�jX=h���7�S��b���>��>½�>�>��s��@�c���xd�=�>�#:>9�����vEG�5����>�H?��^?�˂?.����nq�.mE�������j�ݼD?�Ȳ>�S	?��L>�:�=���w�-�h�c�J����>�o�>��VF�U��D��>�$���>�� ?�A>��?7�R?�?cc?�8-?�5?�n�>2#����¾�A&?2��?��=G�Խ��T�| 9�MF�z��>o�)?M�B����>N�?�?��&?	�Q?�?��>� ��C@����>xY�>��W��b��!�_>��J?皳>n=Y?�ԃ?��=>\�5�ꢾ�֩��U�=�>��2?�5#?F�?���>#��>࣡�u�=�G�>��b?�2�?��o?�q�=0�?�v2>��>��=�8�>��>�?�aO?��s?�J?-��>;F�<�G��0ض���p���M�R�];�K<��{=p��,Zs�b���<�۲;E>�����!����D�6u��m��;Q��>o�r><��V�.>�>þ�,����G>'�z�J�=n���<5��G�=�y>��?؜�>7���=��>�m�>�R�}�(?8�?�v?��7;c�b�5�ؾ,�F����>c�B?�i�=�gl������w�8\g='l?��\?:�Q�ҿ��B�b?�]?%h��=���þ��b�ɉ�\�O?6�
?2�G���>��~?d�q?Y��>�e�1:n�-��Db�*�j��ж=Sr�>IX�N�d��?�>i�7?�N�>&�b>%�=ku۾	�w��q��b?��?�?���?�**>|�n�Z4�i��r��@1p?�k�>���X?�.�P���ݟ�K���RᾯՒ�t���ώ��#��M�P������$�_2=��(?�bL?|�?	iZ?� �5Y��F]��Eo��P��a�r��C?�o�C��XG���e�����Lﾈ���ޠ=sW��׽=��S�?8&?[�+����>tޛ��� �f�Ҿ��3>)����q� �=4g��=�;=��}��Q@�l���@&?Nå>�q�>��;?��Y�P;�G�1��3��9��=�6><c�>��>J��>����.�4+���Ⱦ^���֝ܽ��8>��o?��H?��a?أ꽪�/�+\����a,��C᫾�ef>��c>���>����	'��5���P�ŀ�8^*��%��X��׾=�"?P�>��>��?��?�_��!��π@������<Y��>��p?�)�>�v�>C�w��$�9��>m4m?%
�>p
�>�
��!�B|�[�ѽ@�>�H�>�F�>�No>C�)��U[�����������9����=�g?!�����]��y�>yBQ?��~�#J#<��>&o�� �����n&��u	>��?٪=-�9>#�ƾ�����{�����$u8?��>��ľ�pS���4>z�|?�R?0q�;:�?i,�>����"��3��>�`?<a?s�f?"h�>����'>Y���㕽�=�K�>qx�><����G�=����侃T�><[W>�C �G�<�0��&��< e�G3J=�L�>Amۿ�BK�N�پ�F�r?
��爾骲��c�����a��(��<Xx�����'��V��7c����ָl�χ�?�=�?����d0�����9����������>��q�ۅ����"��m)����n���dd!���O��&i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >VC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾w1�<��?7�-?��>Ǝr�1�ɿc���{¤<���?0�@iuA?��(�"L쾟�`=��>!�?�r<>F�/��v�z����>2ߞ?�>�?�~A=�IW��b��;e?��:<nF�q��x��=�ݧ=' =tc	���O>�7�>us!���@��ؽ�->6C�>Y��{��[���<|�_>�sӽ�6���|�?l\L��Rh��G�h�j��>�>M�L?/��>//>�G/?�`>���̿�W�&xQ?���?a��?��2?�������>�2��{�N?�R,?ZL{>�����%�"N�=�[^�!�]>�Y��;�H��,�>޳�>��1>2�����n�
���;�R7�d�A�ƿ!�$��|�_=&�ݺ9�[��}罕���G�T�_#��1fo���轪�h=���=��Q>Il�>U%W>4Z>gW?��k?�N�>`�>�6�t���ξNx��G�����F���%��n��R�֩߾}�	���������ɾ�=����=Y7R�����8� ���b���F�(�.?y$>��ʾI�M�*,<�qʾ]������%إ��,̾[�1��n��̟?��A?������V�k��H�y���W?TM�_��1㬾���=]����=�'�>���=z�⾎3��zS��3?��?�ɾ������+>� ����=�2+?t��>�=�ٳ>��?��h��爽��>�_V>�c�>|��>�>@���L�T�/v?�3^?�|�p����>y���Ũ�*��= >(0:���5:���=B�=�Ö�eG���Bp��v=8d\?M��<�^3��t'��/	��ꍾ"�>�[�?'�?wN`>�(�?4�E?��½��E���s�l�����=�W?!HW?��>���U���;о5B	?vLZ?��4>#蹾��ʾ��Q�	�x ?'�?�
?H(A�a���;r��v
�U?�z?l�s��ې��T,����3ƺ>��?��j>Fֽ`�/?G��>�佻�~��I��1MI�lU�?���?�{�?>�g�����=��>��y>(/<}�c�v�ǽ����x����$>uļ���h� �5���<�@?��W?�W�>�:��F����=�&K�W;�?���?�X���|o=xA�q�{���}�������{0�x�;6�ھ0�A���Ծ{�
�XX���Z>�y�_>p|@\�޽٤�>)�,�u�ֿo:ȿх�i�Ӿ�몾�%?�v�>o3ҽ�ꈾZDw��È��nY�2�F����P@�>�m=�HὠL`���k�j+5��0<���>�]�˞]>�Ӻ�4�g��� =���>��>y�>S!m��O��A�?��q-ƿTs��+CB�ā#?�]�?f�?`�3?��I>�2�����̽tk'?_�t?�E?޷"�e����>��j?1���NU`���4��`E�x�T>�!3?:N�>�~-�G�|=�k>��>D>PA/���Ŀ�ɶ�E���l��?�}�?X�/��>�x�?V`+?X�R��1I����*��"��QA?(�1>(���Ė!��=��֒��
?H�0?4O��1��_?��a�$�p���-��8ǽ�d�>g;0�rR\��,���(Ve�����Ky���?#c�?i	�?���"��/%?�ү>�M��p�ƾ��<0��>e�>hN>�9c�O�v>A����:��7
>ޜ�?�b�?�3?�p���㦿�>�}?X��>)�?���=���>s��=�E��c���K >n�=`�S�?��N?6_�>���=٤>�rm2��I��/U�����B���>T_?��H?�a>ɰ�Y$4�����4ν��4��a��C6��:9���[A>,u@>J8>��B��ԾC�?Er���ؿ�i���'�14?O��>e�?����t�� ��;_?jx�>�:��,���#��	2�ș�?�D�?��?%�׾�"̼h>{�>�U�>a�Խ-���}����7>3�B?�)��A��I�o���>���?�@@ծ?�i�(d?���S��D@f�E��QV�!.�=`+<?�ʾ��>�?�=�=�`}�y���P6p���>�>�?.U�?� �>[?h?�y\���`���<XG�>�R?�'?�=�
Ѿ �U>Ĵ?��3����L?��	@�E@�`?sG���AϿ�l���⊾|茶c��=6��=G�^>�!���3>ΛQ=��;���=�n>I��>Jhm>ݾ0>���=��#>�V>�}���)�xv���8��ՋC������z�i&
��0��������ֻ��E�39��B���W:�!6��*�WKؽ��m?HI?1�L?%	?NԽ&�����஽e3���
>���>�D?w�Z?��?t�	��޾�r�m~���I���ڍ�M�>�>��>���>zQ�>�+��91>G7+>��>;Б<�ʹ=E:���e�=qǫ>��>5� ?h��>Zp<>�D>d˴��0��,�h��Aw���˽��?�h��n�J�r-����.���w�=-n.?��>����0п�䭿$-H?����-�/+,�S�>�0?V_W?X�>����T���>����j��I>]���^Hl���)��1Q>s?��f>�u>v�3�Cg8���P�+|��ur|>�56?�ⶾ�:9���u��H�ldݾ|IM>�̾>��C��i�����[��ni�5�{=jt:?�~?=���ܰ��u�C>���TR>;\>��=*_�=LM>}cc�¶ƽ�H��h.=&��=>�^>g�?�(+>�V�=�k�>�8���M�5��>o�F>�z!>rA?l%?���B���������&��n{>I��>�> ^>�K�כ�=���>Fyh>�?���㉽�i��@�,�T>�b�x�`��K��Dǒ=�̱�ph�=�Ɛ=չ�w�8�1�=�~?���(䈿��e���lD?S+?Y �=*�F<��"�E ���H��F�?r�@m�?��	�ߢV�?�?�@�?��M��=}�>
׫>�ξ�L��?��Ž9Ǣ�ɔ	�+)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿwi�>�|�`Z�������u�Ƣ#=���>�8H?U����O�`>��w
?$?0b�(�����ȿ�zv�K��>��?/��?$�m��@��s@���>3��?�fY?)ii>�f۾YZ�t��>�@?	R?3�>�9�Q�'�P�?|޶?��?[ȸ=P_�?|�L?C?�K=��#�F��Iw�yUE�
;��=+}D>8��x���Dd���䟿;�����9�j�<���.	�>��=w���7V��7����� 6�=k�>.�>�ӑ>ː�>vz�>յ�>~�>��%�p�� ��Wܾ��K?���?,���2n��N�<l��=)�^��&?�I4?�j[�|�Ͼ�ը>�\?k?�[?d�><��P>��F迿6~��K��<��K>(4�>�H�>�$���FK>��Ծ�4D�ap�>�ϗ>s����?ھ�,���S��IB�>�e!?���>�Ү=ۙ ?��#?��j>�(�>CaE��9��W�E����>֢�>�H?�~?��?�Թ��Z3�����桿��[�t;N>��x?V?sʕ>`��������kE�+BI�8���]��?�tg?`S�.?;2�?�??`�A?w)f>܇�&ؾv�����>�{-?9x���M���@�*�m����>Ŕ?�"?�{ǼZ�R�n8K�Q�d�5a��?2�~?�)?Ĳ¾�0����$�=�y�=���m���'�6=!��>��=��Ľ���=0)>J�>c�ӽ�Z����<�N>	��>knb>�_4�i��<u2?.�e��'þH������m��U>�>~;оϑ?ɤ<�(���h���+��K�K����?{w�?5��?���;@C���A?�ф?�4?�%�>�[Ѿ���X
���оңb�۬��a�b>+�?ښ6>V����՟�����〿����[��3�>J��>��?s�?L!S>�e�>ע���*��6��|	��gZ���:5��[+�K�����U���?�=$��}�t�_Ǘ>������>*�?�o>Mo>¹�>4w���>�F>��}>Fy�>��^>�4>h��=q�1;N@ӽfLR?������'�{��ͬ���0B?�qd?M3�>y_i��������r?�z�?�p�?/[v>�lh�`+�sg?�W�>���7q
?�T:=���|�<�b�����qĆ�* ����>��ֽ�:�-M���f�j
?($?����r̾��ֽ䝬���P=*4�?��&?|9'���N�W'p�a�]�	�S�z�0�tq��0���Z �8�l�ε�������I��W+��'�<�3?�Ѐ?C\�h3�7(���h�0�@�2?r>���>�G�>�[�>��A>ܽ��3��Z�G%���z�b+�>H]y?)��>H/I??�;?��P?wL?+�>/1�>na����>3�{;3��>���>�T9?�-?�-0?&b?�{+?md>=A��j����(ؾ�?ܖ?�H?�G?��?�0������r�������z��ր�~V�=^
�<�sֽ%�t���R='�S>�Z?����8������j>m}7?��>���>�!��h$����<t	�> �
?/C�>�����sr��Z��R�>w��?�	���=w�)>�/�=6|���eں`�=����7��=(��*v;�3�<���=$��=/�t�o����	�:Љ;z��<e, ?>�?=ɇ>m4�>�������/�_��=��Z>r�S>��">�0پ�Պ��x����g���}>U�?1��?��q=���=�[�=�������w��.���=�?:�"?�R?�U�?#�=?��#?^��=�����S����)�?",?~��>���ʾj憎a�3���?�\?�>a�ͮ�
7)���¾"ս(�>�V/��)~�U���D�'ׁ����Cb��y��?k��?�A�I�6�u�0����_��/�C?� �>S�>��>g�)���g�o$��+;>��>�
R?�1�>��O?q�y?&\?�V>�D7�Cv��㲘�
���#q> x=?���?<��?]�x?,��>p�>��/����#����4*�|c���J���0W=�~^>:˓>�E�>�ʧ>���=�ѽa���'>����=��h>��>>/�>�n�>luw>��<�qJ?lz�>��׾�U���˾氘���<Vr�?���?{M&?��>'���U�)�
�dF�>4�?���?=O5?B��>U�H�o�ξbi��]w�>��>���>I�	>C�<�P�=:��>ͤ�>͆
��-"�Y�6�|M5;�%�>��-?�k�=}�ſ&.p��lm�g ��h��<F���R:d�����Y���=�^�����iȧ��@X���${��$s�������|��|�>弅=���=��=�+�<yOؼ��<�N=I2�<�=w|�2(J<��6�ֻ�����G���H<��B=�u���J-�ٿ{?$�,?��?�s?��s>��F;TЁ�L0�=IK�Ԭ�>���>��>*$��H���0ؾ�ξY��q�{�!�^)����<v̂���K>p�J>�M�>Y�J�#��=M�=dm�=�U��;����D���=82�=�'�=z[3>C�=(2w?�ׁ�<띿��R������;9?c�>�!�=$����=?Ȫ*>̓����B�Rm{?[��?��?P_?��i�/%�>j&������BΉ=�����}>���=��#���>t0>M��^=���Q�yT�?�U@�a<?f���Ϳy�7>��8>)L>��R���1�f'^�qNc�r�X���!?��:��̾}=�>䫵=�߾Y�ƾ'2=�7>�c=�K�Ѯ[�n�=nw�[}:=�g=��>�F>��=e:���.�=�OL=WF�=��O>%`��AV4�(�'��4=D�=��b>�A&>P"�>��?w>)?��x?ɇ�>��B�W�\�ʾ��;>�浼�E>�7�=�^3>5޶>�6?R/??K�K?4�>��<�Ŷ>9{�>U�*��+z��8�岪��E>v�?���?���>��v;X��{���0�o' ���?��?N��>��>�U����-Y&���.�����Q5�M+=�mr��PU�#���>m�\����=�p�>���>��>Ty>��9>��N>}�>��>�6�<Mp�=�⌻��<S ��j��=�����<*wżi����t&���+�=�����;��;¨]<B��;�5>e��>��>�O?M��=����ӉJ�B�����`��!˼���8*,�p�6�c�W��3����c�V>-j�>��|ق�>h&?U��>-��>��?��?c����¾�e�� ��6B<M>m	�>�i���[T��
P��K3��Z"��H�>ۊ�>�t�>٠n>&�+���?��1e=}���5�<�>������;����p������n����g���;:��C?$�f��=�#~?|K?��?�=�>�����پ%->)���]]�<�H�,ql�t(��sH?�&?�u�>���eeE� f��`ɓ�ߧE?�.�i�Q�s����[���/�����y��>&���s�Z�'�S���"���A�ڜ�����>�}+?���?8��A՚������8���սM�>>��?h�>��>E?���YO,��5��N[=�.�?+��?L��?C��>�~�=g����4�>H3	?��?{��?�ws?�w?�\]�>���;ǋ >=���FK�=��>���=�+�=n?��
?��
?"\����	�B�� ��$^��?�<�a�=���>lp�>�r>�
�=�=g=Ae�=�\>��>��>.�d>���>[�>U���2�&>+?��=;��>{�0?�
{>:�=���6`�<|�_�c9�Z�&�!ȷ���罛Fn<�)���&=� 	���>��ȿ��?>�R> ��׋?����<�7T>�X>!���8�>�<>��q>O�>�\�>��>UN�>��*>��վ��>#`	�� �*�B���Q�XӾ��p>�˝�(�&�:��1��G��봾�f�Fj�'t��_�=��x�<��?v 
�izi�hL)�}���?�U�>�j6?ꃋ�5�E>�{�>2�>������%G���D߾�	�?w_�?��e>L�>*YV?��?"�'��-��\���t��XC��h��,c�!����������|��P^?qhx?*cB?���;�w>H\?��#�������>Bc*���7��==��>+���"7o�c�Ծ�������^JM>�*n?r�?�?k�V��x���>r?��7?<�?09�>�8T?�XU�
�?���=w�0?�]?�wP?E?���>�~���%车F	��:���������(�=�E�=JA��O���T��<5nT=I�=]�<��	<dN�=K�J>��;��	��3�Y�ĩh=�~�=L8�>�PS?���>�U�>��9?c:�CB?�߸���y? ��#��Cg����I�徂�>�e?�|�?R#]?;�3>B7=���7���>-��>�5>�*{>	�>T)�!�,�v�w=���=�=;�=֡���g[����Z��4|2<o>(�?�H�> ����J>�__�]��ox�>D������D�|=�y��,��fy����>}�F?�*?�0>�`��Q�>�R���B?_	6?�U?��i?��<�����3�K�7��
!��>Y=U�1�^�[G��T^��$�>�b���7�>Zdھ�!��s�b>c��޾Bjn�|�I�c'��MI=1��tS=7���վP�Io�=~�	>����!����֪��3J?z�h=�,��@U������>c��>��>��:��pu�iQ@�Ϗ��=3y�>:�:>�U���^G��!��&�>�nE?J,_?h�?�肾��r�C�B�t����ע�^�ɼ��?M��>t?6^B>��=����2�#e�?G����>jb�>��]�G�Kƞ�����$�8p�>7]?��>�?.�R?j�
?��`?x.*?k?$^�>s~��]"��wA&?>��?��=j�Խ��T�H 9�F���>�)?a�B����>�?�?�&?��Q?X�?��>� ��C@�蓕>�X�>o�W�fb����_>*�J?Q��>z=Y?�ԃ?�=>�5��颾�֩��S�=`>l�2?6#?0�?]��>&?���k|x���>:�P?�?V�X?�_j=��>���<B�>�M]>��<C��>?�"J?'!�?!�\?�d	?E�w���Y�ɫ(=[�J=��� "���=�yo='29��k��-=b�=�"<��d����� 㽖�ƽY�=�8�(_�>��s>�
����0>��ľ Q��?�@>�n���O���ۊ�g�:�a�=k��>��?d��>5W#�=��=ʭ�>BH�>'��s5(?w�?]?��";��b� �ھ�K��>IB?r��=��l����A�u�Ih=��m?ʊ^?^�W��#��o�b?��]?(h�U=�|�þ��b�r�龓�O?v�
?��G�}�>��~?��q?��>�f��?n�����Fb�H�j�͟�=�y�>�U��d��6�>ŗ7?�L�>��b>��=�y۾p�w�q�� ?��?A �?��?O*>��n��3�u�$�9��s�h?,5�>�ww�d�?�6 �ԕ�3}���vվΥ��ξ����[1j��^����]�O��'�����=�&?�X�?
B�?Yok?�D�rX\��Y�u�m���b�=�e#��6A���C�81R�T�b�h�b��þ�������~6�h��?4#?s����>������sؾ��=t���7�4��=�1���d�<:�i<^���X�|����:#?���>��>�w5?��W��$B�h�/�I-��m�R>_�>G��>y�>�����(��>�OI澪&��s�I��*H>��z?�M%?��s?<ּfy-��ֈ��4+�۽��F��>6n>%Ļ>j�Ǜ@�dGK�dCY�ʆ���C�$�� ���R�=�G?k��>��>~?h�>��y��^|��𿾰��r�=\�>Wq?�$?T��>[勻�����>5l?h2�>S��>X��:� �ҳz�-�̽���>W�>�9�>�r>[H&�Q�Z�|���>����y8�ـ�=�h? ���2[����>��P?��;&��;[�>s���U!�V����)��>��?N�=�v5>��ʾ\��2~|�!:��b.?��?�ﲾl�+�[�}>56?���>���>>��?�>
h��ȧA=a��>��U?!EF?S�C?&`?6�=�Q��t߽|���M=9'�>��P>s=]�=��:�Kd�I�G�y=ݻ'>�����e���G�����-=�;�c>�oۿ�K�VDؾ���b���	�����E+���Ǉ�h
��;���|��1�w�I;��4(���V��Ed��ˌ�e�l�]n�?�m�?���7������ ������Lj�>��q�p~�����n���0�����m����`!�l1P��Qi���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�A?|�'����q�V=�&�>A	?�;C>Y�.�|~�e���?{�>�I�?���?�<=DEW��-���e?�S<�WD�
��.X�=��=Q$=��#�C>�t�>�V�D���Ͻ��0>�E�>F����b�=#w<U�V>'�h]���M�?8Lj���g�q�W�8����=jo?D�>.�>�h?Ͷl�z���oQ�-�T?܋ @2/�?!�??o��W��>�p̾%?e?'uF>�����M�G��<s����N�z�	VT�9f��:g>�Or=A�����[K�����=�_�����ƿ��$�G~�2i=Luںf�[��罏����U�.#��co�{u�o�h=��=��Q>�g�>!W>�>Z>BfW?�k?L�>��>�6�X{���
ξF���C�����¦��B���룾�P�ԫ߾��	�$��U����ɾ=�p��=2R�G���A� �z�b���F���.?�$>��ʾn�M��&/<UNʾʷ��

��Ѧ��M̾��1��n���?�B?t򅿴�V���ik�Gn���W?=u����Uì��h�=ڡ��/�=,#�>z�=���)!3�Q�S��Q<?Q�?1]��\@k���!>35>�p�=Pb?~��>�\!���>ޝJ?%�ܾ$�ҽ�-H>op`>��?�o?�8z>����%�_���*?��I?�G��Ӿ%e�>����𾊸0>�>E��f=�>�u�=�� ��Z���1�=&<�S�p���Y?fE�<��+��k�ϔ��ҾУ)>y��?i��>��>L��?�V7?�7�;��D�*kr�u���Q)�=��;?�'c?�'>�kO�/�����q�H ?�oD?e;�=A,�_�z-E�ۘ,���#?<#]?�>rQY�S?d�~��� �{�?xw?�Ya��{���߾y[⾢��=��?#�?[�
�J�>��Y?�*�Hj��}̿!�*��{�?<��?>��?��>"�ʽ��&=���>�`�>�ܚ��9���<ۤ�����=��?'�d������W0�5��=2P?qzu?W?6wݽo,ʾ�4> ��%O�?Xs�?g���| ;aZ�	�d������h=nF�=�x��2��O���<��&Ҿ_B�*����od;Y6`>x�@_	���>���Rh߿��ӿ�ڈ��"ɾ�b��Q	?u^�>H���aߛ��n�E2���OX�R������d�>�K>����!����{���;����J��>F��d�>0GR�c7��P����(<a�>\��>bȆ>3?��첽����?R����;ο�������u�X?�n�?�q�?�f?�j5<-Nv�߅{�a���G?�[s?�%Z?;?$��2]��g8���j?����]B`�1�4��oE�t�S>�3?�y�>Fp-�Bz=��>���>>�t/�e}Ŀ2���N����?q�?<O�T��>�f�?�u+?�'�����&����*��:K��/A?�1>Շ��'�!���<��c����
?Cd0?�������_?��a�5�p���-��ǽ%ԡ>��0�C\�KB���Q��Ze�y��My��?I^�?W�?���?�"��<%?'ݯ>+����<Ǿ�4�<@}�>��>IN>D_�\�u>� �� ;��	>��?�{�?t?*������0>N�}?$��>�?���<3 �>E�=�����;��iμNO�qe[�$�>��8?F�>�c�=e�þ�Ip�&p���t��5#�qP��Q�>��D?�5?l�=4�"�k7���GᾔcP��##�P�=��N潗�+<�e�>`>5~3=g0r������?�t�ߑؿRg��ù'��4?��>g?�����t�D��>_?Np�>�L�*��+���'�閫?BA�?��?��׾x�˼?'>��>�\�>��ԽYQ��*|����7>��B?!��C����o�2%�>���?�@�Ӯ?�h��@?����3��x:|���Pb�����=�yO?Xɾ�J�>t�?^�C=hk�����8Nz�
#�>�>�?���?f��>�Cg?W�p���W���=�aT>�#I?su&?�=��ξ��">H�?�����m��&pM?��@ۜ@�VV?ס��ehֿy���KN��ܗ��n��=H��=�2>��ٽ�^�=��7=h�8��?��U��=��>��d>�q>X(O>!a;>ѓ)>���7�!��q��g����C��� ����Z���Wv�#z��3�������@���4ý�y���Q��1&��:`�q<b��r?�W?{ч?�Y?�C�<�B=>���B
g�Ѵ���wJ��>�~7?��H?�8?���;����Z��G���{ؾ[����>X.�=�*�>v,�>�U�>�|
>�&Q>n�>���=�k����;&�ۼq�F=��>}�>�=�>a�>�C<>��>Fϴ��1��k�h��
w�l̽1�?���R�J��1���9��Ԧ���h�=Ib.?|>���?пf����2H?%���z)��+���>}�0?�cW?�>"����T�5:>9����j�2`>�+ �~l���)��%Q>vl?T�f>�1u>S�3�Db8�x�P��|��_Z|>;.6?����]S9�ٻu�X�H�\ݾ6HM>l��>b#F��o�����,�o�i��{=�u:?��?%<���尾$�u��:���BR>�<\>}=�p�=�RM>8c�j�ƽ�	H�#M.=���=ޡ^>�t?i&>x�}=-�>+���-KX��>��L>�}#>D�:?�%&?�d�p���lJ����9�)|>�D�> :�>%>��J���=~D�>�Xj>Dռ鍂��
��.H��gL>D���a�������=C̋��m�=�~=�D�:�;�T=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾVh�>�x��Z�������u�ڶ#=S��>�8H?�V����O�G>��v
?�?�^�੤���ȿ.|v����>V�?���?b�m��A���@����>9��?�gY?Roi>�g۾I`Z����>һ@?�R?�>�9�|�'���?�޶?ӯ�?+�H>Ĕ�?�us?�g�>�w�\/��/��8�����z=��A;�t�>x�>+����@F�gғ�Gz��Z�j�G����`>h�"=d�>����������=����X����f����>�oq>�bI>�b�>[� ?��>��>,�=�銽�Ҁ�9ܖ�m�K?ʳ�?���G0n� l�<���=�^�c%?H4?��[�:�Ͼ�ը>�\?F?�[?Ga�>S��7>���迿�~��l��<��K>@3�>MH�>4��)NK>`�Ծ�4D��m�>�͗> ���?ھ�,�������D�>kf!? ��>�Ӯ=#� ?��#?��j>y/�>XE��5��0�E�`��>)~�>.N?��~?� ?�����R3�J	���塿s�[�a$N>N�x?F?�ӕ>C����}��-]C�`�I��������?rkg?[?���?Y(�?w�??��A?��e>��@3ؾ�1��q݀>�!?N
�f�A��&�~���X?�?{#�>���ѽA�^O�	���� ?	q\?ku&?�_�D�`�]¾���<��'�qo���;MA�^�>=)>e�����=X>�[�=R2n���6��|`<��=_�>���=��6������(/?�P;zk�(�=4h�I5�`r�>�I>G�پrRX?�&��t_��m��� ����h�� �?��?��?�*?��c��V8?̀?0y?_t�>:Ӿ�J�"�۾񍇾/c$����0�=\�?&4d:�� ��s�������É���Ž�]���>���>G�?�� ?ZP>��>��3�'�Ț�f��]�����*6��n.����nʠ� �(�},�f�þ��{�4��>�𑽈�>�	?�h>.z>\�>�V����>w5R>��}>�ǧ>�UZ> 4>���=k�	<4�ս�JR?������'����5����0B?�jd?_%�>�Ui�����{���?M��?lq�?�%v>s�h�/+��h?�8�>+ ���t
?�E:=c���<�S����P/���/����>�.׽�:��M�kf��h
?�*?'y��0�̾�b׽b�ɾ9�=&^�?'�/?T��!�G���~��+e��4L���ֽe��~���ǩ�i�a������U���[���8���U��7?��k?��ؾ�QѾ.���
�O��d9�W]�>7J�>���>U'�>��D>���_?/���S�w�%��a��/�>��q?Ő�>f@I?!�9?~P?k�L?Q�>m��>Q����[�>��3;�*�>���>.l<?_/?-?k?�(?�mX>]R�v*����վ."?7�?Io?���>k��>a����U��y���sd�{wl���v�J6�=���<����P���ZQ=�hA>׾?*��'�8��:���c>�v5?!��>��>o!��!m��, =�m�>��	?o-�>g� ���p��[�(��>*��?��,=��*>�}�=si�(;���=E����=�Jz�c�?��><b��=�l�=�pN9��9���;D <~��<�??Z��>�>xS��i�Ώ���=��8> qJ>92#>�¾�����p����d��w>F��?��?n��=d'�=̈�=�ۚ�1ֲ�0�}I;d��<Q?A6?�Y?o��?��6?�w0?��>��ܩ��%���������?� ,?-��>����ʾ�憎=�3�o�?Y?�>a�����8)�T�¾��ԽK�>]/�1~�'��D��y������y��ՙ�?3��?A���6��|�꾘��[���C?�>�V�>�>�)�-�g�8&��";>��>�R?�:�>��R?7�u?U5^?h�]>�7�I������D�Ƽ�>*�:?�+�?��?��x?B��>j�>yH:��k龸^���=�Ya��
#���F~=0<f>{�>'��>�q�>-D�=@;ɽ�ֽ��C�zY�=X�d>���>�ϳ>�M�>���>�h<R�R?��>�5�P����n:��$R�=�/c?��t? �?wX�xmE�;q���k�#? ��?�w�?'�_?B�Z���=H�K>�頾w�X�2�?�m?[E7<w��T ��D��}�?V�R?;������v)\��Q�:s8?G/?�>#ƿ<mq��*o�LJ���sh<�����&f�Pږ�[[�g�=�ژ�
��������[�ڷ��kʓ�	s������|��,�>j�=eW�=��=��<�ü���<aDM=3z�<��=�n�O(m<J�9���ۻ1����v0�>�c<d�J=Nໄ�׾a�t?��?3�&?p�N?Ȯ>i�%>^8�|�r>f���>C�>l�m=��y�R�+�v�����S�@�۾El¾����b���}>#���W&�=t�>9�>�{���!�h�<��=�+=�*=�X�=��=#a�=��=�;�=KA=t?L!������FT����m�
?p?۳f>=�@� ak?�~>cǁ��g��o��
�y?�?V�?sc?�3�=/�[>�e��
��?-��޼�;`>�L�=>����>XK�>��a�(¤�±d=D��?P@Ç!?�d{��1ѿד0>ǖh>��=1=R��2�(���ؗ��0�37(?S�-�Ηھ���>2>v�־i������-�V>���=�3̽MC��F�=B\M�N;�=]�=jI�>�x>��=���7�=�i=��=n�A>K�O�V!����<:a=$>�>nk	>��>01?
0?�wd?���>�m��ξ������>���=Aӯ>�D�=��C>��>��7?�]D?l�K?4�>�R�=��>��>��,�Ln�����j�<1ǈ?��?v�>�[<_�@�0��L>��ǽ8?�$1?T?��>I��S��)����O�H�ȼ��K=���q����=.��H��� �uY>3��>�$�>�ϔ>B��=�b�=��>eJ�>i'�=�i;@'�=跏�(\>${�l�F=��->1��R�s���+�(~�������8 ��+S=�=uq=A�>T�>���>��>��>���=����Z>�n��AT�y'>0��pZ.�xF��xp�q�8�X�x��=>��%>5��2����?�y+>�>A��?�b?g��<CMh�W˾e���o�u��k�Q&
>��=�f��P��t�=X����z�>���>6w>CR�>�<� �2�~�������H����>cQ��Ʉ=�֦<sV�`���׼��)�p�:�
�L�1?�̍�3$�>%vS?��?ꐀ?��>��Y��|����=-�ȾYCF=��֜��q�����>�x�>Q�l> �	�Ĕ[��\FZ�t�:?�H��~�R�p��^i��}%=i����?��N�Z��?0�`���)��Y:����R�p>
�7?d�?C�Ǿ�0��b9v�8�{�����/�&?ڎ�?���>A#?��S?�]��c;�M�4��>��?:��?��?IA�>x�=���R �>�}
??�?�֏?)r?��7�!��>Pz�$�>񠢽�q�=�>EZ�=D��=��?# ?�? p���3
�ր�hD���^V�B�<Tl�=Ù>�h�>(z{>UT�=��t=��=��Q>ޤ�>(�>W)e>�4�>�2�>�����E�'?���=��>�!2?7 �>�ZV=�ު��<]L��s?��*�=���3bὝ��<������L=T`Ӽ�q�>H�ǿ!�?�1S>l��q	?O9���q.�S�S>��U>�ݽ���>��E>0�|>�>�>��>ܛ>?��>��(>��羅9>_�˾��f97�Z�D�o|��3>�Y��3�7��d	�Y��`sD�x������m�S@���nD�������?|�{���U�H	3�ВJ��&?V�>�=?񀾦B�<�
>`��>&��>���_������@����}�?���?�;c>��>B�W?�?Ԓ1�%3��uZ�&�u�k(A�+e�V�`��፿�����
�S��.�_?�x?4yA?uR�<':z>Q��?��%�Yӏ��)�>�/�)';� @<=w+�>*���`�n�Ӿ��þ�7��HF>��o?<%�?wY?/TV�̨��K�>��?h�:?<��?	?�$? J��09?�5�<���>E��>��F?��C?��>�?�<��T���ֽ���(�����\��<	''�LG�'����m<��=!�k>��g==Ճ=	�w:=���l��<3=��Y���ٽcc�=,d=>>��>E�Y?x��>�>��5?Z+����4�:9��1-?���<��~���}�m��}�쾮>��i?,�?u�\?SHp>YC��;��Z(>��>/e>h�R>���>:+V�/av=%%>V�!>k��=i�[��ƅ��\
�G��,��<��>�:�>��z>$���n%>����^�y��ge>�P�������R���G�1B2��lw����>fL?��?�	�=�J辦Q���e��n)?K�;?��L?P�?���=�ݾ.:���J�x��oP�>b޺<���r���q���;�ƃ�:d�t>�ϟ��(ƾy�r>��žP�����]�J[�	 �TI1�x���n��1���yƾ�GX��j�=%�=ߵ��=)��U��B"����A?��\=i�����5������=���>}�>�/�;�����.��S��P��=Ҙ�>�2>qv�43�4�N�����>wLE?6m_?of�?����s�|�B������3��FʼZ�?�q�>�b?gB>���=����^�d�t3G���>	��>�����G��0��_����$���>�J?/�>��?��R?��
?y`?�*?c8?���>ڸ��o���A&?J��?JՄ=�Խ#�T���8�d F����>�|)?k�B�Y��>��?t�?��&?��Q?��?��>K� ��?@�v��>�Q�>X�W�hb����_>��J?���>�?Y?փ?E>>��5�W&ߩ�K�=�>��2??4#?;�?Z��>V��>�����=Ҋ�>�c?N2�?}�o?�V�=c�?])2>K��>�ؖ=>���>�?	KO?8�s?�J?�u�>�5�<e?�����s��*Q�(�;�H<�y=�P���s����Y]�<T	�;�I���$��CR��#E�=���K�;yL�>C0t>$��901>��ľ�R���@>����m��<���f�:��=���>�?ߝ�>^j#��z�=;��>3�>]��L(? �?M	?A(;<�b���ھڐK��>��A?f��=�l�C}��l�u�p�g=3�m?*�^?�rW�'�����b?W�]?h�=���þ�b��z�X�O??�
?��G�A�>h�~?�q?��>!f��<n�?��Cb��j����=*w�>T���d�t<�>��7?I�>��b>%D�=|d۾��w��x��?��?���?���?�*> �n�n/�!�l]��v-b?%��>��^�T?U��T���zp������ώ�vʝ�vmu�I�/��!��S?*��,��F#�}$`>	�?Ì?�S�?\ i?�
�[�O�_��X����b������/�"i_�޲\�p�@�K�^�o�����h��o��
�����3�_	�?��'?�)�~��>�C��֘��c��8j>�e������ѱ=^Dr�
�=|�B=����=�<�ɾ��?�_�>���>n�4?ܰT��	F��� ��r-��~Ҿq4>fظ>�4�>���>�畼�.�o���;�����_�M�c>S�k?_�;?W_n?Н��9.�@d����뚽���p$W>�'>���>ř��(��Q-��B���o���$�󭜾,����=F�+?��>�>�>ἑ?[�?8���T��^����9�E��<���>�\?��>8�>���d���G�>	l?���>8b�>�+��W ���w�����^��>V��>J��>�Dy>f �2�Y��u��������8���=>Fi?&T���2Y�/��>�R?�c�&c2<��>�z���:�,�龲�/���=��?*�=m=>E-ž ���{��i��N)?�K?�璾J�*�W<~>%"?�}�>`'�>p/�?`'�>�rþZ�G�Q�?7�^?�AJ?tSA?zH�>�=Q����>Ƚ�&���,=���>��Z>Am=�= ���j\��s�z�D=�r�=��μ�K��y�<�u��x�J<��<`�3>*mۿAK�j�پ���O=
�����xв��b����g������Ox�Ɂ�|�&�7V�`>c�����l���?A>�?�t��=&��T������ ������>��q�������' �h0�����[���m`!�5�O�#i��e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾w1�<��?7�-?��>Ŏr�1�ɿc���z¤<���?0�@G�A?�E(�P��L.T=��>�{	?�A>��.�Q������>�Z�?�Ԋ?D	H=��W�5���?e?ն�;�F�(� ��J�=�<�=P=�4��I>Di�>����@��Խ#3>⻅>���C�T�^�1��<Q�X>8�ٽc���#�?��\���d�m�6�K5����=�7S?��>n�=2H-?.�J���Ͽ�-[�tX^?k�?���?Ώ'?�b���3�>�vؾ��J?�5?�O�>kG"� l�DS�=�������"�ܾW�Q�.��=�t�>H|>�����֢U�H5Ἰ!�=H�.�ƿh$��L���=�?��$�e�B��JĠ�R�W��K���<j��޽�Nv=��=rOO>H��>|�S>��[>9W?�~k?��>�>G/�?Έ���;U�>�]1���r�Pm���%��^���F��-߾�	�_H��-���Ǿ� =�X�=�6R�_���?� �<�b�5�F�x�.?@w$>��ʾ��M�0�-<jpʾӿ��vф�ॽ�-̾�1�"n�R͟?P�A?�����V�w��"Y�������W?�N�����鬾���=ﲱ�ϛ=%�>8��=W�� 3��~S�L2?�d?*�¾%���>&_꽍��=��-?7��>�o�<+ɭ>׫.?����	�-�>kz�=X��>��>��)>,������}�?��R?��
��*��RU�>�kž.O�\=�=���=�VJ��=���>7�<����PgŽ��ѽ͂E=Z?�ی>�r �w��XՇ����=��D>|�?<nA>�**>vSc?��n?$r=����
a�  ��T>ұ1?{�d?s� =�DR=����ʇP��H	?)�)?���>^J:�sܾj��hu�C�?k�?	G=?�,#��p�����e�!�{(?�8t?���Մ������?���V�?��?�?���>��`?ux�d����d���f4�//�?`�?w�?`i�=P�༘�=�0��>�Y�:vM���߾b�\����$���4>s}�m�l�T������#?�@N?}�>�h;�0� ����=�ٕ��Z�?}�?u���!@g<^���l�un��e~�<�Ϋ=���E"������7���ƾ��
����|㿼Υ�>>Z@�U�j*�>�C8�[6�
TϿ!���[оnSq���?N��>#�Ƚ����7�j��Pu�_�G�7�H�	���L��>=X�=!ͽ�奾��s�;�8���g�>�E����>������: ��lM >���>�{�>�w>�C'��Y��S1�?_���ൿ����C�&���E?�հ?6��?4E:?�Y�=�/�ٌ�;v콬_?Ek?_C+?/�C�W�ʽ�k�G�j?%���4�_��g3���D���S>k�3?�> .����=�B>�g�>�>�-��LĿ1߶�lz��޵�?�#�?���z�>���?�+?��������R���+��<�;2�B?��)>��¾���E�:��ܐ��V	?"r,?��7���Z?�t<�{�d�1!#������I>���J�+믾,uP��ƃ�;w��KDs�⒦?v�?z��?����Y�A?��C>�p=\(��@��>��?�
?1����xо7S|=���x!�'��>�N�?��?x&?)Ha�`昿���YsL?\+�>WC�?��]=�r?��E=22������"F>���f=�q�>�bX?��5?�"M>�4����n��Av�Wa�����UY�^p�>��)?K{?%)�>��0���yD��V4���ʾ$[�=�`���U4��pu>�M)>&f�<Ú��N3���?Mp�9�ؿ j��"p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>B�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji���?yE��ԡ���2E��b*������>��B?�°��B�>�%?��=Xp��Sw����l����>�m�?{�?,G
?a�Z?2ng��d��~<5�>SN?7\?�W">��׾��&>�:"?
Y1�i4��I�>�U?��@��@$�^?�^��]Qۿ�矿�p����&�=�s@=�� >��ٽu�>��=��y==$>k��>�Mb>p�J>�P >%� >�Q >y���C���������r�2����v&��#K/� �Ѿ�{D�:����/����ž��Ὗ����Ƥ���Y��`�{▽���=�Nc?2�-?�en?�?ȉ��@=���Jay�Q&������b>`j:?a�F?;�?@}<��n���=V�y{������W��2��>�sF>��>��>�̶>~��;�1>��>7ݢ<N�5�VAD�s9��FsK;��>ٸ�>�?�>W��>:F<>y�>�δ��1����h�?w��̽r �?������J�2���;������p�=�c.?1~>`���>п����`2H?����(�Կ+�f�>��0?{eW?��>���S�T�A>>����j�X> ) ��l���)�n+Q>,k?z�f>28u>��3��X8� �P�j���@S|>36?y�`9�Q�u���H�LݾcTM>���>X�E�$h��������~i��c{=|u:?�?�A��:ڰ�e�u�i>���OR>�'\>�s=��=�-M>��c�y�ƽ_�G���.=���= �^>G2?M�7>�2]=d��>�㛾$�J��@�>w7O>p>�6A?,�!?"�W;j���Zw���I��H>���>7�o>�!>��W�-��=�@�>=�r>�Q ��|��*�	��R��7p>TaS�1�z�^S��r,�=��C�Bh>)wz=2�4��Q�Ӳp=�~?���"䈿��e���lD?+?V��=$�F<��"�G ���H��(�?l�@ m�?`�	�ƢV��?�@�?�
��Q��=}�>�֫>ξ�L��?��Ž�Ƣ���	��(#�IS�?��?Q�/�Cʋ�>l�s6>�^%?�ӾQh�>yx��Z�������u�y�#=S��>�8H?�V����O�d>��v
?�?�^�੤���ȿ4|v����>X�?���?g�m��A���@����>:��?�gY?poi>�g۾5`Z����>ѻ@?�R?�>�9���'���?�޶?֯�?(�H>���?�s?iu�>&x�<f/�7��嘌���=�SP;*d�>8Y>����XF��Г��`��'�j����)aa>��$=I�>�4��&��v�=A����#��qf����>�)q>�	J>�V�>8� ?xF�>՗�>�g=W�������f��y�K?�?���y)n�1��<L��=��^��&?�A4?]�\��Ͼ�Ԩ>.�\?���?:�Z?�V�>����<���迿���F2�<��K>�/�>�F�>&��.MK>x�Ծ�2D��k�>깗>�����<ھK/���ࣻJ�>�i!?ߔ�>u�=� ?��#?{�j>�'�>�`E�9����E���>>��>�H?a�~?I�?�й�xY3�����桿��[��8N>��x?kT?X˕>��������E�LI�h�����?�tg?\>��?�0�?Њ??#�A?g)f>q���ؾ찭���>��!?�e���A���%�����?Md?���>�D��m�ֽ��n��n&��AL?��\?ۍ&?{��a�? ¾<��<��!��9Q�� <��O���>��>�L��^ͷ=�;>_�=K�m���5���h<�Y�=�(�>l4�=��7�N ��Ӣ1?���T_������}�7�U�f�>�mp>5�¾ѢP?t�e�����*��c0��$뽱��?&��?�:�?DHG���[�k]H?y�?@�?Q��>� ����,��J���kzb����Y>{:�>�>̛�5����<��̯��c�< �'>?t��>k�?;� ?fB>�}�>{P���}&��1��{��v�]�T����2��-����a����'�/?R�ӌ¾��w�(��>W}�7-�>�
?�Cn>�Ul>���>��>��>�M>��U>��>�-R>X?>�B>md�;�ܧ�3HR?}.��8�'��N�򿰾9�A?�d?�E�>�n��,��(��[�?@��?�M�?�Kt>}�h�	+�Q?@��>�i��8�
?E4;=���k;�<�)������x��vG	����>�tڽML:��aL��e��a
?~�?�<��r�̾%�Խ�g����u={��?�x)?��(���Q�F�o�
X�W�Q��Z���j�d���$��o�����
��I���()�K�=��*?�J�?���'}�����h�8�=�:f>S�>B��>%��>&�I>l�	��[1�F�]�'��������>��z?#4�>[�I?��;?�kP?\qL?���>],�>�Ư���>XĽ;6_�>���>ˡ9?�-?��/?C-?E+?ޟb>|���C����kؾ&?T�?�?
?
�?m؅��+½
��a�w�53z�����~�=�j�<Pֽ�Bs��T=�fT>s�?�t��H8�Y���g>�6?.��>!��>Y����*~��7=���>�_?���>�L�y)s�k]�t��>���?�|��=b�(>��=㛚�*���4��=���8�=������R��ӝ;kX�=Lb�=W�[��X�EJ��~^����<��
?�?�9>�A>l���!5Ӿ ���
>ۥ>XK�=��<>����ڀ��e��C)[���w>�'�?�'�?�<t=d
�=,�,>��k��v���'����Q�=Ⱦ?��?�AL?䯈?�fd?\y<?�>�J2�4X���{�O{־�=?#,?T��>���T�ʾ�꨿b~3���?�[?�<a�ch�L2)��[¾?Խ��>�b/�7~����FD�&1w���������?!��?6;A��6�cl�F����.����C?1��>F*�>{,�>٬)�/�g���L�:>�\�>m	R?��> �M?�}l?d�`? he>W�-�j[���Р�C,y��>�1?S�w?P�?~[}? ��>�oA>�*�H���D��=�콚a}�w[=5gD>'�>�+�>�>?t
>�~��"���mN�bS�=]a>b�>~��>R��>T�^><�O:��R?�r>3�Ӿ�=N�>�Ծ��Լ��C>�m?��S?�?R��=ע0��k��D�uc9?��?Nܞ?��??�]Y�.��=s�¼�!ľ��f�ݻ>���>>�K2>�1�J�2��?k��>�֣�gh��i���Б5?ƪu?5A1=�eֿvF���Ӽ�� ���e>�5W�Zz��	�3��>�>��L>l#�=*�4>�4޽=0��Z�wP��T����VǾ!M:�=��>�o�<գ�=�d�=�=�_7;`�����<Q����������Sd=���=�?;�B5�[K�z�=x&=3�"=]þ1~?��?�+5?(�U?NWx>��}>���=>�=#�þ��>C� >��7��)w���n�C����P��Ǿ�;�ሾL�����=��W�~>+��>��d>Ɵ>��V>�e7>g�L>��c='�ϻ��=�o�=J'�=���=z�>��
>Lrv?b
��@���"�i�x�n�!� ?��>
 >���2?)�>>���蛹����hp?��?���?��&?��M�:o�>U{����oWɼ?����(>���=Y(�_�Q>�q>8�+�8���O3/=_`�?O@�i?#ۊ�~[˿��P>�g>�n�=�U�e�:�X�g��3.���\�2�!?{s:��뾕��>�J?=�L�$`�=�B>�5>��C��GQ��E�=����S=���=�>r8>��=	½`�=�?�<]��=�=�>�(Y=@[5��*B����<���=]�0>چ%>���>dR?Y
?��[?�Ʋ>�u=�>�������7M>���=�dq>499�4>$��>&eL?NqL?B??���>V��=���>+l>��xG� ����3/> ��?_ݏ?o+�>�к<&u��E �<�<�/J����>t�&?�b�>�r>���[�߿q����*�_"�����@<��e�/�i<-���ʽK�L���">�l�>��>Fw�>w�P>��>&	Y>��>�!>V��<b�<������<�	����=���]�h;@f���i����V<��Q��@و���<=�<�9=���=��>�9>���>���=���*B/>˷��(�L���=�G���+B�Q4d�TI~��/��T6��B>�<X>�y���3��6�?@�Y>�p?>M��?�@u?~�>*"�c�վQ��+Ce��MS�yӸ=��> =��z;��Z`��M�0zҾ�D�>�,�>R��>�o>�}+�d=�ٷ�=.�޾@5��
�>��@�����	n�A򤿞3���(i�Y���|F?G����=6�|?��I?��?��>p]��L�پ�C5>�Ty�,��<����%h�����?Nb%?���>ϕ(C�t����z���'?�웽�Yk��4c�r�����WT��[?���[�L�:>����M��5��>��<��>8R?c��?j�������
���X�5�����>��r?鿼>���>N�7?��������@Ʉ=޶�?|�?y �?�8�>5��=�Π�>��?��?�ԑ?��s?�!?���>G�Y;y�>͎����={�> К=:U�=t[?�/
?u	
?������	��_�P�򾮧]�Z��<x�=���>�`�>�=t>��=ef=:U�=[/^>��>��>%�c>x��>�ƈ>�Ϭ��-
�Q�1?�= >N1�>J�6?x�z>���<����^�D=����U�;�� '�B ��~����/#<���e�<"lG�\��>�ʿ�˖?�2>���y�?��徢�3��?L> x>}�ҽr_�>��<>��p>��>W��>!�>\�>��P>Ѕ��t�>����Ӿk�������־1�[=#�f�ց;�d%� �|���x�������Z�0����L�5d7��ĥ?������(���3�'���FxN?���>�j?ى���,>}�=��?��F>���^��hV���.���Ӌ?��?(>c>��>2�W?G�?�1�L3��wZ��u��)A�e��`�%፿�����
�����_?0�x?�wA?_|�<�7z>+��?��%�2Ϗ��*�>/��&;�?.<=�+�>�(����`�@�Ӿ��þ5��GF>ʕo?R$�?�W?|UV��d�[¬>�t!?�!�>�h�? �N?p�/?�[���?���<���>=��>v�4?w�E?�e�>�=p�Z=J���?��齒�E��S�=	#�;y�[���F<N�~��,���Kh>3�<D�9�@d��E�=GC>��>$,I=к���t���@�=ܨ>S\?��>���>�7?:����=�뾾�%(?��=��������v�������O>,�l?_��?�V?q�m>aX?��?�ؽ>�%�>m,>��]>ww�>�C��B4�]N�=L�>P�>���=��A��8��&���t��?؅<�F>��>�:z>�镽�%>���IUx�\�R>>�_�W���E}W�0{I���1�zwv��f�> �M??�a�=�v�I��ήe���*?g�:?�P?�?.��= �߾ܓ<�$�J��5��>��<�(������t����8�/��� 	k>?9�����K�>�l��-���MY���I�����i��|ݽ&/��J#��Ͼ����+ >سg=��о�fN�,Ŗ�
紿b>?_�=��D��
�Q�\�Q�y>,�>���>��\�.W��6�����˹�<џ>0�=���|d	�?�N���1��>�>JSE?�S_?Nj�?r��.s�&�B�d����d��3�Ǽ��?�~�>j?�B>�ڭ==���d	�4�d��G���>��>��}�G�6���(����$�
��>Y5?�>��?�R?u�
?q�`?u*?�F?s(�> ������A&?��?i�=C�Խ!�T���8�fF����>d�)?��B���>�?��?�&?΅Q?�?��>� �`C@�Z��>Y�>$�W��b��;�_>G�J?���>�=Y?Ճ?7�=>(�5�	ꢾJة��R�=�>$�2?�5#??�?ٯ�>լ�>����u�@=@1�>Fk_?�"�?"Bk?*��=W��>gl*>���>"Ӻ=ׅ�>c[�>��?��L?y?��K?t��>�w<�ǌ�+m����'��+��|��`��<> `='��˗����'E=~f�<��˼<}E��R�lm��?�� �:kV�>��s>����B1>ķľ�?��S�@>~��u��|ي���:���=��>?ذ�>�(#����=Í�>�<�>���T)(?��?�?A0 ;��b�p�ھ%�K��>� B?A��=,�l�L{��	�u�Mh=	�m?�^?��W�����a?&o_?1���9�������j�����M?�&?s�6�f%�>*�?� s?��>��q��zp��*��b�b�лr�$��=0%�>���Kb�\�>~h7?X[�>x�d>�ܻ=�޾iht�_����~	?�1�?�3�?��?B�*>�lk�{0�y����H��^?��>�>����"?�� ���Ͼ�J��6����������B���z��S�$��ヾ�-׽���=/�?�s?D\q?��_?>� �� d�y/^����7mV��$�'#�r�E�� E�w�C���n��a�/������G=|j��Ď7��˷?kw#?�-���>0嗾e�
���'S�=�����!��S�=շz�bm=���<�'��.'a���Ѿ�'?�>O�>�=?USW�g�5��n0���-�d
��qD>���>�%�>K��>C��(�7�3y��ž��x�cpĽ��u>��g?L9D?�Ui?�ལ+.��N�����{�������I>�M0>>�>�D�t�#�L*�pv@���q����>�����{=��/?�É>N(�>�ڔ?o?���������04��NS�B�>m?�y�>�̍>������Y��>�2l?2z�>�E�>��n!��z�}cƽt�>�ޭ>���>��t>ld&�b�[�i叿'ߎ��E9��T�=~�h?6R��[SZ�M��>GBQ?t\�:�|<t�>����[$ �՘��{)���>�\?�W�=-�<>�9ƾ�K��|�r����0)?(B?���W�*���~>�#"?���>�Z�>.�?�o�>�&þ_5�%�?��^?�J?P;A? k�>r	=!j����Ƚ�>&��j-=6u�>��Z>;�m=���=&x���[�����3H=�P�=�	μ�2��U�<�]���E<��<84>�rۿ/K��HپC���c
��'���5�����}��Fr��	��+x��\��)'��V��uc�ݩ���l�dy�?{4�?�A��E���k���4���������>uq��}�侫�)�$��~�簬�1U!���O�i��e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >[C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@6�E?��'�L���l�<Q �>+�?$�6>\���g��V�����>]�?��v?r�	<jT�����m?8�=L(���a�S=>�=r�=�c"�F&�=<�>���A���	��� >��>c[�<�g�2r��M�F�x2>�bݽh�[8�?���4}g��1_������^8���D?���>��.=��K?v�F�"���f���F?h��?"u�?��%?|���EA>�lƾx�J?P�)?�M�>+�/v��25=��2����= ;�o�t��~>Y.?���>P���a���b��I_j�"܉>o�;�ƿ��$�[}��Q=~!���[�l�罹����U�n$��}eo�����h=���=��Q>Ri�>"W>4Z>�fW?��k?UP�>'�>�:�C����ξu���C������������Q��߾��	� ��	����ɾ%)=�N'�=R�~���h� ���b���F� �.?�$>��ʾ*�M��#-<�bʾy���-̄��䥽�9̾ݗ1�B n�cȟ?o�A?�򅿞�V�b�����"��~�W?�O�+��3񬾥�=:V��IZ=��>�<�=��� 3�5�S�|�2?.P?d����ޔ�l�(>�⳽��=K�*?�c�>�;��>@i'?�LH�b���<R>�4>宵>���>�6>n����Iy?7�S?���P���~�>����m�[=��>�4�m+��O>7���s��W��hτ�>ź;��^?�Y>�����
�5ه��1�;N��=?�k?�s�>���=F�c?d�d?\/�<�3��?r����o��=�H?�Wh?DN�=�
>��Vi��/?Z�?��~>
5V�N���U��꾻x�>�?L!?5,?��F���|�����W�?��u?ҵ~��˗�J��� ��'
>3s?��>�� �v�x>�9~?�����잿O-׿�������?��? @��X=�7)<J�=Q}�>qx>�<���:ݽ\!�� k��i%>�T���SR��!��q,�,�h?U�G?��>sY��J�B��=�ٕ�Z�?��?s����Wg<z��sl�9o��NJ�<%ҫ=k���J"�+����7�`�ƾg�
�ڨ��1Ϳ�Ť�>�Y@{S轇*�>,E8�x6��RϿv���Yо-Qq�h�?	��>m�Ƚd���;�j��Qu���G���H��������>�O�=��_����u��	&��r �s�>Mӛ�J��>����hξ�ť�M�N=���>���>vS}>���;��u��?=�"7ǿ&7���m�bN?�Y�?i��?�(?�Rp=@hO�t;{�l�
��n ?��m?��8?�u|=Ʒ�,��Xm?����iQ�X�+�9I6�E�m>}�*?2��>lu)�[�<�!^>?�=�=es-�����﮿#˾CV�?�?[�	�	?
��?L�"?U����������j$��m%<V~8?�9�=����b�!�*��W��qY�>i��>]'A��Z$���_?=�a��j��T�����w�>Mu}�E����E߽N�s��aj�_����N�B`�?H��?ن�?\��8$�+?nV�>%$�K}���%.>O��>4��>��<j�Z���=F�Mk0��v>���?F��?���>�y��e�����=�u?�2�>.g�?�|S=K��>��>��̾=B<�%>#�L<lC>�u�>�/i?��?�� >�n��4�\�xya�q�Y�4)�~<T�g��>��-?�-2?���>��<u���t׾.pP�}���aD��J�z�VzQ��%�<1��>���>%�?>3����q���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Oz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>B�Խ����\�����7>1�B?X��D��u�o�x�>���?
�@�ծ?ji��? ��Fـ�AKb�(��a���@>�j4?��;��>�q	?T�<�9z��\��v�e�5��>��?�+�?���>ߩk?B_�e�����8�vt>�;F?T�6?�	=<���r,>�)?�G8��$����m?��@n�@�<e?�޿����ۀ�<�̾1:B=1`����~=��D���=��+�6:���4=�Ӎ�=6I�>E�9>z�;>M�>H�>>.*>�؀����<�������:�����d�y B���'����
���g���#1��t9�Z炽�IG�=a2�p�'�Pm�=+'\?�dD?�_n?ۋ?���s�'>�ݾ���=�G�,===ɏ>��-?��I?�l ?�=5���|�Y��v��0I��;ߑ��ƽ>g�{>)^�>��>z��>x^�<��9>�F>j5>`t�<�`\�=8��Q=Y>��>���>ad�>gD<>ؐ>1ϴ��1��c�h�"
w�b̽ �?����ۻJ��1��:������i�={b.?�|>����>п$����2H?�����)�h�+�!�>p�0?�cW?z�>�����T��:>+��بj�B^>+ �e�l��)��&Q>Ol?Ĺf>�u>��3��d8�a�P��|���h|>�26?涾�H9���u�&�H��aݾ�HM>rþ>�8D��l�x������si�O�{=x:?�?\2���᰾8�u�B���JR>8\>�S=�c�=�VM>�cc�0�ƽH�a.=w��=V�^>�?�\)>�T�=wn�>zI��2JH��|�>�LE>	W'>J}>?J%?��d���׃��_1��vr>���>d�>�}>�fK�	��=u>�>��a>|��撽�-�UPA���W>�+t�'7^�h�h���=�ە�4��=X��=���d=�t�=��~?3��䈿�*]���lD?�&?�ڐ=(�E<"�# ���I��1�?j�@Om�?@	��V���?p@�?�����=�|�>z֫>�ξ�L��?�ƽ�Ǣ�;�	��(#�fR�?�
�?�/��ɋ�\l��3>�]%?l�ӾPh�>{x��Z�������u�u�#=R��>�8H?�V����O�e>��v
?�?�^�੤���ȿ5|v����>X�?���?g�m��A���@����>;��?�gY?roi>�g۾:`Z����>һ@?�R?�>�9���'���?�޶?֯�?�I>���?��s?�k�>M1x��Z/��6��薌��o=��[;�d�>ZX>����jgF� ؓ��h��t�j����"�a>U�$=f�>�D�G4��h9�=���H��f�f�^��>�-q>��I>�V�>�� ?b�>���>fw=0p���ှ������K?뻏?���b�m�� �<���=3�^�f&?
4?�^���Ͼ1�>ҵ\?��?	�Z?��>W���-��������Z�<T�K>7E�>�j�>�j���K>�Ծ.*D�a܉>�K�>vV��x�ھ����������>&n!?���>���=�� ?�K#?�Ei>��>ME�*	����D��%�>ܙ�>�v?E�~?c�?T·�f?3�g��]���N[��eM>��x?��?�Q�>�������~K�[oU��돽P�?�g?�6ٽ�d?��?͆@?��A?T�d>���Fھ�ŵ�Zр>��!?��r�A��-%��n��?~�?N��>l���ؽ����V"����?a�\?�&?�p�Pa�YH¾I�<����"� ��;fgB�d>]>T$�����=�C>i&�=�$m���6�ŎE<��=Ln�>���=z7������g/?�%�wa����n=̇l���6�3K{>�:Q>�Ǿ��L?�!�r�h�V���?���,~o��^�?���???�?�nR�֎b�{>?���?�R?:��>��ľ#Ӿ7ؾ.�s�[�����(^>���>��ͼ����o��9S��tG���]�Ղ�>�>A6�>�M?:�?�L>�>�ה�IH'�_�>��|\��0N6�Zz-����띾�!�t�	��¾��|�}��>}	��)(�>��?�6f>�kx>�>���:@�>�L>�J}>_�>ܼW>�>>�+>�g<GI���MR?���� �'�f��Ʈ���B?Lhd?s�>�xi��|�������?���?Zh�?�u>ˇh�_0+��Y?SO�> +��5�
?ʌ:=l��j�<�X��-���ㇽW��vߎ>��׽p#:���L�@f�bl
?_?pz����̾rG׽�𠾌�o=a�?�(?�)���Q��o�ɠW��R��*��h�Mz��ƿ$�frp�cߏ�[��u5���(�� $=6�*?�܈?>��6� &����j�F?� �f>u>�>�L�>=־>~�I>��	��1���]�}4'�����L�>?{?��>��J?=`9?N�P?i�L?��>!�>b%��Y��>i6.�aI�>�{�>�R8?Ū-?�-?��?4;(?�~`>�Q�?����پފ?��?�-?H��>�p?rR��������!8ɼ�\��h䒽��t=��<�Ͻ+K���s=Y�\>��?����8������j>Q	;?���>_2�>���2򀾦c:=Ǘ�>Ŝ?�މ>�����m����6G�>���?�1���'=�I5>3C�=3񲼾A�����=A�ټ<��=�,ؼ��%�x��<�F�=���=��ҼI}}�Iɻ���;%��<�?�=?��>s�>$��ǹ���T	�,@�=�>>��%>v�#>@����ӈ�ڗ��*l���d>[j�?�Ȳ?���=���=�>@��Vx��~���ҾT^'=�?�L"?q�O?	e�?Ɍ>?�.?\�>n3��ܕ��Ň��ά��?",?K��>���N�ʾ��ډ3���?7[?;a����9)��¾Z�Խͭ>�^/�61~�=��uD�������d�����?���?rA���6��v辇���1V����C?��>�S�>��>�)�u�g��%�9!;>Ƃ�>�
R?��>YF?cdn?QDb?��b>_�.��s������!I���u	>�3?�u?��?�]�?S��>t_Q>�-�������2�GSϽb�r�O^0=tS>�6�>���>]��>{K�=fu��\C��LX@����=��>>0�>s�>a}�>$Lm>t����U?
�>��	���L�=ϣ�f�
>�#����X?��A?}0*?j
;��>�w�{����m?-��?�d�?�,?�1�<vP�=9dh��ܘ���v�[��>6_�>ܬx>�
K>���=tu =6c,?� ?���ω(�tXO���
��f6?�S?�,�>�eԿ��L�"=�
��?a��6��ܾ��M� ׌� ��������.���k�@��� ���c���᾿+���Km�>��>Tv�=R&>��=�Y��E1�=��g=��=�
>(JI=Y��� �<�.�9WE�<7��C6�:��鼕���Cӽت����s?�º>5T??��a?��S>Nk�>�t>�3>`M5��>�ih>�>�����Ad��U����������]�� ��kߒ�ϛ�=�櫽Fdh=QK>�-�=�����*>좯=3��<��/��s�=B��<� b=U��=_6/>�=��N>�y?}Z���x����m����!�'?�e�>�;J>��۾���>Yy�>���E�ſ�*��\�?���?�@�?�KH?�t��T]v>�B��H#���+ɽ"�̽Cz�=J_0����F��>Ð�>ԝc�Ҳ��{6�[��?ӭ�?�U$? c��׿���=��7>�>>�R��e1�7�[�#b�Z�j�!?�:;�&�˾��>�6�=x߾[rƾ��.=�6>�d=��\�/I�=Kz���<=��j=���>��C>���= ���
�=�3J=���=��O>�����X7��7-���4=y��=��b>'y&>���>�>�M?V�f?ʹ>玽�*�]�)��N9;ӧ�=E1�=��g�s�%>z=�>f�C?\e?��$?B�">͉�=#��>��>���i�����$�V���uZ�>9��?�[�?H��>x�R�oR��H#��Y��ѽ���>��%?�?�֓>�U����8Y&���.�%���k�4��+=�mr��QU�M���Im�2�㽲�=�p�>���>��>7Ty>�9>��N>��>��>�6�<}p�=>ጻ���<� �����=�����<�vżV����u&�9�+�3�����;r��;B�]<��;��=���>�:>D��>Z��=���B/>�����L����=�G��Q+B�4d��H~�/��U6���B>�;X>�v���3��8�?��Y>:p?>c��?A@u?��>�#���վ�Q���De�0RS��Ӹ=�>= =��z;�[`���M�x|Ҿ_��>�I�>���>��]>��$��V?���=�kվ�k(��m?N�{�MB0=Fu漒�c�(m��^̤�{�p��v��]A?UlPU>�p?��A?U	�?�4�>(����ݾs9&>9�'��.������S��p��"?t?�8�>?a���TL�G���TU���:?�e��d�E���L�nӈ<�q�UE�>��V���ca��E��(��N6<�����>�a?U?�?4�������	$�`N��+	�>�I?y/�>�?2�$?�h��ȶ�H��I�=퐃?|��?�I�?���>�G�=�<��@��>r�
?G��?ˮ�?�q?�4�ql�>���;y�>v���9l�=�d>J�=��=".?A�?�	?���	��x�������g����<��=P{�>��>ˍ{>�}�=��T=�:�=O�[>O�>��>+h>��>�:�>���~u�7q.?���=C؉>�a+?��y>EG=�"��D�^�3�����E���"�X��x��d\�;�10��dd<R;�����>��ɿ,�?�]^>��r?����h���$>Ie>�UϽ��>�E>E�h>���>ٟ�>
E>���>i->����� >F��Ȉ��#;���H�'Ծ��n>b����g�}���f'�c���c���{f�B���g�I���6Ԟ?����ªD�o���aO��M?Exq>�1?�z����G=�[>�{?�e�>V��w��:e����ľ#u�?���?kGc>��>_�W?%�?�z1�C�2��Z��u�Y3A�ee��`��������
�Aÿ��_?G�x?$lA?�l�<�8z>^��?��%�ޏ���>/��;���<=�7�>t��F�`���ӾܹþY�@/F>�o?<!�?kW?NWV��������>���>Mb"?z�v?Y�?��2?�Zb=$�=?Hf>4��>-��>��3?�?1[>̡5�a��=(i*���>)�&5+���=��z�o�	������=л��ӽ��;>����b�=���<v�p<�<Q���=��K��<;ѿ=��>C]?	��>���> �7?{K��p8��⮾^�.?_�8=GQ�����1�����B>&�j?���?7Z?X�e>R�A��*B�l�>�E�>'�%>�*[>�n�>d�s2E�>�=�c>��>G�=��N��Y���	�!������<N�>�(	?P�=Cs<��Ҩ>ll���N�>-���$��+K���Y�]4��|�Lh!?�e?�"D?�n=<F��r�=��X�}z0?�?\j?T��?5�>e�0��<��\�������^�>[�=./��i�����p��JW���=�S��7v��ab>��m�߾��n��SI�f+��xO=6��
"W=���;A־V'{�D��=�>ᬿ�K� ��Z��O⪿`�I?��n=}`����U�ҹ��>��>�>�<����(�@��h����=ʰ�>��>>�Z�*�CH�q4�Y5�>fOE?mV_?5k�?���	s���B�����mc����Ǽ�?4x�>�b?�B>^��=`�������d�G�!�>ڥ�>7���G�72���+���$�d��>�8?�>�?q�R?��
?|�`?�*?�C?%�>X-�����*B&?���?���=��Խ��T���8��F����>�)?&�B�㳗>��?�?��&?��Q?�?��>�� ��C@�4��>�Z�>�W�la����_>(�J? ��>]<Y?-ԃ?*�=>�5��颾=ܩ��_�=/>~�2?�2#?�?
��>�H�>K��B�=ڒ�>]d?��?�mo?���=N��>Ɨ�=��>��<���>>�>�?@rM?uYu?M�E?�X�>���;�
ý�đ�����K8i����`=Ω=����aq�r��6�=�#8<��ǼT���`ˣ�F�����`�!��c�>e�s>����0>�ľ�D����@>�v��n��Ŋ�_�:�P~�=:��>W�?��>>0#����={��>-�>����2(?c�?�?gA;��b��ھ7�K���>�B?3��=J�l�y����u��g=�m?F�^?ՂW�&��en?�4?�9"���Y�����]�Ҫ����3?�h?�%k��}�=ZH?|C�?4��>�W���W�
煿#�S�󗕾�=�U�>e�۾p�v��kB>��>?�˖>���>�K>�{���Sn��w����B?���?���?$Ƭ?>8�>�}����B����v��m`?Ĵ�>蠾(� ?F1��H�Ӿ先�d����,پy���{�����������Ow��'ѽ-9�=
X?]kp?�o?�xX?�>��b�AZ_�5�z�h�R�L
����9�B���D�q?�n�n�u�	"��ݫ���VY=�֏���5��t�?;n5? W���>����(��Nk���3>�aq��_��z�<#ߜ�'I9<�c�=�mI���1��u��% -?Bp�>R��>�!?�\�9�7�{!@��&)��a��>�?�>�U�>Ǐ�>X��;��n��ͽ�;پ�5��O�v��7v>�xc?Y�K?��n?4p�+1�����O�!���/��c����B>�j>8��>�W����M:&�jY>�B�r�j��w��A�	�c�~={�2?t(�>E��>�O�?�?�{	�zk��%lx�5�1����<:1�>� i?#A�>�>�н1� ����>�l?YG�>0$�>�p��>!�>�{�.�˽*��>�E�>�j�>��o>�N-��h\��j������\/9�{��=j�h?*w����`�Μ�>��Q?tpp:��J<��>S�v��!����(��>>/p?��=�;>v|ž�/��w{�"I���?%j?�R��K"�
ߥ>��!?&?��>6)g?@�)>BJ�]���I?�D?7bQ?A?C��>�l[=2S����'�;:>O�}>�I>V�=�HT>�,�ʦD������l=0ed=�I;���})�<���<S����vڻ5��=/ۿ��J�Yi׾���LQ��	��b��3���g���N/��U�����y��-�Z�%��U��c�� ��n�
�?^_�?����ʇ������0������eʽ>�p�V�s�0��h��f����޾ګ��F� �1�O��ii��}e�_�'?e����ǿ����:ܾ1! ?�A ?K�y?���"���8�P� >0B�<�1��v��x�����οL�����^?M��>���.�����>䥂>S�X>�Hq>\��'鞾V<�<��?�-?���>��r�!�ɿ]����Ƥ<���?�@wA?��(�Y��o
U=��>�	?��?>��0��_�b���[9�>�'�?���?�&L=ڬW�%��ɏe?p�<J�F��+�(��=�\�={=}�Q�J>�|�>�����@��_ܽ�14>���>� ��e�K^��ܻ<w`]>�Nս(Ô�"Մ?z\��f�m�/�yT��=U>��T?g-�>�*�=�,?�6H�%}Ͽ7�\��)a?40�?���?0�(?�ٿ��֚>��ܾK�M?%E6?~��>�d&���t����=�=�׳������%V�.��=)��>�>`�,���7�O�d9�����=���C���/���
�0=Z��;%���p4���ڽ坍�����I�:�"B��2�<3��=[�=>��t>r�>��0>��[?���?|"�>��?>��e�PF��(��͈�<;{��rｆ������K�ƾ�uо	+޾���! �u>��Hξ:�<���=0bR������ ��Db��HF���.?h%>0�ʾxN�
�<n�Ⱦ�G����r��֣��̾|2�Tn�ޓ�?p�A?�օ���V�=��T������҈W?ߋ�z�~7��.3�=>�����=!E�>٩=���3�8bS�v1?� ?�Lؾ���N�>ܯ���a�<��<?�<�>C�>⼘>�I?,���g��E�V><�m>�f�>y��>#�5=�軾����
�6?_uf?����2���ұ>�pپ�T8��6�=���=�)��, �=3H>>;ԕ��~�>=���>��=' `?��ƽݨ/�A<徦X,��]"���̾P��?til?K��>^s�?F��?􀶾ի���>��vq��1>��r?"�?�)>�<]�޾#��b�?��V?��>!������B~3��ص���S?١6>%�����6���}��?��v?�r^�zs�����:�V�a=�>�[�>��>��9��k�>
�>?#��G��󺿿hY4�!Þ?�@x��?>�;<� ����=�;?�\�>#�O��>ƾOz��������q=�"�>�aev�����Q,�Q�8?̠�?���>�������y]�=�ؕ�uZ�?M�?:x���Rg<A���l��d��^'�<`�=��	�"�s��!�7�~�ƾ�
������}�����>V@�w���>_8�=1�PϿ�	��cSоNGq���?c|�>i�Ƚ霣��j�Ju���G�y�H�����ꝣ>��>"˖�N^��.�{��N;�p��6��>���3�>]tT�x������.<���>.\�>h�>#����ۨ�?�.��Kοj�������X?�D�?�m�?s?EN/<�w�/�{��p�:kG?��s?.dZ?��"��J^�B>�>�j?^+����`��O4��E�n�T>+�2?�p�>�-��p�=�
>�=�>3�>S�/�ĊĿBܶ�4���Φ?%��?��_��>G1�?��*?2z�&��0����e*��b9��@?�P1>������ �;�<����
�
?20?"l��l�\�_?*�a�M�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?ѵ�� #�f6%?�>c����8Ǿ��<���>�(�>*N>mH_���u>����:�
i	>���?�~�?Pj?���� ����U>	�}?l%�>S�?�`�=�[�>�i�=갾�~,��k#>���=Z�>��?�M?AT�>�D�=~�8��/�-RF��DR��#�-�C�9�>~�a?�L?�Pb>.����1��!�jNͽ`h1�Q��rN@�-w,���߽�-5>O�=>�>��D��ӾK�?���}ؿuL����(���3?�>�A?�d��Kt��:�Ś_?
և>4��m%���:�����ӡ�?�D�?P�?<ؾ>`ʼ>��>e�>�kֽj��v���z8>[�B?O��
1����o�7K�>ٸ�?��@�ή?,�h��	?���P��Va~����7�b��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?ZQo���i�B>��?"������L��f?�
@u@a�^?*�Ͽjv���,���>�*1�<���<[G>8�m��pQ=���=i�<������=���>�@b>^�.>���<_8>!A>�B���$$������e�"�P�Q���:��[���)$5�|!����˾�B������������4���m�A3�=�$V?+S?y�e?@[? ��V>uP��eN=`?�o	5=��b>�z2?� K?�y-?ն�=*pb�rn~�!��� �z�<�>��Z>��>O�>/F�>uʖ�L<->��O>2�>�0>Dq=4	�<m@�;B\=>��>��>��>��a>��>^8���U���e��qJ�JZѽ��?MD����D�<���q�� ��մ�=1�2?x0>�ލ��RԿ�έ�9>?V}��ի�LK3�ϒ>�0?�gG?��5>�տ��w��p�%>>�ޡ��5	�=�ٽ�0'�b�$�D<>�*?C�>|�>��=��F�mD��,��)�_>�|C?�~��� ��kh��~L���Ͼ�2>X �>
�=���+���U��ܖx�Oӣ=SC?5g?��׽򴾩y:�����̞$>�X�>Sg=��=�c>�O��뽖�j�-׾=JY>��}>��?2��>�̂;��p>7`��h��N�>J�j>�(C��M?�[?�i��d�=Z��:�#��>K?b�J>��k=���1R>�@?櫊>R�<���;�_U;딣�-٠>�>ڽ���&ZL=��'>A���(��=� �;�T�$�O�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>�-�aj��8܆���u���"=�.�>`�G?_W��D�F�`�>��O
?�T?Vj��ڪ����ȿ�v����>i�?d��?Іm����Q@�:�>1 �?V1Y?f�j>��پnT[��Y�>��@?�vR?i�>���{'���?�?��?�J>1P�?L�r?t��>��t�d�.��j���)�w=̆�;�a�>O�>�����G��ԓ�Ut����j����Ye>$=�
�>�U�Qϼ���=�B��A���~Vg��t�>��o>^?H>}֝>ߺ ?<��> ��>v�=]������^���;7V?�G?� :��P���C���M>�䉾j�?�^?�ֽ�����>;�Q?C�\?��^?���>J��6D������6����c:=��=J��>�}
?p�ZT=�6N��� ��>��?`��.��M���A���>? ?��?���=�.?k�>Ԋ_�EX>{8i��Ǚ�T5V�MP�>�>��?��~?7�C?�T��A�Q'��F���a}�P��>L�?�I?DZ�;�0������Q�� ������Ƣ?� �?.�m���(?˹�?ֶD?Szn?�2�>8�ž��m=�u>���=��'?@���J�)�5�3P3�ڥ?5� ?@��>N����h��6��Sɾ�"?C c?\-?M�bx�/'ھ��<CA�<��vtH�D?�;�[H>���=:�ʼ��@=|N�=G��=g�D�^~���5<�>|�>%Y�=�Ug�v.�:?,?�C�\�����=�r�u]D��>��L>0a����^?ON=���{���l��1�T�U��?G��?�[�?����h�G+=?(�?�/?1�>/���0޾C��I�v�U;x��i��t>f!�>m�n�������{���>��U�Ľ|��:��>'�>��?Je ?mU>D.�>� ���(�L�ξ^l�V�]�����I�ݽ/�����6��d�+�B�<X漾e>l��L�>��½�ۨ>ʱ	?�qt>��l>��>U
���%}>�Mc>�7{>�ޛ>}X>��(>r��=`E�<���MR?^�����'���辪����2B?�nd?�0�>$�h��������{?���?�q�?�Gv>,yh�.++�:d?0�>(���q
?;D:=(��^^�<�F��5��;'��R%���>v[׽�:��M��ef��o
?�7?�^��J�̾F׽�A��/�<��?�?��.�߷E�𨄿bX��1�f�ֽc��Gly���9�3RT�m���$�c�Q(���9���=/�P?��t?$�K�Ri,�L`�͖���N6�Qo�>1��>w�t>+8�>�>�>Z�Pt2�[�d�XN�Տ�n��>G��?�XB>v�]?�)?�?��H?�y�>��%?+{p�E̝>�+(�c��_�>M!P? ?l�H?��!?j�5?���>}P��9�վn#��>�?��?|W ?x0�>�?�`4���L=��{��I�<"�Y�5���U�L>��>qǕ�\�
�!�=��>)�?m|�ϭ;�f�=o>��5?Ķ�>&H�>�S����L� <�
�>+�>>P>���t�`��U�>ﺅ?v?���=�>GQ�=����5<jj�=��ݼ_@�=�;ȼE�w��l�<��=1o|=�@N;�@��S�����<V%<8u�>)�?���>�B�>m@���� �M��j�=�Y>yS>h>UFپ�}���$��!�g��^y>�w�?�z�?��f=�=��=�{��-T�����K������<��?�I#?bXT?<��?m�=?vj#?��>�*�YM��j^��N��خ?�8,?�>!a���˾����0!3��>?��?	�a�ݿ�y�(�`;þ4}Խ5	>"�.�c}������C��û���|җ�W��?�ݝ?��D��6�&D�-�������d	D?��>!J�>F�>�n)�~�g��A���<>8��>�R?�#�>��O?<{?��[?jhT>��8��0��oә�dc3�z�!>k@?���?�?�y?�t�>��>��)��ྂT�����G����?W=	Z>���>C)�>�>3��=CȽx_��"�>��`�=(�b>,��>��>!�>F�w>�A�<�NH?r��>ӫž�i�����97����P��7w?��?��*?HX=P|��	D�����Y�>�#�?.��?+(?�^�	��=1���%�����d�l¶>���>���>N5�=��=9�->�9�>�ɿ>'�+1���8���w���?�H?��=Y�̿�~���#>SR`>��=�|=�h$۽F�ݾ� �����Y|&��*�a袾ց���$E��I8���վm���k�*���>��'>Ý<��=�^>���="��"�<OH��\/�=�����=��*<Ɲ�� �����a=�>�<�]�=�?���	پT�u?��G?��3?�K?4k>72>~c��Xk�>7����?!vc>ȗ���E��f�'�w���瓾�-־�#�W�+�,����J1>�U)<��>�`>>n�G<.��<U(>I�=8>έ;"�&=-��=��c==��=��
>� �=�">�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>|a>�A>��]�*RE�)�7�H�:�b9j��.?i�I������;|>��<(�Ӿe�˾fS=o�i>"z�=����b��?=�e:��&�=��=}�>l>ߌ >
�o�v��;��>^�>�>,�G-=���������m>30�>X�6>��>��?N^0?�Od?B�>��m�Ͼ�0���J�>���=^2�>!��=�mB>L��>O�7?��D?��K?���>}��=O��>��>ٖ,��m��l��ϧ�4�<[��?�Ȇ?���>��P<-�A�����d>��FŽEt?zR1? f?N֞>�\
���ݿ��	�t�V�L�
�=�3c=����/�� )�Ŝ��Z���>�>~��>�F�>B�A>a�o>4=>���>��W>iR�A��<��Q�1g(��f=��=��<�K|=������=]�3���w�<�=2�JL�=]&�=�o+<J��=;��>��>��>&��=6鳾�!/>�Җ���L�1^�=YS��)B�44d�1s~�"/��6��bB>f�W>���B'��.�?��Y>|N?>�z�?zHu?� >z��i�վ<��\�e�cS��a�=�3>��<��m;��T`���M�b\Ҿ�� ?��O>t�=En�>�Y���6�sV|�Djྪ)���?�?��q��Ts��JL���ԭ�Π��	p���Ӽ�|?)c���>��F?��C?�מ?#�/?�w=�,��q�H&="��XX'��ͫ��bʾ
�4?ٞ?�\�>h����J�&%̾���L��>�?I���O�2���׭0��v�Sͷ����>������о�+3�~p��������B�9�r�K�>��O?��?=8b��Y���[O���粆�dn?�g?�2�>W>?�B?t���uG�H���p�=�n?n��?�9�?_�
>m�=9��#��>>��>��?���?�l?���A��>�����'�=�#�bJ�="y>rg>y�> 0?� ?IM?����T����܆��3ve��� ;���=��>u�t>��&>�ܠ=�l�<xt�=�7>o�>�,�>�#>Z��>��e>:����-���2?�В>G��>�/'?��>Eɼ�eM��/=�Q�=���͏]�3��������k%=Q��<�{=/ޖ�i� ?�;¿ׁ�?�F>���n�?���(��]�i>J�>qv����>�1>Ď> U0>n��>�->�V>\>��ξ�P>�J
�!�5E���S�oؾ�Ao>?Қ�l++��c��z彟�V�����}+��/i�����f�=�ˀ=��?e���D+s��"+��^�0��>��>�H9?�9���%v��#>���>���>�D��򾔿P���e⾾��?�N�?:9c>��>>�W?͙? �1�3�tZ���u��&A�N	e�c�`��፿M�����
�����w�_?��x?�xA?�H�<86z>���?R�%��ԏ��'�>�/��$;��B<=y)�>U,��B�`��Ӿɹþ�:��DF>Ǖo?%�?X?"WV���P��� ?�H5?H�?���?4�5?G�D?��Ͻ#�>f�-=Q�q>��i>��4?H�/?i+?��>�f�> ��=R^�����	�����Y��#�y���&��f�ؓ��k�=�v�Q�=��Z:�80��=���;�ޫ��DZ=��>��/>H�>Z�[?�t�>./`>��:?�� �M	!����=)?Q|�Iė�K��F��V��2>�eh?��?]pP?-�@>}AC��\K�k�5>%�o>h.>�F_>ǧ�>"x��:=�0ɑ=}R>�>��=/fb��y�o��G���Y��C�>���>Ŋ>���nJ>�Ȣ���u��a>:D��3���.G�F�#g1��Jn�ݭ�>S�J?/n?��=K���k����e�Ϥ)?2#>?�O?��}?�=i�־�@;��sH��Q�'�>���<�g�����\��UK:�V��;a�p>�&��7v��ab>��m�߾��n��SI�f+��xO=6��
"W=���;A־V'{�D��=�>ᬿ�K� ��Z��O⪿`�I?��n=}`����U�ҹ��>��>�>�<����(�@��h����=ʰ�>��>>�Z�*�CH�q4�Y5�>fOE?mV_?5k�?���	s���B�����mc����Ǽ�?4x�>�b?�B>^��=`�������d�G�!�>ڥ�>7���G�72���+���$�d��>�8?�>�?q�R?��
?|�`?�*?�C?%�>X-�����*B&?���?���=��Խ��T���8��F����>�)?&�B�㳗>��?�?��&?��Q?�?��>�� ��C@�4��>�Z�>�W�la����_>(�J? ��>]<Y?-ԃ?*�=>�5��颾=ܩ��_�=/>~�2?�2#?�?
��>�H�>K��B�=ڒ�>]d?��?�mo?���=N��>Ɨ�=��>��<���>>�>�?@rM?uYu?M�E?�X�>���;�
ý�đ�����K8i����`=Ω=����aq�r��6�=�#8<��ǼT���`ˣ�F�����`�!��c�>e�s>����0>�ľ�D����@>�v��n��Ŋ�_�:�P~�=:��>W�?��>>0#����={��>-�>����2(?c�?�?gA;��b��ھ7�K���>�B?3��=J�l�y����u��g=�m?F�^?ՂW�&��en?�4?�9"���Y�����]�Ҫ����3?�h?�%k��}�=ZH?|C�?4��>�W���W�
煿#�S�󗕾�=�U�>e�۾p�v��kB>��>?�˖>���>�K>�{���Sn��w����B?���?���?$Ƭ?>8�>�}����B����v��m`?Ĵ�>蠾(� ?F1��H�Ӿ先�d����,پy���{�����������Ow��'ѽ-9�=
X?]kp?�o?�xX?�>��b�AZ_�5�z�h�R�L
����9�B���D�q?�n�n�u�	"��ݫ���VY=�֏���5��t�?;n5? W���>����(��Nk���3>�aq��_��z�<#ߜ�'I9<�c�=�mI���1��u��% -?Bp�>R��>�!?�\�9�7�{!@��&)��a��>�?�>�U�>Ǐ�>X��;��n��ͽ�;پ�5��O�v��7v>�xc?Y�K?��n?4p�+1�����O�!���/��c����B>�j>8��>�W����M:&�jY>�B�r�j��w��A�	�c�~={�2?t(�>E��>�O�?�?�{	�zk��%lx�5�1����<:1�>� i?#A�>�>�н1� ����>�l?YG�>0$�>�p��>!�>�{�.�˽*��>�E�>�j�>��o>�N-��h\��j������\/9�{��=j�h?*w����`�Μ�>��Q?tpp:��J<��>S�v��!����(��>>/p?��=�;>v|ž�/��w{�"I���?%j?�R��K"�
ߥ>��!?&?��>6)g?@�)>BJ�]���I?�D?7bQ?A?C��>�l[=2S����'�;:>O�}>�I>V�=�HT>�,�ʦD������l=0ed=�I;���})�<���<S����vڻ5��=/ۿ��J�Yi׾���LQ��	��b��3���g���N/��U�����y��-�Z�%��U��c�� ��n�
�?^_�?����ʇ������0������eʽ>�p�V�s�0��h��f����޾ګ��F� �1�O��ii��}e�_�'?e����ǿ����:ܾ1! ?�A ?K�y?���"���8�P� >0B�<�1��v��x�����οL�����^?M��>���.�����>䥂>S�X>�Hq>\��'鞾V<�<��?�-?���>��r�!�ɿ]����Ƥ<���?�@wA?��(�Y��o
U=��>�	?��?>��0��_�b���[9�>�'�?���?�&L=ڬW�%��ɏe?p�<J�F��+�(��=�\�={=}�Q�J>�|�>�����@��_ܽ�14>���>� ��e�K^��ܻ<w`]>�Nս(Ô�"Մ?z\��f�m�/�yT��=U>��T?g-�>�*�=�,?�6H�%}Ͽ7�\��)a?40�?���?0�(?�ٿ��֚>��ܾK�M?%E6?~��>�d&���t����=�=�׳������%V�.��=)��>�>`�,���7�O�d9�����=���C���/���
�0=Z��;%���p4���ڽ坍�����I�:�"B��2�<3��=[�=>��t>r�>��0>��[?���?|"�>��?>��e�PF��(��͈�<;{��rｆ������K�ƾ�uо	+޾���! �u>��Hξ:�<���=0bR������ ��Db��HF���.?h%>0�ʾxN�
�<n�Ⱦ�G����r��֣��̾|2�Tn�ޓ�?p�A?�օ���V�=��T������҈W?ߋ�z�~7��.3�=>�����=!E�>٩=���3�8bS�v1?� ?�Lؾ���N�>ܯ���a�<��<?�<�>C�>⼘>�I?,���g��E�V><�m>�f�>y��>#�5=�軾����
�6?_uf?����2���ұ>�pپ�T8��6�=���=�)��, �=3H>>;ԕ��~�>=���>��=' `?��ƽݨ/�A<徦X,��]"���̾P��?til?K��>^s�?F��?􀶾ի���>��vq��1>��r?"�?�)>�<]�޾#��b�?��V?��>!������B~3��ص���S?١6>%�����6���}��?��v?�r^�zs�����:�V�a=�>�[�>��>��9��k�>
�>?#��G��󺿿hY4�!Þ?�@x��?>�;<� ����=�;?�\�>#�O��>ƾOz��������q=�"�>�aev�����Q,�Q�8?̠�?���>�������y]�=�ؕ�uZ�?M�?:x���Rg<A���l��d��^'�<`�=��	�"�s��!�7�~�ƾ�
������}�����>V@�w���>_8�=1�PϿ�	��cSоNGq���?c|�>i�Ƚ霣��j�Ju���G�y�H�����ꝣ>��>"˖�N^��.�{��N;�p��6��>���3�>]tT�x������.<���>.\�>h�>#����ۨ�?�.��Kοj�������X?�D�?�m�?s?EN/<�w�/�{��p�:kG?��s?.dZ?��"��J^�B>�>�j?^+����`��O4��E�n�T>+�2?�p�>�-��p�=�
>�=�>3�>S�/�ĊĿBܶ�4���Φ?%��?��_��>G1�?��*?2z�&��0����e*��b9��@?�P1>������ �;�<����
�
?20?"l��l�\�_?*�a�M�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?ѵ�� #�f6%?�>c����8Ǿ��<���>�(�>*N>mH_���u>����:�
i	>���?�~�?Pj?���� ����U>	�}?l%�>S�?�`�=�[�>�i�=갾�~,��k#>���=Z�>��?�M?AT�>�D�=~�8��/�-RF��DR��#�-�C�9�>~�a?�L?�Pb>.����1��!�jNͽ`h1�Q��rN@�-w,���߽�-5>O�=>�>��D��ӾK�?���}ؿuL����(���3?�>�A?�d��Kt��:�Ś_?
և>4��m%���:�����ӡ�?�D�?P�?<ؾ>`ʼ>��>e�>�kֽj��v���z8>[�B?O��
1����o�7K�>ٸ�?��@�ή?,�h��	?���P��Va~����7�b��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?ZQo���i�B>��?"������L��f?�
@u@a�^?*�Ͽjv���,���>�*1�<���<[G>8�m��pQ=���=i�<������=���>�@b>^�.>���<_8>!A>�B���$$������e�"�P�Q���:��[���)$5�|!����˾�B������������4���m�A3�=�$V?+S?y�e?@[? ��V>uP��eN=`?�o	5=��b>�z2?� K?�y-?ն�=*pb�rn~�!��� �z�<�>��Z>��>O�>/F�>uʖ�L<->��O>2�>�0>Dq=4	�<m@�;B\=>��>��>��>��a>��>^8���U���e��qJ�JZѽ��?MD����D�<���q�� ��մ�=1�2?x0>�ލ��RԿ�έ�9>?V}��ի�LK3�ϒ>�0?�gG?��5>�տ��w��p�%>>�ޡ��5	�=�ٽ�0'�b�$�D<>�*?C�>|�>��=��F�mD��,��)�_>�|C?�~��� ��kh��~L���Ͼ�2>X �>
�=���+���U��ܖx�Oӣ=SC?5g?��׽򴾩y:�����̞$>�X�>Sg=��=�c>�O��뽖�j�-׾=JY>��}>��?2��>�̂;��p>7`��h��N�>J�j>�(C��M?�[?�i��d�=Z��:�#��>K?b�J>��k=���1R>�@?櫊>R�<���;�_U;딣�-٠>�>ڽ���&ZL=��'>A���(��=� �;�T�$�O�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>�-�aj��8܆���u���"=�.�>`�G?_W��D�F�`�>��O
?�T?Vj��ڪ����ȿ�v����>i�?d��?Іm����Q@�:�>1 �?V1Y?f�j>��پnT[��Y�>��@?�vR?i�>���{'���?�?��?�J>1P�?L�r?t��>��t�d�.��j���)�w=̆�;�a�>O�>�����G��ԓ�Ut����j����Ye>$=�
�>�U�Qϼ���=�B��A���~Vg��t�>��o>^?H>}֝>ߺ ?<��> ��>v�=]������^���;7V?�G?� :��P���C���M>�䉾j�?�^?�ֽ�����>;�Q?C�\?��^?���>J��6D������6����c:=��=J��>�}
?p�ZT=�6N��� ��>��?`��.��M���A���>? ?��?���=�.?k�>Ԋ_�EX>{8i��Ǚ�T5V�MP�>�>��?��~?7�C?�T��A�Q'��F���a}�P��>L�?�I?DZ�;�0������Q�� ������Ƣ?� �?.�m���(?˹�?ֶD?Szn?�2�>8�ž��m=�u>���=��'?@���J�)�5�3P3�ڥ?5� ?@��>N����h��6��Sɾ�"?C c?\-?M�bx�/'ھ��<CA�<��vtH�D?�;�[H>���=:�ʼ��@=|N�=G��=g�D�^~���5<�>|�>%Y�=�Ug�v.�:?,?�C�\�����=�r�u]D��>��L>0a����^?ON=���{���l��1�T�U��?G��?�[�?����h�G+=?(�?�/?1�>/���0޾C��I�v�U;x��i��t>f!�>m�n�������{���>��U�Ľ|��:��>'�>��?Je ?mU>D.�>� ���(�L�ξ^l�V�]�����I�ݽ/�����6��d�+�B�<X漾e>l��L�>��½�ۨ>ʱ	?�qt>��l>��>U
���%}>�Mc>�7{>�ޛ>}X>��(>r��=`E�<���MR?^�����'���辪����2B?�nd?�0�>$�h��������{?���?�q�?�Gv>,yh�.++�:d?0�>(���q
?;D:=(��^^�<�F��5��;'��R%���>v[׽�:��M��ef��o
?�7?�^��J�̾F׽�A��/�<��?�?��.�߷E�𨄿bX��1�f�ֽc��Gly���9�3RT�m���$�c�Q(���9���=/�P?��t?$�K�Ri,�L`�͖���N6�Qo�>1��>w�t>+8�>�>�>Z�Pt2�[�d�XN�Տ�n��>G��?�XB>v�]?�)?�?��H?�y�>��%?+{p�E̝>�+(�c��_�>M!P? ?l�H?��!?j�5?���>}P��9�վn#��>�?��?|W ?x0�>�?�`4���L=��{��I�<"�Y�5���U�L>��>qǕ�\�
�!�=��>)�?m|�ϭ;�f�=o>��5?Ķ�>&H�>�S����L� <�
�>+�>>P>���t�`��U�>ﺅ?v?���=�>GQ�=����5<jj�=��ݼ_@�=�;ȼE�w��l�<��=1o|=�@N;�@��S�����<V%<8u�>)�?���>�B�>m@���� �M��j�=�Y>yS>h>UFپ�}���$��!�g��^y>�w�?�z�?��f=�=��=�{��-T�����K������<��?�I#?bXT?<��?m�=?vj#?��>�*�YM��j^��N��خ?�8,?�>!a���˾����0!3��>?��?	�a�ݿ�y�(�`;þ4}Խ5	>"�.�c}������C��û���|җ�W��?�ݝ?��D��6�&D�-�������d	D?��>!J�>F�>�n)�~�g��A���<>8��>�R?�#�>��O?<{?��[?jhT>��8��0��oә�dc3�z�!>k@?���?�?�y?�t�>��>��)��ྂT�����G����?W=	Z>���>C)�>�>3��=CȽx_��"�>��`�=(�b>,��>��>!�>F�w>�A�<�NH?r��>ӫž�i�����97����P��7w?��?��*?HX=P|��	D�����Y�>�#�?.��?+(?�^�	��=1���%�����d�l¶>���>���>N5�=��=9�->�9�>�ɿ>'�+1���8���w���?�H?��=Y�̿�~���#>SR`>��=�|=�h$۽F�ݾ� �����Y|&��*�a袾ց���$E��I8���վm���k�*���>��'>Ý<��=�^>���="��"�<OH��\/�=�����=��*<Ɲ�� �����a=�>�<�]�=�?���	پT�u?��G?��3?�K?4k>72>~c��Xk�>7����?!vc>ȗ���E��f�'�w���瓾�-־�#�W�+�,����J1>�U)<��>�`>>n�G<.��<U(>I�=8>έ;"�&=-��=��c==��=��
>� �=�">�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>|a>�A>��]�*RE�)�7�H�:�b9j��.?i�I������;|>��<(�Ӿe�˾fS=o�i>"z�=����b��?=�e:��&�=��=}�>l>ߌ >
�o�v��;��>^�>�>,�G-=���������m>30�>X�6>��>��?N^0?�Od?B�>��m�Ͼ�0���J�>���=^2�>!��=�mB>L��>O�7?��D?��K?���>}��=O��>��>ٖ,��m��l��ϧ�4�<[��?�Ȇ?���>��P<-�A�����d>��FŽEt?zR1? f?N֞>�\
���ݿ��	�t�V�L�
�=�3c=����/�� )�Ŝ��Z���>�>~��>�F�>B�A>a�o>4=>���>��W>iR�A��<��Q�1g(��f=��=��<�K|=������=]�3���w�<�=2�JL�=]&�=�o+<J��=;��>��>��>&��=6鳾�!/>�Җ���L�1^�=YS��)B�44d�1s~�"/��6��bB>f�W>���B'��.�?��Y>|N?>�z�?zHu?� >z��i�վ<��\�e�cS��a�=�3>��<��m;��T`���M�b\Ҿ�� ?��O>t�=En�>�Y���6�sV|�Djྪ)���?�?��q��Ts��JL���ԭ�Π��	p���Ӽ�|?)c���>��F?��C?�מ?#�/?�w=�,��q�H&="��XX'��ͫ��bʾ
�4?ٞ?�\�>h����J�&%̾���L��>�?I���O�2���׭0��v�Sͷ����>������о�+3�~p��������B�9�r�K�>��O?��?=8b��Y���[O���粆�dn?�g?�2�>W>?�B?t���uG�H���p�=�n?n��?�9�?_�
>m�=9��#��>>��>��?���?�l?���A��>�����'�=�#�bJ�="y>rg>y�> 0?� ?IM?����T����܆��3ve��� ;���=��>u�t>��&>�ܠ=�l�<xt�=�7>o�>�,�>�#>Z��>��e>:����-���2?�В>G��>�/'?��>Eɼ�eM��/=�Q�=���͏]�3��������k%=Q��<�{=/ޖ�i� ?�;¿ׁ�?�F>���n�?���(��]�i>J�>qv����>�1>Ď> U0>n��>�->�V>\>��ξ�P>�J
�!�5E���S�oؾ�Ao>?Қ�l++��c��z彟�V�����}+��/i�����f�=�ˀ=��?e���D+s��"+��^�0��>��>�H9?�9���%v��#>���>���>�D��򾔿P���e⾾��?�N�?:9c>��>>�W?͙? �1�3�tZ���u��&A�N	e�c�`��፿M�����
�����w�_?��x?�xA?�H�<86z>���?R�%��ԏ��'�>�/��$;��B<=y)�>U,��B�`��Ӿɹþ�:��DF>Ǖo?%�?X?"WV���P��� ?�H5?H�?���?4�5?G�D?��Ͻ#�>f�-=Q�q>��i>��4?H�/?i+?��>�f�> ��=R^�����	�����Y��#�y���&��f�ؓ��k�=�v�Q�=��Z:�80��=���;�ޫ��DZ=��>��/>H�>Z�[?�t�>./`>��:?�� �M	!����=)?Q|�Iė�K��F��V��2>�eh?��?]pP?-�@>}AC��\K�k�5>%�o>h.>�F_>ǧ�>"x��:=�0ɑ=}R>�>��=/fb��y�o��G���Y��C�>���>Ŋ>���nJ>�Ȣ���u��a>:D��3���.G�F�#g1��Jn�ݭ�>S�J?/n?��=K���k����e�Ϥ)?2#>?�O?��}?�=i�־�@;��sH��Q�'�>���<�g�����\��UK:�V��;a�p>�&��7v��ab>��m�߾��n��SI�f+��xO=6��
"W=���;A־V'{�D��=�>ᬿ�K� ��Z��O⪿`�I?��n=}`����U�ҹ��>��>�>�<����(�@��h����=ʰ�>��>>�Z�*�CH�q4�Y5�>fOE?mV_?5k�?���	s���B�����mc����Ǽ�?4x�>�b?�B>^��=`�������d�G�!�>ڥ�>7���G�72���+���$�d��>�8?�>�?q�R?��
?|�`?�*?�C?%�>X-�����*B&?���?���=��Խ��T���8��F����>�)?&�B�㳗>��?�?��&?��Q?�?��>�� ��C@�4��>�Z�>�W�la����_>(�J? ��>]<Y?-ԃ?*�=>�5��颾=ܩ��_�=/>~�2?�2#?�?
��>�H�>K��B�=ڒ�>]d?��?�mo?���=N��>Ɨ�=��>��<���>>�>�?@rM?uYu?M�E?�X�>���;�
ý�đ�����K8i����`=Ω=����aq�r��6�=�#8<��ǼT���`ˣ�F�����`�!��c�>e�s>����0>�ľ�D����@>�v��n��Ŋ�_�:�P~�=:��>W�?��>>0#����={��>-�>����2(?c�?�?gA;��b��ھ7�K���>�B?3��=J�l�y����u��g=�m?F�^?ՂW�&��en?�4?�9"���Y�����]�Ҫ����3?�h?�%k��}�=ZH?|C�?4��>�W���W�
煿#�S�󗕾�=�U�>e�۾p�v��kB>��>?�˖>���>�K>�{���Sn��w����B?���?���?$Ƭ?>8�>�}����B����v��m`?Ĵ�>蠾(� ?F1��H�Ӿ先�d����,پy���{�����������Ow��'ѽ-9�=
X?]kp?�o?�xX?�>��b�AZ_�5�z�h�R�L
����9�B���D�q?�n�n�u�	"��ݫ���VY=�֏���5��t�?;n5? W���>����(��Nk���3>�aq��_��z�<#ߜ�'I9<�c�=�mI���1��u��% -?Bp�>R��>�!?�\�9�7�{!@��&)��a��>�?�>�U�>Ǐ�>X��;��n��ͽ�;پ�5��O�v��7v>�xc?Y�K?��n?4p�+1�����O�!���/��c����B>�j>8��>�W����M:&�jY>�B�r�j��w��A�	�c�~={�2?t(�>E��>�O�?�?�{	�zk��%lx�5�1����<:1�>� i?#A�>�>�н1� ����>�l?YG�>0$�>�p��>!�>�{�.�˽*��>�E�>�j�>��o>�N-��h\��j������\/9�{��=j�h?*w����`�Μ�>��Q?tpp:��J<��>S�v��!����(��>>/p?��=�;>v|ž�/��w{�"I���?%j?�R��K"�
ߥ>��!?&?��>6)g?@�)>BJ�]���I?�D?7bQ?A?C��>�l[=2S����'�;:>O�}>�I>V�=�HT>�,�ʦD������l=0ed=�I;���})�<���<S����vڻ5��=/ۿ��J�Yi׾���LQ��	��b��3���g���N/��U�����y��-�Z�%��U��c�� ��n�
�?^_�?����ʇ������0������eʽ>�p�V�s�0��h��f����޾ګ��F� �1�O��ii��}e�_�'?e����ǿ����:ܾ1! ?�A ?K�y?���"���8�P� >0B�<�1��v��x�����οL�����^?M��>���.�����>䥂>S�X>�Hq>\��'鞾V<�<��?�-?���>��r�!�ɿ]����Ƥ<���?�@wA?��(�Y��o
U=��>�	?��?>��0��_�b���[9�>�'�?���?�&L=ڬW�%��ɏe?p�<J�F��+�(��=�\�={=}�Q�J>�|�>�����@��_ܽ�14>���>� ��e�K^��ܻ<w`]>�Nս(Ô�"Մ?z\��f�m�/�yT��=U>��T?g-�>�*�=�,?�6H�%}Ͽ7�\��)a?40�?���?0�(?�ٿ��֚>��ܾK�M?%E6?~��>�d&���t����=�=�׳������%V�.��=)��>�>`�,���7�O�d9�����=���C���/���
�0=Z��;%���p4���ڽ坍�����I�:�"B��2�<3��=[�=>��t>r�>��0>��[?���?|"�>��?>��e�PF��(��͈�<;{��rｆ������K�ƾ�uо	+޾���! �u>��Hξ:�<���=0bR������ ��Db��HF���.?h%>0�ʾxN�
�<n�Ⱦ�G����r��֣��̾|2�Tn�ޓ�?p�A?�օ���V�=��T������҈W?ߋ�z�~7��.3�=>�����=!E�>٩=���3�8bS�v1?� ?�Lؾ���N�>ܯ���a�<��<?�<�>C�>⼘>�I?,���g��E�V><�m>�f�>y��>#�5=�軾����
�6?_uf?����2���ұ>�pپ�T8��6�=���=�)��, �=3H>>;ԕ��~�>=���>��=' `?��ƽݨ/�A<徦X,��]"���̾P��?til?K��>^s�?F��?􀶾ի���>��vq��1>��r?"�?�)>�<]�޾#��b�?��V?��>!������B~3��ص���S?١6>%�����6���}��?��v?�r^�zs�����:�V�a=�>�[�>��>��9��k�>
�>?#��G��󺿿hY4�!Þ?�@x��?>�;<� ����=�;?�\�>#�O��>ƾOz��������q=�"�>�aev�����Q,�Q�8?̠�?���>�������y]�=�ؕ�uZ�?M�?:x���Rg<A���l��d��^'�<`�=��	�"�s��!�7�~�ƾ�
������}�����>V@�w���>_8�=1�PϿ�	��cSоNGq���?c|�>i�Ƚ霣��j�Ju���G�y�H�����ꝣ>��>"˖�N^��.�{��N;�p��6��>���3�>]tT�x������.<���>.\�>h�>#����ۨ�?�.��Kοj�������X?�D�?�m�?s?EN/<�w�/�{��p�:kG?��s?.dZ?��"��J^�B>�>�j?^+����`��O4��E�n�T>+�2?�p�>�-��p�=�
>�=�>3�>S�/�ĊĿBܶ�4���Φ?%��?��_��>G1�?��*?2z�&��0����e*��b9��@?�P1>������ �;�<����
�
?20?"l��l�\�_?*�a�M�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?ѵ�� #�f6%?�>c����8Ǿ��<���>�(�>*N>mH_���u>����:�
i	>���?�~�?Pj?���� ����U>	�}?l%�>S�?�`�=�[�>�i�=갾�~,��k#>���=Z�>��?�M?AT�>�D�=~�8��/�-RF��DR��#�-�C�9�>~�a?�L?�Pb>.����1��!�jNͽ`h1�Q��rN@�-w,���߽�-5>O�=>�>��D��ӾK�?���}ؿuL����(���3?�>�A?�d��Kt��:�Ś_?
և>4��m%���:�����ӡ�?�D�?P�?<ؾ>`ʼ>��>e�>�kֽj��v���z8>[�B?O��
1����o�7K�>ٸ�?��@�ή?,�h��	?���P��Va~����7�b��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?ZQo���i�B>��?"������L��f?�
@u@a�^?*�Ͽjv���,���>�*1�<���<[G>8�m��pQ=���=i�<������=���>�@b>^�.>���<_8>!A>�B���$$������e�"�P�Q���:��[���)$5�|!����˾�B������������4���m�A3�=�$V?+S?y�e?@[? ��V>uP��eN=`?�o	5=��b>�z2?� K?�y-?ն�=*pb�rn~�!��� �z�<�>��Z>��>O�>/F�>uʖ�L<->��O>2�>�0>Dq=4	�<m@�;B\=>��>��>��>��a>��>^8���U���e��qJ�JZѽ��?MD����D�<���q�� ��մ�=1�2?x0>�ލ��RԿ�έ�9>?V}��ի�LK3�ϒ>�0?�gG?��5>�տ��w��p�%>>�ޡ��5	�=�ٽ�0'�b�$�D<>�*?C�>|�>��=��F�mD��,��)�_>�|C?�~��� ��kh��~L���Ͼ�2>X �>
�=���+���U��ܖx�Oӣ=SC?5g?��׽򴾩y:�����̞$>�X�>Sg=��=�c>�O��뽖�j�-׾=JY>��}>��?2��>�̂;��p>7`��h��N�>J�j>�(C��M?�[?�i��d�=Z��:�#��>K?b�J>��k=���1R>�@?櫊>R�<���;�_U;딣�-٠>�>ڽ���&ZL=��'>A���(��=� �;�T�$�O�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>�-�aj��8܆���u���"=�.�>`�G?_W��D�F�`�>��O
?�T?Vj��ڪ����ȿ�v����>i�?d��?Іm����Q@�:�>1 �?V1Y?f�j>��پnT[��Y�>��@?�vR?i�>���{'���?�?��?�J>1P�?L�r?t��>��t�d�.��j���)�w=̆�;�a�>O�>�����G��ԓ�Ut����j����Ye>$=�
�>�U�Qϼ���=�B��A���~Vg��t�>��o>^?H>}֝>ߺ ?<��> ��>v�=]������^���;7V?�G?� :��P���C���M>�䉾j�?�^?�ֽ�����>;�Q?C�\?��^?���>J��6D������6����c:=��=J��>�}
?p�ZT=�6N��� ��>��?`��.��M���A���>? ?��?���=�.?k�>Ԋ_�EX>{8i��Ǚ�T5V�MP�>�>��?��~?7�C?�T��A�Q'��F���a}�P��>L�?�I?DZ�;�0������Q�� ������Ƣ?� �?.�m���(?˹�?ֶD?Szn?�2�>8�ž��m=�u>���=��'?@���J�)�5�3P3�ڥ?5� ?@��>N����h��6��Sɾ�"?C c?\-?M�bx�/'ھ��<CA�<��vtH�D?�;�[H>���=:�ʼ��@=|N�=G��=g�D�^~���5<�>|�>%Y�=�Ug�v.�:?,?�C�\�����=�r�u]D��>��L>0a����^?ON=���{���l��1�T�U��?G��?�[�?����h�G+=?(�?�/?1�>/���0޾C��I�v�U;x��i��t>f!�>m�n�������{���>��U�Ľ|��:��>'�>��?Je ?mU>D.�>� ���(�L�ξ^l�V�]�����I�ݽ/�����6��d�+�B�<X漾e>l��L�>��½�ۨ>ʱ	?�qt>��l>��>U
���%}>�Mc>�7{>�ޛ>}X>��(>r��=`E�<���MR?^�����'���辪����2B?�nd?�0�>$�h��������{?���?�q�?�Gv>,yh�.++�:d?0�>(���q
?;D:=(��^^�<�F��5��;'��R%���>v[׽�:��M��ef��o
?�7?�^��J�̾F׽�A��/�<��?�?��.�߷E�𨄿bX��1�f�ֽc��Gly���9�3RT�m���$�c�Q(���9���=/�P?��t?$�K�Ri,�L`�͖���N6�Qo�>1��>w�t>+8�>�>�>Z�Pt2�[�d�XN�Տ�n��>G��?�XB>v�]?�)?�?��H?�y�>��%?+{p�E̝>�+(�c��_�>M!P? ?l�H?��!?j�5?���>}P��9�վn#��>�?��?|W ?x0�>�?�`4���L=��{��I�<"�Y�5���U�L>��>qǕ�\�
�!�=��>)�?m|�ϭ;�f�=o>��5?Ķ�>&H�>�S����L� <�
�>+�>>P>���t�`��U�>ﺅ?v?���=�>GQ�=����5<jj�=��ݼ_@�=�;ȼE�w��l�<��=1o|=�@N;�@��S�����<V%<8u�>)�?���>�B�>m@���� �M��j�=�Y>yS>h>UFپ�}���$��!�g��^y>�w�?�z�?��f=�=��=�{��-T�����K������<��?�I#?bXT?<��?m�=?vj#?��>�*�YM��j^��N��خ?�8,?�>!a���˾����0!3��>?��?	�a�ݿ�y�(�`;þ4}Խ5	>"�.�c}������C��û���|җ�W��?�ݝ?��D��6�&D�-�������d	D?��>!J�>F�>�n)�~�g��A���<>8��>�R?�#�>��O?<{?��[?jhT>��8��0��oә�dc3�z�!>k@?���?�?�y?�t�>��>��)��ྂT�����G����?W=	Z>���>C)�>�>3��=CȽx_��"�>��`�=(�b>,��>��>!�>F�w>�A�<�NH?r��>ӫž�i�����97����P��7w?��?��*?HX=P|��	D�����Y�>�#�?.��?+(?�^�	��=1���%�����d�l¶>���>���>N5�=��=9�->�9�>�ɿ>'�+1���8���w���?�H?��=Y�̿�~���#>SR`>��=�|=�h$۽F�ݾ� �����Y|&��*�a袾ց���$E��I8���վm���k�*���>��'>Ý<��=�^>���="��"�<OH��\/�=�����=��*<Ɲ�� �����a=�>�<�]�=�?���	پT�u?��G?��3?�K?4k>72>~c��Xk�>7����?!vc>ȗ���E��f�'�w���瓾�-־�#�W�+�,����J1>�U)<��>�`>>n�G<.��<U(>I�=8>έ;"�&=-��=��c==��=��
>� �=�">�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>|a>�A>��]�*RE�)�7�H�:�b9j��.?i�I������;|>��<(�Ӿe�˾fS=o�i>"z�=����b��?=�e:��&�=��=}�>l>ߌ >
�o�v��;��>^�>�>,�G-=���������m>30�>X�6>��>��?N^0?�Od?B�>��m�Ͼ�0���J�>���=^2�>!��=�mB>L��>O�7?��D?��K?���>}��=O��>��>ٖ,��m��l��ϧ�4�<[��?�Ȇ?���>��P<-�A�����d>��FŽEt?zR1? f?N֞>�\
���ݿ��	�t�V�L�
�=�3c=����/�� )�Ŝ��Z���>�>~��>�F�>B�A>a�o>4=>���>��W>iR�A��<��Q�1g(��f=��=��<�K|=������=]�3���w�<�=2�JL�=]&�=�o+<J��=;��>��>��>&��=6鳾�!/>�Җ���L�1^�=YS��)B�44d�1s~�"/��6��bB>f�W>���B'��.�?��Y>|N?>�z�?zHu?� >z��i�վ<��\�e�cS��a�=�3>��<��m;��T`���M�b\Ҿ�� ?��O>t�=En�>�Y���6�sV|�Djྪ)���?�?��q��Ts��JL���ԭ�Π��	p���Ӽ�|?)c���>��F?��C?�מ?#�/?�w=�,��q�H&="��XX'��ͫ��bʾ
�4?ٞ?�\�>h����J�&%̾���L��>�?I���O�2���׭0��v�Sͷ����>������о�+3�~p��������B�9�r�K�>��O?��?=8b��Y���[O���粆�dn?�g?�2�>W>?�B?t���uG�H���p�=�n?n��?�9�?_�
>m�=9��#��>>��>��?���?�l?���A��>�����'�=�#�bJ�="y>rg>y�> 0?� ?IM?����T����܆��3ve��� ;���=��>u�t>��&>�ܠ=�l�<xt�=�7>o�>�,�>�#>Z��>��e>:����-���2?�В>G��>�/'?��>Eɼ�eM��/=�Q�=���͏]�3��������k%=Q��<�{=/ޖ�i� ?�;¿ׁ�?�F>���n�?���(��]�i>J�>qv����>�1>Ď> U0>n��>�->�V>\>��ξ�P>�J
�!�5E���S�oؾ�Ao>?Қ�l++��c��z彟�V�����}+��/i�����f�=�ˀ=��?e���D+s��"+��^�0��>��>�H9?�9���%v��#>���>���>�D��򾔿P���e⾾��?�N�?:9c>��>>�W?͙? �1�3�tZ���u��&A�N	e�c�`��፿M�����
�����w�_?��x?�xA?�H�<86z>���?R�%��ԏ��'�>�/��$;��B<=y)�>U,��B�`��Ӿɹþ�:��DF>Ǖo?%�?X?"WV���P��� ?�H5?H�?���?4�5?G�D?��Ͻ#�>f�-=Q�q>��i>��4?H�/?i+?��>�f�> ��=R^�����	�����Y��#�y���&��f�ؓ��k�=�v�Q�=��Z:�80��=���;�ޫ��DZ=��>��/>H�>Z�[?�t�>./`>��:?�� �M	!����=)?Q|�Iė�K��F��V��2>�eh?��?]pP?-�@>}AC��\K�k�5>%�o>h.>�F_>ǧ�>"x��:=�0ɑ=}R>�>��=/fb��y�o��G���Y��C�>���>Ŋ>���nJ>�Ȣ���u��a>:D��3���.G�F�#g1��Jn�ݭ�>S�J?/n?��=K���k����e�Ϥ)?2#>?�O?��}?�=i�־�@;��sH��Q�'�>���<�g�����\��UK:�V��;a�p>�&�����2�_>ث��Y侗_n���K�C���Y=|R�#�`=#l�RӾ퀾L��=~>n��)$���������LJ?�\W=K���^�\�G���*�>3��>Q�>#8�X*��KC�'���=��>��I>�,C���󾷋G��!��>�>�QE?�T_?#i�?v"���s�
�B�����d��D�ǼO�?t�>�i?�B>W�=r���}�Q�d�[G���>_��>B��$�G��6��+,���$�ׇ�>�7?�>��?�R?y�
?Ԝ`?�*?KB?c�>��z����<&?z��?�Ȅ=��Խ۝T���8��
F��>�h)?�B���>��?N�?��&?��Q?�?��>Z� ��D@�)~�>�[�>��W��P���5`>6�J?���>�6Y?׃?�=>s�5�9���h��Vc�=�!>��2?#?2�?ָ�>���>bج�6��>���> k?��v?�~?@���C�(?a��>���>1�=�(�>^��>j�$?��*?�Fz?b�P?Q[�>ڽ=��1���������
���u��{ۼSeO�"K=U�>Ҁ�;$�=�R=�j�B���tu��]�=<s{<� >ml�>�zt>旾*N*>7Cľ�ӆ��?>�vy��l���Ȉ���9����=��|>�� ?u�>�!�H��=k��>]$�>j���(?��?<f?���:�b��xؾ<E���>*A?~�=�Ul��ɔ�\Cu���e=H$m?h._?��Q�ϙ��y�g?�QH?�e����'������ʣ�8s��M?�j?= ���>���?])k?��>�o���x��啿�+N�	����=�H>������[�>�dU?!��>�#�>���=����������?3�g?�,�?��?h>�����tۿ	*������S^?��>�g����"?IM)�b]ξD���۲���ྡྷ)��Qe��e锾w���\#�Ճ��`ʽL��=�)?<jp?Q�o?Ib^?�
��d�Y�_�8~�LwW�X������-D�ǕD��]C��{p��]�r|������1=\~��͊h��$�?��:?_�����?(�����̾�k�D�b>I�>�c�[Q2>�����f��S�=�������K����I?��~>Һ>�%?�􀿐�N���h����6"$���>�'?��>�3�>@"��ө޾d���ȑo�VY��7v>�xc?C�K?|�n?Bp��*1�����0�!�e�/��c����B>�j>^��>��W�X��7:&�UY>�?�r�i��w��+�	���~=l�2?�(�>I��>�O�?�?�{	��k��lx��1����<11�>� i?A�>��>�н"� ����>?�l?|��>H-�>橌��o!�$�{���ʽ.�>O�>���>��p>Ҟ,��"\��k�������9�0�=-�h?fw����`���>a�Q?�KE:?�G<�n�>1�u���!�5���'��>?�? ;�=��;>�Fž��y�{�V��G-?@$-?w�G�����>�a&?��>��>t�h?���=X�쾐�����?$$Z?Ю]?!Z:?��>��=���r���&��È={�8>U>���>��Q���,�˷	���4=W8�=�D�����ؽ�|�;�:=`o=�A>�lۿ�DK��|پ����E
��ۈ�t���^��`���v���9���bx����l'��V��"c����w�l��?9�?WT��������	�������j��>�rq��u~�᫾r��v��Ds�����`!�B�O��i���e�KkA?�0̾�x˿�k��kF	���>!�>���?��dI�^L۾Q]_>8���>л������ҿ����P/M?k��>���3Ly=�1!?�Z>އe>��!>�W�6ݺ�?2�Gc?f�
?���>1	���������C>��?��@��D?�d$�n� ��xi�ĥ�>{N?X�%>1��������SG�>I͚?6�?��<��P��FR�Qb?�r�	�I��2����>2�=��J=~zڽ��@>�B�>���	2o���z�� e>�t>�����Sd�L͎��B�>�ͪ�S�}�Մ? z\�ef�t�/��T���V>*�T?D,�>u4�=��,?�6H�}Ͽ��\�#*a?h0�?���?[�(?vۿ��ך>��ܾt�M?KD6?1��>=d&�z�t�M��=�6�?�����&V�$��=٬�>�>р,������O��K�����=	���}ƿ�"��.�G����;�հ?�m��򐈽u���M���f�����kf�<W�w=��E>O��>��=>o�o>4KR?��i?�,�>�>+>3|��O�����ʾ<s������S"���s����S�����ʾ3ξ����4���|��ɾJ&���c=@�E�wˍ��-��n�-uY�I�"?�w=鮔�Ik�D� =�^�@\��g��e�ٽ����-�Ū�1��?S[I?{t��s�
� �ʬ����O���[?�J�����D���ȇ�=d��s�"=ee�>>�,>��	���D�ݷ_��,7?R�*?�վ%�O�B:�}M<EdM=z�V?�P_>��>rO>� ?!���(�b��M>�ʩ>�_�>���>�Uμ`8Ǿ�r;� )?�b?��*��΢�̸�>����MG� �=k�=h��-�=?��>)z�=�"�5��#��<'=)W?6��>��)�_��g����m =='�x?��?�)�>�zk?Q�B?��<�_��n�S�T ��4w=��W?h(i?/�> {���оw��ƾ5?�e?�N>eh������.�1Q�P"?{�n?�\?y���	t}�P������m6?J�v?v^Z��A������KW��K�>��>J��>��:���>��<?5�'��ؕ�������2�?��??@q��?�Dy;�L3���=�+?6��>�wW��#ɾ�қ��Z���^=^�>t
���ys�Z\!�l�,�N�6?<�?���>�|��\�&��=�ں�Gh�?*݇?x>���YN�%W ��&b����w?�='a->;�'���Z�u���K��NӾ
��ǫ��u�����>��@6�=��o�>�ɜ���-�ӿ�݄��}þN�-�i�(?Q��>ot=��4���m�UIv�"�M�{�H�8´�
m�>��=mx6��߾�-����Q��yu�w�>+��m�>���;v��ä�� ���&>� �>0�»F����/��?n`�8;ܿ�w��ٹ��R�^?�ҟ?��?I!?��n������c��<4?p�?� �?�
|�Ƒ�bL��:n?�c���e�;���?�4ٹ=
?#��>��-��F��SA�>R
�>F������ǿ�@ÿ����ѕ?R��?����?�Õ?��,?�� �W���P�׾��?�uv�=T�N?���=m�O�f��zN�vq�����>I�9?
��`�U�_?��a�C�p�|�-���ƽ�ۡ>��0�e\��P��£��Xe�	��i@y����??^�?c�?���� #�E6%?��>;����8Ǿ��<׀�>�(�>�)N>TI_�z�u>����:�Ki	>���?�~�?Yj?���������U>��}?�1�>i0�?��=���>���=�l��9�*��%>���=ȩE��z?3�M?�6�>���=�[6�A�.�ϵE�V0R�\`�ёC�=H�>M�a?L4L?�wd>(ܷ�uK/�0� �D�ɽ"w4�eZ�]<��..�%�޽h�5>K�<> >�:B�@WҾ��?Hp�8�ؿ j��#p'��54?!��>�?��f�t�^���;_?Gz�>�6��+���%���B�]��?�G�?9�?��׾�Q̼�>5�>�I�>�ԽJ���_�����7>/�B?^��D��q�o�x�>���?
�@�ծ?di��	?"�{Q��&d~�����6����=��7?4��z>C��>Y	�=�nv������s�D��>�B�?/y�?S��>�l?�zo���B��2=bJ�>��k?du?`�i����B>��?���Q����J��f?-�
@>u@͠^?}뢿��ҿ���(W��Sƾ¦�c���w>�0"�=0r>�S����~���Z��,<f��?�=�{>z/�>s_�>��U>,����� �
���I����j�K�'�˻�S�x�9��</��>1��̾
��	ء��'<���&�j/i��mf� �;M�=��X?]�F?O�d?$�>A�;΋>E.征��/R2��x�=��>>�7? (F?�-$?O�=%W��"�[�m"|��*��"�I���>èU>���>���>&)�>$q�<�|>
��=�qa>��}>p��H5<&�z=��<>��>��>h�>���>��ռI���zſ,�d��,[�_p���c�?FI��V+�m�u�r?A�8�v��'�u?�i�>�f�����9����&?}��P 8�^I^��FC>��G?_;G?b�>�����at=�U;&�ý�Q��r>�Y�:Z�i� ���(�>{#?��q>�l�>l~2�&4�P�����bMw>�8?�V��J]��q���G�7;Ѿ�eG>���>��g<���e���߁}�r�u�Я�=Y[6?�?I9�������!t��$��^�F>��2>r�q=쾷=XRs>Ev�˚�;rW��6�<�=;�R>��?�pc>�:=��>O������_�>���>�s�=��B?S�?_��f������0�*��>۳�>a�:>�=ík�>�=���>��u>Z�Q;��2���Q@d��EA>�����,�� E���+>�׼�}>hs=��'��DX���<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>�x��Z�������u�d�#=��>�8H?�V����O��>�w
?�?�^�ԩ����ȿF|v����>R�?���?K�m�nA���@�p��>%��?�gY?Qoi>�g۾�`Z����>��@?�R?��>�9���'�{�?�޶?ޯ�?]I>O��?Vts?���>xy��w/��?��������=�k;��>b>�����fF� ݓ�?�����j���Sb>�z$=��>���H���_�=�@���\���8f�-޷>p�q>*�I>?��>�?�(�>{֙>�T=�؊�����d薾�YJ?C�?<7��j��C�<nļ=�6Z��?�+?X���b�ɾۥ�>t�^?޹}?�P[?Ў�>L�	�	���M���������<��O>���>h��>�Zq�m�I>@�Ѿ1�9���l>�Ж>��?<C�Ծ!
}��ci;�J�>@?·�>&��=�`.?��?1�=?��>5�D�P����v���>u��>�?Q�?��m?�����B4�u��E�ſa[��I�>��?SU?�O�>:�a��*���)�Y��Mk���Ik?�y?��=x�>��?ۈ_?F�?PJ�>��<����Y�
��v�<��!?I]�ǘA���%�Xk�̲?��?���>�����ҽA�ݼm��P(���?R\?�w&?3��~a���þ��<ء��d@��<�����>��>�-��l]�=>���=��i�I�1��6�<��=ȼ�>���=��5�Ӥ��S�,?j'`������=F�r���@���~>L�]>i�ľ�j]?��>�D�y��ݭ��S��þR��ۍ?�V�?�<�?�½Ųg��~<?�T�?�g?[�>jK��$�ؾv޾Ku�`t���b\>x�>�&9�X��Ŕ���
����������"�Ma�>w�>��?�� ?S O>��>��v&����[�E�]���� �6�V[.���5�����#���	�����g�w�&8�>F=���V�>�
?�k>��y>}6�>R>��=O�>c�V>�}>2��>�W>�4>{>1�;<��ѽ�NR?n�����'�N�辁����)B?{dd?=�>HPi�T���ҽ�-�?V��?%s�?C-v>r�h�2+��f?4I�>W���o
?��:=����u�<zQ��Z���A���i�$��>~$׽�:��M�,ff��\
?�'?����̾��ֽ4J���	���:�?	5+?(�6�+Z�
�t*P���l�N�=:�w�ň��>�'�Da�)ћ�Ą������B5��??���?�^!�T��T+ݾj+��R+M���@>4��>{C�>��>�t>���n�#�^ N�t\�j����9�>:*H?��]>�4m?�?*d2?(	M?��>�,�>Lb̽c_�>NN���5=�4�>7�+?�"?$�L?�'?;?:�>����޾�&̾��?��>�E?<�>ٸ>Y���j�u=���+PV�<ξ�ց����=���<b���nʽM��=As�>V?~F�?�8�����Rk>:�7?�v�>��>���F��s�<�+�>3�
?�F�>P����kr�Z��I�>*��?�4��=��)>�1�=F샼�Vں6��=����Mk�=n���`<��%"<�'�=#�=�}q�[�Ƿ�:�C�;TŰ<�t�>}�?~��>�A�>.@��֨ ����m�=o
Y>qS>0>�Dپ�}��h$��/�g�`y>�w�?iz�?'�f=7�=%��=8z��BR��A��0������<��?{I#?MWT?���?M�=?�i#?7�>R*��L���^��n����?Tf<?&�!>E�!�J	���֣��U8�H�>��?i=e��K��(p;�k��Ԩ��ٜz>�U=������SO@�)e>Q,��8^=���?o�?��C=.�+�־���ˢ�e�.?�)�>"��>��>2=/��~z��G+�+c>W �>@�T?��>�O?6{?o�[?8[T>am8�,���֙�qA/��w">�@?⤁?���?�y?���>M�>�T)���3;��-���6�����NV=1Z>�z�><�>L֩>Q�=��ǽ�᰽��>����=NIc>D��>2��>��>Z�w>禮<&�O?���>���*�/������
�ժ��ߴz?�Cr?�z6?9��<���A���>�O�?��?�d?.Ϗ��o�=�j�=��`��D�/�>W��>MB�>8�`>�����)>d7�>�>p���*h�W�,���ǽHP9?Hb?ӌ�=�Jοvu���ܽ{t8��[��޾J�����,���]VV�UV����9����듾�N��f���`I������@�B��>�s>�*�>B�v>Y�>��=�O�xܖ�ά;`>��=�
>1~�=8$l>��|�vt=	���&�K�x��u�о�Ry?�J?nY,?��E?�f{>V{,>.}���>j��0�?rdV>��@�5��y�>�����=���{Ӿ��ҾLA]����[>�A�F�><�0>��>�,�<���=v�k=:�=^u�;g�<�="?�=�x�=�1�=��>�	>M6w?����걝�k3Q�yo�µ:?B8�>Y��=��ƾ@?^�>>>1������c�+?���?�S�?9�?�yi��^�>e ��yӎ�Ȍ�=����92>���=��2�U��>��J>���I��AY��]3�?b�@r�??�ዿ��Ͽ�^/>yI>�=>??N���*��x^��W'��RN���&?�@��ɾ/s�>7Z�=����v��	��=��J>Ӫ=�9��]���<=����x�=_{�=ď�>n�E>a��=���h��=��u8�=i��>�Ub;���pF��Gڭ<]�=��|>�`>��>� ?�f0?$d?�t�>��l���;/v�����>��=t��>�"�='5B>���>�38?��D?��K?_�>�a�=㨺>��>�P,�0Ym��m����L]�<�#�?���?�[�>Ig`<}�?�X{�v�>��Ƚ!Y?�f1?X?��>���ݿۻ���)�����U��! �<�?���E�V\���e��=���=��>k�>�#�>F��>@�>��q>���>��N>��	>E>X`F=]g;�C�<'r�<�ǽ��*�\3�;R����#<q2=s�E=��	=�k��W#��5�Ϡ�=���>�'>X�>��=�P��=/>n0��_�L��b�=󂧾�"B�#Ac��z}��.��1��VD>��S>~1�����k�?5/Y>H'@>�*�?(�t?�r> ��LվhN���a�M�R�K�=�
>��9��u;�h&`���M��'Ҿ���>�]�>��>�zp>o�+�@~?��]i=~���E5��l�>�?������jp�#~���}���Pi����E?��� �=��}?�I?t��?�k�>����Cھ��3>�&�-�='E���l��C��
;?A�%?u��>�龏�D��?̾����ҷ>UI���O�&����0�����η���>������о#3�8g��j�����B�2Ar���>��O?�?a)b�U��QO�n���/��mr?s~g?]�>�K?C?m.��J��]n��vm�=n�n?c��?a>�?|>N21=�kJ;D?vE?�y�?+��?cҀ?���T/�>���<=9/>��A�+)�=GH�=�H>�>y�?�?w�?�D�x��FɾYnپ�����&<D5c=	#>�>�l�>V��=jb=$%�=��>�I�>P`>V�G>��>Ed>��~����9?/��>IY�>fl*?奟>�䞼�����5=T���c�I���.���U=����m�=������=�8��Q�?�]ѿ02?��*>Ȩ�H�0?��.�G�@>��&���J>�Xa=�#{>!M�>�N >@ci>�>��~J�>�<&>!NҾ�K>a?�H�!�":C�˒R��Ҿ=�{>$o���&��3�����I�0����!���i�:U���C=�5[�<�+�?����gk��N)�:[����?��>S:6?���
��d1>���>�W�>.���z���^ۍ������?X�?�;c>�>,�W?�?[�1�k3��uZ���u�9(A�)e�S�`��፿���
�<���_?�x?/yA?�P�<�9z>4��?��%�^ӏ�V)�>�/��&;��=<=;+�>�)����`��Ӿ��þ�8��GF>p�o?0%�?fY?�SV�X�.���>��L?�!?��?0T?�T?�,��W� ?���=瘔>�m�>��?�f ?��>���>��R>�e�=�e>W�P�3�z�7X1��h�W>7= �����E>X��c��=y�=�C�]�������l=��>���=�>B��=�M�<���>8�a?q��>Yl�>I4?�W����$�Wn����)?�</���罎�~Ԕ�+k��:&>A�f?Ž�?
�Z?��U>�fE���M�6�>�X{>��>�O@>�>�>�F�FB�3�=%)>�Y->n��=^ۤ�C*���T�m.���=�a2>���>Jy�>����k&>s�����t�=d>�-L�i3��&R�2G�ɺ1���o����>��K?t?[�=�꾡���h�e�a�(?~�;?�/L?<�?�S�=@�ھh9���I���#����>���<�*����������:��:���t>�ƞ��z����a>���O@޾�n�J��	�>�N=�W�3fV=x���[վ�~�M��=��	>����]� ��%�����dJ?��k=6����V��R��7N>�-�>R�><8�,:v��@�醬�V7�=���>t%:>����_���gG�kf�F�>�JE?�H_?�h�?�'���s���B�%����^����ǼI�?��>;d?d&B>6�=������C�d�G���>v��>~��S�G��=��5����$��z�>�;?8�>�?9�R?��
?0�`?c*?�J?)�>�=��7���N&?π�?���=��ս=�T���8�ZF�C��>�)?B�R��>nf?��?@'?��Q?�?J�>� �(r@�v��>I��>�W��`��2�`>��J?P׳>DY?ă?��>>~�5�[���ʉ��R��= �>��2?�H#?��?P�>s��>��׽'S>>X�g=�Gt?�?,[�?T���3?!G�>_q�>��?�Ov�>r=?��?Z	T?oy?��S?�	�>ŝi=Pȗ��e&���m��(�<�z>����}u=Ҹ�q����E�=Ȅ�=��=�9=�����@=�ܭ��ϯ�)=:k�>�s>�#����0>��ľ�D����@>L����G��W����f:�O&�=�{�>��?I��>�j#�͒=�|�>�E�>����0(?��?:
?� ;��b���ھ��K�h	�>E�A?4e�=��l�v����u�:�g=��m?�^?�W��2��Ӽi?��?��,������Ծ�G|�r�)��?���>�Vu���>$b?Y8K?�	?x�@��U��u��S�|���f�h�=�>�oi������>��I?�>z�ݽ֚<>p5����v�6H�.?�?�7�?�`�?�&y>�~=�7�⿭���Nt��V_?e�>si����!?QD����ξ�O������`�&z��@d��ژ��Τ��= �Q���A ڽ���=e?�'r?]�p?E�^?� ���b�|]�	0|��zT����[�r+D��C��C�b�n��5��B��v}���;%=�_¾�,��}�?��I?�'����>��N�w)���&ǾW�>����h<���������\��;�k�=Vw�iax�na��b	4?���>|�>�C?�UJ�C�3�@�A��������le>@	?�e}>[N�>��Q�"���	#� ������p��7v>�xc?R�K?��n?Up�+1�����L�!���/��c����B>�j>,��>/�W�˝�V:&�rY>�G�r�_��w��<�	�
�~=��2?(�>J��>�O�?�?�{	�kk��-lx�4�1����<11�>� i?!A�>�> н1� ����>�h?x]�>0�>����� ��4{�����>v��>*?�q>d�6��\��	���]���9�p��=|�l?ݿ��u�`�N�t>�U?I<���<���>6V����%�*>�X�1���=}�?�2�=�N>-�ž?���c|��A��lw?��?�݅�Xv=��>��/?���>��v>��m?=׮>j�Ͼ%f���X�>X?�
E?R�C?�?�5�<=�p�սa��^j�=.À>��>B���6v�=^�4�l�e���S��� >M�)>�hG��Ř��M�;�o�<ԃ�<�A=��
>�kۿ�AK�[1پ�����&
�����@���u����w	�𐵾�.���x��$�g&���U�Aic�B���wl�Yr�?&4�?�)��D��&�������w����>��p�~�V׫�;�����Ζ�j���^!�L�O�*�h�X�e�]�'?Ⱥ��˽ǿð���;ܾ=  ?_A ?��y?��#�"��8�Q� >NV�<'+��j��њ����ο�����^?���>	�Y3�����>?��>֡X>mIq>���8螾�1�<M�?�-?���>e�r���ɿf����Ǥ<���?�@��A?��$�)��n�=���>��?��(>�"�h�<����#�>�n�?
%�?^]i=��S�yh#�v�b?{%���C��ܻ!&�=��=j��<����97>ۊ>r��q8��a�p$>��>N{ɼ�a���b���0=�k^>��ֽG(��4Մ?"{\��f���/��T��U>��T?�*�>=:�=��,?[7H�]}Ͽ�\��*a?�0�?���?+�(?>ۿ��ؚ>��ܾ��M?bD6?���>�d&��t����=�4�ڋ������&V����=S��>Y�>��,�ۋ���O��I��+��=; ���ǿ�/��I���;�����3)��`)�k���/߰�OT��x����3��r��!�=�V>
m>�X>bl>��P?1.m?���>ش�={�ҽ��b��4���tW=<9H���۽ |��|f<���������{��%�����,���<��m�=3R����7� ��sb���F���.?�$>�eʾ��M��0<fʾ����˃�$󤽩v˾D�1��(n�3��?(�A?vȅ���V�#��M	�����6�W?���V���笾� �=&|���J=��>�H�=���X�2�A�S��(?��>?n���Z]����O>�O��}�=I?[4->��=[�=gB ??�m��t.�>Ɉ>!��>֝�>��
����:E���?���?ʟi��=��O��>\����4���=�f1>6;����=ԩ<>�C>����D�d��9$>�%>YZc?y��=}4���ľX�
��׋�>v:����?)8?v�����?��p?��3=~��{O��s�W��A��w?{?��
>q������T+ɻ/ <?� j?�zI>����w����ً��OC=>�~�>y��>��p��'(��~g��M�f5?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������5u�=Zߕ�	^�?�?}}���Zf<��*l������֠<��=��"�@����7���ƾ;�
�y��� e�����>cU@�a��>�~8��2⿱VϿ���Ldо+tq���?Ë�>k�Ƚ������j�[Ru�0�G���H�՛��p_�>��>~���͑���{��i;��퟼�!�>���T��>
S�/�������1<HҒ>�x�>���>�>��[���r��?L��u8οͨ����ޱX?�\�?�e�?�g?5�<<p�v��Y{��{��5G?��s?�Z?��$�%u]�A�8��j?ﳪ��r`���3�θE��
R>�Z2?D��>��,�a�u=4�>~��>3>.w/��Ŀ%���P�����?<[�?���֋�>88�?�H+?d��͑��~멾��*���:�@?�2>�9��^�!�*�<��X����
?�0?����]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�"N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?V��>�΄?���=��>5�=6f����Q�&�#>��=.P=�Q�?��M?�T�>��=59�X!/��4F��R�˽�_fC��N�>�Lb?{�K?�Pb>�ظ�z�6�dW!��6˽�Y1�$�����@�^�#���ݽ�3>;�?>�><XD��Ծ��"?�i��DտgL��v�r��?�)Z>|�?Hپٰ��)��<+Bl?ސ�>�$��m���^��� &�N"�?<�?�V?�z̾�C�LG>�.�>/�>|����|ν3�3��k
>tY:??����֋�P�i�O�|>%׼? @�=�?��g��	?���P��Va~����7�c��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?cQo���i�B>��?"������L��f?�
@u@a�^?*	�ĿZ���[*6��A�s���P� >��d�.f�s��:=����=鿽�UR>�3�>9S�>u>���=� ^>wd{��&�ސ�y�f�w�i�r�1�%�A�}+��l�/��~���^��[��7�x��<t�*��rʾP�y�����3�=�X?/P?Q�o?@8?%�6���.>����fw-=���u=��>K�5?,0G?$�,?+��=������b�v����E���>��V��>��R>8��>���>��><h�;�c^>��+>�n}>k��=:f=��p<U��<ΉO>y��>���>=ٲ>�C<>E�>7ϴ��1��C�h��
w�x̽5�?����4�J��1���9��Ѧ���h�==b.?p|>���?пk����2H?���X)���+�!�>B�0?�cW?k�>7����T�f:>Q����j�D`>V+ ��l�Ŏ)�&Q>el?�vk>a*�>��2��:���L� ~��Hpw>4�7?�K���"2��v�bFE��~ܾ��I>}I�>d�������k��#v����g�餀=�9:?"?��ʽ������j�ᔾ�G>�:K>�)=��=bJJ>��X�e跽��F�ַ�<��=�AX>_�?�c6>�}g=b��>8���I��t�>�7E>�>+�??Ą ?Q]μ�"h��o�Mm���p>��>��|>�; >K��i�=���>��a>�ܼ�|��V
��]��|j> ���LNe��$V���=���-��==���J���<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾWm�>��<�c[���w�e���%��r�>��[?=׾�夽aI��ؑ(?�P?*(������Bпzw��D�>o�?R�?��g����po"�A��>���?=T?��>g����Ib��F>�;6? �0?��e>����Ue�O�?r��?�j?�I>���?�s?�k�>�1x��Z/��6��閌��o=~[;e�>�W>|���|gF��ד��h��v�j����2�a>��$=*�>RE�l4���9�=��I����f�+��>-q>�I>W�>y� ?b�>Ħ�>�y=�n��^ှ������P?��?W6-�����>˕�>I��,�W>�>%?�(�>����Z>��Y?]P�?��M?��>5�������N��~u���6+>h^>��>Q�?ĀF=
Xe>>
�����ݕ>���=��=���׾;߽ӛ�>�W?p��>ܷn>%?��>A�=���>��Y��X��-�Y�#?��>��>�׆?�37?�:A�`�0��&��V,���G|�ѫ�>cy?�X ?�=>[���iu���)�c���y� ��Ҁ?�I?y���&	�>���?~�k?�WS?;�>!�Pl�k�Pw�>M�!?#@�֛A���&�k��.�?�%?��>�9��}oӽ-��˱�>H��~�?l�[?|S&?M���a���þ�X�<G��\+���<b�U�0O>p<>t����w�=9h>&�=�l��j6���d<m�=�h�>���=�6���/=,?�G�~ۃ���=��r�7xD���>�IL>#����^?}l=��{�����x��	U�� �?���?Xk�?���<�h��$=?�?W	?d"�>�J���}޾7�ྴPw�~x��w�Z�>���>X�l���G���י���F��R�Ž��R�>���>8�?�(�>�BK>ꨯ>Zߒ���&�����o�\�[�@9��.�<f��Q���� ��+��JL����v��&�>�z��X�>�	?]Nc>D!z>w\�>�,�;�-�>HT>>Ic�>w�m>�7>ٻ>���0m�'UR?����P�'�j~�m�����A?�'d?x�>��e�?����v��?gm�?�Z�?��t>�h��5+�ۀ?�}�>���d
?�.:=���>;�<X ��5��5���A���>��ֽ�6:��M�xf��C
?m1?������̾ֽד���*�00�?��?��0	K���o�P4+�]f���w�_�%=ځ���0��v~�2���ub��1����5����8R?E�?O} �I�*����Vxw���k����=�L�>聝=�	?,D�>dľ0�Im�pR�� �q'?�q?��>Yc`?�/"?etA?�D?[�>e��>����N��>�՟=�'=���>��R?F��>�!D?
9?e�9?7tj>�������=�����?�I?��&?d�>Tj�>�(��(w>-��W@��r����ȼ���=k�F<�������Ი�
��=�x?�4��8�c+��c�h>��6?���>��>E������w�<@��>��
?�,�>QM ���r�7����>,��?���>�=�)>6&�=?�y��HC�:
�=����V�=%���V8��<}7�=b��="�S��!Q:���:#�;�< u�>>�?���>�C�>�@��!� �X���f�=pY>@S>E>�Eپ�}���$��d�g��]y>�w�?�z�?ºf=��=Ö�=�|��OU�����R������<�?-J#? XT?\��?k�=?[j#?ܵ>�*�hM���^�����®?�$,?�w�>���l�ʾ���3��?�]?v,a�w��+)�_¾��Խ#�>�S/�.~�_ ���*D�<^��Z��HY��0��?i��?�ZA�/�6�P�����19����C?��>�W�>H7�>W�)���g��	�h3;>l�>��Q?�#�>[�O?f<{?��[?RgT>j�8�p1���ә�?3���!>5@?��?��?by?�t�>4�>��)�7�]T�����=����]
W=q	Z>g��>�(�>��>���=Ƚd\��r�>�b�=��b>���>⠥>t�>@�w>nC�<��E?a�>|7ʾ�$��!n��(��ۆ��i?��?9 7?���\��&5?�J��>�>w	�?J2�?�,?h���Q��=��);\����9����>��>`b�>�Y>�(����<��>���>��*�k}�T-�����#�?�A?t�=��ҿ*|��mn �l�һ�4�@b��]��V��Y�۾�g�B{ ��X�3�������ܽ�%��+Ⱦs[��t�#��>��H>�*>�t�=��B>��z=��0> X>��p>�l>@��-t�X�q�48�0؅��� �� >N@6>��N��w˾T�}?�7I?1�+?��C?��y>Zu>*�3����>�l���?��U>]�N��r���;�nx��Dޔ��ؾF�׾d�H����l>��H��>~3>W8�=��<a��=Bbr=/��=��c�QZ=�g�=�=sm�=���=w�>�@>�6w?X�������4Q��Z罥�:?�8�>g{�=��ƾq@?}�>>�2������yb��-?���?�T�?>�?Bti��d�>M���㎽�q�=N����=2>t��=t�2�S��>��J>���K��C����4�?��@��??�ዿТϿ5a/>
H9>%�>�eR�+2��Z�1_���Y��W"?�p;�O�ʾ:��>W��=��޾��ž\U4=�)9>'Sw=K���]�J:�=2�y��D=l�=�>�>>�=Ô��I5�=�==���=_$N>�+��x-4�*� ���,=K��=r�e>��%>��>��?*^0?�=d?�I�>��m���ξ0J���O�>rG�=�6�>�t�=�dB>U��>��7?ʷD?��K?p�>ɉ=��>�	�>�,���m��t����ZO�<P��?7Ć?�ٸ>��Q<7�A�U���a>��Ž�u?3O1?6g?S�>`D�A��5g$�*)����ND�a=x���:��J#8�2����(�=�6�>���>J�>�vl>�2>(�J>w�>��>�w�<��=�n<���<	`���=�q�z�=���'k��'wP���P�;��E��;'�;jɗ<b$�;���=h��>'>���>�s�=���8/>T�����L����=�<��3(B�_5d�qL~��	/��q6�۟B>[8X>�4���1����?8�Y>B|?>���?a>u?��>N%���վ:M��FJe��US�/��=j�>7�<��w;��W`���M��}Ҿ���>��a>�J>}ק>-�,�	9�B��<������/�_ �>�b>����b�^�\y|��o���@���m�*�{��Y?�9��G��=·Q?�M?���?���>yiȼ3�Ծ2o�=�D����<u��ۂ�����eE??D_?;��>"����4@�yh;�1Ľ�v�>¯H���O�b���?D0�%�*��뷾�ٰ>c諾�gѾn~3�ࡆ�[ŏ�5B�d4r��B�>/�O?ɲ�?�`�p��}O�����=��[�?2�g?O��>`�?(?�v��Je�?����=l�n?Ц�?#�?��>X'=eD=��>s��>A��?E��?��?�M���>�>K�<�s����R=�+a>�"u>�)�>ܨ$?`�>B��>�ae�Ý�����������7��=4D�=�A>Q�>Z
p>��J>B�:<<����#�>�Ѥ>�B�>�J>A.�>!-�>������vP2?r"+>�e�>a�*?���>���=Ͱf��ҡ<tڢ�KZ��?�tP����i�=��<=~N�
.�>^�¿Aq�?6�p>�B��4,?�^��x#5<�~<>g��>����f�>
J>g�%>~�>��>k�>r�^>�!>�7Ӿ�l>���g`!�n.C��R��Ѿ%z>�����&�ʄ�H���NI��}��_p�Gj��3���5=�C�<$J�?�v����k��)��U���~?�9�>�6?0����P���>��>ߍ>�2��"����΍�kᾊ�?���?�9c>%�>L�W?��?'�1��3��sZ���u�j&A��e���`��፿Μ��{�
�b�����_?��x?�xA?F/�<�7z>@��?��%��ԏ�e'�>a/��&;��G<=�)�>�+����`���Ӿ��þ�2�HJF>V�o?�$�?�X?{SV�iz�%w>T�8?dP+?lz?�0?_�B?�!� '?�1>���>�g�>};>?�`(??�in>�:R>�v���c��E��M��� s��|��#]���C�=�q�=�Q?��n.=s�<��<��m���PF�<�N��=�#=���=�>�t�>:�^?���>�kn>G�7?�� �v�/�w���O)?o�1=y���Q��0I���澙}>i�i?z�?��U?��?>B���D��?#>�4�>�>i4F>�^�>n�ҽ�hH�%�I=�>�V>R��=�%�	r�a�rk��s*$=�g>��>E�|>�����&>�+���~y�[kd>\R��˺�9 S���G�V�1��Xv�RD�>�K?��?���=x龙ٖ��;f�P+)?�e<?TEM?[�?���=��۾}�9���J����7��>鵫<������!��W�:����:H�s>\1���p��;b>�O���޾�`n�oI������N=���A�Z=��־�k�(*�=l�
>xB��!����X����:J?�i=�:��9IT��`���/>�<�>��>�C���w�/l@��R�� ��=��>+�9>����
EG���l?�>�OE? W_?�k�?#��\s��B������c����Ǽ��?�z�>�h?�B>y�=y���t�p�d�G���>��>�����G�A9��2���$���>�7?��>T�?��R?��
?>�`?|*?�D?�(�>�������B&?4��?��=��Խ�T�� 9�DF����>u�)?�B�ֹ�>I�?�? �&?�Q?�?~�>� ��C@��>�Y�>��W��b��L�_>��J?⚳>w=Y?�ԃ?��=>T�5� ꢾ�֩��U�=�>��2?6#?J�?>���>�����=���>�c?�0�?�o?���=.�?�:2>^��>���=k��>��>�?_XO?G�s?��J?���>F��<�6���8���Cs�-�O�6ł;
vH<��y=��54t��J����<%�;�i���N�����w�D����.��;!��>J�Q>�pž,>=��̾����oY>�.=ۣݾ|�]�ۊ��TO!�ww>�?os�>�q�;
��;)��>��>ҥ��)F?:)�>���>ۀu=�CC�}���v�<�O�>�/_?b�>�$��d����}����=�Os?�r?S9����O�b?��]?@h��=��þ{�b����g�O?<�
?4�G���>��~?f�q?V��>�e�*:n�*��Db���j�&Ѷ=]r�>LX�S�d��?�>o�7?�N�>1�b>&%�=hu۾�w��q��g?��?�?���?+*>��n�Z4��h�
���\?E7�>�U��C+?Y����䴾yk*���@����h������(���2��_�x��ޞ��z��S�=]�?θ\?��{?1'\?�	VV�?#r���k�W�b�t���sC�=#2��7�f�?�${g��(�"�羝{��֣@=@���,�,��?�@?��ƾl��>���ڼ
� �u��������N�E)>S�=o�L>SP�:��h{�����@�/?=6>�>ca?��,�G�h�fu�Ն"���(�|�>���>��
?ΰ?��<װ�#ޒ��.x��M���B�.v>|~c?��K?T�n?�K��$1�������!�/��_����B>�Z>a��>��W�����=&��\>���r�����|��	�	��=E�2?O#�>�Ŝ>�M�?1�?�z	��h���lx�e�1� f�<�*�>�i?�B�>��>e8н� ��&�>a�?�$�>?��>�o޽��� nS� +��R�>�e�>]�?E�&>�Cn��0`�R���΍�d<�=�>6�j?���������>��G?��7=h�=�I>�߽���k�Ծ���~�=�}�>%-�=*�X>��׾c���̀��Z���O)?�K?�蒾��*��4~>�$"?��>7.�>d1�?+�><qþmXE�ñ?�^?]BJ?xTA?KJ�>��=� ���<Ƚ	�&�e�,=���>)�Z>�m=F�=����r\��w�&�D=.t�=��μ�O��k�<9����J<���<��3>gۿ��I��׾��������Rb��ױ��R7������t��MŚ�iYy������N�Z��f���t�l�P��?��?B���FS���H�����������>�Gx��7���X��O�
��l���'��{����!�ׇO��$h���d�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >[C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾u1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@	�Q?�uU���Ǿ���>�>�h���J�=���QD�W�E�s�>䚹?+Ѥ?�h�>��L�͵=�b��?20u�,��
��<C��=�Fn���r��~��&;��P>Y�n=������Av#>~j�=���<}"
��0�sF=��=׬�={����҄?4.\��$f�c�/�c<��W>�T?���>Qj�=��,?&H�}Ͽ��\��a?�)�?��?;�(?�ſ���>ЊܾүM?6?]�>w�%��wt��5�=G6Ӽ0LR���|~U��9�=��>s>��,��<���M��A��=�c��Tÿ�4!�J]!�)�=BK�<@9-�d`ڽ�m^�܄��[�����t����β�=��=��A>��|>�tI>�fT>�W?KEi?=��>�>K��q����پf3μ������-�����
&��˝�>�߾����*�[[���ɾ�!=�p�=]5R�\����� �y�b�C�F�o�.?�~$>��ʾ��M�:e-<Fpʾ��������%祽/̾�1�� n�͟?��A?R����V��cR����>�W?�S�����ꬾ���=������=#�>��=��⾶3��}S�D�/?�'!?9uþ�j���5>}�"5A=V�+?G��>/X7<e�>�!?1[5���� D>-<1>5��>�c�>��>4B���>��^?x�S?����V�����>qs����k��,R=��>@0�֪����]>�7
<W���2|���y�����<��V?!��>�<*����u5����&���K=8Mx??l�>^�k?w�A?�1�<������T�W�
�ɶy=��W?'i?|u>�sr��G;S����a5?�Od?�YL>ZRi�1@�P.��m�m�?�n?Ff?�T~��A��9:�?6?y�v?�U^��s��G����V��/�>{e�>���>��9��_�>ϓ>?y#�I��S����X4�bÞ?��@���?�Q><�t�v�=49?AX�>��O��=ƾ�N��꧵���q=��>�z��`Iv�{���j,��[8?���?n�>ń��,����=�ٕ��Z�?��?����rBg<\���l��n���}�<�ͫ=�	�)D"�����7���ƾ��
�몜� ⿼祆>0Z@BV轋*�>oC8�^6��SϿ$��\о�Rq���?���>��Ƚ����G�j��Pu�3�G�9�H�	���b��>ʀ>���`Ӓ�;�{�dk;����#��>�"��"�>�WW�:޶����_|<��> ��>��>�悔�o���v�?���C�Ϳ|�����}gX?�Ɵ?Ǭ�?o�?��<69r��3����[���E?ras?gZ?�O��ua��{>���j?�Q��~U`�L�4�SBE��U>%$3?~C�>��-���|=S*>P��>�Y>�%/��Ŀ�׶��������?���?Op���>v��?�s+?
f��6��^��z�*��i�:A?2>}�����!��*=�JҒ��
?Sv0?��#+�ߐV?��W�R�U����@�F�>僾�H��Hf;6R���s�%���)&z�孥?>��?^��?�i��F���"?7y�>qڒ�~��
2>��>��^>f�q>��ON>��D71�a4Y>���?}q�?�?��楿S_�=f7p?t=�>Kd�?w�=n �>��>���2���$>}�>m�C�Đ?rCI?l,�>
D�=^cK��'1�?�G�t%O�����C��N�>�d?�J?�,b>���F��!��NĽ��-��a���?�I�:�Pv߽N5;>SP8>�Q>RpT��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	? �M��q^~�Q����6�$��=��7?�.��z>��>��=_nv������s����>�A�?rz�?���> �l?^o��B���1=qF�>��k?�q?�ls�w��զB>I�?U��,����J�{ f?�
@u@V�^?�좿��ѿ\p��w���_�վI�>��>��>��R��F>W���X�<b7���]�=�+k>��4>y˒>ab;>��=�n�=�b��
3#�y������}%9���"��3��&p�֋��J��͸��L��@�ƽ
����+��V�*��I��Ǯ�W��=n�U?uR?op?�� ?u�x�ڙ>M����;=��#�t̄=~/�>�h2? �L?\�*?�֓=����W�d��`��B��ɇ���>�rI>&��>�J�>�%�>׻N9��I>1?>��>~� >�e'=���Pa=��N>�M�>���>a|�>!C<>��>;ϴ��1��T�h��
w��̽0�?D���;�J��1���9��Ҧ��	i�=Lb.?	|>���?п[����2H?"���k)���+�Y�>{�0?�cW?�>	����T�:>0����j�F`>�+ ��l���)��%Q>jl?)e><�t>�Y3��z8�L�P�Cٯ��|>H/6?����8��u���H�yZݾ1nM>b�>0�M��u��M�~�bxh�w'{=��:?�w?�#������_�v�/Q���|Q>3#\>�=x��=HM>m]c��Fǽ��H�W:-=���=�J^>�*?e�8>��=2ӡ> ���wU�*��>0:E>�@,>>?\J&?ſ�n��:V���;�@&p>^o�>��>f}>�M��7�=ND�>�=f>���	]��s��:A���_>� |��oX��at��/�=�)��q��=��s=y@��D��)+=ؑ~?�z��ֈ�b�꾦��t^D??�3�=�3F<�"�/ �����, �?7�@�k�?�y	�C�V�U�?�9�?����"��=	o�>�>	�;8M�^�?_fƽߢ��j	���"��Z�?;�?�W/�T͋�~l�Q>EJ%?x�ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?�I>D��?��s?Tk�>�x�aY/�!5��䕌��=�][;j�>mS>Q���&hF�ؓ��h���j������a>�$=�>�0佒3��n8�=�؋�AG��^�f����>�*q>��I>)U�>� ?!`�>���>�|=r���䀾ι����K?���?-���2n��N�<Y��=(�^��&?�I4?k[�}�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��M��<��K>*4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��]S��GB�>�e!?���>�Ү=י ?Ĝ#?L�j>�(�>$aE��9��<�E�ò�>Ӣ�>�H?�~?��?�Թ��Z3�����桿��[��;N>��x?�U?�ʕ>L�������iE�#BI�����S��?�tg?]S�1?22�?�??]�A?r)f>,��Lؾ������>��!?,��A�bR&�^��o?�X?L��>-��[rս=rּ����}���?�1\?�M&?s��|$a�8�¾Xw�<F�KKW��5�;�F@���>�>����"�=7>l�=�Wm���6��a<�E�=��>���=Z07�r�����+?t�<.���(Vb=oc� @�Hg�>��b>Խ�i�V?�;��&w�h����3��F�o�>9�?J��?�!�?Zۃ��9d�K@?���?�>?��>�ٳ��:Ӿ���[i����׍	�-�>���>O���|x��Z��9��l�����������?<�>4%?}7?�E>��>Uj�����~�i���WiW�ŭ�/@�H�9�-�#�U?��	�-��<�<��ξ�&f���>� ���a�>��?y�e>6�H>�ۺ>,aB����>~�5>��c>B[�>��s>�q6>�L�=�m��c��N?$Z񾋔1��ʘ�����ן>΃?�l�>������̚*���?�L�?�'�?㑤>I�0�F%?�}uF?��?�IX��r?W�����q�������x����]�E>�*�pdw>jQ��{u�:J`�Q�ٽ��1?��%?�����'�>������m=�c�?�{(?&�)�O*Q�c�o� �V��R�<�		i�������$�(Mp������}��1���(�r�*=�*?'��?x���|�e����j��g?�32g>�#�>ƈ�>�C�>��I>�	�
2�/�]���&��悾�u�>�-{?���>L�I?;<?)xP?�kL?v��>�c�>�3��m�>S�;@�>q�>2�9?~�-?&80?�z?u+?!4c>������ؾ�
?r�?�J?�?�?^ޅ��sýui���g�.�y�~~���=%�<��׽�Eu���T=�
T>�X?E����8�����jk>#}7?���>���>����,��i�<�	�>��
?V?�>� ��|r��a��X�>n��?���=~�)>��=Yd���Ӻ�E�=�����=B4���^;��Z<+��=��=>�t��J��i��:d+�;��<Ǣ?��1?���=/�6>@���� ���P��>4�)>�O,>�C|>X@־�쉿hu��sKw��.�>QÊ?���?A>k?d=�x>�6��F������پ�K�<�>m  ?� 1?�9�?Y�.?`�*?��$>{?'�Ӱ�����C��ܰ?b!,?7��>�����ʾ��ɉ3�̝?h[?o<a�����;)�ߐ¾g�Խr�>�[/�h/~����!D��䅻�����3��?濝?fA�E�6�y�ƿ���[��a�C?�!�>Y�>}�>@�)�g�g�|%�41;>���>\R?:g�>�pO?�{?�[?c�S>=�8�V���ޙ��X?�Ω">��??Ń?� �?�y?	�>�5>�i(��4ྴ�����#3�`:���RR=��Z>�
�>Z�>K�>��=�#ǽd���P�>�̥=�'b>�$�>�n�>��>��v>?
�<IZM?�[�>*��U����(�7Ϝ��96>۫�?�rU?��J?-� >گ6�5QU�DS�\�?Vm�?�c�?��%?�&��=zD6>צ��AL��?d��>p�T>�	�=�5~>g�W=;�?�w�>8/��X�[�P�]�����G?J�L?��=�hѿ?O��Io�ݜ�UK_>��a;��=K>��)>��W>�f��=s�+��;���K��{���g�p6����>���n��=��=ϥ����=�e������0�=_�T>��ͽ:%�<*-���a�=V��V5��T"��"�=M�����о��?�:?�y�>��g?7a�>Jk�>z���ࡽ> ���-4?�Xy=��U� C�u��3B����־Y����h�����s/;�!>�f��;P>P��>�Eq>�%m=mY>�
�:�/��	�=9�=��%>8�_>��L>/�>���={�=m6w?@��������4Q��]�ֶ:?�7�>�y�=�ƾ�@?��>>�2�������b��-?s��?�T�?T�?�si�'e�>����玽cs�=����O<2>���=��2�a��>��J>����J��~���4�?��@��??�ዿ��Ͽ5a/>s�7>}�>��R���1���\�H�b�0dZ���!?3J;�"@̾�D�>.g�=�	߾��ƾ��-=�~6>�@c=,u��]\�$ޙ=�z���;=�l=�ǉ>��C>f�=�<���
�=3/I=!��=/�O>&7���n7�AJ,�8�3=0��=��b>�&>��>�?kS0?�Md?�#�>�'n�8Ͼ�5���,�>HG�=1�>1��={B>ី>��7?W�D?��K?5��>�މ=�	�>="�>��,��m��Q��ȧ��ɮ<6��?�͆?�>'!V<
�A�����l>�&,Ždx?G\1?�Y?�˞>I���޿��&���.�[�1�u��<u�g=�af�]Eռ������6��Q��=\_�>x��>�:�>A�p>-p>ӫK>��>B�>�L�<:�=�	�<g�=φżSV=ApG�,�_=����i������S�i�fq`��]{��;<��9<@��=$��>X�>��>Uޢ=����<�3>�"��K����=@V����A�Q�c��a~�C�0�"�9�m"?>\�[>v�m��Ǒ�ga?c�a>&C>*��?_�s?ʶ>�?�pо�J��N�_��NR��i�=Ӽ>�D;��{<�UGa��fN�E�о���> 3�>��>1�l>S�+��?��lx=���j<5����>���{h�p��;q��C������i�)ĺ˥D?B��2��=�0~?M�I?�֏?���>#����ؾ�d0>7��_�=| �q��D��7�?�&?�K�>�B쾎�D�_�;��콀�>�7��T�4���d�;�D)�<\a��$e�>����fF˾�1�R���ǉ���E�=i���>	�J?]ث?�r��;o���@���i�̼�
�>�\M?I˝>���>+��>�����ST��;��=X�w?Uk�?f�?0�>���=;���:�>"(	?7��?m��?��s?�p?��><��;�� >�˘��<�=;�>���=�%�=>p?`�
?c�
?�g����	�s�����+^�-��<&ҡ=���>Mo�>��r>���=�g=[y�=2\>�ڞ>��>��d>V�>aN�>�ǻ����o�@?C�=#>Mr5?an�===>���-�=G4��P��^H��
��������?�ʽ˪Ӽ#n��Mt�>�n��g��?u}�>[#�ē?�|
���O��C�=��>�D��l�>��>�8�=E��>g>�>�2z>e-�>.�B>y�Ӿ;2>O���S!�p!C�-�Q��Ҿ��{>ě���#�ֲ�R���I�=��o�Fpj��F��\i=�KB�<�3�?2�%j�#)�D��� ?���>D6?̎�l��څ>��><l�>&1��Xt��I{����nӋ?O��?��,> dG>�B?V�?����МX=��}�V7`�,��^�a���n��5��Q�z��������LS?�x?�G?��S=�]�>�m?X�=���C�$j>� �r|!�,�6�q��> ��q��`7���놾E(=�\�>���?tn?��?�'5�%$r��'>m�:?�Q1?#Ht?5�1?��;?���[%?m�3>�*?<?$5?`�.?��
?%2>��=j�û#A(=����튾�н�ʽ����%i4=T�{=Sd%9��<�=��<~R��)ڼ�0;y���-�<��9=�.�=��=(�>�]?�?�>���>��7?����7������.?�8=�_���G��I���y�[� >�%k?���?J�Z?�Xe>�PB��0@�̧>e�>�&>K�Z> M�>@���	E���=Α>��>���=hoQ� ⃾6n
�'��b�<+>���>1/|>2d��d�'>A}��/Kz���d>ŹQ��պ�2�S�L�G���1���v��a�>��K?��?��=TT�镽p:f�4)?�R<?�IM?W�?��=~�۾-�9��J�����>�>o��<�	�Sâ�# ���:����:
�s>�;���࠾
Vb>���3t޾E�n��J����&CM=0��_V=����վt6����=�!
>'����� ����x֪�-1J?4�j=�v��caU��o����>���>�߮>�:���v�@�S����5�=*��>��:>?_������~G��7�`>�>GQE?!W_?k�?�!��Fs��B�8���,c���ȼQ�?ax�>h?�B>K��=&�������d��G���>���>a��=�G��;���0��@�$�#��>R9?��>��?O�R?z�
?l�`?�*?CE?,'�>V�������@&?��?τ=9�Խ��T�c9�TF�Y�>4})?��B�v��>�?S�?	�&?܆Q?'�?�>�� ��@@����>`�>	�W��a���`>/�J?͚�>�?Y?�҃?>>�5�_T���n�=��>L�2?U8#?1�?���>�r�>��l��d$��[�>�;p?���?Q>t?<g>��?�}I>�!
?%��=�ǚ>���>ˏ�>YrD?�+s?ݯ%?���>9�9<;���#<@C��;=l]�=�z�<L4�Q����9��3��l�'��O��X<�޼򉍽�i��[L�����=���>�a>�B���&�>\�߾�̯�1��=����~ ׾\ ��:?��Y�>_>q?��?�f=_�H�>b��>3���}=?E��>CC>7��<��M�:�������v�Y>/|_?�ؐ�����'ޡ�ŏ���?><�?�ru?涬���־$�b?3�]?Vh�=�L�þ�b�/���O?��
?J�G� �>2�~?��q?���>�e�H:n�9��)Db���j��ζ=�q�>�W���d��?�>��7?�N�>��b>�(�=Yu۾�w��q��D?J�?��?���?!+*>��n�Z4�9��f���?=�?�a>m�7�7?�9p���վ�m5���n������[�Ⱦ�e��Z����#�Xt��̉����>W�)?��m?G��?�V?w�0���T�N>����a���Z��9�4���A�0�:�#�LJ5�Qݾ�h���|h>CH����F�s�?ۺ?��v��3�>*�����ߪ�����=z����3�0�<����[�=3�=2m-��"��A��-�)?���>�+�>�8A?��l��F���O���'����~�= [>�E�>��>e@�=��9�'��o���ߋ���:߼i=v>ےc?�]K?�n?�� ��+1�	l��ٓ!��*1�� ���C> >Zr�>�W��/�wR&�[y>��s�(��g���#�	���=��2?�5�>j��>�<�?	?4-	��j����x��j1�^ك<��>~i?�Z�>��>�uѽ�!��5�>&�?ǔ�>�e>����(�j�N��7/���P>�U�>Ο?��>���0�U�����|�J��ۏ=4�n?�g���<m�b��>ALc?^�>=L]^=��>�m轏��;ξ�����<">�?��>��C>�|従 2��4��9��?�	?'����"�x$�>Pf?�.?�2�>��?���>��k���=S�?�A?�6?
�@?���>j�(��.������	N_=�6v>��V>��=�G�=W�$�[�f���"�&E�<��=��}��S��_��;6
�ng�<�Av=�6>zqۿBK���پ��|�2
��߈�����e������i��V��Ndx�����v'��?V�Nc�Ϛ����l� ��?�8�?,^��� ��Щ��݉������휽>��q�����󫾒���,������ɬ��b!���O�j-i�õe�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾y1�<��?7�-?��>Ďr�1�ɿc���v¤<���?0�@�KG?�2��E˾�a>���>Ƈ�>/�[<����Kq-�y����ͱ>L/�?z�?��V>f�?��:�%G?))>��H��&U��¬=��T=٣
>��}��^c=� �>����սu2���I]>���>���<��2�[.����=�?>����a��Ԅ?�w\�;f�ء/�kT���G>��T?�*�>�#�={�,?�7H�M}Ͽ֯\�O)a?y0�?<��?��(?�׿�ٚ>��ܾ��M?FC6?\�>fb&���t����=����#��|��Y$V����=@��>/s>��,�B��xO�D�����=���r�ĿE�� �y�<�V<��J�B�
�Q����L��i���i��E��
4=�h�=��7>e$x>cV>�F>-V?�/k?Kh�>��>K�½�fs���;��ۼhዾ=�0�u���I��C�����ȕ㾷#	�CL���wþo =���=�6R�ݗ��� ���b��F�3�.? $> �ʾ?�M�ˏ-<Dpʾ~����߄�>إ��*̾�1�_!n��̟?��A?g���W�V����c}�L���X�W?�N�m��+謾@��=N�����=�$�>���=��⾆ 3��}S���(?0V?4�;{���֭n>򿟽qh�=J4?G�?�pC=n��>��?D��$��@>�M>���>	��>�E�=�X��-����?kbF?�x��O����(�>+ӾP����m=��>��+��3�k>hC�<�y���C���E�9U�<[V?~��>gW,��p�^}��l�h���_=@q?@J�>r�>N�h?,�9?d��%��ܺX�9o�Zބ=�0W?p�g?m�=
Lf�[�Ⱦ�����z6?�b?qR>�K���2羇�.�.N�S�?�l?��?�+
�h����y��B��@`7?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?p�;<��V��=�;?l\�>��O��>ƾ�z������1�q=�"�>���ev����R,�f�8?ݠ�?���>������ğ�=ڕ��Z�?F�? ����Og<����l�,n���p�<�̫=-�:I"�����7�J�ƾR�
�䪜�*ؿ�B��>:Z@oW��*�>�E8�Q6�9TϿ ���[о�Tq��?��>�Ƚ������j�WPu���G��H�����J�>��>�i������&�{�Fm;�a4����>��\�>�S�&+��i�����5< ��>}��>���>8+���ӽ�`ę?�Q��b@ο����-����X?]a�?dl�?n?H�8<�v���{�gk�o4G?�s?�Z?,b%��?]��q7� �j?R_��yU`��4�]HE��U>�"3?�B�>^�-���|=�>i��>�f>�#/�z�Ŀ�ٶ�K���Q��?��?�o���>m��?~s+?�i�8���[����*�ų+��<A?�2>���8�!�+0=�LҒ���
?(~0?�{�[.�_�G?��T��K��W!��r���ә>?��1sR�*��=�쾬R{��,>o�!��?�=�?2��?��K�Cb�h�`?X�><�I�;-2�A��>^�P>f�_>N��=�*��^�=*�ﾁ�(����>cb�?��?��?.��Q���j[>��f?���>K�?>��=U�>"� >Z��|�g���>��=��OC?&�H?V��>���= :G�9c1�YVI�ADT�&c�>zD��|�>)(a?��J?&!e>�唽^�*����$���5�2� ��;�?;%��D�&�9>U�E>]t>�mV�ܾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*��οϓ�u���������=-�>�}<>ɽʏ.>I=��Rv<r��=9��>INp>&�^>�~4>":S>��
>7���C3(�'��ѐ��-l[������������8�qM~�W6 �h���P���w�5��.���z�M��U½����=X�U?�R?�p?� ?��x��>6����Z=2w#���=�0�>�g2?��L?��*?��=_�����d�a��]@��hɇ���>hpI>�~�>�I�>�!�>��L9M�I>�,?>��>;>Ll'={��hc=��N>NL�>S��>{�>�C<>��>Fϴ��1��j�h��
w�j̽1�?~���R�J��1���9��Ӧ���h�=Gb.?|>���?пf����2H?&���z)��+���>|�0?�cW?�>!��v�T�4:>8����j�4`>�+ �}l���)��%Q>wl?��f>.u>A�3��]8���P�Rm����|>xD6?ƪ����8�y�u���H�]ݾM>���>��@�KT�������[i�ܠ{=Dj:?;x?_}�����0�u��*���?R>#M\>l�=�o�=\M>�c� �ƽ�G�1/=���=ё^>(f�>m$8>��;m%�>�V��7�:Z�>�>���>X�B?O�0?v�ּJ��ꑾ"4)�UC�>gt�>��>N�=�2����= ��>?cG>0C�8�½�r�q(���5>��/���F��e�簋=T0f�Ŀ�=��=�d��e�&�"=�pv?eʞ�-�g��l���w���6/?T@�>�2i��%ӽ
�>�s�����f�C��?��
@��?��!��mJ�f�$?�[�?Ɏ�̗�G܃>��>��i�4Ո�G�?k�X��� ����)�=��?%>�?�~꼬���7{i��J�=Y�J?�E!�Ph�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?�I>���?�s?�k�>/x��Z/��6�������m=��[;e�>^W>����pgF��ד��h����j����!�a>��$=��>pD��3���9�=��H���f�|��>�,q>��I>W�>k� ?�a�>���>�x=so���ှܸ����K?A��?���q2n�a�<?��=�^�A'?�I4?M=[�C�Ͼ8֨>g�\?���?[?�d�>���4>��.迿x}�����<j�K>P3�>NH�>���`DK>�Ծz4D�_o�>�Η>�����>ھ-���I���A�>Ae!?8��>nԮ=ۙ ?��#?x�j>�(�>=aE��9��S�E����>ʢ�>�H?�~?��?�Թ��Z3�����桿��[�x;N>��x?V?qʕ>_���생��jE�!BI�.���Y��?�tg?yS�2?;2�?�??`�A?t)f>��9ؾ������>@?����'4B��L#�\{۽?�?J�?���>o�ռ���/a�<�
�7��F ?rAT?�'?	� 'e�,�Ⱦ�]�<��*�]�E�9|�Ѽ���=�>tQ���ř=�X>��=
\�Uq(��ߝ<[P�=pv�>���=�+��_��sa,?�Ң�󙆾J��=Kfp�"�D��7�>)�M>��þ�d^?=c;�?U|�~쬿B���ed]��6�?NM�?�M�?Ȱ�J�g�q�<?���?T�?���>�P��R۾v2�ky����Gt�V>���>Di���辞إ�17������c���)n��X:?���> W?o.?:�
>��>����i� �5n��_Ӿ�CW����99���9�!�'���۾R��Fo���3ᾳ4��(e�>������>�l!?< E>r_�>R�	?��I�!>�U>x r>*iv>X�q>���>��><<ǽm�{���W?�?ž�Z�v���x_˾�?�??Ɏ�>pZ޽Z���bs����&?r�?���?�Rt>BS�`�@�E�/?��>_A��]v?&�;<��ýμ�< cJ�<������<���%Շ>Di��Zf� *o��G��)&?��"?�Ur�Cؿ�[ީ=ƌ��,�n=�M�?��(?��)�B�Q�f�o��W�
S�����6h�6j��Q�$���p��쏿�^��%����(�=q*=��*?N�?�����f!���&k��?�jdf>C�>&$�>�>�tI>��	�e�1�O^��L'�N����Q�>d[{?Џ�>ovI?��;?g8P?��L?��>T��>!t��ݗ�>�.�;�s�>��>��9?m�-?0?Rs?W�+?��b>�"�������Aؾ?��?wS?K?��?(���!Ľ����Yl���y�°���+�=J��<�mؽ�Lv�p5U=L�T>�?�����8�	���Wr>+g8?�H�>O��>؍�^���X=i�>k;
?80�>�����p�T�
��c�>�?7��L=��.>��=�`�`��1�= �<��=�}���[3�^�<���=X�=�w��9A��/3�;�<hI?�K-?�mL>�A>"qi�}7�4� ����=�M>'\p>@�>*��zS������[�m�/Wy>塚?�Ʊ?��=�ڿ=�	>.ǥ�Ŵ���rϞ��K=�W�>��?77?lg�?��F?b�?�l�=�_�`���,���ڧ��>?v!,?d��>�����ʾ��ډ3�Н?B[?�<a���;)��¾��ԽX�>�[/�l/~����D�ޅ����S��!��?쿝?�A�8�6��x�ݿ���[��[�C?8"�>7Y�>��>%�)�g�g��%�`0;>^��>XR?��>��?�A[?;�?�w�=�:H�c���Ȝ����ӽe=ck?�6�?�?��?��>��<ozF���@��5�T=���b��Ow�O�>Cv]>��5>��?�Ƨ>�M>>uɽ�(��+�o��u=�iF>��>ѕ�> ׋>(]�>��=�`B?�?;JȾ��������ݾt�z?��P?��J?�E��FsJ��S�6$�ߙ�>E�?7��?�(?�7�g��=d��=8�˾S�Ǿ���>UU�>�ѭ>�Ţ=��U=���=`A?�ϳ>�3N��q8�j�j�PSn���?�???>=��׿�r���=寽���=u��=��.�gd����=�1�<��ƾr��Nʾ���lA۾u�h'��,��^���R?%����>��u��=l�>��C�
(2>�E>X��<[��Iv�HC�{=�:������=`i<�7���=M1����o?��%?K??�D?�\l>�:�>㈊=��>0��<��)?~W>�N(�O����B��p��=�9c��e���/�M�b����=s{f�z>�=8��==9�-;8��=��<M>�=�g3={�g=�=���=�6�=�O�=��=,f�=�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>%;/>��">a&]�"�#�5셽BZ�kT�9¾8?�?�K�<���>�o=>�,��^ZžD��<8�>�2d>Ti��Q�k�{6�=�Ó��}<�Y=&�>�N�>#49;H���U=����9�<cS>S��<����x;���8�<��=�v�>�p7>���>PI?O$?�[?z�>_��Ǿ������P>$s>�e�>�"���>��>N@B?�yR?LH?�&�>k��=U1�>]�>��!��Vv�=�Ͼ���MSg=��?C�??��>m�<�Fk�y&���L������?q�;?��?g7�>�U����6Y&���.�!�����3��+=�mr��QU�D���Mm�/�㽦�=�p�>���>��>0Ty>�9>��N>��>��>7�<|p�=����4��<� ��{��=U���Z�<�vż͘���v&�O�+�Y���~�;���;��]<ơ�;01>L��>�'�=�U�>ϯ=������3>c����O�g��=����kB��Je�$�~��z4�]�?���D>��e>�E��:��"T?_W>*�K>b��?�"r?F$>R{7���Ӿ[Ҝ�R9��5�s�=�>H���D��j�`{Q��þ���>��>3�>hqm>a(�K4?�yׄ=�n⾘�5���>�_��O]5����bp�76��,���k���n��C?. �����=�J}?I?��?l�>Pq���ӾF�>>�恾���<�C�/�m�t����?��&?��>�? G��H̾����߷>yAI�$�O�Y�b�0�����̷�{��>&�����оt$3��g������čB��Lr���>�O?��?�9b��W��UO�����)��q?�|g?=�>�J?a@?�&���y��q��ey�= �n?���?(=�?E>ʎ�=���%z�>0��>�ɗ?4�?�w?�Õ��_?�y=�Nb>tˡ�l��=�A�=+��=˞>�?-f�>R��>�
V����&k��K�,�}����[ ^=lT�>��>y͓>dM>�<=��=�`>R��>>�u>?h>�ʄ>@��)(�('9?�!���>� H?�a>��<�E=7+L=:��3�'�wXP�ѱ���"�b �/s��V(:<k%ټ��>�̿�B�?��=�K���?����a��<���>`�$>_N��@ļ> �>a݂>>ܕ�>��E>9?�>�\>�FӾO>����d!��,C�T�R���Ѿr}z>�����	&����w��`BI��n��xg��j�P.��X<=�l˽<.H�?�����k��)�����U�?�[�>�6?ڌ�����>���>�Ǎ>�J��i���Yȍ�hᾣ�?D��?��\>�w�>�\?ٲ?r�A�X2*�7\��Or�k>��g�SXa��c���u���n	�wQ����^?Xx?Z??7=<�>���?j	&��n��p�{>LK1�!A@�u�]=;��>N;����o��Ծ�O��+8���Y>km?�?�? y?A,F�Br\�Vk2>:�,?#p(?V�s?6(.?�sA?�Ƚy&?�lP>�#?3?7/?�3&?W�?�C>mC>��-�[�:*���[����˽�Ƚ����B	=��7=p�t�ق)<8��<)=��+��}���&<����[��<vȺ<�ԏ=G��=���>-�]?т�>>�>!�7?����7�ذ���:/?��==o���
⊾$����*�ͩ> �j?���?<�Y?>dc>��A�ɟB��'>� �>�&> ,\>al�>z��eIF����=AH>1T>�ޥ=G�K����i�	�5���l�<!�>d��>3�|>Q�����'>������{�;d>:OQ��Z���hR��G�}'2�a$w�=�>&(L?�T?N��=I���f��j)?e1<?�L?_�?W��=3۾�'9��uJ�]����>�&�<G8	��ۢ�����V:�}�R;@hs>އ�������b>���g޾�*n�u�I���ߊT=u^��O=����վ��~�c�=Z^	>b����� � �������J?Fi=�����hU�ni��5O>�b�>��>_k>�}z�Ԑ@��_����='�>-�:>򞼖��2G�\L����>B,E?^`_?D��?�
���Br���A��x�������+����?�`�>P�	?�=>��=�&�����i�d��FF��c�>Hl�>�����G��՛�i[���"�X)�>{?*�>K�?��Q?�?� a?B�*?�?D:�>^N½�&���Q&?���?3,�=��ӽ�T���8���E��E�>O$)?ܗB�Pҗ>ς?��?��&?�VQ?f�?U,>�� ���@�K�>ؓ�>_�W� Y���[`>7gJ?�>�2Y?̓?�<>�5��Ģ�����X�=�>�2?^S#?gy?���>���>5���z��=1��>"�c?E#�?�<o?�=�q?�3>]��>G�=���>��>u ?N(N?��r?�7K?0G�>.��<�&��a5��o�v�S� �^0�;I|.<�g=
���w�����t�<���;õμ,Ls�T���@������j<�N�>�s> ����1>N�ľ�����F@>8����V������:�΢�=Q�>5�?�h�>��#��1�=1ʼ>�6�>D���L(?�?�.?'(�:&�b���ھpdL���>�B?p��=� m�������u��_h=�n?&�^?��V������l?W�U?1����Ǿ��Ҿy��C���R?�w/>�� =\��>��i?ٰ�?��>Ks��e�o���v�'v��6jh=�]�>��'�j�z2?��?I��>,Y�>��=��%�Nhx�ݠ��}?j�?j�?�Ez?�޹>Z�|���`�־zh��k�b?GT�>=���R@?n���p��ԭ�������V��@̨�q��Nƾ�.�������0��0=�b?Tse?�p?gv?�j�Q�f���K�&N��č;�wړ���aeI�YU��I���P���ھ��������,>��y���A�;*�?�2"?��*��l�>5Ѡ�����̾�>$䦾5&��p�=�[ֽ��<��<V&t�-�%��̮��i?�ȸ>��>
�@?A\��=�l�/���>�����~�E>״�>��>wZ�>�����,�h߽H
þ�pq�ֻ��	Qv>�wc?��K?d�n?w��'1�-����!���0�0K����B>�t>ŉ>��W�9���:&�^>���r����xq��Z�	�/-~=��2?*2�>�>�I�?�	?p	� p��4Vx��1����<|8�>�i?�4�>k�>,.нc� �W�>��l?/�>�	�>Lƍ��I!���z��<Ͻ���>8)�>j��>Kxn>��0�y"\�Ou���;��n�9����=?Eg?�~����`�1��>�R?�6:�+x<�+�>ˌf�&7 �b9�R3���>�)	?K��=�-9>��ƾt�pK{��{��EL)?sE?E䒾�*��O~>�"?���>�%�>�+�?�+�>5Tþ��5��?��^?$EJ?%NA?E�>�U=U���u(ȽG�&���,=D|�>�[>M!m=q�=a��cq\�@z�;�D=�ʺ=g�μ�����:<����'L<8I�<$�3>Xgۿ�=K���پz�B��,
�����,���;�����ma�����0Ex����6w'��V�c�æ����l����?�6�?b��|��즚�ꋀ�Q������>��q�MH������;���-��ۢ�>���4g!�2�O�gi��e�.�'?Ⱥ����ǿ氡��:ܾ_! ?�A ?Z�y?��{�"���8�!� >D�<�3����뾪�����ο%�����^?���>��-�����>���>	�X>:Hq>����螾~2�<l�?-�-?Ϡ�>��r��ɿO���+��<���?�@^�A?��(�m�쾘�V=2��>	?�?>*�0�;V�t󰾬X�>@5�?��?�N=H�W�e
�2ce?��;G�X�����=Sߤ=<7=����YJ>9c�>�P�UA�ݽ�a4>�Ӆ>�#�n���^�Wþ<��]>��ս������?� $���a����⒇������t?�X�>u��=$?��W�t!ڿ:�Y�#�Y?�8@��?S3? �����>�0���'B?��?�ʕ>]K�},u� �>%�b���=w8����H��M�=a��>V�=HV$��C�{t0��������=r�|����E�m
G��e�=�F'>s4@�%�='A�>�Ľs����D������=T��<�=>ã�>r�	>w�=�2N?R�|?�!�>�`�>���=?�������VM>�y��(�Ӿ����������x�F��2������'���!=��e�=�7R������� ��ub��F���.?�%>�$˾U�M��,<�Cʾ����܇�O2��5�˾{�1�?n����?�A?	˅�ַV�r����n~����W?��V������_<�='E�� �=[�>�W�=����3��]S��u0?J\?����z_���)*>�� �s�=l�+?#�?-QZ<�&�>(M%?`�*�%9�V`[>B�3>1ף>���>�<	>���T۽ы?ڈT?D��O����ې>�b���z�~a=�/>*:5��꼼�[>qz�<���8V�nL���\�<x(W?i��>��)���(a��0��5Y==��x?��?.�>j{k?��B?wפ<�g��u�S���aw=��W?%*i?��>�����	о{���%�5?ףe?e�N>vbh���=�.�GU��$?�n?._?�|��w}�t��M���n6?��v?s^�vs�����Y�V�b=�>�[�>���>��9��k�>�>?�#��G�� ���wY4�%Þ?��@���?��;<��X��=�;?g\�>�O��>ƾ�z������.�q=�"�>����ev�����Q,�h�8?ޠ�?���>��������=�����X�?$�?Py����z<��d	l��g�����<��=*���R%���d8�@ǾW�
�����E���Ȇ>6K@��x��>��9��6�T'Ͽ6)��O�Ͼm�o�q�?�b�>��˽󨣾=sj���t��G��FH�2���E�>k�>!T_�눋�!ׁ�ќ:�:�ݼ���>c#*��[>7rs���ɾ�f���{�v�>N��>�ä>Τļ�ǭ�9��?����Ͽ쑛�P
�tO@?�h�?h��?�?�<YX{������/<�X?Ws}?o�d?���i􅾑6¼�j?�_��TU`�ߎ4�jHE�U>�"3?�B�>P�-��|=�>x��>�f>�#/�s�Ŀ�ٶ�D���T��?׉�?�o�3��>m��?�s+?�i�8���[����*�S�+��<A?�2>8���X�!�A0=�GҒ�̼
?_~0?�z�M.�2�_?ta�m�p��-��G˽s�>��.�'�\�/k�!���qe��+��\z��ح?eo�?�;�?�����"��}%?H�>N����Ǿ�c�<�ѧ>�ɵ>GzP>�D`���v>��^�:���>�s�?K�??�?�B��0馿�\>��}?�Q�>#�?3Q>s ?�>�ʾb�=p��>V췽����@� ?ɳA?�?�!H>��k�X�*��X-��`~���Y���;� A�>9-O?�4?�b�>^k �|r{��� ���><3|�� �,=�� ��4�C�
����=/4M>-7g>��ȽN[����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Fa~�"���7���=��7?�0���z>���>^�=�nv�໪�K�s����>�B�?�{�?��>�l?��o�W�B���1=M�>��k?�s?�Go���P�B>��?/�������K��f?�
@~u@U�^? ��п�w��s���=�#@u>~��=͔=_����w>�S.>���=�.>kU>�E�>�>C>L�F>	3�=?59>�����%�nG��bߢ�:�B��ܾ�����E⌾�׽�3��žO���)�$X�����c�ܽf+e�+�#�"~#>j�g?�l[?��?��%?4Z%���*>ל�3ɽo��<6�u>��>#�9?[�Q?O��>Q|�<#f����g����芭������>֨a>,� ?q ?@�>M���6�>:��>9&�>)v�=��%���=L��<��N>�j>Y�
?.�?�@<>n�>�δ��1���h�w��̽;�?����J��1��89��O���]d�=a.?Ny>h���>п�����2H?�����'�h�+�_�>u�0?�bW?-�>S����T��7>`��O�j�>]>�* �i�l��)�e%Q>�k?�Gf>Ot>�S3��[8��yP������Y{>He6?�ζ�S(;�S�u��vH��9ݾIL>�,�>��S��_��ۖ�:�~�*�h�|y=U�:?�y?[-���d��v�53���KQ>��[>�=��=�'M>e�g�3�ƽ �H�7�*=���=%D^>�W?d�+>j��=ݣ>�_���BP�P��>�~B>�,>l@?C'%?W��T㗽K���H�-�w>�M�>��>�T>sZJ�/�=~k�>��a>�=����\���?�#|W>�~�wz_�IGu��x=�4��y��=�
�=A� �P=��%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>yx��Z�������u���#=O��>�8H?�V����O�e>��v
?�?�^�੤���ȿ6|v����>W�?���?g�m��A���@����>:��?�gY?toi>�g۾2`Z����>ӻ@?�R?
�>�9���'���?�޶?֯�?B�R>"�?��v?�y�>���/������Ɋ���<4�J�N�t>�l�=�CҾ�E��ܓ�����?/j�/����G>?=8�>7Խ������=�缬3��=�	��9�>Ҝ�>�	�>�R�>`?Aк>���>b4!:g���-(���釾!L?5�?Vg���g�2��<W�=��O��?�N,?�b����Ⱦ�=�>W�_??�?Q�U?��>����̜������P�����<��J>�E�>jK�>l=���J>o�Ҿ�6��>W�>�ҍ�6�ݾ�]y�����+�>Il"?�>�[�= �'?kM?���>^	?�"S���y�=�5�U��>ȻT>J(/?Z�u?d6? ��t�I�"�������o>K/y?E�!?�@b>�uy�<�m��������m�Ӽ�v?	)?>5�O?�)�?�Ȁ?�H*?�Y�>s(�̐Ͼ�d;��j>��!?Q��A�HG&��!��o?6X?���>l%����սy"׼���V���( ?�1\?MJ&?����)a���¾�K�<�L"��YV�/=�;�1C��>'�>8���4��=>j��=�Bm�VC6�_^f<WN�=v{�>��=�!7��w����2?\��=nrr����=6�b�1�X�̳�>B����־ߨ7?�鲾��� ����!��H�e��Ӎ?�?�>�?�@�=�$X�e�1?V��?2��>!F�>Lɽw�*��(�����d��Җ�K��>ˏ>>G��a���괿2���M'��⻂�����z?���>��?x��>z>w�>�)���/������-�V���&�,m7�b_2��[��=���X��u�������Bx���>�����>o?��>%�>�l�>��<�c�>Fx>�u�>	0�>��$>��= �	=��M�N2̽�KR?3����'���辉��� 3B?�qd?�1�>i�������~�?���?As�?�<v>�~h��,+��m?r=�>_��eq
?<R:=�F�@�<3V�����2����Z��>�F׽� :��M�kmf�Aj
?�/?�	����̾F>׽�|��.�={!�?Ȱ*?�z#�ٚF�Y�b��MN�� R�u^=��ɀ�m����p)�i1q��u��H=��1)��@�.���5=��"?�{o?pG�����7���5@�?�<�1d�>]��>�'�>(�?T��>����c�2�xZ�j�(�=0��{5�>\݁?���>�I?�R<?��P?%M?�ێ>a~�>e��4��>��"<֟�>BQ�>�9?l.?�/?6�?�*?)�`>�l��Z���L�پ&�?�!?7�??�f?����,��u|����_��z�t���H�=���<Hٽ��x��g=��Y>�?��v�7�+.��+ap>%�7?���>Ն�>�����(��-.=ڼ�>+?���>B���=r������>l�?V��k�=^J)>9��=^x���N�w3�=�}Ҽ�b�=����?� hQ<�Ҿ=w�=L�u�Ɓ9��/;��;"��<�u�>��?�Њ>(N�>�J���� �f���=�mX>*�R>S�>B<پ\���(���g�^�x>�W�?(U�?f=� �=�!�=EX����-��t���~�<ӧ?-P#?j\T?���?R�=?i�#?�U>�1�hL���h��z��Ʈ?�,?⍑>�����ʾ��3�W�?\W?�<a����d<)�i�¾�!սȕ>_/��.~����iD�P����������<��?W��?�@A�W�6�H}���:Q���C?�4�>t_�>#�>�)�x�g�p&�h;>L��>#R?
�>+�O?]K{?��[?g.W>�8�V���~���B3C�"t#>T@?��?Iݎ?�y?0y�>�
>�)*������\� �����V��6tL=��X><��>�
�>
�>���=H]ʽ2H���?��U�=�b>�
�>��>Q�>��y>���<M[Q?�U�>��ѾO�վ�{Ҿ�V��ڔ>��5?\��?C
?H ��SC��2J���¾
�?Y˶?9�?}�%?�ڝ;꺭=m����|���7R�C�>���>��>��s�^2޺{�,>�v�>���>*�n��L���e�\��	?�W\?Y�=��u\�����8T��Ǩ�=��������/�=������/B���%�a���H@���*���q��:�����r���?s<=�>�t�=^Yg��0R=C�߻��=�����;����C{<F6v�W���)����[̽�݃=8OR�� ž��}?�K?�L/?��G?�C{>I5>�=����>�&.��.?$G^>A��谾�+B�1}������eھ�	ܾYe��S��C��=*��&�>{�;>ٞ�=b�='�>��W={��=��C�=���=8��=�Z�=]��=k�#>�,>�r?�eR��V��m1�8������>��>�,I=�U����?�b<�琿�t����D݊?��?B��?��?*ώ�O�>�&z��*��v��=�_d�5�޽���>�k��A�>��>|��FŞ�C <���?��@�X?Na���8Կ��>2>�� >u�Q�4g1��,U���V�ΐ]�D5#?�8��Ҿ�%�>{L�=��ݾ�Ǿy�=}�.>��X=#D��[�V�=���1�d=�r=D�>/TG>-��=WҪ����=�[3=mu�='O> ��i�O�z�&�=�=�Ƿ=(�b>W�!>��>�?mu0?md?���>qym�ҽξH������>Sh�=���>�ņ=��B>�ĸ>��7?N{D?۠K?�A�>ɵ�=��>�d�>�,��m�s徦}�����<��?�׆?�M�>,Q<��A���0'>�kŽ�<?:1?�?���>>'���nLl��ke� 8=�>3���K���>�>0�^>���=Z�D>J�]=-��>2��>�	{>�_=>\:;>0<>�|�>C>u�:;���;_
A��ov<�bc=
�)>��;Wc�o�E�g_Ľ2B�=&ˤ=�{�<�۫=�7���<��L�b>&��>�E\>p�>��<��ɾ��J>+����K[�U7=׸ξ\W=�Z�u��fu��q1��x4�.�,>�j3>r͡��֋�R�?��>x�2>�?v�m?�6:�ՠ�9_̾������@�e��� W�=%��=k�\���N�JDq���j������>��>��>+�l>V,��"?�
�w= �Mi5��	�>�������wG��7q�>>��|��i�IRݺ��D?B�����=~?p�I?�ޏ?n��>0i���rؾt80>�C���<=] �d�p�z`����?� '?P|�>.,쾏�D���˾����bո>t�G�ƻO�>.��-�0�F�5�Է�3D�>�r����о�/3�_���/폿6�B���r�w��>�ZO?���?��^�� ���DN��_������?�:f?�=�>��?�??�������y��ι=?5o?���?�;�?$T>J��=HYB���>�?Eǘ?僆?�b?x���>�D�=�ȓ>��w���?>gˋ>��;aa=|@�>�?��?]�㽡�$���
�����z��_��=���=
~�>���>:��=� >�֙=ҁ�=�ܜ>?:�>[B>�>>���>vU�>����I��s�?e�~<Ԫ�>?�I?�>�w�>(ڝ���W�6:��Zv+����9�=�yl(�����x�����<Ƚ�4�>�ͻ��O�? �B>�����?FJ���5��P�=��>��d����>�)7>/��=Ց�>U�_>d5�=��>��=��Ѿ} >ҍ�~a ���B��R�>�Ѿ��x>Q)�� 2&�'��x����
K�~Y��3��j�W��a=���<���?� �/k�	(��� ��	?���>F6?i��ʦ}�	w>:��>s>�����g�������*�&��?&��?W|>2 �>�h?��?�n���$ɽ�f�6�u�='�Ac�Mc�y����x���I�DZ���<?"s?U�p?�7�=�9�>��?Ȋ+��
���ݽ�Tq���Tq�=��>z����E!*�d����=vS�>�4�?[�?��?����=����=��?UK?
��?��;?w� ?�D[��C�>[Z~>$A?.?�H?)�T?G?Ƥ�<#2Y=�Q>�=@��g�sJݽ��i�=���=J��݆\�Dq���Ҽ	<#Y4>�XC�*���#,=ld=��=���=�!>��>�]?���>���>nc7?�����7��?��%/?!�9=<��RӋ�&6��g��A�>�Ak?T�?kmZ?�~e>��A��CC�h>�*�>
'>
�\>��>I���F� �=TN>�f>Ju�=(�P�҂�x�	��h�����<��>���>V~}>{���+�(>�&��Q���ql>�W�2��}GS�(gH���2�W�{�8�>�SK?q�?�,�=)
澹���e�t(?�<?pBL?�H?՝=*sݾ�z9�-�K�Z ����>XB�<�Y	�)}��x��h�;�p�-�<gs>�՟�	ˠ��@b>���Y`޾g�n�QJ����>�L=[~�R�V=��U�վ�� ��=�(
>���� ����Ӫ�H-J?��j=�|���mU�>_���>�ɘ>���>��:��Cw���@�૬�)>�=!��>� ;>V�����qG��5�P|�>��D?_?h\�?-r����r���B�}������<]¼�?��>?�?�*B>��=�������%�d�[�F�\��>�T�>���ȖG�4��� ��ϸ$��D�>1?�2>�P?2gR?��
?v�`?̭)?��?8�>[Q������t\&?�I�?��v=tS̽)X�H17���E�9��>�t'?��A�6#�>O�?��?�(?@iO?[X?N>�y���A�z�>_}�>�W� ����+b>��K?Tm�>ԋ[?���?�2>|h6��С�����.�=wi>�.?�)#?��?M��>}��>G���t�=Þ�>�c?�0�?�o?ރ�=9�?�:2>F��>@��=���>i��>�?PXO?;�s?��J?��>���<�7���8��@Ds�D�O��ʂ;�vH<K�y=���T3t�1K�S��<�;jg��|I��I��w�D�����\��;u��>�+�>�Ѿ��ӻ�Տ�]���P1{>���=	���
���nv��x�3�q7b>m�?|��>~ǽ� >���>��>5���$?���>�9?�ۮ=UDi��4����'��)�>t@?� 1>?s�Q��.�����=�܀?�m?�Hp����I�b?��]?=h�=��þg�b�ǉ�.�O?�
?��G���>��~?v�q?j��>��e��9n����Cb�{�j�yѶ=0r�>JX�K�d��?�>��7?�N�>�b>%�=�u۾"�w��q��k?y�?��?���?|+*><�n�;4࿎����C��wj^?H�>뚤��L%?	���s�;K����Ց�ÿ��\�� *��IV�������(��	��@ʽ ��=�6?}�q?D�s?E�^?���b��U`�[0��kT�����L�B�C��oC�*B���k����4񾐵��"�T=�k��hOQ��*�?
?� �v�>w���/��W+��zE<�o���F!=g�f>��޼�u>=[�m=����{:V�����R?̎>��2>��Z?	b�����0�1�!l�U�<�,��>'?��?�D�>�O�xQ����D>'~��[��r�@�r1v>Ozc?�K?��n?�g�s)1�9���ɖ!���/�!d���B>�Z>���>�W�����<&��V>���r�\���w����	���~=4�2?�.�>8��>XL�?t?"y	�Jq��anx���1��x�<W-�>xi?B:�>��>�нm� ��T�>ɪp?��>�>�y�T��Q9^�q�n��#�>��>5e�>z�4>~Y�(U��Ǔ�Y�����/�p��=��Y?� �������>9`?������;L�G>��۽Y��|l��,�Y��=d��>�=b,>9Zվ2e��
���_��EU)?E?����*�?~>-	"?ao�>�?�>""�?��>�þnG����?9�^?�JJ?�OA?b�>��=�3��}�ǽ��&��,=Ph�>� [>�m=�&�=�D�*$\��i��xE=�"�=��Ӽ5��B
<I�� 9U<8S�<�3>Amۿ�BK���پ����>
��爾	���d�����
b��B��*Xx����'��V�V7c�������l����?�=�?���>0��������~���d��>5�q�7���󫾢��7)��Ж�����6d!���O�u&i�4�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >ZC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾y1�<��?7�-?��>Ŏr�1�ɿc���x¤<���?0�@��A?I� ����=��>n-�>���=�H�)�����0��>���?��?�>��:�C����|U?�9�<��L�SR�<2`>��g� $���cG�@V�>3��>\�=�G�	\����<Wb(>,�<?␼��#��5սg�o>��ǻ�o"�
Մ?3v\�5f���/��Q���M>��T?�1�>�=�=��,?9H�f}ϿU�\�(-a?�0�?���?��(?�տ��ښ>��ܾ��M?	B6?)��>`&��t�:��=� ἺL����㾦V����=З�>�e>A�,�	���lO�.[�����=\���ƿ�$�"|��r=�x�:��W����:���Z����	�o��#�r�g=�^�=��O>��>V�W>xkY>��W?`ok?��>�>��[Ɉ�@�ξ����D���~�x����%�	���7j�"�޾7C	�����_���Ⱦ�=��
�=y6R�B���O� �
�b�!�F���.?s$>��ʾs�M�.<�jʾ輪��Մ�Qޥ��+̾��1�V"n��̟?��A?������V����Z9��w��_�W?>P�ݼ�E���=����>�=D$�>�z�=Y��d3��}S��8-?�"?�w������38>�Q�m��=�/?��>���;狛>�t?@�R�Q��Z�=Dc�=�{�>���>��>����
�%?\�^?���w��� N>Ҿ�M}�-�`=#�="X5������<a>R��ͭ�;c˽Y!��滯W?nΌ>I�)�����a��^� ���;=�x??���>;\k?��B?*��<�>���AS�]�
�#�s=�!W?��h?��>b����Ͼ�����5?�pe?7�O>�e�(+��\.�oI���?�)n?�d?ῒ�T�}�t�����6?��v?�p^�rs��5��d�V��;�>�_�>���>��9�^j�>ߐ>?�#��G�������X4��?~�@C��?��;<�%�I��=w<?�\�>�O�*=ƾ!r��2���C�q=�!�>ފ���bv�}��GV,�8�8?��?���>ʒ�����2��=J�W�?h�?軪���c<���,l�UD��k
�<�9�=���W*!�\�� �7���ƾH�
����������><Q@-��9�>m8��4�cAϿ����_оd�p�:�?Ջ�>ϡȽ�����j��,u�;�G�)�H�����1w�>S���{���|��������O�
w�6�>��2���>P=���DK��^U��ۋ>z�?є>B��l�D����?wd�s�˿�"��W�n��22?�:�?X��?1L�>`A�>Ml�<ƒ�kJ)���?�t|?bF?����=ȾV7B>٠j?����2`�"�4���D�\�T>�c3?ԅ�>�a-��{=#�>��>eS> /�]�Ŀ[ȶ�O��c�?vc�?'꾦��>d��?��+?�o�m��骾��*�Sws��A?`�1>|v���s!�v�<�q.��4
?6�/?��p,�]�_?,�a�M�p���-���ƽ�ۡ>	�0�f\�jN������Xe�
���@y����?M^�?i�?��� #�k6%?�>_����8Ǿ��<���>�(�>*N>H_���u>����:�i	>���?�~�?Sj?���� ����U>
�}?���>�a�?���=tG�>D��=����G1��D�%>5t�=��C��?S�I?��>]l�=�iE�Y�0�:dE�A�P�ȑ��C���>	�a?qJN?ݙc>�g��%e�!�;�ԽF�5�(�����E�
�6��S޽O6>\w7>$>D?L�Q�־��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*��ſڔ���lN���3�ӽ|>��>��>�Q𼌳�>�f����n�=�>��==9�>$�>a`>�/<3Eq�K&#��]���#����2��Y��a^�,ao��L���C�܀��,���`v�>U�eE6�߽j�hE�1���A��=h�U?�
R?�p?!� ?��x��>����&=~z#��Ȅ=�1�>�h2?��L?��*?�Г=ҥ����d��_���<����y�>�^I>.z�>�K�>�#�>�3�9��I>~?>w�>� >��'=�ֺ�A=��N>�O�>}��>ni�>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ӧ���h�=Hb.?|>���?пf����2H?&���z)���+���>}�0?�cW?!�>!��w�T�3:>:����j�6`>�+ �l���)��%Q>wl?x�f>�8u>H�3�(b8���P����ɀ|>�26?�㶾�A9��u�ձH��jݾ4M>D��>��F�h�R�������i��|=�z:?�?o5��Lް��u�{L���<R>�&\>�-=�0�=�OM>%:c���ƽ�$H�=�-=�c�=��^>�i?t_d<�}=�A�>�����먾��K>���=B{��}`?
�=?A}�=eoz��&¾$m�:��>��\>܏�Z]�>r+��>3|�>_M>uo+��<h�,��s@�/�^>�"J�ZB���p��}�&>�v$=��=u�<H=�d۽�ý�~?���(䈿��e���lD?R+?` �=�F<��"�E ���H��G�?r�@m�?��	�ޢV�@�?�@�?��L��=}�>׫>�ξ�L��?��Ž6Ǣ�ɔ	�3)#�iS�?��?��/�Yʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�}�#=Q��>�8H?�V����O�g>��v
?�?�^�੤���ȿ4|v����>W�?���?g�m��A���@����>;��?�gY?woi>�g۾>`Z����>ѻ@?�R?�>�9���'���?�޶?֯�?kI>3��?��s?�j�>�x��Y/�U3��%����Z=�Z;M_�>0E>t����eF�kؓ�_i��5�j������a>9o$=��>[1�^'��HO�=�݋��M��S�f�a��>�q>��I>RP�>%� ?�]�>X��>j=v���〾�����K?���?.���2n��N�<��=9�^��&?yI4?�j[�z�Ͼ�ը>�\?k?�[?d�>/��D>��<迿)~��\��<i�K>4�>�H�>�$���FK>��Ծ�4D�Np�>�ϗ>4����?ھ�,��*W��;B�>�e!?���>Ү=י ?֚#?�j>�*�>�aE��9����E���>���>�I?��~?|�?8ӹ�L[3�����塿ɒ[�G4N>��x?$V?�ɕ>Y���7����E�FI���h��?lrg?�D彍?�1�?�??E�A?�,f>���Q	ؾ����>f�.?�e���1�f�ľ,ER���S>�>�P�>�����p�>��>������鸂>��z?��3?�TP��h��t�=ņ=�5�<�M=����t}*����=JQ>����儼
a>`����&�i�k~=>�=��>kV>�*�kb����*?r=�1����3��Q\�z&>�Rܭ>���>f����<P?p�@��7u�.ԫ�F������U�?��?e\�?�qr�j�b�� :?ỷ?�b?-��>���s�޾����Hz���f�:$�<�>���>�����8X��b|��~A��'<ͽ��C���!?#�>�k?�?�!>���>��S�F��m��Mf�iPi�i�1���2�]1D���;�����vCE�850���ʾJ�Z� 9�>c��=��>,�?�9>�R>H/�>֭���q>��1>GY>���>i��>��8>-)�=c]����9�&aS?U���mC������'�>?r�X?�9?���#�}�B�&���?y��?"�? V�>E<f�"��g?7J�>��0��Y?dy��6e�H\6>��ľ�<�.> g=�&`>�Mb��\�	f�%��|,?��?<�!��ĸ���3>����i�n=�L�?}�(?�)���Q��o���W��S��i�'#h��a��V�$���p��ꏿ�[���$��0�(��*=�*?��?�����)��A&k��?��hf>I��>�+�>��>DsI>��	���1�w�]�7J'�{����I�><\{?΋�>8�I?|�;?�vP?�cL?���>�U�>t8��f�>Vs�;���>�
�>F�9?��-?40?y?Vr+?�>c>����������ؾy?��?iI?K?X�?ʅ�Beý�#��Zh�ʨy�Qg��p+�=��<s�׽��t�aU=��S>�s?&��q�8�����j>t�6?���>�I�>�ᐾ��~��{�<�i�>~C
?�l�>������q���s�>/т?S~��A=� *>���=�Ƈ�mF���=L	����=��}�P�>��/"<�t�=��=��x�v]88��:O��;2Q�<Kf?$�!?�a>�=>�q\�G�������>��Z>�@>�V
>weܾ��������g�Go>j��?.9�?5X�=���=4�>0�{�c��
��(���s =���>#"?�<L?Ԡ�?�??�q#?c(�=#e%��S���Z��;ۥ�i�?� ,?��>����ʾ$�3�ƞ?-Z?�:a�/���5)�/�¾Hս}�>+[/�*+~�e���D�tz��z��1f����?H��??A���6�4�边���Z��^�C?e�>uS�>O�>�)�K�g�4&�1 ;>lz�>=R?n�>��?�a6?~GN?Vg�x�2�]t����������ڂ>�?*?_
�?Z,�?b�U?���>���>�"/�:D¾EվGv���Y_=Zׅ��ݗ<��>�H�>��>U1�>Nj>|9���p��b�*���3><B�>o;x>�5�=x��>b?Ep����J?y��>
�J�:������]����>���?�P�?*O?F�S��K/���_��Ҿr��>e��?��?��2?����ɠ=�=�ZY�m���*�>؞>b�>�Z=SW=J\3>�;?���>�p��cH���l�����?p�B?$F�=/�Ϳ��v���N�����nq="z����`=^�z.�An|��O���|;�,��rD�����C���׭��Y�kO���#	?Rf=tn�>��w=L�<�_>=�g˽�/+=o!̼i׋��5��FN=��Y���EZ�����c���/�=���=ڟ�>��?A[!?��?�aP?>́>��d>��=Y�?��t�}�>���xV�G.U�𜖾����9��c������eRQ��퟾Ii�=�H#���6=&P>��B>2	=5ǫ>/�=�p�=|�=�S>�2>��=>Sn>�>?�.>�:>�6w?Z�������4Q��Z罅�:?�8�>�z�=��ƾ~@?��>>�2�������b��-?���?�T�?�?�si��d�>@���㎽�q�=�����=2>���=��2���>�J>���K��⁳�{4�?��@��??�ዿɢϿ�a/>628>��>�R�k>1�A�\��	c�d�Z��Z!?�M;�Ú˾���>k��=_�޾�uƾa1=��6>��^=U���	\��C�=��z��H;=�Aj=�ʉ>VCD>�'�=r���:Q�="oH=�o�= �O>�F����5�0,��1=�(�=�c>E�%>���>�?l90?�Kd?�ٹ>�n�CFϾg���!�>C�=1�>XF�=�;C>d��>��7?1�D?��K?K��>�a�=	�>>�>J�,�c�m���V�����<��?ĸ�?�p�>;�I<�_A��v��.>�AYŽJ9?I1?@t?O��>�\��$࿐�%��.����^/8<�;=�p�^sc�k��ou�bI����=l��>.x�>�7�>�v>��;>�J>O�>$�>�[=��y=:Ļ���<7����U�=M?����<˵ܼ����A�@�=�����uT;<�
:��<�U5<�s�=q]�>�>ϥ�>�=H�����B>"0��[�D��=�]��LD��Je��aw��p9��r�m1->{�K>'5�������%?
�v>�9>�Ծ?�;l?�ܮ=G$��׾F���N�e�GPl�7��=��>��*�I�9��^���P��`�D0�>߸�>p�>B�k>�1+���>��<�=�m���4����>���Dk)�-/�
�p��f������~h�=��ʹC?���X5�=�
~?�|J?�|�?���>H&���پ��->������
=�D�eNq�o�����?��%?/N�>A�,4E��H̾_���޷>�@I�2�O���V�0�9��0ͷ�4��>������оk$3��g�������B��Lr�[��>&�O?��?[:b��W��IUO����g(���q?�|g?.�>�J?�@? &��z�r���v�=�n?˳�?R=�?{>�>�=�u��3�>�/	?���?���?xs?'V?�J�>XQ�;l� >�"��k��=&�>g,�=ϙ�=�d?&�
?�
?)y��O�	�&����_3^���<��=�}�>֑�>��r>�<�=c�g=^բ=_\>��>l��>��d>��>�Q�>��˾�!��_/?^W�=��>�2E?��q>*�n=��D��:�ɽplJ��M$��\ѽ#9��*���䭺`7�=�	��^�>�滿�ϟ?�Z>����g?��G���/c>�:>��Խ#C�>77L>�y>��>>Ԩ>�==>�t�>��:>=FӾe~>����d!��,C�_�R���Ѿ�|z>�-&�s���u��-BI��n��g�1j�[.���<=��Խ<H�?������k��)�����N�?�[�>�6?�ڌ�
����>t��>]Ǎ>]J��/���Zȍ�=hᾒ�?*��?�;c>��>F�W?�?�1�<3�vZ�,�u�n(A�'e�Q�`��፿�����
�u��-�_?�x?+yA?�R�<$:z>S��?��%�Vӏ��)�>�/�&';��?<=u+�>&*��<�`���Ӿ~�þ�7��HF>��o?;%�?|Y?STV���n�f'>��:?��1?�Jt?��1?n�;?�m���$?�53>�;?"W?�;5?��.?��
?��1>���=����	'=e4��z�Foѽ�xʽ<�x4=�#|=��Ӹ��<�o=ɋ�<�yټ��;Ha��OB�<�?:= �=�=�=��>�]?�.�>�@�>��7?�(�Q�7��{���
/?r8=o���b��Z����A�A>��j?��?�Z?��d>B�f$B�̃>C��>�[%>4(\>П�>9��ٷE���=��>�>H�=b!R�c��+8
�)���T�<�@>��>��z>�ꍽ�R(>����0{���b>5iS�0��|HR��AG�1�%�t�8��>��K??/d�=&�ˣ���f�K�)?F<?�M?��?z�=.ܾR�9��=J���Ϟ>��<�9���������:��4;ڲv>@5��	ˠ��@b>���Y`޾g�n�QJ����>�L=[~�R�V=��U�վ�� ��=�(
>���� ����Ӫ�H-J?��j=�|���mU�>_���>�ɘ>���>��:��Cw���@�૬�)>�=!��>� ;>V�����qG��5�P|�>��D?_?h\�?-r����r���B�}������<]¼�?��>?�?�*B>��=�������%�d�[�F�\��>�T�>���ȖG�4��� ��ϸ$��D�>1?�2>�P?2gR?��
?v�`?̭)?��?8�>[Q������t\&?�I�?��v=tS̽)X�H17���E�9��>�t'?��A�6#�>O�?��?�(?@iO?[X?N>�y���A�z�>_}�>�W� ����+b>��K?Tm�>ԋ[?���?�2>|h6��С�����.�=wi>�.?�)#?��?M��>}��>G���t�=Þ�>�c?�0�?�o?ރ�=9�?�:2>F��>@��=���>i��>�?PXO?;�s?��J?��>���<�7���8��@Ds�D�O��ʂ;�vH<K�y=���T3t�1K�S��<�;jg��|I��I��w�D�����\��;u��>�+�>�Ѿ��ӻ�Տ�]���P1{>���=	���
���nv��x�3�q7b>m�?|��>~ǽ� >���>��>5���$?���>�9?�ۮ=UDi��4����'��)�>t@?� 1>?s�Q��.�����=�܀?�m?�Hp����I�b?��]?=h�=��þg�b�ǉ�.�O?�
?��G���>��~?v�q?j��>��e��9n����Cb�{�j�yѶ=0r�>JX�K�d��?�>��7?�N�>�b>%�=�u۾"�w��q��k?y�?��?���?|+*><�n�;4࿎����C��wj^?H�>뚤��L%?	���s�;K����Ց�ÿ��\�� *��IV�������(��	��@ʽ ��=�6?}�q?D�s?E�^?���b��U`�[0��kT�����L�B�C��oC�*B���k����4񾐵��"�T=�k��hOQ��*�?
?� �v�>w���/��W+��zE<�o���F!=g�f>��޼�u>=[�m=����{:V�����R?̎>��2>��Z?	b�����0�1�!l�U�<�,��>'?��?�D�>�O�xQ����D>'~��[��r�@�r1v>Ozc?�K?��n?�g�s)1�9���ɖ!���/�!d���B>�Z>���>�W�����<&��V>���r�\���w����	���~=4�2?�.�>8��>XL�?t?"y	�Jq��anx���1��x�<W-�>xi?B:�>��>�нm� ��T�>ɪp?��>�>�y�T��Q9^�q�n��#�>��>5e�>z�4>~Y�(U��Ǔ�Y�����/�p��=��Y?� �������>9`?������;L�G>��۽Y��|l��,�Y��=d��>�=b,>9Zվ2e��
���_��EU)?E?����*�?~>-	"?ao�>�?�>""�?��>�þnG����?9�^?�JJ?�OA?b�>��=�3��}�ǽ��&��,=Ph�>� [>�m=�&�=�D�*$\��i��xE=�"�=��Ӽ5��B
<I�� 9U<8S�<�3>Amۿ�BK���پ����>
��爾	���d�����
b��B��*Xx����'��V�V7c�������l����?�=�?���>0��������~���d��>5�q�7���󫾢��7)��Ж�����6d!���O�u&i�4�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >ZC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾y1�<��?7�-?��>Ŏr�1�ɿc���x¤<���?0�@��A?I� ����=��>n-�>���=�H�)�����0��>���?��?�>��:�C����|U?�9�<��L�SR�<2`>��g� $���cG�@V�>3��>\�=�G�	\����<Wb(>,�<?␼��#��5սg�o>��ǻ�o"�
Մ?3v\�5f���/��Q���M>��T?�1�>�=�=��,?9H�f}ϿU�\�(-a?�0�?���?��(?�տ��ښ>��ܾ��M?	B6?)��>`&��t�:��=� ἺL����㾦V����=З�>�e>A�,�	���lO�.[�����=\���ƿ�$�"|��r=�x�:��W����:���Z����	�o��#�r�g=�^�=��O>��>V�W>xkY>��W?`ok?��>�>��[Ɉ�@�ξ����D���~�x����%�	���7j�"�޾7C	�����_���Ⱦ�=��
�=y6R�B���O� �
�b�!�F���.?s$>��ʾs�M�.<�jʾ輪��Մ�Qޥ��+̾��1�V"n��̟?��A?������V����Z9��w��_�W?>P�ݼ�E���=����>�=D$�>�z�=Y��d3��}S��8-?�"?�w������38>�Q�m��=�/?��>���;狛>�t?@�R�Q��Z�=Dc�=�{�>���>��>����
�%?\�^?���w��� N>Ҿ�M}�-�`=#�="X5������<a>R��ͭ�;c˽Y!��滯W?nΌ>I�)�����a��^� ���;=�x??���>;\k?��B?*��<�>���AS�]�
�#�s=�!W?��h?��>b����Ͼ�����5?�pe?7�O>�e�(+��\.�oI���?�)n?�d?ῒ�T�}�t�����6?��v?�p^�rs��5��d�V��;�>�_�>���>��9�^j�>ߐ>?�#��G�������X4��?~�@C��?��;<�%�I��=w<?�\�>�O�*=ƾ!r��2���C�q=�!�>ފ���bv�}��GV,�8�8?��?���>ʒ�����2��=J�W�?h�?軪���c<���,l�UD��k
�<�9�=���W*!�\�� �7���ƾH�
����������><Q@-��9�>m8��4�cAϿ����_оd�p�:�?Ջ�>ϡȽ�����j��,u�;�G�)�H�����1w�>S���{���|��������O�
w�6�>��2���>P=���DK��^U��ۋ>z�?є>B��l�D����?wd�s�˿�"��W�n��22?�:�?X��?1L�>`A�>Ml�<ƒ�kJ)���?�t|?bF?����=ȾV7B>٠j?����2`�"�4���D�\�T>�c3?ԅ�>�a-��{=#�>��>eS> /�]�Ŀ[ȶ�O��c�?vc�?'꾦��>d��?��+?�o�m��骾��*�Sws��A?`�1>|v���s!�v�<�q.��4
?6�/?��p,�]�_?,�a�M�p���-���ƽ�ۡ>	�0�f\�jN������Xe�
���@y����?M^�?i�?��� #�k6%?�>_����8Ǿ��<���>�(�>*N>H_���u>����:�i	>���?�~�?Sj?���� ����U>
�}?���>�a�?���=tG�>D��=����G1��D�%>5t�=��C��?S�I?��>]l�=�iE�Y�0�:dE�A�P�ȑ��C���>	�a?qJN?ݙc>�g��%e�!�;�ԽF�5�(�����E�
�6��S޽O6>\w7>$>D?L�Q�־��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*��ſڔ���lN���3�ӽ|>��>��>�Q𼌳�>�f����n�=�>��==9�>$�>a`>�/<3Eq�K&#��]���#����2��Y��a^�,ao��L���C�܀��,���`v�>U�eE6�߽j�hE�1���A��=h�U?�
R?�p?!� ?��x��>����&=~z#��Ȅ=�1�>�h2?��L?��*?�Г=ҥ����d��_���<����y�>�^I>.z�>�K�>�#�>�3�9��I>~?>w�>� >��'=�ֺ�A=��N>�O�>}��>ni�>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ӧ���h�=Hb.?|>���?пf����2H?&���z)���+���>}�0?�cW?!�>!��w�T�3:>:����j�6`>�+ �l���)��%Q>wl?x�f>�8u>H�3�(b8���P����ɀ|>�26?�㶾�A9��u�ձH��jݾ4M>D��>��F�h�R�������i��|=�z:?�?o5��Lް��u�{L���<R>�&\>�-=�0�=�OM>%:c���ƽ�$H�=�-=�c�=��^>�i?t_d<�}=�A�>�����먾��K>���=B{��}`?
�=?A}�=eoz��&¾$m�:��>��\>܏�Z]�>r+��>3|�>_M>uo+��<h�,��s@�/�^>�"J�ZB���p��}�&>�v$=��=u�<H=�d۽�ý�~?���(䈿��e���lD?R+?` �=�F<��"�E ���H��G�?r�@m�?��	�ޢV�@�?�@�?��L��=}�>׫>�ξ�L��?��Ž6Ǣ�ɔ	�3)#�iS�?��?��/�Yʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�}�#=Q��>�8H?�V����O�g>��v
?�?�^�੤���ȿ4|v����>W�?���?g�m��A���@����>;��?�gY?woi>�g۾>`Z����>ѻ@?�R?�>�9���'���?�޶?֯�?kI>3��?��s?�j�>�x��Y/�U3��%����Z=�Z;M_�>0E>t����eF�kؓ�_i��5�j������a>9o$=��>[1�^'��HO�=�݋��M��S�f�a��>�q>��I>RP�>%� ?�]�>X��>j=v���〾�����K?���?.���2n��N�<��=9�^��&?yI4?�j[�z�Ͼ�ը>�\?k?�[?d�>/��D>��<迿)~��\��<i�K>4�>�H�>�$���FK>��Ծ�4D�Np�>�ϗ>4����?ھ�,��*W��;B�>�e!?���>Ү=י ?֚#?�j>�*�>�aE��9����E���>���>�I?��~?|�?8ӹ�L[3�����塿ɒ[�G4N>��x?$V?�ɕ>Y���7����E�FI���h��?lrg?�D彍?�1�?�??E�A?�,f>���Q	ؾ����>f�.?�e���1�f�ľ,ER���S>�>�P�>�����p�>��>������鸂>��z?��3?�TP��h��t�=ņ=�5�<�M=����t}*����=JQ>����儼
a>`����&�i�k~=>�=��>kV>�*�kb����*?r=�1����3��Q\�z&>�Rܭ>���>f����<P?p�@��7u�.ԫ�F������U�?��?e\�?�qr�j�b�� :?ỷ?�b?-��>���s�޾����Hz���f�:$�<�>���>�����8X��b|��~A��'<ͽ��C���!?#�>�k?�?�!>���>��S�F��m��Mf�iPi�i�1���2�]1D���;�����vCE�850���ʾJ�Z� 9�>c��=��>,�?�9>�R>H/�>֭���q>��1>GY>���>i��>��8>-)�=c]����9�&aS?U���mC������'�>?r�X?�9?���#�}�B�&���?y��?"�? V�>E<f�"��g?7J�>��0��Y?dy��6e�H\6>��ľ�<�.> g=�&`>�Mb��\�	f�%��|,?��?<�!��ĸ���3>����i�n=�L�?}�(?�)���Q��o���W��S��i�'#h��a��V�$���p��ꏿ�[���$��0�(��*=�*?��?�����)��A&k��?��hf>I��>�+�>��>DsI>��	���1�w�]�7J'�{����I�><\{?΋�>8�I?|�;?�vP?�cL?���>�U�>t8��f�>Vs�;���>�
�>F�9?��-?40?y?Vr+?�>c>����������ؾy?��?iI?K?X�?ʅ�Beý�#��Zh�ʨy�Qg��p+�=��<s�׽��t�aU=��S>�s?&��q�8�����j>t�6?���>�I�>�ᐾ��~��{�<�i�>~C
?�l�>������q���s�>/т?S~��A=� *>���=�Ƈ�mF���=L	����=��}�P�>��/"<�t�=��=��x�v]88��:O��;2Q�<Kf?$�!?�a>�=>�q\�G�������>��Z>�@>�V
>weܾ��������g�Go>j��?.9�?5X�=���=4�>0�{�c��
��(���s =���>#"?�<L?Ԡ�?�??�q#?c(�=#e%��S���Z��;ۥ�i�?� ,?��>����ʾ$�3�ƞ?-Z?�:a�/���5)�/�¾Hս}�>+[/�*+~�e���D�tz��z��1f����?H��??A���6�4�边���Z��^�C?e�>uS�>O�>�)�K�g�4&�1 ;>lz�>=R?n�>��?�a6?~GN?Vg�x�2�]t����������ڂ>�?*?_
�?Z,�?b�U?���>���>�"/�:D¾EվGv���Y_=Zׅ��ݗ<��>�H�>��>U1�>Nj>|9���p��b�*���3><B�>o;x>�5�=x��>b?Ep����J?y��>
�J�:������]����>���?�P�?*O?F�S��K/���_��Ҿr��>e��?��?��2?����ɠ=�=�ZY�m���*�>؞>b�>�Z=SW=J\3>�;?���>�p��cH���l�����?p�B?$F�=/�Ϳ��v���N�����nq="z����`=^�z.�An|��O���|;�,��rD�����C���׭��Y�kO���#	?Rf=tn�>��w=L�<�_>=�g˽�/+=o!̼i׋��5��FN=��Y���EZ�����c���/�=���=ڟ�>��?A[!?��?�aP?>́>��d>��=Y�?��t�}�>���xV�G.U�𜖾����9��c������eRQ��퟾Ii�=�H#���6=&P>��B>2	=5ǫ>/�=�p�=|�=�S>�2>��=>Sn>�>?�.>�:>�6w?Z�������4Q��Z罅�:?�8�>�z�=��ƾ~@?��>>�2�������b��-?���?�T�?�?�si��d�>@���㎽�q�=�����=2>���=��2���>�J>���K��⁳�{4�?��@��??�ዿɢϿ�a/>628>��>�R�k>1�A�\��	c�d�Z��Z!?�M;�Ú˾���>k��=_�޾�uƾa1=��6>��^=U���	\��C�=��z��H;=�Aj=�ʉ>VCD>�'�=r���:Q�="oH=�o�= �O>�F����5�0,��1=�(�=�c>E�%>���>�?l90?�Kd?�ٹ>�n�CFϾg���!�>C�=1�>XF�=�;C>d��>��7?1�D?��K?K��>�a�=	�>>�>J�,�c�m���V�����<��?ĸ�?�p�>;�I<�_A��v��.>�AYŽJ9?I1?@t?O��>�\��$࿐�%��.����^/8<�;=�p�^sc�k��ou�bI����=l��>.x�>�7�>�v>��;>�J>O�>$�>�[=��y=:Ļ���<7����U�=M?����<˵ܼ����A�@�=�����uT;<�
:��<�U5<�s�=q]�>�>ϥ�>�=H�����B>"0��[�D��=�]��LD��Je��aw��p9��r�m1->{�K>'5�������%?
�v>�9>�Ծ?�;l?�ܮ=G$��׾F���N�e�GPl�7��=��>��*�I�9��^���P��`�D0�>߸�>p�>B�k>�1+���>��<�=�m���4����>���Dk)�-/�
�p��f������~h�=��ʹC?���X5�=�
~?�|J?�|�?���>H&���پ��->������
=�D�eNq�o�����?��%?/N�>A�,4E��H̾_���޷>�@I�2�O���V�0�9��0ͷ�4��>������оk$3��g�������B��Lr�[��>&�O?��?[:b��W��IUO����g(���q?�|g?.�>�J?�@? &��z�r���v�=�n?˳�?R=�?{>�>�=�u��3�>�/	?���?���?xs?'V?�J�>XQ�;l� >�"��k��=&�>g,�=ϙ�=�d?&�
?�
?)y��O�	�&����_3^���<��=�}�>֑�>��r>�<�=c�g=^բ=_\>��>l��>��d>��>�Q�>��˾�!��_/?^W�=��>�2E?��q>*�n=��D��:�ɽplJ��M$��\ѽ#9��*���䭺`7�=�	��^�>�滿�ϟ?�Z>����g?��G���/c>�:>��Խ#C�>77L>�y>��>>Ԩ>�==>�t�>��:>=FӾe~>����d!��,C�_�R���Ѿ�|z>�-&�s���u��-BI��n��g�1j�[.���<=��Խ<H�?������k��)�����N�?�[�>�6?�ڌ�
����>t��>]Ǎ>]J��/���Zȍ�=hᾒ�?*��?�;c>��>F�W?�?�1�<3�vZ�,�u�n(A�'e�Q�`��፿�����
�u��-�_?�x?+yA?�R�<$:z>S��?��%�Vӏ��)�>�/�&';��?<=u+�>&*��<�`���Ӿ~�þ�7��HF>��o?;%�?|Y?STV���n�f'>��:?��1?�Jt?��1?n�;?�m���$?�53>�;?"W?�;5?��.?��
?��1>���=����	'=e4��z�Foѽ�xʽ<�x4=�#|=��Ӹ��<�o=ɋ�<�yټ��;Ha��OB�<�?:= �=�=�=��>�]?�.�>�@�>��7?�(�Q�7��{���
/?r8=o���b��Z����A�A>��j?��?�Z?��d>B�f$B�̃>C��>�[%>4(\>П�>9��ٷE���=��>�>H�=b!R�c��+8
�)���T�<�@>��>��z>�ꍽ�R(>����0{���b>5iS�0��|HR��AG�1�%�t�8��>��K??/d�=&�ˣ���f�K�)?F<?�M?��?z�=.ܾR�9��=J���Ϟ>��<�9���������:��4;ڲv>@5���\���h`>z
�J|ھ��l���H�#L�u#$=3��`_=2.�6f׾��x�&d�=,>!����!������D��K?�Pe=~N����P�t���>7�>K�>�xf���p��@��d���-�=n�>i�>>�ߏ��a���F�w��m>�>RQE?AW_?k�?"��]s�?�B�����mc���ȼG�?lx�>&h?�B>x��=M�������d��G���>���>i��J�G��;���0��M�$���>V9?�>��?\�R?~�
?{�`?�*?GE?%'�>)������ B&?5��?��=��Խ��T�� 9�JF����>z�)?(�B�๗>M�?�?��&?�Q?�?z�>� ��C@�Ô�>yY�>��W��b��D�_>��J?㚳>m=Y?�ԃ?z�=>Z�5��颾C֩��U�=�>��2?�5#?J�?���>d��>]��� �=��>�c?�0�?��o?�y�=��?	E2>���>��=ʗ�>7��>g?hWO?��s?�J?4��>Lэ<�?��9���?s��&P�Vڂ;�VH<J�y=��'t��9����<Ҵ;nK��$9�����D��������;�^�>h�u>����VN->Bƾ�ʇ��%G>��c��5���͌��;�6�=��>8Y?ɘ>L�ΐ=���>O�>�q�5J(?��?��?�_;2.b�e�ݾw&P�� �>]wC?<��=I�l��$��&*u�Urh=�|n?1�^?��]�����8�c?vX?�P����F�Ⱥ�����]���S?��>�|�)��>�#�?6�q?k
?p�F�Կu�+���$�S���*�LR�=>`�>�F�ި^�,�h>��/?�\�>Џn>,�>K��n�u�4��X?ή�?m�?N�?Ҽ>mj��Uݿ�p�*�����[?���>���Ԛ!?�+��1�۾"���������ڷ���o��!?��Jr����(�c���Ὁû=�?8�t?�[r?]�a?������c�\�[�9X~���X�D��>��;U?�|	A���?��1h�}W�����
��i��<�븾m�_�lص?�4?�����>�K����$eþ�]�>���뵇�Dc=G9�<s�=�x�<��_�� 8��JǾ2�,?R��>p�>; -?>i{���X���,�,.�W��[o]=]��>�^�>���>,ͽ+��q5Q�Ѿ��i��)��7v>�xc?]�K?��n?Ip�+1�����U�!���/��c����B>�j>5��>�W����S:&�rY>�K�r�k��w��@�	�U�~=��2?x(�>I��>�O�?�?�{	�sk��lx�5�1�Ǔ�<>1�>� i?&A�> �>н1� ����>��l?Q��>`�>斌�{Z!���{�R�ʽW&�>�߭>��>��o>N�,��#\��j��S����9��u�=5�h?����\�`� �>eR?�]�:��G<�|�>��v��!�����'�t�>f|?
��=e�;>�ž�$�`�{�~7���O)?�K?�蒾W�*��4~>�$"?Ӏ�>#.�>#1�?*�>qþ�D�ͱ?(�^?SBJ?TA?yJ�>9�=� ���>Ƚ�&��,=Ň�>l�Z>. m=��=p���r\�x�/�D='u�=��μP����<]�����J<���<�3>.�ۿ>;H�Ͼ���y��Kh��ʎ�rK���k��F𽔳��B���@AX����V-s�!�^��Ml�HE��L�b����?���?M�x�hb��ᕿ.�~�5m����>���7l�n߷�ksܽ������׾F���- ��7O��i���g�P�'?�����ǿ󰡿�:ܾ,! ?�A ?7�y?��7�"���8�,� >C�<�-����뾭����ο:�����^?���>��/��c��>쥂> �X>�Hq>����螾1�<��?7�-?��>Ԏr�.�ɿ\���ä<���?.�@�A?��(������T=���>�	?�+@>�1��F����Z�>`<�?^��?�MN=d�W���
�le?Nb<��F�é߻���=�^�=˗=k�n�J>���>Mo��7A�^�ܽ��4>�>F"�<��+^�j �<zI]>n�սA���4Մ?"{\��f���/��T��U>��T?+�>?:�=��,?V7H�_}Ͽ �\��*a?�0�?���?#�(?Eۿ��ؚ>��ܾ��M?[D6?���>�d&��t����=�7�l���^���&V�o��=K��>T�>ł,�؋���O��J��	��=���������s���?=�Ÿ=�>���m����=[�<�����Ͼp���Gzn=]y����F>b�e>?�<>}%d>z�c?��}?�y�>^�>"&U�图-|ھka)���W�І ���O�����{ᮾ�վ�����!�l)ž'!=���=�6R�`���2� �Z�b�V�F���.?*w$>F�ʾ��M�s�-<_pʾG���݄�/᥽�-̾�1�"n�q͟?��A?������V�N��HX�����I�W?�P�̻��ꬾ���=����=%�>���=���� 3��~S�!�3?�?��޾`"k��QV>��+�\�V��{-?�U?��=��>_s?�K{��U�1�A>mg>�V�>�f?��->Lؾ����#?/.]?��!�L7��=�)>w��� k���J���=�r�4�ǽ��>z=<���0Ǽ=ޱ��� ���X?���>Ih.�7�>����G=�J�=��z?� �>*�L>��e?b�$?̽=+N־lM=��k�P��=�cF?��y?&�>��������� ����>�pW?�z?�"4���þ��'�=�\2?�h|?MN?��Ǽ�ˊ�ע��?(�2�?�iv?��I�?M���	�,����@�>T~�>i��>�����>�@?H��
������a�0�6Н?���?UU�?�=ܚ����� ?_�?�����5��~�Bˍ��&�=0�>�ϓ�}��f!�^�OI?��l?G�?�����	����=�c��޲�?QƇ?j�e���M��n������.=�"�=��A�!�����>:2�E�˾�h	�*�����+�&��>_@6�!k�>�,b��;濐rͿX����Jþ2�~�Ԙ?�G�>#\ͽi���`k�؂w�J�E�� F�+҂�EN�>��>�������e�{�)q;��*��*�>��&	�>\�S��&�����(�5<h�>֮�>���>�(��潾ř?�c���?οn�����-�X?uh�?�n�?�p?��9<��v�p�{��V��.G?�s?\Z?n|%��?]���7�%�j?�_��xU`��4�pHE��U>�"3?�B�>P�-�=�|=�>���>g>�#/�w�Ŀ�ٶ�>���Y��?��?�o���>p��?ps+?�i�8���[����*�h�+��<A?�2>
���E�!�:0=�IҒ���
?S~0?{�f.�]�_?*�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?M^�?i�?ҵ�� #�h6%?�>e����8Ǿ��<���>�(�>
*N>bH_���u>����:�i	>���?�~�?Pj?���� ����U>
�}?�>\&�?��=$M�>�Y�=/���Է'�̈́#>&��=��B�qy?,>M?���>l��=|E7��.��1F��yR��e�(D��6�>�b?EiL?zb>�B���v0�Q!��.ͽ3d3�H��F�?�}�*���߽C�3>m
=>�4>a�C�Ҿ��"?A��ӿ���Ö�|?h�W>�?\
��n����=r?tfN>��%���rw��M�8��?@N�?. ?��ݾL�ٽdq>\��>Kĭ>P��6���F��|>��-?/��>����bp����>C?�?x�@q�?�dZ�I0?
�羅����������-TX��p�=��/?Q}��]sk>h*�>K->F#t� �����x�jL�>��?��?��?�Y?Mt�y4=�M�>h��>0 h?�< ?J ��ڟԾ���>�?��%��܇�/�뾸�w? @d�@IOr?����hֿ����^N��O�����=���=Ն2>	�ٽ-_�=��7=��8�?=�����=t�>��d>"q><(O>a;>��)>���Q�!�r��\���S�C�������Z�C��Xv�Xz��3�������?���3ýy���Q�2&�)?`����=�Jx?lD9?��W?��>�6=lz>i�þ��e�xϾD�<}�X>R2G?w e?��9?n23>�"��%9p��v|�k�R|j���>29>$��>���>�n�>l��._>\<�Un>�r>�
�=��һ�$�
4V>1J�>�I�>��>�C<>��>Fϴ��1��k�h��
w�p̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��u�T�4:>9����j�5`>�+ �~l���)��%Q>wl?\g>��v>bk3��8�1�P�X$����|>�6?�Է���9�ju���H��xܾ9�N>�u�>�1�7>�>
��?�r�k��~=ƛ:?��?�������� cu�h�����Q>�Z>v[=K��=�:M>��d�1ɽ�cH��<+=��=͞_>��?��->���<��>�L��dh�Z��>�_>��]>��5?�!?�.��_V�tӀ��M'�g��>�i?���>}/>=���ı�=��>_b~>��ͼ�� ���,�a�+�(#>6�｀�i�D�����<V�D�W��=T��=ž����9�Q;=�~?���'䈿��e���lD?[+?� �=�F<��"�? ���H��D�?q�@m�?��	��V�>�?�@�?'��(��=}�>�֫>�ξ	�L��?��Ž-Ǣ�Δ	�<)#�hS�?��?��/�Rʋ�<l�e6>�^%?�Ӿ��>=~��ۗ�|J��X}l��Uż-�>�)G?L)־�畽��(c?��>0������,�ǿU�|�r�>-��?I��?��e�:\���C���
?�5�?��S?��?>�����J��Y>�@?�P?H"�>H�%����?��?j��?bI>���?�s?�k�>�0x��Z/��6������'p=��[;�d�>�W>f���xgF��ד��h��u�j������a>��$=,�>UE�\4���9�=��
I����f�<��>�,q>�I>W�>v� ?�a�>}��>�x=�n��Iှ����a~M?�.�?*"�|i�s�O�5;�=�����Y?��$?�o��cϾ�Yd>�Il?Wf�?��l?�w�>j���*����V��ĝ׾|K�=�O">�O�>=�>����N[A=����a��ӭ�>��>�[`����E����꫼>�#?^=�>�!u�'�?�?#��=��a>A�[�p���V�A�`��>���>2�>F��?-�+?*a��{3�Nw��Jƴ�[dt�;e->sv?��!?�F�>B��ծ���u>���=����? Re?ۼ��j�>p�I?aV?ծ?�B� Z�P�޾7F>�O�>��!?����A�PN&��	��~?ER?���>�5��#�ս�Kּf��P|��� ?_)\?�@&?���+a���¾&�<��"���U�?�;ΧD���>�>�������=>�Ӱ=�Rm� D6��g<r�=���>=�=u37������<,?UR�!��n
�=��h��vC�! U>��\>-{����U?8�4�,|�,���V����P���?��?g�?�/��!�k���<?��?��?�]�>��F'��ھ�戾���@��1� >�ȳ>�o��l߾E�����5��L������)0�>��>_?}� ?F�P>C^�>_���P6'�|���2�,^�vy�K�8��m.�W%�����Q�#�˗�����}��>2����q�>|�
?�h>��{>%�>T`x�`C�>�:Q>��|>�ا>=�W>�g4>9>�;<~�ͽ1OW?oY��qo!�[����Ҿ��E?�!�?�V?[�̼_��A ?��?�?���>g`�ȼ)���>=�>���qA�>��C=�0=�������]���06�}6N=^��>��<�*W����ӟн��1?�62?2ٗ=����xʾe���9��'�?CC?��Z�N%q���l��\���>��=�=��+��JI��8���e���|�b���Mv��0#�ˉ����E?�E�?!�4��&����:��Be7��O�>g;?�+5>2�&?��g>��$�R�.�Bp�[J7��՗����>��?˅�>��I?�;?�tP?sdL?v��>Hf�>�+��U�>K��;���>� �>!�9?2�-?s:0?%}?�p+?�c>N������ؾ.?��?�H?2?:�?�݅��\ýᘼ,�f�J�y��p���=z�<>�׽�1u���T=�T>$?�P��8�� ���j>�:8?��>�L�>���|���=��>�`?u�>����\�s�`����>܂?���/�<DC,>^-�=�lܼ���:���=���v^�=��ۼ��R�Ln�<���= ��=M�<1��3����:��P<�?Ư ?�G>���>t��&"ؾ����>;:>��>�8?>��d�����^aR�-y�>��?.v�?�7>��>,D�=����Z߾w��oX���>_� ?�Y?��K?�%�?�5?�q@?�W>����k���Ƌ��NѾ�??<!,?팑>N����ʾ~��3���?=[?K=a�b��;)�2�¾{�Խµ>�Y/��-~�-���D��������E{�����?���?aA���6�?x�Ϳ���[����C?)!�>�X�>��>�)���g�Y%�/;>��>}R?�#�>��O?�<{?̦[?�gT>q�8�|1���ә��E3���!>?@?��?�?y?�t�>��>�)��ྕT�����?�>ႾGW=&	Z>e��>�(�>I�>��=�Ƚ�Z����>��`�=�b>U��>���>��>/�w>�L�<I�G?���>Z:��K
������*���iS��zu?Db�?�>*?�J=v���F�ͅ���b�>�&�?���?O+?�Q�a�=i����.���5o� Ƹ>kD�>�|�>�n�=�5/=��>���>v��>f���-�7�HK�E�?�E?�s�=#�¿��r�c����ua�u�d=sd��S��G!��vZ�b�>a�¾�1��ş�&�W�>���4p������Wܟ��S��<�?���;�">���=N��<$N�-��<��o=�>�;֟�=��]��ˁ=
�����09X[��l�<x�=��D�˾��}?�;I?֕+?��C?��y>s;>�3�
��>Ѕ���@?LV>��P�͈���;������ ��N�ؾ2x׾��c�Hʟ��H>y`I��>�83>LG�=KK�<B�=s="Î=j�Q��=�$�=�O�==g�=K��=q�>�U>�6w?S�������4Q�@Z罝�:?�8�>�{�=u�ƾl@?��>>�2������zb��-?���?�T�?I�?ti��d�>L��Y㎽�q�=z����=2>;��=`�2�N��>��J>���K��8����4�?��@��??�ዿˢϿ-a/>��7>'->�R�/�1���\���b�w�Z�f�!?kD;�gM̾i7�>~�=e7߾�ƾ�.=��6>sc=6E��O\����=.�z���;=l=v܉>>D>�i�=�4��M��=JI=t��=�O>�2��S�7�'%,�G�3=J��=��b>8&>���>w�?�a0?�Xd?�6�>�n�OϾ?��^I�>��=*F�>�߅=�qB>ԏ�>M�7?��D?��K?u��>O��=9	�>��>5�,��m�Sm�Ģ����<���?�Ά?Ҹ>]�Q<͏A�����g>��/Ž�v?S1?�k?��>2��N�߿��!���6��a����+=��=5.����<�7N��������Y0>}1�>��>7�>��p>�A>��O>�:�>��>��A=H��=�=[�=�����V<��-���8=%J�P�l�ȧ���.����끋����:������;xi�=���>��>��>{�=�.����,>�䕾�/L�nֽ=|����DB�5vd�x�}���.�C�4�SF>�aZ>���h>�� �?bRZ>��?>!Y�?�>u?��>)�_r־~I��OUe���R�`ж=)4>��<��0;��_�"�M��Ҿ���>�ߎ>��>��l>u,��#?���w=��wa5�k�>�{��W���)��9q�c@�������i�:�ѺS�D?LF����=N!~?%�I?��?���>���H�ؾx<0>UH���=���(q��m����?�'?���>.��D��̾�����>�J�j�O�Vƕ��0�l��\~���Z�>_����tо�3��g��X�� �B�$�r�3��>M�O?�߮?�8b��Z���WO�؋��愽,l?�Kg?�6�>	C??al��C>�����Œ�=��n?^��?f7�?�&>O��=�Կ�y2�>�?	?���?��?s?�RA�U��>E�&<	l>�虽B�=At
>F#�=SG�=��?Q.
?7�	?�p���%
� 8�z��^��-=1P�=>��>#��>Q�t>���=(Eo=��=��^>�Ԟ>U֎>��d>B�>'k�>1�
��p4���`?ŋ>�}�>$?/?�Dp>���s����>J4߾=|�<3���j�t�����=�����Ľ~���ԟ�>��ſ���?Ȁ�=A����	?�C��V�=��o>��>�_�a��>ZK��:l�==-�>�M�>J�G>��>��">
6Ӿ�z>���&S!��8C��R���Ѿ8jz>����H�%�E������IoI��v���j�?j�e-���6=��`�<GH�?�=���k���)�&���B�?lU�>�+6?﵌�U���>���>ơ�>�C��0���ō��o�]�?Z��?�=c>��>-�W?��?��1�$3��vZ�֬u�`&A��e��`�x፿o���Z�
�����_?�x?dzA?hc�<�1z>��?s�%�{я��*�>�/��&;��=<='�>�+��e�`�A�Ӿ�þ^8��GF>m�o?�$�?�X?RV�no�*&>9�:?ڜ1?>Mt?o2?܂;?���$?�k4>?a?�5?��.?_�
?q2>'��=]>��ۨ&=ܥ�������ѽ�ʽ�+����3=�Cz=��Ϲ6�<�=�f�<}��tWּc
1;"����9�<):=<5�=X�=��>�yV?ѝ>�7�>��L?�Uҽ�=R�F:�qe?c�a��%1�>���l�ﾁ��q��= �i?��?�ot?oƒ>r����d�
>=�L>?�d>W�>iʝ>�[��"ڎ�mLp=�;3>~��=?_>7��NO����(4Ⱦ	!Ľ3r�>�F�>�w�>E��(�=��ľ��"��>���{p�pDe���#��4.�*�7�?��l?b*/?���=2�'�侾�.��$�!?qOC?�SD? 	Z?�<=�B�Y`]��-P���*�6E�>�a=�b����}����%�=χ���f>:�N�^�shS>���OѾ�Xi�XwG���C��<���B��<����ž5x����=$s>�¾��#�����A����J?n:p=�Ӓ���M�����C�>	��>��>������5�x�B�����E�=��>%�G>q����t�>rD�B��>�>�QE?�V_?�j�?�#���s���B�����wd��Xȼ��?xw�>wh?� B>���=l���S���d��G���>W��>y����G�E;���.���$�ꈊ>�8?�>��?��R?��
?F�`?5*?�D?�&�>#�������:&?��?<��=o�Խ��T���8��F�P��>)d)?�C�i��>�z?��?F'?��Q?��?��>�� ��;@�Iu�>qJ�>l�W��W���O`>�J?4��>�1Y?A˃?U=>�5�ߢ�q��p��=�>D�2?�+#? �?ָ>�|�>�j��2�=��>�a?5�?��o?���=�K?�B3>?>�>�#�=���>�>}�?��O?ks?�SJ?���>x�<�������!�u��_Z��j;4�H< Rg=�8򼁌l�A�
��B�<�`];�ü4p���㼏^A�k眼���;���>��t>���L+>*�ľH����F>afj�����닾�$<���=;x�>?�?�>�$�|A�=I_�>uA�>���@�(?�3?wo?VS\:�b�F�ݾM��\�>�dC?��=uhl��!����t��}k=�Eo?�=_?�,Z�I���4�c?sO[?)��I?��@���7[��Hݾ�MQ?Z~?�T��D�>Y�{?�s?= ?�a���r����<�_�zbZ����=��>�����b�K��>V�4?&o�>Wh>�l�=��ܾ�w�]/����
?��?�$�?�[�??�,>+�r�J��U�ڑ��B�Q?��>J���V� ?ӭ���������奾�-㾝���]'���l�,�*"��o.���=1�?��t?[y?�d?�z��Yf�Nl`���v�~,a������w�u@;���7���<� �h�����8��$����l�<�X��rd�,	�?�??*t��K<?����Q�@������>"����o�=g61�<���R�>c��үV���ى�b�+?��>�r�>�`?K�s��f�
�𾵕=�i4T�>+�>�_>L�>MR(��fk��5�V(���x�'T6>v7v>:yc?�K?*�n?q�x*1�]�����!�9�/��d����B>�i>���>�W�՛��9&��X>���r�<��ew���	�ˢ~=�2?)�>r��>�O�?�?J{	�fl���lx�ԇ1����<�/�> i?%A�>��>� нZ� ����>��l?���>��>󖌾qZ!���{�ƧʽC&�>�>��>��o>:�,��#\��j��S����9��u�=*�h?���W�`�S�>�R?B�:��G<�|�>ݨv��!������'�<�>a|?���=f�;>&�ž�$���{��7����?��?$����d'���h>B�?��>0�>��?��>4i��5�Ҽ�T?�IX?I�E?]&E?���> ke=�g���Խ�M!�v+=x>��W>}�q=��=�G�߿C�C��aw�=�>�=�j@���ٽd��<G�;�n_<�eZ<oS6>�/ۿ%�L�?}߾(l����9��.�������C��r�P�64��L{���v����b�s��`���}��բ�\�|�R8�?�6�?�HH���H�����避'���>d|����k��I¾�ս��w�ߟӾps��,$"��RS�@c��f�W�'?�����ǿ�����:ܾ4! ?�A ?6�y?��5�"���8�� >KE�<1-����뾰����ο*�����^?���>��j/��[��>ǥ�>�X>
Iq>����螾)0�<��??�-?#��>F�r�&�ɿj���P��<���?*�@:�A?D�(����EsU=���>W�	?y�?>�11��L�
��lW�>#9�?:��?XdM=��W�\�
�mqe?�(<��F�V
޻w�=?�=%=3���J>�]�>o�_\A��{ܽ<�4>wӅ>#y"�|�U^���<)l]>��ս]Y��2Մ?�z\�gf�g�/��T��T>��T?^+�>8�=��,?7H�^}Ͽ�\�$+a?�0�?¦�?��(?�ۿ��ך>�ܾĊM?RD6?z��>�d&���t���=6Gἦ�����㾄&V����=���>��>~�,����ՆO��B�����=m~��Ŀ��5�k}��^����==�ͼ��nY�;�I�͇��I��������=��=�=>��L>V̅=jk5>2m\?z�s?/N�>�%�>]���������'W	=��ܾ��[�q#������������ ��$�U�%��.��Sܾ2!=���=�6R�J����� ���b���F�0�.?�u$>4�ʾ*�M��.<~pʾ���e��z好	/̾:�1�!n�*͟?�A?H�����V�����f������W?�]�$��מּ(��=�����==$�>Ί�=d�� 3�Z~S�Q0?	<?�z���s��L*>@}���=��+?�u?d<�[�>��$?�P,��!�#�Z>>�4>d�>�d�>��	>����ؽ4D?��T?���w؛��я>������y� ^=��>��5�.��[>���<�w��M�]������g�<91o?�_#>l�?�H2��#�=��	;-��=�t?�m>?>�H?Y��>�F>YW��a�,c
����\�d?��?#e>>�髽��#����?�G?��8?���%��1�����3?�=�?Z�I?�����ߕ� �7,�K�&?�t~?�G�M7��0���=@��;�>>?���$�>2]O?;��qZ��[����JH���?��@��?���=;���"*>R�?��9?�.��K�R���l�V��=<��>�H~��z��ھ��t;�i?k9P?Q?��Խ̬� ��=a���N^�?r�?b�����i<���l�qa��ꍡ<�ʫ=����q"�Y��,�7���ƾ�
�<�������s��>gX@�J��"�>o8��7�fLϿ0
���Dо�>q���?!��>ˀȽ
�����j�-Ru�ʵG�x�H������W�>
�>=Ӕ�Y�����{��w;������>O��t�>k�S�b������Bu3<mʒ>-��>��>�஽�ӽ��?�e��#@ο����z����X?�d�?�j�?�b?H^7<�w��{�����G?�{s?�Z?�Q%��I]�}�7�Ik?E��Q`�}5�c�C�٬V>�4?�m�>/�.�b�m=��>�	�>B�>�.��FĿ\z��t\ ����?���?������>kC�?��*?���h���[v���0)�~��>P??Z�.>���� ���9��<��T�?��.?��
�Hl�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�#N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>iH_���u>����:�
i	>���?�~�?Qj?���� ����U>
�}?���>�u�?5�=e��>\��=�@���8�~�">���=�,�`�?L?���>��=��2��-��0E���R�<��9D�-�>��a?y�K?�`a>����5k;�`"�	н��;�9r���68�V��~;ֽ�f1>us<>��>wL?�U�ξum!?�����׿�}���`
���'?�5w>j?�����q�Q>���`?s�j>�9��f���H���;�q��?�o�?�E?��۾����>�W�>���>':���M��U����5>l<?p�*Ȋ�o�l�}A�>p�?G2@p�?T�f��?vD�7������\���,�Ǿ�d=�;?�ؾ�g^>B�>��Z>݁��r9���ϕ�;�>���?���?rb?��U?��j���F��_��"N�>��b?���>�5}�>����>��>���艿fK��^V?@ K@�V?�h����ӿ���S9ھ�Ͼ���<(�>�*>�y��v¡>�l4;�抽�,>�A>@f�>)��>C��>4i>>���<h�>���H)�+������pg��YϾJ��g��� ¾���n���C���߾��)��៽�v�:�8����?�D���>��}?�T1?��P?ᣃ>P�U:�#>S�Ѿ�3�nH���L ��9'>m�U?�B|?��2?�S>�+w��X���j��̾}V;���>*6>��>U��>	�>%k`�E�>��F�t��=��#>t�>�ڒ�:*Y�|�u>�ϋ>{n?��?�C<>��>Aϴ��1��f�h��
w��̽2�?����T�J��1���9�������i�=Kb.?�{>���?пd����2H?���u)�Ĺ+���>j�0?�cW?�>���T�8:>T����j�@`>�+ �l���)�h%Q>Ul?j}>���>�2���6�X}P��J��m�>+�8?�Ӽ�2p#�iSp�&�P�+�ʾ�w>��>�cݻ�2��闿d���]�|�=��=��7?Z�?�	ȽԿ���������B>�Y>D=�7>f�A>�2}�����u&�V�y=a}�=.N>���>�Iw>�=H=>��>�>���������>���=��>��C?�:?��H��iٽ ߆������>(� ?�͊>� ><�q��=��>��>���LH<��|�'k��a�>BƩ��V��R�~�\�=�h���=QA=23�F_�=�
=�~?���(䈿��e���lD?S+?` �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��L��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿđ�>�_�������FEu�8S=��>VH?G��Q�C��
9���
?��?T`��&��n�ȿ��u�8x�>[��?}��?��m�z�����@����>�?��X?��g>��ݾ�X_�K5�>�r@?��P?�г>F��q5"��-?�?P-�?\I>���?�s?�k�>�0x��Z/��6������Gp=��[;�d�>�W>d���vgF��ד��h��r�j������a>��$=+�>KE�Y4���9�=��
I���f�=��>�,q>�I>W�>u� ?�a�>|��>�x=�n��Iှ����!R?s��?$'�)Sb�qZ�/��<t��GH?��?	�C=��¾D�=�g_?�Q�?Һa?Qߏ>�a �����V����Ѿd >NlZ>�-?[�>���-#�5�FvY�k��>X{�>�+>�fϾԃ�ʩ<���>[�#?*��>�00=&?ޚ?�U�>9��>j�}��/����.�D�>��?�D?2��?$?f{���O.��q��^��< W�<�>�ր?_�2?Xt>7u���՛�]�>	��O��<�"�?e2;?13�V��>yl?�M�>��?޷A��OY=��������>J�!?�O���A�[&��(�!P?�|?���>������ֽF׼}&�"����/?d#\?�"&?����-a�	þ��<P��ؽZ���<��F��>g�>k���޴=|$>zd�=�Um���6��dd<ߍ�=?�>��=��7�Mꐽ
u,?�I��0���Ȟ=��q�ևD�6{><�N>J���35^?|�8��r{����g��V@U�5͍?c��?��?����Rh��=?�ˇ?\�?�B�>�b��Km߾��-�v���y��9�� >)k�> �e��[�-��kR������=oƽ������>�i�>�t?a[ ?��S>�]�>%��1'������,�]����|6��-�������ɗ#�2/�J¾r�~�>�����گ>��
?��g>+�z>��>i�;�`�>F�N>��y>j�>�YQ></2>�� >��;��۽XEg?7M���� �xC)��ء���*?���?}�&?Ja���GL���p>Y�?�G�?�7�>aˍ�YLQ����>���>�Z�OX?w��=�1�=��.۾��P�������=�C�>�{;��w���7��a�=�3?� F?�b>7A�������6�F<7&�?��-?��T��H0���j���T��+��2�=���D#W�֊��m�^�~�������x��c����=�4??璌?����#ྏ�޾0񏿤� ��?�>+�?�>��?Vw�>��ݫ���i���-�_+���?xo�?N�P>\�f?0�?��??�r>? �>�[�>�ۙ�[�|>uoM�I��=�I�>��F?�.?��%?�b.?ю?;*?>�=(��^��o��B?j+?�?� ?�?$ q��=�A>�"��2ni��pV��/���Z�T����x�<��!>�)?����9��(�Vq>}07?�;�>>7�>5���	����$=��>��?A>�>^��mw�8e�=��>���?e����<�a0>���=��ۼ�>ʸ��=�R�!��=$���T�t�<���=�:�=�Z�<钜�`�R�s���o@<��?�E?:�L>��>ե5�r ����"�N:	>�^Q>t�H> N.>#�[ދ��6��H�]�a�>ᛒ?�?D#�=��>9��=�#�����H��v�����=;��>�e?�kF?�s�?��#?�\9?�j�=����g�����!��˂%? $,?ޕ�>n��6�ʾ�憎و3�z�?o_?-<a�t���6)�ӥ¾�Խ)�>vL/��$~����D�ʚ��������c��?$��?XA���6����h����]����C?�!�>�x�>��>ѿ)�s�g�N��<;>/��>�R?@�>�&P?�{?�o[?�mS>�T8�5��⬙���D�7 >E�??���??�?8[y?���>%>�t)����>��a!����т�%�U=O0[>��>;�>�֩>j��=��˽՚��H�>�炦=�^a>�_�>�ӥ>x��>�x>"��<_.H?�~�>5p���q	��"���0��/���Pu?5�?�)?�5=G��K�G�q]�����>���?j�?M�-?��M��M�=�^�i3���t�^��>�ļ>2��>�'�=G�A=c�>o;�>>)�>)�۲�ď6�j3@��?#=D?�g�=�R���|����=E���!@>,꣼�Bž�)h��Ӿ5⽠�&��L[>��Z���aʽ[�þVz���q�f��>��Ž�>L�=3�>v�,>Y
Ƚ���>�����!>�!k�U������z�:�i
>Bd<N��<��m>�f��*ʾ�|?�b>?��&?�76?�*Z> \J>B6����>:����	?qi>��ۼ���:/�������v��Cľ]�˾GP^��h��K&�=n��s�>L)�=��=M��d%>*\]=���=Ӡ2�'��<�y�=��=]��=�F�=Y�&>l�>�6w?0��������3Q�EW�Y�:?I7�>�}�=<�ƾ3@?�>>�2�������b��-?W��?�T�?��?$si��d�>W��j䎽�m�=����>2>��=	�2���>L�J>Ӄ� K���{��24�?o�@j�??�ዿ��Ͽ�b/>�6>��>fhR��V1��Q\���c�k�X�+ !?K{:���˾N�> ��=7�޾��ž��1=��8>6<i=����[�s��=�]z�Y�:=ݧk=2��>��C>eѹ=�7���z�=�oK=!W�=�3P>]��T�;��)�'F7=t��=�oa>��%>���>�?X0?�Od?w-�>��m��Ͼ�4��1�>ғ�=�-�>ժ�=��B><��>H�7?�D?��K?#}�>oǉ=��>���>q�,�q�m��P�߻���3�<���?*ˆ?}θ>DQ<z�A�[���m>�HMŽ�s?>I1?�h?:�>��1���4���:�\u���sv=/�p=�p����	='�����y9���=}��>���>\�>s�p>CR�=-F>�Է>h>��<�ٿ=4�<k(=�v�F�=ʘ����-�����+���������/�`�N�,�[nM����=���>�:>���>���=��z@/>з����L����=7F��C,B��4d�pI~�
/��T6��B>>X>�|��4����?m�Y>�m?>R��?^Au?T�>�!�2�վ�Q���Ee��XS��˸=͵>��<�cz;��Z`���M��{Ҿ��>�ގ>��>K�l>S,��#?���w=R��a5��>�{��^���)��9q�\@������Fi���Ѻ1�D?GF�����=[!~?�I?z�?���>6��u�ؾ�70>�I����=�+q��j����?/'?��>��l�D��z˾RA����>}�I��P��ҕ���0��������	ֱ>���T�ϾA=3�\l�������B�sr��'�>�O?oخ?=+b�xx���kO��-�R��j7?�ng?WA�>{�?N�?!ܠ�Ǩ��뀾�&�=y�n?]��?��?�_>�{�=�j�����>HT	?�Z�?���?`Os?2�>�ų�>�X;\�>r/�����= �>헛=k9�=�
?Y�	?Id
?�s����	�3��$��K�_�g =�آ=_ё>&�>��w>���=c=��=�Y>,Ӝ>7�>�d>���>�0�>�������/*?�	>Z��>��3?�f>#=��ݽy��<�˷��T!���fL����r�;A�}��<`I����>��Ŀ;ޔ?<L>���w?���0��;V>�IW>7���O�>�;>��t>���>#�>RY>먖>��>�6Ӿ�^>����M!��DC�~pR��Ѿ=Cz>�~��Ժ%�ڍ�����OI�||���]��j�*��i0=�fW�<�J�?B
��.�k��)�`T���^?�]�>�26?���L���J>;��>$��>�+������`ƍ�[|�x�?$��?8?c>��>�W?�?w�1�x3��wZ�¬u�~'A�e���`�|፿y�����
� 	����_?P�x?{A?�Z�<�8z>{��?��%�}ӏ��*�>�/�U&;�(:<=�*�>�)��
�`��Ӿ1�þ�8�VHF>ӕo?�#�?Y?�NV�j*��t�>(R?D?(t?��><�J?�)I�6�3?��>�Q�>$�>��?1�?���>O��>w�k>&C+=�	=�нEe�������0 C�<���gw=ԩ�"�_>¢�=�S>E��;W{��r+���V:=���@A�=?�=�"�=�<�>ȻQ?��>���>��+?�G��;:�����ڒ+?�=o�ɽ��\�ʾ���Ρ�=�h?��?̈g?W�]>܈4��^/��b�=@Q�>�D>��>Z��>�x,����|�=�"˻���<�3�=�I�0�a�@���ٰ�~<Q=�:>�� ?)9�>����7]2>����J���)�`>��!�|�̾�^���;��2���,�x��>��R?��?-��=��������j�a�2?��<?��N?O�j?2��=���eJ�/F�V&�+��>_�>����sj��� ����,����;��>V2w������L>:���M�þ�q��H�#;��TI��H�M=�
�{+Ͼ��u�:һ=,�>�bþV�#�R���۫�ILL?�F=�5��Z/����@�.>�̏>`â>�P���/x�,�>��S��u��=#:�>|uC>����4��-*F�f��n>�>_QE?4W_?k�?"��Hs�9�B�u���yc��.ȼ9�?`x�>-h?B>���==�������d��G���>���>X��A�G��;���0��F�$�ꊊ>E9?n�>k�?d�R?��
?{�`?�*?CE?#'�>�������@&?ԉ�?��=�Խ��T���8�(F����>�)?1�B����>�?6�?Q�&?5�Q?��?�>� ��A@�m��>�V�>\�W��a����_>�J?��>�<Y?�Ӄ?��=>�5�_颾[۩��H�=�>��2?06#?�?���>� �>����=l�>��b?}�?��o?/��=�? 1>�
�>T��=?̟>:��>!�?�/O?��s?H�J?S��>�g�<<��������r�91F��^q;��F<��z=D: �8�p����7��<�w�;���׈������F��铼r�;.��>���>�ܙ�T>���������Y>�	�����򇋾*�;�b�=��>�$?ȣ�>ӹ����=�m�>
ݾ>���yG)?�� ?�_?˴Q���^�z+�^�L���>1E?���=q<l�����u��j�=6+p?
�^?�b����.�b?>�]?�r�==���þ�/b����/�O?}�
?�#H�h�>j�~?r?I#�>c3e�MRn���(*b��'j�Jx�=�Ӝ>WD��d���>�f7?���>E�b>O��=�ھ�w�鶠���?��?[�?��?�**>��n�p?�
7 �g���]?���>�ݩ���?�<��վB���U�����?ժ�⇪�����^���b%����\�c�=?��s?ss?��a?�S���`��]�O:���W�@?�(���KB��IC��qA���j���xv��4��;V=�"ھH�^��`�?�CH?wԶ��8�>�Ӿ	�*�@���:η>����8z���%�=����V4>E^���^A��%Q��2?���>��>ڌ6?�[��}%��Z%�$.�խԾ��j>��M>+��>[,�>~�M��� ��a̾N=��^,��]6v>cyc?J�K?¸n?p��)1������!�f�/��e��
�B>�h>½�>*�W���t9&��X>�(�r����=x����	�Y�~=e�2?�(�>���>sO�?�?�{	��l��Xnx�>�1����<=1�>�i?�?�>z�>5н� ����>��l?̨�>f�>,����Y!��{���ʽ�%�>�ޭ>u��>�o>ߪ,�#\��j�����-9��r�=̩h?G�����`�#�>R?wo�:��G<2|�>ץv�s�!�3����'��>v{?&��=�;>��ž4%�~�{�8����&?#:?DQ��+�(���w>)�"?9I�>Ub�>m�~?��>v�Ⱦ�8:J�?K�`?��J?��B? ��>�==������׽I40���'=W_�>��V>�	`=!�=���R���Pki=��=NP��!�2��:���>�<�%$=�
@>�/߿|Q��ꮾ���f���{{��+����O�d��H���6Ѿ;�����f���>�M�'�cfL���e��D��D#����?V��?-}ѽ(�ӽMc��fc�u���wp>�`����ս��¾�Ρ�M�����ξ�2���%�b+Z��4l���k�Q�'?�����ǿ򰡿�:ܾ6! ?�A ?8�y?��7�"���8�� >�C�<�,����뾮����ο@�����^?���>��/��p��>ܥ�>�X>�Hq>����螾U1�<��?7�-?��>��r�0�ɿc���$¤<���?0�@��A?��(����;T=E��>��	?�R@>��0�Y]����g�>�.�?U��?|N=��W�M��~pe?�m<4�F���߻�P�=��=A�= ��xJ>���>[S��CA��ܽ�4>��>�c ����^��u�<^�\>��ս��Մ?"t\�f���/��S���X>��T?H.�>�.�=>�,?�4H��|Ͽ=�\��,a?�0�?��?e�(?�޿��Ϛ>	�ܾ1�M?wD6?���>e&���t��G�=���>V��A�㾓%V���=]��>Qx>��,����O��W�����=|��ǿ����J<	(���yb��s'�۹!��!f�抪���ahн��<�:�=y(Q>��>��C>�R/>}�[?�qu?v!�>��R>���������ɾ�F����]�H����fK������h�-�۾�,�+J�M��f۾!=���=7R�j���B� �i�b�R�F���.?w$>_�ʾ��M�a�-<�pʾb���
܄��ॽ�-̾�1�&"n�l͟?��A?������V�W���W�����Q�W?=P�һ��ꬾ��=|���>�=%�>���=���� 3��~S�U_/?��?�G���"��K*>-���)�=>I+?�L ?Y�<���>��#?�}(��� �Y>��5>��>S��>��>dׯ�X?���?��S?���{���9��>�ռ�*�v���i=_>A�;�J��V>�lP<i���<sl�Z'�����<)	k?�_�=��G�:_I��A����=�->xy?,'b>��E>��]?�>�܄=Nb˾�wW�>!��zm>�\D?Ǥv?>����󁾙�¾��>+�X?H�.?�;5��"�s�(ԾY�C?C��?�X?q�H:�����^��k�^(?�%�?�<��B��K��+�=1�>h�<��?�־�r>=�a?I���%��GP��Vx�f�?6�@�?h�=����B>­�>�s'?#�p�Y繾�I�4֩��N�^�>�~�`8��\��D�="X?%B?��?�椾�澫��=敾�[�?N�?�����g<t��al�p��w��<��=���"K"�g���7���ƾ޽
�尜�*}��&��>�X@�r轇(�>!m8��8��PϿ����Kо�<q���?>�Ƚ����j�j��Pu���G���H����pl�>�>�_��+���/�{��b;��2���/�>����׈>�mS�]{���Ο�n�1<�>Y��>3�>�L���������?uk��_3ο"���
��ܱX?s�?�d�?�\?r�C<�:w���{��|	�!G?�js?��Y?1�&���]��6���j?0z��8`��5�l�D��GW>64?�f�>�-.�Pfp=r�>��>.b>)�-� Ŀ,]��&��k��?�z�?9��d��>cu�?/v+?�k�*���i7���*��D�:�k@?�r/>���� ��F;�xw��y�
?AA.?�#���\�_?'�a�M�p���-���ƽ�ۡ>�0��e\�EN�����Xe����@y����?M^�?h�?ص�� #�e6%?�>b����8Ǿ��<���>�(�> *N>�H_���u>����:�i	>���?�~�?Oj?���������U>
�}?��>Jև?��=�
�>bs�=:J��$���`#>��=d/�����>mRF?&M�>B�>C���G(�mE�4�T�3����G���>.b?-sG?�_>�f����W��)�M6����z����<}	�B��ɭ�sp>27>��>��B��%��3E-?Qc�^ӿ�Ҟ��7�P!?P[#>�E?sH¾�!?�Q*=~j?$�>:&��A���'��i�+��r�?���?��?�����tY=ap?���>�����F�w��'=�$?�齳5z�݃����> �?��@C��?�dm�4�?������D����� y�#�5��D?񬒾+�N>�R	?��u>�F}�/A���{�~��>��?/�?o!?�R?��a���,�T�=�&�>Lɀ? ��>Ҳ�:�뽾%��=n?4��E%���S?\v@)�@Á?�����ѿhp���ɥ��r��u>�=��=�p!>�&��h)>P�>'��.��w]�=�N�>�~>��>bWW>d��=�>���H�*�EK�����F�\��������I��$�:���	�5䳾�;�ս����g��_8��7�'����:�=R|?�&?RL?w��>�O�=BA>1ھb%5�;�ھ�4���>��L?�5w?��6?u^/>����Ia�aU�9̾�C��H��>qۥ=V]�>Pe�>(��>$����}=ftW=��=*>n.^=p�j;�0��1�>��>��?� ?�C<>��>Fϴ��1��k�h��
w�p̽1�?����S�J��1���9��Ӧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��u�T�4:>9����j�4`>�+ �}l���)��%Q>wl?�bi>/�z>��3�c7��	P��I��u\}>=6?Q��?�6���t��I��pھ��R>���>w�����r���~���n����=[f:?/C?��������&~�#�����N>�ZX>`�=LP�=(L>!�q�_�Ƚr�E�;�+=�m�=�]>�?m�,>!��=���>��`O�2��>&�B>�_+> m??��$?2���U������.�{w>;l�>���>��>��J��ĭ=� �>��a>oy�	Y�����#?���W>iz���^�p�~��_s=�F����=5��=�P�ӧ=�4�!=�~?���(䈿��e���lD?U+?k �=w�F<��"�C ���H��G�?r�@m�?��	�ߢV�@�?�@�?��S��=}�>
׫>�ξ�L��?��Ž3Ǣ�ɔ	�1)#�iS�?��?s�/�Xʋ�<l�q6>�^%?��Ӿx��>t#�ռ��3H���
p�Q���m�>p�P?]������<����=@?R?�>!���﴿�oǿR�|����>���?$��?w:e�	Z��:�H�P}$?6�?��E?�G_>��߾������=/c+?I?/X>�����q�? O�?��w?RI>���?�s?�k�>�0x��Z/��6������p=0�[;�d�>�W>_���sgF��ד��h��o�j������a>u�$=%�>FE�U4���9�=��I���f�:��>�,q>/�I>
W�>n� ?�a�>y��>hx=�n��Tှ������O?�:�?���k�d���y<�;�=?
�[�?L�#?���<��¾�Jf>�Z?HV�?Áj?bn�>���u������J1˾Ш�=�N>W�?a�>��}�w��<���k�8��ٖ>�&>Krȼ��۾����@w�<b�>d�!?J�>(i$��#?��?��k>�W�>�1q�������E���>׃?١D?��?�4@?a���)J$��_��׺���pl��wl>�΃?�w6?���>��������ݝ>�޽���<�*�?,D^?������?��f?�@?2O9?��ܷҽ�b����`=���>B ?�_��E@��%�tF�>	?�?7��>B~�����L�;���~?�c\?$�'?y��Һ_�9����S�<�؎�5�x�f��;��U���>3�>�6w�ٺ=��"> a�=B^o�s�;���x�ǉ�=9�>Ia�=��-�zwk�?|,?3CP�pㄾ��=;�q��)D��T{>��M>X����J]?�,8��5{�vI��+d���AU�e	�?���?̫�?n�����h�j=?X��?��?�`�>Z/���.߾���V�z�O
|�b��e�=���>ҼN��H�8-��<,�����_ƽZI3�Vq?sw�>w�?`�>xOV>p,�>S ��v�7��u����b������%��:,��#�fr����6��<��ľ y����>�Z�wֱ>*A�>��O>߀v>NG�>�F.=mh�>C7�=��*>7��>�$#>\��=�kV=�K_�*t�pd?<���AQ'�E���풾��<?��?�?K��<y�����#T�>zĖ?Ƕ�?�b�>����/:����>�9?�x�c|/?N�=���=(
;���ž��^�����K�*>KH�>[Kh�2o?��3;��6���D?�`G?,ɔ�#���2ؾq`�����5c�?E,D?�f���b���z���Y��8�@��>�yl�"+����ؖh��"q��=��󽃿\y%����v�L?���?�9-��������Қ���~��m�>^�#?�^�>�@;?W&�>�$�qn&���r�;������?6��?�^>�>V?�1?[5?��/?綠>+�>�Q����>�W���1>���>+g<?��.?0k&?�!?��#?�x#>�M������B��p�?M�?N�?.��>�Q�>�?E�%bZ=�߰=	�<�����\�d��������K�i��7g=YR>�V?y��8�^����Li>'�7?`�>��>�������'=®�>�|?�>Ђ�� �u�(��Q�>|
�?�����=�1>E�=�0���л�:�=�ު�q�=�ꑼ�N�a<��=�Ǯ=��5<�  ;$���(�ں6'�<��?��?���=��>���=d�5�(��Q>zW>'�=���>I��[�����m@\�Vh�>�Ś?#R�?���=��&>�6=yמ�!���O�!��xQ>}� ?DT? �j?�{[?)F?�E?��>;��*��*L��!����!?\!,?���>t����ʾR��3�-�?M[?_<a����,;)�)�¾4�Խ�>�Y/�0.~�N��zD��9��}���y��ܛ�?���?/A�q�6��y�����\����C?��>V[�>'�>W�)�1�g��$��/;>���>PR?��>��O?�2{?G�[?�[T>�8�_*���Ι�</6�n�!>�
@?A��?��? y?t}�>0�>V�)� �LH���'��*�pނ���V=VZ>���>
-�>��>��=��ǽ[���>�aF�=nnb>q��>���>�>��w>���<y�G?i�>���!������~���jH��u?�W�?��*?I=����tF�cv����>�\�?��?-�*?yR�h�=�ܼ�����9t�EC�>���>�̙>�1�=��H=>���>���>��,�DK8��:P��R?"+E?�d�=n���������>�:>P�g�]�����Ȝݾ��㾈�C>!���>r��駾����������ݾP��4?G���WL>~7�{�u=n
>��Y�\>h��� >bu	=&�.=� ��=6+Q���<��k=?i>Ok=7zݾ�o??�?�S?��3?�x>M}�>6�S��!�>ǔӽ�&�>FE۽���x���"L��+����{5��ގ��75��m���>б���g>���=؋> ���_>^>�@�=+�=��=��=�u�=���=��=�]:>4<�5w?闁�t���r*Q���۱:?��>���=�}ƾ�@?{�>>�4������ec��#?��?eV�?��?@bi�vc�>���3鎽��=�ќ�=2>O��=8�2��>��J>F���M��[>���/�?9�@ؖ??����1�Ͽ�t/>�r6>��>�KR�B�0�3*[��`���X��T!?�;�#;���>��=��ݾ(2ž5d,=�.7>��g=�x�j9[��'�=������;=x�k=-��>��B>���=�����ٸ=SQ=F��=��J>9��i3B��_2�KT,=�a�=�`>��$>�"�>k?r�/?0�c?���>Dl�kYξ����J��>���=�>��=q�C>�|�>�8?��D?��K??�>4��=O&�>N	�>vO,�wUm�
征���p��<vv�?汆?�_�>'f<��A������>�SxƽJM?UD1?{?m}�>�U����8Y&���.�&�����4��+=�mr��QU�0���Km�8�㽲�=�p�>���>��>8Ty>�9>��N>��>��>�6�<�p�=�ጻ���<� ��}��=h���u�<�vż����yv&�>�+�>����;ۮ�;�]<���;�~�=���>)">���>봖=�볾�d/>�����L��6�=�]���-B�d��,~�
/�fG6�%�B>X>r*���,��_�?t�Y>�g?>�x�?�%u?��>�����վ�<��|e�#�S���=�n>f0=�l�;�RY`�6�M� �Ҿ���>4ߎ>��>��l>�,�`#?���w=2�'b5�p�>�|������)��9q�9@������ii�w9Һ�D?�F�����="~?��I?t�?W��>���Ɔؾ�:0>)I����=Z�J*q�uk����?D'?-��>H쾦�D�|̾PH���ķ>�cI� �O�rɕ��0���_���2��>�Ӫ�͠о(*3�Ge��?��g�B��r����>��O?�?v#b��_���]O��������%e?�{g?��>�.?�9?�ӡ�bs�֣���m�=�n?���?�>�?w>	�=TM��!M�>�Q?�ܕ?�(�?�r?i=��G�>�)ں��>
;��e,�=�>��=Q��=r:?=	?��
?cģ��6
�mﾓ9�-DZ����<on�=��>>ϊ>�<v>�>�=KH=�:�=��S>��>同>yb>���>鞇>�6����v*?P�>+�>,2?
�z>�=��ƽ��<x肽��/��5#��Ƚ^/ս&,�<�ap�Dy$=_:����>�Jƿrە?|&K>��z?��Q���M>)�\>�ͽ�"�>��B>��~>�ެ>3�>b�>�8�>�(>[.Ӿ�E>N���F!��OC���R���ѾkEz>����X%�-������lI�����c�;j��/���/=��'�<�K�?6���B�k��)�4����_?La�>wF6?���W숽|�>���>���>_,��~���CǍ�`i���?���?<c>��>��W?/�?�1�3�%vZ��u�d(A�Qe���`��፿#����
����1�_?D�x?[yA?�S�<�9z>;��?��%��ӏ��)�>�/�';�rA<=�+�>�)����`��ӾM�þ�7��HF>a�o?%�?AY?�SV��j��)��>R?~��>�|�?��>G�N?�ɥ�j�U?��=
;�>�u�>��#?�N?���>���>;�>���__Y��Q��X."���K;��^�D����(:\��_�=��i=�Zw=���=k�Խ �1��]�=�ހ=�>=�"W=��=���>��[?s��>��>G�7?t��[ 9�F���S*?�L�<&�v�P��������𾌹�=��j?�o�?sW[?�Ff>�CE��D���>�2�>V%>��X>�Z�>�޽��;�
�=c�>z��=�֟=�fU�(;��ؗ	�ْ�i�<��>dr�>Ѵ�>Z'�_4>t�������V>�sʽ�ɾȳD��4�S�1��ǽN��>��b?�?>k='\��N
��Br� �"?Y>?��I?-�P?���=<2	��cN���7�⌔� �6> �	>s!ؾ���RO���'�U�o�8�A>�?Y�V��R�T>�� �XȾ1�n���H����[��<���=&2�y޾wi��X�=%�>���������f��!wJ?T�\==���}�]�䷾:">�>,�>��6�.�� 3������=���>�o>>��
�q���E��@�
>�>6QE?HW_?!k�?7"��Ms�Q�B������c���ȼ �?x�>,h?�B>-��=F�������d��G���>���>N��A�G��;��H0��6�$�E��>Q9?�>��?Q�R?u�
?l�`?�*?&E?'�>x�������A&?8��?��={�Խ��T�z 9�BF�y��>q�)?-�B�ٹ�>P�?�?�&?�Q?�?��>� ��C@����>xY�>��W��b��G�_>��J?ؚ�>n=Y?�ԃ?f�=>Z�5�	ꢾ�֩��U�=�>��2? 6#?K�?���>���>'���\�=}��>�	c?M.�?��o?�^�=R�?2>)��>N�=l��>|��>�?�YO?��s?\�J?���>��<�H��[=����s�
�M�_��;��H<i�y=����dt��e�w��<�
�;��������>�
E����(C�;���>�8t>t���%�.>�þ+$����A>͛��p}��*h���3<�ܩ�=6�>I?7M�>~f$����=:��>!�>y��;�(?\�?!�?"�;�b��r۾��J����>L�B?���=�l�n��;Vu�`�p=�[n?��^?-OY�KS����b?��]?.��-=��þ�jb�|��b�O?��
?jI��>�m~?<�q?ڷ�>5�d��Kn��!��r?b��k��Q�=b�>^1�H�d�&�>�A7?���>.Cc>���=Mھ=~w�i����?}�?��?��?_�*>��n��E�r!�쀐��%_?�\�>A�����?n1̼�x���*F�������j��[}��͊��q���7�������P=���>�^?��w?CXp?�R���d�a�r��]���_�����"#�w�2�*�4�NQI�+0V�̑��F뾷���n:��]����V�В�?�eF?r�j��Z�>ɯپ4�3�����>#��i�A�a>Τ�<!�=�7�<�׆��th�����6?���>�4�>{E?��\�[^O�� ^�;�Jɾ-g�>�հ>f�a>X��>���b����S��L��X׾��V��6v>�xc?#�K?v�n?#n��*1�����D�!�5�/��c����B>�j>*��>��W�˜�:&�HY>�-�r�%��=w��Y�	��~=k�2?�(�>��>�O�?�?O{	�'k���kx��1�D��<�0�>h i?�@�>��>�н� ����>��l?���>��>����qZ!���{�ЧʽE&�>�>��>��o>8�,��#\��j��S����9��u�=*�h?���X�`�T�>�R?��:w�G<�|�>ܨv��!������'�@�>b|?���=c�;>&�ž�$���{��7���A)?�]?�ے���*�gS~>
!"?V}�>��>��?	�>LdþJ�.���?��^?�EJ?_WA?�L�>==D����Ƚ��&��~,=�c�>�[>pm=2w�=y��m{\����;�D=z�=߮μiu��Y6<�d��G�H<Ii�<K�3>�kۿ�BK�q�پ���4�b>
���F���i��Ҥ�vo�����Px�Ƈ��&��V�+:c�����{�l����?�:�?	{��"��R��������������>z�q��"�櫾����"�����Z���e!���O�"'i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >uC�<-����뾭����ο@�����^?���>��/��p��>ޥ�>�X>�Hq>����螾^1�<��?7�-?��>r�1�ɿc���o¤<���?0�@��A?&�(��(�c�O=<��>��	?eB>(_1�}�����, �>�I�?0)�?�FK=�W��/e?��<�9F�ɕݻ�4�=��=˟=���r�I>��>�=�/�C�����1>�ڄ>��%�:_�N�^�.�<a�[>Ǉٽ�5��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�󉤻{���&V�}��=[��>c�>,������O��I��U��=W�F�ƿ��$��|��_=j�ܺ�[��7���~�T��#���eo�L��ˍh=���=��Q>�k�>�$W>3Z>gW?^�k?{N�>Ҁ>�7佘��ξ����G�����k���g��g�ZR��߾a�	���������ɾ=��(�=�9R�����"� ���b���F���.?�`$>��ʾ��M�7�*<vʾ�������m���A̾`�1��%n��ǟ?�A?t���V�W�����d¹��W?mQ����xݬ���=tK���=8�>��=ͺ�@&3�v�S�Vy0?@�?��������*>���=��+?�*?|]q<H�>�D%?.�*���>\>��3>M�>�<�>��>MU��k�ٽ�?G�T?�s�藜�Gv�>����pz�`=�>�3��S��\>"ɑ<�ό�OM�_������<�(e?2�>�rH�6Z��3�8S4>R�>�it?��7?��>�%m?�$;?��$>I�"�.4��=��9�C>C�z?��~?�D>��u�\^��9��H�?-XX?[�?���-�b@X�f�"�s�?[��?]T�>�\7>�����Ǧ���3��C8?��{?��I�����K#�V"�WE%>h߶>��$?�{����>�?h?��$����L�ÿ��3����?��@R�?f�=��b�c�f;%�?땿>�u�����w��ݸ�����<Q?�Y.�H
]��q��R4>�\
?djQ?�N?:.���k�gl�=����Ku�?]�?����R�<���]�l�����9�=7��=�&��g$�wz羗6�+pǾ�l�jٟ�3E$�ǌ>��@�R��M��>j2G��㿞Ͽ䅿�ξOf�s�?�j�>�Sٽ)ި�5j�t�t�C�F�]�I�걅�*Q�>��>�Ɣ�������{��w;�.U����>���>��S�b)���F4<WՒ>���>h��>�"��E۽��ę?._��;@οu���7����X?'f�?�n�?!v?�8<��v�c�{�����$G?6�s?( Z?��$�y1]���7���j?����{`�{�4��D��XW>_.4?�V�>z8-�/c=�6>���>7�>��.�`7Ŀ�'�������?���?���"y�>�@�?�+?8���$��4ت�߶*��nŻ�??\M+>	�¾�"�B�;�����c�	?8B/?`
�S�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>W�?�]�=���>Z2�=B��#�Ҽ�->J<�<�-�<�g�>�AP?f��>Kl6>k¾�t���H8��5Q�2��;�F�Fb�>zQk?�X?��4>�*=���6�<(��2��g�k��<B�����l�w����9>��/>�E>=���ϗ��$?� ��Pؿf��Í*��h2?��>di?����s�[���8m^?�*�>��a��V�������<�?$�?&		?A׾͌ݼ�r>Ⱥ�>���>��ս3뜽Om����4>�A?�%�|׊�wRp�}`�>�A�?T�@�֮?�nh�=l?���jn��7u�����>���1�GQ?OP����(>%�?�\>���fͻ�6���8��>c۠?c��?�U?��U?�V��<�S8�<#�?1�?D� ?kc�<D��
]">~��>����./]���`g�?!� @�@�͑?����}�ѿnM��-<���c���P>�_=�Zx>}�^����=k�� ����<��	��=]��>G�q>�т>`A>b>"I*>������$�y��0�k��W�G�!�)u(�a�Ѿ0�|���MO:�._׾jоd]��.7�PF߼�/b�HP!���ͽx�>X-|?6�#?q�s?��>fm�;�&>_E�������Wi=V�?M�+?)�a?3�F?��=7!����Y��]��8վ��5�8 ?˳�>���>}"�>R�>�4
��4>���y̗>,�!>��5=<���1��={o>ǳ�>��>���>L<>ĕ>�δ��1����h�E	w��
̽o �?낝�L�J��1���>��i����s�=�c.?t>^��c>п�����/H?�񔾎'�L�+�A�>`�0?_W?��>����dT��>>>��ϧj�f>� ��il�ω)�(Q>[f?2$�>�Ӊ>��7��Q:�d�>�j&��zۀ>�4?����U,���u�!�H��qھ��i>>�>��N��]!�W����ل���t�g�>5�9?��?����֮���E��H�0>@�>vW�=^��=C�W>D���������g��=&��=�a?>�{?e+>��=�>�I��l�P���>D�D>��->�5@?��%?D��ri�������.��x>q��>$�> ,>jJ���=C9�>�a>�����ܤ�5?��W>�=�M_�(r�/zv=������=�O�=]� �"�<��,&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�/)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�l�>"y��Y�����!�u�i#=��>:H?j?���O�I�=� q
?�?�h����*�ȿ�xv�5��>��?���?��m��A���@�2��>С�?:cY?�yi>GU۾7pZ����>�@?&R?�>�3��^'���?8ݶ?ĭ�?`I>���?�s?�k�>�0x��Z/��6������p=؆[;�d�>�W>f���xgF��ד��h��u�j������a>��$=,�>QE�[4���9�=��I���f�<��>�,q>"�I>W�>v� ?�a�>}��>�x=�n��Jှ�����HN?SY�?~� ��;[��=K�<���+?�9�>� �=h���5x>��6?��?�h?r;�>�]
��]���nǿ�CȾ�]>��>G�3?�{o>%�{��q�=ѐ۾�)s����>�m�>��8>�t����⽾[��{j�>-�??AJ�>��>� ?�?��Q>[��>/�W��ܘ���D��k�>�D�>57?3B�?k?�u̾� 7�>���բ�Z[\���L>�v{?��"?fe�>,n��E=��om4<(�G�K���׆?E�v?����?P�~?pv2?�B*?�E>9���S����K6�'�>�)$?a����5D�i�)�;U޽l�?S�?d��>t������b��/ ��n��kU?��^?�?�{�{�b�a[Ҿ���<P =*��:� �<(����r>83�=Bry���=��R>ή�=E�c���7�(�<2��=��>U�>r7O��)߽�E,?YmJ������=x�r��pD��v>m�L>�����^?w�<���{�q���r���qU�7�?Щ�?yt�?����څh�E=?��?�?���>y1���j޾J��w&w��}x�ko�A�>���>\�g�c��R}������A����ŽG���|�>���>,?F� ?GP>=�>"J���?'�����&c^�8��7�jN.�
Q�_�����#����I¾�}���>nh��7��>"u
?��g>�j{>�d�>(Ȼ�2�>$�Q>~~>W��>?#W>�4>KS >�<[�н�s_?�u��O�B��<�Ұ�K�4?D�?�*�>�'3������)%�	�>v�?	K?�[R>�^����U�sȤ>��>�NI��?m�j=,�O=�>����ݴ����=�Z��ʺ> c���mp�X`��&�=�P6?N�?�!�:d ����׉�b�����?B�;?L�I�&g��5����g��g>��-O>ncx��x�p���O��/���؆��B����0����<`L?��?P�H��b��i������"�Q�>{��>�$V>
p?�l>���TY������m5�B�����?FX�?��0>��|?�/?[H?B�K?�j�>���>0I��¼�=h�C��>��>�,?�jK?eE?�#?�(?�q=��>=�8�?ھ+"�>�.�>u{0?S�>�V�>��=�O뽮S��n���dľ9�ɽ�?z�����E�x� �B4)=��C>�X?S��Ϭ8������k>z�7?{��>R��>����-����<��>L�
?�F�>2 �)~r��b��V�>���?����=��)>D��=���<�ҺZ�=2���.�=F=��\};� `<$��=���=�ht��<�����:��;�m�<٬�>�?��>���>@7���� �Q�����=�Z>��S>M�>�,پd���(���g��Bz>̚�?ā�?��g=g^�=���=�M�������ſ�����<��?�]#?�>T?��?��=?�#?O>�!��(���:��}���q?�!,?��>D����ʾ�憎��3���?'[?	=a���P;)���¾��ԽS�>�W/��,~�?���D��ᇻ&���j��ڛ�?��?�7A�(�6��y�1����[��1�C?�#�>^�>��>^�)���g��#�S9;>d��>�R?�><�O?y-{?w�[?�jT>j�8�$��ϙ�� 6���!>�@?鷁?��?By?���>n�>��)���97��Fx�������V=�)Z>:��>��>t�>5��=�3Ƚ�T��mB?��9�=ub>@��>а�>7�>��w>Fݰ<��M?U��>m�/��S��7u��ܫ���?���?��;?d��>�ܾ��n�HF��	1>T�?�d�?9�U?F%�j�=�<|Ӣ��BL�4��>���>���>}�>��=���==2�>���>��R�e:ξ#+��*�B�>#w5??!=�'���lt�|ͪ>���=������=><��]�P�3l���Ik>W���FWj�w��;g���[��oҹ�L˾/!�Y�?�zY��>�����=O�a> c>�f,>���=�ڲ=~(���K,>�F��]�=��J�,��;�
����=�+���վ���?�h5?�.?�*d?�I|>�>8 ��||Y>�  �>N?jv.>��I�;���9Ԭ�M���w畾�}߾xt��T'v�����`�>��]��*�=��=��>$�<�݁>K*�=�C=��/��K<�֦<���=��=01�=� >c�=�6w?H�������4Q�[�r�:?�8�>K}�=�ƾf@?d�>>�2�������b��-?z��?�T�?u�?�si��d�>%��5㎽/q�=I����=2>���=��2���>*�J>����J�����e4�?��@x�??�ዿ��Ͽ�a/>�7>5 >��R���1��\�c�b�~Z�-�!?,;;�9̾RJ�>��=�8߾�ƾ�<.=Ψ6>�Gc=C7��M\��͙=��z��;={l=Vԉ>��C>4j�=[���=�I=5��=��O>�]���k7��V,�Z�3=���=�b>��%>~��>^�?La0?�Xd?�6�>�n��Ͼ�?��WG�>&�=�E�>f�=isB>}��>��7?ԵD?��K?̈́�>�=��>��>��,�B�m��k�̧����<Q��?�͆?�и>_�Q<œA�Y��/g>�L5Ž�v?�R1?Nk?��>�U����tX&�D�.�i���E��+=wmr�DRU�O����m�ҭ㽣�=�p�>���>d�>%Sy>��9>��N>��>ũ>�8�<�p�=�،�p��<����ղ�=����"�<�ż���҃&���+����h�;ڹ�;#�]<��;���=���>W<>Ĭ�>ґ�=A��2D/>����1�L���=�G��$,B�G4d��H~��/��U6�v�B>S:X>�{��14��k�?�Y>�l?>���?Au?��>m �.�վ�Q���Ce�6VS��ɸ=�>2�<��z;��Z`�J�M�M|Ҿ���>0ߎ>|�>D�l>�,�#?�W�w=��Ab5�Q�>�|��e��(��9q�@�����zi��uҺ�D?|F��.��=A"~?�I?S�?^��>�����ؾ�90>�H����=���+q��f����?'?���>(���D��l��7۽�7o>Aۆ�P���x���_.�b��=Ģ����>��Ƚ uƾ��I����'6���U� -��O��>�a?M&�?����-����z�>9���[�Ho	?�@�?0�?;h�>BY?���W�����9��<��?���?���?�D>xn�=W���\�>�"	?���?���?nas?2�?�O�>pZo;�r >"��=uB>���=��=�I?N
??�
?|坽"�	�������]��W�<�T�=���>��>H�r>E�=�yf==��=.�[>�P�>��>?�d>��>�#�>��о1s���:?�X!>��V>��??D-A>9q5=�7�!�=�4����8�2�½�>+�PԷ���\nW�l�0�����%��>`gɿ���?�%>OK���"?.����\�9�W>:>Ͽ��-�>�N>=�>��n>U�>�t�=���>�oY>
Ӿ�>���#!�bcC�N�R�k(Ҿ��y>ϛ��{%�ʂ�	\����I��y��K��o$j��/��3=�a��<�N�?ӵ��gl�� *����n>?8��>�]6?�\��Zى��>��>k�>#������ѿ��Q[�+�?���?�;c>��>I�W?�?ْ1�33�vZ�,�u�n(A�-e�V�`��፿�����
����.�_?�x?2yA?�R�<-:z>R��?��%�[ӏ��)�>�/�'';��?<=u+�>*��/�`���Ӿ��þ�7��HF>��o?<%�?wY?@TV��(>��e�>��?6!?��~?V�?�B?�����?��z<��>�M�>��?�_(?�x?I�f>ng=��އ�=��ý8
��,P��%LJ����uWr=כ�>{x�=y�>���=��h� !��H;=-/n=�R�].U<���=��=펕=�d�>T�]?���>���>��7??��8�׿��r�.?�;4=�p������-2�����z�>��j?�ګ?��Y?�e>��B�zPC��>k��>��'>V�[>��>���j�E�`��=$�>Id>1�=G�O��w����	�
���<��>R��>�0}>Ha����'>w!��8�y�ϝd>��Q��!����S�#�G���1��	v�H��>J�K?S�?>��=`t龚]���Af��)?S<?KM?ú?Q�=C�۾��9���J��0���>T��<Q������w����:���{:��s>랾�ҾK[8>�t��fVW�Eya��2M�kF���7���&��=p��h)��Eg��C�=f�>0�ʾ�J1��M��访*P?�_�< X��O�_����H>��~>���>0��:<�FD���^��ڔ=���>+�>,��<�Vݾ`93�y��a=�>�PE?iW_?=k�?."��Fs�'�B������c��oȼ��?�x�>�g?�B>.��=R������d� G���>ş�>���B�G��;���/���$�u��>�8?�>�?^�R?`�
?��`?�*?RE?'�>��������A&?B��?��=��Խ-�T�b 9�-F�s��>E�)?��B����>8�?�?�&?�Q?�?��>� ��C@�s��>LY�>��W��b��\�_>��J?͚�>S=Y?�ԃ?G�=>M�5��颾�֩��T�==>��2?�5#?:�?᯸>@��>K��w9�=�N�>;c?�.�?A�o?���=<�?Z�1>v��>�6�=���>�^�>�?LYO?�s?��J?^��>ʉ<Q������r�wHK��'w;%�I<&vx=���{�s�������<�ÿ;w���ƀ��9����E�i[�����;�>�>O&�>�6��?��=�ƾ�Ir��n>�r<�鞾6��K�B��۱���>%
?�>�>����C=Ќ�>f�>�g���4?� ?^�?� <��d�&�,a@�qV�>�[Z?>��=
Ra�ʵ��x6o��L�<(L{?4�a?¤j�E����b?v�]?���� =���þ��a����g�O?�
?{�H�]ӳ>��~?�r?��>#f�T[n��
��+b��,j�q�=�C�>�F���d�3ѝ>�j7?BO�>�b>K�=.�۾ �w����Q?��?�
�?F݊?��)>��n�%,࿊��FD��mZ?\�>Ī���o�>�u_�BD�������t�.���^���p������)���jH;�7K��:M��=j�%?���?0Z|?[&|?��M��$a����E�����'�m)/��}<��xQ�0_`���l�� оߺY����+�R����?	6I?��&�>��ɾr���v���>�!������Y�<\Uc�G�>숩�R���8@s����'E?w��>Un�>�f*?�2n�Z�-�2(1�O�;��v�їi>"z�>��P>J�>OǮ�q�n�R�J���Ҿ�c[�]����6v>�xc?��K?6�n?�n��*1�l���$�!�4�/��c����B>mj>���>��W����
:&�HY>�9�r���Uw��0�	�Υ~=��2?n(�>x��>�O�?�?a{	��j��kx��1����<�0�>� i?�@�>��>�н�� ����>��l?���>��>�jZ!���{�˧ʽB&�>�>��>��o>'�,��#\��j��Q����9��u�=*�h?���[�`�S�>�R?9�:�G<�|�>�v��!������'�;�>c|?�=b�;>,�ž�$���{��7��{=&?�?z\����)��`�>��#?��>���>Ӈ�?��>8�ľW����?��]?�YH?�@?���>�z�<�����۽5�,��E0=R��>l�\>��>=hG�=j�Z�T��R��qL=f�=c+��kꪽ,��;t��,;��<��3>��ۿ'?M�Eɾ��x��w��^�����	��� �}e������~�h��������/V���l�j����s��@�?)��?��r�}I�7���%�w�j���!�>io�աy��Y��{��K��/��#4��s�#��Q�<�m���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >^C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾r1�<��?7�-?��>Ŏr�1�ɿc���z¤<���?0�@H�A?��(���kP=���>;�	?1\A>�1�@���q��]9�>�g�?��?�L=>�W��}�d.e?�\	<nkF�cl�&�=�0�=�=�>�ǱJ>���>L���4B�2��\[4>�ф>ѣ� �$�]�u��<�\>2<ؽn镽Մ?�v\�f�#�/�>T���U>�T?�,�>(�=ױ,?$6H��}Ͽ5�\��+a?�/�?ĥ�?s�(?:῾�Ӛ>/�ܾ�M?�D6?J �>}c&���t�{h�=x:�-Z��@��'$V�"	�=��>W�>��,�d���xO�%�����=R���ƿ>f�s��-��;\���t�Ѽ�� ��Iǽ��%��ɒ��Or�q`����=�>�MR>՛t>�cM>`�8>��Z?�by?ja�>[gc> k߽~{���e���"���5��|��
��K����6���ݾ_�	����>���ʾ!=�%�=7R�m���D� �h�b�Q�F���.?w$>c�ʾ��M���-<�pʾ_���=܄��ॽ�-̾�1�"n�h͟?��A?������V�J���W�����R�W?P�һ��ꬾ��=^�����=�$�>���=���� 3��~S�h�/?:?��ƾ�
��84>2�	=�v*?/H?X�\<���>+"?�)��_��*J>+<B>i��>�3�>�>〯�L����?2�P?��� ӛ�L��>����S���aF=�f>a4�yռp�l>�6�<����������x�pY�<O�j?�Q+>��H��,P���=�5`>��>l�d?S]C?7�f>#�:?Ys?01�p;'��N�&���dX>9Nv?y�}?1ݰ=���Qaþ<n��xd�>^�?[�%?E1羒���@�yL�.Y2?Z��?��0? >
D��le�g(?SO}?��5�1������ɴ��Х>�[=�s?����˘>�c?�^�R���Z���O��ڜ?&�@1�?Z2>Wl۽�&��+�?z��>(��������|�*�6��&��0�>E߈���Y�6�1�m�= ?�U?�*?꽐�����=�ڕ��Z�?��?����Hg<����l�
o��֖�<{̫=��G"�k��E�7�;�ƾ��
�
����������>Z@OZ车)�>�H8�(6��SϿ��z[оIRq���?���>��Ƚ圣���j��Pu�r�G�y�H�ԣ��w��>4�>����*���|�`�;�;P����>�m���>��P�6k������	<_�>3��>���>�ݭ����A��?{���`ο�������[�X?�H�?@�?~�?z�.<� x���z������F?�^s?�ZZ?����^\�
^6�ÿj?�]��&V`�ؐ4�}DE��%U>�#3?C�> �-��}|=�">���>4n>-#/�?�Ŀض�x������?,��?�n꾳��>��?ls+?�j��6��9Z����*���:��4A?�2>����8�!�.&=�s̒��
?A}0?J���.�]�_?)�a�N�p���-���ƽ�ۡ> �0��e\�9N�����Xe����@y����?N^�?i�?ӵ�� #�g6%?�>c����8Ǿ��<���>�(�>*N>oH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�-�>P\�?��=���>���=�#�� �8��O'>��=�\q���>��H?���>�� >fl!�9�'��_@��TP������F��)�>vab?��L?�U`>�⺽��9�X�!�(MȽ��F��4���4�N�+��ͽ�1@>xD1>��>�z+�{�þV�?_n���ؿ�i��!c'�)14?q��>��?h��r�t����:_?Zo�>�>�+��� ���2�ڛ�?�E�?��?>�׾�P̼|>3�>YN�>�Խ���񊇾��7>��B?�!��A��_�o���>-��?F�@�ծ?\i��a?�%��뜅�|�z���19��fA�=J�??�������>,?��0=��y����:���S�>�h�?Z��?J�?Q�j? /c�[Y����;���>�s?��?�`!�<�Ǿ̥>�H�>�J��xJ��U����d?�~@`
@�__?D���ڿ����Y��ѭ�߶=�(<��Y>�p�(�=�q=�����Ww>���>�|y>��d>��N>B�@>>����W �ah�������K��.#��	�״a������~�[�X���M�����ѽ�M��R�O����r���F	�=�Y?�@?�Fa?W��>�-ʼ�0*>���e
/���R���;Ww>��0?��K?CM'?�չ=2��C^�nWj�dߵ��������>9>y��>0`�>ު�>l�ٺ%�f>��L>�<�>z��=�K�<�#�$�A=�A>�:�>ˑ�>L�>�C<>>Eϴ��1��f�h��
w��̽/�?����Q�J��1���9��Ħ��Ki�=Rb.?|>���?пc����2H?����r)���+���>i�0?�cW?�>;��\�T�@:>-��Ȧj�"`>�+ �l���)�w%Q>dl?�|s>t��>�4��7��M��������>e�5?�}��#+�B�q��K�W�Ҿ��b>:�>���;�Q��x���6|�ub�};�=��;?��?�۱�{���\���sb���2>�r>�6&=S��=|�M>��X�^�i�4�A�=�A>��b>V?j�2>ӏ�=�.�>���e�M�P�>�pD>W�&>�>?��#?�Y������〾6)�b7z>~�>���>D�>�cP����=e��>d\b>&>���}� ���IB���T>�z��U�_�l�q��z=]���a��=dq�=�B �X�6��4=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ
i�>"x�eZ�����U�u���#=r��>�8H?lT����O��>�)w
?�?�_����H�ȿ�{v����>?�?e��?��m��A��c@�ׂ�>��?agY?�mi>g۾-cZ���>'�@?�R?��>9���'�p�?�޶?���?aI>���?�s?�k�>�0x��Z/��6������p=҆[;�d�>�W>e���xgF��ד��h��u�j������a>��$=,�>PE�Z4���9�=��I����f�<��>�,q>"�I>W�>v� ?�a�>}��>�x=�n��Jှ�����CM?��?*��n�<2<�P�=c�9��?�)?� �WFξ�<�>Q�X?��?�k]?B�>o�����3���|���я=VkY>��?�%�>7⻽��>]]Ͼ>�k��<�>�R�><e�;�=ؾ�f��b8�͙�>Is&?K��>#�=�!?�?h�g>ʁ�>�xv��?����K����>��>��(?$T�?���>	:�=�7&��u8��B�Z�siy>{ z?�-?~S�>�`��>���*I�=0Q��G;=���?�N�?3j��#?f�j?Z�)?��?��X=(2�=��^���/�'��>7�!?ݬ�6�A��J&����م?O?���>����~�ֽ�׼����M��l? !\?@&?]���(a���¾��<�:%��U�� <�LB�$�>�}>l���=�.>��=�'m��)6��f<X�=�g�>���=tE7��z���?,?�fH�僾Ę=�r�]rD���>PlL>����,�^?O=���{�a��^x��LU���?S��?Yo�?���Q�h�J=?�?��?� �>@6���X޾��ྜ;w�hx���8�>���>^l�=�侗���ϛ���D��4�Žx<���?#q�>�4 ?{R�>5�t> �>n��=,��6�� �(�Y��3�RR'�4!���Kᐾ�n1�Bg�kҾ9���K$�>y���-�>�d?L�\>�m>��>{��<1�>�H?>~,~>Zi�>�4>1�'>8d�=>4S�i<ڽʖ^?9&����<���-��lh?��?Yg�>��Sˣ�PM��r�>��?B��?I�>����t�0�V�>Ӕ?3z���~?�%<�8�<M\����lUR�T\=��N�ҹ>3�͂�\Q�S��=uN?!�!?G�!�9�'���$��+��� �?�i2?C�]��F����[��I�=�7>��*��͎�N�&���d�?�������;���1���e���\?RK�?ݵ0������"�'���P�0�em�>�?v��>�	!?��>>����N�K���.��ï��Y?2]�?>9h>�]?g7?��%?�6<?GJ�>^<�>Z���`�>i&��I5>;a�>�5?:G+?S;(?0� ?S#?��=�xC�n��0 �ǡ�>�'�>H�?m�>��>~��=�<���;W\/��S��m��:�괼":���Ž䚻��M>>�.?X>�c�8�������k>zQ7?Y1�>���>�S��s/��U%�<���>��
?{�>����g�q�<��7�>ˍ�?�%���<��)>�l�=����?��z�=�Zȼގ==���V8���!<r|�=-��=�~0������i�:G��;^H�<� ?]'?@��>�>(O���7 �a]����=��\>�LR>/C>�ھ>�������g�zw}>"�?�Դ?Pg=��=H��=f���/��G�ݢ���=6?�2#?W T?�z�?ԭ=?�~#?r2>���0+��D����s���*?`",?9��>r����ʾ�憎�3��?�\?�=a�F���9)���¾`�Խ>�>�T/�r&~�����D��x��=��+A��F��?@?RA��6��辍����c����C?��>wa�>��>��)���g����@;>Ē�>�R?�#�>��O?�<{?��[?�gT>\�8�n1���ә��J3�Y�!>!@?���?�?|y?�t�>��>�)���zT�������4ႾDW=?	Z>j��>�(�><�>-��=�ȽzZ����>��`�=��b>/��>���>��> �w>�L�<�VN?c.�>ÿ�Q��+���ȿ��&7
�%y?<�?�%(?��%>�l���X�9���@>uf�?��?��??e�нL�>m5~�/�ܾ�������>A��>���>�'<Yvd=�w�=k[>���>Z�ؽ����+�0��f?�dK?���=i���]v����>�J}>���=�t�<���ݾ�ʾw�>Lb����=]-��E��zB�������뾴þ��/�V��>�b��͏M>�(S;��=�5�=����4�v>��E<Z�=RV�=��<�+{���k�<Oqs=��(��>�q>F�;�Xɾ��{?$�6?�W?E?qm�>,�->_�N�ݛo>`�罟�?�?>$��<�ʔ�3��wn��9f����YC���������g�>�S<<L>M�=��=Ce���>�B�=L��=�<���<���=*�= �Q=��=->��>�Jw?d���p����P��׽�9?F�>,{�=�`����>?��C>�_��gq���a�|?���?�\�?��
?�(g�I��>(�������m�=��~9>���=��3�5�>NRM>���ﱛ��什��?m@1�<?������ο��6>�N7>�>NrR�iZ1�0(Y�Y�]��wX�:+!?ĳ:�8;�̄>�=e3ݾ(�ž��/=ׇ9>�f=��v�Z��'�=Vׄ�w6;=E�j=_�>owB>U�=����
��=�xK=�=7O>��F���4��m-��5*=���=��`>r%>L��>K�?�[0?�Qd?s.�>1�m�CϾ;9���4�>���=`9�>b΅=|xB>㗸>��7?�D?B�K?,}�>�։=���>���>��,�ٵm��^徖���ʙ�<1��?�̆?Ѹ>��Q<��A�_���j>��VŽu?P1?Vg?Bݞ>(����࿮1�Ƚ"�X��C��/��=uɊ��cZ�Jk�������sU�=vE�>W�>�[�>�s>+M>>�i/>�3�>��>��k=��=UM��e$�s���[}<�WϽ~n�;�!ݼ
� ����;�7m����^{9�ۼD-1��4\����=���>4>���>Ȏ�=j���1F/>������L����=�J���*B��-d�A~�_ /�~A6�'�B>�/X>�l��%4����?��Y>�_?>���??u?R�>0 �a�վIN��Z@e�VS�"˸=�>�=�Lw;��V`�6�M�:yҾg��>lߎ>�>~�l>�,�C#?���w=��bb5�o�>�|�����	)��9q�@������ei��gҺ�D?�F�����=r"~?�I?\�?��>?��نؾ-;0>�H����=g�p*q��h����?'?���>�쾚�D�rD���ս�ײ>=�N��>u�⌞�5}8��0�=�����>�q�-�Ӿ��?�g���B9����I�K̑�u�>�S?�3�?� �����:Z��/��	�Ɋ?i�{?��>�-�>�?E�Խz�����s
�o��?���??l�L>�ͺ=�G�����>��?�E�?���?�~r?W�<�]�>~8׺��>�0�����=e�>9�=S��=b?��?%�
?M����
�����m�9!Y�&��<���=���>�(�>>s>���=�hi=�o�=K�Y>�>h�>��`>ū�> ��>��i���:)?��>�ь>�/?�&{>=e�ɽ� �<7鎽�>1��L$���`ӽhD�<�ve���=�-@���>�ƿé�?�9F>����?@0�4s��� S>�[>��ֽ	��>�?@>��w>���>t��>��>���>g�">�@Ӿ[S>O��^U!�:3C��~R���Ѿ
Oz>Y���_�%�����|��dMI�Bo���c�9j��-���6=���<�K�?QT��x�k�-�)�r����?�K�>�6?gÌ������>���>q��>�]������ȍ�p��?\��?�;c>��>D�W?�?ؒ1�$3��uZ�'�u�p(A�/e�U�`��፿����
�p��.�_?�x?-yA?$S�<:z>L��?��%�aӏ��)�>�/�$';��?<=x+�>*��)�`���Ӿ��þ8��HF>��o?:%�?sY?CTV���0�_h�>��?��>�gs?�?��??�{$�P�?�>��4��>DD�>s�;?��2?�+?dҘ>z2L=$%(��'>�B�Î��b[ܼ�P��Em<�U���M>�=;:>��<�/=>�T8<J�ɼ,�-=�8)�A��=_�=&6�=���<d�>Y/]?���>��>��7?����48�hެ���.?�4=?ā�e����]���S�[(>�"k?m�?lZ?�e>f�B�y�D�nY>){�>h'>�I\>�ѱ>�b��C�8��=�Y>U>���=�UG����`�	�%��<<K>?8�>k�?ؓ6��>b�����?�>���;��1u� R1��#�����y?4S?��&?�>���K�E��6."?M�B?k�>?pG?�_�=]�߾H�)��-�v���~�2>�6>��ȾȀ�F���E@��_G|=ň�>�W��ɳ����\>!
�[�ܾ��k�T>I�:*��M=J��[=ڭ
�w�վҢz���=��>/���c!��*��6���dI?��v=�����S��ɹ�(>	�>u	�>��M�㜋��y@�����=O*�>�Q<>uJ���s���G�:�����>`�E?��^?y�?�Ň�]�s�t�B�k���?��������?���>��?��5>9��=᬴�Qq���e��lF�@C�>Ɯ�>�N�XmH�����I@𾺅$��߇>��?m!>�_?�gT?�/
?�^?^�(?1?_��>�Խ����E&?i��?8=�ֽj�U�s�8���E���>Ux)?Q�B��˗>�?�?��&?�DQ?�y?�>s�
�@��`�>~�>|�W�FD���(`>�J?aҳ>@jY?氃?��=>�F5����H��� ��=.V>��2?XS#?��?�V�>� �>�+�����=���>H^c?�?��n?_>Ɨ?�H9>���>�"�=;�>w��>L�?�SH?��l?�K?.�>N�<B�������In�$(N���<���<?��=郬��1&�7���%�<�p�:9��O����Ǽ�$A�	�¼˔4�jb�>jt>������0>��ľR����@>)闼T���n��|�9���= ؀>L�?�X�>��#�> �=_��>�>���-�'?֭?>?���;�ab��G۾n�K����>��A?�G�=��l�Ĉ����u��j=��m?^H^?@W�8�����^?�h?��Ǿ��D��9�i���zپ�Y,?�c?�z)����>��p?v Z?W{�>���p?i�4d��GD����ھL��=�*x>�o���a�]2�>J09?K��>ni�>���=����~Z�ȏd��Q&?���?@��?�J�?Q�|>�R��!ݿĉǾD왿a�k? G?���<^0?��?^@��)@�����j)8��ݾ����Rվ|���#o���������<�O<?�6?�?��G?��$���%�R�`�������<�(�
��L"���5o��� �>Q�haؾb�^�Ĉ�;�=k~��OA�Uo�?v(?
-,�G=�>+������M̾�(C>����������=�f���;=�+V=[�g�=.�7�����?��>�I�>�k<?3q[��=��U1���8����d�3>��>D͒>��>��G;n,�f�潒LȾ�˃��SνΧv>��c?�`K?�An?��k(1��`���}!���-�OG��K
C>�>���>q
W����B6&�:t>��@s��^�ck����	��|=�w2?�;�>�ۜ>1D�?�B?�j	�A����w��=1���<2��>�i?�J�>�K�>��ν�� �\��>�@t?X��>R�>�����B�k�e���H��$8>z��>8�>�s�=��M��g^�����Z2K��0>W�C?��~�v_�O��>��A?�J���������>�<��ڛ�>�*;�q>���>)W�=rDO>��ؾ#F�����k��m )?��?+����*�[�}>'B!?���>0�>pC�?�Ϝ>�\¾b��:��?��^?��I?t�@?��>�=ُ��ɽ�W(�;�*=��>~<\>9k=/��=���tZ�|]���A=�[�=�߼V����l<�ش�l8<���<��3>�iۿC@K���پ����"O
�%��k������'����9��1
x��D��(��U�
?c�����Om��j�?��?Fړ�r������`���w��ّ�>~q�����/�� 4�6����ྃ���SN!���O�Bi�d�e�O�'?�����ǿ񰡿�:ܾ.! ?�A ?8�y?��0�"���8�/� >D�<�,����뾫����οK�����^?���>��t/��u��>㥂>��X>�Hq>����螾x1�<��?8�-?��>Ǝr�-�ɿ^���bä<���?0�@;vA?��(�����iU=g��>�o	?��?>R�0��*��ΰ�,y�>�8�?Z��?֜M=O�W��}
�{ee?���;<�F�p����=���=�{=.}��BJ>�8�>�/�2?A��ܽ��4>��>�!����Qi^��<��]>dԽ�g��_��?O+>���k��a@�c�x�(j>�C?��>�$�:DY8?��*���ҿ�o�D�c?d�@s�?�z0?�1ɾf|�>#ϾH�=?��#?,5�>I��bp��n�=���<@ߑ=ҠӾ�tS���=��>&�=&GR��	�wk �[=�c�<�1�A&ÿO'�Ş��Q=o�?�B��
;۽�T���żnZ��(�p��ӽ�m�=���=�J>Q{>`P>H�7>�U?��i?}]�>�">�7ν��h���žP@���T��77�מ����5�"G��)���޾����H�H=���߾�"=����=U2R�A����� ���b���F���.?��$>��ʾm�M��=-<�gʾ�����F��0楽_1̾o�1�'n�qʟ?T�A?���V�}����La��:�W?Q���O����=���ʣ=�$�>uy�=���"3��S�gw-?�?�)�����Q�>'e%��R=^5?.5?y=9<�>`�*?��������;>)>%�>���>��=g����0�Z�?��X?�.�Z����j>:T����>�:7�=Qd�=)�F������UM>��=*���-a廼!��=Y(W?Ǜ�>��)����a��V��\==߲x?��?	.�>X{k? �B?��<;g��K�S����cw=��W?r)i?v�>�����о<����5?�e?f�N>�ah���龮�.�VU�$?I�n?�^?[{���v}������'o6?��v?�r^�{s�����*�V�i=�>�[�>���>��9��k�>�>?�#��G�����vY4�#Þ?��@���?-�;<' �?��=�;?{\�>׫O� ?ƾ){��������q=�"�>���lev����3R,�B�8?͠�?x��>��������3�=�C��U6�?FW�?�����SQ<�T��>k����H��;�`�=i�:���4��[��8�� Ⱦ�]
�;-���@��)�>ƃ@�b彞x�>P4��L⿝�пi���Iվ��z�E9?�Χ>5Fݽ�ʥ��Di�ڟr��lC�l�D�T��0d�>f>���s)����{��J;�3V�����>җ	�v�>��T��p���矾Q�*<��>[�>%@�>a�����?�����Bο#���,[���X?�c�?�@�?lO?6I<�v���{�~Z��BG?'�s?_>Z?�}%�a�]��-8� �j?Z_��xU`��4�aHE�nU>�"3?�B�>S�-�P�|=�>S��>�f>�#/�w�Ŀ�ٶ�7���X��?։�?�o����>x��?xs+?�i�8��m[����*��",��<A?�2>���*�!�$0=�LҒ���
?~0?�{�V.�[�_?-�a�c�p�/�-�w�ƽ�ܡ>#�0�`h\��e�����We�2��Dy����?}^�?��?ݳ�� #��6%?��>q����8ǾY�<��>�(�>�(N>_A_�۳u>����:�wg	>1��?b~�?Mj?㕏�����}U>��}?ͻ>���?	>�>3:8=� ���<�Po>'i>f���?8R?I��>���=͕L���*�`p7�3J�Щ
���;��6`>d�Z?R�R??�>?�޽cM�����ύ���#�{?A�%�)����i�ٽE�0>\b:>�5>�BԽ������?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�e��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=7M�>Μk?�s?�Qo���i�B>��?"������L��f?�
@u@a�^?*�ӿ����������h>dd�=��|=<�3��'?=�4^=�E��d�F�B >���>nw@>��@>zM<>���>-��>I��'�Pˣ�q+���K�W�9��a�������(>������l0��n���Tƽ����lĽB�<��=�4T?"�Q?F.o?�2 ?3���@>����"=4y �2�=8P�>�O2?s�J?-�(?�=r����d�#���e8���6��{C�>��L>�y�>���>|��>v|�GmF>�f?>a�~>'�>�y/=��ٺ#h=J�N>�Z�>�J�>��>�I<>r�>Eʹ��1��e�h�	w��̽��?}��x�J�r/��E5�������t�=_.?�s>���@пl����/H?=����)�o�+���>e�0?�cW?ů>/��j�T�b>>��� �j��j>�$ �Jvl��)�F-Q>ki?5�g>�0v>�3�o�8�MEQ�����S>}>�?6?7����7�K�t���G��ܾ�M>;ٽ>�S��B��������i���u=]:?T�?�]��H����t�.��R�Q>�[>D-=�Ʈ=f-O>)Pd�3�ƽ�HG�a)8={�=�,b>�[?�4>>��=�>^N�����V�>"�>dam>��;?��%?V<=S7��iW���6�o�D>r�>}sf>�2�=��P�^�<���>���>1I�=�}���A���O��@�>lPڼ��q���޽���˕��9�>��=�f��@c���=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾNh�>|x��Z�������u���#=T��>�8H?�V����O�i>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>:��?�gY?ooi>�g۾<`Z����>ѻ@?�R?�>�9�~�'���?�޶?֯�?&�>_Q�?�xl?��>�᥾b�D�kѨ�#?��|o=:��=��>E�=����,�\�M���w�������FK�I�=v8�=�ݵ>�!������#���&=�j��G��e�?�&3>��V>���>o� ?��>o�>�5�=+�2���۾�C��$F?�K�?��<�r��S��-?93���n�?�3(?��=�?���>��S?*n?t&?=�)>���GU��q|Ͽ�<����۽��P>�M�>E �>������l>�҄�*�;�q�>=/�>J >�U�P�Q�V�:>��>��;?k�?S��>K� ? �#?��k>�ϱ>u
F�g��ӻE��>�>���>�k?Ub~?m;?�湾�4�����1᡿�u\�n I>k�w?�?�>ξ��xt�����1�B� g��n�?�hh?
pὫ�?셉?W�>?״@?�he>����Nؾ�
��P�}>S\$?�y����E�(�7������?m�>���>�A��	��/1=�,������?��t?�!;?��羟`b��ۢ�3�=}���K7����K=��>+��= ��\>rF>�0�=jꁾ�}=���;i��=�5p>�M�=hH*�`ʽ(\1?L�>���Ż��@��V*����=�_�=䗶��$@?um��;t�*���}x��<��<چ?���?���?~�
��?[��s"?ކ�?�%?���>0��$��zDȾ��5�U9��0�)�KO>�7?�)꽀�8��¹��ެ���Y��Hl�:���=�>��>r�?Z: ?�Q>Yβ>=-���&����n��*^���kh8���.�.��p��f�#�^g��^����{�u��>gh��nm�>;�
?� i>��|>��>�a��s��>��R>�~>���>��V>@�4>s�>Z�0<��ʽoKR?����E�'�ĵ����d1B?qd?�3�>��h������n�?~��?�r�?:v>"~h�w++�n?W=�>B���o
?�Q:=7���z�<@T��)���2��S��4��>	J׽� :��M�-lf�Dj
?/?���w�̾�4׽�$��j�=���?q#(?�g+�4=T�|~m���V�>\T�*��cEe�����K$��jq� Ǐ��������,�(��=�K)?��?"e���7�$���g�h��u>�c�e>���>���>\��>�X>���S�1�*�[�I�$���&E�>�ow?S�>��B?�9?vkH?��B?�h>�\�>,愾�^?�"=��>���>�9?%�*?��#?�
?��%?��\>�j�`2������j?�"?�"?ޢ�>�A�>������꼮��<m`9�����\	��;u=?I^=�0��P#��	1=�bD>�F?|���7��g��7n>	7?q�>��>P���怾���<x[�>3�?�L�>`P��+�q�����>�?�M�n�=��(>��= �{�.T;%-�=t���#a�=�D���7��<�
�=��=�SY���:8b;�X�;��<�?�V+?�U>��`>�O1���Q���F<:>8->n�=��`/��-���cs�Z\>>숋?��?$�H=���=	�=֗'��G��-������G=�U�>�?s�K?2�?u;%?a8?�M>i���栿��������?�,?袑><����ʾ����ъ3�Q�?md?� a�{�)��P¾	EԽ�>�X/��#~������D��0������ՙ���?i��?_N@�A�6��_辷���$@����C?s�>�w�>�&�>J�)�?�g�F�Go;>���>!)R?�>N3?�?��b?�G�>_Q3��5��I��4�t<�2/>:;?��~?�m�?��k?���>���=�ȿ��ʶ��ޫ��޼�ȍ���<p�=/�k>8��>j��>m�=��B��V-�3�\�ڝ>���>�-�>0��>��>=��>y>T�L?�?v$�c�,�V�������>d���e2?�U`?
k??(?>;;��Vp���޾�?=t�?���?��?p;B��y�=�|�o�Ͼg�#�T��>!�>�iQ>;�C>1�s>R��0>��?*/�=�Y�S���!a��# ?ql?��������<J�Q:=�f0�/��=Gҗ�+��z �=�&j��t�Wי��vཟ%	�ƿI����������}־����c?&#�=�!p>�>v���>k�>�<>��=�$�������y=������4�߅̽\���f���=��=�z��^1?��??�5??F?��L=�^=� >���>v��;��?�f�>R}=�[о:�]��s��|��EH�ž�(��w�jvV>y�=F�>�)G>s��+�۽]K��nB���S�=�dB=s��=>�=,�l=5I�=oL>8�U>�N>�k?"汾�ښ�Cɏ���	�-�b?%(F>y����J����>=�n>����}]ȿ.i�2��?@l��?Ù�>��ͽq�>�z��235�so��X�	��>�0J>p�
���K>d?��\= ���������?��?�3?V����譿8�>Df8>�>�AR�3�1�B�^�ec� 0Y�b�!?��:�\�˾Ά>��=J޾�ž��*=^L5>��^=�a�ͣ\�[��=O�~��b==qxp=Q�>{BC>㍺=&R��i2�= �H=f�=RwP>�G��q7���+�Z�4=���=M{d>��'>Ւ�>��?�c0?-Yd?<�>n��$ϾO<��XI�>T�=F�> �=0�B>��>6�7?	�D?8�K?!��>��=��>��>�,�߭m��m徥ȧ��<8��?ʆ?���>q4P<W�A���[X>�cŽ�s?vM1?0k?u�>�'��̿@;L�������V��������tC��i#>�����ֽg@>��?�>t[>�v>���>�&�>��>9�>>?��=�;�=W�[=�;P����zC�<�ED��0>D�k>h��<��a���r���Yѐ<�K)�3���p�C��=2��>+<>Ȭ�>���=����C/>踖��L����=�G��d,B��4d��I~�W/��V6���B>k;X>�}��;4����?��Y>*m?>���?0Au?6�>� ���վ�Q���Ce�AVS��˸=c�>��<�{;�[`�~�M�G|Ҿ8��>��>��>7�l>T,��<?�&�w=�⾘p5�p�>�i��_��?�.@q��<�������&i��j�V�D?�8��_��=�)~?�I?���?hx�>�<���fؾ1�0>���T�=����q�⓽��?'?TK�>�v쾔�D��>̾�Q��@��>qI�OP�����M�0����෾q�>�����о%3��f��������B�LLr�4�><�O?��?[�a��T���SO����Hx��WZ?�tg?��>�<?>?�:�����}���z�=f�n?Y��?�=�?�>��=խ����>�7	?�C�?n��?WWs?�J9��S�>�;��>#K��:��=�
>�u�=���=��
?�7
?��
?�K��d�	������S�^�;C=(ީ=31�>o�>'{q>2D�=��]=m�=�Z>�*�>D�>�_d>9H�>��>�Ჾ����� ??�>��>!�>?ê>6�=Q��W��n��RK-�[���
����d������k=��;g<�>�ƿ��?Ks>���G?�g��Ƶ�`3F>g44>�7�A0�>]�>�U>�s�>#Ţ>�N>߶w>դ>�XԾ�>�p�� �*�B��.Q�Nо>
{>�ޛ�A(����ڏ��G��˵��q��i�����-=�g�<���?
���>k��?)�����	?�,�>Nw6?q���T·���>2+�>�[�>4���X��tb����N�?���?��>�ک>��U?��?Bk���N�e]�I#r���o�N����J������\��H���)�
�]?��?@R?�%7=J�>Bܰ?8�s�G@3�`�
?S�߾��t�AV��;B�>�E~�<E�SuоF���8����>���?q��?���>N���%e>+���$?��S?Se?z��>�,�>�v�>h9D?,%F>>�>�O?.pW?(�A?��>VkP��,;0�s>�Q�>���.\�z�"����{��:/p>�Pr>Q�>Y�=��=�>q��Q�<zG���^���e�<�<�����F�<bwQ=�ɦ>��]?UL�> ��>��7?P��w|8��Į��/?��:=�u�� ��m������h'>��j?���?�KZ?Mvd>�A�UC��>
[�>?E&>�[><�>���VzE��=�>�(>���=kGL�����w�	�Co�����<eM>���>y8|>H(����'>�z���&z��d>��Q��̺���S���G���1�E�v��T�>�K?�?ķ�=&Z龔2��Hf�}.)?�[<?-PM?��?O�=��۾��9��J��J�)�>9�<9��m¢�0&����:�}�:1�s>4��͢��I�b>۟��D޾K�n��J���羀KJ=T���X=���<�վ�����=�	>����6!�����Ϫ��
J?��i=e+��X-U�F����>7֘>奮>�9�v2v�Il@�o���{�=���>";>�l����G��P��M�>��F?�
O?A'f?�a��A�u���,�-�
�2���&Y=Ru"?�;�>�n?�)#>���<h�ľ��!�����FW���>���>Է�	zU�'m��B¾�����>s[	?��>-�?%C\?�
?�
Z?��!?�?ޤ�>.���1�þ&?�e�?⃆=��ݽGX�dF9��tD���>��'?�:���>Q?��?R�%?w�O?��?��>���A��b�>�ԉ>W�dT���c>6�I?�=�>[?�p�?�?>�3�SF���D��H��=cz >�r3?qO#?�?���>���>4z�����=��>�sd?�.�?Y�n?��=�k?n�6>F>�>�+�=?�>1��>J?��L?I�q?�XJ?��>i�<vY���8ý�-~�	7W���`;z��<ث�={OԼ9�^���ɼ��<"5<���:������qOQ�%�����';!N�>�s>2���h1>6�ľ�v���HA>誟�4㛾%����I:�^�=���>V?���>�#��=8��>��>���6(?*�??�8;�b��۾�K��C�>�B?e�=��l������u�w�g=a�m?&r^?ȂW�2!��ԟb?��]?i��=�[[ľ�Od�����O?wZ
?#fE�4۴>(�~?ީq?�B�>Q(f�% n�&����b���m�?�=_��>�@�g;e����>r7?��>l�f>5��=��ھ��v����cx?��?��?*��?�o+>�m�~�߿�������@�?/4?y��ކN?�	G>��������(ʾ�S"������^���ž^z �1����	ɾ�-I�P��.Q?�s,?�Uh?��\?��������G�H�z�䌍�F)�0r6�dC�Ԏ/�[�=��d��ݾ`���S3��*��>�x�B�[k�?��'?�I3�m.�>�W������ʾ7�A>Š��r���i�=�_��h_3=��L=��i���0�N����!?1��>A�>��<?#]]��=�W1�T18�����->�ʟ>�ړ>/��>N�
:!`.�A
�fMʾ�愾��Ͻ��x>sOc?P�I?�>l?����G2��+����"�j�V�KΡ�BnI>�V>ֵ�>[D[�8"�$�&�x�?��Lt�y����/t	��J�=S�0?+�w>c?�>���?4?����-����u���.�	\�<җ�>�eg?o��>4��>�佈%"���>��o?*q�>���>jJ|�"�'���u�~�?��I>c��>�?z�l>�)'�R�b��(�������8�9��=�gD?����	∾ ��>��G?˭R�d@s�p��>64-���&�?�i��>��V
�=�?@�U>S�>�߾�K<�}I���OȾ�8)?�??���ߏ*��}>�!?��>�}�>>�?�=�>��¾U�9��?��^?
J?�A?���>�=-R��*ɽ.'�EW.=(ׇ>�[>(Tn=��=�(�V�[�����>A=�=�uͼ������<�B��i�K<���<xz4>�nۿ^MK���پ ������ 
�@����W��O�������x��u2���x����X)��`V���c��Ќ�n�l�s�?�$�?꓾��Y���xz��3c��;�>��p�u*~���Ι�R�����D㬾nT!���O�&i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾u1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�|A?]�(���쾫V=���>]�	?��?>�Q1��H�G���kV�>J<�?���?�{M=��W���	�M~e?�D<�F��)޻��=<�=�E=��єJ>ZU�>4}�{QA�q>ܽh�4>�څ>�j"������^���<��]>]�ս	7�����?�sZ�Z�f��0�>Y��:9>��S?4W�>�=��,?�F���Ͽr�]�'`?AP�?l��?��)?�ҿ�(��>�qܾ��L?.5?oB�>��%�C�r�ӫ�=@3¼��%��0��T����=&��>�C>|�0����v L��>e�]~�=5f�#�¿�{!�۽��*�=�83=�1�~އ�I��J�X�ͽ���}����q�=갌=ӈ#>�[>��*>�R>bX?>�i?HD�>��>��ٽ��h��y��b<H=P8R��D齀z��[�0�̾���p^���UR�zA��"�� =���=�6R�a���>� �^�b�$�F���.?�v$>��ʾU�M�Ǭ-<:pʾ=����݄��᥽.̾E�1�C"n�F͟?��A?�����V�"���V�	�����W?�O����9ꬾ���=,�����=�$�>���=6�⾞ 3�o~S�4x)?0D?�����H��9>�7��k|=ON0?�R�>v@5=��>\�0?��uD����>>TN>��>V��>�-�=p���{t�K�?XX?	yȽ�Y���>�؛� I��!:xnM=*�� ;3'�>�/�<%f�����~���{�=&W?���>��)�h��Z��]�<5==��x?
�?�)�>pzk?K�B?66�<�f���S���+cw=��W?�"i?ѥ>����T�Ͼl��/�5?L�e?��N>]Uh����G�.��U��&?r�n?ua?�̝�Ay}��������m6?U�v?'l^��t�����y�V�%>�> U�>J��>��9��c�>��>?�#�H��L����V4��?y�@c��?1<<�2����=$:?�e�>�O��Lƾm�������<�q=e�>/����Yv����`,��~8?���?1��>g���'���w�=S[��w��?�<�?	��>c<F�J�k�} ��ԃ<�}�=l���:#���8���Ǿ$�
��%��E��B=�>�J@/�����>��6��]⿘]Ͽ���"-Ҿ؍s��'?�]�>S9Ͻ�R��43j�
t�H3F��G�%��� ��>�_>n�Wƙ�{|y��:���{��>�+�b�>x�T��T��>া�W�<��>���>��>�ý޽��?L���~n̿�N��w��"�X?��?c��?�M?7=��W�*�|��?���oF?cZu?e	Y?G�C��N]�XѼ$�j?�_��xU`��4�oHE��U>�"3?�B�>T�-�A�|=�>���>g>�#/�w�Ŀ�ٶ�:���Y��?��?�o���>s��?ts+?�i�8���[����*���+��<A?�2>
���?�!�;0=�VҒ���
?G~0?D{�g.�c�_?�`��"q��@.�ǽZ�>w2�V�^��j �z��e��0���i{��ѭ?n�?kE�?���@#��$?���>�%��$/Ǿ,��<�>��>aRQ>TV� �s>f��,�9�e�>�*�?�-�?T�?A���צ���>*~?���>d�w?��	>�5�>d�=�־��u=��K>\��=|�}=)�?��S?�� ?�&>K�D�|�$�9�F�1~I��M�Di=��B>
�Q?1B?nOW>^�3j�;���s����:
�v0ܽ6/#��0���㼉q+>��!>I��=Qa������?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?oQo���i�B>��?"������L��f?�
@u@a�^?*��ݿxW��Γžk1��d
�=ڭ�=�80>v��fh�=���=��L�?-G�R!>N§>9�b>�!b>�F>�}[>|�a>yy���H��i��4p����7� ����/��9���ރ�i�"�C��\J��|S�=֞��8i��D(�B=��fn<CF>H�S?�=H?��V?�x�>�ؽe,>����!=m\˽�X>z��>�/4?�	D?Z�?�*x=3���jg�f��[������_��>$�4>���>\�>w�>�ҕ=�[>�?2>��r>�
>إ=0h�<�7$=��Z>�4�>�s�>?@�>�C<>ȑ>Fϴ��1��g�h��
w��̽)�?����L�J��1���9��ষ� i�=Qb.??|>���?пc����2H?!���x)��+���>��0?�cW?<�>%����T�a:>7����j�3`>�+ �ql���)��%Q>}l?j�f>�+u>��3�e8��P�y����i|>.6?y涾�9��u��H��Rݾy?M>[��>NtD��m�#�����{�i�uP{=Vs:?�?�*��,۰���u�J0���WR>�3\>M=�w�=~gM>2c���ƽ" H�Jq.=��=�^>JH?�/>�L�=�Ϟ>�痾ǝ\�ښ�>rM>��3>��??�4&?(Qq�;�b��hw��~-�F�m>���>y>L��=x�Q�C�=K��>��j>rѼhh������6��m^>^5��zk��!s�*v=l;���\�=�܋=�c����2��H=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?,�h>�R�?Zf?�	�>_��j=�-����N���N+���=ӣ�>�z>�ﱾM:A��׍��뇿�By�E/1�)W�=o.�<�V�>j���1����'=?�[��Z���O9��s�>49Q>�I>��>��?�v�>��>-h�=��`������J���MJ?��?�g��Gn�pK|<�nm=R�S���?[�0?�;4 ���>\?��|?JRU?~�>B�>���|��RQ��[� <G�A>��>M��>�����L>F����(5����>��>� R��;̾��|�����0/�>!?R�>W�=ؙ ?��#?��j>�(�>IaE��9��0�E�?��>���>�H?�~?��?dԹ�qZ3�����桿��[��9N>V�x?�U?Uʕ>M���񃝿�fE��@I�����h��?�tg?ES�,?@2�?��??]�A?�)f>'���ؾ6�����>��"?�:̽��F���.���,�?\,�>TJ�>�̽���)����%�p�wR?�h?v3?v���'ea��������<�毻�=�f�h��'�FH>�F>�������=sH;>HB>�)`��FG��ں���=ꎏ>=m�=� ,�*���~h.?|ͨ=��žԒ���X��5���->y�5>����S;?t,�"�p��>��V����K�"�?���?X�?z���V_���,?H1�?u�,?A�?W����n��#EҾR��}��j��K{�>��?���;�����Ч��b�����/����>���>�?|c ?<BO>�_�>
'���'��3�����^��]�=l8�9�.�2��}���~#����'¾��{��M�>9_����>3�
?wBh>��{>��>�hȻI=�>R7R>�~>fl�>g�W>�
5>��>�<2<ѽ�KR?���D�'���� ����2B?�qd?*2�>i�ɉ��#����?���?Os�?l<v>�~h��,+�Hn?�=�>����p
?\:=��G�<�U������3����ī�>�I׽� :��M��mf�!j
?]/?����̾�<׽=���zi=pe�?�&)?�*�A�Q�[o�W�W��<S������i��y��*�$���p�����^��T%��(�n�*=��*?4(�?���eGج��yk��:?�b�e>���>Ɣ�>nx�>uH>��	��1���]���&�U
��t��>xY{?�><�E?�:?piJ?�F?#��>Dz�>������>Q�<@ӥ>P��>�<?��0?�|*?'�?�!??�^>����x#��Lrھ�?��?Ok?�h�>��>]���򋽜t6�9hA�7�|�Nᙽ;��=+��<�o׽��j��xx=�	R>�.?����8����9Cm>��6?:�>�'�>����x����<Z	�>8/?�(�>�<��M4r��8�n��>\��?��d[ =�T)>`W�=γz�9�����=�>���ْ=��f��t6���<y��=@��=3�u�� ��'�B:�=U;�<�?��,?���=�%R>��%����P� �yw=��R>�s�=�t&>�佾#%���-����a�Y>�Џ?jh�?���=V�D=�g�=$�'�?%\�*��6!ܾ4����`�>���>�3O?\�?'�M?�AE?b>K���L��I���m2ľR� ?k!,?O��>w��r�ʾ���3���?[?�<a�*��O;)���¾��Խ��>�[/�i/~����QD�@�����8���&��?ֿ�?�A�>�6�/x�̿���[��}�C?�!�>�X�>l�>��)�:�g�Y%�q0;>��>�R?W�>��O?��z?��Z?/R>�8�0���t���t�<��#>�U@?-��?4��?��x?���>�!>�+���(���Κ#��K���GJ=2
[>���>B��>z��>�T�=�aƽ2"����<�p�=jc>Tw�>Td�>Q�>dx>.U�<��I?�C ?��"�5 `���Q>�g���y?fo(?N�?�F>�;Q�t���Ų��@?���?ܥ�?��>U��<�O=��������yZ�>��>	�> ��>˦?>���8�>��?��ȽI�Q���X�>��M�?jza?`�>�Ŀ��d���� gC��ƥ=G�Q�긱��d	>Sg�X�=�
����R������
���2���R���ɾ|���f��{�	?�>F6Y>�h�=�y�<���<|�= �>b��<�U=u�X�r��:��8�3eܽ�r���=�h�=M���Aiþn+w?�NC?�?FV:?�S>g',>���'h�>��ۼ=�?��k>E,˼ք���B�e��������ݾ@���ll�ꏡ���>r��;>�o8>�&�=m�\=���=��H= �p=Mƻ;|ml=���=��=W��=;��=�1>ߟ(>�Ho?.�;�����L�`�Q����?��m���>�.�;o$�>��<�ϑ��7���Z��?i��?�G�?;K�>:
��X>�>��;��3V����������1>ڲ�>�V��R��>�v?�+k�6���vw���?S@�I?ࣈ������a�>
9>t>�vQ��1��%]���f���V��a!?��9��,Ⱦ2��>%��=f۾A1ž��(=bz5>��P=�	���\����=_���n�8=�<n=�`�>*�C>^��=O֠�QǺ=	#A=dk�=_�P>ӧe9/F,��)�2C6=�W�=��f>�.+>���>��?�`0?�Vd?�5�>Zn�Ͼ@��iH�>��=�E�>-څ=koB>吸>*�7?%�D?`�K?|��>н�=h�>9�>ۚ,�˴m��l徲ʧ��<���?Ά?6Ը>�R<��A�ܠ�.g>��(Ž�v?~R1?3k?�>G�Q�ڿo�$���A�K=��:�귇=��t��={8�����P ��F��>`9?S%�>��>�N>&%�>��?x;�>`��=�s����=�K=�6=�y�jPh=0�(�Gǎ�O��;����.��G<0�8��m�����_�ֻ	ZF<���=���>�:>o��>���=��B/>���L�޾�=aG��,B��4d��I~�V/��V6�ҷB>�<X>	}��24��u�?(�Y>�m?>G��?�@u??�>U!�P�վ]Q���Be�US��ϸ=)�>+�<�<{;�h[`���M�v|Ҿ��> �>}��>��l>T
,�8&?�L�w=��.i5���>�b����&#�8q�^=�������i��d�+�D?�C��_�=�%~?��I?Jӏ?z|�>$���Őؾf30>k*��}�=�	��q�a��k�?n'?-m�>�;���D��3̾�r�����>S�H��P�������0�o_�e����a�>����о� 3��h��1 ��ԋB��Rr����>�O?.�?��a��[���UO�V��P����O?Xig?Z��>�7?�8?_���ў����y��=��n?T��?�:�?��
>L$�=f�I�>�G	?ʖ?5��?*\s?K>���>���;E!>�/��"��=f>
�= _�=jN?��
?�?W1����	������7�]�E��<�ߢ=GΒ>ш�>��r>���=�Bg=w�=Wp[>��>'��>7bd>��>��>X�ľ���0#?��*>B��>±V?qm�>P��=36�=���= �콳�c�5�8�+0�3�J��>v������[;i�)�6�?��ſ�?;I>a�=�@�&?ܖ��qP�*�>%��="�/�/��>�09>}�b>D�>7�>�b�=��>�i�=�FӾM>����d!��,C�B�R�\�Ѿ�}z>����W	&�ǟ��v���AI�pn��sg�~j�J.��Y<=��ǽ<#H�?]�����k���)�n���I�?�[�>�6?�ڌ�N����>���>�Ǎ>�J��[���Qȍ��gᾝ�?9��?N�>��[>�RN?�y?p¾�4s�@/z�6���e|��Ι��ꊿ�n������4��{h���I?4d�?�4>?�����\>:�?x!��I%����>|n�	Æ�˼E���>�~��2(��g��|0�,#��U?Y��?�@�?N��>���b��=�>�T�1?��M?>��?}b�>�X?sp�>�9? H�>e�?�	??-]T?.�W?2��>Vl,��Y����>e��>?UĽ�K}�*Ư�'�;�pO=Wl_=��=d��VL=�t�=N� �p'ý�-���Լ�U%�|�<r=�<$k�=���=KΦ>�]?��> i�>��7?���}~8��֮�a/?`�9=q����.��x颾�5>��j?��?}`Z?�Sd>�A���B��)>�Z�>h&>��[>�m�>3*ｷ�E�o�=�>�>h�=�SM�!ǁ���	�ߦ��@e�<�I>���>�9|>�,��̤'>�}��"z���d>�Q�<̺�|�S�
�G��1���v��S�>�K?��?���=�Y���	Hf�y.)?3[<??OM?��?���=�۾��9���J�'E���>\�<*��~����$����:�[(�:6�s>3�����e�_>��
���ܾ��m�.J����G�D=�����O=�#�i�Ծ%}�z��=�$>�t��D� ��&�������J?k�v=�i��z�T�	O����>�ʘ>���>�_>�[Ut�BF@�ά�d�=*��>��9>1���P�-G���`�>�F?[�^?�҂?r˃�y�s���D�zV ����Nѩ���?CG�>A8?�$@>���=���A$��zg���I����>���>=o��F�E����-�!�/��>�i?�>Ux?��S?ȉ
?��`?]%*?�w?��>aȥ����@&?���? �=H�Խ��T��9�|F���>�x)?I�B�s×>Έ?͹?�&?)|Q?h�?9�>�� ��M@����>�H�>\�W�)]��7`>��J?N��>�>Y?Ճ?�>>��5�Q̢�`���
e�=�%>��2?�8#?V�?���>��>����`�=Ub�>_�d?_��?L�o?��>��?y�*>w��>A�=ˈ�>���>A"?��I?�p?��I?���>�<�W���
��_[c��k��I:; a:r�c=�3/��5���J����<ɧ�;c���7�r����=8��g��/�<�_�>��s>L
���0>m�ľ2P����@>�}���O��*ڊ���:��=���>��?몕>cY#�巒=[��>�I�>���6(?��?�?X�!;��b���ھ_�K�)�>h	B?��=��l�s���1�u�j�g=C�m?'�^?N�W�W&����b?R�]?�f�q=���þ�b���龻�O?��
?��G���>��~?p�q?1��>$�e�b:n�H���Eb�}�j��ζ=�q�>W��d�}A�>қ7?XM�>^�b>�&�=Jv۾�w�o��4?}�?��?���?�-*>��n�(4࿬��wC���y?V�>)
ݾK�0?W4=����8����}����1��F9���G���ʾ�P�@��4n`�˄�=��/?��?Zr?C02?�##�����Aox��+����v��7/����.�mMQ�l�I��~|��RѾ����0�.��e>���m�A��p�?6�'?A$/��z�>묙�f��<;�%A>�����d���=��9;=�MS=m1i��1������: ?:J�>�*�>��<?b\�&*>�eU1���7��I���2>�ա>�9�>���>X����-�*��E4ɾ�م���ֽ�ƀ>�qe?1�J?��^?��O47��鄿�%�M~���ƚ�ym>N>d��>�v=���2�D�&�J�>�9|�1�!�y����
�R��=��&?N��>/+�>�:�?��?T)����:gj�QF�T�=_T�>��f?���>hu�>��ռ��q��>6p?z�>S��>oD���l-�l/b��`g�#gg>[}�>�>�2>�� ���a�i���7l��4�I�ᆪ=��W? �w���R�#��>Y}8?�7�3>��%(�=���='��x����U�:��6>D�>�C>��<>����#2+�AT����1B)?B(?�ϒ�vt*��~>+�!?1`�>�7�>g%�?�g�>��¾�h�a�?)�^?c?J?91A?��>�p=�{��[�ǽ��&��,=�Ç>�([> l=���=��N�\���sC=*��=�,ͼ��J�<�y���H<sr�<�4>��Y�P����ѽ �K�վ]	��˘� =޽u·�$���Ю��W����S�)��el�GTa��q�{��Yr��X��?��?nj9�\�D�Gߛ��b}�h���>�g���8��ׅ���gҽtk���Lپ�F��O�%���F��Fx���r�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@e{A?9�(�4�쾕ZV=���>A�	?��?>�81��C�:����X�>9<�?E��?��M=��W���	��{e?U <�F�!ݻ��=�)�=�1=-��ڄJ>�D�>E��^A��oܽE�4>i܅>(A"�`��:|^����<��]>m�ս@��ք?���\4���4R��1���-�> $?�� >7}ϼ��6?�/���ݿ_J~�Z-s?�@G=�?v�3?�ϱ��ʞ>������-?5b?cd�>RjC�S|���k>ə�將�Q�%�c��dF=[Q�>;��ԩ�&(���U8����u;�e���ƿ�D��^�R«=����I�����婽g�������T��+�����=5�=4I7>óf>DU>�$>%J?�[k?�U�>/9B>7$�j���<ܾ�~��m���V��N�j�%YֽIo���ھ1����r�p&�CE�4 =���=�5R������ ���b�ϖF���.?�o$>��ʾg�M��~-<�oʾ��������륽G0̾K�1��!n��̟?��A?������V�}��pZ�����&�W?L�T��t款���=�����=%�>C��=���S"3��S��g0?";?LN�����Pr*>X+���=��+?�?N�^<x6�>�Z%?T`*��b��d[>gZ3>d��>j��>�9	>���%�۽}y?�|T?��O휾4ǐ>%B��lsz�0b=�>�a5�H��e�[>Դ�<���X����6D�<�'W?䗍>�)����Z��&���t==�x?��?�+�>C{k?��B?a$�<c���S���<dw=�W?^)i?��>����r	оԀ��M�5?ݠe?(�N>�ch�[�龀�.��U�|$?��n?^?�{��t}�������o6?��v?�r^�zs�����y�V��=�>�[�>���>��9��k�>�>?#��G������jY4�)Þ?��@���?��;<��s��=�;?F\�> �O��>ƾ�z������:�q=�"�>ڌ��{ev�����Q,�q�8?ڠ�?~��> ������#�=����i��?���?e���i8]<B����k�� ���d<bF�=ݧ�*_&�!h��8���ƾ��
���5[���Y�>7}@��뽡��>o�8��h�`jϿbT��QwѾ�t��?���>�8ҽ*����j���s��E�n
G��&���s�>VV>e������۵{��:��Yü_��>�~�*��>��X�������%�;��>�<�>�q�>�8��#佾���?8���g^ο�����X�Y?5�?-9�?w?��g<��r�r�~�_�I�HmG?�1t?�zZ?��!��\_�m�/��j?�'��R`�e4�mCE�:�T>U"3?���>��-���|=ɮ>Ja�>/]>35/�W�Ŀ!Ҷ�����f��?��?0e꾅��>���?�o+?#��S4���x����*��ٹMLA?<2>�[��,�!�b=�����S�
?fB0?����9���_?U�a�]�p���-�M�ƽr�>��0��g\�|L�����`Ue����RKy����?�^�?��?/��A�"��6%?��>~���Q9Ǿ�F�<5��>�$�>�'N>o_��u>C���:�\	>l��?7~�?Tj?���h���GO>��}?
��>���?�v�=w��>̞�=K[��-7��M#>���=�8+�me?��M?��>,a�=�17�ɜ.��5F��R����X0C����>�/a?�_L?A9c>pN���g3�� ���ʽ�m1��⼣�@�T�+��5߽��4>vb=>�>�|C�P�о��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?m��uM��li~����6���=��7?6񾮷y>��>UC�=�v��̪�H�s���>	V�?Z��?Ɇ�>֢l?50o��2C�K,=�R�>��k?^[?^&����� C>��?���X���-��9f?��
@�q@�o^?�ߢ�A�׿�2����W���c>>%Z�<H�>;�j�(=f)�����Oig<E?2>
�>�hK>�@8>>z΂>H�`>"n���@�7J�����[E��<���*����Z� �����p��C��U�ʾ�޼) ƽ�b����U���:�g[h�_)>�NG?��M?=?���>.�T����=6�ླ|1=��H=]FK>���>r?;f7?�s?�J=����˳f�z���Ő���R�����>�*c>S�>���>
��>�s$>���>��>�St>K�w>�r/=��A��8�=@7c>���>���>�p�>�C<>��>Fϴ��1��k�h��
w�n̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?'���z)��+���>}�0?�cW?�> ��x�T�4:>9����j�5`>�+ �}l���)��%Q>wl?I�f>�u>�3�e8�)�P�@}��i|>>36?鶾v@9���u��H��bݾnGM>ľ>�D�l�y����5vi���{=x:?��?�5��ⰾz�u��A��SR>p;\>�]=&k�=KWM>�bc�X�ƽ�H�hc.=2��=ƭ^>��?/-*>�ʕ=�%�>�헾hR�
L�>�1D>��0>w@?��%?���}���.����+�>�s>���>��{>�A>�I��M�=��>ad>K�������u��=�Y>�!��4f]��${�p[s=�藽���=�|�=d���;� �6=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?��>w��?�X?���>m>T���K��b͆��e��H>GC�>���=��vVF��ǒ�S���V����A[�f�0ډ;���>$�<ߤؾMpc>�F���ξpj���̴>|�=,�>��>���>K�>#i�><��=��<����ܚ�q�K?�? ��Z+n��6�<B#�=��^�j?584?��Y�;�Ͼ�ר>*�\?���?��Z?7R�>��>��4뿿�}��v�<O�K>�&�>�I�>��n�K>��Ծ8�C�|�>�ė>�����(ھ����m���U�>~i!?���>�=�� ?G�#?"�i>��>D�E�<���E��?�>���>E�?�~?r?E����}3�����᡿��[�|�L>��x?J?֋�>���!N��܄h�N�M�1왽?7Yg?J'�P�?��?�??��A?�df>��g�ؾ���,�|>G�!?��R�A��&�T��N�?�(?�c�>7���ZԽ2�ϼ]&�����.<?��\?�}&?tY���`��¾Z��<*#&�L�x�pa<��9���>4I>*���M��=*>>J"�=��n���5� .o<Dμ=mi�>�K�=��7��揽��.?d>�Ҿ�=��X���:�C��>4�������A?�C���c�����^2���t��:�?���?	�?ڵc;��[��u)?�`�?�1?�!�>��Ծ�&����羇,v��v�2��!ݷ>�T?��� �/��Ǹ�Ȭ�P\����ד�%��>��>�?�n ?�`O>_M�>�.���'�LO񾎯��^�PR�lh8���.�����࠾ #�����¾
|���>����|��>Y�
?�ph>@8|>�R�>Suƻ�;�>��Q>�K>b�>�W>�4>Rp>�� <��Ͻ�JR?W�����'�Щ�y����.B?!qd?i8�>�h�ֈ�� ���?ǆ�?Dr�?g7v>^}h��)+��n?sC�>
���n
?�p:=��d�<0Q�����o8����Ť�>Ob׽� :�PM�H`f��h
?5,?-����̾W%׽������j=�R�?��(?:�)���Q��vo��W�8:S�
��N�i��b����$�npp���GK������R(�K(==k*?�<�?d�a��Q_��d-k�"4?���e>�1�>�y�>;�>$KH>F1
�T�1��]���&�|��	R�>upz?7^�>�1I?<?�P?�L?#ɍ>4%�>Ҡ����>s!<8ʡ>�z�>H`9?*�-?~�/?�?��*?��`>L�������ؾ�?��?�(?��?�z?���X"��u����A[��oy�.���̀=j��<|�׽�cw�A�S=?0U>�?��$�S�0��ݾ,z�>
[)?��>���>@��!ň�[̶<�W�>W!?��>���`l���2X�>�H�?d���ʀ�<�Q+>U��=����T��i��=o�o�E�=��1< ����q:�fה=���=�<.�Z���hЈ<6\=+�?�D*?<4>���>���`w���羣���S�o=p?>�\=���P���_잿��s��zR>���?� �?ؖ>T��=�D�=tB*��x���y���ξ7-����
?h�%??�\?ナ?�I?�/?7�+>�� ��0��7���C�����?A",?�ϑ>��:�ʾި�T�3�̦?��?aa����T)��¾�սm�>qr/��~��쯿*�C��xg��������}��?Q��?�C��6��v���������C?�	�>���>Rd�>Ѣ)�f�g��s�c�9>L;�>��Q?���>9�P?B�w?8zL?H>�=�G׬�ᖿ�9��*>��C?�Py?:
�?�#q?���>(��=G�E�����c���S��]�`lp��
/=/y>"��>���>f�>[�>Õ���a��s�ؽ�=oQ|>�"�>f}�>U�>lȚ>w��<��G?N��>fq���������d����)=���u?��?�+?�v=���l�E��D��O`�>r�?���?�2*?��S����= �ּhٶ���q�z�>�˹>�7�>�˓=�kF=�z>Z�>��>���[�dk8���M���?�F?m��=��ҿY�U���<��,0=����R��⣽���Q�Ҿ�zؽ�1�:�S��8���ؾ��$�̾O��{? �t=�1�:)lP��-u�|^>䨀>$��>A�>UM�=�cƽ`�J�-�>���'�ǿS�l߄<�����>��=�2���Q?�G?#6?��,?���=���=C�<��>a�e>�A?��>{�-�����］�̓������>�a��$#K�+���¿�=b<�=�rF>�MF>9&^=��	=��0>��0��z�=�(���-�?��=y[�=���=+�<��>��>D�e?�������񣝿�
��ʌ?c�fʽ��¾���>���=�Ҕ�5̿�?�eR�?v#�?b��?X�?4w�=N��>��O�o]�R
��lX���|>�>�>���;�Ȉ>a�?���<�J����ƽ�h�?oS�?j�?�d��t���MZ�>��7>@,>�R�-�1�ɗ\�ʭb��{Z�^�!?C;�7̾�@�>�*�=�#߾��ƾ�.=�~6>�7b=6��Z\�rә=�&{�C�;='!l=Qډ>��C>���=;���*�=�I=��=��O>x斻��7�7�+���3=���=r�b>�&>���>��?b0?=Wd?�7�>�n�`Ͼ�:���R�>3�=J�>���=myB>Y��>��7?��D?^�K?�|�>%��=�>m�><�,���m� h�<ħ��S�<ј�?І?/͸>KfQ<o�A���Vc>�y+Ž|r?*Q1?�k?n�>$V�P�� W&��.��k���&:���*=7lr�dRU�����m������=�r�>���>��>/Ky>��9>�N>Y�>w�>���<.��=gD����<L_��7��=�Ƒ���<x<ż���ǉ&�T�+�+Ȧ�1��;�D�;�\<h7�;6��=���>!7>���>7��=��_F/>!����L�Ͼ�=�I���,B�4d�wJ~��/�	U6�R�B>)>X>v���3���?�Y>�p?>���?�?u?!�>��9�վ�P��De��NS�ظ=0�>�=��|;��[`���M��{Ҿr��>P�>F��>͋k>��,��@��zk=g��6�5�>���%E/����Tq��s���矿�tj��P���C?�<��*��=�,~?;JG?�~�?"�>Ҹ�3�Ͼ8T4>MFz��E=ۋ���q��߇��|?��#?���>�A���bH�9̾����R��>
I��P������0�5%������>;���о�3��a�� ���|B�6�r��#�>գO?O߮?p�_�.S��>LO�o��Q��
?^g?���>��?o�?�x��P	����M��=/�n?���?�G�?>m*�=2ո�V��>�	?l��?��?�?s?«9��;�>x�;��#>td�� ��=��>�o�=�t�=��?;
?D�
?�ș��	�Ob����U[����<�5�=F��>j�>�3l>`q�=}�y=���=]V[>�'�>(��>�!f>���>�;�>�5ܾ{N"�]�?�\�=v�y>�M?��>��>U;�=��d��&�S�Wk(�-'�a���ļ$��<<�-v�2�?lǿ��?i�>��&��E!?ܾԀ7���K>���=Zܲ��>vl>��k>6B�>~��>���=��e>�N�>:dӾVj>���~[!��$C�qR���Ѿblz>�����&����m���.I�#p��xg�Wj�=+��:=����<�D�?���2�k�,�)�������?�p�> 6?2Č��鈽d�>���>8��>#Q���������]�G�?���?�'a>5ا>>�B?H9�>���|j�ah{���v�V�?��ɓ����|����7����N����][?yȈ?��s?���<���>3�?���#�$�Kc�>w�澶@K�2?����>�J���0�����5�)��B���Ց>���?kب?c�?r��2�8>H[{����>��V?o|?3�U>N�A?b2?��H?�17>ת?T�>?�GZ?N�7?mȅ>�5:��?��� >!$�>S<�>�f����=|��=�=�=J7l=����i�����
��'����=;�=[{����<���=��"><�8>;�>Ԥ]?%L�>��>]�7?���^w8��Ʈ��*/?e�9=�������Hɢ����>�j? �?dZ?�ad>��A��
C�*>{Y�>rq&>\>�d�>�w�@�E���=�L>�Z>Jǥ=ReM��ρ���	�m���!��<�'>@t?�<�>D�$�{�=Oz���h��i>q ����ܾB1@��D���?��������>8CP?��*?*o >�ھg�T���`��8&?<�7?� [?pv�?��
;WF��FE?�&hT��N�?7f>��>�:̾77���⭿�F�x䉻���>��ɳ����\>!
�[�ܾ��k�T>I�:*��M=J��[=ڭ
�w�վҢz���=��>/���c!��*��6���dI?��v=�����S��ɹ�(>	�>u	�>��M�㜋��y@�����=O*�>�Q<>uJ���s���G�:�����>`�E?��^?y�?�Ň�]�s�t�B�k���?��������?���>��?��5>9��=᬴�Qq���e��lF�@C�>Ɯ�>�N�XmH�����I@𾺅$��߇>��?m!>�_?�gT?�/
?�^?^�(?1?_��>�Խ����E&?i��?8=�ֽj�U�s�8���E���>Ux)?Q�B��˗>�?�?��&?�DQ?�y?�>s�
�@��`�>~�>|�W�FD���(`>�J?aҳ>@jY?氃?��=>�F5����H��� ��=.V>��2?XS#?��?�V�>� �>�+�����=���>H^c?�?��n?_>Ɨ?�H9>���>�"�=;�>w��>L�?�SH?��l?�K?.�>N�<B�������In�$(N���<���<?��=郬��1&�7���%�<�p�:9��O����Ǽ�$A�	�¼˔4�jb�>jt>������0>��ľR����@>)闼T���n��|�9���= ؀>L�?�X�>��#�> �=_��>�>���-�'?֭?>?���;�ab��G۾n�K����>��A?�G�=��l�Ĉ����u��j=��m?^H^?@W�8�����^?�h?��Ǿ��D��9�i���zپ�Y,?�c?�z)����>��p?v Z?W{�>���p?i�4d��GD����ھL��=�*x>�o���a�]2�>J09?K��>ni�>���=����~Z�ȏd��Q&?���?@��?�J�?Q�|>�R��!ݿĉǾD왿a�k? G?���<^0?��?^@��)@�����j)8��ݾ����Rվ|���#o���������<�O<?�6?�?��G?��$���%�R�`�������<�(�
��L"���5o��� �>Q�haؾb�^�Ĉ�;�=k~��OA�Uo�?v(?
-,�G=�>+������M̾�(C>����������=�f���;=�+V=[�g�=.�7�����?��>�I�>�k<?3q[��=��U1���8����d�3>��>D͒>��>��G;n,�f�潒LȾ�˃��SνΧv>��c?�`K?�An?��k(1��`���}!���-�OG��K
C>�>���>q
W����B6&�:t>��@s��^�ck����	��|=�w2?�;�>�ۜ>1D�?�B?�j	�A����w��=1���<2��>�i?�J�>�K�>��ν�� �\��>�@t?X��>R�>�����B�k�e���H��$8>z��>8�>�s�=��M��g^�����Z2K��0>W�C?��~�v_�O��>��A?�J���������>�<��ڛ�>�*;�q>���>)W�=rDO>��ؾ#F�����k��m )?��?+����*�[�}>'B!?���>0�>pC�?�Ϝ>�\¾b��:��?��^?��I?t�@?��>�=ُ��ɽ�W(�;�*=��>~<\>9k=/��=���tZ�|]���A=�[�=�߼V����l<�ش�l8<���<��3>�iۿC@K���پ����"O
�%��k������'����9��1
x��D��(��U�
?c�����Om��j�?��?Fړ�r������`���w��ّ�>~q�����/�� 4�6����ྃ���SN!���O�Bi�d�e�O�'?�����ǿ񰡿�:ܾ.! ?�A ?8�y?��0�"���8�/� >D�<�,����뾫����οK�����^?���>��t/��u��>㥂>��X>�Hq>����螾x1�<��?8�-?��>Ǝr�-�ɿ^���bä<���?0�@;vA?��(�����iU=g��>�o	?��?>R�0��*��ΰ�,y�>�8�?Z��?֜M=O�W��}
�{ee?���;<�F�p����=���=�{=.}��BJ>�8�>�/�2?A��ܽ��4>��>�!����Qi^��<��]>dԽ�g��_��?O+>���k��a@�c�x�(j>�C?��>�$�:DY8?��*���ҿ�o�D�c?d�@s�?�z0?�1ɾf|�>#ϾH�=?��#?,5�>I��bp��n�=���<@ߑ=ҠӾ�tS���=��>&�=&GR��	�wk �[=�c�<�1�A&ÿO'�Ş��Q=o�?�B��
;۽�T���żnZ��(�p��ӽ�m�=���=�J>Q{>`P>H�7>�U?��i?}]�>�">�7ν��h���žP@���T��77�מ����5�"G��)���޾����H�H=���߾�"=����=U2R�A����� ���b���F���.?��$>��ʾm�M��=-<�gʾ�����F��0楽_1̾o�1�'n�qʟ?T�A?���V�}����La��:�W?Q���O����=���ʣ=�$�>uy�=���"3��S�gw-?�?�)�����Q�>'e%��R=^5?.5?y=9<�>`�*?��������;>)>%�>���>��=g����0�Z�?��X?�.�Z����j>:T����>�:7�=Qd�=)�F������UM>��=*���-a廼!��=Y(W?Ǜ�>��)����a��V��\==߲x?��?	.�>X{k? �B?��<;g��K�S����cw=��W?r)i?v�>�����о<����5?�e?f�N>�ah���龮�.�VU�$?I�n?�^?[{���v}������'o6?��v?�r^�{s�����*�V�i=�>�[�>���>��9��k�>�>?�#��G�����vY4�#Þ?��@���?-�;<' �?��=�;?{\�>׫O� ?ƾ){��������q=�"�>���lev����3R,�B�8?͠�?x��>��������3�=�C��U6�?FW�?�����SQ<�T��>k����H��;�`�=i�:���4��[��8�� Ⱦ�]
�;-���@��)�>ƃ@�b彞x�>P4��L⿝�пi���Iվ��z�E9?�Χ>5Fݽ�ʥ��Di�ڟr��lC�l�D�T��0d�>f>���s)����{��J;�3V�����>җ	�v�>��T��p���矾Q�*<��>[�>%@�>a�����?�����Bο#���,[���X?�c�?�@�?lO?6I<�v���{�~Z��BG?'�s?_>Z?�}%�a�]��-8� �j?Z_��xU`��4�aHE�nU>�"3?�B�>S�-�P�|=�>S��>�f>�#/�w�Ŀ�ٶ�7���X��?։�?�o����>x��?xs+?�i�8��m[����*��",��<A?�2>���*�!�$0=�LҒ���
?~0?�{�V.�[�_?-�a�c�p�/�-�w�ƽ�ܡ>#�0�`h\��e�����We�2��Dy����?}^�?��?ݳ�� #��6%?��>q����8ǾY�<��>�(�>�(N>_A_�۳u>����:�wg	>1��?b~�?Mj?㕏�����}U>��}?ͻ>���?	>�>3:8=� ���<�Po>'i>f���?8R?I��>���=͕L���*�`p7�3J�Щ
���;��6`>d�Z?R�R??�>?�޽cM�����ύ���#�{?A�%�)����i�ٽE�0>\b:>�5>�BԽ������?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�e��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=7M�>Μk?�s?�Qo���i�B>��?"������L��f?�
@u@a�^?*�ӿ����������h>dd�=��|=<�3��'?=�4^=�E��d�F�B >���>nw@>��@>zM<>���>-��>I��'�Pˣ�q+���K�W�9��a�������(>������l0��n���Tƽ����lĽB�<��=�4T?"�Q?F.o?�2 ?3���@>����"=4y �2�=8P�>�O2?s�J?-�(?�=r����d�#���e8���6��{C�>��L>�y�>���>|��>v|�GmF>�f?>a�~>'�>�y/=��ٺ#h=J�N>�Z�>�J�>��>�I<>r�>Eʹ��1��e�h�	w��̽��?}��x�J�r/��E5�������t�=_.?�s>���@пl����/H?=����)�o�+���>e�0?�cW?ů>/��j�T�b>>��� �j��j>�$ �Jvl��)�F-Q>ki?5�g>�0v>�3�o�8�MEQ�����S>}>�?6?7����7�K�t���G��ܾ�M>;ٽ>�S��B��������i���u=]:?T�?�]��H����t�.��R�Q>�[>D-=�Ʈ=f-O>)Pd�3�ƽ�HG�a)8={�=�,b>�[?�4>>��=�>^N�����V�>"�>dam>��;?��%?V<=S7��iW���6�o�D>r�>}sf>�2�=��P�^�<���>���>1I�=�}���A���O��@�>lPڼ��q���޽���˕��9�>��=�f��@c���=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾNh�>|x��Z�������u���#=T��>�8H?�V����O�i>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>:��?�gY?ooi>�g۾<`Z����>ѻ@?�R?�>�9�~�'���?�޶?֯�?&�>_Q�?�xl?��>�᥾b�D�kѨ�#?��|o=:��=��>E�=����,�\�M���w�������FK�I�=v8�=�ݵ>�!������#���&=�j��G��e�?�&3>��V>���>o� ?��>o�>�5�=+�2���۾�C��$F?�K�?��<�r��S��-?93���n�?�3(?��=�?���>��S?*n?t&?=�)>���GU��q|Ͽ�<����۽��P>�M�>E �>������l>�҄�*�;�q�>=/�>J >�U�P�Q�V�:>��>��;?k�?S��>K� ? �#?��k>�ϱ>u
F�g��ӻE��>�>���>�k?Ub~?m;?�湾�4�����1᡿�u\�n I>k�w?�?�>ξ��xt�����1�B� g��n�?�hh?
pὫ�?셉?W�>?״@?�he>����Nؾ�
��P�}>S\$?�y����E�(�7������?m�>���>�A��	��/1=�,������?��t?�!;?��羟`b��ۢ�3�=}���K7����K=��>+��= ��\>rF>�0�=jꁾ�}=���;i��=�5p>�M�=hH*�`ʽ(\1?L�>���Ż��@��V*����=�_�=䗶��$@?um��;t�*���}x��<��<چ?���?���?~�
��?[��s"?ކ�?�%?���>0��$��zDȾ��5�U9��0�)�KO>�7?�)꽀�8��¹��ެ���Y��Hl�:���=�>��>r�?Z: ?�Q>Yβ>=-���&����n��*^���kh8���.�.��p��f�#�^g��^����{�u��>gh��nm�>;�
?� i>��|>��>�a��s��>��R>�~>���>��V>@�4>s�>Z�0<��ʽoKR?����E�'�ĵ����d1B?qd?�3�>��h������n�?~��?�r�?:v>"~h�w++�n?W=�>B���o
?�Q:=7���z�<@T��)���2��S��4��>	J׽� :��M�-lf�Dj
?/?���w�̾�4׽�$��j�=���?q#(?�g+�4=T�|~m���V�>\T�*��cEe�����K$��jq� Ǐ��������,�(��=�K)?��?"e���7�$���g�h��u>�c�e>���>���>\��>�X>���S�1�*�[�I�$���&E�>�ow?S�>��B?�9?vkH?��B?�h>�\�>,愾�^?�"=��>���>�9?%�*?��#?�
?��%?��\>�j�`2������j?�"?�"?ޢ�>�A�>������꼮��<m`9�����\	��;u=?I^=�0��P#��	1=�bD>�F?|���7��g��7n>	7?q�>��>P���怾���<x[�>3�?�L�>`P��+�q�����>�?�M�n�=��(>��= �{�.T;%-�=t���#a�=�D���7��<�
�=��=�SY���:8b;�X�;��<�?�V+?�U>��`>�O1���Q���F<:>8->n�=��`/��-���cs�Z\>>숋?��?$�H=���=	�=֗'��G��-������G=�U�>�?s�K?2�?u;%?a8?�M>i���栿��������?�,?袑><����ʾ����ъ3�Q�?md?� a�{�)��P¾	EԽ�>�X/��#~������D��0������ՙ���?i��?_N@�A�6��_辷���$@����C?s�>�w�>�&�>J�)�?�g�F�Go;>���>!)R?�>N3?�?��b?�G�>_Q3��5��I��4�t<�2/>:;?��~?�m�?��k?���>���=�ȿ��ʶ��ޫ��޼�ȍ���<p�=/�k>8��>j��>m�=��B��V-�3�\�ڝ>���>�-�>0��>��>=��>y>T�L?�?v$�c�,�V�������>d���e2?�U`?
k??(?>;;��Vp���޾�?=t�?���?��?p;B��y�=�|�o�Ͼg�#�T��>!�>�iQ>;�C>1�s>R��0>��?*/�=�Y�S���!a��# ?ql?��������<J�Q:=�f0�/��=Gҗ�+��z �=�&j��t�Wי��vཟ%	�ƿI����������}־����c?&#�=�!p>�>v���>k�>�<>��=�$�������y=������4�߅̽\���f���=��=�z��^1?��??�5??F?��L=�^=� >���>v��;��?�f�>R}=�[о:�]��s��|��EH�ž�(��w�jvV>y�=F�>�)G>s��+�۽]K��nB���S�=�dB=s��=>�=,�l=5I�=oL>8�U>�N>�k?"汾�ښ�Cɏ���	�-�b?%(F>y����J����>=�n>����}]ȿ.i�2��?@l��?Ù�>��ͽq�>�z��235�so��X�	��>�0J>p�
���K>d?��\= ���������?��?�3?V����譿8�>Df8>�>�AR�3�1�B�^�ec� 0Y�b�!?��:�\�˾Ά>��=J޾�ž��*=^L5>��^=�a�ͣ\�[��=O�~��b==qxp=Q�>{BC>㍺=&R��i2�= �H=f�=RwP>�G��q7���+�Z�4=���=M{d>��'>Ւ�>��?�c0?-Yd?<�>n��$ϾO<��XI�>T�=F�> �=0�B>��>6�7?	�D?8�K?!��>��=��>��>�,�߭m��m徥ȧ��<8��?ʆ?���>q4P<W�A���[X>�cŽ�s?vM1?0k?u�>�'��̿@;L�������V��������tC��i#>�����ֽg@>��?�>t[>�v>���>�&�>��>9�>>?��=�;�=W�[=�;P����zC�<�ED��0>D�k>h��<��a���r���Yѐ<�K)�3���p�C��=2��>+<>Ȭ�>���=����C/>踖��L����=�G��d,B��4d��I~�W/��V6���B>k;X>�}��;4����?��Y>*m?>���?0Au?6�>� ���վ�Q���Ce�AVS��˸=c�>��<�{;�[`�~�M�G|Ҿ8��>��>��>7�l>T,��<?�&�w=�⾘p5�p�>�i��_��?�.@q��<�������&i��j�V�D?�8��_��=�)~?�I?���?hx�>�<���fؾ1�0>���T�=����q�⓽��?'?TK�>�v쾔�D��>̾�Q��@��>qI�OP�����M�0����෾q�>�����о%3��f��������B�LLr�4�><�O?��?[�a��T���SO����Hx��WZ?�tg?��>�<?>?�:�����}���z�=f�n?Y��?�=�?�>��=խ����>�7	?�C�?n��?WWs?�J9��S�>�;��>#K��:��=�
>�u�=���=��
?�7
?��
?�K��d�	������S�^�;C=(ީ=31�>o�>'{q>2D�=��]=m�=�Z>�*�>D�>�_d>9H�>��>�Ჾ����� ??�>��>!�>?ê>6�=Q��W��n��RK-�[���
����d������k=��;g<�>�ƿ��?Ks>���G?�g��Ƶ�`3F>g44>�7�A0�>]�>�U>�s�>#Ţ>�N>߶w>դ>�XԾ�>�p�� �*�B��.Q�Nо>
{>�ޛ�A(����ڏ��G��˵��q��i�����-=�g�<���?
���>k��?)�����	?�,�>Nw6?q���T·���>2+�>�[�>4���X��tb����N�?���?��>�ک>��U?��?Bk���N�e]�I#r���o�N����J������\��H���)�
�]?��?@R?�%7=J�>Bܰ?8�s�G@3�`�
?S�߾��t�AV��;B�>�E~�<E�SuоF���8����>���?q��?���>N���%e>+���$?��S?Se?z��>�,�>�v�>h9D?,%F>>�>�O?.pW?(�A?��>VkP��,;0�s>�Q�>���.\�z�"����{��:/p>�Pr>Q�>Y�=��=�>q��Q�<zG���^���e�<�<�����F�<bwQ=�ɦ>��]?UL�> ��>��7?P��w|8��Į��/?��:=�u�� ��m������h'>��j?���?�KZ?Mvd>�A�UC��>
[�>?E&>�[><�>���VzE��=�>�(>���=kGL�����w�	�Co�����<eM>���>y8|>H(����'>�z���&z��d>��Q��̺���S���G���1�E�v��T�>�K?�?ķ�=&Z龔2��Hf�}.)?�[<?-PM?��?O�=��۾��9��J��J�)�>9�<9��m¢�0&����:�}�:1�s>4��͢��I�b>۟��D޾K�n��J���羀KJ=T���X=���<�վ�����=�	>����6!�����Ϫ��
J?��i=e+��X-U�F����>7֘>奮>�9�v2v�Il@�o���{�=���>";>�l����G��P��M�>��F?�
O?A'f?�a��A�u���,�-�
�2���&Y=Ru"?�;�>�n?�)#>���<h�ľ��!�����FW���>���>Է�	zU�'m��B¾�����>s[	?��>-�?%C\?�
?�
Z?��!?�?ޤ�>.���1�þ&?�e�?⃆=��ݽGX�dF9��tD���>��'?�:���>Q?��?R�%?w�O?��?��>���A��b�>�ԉ>W�dT���c>6�I?�=�>[?�p�?�?>�3�SF���D��H��=cz >�r3?qO#?�?���>���>4z�����=��>�sd?�.�?Y�n?��=�k?n�6>F>�>�+�=?�>1��>J?��L?I�q?�XJ?��>i�<vY���8ý�-~�	7W���`;z��<ث�={OԼ9�^���ɼ��<"5<���:������qOQ�%�����';!N�>�s>2���h1>6�ľ�v���HA>誟�4㛾%����I:�^�=���>V?���>�#��=8��>��>���6(?*�??�8;�b��۾�K��C�>�B?e�=��l������u�w�g=a�m?&r^?ȂW�2!��ԟb?��]?i��=�[[ľ�Od�����O?wZ
?#fE�4۴>(�~?ީq?�B�>Q(f�% n�&����b���m�?�=_��>�@�g;e����>r7?��>l�f>5��=��ھ��v����cx?��?��?*��?�o+>�m�~�߿�������@�?/4?y��ކN?�	G>��������(ʾ�S"������^���ž^z �1����	ɾ�-I�P��.Q?�s,?�Uh?��\?��������G�H�z�䌍�F)�0r6�dC�Ԏ/�[�=��d��ݾ`���S3��*��>�x�B�[k�?��'?�I3�m.�>�W������ʾ7�A>Š��r���i�=�_��h_3=��L=��i���0�N����!?1��>A�>��<?#]]��=�W1�T18�����->�ʟ>�ړ>/��>N�
:!`.�A
�fMʾ�愾��Ͻ��x>sOc?P�I?�>l?����G2��+����"�j�V�KΡ�BnI>�V>ֵ�>[D[�8"�$�&�x�?��Lt�y����/t	��J�=S�0?+�w>c?�>���?4?����-����u���.�	\�<җ�>�eg?o��>4��>�佈%"���>��o?*q�>���>jJ|�"�'���u�~�?��I>c��>�?z�l>�)'�R�b��(�������8�9��=�gD?����	∾ ��>��G?˭R�d@s�p��>64-���&�?�i��>��V
�=�?@�U>S�>�߾�K<�}I���OȾ�8)?�??���ߏ*��}>�!?��>�}�>>�?�=�>��¾U�9��?��^?
J?�A?���>�=-R��*ɽ.'�EW.=(ׇ>�[>(Tn=��=�(�V�[�����>A=�=�uͼ������<�B��i�K<���<xz4>�nۿ^MK���پ ������ 
�@����W��O�������x��u2���x����X)��`V���c��Ќ�n�l�s�?�$�?꓾��Y���xz��3c��;�>��p�u*~���Ι�R�����D㬾nT!���O�&i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾u1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�|A?]�(���쾫V=���>]�	?��?>�Q1��H�G���kV�>J<�?���?�{M=��W���	�M~e?�D<�F��)޻��=<�=�E=��єJ>ZU�>4}�{QA�q>ܽh�4>�څ>�j"������^���<��]>]�ս	7�����?�sZ�Z�f��0�>Y��:9>��S?4W�>�=��,?�F���Ͽr�]�'`?AP�?l��?��)?�ҿ�(��>�qܾ��L?.5?oB�>��%�C�r�ӫ�=@3¼��%��0��T����=&��>�C>|�0����v L��>e�]~�=5f�#�¿�{!�۽��*�=�83=�1�~އ�I��J�X�ͽ���}����q�=갌=ӈ#>�[>��*>�R>bX?>�i?HD�>��>��ٽ��h��y��b<H=P8R��D齀z��[�0�̾���p^���UR�zA��"�� =���=�6R�a���>� �^�b�$�F���.?�v$>��ʾU�M�Ǭ-<:pʾ=����݄��᥽.̾E�1�C"n�F͟?��A?�����V�"���V�	�����W?�O����9ꬾ���=,�����=�$�>���=6�⾞ 3�o~S�4x)?0D?�����H��9>�7��k|=ON0?�R�>v@5=��>\�0?��uD����>>TN>��>V��>�-�=p���{t�K�?XX?	yȽ�Y���>�؛� I��!:xnM=*�� ;3'�>�/�<%f�����~���{�=&W?���>��)�h��Z��]�<5==��x?
�?�)�>pzk?K�B?66�<�f���S���+cw=��W?�"i?ѥ>����T�Ͼl��/�5?L�e?��N>]Uh����G�.��U��&?r�n?ua?�̝�Ay}��������m6?U�v?'l^��t�����y�V�%>�> U�>J��>��9��c�>��>?�#�H��L����V4��?y�@c��?1<<�2����=$:?�e�>�O��Lƾm�������<�q=e�>/����Yv����`,��~8?���?1��>g���'���w�=S[��w��?�<�?	��>c<F�J�k�} ��ԃ<�}�=l���:#���8���Ǿ$�
��%��E��B=�>�J@/�����>��6��]⿘]Ͽ���"-Ҿ؍s��'?�]�>S9Ͻ�R��43j�
t�H3F��G�%��� ��>�_>n�Wƙ�{|y��:���{��>�+�b�>x�T��T��>া�W�<��>���>��>�ý޽��?L���~n̿�N��w��"�X?��?c��?�M?7=��W�*�|��?���oF?cZu?e	Y?G�C��N]�XѼ$�j?�_��xU`��4�oHE��U>�"3?�B�>T�-�A�|=�>���>g>�#/�w�Ŀ�ٶ�:���Y��?��?�o���>s��?ts+?�i�8���[����*���+��<A?�2>
���?�!�;0=�VҒ���
?G~0?D{�g.�c�_?�`��"q��@.�ǽZ�>w2�V�^��j �z��e��0���i{��ѭ?n�?kE�?���@#��$?���>�%��$/Ǿ,��<�>��>aRQ>TV� �s>f��,�9�e�>�*�?�-�?T�?A���צ���>*~?���>d�w?��	>�5�>d�=�־��u=��K>\��=|�}=)�?��S?�� ?�&>K�D�|�$�9�F�1~I��M�Di=��B>
�Q?1B?nOW>^�3j�;���s����:
�v0ܽ6/#��0���㼉q+>��!>I��=Qa������?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?oQo���i�B>��?"������L��f?�
@u@a�^?*��ݿxW��Γžk1��d
�=ڭ�=�80>v��fh�=���=��L�?-G�R!>N§>9�b>�!b>�F>�}[>|�a>yy���H��i��4p����7� ����/��9���ރ�i�"�C��\J��|S�=֞��8i��D(�B=��fn<CF>H�S?�=H?��V?�x�>�ؽe,>����!=m\˽�X>z��>�/4?�	D?Z�?�*x=3���jg�f��[������_��>$�4>���>\�>w�>�ҕ=�[>�?2>��r>�
>إ=0h�<�7$=��Z>�4�>�s�>?@�>�C<>ȑ>Fϴ��1��g�h��
w��̽)�?����L�J��1���9��ষ� i�=Qb.??|>���?пc����2H?!���x)��+���>��0?�cW?<�>%����T�a:>7����j�3`>�+ �ql���)��%Q>}l?j�f>�+u>��3�e8��P�y����i|>.6?y涾�9��u��H��Rݾy?M>[��>NtD��m�#�����{�i�uP{=Vs:?�?�*��,۰���u�J0���WR>�3\>M=�w�=~gM>2c���ƽ" H�Jq.=��=�^>JH?�/>�L�=�Ϟ>�痾ǝ\�ښ�>rM>��3>��??�4&?(Qq�;�b��hw��~-�F�m>���>y>L��=x�Q�C�=K��>��j>rѼhh������6��m^>^5��zk��!s�*v=l;���\�=�܋=�c����2��H=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?,�h>�R�?Zf?�	�>_��j=�-����N���N+���=ӣ�>�z>�ﱾM:A��׍��뇿�By�E/1�)W�=o.�<�V�>j���1����'=?�[��Z���O9��s�>49Q>�I>��>��?�v�>��>-h�=��`������J���MJ?��?�g��Gn�pK|<�nm=R�S���?[�0?�;4 ���>\?��|?JRU?~�>B�>���|��RQ��[� <G�A>��>M��>�����L>F����(5����>��>� R��;̾��|�����0/�>!?R�>W�=ؙ ?��#?��j>�(�>IaE��9��0�E�?��>���>�H?�~?��?dԹ�qZ3�����桿��[��9N>V�x?�U?Uʕ>M���񃝿�fE��@I�����h��?�tg?ES�,?@2�?��??]�A?�)f>'���ؾ6�����>��"?�:̽��F���.���,�?\,�>TJ�>�̽���)����%�p�wR?�h?v3?v���'ea��������<�毻�=�f�h��'�FH>�F>�������=sH;>HB>�)`��FG��ں���=ꎏ>=m�=� ,�*���~h.?|ͨ=��žԒ���X��5���->y�5>����S;?t,�"�p��>��V����K�"�?���?X�?z���V_���,?H1�?u�,?A�?W����n��#EҾR��}��j��K{�>��?���;�����Ч��b�����/����>���>�?|c ?<BO>�_�>
'���'��3�����^��]�=l8�9�.�2��}���~#����'¾��{��M�>9_����>3�
?wBh>��{>��>�hȻI=�>R7R>�~>fl�>g�W>�
5>��>�<2<ѽ�KR?���D�'���� ����2B?�qd?*2�>i�ɉ��#����?���?Os�?l<v>�~h��,+�Hn?�=�>����p
?\:=��G�<�U������3����ī�>�I׽� :��M��mf�!j
?]/?����̾�<׽=���zi=pe�?�&)?�*�A�Q�[o�W�W��<S������i��y��*�$���p�����^��T%��(�n�*=��*?4(�?���eGج��yk��:?�b�e>���>Ɣ�>nx�>uH>��	��1���]���&�U
��t��>xY{?�><�E?�:?piJ?�F?#��>Dz�>������>Q�<@ӥ>P��>�<?��0?�|*?'�?�!??�^>����x#��Lrھ�?��?Ok?�h�>��>]���򋽜t6�9hA�7�|�Nᙽ;��=+��<�o׽��j��xx=�	R>�.?����8����9Cm>��6?:�>�'�>����x����<Z	�>8/?�(�>�<��M4r��8�n��>\��?��d[ =�T)>`W�=γz�9�����=�>���ْ=��f��t6���<y��=@��=3�u�� ��'�B:�=U;�<�?��,?���=�%R>��%����P� �yw=��R>�s�=�t&>�佾#%���-����a�Y>�Џ?jh�?���=V�D=�g�=$�'�?%\�*��6!ܾ4����`�>���>�3O?\�?'�M?�AE?b>K���L��I���m2ľR� ?k!,?O��>w��r�ʾ���3���?[?�<a�*��O;)���¾��Խ��>�[/�i/~����QD�@�����8���&��?ֿ�?�A�>�6�/x�̿���[��}�C?�!�>�X�>l�>��)�:�g�Y%�q0;>��>�R?W�>��O?��z?��Z?/R>�8�0���t���t�<��#>�U@?-��?4��?��x?���>�!>�+���(���Κ#��K���GJ=2
[>���>B��>z��>�T�=�aƽ2"����<�p�=jc>Tw�>Td�>Q�>dx>.U�<��I?�C ?��"�5 `���Q>�g���y?fo(?N�?�F>�;Q�t���Ų��@?���?ܥ�?��>U��<�O=��������yZ�>��>	�> ��>˦?>���8�>��?��ȽI�Q���X�>��M�?jza?`�>�Ŀ��d���� gC��ƥ=G�Q�긱��d	>Sg�X�=�
����R������
���2���R���ɾ|���f��{�	?�>F6Y>�h�=�y�<���<|�= �>b��<�U=u�X�r��:��8�3eܽ�r���=�h�=M���Aiþn+w?�NC?�?FV:?�S>g',>���'h�>��ۼ=�?��k>E,˼ք���B�e��������ݾ@���ll�ꏡ���>r��;>�o8>�&�=m�\=���=��H= �p=Mƻ;|ml=���=��=W��=;��=�1>ߟ(>�Ho?.�;�����L�`�Q����?��m���>�.�;o$�>��<�ϑ��7���Z��?i��?�G�?;K�>:
��X>�>��;��3V����������1>ڲ�>�V��R��>�v?�+k�6���vw���?S@�I?ࣈ������a�>
9>t>�vQ��1��%]���f���V��a!?��9��,Ⱦ2��>%��=f۾A1ž��(=bz5>��P=�	���\����=_���n�8=�<n=�`�>*�C>^��=O֠�QǺ=	#A=dk�=_�P>ӧe9/F,��)�2C6=�W�=��f>�.+>���>��?�`0?�Vd?�5�>Zn�Ͼ@��iH�>��=�E�>-څ=koB>吸>*�7?%�D?`�K?|��>н�=h�>9�>ۚ,�˴m��l徲ʧ��<���?Ά?6Ը>�R<��A�ܠ�.g>��(Ž�v?~R1?3k?�>G�Q�ڿo�$���A�K=��:�귇=��t��={8�����P ��F��>`9?S%�>��>�N>&%�>��?x;�>`��=�s����=�K=�6=�y�jPh=0�(�Gǎ�O��;����.��G<0�8��m�����_�ֻ	ZF<���=���>�:>o��>���=��B/>���L�޾�=aG��,B��4d��I~�V/��V6�ҷB>�<X>	}��24��u�?(�Y>�m?>G��?�@u??�>U!�P�վ]Q���Be�US��ϸ=)�>+�<�<{;�h[`���M�v|Ҿ��> �>}��>��l>T
,�8&?�L�w=��.i5���>�b����&#�8q�^=�������i��d�+�D?�C��_�=�%~?��I?Jӏ?z|�>$���Őؾf30>k*��}�=�	��q�a��k�?n'?-m�>�;���D��3̾�r�����>S�H��P�������0�o_�e����a�>����о� 3��h��1 ��ԋB��Rr����>�O?.�?��a��[���UO�V��P����O?Xig?Z��>�7?�8?_���ў����y��=��n?T��?�:�?��
>L$�=f�I�>�G	?ʖ?5��?*\s?K>���>���;E!>�/��"��=f>
�= _�=jN?��
?�?W1����	������7�]�E��<�ߢ=GΒ>ш�>��r>���=�Bg=w�=Wp[>��>'��>7bd>��>��>X�ľ���0#?��*>B��>±V?qm�>P��=36�=���= �콳�c�5�8�+0�3�J��>v������[;i�)�6�?��ſ�?;I>a�=�@�&?ܖ��qP�*�>%��="�/�/��>�09>}�b>D�>7�>�b�=��>�i�=�FӾM>����d!��,C�B�R�\�Ѿ�}z>����W	&�ǟ��v���AI�pn��sg�~j�J.��Y<=��ǽ<#H�?]�����k���)�n���I�?�[�>�6?�ڌ�N����>���>�Ǎ>�J��[���Qȍ��gᾝ�?9��?N�>��[>�RN?�y?p¾�4s�@/z�6���e|��Ι��ꊿ�n������4��{h���I?4d�?�4>?�����\>:�?x!��I%����>|n�	Æ�˼E���>�~��2(��g��|0�,#��U?Y��?�@�?N��>���b��=�>�T�1?��M?>��?}b�>�X?sp�>�9? H�>e�?�	??-]T?.�W?2��>Vl,��Y����>e��>?UĽ�K}�*Ư�'�;�pO=Wl_=��=d��VL=�t�=N� �p'ý�-���Լ�U%�|�<r=�<$k�=���=KΦ>�]?��> i�>��7?���}~8��֮�a/?`�9=q����.��x颾�5>��j?��?}`Z?�Sd>�A���B��)>�Z�>h&>��[>�m�>3*ｷ�E�o�=�>�>h�=�SM�!ǁ���	�ߦ��@e�<�I>���>�9|>�,��̤'>�}��"z���d>�Q�<̺�|�S�
�G��1���v��S�>�K?��?���=�Y���	Hf�y.)?3[<??OM?��?���=�۾��9���J�'E���>\�<*��~����$����:�[(�:6�s>3��`ߠ��Yb>P��`u޾'�n�(J����iCM=4��KGV=����վ�4�J��=2'
>U���� �D��֪�0J?�j=Wu��pbU��q����>���>��>��:���v��@�&����1�=u��>�;>IV������}G��8�]>�>NQE?5W_?k�?�!��Ts�0�B������c���ȼC�?Zx�>h?�B>���=H�������d��G���>���>\��E�G��;���0��B�$���>M9?˩>��?S�R?j�
?s�`?�*?:E?�&�>3������gA&?��?L�=y�Խ=�T���8��F�j��>�)?��B�6��>G�?��?]�&?�Q?6�?��>D� ��C@�e��>X�>��W�b��Q�_>ݫJ?W��>�=Y?�ԃ?��=>��5�T袾�ݩ�N�=?>�2?Q5#?Y�?7��>H�>�`����>��o>�sn?W?rJ�?�_�=~��>�4�<�>��v>*��>GX�>e�?L5?A[}?��??�׌>Ԟ	����+�=Nn��,���VL���,	��(=�=@�U�#����9�mJ=�<��d��.]�7.��.`��ڏ=WL�>��s>-����0>��ľVL����@>>����N��b䊾؋:�%�=ŋ�>d�?=��>=7#�� �=���>j:�>��D6(?(�?�?s;�b�R�ھj�K��><B?ψ�=��l��|����u�4g=��m?/�^?w�W����&8|?�0]?o�$��N]�;����]:�xh	�I�G?aw�>tҽ���>0Oo?��V?���>"���o�H�_����l��oE�_=�<��>n���Z��j�>�QH?$Hf>`O1>�GS�y��ו����UB?h��?$��?��?��>6�r�PM����E�����?r��>�;Ծ>pO?/c%��J�pa��~K^�ϒ��>|�޽��������,�!��
���C@��f�=ʞ;?��9?l�q?*WU?�7;��6�İc�=����N>�����>�vI�Ż*���O���v���
��� ����>8䞾�P_��o�?�u$? ���oj? �ľ�Z�R?���U>�����%�/��=���$�;�+5=����j�)���6?x��>�i�>L�=?��y��_.�M'5��P�%�Ҿ���>a
u>fE>�>P紽�f���z#�������bۻk7v>�xc?%�K?T�n?�o�+1�����S�!�Q�/��c��`�B>�j>)��>#�W����:&�DY>�1�r�v��%w��>�	�=�~=o�2?�(�>B��>�O�?�?�{	�zk���kx��1�U��<!1�>� i?�@�>��>xн� ��=�>�H?�K�>�}�>n�þ%�2��"��Y���p�>�T�>V��>=4�X��]�x����������?�(e�>�y�?5)_� D$���#>�H?M��=6����*>�>N8�q)��U̸<�>?f[>VUi>����)�A�r�3���P[?(�?�����*����>��?6��>��>I�?�Q�>����ٻ<�4?�]?n�K?FD?�2�>���;w�;��d�.�D��=���>�K[>N�k=��D=u3F��}�߫+��2=�p�=sL̼`RĽP��;�4����=��d=5�2>�ۿ�-K�E�׾?z�L]�{�	�Z񈾔���������	�d������s�x�K�$�'��-W�m�b������l�?p�?.��?�T������������� ��?�>��t�Ţ{��R������3���m��Ŭ��!���O�uFi�g�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@}A?�(���쾔V=;��> �	?�?>�S1��I������T�>p<�?��?�|M=z�W���	�.�e?�}<�F���ݻ��=�;�=$F=���ƔJ>�U�> ���SA�'?ܽE�4>Hڅ>�~"�[��߂^�؂�<��]>Z�ս ;��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�O�\2ƿ΢"�q��=k���>_��p�?w��L�b�พ���j����m<a= ��=IM>|ޅ>r�W>��W>��W?$�j?��>P0>K��vh����ξ�}������:Z�Q����������J�i�߾q���c�Y��Kʾ� =�;�=7R�x���� �>�b�I�F���.?�v$>^�ʾ��M��-<)pʾ�����ل�yॽ�-̾"�1�,"n�J͟?��A?������V�O���W����P�W?�O�ǻ��ꬾC��=ҫ���=y%�>M��=#�⾻ 3��~S��,.?D%?�Ⱦ퇚�[.>�R�_��<�&?q ?��
����>�!?��뽜2^�M��>Kf>]�>���>��=P��������J#?�DZ?��ͽ���L�>�]۾�Ϗ���=��.>�l �< һ�b>��S=�?���H��������<U$W?׋�>{M)�������_7���&=�mw?;�?ľ�>�h?3�??���<����n�T�dW��j=��X?Zj?�b>0�y�F�о�*��h�5?�d?BI>;�^��(��/��L��F?R]o?/�?����,L~�������5�5?��v?s^�ws�����T�V�b=�>�[�>���>��9��k�>�>?�#��G�� ���{Y4�$Þ?��@���?��;<��Z��=�;?j\�>��O��>ƾ�z������*�q=�"�>���~ev����R,�f�8?ݠ�?���>��������=	����p�?;�?�<���q|<���Zl�y���9H�<���=�&��"��=�x8�Ǿ~�
��䜾DU��j�>BW@����~�>�9�	@��Ͽ� ��n}Ͼe�o�Ju?#ө>r=ʽU7����j��du�B�G��uH�닾�M�>��>ٲ��6���V�{��q;��$����>���	�>K�S��&�������5<��>��>i��>�)���罾4ř?wc��@οP���ʝ�W�X?.h�?�n�?q?��9<��v�ސ{���7.G?��s?eZ?<p%��=]���7���j?)\��qQ`�K4��IE��T>~3?1L�>��-��}=�>�k�>a>)/���Ŀ�۶�]���U��?���?dh���>a{�?t+?9_�7���_����*�J/�8:A?�B2>"����!�T$=�����\�
?Wv0?D���2�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?Y$�>��?T��=�6�>!��=����-�G7#>���=w@�Y�?.�M?o�>!A�=�U8���.�=F��GR��2���C�1�>�a?�L?,xb>����1�0�]!�z[ν�n1����%H@���+��k߽r25>ǎ=>��>pE�<�Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��)a~�/���7�	��=��7?�0��z>���>��=ov�߻��g�s����>�B�?�{�?:��>�l?w�o�]�B�d�1=[M�>��k?�s?53o�}�Z�B>��?�������K��f?�
@yu@i�^?x�ֿ֘��ܦ�^��}�=J�=��E>�"���">W��=C�;�d=ˏ$>[�>��i>E�>Pn�>��b>a�R>�
���& �3���2��
G�nK����<�B���s��<��#��nt��M5 �6���{����c�T_
�䝑�I�=:5X?�&?fM?"�?�@���Q> �������r<>Ԉ>vJ?ɐY?{�8?BSA>��B��Kk�}o��A�������,��>'8@>�T�>��>&�>��~=�n>�,�>��>� >cM��:ı��j���p>�g�>���>`t�>E<>��>Hϴ�2���h�(
w�̽,�?m����J��1���9��t����k�=.b.?u|>���?пp���62H?~���6)��+�p�>-�0?	dW?t�>�����T��8>D���j��a>w( �4~l�Ѝ)��%Q>�k?~�f>��u>-�3�Dm8��qP��2��8�|>�
6?\��]:��u��[H���ܾ�N>��></����ᖿ�~���i�KNz=��:?[�?\ɱ������v�A���a Q>H[>�=�=R$M>�c��ǽ}xH���0=k5�=��^>�&?��+>�ǎ=}��>���NP��>m�A>��+>�??C%?��D��,;��DQ-�w>�b�>�>\>MJ���=�f�>�a>�d�q��S��X]?��W>
/~��1_��v���v=�G��f��=�l�=�� ��=��\&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾUh�>xx��Z�������u�$�#=G��>�8H?�V��o�O�\>��v
?�?�^�੤���ȿ6|v����>X�?���?b�m��A���@����>8��?�gY?zoi>�g۾D`Z����>ѻ@?�R?�>�9���'�~�?�޶?ү�?f'I>ш�?)�s?~�>_�x�n_/�6��|�����~=�c;�^�>>k����lF��ؓ�<l��R�j�����b>��$=��>�^�#���m�=�#���M��*Mf����>�/q>�J>�N�>l� ?Yk�>���>8�=�����倾�Ɩ��~V?�p�?�3Q�B>��7
�=}�=6(���&?��?����<���v;>�e?z��?�W?���>`����������𷾐�=��>m�?�8�>�Iｍ|}>Цپƚ޽��Q�>F�&=t��� �~�c>G�>��?F�>F1I=t�<?JF�>��<�J?a�/��g����Z�?Ϫ�>{S:?G[�?2ɓ>c8���D����(��2?s�]�>� �?�?�j�>��q�����U>�p�<K�m=�8? �J? ��6?���?���>�`?n�~>L�=V�ݾ__���A=�}!?z��%�A�b8&�s��w8?�K?�<�>���Agؽe>ռM��´���?�.\?G&?�e���`��þ���<�)�q73����;G;F��v>u�>���"��=��>b4�=�l�f	7�rsg<��=�(�>4��=�6������A,?'�I��������=g�r��D�Q�~>��K>J�����^?�3>�|����݃��}V��ݍ?d|�?��?\���mh�|=?��?��?JU�>���̶޾@�߾))x�9�x�8X��6>�=�>�q�������D���$F���Ž�Q#��M�>6�>�?�`?�YH>(�>�T���7(�����]� ���Z����,*2���'�������J�:4�翾�h��E\�>�����l�>hi?�i>wZ{>��>x
A��C�> �R>7t>��>q_>"U.>,��=T�-<�#׽�KR?����%�'���辽���e3B?�qd?T1�>{i�;��������?���?Ss�?!=v>h��,+�|n?�>�>I��Vq
?�T:=�8��:�<V��k��3���/��>E׽� :��M�;nf�yj
?�/?�����̾�;׽������¾�?�49?�[���@�y������NH���>⫩�U۵����`ԁ�6�������ь�oY%�
>�9?�M�?b�;��k��>����Č�uY�P4�=p}?VL�>��F>��(�[)!��KH���}��/��c�F?>��?\K>XB?2�?C�#?�EC?�/d>�&�>����*��>�8���ٯ>~p�>=6?(47?�@??h�?�+?��=��a�~�����ʾȕ?I�#?�!?by�>��>��<Í������;�|��vֽO�N<��ü��v������=cV>�H?[o��8�M����0k>�q7?���>Ͱ�>�,��A���m�<h��>#�
?T�>�����nr�Y�wR�>&��?�	��B=Y�)>ޣ�=M����F׺�m�=�f���א=�!����:�M�<��=�=�i�Rp��.��:�Æ;;ۮ<iA?k%?��~>x��>{о������w�����>,��>���7��&r��+����?�5�>>QX�?�b�?6�y>;�=�>�A���d��L˫�8X��U�ҽ(�,?N�>�R(?��?l�1?�3?Q=�h����l���C"���?|!,?>��� �ʾ���3���?w[?�<a�����;)�6�¾��Խ�>�[/��/~�����D�SӅ��������?翝?YA�W�6��x辴����[��f�C?s"�>�X�>5�>�)�>�g��%�21;>���>"R?,#�>��O?�;{?�[?}iT>��8��0���ә�B]3���!><@?���?��?�y?�u�>/�>>�)�0�(U�����������W=�	Z>S��>})�>��>��=��ǽ=[����>��]�=n�b>Y��>���>��>K�w>�R�<m�G?���>�\��U����ǃ�6=��u?���?��+?�C=�����E�DI���F�>�n�?l��?�5*?��S�	��=�ּ~㶾��q�'�>sٹ>�/�>�ӓ=�qF='a>��>��>g&��`��p8�MM���?3F?㫻=��Ϳ��l��&"�	����=
���%f����y�o�.=����uҽb���qa������䞾�ͭ��苾��~�ë?RT=S�$>!��=.�!����<R�����=H߅���T=����k�[�v��������:�r;-�o��x^ξ��q?��;?h?��D?V�O>݀?>x�uY>-���x?��J>7����2���f��䐾.,���Ծ��^��
���f>�&��)>a:>�O>��=?o>e)5=c��=�=�A=g��=��>Z4�=	ʊ=��>���=�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�'>Fw>��L�n.��>�k�b�`G���?r�<���Ҿ�j�>7�=i��᷾���=/�2>#tc=�f�t�X���=MN����W=��1=���>o>=>��=F=�����=��=�B�=� N>�۸��$�˴Ƽw�=(8�=3\>y>q�>��?�X0?lAd?tH�>.�m���ξ$:���C�>ɞ�=8�>��=ѡB>���>��7?��D?��K?%k�>�m�=��>��>�,�
�m�	s����$�<���?~͆?��>�O<B�A����h>�M�Ž�p?�H1?V?���>AT��࿯T&�]�.��k���>:��E+=�kr��5U�J0��Hp���㽞�=q�>m��>b�>�`y>�9>J�N>��>��>�x�<�j�=�z�����<`���Ą=o:���j�<x�ż���T1%���+������>�;�$�;��\<��;��=�J�>��>h�>�D�=O���,>�u���pL�v��=a����B���c���~��~/�r\7��]A>{[>��x�B䑿�?�6X>V?>�R�?A�t??�>�4	��#׾�P���d�0�Q� |�=�/>�<�6<�'�`�{N���Ѿ0��>�>�>�B�>s�x>/�,��c@���H={ ۾Cv6�Tv�>Ic���[�}��7Qr�N��zޠ���i��� <��E?���m�=ʰz?d�I?��?+��>+���TӾd.>\�~���W=\��z�P����?��!?��>�o��E�B0��fd%�q��>58�<��z��ꋿz�.�㝐��
y�+?f� �����H�{菿\T���C���i� ��>�g?�)�?�[=��R�+�>���&h���i
??�m?aL�>y7�>{��>=tY����hhC����;.�j?���?���?��1>5fl��*�;|�>��>I?�9�?V��?6྽�?�X��� >v�>=��=I��=�1�=�_>��?'2?���>�k�����d�Ҿ2Mþ|}`���(=7j=8q>�V�>��n>R1Z=��=+��=6�?>���>�XO>��7>x��>�c�>G���G���9?�%	>��}>b<?�8>5=�b�(7����zƽ�@�U�����i�M;+r񻦅�<|IG�A>?8ο5P�?2�>�	$�H:?"2��~�:��A=1�>hӹ�zY�>��s>�r>���>[�>��=�M>`3>�FӾM>����d!��,C�Y�R���Ѿ}}z>�����	&����w��]BI��n��zg��j�N.��O<=��̽<.H�?�����k��)����V�?�[�>�6?�ڌ������>���>�Ǎ>�J��g���[ȍ�hᾞ�?A��?gwr>o�>��R?C?��p�""[��,W�F|���2��M��ed�����L��F��'� �w�S?>�u?e+P?��=�A�>"(�?��-���#�>�'3��-7�;��=bZ�>����A�d�Ӿ?i��zK��LG>EFo?���?!�?�L�T�f�5m�=�$
?1o�>K,c?��?a?�C���,?�g����>v�?�)?�� ?+A?'Ƭ>�>�?��<�g���0���7�<����X��C{�=��P>`��=7�=7�>l[��P�<g\��}Y ��E����Ȼ�r�= �>~�9> ƣ>޲\?S�>Xǅ>�A8?���86�!��^z,?v�"=�X��找d���(�$4>��i?�a�?ITY?�`><A��@��>��>��%>+NX>� �>����G�G&�=tg>Du>���=�.L�迀��	�9����Z�<�>��>ۄ|>2���b�&>^���Fy�#�e>
�R�j)��$�T���G�<B1�m(u����>��K?��?^�=�*�����e���(?�t<?�yM?��?��=�ܾ�7:��RK�kC�9�>r��<`���p���ۡ��';�P�$;��u>���������a>[��22޾��n�T�I����3K=���V=�o@־���A��=��
>�Z���� ����p⪿�J?��j=�Y����T�;h����>[Ø>̮>O*;�*�w��m@�����7m�=���>��:>�X����<G��T�W>�>_QE?�V_?�j�?�!��Cs���B�p����c��.ȼ��?�x�>;h?B>���=�����B�d�G���>ş�>R����G�;��/��!�$�n��>=9?=�>#�?��R?��
?a�`?�*?�D?�&�>M������+@&?҈�?�݄=U�Խ��T��8��F��>f�)?l�B�`��>̉?o�?}�&?3�Q?��?�>}� �A@����>�X�>V�W��a����_>S�J?��>7Y?Ӄ?L�=>��5���f�aG�=�>��2?�5#?F�?���>&��>֗���+�=���>&$c?%(�?$9p?�D�=t�?�\1>��> �=x�>RN�>٧?��N?ٙs?��J?���>�}�<�������'�r���F���x;�'X<�Ry=~���=u�v�����<

�;����&������B�w|��[��;�$�>V�t>_$����0>'�ľ�_��~�@>������tϊ��9��e�=ݼ�>Q�?�r�>�#�/�=l��>�U�>��+(?��?��?+��:�sb��3۾f�L�⠰>�A?���=��l�B�����u�S�f=��m?Is^?GW�8���e?%�]?c�	��k��Z˾rNX��Y��t7?��?�g��J0�> }|?e�j?о�>�]��l�����MZm��T�&�F= W�>�6��[�y�>��0?�(�>C^R>Z_����D݄��龾)�>��?�4�?'1�?2�>bJv�N��z��������g?m��>���WJ)?� ���׾����z������H��[3���Ö��(����'�Rπ�͑ν%��=��?�}k?�q?�6]?���^���]��s���P�^� ��W�*�D�s:C���F�D?f��6��ݾ,ꏾ�Q*=�jv���I��E�?��$?iJ���?, ��= ���Ͼ2f>���ۤ�}  =%岽���<�=�=��D���!�Ԓ����*?�"�>�1�>�;?��k�W|7���*�~�:�2�澾�/>���>1r>���>z�
��P���� ���O<g��T��u>zc?pnK?Ѩn?�?�81��o��F]!��/�o����!C>>�>��>��W����)&�H>���r�����s���	��:=�2?7�>	��>�G�?�?�	��d���qx��[1�|��<c�>�i?�#�>}ʆ>�,Ͻ'� �dU�>�l?���>�G�>]v���w!�a.{���Ľ��>4�>��>�q>70+���[�Z��?��Q�8����=��h?߰���[a��p�>��Q?0&;".d<��>�r�Af!�A(�W�'��f>X\?喬=Iw:>/ž<���{�9���h�(?�]?Z-��g�*�!�}>��!?�$�>@��>S�?~˛>��¾�D�7��?��^?/�I?!�@?��>�=�Ӱ�wxȽ�;&��J.=z�>�Z>.j=9��=	��\�ۨ��D=��=�/Ҽ�J���	<ॲ��]Q<���<4>H�ۿ�:K�M�پ����@�W
�-��H��ງ��r�zs��O����-w�j>��'�G�V�.�c�(��a�l�(o�?�C�?ܓ��B��F���Sx���������>"_q�:>������x-�<��d���Yc!���O��`i�0�e�P�'?�����ǿ򰡿�:ܾ1! ?�A ?8�y?��8�"���8�� >vC�<A-����뾬����οA�����^?���>��/��r��>ߥ�>�X>�Hq>����螾�1�<��?6�-?��>Ǝr�/�ɿa����¤<���?0�@�A?��(�Ļ��V=8��>f�	?N�?>[b1��S�s����E�>r2�?��?�M=8�W�WS	���e?	�<�G���ݻ4�=>!�=�'=����}J>bc�>@��%A�SYܽg�4>��>��!�A����^��K�<~�]>�5սc����?��w��hD�Sg���p�5�<�m�>�7>�g=��I?f���ؿ� ��W�b?ߗ�?��?�n4?�-��`z>gQ����2?�(?�ѯ>设8�U�G�	��P�Ț���
�Z� �V=[\5>�>��#��I���3�N���r�Ὀ��}����=�/)�*�S>
�����߽&{����J�$�ݼּ����Y�m�=�.�>��=��J=��>�X�> #q>ժK?���?���>���>�h������vӾ��6�~�28���l�����X�ξh���R�
��	���2���=���=�6R����4� ���b�'�F�3�.?Ax$>��ʾ:�M���-<4nʾ�����ۄ�楽�0̾0�1��"n�p̟?�A?����B�V����h�0v��b�W?�P����|ꬾ��=o���+�=�'�>��=����3��~S��N?��-?�S��fz��cI�=�ވ�?z�=�;?��>�QR�L�>x�%?㉽ͽA��L>��=\�S>c��>�%3>������Խ}�?T�R?F�⼃w��bf>3X�������=*�C>*�����`��7>��v�,%L�N�ọ�,<�N>�F`?ugl>�5/��p%�'�ξ����m�=u�o?��6?ذ?�v?��F?7^�=<5�������L��M?O�s?�w�=�b>���Ń򾼈5?Dm?��	=8k��	4��g=��$�1/?�vu?�Z?����_���ϴ�{�9�� ?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?p�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�ٕ��Z�?��?}����Dg<R���l��n��k�<�Ϋ=���E"������7���ƾ��
�����࿼ͥ�>EZ@�U�v*�>�C8�]6�TϿ)���[оSq���?M��>T�Ƚ����A�j��Pu�b�G�3�H�ť��/�>���=�$8�>��{�}�;4��[����>��
����>nc��й��	���'��b�>�<�>�c�>�-��������?|���[ο�󛿇�
���S?�M�?y��?��?�?<�@|��戾����<E?�2w?�^?ļ�Q_�j;+�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�a�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*��+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�e.�ν_?��a���p�+�-�H!Ƚ�С>�1�;�\�^'��x��ye����~�y���?A]�?$�?P�O#��*%?=�>�|���Ǿ7��<�Ч>d��>C�M>J:]�6du>(���:�(	>0y�?�m�?�e?������ŵ>5�}?�p�>��?���<ި�>t��=.Ͼລ<���>s�>fÿ���?֗E?? ?�;=Y�>�[& ���2��o2��Uξ��-�)Nq>��M?�kP?�,`>?Q��,�,��(�4�-�G�o�!!��ѽz�.��=>��F>(>и���b����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�6�?���W!��W�}�X����1�_�=�h6?%���|>���>$��=�`v�Y����s� ƶ>�&�?0)�? ��>SCm?3o���B��}8=�Š>�k?0h?Z��n��NB>b?�h�Z���|��>�f?f@�w@�k^?����rտ7W���m۾����U�>��>�A>>��E���=*" =�g@�Qf	��\,>��>�ۅ>��=C��=�J�>�F�>w��@�"����������'�0!.�ʗ+���y�&��7���N�� ޾�b�����=ЫH�l�5�g��v�;(�ɻ���=S�U?'�Q?Jp?d� ?q�x��>�f��J=��#�]�=#@�>�h2?��L?�*?�=a�����d��S���>��'Ň�2{�>E�I>S}�>!J�>��>:�t9�I>�?>o\�> >B�'=ԣ�G=>�N>Y<�>���>�k�>]J<>8�>Yδ��2��ӛh��w�S ̽ �?g}��ۿJ��0��m5��D����c�=�`.?!u>T���>пu����/H?�����&�~�+��>9�0?keW?ܤ>����T��9>���I�j��^>& �,xl���)��&Q>Gi?��j>�9s>��2�^8��wP�<r���hv>Z 5?i��+�;���t��tH� ?޾0�N>��>'�
��Q�1���s��:i��=|=� :?�?O��T&���}r��(���DL>:.^>q/=���=sHK>^h���Ž��H��<=��=�Z>{ ?�N>P�I=�?�>j��B�c��>��~>t�>Ď6?ˋ(?9Ƚ���,������#�{H^>Y��>��{>w>l�P�+�=��>�X>��μrP�5�#��&C�.�G>m����k����&<=����(�=��=6*ｺ�0�1�o=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾOh�>sx��Z�������u�g�#=O��>�8H?�V����O�b>��v
?�?�^�੤���ȿ4|v����>X�?���?e�m��A���@����>:��?�gY?joi>�g۾B`Z����>ѻ@?�R?�>�9���'���?�޶?ԯ�?OI>挑?��s?�]�>�Ix�`X/��3��q���/^=Q�U;�b�>�^>J����dF�1֓�g����j�h����a>|$=D�>G�<8��VC�=1؋��E����f�+��>�!q>˻I>�W�>� ?d�>ҟ�>.T=�r��N〾4����L?.Y�?0-� *���� �[�4�L�*)?0i-?ꁗ��˾��>�iP?�M?��E?��1>D�%�����#����y���3="p>�$?dv�>�V���>po��r]�(��>W�>/�Y�c�־������=�W�>��3?��>�"�=�� ?ݑ#?�i>���>�bE�\7���E����>���>�T?�~?�?�~���|3�����㡿��[�>N>}y?Y<?�5�>\���N���,�<�qE�+���/w�?�=g?��罡�?�'�?0�??,�A?`�f>߷�؏ؾ������>N'?��F�VC6�W�����:��>�>���>(W6����z�z��Z+�"��3x?��e?�2?'$�m�n��便��<C�%� #�<+�K=���7�>M)>	���%�==��>��=^�I�S?#���<8I�=3�h>0�=\��a�u=,?��G�rۃ��=��r��xD���>�LL>���ެ^?�h=�{�{�O���x���U�� �?��?�k�?����h�#%=?��?%?T!�>RK���{޾�྽Jw��xx�%v�(�>���>X�l�(�Z������pF���Ž���ӎ�>���>W?� ?��M>E�>ᩗ���&�>�����1�]�}���8�0f.�m��ʠ��G"�����6¾�v|���>�+���c�>�
?:Pg>@�z>���>��˻�x�>�ZR>��>C��>8kV>�3>Lo >4�<�$ѽIKR?s����'�(��~���X2B?�pd?�2�>$i�ۉ�����K�?j��?�r�?�;v>�~h��,+��m?�=�>;��q
?<Y:=j�*�<�U��x���:��g�,��>�I׽� :��M�-of��i
?@/?@���p�̾b3׽T���p�n=�M�?��(?J�)��Q�K�o���W�S���8h��j���$�V�p��쏿�^��-%��z�(�r*=�*?��?��U��h"��&k��?�ef>�>	%�>p߾>�tI>?�	���1�m^��L'� ���(R�>`[{?���>w�I?��:?>,P?]�K?L�>$��>$o��ɐ�>l�;ej�>\��>�9?*�,?�/?H?**?�ec>(%���F��\�׾h|?�?�/?�?p�?
��bTɽ�Z������v��Ii��҅=�j�<_�н�v���U=ӚR>m��>�f�<]1�H� ��$>)�?3'�>W��>��<�w¾�Ǎ=ɷ�>�n	?�z>V���#_����o˟>&�?�/���a��|�=[�A=W�=V��<
�=zH��_>9�9�� ;��=��+>*>�L[�7'���#��	Mz�� s�`?M"�>>Z>u�>[r��EC�B:�^o>�]>��k>exm>��׾{�������_�
Fs>5��?���?�-8���=��i>�������)���ݾX�:>�(? rU?Au?��?�l?_�I?��ֽ��O��d������Ð��M?^!,?)��>U����ʾ;�K�3��?\?�:a�Ͼ�G9)���¾�Խ۩>Y/�".~����LD�$(�����m|����?���?�A���6��t����^��%�C?$'�>.Y�>$�>��)���g��#�33;>��>zR?9�>��O? 2{?I�[?�9T>5�8�	4��ԙ� �<��">@?)��?Yێ?�y?��>Q>Pb)��4�_���D�� ��ڂ�Z�W=��Y>W~�>_/�>��>���=�EȽ~2����>�3��= Hb>�r�>�u�>��>�w>.�<+�O?�~�>����`�Ǿi�����{	�18\?Nd?	�?n
�mK&���S��ݾ�T�>u1�?��?:�0?�YӾ��=�"=`���Ko��Zl�>:�>�=�>��>$�T>/>uO ?���>O�&=<a8���O�n<)�-�?Bd?�Z>��ſ�Oq��Uq�/����g<"ⒾQ�d����iZ���=fV���
�9B���J[��Ϡ������赾2���o{����>�ǆ=��=�[�=�r�<Əμΐ�<�K=3�<$�=�Sn�i�m<�_7��ջ҈��[	���\<�8I=�� ��V��g?�/�>��+?�R)?���=���>cs_>*�g>�´���,?�F�>�{>�=��£1�L���̚���p0�7#�h�M��N���w�=6=:@>���>��
>g&ýG�=��=nL[�W �3�n�{C�=O��=���<i��=ƾ=EV8=4s?)��>�[�1��%ɾ�"J?��>Ԭ�z}��P[?�#�F���B��+���T)�?>)�?��?�$�>\Y�(��>?������ڪ̽@�@=Ve�`Z>N�1=q�>ǀ�=�
��<��w|�����?���?�P?���Kʿ�_�>��8>u�>��O�4�1�2�_� �q���M���#?f�7�YL;½�>�	�=��Ӿ�CǾnm2=��)>N�3=VD�m�S�\��=�Ł�.�D=��=ֵ�>SE>���=�¥�]��=��_=��==�N>S`Ȼ��%��A���0=L��=m�c>3�.>Z	�>��	?�\-?�Og?D�>�!u���վ<ľn>��=�ӧ>>#=��>���>�y:?�E?��O?-@�>9�2<�ŷ>i��>��+��%k��z侕 ����9=���?��?�Ǯ>�x�<h�!�X���D�����$S?�!/?�?�B�>�U����9Y&���.�!����|4��+=�mr��QU�S���Gm�/�㽶�=�p�>���>��>7Ty>�9>��N>�>��>�6�<p�=�������<� �����=�����<�vż����Iu&�;�+�7�����;u��;5�]<��;���=���>�8>B��>p��=A
���E/>ذ����L�縿=8A��w(B�=1d�H~�B/�xV6�H�B>~:X>�j��U3���?��Y>=r?>���?�Au?�>��R�վ�O���Be�QS��Ը=u�>f�<�\y;��Y`���M�%{Ҿ`��>��>i�>�l>�,�|#?�B�w=��+b5���>/{��O���'��9q��?������[i�`BҺ�D?lF��5��=�!~?�I?P�?���>�����ؾ/:0>H��M�=���(q�e��u�?�'?���>��X�D��Ǿ�A���?�w3��KP��y�V�<��!ؽ^ѷ����>��Ǿ�ɾ�m6�v���NY��~6�q�A�?Y�>�<<?�ƴ?�q�B�r�vO;�(G6�݂R�Q�>�OF?�L�>�� ?EC�>�g�÷��坾.�:>Y�?ӏ�?1��?�L�=%�=E��B��>�	?ǖ?�q�?J�t?�>���>�s�\!>n'��v��=4(>\d�=~H�=B_?O?"�?陽D��a��\��9(U��8�<�=aד>)��>�rz>@��=h��=�3�=i�V>)��>'0�>0�a>�ۣ>=��>������t�M?d�.>���>�N?g	�=�8�@mb��=;��qn���k�D�=7d��P�C���O�aX���/�X2.?˃ۿj�?��=��T���C?ú%�%j"�H2_>�L�>>S���>�R�x��5,R>;R�>�ץ>��>��>FZӾ�>����]!��C�#{R���Ѿkyz>w���"&�~��A���>I�)^���h��j��/��	9=�A��<#H�?����k���)�_��ޚ?�N�>�6?�׌�3Έ��><��>���>�U�������Í�2a���?���? �w>7�O>�Wk?a�?ߍ��H���V,_���H<���H� �h�s���ҁ�fx������d?�E�?��??ZDf���>�u?�D3���g��*>�0�9���2�=�Q�>�ǩ�Tv�B��y�����>�?>�?��?�@��4t��0�>�^?�1?�#�?O=?gP�?�Z#��X?͆�=��?Ͽ?x�/?cV�>�4�>H�:=� >{�=>[�9>):���d�x���K�Y�T=R%r=QWI>�U��[�j=�s�<f���&��<���=���=EJ�L�,��b�=��j=�� >O��>ߘ]? (�>7��>ܬ7?H�k8������/?v8=ݍ������t�������>��j?�?IZ?�bd>|�A�h�B�h>_Y�>l&>��[>�c�>���۔E�GL�=�>J�>R��=|�M��΁��	�	u��T8�<>��?\��={(�4@�>Sq��L����5�< ����g�����PG��O��<ؾ	��>�<`?Î4?�G>��^,���M�g�?f�,?ÈJ?�:b?<?3=�<��@��9�:�m�;����>�H�=��پ��2��	�C��C=��>ξ�_��'@�>5+����ԛV�57��ľ4#�<���<� �����ƾƴ��eXW=9�'<U¾��$��p����O�Q?��,=�p��[��ᾸWV>��z>�ô>�^1�\(�SZ(��������=�ا>KHr=a���SV��qY�	�:�>=SE?J@_?yf�?Y���9s���B������{��(�ɼ��?��>�\?WB>�[�=@���}
�8�d��G����>x�>���`�G�&��~��)�$����>/.?��>��?4�R?��
?	`?�*?�A?T.�>�������9&?t��?>��=��ӽ�gT���8��F����>TQ)?�B���>�?�?s�&?}Q?U�?�e>â ��5@��y�>�N�>$�W� ^��'�_>��J?6��>EY?"ȃ?|�=>��5�g��8����j�=� >r�2?�*#? �?"��>�d�>c�����=���>G�c?���?��o?!��=h�?�s8>o��>﬜=��> :�>��?�M?s?y�I?ɸ�>�r�<d����β�e�y�{e[��`�;�D�<&.�=f�㼽M���Y,�HJ�<A��;,����k���Ҽ�V3�g��U��;I]�>%�s>�����0>S�ľLS���@>a����O���ي��~:��=��>�?���>�_#�y��=̬�>IK�>!�� 4(?Q�?}?b9#;��b���ھ�K�"�>�B?���=��l�9�����u���g=G�m?Z�^?ܔW��"��z�c?�|d?=/��e�2��ž>푾�y��W�G?R�?N�V����>ofy?}Gi?z�?Dt��}p�П��_��L��c�=��>M]��Y��È>f�+?�R�>�>���<~�߾|�o��w��p�?|�?�°?�{�?��>Hro�Cݿa���ц�lNg?Ά�>
���{?r	��Hξ%I"�,����1��k��$����������6�|���.)�;a�<�?B��?!ӎ?H�d?5�ݾ�P�޶I���`�a+U�u���F�l�?��V��BG��cr��*�����k��/�����:��4�?�\!?��+���>�������]�Ⱦ�->�ӧ�����Gu=�ߠ��D�<Pm/=:3u�'DX�ZZľ�+#?eֵ>���>?&<?-�]��`5�)0�v@2��$ ��N3>ӯ�><��>mn�>�r�3�@����=˾}���H������>�si?�0?��g?���]C�����#�B�̽0��%:\>�+>��>JO(����)���M��p��8�������N��=��-?�^>��>>��?�'?ܾ�����Y��u�3��=���>M�o?��>�܀>po���)�� �>y6{?�>��>�	�� 8�򮉿r	߽A��>�ԕ>�  ?=�r>�5�7<�p��i.��ƪH��U�=U�j?]���\9���>V�;?<�h�Ђ���{�>�[ܻ�n*�~����?��@`>I�!?�L>e��>K[����!�,���Ú���(?ab?�k��a*��#�>Ӟ!?���>���>��?�u�>�m¾a��9��?�^?�}I?�@?���>��=Q0����ǽ��%��,=ŋ�>&�[>=+m=���=�`���Y�Mr�s�:=���=?�ʼy���W`�;�1����M<z��<B�4>�dڿ��H�g�̾�G��p�����v��r#����ך��Z�����GG�<Y��g� ��پu����?:\�?�/�����C���T|~��B��7�>YA{�%"��d���4k��ś���d���h!��-P��tm� �i�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@B}A?��(����PV=���> �	?S�?>�61�7K����Q�>.8�?���?nM=~�W���	�Ђe?8�<)�F���ݻ�;�=�3�=r?=j�� �J>Q�>��uHA��Eܽ��4>�ۅ>A"������^��#�<�v]>P�ս-����?ǿ_�zJW�?�*�Jى�
Gn>oxN?��>�ϒ>)]?"�e��3޿5�t�w�V?u��?"2�?qK?� ׾	��>�䵾�;=?�O�>R�0>18��*�g�0�}�>��@�
��
��G6>�
n>i�>�9�V'������C>���2����*¿�z�[�<�j�<2*~<��ݦ�3$�<�����ԅ7�;���1�>��>*H]>8~~>�%k>LH0>��N?��v?M+�>��>��B�L���쾖"�;e3t������޾���0j����}E���K�,T���Eq��!=���=�6R�b���1� �c�b�M�F���.?w$>m�ʾ��M�q�-<�pʾC���ބ�y᥽.̾�1�)"n�_͟?��A?������V�W��X�̓��Q�W?�P�ֻ��ꬾ3��=	�����=�$�>ފ�=���� 3��~S���,?��?� �����<:>�?���5="Y)?n�>\���dʯ>m�$?�3$���˽XO>�$>L4�>߫�>�	>�竾'�Ͻ��?E%N?Q��2L��x�>����f���=\�=�/���6yc>��=�8ĉ�U5����+**=�\W?颏>`O*�����=�-���=�dw?z?�m�>�Fk?HB?���<O���}T�����Cl=o.W?d\i?��>�o��yξ$s���4?c?RUN>Լi�1}��l.��g���?tPo?�0?3W��p}����_6?J�v?q�]�����x��llW�A�>. �>
��>�:���>�>=?.�'����)￿W�3��2�?��@p�?��;��� �=�Q?�T�>~bN�o'ľ�������ҳu=���>M��K`t��"���5�p7?Al�?���>M_�����Z��=<ٕ��Z�?P�?(���9Cg<m���l��m���|�<;ͫ=��QJ"�%����7���ƾ��
�0����濼���>CZ@bP�I*�>�C8�;6��SϿ	���[оQSq�D�?e��>��Ƚ%���9�j��Pu���G���H�]���8�>�nZ=�oʻ��'��c���Z�-߅����>��k<�-�>�H��ƀ�|r��#����d>��?I��>
�ֽ�����$�?�o���޿�������`2?�T�?`�m?:(?bʧ=���?�����)�b?��?��?�G>�>�����=&�j?�_��{U`��4�qHE��U>�"3?�B�>T�-�H�|=�>}��>�f>�#/�x�Ŀ�ٶ�6���Z��?��?�o�+��>p��?is+?�i�8���[����*���+��<A?�2>���>�!�10=�]Ғ���
?B~0?U{�Z.�A�b?�	d���i��#���8�Nt�>w����l�'�=Y����oq��p���و��B�?a��?f�?��Ƚr�,�i�3?՜�>M(��~����ԁ�&�>�;�>�w|>���<��>����*����=�q�?��?�?�X������z>�>y?�:�>��?ƾ�ȁ?��=�_,����q�|>�$A��	���!?��K?`'�>��i=�D���~0�S�\��m>��;��1�o��=�D?�T?�>�����Fj<�q⾉"��Z����&�>�[��V��II��S(>��1>܇>��L}����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�g	?'�6@���M~�(����6��4�=Q�7?�$�K�z>���>ܪ=�kv�DŪ���s�⯶>�=�?�q�?���>��l?�zo��C���2=��>9�k?�z?�ہ�����B>��?K��+���A�,f?��
@4y@
�^?ݢ���ҿ�b����^�U���x�=>W>=�>読��'�<[H� �;�l��}�>K�>�`�>]�^>a7'>2^�=�w]>?ׁ�'m"�9`������T���>����\}~�F�"������A�I뙾/"����!Q=��߽e/�`��
s�'J�=q�U?yN?��o?;| ?�U����>����u�<�%�
�=�>��0?�I?(�*?,��=_����a��X��/W�������>[�<>�}�>	��>���>� u;y�H>	�>>U}>e��=G�#=�W��V=��Q>m��>y��>g�>�C<>��>Fϴ��1��k�h��
w�s̽1�?����S�J��1���9��Ӧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW? �>"��t�T�5:>8����j�4`>�+ �}l���)��%Q>vl?��f>W2u>��3��\8���P������P|>e26?0����K9�{�u�t�H�JUݾIM>�ž>�;E��r��������i��E{="v:?��?i���ݰ�E�u��8��u6R>d<\>�=���=gpM>W�c��ƽ�G��.=��=�^>��?�5>.��=�#�>�ӑ���R��2�>�t>>�(>�=?rl%?�QԼwg��u����-�[�l>���>eD�>ů>N�H�u��=���>X>���h���S�Ȏ>��F\>`���i���}�D�_=.��s��=W�=�8�mI:��<<=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?[J>~��?&�r?�K�>?Hs���/�a����(���)y=�A�:���>�T>����՜E�}z���J���j��,��e>��!=���>2��Ż�7I�=+j���H���Wl�-��>�p>[J>Eϝ>�)?t��>o2�>W�=Pٍ�h^������\�K??���n��۾<��=��^�&?&4?��]�5�Ͼ��>	�\?���?w�Z?�(�>����<��(ٿ�����(	�<&�K>�Z�>HM�>]���|K>��Ծ*`D��t�>R��>�u��{�پ�T��堝�lE�>�k!?��>���=\�*?vP1?a�=^&�>a�7��f���f��P�>�>��?yKy?(/?�о�_:��X�����^S��AY>c;z?ٖ?�~�>[�y�>>��
����h�0����|X?|8m?�����6�>�k�?�bL?,�l?O�Q>�m�z`�v0v�v�>��!?�����A��?&�����h?�O?V��>����oֽI
Լ���Ff��P�?T"\?�.&?���9a��¾���<�#��R���;-�B�w�>s�>���lѴ=��>ć�=�Hm��16���g<��=�{�>*1�=�7�J���#-?tuY������/�=�iq��A�tiq>�?[>'Ež��Y?�S<�M|�`L���E����R�x�?���?��?/ý��f��%>?���?�R?N�>�����߾b���t��v�Z���T>�>�>��������9��ێ���Q���굽gs��f�>�y�>6�?� ?�dM>f�>@Ș�'��u������]�K�s�7�/b.�`�����Ԝ"�
*����ۅ{���>q���Բ>�i
?�$h>Q�z>a��>��һ��>P<Q>�h><��>zpW>�5>��> 3<��н�KR?v����'�b�辎���/3B?�qd?B1�>�i�7��������?���?Hs�?�<v>�~h��,+�mn?�>�>C��Cq
?�T:=�6�<�<V��L���3��*���>E׽� :�}M�nf�cj
?�/?�����̾�;׽������P=)�?�&?��)��J���o��U��NR�o��;�p�&衾��$�{Iq�ŕ��і��(���E�-�&�<
/?Ϡ�?�P��G�p��2u`��D���Y> ��>�ښ>�h�>�l>>���/�5�=�]���%��%y���>;�|?��>�GI?�x9?UM?.�M?��>��>�����E�>�0��3[�>t�>��8?~�,?�+?.�?��(?�e>�8�����d&Ծ} ?~�?}�?}z ?���>���ۨ�<����7�ĥs�`r���=.�)<��ֽ�Zp��#_=�[>�?'�㼙e �n־���>�?Y��>�e�>����1���>i�=��>���>�T�>�����f����>�>}��?C�#��H(=	�8>�.�=�;oL�[5�=3�~�h��=r���˹���4�>�_=�$�;s�к&8<=�H����=�f?B&?T�����>>}��+L���,D�OO�>�x�d(��YRn>�����4��t�V�?o/>վ�?�=�?>e�q��=���>��6���ʾ��Ͼ"p�ޝܽ��=zT5?T�e?o�?�+U?�s9?5��=j�%�+��@��������:?�!,?䋑>�����ʾ��h�3�3�?d[?�<a�����:)���¾��Խر>5[/�B/~����iD�������́����?翝? A���6��w�f���\��<�C?�"�>qY�>��>q�)���g��$�
3;>���>�R?*�>6�O?��z?��[?��U>��8��ĭ��l����Q�X� >�n@?Y��?��?Nax?_S�>�>�+�A�߾�K���� ��"�Ɲ��@~Q=�Y>$f�>&��>Pq�>���=�vŽ%����l?�ټ�=0Va>K��>���>��>��v>��<	}a?4!>���C���s�̾��Y��GC�@3�?�`.?~P�>�ߌ��f�0Մ��ɭ�|�?��?]�?;�B?�BѾa:=�o�=�1ʾO�<�!�>�>~�H�7R}>ZO��Z���G?m�
?��o���1�@�;��������>Fw?�.��|	ƿ��q��`o��m��E3g<�w��z�b����Q�X�&}�=Aܗ�V��f���TX�Yj��F��m��������z����>U^�=���=��=��<	̼$�<R�J=��<7�=�bn��Mj<�E7����� ��y�����c<#�I=�����q?��>y�2?D�"?>�<��=�P�=/�(��C���A?Hq�>'����{[��=$ϾƱ龼܅��h�^�Z��cz�e�>�"�����='y>�Ã>��<x��=v��;�%��R������v�=�~�=p	>p�!>}t�=/�=�+y?7���J���ݷ��׾$�N?_��>l���w�s���S?�ӽ骕�v���}����y?@:�?DD�>`W���R�>>����q�莀�3+0��}�<(��>ůV�4��>X(�>s'�J����Ľ@'�?�H@5}?�~t�P˿c��>c�9>U~>C)P��:-��MR���g���R��D"?��;��;~Չ>G��=�Hݾ����:wM=cD0>��X=���,Z��$�=��v�d5M=��K=*|�>0�C>An�=�ʩ�Y�=�=ݐ�=�4N>��O�*�̡s���*=�:�=s�d>mg->���>O�?8]0?�Rd?@�>n�LϾ�D���I�>;;�=$K�>���=n�B>���>�7?)�D?��K?��>y��=&�>!�>��,��m�}e従���Ϭ<Y��?P͆?�˸>"�P<��A�����d>��CŽ4v?fT1?Gf?vߞ>ש�Яҿ�I���m~�7粼{Z:��.>Su���[�=˧Ƚ�p���M)>���>�?'��>�:>�5�=<HA>�>�Q�>�� >�q�!�<��L�?�V=�Le��=D��=y�=LA���	^<VŮ<8o�:��ƽ�d�=��<�I=;�|�P��=F��>#<>��>���=����C/>o����L�J��=^G��,B��4d�FI~�#/��V6��B>3;X>�}��%4����?p�Y>Zl?>���?Au?��>w �s�վ�Q��:De�VS�Xʸ=g�>+�<��z;��Z`�G�M��{Ҿ���>��>8�>�l>�,� %?� �w=�⾢b5�c�>#z��ů�&�x7q�?�������i�B�Ժ�D?/F�����=W!~?��I?D�?M��>���J�ؾ�00>H����=P�J q��m����?'?���>I� �D��[���	e�=�(?ztڽ�vk�^G4�ҨP�	����|��D��>v��ʝվ�-�8�������8�������Y>��?컼?�T���?��8���<�g�$��=���>�Q?���>)�?���>����V���������M>$E�?���?���?8��>n�=�Y�j��>�� ?��?��?�q?y��u�>�4�=#C3>��>9a�=
Y=��=��	?�?��?�`���: ����R��[X��{w=z�=�S�>�>��k>hF�=1�N<τ�=��3>���>9!�>T��>n��>�<u>8���&����K?�ں=oim>p#4?��^>
�T=���zҕ��h��)A�'HD�HN���r�=%;�*��1,
�"�?�?	?|kп@��?�	�>B�!�֌8?���$[B�	4>�2�>�(ӽ�z�>�vT>�>ݐ{>ǜ�>��>�Y�>|�\>N�Ҿ��
>�5����U�B��sK�.Xվ�x>4C����%���	����%M��H��i�
���h������B��/к��?j�;;i��$����?+��>�p1?������Y��>v��>�׌>�I�����?@���'پ�R�?�#�?;=c>I�>��W?��?��1��3�vZ��u�(A�de��`��፿�����
��	��6�_?z�x?�xA?�F�<9<z>
��?5�%��я��'�>�/��%;�V8<=�+�>J)��l�`���Ӿj�þ�4�{LF>��o?�%�?Y?PV���-;2�>;�>��>��?_�>D�h?�pܾ��9?��>���>�v?؉U?��?��	>�J���3�=� �=��c>����y��뜼�,뽄��<Z>4s>9���&QR>�X>hi㼲h=�!>�}�=?1����μq,�[�m<�{=Z��>��]?���>*��>P�7?H(��8��뮾D%/?�7=�p�����^4���m�ì>��j?~ͫ?�CZ?��d>˝A�f�B���>���>O&>�\>-�>����E��Ո=�'>K>���=i;L�BƁ��	�Wz����<�b>�?�b>��I�1>P����p�%�F>d���uľS_���I��7:�v���	�>7�O?; "?lC�=�5־Y�齡_b��s&?}5?�{W?��}?st�=n��Ͻ/�)�V�JI���>8!A=��â�����T�=��4<*��>+������ob>�8
��5۾�*m���J��\羠�A=j��-�M= 3�BվJɀ�<J�=c>����۬ �x ���檿��I?��u=�����`S����6�>�Ҙ>V �>�d:�sL{�|A�,���ܣ�=���>
�4>�7��8-ﾴ G�8�3>�>GQE?4V_?�j�?!��Ns�F�B�����\b��%ȼ��?}x�>�g?�B>���=������H�d��G���>r��>F���G�6;���/����$���>9?j�>��?x�R?��
?�`?�*?�D?�&�>��������>&?��?�Ʉ=��Խ��T�L 9�2F�m�>g�)?��B����>-�?��?��&?��Q??�?7�>ū �1D@�4��>�N�>k�W�s^����_>(�J?*��>�5Y?˃?��=>~�5��袾:©�Y�=>D�2?2/#? �?��> 3�>^W��N�=���>�Ub?���?��n?w��=��?�'3>�m�>�iR=a�>5%�>n.?��N?2mm?��A?��>/�W<�Cǽ8�o��O��"�U<Y�=ǉ9���<@Wϼ��[����n=-9��84V�ѹh��e���8��0��%Ӆ<NE�>
t>������0>X�ľgk��R�@>���Z���ӊ��X:���=GL�>��?d��>�\#��K�=q��>�o�>����(?%�?��?[h;�b���ھ�rJ�nİ>��A?O��=��l�<����u�O�f=x�m?x^?*�W������o?�Vu?P3�f�C�2.�pNžMB�	6m?��
?mhV�H��>)O?0yh?�v�>��P(��G���E���)��v&==���>��D�&���E��>&�)?��'?EQ�>˨>���ѕ���D3A?[v�?
��?l�?�{o>d�h�����X
�o|����\?�G�>%���rq?\!¼g羇|��Tw|��2ؾ##�����z�e���n\���z�������v�?�ք?��q?�Rc?4�ؾ}zk�Y�W��3Y�o�L����m��:>�O�L��kK�X�x��S��e��iͯ�L�(�����A��g�?�(?*.�ic�>Ⱈ��J�9;P�A>����Y%��=�����=7=cQ=�]h��:0�j��4 ?�%�>R��>��<?-�Z�Ap>�3?1���6�����0>��>�p�>��>���c1���x�ɾJi����ս�&v>qc?K?��n?��-1��y��Ό!���.�gb����B>�v>���>��W�e��1&�4R>�(�r�J��~q����	�	w=��2?��>ސ�><H�?�&?$�	�.n���Jx��1�T�<��>i?� �>_�>�нi� ����>��l?3��> �>Ն��p\!���{���ʽ�&�>[׭>���>��o>��,��\�Af��過�y9��t�=��h?���D�`���>R?CD�:�jG<3��>��u�ݾ!�`�򾡻'���>Zu?=�;>�ž	 �ʢ{��1���p?�2?i����&�lD�>q �>���>7�>��?	sP>YE��7�=�
?<�T?n�N?��2?1P�>�\��%��}���6��=�NI>3�>>��=M��=�h>�8x����ӆ=��>=|h<:�ͽ��"=kd�z������<By&>�[ؿ�ZL���'����⾔Z	����@"#������e��?/���ތ��_��#�׽WZ@�J~��%3Q������[��ƅ�?_3�?dV�?-7�d���C灿n��L��>����K������c���3���ʾ�@��GI��j�עp�P�'?�����ǿ򰡿�:ܾ4! ?�A ?8�y?��7�"���8�� >zC�<�,����뾬����οA�����^?���>��/��p��>ߥ�>�X>�Hq>����螾�1�<��?7�-?��>r�1�ɿb����¤<���?0�@}A?�(�����V=���>9�	?��?>�S1��I�t���AT�>U<�?���?�yM=m�W�+�	�C�e?χ<��F���ݻ��=�:�=�D=����J>zU�>:��(TA�^?ܽ��4>Hڅ>�~"�)����^����<��]>�ս�:��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=� �?\ſ�k�AV�Č4=��ۼұ���~޽T�}=�����%;�����t��=��=~ �=�H~><�G>�;I>��\?O�q?��>l�>Ճ�jX�����P7� �p�+/��������S���E:�^�پ�$�b����z��\ =��=�6R�,����� �O�b�s�F�
�.?Mx$>_�ʾ�M�
�-<�oʾ0���lȄ��ޥ�N.̾��1�	"n��̟?��A?������V�����^�q�����W?�S����ꬾ���=i�����=�#�>��=��H 3��}S�r.?�6?7��xu��UOX>T?@���=�.?��&?{�(=/��>�.?q��8g�<��>!>��=��O>�S:=�:Ǿ�)���*?<''?>������X/�>o�\���U�b6�����=��ڽCa)�ϫ�=��6=�XC�D�� �,��-ż�&W?{��>W�)����]��+��[==��x?s�?�(�>�yk?��B?���<De���S�j��Fw=H�W?w*i?Ƕ>ш���о����p�5?k�e?7�N>Vbh���龀�.��R�'?^�n?�_?�p��Yu}�#��Q��Vm6?�&{?�jj��ӎ�������ԾJ2?5�>�>��T�:��>܅�>�f��fЙ�ڹʿ#�3�>Ƴ?k@���?�Ɛ�6��?��=lz�>>p-
��R���ԽZ��{:���Ы>�z��d�t�#�<���,?�z]?�0�>��N���پ��=Е��U�?��?<Z��2`<}���l��j��*�<Ї�=�����#�����7�H�ƾ[�
�p���0ż���>�X@����D�>��7��0⿨CϿi����Wо�q�~�?;[�>@:ɽͣ���j��8u�r�G���H���d�>�t>a��������{��A;��ؠ�!��>pg��<�>ST�LJ��y���
�,<Ò>���>��>����������?�S���Eο������H�X?O\�?�w�?iU?�C:<#�v�t�{��G�BG?:�s?�#Z?��#��]�l�7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�;�>���?��6=��>�	>����p=z�&>GZ>������?#�X?!��>f��=�
<J��bF���H���O@5�?S>S e?]�@?h�l>f�ѽ>��<M��~Q:�`�D�R������9����B ���6>�D>�w�=��
���ƾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�{t?ek���T�<�>;@���<=NU;k�>t����>��+>�蚽����<���j�~�_?L�?�v�?�D�>�G}?i�i�R0f�P.�=2>o�u?�#�>�/>�H��>a�>-�
���u���#��,p?�@ԁ@Äg?������Ͽ�>��k-���vھ�j�=е=��r>�����	+=�b;���<SM�8�[H>��>&,9>Mip>��S>�=>�A>b�����&�.��(����J�s0�3b�Yu��1�C��%������ԫ�t������,ս̔I�����˃��!�=��S?�C?&b?�P?�Eད�?>����'0l=z�0��ڦ=)$�>��)?B2B?ʇ3?���=���H^��v�c����]���c�>�k>�^�>���>Ӳ�>e(���9?>�@>�CL>ɪ>���<�_�9��6</�C>�ȧ>V;�>��>�L<>�>,д��1��,�h��w�F̽��?A|��2�J�f1��m8������~q�=d.?�{>R���>п+���//H?�����(��+���>��0?q`W?̔>u��H�T��+>�����j��\>�! ��sl��)�~/Q>�j?��f>ɵy>Hh3�O8�; O�%C���*~>��6?N}���A��^t��G���۾�}O>�п>G��{��*?��)~�;!k�a_n=��7?�)?r^���_���>s�Q$��w�N>ew\>�a=Mگ=��O>�B`��Ž�zG�:1+=}��=ob>��?`/>3Ћ=Y�>g|���S���>bLE>�w1>ُ>?��$?"M��]��2���N�'���t>�@�>"�~>�K	>?K����=��>$s\>�+
��/��[���8��:R>�`���X]�$�k��w=@���=�=��=�]���:;�E�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�v�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?fI>���?�s?l�>O-x��Z/�~6��ᖌ��n=�e[;�d�>�W>����AgF��ד��h��M�j������a>��$=�>�C�74��Z8�=�񋽍H����f�ڥ�>w,q>��I>�V�>9� ?.a�>���>�v=Jo��>ှ����T?혙?�H[�s���h'L�M/�T߱�-*?O�7?Y��޾D�>syg?��\?\`k?7�`>�Z� T���4���(־������>���>m��>���=�=1>��ھ��0�0��>�.�>iB�=� 辿C&�G=�����>lG?�*?��>�@4?0�$?��7=X��>�L�����������>��>�e?ς�?'�>��Ͼm�I�����˱�~%g� +>��?Ϥ?���>����H�gx�=[Җ��
>��u? <?h��=t� ?��?N�W?�}x?g��>���!����־|ڌ=�| ?+��a�A�&���c�?�f?IS�>q9���轷�¼���3����?��[?�^%?�L���_�i���0��<V�g����Ep;t�&�^e>�_>�^��:�=��>�=��_���,��M<��=#g�>*]�=x+7�.u���v=?��
������a�>���:�t|&=�ix>��+�L�D?k���I'���>���e��������?h��?��?O��QM��R?0TZ?��?���>��� ^	�-􇾓Pu�J3��"�I��Z(�]��>� �=����>���S��Y{Z��5*<�T�@S�>w��>T�?�?Xd?>�S�>�\����#�T��%���Y�k:�<�4���*�?��H����!���|���*���#�>�����f�>��?�hu>ݲ}>8D�>-��8�>��\>Х�>��>8S>�12>�x>�<i�ͽyKR?�����'�y�辍���@2B?~qd?�1�>�
i����J��e�?-��?�r�?2?v>!~h��,+��m?=�>����p
?�S:=|R�5�<^V������.���"����>�E׽} :�$M�Qmf��i
?./?����̾�9׽Y�ʾ� �=߽�?��;?�"�%�e��S��lX�n�F����8��n����,�k\�:ܓ�/��.�v�}4��bݽ;+?��h?m��fپ����c'����֙�=]�>��>%&>Z]`:�G	�4}P��j��H �s����=�>tu?��>nqC?��:?�G?��K?f'�>3h�>����R7�>C�<�&�>S��>�7?�U.?� 1?.P?P�"?�bT>�m��<����־d�?z�?͡?O�?���>A	���<½vZ%��c����j��I����c=Җ8CoĽ_�I�,~=`bV>�s?c5�d8���Rm>�/5?�#�>��>�b��t���=5�>��	?奏>�����q��V���>�:�?��	�l��<�(->���=k������:fG�=�Pۼ��=*9I�0��Ў<g��=�@�=�K������7Z,;�s;2$�<�P?��?2�>�?>���S���L���>�mB�Rb󼍼7>�7�����Q^��.~�g�@>"�?�%�?�!>�7�=�;�>�|׾pM��|��(���7k��>��[?�H2?;�?1�*?��C?�M>P5�4���S����	�M�=?v!,?��>�����ʾ��Љ3�Н?j[?�<a�
���;)�ǐ¾��Խ߱>�[/�_/~����;D��������t��4��?쿝?�A�M�6��x�׿���[��y�C?
"�>"Y�>k�>M�)�y�g�m%��1;>��>kR?d"�>��O?�:{?0�[?nT>A�8��/��ә���2���!>E@?屁?��?�y?�v�>��>�)�A�mP��������ނ�kW=�	Z>���>'�>��>���=UȽ�Z����>��Q�=!�b>H��>y��>M�>��w>�o�<�5H?F�>����������Ex~�pEJ��Ct?�w�?u,?Pi�<RT�J}F�D�����>��?汬?�D+?ؤU�-"�=Iɼ�l����q��S�>�з>�U�>j��=��4=�@>U��>���>T2���ڋ7��6R�.�?��E?�T�=�uĿ/�k�~�Q��톾�G�<"Ơ���b�1$���[i�1yu=�꛾j�� ˮ���S�IL��JM����������Ҏ���>���=ć>�u�=���<�9�.��<aBO=��<<�+�<G���;cɻ��F�'�?�Cɽ;� QW�6y=SJֺ�A���Hq?��7?gw?6�C?��>U@>!)=(��>��ύ?(tk>S�߽�(������Z��k����ɾH���c�U_����6>jὨ��=ٵ;>��?>���=��<��_=� �=�^=�=�>��=!H�=`)�=D< > >�=w?d���������P�d���;?껑>q֫=��ƾZS@?,�<>]@��ɕ��Ź���~?Z��?6z�?�?I�i��d�>����}(��L��=�)��D�1>�i�=Ի0�d�>�aJ>�7�w3������
�?v@��??¯��xϿ{/>�I8>	�>>�O�ۓ.���8�b��pC�<x)?ũ%��Z�$�r>��=�ƾ�2��Χ�=i�G>��	�'�'��9Q�O]=	���\����< ��>�j1>s��=�A���=�B�=f�>s�y>FF=oB*���ü@��<*��=;8?>P�Q>�2�>�?	0?d?�պ>:�n�7�ξ`!��t��>(��=r*�>t�=��@>�M�>@�7?SD?0tK?�e�>��=��>�y�>�,�n�m�s� ����<�ވ?�f�?�A�>�X<_�B�����4>�c�ƽ~?M)1?� ?M�>U;��⿵"����R����<j��<�I%>�ח�#߶�u�¾炔��DF={\�>�Լ>/�Y>�|>�d�>37W>���<�U�>t>�>S2�>e�Q<�ٽ��|�Qr�&��=��>��=�����`w��;q��=P#��)M�;ޒ�<]�x=+��=��>�<>Ĭ�>[��=��D/>������L����=�G��,B��4d�?I~�/��V6��B>�:X>c|��4����?��Y>Ml?>`��?�@u?��>����վ�Q���Ce��VS�zɸ=��>)�<��z;��Z`�U�M��{Ҿ[��>Vߎ>�>q�l>�,�N#?���w=��Pb5�q�>�|�����J)��9q�@������li��]Һ��D?�F��@��=q"~?��I?X�?؍�>�����ؾ;0>�H����=j��*q��h����?'?��>�쾟�D��2���0���	?8���[��|^��$������༾cά>���m��S���杞�P�M�&�m�׼�>�o?���?�C���lU��_*�<4��}�>ìm>�?�=�h?���>�b�>8�����=2F�?�U�?��?[�=VϹ=+����`�>rC?�^�?e��?�cr?��9���>�"k:�{%>������=�>ۼ�=��=]s	?<j?nR?(���ņ	���辵@��\���=��=^�>8��>�p>�^�=�qs=u��=�g\>�ә>^،>8Ge>��>bɇ>q楾��
�S('?*��=�؎>�q/?(��>݈]=�姽E��<9P�)�<�{2�������.Ձ<T[��0�D=dД�ģ�>]�ƿm˖?��J>�8���?���,xB�^M>�Y>O�佘��>'�E>}�z>në>;!�>��>D�>�)'>ɎӾ��>�V��� ���B���R��{Ѿ�y>�����2&�����$��~J�G���4���j�����M=��b�<M@�?�\��-Mk���)���	?1�>�5?p������� >t��>�(�>(����������?�T�?u��?��w>���>إU?E,?5rj�`�罌�Z��x�GGE��gT�P�j�G'��ܸ��62�]佅Sl?�C�?́I?��d��H�>�|?��/�F������>&)��H8�R:�=��>⬾i�Q�܏Ҿ�"��."�daX>�7p? ��?�#??DN�ކ_��>�=M�??���>ȝr?q�(?�wX?!齒�%?�F�>rJ/??�&?7?��?�`&>���E|཈�?'W�E1��灼C�);')�;��#>��i���]�=ڶ=l�^<�
�=�7�K.�=��|=��R�p=h�=$��<�L�=�o�>�p]?r��>{T�>��7?�%�?�7��b��� /?�7=�7�������;��e���>pj?+��?�Z?5�e>��A�
~C��6>j��>8%>��Z>ux�>8��$-G���=��>�>�ɡ=�EM�x����	�����8�<�[>��>�=|>��V�'>so���=z�Ωd>�Q�L���&T���G��1��v��X�>��K?8�?C|�=aY龰"��CEf��()?�Y<?�FM?L�?�=	�۾��9�6�J��I�7�>�é<�������5!��g�:�r/�:��s>'���-��U;�>�W�����1,D��x#�N��>p��' �1\(�I��4���53���!���*��ƾ�f4�*���%��b�??���=`��u=������>ƶ�>�p�>"����,½�	c��;��&H��z�>$�?>I8=�v��rtD���*��7�>8PE?FM_?�d�?'��ks�L�B�����a��]�ȼd�?B��>f?�'B>0'�=ǡ������d�G���>��>����G����E&����$����>3?;�>5�?��R?��
?:�`?�*?�E?$"�>�+��N��]=&?���?=
�Խ��T���8��F����>�k)?��B��ɗ>i�?	�?��&?�Q?Z�?��>�� �}?@�9��>�N�>5�W�(^��	`><�J?�>�Y?dʃ?��=>�5��袾!���f%�=�>:�2?v1#?��?��> ��>����	�=��>�c?�"�?��o?���=�?�1>p��>�w�=���>Ey�>��?�8O?ټs?0�J?��>�z�<�<��I綽�-s���M����;��I<sy=q����s�������<���;Ҷ�υ������D��2��<��;+#�>#�t>8�^[0>�6ľ�E���HA>����}��Sq���9�+��=j�>H�?|͕>�#��X�=��>���>���q (?��?�?*@L;��b�j>۾�9K���>��A?pc�=Ql�=r��m�u��_h=��m?U\^?b�W�6q���i?�o?4�?2E�:��Й�%��ǓD?)�>wrV�IV�>5Ek?e?W?P���Sg�7B��*�Z�bXҽ�5�<��>���eDG�B�h>�48?���>�/�>~2<������	���lX?8�?w��?9ɂ?b9�<��{��)ݿ�D��=����b?�w�>�社ۋ?�fs����%ԅ��Ԑ���ƾ܅n����� L��b�̾�Y��遾�����a=37?J�?݉�?\?�j��8�V���a��p����L������=�9���6�pj?�9Rf�u���������Ύ�A���3�@�g��?�N%?�g1�V*�>%����_󾚤̾O�>>돞�Hd��i�=������=q+?=�%i�	l3�aD��Z� ?I��>2��>�<?�][��><�2��&8��?��*�->@�>�[�> D�>G�9�=�.�0���ɾ� ���ٽ}�u>P\c?�K?�6n?�7 �K81���,� �R�5��֨�{F>"�>��>�UV�-���&��2>��cr���m��r�	��k}=�2?��>Gz�>��?��?22	������x�g�0��o�<�#�>_�h?*k�>���>v�н|!��g�>z�l?c��>B��>�"��p�!�o�{��!ʽC��>�_�>�0�>��p>2~+��y[��j���s���9�.^�=��h?�e����^�<�>�7Q?�&�::{j<�2�>�u���!����Φ*��?> ?�z�=�h<>��ľi��-�{�X�����(?�>?ģ��u�*��3�>%�!?̑�>g�>���?�|�>�¾i�B:�?�^?x�I?=�@?���>�=����ȽK�&��R,=Mֆ>��[>�no=���=�"���[�Y��lWA=F-�=��׼����Hy�;)Ƴ��S<;z�<^f4>�rڿ��I�	泾�4�J��Z��n���\��M|��(�����e���?��R(�L|ҽu~h��}]��V���v�9��?��?j�.�V]�]���;|��:�1ƅ>(�~�)�
�:���׽r������	���)���I��d��[�F�'?�����ǿ밡��:ܾ.! ?�A ?�y?��B�"���8�L� >�C�<�-����뾥��� �ο3�����^?���>��/��[��>祂>�X>THq>����螾�0�<��?)�-?ڠ�>��r�0�ɿY����ä<���?-�@-{A?D�(����V=���>��	?��?>9W1��H����U�>�;�?���?0qM=��W�e�	��|e?@�<��F�^�ݻ��=
@�=B=.����J>�Q�>V��JA�	?ܽQ�4>dօ>�"����̊^�1g�<��]>��ս�!���O�?��^���b��%��=���q
>|�K?V��>�y�=��.?+�O���п�9i���g?��?���?�W/?ٺ����>N�վ�|I?3'?Cl�>�����w��]>]�=��0=mվ߷F��`�=W�>�n>��E����{Q�Q����=/� �L�Ŀ���24�W�=�҉;&��;�=��.�+��<2څ�Q ��@��=p��<UcD>�,l>�T>��!>��T?� ~?8��>��>�3��ʡ�����^���3���W�Oa_�oBd�����DC�ǥᾜh�t��Q�漾Y =�R�=�5R�H����� ���b�k�F�=�.?Ou$>��ʾ��M���-<�mʾT���L��S祽�/̾�1��!n��̟?��A?���o�V���1Q�<{��,�W?�N����묾F��=�>�==%�>؎�=Y�� !3�TS���)?�?�,��������K>�l���<W�?L��>�B$��j�>�{&?���4�׽/)^>w�>A�>���>�g>�ګ��Ƚ�?�L?��޽ո���}�>�	¾��S�	v=�]�=�,�R���P>5�>�(-���<?�a���=�]?;��>?�.���Õ���4+��& ���k?]=?*�>ʙo?�lA?�Lf<;F�;�_�wh�s�<uN?�@r?��=-��<|�־c3ξl.?6[?��7>{|����).�[���\?Ćz?K!4?�`Ǽ�1q�S{���O&��'?(�v?�q^�1]���I�wW�oX�>���>���>�9�8F�>�8>?GQ$�RG��o����4��Ğ?��@���?s�5<�&����=I[?���>k%O� �ž�^�������j=ܘ�>N���&v�D��9$-�G�8?�\�?���>����CJ����=Sٕ��Z�?��?k����g<���Bl�n���q�<vϫ= �v="�8��d�7���ƾz�
�۫��/뿼~��>;Z@&L轡*�>�C8��5⿿SϿ1���[оqUq�w�?��>��Ƚꛣ���j�(Pu���G���H�æ�����>��%=�[���7��I���l$�wp����>���+\�>�2���d��7��F�=��>>|??)�>B�ýq�׾��?ss澾pӿ������о&?�Y�?e֐?�d0?�'=���|]��(��y0X?�_?�S?�vO�)s����%�j?�_��xU`���4�tHE��U>�"3?�B�>T�-�\�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ss+?�i�8���[����*�!�+��<A?�2>���I�!�B0=�UҒ�¼
?V~0?{�f.���_?�a���p�su-���ɽ�ʡ>ˢ1�F�[�9��7��9�e�����{�D�?"d�?t;�?�����"�i�$?�>�o����Ǿ6D�<l��>�-�>�O>Y�U��w>T���s:�A�	>{y�?,h�?? w��4ᦿF�>��}?``�>�-~?�.��D�>�t�=Vq޾����wt>+�N���
�͒4?�cH?���>o�>��=�(�LK�p-��s߾�,���=�R?ShJ?���>ݭ;��v�by�k����ֽ�0'=����N�<�'G��]> �$>��?>����)����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�[�?���*�J�6DM���*�YU>'���'!?4���>@�>5��	�p��T��j�s�դ�>vU�?I��?�<�>y�?�o�5�d��/>���=��@?�/�>1��ە̾�&m>�4�>���m����ձ�5a�?$~@��@�#h?�H��ֿ֬���+�c��:���>��=�ݜ>��.�M)�;��
>��=���=\��=���>�"�>���>^�X>/�=�`�>.���| �ޣ���B���OH�-�!������y�5�)���оy	�@r���+�@����;Tiv=��Ľ�2�����=�e�=�oS?��E?A�i?��?�/��_/%>���Ź�|`6��}�=��>8�2?H$D?��/?
0k=�u��j�[�d"~�%��U��� }�>V�:>�6�>i��>�^�>�����>>US,>�K>K�=�/R=������<�T>��>�}�>Y��>;O<>â>�ϴ��0���h�.w�33̽C �?M�����J�0���3������څ�=�^.?4t>X��a>п����q-H?u����*�ܲ+�I�>ʾ0?�dW?-�>���t�T�R@>�����j�x`>X ��ul�؉)��Q>f?��g>��v>�4�Vi8�.�P��尾�#{>u86?)����:��>u�AH�uܾ3�N>��>��N�H��������~�lj��jx=s:?��?�����߰���s�k���>dR>�^]>��#=%��=�0L>�d���½n�G� 51=%*�=;�]>��?lP/>��=��>MΔ� UT�&�>:s>>�/4>��>?V�$?���n���q����0���o>d��>�>z;>	J��=�z�>oX>7�ּ1Ά������8�G�X>�fh�7^�����g]g=�፽}��=S�=��tN=�f�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾQh�>yx��Z�������u�o�#=Q��>�8H?�V����O�d>��v
?�?�^�੤���ȿ5|v����>X�?���?g�m��A���@����>;��?�gY?soi>�g۾?`Z����>һ@?�R?�>�9�~�'���?�޶?֯�?�H>��?3s?�=�>�[u�'L/�E��a����"�=\D;$x�>�>%���)IF�˓��\��S�j�֫��&b>
:$=��>������ɇ�=z��3D���+g�ŷ>�Hq>�I>X&�>/� ?�X�>pn�>8H=ux��B���롖��)M?�ː?1�:�?lg�S����c�Z����v?@`?��˽V͡�[�>S�Q?��~?��??��A>�)��Й��*������[�*��5>!]?�&�>1XԽ�&�>�/��=���h�>�o�>��:�پ�]��`v>fm�>�?�1�>��[<��&?�$?�5>~�>�A��ᕿhK��0�>��>@Q?z�?�?���*:�U����"��hYR��}>��z??��>�R���礿��g�\�ٽm)��_�g?f�a?���w?�Ï?d�G?��M?�@>�nW�k1�F�D�D��>��!?�$�ñA���%�bL��1?��?Pb�>���I�ٽW�˼0"����Ӵ?c\?��%?R��y�`���¾�<�#�H�Y�QJ�;�`=�s�>q>�����V�=�M>p�=�#m��}6�o�a<gr�=,�>�Q�=�16�簋��7?9Խ�T��5��>��a��X��8�=���>Z�ھ��9?j&w�KɅ���𘿿罜i�?��?��?�⽉�K��WY?���?�?me�>���s���o��_��(���.߾\^>᦬> ��'���X���_���65�&="*��y�>�{�>xo?A?R�N>'��>�����~&�������h]�@��K 8��.��s�Q���6""�1���m��f[{�	ԙ>*���>�t
?X
i>jz>+��>�c����>CN>�[~>��>�V>v�2>|�>N�,<J�˽�GR?������'�������-B?�nd?�*�>�Xi�A���V���?���?Rp�?iCv>�|h�G,+�l?aD�>O���m
?�x:=������<W�����4����饎>�׽Y:�PM�	cf��h
?�+?sč���̾<V׽N,���Hq=��?��%?�(���P�p�n�J�X���Q��S3��Oh��ԝ�d\"�Cp�XV��|D��t����,*�� =�!+?��?y���B�pH��\�f���>�Ra>��>�I�>�D�><�>>��	��H1���\�Hs&���e�>��w?��}>i{H?ӫ+?f\D?�]?�~>���>U$ؾ�!�>�l���>k_�>2�6?��?�;?���>�$?�'�>����Ro��Ⱦ*%?Z�?�s?���>\K?n��}G�<��;=MՑ�F̀���<Q��="E�<I���k]�>��<aCS>���>r�;>�S3�����y->B#�>K�>g8x>���/���i�>�d�>��?��'>k��hO��X�@��>D�v?<q��vt�<dZ�>���:�5�L5���>����=�락�k}<��s:V@�����=�9��ռXJ�=h!=�K>֑?��?��>oT�>�q��9��
��h�>��>Щ�=i�/>d����ڇ��0����9���q>[��?���?�<�=C)�=޵�>�G��EO)�uH����޼�6>��<?ށo?8��?Mv?
]*?�*�=ϋ2�������^��2�(?y!,?L��>���Ųʾ<�l�3���?�[?�;a�1���8)�P�¾&�Խ��>�Y/��.~����ND��9������������?i��?��@��6�y�㾘�J\���C?�%�>�X�>��>j�)���g��$�]2;>΋�>>R?_�>��O?��z?�\[?^%U>g�8�{㭿~���/g7��� >+8@?x��?�֎?��x?t�>��>l�)�۳߾N������m�r���#zW=t�Z>�~�>��>���>s�=��ƽl�����>�*o�=�b>WZ�>:��>���>yw>ow�<�`?p~P��	��X�wq���]�'R��D��?��?v|?��m��_�iT�����X��>4>�?˷�?�T?EM���;=i�<��ɾ�����i?��>k(>}z�>�c���=q�?9��>"�Z>t$C� qD��������>IQ?D �=n�ƿ�%t���d�8Т���<�U���;Q��ޤ���O��8�=�������!����=[�膦�PO��0n��8���	i��e ?��=| >+��=�uM<�����-�;�08=�m�<��<�K@���=Z1�'u�dK���g�C<v�1=��u����Vxu?S�)?k�?УH?HzJ>
��=�����t>\���W?�+�>r��3����"�����31��'���P����.^��猾��)>��e��!%>p�<>�i>#�S���)>�"�=��7;�E��Ɇ=���=I�=��b=�-3>+)>^C>�rw?w˅�(v��&��k׼�V�U?��d=���<�Aƾ5a??���iڔ�v�ĿZd�դ�?d4 @�W�?��?�����>���&?¾ˌ5=�� �Dų�EK:>/��X(�>MxH>����6���l�����?�@=<g?R
b�]�ǿ�|	>p�9>�/>-M��u �$T�ׅQ��eP�5�?�;�JC߾�=�>>ќ���Ỿ?�=�q>�/t�P�sP��Ei=�]w�3�8=a�<��>�~a>ı�=�!�	��=A��<HR@=�4>�͏�a�r��+ǽa�!=���=�t>��Q>�~�>��?�\0?[Ad?%N�>$n���ξzD���p�>�3�=�B�>tK�=ŘB>匸>+�7?ޟD?7�K?�{�>�?�=[��>f��>Ռ,�v�m�G��ͧ����<���?�ʆ?/ٸ>�Q<��A�<��}O>�[:Ž�s?M1?�]?���>7*������ؾ&�E��߹��;��~>r|���o��E��=�Z7�dQ���l>n�>�q�>]{�>��r>���=��R>aX�>�2>�K5;Q1��u�<��=V�8=L�=�/�=�f>Vʒ=ΤZ;ϙ��J�v�s�Qٽ�����ֽ�>s�7��=��>N<>��>���=����C/>�����L����=�G��N,B��4d�}I~�(/�^V6���B>�;X>�}��/4����?d�Y>�l?>���?@Au?F�>� ���վ�Q���Ce�!VS�7˸=��>d�<��z;��Z`�X�M�6|Ҿ���>�ߎ>{�>��l>�,�1#?�d�w=��Ia5���>|��8��L'�9q��?�������i�.�ҺȠD?DF����=�!~?*�I?1�?,��>���E�ؾk;0>H����={��+q��f����?'?f��>��/�D�H{þ8��@b?��
���U���S���9�s�w���Ҿ+��>��վ{%��1�~|��א���JB��.��`X�>j�.?��?X���s�I�.��A���h=\��>�U?�u>.8?�%�>X��⾭>��Q3�=l�{?���?u��?�g>��=�߇�h~�>�< ?��?�E�?�v?DoP��L�>�q�<�">�� �h@>o�>*z�<�Ȫ=�?q�?�G?�F���Y�]�x�����>�K�@<>O�=�>0*�>a��>��=���<C=S�n>�x�>ȓ>�Od>��>6�L>𖺾����H?�>��l>��J?��}>�=����N�om8�諜���_���;���Y�W	R�l���1��^�N�EC?��Ϳ�?ɽ�>FU(�jG?D����=�z
>��>7����>��>��>N��>4��>�i>���>/?�>h�Ծ>���y���A�7�L���ξ#�v>+���T,�l�
�œ��(N�ٸ�v��%�i��(��5�?�#Ǘ;���?���{�g�TJ%�Mc�g�?�-�>�7?.4���h�>���>켊>������#,�ھ�̌?+��? mn>��>�e\?�?JVf�J߽5�a��ks��rD��[��ph�o��Iǁ�Ҧ��)Ƚ�La?[�{?�C?ړI����>��x?��2���{��eo>tk5�� 8�g�=6ޭ>C���f���WE���ھQ;��Ĉ>��~?��?uM?�<_�2����>Ȟ?x��>���?D��>A�o?%w���U?�P>��>z?�x;?� #?�7@>n�޽���=�d=�>����)֊�rˍ��0i�C�k���=/ٴ<j���\����l=�ڝ���"�}��I*=��|��=>��.`���=�x�>�:]?���>2Z�>F�:?�S�k�6������.?Y�=��~��t��񱞾���S�=�f?EM�?�sZ?�p>��A�S�>�S@#>���>�w'>��Z>B+�>�[���P1��m�=P�>E>ٹ=q>�����	O	��&��M�<Χ%>b��>x5|>�����'>�k���(z���d>U�Q��κ�	T���G���1�{{v�R�>%�K?��?d��=GX�+���Df��-)?[<?(JM?��?�=P�۾��9���J��E��>�A�<���񽢿g#��^�:�f��:�s>�!����ľU�>ȟ���޾FSW�B���Ǿ�R���U����:������$���J�=g�=݅��+� Z��ؐ��*|K?��=�t��*��%��� Y>;��>]��>���� W��2��O`���=���>[t�>�fj<����<�9��P:�>�QE?�X_?�i�?6 ��`s�R�B�����e��@-ȼ��?4r�>f?�B>a�=��������d��G�[�>���>0����G�:���+����$����>9?d�>z�?J�R?��
?�`?)*?�E?A&�>e�������A&?;��?�=&�Խ�T�^ 9�F�~��>L�)?*�B���>Q�?��?I�&?A�Q?ߵ?��>ѭ ��C@�1��>�Y�>N�W�Nb��%�_>��J?3��>2=Y?�ԃ?l�=>
�5�颾ש�U�=q>W�2?6#?<�?e��>��>�\��N��=��>��b?�/�?�Oq?���=K�?��/>���>�2�=���>0�>ֱ?��N?*=s?K�I?���>��<���������l�gA?���];��"<D1w=���{p�����<�4�;���5�d�7m鼅?�L���q�<�_�>.�s>�
��a�0>�ľbN����@>����O��܊��:��޷=~��>��?	��>yT#�+��=﮼>J�>���36(?>�?�?{#;V�b���ھ��K�{�>�B?���=9�l�Ȃ����u��h=<�m?:�^?ҘW�y$����f?H>?�[2���,�RD�$ѽ����??Do?ֱ>5�0<��?(7�?m��>�v=�������Fl�������<1z�>�ӈ�,Y?���>w�M?pN�=scl>�b��сھ}�0`���'$?���?_r�?Ø?ⶽ��\���ܿjY��1���Z?a��>����K�?�,c�O�I�����6��1���6����k��z���
K������ ���=�%?m�?�l�?m�R?&�
�/m���d��a����~�(��<����~�p�j���d��&��"�:�k|��������;�ك���=�rȷ?�g4?r�Y��o?����I����ݵ>hf��"����<�3�+!=,��;�Z��Bʂ��Eݾ��C?�R�=$��>��P?�w��-�	�G�������|V>��>ɑh>iO�>��������X˾ޅ!���<8Bv>�wc?��K?�n?�q�A*1�ɇ��ސ!���/�Z����B>As>�ǉ>۠W�zt�R6&��^>�!�r����qx����	��=��2?d,�>/��>�L�?v?~	�s���nx��1��'�<G6�>=&i?�F�>�>��Ͻ�� �,��>*�l?��>��>闌�[!���{�-�ʽ(�>��>��>��o>Ҭ,��#\��j��I���m9�mv�=�h?������`��>!R?��:<�G<�|�>Z�v���!�$��H�'���>�|?��=n�;>܁ž�$�Ƨ{��7���}?+?���q$�+ʟ>�7?�?��>�M�?�VB>	I�VG���z?�7]?��J?g;?V��>�-��.h��kѽ�s#���i<���>��>���u-�<h�n�(��I���3�/=�ƨ=�(���%��@�>=���=�,���߫��e5>ylۿ-@K�@�پ!���(?
��∾f��|q��h���i���5���hx�K��No'��/V�K?c�8���q�l�f��?�?�?�O���'�������������^��>{�q���p����K��J���ྯڬ��q!� �O�\2i�_�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@_�A?9�(���쾊JN=-��>k�?�?=>5-.�$���k�����>���?�#�?�8;=�W�� �(�e?�LL<#F�r0ڻ��=,Z�=V=���E�H>��>�5��c@��8ݽ��3>ː�>�r����e\����<�j\>x�׽�w��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=����ƿB%�3���=]Ш�T \���载M��bYO�����9uo���罥jk=;�=VGR>�R�>��V>��Y>�YW?i�k?-	�>�}>J`�ck���1ξg�<����`��:��U���壾m��=߾�Z	����A���ʾx =�\�=�6R�z����� �2�b�V�F���.?v$>�ʾ-�M���-<'qʾ����k焼�ॽ�,̾A�1�	"n�:͟?d�A?������V����\����}�W?nO�.��9ꬾ5��=`�����=%�>h��=���� 3�J~S�V�1?f�?�����s��>�+>i��24�<W].?�I�><$���?�>��$?��-�s�	�o^W>0�D>�ϧ>���>>H�~�ѽ��?Q�U?.��FT��X��>�����z�)j=2.�=R5>��I"��;R>1 �<�ڋ��9���:����=c`?��>8kC��n־����t޾4�㼂��?��C?�5�>b��?��i?��7����/i�� �W;�=H�1?�`m?���=�{+=L�־��U�?r.?X[�=�_��v����4�I�<E?�v�?�?"M��È�a����3��!?�/}?�&��^x�e�L����c6>�!>�n�>`@�`�>��Q?T3�����4԰�*;_��t`?�Z�?�M�?�1�6(Q���<>�>�?�>~z����	����=�H���(�=�����J��10��)��ww?h��?��>���/����=�ٕ��Z�?l�?z���>g<B�� l��n��G{�<�ͫ=3��H"������7���ƾ��
�C����ῼ��>BZ@�S�9*�>�C8�E6��SϿ�� \о$Sq�n�?倪>ӢȽڛ��5�j��Pu�k�G�\�H��������>ͤ>+9�������{��u;�;���{�>g��@̈>!�S�p۵�
����'<�{�>I_�>��>O����p�����?�;��6ο��������X?%i�?�@�?�?��M<*	v�<{��|��;G?lHs?��Y?�0!��\�]�9��k?����{`��k8��wH��
K>a7/?���>�*�kH�=��>}�>/3�=B_0�$Ŀ�����(����?���?���9��>M�?!s%?j������32��&+�`�;�yE?rB>��þ����q7��D���F?ze2?��H\�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?_$�>��?t�=kl�>'s�=J갾Uc-���#>L+�=}?�^�?�M?AZ�>Щ�=�8�R/��XF��ER��(��C���><�a?|L?�@b>�㸽2��� ��}ͽ�b1�S�lj@�P�,�X�߽�05>��=>t>B�D�iӾ�1?�
�eؿȎ���,+��@3?���>�\?��q�s��t.���^?�"�>���i���-������f��?���?�?��־�`���>m#�>�ԅ>vC̽�x��^˅��=>)�B?wy�̊���n��7�>�^�?��@i��?\�h� �
?���ć�륀�c��p�7���=�3?�N���>���>�Ҫ=1�y��'����t��b�>9�?2��?���>
�i?`(l��<��u=3�>�!m?��?�������T>�?c��N�������V*b?�=	@EB@>`?�����Nտ������������3>�|�=#(�>��c�do#=j�>8�#=�߼O� >�ư>�!>v̆>.jA>��#>U�2>�u��
6����@H��M5�a���w0�i�o����)5W���S�ܾq����fh�p]ӽRIǼ��~�FZ-�ʗ���~>�Qp?iO5?�_�?}?1�����>)��J��=�9!�lY��u�>��@?3�p?�-X?5�>럾j�A��;���!¾���l!�>Ձ">6�>5D?�4�>̯���!�>'-�=o�>���=�t���ݽ�w�NE�=��>3ܾ>ҽ�>�C<>ȑ>Aϴ��1��d�h��
w��̽0�?}���D�J��1���9������
i�=Tb.?|>���?пe����2H?���d)���+���>u�0?�cW?*�>6��"�T�:>w����j�T`>X+ �Il���)��%Q>\l?��f>&u>�3�Aa8�[�P��~��B|>66?�趾49���u��H��Mݾ�QM>[׾>��C��r�������{i�e�{={:?�?#��߰�f�u�?���0R> !\>4@=(�=DM>��b�wƽQ�G�
�.=k��=<�^>�@?C�&>�n=	��>������[��O�>ƜU>�!>�Z:?�:#?m���ƞ��Ȑ��a-�0y�>X�>�+�>G�>��I��۳=<��>�`h>�jռ����k>1��X>�u�c_a�|(���
�=a��
#�='t�=O��D�<��B4=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ*i�>Ax��Z�������u���#=���>L8H?9V����O�~	>�w
?n?�_�ҩ����ȿ�zv�3��>�?M��?n�m�;A���@�r��>��?�gY?ki>�e۾;[Z�'��>H�@?>R?��>L9���'���?�޶?>��?��H>���?u�s?Qb�>z,x�Z/��2������=��Y;�Y�>}'>�����eF�)ד��i����j���\�a>��$=��>�'佊2��XT�=S܋��@��^of���>)+q><�I>(a�>}� ?Od�>e��>E�=�y���‾��ٵG?�L�?�>��,��&�<�W�*ľL�?��>U��=r��O��>s?C~?���?�>6<9�$����h˿Jžӝw=f/�>oS?s{?��b��>#��/`w��:�=�ϑ>���(���I=�*�=n8�>�8,?��	?��ԽF�!?� ?�lX>q�>�yE����CCE��v�>i�>^T?���?��?�_���g3�ܚ�������X��*S>�Fy?��?}�>�W���Ĝ�$��L���]k�9�?&�h?�r��X?�5�?F�;?k�B?*FU>j:.�P�־�Ľ��u>)�!?���4�A��J&�'��R�?nT?A��>�쒽X:ֽ��׼k���d���?�(\?�?&?���(a�C�¾���<�#�tX����;�A�M�>:e>Z㈽&/�=b>�԰=/Hm�<_6��tf<�=搒>y��=Y?7�d��-?)�i�o7��v��=�8q�ƝD��Iw>c1U>���3�Z?"{7���x��{�����l�V��T�?�<�?���?	���g��<?�Ɇ?��?Z�>�y��#kݾU�۾��x��w��N���=�}�>镰�Ƨ߾���詿K����㲽!}�1�	?r
?ط�><�>��>x�>d˾��.���ﾚ��R�x��� ��z)��%�a�*�߁ʾ���:���現=?3�	ћ>l˼�&�>�'?;P>2u�>�N�>61𼧹i>�~�>.�>���>�J�>�c>zp�=z\4<�Nj�.KR?������'�o��Ȱ���3B?�qd?+0�>�i�;�������?���?s�?/?v>	~h�{,+��m?�=�>3���p
?jQ:=�6�X�<sV����:��]����>xF׽] :��M�8mf��j
?R0? ���̾K;׽�����"��-�?��J?U�@��"8��w��?��_����ؽ�J�|�!�b�4���Y�"���}���;����$�I�:=��V?��?���P�P)��8(��5�!*�>@��>?�;>�[�>�Ù>��&�$7_��[��$�M+�s
?rс?z��>�6Q?�Z9?GaQ?��J?s�>Tѥ>�������>��;��>�<�>�x=?��1?[*6?��?M�?,+>}��k��',Ӿ�h?,�?��?qp
?�� ?Dʕ��Jּ5���V���쁽��<�ȼ�������`=��s>5Y?���q�8�����k>X}7?�y�>���>���H4��h��<a
�>��
?�7�>G���Fur��]�[�>袂?r	�`�=��)>���=IS����ӺpL�=�����=�I����;�h�<8��=���=�2s�)o�`��:#�;���<sp?���>P��<�>�>�6��͜����z�>���> �=��>y\��q��J��|9T�X̲> ,w?8�?�F�>���=y��;D����P�D�ʸ�&}>�V�>+�b?�{?�c�?�O?w¹>��>�N+�#����i���־�.�>w!,?��>�����ʾ��׉3�̝?m[?�<a�����;)�Ґ¾��Խ��>�[/�\/~����=D��������:��0��?뿝?�A�Q�6��x�ڿ���[��p�C?"�>Y�>r�>>�)�w�g�l%��1;>	��>_R?�#�>9�O?l:{?ߧ[?
lT>1�8��/���љ��S3�`�!>�@?D��?��?(y?�{�>C�>z�)��ྊZ������ �݂�W=�
Z>���>K,�>��>��=�ȽDP����>��U�=g�b>H��>��>��>��w>ĝ�<HI?}�>�l��'�s签4ۃ�ϳi��s?��?�M'?iY=#�f�H��<��>��?���?�]0?�OO���=��༏ǲ�U�\�sA�>ܽ�>��>[�=�K=��>�@�>g�>�����23�����IW
?�=A?��=��ſPq�0o��򗾵�e<a��/�d�Lҗ�S�[��1�=�옾֚������[��࠾���%H��y,���h|����>?�=7��=���=�G�<�&żIu�<[�M=aԐ<k!=Xlp���|<��7���»�r�����Y?V<�G=W2��G˾wR}?XI?��*?Z�C?��}>��>�:�AƖ>$
��j�?`$U>�E��\]9�Wէ��^��zؾ,־�c�䎟�%�>{XP�w	>Z3>ƨ�=,��<²�=O�k=c/�=�K�eu=K��=j�="��=?��=.�>Fj>�6w?P�������4Q��Z罀�:?�8�>[|�=��ƾA@?��>>�2�������b��-?���?�T�?Q�?�si��d�>3���㎽�r�=ග��=2>D��=,�2�)��>��J>��� K�����i4�?��@��??�ዿŢϿ�a/>%*9>x�>�R�7�1�� ^��jb�k�Z�G!?E/;�&�˾sm�>�-�=m�߾m^Ǿ�(=�Z6>��n=O����[�P��=��z��q==��m=�͉>~	D>q9�=Z1���޵=GH=���=C�N>g`��m7���+�{8=:��=΅c>��$>Ɠ�>4�?:_0?�Yd?m7�>Tn�vϾ_7��;G�>�=�B�>�=�tB>y��>�7?��D?U�K?d��>hɉ=S�>�>��,���m��l�[ɧ�i��<#��?�Ά?Xϸ> R<�A�ƞ��e>��4Ž�t?Q1?�i?q�>�+
�����>@���?�$r�=GQ�=y4&=�2ܾ޴S=Yy�>��>����m&>���>���>���>ۊ#>���=��V=P�>�;>��=��4�����Ü�<�e�=~�=��=�U�I�<9.P�����%컢Ȼ=a�ɼ7.��9V=㕁����=}��>�5>ޯ�>���=�
��};/>�����L�s��=�F��D*B��3d��K~�/�>H6�ڽB>�CX>�c��D3��h�?m�Y>�t?>@��?�>u?�>����վFP��AJe�]S� �=ٯ>��<��y;��Z`�(�M��wҾ���>-ߎ>��>̺l>�,�x#?�c�w=P��a5���>D}��J��(��9q�@��'���_i�'�Һ��D?pF����=!"~?��I?]�?���>���1�ؾu90>9H���=f�l'q�we��3�?$'?��>����D���C�����=!�A��\g��i����N�y �<��2c�=��ž�r��8 k�(��i*��d�J��f��>0[\?
��?�q�<v ����	6��f<��#?n??f?r�?���>�>?���i�����=��1?h��?&'�?aM�=�߸=q���G<�>D�?���?0�?5	t?��@�%��>Z,��3>����J�=>Tp�=d��=R�?TB	?�V
?�q��}2	��c�i���_Y����<bK�=�I�>�5�>�Sp>��=\xh=Oٜ=ٺZ>���>뙑>Seb>�}�>  �>�����1���??�	>�_�>��,?p�c>�݌������"��g��[��# U���M��3��uzR������	r���1�-?L�Ϳ�b�?�>�����)?Y���i�=��>�Z>�/����>H>lr>	�>�b�>���=�>G=(>4�Ѿ�>����U�!�C��nJ���վ]�r>5���:�'��]�g+��P���E��yh�����[#?��:ZO�?K",�'1k�=) ���"�m}?t��>Z3:?Ns����b�l�'>9i�>���>1� �
���n������Nv�?���?K>c>��>��W? �?��1��3�\vZ�ŭu��(A�`e���`�����,�����
����p�_?��x?qyA?t�<::z>L��?��%��ԏ�3*�>O/��%;�:<=�,�>)��Q�`���Ӿ��þ�9��IF>��o?�%�?iY?�RV��l:����>o�+?&	�>�y?zxc?���?4w��l�>ZJ�WBl>ɩ>��$?H?+�?�H�>�>k�̽7pJ>b׽eR���� ����=�]<.+>�qh����<|5�=��=c�;�$���VY�?���,:����=���=��!>x�>��D?�7�>7��>��3?x���<�^���{?'���S�w��Cr�����B)�� >�F~?�H�?�g?���>B3?��q�/��=^֒>��>�vA>���>6埼���M=93 >v'�=6�)>F����^�Y��3�������<�(>���>o8|>�	��*�'>�v��*3z���d>��Q��̺�z�S�Y�G���1� uv��a�>��K?�?-��=�^龐Z���Hf�0)?]<?�NM?+�?��=��۾��9���J��D���>$��<g��뽢�5#��u�:���:��s>+*���Ҵ���g>1����ӾKk��#D���߾OZ"�!��w�S=
���K�������f�=���=�;�.��K���稿<�B?�= *����a�&���z�=�F�>���>�O��hǳ�O�?�������=T�>@>�3e<Ιݾl�D��o��=�>DQE?7W_?k�?+"��Cs��B�����c���ȼ%�?�w�>�g?tB>|�=b�������d��G���>���>2��)�G��;���0����$����>O9?7�>O�?��R?��
?s�`?�*?UE?Y'�>�������A&?=��?��=<�Խ��T�I 9�F�u��>Q�)?ӸB����>L�?��?*�&?#�Q?��?��>� ��C@�n��>|Y�>h�W�wb����_>ƬJ?蚳>c=Y?�ԃ?��=>=�5��颾֩�;U�=1>l�2?6#?H�?=��>}�>	栾rS�=�H�>�&c?�>�? 
p?���=�?z�1>e��> M�=�ڟ>u��>�?Q+O?J�s?َJ?���>�r�<d��񂵽�q���V�y;W?<�@v=R���'q�S��Gd�<�#�;2Q���)��~��6�C�0������;_�>�s>0����0>��ľ�I��O�@>DB���J��`ي�_�:���=���>��?���>P[#�㯒=*��>sC�>����4(?��?i?%!;ܣb�5�ھL�K�E�>�B?��=J�l�!�����u�Sh=E�m?!�^?��W��'���Nj?`?E?�m���Y��������S��F?^�A?h!���3=c�?<��?w?v9׾kC���玿��U�#��a=�ù>� �<�B�6��>7�?ڌ�>09u>���K��t�YɾӠ ?E*�?��?���?�(L>��f���޿������a?{*	?��ɾ�{	?N������#�ܾsGs�'������S��l�g���|�Y�ܽ6���>1��#>TC+?+5�?��?EF?���6�V���w��\~�F	U������{Q��nP�Q�Y�'����6�ы�M���F !=��d���`����?h6?| c�*��>�"���F����I��>�Ò�F�#�=r�=� ʽ��<�>�]���$�$c����:?hu�>��>�29?Ĥv��D�}0�7��@�eZ2>���>Y�_>W��>�J<���b�+��۾QL����3,v>�wc?�K?�n?1s��*1�������!�a�/�ee��h�B>�\>���>�W�m��9&�l[>���r����v���	���~=��2?�*�>ᯜ>P�?�?�y	��m���lx���1�<��<4�>�i?�A�>��>B�Ͻ[� ����>��l?v��>��>����qZ!���{���ʽ\&�>�>��>��o>6�,��#\��j��V����9��u�=,�h?���A�`�Q�>�R?{�:��G<�|�>7�v���!����	�'�R�>m|?ܖ�=K�;>2�ž�$�}�{��7����?}�?h?��z�#�[��>T ??��?�>�L�?j>�u��]���?b]?��G?1?���>�8<v�6Q꽇�;�CI=ͥ�>�RQ>��X�KS�=���V�������=��e=�W,��]d�v^�<9��<#e�<LeG=1��=�jۿZK��Lپ̧�h�
�i��,/��w凾Db	����C���-�x�����#���U��6c�lŌ��;l�rj�? :�?�C��v݉�쑚��n��|i�����>�r���~��﫾mm�]����3�aF���!��"P��1i�F�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@8�A?r�(�I��r�Y=1��>��	?��?>�1�mw�dj��_=�>|+�?!ۊ?6J=��W�;��Ϯe?�V<F�F�� �\5�=֤=p=�s�ŻJ>� �>� ���@�*ܽoN4>/��>��V��6`^�c��<_�\>zC׽|��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=b9���ǿk8%���
���;*�X�#��{/����y������~!���*���=Ai#> ^>���>yE;>�?_>u�V?�o?���>�9>uｖ$p�K=�Shv�*š�ŧ%�+g��#%[������N�ɔ���
�5I������� =��=b6R�K���� ���b�L�F���.?�u$>��ʾ��M���-<Uoʾ侪�ㄼ�楽�/̾��1�3"n��̟?&�A?5�����V�����k��|����W?�R�ͻ��ꬾz��=庱�~�=�&�>Y��=�⾓ 3�0S��u0?�\?N����q��7&*>�� ��G=��+?��?�F\<���>%M%?ͳ*�v�㽚h[>��3>5��>���>�	>����8۽֊?��T?�����>֐>jc����z� a=�7>�O5��(���[>8u�<Eތ��X������<��d?_>&s1��p/�瘿��?�`d���wr?1_?���>�Ix?��`?$������xl���@�����d?G�z?��=A(=�Ǆ�ɯ�46?8Dq?j�u�v������]|V�&�C� !?l$�?�A?�N�ѵ��dږ�C���?�"�?]VE�\,���_̾7*������s> h�>�C�b�M>�qw?�(�򗮿S�������?��@�G@��������>�(�>�S?���>�ᏽ�&�9��>�k����=gWվ?�؅����!��]?�f?�L ?�eɽ����=�H����?�_�?���L{<�L�J�d�1��g�=\��=E�@������K9��&þ��
�"���� �ř�>!z@ա���>�N�29�P�Ͽm����5̾�Ӂ�9�?�>z.ٽ���n��J|���H���A��Ƀ�ea�>z�>�/��<��{�}o;�\󟼾*�>��6 �>�yS�����읟�yt1<ڒ>C��>#��>xᮽ&���پ�?�g���3ο���a��֠X?-a�?sj�?�?eHA<T~v��?{�s?��<G?�fs?��Y?� &���]�e8�.�j?�_���U`��4��HE�U>�"3?�B�>�-�޲|=�>֊�>�e>$/�t�Ŀmٶ�����L��?ĉ�?ro�k��>/��?s+?�i� 8���Z����*�n�+��<A?�2>������!�50=�CҒ���
?�~0?z��.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?3E�>��?���=M�>ݱ�=Z���6�+�#>B��=�H?�iI?z�M?Iu�>Ѻ�=� 8��/�YqF�YYR��_���C���>��a?ԒL?
b>*ɹ���0�k!��ν��1�I��r~@�>-��R߽��5>�>>.�>۪D��Ӿr�'?�I�ӿ����y늾w	?, >�?j�ྩ�g������i?��">�p,��	��3"����#��ʥ?Oq�?߅?Z�[-�k�x=W8�>��)>1�e=�T�0Fv���G>�k3?��Y�(��C�{���>ٙ�?�@5L�?EZ|�E?���7��?��4���þ|O=�_"?���|/�>U�?�G�=�����'�������>d��?�'�?���>��M?�Kh��)�������Y>�OH?^?噟��Nܾ8х>¥-?:v@�=����ž�rA?���?�@N�w?�s���տ`���a��L����=+���rQ=�X���5=t[�=]�7���ʽ)�>v6�>v3�> �t>W��>B|9>��T>oW��B��ƥ�����C�L�?|	���'��5羱���vq��>R��@�������)T��4����u�ɠl�E�k�� >
�z?v0?`�`?���>���=K�>ʜ���ؼc��M��:��>��B?��x?��[?Ó�����=�N�s̈�����J\����>��=�?3?��>pVx=��`>-H>�
>�њ<=?��S&⽗A�=�>��>]?�C<>�>;ϴ��1��[�h��
w�*̽)�?r���4�J��1��l9�������i�=Gb.?�{>���?пg����2H?
���a)���+�^�>H�0?�cW?Ü>G����T�%:>n��Ӧj��_>�* �l���)�N%Q>Hl?4Ug>�@v>T`3��i8��jP��S���z>�6?寶�)9��v�jH�uܾƨN>M.�>g=J�;��4����\��j��V|=�J:?��?�f���ȱ���t�P����fP>ZLZ>�`=���=[$L>:id�s����1F���*=���=�"\>X?7�+>ڢ�=yݣ>�b���AP�v��>�B>]&,>�@?w)%?������� ����-��w>�U�>`�>�]>>ZJ���=�l�>��a>|L��˃�^��$�?�nyW>��}�r�_�wmu�j�x=3��;��='�=�� �(
=�X�%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>�?�;������u�#�!=�T�>�DH?�j��ےR�.�=�g�
?��?Fw�^����ɿ��v�T��>�?Sє?Nnm�y\��: @����>��?,Y?��g>�ھ�|Z�)e�>��@?��Q?϶><���[&���?���?/b�?7�H>&��?۝s?�g�>jjx��W/��2��8���%�~=�I\;�c�>�>����`gF�\ד��h��{�j�����a>�$=��>a7佚6���I�=����-��Xf����>2q>a�I>�g�>� ?3`�>���>'�=k_��'怾8ʖ�(�I?�C�?���s�^�a����Ͻ�Ⱦ��>x��>?-�:�>*�L�>�`?���?
�g?9�">�<��u����ɿK9Ͼ鞯=ef>�j+?]Ù>᠀�4n�>��������A�<��>*����ܾ6��V1�>��>�&�>�P�>x@!��'?��?��>���>+n�荿m�o��Z?���>��>��n?"�%?u���e4�����ư�V�e�L�>��?#�!?V�>�촿3���q�=(4���OE�,�D?�m?�*<����>�2�?<� ?�r�>��S>Z����بm�e\_>��!?t��A�K:&�3��v�?ƅ?���>�v���[׽�-���������?�\?�&?�h�"a�lþ���<��+���Q��:�;|�A��>w�>�Ƈ��!�=��>݈�=�m��d6���p<�$�=x��>Ev�=F�6�2􏽥�-?��a��}��n�=P�j��FA��ۀ>�VM>O0Ͼ��R?�:���w�Z����S���F���?9a�?��?�K��T�e�9@;?�j�?}�?��>gf����߾ ؾ��i��u�_��1�=)��>S���c��)٢�]㪿z^��<h���ᑾ��>�l�>��>���>4g�=v��>�kᾨ�0��������P�q�/h&�[)/�?�3��U�n@�"����6_�{���\FW�Z(�>�C�+�>Z��>�Y�>���>)�>贱��'>�Ŵ>z9�>K��>O�+>Z��>��>C��=�CW��sR?���v�'�q�꾑(�� B?��b?���>u5[�祄�=����?(��?G��?#Zt>Сh�1+��?���>K.���R
?��A=��ܴ�<�w���7�@���+�ث�>H�ٽ��:�ipM���f�v?�~?lP��.;r���t����|�?�9?o�<���>�R�l�jb�%Yq�A�j<*R�����8M1�
b��ȋ�����7I���y%���=z10?���?3�����c��6�_�k�)�!J�>�q�>��3>M��>�܂>.��~iD�u�|�.]H���Ѿ^�>��A?� �>�N?+�<?>lM?bPL?��>Ik�>�7���>��{;2�>���>�1:?G�.?��1?�^?%?L>�������׾� ?�?=�?�?RP?�>������ּ�19��~��d~���=V=�9�ཬCA�ot=�\>�F?�7�٢8������dk>�7?���>-��>u㏾�H�����<��>�
?�W�>`���~or��Q��/�>)��?��T�=�)>���=ꖄ�|�� ��=�a����=q�����:���<�;�= Y�=�,l�)�<2�:���;�%�<��?�j�>饏�Zs�>]x���/㾽����>5)>�#�=2Nx>�F��ms��W��[�(�/(�>�"�?�˩?�6�>+�='��;��\�?�#�]�E��d��Ľ��?��?0��?��?>O?�?���>Y�<�0ב��x���3;��v	?w!,?��>�����ʾ��։3�Н?f[?�<a����;)�ѐ¾��Խ�>�[/�b/~����AD�>������=��1��?�?+A�T�6��x�ؿ���[��n�C?"�>Y�>��>L�)�o�g�m%��1;>���>bR?�$�>�O?:6{?
�[?�^T>�8��.��Gљ���3�l�!>�@?=��?��?$y?o��>}�>�)�X��e������ڂ��dW=�Z>���>�-�>��>
��=�Ƚ�=����>�ti�=��b>���>V��>��>�w>�կ<��G?+��>���+��n���cz=�v�u?���?�+?2=�r�B
F��u����>Nk�?���?AX*?��S�G��=�ּ�¶�u?q��N�>�ҹ>~"�>�=��E=L&>���>]��>N
��H��J8�O�L���?/F?�ӻ=��ſ2�p���k����"tQ<H�����b������]����=�똾w;�Ǫ�J\�ژ��p��SN��%����]��]��>B��=��=>�=��<��ּ�Q�<]=Kۑ<ɑ	=N	v�t�<Wo6��<������Jxȹ��<�=S=Ӡ��mʾ��{?mUE?�$?�E?v{>�]1>�3���>j�z�U?WZV>Å�����_�/�ұ��M��Ϸվ�t̾�9b�i����>�c��a>�	!>���=���<��=.MS=�=��<e=>��=!�= ��=<�=t�>];>27w?R���'���jQ�t��|�:?�;�>ԉ�="�ƾ��??��>>Q,��V����n��+?���?�Y�?��?Mi��Y�>F���I���8j�=�c��sR2>���=��2�L��>n�J>���&F���ʲ�,)�?R�@6�??�㋿��Ͽ��/>F�7>v"><�R��1���\�v�b��vZ�=�!? G;�G̾�7�>T��=.߾�ƾ�w.=��6>�b=�^��V\���=��z���;=�l=ى>��C>/r�=�)����=��I=���=	�O>�"��֯7�q ,���3=���=8�b>�	&>��>��?na0?bXd?07�>�n��Ͼ�>���H�>��=D�>���=�sB>ď�>N�7?�D?W�K?���>��=��>��>��,�̴m�l徭˧���<}��?�Ά?Ѹ>�Q<�A�0���g>�&3ŽPv?�R1?�k?��>����M�2�L��p\��[�E�<v����_Cr���}��N���:�=�\�>���>�c�>{d�>|�=�'8>�x�>>�=˒��G�>�l�����=�>h	^>z����.��W�=P�1d��c���A�<��;�����Ҽg�;��=���>s;>|��>���=���+D/>Ƹ��_�L��=�G��@,B��4d��I~�/�U6�7�B>u<X>}��"4����?��Y>�l?>���?DAu?4�>��^�վ�Q���De�VS�Xθ=ŵ>!�<��z;��Z`���M��{Ҿ+��>Hߎ>��>��l>�,�=#?�
�w=��,b5��>�|��	���)��9q�"@�������i��Һ̠D?mF�����=�!~?��I?E�?s��>�����ؾW;0>�H����=
�I*q��i����??'??��>����D��¾���%�>��G���N�%����0�J@k��~���O�>��ݻ¾�5�������f�C�ӑ~���>\�L?FP�?�1���ׄ�Q�H�����w��?��Y?b�>;?2��>p-t�tr�㆙���=yQo?��?[T�?�-	>��=v�R:���>L��>!�?1)�?�s?�� |�>fV�Ǆ��%��(!.>��(>ǫ�=MG�=Q?c�>���>��ҽ�����i��^"!�U�=b� >�q�>��>=<>?�>=��`<��=�$R>���>�q�>�f|>�o�>�b>��Ҿk�6�,MG?b��>�Si>C?Ǟa><�3=��2�Z�R=��=�1z�'�C�=�L���&���Y=
f<���<٪�;��7?ۿ��?[��>1�"O-?����>�R�=�H�>���Q�?8�>i>G>��>0��>�]5>*�>Ξ�>LԾ�>8��܅ ��B���R�uо��w>���/(�����O����K�'��������i��T"=�j"�<�1�?k���k�A�(�����?ը�>�f6?���,��� ->Y��>+ӎ>Y���)���x��y�߾CW�?E�?�<c>{�>��W?��?�1��3��uZ�Ȯu��(A��e��`�]፿���Y�
�O��c�_?��x?�yA?R[�<�9z>-��?��%�eӏ��)�>�/�A';��D<=�+�>�)����`�m�Ӿ�þm8��HF>&�o?�$�?�X?�QV���g��?�>,�?
�E>���?�J??�C�?+���ŕ?=1>$r>|�k>|�&?��?�*�>�W�>Q�= ���S�=�zʽh�a���;�������"v��cc�=g^��	�;�(>�{7>�%ݼgn����*eǻq)�=<Z�=���=�&#>]��>�[?
�>���>��8?����=6� E��)?}��<
��kቾ�쥾\���r>GWl?��?њ\?�#i>�vA�A�?�^�>�4�>�m*>^>e�>>�߽P�<�*�=��>�x>��=9�[��倾t	�Nk���.<~�,>4��>2|>���)�'>�z���-z��d>��Q��˺���S���G���1�2�v��Z�>A�K?j�?���=6_��2���Hf��/)?�]<?�NM?�?�=��۾��9���J�=���>�[�<��������#��?�:���:��s>�0��|���eb> ���>޾�n���I����"K=_h���U=�8��T־�����=�
>���>� ���ͪ�0,J?�vl=7"����T��=��$>��>�Ԯ>]�:�=�w��@�~���?��=���>��:>&������~�G�:�w>�>YQE?/W_?k�?�!��:s�<�B�7����c���ȼ$�?lx�>0h?LB>���=7�������d��G�q�>���>B��(�G��;���0��%�$�ꊊ>@9?ة>��??�R?r�
?��`?�*?2E?'�>`�������A&?5��?��=��Խ��T�z 9�KF����>l�)?9�B�Ĺ�>Q�?�?��&?�Q?�?c�>�� ��C@����>�Y�>��W��b��7�_>��J?Ԛ�>h=Y?�ԃ?h�=>R�5��颾�֩�#V�=�>��2? 6#?P�?쯸>���>�����=���>hc?1�?��o?)z�=6�?�02>W��>3�=t��>_��>�?�WO?��s?��J?��>#��<�B��^6���>s���O���;�CH<��y=����9t��H�G��<x�;�g��'��٘�@�D�V"��ͽ�;cc�>��s>���P�0>��ľCX����@>���J���ኾ�}:����=j}�>�?✕>h[#����=)��>�R�>&���5(?��?	?�\";I�b���ھ2�K��>VB?���=:�l�������u��5h=��m?8�^?ѓW�[ ��/a?IA?���� �o�����S�=?�Ҿ�@?t�>z$H�Vc>��?�4�?���>p��H������	[�]O1��FM=WP�>�{׾�0/�G��>�]?_L�>N��>�xJ���}���}�v��c�>�N�?��?�.�?RuJ>z�Sܿ��5���D?*��>�����e ?\҈=f$��>W��b��/�	�d8��8�̾'׌������5��	������x=��?��?pJ?�fb?��̾�A��H��ml�^$C��*
����JG�.L��8�tp�1�8B��{����	�;�����[�/��?b8?�
 ����>pة�L�ʾ����W)�>򺷾����kv�=m���a�J6�=������Z�U��D�E?��V>1=�>GE?�Oi���Q�H�F��9پ��o><�?[��>Ra�>�����y�ݽP���F��=�7v>�xc?B�K?y�n?�o��*1������!���/��c��+�B>�j>w��>�W�u��9:&�gY>�1�r����9w���	�a�~=x�2?s(�>!��>�O�?�?�{	�8k��Skx�#�1�O��<�1�>n i?�@�>�>�н�� �3��>R�l?��>,�>.���!Y!���{���ʽ}(�>ح>���>A�o>��,�$\��h��&���9��w�=~�h?p�����`��>�R?��:\:H<rx�>��v��!�����'���>?,��=w�;>�}ž+&��{��/��qF)?�Q?�Ԓ�x�*��\~>�+"?���>Z �>2,�?z�>�kþ|�^��?��^?�CJ?�RA?�H�> =U��5KȽ��&�ݬ,=d��>!�Z>X�l=ZV�=U���t\��z���D=�G�=��ϼ�H��\<�����GK<���<N�3>ojۿ�4K���پ���*�]-
������׳��A��%�������`��ԏx����&��V�Z:c�r��L�l��{�?�;�?�4������{���Ԁ��?���š�>�fq��d��L���R�0j���ྱڬ�'m!���O�Ai��e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���y¤<���?0�@!�A?�d(��M쾣�d=D��>��?��:>�r,��{��:�����>��?A�?�<=B�V�0K���d?Wz<
�D��ѻ���=B\�=Rq =&���I>g�>Z�p�B��	ܽ��7>%	�> &�n�Ҝ`��;�<�W>��ҽ�V��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=ʸ���ƺ�w?.�~���I[<P��;�
�<dw��5l޼��t<�6��) ��-���bx=��=h�^>�f>��|>\f3>�sR?�w?��>�pU>k�Ӽ��4�-6���/弸+`�W�l��s���{���eﾚ����꾬E��A�/a� �˾� =���=�6R�.���� �Y�b�=�F���.?wx$>#�ʾ@�M���-<�pʾ�����܄�ॽ�-̾��1��!n�?͟?t�A?�����V�����W������W?Q�����鬾:��=3���-�=$�>��=��⾎ 3��~S�61?E?M#��'��NX4>�e��0�<��,?��?':�;��>�p%?��.�`p��W [>�7>�U�>Q�>��>����2�ؽ�?(�O?�	�q嚾��>�����{��"[=�S>(0�6Q{��B`>U�_<u���9�n+���J]<� ]?c��=�!������n��!��s½T?�*�>uEf>1�l?s'?�������;]I�8�)����=PDR?�S]?���=z��=Ԕ��j1���=?g�?��E��_�� �MD�@P����>���?�D?��>�l��T���C-��<?N�q?�\�W"���	#������Ƽ��?�9�>����c?vn]?�8������
A��_G����?��@�A�?ܿ/=�w�$Cv�NX�>}\�>�&�M?|�\ 5�_��-�>��3?my�I0������>��?�,?��>�|ټ�����=Kڕ��Z�?o�?�����@g<���pl�1o�����<Ы=$��C"����7���ƾ��
�����*޿�{��>4Z@_Y轂)�>�D8�n6�TϿ����[о5Tq���?��>#�Ƚě��h�j��Pu�O�G���H�餌�qT�>��>����1쑾�{��q;������>���t�>��S�J������4<[�>`��> ��>v���׽�:?/_���:ο����_���X?|i�?�j�?�g?&u9<"�v��{��	��/G?|s?�Z?q&�~.]��e8�=�j?�j���M`�N�4�yXE�s4T>�
3?Bo�>�|-���z=�>3��>��>�0/�G�Ŀ�ζ�9����?���?�K�d��>�`�?^e+?&q�0���ȩ�S�*�>��>*A?�
2>�)���!��S=�����;�
?Ǳ0?�-�+�]�_?*�a�N�p���-�}�ƽ�ۡ>�0��e\�N�����Xe����@y����?M^�?i�?ѵ�� #�h6%?�>c����8Ǿ��<���>�(�>*N>[H_���u>����:�	i	>���?�~�?Rj?���� ����U>�}?	�>"�?�y�=�~�>M�=]ʰ���0���#>��=g�C�j?Y�M?֓�>���=7�7��/��SF�A
R� '��C�>B�>M�a?�YL?�b>�[��r.�,!���̽h
1�\q�I@��r,�!޽�B4>6�=>,�>��D��Ҿ� ?����Կ�����J��!?��y>(L?xB�������=�b?�k>3d����z���&�?Q�?�?��̾�r��&>|�>��n>�
�<1��`{���3>�>?�Ͼ�����*x�r��>з�?�@��?��e�k%?�Z��:��W�r��'����^PK>e&@?��۾�>��?��>��|�48��*���)��>�̪?���?w� ?=�S?<fU�c34�=�b>S�X?ޤ)?����]��v�>���>:X��O_������Uw?o@�%@u?#욿nFԿ.����2f����V-\��Q�>������>Ռ=F�<�`�<�i��@>%9n>���>j�>+	G>ce>��}�9��X\������6l��)�S��#�緉�.�Ž[��ʾ��Tݾ��5�х	���Խ�D���۽K��T��=CN�?(�M?��X?��?i��<2{�=�2��?t�������Zy��9;>e�@?�S�?��M?<������8���p�)ҿ��4�����>Nq>d��>7$�>�5�>Cl.��'�>b-�>�ߖ>l�=�q=�?=�w�|�>e�>��>)��>�C<>��>Dϴ��1��g�h��
w��̽0�?����T�J��1���9��˦���h�=Jb.?|>���?пg����2H?!���x)��+���>x�0?�cW?�>����T�5:>B����j�;`>�+ �|l���)��%Q>ul?7�f>	vu>%�3�yK8���P�r`����{>t86?�"��H�9���u�3�H��
ݾ�M>�>��?��k������&�h�i��y|=�f:?m�?��Oﰾ��u��P��DR>i\>l�=�L�=�<M>b�`�t~ƽ�VH��?/=�3�=��^>�y?q�*>���=v��>�g��uVQ���>S�B>�,>�+@?�G%?�h�J$��G�����.���v>(��>ź>n>#�I�ᥰ=�$�>�a>����΂��j���>��mW>	;���_�	�t��'}=�T��BN�=`̒=�����=��&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿl�>#��X��;��S�u� K#=���>�:H?R���P�t�=�y
?�?�b�^�����ȿ�zv�D��>E�?��?��m�hB���@�>x�>D��?�lY?,ei>X]۾�eZ�v��>�@?� R?�
�>G8�Az'���?�ܶ?B��?jI>���?�s?�k�>�0x��Z/��6������p=��[;�d�>�W>^���wgF��ד��h��v�j������a>��$=,�>DE�\4��z9�=��I���f�7��>�,q>�I>!W�>x� ?�a�>���>�x=�n��Nှ������C?�t�?�eξ��O����=ί>Y�Ǿ��?�ҁ>��[�������>�c?q�o?t?t�>� ����J�ǿJ�����=A >�}?�o�>������{=[ݭ��,�D�=�'y>�y<�����Ҳ���>Ҿ�>��"?��>S��;"�#?�w?��l>�z>��J�����μV��}�>��>o^�>��?i?�о���3��i������\��H>��~?Y@?���>�S������=��D��b�=E�n?E�~?��{�X�?��?�?��?���=�|罝G����G��2�>\�!?����A��V&�q����?8?��>(��O�սTټ����9��?o,\?�>&?����=a��/þ|u�<4$!���V���<!\B��=>M;>u��bF�=s�>�5�=3<m��W6���h<�=���>O|�=�k7�������.?��c��0���{�<��v�b{J�Lu�>PVE>�)��әk?нݽ�6v�� ����k��:̅?�:�?`��?t7����]���;?cH�?��?���>朾���v:ɾyH]����>�I��=ie�>�bO<��۾�➿�p���م���r��Gc��� ? m�>�?��?��}>��>jlǾ̛����q�{��y%�Cc,�>'�S� ��u��h>�-������H*��N�>��{�T�>�0?m(\>�ii>9μ>D.��LC>#�>���> �>h^>�\>2$�=�q��͆�LR?(�����'����!����5B?�ld?U3�>DLi����-���?Ć�?�q�?�Cv>H~h��/+�	h?6�>I���p
?$[:=8���^�<YX�����@���1�/��>�a׽�:�JM��Yf��m
?.5?�Í��̾�q׽8�g�����m�?l�?�E-�0�D�K���sS��o�ll�=���;�*��h��(����x��;���8��Q�=��H??9���b�־`(��J�=���>�5 ?�]�=��?A�>��Ac0���r�mk7�;���D�>��?{�>ؙJ?�;?4P?��L?�Ӑ>��>0𮾨��>i"��A?�>rJ�>*:?��/?��0?�m?:*?��]>�������ֈ׾�?��?�?�� ?�??t臾�1½X發�`��Tz��߆����=Q��<�0Ͻ�p�b�G=�&T>@�?e�m28�'c���[j>��7?!��>���>x��������2�<��>�2?�p�>���Z�s��:����>���?K���Q=X�)>#��=yb���F;���=/�ü�ō=�q�/�G��BJ< l�=RȘ=Y� �a7(:<ҫ9�c�:_��<R7?��?%�>��>hZc����o���
>;�>y�;>E�(>�+���؆�p2���^\���>�݊?-��?�h�=�=�=����8=��G�sW��Ň�=��>"?8�J?`Q�?߇7?��(?QJ2>���cٕ�劉��H��C#�>t!,?��>�����ʾ��ω3�̝?j[?�<a�6���;)�ِ¾��Խ��>�[/�`/~����<D�����'��1��?꿝?8A�R�6��x�ٿ���[��v�C?"�>Y�>��>>�)�x�g�v%��1;>��>pR?�"�>$�O?�:{?$�[?,mT>�8��/���Й�Q_4�,�!>@?U��?��?1y?�z�>h�>��)����U��/��b���ق��W=(Z>͑�>m+�>*�>s��=_�ǽ�K��)�>��a�=_�b>���>ܜ�>���>��w>���<}H?$�>�!��M\����� ��M�J�!�u?���?��*?=����E���� �>�4�?O��?,*?�O���=s�ټ!ɵ�0�t�;��>:�>$��>`
�=��C=78>Y�>��>S����Κ8�ߔV�?�?�E?]��=Gƿ��m�b����ꔾ�:����'Q�I���I7����=��UH2�cG���R�f��Ts��{մ�2ݑ�j�z�p-�>�6�=�>�m�=��(=�.����<Ӯ<=O/,�-��<\6����ͺt�0��N˻�����p�Í;M��<��D�w�˾��}?�:I?�+?>�C?��y>\W>g�3�ٙ�>㏂�=?�V>P�;q���j;�ʩ��S���ؾ�y׾D�c��ʟ��;>�HI���>�D3>�k�=J]�<�-�=V�r=Rώ=�TS��=\�=[B�=�h�=/��=�>`>�6w?6�������c4Q�#X�P�:?�7�>�{�=�ƾ�@?��>>�2�������b��-?B��?�T�?.�?�qi��d�>���㎽w�=�����>2>���=��2����>��J>����J���}��24�?��@��??�ዿâϿ�c/>ݴ7>�*>��R�̇1�@�\���b���Z���!?wJ;��K̾81�>n�=�%߾|�ƾ@�.=�6>Vb=�q�xX\��ә=��z�0�;=�2l=N؉>;�C>tq�=�9��+�=ҝI=���=k�O>�땻cw7�u),��3=���=��b>�&>���>��?�0?�d?/�>-Hn��ϾQ,����>p��=�ݰ>���=��A>h��>U�7?�D?�K?_r�>���=_ٺ>V��>/,���m���g맾���<l~�?���?'��>}h<�&@��B�_	>���ƽ�?��0?o?-��>���Iƿ��`�Y%#�5O���d��c�>U��w�>r�>���e^�Ak�=���>���>��> _+>��%>R>�Y�>X)>kʮ=�>t��=wZ>I�#<��(<:�q��0�J-��M��-e=dND�?���0�a�1�&B'��Ko��:�=���>B�>���>B�=�ݳ�2/>\喾R�L��,�=�~���HB�Bd��5~�8�.�7n6��B>&jX>o��o����?�[Z>� @>\��?W@u?ӎ>���ґվ�M��-�e�BS�y�=P�>º<��o;�P`���M�D<Ҿ���>Jݎ>� �>v�l>�	,��"?�?�w=���_5���>�y��ζ� 1��9q�_?������Ni�J�кۢD?qE�����=& ~?гI?��?Q��>9+���ؾ�?0>;M��a�=!��q��t��t?m'?���>�쾯�D�B4��NJ���>�e���T�>;��.�.���;=��c�>�ǃ�,g���`5�	=��O����5D��cy��-�>[�S?%�?=�D�J{��%�F�&����̽��?��X?�̪>��>J�?΁P�]������=ZNt?�>�?�B�?C�=d��=eX���B�>�0	?���?���?��s?z?��r�>0��;� >�������=>�	�=�q�=p?�t
?��
?�����	�+����(^����<��=X�>CX�>�xr>\��=�g=��==$\>:۞>��>��d>��>i:�>[aо�(��;H?M�>���>��>?  �>�1���؊���G=�������[@ӽ�O;�l?�ѳ�<�J���漌���7?�ݿ˦�?ύ>�g�h*�>ۍ�ω�>H��p��>%2�;QҦ>��n>t�=��c>���>a��=�j>�N>�:Ӿ:<>4���Y!�+C�T|R���Ѿ�z>�����%�ݕ�����t-I�ys��o�3j��-��@8=���<NK�?����z�k� �)�I���{?RD�>A 6?Ԍ�v3��~>��>��>�S��ݑ��QǍ��h���?D��?�Wc>��>��W?��?1R1��3�_�Z���u�$A��e�ϵ`��ۍ�˛���
�;���!�_?�x?rA?�3�<�,z>���?�%����~L�>�/�+);���<=%7�>�)���a�[�Ӿ��þ7H��F>�o?u�?RK?ZV�M��Y�?37?/%?σ?�d?ưY?V�4����>�P��>��>n<?�"Z?��"?vV>�t2>j�N���3��$m��s���?6�Bּ�<e��=�޽��V=��l���=7�2�% �@�f���<=�=@��=����>�)�>��0?P�>a�?�d?.\1��r�s���UD?p1���"��f7.��Z��x���,1>`?���?��4?�!?�F��&� >���>�T�=Yw>f�>�\�=�ꝼO��=I��=R�>mL>�����Խ�־rӾ�R%=R�_=���>N7|>�	����'>�x��B/z��d>=�Q��Ϻ�&�S�-�G�>�1��{v��\�>��K??�?��=�_�V>���Hf��/)?�]<?5NM?{�?H	�=T�۾^�9���J��:�
�>�3�<��ƽ���"��E�:��ޜ:H�s>;,��^M��yb>>���ݾ6Sn�z�I�n��!�G=â�*PM=����־�(��$A�=�1	>_���
!���������&J?�co=jC��<2U�a��39>mE�>]��>k�<��Pw�U@�Ĭ��=ʰ�>Rq9>�ۣ����*�G����k>�>SQE?@W_?k�?"��Ys�>�B�����mc���ȼF�?ix�>&h?�B>|��=L�������d��G���>���>f��I�G��;���0��K�$���>U9?�>��?]�R?�
?{�`?�*?HE?&'�>'�������A&?V��?��=��Խ��T� 9�"F� �>I�)?��B�q��>��?!�?�&?C�Q?��?��>ޭ ��C@��>�Y�>�W�]b����_>j�J?��>�<Y?�ԃ?��=>Ą5�颾4٩�GV�=�>�2?�5#?Y�?!��>��>󫡾��=U��>�c?�0�?%�o?B��=��?z;2>���>��=���>ً�>�?�WO?�s?��J?<��>��<�9���4���6s��O�ɜ�;�qH<~�y=x���-t�=J����<{�;Ra��C�������D���-��;�_�> �s>�
����0>��ľ_N���@>�x��bO���ي��:���=���>��?e��>Y#�Ŵ�=׭�>PH�>1��`6(?��??o!;��b���ھ�K�v�>Q	B?���=��l�Q���v�u�/h=��m?%�^?=�W��&���g?I�D?*��Hw���Y�*����P?4�?Zl��&
}=[G�?���?��?�q,��)��Y��¢y��ͻ,&����>f{ھ��R�X�>�"V?W�>�>��-������S�&e��]��>��?�#�?��w?Ņ=>�<�kݿ����{��e��?Z�?aڥ�_?����q��U�׾T���,(¾���:ᇾ��P�깾�2�ع��N����>ÄC?��u?�RO?	1?$�	�dD��4���Q�]	q������zU���F��b��6j� Q>�Q��^Ѿ�q�=��y���N�5ļ?��&?G��p �>����������F#K>Ϣ���J���=%ۧ��G:��B=�ꍾ<>����B�5?[�>P�>{�3?�o�p�?���6���0����P�S>�}�>��Q>�
�>f	[�c�Z��T���r;Ҡx��?�:4v>Ryc?E�K?A�n?�h��(1�������!�s�/�5e��d�B>�i>��>b�W����";&�	Y>�V�r���� w���	�J�~=F�2?
+�>��>�O�?�?�z	��j���mx��1�Z��<�0�>�i?b?�>��>�н� �ĸ�>��l?��>Y�>����iZ!���{�0�ʽo&�>�>Ӷ�>��o>��,��#\��j��T����9��t�==�h?�����`�H�>5R?�<�:�G<q|�>�v�ӻ!����X�'��>�|?��=8�;>n�ž%���{�g7��vn&?��?������*�b�>��"?qq�>���>ن�?�<�>G����z<�_?P._?<PK?��<?D?�>H=�<�ʽ׽�E#�jVT=���>�`[>���=q�=��'��JV������H='��=���T ��S{�:n�ռ-3�<�R�<f5>maۿ&K���ؾ`��
�
�I��,���Ib����	�v,��4���-x����Gy'��V��Gc�������j��n�?3-�?��"�����aw���6����>7�r�� ��꫾A������xA�٬���!�<P��Ji�Ԫe�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >jC�<-����뾭����οB�����^?���>��/��o��>ޥ�>�X>�Hq>����螾f1�<��?7�-?��>Ďr�1�ɿc���t¤<���?0�@Y}A?��(���V=���>��	?p�?>�P1�WI�m����T�>�;�?���?CjM=�W���	���e?.�<��F���ݻl�=&9�=M=r����J>�V�>�~�RA��7ܽ��4>
څ>�o"�A����^�&|�<[�]>q�ս�9��5Մ?,{\��f���/��T��U>��T?�*�>R:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=u6�����{���&V�}��=[��>c�>,������O��I��U��=Q��muſ�M!�ڴ� �<{���l������⠽e���L���o��u��n�=C��= zU>b&�>��U>aj>W?U4l?��>��>T���!��f�˾M~��I_��Y��S�);!��
����N�߾�_�e�����þQ =�_�=7R�L���Y� �u�b��F���.?w$>��ʾ/�M��-<�pʾ����W愼zॽ-̾i�1��!n�-͟?-�A?����|�V�L���Z�����w�W?4M�G���鬾���=������=$�>\��=���� 3�J~S��?0?��?lD��Z�����*>� �Qm= �+?�i?nR<�Ȫ>��%?H)��$�]>�73>kZ�>�+�>��>RI��T�ٽܠ?�
T?�^�>��A��>⾾/`z�eA_=a>,P4�����"%[>�.�<�)���UL�9Џ�,T�<�F^?��7>z3>�_+�"&���_+� |����b?G�?٬�>��E?�&?|��=�^微�R�Z���n���?ds?L�>�/��N�����8,?C��?1��5�h�n�~�<�b@&��M?�Џ?<U�>����p�������S�%�2?#�q?��d�A�1�����7�ɽ���\?ԏ@?�"��8�p?��?�Ͼ�������3[a����?�L�?Av�?R���E��κ=��>q�>�	�=��ѽ��ռqD{���q��uh><Z<���`Aվ1�1��|-?�Z?��>�fG���ؾ���=�ؕ��Z�?��?����\6g<8���l�r��-��<"ȫ=FI�rc"����<�7���ƾ��
�
����w��֪�>�Y@xQ��&�>�98��2⿃PϿU��E_о=Xq�$�?�y�>��Ƚ������j��Su��G��H�����eܣ>�>{ޗ��|����{�χ;� u��A��>�����>qS�����ߥ����<��>���>�k�>Tܩ�^�����?�0��3ο�z��X����W?G��?���?��?,r<4�s�zz�:T� G?�s?��Y?��"��]���6���j?�����o`�r�4��uE��S>�63?fx�>l-�j&�=2�>O^�>1t>9:/�7�Ŀޜ��	��\��?'s�?0[�Ur�>t�?��+?nm�8��S6���/*�������A?74>���J!��<��В���
?Bw0?����%�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�$N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?ǖ�>���?m�=��>��
>�~���C3;��8>���=/���p��>3�R?��>�}�=���dA+�m�@�P�M�I����A���>pNb?�@A?Ŵn>2\P�Õ!��T)��
Ͻ�/��r���?��֔��J׽�8>^� >�.>P	O���ƾ��?Mp�9�ؿ j��.p'��54?1��>�?��w�t�W���;_?Iz�>�6� ,���%���B�`��?�G�?<�?��׾�R̼�>6�>�I�>�Խp���W�����7>5�B?\��D��q�o�v�>���?	�@�ծ?hi��Z
?ܞ��ԇ�d}����jA���=��6?��?�~>l�>S�=sDw�}ު��t����>s�?���?��>a%j?�fm��LB�`,=��>�Ce?r?I��<�R���N>FV?��h��� �_bd?@
@K�@ �]?q����ٿ�?��X���I!Y��ҝ=_vP<��=�8p��SU>��=�(��2�=G� >���>`l>�Ug>��">��#>I'.>N����@�=��1x|�DH�����H4��ۇ��!��Tl�AO	��h����P�Z�ӱ��C8��J+�bc�� A�<���=�vz?�>?��*?�?K��=9SB>X��}^�=�X�=�K�uɳ> C4?S�X?�:.?�,�D����W��w��X��cQ���C�>kH>>��>���>�>�>�K��΃M>%�>A8>��<��=��r=����&��=dM�>���>5��>�C<>��>Eϴ��1��g�h��
w��̽1�?����Q�J��1���9��Ʀ���h�=Lb.?|>���?пf����2H? ���w)�ڹ+���>x�0?�cW?�>"����T�/:><����j�$`>�+ �kl���)��%Q>pl?��f>YRu>#�3�@e8���P�'[����{>�76?�ﶾ"Z9� �u���H��2ݾtYM>n�>�vE��q��������i�6�{=qs:?��?6�����-�u�=��~aR>�%\>R�=$Y�=%@M>��c�x�ƽ��G���.=���=�^>Vq?3E+>P�=ٙ�>����kiQ��٩>�)C>�1,>�<@?�U%?�������r���?_.�]�w>ϊ�>�[�>�_>�MJ���=f�>)�`>�c��.��ܠ��O?��W>}���^�|t���{=H���!�={ڒ=/����=��h$=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾMj�>>x�zZ�����f�u�n�#=<��>g8H?�Q���O�,>�%x
??d_�s�����ȿ�|v����>w�?���?��m��@��6@�ƃ�>���?�dY?Roi>�e۾�gZ�l��>�@?�
R?��>8���'���?�ܶ?���?�I>t��?1�s?�l�>,x��Y/�76������c=�YZ;md�>%S>����jgF��ד��h��x�j�%��{�a>��$=��>�D佝3���@�=�苽�F��S�f�ޥ�>)-q>Y�I>W�>�� ?�`�>���><{=�j���ှn����3?bn�?��m�d�0�=�S�>f���|/?�O�>{�ֽ܍�jZ�>WW?��i?�0�?5|�="'�����b¿q��}.4>�i�>`�?�Q�>A�j���{>�����ϧ���/>��>�9�<_mھ�ҕ����<+��>EL?L�>Q�ۼ�� ?O`#?i i>'±>�\E��9��Y�E�C��>/��>d?��~?�?�����-3�����6á�nW[�%GN>��x?k*?�S�>�U��򬝿�L�U�G� 㒽s��?�g?��㽠�?%0�?��??V�A?�Nd>���6�ؾ���7À>��!?��t�A��N&�t��b�?�Q?~��>K����ս_uּ����o���?�'\?�;&?����*a�y�¾,��<�9#��1U��2�;��D�l�>��>�������=>���=�;m��U6��e<cb�=���>��=�&7�zd���8?n	q��X��U�H>�\=�[1�W6�>�\>�t�d�2?pj�ML�m��@���Sf��u�?n�?���?!�ǽ��J�m=??�D?�4?�[�>9��a����f���;�;�15�v�=�<�>E����v�D
��:C����t���<����M/�>9��>�!?��?R�>B��>�ܾ�9/��a��Ik���1��C5�I�9�6�;����a_���oH� 9��B4���M�>�?A�RS�>w?R��>37�>Z�>5\�=��L>`ɉ>��>"S�>s�>8Ó>��^>�h�=M����^R?�#��=�'�ޮ쾧����B?�2b?}��>C�j�����?i�K�?��?*��?)z>��h�|�+��b?���>�(��+�
?��<=�ʻy�<���6;���X�0����>��ؽU�9��)M���d�F?~�?�_��p˾�|뽟���Ʉ<���?e3?�� �g�:���c�mI[��fh����3�s�}��7$�@ce�W��r������Ȍ,�7��=�7?J��?.+��X�
v����E�n�(�T>��> ?P>��>�Z>�"��tD���_�/+�����־>'�B?���>�\?��8?P�3?�O?0�>�(�>-����q�>����S�>��>?�5?U03?�3?1?�?�6">�Z2�R� ��վ$�?�1?��?A�>6��>���������۳������D����=>�[�
���p�+4p<Q?X>�W?����8�c���!k>9�7?ـ�>=��>���-�����<5�>Ŷ
?�J�>����5}r�)c��R�>W��?���x=b�)>���=����Ӻ�]�=������=����f;�2�<;y�=0�=BXt��r��X�:���;=|�<w�?��>Tq�4�e>�ַ�W��Q��%(�=�70=�";>(�=-�Ѿrh��c��}�7����>xQ�?�Ȯ?_��>���=}��cؾY�	�VI/��$��i�>�X7?�d?Z��?�͘?�^?6ZF?0V�>�_2�Ĉz�.���߬�c?w!,?��>�����ʾ��Չ3�ڝ?i[?�<a����;)�ސ¾��Խұ>�[/�h/~����>D�>���U��6��?�?KA�W�6��x�ڿ���[��{�C?"�>Y�>��>U�)�~�g�r%��1;>���>kR?`#�>��O?l<{?�[?�iT>��8�1��fә�s:3���!>�@?���?��?�y?�t�>��>6�)���T�����H�����W=�
Z>B��>�(�>��>i��=�Ƚ{\��e�>��a�=��b>��>���>�>��w>�Q�<�H?x�>3c����� �Ⱦ�q�<�O{?���?�:?��>�B��0D�����>I�?N_�? �0?a�i����=���α���u�)٥>D�>�R�>�=�<�<��>f�>�E�>o%��g��5�K"v���?%�<?Gɇ=h˿7�r�sw	��>�=�Խ��e�T���v��F�=,�׽��4�A��<�����ؖ������i̽l���n�������>��=c>��=���q�;���A`Z=/t(�d�������h�q�
^û{o�=?@������=��,<��g=G;ʾ�~?�H?p�'?�HF?)�>��!>��%���>�M��5?�-X>a�)����82�9���͉����پױ׾�f�r����>o�.�˴>ɂ5>���=��@<�M�=�~=�ҏ=	�Q��=��=p��=�5�=��=<�>�i>�6w?���������-Q��a�{�:?�@�>y��=U�ƾ�@?��>>�0�� ���Ye�](?���?�V�?��?�ti��a�>��׎�Q��=�>���d2>���=�2�揹>��J>��WC��'���2�?�@ڙ??�݋�X�Ͽ�l/>ͭ7>�Z>��R��1�҃\���b�pZ��!??@;�G̾D1�>jS�=�߾�}ƾ4/=��6>�1b=cm�%W\����=$�z��L<=��k=>։>|�C>�ʺ=:|��l�=W�I=���=��O>����.�7��\,��x3=���=u�b>�&> ��>�?a_0?ETd?0�>�n��!Ͼ@���C�>� �=
A�>"߅=�^B>���>V�7?~�D?��K?A��>�É=

�>�>�,�F�m��m�ҧ��Ҭ<���?�φ?�Ҹ>eDR<O}A���Hg>��Ž�w?�T1?Kn?�ߞ>ڥ	���ο����r�ݽr
��p
��o��p�n>?���j����\O>�%�=�4�>���>���>�,4>�lC>jE�>�L�>���=�0=���=Y ��+ҕ=J�@�x�^�]吽b�����=_/i;[Os��!��fޙ<��=*8�;�~=��u=���=:��>�U>���>Ď�=K��6/>����L�&[�=/F���0B��6d�3F~��/��}6�G�B>�X>at��V.����?}�Y>5i?>G��?$Cu?Y  >����վeN��EBe��\S�k��=H�>�=�P};��V`���M���Ҿ���>Zߎ>��>��l>�,�#?���w=�sb5�)�>�|������*��9q�@�����ui�eӺ��D?]F�����=("~?ưI?k�?j��>���y�ؾ�:0>�H����=\��+q��k��[�?�'?���>T�)�D�>DP���J�i�>k�:���P��ˁ���C�.u�f����\>afž�}�}�?�L׌��>���|#����̰�>�GV?�w�?�_)����"@t���i�]�O˴><5V?�
?/��>5v�>/h>�A1�8=־[ZI>��f?���?���?�\D<�=Nz�����>�?���?�ӑ?Vos?��=�%��>�#4;��>�n��z(�=9>�_�=ɐ�=�Z?�i	?��	?�W����	��G�]���^�f��<�=�>��>T�s>Y��=9+l=��=u~Y>�d�>�>| d>gã>i�>^�����rK?��n>1�>5?�@�> ��v�g��Z�Q����%�a�,`���U��B�������b��G�a{&?Ʋ�'�?���=_����>A�1�S>R�=n(�>W'��q��>I��>?Rw>��>�k�>�{�ǫ>n�>�FӾ >����d!��,C�D�R�u�Ѿk}z>�����	&����w��1BI��n��~g��j�L.��S<=��̽</H�?`�����k�*�)�Z���D�?�[�>�6?�ڌ�=����>���>ȍ>�J��`���Pȍ�(hᾌ�?7��?<�l>��>˃U??�~:�m5�1\���t��zB�Je�*&`��،��g���D��T۽�z]?�x?�C?�'�<뢀>��?��,��<��VW�>o�0�H[8��]�=�β>犱�4Y��"þ�|̾�(%�I�Q>��o?x?3�?�7_�ʜ#�C�>��"?�Z�> ڐ?��]?�H?κɽ�E9?C۱=��b>�ݰ>{�(?u�V?�4?g����Bѽ�+R��7�/�s���C мrL==飽�8 �3٥=��)�Ø>�3�=~P�=�؃�P]���� =��=�]=$�<:�>�/&>�ئ>�]?t�>-��>��7?���Nb8�ñ��]�.?��8=u����������*$�<>`k?��?�wZ?�=d>l�A� �B��>؄�>�d&>��[>�$�>�
�q�E��D�=��>�>�ۥ=�^M�������	�ǽ��u�<�Z>���>2|>����'>|���/z�V�d>1�Q�T̺�
�S�p�G�^�1��v��Y�>\�K?w�??��=@_��.��\If�0)?�]<?�NM?��?�=�۾��9���J��>���>dW�<��������#����:�Z�:��s>�1���{���8>T&����ɾb	d�I�B�%V۾��<����8�<2 ���꾸���1��=�	>����#�"����������L?3��=�d��H�7�3X��%>?��>ƍ�>��B� V�"�9�;?���M=TX�>�G*>��;>��E(N�t	��=�>oQE?vW_?k�?�!��s���B�����Yc��rȼ��?/w�>�g?XB>%��=(�������d��G��>T��>�����G�H;��0���$�/��>�9?}�>c�?F�R?��
?�`?�*?SE?�&�>���0��� B&?6��?��=��Խ�T�� 9�KF����>{�)?�B�׹�>P�?�? �&?�Q?�?�>�� ��C@����>�Y�>��W��b��?�_>��J?ך�>s=Y?�ԃ?v�=>[�5��颾�֩��U�=�>��2?6#?N�?�>2��>�����=Þ�>�c?�0�?��o?<�=��?*92>���>���=��>��>.?XO?��s?�J?̏�>M��<�9���8���Es���O���;�|H<��y=֒��.t�CI�l��<"�;�l���M��+��Q�D�s������;�4�>��o>3����7>�d���6��j�2>�6���r���֏�=nC�x��=;:t>��>��>��z�=o��>-}�>E��$?.�?�k?��;��`�Ȯپ�E�#�>�&@?���=z	j�����\�u��=K�m?d#a?�T�N
��a�`?JI?N��N^����KJ<1���h?b�?����>�=p?��?Җ�>��d�����䋿����t}�͝2=���>�O�O�U��K�>�3H?(`>3�'>�nӼ�U���x�O��F� ?焖?-�?쵋?>|>�����߿�[���?�X?��>5!|��\?�M=[z��Px����fS�l\��]?��+^q�������6��.��&���bU=g�5?֜�?�b�?e_�?��ھ6�Z�l�Y�G�w���5�@��3���E��	_��ET��h�����b��澝C�0���o�P���?�nO?���o��>g�������ɹ�[��>�A��Vׇ�Di��8����<h1P>��ʾq�^�cp��#�`?��>�>��%?Ra�aT6��=�{������>�>0��>&?,��S��������ξ�c��	=+>v>�uc?�K?�n?�h��)1�������!�Sj/��i���B>�m>���>�W����8&��Y>���r�c���w��~�	��~=Ʋ2?�,�>��>M�??%z	�fl��5qx���1��<�<�(�>�!i?�B�>���>hн�� ��~�>�j?S�>�$�>�L���� ��|���޽��>�B�>#d�>mq>��3�2k]�Ў�xs����9����=} k?�
���Vb��_�>>�S?c�M<b�<���>���2��N��G1�C	>a?s�=A�E>z?���M
��oy��I��HL)?P?ܒ��*��G~>�&"?�z�>�&�>/�?�%�>Ctþ��B���?	�^?�AJ?�SA?EH�>�=` ���WȽ�&��,=>S�Z>�m=c��=x��ik\�s���D=�f�=�μ�W��Ď<�y��tJ<
��<��3>�ۿwbI�^Ծ6���� S�\T����Ͻ����>��������N{��	�C(�3X�'Rk�<ǈ���j�|f�?���?�~��*p�Z������ �U	�>kNo��[���6���8�2����m�4ί�6#�ӿM��k�c:g�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >ZC�<	-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���~¤<���?0�@�A?"�(���쾥�{=o��>Tc?p]5>�y3�E���Q��\B�>��?.r�?��=xXV�J��Pf?�/<tIC�+�����=&9�=6C=m(�q�C>��>�B�_}ƽv�?>�>��2�_����]��[�<S�l>kɽ/z��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�� ��<¿�/���2�8?�=u�=,�=����U[�\˽�����x��L�˽O��=�?>n0>�r4>Q��>X�Y>=Q\??4r?N$?�F�>�ҽ%����辣������(�*7��X�o����4#�/3�%��Ő��G��W;!=�)�= 7R�i���6� �T�b�U�F���.?w$>\�ʾ��M�"�-<{pʾP���jۄ�᥽�-̾#�1�&"n�c͟?��A?������V�G��"X�y���_�W?2P�ʻ��ꬾ���=������=%%�>���=���� 3��~S��+0?�f?uB�������5)>}  ����<�*?�S ?�P<L��>N+%?Y�)�vlά�_>8>�b�>��>��>O���$׽\�?��T?r��(G��	�>'���3}���e=�E
>�m3�]Q��v#X>���<�����@m��a�<�Q?~	��mq���s��\�ܾ�Td>� _?�?�>���?�?A��r��{q��6����=,�C?�U?��=�>>�Cľة��+e?��?x�x���	��B�uEJ��I���?�cK?�u?J��=RI��䎿�1��F:?jq?b�V�^�������h�>��?g�?�G>�K�>�4W?x���)���d¿�k=��C�?�� @���?�=<^�O�X�9�?Mf�>�Zb�8ržyCt��ͯ�"�<�?Zcp��-��B���0���'?��j?��>�L�ӱ���=6ە�=[�?��?z����.g<���l��s��/͠<Zѫ=� �fM"�����7�]�ƾ��
�����P࿼���>�Y@#g��%�>JF8��5��RϿb��BVо�Xq�)�?{��>;�Ƚ������j�xRu�3�G��H����pE�>0K>�R���ȏ���z�kt;����uH�>xܼ���>iR����杢����;|ۑ>�G�>l|�>�p��绾
�?���SͿ��MX	�_�V?M��?Lم?D�?=l�<��k����e��H?�Oq?�sX?G ���W���M��2h?���� Pb�2q%�<zR�m��=��6?�6�>�E����=�8K>��?��=�-=�¿������ݾ�О?���?u�徶��>�K�?�E#?.;%��9��ĒH��d� ��[>M?_u>Eؾ�*�cG�?wo�A�?z�G?���w&�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�$�>��?�f�=�d�>�p�=谾�9.� ^#>��=�?�m�?!�M?BH�>�m�=	�8�[/��SF��?R��%���C�R�>b�a?-�L?�Mb>������1�n
!��~ͽh1�U6�BP@���,�q�߽m5>=�=>�>p�D�AӾ�\!?�h�QXԿ���$i���?W�|>Pf
?�Ҿظ��ï�<c�m?�!I>F��H���W���,��1�?�?��>=5ξRH7�"X>�S>J�>�t=�S�ޢ����{>1C?�����L�|�S�>]��?lc@C��?=�[���?Ur��Lˆ�ɭn�����t�L�0>��C?K��Eȃ>D�?ߙ>��m�1٬���u�!?�>� �?z<�?���>�w\?��n�&,0��=��y>|X?gB?q(=~�%��>�H?���(T����٢_?i�@��@�#Z?3᤿��ܿ����hپ ⾢/
>�w�=&�@>�Vk��y�<��\=�Ǫ�|��C6�=z��>B܊>���>AJh>�>�/>"���a��^��ӑ���~9���
(	�2BV��!��f��!g�I�¾Wݶ���K综�����<�d!+�3�b�^�=��Y?�%P?d�n?'>?���}�>�>��<��<�0�8:=�Չ>m3?aRN?��,? ��=  ��Y�[��Á��6�����u�>��@>>�>p�>p#�>������A>�@:>"}>���=��)=vl�:�H�<�E>���>���>ɺ>�C<>��>Fϴ��1��j�h��
w�w̽1�?����R�J��1���9��Ҧ���h�=Hb.?|>���?пf����2H?&���y)��+���>|�0?�cW?#�>!��z�T�4:>9����j�5`>�+ �xl���)��%Q>vl?'�f>("u>u�3�>c8�=�P��v��'U|>646?鶾NC9��u�ȮH�^\ݾ�OM>̾>OC��h�T���>���i��{=gu:?(�?�6���ⰾ��u�G���GR>{9\>�o=�i�=�HM>�oc���ƽh
H��.=���=��^>N�?s >xG>=�1�>s˾����`��>R�>��>�%J?�7?�ʇ��}�����Ґc�a�\>T��>f-�>�1>z�>���L=���>'F>.�N���[����^V���l>ӷW��I�7��=�"�sY�=�z?=9�����1��D=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ4��>b0�,M�����u�&"=��>�SH?u����V��J=�i�
?V�?��򾴷��ɿb�v���>���?ʔ?�km��H����?�j��>yc�?D�Y?!�h>�ھ�Y��~�>�@?e�Q?f̵>���j�$�m??���?U��?I>o��?��s?�l�>�x��Y/��6��������=��X;U^�>!Y>p���#iF� ד�og��ѻj����J�a>"�$=o�>�;�7,���K�=@틽;L��]�f�u��>�%q>k�I>^V�>�� ?�Z�>ª�>}�=�[��4���⹖���D?a��?c�ܾ�b���=�bg>���-?�Q ?�Jv�.��w�>��^?�~?f�u?���>U��l������H��$�4=��(>��-? �>�|T�{�>R�B�C����&>�-�>��������ޓa>��>�?"+?�m�=��!?��?�+> �>��J��g���W���?���>���>��f?�r9?�̿�Nf/��V���Y��ʖy��o�>�
�?�{?=�>nӦ�ׇ��������!>_�`?�͋?%��xD�>z�?�#�>+�?c�>>����v�Y0X��>��!?��|�A�eM&���Q~?eM?���>�*��w�ս�ּ*��[}����?�'\??@&?����,a��¾��<^�"���T�]��;B4D���>��>�|����=�>�Ӱ=_Nm�~M6��f<��=s��>��=Q-7������C,?�����僾�-�=s��7E�}�>S5P>({��i�_??�3���z�٬�����MX���?�Q�?:��?bz���/h���;?x�?5�?��>��?۾h�޾0<x��!p�ƫ����=���>��U�Ö������9O��2�˽�a$����>_�>�?�� ?7�M>Բ�>�Ҡ���"���������_����&8��E,���<#��B*1�����>��|�m�	^�>�i��R�>�Q	?+�h>�;�>�m�>k�;���>�>X>+ek>�>�-V>��<>�Q>+q��%�LR?�����'���G����0B?zid?�%�>�h�㈅�����?8��?�o�?�2v>�}h�,+��h?�@�>����n
?�h:=�;�;؉<pP�����/?������>�b׽]:�YM�!of��o
?�2?�!����̾�R׽��y��;��?�G??��(�'�G�N�}���0��ew�im>���`���rR�Tej��x��'�y�!Ɏ��k���=��C?���?}40�:����ľ;��#n7����>��?�Z�=�/�>���>���m�8|�mBb�-�t���?A�?!Gf>�&v?��'?m�O?�E?��>���=>����;>=Խ�<�`�>�U4?C�E?�(M?��?x3?�ƚ>Bپ_�!��n�!?���>]_?Q��>'�>~����<�B;3��<�.�����=:�=b����m�����=��`>�Y?h����8�X�����j>�w7?�{�>n��>�
���+���R�<��>گ
?I6�>� ��|r��a��X�>���?����h=�)>��=,)��C`Ϻ`K�=�7¼A�=SV��:�;�� <�d�=v�=�q�6�Z�wT�:�8�;݊�<�?���>ٍK>A�>k;�����B��!B>ˡ�>���>�Ĉ>xӖ�Z}������fs[���n>��?[��?���=���<���<ߪ��A,�f�E�����\g>��?�7?͝�?�?���>*9,?��>�3�����ȇ����]�>�!,?牑>G���ʾ��o�3�J�?�X?�8a�����;)���¾ս��>�[/��-~�p��BD��*��r������
��?
��?��@���6�}�����X��ʑC?�>�V�>t�>��)�a�g�U#��,;>��>!R?+�>^�O?�/{?	�[?S~T>��8��2���ԙ�6�/��!>6@?��?
�?� y?�n�>��>��)��
ྨ-��L��@�҂�Q�W=�Z>W��>$#�>3��>��=|�ǽr:����>���=�pb>˖�>N��>`(�>��w>�ǭ<b9H?I��>��������>�����=�h?��?AZ?��;d6�J�Q��*���>؛�?V��?J(?�����=��x�F��對�,v�>V�>���>�+>ľ%=.l>���>$T�>����|���g7�zUl�1�?��G?� (<��ſ`Zp���l�����{<z��n�b����[��O�=���S���6[��������`����֝��}����>�u�=}��=��=���<��ü�e�<�M={w�</4=�$o�vb|<�}E����u���qcp���N<·7=�,��۾�[�?j�Q?��,?D?��> �9>Y;�����>NW��h�?z��=K�
����#
2�wl��Sਾ�� �
�ƐJ�φ�6>�9��.>W>>@>P1=E>��=�q�=�6=&�;���=� �=
��=�g�=���=���=�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>;�8>~�>F�R�RZ1���_���d���W�E�!?�9;���ʾ���>��=߾btǾ�&=%�5>��h=����[�Y�=�W}��;=��j=�/�>U9D>D-�=�A��9��=1WH=LI�=PVN>j����0�gs,���0=pq�=(b>��&>���>�K?�z)?M�g?�,�>�7u��8ܾVž���>�k=ۚ�>��=��>��>��3?��D?O?�U�>��=�o�>�>��%� �j��"뾖J����R=E�?��?{$�>�X=+�.��8��5��#ǽ��?7<?�	?�2�>���Pֿ:%Z���h����=���=gЎ>����������v���f��Y�=�?ZQ?��>f �>��f>�AI>���>}b�=��=�6V;����F�c��=�}�>�67<3����	����<b�>S��;v�R��������s�(>��=��=���>Q�>r��>Zh�=.����.>�֖��{L����=IO��*�A��6d�XQ~�}
/��O6�;,B>�QX>�.��^&����?�Y>l�?>���?�?u?��>���pվ�L���&f�wtS�@�=��>�<�~O;��d`���M�EҾ.��>��y>�L>�eo>���F36�v��[&�5@��я�>S������;�l��~����*��wm�͝=�Be?���5#�=�fn?�\?$��?���>�Z`�������J>ǣ��K��	�PO��2.Q��1?=`&?���>�P;��5�ʾc������>6E�y1O�}���W�0�,$�jܴ�n�>������;��3�^���<���^�A��uo�u��>�6P?I7�?B�c�р��N��"�����R?�h?�Ҟ>��?�?�����t�F'��?P�=ƺn?m�?ֲ�?b8>$��=r��N<�>�)	?���?��?ups?��?��~�>|V�;�~ >䞘��m�=˭>7Ŝ=ώ�=n?ڂ
?��
?O�����	����G��^����<%2�=v��>W�>t�r>�W�=��g=�	�=�\>oٞ>�>e>q��>�<�>]l��5����=I?�0>���>�?'?�n>ؗ+=���U,�=�s�a=���B��#⦽�#���v�=q���<Co��W?y$ۿ��?X:�>f�n?��?+�=�Z:=�i�>�ձ���>�k~>�>���>��>��=&��>�L>%@Ӿ�d>����Z!��+C�ހR�T�Ѿe�z>������%������[<I�3r��*j��j�D0���9=����<�I�?������k���)������?�R�>�6?�Ό�+=���>y��>yɍ>�G������%̍�ne�h�?���?2�f>��>��U?k�?hD+�7�3���[�|Uv�?F=�7;f�X�a�(���ԁ�ܪ����xf_?�w?d�@?iF�<��v>|d~?��#�U����>�.�Ω9��Z=f��>u{���p\�X�Ͼ��ž����I>+Jo?�m�?,�?7^�������>(4<?�7?��?�,R?o�9?{���K\�>���=	�>q"�>m�_?E�0?[�?�>�}�=�Ѥ��#���+e�?�����r�Zf��|׼�:��b�>�2ʽ����THd=�1�=bՠ;Y��s���8�<��6<��x�bZ=j>�u�>/N?y �>�/�>�9?>$���E�(�Ⱦ�0<?r�+��/����f�L���
��d�=�lg?{i�?��T?�Ù>�H��d�/*3>F��>d�$>�f@>i��>VZ3�tD��m�=��$>o;>m�<t��W�S���D��X"=��==��>�z>�5����)>I���3Ow��^>D�O�pʺ��R�(�G���0��Bt����>��L?�h?��=���z����f���(?��;?�M?si~?f��=(Rپ�;��IJ�{���>NC�<i��`֡����u�:�`]�;�|>���m�����a>A0�^ݾ��j�D4F�b�޾���<����?=���Fz۾Xbx����=~��=�cȾ{4$�����>��?I?��=��`P�do���>	͒>lݫ>4.1���e���<�MP�����=7�>br5>vhn����z�E�1E�TB�>bPE?�S_?"i�?9���s�]�B�����jj��8XǼ��?�u�>.d?�B>$�=,���j���d�)G���>%��>�����G�BL��Y,��W�$�&��>�8?�>��?p�R?��
?��`?�*?9=?7�>�I��o���B&?$��?u�=��Խ��T�� 9��F�n��>��)?��B�i��>މ?�?�&?υQ?��?��>2� �!C@����>�Y�>��W��b��e�_>��J?=��>�=Y?�ԃ?g�=>�5�@颾(٩��V�=^>��2?/6#?V�?��>L�>PS��<\=�>:+i?���?
%t?6�=	�?��N>`�>�'�=x�>� ?i?��K?��m?�OE?1��>���<�谽7ϩ���1���<"��<��O<&�I=^��	~�tOe��� <l"�<����W����K��L?�M��t<>Z�>�t>������0>i�ľ�\����@>N
��z>�������::�6��=a��>?ж�>�y#��v�=d��>n?�>����$(?~�?c?%�;}�b���ھ��K�f"�>�B?�	�=��l�郔���u�ثg=��m?��^?�OW�|�����b?^l?�b�e6R�S:��PӔ�י�0�X?��>]�����>M�v?��j?Y�?���c�����g	_��(�A_=��>����d���>��-?���>�Vr>�
�=�)���N�S}��7i3?���?%Ƞ?���?�s�=��o��ݿ��+�;|u?#U	?�窾�Y=?�=�% �M����ݾHo�0��5�H����ɾ�*��yz����!��G�;�|+?�o?��Q?�t@?��$��2��k�~���p�f�B�1�󾇂�s�M�o�G�O$F��&5�#�̾��Ѿ�Q��-w>>�v�Z�I���?[53?C�"�L�	?��v�����uCݾ���=٪��O����=�NܽC}��9ְ���y�&<���ʾ�*?a#�>kϿ>��6?�C]�D{A��f6�^�5�����>L��>#�b>_��>�_�t��g��O���b���k��1v>xc?-�K?��n?�j�
*1�ń���!��/��]��=�B> m>���>�W�!��!:&�Y>�D�r�����u���	�֢~=E�2?�'�>���>�N�??�y	��i��>fx�ۇ1�ky�<�)�>�i?�B�>P�>;�Ͻ�� ����>��l?o��>��>斌�jZ!���{���ʽI&�>E�>"��>��o>�,��#\��j��I����9�Qu�=,�h?
���C�`�?�>lR?��:�G<�|�>^�v��!�����'�O�>`|?���=0�;>
�ž�$�o�{��7���#%?�
?����*����>�y$?\g�>7�>��?���>���B�=�B?j9b?
�E?}=?�]�>��={㒽Pɽ-�$��'@=�8�>oml>$֑=D�=y�.�^�f�7�?��<�z\=q.��7�����<���r�<4G=��>�]ۿaK���ؾ��������	��G�������뇾-
�-���ou��&�w�F
���,��{W�wd��)��ռl�]\�?�!�?R���,�����槀�����(�>�rp��:}��۫����BJ��;v�3����Q!�#%P�3Qi���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@s|A?Q�(�n��
V=���>O�	?Y�?>MU1�3H�c����V�>�<�?���?�M=��W���	�&e?wi<��F���ݻ��=4=�=�@=f����J>�V�>Ã�aTA�oEܽ��4>N؅>y"�s���^����<��]>��սDB��RՄ?�x\�cf��/��U��
P>��T?2�>�B�=��,?�5H��{Ͽ�\��(a?p0�?��?��(?ӿ�ך>��ܾN�M?�C6?��>�c&�L�t�*��=����ڦ�>��I*V�<��=E��>��><p,�C��b�O�������=����ƿ.�$�p|�Q@=�vպ�G[�2��ܪ��dU�=-���ro�Yf轧vh=�f�=�dQ>h^�>@W>).Z>veW?��k?9M�>�s>7c�}����ξ"P�b;��V��4���k��� M�B�߾��	�3��o��m�ɾC=��,�=r7R�D���&� ���b�<�F���.?Qn$>�ʾ,�M�k�-<�kʾ���uĄ����2̾ڗ1�n��˟?�A?����H�V���EN�{��_�W?�J�����߬�L��=t찼��=#�>���=r���!3��S���.?�G ?�����q����/>އ
���
=0**?A ?U�=���>t�)?R��п��,d>�_$>,"�>:s�>*v>2����=�4G"?��S?�������9�>�=Ⱦzmg����=%q>�LE��JO�ލM>o�O<Z���׺]rT��>=2W?֪�>�*�D���������J;=��x?�?��>9wk?��B?�<\����S���
��Pz=��W?�i?O�>7�y*о���=�5?A�e?ccO>�.h���"�.�XL�15?j�n?�q?�!���m}�������=W6?�w?��\��������\���>���>��>�6�|V�>��>?�Q$�H���f��<�3����?��@���?�&<�$�LN�=)� ?5W�>�QT�!�ľ��#���xQ=���>B ����s����4�%�;?._�?�+�>���9x���=ns���\�?"5�?�����s<���5l��3 �4D�<V"�=�!�T#�>�@�7���ƾ��
�Ah��󒽼*�>�J@Y_�A�>��9�2d��mϿ��6о��q��?�$�>��̽����*j��t�f G�2	H��[��[��>�>����,����{�Ud;�h�����>X��2��>�S��1���%��yH-<���>Qs�>Y�>k	���彾���?Fh��M/ο�������X?m�?�f�?�&?K�G<S�v���z�`��2BG?ٻs?8�Y?�D&��]���6�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?ӵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>jH_���u>����:�
i	>���?�~�?Qj?���� ����U>
�}?��>k�?� �=d�>�d>�ľ�����5>�>N��=HO?�I`?��>��8>(᥽�2.�H=�K�M�Hk�/�A�o+7>T�s?)�I?=�8>�W��R�<=�r8��%;�Ũ=��:=0���/2���0�&L >�F>�C>� qS���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?q��P��a~����7�}��=
�7?�/���z>w��>�==ov�绪�P�s�u��>�B�?�{�?���>��l?U�o�U�B���1=�L�>Ԝk?�s?��n��󾀲B>��?�������K�;f?��
@iu@I�^?�B׿ܚ����þ�˾A<;>��>gkY>E>]���=X{=� =�#'=�@>�6�>�
�=��D>:�>�u&>$�%>�^��֖�����X���<���J��u�D�[�������I�羹h���:	�:O�o+�AM���#�PJ�G>�=��U?�vQ?3�m?U ?T8���>���z�='$��ޒ=[��>�(2?��L?zz*?���=����Qd��D���ȧ��Ĉ�\��>�
L>���>�R�>�j�>;��>iM>�-D>��>���==Ò���=,)P>-��>U�>,O�>�C<>��>Fϴ��1��k�h��
w��̽1�?����Q�J��1���9��Φ���h�=Hb.?
|>���?пd����2H?#���z)���+���>|�0?�cW?�>����T�7:>&����j�=`>�+ �yl���)��%Q>rl?B�e>bCu>�C3��R8��P�i����|>A�5?�����9�%�u���H�I<ݾ�cM>�U�> �O���������Si��[|=&`:?�}?�������;�u������Q>�\>�2=�!�=�fM>�c��1ȽZ�G���0=�t�=OL]>��?3S->7(�=td�>�9��c�O�ݧ�>'P@>�5/>��@?0�%?G���R6��E���1A,���t>2��>V>�k	>��J�:R�=���>Qa>O���~��%
��*B��W>���,y^�|�$t=2������=e�=_����9��T)=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾQh�>xx��Z�������u�n�#=P��>�8H?�V����O�d>��v
?�?�^�੤���ȿ5|v����>X�?���?g�m��A���@����>;��?�gY?toi>�g۾B`Z����>ӻ@?�R?�>�9�~�'���?�޶?կ�?wI>d��?)�s?�f�>E-x��X/�)3�������I=-�W;[Y�>G>����pcF�Dד�{h��P�j�r���a>c�$=q�>v<体/��g@�=�苽LH��q�f� ��>f*q>��I>T�>a� ?`�>(��>��=�Y���ۀ�����F?. �?�� �	�t���==p�;����5?��?�u��S����>Çi?c�~?��Y?��l>��������,���DӾ�䔼;C�>�F?�?�~E�;��>F$�~���@@�>@n�>���=ڿžCq�հ��Fx>��-?���>��}<]($?�i)?kx;>q��>zmC��9��!Y����>|n�>A!?��`?A6?o᩾�&���y��$���P��	>�ax?��?Q��>���h���gbH��c_�/��G�w?�[\?I:��F?P/�?5�\?�[?�<�=QZH��(�]^��v&>��!?���A��K&�����?�Y?ٽ�>!����#ս�Ӽ���W��a?`\?x7&?Ø�V$a���¾���<��"�iTR��R�;��B�p�>��>����7g�=:�>\��=`qm��'6�k<^|�=`v�>X�=��6�p���M><??o�<��ܾ'f�=@Y{�~:H�t�F=���>P����7?����&V�w�������Z[><�?�6�?�?�?�68�"�V���?Y�?�@=?�<?�z��WGѾ �'��k���a�l�L�t��=�S�>~|�<���^����W��+����͓=�B�����>l�?t��>�>S�\>]c�>��˾0A6����o�d�1����d�S��6'��N׾Oɞ��q���nu�jp���1�>1��=�F�>N�?fM>�Wn>�6�>�ػI�>��4>x�r>v+V>��<��1>���>|L%>����KR?�����'����a���q3B?�qd?�0�>Si����������?���?[s�?=v>�~h��,+�\n?�>�>A��2q
?LU:=�5��A�<�U������2�������>#F׽!:�mM�#mf��j
?�/?���&�̾�<׽�����K=`��?F�!?��%�WG��8b�,�Y�e�T�؇��m͆�=����fm�X��ɤ�����(�,��3=O�*?�U�?�����E�c\��"6o��w?���K>{��>���>���>4�'>EK
�4Q,��!V��#�0ǔ�'f�>:�p?J9�>_�H?��8?F�F?�?I?rG�>��>&#��]9�>��P=�.�>�q�>�{8?�[/?��.?��?��#?OPR>U�ǽ�T��ٍھ�$?��?�y?s ?��?}���⚽����+}��ꌾ����x4=�O�<y����>�"��=2#g>ś?�v
� �5��=���]i>�O5?EG�>]޻>��l���A��@�=ߘ�>��?'�>�`��ںj�y	
�4�>� �?O����=��+>���=��	�<�>|3L�!ށ=>�������<G��=��=Trl���"T1��P�<@�w��?��?)��>��>ϒJ�����R� >b>cp>I�=��Ѿ� ���𕿷�K�t]a>㰌?�n�?���=Y��=.g.>�ˑ��`׾�i�ɒ��K���>��?�p\?�Y�?+1G?]�3?J�>&]��:���Eɾ��?" ,?��>���ʾ����3���?�[?�8a�����4)�L¾x�Խ��>�U/��-~�����D�������������?��?�A���6��k�R���uR��ܝC?�$�>�O�>��>�)���g��%��;;>���>R?Y��>=�O?�{?�T[?ьT>7�8�����,���|�#��l#>
M@?*��?<ڎ?��x?z��>�K>��)���E���]1 �|Q��}т���X=��Y>A��>�B�>�v�>&��=$�Ƚ����4�?��F�=�8a>H=�>��>���>B�w>�·<fX?J� ?�����c�� ��aX־ %ƾ���?7Κ?0�>y�-<�v������0�=|�=~�?㘻?��w?�t_��>��L�ȿ󾕇ܾ0�>_��>)	�>�'�>v#�=es>� ?�>R5ɽs�1���$�x�?>RK?t�$?Q�Y�@����G�c{������hl:��u��ѽ	'`��{��(୽�r�~f���8��X�:�mƾDe׾���]�Ȏ���>�%>��>�ϼ=�"=!���@��ڼr=�
�<��H=��4��u�Ͻ�=��}�d�.=�����;�"��˾Y;}?]I?Z�*?suC?��w>�T>J�8�
@�>4wx�'?'�W>�lL�e����9��m��"�ؾ��վ�c����>AD�z�>Z�3>���=��<���=�4m=�k�={8���=a��=i��=0�=���=��>HU>�Tz?��q�}\���T��C@�c�-?��q>)�Q>�j��Q3?��Y>�a~�3Ǻ��/
��Tt?�&�?:��?��?@�e���>�Q��1⾽��=:a�kE'>r�>�^:�܁>��>�����1�W��?��@��$?��e.Ϳga7>�7>�&>��R��1�@�\��b��yZ���!?�H;�sI̾07�>��=�)߾?�ƾ}.=܆6>�Lb=�m�XV\�=�=s�z�I�;=�l=�؉>��C>�|�=�3���=ϡI=���=A�O>�ݕ�Ѽ7��9,���3=���=��b>V&>$��>=�?pp/?8�d?jظ>�Ru���Ѿҿ�:r�>t�=��>0Jz=��9>ժ�>l�7?n E?�FL?Bp�>�9�=x��>�Ǩ>`�-�.�n�b�ᾥ����ي<a�?9�?�E�>�>`<Zy=�V���=��нE?�(2?��?g��>�O����".��I�������=��>Y`��|����C��=��{R��^�x>�X�>�z�>}�N>r�9>|>4[�>���>F�>���;U�*�Zl:�*�N=�=/�>�ZU=Ȗ�$L����[���;J�=���<�����<*��<��=[��=	��>�=>v��>���=^�� (/>����\�L��ҿ=W���)B��4d�kI~�}�.�9Q6�5�B>S@X>�N���1��>�?��Y>�c?>Z��?I<u?^�>�+���վqI��*e��8S��=է>=�}�;�&a`���M�,kҾH��>_ߎ>/�>[�l>�,�C#?���w=��Xb5�r�>�|�����)��9q� @������qi��~ҺנD?�F��E��=l"~?�I?Y�?��> ��نؾ);0>�H��V�=m��*q�i����?'?��>�쾣�D�SE̾7����>u5I�U�O�����>�0�y��WϷ����>q���}�о�$3��g��������B�Jr�Y��>b�O?+�?0b��W��\TO�h���>��	n?~|g?C�>�I?�??�#��~�dt��x�=��n?���?l=�?>_Q�=B೽y�>�?ʙ�?���?��s?X+@���>I\�;N`#>������=߷>+��=���=\?	1
?&�
?������	�� �9�z[��� =ˊ�=4@�>u׈>�5o>���=��V=ɣ=f-^>�E�>���>��e>ۜ�>��>�Ҳ�zn	��??S�>i�>L�X?�Ū>@Zv�>�/�����'U��ޗ�ޫ����sI���/�A�����x��p���M	?m�̿w�?bf�>QG��%?�g����;�D@>��=p��M�>��=*e=���>���>�>�0�>Fm>�FӾx>����d!��,C�9�R�a�Ѿ}z>�����	&����ix��,BI�hn���g��j�N.��b<=��Ž<&H�?�����k���)�����[�?�[�>�6?�ڌ����/�>���>�Ǎ>�J��c���Kȍ��gᾝ�?��?�>�Zx>:�V?��T?#L��]g̾�h�=�_�(_5��t�G�]����ą���G�G�<��R?��h?��W?�c>k֛>�X�?�Q��j̾H�>S�[��v�<��>ť'?�c��!*��d��<4���ɾ�>oŃ?F	�?�H?c� ���c,+>��>k�> �v?pZ?��N?�l���K?��?&�F?ԞD?�`=?��C?��>� >���<�
ӽ�m�>����5+����ܽ��<��8>9��>�b}>'�������u��\Y��=���v�=\J�=M�м��>V=�"=t�R=C֦>b�]?�:�>�Ȇ><�7?]?�O~8�I���b�.??�:=�邾���2ꢾ
1�c>��j?#��?�WZ?��d>��A�&�B��k>�*�>��&>�\>��>�ｴ�E�n�=;�>x�>��=�qM������	��ᑾ$d�<�f> [�>hu{>�䎽+>�b}��a>'�N��Ż��oR��}H��1�n�y�Ed�>�L?A�?��=1��I>���f���(?�k=?^AM?q2�?$�=Bqܾ�.:�&K������>w=�<zn�����U���;��n�t�m>hԜ�����4<M>[]뾫�PGb��2���ʾ�p��}�eh=ř�Ώ�3���8I�=+;>i�о�1� w��G٪��\F?���=����P)���þ�=]�u>��>�&��ܴ����:�jl�����=��>�f>�%����$F���f>�>GQE?(W_?k�?"��9s��B�_���pc��rȼ5�?ix�>!h?�B>��=^�������d�}G���>���>U��>�G��;��>0��"�$���>59?��>��?N�R?��
?r�`?�*?4E?�&�>C������jA&?��?R��=`�ԽQ�T� 9��F�i��>τ)?u�B���>K�?d�?�&?��Q?=�?��>7� ��A@�B��>�T�>�W��`���_>K�J?���>�;Y?Fԃ?w�=>D�5�좾�婽�D�=g>��2?C6#?��?8��>���>M���
?=f�>�7_?w&�?�u?P4�=�i�>��#>=��>��=L��>�$�>�?GK?9h?�??���>�`�<c@��z]ŽkE������<�TԻ@ul=Io��6L��둻�u�<��=r,�:�<����"=��&���65��_�>��s>C	��r�0>��ľ�O��s�@>I���&O��ي�l�:���=w��>��?窕>�X#�c��=?��>7I�>���T6(?��?�?X�!;r�b���ھ>�K�h�>�B?���=��l�������u���g=��m?��^?��W��$��#�e?m�x? `�JNP��)��溾�p��k?�d�>�] ����>=��?�|?��?�O��Jg���,��S�i��6!��z�<	�>K����Y�ǰ�>]�$?h��>YM=H�>y����L�I�.��7?��?s��?�a�?���=�.o���[�;�'���li?z�>P"��A�?{� =�,���.��ɿ|��A���۾�g�������X��jp��A����ǽJ(>�(?xЃ?>�?`D|?�<+�Żz�R�k�Y�c�-[^��]�.����V�i�28;�<|�Ŗ����V��
���>�m��K�A��Ĵ?�V&?c/��X�>����8���̾�j?>�#�����d��=m�����I=�N=i�n��3�!S���t ?��>R��>Y�<?R�\�m/?��w1���5��4��{�/>4�>]F�>���>;¦;u�.��X��Ǿ=�MHݽ�vv>|c?��K?^9n?L����1��.��{� �!g!�v�fdE>x
>���>V�V�4�s	&��=�%�r��b�	���5
���y=��2?\�>��>��?2�? ���į��gy�>�1�Y<'A�>��g?���>j��>E�Ƚ���d��>�l?-��>/�>�����T!���{�Q�ʽ� �>_�>}��>i�o>��,��\��i��\~���9�<J�=��h?:|����`���>*R?6^�:�[I<3��>��v���!����y�'���>�}?:��=��;>�wžk'�F�{�f!��9
(?"�?�J����*�O=}>#?���>C��>a��?��>5���<6;?�m`?�lJ?I�@?��>�t=���=�Ž�(�	%=���>\[>�9~=]x�=����O�|D�kfF=L!�=v�|�=������;a����n<���<��3>��ٿ�G�4t��#��#ݾ�o�<�`��-��+�������ž���f���.������yt�A���u���*l�7��?���?�[��?Z����_ȃ���2��> C>���[i��?\Q������Pž�
��+����R�9p��r�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@.|A?
�(�4�쾚V=��>Y�	?g�?>MT1��H�����TT�> <�?���?͒M=�W�E�	��~e?�G<��F��ݻu�=}<�=b9=�����J>�Y�>����WA�FNܽ�4>�م>�o"����|^����<��]>�ս	4��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=� ���Ŀ��+� v.�=t>�$!>��$=�k���xg���=�3��Cj�5�߽��;w:w>;��=��=�;>w�H>�R?ڀ?��?Z�>s���2�Ӿq�彘����x�H�о�j��5����(�u��҄
���1��.�.UǾ�#=����=y0R�����M� ���b�ߐF���.?�h$>D�ʾ'�M��+<Jwʾ������a���R9͚̾1��!n�̟?��A?��[�V�7�)������]�W?�C�����k��=�:�� �=��>N{�=����!3���S�� 0?�'?<����؏�H'>�Q�]�=f�*?�?Sh�<?e�>�Q%?�(�޽6V>�1>T��>�>�A>�@��/�ڽH"?��S?�� ������?�>������}�M8O=�h>a4�f/߼6K[>���<.����i�ե����<8W?sύ>
�)�Ӣ��9��0%��|6=��x?��?dt�>d{k?��B?F�<����=�S�!�
��=7X?ħh?�m>�S��tlϾ�m���5?�e?��O>ri���꾼/������?��n?W�?`	����}�I2���^g6?��v?	Z]��:�����Z����>Ç�>ER�>�8�9�>�r>?�$�o^��!翿y,5���?ڤ@]��?uS�;�2 ��8�=t�?<!�>��R�͓ƾ_��� ���&%u=D�>Μ���(u�����,�ޕ9?Mc�?���>PÁ�����=����]�?��?�����g<���\l��{��E�<-��=���X"����7���ƾ�
�{����J��M��>&Z@'��:�>�^8�8��TϿ����`о�_q�?�?�f�>�Ƚp�����j�3Eu�r�G���H���� P�>��>K����򑾭�{��s;��v����>���� �>��S��)��՞��2D5<L�>ͳ�>*��>����⽾�ę?�`���?ο�������X?�e�?�o�?�r?�
9<��v���{�����+G?6�s?�Z?*O%��3]���7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�d�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�6�>=�?.��=���>,��==�����+�|�#>�q�=��2���?��M?"�>*�=��7��/���E��XR����ƀC�2�>�a?mhL?8Gc>|ŵ�#q$�� ��ͽ��0��q��@���/��⽨x3>m�>>�#>��B�1mѾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�n	?��CP��A_~����7����=�7?�,�?�z>���>��=�ov�������s�M��>�B�?�{�?���>p�l?��o���B�q�1=.P�>M�k?�r?�)n�@󾷲B>5�?�������UL�f?��
@Su@�^?�@�ѿ���n��'���>7�A>�F>���>�%:>�=$>��<�rW>UV�>(s�>�>t��=�|J>+�^>ʁ�?�!��.��V���S4��l��۟��+��~F˽*����ž҃��A<�S��+��H��v<��Y=u
P?��`?�R?�%?�}����=�����<Piϼ5�t=��H>�$?61?	�?��j�X�˾C�i������P��Q���F�>��>$O�>%5�>��>9�=��B>p�>��[>�~�>��.�[�������{&�>��>��?˴�>�C<>��>Fϴ��1��j�h��
w�n̽1�?����S�J��1���9��Ӧ���h�=Hb.?|>���?пf����2H?&���z)���+���>|�0?�cW? �> ��z�T�4:>8����j�8`>�+ �|l���)��%Q>wl?�=Z>�v>	�/��<8�͒O���E&{>o2?h��r�6��v��L��۾�xQ>�R�> L��z� ��?���$��,Yd����=��9?,?H���䞫�a}��t��ǈN>�b>�)=mʠ=�8Q>�\M���˽>�C��G?=���=�Z>r�?�p3>���=��>�͜��N�Į>N7>��2>��??��"?��}�+�p�g�n�Y�E�;�d>r �>�q>�>@2D�) �=���>�Y>�$��&W���ܽ?�:�_M6>!����[�3�_����=	����k�=^Z�=2�	�[�:�JB=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>zx��Z�������u�s�#=Q��>�8H?�V����O�e>��v
?�?�^�੤���ȿ5|v����>X�?���?g�m��A���@����>;��?�gY?toi>�g۾<`Z����>һ@?�R?�>�9���'���?�޶?֯�? I>���?��s?�k�>�2x��Z/�y6��ؖ��/n=�[;ld�>2W> ���1gF��ד��h��=�j����[�a>�$=�>�D�c4���:�=�����H��ֹf����>�,q>��I>"W�>�� ?b�>D��>�v=2p��Uှ6�����C?ꨗ?�=����o���l=�� ������/?Ǐ5?�">t*]�i�?��y?{�?C�j?�C�=h���.��!��/ɾ���2@�>�l?�?EhJ=�Y�>\��7�ҽ~9�>��>�w�|,۾7,���cP�m�>}�?���>,�>f�'?K�%?R[>ۚ�>T�G����J�Q�)�?��r>U�?G&`?��?-+��p�8��U��%���b�K��l�=論?+-?��>�ޗ�aF���-v���U� l�y?�?N�Y?SY�� B?�?K�`?"�[?Kc�>9Y���)�d�#��hh>v�!?\��z�A�4U&���� �?�?�U�>V쒽8TֽQdȼ�a��|���0?[8\?�=&?�|���`��j¾���<�#)���e�yx�;/L�O>��>KM����==�>v�=�m���4�<�u<�;�=�|�>���=�W7������A?��>�Xk���y>�톿hg�Ԫ�����>�ۃ�r��>E���#S�>���8��;�I��d?��?6��? �>� �B���?1�?a?��>� ���1n�	t
����:�Z�F_��F[=L��>K�<<)�1�`6���ꣿ����H��=m�]����>��>#�?�?6��>�y�>����*�^�־�=�z�Y����`=�G �</��þ-=�ґ1�zU���N��DHw>$����=�>ު
?��>��>I�>p(�:�Q�>ђ>Un>L�c>��3>�1>\;.>��=_M��YKR?w���?�'���辈���3B?\rd?�/�><i�Ɖ������?}��?7s�?q:v>M~h�0,+��m?!@�>���p
?HR:=R_�hi�<�R������3��
����>�D׽�:�zM�zlf��j
?�/?���Q�̾{9׽ޔ���o= N�?�(?��)���Q�b�o�>�W�S����NPh�x��P�$�_�p��菿S]���%����(���)=ˇ*?��?�������!k�Q?��vf>� �>��>�ܾ>8~I>��	���1� ^�PJ'�ʹ��]L�>�Q{?6&�>@�G?�9?.�@?�n@?�qd>��>3���?���=!��>>�?l;?^j#?��?� ?2�?S>���t���|�D�> �?}�?��
?<�"?^愾�z��굽��Y��·��ċ��<�<>M�5Y�T'���>�Ն>��?usƽ+��Pپ;>Ԇ'?!g�>5��>�fZ�t(&���_=���>e�?��>W��� a��}��>@|~?��ȼ�=1v->�ϯ=��ż-�g<�F�=�k
�p»/h��AN2�̜�<�p�=�A�=8���=u��+��Ʃm;R2�<a ?a�?�v�>�c�>W������j-+�bU~>V>v�=�rm�Y9ؾ|��ن����f��s>���?kP�?o�I=9h�=�h�=����]Ͼ'R뾓K��$u�;��	?�@?�]?���?fM?��%?�-(>�Lݾ�]���ۓ�or˾�5#?q!,?��>�����ʾ��Ӊ3�֝?c[?�<a����;)��¾ �Խӱ>�[/�g/~����>D�󅻼��J��3��?꿝?�A�N�6��x�ٿ���[��|�C?�!�>Y�>��>R�)�{�g�o%��1;>��>iR?�>�HP?�{?�Z?�V>R18�d묿�,��^K���.>0-A?X�?�Ҏ?>�w?���>�>*���h���$%+�� �e���|r=vY>b�>���>{B�>��=��̽Wp���D���=��U>���>�֧>���>�V�>�'�<�+[?6z�>�������N�����^�ʾ,�?��?pD�=�t<I�"���n����7Y/��u�?��?[(j?�틾W��=B�+<Ѧ�F �_��>��?Iv>+�>�>o��>�@�>)��>+"齎�'���	��T�$?��Z?b��������c��K�[L�B�>d��j��#�4����6�=V���v^������Fk�Ro�&5��GTپ��� ���' ?ef�;2?=]��=�7<�H׼�A﹌�=�B�<��O<#`������w�:c��=\2@�2�
=�y�<MOԼ�U<��g�X?[I?S�-?[?�}�>�"^>M��Ζ6>6��[�>p�->�:z�[��A~1�����G�����Ҵ���;1��¾nG��G<�.>�)I>]>B^�<V�=���=zŻ==g�=?�=U�>��<o�>�K3>�ig>�6w?X�������4Q��Z罤�:?�8�>i{�=��ƾq@?��>>�2������yb��-?���?�T�??�?Ati��d�>M���㎽�q�=M����=2>s��=w�2�T��>��J>���K��D����4�?��@��??�ዿТϿ6a/>,�7>C*>��R�G�1�>�\���b��XZ���!?$C;�8=̾�6�>_�=߾�ƾ�E.=D|6>�Zb=Kq��L\�&�=��z�M�;=��k=]؉>J�C>��=�0���¶=#XI=���=�O>����.~7�$�+���3=<��=٨b>�&>��>�?�b0?]_d?�ֹ>.�n�WOϾ4������>��=�V�>̈́�=S�A>�M�>Q�7?�D?��K?B��>cۊ=<�>9ڦ>#�,���m�=��씧��Z�<���?�φ?�N�>O�P<�A�ի�y>�7�ƽ��?�d1?l�?��>�6������S�@pG��_e��>�>6M��e��<�0>��йN���W��=�h�>��>�Sl>���=��r>�sx>7h�>��#>cL>9 V>�f=�(=m7=�����^�s!�;��ąM<�h�0j)�Wџ�]٫<C��<y;�;���?e�=2)�>z�>rd�>KF�=������,>�땾 M��Ĺ=<9���B��bd��z~�J�.�5,6���D>׵Y>CH����ʕ?��[>2R?>�\�?f�t?�>���B�־�Ɲ��h���S��X�=�>.�<��|;�S=`�S�N��.Ѿr��>dߎ>�>��l>�,�I#?�t�w=��_b5�B�>�|�����A)��9q�@������Ei��PҺ�D?�F��<��=i"~?�I?`�?���>P��׆ؾ�:0>�H����=c�*q�i����?'?̗�>���D��'̾$྽~�>f�H��P�UǕ���0����Z����R�>������о�-3�xe�����SpB�� r���>��O?��?+b�\[���\O�Ѽ�u>��TU?�g?3=�>6?5@?�����}�9���� �=��n?��?�<�?�
>3�[=��آ�>rW?�/�?��?��q?�,c����>�V�<��>^۞�R��=(�=���=�y�=���>���>�>�>~�F�����������b����<��=�>kÈ>gEQ>	��=��+=7&�=�Ń>�"�>�M�> �X>8ކ>V��>�ܤ��R+�c?�>%>t��>��6?]ѣ>�7O<F{���������;�<��٪����<�W���_�<xN�j����ĽzD?����X�?6��=W�<����>�8�?�*=�Je>�~�=�������>}�>C��>���>��>Ϡn>pI�>��N>dGӾ�>3���c!��*C��R�`�Ѿjyz>Ý���&�@��?{���BI��o��
g��
j�T.��%<=����<�G�?�����k��)�����]�?�\�>�6?ڌ��
���>���>�Ǎ>L������Ǎ�cfᾶ�?���?AR�>u�>?�|?�]?,d��5:Ⱦ`_�u�B���7�ܢ{��@X�Kܟ��9����x��ZG?¨�?��@?
�>��>��?��=�Mr�
ׂ>M�u��腿C$�>S�?���Yzi������򣾜{뽱#x?��?��-?fB�mw5=Y�A>�`�>7�>�c:?�F!?bAf?Y<<�r?�Q>M[?%�%? YC?�=?���>��->Э=p�ѽ���>�1x�c���:�V`$���_)>�`�=�N��M=���<?]�=��h����=^>C�=މ�=�*�=��=���=d$�>�q]?�f�>h�>��5?� ���8�}���J-?��)=&(��L���1���|#���� >�Mj?��?�aZ?��a>�&C���B���>�>i(>B�[>�C�>4�콧�E����=�m>�>c�=��V�V���y�
������<">>��>f7|>����J�'>&���2@z�Γd>V�Q��պ��T���G���1�!�v��J�>��K?��?��=W�/��Hf�`-)?_<?`KM?��?��=��۾�9�>�J�}(�b�>F?�<������j"��M�:��`�:e�s>(������ȶg>\���Ͼ�[�6�C�=ܾ�M�<����=b=��
�>�׾W�t���=k��=��Ǿ��&���,w��`nF?�ƨ=Ņ��R�0�K�����!>�В>a�>[\���Ƚ?I�(&��,x:=T�>|Q6>����Z��J���n>�>SQE??W_?k�?"��Zs�?�B�����kc���ȼF�?hx�>&h?�B>���=G�������d��G���>���>f��J�G��;���0��M�$���>T9?�>��?\�R?~�
?v�`?�*?EE?('�> �������B&?̇�?Ƅ=4�Խf�T��9��F����>�)?��B�|��>f?ͱ?Q�&?��Q?+�?;�>�� �tA@�琕>�S�>��W�{b����_>��J?��>�=Y?�Ճ?��=>p�5��墾�ũ�-[�=�
>%�2?�/#?��?���>|��>L�����=ƞ�>�c?�0�?!�o?��=<�?�:2>N��>&��=���>d��>�?SXO?>�s?��J?��>I��<�7���8��Ds���O��ǂ;duH<��y=��
3t��J�7��<��;�g��>I������D�7������;ȳ�>��t>�ޕ��1>��ľ:���k@>>�b����{����6:���=���>�?�P�>�� ��=�y�>��>��I$(?M�?̓?�E�:�Bb���ھf�M�a�>ZA?��=�=l��E��5{v�Ѱe=��l?=�^?r�U�����7`?�g?e�����E��<��O��/�ѾNsa?u�?�Z��L�>Y>�?�-y?�n�>,.m�ro�Y���TX�eM��=�v�>/�Y_��9�>��<?��>r�m>f1�=3Ⱦ��s��+��#�?�??f�?:�?:>�"m�x�׿�[��H���>V?D�>�N��?o��=�)�,x����4�BK���v�ܿ?��d���ݾ�~u�����p�� ����b?��w?%�p?�Yk?�%���L���^��6|��M�^�,u5��y^�@�L�h;��P�	���<1�D�����g�ZL���$a�W�?x�;?�����?
]��ue��M����A%>��;t�����)>�ʽ?R�:񫽌�{�P�;C�/�1?O#�>�S�>�;?F�9���5��D3�q�H���$��$!>�5�>+/�>틬>,Ռ�>;���y�=�s
��A�DM=��7v>�xc?\�K?��n?.p�+1�����W�!���/��c����B>�j>4��>"�W����R:&�tY>�M�r�n��w��:�	�}�~=��2?~(�>J��>�O�?�?�{	�yk��2lx�5�1�B��<31�>� i?A�>�>н2� �J��>�l?1q�>���>C茾�y!��{��ɽ|�>v0�>���>�ip>�?,��\�Nd��H���9��
�=^�h?ք��X�`����>E�Q?�:��K<�ɢ>эt���!��q�-�'�T\>�?�m�=�J;>ѩž�:���{�e!���4?���>V໾I�0�F�x>X�?�b�>�P�>�?6��=�᧾ː]���>Z�r?d`?�Y?	��><��;��=����ϫ�=�(�>��>I!.>=�L>��:�2���}��Ѱ=v,>��"=��(�hA=W����2��>�;|�<>HmۿBK�ږپ�	���=
��ሾ{���8e��©��[������Kx�G��l4'�C!V��<c�𤌾��l���?�<�?�x��X(����'����������>��q����������_-��Ŗ�����c!���O�'i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@}A?�(����jV=!��>�	?��?>�S1��I������T�>l<�?���?|M=j�W���	�)�e?�<��F�:�ݻ?�=�;�=3E=���t�J>U�>����SA��>ܽ��4>Zڅ>�~"����[�^����<��]>��սi;��Մ?�y\��f�n�/�9T���R>;�T?g+�>�H�=گ,?�6H�||Ͽ'�\��+a?.0�?���?��(?�ۿ��ښ>��ܾ*�M?�C6?"��>c&�	�t���=�Y�jä� ��%V����=���>2�>},�)��Q�O��S�����=|��=�Ŀ��"�G����a=��<J�м����潽!�����M�O
���+=9��=�>>��z>��G>7�:>>T?5Wk?l��>�(->��XΈ� �Ͼ��̼Nׁ��*6��_��0�D����J�n)߾X*����?b��lо�m<��!�=�XR�1���<!��c��F��b.?��#>� ˾��M�.^�;��˾Oߪ�a���١���=ʾl�0�zn���?�oA?�兿$qW����k�eg����W?�������b��x��=n���i/=#E�>��=�2�D�3���R�Ë5?�*?��ɾ&[����2>νZT���M,?e�?�y��oU�>��?*��h�=�M�>I�>8�>�'�>V~Z>����؎��:?�]?QD&��Fy����>0���c8��q��=���=�c��i��\>��7<柤��<<�l��\ڼ�0S?C/�>�\,��b,���۾-7�=cn�?�\�>Q��>n�x?=DV?N��=ݾPN������#�z�P?�a?f��=$t(�� ؾh����?�Ug?�!�>[���\U������i��;�?޾w?~�%?�,��x�Z��f��)n(?z�v?ep^�$s������V��6�>W�>���>t�9�|h�>��>?#��H��?����W4��?z�@���?Am;<��0��=28?�Q�>۬O��>ƾ �������q=#�>֍���ev�'���I,��8?���?���>����̨�_P�=�	���c�?�?`X��K�q<2��� l�����T�<��=��c� ����^�7���ƾ��
�U���|��K�>~S@�w齺@�>��7�32�uUϿ��y�о'q�Q�?J�>��ɽ﹣�O�j���t�@NG�ԨH��ٌ�J�>� >��ǽ�ܗ���|��)?���8�m�>h���{>0�]�g"ɾ���:ㅐ>v�>�.�>M����n¾v��?�]��rq˿�E��H�rBU?d�?�P�?�s&?À7�d�}��_��p,2���I?׷p?�Y?��v���~�K� �%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*��+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.���a?�vH�-Dz�e>@�u�&�<KH>�f�۽[�+>=^���[�����U���bM�?(�?��?;σ��V�#�?��><���������Y=v��>2��>a�W>Żg=�ݥ>u�G ��v�>-�?��?��$?��h�/L��]��< �?>)�>
�?{U�=$`�>�P�=I갾�.��[#>K"�=��>�x�?עM?�J�>��=��8��/��XF�$FR���y�C���>)�a?��L?R7b>��Z2��!���ͽ3_1��4��U@���,�8�߽&5>	�=>�(>F�D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���K��V~�����6�!��=��7?>�X�z>E��>��=�jv�����Ҿs�ҵ�>B�?�{�?S��>$�l?xo�$�B�}�1=�G�>��k?j? r���c�B>;�?H�������L�� f?�
@�u@ʛ^?��п�k����������;J>'M>���>�:��褷=&i >���=z��==�E>9*�>�3>@>J�@>�:>�t>j����!�b��"q��'=&��C�u����O�����I��)��~�������,�����ý��-�<����R�2\�=��U?��Q?�p?&s ?��w�">�����$=�#����=��>B]2?��L?K�*?�|�=��h�d�G��h������}��>,'I>�Z�>�>
�>(�k�m�I>��>>=��>�� >�K&=p�.�=�N>��>[��>�7�>�E<>�>6ϴ��1��B�h�9w�� ̽� �?/����J��1��;������m�=Zb.?>K���>п����%2H?K����(�,�+���>��0?FcW?�>Y����T�;>����j�tb>�' �+}l��)��"Q>�l?�g>��t>A�3��h8���P�V�����{>,6?"���6�9�f�u���H�Mnݾ�M>��>E1;��R�c�}�~�l�i�2I{=l:?��?E���������u�l9��SR>��[>W�= ��=�M>�0b���Ž��G�0V-=Z;�=��^>\`?j�+>�&�=zף>de���P��E�>�<B>(,>��??l%?����������@-��`w>�-�>[�>��>ɪJ��M�=�r�>��a>zF�S���v���k@�W>��}�=__�;�u�<�x=�Ř�T��=ar�=�/ �1�<�ɐ$=�~?|~���㈿�뾒`���kD?R)?��=��F<�"�N����F����?U�@-m�?�	�~�V��?�@�?���9��=�}�>wګ>0ξW�L�o�?�ƽ2ˢ�h�	��)#�MR�?�
�?��/�nɋ�Tl�8>�^%?�Ӿoh�>w�zZ�������u���#=N��>/9H?SV����O�>�:w
??�^�̩����ȿD|v����>8�?~��?*�m�{A���@�"��>-��?�gY?pi>lg۾2_Z�]��>�@?�R?W�>�9��'�+�?�޶?���?UI>���?�s?�k�>�0x��Z/��6������p=�[;�d�>�W>d���xgF��ד��h��v�j������a>��$=-�>HE�V4���9�=��
I����f�:��>�,q>�I>W�>t� ?�a�>|��>�x=�n��Lှ������K?m��?���5n�}Y�<γ�=��^�R
?�<4?�T]��ϾQ��>¯\?@ɀ?[?Nw�>��L8��ӿ�����ܗ<��K>��>$/�>�D��0K>�վ�GD��]�>�ۗ>Bʣ��?ھ�f����S�>dm!?]��>�U�=�� ?�.?��G>�	�>��O�L喿}R>����>e�>"?_G�?�?����/��؏�`���	W��|{>rIs?��?�H�>8M��?����� �����<e�? �]?,ꩼ�	?�J�?�dJ?�UF?�X(>R?Y����-���}>n�%?BY���C�b�)���Н�>r�>���>�u�;�-����<����\�?��a?�?/?�]���`�B+����h<G�z��Ϛ<q�0=y==>�>>oT8>
����_�=��#>]��=��@��d�"r=�m�=�č>���=et>�Hc9��@,?%WD����%�=7�r��D�� >��K>���z^?��=�+|����/n����T����?��?�e�?�ٵ��yh���<?R��?�?.�>�-����޾'Mྞ?v���x� z��c>2��>
�b�����m������sQ���|Ž��{�.?[o�>n�?P�?[��><��>�z����)� ﾊ��/�T����w�D�>n<�s&�jC���p����>�[o���$��}�>�1�����>��?&5>9��>}P�>��<Pf%>�I$>��D>�h�>T�b>Y�>U�>��<MSn�LR?�����'�;������2B?pd?u0�>�i�ԉ��r���?$��?�s�?1Bv>�|h��,+�>m?�?�>���Cq
?�^:=����#�<�T����	D��6'����>�D׽�:��M��nf��i
?.? ���5�̾�@׽O�o=�G�??�(?��)���Q�O�o��W��
S�q��?h��{����$�ɘp�I����[��t.����(�6�%=�x*?��?B^���Ԙ���j��?��f>���>e��>p�>��H>.�	���1���]�@:'�
ă����>�	{?]��>��I?��;?�jP?�EL?˻�>��>Y�� Q�>�F�;o�>���>͕9?�.?T0?��?�W+?x�b>���+"���Fؾ1?0�?�+?2 ?�?E����ý^Q��h�b�e�y�QЁ��`�=[��<CNؽps��EU=o�S>]Y?j�C�8������j>v7?)��>���>C�����c�<% �>��
?�K�>�����|r�;h��P�>��?�#�p�=��)>N��=P����Xº)��=�s��� �=����m�;�i <���=6�=�cr��ꅹ�
�:A�;�Y�<��?��/?�Eb>�>=]������b�>d�[>�*p>�N�>o���*���͔��nK�q�c>���?dخ?��=��=��>Q���о�� �3���
>L[#?"
?��t?\��?^\I?A�'?��=��I�q������[D�H�?�!,?抑>���$�ʾz�j�3�P�?B[?�;a�A��r;)���¾��Խ*�>�Z/��.~����)D��������J}�����?㿝?�A���6�ax�����\��c�C?�!�>�X�>P�>�)��g��%�L2;>ڊ�>�R?/$�>p�O?�;{?d�[?fT>ޜ8�O1���ә�)D3���!>�@?���?��?�y?Mv�>&�>��)��S����������dW=�Z>F��>(�><�>���=uȽuU����>�K]�=E�b>��>d��>��>��w>=�<��F?5�>���$������˛��jl?�Ӎ?�,"?�:=��A�E��{����>�ߥ?4��?}�%?DpJ��v�=����x�������;�>�\�>Y��>�=�=�y=�K/>���>��>������c�?�ݰ��]@?�E?>8�=b�ʿ1�q�����{��J>��I�u����ڽ�Ps���Y>x6ҽ|�8=����Ɇ��Ӿ���щ��(Ţ�(L���k�>|>��T>~<>�0 =Rǵ��w�<O_:'J8������NK�"��������:j˽�ix�4:=�#'���ս;�ѾЈ}?��H?-?A1E?�ˁ>a?&>BW^��Z�>�|��%?��N>Z>���ľkL�!j��1$��{{�8��T�]�M���
>��7���>><>y�=pʤ<�m�=���= tb=����X�=R��=��=\O�=���=�>64>��t?��l�%��V�U���1��;?[�3>o/�=�é�V�&?�$>�}�����1��
�q?���?�?�?U��>	�>�*���ؽ�^.���򡼌�Y>2��< |߽w]�>�]�=f��ۑ��ݼl��?���?��A?�t���Uο��_>��9>@g>BS�)�1��_�te�{n^�!?T":��̾���>%ۭ=́���žiR2=-y9>�Ys=�����[���=�I���W7=��^=�ۊ>�F>Y�=�/���t�=�<=�-�=�4P>Qĺ57%�z�>p>=�=[}]>��(>F��>�Q?v�*?�$Y?=q�>�Xo��6־�����Ì>��=��>���=�,>ܮ>��;?خC?^K?bo�>���={Ů>MA�>�G'��o�_��
���3s�<ms�?E��?N��>���=�<"�7��4;L���*��?�0?5�?黐>$T�%��[&���.�8И��b9ƹ,=�gr�ܸU�;��c��Y�+�=NE�>3��>���>s.y>��9>��N>��>��>���<yÅ=Ê��j��<�X��9��=�:��)g�<.�Ǽ�簺��$���+�ו����;h��;�Z<�d�;k��=���>�a>Գ�>�v�=a����R/>?Ԗ���L��ɿ=G��3)B�q#d�(G~�T/�1�6��FB>��W>�h���(����?M�Y>�?>6��?�:u?��>�,�s�վ�S����e�C�S�59�=@�>!�<�:q;��R`���M�̒Ҿ���>fߎ>r�>�l>�,��"?��w=A�Nb5�O�>�|�����(��9q�&@�������i���ӺߟD?VF�����=Q"~?+�I?p�?���>���ʆؾX:0>�I����=���+q��j����?�'?H��>f���D��;̾hƿ�,�>��H���O�(���5�0���#�n��~�>���>�о:3��a��y��B�r��A�>+�O?��?�a�B[���-O�����a���7?�Hg?e̟>�??&J?;������錀��F�=S�n?%��?F3�?m�
>蛽=52��_@�>�,	?���?��?��s?�y?��x�>�U�;ޫ >�����K�=��>ey�=3�=�p?u�
?��
?�\����	������^����<=ء=��>�h�>2�r>���=�g=��=]0\>Uڞ>��>��d>!
�>�V�>P�8�*��YD?���>0��>2K?��>�A&=��d�Nm��ޞ���H��1�R�.�R�u�>�Y�O<�{Ľ<8/�d��>��ʿe:�?΄F>v���F?����MOR�ɎD>oP>���̪�>33X>��>���>=��>}�>���><��>�FӾ>����d!��,C�0�R�P�Ѿx}z>�����	&����w��4BI��n���g��j�K.��R<=��Ƚ<#H�?������k��)�����R�?�[�>�6?jڌ���ӯ>���>�Ǎ>�J��V���Pȍ��gᾢ�?<��?Ƨ�>͏>\�1?��-?�ak�Qkn���4�9�z��e��6�3C�?0���艿�!�z�O��.I?F%�?��m?��R� ��>��h?Nll�#����<��Z��e�u�=� �>Cƾ3����������Ph>&f�?���?-�>3�;%�m��'>��:?̛1?�Ot?��1?i�;?�����$?ao3>�F?�q?7N5?��.?'�
?T2>
�=�����'=�6���Q�ѽ�~ʽt��V�3=�^{=a�͸@ <�=���<&��ټ{�;�%��	%�<:=v�=�=�ئ>�]?��>�S�>��7?w���8�����"/?\S8=ł������袾T���>�j?���?�BZ?&Vd>�A���B�4�>���>�V&>�U[>�M�>���;E����=��>��>L��=�P�`1��g�	�:h��y��<��>�n?ך>k�̽�n.>ф��z7<�?Aa=2_��O`��ut�s�(�����;0�c>?��h?m�$?��[=9v��5=
�d���"?��5?�b"?��L?�ջB����<��z;�������>�==l��^��h���D8��W >��>7���0࠾>b>͸��_޾��n�<J����hRM=Jx�y�V=���־n9�.y�=�	
>������ ����Ԫ�W-J?��j=�t��Y`U�l����>���>�ޮ>Xh:��Iw�=�@������;�=���>�:>h���ﾡG�i7�j>�>TQE?@W_?k�?"��[s�;�B�y���dc��wȼG�?px�>$h?�B>h��=M�������d��G���>���>c��D�G��;���0��D�$���>S9?�>��?]�R?�
?y�`?�*?GE?''�>�������B&?5��?��=A�Խ��T�b�8��F�� �>Y�)?��B�͸�>Չ?��?�&?ǅQ?0�?a�>� �4B@���>[�>,�W�"b���_>��J?���>�=Y?Ճ?��=>��5�颾Rة��J�=s>��2?�4#?��?U��>��>����k��=?O�>�b?jЂ?��p?��=y�?��4>�2�>F}�=Z�>]�>o?��N?��s?JJ?���>n3�<䳭��r���t��\*��� < a<��p=��"�x����;P�<�_�;{����m��2ܼ@�����՞;��?�4�>Ӥ����<�|���K����:^sM��1�)d��$�~�e4�=Er>p#?��>�"ȽKC�=�>[C�>Ǟ���)?�G?g��>Y�>7-��#��\�)M>�?���<�΀�2���C����=��x?�x�?X��0���d?!�h?����J��I޾|P��پ��r?�?������>�H~?�Jb?z��>�b��{g����ݚh�<,��5�'=��>����Qd���>ϛ)?2�>�v0>�T>����5q�T���?�?ƈ?�l�?xZ�?�}C=o�x�Qm�j�꾷2���9�?W��>f���18F?�>�S������k����r���m��E詾���о�;\��8��Jv���U>G�-?H�t?+!\?��?u?�C{�J�>�Bs��s���i�"��5�ٌK�#�?��T�v��������kA=�̃�D����?In(?E�q?eҋ�<Q�%ȾRr8>����V!����=I�����<�$@=A&r��:�OU��J ?�&�>G�>�./?0�a��`8�^W%��1���� �'> >�>��>f��>=)��#B.��S�.�˾�o�<�_���u>�c?\K?�n?�z���u1�6���~ �N&��:��`�C>g>� �>d<X�����4&�|S>�<s����ސ��	��u�=3?�i�>l��>祘?�?T	�^a����u��70�J��<��>�i?���>��>��ʽ! �u��>��l?9��>���>뉌�]!���{�U�ɽT*�>	�>��>p>ͫ,��\��f��g���V9�|�=�h?�����`�k݅>�R?i��:U�I<0��>)�v�©!����ʚ'�d$>E}?;��=��;>vž�'��{��5��GC)?L?�ڒ�Š*�P6~>A"?1��>&�> -�?F9�>�Mþ�.���?}�^?L3J?LA?�U�>G�=A���B<Ƚn�&�f�,=��>�Z>��m=��=7����\������E=䀺=�μK.��H2<�����K<	�<l�3>mۿ�EK�a�پ��T��;
��ꈾ_ǲ�Z����p[��H���Rx���'��V��1c�������l����?H:�?k|��!������j�������@��>��q����C쫾����'��h��X���Rc!�v�O�z$i���e�ɗ'?�?�ǿ���:ܾ� ?H< ?��y?H�͡"�ř8��� >-+�<]#�����J�����ο������^?L��>���"�����>���>i�X>Qq>c��(䞾q$�<b�?��-?x��>wpr��ɿ5���r��<M��?B�@"}A?��(���쾴V=���>�	?��?>HS1��I������T�>p<�?��?�}M=k�W���	��e?��<��F���ݻ$�=";�='E=�����J>|U�>܂�^SA��?ܽo�4>Yڅ>N~"�S���^����<0�]>��ս<��,Մ?ez\��f���/��T���U>��T?y*�>m3�=ʲ,?n7H�6}ϿE�\�m*a?�0�?Ѧ�?�(?-ۿ��ؚ>K�ܾ��M?aD6?T��>6e&���t�S��=���"��}��t&V�%��=Ԫ�>�>R�,����6�O�eJ��$��=�����xǿ֬%��HѾl�Ƽ�`t=:��v*f���=z�Ƽ�i^���C�떽�-�<q��=��D>�/�>���>5�*>/ka?P�I?���>�̧>�󕼾�c�Z�ݾTco�E�ھ"�/�|��;}�V���d�㾺⾙��v�[
����v<�u�=:R�7����%!�|b��UF�n�/?y^$>RɾHM�{C<g/ʾ�誾-n�������˾�1�w�m�3��? �A?���W��u���5���yW?:i �X�5{����=�ݤ�O�=�>�=�2侯q3���S�QB0?Sl?�,���-����*>�h��=��+?��?�A^<$�>[r%?�*��佉wZ>�D3>Yգ>B`�>�>�(��Xܽ�v?��T?���t.�����> h��+z�3^=�>�4���꼅D[>��<�挾��V��p���P�<�XY?��>+�2?"������$��q%=^p�?|?5�>��g?�GD?�)}<�\���QN�K����=�!I?�{c?���=��������t6?(i_?��_>8R�"&���;�ξ��\u?irp?��?��꼲4v������y ?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=6ޕ��^�?|�?a����h<���l�;|��YV�<�=Kb���"����<�7���ƾ�
�_���<��E��>�Z@���>�58�o7�/VϿJ��Cqо	dq���?�g�>��Ƚߟ����j��9u�x�G�r�H�����ΰ�>�i>����UJ��b�{� i;�������>��
�Wڈ>�2T��p��3$����*<!��>�$�>�@�>�6���˽�v��?N����Sοơ���o��HX?*)�?B`�?f�?��"<�w�^;{���JDG?�s?Z?s�*��;^��:���j?W[��dV`���4�<JE�YU>? 3?�?�>Y�-�LZ|=�>���>��>K/�K�Ŀ�ض�����?��?���?Xn���>���?�s+?�h��7��"_��N�*�`�5��=A?2>�����!��/=��͒���
?3~0?���<+�;Uw?҉1�����7�:���M~���Qؾ�����Ǌ��o����(��g3e�x�?��@,g�?�q����#?��>�U���&ʾs��<<u�>��>�&d>��Ӽ�b>��޾��S����>��?�� @r�=?fș�e4���R�>gq�?G�>�
�?�ʸg�:>O-9>�I쾝�����>�Ez>x�;~��>�jJ?U��>@'t�=�PS�1*A�1�|��.��tH��J>��r?64�?F�>c�H��l��]8�j�ܼh뽏Z==��V�q�Y�mm�����=�
�=2T�=Y$�����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Qz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ca~�1��}7����=��7?�0���z>���>J�=�nv�ۻ��Z�s����>�B�?�{�?��>4�l?N�o�k�B���1=7M�>��k?�s?Jlo����B>_�?1������L��f?	�
@}u@L�^?+u�׿#��BS���I��Ϣ�=
�>>��s>�!���i>+=9>��&=	�[=%��=B�h>v�U>�I�>�5>�D]>�j.>��~��(�L���lb�F}k�j��4A����.���~�N1��a���ǫ�&���Cg��e��:=�I���6q\�f�=t[X?��P?snk?w�?����/ >���==����`�=xd�>)n.?�F?��%?4uv=!&���fe�=���<��@H����>��S>?��>S��>d!�>-��s�F>eB>���>�Z>�t;='d;�oO=��Q>H��>�J�>mһ>�C<>4�>Dϴ��1��g�h��
w��̽@�?X���5�J��1��n9�������h�=4b.?�{>���?пa����2H?���q)���+��>_�0?�cW?��>���!�T��9>;����j�K`>�+ �Tl���)�%%Q>Bl?Fh>LOz>��3�+9�KP���S�y>�7?�ϴ���8���t�pG���ܾ�K>�<�>+3K��p�oS��*���pl��w=�;?M�?�᧽=���D�w������R>k>[> B=�֩=J
K>L4d��ʽ>�G��..=��=�s]>T?�t,>�=�=,}�>t����P�~��>��A>��,>�@?tD%?��u����p��f.�ĸv>���>�>�B>U-J�~'�=0�>�Ea>r��n��
��}@�s	V>�9�� �]��Gt�)�w=�5��3��=I��=k ��$=�`�"=��?qmt�7���������ߺ>�>A����a�ʜ\�������r�&V�?��@�X�?�C��}���d?0��?�Y����)>�5�>��E>�^�����=�E?��/=qW�T����m>���?s�?�β=մ��,����>W�9?|�ɾQh�>yx��Z�������u�w�#=R��>�8H?�V����O�e>��v
?�?�^�੤���ȿ5|v����>X�?���?g�m��A���@����>;��?�gY?soi>�g۾?`Z����>һ@?�R?�>�9��'���?�޶?կ�?_I>���?�s?�k�>l0x��Z/��6������cp=��[;�d�>�W>d���vgF��ד��h��t�j������a>i�$=#�>$E�G4���9�=���H��	�f�9��>�,q>/�I>&W�>u� ?�a�>���>�x=�n��?ှ�����qK?���?���l�s��b<ʑ=B�b�V�?�;4?Y�r�;�ʾ��>�U?��v?"LR?�Ѝ>���Eʝ�N���������<6NY>��>��>�Vɽ��+>���	,�7�e>���>�	�j�ؾnz��{��v9�>��?%�>:C=��#?�(?`#V><�>�LM�s���6hB�0,�>8/�>g?�+z?Z�?ɾ���3�zd������N���:>�u?_�?QD�>����\��[���G��$#��	�?�Ip?���?+��?�C?BgA?PUL>�!�&��������V>g�!?v���A��M&�;�d~?Q?���>�7��@�ս�Aּ��������?�(\?cA&?����+a���¾|8�<��"���U���;�xD���>Ŏ>����Ҍ�=`>hذ=eOm��F6���f<Ak�=��>��=�.7�Cw��?=,??�G�,ۃ���=��r��wD�X�>KL>z��߬^?�l=���{�����x��QU�� �? ��?3k�?�����h��$=?��?	?X!�>K��f}޾m��zNw�l|x�w�Y�>���>�l�U�B�������rF����Žc�$��(�>��>�?xx?�U>tl�>֠��Č#���$�V�^��`��X8�+6/�{�����J7&��>�ܸ����v�/��>����l�>7??H�h>,*~>���>:#����>QW>h�> ��>e�V>��8>��>	�*<�ѽ���b?�1��)_4����龀t?�:?ͻ>��-�����R
���&?l��?߬?��>n�j��i7�EP@?ii ?������>�>vɐ=��]=c7���[����G���.���>����e:��il�/8��#�??�B�=�n��������un=�N�?��(?��)���Q���o�\�W�S�t���(h��u��2�$�#�p�/쏿I]���#���(�m>*=Ȋ*?b�?��}���4%k�{?� bf>���>�>ξ>�wI>��	�E�1�Y�]�BF'�ݲ��OR�>8T{?��>�~I?��;?�P?�JL?�m�>�f�>�߯��y�>�\ <~s�>�F�>Q9?(�-?r�/?#??/t+?f�b>�x�����"�ؾ��?Tw?�-?V'?��?&���XĽ�s���oP���x��`���K�=�d�<2�ս3�s�ۛS=[S>5k"?����G?��R��ZB>r@-?fQ�>I��>���料�����^�>�#?���>�5꾊�t�`����?�?���1�\<S5>��=}.]��Y���=E�2�=�!�;N]�Wq�<\�=D�5=_%��l<��Z<�-P<'Z�;Â?/x,?g�>X�	>R�ľ��Ҝ�GG�>܏�=�S�>�r�=QZž���mo����L�^AY><��?W�?�%�=
�>UhR>��Ⱦ�ɾ	���žno>>i3?H�K?�G?�ښ?�W?-?��=��'������@��ڤ��\c?#,?���>�����ʾ}ӌ3�͕?\?6a�����9)�K�¾��Խ��>,V/�`,~���� D�4J��,�����*��?W��?��@�M�6��{辠���qZ��J�C?>$�>JS�>��>��)��g�� ��5;>$��>	R?�#�>��O?�<{?��[?�hT>��8�M1���ә��83���!>3@?��?��?'y?Ut�>��>��)�)ྷT�����X������W=	Z>ߒ�>�)�>�>���=� Ƚ�Y����>�Sa�=�b>���>���>��>��w>wP�<1�I?��>⣾M��Zd��rR��y �Uuq?>
s?n�9?����!�UR�'=�����>�ӣ?��?~i?o+=����=]�O=SD��xin�IT>���>���>��>9>ZN�>��>M4�>��+�gT1��K���ɽ�H?}W:?�(�=Lб��'����M�F��>��@>Ϲm�=i���Ě��dW=�>�/=t-�4䦾�ۥ����Bk��jׯ�#��)�	�ݘ?�h>ȸm>��L>���=@��T=� >3�H=�[����������x�쫈�4L��[�3躽��Խj"ý_�ľ��"?��4?]�?O�b?�N>��>�>
I?�m�=],?��>m=��eľ�漾�E��s�9�����aľ��.�����=l�=����)�=�b�>�>t2��C���t^
>�7�=�Z��\:=���=z��=��=�7>�c>�*>j{?N�i�@ϝ�/Q�PeC�9
?R&>�_j<���&�?���=Hp��f}��l��dy?D@���?$%�>vf��̈́�>� ���y�(��9�Ϛ�ս/=y���}w轸��>7�=�k&�.������b�?[�@�<P?�����ʿ|D->��7>+>r�R���1�[�\��b�^Z���!?E;��?̾>�>y�=")߾�ƾ�l.=��6>T�b=d�mS\�'��=,�z�H�;=j�k=�ډ>�C>%~�=MG��)̶=��I=���=��O>@>��"�7��,�t�3=���=>�b>��%>@��>Ӆ?��+?�mS?缴>��R���ܾ[�����P>��	>� �>J= =��>aB�>�==?hTG?dZ?…>,̍=N��>(Ƴ>a���cg�����'���<�<�ē?S�?#��>�s<��D���#��}Q�����	?�P9?ۭ?�>����߿ n'�y�#���ƽUJz<b��<������h:6�L�G��~Ľ݂�=�U�>h��>0��>��q>6�V>��J>�>&��=�[<2>�~�F�<�O_���S=f4�ѐn;���Uz���;tL/�îԼh���<���<A�����=f��>�;>F��>\��=���OD/>
�����L�ÿ=zG��,B��4d�kI~�8/��V6���B>�:X>9}��'4����?P�Y>+l?>���?FAu?��>~ ��վ�Q��]Ce�gUS�T̸=��>m�<��z;�[`���M��|ҾD��>�ߎ>Z �>#�l>�,�g$?�x�w=q��d5��>G~��ʩ�n��0q�<�������i���ɺ�D?�E��f��=9"~?ȮI?6�?b��>�3��ŋؾ�#0>�;����=?�?Cq�Č��?_'?���>�#�l�D�-JǾ�Vͽ9��>l�G���S�,����#+�_��lT��i��>�7����Ҿ&*4��x����߂@��i�Ǽ>GO?֤�?�6��Ⴟ�>Q����)Ž�b�>h�^?���>K=?���>=wĽ�����ڂ����=��q?�*�?�J�?���=v��=��.��>�8?��?r�?L�n?��=� _�>��;�/(>����O��=ͣ�=�ia=?��=�
?rw?� ??�������B�~����e��wy�=�>�=ʧ�>O�}>�3j>yX�=6�_=G}�=:�a>h9�>��>��a>�Q�>��>�趾�=��u.?��R>��~>��S?>#�>Y#=^s��{��<Gڠ��-x�С��(	��9���=v@������X�n����>L���cԐ?�|=��3���,?����)tN�ݶw=:�>6�6�O�>�C>3l�>BT�>9��>�2{=��i>Zn�>GӾRt> ���a!�C-C�^|R� �Ѿz|z>����	&�P���~���?I�:n���g��	j��-���;=����<�G�?�����k��)�������?�^�>r6?��������>g��>`č>HI��X����Ǎ�ph�6�?���?W��>���>V~Z?�3�>~����+���E�8oy���_�@�[���c�����拿��y� �Bc?���?�&/?�&�<o�>,�?Slv�1oվ�>5�S���x�Ό���V>U����u¾������N-����>�.�?^��?�d�>�ѿ�;�
�� �>d* ?���>m?��"?��?�\ὄ�?k�>p�!?\y?��? ��>��>e&>�o�>����,�t<�H��X���+Q��ܚF���9���=�3>V����ۼ!�:���=�<��ٻI���~8����=8��=���=2��=m��>H�]?DJ�>��>B�7?.���h8�d���e+/?�:=c�������Ţ���>e�j?���?�_Z?z]d>>�A��C�7>W�>r&>�\>j`�>0��ЗE����=�f>V>S��=�aM�ҁ���	�������<�>h��>�i}>P]����#>4⡾Nvx���_>��U�Zͽ�y�Q���G���1��|w���>A�L?�$?5�=V�t~��.�e��n)?΋<?�8L?��~?��=r۾m7���I�����y�>Iχ<�+
������ء��|9�I�<xo>?k��-�Ӿ���>����о0�f�O�<���¾fϼU��L=ѽ0�-�CV ���w�!TB=��$=��g+/�~A���%��PhD?}��=����E�ڥ�n�W>yɸ>�_�>Q� ��顽
�C��/����@=�j�>ž\>�
�<�"ݾY5>�US��?�>QE?V_?�i�?����s���B�����`���Ǽ��?�z�>�h?�B>d�=��������d��G���>���>�����G�sB��4/��x�$����>O;?f�>��?�R?m�
?��`?�*?C?�"�>"��X����B&?y��?���=� ս��T��9��F�I�>;�)?��B�p��>��?(�?��&?u�Q?ܮ?��>#� �%C@�S��>`�> �W�`���_>��J?���>6Y?V҃?�=>`5��ꢾꩽ/h�=6>��2?k4#?��?���>���>H���S�=]��>�c?�0�?3�o?ԃ�=+�?g92>?��>���=雟>D��>�?XO?�s?��J?���>g��<�6��_8���Es��O�ς;�uH<��y=�l6t��J����<l �;�d���L�����N�D��������;K^�>(�s>Q��+�0>��ľ2Q��l�@>8W��ZK���ڊ�(z:���=���>�?>��>9]#�ʯ�=n��>I�>����4(? �?1?=�#;Ҡb�:�ھ޹K���>eB?���=��l�ԁ��0�u��g=\�m?_�^?��W�� ��4�`?0�a?��_�B�i߾�i��n$�$2m?��?�� ���>+�x?�>r?j_?G�=���l��}���U��1��e�=ֻ>7$��QY�P�>��B?��?�#4>�>�����]�1����>
[�?�f�?���?�#>�\c���׿����&��4p? �?#���Wz>?\�#�����`���򍾌� �㡦�m���h��<�ľ��W��ɣ��,&����=��??GJ?#�T? X?���k؃���p�.�f��;O���Ͼ$�G�[��7��eI�˄P�Z�¾<��o?�S�A>����@��a�?5S3?�"���?'�_�y� �P�=Q夾/,���=q�
�����|����&�f�9*���^6?!�>m��>�*@?�\�gK<�c�D�P�3�����G�>��h>Yaq>���>
q=�b
���˽	ξ�{j����<6&v>hyc?ʎK?��n?�e��(1������!�EM/�9`��x�B>�{>^ǉ>4�W�\��9&�IX>���r����k���m�	���~=w�2?,�>���>3N�?��?x	��n��wkx���1�{�<�(�>^i?�<�>��>�н&� ����>��l?_��>��>N����[!�t�{��ʽg%�>��>F��>�o>��,�V!\�4j��Ѓ���9�>z�=[�h?'�����`�L�>�R?_��:P�G<[y�>b�v��!�_���'�m�>�}?R��=��;>��ž�%�6�{�?:��P)?VL?K꒾�*��.~>�#"?��>�0�>K1�?3+�>"oþP�B���?T�^?�AJ?*SA?H�>}�=���,CȽ��&���,=*��>��Z>&.m=���=����s\�o��.�D=�r�=ŵμMP��e�<Uw���K<q��<��3>@mۿ�BK�t�پ�S�w?
��爾e����c��ݲ��a��6��ZXx� ��N'�kV�k7c������l�Ї�?�=�?"���q0�� ���=����������>~�q���������j)����n���ed!���O��&i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >`C�< -����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾g1�<��?7�-?��>Ŏr�1�ɿc����¤<���?0�@�|A?U�(��쾎	V=:��>�	?��?>�R1��J�����SS�>�;�?��?�uM=��W�R�	��e?�<��F�0޻� �=GA�=�E='��ŏJ>�R�>:x�)PA��9ܽN�4>^݅>;n"�i��2�^��(�<��]>��ս#7�����?wo�1�d���S�Ӻ��=v>.�;?��>��`>a�??lO���ο�Dl��i?�U@���?x�?�}پ>5�>��ξ52?Z�E?>Ѿ)O�~h9�钮�n���`��;��z>E"?r2>�6�;���ő�G�Խ
��e�D�ƿ#�$� }�
_={�ݺ'�[��}罨���G�T�d#��)fo���轉�h=���=��Q>Kl�>U%W>4Z>gW?��k?�N�>C�>�6�h���ξgy��G�����G�����p��R�ԩ߾}�	���������ɾ� =�}�=�5R�◐�� ���b��F���.?�w$>D�ʾ��M��z-<}mʾ_����������0̾��1��"n�a̟?��A?������V�����8�o����W? L�n���鬾��=�����=�%�>[��=��3 3��~S���/?G6?���'���{�&>�9��	=
�+? �?8�><�G�>d�%?�(��3޽X�Y>b�0>��>�Y�>c�	>�簾��۽��?�ZT?,]��yg�����>ܢ��`Pz��5a=��>��4����EZ>�jj<�W���Z8������<�(W?��>�)����a��	�:S===�x?��?�.�>{k?7�B?ɤ<�g����S�(��mw=L�W?�)i?��>���
о����R�5?ۣe?�N>�ah������.��T�$?��n?�_?�m���u}�������n6?�w?tb^�aN��xv �gmU�2Q�>���>=��>v`8���>��<?��)�'����I��B?2�2G�?��@�>�?S}X<� ��<�=E��>���>�K�����b��:B��!э=���>���s�� �#����9?z�?�+�>�2��J������=�ٕ��Z�?N�?f����<g<w���l�o��"��<5Ϋ=��qG"�����7�B�ƾZ�
�~����ݿ�L��>*Z@BT�D*�>fC8�@6�TϿ���z[о�Rq���?�>\�Ƚc�����j��Pu�h�G���H�s�����><��=CZϽ��y��yt��B?�\v���>�7�7�>� I�U��`���1>�D4�>�K�>�D�>��;���H�?�i��Ϳ�������bU?�?�?���?��$?2?=T=L�z'n���>��N?�u?k�[?�wg��W�u�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�b�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.���_?��a�}q��_.�$uϽ\b�>[�.�S�\�Y���,��Ke�9.��K�|��ح?�f�?�O�?�O�"�K�%??J�>����&^ž��<���>At�>t�K>�b�iMu>�����:�bv	>C��?��?��?/.��������>�3}?�E�>��?;-�\�3>q}ļ1Sξ��t�턀>�s�>��u�+�+?�aS?�h
?�ɠ>��J�s�$�	)��T��1˾ ca���">JNh?� c?!ԧ>>�_�"��6(0�������W��3E������t=[�����<��%>�?�=�Yh���Ѿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji���?����ۄ���a�C0��o��=�2?�`��i�_>���>K=D!z�e��1�n��y�>�ߴ?���?���>u�q?��^��O�z�ܼ}Ŭ>��^?��?���=(�¾�tZ>d?���(+��ח޾_4g?Tt@3�@��\?����hֿ����ZN��B���y��=���=��2>��ٽQ_�=��7=\�8�=<��)��=r�>��d> q>(O>sa;>�)>���K�!�r��]���I�C�������Z�B��1Xv�Xz��3�������?���3ý�x���Q��1&�??`�i=�Y?a�Q?��k?Y
?G��jW>đ���H>!�1��G�=�T�>^=A?CO?*?Q��<3���4�^�~o��^��ǀ� ~�>��{>�}�>���>T��>eiʽ�Q>=y2>1�> �>E<GŽ��&;E:>W2�>b�>���>D<>��>?ϴ��1����h�cw�̽C�?������J��1��I9��\���qj�=6b.?S{>����>пV���l2H?�����)��+���>��0?�cW?k�>
����T��:>i���j�e`>n+ ��~l�r�)�t%Q>>l?߾f>Gu>��3�me8�u�P��{��Ll|>�36?J趾%G9���u�<�H�LbݾWHM>�þ>p<D�[l�f���m�	wi��{=�w:?o�?h4��@ా|�u�[D��fOR>�4\>�b=2l�=�UM>xec��ƽ�
H��l.=���=��^>�Q?�,,>�@�=��>7m��eP��{�>�B>7B,>�@?	:%?�������f����-�"�v>�<�>Y�>m>s�J��ͯ=�~�>Bb>��X�#��I�?��hW>�}���_�>�u��
y=����t�=��=�q ��=��	&= �~?���䈿�4e���lD?+?��=5�F<`�"�7 ���H���?f�@,m�?(�	���V���?�@�?��]��=h}�>�׫>�ξ�L���?_�ŽȢ�ٔ	�>(#�vS�?��?p�/�]ʋ�`l��6>�^%?`�ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?�I>���?�s?�k�>�.x��Z/��6��ږ���o=@�[;
e�>X>:���ugF��ד��h��m�j�o��	�a>�$=K�>VF�_4���7�=n��H����f����>O-q>��I>=W�>�� ?b�>Y��>�u=�o��pှ�����J?�H�?>�$�p�_�P��F=C%9��R?A�6?i9<f���X��>P�Z?���?� T?��r>e��^���{��^þ2j=�4->���>ҙ�>�s����w>���
�J��"�=l8�>�@żx���|�#j����>1�?C�>�ȸ=�! ?�� ?��>��m>�1������<b�p	?�s�>]�(?=gz?Ъ?��~�6�)��h���V��D�Z��`>f�k?�{?>�>����B��%�l�D���:��;V�?N�?��;�j
?�q�?`�O?+�N?"6Y>P~����G��U�=��!?���A�uN&���(~?�P?���>�1���ս+Lּ������N ?C)\?�A&?Ɯ��+a���¾�0�<��"�բU����;@�D�*�>��>V���.��=V>4ְ=�Om��D6���f<&o�=��>���=�/7� w���<,?F�G�W��Ø=��r�SuD�F�>�AL>�����^?k=�d�{�^��Ut���T�r��?���?<i�?�촽u�h�r$=?z�?�?� �>�T��m�޾:f�3w�bx��h��>k��>��p��5�P�������x=�� �Ž�,��I�?|��>�?��>.�e>D��>�|��2�"�%��Dp&��9h�ʹ��u;�^7�Ŵ$���¾�4��z.V�yW��X���>PAj�4�>�G?�z�>�|`>\B�>+���(�>9|�>�F>�_�>��y>F4\>/�	>t��<��콢KR?[���~�'�8��/���0B?�pd?�8�>��h����k����?��?s�?f>v>e~h�1-+�\l?�8�>����q
?�A:=G]���<�M��g��DH��h�E��>S*׽:�rM��lf�sh
?b/?�䍼*�̾7׽ӂ��n�l=�Q�?)?��)���Q��o�W�W��3S��5��h�-z���$��p�鏿�T�����׌(�&+=��*?��?ŗ�ix� 4��KLk��%?��vf>�	�>�>�Ծ>h�H>]�	���1���]��'��S�����>�F{?�!�>s�I?<?�mP?�XL?��>��>6-��7��>	��;�>>>�>��9?r
.?(0?FB?�0+?ib>�9��^6���aؾ�	?�?<?�1?4�?�2��@�ý.���SXa��Dy�>����=~�<#�׽!�u�QT=UaS>�X?���Ƭ8�����ak>i�7?��>y��>���,-����<��>�
?	G�>E �!~r�c��V�>���?���Z�=��)>���=����L�Һ4Z�=������=�6�� z;�jf<p��=[��=Ot��!��!>�:ן�;fn�<�I ?#m?ϱ�>��b>p���%�ɛ�>��=@�v>D�>����΁�%m���vZ���\>��?h*�?���=>�=�r">g鞾����	�x(ؾ�䵼�!?��1?:5S??F�?G�K?-�0?D�{=G#*�@/���K���ᖾ��?d!,?~��>����ʾ�񨿾�3�ԝ?t[?M<a�S��0;)�`�¾ �Խ)�>�[/�Q/~����D�}녻���3����?ٿ�?A�E�6��x�ؿ���[��@�C?"�>Y�>X�>H�)���g�V%��1;>��>tR?�#�>��O?�<{?̦[?�gT>s�8�}1���ә��D3���!>@@?��?�?}y?�t�>��>�)��ྖT�����9�=ႾdW=&	Z>e��>�(�>I�>��=�Ƚ�Z����>��`�=�b>S��>���>��>/�w>�L�<�H?�0�>���%��^���넾��H�A�u?��?@+?&=M���XF������q�>�A�?S�?Io+?5�S��@�=(м�J��`Eu�5F�>���>a�>���=$(R=�>���>K�>,y�����=7���B��-?|{E?���=}�ſfeq�j�p�f����}�<x�����b�^b��� Z��;�=�2��F��4慨[5[�����F���`Ե�r_��_�{�#-�>#�=��=G;�=*b�<h�ż���<aRJ=���<��	=��q��ȃ<:�$eǻϟ������s<OK=J��)�쾪ni?s??�&-?�mC?3Mo>[~c>ߓ�{�>�,��Of?��>��`=�C��I�S�i����G��:|;�Kʾf�~��;��ׯ�=��y�آ#>[ >Ʀ>_
I=���=�J�;�()=gE�
����=±�=~y=��=�>��>�#�?%Vl� ���ե8������>���>\e>PEe�L�7?m��=Wm����Ŀ�wܾʿk?���?���?X�$?�V�=�+�>�i��<ʮ��������lȸ>�k�>�΢�g=�>fN�>R'��M��+�J�WZ�?F �?\�M?/o��K�Ͽ&��>|�7>L'>��R�C�1���\�˚b�~qZ�Z�!?�F;��K̾v:�>q�=�'߾4�ƾ��.=��6>-Yb=f�3U\�י=��z�-�;=��k=׉>A�C>nu�=�=��)�=�wI=���=��O>�p��|�7��C,���3=3��=u�b> &>C��>i�?k0?@6d?}�>!)n�jEϾ7+����>�y�=f+�>@��=�,B>�i�>��7?Q�D?��K?靲>���=4Ӻ>I$�>Vx,���m��@��觾i��<���?iȆ?�ڸ>B�X<R�@��{�B�>�,3ǽ+?�+1?Gv?��>�T�ğ��V&�y�.�i]��r���W+=�hr��=U�Z���e�ƃ�j!�=�o�>j��>���>Py>B�9>ϿN>��>x�>�J�<-[�=<2���۵<�������=d���}��<�|ż<���4�&���+��Ʀ�a�;&]�;��]<��;v��=���>�N>��>ϖ=���)+/>B���!�L�Pӿ=8F��)B�n2d�F~�� /��L6��B>�DX>*n��>3����?��Y>�j?>ނ�?�8u?B�> ��]�վ�M���,e��4S���=�>�+=���;��Z`�=�M�BuҾ���>��>��>0�l>�,�i#?���w=��a5�h�>�{��,���'�9q��?������&i�(hҺ̠D?�F����=�"~?]�I?H�?���>M��Ԇؾ�;0>uH��F�=Y��(q�Rg����?�'?t��>���D��`��J�`�T�>!R=�U��Y����K�47�����d�>g�Ͼ���'�kᖿ;͊�0r"��#�����>�0>?��?�#��䌿c�C�i���������>�Xs?��>��>c�?Ξ@�5�.��������=T�|?�g�?�(�?�{=Mw�=!��#6�>K)	?���?]��?��s?�w?�Wz�>�҉;c� >y����b�=��>Yw�=m�='o?o�
?�
?kt���	�����^�x��<�ѡ=׃�>�g�>��r>���=L�g='i�=o+\>CԞ>��>`�d>��>�L�>�_�[Nᾏp5?�ZS>Ta�>M�_?��>j�ռl�j�'��p����.�
�)��_��_`��fr��P������?��ҿCы?c�>\�
��
?���,�j�v=^�>}`�y2�>��>�Ԗ>�F�>��p>	T�=(�l>��>�FӾ}>����d!�l,C��R�]�Ѿ}z>����
&����w��oBI��n��lg�nj�6.��<<=�	Ƚ<H�?������k���)�����+�?J[�>�6?rڌ� 
��:�>��> ȍ>�J��l���bȍ�hᾗ�?%��?�Md>t��>}?W?8?�*3�`�5�b
[��Pu�7sA�ܥd�v�`��΍����N����ýit_?�Iy?TTB?b��<J�}>7��?T�&�����È�>�J/�r�:���O=���>h=��w3\�a�Ӿ ƾ����`G>��o?ܚ�?�?�~W��M�����=��?A6?VTy?`?�J?�I�kE?��=�?5)?�>?�?-��>Dnh��㍼GE�n�x!�񲕾�}	��aX�Qp�<#�v=���=��=�D����V�\��eL�[�ݽ�oX�ء���D���
�=0��=]�=��>�V]?κ�>��>�#8?1S���8�����^p.?��<=Q���|튾�ۢ�Y��p>5�j?J߫?�XZ?��d>��B���A�{�>75�>��&>b�Z>��>bg�o�D�}"�=�>�K>�ڧ=�hW��n��<i
��T��<�g>%?,!
>�<�w<�c���z[��7=�`�����Q���)H4�Y�"�����L�>�Fm?q0?I>,̾���<��`�[�<?I_W?�Q?Ve�?�񐽦�ﾊ�� �a�-��y��>�&�>J�������絿��s�.|�<>��>�@���ܠ�A[b><��i޾��n�[J���羠�L=2}�mTV=����վ�����=�
>޶��n� �8��cժ��.J?%�j=gu��'fU��m��d�>Ø>=�>0�:��v�Ć@����A�=���>�;>�!��3��xG��3�\�>�@D?��]?�q�?�y���0s�;D�/��У�������?�r�>��	?]F>U2�=�ޯ��1�`�d�_�E����>H��>n��}F��Y���6��{ $��9�>��?�7!>�?8�S?�?�_?��(?�W?���>�l��#h��A&?.��?��=5�Խ��T�A9��F�5��><�)?F�B����>��?`�?H�&?�Q?��?��>�� ��C@����>K[�>g�W�Jb��f�_>��J?y��>�=Y?"Ӄ?z�=>u�5��뢾�驽�a�=�!>(�2?�4#?ޱ?	��>{��>��[=�Ѽ>hA]?SԂ?dOj?n�>�	?�\*>ք�>�)=�7�>"��>�"?�T?�>w?�3Q?�_�>�o<�p��\t��~�@��Լǿ�����<&Ĕ=���v�D�P��pO�<|��;��<LJo�i�����s���U����<�o�>�F'>.A����Ƞ�Ԇ�� �>f@�=���0�m�?����ߪ<9U>$��>�;?�gA=^��>_��>hE�$�*?�~?K�?�	��;�o���־}D>��4�>�']?\w�>yh������>p����=�o}?��m?�Ԝ�0��O�b?��]?@h��=��þ|�b����f�O?<�
?4�G���>��~?f�q?V��>�e�+:n�*��Db���j�'Ѷ=\r�>LX�S�d��?�>o�7?�N�>0�b>*%�=iu۾�w��q��h?��?�?���?+*>��n�Z4���(ϛ�cՀ?L5�>�eF��H.?ŕ�ac����-�����%c�K����Г������M���0�������I>��%?��:?��t?�6?L��fL�W!U���S�Z	k��o!��$I��8��<�72N�A˳��Oj��Nk�wH���d�>,R���?��?�h���x�>��ξp �^0�����=�=׾FWW���=:����Cu=�t�=�%'�����%��~�'?h�>_!�=�3?~�W�؃A��-9�zR�_� �qN>���>y�>��?�t1>X�������Ů�c��O��C�q>m�d?�J?��n?&H��v+.�Eā� 1 �B���ѧ��nG>S>>n_�>^��C#��X%�T�>��es�Q���ؐ�(���e�=0?��z>���>V�?��?z��8����b}��0�e,5<�_�>��j?m��>�v�>�������H��>��l?b��>k�>z���Z!���{�K�ʽr&�>�߭>n��>��o>�,��#\��j��@����9�r�=F�h?~����`�s�>:R?P�:��G<�|�>��v�л!�n����'���>1|?K��=>�;>�ž�$�5�{�7���*?��?\���x�(��{>��"?J��>��>���?$�>UG������
?ٓY?l�H?3 D?�K�>bo=��ڽ2�Ƚ5� ��T=�:�>�MQ>�n.=���=_J�ˮX�^��z�Y=�B�=C#μ�t���s<�:�����;N`<��9>9mۿ�BK���پ�
���?
�0舾{����b��Q���a�����Xx�t���'�'V��8c����q�l����?:=�?�~��/��������������s��>O�q�������+��2)��l�ྱ����c!��O�e&i��e�P�'?�����ǿ񰡿�:ܾ2! ?�A ?6�y?��9�"���8�$� >�C�<�,����뾭����ο>�����^?���>��/��k��>ۥ�>�X>�Hq>����螾@1�<��?5�-?��>��r�/�ɿc���f¤<���?0�@jAA?��'�Ô��k��=��>�e�>^,�=r�q��Q$��YѾ�6�>cѥ?L��?�n>XF���q�Z?ū=ԠD�q��<���=��O=�ӿ��S)�Fdc>B3�>eNz���X��eT���;>�օ>�ϧ��޺�܃�'����U>uF��"	��΃?��M�Bg�ŴB��L��k(�;9qd?\�>s�>8?Si@�-�пz�Y��CI?#�?� �?��%?�MѾ��>c@���Q_?��+?�,�>���)�^��u��1���9����þӯ ����<���>R�=uE���龉�ɽ����������.ƿ=�#��0�I=|~�՗g���՗�K-�%ן�
dd��M轢@k=ɖ�=sjG>x�>ZsS>1P[>-X?9gh?L�>�*>��ս���+�̾"���lh�����!���C�C���\�Yr�&2�PS��x��ȾJ =�$�=7R������ �A�b���F���.?t$>��ʾ��M�%�-<.mʾｪ��̄��㥽�-̾W�1��!n�3͟?g�A?����0�V�f���O��}��ٯW?�Q�����鬾\��=?�����=@&�>��=�⾿3�-}S��<?��?�{Ҿ�Ӂ���	>�;���x�=k??��?�ߔ<��>�S�>&���(�{4�>=�>Gk�>�E	?��M�\X����_�"?+�C?;�'��l��H�>%$s�. ��K=�=�BX>1@����'��>���=Kju��	�N�9��=I)W?���>��)�A ��]��6���==��x?>�?��>vvk?��B?�ҥ<W����S���ȴw=�W?�"i?$�>W|��'оǋ����5?�e?��N>2<h�����.��S�N?��n?�`?�ќ��w}���>��r6?4�?���+���rɾ*`3�hU ?�[�>��)?b9��>[sj?k焾9�������B��gw�?v@RT@S�1_���R���g>w��>�¤�~�"�9Q��mD����|>��.>Q�gn�~|⾚�=�y?h�R?�I�>�f���!�]�=����S٫?q�?3���1<]��Zm�2� ��X�<I9�=�����P	�$�6���ž��
�����/M��r:�>�@�}����>�b4�[(�kϿv%���ξ��n��?��>}����j��{t�L�G�?�H�猾�V�>}�>}�������ݓy��p@��v	��a�>�H�R�u>�Y��v��2���=��>#n�>��>�h���Ӽ�6��?�q���|̿�3���'	�2Y?�?�Ά?�?N*�W�m���}�u���1G?R*u?1�P?�2�SJ�X_��%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�3Q?��`��
M�MV���m� Y>�K�����@6����D�R�n�H���n�὿��?��?��?����u�w�,?�:�>�V��1�4��/>פ�>��&>fE=ON���K>Z�þ�@��|~>-c�?���?C3�>�I�i����`�=r�?��>&��?��=��(?{9>z�=�/Խ�(>8!C>��D���*?!�?���>�P�����fE���`�,<s��a�L�N��Ȳ>?<P?gc?v�->}��<������&�r/7�X����n�p���H[�5ï=��)>�=�=� ��˘���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�EC	?����2��V~������6�i,�=g�7?^<��.|>��>�V�=�nv�G۪��]s�^�>�I�?Q��?�t�>pnl?B;o���B�̃2=Z��>O�k??�j����B>Ĳ?�j�7ێ�JG���e?M�
@�m@��^?ﭢ�D�ؿ�U������Z�a�,=�B�<�d=�Ob���?>BA	>֭�<�Ղ=ǐ*>(/�>g�b>��<J=�=XM>f�z>�a���#�Ě��/�����2�ݎ�{!���������IK�I��ڈʾ������;ᄽ�_�)�o�J���+ִ:w��=��X?��P?��o?L�>gA�c}>[����57=����X�=��|>~�.?�E?C�%?��=����d�B���Ʉ��}>����>�VB>B,�>��>�>��/9��?>�zD>��r> ?�=��<�~�;�r{=m�_>ԉ�>��>���>�C<>��>Bϴ��1����h�9w�s̽/�?P���5�J��1���9��ڦ���h�=gb.?W|>���?пX����2H?����l)���+���>b�0?�cW?�>/��3�T��:>����j��_>�+ �1l���)�g%Q>Vl?�xg>1�t>�3�g�8��?Q�3����}>kB6?-���7�L�u��H�9~ݾ��L>�ʿ>��.��'�햿��~���h�G��=W:?�?�W������b�v��q��5(Q>�\>��!=D��=�L>��g�H�ȽG���3=���=�2]>��?��.>#�g=���>�{��
UL��>M`>�+>>�5<?d%?�:z�"5���U��ڂ����>���>��>�b�=JK��d�=�u�>�d>���Aս�{W����2��~E>-^�
�F���f�P�=9�l�;�=�=�o�#�O�p5U=�x?p����ǅ���ľ#Ľ�\'?���>�۪�>?�����-��^%�����?��@���?^"��eS��N?zG�?JB��r >bѣ>L��>���e���e�>;4�o{�6������˽�?��?���\����8^�=��=P�?*��_h�>�x��Z�������u��#=��>�8H?�V����O��>�w
??�^�ʩ����ȿ(|v����>J�?���?T�m��A���@�b��>;��?�gY?�oi>�g۾�`Z����>��@?�R?$�>�9���'�s�?�޶?ᯅ?E�F>!��?�r?��>
�l�h�-������ۋ��È=���:�$�>���=�㿾��F�IQ,���k�����W>��=_��>�ܽǼ�
��=E�Q��Y�h��j�>�Nt>�D> ś>[��>�P�>��>�l3=f����v{����w�K?���?#���2n�O�<���=-�^��&?�I4?�k[�b�Ͼ�ը>ܺ\?`?�[?d�>A��P>��G迿7~�����<��K>4�>�H�>�$���FK>��Ծ�4D�pp�>�ϗ>�����?ھ�,��0K��gB�>�e!?���>qӮ= � ?�#?d�j>�)�>�`E�:����E���>���>�H?��~?.�?�ҹ��Y3�H���塿Q�[��:N>5�x? V?�ȕ>��������E��RI�\�_��?�tg?�I�z?02�?<�??�A?�)f>"���ؾ.�����>$"?x�U�A�$�&�~��?B�?���>������ҽ�k�=i�����C?�\?M�&?��2`��cþ�y�<&���1��J�<��E��>�>>˫���ɲ=$>�=�Ko�ɬ7��i_<Oٺ=��>_��=�i9��U����4?��+=��d�=՝_���L�n��>�ݶ>�?���*N?����1~��`��A����˽(��?4�?j�?�C7��_�A�L?��?�m!?OR�>�ӷ�rPƾ�v �4׋���B��a־��->Jh�>�?������bѤ�kT���\���i��c!�yg?j�>�{?��?�0�>�!�>k|�����"v��ʾ�^\�����=���5�I��)��+���X�$�H]��)���v�>J�ȽjЂ>*<�>�J�>��a><S�>u��=�2>�V'>k5>�%�>m�>���> G>%k�=��=�AV?�۾(�K��m=�5�(�;��>��H?UA�>����[��j�F�UR1?8��?xĳ?�r"?��w���'���?e�$?�.��3�>�M��.���᧾��;:��>�}�>��>��>ҕ��qTy��v��fn��� ?�/?����j�u�=����/�m=IR�?��(?A�)���Q�~�o�.�W��S�f��Hh�3_���$�e�p�1񏿕_���$����(�^�*=��*?Y�?�l�:��^��fk�5?��Zf>���>��>;>%I>k�	�'�1���]��C'����)Q�>�Z{?��>��I?�;?�yP?�mL?_>Tb�>8���V�>���;���>���>՘9?��-?s10?�{?�r+?�c>s��D ��3{ؾj?!�?4J?�?;�?�ㅾM�ýTӘ���f��y������=J��<��׽��t���T=�T>}L?1~�k�8����� 0k>,�7?��>U��>��������<82�>8�
?9M�>"  �{r�%Z��5�>e��?����8=��)>��=�q���/׺Yg�=�Y����=�
���$;���!<�}�=��=�y��ۛ����:_�;��<d 
?jP$?��+>���>�+W����;Ҿ H�=�k�=.^>	G�=��۾����9��l�k���>-~�?���?E�_=p�(>����]��A����4�� ���>��1?^�I?	�u?� �?|&?@t?��$���\ㅿ�#y�}ؽ�	?w!,?���>�����ʾ��։3��?p[?o<a����;)���¾�Խ��>�[/�J/~����?D���������~��)��?翝?A�W�6��x�Կ���[����C?6"�>�X�>U�>b�)�u�g�Y%��1;>ˊ�>KR?���>5?��2?oc?�E>놁�����H��Ι#�b�=���>��?#k�?܉?��>�I>!�Q�2����a���=}����v�����@H0>�|>z�?5?5��=�_��]*��g">.G>�\>ۭ�>?4,=���>fd�>��)�m?T?Si�>)tʾ�����u��z�žg�~>
�{?��l?8mG?e�>EC�3�G���-���>O�?p�?xI@?��8�qc>�=�������U��a�>�W�>\�l>��>�SW��tW>��/?�s�>�|@���1�i���=�;T� ?`�?>�8=U���Ԋ��H�>/�����.>F��=�������\����>�棾��=i~A��S�(���&�������_>$?*�#�3�>Q�>�z5=���=���=v�=qJƽ�u�<�B�O��-�7���/R�r��<S�=���=�Mf=���7W�?dZ?�?�5?�u>��>��j�p>�e�<EM ?�#�>w� �8O;�����t�i���G�2���7�\��t¾S%=��U��>��<w��=�Ҽ��<+��=5�X�{[>�$�=���>R{�=�%�I�>��=��W>��w?Ȗ~�U��+O�e�ݽh�;?b��>ؠ�=@S��\2<?y�?>c���Ji���-��S|?j��?H��?S?c����`�>Ժ��a�{��==Ѫ��l'>�c�=��.�ޱ�>�K>]���ᚿ�;���d�?G�@�->?W튿�xο�;+>�QK>��>ΫS�γ/�-GS��fG��T��1"?��1�˾[��>��|=� �[CξXQD=��N>M�=��ӽKa�j'�=��p���Y=�y=�#�>9�8>W�=�泽�K�=�9]=t�=_J>��5���������DV=]8�=>G>";>վ�>�?
�"?�k?o��>z�_��￾�
ʾ�&R>�\=�ˤ>�yH=�m>7[�>Vl)?'�D?�Q?��>Җ�=@�>��>`d#�Wk��A������ΚJ=J��?7��?���>�G =6zE�$�(h<��6�?�),?\
?�>=��yۿ�W'�!�:����D�*�l(&�����e�1=�{�;%���:����;�=F�>��>��s>��I>3g/>G@k>�>��=v!<V=�<�֧<9����=�t�<JL=̰�;�wK�Er��+��n�E��-j<˂�5܁��&ϻ_�>z��>H��=�p?1L�=K���)>��j��,�R��=�0��i9�q�P��ej��x'�d�4�6��=��=1����g����?�eb>L��>2+�?'|?�<F��~�����3|���K��X�; #>:�=����[�e�qQz��s�ѹ	����>��>��>0�l>�
,�� ?���w=���_5���>�w��.���'�~9q��?�������i�?׺˛D?�F�����=�!~?a�I?7�?Z��>b����ؾ�:0>WH��.�=���(q��n����?-'?��>R�@�D��'˾���B.�>=�G���O�~���/�t���`�����>Db��,�о�$3��_������A�B�o�妺>ufO?���?l�c�� ��]�O��q��m��d�?k�g?��>��?0>?i!����쾘~��%s�=`n?2=�?�\�?˸
>��=N١�%��>�?�X�?�ݐ?�cq?^j>�~h�>�`9<�>_��:J�=�>[p�=y��=?��?i
?5r��?9�����@��,�\�5��<,��=e��> ��>d�u>��=�p�=XO�=mZ>̮�>l-�>ch>���>���>p����9��4?L��=w_�>`�6?<�N>=ހ����p=����έ�1��崽3�`t���j�&�v<GC=���>�����;�?e/7>%龼�?_<߾��U�V5>�2M>������>�M>��a>Ν>iҙ>\�>R>��5>"?Ӿwq>���`!��(C�.�R�s�Ѿ�bz>�����%&����J���I�ZZ���a�j�:,��Q6=�&��<�F�?w���k�k���)������?e�>(6?ތ��O��߮>��>:��>�=�������ʍ�[d���?V��?N�B>.�>9�q?~�?B}[�lp(��^`�Dyf��>M�Bcb�~�l�>Y���qw�s;����R?�'p?��2?����>��?�X8�|��m��=�1�9,C�a�����z>:ɾ�݉�o�ؾ�졾�?�� k�>�ly?���?J?�艾��H�6߈>��!?���>Pov?;<%?:�+?����*@�>o��>��>:�=?�5%?�S,?�g�>��<���=4nO�q9>���U{¾V������㢐<�4�=q]�=\�^=8	����=�do=��>弐=2+=��4s��`k�=͜�<E�= #�>ֶ_?��>72�>�D?����&��Ⱦdv�>6(����y����Sp�����aB�=Կn?�d�?+B?�'I>g�=��J�jg>���>{C>;�)>�U�>ȴ��M5���L=�>Ua>���=Q�r���������b^��z�<h>6�?{�>UU��>ƣ��(�w����>x""���˾!�,�w*���?��r����b>��:?�}D?��C> <ﾾ�'�A1M�ev]?�l?�n�?��?��>`�:b�=Au�+UԾ:��>�1n>6rԾ�)�����&�$��k�<j>EOe��ޠ��Wb>(���t޾Z�n��J�|��IM=���\V=;�	�վ$5�E��=$
>S���%� �'���֪�S1J?y�j=|w��JaU�Yp��,�>还>r߮>�:���v��@�0���.5�=��> ;>�]������~G��8�a>�>SQE?#W_?k�?#"��Zs��B�z���Ac���ȼK�?|x�>7h?B>���='�������d��G�w�>���>M��-�G��;��a0��=�$����>\9?�>c�?g�R?��
?e�`?�*?8E?"'�>���u����A&?;��?��=u�Խ;�T�f 9��F�W��>��)?��B� ��>w�?�?��&?�Q?µ?�>� ��C@�T��>UY�>k�W�]b��J�_>��J?��>e=Y?�ԃ?��=>��5��颾=ة�rT�=_>G�2?�5#?P�?B��>ߘ�>ퟡ��=���>�c?,�?*�o?Ý�=�?6Y2>���>�p�=���>�y�>�?vTO?e�s?��J?P��>*b�<%3��/V��9os��P�Y΄;ԓH<w�y=�~��t�}3��)�<�c�;���bO�����#�D�%���[g�;bv�>s�s>�����0>��ľ4)��n�@>P��Yg��������:�"0�=*~�>?U�>��"��=o��>vJ�>g���'(?m�?��?%|
;��b�:�ھ�=K���>)�A?�z�=��l������u���g=x�m?�^?σW�x)��_sa?%�f?S8�lF�Si�J�>�������z?���>���?��h?-�f?���>����ft�\���m�P<V�'�*�J�?v���@�_F3>��2?�õ>0a=�n/>�[��sL�" �Y� ?��?mU�?�x?��d>���|���>�����f?I��>�Q��t ?�a��XϾ�+��^3�������7Z���皾����Gi���+��$퉽+>� ?�wM?BD�?՜c?�Ͼ�SO���p��,s�2,L�u�뾄�
� I?���F���>��aY������kǾL��􅾮�V��:�?�o.?y�x� r?�ҡ�Ю�A�xzk>� ��tO�(�}�5�!���*<M�<�n�}|н>D����4?���>\�}>U;0?J]P��FP���5���;�s�n��=���>�R>b��>�Z=?��#݊=N�h���F������(v>�{c?Z�K?�n?�{�)*1�C���Ǖ!��2/��[��\�B>�>�ˉ>k�W����7&��W>���r�?���|��*�	�#�~=��2?�8�>���>�N�?j?jm	�ca����x�Ԃ1�#��<�$�>� i?�4�>-�>�Ͻ�� ���>j�l?ߕ�>Q�>ϟ��IY!��{��Qʽs�>y�>P��>p�o>�,�& \�ek��񄎿 #9�k�=.�h?����k�`�{ԅ>WR?���:�I<_m�>�v�U�!�(���'���>=}?���=��;>�~žL)�c�{�%B���)?��?y���H-*� �>Q"?��>'�>�	�?�m�>�þU��9�?�_?޶J?MA?ة�>7�=Y謽��ǽ��&�;Y+=Cц>?Y>U�p=�h�=�P��T[����N�E=,��=��Ҽ�����%<9_����U<L��<�3>mۿbCK�s�پ�����<
��刾᯲��d��ٲ��c������Vx����'�(V��7c�����-�l�͆�?�:�?Lu���)������	��������>��q�Z�����l���,��I��y����f!���O�(i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�|A?(�(�!�쾯6V=2��>O�	?�?>�W1��I�����Q�>6;�?���?�oM=c�W�D�	�ـe?��<��F��3޻J!�=n<�=c=y��F�J>�V�>X���UA��Bܽ��4>@م>�"�����^��E�<�]>P�ս�7��_҅?'�P��^I���7���W�b�=S�2?��>����^?��E���ǿ�}P��j?�n�?A5�?R-?�¾O��>Yξ��3?��?i�y>F�7�;���Y%>�==�)=�9��Z����=�pv>�����Y��J�Ծ����>���j�=�� �ʿ����m6���=�ԃ=��;��\ܽ7�Z��߫�vm*��ɽi=l�>=?��=���>l��>���>i�Z?%pO?(�?��:>��&�VU}������<�垘��O���(���#���F�I�%��,��s���Ⱦ!=�1�=7R�n���J� �d�b�V�F���.?�v$>R�ʾ��M�Y�-<vpʾY���H܄�'᥽�-̾�1�#"n�f͟?��A?������V�T���W�����J�W?!P�޻��ꬾ���=ެ���=%�>���=���� 3��~S��t0?3]?�����_���*>�� �+�=�+?��?�@Z<�(�>M%?��*�f+��a[>��3> ԣ>]��>1	>����]۽*�?��T?	�������ڐ>�d���z��a=->�.5����j�[>e=�<"���U��>���|�<��^?`��>67�11�eѾ{jL��+=���?�,�>��>?��@?Yz<=f��g�e�	N�xX�V�V?=�j?��="׻�u���׹�"�,?�o?X|<o������$�Zk��!?�Ȃ?��!?6Ѡ�􈁿������0�M5(?��v?�r^�bs��>���V��=�>�[�>d��>��9��j�>ϑ>?b#��G������~Y4� Þ?��@z��??�;<�!�e��=�;?�\�>:�O��>ƾ�y������a�q=r"�>����jev����LR,��8?���?C��>m���������=0╾#[�?`�?(x��F�g<a���l��p�����<�=oS�zr"�����7���ƾD�
�ᣜ�ѿ����>�Y@4���!�>MP8�5�CTϿ=���^о�aq��?xs�>�Ƚ{���V�j��Du��G���H�ǡ��N�> �>ۯ������,�{�*q;�Z8����>��n	�>�S��'������5<��>Ư�>���>�*��H罾ř?�a���?οD������d�X?�g�?Tn�?.p?�s9<��v��{�m��D.G?։s?�Z?�l%��>]�h�7�%�j?�_��yU`���4�uHE��U>�"3?�B�>T�-�}�|=�>���>g>�#/�y�Ŀ�ٶ�D���Y��?��?�o���>p��?ss+?�i�8���[����*�`�+��<A?�2>���G�!�A0=�RҒ���
?S~0?&{�g.�1^?�Q�?�N� ����=�n�>v��g�辶�H�U>q�;Y�`͜��b\�'|�?��?m��?���&'��"?��>��7�1�ܾ�Q(;p��>��>��=9��9M>+���W!>t��?FK�?�� ?��p�O�Y9g=��w?]!�>ˈ?�[<���>�ܤ�������=�	>={,>������*?O?7�?��K>L�g��`��pC��]�Z;��"Q��D>��i?�Q?ʰ�>��]����;r%�cV=j�_��+ݽ�&�=�=7�$��}%>`�> B/>�A3������?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ua~����7�b��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=7M�>͜k?�s?�Qo���h�B>��?"������L��f?�
@u@a�^?*�Sҿ+��;w��t���5�>u��={�S>�m��Y��=g��=x��<���>r��>>�`> S>M�m>>~7>��,>Dk����&�D��!ݖ�@>K���_���Z�]��$�T�8��T��}q��1���J���P�Ľ��<�6���J^��!4<��m?	�'?Hh?�>`�S��>������>;��>97�>��T?~�0?��?-��<�料�2O��K���B���Ҥ�z��>	!g>�-&?J��>/Ͽ>I��=��>A�d>�ѽ}>�M��8����;>��= �>���>��?�C<><�>Hϴ��1��|�h��
w�N̽1�?Z���I�J��1���9������di�=7b.?�{>���?пl����2H?����U)�Ϲ+���>]�0?�cW?��>�����T�c:>�����j�p`>�+ �l�}�)�x%Q>;l?��f>ֺv>�3�_8�%Q�K���3}>Y6?{l��mO:���t��aH��cܾi�N>�4�>��A�x�5�����^j���v= �:?d�?�����D��� u�]���ͭQ>\>u=�=ׂN>��c��PȽ.�F���/=�o�=i�^>iB?�%,>h��=��>�V���FP����>�B>��,>:@?�%?O��D$��l����-�"�v>�4�>6��>44>�NJ��Ǯ=nY�>2�a>C�`˃�����?��sW>ˆ}���_���t��Fx=i���+�=~8�=�m ���<�((=�~?�~���∿.��M���lD?F%?��=UF<˂"�:����K����?��@�m�? 	���V���?�@�?���̲�=�|�>%֫>�ξ1�L�#�?��ŽjĢ���	�M$#�R�?�
�?^�/��ȋ��l�/9>�]%?�ӾQh�>xx��Z�������u�n�#=P��>�8H?�V����O�`>��v
?�?�^�੤���ȿ6|v����>X�?���?f�m��A���@����>;��?�gY?poi>�g۾?`Z����>ѻ@?�R?�>�9���'���?�޶?կ�?aI>���?�s?�k�>�0x��Z/��6������$p=�[;�d�>�W>f���xgF��ד��h��u�j������a>��$=+�>QE�[4���9�=��I���f�<��>�,q>"�I>W�>v� ?�a�>}��>�x=�n��Jှ�����K@?���?��0�GSl��q�6H��u�����?|-+?Ը��/��39y>H�Y?�B�?2�1?�PC>�
�� ��Ͽth̾����>���>Υ�>,]�G{�>��
���0��	>�4�>^|<(瞾ZO������>��!?���>We��� ?�#?��i>��>��E�:I��'�E��.�>*��><�?(�~?X�?�۹�b3����_ӡ��J[�+&O>�x?�I?X��>R���!���h�K���H��+����?�9g?$��I2?�G�?$�??ɚA?�e>�O���ؾ������>�#?E��\>���#�����	?؉�>0*�>�	��,�ѽ˓���z�����?;`?�"(?rI���_�=V��-��<�LB�c�e:�.�;ߏ��HU>�H.>��>�-��=��">fz�=��i�ǹ9�ϳc<�F�=8Д>���=r�2�	����<,?�!G�`Ѓ��Û=0�r�4D���>�qK>j%��-^?�>���{�)���r���hU�| �?ޤ�?Wl�?%s���h�.=?��?d6?���>@��,޾Y�ྷ�w��x�tH���>�C�>�`s��K�S������.	���rŽ(K���>��>~$?� ?j+P>3�>�C���&'�q�?���^��y��u8���.�|���Ġ�-�"���'#¾R�{�H�>������>+�
?�h>G�{>���>�xȻ{I�>S�Q>�4>�V�>5�W>��4>��>k�!<�нLR?����־'���ű��w3B?�pd?10�>�i���������?y��?�s�?�?v>7~h�k,+�n?�>�>���q
?�V:=@�1�<�U����U.��<�p��>RD׽� :��M�9nf�aj
?�/?���M�̾�=׽����i�n=5N�?�(?��)�j�Q�.�o���W��S����/8h�yi��2�$���p��쏿�^��%��A�(��u*=�*?��?h���� ���%k�I?�/cf>�>[$�>�߾>�rI>��	�B�1��^��L'�����P�>Z{?G��>�~J?��:?)�P?3oJ?�m�>���>������>B� <|q�>&}�>Ҍ:?��,?'�/?��?"�)?�_>��i\��\vھ�`?r�?<1?b?I|?����^尽�ǌ��6Ѽ�x��p��Zj=�[�<��ٽ�}k��_=�R^>|U?���k�8������k>�~7?��>���>���$�����<3�>n�
?�A�>����zr�rb��S�>2��?��P=#�)>m��=#���5xϺUX�=�����=Y#���o;�!<�~�=j��=Nt�ͯ^���:���;��<�"?ک?��>�?�uľ���	����WC�;o�=�+	�I��=�������=Y��VAm�2�8>�[�?{a�?�tb>��#>��>D���S���G��	��H�=��P?:�<?į�?�Q�?�P?��/?ʎ>@�	�8i����m�xr�	�>>P+?.�>;��i�ʾ-;��2M5��?hZ?ݪ^�����#�m!������i>)/��~{��X��w}E�p�����������?A��?|�(��s6��&��0����B?cG�>��>���>�#)���f�|���c;>��>HQ?]�>�IF?�t?�:V?8�r>Զ,��(�����{���>f�7?��s?؈�?,�?���>�x5>7��4ྉ�⾽Y�hv���ps�_Z=��K>���>�A�>*5�>�o�=������p5����=wXs>|��>Y�>>��>�s>?�<3H?��>:�����uڣ�腾BE�ǳt?Wŏ?73*?���<X��*�E�����;>�>ܨ?ի?�)?Q����=W�м����Z}k�4+�>k,�>2�>�+�={L=��>\��>3��>�@��|��+:���Q�S?EF?�s�=zǵ�'���R>:�N�eK�>�97>�<��0���O����;>�pپ����d�聹�t�ξ�m�f)޾�ϥ���Z��
?�[Ľd�]>�Gz>� >���=6�ȼ�N=�����=p(�bl�#��׋��"���>W�=:��=!|Խ��;��y?ϣ9?(m,?Y:?��Q>�1�>�'� �>�9μ� ?�>�8�<��Ⱦ����I��������оҁľ(�P�n�վe�=j:ӽ��n>��>��=���<��=2��=	.s<�K==��%=�sI=���=yu�=p��=b�>`=�>�6w?@�������b4Q��V�F�:?�6�>_t�=P�ƾ�@?��>>�2������b�.?V��?�T�?��?�si�~e�>����ꎽ�m�=\���q=2>h��=m�2�2��>�J>D���J���|���4�?��@��??�ዿ��ϿEb/>��7>�5>��R�}�1�=�\���b��lZ��!?E;��M̾B�>d	�=)!߾v�ƾ�s.=o�6>^5b=J}�g[\��Ǚ=�{��<=�9l=ى>��C>�y�=�S����=��I=���=��O>�5���7�bP,���3=A��=��b>�&>ª?E��>��%?2�J?�(�>�罞����ܾ�d>� >2w�>�|X��;>��?M5[?��T?d!I?S@�>3�=���>ԣ�>����2g�$v��Ϻ��d>9�?��p?5^�>[��;�^�*��jD���B?�2?��>�[>�����ҿ����@��҉���~=��=�3k�� ��M�:8۽O#�r��=�9�>0�>�mc>�H�>�
�>Ni�>�u�>���=�>����n=� �=�e=U�=��,�-��	E.�T=�������|Xɽ�h9<��HF�=�`�=��=���>/.>���>�=�峾�5/>�Ζ���L�AȾ=�\���0B�`9d�^H~��/�6��
C>�oX>�N���1����?��Y>�?>Hx�?�<u?� >3>���վsM��e��cS�+�=C�>6=��;�@U`���M�iҾ���>0�>w�>��l>7,��#?�U�w=_��`5���>Fy��c���!�Z8q��?��e���ai�+�Ӻ��D?�F�����=1"~?հI?��?X��>+��Ņؾ$A0>�F����=��w(q��k����?�'?o��>���D�KH̾0)��-�>L8I�P�O�������0�����η���>����оx$3��g��-���3�B��Lr���>��O?��?�3b��W���SO�����<��$o?�yg?E�>�H?�@?�7���w�Qp��܇�=��n?���?N<�?�>a˳=C��� �>͆	?��?+��?}�t?!�8���>A
<t�>�t��o�=�>�̩=��=��
?״?�	?� �����w
�����N�G��<'˚=ŋ�>���>Y�t>j��=�=&��=O�T>*O�>ʕ�>7;d>~(�>-��>�Ы�N�
���(?��=k�>$�1?x��>�qW=���G@=����*��S'�F�ҽ�.޽��a;����^Y+=�"ڼs!�>��ƿm�?MS>u���xx?Ϩ��%�%�F>[/W>rI�ad�>W5>�'j>5խ>L��>�>�Շ>Δ1>�FӾl�>���ed!��,C�)�R�X�Ѿ�}z>;���	&���.t��"AI��n��g�_j�4.��4<=�ɽ<H�?������k��)�v����?`[�>�6?jڌ��
����>���>~Ǎ>K��)���(ȍ��gᾇ�?I��?a�s>ޤ$>C?Z?1s?J I��6 ��b��}�#�E�+UV�i�Y�␿��}�nv�m:���]?Uv?�$7?�<�ַ>�͌?ڌO�j��1�%>�r,�~}V�ψ�#"$>Xݾ��/�b���}���g=Uư>elv?Ow?�,�>��F��Tj_>{9?��?��\?}�?�X?��D;_?��>�ʯ>�:A?K?ֽ�>7?�%4>�$=^Ȼ�8�>>ν^ʑ���%�D .��_�Y��=��=��-�a�C<���=�;�<�m��\>��=x�,��	>߉a<궩=�>>���>z�U?+��>\�>#y2?�X�<]2������ ?b�)��ʒ��	��G���6���C�=UBl?��?�:^?��j>��U��B�8Q>��>�>�hf>��>�
��FZ��Q:=�# >�>��<{����꒾����p����=vC&>��?�>" ���[<>�w�O����:�=;z��7̾(�Ҿ�`\��:��;��]�>��<?;�Q?���>�`Ǿ,�h�Ά]�rV)?�?�z�?��J?Lt>Ŏ���OG���2������k>�Z ��) �T���􁻿ŁK��@�=�a�>�����򥾔�R>)����ݾ#i��%E��u�==����=���~SϾo��K�=~��=dʾ:�%�%��]̪��J?��J=�����CJ�%���B9
>�ē>���>�CI���L��`B��������=�,�>�a<>Nм�n~E����g>�>SQE?3W_?k�?"��Qs�2�B�s���_c��BȼE�?kx�>*h?�B>���=C�������d��G���>���>a��N�G��;���0��C�$���>N9?�>��?_�R?~�
?u�`?�*?EE?4'�>+������EB&?���?o�=��Խ��T�� 9�nF����>p�)?S�B�d��>J�?۽?��&?)�Q?��?��>(� �BB@�Z��>�Y�>�W��a����_>�J?)��>�=Y?pԃ?�=>�5�}颾ީ��P�=�>��2?7#?Я?֬�>y��>���{�i=Z'�> _f?��?Y�f?3��=�� ?&>��>+�>�и>� �>�_?>�H?��q?�}D?}<�>��=p�ս�ڙ��ʏ��JǼ9�=��y=ktw=��g�J�м��A��b=��<�N�Ct�����V`z��"M�0�Z?<2f>l��Q�>�Ⱦ�c���r=���� ξB���rv���0��+�>6,?ʐ�>3��<g;�=�֥>Z��>�s�/� ?5X�>	� ?c3�l�W���P��b-� �>[�=?v=�n��o���	���y=0�{?l�c?L]�����+g?��q?n!1�J+����`ھ^��#�A?Ec?V¾\�(?,W?B�R?�a�>�Ů��w�ȩ� �y�:�7�V<+t�>:� ��~4�F{
?\4?N?y�X>D'=���E<a��/�Д?D��?Y\�?ֆ�?���>�vs�mտ#���ɔ���p?��>�C��b3?p��=�B���M���9	�J׾$h����[ئ�5w���}����+�V��d;;�)?��l?��e?�j?1�پ0�Y�H�T�|�J>X�X2����ԟR�@j?�̩'��dB������q��H�b���_<+�y�4H��|�?�~$?���Y�>v���s-��߾"�P>�#���g�K\ӻ����K�<4�;�m�k�O������D(?�R�>%K�>�a=?�LT��4@�	u6��?����A�>N��>�0[>�]�>��=bA׽qꍽA���L�c��D���6v>yc?�K?`�n?�n��*1�څ��Ҙ!��/��d����B>�k>z��> �W�?���9&��X>�q�r�\��Cw����	���~=��2?*�>���>bO�??,|	�l���mx�M�1�
��<{1�>� i?[A�>��>н� �(��>:�l?�&�>/:�>����"�){��nƽ��>7�>,� ?�bn>$-�bg\�H��������:����=�h?1����^���>y�Q?�;4L<��>��|�;�!����t�$�v�	>��?+��=qy=>+HžcM�|�|�g�����?�>?	����.;�5S�>w�*?�k�>@�>�_�?��>�̮��#�=@p?5�K?3??"65?���>�$�=� ;�9��7�����	=�g�>B]>��<�j�=��1��BI����;Ƀ�=s��������~:�#��:	��;�Jr=x�P>�Tۿ)GK���ؾ<I�I��	�Uu��$��������������Ǚ�zgy�{x�8�,�^�V���d�lV���l��W�?a�?:������b���s��������>xat�#y���Z���"�����z��F֬��!�RP�Oi�D�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�rA?O�(�,��(mU=T��>ӕ	?�@>�-1��9�p氾EH�>$<�?m��?�-M==�W�þ	��we?(k <��F���ۻp��=�v�= �=�����J>-k�>�Q�GPA��۽�4>^Ѕ>߆"�����_^�b�<8�]>��ս�S���t�?�.?���X�l--��΂�SM#=�66? Έ>���?�W���ӿ�jZ�4�g?�g�?��?1�0?v�ӾuG�>� ˾��5?��-?px�>�2�f c�Xc!>�6�<*�<�E���D���׼���=L�����T'׾�ƿ�1L�m%�3����¿����Y2�2�c=m�=�^�-�j�$�f�C�w=�'���A�Qt�d�<:�A=�b%>`�D>�>�^>q�V?��n?e@�>>83>]ƈ�J6C�q���D����۾��.�������^��<ƾ]��*I�|r�eM#�T���Ѿ!=���=7R�v���'� �F�b�?�F���.?$w$>X�ʾ��M�:�-<XpʾU����ۄ�*᥽�-̾�1�"n�b͟?��A?������V�J��eW�����S�W?�O����wꬾ���=j�����=�$�>w��=q��� 3�m~S��e%?|?S!���Ę�&X>|���.�;�g&?�d?;�<��>,9&?����xܽ{�X>Md@>�[�>�~�>¢K>�{���ϭ�2?!�f?�½�ܯ�a��>�Ͼ{č����<��=�K$�s�5��W>wp ;8�r�_pn�2�)�U��<�{X?T@�>9�.��9�v�������k=u�w?��?=�>�-t?7�;?�`<�e ���Y�?U���<{S?1�c?��>u-C�H�۾�����<?�`?��V>o�s�����7�����?A�p?γ ?��Թ�y�R����
�/?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?n�;<��U��=�;?l\�> �O��>ƾ�z������3�q=�"�>���ev����R,�f�8?ݠ�?���>���������=.$���a�?��?.���-n<	��9l�����*^�<\]�=�L���%�g��I�7�x�ƾ�U
��|�������>r[@�-����>�8�n$�MiϿg?����о��q���?Ǳ�>J.Ž����Aj��t�Y�G��H��鋾V�>��>����.���b�{�p;��⟼!�>Tk���>v�S�x.�������8<���>T��>ɷ�>^+��yս��?r\��{<ο[������&�X?�i�?�o�?n?J.:<��v��{�ɳ�v$G?�s?Z?�"%��G]��@8�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�GFj?�rD�lN�J���A���>�8�U��Z'���vp�x^��&��x_��P��?���?��? �꽡K���I?�N�>}"����vL���) >a�>��Z��~��tj>C2��� ���F=���?���?w1?��X����">lX�?sA�>5g�?/���?t5<=j���P>��>�NJ>��8(?��9?fq�>Zr>�C'���&�W~�#LO��+�%�K�Ĭm>ۅu?�;;?��>��:���1 �?����^����T��$����8>��2>��g>��`<�u����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?rQo���i�B>��?"������L��f?�
@u@a�^?*�,Կ*��l̾DQ־�=e=i�=5�>���<��=t`>�:�<#v=z4F=C+>>�V>'�I>��E>�3>_5>È��$��^������z�6����l�7�?�F�ھ���m@����M}ƾMz �AJƽֶ`�s޽#�-�N 1��-�=��U?sQ?Kp?�V ?��~�7">%V��t�=�$�#$�=4�>>2?{L?�B*?\D�=�̜�ced��h���ڧ������V�>.�H>h��>��>��>��r��I>,�>>��}>o>^�*=����=�0N>4��>���>��>�C<>��>Fϴ��1��k�h��
w�l̽1�?���S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?%���y)��+���>|�0?�cW? �>!��r�T�3:>8����j�6`>�+ �|l���)��%Q>vl?��f>�Eu>3�3��X8���P�/�����|>66?׶�l9���u��H�\ݾMSM>|��>�D�c������=�i���{=q}:?E�?�Ĳ��㰾��u�a5���OR>*\\>��=wX�=�OM>Kc�`�ƽ��G��U/=��=�^>"�?�K>>@C{=*3�>b��b��9�>S�M>U�4>^?>?��'?n���Ջ���}�[�,���m>N��>��>y��=��U��f�=�-�>�c>��������H F���R>��f�|�n�au}�i��=�������=S�=�x�.�(��Q=�X�?�Ӟ�>ӄ�qw��o����2?=�>�d����/H'�K.���Ͼy�?$�@ES�?�����Q��k?>��?�l���=|6�>��>7��GB]�"�?^��苾����Զ,�卤?�p�?��t�7r���N���&>��?p�ҾPh�>zx��Z�������u�s�#=R��>�8H?�V����O�c>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?roi>�g۾>`Z����>һ@?�R?�>�9��'���?�޶?֯�?]I>���?�s?�k�>�0x��Z/��6������Wp=%�[;�d�>�W>`���wgF��ד��h��s�j������a>��$=)�>PE�Y4���9�=��	I����f�6��>�,q>�I>W�>t� ?�a�>~��>�x=�n��Kှ������K?P��?�����^�s�rcA;G���R	?5?al��D��l�>�U?��}?U R?���>h��P����ʿ��9�����<�Fq>Z��>^0�>�ݸ�3�f>O^��]6��Ǜ>]˅>����Ӿ�#o��!�<�R�>�y/?EI�>��R=K�,?D�/?S�=L~�>�!v��l��rt;�/�>��?��)?�č?�.�>��ԾA�O��۝�_N��h�m���>? \?��?}��>v �������=cp׽��Gg?NU?b1O�Y??�H�?h"I?.�:?Ȓ_>\�Pb�=���.N>��!?����A��T&��?�IW?T
?�]�>�ߔ���ս�uۼ����+���5?q]\?>w&?/c�Pa�U¾���<�����O��)�;�U��h>wV>�Ά��Ҵ=i>�&�=ϼm�[�7�}R<���=�ǒ>���=jZ7�疐��6-?�{+��2��8�=�4s��D��^|>l_@>�þ�Z?��A�L�}�����cW��p�S�-m�?���?L1�?�½��g�b=?�p�?�?�!�>U���*پ�߾��j��v�	M��Q>�_�>�t���8����Oϩ������@����>��>�?:s ?�O>�[�>�혾��&��)񾐖��l^��?��38�Я.����*����^#�]
�&¾�p|����>Fq���T�>��
?Bhg>-{>*��>,��ӯ�>4SR>ߞ>[�>X>P 5>;">��"<B�νdnR?����Y�'�a��܏��>�A?6sc?��>��n�{������T�?���?1��?u�x>��g��+��c?Lz�>���c
?+9=r��ۼu<�c����[C��aI��ʎ>��׽�:��'M���f�+D
?�c?�
��ψ̾M�ؽL{��ea=�|�?��'?�Q(�hP�q@o���W��HS�?��dj��ߟ�oq%�g_p�$���V���q�����)���=y�*?b�?����$6뾓e���k��?�oe>D��>�d�>���>T3L>�	���0���\��'���Yh�>�'x?�\~>�X?��"?iUV?�=?�c>T`�>S�p��?�ܼ��>�
�>K\0?�&?�&?x"�>9Z?��y>
�K����_�<#?7 ?)�/?rG?�s�>�j��
5�p��~R�z<$��æ�ۼ�=y9�<s���EF��|�=3V�>b,?�=�^�3������|>e <?���>c��>�z��s�&�-=�G�>��?2�>8����m�R���=�>��?d��PI=�i#>ʮ�=98c�M'9�{��=�ʼ���=�4;�e�dM:���=c{w=>��<g�ڻ�1�<�=E=R�?�� ?�\>��?!e�4���J������>�h�=�� >^'��������E:u�8�E>��w?��?��r�*y&=��>������X���B�=��r<�5?btl?B�q?`�?��N?�&#?�و<2�H�/#���t���~�x�?\!,?�>����ʾ-�ʋ3���?A\?:a���8)�H�¾b�Խ�>�Z/�j.~�6��HD��+��g���}����?#��?c�@�l�6��v�ݾ���Z���C?/�>UW�>_�>0�)���g�O$��6;>��>�
R?@Z�>��O?,{?��[?�JT>Ɣ8�VG��s♿� =�ei!>G�??q��?���?+Vy?u��>{P>�)���߾�����?�!��₾)~V=�DY>�c�>:i�>t8�>A-�=�ǽ������>���=�Eb>�z�>�ҥ>��>�Hw>'��<,^H?�+�>������T��o����F���s?�q�?�)?���<��A	G������>�ި?]��?�{)?��V���=�qż�紾>j�Jw�>���>�u�>ǯ�=�V=y>W��>F��>	�����:���n��|?��G?�=����B�q��~;>뜤�>_�=���*[���ƽ�������>�龄�Y��XϾn���+��-���40#����u����?��ؽN��>d>n}�<S�=<�=�N>"�d�=cEý\�A=����;=&XS���4=7;��q=Ƨ���ƾ�]|?�kA?��,?n�C?g�>�	>{��@��>�!�us	?�,c>�	]������4��訾MR�����U";��f� ����>�ӈ�)Z'>ԀL>�6�=��Ʂ=¶�<\�=ꕼ�9=�{�=���=�h�=j��=��>-Q>�6w?X�������4Q��Z罥�:?�8�>Z{�=��ƾp@?|�>>�2������xb��-?���?�T�?>�?@ti��d�>I���㎽�q�=N����=2>d��=}�2�R��>��J>���K��6����4�?��@��??�ዿϢϿ:a/>��5>��>h�Q��4�ۍV��:[���X�h"?U9��f˾5��>>n�=`p۾A�žy4=,�4>��{=6��Z��x�=]�z��8=��S=�f�>ssE>R0�=����լ�=��[=f��=IOR>���ME���/� �,=T�=}Za>³*>=C�>�~?��*?�&_??��>p�q��tܾۆ̾,�z>���=σ�>y*=�N>35�>��>?[�H?�<H?ԯ>�[�=�h�>�a�>v�)�5�j�m�9��)�l=4�?���?�e�>�s�;֍J�
H$�m�@�\�Ž_�?�2?��?X4�>w	��jֿg+��cV���4�0q-�ï�ЁL�~>��=�0�;�t�=��=(�K>��>��u>�t>�>I:>�̯>y��=pn�=��Q=�0�<��Y>&�c�){�<Qq��!5>����֝����@��Zi9�eRc�^p��������F��=� �>x>���>6��=����/>����L����=|���B�Dd�8~���.�؊6���B>NX>nu���1��W�?�lZ>�i?>2��?�u?�R>�{��վ=K����e��S��=S�>��<�hp;��\`���M�Ҿx��>��>+��>��l>�,�'?��x=u�HZ5���>Zd��Q���"��5q�?��b���Hi���ںe�D?+E�����=2~?t�I?5�?���>[�����ؾ�00> S����=+��q��5��� ?]'?��>쾾�D��G̾�"����>~?I�r�O�!�����0����η�|��>�����о�$3�4g��u����B�Qr���>ԳO?��?9<b�%W���RO�����%���q?�{g?[�>�H?�@?�2��0{�q���y�=��n?��?%=�?�>|�d=�m��r��>��z><�?��?za?EAν�<�>��<�y�= �)>^�>m�=�U�=u�=OX?�-�>�A?�|</H��ݻ���4��#���yV>
�!>y��>X�>Z>�>�76>��D>��c=���=mHy>[H >�M>q^7>�>&��h��̎G?�n�=Vݚ>w"=?�*�>v8�=�&+�L�>=,ν���.�^�� �՞	���N���7k�+���w�>�`����?���>R�޾�)?|���~�����c>��=���[�>�H�=��r>��>�W�>%d�>n�>%�f>�FӾ�}>%���d!�s,C��R�I�Ѿ�}z>2����&����u���BI��n��ug��j�j.���<=�X��<)H�?������k���)�?���q�?\�>�6?Rڌ����Ȱ>V��>lǍ>wJ��3���ȍ�ggᾔ�?��?7X�>x;>X�k?M'?�:���ٽ�K���{�L�O��2Z���]�����3ă�����ELC���T?~b�?�;3?�-����>>ԏ?��I�쩅��;>��9�du^�|Q�\�A>�*¾ixT�����F�b�=��>���?��w?=n?����	��H�>�-�>�n?��o?�#?-R�>�&<"7?���lH>��?��S?Q"�>�c�>В�=�dM>��V>m��=?���<M���;�D�p=[�Q���D=�"�<�AN��=]��=�=8x$�c��<�b�=��=�L�:�Q�=G��>TZ?ޭ�>Y�~>�:?*���!7�����F�.?�9=Y}��v�w��3��PD��R>%h?�_�?��[?Dl�>�=�~�;��6>!@�>=+,>��:>C��>�=�0�Z�^�M=��=��&>n��=�_I�����M��kp�����<Q�>�?ϒi>G���Y�>�,˾j[����>��� ��1C����S��U��̾"W�>��O?%�L?�/O>2޾��"�;�X��"?��:?��a?��\?��}=�鵾�k6����%Td����>,�=~G�����2����X��j�<�R�>����J���'a>;�A޾�#n���I���羖�L=����T=�(��վ������=��	>n��C� ��"��Ī�5J?�g=>줾0U�|���>���>w�>��:�Fmx�F�@�?���/�=O��>��:>i�����cG��.�h�>sE?'I_?tc�?D�����r��QC����������Ѽ�u?�Ǫ>�;?۬B>YZ�=��������d���F���>��>��=�G�x,�������$�,�>�?�>��?rR?��
?$&a?��*?��?�D�>.���r����P&?�v�?<��=ͳֽ��T���8�m F����>qM)?�VB�Un�>�M?.�?('?e�Q?��?��>�� ��&@����>�q�>��W�!b��.�^>��J?'�>�TY?��?>>bs5��:���F��'"�=rb>U�2?JI#?<�? ��>�}�>����`ڀ=�j�>Kc?r6�?\�o?�N�=�?*?2>���>�=e˟>_b�>@�?�3O?��s?��J?�y�>���<և������s�t��HN���;�*G<�vy=+�*s�[��R�<���;��������f���E�=��#<�;{��>��s>�ϖ��>��ž>.����>>/�������Z��q?�A��={o|>A?ʸ�>d^�e�=���>)��>O
�7�'?A� ?[?��"�Mna���оsA�J��>N"@?���=�rn�<��zw�m�c=ːn?��^?�EV�7����h?��[?�������������-�����?���>sb=k�?D�c?%g�?�t?�����|�|���`N�D�徖JH=��>VN�3�F�u��>ީ]?�>
�>�2�=);�I�a��鍾�Y ?&ו?�?�?ޅ?�Y>T���^���<�f���uxa?�o�>� �U�"?W�;v�ܾ�9���Q���׾� '��ͼ��Ͼ�������Bت�J�a�W�|=�&%??�K?6]�?q�D?��۾��H��M�Da�x�_���Ͼp�!���P�\�C��#�0�T�;o(�9�徑o��|�;AaZ���W�G!�?�0?&�=+�/?�j��+!�Q��x�Q>�{پP�@�?�a�m���8��?�۽C�����aD���>!?��>�}�>ҥ2?��S�f�'��=Z���Z�r��p{9>�>�F�=���> +�=Cuѽ��<�6�Vc><�#�:85v>�yc?��K?'�n?�n��)1���8�!�ت/��d���B>+k>���>:�W�ҝ�:&� Y>���r�}���x��Y�	��~=�2?�)�>��>~O�?�?o{	��j��nvx�Y�1�ܡ�<�0�>i i?g@�>/�>�
н�� ����>-�l?���>��>o����Z!���{��ʽ�&�>�߭>0��>��o>��,��"\��j��0����9�y�=�h?�����`��>�R?͊:VH<�|�>�v�ϻ!�?����'���>�|? ��=0�;>�žN%�^�{��8���/)?�I?�ؒ��*�ә~>V@"?XZ�>��>Q2�?�-�>Yþ}z��4�?$�^?"J?v*A?�>�>�(=Ơ��e�ǽf�&�[Z-=`D�>��Z>Cm=���=���i�\��+��D=$��=�tμH���>�<rg���J<��<�4>�gۿ�GK���پ\�����)
�5Έ�c���`W��4���H��ƽ��*cx�G�FB'��V��ic�����o�l���? �?��k$�����ń�������>5�q��~������oM����n����}!�h�O�0%i�1�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@~A?��(����aV=���>�	?�?>�S1��F����:P�>J9�?K��?�GM=a�W��q	�y�e?4�<��F��޻(�=�l�=��=����J>5T�>&��XFA��?ܽ�4>}�>>"�����^��̽<�t]>Z�սH(��`�?�<���u��bq�b����f�=�gW?]�>Z,j>�?�H`�E�ܿ,�z��]f?݅�?�!�?t�E?{$;���>=i���=&?���>��>�?@���g��~�>��=��m>R`ݾ��(�<�x =hy��P�]�S����xe��=���-� ���ÿ�� �A<�XQ�=�;�e�,%�bN��� ��΄��V�/����e��;C��=�G>1*o>�8>/�O>�.[?�]?���>c�>=ͽ��%���s��������ߖ��ϊ��)��F��n%۾�A�A������v���!=��	�=�6R������ �a�b�>�F�u�.?Lv$>i�ʾ[�M���-<�oʾ����M܄�Pॽ	.̾�1��!n�͟?��A?������V�4���P�����Q�W?nM�ڼ�I鬾���=-����=�$�>ʊ�=x��� 3��}S���0?�?q翾���(>T��Y�=��+?\R?��(<8��>�t$?�Q*����>�Y>B�5>Y�>�9�>�u	>>���A�ٽ��?��U?W����>����y��eZ=z�>$�1�3ӼV�X>F@<Lg��S�W�9��:w�<�AW?<+�>G�)�����O��A3=�k{C='y?3�?rȢ>:l?�B?��<l�����T�I���+b=/�W?��i?"�	>-�z�Z\Ѿd���k�5?��e?Z�L>��a���� �-���Z�?6�o?k?�ċ��F}��x���		��4?�v?�q^��r�����m�V��<�>(]�>k��>R�9��h�>y�>?Y#�sG������Y4�NÞ?��@���?�;<�"����=�<? `�>�O�=ƾ�w��`���B�q=!�>g���cv����|S,���8?��?���><���ʨ���=+꙾��?�Y�?����	�<��"�m��p���<�ȑ=	":��+����77���Ⱦ��	���������ω>H�@�y�����>.>�u��o п��&Bپ�|��?碢>\��K-����e�m�`cC�+�E��������>�R	>S��zн�"�v��.��P�M�>�;��4�>�l}�@Ͼ#����T�=ظ>��>X �>9=��m����?u
���ο]&���X���N?~��?���?.0?�:)<+�u�$��i�� �-?�yk?��_?�-�:�,Y�[,L�%�j?�_��vU`��4�tHE��U>�"3?�B�>S�-�A�|=�>���>g>�#/�y�Ŀ�ٶ�9���[��?��?�o���>r��?vs+?�i�8���[����*��+��<A?�2>
���G�!�C0=�ZҒ���
?S~0?{�d.�@_?8�Q�hgO�z`�5wk��x�>	E��7)�A��3���-�f�b����K�غ?&��?C4�?�c*��7?�;�>�j��wξ8G��O>^�>�v>BzK=��>Ҿ�!��@�=��?��?��.?֫~�}����}=�3v?�К>���?��0?:.=������=is�>�M�>��-�he>?�%??r
7>��V����� ��z�/� �Y�T�g><V?�n,?Iu�>r7�=�G7=�+����Kh�+v�����Q�����>�)>�4�=hl�g�����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*�ҿ=����z������5�=��;fGY>
"��$	��z�>Jt=W$�=d�>�q<>�(>�K>͢O>��>7��>�V}��,(��M����~���Y���>�R:	���l�����Ǽ���ꦾɰ��q���b�b�ɼ^�r���5���r�L?�=��U?̦Q?J�o?\� ?��s�� > ���:!=�w$�݃=4�>�x2?�lL?�V*?_��=�ߝ�÷d�y4���S������y�>m�H>���>6)�>$��>	E���H>�>>.`>�>�
&=6���m=SO>��>J��>�E�>�C<>��>Fϴ��1��k�h��
w�n̽1�?���R�J��1���9��Ѧ���h�=Hb.?|>���?пg����2H?$���z)��+���>|�0?�cW?�>����T�3:>;����j�4`>�+ �xl���)��%Q>wl?"�f>Ou>�3�Je8�W�P�W|��hj|>�36?{趾�D9�H�u�s�H��bݾ$IM>�ľ>D��k�P������vi���{=x:?݄?5���ⰾx�u��C���PR>�9\>�U=Lh�==WM>xec���ƽJH��l.=��=��^>�-?�/>WB�=!��>�X���Q��k�>�sC>��->zB??��%?������=҂��|.��v>Q��>�d�>�>m�L��$�=���>a�b>�>�����#��*�A�(EW>�ɀ���`���r�-Dw=
�����=��=�� ��<�'(=�~?���(䈿��e���lD?R+?Z �=��F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��L��=}�>׫>�ξ�L��?��Ž5Ǣ�Ȕ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾTh�>qx��Z�������u���#=S��>�8H?�V��I�O�K>��v
?�?�^�੤���ȿ7|v����>X�?���?c�m��A���@����>:��?�gY?�oi>�g۾7`Z����>л@?�R?�>�9���'�~�?�޶?ү�?ZI>���?�s?�k�>�0x��Z/��6������Pp=6�[;�d�>�W>[���wgF��ד��h��r�j������a>��$=(�>DE�^4���9�=��I���f�8��>�,q>�I>W�>u� ?�a�>|��>�x=�n��Kှ�����J?Ñ?0&���\�Q��7��;���L�3?Y�/?�!�f�1���>نh?��?ӡ@?�XP>�v������пS�Ҿ��>�:�=�??��>�M�7>�h���GN���>7�>;�ʽ�����7�<��>�BL?N�?H9�>�)?f�?bP>V�>�^�V(���r���>���>�x4?jd�?]?�5���Y=�9����柿'�]����>G�?E�?��>50���)��Wf�<��"��p�����?18?�'_=�J,?hNx?~9n?��R?G>|
���
*�r���~W4>�!?M���A��]&��t� o?�[?���>�|�ս�	ؼB�������?=4\?�Q&?ʃ�]'a�pþ���<\�!��g_���<��F�T�>߶>�U��
�=�>�&�=�&m�f�6�Q�b<nL�=H��>ȑ�=��6������1?��+<m)w�±�=��h�|}7���>U�F>���f??�h3��<u�UP��UH��	�`�K�?���?%��?$'t��y_��'-?�%�?��.?�4�>����ZȾ����0�]��W��F��wb>���>�?��P�:͡�Xޥ�-wo��{�� ����>=M�>�!?�?�sQ>
/�>���ӕ&��$�����]�4��#8�tl.�-����%�%����������|��Ԙ>�~��	ز>p�?[�h>�6y>x��>
����>�PN>�>e�>�X>��5>�->��?<�oн@LR?}���Q�'����5����1B?�od?�4�>�i��������V~?5��?�s�?�Av>�|h��,+��k?)2�>����q
?�2:=���A�<WT��x��+�����+��>�D׽P!:�oM��qf�;k
?P1?�����̾�4׽#���M^m=U�?��(?{�)�H�Q�ݫo�d�W��S�����Th�Q8����$���p��㏿�a���"���(��)=y�*?��?�Z��t�,���nk�S?��f>���>��>V��>V�H>��	�>�1�n�]��S'�t�����>&6{?�ǋ>��J?g�9?�#P?�^K?���>qQ�>�ӭ��x�>v�e:0�>AM�>b�9?-?۫.?�?@�)?��c>����� ��پ1�?t�?�?�F?[�?�c���Ž�[������w��>v�r�=Z��<�{ս9큽[�B=P>+�?�
�K85����`q{>��;?��>���>��	�t�?�<{l�>�Q?�{�><�����q��9	��K�>�݁?�����<�&/>�1�=/�������z��=�ⴼ*z�=���/�W�CG�;=�=��=���:VF�9�a:�ر����<��?!�?���>
?!GҾI.�خw�y''�U
�>��<_�+>ֱ��V�u��T��s��U5t>�͉?ZR�?}'k>��s=U��=*���f���I�.���ȗ��Tt?"�?��s?���?d�=?�,?�==��#�!���L���"v����?v!,?6��>�����ʾ��ى3�ӝ?z[?r<a�)��z;)�͐¾_�Խ��>�[/�U/~����)D�������~��%��?�?�A�R�6��x�ܿ���[��b�C?"�>�X�>[�>V�)�|�g�e%�2;>��>�R?F%�>��O?�;{?&�[?jT>v�8��2��~ԙ�L�3��!> @?���?t�?�y?<x�>i�>��)�X�hQ�������8Ⴞ�V=�Z>o��>�*�>�>���=��ǽ�Y����>�Aa�=�b>��>5��>S�>(�w>�m�<�YV?|��>�:	�;I0��l��N��8S>��b?ˉ�?J��>.-���HF�V*���HξI�?�u�?CV�?�A6?�}>����=D�>|������=ڹ?�!�>�Km>_^]=?�*�t½R�?��,?��=�#"��n�3��m�	?m/s?�$�=����Y���9t=V�t�Bn�>� *��}��_�¼W�|���R�����x>ؓ��oVھ[N��������ܾ���Vt���5?hӽdbA>�G>�D">��>Kƺ=���=�Q�=3ZZ�%M�3<�����k�i�L����g�J�(.�=Ґj��_ھ�;�?r�?��?��4?_��>n�7>�2��#�>�[&�ȯ�>"�>�>Pon�a8�i������.sܾI�þۙl�Il���1+>@䧽h�c>0JH>�7=:����-<:�=�ͼ��>:�;C�;y��=�K�=7��=#�λ�Q$>�6w?U�������4Q��Z罢�:?�8�>{�=��ƾg@?U�>>�2������nb��-?���?�T�?9�?0ti��d�>>���㎽�q�=z����=2>r��=p�2�X��>��J>���K��Z����4�?��@��??�ዿϢϿ.a/>�7>�(>��R��1��\�}�b�e|Z�*�!?�A;��K̾�9�> *�=�!߾�ƾHx.={�6>�jb=�e�vS\���=�{���;=��k=�؉>��C>�p�=9��]�=ӽI=5��=��O>II����7��2,�ײ3=���=��b>2&>k?1��>��$?�?�>�0�8���ڱ=��>)%>�@Ľ�2>�7$?�ia?��B?��C?Iԇ>�OD>�w�>[X�>�N3����������>�ݗ?��?���>GQؼ�\�� 0��cC�@V�??�W7?�?���>����sٿ}�"�S\��"��]�ֽ�����T���+T>����;��>_��>�O�>Î�>u-)>�i�=)�a>=ϰ>˓�=b�=���=Cl�=0�<������=���=�����x�G=�ŭ<����8��:8	�;��J�{�ͼ��b����=�8�>��>@��>D��=0ﳾo/>������L��о=*ܦ�+B���c�~���.�jt6�'�B>
UX>f����5���?CZ>�?>�}�?hRu?.9 >�M���վ)E��B]f�YS�[�=�>��<�d;��Q`�r�M�b�Ҿ;��>�ߎ>��>�l>�,�2#?���w=G�b5��>|����j(��9q�@������Si�J6Һ D?�F��ܜ�=f"~?ǰI?_�?P��>��؆ؾ�:0>�H��>�=A�*q�Vh����?�'?���>�쾢�D��H̾9�� ߷>o@I��O���F�0�c��7ͷ�
��>
�����оr$3��g��������B�,Mr���>
�O?��?Y:b��W��8UO����O'���q?�|g?4�>�J?�@?�&���y�jr���v�=�n?���?R=�?w>���=E����>�/?ޖ?�]�?	q?�.?����>A�;�Z!>V*t�
��=o�>�9�=���=��?o
?z�	?#Ֆ��	�A�쾙X��Q�Z��=}U�=a	�>L�>�Tu>�3�=�w=�a�=�V>���>���>s�`>���>��>���v���k1?i�>v�>4-5?@Հ>��b='�ɽ�C��2��8�aH�F��3H��	���4��ڣ:?jP�R2�>,��\�?��T>D��^O?�T�K�h��W>]�]>WԽ�>�IJ>(�>��>�n�>�	">�ݚ>��">�FӾ�~>����d!��,C�3�R�t�Ѿj}z>�����	&���w���BI��n��qg��j�O.��e<=�ʽ<.H�?������k��)�����f�?�[�>�6?rڌ�A����>���>�Ǎ>�J��Z���Oȍ��gᾛ�?+��?F�w>�G>�Z`?Ц$?}D��큽�g��B����v��`��i�����S�i������V��N?�T[?Eb7?���<���>2v�?W�C�����m)D>+pC�`8V�Ǖ��Kn>���-��6۾�ґ��?>\��>�\�?�Hy?{R�>��'�������>.f?B�>Zx?\�R?">?_� ��n@?��!>�>+0?��M?޹�>�>�Y=�#�=P{�<���<�L��l����]�
�\���=�&>�<��弣æ����=��<�>E��<�������
Eڻ�B�����<�y>�Ķ>r�W?
y�>���>�,?������b��n6'?#,���~�G̊��ڠ����ǣ�=�Bp?��?߀i?s>x�L�3BL���_>�߷>P>�K>t,�>2�`�"��j=���=��Y>� >�<��A(������蠾6#6=��->Y��>�R|>7]����'>����8:z�Z�d>ݵQ�����2)T���G��1�×v�3E�>��K?��?�m�=龀��@f�%')?�f<?�eM?��?�8�=q�۾�9�H�J�[���>��<���ຢ�Q*���:�&��: �s>,���D���va>�v�@�޾$zn�Y�I�J+�sML=�y�H�R=S>���վ������=O�	>����)!�%�� ����CJ?�e=hä�|U��&��iH>SN�>�6�>��<�C�w���@��Q���,�=�.�>�:>�բ��&��G�S�Bf�>d5E?�_?nn�?�Ղ�D�r�*�B��A��$͢�$G̼�?��>�@?��B>M�=���"����d���F��2�>���>e��H��R��������$�̊>�b?��>C�?�R?��
?%�`?<*?�n?��>�H��.E���	'?X�? y_=J��o>V��_:��cH�^��>�%?8�H��_�>??��?�f*?�
U?�?ax>/� ���7�8Ǔ>/]�>�W�rӱ�/�S>��D?��>��[?�t�?u�>>Q26�n����&ɽ�?�=�F >U2?S3 ?��?iļ>��>䮡���=a��>�c?�0�?��o?1��=,�?�;2>��>���=Û�>��>�?XO?�s?��J?���>���<�7���7���As�t�O�Kۂ;pH<��y=��4t�H���<���;%j��1I�������D�<�����;o�>��z>���/>��ȾV�� A>ɍ�cM���#��Q�,����=�>�?	v�>>�"��ڏ=�><%�>qt�7�'?j�??�Q�;,�b�7Dܾ�kQ�8G�>;KA?a|�=�wm�Y���Nu�VDU=�l?
e^?Z�P���^�i?�V?`�J�%����Ě���Ɋ�,�m?���>p�<y?=ʀ?�W�?�
?[���f�p�����#�M��ؾz�=t̴>Z�	�F�N�\��>#3L?J��>=�>��a>�h�p�J��QX�uY�>[|�?���?�?ɿ�>7�e�v���+�:T����v?�J�>�o&���O?U �.G����������߾?8��Z��R!ݾ�b��PL{�_1���ݠ�W/*=�5?��]?K�E?S?G��OoR����h�_�"]g�b�+��+�9o�7lK���0���J�H���s߾�2��7�=����@I�6�?��!?�a	��p?���\���Ⱦ�M>@ٛ����Z�=����'=�%=��j���n{��"�!?;�>^3�>�Z@?=_Z�W_8���4��@;����F�>��>T��>���>r���&��Wֽ�9ľCsp�S�ӽ�6v>�xc?�K?��n?{p�+1�O����!�w�/��b����B>Nk>/��>߮W���<:&�Y>��r�X���w���	�n�~=X�2?�(�>쳜>�O�?�?�{	��k���mx�ʇ1����<�0�>t i?�@�>z�>�н�� ����>Z�l?Ώ�>��>�����`!��{��Pʽ��>n��>���>��o>�w,��\��k��˃��m 9����=Y�h?������`��΅>�R?1)�:�9J<fn�>�:v��!���򾁾'��><�?���=�;>�}žG(��{��N����)?�?8����h+�4|>�J?W��>V.�>8��?���>�3þ#�Y���?{}_?A�K?�2C?��>W:�<ae��,ƽ��'�47=���>��Z>ޕs=��==����Z����"8R=�!�=�ؼ]���H��;�Ѽз�<���<T�,>jܿQ�J�0�ӾZ��F�EN��/��h�����9A�0���A~�i�|�n�%��#�|z^�!�s������l��,�?K#�?ǋf�񉐾�v��͟z������>�/���Ƚ����w�J�wY��5�'��M_&�g�T�;~m���W�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >VC�<-����뾭����οB�����^?���>��/��p��>ޥ�>�X>�Hq>����螾w1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@NvA?��(������Y=���>"�	?��?>J�1��l��_���>��?�؊?�J=p�W��C	�S�e?�<��F�d��Pg�=ld�=K=���B�J>h��>����B�bݽ8y4>�
�>u"�Vc�H�_����<�^>�ҽN`���_�?�1N��^d�N4�|�u����=q�A?ޫ�>�|�=��?TD��.п�2`���f?�"�?���?}�+?��Ѿ&�>�oҾ�B?��/?%�>�8��<g���>x�Ƽ�m�;��ؾ[�N���= ��>%��=�8��t�'P;��?��Bh�=��wK���H$�!y�h<�=� �=<2���<��|μ�p���R��a��z�+=kh>W�3>xm>�>E>��'>Qn`?u	l?G�>��=U*��?[�9v��٨������}N�"��Jo��B���������T�ǯ�KX�ɻ��� =�w�=U4R�P����� ���b���F�b�.?�p$>��ʾm�M���-<�qʾ�ª��̈́��㥽U1̾��1��n��̟?��A?������V���Km�&���>�W?R����z��=����x=k �>y�=��H!3�{S�	*?�M-?�tܾ0�j���/=�S�V_=C�7?\�?D�<c�>��?��X7��+>��>9�>��>QQ�=Nz̾�ø�d�?��O?O��[Х��׎>)Pؾ���c�%>���=��P���<�*>�uL��҉�=#e���m�=@�W?�'�>e�*�������i��JQ=@�x??��>�m?��B?9<=.<��^vV�:��TL=�V?dsh?y:>w���a־�$����4?�Mf?v�=>WU�	-��.��+ �r�?��o?O�?M�.��{�p�����N�-?��v?�r^�os������V�f=�>�[�>���>��9��k�>�>?�#��G������Y4�Þ?��@���?��;<Z �H��=�;?k\�>�O��>ƾiz������U�q=�"�>����pev����R,�P�8?Р�?���>𓂾������=͖��s�?p�?yͩ����<�#��#l�H���C��<&j�=<����"��!�U�7���ƾ��
�󌛾�|ü]i�>?U@����>Dq8���97Ͽ�9����Ѿ�Is�^b?��>�ν_�����i��,t��F�lzH������w�>��>�l���摾,�{� n;�lϦ����>�	�L��>7T�ha��ԥ���F<je�>��>�ǆ>p���	u��'��?��M0ο����:���`X?�J�?Ev�?͆??z=<FXw���{��C��G?�s?VZ?_#&��{]��#4�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�q�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.��^?]�S��k�ݬ���u��I�>?s}�����s�ܽ��B�U�]�lT��~�ԯ?qU�?e.�?v����?Z�>��{��9ܾ�֤���>`�q>{1%>!3�<cȞ>����=�Ў�=�t�?���?��?�{�Ġ�Z�=h��?V�>v�?�~=e��>n�T=�uľu$=��V><d>/S���F?�C?r��>~�>JE���'���2��;A�El�E.J��3~>�]?�JF?K�>����d��D$�ʃ��O(
�OS��JX*�@�����x�>��,>F�>9:��`����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*1�п_���w��6�����=���=�u>������=̄�=�o���U�=��6>���>��_>�J>��5>]�*>_%>|���&�����爐�݌H��������2��Q� �
 Q�k���ҝ�����'�������ҽ?q�j��`.�(k�=�wW?�*O?%p?�G�>ʵ�� �2>Ǹ���w==���L�=b7�>'q6?�tL?�
'?^�=f����b��R���	���m��Y�>�&I>�C�>f.�>�.�>�,Ż�j>>f\.>�k>�)>�lC=��ɻ�p=ؿP>5b�>9�>P�>�C<>��>Dϴ��1��h�h��
w��̽/�?~���R�J��1���9��ڦ���h�=Ib.?|>���?пa����2H?(���v)��+���>z�0?�cW?&�>��u�T�8:>C����j�1`>�+ ��l���)��%Q>sl?:"g>�2u>�3�4m8���P�����|>:56?�����j9���u���H�Ğݾ<�M>��>�=5�+6�����]�~�+Si���z=�s:?ƚ?z貽 ���_	u�5H��z6R>�\>�z=L/�=O4M>e$d��Yǽ�JH���/=���=0^>ܑ�>�,�>��}�Dհ>�%���(��k�>���>��>�.G?P�@?�4��9=!�-�A�K�� B>_?�>��x>\<�=53����j=,�?�ko>�Ɛ=d�
��`���}���5>O�c=�쉾'�\;z�=N ��䑾=��=�����i��`~=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿk�>�s�<Z�������u�g�#=$��>`9H?�W����O�O�=�lw
?+?_����T�ȿ�}v����>O�?���?��m��A��a@���>͢�?5dY?�ui>�j۾fcZ����>��@?a	R?$ �>G7�"�'���?�۶??aI>���?�s?�k�>�0x��Z/��6������p=<�[;�d�>�W>f���xgF��ד��h��u�j������a>��$=,�>RE�[4���9�=��I���f�<��>�,q>"�I>W�>v� ?�a�>}��>�x=�n��Jှ����Q�L?�2�?��$��V��H�qq�<�ˍ�@�<?[6?o�r��Hݽڶ�>9�`?�Y�?T<?C�F>��7�����Ϳ!־���=]�'>���>W�>��#���<�׾�+:=�V�=IO�>�k%��Q
�;���Gd�<���>��.?���>���>�,?�?� >�a�>��r�8 ����� ��>>�>ɀG?_S�?�?�F���6��������֛b�-ߤ>>w?��?Fsf>nȾ���B��u���I���<�?�!?7����#?CL�?��]?��G?�jW>:d� �&��L���Q�=lg2?����|�M���m��2%�B0>���=�S�>��㼒�>��ہ��c��(���*?7a�?v�u?���mk��,>�N=�9�<��_!=8%W=�>�.�>4��=X�3>@��="�>r팾9���a�B�H��;�od>�ND>y�|����'=,?��G�%ۃ���=��r��wD���>�FL>B��K�^?Im=���{�{���x��D
U�� �?��?gk�?D��;�h��$=?��?�	?Q#�>�I��|޾��ྯSw�<x�Qw�%�>v��>�l���M���)����E��.�Ž�Ձ��>���>���>P�?=I�>�s>������$��{�L��yM�c�)���J���1�p�*���Ӿ�Y��D��w���ǝ��;z�>Q���f��>g�?4U�>�i>��>�=�>�6\>=��>(p�>rb>�A[>�V>�n>`��KR?���e�'����ݰ��B?Mmd?�h�>8 h�����ܡ�#�?��?�q�?�.v>�rh��'+��c?��>�.���p
?�8:=���6�<�e���������e����>�ֽ�&:�M���f�a
?�2?�̋�4Y̾�_ֽ�R�� w�<��?$�?��&��uC��s�#�Q���O�rn��Q������4�%�l@w������r���<��2]2�1lo=��.?W6|?��H���#����g��>�=ڃ>�k�>Lً>� �>}��=7��Υ2��^�i�,��m��ڟ�>�jv?�uG>�Y?)&"?W$Q?�2+?�O0>��>⺂�z?w@>V��>>j�>�V?b/?e?Dv�>1�$?3>h��A��C�ƾ��?��?E?��?�m?�����`5��ֽ[9���^�=�71=U�-=YO��{o�w!�=9�F>�X?���ɬ8�����Nk>k�7?	��>y��>���(-��J�<w�>�
?	G�>E �"~r�c��V�>���?���7�=��)>���=\�����Һ(Z�=������=�5��(z;�+e<z��=L��=;Mt��&��5�:��;sn�<�� ?O1?�ӄ>Y=�>��^�_��ed��̢���=�o�=�O�=+�ľ�cz�O]��0Sv��/>'B�?g&�?�D�=1�>�><D�������-h]�.����=}�?N�F?�>�?��? �?k�6?pO>&/��E�����p��Վ'?i!,?��>���*�ʾ���3���?�[?T;a����Z:)�B�¾��Խ+�>�[/��.~�k���D�{.�����n}��͛�?ȿ�?�A�n�6�y�п��=Z��^�C?�!�>�W�>��>J�)�V�g�%�$3;> ��>�R?$�>>�O?*<{?��[?�gT>b�8��1���ә��[3���!>�@?���?��?�y?�u�>��>A�)��ྮS��w��s�ႾK�V=�Z>��>`(�>S�>���=Z Ƚi]��)�>�=a�=݋b>���>��>7�>߃w>$`�<A�I?���>��ľ����G��M�����j��os?kc�?�#?o��<a%!��]J����Ux�>al�?�T�?�?�}/�׫�=3��������K���>e�>��>��`=T�6=��>���>ƃ�>���0��@�8�DΖ���?O�C?Hq=�������5�.=�s����>Pڼ�N��(�$�E�K���=+�ľ�{Y��44¾9����ľʗ���Ͼk�D����>ʭ���]>n�>_>�K�=�~�<�\?;
̼���<4P-�*��� �Ǽ�ʾ�yV�2<=�=4x^�tjӾ�Ā?MA?~s.?j�;?�ip>�uf>0�Pb�>��S�,�?W{j>i�=���APB��ߧ�c8����Ⱦ�hҾ�By������=>}<c�W�'>��]>��
>�;�2�=@�=}y�<�bL<�w�<�+�=���={$�=`��=WR><�>�5w?����ﱝ�n.Q��G罔�:?.�>�B�=j�ƾy@?�>>^2��?����\��/?���?YS�?}�?�qi�9g�>�������H�=/� %2> ��=)�2�q��>c�J>��eI���i��t5�?>�@2�??�����Ͽps/>� 8>�`>$�R���1��\�� c�9�Z���!?�!;�dO̾==�>���=A߾�:ƾrp0=�7>��c=ú�	+\�ʛ�=�{��<=y�m=aى>2�C>}�=ӗ��[+�=	�I=#�=$�O>�����8�A@-�:�2=�o�=5�b>��%>�% ?ʚ?b�?ȪE?�x�>'���q�,� �>�Q)<vQ><y��N�>|G?T�Z?�`?�H>?�>�=P>�w�>CW�>A�)�&&�����k���<B�?"V�?K�>�w����f�}���u#���ּ��?�w?x��>0��>e��sڿ�O-�)�%����;K��=�.�=��48=�n<A�����=�8�=R��>�R�>Z9�>WU>�#6>I�	>,b�>:�>���=���=E;�<>)�=驽��<��%���4<�?���˻X��kZ��I�<hx�<[<�ʼ�CʺH��=���>M>WA�>���=ҷ��YY/>C(��A�L��1�=�f��%�A�d��J~��/�H�5���D>ʌY>2���*��n�?b�Y>�	A>�y�?�=u?�!>��Si־/?��J?e�JR���=�>*?�.�;��_���L��gҾ\��>�ߎ>��>��l>�,�^#?�3�w=��b5�'�>�{�����'��9q�@������[i��^Һ��D?�F�����="~?��I?R�?N��>N��x�ؾ�90>�H����=��	)q��f����?�'?I��>쾴�D�;I̾7���߷>�AI�V�O��k�0���`ͷ�R��>������о�$3��g������-�B�ZOr���>�O?K�?�<b�QW���TO����&���q?�|g?�> K?�@?T&��xy��q��pv�=��n?���?$=�?�>'�=�5���x�>`c?��?<?)�r?�m>�U�>�˸;��>�-�����=��	>I��=6K�=^�?�G
?A�
?�����
����*��7�]��N�<&j�=ꢒ>�>jt>�K�=+�l=\o�=Q]>�F�>���>F�f>���>I��>��۾�d:���R?O%h�g�?{M?�N>���=;�I���>rv(�l|
�Ö���E�;��ަҽ�����<��ɻ���>�跿E�?��2>����
?�����8R;]��>l��>�>��>��>ע�>��>��>��>9M�>��=\Ծ"�>�����!���B�	uQ�MӾHy>�Ϝ�==(��	�4���J�l2��cd��&j�sj����=�v�<�D�?� ��Ej�ۣ)�WT��o�?M�>�W6?Y��T�])>���>n�>���ru���ύ����[�?-n�?�es>��1>tO?'�@?�������h�0�����s�|�u���K�ˤ��Ez��'�d�H<�.Q?�i?��=?���{�>�H�?R�v�u�j�`i~>��S���@��%���#>����G)��ؾ3׾�;>��>4 �?�'x?j��>�������Bhy>�g/?�1?|)g?�V*?o%U?y��(?�NG>�<?o??��G?��%?R&�>��>1��=��';�%=�Խ��q��u����#��,n<1F�=?O�=��~�rX�M�,=>@���<r���r����c<R�<2+�<.�l=���=s��>�ZX?�{�>a��>O�<?�@轔���0ξs�>�ƽ3����{��D���"���=~qY?6�?�Ws?�h">�d��*�)`>P?�>�J>EO]>���>L����V��7=�,�=B->oq=��ͽ0�������d��B>�2>'U?"�>S���>>�oj��ω�&'$>�Sf�L����<��.�9���1��¾�ۗ>k'<?;
-?wC�>��˾�霽<\���?��:?=Us?Գp?o�>�W���X��xa�K����3>���>�������q�N�r��X�=��?pX��䠾kkb>A��"p޾�n�J����reL=�s�n�V=k#�P�վ��~�
��=r#
>:����� �u���Ҫ�i$J?�3k=Q��#U�/`���>6Ø>9Ȯ>j�:�^�v��@������"�=O��>�-;>����i�yG�,:�s>�>�RE?pV_?�h�?�$���s�L�B������`����Ǽ,�??y�>�h?�%B>���=���M	� �d��G��>��>����G�k4���-���$�t��>8?1�>S�?u�R?;�
?N�`?l*?cE?Y'�>b�������A&?7��?��=��Խ�T�� 9�LF���>z�)?�B�˹�>P�?�?�&?	�Q?�?m�>�� ��C@����>�Y�>��W��b��N�_>��J?ܚ�>j=Y?�ԃ?��=>\�5��颾�֩�&V�=�>��2?6#?K�?쯸>k��>O���䜀=8��>��b?�0�?��o?���=��?�%2>κ�>T��=qm�>{k�>u?�^O?��s?��J?Ā�>M�<L���$���cs�}KP�A�;�~I<��y=B��t��'�Q��<�c�;�D�����M����D�h������;�_�>D�s>J
����0>c�ľ7P����@>/���P���ي��:�9߷=/��>��?��>�Y#�o��=���>�H�>d���6(?��?�?<";ǡb���ھ�K���>=	B?���=��l�����+�u�{ h=��m?��^?��W��&���P?��\?�����4�}���,�p�E?��?(���@>hf�?�n?!y�>Hϥ��G��RN����S�CN�g�6�[�>��9�^�_7�>E�0?:|>��~�l����rm�Ѐ��ʃþy�?Am�?���?�hZ? 4�=�2r�6�ٿ[�k���}�e?���>����2?��V�ㆷ�B�������5���B���9����9��@c���2��_���ܽ�=Di#?��\?��d?W#>?����Mo���n�%�{���W��-˾S��c�Q��{E�1�I��c��|�e���6���N�-=����1M�m[�?s�%?��6�$�?�����ܾ�꾲�>"φ���߽m�=+(h��|�<C�=>Nz�#10��糾'n+?���> 4�>��(?�5T���A�!b?��,3��g���W>�~�>a0`>�	�>�x:�%5/��z���˾�o��`��Ov>Q�d?��J?��j?5�S12����r&"�P�&��-����.>n�>���>�I�s;��C(�F[?�Vs�Ee�AD��\��H=�1?��>[Y�>?�?ߖ ?�^�͠��;0x��61���[<�Y�>�i?A�>iI�>EbԽԐ ��6�>�Ll?�R�>�0�>����7"��)|����q��>6��>] ?7s>S�*���[�԰������&i9��t�=��h?����H ^�0��>/Q?~�l;�	V<[�>&���w�!��3�F-�1>Z?s��=0I>>pBƾ3o�"Y{��N���f)?�/?`F����*�a�}>:"?���>���>�#�?m�>��þ����J6?��^?��J?gvA? ��>��#=����Ƚh�&�a-=hT�>^�Z>�Ek=e&�=(��	�\��5��+E=Z�=�4μZ��]�<pz���KF<C��<%4>C�ڿ�K�sоcD��,�T���Ԃ�9lн����-	������v����o��>��9.��V���g�ԙ���#i��N�?�b�?�����f����jw�4D���V�>T�h�⾴��;���<ڽ/E��p�־9W���z ��P�Og�b�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@}A?�(�����V=9��>$�	?�?>�S1��I������T�>u<�?��?|M=��W���	�1�e?(< �F���ݻ�=�;�=�E=���ҔJ>|U�>����SA�X?ܽ<�4>Kڅ>~"�Y���^�<��]>U�ս<;��OB�?�TW�P�h�%�3�l�}�((>]U?�p�>�Y�=�$?�H��tͿ��e�R?�|�?P��?Z1?b$����>uܾ�SE?�1?c7�>�q$���s� ��=\�����R�侙0L�zL�=Q��>�8>��?�>
���V�T�-"�=ј��&��f��>�Y�v=�e{=�Mq�"�s��	������u�ނ�������8= �=[�;>��e>��>ObN>��S?@\s?�Y?�Z�>gbj�"`_�$վ�= T9��LA��~u��E��4���r�վAEȾ�9�l�%�9�{���!!=���=�6R�_���<� �J�b�B�F���.?�v$>R�ʾ��M�R�-<gpʾL���܄�D᥽�-̾�1�"n�k͟?��A?������V�c��>V�j���^�W?P����ꬾ֤�=꫱���=%�>���=���� 3�~~S�T|0?jS?C���Lw��"*>�� �B8=��+?х?cX<0�>�5%?�W+����[>R�3>t�>��>y%	>}��Kc۽��?G{T?���P���А>�U�� �z�/ a=J9>L35��=鼱�[>AƑ<N�����W������ּ<��V?�D�>L�)���e���-��E��˄?��?��z>�$~?{�M?�x=~��sUk�Y��/��;pF?-q?���=��q������%��WQ4?$�L?cּ=�~���3Ѿ���m���?z�~?=_9?�Sa�����z��=E��'!?��|?�E�������5���|9�>�K�>E�?I�󾇭;>rh?~���ݡ�p!�����%�?��@m��?��ؼ��m���X����>	r|>r����`n�C�z=И�O��!��>����E�T���4�0|��a?�h?��>��:�����="ʗ��g�?w݆?J���}��<�x��k����ޚ<�Я=a����{��7�3Ǿ��
�������м�A�>k<@U��~�>�#:��i�D$Ͽ����Ͼl��O?V��> �н����j��Eu�[�G�5H�M��mN�>E�>��������E�{�hq;�`-��K�>��K	�>�S�D'�������n5<��>��>w��>f%��v彾(ř?c��=@ο2���Ν�9�X?h�?�n�?_q?�g9<��v�l�{�k��h-G?��s?	Z?#_%� :]���7��j?M_��cU`�Ԏ4��HE��U>p"3?�C�>��-�ǯ|=L>���>Xg>�#/���Ŀ�ٶ�����(��?ԉ�?�o���>[��?9s+?=i��7��(\����*�K:,��<A?�2>������!��/=��ђ�S�
?�}0?j{�v.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?L�>(H�?3Q�=$�>��=���������>��=̺+�� ?uM?�#�>���=ô6�V0���F�*�R��H	��D���><"a?]K?�5f>_x���%�1i"���̽1+�w��}D�	�5�e)ͽB�:>�{?>�>�qG���ԾZ�?A1���ؿ$_���(��4?M�>%?kP�k�t��z �D�^?��>cL��(��O���?�J��?�`�?H	?�z׾��O�>펭>U[�>��ӽ�ĝ�-����n6>J�B?�$�Q����o���>�!�?��@��? �h��?U9۾cѐ��(s�8�m ����<'�E?�[��a>��?��;���z�>b���s�Fz�>;ȭ?�N�? 0?L\?�r��7V�.H�tq�>�r?bc?��K�q־�	�<1J�>���?���~X�� p?��
@�V@�v?t6��|hֿ����7N��4������=���=͆2>��ٽ�^�=��7=��8��;��1��=u�>��d>	q>(O>ia;>�)>���O�!�r��Z���J�C�������Z�K���Wv�Kz��3�������?���3ýy���Q��1&��?`�8JH=��W?nQO?茁?>/?�˰��A�>�;�:�߽���>n	(�M�?C�??.�m?��8?x�=����r�b�l�|��_�\�;��t>X�>��?�X�>���>ߵZ=R��=H;�H�>�q;=J��<��A���ڽ��>x��>ɝ�>`Н>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?_�f>&Nu>g�3�xf8�U�P�����'|>�#6?�ܶ�k9�O�u�äH��IݾNrM>ƾ>/jH��r���������i���{=�q:?Ā?`����ٰ��u��^���FR>�f\>�
=�=�=M>�1b��Lƽ��G�Ƙ.=M��=P�^>vX?�+>բ�=�ۣ>e��6BP��>�B>�%,>�@?�(%?��G痽������-�Vw>�U�>e�>�\>&\J��=:m�>��a>BI�˃�V��C�?��uW>,~��_��lu���x=(3��n��=� �=� �9=���%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿeh�>Dx��Z�������u��#=$��>�8H?EV����O��>��v
?�?�^�੤���ȿ'|v����>c�?���?P�m��A���@�m��>.��?�gY?�oi>{g۾�`Z����>»@?�R?��>�9���'���?߶?ǯ�?uI>���?�s?Ak�>�3x��Z/��6��󖌿�p=0�[;�c�>X>����gF��ד��h����j����)�a>�$=/�>�D�&4���;�=�񋽑H����f���>�-q>��I>�V�>>� ?�b�>���>iz=n��nှҸ���:?��?�/ݾ6We��N�??�������ʩ>s$?H�*>#���H�>��X?�և?9l\?���=� �g��r^���|Ͼt��A	7>Cz?��?����	�>��qB���>�!�>�����������>*��>��?8�>��o=1�%?��?��>�>�WZ�:��S�;�đ?�]�>���>Ν�?��?@����R9��$��tܛ��P���>�T�?{?�(>����ٌ�9�3���t�������?�|~?Ж��x&?���?O[?\m?��=����NW���88�>��!?i���A��P&���]�?�R?���>I/���ս��ּe��ҍ��Y�?�.\?�D&?����a�w�¾��<O5#�fhU����;��D�׵>��>��y�=�>��=�Qm��?6���f<�Y�=�|�>���=�57�\j���V@?�m/�H��Q硽ICZ�Ǝ�{�>yѫ>�𷾽y�>g�����WD���N����w��?��?Yל?���#Rk��0?��h?T2#?���>�S�X;����]Û�,����8���=��?�L=�(6��ա�=g������n=��g�>���>�?�{ ?��O>L�>�5��('�||�v���^��o��q8���.����kˠ�8#�����D¾��{�I�>ʂ��G�>n�
?^h>��{>�>��ʻL�>�/R>e�>�q�>4X>e�4>ޑ>�<��н�KR?�����'����Ҳ��M3B?�qd?E1�>i�1��������?���?Qs�?	=v>h��,+�on?�>�>^��Yq
?�T:=":�Z<�<V��f���3��Q�H��>~E׽� :��M��mf��j
?�/?���ċ̾6<׽�|��<�Ľ�6�?��?ޤ(�t�(��x{�YG�.r�.�*����]n��yF���[�/|��� ��D`���	� �z=�I?�&�?$���#�Tþ4·��3���R>��?���>�ޠ>��1�"�+��eE�"�V�cY�����$?�Ǖ?p=�>M�F?y*=?�@[?�rT?⾇>�6�>H����>iJf<��>}�>f�;?	F/?S,?Lh?;�%?�l>>�������ӾI?$�?�!?�p?�?-m|�7���!����P����9|��Z=�RC<+�ͽ��=���=�UN>�X?���ɬ8�����Rk>m�7?��>z��>���(-��B�<y�>�
?G�>F �#~r�c��V�>���?���1�=��)>���=q�����Һ(Z�=������=�5��(z;�Ge<���=P��=&Mt��'��_4�:2��;nn�<�?�?�Q!>�9>�Pr���v�#�q:>�=��%=0��=,�u���F���]�g��>>7r�?q��?m�>���<���= �a��߾��6�9$	��O�=�K(?��.?�eN?q��?�vk?��=?��%>����9������,���\?s!,?+��>�����ʾ���3���?{[? <a���i;)�=�¾��Խ�>�[/��/~����0D�煻����~����?Ϳ�?`A�2�6��x�ܿ���[����C?h!�>Y�>��>��)��g�q%�1;>���>R?��>��O?h2{?"�[?�cT>��8�%���ә���2�A�">��??!��?��?Y(y?`��>CL>5*��:ྍ���������/΂�h�X=��Z>C�>�N�>���>9}�=�!ǽ|���>��e�=ȅb>ڙ�>๥>��>g�w>,�<PR?ޖ�>L����� ��Ӳ�Y���W=�|?r��?ҫ?�M�\n"��%j�ї��?"�?�K�?�Q?�n����=I�o�^���������>F��>?��>R;�=���>i��>��>
���m���ԃ����>�(?���=]�ſ�p��;[�	���Z4<ە��d�T��ɹ�!�X�窓=�?���]�W��w�U��֝�M���"ӷ����v��?��=�>F>�P��:�;,p�<��=��<&���K-~�L�[=���<<]��FVO��<�ǉ=QvB��u˾�_}?#jI?�D,?�vD?�Gz>$>>�69���>����/?s�V>��H��D��J;�̹��ɛ��1�ؾ��׾j�d�:l��1�>XEM�%�>�5>���="��<;P�=`s=��=&���_�=Q�=���==�= 0�=d>�7>rBx?$U~��S���yS����S�<?c
�>F+�=����Px8?@�'>2V���|��'��l�?"��?c�?��?�no����>�@�� �{�n�[=	ᏽ�.>RJ�=��&�[�>-�S>X��b��oEĽ���?��@-�9?�Ӊ��˿`(>�W9>X�>��R���1�=]���`�K�X�5�!?��:�R̾�L�>Gs�=ԟ�{QǾ]�<=�8>�n=`��.+\��t�=!!}��5<=� k=}U�>�`B>���=į�M̴=��G=���=O�N>1j��Q�7���.�"�2=�!�=lSa>�8&>u��>z�?�a0?�Xd?W6�>�n��Ͼ�?��SI�>��=F�>c�=�rB>��>g�7?��D?��K?��>7��=v	�>��>X�,��m�wm従̧�O��<���?�Ά?.Ҹ>W�Q<�A����g>��/Ž�v?QS1?�k?��>�8����;/��:�i��=�o�=��>><´��Nn������a��!����>4!�>�Y�>=ɢ>L7.>�I�=a�>d~�>f}>	��;�@�=��Ѣ=�=E=�g�~�� �=�*�=��=@�㽒].�����<$�=`��<�):�~��=.��>?�>���>t��=$�`.>D���7�L�a(�=�d��@=B�>?d�W~�8/�l%6�E,C>�fX>U���&3����?4Z>*?>"m�?��t?#x>�����վ/���ee�RZR���=�w>6=�ơ;��d`�[N�OHҾe�>mN�>r�>!k>�;,��?��/i=mh��Z4����>e͋�nC�J!�rp�p6������Gi��2�&JD?�I���u�=_�}?��H?�ȏ?���>yT���?ھ�->�A��,q�<����n������y?r&?�a�>�s쾞E�Z��ը1��'�>\?���yN�f)��$:���=�I:�n��>9�+�
��ъ+��%��1���:��Ò�j��>���?�q�?�9�:n���\�Y�ɮ���ý�`?ls�?2�?��>�J?s�̽R��R�Ͼ��n=��?Qy�?,��?�#�>���=�
���>�>u.	?r��?���?�s?p~?��w�>��;+� >����8V�=��>"��=�2�=9s?2�
?P�
?^p����	�������#^����<ӡ= ��> l�>�r>��=�fg=�s�=�.\>?؞>N�>U�d>{�>]R�>��־K#�$�5?�ak>j� >w�W?�>�J=�;%�����]���(��o��ܞ�{F ��1��=�ԽR�&����!(2?i�ÿ���?�_K>H����#?�Q���>-�=k�c=1v����>��>Xo{>�>�z>��=0Ǫ>y߾=UFӾ�|>P��d!��,C���R��Ѿ{z>`����&�ٞ�gz���AI�>n���g�Vj�>.���;=�>�<�H�?�����k�/�)�����[�?Y[�>�6?֌�W����>���>�ō>�J�������Ǎ��f���?.��?�;c>��>G�W?�?ג1�23�vZ�+�u�n(A�-e�V�`��፿�����
����-�_?�x?2yA?�R�<(:z>R��?��%�[ӏ��)�>�/�'';�@<=t+�>*��0�`��Ӿ��þ�7��HF>��o?;%�?tY?>TV�a�߽X5�>P�U?`e?0)�?(�=?ҕn?��T����>�F>� ?�i�>ի<?��8?���>Eqp>Sl>0��& ȻY2�� j�u#��#}Q�ARڼ��(>��=q?�=��<���=�0���E���@�!r<�ļFD���J;=�{>��N>��>4�]?;��>�F�>6�7?7^�PK8�<l���#/?k�8=A͂��6���0��j?�[�>�	k?	�?�Z?�d>�A��C�<">�5�>KN&>N�[>�r�>�1ｾ�E�l�=B>�T>���=RM�������	�����0.�<*>E��>�0|>��Z�'>Y|���0z�£d>��Q��̺���S���G��1�C�v��X�>��K?��?L��=�^�+��If�00)?�]<?�NM?��?F�=��۾[�9���J��=�q�>Yc�<F�������#���:�]��:�s>�1���ʾ~�b>c�Ͼ,�d���Z�a�5�dcԾ��9�T�M��f=7z���d3���$C>��L=�����.��v��7���PFP?��=!P���b���W���Dt>���>��>�&7=𙚽��+�������>Mv�>�o�>��=����$�C���Ȇ>�E?��^?f�?Ļ��ar�zC�����!����jɼR?;��>�.?&�@>� �=||���|�5e���F���>5��>���O\G�����~J�i&$��Ɋ>�>?�J!>��?�.R?�?:a?b�*?��?$��>-��8_���A&?8��?��=��Խ��T�z 9�MF�]��>f�)?��B����>F�?�?�&?�Q?ٵ?\�> � ��C@����>iY�>��W��b��e�_>��J?㚳>a=Y?�ԃ?��=>T�5�ꢾ�֩�[V�=�>��2?6#?F�?ȯ�>o�>p6}��� >S��>a�H?�'v?�s?�y
>�((?��!>��>Y�>ˌ>���> G	?=�a?Kj?��??���>�{��������C�+����'��O����(�<�*�sk=V$Q=Q�p�;����i���s��򷽋�ü�
a��_�>��s>(
��u�0>��ľ�O��%�@>1���P��Eڊ�W�:��߷=���>��?;��>EX#����=��><I�>J���6(?��?�?w�!;��b��ھ��K�3�>	B?U��=��l�������u�w�g=��m?��^?�W�U&��Y�W?��v?0�ھ �:�i��x[`��&�9e#?48
?��!���l>��}?i�]?���>�"�'�a�����bo�ɂz����=E�>�֪�JP��]�=V	?_��>TIZ>v�u�U2���_���Ծ	:I?8�?g��?��|?�*>b�i�\߿������`U? ?�p���D&?ɪ7�ߌؾ�Ѯ�Љ�V��\�}����4�w�����D$n��s�]n��-=:D,?-�_?I�?3�k?���9�a���p��L~���i�8Ѿ������H�?�-���3��.z����|�w���ż�����N?�"�?k[,?��:���>bӖ����@��EA:>\���x9��b�=��B�;��FAo�C!A�0a���l*?�	�>0\�>K?%�N��a4�Y�0�G@��u��!?>�,�>b�w>�v�>x.�<�L��&���ؾز�������>�xj?�>F?'"^?��b/�ߋ��.0�0�,�ٛ��	>��>٣�>
.����Z�&���D���v���X���>��G�=S�)?�D�>�'�>�ݕ?���>	�@�{�	���5�8�L�m=��>}gx?���>��>�%ý+��f�>��q? G�>�T�>�w�.4��J���P�'�>.�>���>=�>��R�!Ec����掿�=��
�=�^c?�N��?#U�-�>�`G?��$����<�L�>Iu��m���jھ����f>��?�L
>��e>�ѭ�����'���p���:(?5�?�,��]+���>x�"?���>Y[�>��?ʗ�>����C�H;U`?Q@^?M�I?&A?z��>�=�﫽�,ɽ��&��)=iC�>,�Z>�!q=��=���	�Z�q ��zB=��=�UǼ�I��[[<�Yü��g<|��<��3>��ڿcL��#Ҿ?8���f	��>�����4���L�PQ���怾�`���3Ya��"�+\��U���|��t�?K�?F�e��(�\����ou����\t�>ҥ������[��w�<�u��C�Ͼ3�ʾ7�*�t�Q��vk�u	g�Q�'?�����ǿ򰡿�:ܾ/! ?�A ?8�y?��8�"���8�� >�B�<m-����뾮����ο@�����^?���>���/��k��>ե�>�X>�Hq>����螾~1�<��?3�-?��>Ďr�1�ɿa����¤<���?/�@}A?�(����^V=L��> �	?��?>oT1�cI������S�>q<�?���?�uM=X�W�;�	��e?r<��F���ݻ��=X>�=�C=?����J>5U�>h��oSA��<ܽ	�4>\څ>&u"�����^�'��<V�]>��ս�=��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=7��I�ƿ� ����dލ�_��-=h�z������f�������픽��'�@�=�e�=��>ya�>z|V>�U">�Ud?��u?���>2o>��ֽ[����ھB\��Ⱦ�eR�?�н�¦�?'�C� ������K�	����=��&�=�6R�ڗ���� ���b�V�F�K�.?Ay$>��ʾ�M��.<dsʾŪ��ꄼ%�01̾ї1��n��˟?r�A?����U�V�%�#O�.����W?�M����款Ȫ�=�7����=�)�>홢=J���"3�S�tn0?gm?����f���^*>� ��=�+?�?�PX<��>�Q%?R?+�*�TE[>�J3>���>E��>y:	>\#��=۽_�?�kT?
;�K㜾���>�y���z�R]b=�m>�4�|o��)\>:�<㼌�RZV�O��y��<�(W?x��>�)���c���[==v�x?��?�.�>[|k?T�B?%��<�i����S����tw=��W?�)i?]�>w����о������5?g�e?��N>ch�.��A�.��U��$?=�n?`?ԏ���w}�������!n6?���?z�S�y��Κ��[���}�H;�>�G?�C-��>穈?������YBտ@lM�U4�?��@���?(�>�.���=Em?��>)֖�x�\�y(%=�{���<x��>P��F�����D���&?j5�?HJ?W)����>�q�kc�?�n�?[.���CF=�!�s{\�]R��/�=���bB��N���:�ǒȾY*�e;���\n�^�>�0@�	��tt>����t����ܿ>_z�3��M�R�=t-?L��>���V�޾K�m��hn���V��[R����ݗ�>-�>��p�t����w��5���	�cR�>Fӈ�1�>�+O��C��s*��&��<�Y�>B]�>\�q>�X۽��þ�{�?����˿����'��"s]?~ʞ?<�?��(?ʛ˺G�|��r������<?�	t?*V]?�H��J��={�[�j?�`��'Y`�ʎ4�>KE�,U>�3?II�>��-���|=$->
}�>U>�%/��Ŀ�ض��������?5��?:n�8��>ˀ�?hr+?j��6��(T����*��2�X?A?�2>`�����!��/=�
̒�>�
?%�0?�j�-1�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?C%�>1�?WJ�=(X�>���=���=/��X#>�%�=��>��?V�M?.9�>��= �8�*!/�I\F��FR�"���C� �>��a?�|L?�1b>���C52��
!��eͽ�M1�����C@�N#,�Z߽�>5>��=>{>��D��Ӿ�3'?����Eݿ�����0o�N:?Q�Z>��?t��un�O�?=tI?�c1>���"귿�Ӎ��[����?3��?e�?Hr�@ �$�#>Eݍ>��>�_#��EO������h�>�L?����ӎ���g�o�>���?�@V��?aZs���&?؆	�po��Vps�u�6�Y�Ⱦ`]=��[?����66�>��/?�!��!�����������\>e&�?Ut�?�O?�mB?��f�i
���=�+9>*]E?��?��=�|	��S�>U�%?��4�p����*�i?p
@
@s�f?*���'�޿v��]z����ھ:y�=��=��:>sIƽ��d<����YGY���R����=[�>־o>%�q>�E>�O9>b�5>����������������J@�uZ��y���V�P��Q)�����
�Ѿ�[��( �-D��w+ͽ�S��@���4��n>�i[?��8? �]?K$?bxԽ��{=8���(齜�>��伤]�>�?��M?�F?���=ap�>|��Z��z�¾��5F�>�H�>=3�>Q�>A��>�t%=1I�>�$M=j�n>�>̠�=����6/�C�J>0��>�
?��>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��u�T�4:>9����j�5`>�+ �~l���)��%Q>wl?��f>Q.u>Ә3��a8��P�a|���T|>u*6?�39��u�'�H��eݾ�NM>{ξ>��C��e�������I}i��|{=v:?�?����߰���u�A��"QR>)3\>*u=�{�=IM>�Gc��ƽv�G���.=a��==�^>i=?��+>�/�=i��>7���O���>aB>X�,>@?3%?l��(���Ck����-���w>#q�>q&�>�h>��J�[�=�5�>h/a>������%�(�?�0&W>I�{��_��sw�)Ty=d���� �=�͓=�� �`=��#=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>]������'��Tv�u�=�s�>��H?����\���;�d
?�?���g����@ɿw�v��h�>rV�?}�?m�;Л��?���>p��?�'Z?��n>�Qپ�aX�q�>A%??��P?�`�>��S &�
r?�0�?ae�?��Q>V�?M�e?���>�� ���)��������p=�=p�:���w>#>�G̾`�L�R"��0��:�m�y����a>���<�h�>B}��O=���=��z�ֶ������P��>�s�>E>a>�^�>��?���>��>tw�=r3���H������W�9?4�?�tɾ�xX�Hl(>&�W��dؾ��->b%l>���>Az�J�,>; L?��?JK�?���=v6��� ��݀˿�����)����=�S?�a0?%$(��߶>�������~�>0�>��;���D=i��5�=Y�>:�F?�<�>9�ɽ=� ?�T#?��e>H��>@eE����9G����>` �>S?.=~?��?P�����3��=��R��c�\��K>��y?aO?�>7����jV���\�N拽C)�?��g?~��?���?Z|=?�@?0N_>�n���־I&����>��!? ���A�NG&�&~��u?�;?���>�T���սI�׼����h��n?R-\?i:&?j��6a��+þ���<��$�ŎV��<(�?��>�>�~��Lʹ=�>p�=m��~6�*Cg<��=~�>��=�'7�R����H?O�b�\SԾ1}2=%���bZ�<�a>��?w�i�2�X?��C>k���>��к��Ă���?�T�?B��?��<��Sl��V?�[`?� �>FC.?��z�Fb��n��pMֽ�.оSjM���>��>��Q>��߾-�����>���gи�s��R>�>�.�>}�
?)� ?j}N>���>ك��O�%����Ӱ�(�[��j���9�d*.�I�����&"%����A�¾�qy��"�>����T
�>�
?��d>;es>���>� ��ߍ>�pU>#�>�`�>l`>�;>o >V��[Eڽ�KR?����"�'���辿���g3B?�qd?Q1�>bi�<��������?���?Ss�? =v>	h��,+�n?�>�>H��Vq
?T:=�8�';�<V��x��3��&�1��>E׽� :��M�@nf�wj
?�/?�����̾�;׽�uk��<�ux?O� ?'u(�F�Y�����1I���P��슽���a��`�+�M�u��H�����.����8��>IC>?�B�?e�L�!G�Y����抿�?G�/�>�+?rA>>\�>�V>�3���<�%�l���A�=T��*��>��?�x>��J?��;?Ԫp?��z?u��>���>B�t+�>NI>@;�=Mب>�7?�a/?��A?G��>��;?>&>�*���~�䂾�$M%?_�2?���>�l-?��#?y+B���=F�����%���V;>��=�䯽֝�����KW>���>�?� ���7����Sfl>u8?���>�_�>=׍�������<d��>��
?�ď>�����Xq��S�ń�>h��?���� =�u)>Qe�=���ٻ���G�=پ����=p#��՜;�(<8��=k�=����윺ixQ;�;��<u�>$�?���>�C�>�@��9� �U���f�=�Y>oS>>Fپ�}���$��|�g�'^y>�w�?�z�?
�f=��= ��=�|��yU�����7���U��<�?GJ#?XT?T��?w�=?kj#?H�>+�lM���^�������?s!,?A��>�����ʾ��ȉ3���?S[?y<a�E���;)���¾��Խ,�>�[/�q/~����3D��酻�����0��?ٿ�?A�9�6��x�߿���[��}�C?�!�>.Y�>��>-�)�G�g�T%��1;>���>IR?�2�>hP?�z?�W[?.�U>P~8�����Й�TK�,�$>��??��?���?�	y?C�>j�>,v(��ᾋ�����!���U����+]=�-[>�J�>I-�>4��>��=�WȽP1��A!>���=�^b>��>�ť>�d�>�Mw>��<��G?E��>b����/󤾍ʃ���<���u?홐?%�+?��=�����E��P��|C�><p�?Z��?�7*?��S����=��ּ�޶���q��(�>)ܹ>�/�>�Ǔ=��F=8d>,�>���>Y��\��p8�&VM���?�F?���=3ƿ<�q�1�p�ѱ��|�b<_���E�d��r��4x[�8>�=�����Y�6�����[��������B�������{����>��=���=���=�P�<�5ɼ�J�<�J=xތ<�
=�o��]q<:8��һԊ��]����Y<�I=oC���F˾�8}?I?��*?�C?��z>��>=�1��>[҅��?�V>ÆM��𻾙�:�⧾�u��a�ؾA�־��c�������>�J���>]�3>1n�=V��<!��=�r=z��=��M�>�=3�=}V�=a�=�P�=�>y�>�6w?X�������4Q��Z罥�:?�8�>h{�=��ƾq@?��>>�2������yb��-?���?�T�?>�??ti��d�>M���㎽�q�=I����=2>r��=w�2�T��>��J>���K��A����4�?��@��??�ዿТϿ5a/>��7>k;>��R���1�6v\��b��Z��!?�H;�i-̾�+�>�
�=�.߾��ƾ'/=Ð6>��b=Q���\\��Ù=9	{�(�;=�gl=�މ>��C>�~�=:+����=�qI=���=6�O>���j�7��O,��3=8�=Ǯb>&>C��>��?~�0?4td?�j�>#�k�k�̾�Z��sь>n��=d,�>�'�=�?B>�M�>��7?i�D?��K?��>��=��>�?�>׺,�S�m�z�侻����<x��?��?쳸>үj<!�B�O ��>�Tɽ��?\D1?��?\Ȟ>6l��B�s��&<��������<m��=P�4�����B_���{�`����>��>���>��e>~�k>���=��}>�>Ge=sټw�A>N&��QFʽA�<����V��<�%>�SD=��d>xͯ=i�m�m~��3���N =�Y�����yG>Ɂ ?��S:c�>���=��ξ��=��$���,��j<��S<)�R�h��;���;�0����z�=��>IY��8��9#%?:�\>�I>^��?!�~?�(���(Ҿ�9׾�������ck���od��,�<x}$=�V���x�o(l��]����>���>�P^>)BF>�!��s6��
���r־��$���>(鶾�*[��Iw������� ���%p�{�<$WC?�댿��#>;{?�n1?��?�r�>x������>Gsf�J�Y��t�+�^�3ª�G�1?i�?kn�>m��s�<�c�E��!e��M=W����_��裿��M���>��l���:>SvU�ײ���b��Ë��d��r	r�!/ξ��>�}�?(�?���X���Ҏ=��3�����f*?5π?x�>�N
?�?ۊ���龏	q�h9�0�[?�*�?.��?H>���=Err�V�>��
?�;�?���?4z?���J�>�֖�o>Y�2��!�=P��=�T�=��A>$�?v�?~�	?�CԽvo�����W���d���=6�F=���> ��>�/�>�J>�b��sF=�/>L<�>���>�mh>S7�>�v^>KK�������?,��>� >�G?D�>��w������,��Ľ?����ܽ󷃽j�ν. ���]׽�A��b�����3?�!׿ix?1�J>���VY7?��߾O�>���>N��=s2_�p�>��X�Ko�=���>�x�>�Ӄ>h��>�q�>
���]>����"�#C�Y�X��;l}>(��T�4�����_ٽ)�w�I�þ���Wr������d=��!�=�c�?�p������7�����>���>]�@?rYf�������>�e�>1`>*���8~��'���ܾ���?���?�;c>��>I�W?�?ؒ1�33�vZ�,�u�n(A�-e�V�`��፿�����
����.�_?�x?2yA?�R�<-:z>R��?��%�[ӏ��)�>�/�'';��?<=u+�>*��/�`���Ӿ��þ�7��HF>��o?<%�?wY?@TV��t�g�J>Q6?ja_>P�;?�<I?��M?�ǽ�$?����@�)>�?�(6?��?7�>�\�>J����P=��2>r���<�d!Ͻ�=��x����9<�J=���=0���a��V=�j>�H^�T޼�Ц��P�<$���{�C=�E>;ۦ>��]?�p�>@��>-q8?���B8��0����-?��X=Y��������/��G�>X�j?��?X?h�[>�C���C���>��>�(>�Z>�`�>�F��C��0�=�>�X>���=z#M��B��+��i������<� >���>JQ|>���?�'>;[��6z���d>�R� ں���S���G��1�e�v��a�>@�K?��?A�=v龆Ζ��Ff�i&)?�X<?GSM?��?��=;�۾��9�8�J�O��>�ƪ<������w ��/�:�ȇ�:��s>�&������d4^>W��S�ӾW�m���K��X�
�-=�
�P�C=l��˺ݾ���}�=�	>?�ƾ� �1����᩿V�K?Q��=M���8�3������#>y�>ҷ�>�
�w ���<�����W2�=��>e�<>x�ٻ�S꾇�E��8�&�>�JE?�U_?%k�?�+��s�)�B�����YR��Iȼ��?�]�>@b?cB>���=���;�}�d�MG�5+�>}��>���6�G�kE������$�}s�>y<?��>D�?��R?��
?ј`?(*?dJ?d&�>��������A&?C��?��=g�Խ�T�s 9�IF�,��>-�)?��B����>K�?�?�&?�Q?��?��>� ��C@����>eY�>��W�qb��&�_>��J?��>O=Y?�ԃ?(�=>~�5�ꢾo֩��U�=
>��2?�5#?8�?���>���>.1�����=�{�>�-c?���?)	p?��=�J?v�0>�r�>�=�=�`�>���>;�?IcN?4}r?�BJ?��>X�<�*�����yKz���\�Q�;��J<&5�=tM��}�CU�?��<�K�;�̼���]v��tK�b���M,<�_�>��s>�
���0>;�ľ�O����@>ŉ��:P��Tڊ�	�:��޷=��>��?��>�X#�ӷ�=��>JI�>P���6(?��?�?v�!;�b�5�ھ%�K���>:	B?���=��l�������u���g=��m?��^?e�W��&���Q?���?�1�"=H�R������l8����>��>� F��� ?�ė?Z\^?�>ġ��������f�l��p��p�U��߷>�H�,�y��>M�(?K��>}�> �L�P�Ǿ8$����¾T ?�	�?��?N�~?�>��W�������K����_?�%�>5³�o�?7�ؼ&����m���*��y��{����b������P��Ʒ#�k5��r�����=��?Ȑq?�Rn?M�U?���z)^�~b�(W}���W��#
�����A�e,9��:�b$m��������j���_=D쑾}�W�C|�?V�/?���O��>.���6a���J����=������<�E�=���$=R����|���۫��Z-?���>��>ͩ?��6��a�)�J��=�i�g���~>�{�>}Y?���=A&Y��4�/�ύ��}��;v>=}c?@�K?�n?7P�3+1����!��X0�C>��W�B>�>���>P�W��x��8&�QY>���r�����q����	���~=�2?�;�>V��>!M�?� ?�q	�$\��rx���1��Ђ<:�>.i?K4�>|��>h�Ͻ�� ��q�>R,p?}��>�q�>y��^�"��H��d��h�>R�>W�?���>n��Z�	��{��8V=�J�=h�g?dp���d7��C�>'-I?�^���L�<W(�>���=U"��:�7�e+>x�?��=A�Y>�μ�~���.}��	���K)?�I?)ᒾâ*�BE~>�!"?�~�>n'�>6/�?1%�>&oþ�?��?�^?�@J?�OA?qA�>*�=E����3ȽS�&�Q�,=�>�Z>vm=�}�=ʻ�Gu\��}��D=rx�=;yμ�:���<<����nK<���<�3>�`ٿq^I��}���s �M��L�"�rqa�{]�:>�F���G�"}���+ȾG�����7���6�L���VLr�)����n:��[�?�p�?�����۽������b��r�+�v>�v�����A��� 8�����Z������ �0C���j��>|�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@}A?��(���쾗V=���>�	?��?>T1�xI������T�>{<�?���?ZzM=��W�m�	��e?y<��F���ݻt�=<�=�D=�����J>U�>E��TA�O?ܽ��4>�څ>}"�����^����<�]>��սC<��)ք?ux\�Jf�a�/�U���|>��T?E&�>��=Z�,?04H�Q�Ͽ3�\��a?�.�?��?y�(?ɿ�Vؚ>��ܾ��M?�E6?���>�a&���t���=t^�0ᢻ��㾄 V�1"�=*��>uu>k�,�l��M�O��똼���=� �g���F2�|����M�2�&==7@��6Q=���ߛW���������;���>ߎ>�X?>�/>L%�>�JU?%"h?��>{�L>�=�M��s���15>��~���t�-�о �m�ǾX���ݾ�(�F��U��罾g"=���=,5R�W����� ���b���F���.?"y$>A�ʾ	�M�	-<qʾ����ڄ� ��-̾ޗ1�U n�L͟?��A?������V����<O�Ε��,�W?8P�N���묾כ�=C�����=�#�>/��=���!3��S�v0?�\?����&_��8)*>�� ���=��+?�?ɉZ<'�>bM%?��*��7�3b[>̣3>�ף>���>�<	>����U۽��?7�T?���7���ܐ>�b��Y�z�a=�0>g:5�=��p�[>�s�<����U�1L��Xa�<@\d?`�>�o<���o�ƾ6Ń��,��d�?��?��>�0�?K�9?�"*=�����熿�S9�*��E�??��g?��p�w�I>s�Fv���0S?=�0?�C�.׿��â�;5�A�ۨ4?�~?�/?�l���\��������P�)y"?�؊?�G3�i�����Fs��|<E?���>Ws�>�#�̀��k�?�'�����ÿ�����j�?�R@\��?0�<'x0�o��X�
?a6�>=��V���:�<�-��dh>Ǻ�>L�����	ξ��y���>�X/?�k�>���,`���z�=�׶��L�?/��?^@��0�6=L���b�b;�D$@���+=P�h�;���\9�~ža�Xϭ��:޼-l�>��@�f��Ӂ�>��΋ݿ�οA���$о�Ʉ��(?/.�> �����M�j���|�.�I���@�*i�oM�>��>5���o���2�{�hq;�M+����>-
��	�>ݿS�'������"|5<,�>d��>��>~)���罾&ř?sd���?οު��ݝ�ּX?h�?�n�?�p?Ş9<��v�ܐ{�p���-G?��s?�Z?Si%�~<]���7�v�j?v^���U`�r�4��HE�U>�!3?,E�>/�-�F�|=`%>��>�e>3$/���ĿJٶ�������?X��?�o�+��>耝?�r+?i�N8���]��.�*��:,��<A?�2>������!�Y-=�MӒ��
?2{0?@��d-�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?;��>�9�?�!�=6%�>A�=[�����f��E!>e�=�=��?g:N?t��>pl�=I�<�!�/��F�fIR��t�&�C� D�>5�a?��K?;�a>�����:�tA"�kwн��0�$��u<�Wk)��zܽS�7>y4>>��>(G���ӾR�?[m���ؿ'j���r'�_04?ٮ�>� ?8����t����:_?es�>m:�0-��_%��A�"��?�F�?��?ص׾�ͼ�>n�>J�>�Խ�柽2�����7>4�B? $�iF����o�?�>���?ʷ@a׮?�i�^?S������陃�*t꾳�}�a�¼��h?!� �E��=�Y�>�9�<���Z���B����>]k�?���?al�>��h?zS���s�s�=���>��?�F?^*������f�>���>�;�����I��`݉?j@��@K��?刺�jֿ*⛿�����໾���=4K>=EVH>H�q�q�#����;:v =�΀�ռ>C`�>-nd>�&�>��L>S�>c`l>�҂��6�p��������MU��,�%�
�83���
�n�:��ž�9�%�����Ƚ2=�E�|G��J����!>�T?��8?�M�?�S?�5��qe>�'��cC��ĳ>z
���D�>��$?$k?2	>?�}��򄾺�R��싿�����4����?��?�ɽ>B��>?�=�<C�>=��Qiz>I��=w�����0l+�?�">��>N��>���>�C<>�>'ϴ�2��g�h��
w�{̽�?Ձ��C�J��1��^9��^����j�=_b.?~{>���?п~���v2H?����>)�W�+�o�>r�0?�cW?�>�����T��8>���j��_>+ �k~l���)��%Q>l?M�f>�Vu>�3�"f8���P�����.:|>�6?�
��w�8���u���H�.CݾiM>�Ѿ>`�D��n�����Y��Zi�GQ{=�m:?s�?�l��Uذ�w�u�[T���ZR>�\>=[b�=�3M>W�b�Ϊƽ&�G�r�.=ԡ�=�^>EW?#�+>���=2ݣ>vc��zAP����>́B>,,>�@?�)%?���kٗ�������-��w>�R�>��>�]>!YJ����=�l�>.�a>rE��ƃ���s�?��vW>~�߅_�nou�0�x=K1����=%�=� ��=���%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾTh�>kx��Z�������u��#=6��>�8H?�V��+�O�r>��v
?�?�^�㩤���ȿ1|v����>W�?���?\�m��A���@����>6��?�gY?�oi>�g۾9`Z����>̻@?�R?��>�9�R�'���?߶?Я�?�I>���?s?���>iVy��b/�QA������^{�=�5x;�>��>�=��{PF��ᓿ8}��R�j�k��+b>��!=�/�>�0�e���i�=ŋ�)g��7�l����>��p>�I>��>�� ?d7�>���>\B=�o��)���i��A)?��?�پ�ꄿ||�=��`�N#���#>���<B�>�A�+�>n�b?��?��k?�q3>��(�H��Ōտ�픾�6��E�>m(?��W?1��.�>���a�E�.?��=�Ǚ��վ��E���=�N�>Y�?�o�>o#�=�� ?��#?)�g>ė�>�BE�?���F����>z>�>N?�]?�7?��@63��U���
����[�u�M>�x?
�?�z�>�F���@��ک���F��+����?�g?!���?a[�?�??�vA?�f>'{��پ|!��>��!?���A��M&����N|?�N?\��>�O��W�ս�ּ���2{��,?�)\?�?&?F���,a�aþ�@�<�$#���U����;miC���>z�>�����=�>7Ͱ=/Mm��L6��g<�l�=}�>�=Y,7��o��1T3?�ٕ�%����@r=�u���?�Q�>��>Tڱ�u`?�½ܡr�W��Y|���O��`7�?���?��?#a��͛b�37?�݃?�p?Y��>@�ؾ��뾖���7�p��L;�QW��<>p��>?�=5&�����J�������'6���>
��>#?[w ?��O>�M�>�<��� '�zs���S�^�l��l8��.����Ӡ��*#�_P��5¾�{�HH�>jN���
�>g�
?8h>˕{>)�>�`ɻEN�>�-R>�>ps�>�X>�5>��>�J<`�н�KR?�����'���첰�43B?�qd?+1�>�i�,��������?���?Ns�?j=v>h��,+�+n?�=�>l��[q
?nV:=�B�C�<�U������3����z��>qH׽� :�QM�unf��j
?�/?�����̾�=׽Ԥn�3�����?�Z?�4�I&?�.{����6�=0V�z�?��>Ծӣr��%��g`�lƔ�v������3�1�< >�H2?D�?�>������0�-L��znN��s�>uV�>�̑>S�>�U>�<;�8�^�C�o�|�/�'-�i?�-�?*?�>+}H?ئ;?�rW?��Q?��>�x�>aĺ��X�>p�'=黊>^��>�{9?��1?[�0?�T?r�%?��P>w���O���vվS�?��?�?��?>T?����GX����k*�ٝ���م����=re�<1`˽���>W=�l>�U?���8�C����
k>�7?%�>.��>{
��_6���-�<��>��
?,H�>����yr�!b�!V�>&��?��-�=��)>7��=������Һ�G�=����̐=.���,|;�n~<1��=�
�=tXs���u����::!�;x��<r�?�r? w=�b3>&����J��H�پI>1(�>�vG>�B�>�	��&&���W���n���>��?�U�?��=J�=���=H|������Y�L*%�ܸ��B$&?��?0��?j�?7�7?/LW?Ǉ�>V?.�he���`��
���?q!,?5��>���ͳʾ��щ3�ǝ?[[?�<a�ڸ��;)�Ő¾\�Խ��>�[/�[/~����BD��������k��(��?쿝?kA�R�6��x�ؿ���[����C?�!�>
Y�>}�>N�)�r�g�_%��1;>��>cR?��>�P?��z?G:[?E]U>�8�7��Dޙ��>O��@$>t�??晁?�܎?(y?y��>�Z>�f*�f��������_�������^=rV\>X^�>U�>���>���="]Žhg����>�֢=��b>�w�>��>=�>[Ew>� �<�J?��>�aȾ^�Jl��#�`���"�M�q?�@�?��#?=m���K�� ��>��?�٭?��/?�LO�7��=��Ѽ@j��8�h�Bֺ>s/�>��>/r�=҈�=j�#>�n�>���>���gN�K<���e��-?��G?��=��ÿ�oj��L��{���˼FO��Ro�߿��F1�"4�=Wܗ��=�M����P��ᔾWʜ�l��:���	텾��?�6n=>΄>��
�$'�;��"��<�b"=�B�=��p��0=�J��c�u;�sx�:��<�r�<
�=	鲼�s˾j_}?�7I?�+?�C?b�y>��>�4�"�>�a���9?oV>�N�Q4���;�����$��Ăؾ�8׾j�c�V����j>�I���>?3>l�=�h�<zZ�=�q=�׎=@�Q�#=�"�=Xݹ=�x�=)��=�3>>��?%}_��9��z	O�%%	�[�P?iD{>T�+>��̾��?��=\!����¿+C �J�w?���?t�?s
1?���y��>ɤ��r��]�=�v�aF�>� ;>�E���[�>�kg=�	�!�������~�?��@�L:?W@�Sm���y@>��7>P(>q�R���1�1�\�Әb��|Z�.�!?�J;�
H̾�4�>���=_,߾�ƾĢ.=\�6>�ib=�h�W\�|�=7�z���;=�l=[ۉ>?�C>)y�=�7����=ĺI=���=��O>[���@�7��1,��3=���=��b>�&>/��>c�?�a0?�Xd?�6�>n�dϾ�?��5I�>x�=�E�>D�=�rB>J��>U�7?u�D?��K? ��>F��=]	�>k�>S�,��m�dm�O̧�D��<���?�Ά?:Ҹ>�Q<Z�A�۠��g>�f/Ž�v?&S1?�k?��>�I��q޿_����+�ҽ�����o=�����T��nD��L'=�ʼ�t�=e��>l��>��>�>��A>��L>��>�'%>�Z�]0�=l �&;��k=�=��H>�D�>`�=ڰh�Pa,�R#��>�a��8��[�N���i��v�<���=g��=`��>�:>s��>1��=K���A/>η��a�L�P��=tF���+B�34d�RI~��/��X6���B>K:X>z��;4��V�?��Y>)l?>���?@Au?��>�$�e�վ�Q�� Fe�NSS�N͸=�>��<��z;�[`���M�F|ҾA�>ly�>)
�>yi>dD+���?��EK=Obܾ��1�"�>����9u޼���xp��G��誠���i�E����'E?�4�����=��{?�@G?�)�?%��>�N���8㾟�->����?�<�!��Ii�J ��?$?��%?Z\�>��N�C��,��M����o�>����H�͢��piY��4>s{־��(>�;�N����7��ב����]�J� -���V�>��`?Ľ�?7<i��S����Z���̾����q�?��x?�e�>���>�W+?�ӽ��5�7����X-=,��?Ҍ�?���?���<uQ�=����S�>i�	?䊗?�8�?��w?�P@�;r�>�l�<��	>�ԁ��c�=�p>��=���=T�	?I�?��?�⛽ؔ	�O?����c�=g��=���>馕>��q>�~	>��=���=�3>�>A�>�M>£�>�>�;Ǿ� ���4?��>����?" �=��=��/>`�>D�$���Z���,��K��h��s�=�W��6������
?��ǿ�i�?��">� �R�)?A���2�=Z�=�7g>ŧ
���?��$>��&=a>K>v��>_bE>�$`>b[�>+DӾ�u>?��c!�E-C�сR���Ѿ�{z>�����&�����q��^;I��n�� i��j�i.���<=���<�G�?Œ����k���)�����̏?)U�>�6?�،������>���>���>�N�����Jȍ��e�D�?���?�;c>��>I�W?�?ڒ1�33�vZ�,�u�n(A�-e�V�`��፿�����
����.�_?�x?2yA?�R�<.:z>R��?��%�[ӏ��)�>�/�'';��?<=u+�>*��/�`���Ӿ��þ�7��HF>��o?<%�?wY?@TV��j����=�=?lR?�H{?X#?ǌi?%���� &?_FX=��>[q�>��.?_$?b��>�|�=�L���=K�>/�f���l���������2�t��<~�Ƚ<"z=)�½��8����=Q[��Mr=�D������[=�$!=�@�=[$>-��>�]?�K�>L��>1�7?���Pw8�pǮ�i*/?{�9=z���{���ɢ����>(�j?" �?�cZ?�]d>�A��
C��>�Z�>�r&>�\>�e�>�x�ٓE�$�=DM>�Z>�ǥ=PeM�'Ё���	����F��<'>���>#2|>	����'>�{��d1z�a�d>��Q��ͺ���S���G�z�1�|�v�SZ�>W�K?k�?x��=�_龉2��If��/)?�]<?6OM?�?��=��۾��9�{�J� =�d�>�Y�<��������#����:�+��:��s>�1��|�����_>��	���ھ��n�wG�DJ�Ǵ0=+�=2a=:�
���Ծ��y����=�o>O3¾�"�@閿TR����J?&GO=Z���bR�����>3��>켫>�
J��j��.?��ݪ�ޏ=N��>LR8>��k����H�����>"F?h�]?���?ր��O�s��D�6����ٟ������?da�>�?�9:>c�=�촾Ws���d�F��Z�>r@�>���p�G��	���c�"D"��u�>��?+�)>�?��R?BX?��b?��)?�Y?^R�>Q2��Z����A&?S��?��=4�Խ��T�S 9��F�T��>I�)?��B�칗>��?�?��&?��Q?N�?�>]� �D@�@��>MY�>��W�Rb��}�_>A�J?���>�<Y?aԃ?��=>\�5�k颾�ө�W�=�>b�2?�5#?�?���>���>����΋=`��>�c?�N�?�xp?Q��=T{?u�2>G��>}ܚ=�j�>���>�9?؏N?1�s?��J?�O�>��<�@��_2��̣z��<4��<U�4<�Q}=�.	��{��s����<�&�;Y���ZDl����*J��f��̩1<g_�>��s>�	��H�0>"�ľ}P����@>ˏ��]O��/ي�*�:���=���>��?���>�Y#�ŷ�=���>H�>#��x6(?��?!?Ao!;��b���ھZ�K���>�B?���=��l�{���9�u���g=��m?��^?(�W�^%��>�R?Tu?�E�� �8���c�����2�J?85�>:�e=~?�*�?k?�>�}a���n�e����u��~~�w�=�5�>���ş|�)w>�8?	�?JA�=�ϛ���ƾ~5���<���)?ds�?e;�?J{?��p=%%^�i�����u���YW?��>N��s�?g��}�۾���k�|��cо����D������䱾�<R�fܖ�cq��,�=��"?��g?�zn?��^?1��n�C��j�9�{��>I��������;��>�x�<�Ym���k
��Sԡ��G�M5��]D��گ?D0+?�Yg��) ?����]��:�Ѿ]�R>�4���n���=*aN��){�?��ku���c�֊��[L+?S�>��>�Q3?��F�!K'��j?�?�/����/>���>�q�>���>�Y{�F�J�k�Ƚ�!Ⱦ�[�����Jv>�c?�zK?	�n?wV�� 1�l����!���2�zۧ�D�B>��>s�>0W��q��C&�]>�D�r�e�s��?�	��l~=m�2?�5�>���>*N�?��?�|	��j��=�x�$m1�nń<{�>g�h?�<�>��>��Ͻ�� �c,�>9 o?���>�+�>U�P���)�v
��!�F=���>�%�>u�>��>p�t��݂��H�������H5�
�=��k?�/���R���8�>"�3?��:�#���=1����*��H��������=`�?v�!>��5>�� ���!��>��i�ؾ�P)?�I?w뒾��*�T,~>�%"?�>R$�>�0�?�'�>�rþ�T���?P�^?�DJ?�VA?�I�>,�=���[;Ƚ��&�6�,=���>b�Z> m=ߍ�=���om\�;u���D=�|�=��μ9N����<����EK<���<��3>��׿�I��?о��������|T���ý����������7����`���L#Z���l��o�
����ZI�=�?Ek�?�E��\�`��͖�|	l��g��=�>�Rc���Ԓ�(�?���k�߾�����"��zP�w�d���l�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�{A?��(���쾏�U=���>�	?i�?>W1��N������Q�>W<�?���?��M=�W�y�	��{e?3�<��F���ݻ��=�/�=]k=���J>XV�>���dKA��6ܽ4�4>�؅>["�{���~^�b�<�]>c�ս�<�����?#Z�)�r��HI�b���{��>7??��;?o>i�>�#W��ۿ�xu��Ya?L��?���?3�#?=݇�J�>�����$9?\?��i>�����^���\>M�=�=,�ھ�8>���>�n�>�=鈱�?���.���>�pC=Ȁ�����Wa�j���	3������Ƙ��훽�]轃l���濾X�P��F�����=T@>% >p�N>��2>3ҝ>@�\?ßl?���>��j>��H�]H���ž�~��E�T��������S�|Љ��Qھ>����;�G���6��o	׾� =�K�=�6R�E���6� ��b��F���.?t$>t�ʾ��M���-<oʾ�����؄��⥽�.̾3�1��!n�0͟?Y�A?����W�V�.��&W�e�����W?ER�j���ꬾ8��=����z�=�$�>_��=��⾏ 3��~S��u0?Xb?����L���9*>q�O�=��+?/�?�[<�>�J%?@+�]4彨[>DS3>ž�>���>3u	>�'����ڽ�?�}T?���b��r��>�`����z��a=\;>b,5��ܭ[>搒<w����[�3	��K�<A-W?���>*�;��|����"���7=��x?��?Lӟ>X�j?�B?L+�<����T�< ��w=#�W?ywi? >�5z���ξ2���6?�e?W\K>�dh��꾨..�"b� ?��n?M?�s����}��P���f���5?�v?Ei^�&u�������V��2�>iM�>���>��9�D�>��>?q%#��J��4��� W4�(?��@���?vg;<������=M+?�`�>��O��0ƾ͑���s����q=�$�>É��O^v����pM,���8?��?��>�����ڰ�=�.���^�?9�?�����]n<u�"#l�����u�<`��=���7"����@8���ƾ9�
��Μ�����j��>cL@�(轥��>Y18�D9��LϿ�󅿺Nоֳq�z�?���>��ɽ�ң�X�j��?u�I�G��H��K��N�>�>`�������G�{��q;��'���>X�U	�>��S��&��O����{5<W�>��>˸�>�'���罾/ř?hc��@οI��������X?)h�?�n�?q?�9<q�v�!�{�=��b.G?��s?�Z?�l%��=]���7���j?����Y`��d4��E�fT>��2?���>�]-�n0|=3b>���>K�>io/���Ŀ̶�������?���?���'"�>E|�?J[+?!��'����*�
$ں�EA?�1>�\����!�=�_���;G
?i
0?
���E��h?��]�� ~�qC7��N����>POS�!Ӷ�v�<��v�-�b��Y��M���8ҧ?bb@��?��Ľ�z�ߟ%?m^�>2J���n��p�C�v��> ��>�9�>v�5�I�d>�����'�9@�=:r�?-�?#�	?�'��xF�����=��?B��>�c�?(��=��>��=�����r;2>J���ZYg<��>mR?��>H�=�+�{o.��E���X��R�J3;��cu>MM?L�G?�>d:ҽw�ѻ�!��̽��'�<68�`�1���T����C->_	1>�'=>�$��uվ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji���?�5ؾ�솿��{�>�-o���=�8Z?1f�ԡ�<3? ?�]=����w跿kx�nɽ>��?5C�?;��>F"n?W�C�.~�����9ȳ>0~{?��?��Ҽ�G��2�=o(�>N98�����/��#�?m0@�@4�[?��S�ѿ�f������Ͼ-�>.�=�pa>���c	;>����|�h<�����I>K�>�>��`>���=o��=��=�H���C�H˙��͊��2�C��5��3����������E�оx2ɾ\IO�����5q�.�t�dRD���ֽo>\qj?e�"?nB?nS?���$�>��UL�砂>��T�.U�> QJ?<zN?�K?�?K���t��J��:�����
���m�>҂?'�>��_>�;�>2�<:�?3�=�fs>?]���0�א��=;{'J>�>�>���> w�>�C<>ߓ>�δ��1��O�h��
w�!̽� �?=�����J��1���8��ҥ���i�=b.?�z>���?п����A2H?�����)�l�+�=�>,�0?�cW?ߛ>D����T�y8>Կ���j�:`>�+ �I~l�$�)��%Q>�k?��f>ȗu>Z�3��m8���P�8���g|>\6?�R���8���u�ÁH�bݾ-kM>K��>�G�o������+�Epi�O5{=JW:?5�?5���䰾�`u�/Y��9AR>5)\>o
=�o�=WJM>��b�?�ƽH�%�/=;��=�u^>�P?�,>A�=��>A6��ynP�⩩>�uB>[;,>w@?�(%?���S��l���-���v>�W�>`�>�'>VJ����=Vr�>��a>{���u��ű�D�?�^�W>�~��A_�yu�A{x=�K��o��=�I�=�h ���<�ަ&=�~?���(䈿��e���lD?S+?U �=!�F<��"�E ���H��F�?r�@m�?��	�ߢV�@�?�@�?��L��=}�>	׫>�ξ�L��?��Ž5Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?�j\>%�?�_?V�>��m�0�6�)8��X�w�A�Y=c�=ϣ>��>�ȾQ�T��͓����6i�O3���N>���<^ֻ> �rپ�������&��;<]�W�>re�>��>﹛>p�?�C�>�4�>z� =Z3��~����Ȯ�py=?��?'���Au�{����=+@/��>�L�>��=�����y�>(�a?��q?�B?��A>���n����ɿT���2Dl;�޽=<��>k�?5�ɽ��>��c���]>��h>6��:DA���sC�s�h�)Ñ>�c+?�c�>V#��8?_/0?n V>���>;|?�B���[�Y����>A��>��?P��?X�?�ǰ��q2�{)���(����Y�+�=	�b?�?�"�>Pq��"���?�r��Ɉ<[Bn?#Hd?8��<x�+?v��?>e?�E_?]i�>?S��]iҾs$��/b>c�!?	:�/�A��b&�����?�1?:�>�S��h~ֽ:�ټ�������
?3W\?n&?��Wa���¾(�<�p'���J���;�hC���>N>�������=�7>˕�=��l�k6���j<R,�= a�>J��=W�6�Aƍ�o>?D��<u�޾J�K=nf���4�M\7>J��>�lҽ(!?�7���Y��)��ֱ���봾��?���?n��?��=�d_��7]?�~?�t.?LC,?������jO������;;q��@~�>}N?�d��j�u��������낿��d=���
�>D��>N?�y ?D�O>E�>�1���%'��n񾊳��^��l�Vs8���.�_��pנ��(#��-��=¾��{�N�>�{��n	�>�
?��g>��{>A�>��Ȼ�`�>NR>�>�}�>ZX>�	5>>�>X4<)�н�KR?����!�'��������d3B?�qd?O1�>�i�8��������?���?Ss�?=v>
h��,+�{n?�>�>H��Uq
?\T:=�8��;�<V��l��)3��?�-��>E׽� :��M�@nf�uj
?�/?�����̾�;׽��������?"(,?�*�b~.����[���V�7�L<]:����M�5�\�α��7���
���S(�Y�=�{-?_�?m�����מּ���y�B�ϗ�>mD�>0Z�=���>��k>#�W�J�7e`���JW�q?�d}?���>-.G?$�=?�Z?<�O?�k>���>�B��7Z�>��l=<e�>���>;?q&+?9$?R�?Ê+?.�j>����l��c`ھx�?28?k�?�?���>�ya�5Ɠ������!<��q��ڍ��9;=���<�æ���-���=!�u>�X?�����8�����xk>�7?��>���>���S,��s�<��>@�
?QG�>  �~r��b��U�>"��?����=;�)>y��=�~���Ӻ�Z�=����[�=70���z;�Pc<���=���=�4t�����\��:̱�;To�<@;?�:?��>2%�>dʉ�����)N��к=�b>�(H>V,>�Lھ���Uj����g�XX>h��?V!�?cu=�H�=�2><b��u������lþ��<�?�A"?�[U?���?��@?�u%?B��=���Y'�� 5��T�����?x!,?R��>���p�ʾ��܉3���?�[?e<a����;)���¾��Խ�>�[/�g/~����D��օ�����}��!��?Ͽ�?A�I�6�Xy�ƿ��\����C?�!�>Y�>��>�)�J�g��%�0;>1��>R?��>#P?��z?�[?�U>��8��˭�w����e�G�#>˲??���?��?��x?�8�>��>��)�͋�B���u���d������]�_=�\>��>��>T�>Ů�=��Ž@а��?��=�tb>�r�>/��>h��>��w>��<�T?b��>���j��d>ھ��ڽ�":�gC?��?c�>iݔ���/�x�b�C����>��?�l�?�A?9�����=Ą�=�ʺ�����x��>.4)>�>q�>΄�=��>1k�>�A?���LE=��Ph��fQ�fo#?<oQ?.L�=������}�fW�9�����r�V���pZ�R���F)��[��=�)��?{����y�%�"�32���k�X���/N�����@�?&�=d�<>�H>?Q�oI���.�=��<Y��~<>��]�k7T��ߨ�G�[=?�ս�Ƚ1W:=$��=iQ=�)Ǿ�#|?�bI?�p/?�D?g>j�1>��/����>�A���?ӭ]>����r���,<�����ʋ���Ѿ!�׾��a�������>�9�9�>͵;>7��=h�<.s�=?dp="c�=�J��ޚ=/��=8A�=JZ�=cD�=Ɵ>e?>�9�?{ Y�����R�S��d�x*=?(��="�=Pݖ�O�>��μ\}�����p�����?���??��?!?�Ӓ� �>��s��
Η<{�L�z�>�g=�����'?�L{>�G�0~��~[�����?�k@J�c?s��ͤؿX�>e8>x	>��Q�G�1���[���c��wX��� ?��<���ɾ���>�~�=Iܾ��ľ��,=�3>(Y=P��7�]��?�=�~���2=��w=E^�>��A>��=�����o�=-�K=^��=qlO>����2��[+�c�.=��=�|c>2>%>N��>�?�a0?�Yd?�7�>�n�PϾ�?��rK�>�%�=�D�>��=�wB>���>��7?$�D?��K?ۄ�>ٰ�=��>�>��,�d�m��n�#̧��̬<���?�Ά?dθ>UqR<��A���g>��3Ž�w?�S1?�k?��>���Q�Ͽ��v8���>�Ft<����f���q�=V���2�_�� ��=�ܖ>�*�>B��>�@M�y��;U��>�F�>�J�=<})��qF=�3���!c��G=�<>��S�\>\�޽�k>�0�E��y�; ��<�fü������>�e�=���>�A>'�>��=���t;%>9V��2�I�
л=婾*l?�A�c�׺���0�0�;�ˏ>>�p[>�K�����y?ܫ`>��>>��?+,r?-q>�����ھi꛿Hg�t�O����=�I>G�:��>�5�b�`P�9�վh2�>Gz�>ܡ>>�l>��+�o0?��jn=&hྏ�4�D��>/��5$�]��q�,9��g埿k�h�E�����D?,=���e�=�$~?�OI?ď?=��>����zؾ�r->K��-=��~�o�������?G�%?��>:X�	E��o��\ �	n�> �8���T��͚��mH��J�=�ξ%%a>���©���1��]������F*?�������>��J?�h�?��=����3t��C��n_��Y?�P�?��>�)H>�3?��ƽ��0��gԾ��=f�u?5�?j��?��=zN�=T賽�o�>ǝ	?�ۖ?zԑ?N�s?��>���>Ɇ;ē >Bڕ�e�=/~>+p�=~��=��?2q
?��
?�����	���e���$^�I�='��=�ڒ>���>�q>ߢ�=B�d=��=�Z> ��>|�>�c>-��>}H�>kԛ���WQ+?�pG>�#>�A?i@>'���%� �확=��˼,@�P���Ùd�z�3��%�܎�M���u�ǽ�&?)ȿ�ژ?C�7>d�Ҿ�k?���~xb�E�>�o>$g���u�>ǘ�=�jf>_�>ê>7	�=�_5>���=�FӾ�{>1��Jd!��,C�ނR���Ѿ|z>;����&����v��LAI��m��Ng�:j�2.��G<=�8ؽ<H�?����Y�k���)�������?�Z�>`6?ڌ����T�>���>Ǎ>�J��^���Eȍ��gᾔ�?���?�<c>c�>��W?��?œ1��3��uZ�M�u�(A�Ie�w�`��፿$���՗
����`�_?/�x?GyA?�U�<�9z>L��?��%��ҏ��)�>/��&;�*G<=�+�>4*��I�`���Ӿ��þn9��FF>�o?P%�?�Y?�TV�0X�ڇ>��v?�S�?�?ѓ(?�&�?>����2%?E�>�?;m?��N?�&?���>J_�=5��>�&>�d�=[�߽�������<@�C"�=��>g&�<��<�pн��'��帼*�|���d=wYq<��6<M�=�b=�7b=�S�>5��>��]?�M�>���>i�7? ��0u8��Į��*/?R�9=������TƢ���v�>�j? �? dZ?�^d>�A��C��>Y�>�v&>N\>Yc�>�tｿ�E���=qL>�W>Eå=�gM�d΁�S�	�;���k��<�*>��>'/|>���[�'>p}���-z�J�d>��Q��ʺ�]�S��G�-�1��v�MX�>��K?�?[��=]龴'���Hf�i0)? ]<?�NM?I�?Z�=��۾��9�,�J�.>��>|�<z�����$����:��Y�:B�s>�2�������9c>�|�w�޾�dn�/�I��羔VF=e����]=H�H�Ծ��~���=S>i���P!��"���Ȫ���I?O�i=Q��*mT���{>6�>젮>�<�|�{�6c@�������=G-�>x�:>4!���R��IG����RI�>{\E?LJ_?�R�?Y���r�ȱB��������`jü��?qǫ>�\?�B>�H�=����'�ae��$G�\��>�g�>c��ӵG������=����$����>l)? >2�?��R?� ?}�`?��)?5A?�E�>k������A&?;��?E�=��Խ��T�c 9�F����>��)?�B����>��?Ž?��&?7�Q?��?��>$� ��C@����>!Y�>��W�`b����_>Q�J?���>T=Y?�ԃ?b�=>=�5�ꢾnө�&X�=�>u�2?6#?H�?|��>��>�����Á=��>2
c?�5�?��o?vc�=� ?2>���>�$�=7��>���>�? XO?u�s?��J?+z�>o�<�\��}����]s��O��C�;�G<�z=����Nt�BZ�}W�<��;L���#������D�q���G:�;�_�>�s>`
����0>.�ľ�O����@>J����P���ي��:���=�>��?v��>�X#�Ƕ�=���>I�>O���6(?��?�?c�!;�b���ھ/�K���>	B?`��=��l�}���C�u�P�g=��m?��^?c�W��&���[?{�j?@{ƾ�^�����;��8N�և�>�A�>I�_>��>y�?v�E?���>$8��l��ߥ��t�@��*��t�>�����q@�d�+>%k?�t?��k�º���5��BW��>X}�>>��?���?Tڐ?բB>����(��-����h����^?LJ�>����J�#?U��|FϾ�]���;��:�ྈ���ժ������񥾰�#������׽�8�=��?s%s?��p?��^?�� ��d�w:^�G��m�V�Ē��^�ёE�?GD�|HC�)�n�-X����Z��LG=�f��'U��q�?l3?VY�o�?����I׾�Α�S/	>�jv�|��tk>F<4���v=΍�=+�|��r5�r���5?���>=&�>u`?:�_���N���2���/������A>�>O�j>��>u�3�b�U�6��X�ľ��`½�v>Ŭc?CRK?�m?.M�t�0�%���L8"�%�C��ץ�k5A>[>�t�>F�V��n�:�%�r>��`s� N�-�����	�2�=��2?�݁>�T�>\
�?��?M	�宰���x��l1�wŢ<	p�>q<h?p1�>nÇ>�tͽ�L!�U��>�}s?�t�>�7>r".���^��ð�(��>�m.>�	�>GIP=20����e�q���R핿K�G�!?�=~%�?8ヾ��&��ۣ>�o?k��<��=<��>{�8�3�*��u�K+�	�X>u~?�^�=	�>Fо*�!�\��FF�dO)?5L?�䒾��*�8~>�#"?���>�(�>0�?�,�>�pþ.�>���?'�^?�CJ?(TA?�H�>�=	���>Ƚf�&���,=��>z�Z>�"m=���=���@r\��{���D=%r�=�|μH����<�r��7K<Q��<��3>�fۿ�>K��xپ������<#
�.������Zc��$	����;1��i�w��9�f<'�8^V��Hc�����+�l��|�?T.�?�-��_���s����z��ͱ�����>jwq�U7�)ȫ�;��f㕾Pྍ���9O!���O�W-i��e�S�'?�����ǿ찡��:ܾ)! ?�A ?8�y?��:�"���8�ͭ >EB�<�-����뾯����ο2�����^?���>��/��5��>ϥ�>�X>�Hq>����螾�3�<��?/�-?��>��r�(�ɿ`���f��<���?-�@�|A?z�(����V=��>ې	?��?>�U1�8J������S�>�<�?���?4~M=��W�j�	��e?]<,�F���ݻ�=;<�=L=�����J>�T�>��=SA�Bܽ��4>�م>s"�����^���<��]>��ս�<��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�F �D\ÿ�C!�)��[�=5�V�{�j;Q�	��콥Hս�¾�|����Q��]�=�BT=�:>� �>�wK>�>q�O?�r^?db�>��/>n��-S�"�ƾ�[O�2����\u����I��⏾���(e��"�Jz��������F!=���=�6R�S����� ��b���F�y�.?v$>��ʾ��M�+�-<pʾ׿��!ބ��᥽s-̾��1�"n�K͟?��A?������V����SV�5���,�W?�P����M鬾��=[���-�=%�>���=I�⾮ 3�v~S�
u0?a?U����Z��s.*>� ���=��+?ԅ?��X<��>8G%?�+��u�sX[>�3>�ǣ>���>$G	>r���W۽�?�T?���"��� ؐ>�Y����z���`=5>�I5���i�[>�U�<@���'LW�[l��Β�<�xX?�ė>��(�h�����ӨG��!�:�y?�j?�>�f?.0?�9;(v��9�S��[�^L�<�R?Q�r?��>\ˈ��{Ⱦy�þ�D.?a?y�S>"w������,���%�?V�o?�z?������z�����8�w�7?��~?��3�����P�z���h	>#?��?��Ծ
W�>�ts?Q�n�O����۽���A�]��?�@�@_=kI��j�=[��>�K�>�:����4���νo�۾���=~$�>�R���\�$e������+?��r?vq?d�������=̲����?�y�?��оI��=X��<�Y�z��TB�<I�*>HGּV�n=�ϾK�&����e�
�@~�������>7+@< q��܍>G�}�����JͿ9����b�����t ?��>��#���׾�g�$Iu�2�B��u6��pV��N�>C�>��������D�{�Qq;��P����>����>��S��'�������V5<�>��>,��>�)���佾�ę?�c��c?οK������}�X?
h�?�n�?�p?c�9<��v�B�{��d��.G?��s?BZ?�r%��=]��7�+�j?S^��7U`�@�4��GE��U>�!3?�B�>�-�÷|=E>P��>rf>�#/�7�Ŀ�ٶ�?������?��?�o����>N��?ur+?vi��7���Z��]�*���.��=A?�2>&�����!��/=��ϒ�μ
?�}0?�~�m.�]�_?+�a�N�p���-���ƽ�ۡ> �0� f\�(N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>dH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?�R�>�'�?���=���>	��=N{���%��>D��=�U*��?h�N?���>�)�=��3� �.���F���R��u���C��d�>u�a?�jL?��b>�׼���*��� �_]Ͻ�,4�����@�� ���ؽ��4>#�>>�>D�Y�Ծ(�!?q���׿,
����N��?�|>��?M���(�~�`>�<_�]?�=g>=�������#��_�����?U��?��?��۾>�\�;�>Rv�>U؁>�����^�f#����C>��C?`~$�춋���q�3z>���?��@�ѯ?��i��%?V�վ�Z���y��/���Ծ$�A>��o?U���҄q>R�(?6"�=淄�᰿��ۑ�>Bը?�_�?�K
?=U?Ac���4����=D7>0�k?�$?5Gѽ5�ž�j�>��?�W ��!���sھr}Z?M�@�@b�?,|����ѿwҙ���Ⱦ�B��HW>�1�=Io@>�U�R�=+D|��k���3��"�x>�9�>WgC>Т�>��@>�">e�=���G8��ʡ�����3@�{2�_#��ʄ2�T49��{�_����aה��٠�a����Žq���B�!d�U�2>�K?כG?�-`?�g$?\� ����>��"�/�o��l=��޽α�>̇N?��c?4^T?ŃT>�[?��#c��݌�&S��/ѓ��Q�>�R�>|�?�n�>yK�>{	�=I��>f[���w`>
�6����=
O�>r���6ڇ>i�>���>S��>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?�f>�Yu>�3��i8���P��t��|>�6?�!����8�C�u� �H�zRݾ$FM>y��>u�D��o����8��~i�l�z=>p:?,�?�����l�u��1��|8R>��[>�
=�
�=d�M>��a��&ǽ��G�AT/=W��=,a^>>X?��+>���=�ԣ>Pe���?P�W��>�lB>�,>@?'%?�&�9嗽����	�-��w>�L�>��>�M>�[J���=�k�>X�a>���؃�v����?��oW>�C~�1�_�ڀu�y=�����=x,�=�~ ���<�?�%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ|��>���Y��C����u�I�=�1�>P~H?���tfQ�(=��~
?��?V�򾦯���ȿ�lv����>��?�?/�m�L��.&@�o�>tq�?=�Y?'�j>5O۾�hZ����>�~@?Z�Q?�p�>�M��Q&�!?�׶?���?=�S>ґ?f�h?�8�>�X,��Q+�����)����g=t1M���x>�T�=&�˾��J�b����1���ci���� u>��J=��>�wƽu���N�=�v�񍜾7%���d�>�q>4�o>��>*?�O�>y�>��5<�ϯ�:@��Yx��kF?�?<����p���<�ʑ=%��Mõ>��>�t>�Ͼ���>��J?t\p?~r?V��>�[��
���{���궾�N��7N>+M�>O��>����g>�GǾXU�:>�~>�`7��a�������>��'?��>ʎ��w'?�0*?��=�Tw>�9������hk���>�,�>���>�Kq?l��>FFݾ�:������S����`�+H>��?6&?���>�V���奔`��l_-�J$�=.\�?enh?�����?�FY?}�
?��?��#<�a��R��7�<^��>��!?���A�Ud&�F��f?:Y?�	�>�E��ZXҽ�Hؼ-M��b����?Rh\?%&?����Wa�SAþ%[�<�E&�G%J���<��>���>">����b��=I�>c�=OQm�:95���v<�G�=>��>^�=p�6�J5��)~9?�
�=۾�炼�+n�Wz7�Xl5><.�>�$��E?:��k�[��ⷿ՞��4��֤�?�L�?��?��u���b��:N?��z?fy�>Jn??�҃�.l8��a�U�������\���>E�>��i��Ɯ�n���\㻿-䖿u�"<x���??�W�>�?< ?b\E>�ȏ>����D�"�^��|���`�����k<�IO.����Fv��s��ڻA���E����>�B�����>�h?'r>yh�>g��>�M<U�>jP4>���>N�>@bH>��>���=����ǔ��KR?����!�'���辻���a3B?�qd?M1�>i�5��������?���?Ns�?=v>h��,+�yn?�>�>H��Sq
?�T:=�:�;�<V��d��e3����F��>E׽� :��M�1nf�}j
?�/?P��ŋ̾�;׽Q�z��= �?i="?��5��3R�#炿J�U���U��w=�ђ��Y�v���bg��������Iσ�ʩ!��u=��-?�˙?�L@��A�Y5�����A��3�>V�?���>�O�>�;�>Q26���S���g�%�?�ؐ�}�>aA�?���>��H?(Z=?�hU?��O?��>�[�>u3��s�>��)<��>���>]�:?3?T#4?�?�O)?_�D>���6���pԾ'�?<�?��?��?�?&�X3���J�R=F��9w��1���g�=��<e6���D��2V=��[>Y?!w���8�����
k>�z7?�`�>|��>I��=���T�<���>#�
?�2�>� ��r�e�U�>�?���d=��)>n��=ﲅ� �κ[b�=я��Tސ=0����;�o�<��='�=�t�]�<��:�C�;t�<1{ ?!"?|�>��>�}�Ff��v�o��=��U>9 )>H�>�*⾾7���͗�K7f��ZX>���?���?�'�=�@>t��=}ٜ��ľڬ�ꐹ�1�9=Lt?��"?=iT?ȇ�?|�4?_n$?��/>ک���]��t����?� ,?���>���T�ʾ�憎�3�M�?�T?1@a�^��;)���¾��Խ9�>@T/��,~����D�ʰ��*�������?%��?��@�l�6�v�ͽ���Z����C?,�>FT�>� �>�)���g�R"��:;>��>�R?�m�>��Q?O�w?b�O?��Q>h�4�N/���������;�J>wT7?�g�?$/�?Hct?�M�>O>c;:�T��^J���A����ֺw�-�=�-o>��>G��>f©>��=g�����VK����=o��>� �>䍦>~]�>���>�xһ3H?�~�>	����U��ۦ�B����0���u?ڧ�?K�+?0#)=���6�F�����]�>{��?�P�?|�+?��R�� �=�+Ҽ�R��m�p�hb�>���>��>;ێ=��I=��>*�>K��>�����G�7���F��#?�#F?���=?�ƿ�	y�y����{���M>y�Y�I}�|�>(�D9Q�~r��+䥾?�:��޽�f���2��D��e�p�a0��g?D��=��:>�>��9�x��=��i:�D =�Wf=�� <e����$�=HT<;|�<o�����8�|�(�:��;�˾�}?�;I?�+?��C?2�y>!;>��3�[��>놂��@?QV>��P�爼�J�;�5���� ��N�ؾx׾��c�ʟ��H>�`I�$�>�83>�G�=�K�<M�=�s=�=R��=.$�=�O�=mg�=���=��>aU>�6w?T�������4Q��Z罝�:?�8�>�{�=z�ƾq@?��>>�2������~b��-?���?�T�?J�?>ti��d�>?��z㎽�q�=����=2>$��=��2�N��>��J>���K��7����4�?��@��??�ዿϢϿ5a/>
�7>�B>Q�R��1�r�\�w�b���Z���!?�J;��J̾('�>��=_.߾�ƾ��.=tn6>�a=s��O\���=�){�%�;=l=ԉ>?�C>���=B����=�wI=��=f�O>>B����6��b,��3=���=�b>�&>c��>��?�a0?�Xd?�6�>�n��Ͼ�?���H�>��=�E�>L�=�sB>r��>g�7?f�D?��K?���>h��=	�>��>&�,���m�<m�I̧�0��<���?�Ά?�Ѹ>z�Q<}�A����<g>��.Ž�v?%S1?�k?��>�Z�4ο���qy�O�=/=>�g>.���O��	z�����4���F�^>FI�>N(g>$)>�>c�(>ߖn��q�>ڷ2>'�=Hr%>�?���<ń$=м<n�<g��)����7�E���5���:x�<O��5r��R]�=���=�>Y �>���=m�>nl�=�õ��ؽ=x>��"/=�MC=L���Y�;�)j�3���O-�d�,�B�@>T�s>��������[?�5z>��_>���?�Zl?un�=nn!��&侂���J����d�+
>*?�=5�,���H��Kt�bvW�F���h��>���>-�>�e>�6+���=��	f=H��kG5�C��>�d��}�?����p��a�����9�i�K浻ֽE?������=��}?9H?���?��>x>���Mܾ\!(>�oy�!�
=o��Wo��͌��~?��'?W�>�9�jF��奾_e����>�u�<6V�ޔ��Mt1�O�><Q����>'��HI��a�5�����œ��UM�����{@�>~a?��?T�n�̩����R����j����?��v?���>���>m�?Z
潶� ������ڴ<�x}?���?���?�=8��= ��4Q�>v4	?���?	��?2{s?Qm?�W��>s~�;� >ߓ���U�=��>Ҫ�=JP�=Ol?�
?��
?A1��X�	���,��5�]�m��<S��=�}�>�h�>7�r>n�=�{g=T��=��[>}Ξ>��>��d>��>rL�>0��	�!�A�C?3��>�K�=b;k?��>d5A=w=�O�z�F��#���?��:p�=Rm����=PLս?dO�C�N�l�?r���L�?��>5c��(??� ��P�=�j�>Gw�>$�=���>MI�<3<�>�M�>��>i>6!>?vҾ@�>���<&!�l�B�	gR�%�Ҿ.{>���k '��P�j7���J��õ�)|��3j�*����<���<f8�?�����k��9*������??&��>wJ6?3��Ն�x�>�\�>ύ>�a���u��輍�8X��?��?�;c>��>B�W?�?˒1�23�
vZ�%�u�j(A�1e�U�`��፿�����
����#�_?�x?/yA?zS�<4:z>N��?��%�]ӏ��)�>�/�';�M@<=v+�>*���`���Ӿ|�þ�7��HF>��o?8%�?rY?&TV�����>#�W?HO`?g\�?�L?0�A?M�I�C�&?���=o��>��>��2?,0A?�j.?��>�,7>��	��_��\��[�|P���Ȼ�g�X=+�>�~�<鋺=�v���K�u���*���}.=�Ľ( +����9w�c=��=.�/>���>r�]?y<�>~��>��7?����8�F����#/?��8=-���g��آ�l%�6�>��j?t��?X`Z?�sd>7�A�
C�N+>�\�>�n&>�\>�^�>�Mｸ�E��͇=c>@4>���=	�L��΁��	�X�����<7>���>�9|>���'>Oz��1z��d>{�Q�պ��S��G���1��v��X�>>�K?��?Ȏ�=�c�:E��Hf�r,)?�\<?)OM?��?��=��۾��9���J��J�Z�>��<��������#��j�:�z��:��s>�2���Ǡ�2�b>����ݾ��n��J��{羓vM=�n�FIV=p�S־G��M<�=M�	>���� ����<ժ�J?��k=�G��k�U�D��x�>a��>4�>wU:���u��t@�鉬��=�=���>~�:>�t��	�vG�!2�9��>L?$L?�V�?�n�6�x��X��t������U��=�M?���>���>0	>&��K.Ӿ����Cd�=HJ�(��>�,�>Y�	��D?��aؾ�վ��)���=�~�>(�S>�}3?�s?δ?�m-?^f?ٖ�>8ύ>,}�����:&?㋃?�ׄ=�ս��T���8��F�0��>0�)?�{B�M�>?-�?R�&?piQ?G�??�>�� �<J@��~�>�S�>��W�_���I`>��J?���>4Y?{Ճ?2�=>�{5�梾�Щ���='<>��2?�)#?��?Ȱ�>��>���=��>{c?u.�?�o?~|�=|�?;n2>���>h_�=���>
z�>Z?�QO?��s?3�J?���>�:�<�O��ⶽws���M���;��G<��z=���]�s�%�����<N�;B��������ND��S��?[�;��>��}>�	о=��;�G˾L����C�=�ٙ�8�U��ڰ����eļ#��>�i?���>�a`��d�=�V�>���>�x ��# ?�2�>�!?�l3<Ͽu����䲽,uW>��?R�P>�_M�l2���⃿-��?��u?ʎԾ�>���b?�^?�]�O=�C�þh�b����K�O?��
?��G���>��~?2�q?ɕ�>�,f��@n����[9b��k����=Zm�>�M�:�d��_�>��7?\F�>��b>H��=��۾
�w��m���?��?���?�?+*>y�n��$����L��p?9[�>�թ�@�8?h�^��	#���V��qH��;՘Ӿ|gѾ�������
D�`�Y�Ɯ�l�<�)?�i�?��w?�1N?���K�MN'���Y�2�9��d�?���Hm�t�K�_�:�&*L�x�����g]����C�O��sjB�]��?"�?�9���|�>�։�E�u�O�ƾ�=>=�O>��Y %�$�J��r��<@@o������۾J�6?���>p�>��?�k�S�C��7���*�Ń�i�=ϸ>^З>a��>]�(�c|D�f��ܾ��O�N�3�v>^�c?X�J?��m?�����0��5����!��)�������F>F�>���>r�X�[�ʱ&��>��`r�qd�����#i	��	�=�Z1?�ق>�ٞ>���?H�?�>��f����w�41���<�[�>��h?R�>PT�>vʽ6 �;��>i�l?��>�Ƞ>�����X!��D{�M`ν���>Ԅ�>l��>��r>F�+�m�[�c`�������B9�B�=|�g?>����_�Ŧ�>�'Q?x�:)�o<��>��y��
!�p��O�%�n	>}V?0��=��;>��ľ����z�;����Q)?�K?r쒾�*��#~>�'"?u�>o�>�2�?z"�>�lþ��?���?��^?kCJ?�FA?75�>+�=���_WȽ��&���,=�x�>A�Z>m=��=H���l\�[��čD=�K�=Oμ^����<@���V K<JT�<�3>�hۿ�JK�9mپW���8'
��刾���bX������X������gx�����'��V��)c�V���g�l����?9�?�X��)������ƍ��S���'��>��q��������V�;��w��U����b!���O�i��e�Q�'?�����ǿﰡ��:ܾ2! ?�A ?2�y?��4�"���8�� >�C�<\,����뾫����οB�����^?���>��/��j��>ҥ�>�X>�Hq>����螾�1�<��?7�-?��>Ɏr�/�ɿc���T¤<���?/�@<xA?��(�����WV=)��>�	?C�?>�^1�qD��簾�Y�><�?���?+eM=��W�-<
��oe?�
<X�F�T=޻��===�=7=����J>gJ�>֥�0VA��
ܽ��4>_�>8"����P�^�X\�<`�]>;�ս���!Մ?8y\�f���/��T��%P>��T?S(�>�@�=9�,?�7H��|Ͽ��\��*a?�0�?զ�?e�(?Kۿ�Lۚ>d�ܾƉM?�C6?���>�c&�+�t����=� ἴ��j��(#V���=��>�w>9�,����zO�ộ�i��=^k���ǿ���ʰ�=�߻�G�=����i�<:C�����<Ilx���M��j���<<Bz,=�h>z��>ԆE>�->4�K?Kgl?��>|:>C��[Qo������~��{T��DY������3Ͼw�Ҿmy������&�'��@��!=��=7R�j���9� �Y�b�L�F���.?w$>U�ʾ��M�â-<}pʾd���:܄�᥽�-̾�1�"n�h͟?��A?������V�T��vW�U���`�W?YP�Ļ�mꬾ���=���;�=%�>슢=���� 3��~S��o0?a?y~��BS��zP*>T� �k=��+?]�?��\<r2�>�S%?E�*�;�V:[>��3>\��>ê�>�	>���'�۽P�?��T?������aِ>�Z����z��ya=R8>^5����،[>�Q�<�ꌾ�T�K;����<�&W?Ϡ�>-�)�8��_��U���V==��x?��?�/�>F}k?��B?�<1h����S�$!�%:w=_�W?y%i?Q�>舁�
оA����5?[�e?�N>�\h���龙�.�[T��"?{�n?�^?�I���s}�D��H���n6?��v?s^�ps�����p�V�T=�>�[�>���>��9��k�>�>?�#��G������sY4�&Þ?��@���?��;<��X��=�;?m\�>��O��>ƾ9{�������q=�"�>���vev�����Q,�w�8?㠃?���>%���������=�ؕ�Z[�?�?I���,Bg<����l�o�����<٫=�1��Y"�����7���ƾ�
�����*r��L��>�X@Y���>Sa8��3�BRϿ`��>dоYq���?��>FȽ�����j��Lu�V�G���H�����Q�>�>���������{��s;��؟���>�����> �S�e(������`35<��>��>TÆ>�.��w彾�Ù?�]���Aο������ �X?�d�?qi�?�p?��9<�v��{��6��2G?B�s?�Z?~%�oT]���7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�/�n?Wk"�d(��C��dO�=U_�����E �?�{����D�w��y���S��N׷?1��?8��?��h<�L�j|L?��>�XV�ҟ㾋R�<�
L>��?{��>��:�)?2�r��C%�<�=H��?^_�??=�>�����ʛ�&�M>u(�?��>��?��=[��>B��=j���`D����>��>*T����?��P?$X�>t��=��R�&�2��H��O��@���?����>��[?�>?�/p>��E����Mf��Ӟ�'3���3�gD ����
н�"8>�>>:�>�v)�>ľ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��$	?[���g����x�b4�W�=��E�=W7?�w��U>U��>�=�|t��{��bq�H��>�S�?���?��>[�n?e��[L��}{=�4�>�*^?�w?�6P�=����*>��?�b	�Y������3�n?�n@��@]?+Y����ͿR-���j��S���
�=���=�c>�W����=_ap=����=k�>�T|>�%B>�xQ>Ȉ4>�YN>�;>>U�����%�أ�������?�������r�x�������&�x�������g��LoڽaϽ�W����@�4����=�Z?e�@?��k?PC?bq��U>�t�-6$=��׽a�=���>�?��C?�2?�Z��"���nk�dx���*��������>�H�=%�>6;�>ӣ�>?'8��'>��>��>٭�>!��=����s�;fYA>���>N�>���>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��u�T�4:>9����j�5`>�+ �~l���)��%Q>wl?'�f>�v>Cj3�-�7��ZP�S����1}>��5?i���1J8�#�u�1`H�cݾDqM>��>*�V��������a�`ci��py=Hc:?� ?t쳽�x����u����F�Q>R]>*� =�ְ=�9N>��d��ǽ�G��/=�7�=t;_>�$?��->�m�=�)�>�7���P�B1�>p�@>Jh,>aB@?�M%?���
��ۣ��e/�\u>�W�>C��>��>!�J���=���>&a>	x �]���v���P>��X>FD|� q_�"�q� y=�d���g�=�=�=���A<���&=�?�?%Ɗ�򫆿R�ė.�ڔE?�%�>�-��>���2ɟ���;JG�?j4@�)�?(�C�L��)?T7�?�z�����=���>���=V��^�<�c�>�雽�j����I]����?���?�����P���y�4�=��L?0���Ph�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?GN>�֓?Z�M?�ο>��'��8�����i���	=�z/>A��>���>�ؔ���D�D���3���'h����UM	=��;�-�>�X�W[쾐m�=�^�={`Ͼ�����>�?�=�>aƦ>.��>rÛ>[o�>��<E���`�����K?���?����1n��[�<U��=�^��%?I4?�?[��Ͼ�֨>�\?���?6[?�a�>���>��迿�}��i��<%�K>�1�>�G�>����EK>O�Ծ<4D��p�>�ї>Yģ��=ھ-��Wh���A�>e!?���>N׮=Z� ?�#?O�j>c,�>�^E�V9����E�؝�>̘�>FN?Q�~?0?̹��X3�����桿R�[�� N>$�x?�O?(͕>&���~���IBG�/�H��,�����?�mg?DJ�d?C3�?��??w�A?tf>g��;�׾������>\�!?��ȺA�M&���\}?�P?��>7��W�ս�Pּ@��o����?�'\?n@&?c��I,a�J�¾�5�<z�"�ɈU����;��D���>ԍ>_���ύ�=o>Qݰ=BIm�WC6�l�f<5h�=A�>}�=�,7�6p�� ,?� �v̅��=&r���E��=�>��H>�¾��Z?�`<�]�z�k&���웿Y�S���?���?���?�)���h�/�=?��?�<?C�>ׯ��׾^ྋw��bg��^��>�-�>q���)(�7u��V����Ƃ�*9ݽ����?i��>�v5?���>�R�<��>[ܔ�؏��w׾"���N��<+���'�1��5(�N־/���%���Ӿ4,��w�>�DW��I�>{L?�->L�>9��>V��=��d>k�q>��>��>�@>n��=>50=�Z5�*��h�a?�����y:��% ���Z>A?��?�om>yRL>����T�'����>��?
�?�� ?��Z��s,���G?e1?$G���Y�>��ǽ����=\��4Ҹ��=�g��>Ac�/?�i�C�F����@�>�$?[4�<�Wƾ@5��#���RY�<��?m?8E5��C�3Si��=��V�S����P��/��5L�H�q�=��� ������Z�(�4u<�F2?��?�����;+ol�oI>�27>C�>�U>���>��r>m����,�r{R�C�ΟW��F?��?D��>�	H?VS6?dtV?�`?]<�>���>.�����>��=�^�>�?n1?8 ? ?�O?��&?�h[>p6���o �'/վ4� ?i ?E�?��>
��>M\�{;���-P�l����e�������M=��7=ɯսj����	=�L@>WU?G@�U�8�_���fk>5�7?$��>E��>Z菾*���K�<S"�>8�
? H�>�����zr��k��m�>l��?^���=��)>D��=�<���ź��=ɲ�����=4����;�՗<k��=���=N	p���b���:�Q�;c<�<�t�>J�?���>F�>�@���� ����>d�=tY>'S>�>�Eپ/~���$��K�g�<\y>gw�?�z�?дf=��=h��=
|���T��P��*���'��<��?(J#?�XT?���?5�=?wj#?�>�+��M��_��m���?g�+?���>1��^�ɾt�����3���?!?��`�̇���(�����0�Խ̚>�d/��&~������+D�d�����D����g�?G��?��G�#�6�=��I՘�9x��6�C?{7�>���>2�>��)���g���|,;>���>��Q?/»>C�P?��y?'�Y?��Q>g�7�W��� ˙���|�$>�2A?r�?<��?�7w?�(�>��>(P-�cY߾����1�%�������C=��_>P3�>���>h��>���=�=ҽ y���>�W�=��c>�v�>!ƥ>��>{z>'M�<��G?-��>&`������줾�ƃ��=�Λu?���?�+?�J=���	�E�ME���L�>�o�?���?R2*?��S����=�ּz඾��q��$�>׹>U3�>�Γ=�aF=�]>��>~��>�4��b��r8�yMM�u�?	F?'��=�1Ŀ����퇽q&����v�an׼ǌ5��H>Jy��<>P�~�C�J�B�{���vᢾ��y�������ʞv�<�>'��� >�3�=�T>��&��Ύ�=��<�#�T=膽R����	���o��8�.K-=S�r=�j=���]�|�g�?�?�>��}?`@�>�Q?K�G�[��>_g>>�P?�a(?�!�<�M��h.��0�ʾf��-"��#�4L���3�0>�O�=�T�>�xL>b�>���> �=/@�=�ͽiD���=�a�=��=xB>��)>O�=��>��u?�+j�E�C0�b�ѽ{� ?�ܦ=�;�<��Iy�>M5�=�*{�+��h����?�.@��?ӟ�>[�^�Y��>8͈������;(+>V'=�t<�2��jn�>��p>��5������d漐�?k�@,�C?�2��}�׿W��>��7>7�>��R�j1��W\�D�b�M*Z�-{!?�#;���˾bG�>»=�߾�{ƾ��,=��5>�>`=���^\�n��=	R{�fi<=��i=��><ID>��=Ai��l�=��I=�z�=ZP>5m��=t7���+�d(4=_��=o�b>�D&>"��>��?�a0?�Xd?�7�>�n�BϾ<?���I�>��=CF�>e�=�rB>���>��7?:�D?y�K?ᅲ>��=��>R�>l�,�Ĵm�\l�A̧�爬<ӗ�?�Ά?Ҹ>V�Q<c�A����{g>��-Ž�v??S1?vk?S�>#i
���ٿSn� 3%�FFH���=�Y�=�T���˽<؍���2���(� �>=�_>�v�>�*�>_��>Z�4>˸<>:�>�ˠ=w��<�P�=�Eh<�;T=�%h=��n=9l`�}��;�&ҽ����H��Ro�q->��Z�<#zK;�t�<�rH���>���>g;�=��?p)=1�߾Jʁ>����F���y=�����8���z��Xu�~�,�2�`�e!>N*>�G�N���Q?܁>��;>�Q�?�P`?1>>8�RY��Mσ�4!���B�4�>J�$><��^wK�̛x���?��`�p��>���>>�>�*m>�,��+?��x=��EX5��	�>�t�����n�@1q��<�����Qi���⺐�D?�D��^�=�~?̖I?�ߏ?���>���mؾ�b0>�)���v=>��p�����l�?h�&?Hf�>=�c�D�<d����ڽ06�>S^��.f�D����.-���w=���c]�>zU��+۾,4)�kn���#���<��fs���>x�A?t��?�Z㽢���Pu:�
����i�>�'B?ͥ;>�p�>O�?fݼ�>�u[w���>�Kv?)p�?u�?��K>�K�=�������>E�?N��?��?u�u?�iB���>�<_�*>��k����=�a>=�p�=;�	?=�	?0�?�v��l����뾀e���V�Ȃ�<O\�=��>�q�>�#x>��=mi=@:�=��W>W��>�c�>0�k>C~�>U�>�x��[;���?��^��Q�>��A?/�2=%�>S��=B*>���"�g�K�D�E�"�S���q)��9�)4>g};�ΰ�>����ʢ�?���=\R�FU ?˗5��Zx>�yE=,�>$Je>;!�>��>�)K>"��>�>�~t>��>�
<��ҾX>bk��<!��tC���Q���Ѿ�;|>�;��m�%��@�}P���6I����?��/�i�K1��YE=���<�I�?�����k���)��1�9�?O-�>Z5?VW���Z��ʼ>A��>F�>���hI��cs�����?�?��?c��>�-�>�X?��??���d���\���W�.Lf�W x�r=�u����~��3�����2*g?�
�?�T?>�";�o�>p�q?PwR�;�K����>]@���D����_�z>�r������3���WѾ"��u�>�~�?�ڊ?���>�M��wn�.�1>��8?ז2?��y?��0?H�@?���Z%?��K>r=?k�?�3?\�)?�>?��->���=p&�An=ƍ������i������Q.̼��=��x=O��<�L�<�a)=���;9�,}ݼ�>(��g��
�< �t=#	�=�u�=���>��]?nL�>t��>z�7?���1u8�Ʈ��+/?��9=ޫ������Ȣ�P�}�>w�j?���?�cZ?�`d>��A��
C�� >�W�>�v&><\>�b�>�h�;�E���=�G>�X>¥=�eM�x́���	�I������<&>ʌ	?�>)�����>���xaϾ xE>��Q��̣��f���*�
�+� ��}�>s�K?��3?�q�>-��q�E���d���%?C�@?7[�?A�R?uQ���罀+�DWT��!�j�>�F>�C�T��@����O��ut��_�=Au ��ՠ�R[b>����P޾�n�]J����2M=�z���V=�!���վ<�.��=�
>����<� �����Ԫ��'J?:mj=�o��JQU�`���>]��>�̮>7�:��.v�px@�����f<�=U��>��:>47��a��}G�7���>��>?��<?i�?ES��|���$������4��"@�=4�?�>�{�>:�3>����'P��4���[�j4Q�Y�>:m�>�O���H����A�t"(��߁>b��>��;>u�9?3n?r`�>SXA?�?Ь�>�^>P���Ȃ�qI&?>ك?~8S=�	�kM�%6�s�C�3��>F@*?��9�_�>6�?�?�E%?�QM??^��=@��M?�5��>���>��V��ⰿ�l>-�L?Zt�>��U?�w�?h6>Dg7��e��^���W��=�s">�{2?-"?��?O��>'o�>�e��+[�=���>rlb?yS�?vao?Y��=X�?��3>
�>~�=xR�>�!�>��?+M?��q?��J?�t�>�c�<~����:��OV��ʐ���y:g;<e�l=D����o��f���<�;�;�S��x�i�*�޼�C�]]�����;�}�>kt>dD��0.>�(žn�����C>�"���q��i���j8� *�='�>J�?ۤ�>�_$�n�=�B�>PT�>I����'?c�?��?���9:nb���۾O`J�%��>	�B?�\�=�@l�y����u���g=-}l?�]?��W������k^?��i?d���;�R$���dc����ml-?3	?+ߋ���>�?��m?���>�����r�?`���Q�ƣ���b=��>� ��6��9��>4db?<t�>��>@)>x������M���j3?���?͌�?O�?0�=|t<�R����C �nD���v?U�>-Y��}�8?�ȽJʧ�Q�оwJ�w���3�ƾ��ž~�۾�"��}�� ˾_F��.>ߎ?6��?2O??��M?�)*��^t�n�D������R�2o	�~��&4\��j?��@��
Z�t �=�����e��HY>�m��l��v�?���>��P-?��оG ���� �ey�>��B��V�Zޠ���`�]���tڗ=��оB�i��꾾V�*?���>1�>�w'?Li��@��"��L�(���Q�=���>��9>&��>'��p-���a�";ƾW��\Y�=ܥw>Db?rI?(p?Ճ���~2�@��Y� �r�-�K��>4>M�	>��>�<V�:"�ad'��M=��r�-�o^��Q�	��o=�%1?W��>��>�t�?�q?8O	�&˨�S�j���.�<0}<�}�>�^f?���>��}>�mؽ�� ����>
jh?�>���>�x{���3�4Hn�����4�>�ر>U�><"c>b��Q����������*��f�=jK?�掾>�i�.�>V�K?h�=�ن=׵u>G��j�
�32����	�e�=��?)>;9>y��|V'��*�����E�'?rw?q���1��>bb ?+��>�i�>�V�?�K�>���MJ�:@?��^?��B?H7?���>T=��^�Woѽ�����o=�z>��O>8W�=gO>�����Pb�7(�ʝo='"�=y4V�����?9<5~���@=�W=jOJ>wۿeZK�bپ���
�+
��	��V±�넇��+�c��;��(>x�����'��V�c&c�w�����l����?t,�?8$��
������6w��P����ǽ>Q�q���~�& ���^�(�����_Ǭ�AS!��O�=i���e�t�'?�����ǿ ���i-ܾ�" ?~C ?|�y?��|�"�Ȑ8��� >Ւ�<����@�뾽���9�ο������^?$��>M������>Y��>V�X>!lq>�
��F잾���<e�?L�-?��>1r���ɿ����=4�<:��?��@ikA?Z(���P=��>�	?xK@>ʞ1�����~��G��>-�?W�?�-O=}�W��Y�� e?�<5�F���&��=mm�=%�=r�7K>��>(~��/A��ݽJ{4>;�>s�&����K^�� �<Y�]>�Խ1���Ƿ�?vFX��g��e,�f!~�->xN?y�>�=�=0�%?k�A�g�Ͽb�^��<b?��?���?�w,?I�Ⱦ�]�>�ھ��J?�B5?�ޛ>�%���r����=��j�q��a"�f�T�y�=�@�>��=��9�iA���;�����l�=�����˿@���J8�vX :�=�!���<<�&�=����C�N!ĽM=��=�F=>��j>�8T>�2>�^?L,Q?q?E7>�{���Gw��a¾��=Y)���_���ÿ�� ���������������1F�)��!=�;�=	7R�n���,� �N�b�C�F���.?-w$>�ʾ��M���-<RpʾL����݄�^᥽�-̾�1�"n�_͟?��A?������V�1���U�����E�W?P�λ��ꬾ��=]�����=�$�>���=��� 3�f~S��+,?\�?����ґ�`%>ء�y��=}�*?��?;1=�/�>��%?����DȽ8�B>ky>��>���>��>�|��Xl����?�Q?�罯���F��>HQ��=Հ��=5�=� 0��_ݼwPU>F�l��G����.�9����eT<�V?��>I�*�QI��L���N��D=�v?�S?��>�
j?��B?|�<,��S� q��u_=8�V?�g?��>Vu���ξ)��7C6?�0f?�Y>ҳh�Q��h�.���D�?�l?i�?�`����{����"{���7?��v?�r^�qs�������V�6=�>�[�>���>��9�]k�>�>?1#��G�����^Y4�#Þ?��@���?D�;<|����=�;?s\�>��O�?ƾ~z��������q=�"�>(���Qev�����Q,�W�8?ؠ�?���>����ȩ�E��=�i��q^�?$�?~#��(�u<q���k�� ���<�5�=����t&����x�7���ƾ��Dޜ�Tų�g��>K\@�뽧"�>C�:��C�4"Ͽ"'���eоQ�r��?X�>��ɽ�ɣ���j� ,u�]�F��-H�bɋ�j�>�,>�4���o����|��a<�7�����>
j��z>�Y�z���姾d^;2)�>�Y�>��>�%��'�þ4\�?�:��� Ͽ\^��D���V?n�?\́?�"?�~f<m샾_g��Q��mL?l"x?B _?�j(�X�w�~���j?�^��aU`�F�4�HE��U>0#3?�B�>�-��|=>���>�g>k#/�R�Ŀwٶ�6���5��?��?�o꾗��>���?�s+?gi��7��N[��O�*���,�~<A?2>�����!�+0=�	Ғ���
?.~0?{�;.���d?*�&��Z���j�_�n�8��=N����
�W���ݾT�v�>��������?��@��?='�=|T{�Ϣ�>;,�>PM��������>���>nZ�>�}���?A���xþ8#�<J��?��?e?  ��s��D�f��Z�?�(�>�|�?�{�=�q_>ኃ>�"'�� �>i�>� >A`��W?��G?h?�o>	b���*�Uj;��5'�8y;�u6����=ģ�?�?
��>"�e��e�Ҿiwy���}t�t�g�K5{=��;�V+>��~>2�=$"��;���?p�1�ؿj���o'��54?\��>��?���K�t�����;_?\z�>�6��+���%���B�P��?�G�?#�?q�׾%P̼w>.�>�I�>z�ԽC���{���O�7>!�B?C��D��N�o���>���?�@�ծ?i��Q?��x���fs|��	��;��Y�=F�5?����jNn>C��>^�=Uw�}ϫ�4Wr�Vw�>e��?���?n�>�ul?�Aj�_1E�#'D=S�>|4g?�	??W�������y.>�?���wT���^ ���h?MD@W�@�(^?����y�K{���������>;|=��=��W��\�:qs>|'6<�[껞�=$X�>&JT>�mO>�'>`2�>���>0Â�t0'����q����G2�6���@0�Y��e`*��a¼G��^g�@SӾuK�\���+����V�1��]$�#T�=�T?�M?�}r?�` ?�����!>�$���3�<ʄ�B�a=�s�>�0?��I?�q%?-]=Bh����c��ҁ�
�sq�����><E>��>)�>�w�>���9>>~�@>Q��>	>1u�<C�O:<��<�(E>>��>���>vY�>�C<>ܑ>Eϴ��1��Z�h��
w�L̽)�?f���F�J��1���9�������h�=;b.?�{>���?п_����2H?���t)�*�+���>��0?�cW?�>����T�:>c��Ħj�Y`>�+ �jl���)��%Q>�l?&�f>u>I�3��]8�*�P�⁰�ah|>�/6?a涾�79���u��H��]ݾwGM>
��>��D��j�P������ti�!�{=]u:?˂?�2��eݰ��u�<C��TLR>C\>��=<|�=�SM>1Lc��ƽ�H�r3.=M��=?�^>%x ?��.>�D�=L"�>R����<a�N"�>#L>2fd>N@? ?E��<����'eS�H�2��)L>�S�>F/�>��
>�95�|=�=���>i�S>�_
��殽�a����{FL>���p�:�T��|V<3����=]�[=�3޽�fN�g��<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>�g��Z�������u���#=���>�5H?;N��6�O��>�Gv
?`?�X�$�����ȿ|v�K��>��?��?��m�`?��L@����><��?kY?�mi>�g۾�fZ�!��>��@?\R? �>77�!�'���?�ݶ?���?�xK>��?��p?7��>yLs� �0�v^��j����v=�1F<���>�j>Oξ�i�D�T�������Qj�0���1V>�[)=���>�轗 ��+ժ=�E��ި���e���>L�r>�V>�y�>�:�>���>��>��=9�������7#���!J?U��?��F�s�vc=o|�=��H��P�>}�7?��;ҧ;���>��]?~�|?�
N?���>c��B���D�������2=�eH>��>���>��ȼ�H�>�hӾ�16���x>k�>�r�}���zW�Ϩ�;��>yi ?w�>�&>�8!?�,?��>ۆ�>OC�g���o:����>v�>�"?�v�?� *?X+��?_(�3S���6����Z��(�=XQ?��?@��>�ˊ�����x��b)f=�+��Du?�l?�y�`l?t�?��C?�w?�&@>tཽҕվ����b�> /0?T�'��mg�$��^�I&?���>I�<o��;�᤾���=FJ� �	���=?s0�?�SK?5�_���G���_�<k��]�{=*�b=�v���`>��A>��;c�G>%}5>Y�1>!m��6��o����&=]RG>P.I>M�Z��-��45?q2�=�G����N>�pT�-�a��>�>��=N�ܾ&u?�-���Z�����4���)-��hy?!J�?u�?��^��[�L�!?\-�?�?�"�>uX�/߰��֚���E��>��)��> �-?���=�5�Aչ�%���x�}� ��<	��Hr�>��>�?�{�>�>c��>�ח��q �ۖ־���YU��Q���1���.�$+��(��v4����|���s���]�>6pr���>!?o�e>�W>� �>K�'=�C�>lW>�[~>�r�>,OF>K>ئ�=vߝ��h��O?<՛�Te-��!�����m�B?r�b?�U�>]8�,�{����?�j�?�l�?�N>4g���-�6�?��>1���1
?s>r=�
��rf=5}��>he�d��`:<��br>�R���8�O�Q���<�Zu?>�?�*<%漾�&˼:��c����?�[?%V3�3>?�بl�}�O��D[�aλ]�B�'���W'���x�?V����Ӛ���6'�0�=�j,?K!�?(��g�ھ	T�j0z�	�9�S
>��>��J>ok�>O��=G"��0�'�Q��[#�XD�^�?)L}?��>�NK?�;?�TK?r�Q?E�>ZE�>K��nO�>|��q�>0�>N�;?�5(?�(?�?7�!?21d>Cº�&��������?�:"?�?F1�>��>�fm�q���!�κi��dn{�|ᗽSyL=�f=�+��^�M��T\=��6>��?l*V=��3��,�V-�>��-?�? J�>>�ƽ�S0��~3=�Q�>V�	? ��>v� �{e���E��>$��?e���9>;*�>I�=hܨ���<��>Vl�= ׵�!l��v<M"�=~E�=���=��<��</V�=w��;��>« ?�L?Jl�>偑>�v���:�U�	�Y��=<DN>�E>���=�վ��j��de�#�o>�O�?S5�?r*=kB�=�g�=�����(���w�/��j�d<�?[�#?��\?�ǎ?o�<?:+?B>����?���|�����3�?C!,?L��>����ʾ���3�3�?�Z?z;a�ܷ��<)�}�¾��Խ}�>�[/� /~����ED�K?�����-������?���?�A���6��z�羘�LX��іC?� �>PX�>��>�)�,�g��&�%;>��>R?##�>K�O?�${?��[?�pT>F�8��!���ʙ�rV3�c.">��??\��?�?�y?iK�>o>��)�s� j��������ゾ��V=�Y>씒>5&�>{ȩ>Ԅ�=u�ǽ}��	�>���=u�b>�u�>{��>O��>DWw>܃�<O�R?���>-�]�ƾ{[���/Y��N4����>�5z?�dx>�=�4�јq�u���8�?έ?��?·?*^�E�=vG=r�i�����ё>�F�=�i?���>`�_�51=�>��?�$"���a�Ӭu���6���?�H�?eA�:�ο��L�L> ]޾ �>\
�>l˒��q>x����c�>#7�]�g��Ʃ�D���ݮ��,�o�����q���%��bF?#�W<b��>�l@>`>o^k>�i0<L��<�X�<bΏ��0=W�a7*�4>�7���f����Z��/��쮽�]�o?��5?�:?�JH?��#>�yD>���R�>�5<���>^�W>	�<����h�d�z(¾����}5ʾ�gԾy�S�6����a�=#G=@\ >;$.>�@�=}N
<��=��=!�
>7��=�̩�G%�=�c�=�<%=V^�=^� >b�=2�r?��k��{����2�9���?���=�8�2���?��=Mǉ�}��J����?NW�?��?���>Aү���>ҩ���'p�Hm�=>�m">1��Z[��\�?Ng>�/�o�|�|���>�?%�@�`?Ps���ݿ��=�7>�^>%�R�t�0��A\�pc�SNY��W!?F�:��~˾��>�=ď޾wƾ�+=�5>b$`=~��5G\�y��=��z��I:=C�k='��>JkC>M>�=����ɵ=_�I=��=ݛP>iЮ��U7��O.�j1=l�=�Yb>U�%>u4�>�?$
0?Krc?縸>��m�ؿ;���ˑ�>Qf�=ke�>m^�=�D>�o�>�~7?��C?
2K?�S�>rg�=�>�B�>͆,�Gm��@律���Ɯ<�I�?ϑ�?�Թ>��w<�<B�3@��Y>��Ž��?�'1?в?���>�� ῔�"��l2�##���	�,z�<a�Q ���RB�,��E/ӽ��=O�>]��>���>�Mu>�@=>��S>*��>sw>o�G=���=� f;4=���i�=A�� !=
c�F���ڬ���o�ʀϼ!��;��;p�;؜��*��=z��>G�>֡�>}ؖ=D\����->Y̕�&�K����=y�����@�n�b�+k}�t�.�2�9���C>ϞV>=��Nܑ���?#A]>�A>��?��t?��>�G��RѾ�n���ld�CR�Lm�=��>}�?��<�.�b���O�
Ҿ���>M��>S�>>m>��+�A?���w=���SM5�3�>�Ҍ�����;(q��6���h�K�ֺvD?d@���F�=�~?ګI?ڏ?ܔ�>�)��\cؾL�0>Ǜ��b�= ���'p�O��l�?I�&?���>j�L�D���ƾ<����>,�G���_�AD��}3��Ƽ��о�>:؜����R25��.��l��t>�����rE�>�Y?��?V�׽�΃���A�E��&`�a7�>ݜV?�Ʌ>��>k�?�����)������=Nl?{��?�]�?H�>��=ۭ���>N
?~�?���?��r?��9�85�>���;|�>Y��<c�=��>:��=� �=�?
?Z�
?F�?H��[��~����m�b����<d�=�3�>9p�>�@m>���=Ip=��=�+\>yN�>�x�>��b>�%�>C+�>����3
��6'?���="�>�2?�&�>D�d=^���A�<SE�<��#�Xĸ�v��� �<���7�U=)����>�+ǿ��?�W`>�f��;?�����Z���X>;RW>�V�^��>��@>7y>!)�>,,�>&�>�Ӊ>�M">�<Ӿ��>{��#c!��$C�RR���Ѿ�mz>)�����%�����]���3I�mf���h�j��-��=9=�S��<�D�?T���\�k�s�)�Q����?�b�>�6?�׌������>1��>��>�@��{����ō��`��?m��?��b>"�>��I?
�?���z/��_f��a��P��a�~���*������=����I�vt�fW?�*u?��[?P��=��>�?�5_�F~�M1�>ɫE��:C�h&ؽ�~>%�绡��X��/Z��
GN=��?\ɜ?'�?��>���է.=!�=��>�?��?Cfx>
sI?Z��>1O?G
M>�Ѝ>Ф;?^�Y?<�?;�=���$s��,�>㣂>�Y�������K��G�N����~8��"�������R=�w�=�X�<�Z�����=���=���<��g=��=$L6=[�>�]?�c�>�׆>��7?���p`8�RB����.?[5=W͂�c^���������>�j?C��?�
Z?(�b>��A���B�|f>c�>�s&>_�[>��>����E����=<>��>�v�=/�O�d����	������}�<�>{K�> q}>UF����)>喣�n�s��&X>d�b�ֵ�̴_�lC�4c4�?^��ɞ�>�O?�x ?���=��R<��
d�i�'?l;?��L?2G|?��=��׾��5��J�0�����> =�
���3Q����8�J�_<]�>����Ǡ�2�b>����ݾ��n��J��{羓vM=�n�FIV=p�S־G��M<�=M�	>���� ����<ժ�J?��k=�G��k�U�D��x�>a��>4�>wU:���u��t@�鉬��=�=���>~�:>�t��	�vG�!2�9��>L?$L?�V�?�n�6�x��X��t������U��=�M?���>���>0	>&��K.Ӿ����Cd�=HJ�(��>�,�>Y�	��D?��aؾ�վ��)���=�~�>(�S>�}3?�s?δ?�m-?^f?ٖ�>8ύ>,}�����:&?㋃?�ׄ=�ս��T���8��F�0��>0�)?�{B�M�>?-�?R�&?piQ?G�??�>�� �<J@��~�>�S�>��W�_���I`>��J?���>4Y?{Ճ?2�=>�{5�梾�Щ���='<>��2?�)#?��?Ȱ�>��>���=��>{c?u.�?�o?~|�=|�?;n2>���>h_�=���>
z�>Z?�QO?��s?3�J?���>�:�<�O��ⶽws���M���;��G<��z=���]�s�%�����<N�;B��������ND��S��?[�;��>��}>�	о=��;�G˾L����C�=�ٙ�8�U��ڰ����eļ#��>�i?���>�a`��d�=�V�>���>�x ��# ?�2�>�!?�l3<Ͽu����䲽,uW>��?R�P>�_M�l2���⃿-��?��u?ʎԾ�>���b?�^?�]�O=�C�þh�b����K�O?��
?��G���>��~?2�q?ɕ�>�,f��@n����[9b��k����=Zm�>�M�:�d��_�>��7?\F�>��b>H��=��۾
�w��m���?��?���?�?+*>y�n��$����L��p?9[�>�թ�@�8?h�^��	#���V��qH��;՘Ӿ|gѾ�������
D�`�Y�Ɯ�l�<�)?�i�?��w?�1N?���K�MN'���Y�2�9��d�?���Hm�t�K�_�:�&*L�x�����g]����C�O��sjB�]��?"�?�9���|�>�։�E�u�O�ƾ�=>=�O>��Y %�$�J��r��<@@o������۾J�6?���>p�>��?�k�S�C��7���*�Ń�i�=ϸ>^З>a��>]�(�c|D�f��ܾ��O�N�3�v>^�c?X�J?��m?�����0��5����!��)�������F>F�>���>r�X�[�ʱ&��>��`r�qd�����#i	��	�=�Z1?�ق>�ٞ>���?H�?�>��f����w�41���<�[�>��h?R�>PT�>vʽ6 �;��>i�l?��>�Ƞ>�����X!��D{�M`ν���>Ԅ�>l��>��r>F�+�m�[�c`�������B9�B�=|�g?>����_�Ŧ�>�'Q?x�:)�o<��>��y��
!�p��O�%�n	>}V?0��=��;>��ľ����z�;����Q)?�K?r쒾�*��#~>�'"?u�>o�>�2�?z"�>�lþ��?���?��^?kCJ?�FA?75�>+�=���_WȽ��&���,=�x�>A�Z>m=��=H���l\�[��čD=�K�=Oμ^����<@���V K<JT�<�3>�hۿ�JK�9mپW���8'
��刾���bX������X������gx�����'��V��)c�V���g�l����?9�?�X��)������ƍ��S���'��>��q��������V�;��w��U����b!���O�i��e�Q�'?�����ǿﰡ��:ܾ2! ?�A ?2�y?��4�"���8�� >�C�<\,����뾫����οB�����^?���>��/��j��>ҥ�>�X>�Hq>����螾�1�<��?7�-?��>Ɏr�/�ɿc���T¤<���?/�@<xA?��(�����WV=)��>�	?C�?>�^1�qD��簾�Y�><�?���?+eM=��W�-<
��oe?�
<X�F�T=޻��===�=7=����J>gJ�>֥�0VA��
ܽ��4>_�>8"����P�^�X\�<`�]>;�ս���!Մ?8y\�f���/��T��%P>��T?S(�>�@�=9�,?�7H��|Ͽ��\��*a?�0�?զ�?e�(?Kۿ�Lۚ>d�ܾƉM?�C6?���>�c&�+�t����=� ἴ��j��(#V���=��>�w>9�,����zO�ộ�i��=^k���ǿ���ʰ�=�߻�G�=����i�<:C�����<Ilx���M��j���<<Bz,=�h>z��>ԆE>�->4�K?Kgl?��>|:>C��[Qo������~��{T��DY������3Ͼw�Ҿmy������&�'��@��!=��=7R�j���9� �Y�b�L�F���.?w$>U�ʾ��M�â-<}pʾd���:܄�᥽�-̾�1�"n�h͟?��A?������V�T��vW�U���`�W?YP�Ļ�mꬾ���=���;�=%�>슢=���� 3��~S��o0?a?y~��BS��zP*>T� �k=��+?]�?��\<r2�>�S%?E�*�;�V:[>��3>\��>ê�>�	>���'�۽P�?��T?������aِ>�Z����z��ya=R8>^5����،[>�Q�<�ꌾ�T�K;����<�&W?Ϡ�>-�)�8��_��U���V==��x?��?�/�>F}k?��B?�<1h����S�$!�%:w=_�W?y%i?Q�>舁�
оA����5?[�e?�N>�\h���龙�.�[T��"?{�n?�^?�I���s}�D��H���n6?��v?s^�ps�����p�V�T=�>�[�>���>��9��k�>�>?�#��G������sY4�&Þ?��@���?��;<��X��=�;?m\�>��O��>ƾ9{�������q=�"�>���vev�����Q,�w�8?㠃?���>%���������=�ؕ�Z[�?�?I���,Bg<����l�o�����<٫=�1��Y"�����7���ƾ�
�����*r��L��>�X@Y���>Sa8��3�BRϿ`��>dоYq���?��>FȽ�����j��Lu�V�G���H�����Q�>�>���������{��s;��؟���>�����> �S�e(������`35<��>��>TÆ>�.��w彾�Ù?�]���Aο������ �X?�d�?qi�?�p?��9<�v��{��6��2G?B�s?�Z?~%�oT]���7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�/�n?Wk"�d(��C��dO�=U_�����E �?�{����D�w��y���S��N׷?1��?8��?��h<�L�j|L?��>�XV�ҟ㾋R�<�
L>��?{��>��:�)?2�r��C%�<�=H��?^_�??=�>�����ʛ�&�M>u(�?��>��?��=[��>B��=j���`D����>��>*T����?��P?$X�>t��=��R�&�2��H��O��@���?����>��[?�>?�/p>��E����Mf��Ӟ�'3���3�gD ����
н�"8>�>>:�>�v)�>ľ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��$	?[���g����x�b4�W�=��E�=W7?�w��U>U��>�=�|t��{��bq�H��>�S�?���?��>[�n?e��[L��}{=�4�>�*^?�w?�6P�=����*>��?�b	�Y������3�n?�n@��@]?+Y����ͿR-���j��S���
�=���=�c>�W����=_ap=����=k�>�T|>�%B>�xQ>Ȉ4>�YN>�;>>U�����%�أ�������?�������r�x�������&�x�������g��LoڽaϽ�W����@�4����=�Z?e�@?��k?PC?bq��U>�t�-6$=��׽a�=���>�?��C?�2?�Z��"���nk�dx���*��������>�H�=%�>6;�>ӣ�>?'8��'>��>��>٭�>!��=����s�;fYA>���>N�>���>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��u�T�4:>9����j�5`>�+ �~l���)��%Q>wl?'�f>�v>Cj3�-�7��ZP�S����1}>��5?i���1J8�#�u�1`H�cݾDqM>��>*�V��������a�`ci��py=Hc:?� ?t쳽�x����u����F�Q>R]>*� =�ְ=�9N>��d��ǽ�G��/=�7�=t;_>�$?��->�m�=�)�>�7���P�B1�>p�@>Jh,>aB@?�M%?���
��ۣ��e/�\u>�W�>C��>��>!�J���=���>&a>	x �]���v���P>��X>FD|� q_�"�q� y=�d���g�=�=�=���A<���&=�?�?%Ɗ�򫆿R�ė.�ڔE?�%�>�-��>���2ɟ���;JG�?j4@�)�?(�C�L��)?T7�?�z�����=���>���=V��^�<�c�>�雽�j����I]����?���?�����P���y�4�=��L?0���Ph�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?GN>�֓?Z�M?�ο>��'��8�����i���	=�z/>A��>���>�ؔ���D�D���3���'h����UM	=��;�-�>�X�W[쾐m�=�^�={`Ͼ�����>�?�=�>aƦ>.��>rÛ>[o�>��<E���`�����K?���?����1n��[�<U��=�^��%?I4?�?[��Ͼ�֨>�\?���?6[?�a�>���>��迿�}��i��<%�K>�1�>�G�>����EK>O�Ծ<4D��p�>�ї>Yģ��=ھ-��Wh���A�>e!?���>N׮=Z� ?�#?O�j>c,�>�^E�V9����E�؝�>̘�>FN?Q�~?0?̹��X3�����桿R�[�� N>$�x?�O?(͕>&���~���IBG�/�H��,�����?�mg?DJ�d?C3�?��??w�A?tf>g��;�׾������>\�!?��ȺA�M&���\}?�P?��>7��W�ս�Pּ@��o����?�'\?n@&?c��I,a�J�¾�5�<z�"�ɈU����;��D���>ԍ>_���ύ�=o>Qݰ=BIm�WC6�l�f<5h�=A�>}�=�,7�6p�� ,?� �v̅��=&r���E��=�>��H>�¾��Z?�`<�]�z�k&���웿Y�S���?���?���?�)���h�/�=?��?�<?C�>ׯ��׾^ྋw��bg��^��>�-�>q���)(�7u��V����Ƃ�*9ݽ����?i��>�v5?���>�R�<��>[ܔ�؏��w׾"���N��<+���'�1��5(�N־/���%���Ӿ4,��w�>�DW��I�>{L?�->L�>9��>V��=��d>k�q>��>��>�@>n��=>50=�Z5�*��h�a?�����y:��% ���Z>A?��?�om>yRL>����T�'����>��?
�?�� ?��Z��s,���G?e1?$G���Y�>��ǽ����=\��4Ҹ��=�g��>Ac�/?�i�C�F����@�>�$?[4�<�Wƾ@5��#���RY�<��?m?8E5��C�3Si��=��V�S����P��/��5L�H�q�=��� ������Z�(�4u<�F2?��?�����;+ol�oI>�27>C�>�U>���>��r>m����,�r{R�C�ΟW��F?��?D��>�	H?VS6?dtV?�`?]<�>���>.�����>��=�^�>�?n1?8 ? ?�O?��&?�h[>p6���o �'/վ4� ?i ?E�?��>
��>M\�{;���-P�l����e�������M=��7=ɯսj����	=�L@>WU?G@�U�8�_���fk>5�7?$��>E��>Z菾*���K�<S"�>8�
? H�>�����zr��k��m�>l��?^���=��)>D��=�<���ź��=ɲ�����=4����;�՗<k��=���=N	p���b���:�Q�;c<�<�t�>J�?���>F�>�@���� ����>d�=tY>'S>�>�Eپ/~���$��K�g�<\y>gw�?�z�?дf=��=h��=
|���T��P��*���'��<��?(J#?�XT?���?5�=?wj#?�>�+��M��_��m���?g�+?���>1��^�ɾt�����3���?!?��`�̇���(�����0�Խ̚>�d/��&~������+D�d�����D����g�?G��?��G�#�6�=��I՘�9x��6�C?{7�>���>2�>��)���g���|,;>���>��Q?/»>C�P?��y?'�Y?��Q>g�7�W��� ˙���|�$>�2A?r�?<��?�7w?�(�>��>(P-�cY߾����1�%�������C=��_>P3�>���>h��>���=�=ҽ y���>�W�=��c>�v�>!ƥ>��>{z>'M�<��G?-��>&`������줾�ƃ��=�Λu?���?�+?�J=���	�E�ME���L�>�o�?���?R2*?��S����=�ּz඾��q��$�>׹>U3�>�Γ=�aF=�]>��>~��>�4��b��r8�yMM�u�?	F?'��=�1Ŀ����퇽q&����v�an׼ǌ5��H>Jy��<>P�~�C�J�B�{���vᢾ��y�������ʞv�<�>'��� >�3�=�T>��&��Ύ�=��<�#�T=膽R����	���o��8�.K-=S�r=�j=���]�|�g�?�?�>��}?`@�>�Q?K�G�[��>_g>>�P?�a(?�!�<�M��h.��0�ʾf��-"��#�4L���3�0>�O�=�T�>�xL>b�>���> �=/@�=�ͽiD���=�a�=��=xB>��)>O�=��>��u?�+j�E�C0�b�ѽ{� ?�ܦ=�;�<��Iy�>M5�=�*{�+��h����?�.@��?ӟ�>[�^�Y��>8͈������;(+>V'=�t<�2��jn�>��p>��5������d漐�?k�@,�C?�2��}�׿W��>��7>7�>��R�j1��W\�D�b�M*Z�-{!?�#;���˾bG�>»=�߾�{ƾ��,=��5>�>`=���^\�n��=	R{�fi<=��i=��><ID>��=Ai��l�=��I=�z�=ZP>5m��=t7���+�d(4=_��=o�b>�D&>"��>��?�a0?�Xd?�7�>�n�BϾ<?���I�>��=CF�>e�=�rB>���>��7?:�D?y�K?ᅲ>��=��>R�>l�,�Ĵm�\l�A̧�爬<ӗ�?�Ά?Ҹ>V�Q<c�A����{g>��-Ž�v??S1?vk?S�>#i
���ٿSn� 3%�FFH���=�Y�=�T���˽<؍���2���(� �>=�_>�v�>�*�>_��>Z�4>˸<>:�>�ˠ=w��<�P�=�Eh<�;T=�%h=��n=9l`�}��;�&ҽ����H��Ro�q->��Z�<#zK;�t�<�rH���>���>g;�=��?p)=1�߾Jʁ>����F���y=�����8���z��Xu�~�,�2�`�e!>N*>�G�N���Q?܁>��;>�Q�?�P`?1>>8�RY��Mσ�4!���B�4�>J�$><��^wK�̛x���?��`�p��>���>>�>�*m>�,��+?��x=��EX5��	�>�t�����n�@1q��<�����Qi���⺐�D?�D��^�=�~?̖I?�ߏ?���>���mؾ�b0>�)���v=>��p�����l�?h�&?Hf�>=�c�D�<d����ڽ06�>S^��.f�D����.-���w=���c]�>zU��+۾,4)�kn���#���<��fs���>x�A?t��?�Z㽢���Pu:�
����i�>�'B?ͥ;>�p�>O�?fݼ�>�u[w���>�Kv?)p�?u�?��K>�K�=�������>E�?N��?��?u�u?�iB���>�<_�*>��k����=�a>=�p�=;�	?=�	?0�?�v��l����뾀e���V�Ȃ�<O\�=��>�q�>�#x>��=mi=@:�=��W>W��>�c�>0�k>C~�>U�>�x��[;���?��^��Q�>��A?/�2=%�>S��=B*>���"�g�K�D�E�"�S���q)��9�)4>g};�ΰ�>����ʢ�?���=\R�FU ?˗5��Zx>�yE=,�>$Je>;!�>��>�)K>"��>�>�~t>��>�
<��ҾX>bk��<!��tC���Q���Ѿ�;|>�;��m�%��@�}P���6I����?��/�i�K1��YE=���<�I�?�����k���)��1�9�?O-�>Z5?VW���Z��ʼ>A��>F�>���hI��cs�����?�?��?c��>�-�>�X?��??���d���\���W�.Lf�W x�r=�u����~��3�����2*g?�
�?�T?>�";�o�>p�q?PwR�;�K����>]@���D����_�z>�r������3���WѾ"��u�>�~�?�ڊ?���>�M��wn�.�1>��8?ז2?��y?��0?H�@?���Z%?��K>r=?k�?�3?\�)?�>?��->���=p&�An=ƍ������i������Q.̼��=��x=O��<�L�<�a)=���;9�,}ݼ�>(��g��
�< �t=#	�=�u�=���>��]?nL�>t��>z�7?���1u8�Ʈ��+/?��9=ޫ������Ȣ�P�}�>w�j?���?�cZ?�`d>��A��
C�� >�W�>�v&><\>�b�>�h�;�E���=�G>�X>¥=�eM�x́���	�I������<&>ʌ	?�>)�����>���xaϾ xE>��Q��̣��f���*�
�+� ��}�>s�K?��3?�q�>-��q�E���d���%?C�@?7[�?A�R?uQ���罀+�DWT��!�j�>�F>�C�T��@����O��ut��_�=Au �as���>d>�@
��پ��m�XK�����>I={��Mh=K��dԾ�Ȁ����=�A>����
r!�a���ު�V&H?�1]=jn���IO�O�����>��>DM�>���L�{�~�?��ګ��ġ=�
�>ݓ6>�������q�I��k��>�L?�.M?	��?�.��ju�Bt�����Q��‭=�"?�.�>G��>�>ͷK������e!�2af�0AJ�9��>R�?;����O�B����)ƾ�S��$�=G�>�3M>��M?I�L?���>��??kE?"��>(�> uB=�j�^k"?	��?�=��(� ��j�B�<��y�>?�*? ��}�>�?I;?�?�)?�y�>D��=��l�4�c�>�ƈ>uh[�� ��R.�>��q?��>��[?��?]�'>��?�����}*4�Jp�=H)$>�!1?�� ?�	?�C�>l<�>/�����=���>�-f?Ea�?s�q?d#>�a	?�>?��>��>DƘ>i7�>�?�C?"tt?S#F?���>uo�<�Iӽ
eѽL���kG~�����}�T�)��=ܲA�<���pFZ��^�<蠘;�o�����<N�����������eo<���>�X�>a(̾��=!۾�{��k>�����x�yω��l��q���B5�>�<4?�>�c��vrx=V��>KE�>��%?��>?�,�=��R�c����)��a�>]�P?Q�}>�`�a�����{���u:�[?Zm?f�x�)�
��b?H\_?�U�>��A���EX��F��fN?Ӳ?:8C�̸>A}~?��p?�2�>�k��^o������0`�g*j��&�=G�>����f����>��:?~��>��h>���=��ؾ7y����)�?&֋?��?B��?�C+>�l�\�޿�������� a?S��>{#���&?Z.��Լ�̭��?u��޾���(s���*��,8����&�L8��țɽ�Xh=D�?��n?��o?�6^?t� ���`�[�Y���~�۠R�S���?��G�&E���>�8�i��E��H�ݱ����<@���7�_�N��?3b�>��;�ے!?%;)a�P��vA?�P@��#��P�K��3�;*v��O��,���J�k� ���2?b��>�9�>��1?�}��ON�$�
���;�kl��8�>���>�D=���=������x6���˾H�վ�����P�>Ђd?4�=?�bq?��7�E���g�<�� ������w�=�>�k>>�l�[�C�G�"��MB�[c���E������
�?j�=��/?]p�>G�>	}�?l5?oоJ����tg��$���=Dʽ>f�V?l��>�/@>7b�(�(����>�%o?���>��>�a��U4���f�������>�j�>��>r}>�R��Z�#=��/0���C5�d�=*VL?wُ���p�|�>�R?`#��_���5�>|�<�U��Ѹ־?�J����=U�?5>Ts�=��վ���<��=ܦ�D4)?�t?�,��?,��Q�>m�#?�I�>,�>5r�?a��>PG��`t�U4?�/^?2�H?��?? ��>?:*=p簽c�˽�4*�?M==ֈ>�*]>qt=���=�Z�"�Y��y��JB=w��=��（c���,+<PR���z[<h��<��0>;mۿ-EK�X�پ����P<
�舾����d������b��Q���Tx�u���
'�*V�@5c�䞌��l�υ�?l;�?�|��q.��h���[���-�����>��q���򫾇�� %����о���c!�z�O�>#i�'�e�O�'?�����ǿ𰡿�:ܾ3! ?�A ?7�y?��6�"���8�� >\C�<-����뾭����οF�����^?���>��/��m��>ޥ�>�X>�Hq>����螾�1�<��?7�-?��>��r�0�ɿc���¤<���?0�@1KA?@w'�J�쾌)G=���>� 
?ܜ?>z�0���	������>8�?�Ҋ?�dH=&�W������d?W&<�F�\B���=?��=P�
=���qN>ڬ�>B%�Q=�U�ڽ��0>]�>2�����5]�5U�<~�\>��ӽ\Ŕ���?��W�/�g��1�����7>�NR?��>R	�=�*?�H���Ͽ�\Y�<�e?���?^��?��'?�л���>��ܾ�eL?�5?�2�>�i"��r�n��=�^ּ#�(���۾BO��;�=H}�>��	>�0�,�N�<��Ӽ��=�M��QmɿП�mj/��K�;z�=��E���=��(=e����DL�A/����=�ڨ=�>�m�>�Γ>��S>��T?Z7:?v5?�Q>�ę;�Eƽܷ����<�Ѿ�T޽ ����3�������X�ѾSG��D�����}��� =�`�=�6R�0���.� ���b���F���.?v$>��ʾ��M���-<�pʾ�����ℼ$⥽�-̾�1�"n�*͟?P�A?������V�<���Y�6���u�W?nN�����ꬾ��=+���4�=x$�>;��=��#!3��~S���+?�h$?�U��q��*�r>\���蓬=~V(?��?"�=�>��'?at��x��c�/>_ 
>k�>0��>��=OF������-?Md`?|������%�>�j��/Ԉ��"><���=X1<�P	�p�T>>�O=]S��"��zK��Pn=>�R?{-�>�")�S&�[Y���<��7= o?��?M��>�q?}HB?��-=e����	V�v�:�=��Q?i$\?�n�=ܢ����վ�����9?��q?�[�>37��ܹ��#�b)�Ӯ?D�i?u�?y�����f�3=��8�����-?��v?�r^�<s�������V��;�>$Z�>��>o�9�bi�>��>?�#��G��㺿�Y4�7Þ?��@���?d�;<^����=�:?�\�>;�O��>ƾ���������q=� �>�����dv�6���O,���8?1��?���>攂���.��=å��[L�?��?�]��0]<8��1�k��S��=�<�P�=�|�R<$�0���7�Q7Ǿj�
����Yʼ�Ȇ>�F@}���>9�R⿌WϿ����Uо��p�H?b��>ԪȽ����v�j�gu��sG���H��"��du�>8�>�H��w�����{�k|;��_����>��	�vv�>��S�):��ᱟ��-4<"%�>���>��>Ȯ�7������?�_���@ο�����v��X?�N�?}3�?��?|�A<3�w���{�?��.FG?�s?�Z?W�(�,9^���7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�d�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.���w?�f������3ؾە���}�7P��L�4��>�aA�G���������<x��?��@���?*��G�#�\a?BD�>������	�0�Ծ^�=>��>���>�	W�"}?+	ɾNMG��	J�Y��?��?�?�tb�w4��)<�=+�?K��>�E�?R �=/�>�]q>����W:>
�7>�0O>��Z;���>��G?x��>��������i�&�`�N�m�o�{=�)S1����=fi?SbJ?1��>�����x=�ؾĳ���&L��ε<]���~l�[��y�A>|�0>���=	d(�=i����?Gp�8�ؿj��p'��54?/��>�?��{�t����;_?Rz�>�6��+���%���B�_��?�G�?<�?��׾�R̼�>?�>�I�> �Խ����T�����7>+�B?Z��D��s�o�z�>���?�@�ծ?hi�P	?���B��A~�����V7�l�=��7?�Y�~�z>>��>Yn�=�}v�滪���s����>NE�?��?s��>ʧl?RQo�C��>3=c��>Ftk?�_?�{�%���A>�?��������C�<;f?��
@�w@��^?>颿Пտ�ė��x����־�&�;6-�A�4>�.w��n>[�&>���<�x����=E�I>�,>8�=�NA>9,c>ʉ�>�����d$�U���6����'�5�l�Í<�OX���Y�2,侐Wξ�{�V���Fg�5�H�7��J���]�=X�T?�M?�q?�?�����M?>�P�7=N���XL=���>A�-?:E?(� ?�HV=�°�z�m����<���hM���$�>E:;>o��>���>e�>/NQ�� K>=0L>�א>ė>m�=��f<�!�<(r$>]�>��>���>�C<>��>Fϴ��1��j�h��
w�l̽1�?����S�J��1���9��Ԧ���h�=Gb.?|>���?пf����2H?&���z)��+���>}�0?�cW? �> ��v�T�5:>8����j�6`>�+ �~l���)��%Q>wl?��f>�u>hO3�H�7�cP��ְ�Չ}>g6?������8���u��;H�	$ݾ��L>��>��P�P�����A3�/Ei���{=ft:?L?�汽r����Yv��D��ؔR>~�\>�{=H�=_M>T`�7ǽ�PI��Y-=�c�=f1_>�G?s�->맍=��>���(5N���>�B>z�->o�??S	%?�������̃��/��7u>e��>���>	6>7�J�8��=]��>�'c>m���'���N�6>�˒W>�K�q`�f�u��B{=�����=
ʕ=� �q�=���$=�^�?���$������W��O0?�S�>_��j[~=۴=��P������n�?�,@H�?�Y��#�Z��� ?��?5����S3>ĸ�>^�=>H����i"�`�+?��
f��\��_#-�'��?���?Ѿ�;X����	T�ia>=!?+ؾ�h�>|q�&Z�������u��#=Z��>8H?�S���O� >�+w
?�?�^򾾩����ȿ,{v�{��>n�?��?��m�dA���@�	��>���?hY?�ri>6c۾=^Z����>Y�@?vR? �>�8�p�'�D�?�޶?T��?5�Q>@e�?��j?���>����0����ɲ�����=ti=�y�>n�,>(���!A�+Γ��݌��"h�o��%x9>uH=���>T���־7��=|�D�쪼�1(}�O�>�\>��>qV�>> ?,��>T�>�,R<v�w�Z�U����K?-��?k���2n��4�<G��=̨^��?�H4?%M[���Ͼ?Ȩ>?�\?�À?6[?Yh�>����;��俿�}���<��K>�1�>9K�>-!��_MK> �Ծ�4D�bv�>Rۗ>�ң��Kھ%3��y���>�>gg!?6��>⽮=$�?�j-?hNY>:�>a�4�Y�����B�E�>�/�>Lk?	f�?�%?�j����.�����g,���4W�H�2>2xg?/?Q�>$:��F���K�<�*�=�����|?7�i?����?��?�A;?&�4?s\>V�=���s?D�1��>�6"?S��8bB���&�*o�# ?ؤ?���>�֏���׽J�������+��P�?x�\?>�&?�d� �_�E����&�<:{��9.����;��!��$>�a>����=�=�6>K�=�5n��~;��8<���=H�>��=�7��}�0?�9�=9԰��'�=�M��^B��nO>��8=�L���@?b)��HS��������:-���?\�?5�?����X���/?v��?�>(?v:�>��#X��W���㚾�G��]����>�u�>�5��)�s�������oRf�wi#����9H ?��>�B?���>�~>D�>�����"����f��I�R�u�t7�Z�/�����ﭾ�x� д��-ž,Ɂ���>1Z}�R��>|!?�x>;��>~�>�^b�-,�>�vW>s:�>
��>�R>A/)>�}�=���u�߽�hR?�0��c(��V龿��B?��c?E��>,cf�҄��z$�|�?��?���?}x>��g��)+��?��>� ���{
?j;=����ʍ<o*���H����EL�䓏>ӽyL:�d+M�\pf�
?��?�7��S̾Y�ٽ�f�ﶽ]L�?æ?�#V�$�<�r�o�$�6��f]�H�=�+����or@�K�`�'N������$>����H���C�H�1?ej�?��"<Ǿ�%�ޑp���J�D[+==��>V2>�r�>�ޘ>?����/�^W�#��==�f�?�s�?�׊>\
I?��;?o�I?eDV?F�>� �>-�����?�}ۻڰ�>���>�9?2?�c?�n	?U�$?��e>
}���쾷�?z�&?��?���>��>	k}��p��y�M����I�l������=~&I<�+��F2&<���=f�Y>��?�����"9�[n����>��G?���>i$�>s�=��I��҂=t��>��?3ly>���i t������>��r?�s:�[貼�>>M� >�<��=�'>ר�;���=�-��($�� �<��=bCv=�"�<��l=5%ļF�¡<i?
e"?>e}>���>sF��%��{�	�^��=IP/>�M>��>�&;71���H��M�d��Mp>�(�?.��?�{0=���=Ѹ�=�;��'�U#�zѾ�c=~�? #?�R?�?�)<?-,?�S
>����ܕ�ㅉ��7����?j,?)��>^��H�ʾ�쨿K�3�G�?>Y?�7a�ʱ�;)��¾��Խ��>�[/�-~�����D�������=x�����?��?�A���6�#z辿���R���C?T)�>}Y�>{�>�)���g�l)�$;>���>*
R?'�>��O?}'{?&�[?S�T>�8�2)���˙��h2�3">�;@?c��?��?��x?�;�>A>�)��]U��A��j����ǨT=?*Z>��>W	�>C�>�s�=�=ȽQ��v?����=db>��>a��>e�>d�w>�ְ<�H?+��>����2~�!?�������H?�&�s?���?c+?�J=�\��G�4����>t�?�E�?7�)?5�S�HO�=D.ϼUf���om�o��>b.�>���>��=PD0=ڤ>��>V��>������O9�D-_�f�?��E?L��=v~���G��a6��zž��B��ܛ��߄�E�
>���ݾ>З���J�7�K�� F��א��ϓ��ɱ��.��Ek�b%?t�>���>f	>!E�=Ҩ�=���ɍ�9��{>�n=5[������{���|����<1�����<l��a��}�x??@?�,-?wI?L{>�7y>dp��ܵ�>���
?��{>?�c��)����\�����Ǡ������E��i�n���C�A>�N�;��&>�l+>L��=t��<���=I!=̎�=�<�^=B>�Ʈ=�6=\&>a�:><�)>��t?�5h�p�������2�K_?E�=F���Q\
�O��>8>��ӹ�0�	��?�^�?�`�?��?�7���r�>M^����a����=��=�h:>)F��5��ɻ�>�YQ>�S+��Ќ����= ��?|	@�-M?nY���(ڿ���=q�7>��>L�R�`J1��\�x�b��Y��!?�!;�� ̾B�>���=�޾r�ƾ��,=)6>8_=����o\��|�=?r{�o	==4|k=��>�aD>5;�=�̯�1��=-J=��=7�O>�N����6���+��(2=�d�=Y�b>�:&>���>�?,]0?Qd?N;�>��m�Ͼ==���L�>�$�=�U�>_�=�uB>��>3�7?e�D?m�K?ق�> ��=K�>n�>Ŝ,��m�`����:�<��?І?8θ>D�P<j�A�6��e>��%Ž�v?nR1?;l?�>H7���ҿ�5'��^_�����&ڽ���=���<ˮ =kJ��|>������Q�=�,F>Nx~>"��=��>J�M>?k�>�X�>���=�u�=�P��Ѐ����=�	X=>��>�_�$��X|��D=7C�=A�=Nq �g��;V��3�=Tn���=�!�>��>���>\ߕ=§��̣/>�����L�	"�=�}����A�!d�e8~��	/���6���A>t�V>�M���'����?CLZ>��?>�b�?��t?'� >����Ծ�.���He��S���=�	>9C=�Kl;��o`��*N��Ҿ�>M��>>B3n>��+�з?�./|=��ᾟY5���>����@�\���q�����ş�g
i�qj��ϺC?{/��<2�=��}?F�I?���?|��>�i����־�2>���=����n�fߐ�!{?��&?���>'���D��~��$N̽���>s*���_� �����6�~FK���ʾ�N�>����d׾�(:�c���T萿��A���k��P�>��M?�Ϫ?��ؽ3󆿆�=�1I�Ɂ��G�>"_?`�>
%�>�o ?��꽏��ψ���>��?]8�?ٳ�?2�7>�
�=� �� /�>�{�>�>�?��?�o?G��� ?π��i�g>dڙ<X��=y��=[Cs<,�==i??��?��?�����3���澭��^�[��wU=N6�=x.�>��>^E>U:=s.`=B.�=�RT>L��>�e�>R�5>{?�>*g�>����h��$?/�=�`�>i2?�σ>��=�����=�l�2�8���L5����5̑<{`�P|�=2�����>��ſ��?XH_>�q ��?����5��X�4>ŒT>0�� �>S�C>ɳu>̧�>Ȫ�>8�>���>��>�0Ӿ�>t���H!�%C�ȁR�3�Ѿhwz>䎜��%�E�����=I��f���k��j�Q2��J=��%�<u@�?S����k���)�+����?��>��5?Kь�s����!>Y��>ڹ�>a1��6����ʍ��N���?N��?DL�>�>�)E?��)?�Aɾ,﷾�>m�v�V��{h���u���:�'B���!��މ"�RH�;Y??�z?�|�<�)�>��?r�c��9���� ?�:��oB��	(�~�	>��'��s��F0پ��(���˜?���?	A�?s�#?Dɓ�8ג<�n�=�9?6	9?��v?��?~`?"��>�,R?�<�O?wzM?��3?�>]90>Rp:��V>���=��>��+�S��c�BM��l�ϳ7�8�.=J�6=��j=�>"7�<�t��|���7�v�<�;�&&=�=�`�=
զ>�]?���>Ѓ�>��7?��� b8�0ꮾ-
/?��9=5������!��) �
>J�j?k�?�PZ?wd>]�A���B��d>m��>�&>ޚ[>Pf�>�/�YF�(��=v>w,>`�=�gP�S%��t�	�����@�<��>�?T�>�ŧ��pH�̜��V��>�Y���:��R��\�$�gdH�ݑ����?v.j?V6Q?i�>AA׾[9�;M��?�0?ߎ_?h*�?�*��*#��7����x���ν�9�>q��>ʀ]���ʿG����G9��DO>��>����ՠ�R[b>����P޾�n�]J����2M=�z���V=�!���վ<�.��=�
>����<� �����Ԫ��'J?:mj=�o��JQU�`���>]��>�̮>7�:��.v�px@�����f<�=U��>��:>47��a��}G�7���>��>?��<?i�?ES��|���$������4��"@�=4�?�>�{�>:�3>����'P��4���[�j4Q�Y�>:m�>�O���H����A�t"(��߁>b��>��;>u�9?3n?r`�>SXA?�?Ь�>�^>P���Ȃ�qI&?>ك?~8S=�	�kM�%6�s�C�3��>F@*?��9�_�>6�?�?�E%?�QM??^��=@��M?�5��>���>��V��ⰿ�l>-�L?Zt�>��U?�w�?h6>Dg7��e��^���W��=�s">�{2?-"?��?O��>'o�>�e��+[�=���>rlb?yS�?vao?Y��=X�?��3>
�>~�=xR�>�!�>��?+M?��q?��J?�t�>�c�<~����:��OV��ʐ���y:g;<e�l=D����o��f���<�;�;�S��x�i�*�޼�C�]]�����;�}�>kt>dD��0.>�(žn�����C>�"���q��i���j8� *�='�>J�?ۤ�>�_$�n�=�B�>PT�>I����'?c�?��?���9:nb���۾O`J�%��>	�B?�\�=�@l�y����u���g=-}l?�]?��W������k^?��i?d���;�R$���dc����ml-?3	?+ߋ���>�?��m?���>�����r�?`���Q�ƣ���b=��>� ��6��9��>4db?<t�>��>@)>x������M���j3?���?͌�?O�?0�=|t<�R����C �nD���v?U�>-Y��}�8?�ȽJʧ�Q�оwJ�w���3�ƾ��ž~�۾�"��}�� ˾_F��.>ߎ?6��?2O??��M?�)*��^t�n�D������R�2o	�~��&4\��j?��@��
Z�t �=�����e��HY>�m��l��v�?���>��P-?��оG ���� �ey�>��B��V�Zޠ���`�]���tڗ=��оB�i��꾾V�*?���>1�>�w'?Li��@��"��L�(���Q�=���>��9>&��>'��p-���a�";ƾW��\Y�=ܥw>Db?rI?(p?Ճ���~2�@��Y� �r�-�K��>4>M�	>��>�<V�:"�ad'��M=��r�-�o^��Q�	��o=�%1?W��>��>�t�?�q?8O	�&˨�S�j���.�<0}<�}�>�^f?���>��}>�mؽ�� ����>
jh?�>���>�x{���3�4Hn�����4�>�ر>U�><"c>b��Q����������*��f�=jK?�掾>�i�.�>V�K?h�=�ن=׵u>G��j�
�32����	�e�=��?)>;9>y��|V'��*�����E�'?rw?q���1��>bb ?+��>�i�>�V�?�K�>���MJ�:@?��^?��B?H7?���>T=��^�Woѽ�����o=�z>��O>8W�=gO>�����Pb�7(�ʝo='"�=y4V�����?9<5~���@=�W=jOJ>wۿeZK�bپ���
�+
��	��V±�넇��+�c��;��(>x�����'��V�c&c�w�����l����?t,�?8$��
������6w��P����ǽ>Q�q���~�& ���^�(�����_Ǭ�AS!��O�=i���e�t�'?�����ǿ ���i-ܾ�" ?~C ?|�y?��|�"�Ȑ8��� >Ւ�<����@�뾽���9�ο������^?$��>M������>Y��>V�X>!lq>�
��F잾���<e�?L�-?��>1r���ɿ����=4�<:��?��@ikA?Z(���P=��>�	?xK@>ʞ1�����~��G��>-�?W�?�-O=}�W��Y�� e?�<5�F���&��=mm�=%�=r�7K>��>(~��/A��ݽJ{4>;�>s�&����K^�� �<Y�]>�Խ1���Ƿ�?vFX��g��e,�f!~�->xN?y�>�=�=0�%?k�A�g�Ͽb�^��<b?��?���?�w,?I�Ⱦ�]�>�ھ��J?�B5?�ޛ>�%���r����=��j�q��a"�f�T�y�=�@�>��=��9�iA���;�����l�=�����˿@���J8�vX :�=�!���<<�&�=����C�N!ĽM=��=�F=>��j>�8T>�2>�^?L,Q?q?E7>�{���Gw��a¾��=Y)���_���ÿ�� ���������������1F�)��!=�;�=	7R�n���,� �N�b�C�F���.?-w$>�ʾ��M���-<RpʾL����݄�^᥽�-̾�1�"n�_͟?��A?������V�1���U�����E�W?P�λ��ꬾ��=]�����=�$�>���=��� 3�f~S��+,?\�?����ґ�`%>ء�y��=}�*?��?;1=�/�>��%?����DȽ8�B>ky>��>���>��>�|��Xl����?�Q?�罯���F��>HQ��=Հ��=5�=� 0��_ݼwPU>F�l��G����.�9����eT<�V?��>I�*�QI��L���N��D=�v?�S?��>�
j?��B?|�<,��S� q��u_=8�V?�g?��>Vu���ξ)��7C6?�0f?�Y>ҳh�Q��h�.���D�?�l?i�?�`����{����"{���7?��v?�r^�qs�������V�6=�>�[�>���>��9�]k�>�>?1#��G�����^Y4�#Þ?��@���?D�;<|����=�;?s\�>��O�?ƾ~z��������q=�"�>(���Qev�����Q,�W�8?ؠ�?���>����ȩ�E��=�i��q^�?$�?~#��(�u<q���k�� ���<�5�=����t&����x�7���ƾ��Dޜ�Tų�g��>K\@�뽧"�>C�:��C�4"Ͽ"'���eоQ�r��?X�>��ɽ�ɣ���j� ,u�]�F��-H�bɋ�j�>�,>�4���o����|��a<�7�����>
j��z>�Y�z���姾d^;2)�>�Y�>��>�%��'�þ4\�?�:��� Ͽ\^��D���V?n�?\́?�"?�~f<m샾_g��Q��mL?l"x?B _?�j(�X�w�~���j?�^��aU`�F�4�HE��U>0#3?�B�>�-��|=>���>�g>k#/�R�Ŀwٶ�6���5��?��?�o꾗��>���?�s+?gi��7��N[��O�*���,�~<A?2>�����!�+0=�	Ғ���
?.~0?{�;.���d?*�&��Z���j�_�n�8��=N����
�W���ݾT�v�>��������?��@��?='�=|T{�Ϣ�>;,�>PM��������>���>nZ�>�}���?A���xþ8#�<J��?��?e?  ��s��D�f��Z�?�(�>�|�?�{�=�q_>ኃ>�"'�� �>i�>� >A`��W?��G?h?�o>	b���*�Uj;��5'�8y;�u6����=ģ�?�?
��>"�e��e�Ҿiwy���}t�t�g�K5{=��;�V+>��~>2�=$"��;���?p�1�ؿj���o'��54?\��>��?���K�t�����;_?\z�>�6��+���%���B�P��?�G�?#�?q�׾%P̼w>.�>�I�>z�ԽC���{���O�7>!�B?C��D��N�o���>���?�@�ծ?i��Q?��x���fs|��	��;��Y�=F�5?����jNn>C��>^�=Uw�}ϫ�4Wr�Vw�>e��?���?n�>�ul?�Aj�_1E�#'D=S�>|4g?�	??W�������y.>�?���wT���^ ���h?MD@W�@�(^?����y�K{���������>;|=��=��W��\�:qs>|'6<�[껞�=$X�>&JT>�mO>�'>`2�>���>0Â�t0'����q����G2�6���@0�Y��e`*��a¼G��^g�@SӾuK�\���+����V�1��]$�#T�=�T?�M?�}r?�` ?�����!>�$���3�<ʄ�B�a=�s�>�0?��I?�q%?-]=Bh����c��ҁ�
�sq�����><E>��>)�>�w�>���9>>~�@>Q��>	>1u�<C�O:<��<�(E>>��>���>vY�>�C<>ܑ>Eϴ��1��Z�h��
w�L̽)�?f���F�J��1���9�������h�=;b.?�{>���?п_����2H?���t)�*�+���>��0?�cW?�>����T�:>c��Ħj�Y`>�+ �jl���)��%Q>�l?&�f>u>I�3��]8�*�P�⁰�ah|>�/6?a涾�79���u��H��]ݾwGM>
��>��D��j�P������ti�!�{=]u:?˂?�2��eݰ��u�<C��TLR>C\>��=<|�=�SM>1Lc��ƽ�H�r3.=M��=?�^>%x ?��.>�D�=L"�>R����<a�N"�>#L>2fd>N@? ?E��<����'eS�H�2��)L>�S�>F/�>��
>�95�|=�=���>i�S>�_
��殽�a����{FL>���p�:�T��|V<3����=]�[=�3޽�fN�g��<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>�g��Z�������u���#=���>�5H?;N��6�O��>�Gv
?`?�X�$�����ȿ|v�K��>��?��?��m�`?��L@����><��?kY?�mi>�g۾�fZ�!��>��@?\R? �>77�!�'���?�ݶ?���?�xK>��?��p?7��>yLs� �0�v^��j����v=�1F<���>�j>Oξ�i�D�T�������Qj�0���1V>�[)=���>�轗 ��+ժ=�E��ި���e���>L�r>�V>�y�>�:�>���>��>��=9�������7#���!J?U��?��F�s�vc=o|�=��H��P�>}�7?��;ҧ;���>��]?~�|?�
N?���>c��B���D�������2=�eH>��>���>��ȼ�H�>�hӾ�16���x>k�>�r�}���zW�Ϩ�;��>yi ?w�>�&>�8!?�,?��>ۆ�>OC�g���o:����>v�>�"?�v�?� *?X+��?_(�3S���6����Z��(�=XQ?��?@��>�ˊ�����x��b)f=�+��Du?�l?�y�`l?t�?��C?�w?�&@>tཽҕվ����b�> /0?T�'��mg�$��^�I&?���>I�<o��;�᤾���=FJ� �	���=?s0�?�SK?5�_���G���_�<k��]�{=*�b=�v���`>��A>��;c�G>%}5>Y�1>!m��6��o����&=]RG>P.I>M�Z��-��45?q2�=�G����N>�pT�-�a��>�>��=N�ܾ&u?�-���Z�����4���)-��hy?!J�?u�?��^��[�L�!?\-�?�?�"�>uX�/߰��֚���E��>��)��> �-?���=�5�Aչ�%���x�}� ��<	��Hr�>��>�?�{�>�>c��>�ח��q �ۖ־���YU��Q���1���.�$+��(��v4����|���s���]�>6pr���>!?o�e>�W>� �>K�'=�C�>lW>�[~>�r�>,OF>K>ئ�=vߝ��h��O?<՛�Te-��!�����m�B?r�b?�U�>]8�,�{����?�j�?�l�?�N>4g���-�6�?��>1���1
?s>r=�
��rf=5}��>he�d��`:<��br>�R���8�O�Q���<�Zu?>�?�*<%漾�&˼:��c����?�[?%V3�3>?�بl�}�O��D[�aλ]�B�'���W'���x�?V����Ӛ���6'�0�=�j,?K!�?(��g�ھ	T�j0z�	�9�S
>��>��J>ok�>O��=G"��0�'�Q��[#�XD�^�?)L}?��>�NK?�;?�TK?r�Q?E�>ZE�>K��nO�>|��q�>0�>N�;?�5(?�(?�?7�!?21d>Cº�&��������?�:"?�?F1�>��>�fm�q���!�κi��dn{�|ᗽSyL=�f=�+��^�M��T\=��6>��?l*V=��3��,�V-�>��-?�? J�>>�ƽ�S0��~3=�Q�>V�	? ��>v� �{e���E��>$��?e���9>;*�>I�=hܨ���<��>Vl�= ׵�!l��v<M"�=~E�=���=��<��</V�=w��;��>« ?�L?Jl�>偑>�v���:�U�	�Y��=<DN>�E>���=�վ��j��de�#�o>�O�?S5�?r*=kB�=�g�=�����(���w�/��j�d<�?[�#?��\?�ǎ?o�<?:+?B>����?���|�����3�?C!,?L��>����ʾ���3�3�?�Z?z;a�ܷ��<)�}�¾��Խ}�>�[/� /~����ED�K?�����-������?���?�A���6��z�羘�LX��іC?� �>PX�>��>�)�,�g��&�%;>��>R?##�>K�O?�${?��[?�pT>F�8��!���ʙ�rV3�c.">��??\��?�?�y?iK�>o>��)�s� j��������ゾ��V=�Y>씒>5&�>{ȩ>Ԅ�=u�ǽ}��	�>���=u�b>�u�>{��>O��>DWw>܃�<O�R?���>-�]�ƾ{[���/Y��N4����>�5z?�dx>�=�4�јq�u���8�?έ?��?·?*^�E�=vG=r�i�����ё>�F�=�i?���>`�_�51=�>��?�$"���a�Ӭu���6���?�H�?eA�:�ο��L�L> ]޾ �>\
�>l˒��q>x����c�>#7�]�g��Ʃ�D���ݮ��,�o�����q���%��bF?#�W<b��>�l@>`>o^k>�i0<L��<�X�<bΏ��0=W�a7*�4>�7���f����Z��/��쮽�]�o?��5?�:?�JH?��#>�yD>���R�>�5<���>^�W>	�<����h�d�z(¾����}5ʾ�gԾy�S�6����a�=#G=@\ >;$.>�@�=}N
<��=��=!�
>7��=�̩�G%�=�c�=�<%=V^�=^� >b�=2�r?��k��{����2�9���?���=�8�2���?��=Mǉ�}��J����?NW�?��?���>Aү���>ҩ���'p�Hm�=>�m">1��Z[��\�?Ng>�/�o�|�|���>�?%�@�`?Ps���ݿ��=�7>�^>%�R�t�0��A\�pc�SNY��W!?F�:��~˾��>�=ď޾wƾ�+=�5>b$`=~��5G\�y��=��z��I:=C�k='��>JkC>M>�=����ɵ=_�I=��=ݛP>iЮ��U7��O.�j1=l�=�Yb>U�%>u4�>�?$
0?Krc?縸>��m�ؿ;���ˑ�>Qf�=ke�>m^�=�D>�o�>�~7?��C?
2K?�S�>rg�=�>�B�>͆,�Gm��@律���Ɯ<�I�?ϑ�?�Թ>��w<�<B�3@��Y>��Ž��?�'1?в?���>�� ῔�"��l2�##���	�,z�<a�Q ���RB�,��E/ӽ��=O�>]��>���>�Mu>�@=>��S>*��>sw>o�G=���=� f;4=���i�=A�� !=
c�F���ڬ���o�ʀϼ!��;��;p�;؜��*��=z��>G�>֡�>}ؖ=D\����->Y̕�&�K����=y�����@�n�b�+k}�t�.�2�9���C>ϞV>=��Nܑ���?#A]>�A>��?��t?��>�G��RѾ�n���ld�CR�Lm�=��>}�?��<�.�b���O�
Ҿ���>M��>S�>>m>��+�A?���w=���SM5�3�>�Ҍ�����;(q��6���h�K�ֺvD?d@���F�=�~?ګI?ڏ?ܔ�>�)��\cؾL�0>Ǜ��b�= ���'p�O��l�?I�&?���>j�L�D���ƾ<����>,�G���_�AD��}3��Ƽ��о�>:؜����R25��.��l��t>�����rE�>�Y?��?V�׽�΃���A�E��&`�a7�>ݜV?�Ʌ>��>k�?�����)������=Nl?{��?�]�?H�>��=ۭ���>N
?~�?���?��r?��9�85�>���;|�>Y��<c�=��>:��=� �=�?
?Z�
?F�?H��[��~����m�b����<d�=�3�>9p�>�@m>���=Ip=��=�+\>yN�>�x�>��b>�%�>C+�>����3
��6'?���="�>�2?�&�>D�d=^���A�<SE�<��#�Xĸ�v��� �<���7�U=)����>�+ǿ��?�W`>�f��;?�����Z���X>;RW>�V�^��>��@>7y>!)�>,,�>&�>�Ӊ>�M">�<Ӿ��>{��#c!��$C�RR���Ѿ�mz>)�����%�����]���3I�mf���h�j��-��=9=�S��<�D�?T���\�k�s�)�Q����?�b�>�6?�׌������>1��>��>�@��{����ō��`��?m��?��b>"�>��I?
�?���z/��_f��a��P��a�~���*������=����I�vt�fW?�*u?��[?P��=��>�?�5_�F~�M1�>ɫE��:C�h&ؽ�~>%�绡��X��/Z��
GN=��?\ɜ?'�?��>���է.=!�=��>�?��?Cfx>
sI?Z��>1O?G
M>�Ѝ>Ф;?^�Y?<�?;�=���$s��,�>㣂>�Y�������K��G�N����~8��"�������R=�w�=�X�<�Z�����=���=���<��g=��=$L6=[�>�]?�c�>�׆>��7?���p`8�RB����.?[5=W͂�c^���������>�j?C��?�
Z?(�b>��A���B�|f>c�>�s&>_�[>��>����E����=<>��>�v�=/�O�d����	������}�<�>{K�> q}>UF����)>喣�n�s��&X>d�b�ֵ�̴_�lC�4c4�?^��ɞ�>�O?�x ?���=��R<��
d�i�'?l;?��L?2G|?��=��׾��5��J�0�����> =�
���3Q����8�J�_<]�>���������a> R�Լݾn���I��羘-K=v�o�T=���	־�B��O�=:
>ǉ��&� ����
㪿�IJ?"�j=}?���U������>���>{m�>��9�g�v�S�@��߬�\M�=���>��:>3i��,	�\zG�X@�w>�>PQE?7W_?k�?"��Zs�A�B�v���mc���ȼG�?qx�>"h?�B>P��=^�������d��G���>���>d��H�G��;���0��B�$���>W9?�>��?`�R?��
?��`?�*??E?'�>k������ B&?6��?��=��Խ�T�� 9�JF����>|�)?�B�ܹ�>P�?�?��&?�Q?�?��>� ��C@��>�Y�>��W��b��=�_>��J?ٚ�>s=Y?�ԃ?y�=>]�5��颾�֩��U�=�>��2?6#?O�?���>��>N�����=ٗ�>�c?~0�?�o?'J�=+�?|42>���>��=Ŧ�>'��>�?�TO?)�s?�J?���>��<H���-��q�s��P���;Z�G<(�y=���t��J���<�7�;�\���J��a��%�D��$��h��;�_�>��s>�
����0>��ľ�O����@>����P��7ڊ�>�:���=�>��?���>�X#�D��=��>�G�>����6(?W�??E";J�b���ھ�K���>	B?���=��l�����R�u���g=w�m?��^?��W��%����g?7�Z?Iv�J�>�Pc����P�Q����yM?+�>��j���>�N�?�xr?��#?KD+�}7��G���o�,M��֊�Z��>�����q����>�=?z�P>�>��=�g¾�����E�B�?/Ԋ?R��?m�v?߮�=�\w�mM�֨�����cv?r{*?u�ξ��Q?.%�;����ԅ��b��D���u2���J�:+��%0��)/�1r�������=z�)?��k?_Ut?QlV?,�޾�"b��A�I�n�]&�	����p�0�b�e���/�r�ؙ�K�о�þw
��d����T�@��?Kdd?Q���?i
Q�����0ɾ��3=�V��; {����=\8���{+=��}=����ң�\���K??��>j�>�w?29l�XZ]�76�
lD��]����=�>o>\Ѷ>R��;ǁ���(�9�Ѿ�
���ή6v>�xc?T�K?L�n?Cn��*1������!��/�yc��2�B>�k>V��>J�W�Ӝ�.:&�EY>�@�r�J���w��W�	�ޡ~=o�2?C(�>[��>
P�?�?[{	�`k���kx�]�1����<1�>4 i?�@�>��>cн�� �$�>��d?��>�A�>�bb�:#��D��=|�>�>�N�>���>Nr|>{�`��[��|��M���X02�Ϳ>Khk?鉾�X4�l�{>�E?�t�s�$=p�>/{����	��@ϾD��9v=>�W?��>�!> �ܾ�����}�a�]�O)?�K?�璾C�*��7~>�$"?u��>j,�>1�?n*�>�pþE�C�@�?��^?PBJ?�SA?WI�>m�=0���%=Ƚ�&�G�,=���>��Z>Dm=�~�=+���r\��v�r�D=�x�=�μZQ����<����_�J<���<��3>Xmۿ�BK�՘پ�
����>
��爾v���Td����a������Vx�i��_�&��V��7c�ܡ����l����?B=�?����.��2����������Z��>ߑq������ ���(���ྱ����c!���O�6&i�7�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���z¤<���?0�@�}A?~�(�x���V=��>ʎ	?�?>
V1�IJ�����S�>�;�?��?�cM=��W�:�	��~e?�<8�F�<$޻o%�=	;�=�O=���V�J>%S�>{��<OA�f7ܽi�4>�܅>wb"�X��`�^�H6�<^~]>[�ս�4��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�ޅ�=x6�%���{���&V�~��=[��>c�>��,������O��I��V��=Q��%ſrD"����� =�;��j���������Z��Y��ځe�_�˽�a�=b�>O)G>�>�7g>U�i>�xY?�c?�A�>E�.>�U��Oq��|ƾ��[<1�~�;\�WC����#�����Z��K־%t����Ȅ��7Ǿ� =���=%7R�k���8� �x�b�Y�F���.?kx$>J�ʾ��M���-<�pʾ࿪�aㄼ�᥽ -̾�1�"n�=͟?x�A?������V� ��V�t����W?�N����E묾��=�����=v$�>��=��� 3�a~S�ْ0?-K?@����-��Z�*>n��l�=Hl+?�?�KN<��>::%?�",�B&�coZ>a�1>�l�>���>�z
>'/��.�ٽ�V?pFT?P��0k�����>����[!y��d=��>��3�:�ּ�\>�K�<����Kq�&��b5�<�6Y?c[�>�+��y�Q��Pc��,'�;�!p?G��>#�>�g?�77?��۷��Q�v�u��=�U?�f?���='X	��Rʾ�;��w�3?�_?~�>�r���ξ�z"��"�i�?��l?�N#?c�����/�����V]/?��s?`'T��ʖ��|��Y)��k^�=��?��'?)�!����>ňp?Pp������װǿ��=��Ȣ?���?'��?��켱Ԛ�ĺ��>��>�K!�+����C8�|���zA>($6?av��ـ�G���<t0?�]?-�?���2V�Γ�=�ݕ�[�?��?w���B�g<���Zl��m���M�<ƫ={#�5"�c��m�7�X�ƾK�
�ଡ଼��2�����>�Y@�X�j'�>�H8� 6⿠RϿ���Xо�Tq���?��>�Ƚ�����j�UOu��G���H�¤�����>�>����o��3�{�A�;�2b��v�>g��M�>�R��"�����/{C<ᐑ>]�>���>lC��5��}l�?%����ο՛���R���X?�֞?Oڄ?% ?�jE<�rz���y������G?��r?�Y?y����^�/f7�&�j?�_��wU`��4�rHE��U>�"3?�B�>U�-�>�|=�>���>g>�#/�w�Ŀ�ٶ�<���Y��?��?�o� ��>p��?ts+?�i�8���[����*��+��<A?�2>���E�!�@0=�TҒ���
?P~0?&{�c.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>)�?�J�=*�>�_>������սM>�=�%���>�lX?���>c>����D��a}:�1RN��!���U�&8u>�Sn?�]?�@m>/n��4�����Z7����4��=�c����YϽ��=�A>7E>���w���?�o��ؿ�i��r'��44?x��>��?
��0�t�߻�x;_?�x�>�7��+��r%��"B�N��?zG�?+�?��׾�n̼�>�>$H�>��Խ�)����7>ٟB?s"��D��7�o��>���?�@�ծ?;i��X?	t���ć��yo�Yd�I���Ҩ>�Q>?W)뾿�Z>�
?�1'=�V���A���{�Gy�>A��?�K�?Ţ�>Q�Z?�v�dl>�[�C��ٮ>!sJ?eM'?�Z)>>[۾<w�>�� ?�u.��*����񾕙[?��@'"@�le?����qhֿ|���N��$���r��=F��=��2>��ٽ�^�=��7=%�8�	9��%��=\�>��d>�q>(O>Aa;>v�)>���9�!��q��O���`�C�������Z�%���Wv�=z��3������G?��3ý\y���Q��1&��=`�.}f=�j?�_L?F�N?5�?ѝ:=@�<M��]=���`��=⪴>��&?��R?�)?h_=ꐕ��\���y����*����>Y�>R��>L�>���>��Ｆ��>-�>i҇>�z���	�=��=��8�ֹ>L��>�#�>j��>�C<>��>Fϴ��1��j�h��
w�v̽1�?����S�J��1���9��Ӧ���h�=Hb.?|>���?пf����2H?%���y)��+���>}�0?�cW?�>!��r�T�3:>9����j�4`>�+ �{l���)��%Q>vl?��f>)u>��3��f8�P�P�xy��jV|>�36?�궾�A9���u�?�H�%_ݾ>MM>�Ⱦ>yD�lk�C���F���i��{=�z:?D�?�%��Lݰ�j�u�zB���RR>Z<\>�=�]�=+MM>tc�h�ƽH��.=I��=֯^>�e?�+>���=���>�P���P��:�>ldB>��+>�@?� %?���������9.���v>�V�>'�>�y>�vJ��F�=�K�>��a>�H�N����a�?���W>�|�C�_��"t�ýy=Pw���c�=�=�� �Yn=�x7&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿih�>Lx�~Z�������u�v�#=��>�8H?�V����O�>� w
?�?�^�ک����ȿ1|v����>V�?���?O�m��A���@�Q��>0��?�gY?�oi>�g۾	`Z����>޻@?�R?G�>�9���'�b�?�޶?ͯ�?��I>Tw�?d?s?�;�> �u��^/�WA��م��	�{=S}5;R0�>�>�,���pF�OÓ��l���j�r��7�b>�"=�7�>���RѶ=S抽D��n d��ڷ>Бq>q�I>H��>X?Մ�>M�>�=ԓ���I��)O��US??鵔?�8�J���c�9>�x�=F�վ|�?���>vj@��g��?4Y[?"��?�e?\u,>���ͦ���ſ(���z�=Wã>_�>]�?�
�
>ai��*%8�&�>�~�> �w�����@��m6K=��>th)?�.�>;#���	&?�� ?�8>TI�>�5��U���J����>���>ng?Y�z?v�?:����U+�fŏ�������Y���8>6��?6�?�Z�>3���JH��g ��]�\���;��?X�f?6B����?��?9V?܄O?#�^>��4��e��l�Z��>��!?H�:�A��M&���o~?�P?��>I7����ս5Kּ��������?�(\?wA&?ݜ�#,a���¾�8�<��"�(�U�J��;ÀD���>��>�����=�>�ְ=�Om�{F6���f<�j�=��>m�=�.7�]u��� @?�����ɾ��ؽg>c�q`�.�>�۰>�蒾��5?x��W󃿻ӧ��n��a.����?�T�?Q��?�D=��0��A?�BU?� ?�?���3�7����Mþ�p���1��쒵>VS|>��>V�e��ɰ������f�� �����C��>���>'I?B� ?��I>���>nb��e�'��K�X��\�1����8�Mk.�bo�k6��&w��n伄�¾��u�}q�>�I��\��>�
?p�e>��|>I��>YE���>��U>S��>�ѧ>�S>��+>JS�=�'2;KzȽ�KR?������'����^����2B?od?�1�>�i�׉�����΁?���?�s�?3@v>�h�[-+�tk?�:�>��r
?DQ:=ܐ�Ԁ�<JT��I��t4����Ӫ�>�P׽T :��M�llf��k
?g0?F��m�̾QO׽[s�U>ül��?vsD?�I��=�*)^�:����0:��P��E��m������Vi�FV������΄�g�+���t<bP?D�?�L��`�Eݍ�]k��'@���>�s�>��[>~�>�N�>�0���P���o����7�1�?y"�?��w>��Q?��;?e�F?�S?`[�>+�>���C��>�28�>���>dZ5?��2?˽.?�
?��?�2>����s����g�?ل?�'?��?Q�?y����a���%"�|Y���9� u�=����c�轆&��cw"=>��>�h?�D���8�����pk>�N7?��>D��>� ���4��k��<N-�>F�
?�"�>_ ���r�"d��4�>���?��p�=��)>�l�=����������=䐾����=�����;�u;)<�i�=;K�=<�m�k�6�G6�:��c;�F�<C�?y�?r-x>�҄>P�r�T������=%�4>Y<:>h�>~ξ-��zT���|d���O>���?t��?`'�==�=gq>蝛�����A������)��<X|?l$?|S?��?�u>?[�(?n>fT��ޓ�tǅ�\կ��j?v!,?��>�����ʾ��҉3�ɝ?f[?�<a����;)�Ɛ¾�Խұ>�[/�c/~����<D������-��3��?쿝?�A�L�6��x�ֿ���[��x�C?"�>Y�>}�>R�)�x�g�o%��1;>���>gR?�#�>��O?�<{?ɦ[?�gT>r�8�~1���ә�>E3���!>?@?��?�?yy?�t�>x�>�)��ྋT�����7�=Ⴞ[W=	Z>g��>�(�>M�>%��=�Ƚ�Z����>�a�=�b>P��>���>��>�w>&M�<�H?�	�=���ɜ0��=׾���Q8<R�P?6�?:��?�~��6A���Y�K,z�������?b�?P?5^���=�ы����5�R�� �>�U�>bK�>�
������Nw���a=1��>���N�z�V�y>�>
�4?t|4>��ǿ��q��Qh��x���><�w����d��/�N�g�-�=_֏��������|>E�bM���������� ��/w^��Q?�>=;�
>@>t�7�(�<W =ج�=Y��<��B=�2g��i8��#��=��^S^�Ӳ<�<A,`= �7��T�d�?I<?ޙ?9�d?�7�>Cu�>�D�*��>�q(�{��>h�?>�͔<戏��,������S��w�Ҿ
���z ��QȾ��>�:�|�<N��=,�.>���u��zUܼC��=�/y=�0��Ay�;�>���=e�>�6>��5>v6w?����8����3Q�Li罆�:?J?�>��=~ƾ�@?��>>�3��Ǘ��,e��)?���?�T�?��?�vi�da�>����玽#f�=����;2>��= �2�h��>��J>Ѓ��I���y��I5�?M�@��??�ߋ��Ͽ}\/>5�8>�e>,�R��X1��[�A?c��S\�';!?f;�x�̾��>�{�=�߾Y�ƾmg,=�5>T�a=�����[����=6 w��;=x�m=0B�>OD>o��=26���'�=�BL=U��=jP>/]���5�7.�'n-=�=�)a>@}&>z��>x�?�a0?�Xd?Q6�>�n�Ͼ|?��VI�>��=(F�>M�=�rB>��>e�7?��D?��K?'��>d��=	�>��>Z�,�&�m�wm徚̧��<���?�Ά?AҸ>�Q<�A����g>�t/Ž�v?RS1?�k?��>�$��ؿ�r�RZ&��ca����;�<O<�����b罷�b��sQ���>#:�>P��>�]�>t0W>�Qg>��}>�|�>���=�ZO=��>�����w�=�dS<X��=�����-B=j弳�.�H�ۼ�_�â=�==�L<M��=]��<,/.>�v�>e��=��>���=�OƾΝ�=x�����R�Y'=	��tq4��k�A�{��>)���K��=>��|>C��X�o�?�yU>��h>�4�?�q?��=sN%�#�ʾEi����o����2̺=+��=��5�hqJ�U�b���R�����7��>�ގ>���>ôl>,�&$?��dw=���d5�w�>z��7��<A��9q��=�������i�u˺��D?&E�����=0~?�I?i�?U��>�@��w�ؾW;0>�B����=j�xq��e�� �?.'?=��>O쾫�D�br��ؠ����>�����X�v���.�~d����x-Y>󝾠���k4�3��������4�gv�F��>�DZ?�?s��#ԑ�n���ľ�S�[h?�P�?�F�>��?ٙ#?���$�0D���/�<|?���?M[�?CC>��=y宽��>gA?���?]��?��t?��D�M��>Z�';͕!>Yi��4?�=�b>�%�=�0�=#Q?�	? �?� ��*�	��X�t �۱`����<g�=Ls�>ʹ�>�4s>c��=Rm�=�ì=�p[>7v�>���>�Xc>��>��>?���(��� ?y�c>��>ѼE?�}W>P0���X��M=,�E=g�-���l=`ռ�'>��I=����
>,�T=y�?Lȿ?��?D/�>u-�;[R?^,���H>��>�UX>��@t�>_C�>~_>u�=�#�>�h=��
>�1�=�3Ӿ@>A��=>!��:C��tR���Ѿ �y>˒��F-&��������I�^l��f�j��.���A=��<iN�?���;�k�2�)��
���q?�3�>�6?�Ќ�?)���>O��>���>�e��ȑ��č��Wᾩ�?h��?�;c>��>9�W?�?ϒ1�V3�	vZ�(�u�r(A�,e�K�`��፿�����
�����_?�x?3yA?�S�<:z>T��?��%�Gӏ��)�>�/�,';��?<=k+�>*��.�`�g�Ӿ��þ�7��HF>w�o?2%�?gY?.TV�V˄�x?�>�"?:�>IK�?(2?�j?����1�>>c�<���>��?3?��?1 ?���= ��<&W����~>���P���`���q�j�2�~�ý�N=�S���p����=;��<��=���=*a0��)�<����� <��=���=
�>9�]?��>ۋ�>��7?�.�@�8�Jۮ�+�.? i8=j����������3�Ѻ>��j?��?LZZ?J�d>B�|�B�e>,`�>��&>�2\>�A�>��K;E�bd�=�J>��>���=ŦL��ځ���	�����!��<R>2��>,*|>~��7�'>�e��"wz�$d>q�Q��񺾎.T�	�G���1���v��&�>��K?��?^��=[�w���	>f��A)?�R<?�SM?��?삔=�ܾ?�9�>�J�b!���>�{�<J���������'�:�\�Z:tHs>������<n]>_��umվ�7p��bF�� �c�$=�K��19=,�YGԾ�@v����=oL>s�����!�Œ���L����J?h�^=j/����P���y�>�>���>��F�P�����?���,��=���>}4>y�����=�G��~��=�>�PE?pW_?�j�?�!��1s���B������d��sȼ �?�x�>fh?)B>���=����\�b�d�G���>���>���(�G�k;��/����$�y��>�8?8�>�?Y�R?i�
?b�`?�*?�D?@&�>c��G����A&?8��?��=��Խ��T�{ 9�IF����>y�)?�B�ٹ�>P�?�?��&?�Q?�?x�>� ��C@����>{Y�>��W��b��4�_>��J?䚳>s=Y?�ԃ?o�=>X�5��颾}֩��U�=�>��2? 6#?N�?���>|��> ����r=�q�>��b?��?��o?6��=^�?��1>�!�>駗=yݞ>ke�>^�?@<O?q�s?K K?(W�>K�<�j��U��F0r��U��g|;��F<{�z=:)���t��5�C��<֧�;@���ʈ�R񼗁F��c��3*�;�`�>��s>j����0>#�ľ�O����@>u���Q��Tۊ���:��=��>��?���>�W#���=g��>G�>)��86(?��?�?��!;��b�s�ھӮK���>uB?���=*�l�������u�V�g=�m?U�^?��W��$��u�f?��\?���>G��W|��J��Ƣ�Ro?Nc?}������=�*�?��t?�P?�Tƾ�슿�4���sp��Sݽ�/���?ѣ���`����>�YB?��>�17>��۽�wN��bs��n"?o	�?n��?�ف?���=��c�ۚ�5=�-����T?��>�2��D�'?�ҽ�������Z��'l��
��ډ���x���,��V˒�_�W�o���sƽ5�=K)?mr?�>�?0zz?[@,���E�_v\��v��DD�AY��(�#�?���6�B�7�H�_�?��H)�����6��@���Z6��e�?C\m?��r?R�꾁'�Lv��&-�����Խ��b>��<��<��=�� ׾�Ӿ�y�q�D?���>�6?uA?��l���#$��#�����A+;�t+>��\>���>57l=¼��#�X�.ϣ���Ⱦ7�l��6v>�yc?��K?�n?eh�*1�Ɔ����!�ֲ/��b����B>�m>庉>T�W����9&��X>�y�r�Q���w����	��~=��2?C(�>���>�O�??vz	�j��hx���1�<��<�-�>w i?�@�>��>#�Ͻ�� ����>��l?u��>��>�pZ!���{��ʽM&�>
�>��>��o>6�,��#\��j��V����9��u�=/�h?���,�`�I�>~R?�%�:i�G<�|�>N�v��!����
�'�=�>l|?ɖ�=x�;>3�ž�$���{��7��+a)?��?������*�vz>� ?A��>�=�>S
�?��>�Ǿb<�/�?}�\?�zJ?�B?5�>�=;���`_Ƚ�%��t.=���>� X>��g=n�=�����]�3��	<?=�=���������&<�q���6<���<��3>�-ۿJnK�n
ؾ\���:K�F~���3��cT���;��q���=��}8t����Y"��X���f�����3i�C)�?o��?�1���ǃ��8���\�� �&q�>�n���|����{r�T������o����!�eP���h��e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@#�A?��(���쾞�U=%��>Qn	?k�?>�1�V�U���^��>�*�?ӊ?@�M=�W����"�e?H<?�F�N�ۻIj�=�Ƥ=	�=��]�J>���>e���|A�o�ݽ_5><N�>J�%��x��$_�'#�<�]>�սx�b�?:�^��vX��3��y�|\�<�]l?s�?���>�Y?�*_��)ؿ�:�#�0?��?A��?j!A?�r�����>E˾Sd??[�)?��>���ԭ^�z�=��7�N�<��Ⱦ��R�,ޣ=�)�>
@d>D �����S�M���A�=P� ��Cÿ�6�b%�$"�<�J=_{���� �RI��/{<��҆��_M�����œ=�G�=��0>��a>�4U>2+d>�Y?��i?zi�>��a>v$��l��0ؾ']���P�~�m냾��K������Y�ھ��
���W�Ly��!=�z�=7R�r���/� �Z�b�]�F���.?�v$>l�ʾ��M�2�-<_pʾ;���j܄�a᥽�-̾�1�,"n�_͟?��A?������V�@���X�����T�W?aP�˻�ꬾ��=�����=%%�>n��=|��� 3��~S�$|2?��? Nž���(>�����=��*?R�>�:ٴ>��$?�)N������M>��8>�G�>���>v�>`ԭ�(޽�?l�R?}X�k���y�>����jh�١U=��>$'$���D��dG>l׀�����ȼ%&��>�=�,f?��G>��0�v�i�h�m����m ��lT?�0�>��z>�V�?0;?Q�����u�t�����R�=��??Jj?�H>�vU>-Tξ�Y��g�I?��e?���<C�����8�Z��2��.[?!,V?`�G?��/�p��������!?�bt?�[�2̜��S�_���9@<�	?��?Ȟ>�ԑ�>�zM?e���k��lο�0:��:�?��@�?Q�<[�W��^����?b!�>]����ݢ��J5>����#�S>19?X8��� ��۸þ�85��sO?N��?h?s���3���|��=�ٕ��Z�?��?����Ig<[���l��n���}�<lΫ=��2E"������7���ƾ��
�3����㿼�>;Z@V�k*�>�C8�U6�
TϿ$���[о]Sq�z�?D��>t�Ƚ����I�j��Pu�S�G��H�����6O�>8�>�������� �{�kr;�A䞼�>���/�>i�S��*������5<�>@��>��>� ���彾�ę?�a���>οZ���4��V�X?gg�?Kn�?�q?ͦ9<&�v��{��F�>/G?0�s?`Z?�t%��A]���7�*�j?�_��{U`�ڎ4�`HE��U>�"3?�B�>[�-�F�|=W>���>!f>�#/�n�Ŀwٶ�����Z��?щ�?�o����>d��?js+?�i�8���[����*��Y+��<A?2>׌��O�!�G0=��Ғ���
?/~0?={�F.�Z�_?<�a���p���-��ƽ	ڡ>վ0�~a\��"��'���Xe�_���?y���?�]�?��?���| #��6%?��>ٝ��8Ǿ*
�<΀�>�(�>*N>C_�b�u>�E�:��g	>u��?�~�?6j?��������S>��}?���>9`�?#��=ϫ�>��$>�;��xc��r'>0��=�)a�� �>�M?���>lX>Ⱥ���+�T�D�]�P���G�D�B|�>��h?�~R?j�w>������P��XQv�ӯ�]��<�DK��-�����]�T>7TP>��4>���l�ƾ)�?�o�ؖؿti���q'�D44?���>��?���ߵt����;_?�w�>�7� ,���%��A�v��?�G�?G�?�׾�̼�>�>�F�>��Խ�퟽�����7>��B?�!�E��,�o��>��??�@9֮?mi�??U��������j����������=56"?ͱ�=�B>���>WN�<P��u����x�;��>�ۮ?bQ�?{?�Z?��p�-�J��H��V+�>�~6?
�?�=p>~��OB�>��?%;��)��0��:_?��
@T@�+f?�9���Կ��F����`��>c�c=��->� f�NR���~��hj�=K�<�S:>��>��>�>?�>U�>�����|�/�#���ʹ��iH��K(�4�����]���4?��F�5Z���;��J�*�k����01��]7�E�5�G$����=rt?�r??[�??�� ?/9���|���]޾�m=���8��<��>�?�M?
#5?�1�<�]��ҝM�}.��f���u����>�\�>t�>�%	?��>��=!�h>?�6>��>bL�=D�v=���Ad>�]>a��>C)�>{5�>�C<>��>Fϴ��1��j�h��
w�u̽1�?����S�J��1���9��Ӧ���h�=Hb.?|>���?пf����2H?%���y)��+���>|�0?�cW?�>!��s�T�5:>9����j�6`>�+ �{l���)��%Q>vl?��f>B,u>��3��f8�C�P��{���V|>�06?'궾�F9���u�`�H��_ݾ�TM>�ľ>pD�Zl�������Vi���{=�z:?ކ?V���᰾!�u��A��;VR>�@\>�=4]�=#JM>�_c�d�ƽ. H�*�.=���=��^>�?d"*>埄=�J�>������P�?F�>��C>7�&>܅>?&?������I����/��ax>���>�w�>g%>PSJ�f��=
t�> �b>s��o��99�9<��xZ>�}��Z�Ňe��d=���1��=!i�=k\���=��/=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾQh�>zx��Z�������u�t�#=Q��>�8H?�V����O�e>��v
?�?�^�੤���ȿ5|v����>X�?���?g�m��A���@����>;��?�gY?qoi>�g۾=`Z����>һ@?�R?�>�9���'���?�޶?֯�?aI>���?�s?�k�>�0x��Z/��6������p=��[;�d�>�W>e���wgF��ד��h��u�j������a>��$=,�>QE�[4���9�=��I����f�;��>�,q>�I>W�>v� ?�a�>~��>�x=�n��Jှ�����B?��?gZ#��%����!>yo=e��aP�>�L?�ɽ�)�����>:'R?�m�?��>?5�>�:����@�����f	>��>��>�(?5(��k*>�֫�h)�ā�>���>����r$�d1��&/>���>t�*?6��>.��� � ?��#?�nj>~�>ZE�S9��]�E�]��>���>F@?e�~?T?�乾*R3�U��%塿��[�1N>�y?iP?�ە>��������ęC�ֶH��q��퐂?Tsg?��P�?�1�?)�??ϨA?�f>����&ؾ�����>}�!?�K���A��M&�7#�a?c?��>����Խ�ټ��'f����?1#\?�V&?3t��a�E�¾���<�"��*S�V��;�yE���>��>�W�����=p�>��=y-m�)%6��9i<Q�=#r�>��=�C7��:����,?ʄ�$�����=�r��&E�΂>�rS>����_?)C8�X�{�PX��}���]T�$�?�N�?=7�?�]���xf�\!=?��?�?���>_$��S��"��v��i~�����r>eY�>�+�����P��I/���J����Ž���g��>��>n�?q� ?�qP>ᄲ>E��At'��N��=��2^�����7�Zh.�<��h
���}"�s=�ç���l|�p�>����>��
?i�h>�z>�>�ʰ��>DLS>�>ͻ�>��X>�4>� >
�<�ѽ�KR?����0�'����)����1B?0gd?+*�>z3i�������<�?���?�r�?W/v>f�h��/+��d?�0�>���Ju
?�t:=��8щ<�Y��4��8��a]���>)@׽m:�YM��]f�xo
?�4?Ź���̾Dz׽C�c�UC@�w�?��`?ԇQ���m*o�@Qz�K D���ݽ�M���#}�5��4N�9�����J��Rn>��B=�/F?O�z?�&2��O
���Cȅ��� ��*>�˲>�T�>Z�>��=6��\�g��!s��G#�@�p�'?��?vǋ>��J?��;?�xN?�M?���>�i�>�e�����>�;�J�>׎�>(�8?��-??�0?J�?d*?h�a>Ab�F��fؾЩ?��?y?�;?��?e!��X���������U��Qx�}z�1pw=���<�ӽ��r��X=�U>"q?�5�8�]���A�j>�T7?}[�>ÿ�>�c���N���~�<��>VT
?�B�>���kKr�l%�{��>��?����=?�)>���=�-��Dú���=�>���ѐ=�2���I9��8,<&<�=��=N+��;e���>�:�y�;e��<�n?d?��M>Ñ�>u߃�f��m: ��5>��5>�9>ݵ�>ｾ�`��WK���ln����>$�?�m�?Ge�=�^�=�D�=�c��⓳��{���Ͼ%6|��7?o2?P?���?�A?�W?$��=�X+������'��n��z�?w!,?
��>�����ʾ��։3�ڝ?i[?�<a����;)�ݐ¾��ԽԱ>�[/�h/~����>D�h���S��6��?�?DA�W�6��x�ڿ���[��{�C?"�>Y�>��>U�)�}�g�r%��1;>���>kR?t �>��O?f;{?Ң[?tT>o�8�0��'ҙ���3��!>0@?���?��?�y?�w�>m�>׸)���
Y��^��K�܂��W=�Z>Ø�>',�>M�>��=��ǽ�S����>�Rh�=��b>5��>֟�>���>�w>�y�<"K?_r,>0Ҽ�""�ݖ׾�\�����>���?f�?� ~?�l���h�������[�>�j�?�|�?�.?ⷸ<ۘ>Q6�=0͟�����@�>��>��=�V�-U@������?�?H��nK��j�3�,Q�E��>� 7?SJ��rNƿ�q���m�����u_R<�8���g�?��Þa����=fn���X��n����N�<����5��p���-���w�� ?�=">z�=��<��Yx�;��(=y��<�	2=�y^�`!=<ՌB��W�������ҥ<�!I=6���O˾Lʀ?�XD??'L?�L�>��>ǈ����>b,��+?�lp>�4�_X���⩽���_/��y�����O$Z�뿪��>�Rc�Ɩ>i}>C�B>BN�<M!�=�G=�s�=�<2)S=�:�=Pþ=`��=?=�=�>:>Ӹs?2��̰���V�+�Z��O�>o��>EG}>ִ��ٞg?��>� �������9�)�s?���?l��?�?�d�̌>Dښ�j����4�=�;�G�>��8>��d���?�ѩ>� >��A��L�=���?��?��:?�tz�5�οo�i>wB�>�)�=9W�D�#��{;���h���?�"�?��E��i׾
-�>B��=���N���c�;��=>f�>��ǼDwH� ?z=r�r�X�={��=̞b>�C6>��q=�D���=����s*->%Ő>4���IŽn�)��+%=)�L=lxI>�57>���>Q�?\a0?MXd?<6�>�n��Ͼ?���H�>�=�F�>E�=\pB>֏�>�7?y�D?��K?���>��=,	�>��>#�,�Ҵm��m徨̧����<���?�Ά?Ҹ>��Q</�A����g>��2Ž�v?�R1?�k?��>
����οX%�4|�{t��A->G������؎�����Z0;��p�N�>��>3�>^�I>��{=�F�=7�)>�4�>;�>sŐ=Q#>�E��4׵=uq���0� ��=��{=�=
���;�4=�s�a{B�'���¸:��(�=[%�=N�=0��>
>���>��=R��O/>����z�L���=���>$B�?-d��8~���.��+6��B>�sX>�~���(��!�?M�Y>�?>@��?CEu?�p>ej�R�վ�[��[�d�#�R�X��=D	>�1=�
�;��U`�X�M�ZvҾr��>^ߎ>��>J�l>�,�E#?���w=��Ob5�b�>�|��Կ�)��9q�&@�����vi�uwҺ��D?�F�����=c"~?�I?`�?���>g��܆ؾ;0>�H��x�=l�;*q��h����?'?��>�쾲�D�+�����ӽ���>!����hT�@�����&����Yվ�>����ƾ�?8�X���D����)>�3E`�+�>7.q?�? q�՘��p�����7z��-*?T�?X)P>���>��?cl,��!���澷��=ځ?��?�X�?#�>#�=�ۯ��P�>��?Yu�?응?��r?�+A�s�>]�V;F�#>�G����=S,> '�=L��=K}?��	?�?�����
��H�N�l�[���=4��=L��>�f�>��s>?y�=�v�=q�=��`>��>A�>��]>��>��>�O��e���h'?@3�=�b�>��3?ǀ�>�8/=5�i�<{��k+��}��c����ƽ���;߀<�\Z=�D[�%��>&ſ8�?��<>����?��辄�?�:�?>H�Z>���Y�>��L>�u�>a��>A�>4\>���>Q�&>�5Ӿ�C>0���1!��<C��bR���Ѿ'�y>8���`0&�8���T��aI�U��,l��j��.��}M=��*�<J�?����A�k���)�>}��qs?�d�>N6?�ό�������>���>���>gq�����qǍ��M���?P��?�<c>��>��W?�?��1�L3��uZ�7�u��(A�e�9�`�j፿���N�
��
����_?��x?jyA?we�<�:z>0��?��%�[ԏ��*�>;/��&;��J<=�*�>�)��9�`�ޯӾ��þ:�cIF>�o?�%�?�Y?�TV��}e���?�L0?}}	?k#�?��G?VI"?��<�@?�"��L�>�e�>U?�u?}V;?Q�u��$[�"���D��{� ���Ǿ�����?׼��޽=o8��HY>Gy��u�#�9<��=E����?���{��w�<�a9�<���<.H>֦>�]?��>��>ʽ7?���d8�m����	/?C9=�q��?�������N�>��j?���?�iZ?+Hd>�A�IC��>W�>�2&>�[>�T�>2��UE�y�=u>S�>c/�=w8N����Z�	�U���a�<�>>D�>?{>���ʝ&>���]{�Ue>��P�,����\R��ZG���1��0v����>n�K?��?yk�=�Q辟����e��Z)?�;?YM?��?���='Cݾ�S:�� K���=��>�6�<0N	�
.��)���;�Yˡ97bt>�Q������E,>T ��; �h�ǱA�:�ʾ���;�����=t�c.Ӿ�vN�K�>�Y#>���H�w@������yrJ?jR=��o��1�Ǿ��M>eL�>��>Ah���x���:�ҽ���=$W�>ƫ!>�
���$E�q2� >�>QE?{W_?%k�?�"��s���B������c��vȼ��?�w�>h?�B>��=�������d��G���>N��>1��-�G�<��@0���$�L��>9?ǫ>%�?[�R?^�
?3�`?�*?;E?�&�>��������A&?;��?
�=��Խ��T�f 9�<F����>{�)?%�B�˹�>L�?޽?��&?�Q?�?^�>� ��C@����>^Y�>��W��b��'�_>��J?��>}=Y?�ԃ?>�=>R�5��颾f֩�U�=�>r�2? 6#?F�?���>X-�>�h��A�=��>Z�b?t�?�p?g�=Z�?Y�8>%��>E�=�Ɵ>[�>r�?'FO?��r?s`J?Â�>�t�<
��������z�D�U���<�S<s/w=�����j�� �P�<uд;�𱼹Q��e缷�B�ͷ���B�;,_�>��s>v
��Y�0>.�ľhO����@>�|���N��,ڊ�+�:�T޷=Q��>J�?��>(Y#���=鮼>�H�>��%6(?%�?O?�";�b�?�ھ��K�i�>j	B?	��=`�l������u�>h=��m?�^?�W�%���n?r0A? x��CP�����+����2�*?%R%?�U��Q} �1�s?2@�?��?Ԭ��6������a,f�]dӽk�<(��>�[��^�%T�>.U?yi>��?>M�=)�����* ľ^�*?X=�?X�?�r�?Kj>��L����O	��k����d?�?
վ�1?1V>W�־6yѾWtѾ`Z��Y���B���?������<�����v�?U�=�2?Q4f?�S�?J��?pH�iV-�$k�SH��j/�,/F��-$��Z[��C��=�p�����A���s�Ӆc���p�K ?��c�?�? T�)A?�Us�.�j��N6�0E߾�־����=��缘����>0�����¾��DMD?WG�>��>��#?�T��,�H��p=P�GǾ�f�>��=_�>���>��� �$���0�i�ž'�`�e86�:7v><yc?F�K?6�n?m�W*1�������!�-�/�/c����B>�j>8��>ЮW����9&�qY>��r�!��Rw��G�	���~=�2?D(�>;��>+P�?J?F{	��k��kx��1����<l0�>5 i?@@�>�>(н|� ����>��l?��>��>ǖ��wZ!���{��ʽk&�>�߭>��>�o>��,��#\��j��J���r9��v�="�h?냄�v�`��>8R?��:��G<R|�>�v�̻!�B��<�'���>G|?g��=��;>)�ž�$���{�k7��Z�(?Z�?w���*�@�>��"?T�>�3�>��?�4�>�þ�8Mh?-9^?l�J?�v@?�"�>yM=�쭽�ʽ�
)��*=�7�>|RY>d�o={��=%|���Y��!��]H=p�=	-ȼ�_��a��;װʼ��_<�=�<�5>�lۿVCK��پ<
���}>
��䈾�����e��(���_����Sx�����&��V�@8c�⤌��l�C��?�<�?�~��9,��&���ԓ������k��>�q�Ś���X��i)����������c!���O��%i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >YC�<	-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾x1�<��?7�-?��>Ďr�1�ɿc���{¤<���?0�@��A?d�(����FX=3��>�9	?q�?>q�/���)S��,{�>/�?�Ǌ?�[I=W�����e?��<��F��%�b��=]b�=�<=Q����J>|��>4���@���޽7R3>�t�>;_%�����]�'ò<�']>y�ؽ����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=���ڕƿxf$�=0��� =y���-�U����>����I�l����m��T�F�p=H��=`qS>z�>v�S>��V>YOW?[�j?���>�>��彷Ԇ���̾���E���]� ���g������E��N�߾!��Ѥ���xȾ!=�u�=�6R�T��� � �D�b�,�F���.?�v$>&�ʾc�M��-</pʾ%����ׄ�kॽ�-̾ �1�"n�U͟?v�A?������V�C��jT�p���.�W?�O�����ꬾâ�=#�����=�$�>���=���� 3�K~S�T�1?I�?Yҿ�ꌾn�)>��	�0=1�-?��?ɭ�;v>�>�k%?{2����3V>�+/>���>B��>��>���m׽{?"�Q?ik��b��w͊>B���nav�-=
��=��$��4���K>w��<���h�r٫�iy�<t�n?�о=5�>�e�˾5�~��<Ѿ,���A�?�#?c�N=l�[?�j?�C��O]#��f�E��0ü>�n:?b*s?�&�=��<�DԾVϨ��?Z`U?�M��㾋v����#�߰-?�#d?ل ?q2�����瘿vi'�sh'?�jv?��T�����u)��LP��vb>x��>'��>��L�%V�>�N9?@��Qţ�<�ʿgB��Ī?�@S��?1�妻��Խ��>d��>��8� Q�f���A��C>�s?
%��Oh���ｏn?J�w?ʆ?Qڢ�ͤ����=�ە��[�?(�?�����g<w���l�q���<M��=@��>"�\��y�7�h�ƾ��
�ﮜ��-��3��>uY@iO�,*�>�J8�!5�<SϿi���Xо�Pq�#�?���>�ȽU�����j��Pu���G�y�H�w���I�>��>����������{�[p;�䞼��>�+���>��S��&��ʗ����5<��>���>��>_4���罾�ę?�c��t=οK��������X?�g�?:n�?�n?f9<,�v�ט{����V,G?�s? Z?�w%�5<]���7���j?zo���g`�z�4�n3E�:T>��2?�@�>�5-���~=��>�!�>N>;/�8�ĿM����b�����?��?�?꾃��>w�?Kt+?�5��	��}� �*��;�8ZTA?qc2>y%��y�!�T�<�*w����
?�0?��?"�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�ʶ>��?���=Z��>N�>���{�Ƽ��!>Q��=��3�s� ?�2M?��><��=��,�f�,��E�z�Q������D�s�>��b?��M??l>w����1�0� ���ý��/��Ł�� @���,�
�Y 3>�^=>إ>��>�!̾�!?���Qt׿HQ��h�*�;v)?�tn>g:?M��\��s<~V?�e>"��T����҈������?x!�?�d?.rҾ���o>i9�>��>w����V��rq�=�P>/B?�
��b����[a�)A�>���?�R@��?��e�uI?�x�b"����f�=k�o]��pr�=k�&?�����1>b��>�Ǵ�EV��v����y�n;�>Uܰ?�q�?1��>�+_?�z���N��⢽N[�>i�.?VX?{�9>ŷپtv�>�4'?���c����Q��G?�@�@U�k?�h��JTϿ�퓿}x�����ul =JF���ɇ>3S�����q�9=,^>��2>�Qk>ժ�>D��>yE>�O<>(F>>�c =I�~��S!��홿��F��B�C7�>j����徭�Y���ƾ�wM�^��B�en�&�ƈ�!^E������=Y�|?�QC?x2R?�)?�?�=�G���ؾ�z2=�kɽ�nּ�!�>�|%?{�H?�EA?q��=�S��<T���m��;Bx���`�>���>Sw�>(��>�2�>�d�=��> �=fP�>��=��=�����D]<a�>���><5�>��>�B<>�>/ϴ��1��T�h��
w�=̽�?����%�J��1���9�������i�=Ob.?�|>���?п_����2H?4���^)�.�+���>��0?�cW?r�>*��3�T�:>����j�	`>�+ �Ml���)�T%Q>�l?��f>�%u>�3��d8���P��t���\|>�06?�궾b=9�x�u�îH��]ݾ#SM>Hʾ>��C�uk�����t�V|i�Ю{=�y:?ԇ?s���ݰ��u�zC��&KR>x7\>B�=�_�=�RM>�c��ƽ�H�4`.=���=ƹ^>��?!�>K�s=��>O���K�ޡ�>���>��`>r�@?	4?SB��uԽ��e���P�d��>>��>���>TI4>w�E���>p;�>�lt>O�R��~C�,?�3r2�dz >�|��NTt�d�����=1�kI>%<PR۽\SQ�䮔;�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ*p�>~{��Z��2���u��b#=���>�6H?6G����O���=�u
?�
?�^������ȿ�wv�`��>��?��?��m�O>���@���>���?cY?)Yi>[۾�RZ�q�>��@?r
R?�*�>�4�]�'���?jݶ?���?AI>���?�s?�k�>]0x��Z/��6�������p=�[;�d�>�W>Y���sgF��ד��h��m�j������a>��$=�>E�k4��9�=��I��1�f���>B-q>�I> W�>u� ?�a�>���>ty=�n��Mှ������H?p�?D�%�w��j">O��>�YӾ�v�>�?й��}4���>g�S?��?�8n?�$N>����𔿥�ſq� �`q�>r�>�?�(.?�G��e;�=��Ҿ�ẾL�>���>2-�<�y�d���L>��>��?�n�>\��=�� ?m#?_�i>�>�OE��A���F�ܻ�>���>?~�~?m�?@C��`]3�����֡��\[�~�N>L)y???�ѕ>Dt��d��!�=�nDF����*z�?(�g?-�㽏�?B2�?�y??��A?�Kf>��u�׾����K�>��!?��A��M&���j~? Q?;��>P5����ս�Jּ9��Y~��a�?�(\?�@&?Ɯ�=+a���¾�7�<��"�rqU�N��;��D�&�>��>���Ɖ�=�>pװ=�Mm�}E6��f<0m�=6��>>�=�-7��t��T�2?!B��="��ui=�tr���Y����>���>i����_?�e���v���M���
���3��8�? ��?���?IO����S���%?��}?a�?1H�>uٰ�M0���㾾�B���b�����K6u>���>�C=���P���!9��⯌������N��>���>�K?B� ?�N>���>�m��y>&��j��2� O^�����28��.����Ӡ���!�����k���}�έ�>�����>�;
?��e>{z>���>�����>��R>��>�>��X>�7>��>|	<_�Ͻ^R?(@����'��h��Q���cB?U�c?�<�>��a��o���V��b?&��?F��?(vv>�dh��-+�q�?  �>Q\��K�
?U1;=]��#��<%���f���`����>	O׽W:�M�,e��.?�Y?3i���V̾��ܽ�I�!k�:�b�?:�[?��U���#��
>�Kxu�
Y��;Q���ž'ξ�I�+;\��m��-l��K����]*���;�'=?.R�?�C��o�{���k��N6�NI�>g��>j�h>ߊ�>���=kV-�N��0c��7��@�ʏ+?��?f+�>�P?��:?�gK?p8R?嘚>���>G�����>�	<�"�>8��>{�6?��,?�\4?%?��"?^tS>1����~qھ�?]�?�?"[ ?3h?�_d�( ��'��k_��u��n�c�9=�	�< D�8Y�3�e=��g>�c?���b�8�������j>�<7?&�>[��>���_3���U�<���>�q
?4�>�$ ��nr��C�Fl�>԰�?�����=��)>
�=䭃�*{��g��=��ü���=�p{��L;�ؼ&<1��=ʌ�=
�f�i�n86��:؞�;��<��?�?jrs>��>����Y��م����=�em>҉%>u{">�ڿ�7���.��2�b���Y>X��?�}�?�D�=��=U�=�u���@þ8|�	����&<W�>�2'?'qO?O�?��;??��>�������I��%����?w!,?��>�����ʾ��ω3�ѝ?g[?�<a����;)�֐¾��Խ�>�[/�d/~����<D�����2��5��?�?�A�S�6��x�ڿ���[��y�C?"�>Y�>��>U�)�z�g�n%��1;>���>mR?" �>n�O?�:{?�[?��T>��8�S0��*Й���2���!>�@?��?���?ty?0�>�>��)��ྟN��:	�	$��ڂ� �V=�Z>���>h;�>���>���=xȽ�C����>��`�=�yb>���>Ɩ�>]��>^�w>d��<�W?ج�>�̾�H�꓾�˾�G��4|�?=�?.C<?��>T�M�_�a���C�=�!�?tO�?#�a?j8=Y��=(�f=L����/�t�>�˱>���>�|�>��<Lp>�R�>؍�>��P=Y����.�fՁ=8?F??���Suſ�x�u\�.���~ <����+�������Zw� N>��'���-:$W2��ٽm�&�0�R�{����0�����>P�W=Ӫ�=��=o$B=,~�=M�=��W=�S=ߕ=;�y�Q`ս4�L�� ʻ�$�x>=�F;?�ż�pX<�˾���?1�;?+-?�wL?9=�>��>�?�<��>�
��D?�8>�gg�m����Žp�¾�~������t���F�_�殾���=�^���:�_=7ڮ=�i;�'XT=L�=���=�`���?=FZ�=��O=���=Ƌ�=ۭ>K  >�6w?W�������4Q��Z罙�:?�8�>�{�=��ƾs@?��>>�2�������b��-?���?�T�?F�?Dti��d�>[���㎽�q�=A����=2>p��=W�2�c��>��J>���K��8����4�?��@��??�ዿТϿ5a/>M8>��>��R�zn1�5�\�Y(c�ԲZ�	�!?�
;�W̾P�>�M�=xZ߾��ƾ��,=~*6>&�d=[���\���=� {��H;=��k=>��>ID><"�=P���Tķ=�8J=�A�=�0P>�֘�kl6�Ը+�k�3=|�=�}b>�	&>���>��?Aa0?;Wd?9�>n��Ͼ<���I�>0�=�D�>t�=�qB>��>��7?f�D?��K?[��>�=w�>��>��,���m��l�zʧ�֬<���?EΆ?�θ>'�Q<��A����g>��0Ž�t?�R1?�j?:�>g���2Y���i��#�Kf;�����CY���� y�ý>1=$�>v'�>��>���>Q0�>�S>4��<��_��Ǭ>�3�=��-=g�3>���%�(��=1X�<���]�Q;�qk�(B�A�G=�uO=���<6��=(�*=��U�ڼ���=e��>y5>`��>��=H��N/>ᦖ���L����=�8��'B�!2d��F~��/�/O6���B>�XX>>b���1����?�Y>�i?>8��?�>u?�>n0���վ�S���_e�1S����=Ѝ>��<�@�;��U`���M�$}Ҿ���>Fގ>��>k�l>�,��#?��w=���`5�R�>�{������,�e9q�N@������i���кġD?0F��:��="~?��I?,�?ڎ�>���<�ؾ�=0>
G���=r�(q�^����?e'?��>��8�D��E��\�^Q�>x�*^V�E���W�,��X��	�Ӿ>9�>���M����{=�贋�{/����I��|�Q��>�CS?G*�?b^��ݐ�.�g���Ͼ��N���>�y}?�i>��>$C?� �����¾��_=�+�?au�?ic�?Հ�=��=}�b�&��>��?娖?�?z�s?��+���>�Ú���>�j�����=t�>�z�=z6�=�d?��?�?X^���s���������j���<k¼=��>G�>P�u>PV�=�j=�]�=$�L>��>*��>Hh>�j�>[ш>���y�˾�G/?�����>��?���>ͦ%=�:D��^V>��[;Cã�o5��Ŀ�GX=�>�O^��()<���=9��>�����?�=M�	�K0?=���_W�>��`�>��ܽri�>�%A>�gZ>��>N��>@>�=�WH>��G> =Ӿ�j>��<R!��4C��xR� �ѾHz>����| &�������=I�k��^g�/j�/���>=���<�H�?�{��&�k���)������?�W�>6?ӌ�`戽m�>���>���>P��ۏ��=ʍ�b���?9��?*�c>�)�>��W?��?�2�H[3��lZ�l�u�$=A��e���`�捿������
��<����_?7�x?c�A?��</pz>���?�1&�[���q�>fI/��;���@=oҦ>v2���3`���Ӿ�Jľ�I���E>;�o?�G�?�?�nV�C�ὍV?�.(?���> U�?<O?��]?�<2> �#?R���[��>��>�/?N��>n+?s G��Q�kD��\G>#
'�e���
ǽ,��h�;������s>���5�<<�g�R��=�W���ݼ�㙽R� ��6���!�=(�>���=�ѧ>��\?�@�>Qǆ>{S7?��,�7�[���g/?�H:=7z��)䉾	|�����F>6�j?�"�?��Z?7If>�A�QmA��M>
L�>�2&>H&\>r�>�:�F�q�=s�>>;�=vlU�P���
�$D��뙲<ό>���>ӡ~>.���u&>�W���x��b>TsQ�]㺾[S��&H�Yb1���u�V��>FL?�?\��="�����pf�WR)?7�<?�M?��?eǓ=�ܾ��9���J�
��s�>���<���.���W꡿sa:��
�:��t>��������a>
r
�D�۾�nn��H�m\��y>=s��]Y=���پ��|�05�=}s	>�W��9g!����b��XJ?E�s=���+WP�y(����>��>�ٮ>'!��s��k?�+*���={��>�5<>g3���	�n�F�Ҁ�b1�>ME?dW_?:k�?*���s�b�B�ݴ���Z��a�Ǽ��?�U�> f?�A>��=]�����Y�d��G�3%�>��>���+�G��O�����$�v��>HA?Y�>�?��R?�
?�`?*?tC?��>��������B&?4��?S�=��Խ��T�z 9�HF����>b�)?z�B����>V�?ڽ?�&?�Q?�?!�>� ��C@����>�Y�>��W��b��M�_>��J?Ӛ�>\=Y?�ԃ?f�=>i�5�ꢾ�թ��V�=�>��2?�5#?8�?���>�l�>d�p�V�%>أ>6�\?�%�?s�?�yl=s�>w�b>Hz�>�E>z[	?v,�>�e?�;?�|?��V?+i�>�ě=(�˽vÿ��~"�&�e=��=��U=԰=�o�\B+��Z_��b=����
=��;�l�;ܻѼ�}�����5��>��s>Z����0>��ľ����=�@>=��>��c銾I�9����=�1�>��?�@�>�#��ʓ=�ϼ>���>���j(?^�?�?zK;�b�d�ھmhK�lذ>�1B?K�=�m��{��Y�u�^h=�n?~^?��V��n��*�k?y�P?�l��_�_� ;���J��K�㾖�Y?�c�>�ӯ�2�S>!�?y�:?}E'?�܈��dZ�w���A(n�h8��4�s=뭡>Կ5�(���	��>��D?<b�>$3>cD�<�)�_���ۅ�,r3?O�?���?8L�?�����{�����# �Lp���LX?���>m�6�!?�B����־���}�����޾�[��󼟾�t��6Ǥ�=�� <��
�Y�=��?�=w?K�v?W@`?�����\�#Z��V|�GL�F>��8B���G��/A�<i@�+]h��`���Rˠ��<�G��\6H�X�?�Pc?�i���?� �;���׽ʸ]<�;r�K�����=\��~=kgd>�:��j����۾g�<?�s�>\��>�T?��}���@���S�!������t=<H>i��>�	�>������<�����hˆ����7v>�xc?f�K?��n?�p��*1�����@�!���/�*c��m�B>�h>ۻ�>��W����:&�rY>�(�r�@���v��6�	�ݥ~=o�2?�'�>���>�O�?�?F{	�mk��kx��1�ߐ�<�1�>� i?�@�>��>�н&� �!��>P�f?s��>�כ>x7A���)�M2���8��w�>ѧ�>�U�> I>wa��rJf��턿1��h� �\x>�|?�k���?��ik>�f0?�;��;L"�>���;a�It�Tc2�=�y>K�?{��="'g>��;_������jRb��2(?^�?����*J*�6;�>��"?�D�>Q��>,��?<�>!�¾�aA;�i?�X^?+J?��@?���>M`1=۬��piŽ�!'���;=�w�>��\>0W�=�l�=�$��tb�v��uE==���+B��v�<ͅ��^*X<��<�N3>�ؿN'I�+�Ӿ9���d����型��"罥c�����������4�]�f�$��8���8�ep�ޡ���}Z����?J1�?j��So��2�w��^��D��>��O�<�7��x���)�}���ݾ�ॾ�.��V���h���d�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@tA?͸(�ݏ�m�U=�x�>�f	?��@>W�0��I��ాՉ�>�.�?��?�K=<�W��H
���e?҂<[�F�tg׻���=Ҩ�=�%=���4J>U��>���A�A��]۽S45>���>�"�����^��/�<P�]>�սX���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=S���	�����%�4����	=��=�h��(�(�(.$�	���ʓ��8����>�s�x;��=hZ�>d׌>j>>�oz>��V?s?�X�>�Y>66d��.v�#Ծ�}�-�x� ��猾c�i��[��%�龫 ܾ'�����6�^I �[�ľR =���=7R������� �.�b�<�F���.?/u$>+�ʾ��M���-<Upʾ�����Є�7ॽ�.̾a�1�/"n�͟?��A?����5�V����Q�����׮W?�O�ͻ�W묾ܡ�=B�����=�%�>ӏ�=���� 3��~S��
0?�G?Q=��Yu��v,>�3 ��=��+?�� ?�?T<J�>�]%?�,.�K޽n�\>&�5>�e�>���>4�>ϝ��::޽�?6ZU?����B���
��>`ǽ�	0y��]`=��
>2���̼a�V>���<Z���
;�g���N�<\�h?��>>�=��~�8׾y�ƾ��J>���?�r-?~�->�u?gIA?q0o=��辫 ��$U�؀3>��\?��k?`�A>���[￾6^��d?7[^?����Q˾%��{c?���7��5?��7?S��>�څ>�d���fg�nG �ei?d�v? T\� 1��2��qAd�̙>)"�>*�>{�7�1^�>LdB?~n"��Ĕ������'8����?��@ �?r.< ���p=]l?y��>�N���Ⱦ���Th���t�=���>����!#v�Z�����6?ě�?��>k�{����R��=�[���"�?片?kz���'�<��G�l�UK ���]<zĨ=�+9��[����P7��(ľ���Ea���q鼉r�>�@9���Ds�>!�=�����Ϳ���� վ��m��?�j�>R ��⤦�Ȼl�nu���G���G�蚈�x{�>^�>���J둾��{�8�;��뛼qd�>s�ވ>��R��嵾ɟ��)<�X�>c�>ˆ>0୽�ɽ�Y��?e����$ο}�����{X?�j�?�v�? j?�<<��u��{��x�	MG?�`s?�Z?9�#��]�B1:�΢s?������V��2�J�@���.=�#?�*�>q�����@�w>%��>	c��4��a���V���|����?�a�?�l<�>���?�?v�����.|����(N����o?ޫ�>�����=��ᅾ��<?��*?,�=:C�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?2�>��?	w�=�\�>O��=�谾��+�Hi#>>�=:?�\�?Q�M?|N�>qY�=�8�/�8WF��ER�1"�J�C���>��a?r�L?*Fb>*+��"2��!��iͽX1�[�輏d@�K�,���߽�5>U�=>�>.�D�pӾ1�'?�%��.ҿ����/�~`?+;s>��?��ɾ[o�����:|�`?��U>�P�	����.�������?M��?���>k׾<��tV�=!2�>��j>�8��]���O��,]V>�D?QKp�G����Cg��x{>�=�?NG@��?}%e�(|?׏ ����ELx�3�
�Ggg�u�>��>?�{�ʓe>3�?�"�=��u�8���A|�ׅ�>�?jY�?!i�>�ge?_2q���:��"�<nh�>�![?S�?Sf,=�n�j�h>��?���q/���%�0[?�D@�:@�,^?����8ο0���8���q��+)[>��=Q:>����~ґ��X�>lη;��3��-2>0ě>���>� �>>U�=g	F=��%>��}��� �����#S���W��n����#�����v��\ڇ�g�ݾ�g��b뾌�˽m��<G+=�ş�?0��_�j�|�=�VW?I�P?}>l?�?�P��o)>�����$�<Ĭ'�&Z=V�>�g2?�)K?�)+?Ň�=�ʚ��Wc��Y���!������$�>ӑU>#4�>o�>���>�e+J>�$A>�I�>���=�_;=�`�,��<(�?>��>�B�>�9�>Oz<>:�>�̴�\;���h���v�.x̽���? ���,�J��7��(�����r��=�k.?R�>����Bп~����H?dŔ�"���+�C>R�0?�VW?/^>����]!T���>o	��dj��>����\l�Ѓ)���P>$Q?n�f> �u>s�3��q8���P��d���G|>�.6?綾0>9���u�ȗH�#cݾd�M>�>��=�&_�������a�i�Vs{=�y:?��?�������Ѕu�;���kR>\>ڞ=�׫=�5M>p�d���ƽ�H�ۋ/=^k�=;�^>��?J�
>�|=
��>��a���C5�>��>�K>J-P?j�C?��Ͻ|���,h� ����Q>t@ ?�"�>$�=�Y����=��>l7�>�hi=�qW��X�k9���R>�:�=Z�Y�f����kM=�ͻãL>Q��=A��m���f��~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿj�>Fw�0Z����X�u��#=/��>9H?PR����O� >��w
??�_�멤�B�ȿ�zv����>z�?.��?z�m�dA���@�1��>r��?fY?nmi>�f۾ bZ�ۊ�>��@?R?��>�8�l�'���?!޶?���?oSK>\c�?�9s?C!�>$�n���/� z���싿;�~=Je�;8��>�K>U$þ��F�7z���_��k�i����2�f>�$= ��>��㽾���[H�=WI��9���vfc����>��l>~�H>Y�>� ?o��>;�>�=�W��.̂��╾�C?l��?f�����OgR>:8�=@܁�k�?%��>��.�X�I�|�>q�*?)�?�)o?�j�>��&N��O�ȿdh����N>qp�>I�?/�>��e=0`>��վ��,��2�>{�>:İ��Ǿ㶾�Xٻ��>G|6?�
?)�=(V)?q�!?�d>�e�>aq4�!���h|C���>Ql�>K"?��e?66?����@��sn���D� �H>u|?-�?��y>�!��>���2�XOýB�=��?Y�N?��U���?+��?2�9?zVP?�ux>ة���'��ɺ����=o�!?��(�A��R&�~��}?eM?c��>�H��Vֽ��ּ=���{���?�)\?B&?���:/a��þ���<��!��4V��X�;D���>�>���Ց�=U>���=GYm��=6��Eg<0t�=F��>� �=17�^���[4?��:�W�K�=�N^��uP�pq!>U\�>4�|?q�:�
x�P ���V������wu? ��?���?�Q]X���E?�W~?i�?0�)?f;t���&����zut��:X�Z�;�
G(>���>�뻽]ly����쵤�-d��2N<m��n��>u[�>]?D��>zXP>Ǳ>6���i�&�=����\A_���q8�#u.���$s���$$�z���2��(F{���>v���Id�>|�
?J$g>v�{>�.�>�Wǻ���>�#Q>B�}>���>�dX>{5>eC>�='<�1ҽZR?U�����'������� B?#\d?�G�>�e�ᕅ�d��\�?�w�?iW�?��u>.�h�k+�\a?Ĭ�>��/d
?k�8=�h��3�<�$���<�`	��$:��l�>��׽  :��7M�.�f��k
?�0?P��ϕ̾VOֽ(Y��e<���?��:?Y=P���:��Kp�<�Y��f��ϳ��^G�� ����j�l�P򍿍qk�˚����"�/W=�>?���?��C�Js�at�٦���S��>�O�>iR�>�_�>.�>B�\Q��I���3���½U�?L�?�L>w�d?#�-?��?]�X?��> ��>ӯy��9�>_��v�=��?�+>?��#?�	:?��?m>-?�3N>��n�ط��M��E{?�-?�/?��>��?�@��:�J�h�ݼCa}=��c��>�͞����]�e����-����>EZ?
��ū8������j>�|7?�}�>,��>�	���3�����<^�>�
?A�>j ���r��_��T�>6��?-����=x�)>=��=�d���Һ�B�=�¼��=$T��{|;���<�V�=��=Tgs��Te����:�(�;렯<֕?*�?�>&&�>D����5�3P��p.>GnN>�M>��c>��Ͼ�鈿�U��t��i>}��?�ʴ?Lo"=���=�=��������6tžE�Q=�	?F0%?�T?]B�?Rt2?Z$?3�6>L��܌����|��Μ�0?w!,?��>�����ʾ��׉3�۝?l[?�<a����;)�ؐ¾�Խѱ>�[/�b/~����8D�����j��4��?쿝??A�T�6��x�׿���[��y�C?
"�>Y�>��>R�)�z�g�r%��1;>���>iR?�#�>�O?�<{?¦[?�gT>_�8�n1���ә��G3���!>9@?��?�?zy?�t�>��>ع)��ྑT��q��M�.ႾUW=3	Z>o��>�(�>I�>d��=�Ƚ�Z����>��`�=��b>U��>���>��>�w>�L�<�H?*;�>7p���<����|=��ٗ.��=v?�-�?�+?%*=��E�6E�����>1֧?�ʫ?��*?3(T��,�=<,�����q����>��>���>UG�=5N=#�>�^�>���>N����8���J��?��E?���=F�ƿ�x��!������#�_=�\o�;$a� &�}�z�a>�����s�����>�/Xw���l�:�¾�����z��E�>p��=�k>@P�=;�5�s;`�l: <?o=�<>V���(���je<{����2��dk��9�-��,
=l��=H�R˾[��?�'B?C^#?@�J?��w>&�.>����"�>Z�0��r	?JRM>hFw��\����eF��+;j�7�̾4[����g�W���E�=��w����=S�>恁=z��z_�=�E=��=tf�[Q�7|=S��=3�=Fw>���=Y@>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=J����=2>q��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�[8>�>��R�#i1��]��Kd�{�X�k�!?m;�7�˾+9�>��=e@߾��ƾB&=�b6>F�e=����H\�y��=!=��>=�xk=���>�RC>\*�=>)��D��=R�L=��=/O>Vd���1��b+��,1=�4�=�rb>)�%>)��>j�?�a0?�Wd?�6�>�n�kϾ�>��xH�>|�=E�>���=.rB>ݎ�>��7?��D?��K?Y��>=7	�>��>w�,�Z�m�k��ʧ����<*��?�͆?�Ѹ>��Q<��A�Ѡ�}g>��+Ž1v?�R1?�j?k�>�> ���ѿ�7Y�J��Y�(>�7>&�Y������̽��>�w���|��ӎ���s>>\P�>Q�>#Ԓ>�Y�<u5>���>��>�+�=Y��=;h�ą$�\�$�2<K>�=|�6��^̼��9����=�罂Dl�P�<=��>�_?>z�r=%!�=��>'�>M�>׮�=�w����$>������K���=�	��7�A��he��}���.�,�8���D>�\>
s�䚑��\?�Y>f8?>v��?5�t?}8>�r���վz���o�|
N��ܲ=�=>�[7�=l;�$S`�{�N�*z;���>"��>� �>õl>�,��%?��Ew=��ιX5��>\u�����6U�8q��=�������i������D?C��̴�=�~?êI?��?5��>�e��;�ؾ�)0>�F��]H=W��9q�����Z�?c'?���>i�N�D��=��(�	�>`E��X`�׍�� ��`�=rP��K�Y>� a�䐾k6&�Gz������@���x�֭�>�F?�+�?�;R�񔆿�@]�C��';���F'?|}�?}Ϳ>%]�>N�&?������0�l�%䭽�bV?[i�?���?7�o=	�=�)����>o��>j>�?8Ώ?,�y?p�K����>n$<S#>I�A��},>�f�=]��=�ڮ=pJ?�y?[�?&�h���d����G�A��=Z`�=��>{=r>��>o��=���<��q=P>
��>�G�>�v>R��>-��>cʶ�� ��NA?m�>?�e=|\J?��=	p�.A>�R=S�<���Ƞ+��3ý���sx4>|X��-�Ƚ�O�>�����Ў?�>��ʳ-?I�	�B�X�s0�>�V>;l���f�>a��=>�>�ª>���>��*>b�>j�=h:Ӿ2s>���X!�Y4C�V~R�c�Ѿ�`z>㪜�'&�C�������#I��s��=j��j�2���:=�X޽<�H�?mO��Q�k��)�������?�h�>K"6?'ٌ����Z�>;��>���>�Z������8ȍ�T���?���??c>\�>��W?��?V�1��3��wZ�?�u�H'A�+e���`�#፿����L�
�E	��6�_?N�x?syA?���<f8z>0��?��%�8ҏ�-�>o/�4(;��4<=�)�>s+��}�`��Ӿ��þ">�2LF>e�o? $�?�V?�JV�����`�>��1?��?�4u?5�%?�IO?[���� ?���=Zf�>��?�>?�?�?Zk{=�[2>It =��=r覽q���Q�����X�R�� ��;��<�nؽ@��<�28>_�=�1��s��r��Q��MԽ��=3n>p�<>fO�>)A]?���>��>)8?��&�!/>�13��V ,?d�=�^��݊�QM���g���P�=�c?`ҩ?ܿY?6�{>��?�9);�%�>�6�>� *>�,X>�"�>���6H�u�E=�5 >�V(>}s�=�{�/�w���
��q����B:�G)>���>	߀>IÎ��s">�\��yx��Lc>|O�֤��o\S�ƓH�N�0���w����>?-L?�{?��=�1�a��3pf��r(?o<?�;N?1?�L�=��ھNf9�մI��"�˲�>8��<@���ڢ�򶡿"�:��V�;�mw>�o���Ԡ�̈a>>�
�Wsݾ?�n��I�Y��UH=����]R=��־�i~���=P�	>����W!�@	��v���`J?�h=  ����T����h^>�?�>�v�>f�9��w��h@��ʬ���=�y�>�:>�������ʙG����>�>@QE?+W_?k�?�!��\s�V�B�f����c���ȼ5�?Rx�>�g?�B>���=V�������d�xG���>ʠ�>[��:�G��;��a0��<�$�*��>_9?��>k�?]�R?��
?u�`?�*?4E?'�>�������B&?0��?��=4�Խ��T�� 9�TF����>m�)?��B�й�>E�?ѽ?��&?�Q?۵?��>� ��C@����>�Y�>��W��b����_>��J?>w=Y?�ԃ?]�=>Q�5��颾֩�3V�=~>��2?�5#?@�?�>���>Dv��k�=;��>mc?�?yp?�B�=}�?�0>�1�>���=���>!��>L�?��N?X]s?# J?
��>�}<����J��h�v�BI��J��:�,g<$xj=n��>��9�KQ=c��;�ӵ��6���߼�|F�2r����;�_�>>�s>�
��'�0>��ľO����@>�1P���ي��:���=���>�?���>~Y#����=��>(H�>���	7(?��?K?`w";>�b�y�ھ9�K�6�>�B?��=3�l�r�����u��	h=��m?q�^?��W�>&��M-j?�sV?7�	���8�����>�����q.?�^D?�w�HmF�Y[�?rP?�� ?K����������r�$W��^�9�?�l
�^��,�>��Y?���=��=^���H����r��>����-�>���?λ?�9�?��>�p�sf��S�$o���qW?C�>�����*?�U�b��9����5��e��C���V����X���á��z�@#��*5߽�Ş=��?p?��?��l?K����O�X�\��Ir��!d�)���Y�F���@�mu6���Y������s���m�
��ם���?��q�?(M?N��"?�B�� �.�&��2��蒶��FM���i>�n@<�=?B =�Eľ��s���5���T?/ڸ>�F?_EP?!�v�9\<���2�ř���	��q�<�ؒ>�1�=
IC>���=��?����~ ˾]�¾�����6v>"yc?R�K?3�n?dm�q*1�s�����!�Q�/�1b����B>k>�>��W�t���9&�>Y>�6�r�����w��L�	��~=��2?h(�>鲜>�O�?�?U{	��j��jx�%�1�k��< 0�>D i?f@�>��>(н�� �Ͼ�>��l?5��>��>����}\!���{���ʽ��>�߭>
��>��o>9�,��#\��g��^���9���=�h?����`��߅>�R?�:GH<~�>�pv��!�>���'���>�~?���=�;>ˀž�$���{��0��j%)?e?A�����*�[�~>b&"?���>*S�>U�?�D�>+þ+5��?1�^?SJ?#A?X�>�D=t���ÇȽ�'��(,=RS�>�Z>�dm=���={��k\�O��!(E=s��=�Cμ��<i<�$���N<���<��3>��ڿ��K�N�׾���L��x
�d����½��� 	��X���P�� �m�����p)�]�T�܋e�[X��J�k�p3�?�4�?�+��k1�����"�}�}���E�>a�~�����+�����\����ݾg#����ӎP���g��Rf�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@~A?��(�^�쾈HV= ��>�	?R�?>�P1��K������Q�>�:�?��?�VM=@�W�6�	��e?�<��F�\�ݻE+�=�9�=�E=�����J>�T�>�y�2HA��Dܽ7�4>�݅>�["���р^��^�<�]>~�ս",��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�}��=[��>c�>,������O��I��U��=�����¿Ͳ$�M~!� �<�K�=��/Y^�+<(<⟾�JȾ²E�P^&�^�=^L=��,>�iy> p;>ԛ>>eX?�R?v �>I�>�d��Y�&��cݾ^I������bk��U�D'��>���棾"2� �$������J=��R�=�8R�^���� ��b���F���.?�w$>��ʾ��M�]/<mdʾk����������V=̾ӟ1�A%n��ğ?=�A?�󅿓�V�����u������W?������ެ���=-+����=W?�>^�=2��x3���S��{0?�S?7r������h*>11���=��+?�j?�B^< �>�5%?�8+�z?�6�[>U_3>��>���>y�	>���0۽cv?nT?�<�	䜾�!�>@��z�5�`=ck>�4�w����[>�Ԏ<�匾LY�u����6�<�Kd?��g>��"�{~ϾVl��/@O�Q �=W~?%�?2r>�&R?�J?kS=��ξ+�j�y�,�� :��z'?��?1Ž=D�=�5þ鱾�'?T�w?�>�|��WI'��74�
�&�%C?1��?H�;?�}��W��3�l�+��B$?�{?��l�:%��㑮���Ⱦ��߽t��>�*0?#��>�?0�p?���&����zĿ�.G�Lպ?�i@y4�?C���ּ!T	�G��>@&�>�s�YJ��c�>��h���+>�
�>y0���Wq�Q5��=�� ?��_?��>.a���������=�ٕ��Z�?��?ۄ���Ig<j���l��n���{�<Ϋ=.��D"������7���ƾ��
�<���T迼��>3Z@�V�n*�>�C8�^6�TϿ ���[о�Sq�l�?+��>סȽכ��C�j��Pu�T�G�,�H�@����V�>\�>{����푾��{��s;�L៼ �>�#���>�S�4&��ؠ����4<��>���>ȼ�>���	ֽ����?F^���<οΩ��Z��ݶX?]j�?o�?�u?�9<B�v�Jq{��&��.G?�{s?�Z?8�%��O]��7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�O�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�$N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>dH_���u>����:�
i	>���?�~�?Qj?���� ����U>
�}?5b�>���?>�=���>>.�=�Z����s��M'>��=i�4��]??XM?۟�>/�=Ay2�A�-���E�eR�v�+D�1̅>��a?mN?�cc>5ص����l� ���ͽap-��Ϣ���C��h/�����2>��>>�{>X�@�<�;��?Jp�7�ؿ�i��8p'��54?+��>�?����t�����;_?Bz�>7��+���%���B�_��?�G�?>�?��׾�S̼�>@�>�I�>��Խ���Z�����7>:�B?j��D��w�o�{�>���?�@�ծ?gi�ߟ?���L����]�Fg��؊���>bu<?`  ���>��?�Į<��~�ZS����r�R/�>>A�?��?���>y�]?U��Q�7��6:��՟>��K?��!?y�7>��׾���>�x(?��+������I����^?v�@�p@N1k?��(�Ͽ���"��X���{��=�4Y=3i:>�e��- >�=�@���H�I�4>��>e�`>�߀>IP>��2>!�>���ō$�R����B�J�6�$����A� �ݾGd���VbǾ�����̽]���嗽�!7�Ik���.����=��d?m7N?�T[?�w?����I�=�@;�4����ǽ�Bc=�֎>Pi'?o�R? �/?®�=t�����c�y�h�-ܾ�i4��T��>��>.��>!�>�>�@���D2>]�[>띥>�s=V�e<D���٬<��N>�_�>���>���>�C<>��>Eϴ��1��h�h��
w��̽/�?~���Q�J��1���9��Ц��i�=Gb.?	|>���?пf����2H?���x)���+���>{�0?�cW?'�>(��g�T�8:>8����j�7`>�+ �ll���)��%Q>rl?�f>�/u>�3�Fg8���P��v��?T|>�46?9鶾�A9���u���H�]_ݾ�ZM>dɾ>��C��k�/�������i� �{=�y:?��? #��c߰�<�u�+A��:LR>X9\>y�=Q�=RVM>��c���ƽ.H�k�.=���=��^>��?/�&>�1�=��>�F��̖]��И>��@>>�d>?�"?�'��㽽�����#���j>��>>2�>a�>�I�Ds�=T�>)`>L�ռ��\��N�I_2���a>]󇽸-g�o�:��
�=i��~N�=dY�=���}C���N=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿuh�>ex�|Z��}����u�:�#=^��>�8H?JV��[�O�`>�w
?�?�^�穤���ȿ9|v����>[�?���?9�m��A���@����>A��?zgY?�ni>�g۾l`Z�7��>ܻ@?�R?K�>�9�͏'�O�?�޶?ɯ�?�,I>k��?��s?z�>��w��]/��8��R�����~=P�\;�]�>uN>(����hF�`ғ�2g����j�K��p�a>3�$=��>�=�Y.��@M�=9ɋ��E���ef���>�q>��I>1_�>�� ?�d�>��>:H=�w���倾Ъ��ى=?��?��(㋿�a,>f>r�?�?g�<{G �W�>l�<?�1�?ؙ[?CGn>sC!�O)����������/>?n�>��?C? _���}Y>v2O�eS����q>�1�>⻽��� z���!>�L�>D�2?���>��=Ã"?z� ?w�`>-s�>�D� `��A�C���>�3�>{c?�#}?�t?R���
2�v�젿&�W���M>_1z?��?j��>V
��N"������!?��B/�dف?(Qi?���T�?�ڊ?#�D?9hB?+D>�=�B�ᾬֽՀ>j�!?'���A�M&� ��~?�P?���><��O�սv4ּ����~��'�?b)\?�?&?��^+a���¾�1�<�#��U���;��D���>��>n���k��=x>6հ=WLm��E6���f<ck�=2��>�	�=�*7��s����D?P'?�U.���T>�:X��sr���t<��g>��z}B?fl=�
��B��k8��+����Ճ?:��?���?ዖ���:�A)L?(g?&??Y?��A��b�\�g־�t�cI$�̛�>���>{t���l�> ��ζ����#��=������>*X�>B!?,B?�>>�ɢ>[얾�	*���n����\���o59�9�*�I���̙�\F��Qu�ʶ���k��s�>G ��)e�>|?��d>t�>��>	J7�Ŝ�>�[>K�>U�>ZDW>u}->m��=�*�:�u��LR?2����'����ӗ���0B?�Ed?��>ƛh�{���g��\�?��?�v�?�=v>�zh��<+��C?���>	?��h�
?{�:=g���]�<hO�����t���8*�s��>f׽R:�f"M��:f�Ӊ
?yD?Sϋ���̾�#ؽ�vR��i��MԚ?h�U?��Z�%-�r���x�VB`�6�R�0h��?�¾gD��lHU��ԋ�Tc�zو�lA������M?��?"N�O8ؾ�-`��ԓ�-���\>q�>�v[>~R�>WC>�i'�S�z��b��V�ޱ:���?�6�?��>i]W?�A<?qPD?2�S?1�>ѝ�>>��V�>�#~=���>��>:5.?�4?)03?|?�?�:>?��� ��^྆?�=$?��?*��>n�?as�3�����<w1e=Q��掱�-�&D�<5R̽�G�Rk�=>Lx>t\?���~�8������k>�t7?#^�>*��>o$��g%�����<l�>��
?�6�>�����{r��Y��Y�>���?�6�=��)>���=MU���ʺOY�=��� �=w����;�?� <d��=)�=�t�T��@l�:�r�;� �<��?�H?mX>ƫ>��[�*���� ���>1>�p>?>"WӾN͈������BL��*>m��?�
�?B�=>���=���=�����ʾ�%��谾S9M>�?��7?37?�B�?��G?�=?
J>J�)�Y:���$��|¾W�?v!,?��>�����ʾ��Ӊ3�֝?j[?�<a����;)�ِ¾��Խ߱>�[/�f/~����>D�����X��5��??3A�U�6��x�ڿ���[��y�C?
"�>Y�>��>U�)�|�g�q%��1;>���>nR?�%�>M�O?.;{?��[?,kT>ȝ8��1���ҙ�l�3���!>�@?&��?D�?�y?Iu�>j�>M�)��bO�������x����W=
Z>Y��>�'�>��>���=EȽ�`��9�>�rg�=[�b>���>q��>� �>��w>�k�<yuM?pf�>�+ǾD���3���ݯ�z���Y6x?B�?��?�r�=�2�]K]�1�����>?��?k�?z�A?�UY�d3�=P�������Fm�f�>Ѣ>��$>bc-<qO[=�S��;�>���>1�(����fC;������?t�H?�4�=�ƿ��r����fm����=s�q��4�w���A��:�= E���o���J�}���M��=d���㕾��}��?R�7=��>x�>��F�~`<�%���������ڗ=@����ۧ�E�!M<��P�b�:�ּ��<��ջ&�ʾ�!?R&E?�7#?ROH?|�>�5>v�м�؉>W���L?��Z>�1S��r��<I �濣��玾v�پ{Bɾ9i������=��s��&�=$->��>eB�9���=0�8=A�=� �;~L�<�Ɗ=��=_į=r$�=�q>e�>�6w?^���󲝿s4Q��\��:?Z9�>�~�=S�ƾ�@?!�>>�2�������b��-?���?�T�?~�?ti��d�>���8㎽�p�=���=2>���=��2����>��J>���K��e���y4�?z�@��??�ዿ��Ͽ�`/>	8>*>A�R�$L1�"\���b�$0[���!?�Z;��,̾0$�>���=Xg߾6�ƾ��/=>6>�c=����\�Q��=�;y���;=��k=�׉>�D>OF�=0���{��=N�H=��=/!P>�)��v�6��+���2=[��=#\b>�E&>���>��?P%0?xvd?hY�>��n���Ͼ�������>���=��>�!�=DA>��>u�7?�\D?�K?K��>+ތ=�ź>-�>�{,�e�m�̦待������<t��?�ن?�n�>��R<�}@��&��>���ƽH?�1?^?�>���(˿�49�@dI���5=�$k=�X>܀���*>���
;���k�=��>�ܩ>��e>^�>е�>F�^>�>\o�>t�=NKg<W�$=N� =p6>�Q�<��Z<G�=��x<ֳ���0=(N=s��$jd���	<'E�=1/v�\u�����=�R�>]�>P7�>���=c۵���(>A��T�M��I�=�0��T�A�W�d��G~��.�0�7���D>�GZ>�z������?�VZ>�B>���?�1u?�> �� �Ծ֝�(�i�`�L����=�C	>�V8�]�;��_�2N��Ͼ���>vގ>8�>a�l>,��#?���w=���b5���><|��:���+��9q��?������ki��Ѻ;�D?CF��ޤ�=�!~?ǰI?s�?��>����ؾ�;0>�H��g�=���'q�#e����?�'?h��>��e�D�����HS��a�>Y����`��^��Z,�jۭ���Ѿ��;>������Ѿ,(6��$��=򐿾�4�zC��kv�>�^?
&�?E-�/
���YP��_Ͼ�ቾ�'?�ލ?�N�>?g ?��0?3s�/)&���ݾ8��=��?A=�?���?�#>�M�=P���#�>V��>��?F�?�ls?E;1��|�>B�<��5> �a�CK�=H��=��>��=�4
?g��>��?�E������ᾠ\���x����<���=�Xa>@�f>@>���=�T�=Ö~=�,$>|l�>ݟ>e�>p�>rÂ>٬�~��#?���=� �>cK3?��>==jY����	=Z"o��^8�Ѭ�F]��W�ؽ!��<�ꩻ�@=]M���>�[ſ�͖?�]>��
���?q���
:I�!9>dR>�4Խ�,�>ǫC>�o>��>���>�
>�Z�>�">8FӾ�}>���d!�+-C��R�O�Ѿ'{z>y����
&���py���AI�n��}g�mj�O.���<=�)��<?H�?Ϻ��d�k���)�����^�?y[�>n6?�ٌ�9��h�>|��>6Ǎ>�K��m���Kȍ��g�e�?U��?w�c>$��>�W?z�?&1�m�3���Z�։u�\GA�`�d���`� э������
��B����_?��x?BvA?@��<:�y>���?;�%�����,9�>#�.�;���==�Z�>X-��5Ga�JӾ	gþE���HF>�bo?D�?�+?<�U��v{���?b��>$�9>�
q?��/?'�N?e���S��>P�T>��?��?q�>F:?�[Q?E! =8͊������?�=�
�{¾�ZýK���D���Q*=LvG<�c۽o5$=��=~���x�㺌̹=2�.���ֻ����ڦ�1�=�T=ֈ�>>#S?�k�>H�>_7?�D��kE�Oo��{
?�h=ڑ���ӊ�gڷ�5���:�>��Z?#�?	Y?IL�>�?�����O>aa�>Fl>��g>�P�>y��������B=���=ڒ7>���=�G����� �Ȓ��-?�$�0>���>w;|>��_�'>Sv���+z�әd>E�Q�ͺ���S���G� �1�k�v�]�>z�K?��?���=�`��+���If�.)?^<?>QM?��?E�=��۾[�9�1�J�w9�T�>*�<���f����"����:�'��:)�s>*��࠾PUb>���s޾~�n��J����2M=8~�feV=����վ�6����=�#
>����6� �:��.֪�p1J?�j==w��ocU�6o��G�>���>}�>�:�[�v��@������4�=(��>�:>pY������~G�+8�,�>�\E?�]_?�j�?�7��;�r���B�m���%G���Ƽ��?-`�>�X?��A>��=2������e�
G����>���>S���G��
��Q*����$�7��>2?g�> �?�R?��
?��`?�*?�F?��>*᷽��� B&?6��?��=��Խ�T�� 9�JF����>|�)? �B�ܹ�>P�?�?��&?�Q?�?��>� ��C@��>�Y�>��W��b��>�_>��J?ٚ�>s=Y?�ԃ?x�=>]�5��颾�֩��U�=�>��2?6#?O�?���>[��>9����=<��>�c?!0�?9�o?̊�=��?�<2>���>���=D��>5��>?�WO?��s?��J?���>I��<�;��?���As�q�O����;OH<��y=E��Dt�M�.��<�ֳ;va��^.��%�񼢻D�r���M��;z��>��q>�˗��Q)>�����Ȅ��L?>'/��c㚾	ވ��>=��_�=!+�>�:?|��>Y ��\�=�B�>Z��>v���('?�?��?2�,�Jb�� ݾqsR�)�>$#A?��=a�k�"���u�.kk=��n?�^?+�]����O�b?��]?Ah��=��þz�b����g�O?;�
?8�G���>��~?g�q?U��>
�e�*:n�)��Db���j�&Ѷ=[r�>MX�T�d��?�>p�7?�N�>1�b>&%�=ju۾�w��q��h?��?�?���?+*>��n�Z4�Cm��{�)|P?�q�>Iؾ�?�5�����|#r�y���>ɾ���+ZžI���"�a�+|q�96��tC�W֕=g�@? s�?͔?'<??yN#�lj���m��Ԇ�Qu���"�����M���7��[��!��7����3ڊ���|>���.H�3��?��?�3_�\�>J��|����=�=ZM����νw�>{ޓ<r��=K�=� ��)����˾F-(? �F>�7S>�;?h�E�,IF��'��E�M��eI�=�;�>���>�,?P]>I&���P�����	c�ͪ���l>K�f?��M?%�p?n��-�9i~�5�$�<V�������z->���=	M�>�l�S�-��1)�*�?��)w��3��)�����@�=~+?cމ>��>OI�?=#?k������8�t���+�g��<�̿>	ui?$��>䯄>7϶��	$���>\}�?�?d�?>;���a����A��W��`�>�F>��?>�=2�pzt����(o��"�Q����<8�y?x.����b�Ǘ�>��*?����\o����=�~h�L)��c�#��x���dN>�^�>d+=r>�Y��@��0h���-{�о)?�4?����D,��`�>x�#?�G�>��>�؃?!��>d�ľ�� ���?��_?�K?�A?��>�=C���ʽ��&���=w��>R�V>��c=��=�����Y�y!��I=m8�=0��<�ý�/'<�3P�/�<"�<�/>b*׿̳G�G�پ�
�o��ߖ�=V��˱ҽ�pP�5���_������H������=<X���^���r������:�?}0�?���Yr�;���܃������>3��a��lɯ�|�������+!���
"���D���c��[L�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�)f?��T�:��J�?w�wߊ�+ܽ��Ͻ�Ԅ��:�0R�?3[�?&W�?j��>W�?��>>a�?uѡ��!��j?�;&��=�`���T��,+�=k��>�?p(B>�?��x�6�ց>_�;>~H>�wӼl�a�������>D�ѽ��+����?3;P��sn���D��`�1Ny>
�>?���>0 >_"?�I��&ʿ�b��[?���?5�?��"?��ˡ�>�Ͼm�O?��0?E�>���|��F>.�K=�Y��a���8H��+>���>��<S�F�@o��K޽O�%=&�n=�T���:����+�
���l(=�͊�y��l@u=���:�h��1�Q���t]=D�5>](>^4R>n+�>�+>�6W?�rn?�>j>�����ڰ�}���]��<�ܠ��넾aҖ�K��#����)Sþ�O����ܮ��t��Y"=���=�7R������� ��b���F���.?9�$>��ʾ��M�F�-<Lpʾ6����e���楽Y-̾��1�"n�̟?��A?Y�S�V�������`�����W?-\�g��@쬾{��=g���b�=&�>ტ=���� 3��zS�*�0?)K?}��y����*>[� ��b=_,?*=?|T<̓�>��$?�-��q彺9\>�,7>$�>�>v�	>Vj����׽��?�)U?f*����E�>���r4~�L�_=�U>�W6�K[���Y>��q<�Q�7�a󋽀g�<q)W?���> �)��c���#�8x==��x?�?�>�k?q�B?gʥ<@\��O�S�}���w=��W?p i?+�>t����оΔ����5?�e?(�N>Th�M����.��Y�`?�n?>]?$e���t}�V��{���l6?��v?�n^��r��#����V��:�>Z�>���>��9��g�>*�>?N#�eH��l����T4�SŞ?V�@��?+<<�I����=�>?Cj�>նO�bGƾ�J��Ň���q=��>�����ev���� _,��~8?0��?&��>7��������=�ؕ��Z�?)�?ᅪ��1g<���Al��n���g�<ͫ=C�/M"�����7���ƾϼ
����׿����>AZ@�M�Y)�>jG8�6��SϿI��S\о�Tq���?��>��Ƚ�����j�-Qu��G���H�ˣ��4M�>h�=͔;�ᖾ�wy�̾9�\��{C�>����rU>�^��������t�R<q�>.��>�|�>Sv6�	�����?�N��\ѿa[��5/���=?]�?��c?R0?�N��/�+����C�;>Ťk?b+�?|�]?'�=��o-D�!�j?�_��nU`��4�uHE��U>�"3?�B�>P�-�9�|=�>��>g>�#/�x�Ŀ�ٶ�H���U��?��?�o���>p��?rs+?�i�8���[����*���+��<A?�2>���D�!�A0=�RҒ���
?O~0?G{�c.�_�_?+�a�.�p���-���ƽzۡ>��0�&f\�
Q��d���Xe�����@y����?>^�?_�?f��� #�J6%?6�>����!9Ǿw�<���>�(�>�)N>�J_�I�u>����:��i	>���?�~�?Yj?ߕ�������U>��}?ca�>�1�?���=���>���=�;��o�4��>��=�$5�z�?��L?E��>���=A2<�P�/�Y�F�R�R����C�2�>�xa?�pK?N�b>�?��*�*��� �_�˽fE0�v<�2?��'�xU۽��6>�>>�F>�D��CԾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���E���`~�����
7��V�=��7?M5��z>B��>��=5lv�b�����s�챶>
?�?u�?���>8�l?��o�F�B�2=�M�>.�k?m?q���T|B>�?u��%���`3��)f?�
@�u@Q�^?���п×��n��&�����>/ě='hO>䥽���=���=�<ӄ��t��=H�>�8q>�`k>i�[>�R5>=�>�M���$��m菿�/4�J����#��1��a�ڿS����_����k��%����I�O�����h��uL��[�|�=�<V?�R?�)p?Ƹ ?�
x�y">�;���=ov �J��=R�>�{1?�gK?-�)?+��=hϞ��De�����n����Q���L�>_�I>���>+��>�~�>�V];�GJ>��<>��>� >��'=�k̹a�=��O>r��>`��>{q�>�C<>��>Fϴ��1��h�h��
w�_̽0�?����X�J��1���9��æ�� i�=Bb.?|>���?пg����2H?$���{)���+���>��0?�cW?5�>����T�	:>K����j�B`>�+ ��l���)��%Q>vl?�f>�u>֛3��e8�n�P�f|��j|>�36?X鶾'D9���u���H��cݾQHM>�ľ>�
D�l�|�����'vi�T�{=]x:?߄?
7���ⰾi�u��C���PR>j:\>%U=�i�=�XM>�bc���ƽ6H��g.=!��=֮^>_U?w,>M�=��>l��d3P�A}�>�hB>�,>
@?�%?x�����^���q$.���v>�9�>~�>�>�oJ�+��=�i�>��a>K������^����?�B�W>d�}��n_�Hu�.y=;��k��=�Ǔ=�� �z7=���%=-�~?�~��8䈿��VQ��>oD?�)?_�=4�F<�"������N����?C�@�m�?T�	���V�{�?MA�?-����=�x�>�ѫ>�ξw�L��?�ƽ�Ƣ��	�##�hR�?��?�/�
ɋ��l��;>,Z%?;�ӾNh�>px��Z�������u�f�#=G��>�8H?�V����O�j>��v
?�?�^�੤���ȿ6|v����>W�?���?j�m��A���@����>:��?�gY?�oi>�g۾&`Z����>л@?�R?�>�9�o�'���?�޶?կ�?y'>ZӒ?�u??�K�8��uȢ�H���L�=$��=��7>n�=	z����U�+O�����e�o�Dh<�ۆ�>�MV�#��>Ҵz�%���K��= �Du�����0C�>\ge>��8>Ӗ�>�i�>.��>�u�>�B1=򸦼�Eu���˾��K?���?-���2n��N�<^��=)�^��&?�I4?k[�}�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��N��<��K>*4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��fS��HB�>�e!?���>�Ү=;� ?k�#?	k>���>WvE�l-��[F��!�>��>!?>�~?��?���t3�����f�[��N>t�x?�h?�Q�>�q��zy��pY:�R�G�:���M��?�Yg?
�⽬�?D!�?ar??z�A?�e>@��4�׾����i�>&/?�_.�=\�5$\�X�=�<?S?�>��>��<8;�������B��� ���,?���?�,H?���qV�F����a���<a���8jb�ښ���=�t�<ׇ�0fK>���<���=�B;Ymݾ�kT���>1�?��4>g����}3��.?N�>�O����=i�7�Re)��|�>��o>���t& ?�荾m܃��y���#��D\����?���?�Ɯ?�&ؼXp��uH?B�?��7?A��>�}����=��%���;ަ����1��=s��>>� �wo%�}r���ڜ���E�nϼ���@�?69�>�?Pƽ>�tC>$��>�>������<о!����T�z�,�B�p�6�41(��ľ�El��f�<��Ͼ|xK���>%߿�'ج> ��>NR> <m>2�>�>��P�>�g>^�>�$�>���>N�>-�=f�u8��)i?�����nV��9���>�P�?oH?�~?�X=�uZ���/�1�$>W}�?��?���>��C�Z_�c�9?�E?-�r�	 ?�` =�5ּ>~X>.���g��?d"� �{>��&?��V����胿(�g�O?��?0�o�g뤾<q�>����?�A>��?x?�WO�UiK�|?����0B�q�X��ۂ������<*�����Z��${��%������m>��@?�Ѐ?T���ﾯ9����G�I�@�V�T>�/�>
߻>%~�>7��=r���4��s��'��馾�}�>M9s?*p�>E�I?4<?P?�wL?m��>�z�>6%���r�> ^�;Q��>M��>��9?�-?�/0?6s?Vc+?�b>�T�������ؾ
?�?\Y?<?��?�����*ý�q����e�֮y�v����Ё=���<��׽�u�E�T=*�S>�X?���h�8������k>_�7?��>q��>���j-�����<��>µ
?FF�>~ �@~r�c��V�>���?� ���=��)>n��=*���]tҺ,X�=������=�4���z;��o<���=���=X?t�������:^e�;�o�<��>�6?39�>S�>`�9�}�Ǿis��#ȃ<s�:��0=��-�2�������霿�/r� 5j>ӂ?���?��K>��y< �>����!�Z����ܐ��-����>�-??�@?/�?�0?H�/?��=,�Ҥ�&Y��kW���K?K!,?���>��W�ʾ��c�3���?[?D<a�����;)��¾��Խ��>
\/�z/~����JD�9������������?���?�A�Y�6�#y�࿘�B[����C?"�>Y�>|�>A�)�8�g�#%�L1;>:��>
R?B��>_�N?�z?��Z?�(R>�M9��=�������M�H%">��@?���?��?g�x?���>��>�'��J�����ͦ���������U=�Z>���>$!�>�n�>@5�=r�ý�@��r�<����=�C_>AW�>�ȥ>�{�>�s>6�<k4O?Ŷ�> ��0R+��&�D�սF棽.L�?���?��?,k~��F�B�W�v�޾L�
?�;�?Q~�??�4��g��=B�=�V�wYw=��w>p�=�,�>�P>�64���=bc�>e%�>��Z�>d3��T��Sټt�6?C]?g��Q�ÿ(aw��J��2Et��ý��>��D8�ɓT�D�=G��>��a��,�����-�5��Q���ž����s����?@?�=V=�<��<˚Ի���=%D��k�)<���=#t$�J6ֽ0P�;7���º���9���鼃(<��:<����۾�x�?�s?��R?�M\?G�>��?��F�(>�>D��=�=�>�%>,�l�ﰋ���'��R}�2'��)M-��cC��ۅ���ɾ_����z��o�>��>�M�>V�D>e�|=n��<��)>��=%<��>�d�=��5>Y>�T>�N�=�6w?W�������4Q�vZ罩�:?�8�>n{�=��ƾq@?s�>>�2������rb��-?���?�T�?;�?*ti��d�>M���㎽�q�=[����=2>P��=��2�T��>��J>���K��u����4�?��@��??�ዿТϿ*a/>T8>�K>`�R��e1�G�\���c�w�Z��z!?=T;��<̾��>���=�j޾�4ƾ�,=�6>��f=|��l�\���=��y��(:=��k=̉>�	D>F��=V���]<�=h	I=��=��O>�F��DV8���-�C�3=o�=Q*b>�%&>)��>��?�_0?}Qd?�)�>�/n��(Ͼ�>��@�>��=�T�>N0�=��B>풸>��7?̳D?��K?d}�>�p�=��>m�>_�,�k�m�Ad得Ч����<Q��?�̆?p۸>7�T<=uA����l>��?ŽMv?CS1?�`?.�>t���Ŀ�62�]�ɾ2:J�h4R��9=����z�>?���=ͩ;�:ʼn��=Q		?e�>��=��>�>=��>o��=<��<��=씾�Ҳ=A4�=�;�<ǀ>.n��β������+��;��$=�)����ϗ���o>ޡ�����=?R�>v'>���>�C�=1����0>_����L��K�=���	LB�"Nd�X~�/�s5��C>	�Y>�ɂ�=(����?�Z>s<@>�=�?�'u?k�>���uվ�3��wbe���R�oֺ=I>f�=���;�{�`�L�M�d�Ѿ.�>$�>�x�>Ztr>А,��=���s=$��Xg4�ɫ�>e����2$��>���q�KE��響�i�YqE?14�����=�e}?��H?Z��?���>s����%ھo�1>��|�+�=����m�Ҕ��I?��&?о�>�!ﾙwD��M��d�߼m4?煒�y�[������d����m~����>������<6�/1��~Ғ�l�H�o[��8��>zBM?�7�?8� ���N��*;��\��&����_�>;ˀ?�2>JS�>g7�>�tT=��p�C�F=�>=K�?�a�?l-�?OB����=�m���L�>y+	?˖?���?�s?��>��t�>#��;� >3�����=�>�q�=S�=�M?Pr
?�
?�z��>�	����� �Rl^�E��<��=%V�>�N�>R�r>���=�hg=D��=\>%ܞ>a �>&�d>��>�9�>�f�������&?}M�='��>162?�d�>�Y=�2����<�PJ�H??�kA+�)����t��<�h��h�P=��̼P8�>?�ǿ�-�?��S>$��G?�[���1���S>?0U>�޽���>?�E>Am}>%z�>f&�>�V>�q�>�'>lFӾ��>B��Hd!�<.C���R��ѾMpz>(���a&����~��]FI�q���g��j�n.��_:=�<�<�H�?�����k���)�	����?/X�>|6?vڌ�����>���>�ƍ>TM�����xȍ��j�w�?���?q?c>��>��W?I�?l�1�3�gwZ�g�u��(A��e�z�`�����V���%�
�����_?(�x?�xA?�?�<�Cz>���?O�%�5Ώ�5*�>3/�/';� <=q&�>/����`���ӾW�þ!�YUF>��o?|%�?fZ?0dV����vKU>��>?�3?j��?�&?�`?�ɕ�2�?=�.>%*�>b�? �?�3?���>~8>@1X=��4��=����S���&�1�S�+������9g:�;5�9��b<�(�=
�<�'@�����:�
<�D=��=] �=&�=�c�=d�>�]?l��>#�>ص7?C�z�7������.?��0=�q��5틾"������}� >��j?{��?n�Z?φe>��B�+�A���>V�>��$>�K\>m��>��9�D���=#&>�>;��=��Q����={
�cY����<�� >�E?�?�>�����>JU����n�kl`><�<�����V�OC���3�����"�>�K?R9?߄->������N��d�ʈ.?�BE?ufe?Źc?ٗ����ɳ;�A�c��o��Н>3���g	�����U����?�t�=Q��>�W��砾�Ub>��F޾��n���I���ӑL=_w��U=@���վd:��=
>ڨ��� �s	��wЪ��?J?��k=tO��
mU��s���>(��>�>qD;���v�&�@��������=	��>��:>䫚�����mG��/�T'�>T'D?�k_?�}�?K܅�#�r���C������ѡ�c?��d:?�_�>��?��B>b�=�������d��fG���>o)�>z��/H�[鞾���P�$�7'�>h?�� >5�?�T?�?$`?J�)?<<?�؎>������B&?��?T�=�Խ��T�� 9�XF�q��>��)?ֶB�x��>c�?��?��&?��Q?ص?R�>� �:C@����>7Y�>��W��b����_>��J?���>l=Y?�ԃ?��=>D�5��颾�թ�HU�=V>��2?6#?!�?���>g��>鬡���=���>c?�0�?��o?���=L�?I82>��>���=���>���>�?dXO?k�s?_�J?_��>���<�6�� 9���Fs�x�O����;{�H< �y=ɓ��4t��O����<��;�w��`�������D�x���2��;s�>X3�>����˶�=����<e��1h>�]�� �����4����L���>v�,?}��>_��=�=�e�><��>.�&��u(?�x.?@'?�%���C�ϭ
���PH>�)?�C�=�5c�����x���>�ڃ?ڥV?�b�+ξ�b?�x[?h�U�<�f�ľ�h�D��I�O?�
?��>�Y�>I?�do?�L�>�Db��ll�z✿97b���_�mq�=	��>q���b���>�R8?�v�>d�c>4��=�~۾}�w�Ξ�|?�M�?�=�?��?.�/>�pn�d߿�|����k�-�N?: �>_p���?������d��C0��Un�@d��U���*����#��{ ��w��9��DO���O?��?ܲe?�� ?D��Yr �2U����D�s�������[��B�j6��G��J����gE�����=�r�>��W�?C�#?�PH�IO�>�����H�JF˾�oE>>����!�pđ=�i��
"=��E=�8Z��#�����'�!?J��>�>��4?J�[�2�A�v1�nH3��	��78>UA�>5S�>���>��<-����ԽB�ľ^���[�o8v>Hxc?H�K?�n?r�X+1������!��/��a����B>�k>պ�>îW�w��:&��Y>�)�r�c��&w��=�	���~=�2?�(�>'��>�O�?�?�{	��k��vkx���1����<�0�>0 i?YA�>p�>6н�� ��P�>Dsr?�|�>[�>�������� u�eVŽ�n�>�u�>K��>��K>+-��$]�/������O�7�61�=^Cj?�=��F^�~�>�I?A�"�s��4v�>2�T� ��ڵྼ@(�~�>��?hڼ=0>rӾ i��R�����Q)?4A?ޒ�i�*�U�}>	"?	j�>/�>0�?
B�>�Fþ�)+���?��^?�=J?DA?�!�>W�=�k���UȽ��&��$,=N|�>��Z>��l=yX�=���~\������D=jr�=&ϼr@��E<C���[K<�'�<n4>JTӿ��>��mƾ$�޾���w��𔎾�d����^��s�޲�v����zm�Y{+�S"&<N�)�-`��H����n����?��?)	`�E ��H䒿X�h����߀^>�������Ͳ�QwD�����?�þ�q�����%78���Y���d�b�'?t���h�ǿ����<ܾ� ?V@ ?]�y?����"��8�ϱ >XC�<�/����X�����ο�����^?���>4�G.�����>�>R�X>�Kq>���~枾�i�<{�?��-?M��>��r�u�ɿI������<���?
�@�xO?����Y�����f	?�"?s%�=��=$�����N��>zɤ?ϋ�?U�ż��:�'�>2�V?\4�Q<�v����S>Kg �t���=���>^��>��i�KO=0�����}�=#��>�t>L!����{��&�>��>�9��2Մ?{\�pf���/��T��U>��T?�*�>�9�=}�,?[7H�\}Ͽ��\��*a?�0�?���?#�(?ۿ� ٚ>��ܾ��M?qD6?���>�d&���t�M��=�;�r���`���&V���= ��>��>��,��g�O�.K�����=����;ƿz�$���$ =�w_�[�����ݤ��JV�eß�<�l�LT罯D[=��=�Q>,�>�U>[�W>H�W?�@l?�j�>L>�潯,��N�Ͼ�G������O��ŋ��U�ӕ��V뾉޾I��������h�ɾI�<�v�=�R������� ��b�R�F���.?��$>v�ʾ�M��<:<�7ʾ���W&��x���.̾ǝ1���m�Թ�?��A?H��(�V�'��<��԰��*�W?Kc�w���e�����=�A��Ji=I�>��=��y3��TS�0�0?�J?]X������%>&���=��+?�'?�8�<���>��$?=;-���޽�<\>W^.>�Ơ>��>�>������׽ӎ?�U?I���Y;��Rn�>�K��7�x�c=�!>r�6�\�B�]>��<I���ݽq���F�<{1T?)��=xA����|&ǾDw�����q?v�?�?���?;FF?J4�pa���q#��� �����'?�,z?�
>$��]����ǽdNh?uKj?���>��������K��/�>��\?W�>	�=dlC�h}b������s?��v?s^�us�����>�V�k=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�%Þ?��@���?M�;<��U��=�;?h\�>�O��>ƾ�z������j�q=�"�>	���~ev����R,�`�8?ܠ�?���>������֡�=�֕��Z�?@�?y����wg<���El��m��v�<�ǫ=���G"������7���ƾo�
�'���Fɿ�줆>�Y@�O��(�>FE8��5�TϿ���Zо�Oq���?܀�>\�Ƚ�����j�Qu�4�G���H�Ĥ�����>��<y��=�8˾�茿��6������u�>
淼
ǥ>;�3�)�W�3�7���=�fg>i/�>Q�>	���Ӿ;��?3)��ӿF���l���?�>�ր?�h?
�?��=�>;3=>�*Q>�7?��e?t�D?dJ�ː��ɻ#�W�j?�d���P`��4��ME�\�T>�3?�>�>%�-��V}=%C>̏�>[>� /�r�Ŀ�׶�����-��?���?�k�}��>��?Du+?�c��4��lH��:�*�x���CA?2>������!��)=�wȒ���
?�t0?�W�'�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�E�>���?n/�=rM�>1��=\F���^4��o#>�H�=�Y:���?^�M?x��>�E�=�o8�&/�x�F��+R�����C���>K�a?�^L?Kb>�1��Ȇ3��!�=�ͽo�1�Q���?�p-���߽5>��>>�>��E���Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ta~����7�G��=��7?�0�(�z>���>��=�nv�ܻ��T�s����>�B�?�{�?��> �l?��o�R�B���1=DM�>Мk?�s?Ro���f�B>��? ������L��f?
�
@~u@\�^?)�t׿_��2����ƾ�4�=���<�$>��6�=Y�=��������>sU�>��>I�>�hQ>�v2>e�>]���>C!���������g!���{����"�|���倾%��7C������򪢽�������3�{��c����=�`W?�@Q?�r?s?�7�ǫ">���� <c�(���=I�v>b�+?h�L?��,?k7�=Y����:b��:������W��B��>��X>���>*-�>�5�>�!�;8�@>�7>�Q�>�->��
=�l(�#f=(rH>6o�>�Z�> o�>F<>>�>�δ��1��͜h��w��&̽� �?���O�J�q0���5��z����g�=�a.?�|>����>пe����1H?�����)�C�+� �>��0?�cW?��>���~�T�n?>e��k�j�5\>�) ��~l��)�=&Q>�l?̼f>u>��3�e8���P�#}���h|>�36?�涾bB9���u��H��aݾ7EM>Pľ>3D�-l�>�����Pui��{=�w:?��?�6���᰾��u��B��(PR>=\>�d=�g�=�TM>hfc���ƽ�H��b.= ��=��^>��?��M=.14>�Ԇ>����eپ
�>R$W>P��>��?Q�a?(�_=Uԏ��(��� ֞;��6=��{>H��>�@d�H�=B��>qD�>�A<�8p�x�!�8��>12�)�̛�<�p�(�R;��>!�I>��	�U��ZK>�~?���-䈿 �zd���lD?n+?�=�F<��"�? ���H��=�?t�@m�?��	���V�I�?�@�?���5��=}�>G׫>�ξj�L���?G ƽlǢ�Д	��(#�JS�?��?��/�+ʋ��l�I6>�^%?��Ӿ�k�>���X�����v�u��G#=��>�9H?�I���UO���=�[y
?�
?�T������ȿ|v���>�?�?��m�C��L@���>���?vdY?wi>(p۾�fZ���>��@?8
R?U�>/4��}'�K�?2ڶ?ܫ�?�O>�^�?��?���>̕���!���`��t�=�����Z^>�r�=[n��&�H�x���b��?1j�R8��7�>���<�5�>u!������T�=��������E<���>X�>��@>���>7 �>Nf�>�~�>�&�_E㽊���=����K?���?+���2n��O�<���=�^��&?zI4?�l[���Ͼ�ը>ߺ\?n?�[?d�>2��H>��@迿<~�����<��K><4�>�H�>�$���FK>��Ծ5D�Yp�> З>����?ھ�,��<O��JB�>�e!?���>�Ү=�$?�(�>n~>��>�|g�e�����Z�Fŭ>�y?V+D?v��?K�'?���N
�+0o��[��ˍt��C�=�!�?`r�>�w/>����C�����=Kl.��H�s��?8�N?7�1�j$
?ՠS?�P?�&?��T>=������5��z�|>��!?1���0A��&&����?��?���>�鏽[нo����M�j����?\?V�%?��a�����?�<��.�����?��;��=�8�>W�>kƆ�]C�=��>2��=�;l���5��`<P�=��>�K�=��7�X��2<,?��E��΃���=(�r�/pD���>�DL>z��V�^?z{=�"�{�����x��&U�N��?=��?Hk�?�a�h�#"=?>�?�?��>>M����޾���e3w��ex�@x���>E��>>l�I�i���ԛ��5H����Ž���_?az�>�9
?@��>��>|٭>���1��_T���e����;��C�C�'��\��:�� �<aT¾��q�Р�>9͟>JT�>��#>��>�X�>C�>=��>�|O>�p�>�v�>�9>n�=��<�c��Vs����X?dh����H�,�6�"��7?i.z?��?��!�o����$r�>�_�?Vʷ?��b>�>��㾆�?��>����S�>�@c=78>�ϼ�5徎xܽmj���F����=�����
>�RDg�f���SO? �%?�Q�<�s�HR[>�J��M�=[{�?E�!?d-*��nD�v�n���`�6�V������s�kȱ�w%��jp�����m��+�z�y��Gѻ�6?ƽ�?B��r��k�����Y�o�=���\>d?�>���>�f�>�T>��
��
.�O�`�gO'���W��+�>
�w?J��>k�K?�;?�_T?�4M?߱�>�ܫ>񱽾�R�>�,���Ϟ>B[�>A�1?��-?l�2?�?��-?sf>��Q���D�Ѿiv?��?��?Q=?��?o|���ν͇�'f����i�������D=�÷<Ľֽ� b�C��=�O>�i?�����8�W��w�j>#N7?���>?�>)���=����Y�<���>��
?�ҏ>����	�r��L��{�> ��?]�/="�)>�>�=,�������)S�=.�¼q�=�y�� �;�F�<j˽=�=q&��	���f:��;9�<��>;Z?���>��>�6ͽF���`�+����;76Q�װM�n#��	�LP����T߁��Έ>ʓ?��?��=(yh=v\�=}7�9��(�V�ǫҾ�J���?.a?�l_?��4?P��>7#*?�A�=�L����s}�����$�(?/$,?/L�>(��U�ʾ���]�3�>h?�L?Ma�k����(��@¾jAս�>D/�(~���D� w����#N����?¼�?_@�.�6���F���h	��жC?�F�>��>���>f�)��g�g2�!�:>���>R?7�>�K?�-z?��V?&E:>4�;��ͭ�{���J�;�:>ܛE?3��?LH�?S]w?��>�w>7�B�⾋^�5�6��� �[��X=�W>�7�><��>�d�>�@�=ѽ�*��c�5�&��=��[>��>0��>���>��l>�׽<��G?_�>Ƅ����pࣾ�X����U�10u?Ϗ?1N,?�:3=���/E�������>M�?K��?��'??�J�>�=��ͼ����;m���>��>D�>� �=� "=xz>ԡ�>;8�>T�	���+%7�^-��9?9�C?Ju�=�Ϻ�b!i�g޾�zk=���=�ݼ��KF<��>�z>l+�٘��'�=�!˽��ž�IԽ`�F����s��?���>[Ӟ=��=�+>�����'b����B3l��mj=�2< b�=����j꼩;k=Yũ=Z!���44<	JȽ|;n�{?p�G?�*?�C?�7w>/�>�%'�?�>�����E?�NW>PK��:��#/:�Q���ۂ��+hپ��վ6c�]����	>�H�p�>�5>�u�=P�|<���=��u=0@�=�>/�D�=��=�s�=s�=1l�=�>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�i7>��>"�R�}1�s�\���b��pZ�0�!?�(;��*̾�9�>�o�=H߾�ƾC�.=ς6>�Ba=R���<\���=�	{���;=*l=�݉>�D>έ�=-��á�=�J=���=ղO>Ty���P8�]�+��	4=���=!�b>k�%>%��>�?ɋ6?fJn?Rj�>&��⡾�C׾�R3>@�A=!k�>��=B� >��>��:?�E?��Q?�q�>�%
=BO�>�p�>�� ��h���Ͼ,<��B��=�	�?�i�?$8�>݊������*yF����?̸-?�Y?i�>�Y��EǿG9�$�پ��;=վ�C�=�1=4�>��
�m+-��,���>Y %>�E�>3�>pA�=�7�=,�H>@.�>��=o"���Y>~�*�U���=wH�=|�,=�����KG�,�=��<���='��=���,�@�Y�ػ���=���>?N>���>���=�곾uL/>1ؖ���L�u��=�B���2B�%8d��;~���.�&>6���B>�6X>Qʄ�{1��8�?(�Y>�?>��?�?u?� >��վ�M���#e��5S����=��>W�<��v;�%Q`���M��|Ҿ+��>Z�>�ߢ>�(f>$--�&@�k�b=�R�D%3�m��>�Æ��;��B�P�o�,O���ܟ��i��$�A�D?9�����=��}?^J?3��?�[�>&Ë��8վ213>�G}�v�=��[�v��{���?�D%?��>���gC�6�ƾ����?��>�;F�b�O����
{1��%�>����>�����Uپ��3�����Ր�x=A�J�f�mZ�>Y`F?��?�\�:�x�0O�(��e�T�/(�>$�c?]��>D	?�?�Ƚ����~����=��g?(D�?0�?f�>�=�=�܆����>I�?b��?�ǔ?��?Q�d���>-�a�7�>Ǿ��T=��=R:�=�>�8?C?�H?Q����h��4��qo�AZ�<���=�r�>�ۗ>�Z>���=�=���=lf>g[>|O�>Ǝr>깭>��>(f�
��ȈG?U�=�r�=\�*?��=��½#����;�p$�f,˾t���/H�E+���m���U�=�?->�b�B
?��ѿ���?�L�=�"!��I�>7����>a6�>�1�>~2��<�>��{>0��>�i�>D�>��J>�pN>�uB>�uƾZ+�=�w
�l�&�I�"?W�Ci��ij>����S�������Rx;� ��|G�<Od�������=��a�<�??� ��g���%�����?f�>��7?��x��:���@>G"�>�d>0&��L���^��RTﾱ��?�?Vc>{p�>(W?�?�B2����sX�9y��4D�r.f��"_��F��^M��%N�`�qVZ?�Iw?�	C?�1I�%r�>-�|?��������>i)���9�w.\=F��>�A����c�ygؾF�¾���.>�i?Ѽ�?)?tWF��-p���&>�:?��1?�4t?��1?��;?v.��$?P3>�)?�n?f?5?�.?4�
?g�1>��=k����(=����㊾�1ѽVDʽ%�\�4=j�{=�ud��%	<�=�k�<j�Lhڼ�;�꡼���<!f:=4�=���=�۫>ͭw?H|?3a ?�U?/4�=k�پ������>��㽊�Q��ǾI{��EǾ �>d?-ƫ?�e?�U=��`��u9W>:v�>`0�>���>3?4^�=»,�}$N���>8�{>TU�=o�������i_B���p>�FK>*k?#��>ᩣ=�Ug>U�FRK�s @>4��dm��򦾍�<�+�\�D�����?��w?J=K?�=z>������j���]���*?pw/?wg?��j?�v>�����L�q�U�/4q�>3X���!,����{�������X>��=><�,����s>z�e}ԾRV|�tjI�E��m:P7��=pt�����兾"�=�(�=/?Ҿ�,��똿�T���DE?Me:���8�o�������e>���>L�>\�1�-����C�������=���>�Q>'�;�K߾�uC�(�	���>�]E?�f_?�U�?�p����r��qB�Tk�������齼��?[Y�>,<?�@A>���=�𱾯@�Le���F����>��>d����G�����W�󾡶$�`h�>�:?�] >X�?D�R?��
?ä`?+�)?�S?�J�>�̶�[���C&?ׅ�?kф=_�Խ_�T���8�nF�T�>	|)?+�B�켗>�?B�?o�&?r�Q?�?��>.� �;H@�%��>�X�>��W��a����_>�J?���>=Y?�ԃ?��=>�5�梾�ة��C�=�>p�2?E1#?��?���>���>��C��= ��>�
c?E0�?��o?�~�=��?�52>��>g��=���>�>k?�XO?��s?b�J?��>���<,2���/���2s�X�O�Nw�;ȿH<��y=���2(t�WK�=��<�@�;�~��Pj��O��!�D��쐼'�;���>��m>���ْ�=ו�=�1�
�>_�0��qm��H]���h���f<�:x>`�?�N�>@��t9=7��>��>����D#?S�>�?���<ÐU���|���qڞ>��K?�>��e�e������(�=�|?V�\?�T��8��A�b?G�]?sh�j=�t�þD�b�����O?��
?��G���>�~?W�q?Ӻ�>��e��9n�J��yBb�\�j��ζ=�q�>�W� �d��?�>;�7?�Q�>��b>�'�=t۾ �w�q��M?��?�?���?^(*>T�n��3���#��`��G�M?��?�֭�9��>��/>�����`����^���+���������O������ZX�9���."=��?B�?�n?Ɨ?/���n��v��H���
C��+��Cl3��[R�hOM��KJ��2p�B�%�j��-������=:�N�7��?"?��#��7�>wf�K��ժ�rTI=$���t�<�
>,�<L@>�'�=��ݽ-��<��̾�??�:>��T>��Q?��@�e�R�������a�վ�Ch=���>^�?��V?��>�����1$���������������_>?Wb?٩I?�3j?(
-�5�1������u$��u8���.>%5�=om�>/Y��j3�O&)�8\C�cv�pI
���� �&�b=��*?Iɋ>��>�?�{?�b��,�������8.��]�<�۹>�Bh?M��>�>�޽\#���>tP�?��?�>G�ʾ=�F�+��4�3��>4P�>\��>�;Tр��r�� �������.���ܮw?�G��`;`�%�S>�2-?25��N���;^�>.]�jz��*���-W=د>���>�8>2�=�]��-�� �\��Q*?��	?���@�4�7�>�3?���>�t�>vM�?�t�>i^̾�!��I?n�Z? �\?FK?��>��=%�B����L�	�u��<v4�>��E>�J=ڮ=S�%�
~]�86)����= �=$ײ���6���<&{f=��u=��t;o�>�ܿ�LL�ҮӾ����,�tz��u�ą������:L�������Ǖ�zRy�C��'�-��J���d��Ց�1�d�J>�?u��?L|�2}p�P��Xy����O<�>�u�w,i���_�L���^�ھ\�����!���K��3_��g\�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >_C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾r1�<��?7�-?��>Ŏr�1�ɿc���y¤<���?0�@��K?��5�zY���A�;\��>�lļ��
�J��=ge�a�;���I?�ǰ?�I�?n��>��-b���7\?�T\=H��o뽨�e=}s�e�Z�&��;�:;>��>�*�=�'D�v|H�QP���#>U{��R��}�'��j=uj>�:M�D&E<μ�?n�[���f�z 0��0��>h�S?���>��=;J,?p�G�@ϿY�\��x`?�L�?���?�(? ���8��>��ܾe]M?H�5? E�>c&���t�34�=�9ؼ&Ȼ��侤CU���=��>�> I.�x����J��P���
�=�v��#ƿ�H%�Ȯ��6=���	�L���׽�Ē�e�G�E_��'*h�����xg=�^�=*JU>ۂ>q�J>n{Y>��Z?$;g?؀�>��(>�#�p`���^Ǿ|�ܻ� ���P�����_�|��ON�;v޾0����/!���ɾr<=�O�=��Q�bk���� �+�b��{F���.?O�$>8zʾ��M���<wiʾ����Ɍ������̾��1�k�m�캟?CBA?���e�V��w������M��X?p��]��4���:�=[��ۤ=HW�>�٣=�7⾴�2���S���/?�&?q�վo����\>'}��W"�=n�?��>���%�>�?*&����s���Z>���>f��>�� ?�>��;�AN���)?9�U?K��F:��eX�>�}��,��J/�=��=~�#����;���=�6��t%��,��<M�<r�=�0W?��>�*�����j&��<=>�x?�?�"�>g'k?@OC?��<���d�S���
�D_y=[�W?�#h?�>�����оE?���D5?��e?��O>�'g����I/�{��*�?�pn?�M?-z��QK}����3�ܐ6?��v?�^�i^������6V�5�>���>C{�>��9�9�>�[>?�Y#�L��̵��64���?��@��?bE<z�"�:K�=�V?.��>O�jXƾ�����ʹ�7r=�I�>����1v��� �,�<)8?�w�?���>T����k�{j�=�֕��Y�?l�?,�����e<���*!l��r����<���=�S�Á"�`���7�k�ƾ	�
�櫜�p�����>G[@^C轸�>�g8��4�UϿ����Oо�Aq���?�u�>��Ƚ�����j��Ru�\�G���H������>.�>hL��N��MC|��?:�O�����>5�	��z�>Y�X��t��􈟾�b$<o��>#�>0߂>�(��_��i_�?\F��]Ϳ�	�����Y?�|�?�?�r?�{�;m�z�7�v�A���`�F?H�s?�Y?�-���X��UF�$�j?�_��vU`��4�oHE��U>�"3?�B�>T�-�&�|=�>���>�f>�#/�v�Ŀ�ٶ�,���[��?��?�o���>q��?us+?�i�8���[����*��+��<A?�2>���C�!�B0=�[Ғ���
?U~0?{�a.�N�_?�a���p�|�-���ƽ�ۡ>��0�Kf\��Q��z���Xe�����@y����?<^�?W�?a��� #�56%?s�>�����8Ǿ�<���>Q(�>�)N>�H_�s�u>����:�4j	>���?�~�?Ij?�����2V>��}?���>��?���=v�>���=��C�#��##>�n�=��;��?�rM?\�>��=��9� ?/��wF�bdR�D��ƱC�f��>�a?�DL?)mb>�¸���1��� ���̽��0����Ԯ?�b+��z޽��4>�&>>��>K�D��"Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Oa~����7���=��7?�0�"�z>���>��=�nv�ѻ��7�s����>�B�?�{�?���>H�l?��o�A�B���1='M�>��k?�s?%fo�w�ձB>��?ױ������K��f?�
@zu@}�^?�hֿ�����M��l���y��=��=��2>%�ٽ7^�=��7=\�8��9��]��=��>��d>�q>J'O>�`;>l�)>�����!��q��&�����C�����
�Z�����Xv�Lz��3��/����@��4ýIy��FQ��1&��A`�P��=��U?�R?�p?�� ?*�x���>
����,=K#��Մ=2�>�i2?p�L?��*?f̓=䧝�$�d��`��oA���ȇ�$��>�mI>���>�J�>6(�>6�b9
�I>_2?>��>� >k'=��U=��N>M�>u��>�w�>fB<>�>�δ��1����h��
w�`̽�?N����J��1��:��ꦷ�fh�=�a.?�z>���?п1����2H?%���	)���+�N�>��0?~cW?Q�>h����T�'9>����j�`>�* �~l�.�)��%Q>�k?ٿf>�u>Z�3�<d8�t�P�|���d|>T26?綾F9���u���H�odݾ�?M>���>�#D�wj�����q�Gyi��{=�x:?/�?6��WాѰu��@���RR>�7\>4Q=g�=�XM>�\c���ƽ�H��S.=���=�^>z?��E>5i�=i��>m���1N�ſ�>��;>�t(>19?4�?�?J�:�ƽOё���4��z>���>���>'�>7�`�<0�=�h�>VUp>" �⮗�}=���/�Za>Y�1�MKZ���w��2�=Mj�����=^T=���"v=���9=�~?���䈿��pd���lD?#+?���=��F<��"�: ��sH��:�?k�@m�?��	�ʢV�B�?�@�?�
��з�=�|�>׫>�ξ=�L�ձ?�Ž2Ǣ���	�q(#�bS�?��?K�/�Pʋ�l�j6>�^%?*�Ӿh�>6x�iZ�������u�	�#=��>�8H?�V��0�O��>��v
?�?�^�۩����ȿC|v�]��>=�?���?��m�nA���@���>D��?~gY?^pi>�g۾M`Z�h��>��@?�R?��>�9��'���?�޶?���?I�=
G�?��u?�L�>�_���L(�#늿Aq�>f�=Ƚ,>dc�>2�.=9����D��%���?��� ��W)A��d�>Ӣ	=,:><�g ��o5>�a�<����|hV=4A�>,�>�D�=:'�>�l�>��>#yp>�>3��U	>�G��f�K?q��?���[4n�t��<Ȝ=p�^�#?K4?S�Z���Ͼ�ͨ>�\?���?�[?�j�>8���<���忿��і<G�K>�2�>VE�>8'��nDK>m�Ծ�4D�?l�>�җ>5���fDھ�5���K���H�>�f!?#��>"��=w� ?��#?��j>�*�>[bE��6��`�E�-��>c��>�L?�~?��?Oҹ��Z3�q��V桿�[�8N>�x?wR?���>S���M�����C��-I����E��?�rg?m#�R ?h2�?��??��A?/f>Nn�f�׾�����ր>�%?=����X���@��HY=�8?���>ǌ>�=&?<�׽�a1�����]?#ń?XKC?�9��OgK����E��D�Q=�zb�F|�<J�2��~�=.�=a������=C��=�~:>��Ͻס��Ed���=	�>�d^>
w[��a �}�$?��">�2s�	i�=��3�:.�$׭>��V>z����8?����k�
��N ������Ո?P�?�?̅<Pk��,?m`�?�?T�>M¾p��a���Z_�G�4������==)�>�f����羽
��J���}�����}�i�����#?���>T1?�8�>L��=a.�>:N������?Ӿ���oMX������U�ã2�l�א�H&Q���>Ƽ�yWz����>�Q��Wm>��>�(>b^h>�>� }=̦>��6>2v�>g��>K�8>��[=�r�Ƃ
=n*߽R�S?Y����Y��8?��但eq?�'K?1e.?�>m����\;����>�"�?駣?�{�>XG�"@(��5M?��>(����?T������M�>m�5=m��j�����>��>z[{����o�V罗�b?��?�s�ڡ¾�d�>��ʾ�x�=!�?�'?�oQ�}b�2Cd�gC���L�F~O=��v�!RɾB�*�N�]�쟐�pm���	��7*��Y�=l�2?��?CP��<��F�s�Y���T�m��=@5?��>���>�>5���Z0�?�\���/�m.޾��>b]w?���>8�I?^<?�vP?PhL?���>Z_�>2���p�>$��;���>^��>М9?��-?�20?�v?�s+?D9c>=h�����L�ؾa?��?&G?I?�?݅�[cýؗ�$hf���y��l��4�=��<a�׽9ku�C�T=�T>��?	��x�7����,�a>��-?��>��>��������h*=a��>��?۝>ҽ���1q������>�9x?Pe�f�=�P)>@��=���<k�>��;���=��M�(�A�p�<R�=�H�=�*�
�׻n9���;�22:]�>� ?"
�>PɆ>v8�������}	�"��=��T>�#H>��>Z�ھ$����m����e��7}>A�?h��?�΂=���=���=*薾�t�����ƅ��_l=U�?�!?�T?��?��:?#?� >V.�&m���ჿ����;%?t!,?��>�����ʾ��ԉ3�ٝ?e[?�<a����;)��¾�Խ��>�[/�f/~����:D�c녻���Y��4��?뿝?aA�T�6��x�׿���[��z�C?"�>Y�>��>P�)�z�g�r%��1;>���>hR?D�>��=?�Tx?-�T?o�?>�7�6����Z����L�<W>�	@?�<�?��?�|?*]�>�k>9��=��� �A@�=��k=f=Q>���>c��>�4�>��=*�u���v���,�У	>�^> ��>Oݒ>k��>r�e>}��~iF?
	�>�y�M\)�Oa��v��<��>�9?l��?2w�>�;�7�]dQ�N����?���?c��?ߘ
?Q ���=�<�q��ǽ]w�>���=��>׾=ｍ�'��m�>s4�>���E�*��KV�r�<��A4?T	2?��ξҿ6�� m�^��<\ @=�S��ع=%YJ>
����eS>�Bu�<1i�4�z��Z���xX�z�����ל��5�5�,�?�S�;�#M>�Dh>n�K�����5_W=/4Ҽ��P�AS��a��XJ��ý¢G=�U1��<>W�={�o=�⬽�M��K�{?�N?�''?#2?��W>�c6>��d��/�>�t=�>?�.`>Ӏ\�������|�'X���⭾ D뾽����zW��^����=����M�7>;k#>���=3�;���=7�=���<BR-=eV=x>��=���=>�>�>3�=�6w?X�������4Q��Z罦�:?�8�>c{�=��ƾq@?}�>>�2������xb��-?���?�T�?>�?>ti��d�>M���㎽�q�=J����=2>o��=y�2�S��>��J>���K��H����4�?��@��??�ዿТϿ5a/>@�U>,?�=|<P��`-��S�����e���!?�8>�ыо���>�/>J���Q���`�=V�>PL�=O��j�b��=�T[�!i=���<�>��W>��>�q��=�K=��=MNH>��+<=84���\�{�)=J��=*b>���=���>E�?�a0?�Pd?�-�>	n��Ͼ�4���4�>�0�=�X�>�<�=�B>���>��7?q�D?��K?Ƌ�>�5�=� �>
�>Ѣ,��m�lX��ԧ����<���?�Ɔ?/ڸ>�U<A�.���i>�L`Ž�v?sY1?�W?�מ>R��۟߿�&� �)���d�� %���N=^D\�[m
����Y��ҳѽ�>�="b�>���>�>�gj>��(>�O>V�>F�>v�=5)�=�[r���<�T���i=���޴<���1ۻ�0�[�V{���]<}��;þ0<�D�R��=N�>�>¢�>��=wų��\'>����b�E��4�=[����XA���d�i���I/��&���c>6�N>�q/������� ?��i>��D>ܼ?l?���=Nf�Ŋ������ˠm�2V��,�=�V>X_8�ڜ@���d�*dM��jɾ�t�>qh�>|O�>R�l>��,�-?�js=a�0�4���>
��o&�H���p�=4������ہi��$��+�D?�ᇿt�=,�}?�H?���?�U�>�g��04վ^m/>Uv����=����o�;���z?8'?�J�>%�뾝�D��aʾ`^Ͻ���>9E[�;�H����؝4��ߊ��M��1ص>����^KӾ��3�����֌��P>�L*����>G�C?�6�?i���Hr�LCM�&��������>�Z?�=�>���>D�?��ݼA�پ�bm�3>��t?S��?�o�?��=�̽=� ���#�>`	?��?���?�zs?��?����>0�;�� >���n)�=
�>,�=9o�=�o?(�
?%�
?d���Q�	�������^�^x�<�š=�|�>|f�>^�r>O�=��g=�;�=��[>�מ>F��>��d>}��>�E�>�����ڶ!?+t>�f�=�5?�82>��C>SA��^�=�H���]��bs�˓ͽ��*�t�P��F4����\�r��0R?�0ÿח�?D˕>-6���<.?,����i�=s0���>�f<k �>�E>Aˊ>8'�>���>y�>��? +<WӾ�>����Z!�~=C���R���Ѿ�9z>ƌ����%�h�����TI��j��[o�j�2��LF=��v�<>D�?=��F�k���)�lY�� �?�[�>/6?�ӌ�1��|>0��>Xƍ>a5�� ���3����T��?��?�7c>c
�>��W?��?�1�X�2�xZ��u��&A�x�d�n�`��ۍ�%���
��⿽��_?��x?cvA?��<Xz>���?��%�����>�/��;���;=� �>d9��z�`�%�Ӿ��þ���F>J�o?6'�?�c?QV�*x���>�=��6?�9?�l?rM.?�C?k�߽ח ?�2H>)�
?�	?4�1?��.?�?�E6>E��=E����=���������ʽ��ֽ�o1��=� S=V�c��ᠼJ=�G�<�}��[�Ji:]�����<6�W=b�=���=壹>XZ\?v&�>}�$>K�8?e���� �Iɾt�?J�����󶕾�WݾH��O� >�v?}�?p�T?��T>�*v����X{>�>�ŗ=eM�=�-�>����I���3/�=� >}`>��=���᯺������w�>�WF>�B�>R]�>�*���>����qg��X>�j\�fҴ�b�d�6�E��0�T��_��>�L?M�#?WE�=D�㾧�����d��&?ߩ=?��L?x?�5=81;��7�VO��0"�SC�>�U�<C	��ߡ�WY��<B<�A�8<��>f2�����Cn>_����پ�Uh��6F��~ھP�9=���C�=�
��JҾ��u����=�>\:���d!��Ֆ�7۪��LI?U�=0{��{Mq�\w���%>֖�>%��>򥽲�?���@��`�����=<e�>=/>���&�X�D���]4�>�RE?\Y_?aj�?(���s���B�W����X��s�Ǽ��?_v�>�b?�B>�ݭ=}���l
���d��G��>���>�����G�m1��#1��`�$���>�5?��>4�?��R?`�
?�`?u*?�E?(�>���~�� B&?5��?��=��Խ�T�� 9�JF����>z�)?�B�ṗ>R�?�?��&?
�Q?�?}�>�� ��C@��>Y�>��W��b��G�_>��J?ۚ�>t=Y?�ԃ?w�=>\�5��颾�֩��U�=�>��2?6#?N�?���>5��>����W��=��>c?�0�?c�o?ی�=��?�;2>��>��=̙�>͌�>?XO?��s?��J?6��>���<�0���3���1s��P��&�;�H<��y= ��o@t�8?���<"��;���K����)�D�G ��T��;�`�>��n>7��*>�G���|��8�N>�J���}����rPD����=Zl>�?���>ׄ�8��=k��>�"�>I6��A'?�?��?�Mۼ�gd�]�Ⱦ�#]����>a�;?{�=�k��=��J�u�jP=itl?7`?
J�WZ��I�b?Z�]?mh�/=���þӶb���$�O?��
?T�G���>��~?:�q?��>H�e�p9n���Db���j��Ѷ=Cr�>]X�G�d��@�>�7?kO�>}�b>#�=�u۾�w��q��"??�?��?���?&+*>B�n�4������?��^?���>p#��)�"?}:����Ͼ�Z��$B��+
�C��1��b`��0�����$���)~׽��=Y�?��r?9fq?<�_?m� �M�c��.^�]��7VV��(�i�E�E�}�C���n��U�	��Ƙ�/H=�wa�1�M���?N�?Gv�#��>E��:ܾQ��H=B>���|�ѽ�,>%=��=[x�=��=�qҽ���ľ�LI?��=)@�="P?^�T�F8M�/k.��Z�^����C>���>s[?�!?�.>-	=��ㇽ�Ȓ�Qʨ��a��[�q>e�c?w%L?*jn? �r0��s����!�yv"������B>�C>�!�>�mX�����&�9�>���r�a������'	�U4{=�I1?W�>���>6��?�M?�y	�����{�x��1�\�<��>��h?K��>A�>N�ѽ]�!�d�}>�q{?�?΀�>d$پV��Q�\�@V��^�?�>>/F�>��5=\����zS�ס��@���J�E�s	>'}�?^���OO����>�@?j����,W�T[>0��=��)�s?���t�<��w>���>�X�=9U�=(eξ2�-�󟄿m26�5*?�?����0�e��>��$?�>b��>��?�ݡ>��;{��`�?�Xb?t�W?��>?���>�pd=�X?�����aK	�J�W=���>0<>!d�<���=X����x��9� Ã=F�=��W��b���<���<�D�< �<�k(>]mۿ�BK���پ�
���]?
��爾׫��.d������a��C��"Yx����'� V�8c�B����l����?U=�?1����/��$���,���7���6��>�q�	��/�������(��7��ؿ��d!�`�O��%i�0�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >^C�<-����뾭����οA�����^?���>��/��p��>ߥ�>�X>�Hq>����螾m1�<��?7�-?��>Ŏr�1�ɿc����¤<���?0�@�PN?{W�nx��6���ţ>9��>�n=�Q= �N��wX�6�$?z6�?���?Q�<(%4��Y5>�=?�T��w3K�|�=�XM>ȸ��>��={uG=΋�>�?�F�=4?�=�H�##ٻ�W���=���<5߱���X6�>�k*=9����?]E�`i�<F'���\�g9 >?�a?F��>/<J?c�@�d˿pE\��AV?���?#��?��%?Ē��Pn�>��Ӿ�H?l�G?�'�>tx;���x�K!d>O�*���y�)Ծ��<��m<��>�M^=O'��v>�)R��+=5��=d�B�ƿ�$��|��^=$�ݺ��[�/~�ް���T�X#��&fo����6�h=c��=�Q>?l�>2%W>4Z>gW?��k?�N�>_�>7�n���ξ�w��G�����K�����m��R�ʩ߾{�	���������ɾ��<���=�+R�-���� ���b�m�F���.?$>#�ʾ�M�W�5<Eʾ?⪾�Ń�k䤽�6̾��1�f�m��Ɵ?2�A?������V�������ϸ���W?���¿�z鬾;��=�Ұ�Dz=��>0��=x��3��rS�2O1?��?L�ȾRr����8>�7񽣹^=Fb-?Ӯ�>��L<wޠ>��?�i7�w_½���>սG>��>O��>�o>��%�ƽ�h?��X?�$�ʨ�~��>�Ǿ����B=�>@�g�1���A>�������<��_�&��;^�V?>�?>��+�r�*�g_���w�[��;&j?�?�>P�>ږy?�3Q?1,=wx��/A�X�ؾ��<x8?f�g?��>GZ>��rܾL|���S?��?^׏> ѳ����|4�V�����>1�[?��
?=���p/m��Ɇ��.��&?��v?�r^�ls�����,�V�e=�>\�>���>��9�|k�>��>?$#��G������tY4�%Þ?��@���?��;<� ����=�;?k\�>�O��>ƾj{��������q=}"�> ���aev����JR,�D�8?Π�?���>ؓ��Ʃ����=�ٕ��Z�?�?���IDg<S���l��n��r�<�Ϋ=���E"������7���ƾ��
�����࿼˥�>DZ@�U�v*�>�C8�\6�TϿ(���[о~Sq���?M��>T�Ƚ����@�j��Pu�b�G�3�H�¥���<�>׶.=c+��%�s���:���2]�>q�нr��>w��Á�����ݼ���>��>e�X>2�ڽg�����?�%�T�ʿ�����;�Z?���?z5�?��?�x���
U�:-6��{Z=2�=?c?WR?:���`����%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�e�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�+�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?(�a�P�p���-�O�ƽ�ۡ>��0��e\��M�����Xe����@y����?O^�?f�?ڵ�� #�j6%?�>Y����8Ǿ��<���>�(�>�)N>tH_���u>����:��h	>���?�~�?Rj?���������U>�}?W�>��? ��=��>r�=������@��">n��=��=�
�?eM?f]�>k~�=��9��V/���F��4R�N���C��ڇ>��a?#L?tsb>]R��<�2�Q(!���̽w0�	_�~?��)���޽��5>Ѯ>>
I>�E�4�Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�a��=��7?�0�!�z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B�~�1=9M�>Ϝk?�s?�Po���h�B>��?"������L��f?�
@u@a�^?*��ֿ쎿O蜾�����=� �<�F>0��,j�=���=��:�����=���>�M>��T>�'>) >��.>}�����t����Z����T�	B-��t%����2��^{��X��]e��}Ծ>fԽ3ѽ�˽��\��3F� �P��1=�|Z?�T?�q?��>�}����/>������=��rۊ=���>�+?=�J?.u$?�EV=�׬��Gd�󃂿$Ƞ�hݐ�)�>x1>wZ�>C5�>e�>JZ�<ە>��O>�p>5�=�k=E�W�gv�<�4U>�©>x9�>x��>>i<>tJ>�˴�f4����h���v��3̽���??����J�\�����s�����=^.?U�>���f<пV譿�+H?甾;/��+��~>��0? oW?�
>���1V���>(����j��P>,A �D�l�x)��Q>�\?��f>`u>�3�e8�r�P������[|>�-6?G�09��u�/�H�[ݾMM>T;>�B��h�������si���{=Ht:?C�?R���谾g�u�~E���HR>'$\>�d=�f�=CM>��c���ƽ�
H�,�.=���=��^>��?fP���'>��Ͼ��¾�>���<o+X:�U?&kH?��>IIX=`u�<�!��O�>"��>ѫ�=]D>�F��>�g�>�*�>�-=F*���K�9$��u�>���]�S@�)J��Tb���L�=�=�H
�+�D���>��~?#~���䈿[�vE��zmD?6*?��=��F<�"�����AL��d�?��@�n�?g�	���V�o�?�@�?�	�����=�|�>�ث>�ξ��L���?ƽ2ˢ���	�."#��P�?��?�0�`ȋ��l��8>H\%?P�Ӿ\h�>�x��Z�������u��#=6��>�8H?�V����O��>�w
?�?�^�թ����ȿ3|v����>R�?���?Y�m��A���@�΂�>A��?�gY?�oi>�g۾g`Z����>»@?�R?��>�9�q�'���?�޶?ͯ�?rr�=7$�?��|?>q�>�f5����'���R�w���+>�I�v�>U��= W�_^A������d����x�Ԃ�#��>�$ɼ@ԗ>��i���v�=��_�c{��m��\�>�ߏ>G"Y>�>�c�>B(�>�Э>j��=4cO��.��v�˾��K?���?1���2n��O�<j��=�^��&?�I4?k[���Ͼ�ը>ݺ\?j?�[?d�>:��K>��@迿3~��z��<��K>44�>�H�>,%���FK>��Ծ�4D�Xp�> З>�����?ھ�,���U��LB�>�e!?���>~Ү=ݙ ?�#?P�j>�'�>YaE��9��w�E�ͱ�>#��>[I?y�~?E�?Թ��Z3�}��x桿|�[�k9N>��x?�U?�ɕ>0���ポ�DIE��7I���e��?tg?R�?2�?p�??��A?�)f>r��XؾG����>p''?��"�#kQ�9�?��I<�)?T�>�&�> �H��<+<�Kѽ���c��0?+��?�.&?����(7���@�"E�<o�=� �<� �=�j˽|�;
�->}ŽwU�°E<�
>-v��0��k�^A�=7�>
>��J�5���1,?�XA�׃�77�=��r��`D�a�>8�K>?���m^?��=�P|����`��BfT�;�?���?�h�?$���e�h�)D=?i,�?-?���>~��+�޾��ྚ`v��%y�wu���>���>=z����m���_���$���ŽE�+��p?�]�>	R?:��>�"N>/��>>c��o����ﾣ����Z����T�6�1��� � ����(.�������þq�}��>�3���A�>t�?��U>�Lh>G��>-/�;忎>�'k>m�~>R��>�'`>ڎ:>++�=����v� �0�V?���^�d	�sc>�Tl?s?O�K?��|>\�0�M�2��,�>`"�?=�?�_�>�p�,8���6.?�د>
4n�G�?�׽P:U�O�X=
������v+���P=���>P��^�o�7�[�׽E[e?.A?0��קf���>�Ǥ��p=�+�?�C)?��(��TQ���n���W���R��$���g�塡�c1%��p�A鏿'C�����(���.=��*?V)�?�� ����N���j��?��j>Y��>��>�>ozH>�(	�1���\�b�&��A����>��z?���>L�I?%<??xP?�kL?Z��>�c�>4���l�>T	�;� �>��>�9?H�-?80?�z?1u+?�4c>a~�������ؾ�
?y�?�J?�?߮?Vޅ��rýp���g���y��~��k�=��<��׽�Bu���T=�	T>#c?���o�8��*���j>��6?Oo�>�`�>쏾�?��\�<b �>��
?>���$�q��G����>#��?����M=H�)>S��=����L��=�z¼A�=݄�89�)<'d�=>�=F�B��\�9�S�:�t;Y�<0��>�U7?g�>�1�>ٕ����o��� ʳ�t��>��/�1J�_t�ӏ�n㛿��c�^�>'�?A�?�`�=�X(=��/>�ʚ�ϡ;P�$�I�������f�>:�F?�M?���?��.?M,�>�@A>�w�iL��!ɝ��7����6?�!,?���>�����ʾ9�l�3�O�?q[?k<a�����;)��¾��Խ��>%Z/�.~�*��;D�fԅ����B|����?��?v'A���6��v���3\���C?�!�>�W�>��>l�)���g��$��4;>2��>�R?�>��F?��r?�T?6;>22=�� ��ne��5���?5>��D?Y�?��?2r?�b�>��)>��,��x���ݘ�r��`���X]==�t_>"��>$��>X�>�f�=ؗ½�����,0�F��=Y�J>�a�>�Ң>�j�>�mr>��<N�G?R0�>BB��)r�*r���j��'�5�؝t?��?��*?�p=��4xE�G$����>�\�? O�?��)?�O���=��Ǽ�����m�ѽ�>�O�>���>�=;�;=6.>*�>��>^��C��{8���F�FE?��E?V��=�̿؁b���;���l�^�=�����U�W ｅ�o��M�<�n���� ��ܸ�z�������Þ�a�¾QP����]��D?��.;JC>|��=L?��R��gL�+V>�t�<��B=������ <�J��1;�k�@�+g;�P0=�>L4<��/�鴆?�n?��$?L�>>��=��=�6�y��>�wb�S��>[�!>'ҽaM9�u�*�p,�x���0�Z�C����o�G+Z;�#�ʸ�>���="��>��A�'�#�y�<R4�:��Ի29>XF>߮>�@>n>4�=g����6w?X�������4Q��Z罥�:?�8�>d{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=J����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�l|>�Q���P�%#-����'f�x�����>؂5�Å[����>�>6i�����hn~<�A�>r>V<%Ǘ�|0�p�_=L͋�p�=./�<ʯy>��a>�;�=�'M��'>C\�=;v >�@�>e?����A�CV<J�q<B_�=��@>�oS>��>N�?H_0? Xd?�2�>�n� ϾMA��qG�>j�=$C�>�Ӆ=8iB>t��>��7?/�D?#�K?3��>Mˉ=�>`�>��,�R�m�Ff�§��`�<E��?�͆?ʸ>��Q< �A�֟�ni>�dBŽTu?�R1?$m?�ޞ>�U����9Y&���.�$����4��+=�mr��QU�L���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=#�����<�vż�����u&�:�+�1�����;s��;B�]<_��;��=���>�5>[��>��=���݀/>����L�nQ�=�[��r7B��7d��C~��.���5��C>bjX>���40����?�Z>6�?>�}�?�Bu?٣>�&�2�վ�S��3Se�%1S����=�^>�R=�p;�s<`��M��Ҿv��>b�>5�>��l>�,�?�ףw=�
��Z5���>�w����9�=8q�`?�������i��_׺��D?`E��̎�=�~?�I?�ߏ?��>�)��يؾ�=0>B@����=�C!q��h��(�?�'?{��>��C�D����*꽧�>��[�H=�����'�t)�<Dž���>r����Zо��2�)�������R:�c����E�>f�=?�o�?�~��A�J�3D�+�-��{��z>�{?4�u>f�?��>�4I�p�i��l���z>w�m?Kq�?q��?3i�=�B�=Q���}�>�	?Ɩ?���?(�s?*�=����>\�W;P�>�8��hY�=��>o�=���=ؔ?��
?�_
?z���Q�	���H��o]�|2�<�B�=AU�>t��>��s>A��=hCa=+P�=��\>�k�>�]�>�d>q��>���>)�߾#>ؾ�6?��>֎>�,?���>�Z=�i ��M�=�����1�P����3,�L*ؽ��P;Ґ�t�¼Q���L?�'˿r*�?�E���ܾk�?�ݾHej=L��V>�>"-0�iV�>'�>�~k>ٞ�>�>��;>�&~>�>qvӾ��>=���S!��C�lR� wѾ}Pz>}���s�%�o���b���I��O���`���i��*���C=���<0B�?���Z�k��)�dH��Ǟ?p_�>�#6?l/��7u��|Q>&��>�͍>�M��$���w���~B��?v��?�+b>q��>�NK?К&?���!�r_:��Eo��3/�9ek�N!d�Ȯ���a��7���Dٽ�=h?��?CFK?eh==��A>%�?o��H�Y��>G���?����<ߞ�>�U־LVi�gƮ�J�����g��ʳ=1�Y?�σ?��&?(D���=o�a'>ظ:?]�1?%Ht?d�1?��;?!��^�$?Wu3>j>?�i?�D5?��.?�
?��1>�w�=Ӯ�֛&=q�������ѽ#�ʽ����{4=J+|=o)�8mq<&?=.��<_��ؼx�;�������<HY:=Oâ=d�=�l�>�q^?���>�Q�>�+?�Z��<����þ�&?+[��౾Q����ξ�v�0�J=�p?���?�w?KC.>{S[���潼,G>Bj>�b�=�˙>ΈS>�
��u�����/>�IZ>�W@=r������i���9�=x��=���>�ȉ>�O��~>�ˏ�C�����>��w�M,ľ �I�U�H�V#T��@ľ<&�>�EM?��7?��>�h���=�-Z���D?�zd?�h?DfR?U��=gپ�>���
�%���,?2>x8U�����f瞿g��%����5>���>�s�{���L�b>#y�q	޾��n��J����J=%m�E�X=���־��n�=��	>�#��w"!����٧��&KJ?�'g=�R��NU�"����,>͏�>�T�>y8�^u��@�h�����=���>i�:>6�����u!G���n�>�=E?�u_?R�?�@����r�x�B����SD��#���Ŵ?Kn�>�>?��A>ƈ�=����z���d���F��-�>���>�����G�陞���̛$�G܊>�?MI>��?�R?�'?J�`?��)?c?	�>�J��2s���K&?�i�?;��='9ս�6T���8���E�V�>*L)?�'B�y��>k�?��?)�&?�|Q? �?N+>h� �
m@����>8f�>�W�yw��ˋ`>��J?F�>"Y?��?�=>�w5������u����=q�>��2?�#?c�?L��>���>l���(��=��>ac?�/�?0�o?�}�= �?�>2>���>�==��>E��>-?�YO?Q�s?��J?ē�>ݤ�<�-��`0��@Js��MP�*�;�VH<�y=ګ�Bt��?�B��<�y�;o���Cs��\��Y�D�����<\�;w�>�l>����\�/>U�q�x��>>�>X�=&xJ��H?�ݍ�(�:��M>�+?�l�>}��q�<2��>���>[%��#?�J?��?���Z�	�������>E?H�=�rr�}Ǐ�3�v�
�Z=��~?/�e?F�q�e&�O�b?��]?#h��=�|�þ��b�m�龗�O?��
?2�G�Y�>��~?p�q?��>o�e��9n����/Db���j�VѶ=jr�>tX���d��?�>М7?>O�>��b>�(�=�u۾��w�+q��$?E�?�?���?**>E�n�#4���'��.@?�[�>uF^���?S�=v;H��4'��=}����Ҿaܾ����-���X�9@���st����=-W%?��?�U�?@3P?���e��pq�P����Rc�V�Z6�'U6�!]G�=�P�ߦg������о̤>�S� <A����?D�&?�љ��ϥ>�9 �!��Q� ��:�>�yɾ�tӽ�a�=�>�=�zC>�z/>�Q��ᄽ�_��Y�/?^��=\�	>n6?����\�ڤ���;��ɾx l���>�?��S?�+�>��սK�ýN�m�+�J�}v���t>��c?E*L?n?o.�e0�2m����!��(�Ԑ���XB>��>�*�>
@Y�����,&�v�>��s�`� 菾�
��~|=y�/?��>���>��?>�?�<	�4����y���0�1�<�o�>*9i?�P�>!��>�νfp!�f�>��?1�?]��>������}S�����e�?���>�˭>l�󻇺����t��������F�5��=�$z?B<��S�"���>ZE$?���<�
<Zx>�>���"�}�����2=��>a��>�:�=�;�=+߾j����e��3B���)?x�?8ܖ��[)�uM�> !?0=�>X��>��?Mۜ>��ɾ�3Ļ��?�4`?��L?BM@?���>� =?k���zʽ����H=���>�P>��[=���=%!&�l!_�����7=��=����|Ľ��F<v.�i�<���<+!6>��ڿa�H��}־k���x�+�	�~���a��s����������ء���(��I�b!���U��^d��(��#�g���?���?����(R���U���逿V��J'�>�Xy��p�֌��o�������侏���"�nEQ��wi�B�a�R�'?�����ǿ�����:ܾB! ?�A ?3�y?��B�"���8�T� >`D�<-����뾤�����οL�����^?���>���/��\��>ƥ�>2�X>�Hq>����螾�/�<��?.�-?��>��r�/�ɿ]����¤<���?/�@[,K?W�L��H�T<��>�A�>P��>^D>��P�վ��?D)�?��?/
�>B.#�s
>1Ak?cc��Ɖ�2�~;f�>5����h���=lu�>�L�>�<$>'�>=��Ŭ�<u~>s�D<�mҽԑf��Oo��K>'��`�<��?��I��Qc���"���g��- >��a?�\�>?��=��0?�M��Ϳ�X���^?�q�?{7�?�X$?�#���|�>F޾y�M?7)6?���>�2��Mb�g�=� ڽ�W���bB��+�=J٫>"h'="f^��9�p9Ͻ�W�=Y<]=�7 ����.�'��"����=��t��yq����2���T�$�j�&��>��"��=� >HK><��>4<2>�oC>�aV?ߜv?(f�>):<>F����bl�z�þtػ�lB����2�hj����O�� ��b��޾]���D��р"��N��w=�?�=4R�����ý ���b���F���.?�X$>H�ʾ�M��n/<�_ʾ>���8����å� ̾1�z'n��ʟ?&�A?H���eW����U���H����W?�����謾x��=-���<=M/�>a��=����3��yS�_�0?J?3���	��^->*� ��=M�+?Q�?v�q<z$�>�u$?��*�0gݽ��_>S�4>
�>X��>�w>������ؽ�?,wT?V�?A���֐>n￾�{�k�i=T�>�7���&hY>7�<:튾�//�z�����<p)W?u�>I *�� ��8�����g�>=H�x?��?<�>�uk?u	C?���<	H����S�G�x=˧W? i?Ū>�@���оω���5?�e?k�N>\h�`��+�.�"d�
?��n?�\?����
m}��������n6?��v?s^�ws�����H�V�f=�>�[�>���>��9��k�>�>?�#��G������xY4�&Þ?��@���?��;<
 �]��=�;?m\�>��O��>ƾ�z������(�q=�"�>���~ev����R,�b�8?ܠ�?���>�������d�=�ѕ�TX�?n�?:��	Yf<���l��w���;�<=ӫ=�a�X�"�N����7� �ƾͼ
�㸜��������>5Z@B�罩&�>�n8��5�UϿ���U\о)?q�(�?X��>��Ƚ������j��Ru���G��H�"����N�>6�=����Ր��[e��D:���n�`�?I�ѽ%��> ����j��X�<�ה>?��>U9�>]t-����\
�?)�߾"
˿�0���&پ,Tl?_ٟ?��y?`5?�c��v�X�-������,?}�x?F�Y?�`��m1R�'W�%�j?�_��xU`��4�tHE��U>�"3?�B�>S�-�M�|=�>���>g>�#/�y�Ŀ�ٶ�=���Z��?��?�o���>r��?ts+?�i�8���[����*��+��<A?�2>���H�!�B0=�SҒ���
?V~0?{�f.��_?Ғa��9p�wp-���ȽhQ�>��2�G0]�"� ��m��Ve��Λ��x���?9>�?�?��r�"���$?RR�>�B����Ǿ"\�<�M�>ֵ>�M>�Od���u>z<�kL:���>���?���?~S?�q�����'0>�3}?ө�>�a�?�|�=w1�>���=Ï�� �K���>��=��"�d�?�TM?���>v�=7�?�M/��4G�R��d��C���>a�`?��K?$g>�����C�0�!�S�νe`5������9�O(�e�۽(�1>=�>>�>�uF��wԾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�K	?���N���_~�C��{�6�:��=��7?�2��z>��>��=�nv������s��>�A�?�z�?���>L�l?��o���B�L�1=�M�>0�k?�r?�yp��:�B>.�?3������}H�C!f?�
@Du@֞^?��c�Կ7n���ƾ�y;�� >��<."'>�;��J�>K"�=~�=ŀ��Q�=�{>�M>s<U>h�7>CG�>>�9��:�!�Y��}@����>��t"��{-�RS�K)������B���E���ľ����}b|�`�ڽ��"�!��ҧ�G��=$�U?�R?�p?	� ?B}x��>���OE=Pw#�ʄ=�0�>�g2?��L?a�*?Mѓ=ի��^�d�`���@��Qʇ���>AcI>À�>�I�>&�>gIt9�I>�2?>�~�>�� >hp'=b%��t=��N>�L�>���>�w�>E3=>�o>:���2/��>�g�E"v�sɽ%�?/����~J�ٕ�����ᶾ���=*`.?tq>�ԑ��6пl����G?_����j��@.��>�V1?`�W?�'>���"�^�- >}��Wk�d� > �O�k��)�v�Q>��?��f>�u>�3��e8�W�P��z���j|>�36?Q趾HE9��u�ݱH��aݾoJM>�ľ>�D�Lk�������ui�%�{=9x:?1�?�3���ⰾ�u��B���QR><\>F=�d�=YM>^c���ƽqH�[j.=$��=��^>�[?��+>w{�=|�>�X���bP�皩>�aB>k�+>E@?�%?�j�#旽�m��۝-�Zgw>p`�>�>b>fJ��q�=�k�>S�a>�m���������?�CdW>8�~��B_��u���w=�#���p�=���=�M �\�<��'%=\�~?��fሿ�
� g���gD?�%?9�=�F<�"����rC��a�?��@�l�?�	���V���?�>�?�������= r�>]ի>ξءL�?�?ƽ-Ƣ�C�	�s#��S�?��?	�/��ʋ�Jl�K>>�[%?r�Ӿ>h�>Zx�zZ�������u�6�#=/��>�8H?�V��8�O�H>��v
?�?�^�ܩ����ȿ;|v����>Q�?���?q�m��A���@�~��>=��?�gY?�oi>�g۾'`Z����>̻@?�R?�>�9�[�'���? ߶?ϯ�?�a�=-O�?0
�?��?$�����Ӿ���淍�췀>؊�>ق�>��=����3c���������d��)����>����VM>!~��Ui��>4�>��a;$�f�1(=��G>�OV>s�,>��>��>e/�>��>��> 發	��������K?y��?A���2n��V�<��=Ͳ^��&?�I4?�o[���Ͼ�ը> �\?o?�[?�c�>��4>��*迿~�����<��K>=4�>�H�>%���FK>��ԾR4D�ip�>�ϗ>�����?ھ�,���8��B�>xe!?���>~Ԯ=� ?�#?Ϙj>T)�>�aE��9��[�E�ٰ�>���>2I?��~?�?Pչ��Z3�����桿7�[��7N>��x?V?ɕ>��������E��4I�����W��?6tg?�O彻?2�?ɉ??�A?�(f>A��iؾF���>�>��#?�5���B�� !�z�ýg�?8�?]b�>�)��J��&�w�C�����6K?"pf?X(?ĺ�
�Z�����?�<�6�:��a<�r�<X6��>.>�H��z�p=�,>b��=ͨ���?�G�H�sg�=ܐ�>Æ>v;;�X���:,?�CC�rՃ�t�=u�r��hD���>r�K>����ɒ^?��=���{�z��Is��{�T���?M��?}m�?������h��%=?��??�(�>�*��p�޾f���Zw���x�q���>���>�t��:�φ��y����;���OƽG��z��>C��>#H?U��>�@O>�Ա>߱����&�գ�ބ���^��v��8���.���Ѝ���F#�b���57¾x�{�xI�>��[��>��
?��g>�{>�j�>���x��>�@S>��>�_�>��W>^�4>�p >�<#ZнN�X?�ӄ��1L�}R���Y>��[?��G?��A?���>Mah��sP��~?��?�c�?���>9�[�й羌 "?W��>�&�g��>���<��>m>��	��d�=*��<׹>��>�P��S��u�d�[��NT?z?��u�)��}c�>�n̾��=>�d�?��%?�a2�Àf��nu�T�j��?P���=z̳���_O;�{j�c~��6��6����K����=t�??/�{?�c��Uξ�b ��D�P�C��9l>SK?���>�X�>�w�>�}ʾ�O�oN���/��������>2�^?ȇ�>H�I?!<?xP?�kL?h��>�c�>�3�� m�>��;� �>�>�9?t�-?;80?�z?
u+?V4c>[~������ؾ�
?o�?�J?�?��?�ޅ��týek��g�G�y��~����=�!�<^�׽Du�s�T=a
T>��?��E�9����R-u>:�9?� �>C�>��G�����]<x�> �?���>�W���vr�.��}�>�̀?`j��~=��,>���=�e�Bv�����=�4���P�=�;��8d���;>��=ǣ�=<���aPܺ���;=���>a=?\��>�G�>�o��hձ�#��	氽GS�>V/��XϽB��4����� �c��$�>�*�?5�?�YV>�CX=���=2�|�.�iEJ����;\�E�?z�d?�h?�b�?pr?�q?���=:���䥿�[���-	�Y�.?!,?��>���t�ʾ��ȉ3���?i[?K<a�t���;)��¾T�Խ��>b[/�"/~����D�օ�����~��%��?࿝?�A�I�6��x�뿘�\���C?�!�>�X�>A�>c�)�`�g�%�W2;>���>KR?^�>�0E?�y?��Z?2�C>̾;�OP����������>��;?�Ɓ?���?
}?���>E�>6��o�ؾ����������P����!=��Q>���>���>U��>㥩=%+߽G"~�͂�A��=E�i>�>㎖>7�>Y�d>��ܼ��G?�B�>��ľ�	�������s+J<dh?*��?�<,?��J�����D�������>�|�?�E�?��.?J�)��=
6�;�ӣ�J�y�sf�>�~�>
w�>l�<`��<A�=��>Ƿ�>E�*�I!�i�;�f!���?Y�K?I9�=)ȿ/�s�0��]����=I`��O�Saͼ�BM��:=��g����oq��^�I�D�������Ѯ��+��h=�����>[��=�� >�>�;=�����=�N<=CS:���<�ʈ���:�&�v����;{�Bb�:%<�=�7<<��ƾj��?sT?��?�	;?*M}>�N�=/]��_��>t9�;i:?u�n>�N,��c��j>J�񦧾�A����澿Ծ�vQ��'����=��*)>Ѐ5>�">S�=�V�=�G�=�A%=�,�j�o=gL
>�M�=�4�=wd�=?b>���=�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��B����4�?��@��??�ዿТϿ6a/>��7>E�>	�R���1��z\�4�a���Y��!?�K;�}̾�l�>)2�=��޾�mƾ�g-=��6>ctc=$��:Z\�x��=kz���:=k=J��>�D>��=����-�=��H=<Y�=֞O>/���ǽ6���,���3=F��=l�b>�k&>N��>w�?�Q0?�Nd?�8�>�n���ξ5���9�>�n�=<2�>��=JeB>w��>Y8?p�D?��K?C��>JΉ=���>��>�,���m�5r�A���7]�<���?�ǆ?-��>��R<��A�¡��r>�oMŽ�}?oT1?vp?qΞ>�;��ȿ��B�K��v0�=�d\�n�<p�=��ڻ��.��$L>�f��+�ý�<�>ɵ�>��>	�=�E�>(z�:��>���=|��;�l>��=#4=VH>���=����<<��"=:�O�ʪ���;�<�e=��R<:��<�n���	<���=���>o=>��>ˏ�=���4C/>������L����=ZI��-B��4d�^I~�C/��N6���B>�>X>�u���3����?��Y>�n?>.��?�@u?U�>�!���վ�Q���Be��TS�Cȸ=��>r=�sz;�TY`�>�M��|Ҿ���>�>��>v�l>K,�0?���w=���[5��>�t����+�;q�@��&����i�H�׺%�D?bE�����=1~?�I?��?V��>n/��ۊؾ=20>�L��F�=g��!q�9_��'�?5'?Q��>����D������Y �Y�>B���%ij�ax��I�J��^Tľ�I�>���!�վ��:�#�w�\���4N�PȺ��SU>��=?�}�?	����X5�e(;����f>5��>��i?��>�B�>(�>g��i�����e�/>��~?8R�?��?D�?=�Ͻ=���=,�>�&	?���?���?2�s?�s?�5{�>|��;�� >�֘�UF�=�>Ϝ=�V�=aq?��
?f�
?�s����	����]��)^����<�̡=Is�><b�>��r>���=�Ag=�Z�=�\>�ў>.�>��d>�>�N�>�����d	�E�0?���=�=/>rn.?%Q,>��G=U�^�=�̽�I��\I��ͽ��ݽ�բ<i\Իu=�����O�>U!ȿb�?UJ>����q�	?m�:G���<*>��K>c� �go�>�>���>4G�>	�>��`>�a�>W�=$�Ӿ��>�F������C�/�R���Ӿ��t> F��L�!����9��M���"p�y�j�5���k>����<�e�?���|j��*)����
?�/�>�7?s��P���,>�k�>�a�>G���锿;���Z߾��?	��?�Ie>u_�>klV?d�?�f,��0�}�X��u���?���d�Ja�,��������
�Kw���Mb?G�y?�dB?���<Vcu>h+�?"-#��苾;Ռ>m�,���;��J.=�G�>����!a�"NҾߵ¾an#�)�9>�m?���?ln?$-Z���m�#'>H�:?��1?+Ot?��1?i�;?Y����$?�r3>�E?�q?�M5?��.?\�
?�2>X�=�f����'=�5��{�����ѽ��ʽX���3=6d{=ͦ��A�
<]�=��<���I�ټdK;���10�</:=A�=��=���>Ysf?=�>���>M�>?����7(�cI�k�?j���j��cGѾ%MԾ����#�=t�?��?�Xs?��r>'�_�n��H�F>��>K]�=ߠ�>�T�>_Ľ �Z��p��:9�=X�>��=	�r�@ӾN��i��վ>DZ>��?o
�>C���u2> �R�`�]����>W��G��l�&�ٓU�`�L��ܲ�`ϥ>S�f?�1a?�G[>��4�4Ȗ=n`Z���3?�4H?�'5?��[?^�	>�O��2=��>�����>������>��l���h���U>�)�>I�Ⱦ[ߠ��Vb>���t޾;�n��J�b��oDM=��^[V=��1�վo5�ʣ�=$
>����� ����֪��1J?k�j=?x��%bU�q���>���>�߮>v�:���v�[�@�믬�x5�=���>n�:>�b������~G�B8�m>�>SQE?AW_?k�?"��\s�?�B�����mc���ȼG�?jx�>'h?�B>z��=K�������d��G���>���>h��J�G��;���0��N�$���>U9?�>��?]�R?��
?|�`?�*?HE?&'�>.������B&?4��?��=��Խ�T�� 9�HF����>z�)?'�B�ٹ�>I�?ܽ?��&?�Q?�?��>� ��C@����>�Y�>��W��b��@�_>��J?ᚳ>u=Y?�ԃ?��=>]�5��颾o֩�V�=�>��2?�5#?L�?�>}��>Q�����=8��>nc?�0�?��o?ł�=��?�92>���>9��=Z��>���>�?MXO?M�s?��J?���>鶍<�7���8���Ds��O�wÂ;(zH<p�y=Ș�T3t��J����<��;zj���T��
���D�����!��;_�> �s>m���0>�ľP���@>���M��Bފ��:����=���>@ ?9��>�b#�憒=��>�I�>���3(?�?n?�!;�b���ھ��K��>B?��=F�l�삔�1�u��h=x�m?��^?гW��7����S?�+g?ao�5�@���{�08r�á���[?��>X����-�>2v�?��?W?Y[v�*,v�
;��a�=�(�_=t5�u�e>*���Z��K�>3V!?�B?5�>�g$>�}������}^�����>9t?i�?��?�Ԧ=���QH߿�&�2�����y?k�?jk�
5H?�KнC��V�_��ɺ��i�I�y��g��1s���;�Q\���c�N��?��.�O?OG?��]?��U?�,4��^2��h�U�e���>��rо��^K��P��W�7�\�A*ž�m�����d�<�w��sDD�9W�?MF.?�v�����>Z���9�z˾��>�\�����,��=ֵI���<��=^&k�5�K���[�"?(��>v��>ׇ:?$qV���5��I0���4�գ��B0>'Ś>��>v�>nL�;4J+������Ⱦyv���3v>	yc?��K?��n?k��*1�⅂���!�x�/�ee����B>�q>�>c�W�ɜ��:&��Y>���r�_���x����	�N�~=W�2?�)�>s��>O�?�?�z	�/j��ihx��1����<a0�>�i?4?�>P�>-�Ͻ�� �V��>�l?���>o��>����M!��{���ǽ���>���>ʮ�>Gq>�t*���[�mX������X9����=0i?+Ą���`�ֹ�>O�Q?u�:�CO<F8�>{�w�?�!����${)�0q>�b?%�=�<>��ľ�p��{�g&���)?M?�m����*�:t>��?x��>V�>�W�?���>�KȾ���[?Pg`?]7M?�NC?ai�>b�2=������̽5d.��i+=�K�>�&X>2�z=�A�=���D^�=��q�*=؎�=�d¼�ۯ��;�C����s<��<�_3>Cmۿ�BK�G�پ�+�b?
��爾窲��c�����a��&��4Xx����'�sV�j7c�$���۸l�͇�?�=�?����R0�����5����������>��q������)��i)����r���`d!���O��&i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�|A?|�(����-V=���>��	?0�?>nU1��K�����oQ�>s;�?��?�cM=\�W�G�	�?�e?c�<��F�	$޻��=�9�=�?=���O�J>%V�>0���RA��Aܽ��4>�څ>�s"�Ĭ��^��m�<+�]>��ս�=���i~?TS2��\�d�C��l�iH���u?�?�>�>��8?xrL���п�b��F`?��?�>�?�;$?���}F�>Фʾ�=�>��?�w�>�/���a�>�>Q�=阢=I)��0Q�P�N=G�>��>���a羠���1�0��=��D�ƿ��$����A='���RZ�!��p��i�S������n�5��'i=��=B~Q>gU�>��V>UnZ>`[W?��k?qC�>��>@��vo��cξ+�B3�����������4ף��@�߈߾�t	����z���	ʾ9 =���=�6R�m���r� ���b�<�F�j�.?v$>��ʾ!�M��y-<2rʾU����̈́�ڥ�K,̾��1��!n�͟?��A?�����V����kf�������W?�N���Gꬾn��=!���x�=�&�>C��=)��� 3��}S��w0?jU?�������?�)>4��=_�+?=�?��X<��>�+%?�=+�X=�
�[>��3>
ܣ>���>�F	>����[۽�?�{T?���2(���>�/��]hz�B�a=<�>�\5������[>���<�匾#lW�p��Uݻ<�]P?�,�>,�;��� �o���˽v7�6l�?��>���>��?��D?H�/>�ܥ���d��&�j����Z?9Oz?�װ=�~�=��þ����z>?�H?�:>w��Nb̾�;H�PϾ��=?>�?:*?.��=�v����/���~"L?��v?�r^��r�������V��=�>Z�>���>��9��j�>v�>?�#��G������X4�2Þ?T�@J��?��;<�����=l9?�W�>ԧO��@ƾ�v��d���=�q=D �>󋧾�ev�9���M,���8?���?a��>͔��������=�ٕ��Z�?��?}����Dg<R���l��n��j�<�Ϋ=���E"������7���ƾ��
�����࿼ͥ�>EZ@�U�v*�>�C8�]6�TϿ)���[оSq���?M��>T�Ƚ����A�j��Pu�b�G�3�H�ť���j�>q�>������<�{��K;�t��E��>z��K܈>��S��Z��-���4�(<���>���>���>vw��0ɽ����?}���?οV���/j��_X?n\�?lu�?�i?q4<��v��*|���x9G?��s?Z?f�&��x]� 7�#�j?�_��zU`���4�oHE��U>�"3?�B�>T�-�D�|=�>���>4g>�#/�w�Ŀ�ٶ�I���X��?��?�o���>o��?ns+?�i�8���[����*�+�+��<A?�2>���F�!�>0=�GҒ�¼
?L~0?2{�e.�,�_?-�a���p�M�-���ƽWС>$�0� Q\�I������We�����Ky�r�?^�?��?_����"��4%?w�>Ҡ���6Ǿ�9�<�~�>��>�1N>�"_���u>	�?�:�nb	>��?j}�?�i?�������K>i�}?b�>;@�?��M��>>��6>��x>�>��[>����>�aY?��?)�P>��]1�e-Z�	�w�U�:�E6O�:��=kx?KC?�o'>����8f/��7��ct����,3_:D8�֣+�Ր(�3�>J�*>�r>ܥ���}���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji� 		?>7����D~������5����=�u7?�9�z>�l�>7��=�dv��Ū���s��Ƕ>�<�?t�?�n�>��l?%o�1C���/=t�>�Nk?P~?�!V�S���B>�?8������V�Df?��
@r@)�^?�̢��hֿ����AN��?���g��=A��=؆2>G�ٽG_�=��7=�8�s<��1��=��>��d>q>((O>ja;>��)>���O�!�	r��X���]�C�������Z�;��Xv�Tz��3�������?���3ý�x���Q��1&�K?`����={kW?<�N?z�g?��?�Ĥ�I]>�<����t=$=�B�=�ٗ>�W0?��F?;�#?5=�ϩ��h��#���[���1��:��>VsX>�>"F�>Ik�>Z�D<�@>�9>�!~>�N�=��5=���;��<��C>Pؤ>.f�>m;�>�C<>��>Fϴ��1��k�h��
w�p̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?3�f>�!u>ɜ3�g8���P�Љ���|>�56?�ն��-9���u�̯H��]ݾ�_M>�ʾ>�jC��i���������i��X{=�w:?w�?%9��nڰ���u��O���?R>�5\>A=uu�=�EM>��c��ƽ�	H�u�.=}�=W�^>-X?c�+>듎=��>�f���,P��d�>�EB>�d+>��??��$?b��"U�����;�-��Fw>fw�>��>�D>`|J����=�W�>��a>Tq�AÃ�֔�&�?��YW>�9~��q_���t�my=U��B��=���=a ���<��Z%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾQh�>nx��Z�������u�b�#=K��>�8H?�V����O�N>��v
?�?�^�ߩ����ȿ5|v����>Y�?���?e�m��A���@����>9��?�gY?qoi>�g۾K`Z����>һ@?�R?�>�9�|�'���?�޶?կ�?aI>���?�s?�k�>�0x��Z/��6������ p=�[;�d�>�W>f���xgF��ד��h��u�j������a>��$=,�>QE�[4���9�=��I���f�<��>�,q>"�I>W�>v� ?�a�>}��>�x=�n��Jှ������K?ٳ�?��Kn�m|�<�=�=�]�N8?�=4?�_���Ͼd �>y�\?L��?�Z?��>i�iA���ڿ��ʹ�tT�<QiL>��>���>�/����J>�nվ��C��j�>�b�>~����tھ�=��7T��~K�>�k!?��>��=8  ?WU!?e5>i��>	C�zh��R�E�d��>�<�>Q�%?o��?*%?�w��V-�X���|j����L���d>ųp?YX?;�>����͎��)�<!7j�U�˽&��?��e?E�����?Q��?�M?4�J?\�Z>ϹZ�l]��D舽_<�>�!?��z�A��b&�zu��?;�?jH�>E����Խ<Iܼ �r����?k]\?0o&?�\���`�H�¾Ӂ�<�3+��uZ��<HC�0>��>���=٨>悯=Nm�ǳ5�K�r<�`�=Y^�>:��=��7�9P���;,?[cH��׃�?�=��r��pD��>u0L>9 ��?�^?r�=�B�{�`��y��~�T�~��?���?�h�?3����h�0=?��?�?�>�F��np޾��Mw��x�	s���>���>:�m��"�v���+���1@��ƽ����>��>M�?$��>�O>Ё�>ڛ��,��N������]�Y��p�:���+�6��p���}�"��þ`{����>�9���}�>^?f�j>m�r>{��>�A�o-�>m�S>���>��>�5;>��*>�W>�3�<C+ֽ��Q?`���Y2(����1��L^A?,�d?>�>��h��u����p�?���?�W�?'u>�h���+�l�?��>�:��c�	?��<=��/����<�)������ ��W���R�>-����9��M���e�3g
?��?焼�<Ͼ���W�����n=N�?�(?�)���Q���o��W��S���7h�j��$�$��p��쏿�^���$����(�go*=�*?@�?Ì�̖"���&k��?�Bdf>�>�$�>�߾>tI>��	���1�C^��L'������R�>L[{?`z�>ŋI?�<?�rP?�nL?'��>zg�>x.���o�>�l�;H�>7�>��9?�-?�00?�l?�d+?<c>9p�������ؾ?c�?/M?�?�?�ۅ�ewý�"����g�ιy� Y����=J��<��׽�Du�`U=�8T>�X?�[�g�8������k>ds7?�c�>��>���e.�����<$�>��
?�V�>� �}�r��n��[�>��?;y�р=��)>��=�܄��_ɺb��=93¼�=����<�|� <݅�=�=wSe����f{�:�;U��<�&�>�?6v>z��>������j�����<z�>�n�V>�X�=�0پ~Y|�G���Q
k��Nf>?�r�?0��<� �=�ef>�ݾ	�����ɾH<�� ?�??�?�}�?�/E?�y2?@�>[�;�����bv�a�U���?t!,?��>�����ʾ��؉3�۝?h[?�<a����;)�א¾��Խޱ>�[/�d/~����AD�R����i��5��?쿝?OA�P�6��x�ܿ���[��t�C?"�>Y�>��>U�)�z�g�q%��1;>��>cR?�#�>��O?�<{?Φ[?�gT>r�8�|1���ә��E3���!>=@?��?�?xy?�t�>��>�)��ྒT�����@�<ႾOW=%	Z>e��>�(�>G�>��=�Ƚ�Z����>��`�=�b>L��>���>��>1�w>�L�<&�G?��>���e/��襾�|��'��hv?�̐?К,?1l�<�x��EF������>g��?cS�?0�)?��P���=�n���;��2l���>3u�>���>T$�=	�.={	>�G�>�Z�>����C��7��R��@?sC?���=��ɿ�s�����b���=��n��b�\���a�_L	=�S��K��������>�ў����+ڴ��J�����̶?�>�D)>RS�=�3=������;��<�Um<�=5Z�����<I<���*�<O��h�ʼ�ӻ��l=��ͼ��ξ�`y?ŘJ?ސ?u�Z?�.5>�>fֆ�r�>Dm��R?��>Q��=H_P�<�)���޾��ݾt�	�����I4��&_ľ1�L>��<��>!�>�.M>�9����=䀝=�� =���q>�=��=J�2=�`x=?�=��P>�C�>��o??j_�l*���e��9[�n�?*�0>���=.c��A�	?J�,>��������=7���~?g��?D��?`f?�.*�DE�>��0�Q�P����0=~V��P>"�T=���>��>�G�(������#�?�� @Ӵ/?q������M&>�7>�>��R��T1��\�.vb��Z�&{!?�n;��v̾�>fG�=�E߾b�ƾ�3/=��6>3xd=t�A\��\�={{���;=��k=���>��C>��=B��/�=Z�I=$��=��O>$!��%8�B�.�h�2=t��=z�b>��%>Ւ�>1�?�_0?>Yd?�,�>5n�DϾsB���9�>��=]<�>Qʅ=�`B>(�>��7?�D?�K?���>1��=`�>��>�,� �m��h�qЧ�լ<o��?�̆?	ϸ>�XR<��A�[���d>�q>Ž�t?AQ1?�j?�>h���T�\���N0�[:�<���=��=����ب^=�g2<@+�/Dd�4�>��>+��>❚>�d>�>��o>/�>�>>�=��=Hu�;��<�r�9T�=��#��w=�C��̒:��չ9�J�Xa=�^�;DzU<����S���=#��>{2>���>T�=Mﳾ�/>Ɩ�U�L�f'�=�f��)B��1d��O~���.��6��C>.IX>t����/����?7�Y>�r?>�v�?@3u?��>�N�j�վ�K��$8e�L!S��=?u>�v=��x;��B`���M�T|Ҿ{��>�ߎ>%�>C�l>q,�2#?�7�w=��Hb5���>�{��6��'�99q�@������i�-)Һ_�D?�F����='"~?��I?>�?č�> ��ɆؾW;0>�I����=3�j*q�_h���?)'?%��>�쾽�D��;��=r^��N�>�"1�ݛi��;b��ON�(�$� 禾Ӄ�>�ƾY�ž�-���������a-�a��#�>�:(?�K�?����
��q�>�,�����>�XU?�M`>N�?%��>�J.����FQ���d�=��?���?�"�?m>���=���;�>�+	?O��?���?��s?|?��y�>�K�;�� >����LK�=F�>���=6(�=-s?ב
?��
?�k���	�����m^�F��<�ϡ=2��>�l�>�r>���=�g=y�=�.\>�؞>�>@�d>��>�P�>�о���96?�X*>Ԍ�>y�??v3{>�����E��+���b�����нo�ü7��6良E��
)�<�|���?#�ȿZ�?u0>�K%��R?� �[���X`>�W>�?�d��>#��=�?#>��>���>�>�ї>+>�FӾ0>����d!��,C�A�R���ѾJ}z>�����	&���Yw��"BI�_n��yg��j�L.��V<=�iʽ<3H�?����k��)�����U�?�[�>�6?tڌ�w���>���>�Ǎ>�J��g���Tȍ��gᾤ�?<��?F�>S�7>M?ք?���Y<伮T��Bp���?�0;���N��P��%ց���8�=?���g?3�?[�_?Ӻü|�>�&�?�S�B5ﾹL�>uC�k
��49>%�>Rf��eVڽU�������ܽ��>��{?~qr?��?��
�j���L>/�<?�1?tq~?�f+?��A?+R�M%?��>�?��?�9?�,?�e ?ƺ�=�qH={6K����=TTý�9���>Ƚ�ˣ�!O���=P�=W3f���<5�=��<g�s���R�Iu�:�J꼷��<�Z=�e�=�B	>���>f�U?}��>R��>�t1?����7�S]����?��l<T/��掾昧�$"����>ڂi?�ӫ?�>X?�Z>��K��B�o�>��>�@>Y�R>�]�>�9 �C7@��v=B�>�}>��=��~��%��3H
�ŝ��{=q>)w?�;>����]>y������#�=������B�����T��*A��užl��>C�^?��1?d7t>�ҿ�� ���Y� ��>5�7?��f?��Q?2S�>Ԯ�Af������������>!u�>��Ѿ����)>��R<�(��=��}>qן��ᠾ9Sb>H���q޾��n��
J���(/M=G��/V=	�� ־e6���=}!
>|���	� �����ժ��0J?�j=�r���ZU��n�� �>�>�߮>t�:��v�χ@�5����*�=��>1�:>fq������~G��8���>|VE?�_?S�?kz���Ns��fA�	j���Ρ����?=+�>�*?�A>���=�F��8�)�d���F�b"�>O&�>C����G�,��?,��Ħ%�'P�>�,?�">2?�R?��	?��_?v�)?�%?�~�>���4���?&?B��?���=��Խ4�T���8��F�#��>��)?ܶB����>Ԋ?I�?}�&?�Q?��?`�> � ��B@�ǒ�>�R�>D�W��a��|�_>-�J?���>�:Y?փ?a>>Ã5��ꢾ�ѩ��f�=�>V�2?�4#?�?���>�b�>�J�~=Y3�>��f?���?��r?SG�=�?��x>H6?	�
>��>wY?i?J�J?�i?Ă9?��?���<�7���۸�2v|�[l�ݚ����<��=�W��Y�u�5I�$4�<�q��RƼ�NQ<os��p�����/¼�X�>��s>]����0>�ľU\��YA>�����J����:�x��=�>�?.��>Fl#����=���>$C�>���?/(?*�?L?��$;-�b��۾Y�K���>}B?|��=�l�}�����u�Bh=7�m?��^?��W��&����b?U�m?��+��4?�ν��-x�d4���z?u_�>ܜľp�>r k?k?��><����7��_���|Z����M�<��>o�����]���>�@)?�]	?�>f�@>�	�Jz���W�?b*�?���?�ϊ?mH=�-��'꿃���Z��[~\?:��>ddo��7/?��R�|��1����Ǿ�L4���ھ(���е�4n̾2�P��V��eq(��v=7|*?��y?h��?�y^?����,���0�CtW���L�5����x7�CG��V��\[�!��H��/9���2z�jgź=�����=�.e�?��8?@��yl?�+��Gd��t���L@>�霾k**�tS�=LD�Z.ռG|�;<�w��i=��ž���5?�Y�>7"�>�02?tނ�T����C�8�4��=׾9to>�m�>V�>5��>Cf$<0���߽絰���
�b��18v>n�c?��K?5�n?9:�G,1�u����!�y�/�q��_�B>lm>Xԉ>�lW��Z�<&�T_>���r�G������	�'+=�2?M�>��>M�?W�?�b	�u��{x�i~1����<�%�>��h?)�>	�>oϽʹ ����>!�l?�[�>���>Q���	^!���{���ɽ��>_��>���>~�o>�|,��\��d������>'9��m�=c�h?����q�`�jυ>��Q?�_�:��I<j��>�u���!�/���'�6>:�?�=�!<>�zž$I�,�{�&>��F�'?X?쐾�_*���>��#?��>v��>�)�?�ݟ>� ���<�2?�#`?�I?	�??���>�=�Ӛ�w�ýl�%�
�)=�L�>	�X>@u=��=0�e�b�qX��5O= �=q!Ҽ����$<�ɗ�O�q<&y�<A�4>�lۿ�GK��پ����9
�,������Qf��{���w�����Rx������&�XV�z-c�����	�l�ׂ�?�<�?�b�����O���l���C���۳�>��q�^/��#���:��4��|��dʬ��f!�:�O�:+i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@}A?�(�����V=>��>'�	?�?>�S1��I������T�>s<�?��?v|M=��W�w�	�*�e?�~<��F��ݻ�=y;�=�E=���͔J>|U�>����SA�N?ܽR�4>Hڅ>�~"�a���^�O��<��]>J�ս,;����?�{Z���e�0�/�(J����
>�U?�K�>��=�t,?5AH���Ͽ)�]���^?	�?��?\�)?���O=�>�ܾ��L?��6?+��>��%���q�e=�=�������Q�⾋V���=?;�>@>��%��!�h>N�8����=%���V�ȿ����d�X�=e�p;��(��5���xy���-���KhP��@��H��<i�>#U>P�>7O>,��>��M?Dt?�k�>H�Q>֑(��;"��s;�dԼ�@¾,���П����;�Ҥ����4������H��+���ھ!=��=7R�k���@� �h�b�[�F���.?�v$>o�ʾ��M���-<�pʾf���\܄�=᥽�-̾�1�"n�i͟?��A?������V�L���W�@���Y�W?,P�߻��ꬾ��=��l�=%�>���=���� 3��~S��~0?�V?����~\��f�)>�w�$�=v�+?%^?Y[<�֪>��$?U�+�o�佒�[>�k4>��>���>c�	>
��K�ڽ֍?U�T?���z���?��>ߔ��H�z��`=��>^�4�4�弜V[>V�<�!����S�j����<��\?��>�I��,������|��~'�?��>>т>7�k?D0/?�0b=-vپ�O�B^+�괓�I?'t?���=%�=0tѾ �߾�G:?�{T?��c>L٫��rѾ�X��ؾc�(?L��?�&?�>W\}��ݫ�OF�>�1?Ez?��B����N���]��T�1>ܶ>�,�>NE��|�>�:?�k��>�����¿[ T���?�I@�g�?����λ��>���>=��>�������C�=�R�Z�4��>�V��9x�~�#�͏���.X?WI�?��>�❾�m�����=�ٕ��Z�?��?����"Gg<Z���l��n����<lΫ=��F"������7���ƾ��
�����ῼॆ>BZ@�U�p*�>0D8�\6�TϿ'���[оbSq���?N��>��Ƚ����D�j��Pu�T�G��H�ƥ��ȣ>�>������
|�&t;�1�����>�Y��~�>�R��붾����<�Q�>�>���>����1A�����?	���Cο㷞���x�W?&e�?��?��?Q�+<l�v�&}��@-�;�F?�s?�[Z?a%���]�1/�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?���>@.�?=T�=K��>W�=����=����_>���=����>gM?Ho�> �>�ϒ��E*�y�N�\K^���'�IP8��*U>ڨs?�9W?6r>C�������4����R�h��Z=�_Q�A ���R���/�=d.3>�;>b�޽-����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��f?ei���=e�lYT���*� A+�a�?��??8=���>�>�>��e����ݫ�Tɏ����>\1�?��?p!�>]
c??NC�=�g��$��>��?�\?|W>��#���)>��?c�;����2���FW?X�
@�_@��X?���ҿ��VP��N�|̜=h`>@�0>�Q=�U�;>�}>�=��b=��&>���>/�>�H>}w>�->>4	>���*�.����l���6��$�&��3W���6P������-����ξZ�����a?�.̽���M@Ľ/�>bXg?��J?�op?A�>��m��;b>�#��i�;w;����=��>3y0?��8?�#?��ʽK�羃^k�r�q�O[��)������>�*>��?u?�N�>ϭ����>���=�*>*?=��=�R�;$h����=��>�
?�?�D<>��>lϴ��1���h�Nw�?̽X�?����ļJ��1���8��ȥ��k�=�b.?�y>��?п����	2H?m���z(�ݸ+��>��0?xcW?*�>����T�w8>���v�j�!a>v* ��{l�ҍ)�j"Q>�j?`yh>u{>]�3��8��2P�ޝ��z�{>>�6?�@���h>�`�t�ԭF�dT۾W�O>���>Yi�7K��D��g���j�`Hy=/a<?��?�ղ���P�w�kx���S>�`>�"=vV�=�K>��b��̽y8D��==)��=��\>�o?�!,>�͍=���>Q���@�P��ϩ>Q�B>�I+>b�??z�$?�z��������j^-�F2x>���>Lb�>��>+gJ�^�=b�>��b>���=$�����,j@���V>��}�s�_���s��{=M����=��=�< ��<���#=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿhh�>x��Z�������u�}�#=��>�8H?�V����O�>��v
?�?�^�ة����ȿ<|v����>W�?���?H�m��A���@����>1��?�gY?�oi>�g۾�`Z����>ۻ@?�R?�>�9���'�I�?�޶?ʯ�?�I>)��?%�s?yj�>�x��[/��4�������s=�Y;g�>�^>����eF�֓� h���j�����a>��$=��>�G佟4���:�=.苽�N����f�f��>d9q>�I>�V�>2� ?W`�>v��>e�=�d��>܀�����9�F?~Y�?�/���i�Պ��'�/�����)?�	?�\N���Ѿ��>qQ?2�v?��o?��#>P�0�T:��]�̿���w�=J��>S?�x�>��g��
>%�����p|�> �>��{=(پˢ;��S𼮨�>�*?�2�>��ѽ��&?ު&?���=8�>��G�e��Z.R����>�X�>e3?��v?X�?�y���,�|�������hI���^>��s?��?,�>-���q?��!�=�ꀽ���a&�?�|^?��B��?��?2W?0nN?��r>�����A����8�>c�!?���A�rS&�����{?+O?���>n���ܳս�Tռ#���d���?\?:/&?����#a���¾��<$�>R��@�;CQD�B>�>�=��	��=|�>�T�=�4m��#6�	6l<�Q�=�}�>���=�s7�����A?7��=Gr��n��==x��NL���>BV�>����M}C?���(���쯿D������
�?�Լ?]��?9�h=t M��)?��w?7�A?8��><���E澑���c���~��W	���9>� �>��ѽ�X��m����w��Z��AU� ������><?�?��?��y>�#�>*j���U!�4d��.��9d��*��C���)��������:�m�鏓�/ْ������>�~�<;ա>S
?�>w3�>�}�>��>	E�>�r�>N��>M��>��P>֣>���=H��<`��PKR?�����'�P��7����1B?rrd?�3�>i�����x��N�?D��?�r�?�@v>h��-+�al?�;�>����p
?\:=�K�u=�<�X��$��}<����몎>B׽�:��M��mf�Nj
?�/?4���Ӌ̾�H׽���>�S=���?�*?-2)��wM��<p��X��'R�13+��Xw�W��|2$�Op�?%��.߃�������'��%=(�+?s�?��������ﲾ��i�B=���b>>!�>��>�o�>)+I>;���2��^���%�����C�>xy?�J�>��I?%�;?�DP?�fL?%2�>9k�>����?�>�/�;d
�>��>�~9?��-?�0?��?��*?��a>4������B�ؾ�?;$?� ?pc?�?są�����%��g�n�Hy�-����H�=*��<ma׽�qs�DX=�T>�<?6����8�����NNk>`}7?���>���>R���(�����<b#�>��
?J��>E����fr��a���>���?�����=�)>���=�ㄼ���V�=�qǼ��=����U=��� <���=��=�nw�2ȿ�jF�:�Qh;aŲ<P�?�Z?��r=M2�>̾0���
�FQ�=�I�2Yl>&�=�*�z뇿/���	)^�y�\>s�?�y�?�ۼ���=�R>��ﾠj���ӾGt��yqB��d ?�<.?CH?�Ƒ?VNH?�sI?���>_!&�Y"��刀�B|���o?��+?��>w��oʾN���w4�r�?k/?/�`�J��(�m�����Ͻ/�>h�,�!v}������@E��'��������"�?Y�?|(@��n7�S#�u��x:����C?��>M��>���>)�%�g�`��n*>>(��>�;Q?��>��O?�9{?��[?�zT>2�8��-��Й�4�2�G�!>q@?���?��?Ry?�v�>��>;�)���ES��d���5����w�V=q Z>O��>
�>��>�"�=ܧǽ_S����>�([�=ؑb>���>��>#�>��w>�f�<vqH?P��>E��? ��Ϩ�-y��ˇ,�2Rt?��?��*?���<���PhG�%P��/��>���?�#�?��+?��Q�{R�=������7�h�i�>���>/�>C��=�� =��>�w�>�f�>k��tS���7�>Ek��y?�D?��=A/ƿ~Er�o�m�Q{��k��<슑�.�c��M��p[����=����3��b��g�`��V��?-��}ȴ����B|�Ī�>;��=��=̗�=�r�<�Ǽ�r�<��U=���<�	={a�!�<�<���ɻ������.��D<�D=�/���!p?�l@?E?��G?^�=e�G>H���N�>��H��?

�>Õ=�JK���4��l�ľƱ�'Oо�Ǿ�~[��A���E�=l	�Q��=�j>��#��u�O��>�xh>[��=L��<�TѼZ�=Cؒ=��=U�>*/k>s��=�\~?�JV��4���Y�h�{����>��>�1X>&���L�4?�n+>����5Ŀ�I$�MBG?�r�?x�?�X*?�c�����>�qU�5���uj=^	κ)��=Uj�>�N�ܤ�>z��=jL"�1;��)�����?��@ .?t���th����>A�7>�/>��R�؇1�ԋ\�L�b��RZ�_�!?�?;��F̾�6�>T��=o,߾)�ƾz�.=��6>�Nb=AY�K\��י=�{�G�;=��k=}Ӊ>��C>�d�=��G�=v�I=F��=��O>4ה�cI7�R�+�׵3=���=��b>�
&>~��>	�?6a0?Vd?9�>�n��Ͼ�=���J�>��=jH�>S�=<qB>ώ�>��7?�D?|�K?���>���=9�>�
�>s�,���m�}l循ç��X�<��?dφ?#ٸ>Y�Q<n�A�o��Ed>�42ŽZv?jR1?l?n�>G���d�5�!��AD������]7��4Ѽ�?���D���g[<瀬��'�=���=�Q>4+�>��>�>Q�F>�`>�<�>PǶ=����H6>�fj=a�?<����㨼���"ͽ�?	�e=�ԁ�<�08����4��<��U�+�<�M�=g$�=��>�+>տ�>��=�	���Y/>)�����L�R��=�Z���4B��8d�&O~��.��6���B>skX>�m��0����?ݷY>R�?>�{�?�<u?ɭ> @�7�վ�J���,e��S�x�=W�>�1=��;�|J`���M�ӈҾ_��>^ߎ>�>z�l>�,�Q#?��w=��Yb5�[�>�|��}��)��9q�@�� ���si�diҺ�D?�F��Z��=g"~?��I?^�?ύ�>n����ؾ;;0>�H��?�=_��*q��h����? '?���>�쾧�D�ru��>6��?
��<�`x�ۑd�q�T��-�5C�����>n�Ѿ���o2��]�����h2���E��$�>g}.?�X�?+Oݽ�^x�oL���,����\�>rW?��5>=�?h�?�4�ʩ,�z#Ⱦ7��^�?��?�,�?���<K�=�紽�*�>�?���?���?�Ys?mq?�T��>jy�;�">�����=>ZU�="��=��??�	?	�
?������	��o�B���]�Y��<�~�=i�>a�>-Hs>h��=�Ch=5�=�x[>p�>� �>��d>{��>n�>ԉþ���:?}4w>�e�>3;?zGx>TR�\A��eD�<�wW�\~U�˝!���v��o
������"�.���a�RZ?�z���H�?�pL>�5,���&?�
��h��D\>���>@��^�>��>4��>�7Q>���>;�>쒤>\�(>RGӾ�o>���[!�j)C��vR���Ѿ|kz>U���&���V���9;I��g��Xj�^
j�-���:=�3m�<jJ�?.���v�k� �)��Z����?�G�>T6?kԌ�KÞ>���>�>sL������$ƍ�:cᾂ�?���?yh>��>��W?�?��>�Ѱ1���[��u�^�@��Pa��^�Lp������S���㽴�_?��y?�D?e��;��|>�k�?�u(��J���+�>��1�Ō8�ӌr=���>�����uU���پ��Ⱦ���F>܁q?(�?E�?I�W��U.��(<qa	?�9I>��|?"J?��5??I�T{?
�>��?~�:?��U?2kk?+l?
j�=�a_��@a�)��>�~����p�0r$��Dt��J�<��=��=�M%�8I�=|F�=z@�<"�=H�����=�w=��=
�=�=���=T��>/K]?�U�>TJ�>i5?#��؊6�U��L�+?K9=��rv��vq��������>Zk?r�?��Z?i�c>7HC�A�׉>E��>��$>��]>Q�>�\���J��=k>�>Q�=��]�޹��Y���?����<��>���>��>�X���7>s<�������q>��D��Vž#�M��J��S7��͆�O��>3J?F8"?-b�=Z�׾�σ���c���&?�Y7?>yR?�x?���=�?�5;�8=N��]!�eϜ>��=�s�����}��n�?��V<�v>�
���ޠ�UWb>5��}t޾u�n��J����iGM=��u\V=����վ56���=�$
>������ ����֪�{1J?��j=Jx��QbU�Qp��^�>|��>�߮><�:��v�d�@������6�=D��>��:>�b�����G�(8�w>�>OQE?0W_?"k�?"��Rs�8�B������c��{ȼ:�?Fx�>h?.B>��=,�������d��G���>���>d��-�G��;���0��2�$�L��>T9?��>��?Y�R?r�
?Y�`?�*?0E?7'�>�������A&?B��?E��=� Խ#�T���8�zF����>�q)?��B����>{?Ѩ?f�&?,�Q?;�?R>+� �KC@�u��>DY�>�W�~\��8�_>�J?���>{SY?\̓?��=>pk5��Ӣ�/���[�='�>��2?�8#?��?(ø>���>�����="��>�c?/0�?��o?G}�=��?�;2>���>c�=���>��>r?�VO?��s?��J?���>7��<T@��b4���7s��O�((�;޿H<��y=^��p4t�m=�F��<�R�;�[��I��i��µD�吼�2�;�^�>�1t>���s�0>��ľ�K���!A>����]��튾y:��&�=2��>L�?Z��>I�#���=��>L�>
��W:(?��??[�!;3�b���ھ��K��M�>��A?',�=��l�y���u�@Hh=��m?��^?lX�MW���!Z?2c?̟�0%;�?�Ok�����c?Q��>f���?�>~�}?]Iu?�Y�>y,v�8hr�*��2�7�6�>�=�(�>� �bO��ӎ>N�6?���>��>deX>�>�x��d/��� ?u8�?u��?���?�L)>����f�ڿ#� �#���3}?O
?�	¾M?�A��f�������&�v��,��̘�F������BBB��g�g:��o�;o>?��V?��Y?��H?��A��C<��-e���~�H>P�w����3�utQ��'Z���I��T���g���6ҽ�����䄾5�C�x}�? j*?c�2�P��>�L��a���˾��I>�&�����g|�=���	=Ux<=ӽg�"�,�i����%?�Z�>���>��:?h�a�Ԡ7�n�3��6�¶����A>A��>�e�>��>CJ׻K{'�:�������7ku��ܽnLu>��c?�iK?��n?>k ��k1��=���X!��O-������PD>D)>�܉>!X�Cv��]&�{|>���r��J�S���&
�R�=��2?4o�>��>�Q�?F�?K0	�p6���@w�p}1���<���>�uh?7s�>���>�ͽ� ����>�l?gx�>F�>�M���a!�s{���Ľϳ�>+��>�7�>lNq>4�*��[�^��y�����9�ۓ�=��h?w��� �^�3�> �Q?�k�:�dU<�r�>��v�]!��o����)��N>��?�\�=�P=>�ž`����{�#��'�)?b�?~l���[+�\�}>GG ?(4�>���>,s�?���>�ǾH#��}$?`�_?P2K?	(B?N �>��=غ����Ƚ1q#��h8=�׈>�PZ>�Ts=,b�=��uc���z�H=�ƻ=�Ļ�K�����<�5ż��S<)]�<^E4>@mۿ�BK�s�پ�R�v?
��爾g����c��ݲ��a��6��YXx� ��R'�lV�l7c������l�Ї�?�=�?!���p0�� ���=����������>~�q��������j)����n���ed!���O��&i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�|A?X�(�,��jV=���>��	?��?>Q1��I�?����T�>@<�?���??~M=�W���	�ie?^�<��F�	�ݻ�=�;�=>C=E���J>V�>���4RA�,@ܽ��4>�م>�}"�O��m�^�ǅ�<ч]>��ս�<����?D@U���f�w�3�X�|����=.:?���>>}�=QW!?��M��gο�a��%g?�i�?���?!p&?�^ʾ�9�>��Ѿ�[K?;Q'?�B�>g~��s�?��=�JƼ��	��+�Q�L >��>�y8>�K�/M	�'�T�� ��	>(A�A-ǿ]�$��  ���=F@ͺl�U�+�� 7���$Y������k�7ཤ�m=%�=K�P>�b�>4�W>�LZ>�$W?Sk?�Ͼ>{>������5G̾:��&��p���܊����l��_^�a߾�i	�\������`ʾh =���= 7R�a���r� �5�b�|�F���.?w$>��ʾ��M�Ay-<Hqʾ@����Ǆ��ۥ�9-̾�1��!n�7͟?��A?�����V�����`�(���M�W?�O�����ꬾ2��=ͦ��:�=P%�>���=���� 3��}S�!x0?\?盿��s��/&*>o�R=��+?�{?^�V</�>�D%?��*�ϸ��}[>P�3>���>g��>D}	>��"�ڽc�?i�T?Q���朾u�>hv����z���`=>�95�v[�X�[>��<U쌾�U�ݜ���r�<IS?��>��:�uR)���z�8��V�<sɉ?C�o>�,?=�~?\D?j�>����c�4(�æ^�@��?MiS?p��=���=�[���5��d�(?F;F?^ڌ>�!'�x龾��b��9��B0?<3�?+l3?�Z8=bJ~�e���5���?��v?
s^�js�������V��=�>�[�>���>��9��k�>��>?�#��G�� ���yY4�$Þ?��@���?�;<����=�;?T\�>�O��>ƾ�z�������q=�"�>����ev�����Q,�k�8?䠃?���>���������=�ٕ��Z�?��?����Dg<R���l��n��~�<�Ϋ=���E"������7���ƾ��
����ῼΥ�>EZ@�U�u*�>�C8�]6�TϿ)���[оSq���?K��>Z�Ƚ����@�j��Pu�a�G�3�H�ť��[�>|W>�ߓ�%Ƒ�d�{�n4;�������>Q��8�>�T��X��Iɟ���1<��>���>���>B���a���Ù?o���?ο]���ޛ�b�X?�P�?�d�?ec?��8<_w�||����w(G?Z�s?�,Z?��$��/]�NB7���j?�[���U`�ގ4�>GE��U>�"3?�F�>1�-� �|=� >#��>l>�"/�ǍĿoٶ�p������?<��?�o�1��>���?�r+?�h��6��nV���*�ڢ'�u9A?�2>#���Ʒ!�.=�:Β��
?�|0?;���.���i?X@��<u�<�F��V[����=�ʷٽɧ�;c�T��|��m�����~/�?c��?뢸?]A�z�,��'?O��>2%��48��,�����?a��=/�j�/
v���/=�\!��I�y�>�j�?6�?6��>J�h��茿�¼�1�?�>]6�?I{�<o�/>e�>uUھq>��>��=��a�Ek�>�+L?l3?�U����E��/���Z��M�5�J��8��g>�
m?��C?�Ax>v|I�޷�%/�%>�}�M1{=�W��/��RN��߅=]:	>o�?>9���8���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��S?�
�\�v���j�����L��Ӏ�=�$?E��3�>� �>ta�=x�r��媿�s����>{0�?\�?���>v?��b��I��=��k>#c?L4?�4$�t��P>��>�&�������7,c?D�@j@�a?{ٞ��\Կᮜ��H��O��9�=���=��?>�� �x+�=v�Xfo={=��@>l��>��W>t\>��<>3S>]rG>f����(���������D��$�	!��>����'������\渾���2������z��O&6����8��a�=XW?��O?g'n?�� ?�`���%>�����?=-�0���=��>��0?�yE?�#?s�G=F֥��e�՝��� �����f��>��[>��>���>%��>$?�;%nJ>��8>�,�>,��=�pa=�:�V�<�g=>nͫ>ݓ�>L0�>\D<>��>Eϴ��1��@�h��w�d̽�?a���e�J��1���9��2����k�=~b.?V}>���?п����2H?����n)���+�g�>G�0?pcW?��>���R�T�K9>L���j�W`>�+ ��l���)��$Q>�l?�h>��t>�4���8�EP�N���w>S�5? ۶��z;��Uv�(�H���ݾ'�P>�+�>�c� ������e}�7Xi��h�=�j:?֬?^��6!����t��]��d&N>O�\>�v=�d�=@�M>�b���ƽ�H�2C/=Ig�=��^>X?�+>#��="ۣ>.d���DP�,��>�B>�,>j@?e)%?����ӗ�v�����-�Yw>�N�>��>i[>q\J����=�m�>��a>�F�f�������?��}W>~�܆_��uu��x=�3�����=
)�=� �=�m�%=(�~?`��9䈿i�Vd��+lD?]*?� �=h�F<ʃ"�j ���H����?g�@'m�?с	�r�V�z�?A�?������=d}�>�׫>�ξ��L�۱?.ƽSȢ�V�	�C(#�.S�?��?�/�'ʋ�l��6>�^%?��ӾPh�>xx��Z�������u�p�#=R��>�8H?�V����O�b>��v
?�?�^�੤���ȿ6|v����>X�?���?g�m��A���@����>;��?�gY?roi>�g۾B`Z����>һ@?�R?�>�9�~�'���?�޶?֯�?I>���?�s?�k�>N/x��Z/��6�������q=�[;�d�>X><���zgF��ד��h��o�j�����a>��$=��>�E�N4���9�=]�I���f���>�,q>��I>"W�>�� ?b�>y��>x=�n��Oှ����8�K?귏?A��|:n����<�G�=t(^�%7?144?�l_��Ͼ��>��\?߯�?%�Z?*�>����3���俿<���Ա�<�7L>��>?9�>����%�J>�վ�XC�[d�>���>��:Uھ�U��)����K�>	e!?#�>�h�=�� ?՜#?R�j>�%�>M`E��9��l�E���>���>CI?r�~?K�?�ѹ�6Z3�����桿,�[��DN>C�x?�T?�˕>s���(����RE�/;I��꒽͛�?�sg?�h�^? 2�?R�??��A?�,f>u���ؾҰ��#�>��&?��qI�}b-���0��>�B�>$�>����kE���ܽ�g��y���?1{d?|v/?�1���Lf�aI��{�<>�<�(�<N^=���K# >��>
��6�<p�>���=�R�c]���z<���=Ii�>:��=�8�p�?�j=,?��G�Xރ�K�=��r��wD�~�>�QL>�����^?Vb=���{�����x��@U����??��? l�?�����h��#=?F�?�?"�>$J���~޾���Qw�tx�5u���>��>9�l������o����D��Oƽ�I�z�>���>�?�� ?qcO>wd�>�)��M'��񾗚�?�^�0U�<m8���.�ޫ��䠾I7#��m��A¾�|�>N�>x;���>ӳ
?(Jh>*�{>��>^˻ D�>��Q>ݱ>Ul�>��W>��4>��>c�<��Ͻ��Q?@���(�p�V����@?
�d?���>����y������?�|�?%��?4jr>�h�^-��?K6�>$܀���
?j�I=ǥ� ��<�/��iC���ټn��>]��,�9�O[K�@�c���
?��?�}��|Ѿ�c�9�����n=N�?��(?�)�}�Q���o�θW�S�^��~6h�Hj��H�$���p��쏿�^��%����(��r*=*?c�?��� ���!���&k��?��df>Q�>t$�>%�> uI>��	�m�1�^^�M'�@���dR�>t[{?���>k�I?T<?QxP?�jL?���>�e�>�1���k�>���;b�>��>^�9?��-?m40?qv?7q+?!)c>/������ɇؾ�
?^�?�J?E?�?�؅�Bgý�o��,�f��y�Lo����=B��<&�׽� u�&�T='T>�V?��$�8�o���#�j>_�6?Ӵ�>O3�>Y ��D�����<���>��
?�D�>K���k�r�X&��i�>*��?
��D�
=��*>D=�=���/[7a*�=
ZǼ2�=����1G�x<4��=���=)������:��:z��9Pa�<�,?�?���=m�q>z �������E��ٔj>��<LP�>H�>�2Ӿl���ș�Sa�{jL>aל?���?�1>v;�=!H�=�0���9���������0� J�>�!�>"�p?��?��R?�P?�R=��D�O����)�����8�>�#,??��>+��C�ʾp���3��?nW?�:a�����C)���¾�ս?�>�M/�u ~�����D���~�.���`��Ś�?k��?�0A�s�6��j�t���=m��Y�C?|&�>ET�>�>��)���g�U%��1;>���>R?�'�>)�O?3{?�[?$RT>�8��-���ә�'F5�d�!>�@?���?��?�y?���>m�>Ó)�@ �r^�� ����₾W�W=��Y>���>�4�>��>���=X!Ƚ�����>�=F�=:[b>�~�>(��>�	�>�w>YS�<��D?���>yྮF��1>������44м��z?>[o?��?^D�=W5��Q�$i���>%8�?�۰?��$?�B�MC>�j��Qþ�
��v�>OL�>���>1S>�[����>� �>ݎ�>21�G�>�k\����?�?�`?zr[>��ȿ �q�Bh	��[�*�v=~mI��>��|���`L�"�=ڐ����7�����l�b��
#������u����x�-�?�2m=�A>ܯ'>d�ɹ"�=!5ܼ��=��<���=���[U=>��
d�;��Q�I�$�/"�;�X�<@	��X��)G?5;H??
?�Y?U��=(�?.�Z<f?��Q�-M?_�>4j8>c��=��q��Bk���v����M�������)E>b����<>x�>� >p[�F�>X��=DUI��������=�h&=x� >��=�P4>�O�>6�r?4x�����u�Ծ|P?�_�=�����c����O?e����_���I���z���n?�8�?ޮ�?R��>������>[|��2���z�5��==K�_ =�ŧ=�Q�>�q=�P���>��7D3�Vf�?�@�g8?;���l˿0}S>�7>-&>��R���1���\�9�b�9�Z�ś!?sG;��Q̾:'�>��=�/߾l�ƾ5�.=��6>)ib=�x��L\�ޙ=۵z�u�;=�l=�ى>��C>�r�=�D��f��=B�I=��=t�O>�2����7�7,��3=��=��b>E&>�u�>?�?��y?��>�xv�S.ž*���?M>#"=�l�>��a<jO�=S��>$%A?@??V?�O�>ݏ��D��>�f�>g�1�]`��hҾ����+o�=<o�?�Yz?b�>��=]K�\���rZ���;�d��>8�4?�?�@�>�t��X�0#�d>�7�J�+�{;��=�=���~����
����ػ�bk>*ڷ>��>�ߑ>Dx>��Q>	�R>Z$�>8X�=�߁<���=�w��(Xb=�-�=ё�=�9E=�0�<��/<HV=s��:.����ټ�x`�>w���ļ�<�
��=!��>j<>լ�>K��=���D/>Ը���L����=�G��a,B��4d��I~�N/��V6�j�B>;;X>�}��@4����?^�Y>�l?>���?WAu?D�>� ���վ�Q���Ce�.VS�Y˸=E�>�<��z;��Z`�~�M�a|Ҿ��>��>���>N�l>P	,��!?�x=3�ᾢd5�t�>�s��Yt��94q�:>������4i�%4ƺןD?6E��-��=� ~?ЭI?�ߏ?ʐ�>(嘽��ؾ.J0>�Q���v=D��q�R��� ?�'?���>�$��D�C�Ⱦs��?@�> t4���S�AV��at1�����[8���$�>����էо�2�H펏�b ?�5�b�ڂ�>�eI?T�?W�W����jM��Z�]���% ?�y`?X�>ޟ?9/�>SB佅q��'�����=��u?m��?6��?~�>��=Է����>t4?[ۖ?}E�?�s?�@����>��;��!>����,*�=��	>zY�=ab�=�k?+�	?��
?o:��Ne
�8�����:�[��=��=�Α>C1�>�@r>���=�Ae=K0�=k^>��>���>�.e>V�>�x�>�Ծn�WQ=?4<^>b�>*)J?=�l>�p�������-=��ۙ'�����ݽ5�+�h�J�P����'w��?M��'��?B>f>�&�l%+?�s��g���
>ѩ�>^�V��>Z�>d)W>)�>�٨>�D>�k�>x��=�FӾ�>����d!��,C�i�R�`�Ѿz}z>�����	&����	w��BI��n��xg��j�M.��]<=�pƽ<H�?Z�����k���)�]���[�?�[�>�6?lڌ�}��#�>���>�Ǎ>�J��f���Sȍ��gᾡ�?C��?�iu>��Z>�J`?c4 ?JZ��9O׼��Z����&�<���=���l�_����������`��c?Hj?ͨM?c5:���>�_�?��>���kI>�f3�Z�.��t=���>��� ox��'�PO��H�>�u�?��?E?R�  l�?�M�`�(?��>%F�?4?��5?�@W�{*h?H�8>�j?��#?��9?���>���>�~�<QhO<!9��n�C>�[���ܾ	T1��L�g/�Ǘ�=-��=�ݐ��l=�4a=�=w� �<л�=���<Ny�=���=���=�Q�=w��> �]?��>�m�>�7?=^��8�ٸ��2�.?87=���B������V��>Tk?��?�
Z?�e>��A�I�B�N>���>H&>�'\>G��>�ｷ1F��9�=j�>?t>���=&�N�9Ձ�?�	�N���@�<�>�?��>c6��m>�:��Z�������pѾ��BMf���W��x>�+x���)?�s?��7?�i:>b����5=�
O�NI&?֣F?�?�1?EG>"J���"��A������;
? �F<\�߾+��e:���[F����=��>����٠��hb>1���޾��n�F	J���,�M=�{��gV=�5�վf<��~�=L

>v����� �t���ժ��+J?�j=�m�� FU��q����>k��>�ڮ>��:�zw���@�Y����0�=`��>��:>�њ�%�b�G�V8�h>�>JQE?8W_?k�?
"��Os�:�B�|���uc���ȼI�?Yx�>h?�B>?��==�������d��G���>���>Z��>�G��;���0��=�$����>J9?�>v�?>�R?q�
?n�`?�*?IE?*'�>��������C&?��?���=!ս��T��8�CF����>dw)?ФB����>�x?��?j�&?�Q?��?<�>Ĭ ��7@�ᒕ>�e�>s�W��c��2�_>�J?|��>/HY?�ڃ?��=>��5�P���o>��T��=>=�2?w2#?��?���>p��>A�����=�>�c?�0�?!�o?��=>�?�:2>P��>*��=���>W��>�?PXO?=�s?��J?��>6��<�7���8��!Ds��O�ǂ;�uH<��y=٘�3t�K�1��<�;�g��9I������D�6���^��;��>'�X>���{�=>�w���1���!>�fD�5$���߅��$A�q��=���>D>?��>�o�=pӼ>�J�>c��o.&?���> ?E�7�+�\�Kξ}H�Av�>�xF?���=��q���s���q=]q?c�Z?�r���O�b?��]?Bh��=��þ��b����f�O?:�
?A�G���>��~?g�q?U��>�e�-:n�)���Cb���j�Ѷ=Yr�>EX�M�d��?�>r�7?�N�>�b>%�=cu۾�w��q��d?��?�?���?+*>��n�Y4�w~���K���^?G��>Z>��� #?�2 �I�ϾRQ��P)��-⾯������A���w���$��ރ��׽)�=c�?s?�[q?��_?Ƴ �ud��1^�Y
���kV�0'��%�/�E��'E��C�~�n�Da�v.�������G=']���T�ٔ�?`�E?�wV�$0?�ž{����Ԓ->�}���f����j=Gi=���=���=7q�c=���Ռ���K?���>#z7>CL#?��T��V8��aX���W�~�� >8�$>���>o�?��h>M�>r��=x�վe
�/�J=�5v> yc?�K?ܸn?�p�+1����
�!�%�/��a����B>?j>P��>z�W�����9&�Y>���r�	��!w����	���~=��2?�(�>���>QO�?4?�{	�j���jx���1�u��<�0�> i?�@�>��>	н�� �e�>�Lp?��>�HX>fXd��}���m�fxT�t�>7��>��>]>��@���\�挐�먊�V;��-�=m�R?����4Cd���>k�W?����h=餔>�2��)O�͕���@�J��=V%?��=c�>��Ѿ�3��8�����P)?�K?�蒾��*�g4~>�$"?ɀ�>�-�>R1�?�*�>�qþC�E�ұ?)�^?fBJ?}TA?;J�>Y�=P ��=Ƚ��&��,=���>2�Z>9m=1��=����r\�$x�9�D=�s�=��μ~P��R�<�����J<��<��3>�lۿ�BK���پ���i?
��爾«��Jd��e���a������Wx���$�&�SV�S6c����Ƿl����?�=�?����61�����6�������k��>��q�B����������)��������d!���O��&i���e�i�'?庑�Ͻǿ����m;ܾ�  ?�A ?ۧy?����"���8�� >dW�<Y����뾖����ο���9�^?e��>'�f0�����>¥�>g�X>�Iq>����螾�+�<�?x�-?D��>L�r��ɿT����Ĥ<���?��@�~A?��(�-���^=�E�>]	?�-=>��1�4��.�����>CP�?:�? �X==�V�P��'�d?��=<��E��.⻑�=<2�=��=���b�K>��>P\ �=B�j�ҽ�4>JǄ>�w*�4���]�8b�<z�]>��ٽm���H7�?��N�{m�M�9�F+����=U?r�>���=D�'?��Q��п9	R�UbY?.�?�k�?�:/?"���GT�>�o˾�M?�+?-|b>Ҳ��q�n�5>�̴=@*>M�۾��Q��-=�@�>_WN�pg���6�4�����n���f�F�ƿ$�$�}��^=��ݺX�[��}署���#�T�g#��8fo���轆�h=���=�Q>Ml�>V%W>4Z>gW?��k?�N�>L�>�6�j���ξAy��G�����H�����q��R�ԩ߾~�	���������ɾ�=���=�8R�E���D� ���b�h�F���.?�\$>$�ʾ�M�	�+<"kʾv���|Z��9���>̾9�1�Vn�>ȟ?P�A?������V�j��W��n.����W?��d��6���u_�=�貼)�=%�>���=H�⾪ 3���S�-?!�!?O�ƾ�M��H 4>���,�,=��-?M�?�۫<���>Hs#?�7��}�B�1>Q�!>*�>���>�=�ΰ��⽄� ?&sZ?������܌>*���i�GKV=�> >3RA�h���_>b�<�Ǐ����ѐ ��.<�VM?v"�>2U9���A�(6��f��A�=��{?��?�y�>�Mj?d�A?��n�^��l�Z����2��=�U?��8?=ʱ�; �������J?'�t??��=P�[�t� �B�B���
��?)wm?*(?���CƉ�������S+?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?l�;<��V��=�;?l\�>��O��>ƾ�z������0�q=�"�>���ev����R,�f�8?ݠ�?���>��������=�ٕ��Z�?��?m����Lg<w���l��n��`�<�ͫ=��D"�����7�u�ƾ��
�֪��Y޿�楆>9Z@�V�4*�>�C8�U6�TϿ(���[оKSq�Z�?���>��Ƚ:����j�rPu�o�G�'�H�d���ʭ�>qA>��ؽ�U��q|���7�M�ɻ���>�d��-	�>ݮi��wȾగ��>=�6�>���>ޔ�>��Ľ�Q��r�?��ݾe�̿����x�	�j|I?A\�?��?�*.?�	V��f���:��C���a�+?[p?R.[?>����_���/�j?a��MV`�D�4�6IE���T>"3?�D�>Ք-��&|=">��>�>/�]�Ŀ�ٶ�9���}��?��?�k꾁��>���?�q+?=c�=6��`Z����*��o&� ;A?�2>M�����!�0=��ђ���
?~0?�j��2��Z?��l���5� ������>�>�����S��3�ӽj�L��ى��s��W��?�$�?<��?J���R�Ӿi�1?'��>x��#����w��m�>&=��)>JA����y>��<���L�%K.��I�?��?�l?���汿90>d�?��>m��?�e�<-z�>��=�1���G�=s��>=9]>��
=��?��.?\�>��|����҈!�F�@�/\�I1#�>5��]k>T�?�p?]�={� ��żq���ƽ�̠�p��=\v^����K���V�>�=3>�N>��ɾ^ʾ��?Mp�8�ؿ�i��'p'��54?0��>�?����t�����;_?Vz�>�6��+���%���B�`��?�G�?=�?��׾�R̼�>?�>�I�>B�Խ����Z�����7>1�B?O��D��u�o�w�>���?	�@�ծ?li��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?sQo���i�B>��?"������L��f?�
@u@a�^?*����z��� ���骾�ż+f�=t)>YyI���P�N>��[>��2>�	>��>z>h.�=t,'>��B=E7�=�z��&��������P�R���$�
�%r�u4�b�}�
���������5R�s���F-��?�����u�����=�U?8R?�p?� ?�x�ڙ>4��� E=�z#��Մ=�.�>af2?_�L?��*?jԓ=����R�d��`���A��mǇ���>�sI>F��>.K�>$$�>�+J90�I>l/?>��>�� >8j'=�庄i=B�N>�L�>���>#|�>�C<>��>Fϴ��1��h�h��
w�i̽1�?}���Q�J��1���9��զ���h�=Db.?|>���?пe����2H?%���w)��+���>}�0?�cW?�>��~�T�.:>>����j�4`>�+ ��l���)��%Q>tl?�1f>�w>�3��T8�RP��?����|>�Z6?������7���t��-H���ݾ�J>[��> 7V�{���햿z0�j���z=(;?�y?�P�����@pt���&CR>�\>�!=���=9L>;\b�W�ƽG���/=AI�=�D]><0?�,>���=s��>�_��,�P�g��>�C>�r,>�@?�?%?/������Ƀ���.���v>���>&f�>�)><�J�@-�=���>��b>���⃽a����?���V>��{��^�7(v��w=�㗽���=!<�=�I ���=��$=�x?����y��3Ͼ`��7?�Յ>���~�'��"n�Ls���0̾4��?�@��?� ��M��W�9?9�?N>���1>��>;��>�Ⱦs����E5?>�>���
�!���~>��?��?�ѵ�9ꆿ�n�B��=vi"?���eh�>�x��Z�������u�l�#=V��>�8H?�V��t�O�8>�w
??�^�ͩ����ȿ<|v���>T�?���?O�m�|A���@����>$��?�gY?�oi>�g۾`Z�̋�>�@?�R?��>�9�ߏ'���?�޶?���?hI>���?w�s?;k�>:)x�eZ/��4������wv=`�];Ii�>�U>�����gF�ؓ�`g����j����U�a>ˎ$=��>�.��/��6V�=r닽J��x�f�բ�>y+q>@�I> U�>�� ?�`�>��>w=�o��‾﷖���K?���?-���2n��N�<Z��=%�^��&?�I4?�j[�{�Ͼ�ը>�\?j?�[?d�>=��P>��G迿7~��?��<��K>.4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��tS��FB�>�e!?���>�Ү=ܙ ?��#?~�j>�(�>DaE��9��U�E����>Ӣ�>�H?�~?��?�Թ��Z3�����桿��[��;N>��x?V?sʕ>`�����jE�SBI�5���]��?�tg?mS�1?<2�?�??\�A?v)f>��$ؾX�����>D�!?��/�A��T&��,�?q?�T?{��>����ս��׼����}��o�?�+\?�J&?Վ�i&a�^�¾L�<�E!��EY�.��;��D���>��>� ��kG�=�>��=-bm���6���a<WL�=6��>a�=�&7��玽� ,?(@)=������\���o�}tP��>�|>m��3�c?&*��ۉr��<��4����r�26�?`��?���?^���?_���F?��?�>��?������z̾�&���m������>Yd�>K�2����oS���	���{l���Ͻ�����>�!�>�?q� ?��O>XP�>	��+�&��L�=��ߠ^��y�:v8���.�W��	��<�#��������� |�U^�>������>x�
?�g>k~{>&��>�����>�"R>�>w�>%X>:�4>�>$,<�н�_Q?r1⾋P	�KAc�6��Bm?��?}��>]����_žF\?:��?�?�?�>8��w�'�}�F?�d?�f�ݫ�>�K�>AU>��F>їV<�CľD�þ]X�9?|9��0���^�����~�>�?�x0=C����ߑ����n=$O�?n�(?A�)���Q�e�o�)�W�IS����;h�Ck����$���p�폿_��%���(��e*=͊*?:�?�������$���"k�?�ff>���>�&�>�޾>�xI>��	�T�1�� ^��K'�𲃾�U�>[{?҇�>�I?5<??xP?�kL?���>
c�>)4��Sl�>��;$�>��>?�9?��-?/80?�z?�t+?�4c>?~��p���ؾ�
?��?�J?�?߮?�ޅ��tý�\���g��y����y�=v%�<��׽Eu�8�T=_T>�� ?S�-�z1>�^M߾p9>z?�w�>K��>����)ɾB�=&b�>n�'?q�>6վ%��Gd�%<?ڂ?��ݼH�>=Hi>x(�=Վ=s2�;6l^=����=ؕ�<\{���+�=���=�Ų<�c3�m���b�U=��=,��w�>n�?}w�>�'�>�I��]� �=��C��=�+Y>8?S>%->�Eپ$~���$��M�g��~y>�z�?�v�?�Ff=$ �=v��=gs��Z�����E콾���<w�?�7#?YHT?풒?��=?	o#?�>t3��P��Pa��������?�(,?Z�>+�F�ʾ�꨿�3�E�?%^?9a� ���)��.¾S	ӽC >�4/�@~�b����C�Zk�p���7����?J��?�?��6�zo辒���L:��}�C?�*�>t��>���>ܿ)��g� 3��`;>{��>��Q?B�>R�1?�+t?2i?��j>��#�����������q22>d�3?PLz?�?�k~?�J�>�>`9,�-ܼ�����O���l��\j��qS=��@>F4�>k��>�w>)��=�*c=��s���C�<��e>���>+��>~�>�8�=�d�=�H?���>���9����i���W�>�+g?���?6?����5c�fj[��r���>�M�?��?��>�Ȅ�İ=7�%>��y�%�!�>GHl>W�>h�1>�^>1Ì>��!?D�>\^��U<K�H7g��h���
�>s�<?��)��ƿp2q�,�k��ᕾ�<�B�� �c�|r��<Z�:ܠ=�s������q���]�׳��7���	$��'N��h,|�$��>E?�=�
�=Ɖ�=
�<������<�RN=�;}<��=�]p��O�<�-3�70���녽>����< �T=P�ĻS����?�,1?��>�_?�'8>�Z�>�ϰ>�?�}>�v?I�/>����P� ���.�W����� '3��;"�ܦC��7,�-Dc>a=[�>�q>`��=â�q�2>��y��Ӂ��?����<߯�=�ޯ=� �m�>�4>>P�N>�6w?X�������4Q��Z罥�:?�8�>d{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>q��=w�2�T��>��J>���K��B����4�?��@��??�ዿТϿ6a/>E�7>B">&�R�I2���Z�Web�1�Y��!?U�:���˾Z>�>�ż=O߾�Ǿf�$=�f5>�[=��T`\��=�Q|�P�A=��t=�L�>VE>��=�ܰ��d�=�UF=���=oN>#s��b�3�f</�Q�,=3�=�`^>�$>b��>/�>-B?�X?r�>��A�t���E����� R>ª�>p��
�|>=?i�:?�??�QA?x�>��>�$�>��>�~K�ߠ��<	��t��[�>��?�P�?�Y�>r����žt�4�8;�@s���"?/3?pˍ>�n!>�U����9Y&���.�$����{4��+=�mr��QU�M���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=$�����<�vż�����u&�:�+�1�����;r��;B�]<^��;� �=L��>Y\>3$�>�	�=�V0>�O����K����=vs��h�@���c�*b~��w/��5��"B>r�Y>o��\㑿�? �[>Q?>�A�?��u?�{>�X� �վ@���g�vQ�"��=�b
>%J?�7=<���a��HN�=UҾY��>���>
�>��l>?�+�?�1�v=a���g5�ݦ�>�i������t��q�Q&��i����i�c�d���D?`;��^'�=�5~?D�I?�ߏ?��>�[���ؾ�/>Z���o�=�����q���|�?N'?�>�:쾔�D�҉;���7ǹ>=�E���N�~���<0�a_(�����?��>����#�о�#3�wM�������B�mws���>m'O?0�?�ce�|(����N�q��K_���?��f?3��>k?�?�q�����4?~�Pҽ=��n?���?:J�?D>���="���:�>�-	?h��?���?�|s?��?��o�>{��;ź >	���"U�=Z�>���=�,�=r?"�
?��
?�d����	����=��P^��g�<��=c��>Mm�>l�r>F��=�2g=�b�=�-\>b֞>��>��d>r��><U�>m���]	��,d?�£>Tc�>�Wa?:v>ꠟ��ǽ��B�@�/���D��w�S,��zx��#�.���Ur���X�+,?M~ȿp?�Cc>��6�v�2?�����ԽQ�#<�q�>�т�W{�>"E�>,��>͓?���>���>L��>��>�GӾ�~>����c!��+C�m�R��Ѿ |z>J����
&�)��ky��gCI��n���g��j�l.��^<=�6ǽ<3H�?������k���)�������?O[�>�6?
ی������>���>3ȍ>�I�����ȍ�"fᾲ�?��?�Lc>n�>��W?��?Τ1�*3��oZ�k�u��+A���d���`��፿Y�����
��ο���_?��x?oqA?0;�<A:z>Q��?O�%�1쏾��>�/��;��==@�>�,��a�ιӾ��þ�d��PF>��o?�"�?Q?�zV���m��('>ѱ:?��1?'Pt?��1?m�;?ɕ�9�$?t3>�F?�p?�I5?��.?�
?�2>��=@���'=�8��$¤ѽDyʽ�����3=�g{=lPиvV<��=�ץ<���ټ��;�-��=�<�:=��=��=ؽ�>N�]?�K�>Q��>��7?���Aw8��Į��+/?b�9=���_���ʢ�k���>�j?+ �?dZ?�_d>�A�c	C�>�X�>�r&>�\>�c�>�{�$�E���=�I>�X>�ť=�^M�Dρ���	�Ҋ��8��<;&>��>/|>���i�'>o���4z���d>��Q�˺���S�O�G���1�\�v�MY�>��K?6�?��=�^龊(���Gf�z0)?�[<?:LM?�?9�=��۾��9���J�'>���>�5�<��������"��K�:�֝:}�s>�6���ݠ��_b>����n޾͙n��J����gM=�}�:^V=3���վ�;�ϊ�=�
>����� �W���ժ��.J?��j=�p��E_U�~k����>���>�ۮ>l�:�@�v���@�խ���=�=���>^�:>x������G��6�n>�>cQE?/W_?k�?	"��Ns�#�B�2���Hc���ȼ8�?@x�>h?^B>��=G�������d��G���>���>K��B�G��;��U0��Q�$�Ҋ�>Q9?-�>|�?F�R?{�
?d�`?�*?7E?�&�>�������B&?È�?��=��ԽV�T�e 9��F�(��>_�)?��B�Q��>ӊ?=�?n�&?�Q?Ҵ?��>� ��B@����>QZ�>P�W�Ob��^�_>B�J?���>�=Y?*Ճ?M�=>ǅ5��ꢾ�ө��W�=<>V�2?+5#?��?���>|��>L�����=ƞ�>�c?�0�?"�o?��=<�?�:2>N��>'��=���>c��>�?SXO?>�s?��J?��>R��<�7���8��#Ds���O��ǂ;]uH<��y=��3t��J�4��<��;�g��=I������D�;������;���>��>e�˾R�==C�۾K$w�a�>���=��[���;�:���u�(l�>R?);�>%�#�+f�=]��>T�?�����$?}C�>��>����k�䢿�T������>�%U?P>E�k�r�������Ǳ=���?� w?>���a�J�b?��]?=h��=��þƶb���$�O?��
?��G���>��~?p�q?���>U�e�@:n����Cb�v�j�MѶ=�r�>6X�B�d��?�>��7?-O�>��b>�'�=u۾.�w��q��l?y�?��?���?V**>u�n�&4�
U���$��5k^?ڢ�>I���32#?"�pGоԱ���������3����m�������W��Ȋ$�����ؽ9o�=�^?c�r?ajq?�`?�� �m!c�h�]�b ���V�E���h�l�E���D�]C���m���������t�@=�Uf�"G� �?�9?����u�?����ie�����V@`>ܲ���<]�<-м����<�L�=�Fʽ�a#�̿�449?"Ǎ>��>N�7?Z#|���=���%��L���y�>�mc>��3>4>�>D�=�E�<0�E=�}����Q��e��5v>�yc?��K?�n?�e��(1���� �!�2�/�'\��=�B>�_>0��>��W�����9&�T\>�+�r�����w��r�	�z�~=�2?}+�>���>PN�?�?�{	�0l��]cx�?�1�S��<�0�>Ai?O=�>F�>�н�� ����>t}o?���>䢠>�c��H ��}u��[��1��>΢�>t��>�%`>�.:�A�]�O���������;�s?�=�cc?�����7[��*�>7�L?#�c<	=�<t��>�`��-���� ��>��?[�=/y7>��ľD'���|��熾�O)?�K?�蒾r�*�:4~>S$"?��>�.�>S1�?|+�>qþ�eF�V�?��^?	BJ?hTA?�I�>K�=� ���=Ƚ��&���,=؇�>�Z>- m=�}�=���Vs\�w���D=/t�=�μ%R����<������J<���<��3>Imۿ�BK�"�پ�	����>
�(爾w���	d�����`�����[x�����$'�*V�e3c�������l�X��?m=�?�x��>'��谚�m�������ٳ�>"�q�e������k���(����I����c!�Q�O�7$i�n�e�a�'?E�����ǿ����:ܾ! ?PA ?p�y?���"�?�8�k� >�R�<5�����e�����ο����g�^?=��>�
�1��2��>���>۠X>�Hq>���Y螾<$�<��?և-?��>��r��ɿ������<���?��@4,F?��3�w����׽>I�k=ߔ������Z�����Y�>�S�?D��?�(�>�,$�ܷ��K�K?��>Bz�A�����ҽxf>D>ˈ_�gp=�~��'��^��*�T��U�>*D�>���_�!�Ͻ���<UG�>2�/�Q^���ф?�N\��"f��/��W��X�>��T?�v�>�I�=��,?�;H��|Ͽp�\��a?W#�?~��?7�(?�Կ���>��ܾe�M?"6?��>+P&���t����=�W߼ڙ��c�3�U���=���>��>�,�@^�<�N�G�����=j��Wǿ�+ ���$�^�<�#,��P&������M��G�˼攌�`�`.轑�.=½�=��V>l�>��@>�S>��T?r�j?���>��4>J8ٽ9B���k;�g��D���%�ߝ��%�槾�5��ܾj���-���5ƾ� =���=7R�\���A� �q�b�^�F���.?gv$>��ʾ��M���-<\pʾ4���sڄ��᥽�-̾�1�"n�[͟?��A?������V�4��=U����O�W?sO�����ꬾ���=����ۡ=�$�>���=���� 3�k~S�j�/?��?�L�������v$>�F��B=�-?Eq ?�o<��>��!?��5������R>J74>�#�>w �>�H>�󯾁zͽ��?�MT?h����`��,��>;���Q�w��Q=lV>^�/�/�ż	�T>7U<U}�����	����ʣ<�W?��>��)����А�z3+��'=�5w?��?�*�>��j?W�C?��<���ؑR����#�w=5AX?[�h?�> �u��:Ͼ������5?�lf?W<R>�9d���V2.�v���\?0�n?Li?7�`�|�����-���?6?��v?s^�xs�����M�V�e=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�%Þ?��@���?o�;< �W��=�;?m\�>��O��>ƾ�z������&�q=�"�>���~ev����R,�e�8?ܠ�?���>���������=�ٕ��Z�?��?}����Dg<R���l��n��n�<�Ϋ=���E"������7���ƾ��
�����࿼ͥ�>EZ@�U�v*�>�C8�]6�TϿ)���[о~Sq���?M��>S�Ƚ����A�j��Pu�b�G�3�H�ť��m2�>8�=g��<�Y%�CЋ�^���D��%ư>T�mJ�>�剾r¾����	2;�\�>�%?��>�⪽(����ޜ?�n쾧yҿA@��uA���.?�y�?�cj?�Z?�{F=�,���!��z�<��Z?׆?[Om?�ڈ���H�,�=!�j?�_���U`�܎4�&HE�&U>�"3?gB�>r�-�y�|=>9��>�h>?#/�K�Ŀ�ٶ�����h��?���?�o�D��>K��?�s+?�i�8���[����*��j-�r<A? 2>k����!�0=�pҒ���
?g~0?k{�|.��D\?c�U�9G��P�)l���	�>Ǟ��H4����½��:�������ӌG�P/�?�]�?�t�?ȟ����{*?1��>5���<�Adƾ��?\�=j�K>�9��S>�+�jU-�vV>T��?��?&�?0+������>{�?�>�B�?}��=��>9#�=F簾@h� E&>���=�5�l@?֯L?u�>�#�=$c:��.�y�F��zR�,�>�C�Ƈ>��a?*�K?��c>.δ���:�2�!�fh̽8r.���༠K@��S)�
%ཕ�4>��<>�N>fG��kҾ�?Hp�'�ؿ�i��po'�54?θ�>��?2����t����"<_?!{�>�6��+���%��uB�m��?oG�?�?�׾/S̼�>��>9I�>qս��������7>h�B?g��D��L�o��>���?��@�ծ?si��	?���P���`~�C��/ 7���=��7?p0�M�z>���>}�=�nv�ϻ��A�s����>�B�?�{�?���>L�l?��o�H�B���1=XL�>��k?�s?m�o���
�B>U�??�������K� f?�
@wu@X�^?�Wӿ����xʢ��x�7?C>�*{=��/>`�R��G9>�l+>�-A>W	9=�B >*k>>Δ�=~x>��f>�>��#>]�{�#�!��������H09�_�*�����*��G��!"k������8%��l.����hH�� �O���Q�q��=��U?bR?Ap?� ?�x���>�����A=�~#��Є=�.�>lg2?��L?	�*?ԓ=������d��`��eA���ȇ����>�rI>��>�J�>�$�>��N9��I>�/?>܀�>�� >hh'=&u亟_=�N>�M�>g��>�{�>�C<>��>Fϴ��1��k�h��
w�o̽1�?���R�J��1���9��Ԧ���h�=Gb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��p�T�5:>9����j�5`>�+ �~l���)��%Q>wl?cg>/6~>[P2��x6���O��㰾�q>�j7?�����3��Tt�K�H�ej߾��B>>D6Q����Ė�=~�*�j����=��:?�?�b���x��p�z����FS>��a>�=�ʨ=B�N>��j��&ǽ&I����<^_�=�=^>��?.��>�3G=�)�>�b���!x���>" �>��B>wJ4?2�?gkȽ�4�aʳ���q���X>�O�>��!>�-�=3f�  >Tl	?�OD>�#�<	�b���e��s���u>�J�<q�`���P��s�=��ؽ�v�=]�D<6����^���fX={�w?}����T�����Cʽ'#?��>#����U;�����㩿ٝt��[�?��@�ߙ?�x�_]T��I?�n�?UiO��P�=�z�>}Z�>ט-�?���)r�>b��;�1��������=��?X?�?ϻ��F㘿�߄���">~ A?o�Sh�>~x��Z�������u�C�#=J��>�8H?�V���O�d>��v
?�?�^�ީ����ȿ3|v����>V�?���?f�m��A���@����>9��?�gY?soi>�g۾?`Z����>һ@?�R?�>�9�~�'���?�޶?ӯ�?�I>��?�fs?O<�>�	w�:7/�����B����=���;53�>�W>�����F��Ǔ�"H����j�����Ha>�{"=�͸>�$��8����=����ᓨ�O7m�"c�>��q>Q,J>l�>�� ?��>Lj�>}=���:��������K?���?-���2n��N�<Y��=(�^��&?�I4?�j[�}�Ͼ�ը>�\?j?�[?d�>>��P>��G迿7~��E��<��K>)4�>�H�>�$���FK>��Ծ�4D�dp�>�ϗ>�����?ھ�,��bS��FB�>�e!?���>�Ү=ߙ ?x�#?	�j>�(�>5aE��9����E�M��>��>qH?��~?�?"Թ�2Z3�����桿x�[�J<N>��x?�U?�ʕ>B���߃��
aE�<I�1���^��?�tg?�R��?2�?�??X�A?))f>���[ؾ����>��!?�v�v�A��I&�qC�P[?�a?��>y)��A�Խ�yټg�������?�\?�F&?��*"a�&�¾��<��Ye[���;�iB���>�!> ������=آ>�)�=�Gm��6��ZW<��=���>7j�=m�7��q����)?H��=	쫾J�[=B'`�hZ?���>�%�>�u����S?���W�v�)Ƭ�l����Z����?�1�?#�?[���\�V`7?>�? .'?4��>���Y�оξ����׌�������H>�˳>�������ٙ������x��4�*���8	?��>4~	?Rj�>н:>�L�>ZIh���� Ӿ������\�����5?�a�0���j�����Q�әT�'�¾W�l��u�>>\�����>ba?{;>5?>)�>k�<.�>�XF>B�>��>�H>�>؞�=<����Ľ�R?���#�S���4ݖ��D?o�?���>[���ͱ��W���&&?�љ?Sw�?כ�>�~n������,?��,?E���?�؆�0"�q��<%��>�>Qײ>ȅ�>�K?����{�!t$�1�D���>*V ?�ۘ�ģ���9>n���;�n=	N�?��(?��)�g�Q�`�o���W��S�C��(6h�*j��K�$���p��쏿�^��	%����(��o*=��*?\�?���Ö!���&k��?��df>d�>X$�>�>uI>��	�N�1�I^��L'�U���>R�>L[{?���>L�I?;<?)xP?�kL?u��>�c�>�3��m�>��;<�>o�>1�9?}�-?&80?�z?u+?4c>������ؾ�
?r�?�J?�?�?_ޅ��sýPi���g�.�y�w~���=�$�<��׽�Eu���T=�
T>�r?���ր8�nm����g>��5?���>�8�>����O����&�<%��>2?Ό�>����,�r�_��r��>�y�?����	=0T+>"��=Y���Y��6,�=3`���O�=�R����D��<��=!�=.:�:Ժu ��Q�;kr�<wm�>O?�M�>Mi�>pQ���� ��T�� �=r�X>��R>x�>7_پ�����"����g��/y>�\�?4G�?�cd=� �=wp�=?���������]����}�<2w?@#?)4T?;g�?p�=?c#?�9>�,�C��a~��;�����?>!,?���>B����ʾU񨿽�3��?�[?�;a����C;)��¾7 սJ�>�[/��.~����)D�I������}����?f��?�A�{�6��y�ſ���Z���C?�!�>�X�>w�>�)���g�F%�l,;>H��>�R?,M�>=/%?�e[?�mR?���=g�O���Nƚ�f�{���
�g6>?%Ԉ?�֍?,}?%��>��<�'轍z�� +ɾ�� �	�(��uA��
=RQ>B��>���>���>4�6>u,$���%���-�_gd=r>�>�w�>�6�>*qt>��7=˸H?z��>)>����?�ؾ���6&>�|�?�b�?�G?�7»��9��:N�M����>3��?̥�?ܸ?|ۘ���b=Nz�=�l��������>�c�>�i>�4I=�Ǫ��->=�?L|�>��žE\\�ʿC�R�i��� ?7#,?	B1��rȿ%EY�CGi=.�I�#>Ee�J."�Ed�,�H�ł�<�'W�k�ܽ7�������8 |�̧������K־/4�>ܾ[>i��>���>Z�=��=��=��>Ѧ=�*׻U+<�z�@=a}�6=0/��Ԙ���A���<��1������À?D�6?�o/?�(_?�ӗ>߈>)�>Ƥ�>�+�=�?,v켝������F�}3����<��!�ʕ'���p���>f�=��:>e?u>x�!=xY���A>)��y3>���=lT�=��a>�o�=�:F=��,>g�>a��=&1v?����Ι��nI��`�Y3=?��>E}�=l�žLA?��+>QA��A]����	�f\�?�g�?N%�?o�?��i���>������ֽa�Y=͐�d>�%�=�5�p�>D�F>k���������x�?q�@>�A?oG��Hb̿�C>08>xM>^�R�G1���\��hc���Z�Cw!?�Y;��J̾E�>0��=��޾�zƾZl.=��5>�/`=S,��\�2�=�y��r>=&�k=�ډ>�WD>G@�=�`����=�cI=�@�=yO>|,���7�L>+�(�1=v��=b>J&>���>��?<_0?~Vd?�2�>n��Ͼp?���C�>��=�B�>��=yB>}��>��7?��D?�K?鈲>�Ή=l�>��>��,�v�m�0k��ǧ��۬<���?:φ?zӸ>�jQ<'�A�����f>��.Ž�v?�Q1?bi?e�>�Y�������qZ��I�u-�̆�=�5���+=r��=@=��ܼ��=�Ad>=��>CJ�>���>���=v�$>c��>�A�=s��=�>&�`�E�<~�<�͌=��1� =�7�{:Ƽ�o���v����Z�x<)�y��ᶽ`�Y��{�=fs�>�O>���>���=���7�<>�����I��z�=9R��O�A�5e�V�~�˄/�X73��UC>�fP>훒��&��f?]j>��C>S]�?>�r?��>Ê�`|о�'��B i��M�ќ�=b�>��C��;�`gd��>P��о9��>��>��>�l>�,��"?���w=�	�`5�d�>�{����H.��9q�d?�������i�O�պ��D?�E��f��=�!~?Y�I?��?5��>�&����ؾ=0>�C����=d� %q�wk��W�?''?���>	쾧�D��G̾� ��5�>%3I���O�վ��2�0�Y���ȷ��>?���4�оV$3�g��}�����B�Ar�s�>ĲO?l�?Cb��V��GRO����('���o?@wg?��>AL?�<?8��z��n����=��n?���?�<�?v>]��=���
<�>�+	?f��?ٸ�? �s?S{?��z�>���;=� >����NH�=��>Ȅ�=9)�=as?�
?��
?�g����	�P����A^����<�̡=���>�l�>�r>G��=o�g=fx�=j/\>�ٞ>w�>(�d>�>�P�>ƾ����N?���>]7�>qOj?���=��<���=V��<J�c�6Sҽ�dV�Y��)���4đ��8�;� �F��9�(?Lfƿ{�?a�}>�L�`�7?6U�3���">w�u>ǹ��u�>�W�=�0u>5Y�>fv�>�_�>��>��->�FӾ`>����d!��,C�S�R���Ѿr}z>�����	&���rw��OBI�xn��sg��j�M.��S<=��˽<,H�?x����k��)�����]�?�[�>�6?qڌ����ί>���>�Ǎ>�J��g���Xȍ�hᾤ�?A��?܎c>�F�>C�W?�?c�4���0��zZ�P�u���@��{d��`�׍�ᔁ��u
�����`?,y?7>A?��<B�{>L��?�`&�������>�y/�L�:�N�7=]D�>毰��{a��%Ծ�7þ�����H>��o?��?G:?%�T�'�m�B"'>��:?�1?�Ot?w�1?0�;?���!�$?`n3>�F?�p?M5?v�.?>�
?T2>��=eu��X�'=y6���t�ѽ}ʽ!����3=�W{=b�и�
<ڏ=��<���h�ټ'�; ����<~:=/�=��=�¦>ϧ]?�6�>6��>'�7?���pf8������'/?�:=���F��ۢ��z�>�j?���?�[Z?�Nd>��A�9�B��F>lc�>�z&>�\>XX�>��Y�E�M��=NB>�g>�ʥ=&�M�
ၾU�	������<>���>�6}>�ǐ��&>����W�z�{&f>��O��C��̓R�A�G�l�1�9�w�6��>D�K?�?ߝ=����~#f��()?��<?,bM?��?�^�=ݥ۾�9�B�J�*p��>8α<������E.����:���9M)s>��ܠ��ab>���6l޾E�n�.J����xM=��L)V=����վ�*�6��=�
>v���� �l���ժ�C/J?
�j=�q��'^U�m���>���>:߮>��:��v�I�@�����Th�=~��>��:>���\���zG�[:��`�>�l@?�Y?�7�?��н�'V�n�2�e8��k��*�b�Z*�>�/�>9+?�U�<��<{y��\���q�a�^�	?�>���>��d(4�x�QPӾ["�e%�>/�?Z�5>S��>O1?j1:?�%H?#?mI?ͽ�>�g����4
&?�l�?~��=н�Q�Mh8�j�E�$��>��)?�PA���>s�?.�?�&?��P?J�?��>!Q ��A��y�>"�>|W�	��^>8�I?H
�>Z�Y?��?��@>Ch4��w��ȥ��&�=�!>�m2?��"?]?�
�>g�0?����+Ӿ��>�P0?��{?�8q?�y6>���>��q�8�?���>cq>��M?i�"?��H?�qi?�I?w�"?��=z%<�J����K��C��W]=�"�<}f
���<Gp�����
���|<4f=�>�J=��T��>�wU��_�>s�s>q
����0>��ľ�O��5�@>%����O��Eڊ�:�:��߷=H��>��?ժ�>0X#�B��=P��>/I�>���6(?��?�?=�!;��b�5�ھ�K�C�>D	B?���=��l�k���<�u���g=��m?��^?��W�&��>�b?��]?h��=���þj�b����N�O?*�
?��G���>��~?�q?���>$�e�:n���Db���j�SѶ=`r�>0X�@�d�|?�>^�7?�N�>p�b>D&�=Au۾�w��q���?w�?�?���?�+*>_�n�^4��	�J����E?W�>�۾��?W>=�ؽ���ܾ��,��^��Iپ0�w�wz���w��='ým���E׽*o>��?���?�v?�T?��⡀��>s�� j��k�nW����<�d��8�EyX� ����3�����bо�G�'��� B��I�?t�'?c�1���>
�����1k;��C>2Q���X���=����'C=�K^=�eh��.�����b( ?O�>H��>��<?�[��V>�L�1��U7������3>CǢ>!��>!�>�[�:~M/��齆ʾ�B��W�Խi�->��Y?�7?;�R?�j����D��+���#A�Ge��m|��a�=k�>!�'>����὞��=F�/�I��kj���4�9�j��������D?�V"?|��>sP�?i�2?�ʾ��*D����ž��V��Z�>�jP?�&?��>������!�>=m?3<�>p�>�g�!��b|��eӽ�V�>�N�>]�>-_m>��+��"\��o���Ď��9��8�=v�g?�3��x�a�yu�>�VR?��898�W<�S�>�vr���!�+"���>$��3>~?4W�=�;>[:ľS�F{������w)?Y�?����J>*���>O="?c:�>���>���?���>����:�%?��^?�J?!;A?Y�>|�*=I|��!xƽK�&�F�,=@�>�9Y>6Tr=��=.���[������D=S�=a�μN���%a�;=���&#6<�e�<O�3>Ikۿ�SK��پ����4�Z5
��̈� ���d}��}��������>x�Ms���&�q�U��7c�����|l�f��?�6�?Ga�����9�������������>��q��j��竾�8����3�ྒྷ謾�i!��O�+i�~�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@@^A?�o(����[=*#�>�j	?�J?>��0�I��횱�u��>��?�5�?4�H=N�W�<��Ne?f2�;�FG�E�ֻ��=J��=�o=`����J>?�>dO���?��Cٽ�T5>���>�g�x\�-q^���<��^>�ӽ�䗽5Մ?,{\��f���/��T��U>��T?�*�>R:�=��,?X7H�a}Ͽ�\��*a?�0�?���?%�(?7ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=j6�����z���&V�z��=[��>c�>��,������O��I��P��=������ѿĨ6����D��!�=r�=�{N���ݡ�=���S�,��t����=A�>���>0ه>��>H��>N_[?P�%?D��>�Z�>�Sʾ����ȵ{��>c���h����J �<�G��Tѽ��ľ	���Z־i�'��U�f���!=���=7R�h���D� �h�b�R�F���.?w$>c�ʾ��M�Z�-<�pʾd����ۄ��ॽ�-̾�1�%"n�k͟?��A?������V�M���W�?���^�W?5P�ػ��ꬾ��=ᬱ���=%�>��=���� 3��~S�Ѥ/?i?�g�� k���S>�G
�N�i<��8?`
?���<���>�S-?;m�� �j�g>��?>��>�c?X$>��������|�?�:?</���/�1c�>M�߾@y���ݻ�x�=��4�(-�<B��>��ؽ�̇��0<:Խ3q=��T?��>�"��e�-�x��%�h�)=��x?=�?� �>�4o?��E?y2e����cEL�������=�[?��d?��=Ѝ�4Ͼʧ���2?�o?m�t>�A����.���~?��m?��#?Q�X�u�D�O��f#0?��v?s^�xs�����L�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?w�;<��T��=�;?l\�> �O��>ƾ�z������.�q=�"�>���ev����R,�f�8?ݠ�?���>������K��<&ʫ�é�?�)�?c޾�*��i����[� �4�v=������m�]o���D�z�̾G��1�����;轚>�P@g�D=���>l9���/�;�߿v���V��l���~�?z�>�	y��3���S�������^_�W�i�O ��{L�>��>[���N�����{�	r;�4`����>T���>ӽS��%��c���$25<K�>F��>�>�2���뽾�Ù?+e��i@ο-�����߻X?Xh�?no�?�p?��8<;�v�p�{�����-G?�s?;Z?WG%�*:]���7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�u�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?;�>���?��=o��>�/�=�򰾺�.�c�">��=�fD�5|?m�M?2�>R+�=�>9��/� HF��TR��O�ՎC�E��>c�a?fL?�-c>����@/��� ��ν*�1�����f@��*��`��<5>jT>>�1>�.E�`�Ҿ��?Mp�9�ؿ j�� p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>D�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?rQo���i�B>��?"������L��f?�
@u@a�^?*��пo꓿(#̾F���N�=��>�@>ұ<��>�p
��Ix�kp�=�-鼫��>�8�>x�4>HE�=P	>7f>;���N�}q��Ǝ��$�%������ ������t1�ܬ	����ڕƾ������f�����g���w:��=lfT?�%P?Eq?��?�D���>����u]=KF3��z=�ń>/�4?�G?�"&?K�=����e�G񂿌N���V�����>�@G>�N�>���>���>K�J<x�F>!dF>˨�>���=��4=A;1�=��W>>�8�>�5�>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��w�T�4:>9����j�5`>�+ �~l���)��%Q>wl?��f>�u>Û3�Oe8�M�P�z|��j|>�36?w鶾�D9���u���H�ucݾ�GM>�ľ>�D�l�}����vi�:�{=bx:?ل?w6���ⰾ5�u�kC��oPR>P:\>U=Hi�=�XM>cc���ƽH��g.=���=Ԯ^>I�?��2>�Μ=�i�>H�����L�Hl�>�\>%�E>nz??n�&?2�������눾��)[z>�(�>���>-�	>ScE����=��>�c>������y����FYC��OQ>�����FY�8H�s�V=q��A�=b�=b����9��{x=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?��=���?�.�?Á��`Ӿ__{���ǿUG��������>9!�ā���Y�"��A���թ��P��I�I�/�=�~�=�ъ>}�w��s_�,�'����=�T�L��j��>-ð>���>��>�n�>���>Y>�>�y����ڔz=�p�v�K?���?���2n�uR�<Y��=C�^��&?�I4?�p[�s�Ͼnը>�\?U?�[?d�>��K>��T迿"~��k��<��K>�3�>tH�>�$��|FK>x�Ծq4D��p�>GЗ>�����?ھ�,���O��iB�>�e!?��>FҮ=Ù ?#?1�j>�(�>\aE��9��l�E�J��>���>I?��~?��?�Թ��Z3�����桿��[�(;N>}�x?�U?ʕ>t�����w`E�AI�k���Y��?ktg?�U�>?A2�?��??D�A?\)f>$���ؾb�����>G�!?�`���A�s]&�=�?h?���>i��� �ֽ6�˼����L���{?kD\?�:&? �Û`�>>¾���<�$���m���;��'���>�>'!����=��>���=��m�ڣ5�
�q<��=�M�>�t�=��7�|��0=,?��G�uۃ���=�r�;xD���>�IL>�����^?Cl=��{�����x��	U�� �?���?Zk�?H��:�h��$=?�?N	?j"�>�J���}޾:���Pw�~x��w�`�>���>�l���G���ՙ���F��2�Ž�-�!�>��>�?�P?�E>��>]f���w(����eT ���W�!��h�8���,����U���B��tv��ɸ�9�l���>[a��β>m�
?!{d>mJ�>h�>���-	�>�S>%o�> k�>�T>�?>^�>rߡ��ԽQLR?T�����'���辝���O4B?rd?6/�>�i�X���?��T�?��?~s�?�@v>�|h�U++�%n?^?�>���q
?�N:=����i�<�S������1����p��>7R׽0 :��M��if�k
?�.?��O�̾FB׽zY���>���?��?m�=��s������K�[�n����]��u�Ͼs�7��$���9���N�����	_M�8�= "?�A�?+�C���&�����/��Ӝo�r�>�<?�A�>��>��>�7��Jr��WZ���C�<���y�a>
VN?��>pG?c�7?c0L?HL?7�>��>�E��
	�><�;���>)V�>��3?��*?�*?��?̭+?�ns>�=ؽ(�����־��?lZ?E�?�c
?�?#㍾_�ͽ�ϼ(X��G��O,��O�=�ۻ;�׽�:��Be�<5�Y>�d?'��S�8�*z��}�k>h�7?��>f��>E���a����<�P�>f�
?���>e>��	�q�X�����>̕�?�%��/=C�(>�r�=�ޅ�J�����==ʼ�e�=<�y�j�;�v<���=�d�=�TL�>;:c6;��h;�Q�<݁�>��?x��>�X�>����� �U��#��=L*Z>��S>ӌ>�پ�|���(��%�g��uy> j�?-v�?�g=�%�=^@�=����c+��������tA�<\�?\(#?�'T?�? �=?�3#?�m>��@��)R���Ѣ��?v!,?
��>�����ʾ��׉3�ٝ?g[?�<a����;)��¾��Խѱ>�[/�j/~����>D����V��5��?�?UA�V�6��x�ۿ���[��{�C?"�>Y�>��>U�)�}�g�s%��1;>���>kR?^/�>�*O?+�x?�ra?��>"�,�rǦ��.��_`�<�ߋ=V-?��o?.J�?��Z? {�>S�(>���f��q�6����Ͻ'�`� <=��B>�Ό>��>��>�3#>��;Տ���ʃ����=���>��>A�>���>�R�>}4A���D?٧�>`��� ��'���%���o���?���?�H4?
`>&���	H�r�����>���?M��?�r5?�$6� >@���Ƽ���G����>�e�>�B�>:W�=�F=��=U�>
�>o�z��g��+���V��>�B?��>Yƿέq�x�q��ܗ��k<U���{od�y ��P"[�ε�=R����u�����[��V��YL��
е�ۛ���X{�$��>��=G��=���=FA�<�HǼL��<D�H=Wu�<�=yt��	j<ư7���ֻnʇ��3ʺ��g<V�J=zt�K4��&Sf?oG0?P??�PP?a}<>�>^mӽ�e!>��v�.�?4y?>>�Ľs=Ͼ�r_�]D���ˣ�\M����n�0�dRy�'&�>)�+���Q>�V�>Z2!>�L=�<~�z��;⼮=@�����=<��[�=�]�=���=f6=.S->�6w?X�������4Q��Z罥�:?�8�>d{�=��ƾp@?��>>�2������wb��-?���?�T�?>�?<ti��d�>M���㎽�q�=F����=2>q��=w�2�S��>��J>���K��C����4�?��@��??�ዿТϿ2a/>7�7>.>H�R�W^1��$\�k�b�ygZ�Y�!?q6;��h̾,9�>�k�=�)߾��ƾ<�-=�[6>�b=z��R\�_י=�{��e<=v�l=��>ZD>`%�=e���%�=C�H=��=e�O>�t����7��.,�P}4=
��=�`b>�#&>�g�>�?W9?�pW?��>�6�n|վM0����>�ok>#*�>�C彐+�>2�>�g?G2A?wP?�>�4���ȫ>*#�>��!a��+�d���p�<��?��?�? �r>�L׽��Z�-�)���>�:�>I?�+@?��?�&���ܿ��7�l�K�P�ڻ$-�=bS�=	����ɋ�+E=����@(ǽ��7=��>�,�>f>�>,ea>F,>�}>'L�>g)�=W�����7>`㞽�=-=�f�����-� �*>���|���MB��d;�H�o=V�>��4>�j>�	�=���=���>�7>H��>A��=+���>/>=���;�L�[��=$;��$B��3d��E~� /��P6��B>nEX>�y���1���?�Y>Zg?>˃�?�Eu?��>�*�1�վNP��xHe��`S�d�=G�>I=�w;��U`���M�wҾ��>��>YI�>��l>X2,�5?�,�t=Og�QZ5��,�>[���gm���b>q�d>������ $i��]���lD?7�����=_�}?��I?��? ��>-����(ؾ1&0>����3�=-��CWq��s����?!'?���>j���D�=̾�C����>�@I�;P��ĕ���0�y�&�=ѷ�ޤ�>�����оt3�fh��b�����B�Ѵr�KǺ>��O?/�?X~b��e��)O�����Ʌ��?4�g?��>#?�K?�-�����h�����=`�n?���?�+�?��
>7 �=95��t8�>�>?�I�?D�?�ts?�r8�N��>���;��%>0������=M6>�z�=�I�=<�?U�?cZ?�����	����$��a�f��<��=YҎ>+O�>#�v>�V�=}�Y=RV�=X�\>}�>��>�l>���>�H�>����#���%?�B�=	[�>�42?���>�~K=G����3�<�Fb��p>��1��϶��սL��<��+�Z=����J�>PDǿj�?M�Y>�`�J�?HS�96��N>I�V>���� �>E>G>�>}>
��>�O�>��>�{�>�v*>�FӾm>����d!��,C�_�R���Ѿx}z>�����	&����w��YBI��n��zg��j�Q.��[<=��˽<.H�?�����k��)�	���S�?�[�>�6?�ڌ������>���>�Ǎ>�J��i���[ȍ�hᾥ�?E��?�;c>��>H�W?�?Ӓ1�33�vZ�+�u�n(A�.e�U�`��፿�����
����,�_?�x?/yA?�R�<.:z>Q��?��%�Zӏ��)�>�/�&';�@<=v+�>*��1�`���Ӿ��þ�7��HF>��o?<%�?vY?DTV�_B7�=�+>�6?�$0?�at?r�3?{G:?����V�$?B�'>&�?[ ?��2?x6-?�B?XM1>p��=J��;]=A)�����-�н�����(��Պ=�)�=����f�9���<s�6<�0�h_����<:μ/K�<�B�<��y=���=��>��X?���>o6�>L�1?�9��1��P�
�I?�5�=G����A;�@pǾ�u�y�Z>�]?��?��c?T�w>�81�K��.�=�qu>�a1>��<>��>�9�Q���1,���5>�me>�rr=�W;�������z��L=lqK>��>W0|>���'>�|���0z�^�d>*�Q��̺���S���G���1��v��Y�>;�K?��?ʝ�=V_��,��rIf�;0)?�]<?�NM?��?��=��۾��9���J��>���>�X�<�������#����:�l=�:��s>2��jo�Ќ>�۾�jʾ��o�M}R�N���rн$��6?=����=T˾&�u��7=�F�=��꾖 ?�Md��8R��M�M?����+����l�ٌ���>R>�>|�>�H;Ɩ���5��+z��:>g��>�<.>=�<|�پ�H:��Q��c�>D�J?�1e?�mw?>^��N�|��T���(�>8�qEL��?s��>X?P��=Վ9=�sݾ �6��Å�6aZ�׹�>8;�>M�%�gt;��d�����U��I�>!�?&%�=D�?��[?�	?F[?-c?��	?Fؔ>N)��*ܾ�7&?
}�?�V�=0ս.4T���8���E�p �>e�)?JKB�$��>F`?�?�&?�pQ?��?��>�� �d@��Q�>3O�>�W�P@��П`>��J?�ų>�Y?�ă?]�<>��5�ę��@B��R�=Ԛ>��2?�'#?nL?4Q�>Xd�>M0�t����,�>�+?̀?`f?uV<>��>��\>��>ߦ�=FV?Ɵ)?���>T/?�p^?�7?�A�>�L�=���;o>ɽxNνR"�W����A<�v�=�V =���:�ǽ�]~>�4�|`�	�-�����W�ż������=@�>;jO>����)�<_�ѾŅ����@>ϛe=	��7(1�3�[� >�ޥ>!�?h�+>TN���?>�W�>��>�I�fn?��>���>��콴�}�r���qy�%
f>s�>?�R>�"{�Sk��>+P����=�r?x�e?7��U��D�d?�U?<c�� H,�Ź��~l��*羀&E?l��>�Zy�Hֶ>ir?тu?���>�Gr��;s�XΙ��Fe�󒏾��==�P�>�Q�P_e��ˠ>�k:?���>j(m>��=��s:m�&E{��?��?Aũ?Ӏ�?�	o>�_�.�ۿ[`��h���X?Q�>�H���!?u��;�DϾ����Gև��_��e�����鋾Q��h���G{�.�޽�r�=��?Y|p?��l?�[?� ���a���[�g{�ͅW��m��s�S�G��A�pA���l��!��1쾚t����F=�c�Z@�9S�?�X.?�x����>�R}�����o����B>��ྃҞ��h�=[p�G�m=���=��Q�0X*��ᒾ�&?���>���>K�2?Ya�G�2��� �M<,����5>�Ԓ>q�{>���>��<v^�O��e(������'��jg�>av??��<?e�?"3e=�8��J���),�O�g�9И����>T�V>�6�>N���o����vN��0��iw�֛�f�Ͼd��%6�M�?�I�>�0?�|�?U�?*f��Ī�duO�PH�(ē�eZ�>�K?���>���>r,߹/�f��>~��?�)@?���>.Z@�,H�Q熿2��3E?��*?�FB?���>�UȼBoc�U妿b���uپ	�>:��?��о̵Ӿ��>��c?�>`Ҍ>���>A��*�����P<�4��=�n�>И�=&�D>֚�%� ���^��'�)�'?��?	�z��{;�"xd�|w?<�?�w�>�g�?;�>�pɾ8���|�?>�?�2j?:T?m��>�-�=��,=���W" �D t=���>m�0>_A��C�X�8�PF]�=�ǽB)=�Y%>�9�=��ڼ*�=�9=�:�<�Ǟ;���=;�ڿ�sK��gھ�o�..񾨽��L���̪�7��N�h�������hx��6��Z��V��a������}j����?A.�?���� �������S�����2��>w�l�4�Z�4�^	��]��I�޾��d��	dO�T;h�x�g�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��6�"���8�� >nC�<�,����뾭����ο@�����^?���>��/��o��>ݥ�>
�X>�Hq>����螾{1�<��?6�-?��>Îr�1�ɿb����¤<���?0�@jKF?aQ������>/��>� �>��>~B���l9ؾ���>���?���?D弘�K�{m<G�F?�hǽ�9e��^M��_u>��*>����'7���=�.k>�	��r(�b�e� 5>�S�>����!'4��0Z���>>�)�>��_�W]Ƽ�?1S�·b���4�~��V> \?Y��>��=�k'?!�G���Ͽގ^���f?{�?j�?��'?�����>b�վ�K?z}/?���>�p*��Zq�J�=����{�8��޾�
T��c�=���>?T3>�-��,��sR��ϼ���=I�������ƛ:�T�U��>y=0��=
�<��c��o���|Z�$�>�E'��L������=
��>?ͅ> �>���>�?kA?��%?%��>�>Mx.�ua��]�n��=ǮS�z��<��o�Y���B��5ɾp�� ���Ծ��׾��ؾ_�1���?=�Y�;݌� s�m<I�E�0��/1?r�4>�����R�H��=��♖��V �N�ǽQ}����@jh����?@�C?8K���n_��
�/�۽G����J?�A
�J��."��8�F=h�<B�y=�:y>4��=^.ɾ�+$�t�V���?�
?:
ž_���G>_l
�&Գ���$?��?P9C�"�u>�w ?�)"�Br��O�=���=�Z�>���>@<螼�	 ��� ?T1i?������_�� >��+�������%�=���0<Ò@<s	=D���!�R��?�=�+W?s��>�(�a��!����/���+=�ax?
h?: >/�k?T�B?���<�����T�>���=�W?�i?>56����Ͼ�d��Y�5?��d?2K>�n���羄�-�gJ�>J?(�n?9�?�#����}�&����#���6?F�v?hr^��s��Q����V�;�>E[�>���>�9��l�>��>?�#�G��󹿿>Y4�Þ?k�@;��?��;<� �f��=^<?�[�>I�O�@ƾ;}������ۍq=|#�>����`ev�B��_S,�=�8?̠�?=��>��������|f>����B�?�t�?�o𾂴彪����h�ϲ+����Z=�Y��Y6N��3��S7�h@��CJ$�'[��g��=ɽ�>�y@��>�̈́>7��
�߿L�޿�w���%��KD���c?7O�=BY�����F�_W���j���ƌ���󾃔�>�D>�+��F��Lv�����O�=���>V�=D,s>��i����b��߾=�-�>/?F՞>o�K�ih��G�?#o�`̿3`���r*�,J?���?��?�(?r���@j��cA���S=��`?�Kk?~-I?�؉�GZ{�������j?0_��V`�L�4�vHE��U>"3?C�>�-���|=�>��>h>�"/�5�Ŀ�ض�����M��?K��?Co�o��>c��?�r+?�i�&8���[����*��--��<A?�2>���w�!��/=�3В��
?Y~0?�y��-��o\?�uF��id���<�a�G�6��>�b���Ǫ��9e=�0��}`��֡��ƨ��B�?0��?���?��*����-?{ԯ>Ci��dYܾ�]���I>83�>5ic>�!�;�y>����*8�8�.>���?���?Ao�>w���u����=b�v?�$�>�i}?DK*=�?r�>���
XO��=v�=��*�*��>�LP?A��>�:ۼG�5|��I9��P�I#�O�:�no�>�)g?ygK?w"S>����G!h�	������β�� ߏ��ڽ�>����� >�K�>�;9>�y*�d���0�?�H��ؿ"p��6�'�C�3?���>�?$����s�6��'_?��>u�������M�҅�?���?��?�^׾м�>.$�>"�>,/ֽ���q؇��18>4�B?���&��jo�*�>p��?��@���?P�h��	?���P��Wa~����7�|��=��7?�0�1�z>���>��=�nv�ѻ��R�s����>�B�?�{�?��>�l?��o�I�B��1=M�>��k?�s?�Vo���t�B>��?)�������K��f?�
@|u@\�^?!hп��Ä��0�ʾ�3�=�ڹ=�G>����ao=������Ӽ�c����=*��>�*�>��>��<><v>q%(>MȊ�Z�$�0���u����mI���������|��o�KB���������Rh�Լ�Z���,��+g��������|�=�!U?9Q?�p?�T ?����>�O��T��<�'���=�>Ot2?`�J?Ĥ)?!�=F+��=Je�h���'����:��J��>U�J>��>�|�>�B�>쮢��~I>9�@>@�>8��=r!=�	�-=�O>(�>�k�>�=�> C<>�>@ϴ��1���h��	w�̽�?���ջJ��1���8��7����i�=�a.?z{>����>пE����2H?v����)���+��>��0?@cW?�>���T�*;>v��ɥj��`>~, ��~l�1�)��%Q>�k?�d>ʺr>}�3��|8��O��𯾞Z|>��5?8���a6��Iu��lG��޾�7O>�5�>�zj�<y�r͕���~�#�i�J��=1�9?�?ͦ��@��Pv�o���l%S>K�O>�W=/P�=��L>9�i�[�Խ��L�-!+=���=l�Z>w�>�^#>dj=x�> x���z��%�>�>8�">]�N?�&?�������J%e������0�>���>\�><O�=&�J�0��=L?��=>!�c���(��ٽ#O�H�r>�M/� l��G�����4���6�>0�=>^K��腾.X�<J~?�y���ӈ���꾖���IfD?�?�@�=�aE<�H"�H���6=��s
�?��@@N�?g	�$NV���?W�?m	��vY�=���>X��>ξ	�K�}�?��ƽꊢ�1C	�k#��G�?�-�?C1��⋿q�k���>j`%?��Ӿ:h�>�x��Z�������u���#=[��>�8H?oV��T�O��>�w
?�?�^�ө����ȿ|v����>6�?���?5�m��A���@�h��>��?vgY?]oi>�g۾"`Z�ԋ�>��@?�R?�>�9�K�'���?�޶?���?͋f>!w�?��r?V.�>Yō�.j6��D���팿�=K���q��>$h>���%*H��ڑ�zq���Xr�����C>1�.=.Į>,޽�ٲ���=U���5���F5�p��>kv>�A>ٔ�>���>�A�>��>`9�<�-����q��ʎ��PL?�!�?����l���<=�={�]�S?'�2?�Z��!̾�ȩ>��\?i�~?�:Y?���>�]�����F����K=�<��J>�V�>�W�>��}��#N>�uԾ�hD���>K�>w�N�%�پ~���	9y�? �>�!?<��>Dj�=0� ?cq$?q�m>4�>-�E�aV��CF����>�5�>�?w�~?�?϶����3����U�����Z���O>�x?��?��>�F�����
�,�`nK�6���́?��g?���?c��?�d??��A?�Oc>Qh��j׾�{����>�� ?�e��`A�'v&�s���?�?���>�����ѽ�K�������It?7\?;�%?�?�a�^�Pþ�<ֽ�~:�]<��-�>�>>(���%�=a6> z�=�tg���6���t<��=4��>y��=�G8�����0*?��X�U��W^=��r�k�E�eC{>.I>�|���a?�?��w��o���c��,C=�N?�?�j�?�y�?l!���e�8%;?�&�?�?v�>�����ھ?]޾	�h��>z�����>�L�>��ּe�ھA�����������nݽ)A��(��>���>?�?�L�>ԗ'>�X�>P��/`��~¾�2پ��T���4�Ѷ�G���:��g�0�ܱ�;�uT�/O%>�|ҽ6��>t�?�>5�>���>#��X>�L>��>�X�>H�n>PԐ>W�;>���Zc�=KQ?)���`)��*꾵s���LA?n�c?vR�>`�c�k����� ?|X�?�?�p>�;g��z)�RO?���>��|�M`
?��=9i���G<V��K���0��s���b�>Q<Ƚ�^;���K��a���?��?])�Ѐɾ��׽Iy��2�&>�ۂ?��?C16�V-r�Fp��D�~��n�/Q �W痽wX�n	��kr�����?��f-��ċk��1�8-?��I?�R���¾/f���\�WW8��>`!?�[m>��>���>jxƾ���AB��2�����h��>�G?���>8_B?p�>?�}:?�3U?nx�>
�>����0?�B��p>1��>
.?�?:2?��?�;!?g�<>X���t0���U̾��>��?�w?�T?Fb�>�W���|��9Rܽ:���sU��$�k��=N�=����E���;}�O>��?�[���8�.���tg>w8?��>���>Qr��!vv��m�<ݎ�>�=?V�>�� �Ŷn��9	����>v�?�����z= #>9��=؃��7U;�D�=�ꧼ��=w5<��7��ݵ<j��=L}=|�U�~<�;b�;������<00?�;R?8��>��F>�о]�$��w�$1T>��>�y�>�]b>��(�G&z�W&���^s�&MD>҅?`(�?�Q�=��=q�H>[���Xuվk�����;:�(����>v�A?�FI?��?i��>m ?G3/>ۊ�懝�8Y��	�<?H",?��>�����ʾ�𨿘�3���?Y?q<a�����9)���¾��Խª>�[/�^-~�;��D�)W�����u��қ�?%��?`A�v�6�}y�ʾ���Y�� �C?, �>�Y�>M�>+�)�?�g�u#��2;>��>�R?��>d�K?�v?�_[?H�E>2RA�����DE������A�=:E@?bM�?���?%tj?�*�>NA�=WQv�',��F�F|)�;
������=͆m>SK�>���>���>���=�P��򤩽��H�QI�=�]>7V�>Ȟ>*�>���>l)!=K�E?���>�������B���f{��/U�sys?l��?N�)?���<�� �<�O�����L�>��?D��?�/-?�8,�E��=u�l"žV.�>?�>��>3��=���<{=>��>�>i����()�^9��?�-??��=;���v�TN��I��'Y�=��>GW�=*�>@��IT�>2![�4�n��쨾�8/���1��Jc���8�3m�{s�^��>���=Y:�<ω%=#!I=N���S"�D'�Uz�==*%�J�˼�<X=Igs= ���f�RA���;Z=r-��g}\��!˾�p}?�XI?��+?nD?o�y>��>xG4�\�>�,��p?K[V> %Q�Z���,�;��������9ؾ��־1d�l����=>�~O�K�>"�2>K��=��<Y��=6jt=���=gx��t=N��=��=�ˬ=�T�=5>6[>�'w?��������4Q�����:?Ak�>Y�=I2ƾ3@?M�>>Q<��L���K8�w<?P��?�N�?S�?��h��_�>�iҏ���=V睽�Q2>x��= ;2��p�>VgJ>�l��7���s���/�?��@�??׋�ɑϿF@/>�q>[eb=�uS�F� ������$�Ѹʽ��?�����Ѿ��=Ud=�j������'��=�:�=~k*>W=ѽ�x]����<��<�
�=���=���>���>l�e=�������=�t��.�=y��>ۑ"<�T#�(|Q�~L3=ö4<�[>�r�=��?��*?�??N�R?bʣ>b奾�Ӿ���."m>3y>o�>ޟ}>��J>�&�=�C?�M?K*>?y��>{ϸ���~>l��>|���Â� O#�N��������O�?=��?zC�>}]���>�%�.��?C�p����v�>FX*?��5?I?�(
�zӿ�';�F2Z��i����O=�,�^��|���a�U���S��A$>���>�ޑ>|hj>�u>�=Z>А�>u��>�=3V=:]>aD=x#t=�]��r=hԆ����=���x��<��=��<�$7=@�H=m�>���=/�=�w�>|�#>�o�>��=�Q���(4>s����VC��b�=�)��d�>��b�¥y��U'���,�-	=>��U>��u��Ϗ�": ?�J> @>��?�y?�(>`� �
gʾ�O����y��sI���=�>�6��:5��2]�a�Q���Ծ�Q�>)[�>�Τ>�y>
F(��Y>���U=�l�2����>fO����Kc��Ap�����54����h��j���B?����1�=?x?}�F?��?���>�m�!�о��>�ш��c	=��F�l��#���~?�]&?i�>�Q���D��)̾�Ѿ���>�3I�#�O�����z�0��: ��ɷ�z��>�Ϫ���о}%3��h������U�B�1Er����>_�O?t�?u?b��O���_O�&��Y����h?�ng?'&�>T?0?b��u�
{����=��n?1��?�8�?�>�=L���o�>�W�>aV�?��?wVU?�ս�{�>��!����=>�w�m�;�ډk>#ly>q�<^b�>.��>���>8��Va�BX�����k��B�*�>�>�[�=���=t:��hP�1�
>l�{>U�>���>���>qG>�ȾE��ܴ�>l\�>fړ>��4?��>kW�=S����<����֭�k>�{mG=�N0>n>譞;	>=����?�񛿡�I?4й>��Pa�>��p�F���=�ӥ>��f�>�6&>~6�>�!f>懘>u�'=F�#>k�=0�Ѿm�>�|�� !��5C���R�=�Ҿvx>Y���'��&�Y��$H������|��j�_g����=���<i*�?�. ���k�wa)�0��1J?�ߨ>b6?�׬��Ҋ>���>׾�>����R`�� ����$ᾧ�?��?N:c>��>:�W?�?�=1�x�2�_Z���u��A���d�!�`�Wݍ�����O�
�U����_?Y�x?�qA?i��<E/z>F��?(�%����
�>!/��;�W�;=�	�>�)��n�`�ޤӾ;�þ���kF>Y�o?�?V?V��v��`�>Ұ5?j0?I9t?p_3?f�:?08�Z ?��">��?�	?�2?u�.?�a
?��3>b�=.���=��y��Y����ǽ��̼���<�%=� ����B@=9/=��JR���=C�=���<��@=�%�=3��=�Ĥ>�Z?9+�>`��>>�6?�@�Z7�덲���3?�>=5#z�D샾����Uf�����= d?�X�?7|V?��g>��@�tEK�k>	��>�C>>�X>Ȳ>:)�רE�/b�=&��=ۢ>h�=��0��mX��������5j�<�5>q�>��E>kپ���B>�wҾ��d�2q>:Ku�N`��{�4�q\�x���'u�
<�>s�>?vr)?���=?�޾@%�gN�4?�E:?�uB?tz?�Hl=�Z�^%��9M���\���>\͛��H
��֡�G����<�PE��f>���������a>"p�ۼݾn�~J���羞�J=����pP=�k��վ�X�v��=�[	>����k4!��������I?��l=>#���"U�T6��;L>�>�>5��>C:���x�ς@� >����=H�>,d;>�0����G���ڃ�=�YD?�?�?5u?:���C!��35���),��E�GOg�O�$?i��>��	?F޴��i����)-�������~��>�=�>��}B'��#ӾC~��[�]]�>�?Џ?U2?o7 ?�H�>!XF?�?ܷP?��?�BA��V�&>?&Z�?c�=���P�$�/��M���>~�@?
���J�>�M?e#?�i?�5/?��?�>A|꾋�T�Aޚ>=]�><�Y��Ӵ���$>3PK?+,�>�fX?Ɂ�? ��=.G#��Ȗ��L���t>M^">`?*"?�NF?�B?Ò/?���ш�����>wSN?��:?.x?T�q����>oQ�>#7=������=b��>��'?��Q?1iN?F�>���>&��<OvA��>����gۉ��`���p=M�=��:=�ۼx�G��*�;*`Ҽz����d� @������T�=?7��d�>�vt>�����,2>�G¾������C>vJ���#����=7�CS�=6I>� ?ψ�>h� ���=7�>8�>���i&?��?�?5<��`�^ؾ��J��{�>GxA?	�=c$m��Ŕ��u�H�o=�n?A�\?��]��e��L�b?��]??h��=���þa�b����f�O?9�
?9�G���>��~?_�q?H��>�e�$:n�&���Cb���j�Ѷ=Or�>FX�J�d��?�>o�7?�N�>$�b>'%�=_u۾�w��q��Y?�?�?���?�**>��n�V4࿾�u���y0?��>���� ?��=c�W�ľ�<Ǿ<|꾐����ܽ�E�Wuؾw�e�x���y��&n�>�P?��?H}?��{?o<¾Ʒl�]j}�ځ���
~��O��)��P
^�-�B��7`��i���&�;�*���ma��|���@�mk�?��'?ca.����>䁘���l;�$B>�s��v\��=xʏ�R8<=C+V=({h��90��/���?N��>��>Cz<?��[��>�N�1�y_7������4>�v�>hw�>{��>=�\:��.�Z���8Ǿ�\���k׽�=��B?�bL?c^?B8��HN�	э��a@�T�b��&��n0$?D�>S��<�ɾ�C�[��!��U�78��3�+�}t���� ���d=HT/?�g ?�� ?11�?�??�M���Q����̾��T�ֽRk4>�
M?b��>�؄>C��=�Ҿ�>�	n?j�>{�>���h� �<�z�dn��e��>J��>��>�p>��(�e[��b����^�6�L| >�Ug?=_��6Kc���>�O?�C�;%j<¢�>��Z�+s#�`��8%���>�,	?/ئ=f�9>ž9����x��F���J%?�k�>�у�~|��>(3!?���>�Ҽ>�I~?2��>x��.��V}>��9?�!O?�MK?���>���=Hs�[���ټ�x.�=߰�>�^>���=���<\�l�n����Oܽts=n�<(���5��cvn<�i��r��=��v��-*>:mۿoCK�D�پ����?
�Y刾���~g����oa�����kUx����f'��!V�6;c�:����l���?�=�?�|���,��J���v���K���Q��>1�q���h����7(������¬��d!�;�O�q'i���e����>����+ſu��S��*�?K�-?�zz?g�
�+�4���E���>��>dI�=Cپ�뗿 Pǿ��Z��Oo?B>�>å����<7�>b.>��>��;>x���H������=�$?~�%?=?��V��_Ϳ��=cZ�?2�@��B?��'�4�y=���>�/?��B>q�<�����]���"�>À�?%��?|	e=4�R�o����Cg?6Z�;��C��Ҕ;���=a�z=6�@=����A>W"�>k��:�A�h�ؽd�">�vv>p�/����� a���<Y~Z>�ڽ�˚�Ǆ?Yb\���e��/��0���?>��T?�=�>�-�=��,?27H��|Ͽ7�\�;�`?f�?֊�?��(?X����Ԛ>k�ܾESM?R?6?�7�>9;&��Bt�A+�=s�T`��=�]V����= ��>��>��-�����{O��꛼���=����Oɿ��(�j�$�i�[���y;g�Ҽ�鵽�ѽC���ˤ�8tH��l����=��=9:>�Zx>�h>鿀>G�W?F�h?���>��/>�y��:���8ҾtJ>�������������"��ٛ�g���ﾰZ���'��:���nh��W/�tp��ʝ����b�R�� ��`M?7��=rg�L�U�G���G�վ�"���"��or���徎5	���Z���?��(?�i��o�Q�k�!��k�A];���a?A�'�o��|Lv���>����:��=�(�>�i1� ^�*���|(��l&?�"?�\ž�%��%">�3g�U��=a�+?��>�iq�	��>�1?Eա����j��=5>���>ׯ�>=m>�5��SkF��?��Z?mX<?Y����>�|��h����<m6>4pi� S����)>9�=1���B���y���lK<m�@?<L�>�k��G�jB`��2��<e:H*y?� ?�&~>iyV?�;?�|>d��H�[�̞�.H'>�Ej?��N?<>�8�ߙ���߳�_�?��b?�{�>�>��I��#7���-�?�Qp?@�?<�_=W�X�T$���|¾k3?��v?s^�xs�����L�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?|�;<��S��=�;?l\�>��O��>ƾ�z������3�q=�"�>���ev����R,�f�8?ݠ�?���>�������˖�_a��p��?[2r?�T���X��29p���1����3ڙ=>�<�
�=���H2a�X>
��/+�����@�=�Ր>�@_H>8S�>8s���;�扗�L�̾L�R��?)/�>Q��`����l�������m�w�b��n��>{r>��G/��R�{�e#;�����x��>#/�4�>��S�8��p㞾a]2<��>B>�>yɇ>���O�����?����ο8���U����X?�^�?�_�?��?�T$<�v�b�z���>��fG?i%s?^
Y?1�&�z�X��7%��j?q_��rU`��4�eHE��U>�"3?�B�>L�-���|=�>���>g>�#/�p�Ŀ�ٶ�2���T��?߉�?�o����>j��?{s+?{i�8��r[����*���+��<A?�2>���e�!�:0=�6Ғ�Ѽ
??~0?�{�d.�X�_?�a�=�p���-�,�ƽ�ۡ>��0��e\��L��ۣ��Xe���Ay����?F^�?c�?���� #�a6%?�>[����8Ǿ:�<���>�(�>�)N>�I_�u�u>����:��h	>���?�~�??j?���������U>�}?0�>*�?���=T�>���=����x�&���#>:��=c@���?��M?��>�D�=�&9�j/�MFF�+ R�F��g�C�؇>��a?�L?lc>�F��G�0�0� ��ͽ1�y���@��1�J�߽�g5>�>>�>��E��+Ӿf?���k�ؿֳ��ن)�c�3?&��>��?{7��y�<���_?;I�>�����AN���W�M��?��?�	?��׾�-Ǽ,�>���>�Ճ>�ӽG襽��B$:>'?B?���P�����o�Y�>F��?c�@ȥ�?PYh��	?���P��Ua~����7�i��=��7?�0��z>���>��=�nv�޻��W�s����>�B�?�{�?��>!�l?��o�O�B���1=:M�>Μk?�s?�Qo���k�B>��?#������L��f?�
@~u@_�^?*��˿�������O�þ���=[��=�GN>e�j�=���<�ц�H����o>Ci�>��;>�KU>A1>�_W>��=���9c!������z����G����';���iҽ@���־& �S�ǾٌǾq�"�t��9gF�a�؁���e���\�=+�U?AR?�p?͛ ?;�x�AT>�����=��#�%�=��>�M2?AoL?t�*?���=ȝ�L�d�:b��C,��#������>�FI>']�>��>O/�>��9��I>��>>�3�>�>0�)=dC��
=��N>:��>3��>3�>��;>RY>ZԴ�T7��c�h��w�q�˽*�?���;�J�Q0��A5��%���%��=xZ.?�>��B1п�-H?����7'�T�+���>v�0?_`W?�>N���6U�.s>�r�Ĭj�Rr>y�����l�Z�)�?BQ>�t?��f>�t>&�3�G_8���P�c?��Q~|>G*6?H���k�8�"�u�K�H�ttݾWM>�پ>=�?��N��얿J�~��li���{={y:?��?r���s����u�-O��2R>�E\>n=���=�]M>&ic��OǽW3H��K.=,��=I�^>6?��'>�=CK�>���������>K�D>��7>�a:?�0?�Q����Ͻ�]���i���>J��>>�>(�?���=��>ܺl>4K;y�C��(
�
�3�i~Y>H V��wb�R̝�kO=.���u >�n�=K��4�;�Bc�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>��>�p��f䈿�{���&=J8�>�I?����Ԭ��gW�.?0�?��޾R����Iǿ5Pu�ƙ�>�M�?. �?��q�W ��vJ:����>��?��S?�&R>0X;U$=�@�>Y�B?�Y?	Ѹ>W�#�/��?�Q�?�H�?D�#>ڍ?�o?E$�>G>�^9I� ���G뎿�,��Q8=���>�i>�Xe@�M$��.�@�p���1���=�D=zm�>(��þ��=�P������@�@�>O>��Q>�@>l��>�>a�>��=i2��r��w����K?���?,���2n�O�<`��="�^��&?�I4?�j[�|�Ͼ�ը>�\?k?�[?d�>;��N>��E迿7~����<z�K>#4�>�H�>�$���FK>��Ծ�4D�bp�>�ϗ>�����?ھ�,��8R��HB�>�e!?���>�Ү=�� ?��#?ןj>��>(YE��5����E���>Ĳ�>�C?�~?v�?�Ĺ�'X3����e㡿��[��[N>B�x?�P?ӹ�>x���������C��	I��ݒ����?F[g?��*?�2�?'�??��A?Tf>Ǒ�ؾi[����>n�?��'���8���,��ǽ�t?�?���>d�C<7"��O�[#����m? i?��0?:nɾ�<�d�� E
<|���,&<h�<�����g>�>��ӽ��=R/>�3ݺ�8��8�7�:���\�(=�^H>Q_�=0E���E�=,?��G�+ڃ���=[�r�uD�m�>cLL>@�����^?�v=�~�{�����w��U�� �?c��?Lj�?j����h��#=?$�?�
?�#�>xF���~޾���Ww��~x�<v���>��>�Pl�
徭���a����E��{�Ž5w>��r�>���>G?$G?�,5>���>Rŝ�1f$����E*ʾ39L�u'��mJ�L3!�����˾e�����,�u��=	��͢>�o���)�>�g�>�Ɛ>�o�>��>�sɽn3=Ѝ>�/�>�P�>�?>V\�=o�y>�ds<b�g��1R?�G��G�'�۫�Ň��b'B?Qd?NP�>l�h�iz��`��ah?���?B�?M�u>/\h���*�"�?�k�>��� 
?Y8=����	�<񷶾�z��z�<A�>[�ֽ�:�xRM�nZf��r
?�F?�/���;9Vֽ&C����>�D�?#\ ?��2���k�^�~�ܛk�wod�u�����e��MR�� ���|����Ե��;ʏ��4�j)��ߓ+?�>�?|8����ξ~͔��p�Q�e��
>M�?;J�>���>ۅ�>���nM#���A�O%�ޘx��+�>p�@?r��>*pA?S#9?��O?4�M?D��>��>ສ�0��>p�=i�>%v�>61?�Y+?$�.?�?(.?8O^>�㽭���iϾ�?4/?V�?x�?<D�>����$�4ټ9��<�U�k/P����=U3l=����	��pe=d>.�?8����7�����	[i>�#7?t�>j��>�ҍ�����;�<���>T�?�F�>. �%�p��D
��>�P�?��S�<�;$>���=��+�B�<~��=>���z=�멼�4���f;�T�=���=�1�;v-<�o'�5)/�Ђ�<o�>�H/?/�>js>7]��j���kr����=(�>ALR>P�">��׾����"g��U>�a�?{1�?�cm=u� >M��=�V���o��uC��w!���~=a�?F>?R�=?�M�?4A?��?���=*���L�����˂z�s�?� ,?}��>���)�ʾ��͉3��?�[?�<a�����;)�v�¾��Խ��>�[/��/~�����D�-ׅ���������?࿝?�A�1�6��x�俘��[����C?�!�>SY�>��>H�)�N�g�*%�2;>Ɗ�>YR?c�>��O?�3w?�wU?N>�hK�y����������@>��Q?�{?oҊ?��l?^��>0�>.RY������K�a�gu��e�=ݸr>��>��>�ɣ>��=�l���~��t�I�V=_\D>�>` �>���>�>��=5�D?E��>5'��|8�#
���U���lR���q?�K�?P2+?9:�<���V<C�����W��>)��?Pɫ?Dy)?MY�o��=�տ��[��n�v���>���>f�>Fs�=��S=� >���>��>�R ����GZ5��Q����?lnI?"D�=SnϿR{y�Z�Ҿ����ӽ����x��}��=�T���z�s����I��3.Ⱦ�Ǌ��h;��ξ{gվ�A��1�p4?b�<,>�>7	ａu���g==�Ͻ�~l�&;>�{ؽ�Z�=�0�<R�;��Q1�O��=��=�c=�
�<��˾hZ|?I?^r,?,+D?�)w>(4>]�B���>�i���?�tQ>�_�A�����<�R��������ܾ�پ�>b�����y�>�OH��!>�=3>���=U�<��=��J=��j=R�����:=���=�:�=Gޤ=��=�>Z
>�6w?W�������4Q��Z罤�:?�8�>r{�=��ƾp@?{�>>�2������xb��-?���?�T�?>�?@ti��d�>M���㎽�q�=E����=2>s��=x�2�R��>��J>���K��I����4�?��@��??�ዿ΢Ͽ4a/>��8>R�>YaR��R1��wZ�i�_� �W�	�!?iU:��M˾T>��=��߾_Fƾ@�7=E�8>�g=��.�[���=X�~�j�==�{m=	�>αE>�=�q��0߶=/L=!�=`_K>(׻O�>��(�i�3=jE�=v�`>��$>?v�>��?U,?'�\?[�>�9c���ξq�ľ���>� �=�o�>���=k�L>���>�0?�A?}�Q?:Y�>�0U=߽>|�>cd.��~i��s�p)��V2H=&��?'��?M̧>�P;�jL�Rx �#�1���˽*,?��)?y�?���>�U����<Y&���.�7����4��+=�mr��QU�����Fm�'�㽠�=�p�>���>��>0Ty>"�9>��N>��>��>�6�<�p�=�⌻���<� ��l��=5�����<�vż����Pt&�F�+������;-��;J�]<���;	��=|��>uS>��>q\�=-���?a'>�$����L��"�=󖠾��@���d���~�;�.�U�5��:> �M>r}���p���#?��V>�A>۾�?��u?��&>_���TԾ! ���.s��X��<�=�?>~�;�$�8��_���L�V�Ѿ=��>2��>�3�>��l>�,�U:?���s=@T��g5���>������s��3q�|.���i��8%��UD?67��\��=�~?+�I?q�?�	�>&"���ؾ��0>|;��+^=g����q�D�]�?�'?u��>����D�uJ̾�
����>�>I���O�Õ�`�0�_4��η�.��>������о="3�+g�������B�$Vr�b�>��O?�?<b��V��kSO�<��3'��o?�{g?�>�M?�B?]"��+z�bm��-��=��n?g��?b;�? �
>akM>�+���_�>�$�>��?s(�?[?��
;�V�>8'=)-��b��øx����<2fJ>�ۆ>�)�>��>��>�,ɽ�󾙧�|�-������gA����<K�>ե�>PJk>g��=lX>X�B>��>��>5C�>ď>ܖ�>5g�>bd��,�/ �>�ہ�?�=7#?A׻>D>��(�p�$�5��a.����V�	=\)������Sɒ�4>�E�= V?�uǿר�?��k>%�� ?�U۾�'�*�>l�>D�o�%E?�;�>GRs>g�>�.�>�&6>�j�=E�d>�
��;�=���e1�s|@�GwL�T3��Vi�>>{��a0���(����d�S��Ȏ��/���t�����,����<�ۋ?l���%lg��L'���4�8?�F�>��8?[W��0MĽ^H?>h�?�v�>�n�����'_�������?��?m<c>��>;�W?��?)�1��3��sZ� �u��%A��e�_�`�����ۛ���
�<��>�_?E�x?�uA?l�<�6z>H��?�%�P֏��#�>�/��&;�)L<=/�>&����`�m�ӾŴþ 5��BF>��o?�$�?�Y?	WV���J���>I�;?�5?��m?7�,?�K/?�w3��K?ݐW>Mk�>w�>��'?P2?�?�Oc>Y�>le�:2�=%٠�"H���H���)�ۯ��t�;	w =��;�i�<L�v<���<ܦ�+�<�Ō<�&��R�<��o=���=��=��>Yxp?M �>�=Y>��"?c��m�.����G?��=��d�A����b�ݾ��A=PM?h�?o�Y?5�R>&���z?����=��i> 4>�$L>"B�>
������`ը���<>�P]>^��=.`�ϳ~�4��-��)��=��s>��>5{>d|��D�&>��PUx��e>8EQ����;�R���G�=2�P,w����>$�K?R�?Z��=���=Z��� f� �(?�b<?�gM?_�?��=�ܾF�9���J�	u�pџ>X��<P��l��������:���w:@s>�����T���id>��--ؾ$n���H�\㾵ZE=Y����C=�����Ծ9u�Hb�=�y>���w!�(����w����I?��e=����|�U��=��>R��>�r�>��'���V���?�����ȅ�=���>z�E>Fc���쾑:D�w��x��>��D?:�[?N��?4��f�o�=�����,���H�ݼ�?�7�>*�?Ѫ=>��=�6��@S��c��aL��!�>I�>��iE��ɡ���������>�M?�$>��
?ASO?��?�_^?�h.?�?���>v���p����0(?�"�?�+R=�\S�j�k�6�1���3����>1$?�zM���q>�<?Q�?w?�tO?�z?y�=����-iN��5�>�R�>�|V��h���_=>jw??�>']?�ڄ?�Q>��&�� ����5R�=y�M>!�5?�&??���>��?�W8�{�;���>��?S�?"�h?{c�>C��>�B�>aפ>ɢ\=�S�>|�?1�*?W�D?�?�f<?�6_>v�����.�S���봼.j(>y3�=�6�=hG���r9���+��Z�=͔�>u/���+�j�	=��!=��3��碽�p�>p�s>����61>T�ľ�C���,A>H��@?���׊���:��Ϸ=W��>��?���>�>#�0V�=$��>���>J���*(?�?��?y�;��b���ھ�/K�l6�>(B?�V�=Q�l�����1�u���h= �m?{�^?�,W�+����b?g�]?�0���<���þ��b�t����O?��
?ҊG�A̳>�~?�	r?ܿ�>�:f�A9n�0��CCb�0_k��޶=R4�>}��q�d�YS�>��7?�q�>�hc>���=�۾�w��#����?��?�?���?�F*>��n�x%�[��b˕�[?j?E;��H&?�'�=�8�ȍ��P��,��0ʾ
4��Өi�� ������dI�}s��}@>��?�1l?D�?��b?����k�re���~�_�c��fžz�s�U��1C���+�p`��+��(����þ��=K�y�I�L��$�?*�3?�,a��A�>�]������2����s>g���7���c�=�"�6*
=u�=�d4��p�����e#?m�>��>�6B?�[�H�A�uj2��p=���	�V�>r�>�:>�x�>�S^=�芾����ʾF����,��n�>�7]?��?��[?%�4��2���l�3*�Z2�;��<��=�H?���>S���q��Z��M�.�9?��8R����V2���+{3?�e?>���>���?�?i,��:)���9���a�p�Q��M�=A�o?��?��>E�h<������>��l?��>�
�>}���#b!���{�w�ʽ �>���>N��> :p>Y�,��$\��h��e���f9����=n�h?�z����`���>�R?S[�:*�J<ꈢ>�`v���!�W���'���>�?�5�=��;>�lž���{��D��uC,?�?�����$����>�n!?VZ�>,��>G��?ι�>
f��%�B;�]?c(Z?C�N?�TA?�b�>v��=�c�Y1Ľ��,��=Q)�>d>�=���=��2�_�p�_*$�%�V=ۧ�=�=��鬽����C����|<���;�e.>�kۿ�AK���پ�
�,�:
��刾$���&j�����f��5 ���_x����+'��V�06c������l�8��?x;�?�k���#��$�����������Գ�>*�q�z�w���\��(����ྑ����d!���O��i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�{A?o�(���p�V=3��>��	?\�?>�J1�^A���4?�>�;�?���?��L=\�W���	�le?>��;�G��dܻ��=.(�=�=��y�J>�l�>JU��JA�MGܽ�4>vƅ>��"����K^��s�<}{]>�ս'^��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?X7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=v6����z���&V�}��=[��>c�>Â,������O��I��T��=���ҷ��3��9���=�)>�.�ˍ潮P��+ͽ���8%��v5�0�>�}=O\>8�>(�8>4�>!�J?�\?��>��>��S��l�|軾8Wн��u�.�:����$��������	��	�G����!�`]�����X =���=�6R������� �f�b�2�F�`�.?Fw$>	�ʾY�M��-<�oʾC���݄�᥽.̾��1��"n�͟?�A?����[�V����2V�`���֯W?�O�l���鬾���=ཱ���=l%�>���=��| 3�(~S�j�A?��?c��!��<��>6�����=(�!?��?��<Ԕ?���>����`7�=�5�>�g>0C>�d?�)1>$���B��~?� G?m�=����gϘ>�S羨���e�>��=��Y��!>~�p>�n��� �����=N�RS*�S�\?^֤>�x-��{�|<U��z��DB=l/�?v!@?��E>>�{?&7?B���߾Y&�F�ϾO<�=Zi?�Xa?�P>��{��Ͼ9��e6?C]?em>�e��\F��Kw�\�޾:g�>��[?N.2?R��=���M��/�:	H?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?n�;<��R��=�;?m\�>�O��>ƾ�z������.�q=�"�>���ev����R,�e�8?ݠ�?���>������]�
>�ų����?�{�?�u�@��[)�����閁>����is����T��EP�r"о¼�Ey�� ;�=}��>
@Mב��_�>4W�,������L?����D���R24?�[�>幩����1A����.}��t�"�߽�ݣ>��>�2��N���ϯ{���:�s׊��S�>L��m�>��V�����2�����%<R�>�Z�>wX�>�M�������?���A�Ϳ u��f��IX?E�?�[�?Օ?/_<A*v�"�{���>�G?��s?�Z?���[�Y��8�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?*�a�N�p���-���ƽ�ۡ> �0��e\��M�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>xH_���u>����:�i	>���?�~�?Rj?���� ����U>	�}?�,�>��?L<�=<j�>\��=���A1�Ii#>1�=�:A�1�?,�M?#1�> e�=?	9��/�qVF��WR�2�:�C�/ �>��a? �L?Sb>�x��v�0�H� ��ͽi�1���鼜q@���+����e5>��=>��>�D�:Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�e��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=7M�>Μk?�s?�Qo���i�B>��?"������L��f?�
@u@a�^?*Zr�����aPҾ�Q��̻-�j�j>ƍX>��=Ѹ=�ي�n:��c~'��"
>y>�>���>��>P۔>�ES>F�>4�}�x���J���ߋ���a��
�ʶ��
f�J����u�/�^���
r����e�����L�9�x�1�ȽZs��L�=q�T?��N?��q?���>�ur�Щ,>���ǰ�<�t(���2=Jf�>"�3?�I?J!*?���=%����c�Ci��p��^v��h"�>�s?>���>���>�ΰ>�a;<GR>�MJ>Js>+��=��<�r�;c=��V>���>��>]�>�C<>ő>@ϴ��1��f�h��
w�8̽(�?x���R�J��1���9�������h�=Cb.?|>���?пj����2H?#���{)���+���>v�0?�cW?N�>��a�T�4:>0��ئj�!`>q+ �Ql���)��%Q>ol?��f>�u>u�3��\8���P�_x���x|>�/6?~綾�H9�t�u��H��Wݾ�?M>�ž>��C�0m�������ji�}�{=�r:?<�?[��:߰� �u��8���\R>�F\>�f=,`�=�AM>�Dc��ƽ�G��.=���=�^>}9?��.>��=gĢ>����;$L�Kz�>�B>��+>�KA?	�&?;\&���������$��'x>�u�>��>|�>K�K���=@��>�Qe>6�ؼk�T��W	��M8��/Q>-rV��Rk��i�h@�=�=�����=���=ܮ罯�B�y=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?a|�>���?��?Tw>��Ҿ����ſ�`3�SqW>�{�>3�>>�n����1��㤿;u�����*KM���>�C6=��>o�J�b��R�=4��=�E��O����z>]�>�
>l#�=�>?��?���>"i�="��=Z���Q`�A�K?g��?����m���<�i�=��]�n�?K 4?1�b�5о�Ȩ>��\?���?��Z?U�>����0�������0�� ��<yK>x��>1��>���۱K>3[Ծ�hC���>Bė>7᤼^�ھ�����4r��u�>#a!?���>��=O� ?�#?*n>�C�>˿E�n����G�)I�>��>$ ?��~?�k?�ڼ��4�lT��C��j�\�[G>�{y?�?���>���o�����,�h�W�:���6]�?F�g?�����?j_�?�n??9�@?`sd>$��Ϝؾ$���^f�>a�!?r��vA�;%��_�P?(�?!y�>�S���Q׽;���v�a����?�\?�&?�m���`���ľ�(�<C�(�E���Xj�;H�`�v�>h>8��$�=>Y>�=��m���8�5�t<a�=xؒ>CE�=2�4�zڌ�0=,?��G�ۃ���=��r�?xD���>�IL>����^?el=��{�����x��	U� �? ��?Zk�?_��?�h��$=?�?S	?n"�>�J���}޾6���Pw�~x��w�X�>���>�l���K���ڙ���F��S�Žf�^�65�>���>,�>�?w%�>��>���x���ʾ�	�}3s��:�
5��<$���!v�����WF�f��(�]����>j���?`�>�?�՘>���>���>9֩���>۝>�;�>��u>!s>BI%>L��=�>¼����KR?������'���込����+B?�td?$"�>�i�y�������y?B��?_k�?{Iv>|sh�)0+��b?��>\���j
?��9=������<N�����^↽�z�J��>�-׽ :��M�+Pf��v
?2?:���h̾�:׽L�w�]2�=E�?rG?7�9���l�E ��"{m��/^���m� �@q��$J���z��<���x������P	B��1>�#??a�?m������7��
��Ź_�r�`><�?�7>�1�>l��>�3 ��,;���T���A��̶��V�>��m?�#�>�G?�3?+jK?�xS?�y�>�/�>ڨ����>��>=7��>��>7�5?X.?�72?^?nY,?�||>�齲L��x�׾<?�?�?;�	?i7?��j���۽D�D<����Oh�]��4cO=���&ý�������<B;>kY?����8����ak>��7?��>{��>��	-��tE�<��>'�
?�I�>����{|r�!b��X�>*��?����~=&�)>(��=ko��ҹк�\�=�����ސ=7���z;��a<͈�=��=Gu�����Ȫ�:�v�;�b�<5u�><�?J��>jC�>\@��9� �N��hh�=�Y>gS>�>�Eپ~���$���g��^y>�w�?�z�?�f=��=���=}���U��_�����:��<ţ?1J#?�WT?R��?H�=?)j#?˶>�*�^M���^��P���?w!,?��>�����ʾ��։3�۝?i[?�<a����;)�ސ¾��Խұ>�[/�h/~����=D����W��6��?�?DA�V�6��x�ۿ���[��{�C?"�>Y�>��>U�)�~�g�s%��1;>���>kR?�]�>�W?]l�?+�O?I*>�=��㰿TK���g�Xt\>H�:?�wy?,Ҕ?ӟu?N��>�d�=HbD�I�.����i	�����謾��=�B�>Yf�>�|�>��>��">���u޽2��;��=��w>���>ػ>��>H�z>_值G�N?m��>�NվNf����Ϡ���k�L�?+��?1�?~�I>���9�M�؎	���>���?�Χ? 4?�9��f�>hՀ��_��)��4��>���>�`/>�3!>mL�>���=�E?��>o�q��پ���`�<��	?A"Z?Q��>Rž��*b�P<�n������=J���U�6s���L���I�=ؔ˾)|��yf��*낾���H������Q���A�1��%?�>l��>�">���< ��<5�=�G�=��)=��U=(/��k��� ��z"�>����m��0�<yG�=��D�Ծ�l?/{K?L�$?ZL@?��>�P?>?�;���>���'�?֜F>�R�wuپgB��"���W��j�׾�8ʾ�ZX��祾aL�=}Z�F{>�.>�>�U�=*� >0A=f��=��{=fu=��=[R�=bt�=B��=H��=ش'>�6w?W�������4Q��Z罣�:?�8�>y{�=��ƾn@?��>>�2������yb��-?���?�T�?@�?<ti��d�>L���㎽�q�=?����=2>w��={�2�R��>��J>���K��F����4�?��@��??�ዿ΢ϿCa/>�X8>��>�R�1��F[��7c�s�Z�xq!?��:���̾�5�>9��=߾��ƾ��-=u6>��_=���4m\�g�=��{��=='
o=U�>αD>B��=|'����=� C=$U�=��N>�U����?��,���4=�P�=T�b>�A%>�O�>yX?ʻ?:]a?X�~>�vb��l������n�>�y=$�>�,�=�">S6z>Ճ9?�:?�2?e}�>a��J׷>&S�>]f+�ԁ��s���˾�ͽ���?�˒?��>�qP>���1�ad4�$���W&?ppO?��!?�g�>&���пimS��hb�
����'>6L=�`,��qA�g���x����<^rI<tX�>��>3�>���>Qظ>�Ǣ>���>M�l>(�B=��3>�U<��;���;:�Ӽ�zK��"8<�� f�<�q>"Y�b᪽��<ǀ;Ϳe=���=��>{<>ͬ�>ڏ�=���D/>и���L���=�G��j,B��4d�~I~�=/�rV6���B>3;X>�}��74����?��Y>m?>���?\Au?^�>; ���վ�Q���Ce��US��˸=�>��<��z;��Z`�z�M�_|Ҿ���>��>��>c�l>,��#?�A�w=T⾀b5�V�>^{������"��8q�0@��6����i�}ԺɟD?F�����=: ~?[�I?��?ю�>���d�ؾ^>0>�H����=Y��%q�cb����?e'?��>쾰�D��G̾��}޷>�?I�)�O�z�ޯ0�գ��̷����>������оB$3��g��������B��Lr�;��>d�O?s�?:b��W���UO�w���*��7q?}g?�>�J?A?%��}z�r���w�=8�n?Գ�?U=�?t>�J=w�뽖r�>c��>��?[ő?|�u?��ؽ���>���;�tJ>�c���2>7�y=l}\=��=>��>DR�>��?: g� �������վ����ʧ��v�="Pe>~`�>j�}>�h>=�F�=Ap�=u�>��>1U�>�Pi>t#�>�p�>�θ������?^:>-�9>�32?��>W�*=R�==ҧs="�@쇽�|��F�YQO�^j�=j�=H>c�Ի���>fK���\?���>�t;����>�%��O1��P�>���>����<��>�]>���>ϯ�>��>��>�.�>Hq>�FӾ`>����d!��,C�\�R���Ѿ�}z>�����	&����w��YBI��n��wg��j�P.��Z<=��˽</H�?���� �k��)����T�?�[�>�6?�ڌ������>���>�Ǎ>�J��j���[ȍ�	hᾦ�?G��?�<c>��>��W?9�?��1��3�
uZ�m�u��'A��e�H�`�<፿ќ���
�!����_?c�x?�xA?91�<b:z>��?��%��ԏ��)�>�/�S';��O<=-�>�)����`���Ӿs�þu8��IF>��o?m%�?�Y?�QV�bc���Y>]L<?fH+?�go?�(:?�??�k��)C!??�>m�?�_?K�6?��?y��>R�'>�~�=T�����?=�/���1��vL�P���ň��y�<�J�=���<3��<�&=B&=���<�`Z����<�q��d�D=�<��=g>
��>y]?.�>f�>#8?���7����v	0?��9=��~�Ҋ��飾��mC>n�j?���?��Z?�d>�rA���B�B�>�j�> �(>d�^>d��>���sG��=�4>�6>��=� D��B����	��*����<�!>K��>3|>V��µ'>(t��-z�)�d>0�Q��ʺ���S�@�G���1�B�v��[�>��K?;�?���=�W龡)��=Hf�0.)?�^<?�NM?��?�&�=:�۾8�9���J��0�z�>c\�<l������#��
�:���:E�s>�2���T���id>��--ؾ$n���H�\㾵ZE=Y����C=�����Ծ9u�Hb�=�y>���w!�(����w����I?��e=����|�U��=��>R��>�r�>��'���V���?�����ȅ�=���>z�E>Fc���쾑:D�w��x��>��D?:�[?N��?4��f�o�=�����,���H�ݼ�?�7�>*�?Ѫ=>��=�6��@S��c��aL��!�>I�>��iE��ɡ���������>�M?�$>��
?ASO?��?�_^?�h.?�?���>v���p����0(?�"�?�+R=�\S�j�k�6�1���3����>1$?�zM���q>�<?Q�?w?�tO?�z?y�=����-iN��5�>�R�>�|V��h���_=>jw??�>']?�ڄ?�Q>��&�� ����5R�=y�M>!�5?�&??���>��?�W8�{�;���>��?S�?"�h?{c�>C��>�B�>aפ>ɢ\=�S�>|�?1�*?W�D?�?�f<?�6_>v�����.�S���봼.j(>y3�=�6�=hG���r9���+��Z�=͔�>u/���+�j�	=��!=��3��碽�p�>p�s>����61>T�ľ�C���,A>H��@?���׊���:��Ϸ=W��>��?���>�>#�0V�=$��>���>J���*(?�?��?y�;��b���ھ�/K�l6�>(B?�V�=Q�l�����1�u���h= �m?{�^?�,W�+����b?g�]?�0���<���þ��b�t����O?��
?ҊG�A̳>�~?�	r?ܿ�>�:f�A9n�0��CCb�0_k��޶=R4�>}��q�d�YS�>��7?�q�>�hc>���=�۾�w��#����?��?�?���?�F*>��n�x%�[��b˕�[?j?E;��H&?�'�=�8�ȍ��P��,��0ʾ
4��Өi�� ������dI�}s��}@>��?�1l?D�?��b?����k�re���~�_�c��fžz�s�U��1C���+�p`��+��(����þ��=K�y�I�L��$�?*�3?�,a��A�>�]������2����s>g���7���c�=�"�6*
=u�=�d4��p�����e#?m�>��>�6B?�[�H�A�uj2��p=���	�V�>r�>�:>�x�>�S^=�芾����ʾF����,��n�>�7]?��?��[?%�4��2���l�3*�Z2�;��<��=�H?���>S���q��Z��M�.�9?��8R����V2���+{3?�e?>���>���?�?i,��:)���9���a�p�Q��M�=A�o?��?��>E�h<������>��l?��>�
�>}���#b!���{�w�ʽ �>���>N��> :p>Y�,��$\��h��e���f9����=n�h?�z����`���>�R?S[�:*�J<ꈢ>�`v���!�W���'���>�?�5�=��;>�lž���{��D��uC,?�?�����$����>�n!?VZ�>,��>G��?ι�>
f��%�B;�]?c(Z?C�N?�TA?�b�>v��=�c�Y1Ľ��,��=Q)�>d>�=���=��2�_�p�_*$�%�V=ۧ�=�=��鬽����C����|<���;�e.>�kۿ�AK���پ�
�,�:
��刾$���&j�����f��5 ���_x����+'��V�06c������l�8��?x;�?�k���#��$�����������Գ�>*�q�z�w���\��(����ྑ����d!���O��i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�{A?o�(���p�V=3��>��	?\�?>�J1�^A���4?�>�;�?���?��L=\�W���	�le?>��;�G��dܻ��=.(�=�=��y�J>�l�>JU��JA�MGܽ�4>vƅ>��"����K^��s�<}{]>�ս'^��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?X7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=v6����z���&V�}��=[��>c�>Â,������O��I��T��=���ҷ��3��9���=�)>�.�ˍ潮P��+ͽ���8%��v5�0�>�}=O\>8�>(�8>4�>!�J?�\?��>��>��S��l�|軾8Wн��u�.�:����$��������	��	�G����!�`]�����X =���=�6R������� �f�b�2�F�`�.?Fw$>	�ʾY�M��-<�oʾC���݄�᥽.̾��1��"n�͟?�A?����[�V����2V�`���֯W?�O�l���鬾���=ཱ���=l%�>���=��| 3�(~S�j�A?��?c��!��<��>6�����=(�!?��?��<Ԕ?���>����`7�=�5�>�g>0C>�d?�)1>$���B��~?� G?m�=����gϘ>�S羨���e�>��=��Y��!>~�p>�n��� �����=N�RS*�S�\?^֤>�x-��{�|<U��z��DB=l/�?v!@?��E>>�{?&7?B���߾Y&�F�ϾO<�=Zi?�Xa?�P>��{��Ͼ9��e6?C]?em>�e��\F��Kw�\�޾:g�>��[?N.2?R��=���M��/�:	H?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?n�;<��R��=�;?m\�>�O��>ƾ�z������.�q=�"�>���ev����R,�e�8?ݠ�?���>������]�
>�ų����?�{�?�u�@��[)�����閁>����is����T��EP�r"о¼�Ey�� ;�=}��>
@Mב��_�>4W�,������L?����D���R24?�[�>幩����1A����.}��t�"�߽�ݣ>��>�2��N���ϯ{���:�s׊��S�>L��m�>��V�����2�����%<R�>�Z�>wX�>�M�������?���A�Ϳ u��f��IX?E�?�[�?Օ?/_<A*v�"�{���>�G?��s?�Z?���[�Y��8�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?*�a�N�p���-���ƽ�ۡ> �0��e\��M�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>xH_���u>����:�i	>���?�~�?Rj?���� ����U>	�}?�,�>��?L<�=<j�>\��=���A1�Ii#>1�=�:A�1�?,�M?#1�> e�=?	9��/�qVF��WR�2�:�C�/ �>��a? �L?Sb>�x��v�0�H� ��ͽi�1���鼜q@���+����e5>��=>��>�D�:Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�e��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=7M�>Μk?�s?�Qo���i�B>��?"������L��f?�
@u@a�^?*Zr�����aPҾ�Q��̻-�j�j>ƍX>��=Ѹ=�ي�n:��c~'��"
>y>�>���>��>P۔>�ES>F�>4�}�x���J���ߋ���a��
�ʶ��
f�J����u�/�^���
r����e�����L�9�x�1�ȽZs��L�=q�T?��N?��q?���>�ur�Щ,>���ǰ�<�t(���2=Jf�>"�3?�I?J!*?���=%����c�Ci��p��^v��h"�>�s?>���>���>�ΰ>�a;<GR>�MJ>Js>+��=��<�r�;c=��V>���>��>]�>�C<>ő>@ϴ��1��f�h��
w�8̽(�?x���R�J��1���9�������h�=Cb.?|>���?пj����2H?#���{)���+���>v�0?�cW?N�>��a�T�4:>0��ئj�!`>q+ �Ql���)��%Q>ol?��f>�u>u�3��\8���P�_x���x|>�/6?~綾�H9�t�u��H��Wݾ�?M>�ž>��C�0m�������ji�}�{=�r:?<�?[��:߰� �u��8���\R>�F\>�f=,`�=�AM>�Dc��ƽ�G��.=���=�^>}9?��.>��=gĢ>����;$L�Kz�>�B>��+>�KA?	�&?;\&���������$��'x>�u�>��>|�>K�K���=@��>�Qe>6�ؼk�T��W	��M8��/Q>-rV��Rk��i�h@�=�=�����=���=ܮ罯�B�y=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?a|�>���?��?Tw>��Ҿ����ſ�`3�SqW>�{�>3�>>�n����1��㤿;u�����*KM���>�C6=��>o�J�b��R�=4��=�E��O����z>]�>�
>l#�=�>?��?���>"i�="��=Z���Q`�A�K?g��?����m���<�i�=��]�n�?K 4?1�b�5о�Ȩ>��\?���?��Z?U�>����0�������0�� ��<yK>x��>1��>���۱K>3[Ծ�hC���>Bė>7᤼^�ھ�����4r��u�>#a!?���>��=O� ?�#?*n>�C�>˿E�n����G�)I�>��>$ ?��~?�k?�ڼ��4�lT��C��j�\�[G>�{y?�?���>���o�����,�h�W�:���6]�?F�g?�����?j_�?�n??9�@?`sd>$��Ϝؾ$���^f�>a�!?r��vA�;%��_�P?(�?!y�>�S���Q׽;���v�a����?�\?�&?�m���`���ľ�(�<C�(�E���Xj�;H�`�v�>h>8��$�=>Y>�=��m���8�5�t<a�=xؒ>CE�=2�4�zڌ�0=,?��G�ۃ���=��r�?xD���>�IL>����^?el=��{�����x��	U� �? ��?Zk�?_��?�h��$=?�?S	?n"�>�J���}޾6���Pw�~x��w�X�>���>�l���K���ڙ���F��S�Žf�^�65�>���>,�>�?w%�>��>���x���ʾ�	�}3s��:�
5��<$���!v�����WF�f��(�]����>j���?`�>�?�՘>���>���>9֩���>۝>�;�>��u>!s>BI%>L��=�>¼����KR?������'���込����+B?�td?$"�>�i�y�������y?B��?_k�?{Iv>|sh�)0+��b?��>\���j
?��9=������<N�����^↽�z�J��>�-׽ :��M�+Pf��v
?2?:���h̾�:׽L�w�]2�=E�?rG?7�9���l�E ��"{m��/^���m� �@q��$J���z��<���x������P	B��1>�#??a�?m������7��
��Ź_�r�`><�?�7>�1�>l��>�3 ��,;���T���A��̶��V�>��m?�#�>�G?�3?+jK?�xS?�y�>�/�>ڨ����>��>=7��>��>7�5?X.?�72?^?nY,?�||>�齲L��x�׾<?�?�?;�	?i7?��j���۽D�D<����Oh�]��4cO=���&ý�������<B;>kY?����8����ak>��7?��>{��>��	-��tE�<��>'�
?�I�>����{|r�!b��X�>*��?����~=&�)>(��=ko��ҹк�\�=�����ސ=7���z;��a<͈�=��=Gu�����Ȫ�:�v�;�b�<5u�><�?J��>jC�>\@��9� �N��hh�=�Y>gS>�>�Eپ~���$���g��^y>�w�?�z�?�f=��=���=}���U��_�����:��<ţ?1J#?�WT?R��?H�=?)j#?˶>�*�^M���^��P���?w!,?��>�����ʾ��։3�۝?i[?�<a����;)�ސ¾��Խұ>�[/�h/~����=D����W��6��?�?DA�V�6��x�ۿ���[��{�C?"�>Y�>��>U�)�~�g�s%��1;>���>kR?�]�>�W?]l�?+�O?I*>�=��㰿TK���g�Xt\>H�:?�wy?,Ҕ?ӟu?N��>�d�=HbD�I�.����i	�����謾��=�B�>Yf�>�|�>��>��">���u޽2��;��=��w>���>ػ>��>H�z>_值G�N?m��>�NվNf����Ϡ���k�L�?+��?1�?~�I>���9�M�؎	���>���?�Χ? 4?�9��f�>hՀ��_��)��4��>���>�`/>�3!>mL�>���=�E?��>o�q��پ���`�<��	?A"Z?Q��>Rž��*b�P<�n������=J���U�6s���L���I�=ؔ˾)|��yf��*낾���H������Q���A�1��%?�>l��>�">���< ��<5�=�G�=��)=��U=(/��k��� ��z"�>����m��0�<yG�=��D�Ծ�l?/{K?L�$?ZL@?��>�P?>?�;���>���'�?֜F>�R�wuپgB��"���W��j�׾�8ʾ�ZX��祾aL�=}Z�F{>�.>�>�U�=*� >0A=f��=��{=fu=��=[R�=bt�=B��=H��=ش'>�6w?W�������4Q��Z罣�:?�8�>y{�=��ƾn@?��>>�2������yb��-?���?�T�?@�?<ti��d�>L���㎽�q�=?����=2>w��={�2�R��>��J>���K��F����4�?��@��??�ዿ΢ϿCa/>�X8>��>�R�1��F[��7c�s�Z�xq!?��:���̾�5�>9��=߾��ƾ��-=u6>��_=���4m\�g�=��{��=='
o=U�>αD>B��=|'����=� C=$U�=��N>�U����?��,���4=�P�=T�b>�A%>�O�>yX?ʻ?:]a?X�~>�vb��l������n�>�y=$�>�,�=�">S6z>Ճ9?�:?�2?e}�>a��J׷>&S�>]f+�ԁ��s���˾�ͽ���?�˒?��>�qP>���1�ad4�$���W&?ppO?��!?�g�>&���пimS��hb�
����'>6L=�`,��qA�g���x����<^rI<tX�>��>3�>���>Qظ>�Ǣ>���>M�l>(�B=��3>�U<��;���;:�Ӽ�zK��"8<�� f�<�q>"Y�b᪽��<ǀ;Ϳe=���=��>{<>ͬ�>ڏ�=���D/>и���L���=�G��j,B��4d�~I~�=/�rV6���B>3;X>�}��74����?��Y>m?>���?\Au?^�>; ���վ�Q���Ce��US��˸=�>��<��z;��Z`�z�M�_|Ҿ���>��>��>c�l>,��#?�A�w=T⾀b5�V�>^{������"��8q�0@��6����i�}ԺɟD?F�����=: ~?[�I?��?ю�>���d�ؾ^>0>�H����=Y��%q�cb����?e'?��>쾰�D��G̾��}޷>�?I�)�O�z�ޯ0�գ��̷����>������оB$3��g��������B��Lr�;��>d�O?s�?:b��W���UO�w���*��7q?}g?�>�J?A?%��}z�r���w�=8�n?Գ�?U=�?t>�J=w�뽖r�>c��>��?[ő?|�u?��ؽ���>���;�tJ>�c���2>7�y=l}\=��=>��>DR�>��?: g� �������վ����ʧ��v�="Pe>~`�>j�}>�h>=�F�=Ap�=u�>��>1U�>�Pi>t#�>�p�>�θ������?^:>-�9>�32?��>W�*=R�==ҧs="�@쇽�|��F�YQO�^j�=j�=H>c�Ի���>fK���\?���>�t;����>�%��O1��P�>���>����<��>�]>���>ϯ�>��>��>�.�>Hq>�FӾ`>����d!��,C�\�R���Ѿ�}z>�����	&����w��YBI��n��wg��j�P.��Z<=��˽</H�?���� �k��)����T�?�[�>�6?�ڌ������>���>�Ǎ>�J��j���[ȍ�	hᾦ�?G��?�<c>��>��W?9�?��1��3�
uZ�m�u��'A��e�H�`�<፿ќ���
�!����_?c�x?�xA?91�<b:z>��?��%��ԏ��)�>�/�S';��O<=-�>�)����`���Ӿs�þu8��IF>��o?m%�?�Y?�QV�bc���Y>]L<?fH+?�go?�(:?�??�k��)C!??�>m�?�_?K�6?��?y��>R�'>�~�=T�����?=�/���1��vL�P���ň��y�<�J�=���<3��<�&=B&=���<�`Z����<�q��d�D=�<��=g>
��>y]?.�>f�>#8?���7����v	0?��9=��~�Ҋ��飾��mC>n�j?���?��Z?�d>�rA���B�B�>�j�> �(>d�^>d��>���sG��=�4>�6>��=� D��B����	��*����<�!>K��>3|>V��µ'>(t��-z�)�d>0�Q��ʺ���S�@�G���1�B�v��[�>��K?;�?���=�W龡)��=Hf�0.)?�^<?�NM?��?�&�=:�۾8�9���J��0�z�>c\�<l������#��
�:���:E�s>�2���.��qJd>d���߾��m�k�I���澾8Z=�y�`�c=���/־�W}�!G�=ѫ
>"}���f �2���rҪ�yJ?a_=/��IS����!K>7ř>ؿ�>��E�0�n�f�@�k���+�=X��><>^܏�|��e<G�p�~N�>?ZF?�S^?鳄?�n��)is���B�e���]����5�Q?��>dv?[B>?:�=o���6>�af�τI����>�O�>M@��,H����N�!�nO�>+�?q�$> ?�N?-�	?��`?��)?��?�ݘ>���y���w�?���?

<��m�X��Y=?���8�*��>�>.?�Gq�]_�>h��>�b?'?�>?�H?pb>&��k��ۧ>��s>��g�Qm��,�>9�I?B�?��?���?�>�_P�b�־���ʋK>$T>F�6?q�A?�g.?Nޔ>��?.����^��Y?3G?�FP?�Q?8|c>I�T>��8���%>9=*H>O[?/�"?b�!?��U?ƅF?���>e]'=�f�=�ǽ��=�>� s�
�*<C�!����=��I��l�=��<�SG>h�>>�al���L���0=Φ�<�*[����> r>�P��ek5>��þ���)pB>C0��KȜ�|����t<�Y��=�?�>;
?8��>o"��Ô=&Ǽ>���> H�Y�'?�?��?EA9�1a�|!ھ�AG����>�@?!�=�l� ⓿��t�_h=>�m?id^?dgX�����N�b?��]?Bh��=���þs�b����e�O?:�
?<�G���>��~?g�q?U��>��e�(:n�(���Cb���j�)Ѷ=Yr�>EX�O�d�~?�>o�7?�N�>E�b>%�=pu۾�w��q��i?��?�?���?+*>��n�W4࿢C������n?7E�>geپOO?��]����&���C�姾�����ʾg�|�n����"�.���A��>�?�2�?�{?�g?����z��][��>k���b�;�־ݢϾj��
[W�v�l�K�����Q�����l�q2$>1E~�ǡA� S�?޼'?��/����>:����ҕ;2TB>��������Ν=�3����B=�\]=M�g�;.��	��+�?5�>2>�>�=?�H[�<
>�і1���7����a4>���>�T�>���>gl�9�G.�5 �^�ɾOF��?�ӽQC<>Zk?J]P? b[?���u5�,����7��Kڼ$�ξ�W>�7>�Yu>$����T��!1�Q3B��"{���h���g�����=�\6?��>��>���?IM?�|$��Ӿ��m�fb�g-=��>��c?�_�>��>B�N��R$�q��>�l?)�>6��>������!�'|���н���>'ȭ>�>�>0p>K�,���\��z�����kN9�7��=i?h?�C���f`��>L�Q?B��:�Z<���>!�v�`�!����=(�`0>M9?���=�8<>�ž4��@b{�:̊���.?=�?i�Ҿ��,��>��?/*?���>ۀ?A�>ը��Y�P���?hrS?wD?��;?���>JH1>N�ɽ+�V�^SA�K5 >�_z>9�S>?��=���=g�$�)A���"!�)�!>ٗ�=�A����(�=���=u�<���"%>^nۿKK�D�پ]�1"�@9
�Q舾A���c��٭�B\�����]Xx�Ł���&��V��?c�����2�l���?,;�?�m��R%������Z������3��>��q�l@�z諾+��z9���ྑ̬�+k!� �O��i�{�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >^C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾y1�<��?7�-?��>Ŏr�1�ɿc���y¤<���?0�@�>?H1$�ע�?,>���>�
?N|Y>�y���V�����a�>��?���?� �=k�A�m<\�^?P�;D�B��y�;�v�=��(=�+j=w�佳Ry>��>ʻA�+�#���潛�">o�m>��{�L'�X�b�2)o<�ip>y� �����2Մ? {\��f���/��T��BU>��T?�*�>c:�=��,?7H�h}Ͽ	�\��*a?�0�?��?3�(?�ڿ��ؚ>o�ܾi�M?yD6?���>�d&���t�z��=6ἱ���c�㾭&V����=ѫ�>��>=�,����\�O��L�����=W����Ϳ���F�%�}@�F'=9���B~Ͻf�����<�1n��Ω��r��:T�=P��=nXj>ŕ_>@�C>E�\>]hS?5�f?���>�#<>0���P���|���l�;�4���K˽�]�g�����о����V���^�y%��	�E���i=��9�=A6R������ �j�b�u�F���.?�$>��ʾv�M��Z,<�eʾ=���E���Ͼ��%̾!�1�%n��˟?T�A?N�o�V�Z��\���F��3�W?d`�������\��=�N����=�*�>���=���)3�.qS�i/?՝?4���*.��!p1>=����T=�%-?gB�>Wl�<"ח>&�"?T?)�o0����f>�B>u��>��>�L�=���5����p ?�QW?�罦s��Y��>�ۻ�i؊����<�e>����ڼ��G>��I<(����7Y�p�ͽN~�<&W?���>��)�4���M��Q��j�==αx?K�?� �>ik?��B?�p�<�X����S�R�Q�w=d�W?�i?�>�u��)о�[����5?5�e?B�N>��h���(�.��U��?	�n?�X?a_���l}��������d6?��v?�r^�vs�������V�m=�>\�>���>��9��k�>*�>?#��G��຿�BY4�Þ?}�@~��?��;<��$��=�;?q\�>��O��>ƾ{������w�q=�"�>����Gev�����Q,�k�8?ޠ�?���>-���������=%����?�b�?,w���&j<���<k��� ��9�<��=O��,:�����7���Ǿ8z�M���4��·>�W@�v~�>E7�ּ��yϿ����L%Ӿ�lo���?[Ȫ>DνZ+���6l�7x�Z1H��sH��9���֕>��s>���t����d���:����!��>��F=m>��B�9qᾋ�q��6=�T�>Ŗ�>�(�>�$����?�1��RW��ΐ����ϑ\?d�?���?wI?�<
>W���rQ�΀����T?�_v?�DT?(G��,��5�<%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�P�_?�a�H�p���-�K�ƽ�ۡ>��0�ge\�M������Xe����@y����?;^�?_�?���� #�@6%?&�>x����8Ǿ��<���>�(�>4*N>dH_�V�u>����:��i	>���?�~�?Jj?镏������U>�}?�$�>U�?Il�=Mb�>�h�=�ﰾ��,�jn#>��= �>��?��M?K�>Y�=��8��/�ZF��GR��$���C��>�a?e�L?�Lb>���2�K!�8�ͽ;i1��7�S@���,�v�߽$5>��=>�>��D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?[��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�e��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B�}�1=8M�>Μk?�s?�Qo���j�B>��?"������L��f?�
@u@a�^?*����+����H&��}⾊�ʼ��>YW�=F콊+�<������=����>3��>ڀ>���>kV">���=|8>g#|�&�#� ���?m���ڂ�Z���&*���>���%�tW���ܾ־���b����F�;c���$H����>jI?�2E?��n?�?�ۼ�P3>Y�޾�჻l�)���<��>��0?�D?�W ?��=�T���g��8��������>�"Q>�x�>S��>,h�>p�]���,>�+>�w>�@	>k��=���Wx��@�0>П�>�6�>
�>]<>�7>�������2h��Ww���ɽa�?93����I��4���ݍ�l����=�=�G.?��>�����Ͽ-����(H?����w,�D�*�u�>��0?F�W?b>������L��>>9��l�`J>d���k�ƽ)��JP>T�?tnk>(H>0�0�x�7��GJ�����ﺁ>d�:?�g��6���w��gC�׾��^> A�>�o<{��g���R����R�?,=��>?<�?�5���9��SQ\��,���K,>�S>;��<w
>� 7>Z����Ľ�U6��{�<iΣ=�i>��?6>��`=��>=֐���B��(�> �P>�>��:?4�?�l¼܌��T�{��b���}>�#�>8��>*�>czB�$ǫ=kE�>��y>$����Xk�rl��2L��tQ>hi�E�]���k�Wҝ=7���"R�=j�=����F1���=��~?2��	䈿v��`��|lD?+?L�=2�F<܃"�L ��zF��)�?�@ m�?1�	���V��?�@�?�	��I��=�~�>J׫>ξӑL�X�?��Ž�Ȣ���	�Y%#��R�?��?��/��ɋ��l�8>�]%? �ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?.�#�39�?�}?�@�n5��]��'<ɿ�:��̷�>賽>�*�>] �>���Ŏ������hЃ�̘^�z�>M�=��>�p�La���`�>5^b=��@���х�>S�Ҽȅ�^�>�>�4>�P�>���=<`�=�Ef�n ���K?UL�?jg��m�Ͱ�<tr�=#�Z�c!?4?7Z���Ѿ���>��[?���?�Z?Օ�><c��͚�j���c;���]<KQ>k�>��>{�x���L>�`վ:.I�橈>^��>o@/�;Bھ�4����Իۅ�> & ?SX�>s�=�� ?��#?>�j>L(�>oaE��9��x�E�f��>���>I?*�~?��?�Թ��Z3�����桿��[��:N>��x?V?�ʕ>Y���胝�UhE��AI�h���F��?�tg?�S��?>2�?��??)�A?$)f>����ؾ���L�>�H"?�i���0�.$��n�p8?��?� ?Eؒ�e�A�]��7��"���?O�`?P|(?�A˾*�8��tƾ��<؜���x<�f$<�ӱ���=�ic>T��=밻:�Kc=-7>Jm�-��Y��=��^>��>P��=�����>1=,?��G��ۃ���=��r�9xD���>�IL>����^?Ql=��{�����x��	U� �?���?Zk�?P��<�h��$=?�?U	?o"�>�J���}޾3���Pw�~x��w�j�>���>ʢl���F���י���F��T�Ž������>���>�#?�r ?y_O>� �>�I��<'�{������X^��,��b8���.�:������p�#��.�����V�{��y�>4	�����>��
?�1h>��{>E�>h��i�>� R>��>sU�>��W>Z:5>!>��<�2ѽ��O?pj��µ'�Y�ʾ쒤��]??�+c?�H�>H9��������@� ?���?C��?0�>��a�/$��?�G ?&cs�?͉�=������򖤾fe��,�ƅ�� j>vn��~�6��9B��R���
?�`?:� ;��ҾzνF�˛�<G�?���>�)k�d$q�Xk��˴>��y���2P>d:L>�
w��_W��l��욜����uZ����#����>�}'?���?�Ǿ�뾠վs׏�!�y�0��=y��>�q�>�չ>v��>u̼�̱H�w�|���4��2�<�;K?���>�G?�9?Z�P?�L?Z?�>���>d�����>,�p;$y�>x��>v}9?*-?�/?�j?V�*?�b\>���i���_�ؾ�? �?�/?߅?8�?�Ą��ϽL��J ��du�Wg��{=�"�<F�ӽ�L�]�M=O�O>�?�G�I^9�ur��q>'�6?��>��>����hf���s�<��>��
?�>�����p��l
��R�>��?��"�=��/>`��=�����"���=ʱq��ʇ=}��+7���)<��=׳�=�5�;��׺���:�������<u�>/�?x��>�C�>o@��� �C���f�=�Y>�S>i>Fپ�}���$��X�g��]y>�w�?�z�?��f=��=��=M}���U�����Z������<�?TJ#?"XT?Z��?F�=?\j#?��>+�UM���^��l����?h!,?#��>����ʾ�񨿱�3�؝?�[?7<a�����;)���¾�Խ��>~[/��.~����+D����t��8���+��?�?�A���6�ix�ſ��U\��'�C?�!�>�Y�>�>V�)�T�g�,%�1;>��>GR?�%�>G�O?4{?��[?JzT>�8�c*���͙�CH4���!>�@?���?l�?y?on�>��>/�)�j�)e��X��O"�������V=k Z>���>'(�>��>��=>Ƚ�[����>�/k�=�b>K��>㚥>��>v�w>�ۮ<H?�:�>��Ǿ'���ܛ�Qy����ږt?��?m�&?S=a���?��;�r�>�1�?h�?-?H�L�TE�=M�Լ�E���O��x�>k��>"M�>�x==�f=��,>�q�>�I�>-l�����c3���J�?8^D?�r�=\�ſ��q���p�����|e<璾*�d��{���;[�{`�=����u��������[�����tn��N嵾����ߴ{���>�i�=N�=���=�;�<#,ɼ�=�<n�I=M׎<�V=�bp��l<_a8�|�λ��$a�=jZ<�zJ= ���o}˾M�}?�5I?=�+?9�C?��y>�C>q]3���>Ě��>9?�-V>�?P����7�;�a���v��=�ؾg�׾��c��̟�{@>%oI�Y�>1U3>BG�=ߓ�<H�=��r=���=�QQ�]=�*�=B<�=K�=��=#�>�J>>6w?����K����4Q��S��:?�:�>΂�=pƾ�@?O�>>~1������a��-?s��?�S�?B�?�wi��c�>��+ᎽFi�=�Ŝ��<2>L��=��2�b��>t�J>��EJ�������3�?��@/�??gዿ#�Ͽ[k/>��C>O��=]�M�j(���C��!N���D��["?�:�ɾ$�m>�n�=�6־���<=Z:H>Ѝ=�=(�4'_�v$�=jt����!=DF�=x�>�^[>�L�=]CڽzZ�=/C=�#�=��S>_sX<��K�Fwg�]=���=�&k>(
>�A�>ǈ?�2)?Cze?���>�X�\þyɶ���>{��= �>�VW=@>�ɺ>m�5?��@?
.L?�x�>���=y�>P�>!1��o��tپ>˪�QH�<���?>��?S�>
�<�ZW�r���X<��ȽG?�k+?�?E��>�U����Y&���.������F.�]+=�mr�{RU�����m�Y�㽏�=�p�>���>
�>�Sy>��9>��N>�>�>�;�<�p�=����vµ<�������=A���C"�<}uż'��ܰ&�f�+�����ۍ;̗�;)�]<O��;d��=���>$<>��>���=���_E/>1���h�L�+ÿ=�I���*B�u4d�DH~�L/�HR6��B>�6X>����3����?_�Y>�r?>S��?�Au?$�>�#��վ�Q��e@e��PS��͸=X�>� =��y;�)Y`���M��|Ҿ���>{�>*�>BKl>�,�*5?�1�u=-��P5�:&�>1T���-�D�FGq��F������Ri������D??;����=~?��I?c�?��>gw����ؾVk0>NE���=��O�p��ۓ���?'?M��>��C�D��%;*l���ù>�L��P�	��E^1���E�����.�>@7���ξ�3��}���I���B���w�{��>=9P?;��?�`�����qO�r�t���>?�qf?o�>M�?�n?�����~�6耾W�=��n?h��?]{�?�>��K>!���rm�>F�? E�?�O�?�f?�@��x��>4��B=~<�*(�a3>��9>m��=7�><�?�8?Z�>:������O���&�4Te�֏4=��>~��>�K�>M4y>��=�O��n|����7>�R�>ag�>�k�=h�>bS�>%F��:&���??���=�}�>?�$?��>u��=��Q�"H7=�M��3�Zj���j���H��pO=1�l<'$s=��t��/�>����oy�?��c>Է��?�˾���<Z�=i=4>�j��>v� >�˃>y��>���> ��=�T>�X>�FӾo>����d!��,C�Z�R���Ѿ�}z>�����	&����w��NBI��n��tg��j�L.��V<=��ʽ<,H�?�����k��)�����R�?�[�>�6?�ڌ����֯>���>�Ǎ>�J��e���Wȍ�hᾢ�?A��?�Fc>"�> �W?X�?�1�u3��mZ���u��$A��e�ط`�F���e����
���q�_?��x?zA?穒<�<z>ۡ�?\�%��ۏ�1�>e/�u$;�<A<=x7�>�$����`���Ӿ��þ�>��;F>o?� �?`?�HV��HV��e$>>�8?52?�Cs?�2?݀;?��
��H"?<,>\�?�h?��5?�.?e/
?��4>�Y�=�����
=�b��qω��"սz�нzY����I=��=p�����#<+}#=�٢<W��^��X�;� ����<�M=���=f��=�֦>U�]?��>���>��7?���G8�e���R/?o:=^���w�n������>T�j?��?�=Z?/�c>�A�f(C��<>2r�>��&>�p\>
R�>s��J�E���=�]>V�>�ԥ=`�M�nˁ�T�	��?���J�<^�>Y��>2w>𿅽��,>W����l��r>���m����;��EK��"�Q}�����>-G?�� ?{�=c��u�Y�j�?f%8?<U?��~?�A�=Ѿfd<�WWM���B�#�>�	{=xz���w��࣠��D1�|�=+gE>�����Ԡ��kb>1��X޾�n�8J����k�L=X����U=����վ�!�S��=)&
>������ �f���ת��)J?h�j=;n��lU�gq���>�ʘ>�׮>Y:�ɜv��@�����GZ�=C��>=�:>,������qG�7���>g�L?pF?���?��D;��|3�A�������/�p?l�>��?ߑN>ƪH>��þa���|�Xo���>�9�>�5���>1��g��v9�n
���c�>��?)G->�t�>5N?��?�p?�D?��?��>���;T���c�)?A;�?.��=L�<1Ч��\e��}&�*�?l�N?3�;�VA�)�0?&��>�a,?3�C?ջ?j��=����tO����>�W�>�UG�]����z�;)�-?ӫ�>?(�?��?���=�4��Ko���������ٙ;|f�?,�a?��O?[0D?�W?�g�-���0�>A�`?Oq�?t�t?@ut> +>��>�.0?s�K<�v�>^~?�4 ?<�@?�{?/� ?�ģ>���<�H�-���|E;��;�;�ϼ���o��<ҍ=�9�Y�-� �0=�A=�=�9=��ҽ���<G�>��<Rl�>5t>Y����0>�ƺ��큾�2I>�ts�)'��Ά��'�9��=�Ӄ>DE?6�>y���>�=	{�>d$�>����#?f?��?�ꣻ)8\��Ծ��F��Ϋ>Q�@?s��=�Tl�ov��Q�u��GI=��l?8a_?]�E�Ni��W�b?��]?Ra�=���þO�b�Ï��O?/�
?R�G���>W�~?��q?Ү�>f��;n����Db�-�j�fζ=Pt�>&W���d� ?�>��7?�Q�>&�b>�#�= t۾�w�.v��v?��?� �?-��?%-*>!�n��3����������?���>~>���&?O���߾?���%����˧���������d��������1ॾ̬#<�/4>��?�~?
ZY?ir?�J�b@o�ArW�ׅ��CG��f����D`�{�6�@IH������ ��$�W���e�<�����B\�!.�?�(?λ/����>���z@���Ͼ��>�eu��0��@M�<�A��W%�=^B =��z�[2e�Ȟ��$$?�7�>Q��>�&A?c��n.�T?-���@��徨�c>���>�|b>�K�>�%���_���齔a�����ƽR͚>}gi?H�?x�h?k헼چ=������&�O���ᾳ��=��>��>�ƾ_�7��k6�B�M����u�K�����y羅�=� 5?��h>���=��?]�!?��=���)��o��w�;�%ɻҗ$?�M�?��>��->�~_�L�"����>��l?��>88�>y��o�!�	-�AA���>_��>���>��>��)�*O_�r䏿ك��;�9�`
�=Icc?�V����[�^g�>��P?�\�;Y�;@z�>7mK���"�����!,��;	>ʀ?���=`7I>iþ�{
��y�����bY.?:&?	!���.@��D�>ο/?H�?�4?7mn?ƙ<>��־	n>=V?:<?�+?'�F?�1�>�=H�>z����J��0�׼윩>b�>�c=�>�ʶ�����f��=j�.>��
�c%����=��=�6r�j{	�?����v=��ۿ%�K�jܾ��N�����
���!���<���m�9������BY{�����mV��ja��.���h��N�?�=�?tO������+/�������6��9��>�Qn��~h�]�����S�����૾?� ���N�mf��e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�{A?��(�����T=g��>!�	?�)@>��0��<��߰�/B�>�0�?e�?DbN=�W�R�0qe?�#<��F����u�=���=��=s���oJ>L�>'����A�a�۽�5>�{�>F�#�m;��&^�oj�<'k]>��ս����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=v6�ꉤ�{���&V�}��=[��>c�>��,������O��I��U��=}��n�ſ]�%��!�4a�<�}
�?�M�S�潡E���9�yȠ�0|�������=�b�=h�P>�߆>�`>=^>(�U?��f?d�>[>�.ѽ3��Ҽξ��E������H�o��]������쾣Dݾ�?��B�"����ƾ�;B�%_=UMT��V����%��yc��%C��-.?�*%>inξ[�N����޵;�{���s��M��]UȾ(.��h�>�?!1@?����tZ���Ύ;�^���?MW?2������������=���{k�<{"�>UQ�=�߾\�+��Q�(0?�z?U%�©��=�>Hh��O~>�m-?	�>�r=ǽ�>P}?�/�<F�K<.Ps>��u> h�>X��>,�T>�5����X�8
?�l]?ؒ뽐�u�b��>ڒܾ�����=$[>
���	(�T�t>��=���"�
<|�<B$��t9W?���>�)�.4���x�2�ּ�=��?�#?f6�=A3:?�]??�>���QB���;�>�AZ?��m?�&�=_ӭ��ᨾ@���I?hK�?�Z�>�(���p�I �7f��?HY�?/�?�ߴ�v����+������G?��v?s^�ws�����H�V�h=�>�[�>���>��9��k�>�>?�#��G������yY4�%Þ?��@���?i�;<��R��=�;?j\�>�O��>ƾ�z������C�q=�"�>���~ev����R,�d�8?ݠ�?���>���������=D�پ�y�?�0�?>�۾}�i�<���^u��`	�� �=K��=�鏾�Ce�d��j�E��K���0��೾G��=j|�>k�@B�~�/?:f|��͘ӿ�s��>߾�Iﾐz
?v�>���*���9������yOY��k�XYξN�>��>~�������D�{�$r;�C%����>*�v�>�S�z%��������5<��>
��>��>-��v轾ř?�b���?οv�����&�X?h�?+o�?�q?0�9<��v�3�{����-G?�s?	Z?�c%��:]��7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?*�a�M�p���-�y�ƽ�ۡ>��0��e\�N�����Xe����@y����?M^�?i�?ѵ�� #�g6%?�>c����8Ǿ��<���>�(�>*N>rH_���u>����:�i	>���?�~�?Pj?���� ����U>�}?�*�>=�?���=G��>���= ����3���">R[�=�nE���?[�M?~)�>[��=r7��/��dF�G�R����B�C�o �>��a?�WL?�b>�v��	T,�� ���̽��0����*?�=�'�r?ܽ��5>x�=>��>��C���Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�e��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?VQo���i�B>��?"������L��f?�
@u@a�^?*�ӿOۓ��g־�'���G�;�M<�+>��s�ǃ�=�2�Xä�R�-�5a�=�
�>��>][>߀W>��=z>a��u������Rů�F����K=����-����m������΅о�l7���ͼU7(�.[�+ü���~���=],V?^@J?��s?�?pu���>Ad��ߊ���I����=Y��>��/?ZF?�.?�?=�b��t�l��L���U����s�M�>��F>��>Q�>	[�>�f�:�0U>\I>�~>K�>�(�=z;=/�0=73Q>�C�>��>U�>sC<>��>Fϴ��1��n�h��
w�j̽0�?}���S�J��1���9��צ���h�=Ib.?|>���?пc����2H?#���y)��+���>x�0?�cW?%�>��>�T�/:>6����j�-`>�+ �|l���)��%Q>tl?��f>�u>z�3�d8�|�P�!~��yh|>&36?�붾EH9�%�u��H��bݾcGM> ƾ>:,D�'l��������ui�:�{=�w:?��?6���㰾G�u��B��[OR>�;\>�\=�l�=�ZM>�Tc�y�ƽH�vp.=���=�^>��?f�+>x��=�O�>�8��hF�)�>S�F>�>1�??��%?�&��!����}��N'�_�|>��>�W�>oJ>+J����=�G�>�d>�i�𢁽�{�H?�f+X>�{��[���t���\='t���Q�=㧗=���u�6���=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?���>�}?h�j?cc�>e���(���ſ�ӟ���9=ֺd>NU����w>�՟�N���|��e���v��0T�&����4�=G��>�M��H�����>�GL=_����p�h��>,��>��X<��>��?Y��>�,�>5d/>^�7>�tB��*����K?���?���0n�$��<���=��^��&?C4?�[���Ͼ ը>��\?Y��?�[?�e�>���]<��j俿K}���3�<�K>�7�>�E�>�,���GK>��Ծ�DD��q�>�՗>a����Aھ�"������=�>�c!??��>��=c3?{~!?�%~>��>��H�B��.�I����>���>uh?c��?��?�ʾg;�)���H��F�`��=>�t?�?��>(֎�Բ��3�̼K2-��O��-I�?ܵd?���;?�{�?D�B?��@?��`>��Q�ھ�୽!p>T�!?Z�f�A��%&������?�r?���>�0����ӽpǼw��Q���+?��[?�?&?��qw`�g¾ؔ�<��<��y-���#<�&O�I�>�*>���N��=��>�'�=ūn�Z�7��i<�˽=���>0N�={5�M���0=,?��G�~ۃ���=��r�?xD���>�IL>����^?jl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྾Pw�~x��w�[�>���>�l���K���ڙ���F��^�ŽZ�D�>r��>�?C~ ?��O>!R�>�3���1'��x񾏯�̻^�f�%h8�_�.�����Ѡ��0#�ݵ�y<¾��{�1K�>ZR����>��
?A'h>�{>�>³Ȼ|L�>qR>ۄ>�l�>��W>_%5>A�>Ο<%�н GR?������'����5J��_0B?bmd?�A�>dj��t������k?���?<l�?	Ov>>Hh�[+�gd?Q�>h���;
?�/:=����<�-��ؗ�t����ǰ�>9Mֽ�5:�?M�f��i
?5?_N��v>̾}ؽ2���OUJ=܋?mk>?�=���e�o��R�[���a���Ľ?��O*����T��2�������ړ��m��*I,��/�<�1?x̕?Nh�Fn־����_a�a�S�❈> �>��7>���>[a�>�����4���Z�b�`ߗ����>��H?���>=G?:�6?ţM?r�M?V��>Fq�>����.��>�#�;�>P��>��9?��.?�0?5??ԙ*?i�e>{�7���Nپ��?G�? @?nl?z�?5��X8ҽ�r��,�D�{�6��WY^=m��<ٲȽ/�X��s=��F>��?�&�o�8������n>W�7?39�>ϲ�>�Ǐ�\�����<܊�>r�?Hُ>N6����p�_�.��>|q�?�����<��*>���=6�j��\�8���=ĝܼ�ǋ=�YH��6��\ <��="0�=���R�w%�:lI;��<u�>4�?���>�C�>�@��)� �]��"f�=�Y>HS>~>�Eپ�}���$��s�g��]y>�w�?�z�?��f=��=��=}���U�����O���k��<�?@J#?%XT?_��?|�=?[j#?׵>	+�hM���^�������?w!,?
��>�����ʾ��ԉ3�؝?e[?�<a����;)�ߐ¾��Խα>�[/�h/~����>D�U���[��4��?쿝?5A�S�6��x�ٿ���[��{�C?"�>Y�>��>U�)�{�g�p%��1;>���>fR?LQ�>��O?��y?�\?��V>[f9�Tɭ�:q��~���>>�??��?�s�?�~w?E��>&�>-��%㾴���}��3(�z���Z=�Y>׋�>��>���>���=��ƽ\ŭ�|�:�p��=�ag>!'�>@i�>۪�>��x>��<��H?.l?�����c��7��pɠ��Q-��D�?�ߜ?��
?м�k ��y5�3������>���?�g�?�C/?�j,����=,���ľ�/���8�>���>�(�>�>�Ŕ�l �=�F�>a��>��=�i�Lt=�ira�;?\�O?ob>��ϿL�p�#�ľ������[�Ӿ?�� ��<�ٽ��m=��ǾԆ��
۾|�@^�[Ƃ� b�����5�)��>I��=3]>Y�T<_8�<S���>�M9=��M=�_>�F!���=ǭ��Sƍ���<�=��=rYI>�Y¼Ή˾�}?�;I?�+?��C?޸y>�:>��3�s��>ڈ���@?�V>R�P�Έ��e�;�\���� ���ؾ�x׾��c��ɟ��H>�_I���>�73>I�=MK�<z�=Ss=FÎ="�Q�=�%�=&P�=�g�=G��=��>U>�6w?V�������4Q��Z罦�:?�8�>�{�=��ƾr@?��>>�2������vb��-?���?�T�?>�?@ti��d�>K���㎽�q�=_����=2>@��=�2�W��>��J>���K��L����4�?��@��??�ዿ͢Ͽ8a/>�8>G>��R�]1���[���a�L�Y�E�!?
f;���˾���>��=*�޾ ƾe1=)�6>��c=����\�zE�=��|�HH>=�[o=��>��C>���=�����N�=c�I=r��=�SO>a먻��7�R�*���3=��=�Jc>B6%>v��>!?~30?�hd?��>8�n���ξ_����Ë>}�=Ű>�Z�=B>��>��7?�oD?��K?�ʱ>'߅=&�>�'�>�E,���m��3�I���7�<���?��?t��>9�5<� A�����)>�q�ƽ��?u�1?�?�w�>����)��<]?���O����zF��v�=fg��B>s,�>)����?��	��f�>߯�>m��>���>���>֮�>S��>H�M=�A>V߈>�;�>�4�=�S�8զ�'�ɽ�b�<���`H_9)�=K��;�����$=�#k=~X½��=���=��>z<>ܬ�>G��=����C/>߸���L����=�G��e,B��4d��I~�N/��V6�{�B>&;X>�}��A4����?[�Y>�l?>���?YAu?5�>� ���վ�Q���Ce�9VS�Q˸==�>��<��z;��Z`�}�M�b|Ҿ6��>�>�*�>�l>�%,�� ?���u=�4��^5���>����VR�8��:q�8H��(���s,i��7��}D?�:��r�=�
~?�I?�ُ?��>u�����ؾ M0>�(��C=!�7�p�r�����?��&?��>7�B�D��J̾����ܷ>�EI��O���ʯ0�g��h̷����>������о�$3�=g��I�����B� Lr�7��>�O?�?!9b�{W���UO�����,���q?�|g?i�>_K?C@?�$��tz�s��lv�=b�n?G��?>=�?>��=�������>�?Օ�?�ő?l�s?��7����>/�;�&>�ʒ�B��=Sz>џ=ɰ�=?Z�
?��
?����)�	��C��@^�-��<)�=��>�Q�>�q>#��=ݴI=�#�=ezZ>]��>��>6dh>�>�|�>B޾BU8��0?P/N�̮�>i�!?��+>[�]=	q7�	�>瑝���R��L����J���;�VP<[�=V�O>�}#>�o?}!п�R�?|=>H
��V$?��~��<N0>o �>��D=���>����o=�ƻ>ί>���^\�>���=IӾZ|>����e!��-C���R�ǽѾ*~z>	����&�I���{��DI��m���f�%j��-���;=��׽<�G�?������k���)�����Y�?�\�>�6?�ٌ�a����>Z��>|ƍ>K�����ȍ�ngᾺ�?���?�;c>��>G�W?�?ђ1�)3� vZ�)�u�p(A�*e�S�`��፿�����
����.�_?�x?2yA?�R�<*:z>Q��?��%�Yӏ��)�>�/�%';�@<=v+�>*��1�`���Ӿ��þ�7��HF>��o?<%�?vY?ETV�.��:v�>MN/?�8?��x?/@?�??�.��>�?B��=?4?�1?��E?��-?m�?,W~>��	>��r�ߦ>Ny� 4��>�&��E��ڝ�����=���=����F��?ij=:�=� I=�2��p�����:=Y� =�c�=c�y=�Ѧ>�]?�'�>�`�>��7?����V8��q���(/?n�8=
����ӊ��n����6�>��j?���?�[Z?��d>,�A��!C�E>�c�>�&>�M\>�q�>X'��E��y�=(<>t+>�=��L�����I�	�ߎ���=�<>���>W6|>�,��-�'>"��їy���d>�Q�2��Y�S�ǏG�8�1���u�m��>��K?|�?�ܙ=�)����3f�n�(?�j<?kM?a�?�$�= �۾e�9�S�J������>�ޥ<*	�e������b�:�W��:!`t>�~���.��qJd>d���߾��m�k�I���澾8Z=�y�`�c=���/־�W}�!G�=ѫ
>"}���f �2���rҪ�yJ?a_=/��IS����!K>7ř>ؿ�>��E�0�n�f�@�k���+�=X��><>^܏�|��e<G�p�~N�>?ZF?�S^?鳄?�n��)is���B�e���]����5�Q?��>dv?[B>?:�=o���6>�af�τI����>�O�>M@��,H����N�!�nO�>+�?q�$> ?�N?-�	?��`?��)?��?�ݘ>���y���w�?���?

<��m�X��Y=?���8�*��>�>.?�Gq�]_�>h��>�b?'?�>?�H?pb>&��k��ۧ>��s>��g�Qm��,�>9�I?B�?��?���?�>�_P�b�־���ʋK>$T>F�6?q�A?�g.?Nޔ>��?.����^��Y?3G?�FP?�Q?8|c>I�T>��8���%>9=*H>O[?/�"?b�!?��U?ƅF?���>e]'=�f�=�ǽ��=�>� s�
�*<C�!����=��I��l�=��<�SG>h�>>�al���L���0=Φ�<�*[����> r>�P��ek5>��þ���)pB>C0��KȜ�|����t<�Y��=�?�>;
?8��>o"��Ô=&Ǽ>���> H�Y�'?�?��?EA9�1a�|!ھ�AG����>�@?!�=�l� ⓿��t�_h=>�m?id^?dgX�����N�b?��]?Bh��=���þs�b����e�O?:�
?<�G���>��~?g�q?U��>��e�(:n�(���Cb���j�)Ѷ=Yr�>EX�O�d�~?�>o�7?�N�>E�b>%�=pu۾�w��q��i?��?�?���?+*>��n�W4࿢C������n?7E�>geپOO?��]����&���C�姾�����ʾg�|�n����"�.���A��>�?�2�?�{?�g?����z��][��>k���b�;�־ݢϾj��
[W�v�l�K�����Q�����l�q2$>1E~�ǡA� S�?޼'?��/����>:����ҕ;2TB>��������Ν=�3����B=�\]=M�g�;.��	��+�?5�>2>�>�=?�H[�<
>�і1���7����a4>���>�T�>���>gl�9�G.�5 �^�ɾOF��?�ӽQC<>Zk?J]P? b[?���u5�,����7��Kڼ$�ξ�W>�7>�Yu>$����T��!1�Q3B��"{���h���g�����=�\6?��>��>���?IM?�|$��Ӿ��m�fb�g-=��>��c?�_�>��>B�N��R$�q��>�l?)�>6��>������!�'|���н���>'ȭ>�>�>0p>K�,���\��z�����kN9�7��=i?h?�C���f`��>L�Q?B��:�Z<���>!�v�`�!����=(�`0>M9?���=�8<>�ž4��@b{�:̊���.?=�?i�Ҿ��,��>��?/*?���>ۀ?A�>ը��Y�P���?hrS?wD?��;?���>JH1>N�ɽ+�V�^SA�K5 >�_z>9�S>?��=���=g�$�)A���"!�)�!>ٗ�=�A����(�=���=u�<���"%>^nۿKK�D�پ]�1"�@9
�Q舾A���c��٭�B\�����]Xx�Ł���&��V��?c�����2�l���?,;�?�m��R%������Z������3��>��q�l@�z諾+��z9���ྑ̬�+k!� �O��i�{�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >^C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾y1�<��?7�-?��>Ŏr�1�ɿc���y¤<���?0�@�>?H1$�ע�?,>���>�
?N|Y>�y���V�����a�>��?���?� �=k�A�m<\�^?P�;D�B��y�;�v�=��(=�+j=w�佳Ry>��>ʻA�+�#���潛�">o�m>��{�L'�X�b�2)o<�ip>y� �����2Մ? {\��f���/��T��BU>��T?�*�>c:�=��,?7H�h}Ͽ	�\��*a?�0�?��?3�(?�ڿ��ؚ>o�ܾi�M?yD6?���>�d&���t�z��=6ἱ���c�㾭&V����=ѫ�>��>=�,����\�O��L�����=W����Ϳ���F�%�}@�F'=9���B~Ͻf�����<�1n��Ω��r��:T�=P��=nXj>ŕ_>@�C>E�\>]hS?5�f?���>�#<>0���P���|���l�;�4���K˽�]�g�����о����V���^�y%��	�E���i=��9�=A6R������ �j�b�u�F���.?�$>��ʾv�M��Z,<�eʾ=���E���Ͼ��%̾!�1�%n��˟?T�A?N�o�V�Z��\���F��3�W?d`�������\��=�N����=�*�>���=���)3�.qS�i/?՝?4���*.��!p1>=����T=�%-?gB�>Wl�<"ח>&�"?T?)�o0����f>�B>u��>��>�L�=���5����p ?�QW?�罦s��Y��>�ۻ�i؊����<�e>����ڼ��G>��I<(����7Y�p�ͽN~�<&W?���>��)�4���M��Q��j�==αx?K�?� �>ik?��B?�p�<�X����S�R�Q�w=d�W?�i?�>�u��)о�[����5?5�e?B�N>��h���(�.��U��?	�n?�X?a_���l}��������d6?��v?�r^�vs�������V�m=�>\�>���>��9��k�>*�>?#��G��຿�BY4�Þ?}�@~��?��;<��$��=�;?q\�>��O��>ƾ{������w�q=�"�>����Gev�����Q,�k�8?ޠ�?���>-���������=%����?�b�?,w���&j<���<k��� ��9�<��=O��,:�����7���Ǿ8z�M���4��·>�W@�v~�>E7�ּ��yϿ����L%Ӿ�lo���?[Ȫ>DνZ+���6l�7x�Z1H��sH��9���֕>��s>���t����d���:����!��>��F=m>��B�9qᾋ�q��6=�T�>Ŗ�>�(�>�$����?�1��RW��ΐ����ϑ\?d�?���?wI?�<
>W���rQ�΀����T?�_v?�DT?(G��,��5�<%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�P�_?�a�H�p���-�K�ƽ�ۡ>��0�ge\�M������Xe����@y����?;^�?_�?���� #�@6%?&�>x����8Ǿ��<���>�(�>4*N>dH_�V�u>����:��i	>���?�~�?Jj?镏������U>�}?�$�>U�?Il�=Mb�>�h�=�ﰾ��,�jn#>��= �>��?��M?K�>Y�=��8��/�ZF��GR��$���C��>�a?e�L?�Lb>���2�K!�8�ͽ;i1��7�S@���,�v�߽$5>��=>�>��D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?[��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�e��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B�}�1=8M�>Μk?�s?�Qo���j�B>��?"������L��f?�
@u@a�^?*����+����H&��}⾊�ʼ��>YW�=F콊+�<������=����>3��>ڀ>���>kV">���=|8>g#|�&�#� ���?m���ڂ�Z���&*���>���%�tW���ܾ־���b����F�;c���$H����>jI?�2E?��n?�?�ۼ�P3>Y�޾�჻l�)���<��>��0?�D?�W ?��=�T���g��8��������>�"Q>�x�>S��>,h�>p�]���,>�+>�w>�@	>k��=���Wx��@�0>П�>�6�>
�>]<>�7>�������2h��Ww���ɽa�?93����I��4���ݍ�l����=�=�G.?��>�����Ͽ-����(H?����w,�D�*�u�>��0?F�W?b>������L��>>9��l�`J>d���k�ƽ)��JP>T�?tnk>(H>0�0�x�7��GJ�����ﺁ>d�:?�g��6���w��gC�׾��^> A�>�o<{��g���R����R�?,=��>?<�?�5���9��SQ\��,���K,>�S>;��<w
>� 7>Z����Ľ�U6��{�<iΣ=�i>��?6>��`=��>=֐���B��(�> �P>�>��:?4�?�l¼܌��T�{��b���}>�#�>8��>*�>czB�$ǫ=kE�>��y>$����Xk�rl��2L��tQ>hi�E�]���k�Wҝ=7���"R�=j�=����F1���=��~?2��	䈿v��`��|lD?+?L�=2�F<܃"�L ��zF��)�?�@ m�?1�	���V��?�@�?�	��I��=�~�>J׫>ξӑL�X�?��Ž�Ȣ���	�Y%#��R�?��?��/��ɋ��l�8>�]%? �ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?.�#�39�?�}?�@�n5��]��'<ɿ�:��̷�>賽>�*�>] �>���Ŏ������hЃ�̘^�z�>M�=��>�p�La���`�>5^b=��@���х�>S�Ҽȅ�^�>�>�4>�P�>���=<`�=�Ef�n ���K?UL�?jg��m�Ͱ�<tr�=#�Z�c!?4?7Z���Ѿ���>��[?���?�Z?Օ�><c��͚�j���c;���]<KQ>k�>��>{�x���L>�`վ:.I�橈>^��>o@/�;Bھ�4����Իۅ�> & ?SX�>s�=�� ?��#?>�j>L(�>oaE��9��x�E�f��>���>I?*�~?��?�Թ��Z3�����桿��[��:N>��x?V?�ʕ>Y���胝�UhE��AI�h���F��?�tg?�S��?>2�?��??)�A?$)f>����ؾ���L�>�H"?�i���0�.$��n�p8?��?� ?Eؒ�e�A�]��7��"���?O�`?P|(?�A˾*�8��tƾ��<؜���x<�f$<�ӱ���=�ic>T��=밻:�Kc=-7>Jm�-��Y��=��^>��>P��=�����>1=,?��G��ۃ���=��r�9xD���>�IL>����^?Ql=��{�����x��	U� �?���?Zk�?P��<�h��$=?�?U	?o"�>�J���}޾3���Pw�~x��w�j�>���>ʢl���F���י���F��T�Ž������>���>�#?�r ?y_O>� �>�I��<'�{������X^��,��b8���.�:������p�#��.�����V�{��y�>4	�����>��
?�1h>��{>E�>h��i�>� R>��>sU�>��W>Z:5>!>��<�2ѽ��O?pj��µ'�Y�ʾ쒤��]??�+c?�H�>H9��������@� ?���?C��?0�>��a�/$��?�G ?&cs�?͉�=������򖤾fe��,�ƅ�� j>vn��~�6��9B��R���
?�`?:� ;��ҾzνF�˛�<G�?���>�)k�d$q�Xk��˴>��y���2P>d:L>�
w��_W��l��욜����uZ����#����>�}'?���?�Ǿ�뾠վs׏�!�y�0��=y��>�q�>�չ>v��>u̼�̱H�w�|���4��2�<�;K?���>�G?�9?Z�P?�L?Z?�>���>d�����>,�p;$y�>x��>v}9?*-?�/?�j?V�*?�b\>���i���_�ؾ�? �?�/?߅?8�?�Ą��ϽL��J ��du�Wg��{=�"�<F�ӽ�L�]�M=O�O>�?�G�I^9�ur��q>'�6?��>��>����hf���s�<��>��
?�>�����p��l
��R�>��?��"�=��/>`��=�����"���=ʱq��ʇ=}��+7���)<��=׳�=�5�;��׺���:�������<u�>/�?x��>�C�>o@��� �C���f�=�Y>�S>i>Fپ�}���$��X�g��]y>�w�?�z�?��f=��=��=M}���U�����Z������<�?TJ#?"XT?Z��?F�=?\j#?��>+�UM���^��l����?h!,?#��>����ʾ�񨿱�3�؝?�[?7<a�����;)���¾�Խ��>~[/��.~����+D����t��8���+��?�?�A���6�ix�ſ��U\��'�C?�!�>�Y�>�>V�)�T�g�,%�1;>��>GR?�%�>G�O?4{?��[?JzT>�8�c*���͙�CH4���!>�@?���?l�?y?on�>��>/�)�j�)e��X��O"�������V=k Z>���>'(�>��>��=>Ƚ�[����>�/k�=�b>K��>㚥>��>v�w>�ۮ<H?�:�>��Ǿ'���ܛ�Qy����ږt?��?m�&?S=a���?��;�r�>�1�?h�?-?H�L�TE�=M�Լ�E���O��x�>k��>"M�>�x==�f=��,>�q�>�I�>-l�����c3���J�?8^D?�r�=\�ſ��q���p�����|e<璾*�d��{���;[�{`�=����u��������[�����tn��N嵾����ߴ{���>�i�=N�=���=�;�<#,ɼ�=�<n�I=M׎<�V=�bp��l<_a8�|�λ��$a�=jZ<�zJ= ���o}˾M�}?�5I?=�+?9�C?��y>�C>q]3���>Ě��>9?�-V>�?P����7�;�a���v��=�ؾg�׾��c��̟�{@>%oI�Y�>1U3>BG�=ߓ�<H�=��r=���=�QQ�]=�*�=B<�=K�=��=#�>�J>>6w?����K����4Q��S��:?�:�>΂�=pƾ�@?O�>>~1������a��-?s��?�S�?B�?�wi��c�>��+ᎽFi�=�Ŝ��<2>L��=��2�b��>t�J>��EJ�������3�?��@/�??gዿ#�Ͽ[k/>��C>O��=]�M�j(���C��!N���D��["?�:�ɾ$�m>�n�=�6־���<=Z:H>Ѝ=�=(�4'_�v$�=jt����!=DF�=x�>�^[>�L�=]CڽzZ�=/C=�#�=��S>_sX<��K�Fwg�]=���=�&k>(
>�A�>ǈ?�2)?Cze?���>�X�\þyɶ���>{��= �>�VW=@>�ɺ>m�5?��@?
.L?�x�>���=y�>P�>!1��o��tپ>˪�QH�<���?>��?S�>
�<�ZW�r���X<��ȽG?�k+?�?E��>�U����Y&���.������F.�]+=�mr�{RU�����m�Y�㽏�=�p�>���>
�>�Sy>��9>��N>�>�>�;�<�p�=����vµ<�������=A���C"�<}uż'��ܰ&�f�+�����ۍ;̗�;)�]<O��;d��=���>$<>��>���=���_E/>1���h�L�+ÿ=�I���*B�u4d�DH~�L/�HR6��B>�6X>����3����?_�Y>�r?>S��?�Au?$�>�#��վ�Q��e@e��PS��͸=X�>� =��y;�)Y`���M��|Ҿ���>{�>*�>BKl>�,�*5?�1�u=-��P5�:&�>1T���-�D�FGq��F������Ri������D??;����=~?��I?c�?��>gw����ؾVk0>NE���=��O�p��ۓ���?'?M��>��C�D��%;*l���ù>�L��P�	��E^1���E�����.�>@7���ξ�3��}���I���B���w�{��>=9P?;��?�`�����qO�r�t���>?�qf?o�>M�?�n?�����~�6耾W�=��n?h��?]{�?�>��K>!���rm�>F�? E�?�O�?�f?�@��x��>4��B=~<�*(�a3>��9>m��=7�><�?�8?Z�>:������O���&�4Te�֏4=��>~��>�K�>M4y>��=�O��n|����7>�R�>ag�>�k�=h�>bS�>%F��:&���??���=�}�>?�$?��>u��=��Q�"H7=�M��3�Zj���j���H��pO=1�l<'$s=��t��/�>����oy�?��c>Է��?�˾���<Z�=i=4>�j��>v� >�˃>y��>���> ��=�T>�X>�FӾo>����d!��,C�Z�R���Ѿ�}z>�����	&����w��NBI��n��tg��j�L.��V<=��ʽ<,H�?�����k��)�����R�?�[�>�6?�ڌ����֯>���>�Ǎ>�J��e���Wȍ�hᾢ�?A��?�Fc>"�> �W?X�?�1�u3��mZ���u��$A��e�ط`�F���e����
���q�_?��x?zA?穒<�<z>ۡ�?\�%��ۏ�1�>e/�u$;�<A<=x7�>�$����`���Ӿ��þ�>��;F>o?� �?`?�HV��HV��e$>>�8?52?�Cs?�2?݀;?��
��H"?<,>\�?�h?��5?�.?e/
?��4>�Y�=�����
=�b��qω��"սz�нzY����I=��=p�����#<+}#=�٢<W��^��X�;� ����<�M=���=f��=�֦>U�]?��>���>��7?���G8�e���R/?o:=^���w�n������>T�j?��?�=Z?/�c>�A�f(C��<>2r�>��&>�p\>
R�>s��J�E���=�]>V�>�ԥ=`�M�nˁ�T�	��?���J�<^�>Y��>2w>𿅽��,>W����l��r>���m����;��EK��"�Q}�����>-G?�� ?{�=c��u�Y�j�?f%8?<U?��~?�A�=Ѿfd<�WWM���B�#�>�	{=xz���w��࣠��D1�|�=+gE>�����Ԡ��kb>1��X޾�n�8J����k�L=X����U=����վ�!�S��=)&
>������ �f���ת��)J?h�j=;n��lU�gq���>�ʘ>�׮>Y:�ɜv��@�����GZ�=C��>=�:>,������qG�7���>g�L?pF?���?��D;��|3�A�������/�p?l�>��?ߑN>ƪH>��þa���|�Xo���>�9�>�5���>1��g��v9�n
���c�>��?)G->�t�>5N?��?�p?�D?��?��>���;T���c�)?A;�?.��=L�<1Ч��\e��}&�*�?l�N?3�;�VA�)�0?&��>�a,?3�C?ջ?j��=����tO����>�W�>�UG�]����z�;)�-?ӫ�>?(�?��?���=�4��Ko���������ٙ;|f�?,�a?��O?[0D?�W?�g�-���0�>A�`?Oq�?t�t?@ut> +>��>�.0?s�K<�v�>^~?�4 ?<�@?�{?/� ?�ģ>���<�H�-���|E;��;�;�ϼ���o��<ҍ=�9�Y�-� �0=�A=�=�9=��ҽ���<G�>��<Rl�>5t>Y����0>�ƺ��큾�2I>�ts�)'��Ά��'�9��=�Ӄ>DE?6�>y���>�=	{�>d$�>����#?f?��?�ꣻ)8\��Ծ��F��Ϋ>Q�@?s��=�Tl�ov��Q�u��GI=��l?8a_?]�E�Ni��W�b?��]?Ra�=���þO�b�Ï��O?/�
?R�G���>W�~?��q?Ү�>f��;n����Db�-�j�fζ=Pt�>&W���d� ?�>��7?�Q�>&�b>�#�= t۾�w�.v��v?��?� �?-��?%-*>!�n��3����������?���>~>���&?O���߾?���%����˧���������d��������1ॾ̬#<�/4>��?�~?
ZY?ir?�J�b@o�ArW�ׅ��CG��f����D`�{�6�@IH������ ��$�W���e�<�����B\�!.�?�(?λ/����>���z@���Ͼ��>�eu��0��@M�<�A��W%�=^B =��z�[2e�Ȟ��$$?�7�>Q��>�&A?c��n.�T?-���@��徨�c>���>�|b>�K�>�%���_���齔a�����ƽR͚>}gi?H�?x�h?k헼چ=������&�O���ᾳ��=��>��>�ƾ_�7��k6�B�M����u�K�����y羅�=� 5?��h>���=��?]�!?��=���)��o��w�;�%ɻҗ$?�M�?��>��->�~_�L�"����>��l?��>88�>y��o�!�	-�AA���>_��>���>��>��)�*O_�r䏿ك��;�9�`
�=Icc?�V����[�^g�>��P?�\�;Y�;@z�>7mK���"�����!,��;	>ʀ?���=`7I>iþ�{
��y�����bY.?:&?	!���.@��D�>ο/?H�?�4?7mn?ƙ<>��־	n>=V?:<?�+?'�F?�1�>�=H�>z����J��0�׼윩>b�>�c=�>�ʶ�����f��=j�.>��
�c%����=��=�6r�j{	�?����v=��ۿ%�K�jܾ��N�����
���!���<���m�9������BY{�����mV��ja��.���h��N�?�=�?tO������+/�������6��9��>�Qn��~h�]�����S�����૾?� ���N�mf��e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�{A?��(�����T=g��>!�	?�)@>��0��<��߰�/B�>�0�?e�?DbN=�W�R�0qe?�#<��F����u�=���=��=s���oJ>L�>'����A�a�۽�5>�{�>F�#�m;��&^�oj�<'k]>��ս����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=v6�ꉤ�{���&V�}��=[��>c�>��,������O��I��U��=}��n�ſ]�%��!�4a�<�}
�?�M�S�潡E���9�yȠ�0|�������=�b�=h�P>�߆>�`>=^>(�U?��f?d�>[>�.ѽ3��Ҽξ��E������H�o��]������쾣Dݾ�?��B�"����ƾ�;B�%_=UMT��V����%��yc��%C��-.?�*%>inξ[�N����޵;�{���s��M��]UȾ(.��h�>�?!1@?����tZ���Ύ;�^���?MW?2������������=���{k�<{"�>UQ�=�߾\�+��Q�(0?�z?U%�©��=�>Hh��O~>�m-?	�>�r=ǽ�>P}?�/�<F�K<.Ps>��u> h�>X��>,�T>�5����X�8
?�l]?ؒ뽐�u�b��>ڒܾ�����=$[>
���	(�T�t>��=���"�
<|�<B$��t9W?���>�)�.4���x�2�ּ�=��?�#?f6�=A3:?�]??�>���QB���;�>�AZ?��m?�&�=_ӭ��ᨾ@���I?hK�?�Z�>�(���p�I �7f��?HY�?/�?�ߴ�v����+������G?��v?s^�ws�����H�V�h=�>�[�>���>��9��k�>�>?�#��G������yY4�%Þ?��@���?i�;<��R��=�;?j\�>�O��>ƾ�z������C�q=�"�>���~ev����R,�d�8?ݠ�?���>���������=D�پ�y�?�0�?>�۾}�i�<���^u��`	�� �=K��=�鏾�Ce�d��j�E��K���0��೾G��=j|�>k�@B�~�/?:f|��͘ӿ�s��>߾�Iﾐz
?v�>���*���9������yOY��k�XYξN�>��>~�������D�{�$r;�C%����>*�v�>�S�z%��������5<��>
��>��>-��v轾ř?�b���?οv�����&�X?h�?+o�?�q?0�9<��v�3�{����-G?�s?	Z?�c%��:]��7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?*�a�M�p���-�y�ƽ�ۡ>��0��e\�N�����Xe����@y����?M^�?i�?ѵ�� #�g6%?�>c����8Ǿ��<���>�(�>*N>rH_���u>����:�i	>���?�~�?Pj?���� ����U>�}?�*�>=�?���=G��>���= ����3���">R[�=�nE���?[�M?~)�>[��=r7��/��dF�G�R����B�C�o �>��a?�WL?�b>�v��	T,�� ���̽��0����*?�=�'�r?ܽ��5>x�=>��>��C���Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�e��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?VQo���i�B>��?"������L��f?�
@u@a�^?*�ӿOۓ��g־�'���G�;�M<�+>��s�ǃ�=�2�Xä�R�-�5a�=�
�>��>][>߀W>��=z>a��u������Rů�F����K=����-����m������΅о�l7���ͼU7(�.[�+ü���~���=],V?^@J?��s?�?pu���>Ad��ߊ���I����=Y��>��/?ZF?�.?�?=�b��t�l��L���U����s�M�>��F>��>Q�>	[�>�f�:�0U>\I>�~>K�>�(�=z;=/�0=73Q>�C�>��>U�>sC<>��>Fϴ��1��n�h��
w�j̽0�?}���S�J��1���9��צ���h�=Ib.?|>���?пc����2H?#���y)��+���>x�0?�cW?%�>��>�T�/:>6����j�-`>�+ �|l���)��%Q>tl?��f>�u>z�3�d8�|�P�!~��yh|>&36?�붾EH9�%�u��H��bݾcGM> ƾ>:,D�'l��������ui�:�{=�w:?��?6���㰾G�u��B��[OR>�;\>�\=�l�=�ZM>�Tc�y�ƽH�vp.=���=�^>��?f�+>x��=�O�>�8��hF�)�>S�F>�>1�??��%?�&��!����}��N'�_�|>��>�W�>oJ>+J����=�G�>�d>�i�𢁽�{�H?�f+X>�{��[���t���\='t���Q�=㧗=���u�6���=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?���>�}?h�j?cc�>e���(���ſ�ӟ���9=ֺd>NU����w>�՟�N���|��e���v��0T�&����4�=G��>�M��H�����>�GL=_����p�h��>,��>��X<��>��?Y��>�,�>5d/>^�7>�tB��*����K?���?���0n�$��<���=��^��&?C4?�[���Ͼ ը>��\?Y��?�[?�e�>���]<��j俿K}���3�<�K>�7�>�E�>�,���GK>��Ծ�DD��q�>�՗>a����Aھ�"������=�>�c!??��>��=c3?{~!?�%~>��>��H�B��.�I����>���>uh?c��?��?�ʾg;�)���H��F�`��=>�t?�?��>(֎�Բ��3�̼K2-��O��-I�?ܵd?���;?�{�?D�B?��@?��`>��Q�ھ�୽!p>T�!?Z�f�A��%&������?�r?���>�0����ӽpǼw��Q���+?��[?�?&?��qw`�g¾ؔ�<��<��y-���#<�&O�I�>�*>���N��=��>�'�=ūn�Z�7��i<�˽=���>0N�={5�M���0=,?��G�~ۃ���=��r�?xD���>�IL>����^?jl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྾Pw�~x��w�[�>���>�l���K���ڙ���F��^�ŽZ�D�>r��>�?C~ ?��O>!R�>�3���1'��x񾏯�̻^�f�%h8�_�.�����Ѡ��0#�ݵ�y<¾��{�1K�>ZR����>��
?A'h>�{>�>³Ȼ|L�>qR>ۄ>�l�>��W>_%5>A�>Ο<%�н GR?������'����5J��_0B?bmd?�A�>dj��t������k?���?<l�?	Ov>>Hh�[+�gd?Q�>h���;
?�/:=����<�-��ؗ�t����ǰ�>9Mֽ�5:�?M�f��i
?5?_N��v>̾}ؽ2���OUJ=܋?mk>?�=���e�o��R�[���a���Ľ?��O*����T��2�������ړ��m��*I,��/�<�1?x̕?Nh�Fn־����_a�a�S�❈> �>��7>���>[a�>�����4���Z�b�`ߗ����>��H?���>=G?:�6?ţM?r�M?V��>Fq�>����.��>�#�;�>P��>��9?��.?�0?5??ԙ*?i�e>{�7���Nپ��?G�? @?nl?z�?5��X8ҽ�r��,�D�{�6��WY^=m��<ٲȽ/�X��s=��F>��?�&�o�8������n>W�7?39�>ϲ�>�Ǐ�\�����<܊�>r�?Hُ>N6����p�_�.��>|q�?�����<��*>���=6�j��\�8���=ĝܼ�ǋ=�YH��6��\ <��="0�=���R�w%�:lI;��<u�>4�?���>�C�>�@��)� �]��"f�=�Y>HS>~>�Eپ�}���$��s�g��]y>�w�?�z�?��f=��=��=}���U�����O���k��<�?@J#?%XT?_��?|�=?[j#?׵>	+�hM���^�������?w!,?
��>�����ʾ��ԉ3�؝?e[?�<a����;)�ߐ¾��Խα>�[/�h/~����>D�U���[��4��?쿝?5A�S�6��x�ٿ���[��{�C?"�>Y�>��>U�)�{�g�p%��1;>���>fR?LQ�>��O?��y?�\?��V>[f9�Tɭ�:q��~���>>�??��?�s�?�~w?E��>&�>-��%㾴���}��3(�z���Z=�Y>׋�>��>���>���=��ƽ\ŭ�|�:�p��=�ag>!'�>@i�>۪�>��x>��<��H?.l?�����c��7��pɠ��Q-��D�?�ߜ?��
?м�k ��y5�3������>���?�g�?�C/?�j,����=,���ľ�/���8�>���>�(�>�>�Ŕ�l �=�F�>a��>��=�i�Lt=�ira�;?\�O?ob>��ϿL�p�#�ľ������[�Ӿ?�� ��<�ٽ��m=��ǾԆ��
۾|�@^�[Ƃ� b�����5�)��>I��=3]>Y�T<_8�<S���>�M9=��M=�_>�F!���=ǭ��Sƍ���<�=��=rYI>�Y¼Ή˾�}?�;I?�+?��C?޸y>�:>��3�s��>ڈ���@?�V>R�P�Έ��e�;�\���� ���ؾ�x׾��c��ɟ��H>�_I���>�73>I�=MK�<z�=Ss=FÎ="�Q�=�%�=&P�=�g�=G��=��>U>�6w?V�������4Q��Z罦�:?�8�>�{�=��ƾr@?��>>�2������vb��-?���?�T�?>�?@ti��d�>K���㎽�q�=_����=2>@��=�2�W��>��J>���K��L����4�?��@��??�ዿ͢Ͽ8a/>�8>G>��R�]1���[���a�L�Y�E�!?
f;���˾���>��=*�޾ ƾe1=)�6>��c=����\�zE�=��|�HH>=�[o=��>��C>���=�����N�=c�I=r��=�SO>a먻��7�R�*���3=��=�Jc>B6%>v��>!?~30?�hd?��>8�n���ξ_����Ë>}�=Ű>�Z�=B>��>��7?�oD?��K?�ʱ>'߅=&�>�'�>�E,���m��3�I���7�<���?��?t��>9�5<� A�����)>�q�ƽ��?u�1?�?�w�>����)��<]?���O����zF��v�=fg��B>s,�>)����?��	��f�>߯�>m��>���>���>֮�>S��>H�M=�A>V߈>�;�>�4�=�S�8զ�'�ɽ�b�<���`H_9)�=K��;�����$=�#k=~X½��=���=��>z<>ܬ�>G��=����C/>߸���L����=�G��e,B��4d��I~�N/��V6�{�B>&;X>�}��A4����?[�Y>�l?>���?YAu?5�>� ���վ�Q���Ce�9VS�Q˸==�>��<��z;��Z`�}�M�b|Ҿ6��>�>�*�>�l>�%,�� ?���u=�4��^5���>����VR�8��:q�8H��(���s,i��7��}D?�:��r�=�
~?�I?�ُ?��>u�����ؾ M0>�(��C=!�7�p�r�����?��&?��>7�B�D��J̾����ܷ>�EI��O���ʯ0�g��h̷����>������о�$3�=g��I�����B� Lr�7��>�O?�?!9b�{W���UO�����,���q?�|g?i�>_K?C@?�$��tz�s��lv�=b�n?G��?>=�?>��=�������>�?Օ�?�ő?l�s?��7����>/�;�&>�ʒ�B��=Sz>џ=ɰ�=?Z�
?��
?����)�	��C��@^�-��<)�=��>�Q�>�q>#��=ݴI=�#�=ezZ>]��>��>6dh>�>�|�>B޾BU8��0?P/N�̮�>i�!?��+>[�]=	q7�	�>瑝���R��L����J���;�VP<[�=V�O>�}#>�o?}!п�R�?|=>H
��V$?��~��<N0>o �>��D=���>����o=�ƻ>ί>���^\�>���=IӾZ|>����e!��-C���R�ǽѾ*~z>	����&�I���{��DI��m���f�%j��-���;=��׽<�G�?������k���)�����Y�?�\�>�6?�ٌ�a����>Z��>|ƍ>K�����ȍ�ngᾺ�?���?�;c>��>G�W?�?ђ1�)3� vZ�)�u�p(A�*e�S�`��፿�����
����.�_?�x?2yA?�R�<*:z>Q��?��%�Yӏ��)�>�/�%';�@<=v+�>*��1�`���Ӿ��þ�7��HF>��o?<%�?vY?ETV�.��:v�>MN/?�8?��x?/@?�??�.��>�?B��=?4?�1?��E?��-?m�?,W~>��	>��r�ߦ>Ny� 4��>�&��E��ڝ�����=���=����F��?ij=:�=� I=�2��p�����:=Y� =�c�=c�y=�Ѧ>�]?�'�>�`�>��7?����V8��q���(/?n�8=
����ӊ��n����6�>��j?���?�[Z?��d>,�A��!C�E>�c�>�&>�M\>�q�>X'��E��y�=(<>t+>�=��L�����I�	�ߎ���=�<>���>W6|>�,��-�'>"��їy���d>�Q�2��Y�S�ǏG�8�1���u�m��>��K?|�?�ܙ=�)����3f�n�(?�j<?kM?a�?�$�= �۾e�9�S�J������>�ޥ<*	�e������b�:�W��:!`t>�~���Ԡ��kb>1��X޾�n�8J����k�L=X����U=����վ�!�S��=)&
>������ �f���ת��)J?h�j=;n��lU�gq���>�ʘ>�׮>Y:�ɜv��@�����GZ�=C��>=�:>,������qG�7���>g�L?pF?���?��D;��|3�A�������/�p?l�>��?ߑN>ƪH>��þa���|�Xo���>�9�>�5���>1��g��v9�n
���c�>��?)G->�t�>5N?��?�p?�D?��?��>���;T���c�)?A;�?.��=L�<1Ч��\e��}&�*�?l�N?3�;�VA�)�0?&��>�a,?3�C?ջ?j��=����tO����>�W�>�UG�]����z�;)�-?ӫ�>?(�?��?���=�4��Ko���������ٙ;|f�?,�a?��O?[0D?�W?�g�-���0�>A�`?Oq�?t�t?@ut> +>��>�.0?s�K<�v�>^~?�4 ?<�@?�{?/� ?�ģ>���<�H�-���|E;��;�;�ϼ���o��<ҍ=�9�Y�-� �0=�A=�=�9=��ҽ���<G�>��<Rl�>5t>Y����0>�ƺ��큾�2I>�ts�)'��Ά��'�9��=�Ӄ>DE?6�>y���>�=	{�>d$�>����#?f?��?�ꣻ)8\��Ծ��F��Ϋ>Q�@?s��=�Tl�ov��Q�u��GI=��l?8a_?]�E�Ni��W�b?��]?Ra�=���þO�b�Ï��O?/�
?R�G���>W�~?��q?Ү�>f��;n����Db�-�j�fζ=Pt�>&W���d� ?�>��7?�Q�>&�b>�#�= t۾�w�.v��v?��?� �?-��?%-*>!�n��3����������?���>~>���&?O���߾?���%����˧���������d��������1ॾ̬#<�/4>��?�~?
ZY?ir?�J�b@o�ArW�ׅ��CG��f����D`�{�6�@IH������ ��$�W���e�<�����B\�!.�?�(?λ/����>���z@���Ͼ��>�eu��0��@M�<�A��W%�=^B =��z�[2e�Ȟ��$$?�7�>Q��>�&A?c��n.�T?-���@��徨�c>���>�|b>�K�>�%���_���齔a�����ƽR͚>}gi?H�?x�h?k헼چ=������&�O���ᾳ��=��>��>�ƾ_�7��k6�B�M����u�K�����y羅�=� 5?��h>���=��?]�!?��=���)��o��w�;�%ɻҗ$?�M�?��>��->�~_�L�"����>��l?��>88�>y��o�!�	-�AA���>_��>���>��>��)�*O_�r䏿ك��;�9�`
�=Icc?�V����[�^g�>��P?�\�;Y�;@z�>7mK���"�����!,��;	>ʀ?���=`7I>iþ�{
��y�����bY.?:&?	!���.@��D�>ο/?H�?�4?7mn?ƙ<>��־	n>=V?:<?�+?'�F?�1�>�=H�>z����J��0�׼윩>b�>�c=�>�ʶ�����f��=j�.>��
�c%����=��=�6r�j{	�?����v=��ۿ%�K�jܾ��N�����
���!���<���m�9������BY{�����mV��ja��.���h��N�?�=�?tO������+/�������6��9��>�Qn��~h�]�����S�����૾?� ���N�mf��e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�{A?��(�����T=g��>!�	?�)@>��0��<��߰�/B�>�0�?e�?DbN=�W�R�0qe?�#<��F����u�=���=��=s���oJ>L�>'����A�a�۽�5>�{�>F�#�m;��&^�oj�<'k]>��ս����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=v6�ꉤ�{���&V�}��=[��>c�>��,������O��I��U��=}��n�ſ]�%��!�4a�<�}
�?�M�S�潡E���9�yȠ�0|�������=�b�=h�P>�߆>�`>=^>(�U?��f?d�>[>�.ѽ3��Ҽξ��E������H�o��]������쾣Dݾ�?��B�"����ƾ�;B�%_=UMT��V����%��yc��%C��-.?�*%>inξ[�N����޵;�{���s��M��]UȾ(.��h�>�?!1@?����tZ���Ύ;�^���?MW?2������������=���{k�<{"�>UQ�=�߾\�+��Q�(0?�z?U%�©��=�>Hh��O~>�m-?	�>�r=ǽ�>P}?�/�<F�K<.Ps>��u> h�>X��>,�T>�5����X�8
?�l]?ؒ뽐�u�b��>ڒܾ�����=$[>
���	(�T�t>��=���"�
<|�<B$��t9W?���>�)�.4���x�2�ּ�=��?�#?f6�=A3:?�]??�>���QB���;�>�AZ?��m?�&�=_ӭ��ᨾ@���I?hK�?�Z�>�(���p�I �7f��?HY�?/�?�ߴ�v����+������G?��v?s^�ws�����H�V�h=�>�[�>���>��9��k�>�>?�#��G������yY4�%Þ?��@���?i�;<��R��=�;?j\�>�O��>ƾ�z������C�q=�"�>���~ev����R,�d�8?ݠ�?���>���������=D�پ�y�?�0�?>�۾}�i�<���^u��`	�� �=K��=�鏾�Ce�d��j�E��K���0��೾G��=j|�>k�@B�~�/?:f|��͘ӿ�s��>߾�Iﾐz
?v�>���*���9������yOY��k�XYξN�>��>~�������D�{�$r;�C%����>*�v�>�S�z%��������5<��>
��>��>-��v轾ř?�b���?οv�����&�X?h�?+o�?�q?0�9<��v�3�{����-G?�s?	Z?�c%��:]��7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?*�a�M�p���-�y�ƽ�ۡ>��0��e\�N�����Xe����@y����?M^�?i�?ѵ�� #�g6%?�>c����8Ǿ��<���>�(�>*N>rH_���u>����:�i	>���?�~�?Pj?���� ����U>�}?�*�>=�?���=G��>���= ����3���">R[�=�nE���?[�M?~)�>[��=r7��/��dF�G�R����B�C�o �>��a?�WL?�b>�v��	T,�� ���̽��0����*?�=�'�r?ܽ��5>x�=>��>��C���Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�e��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?VQo���i�B>��?"������L��f?�
@u@a�^?*�ӿOۓ��g־�'���G�;�M<�+>��s�ǃ�=�2�Xä�R�-�5a�=�
�>��>][>߀W>��=z>a��u������Rů�F����K=����-����m������΅о�l7���ͼU7(�.[�+ü���~���=],V?^@J?��s?�?pu���>Ad��ߊ���I����=Y��>��/?ZF?�.?�?=�b��t�l��L���U����s�M�>��F>��>Q�>	[�>�f�:�0U>\I>�~>K�>�(�=z;=/�0=73Q>�C�>��>U�>sC<>��>Fϴ��1��n�h��
w�j̽0�?}���S�J��1���9��צ���h�=Ib.?|>���?пc����2H?#���y)��+���>x�0?�cW?%�>��>�T�/:>6����j�-`>�+ �|l���)��%Q>tl?��f>�u>z�3�d8�|�P�!~��yh|>&36?�붾EH9�%�u��H��bݾcGM> ƾ>:,D�'l��������ui�:�{=�w:?��?6���㰾G�u��B��[OR>�;\>�\=�l�=�ZM>�Tc�y�ƽH�vp.=���=�^>��?f�+>x��=�O�>�8��hF�)�>S�F>�>1�??��%?�&��!����}��N'�_�|>��>�W�>oJ>+J����=�G�>�d>�i�𢁽�{�H?�f+X>�{��[���t���\='t���Q�=㧗=���u�6���=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?���>�}?h�j?cc�>e���(���ſ�ӟ���9=ֺd>NU����w>�՟�N���|��e���v��0T�&����4�=G��>�M��H�����>�GL=_����p�h��>,��>��X<��>��?Y��>�,�>5d/>^�7>�tB��*����K?���?���0n�$��<���=��^��&?C4?�[���Ͼ ը>��\?Y��?�[?�e�>���]<��j俿K}���3�<�K>�7�>�E�>�,���GK>��Ծ�DD��q�>�՗>a����Aھ�"������=�>�c!??��>��=c3?{~!?�%~>��>��H�B��.�I����>���>uh?c��?��?�ʾg;�)���H��F�`��=>�t?�?��>(֎�Բ��3�̼K2-��O��-I�?ܵd?���;?�{�?D�B?��@?��`>��Q�ھ�୽!p>T�!?Z�f�A��%&������?�r?���>�0����ӽpǼw��Q���+?��[?�?&?��qw`�g¾ؔ�<��<��y-���#<�&O�I�>�*>���N��=��>�'�=ūn�Z�7��i<�˽=���>0N�={5�M���0=,?��G�~ۃ���=��r�?xD���>�IL>����^?jl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྾Pw�~x��w�[�>���>�l���K���ڙ���F��^�ŽZ�D�>r��>�?C~ ?��O>!R�>�3���1'��x񾏯�̻^�f�%h8�_�.�����Ѡ��0#�ݵ�y<¾��{�1K�>ZR����>��
?A'h>�{>�>³Ȼ|L�>qR>ۄ>�l�>��W>_%5>A�>Ο<%�н GR?������'����5J��_0B?bmd?�A�>dj��t������k?���?<l�?	Ov>>Hh�[+�gd?Q�>h���;
?�/:=����<�-��ؗ�t����ǰ�>9Mֽ�5:�?M�f��i
?5?_N��v>̾}ؽ2���OUJ=܋?mk>?�=���e�o��R�[���a���Ľ?��O*����T��2�������ړ��m��*I,��/�<�1?x̕?Nh�Fn־����_a�a�S�❈> �>��7>���>[a�>�����4���Z�b�`ߗ����>��H?���>=G?:�6?ţM?r�M?V��>Fq�>����.��>�#�;�>P��>��9?��.?�0?5??ԙ*?i�e>{�7���Nپ��?G�? @?nl?z�?5��X8ҽ�r��,�D�{�6��WY^=m��<ٲȽ/�X��s=��F>��?�&�o�8������n>W�7?39�>ϲ�>�Ǐ�\�����<܊�>r�?Hُ>N6����p�_�.��>|q�?�����<��*>���=6�j��\�8���=ĝܼ�ǋ=�YH��6��\ <��="0�=���R�w%�:lI;��<u�>4�?���>�C�>�@��)� �]��"f�=�Y>HS>~>�Eپ�}���$��s�g��]y>�w�?�z�?��f=��=��=}���U�����O���k��<�?@J#?%XT?_��?|�=?[j#?׵>	+�hM���^�������?w!,?
��>�����ʾ��ԉ3�؝?e[?�<a����;)�ߐ¾��Խα>�[/�h/~����>D�U���[��4��?쿝?5A�S�6��x�ٿ���[��{�C?"�>Y�>��>U�)�{�g�p%��1;>���>fR?LQ�>��O?��y?�\?��V>[f9�Tɭ�:q��~���>>�??��?�s�?�~w?E��>&�>-��%㾴���}��3(�z���Z=�Y>׋�>��>���>���=��ƽ\ŭ�|�:�p��=�ag>!'�>@i�>۪�>��x>��<��H?.l?�����c��7��pɠ��Q-��D�?�ߜ?��
?м�k ��y5�3������>���?�g�?�C/?�j,����=,���ľ�/���8�>���>�(�>�>�Ŕ�l �=�F�>a��>��=�i�Lt=�ira�;?\�O?ob>��ϿL�p�#�ľ������[�Ӿ?�� ��<�ٽ��m=��ǾԆ��
۾|�@^�[Ƃ� b�����5�)��>I��=3]>Y�T<_8�<S���>�M9=��M=�_>�F!���=ǭ��Sƍ���<�=��=rYI>�Y¼Ή˾�}?�;I?�+?��C?޸y>�:>��3�s��>ڈ���@?�V>R�P�Έ��e�;�\���� ���ؾ�x׾��c��ɟ��H>�_I���>�73>I�=MK�<z�=Ss=FÎ="�Q�=�%�=&P�=�g�=G��=��>U>�6w?V�������4Q��Z罦�:?�8�>�{�=��ƾr@?��>>�2������vb��-?���?�T�?>�?@ti��d�>K���㎽�q�=_����=2>@��=�2�W��>��J>���K��L����4�?��@��??�ዿ͢Ͽ8a/>�8>G>��R�]1���[���a�L�Y�E�!?
f;���˾���>��=*�޾ ƾe1=)�6>��c=����\�zE�=��|�HH>=�[o=��>��C>���=�����N�=c�I=r��=�SO>a먻��7�R�*���3=��=�Jc>B6%>v��>!?~30?�hd?��>8�n���ξ_����Ë>}�=Ű>�Z�=B>��>��7?�oD?��K?�ʱ>'߅=&�>�'�>�E,���m��3�I���7�<���?��?t��>9�5<� A�����)>�q�ƽ��?u�1?�?�w�>����)��<]?���O����zF��v�=fg��B>s,�>)����?��	��f�>߯�>m��>���>���>֮�>S��>H�M=�A>V߈>�;�>�4�=�S�8զ�'�ɽ�b�<���`H_9)�=K��;�����$=�#k=~X½��=���=��>z<>ܬ�>G��=����C/>߸���L����=�G��e,B��4d��I~�N/��V6�{�B>&;X>�}��A4����?[�Y>�l?>���?YAu?5�>� ���վ�Q���Ce�9VS�Q˸==�>��<��z;��Z`�}�M�b|Ҿ6��>�>�*�>�l>�%,�� ?���u=�4��^5���>����VR�8��:q�8H��(���s,i��7��}D?�:��r�=�
~?�I?�ُ?��>u�����ؾ M0>�(��C=!�7�p�r�����?��&?��>7�B�D��J̾����ܷ>�EI��O���ʯ0�g��h̷����>������о�$3�=g��I�����B� Lr�7��>�O?�?!9b�{W���UO�����,���q?�|g?i�>_K?C@?�$��tz�s��lv�=b�n?G��?>=�?>��=�������>�?Օ�?�ő?l�s?��7����>/�;�&>�ʒ�B��=Sz>џ=ɰ�=?Z�
?��
?����)�	��C��@^�-��<)�=��>�Q�>�q>#��=ݴI=�#�=ezZ>]��>��>6dh>�>�|�>B޾BU8��0?P/N�̮�>i�!?��+>[�]=	q7�	�>瑝���R��L����J���;�VP<[�=V�O>�}#>�o?}!п�R�?|=>H
��V$?��~��<N0>o �>��D=���>����o=�ƻ>ί>���^\�>���=IӾZ|>����e!��-C���R�ǽѾ*~z>	����&�I���{��DI��m���f�%j��-���;=��׽<�G�?������k���)�����Y�?�\�>�6?�ٌ�a����>Z��>|ƍ>K�����ȍ�ngᾺ�?���?�;c>��>G�W?�?ђ1�)3� vZ�)�u�p(A�*e�S�`��፿�����
����.�_?�x?2yA?�R�<*:z>Q��?��%�Yӏ��)�>�/�%';�@<=v+�>*��1�`���Ӿ��þ�7��HF>��o?<%�?vY?ETV�.��:v�>MN/?�8?��x?/@?�??�.��>�?B��=?4?�1?��E?��-?m�?,W~>��	>��r�ߦ>Ny� 4��>�&��E��ڝ�����=���=����F��?ij=:�=� I=�2��p�����:=Y� =�c�=c�y=�Ѧ>�]?�'�>�`�>��7?����V8��q���(/?n�8=
����ӊ��n����6�>��j?���?�[Z?��d>,�A��!C�E>�c�>�&>�M\>�q�>X'��E��y�=(<>t+>�=��L�����I�	�ߎ���=�<>���>W6|>�,��-�'>"��їy���d>�Q�2��Y�S�ǏG�8�1���u�m��>��K?|�?�ܙ=�)����3f�n�(?�j<?kM?a�?�$�= �۾e�9�S�J������>�ޥ<*	�e������b�:�W��:!`t>�~��ߑ�v4�>�����	�Vwc��)<�M&��^�����$^�=���n��VeA��A>��=�����,������Ʈ���B?9��=%�ž��v��7���K4>v�>*�>|p\�h�����E������ž=��>گ|>Üϻ[��z7�5����t>��J?��`?��a?�=��H<o�}�;�U$���ؾ˽=�d%?�R�>���>�E>$#���������3X���J����>
�?�a!�fo`�����	��S�3��-�=�!8? �u>v��>�o$?�]?`�e?e�;?�?��>>��=�Ǿʕ%?�
�?��=�W���T��=7���G�q��>)�(?7���>D9?ZS?z�(?	�N?H?�?>-� ��_B�`�>~��>\7Y����2wc>'�J?@�>ӋV?؈�?9B>"v6�,o��蕠����=�(>�<2?��!?U�?}ʶ>�F�>f���Ϋ>$j�>:�\?I(r?�j?il�>h�>��u�pk?��d����>�0�>QN6?��v?<�j?l&?���>���<���|p����ҽ��H<�Қ=N��<`۞;�t�<h�'���� k����
�\jz������#�48==��=G\�>�t>����31>��ľ�e����@>�ϣ�h`��������:�o
�=Tz�>W�?܀�>�#� ђ=���>%J�>����#(?R�?�?�z;��b��ھ��K�?�>I�A?���=��l�Vx���u�g=��m?Ҏ^?��W�]E��1nN?z�m?��¾�Hc�Q����N�!f&��!�>
~�>�H����>^?.�k?��?�V���^�2x���r^�gyѾ2 >�k�>�#;�C����>FbG?n]�>q��=t�W>W[���y����Ǿ�o?��?O�?g҈?��=c�E�ֿ̬�����K_?��>ԡ��X�&?�8��̾f腾�S�����#������r@��������U·�f�(z�=B�?��k?��v?�J^?@I�'c��a����opY�d��O���B�� @�5�A���s���6��l��V�:==ԃ���m�M�?�% ?7؍� �?����VؾF��PF;>�(��4B�%=��+=Kx9<�� >�Q��Dg�E��jB4?�5�>N7?\�7?ݶu�g�I�K�O���E��;$�✃>n��>�ǆ>���>�ۼ�ƾ��-�֘Ӿ�Ͼ\���A>ʧw?@K$?C�A?���=�a�# �����@[�=�/�4�u�J�>�g�>s!���	"=����m��9�����0���_�<=I>T�h?-W>	x=)C�?�/@?G��4�W�C����j��x��&>g�3?�=��I>コ�����>��l?ry�>ʩ�>�����"��y�w�ǽ�j�>��>P�>+�o>y�.���]��������5�6�ݵ�=}h?�����a�N��>�7R?��:d <~�>~���^!�qR��eI.���>� ?4��=d�3>�%ľl.	���}����(?Ƣ?�ؔ���1��P�>".#?%��>DW�>�I�?ь�>��ľ��S�
�?߀b?r�F?�=?��>��=O޽�uŽt>'�0�+==L�>��`>(�x=7��=��5�U��"���&=�@�=8{��½?m<n��Ҕ<���<�=>;mۿ�BK��پ�
���&?
�C爾����c������a������Wx�6��F�&�TV�97c�����#�l����?~=�?����60�����甀������>2�q�?������ ��;)�����G����c!���O�t&i�V�e�~(?
�����ǿ���,oݾtv?"5?��y?B���!���8�b'>��<NZ����ך�Q�οpҙ���_? ��>/��Υ�.�>���>�K\>ˍs>�����蝾}��<ʄ?�f,?���>H8q�'Pɿ����>�<���?A@�A?
'�r�V2>=e�>�?O9>�*4�j!������>.��? �?�O=p�V�����c?^�E;J�F����.��=��=��3=]���hB>���>����-@�����~2>�T�>I}�R����Y�'��<��Z>&G���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=��l�ƿ�#��+�0.�<��tZ���0����d��f��sr�2I�v�w=�E�=��S>���>��U>�X>�W?�k?tѾ>�6>�I�a/���;� �����n���a��p��nB��q�C�ݾ���O�5���3ʾ֜<���=�Q����� ��ob��G�c.?`�%>�˾��M��$v<��Ⱦ�>���󀼪l��;'2�N�m�:f�?rlA?�����[U�A|�����軽�MX?_��
��M�����=�����<2�>��=��⾔�3���R�zf0?oj?F���.��C*>�&�ɾ=��+?rq?�L\<��>�E%?G�*��n�I�[>��3>hģ>	��>�> ���}۽7�?فT?�������̀�>��z�A~a=�Z>�-5�2���[>i,�<Ǧ���4Q�`��F�<B[?�k�>��1����Z�����;(FI=v�y?$�?d��>�n?Q�9?< V:�&����T�y��[k�=��^?5�j?��=�����ɾ�P���;?v�X?�gK>�-\� �{�'�7� ���?�'p?D/?�p��g~�t ���z��_3?��?��B��w���i	���߾�/?F��>e#?����@�>L�T?~-��������^�@�q\t?� @�D�?�S>�̥��<>@��>՛�>�H�=�|�ᣗ�ƺ+�0;�����>+n��	g��LG�]�= ?m�W?y�
?��g�0>����=��ӾT��?Nb�?N6�^#��`�/��^w���1�I�>p��>��=�6w<7�s��mP��D���4�����}��i�>��@��3�O�>�I�s�������:��P4�ҳH?�S�>6�P�����y�������0�9H/�H	���K�>4�>a��������{�m;�r������>o:���>>�S� #�������7<&Ւ>֟�>]��>�V��5���2��?�M���>ο����0���X?te�?vg�?Au?�l;<cw���{�����.G?f�s?KZ?ĭ%��]�q8�c�j?����a�_73���C�YRL>T33?�a�>uw-�ǂ=�>���>��	>-A/��Ŀ�𶿸u�����?�i�?C���-�>���?(-?����Q���s��О+������=?�$>^j���` ��=�I���+,	?��-?�V�A'�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?$�>��?D�=�]�>>��=}��M�.�fb#>��=��?�x�?��M?�N�>'	�=��8�w/��ZF��IR�$���C��	�>��a?D�L?�Fb>�d��	
2��� ��|ͽ�1��D�^@��,�|�߽+5>��=>�>�E�Ӿ�K]?N�
�*Pۿ ㆿ�h1�tp#?�>�� ?�ҕ=�_3�fC����T?DC����>�U赿�蚿a�H�߮?�� @F��>����9<4�L
>�w�=e�>��C>{DL��쾪[D>A�>?#�����v�D�u��>�?n�@�u�?p�[��?�y�U���#�y�~t�Q?�v�=Ÿ4?�K־{͋>��>c��=�σ��ӫ�K�t�PT�>�l�?��?˺ ?��`?8Td��=��-/=��>�h?
?j��<����;>=�?��	�	#��(b��z`?�@}@��X?�5��d�ٿS�������UO���g�=��="#>�\�MC=�g'>(n�}3�X�k�ojk>u�>%ђ>RZ+>��>��9>�ۂ�����1��S퍿r�B���	�E����,�h��\u�}$��w�þ�zվ�ս�&g�w񧽿�J��
��}x�J�=J.V?,6R?��o?G�>���("+>� ���8�<�����=�V�>ew0?��H?-�*?��=����?a���U]��k݇��&�>g'I>�U�>�q�>D��>;���
\>�?H>B}�>Um�=y=�_�<SM=�[>;��>4�>F'�>�?<>v�>̴�*.��Ėh��w�(1̽R �?����J��3���A������Za�=�a.?�t>U��_?п����{0H?8 ���(�+�+�.�>��0?6eW?^�>����T�5>u��նj�R>�9 �:�l�ي)�S6Q>�k?��f>��u>�k3��(8�&�P�۰��{>46?z඾-b9���u�c�H�^Uݾ�
M>!о>ŬG�Պ�������?i��Dy=�P:?�}?��������
�t�����~�Q>��\>��=�ϩ=�SL>�4e�&�ǽ��H�B[/=$Y�=��^>��?�n2>�:�=e��>f]����R�æ�>jB>��$>�??$?�Y������	��D'�P�x>K��>�ʀ>X�=i1I�}p�=��>l�a>��洀��o��SH�
c>k#_���X�TFz���=ؙ�V]>��=�r��\�/��*=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿp�?6D�����7���t���ͽ#�,>�1O?�b����F=	:|�ݫ[?��>�r�P����пLˁ����>�D�?V�?o�^��)����?����>�$�?�K?��^>��R������e>&�!?�4?W�>0�6�˸D���>���?�g�?$�H>ӓ�?�Js?g��>��|�@//�����{��rc{={��;ｑ>52>�_���D��ߓ��?���	k������\>)=���>���}����=Ę��FZ��B�m����>`"r>bUE>��> ?��>>s=b����*����� a,?S�?oh�;P���>c#f>���FD��-?d��>Aa뾐p>@�a?���?�?�F[>!TC�}��ʓ��]���jn���>څ?���>!�9���=7�T<	ߝ��ν�z�=�`�>�T�S�M>aU�>(~�>���=�4�>�J$?P?+6&>Ds�>8L��!���fI�>�>3��>�F?��j?�)*?-E���z<�#���g���z�^���;>{q?p�.?\Xu>e������]�ý�쭺Yj��2ir?��|?{����?u�?:?O�9?*��=]|U�e�Ӿ�����Ϩ>��!?|h�ĵA��{&�)��a�?E&?(T�>�В�SԽ��׼ ��#>��v?�\?�,&?����a�/9þ�1�<�3#���Z�{��;L�@���>��>����Y��=��>h�=�m��J6�!:f<���=�>�5�=!7�[鍽�iA?bz�=c��������R��N!�;�>���>���5�h?��ջR�{������뒿h(��d�E?iP�?�?#�="�j�66]?��n?��%?G�?�1�Cz����?���3Ym�j55�]�C>��>KkH=�¾�W���|Ŀ����D���_�p��?[�>y/?8�>�+���?��<��y���/�n�����h��XJ�#�@�0la�֦��3���t�-�7��>�l���>C��>b��>�]y>9H>��2>J�>��;>�@�>/�?��?��>(�;�Р=�ҽ�iJR?_����'����«���0B?qid?D(�>�h�9���>����?���?�q�?%<v>�zh��.+�Ah?�8�>����n
?3e:=FX�Lg�<�a��,��{�����떎>vN׽I:�)M�G�f��l
?0?�G���̾�׽l;��a�=��?^�%?d,���V�{�w�|\�]�U�"f��0�����,��eid�ଐ�v���K'����+�k��<-l)?���?Ru��O�$�����b�~<E�r�E>��>D��>N�>��I>�1�S�+�v�X��G(�Y㈾)S�>v�p?��i>�<?��D?f�V?�43?1	�=k��>hK���Į>�W�=#��>B��>2Ra?�?�=?�p?vf@?,}�>�7�y���o����>b?��,?o��>q��>������<.��B;Ž-�2>�h�>��<fH��N>��.�>�X?���Ӭ8������k>��7?��>|��>���-���<�>�
?�F�>+ ��}r��b�W�>���?;��}�=��)>���=N�����Һ8Z�='�����=�7���y;�Tc<���=��=�Ht������9�:���;{p�<'w�>��?���>`A�>\A���� �v���p�=�Y>�S>�>{Gپ�}���$��|�g��Xy>x�?({�?0�f=��=V��=g|���S����+���?��<Y�?�H#?�WT?[��?�=?j#?۹>@*�}M��F_����Q�?�#,?qő>��m�ʾ�ب��3���?�Y?1a����+6)�Wd¾uHս b>�\/��7~�:�����C�(kk����T.��3��?$˝?�w?�S�6��[�����(r���EC?L��>���>��>l�)���g���ֺ:>U��>i�Q?��>0P?�
{?�,[?�KT>�r8���ԙ��W1�
�">��??@��?��?��x?�a�>�>�%*���߾���w�X���jW={^Z>�h�>x��>�v�>{"�=g�ǽ=�����>�oѧ=S�b>���>D��>4�>�w>jβ<�G?��>�d�����*����l�<�E�u?��?.�+?&{=R����E��K��OD�>Fm�?���?=7*?��S����=��ּT߶�Z�q��*�>�ܹ>�/�>ѓ=�iF=�_>O�>f��>I��]��n8�q3M���?XF?ݞ�=۶ſ?p��ae�J����S�<�W��bM�l5���V�p��=�����-�����"�9�����ۃ��==���Қ�ĵ��-j?$�X=�7>��=����/���Lu<�=��=7S<_���h:�<WL5���l<�u��|H<6�;��V=6j���˾ԏ}?�;I?�+?��C?�y>�;>k�3�B��>�����@?+V>��P�҈���;��C ���ؾx׾��c�%ʟ��H>5`I�A�>�83>�F�=AL�<��=s=�=zR�/==$�=�O�=�g�=��=�>HU>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=J����=2>r��=w�2�T��>��J>���K��B����4�?��@��??�ዿТϿ6a/>]�7>H9>��R�Ɓ1���\�S�b��[Z��!?�L;��D̾�0�>���=�(߾��ƾ��.=��6>�^b=zo��U\���=I�z�<=�l=�Љ>�C>�I�=�=��<4�=;J=E��=/�O>p��R7��+�h4=���=W�b>�&>��><�?�e0?Td?�%�>�#n���ξ��B�>%F�=2�>|��=�nB>�g�>M�7?խD?��K?�u�>"�=j��>o��>>�,�Y�m�:c�ߵ���m�<Y|�?׆?k�>��U<�A��r��5>���ý?EK1?2�?WԞ>�7��h��<���+��<�A=@1�:x��=��B0S��S�����d��y�.����>�&?X�>�,]>�R�:q�u<���>[-:>J<e�>b��=z�={��=b2"<�{=���=S& �aY�<S�=���=ʠ�%�@�I���������rs�=���>�>w��>{P�=ꟺ�H�5>����3�L����=�Ҩ�g�?��c�l-~�7�/�:F�+l?>l�_>��I�7���A?�;k>�O>�m�?<�o?�k!>��)ؾ�����w�wG�c�=q��=�>�]k:���_��R��4Ҿ���>���>r��=9��>w��?c[�B�>�����_B�~0z>�-۾��=GV�Vǁ�_�������@�j��<�R[?�އ��I=�%�?�:l?�
�?@\�>�y����5�=���uem���澔'!��u��Ӥ�>e?m�?�R�[oR��/̾��ŷ>�I��O��ƕ�=�0��������t��>c����о 3��i��s�����B��{r���>E�O?��?�Hb��]��0WO�����;���f?Jig?�:�>nT?�J?B��/a�/���U�=�n?֫�?�=�?DT>1Ǻ=���R�>T
?~��?�@�?�8s?Ԇ4����>�`��Б>�����=�!>�=���=]�?dx	?�	?� ���?	��������_�=F=è�=�a�>ѕ�>vCq>���=O@z=w��= 4R>��>Ƶ�>�`>���>s �>��پ�3 ��a?n�>��k>��:?=I�>��d=�੼C����ڽz*��+�RN�=�E���=��[����<�ѿ��?�5̿b�?�L>��6��p%?�d���&;�y>$��=�H@�B?�~�=[��>[6>���>�K==&^;>,$>2H��yP>�f���>���!��K��� ���>�(�����c9�'�P���^�1���|�辕Ip�"�����B�5����?�Er��B��o�-����؎�>�m>�?�i��j�$>>e$@?"b�>'�������Ӗ�j�����?H��?�:c>a!�>7�W?A�?K�1��"3��iZ���u��(A�~ e��`��ލ������
��濽S�_?]�x?�tA?���<�3z>��?��%�\͏��#�>�/�:+;�"�;=�>�>�����`�e�ӾS�þ��)kF>�o?w#�?A`?~PV��B����b0?P*?%ap?�2?:iB?��=��
?=J�;�?x=�>jo;?��?e�"?�
�>]fw>f�=��(=i蕽3���W3��!��>H=�h�=;?ɼ\=�B���Q�G(0=U������d7н��k_�=&0==<��<0�<��>�]?�W�>䯆>Z�7?���@_8������/?':=̣�����������>�j?���?^\Z?U/d>��A��C��>�P�>'v&>�\>T@�>����XE���=�d>E>;m�=�L�M���I�	��_���I�<%>���>�K|>J���Q�'>1j���Tz�X}d>��Q�Uɺ�� T�c�G���1��v�EM�>��K?
�?$I�=t�$W��1Bf��#)?}X<?�MM?��?	��=��۾��9���J�	/���>ь�<| 	������!����:�J��:.�s>x+�������>� ���%�x'9��V�ծ��F��w �e�G>��Ͼ8"侭�#��8�>�|�=ُ������タ������<?|��=��s[y�|y�����=�>�>P��<N���E�W���<�I�>N�S>��w=i]ž�<�����&w2>KD?��Z?�)]?�q��p��c�C�$��9��Era=��?2��>`�?m�7>1�0=%���y�!�a���J��T�>�x?�??�l�l�t�+���{�������=p3?e�q>`9?M"?�\�>�/J?��?G�>��>���="����+?�l�?��= 4�GP0���(��R���>5�?"�޽]��>�?�?��(?�%E?3�?ķ�=_��D�_T�>��>�~^������y>7�Q?ݑ�>�I?N��?��P>>+�Cd��DV���:%>��>ϵ!?�
?:?�?�>�e�>c1ξ��P>3��>e�Q?,�n?��q?���=2??�L�=�?��=�l>�w?��)?ߍc?|y?R�.?Y%�>4� =d��b/ҽ��%�Q����:%�q��Ӱw=����$*���<e�4=�p�<�&D��,0��qC��ݗ<�c/�f�ȼ�]�>�du>�x��d'/>��þp���ѨA>���?P���슾�<�?��=���>�k?�ה>�L$�¸�=^��>�s�>�����'??u>?�aB;5�b�0ھ��I��o�>�A?���=�Dl�>��\�u�SPi=-�m?�b^?�gZ�
��H�b?{�]?�f��=�(�þ�b����y�O?��
?��G���><�~?��q?���>��e�9n�~���Ab���j��Զ=;r�>MX��d�@�>��7?�O�>��b>�-�=�u۾��w��p���?��?�?G��?j,*>G�n�)3࿄���R���^?$��>`D����"?�1��Ͼ�X���펾�⾠������ $��:L���u$��΃��׽	��=x�?�s?�[q?��_?� ���c��<^�<���vV����!�j�E�k�D�ytC��n�Se�f��C"���G=�,־��r�x?�?�5-?,Nm����>Z��˭�A 龙��>!�ȾAuG�!n
>���;�U*>'�><�F� ����þ��:?� �>��>�?ze��>�D]���6�����>"�T>CX�>��&?���=U���:�b�-�RP��Z����9X>��c?kC*?j5?>S���iJ�|ۀ���侭�Ӽ[ ̾B��=��r>��n>�>W��p<	o��̙&��-v�=���p����*�v��=�Uh?��>�>��?#PL?	��?�������@�[F��/?>�N\?��>���>O@�I��[�>sl?�\�>�\�>Z����3"�5ys�Aռ�D&�>�ϧ>���>�kq>�'&�Q]�����M��Z�8���>Yk?"뇾S`^�u�>;�Q?��;6X<T��>����N� �M���	@/�� > k	?mۆ=��0>ؾ�A��"�E&��� ?�U?�Ϗ�M?�tW�>�)#?��>P�k>��~?���>����ST���?�mg?@?�y8?���>�=���)���'��6=x��>��O>�����=�'���8�D&F��6��	>)�S��I�J�;=X�<^Y<΍��om7>�dۿHBK���پ�����09
�����y?��au��c�uk��c1��spx�2��)[&�		V��$c�O�����l���?L0�?���H<��g���@���������>XVq�]y}��߫���pߕ����/ܬ��Y!��O�~i��e��<?�S����Ŀ靛�I���1?Ő?�Cx?Ն��\��}d!�.��>�+�� Ue��D��S����ͿЧ�I�r?{��>��� X����>f�"=��>B��>@����?���"�c?i]
?�ִ>,��Y.�������T=+�?f��?�^A?E�(�K��]U=���>)W	?/�@>6[1�jG�r�����>��?��?$�G=
�W�\"��Me?���;#�F�+'커?�=��=A�=��iJ>��>��<�@��ݽ��3>g��>�� �(�\-_�4ӽ<4_>bnؽ{��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=����ƿ�m�&K�!F;=$g< \���׽De��3y�����^�pA�O�r=��	>�o|>��>E�5>��H>��Y?ׅ_?r��>�%>%��:��yؾ�.3�:�p�ae�������	��я��D���ᾳo��A�c6�^�ľd�7��=�M�Y듿���3�]��PJ��$$?��)>����wI����<*0þ��򜭻A!��/%ξ!�.�Zp�v<�?Xu8?�����E����])��ˣ��d?����h
�!����>��%:^��n�>��=��ܾI7���F�ڐ0?��?�Ⱦ^m���;>�_��K�=Dg*?�|�>n<��>�Z$?�$����d�F>ڍ>�-�>�)�>Z�.>�賾_hҽ� ?��T?��"���v�>^��cQ��2��<3��=�4���S��a7>b�a<�����ź��b�8<��i?�>ݑ=���+��|�y��=�@����{?
u(?��>֐V?�Z?B8q�����d�5P��s��a�N?��|?g�=>)�1X��񆾴�?��m?~>�>I�u����	7-�*��k?4?:�3?bL!���y�$�����W��TC?��v?s^�xs�����S�V�h=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�$Þ?��@���?��;< �Y��=�;?k\�>��O��>ƾ�z������!�q=�"�>���~ev����R,�f�8?ݠ�?���>�������p�<_��7�?�P�?��Ѿڿ޽Y]"���h�˭&����=v,�=w�=O��=W��.*�w�����_Ͼ/����e�>Ђ@����ة>�潍�ٿE�ϿҢ��	�̾ ˠ�ҧ,?�6�>��;�!����Yj���c�e�D��=��ܖ��΢>u�>�哽����~4{�&!;��{��3,�>��
�'"�>}dR���q���01<ق�>�>��>�ү��T�����?�����8ο-Ğ�\.���X?#�?I�?��?ȵO<<Eu�TS{�����G?3�r?1pY?ܨ%��[�S�5��v?�PM�__���J'�[N:���>�
=?^��>I$�"�<9��=�[�>�E~:�&�貲�����!f��v�?5=�?Q� ��:	?�s�?�?�׽�E���qx�{���)[��?�,�A"z�����05�]�>��B? $?��W3�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?���>��?�%�=��>Ӯ�=i%��f��y$>ƚ�=l�C��?:KM?;��>F��=��:�(n/�=F��P�����C��l�>�0b?ЕL?�xb>v ��);*��� �kϽ�@6�X����@�á��&�f�2>'�?><>�.L�y�Ӿ:8.?ǂ��	׿�������R�B?���>�?������\����<ݣX?��+>�}�1���a��m�9���?���?	?R^ܾ�섽Y@$>��[>��>�ԏ�I�nT����>��??NmA�(v���a�D��>QT�?{� @J�?�b��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?rQo���i�B>��?"������L��f?�
@u@a�^?*��ٿ�����F��[F�����=^4�=5�M>P�ĽX��=꼓./=<�|=��=ج�>�&�>�н>+�>+c>��>�8���X� �������|/��	����鋅����v�I�����XD�����2�o����<�{�)�I�!�����=!�K?�Q?�Hu?��?��*��~c>& �{�P=�u�v��<�FL>��9?�C?��9?rB>OB�L_\�|�x�K��Sw�}2�>��K>;�>��>�Ģ>�L�;1�H>p9W>`��>d<>�ē=��y=��*>���>�*�>tG�>�x�>�A<>��>�ʹ��0����h��w�8$̽� �?�����J�81���7��l����c�=�b.?�|>���d>п����Z0H?z ��(�u�+�}�>��0?eW?��>���p�T��3>���[�j��X>�' ��l��)�	!Q>Sl?d�`>�n>b�1���5�M�8 ����|>��7?���f>=�6�u�>iL���侌G>:1�>�����2h��'~��g��!n=�Q9?P�?0���������p�;����J>9Si>:�=�=6@K>F끽�ʽ+I���=l��=�%_>�W?�,>p��=���>���9�P��˩>0�B>%�+>M�??��$?������������.��fv>V�>�9�>��>H�J�#�=|��>Hb>i��넽oO���?��W>"-��_��t�o�z=����=&-�=n2 ���=�w�$=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ(�>��jp���φ���t���K=�b�>x�H?*7��@�m�9��?�� ?^�ᗤ�O�ǿ�yw�R�>� �?�,�?��m�(����&=�H	�>���?Y�Y?�a>��׾Z0\�.Ȍ>��=?0GN?�a�>����4�n�?yT�?'�?�h5>	(�?��j?td�>4��������f6����)=�8�=hѠ>�!�=β���3�����]e��a�i���	*>��V=D�>s��?ؾz��=�������[����>cGs>D�?>#�> E�>]T�>쑓>�u�<�I�}V����mkD?��?���v�y��ڃ=�="����>9�0?W�<�t˾Υ�>#U?	�?U�V?P�>E���Ė�����������H>�t?KN�>S��-gP>����9�9�<�Q>�U~>��=0۾F����0=�q�>:?#	�>p�=�=%?6
"?\�=�^>T�2��R����H�ó�>��>:�3?�X_?D�?�@���^�Ί�o��YN�je�=طf?�i5?�L�>��������չX;�:�=V�$�p;j?�u�?7[�	�?ǝ?d�6?�8?�b��RB�YW�"���y	?�g!?���xjA�Cx&���
�?��?2+�>j����[Խ��ؼ�\�y����	?"�[?��%?.m���`���þy:�<��$�
]��r�;�]A���>e�>>���os�=��>�ܭ=��l�`Q6��4S<C��=H��>�Q�=I"7�Z�>=,?��G��ۃ��=t�r�xD���>�IL>����^?pl=���{�����x��o	U�� �?۠�?ck�?�
��9�h��$=?�?C	?�"�>^K���}޾���@Qw��}x��w���>���>G�l�x�+���ř���F����Ža�	����>ъ�>w�?�	?=f�<z��>�'*�]%�rJ:��U��w��Pľ`o?���2�3�(���,=៍�g߶�$|���@�� }�>��z=�gx>N �>�=,�1>鳮>^w6>��_>�l�<�d�=�s�>�)�>��>֏�=�����¾�*S?���6T)���}-���C?u�c?"��>�X��ل��S�^[?�?�4�?�n>�i�++���?d� ?�����
?>E=�B�d��<�3���H�����~,�G��>��潘�8���J��Ag���	?��?������̾�xѽ9��3�u=x�{?��?����]�=�p�v�=�(�e��7�=�zZ�r^���q�I�h�:�|��lf���}�	�-�Z$��t2?���?�'�lh�d~��(�Y�)�X����=�"?1��>w��>���>�׾@�;�#!a�E!�ls�p�>t�n?�7>�H-?]P?�6a?��F?�TU>�>Z<P�>��:��b�>���>�Y?MP9?�pP?2?G�d?�b>~ܽ`5�>e�%?n	?}V?��?���>h���c�L�=��<��>;�P���ؽ���=��/=첺=��-=�F%>���>i;A?�0M���]������O�^�d?~�>Yo�>��ĺm‾�M>�ͭ>���>:'z>����� �֟/?��?Ѕb��5D=�S�=e�=�2�mі<<C	>�R]�ޘ8����������	��=!k�ۙ�;l���D�=�<!d��	q�>\�?w��>�>�>A?��� ����~��=�X>!ZS>��>�Uپj{��)���g�DKy>�o�?xp�?W�f=B��=���=����p�����G������<��?9]#?�VT?T��?��=?q#?�>9��B��q\�����g�?]#,?&��>���)�ʾ�䨿��3�Q�?�Y?>7a�����?)��~¾�Խ�u>*]/��1~������C�mCu�,���O����?��?�@���6��X�!���}c����C?R��>�N�>&�>��)��g�$��D;>�P�>�Q?��>5qS?H[v?>M?��]>�M0�Sͮ�Ҝ�N���A#=>�A?��{?��?lMz?^��>?}>�5��پqT �r� ��jٽ�����<��`>
�>���>��>�>�=�'Ž̡���2G����=�r>v�>�>E��>�Mz>��<��G?���>U]��Q��ꤾƃ��=�؛u?���?y�+?�P="��q�E��E���J�> o�?���?3*?ݿS�k��=�ּ�ᶾ~�q�Z#�>�׹>B2�>�ړ=�wF=�\>w�>���>�*�b�p8�IM��?�F?���=��Ŀ�-q�@kl�_����^�<�V��w�^�y�p�$i�$�=����/�������_�0��h͔�,���N������>+Ղ=���=�$�=�b�<�ʼU1�<�/=��L<��g=`Uv�Xz1<P �}��4x��Թ����<;�D\=4疻'�˾�}?�;I?��+?��C?y�y>�:>֗3�9��>�����@?V>5�P�����i�;�I���� ��.�ؾGx׾��c��ɟ�uH>bI�I�>�83>�G�=3N�<��=9s=@=�R�5=�$�=�O�=�g�=V��=��>U>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>`�,>Zx�=5O��,�eJ�q.V�f�Q�B�$?|!?���;-,x>��F=-��m<Ⱦ�f=�y)>�p=�;�3�[�w�=g���A=��m=���>.C>�[�=)Y��")�=���=a��=o�B>����+t��nC���=;��=ݱh>r�'>f�>4S?)S/?Q3`?�<�>&ml��Ѿ`,þme�>���=��>%ن=�kB>~��>�S7?6D?�$J?
�>��u=�ƺ>p��>�+��j�J�徎>����<~��?jB�?r��>��;�l9�u��?�g���7?�S0?�?�2�>���g�(��{~$��VR�&�<���=��g��L�v�|L���	޽Q+�=aQ�>V��>��>�s>��>� A>�9�>a0>j=<��T=H��8�5�`����z�=��<���<u�� ��;	��gQ����U��] <�=�<��=��/<c�=�a�>�">���>��=�&���C,>.O��d�L�n��=���D���e��|���)��7�~KG>�TH>����&p���#�>��[>�*L>�D�?�w?��9>1C��3Jݾ�֛�`�k�[qu��!`=_�>X^;��=��h[�;�I�!�о']�>y��>��O>��a>DX�g=��sI>¾j�6��$�>�d���������E#��c����՚��=X���<�R?Ou��QL�=�?��E?���?w��>�i���>XE��8�������y��d�>`�?l/?�i�Ҡ_�:̾�񾽔ѷ>c8I���O�I���3�0���׷�m��>v���0�о�"3�k������}�B��Tr�@�>`�O?B�?��a��[���]O����*@��W[?�qg?�C�>;N?�I?�u���V�w��4�=��n?��?�3�?�G>�C�=1������>lS	?}��?v��?�ts?�F?��_�>�*�;�
">����)�=[8>��=�Z�=Ѽ?V
?Sb
?qל�Q�	��p��k�E�]�=&�<�x�=10�>�A�>w�r>��=��g=�|�=��[>���>���>��e>�ţ>E�>i�ľ����Y'?��>A4�>#V-?u˂>�o=�@�����<L��1��4��Q���:���Iv=#&�<�M�<�(�!��>WSſ���?G�T>�_�&??$	�|KR��D><:�>����m��>��v>���>6G�>��>���=��~>��>�Ѿ��>��!�7�B�o�R���Ҿ��{>@՜����p)�N�����I��׷��+��7i��쁿=�}��<uR�?g*��s�l���*�%i���S?��>�H5?�R��3τ��r>�?�>̎>?E������U�����u��?���?18c>l�>��W?`�?�1�}!3��qZ�S�u�('A��e���`��፿.���Ö
� ��U�_?��x?�uA?f#�<�8z>"��?]�%��Ϗ�(�>y/��%;�$N<=R,�>�$����`��Ӿ��þ0�(_F>u�o?�"�?�W?"UV�-'��b�="K?4�=?;�^?�s?��??�aؽ�7 ?���=t�0?��?�o?��8?��!?!��>x�>"Y���o,�R�}�1@b�R���M��<�,<�܋=�Uj=>�R<.�k��B���=�P��� &�J_`�[]�DZ�=���<��=z��=f��>'�]?�:�>�_�>��7?*��Jo8�Ю�E/?ǫ9=5�������&���>��j?��?�EZ?g�c>��A��!C�'>i�>�O&>��[>kd�>�e�5{E���=�>�_>�X�=s�M�������	�zf��X��<H.>rj�>��l>����Z4>O(��Z���R>L꽧�ž<N��dH�c-9�◾��>�M?�?�\�=���b�׽w�c��{?Ȼ6?vQ?�~?�o>4e����#�T���,��>���	G#�6E���5���?D���<&��>���ߑ�v4�>�����	�Vwc��)<�M&��^�����$^�=���n��VeA��A>��=�����,������Ʈ���B?9��=%�ž��v��7���K4>v�>*�>|p\�h�����E������ž=��>گ|>Üϻ[��z7�5����t>��J?��`?��a?�=��H<o�}�;�U$���ؾ˽=�d%?�R�>���>�E>$#���������3X���J����>
�?�a!�fo`�����	��S�3��-�=�!8? �u>v��>�o$?�]?`�e?e�;?�?��>>��=�Ǿʕ%?�
�?��=�W���T��=7���G�q��>)�(?7���>D9?ZS?z�(?	�N?H?�?>-� ��_B�`�>~��>\7Y����2wc>'�J?@�>ӋV?؈�?9B>"v6�,o��蕠����=�(>�<2?��!?U�?}ʶ>�F�>f���Ϋ>$j�>:�\?I(r?�j?il�>h�>��u�pk?��d����>�0�>QN6?��v?<�j?l&?���>���<���|p����ҽ��H<�Қ=N��<`۞;�t�<h�'���� k����
�\jz������#�48==��=G\�>�t>����31>��ľ�e����@>�ϣ�h`��������:�o
�=Tz�>W�?܀�>�#� ђ=���>%J�>����#(?R�?�?�z;��b��ھ��K�?�>I�A?���=��l�Vx���u�g=��m?Ҏ^?��W�]E��1nN?z�m?��¾�Hc�Q����N�!f&��!�>
~�>�H����>^?.�k?��?�V���^�2x���r^�gyѾ2 >�k�>�#;�C����>FbG?n]�>q��=t�W>W[���y����Ǿ�o?��?O�?g҈?��=c�E�ֿ̬�����K_?��>ԡ��X�&?�8��̾f腾�S�����#������r@��������U·�f�(z�=B�?��k?��v?�J^?@I�'c��a����opY�d��O���B�� @�5�A���s���6��l��V�:==ԃ���m�M�?�% ?7؍� �?����VؾF��PF;>�(��4B�%=��+=Kx9<�� >�Q��Dg�E��jB4?�5�>N7?\�7?ݶu�g�I�K�O���E��;$�✃>n��>�ǆ>���>�ۼ�ƾ��-�֘Ӿ�Ͼ\���A>ʧw?@K$?C�A?���=�a�# �����@[�=�/�4�u�J�>�g�>s!���	"=����m��9�����0���_�<=I>T�h?-W>	x=)C�?�/@?G��4�W�C����j��x��&>g�3?�=��I>コ�����>��l?ry�>ʩ�>�����"��y�w�ǽ�j�>��>P�>+�o>y�.���]��������5�6�ݵ�=}h?�����a�N��>�7R?��:d <~�>~���^!�qR��eI.���>� ?4��=d�3>�%ľl.	���}����(?Ƣ?�ؔ���1��P�>".#?%��>DW�>�I�?ь�>��ľ��S�
�?߀b?r�F?�=?��>��=O޽�uŽt>'�0�+==L�>��`>(�x=7��=��5�U��"���&=�@�=8{��½?m<n��Ҕ<���<�=>;mۿ�BK��پ�
���&?
�C爾����c������a������Wx�6��F�&�TV�97c�����#�l����?~=�?����60�����甀������>2�q�?������ ��;)�����G����c!���O�t&i�V�e�~(?
�����ǿ���,oݾtv?"5?��y?B���!���8�b'>��<NZ����ך�Q�οpҙ���_? ��>/��Υ�.�>���>�K\>ˍs>�����蝾}��<ʄ?�f,?���>H8q�'Pɿ����>�<���?A@�A?
'�r�V2>=e�>�?O9>�*4�j!������>.��? �?�O=p�V�����c?^�E;J�F����.��=��=��3=]���hB>���>����-@�����~2>�T�>I}�R����Y�'��<��Z>&G���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=��l�ƿ�#��+�0.�<��tZ���0����d��f��sr�2I�v�w=�E�=��S>���>��U>�X>�W?�k?tѾ>�6>�I�a/���;� �����n���a��p��nB��q�C�ݾ���O�5���3ʾ֜<���=�Q����� ��ob��G�c.?`�%>�˾��M��$v<��Ⱦ�>���󀼪l��;'2�N�m�:f�?rlA?�����[U�A|�����軽�MX?_��
��M�����=�����<2�>��=��⾔�3���R�zf0?oj?F���.��C*>�&�ɾ=��+?rq?�L\<��>�E%?G�*��n�I�[>��3>hģ>	��>�> ���}۽7�?فT?�������̀�>��z�A~a=�Z>�-5�2���[>i,�<Ǧ���4Q�`��F�<B[?�k�>��1����Z�����;(FI=v�y?$�?d��>�n?Q�9?< V:�&����T�y��[k�=��^?5�j?��=�����ɾ�P���;?v�X?�gK>�-\� �{�'�7� ���?�'p?D/?�p��g~�t ���z��_3?��?��B��w���i	���߾�/?F��>e#?����@�>L�T?~-��������^�@�q\t?� @�D�?�S>�̥��<>@��>՛�>�H�=�|�ᣗ�ƺ+�0;�����>+n��	g��LG�]�= ?m�W?y�
?��g�0>����=��ӾT��?Nb�?N6�^#��`�/��^w���1�I�>p��>��=�6w<7�s��mP��D���4�����}��i�>��@��3�O�>�I�s�������:��P4�ҳH?�S�>6�P�����y�������0�9H/�H	���K�>4�>a��������{�m;�r������>o:���>>�S� #�������7<&Ւ>֟�>]��>�V��5���2��?�M���>ο����0���X?te�?vg�?Au?�l;<cw���{�����.G?f�s?KZ?ĭ%��]�q8�c�j?����a�_73���C�YRL>T33?�a�>uw-�ǂ=�>���>��	>-A/��Ŀ�𶿸u�����?�i�?C���-�>���?(-?����Q���s��О+������=?�$>^j���` ��=�I���+,	?��-?�V�A'�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?$�>��?D�=�]�>>��=}��M�.�fb#>��=��?�x�?��M?�N�>'	�=��8�w/��ZF��IR�$���C��	�>��a?D�L?�Fb>�d��	
2��� ��|ͽ�1��D�^@��,�|�߽+5>��=>�>�E�Ӿ�K]?N�
�*Pۿ ㆿ�h1�tp#?�>�� ?�ҕ=�_3�fC����T?DC����>�U赿�蚿a�H�߮?�� @F��>����9<4�L
>�w�=e�>��C>{DL��쾪[D>A�>?#�����v�D�u��>�?n�@�u�?p�[��?�y�U���#�y�~t�Q?�v�=Ÿ4?�K־{͋>��>c��=�σ��ӫ�K�t�PT�>�l�?��?˺ ?��`?8Td��=��-/=��>�h?
?j��<����;>=�?��	�	#��(b��z`?�@}@��X?�5��d�ٿS�������UO���g�=��="#>�\�MC=�g'>(n�}3�X�k�ojk>u�>%ђ>RZ+>��>��9>�ۂ�����1��S퍿r�B���	�E����,�h��\u�}$��w�þ�zվ�ս�&g�w񧽿�J��
��}x�J�=J.V?,6R?��o?G�>���("+>� ���8�<�����=�V�>ew0?��H?-�*?��=����?a���U]��k݇��&�>g'I>�U�>�q�>D��>;���
\>�?H>B}�>Um�=y=�_�<SM=�[>;��>4�>F'�>�?<>v�>̴�*.��Ėh��w�(1̽R �?����J��3���A������Za�=�a.?�t>U��_?п����{0H?8 ���(�+�+�.�>��0?6eW?^�>����T�5>u��նj�R>�9 �:�l�ي)�S6Q>�k?��f>��u>�k3��(8�&�P�۰��{>46?z඾-b9���u�c�H�^Uݾ�
M>!о>ŬG�Պ�������?i��Dy=�P:?�}?��������
�t�����~�Q>��\>��=�ϩ=�SL>�4e�&�ǽ��H�B[/=$Y�=��^>��?�n2>�:�=e��>f]����R�æ�>jB>��$>�??$?�Y������	��D'�P�x>K��>�ʀ>X�=i1I�}p�=��>l�a>��洀��o��SH�
c>k#_���X�TFz���=ؙ�V]>��=�r��\�/��*=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿp�?6D�����7���t���ͽ#�,>�1O?�b����F=	:|�ݫ[?��>�r�P����пLˁ����>�D�?V�?o�^��)����?����>�$�?�K?��^>��R������e>&�!?�4?W�>0�6�˸D���>���?�g�?$�H>ӓ�?�Js?g��>��|�@//�����{��rc{={��;ｑ>52>�_���D��ߓ��?���	k������\>)=���>���}����=Ę��FZ��B�m����>`"r>bUE>��> ?��>>s=b����*����� a,?S�?oh�;P���>c#f>���FD��-?d��>Aa뾐p>@�a?���?�?�F[>!TC�}��ʓ��]���jn���>څ?���>!�9���=7�T<	ߝ��ν�z�=�`�>�T�S�M>aU�>(~�>���=�4�>�J$?P?+6&>Ds�>8L��!���fI�>�>3��>�F?��j?�)*?-E���z<�#���g���z�^���;>{q?p�.?\Xu>e������]�ý�쭺Yj��2ir?��|?{����?u�?:?O�9?*��=]|U�e�Ӿ�����Ϩ>��!?|h�ĵA��{&�)��a�?E&?(T�>�В�SԽ��׼ ��#>��v?�\?�,&?����a�/9þ�1�<�3#���Z�{��;L�@���>��>����Y��=��>h�=�m��J6�!:f<���=�>�5�=!7�[鍽�iA?bz�=c��������R��N!�;�>���>���5�h?��ջR�{������뒿h(��d�E?iP�?�?#�="�j�66]?��n?��%?G�?�1�Cz����?���3Ym�j55�]�C>��>KkH=�¾�W���|Ŀ����D���_�p��?[�>y/?8�>�+���?��<��y���/�n�����h��XJ�#�@�0la�֦��3���t�-�7��>�l���>C��>b��>�]y>9H>��2>J�>��;>�@�>/�?��?��>(�;�Р=�ҽ�iJR?_����'����«���0B?qid?D(�>�h�9���>����?���?�q�?%<v>�zh��.+�Ah?�8�>����n
?3e:=FX�Lg�<�a��,��{�����떎>vN׽I:�)M�G�f��l
?0?�G���̾�׽l;��a�=��?^�%?d,���V�{�w�|\�]�U�"f��0�����,��eid�ଐ�v���K'����+�k��<-l)?���?Ru��O�$�����b�~<E�r�E>��>D��>N�>��I>�1�S�+�v�X��G(�Y㈾)S�>v�p?��i>�<?��D?f�V?�43?1	�=k��>hK���Į>�W�=#��>B��>2Ra?�?�=?�p?vf@?,}�>�7�y���o����>b?��,?o��>q��>������<.��B;Ž-�2>�h�>��<fH��N>��.�>�X?���Ӭ8������k>��7?��>|��>���-���<�>�
?�F�>+ ��}r��b�W�>���?;��}�=��)>���=N�����Һ8Z�='�����=�7���y;�Tc<���=��=�Ht������9�:���;{p�<'w�>��?���>`A�>\A���� �v���p�=�Y>�S>�>{Gپ�}���$��|�g��Xy>x�?({�?0�f=��=V��=g|���S����+���?��<Y�?�H#?�WT?[��?�=?j#?۹>@*�}M��F_����Q�?�#,?qő>��m�ʾ�ب��3���?�Y?1a����+6)�Wd¾uHս b>�\/��7~�:�����C�(kk����T.��3��?$˝?�w?�S�6��[�����(r���EC?L��>���>��>l�)���g���ֺ:>U��>i�Q?��>0P?�
{?�,[?�KT>�r8���ԙ��W1�
�">��??@��?��?��x?�a�>�>�%*���߾���w�X���jW={^Z>�h�>x��>�v�>{"�=g�ǽ=�����>�oѧ=S�b>���>D��>4�>�w>jβ<�G?��>�d�����*����l�<�E�u?��?.�+?&{=R����E��K��OD�>Fm�?���?=7*?��S����=��ּT߶�Z�q��*�>�ܹ>�/�>ѓ=�iF=�_>O�>f��>I��]��n8�q3M���?XF?ݞ�=۶ſ?p��ae�J����S�<�W��bM�l5���V�p��=�����-�����"�9�����ۃ��==���Қ�ĵ��-j?$�X=�7>��=����/���Lu<�=��=7S<_���h:�<WL5���l<�u��|H<6�;��V=6j���˾ԏ}?�;I?�+?��C?�y>�;>k�3�B��>�����@?+V>��P�҈���;��C ���ؾx׾��c�%ʟ��H>5`I�A�>�83>�F�=AL�<��=s=�=zR�/==$�=�O�=�g�=��=�>HU>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=J����=2>r��=w�2�T��>��J>���K��B����4�?��@��??�ዿТϿ6a/>]�7>H9>��R�Ɓ1���\�S�b��[Z��!?�L;��D̾�0�>���=�(߾��ƾ��.=��6>�^b=zo��U\���=I�z�<=�l=�Љ>�C>�I�=�=��<4�=;J=E��=/�O>p��R7��+�h4=���=W�b>�&>��><�?�e0?Td?�%�>�#n���ξ��B�>%F�=2�>|��=�nB>�g�>M�7?խD?��K?�u�>"�=j��>o��>>�,�Y�m�:c�ߵ���m�<Y|�?׆?k�>��U<�A��r��5>���ý?EK1?2�?WԞ>�7��h��<���+��<�A=@1�:x��=��B0S��S�����d��y�.����>�&?X�>�,]>�R�:q�u<���>[-:>J<e�>b��=z�={��=b2"<�{=���=S& �aY�<S�=���=ʠ�%�@�I���������rs�=���>�>w��>{P�=ꟺ�H�5>����3�L����=�Ҩ�g�?��c�l-~�7�/�:F�+l?>l�_>��I�7���A?�;k>�O>�m�?<�o?�k!>��)ؾ�����w�wG�c�=q��=�>�]k:���_��R��4Ҿ���>���>r��=9��>w��?c[�B�>�����_B�~0z>�-۾��=GV�Vǁ�_�������@�j��<�R[?�އ��I=�%�?�:l?�
�?@\�>�y����5�=���uem���澔'!��u��Ӥ�>e?m�?�R�[oR��/̾��ŷ>�I��O��ƕ�=�0��������t��>c����о 3��i��s�����B��{r���>E�O?��?�Hb��]��0WO�����;���f?Jig?�:�>nT?�J?B��/a�/���U�=�n?֫�?�=�?DT>1Ǻ=���R�>T
?~��?�@�?�8s?Ԇ4����>�`��Б>�����=�!>�=���=]�?dx	?�	?� ���?	��������_�=F=è�=�a�>ѕ�>vCq>���=O@z=w��= 4R>��>Ƶ�>�`>���>s �>��پ�3 ��a?n�>��k>��:?=I�>��d=�੼C����ڽz*��+�RN�=�E���=��[����<�ѿ��?�5̿b�?�L>��6��p%?�d���&;�y>$��=�H@�B?�~�=[��>[6>���>�K==&^;>,$>2H��yP>�f���>���!��K��� ���>�(�����c9�'�P���^�1���|�辕Ip�"�����B�5����?�Er��B��o�-����؎�>�m>�?�i��j�$>>e$@?"b�>'�������Ӗ�j�����?H��?�:c>a!�>7�W?A�?K�1��"3��iZ���u��(A�~ e��`��ލ������
��濽S�_?]�x?�tA?���<�3z>��?��%�\͏��#�>�/�:+;�"�;=�>�>�����`�e�ӾS�þ��)kF>�o?w#�?A`?~PV��B����b0?P*?%ap?�2?:iB?��=��
?=J�;�?x=�>jo;?��?e�"?�
�>]fw>f�=��(=i蕽3���W3��!��>H=�h�=;?ɼ\=�B���Q�G(0=U������d7н��k_�=&0==<��<0�<��>�]?�W�>䯆>Z�7?���@_8������/?':=̣�����������>�j?���?^\Z?U/d>��A��C��>�P�>'v&>�\>T@�>����XE���=�d>E>;m�=�L�M���I�	��_���I�<%>���>�K|>J���Q�'>1j���Tz�X}d>��Q�Uɺ�� T�c�G���1��v�EM�>��K?
�?$I�=t�$W��1Bf��#)?}X<?�MM?��?	��=��۾��9���J�	/���>ь�<| 	������!����:�J��:.�s>x+��`!Y�c�>w���@�~�N�	2�)�,U�������7>����Ñþ+��RF�>j�>"⾧hI��
���F����3?�k�=�fþI_���N�e
�=Jl�=@*�> �h=�H=�]/�3������<���>�77>���z藾�%�b����q>�8?�GR?��d?a)��e�{��"K� ��X¾�;��q?�o?�-?�[�>m�$�)����E$�ks�2zG�`7�>T?��:�kM_� v��R���;��Ⱥ=G�?�d�>���>��$?�z�>�*M?{;?��?�:+>'�!�r �g�?��?1�<�97��g���
2�'�R��T>��?�#�_l>W�#?��?��0?ȝ6?��?P�!��
��!R����>���>��e�׍���l�>�QO?�͇>�.4?��t?�8�>��,���Ծ�`��gL�=t1�>Q�?9N�>O�+?Lfr>���>`���&�P>��>24?��?�?7�)>;��>�X��� ?$��>���>��>�-?Uza?�j?�t-?���>�9=���5�����[=�hѽj��� ٽ{����>?\�=�!�=�;�=K�=b����s�=�~�;(�;��S�=H�z=�B�>8�t>��X�1>�ľ����xnB>H㡼ɞ���F���X;����=@��>ɖ?���>}�"�4z�=�K�>�
�>ݶ�3�'?��?!?ӆ;�>b��۾��L���>��A?���=�l�DX��	�u�I d=��m?�^?+�W�lD��%�b?��]?>6�M=�ľjWc�n�)�N?kw
?�H�Ԗ�>y
?s�q?7$�>�;f�K�m�����Rb�)Sl�Է=Ӝ>���me�|Z�>Ţ7?���>�a>�e�=��پ�w�HѠ�J?濌?;��?jފ?0)>�3n�T�1��V^���w]?+��>i ����#?ݼ�\^ξ����+����5���m7��i3��1(��Ή$�����k�ؽ1w�=�q?^�q?�rq?��_?�� ���c��#^����LnV����q���dD�ilD��'C�Υn��{����������~J=�%���^�]x�?a?���O�	?�����F;t�Ӿ����N�����F���=i�{����i,�=�����~n�?愾I5?A
�>Z_?�\B?<+q��yb�F�+�Y�O���%�S,X=�ۣ>���>@1.?k�>�Z���R�4�þ饮�.Q���k>}BU?l�?�O?C"�.-J����T���Ĩ5�ѐ���;o<ܛ=(��J���X���*��uI��zh��)�%%������ >��?e�>' �=U��?a?�/���ľ�K=���Z�%qؽ��i>��-?�5>�V�>����}�ܾ'��>��l?���>���>����!��|�Cw̽��>��>س�>�ar>��/��[�������}e9����=R=f?�D���]b�[��>�4T?�� �~�<���>I]Z�!�"��#���3$�a�>;?���=Jw:>��ƾ3e���z�n����(?�?�����)��k�>a
#?ۢ�>}�>�Ղ?�8�>^i��Y�;;��?�B_?�K?})A?���>֥=񵽦M��j'��=~��>O+P>�x=˹�=�c���_�:y"�i�R=|�=�^�����_[+:�ļ �~<a�=��5>�pۿZvK��iپ�P�k�/
��و��Ʊ�SM��1g�/���B��dx�VC��p!��TU�>�c�����MSl�YR�?���?�=��T��a~��kV������Oa�>��p���������������6߾�a��'�!�t�O�S�h��ae�J�'?�����ǿ��:ܾ5! ?�A ?<�y?��;�"���8�� >(D�<,����뾨����οA�����^?���>���/��i��>ȥ�>�X>�Hq>����螾�0�<��?1�-?��>Ҏr�0�ɿ`���1ä<���?-�@��@?�/(���꾅�S=���>ܻ
?h�H>f�*��2�����>�О?��?�_U=.]V�������e?�&�;�E��͊�=t�= ��=Y�"=_[�GFI>���>��!�5#<���ҽ��7>%��>4����Gta��P�<C�_>�ʽ�M��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=����M���e
�X�D�%$�g@�<�A����<����Ě����!���K W<>Bh>���>�$>���=���=(�(>~E??�)L?( >Ǵ�=��=���|ʾ���U�Ԟ�������Ϫ��N��~���BwɾT0�����¾�����=��4�={�Q��䐿P!��a��GF��G-?Q #>j%ɾ��N����;ݫɾ(���%,�;尿k�;[�0��Fm�L��?�@?����0V�,�̀���p����V?�������̭���=������.=G#�>f?�=���ϲ0�V�Q��&0?��?.%��������)>�����<t�*?�?��u<>A�>$�%?p-���]�X>��2>�j�>	q�>��>�e���޽��?�iV?������m.�>����u~�H{I=΂	>,x7��T���S>��<�F���K`�w���O/�<Q�r?��@>)=G�\1�_��U؜>�����a?,S!?�g�>[D�?P�>4Q���v$�b'J��y�HĤ>i@�?Ԉ�?��o��8�>�e�H&��|D?�� ?1��>�&�<�'���޾\`�i"?Z�l?�?��%���k�x���]�+��4??~:�?$9j����y�񾝜2����>p>I>=q�>����n�>u�?#߾����N�����;f?�G@�@^*/>��j��h=�ߪ>3z�>#^ݽD=o�ι��}��̡�ʶj>gS��la]���˾�.�H��>3�Y?٧�>�/�������=V.���H�?6�?�þ������<�g����a���/_�=D�W>n��>����W!F���Ҿ=g��=Ծ������>��@$&��R��>Gϑ�����Cȿ�|��;;���oA?q`�>�|=����d�[ht�|09�[J�`(þ�#�>�0>�B�����-�{��4;��e��
=�>��	���>~�S��x������bK<V�>>m�>h܅>.���j��0��?����6ο�������X?y<�?�?�?w4?d�N<zxv�Sg|�(D/���F?�Ms?��Y?x�&���[�~-8�ƽj?����`�+L4���D���T>��2?\��>V-��ˀ=��>�G�>-�>�Z/�g{ĿǾ������I�?؝�?x>�{�>U9�?��+?-U�����%����*�~B�ԝ@?|C->�o��^!�-=��Y��N�
?7/?����&���_?ݙa��p��-���ƽ�ݡ>��0��Z\�XY������Ve�����8y����?E^�?��??��� #�N4%?N�>u���h=Ǿ���<{�>�)�>7N>z0_���u>/
���:��c	>��?d}�?�g?���������T>��}?�(�>#�?y��=���>��=�	����:�I�">��=_�<�a?��M??�>�F�=L=9��	/�v^F��BR��B�ѸC���>��a?��L?)�a>�|��R�0��� �B=ν��1�����<@��b.�Ѕ���4>��=>��>- E�|�ҾF05?���D�Կ�܅��6��"?EV5>�G?�f���"��R�=]�W?)7:>Ѭ*��d��t���ZX��y�?���?�(	?�ݾ��<c�q<��>��>\���f��r/��7�=�YH?�RC������Y����>���?@���?�c���&?]m����5�i���	��њ���,=�.?���7؞>�� ?-�~=_�������0H_���]>' �? O�?�?1�X?��i�:��щ5�p�>B�n?�
�>?|'���Ҿ.:>v
?� �΄��]xԾ��k?�@
�@0�u?�謹�:ӿ2���}���;ݾ��K�Q�Խ�>|T���<Sd�>�� >9�>�[D>E�>
�>�>�`�=0�=m�>�%����w���	��H�a��#!�#�Tf���	�����H�,������
 '�ޠ��k�߼��b�8ē�f������=�Z?$�V?5�r?M�?h��TM$>�c��ptl<�R��ݠ=>]k>��-?e�G?�T'?ơ�=�̃��u_�J��������-���6�>�
\>]��>��>���>��<DE>�;>�Ԉ>�:>�=��=L&�=Aiw>�ۭ>�h�>�z�>]�;>6�>�Ĵ�A3���h�q�v��4̽?��?�l����J�&=��y��c���Ň�=o.?	V>|��?,пR䭿3#H?)ꔾ�>��+���>|�0?FW?��>)߰�QV�$�>�?	�nUj��>�B ��3m���)��vQ>�b?�j>��>�2�Q%<��FL����Y>-�/?������%�a0w��:B��߾/wO>���>��Y�M �f(�����]�j���\=�;?A?mj���S���i�#̌��ZC>xYF>�&=䉫=r=>t����ս�kE��)=+��=Pdj>'�?�o4>���={��>vߕ��yL��8�>�@>��&>cI??��#?/j&�����%��D�/���w>l��>S�>6� >&I��%�=<��>KQi>�)�cX��.l��;��[>(ZG�JU�>}y���=I�>l�=%��l<���=�~?���䈿���d���lD?h+?� �=-�F<��"�= ���H��D�?o�@m�?��	�ҢV�3�?�@�?�
��4��=�|�>׫>�ξ�L��?��ŽEǢ�ʔ	�)#�aS�?��?+�/�`ʋ�8l��6>�^%?�Ӿ�M�>�V �����5>k�����SF��P�>/�_?[і��A=��ƽ��?F��>��	�hB���ο��l����>g��?�-�?@�l��ٖ�kKE�w��>+��?NW;?�0>�Α�$7u���>!�=?�BD?��>[
����<���?˜�?L��?̙O>nL�?c?�˪>����__)��h�� �����4=�_=�1�>U[�=Q	Ѿ]3�@n���c��V~s�g�S>��C=���>?�O%ƾ��=o撽d}���s�<z�>qiz>��>>���>��>F7�>%��>��><P"�`u�*䘾9�??h��?8�j���=�暼���ur>b�%?6�7>����H�>-0?lfx?Q�1?��X>���*h��Vɿ����� ļ{o�>�?���>\�0w>$I����+�_/7>o��=Z��=����� �/����> �?<��>IH>L�'?bS?���=Ӄ�>�Z��^��C;���?d��>��$?��n?d_?�rξL�@�e�����'P��L@>�n�?=x<?#�D>�ϒ�k���h���k������T=�?���?Z�sj)?
��?c
<?"$?��t>+ȩ��CӾPD�=p�>֍ ?j���KLA���)��=��6?,��>�E�>d���L���ڼ���i���I�?�$Z?b' ?�
� ^���;���<��o�IT��Rû�ܯ���>��>��h��,�=��>���=Ns���8�E��<y��=`�>I�=U1�3���d/0?� �;���T�t=x4m���4�g5s>|Zh>M����"^?w8���v�Kڧ��X����l���?��?� �?�3Ҽ��k��J?��?A�?L|�>�RվPl����Ծ�s��2:n�]��� >���>a.M�&�㟿S���s��d{��ৄ���9?���>��"?�M/?�ʼ���>N�þkOM�疡����)!Q������=�l[�\~��κ씾	�D�IJ��-�D���?ؽٕ >m��>�+=7�>_�>�Y>T��>��<��p>4�?!��>��>P0>��+<G�N�>BR?�����'����֮��.B?�id?��>b�i��������?`��?aq�?n?v>Voh��*+��]?H�>��4m
?_?9=r��Dˈ<~8��G��wj�����3ǎ>$׽�:�&M��f�4c
?%?����Y]̾�B׽�Δ� �z=L|u?��3?.�)Z�t�i� $=���V�`[�����dӾ�/�k�j��j��@8��pz�b,��OV��c0?�5�?�/	�Ө�L�Ⱦ�7[��:-�Ϋ�>��?��>��>��S>��񾶐>�xb����g���>���?3G>�bb?
u?��n?�[j?Oo>&J�>�!���C�>��>�E�>���>��2?#?P�;?��8?4;?<k>�SJ��~�ۗԾ$�-?��?��?��>'�?��/�����&\���%�23�;���=�G7>��>V��=����_�z=��>�[?ס�ʭ8�����k>�7?$y�>���>�	��0,�����<��>'�
?�=�>�  ��{r�]�$a�>š�?=��=)�)>���=ǧ��v�ϺIS�=����ߐ=OV���;��<W��=�=��t�"����
�:ia�;-��<� ?�u?#��>0̈>:7��&��������=�[>��R>�1>4�پ�v���1����g��?x>z��?���?`Ql='5�=��=�b��y8��3�����O��<��?#�"?�@T?�V�?��=?�r#?��>p"��A���>���ã�a�?�,?w��>�����ʾ*⨿�3��k?�D?�'a�	j�5J)��Z¾v\ս"�>�Y/�~�>��<D�(ו�Z��Jƙ����?�ʝ?iB���6��;� ���z��!gC?D�>+A�>m��>��)���g�O#�K;>�o�>�R?���>.�O?�w?5W?dM>�_7�<���2��Z����g&>:=?\�?yT�?�*y?W.�>�>��9���������ԯ齊��)=�4^>m��>��>��>��=�������HK�r*j=Fva>{,�>ƥ�>D�>X��>�@w<}�G?��>�־�S�cB��R��d-�K�u?dA�?gF*?od=8A�gE�.{���?�>9�?D��?�8*?buR��[�=�Kռ���p����>�>e?�>�o�=�MG=��>7�>��>�����
�8��LI�R?��E?�N�=� ƿ`lv��Io��˹�Mm��1$��%D��9)=^V9�˽6<Y���;$z��(z��0�1�r������Ѿcc���V��?��y9���=�J1>B?C>��=SjA�&�=��N=v;ݽ�Ւ���$=�H�P����U�&=����'1<`��<�n˾B�}?�/I?G�+?*�C?�y>;z>�K4�ON�>Ԓ���$?��U>.GQ�H���/�;�߹������4�ؾ�{׾�c�o����>��H��h>33>'��=Ka�<0��=��t=��=��[�kx=3 �=pO�=t�=��=��>�'>�6w?X�������4Q��Z罥�:?�8�>d{�=��ƾq@?��>>�2������yb��-?���?�T�??�?>ti��d�>L���㎽�q�=K����=2>q��=v�2�S��>��J>���K��A����4�?��@��??�ዿТϿ6a/>��7>�G>޷Q��1�N�[�=[d��a�[?WX;���Ǿ���>�Ԯ=�W�����?+=jP->Uz/=Ϙ���]����=�s��J=�FW=��>��B>F�=0����f�=#b=���=*3F>����=�5/�ɖ(=��=bc>�U$>���>z`?�.0?��c?{�>Wvi��(˾�[��d~�>��=Ű>b�=��D>�4�>��7?�YD?��K?XR�>�ه=E��>Z_�>��,��l��|澅����/�<��?�{�?e�>�tn<)$?�L��	�>��)Ͻ0?��1?��?��>���iؿ�f���Z�R�̾�� �&��;k��e���Dw��qľ .���Ռ>��?H8�>��P>@�= l�=�v>�߮>�%0>�)�=�E=�� >"�(>�����?>��b��"�������;���=�ঽЃ��ʽ�|߻�=������=r��>�>���>���=/�����0>���ҾL��I�=W��:A���c�e�	0�ti7��C>�HW>��}����S�?��^>��A>��?��s?�!>b����־[ԝ��>h�{�U�k�=+g>��?�4W:��;^��O���Ծ��>xk?%��'�>ɟ����O�C4>�����y-����>�;ʾ>�=x��❇��D��su����R�Hj�=@[\?�j��$U>KB�?�
i?�?�a�=u��=��(��Ø�Y�ɾ(�¾:9��X$���G����>��&?}��>W�@�u��8Ⱦ�Ϻ��t�>;+<���O�c��Q0� ;�#����>��QmԾ	4��V��3K��_zB��Jr��>eAN?y"�?��a������N�}+�^o��*�?�h?+�>�?�?������c���i�=�j?���?���?t >W��=��Ž��>�J�>p��?���?�t�?�5c=��>D�u�^�>���\E�>Dd�>�˃>��<>�?��>��>{��<�%���a����z%���>�=[E,>|�k>��,>$>Ʌ5>h��=L�>X��=Ү�=��b>�E�>Jv�>8|�>�*ƾ��i�?��=���>�H?�c>���=I�-���޽Md��.�I�BTN���ݽ�׽��X<�&���
<U�$�}o?	�ÿ� �?E��>�6���?b��rõ�>졆=�����?a�C>��T>�ӄ>�N�>L>mC>��6>����R>��T'��;A�qg^��wҾ%٣>���D��O	�H\]�����/Ѿ�H�&sa��u��@<���<Jy�?z���Ȣs�XN'��d��� �>n��>��D?�,�9@�<�V>��?�՛>d�F���n�پ��?@��?�/c>�7�>K�W?ϡ?�S1�'3�ubZ�'�u��&A�O�d��`����������
�]`��|�_?��x?�bA?�}�<�+z>���?��%�����%�>K/�);��==�<�>�氾�`���Ӿɕþ(��F>٤o?Z"�?]I?vMV��*ٽ��N>]҄?�VH?=�?rt?K�N?�a�ё�>�<Ƚ�>6�?�/?��-?��K?��??.�n>j ��?�=0v?��'����X�靄�%a�΀=i�m�?;j�=Q�7=�Q4<2��.��"=�m���L���y�<�~�<�cg<ɭ�>G�]?7p�>ӆ>��7?����H8�)�����.?�<=����5������4��S�>��j?��?+Z?:�c>r�A���B���>Fy�>��&>E�[>QO�>�olE��@�=��>rj>`�=��J��&��\{	��2�����<\�>��>{�|>i��&�%>@���jz�H�b>\�Q�l���#;S���G�h\1���v��$�>��K?�?�3�=@��􆙽f���(?Pc<?��M?�,?ƒ=�ھ�*9�^�J����k2�>�;�<D	��٢������:�H$�:6as>"?��e��ml%>)�li�� <�iF�M�1�d�����־�a�> ������ߕX��=f>Y�����dS(� �����A? e<I����5��{���!(>Tҳ>���>��K=�<"�%��ꤾcS�>�-k>8�>�q�܃�����z���˄>f/E?Ѳ^?�˃?�Ѐ��_r�t�A��m���m��O����?o7�>�w?3�B>D�=VM����%�d��UF�c��>R^�>���1fH�.���qj�w#�ы>��?�>%�?��R?��
?��_?��+?D�?�K�>뷳����<A&?w��?*�=��Խ��T� 9�F�A��>�)?��B�|��>��?��?��&?p�Q?��?y�>ƭ ��D@���>�X�>V�W��a��#�_>��J?���>�<Y?bԃ?�=>ń5�袾�ͩ��O�=�>,�2?�5#?��?b��>���>�&���؃=���>Pc?_\�?)p?�B�=�X?�K1>���>���=w�>.�>"o?wAO?�{s?�J?���>#��<�S��]鶽W�q�y�U�9�;�F<�x=�j���q�}�e��<ă~;���Rz�Ǳ��i F�쐼���;u��>��>���	4>gý�*��׃A>wT���"�����(6>��{�=Hpy>M��>/n�>��'��=�w�>���>���>�%?P+?Z0?Ț��J�_�پ�jS���>xe;?��=JDk���$�w�άV=�#k?c\?"�h�*���g�b?.�]?�n�m=���þ�b���龌�O?��
?��G�B�>`�~? �q?r��> �e��:n����@b�k��߶=-m�>�W���d�;�>p�7?`F�>�b>?/�=�q۾^�w�ji���?��?���?��?*8*>U�n��1࿳'�YZ���g?���>����X*?Q��<�վ'���!,���¾�k{�~F��Ma4�Q���
ҽ�v���8R�7�r=�?+�S?.,�?��q?�%�dko�􉃿�-��)Fn�꾠��g��X:���.�SZ������6 ��R���<=n���7
V��T�?�/?�N�o��>�������ﾳ�m>�Һ��d�=1��f��<�w|=pv��t�h��&���,%?�R�>gv�>�@?	5U�H�S��qZ��vH�&�	��� >=�>7��>�l�>\Ԁ<<������2ξ�w�������3>�SN?"�,?t�Z?�����1������R����i���>I0>6t�>��4�Z뽿�0�h;B�n�4��lE��h�����=�`;?jsL>���>u�?�
?a���˾�X��xE������a�>�qm?x��>�:>x��g�
��I�>K�m?M��>F{�>����A!�Fx��KȽn>�>Mp�>�t�>�Is>m�/�]�ſ���u��:7����=F�f?O���q!a��ڊ>[�T?ȵ�*D<�>�E����������9���>"1?���=��2>Ԟľ��	��}�Z����)?��?	͓��+��Q}>mr!?���>B��>P��?�r�>p�¾Bؠ:�%?��^?�xI?�!@?z7�>�L=����6�ǽ�b&���*=�>[>~�c={��=�"�8]\�c �U@=r��=��̼����<� <�S���]X<)F�<�2>�gۿ�8K�f�پ3����D
�6��++���g��_��eM��'�Kx�tf�A�'�V�.ac�m�����l�r��? 5�?_���zH��먚���������<��>�[q��������������Z���r`!���O�;i���e�N�'?�����ǿ񰡿�:ܾ4! ?�A ?7�y?��8�"���8�� >KC�<-����뾭����οB�����^?���>��/��p��>ܥ�>
�X>�Hq>����螾z1�<��?5�-?��>Ȏr�1�ɿa����¤<���?0�@V�@?�%(����n8=��>[�? :7>�X7��f�]X��� �>+�?[�?@U=�lW����c?п;g�H����y�=��=�p=�*���C>D3�>�����B����92>�9�>t�*�C?���]�<y�<t\>q�׽�M��5Մ?,{\��f���/��T��U>��T?�*�>V:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=n6�����z���&V���=[��>d�>,������O��I��W��=���ƿ��$��{��V=��ݺ�[��|罤���U��"���ho�Շ轃�h=���=�Q>Xi�>� W>�2Z>�eW?v�k?�O�>�>�7�F}���ξ�E�zG��N��������r�R��߾?�	�'��(����ɾ��;���=�N�'��(���	d�FM�Q"?M�>�꾾�RG���=\�¾ۙ��>h'��w����Ҿ �1��bj��?�n>?�p����W�y�
��w��놊��cR?C潁?��uͭ�U��=~"�����<X��>qS�=i۾��+�/�R�}�/?�e?/4��Ni��D�*>0��[s=�*?- ?ׇQ<ְ�>��%?h)�����X>*a0>*N�>Ð�>N�>�㯾<�۽M�?f�U?�>��@��>b����y���L=8�>��5���3�V>g?�<����)�i������ݷ<�;j?/��>�
=�9�@�P���V��=���=��r?�m?k��>��^?��?8@w�׭�MTO�1���m�<>	�n?�}{? �@�L�s>0CӾ��n�i?��9?z��>���L)��V۾�ä�\� ?���??Q7?*���ʙ���������]^?讘?��o��Η�H��x�{��="��>�>6���F�=Ģ?��7���a���� &����?�@5�?{k<��
=��)=��>e�$><1=��Sd<�ۦݾZ>>rZ�<���vo3���ʾb4��k?o�M?�k?}��j��+�=�3�� ��?�.�?�9��f�[<M����l�� �~�<o��=�3����%�G�7�Uƾ_�n���ü��>�^@*P��E�>)�7�rZ�6п�(���о�pq���?���>��̽m����k��u�-kG�Y�G�%o��{ȡ>2>�疽�L����z�~�;�ڼ��>*���>�P����|����\<�}�>9�>�$�>���@����˙?T����~οt{����dX?C\�?�?��?֟<[yw��~�͟����E?��s?�3X?����iW�>J���i?�à�-Va��6�@{@��hQ>O3?#S�>k�.�<��=�>Ǣ�>>(R.��zÿ�����8��?Ĉ�?�\���>�<�?
0?�
�e��D����%+�* ��)<?�$#>R����� ��1>��돾��?N,?�[�gs�\�_?*�a�J�p���-�l�ƽ�ۡ>��0��e\�)N�����Xe����@y����?N^�?h�?ص�� #�f6%?�>e����8Ǿ��<���>�(�>�)N>nH_���u>����:�i	>���?�~�?Qj?���������U>�}?�ޗ>�aw?]I��&�>==$>���*�۽L��=	��nк��>�1Z?j�>��U=Nc���-���5�F�/���޾QD���X>+m\?S5y?c��=s���ѹ�9�Z��;����1��o���U�����)�U>��>��W=>�������?Vp�0�ؿ�i���p'�i54?C��>+�?���ٳt����;_?�y�>7��+���%��-B�a��?�G�?K�?��׾U̼�>%�>�I�>@�Խ����.�����7>�B?S��D��m�o�v�>���?�@�ծ?[i��?x
��H����l���n�iK>7�M?I7ϾZ�>%?��<�c~�d.��K6t�g �>�	�?>�?�q?u?��r���I�@/L���p>��W?k?�y�!�;�5g>�I ?D^�������WW?n�@�Q@PRo?�i����Ͽm㚿/��鄼�1�=�f9>��}>x$O���>hw�=�6�=u��5>���>�ߊ>[)N>O>�h�=S�>����Y%��������L3V����9F�D"��>� �`=�Q���Ə�86;0����<���2�G�������u����Ɂ�B�b?)�b?:S?�Q?m�<߽u>�}��A�T���:>n����>��:?�m8?!mS?��T�n� Y��\�{��"O:�H��>ٌ�=П�>�%�>�B�>3�3=7X�>�k�>M�?p;`;�=�0>z�<>j��>Q=�>�� ?���>@<>�>�δ�71��Ǜh�Ow�p"̽6 �??���λJ�11��8��A���0j�=�a.?w>���}>п���� 1H?����(�Y�+�)�>��0?dW?��>���"�T�V:>8����j�"\>G( ��}l�V�)��#Q>hl?®X>�]k>��3�O�6�S�M�?U���>^>� /?������6�8�p���B���Ӿ�M>�o�>x���}��}��O�}��m�Cts=��9?�?z�թ��\����DD>�E> 6=��w=p�->����m��c�<��=�+�=?�g>�?�b,>��=�H�>�����pQ����>uA>+>��??,�$?�}
��p�����EN.���u> ��>���>�>B�J����=�x�>�c>�`	�_��dv��)?��xW>ȁ� �`���v��'t=a���@��==�g �w7>��;$=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿh�>]x�vZ�������u��#=¨�>�8H?�V��j�O�!>�w
?�?�^�ܩ����ȿ7|v����>6�?���?N�m��A���@�k��>(��?�gY?oi>�g۾�_Z����>��@?�R?��>�9��'���?�޶?���?��H>�B�?<~r?3��>ew��/�Y��������=M?�;Y|�>l>�"����E����ab��Qj������\>&$=�}�>��㽧
��G2�=o���d;���q`�u�>�$p>.�G>�Q�>(� ?���>���>d={D��U6��|��K?�Ԏ?!��{o����<K&�=Q�f�1?��3?�	ѻ��ξLl�>�I]?\�?��X?x�>+��{���ht��R��p�<�#K>b�>�K�>����J�H>�оf�E��'�>;ߕ>xv�ھK?���oǻ��>�| ?�o�>aG�=Θ ?(�#?g�j>&�>b`E��9��Z�E����>���>[I?z�~?W�?Rӹ�+Y3����t桿̒[�K8N>��x?�V?�ɕ>ҏ�������nE�=:I��뒽���?ktg?EK�@?E1�?��??;�A?L-f>݊�eؾߡ���>��!?T����A���&�"���??��>~А�.�νA�Ҽt�~[����?Kf[?+%?���l�`���ľ��<#��x�U��;�r;�A>)N>;�����=i�>mr�=]k�!#5�M�S<�ں=�	�>���=�D7�v%��.>?��k��`�������o��y,�D�p>��c>�v��E?]W5�bUy���������p�u��?�{�?�{�?�f���Eb���G?Q�w?�D ?]g�>z!��|���䳾�+��s�޽({羰wT>��>^D�=�O�ƣ��m�������D�<�)F�� ?X��>�8?��>�T=ٗ�>2w}���������\�!�0�O�־"j/��m!��G�t���պ����5�l���!�w���>�!6�r I>9��>�v�>=�>]�>�Z~�%�=�d->���>���>`,�>�2����.���콉?R?����'�'���辇���sB?�Td?9�>�ui�_��������?���?Wm�?F#v>�}h�(,+�}a?�(�>�(���i
?:=�
���<GH��B���Ά�#��G��>�7׽�:�wM�f��m
?�%?�^����̾a�ֽ��v �Jd�?~?�O ���R�7Ώ���v���`��.=����z��	��*&�p]����h��H��p�3��k�=�`8?~��?��H��J.�����t�g�T��z!>1
	?�1h>���>؀>Y����&�>Ac��n�����Xz�>(�X?���>�I?nH<?)gP?��L?��>�0�>���A��>��;mӠ>���>:�9?'.?�0?�z?#++?|+b>�#�������Sؾ|�?W?�?u/?��?������Ľ� ���T�GHy���{�t�=��<Gֽ�q���W=�T>�&?:}���8������@j> �6?���>���>�W���9��p�<2c�>�?�y�>D�����r��T����>�?����:=�)>T��=���8�EH�=ZƵ����=k����>�d]3<|B�=ϒ=^ы�����q1;��n;���<N|?H�?�&�>횅>�V��������<
�=�Sb>��M>�>��ھ����V���bg�?�>�?���?$�]=�;�=�U�=�D���뿾�R�ȯ��t��<�?R!?c�U?̑�?=�>?�$?�w>����D���؅�����kF?�,?���>��ܹʾ*�6�3�p�?jZ?�<a���7)�j�¾��Խ��>�Z/��-~�J���D����g���h�����?���?��@�?�6�ko�4����_���C?��>1W�>4�>��)���g��$�9;>%|�>�R?R�>�cM?��u?�U?��P>t 8�db��Ȅ���{�J�.>uQ>?nn�?��?m�w?�(�>�>��,�X�߾�� ��Jn�㇂��^J=ʇX>���>�@�>�I�>���=gν?ݵ���6����=�g[>p��>n�>���>��r>ʔ�<��U?�k�>3$վ#9��׾�-����X���v?�[�?^
+?
�=�� ���V��&
���>5X�?�a�?�#;?^��|u>�<��{���:��D�>���>ҍ�>�V�/��=�&>���>���>5��,	��(��罿�?"�B?�ʺ=�'���bZ��Ȅ��e���ͼ����J䇾iU̽s��a�>;I����d�������1��������P�־�����o��?!�>�n�=W=>&/�=�2�<�v�<]�>�8 >|�_=��������ؽ&'��|�I ���t=~8|=�j�=��<�˾y�}?�,I?>�+?��C?�y>�>�K4���>zM���8?/$V>��O��u��ou;�3����%��ѷؾ�׾��c�0���H>ruI���>�&3>�A�=o>�<7�=c�r=�Ŏ=�%R�J=� �=�1�=%��=��=V�>[A>8w?h���β��5Q��f�յ:?�7�>�|�=Lyƾ�@?s�>>3��͗��{d�w+?<��?�U�?_�?Oxi�c�>E���⎽l�=N����@2>���=��2�䠹>��J>u��I���o��4�?��@��??�ዿݡϿ�f/>B#>�q�=��R�ud7��W�Kń�jj��ʌ?��2�k���-r>@�>,Ǯ�#���5�<�#�=o��;�6���g�ߙK=�Et���=���=��x>�j>�6�='»�>d=_�"�=��>>��e��U�����L�f=_t�=1�@>*?>��>��?�^0?�Vd?r0�>�n�_Ͼ�5��?�>���=�C�>���=odB>,��>��7?�D?E�K?�|�>Nω=R�>��>�,��m��t��ӧ���<���?�φ?hٸ>�kS<@�A�ݡ��i>�VfŽ�{?�V1?�q?l�>�U����6Y&���.�B�����4�]+=�mr��RU�����Cm���㽉�=�p�>���>��>Ty>��9>��N>z�>��>�7�<�p�=*������<����δ�=������<hvż������&�t�+�!�����;���;Ǩ]<���;a�>Q �>D�=�0�>�i�=�f���<>�N|��RN�2B�=�S����8���[�èx�\0�Pv8�t::>�Px>���< >��^�
?��f>�t>
�?�V[?�q->I�{c��͚�9f|���0��%�=�|�=5�5��@�Kd���R�j�Ͼ��>ٲ�>�)~>�L>�z��+=�\�=\Ǿ'�=����>}��|���gl�E��'���_`����<lL?u���xr�=A
�?�*c?㢈?�ۭ>��������!>_Ѥ��*o�7#
�N����"��?�?���>�T�b�O��^���Ľ�q�>�&��uNW�H势����v>�}��
ڋ>�tʽ���`H9��Kw�����01	��^��;�>��[?i�?E�������1:�ٿ[����q?b��?#+�>��E?ȝ:?K��= "����TX��f�?�X�?��?H�>��=��o�?t�?���?,�?�no?)H���>]�6�Q�>T����->��e>E�9>lt�=���>�k�>1�?n����
������8WF�>�0=ч�<ҧ�>�r>�@v>�R�=$���\��=��>���>�$�>-MG>`�>��j>�Ǧ�_��&?B6�=��>!22?�r�>�\=�k��0{�<�{K��A�� +��t����ܽ�ҳ<�Ȼ��G=�ʼLV�>
ǿ��?J�S>�g��?�=���&��T>�U>�Eܽ�s�>��C>t�|>/X�>���>>�n�>@�(>�Ӿ�>}�Q|!�bB���R��վ7s>0����$�mr�ߣ�Z�G���)��$i�1���N=�y�<��?d�����l�O�*�����ݪ?h�>�p5?�,��Խ��
�>�3�>�P�>"���߻��0���`�/��?���?�7c>6�>�W?]�?�1��3��tZ���u��(A��e��`�p፿������
�|��l�_?��x?iwA?-S�<c;z>���?��%��Џ�?'�>�/�o%;�N<=�.�>�(��$�`��Ӿ��þ�:�{@F>�o?%�?�X?uRV��:)��D�>��k?f|J?�T�?�{?�TV?���=��>�F�=J��>��>4�L?��W?�\k?lՏ>�=�ܺ����=�l�;����J�	�P;h��qR;�1>�G�=�ƚ�YQ+�
1�=6�d=����P?=�[>Q�J<���<+$=*+=��I>r��>�]?A�>��>ʾ7?��QK8������/?@e6=�>��e튾&ߢ�tn�i#>��j?��?�3Z?��c>�A�[&C���>>��%>�"\>�,�>(��ND���=%/>�>ς�=+*L�-����	�.L��7¼<B[>���>hC}>^���Y+'>0颾�>z��d>�2Q��1���S�N�G�Ȝ1�.v�_��>�K?'�?��=����=��MMf�$)?]q<?L�M?o�?�,�=Ơ۾�9�L�J�b%��3�>��<Y��/�������}�:��yR:� r>�����䠾Rb>����p޾��n��
J����.M=-~��jV=\���վ�;����=�
>����6� �L��7֪��1J?��j=`t���^U�on��8�>-��>�>ӹ:���v���@������,�=��>�;>z��~ ﾦ}G��7����>�C?|�^?�f�?�kz�Js��&A��Z ����1���K?E�>��	??H>(R�=r����e�y%b��E����>\V�>���iAG��e���T����"����>�r?|�>�?�IQ?(=?_�_?u�(?�?��>jݝ�Â���A&?<��?��=c�Խ��T���8�+F����>��)?ϸB�y��>��?ܽ?J�&?��Q?5�?��>� ��B@����>gY�>b�W�Jb����_>-�J?���>�=Y?�ԃ?m�=>�5�颾�ҩ��S�=�>�2?�5#?�?P��>RQ�>O�����=A��>�c?(@�?_�o?H�=��?��1>��>�6�=� �>��>��?O?ls?�J?��>t�<X<�����S�q�oD�eD�;y\G<qXw=�+�^�s�j��Ev�<� �;���S+��c����D�	L����<%��>�Xt>e]����/>�ľW���t%@>A㟼�f����$�:��!�=:��>�?Ӈ�>�>"��|�=S�>K��>�����'?s�?�)?�/�:�b�}zھ�2L�E&�>|B?��=��l��k����u���c=־m?�Q^?��V�y��f�f?y�P?C����?�f&Ӿ^�B�0?���CV?��?5�W�Ae�>���?��{?mL?��v���w������W�w�)� ��=���>gw���b���>�SH?���>�V>��>ɐ��ϳ�A���+?34�?a��?(#�?��
>�wp�g��ծ��?��MW?�Ƨ>g���&#?�񽃇۾(E���r\����_�����2䮾������l��7����g��>.2?�U?P.V?��/?D�+���j�D�B�.�@q��%�o� ��b���E���E��KG������Ҿ����C;>j}���A�c�?��'?��.��V�>�����𾎮;KkC>����B�;�=�_���<=%W=�h���,��୾�  ?q�>{*�>�<?Ѳ[��>��)1���7�BA��x�2>hˡ>�u�>66�>�h�:�F.��U�)	ɾ�����н�v>sc?��K?��n?��w	1��}��	�!�\�/�e��3�B>[�>pω>�iW�/��2&��a>�A�r�L��ln����	�h�~=;�2?�$�>k��>J�?)?��	��S���"x���1�nC�<��>�	i?
C�>�>�tϽ�� �V��>��l?��>��>陌��Y!���{� �ʽ�$�>s�>C��>2�o>��,�� \��i��~����9��Z�=��h?����G�`�E�>]R?X��:S�G<�q�>�v���!�r���'�#�>�|?|��=�;>S�žN'�8�{��:����,?�?&�˾��9���`>�<?���>:}�>3Px?(�">YZ��M`۽U�?�$i?�}?�N??��>���&�=Qg����)�t=C�>�!�>U��s�T�g"�=�����5�}v=_	>��==�:���e=�~����
=������{>�tۿ�RK�?�پ�����
��s��n紽�!�����h���S��6�y�/	�g-���V���a����� m�U]�?:&�?Qm��:5��d��"k��G������>G,q��y����l4�¯���䞬���!��O�Ki���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >`C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾}1�<��?7�-?��>Ŏr�1�ɿc����¤<���?0�@:A?��(����]�U=���>·	?r�?>�1�/E��᰾�5�>:9�?���?�"M=9�W�W�	��{e?̀<��F�.��)�=yc�=:�=��luJ>�A�>[l�4qA���۽S�4>�݅>8�"�����^�Y�<��]>�iս���r�?��X��Uf�BD0��~��3>	�Q?�o�>I�=Yl)?�bG��Ͽ�Z�n�a?���?�_�?T>(?�¾`��>�]۾��J?a6?ւ�>?V%��t�:5�=&B���s�)+�qU��,�=���>�>�w-��%�JN��凼u��=��&�ſA�7�����+D>-��;M�n��ƀ�cw��J �E�����y�LB�]�ܼ@��>9n�>n<p>�6>��U?p��?nu?���>a���繀��ﯾ��0��=?�J�<ɏ��M�������Ѿ�쾔�"������1�&��
!=���=�6R�R����� ��b�,�F���.?�w$>��ʾm�M�
�-<�pʾ/����݄��᥽�-̾�1�+"n�T͟?x�A?������V�'��"Y�K���A�W?GP����Sꬾ"��=����ȟ=%�>Њ�=?�⾰ 3�D~S��A?��?����uȾ;�=&t:�H�I>jC?z��>��Y>x��>�n ?����O0�;>W��=���>�O�>}_�=;X̾K�X���/?�Pq?&Z����o4<>c���舾t�3>��<�S����U��=�{��/�Q���b �h�H>Lc?tWj>�,�W-!�_jľ��"��_@>�?q~?���>�nt?biF?E >=�ݾ��X�<�.����Oa?!��?��?>��DZ侯��k�1?� �?��>�O*��ϴ��uh��
�~�/?:�?hC?�==�ɂ�˕����#�"?��v?s^�ws�����M�V�e=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�%Þ?��@���?y�;<��T��=�;?k\�>��O��>ƾ�z������5�q=�"�>���~ev����R,�f�8?ݠ�?���>������q��=�ە�Z�?s�?k���D�f<����l��q���v�<,ū=�$�vd"�\��^�7���ƾ�
�g����������>PZ@aY�)�>�G8��6��RϿW���[оWq�,�?�v�>��Ƚ垣�X�j��Lu��G�X�H�����jU�>9>'ך�a���`y�®<���뼈��>Frμ��>q�W��绾Sޢ�Ɋ��>��>1 �>1➽�S���x�?�����+ο՜������dX?���?.��?�� ?vD<�r�N|��wN���H?ؕv?W�\?|/���n�WhE�*�j?G_��mU`��4�oHE�QU>#3?"C�>+�-��|=1>���>@g>�#/�`�Ŀrٶ�����7��?���?p���>y��?�s+?�i��7���[����*�p�+��<A?�2>����<�!�=0=�vҒ�ü
?~0?
{�$.�v�P?�X���|��KD������U�>8�D�����=T��}�J��N��Pd�?x@�)�?"���B*���'?_@�>�K��Q���� =+F�>���>�؇>��#=(B�>�[ѾG��>�C�?Ͽ�?�H?�υ�=ϙ��0�=kLp?OF�>w�?��Z>�9?sw��嶺�%z=|�|>2k�=b�=6��>ԻF?A2�>���=T<Z�O��_sD��e�T���K� ��>�w?�/V?UiK>&἟<�����a���ؾ���;��~"�=�	����<>P8 =��i�}��B{߾��?Mp�9�ؿ j��"p'��54?0��>�?����t�����;_?Qz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>@�Խ����[�����7>1�B?Y��D��u�o�y�>���?
�@�ծ?ji��	?���P��Wa~���7����=��7?�0��z>���>��=�nv�Ừ�C�s�۹�>�B�?�{�?!��>�l?t�o�^�B�F�1=KM�>ǜk?�s?*Do�;�#�B>��?#�������K��f?�
@u@C�^?#_׿vѨ�O���$���DE>/��=�q�=h�o��>T-��XN/�!]�¸7>�܀>�>���>q4>5��>��>�"������:��R������
���.��u��Y>��ߤ�����/���Ӳ�;�ͽ�%�7o(�rè�d1�;���5�=��T?>W?p%o?V� ?%�$���>��G��<[�0��Լ=���>�:3?�I?��?L[=�w��?�_����]O���ʏ�C$�>I4I>��>�<�>P�>*��<[*1>��7>
˃>��=W�<఺���<�5U>V֫>p�>�/�>cR<>3�>Cϴ�c2��h���v�?�˽� �?v����J��/���1��A���{��=Da.?�x>
��&?пe����/H?T�`(���+�\ >û0? \W?��>|���T�+H>����j��S>�% �M|l�Շ)��)Q>k?�3j>u>O4�y9��P�q��>\�6?��'�7��ft���G�.o۾�uO>R*�>؁G�@i�9ꖿ�
�#�i��8�=�%:?�o? V��������v��~��1�M>�{^>�=�٦=%�K>��k�O�Ƚ�kG�9�6=A�=�>`>�p?��F>��"=Y��>1s���Qa��p�>4mk>	R4>0�R?R�$?�v�0nV���o��@�Ůd>2�>�7e>��>����)��=��	?�g�>��/���\��rT�tn��1L>*��lǄ��mo�vD=�sҽH]�=�"�=��F��DH�[��=�~?���'䈿��8e���lD?P+?� �=p�F<��"�= ���H��C�?n�@m�?��	�ڢV�1�?�@�?��ѷ�=}�>׫>�ξ��L��?��Ž>Ǣ�̔	�[)#�cS�?��?i�/�Sʋ�-l�i6>�^%?�ӾCR�>g�!�M����冿��y�{�=��>Z1Q?�Nݾ/���{��?�@?��ؾ�p��@U̿{�x��G�>��?���?~,p��;��.VB��x�>���?�h?��b>"���*����D>{�I?[�P?]�>������T�>���?2	o?��H>^��?�s?���>�tw�a/��)������=~=�P;9��>�>C���BGF��ѓ�j^��P�j���1�a>G�$=��>EC佨>����=/9��D����f�@��>>q>ȲI>�V�>�� ?�d�>R��>r�=2M��ϱ��d���~c?'r?`D2�����ڢ�0϶=�<=��&?�,H?Q3	=3%i�@��>m!W?�}?��E?�J>Wʾj����ſ�,��@	>(D6>(�>&?��n����<*Xu�$��*��>���>�9ؽȯ˾iϦ�:�<�]>�6?2s�>��@>�>)?ѱ�>��I>��>v�f����ٰ�W`�>�P�>b@j?�m?ʼ
?������M�A͓�ۃ���M8�U��>��?-G??u|�>�T��Ƈ���7�څ��}H>$�?E/�?.�-�J"\?k|?5�l?�bZ?Z�>�Ⱦ�0׾���3G�>M"?ܽ�oD���(�!���?sz�>���>
u�����D���u�b�꾼W?Z�f?w�)?W�����c��'����<Й���!<�R�<������=d>Xj��o=a�>��=��r�K�4�g���V�=��>#�=��'������)?�(¼�_�|%�=��p�NpA�ik>��?>�,Ծ	�^?!~��)r�V����Þ���C��5�?�I�?��?�벽�f�R96?ֵ�?Z}?F�>�U��ݾB�Ծ~�~� @y�'���<>2b�>��v�Ֆ���1��b�y�Z�Ͻ8	#�!o�>���>0l?�;?�3P>o��>�����&�'�uw�)�]�����8���-��]�)���V|�������-|�I�>e���렲>=C
?/h>�|}>�V�>��˻-�>PT>|~>돤>�-W>V.3>%��=nU<v$ʽN�r??j�y@��4%��)��rv?�X�?Eu$?��>]Y������o,M?R�?���?�k>jf��FL�ؠ�>��_>~�W��?G����,�&�<W���b�|��8�h �=A܎>�佉�.��mQ��'�s<)?�E?�>�*��� ��������<}܃?�'#?M(�=CQ���n�?\��W�q���s�Tɪ��#(��Pt�����;���3��,�&�OQ�=Lu+?Ў?I���`�/1����s���;��e<> 2�>���>�`�>.�=Y��;6�;DS�͌��,B��� ?Y{w?�f�>�xI?�<?vP?mtL?���>P8�>�����#�>w��;�?�>#�>I�9?��-? 0?[Y?y/+?"c>�w��!���y�ؾ��?�?"/?�?��?�_��,^Ľ ���a�F�y�񘂽�x�=��<��ֽ�s�ޔV=�S>W?%����8������k>��7?l��>���>]���$��IM�<a�>�
?�D�>�����yr��]��O�>���?��,�=��)>�!�=����߄ۺ��=O�¼���=@���hY;�R�<$��=j�=��w��Y�����:vJ�;�P�<��>�<�>s�>���>�⍾��gb ��]��y<$��%�>�Ŋ�P��Cd���f��%�M�T0+>>��?OD�? C>�2>�{>�۾{ ��_��*���&<>r��>��7?��i?�ƨ?�a?��0?w�1>�H�;����|s�)���z�:?"",?���>���{�ʾ쨿-�3�H�?(V?A=a�u���7)�¾��Խy�>�@/��~�����eD��̀������-��?���?��A���6�L_����pm����C?���>�U�>���>��)�$�g�P��;>���>x�Q?\{�>�M?�Yz?�Q]?�iW>�:��f���f��>ؼ�P>��A?q�?��?��x?��>�>a9+�� ھr�����M��]h����6=�S>���>r�>)��>�1�=�ý�*���9�{��=�e>��>�ͣ>:��>��><�<��G?���>�s�����ा9ۃ���=���u?���?�k+?hL=�w���E�������>e�?7�?\*?�KS�C~�=��ؼz����mq���>�}�>,)�>'ɓ=�2C=Z�>���>���>�H�Uh� s8�F*N�_�?F?���=��ǿ��;�li�eg��=��>�4���	ξ3��nԁ=��p>�U� ɾii�G0���$ɾQs̾�؅�*[O�B���5�>δS=�B>���=hn=��>R�=�f>s�)>�3�=���p�;�7�<�uE����=�*5=5��oV�=YJ:݋��mYT?�g?��J?��+?x�>	T�=�A�=��>�ii�o�?��>��p>�T��eÙ��#��d��Zľ0��zU5��灾8_=�U�+0�>Ʈ=�)ѽ�J����=k�~<�>S=�=C�
>$�#=���=� �==�C>��=V�Z?�%����3to�����{`�>�U>=,񪽣�G����>�_�==������)S�ɇ?"� @���?�7�>{��M��>nq����e�]�m=a���T��>o�>�؂��s�>Hz>�� ��͊� Z^�_��?�@q�L?q5��{:ӿ=��=w B>|&>��S�8�3��9a���c���L���#?�7�K�Ǿ�+�>���=��ھ-����5={U0>��=�A���]�%3�=��i�k�J=���=L��>��<>�m�=N䪽���=��o=�`�=R�I>Z�һOH��F�g�(=��=ϲf>D�0>���>��?+b0?�Zd?�4�>y"n�AϾaD���6�>��=�F�>B�=�zB>֎�>�7?j�D?��K?.��>vÉ=;�>��>��,���m�ue�Hɧ��L�<���?s͆?θ>�!Q<�{A���2c>�Ž�p?�N1?�m?}�>���v���K6�� /����$<uZ=�����ֱ���)��?���"½9x�=^��>�>��>ϋ>�f>2�I>���>�">#�Q=ށ�=�S�<�Қ<����l�<\B��%=��ɼ����(�c������(��*�u�[=��T����<���=��>�#>.��>�c�=!���y�(>�Ɩ�+O���=*����L?��d��"��F�,���0�]�D>��f>�"��E���k� ?e�_>k
B>]��?�=t?��>���
E־DV��2�p�#�=��=�;�=�D�+�=�ؘ]�YsI��Ҿi��>���>d�>��l>#,��!?�E�w=	��_5�s�>A~��!��X)��7q��=���򟿯i��ZϺ��D?�F��2��=e%~?��I?�ߏ?a��>zH����ؾ10>=O��$�=��(q������?0
'?z��>��n�D��dǾ�-㽲��>�<��
O�ɣ���;/��n��6ľЮ�>
����Ҿ6�3��?���f��t�@���z�۸>�AR?���?�&��� �K�#Y�B��M>?m�`?�g�>[p?З
?����Gܾ�ޅ��=��j?-�?_�?	>>���=Rµ����>�m	?4��?<ʑ? 7s?�7<�QB�>ȹ};�">�\�����=5>¼�=v��=�?(w
?�'
?���L�	�|����d�\�pd�<`�=�>r��>e9r>Ә�=�Df=K��=0�Z>�0�>�-�>Y�d>���>���>1�¾����@#?Ӗ�=r�>�2?Sj@>f�<�2�x=�N�Y�*�܊+�����?���~�X>��X;Y=~���H�>��ǿ�f�?���=&�V�?��꾾|4�?V>��->4�,����>�#�=j�x>�ѡ>�>e� >�G->rUQ>�FӾ>����d!��,C�L�R���Ѿ`}z>����F	&����vw��dBI��n��zg��j�H.��D<=�J̽<1H�?����k�%�)�����A�?�[�>�6?�ڌ�r���>���>�Ǎ>�J��c���Tȍ��gᾒ�?>��?a� >ͯ�>�B?v�>uq/�CFҾJ_�Sǂ�x7��e�`�U�����Y�Ց=��ί�0M?��?�8W?��>���>���?��;�����C��>�#���,�"��=�I?Y"�4JF��n��t��������>9��?���?G�?�'\������2>�]H?��O?k�q?g|,?j?$=�;�D�>�{=ԃ:?0Q?%?�?E>e>��=��ȽE�=�߽�w~���H�1�9������_;<��=/gS<��<��-=Z�=b��x��ˀc�����=�4�=��={U>|��>��F?�?, �>Qd&?��"�,8���� �?w{�=T�پr�Q�����f�X�>��]?�V�??�m?V>��H��DG��| >�5s>B3J>�tI>У�>6�Խ*T�*"M=YZ�=�rC>�zI=;̽����P��L���	p=-�*>��>��C>�ȼi�>P���FԾ��r=�]���	"�K���ye���;�ƂU��g�>Wy?y??�_�=^]��+��=��H�7��>�%�?y�?wd?G��=�|~���%�3U�T�>������>��3��Դ�0���o6�u�<�F?�o���ޠ��Wb>��<t޾h�n��J�D���GM=���]V=}�U�վ6�o��=/$
>���� �"���֪��1J?=�j=�w�� bU��p����>ѿ�>�߮>�:���v�i�@������5�=��>��:>�_������~G�J8�~6�>^WE?#T_?n�?"*��?s��B�6���1c���Eȼz�?w�>�^?��A>ѭ=$���i
���d�`G���>��>�����G�5���)���$���>H=?�>�?)�R?Z�
?��`?j*?�D?�%�>���b��oA&?���?���=Y�Խ	�T�B9�{F����>��)?��B�c��>O�?h�?M�&?]�Q?^�?��>v� ��A@�J��>�Z�>��W��b����_>ڪJ?��>�>Y?'ԃ?�=>ڃ5��詽�S�=�>j�2?�6#?��?d��>}��>M���~�=���>�c?�0�? �o?���==�?�:2>R��> ��=���>X��>�?UXO?A�s?��J?��>G��<�7���8��.Ds���O��ɂ;iuH<��y=���Q3t��J����<�;�g���I������D�����\��;q��>%�>9� �>Aﾙ����a>��{�b�߾�`������gh>֎�>R?���>��ڽ́>�v�>��>9����$?��?$k�>\+���}E�J|�����>77?�a,�.숿F���o��^�>P�?H�3?��g���Z���b?��]?c��?=���þ�xb����P?߱
?�NG�F�>B�~?�q?b��>�8f��<n�\���Sb�j�i�X,�=���>�
�{�d��؝>�P7?so�>�b>���=��ھ�w�V(��$�?"Ԍ?��?C��?�)>��n�`'�� ��F����m?;v�>��ξ�{?�+��s˾�F��)^�� ��y�����O���,��V�b�J��*���y�=394?Cԃ?�No?�zJ?�� �?q�&�e�l���}>�z�,���9X���/�O�-�ܧ9��¾T���n='��'�=Nـ���B� �?��"?��B��>y���H��"A̾��B>b��o)�p��=�b����S=+��='�Z��~'��g����#?i��>���>�[;?m�\��A�y3�+<�B�����>�@�>�>>��>���;AK��ٺ���¾q�u�x��'�u>״c?GbK?i o?<���1�K��[�!���5�W.����B>�>�	�>�cY�a��us&��u>��
s�i������ۺ	�O+=��2?��>�ۜ>l�?�?w%	�x���%iw��1���<��>��h?���>=�>,н�� ��>�p?�_�>�!�>�����'u��j�2ݿ>���>�k�>Z�q>/�9�ڻ_��'��U����:�
��=��f?�ԇ�2�Z�D��>*W?�~�:P��<�z�>}	����r8�����)]�=Cc?��=!Y5>�Ǿ.��`w��$�� O)?�G?�ڒ��*��6~>�"?r�>I0�>1/�?�'�>�yþ2�D�8�?D�^?�?J?UA?�R�>��=���5Ƚ��&���,=|��>��Z>Im=ʊ�=P��
l\�m�,E=gl�=g�μ�_��Ql<*a����K<J��<��3>[Lۿ�K��ؾ1&�70�t
��׈��W��w�������������x�y����&��U�o�b�����7l����?��?�����D���ؚ���������Q��>��p�؀��b��G(����8L�0��S� ��pO��h�9Ke�?�'?������ǿ簡�L:ܾ�  ?%A ?q�y?�П"���8� � >�P�<���כ뾙�����οS�����^?���>;�82��E��>[��>֢X>Hq>��^螾$>�<g�?��-?/��>h�r�>�ɿo���Ť<���?��@�9?J3D�:���L�=	�?%>���(0�����`ž�=p��?"]�?��
?>o�)��0n?�1�>�<���59��>U>_>ʀ>tl��m�=���>��9�}!���! �}.>�ة>*��H(�2� ��A=p��>��`��N�5Մ?+{\��f���/��T��U>��T?�*�>N:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=c6�鉤�z���&V�x��=Z��>b�>Â,������O��I��S��=��\�ƿ��$�d}�h=�׺.�[��f罷˪��T�'��ho���轐sh=ƕ�=7�Q>f�>|W>�0Z>yoW?��k?q[�>�a>���򆉾�ξ�|��<��G��0�������飾+G�{�߾\y	�������u�ɾ!=�u�=7R�k���7� �c�b�U�F���.?w$>P�ʾ��M���-<npʾJ���z܄�᥽�-̾�1�"n�i͟?��A?������V�W���W�����R�W?	P�ʻ��ꬾ%��=F����=�$�>��=���� 3��~S��w0?�R?Z����c���*>�� ��]=�+?�y?��Y<�(�>3O%?S�*����I[>L3>���>Y��>�N	>�����ڽ)�?	�T?�����y�>8g��{�b=2�> 5����-x[>�G�<�֌���W��ѐ�Iݻ<Zk^?}��=؃@�/
P��2���	?�d�>$vu?�a?+1�=��?2�/?V���a ��W������P?>r�t?;�z?�N�=	�3�\�ξg�z�^?64?c��=D�C�☴��D�T��\?��x?,NP?����o��ﱿ�.�]?��v?�!^��W��~���-U��Z�>���>N�>͵8�I۳>��??�0#�m/���꿿�4�l��?Z�@Ջ�?ȳK< �!����=�?t;�>.%O�
g¾�볽�ʵ�4q=I��>3å�x_t��C�+��6?]��?\��>'H�������=�ٕ��Z�?�?߅��^,g<r��l��n��=y�<ʫ=h�KI"������7���ƾ�
�3���5׿��>EZ@!X�g*�>�C8�V6��SϿJ��\о�Vq�h�?��>�Ƚ������j��Ou��G�f�H�ɤ��U��><:>�>�����ψ�J"=��4�=7�>����B�>U���־�x����l����>&?x#�>!ǽ�������?s9�-ҿwã���,�Ȫ}?��?���?��P?Vz�>3V�=�|��	�:7�>\Y?v�<?.7V�q����(�<��k?��t���i���8��0��rq>�B?�w&?�{�=xb�>���>;�=��ϱ�/���$�"��Ev?l��?jվ֨?oԛ?�*?k �yg���w�����EB�Y[?�(�_a����&1�6S�?�?3�?$�Ӿg�(�c�A?�V=�[W6���0�qK6��9U=.���D����$��tܾC�[�Al��D�G?�?$\@���?'�)�v��.?�R�>b:��-��g�S�IF?�Un>��I=+�޼!��=B�3��^���e>�P�?2; @�?����tि�PN>�h?��>���?.�=�)�>� ��'�����R>LK�>N�ν��>~u�>ψB?�_g>�ɣ�X���ۓ.��g��o�x����P�J��>��T?�>y?�=>Qt	�K�2�b�\�)�S���Y����I�ѽ2��B�����=/��=��0>�y���c���?Np�8�ؿ�i��p'��54?%��>�?����t�c���;_?Xz�>�6��+���%���B�`��?�G�?=�?��׾�R̼�>=�>�I�>@�Խy���Q�����7>-�B?J��D��t�o�l�>���?	�@�ծ?oi��	?���P��Wa~����7���=��7?�0�/�z>���>��=�nv�޻��T�s����>�B�?�{�?��> �l?��o�P�B���1=@M�>ќk?�s?�Ro���[�B>��? ������L��f?
�
@u@f�^?(�
ʿ����l�6�՛e>M>��=-@����=���=�D�=�t%�6�=��p>�
:>��k>���=6�A=���=ġw����g�������*x�ς$�3�����C�L��H �7+� ����C��u�_aA�'f�nae�vg��U�=W�U?R?�p?�{ ?%y��>á���=D�#��ڄ=�,�>G2?!�L?v�*?3��=\�����d�`��s:��N������>�`I>ŀ�>&0�>��>���9��I>9 ?>S��>�� >�'=�%ź[}=�O><I�>��>qC�>�C<>��>Eϴ��1��m�h��
w�O̽1�?y���M�J��1���9��צ���h�=Ib.?|>���?пe����2H?(���})���+���>�0?�cW?(�>��h�T�C:>7����j�+`>�+ �{l���)��%Q>vl?�Eh>E�v>fC3�(`8�x�P��T���>h7?�5���5�r'u�P�G�xrݾ��K>���>t�Z���
"��ܢ}�)�k�5��=�:?|�?_I���ֱ���u������cO>_]>A�=d�=U�J>�ml���Ž��E�ϐ-=��=��Y>9l?�{,>r[�=M�>����P���>0�D>�*>�@?Q�$?���8g��6S���0.���u>�1�>�>ː>a�J��Ѳ=��>�Sb>d�
�2L��V��&�@��V>Kw�'a��Oq��s=zz��8�=W�=� �rt=���=�j?0z��|�{�3o��K�<���><A#>�;��>��A�s!��)����9�?H	@��?�m��>�ǫ:?f�?v�"=�;���}>:q�>(RO���S��A�>��=MO�v��T����?�R�?���pq���;N�|Ym>أ(?���Rh�>x��Z�������u�|�#=N��>�8H?�V����O�c>��v
?�?�^�ߩ����ȿ4|v����>W�?���?g�m��A���@����>9��?�gY?yoi>�g۾2`Z����>һ@?�R?�>�9��'���?�޶?ԯ�?��/>H�?l[k?���>��ν�#'���������<#O��ݟ�>/h>K̾Y�L�0㐿"����-l��#�
d>��<��>R���j����=��`�W����3�I��>N�L>7�A>8�>�T�>�g�>��>3�J=3Z�`<~�uO����K?���?+���2n�0N�<H��=�^��&?�I4?qi[�{�Ͼ�ը>ߺ\?h?�[?
d�>B��Q>��A迿>~����<��K>/4�>�H�>%���FK>��Ծ�4D�cp�>�ϗ>����?ھ�,��BS��HB�>�e!?���>pҮ=ۙ ?��#?��j>�(�>BaE��9��U�E�Ĳ�>آ�>�H?�~?��?�Թ��Z3�����桿��[�p;N>��x?V?uʕ>`�����kE�`BI�8���]��?�tg?cS�-?;2�?�??_�A?{)f>ׇ�*ؾ������>?�!?r�a�A�QN&�	��}?�Q?���>17����սּ����~����?�%\?y=&?c���+a�|�¾&�<W5"��LS����;q�D�޶>��>/����{�=�>1��=@Lm��I6��f<l�=���>|��=�:7�_����=,?(�G�]݃��٘=��r�LtD���>+LL>* ��Q�^?�`=�	�{�i��6y���	U�l�?{��?�k�? ��[�h��#=?��?9?!�>�D��-}޾p��[Ow��x��u���>d��>��l���{���z���$E����ŽD��H�?J��>��$?���>(~3>yѷ>e����q0���ᾲh��ԶM�����F�q�3���'��ϻ�|vn��j;�8þۑm��ߕ>)�*:��>P%
?��M>׿Y>�L�>#d ��1�><(>pv|>.|�>�fY>,7#>f
>$B�N;ֽ�WR?�T(� b�s��b@?� c?Ay�>�+h�ϲ�����[9?{��?�p�?2qm>?'i�}�*�8?>Z ?��}�L�
?A\=���:-<����=��0x��C\/�_�>�����69��MM�bi�,
?�x?�*����о޲׽����0o="M�?l�(?��)���Q���o���W�rS�M���5h� g����$�T�p��쏿�^��3%����(��*=φ*?��?�������#k�p?�/Yf>��>��>!�>�lI>��	�N�1�4^�9M'������P�>Z{?Ӈ�>��I?�
<?�rP?�dL?ԥ�>�Q�>�+���V�>2��;>�>z��>2�9?�-?P;0?X�?`{+?�3c>�y������ؾ�
?��?~D?�?˰?5م�`iý?i��Ff�)�y�g����ہ=��<_�׽vQu�~U=,�S>��"?���s�M����+^>�7F?�N�>��?e^$�����
)8>ӵ�>�_�>Q�>1e��'~�����>��?��Ӽ��=��>�>�<=� X'��o=Dߘ<YK
=A(L=����9�ˈ�=a�
>i��<�m����������>�<u�>��?^��>�B�>�@��� �ߵ�,e�=�Y>�S>�>�Fپ�}��L$���g��cy>�w�?�z�?��f=F�=���=?}��fU��Q�����'�<,�?:J#?�WT?W��?��=?�i#?#�>+��L���^��o����?Y�+?ɷ�>�7�\�ʾ9����23�W�?E?�0a��	��(�翾�ڽW�
>�"/��}�]��~E�R��M���k��v�?��??@�f�6��9�;C�������?B?̨�>���>�#�>X�*�6�f�|��;>���>8�O?$}�>�N?@�z?d�[?��P>��8�)�������R�����>��>?V�?��?�>y?�M�>7>��%��o޾����p� ����
���ZCe=�V>�͑>�R�>8�>|�=5�½	ν�W�B�K,�=�3^>U[�>n��>(��>��w>_��<��V?�͇>�4޾޵;��?ɾ-�:Y��>ý�?i�?�r?���>d!��S\�sQ$��r�>:�?�y�?��?�_콅k>���dW�?/��Gc"?��9?��=�{Y=�?j:{���8?~��>f�ý�bA���K�
Cm��(G?Ͻ�?��=Y�ۿ��G��g��� ��\?��-=�2V��3��yؽq�>=�ֽh�w~̾m��|ﭾ�h���v��ads��I���>#��=F��>'� =��!>m״=/�>��=��=��=�a$���=����0�\�x�N��)�w��=R>9��=B�־�]�?=�A?�j?�m�>]�=�pT>��Y�la�>`�a���>�s>�E��խ�����پ� �C=�R��sc�b<,�Yk>��+`>=��=��<v|�=��w>,���Ps>��V��=���>_�9>��h>w��=EC>Tٽ�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>֭7>#>d�R���1�*�\��b�f~Z�(�!?KI;�J̾�5�>A�=<,߾͒ƾ��.=��6>zpb=Yg�+V\��=�z�w�;=�l=�׉>1�C>�w�=0����=�I=��=��O>�A��U�7�5,���3=U��=�b>&>���>U�?g�A?`�[?�ϓ>K����޾��Ǿ(�>Q�=��)>��<x�!>�z�>ޡG?]�R?e�R?�^�> X�=?��>�Ʋ>���.r�V����᜾Y%U;�:�?jz?N�>d^<).���X2���4���Y��2?ہ-?[<�>���>KT�e�࿝m&�iy.������:j�*="r��T��������9�=�-�>���>n��>��x>x�9>�tN>���>��>�A�<O��=�5��1w�<���"��=뒐����<EPļl�e+��+����9��;�΋;�__<��;���=k�>yZ>�>"ʓ=+9��A(0>ᖾ�M�8U�=�;��mxA�p1d�z~��/��7��?>�zU>�+���*����?s�Y>�	D>|F�?��t?�>zP���վwE��e�c�G2T�Tq�=u�>�=���;���_�F]M�@�Ѿ��>U��>o��>�q>Λ,��Z>��G�=ō޾VK8���>x>���.��	� ��^r����Oɞ��Hk����`�A?�c��Vq�=K4z?�R?�v�?I��>�ý���C�>>6���=
����t�$�ҽ�?�?���>��?�@��H̾�� �>BI�S�O�Q�$�0�2��&ͷ�3��>�����оD$3�kg������K�B��Kr���>�O?��?p6b�CW���TO�X��1.���p?u{g?��> J?!@?�+��my�r���{�=G�n?���?,=�?�>��=����:�>�+	?u��?ظ�?Ƀs?z?��z�>��;� >��II�=V�>��=�*�=�s?a�
?��
?i����	������D^����<�Ρ=Ʉ�> m�>b�r>���=�g=/x�=v/\>�ٞ>�>R�d>J�>YP�>�����%�^�&?�t=Y�>��'??W>m��=��:�h�=%����+0�JCH�[m��>2���<�!������Ɯ ?�qϿ�ȏ?��X<�UD�C��>a�Ծ!_��F[>��v>�������>�5'>���>��> ,�>6�S>��r>y�y>�FӾ`>����d!��,C�]�R���Ѿ_}z>Ȝ���	&����w��@BI�jn��hg��j�O.��Q<=�t̽<+H�?�����k��)�����U�?�[�>�6?�ڌ�p���>���>�Ǎ>�J��l���]ȍ��gᾤ�??��?�O>�ǈ>J�p?˙?݂��VP��]9[��rn�#SE�ĄS��t�����j���Ѿw��=�q?��y?%�*?7ˑ=)��>_�?���]^����>s5���:�q��=V��>>ƺ�Z��t�2̾���M-�>Ul?bp??���1�m��'>��:?1?�Ot?��1?[�;?i����$?�o3>�F?�q?N5?��.?�
?A2>�	�=����'=�6���ݩѽ�~ʽ����3=�^{=��̸} <��=Q��<��)�ټ�;�%���$�<
:=d�=8�=��>>S?�2?;�z>8�&?��~��<�����%?� :=h���w���>���ľ�	T>:�v?i�?|�O?9#P>�����;�;�.>�7�>��=�Q>��>�	��!�&���%>V5>�e�=ȻA=���oE��c��2A���0�=,�=�s�>��>�E����%>�k)��Z�n>P�J��N��UnC�Y�F�8�,�2~�>�/G??�?�b=�Yﾗ����Cg��^*?�5;?FRR?G*~?)*�=}��7�?��J�wM&�B��>��<`"	�ag��������:���<�2x>�/��!٠�KUb>M��x޾y�n�MJ����I{M=+z�$9V=|���վ6����=�"
>w���:� �����֪��.J?�j=mq���XU��u���>���>�>�:���v�-�@�r���k8�=y��>�	;>������}G��;��E�>w�E?�o_?ox�?������r��A�O��������׼�?�>k�?�@>��=-���#��Ee��G����>m��>P��3IH��T��A����%���>�?�> �?z\R?p�
? �_?Ş)?J?iĐ>�
��Eѹ��A&?4��?<�=l�ԽJ�T�� 9�CF�l��>o�)?��B����>I�?ѽ?��&?�Q?��?��>� ��C@�˔�>yY�>��W��b��*�_>��J?>x=Y?�ԃ?��=>J�5�ꢾ�֩��U�=~>��2?�5#?L�?ﯸ>��>C���%�=���>1cc?c�?�o?���=�;?9�3>���>j��=�֞>o��>�?.>O?+(s?�mJ?NK�>)ے<�*��S��Rw��c>���y;|�B<�-t=�E�e�q��A���<?s�;",���Mn�yw�(,D�U#�� w�;P��>�j�=W����}�>{�������?�=�I����̾�����̾hYz>��>�,?���>n��<�S>8�?���>�)��5?��7?�&�>�^��^,��=j�*`g����>e0`?���>쁿\eʿ~��]��>�s�?{?�#�@ �̺m?Z%1?L~��e�+��=���8��(e?G�?�g���߅> �o?o�=?E�>
���kw��ܛ�*^�ZX.�ӿ =�Q�>=NѾ���Ziͻ�a>?<:?�@k>og�>�+㾛r�ߥξ(��>]�?J�?.?@>�>�Rr�"���d�����<Mr?�ϴ>>���5�3?����柾��վ��ǽ>�����/���쳎��$��56�M�D��v��p>d9G?��?/�T?c�L?SJ?�"�v��I��<��"_�v����1�\�RY1���@���6��ֈ��葾3���>і���mB�0��?��&?ԗ0��}�>�������r�Ͼ`�G>�����4E�=<��ӟ6=�Xe=��d��~.�~���N�!?z�>���>�b<?I\]��@��{1�x�9��J����->��>�؍>���>D�����&��$ӽ<�žai��߇˽J�u>�c?��K?��n?)��#1�9h����!�z�/�Dj��'�B>h�>��>��W�=��z1&��[>�s���ԃ���	�1M�=�2?�>�>fÜ>c9�?��?Wo	��P����w�$e1���<E2�>�i?��>���>�ν%� ����>ܰl?�g�>���>�k���H!�Z�{�g�ɽ5�>1ح>��>�?p>��,�L*\�@l�������(9��F�=b�h?�~����`�U݅>�R?>}r:��F<ԉ�>�v�O�!����(�ڕ>Uw?i�=	z;>�rž�2���{��U�� P)?�D?钾��*��A~>�'"?�v�>*�>/3�?'.�>Nsþ:}9�յ?i�^?�:J?�OA?BD�>��=���<Ƚr�&�G�,=g��>��Z>�m=�v�=[��{j\�_w���D=*��=~�μ+W���<e]��z�K<���<r�3>mۿ:CK���پ�
���>
�\舾
����d�����qb��`���Xx���R'��V�}6c�$���P�l�ׇ�?�=�?�����/��W���N����������>5�q�����������N)�����r���Qc!��O��%i���e���'?ް��q�ǿ����v7ܾO ?�3 ?��y?,��"�(�8��� >��<Pg���w뾇�����ο�����^?���>�`.�����>أ�>��X>UTq>���՞�}ӕ<�?��-?3��>I`r�&�ɿ�������<���??�@K?�yE�������=�$	?KW�>�ǖ���I��Ӿ����F>^&�?�G�?�b�>�F_�&V¾Q�>?H&�>�"�t �Չ^>��>o�L>����E4�;	�>yщ�5���Ɨ�9٦>�6�>�M���L��Xx�i���F>n�,>W>�5Մ?,{\��f���/��T��U>��T?�*�>U:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=v6����z���&V�{��=Z��>b�>,������O��I��S��=����ƿ��$�Bi���=��$�[��N罦S����U������o���h=�>�=}Q>T[�>�'W>'Z>�WW?�k?�p�>r>���Tf����;���kf��ّ�������A����W��߾�u	����y��4�ɾ� =���=7R�s���>� ��b��F���.?�w$>��ʾ��M���-<�pʾH���@܄�p᥽�-̾�1�/"n�R͟?��A?������V�z���V�Ѓ��J�W?*O�����ꬾ���=����r�=J%�>狢=C��� 3��~S�y0?VR?Ǝ���c��T�)>� �aJ=��+?�?X)X<��>R%?p�*����&T[>�h3>�£>��>��>"��F�ڽG�?��T?E�E���ސ>�{����z��b=.>�N5��3�L�[>%Ò<Oˌ��dV�3���g1�<��n?+�2>��U�z�w���ƽ�`>��H>'�}?�T�>"��>�l�?��`?�b��(6�P{d�y����>��T?�L}?��=���������skL?�6?����I*��몾��G�'�!��8?�yP?#??�5��b�������$�?�N?��v?�r^�xs�����S�V�n=�>\�>���>��9��k�>&�>?�#��G�����~Y4�Þ?��@��?f�;<��\��=�;?F\�>e�O��>ƾ�{������o�q=z"�>Ռ��Jev����R,�I�8?ɠ�?���>�������Q��=�㕾m[�?O�?ψ����g<h���l�|���B�<ُ�=�j��}"�����7�N�ƾ/�
�����P��ܴ�>/[@���,�>�n8�59�PQϿ����aоtq���?�b�>�Ƚ񞣾[�j��<u�	�G�u�H�a������>�f'>#��;lS\��󍿐w7�Ll�=y��>��G�f��>��p�"ϾmP�еK���>��(?���>&�$�4�ʾ�O�?B��tԿ���g� �ǡ8?���?)$�?��.?"�?>%�	<C��,|�=�#
?
�[?��3?Ǖ����2e,=G�j?Y%��X�`�Sc5��4D�QU>��2?B�>w@-�'i|=Ld>��>��>�d/��zĿ��������?t��?.���_�>)�?{�+?�l� ۙ�����zq*�y0:ek@?��.>E����6!��<�ԯ����
?�X/?f�
����w�<?O�n�x��'+�\�����@߾0�����о�&w��۞�|����?�d	@ǘ�?j�������N?	��>�鎾�w�����(��>*M ?��>�P����>��ؾ�n0�a	g>���?t�@��?Lƪ��T���ܿ>rn�?��>+ҍ?��>�
?�y��ھP�=��@=���=�x��s�>�9?6t�>���;�e��?� �=��������HB��>�U?�X?�Qm>r�i�3����B�[�p�������=b�ǽ�������_\�==��=��:=�@�d'�� �?cp�)�ؿ�i��jo'��54?ɸ�>��?�����t�w���;_?�z�>�6��+���%���B�U��?�G�?,�?|�׾^O̼�>�>�I�>�Խ��������7>�B?o��D��h�o�9�>���? �@�ծ?�i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?oQo���i�B>��?"������L��f?�
@u@a�^?*�(ڿ\Қ��:����ii�=�T>b�>Rk��'7��k�8�.D=U�Q��=LR>�=2>(,y><��>P�=>���=����D��.��[���X�J�u���	�I-ӽa��2Ǿ����O������ea�8��*���[gG�J�W��Ք��I�=#IX?��Q?*Dq?�R�>���6E&>�w ��,=��'����=��>^�-?4�G?�c'?�Q�=:��<`h�;퀿=������c4�>3M>�b�>���>(_�>U#z�D>��=>"�>0��=�f!=dU;==WbI>:�>��>�-�>;H<>��>ϴ��1���h�: w�Q̽`�?%{����J�v1���7������Ti�=Va.?�x>����>пM���	1H?@���'�c�+�J�>8�0?YcW?k�>.
��C�T��5>���Y�j��d>�# �/xl���)�,#Q>�h?���>�+v>��2��>�AS�4OZ�\��>�D?[�'�p�9�ҕp�i�4��~ԾB]M>�h�>]���"���T��/���UÃ��F>�E?��?��$�ۢ��>s��f���\b>�J�>w@�<\=��Q>S�#�}X����ͣ=�Cp=�_>�W?��+>㦎=�ڣ>"n��^AP�-��>c�B>�7,>�@?�#%?~c��ܗ�̂����-��w>~L�>L��>�<>6fJ���=�q�>f�a>-w�7܃�����?��dW>t�}��s_�?qu�?�x=OB����==/�=Ç �m=��%=��r?wՖ�xK��0ђ��(>��.?˱F��ϸ���?>[D�Z������)��?=
@�)q?~m)�&I� �;?��?���=�KZ����>G��>j���	�=�>���<ђ�=}:�з�����?
�?��H��Ԟ��&�I�#>�3�>���hh�>zx��Z�������u�̷#=R��>�8H?�V����O�M>�w
?�?�^�੤���ȿ>|v����>X�?���?X�m��A���@�q��>/��?�gY?foi>�g۾Y`Z����>��@?�R?(�>�9�f�'�r�?�޶?¯�?��H>뒑?Οs?K��>f�x�L_/�,"��~����\=?hK;�z�>�>�����_F��ʓ��`����j�!��݄a>x�#=��>�H�A\���=򈌽�d��(�e�H��>�q>��I>�L�>�� ?�9�>���>f
=�^�������Ӗ�
EL?zߊ?���<4m��Mt�g>��׽W�?�U?�%�<�9ؾ�ۨ>S�L?��s?�V?Kя>Sv��9���*¿عžܛ�=�ي>
 ?b��>1�,�8�>*-�7�n�i��>P��>�5�	sƾ5���z���r�>��?���>�J�=ܙ ?��#?��j>�(�>@aE��9��V�E�ò�>ע�>�H?�~?��?�Թ��Z3�����桿��[�r;N>��x?V?rʕ>a�����kE�<BI�.���]��?�tg?yS�-?:2�?�??a�A?x)f>ׇ�,ؾ������>y"?���g�A�`�&�5,��N	?g?)Y�>����GڽOI�O2�1��F�?n�[?F�%?����4a�'4ľ=�<����YI�79l#<"V��-k>qt>�X���s�=DJ>@�=�Vm��65�ǻ�<#��=���>��=Z]7�f���,=,?�G�Eۃ��=��r�3xD���>�IL>(����^?�l=���{�����x��rU��?��?Ok�?���2�h��$=?�?/	?d"�>�J���}޾���Pw�6~x�ew�K�>���>§l���;��������F����Ž�e��>���>�!?)w ?��O>`d�>�$���'��n�����^��l��k8��.�����頾Ff#�F��2¾�{�u@�>*�����>ڞ
?7�g>��{>1�>ʻ2G�>��Q>�s>'Y�>��W>"5>?�>�!<yXн�S?����c(���޾z��bF7?Z?��>���I����� ��'?��?�җ?>P>��d���%��?b=�>�����?m9�=&U�=����U.��<��EY轨ķ<�U�>{�@�5�XCH�+Q�B?Vl?J#��̾�	�/���h o= N�? �(?�)���Q�M�o�ƸW��S����5h��i��C�$��p��쏿�^��%����(��p*=��*?]�?Ì�h��D!���&k��?��df>P�>/$�> �>uI>��	�o�1�D^��L'�2���}R�>)[{?���>[�I?:<?4xP?�kL?O��>�c�>4���l�>��;Q�>u�>�9?X�-?	80?�z?�t+?3c>��������ؾ�
?��?�J?�?
�?rޅ�.tý�h���g���y��~����='�<�׽�Fu���T=�
T>�&?ݲ�ןC�;3��&�>s�2?fB�>">�>�����Y�[�=���>x�?�8>���=4�����n3�>�I�?}����=h�+>O�>��I��t��_�>�;W�:��=!mq�g��"�X�Vi�=�`>����T��`)��o�3Ŧ�4^�>��?���>���>�چ�J� �Y��Yծ=�wX>��S>�>�پe��������g�V{>C��?�X�?=cc=���=w��=��$���c���ͽ�C�<�?�k#?XmT?>��?�h=?0R#?�>�*�����O��|ˢ�6�? ,?W��>����ʾ�񨿀�3��?"\?*a�K��e8)��¾��Խ��>xU/��%~�"���D�=n�����A0�����?�?r6A�'�6�{�辴Ø�fw����C?�'�>VP�>g�>E�)�3�g��!��);>Rj�>�
R?$�>y�O?�;{?��[?~gT>z�8�,1��mә��[3���!>h@?#��?�?5y?�r�>�>��)��+T�������߂�W=�Z>萒>,)�>��>���=�Ƚ�V��1�>��\�=��b>Ï�>$��>��>��w>lG�<�W?u��>�	ݾ�B1�����=�����x>���?ZP�?k�u?�5>� %��^E��l��O�>�?�?�ַ?SZ'?��F�9�Q>��I��	�����$?�M�>�ǒ>�u>G/��іa=�)?�?��V<��4��M�� ��[�?rXT?Q!^>]Eƿܡq���m�t���`��<l����!e�*����;[�r�=���7/�$�����[����o��kZ��6���(�{�+��>��h=,��=U�=69�<��J[�<�qS=΁\<��=�P�����<f1��<����NL��PP<��A=_{�j
��;x?��Y?�w#?J�?y
h=���>T���p]>�3��<?��
����r羋�>�WT���	�k��I���+�o�|�x�=Ga�D��>��3>`L�<��x>S�>]M�=v}=����D<05=q�}=�ç=�/>�Z�>\R(>�6w?W�������4Q��Z罡�:?�8�>S{�=��ƾn@?y�>>�2������yb��-?���?�T�?=�?:ti��d�>F���㎽�q�=B����=2>Z��=|�2�S��>��J>���K��6����4�?��@��??�ዿϢϿ9a/>�7>Y$>d�R�8�1��\���b��zZ�^�!?ZH;��I̾�8�>7�=�+߾ϓƾ��.=�6>�`b=i�V\���=3�z�k�;=k
l=�׉>�C>sv�=q6����=N�I=���=��O>, ��z�7�H',���3=���=~�b>�&>6��>�?ra9?�Ad?Bƀ>qw� ǾB�Ͼ2�e>��>�>�g=]��=�l�>np0?�V?(c?��>��t<���>��>c�2���l�B㾲l��%��=j�?��?C!�>zӤ=(ef��6��<�Tf�x�?�I'?�[?y:�>)���F�,;�D�ô���.���T�<������M�c�� ���@�:Q=�Su>Ԃ�>�z�>T8q>�$>��>�͝>�>/��=���=�x�=�~���¶;j'�-_�Lo>�~d���༞�#�Cd)�n�T��μ{ڙ�Oc�<�=<��=n��>�<>���>�w�=�
��;H/>U�����L��Ŀ=jF���*B�d3d�WH~��/��U6�p�B>�(X>n���4����?��Y>�v?>(��?#>u?S�>�0�0�վ�Q���:e��RS�Yø=ԭ>!=��z;�Z`��M��xҾv�>��>��>�^n>V�+��L?���t=Ɋ�Jv5� 9�>ti��MK�&����p��#���ǟ��h��\a:o{D?�$����=�h~?��I?�[�?[�>����ːپ��0>/Ӏ�~ =�@�z,t��AS?��'?xu�>���aUD��H̾G�� �>?I���O�����4�0�,��з�ʑ�>����#�о=$3�Eg��d����B��Hr�`�>�O?��?�*b��W���SO�T���B��p?�xg?4�>vH?$@?M9��Cy�ts��Ђ�=�n?o��?�<�?�>A*�=ኴ�[{�>j�?'Ė?/��?FVs?�J=�	��>���;��!>cߚ����=��
>+��=���=b.?:d
?X�
?'����	�������#]�d��<��=CO�>�'�>A�r>�6�=m=�C�=ZO\>F�>J#�>ƹd>��>�4�>_=��	���A)?G�=��>Ϫ;?��$>��=q��ח=�j�g�6��*G�9#��V��v����Ke����',%���?6̿�C�?
��=_���?S�O��2�=�c�>�����<�>�OH>#܎>���>܀�>�L>��O>GC�>�FӾC>����d!��,C�N�R���Ѿ�}z>�����	&����w��ZBI�tn��pg��j�L.��T<=��˽</H�?����k��)�	���Y�?�[�>�6?�ڌ�g����>���>�Ǎ>�J��g���Yȍ�hᾠ�?B��?��0>�i�>S�f?9�?[�۾_k��K�R��o|���d�_&�r�r�&'��u�� ����">�)�?�j�?l#?��:B�>�Б?�6K��;��
�A>�+A���8�7,���~>�4 �)�i��:��⻾߬f���7>$|m?�r?���>�]���9����=uM7?��>�?��?�0?���=9�+?9��>�/?֐�>�S?X� ?
K?/t�>Ԯ�=�;�P�=Y����!ؽ�9��LE<@N�<�*0=�Iս�,7���_=��=�P)>�G�;�/�=8[=cb�=��`=��=�%�<7��>ț]?ݘ�>Vǆ>	t7?.(�Wh8�����F�.?:;=L������+�����4>�k?O�?KZ?r�c>��A�x�B���>��>�O&>�\>C~�>��p)E�d=�=�>X�>#�=��N��L����	�)B���D�<u�>���>���>yg@�l�>)	۾_=z��9�>L�뽳�9�6����=�L�sn�T��>�>?-(?>�]=ϥ���O��l�fF9?�B=?I_j?��_?�1���]��cp��P%��4�>����¡��؞�X|��Pb-�ѭX<L<=e]��䠾Rb>����p޾��n��
J����.M=-~��jV=\���վ�;����=�
>����6� �L��7֪��1J?��j=`t���^U�on��8�>-��>�>ӹ:���v���@������,�=��>�;>z��~ ﾦ}G��7����>�C?|�^?�f�?�kz�Js��&A��Z ����1���K?E�>��	??H>(R�=r����e�y%b��E����>\V�>���iAG��e���T����"����>�r?|�>�?�IQ?(=?_�_?u�(?�?��>jݝ�Â���A&?<��?��=c�Խ��T���8�+F����>��)?ϸB�y��>��?ܽ?J�&?��Q?5�?��>� ��B@����>gY�>b�W�Jb����_>-�J?���>�=Y?�ԃ?m�=>�5�颾�ҩ��S�=�>�2?�5#?�?P��>RQ�>O�����=A��>�c?(@�?_�o?H�=��?��1>��>�6�=� �>��>��?O?ls?�J?��>t�<X<�����S�q�oD�eD�;y\G<qXw=�+�^�s�j��Ev�<� �;���S+��c����D�	L����<%��>�Xt>e]����/>�ľW���t%@>A㟼�f����$�:��!�=:��>�?Ӈ�>�>"��|�=S�>K��>�����'?s�?�)?�/�:�b�}zھ�2L�E&�>|B?��=��l��k����u���c=־m?�Q^?��V�y��f�f?y�P?C����?�f&Ӿ^�B�0?���CV?��?5�W�Ae�>���?��{?mL?��v���w������W�w�)� ��=���>gw���b���>�SH?���>�V>��>ɐ��ϳ�A���+?34�?a��?(#�?��
>�wp�g��ծ��?��MW?�Ƨ>g���&#?�񽃇۾(E���r\����_�����2䮾������l��7����g��>.2?�U?P.V?��/?D�+���j�D�B�.�@q��%�o� ��b���E���E��KG������Ҿ����C;>j}���A�c�?��'?��.��V�>�����𾎮;KkC>����B�;�=�_���<=%W=�h���,��୾�  ?q�>{*�>�<?Ѳ[��>��)1���7�BA��x�2>hˡ>�u�>66�>�h�:�F.��U�)	ɾ�����н�v>sc?��K?��n?��w	1��}��	�!�\�/�e��3�B>[�>pω>�iW�/��2&��a>�A�r�L��ln����	�h�~=;�2?�$�>k��>J�?)?��	��S���"x���1�nC�<��>�	i?
C�>�>�tϽ�� �V��>��l?��>��>陌��Y!���{� �ʽ�$�>s�>C��>2�o>��,�� \��i��~����9��Z�=��h?����G�`�E�>]R?X��:S�G<�q�>�v���!�r���'�#�>�|?|��=�;>S�žN'�8�{��:����,?�?&�˾��9���`>�<?���>:}�>3Px?(�">YZ��M`۽U�?�$i?�}?�N??��>���&�=Qg����)�t=C�>�!�>U��s�T�g"�=�����5�}v=_	>��==�:���e=�~����
=������{>�tۿ�RK�?�پ�����
��s��n紽�!�����h���S��6�y�/	�g-���V���a����� m�U]�?:&�?Qm��:5��d��"k��G������>G,q��y����l4�¯���䞬���!��O�Ki���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >`C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾}1�<��?7�-?��>Ŏr�1�ɿc����¤<���?0�@:A?��(����]�U=���>·	?r�?>�1�/E��᰾�5�>:9�?���?�"M=9�W�W�	��{e?̀<��F�.��)�=yc�=:�=��luJ>�A�>[l�4qA���۽S�4>�݅>8�"�����^�Y�<��]>�iս���r�?��X��Uf�BD0��~��3>	�Q?�o�>I�=Yl)?�bG��Ͽ�Z�n�a?���?�_�?T>(?�¾`��>�]۾��J?a6?ւ�>?V%��t�:5�=&B���s�)+�qU��,�=���>�>�w-��%�JN��凼u��=��&�ſA�7�����+D>-��;M�n��ƀ�cw��J �E�����y�LB�]�ܼ@��>9n�>n<p>�6>��U?p��?nu?���>a���繀��ﯾ��0��=?�J�<ɏ��M�������Ѿ�쾔�"������1�&��
!=���=�6R�R����� ��b�,�F���.?�w$>��ʾm�M�
�-<�pʾ/����݄��᥽�-̾�1�+"n�T͟?x�A?������V�'��"Y�K���A�W?GP����Sꬾ"��=����ȟ=%�>Њ�=?�⾰ 3�D~S��A?��?����uȾ;�=&t:�H�I>jC?z��>��Y>x��>�n ?����O0�;>W��=���>�O�>}_�=;X̾K�X���/?�Pq?&Z����o4<>c���舾t�3>��<�S����U��=�{��/�Q���b �h�H>Lc?tWj>�,�W-!�_jľ��"��_@>�?q~?���>�nt?biF?E >=�ݾ��X�<�.����Oa?!��?��?>��DZ侯��k�1?� �?��>�O*��ϴ��uh��
�~�/?:�?hC?�==�ɂ�˕����#�"?��v?s^�ws�����M�V�e=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�%Þ?��@���?y�;<��T��=�;?k\�>��O��>ƾ�z������5�q=�"�>���~ev����R,�f�8?ݠ�?���>������q��=�ە�Z�?s�?k���D�f<����l��q���v�<,ū=�$�vd"�\��^�7���ƾ�
�g����������>PZ@aY�)�>�G8��6��RϿW���[оWq�,�?�v�>��Ƚ垣�X�j��Lu��G�X�H�����jU�>9>'ך�a���`y�®<���뼈��>Frμ��>q�W��绾Sޢ�Ɋ��>��>1 �>1➽�S���x�?�����+ο՜������dX?���?.��?�� ?vD<�r�N|��wN���H?ؕv?W�\?|/���n�WhE�*�j?G_��mU`��4�oHE�QU>#3?"C�>+�-��|=1>���>@g>�#/�`�Ŀrٶ�����7��?���?p���>y��?�s+?�i��7���[����*�p�+��<A?�2>����<�!�=0=�vҒ�ü
?~0?
{�$.�v�P?�X���|��KD������U�>8�D�����=T��}�J��N��Pd�?x@�)�?"���B*���'?_@�>�K��Q���� =+F�>���>�؇>��#=(B�>�[ѾG��>�C�?Ͽ�?�H?�υ�=ϙ��0�=kLp?OF�>w�?��Z>�9?sw��嶺�%z=|�|>2k�=b�=6��>ԻF?A2�>���=T<Z�O��_sD��e�T���K� ��>�w?�/V?UiK>&἟<�����a���ؾ���;��~"�=�	����<>P8 =��i�}��B{߾��?Mp�9�ؿ j��"p'��54?0��>�?����t�����;_?Qz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>@�Խ����[�����7>1�B?Y��D��u�o�y�>���?
�@�ծ?ji��	?���P��Wa~���7����=��7?�0��z>���>��=�nv�Ừ�C�s�۹�>�B�?�{�?!��>�l?t�o�^�B�F�1=KM�>ǜk?�s?*Do�;�#�B>��?#�������K��f?�
@u@C�^?#_׿vѨ�O���$���DE>/��=�q�=h�o��>T-��XN/�!]�¸7>�܀>�>���>q4>5��>��>�"������:��R������
���.��u��Y>��ߤ�����/���Ӳ�;�ͽ�%�7o(�rè�d1�;���5�=��T?>W?p%o?V� ?%�$���>��G��<[�0��Լ=���>�:3?�I?��?L[=�w��?�_����]O���ʏ�C$�>I4I>��>�<�>P�>*��<[*1>��7>
˃>��=W�<఺���<�5U>V֫>p�>�/�>cR<>3�>Cϴ�c2��h���v�?�˽� �?v����J��/���1��A���{��=Da.?�x>
��&?пe����/H?T�`(���+�\ >û0? \W?��>|���T�+H>����j��S>�% �M|l�Շ)��)Q>k?�3j>u>O4�y9��P�q��>\�6?��'�7��ft���G�.o۾�uO>R*�>؁G�@i�9ꖿ�
�#�i��8�=�%:?�o? V��������v��~��1�M>�{^>�=�٦=%�K>��k�O�Ƚ�kG�9�6=A�=�>`>�p?��F>��"=Y��>1s���Qa��p�>4mk>	R4>0�R?R�$?�v�0nV���o��@�Ůd>2�>�7e>��>����)��=��	?�g�>��/���\��rT�tn��1L>*��lǄ��mo�vD=�sҽH]�=�"�=��F��DH�[��=�~?���'䈿��8e���lD?P+?� �=p�F<��"�= ���H��C�?n�@m�?��	�ڢV�1�?�@�?��ѷ�=}�>׫>�ξ��L��?��Ž>Ǣ�̔	�[)#�cS�?��?i�/�Sʋ�-l�i6>�^%?�ӾCR�>g�!�M����冿��y�{�=��>Z1Q?�Nݾ/���{��?�@?��ؾ�p��@U̿{�x��G�>��?���?~,p��;��.VB��x�>���?�h?��b>"���*����D>{�I?[�P?]�>������T�>���?2	o?��H>^��?�s?���>�tw�a/��)������=~=�P;9��>�>C���BGF��ѓ�j^��P�j���1�a>G�$=��>EC佨>����=/9��D����f�@��>>q>ȲI>�V�>�� ?�d�>R��>r�=2M��ϱ��d���~c?'r?`D2�����ڢ�0϶=�<=��&?�,H?Q3	=3%i�@��>m!W?�}?��E?�J>Wʾj����ſ�,��@	>(D6>(�>&?��n����<*Xu�$��*��>���>�9ؽȯ˾iϦ�:�<�]>�6?2s�>��@>�>)?ѱ�>��I>��>v�f����ٰ�W`�>�P�>b@j?�m?ʼ
?������M�A͓�ۃ���M8�U��>��?-G??u|�>�T��Ƈ���7�څ��}H>$�?E/�?.�-�J"\?k|?5�l?�bZ?Z�>�Ⱦ�0׾���3G�>M"?ܽ�oD���(�!���?sz�>���>
u�����D���u�b�꾼W?Z�f?w�)?W�����c��'����<Й���!<�R�<������=d>Xj��o=a�>��=��r�K�4�g���V�=��>#�=��'������)?�(¼�_�|%�=��p�NpA�ik>��?>�,Ծ	�^?!~��)r�V����Þ���C��5�?�I�?��?�벽�f�R96?ֵ�?Z}?F�>�U��ݾB�Ծ~�~� @y�'���<>2b�>��v�Ֆ���1��b�y�Z�Ͻ8	#�!o�>���>0l?�;?�3P>o��>�����&�'�uw�)�]�����8���-��]�)���V|�������-|�I�>e���렲>=C
?/h>�|}>�V�>��˻-�>PT>|~>돤>�-W>V.3>%��=nU<v$ʽN�r??j�y@��4%��)��rv?�X�?Eu$?��>]Y������o,M?R�?���?�k>jf��FL�ؠ�>��_>~�W��?G����,�&�<W���b�|��8�h �=A܎>�佉�.��mQ��'�s<)?�E?�>�*��� ��������<}܃?�'#?M(�=CQ���n�?\��W�q���s�Tɪ��#(��Pt�����;���3��,�&�OQ�=Lu+?Ў?I���`�/1����s���;��e<> 2�>���>�`�>.�=Y��;6�;DS�͌��,B��� ?Y{w?�f�>�xI?�<?vP?mtL?���>P8�>�����#�>w��;�?�>#�>I�9?��-? 0?[Y?y/+?"c>�w��!���y�ؾ��?�?"/?�?��?�_��,^Ľ ���a�F�y�񘂽�x�=��<��ֽ�s�ޔV=�S>W?%����8������k>��7?l��>���>]���$��IM�<a�>�
?�D�>�����yr��]��O�>���?��,�=��)>�!�=����߄ۺ��=O�¼���=@���hY;�R�<$��=j�=��w��Y�����:vJ�;�P�<��>�<�>s�>���>�⍾��gb ��]��y<$��%�>�Ŋ�P��Cd���f��%�M�T0+>>��?OD�? C>�2>�{>�۾{ ��_��*���&<>r��>��7?��i?�ƨ?�a?��0?w�1>�H�;����|s�)���z�:?"",?���>���{�ʾ쨿-�3�H�?(V?A=a�u���7)�¾��Խy�>�@/��~�����eD��̀������-��?���?��A���6�L_����pm����C?���>�U�>���>��)�$�g�P��;>���>x�Q?\{�>�M?�Yz?�Q]?�iW>�:��f���f��>ؼ�P>��A?q�?��?��x?��>�>a9+�� ھr�����M��]h����6=�S>���>r�>)��>�1�=�ý�*���9�{��=�e>��>�ͣ>:��>��><�<��G?���>�s�����ा9ۃ���=���u?���?�k+?hL=�w���E�������>e�?7�?\*?�KS�C~�=��ؼz����mq���>�}�>,)�>'ɓ=�2C=Z�>���>���>�H�Uh� s8�F*N�_�?F?���=��ǿ��;�li�eg��=��>�4���	ξ3��nԁ=��p>�U� ɾii�G0���$ɾQs̾�؅�*[O�B���5�>δS=�B>���=hn=��>R�=�f>s�)>�3�=���p�;�7�<�uE����=�*5=5��oV�=YJ:݋��mYT?�g?��J?��+?x�>	T�=�A�=��>�ii�o�?��>��p>�T��eÙ��#��d��Zľ0��zU5��灾8_=�U�+0�>Ʈ=�)ѽ�J����=k�~<�>S=�=C�
>$�#=���=� �==�C>��=V�Z?�%����3to�����{`�>�U>=,񪽣�G����>�_�==������)S�ɇ?"� @���?�7�>{��M��>nq����e�]�m=a���T��>o�>�؂��s�>Hz>�� ��͊� Z^�_��?�@q�L?q5��{:ӿ=��=w B>|&>��S�8�3��9a���c���L���#?�7�K�Ǿ�+�>���=��ھ-����5={U0>��=�A���]�%3�=��i�k�J=���=L��>��<>�m�=N䪽���=��o=�`�=R�I>Z�һOH��F�g�(=��=ϲf>D�0>���>��?+b0?�Zd?�4�>y"n�AϾaD���6�>��=�F�>B�=�zB>֎�>�7?j�D?��K?.��>vÉ=;�>��>��,���m�ue�Hɧ��L�<���?s͆?θ>�!Q<�{A���2c>�Ž�p?�N1?�m?}�>���v���K6�� /����$<uZ=�����ֱ���)��?���"½9x�=^��>�>��>ϋ>�f>2�I>���>�">#�Q=ށ�=�S�<�Қ<����l�<\B��%=��ɼ����(�c������(��*�u�[=��T����<���=��>�#>.��>�c�=!���y�(>�Ɩ�+O���=*����L?��d��"��F�,���0�]�D>��f>�"��E���k� ?e�_>k
B>]��?�=t?��>���
E־DV��2�p�#�=��=�;�=�D�+�=�ؘ]�YsI��Ҿi��>���>d�>��l>#,��!?�E�w=	��_5�s�>A~��!��X)��7q��=���򟿯i��ZϺ��D?�F��2��=e%~?��I?�ߏ?a��>zH����ؾ10>=O��$�=��(q������?0
'?z��>��n�D��dǾ�-㽲��>�<��
O�ɣ���;/��n��6ľЮ�>
����Ҿ6�3��?���f��t�@���z�۸>�AR?���?�&��� �K�#Y�B��M>?m�`?�g�>[p?З
?����Gܾ�ޅ��=��j?-�?_�?	>>���=Rµ����>�m	?4��?<ʑ? 7s?�7<�QB�>ȹ};�">�\�����=5>¼�=v��=�?(w
?�'
?���L�	�|����d�\�pd�<`�=�>r��>e9r>Ә�=�Df=K��=0�Z>�0�>�-�>Y�d>���>���>1�¾����@#?Ӗ�=r�>�2?Sj@>f�<�2�x=�N�Y�*�܊+�����?���~�X>��X;Y=~���H�>��ǿ�f�?���=&�V�?��꾾|4�?V>��->4�,����>�#�=j�x>�ѡ>�>e� >�G->rUQ>�FӾ>����d!��,C�L�R���Ѿ`}z>����F	&����vw��dBI��n��zg��j�H.��D<=�J̽<1H�?����k�%�)�����A�?�[�>�6?�ڌ�r���>���>�Ǎ>�J��c���Tȍ��gᾒ�?>��?a� >ͯ�>�B?v�>uq/�CFҾJ_�Sǂ�x7��e�`�U�����Y�Ց=��ί�0M?��?�8W?��>���>���?��;�����C��>�#���,�"��=�I?Y"�4JF��n��t��������>9��?���?G�?�'\������2>�]H?��O?k�q?g|,?j?$=�;�D�>�{=ԃ:?0Q?%?�?E>e>��=��ȽE�=�߽�w~���H�1�9������_;<��=/gS<��<��-=Z�=b��x��ˀc�����=�4�=��={U>|��>��F?�?, �>Qd&?��"�,8���� �?w{�=T�پr�Q�����f�X�>��]?�V�??�m?V>��H��DG��| >�5s>B3J>�tI>У�>6�Խ*T�*"M=YZ�=�rC>�zI=;̽����P��L���	p=-�*>��>��C>�ȼi�>P���FԾ��r=�]���	"�K���ye���;�ƂU��g�>Wy?y??�_�=^]��+��=��H�7��>�%�?y�?wd?G��=�|~���%�3U�T�>������>��3��Դ�0���o6�u�<�F?�o��tᠾ�Tb>-��s޾2�n��J���羲EM=���PV=(�Y�վ�5����=�"
>���� ����7֪�Q1J?��j=�v��qaU�0q��E�>���>�ޮ>��:�[�v��@�ů��~5�=Q��>L�:>�[�����d~G��7�.=�>SE?�U_?�k�?�&���s���B�����X`��/ȼA�?�u�>�e?ZB>��=����v���d��G���>��>��Y�G��7��/*��Q�$����>p9?h�>�?��R?��
?$�`?P*?�D?h&�>���V����A&?1��?��=��Խ+�T�� 9�FF�n��>h�)?#�B����>M�?ݽ?�&?�Q?�?��>� ��C@����>�Y�>��W��b��,�_>��J?ٚ�>k=Y?�ԃ?��=>U�5�ꢾ�֩��U�=�>��2?�5#?E�?���>���>g��8�=C��>#$c?N�?�~o?��=oJ?V�4>�D�>�u�=:�>!��>!�?[�N?"Ls?:J?��>�}�<鬭��ٹ��Jt�}x;��.�;�N\<��u=�V�Az�	��5��<���;�������Ț�G2B�1m��;Y�;N��>l�=,';��\]>o���߳��7>W�K��3ݾ�ɒ��>(jW>'v)?�?�(�=�O>W�>�ú>�(�ED?���>\ۿ>�啼�8<���۾Be*��">��'?��A�� i�:7��W�<�jɡ>柀?x?�ޑ��n��*e?�IV?����<���žYK�i!��qe?N?��I��.�>��q?� c?ji�>,�~��Ow�rߙ�sNT���n�U=B��>0��(�P��N;>��)?�1�>:��>�i>��Ᾰ5~��C��l!?�	�?��?=Y�? T.>'[f��l�=�����nX?�>C���d?�Y�.Ѿ�f�ѓ������ڼ��/Й�������������� z�=��&?Dn]?�_q?�#D?l\���o��]Z���{��\:��Q�&���W��8;���7�ƛ[�$˾���j���?�=K��A����?��'?La0�7n�>�˘���;n�B>/ٟ������=�a���A=Sk]=Vh�m.����W+ ?�I�>1)�>u�<?Ž[��,>��1���7�ͱ���!4>^��>�>���>�p�:Ğ,�@X�a�ɾ=�����ҽ��u>@�c?$pK?��n?j�rG1�z`���!�t/� =��]jC>9>�_�>�
X�����;&��`>��s����$����	��K�=�2?M�>D�>5"�?��?:<	�7 ��+�w�/d1����<��>�h?�(�>(�>%�Ͻ� �/��>��l?��>�͠>+猾�N!���z���ƽy*�>s��>�7�>��n>O-��[�S��
���&?9����=&�h?���ɂ_��f�>�OR?�a��Y<��>�	t�-� ����%'�_�>2t?UT�=�<>P�ľ-��6;{������Q)?n9?8�*��T~>�"?f\�>-�>�/�?#�>	nþ��й2�?��^?7J?~SA?nV�>�=�L��f9Ƚ�&���,=g�>��Z>�_m=���=���?M\�ux�[VD=�i�=ީμ�$���<�ϵ�7�J<��<5�3>|�ڿl�K�(x׾y,�Ȑ���	�	���Z��u���]	�ﵾ�����ox�j��l�1�y�T�a�d�%���
(j����?p��?
j������;嚿���1���e�>o.n�k}�&��� ��1��L;�:����!N�ǥg�wBd���'?T�����ǿ���S9ܾR! ?�A ?��y?c�L�"�ّ8�r� >h;�<{>����뾯�����ο������^?���>{
�(.��=��>Z��>��X>�Fq>8��D螾�E�<��?h�-?ڠ�>t�r�˕ɿw������<��?�@�>I?�|�Y�S=(i?0O>���V6�L��GȾ9��=8��?挼?U��>b�R��B$���?�(e>�!������+>Jm~>��>�����=��>����Xr�O�����?>i/�>�jb���C�αg��{p�� B>n�N�Ub���Ԅ?�z\��f��/��T��S>�T?R)�>�0�=v�,?�8H��|Ͽ��\�<+a?1�?��?l�(?�ٿ�pٚ>��ܾ��M?UD6?��>Vd&�R�t�d��=$=�sp����㾯&V�i��=��>F�>�,�����O��T�����=���ƿ �$��q���=����1]���罅4��NMV�g��TVo������g=\��= Q>�>�V>�-Z>��W?tQk?���>ʿ>���勉��ξ�\��́�J��=���P���У��M�x�߾
D	�q�����^ɾ=�Ѝ='!R�����
� �q�b��F���.?�$>��ʾY�M���(<�oʾ�����������4̾��1��
n�Gӟ?OB?������V�T��O@�V��W?8q�����笾�+�=����5=g�>
K�=��R3��eS�/�0?��?�����̒�;�(>�'���e*=�b-?_?�`<�,�>��$?+��@彋W>�*>T�>)�>�>{_���ս�?=�T?�7
�~v���ē>���:u�0�L=�+>b�1�ORѼ��[>�u�<����pH4�T~��P�z<��k?�|>G�c��Ug����ڰ>�dk>���?���>��>]��?�f?�����?�5�i��	ؾ�>�B�?��?�"�=x�=<:��3�6��A??��ս�Cx�|羃8��t����>��v?�b%?njӽȠ���ṿ\r��!W?��v?L[^�(���{�Z�V�z1�>|��>��>>\9�ӯ�>��>?\�#��K��iѿ�ut4��Ϟ?ח@��?�K<���D��=�3?'e�>e�M���ľVG��"�2m=*�>J����eu�)�#],���7?&�?~M�>�ف��;����=�ٕ��Z�?��?}���|Dg<R���l��n��j�<�Ϋ=���E"������7���ƾ��
�����࿼ͥ�>EZ@�U�v*�>�C8�]6�TϿ)���[оSq���?M��>T�Ƚ����A�j��Pu�b�G�3�H�ť����>��~=a��c���灎�f���ȗ=?؅>� �=	P?���� �ݾ�־J�3>��0?,�J?�L>�7M��\�^ �? ����Pڿ�+�����D`E?!q�?��?�qb?byE>"Y�=M]��ؽ��?��R?�+6?	
�4w���m<��n?�͔�Bqd�E�<�4�1�o�U>�=?�h?� �vW�=�R>c��>��=إ'�.h��{̺�������?���?��*�>�=�?�w/?�-�����^@��c�s2�=��?�J�=�]����k_&��g��,?XW)?��(�#+��M?�M@��Aq��1��1�ҵ<�D���K����^�������f�>��w�;���?�/@�ͳ?h��P�	�;?��><�~�fe5�r=Ȏ�>��>}'�=�ҫ���=�+��z*��e�>Gg�?��@
�?�W���N�>�o?��>�*�?FT�=�?u`%��F����='�=�uS=<!h��0?z�!?�w�>lF�b(���i3�͋Q�]j�GT׾;zG�[��>5�[?�?M�V>h�<8k(�G�=�H{=z5�,�1>/�}%���ͽ�>>2>u%1>�	;��8��!�?	p��ؿj��=o'�i54?���>z�?���6�t���{;_?�y�>�6��+���%���C�0��?�G�?��?��׾\I̼3>��>�I�>��Խ����������7>��B?��aD����o���>���?�@�ծ?�i��	?���P��Xa~����7�u��=��7?�0�.�z>���>��=�nv�޻��U�s����>�B�?�{�?��>"�l?��o�Q�B��1=@M�>̜k?�s?fRo���[�B>��? ������L��f?
�
@u@d�^?(14ۿ{p������d��á&>+�=�?>�?�;﮼��5�pݝ�Yd��Z��=�\>��)>�k7>�g>vw�=�	�=���p��9����?���*1��������bn!��𠾰�S�ξ����y���ێ�G����a~�X��1B�	��=W~V?h~R?e3p?�O ?À���>�&���G�<��"�R�=�m�>��0?�IK?�*?@V�=�+�� $e��P�����*��m��>�wH>�e�>� �>;�>�H�:�TG>�<>M�~>x�>�;!=�����0=j�N>��>%��>�h�>�C<>��>Fϴ��1��l�h��
w�f̽1�?|���Q�J��1���9��զ���h�=Ib.?|>���?пe����2H?&���{)���+���>|�0?�cW?$�>��r�T�9:><����j�/`>�+ �}l���)��%Q>wl?fih>�x>h3�(L8�=�Q�
���\��>�$7?]����6�)Iu��"H�&ݾ��J>X1�>�<u�{��O����~�o�n�z4�=��9?vH?�(��+���"|z�������J>��[>�=h�=�5H>�?i�M�ƽ�:F�	�'=���=lh\>�?��,>p�=�>U���P�p
�>	�F>B'.>NR??P�$?�2�Ѿ��W��(.���s>I��>&��>Z>�K�pʳ=���>sHb>���Ƅ�.[�h�>��nW>�x�lb�S�w���w=�~���!�=�o�=�� ��Z=��	=�aj?(���^疿�8�4pŽ�>��)>TF������I�z���K�����?s�@8!�?lT���46��DT?�\�?6_=�պ�� �>8�>-z�	�>�b�>�	��$���)�ٌS���?#˾?����࣫�^<a��%h>��+?�?��i�>;w�sZ�����i�u��#=ު�>�9H?yT����O��>�Ev
??u^򾨩����ȿB|v�t��>�?���?��m��@��	@�~�>o��?�hY?�ri>�d۾odZ�[��>�@?�R?�>�8��'���?޶?���?5�H>*��?u2s?���>�����w/�����߄�����=}�;O<�>fv>���JF�z����J��g�j��&�{�a>ݒ =�>ۨ�HW��^��=I5�������1j��η>W�q>��I>O��>[� ?2>�>H��>�Z=�슽"���C�����K?���?&���2n��:�<���=ү^��'?�I4?�_[���Ͼ;ը>��\?(?N[?/c�>o��>���翿�~����<n�K>�3�>�G�>�*��XDK>1�Ծ�7D��p�>Qϗ>��
@ھ-���D���B�>e!?U��>Ϯ=�� ?�#?g�j>�$�>`E��8��Q�E�;��>��>�H?��~?��?VԹ��Y3�x��[硿��[�c;N>
�x?�T?&˕>���V����F��@I�%ᒽ}��?�tg?�`�Y? 2�?͉??��A?Q+f>0��Nؾ歭���>[�!?���@A�'�%�/�"?�?��>Ƒ���n׽]������p���G?�\?x�&?/�Ɗ`�+¾^}�<����$��N<H�I��t>��>=���d0�=�q>��=��m�Y�7��_<3�=lʒ>C��=��7����E,?McJ������=J�r�"KD�.	�>vL>~����^?T�<���{�K��S���EU���?���?+s�?՛��ώh��=?��?�?2�>X����޾9r྽qw�u
y�zc�{`>�	�>��l��&�l���o���9��	yŽ]N�K��>��>�?���>��M>�C�>g��`�&������Ƃ^��p�RZ8�n�.����A��`%��@��,¾��{�ݛ�>J���}�>��
?��f>��z>1��>�Z���:�>�#R>� >�O�>��W>|�4>�>8<#<X�нg+T?�+���(�Ͼ!v�w�?��q?��?�w#=�i�_���?A�?��?Yl#>lka�����?O��>��J?��> e�<��F�:�;ج$��;����I�>)׭��?�tI�J?/�Y�?_V+?(����ǷJ�򌠾�n=�M�?��(?��)�&�Q�E�o���W��S����6h�^j��!�$���p��쏿�^��
%����(�s*=�*?#�?<����"���&k��?�cf>��>L$�>K߾>sI>��	�H�1�^�PL'�~���qR�>8[{?M��>�I?�<?=wP?�iL?���>�a�>=6��e�>��;M��>F�>�9?Q�-?:0?+|?�t+?o2c>u��8����ؾ�	?ڥ?�H?�?ͮ?݅��cý���<�f�e�y�d���
�=?@�<��׽R[u�\�T=�T>�20?k��R�Q��&'�h�>`�!?�S�>�T?ܙY�y�b�%�>��>��>��$>O�������+�t�>�3�?i�t��n�=���>��T>���yϽℑ>�Y=�>�b��������=$M�=�v1>�r=�8ʽ���<�H
�K��'u�>�?E��>DC�>�@��� �0���f�=�Y>KS>H>�Eپ�}���$��}�g�3^y>�w�?�z�?C�f=��=��=�|��ZU��~��������<��?J#?�WT?S��?��=?uj#?ӵ>+�|M���^�����ɮ?N4)?�ۣ>B���Vľa��7�<�^$?9=?�a�<�?;%��¾˫��tW�=��-��]|�`���z8H�����C���7%�	��?��?.VW���9�W��� ���O��(�6?3��>��>�d�>#(�Wd��c�=�6>�e�>��N?Z)�>��O?�2{?��[?�>T>ۙ8��+���ҙ�k�7���!>��??.��?G�?.y?��>v�>I�)��߾�D�����r��͂�AW=��Y>	��>�"�>Zݩ>��=?�ǽ�����)?�V��=��b>w��>���>���>�w>)K�<kZ?�z>�>�)�d�_���������>t?�ә?J��?Ѧ>8�:���g�� ��>��?U��?,?Y�[��/>O�p��3�E���96?��>6��=_"�=����ս&�N?վ>�����U�a��lG
��S?��u?'&�=�+Կw�*��A1>~�.��c�>�͘�#\�z��SI׾9�����W�c#P��ҋ��\��|��p��&~�;���@|?�/�w��=zpV���u��M�q+��^���="�
=*����U�=�kһ��������7=A���Q�=O�m=UӾX��?�vi?�=G?*�>~>V6>?-C����=��>߬+?���8��<�������i���B6�F�Ǿ'�w��Q��D�I>0sZ��G�>��>Vf�<D�>��R=k��=�(ͼߚ����=�´=Xf�=��=4U>�D>��=|6w?4���ò��Z4Q�r\�C�:?r8�>Zx�=i�ƾ'@?�>>2�������a�a.?���?�T�?L�?�ri��d�>����⎽{r�=����>2>��=��2����>��J>K���J��僳�A4�?��@��??�ዿ��Ͽea/>�<>���=��R�yb0�D7S�I2d���d�}�!?:��\;a��>�=��ؾ��ƾT�=�7>O��=�>�8V\����=8�v�jM?=��=���>"�C>45�=M����-�=W�==9��=6#P>C�C<���(��48=��=��e> �&>ZT�>s�	?i0?�t`?���>Eow�u̾�&վ�2>n��=�AU>)�=�� >�6�>�hK?]�Q?�zK?L.�>!��=�>��>��#�ɥ`�������7�k=���?H�?]��>�^=��i�J�%���8�B抽��?�i?��>�O�>7<���4�%��C.�"���vuI���(=�"q��6W��6 �- ����@�=���>���>�A�>�fw>�D9>�M>1�> [	>���<���=��g�n}�<*f�����=�~�����<�MƼ���,�,�"�)��G��-�;�z~;��b<?��;[��=���>0>��>�O�=���GS/>\����L��ǿ=pF���*B�N3d�^G~�S/��a6�ϛB>�X>�|��65����?��Y>��?>���?�7u?��>�O���վlP���%e��SS�顸=Q�>=�%x;�~V`��M��tҾ�T�>���>���>�]>y�2�`E�C�=77о��4�4��>X��u�E�v]�I�m�<ܡ���k���I�=?&`��-�>aIy?4bT?p��?H��>�D�L��]�>	B�����=S)�50��Ҫ��dx?�.!?C,�>7,���<��Xξ'�/�V5�>�{��2N��^��\�2�� ���*m�8�>�)ƾ~���+����ش������!W����>NJ?�к?#��
M{�4�A�9�����y��>fwE?��>B_�>�x�>8T���վI(,��}>�J�?M�?�
�?p�F>@��=�<����>g	?���?kő?`s?�U>��;�>5Ԣ;f3!>ՙ���=
`>b"�=\&�=+M?vQ
??�
?	����	���� �5o^�D6�<m��=�ƒ>�j�>"�s> ��=�g=D�=�h\>m̞>��>îd>3�>�s�>����O��%??��=�Q�>W1?*@y>��J=�P��ӂ�<�S���>��*��Ժ������<�
��k�3=����O@�>�ǿe�?��E>	
�AJ?�"���qO���\>2aS>C���X��>�&A>ZAr>���>�m�>.J>s��>�51>GӾ�~>����d!��,C�'�R���ѾA}z>�����	&�֟��w��SBI�pn��ng�qj�L.��G<=�u̽<:H�?<�����k��)�����1�?x[�>�6?/ڌ�s��A�>G��>�Ǎ>�J��`���:ȍ��gᾉ�?,��?ք^>�M�>�@V?]_?u@���M��8Z�ҭu�p<�Dc��Tb��͍�����Y�#]���nd?�'w?��@?�, =�щ>ѽ�?��,�s܏�Aĉ>��3�z�;��KA=���>k���u�d���־�w�����v>��q?b�?�/?#^>�>�*�AzO>kyK?��?��u?�O?�+-?F��<<�(?�¬>�B?�U�>$�>aa�>d�>��C>H>�ػ)�=�2ɼ�މ���I��Ǿ����<�J0=�j�=-�ټJU�=��;�D}���:;���<�=K�������<`�z=�=bB�<N��>�Y?6��>f�>}*1?�!���6�+���du$?|%=ed���X��s ���Y�"'(>�'o?���?��Y?�5n>;�L�:���>:��>t�>��e>�b�>�=���@4��]�=��>�>dcr=�\�D�v�C|�쇘���O<��!>�>��>�鹽1>p�¾�8����>����ҹ���+� F�-�,��|�<G�>ga??K ?+LT<�����n�)X1?]�4?~9X?`9n?��d�[����:V��@U�������>J� ����oJ�������0�1zr���>A����۠�HWb>.��Fr޾~�n�5J���羣#M=��YVV=����վ�1�|��=�#
>���� ����Uժ�s/J?��j=#z��]U�#p����>X��>v�>V�:��v�Q�@�P����:�=W��>� ;>.[��m���{G�(6��U�>��D?_?@Q�?ma��F0r��~B�b �����ſ��!?�J�>Y?�x@>fU�=�^���}�_De��F�/4�>���>�>�+G�����(�D�#���>p?�I!>�*?�"R?�6?[�`?e�)?(1?z��>	����n��Z@&?���?%�=�0ս��T��9��F�s��>�z)?h�B���>�}?�?i�&?s�Q?&�?7�>�� �K8@�d��>�Y�>��W�T]��m�_>��J?��>y;Y?ZӃ?��=>��5��⢾zϩ�9�=�	>M�2?�2#?q�?U��>s%?�8k��5>?u�?�jq?C�]?=�����>��=BA�>��=��>���>V?\8?YDh?F�]?J1?K�b=8^�=�&
>� ����J/��AӼբG�/�)���ݽ:A�:#`=���������=��>�T9>[>N��<�Y�>�s>�ꕾ-=1>��ľ�/����@>�"���N���ϊ�d:��|�=���>z�?��>cb#��&�=�z�>T�>=���)(?ʼ?�?j�G;�~b���ھ�`K�V�>��A?H^�='�l�0v����u�*�g=?�m?�x^?AW����'`?Ҳ�?��U���j�q�辨,���J���e#?��\?`!�=���>���?��~?�?����8}�
!��(h��Aګ�2��=r��>���-Z�م�>25?��"?��>ۊ<��ގz�ޤ��;.?S��?ө?��?o��=8ꁿR<���=����c�[?��>� ���8?8���w�`���ִ���K��i<��Ā��a5���ћ� �b��y=_��=| 6?��?ލ?$�?@�'��d����\� d�B\�����KF��n�Ez�UH��3M��(����Y�u�d�\�>������A�#v�?E�'?�#1��F�>����1�G̾�lB>q��}���#�=Em����?=�Z=@�g�ה-����W: ?��>^��>&�<?�\��'>���1���7��
���3>
��>�*�>Y��>�Ad:��-�����Aɾi�����ӽ�Ԇ>4	S?<�T?��c?i��-��m��Kg�EXu�Kw��7��>��>�i�>ŧ��^(��3:7���X���|� ��P���|(��y˽�f?�7>�?���?���>y������>I���O+���>���>9�<?��>h�>��;pҟ�=��>��l?-��>L�>�{��<h!�|�{�I�˽���>��>��>�op>��,�+\�&f��z���b(9��*�=�ph?����a�U�>lR?�e�:��Q< g�>�x�|�!����J�'��>=l?,�=�Z;>�gž����{�[ډ��$)?5?�����<+�m�|>g!?���>�ԣ>P��?9$�>��ľ�p��Y�?�'_?cK?��A?|d�>��=8����ǽl�%�#o%=ч>5Y>/�q=���=4��'[�8���A=3�=��ͼڰ��]�<�#��S�T<8��<�r3>�lۿ&CK�(�پ�
��>
�_舾����Ec��t��ja��D��DXx����'��V��5c����l����?�=�?���+1�����j���r������>p�q�����������i+��M������c!���O�+&i�*�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >^C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾r1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@FtA?��(����W=y��>@�	?��?>��1�;C��㰾�c�>G8�?���?y�M=��W�Y�
�0^e?ݻ�;g�F��޻��=���=͑=����J>�a�>�7��:A�r<ܽǞ4>�̅>��!�|n�aU^�K�<O�]>Aս�Ɣ�8?�-\�Ьe���/��G��W�>'lT?�>���=�1,?�nH�$~Ͽ��\��Ja?;:�?|��?;�(?�ſ�A�>��ܾcmM?�5?2�>�a&�ht����=��ݼ,f��k��k V��J�=�{�>\�>�,����3O�Q���Ss�=Q���ƿ
�$�*4��C=u]��ZX���Nm��l�X�x����%o��T归�k=V�=�GQ>�s�>��W> �Y>�qW?�k?Ψ�>�>6�罼���|QϾހ��逾�8� (��l��(��(��q�߾�b	����T����ɾ� =�J�=�6R�����H� ���b���F���.?�u$>E�ʾ�M��~-<2qʾS���RÄ�Xۥ�-̾�1�m!n�6͟?��A?����d�V�?���U�R���E�W?O����SꬾX��=^���ڜ=�$�>��=��⾲ 3�y~S��s0?)U?Ą��rL��aG*>�� ��	=-�+?Y�?Q.[<>(�>I%?-�*�a:�b[>��3>G֣>���>F	>���+۽�?�T?A��>����Ő> n����z�6�`=�>�25�3��%�[>��<�挾0T����ɉ�<�(W?m��>��)���ka����Z==��x?Œ?b.�>_{k?��B?�פ<h����S���(_w=��W?*i?��>�����	о����C�5?ۣe?��N>bh����)�.�GU��$?�n?,_?T~�� w}�x��}���n6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?p�;<��U��=�;?l\�>��O��>ƾ�z������1�q=�"�>���ev����R,�f�8?ݠ�?���>���������=ڕ��Z�?h�?����xLg<b���l��n���w�<�ͫ=�SH"�����7�f�ƾO�
����㿼c��>NZ@T�p)�>�C8�s6�TϿ��N]о�Sq���?��>y�Ƚۛ����j��Ou���G���H�����ud�>Y<>��h�f����zz�$�=�"��I�>� <��z>Eh���� ~��φY<i
�>�D�>���>�x���f�����?�X��LU̿�7��XL��WS?,7�?fd�? �?��:x��	w�!b9�!J?5�u?(UY?�xN�1Qf�DO!�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.���I?%�,����d_�,�۽s%)��Ӿ3��j�q�w��8����K��e�޾�̪?Q*�?/ھ?��[=��B"-?�,�> (C�Bþ���c`�>��p>�2�>�vD�Q�>T���2�)��=��?H��?5/#?-�h�'���_=��zd?H��>o��?��>�%�>	��<p��ՠ��e�b=�Kc;J���?W~d?.T�>؛>+�N���C�$$`���j��v^�)�2����=tݎ?�pi?.��>UT���]1�ޘH��k����_�>�0)�
ﭽ:݆����=P2�=���=u>������?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ta~����7�W��=��7?�0��z>���>��=�nv�ݻ��W�s����>�B�?�{�?��>#�l?��o�M�B�T�1=7M�>ɜk?�s?Ro���e�B>��?%������L��f?�
@u@`�^?)�Y޿�����B�������'�<�E.=M͊>@��=6^=��e=��6=I�=�f>b�>f�>ԡ;>�5>��@>��>	�����%����J#����B��c���e�8�9�߾�I�[���H�7�v���T���hh��=+�D�����a��=$�K?�K?i�o?���>/��^#>~?�丏<_�����=p�>+�2?soI?�~?Ξ$=�੾!�d��B|�J����͕�G��>{0N>���>G�>Z�>l`C=��N>n�9>~�t> �=;�e=���<�4=k�L>�C�>�v�>���>�C<>ӑ>Gϴ��1��g�h��
w�]̽-�?o���L�J��1���9��ɦ��$i�=Ab.?�{>���?пj����2H?'���m)�ʹ+���>o�0?�cW?"�>1����T�M:>3����j�$`>�+ ��l���)��%Q>nl?:<g>bv> �3��u8�R�P�7��{>�6?N����Z9���u��bH��0ݾ�QN>���>��J���,����]�!�i�rVy=B�:?��?���ip��%�v�����.aP>-�Z>[ =˗�={ML>��g�&MŽЕH���,=M��=�!^>�H?� >rх=�u�>���9�A�X��>��=>��$>'�>?�%?��`2t��]z��B0�1/c>�n�>�u>u�>%�E���=S�>��\>�K@�x�������c3�>�W>cy��k�b��_��b>X=a
�����=���=#��H,��s=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾQh�>tx��Z�������u�v�#=P��>�8H?�V����O�b>��v
?�?�^�੤���ȿ5|v����>W�?���?f�m��A���@����>;��?�gY?zoi>�g۾:`Z����>һ@?�R?�>�9�|�'���?�޶?ԯ�?C/M>���?I�v?���>��;�
b/�5I���ӏ�D�< I����>�� >0c���qF��ɒ�]���9m�i��2�D>�f=���>)��.������=~ҼM|��1铽��>Yi�>�8>#��>J{�>A^�>Qn�>1�-=cz���]�����QL?P��?��E�3Yx�o���6�<dm ���>^�N?��i=`ҾSy�>�Z?^�?j�&?&�>�}"�`���%�ҿM'����뼭z�>��?~K�>����H�<&���OǾ�З=�t�>��
B	�vБ�.02>�t>H� ?\�>ڀ����?� 8?�o=	�t>��R�å����L�H�[>��$?�T(?�'f?�Z?4�о�M�����V���h[T��?]>��s?,H?!�>ˮ��⭦���gl=��=�r?�4u?<o�=�/?gǟ?̄?ya?5}=����wP>�y���F�C>�� ?S���;�E�*�N��:?G ?��>(|��U{ ��M��������5F?&/a?5�*?��Z�^��(���+�<_����ρ��5�<8۝�p*#>�>�1p�@\�=�>�=9�f���3��e�;���=Ac�>~��=P5�W��<:,?oF��у��ߘ=��r�4xD��>�GL>%���H�^?��=���{�{���{��	�T�� �?��?fj�?����h��!=?��?�?n1�>vH���w޾ӌ�xPw�)[x��r�6�>���>��m���򐤿����<����Ž�����>��>��?a� ?��P>?�>򗚾B�&�)��8K�C]��4�\�7���.�w����eA%�e�����x�}���>�⌽�|�>4�
?$i>ؒ}>��>�Ɂ��z�>�Q>%6�>�1�>��W>�6>��>�\b<k�ɽ<R?����r�'��M�𗰾Q'B?;pd?2�>�ii��t������t?�~�?Qi�?y�u>2�h�:5+�TI?\%�>����j
?��9=��Y�<�G��4��.���c�^d�>��׽=:��M�=�f�O\
?�"?7s��2F̾��սK}���so=�O�?��(?��)���Q��o�n�W�`S����g�QC��Q�$���p��ꏿv_���&����(���)=�*?L�?r��b��6
��k��?�F*f>*��>W/�>C׾>�VI>��	�ڽ1���]��C'������C�>�a{?�΍>�6I?��;?�|P?*�L?�> l�>�#�����>ǽ�;�>���>��9? �-?W60?�o?��+?F�d>p����q��,�׾?�u?"�?͑?	�?�~��t�Ľ8����q��y��能߼�=m��<�ֽ��r��~W=U�S>��?�,�l�%�LȐ���>D0?}D�>Bѫ>�ᇾ��*�6��=�&�>�?�(m>���9�e�[?��V�>szy?�Z��(Y=�Y�=D�@=&\�=��;8�x=�N�T�=9�=8$��뼮��=E䨼A]��Jk=�g=��=셸=?��>�/?7iu>�ca>��V�=��P�%�nGT=�hz>�F>ފB��4�d����}��`�c���B>�?ie�?P��=��>Y�)>�y߾��޾�� ���(��<�[�>�]F?�#|?��?�p?�w,?�
*>�\Q��V������xe��>�&?Q�+?潱>�*��̾�ۢ��1<�U�?Yr ?Z?T������N瞾z���}2>�X(�X�~�t���L���g��t㽡a�?F�?Q#f��F@�a���$����}Ծf�%?�v�>�U�>�?�>F�.��V��h�
� >��>`�I?^.�>�H?�Ax?��Y?�U^>|-������������K>��F?�W�?\�?�\b?D�>]i�=�q��|�tQ��?��,B��!���d�=l�:>�;�>�b�>��>��=�\��
�ٽqvM���=*�x>���>8ץ>��>3�>��=��5?!�>��F�����亾�~�+X?j�v?ښ�>�%p���=�Jp���9<?��?,s�?��?����=2��=%8��~~�=���>�:�>cO�>��=��>��>���>�2�>�VA��!T���o�#�h��("?�Q?;��ſ(�q���q�D��W�{<x���:�b�F���b�Z��_�=�����#�`5���Z�#��FV��ez��>؛���z���>[��=x,�=n��=��<�����<Y�N=�=�<K=��n���Y<|�;��Y��,Ή�xk+��me<$tL=zF�ɥ¾g8u?�'B?=V-?��D?�z�>K['>!fE���>��"�n ?�&W>٬�-O��#	@��s������Ѿ��ɾK,_�Sk���>��V�l�>Ǖ5>Lr�=�ޮ<���=?��=#�=aVb���=��=�+�=8�=��=~>�D>��v?�4���Ӝ�ǎQ���TE9?T.�>��=��Ǿ�S>?��8>Vc��ы������}?���?�H�?X�?�g�-W�>�꡾.���Fk�=1���U@.>�<�=!w1� �>�}G>5o��Ԝ����@U�?�@�??����h~ϿV0>�7>�>)�R�:k1�@|\���b�THZ�܋!??;��?̾R+�>���=>߾~^ƾd�.=�f6>�a=���d0\��ә= Yz��;=>l=���>��C>�=ů�/�="I=օ�=�ZO>�/��,9�?,���3=u�=o�b>�Q&>p"�>\k?P�0?�Kc?.r�><�m���̾�^žM��>��=�~�>�= 4?>M�>�c8?��D?jL?3h�>���=F4�>gӦ>J^+���k��l������<�:�?z"�?X��>TV`<ts=�����6>�xɽ�?�1?L�?�u�>��6�ۿ��8��
�]�
�Mp >hPl>��=�=���=i�N=.�V=L3�>oc�>%ġ>�e>f9>�
>��>3��>`��=�U��n��=e�!<��>9>���<�=���=�5����<)�y�@y���]�<��=�$<��;�R<�b̼��=��>|<>ݬ�>C��=����C/>ݸ���L����=�G��c,B��4d��I~�K/�~V6���B>#;X>�}��>4����?X�Y>�l?>���?UAu?-�>� ���վ�Q���Ce�>VS�<˸='�>��<��z;��Z`�t�M�T|Ҿp��>��>.�>>�l>y,��%?�N�w=�⾹d5�m�>yj��y5��#�6q�V>������ki�c����D?<D���v�=�!~?��I?[�?t��>�!����ؾW(0>xD���
=�
�M*q��t�?�'?���>����D�wH̾W��+�>�>I�]�O�����j�0�m��Tͷ�D��>�����оO$3�lg������J�B��Ir����>/�O?��?�1b�W���UO�{���5���p?�{g?)�>/J?H>?�5��0}�s���x�=��n?߳�?�<�?>R�>yL
��U�>=l?E�?Oה?��?Ȃ��[��>>5�=4$V>�:���>�Y�=�8=M��=��>�� ?��?b팽�#޾;���r㾝�D�� �3�I=�'D>Վ�>�dE>�J�=U��=P��=)d$>���>�>�z�>���>s�>����%��?��>��X>�zD?�$L>��G>_3=�`*���;10&������Qڼ}{��̸�<���<��=���ԕ?�¿/��?�[�>W�;�wC?߇&��,켂e�>��!>�E6��<�>��=u�K>[Rc>�|�>�J>Zn�>�>hEӾ�~>?��uc!��+C�X�R���Ѿpxz>����&�����q���?I��m���g��j�Y.���<=����<�G�?�����k�a�)�����N�?:\�>$6?�،��
��N�>���>ȍ>5I��Ώ���Ǎ�xfᾔ�?���?��P>�v>��n?�ټ>���_$����~�#W+���j��Ku��!}�d���V���>n�;��s?��?{OH?�Y]=�8�>���?�����k�6�?�]e�(rN�-�>%�=��������
�F�ھkԼs��>4�?řq? o�>�4���:	>j.ɽ���>N�O?աL?4?��S?3B����>HG	?��"?���>X.%?}
�>���=U�"��]d��w�=�;>ۜ0��U��&u��L`�7�=j�2>�c>�͖>(8h=�h��-!��kT�?⼈�=u3o<���$>��h��=�D�<dg�>ƏN?i�?���Y)�>�a׾�yP�M���3��>[���
����?��������>�6�?�¢?�3?=r�>�&�E볽��<�B�>�>
~>{��>"��Qͽ�O1>f>�">^C�=d}�x����v������=5�>_-�>>؋>�V�.��=�[���M��jI�=�i)�(m��_g��+hW�	�?�V��,L�>sw]?��/?�.>���O���W�e�%?=?$?s�^?"�g?s=�=�]˾�+���-���н��>�=(	�k����֤�%n=�鹀=��>�8��������b>7�	�y(ܾ�m� �F�%��C=�}�(�+=��
�)�Ҿ�fu�j�=)��=y�žo!��S���_��;I?)K�=]�����R���{2
>��>���>8�M�ܲ��{�<�����ǝ=�O�>��6>�ټ���IAI��3�w,�>�_C?��S?(jy?�;��{�k�|*1��:��(����o���?KϮ>��	?�E>�����־e��>.o���:����>�� ?��YK�?s���	���&�fH�>��?�� >�	? :M?�?߇g?��$?���>,wn>6��ܼ���A&?+��?N�=��Խd�T�� 9��F����>'�)?��B����>��?@�?��&?	�Q?@�?��>έ ��C@����>�Y�>��W��b����_>o�J?ך�>�<Y?�ԃ?��=>��5��颾թ�qT�=l>�2?6#?2�?p��>�&?l���xϼf�>�Do?éw?y)g?q=�=�?u��>tF
?`�=>�`�>��?�|/?0h7?��C?��G?z�?��f=�z~�0[*�����ږ;׿��ك��9��=���<��>�I�m���=s�f<�q��*�=��~=6)��7� `�>R�s>���a�0>��ľP��4�@>ˣ��tP��؊�t�:�}�=���>m�?@��>�Y#���=ĭ�>"H�>���X5(?j�?>?�	";Ġb��ھ*�K���>�B?g��=}�l�����a�u���g=��m?^?�W�)#����X?َq?��L�C�Ѿ���@�Ͼ^-3?13&?e�}��W�>��e?l�n?�#?����y�������ل� -��q>!>�q�>�]0�JE~��	�>��?�ˁ>���=0�f>3#d�[r�þ>��>�9�?�ֹ?Jr�?7�	>��Y�e���2�������?��>�C
���S?�����p@��툾ϝ־/豾}��뫞���t�Ɨ{�]�v�?����VX�=�)?k�z?�?��S?�����p�r���
p�X‿v����4�XӀ�"*��\l>�	��ha��n���F�o�p�j;����?���?�&?��1��T�>�x��>qﾠ|;�1:>������d`�=7Д���	=�c3=�l��36������?���>-��>W<?U�\�Z>�ڿ.��'7�����a6*>�M�>�^�>[v�>yu<��-��F��̾c/���ս0v>�nc?ÊK?~�n?�Y��"1����H�!�R/0�vY����B>>3��>��W�����:&��Y>���r�N��q��0�	�~=5�2?(�>���>aN�?~ ?J}	��s��phx�ʃ1�#�<7�>�i?GA�>��>��Ͻ_� ���>�Y?�5�>�^>_m�N��F^�ܶ[�R�>\��>} �>��6>$� ��Di�~��m���L*����=d�R?��h�&��~X?>m~Y?<�_>��
?)V6�i�9�����"=5$w>v1?Xܒ>N��=œ��n�F�长^���-�)?P�?S^���*�Hp}>kM!?��>2+�>˃?��>�x���;8�?� ^? eI?�C@?�'�>�=m岽-�ɽ�K(��;=�-�>^Z>�k=���=���'�[��$���G=���=:�̼�ɼ���;�r��-�R<e�=�:>Oiۿ1=K�1�پ����K:
� ݈�L���yg��=��|\�����\Cx�����'�s5V�'Ec����ڷl���?�:�?(����.��������������>��q����[諾s��T#�����w���;e!��O��(i���e�Ӗ'?��� �ǿů���7ܾ] ? A ?,�y?����"� �8�ζ >e��<x����뾻�����ο����+�^?n��>�������>��>��X>xPq>���b垾c��<��?C�-?=��>l�r��ɿ$����Ӥ<���?�@"A?��(�f�쾔LU=���>cy	?6@>��1��6�Υ���a�>�3�?s��?�mM=��W��z
��Ke?�� <�F��K�4t�=m�=��=���zJ>�t�>"��0GA��Zݽh�4>��>YI"������^��־<�~]>9�Խ�C��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�#�ͫƿ*�$��!��s�<Ng/��W�#��|쩽|�T�枾��m�z��Tck=���=G�Q>��>��W>�Z>clW?��j?�u�>�>��U����ξ�#������yk����9���-��mI�sd޾Ս	�ci��B��ɾ�=��.�=�.R�����2� ���b��F�O�.?c$>��ʾ�M�^o.<x\ʾ�ª�!��aL���7̾��1�"n��ɟ?��A?�����V����0�����W?�D�Z���ܬ�q��="S���c=�!�>MW�=����$3�SyS��:5?*�"?��꾽'���#>�P�m��=Z ?���>�X=0�>��,?G�����59>��=�1c>I��>�>h�U  ���1?�C^?�%ҽ<X���D�>2��񏈾�9��d�>�q��tKмn�j>Rg�_����ʺ��ۼ�=�]V?��>�=)�U������!��7=m`x?�?%��>��j?;?B?6��<����1tT�N��w=x�W?�h?��>5����Ͼ���*w5?*f?�S>:�j���꾄O/�6���`?u�o?z?l�����}��Y'	�P6?��v?s^�xs�����L�V�e=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?b�;<��U��=�;?l\�> �O��>ƾ�z������4�q=�"�>���ev����R,�e�8?ݠ�?���>������d��=�[����?f͆?�8����u<�F�Y�k������>�<qޫ=��:�'���z8���Ǿ��
�'ǝ���ü��>`-@o��51�>7X;��-⿠�ο%Å�9fо��q���?h��>��ɽ�+��*$j��t���G��I�jB���J�>3�>����`�����{��s;�y~����>�f���>X�S��6�����=u4<��>_��>Ć>#���彾_?�S���>ο����ۍ�o�X?�d�?�j�?�v?�:<#w�Ά{�����&G?"�s?NZ?�(%�F<]�!�7�%�j?�_��xU`���4�tHE��U>�"3?�B�>S�-�e�|=�>���>g>�#/�x�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*��+��<A?�2>���I�!�B0=�UҒ���
?V~0?{�e.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?���>�Nr?x&�=��?��>�3ž�l�=gY7>�=��<��?	X[?���>j(>�0���)��@��SK�����8��>hht?��k?'�>2 ���ǽQ76�M�齒埽V]=դ9�[�ĽP��a�>�r1><��=խ�[����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*��ۿ�J��fyʾE���1��=��<c9>:um�S��<J7�! r=�3�=v$>�5�>�?>��p>]*J>c*>$�9>fc����v뢿u.��/"G�e���E��w���m
��]���� g��~��߽��Ͻ�~���:�X�&�xL �+h�=`S?�"Q?�q?>?�Rv�S!">���2B�<��ߟ�=�A�>u�1?P�J?.o)?���==���id�j������ሾ��>D>��>�$�>�w�>Z%�:��C>��8>5�x> A�=Z�%=1V�:�J=�=W>̫>���>1��>�C<>@�>Gϴ��1��T�h�+w�e̽�?'���>�J��1���9������&j�=6b.?�{>���?пp����2H?���v)��+���>z�0?�cW?h�>E����T�d:>R��ͦj�a`>+ ��~l���)��%Q>Hl?j�f>�.u>;�3��`8�R�P�Yq��{|>�6?�䶾�/9�t�u��H�1Fݾ�0M>���>��F��m�����<��ei�c�{=�q:?��?Uy���氾��u��%���;R>��[>�=���=XM>)Jc�0�ƽ]H�L	.=���=��^>Z�?��->�"�=�բ>�u���+P���>B>>X+>�@?W,%?���&���Z��$�-���t>��>�n�>� >��J�1�=�[�>�hd>�p�d9����	���7�ҹU>�U��y)^��qj��x=�Q���B�=(Z�=�����59�}==�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾKh�>rx��Z�������u���#=Q��>�8H?�V����O�c>��v
?�?�^�੤���ȿ3|v����>T�?���?f�m��A���@����>9��?�gY?joi>�g۾T`Z����>ӻ@?�R?�>�9���'�}�?�޶?ӯ�?��G>��?�Yr?��>֒��t�.���������vq=�y>�p%�>>᰽���E�(r���̉�y�j�,G��m`>�1=���>4��E[��j�=㝽�˨��c���>��o>�nK>�>oA ?��>��>�=�F���傾� ���A\?v͕?�<T��Ȅ�Q�p<r玽�l���ȯ;b!?�}�>�y��H�>ןN?5��?��0?+5X=�7!��Ҝ���ɿ��佢Q2>ۃ?��>A�"=jy�>�XӾ����b�>���>�W�=y�ȾM����<@f�>��?�?[�x>J	?�n%?=^>�G�>�lG��Α�i?�w>�>���>�8	?فz?��?�H����/�0[��❣��J]�E�>N�s?
x?|t�>�����n���A5��\��$�ǽm�?ȃj?Qƽ�w	?ǥ�?��;?�FH?O�v>�K��5ؾ�tǽ�Ok>��!?(��}�A��J&�U��w?�P?Q��>�:���ս�ռ����j���?� \?�8&?��&a���¾!��<�*$��P��� <�yD���>ӡ>��O��=��>Sܰ=1m�`<6��Ce<�P�=ƀ�>��=}�6�؍��9,?	�F�Zԃ����=��r��yD��>�WL>�����^?;�=���{�����z���U����?���?Gl�?���#�h�O =?�?x?��>D��wq޾���aDw��px��m���>4��>I�l���ڑ����:E����Ž^�"�9��>3�>�	?���>��Z>$�> � �%�����D��d)Y����"n8�)5��:��M���:�d��hɺ���q�N�>D�Y�dM�>H? �>�lj>)�>����~�>\�b>䎆>��>�J>�>@��=��
��>۽�KR?����\�'�4��+����2B?�qd?�/�>�i�ɉ��;����?{��? s�?O<v>�~h��,+�6n?\>�>H���p
?S\:=��9�<�U��P���*�������>�C׽ :�1M�Dmf�j
?T/?�����̾U5׽XC����=�=�?��"?"�*���H��i`�`�Q�Q��'��'�Y��ڔ�E�\�l�m���ꆆ�����I�0���=B)?��?q���,�Y��׭p���9��V]>�j�>'�>��>�]>U���� �c}V��(��Ս�M �>��q?ɉ�>уI?d�;?�xP?]hL?;��>ll�>M4��Y�>�-�;��>��>�9?C�-?�10?�q?�h+?7c>6������$�ؾ�?˫?BJ?�?��?m䅾�vý#@��Zpf���y�����G��=�C�<w�׽=Hu��kT=�T>0?��-8��^���Np>��7?���>^d�>���M�~��0={�>�?C�>(����q��g��a�>�a�?�O��x =�F+>su�=+5��0���m�=�Ю�㲊=�ժ�vw/�%fK<y��=U2�=���}�?�Y5;�y�;�1�<���>b-?y١>n��<c����m�t�(�� �>Δ�>8��>٪1������e��=!��(�x�C��>W��?D��?g)b�ؐ8=�vj=&Q��!w��g�S�q��E.>[�>`+?�B?�,�?�^G?m�@?X^�=��@����������@���*?'",?>����ʾQ�Ј3���?�V?0:a����8)�(�¾<�Խ_�>�Z/��-~����D��s��
��<���Y��?Ϳ�?�A���6��s辑���0Z����C?�!�>�[�>��>��)���g� $�"1;>��>�R?�
�>W�<?z�q?c�f?+�w>]�-�0Ο�,֝�̮��Q@>U=C?�?K�?6xh?���>z-�=�1Q���:�澕P��V��������<��,>v��>ł�>�N�>Yً=s���x��Ei�r�=�0{>��>@1�>z��>|X�>1�#>��0?o�>l���!�&����׵�m���:!q?�{?.S�>��p�C->��lf����<p�>���?�w�?R'?k�����=q��<�<Ⱦ^�����>=�>�,�>����^+>)�>L�>Wv�>ә��Y���P������M?
	I?8<�6ǿOpq�~n�!���FE<�N���_��&���._�]��=�Ӕ����N��9�V�	R��}5��_Ե�����8�x�,?�>	�t=�d�=��=���<�D��w��<B�a=��<\�	= �j�w<�(����m���ƃ��Df<|�Z=��λ��ʾ��|?�I?�,?��C?�Ny>n�>!�@��P�>#�"p?ЃW>�M��a��I;��˨�5���N�ؾ�-׾�c������>�ML���>�&3>M�=1ʊ<���=��n=��=k����=�\�=4�=g�=N"�=4%>4O>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>d�7>TR>c�R��1��\��zb�x/Z�4x!?r9;��-̾^7�>pM�=�޾k�ƾ2�,=�(6>I/a=��F\�'ٙ=,�z�e<=�"m=���>��C>K
�=lr�����=y�G=!�=pP>J-���W7���,���2=q�=�b>]V&>g��>��?&V0?gcd?E�>.�m�r�ξ�o����>VF�=�]�>Bj�=rB>x��>o�7?��D?��K?�l�>�O�=��>W�>k�,�Ům��j�֬��g��<��?h��?լ�>{:M<!�A�č��6>��nĽ�?cU1?}{?�K�>����!ۿ����%�%��H4;�x�=}��+>���l'�F(ɽC
i����=\��>���>9�> �]>�5>C�N>"��>Pr�=m=0�="�k���=n�J����=Eq�<}H�<T���|:�^�<�1Z�ԉ�ƭ���v<��q=�<d5�=���>�>n��>�q�=糾[Q.>#���
L��C�=�O����A�0�c�J~��t/��t7�=UB>�X>�₽c ��2J?�Y>=�@>>�?9su?%&#>7��x־�[���Kb��~Q��L�=>?>GV=�R�;��a���N��%Ҿ6��>(ߎ>B�>h�l>�,�-!?�E�w=Z�?a5�]�>�{��Թ��#�K9q�`@�������i�5fպ\�D?�E��ҙ�=� ~?�I?���?ٌ�>e���ؾ]20>iL����=�
�I"q�ZW��&�?�'?���>�쾾�D��H̾T���޷>�@I�2�O���S�0�U��2ͷ�4��>������оk$3��g�������B��Lr�Y��>&�O?��?]:b��W��JUO����_(���q?�|g?/�>�J?�@?&��z�r���v�=�n?˳�?S=�?�>��=����q�>�?đ?3��?�kq?kـ�&�>7��<O>:u�� �>mJ>���=��=��>�@ ?��?�'������J�¹���f���h=�0>EG�>s��>g[M>r�n=�� �H5�=�>��>�n�>uɅ>;��>���>��
��S*��?ak�=C3>��??B�>k>�c�y�:D�/=���x5ͽ��,��*��.4=�9E����=4�<���>��ſ��?X��>��)�:�<?oe��>���>���=M��,Y>1�.>�".>���>R�W>'94>h��>a� >�Ҿ��>���Ab!�~C��hR��wѾ��y>M����n%�x�����S�H�oV��Pf���i�L(���3=�K��<k0�?����V�k�-�)�m��&v?l�>�06?�Ì��?��b�>��>���>�L������X����Kᾈ�?���?��>]Px>��?�#�>�j���G���`��<]�`r������k�ɚ��d�������.>�z}?N��?.I3?1晻���>%��?��=������>;�R�E�N���=��>�Le�k�a�ھ�������2>4��?/�?���>�
^��M�=l 3�`�>��P?��?��R?)�X?�%<��"�>�>��?�?Ո2?P�/?ʈ?kB�=�ɨ��3=G��>M輡�B�I_����ݽ��C=*�0>M��=�?�=M��=۟3��Z����O=10=���<������1''=�*/>X;H=j��>�]?���>sC>D�1?J�k��BI�^6��=5&?��"=�lھ�2žp㾴��pH�=��~?�d�?_c?!��=�H7�P�#���>7��>!>#�F>?�>����M��,>>I~>O�c>�q�=���H%о*
���O�w��=���=F��>�1|> ��,�'>6|���1z�ڣd>`�Q�̺��S�<�G���1��v��X�>��K?��?杙=�^�/���Hf��/)?�]<?�NM?��?�=E�۾��9��J��>�<�>kg�<L�������#��Q�:�|��:N�s>i0���ڠ�h^b>����y޾M�n��J�����BM=~~�0V=��վ8.�G��=�+
>����� ����Iת��0J?�j=Bz���eU�Ol����>t��>eܮ>N�:�k�v�|�@������<�=���>;>���Z���}G�9���>"`E?�4^?В�?1ȃ�Er�FB�3_ �$����!?٪>�?�<>�_�=�h���l�I�d�J`D�l��>k�>n(�3FI�Ĩ��e��,$��t�>/??@>|�?��T?nM?#Ea?_ )?U�?�>�?ɽQ���B&?7��?p�=1�Խ�T� 9�HF����>z�)?E�B����>K�?�?�&?�Q?�?<�>�� ��C@����>Y�>��W��b��S�_>��J?ۚ�>i=Y?�ԃ?��=>Z�5�ꢾm֩�V�=�>��2?�5#?K�?⯸>$?n7�����<?qZ?�
�?���?A�3>��|>���>"�?�m�>:j�>%7?"�?�!,?�X?�O*?�6�>�h�=��[��u����;QȌ=.��<g���8<��+=���@B�<�躻�Z���[��,�O<;%7�X��;;o�6>�_�>s�s>�����0>��ľ�L����@>�p���Q��V׊���:�<۷=҇�>��?^��>QU#�=���>�I�>D���6(?�?}?�R";�b���ھb�K���>e	B?���=v�l�.���'�u���g=J�m?��^?�W�C%��El^?�l?���D�Q�grȾ����R��߬?PE?��ɾg?<>"�l?Ζ_?��?S�f� ���Q⤿UU{�۞žr31>���>tC8�	ن�V�>�;?Ҁ�>���>4�=�о݅�����؉-?/ʣ?Y5�?ͺ�?!UX���h��1�I�����?cJ?�>�� ��?�Paľ�¾���R���˯��Ȏ�)u��d���E�9(%���ͽ�?n>�Q?*ł?�e�?��W?�X �=���N\m��7q���V��	������C��W}�|�e���fM��v���8.�=|y��@��k�?�)?�~"�){�>E�������о��I>�.?���=����B�@=��o=T�i��?/�*��|�?�>ً�>�;?�X�zFA�h'2��*8�����ec=>o��>���>�q�>�Eg<��+��콸yǾ����K9нa�w>�c?�K?#0n?M�����0��-��6D#��1I��.���5A>�u>�@�>�RT�3�ɻ%��4>��rs�y������F
�歏=&�3?�ހ>��>:/�?�d?�	����R�w��P0�!��<��>�>h?h�>t�>��Ƚ� ��#�>��X?�[�>s��>�ƴ�Z,�I�z�d󻡭�>�md>���>�d:=�0N�X�@ߐ�p����@��m�=k`?5�d�X�y���>H]J?�����> �>��)�Z]7�Ӂ��&=�U�>9�?�>N��=`��,��>F��{�Q�PO)?�<?nђ�1�*�P~>�0"?���>v>�>7%�?,�>Vþ*�7�@�?�^?�BJ?VUA? 7�>�)=Cñ��$ȽV�&���,=/��> [>X�m=1��=��$�\�8t�a�D=��=3%ϼר��Ԁ
<�崼SK<O��<�	4>��ֿOI����BS�2����-��r6���O��Ο���ӽ�"��.J��J�Tݽ��;TP��@��X��kx3� �?Q�?�o�����ˢ�J�����C��>���[����ۯ���I�����e�徘!���6,��&E��_�%@O�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�{A?��(� ���V=a��>��	?C�?>!R1�NO��T�>�7�?x��?ύM=)�W�n�	��ue?�h<�F�މݻj�=�I�=8�=��~_J>�H�>(���MA��ܽ}�4>��>�"�ƌ��}^��9�<��]>b�ս�8��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=����=�����մ�ݎ�=���=X�]=�([�Nϴ������8F�c :�a�8<���=܁>���>iV�>�f7>��c>�I?��|? _>�Ɩ=]��u<���~��Z=�F���P�F����[�鑾Z����ƾ��� `⾢���?��!=�c�=d6R�ܗ���� �O�b�C�F���.?�y$>��ʾi�M��-<�mʾ��������!إ�?,̾G�1�� n��̟?��A?������V�����`�T���®W?�U� ���쬾���=񳱼��=�#�>��=��Z 3�l|S�v0?*\?�k]���**>�� ���=��+?B�? �Z<�'�>	M%?��*�*7��a[>ˤ3>�֣>ط�>�=	>Z���S۽2�?��T?�������ڐ>�c����z�#a=�1>x75���G�[>�w�<����U�O���a�<["W?��>��)�P���f��Gy��<=r�x?�?*�>�gk?��B?eu�<hr��%�S�-��pw=��W?7&i?ǯ>�ׁ��о"[����5?(�e?�N>[h�8����.�O<�B*?��n?�b?>/���}��$�����ks6?��v?�r^�(s�������V�V<�>[�>M��>0�9�l�>[�>?#��G������Y4�$Þ?��@���?c�;<��B��=V;?\�>�O�`>ƾTx������M�q=)"�>>���3ev�����Q,�X�8?䠃?,��>Ó����;��=蓾,٫?=��?~���
@<�z�=�j�� ���^<)��=��&���0�ܴ��48���ʾlo	�@D���y�Ak�>S�@ymؽ-@�>�88���$�ͿEp���]о��m��h?O�>����:����l���v��xF�6�G�#����K�>�>A�������{�i�;��ݡ�r��>�4�~�>K=T��h��[۟��-<���>.��>H�>뭽彾J��?Q���7ο.���˨���X?�g�?Qn�?�d?��6<�w��y{�n�v%G?߁s?z#Z?·#�E]�C9�!�j?�_��qU`���4�yHE��U>�"3?�B�>W�-�I�|=�>���>g>�#/�x�Ŀ�ٶ�9���X��?��?�o�#��>r��?ts+?�i�8���[����*�!�+��<A?�2>���P�!�I0=�bҒ���
?R~0?{�e.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?J��>��?#I�={c�>z��=�毾�XL���>H�=Q��?˵L?R��>6��={�4�O�-���E�)�S�2�	���B��2�>5�e?I�O?��a>Q���#��� �r�ٽ��;�K�fs8�]E�(�콈82>�;>�>�<�^mҾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��?"���
���~�/8��>�GZ�=�6?2^쾨�~>�p�>yv�=��w�8���t�Ҷ>��?ܡ�?>�>��k?wBn�\B�Xy+=�o�>�'k?��?ũ��Si���>>L?L�����V��he?;�
@v@�a_?�u��p������۾66��nPt=p3�=��Z>:�=���=��b>���<ր7>y�>S3�>��>�nf>��>s�'>><�<�F~���!�����,��SPa����2�����t=5���n�нt�߾(n<��Y���ʽ@�νF��R�̽�hJ��:����2>�W?�H?��d?`&?��h���>ޯ4��	3��S��� =�J�>c2?�K?�� ?<r=<㮾Dt�r����髾���Z�?̧�>@;�>�5�>n0�>?��G�>�}=��c>DI>���=A붽4K\<_0:>�Z�>��?��>�X>d�D>]���u��:�c��o�A0���?����w`R�G
���������͎	>�7?�u�=���A�пfa���C?�����wB� '>�2?�T?u1 >__���k!�e�>f�%�܍Q��t>����j_,�r$� G>+?	?E�f>�0u>�3�d8�*�P�|y���Z|>6!6?�����H9�սu�!�H�Xݾk^M>�þ>��C�Xk�B���3��wi��^{=~�:?e�?�(��ް��u�DI��`,R>�\>�R=���=�RM>��c��ƽDH�چ.=#��=�^>�Q?�l)>U�=GG�>2Õ�ԔG����>�E>'N$>%�@?�+%?����.��肾��,��My>���>�>�>}6H��=��>Ρb>[C����������GD��W>��`�juY�9M�@�m=mꆽ>�=Z��=�U��>�?���%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�w�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?`�N>f�?�Ii?2��>����(�G秿(�����E=}���>=�==9����?������k��f�A�t��>qʷ=���>��I��t��?>�ط����N�$C�>]/@>�P>>��>��>h��>Qh>l�=��~���xE��rT?�ے?�d�'<��U;>%{a=������;R��>?7��g���G>�KV?�ы?E%U?ml�>;�?�2���Oʿ�D���k���q�> �0?O~?��j��s>�"�%�ؾ�>-��>Qߴ=��ξ���+%�_��>�9?���>ON>�?��'?�}>9�>^�D��<����F�n�>T��>[k?��p?w�?��ľ��6�
A�����'.V�o�>�;v?Un?j��>�����ќ��L=]½V���$hd?�Pn?�ѣ���>��?�S=?`�C?��{>��)ؾ"ܽ��3>��!?�����A�)T&�
��}?�K?���>E6���1ֽi+ؼ����c���?�-\?�<&?���.a��þ�e�<�"�[�\�H�;�[B���>��>s����_�=�)>�ɰ=�hm��76��8g<��=W��>���=�(7����{�+?�9�5���ړ=>�r�"E���z>�M>�C���[^?s�D�o�|�_��B���"�V��#�?���?r��?�����g���;?�[�?��?]��>�k���zݾx�ݾCx�ʒy����q>p��>r�/�Y��������񩄿=㼽S��r��>�@�>�K?���>'VO>A��>�����&����i� �^�*Q�g8��/�����8���9#���������z��>������>BF
?2i>�ay>�N�>:��dR�>5eT>;@>�w�>b�V>{4>l�>���;�н�KR?����!�'���辬���g3B?�qd?Q1�>�i�7��������?���?Qs�?<=v>�~h��,+�qn?�>�>=��Qq
?T:=(9��;�<V��j��;3��C�?��>�D׽� :��M�'nf�sj
?�/?�����̾�;׽�C��l��=6�?���>�c^�A�^�
�l�H,�P�n�,!��ʞ{������w?��}�h��� ����T�/�
��S>kc?�c�?(o��zi��"K@��L��[�*�\g�>\z�>�a ?�[�>�A>hm0��Kc�k�t�N��G����>�W?D��>'uI?��;?�jP?$sL?�ߎ> e�>0y��X��>oW�;/�>��>��9?��-?c/0?�p?�:+?��b>[?������ �ؾw5?M�?G<?�?��?YŅ�OĽ�?��	�h�s�y�� ��W|�=_�<3{׽�\u��uV=	�S>-q?Ǩ���8�#����k>ϥ7?���>���>���������</<�>��
?}�>;g���]r�m:��<�>J��?��i=�|)>���=҄��u��r)�=&̿��Ґ=I����V<��<✿=R̔=�4q��0��D�:�H�;:��<�`�>�)?C%�>�)7>�ѻ����9#��6>���>�p>R�,�-H'��?��������`��0�>�(�?.T�?�=�g�=��ڼ�-��-|����Ǿ�:��U�0=�?n6�>,?��?�hE?@aT?+��>��m���Gע�+����/?�!,?���>����ʾ�憎Ј3�b�?UV? >a�k��;)�}�¾�Խ_�>)Z/��-~����D����X��<�����?���?�A���6��t�J���^����C?u �>aZ�>�>��)�I�g��$��0;>���>�
R?$�>y�O?�<{?��[?iT>�8�71��ԙ�t3���!>�@?걁?��?Uy?�t�>B�>�)���0U�������n߂��W=�Z>���>%)�>�>��=�ȽZ��K�>��b�=l�b>Ӑ�>S��>0�>M�w>dF�<��B?���>n�������X���?���̻���f?s�?�-?n�A�I�'�:�S���	��˦>�+�?�?k:?�Z����=�˼����Fo��1�>3d�>��>k��=�3'=��=@�>�K�>�E�2���x,�������?&A?�H=ApƿM}�T�R�8���1Ð=�nu�۵*��e������ͻn�h��������iJ�����	9o�Dx������m��ȩ�>�DE=�>B�= =�L8��C=<7�$=6�n=���<d�m���r�$����i7��Ҋ;,�<"W]=��<A�˾��}?@;I?��+?�C?�y>�=>՗3���>1���F@?�V>r�P����ă;�˪��� ����ؾ�v׾��c�Nʟ��G>�lI���>�93>�L�=y��<4�=�2s=�ǎ==/R�+=�$�=�Q�=e�=��=��>U>�6w?X�������4Q��Z罤�:?�8�>e{�=��ƾq@?}�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>s��=v�2�T��>��J>���K��A����4�?��@��??�ዿТϿ6a/>%�7>�">q�R��1�N�\�y�b��{Z�l�!?bI;�{J̾�7�>��=n,߾"�ƾL�.=k�6>�cb=�h��V\�&�=��z�.�;=�l=$؉>v�C>�u�=R2����=`�I=W��=��O>�����7�H/,�g�3=���=!�b>�&>���>}�?b0?XWd?	7�>\n��Ͼ�=��`H�>3)�=�A�>�΅=�jB>���>4�7?��D?��K?+��>�=$�>��>6�,�۲m��l�2ͧ�㱬< ��?@͆?�Ѹ>��Q<!�A���\d>��*Ž�v?tT1?�k?vޞ>�>�M�ܿ�-��%����]�=<�T>ͯ�=^��<?���2��<ۘ�=6�l>0��>�
�>�"�>l��>���=IT�=`V�>�%'>V8(=$�6<�9>a�H=�>��ݠ�����k��6��u=s�<$X�;cz@=ߩ7�h><_�;=���=|��>�]>���>d��=�#��y�.>}����L�Y��=!x���EB�{<d��J~�{/��I6��B>��X>�	���&����?u�Y>l@> u�?�\u?A�>��a�վ7N��-<d�$�R�п�=�	>�.=���;���`��N� &Ҿnn�>C�>j�>�Sb>2,��)C���%=��ܾ�0���>F���r�S�m�$��wt��k��b7��t�f���
<�G?���R�=��z?�eG?fא?f%�>򭭽����K>Q��3&p<��ߪz�Vԉ���?Jb)?W��>vܾ�NE�B���V�<� �>x%��v\T��o���~N���=:�e�$s?E��g����%T��'��1񖿎.I�A�b�_��>�yl?�o�?���u"e���3�-$���tǽ��> �?�?�S�>��a>�N���~�q�X�` >^"�?6��?��?
�F=��=X#ȽDy�>P ?���?�'�?{ct?o	#�P�>C=��3>���E>��>�ܠ=f@>��?E�?�?m֊�T�1��9��bL����l�I=�Ȁ>Ze�>2h�>P�>_W�=�P�=ͭ~>�T�>�>W�`>\�>���>����Xa/��?���=p�>'�)?<��>5��=Ɍ�<Wd5���=���6��f����_O����=����=�ܽP��>P�4��?�=�վ��?a�<W���v�>4Γ=d'��dV>B�7>��N>J��>�o�>���={��>KH>�FӾ�>����d!��,C�Q�R���Ѿ`}z>�����	&�؟��w��uBI��n���g��j�L.��Q<=��ͽ<&H�?�����k�%�)�{���-�?�[�>�6?~ڌ�����>��>�Ǎ>�J��h���Xȍ��gᾋ�?/��?<g>V!�>5Gg?P��>2h8�/߾��r��7s�na��"&���t�����?���	�.�O�g���M?�x?Q�c?�=��l>,�l?���g�����S>2��������б>}�ɾZ����z����ҾL�ӽ �J> Ӏ?��?O�8?��⾜,�=��Ѽ�;?�D?Q�s?��P?��Q?~�<n�>@�>��
?P?�1?�e?�M?r�>��_<f6=�#>��лf��-���_S1���H���k>��z>���>�q�<��G>���=���Ň��?= �UAf=9�=؎�=��>9�<>�M�>jG`?ح?%�4>�u?�z��^�@�GĬ��nA?��=ξ�zӾ�U�j��>l3=��t?/�?��t?4.>g�5��;;����=��>f�=�|>G��>�>��C���<>��=?P2>���=�����F�>"羪�T�	0;TI�=��>Cm}>����yn'>7W����y��c>W�U�#��L�T���G�u1��Nu�J��>��K?��?���=0N꾿3��ef�S�(?	=?��M?�z?iӔ=�ھ��9��J�7���>U�<w�����:롿h�:�8q�:�t>c'���ݠ�kYb>`��Hu޾%�n��J���羶CM=���TV=����վi5����=%
≯��2� �-���֪�1J?{�j=7x���_U�p��.�>���>�߮>��:���v��@������6�=O��> ;>wZ������~G��8��@�>$FE?oW_?Xl�?�	����r��B�%���4U���jȼ��?Db�>?b?WB>���=������d�fG���>o��>&����G��#���-����$�Ku�>8>?��>"�?��R?��
?�`?�*?iF?>6�>G��F޸�B&?���?^�=��ԽL�T��9��F����>x�)?,�B�Ѷ�>��?��?�&?�Q?��?��>b� �nB@����>�Y�>��W��b���_>��J?+��>�<Y?�ԃ?>�=>K�5��ꢾ�ԩ�fZ�=>|�2?:5#?��?T��>�'�>������w=C�>��l?s}?��m?�٥>�?��d>`?H�>g��>��>��>�]#?�Hj?��;?�g�>&�<�v�hy��.������<�����s�=���v���~%�{�<#9>���=|#� �<a2S< w�<~?�;��>Bau>&�n2*>��ž�����x9>�f���>��1!���@�/P�=�X|>H	?	�>d��κ�=�_�>ɽ�>$`��d(?�?��?��;�a��hپ:jI��`�>gB??	�= $l��͔��x�9�M=��l?E�^?b!V�hY��mWh?�{?���']S�����؆���ž`�?W��>q6����>�7d?
[?h��>�)ʾ.(���Ӫ�}�r��Ή�>s�<]h�>(�d</�y��>? ̴>���>���=�I��g`�����i?~Z�?jڸ?�ֈ?dQB>�^���O�@�/З��T]?X��>5(%���F?�÷�aİ���0��x���[���%1�����`x�߽��g�$?���= 4?X�~?�A�?�,T?��%�d�����H���Kr�I��M&�p/|�_�3�%� ��pC��^	�l�ᾈ&-�:|X=�^�J�A��h�?��'?�2�G��>����<l�I;̾L\B>�#���M�7D�=�B��A�A=�]=w�g��.�Q=��\c ?��>��>��<?�M\�(>�w:2���7��.���P2>衢>�I�>�+�>&�:�,���꽜�ɾ�@��4cӽ�u�>�g?�#V?Y"l?�l:���'�p t��~9���L��G��v�j>�^6>�Ld>�����W�W+�sP��hn��"��|��[N�>j�4?A�>�;�>�J�?ej?:��;l�������=�w��LÍ>cL?��>@Bv>��=���dA�>Im?��>>�>���V+!�6c{�
�ս"g�>�ʮ>��>Y�o>}\,��[�l ��|*��N�:��N�=T#i?4���mC]�ك>�<P?��4��j<��>�j�lT#�[��� '���>r)	?���=�R>>iƾU\���}�e���TO)?�H?>咾/�*�7C~>%"?փ�>W5�>�0�?,�>�gþhu2�8�?&�^?�>J?�OA?4J�>)�=K𱽀7Ƚg�&�M�,=鄇>M�Z>�3m=�t�=����p\�4y���D=�w�=�zμ�M��z�<�f����J<��<�3><mۿJCK���پ�
���t>
�u戾�����b������`��P��Vx����O�&�PV�5c������l����?f=�?e���A/��̲��ؔ������K��>�q��������&+����r����c!�\�O��&i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�|A?��(�[��CV=���>$�	?��?>�R1�DI�>����T�>m<�?���?wyM=O�W���	��e?~<��F���ݻ��=�:�=�E=%��%�J>�T�>����SA�AܽQ�4>Iڅ>%}"�H����^�3��<�]>I�ս*;��ī?�$\��e��	0��G��e>� T?�j�>��=d�+?��H�0�Ͽ��\�նa?>�?��?�(?\����m�>�ܾ(vM?��5?��>�n&�z9t����=}Rڼ˭��F��_�U�<��=cP�>�>�!-�5�� O�������=�� �!�ÿZ=�x��k+��/��=G\=�������J=#�^���-�����?b<�1�=@�@>艜>t�x>iu�>��\?�_?:�Q>P�8>垶�n�a����;{�K,���b���?���h�������Q�O߾AL�����W��� =���=�6R�y���3� �V�b�^�F���.?v$>��ʾ��M��-<�pʾ�����ф��ޥ��-̾ۗ1��!n�J͟?~�A?������V�f���R� ���1�W?BO���tꬾU��=�����=�$�>芢=V�⾴ 3��~S��u0?H[?ʄ���Z���/*>k� ���=��+?��?�Z<)�>RN%?��*�<佊_[>��3>�ף>���>)?	>���pW۽��?P�T?w������Iِ>�a����z��a=�0>�75������[>�z�<�{�U��J���^�<��W?P��>�*��*�Rd����6��W=ǘq?�?`v�>j?�R@?���<L��K#X��@�9=?�W?�6j?$�>C)a��XѾ�����=0?��d?��h>�`�����0�bl����?X�r?�)?��m�^~�t��3��4?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?r�;<��U��=�;?l\�> �O��>ƾ�z������3�q=�"�>���ev����R,�f�8?ݠ�?���>��������=�?
a�?Ax��]��<r��l�j��8 �==<x��=k�;�/Y/����G5�9�þ�E	�4��+���G��>"�@T�̽@��>I*��\保 п������پ��b�?���>:\ܽ���t�e� �p�ۇD�O�G����\k�>f�>����H7����{�U�;��ʩ�3��>�'���>q�T����n����G<׉�>�8�>�چ>2j������r��?�����9ο'ў��[HX?0P�?�_�?�8?��:<��w���{�q��#^G?w�s?�?Z?�t&�\]^�=�4�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�/�S?�F����A<��eւ�����S���ި���F.����ױ���v�]�?I�@�5�?s����B7���R?�y�>����KU��X߈>���>s>�e�xd>~����!�\��<X �?���?ܭ?dN��a���z/>W[?��>!f�?�o�:��>C*�=�"޾�'�?�ֽ�+=z����#�>CEC?��?5';=\8���4�+[m��*��٠m�g�*���(=Hs�?��g?7c>��n��v�T�.������b��V7=�<�<��c���@��>b�f>�y�=���������?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6��+���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>F�Խ����Z�����7>0�B?[��D��t�o�z�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?sQo���h�B>��?"������L��f?�
@u@a�^?*�!׿���Ծ���^P=ǉ=K��>��=D+�>��I>4��<�]>��>���>^n>^R>��>Qy>��>!p��a�&�����婒��K���.��푎=U�ž�,��A�4���Z{�E�C�&�	��d�<>��6Iؽ�2N=��=BIW?�6S?1{n?5��>�����=>F\���<�"�㺣=�e�>��/?�D?�"?�S=Js��[Ah�����Dd��G
��T��>!�X>n��>�d�>3۬>�����M>�jA>��t>o��=��;�/_���=[�E>�T�>��>�K�>�C<>��>Fϴ��1��j�h��
w�v̽0�?����S�J��1���9��Ӧ���h�=Gb.?|>���?пf����2H?%���y)��+���>|�0?�cW?�>��s�T�3:>8����j�3`>�+ �zl���)��%Q>ul?w�f>/ju>ǥ3��i8���P�A���g7|>8'6?Wݶ��Q9���u���H��Kݾ�cM>o��>�F�.u�� ������i��{=�t:?
�?����ٰ�w�u�K��bVR>X9\>�<=���=�aM>�c�k�ƽ��G�1�.=�r�=�k^>V?u�*>ޖ=m�>V���mM�/��>��E>T�.>4@?�:%?�������:��4/�ޭq>J��>���>]H>��H����=2��>��_>�������J�D>�!Y>?}���_�e#f�Tq=W훽+��=���=�� ���<�S#=L�~?~p��_ۈ��P뾨���}LD?%�?�b�= 3><��"����|��	��?��@[w�?�\	��V���?�C�?8�����=#O�>���>q'ξ�8L�Ф?��Žv���Β	�>#��G�?���??�1� ǋ�%l��6>I_%?V�Ӿsh�>�w�}Z�������u���#=��>�8H?~V��V�O�>��v
?�?�^�멤���ȿL|v����>S�?���?A�m��A���@�L��>-��?�gY?�oi>*h۾�`Z���>��@?�R?F�>�9�Ϗ'�0�?�޶?ǯ�?)I>u��?/�s?�|�>R�w�\K/��*��d���
O=��X;Gr�>�G>s���2]F� Փ��e���j�P����a>5l$=��>�K��#��ON�=�����K����f��>�6q>�I>�[�>y� ?�J�>ˬ�>��=&7��8Ӏ�6���ٕL?g��?���k:n�6��<^�S=w�g���>>1?������ƾj�>��Y?`	}?;�O?Ox>����2������d᷾�<�S>�T ?�;�>ڤ��Y�>��پ�2�_�>�/�>���w�̾����q�<"��>s�?�~�>�KG=F�*?�5?}N>PI>[�I�f�����F� �e>�t�>C�?��m?��>�P¾p1�ߟ�ì��'�g��h�>�<}?>�?�Z�>�%��S]���]��˙�<�">J�r?b;?��7�,SB?���?��b?g"V?cL>����6�g�����>�"?c�,�@�8r(����K?��?���>oA��m�����ؙ��@U?�<^?o�'?�Y���_�o����<��컢���z<`���&!>o�>;~��:�=O�>�?�=��k�=�6���;�X�=�l�>^��=[�2�趛�2=,?ѺG�wۃ���=m�r�MxD� �>8IL>�����^?9m=��{�����x��	U� �?��?]k�?���*�h��$=?�?=	?]"�>�J���}޾#��qPw�<}x�nw���>���>�l��W���ʙ��vF����Žs��ud�>���>�(?R ?L�U>���>k���qv%�u�� ���\��Q���5�[1/���h���e$�T�}���eE~�~�>.���	�>0�?�cd>Q}>'��>��M�(>�><�Q>켃>I|�>[[>�8>Hn>�>G<�A���KR?�����'���ϲ��83B?�qd?1�>Yi�J�����H�?���?is�?�=v>�~h��,+�sn?�>�><��Vq
?S:=e/��8�<�U�����k2������>�D׽� :��M��nf�Uj
?�/?:����̾�<׽ӊ���	o=N�?�(?��)�2�Q��o�d�W�~S�����3h��h����$�ěp��쏿�^��A%��֡(��`*=��*?h�?���� ��m%k��?�Tef>��>�#�>�޾>xpI>r�	�C�1��^��L'�ƹ��U�>b[{?Ĉ�>��I?<?|P?mL?�>�f�>2��|j�>��;�>[�>g�9?��-?�+0?�n?�h+?�c>&x�������}ؾ�?	�?XJ?�?b�?qޅ��hý�b��V�g���y�2c����=���<�׽�t�T�T=T>�M?l���[8�����Zl>h�7?���>�i�>�V��<���<��<���>2�
?��>R����Hr�~��C�>ℂ?d�u�=�o)>ur�=�����.����=�Yɼӌ�=���f;��� <d!�=f��=��t���b��٠:�};�u�<�?o�/?vs?>cR4>�xB�?���^)�*
����>�t>��,�s%�����\G���ur�2�[>%/�?���?F��>>dV>>���@�
�\��R[�?�>k�?;��>�K�?���?�H?�/I?��g>��g�h;���ʠ��J���V?{!,?B��>n���ʾ$�ĉ3���?nX?y:a�ͷ�G9)�w�¾��Խ_�>W[/��.~����MD�[��������ɜ�?&��?�A���6�ew辀����]����C?"�>�^�>��>U�)���g�<"��0;>/��>
R?'H�>g-P?aL{?�[?�GU>�p8��ѭ������;�`:!>@?<��?⏎?�w?���>�>x�-��������� ��v���뀾lYa=�7[>��>�:�>�n�>���=�FƽDѱ���A�bU�=91`>��>3ˤ>]R�>Z}>R�<�G?��>���y ��%��������Y�]4?��?H��>�pa���1��Ux�8C�j�>�%�?0��?g#?������=�l�;�A��`�����>�w>�0�> aT�{"{>o �>qq>N��>:=�g�B���k�g/�cp5?��X?؉���ÿ͙s�*��k$��x@���6e��(����PG~��o�=
X���'�jw���j�1O��ȉ������菾�-���>���=�R
>Ͷ�=��=*�:�U[:��=�A2��<̻='��.'�<*�׼�3 <����y�I��9�<X��=t:1�G��C�9?��m?�)R?ur9?$�>�Hx>&�W�JH�=H� �&?%C(>�Q ��F������ƙ�,��A��]��T<�-}��V/�<�d��}�=��a>�o�>��&>��U=���=6��=�����=�8>'
�=�R�=n�.>N��=X�S>�6w?N��������4Q��Z�v�:?�8�>u{�=��ƾ>@?�>>�2������Yb�
.?���?�T�?'�?ti��d�>%��#䎽Yp�= ����=2>���=W�2�:��>��J>���K��3����4�?��@��??�ዿѢϿka/>�77>��>��R�ׄ1���\���b��IZ�8�!?]6;�$̾A<�>�	�=�*߾��ƾŇ.=��6>�*c=#	�,6\�3��=��z��s==l=C��>�D>w@�=����x�=�KH=�h�=�O>B�����7���+��05=s��=�ob>��%>��>��?z^0?wLd?s.�>�n�[(Ͼ�C��9�>���=�3�>͢�=�dB>^��>O�7?�D?�K?���>}�=��>e�>��,���m�@n�;§�B��<���?AΆ?�͸>��Q<��A����:l>��HŽ�r?�Q1?�k?^֞>B)��eiǿ9�k�a��	�@�\)>�ٴ>�>+�G��{J>j$��D�=�m�> �>�=`>q s>*#�>a�>*�>�U�>��C>W�W=A����<�\�</�ܽ���=Th�_5=s`�;��ཛ|뽛���S�<��y=N� =�~�=�Iv����=��>}<>ܬ�>Q��=���D/>߸���L����=�G��e,B��4d��I~�N/��V6�z�B>';X>�}��@4����?Y�Y>�l?>���?XAu?6�>� ���վ�Q���Ce�7VS�G˸==�>��<��z;��Z`�|�M�_|Ҿ���>�ߎ>7�>b�l>�,�*#?�^�w= �>b5�E�>L|����)��9q�@�� ����i�#�Һ��D?~F�����=3"~?�I?B�?��>���,�ؾ�:0>�H����=T�*q��h����?'?���>}쾅�D��H̾J���޷>�@I�2�O���U�0�)��0ͷ�5��>������оl$3��g��������B��Lr�\��>%�O?��?a:b��W��JUO����[(���q?�|g?.�>�J?�@?&��z�r���v�=�n?˳�?T=�?y>S{�=z����>�?~�?Y��?lYt?����>p�L=�vS>p�����=��=F#o=g!�=_?@?��	?p���pl
��m��l��b@b�O��<Lڟ=T��>���>i~h>MP�=�
�=�V�=F
I>卙>�ʚ>�h�>ޛ�>�K�>��׾�%����>��=��>�G?���>,�=>�u+=���<���f��"�b��E���o��>v�=YF�=҆ż�g?r⽿7`�?���>-�L��I?3�U�]�@�>�����J޽F9�>��1>��4>]c�>Y]v>`��=��>�T=�FӾl>����d!��,C�Z�R���Ѿl}z>�����	&����w��\BI��n��xg��j�Q.��Y<=�˽<,H�?�����k��)�����V�?�[�>�6?�ڌ�����>���>�Ǎ>�J��i���Zȍ�hᾨ�?E��?y��>�3o>fv}?j` ?$���]`����x���a��@]������:b����)=��w�˾�D�=��c?4�h?Kj7?ua�<R�>;�?n ��O��"?�B��1�S�E4�=��ʹ�^�/F�O^�(V���[>Vl�>a��?�2s?&�>�ý��>	�E=4�!?��]?��?fa-?)Q?��H>Ȳ?���>�p"?-X?H�2?gs�>�y1>������=���=DQR>Tf���!��'��A��
,*=	m�<��=AJ=��=���=y�;6�>f&�<�PZ��s�=8B�<�=�r=*s�=�!�>��]?��>��>6s6?aP0��-;�M�����1?,�=~�������;��{����?>��l?Ԡ�?`�Z?>F>)4>�9�=��v>�>�l+>ekU>5�>���<�2����=��>ȣ(>�˭=ߡ���
�����e����N=Z�>��	?u�> pŽ�)��7;�j�����9훾���������u���m��ξq�?��|?[K?Mv�=E�����=8>�V�+?pF?XÅ?�*T?\ѭ=R����d�Ә����p�u>Y�G=�86��/ƿMᨿ{~!���Y>�k�>Б�Oܠ�]b>̾�Yw޾l�n�YJ�:���+M=}��+CV=R���վ7�l��=�(
>����� �r���ժ�`0J?E�j=w��s`U�qo��R�>���>�ۮ>��:���v��@�����*�=;��>6;>�G����~G��8��A�>mNE?�]_?Rk�?����s���B������i��Q�Ǽ��?�v�>lg?��A>(��=����d��G��>���>�����G�76���&����$�㠊>#9?��>*�?�R?��
?��`?T*?6@?m*�> ͷ�0긾f;&?z��?r�=�׽~�T��)9�	/F�f��>�)?+�C��9�>�1?p?{'?r�Q?^�?i>|� ��?��}�>��>��W�W����_>�J?��>p�X?|̓?$?>�E5�	9��%ɪ�t��=,>z�2?�$#?��?悸>��>,���m~�:�d�>Bg[?�v?�H�?�Fk>�R�>,��>(T?�A>��>���>�b?$�'?*�W?VD?T�>\��<|9�L^������K*���q<�)=�?=�Vv�(�ǽW������<�N=&6=��<�D��f�D�ޅ�F�a<Q`�>yt>/��N�0>��ľ~`��~�@>��d���犾�:��U�=}e�>5	?H˕>S#�pݒ=Α�><T�>,���5(?��?Q?�;9�b���ھ �K��"�>�B?���=��l������u���g=X�m?�^?�W�1!���K\?(�t?��"�Q?��ݾ$��op����-?��?,,����*>W�o?-҂?��>�4��	������Gw_��Ď�� �=�Q>+�'�=�l�>١1?2�U>�I>>�j<��Ѿrh��ol�ϛ?��?��?yʌ?\?�=;�x����ݾO���_�f?���>����%G?�
�"=5��|�I�������h��G&��5��59����3��+��D��Yb�=��5?�o|?G�?уL?��=���y�D���g�y�=J�������.��ct�=>M��>�tXA�:���������Ee
���~�v�A�W�?G�'?Pd2���>���G��9̾�B>�������=�X����?=�9Y=�g��`.�����m ?]�>��>g�<?�U\��@>��A2���7������2>�>�A�>��>���:ɼ,��p�1�Ⱦx��ֈԽ�҂>*�]?K Y?��o?㴡�8�%�(~�q�+�+���j��hE_>��>W��>�0w���=�O�'��hI�bn�͖��ʊ����/�3=�R0?�~>�њ>�ݕ?��?����:��AU`� &1��븼�D�>��[?�9�>G��>����{�^p�>}uo? "�>�
�><Z��XV#��z�c���ŭ�>Yq�>���>��h>��*��Ra�`ꐿ�~���\;� 3>l?�逾~{U��z~>ޓI?"Jb�t��:3�>C�8� A��W��M��-<>T�?e�=��#>�p˾%���}��;���N)?Z=?�쒾3�*��L~>�"?���>p>�>�(�?�5�>!Hþ+��y�?E�^?�8J?xDA?�:�>Ng=����k3Ƚ�&���,=t�>��Z>��l=L!�=5��W\����4�D=���=��̼�帽�`<Ʀ����J<���<{4>�lۿ�CK���پ�
���=
��爾S����`������_��f���Vx�߉��'�V��4c�"���Ŷl���?�<�?|��!.��Q���K��������>M�q�֜�x���"���)���������c!��O�p%i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���z¤<���?0�@-yA?��(����u;W=��>��	?p@>=Y1��K�Q�T]�>y7�?���?�<M=��W�l4
��pe?��<s�F��ݻ`��=�=�=[����J>�e�>-c�#JA��ܽ��4>��>rW"�7��'t^���<��]>��ս*����y?����U�z-R���~�\lr;	~&?�r;>jļ�R?�[Z���տݺ���Ha?9��?ui�?|}(?l�����>���raB?��-?�V�>8}+�KP�AT&>X�<�dL>a��ͱI����=��t>M�󚃾��񾳲�x

;}�1=D���ƿ��$��q�)9=2�+�S�}��x���5�M����?gm����Zi=�C�=`�P>�x�>�5W>e�Z>�ZW?��k?+w�>:U>佝q���:ξ��&��m�����l���s�)����U��߾�R	�{���}rʾ� =���=7R�x���=� ���b�b�F���.?>v$>��ʾ��M���-<�pʾ򿪾3Մ�]ߥ��-̾(�1��!n�]͟?��A?������V�B��GV�R���*�W?�O����]ꬾ��=����e�=%�>ꊢ=}��� 3�t~S��r0?�@?���p��]i*>.� �Y9=U�+?8|?��]<�K�>
S%?��*�����\[>p3>���>z��>m	>1���ڽ�?�jT?��|�����>/����z��`=��>E�4�x���\><��ǈV����ۑ�<Q�V?D6�>��)����ߐ��c\-���*=��u?�d?T[�>�j?�A?��<	�����T�f����f=�X?��i?d�>�w�@�Ͼ)�����3?H
d?^<V>y�g�	��`�.��e��?(:p?�F?�Lȼ/~��'���z���6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=啾h`�?��?����_ih<D �'
l������<���=����r"�����7���ƾ��
����^Z����>�[@���4�>�<8�EB��QϿy��$�о��q�Z�?TG�>�Mɽv���!�j�&4u���G�y�H�j����ã>*%>I���y��X|��Q=���企��>4�{�>޳]�l�������;�<ޗ>��>�n�>���"ﺾ��?2����ο^��_�ejV?�˞?cރ?�
?83<r�x��={���@�x�G?�%t?6�Z?n�5��d�@"�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.��M?CQ���:���Z���:������о�� �ľ�b*�]m��MQ�����d��?J�@��?W6M�g�K��;?���>8�mn1�Ł��ɀ?X�>�>�c��2w>@W��\:��P�<�i�?���?:�?�S��_��cF���}?�A�>Q�?�|6>C�>��=�ƾg�5�ɫܽYl�˶ǽZ�?ʵM?n�?�4=��5��'T`�ۀ��4w`���+�.�[=�?	W|?�[�>}�2=%9ü^�%�>t��a�T;N>�轤�뽠�m���!>$G>��>_��qɾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?xQo���i�B>��?"������L��f?�
@u@a�^?*ֿGڟ�v��P���G>�#>׆�>�#�=�|}>"�=�q0=��i=���=���>��5>_j`>�>BV]>��x>���{!"��E��i~���J/��&��{>׾��Uw���X�]�Ծ����_夾�邽Jp���*6�$(���)�D�����>��S?�YZ?�
o?���>s^��>k
�W0:�A�����=���>�c2?�A?ʴ?��Y=�믾k�e���������ύ��C�>^$h>���>'��>sW�>�#S�)�E>t�E>Q~p>q{�=K��<\�����<��6>�+�>�z�>�I�>�C<>�>?ϴ��1��V�h�w�b̽�?Á��k�J��1���9��醴�Cj�=^b.?�|>���?пM����2H?����w)��+���>��0?�cW?��>��m�T��:>�����j�V`>j+ �Il���)�k%Q>Vl?+�f>��u>ǘ3�R�8���P�������{>��5?2��@�9���u�x�H�z�ݾM�M>"%�>d6�_L�3���~��Zi�ME|=fk:?]�?ʵ��l����Fu��3����R> �\>��=)*�=��L>�e��ǽ��G��.=̓�=Ij^>�b?�d$>!�=���>5p��xmG�}'�>nL>�C*>�!@?J<&?�׼}���⁾��,�:�o>Uz�>�>�X	>P,H�BX�=�2�>- [><��3w����%B���V>B߂�nN^���g��Q�=u函�t�=ב=���n�9��*:=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾRh�>bx��Z�������u�'�#=K��>�8H?�V����O�a>��v
?�?�^�ᩤ���ȿ7|v����>W�?���?d�m��A���@����>7��?�gY?�oi>�g۾M`Z����>׻@?�R?�>�9�~�'��?�޶?ѯ�?��I>	f�?{/t?�
�>�q��.����،���u=V�~;�̐>|D>R����iF�ֽ���M���!k����]>+)#=c�>Z佚����=�o��-g��nb^��Ϸ>��p>[�H>Tϛ>'Q ?_��>�/�>hz=�����W����p�K?`��?���`:j���T<�"=`:����>X�(?AD��Ҿbx�>]�_?��w?�NB?a�h>0e ������¿�孾��O��>�>�T?�]�>��B��+(>3�����>9 �>$����Έy��!~=E�>�u?!�>���<��!?�A;?��>m�v>6DB��3���2@�	�K>~��>��?@�h?��?� ����R��Ҝ�Y���0�i�ɾ�>��?�?0H�>����q���!��m�ҽaH�=ݜ�?�	Q?�v��c�>�K�?c�v?D?(��=N*>�>�mB��\�>X�?WjA<A�A�m�R�{�(�⶛>���>��\>ב��n-{�1�8�"I���%��79?� �?��O?��¾��s�GT� �<�
�=����,<VѶ����>�{v>��ýe�`>K��>��>g���d)���3���щ=�v~>��=y�3�R����<,?^!G��܃���=��r�FyD�M�>�EL>]����^?�z=�E�{����}y��{U�� �?��?,k�?��ڜh�d"=?�?�
?�$�>xI����޾ْ��Kw�frx�u�J�>i��>"5m���Q�������D��o�Ž������>�6�>Px?�� ?�KV>��>�n��X�&��|�4���Z�Y��	�t9���.�u���禾���6�S�ot�������>��c�>?	Dr>�{�>���>�vI���>hQ>��u>�Ҡ>v�S>Ā<>Ҹ	>�"�<��Ľ�KR?�����'����(���3B?�qd?g1�>[i�ǉ��G����?z��?s�?�;v>�~h�u,+�Yn?>�>���p
?	R:=�1�=2�<V�����,��
����>#B׽j :�LM�mf�gj
?o/?m��p�̾%8׽�p���o=V�?��(?��)�=�Q�&�o�<�W�S�VE���g�<N����$�Z�p��鏿�[��^*����(��(=J|*?�?3���q�~��0k�?��f>i�>v�>oɾ>�I>��	�0�1���]�XJ'�Y����a�>f`{?���>GlI?��;? �P?IlL?�ڎ>�{�>)���/�>r#�;K�>L�>��9?#�-?�0?�[?RX+?�Nc>bA�������gؾ��?s�?�G?��?��?g���*Ľm*��3�k�,y�!���L�=��<�
ؽp�s���S=��S>�?�: �Ӊ6�43Ծ�R{>T�2?�R�>W�>�Ƈ���I�P��=� �>��?� �>~��j��I�ճ�>4�?����^>=�Q,>���=ל|����y�=éf�LN�=&�=��B�F�<)$�=�=o�p<���:\�ûy3D<�=�?��;?�B�=�P:>1�n����xP5�����{ǵ>��>�'���������쯿�!n��m�=}��?O��?�>[�>�t�=����wx���%޾3v����=δ�>���>a�\?fr�?'u?�M>?�L�=zJ��n��$��B�1�E�B?�!,?��>q��%�ʾ�憎��3�q�?>V?�;a����8)�,�¾��Խ�>X[/�I-~����wD��!�����m���Ӝ�?���?+A���6��v辧���`����C?*�>�Y�>g�>��)���g�i!�6;>'��>BR?�|�>!J?���?�^?��{>�T ��e��裿��Խ�+>��>?v�y?ʼ�?��P?J:�>�i�=S�����+���F��H!��l����=nrx>"L�>�/�>��>U�>�g��g��SЈ�/z�<�*/>+t�>e{>=z�>5�>�o>N;?؉'?=<¾�A%���l,޾?LS���?�˃?@�>�����*U�3�������x�>(��?fr�?� �>�,�	Ǫ=��_����
�>��>*�}>s@�=��:>���>�!>��d>I�>]�M>C�_�ė��e���V�<?牄?�4׽�ƿ�q�0"r��/����|<O����j`��ȍ�՘U�/�=���������X�����������E��u�{����>⥆=Y��=��=6��<�Ƽ�%�<%=P=I�<};=
�j�,j<;���Ȼ��-�<��sP<��I=-���',�E�4?�Vj?}ZI?�}5?mo�>���=��H�=��L��5?�k>��<�	������b�����6XO�i�ch>�X̾��j�����ؠ=��>y�>R��>�I>�*����=|O�?�d�o:�=9��=R�'>F�e>VY�>���>�6w?,���˲���4Q��\��:?�7�>�z�=H�ƾ�@?|�>>�2������b�5.?���?�T�?��?{si��d�>v���玽4m�=)����<2>���=f�2�O��>��J>����J��ׁ���4�?��@Ǟ??�ዿӢϿ|b/>�7>�)>�R�B�1��\���b�h|Z�:�!?�I;��J̾R3�>,�=t0߾r�ƾ��.=��6>mb=p��Q\���=��z�*�;=�	l=�Ӊ>-�C>&��=�6�����=��I=���=��O>�#��Y�7��,,���3=���=��b>c&>��>;�?]0?�Qd?�5�>Sn�2Ͼ;A��39�>��=�>�>پ�=|]B>��>��7?*�D?r�K?&|�>	ˉ=��> �>ř,��m��m�I§�5	�<���?`Ά?ݸ>��R<�A���_e>��+Ž�s?P1?Cj?��>g�1����$�r
�ٰ�=<��>���>��W>B4�>�F�>2㼳�x=�G&>�x�>f��>h�*>9�#>��^>i�=~}�>�mF>�nF=�j=�5/��/=YNW���;M���0s=9���ۣ�9�޼(�u�r}�p~���K�8���bGѽ��=��>�<>��>{��=���D/>߸���L����=�G��],B��4d��I~�L/��V6�p�B>0;X>�}��<4����?@�Y>�l?>���?OAu?Y�>� ���վ�Q�� De�VS�\˸=B�>��<��z;��Z`�z�M�_|Ҿ���>�ߎ>��>�l>�,�7#?���w=�8b5� �>�|������'��9q�@�������i�vӺA�D?vF��ě�=X"~?��I?>�?��>���Æؾd:0>�H���=-�:*q�oh����?'?���>�쾥�D�cH̾$��߷>5@I��O���J�0�$��:ͷ�,��>������оW$3��g�������B�@Mr�R��>��O?��?�:b��W��9UO�����'���q?�|g?1�>�J?�@?�%��z�r���v�=�n?³�?O=�?t>�q>������>1>!?�~�??��|?m��K2�>�k"=�gV>Y�`<H�>� 	>���<>sy=��?��?}/�>�]���%�^���A�оK�v��Nȼ��=��>Z��>g��>V��=?�=�\U=ӑh>Mk�>,x�>��;>��>�G�>!ƾR�$�"�?��=��D>��F?��w>��]>%�7=!8�=J�=M����׵�C�˽Ǌq<2�<���<������?������?ԃ�>1VN��*?N,C��=ђ�>���<�����r>d*>�U�>���>�7�>)�Y>�g>Ď:>�FӾh>����d!��,C�Y�R���Ѿk}z>�����	&����w��OBI��n��xg��j�Q.��X<=�˽<,H�?�����k��)����R�?�[�>�6?ڌ������>���>�Ǎ>�J��i���Zȍ�hᾥ�?F��?X1�>=[>�֌?��>S"��0���gz���9��v����0�g��y��S���xپ}�=��\?�T�?��6?YO��Ë>"��?�,�+.	����>����k1�ZO8����ON1�+��N��Y��lR��,�?C�?8xZ?s�>�r���tc>��{�p{�>�b?��i?s#?H�]?�/L=�ݧ>
��>�?�\,?��,?{� ?M�`>a������=K�>z��>JT���8����sھ�S[�=%�(=Z^>��.���L<��=u���G��=�C,=��=�8<5A�<|�0>�ԫ��*�=��>~�]?�%�>I��>h-7?͋��8�F����q.?�	0=f5���ό�f:��O�y�>tbk?M��?@�Y?Ie>v�A�1HB��n>���>�"&>`�\>N%�>LA�4#C�;]�=>;�>�ڤ=\�U�b���	����a��<�g>3�>�J�>����C��=�r��g����N>��h�C׻�{�]���K�99�������>nR?Ɓ&?J\�=�p��� U��a��n(?=�8?�O?��w?�ؗ=��վ�>3���<�o���/�>���<*��A����*��\8���<ͳ�>]A��ݠ��Wb>>���t޾��n��J���� 2M=�~��SV=D�(�վ|4����=�$
>���_� �����ժ�70J?!�j=cu��r\U��l���>��>�ܮ>x�:�g�v�R�@�����Y8�={��>��:>[������}G��9��͆>�D?n�_?/׃?%���r��TE��>�<奾qc ��g?�!�>&�?*�L>���=O���7j��;d�E�i��>gG�>Q���pH�.E��H���67$�؋�>29?b�>,u?a�S?C+?�a?F>'?�w ?��>:���ȁ��JB&?舃?O��=F�Խ#�T�� 9��F����>�)?V�B����>C�?�?��&?�Q?H�?��>�� ��@@����>\T�>��W��b��|`>�J?ߕ�>�?Y?�ԃ?�=>~5��颾�𩽢E�=A>�2?�8#?��?���>��>5s}����R+�>��O?~Έ?��l?��M><�?��`>��?!^*���>?�>	��>y�E?2xd?M�0?E�?Xx�<����ͽ�v<���ؤ<Pa>�#c�����7��j��=#��G9k��덽�hk�Q�=�0=>i_�>��y>��Ǿ ��=)
�E����J>8N�<�YH�&����$����Js�>���>���>ޞ�����=��?��>�5�t�H?L?���>k�
TI�}��$:=�Q�>�_P?���=P����W���6����>O"�?�	e?n]�Ǿ�xc?G�b?;U���e�dݴ��9B��.���M??r�.?�0����>@{?iC_?Vl�>�/��E��+���cd��t.�;�t=Z�>�����W4�+ӵ>�E.?�w�>R>��%�@	�7̇����p��>7K�?���?��?z,>C��d��2�@ܜ�AgX?�y�>�?��?no=C���w�I��,��I�ؾ�Y���/��EL�5�����,��l�=�?�b?��?Q�N?����{���q�ѯ����U��/�J$�ݲ!��<�0`&��$=��mƾs���� ��`>����"�E��1�?5?CQ=���>ᶾ#B ��fᾠ!�=+�ɾ@���~n����)�=� >�X.�[����l��n)?�?�,�>��$?�E���;�٩`��"A�J"�'��=i��>?[�>Ǌ�>�J0>B�4=�E+��˞�c~���S��9v>�xc?#�K?g�n?qp��(1�������!��/�:\���B>pf>*��>�W����8&�`W>�n�r�����u��1�	���~=Ǳ2?�%�>ɸ�>QN�?6?�{	��i���`x�t�1���<�.�>�i?�@�>R�>�нr� �r��>�Gm?���>k��>2��9h�q�w��$�����>&ϴ>���>q�z>�M&�z7[��͏�>���#:���=սh?�ك���`�D�>.�P?��)<ܩ<�j�>�˒�{"��i��iC���>�?bR�=��?>l!ƾ���5���ɗ�P�(?��?������)��w>�� ?q��>;��>���?V�>����9�a���?��\?�kI?��A?-��>�Z=�M���ǽ��%�Y�==|^�>�Y>�Ur=C��=�b�B ]��.�ʈ\=k#�=��μ9��S
<�㳼�x[<i=>t3>�mۿODK�Z�پK	���T>
��戾����d��۵��a�����2Yx�R���'��V��:c�Ƥ����l���?&<�?X~��5.������O���t������>t�q�ܥ���������)���������c!�-�O�%i�/�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�@?u�(���;_2=E��>�?�%>�_M�yv �᷾�\�>-��?�)�?k�=��W��RZ� 	_?v�<[J�y���s��=���=DS$=.a���M>��>���2��v���O5>�Sz>a�/��r�z
V����<�K]>�L������̄?@Y\� f�-�/��d���>��T?'5�>�z�=z�,?�2H�XxϿ�\�wa?`,�?��?��(?❿�߿�>C�ܾ��M?<_6?���>�j&���t��E�=���3�����:V����=�v�>J>a�,��k�?'O��}���b�=7�q�ƿl�$�!w�|o=�(غ�[��g�k���(U��$���no����sh=���=3Q>�b�>�W>�&Z>�eW?��k?�V�>�{>bE�큉�ξ��D��x��ث��+��R�N�;�߾�	������~�ɾ!#=�%��=8R�,����� ���b���F���.?�q$>��ʾ��M��?-<�oʾʿ���΄��䥽�.̾A�1�p"n�R˟?=�A?����@�V�����o�f���V�W?P�w��쬾	��=]ı���=�"�>懢=��⾱3��~S���(?Fr0?�6���3��b�7>_H=���=8$?R�?k>�'�>�R?��G��8�6�Q>��m>�v�>��a>�46=�j��w%���$?�*Z?q(��,��Y�>�-��VWc��=�=[:�>�?��;��N�A>�(U=z?7�K��<R�<�:=Z�[?���>@5��_J�庚������<��r?BK6?U�?=a?J�B?��H����ٱg�0���pJ=��[?h�?�<�=�����ھ3�����?�%e?ϼo>L���$���&�)�a��1y?��?%I)? �ؼ�������\�M��%?��v?�r^�is�����#�V��<�>�[�>0��>��9��k�>�>?�#��G������vY4�Þ?��@���?W�;<I�=��=s;?�[�>��O��>ƾ�{��c���ԙq=m#�>����Nev�����R,��8?Р�?��>������� ��=������?a�?�����mT<�c�t l�� ��<9Ѧ=���Ǟ,���>�6�.ž#)
�����Y����h�>@I@xH���>9L7�y��	�Ͽk��Z?Ѿ$�q�Hh?���>K�Ž�����(i���t��G��H�]����>�J>Z6���ϑ���{��;�������>�P��ۈ>I�S�.浾l៾��2<|�>R-�>�V�>�g��b���-��?1U���8οȻ���N�bX?�:�?V��?��?��I<�Ju�\|��C)���F?�@s?�Z?w:��\��5�%�j?�_��xU`���4�tHE��U>�"3?�B�>S�-�i�|=�>���>g>�#/�y�Ŀ�ٶ�?���Y��?��?�o���>r��?ts+?�i�8���[����*�e�+��<A?�2>���I�!�B0=�TҒ�¼
?V~0?{�f.��=9?�qG����0� �����L9>�'���=Ǿ^�z�����2r���~�A욾U�?h@��?��o��K'��4?�=�>&6@��GӾu�+�9�>��u>�� ��j����=�:�O�#���>���?>@��?Y���)�>a�=�u>?ec�>m��?+�=�n�>Z�>����0�<ʆ>��)>�uǻ(R�>��F?&~�>��=��T�:W0�5MA���[�a�
�Ut>�'I�>��`?�]Y?�p>=�㽵漴���+�H�&���뼜�b�Wh���gѽ��Z>��>˯4>b�kE���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?V��P��a~�!��a7����=��7?}0���z>���>��=!ov�������s��>�B�?m{�?#��>�l?o�o���B�d�1=�M�>-�k?gs?�yn��󾭴B>��?.������6L�%f?��
@ru@X�^?���޼������徿�/�\y�=܅y>���>�밸^j\<��=��=�?ѽ��=�r>ไ>|S,>�->IP|<|�{=�[}�G�!��ߜ�``�N�=�86�r�#�������g�$�*��۾����QF �	?�!y��*��ذ6�t���l�=�4V?�Q?�m? ' ?vd���L#> ���:d=��w��=���>Y�0?mzJ?��)?�G�=B��i�d��ɀ�Z����[���7�>.�N>p��>�>��>��5�ZJ>n�?>��>���=V8=|\ �J<=�M>k��>���>/�>�C<>��>Eϴ��1��f�h��
w�^̽/�?v���M�J��1���9��Ԧ���h�=Cb.?|>���?пe����2H?"���u)�ֹ+���>x�0?�cW? �>(��j�T�6:>C����j�3`>�+ �dl���)��%Q>ql?�Up>�5�>C�0��~9�G�(m���r�>�3?/�����o�/CC�F�޾^G7>�U�>�~�;g��������|��o�#z=E:?g�?����Iη�[�g�ɉ��TUD>�If>ɰ�=/
�=;iF>Lq������Q&��:P=1$�=y}X>���>vF�>U�6>���>�྾��ս���>-">4Ae>�K?��@?��Ὅ���Y댾�����>���>ސX>���= 6�����e�>��>՜��3?�>� ��l�k�=dN��kI����j����=U�����=w��<���ef��z�=��{?�ʥ�������羥��n�=?��?��=�50���%��¦��ì�� �?@��?���qNY��?��?�W��6��=Dz�>��>�+þ؀Q��??�Jݽܺ�� �	�k���#�?�%�?�������n��>�
'?`�߾Ph�>zx��Z�������u�y�#=R��>�8H?�V����O�e>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?roi>�g۾>`Z����>һ@?�R?�>�9���'���?�޶?֯�?1I>���?��s?Hl�>�Xx�,Z/�5�������\=�O[;a�>7Y>����fF��֓��g����j�]���a>i�$=��>�S� 4���G�=g����I��	�f�ɤ�>�*q>��I>�W�>:� ?-`�>A��>>M=�c��a‾7���pJ?�.�?�7�xhs�m�B=:|=1�$�>@e4?�P=09پ��>%�H?�l?O�F?n�>�+	�V������������ =�Rl>�?+S�>�S۽��K>ތ��y�ō>C�>��s���ݾ�1���O=)�>S!?!�>T-=M� ?�#?��j>�'�>�bE��8����E���>��>�F?M�~?4�?|ع��X3�<��桿%�[��GN>��x?[U?x��>k���9����D��yI�������?sg?A��
?�/�?��??�A?G#f>[����׾㺭���>M�!?t���$A��`&����-�?2a?Ξ�>پ��yʽb�ҼeR�	C���?�[?�&?p �+�a��tþ9�<� �5#�E~O<m�A��>�>�4���]�==8>]��=l�m��H5�EmY<��=H��>�x�=�}4�FҌ��,?Gj�`��V'�=^�s� `D��ـ>�WJ>#���j�]?Z�?�VS{�.���9��Q��F�?jg�?�g�?�-���\g���<?�	�?Sr?��>࿭�,�ݾ"@��`y�7�x�Ǔ�>���>ƈ��S�ܨ��~��o���_�ǽ#-�
\�>lI�>q?5��>eO>�o�>K���&������5k^�(N��S8��r.�1f� B��&/"�n��J���r|�x��>	Ƌ��E�>͇
?�Lg>t�{>-��>�һAތ>!R>��~>�%�>m�W>(�3>�>r<ƗͽߚJ?��˾�!��s׾�`>��f?�S/?n؈>�.�Ut��9�
��a;?��?�~�?\>��k�5s+���?���>o�{��3?<@���5=��d���p����>��D>~ޯ><�����q�T%a��Ѿ=q0?W�?�]=�����P=s���"%o=�N�?��(?L�)�j�Q���o���W��S�О�=h��f��@�$�x�p��ꏿ�]���"����(��^*=�*?��?e��]��"��&k��?�Ijf>��>L"�>F�>�wI>m�	��1�^�;O'�ô���L�>G\{?��>hI?��;?�L?�F?L�>��>h����c�>c��<̶�>���>�f7?#�(?�E,?|?_:)?j^[>m#����ԡܾ��?ͺ?[?�#
?��>>�Gi̽^��� ,1;bMz�BF�\j}=8�<y�ٽ��v���o=��W>�?�2��{�,�������>�P?{�>���>��v��3_�[Hf>���>��?��>��
�g[Z�_Ѿ���>p�?�G3��=�0>��=���<Q�=��>�����z�V�(�=�K=�V�=l��=ZY=
����*�<�A=w;>X	?�7)?�>��
>�������)��V�	>���>�v�>��>oZľ�n��n�����_��B�>���?��?,�a=P�>d� >y������^���ѕ�ɳ�����>�3?�5`?Z�?�>?��?M�=���ƭ�����v��Ւ)?p!,?3��>�����ʾ��Չ3�۝?c[?n<a�ø��;)��¾��Խ��>�[/�#/~����)D�}�������~��2��?꿝?BA�K�6��x�Ͽ���[��o�C?"�>Y�>O�>I�)�f�g�U%��1;>ߊ�>BR?���>�G�>?�m?�?#?əP��S���F���~ʾo�a����>��?��?�a�?��t>t�z�=M�������#���=Q�3�s���\���h>�uV>}5?wɣ>�B�=(�6=4�;�I�;η�>�b�=�H=�2}>���>8�>���6@G?ϒ�>ze�����k�˾D���sY;�v?&v�?u�'?+�g=���k�V����>�ţ?� �?<�F?lC�C>��7=,���\Ͼ�Ȼ>W��>�<x>d��=AcW>�I�>9��>Ǘ�>�R���#��1F�N>�<W��>ثF?a�a=mfؿ��o��jZ>>hMO>�^!��"s�bd�>�
>���.�)P��H���⸾�`��L����ס�c��g>� Fž^�>�t�=S�f>ȵ=\��=�	N=��=j����Y>�pl=�Se�ck�=w �=��CZ��o	�<`�_�m����>�=���o�z?�rA?�� ?"�7?��>|�1>G����>�3�!?:7>ϖ�����:�2�UÎ��ȋ����Aʾ�wZ�W���S
>�&��>_>j'�=n�<���=� =���=�	��=���=d�=�Ɵ=%��=W�'>��&>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>И8> _>�$R��1�&aZ��Od�%)W��n!?r:��aɾ�l�>DY�=�*߾��ƾW�0=�p8>|�a=���!\��ɖ=�n}�ߒG=-�x=Ԉ>k�A>��= ���C�=��N=���=�3N>*Xb��6���'�*�8=��=�Oe>.�&>�v�>�'?�T*?��N?f�R>�ޡ��l��������>>�5�=��>�=�f==���>�2?�[?�{d?�&�>u��=��>�U>lG�(̓��|���ľ���_0�?���?<��>�hY>}�Y��1��9�����?FO?b��>妱>�T���࿳_&�\Z.��ۘ�m`9��+=4�q��}U���w������=�5�>��>�ϟ>/�x>��9>�SN>��>��>���<ȱ�=����<]���Qt�=�����<�IƼXĕ��,�J�+�R��N]�;�ـ;u�Z<���;���=/��>\>��>P=�=���[N/>ݻ����L�п�=	M���(B�2d��E~�" /�?6�h�B>_SX>棄�F0����?Q�Y>�t?>��?�=u?��>m*���վXO��Ae��?S����=�> =� �;��V`�y�M�(sҾ���>T�>��>Y�l>�
,��!?�v�w=��^5���>�~������)��8q��?�������i���׺<�D?�E��l��="~?�I?��?��>f��7�ؾ;.0>pH����=��.q�>f��t�?�'?��>�쾾�D���˾�L���ѷ>�)I���O���k�0�,���˷�Ey�>�۪�Ӻоv63�\��p⏿�B�6q���>ìO?��?jqb�C`���O���oن�YS?�g?�f�>�e?�f?��������%��=E�n?���?)-�?�>d=�=�ǯ����>��?Xٕ?�|�?�As?M�;��T�>BU<"�+>_C����=��>^�=h�=4v?�?5�?Z8���^	����c��X���<�"�=-"�>���>�in>��=�d=,՝=��Y>+��>I��>T(g>Z-�>C��>�Ģ��P�@%?�j�=��>,�,?嗇>O�n=.�H���o=���:�J��)��fн������=Se&���<�P��|��>� Ŀ��?U�p>=�
�[Z#? 4�����ކB>�E>n�����>~R>�t>-8�>�3�>��>���>�2>�FӾ�>����d!��,C�P�R�t�Ѿ}z>Μ���	&���+w��|BI�mn��Vg��j�<.��&<=�ʽ<$H�?ѻ�� �k��)�����2�?�[�>�6?vڌ����V�>���>�Ǎ>�J��^���aȍ��gᾐ�?7��?a<O>�Õ>�ea?��?4�H��SA�moY�ԉt�_�B�m@c�Ib�����kF��]���p{�:�a?�}w?0=?�=��>���?�C!��*����>�c+��H�2��<~��>�㰾��X���ž۬�����L`>��f?<�~?U?w�<��� �Y�=>Q�"?��&?jQ?�sd?��9?4��L?�
m>�,?���>��:?�?�?�>9CU>�j�=Qi��>$k�Ԩ��*�*���ʽH�=h={�>���=Ź=�/K�b�j�죹��
����;�6����<ʴe=�b�=�>���>�D`?��?O��>Ɛ?xb1��I#�������?o==����>c��]c���>�|=>�sl?�Ш?v�b?�><6!� -�;�>�L�>��P>�J]>�r�>���9Z�^�/=	��=�F>�r=�`����T�#.�����<qq/>C�>���>��<9">D羍���U��>+nA����r9�5&D�!�/��Pn�(9�>�M?�s4?^R>����C�����O�v%?	�H?�oQ?M�w?�L�=_)��Q�C�`�K����=�>���=�{�뎜��g���>��W<��r>�]��H_���E>����߾��c�?:�M޾��!=�
���=�P	�{G�UMu�U��=�&>����w"�d7��kq��7�G?� �=���֖$�:6��fa(>斧>+h�>%k�0����b@�+��\�m=�L�>��'>:��[���ՑG�7e�`X�>hrE?�U_?\^�??����r�L�B�7���k����ļ[?�_�>�g?@�@>%��=Wб���}�d�{�F����>�p�>�F�G����r�����$�ކ�>�n?f� >E�?h�R?�
?�q`?L+*?5G?9�>z���\����@&?���?K��="Խ!�T���8�&%F����>8^)?�C��n�>�?,�?j�&?�Q?z�?��>�� ��@����>�=�>M�W�5P��Z�_>�J?~�>�aY?a˃?^�=>��5����W>��k��=f�>��2?�K#?Έ?Yk�>���>����V�=��>�c?�/�?��o?k��=�?<82>���>1��=���>܊�>�?�XO?��s?�J?��>���<a8���:���Js���O�n��;[�H<�y=	���,t��<����<�޳;_��3I�������D�������;1�>��>R����ON>�G��E���|">D��ॾ$���	�y�i�=w�z>�\?X�>\ǵ�%�=�ط>=�>cR�(:?���>�~?�0��Zb��<�������w�>�8?;�^=]Tt�ϙ��~����s?�j?�OK�s��z�e?�VS?ɜ�-8�V�ؾk|���ܾ^�I?���>D��Ac�>o��?v?���>B� l�f뙿�c���%�\�=7E�>�Z��v|a���>vI?��>�$[>�<s'վ�q�����Z?� �?�d�?~��?�I>Ģ`�3��Y���Ӕ��x�d?��?���?#?R��<e�ྱR{�} �����(p��u�¾F��Ϧ�z�h�tꞾ�a=�⨸<ē?Ѻ`?��r?�;Z?fO�^e��u\���s�a�d�������'�"{N���;��Ok��t�?ؾ�y����=Qܐ���E�%��?SW>?79��K��>-�p�����6���&�>���1�M�2n><$o�Ge�<���Pё������Y˾�m%?:�>���>�;?Z�e�%�=�d�1�W�6�20����=�Ds>�L�>נ>����Z���|����Z��Ѽ�Bv>�|c?�K?�n?�~��#1��~��O�!�H�.�'Y����B>�f>�Ɖ>��W���>&��Y>���r�d��!t��J�	��1=k�2?0*�>6��>�F�?�?cj	�?W���Vx�v1�z��<*(�>v i?�F�> �>1�Ͻ=� ����>��q?i�>^p�>	�����,T�qq�E@�>���><J?':k>jsc�Lt]�9������A�s�=Cj?�v���k�M�>{�J?���=�.�=�x�>�[������9��|e��w">�?׽�= �1>����.% �rp�gz��{b)?�<?�ג��*���|>�"?a��>���>B�?��>��¾&��:��?��^?r�I?pA?��>�=}f��q�Ƚ2V&�EA-={u�>5�Z>��o=���=;��s�\�^N ��PJ=g��=��̼�R���<�����QN<���<�H3>�)ۿ�{K�I�ؾ�4�I����g���ڳ��i��dE�Tp����&�v����9���V�d����2s�N��?��?z���OX��9Ǚ���~�������>r����29�����]��z�ྼڬ�(!�)�P��i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��6�"���8�� >gC�<	-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾r1�<��?6�-?��>Ŏr�1�ɿc���}¤<���?0�@ʕA?�V'�(�W2C=�X�>��	?��C>�,�
�S���F�>@b�?ފ?y�I=�(X�G��jc?�?<W�F������=b֥=�X=F+��O>r��>�t� AA���彔�8>��>Y����0^��<�T^>�սH��,Մ?�z\�uf�X�/��T���T>��T?�*�>;9�=g�,?v7H�T}Ͽ�\��*a?�0�?���?7�(?�ڿ�ٚ>s�ܾt�M?\D6?���>�d&��t�A��=�3�Z���L���&V����=���>��>N�,������O�[F����=�O��mĿ߹%��|'�*�=�Ϧ=����b��h拽-+k��|��g��	Ē��d�=?N2>�2>
Vt>��.=*�U=��N?%r?��?�tQ>�޽Ͻ�l��ڧ*�k�X�\������Zr���$���b�0�Ӿ��
�ı �`@��(�""=�d��=$5R�ߗ��� ���b�w�F���.?Xv$>��ʾ��M��,<nʾ��e����好l.̾��1��#n��̟?]�A?������V����X)�l����W?�R�9������=`ʱ�]�=�!�>~��=���7!3��~S�YD3??gd���l�����=���Ѹ=�.?{��>t-�=��>�4?)���o�� � >^>R�{>B��>���=���H����?#�H?���0�n��_�>P|����{�g���O>�+o�T����1>�N�<0?�� I�;P�����t��I`?���>.:�F��C����|ȼ�ib?7�"?��?�+\?�j?ڥ=D���^�S���Z>�%m@?�;�?�o�=��ƽ;��'.�OM?�0b?�g>|�v�G)��]M����io?6َ?|R!?�2!�9�������;K���>?��v?�r^�os�����h�V� =�>�[�>��>��9��k�>	�>?�#��G������tY4�(Þ?��@���?[�;<z�B��=�;?3\�>Q�O��>ƾB{������ԕq=�"�>ˌ��^ev����UR,�C�8?Ϡ�?i��>퓂������=���%c�?�&�?�k��q?f<����l�z���w�<��=�o��&���7��&ǾP�
��ٜ�^���Ά>�R@�t�& �>�%9��?��QϿ������о&�q�y�?@|�>�ʽS���V�j�wu��ZG�c�H�!i��a��>K>?W7�@��g�u���=���p��_�>��g�$�b>OHy��pƾ�߬�~<�>@:�>o{�>�;��,i¾8!�?�e�~�ɿ�)���y�<b?[��?��?�?J��<�ێ���Z���=k�R?�~?�9\?{"��Vu��L��j?�7��JG`�[�4��PE�zOU>�,3?aJ�>*�-��#}=_u>���>�>2$/��Ŀ�ֶ������?�z�?_k�/��>y�? s+?�g��2��O����*���Źh9A?!*2>Ǿ��/�!�Z/=�~�����
?Ir0?�o���2H?GP��6
�%#��D�=�Z�>c����?��ϙ���~�����Fv��f�K��?��?�Q�?B��,�&��\?c�>In��H����ʽ��?�~?i����F߾2�>H7��GL�@��>�
�?�@�!8?H5���t�����=�?�J�>���?i$ >�>�{5���9�) >}��>~�H>:[n<�c%?0??��?V�T���j�@�vfF�}�3�51۾�2�,�v>�X?�(H?o3�>x���h�c��U�t�d�5�����-~^�����9�Q�R>'�9>}�9>̱$��վ��?Lp�9�ؿ j��#p'��54?/��>�?����t�����;_?Qz�>�6� ,���%���B�_��?�G�?=�?��׾�R̼�><�>�I�>?�Խ����\�����7>1�B?Z��D��t�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?VQo���j�B>��?"������L��f?�
@u@a�^?*��ѿ���z��(٪��4>���>��->�c��$>��b=(:�=��W=�)>���>	�>4�>E�H>y_l>-��>sւ��	(�ڳ�Z3���8������b���"�'�;Y���*�w�پ����Ktʼ"O��N<�E&�=v�g;Q=n@�=S?hR?�o?O�?rY��%>�?�����<�&�I9�=���>�Y0?��J?��)?n��=�����f�J������ꬆ�(�>/�V>��>��>P��>2�T;�Q>��A>��>���=��=��һ�b�<|�H>Z��>A��>�Ǻ>\B<>�>ϴ��1���h�`	w��̽� �?{���0�J��1��:�������h�=&b.?a{>���?пy����2H?k����(�n�+���>|�0?�cW?N�>����T�{9>����j��_>�+ ��l���)��$Q>l?`�[>�@o>>�0���6�o)M�h�����>"4?�����Z=��Tt���I�ڧ۾k�K>���>�������f��g���zf��1�=�;?6?�ᗽ	���%,j�3���H�Q>߯X>��=K*�='BG>$q��̽�K�BQ&=��=��[>�w	?c��>W�=���>��羷_�����>�H�>.ɥ>[ <?��M?���A"�=��žnٝ����<Z�p>�I]>�>�dF��>���>�!g>�*q��^��&�_����>�q�=�j��I?2�4[���Hܽ�$A>!�]=����M�ս=��=��~?m���㈿T��a���lD?�*?B��=��F<��"�9 ��.H��3�?~�@(m�?j�	�ߢV�I�?�@�?G
��E��=|�>U׫>�ξ
�L�ױ?��Ž�Ƣ���	��'#�BS�?��?��/�,ʋ�#l�m6>._%?��Ӿ8}�>Ea��[�����b�u���"=��>�2H?�F���N��>��
??�Z򾌫��d�ȿixv�½�>n�?��?��m��7��L@����>��?XfY?�ei>A�۾}�Z��R�> �@?�R?%*�>x8�/�'���?{ʶ?���?�M>�?�ps?���> ���E/�rW���0��fE�=1K<���>%>�C��2H�ޒ�$툿N&j�7=���a>� = ��>I�нP���2�=q���/ר��V��M�>ӏ}>D*P>Y�>�G�>7�>*�>��'=�W����w�ؒ�3�K?���?���j2n�ؖ�<ө�=��^�R'?�B4?�`Z���Ͼ��>��\?տ�?X�Z?>Z�>s���;��z忿�~���ʖ<l�K>�+�>�G�>툽QQK>��Ծ�0D�qi�>%֗>�x��N=ھ�+��]㢻�<�>!c!?��>���=� ?��#?�Nk>a�>�vE����oE�4�>���>�p?�?��?���K�3���֡�`�[�BUN> �x?�?���>�G��QP��S�E���N��ٓ��t�?�g?V!�?L��?6??{iA?U�f>�!���׾;W��_�>��!?���ݯA��I&��\��z?�S?��>8c���mս��Լ���>����?��[?#&?���a���¾�<�p �.*J�Y�;�/D�|�>(�>�T���ʹ=�>w7�=�m��Z6���c</�=o�>E2�=<�6�����!?,?aG�?݃�5��=��r��{D���>�TL>���&�^?�_=���{�����w��U�8�?I��?�m�?���ɗh� #=?��?�?k�>dF��ׅ޾���;Fw�sx��n��>��>��l���̑��y���kG���Ž1*��9�>|y�>�_?4'?��X>�ҵ>�w���"%�g}�E��@`��:���6�b�+��i�~줾��8�tg�|��! x��-�>��9���>rx?��k>$d|>��>
����U�>�N>4�t>泡>��O>��+>�>�O�<�Ľ�JR?���^�'��辊��3B? rd?�9�>��i��l����m�?!��?X�?Jtu>�xh��++�E[?S �>+*���q
?z�:=:�뽉<����H:�7D����Nf�>&ֽ�A:���L�+�f�rS
?0?�{���o̾�g׽����-������?��??�n��1E�{ ]���U���R��ν�d���O���7�~q�䋿$ن��5���.�l�,<��-?F@�?F�ھךվ?�߾Ю����J���>���>��?>��>NR>��~G+���S���ҷ �O�?�*v?Ĉ�>W�I?4<?�wP?[kL?5��>uc�>�3��i�>Ӹ�;���>��>O�9?j�-?:70?�{?�u+?b7c>>�������ؾ�	?�?�J?�?��?�݅�sý3`����f�n�y������=<�<��׽=u�m�T=_T>��.?솎=��<��\]��?��>��?�|Խ-�!>fz>?�"!?&��=��1�rb��d"��v�>WP@?*�н�9�=�m�>���=��9>V�4>�R�<��A>ߪ<��I>���>E�=k�<���=��<�T����=���<�?3?�KG>�2�=0��=����kZ0>?a�>���>C�B>���U���ڝ����_��ѱ>�D�?���?�Ӭ�A&>��>���4���FW�`���fL�"˽>~� ?��P?���?EnO?Z0?Q�=c]�x���䒿��Ӿ:9??�!,?���>S��$�ʾ�񨿤�3�#�?�[?�;a�x��F:)�Ɏ¾��Խ�>A\/�R/~�s���D��
�����M{�����?}��?VA�m�6�{w�Q���VZ���C?�"�>]V�>��>�)���g�2%�P1;>���>�R?P
�>J�D?�[~?q�O?c �>�����ȿ�����(L��=��?X�n?M�?- �?��?�*>�>��sPp�,��F�<�$�b4��7>���=L�a>��>��>	 >̽߶�=AU��LD>0M�=u7�>�Uj>���>��>�!Q=�tK?.��>c���4]�BX��
}꾦�=�yy?�/�?��/?n'��xn�� y]��^߾+-�>
��?[��?�1Q?6c���"$>_�Ө�!�;���=]B�>2�}>	�=>��>~��>/2�>�:�>ҍ(�v�%�@4G��L�5q ?T�S?ߙx;�7���a�1*ɽ7<��QZ>��*�r�YV�1*�`��\���Խ��a��j�I���F��&�������Be	�ʮ�>�!�=��>ׄ�>9>N�껈�>��8={�=��<�qʽ�>�������/�@���?!��!=Ã�k���lq?a�M?�{+?O9?�\R> |K>e}3=jf�>�)x��X?�w�=]�$�X�־҂9���Ⱦv֭�K(ݾȠ�
IB��Ӝ�h+>�Ǔ<3>-b�=���=h�a<��e>��>���=[�;�j��IR�=,��=��=�`�=��=>$>�0w??���䩝��%Q��S�Ǩ:?��>���=s�ƾu	@?��>>`5��k����^��+?���?�T�?d�?��i��j�>���厽jď=�@����2>kv�=�2����>��J>���(B��l���9�?�@w�??�ዿY�Ͽ�o/>�C>aS>��Q���1�I�f�9�\��]Q�(3!?2�:�6Yþ��>�<�=?�־�wþ��<�*>f�4=w9���Z���=�q�.i=�sO=���>�R>���=0n���f�=�K=��==�E>�
�_3��)��L3=�=P�h>LL>�y�>_	?�K?��S?&��>m������3���_=�p*�d{ >�	I=�,>�>&�[?�Q?kT:?��>~H>~��>Z�>�FA��U�c2�Y�����>$>�?$��?�h�>����K8M���6��yW�\��!?�D?-׾>�i�=����t߿~ky�m�Z�,�>��k>���=Uf۽�i�V��!�������$>��>�>�ٌ>vN�>�N���9>�>4�#>���<��<�9+=y�սp[ʽ��=��*�������u��Ix;��<¤=6�Z=?���7�<ؓ��;0� ��=_��>V:>��>"z�=��� J/>����Z�L��ƿ=1B���'B�1d��G~��/��X6�\�B>�:X>�����3����?��Y>Ok?>{��?�Au?��>�"���վ�Q��y8e�`S�3˸=u�>��<�@{;�8X`���M��|Ҿ��>��>�z�>.!l>�(,�i?��4x=����J5�s:�>O������@q��A���響;i�P
�3�D?�0��w#�=w~?zI?�؏?��>Ɨ��Xؾ��.>{���*=��j�p� ���4�?��&?*S�>���D�	�˾D�ƽ���>�J)� �N��V���^/���J����cM�>gA��̃Ͼ�c8�|��/+����B��m����>cL?�8�?M�C����mL��������y�>�6h?�z�>�7 ?j�?����"��"Y{�ּ�=t?tH�?�>�?�>���=N괽�5�>�+	?���?3��?>�s?��?�i�>�;�� >7☽��=׽>ԉ�=�\�=@w?�
? �
?�S��i�	���� ��^��/�<[ڡ=É�>x�>u�r>e�=��g=�Z�=4/\>�מ>��>x�d>�>�M�>^�������*?I}:>���>]�2?;A�>o)=��؉<3hz�F�q��<�~t��8ݽ}~���~%�CV�/���Um�>�ſNo�?��{>��	�u�?*��ϥ����5>U;;>�%�h/�>�� >��e>K��>�I�>��>���>+�B>�FӾ�~>����d!�s,C���R��Ѿ&}z>d����	&�Ο�#y��^BI��n��bg��j�N.��~<=����<H�?׻����k���)����'�?�[�>�6?�ڌ�>��k�>���>fǍ>�J��V���Gȍ��gᾉ�?��?*�J>$�>[�d?UfS?,Z9�����Q��?8��D�L|����k��2��ꑕ�[r
�f�N��Z?�A�?NT=?��z�v �>���?A���}�Q��>�3���L���=(g%>��/Oþ���O�k�2u=�}�>2��?��?A}?g�{���m�� '>��:?��1? Ot?:�1?R�;?C��d�$?1p3>�F?�p?�M5?O�.?`�
?j2>��=�>��S�'==6����ѽByʽR��f�3=w[{=l'θ'?<�=P�<���&�ټA�;	���'�<c:=��=��=�>:^?Ld�>U��>�=?����3������d�>E���i��jŰ�7ؾϕҾ��=0t�?���?3�b?�5>���q�l+�=]>�Y>�>��>Ȳ�k@�RC�=yk�>�Z>д[<a0�/�������q�k�M="�=m�>�+�>����<>�j��fW���[>�oO��¾�c���M��!4�x��/��>EO?\&?G��=��ھ`n^��_��b%?��;?��G?�{?�(=ǡþ��0���F���Zt�>�*�_��p������F.�Q�A=�W�>����쫾5�V>R���^پ��i���A���ܾww=6�֦<�u	��(޾�~��C<�=��=�ھ��T!������⫿5J?#R�=�m���tM��n���v>Y��>/�>ک����q�؟;�7���o=��>q~'>:Լ&���I��I��?�>�PE?xU_?k�?�"��;s���B�Ȭ���f���ȼ�?~q�>�g?�B>���=|�����F�d�fG��>���>[��w�G� >��=*��(�$�ъ�>7:?'�>��?��R?��
?$�`?�*?uC?�(�>������dD&?���?Ä=��Խ��T�i	9��F�q�>x)?�B���>6?��?��&?�Q?��?->Z� �UA@����>qP�>��W��d���_>x�J?A��>1AY?�܃?��=>�o5��Ƣ�q��]<�=1>��2?c;#?ɭ?��>'e�>IӒ��E=���>A�W?�?��o?J�	>��?`tm>�U?�3=�k�>l>�>��?ٽE?�Mh?78?S�>YmM<�l�����i�W�U��<�=@h�<ڱo=����7P�)����<�>ƺW�|�O+�ർ�?��:���73;}x�>Ο�>*����8>@.��f�����=W��<ᾥ�����ϾM��<�Ӣ>L?�>L5/��3{=}�>�c�>7�˶1?1�>�K?o�]5���^*=Jā=<R�>�T?1��=�!��)o���
���rg���?��g?��ѽ����q�b?;�]?��`=�2�þ}�b��&�g�O?�
?��F����>�0?d�q?���>8g��Mn��%��*b�e�h���=S��>���TJd��>�?7?���>��a>��=�|۾ƿw�������?�׌?C��?Lˊ?�*>H6o��b���xß�ž�?B
?��־�&?�n�=����F����`�/�	�գ���꾢>���澨�n�_����7;�p�=��&?|=?yw?~�c?�񾖘t�U�]�X,u��n�g�fe �8��y&3��	-���^�������ξ���mR5>%�/"N�E�?HD/?/SS��U�> M������;Ѓ>>;汾j�
��
�<X���x�2�@�<�f��]�@�����7#?+�>9\�>��??8�S�)^F��4�rD3�������=_}�>�'�>�N�>0-��$�%��Sѽ���Q�`v��8v>�yc?�K?,�n?2p�i'1� ����!�^/�MU����B>;q>ۻ�>@�W����9&�U>���r�Y���{����	�&�~=C�2?�$�>^��>PM�?1?�u	��i���Nx�2�1���<�.�>�i?�7�>��>��Ͻ�� �Y��>��o?[Å>fs�=wK~��~�
�d�$����>��>W>�>i�>�;|�/Y��	��r���ǗP�rz>��?(N��{����>H#V?���<���<��>+���m*�'q�]��_$�=�M?�&�=��=�kƾ��	�������))?H;?˥��~D*���}>K "?���>�:�>"0�?�R�>��¾����/�?�t^?��I?�GA?"A�>��=j>����Ƚ=*'�=M,=?��>��[>(-p=p��=���>	]��e �6�A=���=Q�ͼ�d����<8�����I<���<d;4>��ڿ�%J���Ҿ �	�i������z����tY��);�����צ��s��H����A�w(Q�W6k���������=�?���?��R��!��β����w�ql޾ms�>��?�١�����Z�$��������M����)�O�/�m��h�P�'?�����ǿ򰡿�:ܾ4! ?�A ?5�y?��8�"���8�#� >�C�<�,����뾭����ο>�����^?���>��/��r��>ޥ�>�X>�Hq>����螾`1�<��?7�-?��>Ǝr�0�ɿb���¤<���?/�@ǡA?�=(����ˀ6=�d�>�?�r1>�9�����[����>���?���?֨�="�U�L7��Gb?�W\<||G�n���l#�=�W�=Q+4=,-��*@>�]�>2��.,@�9��"S5>���>aP,�m;��^���<� ]>�"ҽ�B��Մ?Nz\�Bf��/��T���O>��T?2+�>.5�=H�,?�7H�j}Ͽc�\�{*a?�0�?��?*�(?Zٿ��ؚ>R�ܾ?�M?qD6?y��>�d&���t�v��=�.�u���	��&V����=��>��>��,� ����O��A�����=4 ��i¿}�"�N��e�=��=t�?����������������7н��=�x�=q�I>vr>�#>]��=�uY?�
z?#3?�5>�<��dc��Λ�+�=�E�\nq�]����\�K˾{D��p��\��w��N=%����V(=�S�=�,R�;����� �U�b�*�F���.?jg$>��ʾ��M��|*<�{ʾ�ª��Q���祽�3̾7�1��)n�#˟?+�A?z酿o�V�6���W�J��i�W?�����ެ��e�=e���AB=��>Id�=��⾆'3���S�#S/?� ?:#����L� >y��9T6=N�)?�^ ?���<���>p"?��)�+@��
�C>��->���>���>D� >C���uν�I?�5V?����4-��+�>Ʀ��dVm���Q=�">�5�:I���
Q>�F�<rC��>�R�Q@���=�\_?���>Ѿ9�z�Z�?E�����s�@�V�?ڐ'?��?�a?^7]?8�����
��R�&����>Z�?I�?��=(�ܼ����I���54?>�c?'�">�V�	��.'���
�G�%?�?C�?;������K��27�x�m?��v?�r^�Xs��n��J�V��;�>\�>���>��9��k�>~�>?�#�oG��Ⱥ��$Y4�CÞ?m�@s��?��;<� ����=�;?�\�>�O��?ƾ�x��/�����q=�"�>Z����ev����S,��8?ݠ�?���>�������#1�=s����?\p�?^�G҄<�Y���l�B2��'<d�=~Y���m�he�:���ɾ2���?��%���@j�>B�@Ҫ��"��>�L2�q��ο|X���8پ0<���T?y3�>g�ҽ$Y��i0c���o�I?��#@�3Ԅ�^B�>2�>tٖ�K ��n+|��"?�4�м�?�>>YF��>TV��A�������8<�>!�>㏑>&^��hμ�n��?���k̿uU��h	��,\?�s�?�y�?��%?J�n<��W���^���K.E?ܔr?)U?��ټ��]�8�U���j?�%���\`��4��5E�t�T>�3?pB�>1w-�dF}=-�>m��>$�>�$/��Ŀ�ֶ������?=��?z�H��>�?�~+?�Z��-�������*���~�A?*�1>������!��=�R֒�ŭ
?n0?aQ��d�)�L?� �G�V �wI����>�}���T��烾�}���i�*K���y�B��?p	@L�?JQE�|���,?���>�������/^�+?O|�>;������v��=t:W�bQ�j��>^4�?�(@�f?�a��
���f�O>�tR?s1�>��|?��B��\,>��
=Y�n��=�I>��)>�>Q��>��??�U�>�N��]�Ҿ!�)��7:�,�_��
���=�B�Y>��]?��V?�>�Nڽ9�K=<��������:���m>�C����������7>�/d>�u�>	獾�	ؾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ua~����7�c��=��7?�0��z>���>��=�nv�޻��W�s����>�B�?�{�?��>"�l?��o�P�B�}�1=7M�>Μk?�s?Qo���i�B>��?!������L��f?�
@u@a�^?*V޿l���,����k�����=�G>��A>����OP�=^�>3L=Bjh�E>VZz>\�[>Pv>�<s>t�I>��>m��Ix�'Ѡ���K�*5%�����h����룾��R�¾9���{�����_��l&��q8��}�I��=U�U?��Q?��o?Gc ?�Jw�& >�k��"�=��"��Ԇ={�>Z2?ZL?�n*?���=~�����d��H���A��=ۇ�a�>@BI>#0�>;Q�>��>m����I>�C?>�t�>�� >}q&=f���=�3O>�N�>���>��>eC<>��>Aϴ��1��e�h��
w�L̽/�?���X�J��1���9��ۦ���h�=Ab.?|>���?пg����2H?���j)��+���>x�0?�cW?5�>��y�T�6:>E����j�$`>�+ ��l���)�v%Q>ml?��f>��w>�2��]8��P����e{}>��5?������5��/t���G��cݾ܌H>�>�vh���ܖ�S{���j���=t�:?�?�������t���sS>��\>��7=Ӈ�=}�J>ѧk�/�½�4D�]y==P��=w�^>�?s�S>��}=?�>�֖�x�1�>S>�>O�;?1}?Vý�G��
��e 2��A�>'y�>x>�(>��J�!��=R=�>Am�>����Ƽ�����'�|WP>������6�B�K�x=W���G\�=�,J=tS���2�MB`=M�u?����7b�p��;��>�'/?� =# ��#����T-�����/�Q�f��?	E@���?E�5���m�J�$?��Q?�μ�	����=��g> ��/ھ�d�>Xa�=C����f�G�U��?��?�6�<Z��n�r�>A�,?�	�Vh�>^x��Z�������u�Y�#=J��>�8H?�V��j�O�a>�w
?�?�^�ߩ����ȿ8|v����>[�?���?h�m��A���@����>8��?�gY?Toi>�g۾Q`Z����>λ@?�R?�>�9���'�{�?�޶?Я�?qI>���?��s?�k�>=1x��Z/��6��ږ���q=�[;1e�>X>!���rgF��ד��h��W�j������a>X�$=�>�D�4��U9�=�����H����f�#��>�,q>P�I>�V�>p� ?�a�>���>�x=�n��ှ����H�K?��?����2n����<�T�=ڠ^�*%?AD4?m�Y�|�Ͼk֨>��\?�?�Z?V�>F�� =���濿������<��K>�7�>�>�>GF��[<K>)�Ծ�0D�_o�>F�>�夼Aھ�-������1H�>h!?���>�ɮ=ڙ ?��#?��j>�(�>AaE��9��S�E����>٢�>�H?�~?��?�Թ��Z3�����桿��[�f;N>��x?V?pʕ>`���택��kE��AI�,���]��?�tg?}S�2?;2�?�??^�A?y)f>߇�%ؾe�����>��!?C���A��F&����|?�Q? ��>���"�ս�[ռ����u����?!\??&?}���(a�u�¾��<�M#��U�0�;�bD���>-�>F���Ύ�=�>�ذ=�Rm��I6�k�f<�j�=�>��=J"7�Re��p=,?�kG��ۃ�X�=��r��yD���>�OL>�����^?�l=���{���=x���U�3�?ߠ�?�k�?S��&�h�J$=?	�?c?"�>�I���}޾@���Pw�zx�qu�1�>��>��l�<�菤�y����E��e�Ž�M"�{o�>�_�>�`?&,�>�mQ>�+�>����%�6����^�[�[8��
/�!��a����+���(�֏���w��g�>zƂ��N�>O�
?e�i>��{>HQ�>���E�>�@Q> �>��>�U>1>��>k@<U�̽_�Q?���&m$���來�=0�
?q��>v�S>����֋��*�}@Z?�:�?���?�Y�>i`��,�;��?)�>-߄���>@SF��8H>������.q�=^>�;�<�u�>~?���I;��fO��۾��?r�?=u7=蟤���><�i����a=D��?�j)?	*�muQ��1o�_�W��S�����i�����"%�pp�� ��-P��%��k�(�_�,=:�*?l6�?
��_r�d���|k�yY?�B�f>NZ�>W+�>�>I>�	��1�@]���&�Eb��Y.�>�D{?�̌>�G?,:?�O?%-I?G3�>�t�>�̫��>�>���;H�>/�>��6?S)?��-?�?�P*?�[>B�꽒���iپ4_?��?T?�?� ?�ˇ�,�ݽ�c�����E�r�?�h��I�=[�<�`߽��~��(=PD`>�?���n8��P���/k>*�7?��>k��>EU��:�~�\� =�V�>��
?CՎ>i����r�T��Ȇ�> ��?�K���=d?*>=!�=m�{�>����d�=jǼ�2U�=DJp��A:��w<J�=�*�=����x'$8ٻ�:*��;��<j!?HI ?aU�>}>L�����^0�G��=P1h>�a>� >ΙӾ&势�����:g��`~>q�?Nյ?�d=:I�=zq�=MU���e¾��lȸ�	ܷ<3�?;� ?x�S?;ܑ?!4??�8&?+W >�(�:ʓ��چ��Ƣ��i?q!,?���>�����ʾu�P�3�̝?Z[?G<a�����;)�ڐ¾��Խ��>�[/��.~�d���D�������m~�����?ҿ�?=A���6��w�v����[��M�C?�"�>GW�>��>A�)��g��$�83;>9��>�R?=.�>R�O?5,{?�[?�T> �8�5��ՙ��m7�߭!>�@?x��?���?K*y?�s�>`y>�)��߾�`�����J#��낾�W=��Y>�m�>�,�>��>n��=�Ƚ�9����>�Q.�=Yeb>���>	��>���>t�w>��<�VU?��>u{ž��T��i
�������?ût?�j?:X�<8�	�oI`�`�����>鬪?y��?E�_?9���H�>��r=�������e��>�Z?HT>r�>hF?kw�>^?�5?h4��d��C�2�Ϯ�{?aQ?�8�=k¿��U�]��6�u�	e�<K�se��հ�<�&�6Ԑ�ݺ~�����8ʾ�I���f��7앾I�˾k)���쾯/?� >괇>��=��<L}���=���=�< >��>�3���(�q>�rx�bLս�"3�ca�<�U���޼�	k�̧b?��?��?$�>q�>?�>H��=��?:>�qE?:��=+��=���Cr���x����f���j1����P�Ū�X��=��<q��=؀�>*�s=��,�1�=7�=��$<�Qp���9=�2�=�<>���=���=��[>* >��v?�M��L$����P�D��Ä:?O�>�%�=I'Ǿ��>?��=>�'������)����?���?�K�?�n?��h�`��>�꡾�瓽q}�=���� D4>��=	5�K�>�qL>3{�����B��o�?��@|�??�����Ͽ80>|'9><f>�ER��41��]��
g�+�X��j!?�:�{�ʾ*o�>�>�=an޾��ƾ��$=c�6>,b=����4\�E��=-Sx�(�A=�Ou=��>�C>��=E�2��=U�J=6W�=�M>���#�<���'�\c7=ja�=��`>ª&>�j�>�3?�Y!?�g?$י>�q����žBy���{G>�`�=Y�>�P�N�D>4��>�4?}M?q�R?���>f�S=p��>�{�>},�O$l��q��fMe�)s�@~�?C�?�ө>�� >ħ����/�J�4������u�>d:7?�E�>L�>1��Q⿄�E���b����Z�=v|�=��f��À�S۽4�Z�!�3��\ >$Ċ>Y�>�o�>�>s>�S�=�ga>Ks�>�~B>�9�=��6=�O��`]�=Wp�YL�<���^��A�ʽNm�;�k������ƼO�;�V鼯���%�����=���>':>"��>4��=i���I/>*�����L��ҿ=0>��;)B��1d��H~��/�|T6�n�B>&X>x���3���?��Y>~?>u��?QBu?��>U���վ6P��$-e��NS�*ٸ=�>m�<�xy;��V`���M��qҾ���>w�>ڢ�>\�k>|�+��?�Dx=l�ᾎ55���>�t�������0q��>��i��)i�˱���D?�>����=�%~?,�I?̏?�G�>ꮗ�*�ؾ$�/>�M��g=���Qq�쒽��?��&?v��>���PE�09̾�4�>lyH���O�����+�0���!�T뷾�Y�>T���о�63��b�������B�V7r�'�>i�O?��?uUa��Z���BO�X���͆��A?�tg?��>i?�N?0s���z�0Y����=��n?���?�:�?j>˸�=����%d�>��	?af�?6ő?�vs?�=����>�;&>����N�=H+
>#�=&��=��?h	?V�?쑜�Bu	�Uh񾄎𾑁_�ɾ�<�)�=���>@�>�!w>��=��h=�u�=��\>��>��>.6d>�ѣ>M؈>��Ѿm~��O;?�W9>n�M>U�@?oU�>8M=�~�)+%=�?���=���������f"�f'��h����ܽvK���?<�ο;:�?��>���8�>�_־�%�����=
��>�a�����>� �=/2�>��> ��>H��=�T�>�E�>�FӾ[>����d!��,C�O�R�}�Ѿ�}z>�����	&����w��nBI��n��xg��j�M.��_<=��ɽ<,H�?�����k��)����Q�?�[�>�6?uڌ�i���>���>�Ǎ>�J��f���Xȍ�hᾠ�?@��?��J>�n9>�U�?�tC?���-�jtH���o�k8Q�p���؉Y��Rw�����<%��G���4�P?+~?%�0?��=���>s�?&:L��w���z>]��f;o����<�Y9>�3�u�����ȏ����=�~+?���?_�?���> �&��K�:�V>{�>D9?6gC?H�M?��H?B�t�5�E?Q��> �F?X>�>��$?�1�>��>]/0>�7	>�4ܽ	$�>?�T�;�{�霽�-��f�7</�=�M�=ԓA=r�=�w>�Y�=[vb�Ijo� �j<"o��=a�p=��=��Y=o��>�\?�'�>���>N/?�~�l,��Ý�B�?v�[=�n���I���e�����u
>��v?�è?�_?$�\>�3��_H�'w$>�͗>�`>�B>���>x�ֽ4�I���=��F>I>ҳ�=kq���Ȃ�����Q}��)�<[�>���>��|>�q��W�'>*q��*�{���d>>jQ������S��G�N2�]v�_:�>��K?�(?�w�=м辏䕽Z(f��)?�^<?xSM?�?�Ǒ=�{۾��9���J�����K�>�
�<'��M������3�:�@(�:��s>W��1��a^c>�F
�&�ݾ��n���I�]b辞�"=p��#�9=��	�׾���V�=�
>:������^���k��JI?�(m=�~��q�[�꺾�F>Yr�>bR�>��5�`�q��c>�� ���J�=�&�>�D>�{}�Bt��2G�2���\�>)E?�f_?#k�?Y�D�r���B�Ķ�����I�ɼ��?���>�q?q�A>��=�α�^���d��$G���>ן�>
����G��#��l ��;�$����>�#?��>��?��R?��
?@�`?�"*?G?I%�>{(������@&?#��?y�=��Խ�T�� 9�iF���>b�)?&�B�B��>̈?ռ?�&?�Q?�?��>ڭ ��B@�|��>WZ�>��W��a��[�_>��J?ҙ�>�<Y?aՃ?�=>�5��ꢾ]ҩ��K�=�>��2?`6#?°?���>Y��>1����N�=C��>�c?�1�?f�o?�m�=��?F2>���>�ޖ=}��>���>�
?�NO?Q�s?��J?��>�B�<:[���綽�Jr���N��v�;$J<	+y=���}t�����<@��;�<���р��f�!qE��%��!��;�Z�>�t>����0>��ľOT��O�@>b��yF��a���3~:��6�=l��>�	?6��>�3#����=Ǌ�>n6�>]���9(?��?H?V;�b��ھI�K�M�>*�A?���=��l�w|����u��Yh=�m?��^?�uW�~��EB]?3�5?���nh�U|�
0p����Tc?9*�>ɡ<�h>���?�Z�?=�?� پ�Qx�������`���:�7 _=0F>>�k,��B6����>��F?!��>�>��9>X����i�_q��[, ?��?tĬ?Cy�?�@>,@���y��N,��Y����<?"0�>�?��V	�>L�:>����+Έ�Hؗ����Ⱦ�p�L���K^þH�Pqi�~�0�e�P>?X�>��q?��:?�-H?jm��=T�ý�������:i��}4��/��{B��C�R�?��	Y���Ͼ*��2��>��ܘM��BJ�S�?��-?T�ɽsV
?�?F�"�f����E>��5��� ���#>=��V�=*��;)����>��^����?��>���>��E?�G�Z�"���#�d�1�H����=��>���>?�>�nz���E��U@�|�Ҿ/{�b���9v>�wc?�K?��n?�m� )1�&���@�!�~�/�ec����B>{l>���>F�W�]���:&��Y>�[�r�0��v��[�	�	�~=/�2?�(�>���>�O�?�?�{	��i���kx���1�s��<�1�>� i?�A�>A�>н#� ����>��l?W��>�
�>�����[!�0�{��ʽ�%�>�>O��>�o>
�,�V"\��k��*���l9���=��h?����`���>�R?���:��G<~�>K�v��!����~�'�.�>V?���=d�;>C�ž'�è{��5���B)?�4?�Ԓ�y�*�lg~>� "?�u�>/2�>�)�?7M�>.þ�s��?��^?x7J?�?A?�>k�=Z��Ƚ��&��U.=�ʇ>@�Z>�m=i��=b���\�r��ˉE=Z�=μ`���g[<�!��H<Ӫ�<��3>4hۿlaK�7پ��:��k�
�C҇��%���ۈ�3:��������\�{��y��]5���S�h�`���#�h�W��?�N�?�J���?���d��D�~����.�>hAw��6��Mʭ���Fܑ��߾3�b��  M���g�'�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�yA?8�(����2�Y=��>��	?-�?>��1����尾���>Y�?��?�HL=Y�W�e��b�d?�'�;��F�P�ӻ��=�1�=� =����J>��>�Y��@�@kܽ��4>'��>ef"�`"��]�W+�<!�]>bֽ���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=����ſ&$�L���g�<��W��f�g���ty��=����s�Z�����N=���=7�R>�*�>��X>�]>4�V?��m?lk�>�D>�Yҽy����]վ�)Ǽ�憾�(�;����> �qۜ� ��Lzݾ����@�i���˾�B=�h��=+R�Gh��:� ��b��}F�Ft.?0�">�j˾��M���<�ʾ����i�������t˾�Z1�I�m�װ�?XB?�t�V�����]�lϻ��5W?v�������v�=7y���=�'�>Ri�=���z�2��iS�x�.?Ǌ ?XL���I��NZ*>�,��Z�<�T,?$� ?U6
=D�>Oh&??�����o�d>��:>�1�>���>��>�7��J��¾$?�MX?�� ����"�>'��2�t���<0�*>��I���ȼ'dJ>Y�<l��?8�Z�z��	 =bzT?���>G����;�5椾7�b�<x6�H&�?C��>{~�>W�P?,�R?H�<��ľ`�|��a�7�Q?�̎?�=>����-��;���aR?X?SF�>g�s������������=?��?�K?^�t����$��5�X�?��v? s^�xs�����N�V�\=�>�[�>���>��9��k�>�>?�#��G�� ���vY4�$Þ?��@���?��;<��4��=�;?a\�>�O��>ƾ�z������V�q=�"�>����sev����R,�b�8?ڠ�?���>
������u��=0敾�Z�?��?x��h�i<����l��a��
q�<� �=�	��!�%����7�j�ƾ��
�7����ڿ����>�V@e[�i*�>1A8�f/�=QϿ���wHо�`q���?߆�>$�ȽK���k�j��Qu�ʬG���H�褌�Iߟ>�b>�3��M���`�{��E;��E���.�>��1��ͅ> �W�κ��Ю��Pa<�>���>�׈>���0̼��%�?��� Ϳ"��� ����V?���?N�?Y�?Γ\<�r�lw��2-��G?	t?
�Y?"u'���^��j&�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.��_?�a���p���-�)'ǽ�ʡ>r�0���\�����y��Xe�*��^y���?Z^�?��?x��! #��5%?S�>㓕�tDǾ4B�<`t�>q�>TN>��^���u>��
�:�k	>���?�w�?�l? �������eG>��}?��>_��?�G�=���>/�=>����Ҽ�(?>[�>��<_�?�&N?L2�>_v>�D��9 �[�?�� U�b���@���>f�r?�'W?x7>�ʽ�G;���V����'r��N�=�pw�4�=��r4>v�=>H�>�x%�A�����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��2a~����7���=��7?�0��z>���>�=�nv�ػ��P�s�¹�>�B�?�{�?��>�l?i�o�J�B�R�1=KM�>Ԝk?�s?�no����B>y�?�������K��f?�
@zu@Q�^?$���&��������q��&>�c>�>yD<p�B>��=�s=�+&<i�A=
�>��^>�
Q>7�6>�(>�X�>_~�s$�/���)�n�0���6T�n���_�-C�����R/����b%�ZPS��3o������Q��\�����<;�>=-?ZCz?z�?q<#??�~>pʏ>�Ҿ}�=y���>���>�~;?O.?�,?�r
���߾N�b��H���vN�qJ۽��>�,e>
P?�P�>S�>E��=i�=��>��#>��n�F1<��/=�Jf>gɺ>
l�>2Ӽ>D<>l�><ϴ��1��՛h��
w��̽+�?�����J��1���8�������l�=�a.?R{>���?пb���h2H?����})�Ÿ+���>7�0?�cW?��>����T�1;>��9�j��`>�) �$}l�(�)�%Q>&l?,e>��u>>C3��H8���P�9���L�z>Mr5?P=��Ӛ9��u�5�H�o�ݾ��N>��>@�����iؖ�B~~���h�(�}=�2:?$?dm��I����Cu�Gi���jR>.[>�=
�=�M>}s`��1½cG��./=�,�=b�_>6�?l�>�X�=��>�I���w?�A�>��<>��/>��>?
'?g�|y��	|����,�hm>��>��z>D�>z}C�[�=��>s�j>�7��i�k��L���B���T>$����_��u]�Ux=����=,��=���ݔ=�&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>@��F��s'��a�u� =i�>�XH?�V��,�K�>�ع
?%?Z�񾘺����ȿxv����>~�?^ڔ?��m�?��
@�G�>���?G�Y?�i>�<۾F�Z��ŋ>y�@?�KR?�p�>E���'��?���?�f�?�I>��?T�s?�l�>�)x�(Y/�/6��Ζ���y=Y6[;Sf�>�X>����)gF��ד��h����j����Z�a>
�$=W�>�B��3���8�=�����H����f����>p,q>=�I>�W�>f� ?Eb�>$��>�z=m���ှx���T�??��~?�(��~��p�:>|�w;�b�6C?�!??R`>b�Ǿ5m�>_�[?}��?�aH?#�>�����Y��^h���	>"��>�3?d��>�սP�3>�H;k'��3o>�Y?@�/��׾�U��p�5>ȟ�>u�+?���>��?>Ǐ ?��#?h>(�>C�E��V��d�G�<U�>D��>I�?��}?�=?pغ�b�2��������߶Z���S>$�z?Ô?B��>����������3X�����?��c?��߽�U?3��?¦A?��C?��_>{���-ݾ˔��Μ�>n�!?���*�A�Ŧ&��x���?��?`��>zÓ��bѽq����Y����?��[?2&?c|�	Sa�8�þa��<ǝ��҄��8<NcK���>oc>�d���v�=�>%��=dn���6��8w< ��=�Γ>��=��6��y��$=,?��G��ۃ�<�=��r�?xD�#�>1JL>�����^?Fl=���{�����x��]	U�� �?���?^k�?����h��$=?�?+	?S"�>K��~޾	���Pw��}x�ww���>���>��l���L���♪��F��V�Ž�i ����>���>և?�r�>אR><��>�����%�^���G���]�����8�.-�e���^������t��{��2nu�Ty�>𭓽G�>��	?q�^>#=w>���>�֥��;�>_!W>��w>���>N]\>S�4>��>�<xֽGR?������'�#�辛O���B?kQd?�X�>P4h�)j�������?�?�w�?��u>�{h��2+�7?/��>���?e
?�t8=�M	�	�<�E������k��Uu�LÎ>��ֽd':�M�?�e���
?�R?�L����̾�Jؽe����n=yN�?��(?��)���Q���o���W��S����6%h��h��\�$��p��돿�^��t%��K�(�#t*=؈*?��?ǋ���,���!k�E?��_f>R�>��>�ݾ>7|I>��	�T�1�� ^��N'�浃��L�>W{?wt�> �H?F*<?q`P?�gL?ޟ�>�ѩ>5گ�:}�>!��;�%�>�Z�>�9?I�-?�0?�?|�*?(b>�k��9��z�ؾ5?I?�I?�L?*�?@�����ƽ����{��y�[���=u,�<[ؽ��|��JS=$�R>�[?���rw8�N{��~Ak>
�7?/v�>���>�ӏ��'��,��<��>�
?%$�>6�����r��u�k�>���?�k�6=��)>��=����tݾ����=������=�j��Ų:�i�#<�S�=�J�=e�jn¹�;��;���<Nɦ>N�?���Wy�=E��i��-���U�>|��>�4�>�>����5���X�K��I>��?��?X�>8τ>0_=)6��B~(�����þ04Z��>P?��?��~?Q��?��S?�!�>`R>��4��Î�|��_ ���kM?W!,?���>����ʾ����3���?[?4<a�d��=;)��¾��Խ �>c[/��.~����VD��������0}��O��? ��?A�)�6�\x边����[��ȓC?"#�>X�>b�>_�)�(�g�/%��1;>���>xR?���>�M?�|?�\?V�V>�5�����V����ƻ?<>��@?�f�?+�?S�w?�|�>>�/���������D����I�����\= nZ>	k�>���>��>���= ������?>����=C�d>���>ƻ�>P��>$Ev>-q�<EF?B��>o�����jK������J���s?��?6i)?c�<�3�"�E������P�>Y>�?�"�?^H*?e�T�8�=�aҼ]����Oo�Ǹ>��>,t�>��=�g=s� >>��>�l�>�U�e����8���\�`�?{HG?rc�=�ÿ�q��b����E	�<ꇋ��]]�T����@X��(�=`8������x����^��٠�����Q'��-����z����>��=FC�=-<�=��<�����h�<[�>=���<��<j�o���<VB��_�|��Ve(��m<:>==!�'@��o�r?a�L?��.?3 C?/��>J�>q�a��{�>�i��/Q?�"[>�|�*=���9��a���=���%޾�ܾ��V�!���,>>QH��8>r�3>��=��<_��=Xwm=�ߕ=�9<�8=���=�#�=`�=��=�h>ey�=�6w?V���
����4Q��Z罢�:?�8�>F{�=��ƾm@?s�>>�2������vb��-?���?�T�?<�?>ti��d�>K��~㎽�q�=V����=2>s��=o�2�Q��>��J>���K��J����4�?��@��??�ዿϢϿ=a/>��>�>��Q�B*-���c���n�#�]��J?�V9�S�ξ�u>�=�_徶̾bl=��L>���=��V Y��ۡ=m,��'�=
p.=u~�>5�:>�{�=K�=���=zq�=�>��k>C^�1y?�E���5*=fc�=!Br>q	*>Q��>��?[&0?-�c?lM�>c�n��>Ͼ������>)n�=H��>;Ƀ=;A>ڿ�>�C8?< E?]�K?>4�>�(�=��>�
�>|�,�?�m�k8�vѧ��W�<���?�Ά?�m�>cZR<B4A�gX��>>�vKĽ�)?�C1?�Y?xΞ>�U����8Y&���.�3���O�4�n+=�mr�RU�����Ym�O�㽤�=�p�>���>��>DTy>�9>��N>��>��>�6�<]p�=������<� ��n��=Z�����<�vżb���,u&�	�+�������;簆; �]<à�;���=���>�:>#��>���=���B/>�����L����=�I���,B�>4d�CI~�r/��S6��B>�;X>�z��_3����?|�Y>Wi?>Y��?�Au?'�>I(�S�վ�Q���Ee�"XS�YӸ=�>��<�
y;�PX`���M��}Ҿd��>Jߎ>�>n�l>�,�G#?�[�w=��Xb5�~�>�|��a��)��9q�%@�� ���qi��dҺ�D?�F��i��=f"~?��I?_�?���>��نؾ6;0>�H��|�=d�`*q��h����?'?��>�쾮�D��;�����>�YG��P�՟���P0���2�ܻ�����>���2bѾ(3��S���ޏ���A�4p���>�rO?���?J�]��4���*O�������?�?��e?2�>�.?�q?�N��lk�����9�=��n?��?���?}�>o�=�k��@�>q?�+�?�'�?�o?`�M�uC�> :`oE>z䑽ܴ>�H�=G�n=��y=� �>4?�?��p��E�����J��XX�n�5=�M=��>!3�>0LN>]_�=P�=�{�=�S>v�>�lk>*e>���>�Q}>t����,���0?�0'>���>��>?�{�>���<�:8��U�=5\�=�EO�ih�jV�MG��֤;�.��"��<S�{���>�ݻ��X�?8Ŭ>O����?s/���� �ڇ�=�
>o)����>!�Q>t�>鮆>��r>���<R�o>�B�=�FӾP>����d!��,C�U�R���Ѿ~}z>�����	&����w��QBI��n��vg��j�O.��T<=��˽<-H�?�����k��)����R�?�[�>�6?|ڌ������>���>�Ǎ>�J��i���\ȍ�	hᾣ�?D��??iC���>~��>zq�>�D�h�����P��ɂ����@���{����H�[��ㄾ0m>���?���?�l�>��ۻ ��>�(\?U��k���\v>^ݾy�H���>��`����&zþ]<d�٫��X��>i�8?*i?��>m�?���=���;w1Z?n�H?Il?6Z?��/?M6B��q%?��=X�(?���>T :?��?���>�Ŧ����:�h���1:L���+J�l�(����;�	�=�[=��c<��f=����<	2+=�,����0=x"=t�G����==�<R�r;u�>zq?�a>�h^>�?�j�t�,�������&?)\��S��9澬�Ǿ���]&>��b?�^�?�Al?�4�=�K�E惾~\�=�@�>�-;>��Q>�T�>�^x���z����>���>�y�>��8��C�+���-��E̕�!}�>1>�	�>k�}>���&'>N֣�P{��b>K�R�⺾\�U�H�2���v�V �>BL?@?đ�=�龔�����e�h+)?j�;?FM?O�?���=�c۾��9�1�I�yl��Ο>�f�<F��Sݢ�%��e�:��^;��u>`O���ᠾ b>U�7�޾m.n�K�I�#��L=�q���S=O]�fM־���dV�=��
>�>��d� �g��=Ӫ��J?DCj=�R���V�������>���>��>8>�B?u��J@�����4ǘ=���>v6=>�S��H&�L�G��r=�>4PE?KW_?�k�?v"��$s�e�B����g��*.ȼj�?Hp�>ld?B>��=����%�d��G� �>���>��;�G�@���,����$�O��>x<?W�>��?O�R?��
?x�`?�*?�B?�'�>��������A&?ň�?��=`�ԽT�T��9�F�� �>?�)?7�B����>��?m�?��&?a�Q?��?�>� �iB@����>Y�>c�W��b���_>a�J?���>�=Y?ZՃ?0�=>=�5�&梾!֩��L�=9>v�2?�5#?�?Z��>���>b���s�='��>nc?"0�?��o?̈�=��?<2>I��>��=���>5��>'?lVO?P�s?��J?��>`��<�J��27���Fs�гO�a΂;��H<�y=���{Mt��Q����<�;�I���E��q��˽D�������;���>Z�x>���r�b>m���Ф����C=���1qǾ�����t{�� "�d�y>p?5�>?�)T����>9k�>(R �#.?:l�>b?p�P��4��P����E	>�Q$>l�>?�V>#����!���Z���?��E_?��n?��ؽb{�Q�o?P�L?�c��9U�����+�޽����I?���>m�;�Ϣ`>²�?l�|?]B�>�x��ңp�����N�U�	EP������<>�w���+�+I�>�g?0b�>ݏ^>��'>&�ľ<Z~�nܡ�NB�>e�~?Y�?���?�?9>u����)�d>S�����^i?qR?rBE��?�3>�3��;䍾Nq�6�޾����,�JW��:�Ӿ6����\���g�]�½f?b�K?o�^?D�@?B�"�����Zq���_��W���+�*<�If��S5�B"�h-N�a����B����ټ>?���hA�Ä�?��'?g�.���>��ض𾲌;�>A>��
|��̚=����/�B==b=�@g��d.��X��� ?��>X�>�M<?�Z[��=��{1�ɦ7�:����3>�b�>p�>@@�>)&;ɛ+�b�罉�ɾ���ҽ�7v>�xc?G�K?��n??p�"+1�����+�!�t�/�sc���B>Hj>)��>�W����-:&�:Y>�!�r�[��7w��5�	�ץ~=�2?C(�>\��>�O�?�?�{	�Uk���kx��1����<�0�>x i?�@�>/�>6н� �>N�>(hl?P!�>�g�>D!��,g �9�z���ƽ���>s��>x��>��u>@J(� �[��|��I����J9��C�=��i?]���%b��$�>�Q?jU�;�l<���>��v�*�!�����.�\�	>��?��=�<>+�þ���3�|�x��pI)?�D?rޒ�ɤ*��m~>6)"?�Q�>x��>Z'�?��>Dmþ �^��?��^?ZIJ?UKA?�!�>��=�����4Ƚ��&��K,=4��>��Z>Q5m=iq�=N��Zj\�����D=���=��ͼ B���P<�q���3K<�%�<�4>�mۿsDK���پ�	����<
��䈾%����b��ŵ��`��u��;\x����O'�`V��5c�i�����l�/��?�;�?+���O.��겚�����A�����>�q�[����������*�����>���id!�o�O��%i�O�e�G�'?�����ǿ𰡿�:ܾ;! ?�A ?�y?��9�"���8�� >1E�<.)��s�뾣���
�ο0�����^?���>���/�����>ۥ�>(�X>xHq>����螾/1�<��?5�-?(��>��r�&�ɿd���O¤<���?-�@[�A?��(����[kT=���>��	?@>V�0��-�����r�>�?�?���?�M=��W�n�
�be?���;��F�{@�}��=��=%=���8J>Aa�>�f�|A���۽.�4>��>�#�9��0^� ��<�]>
tֽ�̖�5Մ?,{\��f���/��T��U>��T?�*�>R:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=q6����{���&V�|��=[��>c�>,������O��I��T��=p�S�ƿ��$��|�c=�ܺ��[�7}������T�&#��qfo�3��&�h=���=0�Q>El�>h$W>3Z>_gW?��k?N�>��>�7�����ξ�{�
H��G��զ��L����'R��߾��	�������_�ɾ'=���=D4R�ė��� ���b�{�F�d�.?Ow$>��ʾ�M���-<�mʾJ����ۄ�X¥��)̾��1�L"n��ʟ?m�A?������V�p���l�]}���W?�P�a���嬾b��=I�����=`.�>œ�=	�⾳"3�0S�mY2?J/?+�Ǿ�ϗ�c�!>���g I=MU,?�?
=��>�)? ���j��H>;%>]��>�h�>U��=ݶ�V�ཛ�?fS?�d������G�>�2����l��s�=|>p�@��E�=�X>&�=҇�?|�����e9��d?qȳ>�4;���K�H��E��K-=3-r?FZ?~/?X=`?0�X? ��<����xk�o�(����<|l?ۻ�?&��=��=I���ý���`?H`f?ƺ�>e>�����T�%�����7?H�?UH#?�ђ��O|�/��)3,��<I?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�ٕ��Z�?��?~���LDg<Q���l��n���<�Ϋ=��F"������7���ƾ��
����ῼϥ�>EZ@�U�r*�>�C8�[6�TϿ(���[оzSq���?J��>T�Ƚ����?�j��Pu�_�G�0�H�ĥ���̏>D�>'d���N����c���7�xv����>�EK�S&_>L
����ʾ�}����<�7�>G?�͗>7���BԾj�?|��َÿ�����پ�iO?oF�?Fh?�3?[s=V�b��ŀ�I�=L�Z?��? �W?�;�3���3�4���j?:S���U`�8�4��BE��U>:3?xD�>�-��}=�>���>�>"/�b�Ŀ�ٶ�����H��?̋�?�m�.��> ~�?�r+?�\��1��bM����*���2��0A?T�1>w���٭!��&=��ƒ��
?_x0?W���5���(?�9�����G����>o
�>l���_�
y�)R��l�g��唿,��ܺ?e8�?)ζ?��߾֬"���>s�>Լ���	׾�Y,<���>�� ?������2Z<Nf��h�־�>N_�?}��?��?������+�>τ?i1�>I0b?$��{�^>����׾Bp>Vc>9t�>��l>��?��`?��?�k=�~s�5��x��Tyc��/�j�l��y�>a�X?�mC?�>�,V��9=��>gc�H���4ҧ>����
��X��>o$>%>	E��.m����?Gp�7�ؿj��p'��54?.��>�?��q�t�����;_?Xz�>�6� ,���%���B�]��?�G�?:�?��׾hR̼�>F�>�I�>&�Խ����^�����7>#�B?L��D��m�o�{�>���?�@�ծ?li��	?���P��Ta~����7�^��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B�q�1=9M�>Μk?�s?)Qo���m�B>��?"������L��f?�
@u@a�^?*�sֿ����9#���������=~�=��2>p�ٽ��=�7=��6�o���_�=�Η>7�d>��p>�(O>*;>�N)>8��k�!�q��֘����C���'u�{�Z���œv����������X'��Jý�Ҥ�lQ��+&���_��
�=�U?��Q?�o?���>�y�?�!>�����u=a"�|ǋ=/��>"�2?�L?g�)?ꕑ=�����d��8��\0���>��M �>��J>�%�>�{�>eG�>���8��H>�I>>o��>��=Lb)=@���
=�M>H��> ��>�S�>�C<>��>Dϴ��1��b�h��
w� ̽.�?f���:�J��1��{9�������h�=7b.?�{>���?пc����2H?%���w)�ҹ+���>g�0?�cW?�>����T�\:>W��֦j�5`>{+ �hl���)�{%Q>Zl?�o>��t>4:5���8���O�0�����>�{6?r谾=�)�t��C��1ؾɜH>u�>����>x�i�����as���t=�\8?\?ze��{����o�fT��3�S>[�^>�=V=!6�=bA>B.^�U�����D�M(4=�y�=��O>D*?v�1>��=���>�+��uje�)�>�KD>)�>֜;?�"?�_�*U��y<���'�{*|>��>O��>�v>�dJ�V@�=F�>�wg>�V7����
R���2�9�a>{�y��)`�N�M�E�o=����A��=��=�m轮yB��2=��r?>���岀���澓��:��J?���>|x6�mc�4�%��~���J��7�?��@5��?�J��Nd��? �?Τ���n�=�f�>RJ�>Y5��R�l�?>�֍��w��[$����?�?�§�ڄ��b��!>|o!?�ؼ��p�>l�	Z��0����u���#=/��>�7H?�T��O�G>� }
?!?<_�쩤���ȿ�{v����>��?|�?��m��=��q
@����>��?ufY?�hi>�i۾�oZ��w�>��@?�
R?a�>45���'�b�?Y׶?�?`I>���?�s?�k�>�0x��Z/��6������p=y�[;�d�>�W>g���wgF��ד��h��s�j������a>��$=*�>KE�Z4��v9�=��
I���f�?��>�,q>�I>W�>v� ?�a�>{��>�x=�n��Jှ�����0M?�i�?�B�Hn����<4��=�K���?ʉ4?�)<�Ҿ�ײ>^�[?}{?�S?L�>�j���������]���z�g<#~B>$V�>G��>pg����N>1oҾ��8��!�>{0�>J�,=�,�}�Πf<`��>�F?���>�Db=�� ?�#?͒j>�*�>�aE�4:��v�E����>[��>BH?��~?)�?>ֹ�jZ3����O塿n�[��BN>W�x?W?Bʕ>��������gF��(I�X ��m��?�vg?79彪?�2�? �??ݡA?hf>����ؾܓ��w�>X�!?���A�QN&���?�L?���>�>��&�սكּk��#v���?.(\?�>&?����*a�O�¾��<+#� DW�g:�;j�D��>��>����꒴=3>!ٰ=�Lm�DG6���f< u�=�|�>��=q-7����G9,?\�F�?؃���=��r�'}D�v�>�IL>���^?n=�w�{����bu��h�T�Z �?_��?k�?	��z�h��=?� �?9?�>�K��as޾�ྔNw��xx�u���>S��>�nm��徳�������E��x�Ž���\#�>ĝ�>�*?J��>M]�=�O�>侌�M�2�@򾽼���f��I��u1�>##��J�$~���� �o/ü�T���%���.�>v�.�+E�>�?B�h>"�>oI�>����ry>��m>m�r>5Β>�'5>��>'�>{�~�y ���O?�=���&�`�@%��@hC?H�T?���>�����;��-�í?�В?��?S3�>yc�k�0��??ծ?g@~�	?S�;{_h<�s���b����ҽ�¼P���}Ǌ>0�ֽ��4�K�O�}p���?�?a�?;�ƾ�d轿�����l=Y�?�)?z�)�~�Q�z�o�l�W��S����
[h��c��N�$�i�p��돿�[������(��`*=\�*?�/�?�}�U��U ���k�6:?�&Kf>���>+1�>}��>�,I>��	���1���]�!'��i��	�>M{?/�>�zI?�;?�P?��K?.��>���>�j��2^�>��;��>���>�8?�k-?��/?Z?v\+?Qec>{���0%��ftؾ^�?��?Z�?*�?l?����m�������h���x�w~=Q.�<��ؽ�n�B�O=/)T>��?���E�9����g>�6?�!�>�N�>����
�r��H�<Q��>`�?�ʉ>_���t�^��J��>m�?���<D->Ǔ�=�M;��<�@�=g�ƼA�=�3��Qc��Q�<G1�=�^�=�P,;���;�Hʺ�¼'�;Y?7�?[�=/�H>5������
W��/ʠ>W.�>=�>l>����{��K��G7\���t>f��?��?ߑl=�fI>&�>��Ǿ�&�+����+� ��>D?�x?�?�Zh?$�
?�7;e:��h��Syr���,��7?"!,?���>���D�ʾ�F�3���?F[?�<a���Q;)���¾��Խw�>�Z/�H.~�.��DD�.(����+��^��?ǿ�?A�d�6�w�I���V\����C?^"�>wW�>f�>.�)�I�g�%�{3;>։�>vR?4k�>��<?��n?ŒC?�S�>N���P��vߣ���߽�j�=@r'?:e?r�?J%�?�?e>~<��L��*��a!�Ķ��A���c>fI�=�Z�>ר�>�u�>�/�=O�������U꽝��=�a1>Q��>A{�>]�>��>{��=#�G?r��>7����`�vh���S��tE<��]w?D�?��*?H��<�(�5@F�i���p�>�ۦ?ݫ?E�,?`MP��>=۩����nօ��'�>cs�>�֒>g��=�I�=�1>9	�>��>ə����k;�KS\�_:?�xG?*��=�iҿ�z����Ȫ��,֯=�
�"�21D�3�6�TƑ=_�|�]�8�nѵ�7����u��U���3��ev��zȓ��y�>��d��.=k{�=.T�<��5��S=��t=.�p<6=��'R���	=�(�J��6[a���N��(<�)=��4<�ߊ�7�n?l�?u�?
��>Iݪ>���>�#�<�|?�( >�Wc?��l>�G]>�4̾o\�ڡ�%̽N����Ǿ`)������V��=��7���>�At>\�A=�F9=�	>p��8�U�=/�~����q5<a >q��=��=�3�=�y>[�s?�g�������DP�l�ս�7?�N�>�*�=",ƾ�{<?�o,>D��h ��� 
�oi~?���?�|�?N�?lSs��s�>�堾ɱ���\Z=��y��
2>��=L�?���>�$N>����M���;��f�?��@�??Yڍ�r п��,>��7>�)>��R�}�1�ǣ\�)�b�/<Z�מ!?3;��̾��>}��=�߾}�ƾ��-=�`6>�)b=���fX\�O�=1{�N�;=Dxl=�ǉ>��C>���=�7��z�=�J=�X�=d�O>6͝���7�#<+�W�3=���=/�b>e�%>p��>b?�&(?8s?�(�>���
*�������>"-V=6�`>�����=r��>o�0?��6?GL?O��>>��>�ш> �;�gTi��,������;�-�?-�?S��>~(�S�����E�80=��$�>��&?�?�A>�U����9Y&���.�$����{4��+=�mr��QU�M���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=$�����<�vż�����u&�:�+�1�����;r��;B�]<^��;~��=;��>�>}��>��=@:���G/>����Z�L��}�=vF��fBB��6d�g3~�`�.���5���B>M�X>v����/���?o�Z>-�?>:t�?�"u?� >.��I�վ�D��H1e�cgS�#:�=O|>>=�vp;�8`��M��pҾ���>,�>��>O]l>�,�2?��1x=`���U5���>����"�I��1q�X>��<���2i��w��D?�C���V�=~?b�I?�ݏ?�~�>�ɘ��wؾ�>0>�F��8=���q�&9��h�?N'?���>6� �D�CϾ�XϽ�T�>.�;�.�O�����E0��g.��m��d�>����kо�4��������z�@� 4d��,�>��M?;��?��E�%�����O�����r�d��>z�e?� �>V�?��?ܮ����\���9T�=%�q?e��?��?��>���=����;�>�*	?3��?͸�?�~s?��?��t�>��;Y� >'Ø�cd�=*�>���=��=0n?V�
?��
?�j�� �	�0�����1^�R|�<�̡=և�>�r�>J�r>���=��g=0p�=(\>?ٞ>��>|�d>��>nQ�>�������%'?1��=�T�>J0?$��>ہ]=6�����<T�N��HD���.�򄸽�ݽ9i�<^�6��-W=��ļ���>-ǿ0�?q�T>�!��}?~�p�#�LX>�U>�9���>�E>��y>ͬ>x��>��><��>�)>�FӾS>����d!��,C�Y�R���Ѿ�}z>�����	&����w��aBI��n��ug��j�M.��W<=��˽<0H�?����"�k��)����Q�?�[�>�6?~ڌ�����>���>�Ǎ>�J��j���[ȍ�hᾥ�?D��?��=:�\>�j?d�?�+���/��`�p�U��6���o�4	o�����A���3
���	��.j?��?�t@?������>?/o�d��C��>[��!�N��9&=���>�M�l������t��Ա�<��>m9�?��f?R&�>�>�� |y��G�=��6?�3?e�a?>?��C?-}�ƌ'?�s7>z?�??��3?`?u�?��>���=��S�>j�=�e��^뙾$�����Q��J�<�,	=\|g<���=R��=UD><�g���	K��$�;+��<F��<�^=E�=���=v^�>�Z?�&�>�X�>�q4?�HU�(0�G񤾁�?��<�������W���*���>(�i?��?AKY?{�^>��@��R��X>ڑ>�e>:`R>G��> ���x#���=�Y�=��*>�f�=���@P��:��r���E81U$>�8�>���>z����_>d��:ש���b>��6�)>�@Y��?���E��S�� e�>7=K?#?4ū=���
����{f�$?�\?�+Q?h�o?�������6���R��b �2O�>�Dp��`�2ߞ�0����.�1�=$"I>\f��ʔ���Y>��r�ؾ��m��1G��w�'jp=�h�K�$=:��-�ҾC�w����=zJ�=�ž-� �G䕿v`��ٱI?ue=T���ݏM���q�>GF�>%a�>EJ<������'=� ���⬨=t�>��7>G�ټf���F��y��8�>MLE?8V_?�g�?\,���s���B�$���%]��\ɼ��?�z�>�f?�&B>��=T���7�}�d��G�`�>A��>g��>�G�'0��~��A�$����>�3?��>��?q�R?��
?Û`?�*?�@?&�>�+�����A&?7��?��=��ԽW�T�� 9�F�o��>v�)?7�B�깗>Y�?�?�&?�Q?�?R�>� ��C@����>�Y�>��W�b��c�_>��J?���>p=Y?�ԃ?��=>]�5��颾�֩�TV�=�>��2?6#?F�?Я�>52�>�����7|=�"�>#!g?�Ʌ? Je?Ð> W?>	��>��=�>R��>?_?��E?�Zg?_�@?R��>+c=� ��@����#�i��<t���w�<�4�=w ��:�2���=���<A�/�3n�<�a/��7��%���?�<9��>T�u>�ߖ��.>�ž�����C>"d������������5���=�%�>$?]�>io#����=�g�>��>�����'?26?�?�&=��b���پ��N�U��>B?��=�5l��$��j�u��rb=n?��]?�=U�����ƚv?��L?2+�[�N���,��@S�M�c?_L�>��m��4�>�v?3�u?C�?0���ko�Y���5��{��C�
>t�r>7Y.�~c�m�9>�]k?N&?��>C[�>��%��S����#�R�?閗?e?�?���?�<>�JS�ݾ뿎7�^c��0>f? 5�>���#�?���U����9n���%�&n���q��ʖ���b���J�ꖾ�uǽ�PT=~�"?��V?�Z?m�[?�f�T�h�:Ba��s�{DZ�^ ����� 1�O�1�v�\���{����pž��O�.k�=������6��	�?
�?8�*����>���ᢾ�������=�������7��=����st<Q�޼���Α5�����Q�(?��>{º>�`;?�e�px:�5�(���)�# ����=TS�>��>�_�>0����@���3�����yo��@���0v>vc?��K?>�n?͈�(1��~����!��/��m����B>�>��>��W�%��~5&�:W>��r�����w��@�	�t�~=m�2?�-�>i��>G�?
?|x	�l|��}fx��{1�X̓<F;�>Xi?�:�>��>�нh� �_�>�b?`�?�>=�����)�� b��ա>�.�>x��>��Q>	|��XZ��g������� <��k'>�mf?�q��C]��$�>�#7?���<������>����}������#��93>A�?��=��>1���:3z���:�$I)?�Q?�ے��*�v�}>�"?���>��>z,�?�>�?þ����?"�^?�BJ?�KA?�#�>�_=���[�Ƚ��&���-=2��>&[>�m=2 �=�}�'d\������C=Sں=�.ϼ$⸽�<Im��[�L<ֱ�<��3>SۿWBK�(,پ+�����
�U�~�������=�W���E���w�����>&�5�U��c�C����m�Oh�?���?j/������Ԣ���q��'��e�>�jq�Qs���2��}���Е��x�����~!���O�5�h��e�P�'?�����ǿ򰡿�:ܾ3! ?�A ?7�y?��6�"���8�� >uC�<�,����뾭����οB�����^?���>��/��t��>ܥ�>�X>�Hq>����螾�1�<��?5�-?��>Ύr�1�ɿa���{¤<���?0�@�}A?�(�j�쾍�U=9��>�	?`�?>MV1�HK�����\\�>�:�?c��?i�M=t�W�Z�	�\}e?<P�F��޻w�=TR�=�=����J>�U�>]���NA�Z%ܽ�4>,م>�o"�޴�n�^�Lվ<�~]>�ս���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6��{���&V�}��=[��>c�>,������O��I��U��=��t	���G)���	�J�='p`=3&;�J�����[�>Qܑ�
�c�S�>=�&��k�>)zf>�n>&�=):>�S?��b?)�=>a�>�#ֽ
�!�N/�����������Ѿ�O>�����[��N����m�����ʾW���i!=�?�=r6R�痐��� �P�b���F�b�.?�v$>�ʾS�M���-<�nʾT���xބ��ॽ0-̾��1��!n�3͟?m�A?������V�1���S�����q�W?N�/��묾'��=|���o�=�#�>I��=&��  3�Q~S�f�0?5k?Ft��m:��zH#>�����==X�(?
��>�y�<�r�>0�$?g$�|mؽ4�^>�3>�B�>W��>9�>��� �ֽ!�?��U?����P��滐>����s�bb=�/>��/��k�HX>��<�ۇ����7R��{��<�(W?u��>��)��xa��k��Y==��x?��?.�>j{k?��B?dդ<$h��|�S����aw=�W?0*i?��>����	оW���B�5?�e?~�N>�bh���;�.�[U��$?�n?5_?�}��'w}����p���n6?r�v?�,^��_�����U��ԥ>���>���>��9�
�>J2>?�#��h������K4��؞?N�@���?�V1<$0�M�==?��>�YN�L�ž������=u=z��>L茶�Ev�)��.,��\8?/��?���>4��������=&ڕ��Z�??�?����Rrg<��l��i���;�<EΫ= ��H"������7���ƾ��
�0���]������>Y@pc�-*�>�L8�~6��RϿ���,aо%Kq���?�|�>��Ƚ������j��Ju��G���H�Ȟ���z�>$,#> ��8���J�-�T��ć=-=�>�$ʽ���>bfƽ*R����z����=o�v>*�>*�4>��K��t���ј?X����տ�������j?jƫ?��?�L?�=��򀾴5���=��j?5ݎ??�W?�D������3�s�%�j?�_��xU`��4�uHE��U>�"3?�B�>T�-�g�|=�>���>g>�#/�x�Ŀ�ٶ�>���Y��?��?�o���>r��?ts+?�i�8���[����*�M�+��<A?�2>���I�!�C0=�UҒ�¼
?U~0?{�d.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�0�>O��?6�<3`�> ;�_�s>ne�;�=�=��9=H(?��G?���>cOS>��������9�ԾA����`F���>��n?��]?f�>G4���ѕ�k�
������*�(�&�I�	co���>���;>`O�>� >�������?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�	?p��>���E~�C��VP7���=4�7?�K��z>l��>)g�=Ksv�8�����s��ض>>�?'}�?��>�l?Mo��B�+/=���><uk?qT?�r�_�n�B>��?�����S��f?��
@�y@;�^?��`¿	z������Uۜ�O&�>��=��>2��=n�E�v��=RS�=	�;��ڃ>�S�>��>���=�7>1��;�@�>Lm|�0�%�������)�;���~ؽ��h��a��������u6��Ņ���<�M�J�7����u=���=��d?b�F?�6r?�E�>�����w>��Ѿۓ �鴾+z>� �>e/?`�Z?��>?�
>S���'�Y��ep�-��O����ſ>3�>i��>͊?�4>Õ�<٫	>wF�=f��>6�'>�H="�=t�=1>υ�>M'�>�f�>t�b>�>�ﵿ2�����r�Tc�nO1�� �?����f�N�q����r�'����>�7?���=�&���dп<б���A?핉����@�U>��3?2ZR?H�>���Մi�c�>�����{� ">�����U�� ��8i>� ?k;g>S�u>�3��h8��P�X���K*}>p6?W
����8�qIu��wH���ܾ��M>�ܾ>�aI��_�Y���i�|=	�:?k�?�t��Mݰ��+u����®R>1�\>�]=ba�=>JM>We�.ǽ�&G��,=�T�=��_>i?I�k>�
=N��>�w������L��>���=�'>42C?Y�3?�g;;�C�M��J���>�*�>	�Y>�>vr�/�=�w?�e�>�~���������u�;�`�>�'ؽ�����U���=��&�'�>���=��O���G=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾXh�>ox��Z�������u���#=V��>�8H?�V����O�E>��v
?�?�^�੤���ȿ6|v����>W�?���?d�m��A���@����>8��?�gY?�oi>�g۾a`Z����>λ@?�R?(�>�9�r�'���?�޶?̯�?%Cb>�ʃ?���?��>m�'�Rv%������x������=�>э�=m��t+C��7��)���^j�Q�ϾE$�>��^=_��>8է������:>S�B���ԽD�|����>�r�>���=���>���>��>�@>E��� ��"����ǽ>hj?c��?lM�O��%8½�L=OLF>�& ?_k?V��<�����>s�J?An�?ԑ�?r��=U<�xۖ�ܷοo�ؾ��\>wDU>�,�>*!?�_Z�%��:���YҾG��>�.?*G�iճ���g�>�l��>�?���>��>�<'?"�?,B�>���>��A�p����!��۬<�{�>��a?.�]?�J?����y�)����@;��Akm�/� =e�?0j3?T�p>U+��TR��׮���O�1��>Jr�?�!?��B��I?��X?�Qn?bO\?'!�>�ד�bo��,�ɾ�M*=�"?����B���&�K��p~?>�?���>�x���%ٽp2ؼBV�'����r?��\?k�%?R��ha�Pľ���<���,�m�D>�;	�0�j�>�k>�ň�� �=N�>룱=��l�i7�^�k<��=���>���=ߔ5��א��e1?Y�<��]����=��g���E���=��1>���ׁ??mn�j]v�zԯ��a��.���"��?J��?��?O}ֽ�ok�6�5?զ�?�J?;��>�R���M˾M���U��L��ԾK��=��>tj��c��Z���4���n�m<�a����>�M�>��?� �>6U>2��>������!�"������\U�0�,O1�Z�.�� �;F���0�4��}w���>n�V��>����#ӫ>`?4{>5�>f��>i����p�>��E>y{�>�M�>�v>��$>u��=]���w硽!FS?w��)�_j�G�����A?��e?��>�J������T��4 ?/D�?�?H>��g�]+�w�?���>�$��,�
?��3=t�Z����<�J��\�X���#��=ٍ>��н;9�e"M�ޥd�s�
?J-?]���ȾU_߽M͓���=P�?f$?q)�=|Q��;m�l�c�5�I�;��]Ox��ɗ���'��m�u ��ް�� Ƅ�9� ����=�c)?�:�?g���,� ���Cp�ܶ-�&�Q>���>2�>���>�nE>i�����-��^��!�K������>(`{?�,�>�BV?!�2?��Z?�|5?}��>��>���/@�>�����>��?�6?�P??�WA?*?pD?��!>�� �8D��©ݾX�
?�o?��?�@?hW�>^&`�i�Ž?�������Tm�
�1�h�=�&=q)!��KA��=A~_>IW?<��L�8�?���=k>g�7?x}�>'��>���3/���I�<]�>/�
?�E�>x  �xzr��a�1R�>���?����=��)>���=X�����к�Z�=�����=�4��Dt;�E]<r��="��=�qs��v��>�:J��;"��<�=?��?�6>�>(��&��A`Q����#�s=���>�/��R
��	��Q6���6�[��>b�?�B�?p����>�7�&�-�^V��"x2�[�� Z�<���>�G|> �6?���?=,?�Z"?��0>�Ʋ��ꚿ�]��OҾ�x?�-?��>�>���Ҿ_y����4���?R ?�rc�2�"���໾×��6�>�P(�YF{����!D�����z.�v,����?L��?�����%7��Oᾢ��Ȧ� �E?1��>��>s�>Am,�ߛg����.>�N�>!W?��>��O?�6{?Y�[?`^T>a�8��%��Ι�3t4���!>d@?���?��?y?1��>f�>�)���I�����<�3؂�C>W=�Z>欒>I�>��>/��=��ǽa��?�>_�=ؠb>��>b��>��>�w>"�<�$D?�h ?aȽ����*�$�2���^����]?��?W�?|��g$� l��N��!�>=��?�?�>J?�����=�cW=2̾CE�����>R��>�_�>� �y�8>[��=��>���>�������S�@�
��?��%?�y?=�$��P�b��^��Q�$�\sG;��ڼ(�N�o����w"�|�j=
����E>�ý~7�zX��$䂾����݁�Bv���>;�g>���>�Q��g�	<η�<L�=���=���=:�q=\8;*:h��R���њ=���>�������"�=.�U;���}?a?7$V?��&?[�'?ߞ>���=��=�}�>?����I�>�S>>�:Ի�����.�����s߳�)�����k4��.����>�2(�>>;�U>4 >quu=�>W v=�s>��˼��$<q��=�>���=��=?#>�P>�6w?��������4Q�&X罌�:?�7�>�x�=�ƾ�@?��>>�2�������b�X-?|��?U�?y�?�ti�e�>@���⎽�t�=�����=2>���=��2�D��>��J>���J��;��]4�?��@�??�ዿ��Ͽ�a/>�}7>�>n�R��v1�Y�\��kb��Z�9�!?�6;�L̾)�>E�=�߾��ƾ��-=.I6>��a=�w��R\�e��=q�z��<=�k=?ˉ>�D>���=������=��I=#��=��O>\����6�v�+�"�3=���=��b>�&>���>��?b0?�Xd?A5�>	n��Ͼ�<���J�>W�=�E�>��=KrB>���>��7?;�D? �K?2��>~��=
�>q�>��,�Գm��m御ͧ����<�?�͆?�Ѹ>��Q<B�A���kh>��6Ž�v?RS1?Dl?��>���ݾ�|�C�,���>�ݶ<���=�HX��>���>m,�t1;��>?�=^ �>�M> >� ~=@P�>�>n5�=�Z�=�Ǔ=7���=w�=�s�<uP���>�ݻ���WT�;"M����O�Q>i�<�#���*����=$��>�`>n��>Z��=������,>�ʖ��M�C�=�7���-B��Yd��Y~��;/�&�5�PB>WnY>�샽,#���?��[>��>>�4�?@*u?� >��Bվ��ϋd��cR��J�='i	>@�<�s�;�1�`�y�M���Ѿo��>���>%�>T�l>A,��"?���w=��a5�Y�>�|�����/��8q��?������Di��-к�D?_E�����="!~?��I?3�?���>}����ؾ5?0>~E��q�=�
��$q�-^���?A'?j��>��S�D�픴��5ҽnv�>���I\��w.��锺�㲾*`�>����Ҿ��,�����eڏ�$l=��"~��]�>��P?2�?r��[9�g�H�� ��R6�(��>l�C?hRH>��?ŧ�>�����	�q���(��<���?:��?pH�?Q�>��=Kc��ߙ�>X�
?���?���?ZQr?X�:���>��C;�$>:�����=��>���=ȕ�=n�?��	?)#?�P��u��9G�h��,�Y��_�<"t�=�ݓ>7�>iq>���=?Gu={�=�[> @�>���>P�c>���>7~�>~ݦ�_S� 4'?� �=�]�>/2?��>t�g=�D�����<6gT���>��;*�ƣ��T�߽K��<|�˻]LL=�HݼA��>��ƿZ��?7�T>�B��F?)q���z,�xYR>��R>��ܽ�E�>�D>laz>7k�>[�>Q>�Љ>
�'>�>Ӿhe>˻�	V!��(C�-oR���Ѿ��z>E����(&�ܜ�K{��L1I��b���b�Nj�.���6=�]�<%F�?ѵ��-�k���)�����?Q�>\6?J������>���>���>*\������	����Vᾱ�?���?���>)��>^�F?*�>�T�2;�/f�eiJ�.sP�F�F�F[_�1]������,9��-a�O�?TT�?]-�?$���4}>Ub�?�|>�\.�XJ$??#�IX:��1��Ԓ>�G��K��&�=AH�1P�<iv>��?�a�?7�J?�2پ��(�!�>�N�>�kv?:`?�~?C/?�Լ<�PP?nZ���t?`�>�"?;C8?4
?7�'>7>=�܇�\��>*�*<Z:n�hF�zڧ����ň=X�̼��&=�>�0�=��i���?�@"ǽ�2��0Ͻh�Ȼ1F=�>i.�=�ֱ>��h?��>��>4�P?Ǌ ��jE��3˾��5? � ���ܾj����龯�ac�;L�?lN�?D�p?��=ǂ��VE�#�=�p�>4 >���>�H�>��5�S/���"0=��>�.> �m>�2c�)ѧ�ʮ
�gׂ�����&�&>���>p�|>x&���'>��lz�A�d>��Q��ʺ�6	T���G�-�1�8Rv��t�>n�K?�?�h�= Y�a}��NGf��+)?�_<?�WM?;�?�@�= ܾ)�9�J�J�-�����>9.�<������3��[�:�z�:8�s><(������3%>i�ܾ�vҾ��^��?�����k<)��CΔ=Ҡ��M��"��nu=��=��ؾQX&��o���2��<�N?� �=��z�EVk�������=���>�ړ>d���<���6M@�CNȾVf=FS�>~�K>|�	���
�u6N����j>�>MQE?CW_?k�?"��Hs�/�B�����zc���ȼ(�?�x�>�g??B>��=������U�d�yG���>���>?���G��;��N0���$���>R9?c�>��?:�R?��
?h�`?�*?+E?�&�>~��o����A&?4��?�=p�ԽT�T�� 9�`F����>_�)?�B����>�?��?��&?1�Q?�?H�>� ��C@����>�Y�>��W��b����_>t�J?���>N=Y?�ԃ?�=>I�5��颾'֩��V�=>}�2?�5#?"�?į�>�R�>8^ �=BF�>?`?���?�4_?4>x�?!;=/��>��>���>j��>þ�>ƒ=?+�i?S�a?-�1?ˎ=�i�ղ�����?�K=*H�='7��ʑ=�_3�_,���^�/�>�[6>w@�:�
�=����b�+���<�ŕ>��>ivt>M�� P.>�ž{��fB>� ��[Ԛ�d����9�43�=��>�?�>G�"����=ɳ�>���>S����(?:�?�X?��;x<c��/ܾLK��>R$B?�U�=�/m��S���v��a=|dm?Y�^?W�����u�n?��H?����s@�m�������f���s?�I?o8����>�v?i/�?��?��c�7�p����d�_��W���#>�;:>?h;�ۑK���/>R`?,T0?#�>�c�>�+��H��#A޽1g?�T�?{l�?��?R�>�7p����4�J����K^?T��>� ���I?�W�jV̾�ӌ���l��߾Χ������uT��1�H�"u����1�=��?H2s?��x?�\R?���n�e��,Q��s�l8S�D{�� ��AN�ΊA� �<���h������
���ľv��]퀾�vA�o��?��&?��.��]�>><��ߠ�$kϾ�D>.g��D3�8p�=sA��}�(=�g<=�o�"66��Ա��B ?�.�>Ri�>�k;?0�Z�N;=�*�0��7����5�4>,�>���>7��>�E��,�I꽽�ʾ*2��)ֽ
$v>t�c?�yK?��n?"E�?1��d����!�א-�D_���C>e�> ܉>2W�#O��&�0T>�M�r�B�������	�b/�=�2?��>e-�>�?�?�?p	�9���iux�<X1�6�~<�&�>i?���>`ކ>sϽ�� ��w�>2�l?@c�>��>'X���!�C�{��нq�>�3�>'1�>�q>��1�T^\��/������e�8�,��=�h?v����5`�CO�>b�Q?�yN:��:<1_�>m���	!����Rw%��K
>�Z?׫�=�p9>{gƾ\��z�Eʈ�kJ)?�k?1����$+�$o�>�a!?��>���>��?骚>G	ľv�$��?��^?��J?:�A?!=�>�@=xɲ�>ǽ�&�/�.=�߇>Q�Z>x�i=���=~��g[��T ���H=JB�=f�˼P��f�<Z���C<<�^�<�83>D�ٿ}L�a�ƾ.[	���>����x��N����h�8ȷ�@����}�Ͽ!�]C��C�g� �a�����p����?fH�?�}�������������/�����>�{�	J��;��N�.�����!ܾ|ī�
�"�"MV�io�n�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >[C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾w1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@|A?��(�:��\�U=���>��	?,�?>�(1�A�����j�>9�?���?c�M=p�W���	�{e?��<��F�IR߻#�=�a�=9�=���yoJ>�A�>��-fA�Eܽ��4>Fօ>�M"����$�^��N�<�r]>��ս��Ԅ?�x\��f���/�2S��QN>��T?=+�>�4�=ܮ,?x7H�*}Ͽ��\��)a?1�?,��?e�(?ۿ�>֚>;�ܾ�M?&D6?T��>Be&�?�t�׀�=V�ꊤ����q%V�)��='��>�>�,�ʋ�P�O�fS�����=����ƮÿZ�	��(=���=�.��V���=��<�=;�~���N�����6ܻ�$F=�>`�>���>@��>�L_?j[b?�l�>�eP>����话��*˾��f=﬒���O�)����i��f��O~��^�����R�nS%��뾚=�U�=�5R�1���^� ���b�טF�R�.?�p$>5�ʾ"�M���,<	uʾ����D]��Rƥ��$̾��1�� n�!̟?]�A?����f�V�h��Z~�����ϫW?G�+���鬾��=A����=�'�>V��=���"3��~S�Qd0?��"?e:Ѿ������?>�q'��3=�,?���>f��<��>�Y?��)����=>:�!>Š>r��>6�=����	ڽ[�#?�KZ?T=�OK��9q�>�/־�]�Yk�=�O�=�6���ܼG#]>E˹X�����O닽�	�=��V?�%�>#@)�<��~z��u���F=�x?]�?���>DCk?�'C?'��<Q���,�S��0
�^ځ=�{X?��i?�~	>����v6ϾYG��Uk5?��e?ГM>��f�v���$/����x�?�o?z�?�鉼9�|������H�D6?��v?4r^�s�����)�V�)<�>?Z�>���>6�9�>k�>C�>?�#��G��躿��X4�YÞ?��@���?�;<a����=:?'Y�>��O��=ƾ���������q=��>l����dv���.O,�ĉ8?���?ĕ�>����۩�6��=�ٕ��Z�?p�?y���gBg<^���l��n��k��<Gͫ=��I"�I����7���ƾ��
�����忼ƥ�>,Z@U�Y*�>�C8�46��SϿ!���[о�Rq�w�?l��>ġȽ����-�j��Pu�Q�G���H�f������>�|>a��C���	�|�}�9�@Ck��{�>�@�2c�>"*H�X��������R�<eS�>5��>}w�>�X���R��k~�?�����ο�Ǟ�8��8Z?���?2Ԇ?J&"?��?�|���r�:�:kBK?>su?O�Y?P�?�i��}s�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�d�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�0�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.���_?΃a�W�p���-�{�Ž���>�1��%\�~������@]e�W��A|y���?�`�?��?�K���"�2*%?	�>����}/ǾT^�<r��>��>9N>��_�{�u>
���:�\|	>���?w�?~g?e��������*>��}?;N�>O?�?�����-�>չ6>�f�$�=�W�=�_y>��=_�6?�x-?D ?��>E��k^��v1���N���ʾ,�7�vs>.C}?��h?�!�=UNӽTg����/���B=�41� �B�k�m��Ľ|�$�x�k>���>`��:��Y�j`Ͻ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji���?������Lty���CQB���=X_4?�9��GN�>�>�H=@w������s�
ٽ>(�?��?��>�}l?dhh�`�G��f�<�
�>��h?��?V�=���@M)>��?�B�7����0��8Ik?�[@\h@�%_?����ƿ6ӡ�s����7�[�=륙=�Z>�A�1�{=�e<>�͓=���=d\H>���>k�>!�
>2=5>K�p>�m�> +{�]'������.���\A��E$��`߾:>O�����.��O	� ��+X��+�w����U��}��	��/�����=u�U?��M?�(t?���>Qm���.>'3��y�a=�~��o�=��>$�1?IqP?�P(?�w=]N���`�Rw�m8������;�>�I^>�B�>Ů�>/E�>^V��i6>x�3>�>�>��<�I
�Q�=�tC>뚧>O��>Dֻ>I�<>�~>?ϴ��(��Яh���v���ʽj�?=����J�=5���	���w���L�=,g.?.b>-���9п����*H?0���0�=�+���>��0?�eW?Sz>̰���U���>v���j��Z>���@l���)��Q>�P?��f>KTu>;�3�nd8��P�1���#�{>�6?$涾��9�H�u�{�H�?�ݾ:TM>��>h�7�<��񖿇
��fi�4�z=D�:?��?���L����u��g����Q>y\>9=Y��=� M> �d���ǽ�[H��,= ��=�|^>W?�5>UWw=t�>
r����[����>�?A>��.>(@@?��'?ǯ������3{�PY3�hr>�%�>E�w>�I>�dM����=���>�l>��+�����dK�{+_>R�l���f�I'b�3Mx=}��X��=\��=5��48��Bc=<�~?|��5䈿��cj��>mD?�+?�=Y�F<܃"�S ���G��7�?q�@m�?��	���V���?y@�?m
����=&|�>(׫>�ξ�L��?��Ž�Ţ��	�~+#�dS�?d�?Q�/��ɋ��l�}6>�^%?��Ӿ�h�>x�eZ�������u���#=K��>�8H?sV��z�O�A>��v
??�^�ߩ����ȿ8|v����>;�?���?U�m��A��@���>/��?�gY?Nqi>g۾`aZ����>��@?	R?�>|9��'�f�?�޶?���?ўJ>>c�?o�s?7m�>(Q����)��۱��8��S8�<��
=A�>�E>���rJ��U�������a�O��V�_>��@=���>W��XP���r�=rJ���ጾ�̰����>���>��[>l�>�?2��>o݆>cX�:?A����C������S?��?��K�����>:��;�5���9?�V*?\�=�u�D���>�`?Qq?�T:?�K>��Ѿ;���6)���EоB�9>��v>��>?�x2��5P����U��>��?9_�EþC�b��7�X;>\�?���>��>+d$?P�?Y��>��>�R������.���>��>�E?6p?��?(C����'�"3��L⡿_
^�!\�>�og?8^4?�EK>g���O���ʈ*��A�<�>n��?�vw?��
��{ ?:�W?XM�?�'{?�.R>jFK�(�ھA��>��!?��5�A��{&�>��PA?Q?D��>Mْ���׽x�ۼ���������?^\?o&?R�da�þ���<��"��M��<�C��i>�w>������=1�>�j�=��l��6���k<&i�=�>�O�=Q7�͎��;,?�F�1΃��=�r�prD��>I@L>%����^?n�=�E�{����hx��r�T����?���?Qf�?�A����h�<=?s�?�
?��>@@��]o޾T��Uw��Dx� s��">r��>�p�\ �H���˖��Y=����Ž�@��Y�>���>
r?���>��K>L��>����K(�B��33���[�]�F�9��,.���b���u�����Q_��&�w�k��>Pf��G@�>l�?�9m>s�m>m'�>�/<�̍>��\>� y>f�>�P>'Y$>�x�=;��<�����n?=ɟ��CY�h���-��I}?�m�?�`7?���>Ὂ�p6�<�F?<9�?Ex�?y%�>,5�
�3��R�>�w�=�n�׫?~ܽP�6���w>�T̾`���o��hvL���>�@=�`)�v�D��оH��>c�?O�D>JĜ����Tr���M�u��?�?�!&���3���U�wxs��mh�[*�=�����.վm���������O��_����k6��R���L*?�d�?+H�RC��1�侠LM���<�Ĕ>�B�>.�>��>�w�=��ix/�:�O�� �����?e��?qR�>�R?*�3?�.]?.�>?�?>)X�>����:?�?ؼ�T�>U��>H�6?&,?�2*?�*?�w?	C>-M��z����H׾��?+s?�?�?K� ?�0����ս��v���EX�:��O��=R��=���7(?�B�v=!�$>��?X@�6����w�}>��<?T��>l��>ꏄ�����T��<�a�>36?�c�>� ��n�@	�}-�>��?����=�T >>�=V]�	h;M�=�e�ދ�=��Z�0�]�T;?F�='x�=�@ڻ�:���&�:��9M��<��>u(?t:�>��>-�qt�&(�{䐽�P�:�{Z>.�!<K���jf��l��6U��.<�kh?#�?3=��=&r�=+�0�E�}�-Gݾ���`4>�>En?sBt?��?��N?�[?+��=�c�ґ����t�h3����#?� ,?i��>���ֱʾ3樿(�3�ِ?s[?"5a�Q��$)�Z�¾��Խݱ>PX/��#~�*����D�~�������u�����?ʿ�?�;A���6�[q�����M��
�C?��>]�>=�>̺)�s�g�B'�=;>͇�>5R?!�>��O?�8{?B�[?*fT>��8�,��Wљ��<2�h�!>�@?���?p�?�y?*s�>��>�)�\ྎJ�� �`�ւ�'@W=�Z>+��>�(�>0�>���=Ƚ�b��j�>�2=�=	�b>i��>-��>��>�w>'�<��D?6��>�-վ\�(��<�a������b�v?,P�?:�	?"�G��$��OO�u��4?0�?�P�?��?��X��d�=�(N������V�:�>��>ŉ�>���<W��=���=�c�>j�>�������&����[�>��.?�0m=∲��gg���=o���/�<�N����B�)W�9�����=Nܾ������������鸾� ξA�����}D�fo?>��=*�/>��=z�a��'*�(�+=4���(Һ�vE�=!Z�<�#�7xH��0��3I��<!N��aY=I\���qʾk�}?5�H?,�,?N�B?u>��>��9��>�����H?�Y>e[E��C��k�8��r��Jו�sؾ��վz�d������	>B"D���>6=>�M�=�jg<�e�=�f=,�=��S�yk=��=x��=4L�=���=�J>I�>�j?\sF�ϒ��Jt�85=�G?��O=-F�>I4�E�?4�¼a���<���]�V�?
v�?c��?��?ՃD���>�0(�ݒo�/�%��01>�=͔�r&۽�i�>��<X��/s�Q���V�?#@�/?2�w�I�ο�:\=-89>_1>�S���2��OT�g�W�_���!?�:��XξaX�>S)�=�ྨ;ƾ*ZQ=�E=>��|=(^��[���=� y��<=$br=�"�>�C@>ѹ=~���Jƻ= �>=�9�=��P>�\��u,��(���6=�y�=��_>�=$>x��>n�?�a0?[Xd?6�>�n�3ϾG?���H�>Q�=�E�>T߅=rqB>���>=�7?��D?��K?���>���=x	�>��>T�,��m�m�Ķ�P��<���?�Ά?�Ѹ>r�Q<��A����g>��-Ž�v?RS1?�k?��>VW�u ��!�̦ �A/ ��`�;���=XX���Ѱ�G)X=r�p@��}/>�E�>倦>��>�S>��t>�t>6۫>�X>
g�<�N�=|�<�$>�B��Ub>�³�Y�;C爺�Y���\��ν�횽��ۼ&�=�@�=��e��=2��>�R>z��>�F�=�����.>ɳ����L��z�=�V��V&B��:d�BO~�X/�U6�D�B>�@X>.����0��[�?��Y>1{?>R��?Y6u?��>�9��վB��Z/e�8�R��~�=]�>](=��;�+W`���M��XҾ6��>�ߎ>��>̼l>},��"?�)�w=$⾈b5�?�>'}�����,�:q��?�������i��5Ѻ��D?UF�����=:"~?ðI? �?&��>�����ؾ.;0>�F���=H��*q�*g��3�?�'?���>�쾯�D��c��+�����>k�k^����L"1���g����7�>Ȏx�H��"�2������ܔ���1���q�y�>��H?�©?ԅ��ʁ��<��C��f�����>��z?P�>��>�?t�u�����V����=ږ�?�?*-�?��j>��=�U��,��>D�
?���?ݓ�?߮q?7�b�>t�J�c*>�d�5��=!i>��k=���=�9?_p?�?}������쾩�ﾔvS�/�==���=��>�v>��X>��=�6�=gd�=�V>9��>�>F�S>+��>��>Vg�������&?Lq�=(Ǎ>@=2?Lx�>�4Y=�:��P��<��I�u8?��9+�c%���0ώ��<�c��*�P=g̼-�>
�ǿ�4�?��S>��w	?�V����0���S>�AU>2�޽���>#�E>�>}>p�>E�>�;>�l�>�'(>jAӾD�>i��V_!��+C�C�R�e�Ѿjqz>m����&�������OTI�\x���f�g	j��,��9=��e�<E�?����k�g�)�7���ݑ?�[�>o6?*ٌ��؈���>��>h��>�L��ݏ��@ʍ��gᾴ�?���?���>٭�>L?8�?�X���n���W���P�*�Q�U�A���K�ο������	����#q?Њ?�i?�̆=���>>Yz?�6F�+p׾��>d+��-:����>Xh�>��Ss����Ծ�[�rc�:?�>���?xp�?5{?@w��>Լ���>�<?�U?8Y?�M?<�1?D��U2?ȱ1=���>yo ?@�9?��L?�g�>�\="�>�h��@ږ>����k����J����V�*��=�Q%>rB�����5�=��>+&W� JQ��Ix���=���t�Ƚ�0=�?=tZ>2Q�>:[?���>�ۄ�-|g?�!���_�<uK�'5?�ќ�����Q�-'��ι�?*-�?�'�?]"?���=����y^�Qk�>/C�>7t5�}�f>?��>�؊�r�=��[W<��`>�4>6JL=�k�;�l������<��u��v1=�?�H�>Ȗ�;>/Ǳ� ʁ�3�����O��׾*�ӾuF��b=��پ�'v>(�P?�6?�!>׾J�^���O��?�I?w�_?-?��4>6ֱ�y�%�s�G���=�
l>5N>����͇�� լ�%�m��k��5�>�0t�	;���a>NB���޾rn�� J���羈RM=c��7W=4Y�:־.��� �=�X	>6���� �L��f����&J?�Ql=�S���tU�W���1>���>��>�q:�p9x��w@��b���p�=7��>}j;>����}��\bG�P-����>o�E?˨^?hZ�?����Is��iA��� �`���ͼ,�?��>�$	?IE>��=���\��N�e���F�@
�>�8�>�����F��������:�%���>��?�>=�?r�S?�c?�a?��)?W2?��>,��������A&?:��?�=4�Խ$�T�� 9�8F�U��>p�)?F�B�ع�>\�?�?�&?�Q?�?B�>�� ��C@����>�Y�>��W��b��]�_>��J?���>z=Y?�ԃ??�=>F�5��颾�֩��U�=�>~�2?6#?W�?�>�G�>�Ρ�:<�=!&�>3'c?b��?i�n?�"�=��?w2>�E�>g[�=j�>l�>J?��N?�Vr?A]J?l�>�2�<9h�������t���@�qs;|i4< xo=����t�����<ο;;e�Kg� %�XD�������;0B�>!Gt>�@���u/>Cž���m�C>�&���v���d��S;��c�=�[�>1L?��>��"�9ۏ= �>���>��,')?8?k�?)��;X�c�|1ܾi�M�:��>#C?�!�=��m�:����v��>\=h�m?It^?"Z�������|?{4T?�{=� �v��S��-ƽ�N+��}?o/ ?;�w����>@�o?�l?,�>�'�ei��Z=��u�V�cJ>�>i@>� +���*�o3'>�u�?��??a�n=x�>~�)������5�=��?lW�?<��?�?ݞ>~z�U�ѿ�-!�����h?� �>����у?�G����Ҿωžw��Պ��7��\�о8���ܰ�����y�����>�m4><%?S]u?N��?3�U?V���]�n�ѧH�F`�u�O�7����.�8�e�HwI���V�0���-�ӱ�ُ��Qֹ�I��E�A�?z'?zx0��R�>m☾E��2{;f;C>����0�h�=�|��� >=�V=�h�%/�]%��p ?�W�>�>r�<?��[��
>�.�1���7�����x3>Ң>Z�>0�>��:I-�bT齩�ɾʊ��q�ѽ�8v>^yc?j�K?�n?�r��+1�Z����!���/�c��V�B>�m>ƿ�>H�W�L���8&��Y>�(�r�U��Ey����	��~=�2??(�>Ნ>�M�?@?ky	�On��Khx���1��9�<�3�>�i?S>�>:�>'�Ͻd� �|��>��l?թ�>=�>"���nZ!���{���ʽ�%�>a�>��>v�o>T�,��#\��j��%����9�!v�=�h?􃄾��`�6�>�R?6ۈ:U�G<*|�>A�v���!�b���'���>�{?헪=��;>U�ž5%�W�{� 7��sO)?�K?�璾T�*��6~>y$"?���>K,�>:1�?�)�>�oþV-B���?�^?�AJ?TA?[I�>i�=}���R=Ƚ��&�'�,=���>'�Z>�m=T~�=����r\��v���D=�q�=�μ�Q����<݄�� K<��<��3>�gۿ'�K�'�ؾ��t��B
��'������g�����6޵�V��vRy��Q�v%*��`W��c��򌾳�k��j�?�?}Z��w���}���񖀿����b��>�r��������� ��1[�����_��q�!�d�O��i�0�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >ZC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾y1�<��?7�-?��>Ŏr�1�ɿc���}¤<���?0�@}A?9�(����TV=��>&�	?��?>�X1�J������R�>�;�??��?�|M=��W���	��~e?6'<m�F�!5޻]�=�G�=�Y=���<�J>AR�>���_QA�Fܽ��4>�܅>��"�M���^�n|�<ۂ]>�ս /��5Մ?+{\��f���/��T��U>��T?�*�>N:�=��,?X7H�a}Ͽ�\��*a?�0�?���?$�(?;ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�ۅ�=�6�w���y���&V�w��=\��>`�>ǂ,�ߋ���O��I��W��=�� �̿I����(�["=�5=�+��]���"��@�<�ْ�-�4� ���I%=-� >�N(>kGm>��>�r>jqX?�b?{��>>�>K��� ��~ʾ�9�����`t��<����H�ofξu��y��#�����Y���� =�=�= 7R�n���� �m�b�k�F���.?�v$>v�ʾ��M�˗-<�pʾ����,����ߥ�C-̾ӗ1�5"n�`͟?��A?������V�X��iX�"���F�W?jP����oꬾѣ�=���l�= %�>늢=���� 3�i~S�7�0?H?�@��R���?�'>��s�<څ,?A*�>�<�ϩ>�w ?� (�%����V>�'A>༧>qL�>b]�=ɩ��*~��?�W?� ��[��ʕ>����;���#�=(�>7�3��rƼN$^>��Y<����$ɼK䏽` =�x_?X�>Tp1�UB.�k�� ��z=���?7��>��>m�s?5�-?�3=��/4S�&i+��P�:_�O?��?�&>�缅o�&\ƾ�K? �l?K�>�G"���־�?D����q�)?�}|?�v+?�=��n����&+#��<?Nor?�}S��i���D
���5��ؚ>(�>x�>�-��$�>�F3?�7>�٪�����B�9���?�@���?^�ڼ���	��=�)�>��>�'�hۼ�
�Ͻ8Bľ)�=���>�w���n�����h���2?��???�(��QX����=�ו��Z�?��?<���Rg<���*l��o��٩�<�Ы=� �jv"�����7�e�ƾ�
�����Ϳ�6��>tY@�Q转$�>|D8�)5⿅SϿ����Xо~Sq���?��>J�Ƚ٘��_�j�Su���G���H�ۢ���[�>��>L����	��w�{��i;�����F�>����>��S�?$������4<��>���>?��>a���aս�5?�f���<ο7���Ƞ��X?�i�?�j�?�v?O�7<@�v��e{�����1G?m�s?�Z?gW%�]0]�&88�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�w�_?�a�{�p���-���ƽ%ܡ>��0�;e\��F��Ф��Xe����@y����?K^�??�?.��� #�j6%?�>��8Ǿ��<��>X)�>=+N>AH_�W�u>��$�:��i	>���?�~�?ej?˕�������U>��}?�C�>�7�?�.�=�6�>&��=�h���I�(t>^��=4�B���?��M?���>z��=�v6��.��F���R�:���C��Ȉ>5b?�L?�Cb>����D�� ���Ľ�N5�'�ۼɕ9���B��N׽*-5>i�;>�7>�\?��Vо��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji����>�	о_�l�z"p���
�>���#�%�a?6����>ƒ?Ƙ+�܌�����<��>ٮ�?���?Qt�>�md?Qj4�~�j����)�?�5?�\�>���;"}�R�ýA�>���(�<2(�0�'?{�@��@�m?��Xҿ���/���O����=g:*>�6>������=}n)=��/��z����=i��>+�)>�>�>��>>5>�{F>0����'�=����u��|:�W�����M���q���m��\���������ļ�K����ma��Ľ�ѻI	>�r�?zg8?�q?Iژ>�y����c>��$�F�g<�������=q��>�j;?pUY? ?I-�=7�پ\j���Q��}߾�/��gm�>�Z?>�r�>П�>�*�=��)>�R�>�s�����>0=�>��+��Uu=�=�;�=���>�?GҰ> _<>=�>1Ѵ�1����h�6�v��˽� �?�n��@�J�I2��&��M�����=�g.?�h>���/=п��P/H?Z���&��+���>#�0?JjW?՚>j���`8U�>[����j�,�> �^l�g�)��%Q>�_?%�h>Q�w>ܙ3�7�7�j�P��s����>�4?1E��Ҝ5��<u��TH��iپe�M>ͽ�>�e&���XJ���x�ߍk�zR{=�;??ͼ��@����9y�����Q>:�Y>F�='�=[�L>�\��ͽlG�x�"=���=C~a>-�?1B->`�=���>j,��Q�V��>�F>� >��@?D$?I�?�����E����(2�oq�>�p�>��>���=C!L�V/�=��>{lo>ZV+��[l�3����C���Q>�`�(�[���h���a=HՕ��8�=%��=���#K=���E=�V�?Sѥ��ۊ�M��w޽��J?D?$�==�w&�	q��r����M�?�@D��?�F
�hV�r�?�?�ܚ����=U��>ヶ>�׾3�P�
?A���L�����lF@�"�?�J�?��g�"��4�c�n�>$?V�޾|O�>iP�>Q��Z9��4�u��=Q��>��H?I���p�D�i�:���	?]�?�������)ɿbv����>&�?Д?-8m�[r���H@�J��>���?�"Z?��j>�ھ=�]�6ˋ>�RA?�yR?�-�>���'�'2?��?��?�I>�g�?^�s?���>o�{��S/�&������k{=�F�;UW�>��>�"¾t�F��Փ��<��]j����Pb>K&=���>���6���̊�=9?���a���e�Mз>�,q>I�I>�>ё ?̺�>�ؙ>��=AU��#����<���L?���?����l����<	g�=�>X��?yN2?|�'� �ξ��>H�]?��?Z�Z?�ݔ>�f����׿��ߵ���<��P>�]�>��>�ّ�?�D>�z׾>aE��߉>�3�>�ʖ�alپ�{��q�/��ɜ>_6 ?֜�>gɶ=��*?��?�oJ>x4'>�?m�.ԕ�@�B�!��>�8�>�>J?z.z?.��>���wS/�����;��B�>��ǧ>��q?U�6?�~�>�3��#᭿�U����r j>Z��?kQ?��)��]?8w?�{?^4V?�S>�.پ���6���Fw�>��!?��e�A��M&����~?Q?���>T5��j�սWּ���S��+ ?+)\?eA&?��&,a���¾�7�<�"�]�U���;n�D���>��>I������=Y>�հ=�Om��F6���f<�k�=��>�=_.7�&x��(?��<�l*�YX�>#~k�[C���>�}^>Fx�ޏl?W)��l���Ȝ�8���<���[W�?��?��?"I
���e�:�?|C�?�Y&?���>F�P���ʾ��
�$:�� <����{gf>��=��;�%���m���J��۷���Ӭ=�A����>p��>�?!n ?~O>7�>-4���/'��Z�"����^��v��s8�5�.�o��jР��1#�_A��0¾��{�+?�>�،����>�
?��g>w�{>��>6λ�A�>X:R>x>�t�>�X>~�4>[d>�"<�jн��}?�Ͼ{��<�k�.����?���?\5.?���>��=�m�4�[?؎�?�u�?��=?)DA��5� Z>�E9>�Q�����>
�>#�>�k�<�ľ-#��J��6���}�>�'�� �2�ȇ�lJ�F�?�P)?�b�<�������跾S_���A�?�}?�4���G���j��V@��y^��"�}С���@&�:ts�iׇ�BІ�*d��ш,���=�b/?2�?����#Ⱦ��ξ��U���?��p~>��>�C�>S+�>�n>�����*�n`H���!�x\�
�?q^�?�	�>,"J?��;?��P?3L?Z�>�W�>7�����>��;��>�>��9?�.?��/?'<?��*?4�`>�g��$���moؾ�?<?��?N?�.?h���½[�����Y��{��8���v�=�Z�<��ֽ�(n���X=/{R>X?����8������k>q�7?��>���>r���,���<�<��>۵
?�G�>} �w|r�/b��U�>3��?��ǂ=E�)>���=R����\Һ"R�=������=�'��$�;��V<=M��=ߜt��}�.e�:���;x�<�R�>��?�;x>�r{>�OJ�7^�0a2���w=B4Z=o{b>��=VP�ݎ�Pa���se��{�>.t�?�'�?o����> :m=q�+�����z2�eþ5��=�(?�ǣ>��Q?-ƀ?3�	?�?���>�	���5���m���盾�@?4?k��>���'���m��G�;��~/?kȎ>|�o���-=yF�ş���r>�"7>�����A��'��ts�z��J�+>��.�??Ҫ�.JB�..�����2��� ?��~>�i�>u:�>	���I��F����j=<��>�Z?��>��O?�4{?��[?�NT>��8�$���љ�+�2�Գ!>>@?K��?��?ay?�x�>��>c�)��$�K���w�S��6ς��W=�3Z>�>��>/��>m2�=�"Ƚ���y�>���=r|b>��>��>Y�>��w>?=�<W8?��>�ݾ�'��X�텢��T�KLq?���?���>8oK���+�W%f��?.���$>z��?�?k�^?>����>H/ =վ���Z ?��>�>X>���V��>t6�<�3>W��>��M�B���&�Z:
=�!(?�M?h����g��)>����ͥ�����n���H��L���7�=��������þ�賾�ƾ��IF�7������?G�1>�,�=Ў(=�m�4}=�[;] >�<���D�����=�I�=Z3"�$f�=��<4O�����<"@=��Ⱦ�K?)tH?�-?��B?ɳr>y�>�Hb�>͗��?�c>��4������3��I��`����پ,)վ��d�[Ş���>�D�>�C=>��=&��;.z�=~�=���=9_��;��<���=l��=���=��=�>�3>�0w?�������N9Q����`�:?��>Ao�=�eƾ@?̖>>Q6��{����q�]?2��?�[�?�?��i�ie�>���収���=,����1>k�=�2��a�>�K>wq��F����e0�?	�@ʕ??�狿ܝϿoa/>�7>Ro>��R�ơ1�^�[���b�$/[�1�!?�;���̾�>Gù=|o߾N�ƾ�+=OC7>��h=�K�=j\���=��y�A<;=�k=��>��C>l��=,M�����=��I=���= �O>H)���6�c',��74=�P�=[b>�%>M��>��?�a0?�Xd?�5�>�n��Ͼ @���H�>C�=F�>z�=prB>T��>?�7?U�D?�K?^��>V��=��>$�>��,��m��l�+̧����<���?�Ά?�Ѹ>�Q<D�A����Cg>��.Žkv?6S1?�k?��>�M�(��g}��B<�WܽF�μ=Ƚ�	s�J��`,�=8�0��/)�8��=i:�>~�>�&O>��)>�8�=>6>2��>�D3=�c>�-�a�<���=kk���>>�����>Pg�<�@�=�(���p�}S�;ڴy<�y=���W~��
�=r��>�>�u�>�1�=�v���*>U���� M�w�=���~B��:e�s�~�5�/��=2��E>��Y>߁��ᑿ�[?#�[>AT:>q��?5t?��>(��+Ӿӝ��8d��QN���=	
>�;�(�=�ga�� N��sϾ���>2��>���>N�l>�,�u)?��|x=`<��e5���>1����b����!q��4��響i�C���D?�F��[��=])~?�I?{ُ?b��>9љ�U{ؾ�k0>�o��t=���b�q�������?I�&?���>���D���ξ��].�>9kG���n�j���(D�f>�E�/�>2����n����<�h톿ۨ|�buY��������>��o?"}�?a�<�؄�u) �����X��wv�>�q?ٗx>?A�-?_!����|2���s{��y? �?W��?o8O==S�=�����&�>�3	?ü�?;��?wbs?H�?����>D|�;!>�#�����=%>c�=��=_O?�q
?�
?�_����	�G��,���o]�צ�<�f�=�P�> �>� s>s�=t�f=w�=�[>�H�>M�>M-e>�*�>AF�>ai��Ά���&?-b�=%ƍ>-<2?�w�>>FY=o<����<PJ�P>?��:+������Ǿ<Kɇ���P=8�̼�,�>�ǿ�5�?��S>����	?/Y����0���S>KU>7�޽b��>d�E>�B}>%o�>� �>LF>�p�>="(>M�Ծ��>m!
��!���C�>�Q��fҾ�7{>r{���e$���	�.<��aK��Z��*��|j�%3��=����<O�?�3��{�k�b(�64��1?�M�>��5?�Z��O⁽;�>��>��>�
��Y����(����߾�=�?��?\cc>EE�>��V?ڦ?�$0�4�#�Z���t��@�x*e��w`��捿�́�O�D5Ž`?1�y?�9B?x+�<�z>��?P&��'���g�>t.�K ;���.=�Ȩ><���c��Ҿy�¾!�:uE>Pno?s9�?i�?��W�R���>�?�5T?��?��?���>����|)#?&��%�*?��?���>�m"?�>�){>U��[��<u?0>-�S����%Z�kQ��<�8;D�6=^��;���=R��=�@�ӽ���X���e���<+��<]i�= V�=}\�>S�U?7�>�s=LA?�{����U�u����"+?�O��aZ����쾞9ž�+�͊Ͻ�]�?F��?�v?~]��O��]-#�VZU>z�>�^�=X�=�t�>��ѽ����lD;>��>L�2=L_c>)?^=�	 ��V׾���=��t>��?է�>�Q��z�=�����KH��`�>~��������CJ���2��9�����u��>�.o?�?<�k�����Y[e��M?)jC?�E?�t�?�sX��A�)V�K�y����=vU�>��:���¾���e૿�V���=��=�6��p-��ABa>>B�f[޾C]n�R�I����RL=7��ҐV=	D�"־_����=j�	>����!�(��LǪ��.J?օj=�夾b�T�g<����>XԘ>��>;�-�y�s@��֬�u�=�V�>�u:>n����ﾎsG��;�d>�>aQE?�V_?k�?�!��:s��B�����c���ȼ6�?Lx�>h?�B>i��=Ӝ������d�rG� �>l��>����G�w;���/���$���>g9?j�>��?X�R?>�
? �`?�*?E?'�>L��3���#B&?���?I��=��Խ�T�A	9��"F����>�t)?��B�(��>u?�?��&?��Q?"�?i�>!� �{8@�(��>r\�>_�W��V���`>��J?ً�>�*Y??׃?.�=>��5�zƢ��䩽W�=(>A�2?.4#?Ϡ?ܳ�>�x�>t���R�=Q*�>��b?�,�?]�o?"�=�? J2>;4�>�͖=[��>���>�	?TBO?��s?�J?oY�>@��<oʭ�]���9lq���P���x;��H<��{=�5�"u��<�ݟ�<V��;�׷��y��y���E��n�����;��>./t>����g/>�@ľjƈ�~�A>����ؾ����u9�Q̹=Il�>�?�>��#���=(�>���>���G�(?ç?Z�?yf�;��b��۾(M��>*=B?���=%�l��a��v�w4h=2�m?�y^?��X�R����g?hGU?HL��I���ӾL����ΰ��V?�?�O?���>���?9�|?��?o�t�T�w�ќ��P���Ž:G�=��w>�X���M�C�m>I�S?)<�>��d>�3>E ���z���;�Sz�>|��?B��?�a�?��,>�k��d�̹�l���^?�j�>����w�?���Fvξy쑾��i��]�6���Gc��g���=�J@��F��6L�Xc�=�w?��o?Cy?�YZ?z��ev^���S�S�y�uV�����+ZC�=sA�CE��&l�� �+���>�� r�;[	���eB�yõ?��#?�5�'��>s����F�+�;�;>�j��z��5��=���r=*N:=��y�2:�$T��9� ?,��>`5�>C�:?�[^��^>�q�0��=7������%8>�T�>���>���>�^	�iH2�e�齠���#�u��v½�v>ȇc?naK?v�n?�\�;1�;W����!��A0��[���%C>�>�3�>�V�����'&��f>��r�f��"�����	�.��=٪2?�>f؜>�'�?�*?�H	�g���xEy��@1����<���>�h?���>��>��Ͻ�� ���>��l?���>U!�>g���cZ!�=�{�:�ʽ.%�>�߭>��>q�o>V�,�]%\��j��4���:9�%��=ըh?������`�Q�>�R?L��:��G<Z~�>uw�E�!����+�'���>Zx?���=��;>�ž����{�z)��sP)??P?h����*���~>��!?Q%�>?�>9!�?nӛ>U}þ����~v?��^?�jJ?�rA?�x�>*�=����%Ƚu�&���,=�w�>��Z>�m=�j�=ތ��:\��_��E=���=m�ͼ+���<�鵼�|N<.��<��3>^Hۿ\uK�[�׾v�=3�+�	�œ���6���Ӈ�]n��	���D��R=y��6���'�1�W�Frd�K����l��:�?��?k���o;��
6��X��E���2��>wHs��f���Ŭ��4�!m���HᾹL��x�!���P�k?i�U�e�L�'?�����ǿ񰡿�:ܾ3! ?�A ?7�y?��7�"���8�
� >�C�<r-����뾬����οG�����^?���>��/��n��>Х�>��X>�Hq>����螾�1�<��?5�-?��>ώr�/�ɿa���
ä<���?/�@�|A?��(����>�U=���>O�	?E�?> N1�jH������W�>�;�?d��?��M=��W�A�	��~e?]8<s�F�J޻D�=BH�=Vf=�����J>jS�>Ј�TA��@ܽ��4>�ׅ>�z"�V���^�!m�<(�]>��ս�?��ö́?�C\�yf�Ԓ/��4���X>L�T?R��>0�=�g,?#0H��wϿ>�\��a?<�?���?��(?���AĚ>7�ܾ7|M?��5?�>�%&���t����=����!�����bV�B��=�b�>t�>�+��y��XO�JT���y�=���3<ÿ�0�;�:ҹ<p6�<wh��Gͽ���Y�=�f���)x�nw�/�9;-N�= 	>ц>b�>P�<>sY?GHa?�T?�%	>�z���Z�R_;�@�\�����i��|�f�LǾX�����U��+z2�=� ��*��� =���=�6R�H����� ���b���F�I�.? u$>�ʾ��M� |-<�qʾ���𼄼�٥�-̾J�1��!n�7͟?��A?����P�V����Y������W?M����ꬾ��=������=&�>���=@��!3��}S�ye/?��#?>ʾ����l?>�l���=�O)?�Q�>ȸ�<�$�>\�!?�q ��򶽓3W>%N*>�m�>���>��= A��5��}�#?��W?e[%�����}�>�Ͼ�w}�\{=F��=��G�Ʈp���U>}R��q���缫":�o}=pF^?Rȍ>�(���3�߄��'
�L�>1�?! ?v�>�v?g�@?��<>P�ԾGcY��W�+���^?��?A,>X��`��9���%?�?�?Xg�>`k����xN�y�׾�O4?�hb?��4?�:=ǁ�b��"��V)?��v?�r^�ms�������V�B=�>�[�>���>��9��k�>�>?(#��G�� ���uY4�%Þ?��@���??�;<!�ќ�=�;?P\�>��O��>ƾ7{������Ǔq=�"�>񌧾}ev�����Q,���8?렃?���>)���������=�ٕ��Z�?|�?����YDg<P���l��n��:�<|Ϋ=��E"������7���ƾ��
�����࿼ӥ�>CZ@�U�u*�>D8�[6�TϿ(��\оnSq���?J��>F�Ƚ����?�j��Pu�W�G�'�H�����sh�>��>q���ؑ�4�{�"};����W��>�H
�g�>�T��d��M����,<���>���>��>����a��m��?���<ο����h��X?�b�?Be�?n�?W]9<�u��{����TG?��s?�Z?��(�G�]�>14�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�l�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.��^?S�[��o���,������>r�C�� b��	B�j�0��c�G���<���{�?�3 @澴?�h�H3%��e"?�î>�#��j;}L=W�>��>D�A>x���K�>�;�*�:��>�G�?���?��?B���������=*�{?��>� �?����A�>��3>Q�ʾ��b=�c>��D�<6�=:"*?h�4?#�?��>U�D�WL�G�4��?���#�b�:��>��w?Ya?dY������+g��?@��ҽ�F�T��>�
�
0�=q����^c=�	><rϼ.�ӽ1�	���?Gp�6�ؿj��Vp'��54?R��>�?����t�+���;_?gz�>�6��+���%���B�\��?�G�?:�?��׾S̼!>�>J�>��Խr���6���a�7>�B?��D��\�o���>���?�@�ծ?zi�Z?���UK���'|�^�Q�;�.��=k�5?<d��I�}>{�>"��=�'t�!\��T#t��x�>�?�>�?���>P<m?��j��E���0=���>��g?
�?�(�b��n�?>'	?zH�X�����یg?@q@]�@��^?�꡿K�Կ�V��qv��S���<�>6)P=�� >�d��c�*��=�4>&�<um>�_�>�(4>�'q>QV�>+��>�i�=����$�t���ט���,����|���ڍ����(�K�ɳ�| ľ�#���f ��pO�
6�����Z� ���.�p%�=��Z?�BE?�6m?��> w���B,>�����<.�y�=���>R:?-�K?��?�=S�y_�su��㬾�������>�j>�>A��>���>�#�=C�C>l{�=`q">&�
>}_�<�8��V9=>�/>�,�>M�>Y�>�C<>��>Fϴ��1��j�h��
w�x̽0�?����S�J��1���9��֦���h�=Ib.?|>���?пf����2H?%���z)��+���>|�0?�cW?�>���T�2:>5����j�6`>�+ �}l���)��%Q>wl?��f>Ԕu>a�3��V8���P������{>�6?�B~9�h�u��H��ݾDmM>a�>��9��7�R�����1qi���{=Va:?�?Zj���䰾F�u�����R>�[>��=���=�GM>��b�лƽ�H�<.=��=X�^>m<?N�->��=��>O���Q�#�>��@>��+>��??V%?��ֻ�����x.�w�v>��>���>�^>rK��L�=F�>�c>����ǂ�!R�,/A��uW>s�~�6�`���m�WT|=hw��6d�=���=h��%<<�|�.=(�~?���(䈿���g��6mD?�+?��=0�F<ƃ"�1 ���G��7�?p�@�l�?��	�ܢV�H�?�@�?�
��v��=�|�>^׫>�ξ��L��?��Ž�Ƣ��	�7*#�XS�?��?��/�2ʋ��l��6>�^%?˱Ӿ���>����r0������s����=�>��O?��ξ�S=��Ͻ��?�$?�ؾ������ƿ��v�G�>���?!P�?�g��p���>A���>���?�Sh?_�>�����b��E��>Q�V?@�J?[�>����[��� ?I��?��y?tI>6��?�s?Zn�>�-x�vZ/�F6������ju=4)\;Ja�>�X>�����gF��ד�h��͸j�b����a>��$=C�>e<��4��e4�=<���yF����f�֡�><3q>%�I>]U�>�� ?rb�>饙>�a=�l��\ހ�䶖���N?�p�?�LG������ܼ>�G�=�鏽h�?_ ?_�=��lw�>��D?�Pu?�Q\?YW>\/ �>�������a:۾KoP>Y�u>0��>���>�����U�ȡ���.��Q�>���>��D�(b������b��9>�>�g3?n��>�ؽi�%?�?��>t��>ON����/l��@�>j��>b1V?��[?���>��A��a/�o��2����ZB�i��>}�?c8?�Lp>(���a(��C7)�� �=�}�>yg�?r?)�����G?F̃?g�?�WW?q�7>�	g��C��̽T�>�
"?���4�B��r"��.�ʮ�>l��>a��>�����t�2��W�G6�kj?,�e?�-?wE��'�c�쐻��;�<�&V��6q�[WG<��:��>Z�>��%�=�8>d�=NX�32���o<U�=�Ɍ>���=m�6�F�{��;+?��9$���5W�=��o�ʓB�xj>X�O>�m���>X?��E��z�³���G��x#Y�u��?=�?l�?Bا���g�=�9?�̇?ց?�Q�>�	���4پ�۾S
]���s���Fl*>L8�>�Z�qQ�X8��?������gi���]�،�>�i�>�1?�] ?O>���>�蘾��&�nH�F��э^���!�8�'�.��y�嗠��E#���������{�)��>T���v޲>�x
?#+h>�5{>V��>}�����>u�Q>��>$.�>� W>۠3>�Q>�h%<1�ν�my?HuɾuhX�'$�ׁ�>��?M��?�p?gp?Oy���Ⱦ^�x?��}?��?�T�>Pn��;4�.��>c�>�FT�!�?�����<T�>�侟Ŭ�tɲ�m�"�<�w>�~0�����L�jS��9?E�%?�p�==���9���h���|�;;n�?��?:�*���H�UTe���C�b"O��y�e���S��G���,r��.��Z8���눿d�/�ع=�-?¢�?r��f�� Ծ)Dj�ƴ<�|%=>�/�>콟>(��>�H>�o��m45���Z��� �e�5�K?"�w?<h�>3�I?.�;?GbP?rL?P5�>�a�>N������>�Q�;�^�>d�>�9?.?��/?�?��*?�b>����c���aؾ�&?��?�?�?�?����,�½PV��
?y���x�Sۀ��=�h�<��׽�Qu�YT=��T>�X?җ�~�8������k>�7?��>b��>���-���<��>M�
?iG�>7 ��}r�*c��U�>a��?I�B�=��)>���=����KtҺZ�=����+�=�?��e;��q<M��=���=�>t�Ӏ��5j�:}��;[s�<c��> �?��>q�>�7��=�4��&��;#�>�J�>�m��1o��2���ez���l�
�*>e��?Δ�?�cS>FSA>���=o��v��*������mg>@]�>��>�ml?5o�?�%?e�G?��/>������'�{�,�D<?� ,?ߓ�>����ʾ��̉3�x�?�X?=:a�����3)�y�¾�Խ]�>�Y/��,~�����D�툻������	��?��?�`A���6��v辩���-[��D�C?��>�R�>�>��)���g�J#�;>��>wR?;�>J�O?0,{?>�[?1VT>��8��"��?ә�f<4�`�!>5@?쮁?�?qy?�^�>�>��)�N ྏL���[��
�H����W=g�Y>���>��>X��>Z��=}zȽg߰�j�>��Q�=h^b>ˇ�>���>��>lw>���<+E?>�>�6̾���Qg��Σ�G�U}X?��?�S?X$�<��#�g�X�P�޾_,�>��?���?5�
?+�>�W	�=G��������'�,��>���>|s�><"�=�=��,>S��>s��>�|ѽ���g�E������?B?��=�`����z�+�>â���Ɗ=m�5� ~��k˺Q������;����S���$�� �پ�?ľ�Zɾ�%���$�Ծ��?z4=�8>�=7@�"Ӟ��g>��G>T�A;�����ؽ�)�Q��=Ů��'�*��z=6�ս��#�!��<�٭��p?&-6?;b?�0?J~>�S>Z)J�] 3>'����?˚�>7��=�g�#yn�����s���>��������a��4���O>�\=m�H>_�O>W�==$�9;ac/>���=-0�=n�<�_�����<��3=u��=/��=�D>;�v=ތj?��T��:��T�H�@.����>���=�r0=t���?Z>P����η�Vu�Ƃ�?��?ȷ�?�D�>тZ��>�=�F�u�E@O=7>ۧ�=��)�lj�
�>�*�<Z�d7y�3����=�?�Y	@\8P? Ł�: ڿ�VM>s;>�>k�R��l0�=�T���j��=b��?��:�Ͼ��>���=���f�ľֈr=��C>i�=>6 ���Z�[�=}]q�ݙ+=�v=n��>�tD>'��=�Ȳ�&��=�A=B��=��S>�Ý�q26�/[*��2,=E�=i�_>^'>��>��?�<0?_Ad?NJ�>Pyn��JϾJQ��;#�>�	�='�>��=o�A>c��>�8?9�D?��K?V:�>�̉=���>g�>r�,�A�m�\D�p����H�<ᆈ?-Ά?���>qP<(A�I���X>��-ŽK`?^J1?�X?��>\���࿄���x&��`���w�lR���T��9�Z�=�T0��JӽpO�=99�>�`�>�Y�>><�>6S�>�� >���>
�>>��=|�Ѽ�'����;s�B���s>�ܺ=<Z�=uu���a̽��5�<���RR�R����P���.|�Kl�=��=X��>�,>���>�G�=R
���.>����j�L���=Wz��B�]<d��Y~��/��5�G!C>@X>僽.����?�RZ>��?>#o�?vu?��>�,��]վ�;����e�o'R��߸=9�>`�=�>�;��A`���M��Ҿc��>Zߎ>�>��l>�,�M#?���w=��[b5���>�|�����!)��9q�$@������qi�|aҺ�D?�F��`��=s"~?�I?]�?��>(��چؾ8;0>�H����=g�z*q��h����?'?���>�쾢�D��1��>++�.��>�Y�m�}����P)��8=<�~߾R��> �Ѿ� ������d��p��m,>��'��)��>�6? �?5S�����J
$�������ح>S�,?N��=��?��?���y��E��e��=�g�?���?*��?�1�=���=����;�>J,	?/��?���?��s?o|?�Jz�>Ӂ�;x� >-���'I�=z�>
��=)�=6s?F�
?	�
?�i���	����&��X^�<��<�͡=E��>
m�>��r>$��=�g=�v�=n/\>�ٞ>%�>��d>��>�O�>�k�����n�&?fW�=�č>Q:2?7t�>\Y=kH�����<NQJ�$L?��;+�17��3�ֆ�<����WP=4
ͼ�.�>��ǿ{4�?:�S>��q?8T���0�4�S>nCU>��޽���>�E>j?}>Zk�>��>B>�p�>�%(>�`Ӿ�>��3r!�HC��R�2iѾ��{>������&�^&	�����E�G�!��|��\�i�c����=�r��<j7�?e����k��)��O���?/��>O�5?���⌆���>x��>�"�>n����m��#���B�߾�(�?4��?!r>}�>�BM?�=?vף��5��i[��b��`��B���S�&u����n���&�����b?~<�?ݒP?_���/��>�z�?�SI�������>��1�$;�q�e;%Hg>���O�1l�o����<W+�>�?���?2d�>Ü9�阠�y�@>7#1?�W?5�i?^�)?�+?�I���?�x%>�?j�?�*?.X'??��>!�
>/x>=r8=���f�������=z����n���W=�D`=[�h=�@�=ד3=�s=�h���g|�n������2=۷�<�O�=�Ǒ=��>�LJ?F/�>�R�>_�+?u�ƾ:]�QO��4��>�U��Ծ�ڼ��b4�޸��?��>`�?��?�� ?[�>��@���'�u٘>Ak>�҉=�Pb>�W�><�������8w>*~�=��^>D��=�����
%��C�O�l>��)>:�>6�>'3����b>����sl���>��,��,��.�e�L�>�i<4��������>��;?Qe/?�>1*׾XJ��9b��`?��=?��Y?�*f?���=|uþ?�(��+�X���B8>(>p�t���K?��q�K��r��^�>�fb�g ��ta>�W�]޾�Tn���I����L=�����W=O0��/־c2�r3�=��	>�����!�������<<J?�@l=na���*U�ॺ�3>2��>��>+9�N
v���@�%����З=,��>g;>k��~+�tzG�H;��>�>LQE?�V_?k�?�!���s���B������b��1ȼv�?�x�>�h?,B>��="�������d��G���>}��>���Z�G�Y;���.��1�$�H��>�8?��>�?`�R?B�
?�`?�*?�D?G&�>=��[���B&?0��??�=w�ԽF�T�� 9�iF����>V�)?v�B����>�?��?��&?F�Q?�?O�>� ��C@����>fY�>��W�zb��>�_>��J?���>@=Y?�ԃ?�=>V�5��颾�֩�XV�=�>u�2?�5#?�?ܯ�>�]�>�����=�z�>��f?��?#�j?���=&'?L�$>��>_^�=�ӗ>���>�m?ȎI?9�l?�pM?k��>�õ<V;̽m����@���^�5U=+)�<�+:=D!̼Uܛ��}w��S�<Q�<�;��[��=Y�A����V���:̬�>��t>���i�.>0�ľ㈾"�A>�Y���������=1:���=�C�>N?C֕>]�#� V�=�t�>H��>
���(?��?B�?1$�;�b�&�۾tM�V��>�pB?{\�=rm��W���v�g�h=��m?}q^?&�X��4����o?c�P?���U�K��־.���|��:g?��?0�n�Yf�>ވ?`�z?��?��}����w˞�,QC�0<t=�ٲ=l|/>�����5���>@�c?#�?|×>�wu>��#���x��������>�B�?���?Q�?�#�=[�`��>��-�9��4m?�޽>^Z�V�,?�r0�t=ƾ>����S�g�;*��%ݨ�1$���\��ce��B���-��XA�=�d?�Yz?}�m?+Z?�b���I���B��k�H`H�*Y�m6���V�j&8�`-�H7_��`� ��'G���˻�5��d�B����?�$?��+�pm�>[����SҾ5�L>	����)����=����/I-=�0=�|�(3�������"?��>�ܼ>�;?�]��WB���.�W'/��k��Cg5>#^�>(k�>�}�>KW���z1���ڽ�*����q�Ž�<v>2wc?h�K?�n?�j��!1�u����!�!�/�~f����B>��>�ω>�}W�a��~6&��Y>���r�{���y��R�	���~=�2?P%�>e��>�H�?? w	��j���ox�Zz1�³�<)*�>�i?4�>3��>��Ͻ�� ���>��l?��>�>1���[!���{���ʽ�%�>�߭>��>�o>��,�$\��j��񃎿�9��z�={�h?����e�`���>9R?��:�G<�|�>��v���!�����'���>�{?���=�;>"�ž`$���{�;5��_Q)?�K?������*���~>�"?X2�>�'�>"%�?H��>|þ������?S�^?�cJ?!hA?Cv�>}�=;2��&Ƚ3�&��r,=~��>��Z>��l=q_�=����R\�h�uuD=K��=�sϼw4�� <G�����H<�*�<��3>piۿFK��oپ����2
��舾0����u��Ŗ��i��u ���Sx����L&'�<V�GTc�֣����l����?e8�?�x��#�������������Q��>w�q�8l�����_�������>����_!���O�! i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾u1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@A{A?��(����e�U=��>�	?�?>ы1��C�E����Z�>8�?���?D N=!�W�%�	��ue?s�;cG�b�޻��=�ԥ=Y\=���ғJ>B�>@���.A��iܽݽ4>܅>�"�����^��D�<�s]>D�ս5��1��?_h[�=�e��/�Jj��F>�"S?F��>�	�=��+?�ZH��oϿ��]��`?�;�?���?ju)?A_����>�ܾ]�L?!�6?uߙ>,'��fs�F��=#�ؼ�Z�r:��U�tl�=#��>�>�22��g�5cQ�V�[��g�=�����Ϳ�)��5$���=��=��ǽYݽ(;�'Y=��E���c�'(㽈"L����=��>7:�>R��>��Y>:aQ?<k?|E�>��>���0��A�����4���n�tݮ�8"��֎�����R�[������{�N0Ӿ� =���=7R�j����� �m�b�w�F���.?v$>�ʾ��M�{�-<�pʾI����̈́��ޥ�G-̾>�1�"n�W͟?��A?������V�:��_Y������W?�O�ɻ��ꬾң�=+���ߡ=%�>���=���� 3�h~S��v0?"]?����l_��y>*>�	��=@�+?.�?"Y<)�>?%?+�!'�O�[>/�3>��>���>	&	>y���_۽�?	�T?!��U�����>c����z�*Ta=Z&>�*5��2� �[>T�<K񌾿�V�����N�<da?$��>+�/�;T/�$¨�I6t�m��=��}?�4�>%�>�:f?I�??T�>2,�"?d�%�,���
��CV?t��?�b2>S�����o�Ҿ��<?:�{?�>�q�����nO���Ѿq�J?��f?��>?��=i��跏����xH7?0�v?�p^�Or��V����V��8�>�X�>Z��>��9��k�>��>?	#��G������0X4�XÞ?��@2��?j�;<�	���=8?W�>#�O��<ƾ����������q=��>�����dv�0���H,���8?��?���>s���^��z��=�ٕ��Z�?}�?~����Cg<Q���l��n����<eΫ=F��E"�����7���ƾ��
� ���5ῼ֥�>BZ@�U�y*�>D8�\6�TϿ#���[оoSq���??��>5�Ƚ����@�j��Pu�R�G�#�H�����$��>�D>������{���;��%�����>]�!�%�>��S��t���ޠ�c��;=��>E{�>嶊>z���ᕽ�ɥ�?�5���`ο����w^�P@X?9n�?"�?�a?D��;��v�~y|��(����G?fau?��[?<���^b�I�:�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�ٶ_?N�a���p���-�uPƽ.��>/ 1��L\����ɿ��Ve���ty�r�?b�?��?�i�T	#��,%?c�>-���;Ǿ$*�<��>:�>��M>��_���u>�	���:�hm	>���?�x�?�m??�������y>�}?��>�ˋ?
�:5�>	>}ҵ����=�N����=�l�Ւ?2�@?y��>)+;>�m8�Ɗ�q�8�	Hg���'�I}8��>��?�"j?(��=nR���lŽ97�-��&CL���<�&"��_v=r1��8x[=Ȗ#>�=>;��������?Lp�9�ؿ j��"p'��54?1��>�?����t�����;_?Qz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>:�>�I�>8�Խ����Z�����7>0�B?T��D��s�o�{�>���?
�@�ծ?ki�J{?Z����x�iq��8� em�96�=?\8?�
��_�>��>"7�;��n�|6��aHq�Lg�>ų?8�?)4�>vUo?U��qN��H�xξ>e_?.��>%A;�m����>��?���)~���p���1q?�1@1	@�R?�Ϝ�y�ؿ�e��p����ᘾQt=����T�=f���gV<�<}�E=8��<��>�&~>G>��>��\>��/>ט�=�+��E������k��w�?��0�G��x�����)�i�V���?��T���԰�/����g��2�l浽�O̼�1>%sP?ϗ5?%�d?��>��%;�E>d�T��~�=��i�hun>�b�>�[S?��\?c�>T ���ξ�=^��3��_h���������>c'�>���>O��>�6>���=��.>(��=�{>�R�>(�R=�7��m_=L��=f�H>���>T�>�C<>��>Eϴ��1��e�h��
w��̽/�?����S�J��1���9��ۦ���h�=Mb.?"|>���?пe����2H?"���w)��+���>z�0?�cW?�>%��L�T�3:>8����j�2`>�+ �yl���)��%Q>ul?�cg>אv>��3��R8��DP��Ȱ��{>զ5?����C29�[bu��H�/ݾ��M>�*�>�w1�������+��ki��{w=|�:?��?�������9u�PԞ�>R>��[>��=�d�=��M>\]b�Ҿɽ�G�d-=f�=�^>�V?�,>��=Iߣ>`���NP�҆�>(B>�',>�@?1'%?�X�}����q����-�.w>$E�>G�>�>�]J�3��=i��> b>U��ע�����h�?��W>c~�nn_�p�t�z y=i�����="�=s� �V�<�X[&=/�~?���2䈿�뾑i��CmD?�+?��=��F< �"�8 ���G��.�?o�@�l�?��	��V�0�?�@�?f��ڵ�=�|�>1׫>ξs�L��?B�Ž^Ƣ��	�m+#�,S�?|�?��/�-ʋ��l�7>�^%?H�Ӿ4X�>p���AD���W����t�>=���>BK?ݯ꾢t��#�5?�+?w��Bn��Evʿ��v�I�>�?���?�h��̙��C�m6�>�a�?/�_?S�>��ھ Z��l�>��Q? hP?)��>���K|C���?ح?�?�I>���?T�s?ɕ�>��y�4q/�v1��r���B�=��`;3�>�>x����qF�(ד�]����j�!���a>�$=��>]e����0�=+�&��F6h�h·>�gq>�$J>�F�>�� ?���>'��>��=W@���Ԁ�kf����J?o��?3�F�:����>�a!=ԇ/����>��?	$�<�݁���>D?��x?�^M?c�g>������������(ξi�>8l�>MK?Uk�>�y�pX�=�V�w��� �>5��>����j-�󧃾(���4��>\u'?��>N�ý�(?��!?�@>���>':b��U����&��-�>�A�>o3>?N�a?�%�>]����v<����i0��X�L�X��>h�?P /?��_>̗��HЯ���:�5����=�v�?f�J?F�����)?�?�}?s�L?���=9�^�������>��"?�� �ssA�'�&��.ڽ��>�k�>Q3�>���n��.�1!!�����?��f?�p-?����3f�v#þn��<l�V�'���I	�<.}��@�>ș>��䱲=��>
��=v�c�s=�nU�<��=lR�>���=�v>�93���H$?Zn>=\�M�=�(q��I>��>ڨj>����K?�����,s�=���+����@�G,�?g�?V��?Ĥ��uj���2?|�?��?��>R���о��Ҿ{���[�Q�#���c>���>��%�9q�|���ӵ��"S���K�X�.�>��>�'?oZ ?�O>��>�0���'��\���[�^�u|�q8���.���`�����"��'��3¾��{��<�>8��, �>��
?h>�;{>`9�>��Ļ\�>%	R>8{>,��>p�W>�4>��>xQ<��Ͻ�p?���t�!��L;���?۟�?�ON?|�>�3���� �g�[?��x?Ӌ�?�U|>�`�ǲD�%�>�&�>����g?��j�!���w>�߾Y(��i���2�����>=��lV�g�X�~�Q�b�?�S-?B�n=}�-m��6	���G5=S��?�&?Xz(���O�$<m�ZkQ�DS��kּo�q�h����I!�	q�s1���L��逄�q�&�w5=+�,?���?W��'D澯���ŉn�u�=��o>��>�,�>��>�<>α��'1�OB]�+�"��gk�}�>I�y?]��>��I?��;?YnP?&L?'��>pm�>�D���Z�>(��;�k�>�+�>�9?d.?c�/?�4?v+?o�a>�L��b���V�ؾ-/?I�?b?�?�R?�����_½����g��mx�Ȁ���=���<��׽��v���W=��T>�X?�����8������k>z�7?��>6��>>��'-��m
�<q�>�
?G�>G ��}r��b��V�>���?[����=��)>��=f���śҺ�Y�=F�����=7���z;��i<���=���=�Tt��*��J#�:ͣ�;�m�<}��>�$?���>M�>P;���,��r�|���}Q>��>�Q��Mq߾�t��TI�j���=}��?�.�?}�>��C>���=�Sݾz���@�Aq�s>1�u>�')?d�X?Bܐ?¯?�/6?�aZ>Τ	��S��g�b��8H�%WG?
,?��>���n�ʾjᨿ9�3�O�?03?`.a�&��x!)�w¾�YԽ��>�Q/�}~������(D�[������(��<��?�ȝ?IjB�|�6�x{辇Ø�#1���xC?#�>�O�>�-�>��)���g�>�C ;>e��>��Q?�"�>��O?O�z?"�[?)T>=�7�-������i)��] >M0@?I��?
�?+y?oG�>��>�H+��g������"���~%��9?Z=mZ>K(�>yS�>8��>Hf�=ȻȽa1��ħ<����=��a>�w�>���>g>�>Ȼw>���<+JH?�!�>?ľ��
�(ق��Ŝ�,���!�i?�߃?��?�V���#���T���5��>[��?�>�?�?o^[�?��=ݕ�lܞ�^-8���>2V�>�`�>���=�$�:�>>h��>z��>W�"�b���%?��N�� ?��F?6�=&��Ŧ|� ��='f��)�=���uw�xl�Ǚ��CB>|ݽ�u������.�������ɾ<�} ��*.��f�?�{>p��=�+>�+�f�:��A=�P5>AoT=��U=�E��)� ��..=ņ0�J��>��g���A�<HȈ��Ǿ0�t?��A?�0?��C?��l>��>�ir�iR�>غ��z�?q r>�ૼ�ɧ���7�Er���d��#̾jپ�h�l✾.j>!�B���>�$>���=��L=$�>U��=�9�=մ2�T۱<��=[��=3��=O�>�>�+>_Gj?Z�?�a��MS�ϥ�=L�>���<@�X><��h?a��=\E��L@���j��ڗ?V��?�?7X�>FAw�෨>y���\�g�ݾ��p>�>�v2��ss��?�u;խ��킿�?R�k�?w�@�b:?4聿d���e�=l.A>)�
>RQR�3�1�A��s��@v�?�?�0:��ZҾU{>
Մ=���ľg�=i�S>5�=�`3��vZ��=:����w1=��==�>��>>�n�=C�����=O@=�t�=W�O>QSK��-�o�-��q0=�+�=��V> [$>l��>c�?Va0?;Xd?�6�>=n��Ͼ$?���H�>��=vE�>�݅=�oB>���>��7?ҵD?��K?F��>u��=
	�>u�>�,���m��m�-̧����<{��?UΆ?�Ҹ>�Q<�A�͠��g>��1Ž�v?�R1?�k?��>��	��-����O�[������<v1��Z���V�>��<K�½2��=z�	>���>��}>� +>��>
�>@I�>b�*��>�."����<���=������U>�ww���H>���<�o=:�<@�.�_1=���3�e=ݹ3=���;���=Q��>EG>���>�v�=�	���6/>ʴ����L�_��=�R���+B�.6d�L~�D/�fM6��B>AEX>����3���?��Y>�r?>���?�;u?��>�$��վ�O��%Me�XLS�ܸ=Ԭ>c=��~;�>X`�U�M��uҾq��>rߎ>��>!�l>�,�B#?��w=��Pb5�n�>�|��l��1)��9q�@������qi�ŐҺݠD?�F�� ��=o"~?��I?b�?���>����ؾ�:0>�H����=r�V*q�8i����?'?��>�쾦�D�2罾0�� � ?��aR��	F(�~o�=�A����>�ȹ�=�
�� �����kz����?��~k���>K/?T��?�<��t�k�/�{��q�o���>\xN?	��=�s�>:x?��-��T �LE���X�<�?�,�?o=�?Z�2>���=�P���>Zc	?���?��?�`s?�e?����>[�;P!>*�����=��>Ry�=���=b?ͯ
?��
?�	���	�kn𾨛���]�Ԟ�<���=�:�>qN�>��q>��=��g=`*�=M�[>s��>ď>zd>D�>@$�>�/��OH�ѿ&?DX�=U��>l2?ј�>�/U=������<AH�(?���*��
���ὢY�<zK���nM=WlԼ�>h�ǿ0F�?O�T>��x�?�s��j�3�P,T>K�T>Q޽u��>��E>�E}>��>���>V�>���>�[(>�FӾHv>0��c!��+C�T�R�T�Ѿ&z>R���K�%�ʠ����(?I�r���f��j�d.���:=�.��<SH�?(���$�k���)�����Վ?=Z�>)6?�،����ϵ>}��>�̍>�I��l����ƍ��bᾂ�?|��?qp>~��>�TQ?٪?��6�4����U���S���W�eM�BT��@��\�����T���E�g?�+�?tP?��;4�>Y�?9�;��g��I7�>c���0?�0�=�]�>#�˾��X��ھ2�� �v�W��>\f�?�f�?�W�>~Y�ئ��2>��>�-o?��h?��?�P?���K?_U��./B?��?ɑ?�y?9(Q>�)>Fɽ�t�=&�(�M3�8�t�����d @����=9�=�}�W;4=�3�=�=�<,To=������׽����ȼ�k�=us�=��>{
>���>�Q?�.�>U)>�[H?ƪ��!`]�6����� ?$
нZ6��N���F���Ծc*�>���?�=�?��>��>3.�m�8��N'>�ǯ>��}<�J>i�>ʈ���n�V�=�
�=*Q(>��`�6i"��=��6������F�;=��>Y�?���>�׋��8>^[������\C�=I�!�������?���Q�(�A������>��W?t�C?�@@>I���ҿ_��?�tS?�?G?�:4?�*>n"��I�4�8���,��*>�s4>��վ�6��Sr���VK�L���-��>����թ�R�E>�j���ھ;�o��NF�!��a=/��B=�����׾}����=j�>�t���!�՗��w���2Q?�C�<F����1R������H#>�	�>��>�D{�s����@�&>��� �=.�>uR9>-Ժ�e���H��| ��8x></0?�w?���?��'��C����/�B᡾���~=�W5?�1�>1�?˄>�5�=�D�����a%c��p�d'�>��>N����;�ᦾ���:J�/
�>ێY>�{u>�I?*|?�<?yv1?k�[?Zk?�5*>��v�}��UO$?#�?���=V���R��[jG��UK�
-�>o?1��ˎ�>2?��$?��&?ϼS?l?'�=	��C[I�2'�>�9�>= Q�欿+��>��V?�>'�K?�(�?�r.>��<��딾�ऽ���=�<>��2?��?$?���>�?�
��[�:	al=�R?�a??s?�/�>��?��>�"?2��>���>�&?Fw$?zMH?�c?�9&?).M>����D��;�^�b����X�y :.N=n~=��.���#.��9u=��]= L���I�=�ᱽ` �ά�=	�缻x�>r7s>[Ε�E�0>��ľP�����@>5���ǘ�������`:�#Ҹ=d�>��?j#�>5�"����=UN�>՜�>��(?��?� ?A1`;)�b��ھnNL���>w�A?�-�=�l��]��w�u��:h=C�m?r3^?X��#��V�b?�]?P`��=���þ��b���龙�O?^�
?z�G���>s�~?��q?���>e�e�#7n�B��TDb�}�j�Bö=�r�>;W���d�yG�>E�7?�K�>-�b>TF�=lt۾�w��m���?��?
�?q��?T(*>��n��1�։
�yq�����>!�>�����>t�$>�+Ѿ�X����վ*�%w���<+�4�˾��������־%�=ӿ<?Na?J*}?AHh?1�_���Z�2�;��U��?i����y��j�a��X[�b�X�E�����9�e�Ҿ0l!��b.>En~�T�@��W�?��(?X3�{[�>R�6���;YA>C.���[����=rz��Qw>=��V=��g�I1�3��;�?k�>���>�U<?F�[�!�>���1���6�Ԣ��
84>ba�>�>���>�e;0�(�= �iHɾ{����Qٽ�2B>g[?"�N?��w?c$��!M<�O�_�!��ȿq�gl��!�S>_$�=�_>b_���QR�]���,��u�$���ݡ���K�=KL;?��y>>���?�
?����{���2�w����>��?�Hs?���>���>������|<�>+�?h�c>����V�jξ Ǌ�Ғ�qTr>M��>�w�>�B�׎d�olH�A֕�O����
E����>���?����T���⢜>rI?�#���L=�+�>RG�x��`1�O���P�>A��>h�$�c�>n����I5�ۇ�j˾r�-?�I�>����`�&��8>/9%?��?���>�P{?s0�>.<_�w	>&W?>�W?�I?3-??�Q?�ۡ=���>�
��ƺ���g=��Q>#�>t��=�բ=ǚ'�G��O��)����N;Մ�<7L����S�q���m<�ީ; J�=`q��NO��_ �7R �
�׾��7�F��<����?��%𾾃����ٶ��X	���˽xG�L����P���[���?��?\����d�?j����g����>�*�K� ��_�鼽[���3Ծ~�����Z���{��a�%�'? ���˽ǿ鰡��:ܾ!! ?LA ?W�y?��_�"���8�Ь >^5�<�5��Z�뾹�����οu���:�^?[��>�
�0��I��>쥂>A�X>�Gq>|���螾�B�<��?Æ-?���>��r���ɿX����Ȥ<���?"�@�wA?��(����?�U=K��>[�	?�@>91�2��۰�b[�>�5�?L��?0JN=�W����w�e?R<��F�3�:2�=�*�=`b=x���J>gj�>�s��MA�V0ܽ*�4>څ>��"�`��U�^�؜�<-�]>PzսAꔽ5Մ?,{\��f���/��T��U>��T? +�>W:�=��,?X7H�`}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�ޅ�=|6�剤�z���&V�x��=[��>a�>��,������O��I��Q��=������2e�m�%4=�Y����;*�|����ɉν�����l���9@�-�==��A>�$�>�X>hW>�T^?��X?P��><�>�4ҽC��b�;���E]B�B[ǽ���_p�����`ʾ����=�wv!�����¾ jS�p>�1xk�)H��bt$��?Z�S�7�Nx?L�+>�����R�����о7�(9��Hm���߾�C<�v.g���?��?�炿�D�&��sF=⟍�_D1?α3�����ZȾ�o�=< 7<�S�Z��>%� >[vɾ��D��G��0??V#�������a(>�ғ�U�L=�F+?M	?�����>W%?H��2����̈́>�\P>*�>�N�> �=����걽��?��M?ӫǽ�á��Ȅ>�|Ǿ��d�P9�=H�=Qgk�w?�1�J>I9�<�|��h8������\ߪ;�#W?��>5�)�L��Q�����/�<=��x?U�?�@�>�lk?��B?V �<N[��F�S��+��Fw=�W?3i?۰>Á��оJ~��߷5?��e?��N>Ih���龓�.��L��?\�n?�V?Xz��ds}��������e6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�֖�s�?�@�?� ��a�D<���8�k�' ��n�<�`�=o%���,�_3�yA8�.�ƾ��
��s���۾�t��>�n@8����>�z7�����~ϿBV��Qaо��r��?p��>E�ɽ?���k��v��G��H�j⋾�&�>�>�����ۑ�F�{��y;�c �����>��h�>�S�e���R��� 8<��>Ƕ�>#��>xM��!��{��?<p��O#ο����4R���X?o^�?�T�?my?�	4<C�w�`�{�cp�G?�ps?�Z?�k$�(e]��i5��xj?Ш�UV`��5���D���V>o2?u�>��-�}�x=E2>��>�5>V/�̋Ŀq	�����\��?ރ�?b����>�p�?[�+?\����AѨ�nO*���˺�??"3> ���)�!�L�=�����z?�{/?��
�F��]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�6�>�]�?+��=�v�>���=}����w���&>�3>X�5�6�?�SL?$��>Q/�=n+�.�+��E�ISQ��m	�`�D�ᖆ>�`?�L?��m>�gɽV�3��!��vʽ@+�����I���8����jH5>�n>>�S>��G��Ѿe�?hm��ؿ�j���k'�A54?��>d�?��C�t�_.��8_?�v�>�5�	,��w&��C��?�G�?a�?J�׾ h̼�	>��>�J�>��Խ�����+�7>R�B?�!�AC����o���>g��?T�@Gծ?�i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*�oֿ����B��r������=��=��2>`�ٽ�d�=٧7=�$9��#���P�=<�>#�d>�	q>d-O>�f;>��)>\���!��u��1�����C�2���C[�а��'v��v��:�����1��-`ý􅤽41Q��<&��x`��L>~??��Z?��]?�Z�>j��	==]�Ǿ�ծ=)����=�>��E?v�<?��>?��$>�a��	�b��:���_�<ΐ����>��`>SJ4?�?�E�>X��K%�>*�#>�U�=��=�t�p��<˽��E`>9�>�v�>���>]<>V>�Ѵ��,����h��v��̽���?l|��*�J�42��"@��4����K�=�\.?3�>���"?пj󭿟@H?��� ��+���>��0?�dW?��>"���AU�� >���.�j�D>m+ ��Vl��)�� Q>�l?2�f>��t>�{3�!K8��P�*!��GV|>�16?%���?9�(�u��H��ܾ�BM>���>N�>��T�ꖿ�
���i���{=�g:?��?Fձ�N��H�u��s��:NR>=J\>�y=t۩=�.M>l�d��rƽ��G�A�,=x��=	-^>k?�@>���=T|�>���J���$�>/�\>&&P>�8?� ?0�ٺ-O��[��x��1�>�>�r>Զ�=s*f��p�=pL�>;+m>�P���¡�
-��mM�<�P>AR%��\}��|���^�=.Ľk$�=E�s=���N��zb<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�a�>�D��W��%����u�F�#=��> H?=f���
P��B>�od
?��?a������ȿPwv����>�	�?��?Q�m��=��q@���>w��?\Y?x�i>re۾��Y�`��>��@?2R?�3�>�1���'��?`߶?
��?�8>�T�?t�+? _�=�(�;����Ѻ��ǟ�G%�`�<͢e�Eh�k�
�[�0����6����T��|L�#�?R�<#��>T=@�Ҩ���*>��T������=���>)0?ܛ>�ؐ=[u?��
?V'�>����KK<u���]�A���K?Ʃ�?����
n�B޾<F��=�_�0?r,4?��V�׉Ͼ��>��\?���?�[?'w�>,���8��V濿�����r�<H�K>a+�>r��>LD��<^K>�
վ2cC��N�>/^�>�����Aھ������D�>�Y!?�e�>�ϯ=� ?ѥ#?�_j>��>RE��/���E�oj�>\n�>�??�~?�?�����T3����J롿�[���N>�y?�K?�ݕ>����ო�F�B��I��	��l��?�dg?�/�"?� �?��??%�A?�2f>��&�׾������>~�!?>u�G�A��%���
��?J?*�>p��"��%��`��(���'z?�(\?:�&?���	_�J�¾�Q�<�T
����];�L���>K�>f���JV�=jo>�ػ={Kp�`�5��&�<���=4�>��=��5��L��0=,?¿G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Y�>���>(�l���K���ڙ���F��_�ŽK[�� ?>�>?i��>�F>�-�>5̢��'��������Y`����6�%2�x�"���ǭ�7[!�����~�v�C�>|؃����>�$?_f>�]�>
��> E�<�:�>@F>��>���>n=e>�Y.>o>mHW<�ٽLFR?������'�Ю�zȰ�i@B?C[d?4R�>�Rf�Nv�������?���?k�?��v>Ah��+�vS?���>EJ���g
?��:=p*
���<WS��=���ч�V���>��ؽ�):���L���f��]
?.?&����̾ؽ۔����=qM?t:&?����QB�!�r����ci_�C^��7���X��1M� ���w��������Յ�E���E>��?#��?�5Ѿm�7������#���y��4���>A,]><�p> �>������i�V� YR�_;y���1?���?�υ>��7?$[Q?��G?(-e?�>t�p>#�_�	�	?�.b=.�>U�?��D?t1)?Ut5?�"?�?L��=��"��*
�޼񾑶�>��
?&21?��?��?�ܽ"�=Z����Fl��H��/!�$�w=�$½z���J<=��>8��>Ѿ?;~H�wOA��p�\�>n�6?p�>K"�>93��.o+�c��>-��>��>.���������?���?�.*���=��>,2�=����p�<f��=���:��=h�z����`�wH>�_P=I���������z���%;�H�>�?&�>�}�>f���� �C��!��=��W>��R>S�>ĳپV���3��h�%�w>cN�?!��?�n=���=���=�������޳����q�<��?!#?٤T?���?&_=?=u#?��>����J��x5��7f���?e!,?=��>�����ʾ��ǉ3���?=[?�<a�1���;)��¾�Խ;�>�[/�d/~����(D�>������)��??A�8�6��x������[��U�C?�!�>/Y�>`�>D�)�S�g�9%��1;>���>8R?YG�>��O?L�{?iZ?�C>�9<��%��������n�'>�XA?V��?�b�?�\x?Q��>�>ô*�
⾈p��*f3�D}�T����,>=A�g>��>���>���>���=��ɽ�ý�9�:�=�e>�a�>+ǧ>Y��>uxq>�V�<�D?�n�>�¾R�䕾<�t�[.���r?-�?�-?8b=����<�R�DC�>���?g��?ȡ"?��V����=��j��9���:��-~�>槺>��>�[�=�=/�>��>q��>M/��d��=A���W��W?b�C?�H�=��ȿalr�Nt����V,<'H���GZ������Z�Ƹ�=:q������s���4`�K➾������
1���.y�/�?��k=� >oP�=�8�<�(��Ys�<[�3=:=U<��<8�|�# ��a����:O˕�35�X^1<�9=�1i��l˾&|}?�6I?��+?8�C?�y>�:>m$3����>�d�� 4?�V>�O�h���,6;�ؒ��S$��R�ؾ	�׾�0d��ğ�0E>8�H�~>��2>Z7�=�v�<���=
�s=�Ў=b�a�%�=��=�\�=���=���=?�>�L>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��8>/�>��R��71�P[�=�`��Y��!?	�:�U�̾�g�>E �=�޾ƾ�4=��7>�b=���;\��)�=�x�QP>=�7g=ix�>�tC>�y�=���Eݶ=��H=��=T�N>�љ�W�4���,�E�1=�&�=�wb>=&>�'�>��?TU.?��b?n��>��k�7wʾ�m��7x�>���=z`�>�=�=l�H>���>�Z9?�fE?��K?�٭>��x=��>|��>��-���m���⾻a���=���?2�??��>ȿ�<��<��w ���:�1�ؽ�R?�V4?
�?�2�>�*�t�ݿ�,!�)�������1��ep=�S�VJw�m���ϱ�aa۽($�=6՜>;��>c��>T�~>͡6>�)M>���>m!	>k�<=EK�=��Y:�f�<�I���^=Aޥ���<�-ټ��z�	�� ���2"����F���ٍ<5qT<���=m��>I?>���>V��=	���=/>Ӹ���L�ſ=yF��<+B��2d�H~��/��U6�޴B>X8X>����14��'�?:�Y>�l?>-��?�Bu?��>�!�R�վZQ���He��TS�Gȸ=ʵ>6�<��y;��Y`���M�CyҾꝩ>�l�>��l>��=]�SV�U��e��i=��A>w���=9�҄�����֤����q��q����1?���%�E(�?M͆?�M?���=m�a>�#�'>�>�g{�4�[>jl���!|���
?��`?\�?��1���~�ƾ�o|�Xl�>��d��J��b��&8��k��s�þVk�>>���Fܾ�:��م�:y���I�͡{����>��Y?Uũ?ث;��~���U����4Wc�b��>ĵc?�ԓ>�
?T1?B�����C��t�=�{_?[��?�<�?%P%>���=��콯��>��?ET�?҆�?�wc?�I���+?�<�2>�:!��>TJ>��>�%?>�o?���>���>����c���!
�3�/�l��e�=�/>GH�>�
M>�F>ԩ=��=�8{��4>��y>H��>ڤp>���>��>kS���7��#?3p�=P�>[�1?}e�>%�F=ѕ��Z��<��c��lA��$,�t��y�߽��<�&����*=����1�>��ǿz��?O�R>�>���?`��a�4�/4K> �M>:M��Y�>�D@> w>}B�>=}�>[>��>k"*>aӾ�%>��� N!���B��5R�$�Ҿu$w>�	����(�W	�����7HK��Y��J���/j��.����<����<��?TH����k��j*�s����?�W�>~5?�Ō��셽*�>�w�>]t�>����o���ˍ�����9�?1��?c>�[�>łW?LG?�w1�ڮ2�֡Z���u��:A�/e�
�`�����t�����
���½�F_?ؠx?��A?�8�<` z>ئ�?0�%��t���8�>2�.��;�r�<=.Ӧ>w��=M`�
�Ӿ�pþ��NF>�(o?5 �?��?t"U�5�:�+>NhN?o�+?��?o�?��?�X>-L?-B8>^??,?�<?�1?~?56i>�F>��==&�
=�(�����]sZ��*��>D�������=���=F٩=)��z�M=�m� �a�#=lЏ�Ծ[=PS��X��=?�>2��>�]?���>R��>��7?�/�Yg8�~鮾@�.?�v>=����W��_Ȣ�م�>�wj?m�?��Z?vwe>n�A���B��>��>�%>t\>_\�>�����D�]��=��>�'>7>�=t�L�.ہ�X�	�hj���
�<�>R��>��{>⚊� �'><��5�x�j7c>�:P�O�����R��>G��0�M s��.�>�&L?��?���=E���>���jf��(?/<?|FM?G4�?X��=�۾��9�(�I�y���R�>�*�<	��Ar��?����J:�@�l:�r>�q���թ�R�E>�j���ھ;�o��NF�!��a=/��B=�����׾}����=j�>�t���!�՗��w���2Q?�C�<F����1R������H#>�	�>��>�D{�s����@�&>��� �=.�>uR9>-Ժ�e���H��| ��8x></0?�w?���?��'��C����/�B᡾���~=�W5?�1�>1�?˄>�5�=�D�����a%c��p�d'�>��>N����;�ᦾ���:J�/
�>ێY>�{u>�I?*|?�<?yv1?k�[?Zk?�5*>��v�}��UO$?#�?���=V���R��[jG��UK�
-�>o?1��ˎ�>2?��$?��&?ϼS?l?'�=	��C[I�2'�>�9�>= Q�欿+��>��V?�>'�K?�(�?�r.>��<��딾�ऽ���=�<>��2?��?$?���>�?�
��[�:	al=�R?�a??s?�/�>��?��>�"?2��>���>�&?Fw$?zMH?�c?�9&?).M>����D��;�^�b����X�y :.N=n~=��.���#.��9u=��]= L���I�=�ᱽ` �ά�=	�缻x�>r7s>[Ε�E�0>��ľP�����@>5���ǘ�������`:�#Ҹ=d�>��?j#�>5�"����=UN�>՜�>��(?��?� ?A1`;)�b��ھnNL���>w�A?�-�=�l��]��w�u��:h=C�m?r3^?X��#��V�b?�]?P`��=���þ��b���龙�O?^�
?z�G���>s�~?��q?���>e�e�#7n�B��TDb�}�j�Bö=�r�>;W���d�yG�>E�7?�K�>-�b>TF�=lt۾�w��m���?��?
�?q��?T(*>��n��1�։
�yq�����>!�>�����>t�$>�+Ѿ�X����վ*�%w���<+�4�˾��������־%�=ӿ<?Na?J*}?AHh?1�_���Z�2�;��U��?i����y��j�a��X[�b�X�E�����9�e�Ҿ0l!��b.>En~�T�@��W�?��(?X3�{[�>R�6���;YA>C.���[����=rz��Qw>=��V=��g�I1�3��;�?k�>���>�U<?F�[�!�>���1���6�Ԣ��
84>ba�>�>���>�e;0�(�= �iHɾ{����Qٽ�2B>g[?"�N?��w?c$��!M<�O�_�!��ȿq�gl��!�S>_$�=�_>b_���QR�]���,��u�$���ݡ���K�=KL;?��y>>���?�
?����{���2�w����>��?�Hs?���>���>������|<�>+�?h�c>����V�jξ Ǌ�Ғ�qTr>M��>�w�>�B�׎d�olH�A֕�O����
E����>���?����T���⢜>rI?�#���L=�+�>RG�x��`1�O���P�>A��>h�$�c�>n����I5�ۇ�j˾r�-?�I�>����`�&��8>/9%?��?���>�P{?s0�>.<_�w	>&W?>�W?�I?3-??�Q?�ۡ=���>�
��ƺ���g=��Q>#�>t��=�բ=ǚ'�G��O��)����N;Մ�<7L����S�q���m<�ީ; J�=`q��NO��_ �7R �
�׾��7�F��<����?��%𾾃����ٶ��X	���˽xG�L����P���[���?��?\����d�?j����g����>�*�K� ��_�鼽[���3Ծ~�����Z���{��a�%�'? ���˽ǿ鰡��:ܾ!! ?LA ?W�y?��_�"���8�Ь >^5�<�5��Z�뾹�����οu���:�^?[��>�
�0��I��>쥂>A�X>�Gq>|���螾�B�<��?Æ-?���>��r���ɿX����Ȥ<���?"�@�wA?��(����?�U=K��>[�	?�@>91�2��۰�b[�>�5�?L��?0JN=�W����w�e?R<��F�3�:2�=�*�=`b=x���J>gj�>�s��MA�V0ܽ*�4>څ>��"�`��U�^�؜�<-�]>PzսAꔽ5Մ?,{\��f���/��T��U>��T? +�>W:�=��,?X7H�`}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�ޅ�=|6�剤�z���&V�x��=[��>a�>��,������O��I��Q��=������2e�m�%4=�Y����;*�|����ɉν�����l���9@�-�==��A>�$�>�X>hW>�T^?��X?P��><�>�4ҽC��b�;���E]B�B[ǽ���_p�����`ʾ����=�wv!�����¾ jS�p>�1xk�)H��bt$��?Z�S�7�Nx?L�+>�����R�����о7�(9��Hm���߾�C<�v.g���?��?�炿�D�&��sF=⟍�_D1?α3�����ZȾ�o�=< 7<�S�Z��>%� >[vɾ��D��G��0??V#�������a(>�ғ�U�L=�F+?M	?�����>W%?H��2����̈́>�\P>*�>�N�> �=����걽��?��M?ӫǽ�á��Ȅ>�|Ǿ��d�P9�=H�=Qgk�w?�1�J>I9�<�|��h8������\ߪ;�#W?��>5�)�L��Q�����/�<=��x?U�?�@�>�lk?��B?V �<N[��F�S��+��Fw=�W?3i?۰>Á��оJ~��߷5?��e?��N>Ih���龓�.��L��?\�n?�V?Xz��ds}��������e6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�֖�s�?�@�?� ��a�D<���8�k�' ��n�<�`�=o%���,�_3�yA8�.�ƾ��
��s���۾�t��>�n@8����>�z7�����~ϿBV��Qaо��r��?p��>E�ɽ?���k��v��G��H�j⋾�&�>�>�����ۑ�F�{��y;�c �����>��h�>�S�e���R��� 8<��>Ƕ�>#��>xM��!��{��?<p��O#ο����4R���X?o^�?�T�?my?�	4<C�w�`�{�cp�G?�ps?�Z?�k$�(e]��i5��xj?Ш�UV`��5���D���V>o2?u�>��-�}�x=E2>��>�5>V/�̋Ŀq	�����\��?ރ�?b����>�p�?[�+?\����AѨ�nO*���˺�??"3> ���)�!�L�=�����z?�{/?��
�F��]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�6�>�]�?+��=�v�>���=}����w���&>�3>X�5�6�?�SL?$��>Q/�=n+�.�+��E�ISQ��m	�`�D�ᖆ>�`?�L?��m>�gɽV�3��!��vʽ@+�����I���8����jH5>�n>>�S>��G��Ѿe�?hm��ؿ�j���k'�A54?��>d�?��C�t�_.��8_?�v�>�5�	,��w&��C��?�G�?a�?J�׾ h̼�	>��>�J�>��Խ�����+�7>R�B?�!�AC����o���>g��?T�@Gծ?�i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*�oֿ����B��r������=��=��2>`�ٽ�d�=٧7=�$9��#���P�=<�>#�d>�	q>d-O>�f;>��)>\���!��u��1�����C�2���C[�а��'v��v��:�����1��-`ý􅤽41Q��<&��x`��L>~??��Z?��]?�Z�>j��	==]�Ǿ�ծ=)����=�>��E?v�<?��>?��$>�a��	�b��:���_�<ΐ����>��`>SJ4?�?�E�>X��K%�>*�#>�U�=��=�t�p��<˽��E`>9�>�v�>���>]<>V>�Ѵ��,����h��v��̽���?l|��*�J�42��"@��4����K�=�\.?3�>���"?пj󭿟@H?��� ��+���>��0?�dW?��>"���AU�� >���.�j�D>m+ ��Vl��)�� Q>�l?2�f>��t>�{3�!K8��P�*!��GV|>�16?%���?9�(�u��H��ܾ�BM>���>N�>��T�ꖿ�
���i���{=�g:?��?Fձ�N��H�u��s��:NR>=J\>�y=t۩=�.M>l�d��rƽ��G�A�,=x��=	-^>k?�@>���=T|�>���J���$�>/�\>&&P>�8?� ?0�ٺ-O��[��x��1�>�>�r>Զ�=s*f��p�=pL�>;+m>�P���¡�
-��mM�<�P>AR%��\}��|���^�=.Ľk$�=E�s=���N��zb<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�a�>�D��W��%����u�F�#=��> H?=f���
P��B>�od
?��?a������ȿPwv����>�	�?��?Q�m��=��q@���>w��?\Y?x�i>re۾��Y�`��>��@?2R?�3�>�1���'��?`߶?
��?�8>�T�?t�+? _�=�(�;����Ѻ��ǟ�G%�`�<͢e�Eh�k�
�[�0����6����T��|L�#�?R�<#��>T=@�Ҩ���*>��T������=���>)0?ܛ>�ؐ=[u?��
?V'�>����KK<u���]�A���K?Ʃ�?����
n�B޾<F��=�_�0?r,4?��V�׉Ͼ��>��\?���?�[?'w�>,���8��V濿�����r�<H�K>a+�>r��>LD��<^K>�
վ2cC��N�>/^�>�����Aھ������D�>�Y!?�e�>�ϯ=� ?ѥ#?�_j>��>RE��/���E�oj�>\n�>�??�~?�?�����T3����J롿�[���N>�y?�K?�ݕ>����ო�F�B��I��	��l��?�dg?�/�"?� �?��??%�A?�2f>��&�׾������>~�!?>u�G�A��%���
��?J?*�>p��"��%��`��(���'z?�(\?:�&?���	_�J�¾�Q�<�T
����];�L���>K�>f���JV�=jo>�ػ={Kp�`�5��&�<���=4�>��=��5��L��0=,?¿G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Y�>���>(�l���K���ڙ���F��_�ŽK[�� ?>�>?i��>�F>�-�>5̢��'��������Y`����6�%2�x�"���ǭ�7[!�����~�v�C�>|؃����>�$?_f>�]�>
��> E�<�:�>@F>��>���>n=e>�Y.>o>mHW<�ٽLFR?������'�Ю�zȰ�i@B?C[d?4R�>�Rf�Nv�������?���?k�?��v>Ah��+�vS?���>EJ���g
?��:=p*
���<WS��=���ч�V���>��ؽ�):���L���f��]
?.?&����̾ؽ۔����=qM?t:&?����QB�!�r����ci_�C^��7���X��1M� ���w��������Յ�E���E>��?#��?�5Ѿm�7������#���y��4���>A,]><�p> �>������i�V� YR�_;y���1?���?�υ>��7?$[Q?��G?(-e?�>t�p>#�_�	�	?�.b=.�>U�?��D?t1)?Ut5?�"?�?L��=��"��*
�޼񾑶�>��
?&21?��?��?�ܽ"�=Z����Fl��H��/!�$�w=�$½z���J<=��>8��>Ѿ?;~H�wOA��p�\�>n�6?p�>K"�>93��.o+�c��>-��>��>.���������?���?�.*���=��>,2�=����p�<f��=���:��=h�z����`�wH>�_P=I���������z���%;�H�>�?&�>�}�>f���� �C��!��=��W>��R>S�>ĳپV���3��h�%�w>cN�?!��?�n=���=���=�������޳����q�<��?!#?٤T?���?&_=?=u#?��>����J��x5��7f���?e!,?=��>�����ʾ��ǉ3���?=[?�<a�1���;)��¾�Խ;�>�[/�d/~����(D�>������)��??A�8�6��x������[��U�C?�!�>/Y�>`�>D�)�S�g�9%��1;>���>8R?YG�>��O?L�{?iZ?�C>�9<��%��������n�'>�XA?V��?�b�?�\x?Q��>�>ô*�
⾈p��*f3�D}�T����,>=A�g>��>���>���>���=��ɽ�ý�9�:�=�e>�a�>+ǧ>Y��>uxq>�V�<�D?�n�>�¾R�䕾<�t�[.���r?-�?�-?8b=����<�R�DC�>���?g��?ȡ"?��V����=��j��9���:��-~�>槺>��>�[�=�=/�>��>q��>M/��d��=A���W��W?b�C?�H�=��ȿalr�Nt����V,<'H���GZ������Z�Ƹ�=:q������s���4`�K➾������
1���.y�/�?��k=� >oP�=�8�<�(��Ys�<[�3=:=U<��<8�|�# ��a����:O˕�35�X^1<�9=�1i��l˾&|}?�6I?��+?8�C?�y>�:>m$3����>�d�� 4?�V>�O�h���,6;�ؒ��S$��R�ؾ	�׾�0d��ğ�0E>8�H�~>��2>Z7�=�v�<���=
�s=�Ў=b�a�%�=��=�\�=���=���=?�>�L>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��8>/�>��R��71�P[�=�`��Y��!?	�:�U�̾�g�>E �=�޾ƾ�4=��7>�b=���;\��)�=�x�QP>=�7g=ix�>�tC>�y�=���Eݶ=��H=��=T�N>�љ�W�4���,�E�1=�&�=�wb>=&>�'�>��?TU.?��b?n��>��k�7wʾ�m��7x�>���=z`�>�=�=l�H>���>�Z9?�fE?��K?�٭>��x=��>|��>��-���m���⾻a���=���?2�??��>ȿ�<��<��w ���:�1�ؽ�R?�V4?
�?�2�>�*�t�ݿ�,!�)�������1��ep=�S�VJw�m���ϱ�aa۽($�=6՜>;��>c��>T�~>͡6>�)M>���>m!	>k�<=EK�=��Y:�f�<�I���^=Aޥ���<�-ټ��z�	�� ���2"����F���ٍ<5qT<���=m��>I?>���>V��=	���=/>Ӹ���L�ſ=yF��<+B��2d�H~��/��U6�޴B>X8X>����14��'�?:�Y>�l?>-��?�Bu?��>�!�R�վZQ���He��TS�Gȸ=ʵ>6�<��y;��Y`���M�CyҾꝩ>�l�>��l>��=]�SV�U��e��i=��A>w���=9�҄�����֤����q��q����1?���%�E(�?M͆?�M?���=m�a>�#�'>�>�g{�4�[>jl���!|���
?��`?\�?��1���~�ƾ�o|�Xl�>��d��J��b��&8��k��s�þVk�>>���Fܾ�:��م�:y���I�͡{����>��Y?Uũ?ث;��~���U����4Wc�b��>ĵc?�ԓ>�
?T1?B�����C��t�=�{_?[��?�<�?%P%>���=��콯��>��?ET�?҆�?�wc?�I���+?�<�2>�:!��>TJ>��>�%?>�o?���>���>����c���!
�3�/�l��e�=�/>GH�>�
M>�F>ԩ=��=�8{��4>��y>H��>ڤp>���>��>kS���7��#?3p�=P�>[�1?}e�>%�F=ѕ��Z��<��c��lA��$,�t��y�߽��<�&����*=����1�>��ǿz��?O�R>�>���?`��a�4�/4K> �M>:M��Y�>�D@> w>}B�>=}�>[>��>k"*>aӾ�%>��� N!���B��5R�$�Ҿu$w>�	����(�W	�����7HK��Y��J���/j��.����<����<��?TH����k��j*�s����?�W�>~5?�Ō��셽*�>�w�>]t�>����o���ˍ�����9�?1��?c>�[�>łW?LG?�w1�ڮ2�֡Z���u��:A�/e�
�`�����t�����
���½�F_?ؠx?��A?�8�<` z>ئ�?0�%��t���8�>2�.��;�r�<=.Ӧ>w��=M`�
�Ӿ�pþ��NF>�(o?5 �?��?t"U�5�:�+>NhN?o�+?��?o�?��?�X>-L?-B8>^??,?�<?�1?~?56i>�F>��==&�
=�(�����]sZ��*��>D�������=���=F٩=)��z�M=�m� �a�#=lЏ�Ծ[=PS��X��=?�>2��>�]?���>R��>��7?�/�Yg8�~鮾@�.?�v>=����W��_Ȣ�م�>�wj?m�?��Z?vwe>n�A���B��>��>�%>t\>_\�>�����D�]��=��>�'>7>�=t�L�.ہ�X�	�hj���
�<�>R��>��{>⚊� �'><��5�x�j7c>�:P�O�����R��>G��0�M s��.�>�&L?��?���=E���>���jf��(?/<?|FM?G4�?X��=�۾��9�(�I�y���R�>�*�<	��Ar��?����J:�@�l:�r>�q��Kʦ�-+j>���־GQl�NK����ηA=2���CI=���9\ھ.4��_��=F;>���ܣ#�b����Ԫ���G?��G=|.���/@�����)Y>��><��>�rW��n�y�:�m9�����=�V�>��:>�������F�������=	`\?�e�?_�?�ܾل��X<S�ݦ徬�Ⱦ�<4�F?��>o��>I�
>c�=�3��7� ���v���o���>\�?_3����J������]�f�E��hz><g?��!>�M�>q�t?�8$?V?�wY?��?��x>X��������?f(�?2�f>����R4�x�?���R����>�R?�o2�>׷?�W?�1?,�M?�
?�E>���3�G��O�>�SQ>?j�夿]�>%�x?5�>�e?x4�?EU�=��K��ih�����5=aK>�e=?�^?M?���>O�?������Q�h˧>nm$?:�n?y�r?y��>j?���>���>5�]>i!�>	��>��>i�<?j�5?`P?�,�>aAY=>�	�s��g�ݽg��=uf�G
�<��>���<�T+��Q$�0�<A�A>���=�Q>z���}G��ɶ�򨊽���>@ks> ���l0>��ľ8��*MA>Ϧ������p\���:��}�=���>W?���>+�"���=��>z�>v����'?��?/?��:�ub���ھ_L�Z�>�B?���=ixl������"v�`�g=K�m?�^^?�PW�Х��O�b?��]?@h��=���þy�b����h�O??�
?"�G���>��~?i�q?W��>��e�#:n�(���Cb���j�'Ѷ=^r�>GX�R�d�~?�>f�7?�N�>7�b>J%�=ku۾�w��q��c?��?�?���?�**>~�n�T4�=8��R��ڽk?e��>���1�?�,�x��ȿ� �������ľy�ž�k��Io;*\�L����1��o�=R�.>�5:?�|F?�Y?bK�9Q]��W�2�������ي:�Q@���a�D�a��BP��Ɋ���M���c��n)�=񛧾o(�/԰?e�2?~Ti�"!�>wƅ��	�I�߾��%>9����-?���f=Cq��2�����<(V������n�о��?Q/�>h��>G�:?��\��I�*"-���#�4�W�>>���> �>}��>�6 �!��q�m���l�6��0�\>�He?��L?�k?�|޽�c1��������=�_s���/@>&>Zm�>1�T�C��z!�2h=�!�u�9��f��	���/=��6?0��>��>�I�?NE
?���Uz���l�-�&��w`<�v�>KDd?�X�>ߎ>b�ݽ&��e�>�v?(޶>{-+>٭Q�8�](~��_�8��>�T�>H��>ǝ=t�M�"g����yp���X3���y>��y?��w�ulE����>��e?wE{�6}4����>K���N��پQ���2>x�?�=�B>��;E<�ٞ��P,����J?N?�>&�g�d
<��p>.\�>��?a�?��?#��>��@�>Ϝ>\i<?��r?p�|?_^?��>g��=D��j�B�v�H;}\>�v�=���=Eـ�	�4�a��6�j�ِ��P�
>pcC=�Q��E=��=Gq����1=��K=E�>�lۿ=@K�a�پg���^C
��䈾(����g����R[�����Wx����''�V�}5c�릌���l�5��?�;�?Pz��K.��F���7����������>��q�.o�X竾���+.�����X����a!���O�I$i�5�e�P�'?�����ǿ񰡿�:ܾ5! ?�A ?7�y?��5�"���8�� >EC�<0-����뾬����ο@�����^?���>��/��q��>ܥ�>�X>�Hq>����螾�1�<��?7�-?��>ǎr�0�ɿb���o¤<���?0�@�A?-)�7r�$K\=���>��	?�B>�A0��K����j|�>^ �?���?*A=��V����S�d?� <�TF��E��2��=>��=��=e���I>e��>���W�B��ٽ�5>���>�`"�C�_�I��<��\>0�ֽAݐ�6Մ?{\�sf���/��T���T>��T?+�>�:�=��,?G7H�Q}Ͽ��\��*a?�0�?��? �(?&ۿ��ؚ>��ܾ��M?dD6?���>�d&��t����=7�Ί��L���&V����=3��>�>�,�����O� I��[��=V�'�ƿ.�$�	}�K_=�yݺޤ[�c~�`�����T�n#���fo�+�轒�h=��=��Q>ml�>�%W>Q4Z>gW?j�k?�N�>��>�7�U���ξL|��G�����������]��R��߾{�	������g�ɾ�!=�!�=�6R�����|� �Y�b���F���.?�o$>-�ʾ9�M�0�,<{rʾ�����	�*̾X�1��n�N̟?k�A?������V����Pg�os��_�W?�P����|款z��=(k��^�=�#�>i��=���@!3�X}S���3?�?����9��'>6����^=�-?�x?��=�ʩ>�'?L����U�>2vS>?W�>
�>��>Jڦ����Ӊ?c�M?)b���%���_�>֖��\˂����=�8>?6�:��\�[>�4/<t������5p��"Ǡ<X1W?V��>*�C��J���,�B=_{x?��?wĠ>�bk?C?F$�<����=S���
���v=ˋW?�i?&	>sj���Lо�㦾+\5?�Qe?�JO>��h��܇.���Q0?|�n?0?�����|��풿f��x6?:�v?zr^��s��/���V��=�>yZ�>Y��>��9�
k�>C�>?�#��G��ĺ���Y4��?��@���?<<�����=:;?�[�>��O��>ƾ�z��񂵾ƚq=�"�>&����ev�`���O,��8?ɠ�?���>ܓ������~�=����W�?
�?�ê���S<����l�y���J�<x�=l��Z#�/���7���ƾʩ
�����9�ż�>lO@'��!�>�W8�W4�R_Ͽ\����оB�p���?ȅ�>�tɽ������j��$u���G���H�ӓ�>FQ>1������:B{�I�;�����S�>@P���>?�P��������=<T)�>Y@�>˽�>�
��t��ގ�?�.���1ο�o���,���Y?�s�?�v�?��?*<ay�Źy��c�;�F?�Ls?;8Z?Z� �$\�w�-��j?h_��|U`� �4�_HE��U>�"3?�B�>V�-���|=}>J��>�f>�#/�x�Ŀ�ٶ�!���_��?��?�o���>w��?}s+?�i�8��k[����*���+��<A?�2>����,�!�G0=�OҒ���
?&~0?`{�^.�]�_?+�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>c����8Ǿ��<���>�(�>*N>_H_���u>����:�i	>���?�~�?Qj?���� ����U>	�}?\$�>��?o�=�a�>`d�=B�*-��k#>�"�=b�>��?��M?L�>EW�=z�8�~/�:[F��GR�]$�5�C��>y�a?�L?Kb>���q2��!��uͽ�c1��P鼜W@�=�,���߽6(5>��=>�>Q�D��Ӿ��?�9�:G׿1ѝ�O ���3?��>y۶>�� ,��39?��	>����,��䍿�~
=,��?>F�?��?&����j2�=#��>�>?��ʀ+���4�I�x>]�D?PF^���x�8?D���|>��?+�@7�?�5b��h?��j����~��3���5����=k�6?�*�~�x>���>PZ�=u�v�.���t�s�0M�>$n�?>��?���>p]l?o��C�Ud,=>]Ok?�?��C�*��|�D>��?��S����C�d�e?�
@�e@H~^?Kâ�v���h���-*#��q��0S�=\y�=���=��ʽ-"�=���;c�<{�"�I��=,p�>M�O>�$l>��Y>�n">o�4>%���Hq%�D��^%w��B���	��{%���'�:�;D
�1�/�9��������R��혾�]�0Г�gIt���W��~�=�S?h�K?"i?�?��D��a0>�Iž1D=�#�g�>��>�+?��2?�+?�J�=�q}���h�������h����t>5��>	^�>ˢ�>�p�>���=OD>��Y>k�n>#�>�>G=�-=@5^=ajT>�\�>+��>+�>�C<>��>Dϴ��1��l�h��
w�;̽.�?j���F�J��1���9��צ���h�=Hb.?|>���
?пa����2H?/���)�˹+�w�>z�0?�cW?��>$����T�::>��Ħj�`>�+ �bl���)��%Q>zl?�e>�u>�E3��8�E�P��ְ�Fc|>k6?�	��mO9�a�u�)�H��HݾJM>z�>�I� �������&=i��y=dP:?%�?����43����t��؝��Q>�,\>�=pѭ=jTM>P�a��ƽ�G���2=�i�=T�]>f}?��;΁_�!��>��̾�a���c�>0�h>)��>z�I?!?��=i�Y�������޽��>���>ɟL>s>s��2}=h��>1�Z>҃�</l`�0j���
��>�2����^�ɾ/��B�=�潦)�<��=g ���dG�� �<�~?���(䈿��e���lD?S+?c �='�F<��"�E ���H��G�?r�@m�?��	�ߢV�@�?�@�?��L��=}�>׫>�ξ�L��?��Ž6Ǣ�Ȕ	�+)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿg�>bw�`Z�������u�D�#=���>�7H?�W��S�O��
>�Ov
?�?%`����ȿ�{v����>`�?{��?��m��A��F@�g��>��?gY?'ni>�g۾�]Z�#��>c�@?�R?��>u9���'���?$߶?ȯ�?�I>���?5�s?�k�>�2x��Z/��6���yn=��[;e�>�W>`���_gF��ד��h��l�j������a>��$=0�>�D�C4��y9�=s�I���f�/��>�,q>`�I>zW�>�� ?b�>���>�y=0n��>ှ����/L?:��?��>An�T��<-�=:*^�N<?�C4?��Q�)�Ͼ�ۨ>�\?�ր?[?
��>����#���ѿ��d��A�<�;L>��>E�>I����J>��Ծ	%D�#��>A"�>DL��Rpھ��������Ϝ>�X!?Ǚ�>L��=ۙ ?��#?��j>�(�>CaE��9��X�E����>٢�>�H?�~?��?�Թ��Z3�����桿��[�s;N>��x?V?sʕ>b���񃝿bkE�/BI�9���^��?�tg?rS�0?<2�?�??`�A?|)f>ׇ�)ؾn�����>�$?*4%�'B����!���?��	? ��>R%�В���&t�?��4o��	?�[?1�'?�z�+Z�)��S�
=�"޻|+�0�;'�輺�	>�m>�`���1�=�>{u�=��]�v�.��
�<a$�=9�>�F�=B+2�~�L�W�+?� 6� F��H��=�ir�$3D�/�~>��J>m,��X^?�N>��|�k��_r��:�U�潍?���?Ǆ�?H��Jgh��=?4�?@-?���>	J��K�ݾhe��|w�oPx��F�E=>�^�>�[|����񐤿Ū�LM���Ž�l`�1M?s4�>���>��>ea,>��>�Ϋ��)����g0��Fh�����-�p	1����E���3��@ϼ����{��3�>�Q��Ϙ>^��>���>,�>�=�>�� <Z!�>Ωm>q��>՞�>�F>��H> >�.�����>OR?o�����'�L��T���B?Bod?�q�>�e��d������?���?]g�?�v>�2h��+��V?�>���ln
?!j;=i��o�<����xF������V�Na�>��׽N�9��M�ZGf��r
?�H?�Ў��T̾|�ս֝�N��u?50?<�Y�M�Z�k`��\f��tq�=1��=�����*F�fj���4o������z&���=�i?I��?
��(��\�Ҿ��K�O�?��D�>��>��>{%><H.��.��@��1�1c?�D�?vk?���>(L?��:?txK?�FV?k��>�F�>�����9�>F�Q<Lp�>�J�>T�5?P ?�_0?�x?�1)?ta >�%�������h�>�T!?c?�(?L�?�)=�F���n)�<f��y	`�}w�����=��<�����K��-�1=�/>E?�$��9�G��_>��7?�	�>*�>`󄾾�i���=��>DW	?���>���,�i��t	��3�>���?0����v=��)>��=�֦��v�:<��=[��r��=�ǼiHZ��ܹp/�=��=wz$��)��o�;ϒ<�͋<_�>�� ?7i�>-�}>�n��X���w�&T�=lP>��I>,�>ճ��m��I嗿�i�1i>�5�?@Z�?r�=�)�=�(�='#���ҷ�
���ͽ�[�!=�?�� ?�lR?8��? b=?��%?�J�=q��{������q����?!,?܏�>a��ȹʾp憎&�3�&�?�V?�<a�3���<)�b�¾�ս��>9]/��0~���gD�
��_��fy�����?@��?75A��6�3q����#\���C?�"�>�Z�>�>��)�`�g�*&�x;>L��>�	R?
��>�P?�{?��Z?a�S>��8�U��F�� �:��J">��@?��?	��?dx?���>u�>h�(��ᾊy��m��4#��6���+P=�s`>Tܖ>q,�>���>���=�ʽ���T�;�Z|�=�m`>���>�>q��>�w>jy�<��G?U|�>9:þ�,�&����`��O���q?��?�.?Y]E=!��XyB����XW�>Z�?u�?a,&?�0M��>�]�&�¾)�D�;֛>s
�>���>�X)=�0=u�:>��>��>��8����2��	�-W
?N�=?[M�=�Ŀ6Q^���7��WR�D�@��渾��8����ں��2@�=�Є�|p(�f.���A��Ϯ�24������ ����l��D��>])=/��=$#�=����
˽s��;_1=���f�G=�S�==6�= Zt���#�����r<aǕ=�آ=�����ʾ�}?*�H?��+?��D?��y>eW>�&��>R{��?�rY>0+I�� ��D7�����G���yeھ��ؾ0�`�~S��"V>�.��o>��7>5��=��<���=�%=m��=3+ں�#=��=���=���=e��=.�>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>s��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>g8>��>��R�@L1��h\��:`�JiY�r%!?f�:�,˾~��>��=q,߾Ъƾ��-="�6>��i=`n�j[�(�=��z���7=��m=N��>�`C>��=3����=�L=��=�5O>"w����8�_6.��7=�x�=Mb>�J&>2��>M?�\0?#�c?T��>òm�"�ξ�ٿ�c��>Qf�=�ӱ>�	�=NC>)Ʒ>*�7??{D??yK?�ݰ>V�=5�>�>�%-��fl�E!㾛����+�<苈?���?K��>�)<c"?�K����>�b�½X�?��0?^�?�k�>�U����7Y&���.����ۀ3��+=�mr�dQU�����Fm�-�㽰�=�p�>���>��>,Ty>�9>��N>}�>��>�6�<ep�=~ጻ��<f ��a��=Þ���<@wżÛ���q&��+�&�����;���;N�]<[��;)?�=�}�>�j>J)�>�=p���d->3���(�L���=E䧾��B�5?d��G~��>/�8���C>�Z>"-��������?\>`�@>5#�?��t?�U!>T��l�վ� ��|{d�XaR� ��=��>?�<�o�;�Ea�sN�PҾuk>֕�>�9�>�;>fa�� -���O;l���+>�v��>�g��k�^�z��kKr�����)��+튿���<�EJ?��}�tA�=�i�?�8?�"v?}�J>�]�=���Nt>��*�6#�=2k߾��%�'�=ϔ3?��A?Sߏ>3J�.5��>��i�<Cw3>32þ��Z�]�f��4W�C-��B���,�'�!�t��_�n��M��?t��)m�����+?�Z}?�Ɨ?�ͽ������t��bH�c!�=��>��0?��>�b'?���>�j��/���[
�&[�=ܥq?�{�?+��?<�G>y��=7޶����>JT	?n�?��?��r?��6�,&�>��"<'�%>�Ӊ�I$�=��>M�=���=�A?�g?\�?�唽�Y
�Α��u�y�a��=�r�=̡�>���>֌t>"D�=�zq=�#�=݆Z>횞>��>L�_>?a�>#&�>Yc��Ъ���?v,�=�Aj>�4?��>&�=��`����=�r��8�t 1��%߽Nd��2�<=ۥk;<�Y=�`����>0�ÿ���?q��>w&�֕?]Ҿ�a��Z�H>��>����J�>�k�=+�>�y�>郦>�2>' z>��J>�]Ӿ�>S��S!�1C���R�L�ѾPz>ǰ��-&����H���vVI�l��l��j��,��#?=��L�<�B�?�����k�?�)�V���?U�>|6?i㌾A숽>�>���>>IG��=���<����;�9�?M��?)�^>��>��U?7?J�-�J0��H[��gv���A���d��na�s������
�%`ɽ��]?��z?��B?wj�<��y>@X�?��%�P	���n�>��.���:�3F=��>�.����\�d�վ�������GE>w?o?]�?��?e�W��H�=����k�>��,?��e?}8?
�5?e�_>�n'?��>��?w�?�~#?r�G?��?��>�-`��U���@J��K�<�u����Up�A��I�=1�<X�����%>��\����Դ(��q]���\=|���*<U:t2=??>AW>�	>�nd?ԥ*>�\��iWN?LO��Y�GT���>�큽�վ�����S�־}ഽ��?���?�o�?`�>bw�kF��b�h>eY�>w%">��(>��>�d��L���k=)�I>Z�B=U>ԝ ��q�ʞ�A���b6�v��=Al�>4|>�Y��$%>z���ELz���e>��O�*���Q�s\G��i1�.�t�Z��>�8L?w�?���=C��2���H�e�9)?{<?��L?9H?�	�=!ܾU�9��J�����>�;�<E=	�`����;��'�:�:t>ɾ��������`>��	��)ھ3l��1J�C��.=�.�TQ=��
��2վ�}�N��=�	>+��+ ��Ö��n����I?�Tk=頦��}S�������>o��>�M�>f)B�}|�w�>�9�<��=��>E@>t�{��G��F��&�ي">�P)?�!M?�N�?>���`�u'������7����&,?��q>}'�>:Ή>�,->0/������zU���j�K��>'�
?g�
�:7���龼���#����>�)?]�N>F:?��8?���>)�N?��??lP?S�>N�B<��ʾ�?@G�?��>�\���?���.-���;�%��>=f?q����*�>�O?B?�+?��U?�?xD->�+ξ7�H��ɒ>�>P]0��#����>T�z?�#�>.f?���?8>ƩD�_Ú��i�=�>�=�;">�C3?�/?0A-?x��>=�>�b񾲂d>"�>�d�?��?]�?���>���>$2�>��>|q�>���>�M?�F(?2�Z?>ut?�gI?<S�>3��=
��=��<�'>�[C1���q��=w�>���;�4�<J>C��Ҽ��߼.���y=J$=������ͼ髷=#\�>��s>�
����0>>�ľ~R����@>Տ���R���ኾk�:��ʷ=��>v�?6��>a#�G��=ٮ�>�G�>(��5(?G�?u?�S!;i�b�k�ھ_�K���>�B?Y��=��l�������u��&h=M�m?�^?�W��(��O�b?��]?@h��=��þz�b����g�O?=�
?3�G���>��~?f�q?U��>�e�+:n�*��Db���j�&Ѷ=\r�>LX�S�d��?�>o�7?�N�>/�b>'%�=iu۾�w��q��h?��?�?���?+*>��n�Z4�[��q����B?R	?J|���?��Ǽ�a¾�.0�+Q���g
�I�־�?Ͼ�]8��ݢ���^u��{T\�k�:���>M�K?�C?�6?�U��'^�O-g�����ecY�i��T>�<|U���k�e�`�����+�3���)�8��e;�ㄾ�<��H�?*?�)�ߨ�>�ѐ�\�����ؾ��>>��������=�|��-n0=4Y7=8+a��:�i	��^?���>��>��:?d�R�N8���2�S�7��M��x�7>X�>���>1�>�=/���R���¾�拾p����(s>�c?�`J?��m?����a1�����6W!��>�9��B>�S>��>`T[�����&�b�>���q�]��揾��	���=/Q3?��>��>&|�?��?��	��w����u���0��%k<��>�i?b��>A��>�3ͽUa!��|�>�5m?�)�=A�={K�ZJ	�~Ԉ�]�۽#��>���>整>p�>Z[I��mx��˘��a���B�dbY��_v?ei7�mA��a>^�]?�C����Z��>8�A�$���'�(�������>ۧU=,=>U���L���B�(�ؾN�>?��>:$��<B,�OI>=?��	?u��>�i�?_�>�t��B�>��?�X`?��S?POO?�r?h�;>� B<R M�z��[���>�>��g>�4N<��[=����9�Fl��{�=@�=�ep�� N��'��;�\�=z}�=-?>�cۿ�AK�G�پ����F�C
�W���?Բ��B���	�KԵ��N����x���c$(��&V��c�������l��g�?;�??�������`���~r�����\W�>��q��I�V���Z���N��|ᾧ���!��O�[i�U�e�Є'?������ǿĴ���ܾE% ?�' ?��y?P���"�4�8�"� >��<ka�����t�����ο1���9�^?���>���Ԕ��G��>Q��>��X>*q>L�������<)�?H�-?j��>��r��ɿ����vڤ<���?��@t}A?��(�N�쾇V=���>�	?��?>KN1��H����U�>�<�?��?2�M= �W�Ǹ	���e?C�<��F�7�ݻ'�=i9�=D=K��&�J>*U�>��TA��<ܽǸ4>yم>�|"���Q�^�{��<��]>�ս7��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=���ƿ��$�"{�o@=c�ߺu�[���Ǭ��U��(��4lo����R�h=g��=��Q>lg�>W>$/Z>�eW?��k?$L�>�t>5�%{��Wξ���I��k��⦋�P��		X�Ȭ߾�	����Y����ɾ�=����=�MR�֘��[� ���b��F��.?-7$>��ʾ
�M���)</�ʾ���(㌼so���h̾ʣ1���m���?f�A?�腿1�V�� ����G���W?��&���ͬ�+|�=|_��^e=���>�9�=���i 3��eS��s0?�\?����`��S!*>� ���=��+?Ή?�|Y<�$�>zI%?��*��P�jU[>?�3>�У>{��>E?	>���Y۽��?��T?���} ��1�><b��Z�z�A�`=u3>�>5�<��[>sȒ<X󌾏�U��8��2�<YEW?�S�>$*��wF��u��p>=��x?�?�5�>�jk?�C?X��<�%����S�5�
���z=�W?F:i?��>
"��-о�O����5?�e?&�N>
�h�#�龈�.��!��?��n? K?i���z^}�������b6?
�v?s^�xs������V�B=�>
\�>?��>��9��k�>
�>?#��G��ế�JY4�,Þ?��@���?[�;<����=w;?|\�>��O��>ƾ<{������+�q=�"�>����lev����R,�?�8?Ѡ�?���> ������)��=�ٕ��Z�?~�?���KAg<K���l��n���~�<aΫ=D�uF"������7���ƾ��
����⿼˥�>?Z@V�Y*�>�C8�L6�TϿ&��\оkSq���?H��>C�Ƚ����4�j��Pu�Y�G�.�H�å��N�>�>����_���r�{��q;�%%����>��
�>>�S�d%������U�5<��>���>���>q'���轾�ę?!a��T?ο����g��y�X?�g�?�n�?�q?T�9<��v�e�{��e��-G?:�s?qZ?�e%��9]���7��j?�]��?V`��4� HE��U>W!3?B�>5�-�e�|=�>���>3e>�$/�h�Ŀ�ٶ��������?\��?�n꾌��>���?Et+?=j��7���V��"�*���/�:A?�2> ���j�!� /=��ϒ�*�
?g}0?v�?/�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�#�>��?Gn�=�a�>@d�=���-�j#>p�=?�>��?5�M?cK�>�T�=��8��/�[F��GR�$���C���>1�a?�L?BKb>���� 2��!�Pxͽ�c1�bM�ZW@��,���߽�(5>��=>�>��D�Ӿ��?�o�4�ؿ	j���o'�q54?`��>��?����t�f���;_?�y�>77��+���%���C�$��?�G�?*�?O�׾�O̼�>��>9I�> �Խ����������7>�B?���D��(�o�S�>���?�@�ծ?_i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?Qo���i�B>��?"������L��f?�
@u@a�^?*C�������@���?S�:��=�z>�j>ʓ�V1>t��=�={�<Q>>�`�>.�u>.!�>n�>ÓA>��>� }��3 �x����Cx��yB�F�"��2�(����J��Wɾ{/�\����U�8v߽��p��&�%)ξ���֔��>&�=�~R?^nR?�Lp?���>�C��D">*���<#�����=��>0?��J?�,(?6.�=�9����d� ΀�'���·����>�`K>���>���>L�>��g���6>��9>��>K�>��[=oE�<�?=}X>hp�>ڷ�>)��>IC<>Ñ>Fϴ��1��b�h�w�̽!�?����Z�J��1���9��ষ��g�=b.?�{>���?пR����2H?���X)���+�;�>d�0?�cW?�>;����T�2:>u��צj�`>�+ ��l���)��%Q>Tl?Pif>Vu>O�3�b8���P�������{>�6? ���(B:���u�y�H�bhݾ�PL>�O�>��O�J���薿J�~��Yi���z=1�:?*�?�B������Mt��<���Q>�[>�T=~��=�L>�[a�]RŽ��G�ow.=���=��]>cP?��+>�ێ=��>�a���\P�_��>�[B>�,>>@?�(%?Ӕ��◽恃�1�-��	w>�P�>(�>�K>zNJ�ٯ=�f�>��a>���&�������?�]W>ݹ}��s_�Du�I?y=S㗽!�=Cb�=?} �(=�ߌ%=�~?���(䈿��e���lD?S+?d �=2�F<��"�E ���H��G�?r�@m�?��	�ߢV�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž5Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ ]�>Kg��Z����M�u���#=���>w0H?�P���O��>��u
?z	?�i�v�����ȿ�{v����>�?��?R�m��@��0@�I��>ʜ�?H`Y?�xi>j۾LZ�J��>��@?R?��>#;���'�`�?(ڶ?���?��@>�?��l?��>�m:�ǐ+��{�������u=H2<��>O�>%þ�"H��������pj����+�t>��7=�a�>���K����ˮ=	�������U~A��ͱ>n�r>�~I>~��>R�?"4�>T��>�=z���G����N����K?���?-���2n��N�<Y��=)�^��&?�I4?k[�|�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��L��<��K>*4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��TS��GB�>�e!?���>�Ү=�� ?��#?֔j>u'�>�`E��9����E�N��>���>�H?��~?��?�Թ��Z3�����桿��[��:N>��x?	V?�ʕ>\�������hoE��EI�����T��?2tg?�R�?2�?�??!�A?&(f>	���ؾK�����>��!?/�9�A�N&�6��~?�P?B��>u7����սzJּ��������?�(\?lA&?��,a�Q�¾\;�<&�"�&�U����;��D�)�>T�>抈�m��=�>װ=�Om�dF6���f<�i�=��>��=E.7��u��0=,?��G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>$�l���K���ڙ���F��_�Ž��d���>���>��?cX�>���;"P�>�+��`p7�]d��:վԀX�$���0�Q�'��/"��A��dZ�W��������;�>��=!A�>��>�o>5��;k��>�C2>,L�>��>r��>��?��>�j�>���>���+j;�!PR?����W�'�ϻ辤���a1B?'ud?�A�>Ǜh�������$�?���?�r�?�Ov>�th�`#+�.t?�D�>8��<n
?�#:=a��	K�<Z��t��t%�������>?=׽�:��M�5\f�e
?Y/?�G���z̾�*׽X����A�<��v?%?��/��"L�^�j��P���C��l��٨�௼�K�0�Ri�.m���9�?����4��9/<P"?mԍ?�� ���	�N����K� �@��{>J��>��>h��>O�I>�
��(F�I�c�);�O]�����>�{?�G�>�FH?�CE?H<?��J?���>��>��u���
?�O=���>L��>ΩN?D�.?#O=?��?�c2?���>�n�b�5� �>�?�(?e�$?W ?h~?f~ ���;���-�ݮٽ�x�8ھ<8h�<�m�=Mo����%��=��O>�?����9�������m>zd7?���>���>)񏾪����<V	�>'�	?��>�� ���r�m����>��?� ���=��&>���=[G������B��=����a�=6P}���9�mx<�Z�=���=��л~����b�:��;;ԇ�<�t�>6�?���>�C�>�@��(� �i���e�=�Y>CS>p>�Eپ�}���$��x�g��]y>�w�?�z�?m�f=��=��=}���U�����L������<��?8J#?(XT?^��?x�=?`j#?˵>+�hM���^�������?�Q+?��>�b�:�ʾ'���C�3���?x�?h%a�����(�ľ��׽��	> �/��p~�@���~C���b��v�u蚽X��?�ߝ?�>K���6��P�gn������=�A?:L�>�.�>���>�t(�36f������;>�F�>|pP?m�>��O?�:{?a�[?�NT>ϝ8�5$��ҙ���8���!>. @?ާ�?��?Oy?q�>.�>M�)��྿c���L�����₾��V=�Z>&��>��>o��>3��=�Ƚo���>��ݥ=�b>4��>ܯ�>%��>�zw>���<��e?_e�>��ܾJF�ر���[����t=�y�?u�?9�?�N�<��ľ����a��v��>߯�?�״?�S?-0e�H
'>$���E5߾������>�Γ>��X>�a�<�m(=�<a>�>J&�>6����388��n��'?Z�:?��=�н���Y��Q��'���=�j���Ȑ�yU�?�p��O�= ���$�轪@���w��l��r*��/����N��J%�w��>��=qXf=m�=��<�|����=*廼r/b=
���1<�1m;<2�;����͡�B1<�A^<fh��N;��z?�I?_p,?�B?�Xl>+�>�Ep��Ҍ>�"|�]s?��S>UJ�&Ӹ�k59��ͧ�����#�ھ�پN�]������>�7:��>��3>���=eo<���=��g=R��=4�l:PM==���=���=�ܺ=��=�@	>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�b7>sh>��R�6�1�� \��Fb�[�/|!?�9;��̾e�>lV�=:>߾��ƾ"N,=��5>��`=J���\��9�=e�y��*:=�!l=���>�zC>&�=����PG�=2J=���=1�O>`͊���7�'�-��13=���=�cb>��%>!r�>�?[[0?<d?Wa�>��n��Ͼ�O��F�>��=Yձ>���=��B>%��>�8?��D?��K?�]�>��=�>�f�>Xa,�J�m��8�E���s"�<��?6�?�ڸ>� P<M2A�dH� 1>�`Ľ�?%U1?ߏ?$�>�U����9Y&���.�$���Ă4��+=�mr��QU�M���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����='�����<�vż�����u&�8�+�-�����;p��;?�]<O��;���=W��>?@>��>���=<
���E/>7���]�L�T��=�E���+B��3d�|H~��/��X6���B>J7X>����J3��a�?�Y>�o?>��?@u?��>�'���վTP��O@e��PS��ո=�>��<�x;��X`���M�M}Ҿ8�>�W�>�X>7�:>2�ɳ@���=�_Ҿ�R:���&>���-2�}}K�u4}�,���ݠ��Cr�)�<�3?�rv�\�=mZ�?Vz]?epq??r�>��#>�ᾒd=����N��=�	�oe��� �=� 0?��!?�U?�����O��I̾FC���o�>��I�z�O�մ����0�T ��ڷ��>���� Ѿ� 3�8o�������B�f�r��Ϻ>(�O?�ڮ?�)b��.���O����Ș?8\g?�>�?c>?�}����Q2���(�=m�n?��?s/�?�n
>�Խ=�ݵ���> �?���?��?Vss?F�;�C �>!��;4 >���M�=b�>8��=s��=��?��
?_>
?L���!
�;�����i\�M��<I�=I}�>8t�>�Lr>�Z�=��q=nk�=�YZ>aϞ>��>*d>1��>?;�>�R��C��"q'?���=yp�>̴/?�L�>�y?=�4�����<��?�bu?�-,��9����v٪<I�q��F=�Z�b�>��ƿV��?_V>ϗ�E�?���L�L���N>��X>��ٽ!,�>^�J>�>�)�>�Ŧ>ҷ>}��>M�#>�(��j�>7�K3�Y�/\�����R�<TS���@�=�*�8�U��4Ͼ���H��5�l�H�R;@�0'>�c�?���=T�i��W�*8>lh?L>�=��?ǟ��x�M=}�>[b ?��>��r���׎�����{y?*0�?�:c>��>L�W?8�?ɒ1�@3��uZ�0�u��(A�e���`�o፿����ӗ
������_?��x?�xA?�L�<>:z>)��?��%��ҏ��)�>�/�';� =<=+�>�)��|�`���Ӿ��þ`6�JF>��o?)%�?Y?UV���_�+0>g@?<7.?~�u?�7?:�<?���s�%?�`<>E�?1?��<?��.?��?5�E>��
>lg�<Q�=38��᱑�����n������*=0߰=�$�<�j�<�@=~�<~G��R�����}���ۭ<cj:=�9�=w�=U��>-�]?$U�>���>��7?���r8������./?��9=�������������>��j?���?�eZ?r]d>�A��%C�,>�[�>و&>�\>�n�>fG��E�*؇=�.>�p>�=\�M��Ł�!�	�t���N�<�&>:��>�-|>���{�'>v|��0z�{�d>�Q�˺�?�S�b�G���1��v��Z�>��K?��?E��=U_�`.���Jf��.)?�\<?sNM?��?��=��۾��9���J��A���>P8�<��������#��6�:��f�:H�s>�2��Kʦ�-+j>���־GQl�NK����ηA=2���CI=���9\ھ.4��_��=F;>���ܣ#�b����Ԫ���G?��G=|.���/@�����)Y>��><��>�rW��n�y�:�m9�����=�V�>��:>�������F�������=	`\?�e�?_�?�ܾل��X<S�ݦ徬�Ⱦ�<4�F?��>o��>I�
>c�=�3��7� ���v���o���>\�?_3����J������]�f�E��hz><g?��!>�M�>q�t?�8$?V?�wY?��?��x>X��������?f(�?2�f>����R4�x�?���R����>�R?�o2�>׷?�W?�1?,�M?�
?�E>���3�G��O�>�SQ>?j�夿]�>%�x?5�>�e?x4�?EU�=��K��ih�����5=aK>�e=?�^?M?���>O�?������Q�h˧>nm$?:�n?y�r?y��>j?���>���>5�]>i!�>	��>��>i�<?j�5?`P?�,�>aAY=>�	�s��g�ݽg��=uf�G
�<��>���<�T+��Q$�0�<A�A>���=�Q>z���}G��ɶ�򨊽���>@ks> ���l0>��ľ8��*MA>Ϧ������p\���:��}�=���>W?���>+�"���=��>z�>v����'?��?/?��:�ub���ھ_L�Z�>�B?���=ixl������"v�`�g=K�m?�^^?�PW�Х��O�b?��]?@h��=���þy�b����h�O??�
?"�G���>��~?i�q?W��>��e�#:n�(���Cb���j�'Ѷ=^r�>GX�R�d�~?�>f�7?�N�>7�b>J%�=ku۾�w��q��c?��?�?���?�**>~�n�T4�=8��R��ڽk?e��>���1�?�,�x��ȿ� �������ľy�ž�k��Io;*\�L����1��o�=R�.>�5:?�|F?�Y?bK�9Q]��W�2�������ي:�Q@���a�D�a��BP��Ɋ���M���c��n)�=񛧾o(�/԰?e�2?~Ti�"!�>wƅ��	�I�߾��%>9����-?���f=Cq��2�����<(V������n�о��?Q/�>h��>G�:?��\��I�*"-���#�4�W�>>���> �>}��>�6 �!��q�m���l�6��0�\>�He?��L?�k?�|޽�c1��������=�_s���/@>&>Zm�>1�T�C��z!�2h=�!�u�9��f��	���/=��6?0��>��>�I�?NE
?���Uz���l�-�&��w`<�v�>KDd?�X�>ߎ>b�ݽ&��e�>�v?(޶>{-+>٭Q�8�](~��_�8��>�T�>H��>ǝ=t�M�"g����yp���X3���y>��y?��w�ulE����>��e?wE{�6}4����>K���N��پQ���2>x�?�=�B>��;E<�ٞ��P,����J?N?�>&�g�d
<��p>.\�>��?a�?��?#��>��@�>Ϝ>\i<?��r?p�|?_^?��>g��=D��j�B�v�H;}\>�v�=���=Eـ�	�4�a��6�j�ِ��P�
>pcC=�Q��E=��=Gq����1=��K=E�>�lۿ=@K�a�پg���^C
��䈾(����g����R[�����Wx����''�V�}5c�릌���l�5��?�;�?Pz��K.��F���7����������>��q�.o�X竾���+.�����X����a!���O�I$i�5�e�P�'?�����ǿ񰡿�:ܾ5! ?�A ?7�y?��5�"���8�� >EC�<0-����뾬����ο@�����^?���>��/��q��>ܥ�>�X>�Hq>����螾�1�<��?7�-?��>ǎr�0�ɿb���o¤<���?0�@�A?-)�7r�$K\=���>��	?�B>�A0��K����j|�>^ �?���?*A=��V����S�d?� <�TF��E��2��=>��=��=e���I>e��>���W�B��ٽ�5>���>�`"�C�_�I��<��\>0�ֽAݐ�6Մ?{\�sf���/��T���T>��T?+�>�:�=��,?G7H�Q}Ͽ��\��*a?�0�?��? �(?&ۿ��ؚ>��ܾ��M?dD6?���>�d&��t����=7�Ί��L���&V����=3��>�>�,�����O� I��[��=V�'�ƿ.�$�	}�K_=�yݺޤ[�c~�`�����T�n#���fo�+�轒�h=��=��Q>ml�>�%W>Q4Z>gW?j�k?�N�>��>�7�U���ξL|��G�����������]��R��߾{�	������g�ɾ�!=�!�=�6R�����|� �Y�b���F���.?�o$>-�ʾ9�M�0�,<{rʾ�����	�*̾X�1��n�N̟?k�A?������V����Pg�os��_�W?�P����|款z��=(k��^�=�#�>i��=���@!3�X}S���3?�?����9��'>6����^=�-?�x?��=�ʩ>�'?L����U�>2vS>?W�>
�>��>Jڦ����Ӊ?c�M?)b���%���_�>֖��\˂����=�8>?6�:��\�[>�4/<t������5p��"Ǡ<X1W?V��>*�C��J���,�B=_{x?��?wĠ>�bk?C?F$�<����=S���
���v=ˋW?�i?&	>sj���Lо�㦾+\5?�Qe?�JO>��h��܇.���Q0?|�n?0?�����|��풿f��x6?:�v?zr^��s��/���V��=�>yZ�>Y��>��9�
k�>C�>?�#��G��ĺ���Y4��?��@���?<<�����=:;?�[�>��O��>ƾ�z��񂵾ƚq=�"�>&����ev�`���O,��8?ɠ�?���>ܓ������~�=����W�?
�?�ê���S<����l�y���J�<x�=l��Z#�/���7���ƾʩ
�����9�ż�>lO@'��!�>�W8�W4�R_Ͽ\����оB�p���?ȅ�>�tɽ������j��$u���G���H�ӓ�>FQ>1������:B{�I�;�����S�>@P���>?�P��������=<T)�>Y@�>˽�>�
��t��ގ�?�.���1ο�o���,���Y?�s�?�v�?��?*<ay�Źy��c�;�F?�Ls?;8Z?Z� �$\�w�-��j?h_��|U`� �4�_HE��U>�"3?�B�>V�-���|=}>J��>�f>�#/�x�Ŀ�ٶ�!���_��?��?�o���>w��?}s+?�i�8��k[����*���+��<A?�2>����,�!�G0=�OҒ���
?&~0?`{�^.�]�_?+�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>c����8Ǿ��<���>�(�>*N>_H_���u>����:�i	>���?�~�?Qj?���� ����U>	�}?\$�>��?o�=�a�>`d�=B�*-��k#>�"�=b�>��?��M?L�>EW�=z�8�~/�:[F��GR�]$�5�C��>y�a?�L?Kb>���q2��!��uͽ�c1��P鼜W@�=�,���߽6(5>��=>�>Q�D��Ӿ��?�9�:G׿1ѝ�O ���3?��>y۶>�� ,��39?��	>����,��䍿�~
=,��?>F�?��?&����j2�=#��>�>?��ʀ+���4�I�x>]�D?PF^���x�8?D���|>��?+�@7�?�5b��h?��j����~��3���5����=k�6?�*�~�x>���>PZ�=u�v�.���t�s�0M�>$n�?>��?���>p]l?o��C�Ud,=>]Ok?�?��C�*��|�D>��?��S����C�d�e?�
@�e@H~^?Kâ�v���h���-*#��q��0S�=\y�=���=��ʽ-"�=���;c�<{�"�I��=,p�>M�O>�$l>��Y>�n">o�4>%���Hq%�D��^%w��B���	��{%���'�:�;D
�1�/�9��������R��혾�]�0Г�gIt���W��~�=�S?h�K?"i?�?��D��a0>�Iž1D=�#�g�>��>�+?��2?�+?�J�=�q}���h�������h����t>5��>	^�>ˢ�>�p�>���=OD>��Y>k�n>#�>�>G=�-=@5^=ajT>�\�>+��>+�>�C<>��>Dϴ��1��l�h��
w�;̽.�?j���F�J��1���9��צ���h�=Hb.?|>���
?пa����2H?/���)�˹+�w�>z�0?�cW?��>$����T�::>��Ħj�`>�+ �bl���)��%Q>zl?�e>�u>�E3��8�E�P��ְ�Fc|>k6?�	��mO9�a�u�)�H��HݾJM>z�>�I� �������&=i��y=dP:?%�?����43����t��؝��Q>�,\>�=pѭ=jTM>P�a��ƽ�G���2=�i�=T�]>f}?��;΁_�!��>��̾�a���c�>0�h>)��>z�I?!?��=i�Y�������޽��>���>ɟL>s>s��2}=h��>1�Z>҃�</l`�0j���
��>�2����^�ɾ/��B�=�潦)�<��=g ���dG�� �<�~?���(䈿��e���lD?S+?c �='�F<��"�E ���H��G�?r�@m�?��	�ߢV�@�?�@�?��L��=}�>׫>�ξ�L��?��Ž6Ǣ�Ȕ	�+)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿg�>bw�`Z�������u�D�#=���>�7H?�W��S�O��
>�Ov
?�?%`����ȿ�{v����>`�?{��?��m��A��F@�g��>��?gY?'ni>�g۾�]Z�#��>c�@?�R?��>u9���'���?$߶?ȯ�?�I>���?5�s?�k�>�2x��Z/��6���yn=��[;e�>�W>`���_gF��ד��h��l�j������a>��$=0�>�D�C4��y9�=s�I���f�/��>�,q>`�I>zW�>�� ?b�>���>�y=0n��>ှ����/L?:��?��>An�T��<-�=:*^�N<?�C4?��Q�)�Ͼ�ۨ>�\?�ր?[?
��>����#���ѿ��d��A�<�;L>��>E�>I����J>��Ծ	%D�#��>A"�>DL��Rpھ��������Ϝ>�X!?Ǚ�>L��=ۙ ?��#?��j>�(�>CaE��9��X�E����>٢�>�H?�~?��?�Թ��Z3�����桿��[�s;N>��x?V?sʕ>b���񃝿bkE�/BI�9���^��?�tg?rS�0?<2�?�??`�A?|)f>ׇ�)ؾn�����>�$?*4%�'B����!���?��	? ��>R%�В���&t�?��4o��	?�[?1�'?�z�+Z�)��S�
=�"޻|+�0�;'�輺�	>�m>�`���1�=�>{u�=��]�v�.��
�<a$�=9�>�F�=B+2�~�L�W�+?� 6� F��H��=�ir�$3D�/�~>��J>m,��X^?�N>��|�k��_r��:�U�潍?���?Ǆ�?H��Jgh��=?4�?@-?���>	J��K�ݾhe��|w�oPx��F�E=>�^�>�[|����񐤿Ū�LM���Ž�l`�1M?s4�>���>��>ea,>��>�Ϋ��)����g0��Fh�����-�p	1����E���3��@ϼ����{��3�>�Q��Ϙ>^��>���>,�>�=�>�� <Z!�>Ωm>q��>՞�>�F>��H> >�.�����>OR?o�����'�L��T���B?Bod?�q�>�e��d������?���?]g�?�v>�2h��+��V?�>���ln
?!j;=i��o�<����xF������V�Na�>��׽N�9��M�ZGf��r
?�H?�Ў��T̾|�ս֝�N��u?50?<�Y�M�Z�k`��\f��tq�=1��=�����*F�fj���4o������z&���=�i?I��?
��(��\�Ҿ��K�O�?��D�>��>��>{%><H.��.��@��1�1c?�D�?vk?���>(L?��:?txK?�FV?k��>�F�>�����9�>F�Q<Lp�>�J�>T�5?P ?�_0?�x?�1)?ta >�%�������h�>�T!?c?�(?L�?�)=�F���n)�<f��y	`�}w�����=��<�����K��-�1=�/>E?�$��9�G��_>��7?�	�>*�>`󄾾�i���=��>DW	?���>���,�i��t	��3�>���?0����v=��)>��=�֦��v�:<��=[��r��=�ǼiHZ��ܹp/�=��=wz$��)��o�;ϒ<�͋<_�>�� ?7i�>-�}>�n��X���w�&T�=lP>��I>,�>ճ��m��I嗿�i�1i>�5�?@Z�?r�=�)�=�(�='#���ҷ�
���ͽ�[�!=�?�� ?�lR?8��? b=?��%?�J�=q��{������q����?!,?܏�>a��ȹʾp憎&�3�&�?�V?�<a�3���<)�b�¾�ս��>9]/��0~���gD�
��_��fy�����?@��?75A��6�3q����#\���C?�"�>�Z�>�>��)�`�g�*&�x;>L��>�	R?
��>�P?�{?��Z?a�S>��8�U��F�� �:��J">��@?��?	��?dx?���>u�>h�(��ᾊy��m��4#��6���+P=�s`>Tܖ>q,�>���>���=�ʽ���T�;�Z|�=�m`>���>�>q��>�w>jy�<��G?U|�>9:þ�,�&����`��O���q?��?�.?Y]E=!��XyB����XW�>Z�?u�?a,&?�0M��>�]�&�¾)�D�;֛>s
�>���>�X)=�0=u�:>��>��>��8����2��	�-W
?N�=?[M�=�Ŀ6Q^���7��WR�D�@��渾��8����ں��2@�=�Є�|p(�f.���A��Ϯ�24������ ����l��D��>])=/��=$#�=����
˽s��;_1=���f�G=�S�==6�= Zt���#�����r<aǕ=�آ=�����ʾ�}?*�H?��+?��D?��y>eW>�&��>R{��?�rY>0+I�� ��D7�����G���yeھ��ؾ0�`�~S��"V>�.��o>��7>5��=��<���=�%=m��=3+ں�#=��=���=���=e��=.�>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>s��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>g8>��>��R�@L1��h\��:`�JiY�r%!?f�:�,˾~��>��=q,߾Ъƾ��-="�6>��i=`n�j[�(�=��z���7=��m=N��>�`C>��=3����=�L=��=�5O>"w����8�_6.��7=�x�=Mb>�J&>2��>M?�\0?#�c?T��>òm�"�ξ�ٿ�c��>Qf�=�ӱ>�	�=NC>)Ʒ>*�7??{D??yK?�ݰ>V�=5�>�>�%-��fl�E!㾛����+�<苈?���?K��>�)<c"?�K����>�b�½X�?��0?^�?�k�>�U����7Y&���.����ۀ3��+=�mr�dQU�����Fm�-�㽰�=�p�>���>��>,Ty>�9>��N>}�>��>�6�<ep�=~ጻ��<f ��a��=Þ���<@wżÛ���q&��+�&�����;���;N�]<[��;)?�=�}�>�j>J)�>�=p���d->3���(�L���=E䧾��B�5?d��G~��>/�8���C>�Z>"-��������?\>`�@>5#�?��t?�U!>T��l�վ� ��|{d�XaR� ��=��>?�<�o�;�Ea�sN�PҾuk>֕�>�9�>�;>fa�� -���O;l���+>�v��>�g��k�^�z��kKr�����)��+튿���<�EJ?��}�tA�=�i�?�8?�"v?}�J>�]�=���Nt>��*�6#�=2k߾��%�'�=ϔ3?��A?Sߏ>3J�.5��>��i�<Cw3>32þ��Z�]�f��4W�C-��B���,�'�!�t��_�n��M��?t��)m�����+?�Z}?�Ɨ?�ͽ������t��bH�c!�=��>��0?��>�b'?���>�j��/���[
�&[�=ܥq?�{�?+��?<�G>y��=7޶����>JT	?n�?��?��r?��6�,&�>��"<'�%>�Ӊ�I$�=��>M�=���=�A?�g?\�?�唽�Y
�Α��u�y�a��=�r�=̡�>���>֌t>"D�=�zq=�#�=݆Z>횞>��>L�_>?a�>#&�>Yc��Ъ���?v,�=�Aj>�4?��>&�=��`����=�r��8�t 1��%߽Nd��2�<=ۥk;<�Y=�`����>0�ÿ���?q��>w&�֕?]Ҿ�a��Z�H>��>����J�>�k�=+�>�y�>郦>�2>' z>��J>�]Ӿ�>S��S!�1C���R�L�ѾPz>ǰ��-&����H���vVI�l��l��j��,��#?=��L�<�B�?�����k�?�)�V���?U�>|6?i㌾A숽>�>���>>IG��=���<����;�9�?M��?)�^>��>��U?7?J�-�J0��H[��gv���A���d��na�s������
�%`ɽ��]?��z?��B?wj�<��y>@X�?��%�P	���n�>��.���:�3F=��>�.����\�d�վ�������GE>w?o?]�?��?e�W��H�=����k�>��,?��e?}8?
�5?e�_>�n'?��>��?w�?�~#?r�G?��?��>�-`��U���@J��K�<�u����Up�A��I�=1�<X�����%>��\����Դ(��q]���\=|���*<U:t2=??>AW>�	>�nd?ԥ*>�\��iWN?LO��Y�GT���>�큽�վ�����S�־}ഽ��?���?�o�?`�>bw�kF��b�h>eY�>w%">��(>��>�d��L���k=)�I>Z�B=U>ԝ ��q�ʞ�A���b6�v��=Al�>4|>�Y��$%>z���ELz���e>��O�*���Q�s\G��i1�.�t�Z��>�8L?w�?���=C��2���H�e�9)?{<?��L?9H?�	�=!ܾU�9��J�����>�;�<E=	�`����;��'�:�:t>ɾ��ݠ�=Ub>O��$v޾��n�J�?���rM=C��/V=��g�վ�0�կ�=%
>������ �`���ժ�b/J?��j=�z��X_U��q��h�>��>�֮>��:�h�v���@�����-�=��>�;>�8��% �~G�w4��C�>ILE?�U_?_j�?&��Us���B�͕��Y��>hȼ��?�{�>-l?�*B>�
�=*�������d��G���>A��>5����G�B���*��S�$�g�>�&?�>��?O�R?��
?��`?� *?d>?&�>V/���긾bB&?%��?G�=�Խ��T�4 9��F�S�>|�)?��B�[��>݊?��?��&?|�Q?��?X�>k� ��D@����>eY�>d�W�)b��� `>ìJ?3��><Y?�Ӄ?��=>��5�Tꢾ4ѩ�Q�=N>��2?T5#?��?M��>wJ�>`ͳ�;מ=0�>��U?ъ�?�_?)�>՜�>)��=y �>L�{=�1�>�-?A*?vI??�f?g<6?j�>�;�<���᳼�I3�uR�<:��P=�>k��&�Ӽ�:���<��Z�&J =f�=�_���X�Ϻ\��U��DW�>*�s>��� �0>��ľ�L��m�@>���<T���֊�I�:�^ٷ=ׇ�>`�?쬕>�S#��В=ȭ�>nG�>D���3(?-�?�?��;��b�E�ھ��K���>IB?���=��l�|�����u�u�g=��m?�^?��W�#"��)�r?�/n?�-���<�	Q�S�����.�T?.�7?�~1�0ߤ>Ц�?�r>?`��>|x�����裿w���m��0�=J��>���ڜ� ��>!GR??f�>���>��2�MM���Y�Ϭ��*X>W��?U�?y�?L��;�~p�{ݿ_�߾֚���3R?�:?���G:?�Xz<������R�q�כ2���˾Xr�ڝ��,�u;���-�r�0>��+?��_?<�?�\?� ��eT�^=P�`���]R?��������ܬG�/tP��rY�E��(P'�	8 �1_��{��<��۠A��#�?��'?V3�1�>�������d8˾��A>�~��|i�S��=����=xA=�+[=j�g�F�.����X ?X��>�\�>��<?�B\��Z=��L1���8�Ao���6>|��>hy�>�8�>u[[���0����1�ʾ�*����ѽL9v>Sxc?,�K?�n?n�*1�����[�!���/�|b����B>�m>伉>!�W����	:&�CY>���r�����w��T�	�-�~=��2?9'�>���>�N�?4?(|	��j���hx�P�1�b��<1�>� i?�?�>=�>oн�� ����>�ko?I��>�#�>T엾�C��d�y��y�>e��>a��>&��>2�U��5o�*��U��#�6�mN�=4�l?f����O��ܑ>e5B?����uM��Hl>݅��i�꾑\޾����i�>�r?�	�=���=�U��w�-�n흾�1)?�s?�F����)��K~>��!?0�>�=�>��?� �>�����;i�?�	^?|�I?B�@?�	�>��=����	"ν�(�<k0=%��>!E[>�,={
�=,��]��N#�vAU=G0�=�'Ƽ�(����<2ʼ_�Z<;_�<�7>8lۿ2BK�;�پ\
���-?
��刾����e������a������Ux����N�&�+V��2c�W�����l�v��?<�?.����.��%�������`���ᱽ>�q�@�������*��W��l����c!��O�&i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�}A?]�(����	aV=���>�	?|�?>�M1��E�w����R�>�;�?9��?y6M=��W��
��{e?�T<��F�ό޻��=�E�=_@=���[�J>(O�>E��%CA��;ܽ�4>�>oZ"�_����^�G�<͂]>.�ս�E��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=���d,ƿ�$����Z=Z>�f�Z����j���9 Y��ꟾ,p�͆���u=~Q�=�S>�ۇ>��W>�KZ>�tV?��j?%"�>Z>dX������ ξr�#�����8��7��6������E�8߾4������L���Ⱦ� =���=�6R�/����� �*�b���F���.?vu$>�ʾ[�M�W�-<�oʾ/���,ׄ��ߥ�Q-̾�1��!n�͟?��A?����O�V����DN�+���
�W?�O�����鬾.��=�����=+%�>���=���� 3�p}S�k11?�� ?5	�����\X2>f�ݽ�˦=E\8?,?Ԛ[=k[�>�k,?�,%�Z�ͽ��c>݄:>�v�>(��>���=�_���q���? �Q?���|�Q��>�	Ǿt�����<�8>+��w^��^>�=֑���;_h����=)7W?Q֍>u**�ݧ�m��Ut"��i>=Ӕx?�v?9f�>+Fk?��B?�ݨ<������S�i+���u=мW?I6i?@>�����Ͼ Y��ؒ5?EDe?&�N>�\h��R龌�.�7�j[?�#o?�??�Ҥ�p�}����%��`6?m�v?/W^��f�����lV��4�>		�>G��>��9����>�d>?�#��M��G���vo4�N��?Ϙ@j��?�54<U����=�8?mv�>ƁO��.ƾ�3���e���p=j��>�����fv����t,�U~8?餃?���>��������>����?\�?����^�<�������yܾ�Z>�����n����fX�3X�2k��8O)��㷾�{$=��>N@��>'}�>��>���￨�ƿ��`�ˡ#��+L�{�9?n�=n]�2��?���e��X�!'7���g��S�>��>ޭ��q�O�{��p;�>ҟ�]
�>j��
�>��S��-������>3<Nܒ>���>��>�Ү��齾�Ù?e��@ο줞�{����X?qh�?�l�?�k?C'9<a�v�n�{� .�a+G?��s?�Z?۴%��C]�Z�7���j?�w��ӱ`���3�59E��	R>.3?� �>�]-��]�=��>��>Q�>��/�5xĿ�ζ�����Ц?�{�?t�꾞��>�V�?+O+?_��E��2O����*�`��:�1A?��2>ཾ��� �=�����	?�90?�
	���]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?7̿>T}}?�
>�j?��>������=>�>{�$>������?2)G?i��>��=+ �A�.�h�D�MvJ�1���F@��'>�Z?��8?�>>����*��6��_O����o�<�.����4e�,�@>�1�=�>d������?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�{.?M��s_�&����;��D�5��i�K�>!�v�?��{>,W�F��S7��n����>�ѳ?�'�?��>ݪb?gt��s?���>���>rf?1�>�DH��0��J��B>Fl/��݀�f���@?Y�@��@ʳ^?P���4п�ڗ� X���&ƾAb�=�כ=�|:>ǎȽ�i�=��k=<��м�>��>�|u>''�>f�A>�9>N\I>�@��u�&�����G��
�K��.�m���:}���
�G�����,վ-�վYM���񒽭�k���@�ˇ	��զ�ݦ	>.aU?�zQ?�e?P��>�"$��>>��ݾ�+ =y�����=P��>DN*?�G?]*?�ܩ=&���`c���ŭ�ͽ�����>��f>t��>y'�>%�>U)����=>M�>l�>���=��O=���9�D3=��7>��>x��>���>6h>>`�>k״�q_��,;h�__x���ͽ�
�?-��.DJ����;������(�=_
.?ܗ>�I��jcпSJ��5�G?���a���*-��
>��0?
DW?J`>�P����V���>#q	���h��  >����6g�&)��|P>W�?��f>�qu>Uu3�u8�
�P�L����I|>�M6?¶� �8���u�iH�[ݾxhM>P��>X<�@k�(��%��i�L�x=R�:?K�?d��,n����t��%��.HR>��\>S�=C}�=��L>��e���Ž� H��.=	�='9_>��?�k->�ۗ=D��>9����L� J�>�L>)->��>?�p%?i8�U���%Z���!)��s>
�>�|>� >
M��b�=�>��a>���tᆽ��G�G�i`P>u�����Y���m�D�x=�ʏ�L��=�L�=�����=�Q�4=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾQh�>wx��Z�������u�`�#=R��>�8H?�V����O�g>��v
?�?�^�੤���ȿ5|v����>X�?���?g�m��A���@����>:��?�gY?roi>�g۾9`Z����>ӻ@?�R?�>�9���'���?�޶?֯�?�I>���?y�s?nr�>�>x�k^/�h5�������=�l];,c�>�a>�����iF�"ؓ��i��S�j����4�a>ۓ$=��>�<佟8���.�=G닽�M��¾f����>h)q>��I>�\�>� ?�f�>+��>�a=v���瀾������\?�l�?=���B��u�=p���]?���>?��?��>�ђ�n\?��?^{_?)n+?A��>W1<��ۣ���ӿB��򽥗�>T�?Ǐ�>$�=S��>#䐾|H�K��> 6�>��Y<����;N�=&P�>- ?�?��d>��1?<;4?*%:��?�>�yA���u+��W�>4�?�('?O4R?��?R�x[�閕�苮��9Y�o�
>�7r?r��>��>=
p�i)���z����z2g�;.[?l��?��{��?+d�?J&?!�I?�1>a`��@ȾU����=��!?����A��&�aR�%�?bO?���>�+��� ؽ4�ͼʞ�j�����?�.\?p�%?����a�׬¾��<�l0��4�����;h6�޳>�<>ʉ�[/�=�>,��=KEm��6�N-[<8��=ܩ�>��=8�6�ַ��3E,?;�C����㲙=N�r��D���>�HL>����_�^?i�=���{������|��X-U���?֑�?_f�?0s���h�$=?1�?�?��>�q��$n޾���j�v��>x��_��]>Z4�>!�m�1� ��������O����Žg�N��>[��>~�?�b ?�0O>J^�>Bݘ��'�e����<�^�0J��>8�w�.� |������#�K���¾��{��ޘ>���u�>z�
?6.h>Q�z>$��>ڕѻMa�>��R>M�~>�>m!X>��4>�� >��<�Ͻ�JR?������'�ɫ辉���~1B?nsd?�8�>��h�l������v?���?vq�?R<v>�}h��,+�~j?F;�>����j
?/k:=�f�0�<�X�����9c���f����>=/׽:��M��cf��g
?�*?\��S�̾�0׽�u��a>�S�? �"?��b��rY�f��s��~k��Y=Y>N�d6��l�L�6z�� 4��y���x�F�#�m�$>�'!?��?r�����%�D �@�s�E�j�k�>ĳ�>O�>���>�=0��'�~�(�>�O���5��Q:��� ?GQl?��>�I?��=?�t3?XbI?܂�>���>�,���>�6�=�F�>�?�F?#?K�.?v?Į?�m�=[�1�G�!��9(�>pX1?�v;?�?���>���o���|[�ҫ =І��D�<j�=�K�<�<�F���<?�>�?�7��8����Jo>.l8?�;�>���>�̑��X����=���>:A?c��>e����p�Y����>f��?�D�	I�<��'>���=g�%����:���=漬�=7Qc�v4)��8<p5�=p�=e�)�h;/�N;�6�;�e�<�\(?��2?�+�=+�?��`����~��U=�A��`�=U� �����������Q�{G�>Y4?�u�?���04>�@=o�6���<5��҄�p2�>0?�:�>��M?Y��?��P?d#{?�TH>��e��&�����M���v?RR.?�&�>4��m��uT��]	9�*y?�?w!^�(��*O(�VþﭽaA�=J0�c~�[i��'e?�i��<6��9m��~?�?뷛?�_�n�:�G	�D�������C?56�>cʵ>V�?�y(�> k��� �6>�N�>�mO?�$�>��O?�:{?Q�[?�gT>�8�v.���Й�Q�3�J�!>g@?^��?��?ay?-y�>"�>#�)��N��,�����悾��V=eZ>F��>,$�>��>ٽ�=�Ƚh��+�>�^�=��b>���>��>y�>��w>-I�<��H?q�>�m��-��7�n�%�z�,:(���Y?�Œ?�e4?����,��zU�3;����> }�?��?�<@?~���Y>���ئ�/�#�A2�>��><��>���=����dm�4�>�'�>q��C���0��<c!?d9?�G �?���hl���\��O��t��<����g.O���=��@p��'=c"��[���t��+O9�S���q��]��3��	�f��;�>
|=�
�=l�=c`¼kF��	�<�
�<���<n0<<<�h��f=�Ҏ�6��t�{�D���1�L��<�l<wiȾk�|?��H?��+? D?([{>�>�����>Ʌ��X?,�X>�[>�=����7��5��zݕ��پ��վ�e�������>-G��Y>2�/>��=��$<6��=�[q=��=���ք$=Ь�=���=`��=�K�=��>�>�6w?W�������4Q��Z罤�:?�8�>e{�=��ƾp@?{�>>�2������zb��-?���?�T�?@�?@ti��d�>M���㎽�q�=L����=2>���=u�2�S��>��J>���K��2����4�?��@��??�ዿТϿ?a/>n'> ��=vL��6.��@X���f��zJ��!?�W:��ZԾ2�~>��=�bؾ�,�� #C=�b8>jn�=�m�y�V�DŢ=b����s�<�}�=�,m>�wR>T��=Y�㽞��=_�.=u��=��k>�9��$u����R�=��=�6N>�9>���>�?�a0?$Xd?+6�>sn�sϾ�>���H�>��=�E�>=�=�rB>S��>P�7?I�D?��K?���>���=5	�>��>�,���m��m��̧�J��<`��?�Ά?IѸ>��Q<h�A���fg>�20Ž�v?S1?�k?X�>��ڿ,k��)���S�l%9���j���
���Ѿ�B־uF��B���a���a>{(�>�T�>��?��>2'X>6}�>H��>�>���<sG�=R�<J�=��d;��=�+�<��<��y����=e=ʽ�A�q��<v�e<��<7+����=���>�6>���>m��=�	��E/>+�����L�@ƿ=H��-,B�v3d��I~�\/�9X6���B>�;X>w��#4����?��Y>-m?>���?�?u?��>� �^�վQ���@e�PS�ڸ=
�>L=��{;�pZ`�b�M�x{Ҿ+o�>
��>9a�>��s>u�+�m�@�C�~=	�ྪ�4�2��>~e������4�W0r��%�����Ǹh�{ꃺ#E?����>�=�q}?�I?��?��>�L��_iؾ^�6>̀�U`=A��уg�Ԝ���?�o$?08�>�f��DD�i���i�>�?�/��`N�����g�Dw�)�)E)?[n��� �S�j��J��E����Mz�[����>��]?���?��E?��2li��0�jE=6+#>TF?�?�P5?z�l>|�n�3ᴾ�|Y��,>���?i��?G9�?
/-<��=����`��>�	?m��?T��?4�s?
:;��'�>�7;�'">ꠖ����=��>P7�=�?�=��?7 
?�p
?w��(�	�R��#��^�V��<@��=8��>�[�>��p>V��=�jg=4?�=�E\>��>̬�>7�c>O2�>4�>7������?\�>��=��%?��>��;<�����ݽ�-潛�����-���S�0KE�j*=�j�<�,d<W�=�*�>��Ŀ��?>0�6��D??�J徿nھ��>H��>�\y�4�?���<�?F>.�>=}v>�<:8>�y>�EӾP�>]���c!��,C���R���Ѿ�}z>ќ���&�ݟ�4y���@I�No��eg�Fj�.���;=��ڽ<�G�?������k���)�L�����?�[�>6?*ٌ������>W��>�ɍ>�J��[���rȍ�h���?���?/�c>~��>J�W?�3?ð/��2��Z�	�u�ҍ@�id�2a����S�����
�V�Ľf�_?�y?z�A?��}<d�z>7T�?ǧ%��펾JR�>��.���:�{G?=��>�в�~Xb�Ծw�þH��F>��o?�=�?$?Y�I>�}�=�2�>m�?�a?ىN?�8?�<�>�&�>�۽��I?���>A�=? �?�`?�X=��=�����T>���>�Y��΍��x�����ޏ<N�=�=E<�If=�3ƽu��V���3EE=ޝ=��e�}� =�nu=6��=�Q�=�|�>!�a?�?��A>�hJ?�0��e�;dʾ�v'?���;ը�����a����#�K��m.p?���?s�|?�%ǽ8��Tc�o>�x�>�v�<�0>��>-=�o��1�'���`>�u>G4�=BW��������3d��0���>���>�0|>����'>t{��P0z��d>��Q�]˺���S�g�G���1���v�eY�>��K?��?H��=_龃,��If�/)?k]<?hNM?��?�
�=�۾��9���J��=�G�>�c�<���y���m#����:�Q�:�s>�0��L͠��gb>��!E޾�n��J����5�M=A���V=%��վ�L�y�=�
>������ ����%˪��-J?�/j=L^��vU�ǅ���>��>�Ѯ>��8�@�v�"�@��y�����=���>M;>�A����'oG��6��K�>AB?�9Z?G�?j���3r�179���"&���c�-i?l�>���>9.>���=y׾�B�Е\�c�=���>o��>���KvI�K������ ,�߇�>��?%n0>N�?�_?�?�6V?��$?vb?W��>���f㽾B&?3��?��=�Խ4�T�� 9�JF����>z�)?��B�ѹ�>_�?ڽ?��&?��Q?̵?&�>� ��C@����>�Y�>��W��b��u�_>��J?���>�=Y?�ԃ?�=>T�5��颾�թ�W�=�>��2?�5#?8�?���>�~�>������ƾMo�>׍�?
?r�{?gQ���>��:��%J?�=��>l?���>h0?�M?�?ˋ>X��<���ʡ��⻽�f߽i��; *=t3>|�:O�F��/��;�<���<�؃=3;>���=��ݽM�6<��潤_�>��s>{
��{�0>;�ľ�O����@> ���IP��pڊ��:�H޷=ↀ>��?���>�Y#�q��=��>MI�>/���6(?��?�?5�!;ơb�L�ھ�K�3�>'	B?~��=��l�~���s�u��g=��m?~�^?�W��&��c�k?/�]?jf߾��[���Ͼ=����� �/��?��
?�w����>�?\/\?B��>V�>�h��妿��O��V��n�k=��>�������>ªF? ��>%0�>��={�!�E�}��跾pC?$e�?���?���?M
�<8䈿N�ֿ��~���&�m?/?�F��h�#?�W�=�:�]t�� _�<�������9��Ę��`�}eԽ��d�k�`�"0l>A0?��?J�?��\?�Q���r���V�&�N���i�EDվ�Ϋ[��A^��7j��ɇ��*���ﾬ�����h=q:��;�E�-$�?<(?��:��A�>m���Y�n�ɾ�Q>!������k��=	=��QU=�.s=K f�w'(��`����"?t��>��>w�=?1)]�D\<�o/�<l5��X����D>��>|�>ӫ�>X�����2�Z��!�ƾ����ӽ47v>gwc?f�K?l�n?�z�.1�炂���!��U0��a���B>\b>,��>�W����C&�&Y>�t�r�����s��{�	���~=x�2?��>M��>M�?� ?Oq	��m���vx�k�1�!!�<X)�>�!i?�6�>)ۆ>��Ͻ�� �6��>Y�j?1��>�3�>�2���0���l��`�$�x>j.�>�[�>�S>Ě`��[��o��]���o]-�\+�=�Z`?�E���m��Ԍ>��I?�O�!:Y=���>������c������� >�Q?̒�=��c>�>꾆�5\v���h�� )?�?�ϑ�5c*���>�^"?#�>��>��?pq�>¾��:��?!�^?2+J? �@?ʤ�>\�=�϶���ʽ��%��1=�͇>Z>�Vn=k��=؜�LZ��� �?N=U�=��̼�Գ�"�<�|��KC<��<��5>2mۿvCK�
�پ�
����>
�+爾U���wc������a������Ux��� �&��V�7c�s����l�Ǉ�?T=�?Q��//��3�������7���Q��>��q��u�F���9��L(���ྻ���xd!�x�O�G&i��e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@vA?��(����D�V=9��>ޔ	?S@>��1��D���@��>53�?���?�BN=��W�ۖ	�V{e?<<��F�^aܻ��=�Ť=�=���|J>�>�>ǉ��EA�t�۽P�4>Y�>"�!�Hc�^P^�0��<�c]><�սrv��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�����ǿf"�cm�	�`<�s(<��:�8��G���AwE�&7���d��)ǽ���=��>F�f>���>;�W> u>��Z?t�^?M��>��)>�q�P�����ľ��&v��3��Jy���t�.��v��z��0����e��k@��!=��=7R�l���G� �l�b�X�F���.?w$>Q�ʾ��M�H�-<�pʾk���T܄�L᥽�-̾�1�!"n�j͟?��A?�����V�L��AW�Ԅ��b�W?P�ۻ��ꬾ/��=f���)�=%�>&��=���� 3��~S���.?Y�?�+���<���C>�p߽+�<�0?p�?A�G<N��>��(?���e�߽f�i>��->>q�>=/�>=�=�󳾞2轱�'?��S?��������w�>$a̾t�{���=\m>��.�$�p�r>��<�/��ʺ<̜N���#=�W?ֳ�>5�)����aX��A� ��:==��x?^D?|=�>,bk?��B?�,�<fz��B�S��8���w=��W?i?�x>ܾ��(�Ͼ@e��n�5?��e?�EO>��g������.��;��?��n?�c?�*��$�}�M%�����Sn6?�sv?��\�>ʟ�T����W�尥>���>�/�>N8�b}�>��<?�{+�����Wÿ�(5����??�@���?��<9! ���=)�?� �>��M���ž����K˴�K�v=�h�>:��h�t��E ���*�?n7?"��?w?t��<
���=̢����? ��?�{Ѿ$�¼�
���f�o��;�=X��<�1���o0�l ��;�/оl�
������y=%ט>mQ@������>$k�n��?/ҿ�Ft�/yӾ?���� ?o>H<��񮿾hI���|���L��TI�<�V��M�>��>.�������_�{��q;��$���>��	�>��S�n&��l����Y5<�>���>¶�>E)���潾ř?'c��c?οA���ܝ�X�X?Zg�?�n�?�q?��9<��v�݋{�Sr��-G?N�s?-Z?1q%��;]���7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�d�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*��+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?)*�>Ĥ�?�b�=J��>h��="����A,���*>f`�=��.�� ?PN?:��>H��=�0��.�U[D��\R��P
�igC�c�>�Pc?"L?E�Y>����­����"��!ͽ�+�[^��|-A�f!"��Ž�E5>69>0�>�?@��w̾��?h�|�ؿ�i��c�'�-4?���>��?�����t�c���)_?Eg�>�<��+��y"���C����?TE�?��?)�׾ Y̼b�>���>=a�>y,ս�����w��{�7>n�B?^-��C����o���>���?��@�خ?�i��
?�#Ͼ��z��0���H�bA����#�?����<�>e6�>7�۽���3>���%{�|,�>�7�?�}�?^�>�Y?ZKM�Ou/���3��W�>9hz?}��>��;��ƾ�d>\��>Q��(��S���.�T?��@�r@�n?fo����п�癿�宾�P��\��=�E�=Jo:>�Z�^n�=�=>=}Q�<���l�>c��>�!�>�s>V�<>%�K>9IB>{���$�m���돿�H��3����8w�J��V�p����!ֵ�P�¾T���6���M��vsU���xv�<�*>n�O?ίd?�.?�f?<a�=$)V>�M��R��=F���Y'�<���>�[2?t�L?3�1?~�#=�Ӏ��d�����﻾��]����>_�>��>��>�1�>_�>�%�i>�
�=�r�>�*	=�G=`�;>.�v=y�[>ܝ�>��>���>I<>,�>�δ��2��[�h�4w��̽�?�����J��1��Y5��M���Lr�=1c.?�|>���S?п����40H?O����)�w�+���>��0?>bW?��>G��[�T�.>\��:�j�IY>' �Twl�(�)��Q>�j?gg>�u>�T3� �8�>P������{>�_6?\i��� 9���u�F H�.�ܾ��L>��>ߒD��@��񖿜?�8�i�N�y=��:?C�?N�������/t�Zޞ�,�Q>�0]>V=L�=U�M>�N_�O_ƽ��H��32=[&�=4_>p ?ZE->��=8�>�ʚ���S�R��>5 D>U%>}??�[$?3y��ʜ�L]���~.��)o>u��>s�>�>��I�f۫=��>��`>V�E�z������?�][>|���X�`��l�'܁=�c��os�=j�=,.�#x<�F�%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>ux��Z�������u�?�#=K��>�8H?�V����O�i>��v
?�?�^�੤���ȿ5|v����>W�?���?d�m��A���@����>;��?�gY?poi>�g۾6`Z����>л@?�R?
�>�9�u�'���?�޶?ӯ�?EI>�k�?�Xs?��>tW~�(u/��۳�K���w=�E@;,|�>��>�����F�-���i���U�j�Ӝ�1�a>�(=zs�>&3�Ej�����=�����ި�� g�`�>�@q>m�H>�q�>Y� ?N��>�>�;=E���Ic���ٖ�s�H?�,�?��������b>֘>[���L?��%?%����Z�>-aB?B�R?˃^?�5�>ٟ*��{��sCſ2rھ+<x��G�>"��>��?�h=�N>��G���)�>��M>��q�Xm���E�� '��r>�tD?���>�6�=��$?f�?��t>�ʽ>�AM�ˏ�x?9����>�S�>5,?(�U?e "?�D��D�=�dޅ��ט\��JN>�Y?�5$?ol�>U����Ѧ�
��<�^���m��[�?�w?��t�T?E�?�@D?�R??{F>�-ʼ��׾�E�&�>�!?��� B��%������?O�?&��>W̒��ٽs˾�����n��<4?<�[?�L&?	S�t�`��þ�@�<� ��Y%����;j&M��>U>�z��O��=J�>M�=1�m��C6�{Af<Nɾ=l��>�a�=��6�������+?uo⺉H���_�=�q�DKG�.�m>�E>&���W_?�K�k�z��H��1�����a���?93�?�:�?U����f�z{:?���?v?mK�>�H��@�ξ�־�I����u���
��>�A�>r��5
ݾ(񥿶�������K����5 ?ƴ>��?3��>.K=$$�>F�N���J�$m޾.����O� �T;�%E%�� H������q"�6�<Nz��������>ќ���<>�?l�P>��D>�� ?=���j~3>�s�>�7�>�!�>���>>��=u�5�=�U<S���KR?����B�'�w��R���h3B?�qd?#1�>di�@������z�?���?Ls�?)=v>�~h��,+�Nn?D>�>?��9q
?�S:= ;�=�<�U��8���2������>�E׽� :��M�+nf�{j
?�/?����̾(<׽�����	=�Ȉ?�?>?l�>��n��g���I�v�\�,>0=n��yǾ��-���w�;I������q��PA$�~�b>4.?^�?.�.�.���j���{��-h���i>%�?�`>$h�>�44=J#�p�-��m�i������>�u?|��>�oH?`D?T(=?a�K?�o�>�>W����2�>*�v<�7�>���>z79?R�1?ߕ2?�^?h"?F$>�6#�#D ��ʾJ�?F0?z�?&��>�R	?����
z� ��v��=�^���ZH�Nw�=�e= [��r�q�dGP=�1�>�2?_b��U9��&��[n>�7?�X�>R��>4��9K��d�=���>"�
?T�>������q����aN�>�6�?m����<��'>�%�=
���źk��={����%�=��v�Rk8���)<n��=a��=�ۤ:�4U:ݦ�;���<m�?a�#?��9>���>����&�x�&�O�<�(>p �>A?��*]��.����H��B�s�f��>���?��?�U�A�=��=���M����Ⱦ�6����>Z�?T >V1?���?c�]?�?L15>r����𠿢����^���.?� ,?/��>w����ʾ&񨿐�3���?�[?�=a�6���;)�0�¾nս�>�Z/��1~�8��WD�㲅�����������?���?�>A�Z�6��w�Q����T����C?��>�Z�>��>��)���g�%��);>��>�
R?�#�>z�O?�<{?��[?9hT>&�8�K1���ә�:>3���!>@?��?��?{y?�t�>W�>�)�
ྯT��c����ႾcW="	Z>V��>
)�>��>���=Ƚ?X��1�>��`�=��b>=��>���>��>��w>wS�<M`E?���>{��GD�����c�r��mB�-`?���?��.?�3��2�o�W����v�>�z�?��?7^J?��y��-�=�c��৾��.��Ƴ>��>�`�>1�=w%�=���=���>�/�>G�N�`���21����<d�)?�W5?���ƿ'�q���p�����8e<�V�d����[�I�=����B���©�K�[�ۨ���{���`����{���>-4�=^��=#�=�F�<�kɼ��<��J="-�<f�=�Hp�Eo<"U8���ѻ}Ĉ����`�\<��I=���}˾��}?�6I?1�+?�C?��y>�[>y�3����>����=@?�"V>�9P�xr��8r;�§�����O�ؾ�u׾��c��ǟ��/>xI���>b(3>�r�=E�<��=�r=��=˒R��=�L�=�A�=q��=��=��>�b>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�7>�> �R��1�Gy\���b��[Z��!?�F;�_R̾�?�>^�=m!߾�ƾ�d.=�w6>�yb=�l�=P\�@�=�{��;=��k=Qˉ>}�C>ue�=�9��q��=	�I=��==�O>ǔ�0�7��
,���3=���=z�b>m�%>s��>r�?�a0?�Xd?6�>n��Ͼ[?��I�>S�=�E�>���=<rB>���>I�7?8�D?��K?��>���=�	�>��>;�,��m�}m�Y̧�֎�<���?�Ά?>Ҹ>7�Q<�A�̠��g>�//Ž�v?7S1?�k?b�>�3���߿t�#����f!����<��=x��������[�X����=���>���>B�>2�>��[>nŘ>v �>= ==��=�d����<~��ɋ���~�iw�=�.��|J�=�qW��Ƚ���3�<]V��.D<~WH<�{>���>��=��>Zu{={=��>< ��#�f��
>h�����:���k���~�#�2�O q��d>[�P>X�\��s���W�>�W>��M>@�?hj?��r>!�K�Q2��d1��X?���>�8~#>S�:>���=S�K'p��Q�R���Y��>k�>P��>��l>,�-?��$x=��ᾮw5�<�>G����'��]�O8q�o8������Ci��Ӻ\�D?!=��H�=,~?5�I?{Ώ?j��>�
��u�ؾq�0>U��=#����p����
?H�&?�a�>[�c�D�\Օ�����ȝ>]�6�ִZ�j	���N�Y�j��1��v�>h����z�c�?�.����?��mn=�[������>��o?�͠?��v�ʉ��l�w�Aj���J>zɅ>��F?�U�>" ?��>�U[��������A>�
v?�c�?��?O�+�l��=�U��:��>>,
?8z�?Ր?=Ou?�)^�L>�>e.6�2�N>�h��Qt�=��>��d=��=��?
?Z�?nUz�F�	�!����gUZ�'�W<�j�=u�>�%w>{�q>6�=�٘=(��=��\>D#�>���>�V_>%�>��y>������2�}f?,�>��%>-?VA�>��M�T�t��=A\�����!ٌ���b��ƅ��\>����8"�=q�=0�?"Ŀ��?��>+�'��?:���--��<[>�>�>����>d�>�8�=u�~>�k>_�>�Қ>JvT>,FӾ�>���*d!��,C�i�R���Ѿ�}z>q����	&����w��CI�o��Bg�j�M.��<=��ν<H�?x�����k��)�����\�?�Z�>�6?�،�|
��4�>���><ȍ>�J�����ȍ�hᾁ�?���?��e>���>�ZV?O�?[H4��C3��I\�6�t�[?���a��z`����Y���_'�pUϽ�/_?��x?��C?_~�<��x>Z(�?h�$�-����>Ld,�D�:��==�>f;���e�	#Ӿ^�ž�
�FAE>;p?�:�?�$?�Ud��)H���\>�_+?:H?Ǖw?\�H?�Y?�z�:�D?��<�ـ6?,��>5FD?FN?/�?�8�>9�	>_��>=<��B���@/E���0<��=o�7=�˱=�?轎d�À`��x�=��O�~����`�S����<A��=���=R{->��>��\?\��>?VL>�(?k��v(L�����	4?:�=Ɏ��������Ѿ�	���=@�q?�"�?C�n?a�>%�?�+0K�'	>dͫ>�2
>�B>�Ϳ>rZ���@��t=�=GY>-5=�!&���u�d���W�k�� �=��>}0|>���d�'>a|���0z�'�d>��Q�l̺���S���G���1���v��Y�>;�K?��?���=x_��-��rIf�)0)?�]<?�NM?��?��=��۾��9���J�>���>�X�<��������#����:�8h�:��s>�1���s����e>'x��ݾK�n��VJ�����==Ǐ�m�W=���'�Ӿ�~��w�=��>�nľ�� �ޖ��ߪ�эI?�`h=�Ӥ�]^��e��Z>�ǖ>�>o�<�zY���?�������=�N�>�=>���M��ZKF�N��P�>�=E?b-^?�'�?_؃�g s�v�B�����y���W¼x�?��>3�?}><>8æ=xW�������d���G����>���>#=�CI��D����s�$����>��?I>|�?wsR?��
?V0a?L"*?0�?���>�s���>���A&?��?��=��Խ��T�� 9��F�� �>��)?��B����>P�?Ƽ?K�&?)�Q?ŵ?��>"� �~C@�蔕>@Y�>��W��b��.�_>��J?c��>�=Y?�ԃ?��=>��5��ꢾ�ѩ��Z�=�>�2?�6#?�?}��>�>[�����=�I�>��L?)'�?Z�j?~��<y�>�1=s?�[C=�:�>��?�~?~j)?�IR?b8M?A��>�-���	��S��g�<�Z�<�Ӏ=E=?ⶽĐ��|&�1
=^�
<s�н=������u���� ��8�<�^�>R�s>����1>Ͻľ=7���@>�ۤ�XK���):���=y��>�?_��>�j#�cy�=P��>�<�>.��r7(?��?�?F@	;ʗb�<�ھ�K���>B?Q��=��l�eo��V�u�%�h=��m?7}^?#�W��U���Z?d�d?����w��@¾�x��(�;�a?��U>Hr��ҍP>u?*G?�,�>/JR��(���C���f�0ᾙ\�=�y�>|s��L��<9?�D?�H�>�w�><��<����@�k�F���>�&�?A��?��?*��<��t���ɿ����l��ޗ[?Ee�>`|���?�!��/�پן��^�\=����u�$pe�]dx��Fb��A��X����߽��>k�(?L�r?���?�tL?"�"z��GH��Lv�h�W��K/�o�w��u_�B'U�R��D6����m���D<�}�j�A��?Z�'?�]/��h�>�㖾��R�̾��?>eɝ��F���=�ˇ��<==�R=��g�4]-��⫾	] ?5<�>��>��<?/[�>�=�?d1�"7��H��pP2>Sՠ>���>q��>�H��Y�.�l�q�ɾU̅�8(ѽ�:v>�{c?�zK?��n?r���51����c�!���0�=��DXB>�|>쯉>�0X����J&��L>���r�;��r��7�	��9=܌2?6�>�Ҝ>,@�?$?Zf	�����Ox�'q1��Q�<M�>i?��>V��>r�Ͻ{� �%��>�To?
��>Bܾ>Tt��281�{�t�9i$���>T�>X��>��h>QE��'p�t���������)�/چ=l�_?�p���V���>&�D?W��;�{�<�Ù>>y����ޢ��a]��>5a?T�7=�>0>��������⯾�#&?�(�>�:��uO%�B�>,K.?y;�>�ȃ>[3~?�C�>����}.7=�:?O�a?��G?��7?D��>)��;q���η�T���=��>�H�>���=�b�=�)��b������=�Q�=�#<Q'o��<;�<��<�=�N>peۿ�K���پ@���:�
��㈾�G��=��?v�Y��8����[w�g$�e�"��V���b��|���k�A��?5��?W*���[ٚ�S���Y������>��p�5�v��������@��	��ꬾOa!�z�O�Wi�k�e�P�'?�����ǿ򰡿�:ܾ4! ?�A ?8�y?��7�"���8�� >UC�<-����뾭����οC�����^?���>��/��r��>ޥ�>�X>�Hq>����螾�1�<��?6�-?��>Ŏr�0�ɿb����¤<���?0�@�OA?u�(�N��E�W=�P�>1�	?P@>f 2�r�<J��\�>��?gߊ?�rS=D'W���
��d?�E�;�F��
޻'f�=�Ф='�=�����I>O�>���:�@�7ٽI5>��>?i�.m��e]����<�]>��ս�+��5Մ?,{\��f���/��T��U>��T?�*�>U:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=x6�����{���&V�~��=[��>b�>,������O��I��U��=t���ǿF����ԑ<�=!=����#��ͽ�v���o��[^-��u���=1�K>��G>1D�>M&W>��>��g?�A?e��>��>]���4���P�@G=�8(��<=GѾ
ĽEI���&�C�ܾ����o���b4���7:��۠=�P�ُ��"��b���G��,?��>�hʾ�SN�Oы<�0Ⱦۮ��"W�1b׽�оow1�ԙo����?��??^����[�FH�g*���f��ai[?M����j�����=� ¼�Ba=L@�>G��=�S�1���Q���.?3J?���~���t/C>�O��<��*?��>���<j�>��%?��&��q ��\e>xf(>��>6Z�>vO�=򥲾v��}@'?j�Y?m��ѡ��w��>|vž�l���Y�=�>�%�b�t;�ec>\�m<Yj����<�E�Y��=S%W?�>�)����i��S?���<=b�x?f�?�&�>pk?��B?��<�q����S�r*�$�v=\�W?^i?1�>Ћ��Iо!�����5?%�e?�N>8+h����e�.��L�}$?�n?�e?�����r}����C���i6?[�v?�I^��}��G��>W�4�>?x�>���>ު9��j�>Bk>?F�#�IJ������9V4��Ҟ?��@��?�
7<^^�0.�=j3?p��>P}O��UƾI��D����pp=���>'8��$1v�c��B�,�~p8?��?�R�>�u��r��Ƿ=���AT�?��?+>־.ɿ�����-s�x��M�/>����]��!��7cﾣEC���о��R]���=��>�V@G���A�>��.�����bͿ�}�:ھ�{���#?�:>'܌���ھ���ދn���D�6}%��#��	f�>��H>�W��m��Ѓ�v�N��g��'?��>q��>�+����	��������>���>�F�>A�=�����x�?��澒ɿ�����C�h�c?���?<��?�b/?�y=���E���/{>��V?a;x?
�u?c�O>��A�N�+�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�f�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ���
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>�^�?\�=/��>i� >
���8G��4>S��= #��,A�>v�M?+�>ZK�=7� �(��D�X�V����UA��lz>�Zm?��S?L�b>�����)�<t�#��������| 	���%���4<e���e�'>a�&> �<>@� �������?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�	??��DɆ�H�{�=u�ˊC��Y�=5�9?=뾡�y>���>Sא=�Iy������t�q��>)ί?��?y+�>�Ml?�&m�^C���=��>�k?��
?CHa<��@E>>y�?+�5���G���cg??�
@��@~j^?W9��+߿�A���8{�-�¾�v�=��>Ǟz>m@ӽ�F>{��;��><i��<3qA> ��>I��>\�>�b>�3>�_�>� ��p�"����u��mN<��u�	���Vs��0�s�\��'�VZԾ��ž��ӽ<�<7�b;?���}�=p��=�.R?�W?��B?H�?�����>�Ͼ	TԽU{��i�/=wL�>��,?/?} ?��8����r�4	g����R��	?�/�>�$�>,?Z4�>A���>h�=�6�>�ݽ���= V�>tU���k>2Ǩ>���>�?dD>t5(>�������G"c�gqu���߽x��?E�����J�����B��|��l��=�.?D��=k����hпiG��R(E?���';�$�%�a�>@i/?��V?6�>sܦ��2�`�>�~��	l��Y>X�޽��M�3&$���@>�?��o>@�>�43��;���F�����n>�<6?s贾-�6���r�j�?��۾��;>"#�>*�o����z��yi��*in���M=f.??�	?7���YǮ�VZ��֣��J>Rm>�%+=�M�=a
Z>�d[�W^˽�dD�H��=2�>��u>��?��&>��=jΣ>x떾��J���>�|<>*�)>\;=?s)&?�q
�7��˗�18(���r>�h�>��}>
�>�CI����=e�>Q X>�!�7�����Q>���W>��i�+�^���m���=&s��2��=��=�S ��i>��_�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾXh�>Jv�LZ��s����u�x�#=���>o8H?�V����O��>�w
?�?�_�ש����ȿQ|v����>��?z��?��m�XA���@����><��?�fY?{si>lh۾ScZ�S��>��@?IR?��>�8���'�;�?�޶?���?�R>q�?��E?���>�,�L�,u���C���;��n��=��m=�e>֪�v�c���oŒ��I���'��N=�P�<�ٖ>��?�������_��l�=8o��{ =8�>�j�=�*>#^�>��?�d�>I8�>��#�C/��Z�>�S���t2H?zS�?̤!�����S�>4�8=�.����?��?�⛽��ھϝ�>�"0?5�L?1�X?�c>#�+�,Q����ȿ3i����O���>2?�?�>�Д��O�>�{� T.��֭>��>��-��㩾��i�a�:��>uS8?Y��>�F>�;?I!(?��S>�(�>OK��@����K����>���>��	?v�d?q??I��X�>�ᓿ����<l]�R$>��Y?��?���>���NӦ��5t�Gc=�}ƽHʊ?��P?�N��?���?�:4?͠P?�ϊ>T�%�(D��ℽo�m>��?�(�c�@��)��6��$?
?
��>�m��O�}=���|Ծ͹?��Z?�6?OF��X���ž�^�<Ȯ=�C��M#��V���>~�>�0v�@��=��K>C�=�<N�ᆺ�-�m='t�=���>���=3�:�`R"��:?�O\>���w>�|p�܅g��Z>Hւ>�ZK��GR?��anu�"���L������o�?q��?�`�?}B��ASZ�K�$?|��?�s&?MQ�>�s�����}P�\4���8�U��>��>��žn�U���b��������=Ԫ����>N�>;%?|�>�jI>��>ͬ���(�+*�d��\��o�o29��|/��5�QE��w�&�r	��&��H�z��٘>l����>�R
?bd>�jw>H��>~@��M�>��T>�>��>+aV>��,>\b�=��;�3�`�Q?����b�'�gn��ܬ�R�A?K�c?=��>�gk��Z������?���?��?R�y>/�g���*��?���>�~�d�
?�K0=xћ��,�;u����������	��W�>��ֽ�+9���I��_���
?�?Ѹ���n̾d��	 ���)=l�?Н5?�/@�d__�!$z��u\���Y�N`�=(e����Ӿ��7���q�$��RL������G�	��>ǩ(?���?��BȾ$7M��~�c�;�>*��>��=i+�>�4>��8��cC�9�f�����3���?g�U?�'�>-�I?��=?yN?yM?�z�>k�>�̫�J��>�D:<.��>�k�>��8?��-?��.?Hj?W(?2�O>9������Ӿ�?&�?X�?l?u�?n������ޗ���Ր��JՈ�G��=�H�<������h�pr=��g>�-?�)��8��[��>D�<?��>��>s6��pU��4>���>�?x��>AѾRX_�tz	����>��g?�.�Zx=�+>�}=`��
��;r��=��'�V+�= m:=ޜּCά<��>`�=���:Q��<�x;;��;
��<�y�>��?6��>@D�>jE��>� �����z�=�Y>yS>1>aNپ�~��$����g�Lxy>�y�?b{�?h�f=�=���=Fv��fI��n��������<g�?PC#?�TT?啒?3�=?�e#?-�>�*�~M���^��+��A�?� ,?j��>���/�ʾ�쨿�3��?�[?�9a����:)��¾	�Խ}�>_V/��+~�=��ZD�xA�����M���L��?���?F	A�@�6��j�����"]��G�C?� �>�W�>5�>N�)���g��#�A;>Ռ�>uR?`#�>��O?f1{?�[?�yT>h�8�U*��љ�Nt3���!>�@?���?��? y?�w�>��>+�)���N���������ނ�^yV=��Y>���>� �>e�>u��= �ǽmS����>�鐥=��b>��>���>I��>�ww>�8�<��Z?���>���d��(���|ž6ܽ�k�?ɓ�?�(?�䌾Q\r�=ZT�>��x>�ݾ?|��?��]?*v��TN>��F=O���н:��>���>�]3?h;%���@;x#�=Eh�>�v�>��޽����2 ��H��=��>��"?�|
=K�Ŀ�Rq��hm�U��&0�<����j�]�����7]��j�=K%�����,q����W����=-������|��V0v��>�'�=v3�=o��=O/�<�+�U�<riG=Ҍ�<�:=?nf�9Ք<^:��G"�dށ�K��^'<�5=�类F�ʾAV}?�J?�E+?`�C?C�{>6>�g(�{e�>+ ����?XS>�3G�O���`9����Ԕ�y�پDdԾ�d�Lb���>��A��>:63>4��=l�<]��=�L=w�=�~��Js=���=�ػ=m�=v�=`�>�>�6w?S���	����4Q��Z罙�:?�8�>�{�=k�ƾp@?I�>>�2������xb��-?���?�T�?F�?Kti��d�>K���㎽�q�=;����=2>���=��2�S��>��J>���K�������4�?��@��??�ዿ̢Ͽa/>|=>�3
>�)S��-5���P��]�w�Z�T�!?6�:�o;�J�>7A�=�cܾ�þ<iZ=��/>Z:=1X)���^�8�=���:=$��=}�>qEF>k�=랺�>�=�(k=�u�=CP>4 �Y�+�e��%Nj='<�=�\>[�!>���>��?�Z0?�Sd?�@�>6�m�
Ͼ�=���D�>��=�Q�>�م=�tB>u��>��7?�D?��K?�s�>Bĉ=���>��>Ô,���m�_~��Ƨ�	��<0��?͆?�̸>R<�A�����W>�'�Ľv?CL1?f?2Ϟ>.���ٿP5 ���A��dG=���=[����K	�`/
���@������7>�>W��>H��>\o>�@9>��>�!�>��
>><�x[�=#r�����i��>?��<�k�=*��=���<"�/=N�"��4̜�	V��-��h9����>P-�>4X�="��>`=^Ծ��>
f��{X�x$>:����8���d����n(7���I��#P>�3>�0�h���OR�>�l>U_9>x��?��k?�f>]O�7t� ���P���75�`�$>�P�=��:���F�^�`��\��v�%��>v��>�-�>Go>��+�3�?�5$t=��y6����>�W��������q��J��Jݟ�soh��A[�I\D?�&���#�=��}?�9I?��?̅�>Ԙ�.wپ�/>,?��5�=N���lm�Eo��i�?�&?�Z�>(�
;E��i��)ͺ����>������e�`l��6�g�ˤ=�陾���>�!��(q ���a�;������8�\��7�>�*K?���?�&��`��:�R�M6���X��˺�><��?���>��>,��>�/��$ ���h��I>5��?��?��?�i#��O�=-T�x��>ӄ#?��?�?��f?�%o���>�v�ܓ�>�6<q7�=�Z>��=h��<{��>�<�>�?�:�����	�:��6�O�����ډ7�n�[>Li|>/�>">f�0<�$#=e�^>�k�>'�]>9'1>�b�>��">Ҿ��%�od?M�	>Q�W>O/?նi>�KT<1ܛ���=�@��(ս������U���μ�D�;���zlc=���=M�?��ſ-��? ;^>�*��G?�s�@�ػ�3h>i�>g����>A >�gO>���>~�|>��=�X>�>47Ӿ^�>���a!��1C��R��Ѿ�^z>N���&�Υ��6��9I�����Go��j�%.���;=�%Ȼ<�D�?�����k���)������?�H�>&)6?h猾O�����>m��>U��>�������ō������?���?Q<d>��>�dW?%�?DQ9��{<��M]�L�r�Y&?��c��`�*������y��s�ӽ]�^?�8x??�B?��<*}>Wb�?07&��z���#�>7�-�Z�:�CQs=��>���ڮh��վ�z¾���'BM>;q?*}�?�?V�]����q`�=�;?^��>�0[?܀M?�.7?�f7�}S	?�G�dT;?`r�>iC??]I?��?�W>.�d���ř�=�`/��p��������g=�z&;���=q"�<���L䉼W�� T�=&t�=���<bʔ<Y��<��<Yz=�H�>-�>�>b�]?PJ�>	��>��7?���v8��Ů��*/?h�9=ۭ��k��hʢ�$�K�>�j?' �?dZ?Had>v�A�TC��>ZZ�>�r&>�\>�d�>�ｃ�E��݇=�M>�\>ť=�rM��ρ�L�	�w�����<&>R��>x/|>E��T�'>�z���.z���d>�Q��̺��S�`�G���1�Z�v��X�>;�K?��?���=�^��-���Hf�|/)?�]<?OM?T�?��=��۾e�9���J�$?���>�t�<]�������#����:�!�:'�s>E0������rVb>����/޾�wn�,J�l���DL=̛��U=L8��8־�	��=�
>�*��^� �i��HЪ�� J?V�h=�{���9U��`��>���>�j�>y�<�q�u��h@�O�����=���>�a;>�6����?�G�+��<�>PE?�W_?lj�? ��k	s�M�B�:���9^���&ȼ!�?�w�>bi?�B>��=䝱�'�/�d�G���>��>�����G��;��^,��R�$����>�9?��>��? �R?I�
?�`?*?.D?�$�>������B&?)��?��=��Խ�T�� 9�,F�4��>K�)?��B����>,�?ӽ?�&? �Q?��?��>�� ��C@�Ĕ�>]Y�>��W�pb���_>��J?	��>b=Y?�ԃ?��=><�5��颾ש��T�=G>b�2?6#?[�?���>���>�f�����=
u�>��b?�,�?��o?2@�=�?G�1>���>�}�=���>q�>�?�/O?[�s?��J?	��>(�<ﭽUQ����s�F.Q��N~;/�E<V{x=��ݍt�� �`W�<�k�;����}�S�;E�xE���o�;���>5�>� Ǿx�>Zô�����<>ߡ���Ӿ�펾
�����<�6�>.*?��>�Ң:'�=�Ng>4��>���]6?��>��4?���!l�A��<� ��"�>�7f?k	>I�|������Pa�����ZQ?�x?Z-�0��o�i?��Y?�6�Ě\�! ���.��iҾU!n?�?Q��ɷ�>�?�?i?�*�>Ʋ� ����;uH���C��#=�v��>?C���I�X��>��?�̢>��=u&ʽ���p�t��Yھ���>8�?�ح?Ρ�?��<A�j�v���b���O�?r��>z�"�R"(?����9ľ=�ľ\j����ӷ������i����s���[ͽ��[�Xa)��?�=�=9?��?�A�?�4O?�'����+i���[���N�0ɨ�D6�9iq�m�y������b��N��8�̾-��ErW=����
B�ń�?ϴ'?�=1�d4�>���T��G;#$C>������|ȟ=�y��PjA=��\=h�g�A�-�t$��j� ?[n�>z��>Q�<?4\�$>�۰1�SG7�����5>�l�>:��>^��>��/�U�-�����ɾ����ӽ98v>0yc?��K?зn?te�\)1��̗!�d�/��a����B>�p>o��>n�W�0��;&�PY>�o�r�4���w��R�	�<�~=,�2?6*�>n��>�O�??�x	�dl���_x�r�1�⡃<W/�>�i?�?�>��>P�Ͻ�� �B��>Y�l?>p�>LĠ>my��G!��{��[ɽ�1�>W�>���>S�p>�Q,�y \� n������m*9��y�=4�h?
����b`���>��Q?m��:N	K<�^�>�fw���!�]�e?(���>�~?�Ū=��;>��žb.�A�{�bj��;O)?�K?�撾��*�z5~>�$"?���>f-�>/1�?F)�>nþ�C�ױ?A�^?�@J?(SA?�I�>��=�����=Ƚ��&�}�,=��>��Z>�m=�|�=����q\��x�H�D=iw�=(�μ�P����<Zw����J<��<��3>	mۿlCK�Z�پ�
���>
�q爾���Jd������a�����Vx�M��P�&��V�"6c�x�����l�܇�?%=�?�~��l/��b������R������>��q�ax�����X���)��͗�E���;d!���O�^&i��e�Q�'?�����ǿ밡��:ܾ'! ?�A ?%�y?��@�"���8�$� >lC�<�*����뾤����οN�����^?���>��/�����>Υ�>��X>	Iq>����螾�1�<��?6�-?��>��r�,�ɿc���Ĥ<���?.�@=}A?b�(����A2V=���>͎	?e�?>4W1��I������Q�>�;�?l��?	�M=��W�Z�	��e?�S<��F���ݻR�=�9�=�M=���L�J>�U�>���MA�E9ܽø4>ۅ>��"����^��Y�<'�]>��ս,?��.Մ?�z\��f�â/��T���Q>��T?a*�>_7�=��,?|7H�M}Ͽ��\�$+a?�0�?��?(�(?�ۿ��ؚ> �ܾ(�M?D6?C��>�d&���t�k��=�<ἂ���B��w&V�0��=ī�>��>N�,����ׅO��I�����=��?�ƿ��$�.c���=^X��h�Z���+��]V�����Uo����)<k=���=�Q>��>QW>�%Z>a|W?�k?
��>�>C��2t���ξ�����l���v�������pǣ�\5�Mv߾+^	���������ɾ%=�#�=�5R�㕐�̼ �w�b�5�F�K�.?�[$>_�ʾP�M��A+<�qʾ]Ī��������#̾&�1��&n��ʟ?
�A?������V����]0�����B�W?�l�Է��묾���=P����=5;�>-��=���V*3��wS�]p0?�e?Uz��"a��)x*>�� �֑=9�+?�?��[<G,�>�T%?E�*��{��-[>D3>u��>X��>Z�> �� ۽y�?��T?U���՜���>�[��lwz�e`=��>�e5�:��k�[>���<nጾ�S�� ���H�<�Nr?�go>RI��f%����#Q��t&�=�]�?0�0?L�?��c?�
r? F��
��}��}*�`c��z|A?�2�?��=k��=��������N?�/d?Fy=�L � ���T"�����F?t�?�?����Qo�������y��c?��v?s^�xs�����L�V�e=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?G�;<��V��=�;?k\�>��O��>ƾ�z������4�q=�"�>���~ev����R,�f�8?ݠ�?���>������AL�=����3��?��?O嬾��h<���B l��������<��=�c#�8�*�f���7�g_ƾ�~
��z��z0��=B�>�u@b����>�F8��x⿖5Ͽ�ׅ��jо}r�nR?���>�qҽ
���H�j�a}t�aG�]�G�����Wң>�>�ؕ�'��@y�:�;����`��>���`�>��\�$»����Ø;;W@�>X�>X��>�$�� ľ��?'"����ο)����X?�&�?1�?[?�s*<<<{�.u���;�[H?�Qu?�b[?s><��j��E�_�j?tY���U`���4�RDE��U>�3?�M�>P�-���|=#>���>�r>�#/�X�Ŀwڶ�����U��?���?�r����>H��?On+?�c��4��Z\����*�3�E�4A?��1>�����!� ,=��ǒ���
?�w0?�~��1���O?p�'�Q�g�S���%>u��=��2���Ҿ=K������`k��i��ꆇ����?'@�R�?>lξ
cZ���>^�>����5����>��z> �*>`K�>J���%��=(��
�}4�>�Q�? l�?x�?萈�렕��SD��ه?���>^�?Z�<�!4>�>ĵ����,���>���=& =��>��`?�ٓ>#�*�~f��6�G��t��g�nlA��C����>�pU?��Y?�X�>��<?7"��x��~ؼz���8>.�|�$.A�� ��d>�z}>�B�>i�=�{�����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�^��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�Q�B�{�1=:M�>Μk?�s?�Po���f�B>��?"������L��f?�
@u@`�^?*0�Ͽ_���C���+ž!w=[>փ4>��>����=(�@>�ď<�� �̨:>A�>�V)>0�Y>+e>jm>��>Z��� n �X���س���2Q��C�XB��������C����"��괾����U��Z� H��#�fѽM�ݼM�=/�U?��Q?H�o?� ?LOw�,�>c8���=�(#�,��=�]�>@O2?�fL?nm*?F�=-�����d�4V��?�������b�>R�I>��>���>�V�>i-8�fJ>0�>>���>�f >&�'=au��VO=��N>�k�>8��>Ny�>�V<>�>�˴�+����h�!w��ͽ��?������J��4��T�������b�=4t.?�>z���;п���J+H?���Y$���+���>ܽ0?SW?y3>�9��<�T�::>��3�j�ů>�����~l���)�8�P>�p?2�f>/u>d�3��e8��P�U���f'|>..6?����{B9���u���H�dݾ�NM>�ʾ>;mC��z�[�������i�F�{=�u:?��?g��7۰�?�u��T���7R>�.\>f�=���=�BM>C�b��ƽ� H�`�.=u�=۰^>AS?��+>���=��>\���9P����>�[B>�2,>�@?�&%?ƫ�v��"t����-�Fw>NK�>���>oI>@J�?ϯ=V�>v�a>�g�����-��/�?�c�W>s�|��R_��eu�~ux=�K�����=_!�=Vl �p�<�.%='�|?�q��ᕇ��(ݾ�j��`�7?d�>��<G�˼	*��'��E	��Z�?B�@Z�?�"���<Y��?���?Aq����=��>�w�>S�Ҿ����H?{H��܈���{�$����? �?w3�鐉��o���:>�+?�ż�eh�>cx��Z�������u���#=H��>�8H?�V����O�T>�w
?�?�^�ᩤ���ȿ9|v����>T�?���?P�m��A���@����>6��?�gY?Soi>�g۾s`Z����>ͻ@?�R?�>�9���'�q�?�޶?ɯ�?<I>���?�s?�k�>y.x�\Z/��6������Ar=�y[;-e�>X>����hgF��ד��h��Y�j����e�a>��$=#�>�E�4���9�=�����H����f�c��>n-q>��I>�V�>_� ?�a�>��>�x=�n��>ှ������K?���?���P?n�'�<}=�=ל^��F?�(4?L\Y���Ͼ�>�\?���?|�Z?e�>G�<��b쿿̦��͗<�%L>�T�>�?�>Y����K>sվ�SD��X�>�ח>�ͦ��Nھ���#����z�>�f!?�A�>P��=^� ?o�#?=yj>F&�>�dE�g8����E�!��>���>O?p�~?��?&߹��[3��	��:塿x�[��HN>��x?&U?Pȕ>���׆��Q�D�_�H�n	��U��?rg?-:彞?5�?�??h�A?�f>l��=ؾ٭�#��>��!?%��A�w@&����Z?C?���>O���Rֽe`ۼ���z���?�K\?(d&?ʭ�"Ea��þ���<�h$��?U��&<��C�3�>`�>۫��.-�=��>� �=�l��T6� �q<'��=�@�>l[�=Ik7�Ю��3=,?��G��ۃ�$�=��r�AxD���>�IL>	����^?xl=�	�{�����x��	U�� �? ��?[k�?���2�h��$=?�?<	?V"�>�J���}޾�྄Pw��}x�qw���>���>�l���I���ڙ���F����Ž����>���>�?|� ?��O>fU�>�!��J'��q񾊟�-�^��Y��l8�U�.�©�jԠ�yF#�Of�K7¾ �{�9�>� ����>A�
?�%h>@�{>�!�>7�Ȼ�i�>r�Q>L�>�i�>�X>�	5>_�>��<�wнMR?�����'����h����)B?fd?�;�>�$i�����u���?��?n�?�)v>u�h��7+�Ne?�5�>!���q
?al:=�����<�d������6���o���>�Z׽V%:��M�8\f�.m
?.1?���<�̾?�׽[���)n=)V�?�(?��)��Q��o���W�lS�����`h��z����$�֠p�鏿�Y��� ��Г(�+�*=�*?�%�?"��:��-��7k��?�[Zf>���>��>�Ѿ>�I>Q�	���1�{ ^��@'�穃�Fi�>!Q{?���>��I?I<?!oP?'kL?v̎>�q�>�!���r�>�:�;W�>j��>]�9?J�-?�&0?Wl?�n+?�3c>�I�� ���^�ؾ(?T�?�??k? �?	܅�`uýل����g��y�BV���@�=�o�<&�׽�u�=
U=�T>�D?�a� �8������k>�7?r��>w��>�؏��D����<�>��
?�2�>u ��sr��\�G�>ᜂ?� ���=��)>@��=�І�&�ߺaM�=����q�=,:��˲;�&�<A��=-��=,2t�$ʹ���:� �;�߭<�X?MP?���=��>�ĺ��	�
�ؾE D>�>̟�>UB6>���{�������4/\�.N>_��?�e�?Ϳ~=��5>�'�=1����#�C��K0��v�&�9?��E?/�K?�'�?��S?�o?�̬=�:X�O����O��Bѩ���8?�!,?��>���G�ʾE樿�3�w�?�G?�Aa�����B)�¾^�Խs>�?/��~���D�
�|�P���P�����?Hŝ?��A�i�6�90�A����4��q�C?��>�]�>c"�>E�)���g��-�}j;>ݞ�>�R?88�>��O?{?��[?�T>&�8�F5��t֙��<�.!>��??���?��?�7y?���>P@>!*��@�D����s���w߂���Z=��Y>z��>��>z�>��=l�ǽIh��X�>���=4bb>�^�>1A�>�A�>Jx>��<sO?Z��>����k�
(��x;5-=��N?CO�?��??��_��<��5X�����ؤ�>~��?��?��3?�����s>���3������7��>��>{H_>
&�>�%�>R;>�??kU�>�m��j�>�H3^��&c��?�(m?x�>i�ſ��q���p�����yAg<t��O�d�nO�Z�9�=.���9���x����Z�����`X�������`����{����><<�=B��=���=���<1aɼ�<�M=�ߊ<S�=R�r�/bl<�7�������J�D�]<dI=����M)|�0�g?h2?�A�>�7?�m�>|
�> �=�?k�m�G?b�d>0�A>"�Ǿ�ߘ�P�;�i��!׾0ӌ�	!-���?�a�C>^�=���<�>�rc>N��>�,�=,8�=Q���b�=)�>oB�<?�8>�Q>��1>z>�=�fi?P�V�c���[T?�G�R��L?�<�|>u#߾�A? Q��ڎ��C����Nnx?�X�?K�?�?��ھ��>�Φ��w�<�M=6�\>i�ܼ����j>�M>x���$��8�>�,�?V�@q�N?%
���-ۿ�X'>w�7>2>��R�1���\���b���Z���!?yG;�JD̾�4�>�!�=�*߾��ƾ�v.=L{6>�b=�|��X\��̙=��z�`<=�Gl=Zۉ>��C>�w�=�C��Y�=\�I=b��=޾O>,ȕ��7�x,���3=2��=[�b>@&>��>�?�~?�m?�ϸ>����i-ξ�1;�3d>�_�=�ߌ>�/�=J"<>0��>�EB?�E?'\D?.<�>���=T�>�ң>�
)��DU����p���=��?��?���>��<K	B�E���B��M�b]�>^�:?��?J�>�0	�6fֿ�J�.�>�U�z�&I�=� *=������+;#�e�P�+E��z>g�>�#�>��>���>��>�/�>���>N�p;k=9=l�>9<�=E�x<M���P���������m]��J�7ټ�G�=�M=U<�=C�r<��=��>��="��>n<>Ь�>q��=����C/>ϸ���L����=�G��[,B��4d��I~�N/��V6�l�B>;X>�}��?4����?X�Y>�l?>���?YAu?4�>� ���վ�Q���Ce�:VS�`˸=>�>u�<��z;��Z`�z�M�_|Ҿ���>��>���>��l>�,�p?���w=��ᾬZ5���>yy��k��h�8q�Z@�������i��aѺ	�D?F�����=�~?�I?��?q��>�&��,�ؾd0>�W���P=X��q�gS��?t
'?��>�쾭�D�XG̾?!��a�>�:I���O�����D�0�2��Ϸ���>����t�оF%3�h��S�����B�4Kr�I��>��O?G�?�(b��V��ATO�����C���o?�{g?��>.I?�??�;����w���p�=�n?F��?�=�?�>�W�=`����*�>�-?�3�?P��?�Ls?�>�.��>�k�:��&>�������=,t>H��=gW�=��?��
?.5?�i���
��&���Oj_����<Ɛ�=4��>��>��o>���=�O�=���=QX>7�>(&�>Y�b>�!�>�Q�>O�Ѿ��,�j�?�>�Fe>��=?F�>
��������f����.�|���V<=������=��v=�Ѿ=21����?lȿ��?w�>�!*���?�b��/�>��=v�>����A��>7
.>��>�m�>��>	�=�Xb>�>�FӾa>����d!��,C�]�R���Ѿ�}z>�����	&����w��YBI�|n��ug��j�P.��Z<=��˽<.H�?���� �k��)�
���Q�?�[�>�6?�ڌ������>���>�Ǎ>�J��k���\ȍ�hᾦ�?H��?�Oa>�߄>[�?�?��ʾ�맾P�l��'?�P1R��K���q���������P�/,ܽ@zd?�H|?)�?Zc����>���?�m���¾�� ?#�6�a�W�h�>��>�����`�Abؾw���߀��%�>}Ў?&��?��?]�վ�蜽�Z�>׏6?��>͜G?�EG?N�J?K���l�/?̇��s>?��>��3?���>�Z�=����t�=�i�=JՈ>-c��鱹��w���d����H�=L<=���>=�}�:�4��=�<MP�]�@:�#�<b�ļP�<q��<��>f�]?�@�>���>��7?���=|8�OĮ�#/?/�9=������3Ƣ�R�>z�j?��?_Z?�Ed>��A�dC��>�T�>vp&>%\>�]�>%��ǭE����=�H>d>�ե=�"M�*�����	�ԕ�����<�*>�u?>k>��2���>~u��h[��#�>8g����߾V�ѽOKN��9��JQ����>x�]?�+?,�4>T�Y<�!�E��K?\[#?U"I?!m?�6>���t�+�����|�>y�e=����y���Z��XQ@�A>Ȑ�>��Ѿ#�����S>������־OMm�b�D��bݾZ�<����)=ܧ
�iM꾇"��˽�=���=_G¾�("�ꗿ0����pK?a��=W����DA�sg���>b�>7��>>��p�>��I?�����Ef�=��>�6>�z��=�~�G����l>�>TQE?@W_?k�?"��Zs�=�B�����kc���ȼG�?ix�>'h?�B>r��=K�������d��G���>���>g��H�G��;���0��L�$���>W9?ߩ>��?[�R?��
?{�`?�*?IE?''�>+������ B&?4��?��=v�Խ�T�� 9�JF�{��>z�)?�B�ѹ�>M�?�?��&?�Q?�?��>�� ��C@��>�Y�>��W��b��2�_>��J?ۚ�>t=Y?�ԃ?��=>W�5�ꢾ�֩��U�=�>��2?6#?P�?篸>���>3�����=���>O
c?�0�? �o?s�=��?y/2>���>��=힟>υ�>>
?�SO?�s?(�J?���>�y�<�P���.���0s���O��X�;�H<j�y=���Dt�g����<,C�;�[��3+�����h�D�H6���=�;��>W~�=��ھ{#�>?���qz���;|�g����:ľģ�9��>g�>�i&?f<#?�E�;1��=��M>��?T�#�^�?(?��Q?�L>4n[���c��G��ɓ�>�N\?�Г<�AD�p�q�1,����=j^?'�?0�S
�O�b?��]?@h��=���þx�b����i�O?3�
?�G���>��~?d�q?J��>�e�.:n�)���Cb���j��ж=br�>DX�M�d��?�>j�7?�N�>�b>%�=iu۾�w��q��c?��?�?���?+*>��n�Y4�,��󐜿�3�?]�>�Y��;d ?`n5<����-����,����������u����ݣ��o_����,(����=wT,?��j?��T?�H?�S�v|���g�4�y��'X��vӾv����;���>��]G�T>h� �󾅪�����X>	(����H��o�?�)?�X����>�ᑾ����˾JTQ>�������=�H��_D,=/�= �q���E��@��H�'?�~�>�}�>;8?Uq\�@�,0�7�6�0���TE>�Ì>4F�>��>QE����4�>���Ⱦ�@c��k]��7v>�xc?U�K?��n?p�+1�����M�!�X�/��c����B>�j>5��>1�W�ŝ�S:&�pY>�F�r�n��-w��0�	�~�~=��2?w(�>A��>�O�?�?�{	��k���kx�2�1�6��<>1�>� i?:A�>%�>�н'� ����>��l?���>��>����1U!�~�{�gkʽ2!�>��>׸�>� p>�,��"\��j������9�=��=��h?�����`�3�>�R?Y��:��F<p�>i�v���!� ���'�.�>�|?ה�=u�;>��žQ%�h�{��:��KN)?�L?�璾��*�9~>�%"?���>�+�>�0�?n(�>�kþ�RA��?Y�^?C@J?}RA?�I�>n�=���.CȽ��&�g�,=l��>��Z>/m=΄�=���Vs\��y�e�D=�u�= �μyL����<Y�����J<��<��3>�dܿ�K�.�Ǿ��T��mJ�h�������݊����U���x���6��
��r�<� �W�J�c��]��sو�ģ�?ћ�?Rp��w�鐙��`z����j�>�^j���R���?a(�ve��D�־a���H�!��P�K�g��f�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��6�"���8�� >hC�<-����뾭����ο@�����^?���>��/��p��>ޥ�>�X>�Hq>����螾�1�<��?7�-?��>Ďr�1�ɿc���p¤<���?0�@�|A?�(�K�쾕pV=���>͊	?��?>�_1�BI�r���hJ�>�:�?���?�sM=�W�N�	�M�e?��<��F�I�޻u�=L@�=TL=���w�J>yT�>-}��EA��"ܽ��4>�υ>�"�a��g�^��s�<��]>V�ս\f��5Մ?,{\��f���/��T��U>��T?�*�>R:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=u6�����{���&V�~��=[��>c�>,������O��I��U��=c���ſx�!�']���<p�Ϻ�]�����V����>h��+����z����n�`=N�=%4M>B�>?�L>ajI>1�W?m?w��>.�>�F�
G����Ⱦ����3��e{�c����%������}8߾��	���N���̾!=�[�=�6R�V���9� �x�b�p�F���.?�v$>o�ʾ��M���-<�pʾl����ۄ� ߥ��-̾�1�0"n�j͟?��A?������V���U�=���?�W?P�����ꬾ���=+���"�=�%�>!��=���� 3��~S�q2?k�?&Zþ.���h�*>�����=c�-?�� ?�n�<R�>�f'?@r#�����O>��)>�@�>	U�>f�>�2���н�U?/S?u��	I���>)��O���A#�=�>.�3�����Z>
ya<3����[��`8��mV�<ǅw?�>�C��G������N�=3�T=��?�K-?hL�>+�h?�OX?�%ڽ΂��T�������w<��|?��f?���=tb>�Ǖ��������M?8�B?�.&>m>�������������*?��|?���>hӽϦ��;������-?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?n�;<��U��=�;?l\�>��O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������=������?u҆?���u�;D����k��K ��M�<"B�=����,<��\𾨹7��kǾ�#�>R���U;����>��@������>��1�r�㿨ѿ���.оNs��`?��>�%����Yj�:�o�*rC�֔C� ���ݳ>��=�X	�����f�R�E��!�;��>��"=Į�>�g�����G�~!��=�>x<?�i�>�X̼ ���?�{��ƿ�B�����B�h?[�?W(�?.#?��t�Y��IT2��ջ|�5?�XO?K_O?�e�@���	��B�r?O��b���B�[����]>��/?*?J{4�P��>�;U> q?��b>��,�S@����q5�~9�?��?���� ?Oě?�K?��澂e��2����F�ks����N?�g >�������w
'���%´>�i?��U�J�(�|rN?��W��)l�>��� =�;>���Q=\�
.��Ծ�n������Ͻ�:�?;�?F��?=ҁ���f?�1�>�*��~�Ӿz��WED>@ �>�;>>���]�*=�����CRa>H9�?i@~R1?�����X���>Pw�?`	�>���?�-�=��>�ď>�7��uc�=��>�6%�-��=�-?�E?q+�>,��`ޒ�mlD�{F���A�����h����>g�T?�	]?��~>ٺW�z|q<'�?!>SV����j��:��7j.�e���F�u>c��>�3>�7C��#پ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>B�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?I�4O���]~�x��7�\��=��7?�1���z>���>���=�rv�s�����s�d��>bB�?L{�?ۿ�>�l?�~o�g�B���1=.S�>ߚk?Ro?��m�����B>0�?d�����J�. f?=�
@u@�^?��hֿ����^N��R�����=���=ۆ2>�ٽ4_�=��7=\�8�5=�����=s�>��d>q><(O>�a;>��)>���P�!�r��[���R�C�������Z�B��Xv�Xz��3�������?���3ýy���Q�2&�?`�Ӝ�=�U?��Q?�p?ƿ ?��w�	$ >5����=K>#���=	�>fW2?�[L?�Z*?!�=����?�d�vV��n���.o��m�>�xI>qc�>�-�>��>0C�:��J>@#>>b��>�>d�(=JO���=��O>�r�>���>���>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?��f>zu>e�3�Oe8�v�P�g|��#j|>�36?Q鶾@D9���u��H��cݾDHM>�ľ>1D�l�����-�Eui�̙{=ix:?�?�7���ⰾʰu�)C��QR>�:\>T=-j�=wXM>bc�|�ƽQH��f.=Ļ�=��^>t\?��+>�f�=�ģ>�O���1P����>��B>�,>�@?�)%?���N�������.���v>R:�>��>�k>T�J�P%�=�t�>��a>-��������?��;W>֮}��~_��u���x=�)����=��=(� ��=�R%=��x?S՞��<��$+�b��ɕ?��>m�<��#��UA�B7��W���AG�?�@x�?�ܾm�f�Q;%?���?*rB�"��=�`�>:��>�3�%���$?�l�vA��I0ﾵv���0�?���?����|��}u�\�:>o�?�͒�]h�>{x��Z�������u���#=R��>�8H?�V��2�O�N>��v
?�?�^�ߩ����ȿ2|v����>W�?���?_�m��A���@����>4��?�gY?hoi>�g۾`Z����>ͻ@?�R?
�>�9���'�}�?�޶?ѯ�?aI>���?�s?�k�>�0x��Z/��6������ p=��[;�d�>�W>f���xgF��ד��h��u�j������a>��$=,�>QE�[4���9�=��I���f�<��>�,q>"�I>W�>v� ?�a�>}��>�x=�n��Jှ������K?���?-���2n��N�<Z��=)�^��&?�I4?k[�}�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��J��<��K>*4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��QS��GB�>�e!?���>�Ү=ܙ ?��#?��j>�(�>DaE��9��V�E�ɲ�>ޢ�>�H?�~?��?�Թ��Z3�����桿��[��;N>��x?V?qʕ>a���񃝿:kE�BI�I���^��?�tg?wS�3?=2�?�??^�A?s)f>���.ؾd�����>��!?V�9�A��M&���m~?�P?��>�8��%�սlLּ������) ?)\?~A&?��,a���¾E9�<��"���U�� �;�D�I�>�>ы�����=�>sְ=cOm��F6�a�f<�j�=��>��=�.7�[u��5=,?X�G��ۃ���=��r�7xD���>JL> ����^?Ml=��{�����x��.	U�� �?���?]k�?H��8�h��$=?�?D	?o"�>�J���}޾&���Pw�~x�yw���>���>��l���J���ۙ���F��*�Ž۔��F�>}u�>U?� ?`�O>���>�ʘ�ԡ&����!	�1^�����^8�4�.�f��Z��J�#�.��ntþ�Dy��G�>������>�K
?*|h>�P}>c��>=��,��>j�P>�>Ł�>^�X>��7>i>�� <n�ν�TR?�N��{<(�;Q羕��T@?�b?��>�^y�ǅ�/���?8?�?})�?�{>�fg��i+�vv?OV ?�K���O
?֋6=��޺ ��<=���<��`=��ͣ��>�߽�"8���L�trn�0�
?�
?��E�!3ξs�ս�������:i�?�+?ر<�Y1P�̇i��U�5#R��+�<^V���&����%��Vq�G��(���Z�����g�=:T-?r�?��O�侻���̃�	�]�N>�w�>�>l��>�Ѯ=Sx�{1�L<\�f�	��]A�I�?;�r?�C�>^�I?��;?4>P?�yL?��>���>
��/��>I@�;�S�>��>3�9?��-?�0?lQ?&]+?IGc>���b����ؾe�?�s?*!?�?G�?�%��6�ý�ޗ�E�a�O�y��-��E�=���<��׽+rt�"7U=�S>2l?{��X�8����Z�j>�7?�r�>�>�Џ�����g��<�@�>ԩ
?��>c ��sr�+\��m�><��?�� �=��)>��=Y���'AϺ)'�=�ļ�~�=��~��b<�+-!<n��=��=�K|��� ����:U�w;�	�<��?��?��c>�={>�������Q.�a�2>HӋ>_a�>�@>#e۾a����ԓ�tTc�Uυ>�ȑ?�f�?H�*=<>l��=�����k�g
�ay�����<�"?�'?#�M?G�?dE?��?6 �='��|呿�ފ�[gm��?�.,?�z�>���E�ʾ�Ԩ��x3��?1y?�Ja�����)�^ ¾�Խu�>�_/��8~�v��q�C��;q�����ǘ���?t��?y�?���6��a辡������S�C?���>�>�>���>�)�|�g�/-��;>1*�>��Q?%N�>�7O?�jz?��\?��U>�+9�8	�������G�qG!>r�>?g�?2ߎ?v�x?��>�>��$��X�-��k� ���p���W=�JZ>U�>���>���>���=�RĽbL��B�3̟=%
a>#%�>�j�>b�>�Tw>o��<SuO?��>�rо=v��B;��'���:�?o��?�O8?l�=����Q��������>��?0"�?c�6?�`�g2>��6�3���Aþ�:�>8��>��>-�p>�`=��3>9,?���>)�0������D�b�ֽA��>rY?B�>��ɿWX���;�p��C����������7���]�Qw}<��[�;�]��]�'����ۢ��ھ�K���;��g�?�>(�>�V0>wZ����c���[��^�=���=�r�=t|�Q�<����?�<I�U�-PO��ok�R���(l��H���ގ?��>�@>�Q?s?��?;Hн���>~}��xP?+��>[�1>Mգ���������佢Q�Ţ��4�˾�ƾc�>���-Ѽ�h >=m��JM>�t��%c=��	�-�Q=!��=�!�=�p�=&>|b�=��=�Mq?�=��F���[G��ݽ�+?�3_>>�=>�Ⱦ��2?�)>j���Vк���j�y?i �?�:�?$�?����pm�>mԩ�o����J=�� �^h> ��=�5�p^�>�V>+���ɒ�	0����?Y�@�"E?_i��4ѿ߫->e�7>�%>P�R�8�1�ݜ\�D�b�uzZ��!?�H;�PJ̾�8�>E�=�+߾�ƾÄ.=�6>�eb=�f�^V\�M�=��z�0�;=�l=g׉>��C>�v�=,4��
�=9�I=���= �O>�&��;�7�X/,���3=���=��b>4&>���>C?�>?e�?R��>R�þx�q��q�>���=b>�)r�@>xW�>��L?�xO?��?"�>S7-=>SX�>M���^p�-_�����l >�r�?�8�?���>3_5>�#����=�+�.� ���~�>#�6?��?(�g=�/������O6���(����-�q=@���;1��%�\溽'%���i>uB�>ᨾ>���>�HH>!��=O{�>��>�Z >?��<2%=:��xв�Ļ%�K�J=[�M��=qӼ� Q�}!�����6���R;_�y<�ޒ<�7=.?�=i�>9�>���>:~�=	j����/>�����%M����=yc���gA��c�x=~�Q&/���8�b�@>QW>�̆�K^���P?PZ>��A>�I�?�u?xb >�����Ӿ�|���e���T����=3w>Tn;�)�:���_�j�M���Ҿq��>���>܀>�A�=�����Q-��&�=����n�Y��l?�w-���=�����Qk�,����Z��Cj�?S��(?>V���w>A�{?��G?xz�?ڠ�>��������05>�ľ0�<t��s���۲�ũ?qm?���>���*�P�Q	˾ڽ�Q�>��8��uT�J����,1�~������̶>N����SѾq5�o�����@�,u���>]�Q?V��?�[8�/���L��P��۽T��>�d?{��>UV?y?�;潂������ȣ�=C�r?�t�?�N�?:��=�}�='�����>��?[��?ҿ�?тs?��?��|�>T�u;#2">�3��h��=�G>�$�=w��=WZ?�
?~�
?zߞ���	����W^�9��<�֢="ԑ>A��>U�q>��=(�g=0��=�J\>���>��>��d>�ӣ> �>J.�O���X?7�e>��r=c�)?�M>�gV=H�k���F=~���}���w�����u��͞��������u�r���#?Psܿ�+�?�M�>����{?�yξ�kC=S�=�b�>sD��5�?�[,>�(>�!�>_tp>��(>^��>D�>?PӾ�A>O��V!��3C�buR��Ѿ9~z>J�����%�=���s���SI��g���c��	j��+���C=�١�<ZL�?�^�� �k���)�; ����?S\�>
6?挾ϳ��k>���>~ƍ>BL��=����č��b�b�?���?Qe9>5rg>êY?o�?%��0�Ծ��p�S�W���?��7�^��B������o;�<U0���^?O�p?f�P?sw4={ҟ>�v�?A�p������>�/� 8j�4�=���>��=���~j�ɟ�)L��+��>��?���?�B?�c׾������>o�+?��?��c?�qA?B�P?�o=��>,?"C�<�X?��?(*5?x?���>p�=�t�=\��<��<���$���&�cLf���f�.=�<�~�=��=�_�"<�N���I�Y���")�-��:~�\�.Q<�Ƶ<�=ǭ�=BȦ>f�]?�>>�>��7?����x8�=��I
/?Ey9=|낾�	�����(�񾀩>\�j?�
�?�%Z?C�d>��A�2�B�W>fL�>q�&>�a\>�O�>(���D��u�=��>��>̹�=�N�s���	��#��KS�<]O>$��>��m>�ࣽ��Y>����/��rO>�}q�W����R��L��z,�QlX��-�>��R?�. ?w��=�&��0�O�մd��+%?.4;?#�L?z�~?��=��׾ؖ6��{?��x�-ߣ>^�V�³	�������5�HY4=��d>����Ƞ��Lb>X���k޾��n�JJ����M=s��aU=6��־��~�1m�=)S
>����X� ���vѪ�+J?hk==�����U��/��a�>���>]�>:�[qw���@�Ȋ���K�=��>;Q;>3}��w�݂G�(.����>�p>?��^?""�??�~�ieu���/�[��������F<�=
?�@�>� ?���=��q=ؚ�������_��l@�9R�>M�>���x�D��DǾX����*��R�>�.?�m>�8%?/�M?�#?��\?Md?&?�>�K�>P��`䜾g( ?F*k?��g��C�Y��a{0�)h�[��>%�&?.���灒=a��>��?@�&?	�r?J;?>���E���%�cV�>.0�>9�Y�;8��B��>Y�!?���>a?���?�u�>�*2���+���ؽc^��*c>}W?ZQ"?	��>�O�>.%�>W����+�=R��>�+f?�^�?#L~?kտ=��?�&�> *?��W>��>��>r�?y}C?��|?�KS?���>�/=��tkp�;�;\�<�]��3�@=V��=t�r^:��3��Z�<�M�����J�>������������<c�>��s>�'���0>%�ľ(g��HV@>i0��w���\���N�:�$�=��>j�?��>��"��c�=b�>�Y�>���7(?.�?�?9�);�b�]�ھ�K��;�>�B?m��=��l�Vx��+v���g=�m??�^?ӳW����֎m?®Y?���Q0�R�Ծo�I�9oӾ��^?�~?���G)�>ikU?��x?x�?҅�� �u�@��y�(�g�ؾ�N�=a�f>X��pd�$�>�$?[E�>���>H����N�n�Jݺ����>阎?;��?��i?ӽ>��\�I������ت�� �x?��>���%O?{*P�(ھ&�m�Tޫ�%E��_;�����g���5"���/��꘾{\���>��!?�t?G<g?�}n?��� cq��b�9m��u&�>����D4��*O���F�b4�WfD��엾G����ѽ��-=��~���A��o�?Q�(?�I2�v��>���j)�̾`�A>�m��)B���=�ѓ��o1=b�R=�g���.��&���? ?+��>�G�>d�<?��\��W>��1�{�6�$��!O6>�l�>���>P�>m�;��-��D�X�ƾ炾��ν�7v>�xc?��K?A�n?mp�%+1����!���/��c��{�B>�i>%��>�W�l���9&�Y>�[�r����v��=�	�a�~=j�2?(�>j��>�O�?$?�{	�_k��4kx�ڇ1����<2�>( i?R@�>\�>�н�� ����>��l?ܧ�>��>+����Y!���{�"�ʽS(�>��>˹�>��o>�,��"\��j��$����9�e��=ʨh?������`� ޅ>�R?CS�:�H<�z�>�v���!�U���'�`�>�}?Ġ�=.�;>��ž~%���{�D=���)?Gu?�&8&��>�>i�?��>�>lŁ?q�>T���s�?�{\?��V?��O?�H>?���>ǀ	<sܽ)ɽ�%���*=�_�>9YP>,=�=��=�]���Z�+��-~�=�=⼡��/��Q7������=�6�;�YC>>mۿ�BK���پ9��2?
�H爾���.d�����a�����Wx���	'��V�68c�����l����?�=�?����|0�����������i��>��q�u����w��X)�����{���_d!���O��&i�F�e�5�'?�����ǿ󰡿�:ܾ>! ?�A ?/�y?��6�"���8�)� >3E�<4-����뾩����ο?�����^?���>��v/��X��>Х�>'�X>qHq>����螾|0�<��?'�-?��>��r�+�ɿ]���k¤<���?-�@%�B?�k�7����*�<���>U�$?`��>3x;�"��b�H��>�ê?�V�?	��=�aN��S�ٝs?�@�=�6�?=�K<>��=���=�PȽN�3>�o�>�c���y*�������N>~{s>��P���%�F�L�slU<��B>N����6� Մ?�z\�qf�x�/��T���S>�T?,+�>�;�=%�,?h7H�B}Ͽ��\��*a?�0�?��?�(?�ۿ� ٚ>[�ܾI�M?#D6?���>�d&���t���=�Dἳ���U�㾐&V����=d��>��>9�,�����O�5N��A��=��u~ƿT�%��� �ʷ=��<�X+��ὺ鹽L�c��՟�қj���Խ��c='�=qL>(�>�UT>%_>C�V?�|k?��>��>�H�`݅�R�о�N��h����������� ��ע�N�fQྨi	�q��
u�&Fž��<��)�=�R��u��ώ ���b�U�F�N�.?�n$>��˾��M�S�#<-�ɾ؞���b�2~��x�̾˜1��m�r��?�A?1���E!W��4�	�t	����W?�)�M��H�����=���4
=麝>Q!�=<�>63�R�R��<?�1?��˾	N����>��K��j��m:?�V?ȏc>�Q�>�$?�У��&h=��|>Dn�=y��>)��>�nC�:�c��:S�*?�/?�i���["���>P�ྞ�f��rW<5!>׃��Y�0�=���}���&$�=�c_:ay�>��W?.�>� )�H]�n���	�"��J3=�w?Q-?��>o-m?MdC?���<Pr���IT�'��=s=��X?/`g?8�>L�}�CuӾ@譾%/6?��e?�7I>UW����I/�&.�t�?�p?�H?#i��-}���Q����/?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?r�;<��V��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�╾�Y�?9�?UЪ��Ed<����l��u���}�<.8�=���B"����7�o�ƾA�
�N���+뿼D��>�U@U�l��>S�7�Y4�9RϿ1���gо��q�a�?�y�>��ǽL��4�j�Tu�'�G���H������>��
>����ƌ���|��K;���h�>ɳ4���y>��]��Y���W��>I=��>�\�>��>c౽�U��޴�?]��ٰο���!��&�T?#V�?�8�?h#?��Ի/+~��}l�%��;ѫE?m[w?��Z?�N��5�m��$�%�j?�_��wU`���4�tHE��U>�"3?�B�>T�-�k�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*�F�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�\TS?N�R���W��#��*���p>
�������;ν���;�g��+��3�/�QG�?s_�? ��?��d�����?�]�>��I���TC���>Nڬ>b�&=9�$=��>r���;�#�X>���?�~�?�f(?�Vx�B�����g<�"w?�>���?(j�=ď�>��	>mq���K���/>��>,¸���?� N?���>��=�:5�Q./��ZA�d�L�O��A����>1<b?#J?ڱ]>y����� ��˽��.��̼�NA�.�)�&���'>+�H>��>�t=���ľ��?Np�7�ؿ j��p'��54?5��>�?����t�����;_?Gz�>�6��+���%���B�^��?�G�?<�?��׾�R̼�><�>�I�>1�Խ����V�����7>)�B?i��D��l�o�{�>���?�@�ծ?ki��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*i�̿抿�浾H����>���=_W>�\�w
i��e�=��<_�x�MR>��.>� �<�`�=�Iu<�ټ>L��>'|���>�F4���"��es;���>��M����3�����5��W�`�T�0��3a�)m��*1;��7ʩ=�X�=D�U?��Q?p?h� ?B�x�7�>4u��	8=#�Q��=C�>�[2?*�L?ݒ*?x�=����r�d�Vc��gC��1���}��>�jI>�a�>!N�>9�>-8X8r�I>?>���>�� >�Q'=Vx��sf
=eO>�W�>���>˚�>3G<>8�>zδ�*1��u�h��w�@=̽� �?<w����J�62��28��X���%\�=�e.?��> ���>п2�K0H?����?(�ߺ+�G�>X�0?�aW?��>���ѦT�76>!��^�j�rL>) ��|l��)��Q>�k?�$j>�h|>��3�l�8�k�K������"c>��9?Y/���yE�X^w���E�A׾�6>��>�SM<������~�x��h����=q?9?��?"��2h����q�� ���N>�`>��)=�}�=�;S>�	����Ľ��C�$Kl=$�=��Y>�[?��4>ו=`�>�k���I��>�yE>@1>g�A?@G'?Q<��+����Y~���.�i7p>c�>�j�>��=S�J��e�=�C�>�ta>�W�Fs��� �7�B�MS>�~���X�r�b���t=#&��$��=V�=K�(6�7�O=�~?���(䈿��e���lD?S+?] �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��L��=}�>׫>�ξ�L��?��Ž5Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l�6>�^%?��Ӿeh�>Bx�}Z�������u�H�#=@��>�8H?pV��e�O��>��v
?�?�^�ީ����ȿ(|v����>L�?���?Y�m��A���@����>6��?�gY?�oi>�g۾e`Z����>��@?�R?"�>�9���'�o�?�޶?���?�I>���?
�s?�r�>�x��Z/�4��T���"f=LK\;_�>_> ���iF�ד��g��&�j������a>N�$=j�>�M你2���#�=J��I����f����>54q>��I>K\�>Z� ? a�>���>�W=�p���䀾�����kP?zd�?͖��i��tb=g�u=� [�1?�+0?�@=WB��Mԭ>-�S?�5�?.Q?WB_>����Ԏ��ǿ�k��~o<�@>�>��>hꎽ��>>B�ҾAo*����>Ӯ�>\&=�E�ܮk�l��<v�>��?l~�>պ�=4�*?��%?M�n>7�>��g��u����&�>�>C�?��3?��?��+?�����.�]�������{*�_��>3�_?�_,?u��>m����t������} >��~��?T�@?)�b�z;?�vF?B�M?�wE?�!>���F����6�=W�=H� ?93�� �C��&���;��>���>n:�>�C�<���������\�ݾm��>C?h?bf/?�3���f�
7���(�<@9�;�?z�o�< y;���=�)>�{�f�=�*>���=�nM�PGV��fֹ��=F`�>�i2>�bH�$���/,,?�8B�!y���|�=��r�DoD�W�>
RK>q'��2�^?E�=�} |��'���o����T����?��?'_�?�д��h��<?�+�?g"?44�>�箾�ݾ�྆�w��Iw�����>���>��|��I�=���������~�ƽ�!�#��>���>!�#?v?��B>���>[�ξ� -��ԾO���D^�S�6�h�D��~&����,u��:��ٷ�'��������A�>,'����>g7?n��>U�Z>}��>4S <(�_>��>/!�>�\�>�v5>t� >�|p=���^�zPR?�����'���
����'B?�dd?I�>��h��|��ǵ�4v?B��?�s�?�.v>h�1&+��o?���>&���g
?�9=`�Z��<O��x��%������>T׽�:��M�h:f�r
?*?[:��X�̾��׽�ڟ��Wp=!B�?o�)?��)�#R�?�n���W��QR�K��0h�����s�$��p�gƏ��0�� ����v(��	)=ث*?�?
����"����j��t?�X�g>�C�>��>���>@nI>)	�u1�^��h'�܇���e�>]Y{?���>��Q?�<?��??�JN?�d�>mұ>OL��ٝ�>]��=;��>�>u-?��(?�?YF?��2?^
�>vp�H� �5�Ծ	� ?�]?B�?@�?�5?"I��rν�^.��;�X%��9�T�F=����s���˺y>�=�r�>�w?���ڽ8�(�����k>�>7?K5�>_&�>^����b����<l�>Ζ
?Ǐ>s���f}r�o'�-Q�>�7�?���M�=o>*>4W�=
����غN�=5�ż�t�=V���_&;���"<
�=��=�<~�I��9�;��;[�<�b�>�n?���>��?� �4��{0��kX�+/%>y�|>�%���b��h���L���HR��9>E��?`�?P.�;�x>9��=�׵�Z\���"�&྘�?��/
?"�:?�^?�Q�?�GV?RF?�4>.��>��R8k�'H����?v!,?��>�����ʾ��։3�؝?e[?�<a����;)��¾'�Խѱ>�[/�c/~����<D�U���]��5��?쿝?%A�R�6��x�ڿ���[��}�C?�!�>Y�>��>V�)�~�g�s%��1;>���>gR?I$�>��O?d7{?S�[?�aT>Y�8��1���љ���2���!>@?K��?`�?7y?F}�>��>k�)����M��\��D��₾W=�Z>k��>'*�>ީ>���=4Ƚ/N��-�>�+0�=ʖb>���>���>9�>iww>>d�<�B?Mz�>�;����v���r��y��WЀ?s��?�?��Y�~�/�
����>Cū?��?��?
S�w��=�<&���JO?�	�>nט>�s�>U�=�K)=�0>?�>��>�ܽ���ޅ,��B���?�8?�4�=��̿5~�ܢ߾)�
�Y�4>��^��@F>�F�<�����������[[��P�0Č��\����{���4���_N=(��>������>`N�=4����r>��S=�s��t�<g�%��V���Mu��=i\�=��l<F*�=$�@= �S�I��f*˾"�}?*I?t+?K�C?g�y>�Q>�2����>�����_?�}V>o�P� F��^�;������̔�P]ؾ��׾<%d�	����	>NI�B�>�o3>Bm�=%��<ѝ�=�r=��=p�;�v5=��=�y�=�̬=���=�K>�>�6w?X�������4Q��Z罤�:?�8�>^{�=��ƾo@?|�>>�2������wb��-?���?�T�?>�?@ti��d�>J���㎽�q�=@����=2>g��=u�2�R��>��J>���K��;����4�?��@��??�ዿТϿ4a/>�~x>��)>�kY���/���"��a�7�V��k-?m�'�������>���=̰ɾ�އ�X=$k�=�s=��ν]uz�fJb=�x���-=.*C=�X�>��.>_��=��གྷ��=�_�=:��=��>��E�V���~��ڇx=T_>}�@>8>'>UL�>#]?0
0?�e?y��>��r�l�;��¾�/�>Xm�=Ԯ>ʿ�=VB>���>�6?��C?��J?�ׯ>$ʉ=%p�>o��>܍,�0�m����;h��1+S<��?�E�?�c�>�J�<�>>����&F=�}ɽ,�?��/?��?�&�>Jj��+�-)�T�/���a��~�<�ީ=k�b�޲����(�E��ڽG��=�d�>��>-/�>YnW>8�&>0�M>#�>�>���<�F=&r��FB=p��;qu="���
��<A۔��~�<�n =�-5���>�R>D<!r�Z�Y<-��< �=���>��>��>�=h����$1>���� M�sv�=����@�B�D]e�߉~���.���4�"E>��Z>�����ܑ��
?vQ[>��A>=$�?��t?g"#>8W�r@վ�����Sg���M�2�=�>4�=�/G;��y`���L�<�Ҿ^��>Yߎ>+�>��l>�,�J#?���w=��_b5�|�>�|�����)��9q�@������Ui�KNҺ�D?�F��&��=y"~?�I?^�?��>q��݆ؾ�:0>�H����=f�z*q�}i����?'?���>�쾨�D�q5̾����>x�H���O���D�0�� ��������>s諭��о�3��g�������B��r�@�>��O?W�?b�gT��XVO����i���W?(|g?�:�>k[?a?���'b��[��/�=S�n?��?9�?�1>:k�=�����U�>$	?D��?xّ?E t?�>A�{��>"�<P}">$����=u�
>*��=��=�&?O-?�l
?!Z����� �ﾽ�ﾳQ\�Q�<�n�=ԝ�>ɉ>�t>�z�=��n=탤=�~Z>[D�>J��>�b>�¡>F=�>�$ྔ�5�Z�8?	�5=S�>�\?�Y�>��wQ����+����=�d�Γ�����O�Z�.����L#���Ƚ��C={w�>Dѿϗ�?C��>�n(�q(?{|�8��&�>�%!=/n�% �>��7>ty�>��>�W�>�ּ=X��>�d�=�4ԾYt>�����!���B�oR��JѾ�0z>i=��^�%��v�����*I����}��;j�wA��M�<�\�<�ۏ?������k��)����1?xb�>�6?�l��N~���>�`�>��>�0���s���Ѝ�a��C݋?���?�9>�`>�z?�j4?�;�Wi	�~M�"s��u�-�JQe�k�V����F7h��K���D���:b?��x?^�G?�@:=���>�:�?/9�����)՜>�js��qD�9��<I>Ru�����S����=o[�>�f�?7�Y?��>ڤ���Il�7_'>�:?1?OUt?��1?�|;?(T���$?	�3>W?�x?^A5?��.?��
?��1>f9�=�^��n	&=Tb��̊���нnBʽ�t��Z4=x|=��u���	<%]=���<�e�hyټ[f;N����?�<:=�'�=���=�N�>�`?�G�>�6�>�1$?�k���2A��b:��%?䞇��dɾQǾ���|o���>i�y?T��?�?k�>�9���%�V7<>=o�>M��=x˓>�>����aN�����=?#�=�N�=�NU=̉O<�_~�$�b�����=� �=_/�>|��>���Ո�>�Ê��ǰ��~�=5K���O��r�����>�Q�:�1��U?�>�HI?#?��><<�,��<�nF����>�X?)3`?<c?4W
>��Y=��Q�/�X�@;q> %P>hY����:�����s��TpX�>��=T�>H���ޠ��Ub>���s޾5�n��J����6HM=���YV=F�t�վF4� ��=�#
>θ��j� ����I֪��0J?ڥj=�v��z`U��n����>��>�ޮ>�:���v���@������2�=Ҷ�>� ;>_������~G�48���>-�F?�h?�?��_�!,d��A*���X҆��$q=��?5a�>+��>�>W7=7�Ǿ����X���2���>8��>(��O6�2mľ���PV.�S��>;�?���>��?�lO?�?�fP?�?�"�>g+�>=�3�,g��ѳ*?�%{?�̇��:����ă7���r�rj�>��>SX־u��n�>B4;?$m=?�׉?!K?  ��lw��n��-u>�6�>��H������q>T99?�?��l?�A�?�IW>3�!�M���l�L�t�_�"=�,?�j7?��?�OM>œ�>E���.��=n��>	c?�0�?a�o?[Z�=��?52>A��>�Җ=n��>I��>�?�PO?;�s?��J?��>i��<S0������1s���N��ք;�rJ<Ӽy=���u&t�J��l�<�O�;!�������3�IE�T0���n�;��>�qv>���X->�þ�͉��A=>i#���G��嗍��A���=V}�>�s?L��>,��0B�=ʥ�>�<�>�m���'?K6?W�?�]ʺίa�y�վ4E�@>�>%�A?��=>m������xv��J=�0l?K$`?��N����Q
r?��m?���K'-�����i־t�۾��|?:�>r���S�>���?4$�?�?�>��]�wk������\��*��� �=|E�>��!���f�%��>�=8?kl�>N{�>��5�/+����.˲��t�>�E�?9j�?�w?:L�=0z�I�W|ھ�0���FL?md%?�� ���D?O���:�������W~��������~�1���?�H�ǭ��(c(�Ϊn�:c$���P=w?�Yy?�w?v\V?�v�m��i�j���q��^��
�w��IX��6�ި2��XR�F���y���fሾ��>|�q���=��;�?8,?O2��B�>_G���s�����>�A>�o��������=����4h�<˄�<>Br�~ 8�9~����!?���>�>J�>?��a���>���5�̖7�ڭ�·@>��>�%�>ۭ�>T:�;��/���޽�����y�.C���8v>�xc?ԏK?�n?k�'*1�m���7�!���/�b����B>Sl>���>|�W����.:&�Y>��r����8v����	��~=߯2?�'�>ݲ�>O�?3?@{	�	g���ex��1����<o0�>i?�=�>��>�нR� ���>v�l?�U�>�S�>�A��f(!�y$x�;MϽ�^�>uK�>��>Zon>��7�B%]���������_�7��[�=/�f?)H��:a���>��O?��e<�}�<�ƣ>�y�_*#�����>�8	?�H�=�7>��ɾ���(�{����sP)?7L?�璾�*�d:~>;#"?��>	0�>�0�? *�>YqþDD�R�?��^?"BJ?GSA? F�>��=���M?Ƚ@�&��,=��>%�Z>a+m=b��=���2n\��r���D=�u�=�μX���<�p���K<D��<��3>&mۿ�BK�}�پ�
��� ?
�z爾E����c�����/a������Xx���('��V��5c�����p�l����?�=�?P����/��ղ������������>�q�����������5)�����ӿ��Bd!��O��&i�<�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >ZC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾x1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@}A?��(�,���V=���>�	?��?>�S1�&I�	����T�>`<�?���?-{M=5�W���	��e?/j<�F���ݻ��=I>�=�I=[��;�J>�U�>ك�SA��<ܽ��4>�څ>K"����/�^�'��<7�]>��ս�7��0Մ?�z\��f���/��T���T>��T?/+�>�9�=Q�,?|7H�R}Ͽ�\��*a?�0�?���?�(?1ۿ��ؚ>|�ܾ�M?MD6?���>�d&� �t����=3��k��/�㾶&V�Y��=ӫ�>��>��,���^�O� C����=P�#��c�=���0��g�<&#>��!=��o������<��+����ё��v�_�ؽ]��=��?2��>0;�>u�8?��<?���>��>�=������䶾-��B~���k���m�\X;��E\����������[��ڇ
�j6J�^��� =���=�7R������� ���b�v�F���.?At$>M�ʾ��M�v�-<znʾ0��������ԥ�|+̾�1��n�0̟?7�A?����k�V�+���R��r��įW?I�'��T묾C��=�ݱ��=� �>��=���=3��}S��0?��?�#�������%>?��L8=�E,?�?k��;�q�>D"?b&/�X8罅�]>�39>�/�>��>��>K�����ٽI&? �T?}��蜾�=�>)���&s�V=r�>�~5�"��V>H��;	x��=��������<j(W?웍>+�)����`���]==>�x?Ȓ?�-�>{k?��B?KƤ<�h��k�S����`w=a�W?�)i?ֹ>�����оr�����5?�e?�N>]bh������.��T��$?E�n?�^?B���Jw}��������n6?V�v?|s^��s�����c�V�>�>"\�>T��>R�9��k�>O�>?�#�~G�������Y4�&?W�@���?�#<<��⛎=�;?D\�>A�O�x;ƾ��������m�q=��>≧��cv����@U,��8?���?���>�������t�=@��`U�?8=�?����:m<���Ql������ܘ<�I�=#n�)j&��B�g�7�a6ƾ�X
�7���㙺�,�>6_@�?�y�>�g8��f⿨6Ͽs�Ѿ)�q�<<?�ݨ>��ƽqZ��I�i��t�(.G�NlH�ц��U`�>��>G���󏑾�|�b�;�h0���_�>Ek��Z�>�]T�PǶ��x����M<�"�>�>�>����ݎ�����?Р��^?ο�����_��_X?�0�?m\�?��?*�)<;w�9~{�F���pG?��s?�5Z?�c)��]��6�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�znT?��"��f?�¿��3����<g�!�پ����x����v������Y�;���?%��?.�?p���_G&��+?��>�h�@��9}��?]l�>�M߼n?�=;�/=w����>�2)�>�0�?'�?�V?�w4�ݮ�|�V=-�u?)q�>���?��>���>�>�:���<<��<>#>���3?��I?���>���=��1��?-�P�H���S��M�^�?�On>�e?�Q?��Y>���*��&�=����N�)��<�P�2?]��F����>K�J>Et(>�5,�W��	V?�����ؿ�x��C�'�O�3?�T�>��?c9��r�Ll��h�^?�ц>�^�e���O����������?�(�?��?�H׾B�ļ5 >�;�>�,�>�ԽX���ň�L�4>JQB?}c����?yo����>�u�?mo@�O�?P�h���?�&�%T��yd~���&�6����=N�7?�#��z>0��>�5�=unv����c�s���>PB�? �?R��>�l?qxo��B��(2=�P�>��k?�l?�-s��f�B>�?��������K�f?��
@�p@P�^?U좿!&ʿ\G��A���+�Q �W�g<��P>�Ľ�.>�wh>A�_>fPۻe:>�O>��>�R> ��>�#�>���>w����M�2ٱ�rӡ�6kR���!�Dy
�<*�"(�P	����,ʾ'��R@�Œ�xQi�b����=�x�=O�O>�R?�`?[�j?�1?j&��=Q>�Ҿ$>do,�E(>8��>s�*?��6??Z?I1�<>����c��c��/]����J�?>�>�S�>Z�>�>X6�z�D>+:>
g�>��}>�w\��Sټ�m0��Ch>��>q�>p�>�^<>��>�̴�.���h��w�to̽d��?���v�J��6���;�������v�=�s.?�>O���:п�ꭿd'H?L씾�%���+��>ջ0?ZuW?7�>�۰�a~T�F=>�����j�G>�s �ӗl�Tk)�6hQ>$V?��f>�1u>��3��d8�}�P�?~���M|>�56?�eh9�5�u���H�~Mݾ�FM>R۾>�=A�Sk�����	�Yti�a�{=er:?B�?y^��vذ��fu�9,���R>�C\>v�=�,�=l(M>2 d��&ǽ�H�k/=�=!�^>SO?38->��=i�>�e��X�O�S�>ݰ?>�,>�??��$?��>똽������.���t>�,�>�1�>�>#I�}�=�!�>�4b>��&���H���A�drX>ul��\�C}p��1�=�|��K2�=[3�=P��� �:��+=��~?�`��&݈��׵��9D?��?XO�=85<��"����h<����?��@u��?�-	�Q�V�G�?�B�?락J�=�>�>��>ޫ;�=L���?��Ľf����u	��Z#�UO�?v�?�w3�����o�k�;>L>%?ӐӾIh�>�x��Z�������u�l�#=R��>�8H?�V����O�_>��v
?�?�^�ߩ����ȿ2|v����>X�?���?g�m��A���@����>:��?�gY?voi>�g۾?`Z����>ѻ@?�R?�>�9��'���?�޶?֯�?e�J>�K�?+t?���>;�e���-���������m�~=O�;�>~F>G��E3F��H��?��4sj�h���`>��/=]q�>*�����%��=9�������{��D�>�f}>�O>���>8�?���>�ԗ>��=�s����y�����u�W?��?����Y�pYx>�ҼT̽ʚ:?
�!?�T=aSξ�b�>o�d?�i?ʞ??�B�=?�"�vA��2aο̗��F~�MR�>��>T��>�һ=滍>b���܏��/�><��>F7��\>����~���'����>O�?t+�>#���4(?�0?a�>��>�<@����'x6�k�>w��>*)-?�ۀ?vM'?j�f�U�1�W��%��ՙL��A>�i?�T#?�w�>���ta��C�Y�3�U�ɮC�V��?�?N?�
�t?�܄?1�W?[)4?�E>��d��ӾQ.��[�>["?tw�x�A��&��� �fn?N��>ߴ�>��ν�0��8a�z'�-��ye?�c?S�+?�	�yZa�/t��
��<�s���*�N���Y��>==2>~�;��`�=�>n?�=�ge�a�@�������=� �>���=SP6�*����#,?\[8=�#��+�=�$q�_�F�ס|>c`L>�l����H?�1h�N������yV����O�Փ�?���?v�?��׽�Pb���/?�O�?�?���>\���w�� .���e\�; ����]�3>�[�>����v]�;묿-���ˇ��Mh���"���>�^�>eM	?آ?��P>s��>?֚�R��X[�H4��[��y���9��-�%��Ꝿ�*���@�����v����>�Ր���>��?sr>˝q>���>�UX<���>&�^>�b�>f�>�N>��>�=�vֻ�H���KR?����$�'����󰰾2B?Tod?]0�>�,i�i�������?ۆ�?ys�?;Dv>�|h��-+�>m??�>��� q
?�N:=�b��T�<�T�����:,����C��>hG׽�:�}M��rf�j
?0/?F����̾3>׽���� �=(��?ݣ)?��'��pP�9�l�eY���P�Vh�ʀe�����#���o��7��C:��񯃿��'���/=h*?�Y�?���,���᰾˶l��?�&Nc>���>�ל>;�>��L>j��50�!�\�QC'�X���Uk�>g�z?�>�pI?�<?��P?o�L?�ώ>_��>�鯾��>)s<���>e��>)o9?Ө-?��/?
?��*?�<a>��������H�ؾ m?f�?��?�^?��?�z����ý૙���>���v���3�={8�<#�ֽ�o�}X=�aV>�X?X��]�8�)����k>n�7?_��>��>����,����<��>��
?`F�>A �~r�c�7V�>m��? ����=��)>���=r���l�ҺCY�=N�����= *���x;��o<��=���=
Nt�恹�$�:���;�r�<'��>��?�n�>���>����@����w˰=A�^>�7N>��>�/ܾ�������w�f�[Zz>6��?x��?��\=�`�=���=����S켾_9��¼���=��?�"?zU?�ђ?I2>?�!?���=���;��O���>٦�|{?{!,?5��>n��x�ʾ�񨿿�3�ܝ?f[?`<a�����;)���¾s�Խ��>�[/�T/~����BD��
��������+��?꿝?�A�7�6��x�ٿ���[����C?P"�>5Y�>b�>K�)�w�g�V%��1;>��>nR?�!�>�vO?*w?�`X?��W>��8�ΐ�����K�u�>��9?%P�?���?�v{?���>]->N(8��q�Q���'<��*���/=��c>'|�>���>c�>�m�=ˋ�������_3����=wsM>mD�>���>a��>"q>�˧<��D?"6?z�Z��jȝ�󢾟>v�D��?M�?(��>��_�l6+��-��r���>v�?e�?#'?�g>�W��=i?<�W��ن���$>Q��>�-�>9��<4:�>�;�>\�>1�P>��Ծ!���Fj������fA?��Q?�4�����͜x��<ӾL�����=�H�<�e>V�M�IĽ�B~>?%������X
���Ծ転�J�ٽ�<>(�	=��>�"=��o=}>&rn>@� >{B>�I�=�X�[&&=􅰽�������$��([���u½M���Y�>§=(m�.k?	�p?C1?�E?^��>���>�ֽ>��	�?�޵>qͻ��"ľ�X�#:��ۧ��=��w�پ��/�������->��=�-�<2a>L�=�W
�F}>=�t>�@=2�K<���=�>��>Vl6���=��w>o[>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>Hj5>.C>��R���1�n%\�aJa��Y��e!?�;���˾ģ�>m�=��߾<Ǿ5G)=��5>��h=����[��s�=��y�݊?=�+p=��>B3D>W�=�q���{�=�oG=�=�= �N>�����~5�3m+�A�1={��=r`>S�$>���>|�?z,?U�`?���>�p�[(Ҿ ���P��>>W�=��>A�}=KI>�T�>Z9;?�F?��H?7Ĭ>���=8ȸ>�:�>f�+�Xdk�#��찥���%=C$�?a��?���>O�o<�G����n�@��߽�u?�4?{
?��>�s�m7߿�w&���-�)딽X<��L=c�q�ݪM��ҼV�����K�=���>��>�ޛ>�]�>�E>5T>�Ӿ>��>]��<��=!��;���<�&���V�=8.��t\�<�!�&�~���4�p3��X�v���	��US<�^�;�
�=���>��1>�6�>�q�=�y���XE>����Y?�ݏ�=�����:�.ri����l.���8�k09>�.>o�v�b����>i�v>�l,>��?o�u?E�0>ƹ����؁��{�9��"��Y	>���=�?�K�A��k���P��]��c��>qߎ>=�>��l>�,�F#?���w=��=b5�d�>�|������)��9q�@������`i��Һ�D?�F��1��=p"~?�I?a�?���>���φؾ�:0>�H��V�=<��)q��h����?�'?���>�쾄�D�Mm̾}�����>��I�� P�۽���0����������>Pت�f�о�3�>e������ �B�r�E�>�O?��?rIb�	Z��JO�������o?lzg?��>�=?*?�����x��,�=��n?���?�=�?	>���=C;�����>B�?궖?sؑ?+�s?�j@�J��>W�<��!>�V��_��=�>���=�=�9?�Q
?
B
?�ؘ�!\	����C�* _�� =�.�=�̐>���>Us>��=��u=Bi�=(r^>ì�>'o�>�d>�U�>겉>>g̾��$�R?TK>���>=�^?��>8dS�Ō=�Կ=�W=���}3v��>7�mHG��&���3���=��:V'?"�����x?Y��>�@�U�
?)�#�����ݷ> 砽���N<?鞇>��>�C�><٭>�0,>oi�=?@�=EGӾM~>����d!��,C��R���Ѿ	}z>"����&�q��`w���BI��n��xg�Pj�.���;=�yֽ<�G�?����k���)�������?s[�>�6?�ٌ��	��;�>���>�Ǎ>�J��E���6ȍ��gᾰ�?��?E�f>B$d>Eij?�+6?ib����=�J�c�Q���a�7��e�(�Y�ޔ�[�|���Ѿ�q���`?)r?z�&?`J�=�)�>_W�?��s=Ͼg�>%�k�v�E�� ;`m<�8澶5��������H�=��>.�?��n?��?�)����en)>�6F?��5?��p?�6?�??xN�("$?>�A>f7?�U?r�/?ٽ)?j?�$>J�=���8W<3Ė����Ѹ������1�-c=���=�0��klݻ�	`=�x�;����������;9^��@�;ӡ�< ��=��>ߔ�>3�]?/a�>%��>Z%6?�d��Y7�$_���/?AP'=�������[-��'N򾃐>��j?x3�?A�Y?Q�a>��B��nB�_&!>=T�>�0&>z�Z>�W�>֙��B���=l:>�@>�$�=9 Y�xz�����pr��.�<�>�7�>^
�>c6����>�Z����vL>P%6������w���N���1���f�W��>,�Q?Ɍ$?�Ҟ=�J龾烽�0a�g&?�8?2J?��s?�'�=�G��"l/��1:�?�SI�>��<�Oe�>���ˣ��=�7L=�م>|���Ƞ��Lb>X���k޾��n�JJ����M=s��aU=6��־��~�1m�=)S
>����X� ���vѪ�+J?hk==�����U��/��a�>���>]�>:�[qw���@�Ȋ���K�=��>;Q;>3}��w�݂G�(.����>�p>?��^?""�??�~�ieu���/�[��������F<�=
?�@�>� ?���=��q=ؚ�������_��l@�9R�>M�>���x�D��DǾX����*��R�>�.?�m>�8%?/�M?�#?��\?Md?&?�>�K�>P��`䜾g( ?F*k?��g��C�Y��a{0�)h�[��>%�&?.���灒=a��>��?@�&?	�r?J;?>���E���%�cV�>.0�>9�Y�;8��B��>Y�!?���>a?���?�u�>�*2���+���ؽc^��*c>}W?ZQ"?	��>�O�>.%�>W����+�=R��>�+f?�^�?#L~?kտ=��?�&�> *?��W>��>��>r�?y}C?��|?�KS?���>�/=��tkp�;�;\�<�]��3�@=V��=t�r^:��3��Z�<�M�����J�>������������<c�>��s>�'���0>%�ľ(g��HV@>i0��w���\���N�:�$�=��>j�?��>��"��c�=b�>�Y�>���7(?.�?�?9�);�b�]�ھ�K��;�>�B?m��=��l�Vx��+v���g=�m??�^?ӳW����֎m?®Y?���Q0�R�Ծo�I�9oӾ��^?�~?���G)�>ikU?��x?x�?҅�� �u�@��y�(�g�ؾ�N�=a�f>X��pd�$�>�$?[E�>���>H����N�n�Jݺ����>阎?;��?��i?ӽ>��\�I������ت�� �x?��>���%O?{*P�(ھ&�m�Tޫ�%E��_;�����g���5"���/��꘾{\���>��!?�t?G<g?�}n?��� cq��b�9m��u&�>����D4��*O���F�b4�WfD��엾G����ѽ��-=��~���A��o�?Q�(?�I2�v��>���j)�̾`�A>�m��)B���=�ѓ��o1=b�R=�g���.��&���? ?+��>�G�>d�<?��\��W>��1�{�6�$��!O6>�l�>���>P�>m�;��-��D�X�ƾ炾��ν�7v>�xc?��K?A�n?mp�%+1����!���/��c��{�B>�i>%��>�W�l���9&�Y>�[�r����v��=�	�a�~=j�2?(�>j��>�O�?$?�{	�_k��4kx�ڇ1����<2�>( i?R@�>\�>�н�� ����>��l?ܧ�>��>+����Y!���{�"�ʽS(�>��>˹�>��o>�,��"\��j��$����9�e��=ʨh?������`� ޅ>�R?CS�:�H<�z�>�v���!�U���'�`�>�}?Ġ�=.�;>��ž~%���{�D=���)?Gu?�&8&��>�>i�?��>�>lŁ?q�>T���s�?�{\?��V?��O?�H>?���>ǀ	<sܽ)ɽ�%���*=�_�>9YP>,=�=��=�]���Z�+��-~�=�=⼡��/��Q7������=�6�;�YC>>mۿ�BK���پ9��2?
�H爾���.d�����a�����Wx���	'��V�68c�����l����?�=�?����|0�����������i��>��q�u����w��X)�����{���_d!���O��&i�F�e�5�'?�����ǿ󰡿�:ܾ>! ?�A ?/�y?��6�"���8�)� >3E�<4-����뾩����ο?�����^?���>��v/��X��>Х�>'�X>qHq>����螾|0�<��?'�-?��>��r�+�ɿ]���k¤<���?-�@%�B?�k�7����*�<���>U�$?`��>3x;�"��b�H��>�ê?�V�?	��=�aN��S�ٝs?�@�=�6�?=�K<>��=���=�PȽN�3>�o�>�c���y*�������N>~{s>��P���%�F�L�slU<��B>N����6� Մ?�z\�qf�x�/��T���S>�T?,+�>�;�=%�,?h7H�B}Ͽ��\��*a?�0�?��?�(?�ۿ� ٚ>[�ܾI�M?#D6?���>�d&���t���=�Dἳ���U�㾐&V����=d��>��>9�,�����O�5N��A��=��u~ƿT�%��� �ʷ=��<�X+��ὺ鹽L�c��՟�қj���Խ��c='�=qL>(�>�UT>%_>C�V?�|k?��>��>�H�`݅�R�о�N��h����������� ��ע�N�fQྨi	�q��
u�&Fž��<��)�=�R��u��ώ ���b�U�F�N�.?�n$>��˾��M�S�#<-�ɾ؞���b�2~��x�̾˜1��m�r��?�A?1���E!W��4�	�t	����W?�)�M��H�����=���4
=麝>Q!�=<�>63�R�R��<?�1?��˾	N����>��K��j��m:?�V?ȏc>�Q�>�$?�У��&h=��|>Dn�=y��>)��>�nC�:�c��:S�*?�/?�i���["���>P�ྞ�f��rW<5!>׃��Y�0�=���}���&$�=�c_:ay�>��W?.�>� )�H]�n���	�"��J3=�w?Q-?��>o-m?MdC?���<Pr���IT�'��=s=��X?/`g?8�>L�}�CuӾ@譾%/6?��e?�7I>UW����I/�&.�t�?�p?�H?#i��-}���Q����/?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?r�;<��V��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�╾�Y�?9�?UЪ��Ed<����l��u���}�<.8�=���B"����7�o�ƾA�
�N���+뿼D��>�U@U�l��>S�7�Y4�9RϿ1���gо��q�a�?�y�>��ǽL��4�j�Tu�'�G���H������>��
>����ƌ���|��K;���h�>ɳ4���y>��]��Y���W��>I=��>�\�>��>c౽�U��޴�?]��ٰο���!��&�T?#V�?�8�?h#?��Ի/+~��}l�%��;ѫE?m[w?��Z?�N��5�m��$�%�j?�_��wU`���4�tHE��U>�"3?�B�>T�-�k�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*�F�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�\TS?N�R���W��#��*���p>
�������;ν���;�g��+��3�/�QG�?s_�? ��?��d�����?�]�>��I���TC���>Nڬ>b�&=9�$=��>r���;�#�X>���?�~�?�f(?�Vx�B�����g<�"w?�>���?(j�=ď�>��	>mq���K���/>��>,¸���?� N?���>��=�:5�Q./��ZA�d�L�O��A����>1<b?#J?ڱ]>y����� ��˽��.��̼�NA�.�)�&���'>+�H>��>�t=���ľ��?Np�7�ؿ j��p'��54?5��>�?����t�����;_?Gz�>�6��+���%���B�^��?�G�?<�?��׾�R̼�><�>�I�>1�Խ����V�����7>)�B?i��D��l�o�{�>���?�@�ծ?ki��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*i�̿抿�浾H����>���=_W>�\�w
i��e�=��<_�x�MR>��.>� �<�`�=�Iu<�ټ>L��>'|���>�F4���"��es;���>��M����3�����5��W�`�T�0��3a�)m��*1;��7ʩ=�X�=D�U?��Q?p?h� ?B�x�7�>4u��	8=#�Q��=C�>�[2?*�L?ݒ*?x�=����r�d�Vc��gC��1���}��>�jI>�a�>!N�>9�>-8X8r�I>?>���>�� >�Q'=Vx��sf
=eO>�W�>���>˚�>3G<>8�>zδ�*1��u�h��w�@=̽� �?<w����J�62��28��X���%\�=�e.?��> ���>п2�K0H?����?(�ߺ+�G�>X�0?�aW?��>���ѦT�76>!��^�j�rL>) ��|l��)��Q>�k?�$j>�h|>��3�l�8�k�K������"c>��9?Y/���yE�X^w���E�A׾�6>��>�SM<������~�x��h����=q?9?��?"��2h����q�� ���N>�`>��)=�}�=�;S>�	����Ľ��C�$Kl=$�=��Y>�[?��4>ו=`�>�k���I��>�yE>@1>g�A?@G'?Q<��+����Y~���.�i7p>c�>�j�>��=S�J��e�=�C�>�ta>�W�Fs��� �7�B�MS>�~���X�r�b���t=#&��$��=V�=K�(6�7�O=�~?���(䈿��e���lD?S+?] �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��L��=}�>׫>�ξ�L��?��Ž5Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l�6>�^%?��Ӿeh�>Bx�}Z�������u�H�#=@��>�8H?pV��e�O��>��v
?�?�^�ީ����ȿ(|v����>L�?���?Y�m��A���@����>6��?�gY?�oi>�g۾e`Z����>��@?�R?"�>�9���'�o�?�޶?���?�I>���?
�s?�r�>�x��Z/�4��T���"f=LK\;_�>_> ���iF�ד��g��&�j������a>N�$=j�>�M你2���#�=J��I����f����>54q>��I>K\�>Z� ? a�>���>�W=�p���䀾�����kP?zd�?͖��i��tb=g�u=� [�1?�+0?�@=WB��Mԭ>-�S?�5�?.Q?WB_>����Ԏ��ǿ�k��~o<�@>�>��>hꎽ��>>B�ҾAo*����>Ӯ�>\&=�E�ܮk�l��<v�>��?l~�>պ�=4�*?��%?M�n>7�>��g��u����&�>�>C�?��3?��?��+?�����.�]�������{*�_��>3�_?�_,?u��>m����t������} >��~��?T�@?)�b�z;?�vF?B�M?�wE?�!>���F����6�=W�=H� ?93�� �C��&���;��>���>n:�>�C�<���������\�ݾm��>C?h?bf/?�3���f�
7���(�<@9�;�?z�o�< y;���=�)>�{�f�=�*>���=�nM�PGV��fֹ��=F`�>�i2>�bH�$���/,,?�8B�!y���|�=��r�DoD�W�>
RK>q'��2�^?E�=�} |��'���o����T����?��?'_�?�д��h��<?�+�?g"?44�>�箾�ݾ�྆�w��Iw�����>���>��|��I�=���������~�ƽ�!�#��>���>!�#?v?��B>���>[�ξ� -��ԾO���D^�S�6�h�D��~&����,u��:��ٷ�'��������A�>,'����>g7?n��>U�Z>}��>4S <(�_>��>/!�>�\�>�v5>t� >�|p=���^�zPR?�����'���
����'B?�dd?I�>��h��|��ǵ�4v?B��?�s�?�.v>h�1&+��o?���>&���g
?�9=`�Z��<O��x��%������>T׽�:��M�h:f�r
?*?[:��X�̾��׽�ڟ��Wp=!B�?o�)?��)�#R�?�n���W��QR�K��0h�����s�$��p�gƏ��0�� ����v(��	)=ث*?�?
����"����j��t?�X�g>�C�>��>���>@nI>)	�u1�^��h'�܇���e�>]Y{?���>��Q?�<?��??�JN?�d�>mұ>OL��ٝ�>]��=;��>�>u-?��(?�?YF?��2?^
�>vp�H� �5�Ծ	� ?�]?B�?@�?�5?"I��rν�^.��;�X%��9�T�F=����s���˺y>�=�r�>�w?���ڽ8�(�����k>�>7?K5�>_&�>^����b����<l�>Ζ
?Ǐ>s���f}r�o'�-Q�>�7�?���M�=o>*>4W�=
����غN�=5�ż�t�=V���_&;���"<
�=��=�<~�I��9�;��;[�<�b�>�n?���>��?� �4��{0��kX�+/%>y�|>�%���b��h���L���HR��9>E��?`�?P.�;�x>9��=�׵�Z\���"�&྘�?��/
?"�:?�^?�Q�?�GV?RF?�4>.��>��R8k�'H����?v!,?��>�����ʾ��։3�؝?e[?�<a����;)��¾'�Խѱ>�[/�c/~����<D�U���]��5��?쿝?%A�R�6��x�ڿ���[��}�C?�!�>Y�>��>V�)�~�g�s%��1;>���>gR?I$�>��O?d7{?S�[?�aT>Y�8��1���љ���2���!>@?K��?`�?7y?F}�>��>k�)����M��\��D��₾W=�Z>k��>'*�>ީ>���=4Ƚ/N��-�>�+0�=ʖb>���>���>9�>iww>>d�<�B?Mz�>�;����v���r��y��WЀ?s��?�?��Y�~�/�
����>Cū?��?��?
S�w��=�<&���JO?�	�>nט>�s�>U�=�K)=�0>?�>��>�ܽ���ޅ,��B���?�8?�4�=��̿5~�ܢ߾)�
�Y�4>��^��@F>�F�<�����������[[��P�0Č��\����{���4���_N=(��>������>`N�=4����r>��S=�s��t�<g�%��V���Mu��=i\�=��l<F*�=$�@= �S�I��f*˾"�}?*I?t+?K�C?g�y>�Q>�2����>�����_?�}V>o�P� F��^�;������̔�P]ؾ��׾<%d�	����	>NI�B�>�o3>Bm�=%��<ѝ�=�r=��=p�;�v5=��=�y�=�̬=���=�K>�>�6w?X�������4Q��Z罤�:?�8�>^{�=��ƾo@?|�>>�2������wb��-?���?�T�?>�?@ti��d�>J���㎽�q�=@����=2>g��=u�2�R��>��J>���K��;����4�?��@��??�ዿТϿ4a/>�~x>��)>�kY���/���"��a�7�V��k-?m�'�������>���=̰ɾ�އ�X=$k�=�s=��ν]uz�fJb=�x���-=.*C=�X�>��.>_��=��གྷ��=�_�=:��=��>��E�V���~��ڇx=T_>}�@>8>'>UL�>#]?0
0?�e?y��>��r�l�;��¾�/�>Xm�=Ԯ>ʿ�=VB>���>�6?��C?��J?�ׯ>$ʉ=%p�>o��>܍,�0�m����;h��1+S<��?�E�?�c�>�J�<�>>����&F=�}ɽ,�?��/?��?�&�>Jj��+�-)�T�/���a��~�<�ީ=k�b�޲����(�E��ڽG��=�d�>��>-/�>YnW>8�&>0�M>#�>�>���<�F=&r��FB=p��;qu="���
��<A۔��~�<�n =�-5���>�R>D<!r�Z�Y<-��< �=���>��>��>�=h����$1>���� M�sv�=����@�B�D]e�߉~���.���4�"E>��Z>�����ܑ��
?vQ[>��A>=$�?��t?g"#>8W�r@վ�����Sg���M�2�=�>4�=�/G;��y`���L�<�Ҿ^��>Yߎ>+�>��l>�,�J#?���w=��_b5�|�>�|�����)��9q�@������Ui�KNҺ�D?�F��&��=y"~?�I?^�?��>q��݆ؾ�:0>�H����=f�z*q�}i����?'?���>�쾨�D�q5̾����>x�H���O���D�0�� ��������>s諭��о�3��g�������B��r�@�>��O?W�?b�gT��XVO����i���W?(|g?�:�>k[?a?���'b��[��/�=S�n?��?9�?�1>:k�=�����U�>$	?D��?xّ?E t?�>A�{��>"�<P}">$����=u�
>*��=��=�&?O-?�l
?!Z����� �ﾽ�ﾳQ\�Q�<�n�=ԝ�>ɉ>�t>�z�=��n=탤=�~Z>[D�>J��>�b>�¡>F=�>�$ྔ�5�Z�8?	�5=S�>�\?�Y�>��wQ����+����=�d�Γ�����O�Z�.����L#���Ƚ��C={w�>Dѿϗ�?C��>�n(�q(?{|�8��&�>�%!=/n�% �>��7>ty�>��>�W�>�ּ=X��>�d�=�4ԾYt>�����!���B�oR��JѾ�0z>i=��^�%��v�����*I����}��;j�wA��M�<�\�<�ۏ?������k��)����1?xb�>�6?�l��N~���>�`�>��>�0���s���Ѝ�a��C݋?���?�9>�`>�z?�j4?�;�Wi	�~M�"s��u�-�JQe�k�V����F7h��K���D���:b?��x?^�G?�@:=���>�:�?/9�����)՜>�js��qD�9��<I>Ru�����S����=o[�>�f�?7�Y?��>ڤ���Il�7_'>�:?1?OUt?��1?�|;?(T���$?	�3>W?�x?^A5?��.?��
?��1>f9�=�^��n	&=Tb��̊���нnBʽ�t��Z4=x|=��u���	<%]=���<�e�hyټ[f;N����?�<:=�'�=���=�N�>�`?�G�>�6�>�1$?�k���2A��b:��%?䞇��dɾQǾ���|o���>i�y?T��?�?k�>�9���%�V7<>=o�>M��=x˓>�>����aN�����=?#�=�N�=�NU=̉O<�_~�$�b�����=� �=_/�>|��>���Ո�>�Ê��ǰ��~�=5K���O��r�����>�Q�:�1��U?�>�HI?#?��><<�,��<�nF����>�X?)3`?<c?4W
>��Y=��Q�/�X�@;q> %P>hY����:�����s��TpX�>��=T�>H���ޠ��Ub>���s޾5�n��J����6HM=���YV=F�t�վF4� ��=�#
>θ��j� ����I֪��0J?ڥj=�v��z`U��n����>��>�ޮ>�:���v���@������2�=Ҷ�>� ;>_������~G�48���>-�F?�h?�?��_�!,d��A*���X҆��$q=��?5a�>+��>�>W7=7�Ǿ����X���2���>8��>(��O6�2mľ���PV.�S��>;�?���>��?�lO?�?�fP?�?�"�>g+�>=�3�,g��ѳ*?�%{?�̇��:����ă7���r�rj�>��>SX־u��n�>B4;?$m=?�׉?!K?  ��lw��n��-u>�6�>��H������q>T99?�?��l?�A�?�IW>3�!�M���l�L�t�_�"=�,?�j7?��?�OM>œ�>E���.��=n��>	c?�0�?a�o?[Z�=��?52>A��>�Җ=n��>I��>�?�PO?;�s?��J?��>i��<S0������1s���N��ք;�rJ<Ӽy=���u&t�J��l�<�O�;!�������3�IE�T0���n�;��>�qv>���X->�þ�͉��A=>i#���G��嗍��A���=V}�>�s?L��>,��0B�=ʥ�>�<�>�m���'?K6?W�?�]ʺίa�y�վ4E�@>�>%�A?��=>m������xv��J=�0l?K$`?��N����Q
r?��m?���K'-�����i־t�۾��|?:�>r���S�>���?4$�?�?�>��]�wk������\��*��� �=|E�>��!���f�%��>�=8?kl�>N{�>��5�/+����.˲��t�>�E�?9j�?�w?:L�=0z�I�W|ھ�0���FL?md%?�� ���D?O���:�������W~��������~�1���?�H�ǭ��(c(�Ϊn�:c$���P=w?�Yy?�w?v\V?�v�m��i�j���q��^��
�w��IX��6�ި2��XR�F���y���fሾ��>|�q���=��;�?8,?O2��B�>_G���s�����>�A>�o��������=����4h�<˄�<>Br�~ 8�9~����!?���>�>J�>?��a���>���5�̖7�ڭ�·@>��>�%�>ۭ�>T:�;��/���޽�����y�.C���8v>�xc?ԏK?�n?k�'*1�m���7�!���/�b����B>Sl>���>|�W����.:&�Y>��r����8v����	��~=߯2?�'�>ݲ�>O�?3?@{	�	g���ex��1����<o0�>i?�=�>��>�нR� ���>v�l?�U�>�S�>�A��f(!�y$x�;MϽ�^�>uK�>��>Zon>��7�B%]���������_�7��[�=/�f?)H��:a���>��O?��e<�}�<�ƣ>�y�_*#�����>�8	?�H�=�7>��ɾ���(�{����sP)?7L?�璾�*�d:~>;#"?��>	0�>�0�? *�>YqþDD�R�?��^?"BJ?GSA? F�>��=���M?Ƚ@�&��,=��>%�Z>a+m=b��=���2n\��r���D=�u�=�μX���<�p���K<D��<��3>&mۿ�BK�}�پ�
��� ?
�z爾E����c�����/a������Xx���('��V��5c�����p�l����?�=�?P����/��ղ������������>�q�����������5)�����ӿ��Bd!��O��&i�<�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >ZC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾x1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@}A?��(�,���V=���>�	?��?>�S1�&I�	����T�>`<�?���?-{M=5�W���	��e?/j<�F���ݻ��=I>�=�I=[��;�J>�U�>ك�SA��<ܽ��4>�څ>K"����/�^�'��<7�]>��ս�7��0Մ?�z\��f���/��T���T>��T?/+�>�9�=Q�,?|7H�R}Ͽ�\��*a?�0�?���?�(?1ۿ��ؚ>|�ܾ�M?MD6?���>�d&� �t����=3��k��/�㾶&V�Y��=ӫ�>��>��,���^�O� C����=P�#��c�=���0��g�<&#>��!=��o������<��+����ё��v�_�ؽ]��=��?2��>0;�>u�8?��<?���>��>�=������䶾-��B~���k���m�\X;��E\����������[��ڇ
�j6J�^��� =���=�7R������� ���b�v�F���.?At$>M�ʾ��M�v�-<znʾ0��������ԥ�|+̾�1��n�0̟?7�A?����k�V�+���R��r��įW?I�'��T묾C��=�ݱ��=� �>��=���=3��}S��0?��?�#�������%>?��L8=�E,?�?k��;�q�>D"?b&/�X8罅�]>�39>�/�>��>��>K�����ٽI&? �T?}��蜾�=�>)���&s�V=r�>�~5�"��V>H��;	x��=��������<j(W?웍>+�)����`���]==>�x?Ȓ?�-�>{k?��B?KƤ<�h��k�S����`w=a�W?�)i?ֹ>�����оr�����5?�e?�N>]bh������.��T��$?E�n?�^?B���Jw}��������n6?V�v?|s^��s�����c�V�>�>"\�>T��>R�9��k�>O�>?�#�~G�������Y4�&?W�@���?�#<<��⛎=�;?D\�>A�O�x;ƾ��������m�q=��>≧��cv����@U,��8?���?���>�������t�=@��`U�?8=�?����:m<���Ql������ܘ<�I�=#n�)j&��B�g�7�a6ƾ�X
�7���㙺�,�>6_@�?�y�>�g8��f⿨6Ͽs�Ѿ)�q�<<?�ݨ>��ƽqZ��I�i��t�(.G�NlH�ц��U`�>��>G���󏑾�|�b�;�h0���_�>Ek��Z�>�]T�PǶ��x����M<�"�>�>�>����ݎ�����?Р��^?ο�����_��_X?�0�?m\�?��?*�)<;w�9~{�F���pG?��s?�5Z?�c)��]��6�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�znT?��"��f?�¿��3����<g�!�پ����x����v������Y�;���?%��?.�?p���_G&��+?��>�h�@��9}��?]l�>�M߼n?�=;�/=w����>�2)�>�0�?'�?�V?�w4�ݮ�|�V=-�u?)q�>���?��>���>�>�:���<<��<>#>���3?��I?���>���=��1��?-�P�H���S��M�^�?�On>�e?�Q?��Y>���*��&�=����N�)��<�P�2?]��F����>K�J>Et(>�5,�W��	V?�����ؿ�x��C�'�O�3?�T�>��?c9��r�Ll��h�^?�ц>�^�e���O����������?�(�?��?�H׾B�ļ5 >�;�>�,�>�ԽX���ň�L�4>JQB?}c����?yo����>�u�?mo@�O�?P�h���?�&�%T��yd~���&�6����=N�7?�#��z>0��>�5�=unv����c�s���>PB�? �?R��>�l?qxo��B��(2=�P�>��k?�l?�-s��f�B>�?��������K�f?��
@�p@P�^?U좿!&ʿ\G��A���+�Q �W�g<��P>�Ľ�.>�wh>A�_>fPۻe:>�O>��>�R> ��>�#�>���>w����M�2ٱ�rӡ�6kR���!�Dy
�<*�"(�P	����,ʾ'��R@�Œ�xQi�b����=�x�=O�O>�R?�`?[�j?�1?j&��=Q>�Ҿ$>do,�E(>8��>s�*?��6??Z?I1�<>����c��c��/]����J�?>�>�S�>Z�>�>X6�z�D>+:>
g�>��}>�w\��Sټ�m0��Ch>��>q�>p�>�^<>��>�̴�.���h��w�to̽d��?���v�J��6���;�������v�=�s.?�>O���:п�ꭿd'H?L씾�%���+��>ջ0?ZuW?7�>�۰�a~T�F=>�����j�G>�s �ӗl�Tk)�6hQ>$V?��f>�1u>��3��d8�}�P�?~���M|>�56?�eh9�5�u���H�~Mݾ�FM>R۾>�=A�Sk�����	�Yti�a�{=er:?B�?y^��vذ��fu�9,���R>�C\>v�=�,�=l(M>2 d��&ǽ�H�k/=�=!�^>SO?38->��=i�>�e��X�O�S�>ݰ?>�,>�??��$?��>똽������.���t>�,�>�1�>�>#I�}�=�!�>�4b>��&���H���A�drX>ul��\�C}p��1�=�|��K2�=[3�=P��� �:��+=��~?�`��&݈��׵��9D?��?XO�=85<��"����h<����?��@u��?�-	�Q�V�G�?�B�?락J�=�>�>��>ޫ;�=L���?��Ľf����u	��Z#�UO�?v�?�w3�����o�k�;>L>%?ӐӾIh�>�x��Z�������u�l�#=R��>�8H?�V����O�_>��v
?�?�^�ߩ����ȿ2|v����>X�?���?g�m��A���@����>:��?�gY?voi>�g۾?`Z����>ѻ@?�R?�>�9��'���?�޶?֯�?e�J>�K�?+t?���>;�e���-���������m�~=O�;�>~F>G��E3F��H��?��4sj�h���`>��/=]q�>*�����%��=9�������{��D�>�f}>�O>���>8�?���>�ԗ>��=�s����y�����u�W?��?����Y�pYx>�ҼT̽ʚ:?
�!?�T=aSξ�b�>o�d?�i?ʞ??�B�=?�"�vA��2aο̗��F~�MR�>��>T��>�һ=滍>b���܏��/�><��>F7��\>����~���'����>O�?t+�>#���4(?�0?a�>��>�<@����'x6�k�>w��>*)-?�ۀ?vM'?j�f�U�1�W��%��ՙL��A>�i?�T#?�w�>���ta��C�Y�3�U�ɮC�V��?�?N?�
�t?�܄?1�W?[)4?�E>��d��ӾQ.��[�>["?tw�x�A��&��� �fn?N��>ߴ�>��ν�0��8a�z'�-��ye?�c?S�+?�	�yZa�/t��
��<�s���*�N���Y��>==2>~�;��`�=�>n?�=�ge�a�@�������=� �>���=SP6�*����#,?\[8=�#��+�=�$q�_�F�ס|>c`L>�l����H?�1h�N������yV����O�Փ�?���?v�?��׽�Pb���/?�O�?�?���>\���w�� .���e\�; ����]�3>�[�>����v]�;묿-���ˇ��Mh���"���>�^�>eM	?آ?��P>s��>?֚�R��X[�H4��[��y���9��-�%��Ꝿ�*���@�����v����>�Ր���>��?sr>˝q>���>�UX<���>&�^>�b�>f�>�N>��>�=�vֻ�H���KR?����$�'����󰰾2B?Tod?]0�>�,i�i�������?ۆ�?ys�?;Dv>�|h��-+�>m??�>��� q
?�N:=�b��T�<�T�����:,����C��>hG׽�:�}M��rf�j
?0/?F����̾3>׽���� �=(��?ݣ)?��'��pP�9�l�eY���P�Vh�ʀe�����#���o��7��C:��񯃿��'���/=h*?�Y�?���,���᰾˶l��?�&Nc>���>�ל>;�>��L>j��50�!�\�QC'�X���Uk�>g�z?�>�pI?�<?��P?o�L?�ώ>_��>�鯾��>)s<���>e��>)o9?Ө-?��/?
?��*?�<a>��������H�ؾ m?f�?��?�^?��?�z����ý૙���>���v���3�={8�<#�ֽ�o�}X=�aV>�X?X��]�8�)����k>n�7?_��>��>����,����<��>��
?`F�>A �~r�c�7V�>m��? ����=��)>���=r���l�ҺCY�=N�����= *���x;��o<��=���=
Nt�恹�$�:���;�r�<'��>��?�n�>���>����@����w˰=A�^>�7N>��>�/ܾ�������w�f�[Zz>6��?x��?��\=�`�=���=����S켾_9��¼���=��?�"?zU?�ђ?I2>?�!?���=���;��O���>٦�|{?{!,?5��>n��x�ʾ�񨿿�3�ܝ?f[?`<a�����;)���¾s�Խ��>�[/�T/~����BD��
��������+��?꿝?�A�7�6��x�ٿ���[����C?P"�>5Y�>b�>K�)�w�g�V%��1;>��>nR?�!�>�vO?*w?�`X?��W>��8�ΐ�����K�u�>��9?%P�?���?�v{?���>]->N(8��q�Q���'<��*���/=��c>'|�>���>c�>�m�=ˋ�������_3����=wsM>mD�>���>a��>"q>�˧<��D?"6?z�Z��jȝ�󢾟>v�D��?M�?(��>��_�l6+��-��r���>v�?e�?#'?�g>�W��=i?<�W��ن���$>Q��>�-�>9��<4:�>�;�>\�>1�P>��Ծ!���Fj������fA?��Q?�4�����͜x��<ӾL�����=�H�<�e>V�M�IĽ�B~>?%������X
���Ծ転�J�ٽ�<>(�	=��>�"=��o=}>&rn>@� >{B>�I�=�X�[&&=􅰽�������$��([���u½M���Y�>§=(m�.k?	�p?C1?�E?^��>���>�ֽ>��	�?�޵>qͻ��"ľ�X�#:��ۧ��=��w�پ��/�������->��=�-�<2a>L�=�W
�F}>=�t>�@=2�K<���=�>��>Vl6���=��w>o[>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>Hj5>.C>��R���1�n%\�aJa��Y��e!?�;���˾ģ�>m�=��߾<Ǿ5G)=��5>��h=����[��s�=��y�݊?=�+p=��>B3D>W�=�q���{�=�oG=�=�= �N>�����~5�3m+�A�1={��=r`>S�$>���>|�?z,?U�`?���>�p�[(Ҿ ���P��>>W�=��>A�}=KI>�T�>Z9;?�F?��H?7Ĭ>���=8ȸ>�:�>f�+�Xdk�#��찥���%=C$�?a��?���>O�o<�G����n�@��߽�u?�4?{
?��>�s�m7߿�w&���-�)딽X<��L=c�q�ݪM��ҼV�����K�=���>��>�ޛ>�]�>�E>5T>�Ӿ>��>]��<��=!��;���<�&���V�=8.��t\�<�!�&�~���4�p3��X�v���	��US<�^�;�
�=���>��1>�6�>�q�=�y���XE>����Y?�ݏ�=�����:�.ri����l.���8�k09>�.>o�v�b����>i�v>�l,>��?o�u?E�0>ƹ����؁��{�9��"��Y	>���=�?�K�A��k���P��]��c��>qߎ>=�>��l>�,�F#?���w=��=b5�d�>�|������)��9q�@������`i��Һ�D?�F��1��=p"~?�I?a�?���>���φؾ�:0>�H��V�=<��)q��h����?�'?���>�쾄�D�Mm̾}�����>��I�� P�۽���0����������>Pت�f�о�3�>e������ �B�r�E�>�O?��?rIb�	Z��JO�������o?lzg?��>�=?*?�����x��,�=��n?���?�=�?	>���=C;�����>B�?궖?sؑ?+�s?�j@�J��>W�<��!>�V��_��=�>���=�=�9?�Q
?
B
?�ؘ�!\	����C�* _�� =�.�=�̐>���>Us>��=��u=Bi�=(r^>ì�>'o�>�d>�U�>겉>>g̾��$�R?TK>���>=�^?��>8dS�Ō=�Կ=�W=���}3v��>7�mHG��&���3���=��:V'?"�����x?Y��>�@�U�
?)�#�����ݷ> 砽���N<?鞇>��>�C�><٭>�0,>oi�=?@�=EGӾM~>����d!��,C��R���Ѿ	}z>"����&�q��`w���BI��n��xg�Pj�.���;=�yֽ<�G�?����k���)�������?s[�>�6?�ٌ��	��;�>���>�Ǎ>�J��E���6ȍ��gᾰ�?��?E�f>B$d>Eij?�+6?ib����=�J�c�Q���a�7��e�(�Y�ޔ�[�|���Ѿ�q���`?)r?z�&?`J�=�)�>_W�?��s=Ͼg�>%�k�v�E�� ;`m<�8澶5��������H�=��>.�?��n?��?�)����en)>�6F?��5?��p?�6?�??xN�("$?>�A>f7?�U?r�/?ٽ)?j?�$>J�=���8W<3Ė����Ѹ������1�-c=���=�0��klݻ�	`=�x�;����������;9^��@�;ӡ�< ��=��>ߔ�>3�]?/a�>%��>Z%6?�d��Y7�$_���/?AP'=�������[-��'N򾃐>��j?x3�?A�Y?Q�a>��B��nB�_&!>=T�>�0&>z�Z>�W�>֙��B���=l:>�@>�$�=9 Y�xz�����pr��.�<�>�7�>^
�>c6����>�Z����vL>P%6������w���N���1���f�W��>,�Q?Ɍ$?�Ҟ=�J龾烽�0a�g&?�8?2J?��s?�'�=�G��"l/��1:�?�SI�>��<�Oe�>���ˣ��=�7L=�م>|���ޠ��Ub>���s޾5�n��J����6HM=���YV=F�t�վF4� ��=�#
>θ��j� ����I֪��0J?ڥj=�v��z`U��n����>��>�ޮ>�:���v���@������2�=Ҷ�>� ;>_������~G�48���>-�F?�h?�?��_�!,d��A*���X҆��$q=��?5a�>+��>�>W7=7�Ǿ����X���2���>8��>(��O6�2mľ���PV.�S��>;�?���>��?�lO?�?�fP?�?�"�>g+�>=�3�,g��ѳ*?�%{?�̇��:����ă7���r�rj�>��>SX־u��n�>B4;?$m=?�׉?!K?  ��lw��n��-u>�6�>��H������q>T99?�?��l?�A�?�IW>3�!�M���l�L�t�_�"=�,?�j7?��?�OM>œ�>E���.��=n��>	c?�0�?a�o?[Z�=��?52>A��>�Җ=n��>I��>�?�PO?;�s?��J?��>i��<S0������1s���N��ք;�rJ<Ӽy=���u&t�J��l�<�O�;!�������3�IE�T0���n�;��>�qv>���X->�þ�͉��A=>i#���G��嗍��A���=V}�>�s?L��>,��0B�=ʥ�>�<�>�m���'?K6?W�?�]ʺίa�y�վ4E�@>�>%�A?��=>m������xv��J=�0l?K$`?��N����Q
r?��m?���K'-�����i־t�۾��|?:�>r���S�>���?4$�?�?�>��]�wk������\��*��� �=|E�>��!���f�%��>�=8?kl�>N{�>��5�/+����.˲��t�>�E�?9j�?�w?:L�=0z�I�W|ھ�0���FL?md%?�� ���D?O���:�������W~��������~�1���?�H�ǭ��(c(�Ϊn�:c$���P=w?�Yy?�w?v\V?�v�m��i�j���q��^��
�w��IX��6�ި2��XR�F���y���fሾ��>|�q���=��;�?8,?O2��B�>_G���s�����>�A>�o��������=����4h�<˄�<>Br�~ 8�9~����!?���>�>J�>?��a���>���5�̖7�ڭ�·@>��>�%�>ۭ�>T:�;��/���޽�����y�.C���8v>�xc?ԏK?�n?k�'*1�m���7�!���/�b����B>Sl>���>|�W����.:&�Y>��r����8v����	��~=߯2?�'�>ݲ�>O�?3?@{	�	g���ex��1����<o0�>i?�=�>��>�нR� ���>v�l?�U�>�S�>�A��f(!�y$x�;MϽ�^�>uK�>��>Zon>��7�B%]���������_�7��[�=/�f?)H��:a���>��O?��e<�}�<�ƣ>�y�_*#�����>�8	?�H�=�7>��ɾ���(�{����sP)?7L?�璾�*�d:~>;#"?��>	0�>�0�? *�>YqþDD�R�?��^?"BJ?GSA? F�>��=���M?Ƚ@�&��,=��>%�Z>a+m=b��=���2n\��r���D=�u�=�μX���<�p���K<D��<��3>&mۿ�BK�}�پ�
��� ?
�z爾E����c�����/a������Xx���('��V��5c�����p�l����?�=�?P����/��ղ������������>�q�����������5)�����ӿ��Bd!��O��&i�<�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >ZC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾x1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@}A?��(�,���V=���>�	?��?>�S1�&I�	����T�>`<�?���?-{M=5�W���	��e?/j<�F���ݻ��=I>�=�I=[��;�J>�U�>ك�SA��<ܽ��4>�څ>K"����/�^�'��<7�]>��ս�7��0Մ?�z\��f���/��T���T>��T?/+�>�9�=Q�,?|7H�R}Ͽ�\��*a?�0�?���?�(?1ۿ��ؚ>|�ܾ�M?MD6?���>�d&� �t����=3��k��/�㾶&V�Y��=ӫ�>��>��,���^�O� C����=P�#��c�=���0��g�<&#>��!=��o������<��+����ё��v�_�ؽ]��=��?2��>0;�>u�8?��<?���>��>�=������䶾-��B~���k���m�\X;��E\����������[��ڇ
�j6J�^��� =���=�7R������� ���b�v�F���.?At$>M�ʾ��M�v�-<znʾ0��������ԥ�|+̾�1��n�0̟?7�A?����k�V�+���R��r��įW?I�'��T묾C��=�ݱ��=� �>��=���=3��}S��0?��?�#�������%>?��L8=�E,?�?k��;�q�>D"?b&/�X8罅�]>�39>�/�>��>��>K�����ٽI&? �T?}��蜾�=�>)���&s�V=r�>�~5�"��V>H��;	x��=��������<j(W?웍>+�)����`���]==>�x?Ȓ?�-�>{k?��B?KƤ<�h��k�S����`w=a�W?�)i?ֹ>�����оr�����5?�e?�N>]bh������.��T��$?E�n?�^?B���Jw}��������n6?V�v?|s^��s�����c�V�>�>"\�>T��>R�9��k�>O�>?�#�~G�������Y4�&?W�@���?�#<<��⛎=�;?D\�>A�O�x;ƾ��������m�q=��>≧��cv����@U,��8?���?���>�������t�=@��`U�?8=�?����:m<���Ql������ܘ<�I�=#n�)j&��B�g�7�a6ƾ�X
�7���㙺�,�>6_@�?�y�>�g8��f⿨6Ͽs�Ѿ)�q�<<?�ݨ>��ƽqZ��I�i��t�(.G�NlH�ц��U`�>��>G���󏑾�|�b�;�h0���_�>Ek��Z�>�]T�PǶ��x����M<�"�>�>�>����ݎ�����?Р��^?ο�����_��_X?�0�?m\�?��?*�)<;w�9~{�F���pG?��s?�5Z?�c)��]��6�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�znT?��"��f?�¿��3����<g�!�پ����x����v������Y�;���?%��?.�?p���_G&��+?��>�h�@��9}��?]l�>�M߼n?�=;�/=w����>�2)�>�0�?'�?�V?�w4�ݮ�|�V=-�u?)q�>���?��>���>�>�:���<<��<>#>���3?��I?���>���=��1��?-�P�H���S��M�^�?�On>�e?�Q?��Y>���*��&�=����N�)��<�P�2?]��F����>K�J>Et(>�5,�W��	V?�����ؿ�x��C�'�O�3?�T�>��?c9��r�Ll��h�^?�ц>�^�e���O����������?�(�?��?�H׾B�ļ5 >�;�>�,�>�ԽX���ň�L�4>JQB?}c����?yo����>�u�?mo@�O�?P�h���?�&�%T��yd~���&�6����=N�7?�#��z>0��>�5�=unv����c�s���>PB�? �?R��>�l?qxo��B��(2=�P�>��k?�l?�-s��f�B>�?��������K�f?��
@�p@P�^?U좿!&ʿ\G��A���+�Q �W�g<��P>�Ľ�.>�wh>A�_>fPۻe:>�O>��>�R> ��>�#�>���>w����M�2ٱ�rӡ�6kR���!�Dy
�<*�"(�P	����,ʾ'��R@�Œ�xQi�b����=�x�=O�O>�R?�`?[�j?�1?j&��=Q>�Ҿ$>do,�E(>8��>s�*?��6??Z?I1�<>����c��c��/]����J�?>�>�S�>Z�>�>X6�z�D>+:>
g�>��}>�w\��Sټ�m0��Ch>��>q�>p�>�^<>��>�̴�.���h��w�to̽d��?���v�J��6���;�������v�=�s.?�>O���:п�ꭿd'H?L씾�%���+��>ջ0?ZuW?7�>�۰�a~T�F=>�����j�G>�s �ӗl�Tk)�6hQ>$V?��f>�1u>��3��d8�}�P�?~���M|>�56?�eh9�5�u���H�~Mݾ�FM>R۾>�=A�Sk�����	�Yti�a�{=er:?B�?y^��vذ��fu�9,���R>�C\>v�=�,�=l(M>2 d��&ǽ�H�k/=�=!�^>SO?38->��=i�>�e��X�O�S�>ݰ?>�,>�??��$?��>똽������.���t>�,�>�1�>�>#I�}�=�!�>�4b>��&���H���A�drX>ul��\�C}p��1�=�|��K2�=[3�=P��� �:��+=��~?�`��&݈��׵��9D?��?XO�=85<��"����h<����?��@u��?�-	�Q�V�G�?�B�?락J�=�>�>��>ޫ;�=L���?��Ľf����u	��Z#�UO�?v�?�w3�����o�k�;>L>%?ӐӾIh�>�x��Z�������u�l�#=R��>�8H?�V����O�_>��v
?�?�^�ߩ����ȿ2|v����>X�?���?g�m��A���@����>:��?�gY?voi>�g۾?`Z����>ѻ@?�R?�>�9��'���?�޶?֯�?e�J>�K�?+t?���>;�e���-���������m�~=O�;�>~F>G��E3F��H��?��4sj�h���`>��/=]q�>*�����%��=9�������{��D�>�f}>�O>���>8�?���>�ԗ>��=�s����y�����u�W?��?����Y�pYx>�ҼT̽ʚ:?
�!?�T=aSξ�b�>o�d?�i?ʞ??�B�=?�"�vA��2aο̗��F~�MR�>��>T��>�һ=滍>b���܏��/�><��>F7��\>����~���'����>O�?t+�>#���4(?�0?a�>��>�<@����'x6�k�>w��>*)-?�ۀ?vM'?j�f�U�1�W��%��ՙL��A>�i?�T#?�w�>���ta��C�Y�3�U�ɮC�V��?�?N?�
�t?�܄?1�W?[)4?�E>��d��ӾQ.��[�>["?tw�x�A��&��� �fn?N��>ߴ�>��ν�0��8a�z'�-��ye?�c?S�+?�	�yZa�/t��
��<�s���*�N���Y��>==2>~�;��`�=�>n?�=�ge�a�@�������=� �>���=SP6�*����#,?\[8=�#��+�=�$q�_�F�ס|>c`L>�l����H?�1h�N������yV����O�Փ�?���?v�?��׽�Pb���/?�O�?�?���>\���w�� .���e\�; ����]�3>�[�>����v]�;묿-���ˇ��Mh���"���>�^�>eM	?آ?��P>s��>?֚�R��X[�H4��[��y���9��-�%��Ꝿ�*���@�����v����>�Ր���>��?sr>˝q>���>�UX<���>&�^>�b�>f�>�N>��>�=�vֻ�H���KR?����$�'����󰰾2B?Tod?]0�>�,i�i�������?ۆ�?ys�?;Dv>�|h��-+�>m??�>��� q
?�N:=�b��T�<�T�����:,����C��>hG׽�:�}M��rf�j
?0/?F����̾3>׽���� �=(��?ݣ)?��'��pP�9�l�eY���P�Vh�ʀe�����#���o��7��C:��񯃿��'���/=h*?�Y�?���,���᰾˶l��?�&Nc>���>�ל>;�>��L>j��50�!�\�QC'�X���Uk�>g�z?�>�pI?�<?��P?o�L?�ώ>_��>�鯾��>)s<���>e��>)o9?Ө-?��/?
?��*?�<a>��������H�ؾ m?f�?��?�^?��?�z����ý૙���>���v���3�={8�<#�ֽ�o�}X=�aV>�X?X��]�8�)����k>n�7?_��>��>����,����<��>��
?`F�>A �~r�c�7V�>m��? ����=��)>���=r���l�ҺCY�=N�����= *���x;��o<��=���=
Nt�恹�$�:���;�r�<'��>��?�n�>���>����@����w˰=A�^>�7N>��>�/ܾ�������w�f�[Zz>6��?x��?��\=�`�=���=����S켾_9��¼���=��?�"?zU?�ђ?I2>?�!?���=���;��O���>٦�|{?{!,?5��>n��x�ʾ�񨿿�3�ܝ?f[?`<a�����;)���¾s�Խ��>�[/�T/~����BD��
��������+��?꿝?�A�7�6��x�ٿ���[����C?P"�>5Y�>b�>K�)�w�g�V%��1;>��>nR?�!�>�vO?*w?�`X?��W>��8�ΐ�����K�u�>��9?%P�?���?�v{?���>]->N(8��q�Q���'<��*���/=��c>'|�>���>c�>�m�=ˋ�������_3����=wsM>mD�>���>a��>"q>�˧<��D?"6?z�Z��jȝ�󢾟>v�D��?M�?(��>��_�l6+��-��r���>v�?e�?#'?�g>�W��=i?<�W��ن���$>Q��>�-�>9��<4:�>�;�>\�>1�P>��Ծ!���Fj������fA?��Q?�4�����͜x��<ӾL�����=�H�<�e>V�M�IĽ�B~>?%������X
���Ծ転�J�ٽ�<>(�	=��>�"=��o=}>&rn>@� >{B>�I�=�X�[&&=􅰽�������$��([���u½M���Y�>§=(m�.k?	�p?C1?�E?^��>���>�ֽ>��	�?�޵>qͻ��"ľ�X�#:��ۧ��=��w�پ��/�������->��=�-�<2a>L�=�W
�F}>=�t>�@=2�K<���=�>��>Vl6���=��w>o[>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>Hj5>.C>��R���1�n%\�aJa��Y��e!?�;���˾ģ�>m�=��߾<Ǿ5G)=��5>��h=����[��s�=��y�݊?=�+p=��>B3D>W�=�q���{�=�oG=�=�= �N>�����~5�3m+�A�1={��=r`>S�$>���>|�?z,?U�`?���>�p�[(Ҿ ���P��>>W�=��>A�}=KI>�T�>Z9;?�F?��H?7Ĭ>���=8ȸ>�:�>f�+�Xdk�#��찥���%=C$�?a��?���>O�o<�G����n�@��߽�u?�4?{
?��>�s�m7߿�w&���-�)딽X<��L=c�q�ݪM��ҼV�����K�=���>��>�ޛ>�]�>�E>5T>�Ӿ>��>]��<��=!��;���<�&���V�=8.��t\�<�!�&�~���4�p3��X�v���	��US<�^�;�
�=���>��1>�6�>�q�=�y���XE>����Y?�ݏ�=�����:�.ri����l.���8�k09>�.>o�v�b����>i�v>�l,>��?o�u?E�0>ƹ����؁��{�9��"��Y	>���=�?�K�A��k���P��]��c��>qߎ>=�>��l>�,�F#?���w=��=b5�d�>�|������)��9q�@������`i��Һ�D?�F��1��=p"~?�I?a�?���>���φؾ�:0>�H��V�=<��)q��h����?�'?���>�쾄�D�Mm̾}�����>��I�� P�۽���0����������>Pت�f�о�3�>e������ �B�r�E�>�O?��?rIb�	Z��JO�������o?lzg?��>�=?*?�����x��,�=��n?���?�=�?	>���=C;�����>B�?궖?sؑ?+�s?�j@�J��>W�<��!>�V��_��=�>���=�=�9?�Q
?
B
?�ؘ�!\	����C�* _�� =�.�=�̐>���>Us>��=��u=Bi�=(r^>ì�>'o�>�d>�U�>겉>>g̾��$�R?TK>���>=�^?��>8dS�Ō=�Կ=�W=���}3v��>7�mHG��&���3���=��:V'?"�����x?Y��>�@�U�
?)�#�����ݷ> 砽���N<?鞇>��>�C�><٭>�0,>oi�=?@�=EGӾM~>����d!��,C��R���Ѿ	}z>"����&�q��`w���BI��n��xg�Pj�.���;=�yֽ<�G�?����k���)�������?s[�>�6?�ٌ��	��;�>���>�Ǎ>�J��E���6ȍ��gᾰ�?��?E�f>B$d>Eij?�+6?ib����=�J�c�Q���a�7��e�(�Y�ޔ�[�|���Ѿ�q���`?)r?z�&?`J�=�)�>_W�?��s=Ͼg�>%�k�v�E�� ;`m<�8澶5��������H�=��>.�?��n?��?�)����en)>�6F?��5?��p?�6?�??xN�("$?>�A>f7?�U?r�/?ٽ)?j?�$>J�=���8W<3Ė����Ѹ������1�-c=���=�0��klݻ�	`=�x�;����������;9^��@�;ӡ�< ��=��>ߔ�>3�]?/a�>%��>Z%6?�d��Y7�$_���/?AP'=�������[-��'N򾃐>��j?x3�?A�Y?Q�a>��B��nB�_&!>=T�>�0&>z�Z>�W�>֙��B���=l:>�@>�$�=9 Y�xz�����pr��.�<�>�7�>^
�>c6����>�Z����vL>P%6������w���N���1���f�W��>,�Q?Ɍ$?�Ҟ=�J龾烽�0a�g&?�8?2J?��s?�'�=�G��"l/��1:�?�SI�>��<�Oe�>���ˣ��=�7L=�م>|��oSp��x�>U}վ���{���A�K&�w�!>0�7����>��M��3!��.�\����V�'�|�D��ͦ� (���@?���=A˾i�ʾ!���I�>R�>�9?��<=���D`�J�~5~>H?� �>к:=Y���D��48�+�>b�E?�:d?z��?�ہ��1s��HB����ࠜ�pv��?�K�>��?,&I>���=T���%���P`�nWI�9f�>��>W���H�	៾���Z0�Ϧ�>��?�>��?�EV?!f?>?\?�'?�?��>X�`�����%L ?�-�?f,�=)�ý�HV���8�.E@�y��>.k)?/Qv��ĝ>�$"?I�,?�.&?]K?��?�3>8� B��̓>�>[Sb�3>����l>�J?�9�>�P?Z}?�>-�%�J*w�����>.H>�,?u4?��?=.�>��?)L��>ϖ?n/?��s?���?���>���>a��&޶>��=���#�>F��>al?���?��_?*�7?v鲼{��=�j�;2Xy�KC!>/�*�ڠZ�ߴ����g=�J�����r%g;[Щ��>`=�E�='��=z�ɽ�c����=%R�>��s>������0>�oľ^����A>�駼�W��Ғ��l�9�ȧ�=�y�>�?���>A@#����=�>�<�>�����'?�?�?G�;�nb���ھ8�K���>�0B?!e�=��l�����1�u��vh=��m?h^?F5W�I���
qb?�^?g��^�=��Hž�"c�����O?	?�/C��>-j}?l�q?ږ�> �g���n����"�b�m�l�=���>�n��6e��۝>�C8?�U�>�af>b��=��۾#x������?v$�?�?�׊?A<+>�n�I�	��������.]?�=�>������?G[�-ξ���������M�崧�����d���Ã���F��w�<�۽&��=Ɏ?��v?<�n?��_?0��xh�t�c��>y�q�]�E��?��%C���<��
D��$v��W����E��«�<�H��}�B�
�?x'?j?0��h�>Ӏ������ξqYE>�|������c�=k��T=�`=�oc�lD.��8���6 ?���>���>��<?*$Y��6?��,3��'6�[���L�,>Nǣ>���>/��>Ds���8�&���0̾0ʇ���߽:l>N�d?�dW?f�i?啽���8�����0+�2߽y޵���5>��>C �>/�*�?�%�'��	E��m�jX�|E��r"
�Lr1>��@?�Ճ>i�>�W�?Q?#������qu��u%�G��=W��>5N?�Բ>3�>��,���>��l?���>W�>����[!�f�{��ʽ�#�>�߭>���>&�o>��,�o#\��j��h���`9�Po�=�h?������`�W�>�R?3��:��G<|�>�v��!������'��>�|?���=��;>m�ž$$�1�{�^8��xW)??�?О��KH*��[}>g"?���>`��>��?o�>n�¾ď�c?��^?�J?0#A?�w�>�P!=]�����ǽ}D&��.=+��>�R[>��o=���=���\������C=�!�=�VӼ������<����<�T<��<=y5>LWۿ��K��%پM��$s��
��L���\������@��,��[U��3�y�\/��^�8�U�9�_�����p4i�)��?_��?�z��Fꉾa���,5��v���"�>�y������ޫ��P��[��-G��԰�Y�!�ƦP���i�:f�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >^C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾u1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�>@?��$����W=��>��?ܦA>"�4��H��%��߮�>���?9��?Pjy=��V�7��c?X3L<̒D������=��=i�=Z3���^>��>���LqJ��.̽n}7>�}�>D�s��"��[]����<�"R>k�Խ�q�5Մ?-{\�yf���/��T��"U>��T?+�>Y:�=��,?Q7H�[}Ͽ�\��*a?�0�?��?)�(?"ۿ��ؚ>��ܾ��M?dD6?���>�d&��t�Å�=87�%�������&V�a��=V��>a�>Ă,�Ӌ�t�O�J�����=����@����=b�;=���*輹{ͼ��9���M���=%p��gnE�I3���۽I�l>43>�p�>��Y>���>�PW?uWU?�³>F��=Fǽ�]���ݾ.[�=!ȾW�d��T���T���9���x��G�
��Z�z_,��ʾH�<��=��Q�B���"X!���b��G�'�.?�� >�Ⱦu�N����;pɾ��4Y���q���{;nS2��Hn�{��?S�A?�兿n3W�c���4���SX?���8��������=DV��L�"=?�>+G�=|���3��S�hl0?l[?�}���R��^^*>� ��?=��+?;�?�FX<ZB�>a_%?��*�Pp��T[>�3>�ɣ>H��>M0	>�����۽��?V�T?�������Ӑ>ya��d�z��Sb=!r>�45�����q[>V'�<�ތ���W�������<W?Y��>��)�U���E���S��>=́x?R�?���>�nk?C?���<�����S���sax=�W?�i?L�>\j���%о}����5?��e?rhO>�5h���龺�.�;7��?��n?�\?�S��D}��������6?�v?�y^�Oi������V�WF�>ӆ�>� �>��9��_�>��>?��"�XF��Y����I4�B��?��@O��?��=<�����=�<?�@�>�P��#ƾ�����`����p=���>�����Qv�u���',���8?̙�?R��>n���Ӡ���<H��G��?k3~?/댾�])��Q#�S�Y���7�� ��T�=ب���*�$���=�/�þ�D�W«�^D���^�>��@����ӹ�>M��)��T�ۿ�yj�H?�: ��\�?7�>�Ѡ�EK���� ���3n��'�f���о���>^@>�䆽�㚾ڍ~�dD<�j�L����>�gn��8�>Ao������zp����>��>�lm>>�齝¾Bl�?�8�1̿��?��J�]?�x�?EI�?XN?7�<����R��Ȍ	<��I?)�s?&nV?�$��l�Yl��%�j?�_��sU`��4�nHE��U>�"3?C�>G�-���|=�>~��>�f>�#/�s�Ŀ�ٶ�3���[��?���?�o���>m��?hs+?�i�8��n[����*�C�+��<A?�2>���H�!�80=�=Ғ���
?[~0?'{�h.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>��?�H�=�]�>^��=8���DZL�ӟ >���=��C��a?9~M?R]�>�=�=�8�&/���F��*R��\�،C��J�>ǂb?!�L?7�b>���� 6�7� �F�ҽ`C2�S�I�?�G� ���^�2>��:>�J>�#D�J�Ҿ��?bp�$�ؿ�i���o'��54?C��>4�?���]�t�����;_?z�>�6��+���%���B�b��?�G�?C�?��׾�R̼�>��>�I�>m�ԽV���`�����7>�B?1��D��Z�o���>���?�@�ծ?}i�	?](��L��)M~��x�w�6���=��7?:�|�z>���>���=�lv�J�����s�S��>�:�?5z�?���>��l?zo�J�B�F�1=��>(�k?@�?/�b����B>��?k������ME��f?(�
@er@,�^?���ڿ�����Ծ����,�=��i=��>�sC��J=�J�=;�i=.�<���=��>��=�¬>��>?�3>+�9>yn���z"�����͔��zG����}�K#��IH�c���Y����྇]��ԛ@���5��c(��%���b���)����=]�U?�X?n?��>}���>�D�4��;�G4���=�X�>��8?f�J?T�$?ۗS=+-���Zb�IB��E��>���7�>��Q>���>�
�>�R�><^<WG>��2>y>x>�p=���8�<?�;>喝>��>	ҵ>Y�u>�Û>S���g����x�p^O��/o����?���� 5�޷��)M	��=�@�=�8?�sg������ӿ[l��ż9?�L[���-�����U0>�?ӎL?f�=�=��Z�fB�>
eS�x�?��S�>�@�;��&�����0�>��?G�g>@w>�3���8�
Q��G���z>�q6?,W��zV9��%v��AI�d/ܾ��M>-��>��a��������I���h���|=��9?�Z?D>��e۰��Ot�؞��YT>�D[>*� =���=��L>��W��ý��E���/=֬�=?u^>Q?��'=��<=��>�+��D��7��>Z��>YpS>��/?��#?�I!�ۚ �!a���S!�M�h>�#�>�X�>�*>���c��=B��>׼3>m�)�t��f������i{>ɱ�����ĥ?���G<9��A4>�)�=�?:*�_�?�Z<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾQh�>�x��Z�������u���#=R��>�8H?�V����O�\>��v
?�?�^�ߩ����ȿ3|v����>V�?���?f�m��A���@����>9��?�gY?{oi>�g۾5`Z����>л@?�R?�>�9���'���?�޶?ӯ�?:�H>�~�?��s?<��>�px�;�/��9������nv=��O;�>��>�p��AF��ғ��q��~�j����<9`>V%=s�>t��kR�����=<��������`���>F�q>ITH>�ߜ>�� ?��>TS�>J=cH��0���o���1@??O�?_"^�*?���v�0l?�k�v�G��>�Z?w ,>	���$�7=U�U?^Љ?�xg?���>dQ0����Y@������d܆<BX>t�>�Q�>Oq��~>�G6��W�����><�?��>m�����н�L<=�7�>[��>��?�?(>Qe ?��#?#=k>�ұ>�uE�`���[F�3Q�>��>؁?ja~?�?:���D�3�n*�����C�[���L>�x?bV?�3�>�|��֭����^��{D��O��Y��?8Pg?�Tὁ8?�ʈ?�W??��A?�of>�'�� ؾ!O���$�>��!?%���A�o&������?��?���>a命�gֽ,QԼ���N�����?�\?�&?AH�Ү`���¾�!�<I���x�F<�vM���>A�>����D1�=�>���=�/m���6���l<�/�=8ƒ>���=��7�Ĺ��>=,?D�G�!ۃ���=z�r��wD�p�>�JL>
��]�^?Ml=���{�����x���U�� �?���?Uk�?�
���h��$=?�?Q	?�"�>�J��~޾���Pw�5~x�|w�H�>���>�l���"�������wF��)�Ž>�E��>��>�?&� ?'�O>S�>����'�x�����^��l��i8�W�.�Ŝ��Р�g�"�_��k'¾m�{��C�>�q��(�>��
?^.h>D�{>��>�xȻ�C�>=R>�>N]�>�X>�5>��>y <��н��Q?M����N'���������A?G�c?� �>�ao��م���� ?P��?Hn�?W�r>�g�:�)��?g��>;�zR	?�2=����2�<찾Q��鉽6�!�BE�>Rsν}09��jO�=e���	??����s˾�Sʽ�랾@��=/�?4?��(�+g{��3��!6O��O`���=t2���3��SQ�p���(��@5��ұ��4S8��=<q�(?�B�?m���H!����ON���E��!�>��>���>g�=T��<����� ��tK�X<O�A����MT>n�E?�N�>�DH?G?�q,?�kU?x�>�b�>tV߾gW�>}ǽ+��>�1+?ΟA?�>?��?3Z�>B�?$d`>D}Ľ��߾����>�?�}*?�w,?���>�O�� ����>�60>ocs����|Ed<i[=PC�����"�=�L�>�i?�d�ː8��K����j>Ru7?���>.g�>۳�����O��<���>�h
?�>Q����Fr��+���>���?�W�nK=�*>�T�=���؏���c�=�Y���ݏ= ���j�=�g <z�=�t�= .L��@�6&?3;�i;�F�<Du�>��?吊>�G�>[9���� ���݁�=Y>�S>_>:Eپ�}��$��K�g��]y>�u�?�z�?��f=�&�=���=�{��U��L��c����Z�<(�?�G#?LWT?���?'�=?pj#?��>�(��L���\�����z�?( ,?� �>����ʾ�¨�L�3�
E?b�?��`��a���(�¾Q^ҽ��>��.��}�C����D��ϫ���a�����?��?:�.�6�A��젘�Ѥ����B?��>e�>���>h�)���g����;>��>F�Q?֦>֡P?�6�?��J?��,>�%C�y͝��͒����5�߼��+?g�?WI�?��h?��>NL<�ʽ�ɾ��m6N��	ݽ���d��u�@>�3�>�t ?���>#�>>�?�u�H;�E�;,�=�q`>/�>s9�>W�?��>{��=EH?-�>5󾾤���դ��˂��f1�bv?Pq�?�+?�=jF��F�B�����>�&�?�«?Q�*?��Q����=,�Ӽ�⵾�pq���>竹>lϙ>^��=֟A=io>[��>B5�>�	�l��5�7��kJ�xA?��E?���=�Oȿ��h�r萾m���2<;]$��8S�X�Ľ�Dx���ͼ4���
�ʙ��Υ}��~��!쬾����~՛�]�n�B��>9�=>�C>�%)>Ѭ=���A�Լ�.=����Yw";���W4=��ؼ��<e���c=�tS:��"<��?��˾��}?}>I?r�+?w�C?/�y>d/>��3����>�{��1B?e'V>�GP�Z����;�j����!��۳ؾlw׾*�c��͟�~O>&"I���>�,3>�D�=���<�%�=�s=l؎=;�Q�g-=.�=2E�=o[�=(�=}�>uT>�6w?X�������4Q��Z罥�:?�8�>�{�=��ƾo@?��>>�2������yb��-?���?�T�?@�?:ti��d�>I��x㎽�q�=b����=2>���=r�2�O��>��J>���K��R����4�?��@��??�ዿϢϿ9a/>Z�7>�">=�R�L�1�}�\��b��NZ�v�!?�9;��W̾�0�>�=J߾~ƾ�q.=�j6>�b=�P��K\�y��=��z��;=�k=�Չ>�D>�պ=l/���Ķ=�yI=:��=Y�O>.���37�l�+�	N4=��=g�b>�2&>���>i&?�0?�c?D6�>�Up��`Ͼ���睌>��=Ef�>��=��G>���>[�7?�`C?1�K?��>fA�=�պ><��>�p-��m�f�例4����<�A�?�?nж>�q<��;�����[=��ý$?��1?�"	?��>�����t\=��,��l���<4�=d�v�臽|��<NA��"��b�=k��>ף�>��>���>U�E>cm�>���>��>��X=\�<=q1�qpy=��y�;��=N�=\�)=��O���9=��<1R���ݎ;�麛ڰ;�=*㺼��=!��>}<>ج�>N��=����C/>帖��L����=�G��a,B��4d��I~�I/�}V6�s�B> ;X>�}��?4����?{�Y>m?>���?TAu? �>� ���վ�Q���Ce�/VS�o˸=-�>��<��z;��Z`�z�M�[|Ҿ���>��>�>��l>�,��$?�_�w=��c5�G�>~������]&��;q�k@�����ii��Bں~�D?�D����=�~?K�I?��?��>��I|ؾ�60>/E��΄=_�!q�:T��H�?H'?��>�h�D��̾�0��H��>��H���O�*���݊0���R����~�>�����о�%3��b������sB�Gr��2�>�O?(�?�Wb�H��cKO���[���?��g?%��>�J?$?����<L�g��c�=5�n?o��?*�?>
>�	>.�?�s�>�)?�ޡ??�?PW?q�9�p?������>�f��_����=
 �[�>���>�-?Y9?+�<T�!)Ⱦh׳�h�۾��T=?k>��>~�M>�܈>+>��8��
�=@S�<r�a>��H>�$>e}�>��=�޾8�ߠ?ş>2�>}�?&^�>�=>@���L���UVL�u��!�[v=;��=��)�q�>��n=1�>ӪÿT�?	FB>���X�?�����ü���>U=�>����>,"h>>M8<���>�n�>az�>��>�gz>�FӾ~>����d!��,C�a�R���Ѿg}z>�����	&���Sw��"BI��n��|g��j�M.��V<=�!˽<*H�?R��� �k�#�)����\�?�[�>�6?�ڌ�d��į>���>�Ǎ>�J��d���Xȍ�	hᾛ�?>��?�;c>��>M�W?)�?��1��3��uZ���u�c(A�/e�A�`�~፿�����
�|��-�_?�x?9yA?�U�<:z>K��?��%�=ӏ��)�>�/�(';��=<=b+�>*���`�f�Ӿb�þ�7��HF>��o?5%�?uY?TV�A�Z�>��*?	d4?Y�m?�E?�3?
����c??��>xX3?�I!?G( ?]�4?�i ?Y�9>�s�=$�*=']�=y�Ƚk��·��c<VS���n��ě =�]=��=�X�:3�=��nxO��(=�?<�I�;���=�?�<[>�=<��>��]?�@�>��>��7?q���i8�{Ʈ��(/?��8=����(芾1�������>I�j?���?�^Z?�`d>��A��C���>�N�>%�&>�H\>l�>#k��E��߇=�Y>f\>sV�=�(M�~ׁ�R�	�ᔑ��c�<�^>��>1ϴ>����b�=�䖾Hp����	>ݰ��쟄�C�2���-���V�޽�b�>_�N?HH?(Z0������.��Y��v
?�xp?Cz?�<�?sJ�<�3�/�A�y�P���v��>�En=9@��򔡿|���nZ���;?c>>fDq�$v�6�>�[�� �$~��T��9��-�>�$���=u>4��Q�^��/a����-��"���Z�����Ƭ��d9?T��=_���-�ƶ��v%�>��>��>�ؼ����`l�����<W>�?�>y]�<j���R_6�e����.�>�HE?��a?K�?�w����r�d�B�I� �x2������M�?���>�?� G>��=����}����d�l�H����>h-�>�s���H��f������"����>9�?�>��?�N?J?9�_?��)?��?��>���A����9(?�U�?p�>l�	���� 2#��5+�S��>[T?g�&�d��>ud??�d2?�@?J��>�(>g%ھ�6��-�>d��>�y�Lӷ��o�>�+V?���>G�X?��^?
6>s��\Y���v={�
=8��=u�0?�j9?��&?�?��?&�0�¡>i0�>Lr\?!IG?�_d?�ig>=�S?Y(+��q�>P�>�߻=�{�>�,?��E?ʵa?
�<?�F?�*:=؎,�t�<�22���3<�J���z=���=�9A� �]�s�ӽ�0>��=[R�=η>��<��P0+=rG�	�>u>���e`2>%���;��g4C>���������G4��=�>�K?�ْ>�j!�qَ=���>g��>����&?aM?�u?��^�%c��ھ��E� Z�>$B?�'�=�am�������v�8�O=EJl?�^?k�X�������c?g�g?�۾�Cr��;����e���Dr?�#�>��߽wS =�\@?��e?�¡>�p��9����g��ߟ{�lM��K��=�?�>�q�p�X�anS>�;?? ��>�8>Ze>��侼�x�+쥾�?�|�?���?��?�48>��S��տ��������[?�3�>����mt!?�|����ʾ�����1���ݾ�����N��_���Wס�?W�[E��㽑��=�U?�t?��u?��^?� �Td�yvb�=*��x�Z����k)���B�$}?��rD���s��5�#����p��7F�<�T}���F��İ?�'?��4�d3�>F`�� -得Ѿ�k>[���,���=����3z=܈�=��\��T3��>��ݫ ?�M�>3��>f;?Q�X�o�=�]�5�Ϋ7�և�>�.>%ˡ>��>'��>:d��8R�I��v�Ҿ�t�������>d1a?]�W?2�r?�7�<�9� I��(Q>�?�����b��NK>�0�>7�>h���M(�<'��l;�gu�°"�ꌾR�	���b>F�O?Zդ>=�>��?���>���������'���$����7<�>.eX?��>өf>���� F����>��l?l��>N�>v���mZ!�?�{��ʽ&�>gޭ>���>��o>L�,�h#\��j�������9��q�=	�h?[�����`���>�R?o�:�G<(|�>��v�~�!������'���>({?J��=�;>�ž5$��{��8���)?��?����#'���>(#?���>~`�>f��?BX�>a�����<�m?NI^?�I?�"@?��>w�4=�q��eĽ�F&��=Hׇ>[�n>c�=���=>���Ge�L6���^=���=�i1�Т��$�:,E���ɐ�K��<�>>riۿ�FK�M�پ�����;
�]ވ�����i��t���]�����x:x������&�3V��+c�b�����l����?;�?j��3)������p���P���I��>޵q�~������Y��|�ྷЬ�Th!�g�O�.*i�2�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾w1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@��A?8�!���� �=��>�m?��=>E�3�q��K󧾊e�>�J�?`�?$��=�T�E��3�b?��;��B�����=��=w�)=k
���a>���>P�-�+X��þ��k.>ԇ>?5� ����a��!=�WT>�P�O�Y�5Մ?,{\��f���/��T��U>��T?�*�>Q:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?aD6?���>�d&��t�݅�=y6�p���z���&V�}��=]��>b�>Ă,������O��I��O��=&�=���W^��z۾'�='�V��&=[B�����>�e}���� �a̜=�Ӳ>܊�>���>���>��>TH9?O?���>O	1>`��:�ֽ��a�н����1M����_���C�H���������۾�E"��k:�%�����9�2��=�ZP�ǩ��(!"�KQd�j�I���/?��>�ɾC�N�k+�:�˾`�����Nǽ��Ӿ�&4�So����?�@?F腿ՁY�	L�5��Mb��b/Y?�z��3�������=�^����-=�@�>1��=�D߾i�2��'R��N0?��?%���b/���0/>����;%=�/+?2�?Og<v�>�&?��(��dݽ�P[>�4>�> (�>,�	>�֭�˰ܽ�h?۱S?�.���p��ޓ�>S���Rx���n=��>��3���ݼnY>3g<�����=��8̖�	�<pV?f�>�=!�6W"����� �:٧1=l�l?���>���>�Pr?�pH?].�=L�Ҿ�mF�5��aŸ=�gN?'#]?��> ���Ծ&����-S?y o?6vL>F���#�R��i��C?�s?�?�;5�&]a�1��e���l??��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?x�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������-��=}����?N��?����ɽu��s-\�`b=��O�=��=�1N��i>:����K����l����ӾH��iF�>z@��*>�9�>�y���(�R�1����������&�>�f�>~	]�@���󟿄���}�~�֘`�##
����>��>���Pv����{�Ol;�䧭�6[�>�k
���>vuT�ɇ��������<�>�u�>A��>�c���o��㣙?�����"ο�ƞ���Y?m[�?�}�?�U?��<<��w���{��i
�FG?
qs?\�Y?0� ��v\�:�3�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�a�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�[�_?+�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?M^�?h�?ѵ�� #�g6%?�>f����8Ǿ��<���>�(�>*N>OH_���u>����:�i	>���?�~�?Pj?���������U>
�}?���>c�?�>wB�>0��=����C.߼/C�=o��=�@_��?TbS?�C�>g]�=�<�UA/���D��S��z�KA�ky>P�k?�#X?�>a��*`��"�����W�%�Dپ�oa"��#�WнO�*>y�B>��>��&��QѾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ta~����7�i��=��7?�0��z>���>��=�nv�ݻ��U�s����>�B�?�{�?��>!�l?��o�O�B���1=4M�>̜k?�s?2Qo���h�B>��?"������L��f?�
@~u@_�^?*lѿϘ�G�𾟰ԾP�>rN=�_>�'&>��8�^w������-�u��=�?�>���>~�~>���>>}�>��q>غ����!��{���1k>����{����d�T�)���u�����=���Y����=(F�=�������C�q�<l1�=�WU?kU?�=p?E��>�ҳ�9	>T�� ��<�� ��#�=�ߘ>�8?:�M?#�$?aa]=Kޠ�3�e���������k�����>�?~>4��>)��>��>�B�d0>~=><܉>w(>�p=���::� =��S>�٥>���>��>��E>U�(>�������Pk��Op����\��?є��BI���������W|��?�~=�%)?J��=�8����п$���d$E?,��	����'�z?�=J�-?�)W?_�>����y�m�tR>N�:�c��j>�bݽ�^�8�%�5�N>��?N��>^n�>*�)���Y��e��W��s >9?u?���Fv�ۉ�cZ�<���c�>�>�Ľɧ3����h����){��$=s�*?��?	ͽ��澮8�?����>�?>�,A>V� >PR>>��=�L�^<��(��='s�= �>M3?�->��=(�>�ɖ��O����>�0D>�1>�R>?�9%?e��@{��FĂ���0�>w>�l�>c��>'�>�+H�[g�=�`�>ja>���뉃��Q���<�VY>Yh��`��P����j=����}_�=T��=a����,:�+-=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾWh�>Rx��Z�������u�>�#=/��>�8H?�V��n�O��>��v
?�?�^�ᩤ���ȿ;|v����>M�?���?a�m��A���@����>=��?�gY?�oi>�g۾(`Z����>ʻ@?�R?%�>�9�o�'���?�޶?ү�?e2e>��?>�t?v�>�1R�cgX�0ݿ�<���d�ɼ�(N=�m>>=I�Ǿ�6n��ˢ��ʔ��R��W.����=oܨ=�*�>Q[��H� ��=�y�4����5�=Y��>3�L>���=�Y�>tV�>iӓ>�x�>�ϫ=��ڽ2|�������K?S��?���i�t�I"�飀=_�x�p��>�y.?�ż�M�H�>|�Z?SMz?�hS?́>28��0�������)���}�;�<W>��?��>y���S>�N�%�^�>f��>�f=�"ξP�E�%+<���>�_$?@��><k�=�� ?��#?��j>b��>WxE�FL�� 'F�B��>�F�>V??)�~?3�?l߹�r�3�A���񡿒�[�m?M>�x?�R?�ߕ>w���.���)�?���F��ݒ�]��?�Sg?8~�I�?��?qb??�{A?Guf>�I�0�׾�b�����>Q�!?	�E�A�TN&�P�J}?�N?T��>�,���ֽ��ּe��_w��c�?W%\?==&?3���(a���¾�F�<��"���W��o�;��D�ȼ>��>_���U��=F�>{Ѱ=�Pm�/?6��tg<�{�=Z��>��=(7�����#=,?K�G��ۃ���=��r�1xD���>�IL>����^?Zl=��{�����x���U�� �?���?Qk�?��)�h��$=?�?O	?["�>�J���}޾2��Qw��}x�}w�S�>��>�l���E���י���F����Ž�*����>x��>E ?u ?$gO>�h�>i��|�&����~��h�^�T��aX8���.�|}�����^�"�3?�w����.|��>F���ز>Ś
?�)h>V�{>O�>a����'�>�vQ>�>��>��W>U�4>��>{<�VϽLR?]���߻'�T��\���75B?�nd?&+�>ai���������?$��?�q�?K>v>cuh��$+��k?>�>����l
?Y:=^�㹊<ZG��1���F��+��>��>TV׽�:��
M��hf�ye
?92?�Ս���̾t׽�Ǆ����=?@�?�i&?�6=��p��#����^��'b��fa���U�r����l߄�B䟿�Z��mꌿ�z7�`��!&%?z��?{Y��]&��iо2�s��V��[�>�{?�'�>���>)�>>���^�>���X���$�q�����>6hZ?��>>�K?{�$?6)?��W?k!?��>��U0`>X�(>�Y?s�?��R?�A??�?�?�A!?�->�c<���n��n?v�?��??�f	?a�?Y̧��5�^�ӽ��'���J�dn<��
Z=%��h�;���:�>�T�>�a?X�ђ8��{��M�k>��7?ު�>Ƿ�>N����C��-��<��>ʸ
?u�>����yFr�P��T�>��?����H=h�)>q.�=��}���ź4��=~&¼X
�=��]�9��{<�.�=k��=�b���k6�Lּ:�5|;��<�t�>��?d��>�D�>�>���� �;��'i�=�Y>�S>\>nEپ~��h$����g�#^y>�w�?rz�?x�f=�=��=0}���T�����;������<��?�I#?aXT??��=?�i#?F�>�)��L���]�������?S�+?���>��������w���?�CB�>�в>�F=�t���:�.�&����J	;;�F>�^���{���ҡ\�ۋ_��/��O�v��?���?{p�=
�J�a��ͤ��Z���Q?�>$?��?D�?�qƾ�>M�����1z�>�P?�vO?>S�>�)M?^�?�]{?�W�=��6��V���㣿�7H��i>�58?y�z?�$�?��y?���>Gԭ=�y�O%��T�&�]����@ȽK
[����;��(>�r�>���>�Z�>3�$>)��ҿK<8�������g>��>D:�>y��>e��>�V�={�G?C��>E-�����Z뤾����I<�I�u?ϓ�?�u+?�v=C_�R�E�0��g#�>YZ�?7�?c%*?1�S����=�ּ���r�E�>��>�-�>ļ�=�E=��>{��>N��>G��EY��^8���K�E?�F?|��=������t�R����xi���o<������4�ֹҽ9oG�! ݻ[G���]�XrҾ�BI�>p��GT�BE��̞[��2���?\R'=g��=���="��<vp���� =qm�=�� <t�H=S�V���Ӽ��<��������;�ud�<�7;^�<��˾Ѝ}?�;I?��+? �C?��y>%C>=x3�J��>w����@?V>μP�����ʎ;�����c���ؾs׾H�c��ʟ��C>SI�˶>W53>�G�=ok�<D*�=�>s=;��=JU���=L�=@O�=�h�=���=��>/Y>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>q�0>�G�=�]S��B/�~�]�J�b��V�?�:��z;��>&k�=����ľ*�C=��;>�~u=����rZ�v�=�"��a�5=#�l=+4�>-�E>�,�=�ק�E��=��F=�U�=*�I>��y:e@��B/�Ӫ=J��=rPX>=�)>�k�>{�?�A?�\?�Ƕ>*�|��F���򫾬��>J0=}Y�>��=N�>!��>��?$q-?��,?��>���<	y�>�ږ>_V3��l�K��F��H��=n�?N?m��>���<d{��_�%�y�B���;�?0F?��?��>�& �4v̿A�E��B���=���<�s=�&F��|ͼF�9�p#��^ U��׽�O>< �>�F�>�j�>7��>�W�>?)�>�V>�k�=�	>�$!�R�ǽW��:|b<��>P�=�բ��,= �ܼ�g���=
�=���=q>)������=��>e<>۬�>>��=���D/>㸖��L����=�G��f,B��4d��I~�H/�mV6���B>0;X>�}��=4����?T�Y>�l?>���?WAu?3�>� ���վ�Q���Ce�<VS�\˸=5�>��<��z;��Z`��M�Y|ҾJ��>~�>��>̿l>�,��,?��w=�=�H[5��,�>�m���6�����q��8��F�5i�g���B~D?A��}8�=8~?�I?��?y��>�옽M�ؾ��/>�2���'=Q��!q�.��m�?�'?���>��B�D�F̾����>Q=I�^�O�!��0��l� ɷ� ��>����$�о�$3�ig������B��Jr�X�>�O?��?;b�iW��DTO�)���!��|q?R|g?N�>uK?�>?�1��{� s���w�=��n?̳�?�<�?�>O�>lm7�e��>!:?��?5+�?Lp?O�ֽn?���-�D>�s\���<��s�=�-`�l�>Q�?`l�>�
?ifG����	R뾷V;̚���%=�I�=�S�>�>%q�>�{=�2�p���]%>+�>���>��>k�>%w�>�﮾�� �q��>�s$>Fwf>&T#?`1�>]��=�Ζ�I�h=�e�K���ϴA�L,���
��)�=��i=���=�3u=C��>fĿka�?�)5>3��l�?}�����=k��=ۚ�>Z��gC�>���>xY�=��>VI�>��=s��=��V>�BӾ:�>����e!��-C�'�R���Ѿ2�z>-���k&�������~EI�|t��Mi�(j�/���==��~�<�G�?t���<�k���)�����Ȗ?�\�>16?�ٌ�K���>���>vȍ>F��ώ��tǍ�{d�{�?���?>;c>x�>	�W?�?��1�M3��uZ���u�(A�e��`�u፿����
����&�_?�x?yA?�T�<f:z>'��?��%�!ӏ�)�>�/��&;�u@<=A+�>�)����`�ϯӾ��þ8��HF>E�o?6%�?DY?zSV��[v=�A>t/?��.?$;�?��<?e�=?��߳0?	>Yx?�P0?.�)?e�.?L?
�j>;�=+��=-�>�����ds��Q��5 ���1=��!T�<NSO=�:�=���<�,<���F.��s��9EF��ɓ;�#h=��=�� >~ۦ>:|]?_�>�Æ>h�7?�p��8��X��P^/?�8=�H������������5>E�j?	�?j>Z?R�d>D�A��AC��>t=�>�%>g\>=O�>���YE��u�=�>q >��=,pL��r��7�	����<w�>Y��>� |>���6�'>2}��u-z���d>��Q��κ��S���G�b�1��rv��U�>}�K?��?Z��=�_龲$���Ef��/)?Da<?gNM?=�?: �=��۾��9��J� >���>{s�<���K����$����:���:�s>j9��oSp��x�>U}վ���{���A�K&�w�!>0�7����>��M��3!��.�\����V�'�|�D��ͦ� (���@?���=A˾i�ʾ!���I�>R�>�9?��<=���D`�J�~5~>H?� �>к:=Y���D��48�+�>b�E?�:d?z��?�ہ��1s��HB����ࠜ�pv��?�K�>��?,&I>���=T���%���P`�nWI�9f�>��>W���H�	៾���Z0�Ϧ�>��?�>��?�EV?!f?>?\?�'?�?��>X�`�����%L ?�-�?f,�=)�ý�HV���8�.E@�y��>.k)?/Qv��ĝ>�$"?I�,?�.&?]K?��?�3>8� B��̓>�>[Sb�3>����l>�J?�9�>�P?Z}?�>-�%�J*w�����>.H>�,?u4?��?=.�>��?)L��>ϖ?n/?��s?���?���>���>a��&޶>��=���#�>F��>al?���?��_?*�7?v鲼{��=�j�;2Xy�KC!>/�*�ڠZ�ߴ����g=�J�����r%g;[Щ��>`=�E�='��=z�ɽ�c����=%R�>��s>������0>�oľ^����A>�駼�W��Ғ��l�9�ȧ�=�y�>�?���>A@#����=�>�<�>�����'?�?�?G�;�nb���ھ8�K���>�0B?!e�=��l�����1�u��vh=��m?h^?F5W�I���
qb?�^?g��^�=��Hž�"c�����O?	?�/C��>-j}?l�q?ږ�> �g���n����"�b�m�l�=���>�n��6e��۝>�C8?�U�>�af>b��=��۾#x������?v$�?�?�׊?A<+>�n�I�	��������.]?�=�>������?G[�-ξ���������M�崧�����d���Ã���F��w�<�۽&��=Ɏ?��v?<�n?��_?0��xh�t�c��>y�q�]�E��?��%C���<��
D��$v��W����E��«�<�H��}�B�
�?x'?j?0��h�>Ӏ������ξqYE>�|������c�=k��T=�`=�oc�lD.��8���6 ?���>���>��<?*$Y��6?��,3��'6�[���L�,>Nǣ>���>/��>Ds���8�&���0̾0ʇ���߽:l>N�d?�dW?f�i?啽���8�����0+�2߽y޵���5>��>C �>/�*�?�%�'��	E��m�jX�|E��r"
�Lr1>��@?�Ճ>i�>�W�?Q?#������qu��u%�G��=W��>5N?�Բ>3�>��,���>��l?���>W�>����[!�f�{��ʽ�#�>�߭>���>&�o>��,�o#\��j��h���`9�Po�=�h?������`�W�>�R?3��:��G<|�>�v��!������'��>�|?���=��;>m�ž$$�1�{�^8��xW)??�?О��KH*��[}>g"?���>`��>��?o�>n�¾ď�c?��^?�J?0#A?�w�>�P!=]�����ǽ}D&��.=+��>�R[>��o=���=���\������C=�!�=�VӼ������<����<�T<��<=y5>LWۿ��K��%پM��$s��
��L���\������@��,��[U��3�y�\/��^�8�U�9�_�����p4i�)��?_��?�z��Fꉾa���,5��v���"�>�y������ޫ��P��[��-G��԰�Y�!�ƦP���i�:f�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >^C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾u1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�>@?��$����W=��>��?ܦA>"�4��H��%��߮�>���?9��?Pjy=��V�7��c?X3L<̒D������=��=i�=Z3���^>��>���LqJ��.̽n}7>�}�>D�s��"��[]����<�"R>k�Խ�q�5Մ?-{\�yf���/��T��"U>��T?+�>Y:�=��,?Q7H�[}Ͽ�\��*a?�0�?��?)�(?"ۿ��ؚ>��ܾ��M?dD6?���>�d&��t�Å�=87�%�������&V�a��=V��>a�>Ă,�Ӌ�t�O�J�����=����@����=b�;=���*輹{ͼ��9���M���=%p��gnE�I3���۽I�l>43>�p�>��Y>���>�PW?uWU?�³>F��=Fǽ�]���ݾ.[�=!ȾW�d��T���T���9���x��G�
��Z�z_,��ʾH�<��=��Q�B���"X!���b��G�'�.?�� >�Ⱦu�N����;pɾ��4Y���q���{;nS2��Hn�{��?S�A?�兿n3W�c���4���SX?���8��������=DV��L�"=?�>+G�=|���3��S�hl0?l[?�}���R��^^*>� ��?=��+?;�?�FX<ZB�>a_%?��*�Pp��T[>�3>�ɣ>H��>M0	>�����۽��?V�T?�������Ӑ>ya��d�z��Sb=!r>�45�����q[>V'�<�ތ���W�������<W?Y��>��)�U���E���S��>=́x?R�?���>�nk?C?���<�����S���sax=�W?�i?L�>\j���%о}����5?��e?rhO>�5h���龺�.�;7��?��n?�\?�S��D}��������6?�v?�y^�Oi������V�WF�>ӆ�>� �>��9��_�>��>?��"�XF��Y����I4�B��?��@O��?��=<�����=�<?�@�>�P��#ƾ�����`����p=���>�����Qv�u���',���8?̙�?R��>n���Ӡ���<H��G��?k3~?/댾�])��Q#�S�Y���7�� ��T�=ب���*�$���=�/�þ�D�W«�^D���^�>��@����ӹ�>M��)��T�ۿ�yj�H?�: ��\�?7�>�Ѡ�EK���� ���3n��'�f���о���>^@>�䆽�㚾ڍ~�dD<�j�L����>�gn��8�>Ao������zp����>��>�lm>>�齝¾Bl�?�8�1̿��?��J�]?�x�?EI�?XN?7�<����R��Ȍ	<��I?)�s?&nV?�$��l�Yl��%�j?�_��sU`��4�nHE��U>�"3?C�>G�-���|=�>~��>�f>�#/�s�Ŀ�ٶ�3���[��?���?�o���>m��?hs+?�i�8��n[����*�C�+��<A?�2>���H�!�80=�=Ғ���
?[~0?'{�h.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>��?�H�=�]�>^��=8���DZL�ӟ >���=��C��a?9~M?R]�>�=�=�8�&/���F��*R��\�،C��J�>ǂb?!�L?7�b>���� 6�7� �F�ҽ`C2�S�I�?�G� ���^�2>��:>�J>�#D�J�Ҿ��?bp�$�ؿ�i���o'��54?C��>4�?���]�t�����;_?z�>�6��+���%���B�b��?�G�?C�?��׾�R̼�>��>�I�>m�ԽV���`�����7>�B?1��D��Z�o���>���?�@�ծ?}i�	?](��L��)M~��x�w�6���=��7?:�|�z>���>���=�lv�J�����s�S��>�:�?5z�?���>��l?zo�J�B�F�1=��>(�k?@�?/�b����B>��?k������ME��f?(�
@er@,�^?���ڿ�����Ծ����,�=��i=��>�sC��J=�J�=;�i=.�<���=��>��=�¬>��>?�3>+�9>yn���z"�����͔��zG����}�K#��IH�c���Y����྇]��ԛ@���5��c(��%���b���)����=]�U?�X?n?��>}���>�D�4��;�G4���=�X�>��8?f�J?T�$?ۗS=+-���Zb�IB��E��>���7�>��Q>���>�
�>�R�><^<WG>��2>y>x>�p=���8�<?�;>喝>��>	ҵ>Y�u>�Û>S���g����x�p^O��/o����?���� 5�޷��)M	��=�@�=�8?�sg������ӿ[l��ż9?�L[���-�����U0>�?ӎL?f�=�=��Z�fB�>
eS�x�?��S�>�@�;��&�����0�>��?G�g>@w>�3���8�
Q��G���z>�q6?,W��zV9��%v��AI�d/ܾ��M>-��>��a��������I���h���|=��9?�Z?D>��e۰��Ot�؞��YT>�D[>*� =���=��L>��W��ý��E���/=֬�=?u^>Q?��'=��<=��>�+��D��7��>Z��>YpS>��/?��#?�I!�ۚ �!a���S!�M�h>�#�>�X�>�*>���c��=B��>׼3>m�)�t��f������i{>ɱ�����ĥ?���G<9��A4>�)�=�?:*�_�?�Z<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾQh�>�x��Z�������u���#=R��>�8H?�V����O�\>��v
?�?�^�ߩ����ȿ3|v����>V�?���?f�m��A���@����>9��?�gY?{oi>�g۾5`Z����>л@?�R?�>�9���'���?�޶?ӯ�?:�H>�~�?��s?<��>�px�;�/��9������nv=��O;�>��>�p��AF��ғ��q��~�j����<9`>V%=s�>t��kR�����=<��������`���>F�q>ITH>�ߜ>�� ?��>TS�>J=cH��0���o���1@??O�?_"^�*?���v�0l?�k�v�G��>�Z?w ,>	���$�7=U�U?^Љ?�xg?���>dQ0����Y@������d܆<BX>t�>�Q�>Oq��~>�G6��W�����><�?��>m�����н�L<=�7�>[��>��?�?(>Qe ?��#?#=k>�ұ>�uE�`���[F�3Q�>��>؁?ja~?�?:���D�3�n*�����C�[���L>�x?bV?�3�>�|��֭����^��{D��O��Y��?8Pg?�Tὁ8?�ʈ?�W??��A?�of>�'�� ؾ!O���$�>��!?%���A�o&������?��?���>a命�gֽ,QԼ���N�����?�\?�&?AH�Ү`���¾�!�<I���x�F<�vM���>A�>����D1�=�>���=�/m���6���l<�/�=8ƒ>���=��7�Ĺ��>=,?D�G�!ۃ���=z�r��wD�p�>�JL>
��]�^?Ml=���{�����x���U�� �?���?Uk�?�
���h��$=?�?Q	?�"�>�J��~޾���Pw�5~x�|w�H�>���>�l���"�������wF��)�Ž>�E��>��>�?&� ?'�O>S�>����'�x�����^��l��i8�W�.�Ŝ��Р�g�"�_��k'¾m�{��C�>�q��(�>��
?^.h>D�{>��>�xȻ�C�>=R>�>N]�>�X>�5>��>y <��н��Q?M����N'���������A?G�c?� �>�ao��م���� ?P��?Hn�?W�r>�g�:�)��?g��>;�zR	?�2=����2�<찾Q��鉽6�!�BE�>Rsν}09��jO�=e���	??����s˾�Sʽ�랾@��=/�?4?��(�+g{��3��!6O��O`���=t2���3��SQ�p���(��@5��ұ��4S8��=<q�(?�B�?m���H!����ON���E��!�>��>���>g�=T��<����� ��tK�X<O�A����MT>n�E?�N�>�DH?G?�q,?�kU?x�>�b�>tV߾gW�>}ǽ+��>�1+?ΟA?�>?��?3Z�>B�?$d`>D}Ľ��߾����>�?�}*?�w,?���>�O�� ����>�60>ocs����|Ed<i[=PC�����"�=�L�>�i?�d�ː8��K����j>Ru7?���>.g�>۳�����O��<���>�h
?�>Q����Fr��+���>���?�W�nK=�*>�T�=���؏���c�=�Y���ݏ= ���j�=�g <z�=�t�= .L��@�6&?3;�i;�F�<Du�>��?吊>�G�>[9���� ���݁�=Y>�S>_>:Eپ�}��$��K�g��]y>�u�?�z�?��f=�&�=���=�{��U��L��c����Z�<(�?�G#?LWT?���?'�=?pj#?��>�(��L���\�����z�?( ,?� �>����ʾ�¨�L�3�
E?b�?��`��a���(�¾Q^ҽ��>��.��}�C����D��ϫ���a�����?��?:�.�6�A��젘�Ѥ����B?��>e�>���>h�)���g����;>��>F�Q?֦>֡P?�6�?��J?��,>�%C�y͝��͒����5�߼��+?g�?WI�?��h?��>NL<�ʽ�ɾ��m6N��	ݽ���d��u�@>�3�>�t ?���>#�>>�?�u�H;�E�;,�=�q`>/�>s9�>W�?��>{��=EH?-�>5󾾤���դ��˂��f1�bv?Pq�?�+?�=jF��F�B�����>�&�?�«?Q�*?��Q����=,�Ӽ�⵾�pq���>竹>lϙ>^��=֟A=io>[��>B5�>�	�l��5�7��kJ�xA?��E?���=�Oȿ��h�r萾m���2<;]$��8S�X�Ľ�Dx���ͼ4���
�ʙ��Υ}��~��!쬾����~՛�]�n�B��>9�=>�C>�%)>Ѭ=���A�Լ�.=����Yw";���W4=��ؼ��<e���c=�tS:��"<��?��˾��}?}>I?r�+?w�C?/�y>d/>��3����>�{��1B?e'V>�GP�Z����;�j����!��۳ؾlw׾*�c��͟�~O>&"I���>�,3>�D�=���<�%�=�s=l؎=;�Q�g-=.�=2E�=o[�=(�=}�>uT>�6w?X�������4Q��Z罥�:?�8�>�{�=��ƾo@?��>>�2������yb��-?���?�T�?@�?:ti��d�>I��x㎽�q�=b����=2>���=r�2�O��>��J>���K��R����4�?��@��??�ዿϢϿ9a/>Z�7>�">=�R�L�1�}�\��b��NZ�v�!?�9;��W̾�0�>�=J߾~ƾ�q.=�j6>�b=�P��K\�y��=��z��;=�k=�Չ>�D>�պ=l/���Ķ=�yI=:��=Y�O>.���37�l�+�	N4=��=g�b>�2&>���>i&?�0?�c?D6�>�Up��`Ͼ���睌>��=Ef�>��=��G>���>[�7?�`C?1�K?��>fA�=�պ><��>�p-��m�f�例4����<�A�?�?nж>�q<��;�����[=��ý$?��1?�"	?��>�����t\=��,��l���<4�=d�v�臽|��<NA��"��b�=k��>ף�>��>���>U�E>cm�>���>��>��X=\�<=q1�qpy=��y�;��=N�=\�)=��O���9=��<1R���ݎ;�麛ڰ;�=*㺼��=!��>}<>ج�>N��=����C/>帖��L����=�G��a,B��4d��I~�I/�}V6�s�B> ;X>�}��?4����?{�Y>m?>���?TAu? �>� ���վ�Q���Ce�/VS�o˸=-�>��<��z;��Z`�z�M�[|Ҿ���>��>�>��l>�,��$?�_�w=��c5�G�>~������]&��;q�k@�����ii��Bں~�D?�D����=�~?K�I?��?��>��I|ؾ�60>/E��΄=_�!q�:T��H�?H'?��>�h�D��̾�0��H��>��H���O�*���݊0���R����~�>�����о�%3��b������sB�Gr��2�>�O?(�?�Wb�H��cKO���[���?��g?%��>�J?$?����<L�g��c�=5�n?o��?*�?>
>�	>.�?�s�>�)?�ޡ??�?PW?q�9�p?������>�f��_����=
 �[�>���>�-?Y9?+�<T�!)Ⱦh׳�h�۾��T=?k>��>~�M>�܈>+>��8��
�=@S�<r�a>��H>�$>e}�>��=�޾8�ߠ?ş>2�>}�?&^�>�=>@���L���UVL�u��!�[v=;��=��)�q�>��n=1�>ӪÿT�?	FB>���X�?�����ü���>U=�>����>,"h>>M8<���>�n�>az�>��>�gz>�FӾ~>����d!��,C�a�R���Ѿg}z>�����	&���Sw��"BI��n��|g��j�M.��V<=�!˽<*H�?R��� �k�#�)����\�?�[�>�6?�ڌ�d��į>���>�Ǎ>�J��d���Xȍ�	hᾛ�?>��?�;c>��>M�W?)�?��1��3��uZ���u�c(A�/e�A�`�~፿�����
�|��-�_?�x?9yA?�U�<:z>K��?��%�=ӏ��)�>�/�(';��=<=b+�>*���`�f�Ӿb�þ�7��HF>��o?5%�?uY?TV�A�Z�>��*?	d4?Y�m?�E?�3?
����c??��>xX3?�I!?G( ?]�4?�i ?Y�9>�s�=$�*=']�=y�Ƚk��·��c<VS���n��ě =�]=��=�X�:3�=��nxO��(=�?<�I�;���=�?�<[>�=<��>��]?�@�>��>��7?q���i8�{Ʈ��(/?��8=����(芾1�������>I�j?���?�^Z?�`d>��A��C���>�N�>%�&>�H\>l�>#k��E��߇=�Y>f\>sV�=�(M�~ׁ�R�	�ᔑ��c�<�^>��>1ϴ>����b�=�䖾Hp����	>ݰ��쟄�C�2���-���V�޽�b�>_�N?HH?(Z0������.��Y��v
?�xp?Cz?�<�?sJ�<�3�/�A�y�P���v��>�En=9@��򔡿|���nZ���;?c>>fDq�$v�6�>�[�� �$~��T��9��-�>�$���=u>4��Q�^��/a����-��"���Z�����Ƭ��d9?T��=_���-�ƶ��v%�>��>��>�ؼ����`l�����<W>�?�>y]�<j���R_6�e����.�>�HE?��a?K�?�w����r�d�B�I� �x2������M�?���>�?� G>��=����}����d�l�H����>h-�>�s���H��f������"����>9�?�>��?�N?J?9�_?��)?��?��>���A����9(?�U�?p�>l�	���� 2#��5+�S��>[T?g�&�d��>ud??�d2?�@?J��>�(>g%ھ�6��-�>d��>�y�Lӷ��o�>�+V?���>G�X?��^?
6>s��\Y���v={�
=8��=u�0?�j9?��&?�?��?&�0�¡>i0�>Lr\?!IG?�_d?�ig>=�S?Y(+��q�>P�>�߻=�{�>�,?��E?ʵa?
�<?�F?�*:=؎,�t�<�22���3<�J���z=���=�9A� �]�s�ӽ�0>��=[R�=η>��<��P0+=rG�	�>u>���e`2>%���;��g4C>���������G4��=�>�K?�ْ>�j!�qَ=���>g��>����&?aM?�u?��^�%c��ھ��E� Z�>$B?�'�=�am�������v�8�O=EJl?�^?k�X�������c?g�g?�۾�Cr��;����e���Dr?�#�>��߽wS =�\@?��e?�¡>�p��9����g��ߟ{�lM��K��=�?�>�q�p�X�anS>�;?? ��>�8>Ze>��侼�x�+쥾�?�|�?���?��?�48>��S��տ��������[?�3�>����mt!?�|����ʾ�����1���ݾ�����N��_���Wס�?W�[E��㽑��=�U?�t?��u?��^?� �Td�yvb�=*��x�Z����k)���B�$}?��rD���s��5�#����p��7F�<�T}���F��İ?�'?��4�d3�>F`�� -得Ѿ�k>[���,���=����3z=܈�=��\��T3��>��ݫ ?�M�>3��>f;?Q�X�o�=�]�5�Ϋ7�և�>�.>%ˡ>��>'��>:d��8R�I��v�Ҿ�t�������>d1a?]�W?2�r?�7�<�9� I��(Q>�?�����b��NK>�0�>7�>h���M(�<'��l;�gu�°"�ꌾR�	���b>F�O?Zդ>=�>��?���>���������'���$����7<�>.eX?��>өf>���� F����>��l?l��>N�>v���mZ!�?�{��ʽ&�>gޭ>���>��o>L�,�h#\��j�������9��q�=	�h?[�����`���>�R?o�:�G<(|�>��v�~�!������'���>({?J��=�;>�ž5$��{��8���)?��?����#'���>(#?���>~`�>f��?BX�>a�����<�m?NI^?�I?�"@?��>w�4=�q��eĽ�F&��=Hׇ>[�n>c�=���=>���Ge�L6���^=���=�i1�Т��$�:,E���ɐ�K��<�>>riۿ�FK�M�پ�����;
�]ވ�����i��t���]�����x:x������&�3V��+c�b�����l����?;�?j��3)������p���P���I��>޵q�~������Y��|�ྷЬ�Th!�g�O�.*i�2�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾w1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@��A?8�!���� �=��>�m?��=>E�3�q��K󧾊e�>�J�?`�?$��=�T�E��3�b?��;��B�����=��=w�)=k
���a>���>P�-�+X��þ��k.>ԇ>?5� ����a��!=�WT>�P�O�Y�5Մ?,{\��f���/��T��U>��T?�*�>Q:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?aD6?���>�d&��t�݅�=y6�p���z���&V�}��=]��>b�>Ă,������O��I��O��=&�=���W^��z۾'�='�V��&=[B�����>�e}���� �a̜=�Ӳ>܊�>���>���>��>TH9?O?���>O	1>`��:�ֽ��a�н����1M����_���C�H���������۾�E"��k:�%�����9�2��=�ZP�ǩ��(!"�KQd�j�I���/?��>�ɾC�N�k+�:�˾`�����Nǽ��Ӿ�&4�So����?�@?F腿ՁY�	L�5��Mb��b/Y?�z��3�������=�^����-=�@�>1��=�D߾i�2��'R��N0?��?%���b/���0/>����;%=�/+?2�?Og<v�>�&?��(��dݽ�P[>�4>�> (�>,�	>�֭�˰ܽ�h?۱S?�.���p��ޓ�>S���Rx���n=��>��3���ݼnY>3g<�����=��8̖�	�<pV?f�>�=!�6W"����� �:٧1=l�l?���>���>�Pr?�pH?].�=L�Ҿ�mF�5��aŸ=�gN?'#]?��> ���Ծ&����-S?y o?6vL>F���#�R��i��C?�s?�?�;5�&]a�1��e���l??��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?x�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������-��=}����?N��?����ɽu��s-\�`b=��O�=��=�1N��i>:����K����l����ӾH��iF�>z@��*>�9�>�y���(�R�1����������&�>�f�>~	]�@���󟿄���}�~�֘`�##
����>��>���Pv����{�Ol;�䧭�6[�>�k
���>vuT�ɇ��������<�>�u�>A��>�c���o��㣙?�����"ο�ƞ���Y?m[�?�}�?�U?��<<��w���{��i
�FG?
qs?\�Y?0� ��v\�:�3�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�a�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�[�_?+�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?M^�?h�?ѵ�� #�g6%?�>f����8Ǿ��<���>�(�>*N>OH_���u>����:�i	>���?�~�?Pj?���������U>
�}?���>c�?�>wB�>0��=����C.߼/C�=o��=�@_��?TbS?�C�>g]�=�<�UA/���D��S��z�KA�ky>P�k?�#X?�>a��*`��"�����W�%�Dپ�oa"��#�WнO�*>y�B>��>��&��QѾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ta~����7�i��=��7?�0��z>���>��=�nv�ݻ��U�s����>�B�?�{�?��>!�l?��o�O�B���1=4M�>̜k?�s?2Qo���h�B>��?"������L��f?�
@~u@_�^?*lѿϘ�G�𾟰ԾP�>rN=�_>�'&>��8�^w������-�u��=�?�>���>~�~>���>>}�>��q>غ����!��{���1k>����{����d�T�)���u�����=���Y����=(F�=�������C�q�<l1�=�WU?kU?�=p?E��>�ҳ�9	>T�� ��<�� ��#�=�ߘ>�8?:�M?#�$?aa]=Kޠ�3�e���������k�����>�?~>4��>)��>��>�B�d0>~=><܉>w(>�p=���::� =��S>�٥>���>��>��E>U�(>�������Pk��Op����\��?є��BI���������W|��?�~=�%)?J��=�8����п$���d$E?,��	����'�z?�=J�-?�)W?_�>����y�m�tR>N�:�c��j>�bݽ�^�8�%�5�N>��?N��>^n�>*�)���Y��e��W��s >9?u?���Fv�ۉ�cZ�<���c�>�>�Ľɧ3����h����){��$=s�*?��?	ͽ��澮8�?����>�?>�,A>V� >PR>>��=�L�^<��(��='s�= �>M3?�->��=(�>�ɖ��O����>�0D>�1>�R>?�9%?e��@{��FĂ���0�>w>�l�>c��>'�>�+H�[g�=�`�>ja>���뉃��Q���<�VY>Yh��`��P����j=����}_�=T��=a����,:�+-=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾWh�>Rx��Z�������u�>�#=/��>�8H?�V��n�O��>��v
?�?�^�ᩤ���ȿ;|v����>M�?���?a�m��A���@����>=��?�gY?�oi>�g۾(`Z����>ʻ@?�R?%�>�9�o�'���?�޶?ү�?e2e>��?>�t?v�>�1R�cgX�0ݿ�<���d�ɼ�(N=�m>>=I�Ǿ�6n��ˢ��ʔ��R��W.����=oܨ=�*�>Q[��H� ��=�y�4����5�=Y��>3�L>���=�Y�>tV�>iӓ>�x�>�ϫ=��ڽ2|�������K?S��?���i�t�I"�飀=_�x�p��>�y.?�ż�M�H�>|�Z?SMz?�hS?́>28��0�������)���}�;�<W>��?��>y���S>�N�%�^�>f��>�f=�"ξP�E�%+<���>�_$?@��><k�=�� ?��#?��j>b��>WxE�FL�� 'F�B��>�F�>V??)�~?3�?l߹�r�3�A���񡿒�[�m?M>�x?�R?�ߕ>w���.���)�?���F��ݒ�]��?�Sg?8~�I�?��?qb??�{A?Guf>�I�0�׾�b�����>Q�!?	�E�A�TN&�P�J}?�N?T��>�,���ֽ��ּe��_w��c�?W%\?==&?3���(a���¾�F�<��"���W��o�;��D�ȼ>��>_���U��=F�>{Ѱ=�Pm�/?6��tg<�{�=Z��>��=(7�����#=,?K�G��ۃ���=��r�1xD���>�IL>����^?Zl=��{�����x���U�� �?���?Qk�?��)�h��$=?�?O	?["�>�J���}޾2��Qw��}x�}w�S�>��>�l���E���י���F����Ž�*����>x��>E ?u ?$gO>�h�>i��|�&����~��h�^�T��aX8���.�|}�����^�"�3?�w����.|��>F���ز>Ś
?�)h>V�{>O�>a����'�>�vQ>�>��>��W>U�4>��>{<�VϽLR?]���߻'�T��\���75B?�nd?&+�>ai���������?$��?�q�?K>v>cuh��$+��k?>�>����l
?Y:=^�㹊<ZG��1���F��+��>��>TV׽�:��
M��hf�ye
?92?�Ս���̾t׽�Ǆ����=?@�?�i&?�6=��p��#����^��'b��fa���U�r����l߄�B䟿�Z��mꌿ�z7�`��!&%?z��?{Y��]&��iо2�s��V��[�>�{?�'�>���>)�>>���^�>���X���$�q�����>6hZ?��>>�K?{�$?6)?��W?k!?��>��U0`>X�(>�Y?s�?��R?�A??�?�?�A!?�->�c<���n��n?v�?��??�f	?a�?Y̧��5�^�ӽ��'���J�dn<��
Z=%��h�;���:�>�T�>�a?X�ђ8��{��M�k>��7?ު�>Ƿ�>N����C��-��<��>ʸ
?u�>����yFr�P��T�>��?����H=h�)>q.�=��}���ź4��=~&¼X
�=��]�9��{<�.�=k��=�b���k6�Lּ:�5|;��<�t�>��?d��>�D�>�>���� �;��'i�=�Y>�S>\>nEپ~��h$����g�#^y>�w�?rz�?x�f=�=��=0}���T�����;������<��?�I#?aXT??��=?�i#?F�>�)��L���]�������?S�+?���>��������w���?�CB�>�в>�F=�t���:�.�&����J	;;�F>�^���{���ҡ\�ۋ_��/��O�v��?���?{p�=
�J�a��ͤ��Z���Q?�>$?��?D�?�qƾ�>M�����1z�>�P?�vO?>S�>�)M?^�?�]{?�W�=��6��V���㣿�7H��i>�58?y�z?�$�?��y?���>Gԭ=�y�O%��T�&�]����@ȽK
[����;��(>�r�>���>�Z�>3�$>)��ҿK<8�������g>��>D:�>y��>e��>�V�={�G?C��>E-�����Z뤾����I<�I�u?ϓ�?�u+?�v=C_�R�E�0��g#�>YZ�?7�?c%*?1�S����=�ּ���r�E�>��>�-�>ļ�=�E=��>{��>N��>G��EY��^8���K�E?�F?|��=������t�R����xi���o<������4�ֹҽ9oG�! ݻ[G���]�XrҾ�BI�>p��GT�BE��̞[��2���?\R'=g��=���="��<vp���� =qm�=�� <t�H=S�V���Ӽ��<��������;�ud�<�7;^�<��˾Ѝ}?�;I?��+? �C?��y>%C>=x3�J��>w����@?V>μP�����ʎ;�����c���ؾs׾H�c��ʟ��C>SI�˶>W53>�G�=ok�<D*�=�>s=;��=JU���=L�=@O�=�h�=���=��>/Y>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>q�0>�G�=�]S��B/�~�]�J�b��V�?�:��z;��>&k�=����ľ*�C=��;>�~u=����rZ�v�=�"��a�5=#�l=+4�>-�E>�,�=�ק�E��=��F=�U�=*�I>��y:e@��B/�Ӫ=J��=rPX>=�)>�k�>{�?�A?�\?�Ƕ>*�|��F���򫾬��>J0=}Y�>��=N�>!��>��?$q-?��,?��>���<	y�>�ږ>_V3��l�K��F��H��=n�?N?m��>���<d{��_�%�y�B���;�?0F?��?��>�& �4v̿A�E��B���=���<�s=�&F��|ͼF�9�p#��^ U��׽�O>< �>�F�>�j�>7��>�W�>?)�>�V>�k�=�	>�$!�R�ǽW��:|b<��>P�=�բ��,= �ܼ�g���=
�=���=q>)������=��>e<>۬�>>��=���D/>㸖��L����=�G��f,B��4d��I~�H/�mV6���B>0;X>�}��=4����?T�Y>�l?>���?WAu?3�>� ���վ�Q���Ce�<VS�\˸=5�>��<��z;��Z`��M�Y|ҾJ��>~�>��>̿l>�,��,?��w=�=�H[5��,�>�m���6�����q��8��F�5i�g���B~D?A��}8�=8~?�I?��?y��>�옽M�ؾ��/>�2���'=Q��!q�.��m�?�'?���>��B�D�F̾����>Q=I�^�O�!��0��l� ɷ� ��>����$�о�$3�ig������B��Jr�X�>�O?��?;b�iW��DTO�)���!��|q?R|g?N�>uK?�>?�1��{� s���w�=��n?̳�?�<�?�>O�>lm7�e��>!:?��?5+�?Lp?O�ֽn?���-�D>�s\���<��s�=�-`�l�>Q�?`l�>�
?ifG����	R뾷V;̚���%=�I�=�S�>�>%q�>�{=�2�p���]%>+�>���>��>k�>%w�>�﮾�� �q��>�s$>Fwf>&T#?`1�>]��=�Ζ�I�h=�e�K���ϴA�L,���
��)�=��i=���=�3u=C��>fĿka�?�)5>3��l�?}�����=k��=ۚ�>Z��gC�>���>xY�=��>VI�>��=s��=��V>�BӾ:�>����e!��-C�'�R���Ѿ2�z>-���k&�������~EI�|t��Mi�(j�/���==��~�<�G�?t���<�k���)�����Ȗ?�\�>16?�ٌ�K���>���>vȍ>F��ώ��tǍ�{d�{�?���?>;c>x�>	�W?�?��1�M3��uZ���u�(A�e��`�u፿����
����&�_?�x?yA?�T�<f:z>'��?��%�!ӏ�)�>�/��&;�u@<=A+�>�)����`�ϯӾ��þ8��HF>E�o?6%�?DY?zSV��[v=�A>t/?��.?$;�?��<?e�=?��߳0?	>Yx?�P0?.�)?e�.?L?
�j>;�=+��=-�>�����ds��Q��5 ���1=��!T�<NSO=�:�=���<�,<���F.��s��9EF��ɓ;�#h=��=�� >~ۦ>:|]?_�>�Æ>h�7?�p��8��X��P^/?�8=�H������������5>E�j?	�?j>Z?R�d>D�A��AC��>t=�>�%>g\>=O�>���YE��u�=�>q >��=,pL��r��7�	����<w�>Y��>� |>���6�'>2}��u-z���d>��Q��κ��S���G�b�1��rv��U�>}�K?��?Z��=�_龲$���Ef��/)?Da<?gNM?=�?: �=��۾��9��J� >���>{s�<���K����$����:���:�s>j9��oSp��x�>U}վ���{���A�K&�w�!>0�7����>��M��3!��.�\����V�'�|�D��ͦ� (���@?���=A˾i�ʾ!���I�>R�>�9?��<=���D`�J�~5~>H?� �>к:=Y���D��48�+�>b�E?�:d?z��?�ہ��1s��HB����ࠜ�pv��?�K�>��?,&I>���=T���%���P`�nWI�9f�>��>W���H�	៾���Z0�Ϧ�>��?�>��?�EV?!f?>?\?�'?�?��>X�`�����%L ?�-�?f,�=)�ý�HV���8�.E@�y��>.k)?/Qv��ĝ>�$"?I�,?�.&?]K?��?�3>8� B��̓>�>[Sb�3>����l>�J?�9�>�P?Z}?�>-�%�J*w�����>.H>�,?u4?��?=.�>��?)L��>ϖ?n/?��s?���?���>���>a��&޶>��=���#�>F��>al?���?��_?*�7?v鲼{��=�j�;2Xy�KC!>/�*�ڠZ�ߴ����g=�J�����r%g;[Щ��>`=�E�='��=z�ɽ�c����=%R�>��s>������0>�oľ^����A>�駼�W��Ғ��l�9�ȧ�=�y�>�?���>A@#����=�>�<�>�����'?�?�?G�;�nb���ھ8�K���>�0B?!e�=��l�����1�u��vh=��m?h^?F5W�I���
qb?�^?g��^�=��Hž�"c�����O?	?�/C��>-j}?l�q?ږ�> �g���n����"�b�m�l�=���>�n��6e��۝>�C8?�U�>�af>b��=��۾#x������?v$�?�?�׊?A<+>�n�I�	��������.]?�=�>������?G[�-ξ���������M�崧�����d���Ã���F��w�<�۽&��=Ɏ?��v?<�n?��_?0��xh�t�c��>y�q�]�E��?��%C���<��
D��$v��W����E��«�<�H��}�B�
�?x'?j?0��h�>Ӏ������ξqYE>�|������c�=k��T=�`=�oc�lD.��8���6 ?���>���>��<?*$Y��6?��,3��'6�[���L�,>Nǣ>���>/��>Ds���8�&���0̾0ʇ���߽:l>N�d?�dW?f�i?啽���8�����0+�2߽y޵���5>��>C �>/�*�?�%�'��	E��m�jX�|E��r"
�Lr1>��@?�Ճ>i�>�W�?Q?#������qu��u%�G��=W��>5N?�Բ>3�>��,���>��l?���>W�>����[!�f�{��ʽ�#�>�߭>���>&�o>��,�o#\��j��h���`9�Po�=�h?������`�W�>�R?3��:��G<|�>�v��!������'��>�|?���=��;>m�ž$$�1�{�^8��xW)??�?О��KH*��[}>g"?���>`��>��?o�>n�¾ď�c?��^?�J?0#A?�w�>�P!=]�����ǽ}D&��.=+��>�R[>��o=���=���\������C=�!�=�VӼ������<����<�T<��<=y5>LWۿ��K��%پM��$s��
��L���\������@��,��[U��3�y�\/��^�8�U�9�_�����p4i�)��?_��?�z��Fꉾa���,5��v���"�>�y������ޫ��P��[��-G��԰�Y�!�ƦP���i�:f�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >^C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾u1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�>@?��$����W=��>��?ܦA>"�4��H��%��߮�>���?9��?Pjy=��V�7��c?X3L<̒D������=��=i�=Z3���^>��>���LqJ��.̽n}7>�}�>D�s��"��[]����<�"R>k�Խ�q�5Մ?-{\�yf���/��T��"U>��T?+�>Y:�=��,?Q7H�[}Ͽ�\��*a?�0�?��?)�(?"ۿ��ؚ>��ܾ��M?dD6?���>�d&��t�Å�=87�%�������&V�a��=V��>a�>Ă,�Ӌ�t�O�J�����=����@����=b�;=���*輹{ͼ��9���M���=%p��gnE�I3���۽I�l>43>�p�>��Y>���>�PW?uWU?�³>F��=Fǽ�]���ݾ.[�=!ȾW�d��T���T���9���x��G�
��Z�z_,��ʾH�<��=��Q�B���"X!���b��G�'�.?�� >�Ⱦu�N����;pɾ��4Y���q���{;nS2��Hn�{��?S�A?�兿n3W�c���4���SX?���8��������=DV��L�"=?�>+G�=|���3��S�hl0?l[?�}���R��^^*>� ��?=��+?;�?�FX<ZB�>a_%?��*�Pp��T[>�3>�ɣ>H��>M0	>�����۽��?V�T?�������Ӑ>ya��d�z��Sb=!r>�45�����q[>V'�<�ތ���W�������<W?Y��>��)�U���E���S��>=́x?R�?���>�nk?C?���<�����S���sax=�W?�i?L�>\j���%о}����5?��e?rhO>�5h���龺�.�;7��?��n?�\?�S��D}��������6?�v?�y^�Oi������V�WF�>ӆ�>� �>��9��_�>��>?��"�XF��Y����I4�B��?��@O��?��=<�����=�<?�@�>�P��#ƾ�����`����p=���>�����Qv�u���',���8?̙�?R��>n���Ӡ���<H��G��?k3~?/댾�])��Q#�S�Y���7�� ��T�=ب���*�$���=�/�þ�D�W«�^D���^�>��@����ӹ�>M��)��T�ۿ�yj�H?�: ��\�?7�>�Ѡ�EK���� ���3n��'�f���о���>^@>�䆽�㚾ڍ~�dD<�j�L����>�gn��8�>Ao������zp����>��>�lm>>�齝¾Bl�?�8�1̿��?��J�]?�x�?EI�?XN?7�<����R��Ȍ	<��I?)�s?&nV?�$��l�Yl��%�j?�_��sU`��4�nHE��U>�"3?C�>G�-���|=�>~��>�f>�#/�s�Ŀ�ٶ�3���[��?���?�o���>m��?hs+?�i�8��n[����*�C�+��<A?�2>���H�!�80=�=Ғ���
?[~0?'{�h.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>��?�H�=�]�>^��=8���DZL�ӟ >���=��C��a?9~M?R]�>�=�=�8�&/���F��*R��\�،C��J�>ǂb?!�L?7�b>���� 6�7� �F�ҽ`C2�S�I�?�G� ���^�2>��:>�J>�#D�J�Ҿ��?bp�$�ؿ�i���o'��54?C��>4�?���]�t�����;_?z�>�6��+���%���B�b��?�G�?C�?��׾�R̼�>��>�I�>m�ԽV���`�����7>�B?1��D��Z�o���>���?�@�ծ?}i�	?](��L��)M~��x�w�6���=��7?:�|�z>���>���=�lv�J�����s�S��>�:�?5z�?���>��l?zo�J�B�F�1=��>(�k?@�?/�b����B>��?k������ME��f?(�
@er@,�^?���ڿ�����Ծ����,�=��i=��>�sC��J=�J�=;�i=.�<���=��>��=�¬>��>?�3>+�9>yn���z"�����͔��zG����}�K#��IH�c���Y����྇]��ԛ@���5��c(��%���b���)����=]�U?�X?n?��>}���>�D�4��;�G4���=�X�>��8?f�J?T�$?ۗS=+-���Zb�IB��E��>���7�>��Q>���>�
�>�R�><^<WG>��2>y>x>�p=���8�<?�;>喝>��>	ҵ>Y�u>�Û>S���g����x�p^O��/o����?���� 5�޷��)M	��=�@�=�8?�sg������ӿ[l��ż9?�L[���-�����U0>�?ӎL?f�=�=��Z�fB�>
eS�x�?��S�>�@�;��&�����0�>��?G�g>@w>�3���8�
Q��G���z>�q6?,W��zV9��%v��AI�d/ܾ��M>-��>��a��������I���h���|=��9?�Z?D>��e۰��Ot�؞��YT>�D[>*� =���=��L>��W��ý��E���/=֬�=?u^>Q?��'=��<=��>�+��D��7��>Z��>YpS>��/?��#?�I!�ۚ �!a���S!�M�h>�#�>�X�>�*>���c��=B��>׼3>m�)�t��f������i{>ɱ�����ĥ?���G<9��A4>�)�=�?:*�_�?�Z<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾQh�>�x��Z�������u���#=R��>�8H?�V����O�\>��v
?�?�^�ߩ����ȿ3|v����>V�?���?f�m��A���@����>9��?�gY?{oi>�g۾5`Z����>л@?�R?�>�9���'���?�޶?ӯ�?:�H>�~�?��s?<��>�px�;�/��9������nv=��O;�>��>�p��AF��ғ��q��~�j����<9`>V%=s�>t��kR�����=<��������`���>F�q>ITH>�ߜ>�� ?��>TS�>J=cH��0���o���1@??O�?_"^�*?���v�0l?�k�v�G��>�Z?w ,>	���$�7=U�U?^Љ?�xg?���>dQ0����Y@������d܆<BX>t�>�Q�>Oq��~>�G6��W�����><�?��>m�����н�L<=�7�>[��>��?�?(>Qe ?��#?#=k>�ұ>�uE�`���[F�3Q�>��>؁?ja~?�?:���D�3�n*�����C�[���L>�x?bV?�3�>�|��֭����^��{D��O��Y��?8Pg?�Tὁ8?�ʈ?�W??��A?�of>�'�� ؾ!O���$�>��!?%���A�o&������?��?���>a命�gֽ,QԼ���N�����?�\?�&?AH�Ү`���¾�!�<I���x�F<�vM���>A�>����D1�=�>���=�/m���6���l<�/�=8ƒ>���=��7�Ĺ��>=,?D�G�!ۃ���=z�r��wD�p�>�JL>
��]�^?Ml=���{�����x���U�� �?���?Uk�?�
���h��$=?�?Q	?�"�>�J��~޾���Pw�5~x�|w�H�>���>�l���"�������wF��)�Ž>�E��>��>�?&� ?'�O>S�>����'�x�����^��l��i8�W�.�Ŝ��Р�g�"�_��k'¾m�{��C�>�q��(�>��
?^.h>D�{>��>�xȻ�C�>=R>�>N]�>�X>�5>��>y <��н��Q?M����N'���������A?G�c?� �>�ao��م���� ?P��?Hn�?W�r>�g�:�)��?g��>;�zR	?�2=����2�<찾Q��鉽6�!�BE�>Rsν}09��jO�=e���	??����s˾�Sʽ�랾@��=/�?4?��(�+g{��3��!6O��O`���=t2���3��SQ�p���(��@5��ұ��4S8��=<q�(?�B�?m���H!����ON���E��!�>��>���>g�=T��<����� ��tK�X<O�A����MT>n�E?�N�>�DH?G?�q,?�kU?x�>�b�>tV߾gW�>}ǽ+��>�1+?ΟA?�>?��?3Z�>B�?$d`>D}Ľ��߾����>�?�}*?�w,?���>�O�� ����>�60>ocs����|Ed<i[=PC�����"�=�L�>�i?�d�ː8��K����j>Ru7?���>.g�>۳�����O��<���>�h
?�>Q����Fr��+���>���?�W�nK=�*>�T�=���؏���c�=�Y���ݏ= ���j�=�g <z�=�t�= .L��@�6&?3;�i;�F�<Du�>��?吊>�G�>[9���� ���݁�=Y>�S>_>:Eپ�}��$��K�g��]y>�u�?�z�?��f=�&�=���=�{��U��L��c����Z�<(�?�G#?LWT?���?'�=?pj#?��>�(��L���\�����z�?( ,?� �>����ʾ�¨�L�3�
E?b�?��`��a���(�¾Q^ҽ��>��.��}�C����D��ϫ���a�����?��?:�.�6�A��젘�Ѥ����B?��>e�>���>h�)���g����;>��>F�Q?֦>֡P?�6�?��J?��,>�%C�y͝��͒����5�߼��+?g�?WI�?��h?��>NL<�ʽ�ɾ��m6N��	ݽ���d��u�@>�3�>�t ?���>#�>>�?�u�H;�E�;,�=�q`>/�>s9�>W�?��>{��=EH?-�>5󾾤���դ��˂��f1�bv?Pq�?�+?�=jF��F�B�����>�&�?�«?Q�*?��Q����=,�Ӽ�⵾�pq���>竹>lϙ>^��=֟A=io>[��>B5�>�	�l��5�7��kJ�xA?��E?���=�Oȿ��h�r萾m���2<;]$��8S�X�Ľ�Dx���ͼ4���
�ʙ��Υ}��~��!쬾����~՛�]�n�B��>9�=>�C>�%)>Ѭ=���A�Լ�.=����Yw";���W4=��ؼ��<e���c=�tS:��"<��?��˾��}?}>I?r�+?w�C?/�y>d/>��3����>�{��1B?e'V>�GP�Z����;�j����!��۳ؾlw׾*�c��͟�~O>&"I���>�,3>�D�=���<�%�=�s=l؎=;�Q�g-=.�=2E�=o[�=(�=}�>uT>�6w?X�������4Q��Z罥�:?�8�>�{�=��ƾo@?��>>�2������yb��-?���?�T�?@�?:ti��d�>I��x㎽�q�=b����=2>���=r�2�O��>��J>���K��R����4�?��@��??�ዿϢϿ9a/>Z�7>�">=�R�L�1�}�\��b��NZ�v�!?�9;��W̾�0�>�=J߾~ƾ�q.=�j6>�b=�P��K\�y��=��z��;=�k=�Չ>�D>�պ=l/���Ķ=�yI=:��=Y�O>.���37�l�+�	N4=��=g�b>�2&>���>i&?�0?�c?D6�>�Up��`Ͼ���睌>��=Ef�>��=��G>���>[�7?�`C?1�K?��>fA�=�պ><��>�p-��m�f�例4����<�A�?�?nж>�q<��;�����[=��ý$?��1?�"	?��>�����t\=��,��l���<4�=d�v�臽|��<NA��"��b�=k��>ף�>��>���>U�E>cm�>���>��>��X=\�<=q1�qpy=��y�;��=N�=\�)=��O���9=��<1R���ݎ;�麛ڰ;�=*㺼��=!��>}<>ج�>N��=����C/>帖��L����=�G��a,B��4d��I~�I/�}V6�s�B> ;X>�}��?4����?{�Y>m?>���?TAu? �>� ���վ�Q���Ce�/VS�o˸=-�>��<��z;��Z`�z�M�[|Ҿ���>��>�>��l>�,��$?�_�w=��c5�G�>~������]&��;q�k@�����ii��Bں~�D?�D����=�~?K�I?��?��>��I|ؾ�60>/E��΄=_�!q�:T��H�?H'?��>�h�D��̾�0��H��>��H���O�*���݊0���R����~�>�����о�%3��b������sB�Gr��2�>�O?(�?�Wb�H��cKO���[���?��g?%��>�J?$?����<L�g��c�=5�n?o��?*�?>
>�	>.�?�s�>�)?�ޡ??�?PW?q�9�p?������>�f��_����=
 �[�>���>�-?Y9?+�<T�!)Ⱦh׳�h�۾��T=?k>��>~�M>�܈>+>��8��
�=@S�<r�a>��H>�$>e}�>��=�޾8�ߠ?ş>2�>}�?&^�>�=>@���L���UVL�u��!�[v=;��=��)�q�>��n=1�>ӪÿT�?	FB>���X�?�����ü���>U=�>����>,"h>>M8<���>�n�>az�>��>�gz>�FӾ~>����d!��,C�a�R���Ѿg}z>�����	&���Sw��"BI��n��|g��j�M.��V<=�!˽<*H�?R��� �k�#�)����\�?�[�>�6?�ڌ�d��į>���>�Ǎ>�J��d���Xȍ�	hᾛ�?>��?�;c>��>M�W?)�?��1��3��uZ���u�c(A�/e�A�`�~፿�����
�|��-�_?�x?9yA?�U�<:z>K��?��%�=ӏ��)�>�/�(';��=<=b+�>*���`�f�Ӿb�þ�7��HF>��o?5%�?uY?TV�A�Z�>��*?	d4?Y�m?�E?�3?
����c??��>xX3?�I!?G( ?]�4?�i ?Y�9>�s�=$�*=']�=y�Ƚk��·��c<VS���n��ě =�]=��=�X�:3�=��nxO��(=�?<�I�;���=�?�<[>�=<��>��]?�@�>��>��7?q���i8�{Ʈ��(/?��8=����(芾1�������>I�j?���?�^Z?�`d>��A��C���>�N�>%�&>�H\>l�>#k��E��߇=�Y>f\>sV�=�(M�~ׁ�R�	�ᔑ��c�<�^>��>1ϴ>����b�=�䖾Hp����	>ݰ��쟄�C�2���-���V�޽�b�>_�N?HH?(Z0������.��Y��v
?�xp?Cz?�<�?sJ�<�3�/�A�y�P���v��>�En=9@��򔡿|���nZ���;?c>>fDq�A���c>ce�@l޾�n�hJ�s�b(I=R��? W=N��h־|��_T�=D3	>� ���!�:���Ԫ��J?k=\M��M�U��h��\>�>�Ů>;��Eu�L@��鬾�Õ=�;�>|=;>��������jG���%�N>ߕ&?��Z?��?r�¾yg�Ә'�t�ᾫ�i���>8^�>'��>?0��=��>9���H\"�K�V��tU�A��>i��>#L��F��Ͽ�����M��X�>���>MX�>zn?�<R?�"�>�c[?�,?� ?t>#��;�\��?�π?K��=�-���ɾF�Q�#�"��
�>x�+?c���'>[?�k�>�1?��M?��?��=�.����F��;�>Y��>�PO��gƿ��V>��A?(��>Ek{?z��?���9%�3�����>�����>M�k?�^?�� ?z4?
����˾C�>�h]?t�?W�a?3��>�y�<T��R�?�~"=I�>W~3?�H-?��3?z�d?��.?G?t��;�q�nR޽,����1<���ܼ$��<3S0�(����&��7���@Tv�K��<:�=�:~<���<Z�ʻ��=��<�_�> �s>����0>�ľ*N��`�@>lv��vH��'Ԋ���:��ڷ=��>g�?r��>RX#���=���>�K�>s��d4(?��?�?�>#;��b�z�ھ#�K���>-B?@��=��l�������u�i�g=��m?;�^?Q�W��#��O�b?��]?@h��=��þz�b����g�O?=�
?3�G���>��~?f�q?U��>�e�+:n�*��Db���j�&Ѷ=\r�>LX�S�d��?�>o�7?�N�>/�b>'%�=iu۾�w��q��h?��?�?���?+*>��n�Z4�1
�L&���oO?ި�>"4þf�?1Q�?׾�q��m���]�u�w��4��'4��R���	��B��:��'W�=�'?&)�?��?^e?(�ɾtw�D�m��Q��2Oh�O꾴����;�*�6�T=�?x��d�i���վ����f�~���>�y]�?I7+?�b=���>�Ȕ�1c�6!ľ<�F>���$ �l��=�����=�Η=��t��G4��ѷ� �?���>oS�>~�;?"�Z���=���0�.n1�g���Q>�3�>�Š>~��>�,�;�)
�0��̾͘p}�ͯ���w>�Sd?��b?g6S?���2�X�e�Ʋ4� ���٧��>=9?���U>D���<a>��-3��&T�����A�/�j,��ڴ���=�:+?�i�>��>& �?&?I����]n��'�������>��?z}?W�?�-�>h�<J�C���>�/l?&��>���>�9��F� ���{�T�ŽK��>�J�>Z(�>ap>�(�hY[����������7����=��h?�\��.�b�0T�>*rR?$�;kCR<鷢>txj�P�"�ˡ���1�
>8g?��=)�:>Ȟľ٭�RI{��ڊ��r?>~?����F��Z�>��?,j�>$J�>G��?^�?ҍ
�����j-?Q?-�	?��
?N%�>��L>�6>(�|���K�����>>�>���}Į���>��Ͻ��ֽa�=��'>�@t<lK�h����jR==���MK�<��>Q�ۿ� \��������������zFn��y��Xa��x�s��;�K�9�u�B[7�����@s���p�{퉾�V�|��?�e�?n����#��Ԑ�n��=4
��v�>��Y��Qޥ�oҽõ��q���"��r�"���e���{�C�v�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾x1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@JoA?'�(��쾃HX=s�>͆	?'�?>��0�*!�������>P8�?v��?h�M=��W�f
��re?�4<��F�*���S�=��=M ==��U�J>�ϓ>�8��:B��s޽�q5>�>@�#�q�ސ^���<�]>H	սӕ�5Մ?,{\��f���/��T��U>��T? +�>R:�=��,?W7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?aD6?���>�d&��t�݅�=^6����|���&V����=[��>b�>��,������O��I��R��=)��Àο�E�DB'����̄=P�=�+"������=F�ݧʾ��&�)C�=�j�=�)�>)�>��Z>b�>��o?evB?���>rӐ>�_�� ʾ��Ⱦ��� ����޽,��:�)>)<r���:��x����־7�8���*���߾�=��#�=30R������� �R�b�^�F�4�.?�t$>��ʾ��M�)J/<vnʾ���?������1̾�1�8#n�˟?��A?*����W����@���m����W?\5�����מּ��=����@�=;�>�G�=��⾢3��wS���&?�? ^��k�B�w��>�eؽPr����(?F#??!r>��>�� ?_g���߽P��=�>���>�]�>���>�O��X;���?'`Z?�P��ٌJ��b�>A�k��m���s�2m�>j��090>�]���1��[Ҧ::w��dO?ߙ�>8#�p�<�{����ػ;��=sx?R�?���>�0F?�4'?��=��̾��J�;��� >:Jh?H�c?���=uB���-ɾK���L?�~w?J[>�z��&Ҿ�y���R���H�>W'w?��?{נ��Ar�/��F!���>?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������f��r���ȣ?}a�?������bm��q�s	���><^fS���=xL׼c����~3��������Ǿ�'��*��>�	@�K=���>��;���D�ۿ�`��nt��qF�&�!?�6�>��窎�Ϙ���*���XP��@_��3ƾW6�>�>Qʓ�������{��};��v��#��>����#�>��S��ŵ�@���t4<K�>���>z�>	��j*�����?���/+ο����s����X?�R�?�s�?$?I�5<D�v��{�����G?�Ks?��Y?�6!�H�[��#5�$�j?�_��wU`��4�tHE��U>�"3?�B�>Q�-�|�|=�>���>g>�#/�x�Ŀ�ٶ�<���Z��?��?�o���>q��?ts+?�i�8���[����*���+��<A?�2>���G�!�B0=�UҒ���
?U~0? {�e.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>hH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�$�>T�?�c�=�b�>|��=W��-�8s#>B�=��>�(�?.�M??N�>�Q�=�8�d/��VF�|CR���8�C���>w�a?�L?�Nb>~
��)�1��!�8�ͽ�p1�q�J@�l�,��߽�#5>��=>>0�D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*$"Ϳ����x]��!�Ծ�ܟ=΢�=��/>����EZ
>�;F=uk��}����=/$x>�>>�[�>�P>7�5>T�*>Ym���#�t$���>��@<L�
�����*�0��S�W:K����=;ݾKо�u���(��E_��6���)�cN�
��=n�N?�IY?"&m?���>�6��d�&>J2��
=9=`9 ���<��r>�/?<??[(?�٥=Y量^�c�����ݜ����yo�>��i>��>��>�k�>�ρ=?�`>�`_>
Q�>��G>�Y=�/��%�=V�>�0�>�J�>d��>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��w�T�4:>9����j�5`>�+ �~l���)��%Q>wl?��f>�u>a�3�!e8�q�P�v|��j|>�36?鶾�C9���u���H�cݾ�GM>ž>�D�l�o���&��ui���{=x:?�?�6���ⰾD�u��B���PR>5;\>QW=l�=�XM>�ac���ƽvH��g.=^��=F�^>\"?�->���=�S�>]0��1�K�#��>�E>�D2>d�@?��$?���䋽�=����/��s>���>gy�>+>@�J���=���>F�d>}&�},y��L	��0?�ܙO>�$���:X�*	d��;v=����IZ�={�=������=�'"=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>gx��Z�������u�y�#=S��>�8H?�V����O�p>��v
?�?�^�ީ����ȿ.|v����>V�?���?e�m��A���@����><��?�gY?coi>�g۾#`Z����>ͻ@?�R?�>�9���'���?�޶?ׯ�?���<��?8��?��H>����3� 5���ߞ���p���1<O��>wF��|7R������6��}-���@���^[�ݏ�<T�M=�z[>�l��S�F�
-��0,=I����'�;�Z�>�5H==v	�n%v>�?
�>���>Z��=�꽌;b�t�<���K?���?,���2n�O�<_��=*�^��&?�I4?Uj[��Ͼ�ը>�\?k?�[?d�>;��N>��E迿7~����<��K>,4�>�H�>�$���FK>��Ծ�4D�dp�>�ϗ>�����?ھ�,���S��FB�>�e!?���>�Ү=ڙ ?��#?��j>�(�>?aE��9��W�E����>��>�H?�~?��?�Թ��Z3�����桿��[�z;N>��x?V?nʕ>`�����jE� BI�+���^��?�tg?�S�1?:2�?�??\�A?q)f>ׇ�#ؾg�����>��!?�b���A��4&�����?�Y?���>rg���{ֽ�Ӽ��:Z���?{%\?�9&?;}�a�>�¾�$�<��"��M���;,F�ך>�t>F��qb�=��>
İ=�m�|/6���g<���=l^�>˖�=�7�{��/=,?�G�ۃ�h�=��r�9xD���>�IL>����^?{l=��{�����x��	U�� �?���?[k�?F��=�h��$=?�?S	?{"�>�J���}޾A�ྷPw��}x��w�Q�>���>#�l���I���י���F��,�Ž�%'���>��>?U��>7!>>�>�럾��!�;j�3
�YB`����5�|(���A���
�=��0��|û�L1���>/�/��!�>�;?��m>Ӓ>���>"<�|�>iat>�7�>\�>��>
�r>��>�u%=�:ڽ�KR?U���ǿ'�������3B?�od?D3�>O�h��������{?م�?�r�?^<v>�{h��&+�iq?�@�>n��qm
?V:=.��Y��<�P����sX�����'��>�Q׽:�DM�pcf��f
?�,?1����̾� ׽�5���>)&�?$��>-�X뉿�k��,��.Fm��_���5�a�J��0:�H!y��q��?$��ߟ��F�W�ay��K�?�b�?�d�dU!�VMʾ��@��8�=!{�>��>g
?�w8���;���O���R��*�ńm�"(�>U3?e��>,PD?�6?2Q?��O?��>ȡ>Jr���t�> �#=��>� �>7�7?S)?0�&?/c?��*?�f>y�Ž���<پ �?�?Dv?hX?��?!{�Z|�������<�Cb�H���E�=�
U<�Tڽ�8E�+̀=�S=>I�?�p��,:��N��:�t>�P8?U �>L�>k�������u�=���>��
?Ey�>�R��9�n����q�>�X�?n����<�'>���=§���(�^�=rnϼ���=�� ���S�x��;�W�=�+�=�o����G;>�<1%�<�t�>A�?���>mC�>�@��(� �T���f�=!Y>jS>0>�Eپ�}���$��g�g��]y>�w�?�z�?^�f=��=Ŗ�=}��qU������������<�?5J#?.XT?V��?d�=?jj#?�>+�cM���^�����ͮ?u!,?��>�����ʾ��ω3�؝?h[?�<a����;)��¾��Խܱ>�[/�g/~����2D��녻���o��1��?쿝?�A�L�6��x�޿���[����C?�!�>Y�>��>N�)�|�g�q%��1;>��>lR?���>&�O?�"{?+�[?)�Q>8�$߭�ː���b*��#>�??���?�ʎ?]ox?�a�>"> V+�[.�����=��Ev�Q����P=MPX>�j�>[��>,��>��=^�ĽH���r=�n5�=ʄc>���>E��>��>'Ax>�·<xB?� ?w��]�2�<���Ɍ��!���z?���?��%?�ʳ�3j��9����i��>&��?���?�e=?89���=D1!�t�ľ �w���>P�>��>��=�ѱ=��\>�ޱ>�͑>����-���C)C��(��t�?�J?��e>_ƿ�q���p��Ɨ�_d<����
e�Ҕ��[�u��=繘����F˩���[�����a���2�������K�{�U��>~|�=��=N�=�c�<n�ɼ0ڽ<-K=�<_�=�p��Qm<��8�+ϻ����+��ۆ\<��I=���˾�L}?�I?��+?r�C?�z>b�>.�/�0s�>4���А?]W>?O�s5��i/<�ߨ��A���44ؾ,�־n d�蟾�(>�6I��M>�3>���=Jǉ<{��= �j=�a�=/V��=P��=gܹ=���=]�=�e>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��7>�>^�R�#�1�ؔ\���b�YsZ�Q�!?�G;��M̾V9�>��='߾P�ƾδ.=�6>}b=�`��S\���=�z��;=� l=<։>T�C>�q�=h2��D�=?�I=���=��O>�ϕ���7�a,��3=C��=�b>�&>t;�>a�?w�/?v4b?w��><�z�1;������>��=�!�>�¡=!V?>��>�<9?�fE?�G?P�>X[=3�>@J�>e�+�r�r����©��K�<�s�?��?�8�>�5�;-VD��D ��6:��a޽I?�4?�/?Ł�>_V�����Z&���.��|��|%��[$+=knr��qU�=0��Ai������=9r�>���>(�>RTy>]�9>��N>"�>ۦ>%�<�u�=���q��<J�����=%�����<�
Ƽ��{�`%�H$,�PU���D�;<T�;� ]<�s�;}��=���>�;>)��>���=���B/>����#�L�+ǿ=TF���+B��3d��H~�6/��V6�p�B>�;X>Xy���3��$�?�Y>�m?>J��?JAu?~�>��{�վ�Q��Y?e�TS�ȸ=O�>�<��z;�4Z`���M��|Ҿ���>���>��>��l>�,�:$?�ыw=�#��b5�N��>}��%R��M�;@q��>������Yi�j��D?OB���V�=�~?��I?�ޏ?ŉ�>�Ҙ�mؾ�X0>�D����=����p������?�'?p��>M���D��H̾=���߷>�AI�H�O���ϰ0����`ͷ�Ǐ�>������о�$3��g������<�B�xNr�(�>�O?T�?�8b�{W��|UO����#���q?�|g?�>�J?�@?8+���z�Qs���u�=��n?~��?=�?�>���=h���!��>�	?��?/�?��r?;7�aK�>	[�;�{.>e��'O�=(9>h�=4�=s�?��
??�����	��%��ۆ^�L�=��='G�>��>��d>���=��W=n��=�_>���>�t�>r�f>֜�>*	�>���a���l,?L	>U6�>/@,?�߂>z�2=�r��;[�<6��i0=���aɽӠ���m
=�Į����<�d����>��ſ�a�?��h>����]?�/�Qޛ�k^>��k>���G�>��G>�?r>�T�>2ؽ>�>�k�>�A<>�FӾ�>����d!��,C�q�R���ѾD}z>����N	&����v���BI�yn��dg�vj�G.��B<=��ǽ<!H�?U����k�N�)����W�?�[�>�6?:ڌ���ɯ>`��>�Ǎ>�J��j���Xȍ��gᾬ�?5��?�;c>��>O�W?�?R�1��3��uZ��u�L(A��e�Q�`�p፿�����
�����_?��x?yA?�K�<,:z>?��?��%��ӏ��)�>�/�';��B<=�+�>*���`�;�Ӿ��þ�7��HF>��o?@%�?�Y?�SV�\��;@��=߫$?��2?.�x?^S0?]8?�|���^?�->�=?��?R�:?9*?(��>��)>�S%>G=Λ�=�� ���\;�k��{��ݠ�=�/>?�������ɽd0j=X�Ƽ�eM��=���:���<��=s�>u��= ק>z�[?,J�>�Ci>��6?a���u7�������8?���=4ߌ�}���t��}��ɻ�=Q�a?�Ѩ?G�Y?d��>u�A��T�k>И>"�>>�qT>%��>���D�K�/,�=Ś#>W;'>��=������ԓ����:���>���>�1|>P��x�'>q{��p/z�_�d>��Q�[ɺ�h�S�z�G�f�1���v��Y�>.�K?�?䠙="]�`&���Hf�5/)?p]<?�NM?�?��=^�۾q�9���J�U<���>@b�<8������#��f�:�`��:�s>�1��A���c>ce�@l޾�n�hJ�s�b(I=R��? W=N��h־|��_T�=D3	>� ���!�:���Ԫ��J?k=\M��M�U��h��\>�>�Ů>;��Eu�L@��鬾�Õ=�;�>|=;>��������jG���%�N>ߕ&?��Z?��?r�¾yg�Ә'�t�ᾫ�i���>8^�>'��>?0��=��>9���H\"�K�V��tU�A��>i��>#L��F��Ͽ�����M��X�>���>MX�>zn?�<R?�"�>�c[?�,?� ?t>#��;�\��?�π?K��=�-���ɾF�Q�#�"��
�>x�+?c���'>[?�k�>�1?��M?��?��=�.����F��;�>Y��>�PO��gƿ��V>��A?(��>Ek{?z��?���9%�3�����>�����>M�k?�^?�� ?z4?
����˾C�>�h]?t�?W�a?3��>�y�<T��R�?�~"=I�>W~3?�H-?��3?z�d?��.?G?t��;�q�nR޽,����1<���ܼ$��<3S0�(����&��7���@Tv�K��<:�=�:~<���<Z�ʻ��=��<�_�> �s>����0>�ľ*N��`�@>lv��vH��'Ԋ���:��ڷ=��>g�?r��>RX#���=���>�K�>s��d4(?��?�?�>#;��b�z�ھ#�K���>-B?@��=��l�������u�i�g=��m?;�^?Q�W��#��O�b?��]?@h��=��þz�b����g�O?=�
?3�G���>��~?f�q?U��>�e�+:n�*��Db���j�&Ѷ=\r�>LX�S�d��?�>o�7?�N�>/�b>'%�=iu۾�w��q��h?��?�?���?+*>��n�Z4�1
�L&���oO?ި�>"4þf�?1Q�?׾�q��m���]�u�w��4��'4��R���	��B��:��'W�=�'?&)�?��?^e?(�ɾtw�D�m��Q��2Oh�O꾴����;�*�6�T=�?x��d�i���վ����f�~���>�y]�?I7+?�b=���>�Ȕ�1c�6!ľ<�F>���$ �l��=�����=�Η=��t��G4��ѷ� �?���>oS�>~�;?"�Z���=���0�.n1�g���Q>�3�>�Š>~��>�,�;�)
�0��̾͘p}�ͯ���w>�Sd?��b?g6S?���2�X�e�Ʋ4� ���٧��>=9?���U>D���<a>��-3��&T�����A�/�j,��ڴ���=�:+?�i�>��>& �?&?I����]n��'�������>��?z}?W�?�-�>h�<J�C���>�/l?&��>���>�9��F� ���{�T�ŽK��>�J�>Z(�>ap>�(�hY[����������7����=��h?�\��.�b�0T�>*rR?$�;kCR<鷢>txj�P�"�ˡ���1�
>8g?��=)�:>Ȟľ٭�RI{��ڊ��r?>~?����F��Z�>��?,j�>$J�>G��?^�?ҍ
�����j-?Q?-�	?��
?N%�>��L>�6>(�|���K�����>>�>���}Į���>��Ͻ��ֽa�=��'>�@t<lK�h����jR==���MK�<��>Q�ۿ� \��������������zFn��y��Xa��x�s��;�K�9�u�B[7�����@s���p�{퉾�V�|��?�e�?n����#��Ԑ�n��=4
��v�>��Y��Qޥ�oҽõ��q���"��r�"���e���{�C�v�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾x1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@JoA?'�(��쾃HX=s�>͆	?'�?>��0�*!�������>P8�?v��?h�M=��W�f
��re?�4<��F�*���S�=��=M ==��U�J>�ϓ>�8��:B��s޽�q5>�>@�#�q�ސ^���<�]>H	սӕ�5Մ?,{\��f���/��T��U>��T? +�>R:�=��,?W7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?aD6?���>�d&��t�݅�=^6����|���&V����=[��>b�>��,������O��I��R��=)��Àο�E�DB'����̄=P�=�+"������=F�ݧʾ��&�)C�=�j�=�)�>)�>��Z>b�>��o?evB?���>rӐ>�_�� ʾ��Ⱦ��� ����޽,��:�)>)<r���:��x����־7�8���*���߾�=��#�=30R������� �R�b�^�F�4�.?�t$>��ʾ��M�)J/<vnʾ���?������1̾�1�8#n�˟?��A?*����W����@���m����W?\5�����מּ��=����@�=;�>�G�=��⾢3��wS���&?�? ^��k�B�w��>�eؽPr����(?F#??!r>��>�� ?_g���߽P��=�>���>�]�>���>�O��X;���?'`Z?�P��ٌJ��b�>A�k��m���s�2m�>j��090>�]���1��[Ҧ::w��dO?ߙ�>8#�p�<�{����ػ;��=sx?R�?���>�0F?�4'?��=��̾��J�;��� >:Jh?H�c?���=uB���-ɾK���L?�~w?J[>�z��&Ҿ�y���R���H�>W'w?��?{נ��Ar�/��F!���>?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������f��r���ȣ?}a�?������bm��q�s	���><^fS���=xL׼c����~3��������Ǿ�'��*��>�	@�K=���>��;���D�ۿ�`��nt��qF�&�!?�6�>��窎�Ϙ���*���XP��@_��3ƾW6�>�>Qʓ�������{��};��v��#��>����#�>��S��ŵ�@���t4<K�>���>z�>	��j*�����?���/+ο����s����X?�R�?�s�?$?I�5<D�v��{�����G?�Ks?��Y?�6!�H�[��#5�$�j?�_��wU`��4�tHE��U>�"3?�B�>Q�-�|�|=�>���>g>�#/�x�Ŀ�ٶ�<���Z��?��?�o���>q��?ts+?�i�8���[����*���+��<A?�2>���G�!�B0=�UҒ���
?U~0? {�e.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>hH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�$�>T�?�c�=�b�>|��=W��-�8s#>B�=��>�(�?.�M??N�>�Q�=�8�d/��VF�|CR���8�C���>w�a?�L?�Nb>~
��)�1��!�8�ͽ�p1�q�J@�l�,��߽�#5>��=>>0�D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*$"Ϳ����x]��!�Ծ�ܟ=΢�=��/>����EZ
>�;F=uk��}����=/$x>�>>�[�>�P>7�5>T�*>Ym���#�t$���>��@<L�
�����*�0��S�W:K����=;ݾKо�u���(��E_��6���)�cN�
��=n�N?�IY?"&m?���>�6��d�&>J2��
=9=`9 ���<��r>�/?<??[(?�٥=Y量^�c�����ݜ����yo�>��i>��>��>�k�>�ρ=?�`>�`_>
Q�>��G>�Y=�/��%�=V�>�0�>�J�>d��>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��w�T�4:>9����j�5`>�+ �~l���)��%Q>wl?��f>�u>a�3�!e8�q�P�v|��j|>�36?鶾�C9���u���H�cݾ�GM>ž>�D�l�o���&��ui���{=x:?�?�6���ⰾD�u��B���PR>5;\>QW=l�=�XM>�ac���ƽvH��g.=^��=F�^>\"?�->���=�S�>]0��1�K�#��>�E>�D2>d�@?��$?���䋽�=����/��s>���>gy�>+>@�J���=���>F�d>}&�},y��L	��0?�ܙO>�$���:X�*	d��;v=����IZ�={�=������=�'"=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>gx��Z�������u�y�#=S��>�8H?�V����O�p>��v
?�?�^�ީ����ȿ.|v����>V�?���?e�m��A���@����><��?�gY?coi>�g۾#`Z����>ͻ@?�R?�>�9���'���?�޶?ׯ�?���<��?8��?��H>����3� 5���ߞ���p���1<O��>wF��|7R������6��}-���@���^[�ݏ�<T�M=�z[>�l��S�F�
-��0,=I����'�;�Z�>�5H==v	�n%v>�?
�>���>Z��=�꽌;b�t�<���K?���?,���2n�O�<_��=*�^��&?�I4?Uj[��Ͼ�ը>�\?k?�[?d�>;��N>��E迿7~����<��K>,4�>�H�>�$���FK>��Ծ�4D�dp�>�ϗ>�����?ھ�,���S��FB�>�e!?���>�Ү=ڙ ?��#?��j>�(�>?aE��9��W�E����>��>�H?�~?��?�Թ��Z3�����桿��[�z;N>��x?V?nʕ>`�����jE� BI�+���^��?�tg?�S�1?:2�?�??\�A?q)f>ׇ�#ؾg�����>��!?�b���A��4&�����?�Y?���>rg���{ֽ�Ӽ��:Z���?{%\?�9&?;}�a�>�¾�$�<��"��M���;,F�ך>�t>F��qb�=��>
İ=�m�|/6���g<���=l^�>˖�=�7�{��/=,?�G�ۃ�h�=��r�9xD���>�IL>����^?{l=��{�����x��	U�� �?���?[k�?F��=�h��$=?�?S	?{"�>�J���}޾A�ྷPw��}x��w�Q�>���>#�l���I���י���F��,�Ž�%'���>��>?U��>7!>>�>�럾��!�;j�3
�YB`����5�|(���A���
�=��0��|û�L1���>/�/��!�>�;?��m>Ӓ>���>"<�|�>iat>�7�>\�>��>
�r>��>�u%=�:ڽ�KR?U���ǿ'�������3B?�od?D3�>O�h��������{?م�?�r�?^<v>�{h��&+�iq?�@�>n��qm
?V:=.��Y��<�P����sX�����'��>�Q׽:�DM�pcf��f
?�,?1����̾� ׽�5���>)&�?$��>-�X뉿�k��,��.Fm��_���5�a�J��0:�H!y��q��?$��ߟ��F�W�ay��K�?�b�?�d�dU!�VMʾ��@��8�=!{�>��>g
?�w8���;���O���R��*�ńm�"(�>U3?e��>,PD?�6?2Q?��O?��>ȡ>Jr���t�> �#=��>� �>7�7?S)?0�&?/c?��*?�f>y�Ž���<پ �?�?Dv?hX?��?!{�Z|�������<�Cb�H���E�=�
U<�Tڽ�8E�+̀=�S=>I�?�p��,:��N��:�t>�P8?U �>L�>k�������u�=���>��
?Ey�>�R��9�n����q�>�X�?n����<�'>���=§���(�^�=rnϼ���=�� ���S�x��;�W�=�+�=�o����G;>�<1%�<�t�>A�?���>mC�>�@��(� �T���f�=!Y>jS>0>�Eپ�}���$��g�g��]y>�w�?�z�?^�f=��=Ŗ�=}��qU������������<�?5J#?.XT?V��?d�=?jj#?�>+�cM���^�����ͮ?u!,?��>�����ʾ��ω3�؝?h[?�<a����;)��¾��Խܱ>�[/�g/~����2D��녻���o��1��?쿝?�A�L�6��x�޿���[����C?�!�>Y�>��>N�)�|�g�q%��1;>��>lR?���>&�O?�"{?+�[?)�Q>8�$߭�ː���b*��#>�??���?�ʎ?]ox?�a�>"> V+�[.�����=��Ev�Q����P=MPX>�j�>[��>,��>��=^�ĽH���r=�n5�=ʄc>���>E��>��>'Ax>�·<xB?� ?w��]�2�<���Ɍ��!���z?���?��%?�ʳ�3j��9����i��>&��?���?�e=?89���=D1!�t�ľ �w���>P�>��>��=�ѱ=��\>�ޱ>�͑>����-���C)C��(��t�?�J?��e>_ƿ�q���p��Ɨ�_d<����
e�Ҕ��[�u��=繘����F˩���[�����a���2�������K�{�U��>~|�=��=N�=�c�<n�ɼ0ڽ<-K=�<_�=�p��Qm<��8�+ϻ����+��ۆ\<��I=���˾�L}?�I?��+?r�C?�z>b�>.�/�0s�>4���А?]W>?O�s5��i/<�ߨ��A���44ؾ,�־n d�蟾�(>�6I��M>�3>���=Jǉ<{��= �j=�a�=/V��=P��=gܹ=���=]�=�e>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��7>�>^�R�#�1�ؔ\���b�YsZ�Q�!?�G;��M̾V9�>��='߾P�ƾδ.=�6>}b=�`��S\���=�z��;=� l=<։>T�C>�q�=h2��D�=?�I=���=��O>�ϕ���7�a,��3=C��=�b>�&>t;�>a�?w�/?v4b?w��><�z�1;������>��=�!�>�¡=!V?>��>�<9?�fE?�G?P�>X[=3�>@J�>e�+�r�r����©��K�<�s�?��?�8�>�5�;-VD��D ��6:��a޽I?�4?�/?Ł�>_V�����Z&���.��|��|%��[$+=knr��qU�=0��Ai������=9r�>���>(�>RTy>]�9>��N>"�>ۦ>%�<�u�=���q��<J�����=%�����<�
Ƽ��{�`%�H$,�PU���D�;<T�;� ]<�s�;}��=���>�;>)��>���=���B/>����#�L�+ǿ=TF���+B��3d��H~�6/��V6�p�B>�;X>Xy���3��$�?�Y>�m?>J��?JAu?~�>��{�վ�Q��Y?e�TS�ȸ=O�>�<��z;�4Z`���M��|Ҿ���>���>��>��l>�,�:$?�ыw=�#��b5�N��>}��%R��M�;@q��>������Yi�j��D?OB���V�=�~?��I?�ޏ?ŉ�>�Ҙ�mؾ�X0>�D����=����p������?�'?p��>M���D��H̾=���߷>�AI�H�O���ϰ0����`ͷ�Ǐ�>������о�$3��g������<�B�xNr�(�>�O?T�?�8b�{W��|UO����#���q?�|g?�>�J?�@?8+���z�Qs���u�=��n?~��?=�?�>���=h���!��>�	?��?/�?��r?;7�aK�>	[�;�{.>e��'O�=(9>h�=4�=s�?��
??�����	��%��ۆ^�L�=��='G�>��>��d>���=��W=n��=�_>���>�t�>r�f>֜�>*	�>���a���l,?L	>U6�>/@,?�߂>z�2=�r��;[�<6��i0=���aɽӠ���m
=�Į����<�d����>��ſ�a�?��h>����]?�/�Qޛ�k^>��k>���G�>��G>�?r>�T�>2ؽ>�>�k�>�A<>�FӾ�>����d!��,C�q�R���ѾD}z>����N	&����v���BI�yn��dg�vj�G.��B<=��ǽ<!H�?U����k�N�)����W�?�[�>�6?:ڌ���ɯ>`��>�Ǎ>�J��j���Xȍ��gᾬ�?5��?�;c>��>O�W?�?R�1��3��uZ��u�L(A��e�Q�`�p፿�����
�����_?��x?yA?�K�<,:z>?��?��%��ӏ��)�>�/�';��B<=�+�>*���`�;�Ӿ��þ�7��HF>��o?@%�?�Y?�SV�\��;@��=߫$?��2?.�x?^S0?]8?�|���^?�->�=?��?R�:?9*?(��>��)>�S%>G=Λ�=�� ���\;�k��{��ݠ�=�/>?�������ɽd0j=X�Ƽ�eM��=���:���<��=s�>u��= ק>z�[?,J�>�Ci>��6?a���u7�������8?���=4ߌ�}���t��}��ɻ�=Q�a?�Ѩ?G�Y?d��>u�A��T�k>И>"�>>�qT>%��>���D�K�/,�=Ś#>W;'>��=������ԓ����:���>���>�1|>P��x�'>q{��p/z�_�d>��Q�[ɺ�h�S�z�G�f�1���v��Y�>.�K?�?䠙="]�`&���Hf�5/)?p]<?�NM?�?��=^�۾q�9���J�U<���>@b�<8������#��f�:�`��:�s>�1��A���c>ce�@l޾�n�hJ�s�b(I=R��? W=N��h־|��_T�=D3	>� ���!�:���Ԫ��J?k=\M��M�U��h��\>�>�Ů>;��Eu�L@��鬾�Õ=�;�>|=;>��������jG���%�N>ߕ&?��Z?��?r�¾yg�Ә'�t�ᾫ�i���>8^�>'��>?0��=��>9���H\"�K�V��tU�A��>i��>#L��F��Ͽ�����M��X�>���>MX�>zn?�<R?�"�>�c[?�,?� ?t>#��;�\��?�π?K��=�-���ɾF�Q�#�"��
�>x�+?c���'>[?�k�>�1?��M?��?��=�.����F��;�>Y��>�PO��gƿ��V>��A?(��>Ek{?z��?���9%�3�����>�����>M�k?�^?�� ?z4?
����˾C�>�h]?t�?W�a?3��>�y�<T��R�?�~"=I�>W~3?�H-?��3?z�d?��.?G?t��;�q�nR޽,����1<���ܼ$��<3S0�(����&��7���@Tv�K��<:�=�:~<���<Z�ʻ��=��<�_�> �s>����0>�ľ*N��`�@>lv��vH��'Ԋ���:��ڷ=��>g�?r��>RX#���=���>�K�>s��d4(?��?�?�>#;��b�z�ھ#�K���>-B?@��=��l�������u�i�g=��m?;�^?Q�W��#��O�b?��]?@h��=��þz�b����g�O?=�
?3�G���>��~?f�q?U��>�e�+:n�*��Db���j�&Ѷ=\r�>LX�S�d��?�>o�7?�N�>/�b>'%�=iu۾�w��q��h?��?�?���?+*>��n�Z4�1
�L&���oO?ި�>"4þf�?1Q�?׾�q��m���]�u�w��4��'4��R���	��B��:��'W�=�'?&)�?��?^e?(�ɾtw�D�m��Q��2Oh�O꾴����;�*�6�T=�?x��d�i���վ����f�~���>�y]�?I7+?�b=���>�Ȕ�1c�6!ľ<�F>���$ �l��=�����=�Η=��t��G4��ѷ� �?���>oS�>~�;?"�Z���=���0�.n1�g���Q>�3�>�Š>~��>�,�;�)
�0��̾͘p}�ͯ���w>�Sd?��b?g6S?���2�X�e�Ʋ4� ���٧��>=9?���U>D���<a>��-3��&T�����A�/�j,��ڴ���=�:+?�i�>��>& �?&?I����]n��'�������>��?z}?W�?�-�>h�<J�C���>�/l?&��>���>�9��F� ���{�T�ŽK��>�J�>Z(�>ap>�(�hY[����������7����=��h?�\��.�b�0T�>*rR?$�;kCR<鷢>txj�P�"�ˡ���1�
>8g?��=)�:>Ȟľ٭�RI{��ڊ��r?>~?����F��Z�>��?,j�>$J�>G��?^�?ҍ
�����j-?Q?-�	?��
?N%�>��L>�6>(�|���K�����>>�>���}Į���>��Ͻ��ֽa�=��'>�@t<lK�h����jR==���MK�<��>Q�ۿ� \��������������zFn��y��Xa��x�s��;�K�9�u�B[7�����@s���p�{퉾�V�|��?�e�?n����#��Ԑ�n��=4
��v�>��Y��Qޥ�oҽõ��q���"��r�"���e���{�C�v�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾x1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@JoA?'�(��쾃HX=s�>͆	?'�?>��0�*!�������>P8�?v��?h�M=��W�f
��re?�4<��F�*���S�=��=M ==��U�J>�ϓ>�8��:B��s޽�q5>�>@�#�q�ސ^���<�]>H	սӕ�5Մ?,{\��f���/��T��U>��T? +�>R:�=��,?W7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?aD6?���>�d&��t�݅�=^6����|���&V����=[��>b�>��,������O��I��R��=)��Àο�E�DB'����̄=P�=�+"������=F�ݧʾ��&�)C�=�j�=�)�>)�>��Z>b�>��o?evB?���>rӐ>�_�� ʾ��Ⱦ��� ����޽,��:�)>)<r���:��x����־7�8���*���߾�=��#�=30R������� �R�b�^�F�4�.?�t$>��ʾ��M�)J/<vnʾ���?������1̾�1�8#n�˟?��A?*����W����@���m����W?\5�����מּ��=����@�=;�>�G�=��⾢3��wS���&?�? ^��k�B�w��>�eؽPr����(?F#??!r>��>�� ?_g���߽P��=�>���>�]�>���>�O��X;���?'`Z?�P��ٌJ��b�>A�k��m���s�2m�>j��090>�]���1��[Ҧ::w��dO?ߙ�>8#�p�<�{����ػ;��=sx?R�?���>�0F?�4'?��=��̾��J�;��� >:Jh?H�c?���=uB���-ɾK���L?�~w?J[>�z��&Ҿ�y���R���H�>W'w?��?{נ��Ar�/��F!���>?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������f��r���ȣ?}a�?������bm��q�s	���><^fS���=xL׼c����~3��������Ǿ�'��*��>�	@�K=���>��;���D�ۿ�`��nt��qF�&�!?�6�>��窎�Ϙ���*���XP��@_��3ƾW6�>�>Qʓ�������{��};��v��#��>����#�>��S��ŵ�@���t4<K�>���>z�>	��j*�����?���/+ο����s����X?�R�?�s�?$?I�5<D�v��{�����G?�Ks?��Y?�6!�H�[��#5�$�j?�_��wU`��4�tHE��U>�"3?�B�>Q�-�|�|=�>���>g>�#/�x�Ŀ�ٶ�<���Z��?��?�o���>q��?ts+?�i�8���[����*���+��<A?�2>���G�!�B0=�UҒ���
?U~0? {�e.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>hH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�$�>T�?�c�=�b�>|��=W��-�8s#>B�=��>�(�?.�M??N�>�Q�=�8�d/��VF�|CR���8�C���>w�a?�L?�Nb>~
��)�1��!�8�ͽ�p1�q�J@�l�,��߽�#5>��=>>0�D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*$"Ϳ����x]��!�Ծ�ܟ=΢�=��/>����EZ
>�;F=uk��}����=/$x>�>>�[�>�P>7�5>T�*>Ym���#�t$���>��@<L�
�����*�0��S�W:K����=;ݾKо�u���(��E_��6���)�cN�
��=n�N?�IY?"&m?���>�6��d�&>J2��
=9=`9 ���<��r>�/?<??[(?�٥=Y量^�c�����ݜ����yo�>��i>��>��>�k�>�ρ=?�`>�`_>
Q�>��G>�Y=�/��%�=V�>�0�>�J�>d��>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��w�T�4:>9����j�5`>�+ �~l���)��%Q>wl?��f>�u>a�3�!e8�q�P�v|��j|>�36?鶾�C9���u���H�cݾ�GM>ž>�D�l�o���&��ui���{=x:?�?�6���ⰾD�u��B���PR>5;\>QW=l�=�XM>�ac���ƽvH��g.=^��=F�^>\"?�->���=�S�>]0��1�K�#��>�E>�D2>d�@?��$?���䋽�=����/��s>���>gy�>+>@�J���=���>F�d>}&�},y��L	��0?�ܙO>�$���:X�*	d��;v=����IZ�={�=������=�'"=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>gx��Z�������u�y�#=S��>�8H?�V����O�p>��v
?�?�^�ީ����ȿ.|v����>V�?���?e�m��A���@����><��?�gY?coi>�g۾#`Z����>ͻ@?�R?�>�9���'���?�޶?ׯ�?���<��?8��?��H>����3� 5���ߞ���p���1<O��>wF��|7R������6��}-���@���^[�ݏ�<T�M=�z[>�l��S�F�
-��0,=I����'�;�Z�>�5H==v	�n%v>�?
�>���>Z��=�꽌;b�t�<���K?���?,���2n�O�<_��=*�^��&?�I4?Uj[��Ͼ�ը>�\?k?�[?d�>;��N>��E迿7~����<��K>,4�>�H�>�$���FK>��Ծ�4D�dp�>�ϗ>�����?ھ�,���S��FB�>�e!?���>�Ү=ڙ ?��#?��j>�(�>?aE��9��W�E����>��>�H?�~?��?�Թ��Z3�����桿��[�z;N>��x?V?nʕ>`�����jE� BI�+���^��?�tg?�S�1?:2�?�??\�A?q)f>ׇ�#ؾg�����>��!?�b���A��4&�����?�Y?���>rg���{ֽ�Ӽ��:Z���?{%\?�9&?;}�a�>�¾�$�<��"��M���;,F�ך>�t>F��qb�=��>
İ=�m�|/6���g<���=l^�>˖�=�7�{��/=,?�G�ۃ�h�=��r�9xD���>�IL>����^?{l=��{�����x��	U�� �?���?[k�?F��=�h��$=?�?S	?{"�>�J���}޾A�ྷPw��}x��w�Q�>���>#�l���I���י���F��,�Ž�%'���>��>?U��>7!>>�>�럾��!�;j�3
�YB`����5�|(���A���
�=��0��|û�L1���>/�/��!�>�;?��m>Ӓ>���>"<�|�>iat>�7�>\�>��>
�r>��>�u%=�:ڽ�KR?U���ǿ'�������3B?�od?D3�>O�h��������{?م�?�r�?^<v>�{h��&+�iq?�@�>n��qm
?V:=.��Y��<�P����sX�����'��>�Q׽:�DM�pcf��f
?�,?1����̾� ׽�5���>)&�?$��>-�X뉿�k��,��.Fm��_���5�a�J��0:�H!y��q��?$��ߟ��F�W�ay��K�?�b�?�d�dU!�VMʾ��@��8�=!{�>��>g
?�w8���;���O���R��*�ńm�"(�>U3?e��>,PD?�6?2Q?��O?��>ȡ>Jr���t�> �#=��>� �>7�7?S)?0�&?/c?��*?�f>y�Ž���<پ �?�?Dv?hX?��?!{�Z|�������<�Cb�H���E�=�
U<�Tڽ�8E�+̀=�S=>I�?�p��,:��N��:�t>�P8?U �>L�>k�������u�=���>��
?Ey�>�R��9�n����q�>�X�?n����<�'>���=§���(�^�=rnϼ���=�� ���S�x��;�W�=�+�=�o����G;>�<1%�<�t�>A�?���>mC�>�@��(� �T���f�=!Y>jS>0>�Eپ�}���$��g�g��]y>�w�?�z�?^�f=��=Ŗ�=}��qU������������<�?5J#?.XT?V��?d�=?jj#?�>+�cM���^�����ͮ?u!,?��>�����ʾ��ω3�؝?h[?�<a����;)��¾��Խܱ>�[/�g/~����2D��녻���o��1��?쿝?�A�L�6��x�޿���[����C?�!�>Y�>��>N�)�|�g�q%��1;>��>lR?���>&�O?�"{?+�[?)�Q>8�$߭�ː���b*��#>�??���?�ʎ?]ox?�a�>"> V+�[.�����=��Ev�Q����P=MPX>�j�>[��>,��>��=^�ĽH���r=�n5�=ʄc>���>E��>��>'Ax>�·<xB?� ?w��]�2�<���Ɍ��!���z?���?��%?�ʳ�3j��9����i��>&��?���?�e=?89���=D1!�t�ľ �w���>P�>��>��=�ѱ=��\>�ޱ>�͑>����-���C)C��(��t�?�J?��e>_ƿ�q���p��Ɨ�_d<����
e�Ҕ��[�u��=繘����F˩���[�����a���2�������K�{�U��>~|�=��=N�=�c�<n�ɼ0ڽ<-K=�<_�=�p��Qm<��8�+ϻ����+��ۆ\<��I=���˾�L}?�I?��+?r�C?�z>b�>.�/�0s�>4���А?]W>?O�s5��i/<�ߨ��A���44ؾ,�־n d�蟾�(>�6I��M>�3>���=Jǉ<{��= �j=�a�=/V��=P��=gܹ=���=]�=�e>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��7>�>^�R�#�1�ؔ\���b�YsZ�Q�!?�G;��M̾V9�>��='߾P�ƾδ.=�6>}b=�`��S\���=�z��;=� l=<։>T�C>�q�=h2��D�=?�I=���=��O>�ϕ���7�a,��3=C��=�b>�&>t;�>a�?w�/?v4b?w��><�z�1;������>��=�!�>�¡=!V?>��>�<9?�fE?�G?P�>X[=3�>@J�>e�+�r�r����©��K�<�s�?��?�8�>�5�;-VD��D ��6:��a޽I?�4?�/?Ł�>_V�����Z&���.��|��|%��[$+=knr��qU�=0��Ai������=9r�>���>(�>RTy>]�9>��N>"�>ۦ>%�<�u�=���q��<J�����=%�����<�
Ƽ��{�`%�H$,�PU���D�;<T�;� ]<�s�;}��=���>�;>)��>���=���B/>����#�L�+ǿ=TF���+B��3d��H~�6/��V6�p�B>�;X>Xy���3��$�?�Y>�m?>J��?JAu?~�>��{�վ�Q��Y?e�TS�ȸ=O�>�<��z;�4Z`���M��|Ҿ���>���>��>��l>�,�:$?�ыw=�#��b5�N��>}��%R��M�;@q��>������Yi�j��D?OB���V�=�~?��I?�ޏ?ŉ�>�Ҙ�mؾ�X0>�D����=����p������?�'?p��>M���D��H̾=���߷>�AI�H�O���ϰ0����`ͷ�Ǐ�>������о�$3��g������<�B�xNr�(�>�O?T�?�8b�{W��|UO����#���q?�|g?�>�J?�@?8+���z�Qs���u�=��n?~��?=�?�>���=h���!��>�	?��?/�?��r?;7�aK�>	[�;�{.>e��'O�=(9>h�=4�=s�?��
??�����	��%��ۆ^�L�=��='G�>��>��d>���=��W=n��=�_>���>�t�>r�f>֜�>*	�>���a���l,?L	>U6�>/@,?�߂>z�2=�r��;[�<6��i0=���aɽӠ���m
=�Į����<�d����>��ſ�a�?��h>����]?�/�Qޛ�k^>��k>���G�>��G>�?r>�T�>2ؽ>�>�k�>�A<>�FӾ�>����d!��,C�q�R���ѾD}z>����N	&����v���BI�yn��dg�vj�G.��B<=��ǽ<!H�?U����k�N�)����W�?�[�>�6?:ڌ���ɯ>`��>�Ǎ>�J��j���Xȍ��gᾬ�?5��?�;c>��>O�W?�?R�1��3��uZ��u�L(A��e�Q�`�p፿�����
�����_?��x?yA?�K�<,:z>?��?��%��ӏ��)�>�/�';��B<=�+�>*���`�;�Ӿ��þ�7��HF>��o?@%�?�Y?�SV�\��;@��=߫$?��2?.�x?^S0?]8?�|���^?�->�=?��?R�:?9*?(��>��)>�S%>G=Λ�=�� ���\;�k��{��ݠ�=�/>?�������ɽd0j=X�Ƽ�eM��=���:���<��=s�>u��= ק>z�[?,J�>�Ci>��6?a���u7�������8?���=4ߌ�}���t��}��ɻ�=Q�a?�Ѩ?G�Y?d��>u�A��T�k>И>"�>>�qT>%��>���D�K�/,�=Ś#>W;'>��=������ԓ����:���>���>�1|>P��x�'>q{��p/z�_�d>��Q�[ɺ�h�S�z�G�f�1���v��Y�>.�K?�?䠙="]�`&���Hf�5/)?p]<?�NM?�?��=^�۾q�9���J�U<���>@b�<8������#��f�:�`��:�s>�1��ci���� >o{򾺳��1X�>�F�����Y�Ȕ
�"��=
���V�:}����=>v�=y Ǿ^Q'� ��৿p�I?;�>�˾v���N��(�J>&�>�ɩ>
B=���M�6�1����>��?uԂ>���=��𾐩O�	�	�F��>\�A?��]?R��?�N����q�
�D�ϟ��B������5	?Ys�>�?a�@>�@�=�x��˅��de�c�G�`=�>��>g.��zK�忠�q�쾙�!��.�>�?�b>{
?t�O?c�?h�d?d,?�?�0�>gҽ7Q��`#?ޢ�?Q;�;�%"��Pl��{0�EyC�r�>)Y/?W�+�߄>1�>��?��3?��T?�?�B�=i���G�@�>�1�>�n`������;@>��K?��>Y�a?� �?��V>�07�?f�����<>tL>yT7?ʞ0?��?3�>|�?:�s>�B	?�5T?6�?�6~?!;�>D�����ʼ�H?Ǽ�=�.�>ù?D� ?qd=?�q?,{?껫>��<=�-�7GT;M�.=G,�=���<L��<��5:�5��K�C�F>~=��W=K��y�n���T�}��r&�Փ�=g�T$�>Rq>�=���?2>�xľ���[=>�M��e���D���qz;�f��=~��>�4?��>nQ&�Ɍ=xR�>'9�>	\��B'?/�?ٌ?5��;FAb���ھzNO�Z�>@B?X~�=�m�<1���Ju��p=��m?f�]?O_W������b?��]?�k��=���þ޳b�׎���O? �
?�G�R�>��~?7�q?N��>��e�b4n�T��,Ib��j���=�}�>+`���d��3�>Ý7?�Y�>��b>�]�=)p۾4�w�%y���?K��?�?��?\:*>V�n��1�Lc������N?%��>t![�L��>\��ܾ��"�xǢ�)���E���h����!�����o��q�����J�=�>��3?�`\?�iC?������ch������'B�b���P�$���A�b�<���=�4w��q"���zʚ�%A�;��J�(UP��7�?��1?Ÿ�Xu�>(!��(ܾD��D�=Ȣ�3�7��D�=�|�:A�=�<
�G��{��꠾�$?�&�>�R�>��?4�I���;��k+�M�8�T���LȐ>�Ɩ>+�V>�t�>�]�<Z;��9�@����b�t�� �u>�gc?�K?�n?���(1�`���$�!���.�c���'�B>��>y��>�W�����E&�V]>�)�r����}m����	�,~=m�2?C�>)��>0B�?��?�i	�����vx���1� .�<h3�>�i?�6�>'߆>*�Ͻ�� ��n�>�@Y?��>��o>z�Ǿ�e�ws�s�Z�x8�>Cx�>��>>�>i�}�r�g�)��B;����?��MO=fx?T�Y��w��$>S�S?��=�|�<�F@>�4��9��m�$��^{�&A>q"?LP�=�p0>%�ξ���ǋa�ޱ����"?�%?sO��&�A���>X�!?�
?V�>!qt?G��>�	��0�˻��?��6?C9E?��T?R�?ì�=Q�������
��m"
>���>d�>�t�;z]8<g^�=-�Z��≾>YJ>�o�>l��="�Z���	��t"=�79>��=0!�>�lۿ!CK�ܗپ@	����?
�\ꈾb����b��r���a��x���Yx�	��L
'�  V�A;c�͢����l���?�<�?6���/�������������;��>5�q��l��e��u(�������Jb!���O�U&i��e�O�'?�����ǿ򰡿�:ܾ4! ?�A ?8�y?��7�"���8�� ><C�<(-����뾭����οA�����^?���>��/��q��>ߥ�>�X>�Hq>����螾?1�<��?7�-?��>Îr�0�ɿc���s¤<���?/�@4.C?C�&�)��}:i=yq�>�$	?�`E>�%��5��?�����>�V�?�P�?��=�MT�\b��Ae?�Ԅ<��C�!�W;W�>�n�=�=]���A>H��>�z!�V�7�{�ֽ<}'>�>1<�\u���f��<4YT>��������5Մ?({\��f���/��T��U>��T?�*�>W:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?:ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=�6�⊤�y���&V����=Y��>\�>ł,�ߋ���O��I��V��= ��ƿ.�$��w�DI=Q���[���b����jU��'���bo�v��Oh=p|�=upQ>a�>�!W>15Z>�cW?��k?�S�>��>��Q���P	ξ���L���������;	����N�z�߾�	����P����ɾ�S<��7�=��Q�o?���{ �?�a���F�%D,?%�'>�ʾ�kM��q�;d�Ⱦű����s�I����Gξ��2�}n�i�?(aB?�����W�������
ϭ�W�W?�Q���G�����)�=�����5=�3�>�p�=��߾��2�V`S�T*?0�?#E�TP����>�X8�@Q�=5VP?(��>�n=+	�>* ?u���bx=��Ϙ>�T�>o�>� �>j��=������9�M�8?�]?����<�*�7��>�a���jɾZG>s��=�^�
��< U>%�t=R���2&�N��qYN>.X?:w�>I(����3���^��H=p�x?Wi?m0�>DEl?��B?Ld�</��R���
��9~=ȠX? �h?��>r�h���о~���)P5?�Td?>EK>|�j��*�A�-�2����?�n??xE��ѡ}��쒿�L���5?��v?s^�xs�����I�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�%Þ?��@���?I�;<��Q��=�;?m\�>��O��>ƾ�z������2�q=�"�>���~ev����R,�f�8?ݠ�?���>������\=�=��5X�?��?h��ݨk<%��5�k�«��D#�<sv�=/���w!�T��N�7��ƾ�
�6����e���ц>�[@�Z����>Ǡ8��0�JϿ����0о�q�ǻ?cz�>�0ǽ僣���j��Vu��G���H�[����Ï>A�>�+�G'���f���+�����6`><+I=K�>s&i�f��G�n��>S��>��>;��=����t��0֔?;����׿.9����`C]?_�?iY�?��??�u|<�
������=��j?�j�?($s?_A=ێ��s�Խ%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�Z�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�u�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�[�_?)�a�K�p���-�n�ƽ�ۡ>��0��e\��N�����Xe�
���@y����?L^�?h�?���� #�f6%?�>e����8Ǿ�<���>�(�>*N>�H_���u>����:��h	>���?�~�?Pj?���������U>�}?L3�>c�?q�=�b�>os�= 氾^W,��l#>;��=��?�1�?z�M?�Q�>Zq�=��8��/��UF�n<R���k�C��>q�a?�L?Mb>%���I2��	!��Qͽ�r1��輸K@�I�,�'�߽ 5>��=>�>1�D�oӾp�?Yp���ؿ>i���q'�D44?쵃>e�?Z����t����;_?�y�>:7��+���%��yF����?	G�?��?��׾�Q̼L>��>?H�>�ս �������7>��B?�'�D�� �o�{�>D��?~�@Fծ?Oi��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?}Qo���i�B>��?"������L��f?�
@u@a�^?*E䬿Ϸ����_���l��P^>,��=XLA>����I�=�k�;:��<�dX<t�="�>�`>�u>CRN>)�>>�h>q������O���,���3A�D�cp/��>���Ծ�3O��5�<󝾡*�����|�y�a������X���B�6��=|�U?�R?�p?Џ ?^vx��>j���n.=�{#��̈́=)/�>*i2?�L?��*?�ܓ=襝�j�d��_���A���ɇ�L��>�tI>�~�>YL�>�&�>��=9��I>q2?>S��>�� >�k'=���e=N�N>KM�><��>�|�>��>>s�'>-���P�����h�O&p��VȽA�?�+����F��7����3ǲ��M�=9J0?͓	>�
���cпc���kG?�@��W���s0�Qz>�0?V�Z?�)>����(��>�p
���m�v{�=����Qa��!���X>�4?�f>S�t>Ν3�9X8���P�8~���|>b$6?_���Ѣ9��u�S�H�hOݾ"M>Ϣ�>��G�:o��򖿲�~��ci�]�z=r:?�?򘲽Pⰾ��u�X\��U4R>*X\>�=�k�=�=M>�ac�<fƽ��G���.=]��=Y=^>x�?M0>�ԕ=��>݁��yB��>V�Q>��>�;?��'?5�߼��G�v�T�!���x>Z�>��>{�>�1?�.�=��>5wb>���ml������I�\1O>��f���g��8q�L��=a��*��=~�]=)����.�8<;=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�,�>�e�=J�������u�X�"=0k�>-H?m&��J�Q��M>�@�
?��?��򾥩��0�ȿ"}v���>�?��?��m�?����?����>F��?6Y?�.i>."۾]([��I�>ߟ@?R?� �>�$��'��?�ζ?T��?č3>�?nnp?&�>���T�.�/ױ��͈��z�=ҵ�:�ډ>��>�˾�.I�R���މ���j�
����~>07=�Ų>q �������=������_�&��>�VA>��3>{՝>?CS�>a��>!�<"���(~�����ZD?�?޹5����QEO��>����z�>6`??���=�W���ǘ=�HQ?��?��h?���>�(��eA����� ���� �=G$>R��>�d�>lMO:��>؂��#|`���>���>p�<BF뾇y��xtʼyG�>�hK?�  ?�9�=4� ?�#?��j>N!�>RdE��8��%�E�ܲ�>���>�F?��~?� ?�۹�
]3�����桿��[�/N>p�x?�T?ƕ>Ҏ������nD��1I�4��k��?Wrg?+��< ?�0�?�??V�A?~%f>��`ؾ���m�>�!?(��٭B��M'�{H�B�?D\?A�>������̽��� ����9�?#�\?�s&?��Ba�f�ľ��<�
�j�c�˖�;���8�>G>3s��K�=<7>��=_ij�`�7��^+<�=�2�>�,�=��2��,��0=,?{�G�{ۃ���=��r�>xD���>�IL>����^?kl=��{�����x��	U�� �?���?Yk�?b��C�h��$=?�?R	?i"�>K���}޾8�ྻPw�~x��w�Z�>���>]�l���K���ڙ���F��[�Ž�%����>��>�?���>y�C>��>t�����$��	�����\�e���R9���.��Z������7#�5���m���ez��Ę>y~��'b�>T(	?�Sa>��l>���>|�>9�>ƃD>~�>��>�^>��:>�\�=�̶;(�qR?˃����'��^辗o���'B?0fd?�2�>Cl�ˉ���r�ք?���?�n�?=Dv>�_h��+�x�?w0�>�����
?I>9=�S��=�<�=��������Č��o�>�H׽��9��L���f�~A
?_?[b����̾�׽5ܾ�b-�q?Z?!�&��Fl�uTu��QT��y1����������c�B'�7}j��o����ꄿ�����=�z?�l?���Dm �������X��s&���U>h��>;�>�=�>a`>�n��U,���^��&������S�>Ͱ�?��>,�>?�1? cJ?��K?�B�>>�@���Y�>S`=r>f�>�j??��"?c�2?�9?�71?�}/>
>ý�D����ܾ�t?�W?Z'?��?�}?'�����7�N�;�����4���'�8��=�= .	�ˋq��
�=��`>O�?X��X�4���'q>7?��>�Y�>�������<�C=� �>`�?ݔ>������o�'I	�\3�>�t�?�߼�%-=P�">	��=��R��a�����=�^�y�=.]ȼs3��
�<���=�3e=��c�� 5,�>��YC< u�>6�?���>�C�>�@��/� �c��f�=�Y>=S>|>�Eپ�}���$��v�g��]y>�w�?�z�?ͻf=��=��=}���U�����H������<�??J#?(XT?`��?{�=?_j#?ϵ>+�jM���^�������?� ,?É�>�����ʾ��ى3��?�Z?z;a�ϼ��;)�X�¾��Խͯ>�[/��/~�����D��ԅ�n��������?���?�A�:�6��x�꿘�5\����C?S"�>AV�>��>��)���g��$��1;>���>R?�#�>t�O?�<{?˦[?�gT>o�8�z1���ә��F3���!>;@?���?�?py?�t�>f�> �)��ྒT��c����HႾ�W=$	Z>h��>�(�>9�>C��=�Ƚ�Z����>�a�=�b>[��>���>��>��w>VK�<��C?�?e��e�vّ���C�~�<��b?�{�?�J6?u��;8� ��G>� �ݾ ��>ț�?
�?�� ?YȒ���=����� ���/�50�>T�>l�>V˛=�%<�.�=ճ�>M4�>���t�!�%�;�s~���?��J?a5�=�����
R�𵾽[��Xb��T/о�Y��>��!L ���=�����u]�f�m�Ծɞ��d����ƒ��c$=�.�>�)�=,�=��>�q�=f�=
D<ΰ�;7H�_��<\�=������<uy�;�Ԅ=��)=]��E�׼��߽5�˾�}?�;I?ӕ+?u�C?�y>
;>��3�V��>�����@?�V>ڞP������;�Z���� ��M�ؾ x׾��c�ʟ��H>,`I�>�>�83>eG�=�K�<%�=&s=�=R��=$�=�O�=dg�=���=��>*U>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>o�8>�>��R�Fz1���Z��a�Y�X�܀!?A�:��̾/�>#�=C	޾K=ƾ��1=Ǣ7>םi=����\���==[~��?=��s=*�>|�B>wT�=��z�=l&B=��=�'Q>��_�-=�3+,��4=|��=�Ga>��&>q �>]l?�:2?!a?/��>�Y�+H��|Q��H0]>���=d��>7ͬ=̇k>[�>�5?)@?��K?�[�>9��=�,�>]:�>��,���i��/�gĮ��I&��y�?��?�͵>
�}0�s��-[9��u��>%?��?H��>�U����9Y&���.�$���|4��+=�mr��QU�M���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=$�����<�vż���u&�:�+�1�����;r��;B�]<]��;�{�=���>�F>��>�=��� %/>稖���L�鶿=oG���B��:d��M~� /�=�6�'�B>�X>�؃��+����?u�Y>�?>(��?r8u?��>s�(�վ�V��de�8S�SS�=m�>Z�<��z;�DT`���M�ǂҾ��>�
q>0��>=i>�,���<��ӻ��׾o5����>�ޠ���<<\���q�U������j�i :��D?����n�r=,�n?��P?��?U�>��̽���ۘ:>���� =t�#���K��YO�ds?�!?ԏ�>Vxپ��P�x����"��X�>�a�6�e��>���/��aX�nх�y�>��;�_����F�0Ѓ�������J�����N�>�]?_��?^�$�m�b��Q��]'�ݴN=N�?��_?L�>�s?>�?���8
�����s>��g?g�?|h�?&{w>;��=]����<�>��?�3�?�M�?�	w?�%����>4s��D�8>�h�����=3>w�=V{
>?$�?(�?�����q���0o�"CH�-�<��=�m�>��>Jf>:��=?v=���<��U>�K�>�>�HJ>�K�>H�>������e#%?�h�=,��>�?1?r��>�!`=nŧ��X�<7Q���=��B&�����OB߽��<��q��B=���-�>ڴƿ,5�?,�Y>h����?Y"�8�T�H>�wZ>��ؽ�M�>J�C>��>���>ֶ�>0c>xߋ>͚!>c��,�=�l�,h��$=�Zo]��-㾜lW>>���� �'��2�ý�pQ�����=���l�����{O;�G6=w��?cB���d�B)+� �A���>B��>�
-?=���YJ�Y��=���>KK}>!���)����w���W�C��?���?�9c>^�>/�W?N�?��1��3�MvZ�ٯu�F(A�Ee��`��፿朁��
�[��?�_?
�x?�xA?-C�<;z>D��?��%��ԏ��)�> /��&;�y<<=�+�>s)����`�/�ӾT�þ�3��JF>�o?�$�?�X?�UV���^��r(>w:? �1?Vt?J�1?��;?�����#?3�0>:�?��?�s5?_�.?��
?�1>�a�=��[�e(=�"�����vѽ�oɽ��pO3=D�w=�3ƺ/
<X =�~�<ޑ���伝��8�����Ŭ<�h;=�F�=��=�ݦ>�]?=��>cm�>t�7?�(��-8������.?�;=�R��Lˊ��6����	�><k?6��?� Z?eAd>��A��WC�_>͝�>�B&> �\>^�>P���F����=�>��>8`�=�K�����'�	�p�����<V�>d��>I�|>�+���'>�좾��y��yd>��Q�������S���G���1�uov��G�>F�K?}�?`��=�@龋�����f���(?~*<?:M?�?�~�=`ܾ:��J���H�>jϬ<~��W���5����:����8�Ss>����6�۾R�>��-�$_�ؗj�_�Q�e�@��oϵ����=uP����n-���>�␽P��m#��φ��Ǖ�K0?�-������Q�'��� >(�a>x �>b�PK���*�����%6�>���>�3~>L�<Eվ��D���Ӿ��>�D?ш_?���?�j��E�p���A�	B��΅��L�ü��?���>(�?��>>o�=i������)?e�K�F��w�>M8�>!*�X�F�5����3��M_#�~�>�[?#�>
�?��Q?��	?�`?�<*?=�?P�>���@���B&?ׅ�?cd�=1"ս��T���8��E���>}V)?FC��З>
v?9�?��&?�xQ?��?J�>�� �T8@�%��>yi�>��W��Y���_>t�J?���>rY?'؃?�G>>Wx5�e������1y�=w>>��2?v #?��?���>�c�>u���Ho>���>12V?�e?��}?��ἇ��>9�>	�?���>�l7=�O�=�2?��b?�P?`A�?��:?)rE�k�=��޽ѳ���Z��Y �=�2N�sv>9��=E(�p�{=�m���B�=��=��"<�0��������u>��>�=l>����q>]�˾���5%2>�.�w��� 냾��4�Ǹ�=Z({>!�?���>�f�H�=#S�>)"�>���y*?��	?jY?]A�<�>b���ᾍ�h�=F�>��<?;3�=<lc��h���Xp�&c�=4(m?}F[?c�T�@:����c?k�^?L[��H�;�]��6�`����cO?m}	?pM���>��~?�-r?���>�f���l��Ü��/a�G�i�G��=S��>���c�+�>�;7?uC�>ok^>���=]|ܾ��v����?�Č?y��?M͊?��->�m���޿��	`���Y?���>���>[d�,��6�g�{����y���t���ˬ�J�������΍���¾��E����<\Xh>o�;?۟U?K�a?!=�����s����8N�p�����=���4��4���r��9��	��?��KM���T��]�~"�?eO?f�G��>�����:�������>��>�����7<��'I=,C>���l*Y�o���Q�?�q�>>��>M�?�t@�~P8��)��3�3��ka>0��>�ˬ>#�>}k9>�%+=ڬ ����G�Ͼ#
��:*u>�c?��K?�n?����v0�LT��{�!�\�?����*D>��>E��>��W���4�%��5>�V�r�x��t���
���y=g]2?��>�Ҝ>�:�?:�?W"	�p#���w�T�0��v<�¹>�;h?1��>B�>O�˽|i ���>��l?ʫ�>x�>ӎ��W!���{�~�ʽ��>٭>���>��o>ީ,�l\�_i�������9�lu�=]�h?ۄ���`���>$R?�O�:�G<g��>��v���!����'���>�z?�>�=`�;>}ž�!���{��0���s+?-f?����w%��h�>�!?��>Y��>Sh�?�r�>���9����6?sa?�wG?U�>?���>^==�3��
ͽ������=2�>�\>��`= ��=�����U��v�� =��=3l��Nћ���+<$?|����<2�=��;>L'Կ��I������T���%�l�q�R���L��mJ�����)���9J��3S!�����xB�i�t�~�k��O����?].�?�劾'a���x��>�}�J%�����>��'�Uͽt0��>����}�|�Ǿ酯�
�."?�H�f��Z��'?����ǿQ����7ܾ ?%> ?Шy?�-�"�i�8��� >�w�<�g���������*�ο�����^?&��>�C����>���>N�X>�Tq>���=I-�<��?E�-?���>o�r���ɿ����J��<t��?x�@8bR?���$0����>̫?N	?Z:#>i,��)�G{𾛆�>yu�?T��?w�=X"T�v?Z=\�l?Jbл�7���K��l$>��>�Z�=m&��+>v�>o[ѽ�B^��&ͽ�0�=225>R>� u����bVg<�n>���u���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=t6�剤�{���&V�}��=[��>c�>,������O��I��T��=�������!��V"�*�*�s��q���P�½-��H,��BN���e��6K���1�=��=�_U>_��>Hg>��Z>m7R?��k?F��>��>!ǽ%��gݾ�N�|���3�;d��-?�N��� �۾�7��N4��6��.�ɘƾ'?&�G_>��U��G���6��U]���>��-*?�-W>[�����4��}Ͻ�Jk�^�W��}��&�H��Q�kQT�Xn�?�<?0P��h^I��Z�ǅ�<3���&r`?����O��v;��L5>íE<�%�;�p>Nc�=J�¾�I,�׺)���O?�dC?�����S�>\<l��Z�ű$?cf�>��x�-�>�?�=��=��>`%a>l°>-�>��	>���i���~'??d�I?Ia˽�'��ڪ�>�����&X�/T]=
��<�/F�I$<	�c>�|��%�J�no�=WS��K<~YY?��>%|,�T�;*��$���h,={�x?��?(��>�!m?�7C?a�=�F��T��E	�e=�3T?үe?�a>�t}�C�׾x���L5?��d?�	G>o�g�+'꾀�.�n� �7?w�j?�?&���az��~��+��J�3?��v?�u^��o��y����V��>�>b�>���>��9��h�>'�>?��"��H�����V4��?��@.��?��;<<!�竎=�9?�Y�>]�O��?ƾ����g���'>q=� �>�v���`v�����O,���8?��?���>\������+">���A�?X0�?d������<Qi��O\��Zؾ1�M<��=Q�:��/Ѽ�
5��l������%��@��<]ʧ>��@Ϯ�Lq�>�57�H��XͿs�o����8�����?�r�>��ɻ��� h��G{�^�M��O��L��.6>�,>�%�(ξ/�����R�����>'��=o]�>x�Ϫ��?���(�n=�%>B��>���>����6��?�����eͿgw��/���o?q��?s1�?&�(?W����O��ݧ��Ij����>?�vZ?��Q?J�S��\[��>&�j?�_��wU`��4�pHE��U>�"3?�B�>S�-�$�|=�>���>"g>�#/�x�Ŀ�ٶ�9���X��?��?�o���>r��?ss+?�i�8���[����*�X�+��<A?�2>���G�!�A0=�TҒ���
?U~0?{�d.�Z�_?+�a�D�p���-�j�ƽ�ۡ>��0�f\��M��$���Xe����@y����?N^�?g�?��� #�g6%? �>o����8Ǿ��<���>�(�>*N>|H_���u>����:�i	>���?�~�?Rj?���������U>��}?$C�>sV�?�9q=��>s�>�5���$�M�3>O�=���3�
?uSH?:��>���=�E���'��6D���H�>����@��{d>lA_?�EC?��L>�렽S�ü[#����e��y(����$��O��Խ9\X>#�E>+0">CK��#����?Hp�8�ؿ�i��p'��54?,��>�?����t�����;_?Nz�>�6��+���%���B�]��?�G�?=�?��׾HS̼�>4�>�I�>F�Խ����X�����7>.�B?f��D��p�o�w�>���?�@�ծ?fi��	?���P��Ea~�	��w7����=��7?�0��z>���>��=�nv�ڻ��O�s����>�B�?�{�?	��>�l?��o�D�B�_�1=)M�>Ük?�s?2Oo�|��B>��?#������L��f?�
@xu@Y�^?A˿e���c���p���I�;؎�<"�->������=כN<��$���<X?�=@o�>��R>�wL>�! >���=!>�k��12 �80���u�� `�X?�E��n������}l�����Ͱ��;ľ�ٵ����je�����Ji�i�m�>>"mZ?�]?�,c?�F�>����u�(><�˾�I��[�~� >Fb>e�"?�>P?��#?��<]
���D]��Bk�����s�����>2+H>QP�>E��>��>"�W�鲀>�|>��~>��
>:f���\��L�=�ݵ=o�>O��>��>�/>Nh>p���򰿱�d�.W��]$ｲ6�?`���C�D��V��B��䫾7�=*�,?��=�T���*п��D�E?&�����%��4L	>�h0?��V?7$>�~����Y�� >彪Nu�0��=b����lj��)��ZI>N�?]��;��L>}�I�:4d�?/���,��;�5H?Ҏ�n\]=C���N	]�l�����>�K�>c5��+7����9�L�6C��oҽE1O?�#?Yͮ=ce��䭣�t��(�>7�s>z�N<e��>�e>�1��L�(=�:ܽ�$=P�P�V�?>jw�>�>�o�=J�>h���T�sT�>f�^>0C�=�,?��*?�T��i ����e����V>��>�Co>T>�p#���=<��>�GF>j��o��A穽~��c��=Hf��G3��򯼥N�=����(�=^��=�"�JUK����<5�~?���}∿��^X���lD?2,?��=��F<�"�����LE����?��@�m�?�	��V���?�?�?
��^��=�{�>F׫>uξ��L�D�?�ƽĢ�\�	��7#��R�?3	�?�0��ɋ�:l�.:>�_%?_�Ӿ�X�>ed��\�������u��r#=��>�3H?�B��m�O��>��l
?$?�N�\���R�ȿjxv����>�?�?��m��@��	@�d��>���?�hY?�ji>�i۾V_Z�소>�@?�R?W!�>�5���'�[�?Iض?ѱ�?9I>��?��s?Nk�>@-x��W/�:5��%����,=f�[;1f�>q\>�����eF�	֓��f���j�n��	�a>!�$=z�>�<佣2���&�=�����C����f�E��>�0q>�I>OV�>d� ??`�>⨙>8I=�z��g߀�������L?׏?|K�F�l�w\�<p�=�b���?dJ3?t����˾�>��\?ɝ�?d*Z?��>�%�N����﾿-���W��<�O>�2�>]��>OQ��h�K>��վhA�QJ�>QQ�>����҄׾�7}�Z�G9��>�;"?�<�>A��=v
&?�(?�fi>ڕ�>ז;�Yj���F?��<�>���>�%	?�|?m�?,�����*�������ZBV���L>��r?bV(?@^�>U��A��<h����|ݽq�?�L?ӈ*�֑?���?�bD?~@?��@>¤���ݾǧ��CJ>` ?�=�)�;��7(�`�'��?=�
?|_�>�����j���߻�Y�&���G?6�[?GJ?o>��>�V�t=��=z=b�m</䟼�)ͼ؅���"->]J$>9(��Kw>��R>���=�����U:��&�<!��=^]�>op�=���K�M�c8,?z?O��Y���A�=�!r��C�o��>�qK>避�3^?.�;���{��Ҭ�H��pU����?ra�?�W�?hW����g���=?f�?X�?:�>Vΰ�F߾�}߾Zx��;{���֨>���>l�V����������cD��P�ɽdm�P�>���>�>_<�>D@�>�#�>�*n�i�0��R;�*��8�9�1�5���9��	��n������%��*༐�퉗�#�\>a�H�u�>�{?�~_>���>��>��T�j��>�><F>�zU>�M>t� >C`>mC�=Ϊ�"R?n����U'��e�98��)B?�Ed?���>�Fi�	}���w��P?PR�?�W�?��x>�g��"+���?���>p���	?�V9=Ԛ����<*������!����~`�>ܽ��9�M��8g�-[
?�
?������˾+Rؽ������<�	{?{�=?5�U��{��Ӕ��x�~���7���/<�ѷ����]�n*]��-���Н��2����L�-C`���?w�a?^���g澑SZ�EWi�U�Y���<�>k�>�7�>v<<>y3���<��]^��	��0�OM�>y�?�[�>��L?L�;?��P?e�K?�.�>�f�>䢦�$��>s�X8�`�>"��>�49?�\0?�i,?aI?��)?k�[>~���W���tվ�?��?�?(��> ?�����?��� ��+�a'n�'1��
1a=�6�<��ֽ9�{�6�l=]%\>�_?Iq�/�8�I>����j>Dp7?���>��>KZ���u���t�<���>�
?|��>�4��*Ur��5��>c�?w7�|��<�6)>���=�[����(�=,ü/א=�ه���9��� <��=��=g��Z�:��,;f֍;	�<��>ϳ?y��>�-�>����^P�������=o~[>��Q>i�>Y�ؾz0��\ߗ��g�~�{>�9�?X'�?�Y{=��=��=�����_�����۶���m�<:�?j�!?��Q?��?	5>?�$?G
>����m���f������?�v+?�1�>���P�ʾ5˨�u�3���?�^?��`�^���)��[¾Ϡҽ��>�,/�?~����WD��Y��d���0���{�?5ѝ?|�@�X�6�^��V���0����oC?Zu�>���>��>��)��g�XE�':>�,�>U�Q?wE�>!I&?ˑ{?SP?&�n>H������G��m��M=�v6?��z?h��?-��?�	?�iU>Հ���|�([����<^Ok��kw��=}�>���>���>"�>��'>�vɽ0����A���ِ�I)>��	?��>�N�>*� >6c���G?���>/������h8��NR���-��Nt?�@�?[�*?�=���GF�C�����>�;�?���?�e*?#�S��v�=��Ҽl����p��l�>�&�>�t�>>�=+B=J>3B�>�'�>�5��~���8��K��<?�rF?LO�=���z>h������Oפ�OUf�Σ�w�;;oQ�+�t>՚[��S���6Ѿp�x��9��}D���ڵ��~H�S ��J�>y^=�_=Q�<x�Ͻ.�<��2�$��.2=8�r��+��н�wX;��='A�|+>�>j0�=� 2�ƺɾ6�}?�.I?�+?�^C?P�y>��>C.���>vہ��z?�NU>:�Y�~��C�;��+��������׾��־�1d��B��#�>RiF��>1L3>x_�=!b�<���= �|=�q�=����o�=!f�=ȹ=G��=�`�=e�>hW>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�??ti��d�>M���㎽�q�=J����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��>���>��M��y�V{(���)O��ݩ/?��W�i@�;A�>�:3>l�����׾wg���$>��=x�A�r�2����=J�����x��_>�G�>��=���}Y>g�<��m�(1=3�����;@�>��=ʷ�=�̏>	�B>cL�>�?�0?-�c?=/�>	]k���;�z��hǋ>8��=�Ȱ>A�=ؘA>�#�>t�8?�mD?��J?%Ѱ>}��=��>�ߤ>Z>,���l��㾨󦾉��<�.�?2��?��>��
<��@���G�>�U�ĽI�?�1?c�?���>=E�\��@O&��.��㛽�㪸�.+=�#q��S�|����[�B�4��=�f�>��>�>��y>I�9>}�N>��>>h��<�݅=>o�����<�����x�=Q������<2Kļ��c����(�$;�� �;��;�e`<q3�;��=S��>�>���>wf�=�_��_v->�{����L��a�=F����~A�$Bd��0~�Sf.��5�01B>��V>ٟ��R둿�G?\�W>,�?>�-�?QUu?��!>(����־'F��k f� eP�8c�=^T>�v@��I;��`��wM�!EҾ�W�>`@�>��>�,r>b�.���A�U\=`��/
4���>+ɐ�4e�4��4p�����q��(ck��?��AA?!R����=}|?�IJ?iԎ?p��>˪���yݾ$,>$�|�� =��R�l�����=?Y9#?{��>��H^F�b��[�ýe֥>��J��\��'���K�Q�(��@��_g�>���Qx��&��ép�ms��s�I�b�� �>�?[�?�*����@��!�H7��?'ws?o�>(k�>C��>��ٽ5lپa�'����=9�}?%��?W��?�%>�'>����/?��?�I�?´�?/�?/������>Cz�<�R]�B�=��,���{>�Xa>Ȫ�>`?D��>��M�7����1��6����(��ؿ���w=f�P>��>D��>+>}>)��=��H����8��,=��e>ҡ�>l��>��~>+]����f�?l��=��>�+?�1�>3w��2xսX�0=�%%��x��G{�-��t�>=�͠<J�½I�`;�N�;iz�>�J���Ru?�A>M�Ѿ��?<�����H��#J>�1>�(L�s��>���=fA�='B>�?�>��9>^�>�ּ=� ��8>��]@�o�9���S��J ��A�>� �w3'�y�[�'���4��o���	���\��Sa�=�'��=�<��w?G�=xY��q���J4��h.?�*	?D�?Nhþv�ν .>���>�-�=��ܾ����a���z��v?ۘ�?�QN>Q��>��U?�?II�i�A��D[�TAo���:��.^�Ka[�z.����+����ֈ_?�z|?�b@?Ľ�<`�{>)߁?���ט���=�>o 1�^�>���;�Q�>�T��4uS�M�����̾�����l>�rp?F�??�/X���D���">dq:?˲1?�ct?@C2?\<?�[�/�$?v�:>�?��?�3?6�.?�w?�5>Z+�=}q�k�U=�r��'̆���Ľ��ʽ����=
0�=��;�h�<Bn=���<n��C켝CY<����u<|�B=�Ƞ=6��=�E�>E�i?w{�>�z�>��7?������K�F��8�>���}ݘ�;%Y�(k\��_;8���d`?jk�?��5?��9>F?2��� �н�>f�>�>�)5>�>9경c�Z�>k*>��=��q��D��y�k����^|�����<[�=k��>!v@>�r�.�4>�����T�,�>g.o�7料�tP�\N�q%��9n�i��>�T?�w ?	H+=?|꾈#�Z��?�6?��K?l�?2e�=���9��DC�� ���|>i�={.� #��{���xe2���=�"�>Bԧ�Χ׾*R�>���}�$��j�L�^��y�5~��e(���E>[Ǿ!���ž/���ġ�d����8Ԟ�:��-
-?-&�=kk�d���ž�q>��>�֬>�=Q>����M�����<�?9>(��>�����^�D��u����H>0:?�iU?m�?�u���I��(�Ǿ�����Z߻�@?�b�>�?��q>�I>����<�&�N�,���>��R�>u�>ㅰ��gS�Lݙ�d���g�⾡��>��?��=�%?�W?8�I?%��?�L,?q)?��>�'�g��`]$?�À?0q�=�?ƽ&~R��U7�iU?�}C�>��?��G���>8�?7�$?��)?xCR?��?ʃ�=���7��l�>K
�>��N��`��[Y>ڡU?���>�`?炅?�/>|�.��A���n�����=��>��;?��-?�	?�~�>K	?�Ԟ�k�<�Y�>]Ma?p�?�2}?���><$*?t<U��k�>���>�x�><�?�1+?�U?su?��V?��$?�	�=����_�H�ˉ=�>��=�3��Gƅ�+ҽ�i��C�=iU���+��6�ZD���$'�{��a�e=IA= R�>��s>����1>��ľOJ����@>+{��<I��V�{�:����=�s�>h�?«�>�f#�w|�=֖�>^:�>����)(?}�?S ?��3;��b�A�ھĉK���>� B?N��=?�l� �����u��h=9�m?#�^?@GW����O�b?��]??h��=��þ{�b����g�O?=�
?4�G���>��~?f�q?U��>�e�+:n�*��Db���j�'Ѷ=\r�>LX�S�d��?�>o�7?�N�>1�b>)%�=iu۾�w��q��h?��?�?���?+*>��n�Y4࿹���`����i?`�>�lk���?�=�6E���1a�A��m�ƾ$n�����'EV�\1�����p����[5�N�=���>-S?5?Hb.?���ܥ��ֶ������Y8�ݶ��=�V�*/F��s)��0n�(�3��"�Gz����.Y���A���?��'?�0�Ù�> ͘����;��B>𤟾2!���=8\����?=�Z=W�h�D�.��X��l ?�&�>P6�>��<?��[�cF>���1�8�7�������3>�բ>���>w;�>���:�>-���Q�ɾ���Խ��m>�T`?,F?vn?,b�Y�/�B瀿��#�u�6�Nԯ��!>I�>-{�>�l�x���?'��U@��r�Cj�yY����	�垜=�C9??;�>�`�>ִ�?��?���]$���r�9-�@F�;�V�>��g?�:�>��>]L���� ���>��l?i}�>yݠ>���?X!�4�{�� ˽V��>��>��>!�o>��,�V/\��f��a����#9�#��=��h?�n��^�`�݅>�R?p��:mpJ<Q��>�v���!�����'�E>4y?B��=��;>lž��{�?+����'?u?R��&���M>�$?�?/
�>�E�?��`>79�����=�?qR?�D?C�D?��>�χ=��g�	���H�HoB=0��>´�>H^=���=U�꽙XU�W�.��`���;=�<�y��^��<,��G6/<��Q=x�>�ٿuVO��MҾcp���侑Y�U`�����E�B�)k��*w��j0��������N5ʽ/{�Ӥ������d�?��?�����˾��v������(N>iz��O>�����@u�0xR���ξ%1���F���;�->����L�'?�����ǿ򰡿�:ܾ2! ?�A ?1�y?��3�"���8�� >C�<�-����뾭����οH�����^?���>��/��w��>ޥ�>�X>�Hq>����螾1�<��?8�-?��>��r�-�ɿ`����¤<���?.�@�{A?��(����ƧU=P��>T�	?b�?>�.1�C�a���\�>+=�?���?��M=5�W�T\	�"�e?x<H�F�Hܻ��=7T�=��=���9�J>�b�>�E�4A�	Eܽ��4>�܅>R�"�@����^��<Ҵ]>z�ս���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=M��ƿ}�$�=}��Z=9�޺��[��罼���d�T��"���eo����؈h=���=�Q>+l�>�$W>�1Z>�fW?w�k?�N�>C�>�5佟��qξ&���H��e���������죾^S��߾�	������i�ɾ�'F����=��[�1����`"��+g��JT�L�
?&w>��Z��Y�%����ݾ[���K����d7�m�׾�;&��vy���? �S?�F��"WZ����|��I����7?��p�tԿ�i�D��k>�4=��$�|Nn>\J<�Ν���ԺW�Ri0?�7?�����n���@)>�c���`=w�+?��?xu@<٪>p%?��(������[>ü4>�^�>���>)�
>�⮾X�ڽ]?Y�T?2����̜���>Fٽ���z�_=�>��5��C㼝\>w��<V���2V�*��	�<�(W?[��>`�)���Ra�����f]==��x?ے?n-�>/{k?��B?�ޤ<�g��3�S�k��ew=��W?E*i?��>�����	о򀧾k�5?��e??�N>�bh�N��6�.�MU�F$?�n?#_?�z���v}�b��9���n6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�ٕ��Z�?z�?u���i@g<b���l�fn���~�<sͫ=)��G"������7���ƾ��
�/���w⿼ƥ�>DZ@W�1*�>9D8�^6�TϿ.���[о�Rq�f�?N��>�Ƚ����+�j��Pu�U�G��H����I�>�>Ty���͑�߽{��m;��k�����>�)	��و>J3S�ɵ�L��?<(�>\p�>Oj�>$���B������?IY��kο �������X?�]�?(~�?��?�16<8�v�J�z�1�XG?�gs?�GZ?�{ ��']��3�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?z!�>h�?a�=�_�>�Q�=���9-�b#>��=��>�*�?��M?FH�>]A�=��8��/��[F�!HR��$�q�C�<�>��a?�L?^Qb> ��'2��!��sͽMj1��l鼜R@��,�w�߽)5>��=>>M�D��Ӿ��?Gp�9�ؿj��0p'��54?!��>	�?��W�t�����;_?Hz�>�6��+���%���B�]��?�G�?=�?��׾�R̼�>;�>�I�>5�Խ����j�����7>8�B?=��D��x�o�k�>���?	�@�ծ?gi��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*&����J��%0�F3���9>A�>�;>\˚�v�=�jݼ��	>'�ȹ9�=�ץ>a�d>Ǭ�>J��>]�o>Fb>��~���!��}��&"��c<��)��!3��ng�FF��~݀�ܱ�~����9�����Y�+����4���R�������=��U?.R?�p?ċ ?	�x�7�>������=҅#��΄=1�>�l2?��L?��*?,��=�����d�<^���8��Vɇ�҇�>�]I>-~�>JR�>�'�>��9��I>/(?>݁�>&>��'=@�ݺ�z=��N>�U�>t��>2��>b+<>��>�˴�#1����h�Iw��:̽���?�����J�4-��.I�������ޞ=DU.?�K>����?п���.H?� ���%�ː+���>S�0?`dW?��>���U�� >F��&�j��k>Y����tl���)�9Q>j?.31>�D�>J5���,��^������F>�?�Ų�ܓ^�B��=�?����Dy=���>�Vҽ33��K����u�',:�{����7?�@1?[�X<�����5;�偘�8�\>�e�=0u�q>z�,>��ȼ%x>�`�,��V�=T�m>�>;b?ȣ+>S�=s0�>S����O��֩>K�C>�->�??�!%?��	�E���,����,��x>���>.�>��>��I��\�=>v�>��a>�)�p��*U��/>� �X>$/���`���u���y=ݛ�����=�Y�=',���<�2e&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾEh�>mx��Z�������u�0�#=E��>�8H?�V��#�O�d>��v
?�?�^�ߩ����ȿ2|v����>Q�?���?a�m��A���@����>7��?�gY?joi>�g۾:`Z����>ջ@?�R?�>�9�x�'���?�޶?ӯ�?��?>��?0�o?L�>�͘���/�o8���G��cV=��<���>��=`�ľ�I�!Г�X`��VSk������U>ȵ6=m�>��������.�=�Gh�7��YT�f��>;�n>�jF>�ؚ>��>���>5#�>�d=7;���(}�������K?���?-���2n��N�<Z��=)�^��&?�I4?"k[�}�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��F��<��K>*4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��NS��GB�>�e!?���>�Ү=B� ?��#?��j>W)�>�`E��9��q�E�H��>c��>H?��~?��?�Ϲ��X3�����桿��[�g<N>��x?@V?+ɕ>a������KmE�N%I�����?ug?�U��?=2�?A�??}�A?*f>�~��ؾ�������>&�!?��A�/N&�m
��~?�P?���>*6����ս�!ּ.��w}����?P(\?�@&? ���*a���¾�H�<.�"�fU��?�;߰D�#�>,�>�{�����=`
>@Ͱ=�Jm�jG6�
�f<Ii�=n��>��=�)7��n��/=,?��G�ۃ���=��r�?xD���>�IL>����^?il=��{�����x��	U� �? ��?Zk�?f��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>F�l���K���ڙ���F��_�Ž�W&��K�>O�>Kh?��>W�1>Ā�>������"�#���Q�,�Y�7z��[B�?(��=��@��n�M�c�|������c���:�>���<~D�>��>^>IYn>KN�>O�ܺ� �>��T>�3Z>Ť>��m>i9> �>���=�6JR?������'�´�˯��I3B?�rd?6�>��h�������d�?���?<r�?�Dv>yh��'+�o?�A�>���o
?5D:==��q�<9T��-��?)��z(����>R׽� :�JM��Xf��m
?O/?��}�̾E׽�-��`r=4�?P�'?��)�uR���o�	X��HR������m�����\(%�Wp�����NW��	���j�(���=f**?��?��ly�"u����j�t>��b>���>�H�>ma�>�PK>� 	��x1���\�n�'�K������>Y y?��>F?��<?��K?�>H?���>t��><��v\�>\Ƽ[��>T��>߉??,D,?��0?�"?et-?�~m>r'ƽID����վ?C?ک?Y�"?���>A\?�7���)޽Q)�[��8f��g����C�=p�n=��ý{���p��=41D>jZ?9����8������k>}�7?˂�>���>���,�����<��>��
?�I�>����zur��]��Z�>x��?7��!�=|�)>f��=�6��-�ֺ f�=+�����=�ā�1_;���<끿=��=�\t�IЂ�Ri�:�@�;"�<�t�>6�?���>�C�>�@��/� �c�� f�=�Y>>S>|>�Eپ�}���$��v�g��]y>�w�?�z�?̻f=��=��=}���U�����H������<�??J#?)XT?`��?{�=?_j#?ϵ>+�jM���^�������?��*?�Ր>p���-ƾ���d(3�P�?�=?S`���!�*��E¾G�ܽ�U>�t.��~�vۯ��1D����������xA�?`H�?<e�Cb7��羞��Fԭ��C?�H�>j�>���>��(��6f�H|�T<?>�R�>�?P?پ�>�O?$4{?&x[?qS>6�8�[����|���+h�� >��??���?8<�?� y?u7�>�j>�,���޾�T���Z�2���s��F=ZSY>:��>���>��>O��=;�ɽ�B���<;�:��=�<d>�k�>=�>,Z�>��v>��<&�G?W��>բ������n��7$;�y�u?���?�_+?7�=n%�{�E������y�>Ng�?���?y(*?"�R����=��ռ�����q�mͷ>��>y�>Қ�=�8K=
>���>���>�d�Sn�p8��J��?� F?3)�=��ÿ�g�K���q����Իi����
��ν��q��>�h�����S����a�\���D��((��T����u�����>E��=�h	>C��=�==0��I�<b�*=ʛL�	g�<mݣ��!=�2�Ւ1�D�Ƚy�%<G��<��=��"�)�˾��}?�;I?˕+?t�C?�y>$;>�3�J��>�����@?RV>G�P������;�Q���� ��a�ؾx׾��c�"ʟ��H>�_I�>�>�83>�G�=�K�<2�=�s=P=j�Q��=;$�=	P�=tg�=���=�>DU>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>.��=h5>*�\�!�;��_��,ݍ�V�����?ErA�v����>�=ʞ��QԾ:�	��-�=Y�
=)�/���a�j��=W� ���=�է=�>�>H->��=�+½��=޿;�%>vv>��<��7��h��=Rq�=P+4>��>���>�?�5?�??�֘>H3F�.������T�S>��]=��>�F>��>	��>N�>?D�9?#P??���>��>:��>[��>�O�$�o���������=���?��?���>�L�<)w����)�-�6�4˽�B/?L'V?Bb�>>��>�U����9Y&���.�$����{4��+=�mr��QU�M���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=$�����<�vż�����u&�:�+�1�����;r��;B�]<^��;��=���>�>3��>~p�=��� />�Ŗ�X�L����=�;��K&B��1d�vI~�_/��j6���B>f(X>�����/���?� Z>�u?>q��?,8u?��>e�]�վQ���4e��NS����=А>?=�s;��T`�(�M�[wҾ��>!��>ӡ>��o>�5,���>��t=o%㾴�4��_�>���x:���q�m¤��֟��;i��?����C?�؇����=�.~?��J?g&�?�F�>N♽
�׾�U->Q����9=�u�F�r��<����?!�%?�J�>$�ӤD�CҾLª�7�>x`�
CP�����$�3��.��q���4�>�����EӾ�f3������6��DLE��`u�v��>E?)�?^9I�~����gN�.�����y?M%a?��>/?��?xJ�N��∾I��=�i?n�?yz�?L�=R��=3���<�>{�?�@�?�]�?��s?h4��o�>?����>6���X��=�>~�=E]�=�K?`.?��?����E	����	��L����<"��=��> �>Z�x>�U�=�aX=߾�=+nf>j�>�b�>CEb>q��>+~�>�Z��Hi���&?�g�=vt�>u2?a`�>��W=������<��K�h+?�f+��Ҹ�n����<ڰ��\&O=��ͼ�$�>o�ǿe.�?�T>�o�:�?g"����/�'�S>(�T>��޽���>JhE>�G}>S��>�&�>��>3��>�(>c5׾О>@��� $�ÄC��IS��q׾ �j>N����c�	�(���(P�}��*)�7ok�
N����:�Ú�;_�?��޽�k�Ʋ)�[��:??>7�>�d2?�U��@Uk��C&>r��>_�>�Z������{��^�־ˍ�?��?}5c>��>p�W?��?1��3�,tZ�̯u��&A��	e���`�B���՜����
�R����_?��x?ZtA?��<�7z>[��?��%�ŏ��3�>p /��%;��<<=�#�>�%��5�`�.�ӾW�þt4��KF>�o?,%�?\?YV�E�i���&>��:?�j1?�t?�2?u�;?K��vE%?'�2>d�?�?�l5?W�.?5�
?��3> �=��x�/�,=�t��{���p�ѽ��ǽ��ֲ5=��}=Շu9(D<w=�$�<_�\ؼ;8q��]/�<�	;=3ף=C'�=�Ȧ>d�]?�p�>w}�>V�7?�t�9?8��b��J5/?$7=����Ί��T�����>�j?a��?�[Z?��d>!�A���B�|�>�|�>�/'>[�[><g�>�ͽE�۷�=��>s�>��=�K�������	�f�����<u�>�F�>=�{>/$��h�)>�ޣ��lz��c>�eS����=�U��SH�&�1��vw����>˜K?�R?A�=���[���e���(?��<?��M?��?.�=S�۾��9���J��g�ʃ�>��<2	�s|��|ѡ���:���.;U�u>�l���*��uef>�J
�߾��m�"�I��v边G=�^�5�P=�
�
Ծkm��v�=�w>�����f��e������5aI?Q�c=d<��S�4���U>퇛>���>J�b�l���?9>��q����=H��>�D>��N��z�F��a����> �M?��A?`�[?��9�{���,@��{��e��i�=>Y�>��>���>�RA�/��y�޾���V�f��C��c�>S��>�ɾ�[���������7�͸?]{�>6��=�G?��(?���>'d�?iIa?'�>7 �>^Z��.�NA&?���?��=�Խ2�T�? 9��F�?��>"|)?�B�(��>Ҋ?��?��&?��Q?��?��>w� �)F@�#��>�V�>��W��_��w�_>�J?��>�;Y?�у?��=> �5�!袾nݩ�]l�=-!>b�2?�3#?Z�?�>���>���>�?cU�?d�,?�$t?��>w�>�ʽ�d?��>+�}>�L?��J?�R?%�?nVL?ehQ>��
>�Q�v=�SA=Ѥ�����ǘQ=/��>��=�޽����G��٭r</O�����K=a)�J2���N���s�>(�u>���.>;�ľD<���+?>r����E��&���_6;���=��>�?W��>�%�ݑ=���>>��>xt�$�'?�?��?���;%}b�.۾��K�@Y�>�B?X��=Pkl�m{��o/v��Ui=��m?UT^?)X��w��h�b?� ^?�a=���þ�jc����z�O?ٍ
?ZFG��>��~?n�q?�W�>ϥe�/&n�	✿�pb���k��Z�=�4�>$�H�d�=J�>7?�V�>ɢc>ݫ�=��۾�@w�Mo����?*�?v�?X��?�8*>4�n�['࿖��A@���gc?z�>�,���%?��<��i��||�;����h������i��(���e��<������=��?�h?�9t?Tf^?�*��ݽb�G`d��\{�;�[��
�����@��<��@���p�������<R��%'n=u���S����?��)?)�~����>h|���7�� <��ĵd>����#�r\}�ͅ�����<�Q�=X�����Z�J˥���$?*�>B��>�9?��N��v?�+BG��C.�����fW=�l�>��>)1�>�1�x�H۽:����"������x��>~!a?,5;?P>?�O���/�:t�����c�]��J
_>��>�S>4�Kw��[��ޕ�v˂� E+��@a�y� �ޱB=i�)?��w=���>���?+��>:�*�p׾U~���{�=K�>&l?8?Zm>#Y޼h�2�Nq�>�o?ib>�E>���F� ��Ox��:�����>��"?	P>����ie���{�jʇ�Xŉ�1�;����>U�u?����@��ru�>0>�?�#`=x���sM?�ɑ�)�'���ҾL�\��>g��>3�T=9�\&F��$�����}�UP)?�H?���*�w4~>�$"?o�>#.�>/�?2*�>�Xþ��|�Ӵ?��^?�:J?�GA?�N�>��=�Ա��Ƚg�&���,=��>�Z>5�l=�a�=в�=e\� F��BD=$j�=$ϼ5����<iJ���J<1l�<?�3>�-ܿE<=�չ���>���r���7�P���:��j�LT�[��.�����������6m�oC��&p�)ȅ��w�1<�?��?\����ɑ��;����w��y�Q/�>��� 20��$������Gl����¾���K��h��Zb�xU'?f^���ǿ������޾)"??�?ۆw?;����!�tO8���>���<X�ȼ��:����ο�M��[`?���>
��0ˮ�e��>9Ԁ>�Kb>0q>�0�������(<:�?b�(?<,�>��h���ǿv����Ax<C��?/�@TxA?�(�	���*V=���>S}	?��?>B�1�7\�9��|M�>�8�?��?�iM=ĳW�b�	�Ewe?\��;�G��޻��=mK�=�=����J>�h�>���XA��_ܽ��4>~�>f�!�#���J^���<H�]>mս�x��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=��^�ƿϰ$�F��O=]R���W��$�Aԩ�ыV���Hp�rH콙<i=�[�=9xQ>��>��V>\�Y>G~W?��k?A�>�>ē�&����;���h�����h���q�T�������B|	�������iʾ'=�&��=�R�����Ѯ �E�b�ktF�e�.?�j$>��ʾ��M��P(<?�ʾ����ڧ����^̾Г1� n�]Ɵ?��A?�݅�u�V�AD��4��`����W?r�L��S���Ҁ�=����R�=�>�=#��M*3���S��j0?�k?$>���z��7#)>g� ���=m+? ?�XQ<�?�>E%?D�*��_�>�[>�&3>$ۣ>�C�>��>Ԯ��P۽�q?ڄT?���0윾�#�>4q���{���b=4�>��4�C�� �Z>ݦ�<xa��R�Y��׎��3�<��V??�>+B*��s��7��8�_S5=�&x??O?T�>v�j?Y�B?��<����4T����W�l=3W?�{i?v�>�W����оHƧ��5?�Jf?ErO>�i��D�./�����?��n?{?j���o}����L#���6?��v?0r^�rs��=����V�X>�>�Z�>@��>�9��l�>�>?O#�FG���]Y4��?S�@���?��;<b����=�;?�\�>i�O�_?ƾ|��������q=m#�>����0ev�����T,�$�8?Ӡ�?C��>2������K��=w�ܾ��?p�?�aپ�p��#�(���-������ҽy�=��W���@�5���E>��H��A�(����?�+p�>H�@�:�XL�>|/P��g꿎�ؿ������
����$?���>�=��̾�ǆ�k6��9�D���H�nP��^�>�Z>NE�������{���;�ُ��s��>���$�>�S���ӝ���
0<P͒>�N�>��>Q갽I����?*D���ο����,��4�X?�M�?�x�?:?�1<��u���{�v��HtG?��s?�Z?�M$���]�_;��h?�s�G?d��G�x�B�X~�>,4?I��>����@>��>[Ϝ>�:>�6�g]�������]񾼘�?���?�Ҿ��>u*�?�f.?2m�?�������%���	�I?⺾=q��� 5$�+�L��r���?��&?v3�42�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�8�>P�?��=3�>l3�=�����,���">5��=T�@���?əM?�#�>�B�=!{8�@/��8F�RR�]J��C����>��a?��L?��a>C︽�h.�B!�Zuν��1��w�)�?���)��^߽��5>nc>>�>�3D��+Ӿ/?r&���ֿ�2��Z���7v?GM�:-�>�u �>T3�_�X=p��>n��>�5
�����S��!s��L�?��?���>�y��т�=�ay=��>��> 	 ���%͛�+��>5�2?�ǂ��<W��+c�	>�>Z4�?h@��?��d��	?���P��fa~���87����=��7?t0�T�z>���>��=�nv�ۻ��P�s����>�B�?�{�?,��>�l?��o�7�B���1=9M�>��k?�s?CQo��󾵲B>|�?!������L��f?�
@{u@U�^?%�������� ��g;�X>�54=¬]> �f�_�)� {�����=�����)9>MY�>8æ>*7�>�f>&�U>�6>�����7��?����:�7 ���	�p�����*Z�����R���^��b���U&߼�>�2h���^<����<њ7>�N??�4?	�M?/~>ju;��o�>�s�u4��ԾX>�	?\�S? G-?�1?�=d>�%��O��	�������k_�H��>�n>�l?a�>���>�V�=�"�>פ�=w��>-�1>��'=���=�Y����>a��>J��>S�>�C<>ݑ>8ϴ��1��h�h��
w��̽#�?����L�J��1���9��Ҧ���h�=Ab.?�{>���?пd����2H?%���t)�ȹ+�?�>|�0?�cW?�>L����T�F:>+��{�j�a`>G+ �6l���)��%Q>\l?�Jg>o�u>7P3��?8���P�����
|>�5?�߷�':��Tu�xYH�>ݾ�M>���>�uG��(�����ZD��i�b�y=[-:?+�?봽����C8s�����ӫP>nH[>��=�)�=ʞN>_�b�p�ýwF�?�.=7�=�A]>#]?�]->�ٌ=���>�\��ȅN�O��>ӉA>��,>_@?�%?)B�P��7����-� �u>m�>؁>/�>ڱI����=���>{�b>}>��������?��V>��t�;N`��v�G�r=wD���?�=�p�="� ���<���%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿv3�>/|w<@���y��-����>tk>o�?�߾�N<��������>k/�>��
����!�ѿ.����D�>z�?��?�8��ɗ��+7����>�?ygD?�=n{���9��[��>��>}�X?��>�;2`��,�>�0�? ��?{D>X?�?ld`?�l�>8�;�42�����g��_k8=� =�&#>�<>������S�M������6Lc���v�Z>F�U==G�>�AP�]Wվ��=�!��XkǾd�^��8�>FiS>�Ɵ>�>]�>C �>p;�>i����<S���,)о�K?��?6����m��L�<6��=3X^�4�?�V3?��n�d0Ͼiި>�_\?��?��Z?y�>��:���￿W9�����<�9K>ɍ�>�y�>��sM>pQվ�lE�m�>س�>�B��پ3聾%�a�xԝ>�;!?��>�=��?�$?�b>�[�>�D��L����J��T�>�b�>�a?��s?�?`����5��ה��硿ç\���6>��w?X�?;F�>����ˣ����ߘ���@��l|??�a?|Ͻ�?�`�?P�??��=?�ra>WJ?�.׾�{��W��>#�!?�&��tA�D3&�V���1?v(?LA�>�"���w׽�tҼ'��`R����?�\? &?�g��Aa���þr�<`'��9b�[�<��Q�p�>A=>�]��n�=bB>��=Gl���4���i<�ž=��>��=5�5� Q��6=,?��G��ۃ�>�=��r�xD���>�IL>���Ŭ^?~l=�8�{�����x��B	U�� �?��?ck�?K��$�h��$=?�?w	?5"�>FK���}޾O���Pw��}x��w���>���>�l���.���ڙ���F��C�ŽW����>��>�?�?�a0>��>z@���.$�A�޾��V�U��Z��j>�W2��������,��P|����&e��7�>������>ʝ?A'U>��i>@�>�H�����>��Y>A\>'B�>/IY>+s >��'>�FW���$�,IR?B�����'����l°��@B?6_d?��>3�h����$��Pj??7l�?bv>��h�h6+�qq?�U�>���Wq
?$a:=��້<�O��Ĺ��9��`�����>� ׽�$:�HM��Gf�o
?+/?�-��!W̾WR׽e}���+=◅?��$?��'�>Lt�]l��˃3�>�5��k�E&��Mq-�)�.�|?t��W��T�r�m���-�@�\�e=B�'?=X�?�W6�����]z��r`�8�Pa�<]�? ��>ep>/�>G�оYC���p��b� L�&��>� y?��>ۖ??7??{>J?�<?pu<>���>����X��>#����R�>�
?s?F/?��2?��?��.?>>�퉾�	�4���j?��?>�.?�_�>���>�@���=��*>B�O=kB��D����	��2d	��)��S��S�=�>�w?���
9�>���@h>�68?r��>��>������}�D�<���>��
?X�>������r������>籂?%���~1=�,>8�= ��������=�yȼx��=�MA��2H��<�_�=ۉ=��Y�,^;�;9l;���<,u�>[�?(��>�B�>�@��ϩ �����d�=}Y>�S>>�Fپ�}���$��_�g��\y>�w�?�z�?��f=��=0��=y|���T������������<��?�I#?#XT?��?��=?j#?��>+�2M���^��$����?�!,?��>7��F�ʾ+��3���?pY?z9a���4;)���¾��Խ��>�[/��/~����D�K���������p��?$��?�A�f�6�Iv�����\��B�C?�>�Z�>��>��)���g�5#�y*;>V��>�
R?�Q�>`QO?��x?��Y?MG>n8�׏��c��%0	�X�>�P???�Q�?I�v?���>X>�#��0⾿G ��2&��p���ǀ�n?x=n:Z>惑>.o�>�>��=/�˽&��,#2�ö�=z�d>`c�>�Ū>��>��}>l��<��G?���>�e�����&菉����z=���u?;��?��+?�g=#��@�E��N���A�>Lh�?��?�;*?>�S����=S�ּ7Զ�.�q��#�>�˹>�)�>���=�?F=R}>)��>Ԛ�>�8�3h�zm8�EM���?\F?m��=hƿ��q���p��җ��d<Q풾=�d�t����Z��_�=�����M�����[�ǡ��r|������2���w�{���>��=E��=���=C��<��ɼm�<�*L=�n�<h�=hp�"'n<.69�hy˻N(��>��C�Z<h�H=�`���ƾ"Wy?��K?�,?�jE?��d>�(>�D�(�>�NH�5^?:�[>���5W��T"(��Ꜿ�X���2Ҿ�۾Ɏd�d���>�F`��>�72>��=z8=n>p�=s�^=er��h0�<�j�=x=�h�=|A�=.>�43>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��=>��>�[O�+�/�
g��g���U�H�?9F?�v�Ͼ!P�>���=a2ܾ��þ��S=�93>f�m=l�#��_�L'�=�����D3=�m�=� �>_B>
��=if½�D�=h3=|�==X>�I<�;0�
N�I�k=m��=��m>A`>�Q�>F�?�Y0?8+d?߹>�Qn���;�����>���=C��>�[�=��B>��>V�7?��D?@�K?�ڱ>R��=��>p��>�
,��7m�'#�`������<Y��?�Ն?&I�>=�c<ӝB��h��r>��Ľ�?�0?RJ?i�>jv�	�9!>�%�6����;���<��=�������je�^u��KԽZ�#>���>���>���>�	O>��>�Ee>3��>�*>_C�=�#M=��Y==�=�*��z���!�<N��=�q.<^kr=+P�����)ƨ�5�߼q��t���<.��=���>��>���>}�=�����1>#B��ˬK���=���@�t.b���~��/���8�c<>�bU>�bt�Ա��	:?:�Z>�@>��?:�s?�I">p��Kg־W�΁a�CXM�';�=.;>��<� �:���]�^�N�7	־��>̉�>�0p>���>2��C�I��=s6���$�{�>^r��X�o�M)���{�8��� �;j�0����%G?B��ߙ�=+
o?,3A?Pd�?Y�>�fW��&�=&і�;p=+�侁����ӽ,�
?ޮ?
�?`l	���W��C̾�����ڷ>*<I�(�O�-�&�0�����ȷ����>������о�"3�^h�������B�Rr���>��O?��?�(b��U���WO�����$���k?:|g?*�>NJ?�D?�&���y�k��=��=��n?��?m:�?��
>�Խ=�t��sT�>�7	?���?K��?z�s?��>�^�>�s;�O!>7���Fv�=��><��=�>�=߈?ו
?��
?X	��X�	����񾂴]�A�<�'�=|
�>��>�r>��=�f=�n�=;�[>q��>��>2=e>���>KM�>��۾��%-?���=	��=�)?�D�>Ya�>|I>�<>��
�3h�U���^��@����=e숽pE��u��5	?�Aҿ)��?���>v���?l���wϽ�MF>�(�>E�]����>���=��=1�>���>T�ú��>�i>�߮�c]O>����)��iB��RV��	�i�Q>70�Ef<����;�4l���޾V�'�]�t��n���[C��0�=<��?[Ǘ��@���aK�\�P�߅=?d��>j�?zG��lO"����=���>0{�>l�߾�䅿������?���?�;c>�>��W?�?o�1�I3��uZ���u�:(A��e���`�H፿霁�V�
��	����_?��x?�xA?�Q�<M:z>H��?r�%�ԏ�g)�>�/�k';��E<=U+�>*����`�2�Ӿ��þ�6�6JF>�o?O%�?Y?�VV�E3s���>
�H?h@.?�u?D�
?lL??�>��d^?�x-> �?�?}�?l�.?sP?<r>�WW>�I=DM�@a���땾$ᱽ����[�q�xe}=��=g�>ė=���_�P�������f�=k=��:{}<���=��=�c>궦>ĝ]?�U�>	��>�7?���MV8����
/?�9="g��1ꊾ����t��->4�j?���?hKZ?��c>��A�V�B��\>�]�>:�&>��[>�D�>�=�	&E��=dE>�>��=�:N�Oց���	�O����&�<��>���>�=|>J���b�'>�i���Kz�3�d>h!R��Ӻ�M�S���G���1�dv��<�>��K?��?o��=_龹V��\>f��))?�[<?NDM?]�?C��=`�۾9�9�K�J���*�>�ܩ<|	���� ����:���:��s>53��Χ׾*R�>���}�$��j�L�^��y�5~��e(���E>[Ǿ!���ž/���ġ�d����8Ԟ�:��-
-?-&�=kk�d���ž�q>��>�֬>�=Q>����M�����<�?9>(��>�����^�D��u����H>0:?�iU?m�?�u���I��(�Ǿ�����Z߻�@?�b�>�?��q>�I>����<�&�N�,���>��R�>u�>ㅰ��gS�Lݙ�d���g�⾡��>��?��=�%?�W?8�I?%��?�L,?q)?��>�'�g��`]$?�À?0q�=�?ƽ&~R��U7�iU?�}C�>��?��G���>8�?7�$?��)?xCR?��?ʃ�=���7��l�>K
�>��N��`��[Y>ڡU?���>�`?炅?�/>|�.��A���n�����=��>��;?��-?�	?�~�>K	?�Ԟ�k�<�Y�>]Ma?p�?�2}?���><$*?t<U��k�>���>�x�><�?�1+?�U?su?��V?��$?�	�=����_�H�ˉ=�>��=�3��Gƅ�+ҽ�i��C�=iU���+��6�ZD���$'�{��a�e=IA= R�>��s>����1>��ľOJ����@>+{��<I��V�{�:����=�s�>h�?«�>�f#�w|�=֖�>^:�>����)(?}�?S ?��3;��b�A�ھĉK���>� B?N��=?�l� �����u��h=9�m?#�^?@GW����O�b?��]??h��=��þ{�b����g�O?=�
?4�G���>��~?f�q?U��>�e�+:n�*��Db���j�'Ѷ=\r�>LX�S�d��?�>o�7?�N�>1�b>)%�=iu۾�w��q��h?��?�?���?+*>��n�Y4࿹���`����i?`�>�lk���?�=�6E���1a�A��m�ƾ$n�����'EV�\1�����p����[5�N�=���>-S?5?Hb.?���ܥ��ֶ������Y8�ݶ��=�V�*/F��s)��0n�(�3��"�Gz����.Y���A���?��'?�0�Ù�> ͘����;��B>𤟾2!���=8\����?=�Z=W�h�D�.��X��l ?�&�>P6�>��<?��[�cF>���1�8�7�������3>�բ>���>w;�>���:�>-���Q�ɾ���Խ��m>�T`?,F?vn?,b�Y�/�B瀿��#�u�6�Nԯ��!>I�>-{�>�l�x���?'��U@��r�Cj�yY����	�垜=�C9??;�>�`�>ִ�?��?���]$���r�9-�@F�;�V�>��g?�:�>��>]L���� ���>��l?i}�>yݠ>���?X!�4�{�� ˽V��>��>��>!�o>��,�V/\��f��a����#9�#��=��h?�n��^�`�݅>�R?p��:mpJ<Q��>�v���!�����'�E>4y?B��=��;>lž��{�?+����'?u?R��&���M>�$?�?/
�>�E�?��`>79�����=�?qR?�D?C�D?��>�χ=��g�	���H�HoB=0��>´�>H^=���=U�꽙XU�W�.��`���;=�<�y��^��<,��G6/<��Q=x�>�ٿuVO��MҾcp���侑Y�U`�����E�B�)k��*w��j0��������N5ʽ/{�Ӥ������d�?��?�����˾��v������(N>iz��O>�����@u�0xR���ξ%1���F���;�->����L�'?�����ǿ򰡿�:ܾ2! ?�A ?1�y?��3�"���8�� >C�<�-����뾭����οH�����^?���>��/��w��>ޥ�>�X>�Hq>����螾1�<��?8�-?��>��r�-�ɿ`����¤<���?.�@�{A?��(����ƧU=P��>T�	?b�?>�.1�C�a���\�>+=�?���?��M=5�W�T\	�"�e?x<H�F�Hܻ��=7T�=��=���9�J>�b�>�E�4A�	Eܽ��4>�܅>R�"�@����^��<Ҵ]>z�ս���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=M��ƿ}�$�=}��Z=9�޺��[��罼���d�T��"���eo����؈h=���=�Q>+l�>�$W>�1Z>�fW?w�k?�N�>C�>�5佟��qξ&���H��e���������죾^S��߾�	������i�ɾ�'F����=��[�1����`"��+g��JT�L�
?&w>��Z��Y�%����ݾ[���K����d7�m�׾�;&��vy���? �S?�F��"WZ����|��I����7?��p�tԿ�i�D��k>�4=��$�|Nn>\J<�Ν���ԺW�Ri0?�7?�����n���@)>�c���`=w�+?��?xu@<٪>p%?��(������[>ü4>�^�>���>)�
>�⮾X�ڽ]?Y�T?2����̜���>Fٽ���z�_=�>��5��C㼝\>w��<V���2V�*��	�<�(W?[��>`�)���Ra�����f]==��x?ے?n-�>/{k?��B?�ޤ<�g��3�S�k��ew=��W?E*i?��>�����	о򀧾k�5?��e??�N>�bh�N��6�.�MU�F$?�n?#_?�z���v}�b��9���n6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�ٕ��Z�?z�?u���i@g<b���l�fn���~�<sͫ=)��G"������7���ƾ��
�/���w⿼ƥ�>DZ@W�1*�>9D8�^6�TϿ.���[о�Rq�f�?N��>�Ƚ����+�j��Pu�U�G��H����I�>�>Ty���͑�߽{��m;��k�����>�)	��و>J3S�ɵ�L��?<(�>\p�>Oj�>$���B������?IY��kο �������X?�]�?(~�?��?�16<8�v�J�z�1�XG?�gs?�GZ?�{ ��']��3�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?z!�>h�?a�=�_�>�Q�=���9-�b#>��=��>�*�?��M?FH�>]A�=��8��/��[F�!HR��$�q�C�<�>��a?�L?^Qb> ��'2��!��sͽMj1��l鼜R@��,�w�߽)5>��=>>M�D��Ӿ��?Gp�9�ؿj��0p'��54?!��>	�?��W�t�����;_?Hz�>�6��+���%���B�]��?�G�?=�?��׾�R̼�>;�>�I�>5�Խ����j�����7>8�B?=��D��x�o�k�>���?	�@�ծ?gi��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*&����J��%0�F3���9>A�>�;>\˚�v�=�jݼ��	>'�ȹ9�=�ץ>a�d>Ǭ�>J��>]�o>Fb>��~���!��}��&"��c<��)��!3��ng�FF��~݀�ܱ�~����9�����Y�+����4���R�������=��U?.R?�p?ċ ?	�x�7�>������=҅#��΄=1�>�l2?��L?��*?,��=�����d�<^���8��Vɇ�҇�>�]I>-~�>JR�>�'�>��9��I>/(?>݁�>&>��'=@�ݺ�z=��N>�U�>t��>2��>b+<>��>�˴�#1����h�Iw��:̽���?�����J�4-��.I�������ޞ=DU.?�K>����?п���.H?� ���%�ː+���>S�0?`dW?��>���U�� >F��&�j��k>Y����tl���)�9Q>j?.31>�D�>J5���,��^������F>�?�Ų�ܓ^�B��=�?����Dy=���>�Vҽ33��K����u�',:�{����7?�@1?[�X<�����5;�偘�8�\>�e�=0u�q>z�,>��ȼ%x>�`�,��V�=T�m>�>;b?ȣ+>S�=s0�>S����O��֩>K�C>�->�??�!%?��	�E���,����,��x>���>.�>��>��I��\�=>v�>��a>�)�p��*U��/>� �X>$/���`���u���y=ݛ�����=�Y�=',���<�2e&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾEh�>mx��Z�������u�0�#=E��>�8H?�V��#�O�d>��v
?�?�^�ߩ����ȿ2|v����>Q�?���?a�m��A���@����>7��?�gY?joi>�g۾:`Z����>ջ@?�R?�>�9�x�'���?�޶?ӯ�?��?>��?0�o?L�>�͘���/�o8���G��cV=��<���>��=`�ľ�I�!Г�X`��VSk������U>ȵ6=m�>��������.�=�Gh�7��YT�f��>;�n>�jF>�ؚ>��>���>5#�>�d=7;���(}�������K?���?-���2n��N�<Z��=)�^��&?�I4?"k[�}�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��F��<��K>*4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��NS��GB�>�e!?���>�Ү=B� ?��#?��j>W)�>�`E��9��q�E�H��>c��>H?��~?��?�Ϲ��X3�����桿��[�g<N>��x?@V?+ɕ>a������KmE�N%I�����?ug?�U��?=2�?A�??}�A?*f>�~��ؾ�������>&�!?��A�/N&�m
��~?�P?���>*6����ս�!ּ.��w}����?P(\?�@&? ���*a���¾�H�<.�"�fU��?�;߰D�#�>,�>�{�����=`
>@Ͱ=�Jm�jG6�
�f<Ii�=n��>��=�)7��n��/=,?��G�ۃ���=��r�?xD���>�IL>����^?il=��{�����x��	U� �? ��?Zk�?f��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>F�l���K���ڙ���F��_�Ž�W&��K�>O�>Kh?��>W�1>Ā�>������"�#���Q�,�Y�7z��[B�?(��=��@��n�M�c�|������c���:�>���<~D�>��>^>IYn>KN�>O�ܺ� �>��T>�3Z>Ť>��m>i9> �>���=�6JR?������'�´�˯��I3B?�rd?6�>��h�������d�?���?<r�?�Dv>yh��'+�o?�A�>���o
?5D:==��q�<9T��-��?)��z(����>R׽� :�JM��Xf��m
?O/?��}�̾E׽�-��`r=4�?P�'?��)�uR���o�	X��HR������m�����\(%�Wp�����NW��	���j�(���=f**?��?��ly�"u����j�t>��b>���>�H�>ma�>�PK>� 	��x1���\�n�'�K������>Y y?��>F?��<?��K?�>H?���>t��><��v\�>\Ƽ[��>T��>߉??,D,?��0?�"?et-?�~m>r'ƽID����վ?C?ک?Y�"?���>A\?�7���)޽Q)�[��8f��g����C�=p�n=��ý{���p��=41D>jZ?9����8������k>}�7?˂�>���>���,�����<��>��
?�I�>����zur��]��Z�>x��?7��!�=|�)>f��=�6��-�ֺ f�=+�����=�ā�1_;���<끿=��=�\t�IЂ�Ri�:�@�;"�<�t�>6�?���>�C�>�@��/� �c�� f�=�Y>>S>|>�Eپ�}���$��v�g��]y>�w�?�z�?̻f=��=��=}���U�����H������<�??J#?)XT?`��?{�=?_j#?ϵ>+�jM���^�������?��*?�Ր>p���-ƾ���d(3�P�?�=?S`���!�*��E¾G�ܽ�U>�t.��~�vۯ��1D����������xA�?`H�?<e�Cb7��羞��Fԭ��C?�H�>j�>���>��(��6f�H|�T<?>�R�>�?P?پ�>�O?$4{?&x[?qS>6�8�[����|���+h�� >��??���?8<�?� y?u7�>�j>�,���޾�T���Z�2���s��F=ZSY>:��>���>��>O��=;�ɽ�B���<;�:��=�<d>�k�>=�>,Z�>��v>��<&�G?W��>բ������n��7$;�y�u?���?�_+?7�=n%�{�E������y�>Ng�?���?y(*?"�R����=��ռ�����q�mͷ>��>y�>Қ�=�8K=
>���>���>�d�Sn�p8��J��?� F?3)�=��ÿ�g�K���q����Իi����
��ν��q��>�h�����S����a�\���D��((��T����u�����>E��=�h	>C��=�==0��I�<b�*=ʛL�	g�<mݣ��!=�2�Ւ1�D�Ƚy�%<G��<��=��"�)�˾��}?�;I?˕+?t�C?�y>$;>�3�J��>�����@?RV>G�P������;�Q���� ��a�ؾx׾��c�"ʟ��H>�_I�>�>�83>�G�=�K�<2�=�s=P=j�Q��=;$�=	P�=tg�=���=�>DU>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>.��=h5>*�\�!�;��_��,ݍ�V�����?ErA�v����>�=ʞ��QԾ:�	��-�=Y�
=)�/���a�j��=W� ���=�է=�>�>H->��=�+½��=޿;�%>vv>��<��7��h��=Rq�=P+4>��>���>�?�5?�??�֘>H3F�.������T�S>��]=��>�F>��>	��>N�>?D�9?#P??���>��>:��>[��>�O�$�o���������=���?��?���>�L�<)w����)�-�6�4˽�B/?L'V?Bb�>>��>�U����9Y&���.�$����{4��+=�mr��QU�M���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=$�����<�vż�����u&�:�+�1�����;r��;B�]<^��;��=���>�>3��>~p�=��� />�Ŗ�X�L����=�;��K&B��1d�vI~�_/��j6���B>f(X>�����/���?� Z>�u?>q��?,8u?��>e�]�վQ���4e��NS����=А>?=�s;��T`�(�M�[wҾ��>!��>ӡ>��o>�5,���>��t=o%㾴�4��_�>���x:���q�m¤��֟��;i��?����C?�؇����=�.~?��J?g&�?�F�>N♽
�׾�U->Q����9=�u�F�r��<����?!�%?�J�>$�ӤD�CҾLª�7�>x`�
CP�����$�3��.��q���4�>�����EӾ�f3������6��DLE��`u�v��>E?)�?^9I�~����gN�.�����y?M%a?��>/?��?xJ�N��∾I��=�i?n�?yz�?L�=R��=3���<�>{�?�@�?�]�?��s?h4��o�>?����>6���X��=�>~�=E]�=�K?`.?��?����E	����	��L����<"��=��> �>Z�x>�U�=�aX=߾�=+nf>j�>�b�>CEb>q��>+~�>�Z��Hi���&?�g�=vt�>u2?a`�>��W=������<��K�h+?�f+��Ҹ�n����<ڰ��\&O=��ͼ�$�>o�ǿe.�?�T>�o�:�?g"����/�'�S>(�T>��޽���>JhE>�G}>S��>�&�>��>3��>�(>c5׾О>@��� $�ÄC��IS��q׾ �j>N����c�	�(���(P�}��*)�7ok�
N����:�Ú�;_�?��޽�k�Ʋ)�[��:??>7�>�d2?�U��@Uk��C&>r��>_�>�Z������{��^�־ˍ�?��?}5c>��>p�W?��?1��3�,tZ�̯u��&A��	e���`�B���՜����
�R����_?��x?ZtA?��<�7z>[��?��%�ŏ��3�>p /��%;��<<=�#�>�%��5�`�.�ӾW�þt4��KF>�o?,%�?\?YV�E�i���&>��:?�j1?�t?�2?u�;?K��vE%?'�2>d�?�?�l5?W�.?5�
?��3> �=��x�/�,=�t��{���p�ѽ��ǽ��ֲ5=��}=Շu9(D<w=�$�<_�\ؼ;8q��]/�<�	;=3ף=C'�=�Ȧ>d�]?�p�>w}�>V�7?�t�9?8��b��J5/?$7=����Ί��T�����>�j?a��?�[Z?��d>!�A���B�|�>�|�>�/'>[�[><g�>�ͽE�۷�=��>s�>��=�K�������	�f�����<u�>�F�>=�{>/$��h�)>�ޣ��lz��c>�eS����=�U��SH�&�1��vw����>˜K?�R?A�=���[���e���(?��<?��M?��?.�=S�۾��9���J��g�ʃ�>��<2	�s|��|ѡ���:���.;U�u>�l���*��uef>�J
�߾��m�"�I��v边G=�^�5�P=�
�
Ծkm��v�=�w>�����f��e������5aI?Q�c=d<��S�4���U>퇛>���>J�b�l���?9>��q����=H��>�D>��N��z�F��a����> �M?��A?`�[?��9�{���,@��{��e��i�=>Y�>��>���>�RA�/��y�޾���V�f��C��c�>S��>�ɾ�[���������7�͸?]{�>6��=�G?��(?���>'d�?iIa?'�>7 �>^Z��.�NA&?���?��=�Խ2�T�? 9��F�?��>"|)?�B�(��>Ҋ?��?��&?��Q?��?��>w� �)F@�#��>�V�>��W��_��w�_>�J?��>�;Y?�у?��=> �5�!袾nݩ�]l�=-!>b�2?�3#?Z�?�>���>���>�?cU�?d�,?�$t?��>w�>�ʽ�d?��>+�}>�L?��J?�R?%�?nVL?ehQ>��
>�Q�v=�SA=Ѥ�����ǘQ=/��>��=�޽����G��٭r</O�����K=a)�J2���N���s�>(�u>���.>;�ľD<���+?>r����E��&���_6;���=��>�?W��>�%�ݑ=���>>��>xt�$�'?�?��?���;%}b�.۾��K�@Y�>�B?X��=Pkl�m{��o/v��Ui=��m?UT^?)X��w��h�b?� ^?�a=���þ�jc����z�O?ٍ
?ZFG��>��~?n�q?�W�>ϥe�/&n�	✿�pb���k��Z�=�4�>$�H�d�=J�>7?�V�>ɢc>ݫ�=��۾�@w�Mo����?*�?v�?X��?�8*>4�n�['࿖��A@���gc?z�>�,���%?��<��i��||�;����h������i��(���e��<������=��?�h?�9t?Tf^?�*��ݽb�G`d��\{�;�[��
�����@��<��@���p�������<R��%'n=u���S����?��)?)�~����>h|���7�� <��ĵd>����#�r\}�ͅ�����<�Q�=X�����Z�J˥���$?*�>B��>�9?��N��v?�+BG��C.�����fW=�l�>��>)1�>�1�x�H۽:����"������x��>~!a?,5;?P>?�O���/�:t�����c�]��J
_>��>�S>4�Kw��[��ޕ�v˂� E+��@a�y� �ޱB=i�)?��w=���>���?+��>:�*�p׾U~���{�=K�>&l?8?Zm>#Y޼h�2�Nq�>�o?ib>�E>���F� ��Ox��:�����>��"?	P>����ie���{�jʇ�Xŉ�1�;����>U�u?����@��ru�>0>�?�#`=x���sM?�ɑ�)�'���ҾL�\��>g��>3�T=9�\&F��$�����}�UP)?�H?���*�w4~>�$"?o�>#.�>/�?2*�>�Xþ��|�Ӵ?��^?�:J?�GA?�N�>��=�Ա��Ƚg�&���,=��>�Z>5�l=�a�=в�=e\� F��BD=$j�=$ϼ5����<iJ���J<1l�<?�3>�-ܿE<=�չ���>���r���7�P���:��j�LT�[��.�����������6m�oC��&p�)ȅ��w�1<�?��?\����ɑ��;����w��y�Q/�>��� 20��$������Gl����¾���K��h��Zb�xU'?f^���ǿ������޾)"??�?ۆw?;����!�tO8���>���<X�ȼ��:����ο�M��[`?���>
��0ˮ�e��>9Ԁ>�Kb>0q>�0�������(<:�?b�(?<,�>��h���ǿv����Ax<C��?/�@TxA?�(�	���*V=���>S}	?��?>B�1�7\�9��|M�>�8�?��?�iM=ĳW�b�	�Ewe?\��;�G��޻��=mK�=�=����J>�h�>���XA��_ܽ��4>~�>f�!�#���J^���<H�]>mս�x��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=��^�ƿϰ$�F��O=]R���W��$�Aԩ�ыV���Hp�rH콙<i=�[�=9xQ>��>��V>\�Y>G~W?��k?A�>�>ē�&����;���h�����h���q�T�������B|	�������iʾ'=�&��=�R�����Ѯ �E�b�ktF�e�.?�j$>��ʾ��M��P(<?�ʾ����ڧ����^̾Г1� n�]Ɵ?��A?�݅�u�V�AD��4��`����W?r�L��S���Ҁ�=����R�=�>�=#��M*3���S��j0?�k?$>���z��7#)>g� ���=m+? ?�XQ<�?�>E%?D�*��_�>�[>�&3>$ۣ>�C�>��>Ԯ��P۽�q?ڄT?���0윾�#�>4q���{���b=4�>��4�C�� �Z>ݦ�<xa��R�Y��׎��3�<��V??�>+B*��s��7��8�_S5=�&x??O?T�>v�j?Y�B?��<����4T����W�l=3W?�{i?v�>�W����оHƧ��5?�Jf?ErO>�i��D�./�����?��n?{?j���o}����L#���6?��v?0r^�rs��=����V�X>�>�Z�>@��>�9��l�>�>?O#�FG���]Y4��?S�@���?��;<b����=�;?�\�>i�O�_?ƾ|��������q=m#�>����0ev�����T,�$�8?Ӡ�?C��>2������K��=w�ܾ��?p�?�aپ�p��#�(���-������ҽy�=��W���@�5���E>��H��A�(����?�+p�>H�@�:�XL�>|/P��g꿎�ؿ������
����$?���>�=��̾�ǆ�k6��9�D���H�nP��^�>�Z>NE�������{���;�ُ��s��>���$�>�S���ӝ���
0<P͒>�N�>��>Q갽I����?*D���ο����,��4�X?�M�?�x�?:?�1<��u���{�v��HtG?��s?�Z?�M$���]�_;��h?�s�G?d��G�x�B�X~�>,4?I��>����@>��>[Ϝ>�:>�6�g]�������]񾼘�?���?�Ҿ��>u*�?�f.?2m�?�������%���	�I?⺾=q��� 5$�+�L��r���?��&?v3�42�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�8�>P�?��=3�>l3�=�����,���">5��=T�@���?əM?�#�>�B�=!{8�@/��8F�RR�]J��C����>��a?��L?��a>C︽�h.�B!�Zuν��1��w�)�?���)��^߽��5>nc>>�>�3D��+Ӿ/?r&���ֿ�2��Z���7v?GM�:-�>�u �>T3�_�X=p��>n��>�5
�����S��!s��L�?��?���>�y��т�=�ay=��>��> 	 ���%͛�+��>5�2?�ǂ��<W��+c�	>�>Z4�?h@��?��d��	?���P��fa~���87����=��7?t0�T�z>���>��=�nv�ۻ��P�s����>�B�?�{�?,��>�l?��o�7�B���1=9M�>��k?�s?CQo��󾵲B>|�?!������L��f?�
@{u@U�^?%�������� ��g;�X>�54=¬]> �f�_�)� {�����=�����)9>MY�>8æ>*7�>�f>&�U>�6>�����7��?����:�7 ���	�p�����*Z�����R���^��b���U&߼�>�2h���^<����<њ7>�N??�4?	�M?/~>ju;��o�>�s�u4��ԾX>�	?\�S? G-?�1?�=d>�%��O��	�������k_�H��>�n>�l?a�>���>�V�=�"�>פ�=w��>-�1>��'=���=�Y����>a��>J��>S�>�C<>ݑ>8ϴ��1��h�h��
w��̽#�?����L�J��1���9��Ҧ���h�=Ab.?�{>���?пd����2H?%���t)�ȹ+�?�>|�0?�cW?�>L����T�F:>+��{�j�a`>G+ �6l���)��%Q>\l?�Jg>o�u>7P3��?8���P�����
|>�5?�߷�':��Tu�xYH�>ݾ�M>���>�uG��(�����ZD��i�b�y=[-:?+�?봽����C8s�����ӫP>nH[>��=�)�=ʞN>_�b�p�ýwF�?�.=7�=�A]>#]?�]->�ٌ=���>�\��ȅN�O��>ӉA>��,>_@?�%?)B�P��7����-� �u>m�>؁>/�>ڱI����=���>{�b>}>��������?��V>��t�;N`��v�G�r=wD���?�=�p�="� ���<���%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿv3�>/|w<@���y��-����>tk>o�?�߾�N<��������>k/�>��
����!�ѿ.����D�>z�?��?�8��ɗ��+7����>�?ygD?�=n{���9��[��>��>}�X?��>�;2`��,�>�0�? ��?{D>X?�?ld`?�l�>8�;�42�����g��_k8=� =�&#>�<>������S�M������6Lc���v�Z>F�U==G�>�AP�]Wվ��=�!��XkǾd�^��8�>FiS>�Ɵ>�>]�>C �>p;�>i����<S���,)о�K?��?6����m��L�<6��=3X^�4�?�V3?��n�d0Ͼiި>�_\?��?��Z?y�>��:���￿W9�����<�9K>ɍ�>�y�>��sM>pQվ�lE�m�>س�>�B��پ3聾%�a�xԝ>�;!?��>�=��?�$?�b>�[�>�D��L����J��T�>�b�>�a?��s?�?`����5��ה��硿ç\���6>��w?X�?;F�>����ˣ����ߘ���@��l|??�a?|Ͻ�?�`�?P�??��=?�ra>WJ?�.׾�{��W��>#�!?�&��tA�D3&�V���1?v(?LA�>�"���w׽�tҼ'��`R����?�\? &?�g��Aa���þr�<`'��9b�[�<��Q�p�>A=>�]��n�=bB>��=Gl���4���i<�ž=��>��=5�5� Q��6=,?��G��ۃ�>�=��r�xD���>�IL>���Ŭ^?~l=�8�{�����x��B	U�� �?��?ck�?K��$�h��$=?�?w	?5"�>FK���}޾O���Pw��}x��w���>���>�l���.���ڙ���F��C�ŽW����>��>�?�?�a0>��>z@���.$�A�޾��V�U��Z��j>�W2��������,��P|����&e��7�>������>ʝ?A'U>��i>@�>�H�����>��Y>A\>'B�>/IY>+s >��'>�FW���$�,IR?B�����'����l°��@B?6_d?��>3�h����$��Pj??7l�?bv>��h�h6+�qq?�U�>���Wq
?$a:=��້<�O��Ĺ��9��`�����>� ׽�$:�HM��Gf�o
?+/?�-��!W̾WR׽e}���+=◅?��$?��'�>Lt�]l��˃3�>�5��k�E&��Mq-�)�.�|?t��W��T�r�m���-�@�\�e=B�'?=X�?�W6�����]z��r`�8�Pa�<]�? ��>ep>/�>G�оYC���p��b� L�&��>� y?��>ۖ??7??{>J?�<?pu<>���>����X��>#����R�>�
?s?F/?��2?��?��.?>>�퉾�	�4���j?��?>�.?�_�>���>�@���=��*>B�O=kB��D����	��2d	��)��S��S�=�>�w?���
9�>���@h>�68?r��>��>������}�D�<���>��
?X�>������r������>籂?%���~1=�,>8�= ��������=�yȼx��=�MA��2H��<�_�=ۉ=��Y�,^;�;9l;���<,u�>[�?(��>�B�>�@��ϩ �����d�=}Y>�S>>�Fپ�}���$��_�g��\y>�w�?�z�?��f=��=0��=y|���T������������<��?�I#?#XT?��?��=?j#?��>+�2M���^��$����?�!,?��>7��F�ʾ+��3���?pY?z9a���4;)���¾��Խ��>�[/��/~����D�K���������p��?$��?�A�f�6�Iv�����\��B�C?�>�Z�>��>��)���g�5#�y*;>V��>�
R?�Q�>`QO?��x?��Y?MG>n8�׏��c��%0	�X�>�P???�Q�?I�v?���>X>�#��0⾿G ��2&��p���ǀ�n?x=n:Z>惑>.o�>�>��=/�˽&��,#2�ö�=z�d>`c�>�Ū>��>��}>l��<��G?���>�e�����&菉����z=���u?;��?��+?�g=#��@�E��N���A�>Lh�?��?�;*?>�S����=S�ּ7Զ�.�q��#�>�˹>�)�>���=�?F=R}>)��>Ԛ�>�8�3h�zm8�EM���?\F?m��=hƿ��q���p��җ��d<Q풾=�d�t����Z��_�=�����M�����[�ǡ��r|������2���w�{���>��=E��=���=C��<��ɼm�<�*L=�n�<h�=hp�"'n<.69�hy˻N(��>��C�Z<h�H=�`���ƾ"Wy?��K?�,?�jE?��d>�(>�D�(�>�NH�5^?:�[>���5W��T"(��Ꜿ�X���2Ҿ�۾Ɏd�d���>�F`��>�72>��=z8=n>p�=s�^=er��h0�<�j�=x=�h�=|A�=.>�43>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��=>��>�[O�+�/�
g��g���U�H�?9F?�v�Ͼ!P�>���=a2ܾ��þ��S=�93>f�m=l�#��_�L'�=�����D3=�m�=� �>_B>
��=if½�D�=h3=|�==X>�I<�;0�
N�I�k=m��=��m>A`>�Q�>F�?�Y0?8+d?߹>�Qn���;�����>���=C��>�[�=��B>��>V�7?��D?@�K?�ڱ>R��=��>p��>�
,��7m�'#�`������<Y��?�Ն?&I�>=�c<ӝB��h��r>��Ľ�?�0?RJ?i�>jv�	�9!>�%�6����;���<��=�������je�^u��KԽZ�#>���>���>���>�	O>��>�Ee>3��>�*>_C�=�#M=��Y==�=�*��z���!�<N��=�q.<^kr=+P�����)ƨ�5�߼q��t���<.��=���>��>���>}�=�����1>#B��ˬK���=���@�t.b���~��/���8�c<>�bU>�bt�Ա��	:?:�Z>�@>��?:�s?�I">p��Kg־W�΁a�CXM�';�=.;>��<� �:���]�^�N�7	־��>̉�>�0p>���>2��C�I��=s6���$�{�>^r��X�o�M)���{�8��� �;j�0����%G?B��ߙ�=+
o?,3A?Pd�?Y�>�fW��&�=&і�;p=+�侁����ӽ,�
?ޮ?
�?`l	���W��C̾�����ڷ>*<I�(�O�-�&�0�����ȷ����>������о�"3�^h�������B�Rr���>��O?��?�(b��U���WO�����$���k?:|g?*�>NJ?�D?�&���y�k��=��=��n?��?m:�?��
>�Խ=�t��sT�>�7	?���?K��?z�s?��>�^�>�s;�O!>7���Fv�=��><��=�>�=߈?ו
?��
?X	��X�	����񾂴]�A�<�'�=|
�>��>�r>��=�f=�n�=;�[>q��>��>2=e>���>KM�>��۾��%-?���=	��=�)?�D�>Ya�>|I>�<>��
�3h�U���^��@����=e숽pE��u��5	?�Aҿ)��?���>v���?l���wϽ�MF>�(�>E�]����>���=��=1�>���>T�ú��>�i>�߮�c]O>����)��iB��RV��	�i�Q>70�Ef<����;�4l���޾V�'�]�t��n���[C��0�=<��?[Ǘ��@���aK�\�P�߅=?d��>j�?zG��lO"����=���>0{�>l�߾�䅿������?���?�;c>�>��W?�?o�1�I3��uZ���u�:(A��e���`�H፿霁�V�
��	����_?��x?�xA?�Q�<M:z>H��?r�%�ԏ�g)�>�/�k';��E<=U+�>*����`�2�Ӿ��þ�6�6JF>�o?O%�?Y?�VV�E3s���>
�H?h@.?�u?D�
?lL??�>��d^?�x-> �?�?}�?l�.?sP?<r>�WW>�I=DM�@a���땾$ᱽ����[�q�xe}=��=g�>ė=���_�P�������f�=k=��:{}<���=��=�c>궦>ĝ]?�U�>	��>�7?���MV8����
/?�9="g��1ꊾ����t��->4�j?���?hKZ?��c>��A�V�B��\>�]�>:�&>��[>�D�>�=�	&E��=dE>�>��=�:N�Oց���	�O����&�<��>���>�=|>J���b�'>�i���Kz�3�d>h!R��Ӻ�M�S���G���1�dv��<�>��K?��?o��=_龹V��\>f��))?�[<?NDM?]�?C��=`�۾9�9�K�J���*�>�ܩ<|	���� ����:���:��s>53���h���	c>_e�<<޾^%n���I�ߐ�o�B=`����V=A
�z�վʒ�Jy�=��	>����� �$���̪�oJ?ԟj=uG����V�(�����>S�>�H�>�6�љ}��@����t��=�m�>;>y� G��A���>�^G?-^?o�{?h�_���h���;��r���žx���i�	?k��>v�>�y�=cӄ=+p�����=>l��^K����>,Z�>�l�P�(?����վM�0_�>�W? ��=�V�>[xR?�
?`�n?��(?mF?f�>�*'�=x���*?_�?�A�=�����H�<��H��*�v>,�?��!����=�^�>�"?��?u�=?�O?�wC>�e��>\��I�>���>:�S��C����=F"1?�F�>Aj�?��?HU>�h��ιbU����>���>��N?|D?,dE?mwz>ar�>���m��=��>��e?��?��r?�S>Q�?T�>]u�>�<�=�K�>���>��?o�N?��t?��J?ʧ�>HB<�x��oј���J�Q� <g�<��<�=<y����f������<qa���f1�����@#��yj�_���q8;��>H�t>�͕��31>�xľ<ሾ�<@>G���윾m����;����=�M�>�e?�S�>�e$�s|�=�%�>:*�>���S(?8�?�?��;_�b�o۾X{M��q�>R8B?���=��l�������u�(�m= �m?��^?��X�!(���b?L�]?�[��=���þ�Oa�-��'�O?��
?�aF���>�~?;r?���>��f�o{n�0��O�a�
�h��k�=�&�>;��id����>�b7?)R�>��a>J��=�۾z�w�Nğ���?G��?t��?��?��)>=�n�A.࿙����鑿�^?��>k��J�"?�λ�o;�m��`p��x�߾檾�7��b��
Q��#� �' ��w��>��=�?Z�q?6�r?V�^?Sh �x�b���_��b�l�S�G�����D��)E��B�?o�q�����pĝ�&�4=�\�?F�,��?1I ?����Z�>9����Ⱦ93ƾ[�>�`���q=�#�=Q��>B�<���=E��`mv�N����m5?O>�>�\	?�0?�r���K��yi�IG0�C��e��:�7�>�g�>�9�>6D=���4������Զ�����z>�c?@K?��l?#~�60�Ϥ��	6&��|�����3@>��>�N�>��d�4 �K&�^<�:�t�[�0����� �=Ƭ.?�Iy>�Z�>�?�,?n��������-��,�<'Ǿ>��f?��>>�>C�Žw#!���>9m?s5�>�r>f3������y�v_ҽ�?�>��>DU�>�3>�j��;Xb��C��������B��>1�w?p,v�@�c�C��>� O?#�:=��<'��>�D^��'�W���b�iG>V5?j=D�h>E ���r��sl�𒾼�.?G	$?7�`��UD�ӄ8>Br?~/?n�>>y?��>(����s��+�>�([?>�T?��??hr?�a2>���D鉽 �k�k�l=�)?��=>̣Լ��K>f/C��AP���p�a|>�n�>ne=-�'�[��<=��=��=� <>�>�hۿv?K�R�پ���w3
��ǈ���������s	�m;�����cAx�eu�-&��V�@(c�u��� �l�5{�?/1�?F�����񠚿ӂ�����ʋ�>րq�M~��뫾�B��U�����ˬ��d!���O��5i���e�͜'?9Z��*�ǿǲ����ܾ�3 ?��?fmy?����r"��V8�>���<?^����ģ����ο���_?$��>=��nt�����>�т>@�X>��q>ġ�J��Д<��?�q-?%�>�lr��nɿ;����1�<���?�@}A?��(���쾵�U=���>E�	?��?>�y1�gK�Z����E�>�8�?C��?�M=g�W���	��|e?��<�F���ܻ��=��=�=�����J>N]�>j\��9A��ܽ�4>-�>��!�E���k^�N>�<��]>?�ս�'��5Մ?*{\��f���/��T��U>��T?�*�>Y:�=��,?X7H�a}Ͽ�\��*a?�0�?���?&�(?7ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=V6�щ��{���&V�~��=Z��>b�>��,�ߋ���O��I��W��=���Ƶ�>�%�H"���&	=aY��e=4�~����\ꕾ=)���ֽUa�;[>�\k>jke>'|>�Tc>�C>�@?�hX?���>S>	�����ν׷���R���k�����>�c��ǅ����3�M�侭����@�:�jB �~!=�d�=�6R�	����� ��b��F� �.?Ay$>��ʾH�M�4�-<�pʾ����9΄�7ڥ��+̾ǖ1�i!n��̟?I�A?������V�A���W�E��z�W?�L�ݺ�J묾���=,���ե=?$�>,��=�⾀ 3��}S��1?w�?��.A��e$>���G�=�o)?�B?˷�9 ��>�(?���U�ýN n>��E>C��>(f�>kS�=[ ���^��x?(K^?-��T՛�mS�>=Ѹ��Dz�1�<==�>��e�6;��H>mS<!܁�����T�h��F=d�W?͍�>��(��'�O�Ǿ�=/���^?`R?��>�j?�^?dLֻ�����d����3'&�j�E?��|?�i>�^��s˾�V��n�6?ؒd?o��>ܓ1����%�CI��a
?��?�?;(�<��{����m�Ǿ�V3?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>��������>`圾���?	��?���'��4�qdO�A�ɾd�%�GH!>��ջ�����;/K=����O9�j�ܾ1#�/��>�@�#{�g[�>�8�qx�Kj�`@��^m{���N��L?���>`v7��)�(+���Ό���Z���=��<P�s��>̮>-x���ē�Vzy�Az9�,����~�>"�)��%�>ͻY�-[���ϟ���; k�>��>8ˆ>I���h%�����?��&�Ϳ{=�����lX?�?e|�?P�!?(��;m�z���y���»�J?ځt?]�[?B%���P�&yD�GTk?6��<�[��`6���C�t�z>��'?�G�>�)+����=5��=�&�>ThX>��6�2�¿�c���P�J��?yr�?��"�>hH�?�.1?�F
������q����,���,�i�-?9>�ڥ�*v �R�;��jl�B ?��&?m(�S&�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�$�>��?cn�=�a�>Lc�=h𰾐-�[j#>��=!�>�J�?U�M?oL�>�R�=o�8��/��[F��GR��#��C���>m�a?�L?�Lb>����2�
	!��xͽd1�LL��W@���,��߽�)5>g�=>8>�D��Ӿx�?
j�Ɣؿ�i���y'�84?p��>2�?����t�ɇ��6_?���>>:��+���'��	X�\��?�G�?0�?��׾/̼�>��>G�>2�Խ����{�����7>��B?����A����o���>a��?��@7Ү?�i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*�������f�־�����W>��>i�Y>*Q2=��2�����X�+>�">���>�?f��>2�>>;�>)�>հ�=��{��� ����놿^�;�r�=���Y�ܒ$�2�c�ݾ�.��A��]���'�۽���=c�B��`�=��8�G�=��U?7R?8p?�� ?_�w���>1����G=�#�q��=+�>�N2?ϚL?�*?�̓=՟��>�d�x]��[)��Y������>~|I>���>�J�>��>���9��I>@R?>�p�>� >�&=��꺟�
=�N>�a�>���>�w�>�C<>��>Fϴ��1��k�h��
w�p̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��t�T�4:>:����j�5`>�+ �~l���)��%Q>wl?��f>u>��3��d8���P�<z��l|>�26?t궾�D9�ݿu�]�H�gcݾ�HM>�ž>�D��j������gri��{=�x:?�?:+��5ా��u��B���QR>n=\>�[=�]�=�PM>	ic���ƽ�H�t.=\��=ש^>a?`B,>(��=@У>�1���`P���>BB>��+>f@?�%?����e��_{��,n-�6w>4s�>��>J�>�-J�� �=�F�>e�b>RA�Ã��t�!�?��?W>n�~�z_�Qs��z=HI���Z�=�˔=6< ���<�˽&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿh��>���:�p���T��؄�<88>�^>�#?��vE{=d/@�=QW>T4?���������οj��y(�>=��?Cs�?V�V�������&��B?:[�?��b?���>�E�����Y$�KV?�]w?۱�>Q�Ҿ�x�
.	?��?DEo?A�t>�?�$c?���>�f=�*��*��+D��O ��|>#]�>��5<��~+Z�A���Yۈ��
`�e2����=�A=��>��g�M����\�=쿵�:������A�>�R7>/u>��>ȕ�>��>��><�=�%I> ś�������K?忏?R*���r���<�_�=�,V�h3?��4?¢m���Ѿ8�>��Z?��?>�[?�!�>�B
�.��v��d�����<'�F>LC�>���>l͓�8T>hƾ�/��<�>>� ���پ$�r��p<:��>��%?ea�>��=i&?d�.?`P'>!5>�vu�K��;Fu��{>cE?e5?Kr�?Fy>��*�!#C�O]���|����s�%����?�?)�>r'���ۜ��{{����>k�=0�U?��B?��=���>��?]�%?�i?H9>o��:ؾ�Z=�?��!?��*�A���&�n���i?vQ?�}�>sU����ҽ�.ݼG
���==?=\?+8&?���m�`���þ��<���HP�w��;�aN�ۥ>F�>�B��汷=7>�3�=D�m���6��x<T�=fВ>���=ib4����0=,?��G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>$�l���K���ڙ���F��_�Ž�4߽�5?)?�>e?��?�/>|T�>��ݾa�;��������X������D���'��M����`����g��꿯��m�Jؘ>���7=�>�J
?n�>��>�N�>1?���U>�}>6O�>�#�>]A>��}>{g>��<���GLR?�����'��辉���w4B?�nd?�,�>K/i�g������]?J��?�o�?0v>��h�/+�qm?�C�>o���o
?{l:=�8�ΐ�<�V��a���S���@�A��>�C׽�:�AM��pf��l
?`2?�����̾�g׽ WZ�r��=���?�Z$?M.�xe��礍�-�P������s��Jҽ�wM�z�.��|o��i�������G����=��9X=�#?�m�?{�>�� �L�̾X.[��w/�'�=�n�>΅�>�q�>'�=����?� �y��kU�ej��1S�>dm�?�>�>x{9? �?l�j?��@?9�C>	 ?1�\��K?v���0�>�3?��J?��!?e�4?��)?#�B?�>�\�% ׾����?"NI?3-?��>�P�>� �iYI��OH�㉚��Q[����=$�����	� ���Q�0��g}>,`?}ͽ��6���z-A>��=?`�>-��>⁍��0���(�{�>�?&a[>h���$�eZ�h��>!�?��1R<�F4>\�>*�<S/���	�=RS���=�<�B��z��#P�=4.�=߄E=ځ-=��<}���Ek�!��� u�>6�?���>�C�>�@��/� �c��f�=�Y>=S>}>�Eپ�}���$��v�g��]y>�w�?�z�?лf=��=��=}���U�����H������<�??J#?)XT?`��?{�=?_j#?ϵ>+�jM���^�������?c#,?��>�����ʾ��<}3��?=W?6a�u���?)�Y�¾h�Խ�>x`/��6~�����D�>E~�7��Ȏ��ӗ�?���?��@���6�i辶����h��͐C?&	�>sn�>�!�>��)�(�g��!�N.;>+��>�R?�z�>?P?��z?L#[?�V>�j8�ޭ�SJ��PℼL%>\�??�'�?�S�?�]w?��>E>*)����C���_��������M=��W>uВ>H��>ũ>-|�=W�ѽ�߳��;�O�=Uod>Y��>���>��>G"w>�y�<��G?��>"a��iG�����A_�������s?E�?�2*?��=M�g8E�M��O��>���?x��?$]*?!�a����=����Ɗ��q�]����>^&�>dݛ>?ѝ=_�==�>�3�>�=�>�@�v/�� 6��3�e?��F?x�=4�����a��(�U[e��I�=��5�0�bE��Pr��b-�<�|`�aFQ���ƾ�WD��g]��K���R���¾����F�>o�>}�o>��=xE->͉5=�vh<u��=A9�=`��=G������ٌ�v����F�< X�=7�=voۼ��˾V'}? .I?��+?��C?�nz>J�>G�3��ԕ>��8?CU>�FU�;X����:�Kz������4 پ}�׾�c�d(���D	>�hG�,8>��3>�
�=��<�(�=�~v=�=��w�P=�e�=��=�t�=�=� >�n>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�67>R
>1�R�{1��U\���b���Y�	�!?�5;��i̾�>�>&
�=��޾k=ƾH�0=/�6>��c=�"��E\��=�nz�a7==�n=���>@�C>�Ѻ=%,��KT�=VI=�=?�O>^���9��,��3=i��=��b>��%>~��>?�J0?d?N)�>}�m���ξ^?��uR�>��=�>=�=�mB>C��>�7?!�D?�K?�l�>:k�=X��>��> �,�U�m�7p循ʧ��s�<$��?dԆ?vи>O�V<A�A�����0>��ý؁?Yq1?��?�̞>���0�ɿ��M����#_�-<J�#�>0�>���= � jM��YM>4���A� ?�?�<?��>��>\p0>^E�>G}�>�<=xe���������W��;�{=9͹q-����g���#<m�y=NϼJ��=���_���G����=I��=t��>�<>���>���=���"C/>)���f�L�4Ŀ=�G��`,B��4d��I~�"/�zW6���B>�8X>Z��4����?��Y>l?>i��?�@u?d�>$!���վ�Q��=Ce��US�kʸ=Զ>!�<�cz;��Y`�g�M��|ҾQ]�>���>u��>�`>l���龯���/��	�L���>����ӯ�]
��Z��*q���'��J/��蜽!�:?��k��X�==%g?u�G?���?i�)>�߽��/�ki2�Y$��tbW>�f�����!Y��XXA?�5?R�?��#��'���C̾X���ݷ>�CI���O�g��0�
D�.ʷ�/��>����о�%3��g��������B�aSr���>�O?��?{4b��W��LVO����v���r?�{g?��>kJ?A?? 6���w�p���t�=~�n?1��?�<�?>=��=����;�>�.	?���?|��?t�s?�h?��w�>�x�;� >�����?�=*�>c��=�;�=6t?;�
?��
?�T����	�a�����^�z��<̡=���>�o�>��r>���=�mg=�r�=�0\>�ў>��>�d>? �>�M�>���Ή��1?�T">0/�>�1?�Ӕ>@��=��	��0�=5*��耾��K�/��� 핽�g,=~��Q��<4!��?�bÿ�J�?�W>=\�3�?��x�E���^>�>�$���>�T�>)E�>:�a>Y�>�u#���>�(>��о�>�b��!��ED�z-R�B�Ծ��u>7���9y!�1�p� ���N�@�����x�j�}m��J�=�� �<�ُ?g�����k��+*��� ���	?6H�>�d5?$��_V���_>y�>t��>���� �����r���?��?�Kc>�#�>��W?T�?�x1�^3��oZ���u�b2A��e�h�`��܍�E�����
�G��2�_?��x?�eA?6�<O;z>@��?��%�cꏾ1�>]/�;��==t<�>q<���a�؜Ӿ��þ���~[F>R�o?�$�?�]?�aV��A=�A >�1?�qg?��?-�(?�&V?��=ˀ:?I��=���>�S?��2?��/?2c?�Z�>��v>�ӈ=A����Ϣ��7��c\z��Iǽc�<���=�g�<�<�G��>�s�=��$n���<i;��+��<m�a��xX=�R�=R��>*�]?��>�6�>�7?� ���6������/?2{4=�����������GB�a�>0�j?=��?L�Z?�_>��@��JE��$>g��>T'>�uZ>���>|���E����=tX>u8>ث=�yT����X���O�����<�!>5��>�1|>���Ͷ'>%|��p0z���d>��Q��̺���S�[�G���1���v�HY�>!�K?l�?t��=�^龒/��If��/)?�]<?�NM?��?u�=Q�۾��9���J��=�o�>�a�<��������#��d�:�A�:�s>#2���ݠ�aWb>7��#r޾n��J�
��8M=���SV=�U�վ�0����=�$
>#����� �H��v֪��0J?��j=w��+aU��p����>	��>f߮>��:��v���@����� >�=��>� ;>�T����~G�:8��>��X?ʲL?:{?c�����~���D�q�#�������C��3?� w>?w#?	{�=�;��"Ͼ�t���_��6�>�>�N�>�l&�PM`���W�s��*^4�A�=9��>#��>��?�xd?^�O?��?��H?�˯>
�>�D�=��־`&?%ւ?�ф=g�˽Z$Q�̫7��C�|N�>s(?�H�喖>,�?��?'�'?��Q?Gs?�\>~� ���@�K�>;͊>�W�S˯�X�b>^>J?Rܲ>9qY?_��?j�<>k�4�'���Yq����=�>��0?�o"?t�?1�>�?[tU�{���+�>��_?�@t?�Ǉ?�>Q@V?�_$��u�>��Pm��Q�>�'?�x?��~?��N?��?F�O=L�;�{�<#�f��j�;�0��竽Z[�������+�>Y�E>����2��.my���S���w�
<�Z>�[�Ld�>v�s>W���u�0>��ľD7��A>�>���A��t9�:����=ǁ�>b?ݵ�>�6#�mْ=F��>�,�>����,(?��?�?t});C�b��ھ�K�V	�>J�A?{e�=4�l�^���Y�u�!bg=��m?<�^?�bW���+�b?��]?#e��=��þ�b�Ћ���O?[�
?^�G���>_�~?��q?���>��e��9n�4��KCb���j�/ζ=�q�>&V���d�>�>ݜ7?�R�>��b>��=�u۾��w�.m��`?�?�?v��?<,*>��n�D3�X5	�����K?�W�>�Y��l:?ؓļ(f����5;�շ�<�������T�� �P˽b�8�W��=F�=�?g:~?T*�?�\a?��3xz��d����/K��<�90�W�I���B��$Z����y'_�(�����`@k>m=��A��z�?b�'?s/����>w���"���@;�YC>y����Yܞ=&����A=ٸ\=#(h��j.��l�� ?��>�r�>��<?��[�>�v~1���7������N3>Kw�>�B�>��>lT�:��-��齩�ɾ�W��q.ӽ���>��q?FNM?�`Y?�������`�-T��P�_#��‐>�@�>�^�>� ��B+��-���f�b�h���������=�d9?d5�>�"?�?*��>�t��O-�`�ؾ�]����mT�> F/?x�>�>Rah��@*�:T�>��_?��>m�{>S�
�>R�my��"�=B?�|�>�KQ?zKJ>�.ƾ��h�����$����N��!>VH�?��d�����F�>~q�?>�=�Q����>�Ħ���W���#�f���'�;a��>��;�U�=�����j ���x��E�G�(?�E?��&��U�>��!?�"?���>c�?�p>ž�U�U<��?�`?�BJ?uk@?L��>�ύ<� �������W$��_M=;5�>�fm>���=�z>����(�J� ��D�<r�<����%� ��/����
�=[Tv=��I>5mۿ�BK�m�پ�	�5?
��爾ʨ��(d�� ���a��I��$Xx�����&��V�7c�ʢ��	�l����?�=�?����K0�����%����������>��q�Ɔ�c������2)���ྻ���fd!���O�g&i�\�e�P�'?�����ǿ򰡿�:ܾ4! ?�A ?8�y?��7�"���8�� >MC�<-����뾭����ο@�����^?���>��/��o��>ޥ�>�X>�Hq>����螾x1�<��?6�-?��>Îr�1�ɿc���}¤<���?0�@�lA?]�(�[@�ڦY=H��>�~	?2O@>�2�;��s����>-C�? �?~R=�}W��U�We?�s�;8G���ໞ�=פ=��=^��1sJ>cF�><��?�@���ܽHa4>�̅>�`"��(�e�]�̆�<�v]>��ս;i��5Մ?*{\��f���/��T��U>��T?+�>t:�=��,?U7H�`}Ͽ�\��*a?�0�?���?&�(?3ۿ��ؚ>��ܾ��M?aD6?���>�d&��t�ǅ�=�6����q���&V�f��=W��>X�>��,������O�J��H��=�^����ƿu�)��"����=��=C�b�����	�)��<O����.��TFֽ�!|=��>��q>?u�>��r>�>DO?�&[?dq�>�� >]�˽~ui�B�Ǿj�;j����g,�K�����E��I���侬;� w��A��e��w��4!=�g�=7R�p���(� �<�b�E�F���.?�v$>��ʾ��M�6�-<�pʾW���Mۄ�*᥽�-̾ח1�"n�S͟?��A?������V�6��W�����C�W?OP�����ꬾ���=����c�=�$�>���=���� 3�c~S��u0?�!?m����'+>�P����=��+?V�?��J<��>��$?�1+��H�)(\>,5>�F�>ñ�>Zg	>�Ѯ���ڽ�~?:aT?�� �t���y{�>S��OUz�z�f=�:>�7����z"Z>��<�쌾`[��#��Gs�<?W?\>�)��2�y���%�!�c-9=Ƶx?��?4��>��k?��B?1֞<������S�6"�Su=��W?�ui?V�>@���оTΦ��i5?�le?m�N>,Pg�Y���.�G�>Q?��n?�F?�T��GJ}��������086?��v?s^�vs�����4�V�l=�>\�>���>��9��k�>�>?�#��G������rY4�&Þ?��@���?��;<��X��=�;?n\�>�O��>ƾ{������6�q=�"�>�����ev����R,�c�8?ڠ�?���>�������@=@v���7�?W�?�ɾ��f;����1Y�l�$�P��=�ϴ��:�jO� ��1�>�+U��j����M��;��>�@���=e:�>�t߾������޿�̔����t�+�0?���>��o�<�������ϥt��[�����M�>r�>�������l�{��q;��+����>C��	�>~�S��&��_����z5<��>A��>y��>�)���潾ř?�c���?ο>������O�X?h�?�n�?.q?J�9<��v�ɐ{����U.G?ĉs?rZ?�k%�=]�J�7��j?�^��IU`���4��HE��U>"3?HC�>��-���|={>w��>�d>�#/�Y�Ŀ�ٶ�����$��?��?�o���>���?st+?i��7���[��J�*�+�/��;A?�2>ۍ��p�!�-0=��Ғ�;�
?�}0?Q|��.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�!N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?C�>��?D��=q@�>z�=v��I�3��K">�i�=�<�	�?$�M?=��>�'�=.�8��/��DF�ER����C�s��>q�a?�fL?)�a>����f.��� �*�ͽֳ1�N���?���,�a�޽#/5>-J>>�	>��D�;Ӿ��?Fp�5�ؿj��;p'��54?"��>�?��|�t�����;_?Az�>�6�,���%���B�^��?�G�?<�?��׾S̼�>>�>�I�>:�Խ|���L�����7>:�B?S��D��k�o���>���?
�@�ծ?bi��	?���P��Va~����7�c��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?RQo���i�B>��?"������L��f?�
@u@a�^?*�ԿSޗ����H�־�&�=�u�=��s>#�y�K>��>�ѽ� �Հ=�B�>��p>��~>�ɹ>S��>
!�=����#���4Z���� ����[�
���]��T⾌�Ὣ$�gC羔����e�=��t<��'�����ʽxr6���>�d?��/?�2g?���>�E�="��>�.�<a3������7B?�Oo?���?��?�W�>�Y�&��R�w�0S��◾���=y�=�;>..X>���>tg{> �>1�=�r�=\k�=��=���=Ti>�F>�l>CJ�>
^X>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��w�T�3:>:����j�5`>�+ �~l���)��%Q>wl?J�f>4u>3�3� e8���P�y���i|>(46?붾�@9��u�S�H�DbݾHM>�ž>��C��j��������si�C�{=�x:?��?}4���ాR�u��B��|OR>�6\>�3=�[�=�YM>0mc���ƽoH��_.=���=w�^>^?��+>^��=.�>O�����O�ͥ�>;bB>�,>x�??�%?�������A��E�-���w>�`�> �>�e>`AJ�l��=�q�>��a>_y�Kۃ�����?�NSW>c�{��$_�EMv�	�x=��� ��=H�=J� �8>=�~�$=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>�`�$W��9���u�t@#=���>d5H?N��C�O�e>�o
?f?j�*���x�ȿ�v�7��>��?�?��m�@���@�-�>���?EeY?�wi>IZ۾pKZ����>�@?R?�%�>�0��z'���?�ݶ?j��?��w>�u�?s�h?��>��e�D�V�����k�}�O��<
����=�����㾁qm��?��v"���ֆ��5�]�>0�{=�ԩ>�HW�Gx��<]��<R���3��'%�>��s>�u>0�V>^�?�r�>���>�D>M�:v�R����K?0��?���)n�]��<?Ȝ=�$^��?�04?|�b�W�Ͼ(��>Ż\?UĀ? [?�r�>k��O2��ڿ��]�����<
�K>&�>wE�>�,��кK>$�Ծs�C��I�>���>E����ھA]��I]��e�>n_!?^��>	��=v?+�1?��S>e�*��_�痿�f��t�>��?�?`?�b�>?����U�|���z顿�{�|�>劓?\�?G�9>�c��e��ｮ=j	�����P�? �?d��<��A?�5�?�+?�H5?܁�>>^�=��g|��+�>Ӽ!?/��I?��#�d����?|?^�>(w��a��B�缦������
?w\?G&?'���_��0ž-��<.�s&$��� <ז���P">-K">�	}����=��>���=��~���E�'�q�^�=��>�y�=E�-��/}�1=,?�G��ۃ���=p�r�+xD���>JL>�����^?Al=��{�����x���U��?���?Xk�?���4�h��$=?�?U	?y"�>�J��~޾J�ྺPw��}x�}w��>���>L�l���G���ؙ���F����Ž0��L�>N�>�W?4?5�P>�p�>6����'��������]�4��]�7�"b.�;���K��+�&���
�����Cr}��r�>�ꊽ��>�
?ig>n�|>���>"F��a!�>�"P>�Ԁ>�>�>UX> �6>�=�$�;>�̽�JR?����s�'�2�辰���)2B?1rd?.�>Ni�����q���?!��?Gs�?�Fv>�xh��)+�vj?4�>���0o
?�S:=7{�J��<EN��β�s$��������>SK׽%:�M��wf��f
?�+?�썼��̾�&׽Vm��O	>�N�?�^?@�Z��8l��M���!H�IQ��=�/��rǻ��t3�͗�����������q��.���v\	>�4?�ߡ?�)�-��&�����~�>�K�p�h>��0?ъ>a��>���>[Cܾ��D�nSu��$�	ӾGu>��?!Ý>�c>?��2?LyI?G�P?���>O�>��&�>eӽ��>�#�>�2?��2?Iu'?��?�^?#��=��A��1ھ@�?G�
?�V?���>�?�9���s�����{o�.��\�޽�ż�i��;A!��b"|�U~ =:�o>�X?���2�8�R���� k>��7?���>r��> ��11�����<	�>�
?oJ�>�����{r�Ja��Q�>,��?���Ry=?�)>���=����FԺ�V�=���r�=&3��fr;��O<_��=���=}ht���x���:Cs�;li�<2u�>B�?��>�?�>�A��� �#���m�=�Y>� S>k>�Dپ�}���$����g�FZy>�v�?tz�?��f=��=��=�}���Q����������<Ĥ?�I#?�WT?0��?d�=?�j#?�>s)��L��^��2���?r!,?a��>w����ʾ��:�3��?q[?<a�����:)�t�¾��Խϯ>�[/�}/~�����D�������}��B��?D��?"A�L�6��x�#����]��Q�C?[ �>uW�>a�>L�)���g�m%��0;>ŉ�>�R?��>��L?��c?бD?�">��2�������&����>b<@?f��?�ۙ?�e�?���>��>o\������txT���齝v�<��<��H>��>3W?7Dj>;�׻�X�� ����왼-*9=я�>��>!��>O�>�C.>�.����G?��>���n��e���r����$��Ou?]�?B�)?��=�k�9�E�;��R��>�<�?6��?��)?�hS�i��=��߼�����o��F�>nԹ>dF�>;W�=�H=2>�f�>S��>�
����38��mE�/�?
RF?O/�=��ſjv�eX���z���m�<����oa�f38���h�A:�=��0���|��0S��ӏ��	��\}���M�������_�>��=��>M��=&��<��f��g�<5kY=�s�;ײ=�[��%a�;��������ɓ��Z`;�sd;lS\=C�r�ʾ
z}?�*I?�+?�D?�tz>ĭ>�e;��>׋����?��V>g�N��껾�c;��H���˔�'aپď׾��c��"��u>��G�ʬ>�z2>$j�=�!�<V��=8w=b�=����=���=��=Si�=���=�u>V�>�6w?N�������4Q��Y罨�:?9�>E|�=1�ƾ[@?��>>�2������eb��-?���?�T�?K�?�si��d�>8�� ㎽&r�=b����=2>���=��2�B��>K�J>���
K��΁��p4�?��@��??�ዿŢϿa/>?S2>��=�oR��B1���X��\���Y��$"?
<���Ⱦ�:�>2��=c�޾��ž(�?=�4;>N�m=cK�K\�6�=��w�p�N=R�t=3�>�#E>d�=�L����=�>>=K��=�oI><�a9jJ5��B��p4=G�=��h>�&>���>�M?��/?��c?A?�>q�h���ɾܹ����>N��=�Ǯ>�ʍ=�E>��>��7?�D?�K?��>a�z=Cܹ>�/�>t),�2�k�KK�b���I�<��?�b�?�	�>�<;�B�g����>��̽k3?Po1?(�	?��>���4ڿ��t��\����=]S�>���⬩>aO����>�ʽ�i�j�R<4k�>֧(?�/D>d��>�
�>l&1��#�>a��<tYt>
O�=��<�">�x���W>���tǀ=r_C=C�P=��;o��+��<Jr>�n��������P��=5��>JV>���>�]�=y��0/>n���&�L����=�2���%B��5d�~G~�|
/�5u6���B>%X>�I��l0����?^Z>L�?>��?v@u?% >�g���վ�R���se���S����=Y�>�=��o;��N`���M�:�Ҿ���>��>�M�>�L�>��1�eL�܃��/پ��-���>_�S�]��`�`�	}u�(C��🟿��o����-OK?Cۃ�r�>��?ĻW?�n�?��>��<�;��)V=K������6�$��kk�r*��sU?��?�w�>�� &L����$����"�>�D��i�]�����:���_�q ���W�>�c��1>��>?�����՘��wN�q����_�>Xa?f��?�?o���{���F����Z̼e� ?tMc?Ͷ�>��?��(?O�ǽ���W��c.>:cn?�U�?A^�?� ;>��M>�ߣ��	�>C�	?s��?�/�?�ǈ?	���>Yb��O���6��ܼ��(=V�>�ǅ>��?nS�>p�?�i��-�-t	���Ѿ'H���6=sȖ=���>+�>�O->��=-�>�b�=�ȹ=< r>���>�J�>܆�>�0?+���f�<#?cS�=��>jy4?!�~>E�=�7Խt]*=�XT�>E�U�'��R��?.ɽ�X"=�G�;TXm=�V��}�>�\Ŀ/��?`�V>J5�M(?�j�޿7��O>��G>���>?TQ>l�t>��>7��>��
>u>��,>�BӾv�>���Df!��.C���R�_�Ѿyz>����&�����z��TJI��w��:l�Sj��/��:=�?=�<&G�?s�����k�x�)������?2\�>E6?1Ռ����_�>���>sč>PI������pō��h���?[��?Q<c>��>�W?�?��1�|3�#uZ���u�(A�Ye�e�`�z፿����ϗ
�����_?��x?�xA?�M�<�9z>��?��%��ҏ�*�>^/��&;�.E<=)+�><*����`���Ӿ��þ�:�]GF>c�o?%�?�Y?�PV�����Ij*><�+?�-?��k?�+?6=?����?�Qr=���>4"?�~<?t<?��?Kg>x�=K����
���p�}6���������v��;�v�=X$�=TA�<R�=h�D=���<��,��1Ľ�ܐ��+��Ke��Q=z�=� >�ͦ>��]?C�>��>�7?ъ�SI8������#/?P8=ں��R"��tɢ����>��j?7��?�LZ?/d>6�A�
C��>�`�>)�&>�\>'b�>��z�E��և=l�>7>�H�=�yO�	݁�t�	����Y�<G�>�`�>y{>󒈽l�(>������r�1�l>Z	O�ճ���Z� ]G��1��v�i��>ԨK?��?�u�=R_�~Ɵ�,�d�χ'?�B;?T�L?iN?Y1�=�׾{o7���I��h�X
�>Z�P<�
�����^ա��~9����;L�y>Lʙ��젾:�a>�n��޾��n�7�I�5�羜qK=����	T=���,־:'����=%�	>�~���� �G���ƪ�a"J?�|j==o��A^U����e�>���>���>��=��w��c@��)��YO�=���>F�;>W��7@ﾀ�G�V@�/�>��Z?S�:?��J?�͓�	؈�w`c�F��UH�����=F?��K>�q?V&ϼ.��=�1ݾ���<S� �<���>�F�>���=�^��X�2�ƾ��M�C��=h!?�6�>�?��U?��9?)1�?��I?ϛ?�'?k^��c����'?'��?�i�=Ў���P���=��ZL����>C�&?���c�>8�?�� ?t�$?�P?�a?�.>�� ��<?����>>/�R�������n>�dI?�Ӵ>i�Q?�Z�?'�J>�.�O撾c��ۍ>9�0>73?}�'?!�?��>�p�>/3����Bf>�u?��m?�ކ?h�>��?��W>��>�����e�=o��>�=?ǫI?�]?��L?~�?$�=����I =��j=�lC�ݙ.�A/ӻ�#W��;��\ƽA��;x�=�k������j�����Wڽ�N>��3>���>�ix>]֚�}IO>c亾j+n��cC>������3���3����=E-v>$�?Ǒ�>I�$�d+�=�V�>2 �>}��v!?�?��?�y+=)e�^���B���>ױE?9��=;p��`��\�k�G��=3�m?VGV?rDP�M��Q�b?q\^?���[=�}xþ�2f�uk�ĹN?Ո
?�pC�j��>�P~?v9r?y9�>��c�
n������	b���k��	�=%��>l����d���>~u7?��>ξ`>K��=��پ��v������?�h�?.�?���?��->�Pn��߿"�����mgg?O
?n$���C?��p�[8������)ɾ�b�����o 5�r9�(tȾ�>i�)2����=�9'?��n?n=�?1K?J*��_�>#�\�y�:�X�èѾ��	�^�O�ȑ`��?��T���C�� :���̾=�������\�C��?�6?�ﾑ?Ą��:S�V��������4���o�6>FH�=��<�},>R���!��ؾHy?���>��>��?#��_�6����i��e��5�M>^Ȭ>���>�V?pc�<�+������+���*S��B���.�>a�f?KzG?\�d?ܝ�Ц0�!s��T$���^�+��� X>��">1J�>	B��#���"�φ6���p�C�>���c���X=]7?P�q>$Ƕ>FJ�?H��>Q���ƾWv����&��ڼ��>��_?|D�>a`�>�oٽ�o�]�>��l?�y>�=�=p����]��7���r>�d�>�?��>��
>�mھW}�i��렿D�R����>	�?��t��9��e>�=�?��(>�������>��A|b�^�.�n�ﾝ�4�-?{�_��=k�:�d����T���볾�H'?�?�3���$)�rڊ>2"?���>٥�>K��?(�>�����C����?�U^?��N?��A?�<�>w�l=w����#������=�݈>�V>��5=�R�=���X�V�1T%�B�T=�n�=��e�����'9u�C����;��=Y�G>mۿ�CK��پ�	����<
��爾����'a��5���_������Qx���	'��V�4c�
���;�l�R��?�<�?.z���-������Ҕ��J���Z��>�q�.��j���U���*�����Y���d!�	�O�&i�%�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >XC�<-����뾭����ο@�����^?���>��/��o��>ޥ�>�X>�Hq>����螾u1�<��?7�-?��>Ŏr�1�ɿc���~¤<���?0�@��C?�r�"L�J��=a��>�?�^f>�궾��.��Ծ���>.ܩ?soZ?�I>��/��g�ݝd?<N˽�pP�o{$�oc�����v>;�ּ���>�-�>w*o���-�+�x��Ǆ=��>1됽o������il���d>��轋C5<�΄?Bt\�f�r�/��A���>.�T?�_�>�
�=@�,?�H�={Ͽ��\��$a?�1�?[��?��(?������>��ܾe|M?YA6?@�>l&�Y�t�R�=�)�z]��h���V����=���>B�>�,�R��loO��ƕ��k�=� �j�ƿ�+���"�b����=�Z��T���oKs<:lнKl��.Y����;�>���="�>�<�>�?>-�=>�?W?J�L?��>B�>o㌾v|ݽ��Ѿ�[��Ft�Z�S���l�JQu�n�����վl@������,��A�w��� =�|�=�6R�Z���3� �d�b�F�F�y�.?Uv$>)�ʾa�M��-<^pʾ\���Uل��᥽�-̾�1�"n�P͟?_�A?������V�j��R������W?GP����iꬾ ��=���m�=�$�>��=���� 3��~S�p0?�J?/z���ܐ���*>������=�l+?oZ?�cP<B�>�_%?8�*�rx⽎d[>�l3>��>�Z�>��>^���'�۽t?�yT?�����ń�>)��(�y��}b=I�>}�5������[>�9�<~�����_�tw��q��<>*W?ŝ�> D*�%��đ��-K��P=cgz?�?���>�2n?��B?�d<l���s�S��Q���[=�1Z?�*j?�X>x���&о����5?�c?4_N>�t���4�/�þ�QQ?<Un?�o?8����z��'��"Z�m=3?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������O_�=�=��ᨱ?u�?.RҾ� �<Q���zi����]��D{>jϢ��g�<�	߾RC9�����ݭ��	��W��>��@,������>j0c��,�[cͿ8�w�HV��W����Q?�Qx>ƪP�*�ӾTu}���w�&0B��s2�=�6��T�>4*>���������1{���:�۝�z�>ƺ�hJ�>vO�I����퟾��c<��>s��>Q��>�����㿾'�?M`��3�Ϳ���z7�H[??�?"o�?V�?虔:�{�G�t�앇�� F?Vfq?�2Y?8F�{`^�D�7���j?�F���S`���4�-CE�0�T>S3?SL�>��-�B_}=�&> �>k/>�+/�B�Ŀ4۶�i������?Ɖ�?�h�P��>|�?�t+?Ge��4���U����*��M�A1A?�2>�����!��+=�������
?}x0?v��j2�>�_?�a�Z�p���-�g�ƽ�ۡ>u�0�>d\�9D����(Xe���mAy����?N^�?d�?��� #�c6%?��>G����8ǾZ�<2��>�(�>�)N>�F_�,�u>Z���:��i	>���?�~�?'j?䕏�����W>�}?�H�>�?�f�=��>���=li��Wp)��">��=�h@��?�M?��>2/�=��8�$/��F��;R��$��C��χ>M�a?{L?�3c>ҙ��L5�l� ���ʽ�m0���!A�FG*���޽�^5>8a>>X�>T�D���Ҿ��?i�ݔؿ�l���x'��*4?f��>�?���t�t����X<_?f�>@8�{*��(���Q����?�G�?��?0�׾t�̼> �>_?�>�սC���x�����7>�B?L�mB��u�o���>���?�@�Ү?�i��	?���P��Ya~����7�L��=��7?�0�1�z>���>��=�nv�ݻ��W�s����>�B�?�{�?��> �l?��o�P�B���1=6M�>˜k?�s?3Ro���h�B>��? ������L��f?
�
@~u@_�^?*��տ��w��+ξ�D�=���=� ?>�Ԅ�
�|>�+�=U~.��T��|$>�O�>覒>��>��>R�>� >���H$�*s��I���zHD�F,�#8�@�|����[W�w��.g�t�S�v��.޽5%���洽
ힾ�4� ih>��3?D?Sz?�?��=�os>ʢ#�y�=	���g��u<?u�/?G�S?�?q��=ɋ< [�����v����W����>���='�>��m>�6�>�Q>�|�=���< '><��=X3>ijȼ����UT>��>���>��>�C<>��>Eϴ��1��j�h��
w�m̽/�?����R�J��1���9��զ���h�=Hb.?|>���?пf����2H?+���z)��+���>��0?�cW?�>#����T�,:>1����j�3`>�+ �}l���)��%Q>vl?~�f>u>-�3�Xd8���P��z���j|>�26?*궾gF9�@�u���H��bݾ}IM>�ľ>D�xk�k������ui�Д{=�w:?̈́?3���ⰾ��u�:C���QR>E;\>�U=pf�=ZM>�`c���ƽ�H��b.=A��=`�^>�(?u3>��F=�<�>�����d(��>uE>��,>@�6?'�?e!(��Q����g�oR)�L�j>���>|Bi>W�=k$M�͝�=��>��l>	�<��Խ�.�p�/���>U|���q���Ž���=~�S�y�>!��=�
��8����<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�p�>RJ��R�������u��&#=��>�7H?35��p�N�	[>�)v
??��P����ȿU�v�A�>��?x�?�m�0C���@����>���?�bY?'�i>#=۾
KZ�M��>B�@?]R?�"�>4�"�'��?+߶?��?}�{>�`�?�NR?�C�>!���KI����'م��k���j�<��[>��<Z�ʾu<f�:'��Д��W�p���,�>��6=�ջ>/k��KԾ�:��鬽�Jܾ�D��Kú>}+�>�T�>h�>2�?�h�>���>1��=}��=#���6��DK?�4�?k ��pv��<�8��&��ơ�>��?���=r�i��0�>~�]?
2?�Q_?+�u>v�羶���N������[K��)1>��?fl�>�5�=$ �>^eɾ�^��ۀ=Жy>M��=?2��V[��JJ���>��'?4�>kT�3�*?];?+�	>��J���W��Z��d`k��� ?� ?0KY?�?��? ���"~�[q���t��$e���0?�?#�?���>^������<�j>��ݽ�4 �)�?N�h?:��=�cO?�h?!.�>��F?�K�>UF�f���W�U>�>�>��!?n*���A�N&�:��۞?��?���>���*ս��ϼ��!���S�?}\?�S&?��Y�`�U¾��<0�+��]u����;��S��&>�>J���9�=׷>@��=L�l�,�4��"v<w��=�i�>�<�=��4�}Ɋ�1=,?��G��ۃ���=��r�FxD�o�>�IL>����^?il=�	�{�����x��B	U�� �?���?\k�?��:�h��$=?�?a	?�"�>�J���}޾g��Qw�X~x��w��>���>��l���D���ؙ���F��Y�Ž/��ƪ�>���>o�?{� ?G)Q>��> ��=�&�S��Z���]�s���7��-��)��џ�t�#�w	�C���Y�|�]��>Բ��-��>+�	?f>�	|>���>Mj��@�>��N>z^>�}�>Z>��6>v��=p�<xѽ�AR?�b��6�'�a������B?$d?(�>�qm�%u���:�@ ?4�?H"�?��t>��g�L�)��j?�x�>'���v	?��8=O௻�n�<�I��Oe����*�鼩r�>�׽T�:��K� 5d�;
?�6?����<˾gfս��[��͉=��?Ś-?�HU�*�[�w���F�o-c�D��=`�d�U�̾��#�܀����
�t�ד��j�k��=�d5?W˥? q&�YW�͆��{ow��i^��>j�?H�>��<�͔>��-���t� Ty�2\���L��[f6?���?�á>��8?��#?5�V?�I?V��>n{�>�AϾ$��>�����A>{�?�-?C�6?D�?�� ?N�.?M��=8xd��r�(>Ǿ��?cI�>R	?}ܶ>���>H���� ����<t� �i����_�"��=��==����b�9=�p>�]?tU�˦8�w���k>��7?_��>�[�>�1��:b�����<d]�>�
?�V�>����
er��3�[�>��?u+��=.�)>��=Ӏ���Ѻb��=��ü�(�=�E��f&;��<��=2ɔ='���iA�����:�0�;<K�<u�>7�?���>�C�>�@��0� �d��f�=�Y>GS>~>�Eپ�}���$��w�g��]y>�w�?�z�?�f=��=��=}���U�����H������<��??J#?(XT?`��?z�=?]j#?յ>+�iM���^�������?{!,?w��>���=�ʾ���3���?7[?�<a�����;)�7�¾��Խ}�>\/��/~�����D�й�����D~����?鿝?�A�0�6�)x������\���C?6!�>aX�>x�>t�)�4�g�3%��0;>���> R?���>-c?S�a?�^"?q�H>="J��:��4?���;�>T+J?^�t?wM�?�t?�A�>f��=���|�羟b�g�7�:ힽ�f���"=�7D>��>P7?ˍ>��=E{��,�QC�	�-;,��>7��>��>�N�>l�S>o@�|G?-��>V¾pV�<M�����
���v?���?f,?�{.=��h�E�'1��7�>o<�?_�?)!*?-�M��^�=D2ܼ)=���(q����><�>;��>G�=��Z=�" >�>�=�>�����s�7�5�T��^?�'G?8��=#ſ�Ar�sf��W��䌺;���WVd��Ŝ�� b�≕=�������T��*WU�#-��Ҍ���$��=!��q��I]�>ZȈ=��=Ī�=)n�<i�༃[�<M�B=��Q<��=A�W�&��<Q��S*��@�����7-TX<_�_=��W�ľ�z?TcI?�*?��E?o��>�&>/�e��>)��q3?+<><�e�j����J.�ߡ��B���Nؾ!�ؾ6e_��M����>WC%�-�>/J/>�s�=x%�<H�=au=��=&+y��V�<�*�=�A�=17�=���=��>�
>�6w?X�������4Q��Z罥�:?�8�>j{�=��ƾp@?~�>>�2������yb��-?���?�T�?>�??ti��d�>M���㎽�q�=I����=2>t��=u�2�U��>��J>���K��A����4�?��@��??�ዿϢϿ6a/>x8>�>=�R��1��7\�NV`�EY��� ?\c;���̾|�>H��=�*߾e�ž��-=��5>ݙf=�*��J\��W�=����8=��q=9Y�>ZD>�8�=�����=/�K=j��=�*N>S�w�f�7��#/�Zj3=��==�b>��&>���>��?D;0?�]d?�N�>�mm�C�ξ�}���$�>�D�=�#�>���=K<B>)��>1�7?2�D?��K?47�>�҈=Ӻ>�ʦ>�q,�}m�q���秾��<#��?�ʆ?�޸>�gJ<7B�G}�a3>�eĽ��?� 1?Q?���>�E�ֿ�l�|FN��\=�Em��=c�z�Fv�>��=;W&��I�=�׿>�=�>�)�>�!�> �>��`>��<!)�>*�=vI=䥱=+�����%>�[t�P2�=�YE�?$����=� �<	��=�����*��v��;�ݽ&��;�w��u�=�8�> >�O�>��=���8�->�i����L���=�X���B��1d�;]~�(/���7�MsA>�rY>���j��\�?9�Y>��A>��?�u?Wa!>H7���־Cp�� h���T��ǹ=7�>x>��8;��L`��=N�H2Ҿ���>�W�>�h�>Lk>�*)�$�B��:=�.޾�!5�^�>���WRV�����u�)]��.ʠ�p�j���b<��F?kr��i�=�|?AK?��?
��>��|�&T��b>杋��ZA<���da�%E��L;?��%?w~�>�d���jC�0t˾�1��%��>w�J��)P������0�����ն��2�>o���HоI*3�����K8��n�B�,�t���>P?nî?��`��l����O�`K�)��^c?��g?b�>>8?�l?j������K�=+[n?`��?�7�?T>o�&>.rܽ��>E�?	�?�?н�?���=�>A�8��'q=�lѾrE����=���>mW>���>^+�>"��>j꛽�P��g:���,I���z�=�kF>�%�>h�>a��>�FU=����e�=,vr>R��>SY�>!g�>m/�>�)�>�ܾ@�!�^/?���=�c>�tD?A�L>��j=Z��;{M���p<5�7�<De�����潖l>�Z�=-Z�<�+��'�>�P��$`�?z/�>Y)��8(?�v��1!��}<>G#>իƽ�4�>"H=>!�f>��_>=�>�h�=��E>0Sp>�6Ӿѐ>��`!�3C�φR�|�Ѿ�rz>ʜ����%���q��u`I�Q���ot��j�c2��#0=��C�<�F�?�M��U�k���)�^����?�K�>�6?k���7z><��>�Í>V�������ˍ��dᾷ�?���?N<c>��>��W?K�?H�1��3�xuZ��u�%(A��e��`�W፿������
������_?��x?�xA?sM�<�9z>��?��%�ӏ�4*�>�/�';�-B<=,�>")����`��Ӿ�þ7��IF>~�o?%�?0Y?�TV���=}R>�>?�d'?�]�?�?g�S?����:>+�H���u>���>�&?�?�x?S�>�_q>�E��!ǽ��_���n�pS�9v��g=���=�b�<Y�O=$���H�=�p�=zp\���,�dT����<f��;8B�<Xe�=9��=��>ڇ]?~�>��>��7?����8��(����.?��5=ւ�21��'���v��>��j?q�?��Y?>+c>�A�IFC��>^n�>�&>_�[>�O�>��:?E��{�=�Z>��>�=$(M�с�c�	�5w����<�t>h�>ǘ�>����Ii>S�f[u�^b>�j�!����U��`@�m#&���~�¬�>�tK?��?$��=>��˽a�`��`?ڒ4?�R?�sz?\>�]��S�:�WbL��K��>�-F=������ȡ�o7�4�<@c>�G��d顾�]>��	��ܾ��n��pH�		�73==����H=O���Ծ�v���="�>����	!����j���I?�
\=:{��#U�pF>�B�>�ݮ>20�v��@�2=��>��=��>B)?>�i��"��8G��F��È>[�E?��\?Z�?��:-t�gC��$ �Ej��V8���]?ѱ>��?��<> �=����Ŷ�ѿd�fIG��Y�>���>���zVG�hʠ��U��a�$��Њ>͑?��!>MF?��P?C�?��a?��+?nZ?���>]Z��󿾾''? 4�?��<=7��B�\���A��dK�Q�>�%?p�9�jj�>��?�[ ?��#?}tW?�u
?��	>L���vG�qz�>*ω>N�@m���>��H?�M�>�Y?��z?cf>Q)/�E����:a�>�WB>F",?~�(?Lj?�ܮ>�4�>�0��R�G�9�>4�H?�Ae?�ݐ?�?KN?��ռ���>���������>��?6
 ?ᤄ?U�i?<�>���<q���x�7.��н�^.<���;��>>s��=AKɼ���.}�1����^���Xҽ<a�|_^�p >_�@>Q�>��s>����1>f�þ3���zAA>I����5���׊���;��ж=+��>�Q?p��>C#���=H;�>z��>p����'?[?'�?B%}:��b�*�ھ��J�[�>��A?���=�jl��:��*mu���i=�m?^?d�X�~}����\?Z�j?�p�>,����ǃ�2���B?+ ?������>�m�?1]?��>6��+d�#����y_��߻��1�=���>Z�cwZ��xb>��?�i>�K�>H3�=B/c�&�c�rm��^�7?��?$w�?sz?�jz>N2]���a���͖��]?���>M���,?Уg����Y.��-���������F���6��K`Ѿa�1����:�).C><�?(�u?���?�Y?9���Y�<�Z� Yt�W�_��߾��	��_#�
�6�LD�a n�5��?��H����˻bkھNV��c�?��&?�:���	?������d$־]�D=~R��Dm�����>��	�]��Rj>b����*���fd��]!?2A�>�	�>a> ?f)N�i�����!<@����6��=F�>���>�q
?�s,>��Ǳл�虾dʮ�8�x>��c?"�I?;}m?��G62�ʌ���""��K/�F���v5D>
�>�|�>:�[��X�c|&���=�J�r�(���7��jj	��ʂ=��1?�|>�[�>�z�?��?�`� ���Wx�B�/�,�<���>��i?|�>���>5׽��"���?��}?:sS=�S�Yc���rl����kj^=(A�>D2?��8?y��>0l��� ��٭v��됿K�7��6�>B V?��i���� �>�$�?���=A/�<� >!a徴�S�|�x�'�ƾ�N>�� ?�ϻ�9�@>����`u���a��I��C�(?��?`]���\(�.l�>� "?��>�P�>K�?훙>k�ľz�ɻ	r?&�^?7J?{??�e�>��/=�3���dǽ�$�&=E=\Ņ>gmS>\tN=���=��9)Z��� �Y�]=R��=tż�f��v<C�����;�t�<>�0>�kۿ�TK�27پL��U&��
��#��������	��x���՚�6x���h�*���U�P0c�������k�3x�?",�?_���굉�B���c�������(�>�}r�s��嫾��V�����# ��d!�9)P�i�?�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >YC�<	-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾x1�<��?7�-?��>Ďr�1�ɿc���z¤<���?0�@�@?�%�J��F7c=�0�>
?�yC>A����j_��m��>�\�?	�?A�c=R�U��N%���d?$x<)�F��U���=h�=�:=����8eS>/C�>޽��4?��E׽��+>H��>3�<a���]�X=n<�=Y>s�Ͻ�f�5Մ?+{\��f���/��T��
U>��T?�*�>U:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�܅�=c6Ἴ���z���&V����=[��>f�>��,�ߋ���O�J��L��=�*�Vſ��,������B�.�o=�����"y�=x���q�@��T�$/��Hm=dK=ϊ�>G7�>���=��>�BY?N�X?�� ?-��>��7�"���E��A=���L���m�qv���0��� �����s��"����et(�_ =��=�6R�1���+� ���b���F��.?w$>��ʾ&�M�#�-<�oʾ����҄�=㥽�-̾�1�!"n�͟?C�A?������V�T���Z�?����W?�O�]���ꬾ���=������=V&�>���=���� 3�S��t/?0?h��������4>�j��{+=^h(?�~ ?�j<��>+�"?��&�i׹�4d>f1>�6�>p�>�>�W���ݽ� ?��R?���RD����>&��l x���2=�3>�F&������b>�G�<|���򙼮稽v8<1W?�~�>��+�0/ �9����3l�9s=�y?��	?@į>�Ho?�JD?��;�����1R��.��P=MZ?!gi?��>P�p�G�;Vq��]u4?��a?�_F>�6m� C�@0�!�l�?F�p?�?�����y�{����
�~?1?��v?s^�ws�����9�V�n=�>\�>���>��9��k�>�>?�#��G������vY4�"Þ?��@���?��;<��^��=�;?g\�>�O��>ƾ�z�������q=�"�>����ev�����Q,�b�8?נ�?���>�������~=dc���?E}?�E徝D=��KT�\��oL�=��Ͻ^��WV<;��6[$��	d�ē+�X�������)%�>.�@]�\����>C߾w�����	}�����¨޽��>1��>�ǰ�F쾍^Y��ꑿ]zr�� K�٫7����>c>�푽g�����{���:��������>���:��>A�S�����X���><<@ڒ>�C�>��>�2��R���	��?+���)οv����!�	�X?�q�?�t�?�W?0�J<��w�t7|�,b4�+�F?v]s?+�Y?˨&�~�[��1��j?�^���U`�u�4�eHE�?U>o"3?�C�>\�-���|=�>��>�d>�#/�H�Ŀ�ٶ�����t��?Չ�?`o����>1��?�s+?Di�	8���[����*�-��<A?�2>������!�_0=��ђ��
?e~0?�|��.�K�_?�a�D�p�Z�-���ƽ�ۡ>��0�vf\�fN�����Xe����@y����?;^�?N�?���� #�H6%?��>l���h8Ǿh�</��>k(�>�)N>+F_���u>����:�Oi	>���?�~�?Vj?ҕ������U>��}?�E�>G�?��=�^�>��=�4���x6���!>��=5D��W?8�M?���>��=8�y/�F�5@R�C�=�C����>��a?�TL?5L`>���2��� ���̽�3���弅6>�.'��oܽ[6>�>>0�>�|F�gԾ��?j�{�ؿ�l���v'��,4?ᰃ>s ?���t���3=_?Yh�>[7�a*���&���R�4��?�F�?��?�׾}�̼�>���>�<�>. սI���~����7>	�B?��)@��'�o�m�>^��?�@�Ѯ? i��	?���P��la~����7���=��7?N0���z>#��>^�=ov�ٻ��O�s����>�B�?�{�?6��>�l?��o�Q�B�<�1=HM�>��k?�s?�Uo��󾓲B>��?������
L��f?�
@zu@E�^?*Ͻٿ=ך�����B�վo�5>�f�<�>��"�#D>@��=]�=�qI��F�=z�>c��>�)�>��O>���>W�Y>����ă$�!����@��"+���l��o	����̾����M���x��?2�����S��̃�.I���ሾ�J�{�J>c�*?��9?�Sy?�z%?�8-<���>���A7�sо.�+����>'�?o�o?Ee?��=DA���a����BOV�|�K�9+�>$1>�.]>:�>{��>[+7=�t�<hZ=���>l�P>t�ٽT���>1���k>��>w�>�2>�C<>Ñ>Cϴ��1��h�h�w��̽-�?}���M�J��1���9�������h�=Nb.? |>���?пg����2H?!���s)���+���>~�0?�cW?-�>'����T�8:>[����j�Q`>�+ �~l���)��%Q>tl?��f>.u>�o3�n�7���O�������|>��5?�����}9���u��iH���ܾ�P>qK�>�eC�}�kޖ���~�[�i���y=��:?8v?�}��
۱���u�l��� R>JZZ>�=��=��N>7�\���Ž��F��(=���=t\>}??�,>=�=�y�>U:���.I����>�!<>P�*>D�=?��!?@t�����3�w�;%�J�t>���>w�}>�M>qxJ�pi�=���>�Ub>C�*����V2�9:��gV>~��lZ�z�W��[�=&���=ՙ�=����C��V=@�~?�~���㈿��0X���lD?3+?���=O�F<1�"�! ��H��h�?W�@�l�?�	���V���?�?�?&�����=#��>#׫>Zξ��L���?�Ž6Ƣ�>�	��%#�IS�?��?]�/��ɋ�Jl��1>�\%?S�ӾSi�>�o�=Y��m��0�u���#=���>�9H?sQ���O��
>��u
?�?�b�#����ȿ�}v����>s�?���? �m�qA��@@�ہ�>ơ�? gY?�wi>b۾�[Z�*��>Ϲ@?8R?p �>9�U�'���?߶?���?�rX>�ޑ?��f?|c�>�߃��d6�?��'���0#y=��༲��>��?>����}J�.��_��؂g����|�X>@2=�e�>��Ž�����1W=%M�����Q_���8�>vsP>��<>�.�>��?���>b��>��=�ۂ�Lɋ�ᱱ��cJ?~��?77��}`�f=��4�v�־	�>k�>&��=	�C��x�>ih?+�u?F�?K��=l��ؐ���տ�\m��[Ҿ<���>���>�3?���>T��>5��{f��� o>��>��C���Ծ�R{�������>_�+?	��>y�=c>$?�B?嫘=��\g|�Z����i� j$?�O5?&_e?��<?�6?U#Z��_�HK���G�����6<,?���?��?W#�>�����򜿥�>y7@����=Vl? P|?6]>��c?��V?���>�zA?���>����=�C��>[�H>п!?���j}A���%�����?�?��>C���b�ֽ	y�>�_���?.�[?��%?��ol`��&¾e��<�\����W�;CY��4>��>����ӳ=��>^��=�nl��s6��Hh<�Խ=�$�>��=@-7�Iq��/=,?��G��ۃ���=t�r�'xD���>JL>�����^?�l=��{�����x��	U�� �?���?Zk�?���1�h��$=?�?K	?U"�>�J���}޾;���Pw��}x��w���>���>0�l���M���ۙ���F��:�Ž]+��N�>���>�?ص?
2d>���>ȴ���u+��I�Qs���Y��Y���-�d)����`딾�����.���qh���#�>�a�j�>@�	?dob>�΀>�9�>(;j&{>_<>;�v>ۭ>'ja>!�9>�t�=Ap:�����Q?������'����gέ��]B?�8d?P��>�vp��:��Z����?�'�?��?�Fw>7h��e*�,?�@�>j-��#�	?�fA=�񻇘~<z�����������v�>3�ڽݏ9�L�X�b��k
?�5?�����5;�׽����z�=b��?� ?�FO�g�]���~�y8U��Z�t>%�ľ�Hq��+%�-��	^��괃�c��;�'��v>�0?��?�� �;Z*�z����\��TT��R�>0m?��>��>�{�>l�4���E��'��k�=�L�?*�?�>�>t$K?G ?�o3?]R?�1�>���>����?�=n�ܽ��>7��>(�#?P7?�� ?�Q�>�|(?�M>�þ�8׾����>��%?^c??h"?��?����U)���W����B`���Խ��=�d�ۃ)��kH����=Ч�>��?��z�6�yS���Er>2�6?�7�>�5�>߷w��w����<:��>��>�ۍ>��龤nm�[��׬�>���?Bv�/�=�3>/ʮ=���sP���u�=��4��a�=�7ȼ��Ż�`=��=hW�=�>�o�<�7[<R��<���<u�>2�?���>�C�>�@��)� �Z��6f�=�Y>;S>s>�Eپ�}���$��q�g��]y>�w�?�z�?�f=��=���=}���U�����E������<�?;J#?'XT?[��?r�=?Zj#?ѵ>
+�jM���^�������?t!,?��>�����ʾ��͉3�ٝ?_[?�<a����;)�ڐ¾��Խ�>�[/�a/~����=D�����`��6��?꿝?�A�]�6��x�տ���[��m�C?"�>&Y�>��>H�)�u�g�j%��1;>݊�>[R?>4�>PqO?{gy?9�Y?�R>.P8��<��i)��]�n���>g�>?O�?�ڎ?&�x?#{�>�*>5%�W&������o�����T=]�^>Ⳕ>�J�>Ȉ�>��=�����<��H�A��D�=�b>�3�>��>��>9�w>;¡<��G?���>�\��R���ɤ�9���ܡ:��u?���?1w+?=�=�|�K�E����T�>�]�?���?OL*?DS����=X׼nѶ�~�q����>D��>�!�>C�=��E=�>��>��>j(�jI�m8�AaK�	?xF?ԃ�=��ÿ�tv�gI��!���)�;�|w�B�V�Иd��)N��#�=�>���s/������e��{��ڟx��h��'���&Fj�I��>�:�=�,�=#��=@��<&�ür��<J�p=�n<�J=��n�8Ѭ�;{��{����퐽��以��<W�}=b���Y��v�q?�wK? 01?\EG?_Sz>�CT>����ۇ@>L�ｾr?�x2>�N��������̍�&�N�ؤ�@�ϾϦM��Ě���=Ĕ�pŽ=��C>���=z�<��=o:�=�
>�'�/�<q�=�~�=�A�=��">;#>��>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?~�>>�2������yb��-?���?�T�?>�??ti��d�>M���㎽�q�=L����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�
8>ű>�R�RS1�*�[��6b�A�Y��A!?7R;�U̾�'�>&p�={�޾\'ƾI10=^6>�'e=�h�e\����=�?|�vG:=�sm=�%�>�mD>ue�=]а���=�[I=�g�=�O>�圻�'8���-���2=ެ�=G�b>u�&> Y�>�i?eQ0?��d?Ow�>��j�@˾ O���_�>���=�S�>߉=�QA>DR�>�7?�D?i�L?�>�p=�M�>ڙ�>5,�}�l�e��뉥��м<:*�?���?us�>�g<�b;��D�>���ƽ��?�"2?��?�i�>e�j�޿��P���.���������=:�F���=�(t=��=
�u=jǎ>���>�J�>�'�>dx>?4)>���>��=�e�=���=�[E��6�=��7�<	�ļ_d����e�U�ս�s�<�g�Q�����G=i�=��@{��o��=���>�&>��>�֖=A���,N/>�͖���L�v��=w=���$B��.d�%?~�E/�hh6���B>�<X>�����1��?�?��Y>e�?>b��?�Bu?��>�#���վLM��sUe��]S����=��>M�<� |;�W`�&�M�z`Ҿ���>/�>��>ʭl>d,��)?�Nw=���]5���>*o����q7��>q�P=��L���3i� Ժ�D?�C�����=�~?�I?�ޏ?���>�����ؾ,(0>�i��ig=B�xq�D��S�?�'?���>�*�f�D�� ̾Cg����>�}I��P�$���;�0��ظ����>�"����о�73��t��}��g�B�<�r����>�O?|�?�a��_��h�O����o����c?ǒg?�_�>�5?4D?�!�����JO��8y�=A�n?ۡ�?�C�?�Y>�^E>�q��K1�>~?�Й?Ͱ�?n�p?����)�=?ޗ���=�(��ɼ�"�>�M>��4=F�?���>Sз>�-���v���7o����F��=Z��>��>'
`>t!D<�l�=צ>�ѭ>�%�>��>��=1�>��8>��� �E�E~S?�^>��[���M?�	>��N��U�M���C��)�W�>��;�b�1��>r�^��\��Z���>�쭿��a?@�b=��4�@?�9Ƚ��S>���>]Ӣ>17���:>���y=t��>���>�t�=��>iu>SӾ �>����a!�iHC�ƅR�<�ѾbEz>�����h%�q��x�����I��⵾���'j��5���$=�yn�<C�?�M����k��(*������?�7�>?6?;\��T���D�>���>�q�>�$������<э�tI�W!�?���?�<c>��>8�W?q�?��1�<3�ntZ���u��(A�e���`�$፿����F�
�_����_?��x?xA? F�<�9z>Ȣ�?\�%�Yӏ��(�>/�P&;��C<=�*�>�(��O�`��Ӿ4�þ�8�IF>��o?;%�?�X?�RV��<�<5QB>�a7?g{??��q?�?!?�s@?��B��=�>��X;V��>*F?�%?.+?�r�>�^>��Q>.b�Wd�B�,��'d�h=��Z�Z���ń=?aP=���<}	��{�9=�'j=iMɼ�m���A�H�Puf<-V={i�=��)>_&�>M�]?E�>���>:�7?�Y7����p�-?2=�����.���㡾�=�G�>�j?«?�Y?��_>��A�h�D���>SP�>��*>ğ^>�*�>-]�
0F��C�=pz>��>�ˢ=�M������	�����O�<�Y">���>�R}>�����'>�W���y��e>�T��G��CT�tG�܇1�\bu���>�K?q�?���= *龀P����e�g�(?�;?�NM?Y�?[a�=j�ھ�9�N�J�C!����>i+�<I���l�������}:�`��9}Rs>Ϭ��M��[^>*�
��ܾ�n���H�iF��pN=���>?=�0�;�Ծa@|����=l�>̾�� ��▿8��y�I?�Fc=������V��I��j�>*��>	��>�+��Yn��W@�`����=`�>L;<>'X��x��F������>I�A?_'1?�:o?*����;{���C�<����-���?�|�>5��>1�=��/>�����-�F�q�� 2����>���>2��O<�<,c��r��G��X�>R�?�{�>���>.�)?��+?�r?D�C?e�>x��>{mѽF���9/&?��?˔�,�Ͻ�6�3O�S*^��ī>PU6?�����&>TK?b� ?y?Z]?��>���=:���Y(��9�>�l�>��8�h:���´>$5?q32>�A?���?��>A�0��_Ѿ0�f=ױ�>GZ�>�.?�K ?�T?vD�>���>N�njּ�l�>|?.��?r�?_Dh>��>��;>H��>6�!���q>i�>�?mD]?�ف?�9F?�G�>d�<a����ν�1�$�̽	�h=�Ұ=��>>> �=��k�Ja�<����P�./�=-�|;:Q���?>h2�=�b�>�s>�����0>��ľoC����@>؛��\���݊��w:�c·=x�>2 ?䲕>1Z#��Ò=b��>�1�> ���-(?d�?�? �';ǔb���ھީK��	�>r B?I��=�l�8����u�G�g=3�m?x�^?�W����0pb?o^?���>><��}�� zk����L?�9?k�?�䑮>�~?�r?:��>,�Y��m��e���b�V)g�o]�=c �>O^�t�d��j�>Q�7?�R�>��[>��=�Ӿ��u� N��q�?zR�?7��?���?�,>��l�i߿Ҳ�!����W?�2�>ړ���9!?p!�����h�]�]���:�徫�Ǿ�U���o��8C��a:��kc�������=i?7�m?�t?4�\?a��oU��zY�A<���Vd��V �4�H;�!�I�(�@��Lc��6�u����N�;ί��^�R�?�9%?otӾ`?��u�[�+�s�U��>�*f��iH���M�>��>6�j���n>��#�W���&�~�-�"?ݚ�>�z?��%?��[�H�0�1����*�[S+�a�>a��>�=_>���>����`���W����i<y�َ$�'C�>�a?��7?-�c?�����4�ay��"'�n�����ʾ��=>�gW>j�3>�4�����i��� =���o���?j��;�iϳ<R.?� %>��>��?��>���ø���;m���$����;��>DOy?]��>kI>
�M���.�U9�>�X{?�A�>�Vؽ�.��aHI���a�
9]>)8�>���>��=?Ȋ?~���i��倿^����,�<�>�?�?�^���I���8�>J�?��U>)5��}�j>� ����4�'��4���`>�D�>k�=�M�>biy<�������ľH�(?��?�����*%�b}�>=9"?�@�>�?�>��|?:��>c��&}޼I�?a?R�J?��;?ņ�>\$B=j��`½�,� ��=�Ƀ>��Y>�Օ=f�=J�Y�b�����7=Ov�=6��c����֑�����Y��;�(=�-:>�eۿpkK� �ؾy)�̍򾎩	�����]��`���&
�5���=\��}�y������)��
V��ea�e���}�k��5�?���?{����1�������������1�>�u��?��O��CD�nB��t�*B���*!�\�P��]i���e�P�'?�����ǿ򰡿�:ܾ3! ?�A ?7�y?��5�"���8�� >(C�<)-����뾭����ο=�����^?���>��/��n��>ޥ�>�X>�Hq>����螾u1�<��?6�-?��>Ďr�0�ɿb����¤<���?/�@u>?Sd���Ѿ���=�w?��?�o>F���%�����e�>��?X��?dE=nN��#�;��j?v����M�qb��v�=:��=�̃=D�+��t>�N�>Fq�ד!�<����>�)�>�(�8��{X���=f�K>#�����5Մ?*{\��f���/��T��	U>��T?�*�>H:�=��,?X7H�a}Ͽ�\��*a?�0�?���?$�(?7ۿ��ؚ>��ܾ��M?aD6?���>�d&��t�ۅ�=g6�;���x���&V�{��=[��>c�>Â,������O��I��V��=[ �.���TV0���ྻBL=Z�=���;�y=E+�>�罋��91��t=��=�	�<�hL>��? S>��9>!sN?�_V?��>�>51��E���r� �u4h�� 9�
w`�kB���l���b�8�ھ[��D��J�+�s'�o���!"=���=HR�1����� �*�b� �F�A�.?%>L˾i�M��i(<  ʾF|�����1���̾�1��n�Rş?�A?��W�V������I��ϰW?c���S���k��=�Ҭ���=��>���=+���3��LS�0?c{?=ҿ�aݐ���,>����u=��)?Y��>��I<�[�>g)$?��.���ܽ��]>w1>K٢>�>�>`î�f�ݽR^?�S?�� �S��}Ώ>$�����{�9/_=;>�x3���ۼkdZ>`�<�-��mQM��鐽9]�<��V?���>�j*�&�!��f��զY�¹!=��x?b ?���>�.n?:�A?+�;���NST�����-=�Z?Bk?�<> �u��˾K�v�4?+�a?=�M>��[�<���U,�����=�?6n?�~?K�ӻ�py�3�����{4?��v?�r^�|s�����I�V��=�>�\�>2��>��9��k�>�>?�#��G��ế�HY4�%Þ?��@���?y�;<�����=|;?K\�>��O��>ƾ z��T���r�q=�"�>댧�Rev�����Q,�s�8?Ѡ�?D��>�������a�=����m6�?f��?nP����g���G�zj�O�>�C�T w�J�K>�rϾH=�l�W���������I����>w�@������>��3�������ѿ������5��=�� ?��>}΄��+�xR����z���h��B��U�e��>�� >�9���;���y|�~7��ٵ���>����M�>q^�s,���������<�P�>���>e�>�꼽������?O4��/Ϳ������g�U?��?���? � ?��q<ދ~�Z��6p,<_�G?Vp?>?\?V��gW��T��j?�㧾sp`��5�لE��P>	&2?}��>R-�ą=�>�;�>�
>��/��eĿ�&��B����'�?���?���}��>g��?�T*?����󙿬Ш�*��j��
�@?��4>����)� �[�<�����
?�0?���E��Z�_?�a�M�p���-�j�ƽpۡ>6�0� f\��L��
���Xe����@y����?I^�?^�?��� #�^6%?�>R����8Ǿ��<Ѐ�>�(�>�)N>NH_���u>����:��h	>���?�~�?Vj?���������U>�}?�,�>��?`8�=�K�>�V�=m����/�uK#>g�=�M?�?&�M?()�>�=o�8�v/�VF�#=R���R�C�%��>6�a?�L?�>b>�츽� 2�e!�Xtͽ�o1�#꼃^@��,��e߽�i5>s>>]> %E�#Ӿ��?&e���ؿ�m��݄'��)4?Y��>��?/����t��5�S5_?�f�>�<��*�� )��Qf� ��?iF�?j�?-�׾�#̼��>E�>�A�>]�ԽBܟ��~��a�7>��B?�?��M�o���>?��?��@QҮ?� i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?lQo���i�B>��?"������L��f?�
@u@a�^?*�ֿh���}��a���v>̏
>��>���G~�=2y=W�=6�<1�=�*�>G˰>j��>�o>�_�>�*)>uȂ�j"�4���'w��C�_��5A�<��������Ͻ�F�������m)��OY ����\;Z�z����	>kK?�oL?P�n?#�?�O��yV>p���mм�(H��T=<�>�(?$QK?*?���=%���v�b�;�� ٣�����S�>|Y1>��>6��>|ة>��<��I>� F>:+�>���=m�=�A<�C{=��m>W֚>��>�>!C<>�>)ϴ��1��\�h�@
w�O̽�?����V�J��1���9��X����j�=(b.?t|>����>пV����2H?(���x)��+���>o�0?�cW?��>�����T��9>�����j��`>�+ �a~l��)��%Q>�l?{�f>^u>Ö3��,8���P����Ki|>�5?Dʶ��o9�V�u�p�H�w@ݾZ5N>M�>�B�C=��Ԗ�1�i���z=��:?kS?�!��,�����u��흾��Q>�\>�8=L��=��M>��a���ƽ��G���-=�=�^>q�?�.>�D�=V�>����Q�I����>�k8>�">GO>?gf$?F'����]�}��&�u+t>g�>l$�>v�=�8J����=څ�>2O`>�U���u�[C� s<���R>f�x�*4\��l��ׂ=)������=��=/���6;�8�&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�l�>�Y��X�������u��B#=��>�8H?�N���TO���=�hv
?�?�j�`���S�ȿ�v�	��>��?��?��m��>��,@�A�>���?�dY?h~i>�^۾�]Z�U��>��@?�R?��>0���'���?'ܶ?ì�?yfR>TV�?��e?2'�>B�����1�`�y`���P7=�A=���>iF<>��о;�H�ً�eԄ���j�����MZ>N�)=)�>�� �f��]/8=�V���谾�Q��>��>�P�>4�;>���>�{?@��>R6�>�@=�����x������N�G?��?w�
�,X��3�=�5ν/Ӿ��=��?QK>X���>��??(߄?���?���=��辪Í���r����<Im=s�>�"�>>X�?�˾T�羦.d<�?݄�ǂ���8�9�A�ȥ�>�w%?�* ?Sĝ�w	%?>?�1�<(=���GU������N���>�I�>�_=?rA?8�?�G�++s�O1����������?�S�?Y�>�U�>�%�����E&�<Q�g�ׁ�=Kv?�fI?z''�-_E?��J?���>K�%?�¾>)�ݾ�X=���_>7�t>4�$?�S)�%WX��4��P��N?G>?��s>R]+��8*���<rM"�I��?0�b?��?ؽ�p&=�ę��.�<o�����=��#=�=��k>�vH>��H���O=Q�*>շ�:�Մ��;�֏/=}��<@��>Z?b=����N�;0=,?��G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>$�l���K���ڙ���F��_�Ž��޽;�>#��>�|?Aw?+�>��>W����3������Eq[������!�z�fu����������ֽ�V���M��2��>|��*�>�?�n>L2�>Qn�>P2�����>{cw>�h�>&4�>��>k�P>�u6>�HɼС��rKR?����S�'���辍����0B?od?�>�^i�������z?1��?�r�?�Qv>s{h�>(+��l?�(�>���/k
? :=|����<�D�����,���:���>�R׽�:�\M��gf��d
?).?@��[|̾+׽�[w��y�=|�?��%?p#6�k.a�?�{�O�a.g��7q>�
��g��A���h��¨��I�b�O3��L� ��f>�]*?�v�?,�*��T&�G��b��.=��6a>��>�ř>wq�>��>�/&�{�J�R_p��L��
���?��?���>�5>?�.?#�>?�a?�-�>g�>�@�Q=>c����@�>�c�>D�?S�/?x).?���>J$?�}>b��?���⾩�?4?X2?-�	?A�?��.�|Խc���A��� �����,=1A����1�=�>������h>��?��}9����/1k>�w6?�
�>�>@L��M9���=Wk�>�,?���>��W�r��z���>Bǁ?g6��0 =�.>A6�=���u0�GW�=����_��=�\^���2���%<���=Q#�=\%��⳺s��:���;H�</u�>h�?���>�A�>6A��g� �q��
h�=zY>�S>#>�Eپ~���$����g�<Zy>4w�?�z�?=�f=j�=.��=1}��$V�����l���=��<ˣ?�I#?�WT?���?��=?j#?Y�> *�_M���^����n�?|!,?H��>�����ʾ�񨿖�3�ϝ?[?�<a�ʸ�V;)��¾��ԽJ�>�[/�T/~�����D����������0��?Ŀ�?9A��6��x辨����[��S�C?�!�>!Y�>��>-�)�F�g�Q%��1;>̊�><R?�>r�P?�u?�V?}VW>��:��������+<P5>��8?$�?�Ҏ?9"y?0��>-�>\�-�oS��������ֽ`z���!=�8b>��>?��>x��>mZ�=h͛�~ ��5S���=�t>��>�o�>��> 1z>��;��G?3�>ൿ���s���S���#�;��+u?nj�?wT+?�W=�v���E�s������>?J�?��?�*?��T���=@ۼ8���q�Ϗ�>qO�>��>��=#D=�d>���>;w�>V���H�/o8���K�k�? 6F?��=��ÿ?�s��6Y������r���ꂾH�d��W��n6��6F=ݾ��7�"�����%=�g/���Ɇ��@��� ��@l~��� ?��h=$��=9�=��hx�����<$ �=��<{=s){��*K<;�"���z<�ǌ�+��<��;0V:=ט�;�`˾ҁ}?x.I?Ԕ+?t�C?V�y>�>�u4��]�>�Ђ��3?�U>�
Q��c��BF;�����L���9�ؾ`�׾u�c��̟���>I,I���>e:3>�-�=l^�<��=��r=���=w�M��=�=S%�=�h�=8��=��>@S>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>
{^>cz3>�#[���$�t
��3��1����>�g@��:Ӿ�^�>^3=�C�����ps�=W>�l�=`�s[h�,k�=[�ɽv>O=��=��>�Z�>!>�h��\�[=z�=�Ҙ=E2>sr��+��iD����H=���=��>L7>'��>��?�L0?jId?���>Im�ͥξ�{����>	��=iB�>:��=�B>�>�7?�D?��K?�N�>�̇=�ֺ>���>�,�.hm�������Cӱ<��?W��?:~�>�#M<U�@��v�e>��$ƽ%�?�W1?�6?���>���-޿�*��%��<	��=��=��޽p= =�a;����*h�L�+>�ۭ>��>=͸>^-�>�=d>�K>C��>�T�=�Ի �R=3>4�T�]<�����=��=^�=���I�=�u�=PS��F��T���`y>��;�:��=���>,3>Щ�>\��=E��j?/>����6�L���=�?���%B��4d�bF~�K/��\6���B>�:X>����d2���?:�Y>�?>���?�@u?d�>�=���վ�Q���Me��QS�K��=��>��<�Cq;�X`�F�M��ҾHM�>Y�>�T�>6h>��(�ceA��FL=�)ܾ�3�T��>"��>�f��p�RVr�?ࣿ�����f��U;�E?�V����=Sy?�\M?"f�?�M�>�Æ�oW�9>)>�F�s<��.iy��i���?S'+?���>B?���CI��!̾]~��÷>��I�� P�����´0���*÷�x��>�誾X�оX,3��l��V��G�B�W�r���>7�O?&�?��a��X���bO����
4���s?!xg?�"�>U=?ON?@/�� x��a���Ҹ=�n?��?~9�?�>��>Jm����>1�?`�?�j�?�Zz?��p���>�������=y�;�zH�=�>��=��6>��?aK�>t�>[o���?�İϾ�_���VS��謁�]�=/4�>���>(G>��=�f>]O	>�F>g��>U"�>��k>�jM>w>�e龘�0��.*?�{>�(��>?�>U#> �>/�\��+��at�Kw<l��=��6�~�=��=���ݡ�K��>���*�f?[`d=�\���>:����[�=��>N!N>��\�7�>���>�X�>k�w>UH?�B>�p>o�i>�	Ӿ��>ڦ�PZ!��8C���R���Ѿ0z>�Ĝ���$��������o[I��������i��;���=��w�<�?�?V���A�k��*�������?:H�>�.6?%@��>0���k>�=�>z�>m��哕��ٍ�;A�\�?���?�<c>��>��W?+�?l�1��3�;tZ�K�u�')A��e�R�`�፿Ŝ��/�
������_?�x?�xA?)1�<48z>���?�%�=я��*�>�/��%;�KH<=+�>�)����`�߫Ӿa�þ�;�uCF>
�o?w%�?�W?�RV��`�;���=_�<?�>?#}?�c-?JIU?ƽ�{�>��=���>���>�(?� ?
C?(��>D�?>�f��V����#�o���ҽ��ġ"<�o>��=E�A=w��<�P�<oU��ֆ���LE��A��N��⼝�w=6�>���=���> (]?A��>�Ԇ>u�8?{M��@6�^��R6,?�y-=�5��k������g?>ɥi?�W�?h�Y?�([>oB�5�D�X2!>���>'>Z]]>p�>���'�E����=�M>b>��=NWV�G����b�cq��G��<� >`��>��>^<���f&>�ȟ�(�u�� f>^�X����WU��kE�f�1���z�!V�>�hL?��?؈�=�������e�?`'?s�;?��L?��?z��=�$׾��8�0�J��?��{�>.��<�������]����U9�C;�Dv>	6���󠾦+b>����ݾ�on�� J����{pN=ur���Q=Ӳ���վ�]�5��=<
>���.� ����������I?d�i=\1��,�T��A����>|��>��>�99�Lv���@�+E��ٙ=�>8�;>3ꑼ���F)G�x�/i�>��G?�i7?a�m?�2�����.Q�Fn��ui_�77����>5��>�%?�z�=Y�#>����T��gs���O����>`.�>]����C�O�𵨾=�<����?�y�>(��>q�(?�3?�=�?.�/?���>�x�>4���w����%?5X�?&(!=�����c�.!E���_���>��7?�0"�V�y>�?�/? J+?҉\?���>-��=���a�<�>��>t��>΍2�W������>IM?�\>>a<?!}?�I�>mc#�ڗ����?=�"�>�}�>>�?K$%?t?�-�>��>�B���a��6Y ?�`?N�q?��?$��>^�L?�Vh�B�/���=�a�=Ú�>���>��;?!ϕ?�(?ś<��=���Kٷ�Љ����a�d7�0	��v�?>�u(�-?"��/I���=��=�<׹��L1��DŽlg >:W��1�>+�r>�T��s�5>� ��:p���C>F�м)����L����<�2�=м~>�U?Ӌ�>4T����=���>iO�>.g�%!'?��?B�?�<:u�b���ھa�F���>�A?�h�=�l�����?u���t=�7n?X�]?J�^��j��^4a?��]?=c�dx8�\�ž7�~�|]�rN?��	?3�_��k�>9}?wQn?q��>��R��>j�����nwf�@�m���=�f�>���]��I�>[�/?�ɼ>�CS>]a�=��Ѿ*�r�O���a�?]�?��??�.>�gl��}�<*��M����%^?
��>�����"?�B0�^�Ͼ5R��^�����ݾB����Z���������������Aeڽ�E�=�?�0t?ָr?/�`?� ���e��^�2���W�j/��Q�	F�k�D�i�B�/�n�¯�����<b���/8=�����^���?�@?����4��>$s��?{Ǿ�j����> Q��f��<v�>S�K�D�j=l{v>u���}~1�p7g��-?�d�>>?0GY?�S@�GSH���$��;Q�����>�WY>g�>���>�}����V�����Q�о[hG�'�5�*E�>�pb?�M5?kEZ?��8�k>�����8���X�W+���>>�>>��Z>B���.��f� ���?��){�y���&葾��
��*��cC?Ԡ>�9>�֋?10�>���Êվ��U�H"���=��>��n?�?e�>��U��D�/s?Ç�?k��>��v�jy�)jU��uu�%>�u�>�>�>Z��>�&#?�7���-_�#H��wK����I���>s�g?KB�������'>� x?��z=�x=h6>�:�����#>��� �k8���p?�z��/�>]}�������J���H�(�&?]�?�ە���x��>�%?O��>�E�>C4�?=�>�Ͼlc��ǔ?�b?x�G?+�??��>A =�M���Ž�$�V.�=J�>e@>o�=�C�=V�뽫�L��8���_=���=�Tļ�N��@��<��.��w�;�I����;>�ۿ�K���پt�������	�~��	X��lӉ�&w�&���Uĝ�ɼ�����x�@��W���f������b����?���?KC��A�������O������W�>�,s���r�֣���^������ݾh���{!��lQ�Ii�8Fe�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >[C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾u1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@��6?�C�������=3�?3� ?���>����@�N�
���&i�>��?Ձ?f�;=>�J���ϼ%pg?�e$��"Y�����@F<��8���=��>�S�>[9�>�{(�|���Iؽ�>k�j>�|P��t����
�5<dV>��2��R>5Մ?,{\��f���/��T��U>��T?�*�>V:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�ޅ�=q6Ἱ���z���&V���=[��>c�>��,������O��I��V��=d��ؐÿ>A������=�	�mѽ{�+��-��u>���&=����bž{�׼�J=>�*>Hd>6z�>h�Q?�q?��?�bn>.Ei�Y_����н8���K�y��)Pn�Ȝ�����E��p��":�%�)��@��c=��X�= 0R�􍐿�� ��b��F���.?8m$>�˾��M��0<�jʾ�ા>��=ܥ��9̾=�1�|n��?<�A?^􅿁�V����gh�㋹���W?�+�|��;款r��=�����=�7�>.��=����3���S�J]0?�j?����q����(>w'�ą	=$�+?�K?�0<�L�>�h%?��*�ԛ轚\>��3>���>�A�>>�ˮ���ڽ?8T?j���%n����>~�����x���e=�]>p�4��ݼ��]>n�<m񋾔J����Q�<�W?C�>�K&�u�#��h��̓~��0=A�y?��?��>�ah?
�H?��	��v��2ZV�����)="�^?�h?�p>��r��̾'����2?
�_?hO>3b�D��/���:?��k?̬?�2�J�x�/K���U���2?��v?�r^��s�����c�V�y>�>i]�>w��>f�9�Sj�>.�>?
#�nG��R���fY4��?��@Q��?,�;<F����=l;?'[�>��O��?ƾ�{��ـ����q=_#�>}���nev�����Q,�;�8?���?���>7���������=�]��P��?�"�?���>	�Z��L�^�Um�p\$>xN�=�Ľ��K>�)��1)�Ս�X���E������>��@P����>A�O�N\��ɿ�Xu����c�����>�Q�>�ת�����o�W����]F�)Q@�O��,J�>V�>ꮔ���(�{��m;��۞��>��?�>�S�'*��ǚ����5<<�>���>h��>�)���彾fÙ?vd��!?οS��������X?=g�?n�?pq?�9<H�v�I�{��[�H+G?&�s?@Z?�+%�`7]�J�7�b�j?D���M`�$�4��JE���T>3?LO�>�-�j-}=v>K��>42>$/�׍Ŀ;ܶ�������? ��?�h�A��>Y}�?�p+?�d�.5���U���*�x�;��0A?��1>҄��-�!�@(=�5Ȓ��
?�w0?Հ��)�Z�_?&�a�L�p���-�S�ƽ�ۡ>��0��e\�kM��%���Xe����@y����?I^�?g�?���� #�a6%?�>c����8Ǿ��<���>�(�>�)N>�H_���u>����:�	i	>���?�~�?Rj?���������U>�}?l»>�ƃ?���=K+�>2Ȭ=v�ϾDI��C>�=oz���t�>��O?�'�>�d=�=�G�&�DF�o�\�m��=�n��>_�T?I?4">�����s��)�k�����c�L!/���=������O>��R>S�>�#F��-����?Hp�7�ؿj��(p'��54?*��>�?��v�t�����;_?Hz�>�6� ,���%���B�a��?�G�?=�?��׾�R̼�>;�>�I�>5�Խ����[�����7>1�B?T��D��q�o�{�>���?	�@�ծ?ii��	?���P��Sa~����7�s��=��7?�0��z>���>��=�nv�ݻ��W�s����>�B�?�{�?��>!�l?��o�R�B�n�1=7M�>Ϝk?�s?�Po���i�B>��?#������L��f?�
@u@`�^?)��ؿ�}���� ���޾'�C>��=�Y>E����*�=��=O�6>/�D����P��>:W�>}Z�>.@>�5�>�c�>���8$�%�����Ke3����e5��{��B���+m��{�� _��YJ��Qq�B���ۂ�,�ȾaJe�o>�={�>P�E?tD?q�l?s�?@j�<S�V>�)	��1=JK���<�#D>�!?,+Q?��,?��>H�q�-a����	����j��c��>�X>L�>�$�>���>��=)��=g">Q-�>�$<>gx�<�[ý�����r>%p�>��>gI�>�C<>�>1ϴ��1��]�h��w��̽(�?]���|�J��1��:9�������f�=?b.?	|>���?пU����2H?���m)���+��>>�0?�cW?�>����T��9> ���j��`>!+ ��~l�}�)�\%Q>	l?�Mi>qy>�3��Z6�=AP�����s>�A6?	����C��qt��UE�p�۾�B>%Y�>�y0���}{���~�|�h�|�z=�8?r�?Wᦽ�@��jx�?��!U><�`>��=iϬ=�iQ>:&=�Q»��D���:=�S�=�MP>'9?�?+>�=�(�>�,��M�O�>��?>��,>:�>?�O$?�e�F ���N���*���x>��>�C>��>��I��7�=��>��a>�<
��j��Q���;��GW>A|���\���t�u=�ܙ��2�=Ra�=�����;>�o}&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿvh�>zw�eZ�������u��#=ݨ�>�8H?VV����O�d>�(w
?�?_�쩤���ȿ4|v�H��>I�?���?2�m��A���@����>��?�gY?�oi>�g۾5`Z����>̻@?�R?*�>�9���'�m�?�޶?���?�J>�~�?\�r?O��>y��H00�����̋�F�=t�:qv�>jX>����z�F��l��s3���j�!��W^`>�H$=\Ǹ>�l�Tһ����=,����e���u�E�>)Or> �I>�(�>Y� ?��>�K�>��=����R��� ��f<C?� �?��ξ�X���=%~�����=��-?�FX>������A��@x?T��?��?���=��Ҿm+�����_3���<�5W>kn�>Z�?RA�>O�)?ҵ�%���%�=���>]��)��7P������>�=(?�>��ƽ�B)?��N?��>y\��,m�= ����[��1�>H�>7�O?��?�L?�쾑�h�ֺ��(f���k�a�?�8~?�
?ގ�>��H����*�>����Ҽ�Dc?��[?%;����'?_�|?QG�>�d6?Mn]>��"��dr����>~X$=�� ?B���>�LB ������	?,�?��>���h{��g �p�*����?��\?Ӳ&?;��1�`�Rľ�n�<�+S�b�<�oM<�Ɏ��%>>�Z�ղ�=�>"��=ɔi��U6��=<"��=�"�>��=r�D�X��0=,?�G��ۃ���=��r�;xD���>�IL>����^?vl=��{�����x��!	U�� �? ��?Zk�?i��>�h��$=?�?P	?m"�>�J���}޾-���Pw�~x��w�Q�>���>Ǣl���I���ڙ���F��h�Ž ��y��>���>��?� ?�S>8˲>{ ���#(����dN��^��{�[�6��L.�U��럟��-#��������k~��Q�>ڷ���	�>�
?Tg>΢}>r��>�|ѻg�>t"P>��>���>��Z>x8>97�=5�o<lȽ��Q?��'�Ic�����I�B?�;d?}x�>kMf��b�����I�?y��?���?�w>�hg��z*�,K?��>)��,�	?W�>=�û��n<�举����i�����>sؽ.�:�XxL�N�a�Ne?�[?Z`���{;Fv׽��c��E�=���?kO?�~U��n_��o���7��gk���>�q��~�v��t���Xh��%؉�UK���� ��R�>�c-?t��?4�&NM�e#ݾ��]��M@�){�>���>嚖>�-,>h��>H,�53�w6x��NY�(	��� ?�W�?��>b�D?;�-?�!>?�J?1l�>��>],龍��>'�G�H�>��>��'?��0?kT0?��?#�'?3,+>䋾�꾁�޾��?��?��?�?�� ?�`9���L�*R�A�A�fֽH���_���\��g����<8v�<x�H>
_? ���8�J�����j>�W7?6f�>	�>����z����-�<BE�>�y
?�)�>� � }r�pM�u��>Ə�?D��ί=��)>���=�������`[�=���螐=�	��X�;�C� <B��={g�=!t[��@���:���;jA�<;u�>D�?9��>yB�>�@��6� �9��i�=�Y>KS>�>�Dپ�}���$����g��[y>�w�?�z�?��f=��=��=�|���U��b��F������<�?�I#?�WT?C��??�=?�i#?��>�*�7M���^����]�?w!,?*��>�����ʾ���3���?m[?|<a�H���;)���¾1�Խi�>�[/�_/~����3D�x򅻴��7��#��?῝?~A�J�6��x�߿���[��s�C?�!�>Y�>��>/�)�^�g�^%��1;>ي�>HR?�>��O?FLy?�Y?VfT>(8�Pޭ�@������)#>�j>?�>�?zǎ?"�y?�!�>	>��'����in�����J�뽅��CD=��`>	z�>���>3q�>P��=;P��?��/<E���=�]h>Z�>5t�>Sl�> �v>�(z<fG?��>z+�����꡾����Su?$��?�Q)?�C�<-��E�pj��Wf�>O9�?'R�?M�)?f�R����=�s߼������r�g��>�߸>���>���=�![=��>��>��>F���2��7��Z�>?��E?��=yvɿ�l��3=���W��6�\r��,���`�ٽ�u���Q�=뗠=װ��
־W�@�c����3��_�ྦྷj��2uֽ38 ?!^=ϑh>P0�=�U��[=k��=�)>79T<đ0=�s�s�=@C>�B�=�#�=�=do�n��=uk����˾��}?*;I?͙+?��C?�y>$S>�:3���>T����9?�V>��P�-����;����������ؾ�x׾��c��ǟ�(M>�cI���>�/3>�M�=� �<��=s=��=MW�{�=A��=T�=�u�={��=c�>�n>�6w?V�������4Q�qZ罧�:?�8�>W{�=��ƾl@?q�>>�2������tb��-?���?�T�?>�?Dti��d�>M���㎽�q�=[����=2>g��=q�2�[��>��J>���K��<����4�?��@��??�ዿ΢Ͽ0a/>œ9>Ï>�.R��0��^�Rdj���]�)�!?-:�:aϾj�>ȓ�=_�ݾ7�ȾD�8=��6>S=�f ��2\�K	�=�By��7=�o=h�>W�@>@ǳ=�p½�?�=fAY=	��=��O>�>�����k��c9=���=� b>�>�{�>�?xc.?sj?���>|f9���jg���G�>;��=.w�>�E/=^�> ��>��>?ON?�E?��j>9=��>��>�}��|`�9�e�����b<�C�?�Lx?�)�>E�=Uҿ������B�Ϫؽc>?peI?��?�(s>6����޿��0��~'�˺�����<V�'=��@������;TB�<eJ�gʜ=�5�>-X�>�<�>�t@>'(K>���>��>���=���=� �=�� ���^<
 }��A�=���<�'�="�<� �=�ݨ<�b��7Ϝ��&X��4=cļ���4��=���>�D>���>$��=�򳾯]/>�˖���L��y�=�A���"B�;-d��A~�j�.��M6���B>M,X>O����/����?=�Y>��?>���?}Bu? >��b�վ�R���e��S��׸=1�>	'=�Lu;��L`�;�M��mҾɣ�>��>��>j\h>�l,��o?�t�b=��o�4�� �>~B���o�����q�
����ğ�B�h�;�*�D?d臿c��=��{?a~K?Ʉ�?�U�>�l��j=׾_/>Qh��Y�=�w�Zq��-��b(??�'?��>V��;aE�ވ˾>份���>|�J��gP�9�����0����f ���]�>¨���Ͼx�2�[���4(����B��t�R��>� P?�Į?v�_�CZ����O��J�����?lg?-�>�6?
?������=��j�=�@n?	l�?A�?��	>)�F>[/��G�q>��$?kX�?��?�S�?SV�p�c>���0����a��y�����>c��=�;�>=�#?���>�@�>�5�����v������m]2�Z]0=V=�<�>�Y?[�>s���d��b��� �>���>$�>x�P>��f>��>o���1�e�?�d�=�g�t�?�
>8)5>���u7>��v>� u�[I����BM?���>��?�~�a����=%��>����AÈ?V��=A�2��?�Y��L�=�;�>^��>@��=1�>'��>��=~�>��>�`�=(l>�V9>K=ӾɊ>���5d!�~3C��R�D�Ѿ�~z>������%�K��a`��T?I� ���m��j�'/��Z9=�H�<�F�?�f����k�4�)������?&R�>26?�ˌ���۟>
��>���>L�����Sȍ�rd᾵�?���?�=c>��>��W?˜?y�1�|3�coZ�v�u�P&A�e�-�`�����B�����
�����_?��x?{vA?&�<�5z>���?��%�<ԏ�|)�>M/�'#;�g\<=�/�>�&����`�G�Ӿ��þF:��LF>��o?�%�?�W?�KV��7�D�	>K�4?��B?�mq?�8+? �D?a���_�?wM=��>7i?��%?�*?���>�(g>�E>����q��3|�@Ow��/��+��������=w��=ෲ=�м�X�<8� ������Ba�6����KV�|]�<�8=�!�=�:/>:H�>`]?���>|�>�k7?�b�J�4��۲��C+?M�=<����懾��Fo� >>Hi?q�?��W?�hP>'�@�\G�d>�s�>U�)>��b>/!�>[|���U��^=r�>��&>c!�=�l���̹��$���E�<w�">�+�>�X�>5�7�0�>��gC=�|>����k����g� �>��',�SMk�)�≯J?�h?��=Y�߾��1���[�&?��4?�-O?08p?� >}@���~'���Z��{���>_�>�&�����/����u.�ĩ�=!Z>I�����Oa>xT�5G޾n}n��I�ƹ��7T=���U=W<��վYZ�_ �=��	>0h��F� �'���Ӫ�^kJ?�h=����U�R����>8u�>�2�>U�9�..t�x�@�RF��=/D�>�3;>�x��x�WRG�sa����>dWS?`LM?܃?��p�
�Y��0�c:��|ǘ�3���J?�_t>$G ?	�s>w�=�y��ւ��x�ߝJ��>Y9�>���v�H���#��tѾ�� ��J�>���>�
<4�?�GX?��?Q\?qy-?5?G�>��zw��6&?ꍃ?�ф=DIԽ�T���8��F����>4k)?�AC��Ǘ>0v?�?��&?�qQ?�?D�>�� ��L@��n�>Kk�>��W�nV���j`>(�J?[z�>�:Y?���?�u=>�k5�~����O����=�f>��2?-S#?��?P�>��J>y�ؽc�A��D�>{G?�;�?�V?����:&?p ��&C?hj�>��1?�EJ?rc?烈?��?�f�>:>��O={�������[�;���#a��a"8�;^d=J�8=��<�v��	�Q���o=1}=-%��C^�=�x�� ��"Z	=�m�>_�s>Aŕ��0>cfľ�[��D�@>Q����Ȝ�΢����;��*�=x)�>{�?"�>ʏ#�>ɒ=Y�>E��>���J(?4�?�?M`I:ڬb��۾?K�t��> B?-��=�l��S��G�u��Zg=��m?0r^?� X�����s�`?�x_?�Z�_3��žJG\����4QG??�?�JO�q��>2Ov?-Ln?���>Ѱd��m�l󝿾e�qkj��E�=��>���+e���>~�4?H*�>
n>�q�=j8羚�r�"����?̌?��?~S�?�<>�m�/��.��Ṓ��za?���>.ݧ�l8#?����FqǾ����儉��;�!v���7��RY���p��'x#�����<轑ŗ=�R?X_p?�Ut?�
^?�2��da���`�ƹ|� �S�� ��{���E��]C�
@D�ېm��V������e��Oi0=p�a�����?�l?{Ȝ�z�?���5z��zy����>���⣶<a@=Ya=�
K>A���
��/���,���3?�z>�W?<:?:�2�=���<2�xx��ݾ�,�>$��>o��>��>i���*0/�����4;HoĽ�TĽj�w>"�d?�I?e�o?���D).�󄀿9A"�X�,��V����F>��=�Ԉ>�qK�-�^�%�K�@�8au�$������u=E�,?g>P��>��?v%?q�	��(���Ir��=-�}��<���>9�h?,�>fА>t�ݽWP(�0�>iY[?�>�;�>,5��D�2���q�ʀ >���>Qva>� ?��;>7Ђ��$K��������Q�U���>��g?A􈾘q��&b�>,:m?Nݽ�Sv=M(�>��|�i��h���@,�`�>#?���=j5>U�����B����9��?	b?�堾�$�e�p>��(?u
?_��>�ރ?PWv>Tʗ���=!_!?1g?��X? �J?��>�e�;�u��ݴ�<�6���=�y>S> :�=ֽ�=?$3���V���S�p=�CJ=P=1?R�yu�;���( �<�D�=��>0׿�AO�߉�����~�M� [q���;�J�����Fо�1�c��[��%�1���%���"�sf�ɧ��(p��O��?� �?#P��#;]����
hj����� ?F:���f� �Ҿ-�7�Wט��5�����jY"���_��dd��8e�S�'?�����ǿ񰡿�:ܾ"! ?�A ?I�y?��@�"���8�� >[B�<.����뾱���
�ο.�����^?���>��l/��v��>̥�>�X>�Hq>����螾�1�<��?7�-?��>{�r�/�ɿa������<���?-�@��A? �'�Ѫ��A=���>Xx?�C>�-�w���H��b��>��?Fs�?T'D=�X��3�6xe?'�<x�E�������=.��=�D=��
��M>ђ>�%���A�k�ٽ��5>�;�>�������[�V]�<;.^>7]˽� ��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=0��FſCV�Ӱ�
��<��!=|�򼟀뽈����)����J;����XN-=���=�l>�'�>�[">��>�W?��g?�
�>1FG>(����B|��"žO=>�R�rR-��T���G�x���_�n�ݾJ&���Y-�?"���ξ=�+)�=h-R�d����� ���b��F���.?�@$>!�ʾ��M���/<tʾ�Ϫ�3��f���̾5�1�fn��ʟ?��A?!���/�V������1����W?�f����&�����=
ű�+=��>��=���A�2�ЇS���H?� ?;ھ��־a��>7iA�q >��?s�>y26>�g�>�	?n4��ꖼ��M���j� 6�>��?u��>���+!��?��?�\��Ge��w>�1��V��	�<��>�@���׽��?���[� ���w�x倾[��=��m?CS�>�;,��a��A�����t�K����?3�>N�C>�E?���>����(��b�߿$��<~r?��J?I��=/��ݺ���iվ��?~�_?o>�k�R�<n-��D���~%?s�H?��%?n���<j�W��~����2?��v?�#^��l�����ʲV�է�>'��>���>Ǭ9�y��>�d>?p�#��P�������g4����?$�@Q��?�^A<f�����=?o��>�O��cƾUG���V���<u=0m�>#m��f[v�8����,�ף8?ƛ�?"E�>fM��@�����=��ľ�k�?��?L����C=����v������>���<�< �V�,���7.0�m۾���l��ES� ߊ>��@�Y9����>T�O��+�UL¿�H���yѾ�us�!n?��t>)�Q��о����At�-&J��u0�Z!�ߤ�>Z�>�[���}�� o{��w;��:���j�>�2�?�>$V���������<8��>�#�>���>�������˰�?za���ο������W?\-�?�G�?�?��J<��r�u{z�M��;�F?^�r?�Y?`��Q[���:���j?���`��_4��pE��DS>��2?��>X-�a�z=�^>�6�>bZ>�/���Ŀ���x��AǦ?�k�?�V꾭�>�p�?5�+?�v��홿uY��w:+��ܠ��xA?F�0>J%��*!�w�<�����/�
?�x0?���)��]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>�`�?v��=��(?�i��덌��xm=Q����=%f@<Ӹ ?Z�,?�v�>�=�3i�WI5�z�e��^�����I��î>��K?��7?��!>�갼Q./���$�_��? ���QO��)��Pc=N��Ύ>g��>�X�;����֊,�W?D,�~ؿ�w���y'���3?�>�?���nt�)I��_?1�>/:�/(��|��v���?!$�?%�?�U׾�Ѽ4l>�w�>d��>w|ս�y���x���)8>�B?:J�5����o��x�>D��?�@Eޮ?��h��0	?"��J���n~�	|���7�c�=>�7?%��Y�z>�|�>���=�v�u���	�s��,�>�*�?Yv�?���>��l?�Mo�� C��23=���>�Uk?K"?.�i��V򾎇C>ǫ?����ێ��4�1f?��
@<a@��^? ע�N�ܿ�����о�Aþy�>���=�#w=8�����<�����}�J;	;8e�= ��>�>W��>��)>�>,>'_�=���d �iʞ�;a��A5@�@�3��g3�<���6�%�ls������ݐ��F(�܎u�UBZ�}�W�b�;�P��������=�
?-?��?� ?Y�@=>�">5�˾��=}����M>���>>,?ڸB?�~?Z>��w���o��j��҆��md�3��>�D�>!o�>��>���>�=�4�>�#k>&�v>՛z>�2>.�.���%>zda>���>�!?<k�>�C<>��>Eϴ��1��l�h��
w�e̽1�?����R�J��1���9��Ԧ���h�=Fb.?|>���?пe����2H?#���{)���+���>}�0?�cW?�>"��w�T�::>7����j�9`>�+ ��l���)��%Q>tl? �f>�u>��3�Ke8��P�Q|��Tj|>�36?�鶾�D9���u���H�Rcݾ�GM>�ľ>4D��k��������ui���{="x:?��?f8���ⰾX�u�$C���PR>�:\>rX=1j�=YM>.dc���ƽGH�l.=L��=��^>!�?��1>��=�K�>����Q��-�>CC>��&>̴??��$?����C����}��d5��Wg>���>{�>�r>��N����=�2�>5�q>�%��W�Ҵ�`�K���Y>p�z�nM]��j�엄=�������=��=5>���N��>'=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ/E�>�2�l���M���v�7�b<��>�uJ?B���fDK��(9�߫?	��>B���U���Uƿ��m�#��>)d�?=��?�nc����`�@��;�>���?ѼX?a>�g�vT��h�>��<?��N?&��>_���9��?+��?M?�CI>h��?�~s?�c�>N�x�Qc/�Q6��r����X�=�d; T�>՟>�����gF��ԓ��e��װj�	����a>v�$=��>�z���)��=3q���^��7�e����>;:q>��I>n,�>I� ?�Q�>�ř>*}=P����ˀ��㖾Z�K?я?r��%Qm��T�<E��=�=^���?�3?!P����ξ3��>�r\?«�?ѤZ?�m�>���8k��⿿�������<�uJ>���>4�> Ɔ��J>�Ӿy D�G��>��>OV��پ���^�d�>�!?s��>�m�=��"?�4#?6\>�Ӣ>�{G��D���RC�p3�>���>�n?��x?�B?���8�6�u��x+��S_V��Y>�)w??�P�>4���r3��=/#��>��\����?49`?L���Aq?ᄈ?�<?��@?TcW>�(��ӾZ���&j>��!?H����A�K7&�	9���?�U?���>Ւ��fֽ�gּ0������?8'\?sG&?�c�2+a�)�¾��<m�'�m�a����;��N�R�>��>���Rv�=b�>���=�0m��y5��m<.b�=���>;�=�!7�����B,?FME�1�l"�=��r��D��->	.L>������^?/q=��|�����z���4U���?���?Kr�?�紽�h�0=?��?d?b�>Kr����޾Ci�v	w�x�g���>���>o^o���/�������Q9��hNƽ�ν˃�>�.�>f��>�Z0?� )>�m�>ap��W����|�N�KI��8��6�Z	1��%�I��Ev��S>;����rn��>��1�E�v>��?�_>H�>{��>�*�=�d>8��=2#�>RR,>��
>�{Z>��>i<��+=�LR?����|�'������4/B?�qd?�.�>=.i��������~?���?�q�?M,v>{h��++��k? F�>����o
?t^:=��w��<_K��:���P�������>�A׽u:��M��yf��j
?p0?娎� �̾@׽3�J�����17�?4/?�@��@��Xy���v�mZ�TiP>'D��69��@&C��I��p���?e��=x���H��`��:�_0?S�?_la����B�����e$�3��>�,?j%�;��>� ��Uk]���3�~��$6����1[?L
�?��>�)R?JK-?��\??�X?4Ğ>��>�碾J� ?��E��{�>v��>jW:?��,?�0?-�?�&?_]K>���@Q���S�8�?�w?��? �?��?E1x�w����J�=���_���F��h��=��	=h��C���%�=�Xq>~�?�
�j�8���%�o>�5?Z��>Ï�>A���ay��V�<�>�>~Q	?̎�>dU ���p���	�+��>��?��
�1�<lD)>���= �m���;�˱=-�޼砩=��a��Y?��,< �=h�=�Wߺ�Y�����:��<�8?�Y?�s�;�;�>w���l�a���r�f��=3�?ק?J
�=.��ft���9���OZ����<�pR?�^�?}�C=�;�=x<Gb�*ux�&�;]�����0=��+?D?u�$?��?4?�E?�K��+����_��nd�*<P�l��>�-?^�>�x���ʾ$�����6�"	?o�
?��\��p��^ �C濾����>(4�����z#��	�?�]�	<\Q�􊽽���?B��?��q�tV1�uwվ<�� ���H?=,�>7դ>�??��#��sd�m��N>��>��R?��>�/P?=�z?[�[?��T>c48�筿���K�8��>D@?�r�?|Ŏ?��x?!4�>
�>��*��F�_����!��l������T=M�[>ȶ�>��>�\�>�s�=D�ʽ�𮽂�;����=�zb>���>���>�)�>�nw>b�<s�H?���>�K¾a��}���]O������2�r?�6�?��-?�~	=֢��4I��8 �兺>ä?�Ʃ?��.?��L��=�=�ڼ�5��c�j�N��>��>O�>�k�=)�W=�">%��>��>	.��x,2��9@�ܾ?vvF?v)�=�]ƿpbr���u�}���\!3;a���=F`�]B���,f���=񁗾Z���9���$\����2S������J<��`3��b�>�{=���=���=���<���o?�<M=O=�^�<�7=+g���<��4���9��@:�n�<��`=/�6�#�ʾ;~?CLH?�,? �D?�v{>=>hY2�9S�>E���#r?S:X>*�D�Nƺ�eM8��u�����:Jؾ��׾�Je�3䠾�>�K��s>&�5>E�=Uʊ<��=jl�=���=����k=��=`]�=���=G��=B|>5>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>q��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��E>��>YrR�e6�UKV�`i���E��0"?�>�
Ǿ	�>���=�Iݾ1Ⱦ�>�<�->�9�=S@�ĄW�kP�=��b�C=?�C=ϔ�> PT>W�=�������=��d=s��=�J>��;P�6�����X=Z��=Zo>jG->{��>�?v0?;`?�ֿ>�m��Ǿ�q���u>.-�=5��>�<^=�P>>��>��2?��A?D�J?f\�>ts�=�#�>��>G�+��Tn�������:��<��?kć?E��>� =S]=��!��?�q@ֽ��?ۦ2?��?���>w	���տCt)�A�M�a��>j=�i_=��/\��N~��ph��z4�{�1=��>�D�>� �>��X>�t;�y<[�>O��=�e >��=>�=��B>�J�=��=����=÷���>w=<���/U��"h�=xY�<��=�P��(?$><�>!�R>ɸ�>�nU>�Ⱦ��N>��h���[�'J����A)-���^��tm��+�aG����=.�>c��=�U��u��>T�W>
� =K��? �x?�o�>`rѽ�7�������p`8�=�Ƚ�>�ѽ���0(C���>�:��&��>��R>�D�>�2�>�O���J���<sˡ������>ƒE��c!�����`��𥿔���f�����[?r|����<�r?U~T? ��?��>o/W>���n�b[;�Nվ�� �ք���0� �<?+d?�?��������P=u��>�ʾ5
Q��t��MO�t�R=ǋ¾<�> ���� ��U��I��'���/�;��P�>C�m?{�?�Q�=� ��p[Q�L��pյ�ӂ�>��H?a�!?vq�>iN?k>齹����������'?팻?�s�?����mL=����G�>s��>]ӕ?�D�?��h?Nz�6��>1��_> ov=�S/>��F>��:>?.E>v?�K�>\U�>�����I�5�����]��W��=�}�=I>>⭀>��'>�1=�;~=��>nB�>�B�>(u�>��>�U�>q>h���E0���A?���=5~S>��4? n3>�cG>˜��XcM=�����Z0�fV��_˽P�</9����]��Q��N	?�jĿ��?�]>3�/ ?�� �x�^�E>�ǐ>� �|�>5�c>ir>�c�>Be>>�T=��>���=�?Ӿ�>��;f!��-C���R�@�Ѿ��z>à��F&�Ҡ�n���DI�Cr���i��	j�`,���<=�
A�<�G�?£��&�k���)������?_�>�6?�،��	���>R��>�ō>�E������ȍ��bᾌ�?���?'i>'��>5rT?>�?��5���;�sE\�\ u���=���b�}�_�I������N$�.ٽ�@[?��v?��C?}�<+�}>+�?+C(��^��ģ�>�/��D<�yLH=���>����0�Z�� پ<�þ�&���K>��n?��?2?� W���v~�>��>��?��g?�bK?��H?�4"���2?2Ɖ=��<?�?0�a?b�\?��<?���>V��>�A�;^0�dkc�X���Ĉ�LdW��C2��k�;����5=�����,=M�_;��=�nF�#F�P	�;�����#�=kOp<`�C>F��>�\?$-�>�*�>�6?bK*��:�����,�0?JQs=E`���q������"���>T�=�`h?*��?<�\?m�d>і@�v�C��#>�R�>;l&>%RX>�>zཱུP@�:��=�^>r�>^	�=JIQ��	{�|�������<��>���>�-|>+�����'>_r��*3z�g�d>�Q��Һ�\�S���G�"�1���v�,V�>��K?;�?���=�_�����Hf��.)?B\<?3JM?��?� �=<�۾��9�>�J��C�p�>�Q�<���￢�E"��x�:��:��s>Y/������?b>2���[޾��n�IJ���q�M=@��mvW=��C�վ�s��=�E
>=����� �����ɪ�� J?��i=�Y���:U������>�ݘ>c��>rE;��'u�vr@��#=�=o��>z�:>�җ�S�tG������>a�E?.�\?Pc�?\6���q�-�@�6j��9o��#�󼔜?�>,?�>A>�F�=�Z������Fe��KH����>P��>����qH�������#���>�?-�>&d?Q?ZJ
?�_?\(?x�?[��>��Թ��=&?y��?�(�=!UӽT�S�#�8�o�E���>#)?��C����>u�?�?N�&?KQ?!|?��>�� ��h@�`I�>��>��W�T����`>9�J?>j�>�OY?���?Z*=>T5�g������� �=�>h�2?�F#?]�?❸>�EO>x���0Ĩ��\>(b?��f?U�q?���=NN[?+l���>{,��!�?�^V?�I? �o?J`}?�8D?w���=ƫ��B��eǟ<�'���nR�`Ӽ/ I=�X>�3z��rɽ����9m�dV	<
Ǯ==)�=���_�ϽS������>[�o>������4>�º��|��ԐH>od�����H%s���3�� �=$Vz>��?Dߔ>*�-���=�q�>�F�>3�|�'?9d?�?���W�]�fSھ�']����>�m>?���=[!k�����S�u�_My=�jo?[�Z?dhf�YM�*�d?Ӱp?׌ﾆ�@�������5���q?��>�e��M?@�? �?]	�>9Ik=�O|������a�������=��=�X�h,>�%&�=7��>��>��`>~��h��]�u@6�	q>?� ?�}�?%��?�LZ>@W���пdA	�љ�m?�>&ʾ�#?����ɿ��8���r�/�ܜ�ck��o�[�rM��wEG�%�~���|��q��e(?�\?�,�?P�d?0z����������r�M�g�`޾���\H!�EW��(J��y���.�����������������R���?�!?����~�?�|������Ծ��K>&?��3� �m/�(������!L���q¾����+/?,G�>g�?*A?_�a���mz\���A��^���8>�X�>�,�>=Q�>w,�����ZK�/���?��,�|��X|>2b?B�J?F�p?��_4�I.���J��VS��*���=M>�>�a�>7(`�Q��V�"�K�?�h�q�����8����ϼ�=H�6?�-�>�Ԭ>E�?Zt ?�E��w�������8���G��U�>޸^?�+�>#��>7�����H��>ٹl?B��>�>*m��GW!��{��nʽ�	�>��>u��>��o>j�,�R\��a�����9�7>�=үh?҅��>�`��߅>�R?u�:R�G<�p�>��v���!�����'���>3q?�U�=�;>�_žr'��{��C����?'A?�s�<(�i�>&n'?H��>��>` �?2��>%Ȩ���O��?�Ze?�pK?�?Q?�d�>t�5=�$��蜽j	��H=v��>��A>I��=O4�H3�B�\���x��=�>w߯���P�	���q����&��Q�=���>iJۿ�K���ؾ<��v�H�	��戾�T���n��:����������z��&�Yc&���U���b�����'(n�1M�?���?���rk��H��$ �kC�>H�r���}��!���|�����_��M��]�!�E�O�'�i���e�P�'?�����ǿ򰡿�:ܾ4! ?�A ?8�y?��6�"���8�� >]C�<-����뾭����οA�����^?���>��/��q��>ޥ�>�X>�Hq>����螾�1�<��?7�-?��>Îr�1�ɿc���r¤<���?0�@�B?w
'�~�쾶ea=?��>U	?;C>*23�z������*��>�=�?���?�?Y=|@V��%��Rc?�\�;�AD�:�3��\�=:�=#z2=�D���M>n��>� ���B���߽z�5>� �>��~>��Y�(i =M�[><J�VԬ�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6��{���&V�}��=[��>c�>,������O��I��U��=�o��5�ȿ6�$��@5��("��'�;��˽bI��:Ž#���T޾#
��.)��<�=Z��=��@>(t>_�s>9?�=�&K?�3d?��>eQ>�J��O�����߼ن`�"�'��BT�~��AȾ?1꾬�ؾ~��u�V�%�m=ƾ#=���=86R�Ǘ���� ��b���F���.?�p$>��ʾ
�M��B.<qʾ����榄��楽/̾Ԙ1�U!n�@̟?W�A?������V�>��|\��}��Z�W?S�����謾��=�k��X�=$�>j��=���m!3��}S�7X<?Qq?H̾%�����>���2��=��"?J��>��>L4�>�3?3�G��B{���@>�V=�n�>ձ�>KΉ>籾f ��hy?�h?�)�Ei���>c�(�g���>�}/>` 4����8DE>��=e
'��3���6B�.�c����?�ψ>sI��z]�0���wMj�>��>R(�?A(>���>�2C?�37?v	=������,?��6�>��?��?�	>�XS���ʾ��̾3�w?R�T?�+>a�پ�O����L�!�U=D?��?��h?��>E���ԓ��@�B�?��v?s^�xs�����M�V�d=�>�[�>���>��9��k�>�>?�#��G�� ���{Y4�%Þ?��@���?��;<��P��=�;?h\�>��O��>ƾ�z�������q=�"�>���|ev����R,�e�8?ܠ�?���>������s\�=�����d�?��?����@aj<�
�Cl��q��]��<��=����#����L�7�p�ƾ�
��ۜ�܇¼ƽ�>|U@Ƌ��6�>Kt8��(�jWϿ"��Jxо�8q���?�t�>lmȽ}�����j�<Nu���G���H�|���L�>�4>ժ��������{���;�+]�����>��?�>F\O�oK���u�� R�;1g�>n��>I�>K����绾���?�|���2ο�Ş�?:�Q X?�I�?���?�f?N�B<W t�vHw��ѻ��F?�r?�:Z?؀�?�Z�1��n?�g����_�`r4�b�3�A=N>�]3?sM�>��'�6��=A>q ?�3�=��&�M@���W������OU�?���?���)�>&Ǜ?��3?�h�Wӓ��稾.0�Ah�;��F?2l>>�麾<��6�6���r��?Rh%?E2���]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�I�>7�h?g�=��-?��>�J��Z�=yW��V$<��4><��>��b?ڻ�>���=��׿+�*�/��SQ�����lQ��,�>�A6?�7?'��;�Q���3��I꾾������}Z|��$�^�h�H���8�=�s�>��>!5��R���?�o�ٖؿ�i��h'��44?��>��?m��l�t�T��p<_?�x�>�5��+��@&���B�;��?�G�?r�?|�׾�>̼o>��>�J�> սt��^�����7>/�B?�gD��'�o�s�>���?R�@iԮ?�i�A�
?*#��L���V{�o2��&A����=�;?��ʂ>���>��=�`t��g��P�u�A�>�7�?�f�?tB�>6n?L2n�y�E�PY�<�å>�-i?ʾ?3��<������>>BT
?���u���j� ��[a?h
@��@�`?BM���ֿ�>��r*־D���1/��Z6���>�1���;Hż����|z����>�V�>N��>~�>�L->,��=C58>�P����%��*������?�Q�?7!������~.)��G����-��]u�٬h�8F�����༊Q������[@�ArA>p?U� ?e�Y?�p?ӡ�=�I6>�yľ��H��o��=ii=�C�>K$1?]C? )?�#�<���-�_�z��\>��-V�Ľ�>�0�=O�>���>S�>=|qR>P;g>�d> �
=al�>��>7�=&��>	u�>S��>���>�H<>��>pδ��1����h��w�=/̽l�?U���N�J�D/��51��P���Ic�=:d.?�w>��4?п-���1H?�����'��+�5�>�0?�dW?ݕ>����T�v;>�����j��c>{, �ql�I�)��Q>�k?��f>�u>֐3�P8�N�P�P����_|>v46?����w:9� �u���H�biݾ M>���>�E��s������5ki���{=�s:?��?�������u�U/���KR>IH\>�=�N�=�eM>�dc���ƽH��.=���=��^>��?tq+>�܊=F�>Ȏ����M��G�>�N?>g�+>FbA?��$?�D��R����-���R,���r>�y�>e�>8�	>G;L���=-��>��g>�S&���}��`�wD��HU>���i^��xz�){=�����=gO�=5� ���@��� =�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>�w�qZ�����e�u�ȳ#=}��> 9H?1V���O�U>��v
?�?-_�𩤿{�ȿ�{v����>_�?���??�m��A���@���>��?jgY?�oi>�g۾�_Z�ʋ�>�@?�R?g�>�9���'���?�޶?ӯ�?�BI>
��?Hxs?#��>�Zw���/�p���W��>;{=N�V;�%�>0 >w��=�F�����ri��^�j�v���wb>΂%=��>��㽀���6�=�э� @��>^d��n�>�q>=�I>ma�>
� ?�K�>Mՙ>N=�������c����K?R��?����n�Y��<��=}�^��?�04?6M]���Ͼ��>��\?#��?R�Z?^S�>����<��濿���m��<��K>U�>M�>��CK>��ԾI<D�S�>͗>���8 ھ������CE�>hh!?׎�>_Ȯ=sz#?�O?��Z>>�\>��?�����ޅh��1�>���>���>�h�?�*?,���I�[��� )��ך����=��?+?���>0���⚿{"�>:rҾ��D��l�?��?�B����E?��?a�?"[?��?W�M�Ƴs��q�#[>#�!?���ūA�
>&����Q�?xS?���>ă��U$ֽ7�ռ����M���?�"\?�E&?0��sa��þ��<l\!��T�)��;��C���>�8>�����g�=�>u(�=�m��6��{d< �=xj�>5��=w17��_��1=,?��G�ۃ���=��r�?xD���>�IL>����^?jl=��{�����x��!	U�� �? ��?Zk�?X��?�h��$=?�?R	?n"�>�J���}޾7�྾Pw�~x��w�]�>���>Ңl���K���ڙ���F��]�Ž�����>���>�n%?���>*��=`%�>��[���9�2��i���be����|J�zL �c��:Gξ���Ć�w³���X�N�>�-����>=��>��p>m�>�]�>�>;�U>M&>�Zv>�T�>'41>�o>���=q0�<��<��U?d���g�(�h���]��op=?M�c?S��>�P��n{����[$?x��?͚?�.d>/^n��(��)?"�	?�ց��?!
v=m�=�<�������ʽ��^ĝ>鑵��A5�X[J��Y��T?�=?J�*�
/ݾ����#g�ͮ��(��?E\>?�i���/���`���&m�Y�H�0�6> 2ž���� t�{���)������L���CLZ�h����(?�!�?\/�뇒������y��ԍ�e�R>(f ?lC�>3��>ȫ<6>��vy7��>�55⾽i̾�g?)�?��>M?�Z/?j�K?��M?��>+ǵ>d����>�(�����>���>�D?�
0?n�%?�?�/*?�8W>�W�B���$H侖w?�z?�E?��>��?��c�|�(�����߹uJ����9�;�-=��L<҂��d9����=�Xm>�s?�d���8�g���	l>�b7?J��>w��>����<ǀ�դ�<�[�>M�
?b�>� �v�r��P��s�>i��?�����=�*>��=�=��X�����=ւǼ3�=.�t���9��,!<�=.��=��1��!Y9;��:w�Q;Vg�<x�>F�?;��>�B�>�A��j� �5�����=NY>|#S>>�Gپ�|��4%��d�g��cy>x�?M{�?��f=x*�=ύ�==���\��������{�<r�?{E#?�UT?���?g�=?�j#?��>�+�IL��S\�������?��3?�Y�>����žɝ��2&w�|��>9O?��`��RN>�s�BF}�#�L=T��=���P�T��]���f���c=\o������?m�?(.]�L��Sd�냢�D�7�F=?���>�c�=F�.?�6���y�b��F�F>!�?�A?V5�>m�O?5{?�[?q�T>t|8����{���L@��t!>|@??�܎?1�x?M�>>��)��?����o �S�î�|U=�BZ>F��>��>G+�>�m�=_ɽ��?�>�j(�=x�b>:]�>i��>b"�>̦w>@`�<E�I?ԃ�>�6��u��w��}��f�%]z?���?ɜ-? �u=����.C�K���l�>��?9�?TX.?.�5��K>��rR��Cֆ��6�>�>|��>�w�=��<v3>1��>���>o����9��9��n?�kG?�O�=]�ĿM�x��y����n�����`V��6�6����X=b��L^=�.X��K�8��O��-�k�pƬ�3������?�>�9o|e>F >p�}<�=鳃<J��=��x=�L�=��V��.=J
���c<gQν�
��i �Hx';�������Y?>?d�+?�B?�sx>�%>�����k>��5_?1}>�4t��⳾�M=��ު�?k����ྋ$���f�3J���>\���/>xM>U��=ëy=2x�=)�=��=ڷ<�x�=�C�=��=RE�=��>e�>�P>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>RK;>�s>��Q��{.�ղS�i^�ÌW��� ?Ɯ<��о��>.+�=9޾�)ľ�?&=4p1>G�n=����y]�F7�=�q^��KC=��N=."�>�	L>���=�+���=�OB=�=��P>���;� �����B=�S�=��a>r�)>�>�>IX?�/?. d?,��>�j�!�̾1&�����>�x�=64�>�݉=�G>L6�>7?�2D?�K?��>[�=��>_1�>��,�ުl����]����<�<W��?��?�g�>��Y<�nB�^����>�l�Žj�?/�0?$�	?̽�>2���tٿ,�?�sIt��*��(e��0�A���	�DҼ�O��>`
���J��Y>F�j>� �>\�>{5�>fN�>E'���8�>��=�Z>��>=��,��<�Bz�h~�=�G>ޞ�=�l���0��T�	� ]K=l	��%p�nm�TJ=@����>��>�q>��?��W�9����U >{V��:yN���>�򸾂A�w�P�􂿇���NN���=攠=+o��؏�_��>h�6>ob>b�?(�w?OI�>��U<e���^������|�%Y`���ؽ�Qb�x�H��GX��^I�����U�> Œ>"��>���>^��<�>���O=͡۾p�!��@?O�$��o�=Vy����U��_���D��# d�ܽݼa�L?27���v�=��{?�wl?�v?��?�
T�����&>����mnʽ4�.�W���N�B�Z�?�?J��>�����Q���)�Xu�=�a�>��=�=��㖿��羪�:>C�x���>0��{.��b$��앿`鎿r��4�F�V��>�)l?=��?���F���"wm�A�J I��G?�n?ƌ�>5�?lhY?]����� �q���o��&�?�?W��?�u�>��=�[.<`��>#�?�ԑ?��?I�s?�R��A^�>�����<>�	��%?�>M{M>��j=�>j�?"�?"��>^꽇��ֹ��M�Ҿ(KW��/ �B�=���>��>�A>�D�=h�<�WC����=�>E��>F�Q>p��>��>����C��k%?�u�=��>7/?7j�>�'J=�?���9�<�,����B�cE3������ܽ�T�<��4�<=k��D��>G^ƿu6�?\�Y>���?]y��m+�� O>OHW>�{ٽ�m�>��->l\}>k7�>�җ>�$>wy>7�>p7Ӿq�>����A!�� C��R�@�Ѿ�z>�����%�y������/cI�ו���`��	j�g2��aC=�6�<�A�?������k�-�)����{y?�Z�>�6?Ȍ�㹈�Ѣ>���>�͍>�=��"��������\ᾍ�?��?�;c>�>S�W?�?�1��3�^uZ��u��(A�Ae���`��፿֜����
�@��,�_?��x?QxA? f�<{;z><��?7�%�hӏ�j(�>�/�e&;�I<<=�,�>�(����`�ǯӾ��þ�6�]EF>a�o?y%�?Z?�QV������hX>��>_�?po?;�R?N�??�HO���M?�n���>	��><g??��'?�?�ȳ>J/a>�r�=�Q��䊽HVa�V<��E9��z��x�>��<��T��㵚<[�=-��X�\=�>�Ú=��>��ݪ=��>xt�=���>�T]?��>�:�>X�7?�
�~�7�/x����/?Xr8= ��<��u����p�j>�7k?��?��Y?�nb>RMA��mB��u>y��>["&>�(\>��>lW��3E�N�=ٖ>>�(�=��X�н����	�`5���<$\>t��>�#>0"���0>N7��zF�W�_><�S���'�G���D���/��2l�V7�>�K?�|?�N�=Yc龷���hf�wd'?� <?��N?$Y?ㆴ=C�׾�~9���I��p&���>���;��
�%�����g�:���;�,s>އ���`e��jh>=[�[�����S�|E
��F>�y&�� >�������X��1>u�J>�t��'�+�ĥ���ί�%�;?�ڎ<Z�����J��1���T0>u��>�g�>��b<s�
��HQ�� ��%=.>�U�>X�a>�==�޳�>�G�{@����>1;E?��^?9�?N��;gs���B��T��갣�DO���i?�ǩ>�U?�T>>���=���-�� e�ݾF�Q��> �>�[��G�����J"󾤯$����>l�?K�>��?ISQ?�
?վa?Z+?vl?E��>m���[d��\B&?���?Cׄ=b�Խ��T��9�F�|�>h})?�B�H>�?��?��&?�Q?d�?�>]� ��E@����>�U�>p�W�Ha����_>&�J?���>�>Y?�Ӄ?}�=>l�5��ꢾ����"w�=S>��2?�7#?�?D��>�@�>*�$�٩%=�P�>��d?Y�~?R�V?O+=��C?o�;��?��?�>ȉ�>�+?8qh?�h?#*0?ⴃ>؀<����tG�D�2��+)=��;F��:�	�=�r���\!�掍�C����Q�*:ͽ����ŕ=�u=�8����o��~�>�%t>����1>��ľ�����@>���W0��̦���]:��ȸ=�}�>)�?���>�w#�b��='��>nE�>U��+J(?��?�?^K;b�2۾t�K��ް>��A?��=��l�+n����u���i=�n?so^?�@X������c?E�T?�~ ����7���P�q�E��Y#=?n~�>4:����>��S?G�]?���>���T�c�Ğ��2]�"jx�J�=Ğ�>��FLT���K>9�%?�݄>���>|�S<?]��hS�'����Y?��?� �?XU�?v�t>�J~���������w��\V�?6:�> �z�I�?w��=�0��F��q��|��)/F���	�����}t�����?Q��>�9>H=Z�?tK�?��k?�-�?���.�t�n~s�oE���2������(�4�E@_�2�l�a#��Ō �@�4��>���/�=k���w�J��D�?!*?�$����>ˌ����7*þq�B>B����cҽmCv=��V���=ahc=؈R�y 3�Z���[i!?���>}��>z*A?�YV�
�:���.�9�3�K@�[�#>,�>.��>Uj�>]O��Q�>��0����ξ�x���CĽ3�u>,�b?�K?1�n?{�	�X�3�c��*�!��r@�x᥾��<>�]>��>�R����5&��v>��r�6��:���[�Yɂ=�2?#�>[��>�F�?|�?B�
�ַ���$���0��R;��>�qd?��>:q�>�ǽ����,�>�l?9F�>`��><Y���!��l{��ɽ��>M��>���><#q>��,�L�[�DQ��k���s9�;A�=T�h?C�����^���>�%R?�@%�F�d<��>[m{���!���N�&�B�>�?���=�D=>j�ľ�m�"�{������&?ɥ?�̑�Z�'�䜁>��"?g`�>���>&��?Gp�>���wV�/�?�U_?TlK?��A?�>l?=Rޭ�"ƽv<(��/=R�>\�]>�	x=[u�=����hZ��b"�,V==��=J����½|<�bH�v�|<�m�<�,>@mۿ�BK�x�پ7�O�O?
�舾����c������a��5��=Xx���=�&��V�A7c���Ըl����?�=�?À��g0������0���k������>r�q������g��o)�����b���/d!���O��&i�\�e�Q�'?�����ǿ񰡿�:ܾ2! ?�A ?8�y?��3�"���8�� >JC�<x-����뾭����οA�����^?���>��/��j��>ܥ�>�X>�Hq>����螾j1�<��?7�-?��>��r�1�ɿd����¤<���?0�@�A?�(�����$[=���>�	?Q}@>��0�I�f��7�>�<�?L؊?`�M=@�W���*e?W�
<>OF������=��=~�=g ���K>�ɒ>�V��@��߽�V5>b,�>���0���\�A,�<��[>g4ٽٗ�5Մ?,{\��f���/��T��U>��T?�*�>Q:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?:ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=�6Ἶ���{���&V�~��=[��>b�>,������O��I��V��=���`�ƿ%l$����� =8���Z�[���1]�]l��Sn��*�k=:��=0R>���>IV>��X>zKW?F�j?k�>o�>����V����̾���с����D`��ko�.L������=߾A	��k����`ɾ �<��{�=F5R�j���~� ���b���F���.?��#>?�ʾYsM��e"<�1ʾĪ�3��~��_�̾@�1�� n����?:�A?d���)�V������-չ�#�W?>��.��બ�{��=ꬮ�i�=�y�>--�=�R��$3�ǪS��o0?GM?����:C��|*>� ��=��+?ԓ?��]<�8�>>?%?�!+���5[>X�3>���>���>�[	>{
��n'۽�?�T?%
����#�>�X����z�_b=5>FG5������[>14�<w)����Y�۾��^�<Slg?�->i�#�+�`a"��e>>9v?�_�>��?#9?�2?Xo����&�e�b�,��C�=bHr?铅?'Ģ=(�^=�ȑ�����?�h? !�>��]�q���	V�����?�n�?��$?-Q�=b|�����1:�C�;?C��?f�P�堿0>	�� 	=\"n>Ï�>�q?+�?�b��>@.�>�)>��7��
F��Q�P�Y�s?r9@�	@6�`>?S�	_{��3?��>����������ؾ��X>�2 ?�־ o�a���L�Z�+?N\k?M��>A�#�7�ξ���=�߸��O�?Bp?LT��'Fv�Z>��%���C��c�U�F����{>�򅾱��d\G�Eؾs���`�������D�>��@��Y�H% ?�Oھ���տ�1��ޱ���͒���?�F>��p=b��ڰ���k���z�j7���!�9��>��+>�F��_p��3�����K�6����,�>C&�����>[���(2оJ���"��?$�>J��>Gp�=���F$��rؓ?�	�`�οMa��'����Q?[f�?PT�?e��>��<�ǽv���`�<��h?4�?&�V?V]=3J��AF�i*k?����ǀ`�s 4���C�/T> 3?Ӳ�>��-��Ȇ=��>���>ˑ	>��.���Ŀ�����'���:�?Gz�?���O��>�"�?F�+?7����������_�*����:k�@?�P0>�{���{!���<����h+?ʓ/?#�����]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?&��>��?��9=��?�i�=����H@�;o�T=��=�
����><]P?J��>���= �ܽRm�J�J��NR��.��J�泶>P?-?�>|�I�������-cF�t������UT&�u軒!�;�jh>Sx�>�Od>v�������cA?���Q�ԿQ3���D���=&?
��>��L?�W5��̪��(=��x?a��=Q���Ž�F�����=��?���?/��>�6þ�׽>� >0�?���>G;d�|2�Or����>��?��8���>0��>�;�?`� @.��?"�u���	?��n���D~�!���"6���=�<8?M�uz{>�2�>��=G�v��{���t�"��>�R�?b��?
X�>�Pl?�5o�:xB���5=-@�>��j?��
?�崻|���C>�?���!���w�Sf?��
@�M@ë^?ἢ�TԿ*m���ݾ-�վ(�=�k;>$�<|�N��r
��F�;�M�>�A�>�І>Xb>P->K�=���=����� �Cͤ�+��U/T�w�,�j|I��f�+�6�����z���~L��������B���0�px8�n#���J�(-����)>V�m?��6?%��?�?����g�X=��վ`���?��Y�=�>gJ&?rQ?%,?�Q_>ڢ��W5d��w�o0��:�Q�̗�>�*e>�?�S�>���>~M=o�2>�H�>(��>��=��=\>�B`=��J>�U�>�+?_<�>��<>��>�ʴ��&����h�f�w��oν��?���|MJ�-𕿄ڍ�<ζ�㿠=�t.?�+>`���Cп?���H?��������B+��>�0?�YW?�>�c��c[T�ZV>H��~ni��>����5�k�P)��vP>�<?S0�>*u>��;�s�9��Zr���پ��=�F?/�վ�Wh���S�P~_�\N�B"b>�?�>OzN���(�-柿�p��_���T=נD?D	?j�z�O���V��O
�;'�>b�=>�;�Q >|>w�����D�����<���=�>q�?#,>Ъ�=���>Q'��=O����>�WB>�,>U@?x%?v�	�|���^����-��u>�h�>��>h\>�K�H�=��>��b>����@�������@���V>�ք���^��Lr�wl{=�r��%��=��=����S?���=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾK��>������Ly��.l�������>˲`?�|���=FMX�)�>�<�>����"����ֿ:�^�H��>	�?�Y�?!f��Y�� 2Q�ƕ�>�x�?G8h?�/�>��ym���g�>g"[?P�B?� �>j�mȾ��?CT�?�mz?�G>��?
�s?���>��w��/����˽��),W=H�	;e��>N��=ou¾8F�m���j��c�Vc\>��&=���>��׽R��̽=]������n�[����>h�u>/�C>���>;\�>\��>��>i=���{Y��A���S�K?u��?+��Ƨk�rñ<�?�=��_�&?|n2?��|�~�ξTO�>"8\?e_�?�Z?�~�>���3_��Į��֔���i�<��N>(b�>j��>���+G>l�Ҿt|E�ڋ�>���>ˊ���׾����V�W��>�"?���>���=�}?N�?�щ>[Ӄ>{nh�x����QQ���=F�>'i?Ozd??2�>O���Io��֓��������Ć='gr?bj(?ӯ>�鞿3��V����WH���L����?�?(����)J?ҍ'?>P?^�N?zl�>1��q���W޽��>@�!?�H���A��}&����;�?uE?�c�>4���ަн����q�ב��g:?M9\?��%?�����a�[�ľ���<�s/���X��[<�N��2>#;>輇��8�=b>���=+
m��C3���p</�=��>¹�=�H8�j吽�/?�/ռz���=j��D�a�{>nV>z����Dd?�N�W+w�wĮ��'��\;j�L�?��?�\�?�р��Pe�?�9?�Z�?'L?�J�>v���ʾ��۾+�e�g�[����y� >�(�>D*n<',㾪���Ƣ�����>%���p����>�Y�>
@?��>$N>爗>�v���[7�,!ﾔ��-:d����b2���8����'��.�Y��Ž�弾͗���d�>�V�����>�[?Po�=V��>:Ο>[�N<��W>�@f>/X>f�d>�+>�	3>*�=}�#��[i�W`R?ؕ��D�'�u��6����6B?�Zd?E�>�og��>�����H�?�c�?�G�?�u>@�h�u7+�a?r��>4K��Ȳ
?�9=��k�|<8����u��I��~�_��>W/ֽ�9��L���f�-�
?Zi?d���/;�I۽��i�#��=^1�?�+?0� �4UX�4%��b<N��<�g��=6��4V��5������3��Qqz�⢋��J:��Pv=?�@?6�t?,t���-߾F���0�f� "!��`>���>�&?�a�>��'>��L��O�}:�~��������>-�?�]�>)�\?T�?��m?�jV? ;�>�?�>ix��=��>Os-;A?�>���>ч*?&�Q?�-?�Z-?�9.?�@]>AO;�"y�Er����>��?r? I$??�(�:*����ݽg����<��G۽#��<�%����۽�Z<M�=5�5>�X?���V�8������k>�7?�~�>��>[��,����<��>3�
?2G�>�  ��|r� a�sY�>]��?S���=d�)>���=������Ӻ-]�=m���2�=��Ax;��l<��=���=�t�Z�����:���;'u�<s�?�6?(�n>�u>c�a�RS�,!��	�= 2A>:��>�=�=LVѾ5
������v�k��FP>�4�?V�?���=Mv�=O��=�������yK
�?#����=�M?�#?'CX?�E�?�6?N�+?H9>T8�{��B��������?��.?���>/���W���=��wiV�T��>`��>�8H���D�t��RU�7">�=T
��Z�X#���l]�{��#��H����?�ʤ?��=��C�K����4��KP]��"?���>�b�>���>Y.�]p�q��7%>57?��X?1$�>H�O?2,{?��[?�T>��8��%���ř�͏5�S�!>v@?��?��?Cy?̃�>>ǌ)���a��7w���΂��}W=�AZ>���>�A�>�֩>n�=�Iǽ#���?��|�=��b>I|�>y��>��>�w>���<��G?X��>F^�����ꤾ�Ń��=���u?���?��+?�N=�����E��G��nI�>!o�?���?�4*?h�S���=��ּgᶾ��q��$�>#ڹ>S2�>�Ɠ=7{F=�c>��>���>�'��`�pq8��WM���?%F?���=��ǿvOv�~6���������%�������t��|����;����˲��^����V������m������'���]����>@k�<; >f3�=u��<��i��`"=ܖX=ڿe<'��<�M^�'�=ݗG� ZH<��t�v��<+%�<4"S=�7��x˾�}?,)I?!�+?��C?�z>z�>�A3�4��>� ���D?��U>��O�[���P;��}�����ؾ?r׾x�c��ȟ��;>#7J�=�>4=3>��=�|�<P(�=��r=Yю=��W�r~=>��=�`�=Z�=��=�>]G>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>U8>:.>��R�ؕ1���]�k5c�eN[�P�!?sj;�J�˾���>���=u�޾�%ƾ�1=�E6>3�_= z��\�Oۙ=�{�J�<=]�l=���>y�C>H0�=Q����R�=%�I=7�=��O>��z��8�jv+�R�5=�k�="b>$�%>g��>��?a0?Xd?m7�>�n��Ͼ9?��"K�>Y�=!G�>X݅=ytB>���>j�7?�D?��K?>��>-��=~�>��>��,��m�hl�l˧����<��?9Ά?^Ѹ>!�Q< �A�U��g>��-Ž�v?�R1?k?��>7��Gl���/'���C��.z��?H=��T�Ծ�"����f���z���b=	@,><��>k�>-�>���='�%<n�>?v=�W>'=�s<
����]>2%\=���=���Jo¼t=5=����� �=�<��U<�߷=���;	;�����=���>X�`>XW�>��a��4�3F>>G>��5jO��Β=6ɾ��I��I�]�x<3�\�r����=F�	>�r�����,.�>��R>,�!>H�?jF�?���=[�O�����5]���8e������i:=ꑒ�4r5���F�uB��k¾$��>sm�>�$�>S �>ģ���!��>�f������?{Dg�s��=?w�s�T�ȇ��3¡�La��I=��c?���R4�>��b?}�V?�G[?�
?��"�Ϭ��a�">#վT��='پ_��e��K3?�!0?��>f�pY�X\���P�����>b]:��/N��P����0��:<�$���\�>Qž��ʾ�E2�"���
����B��Hy�HŪ>2_S?#��?��k�1V���P��;������?�e?;��>w�	?�N?q͑��ܾ���.�Y=V)Z?u��?r��?��Q>�2�=�����0�>�?HҖ?e�?�t?5�8�7��>�:(�Z�*>R���]�=��>���=S��= �?8�?�?�Y��`?���C��d�a�:�<�}�=�I�>X)�>C�`>�r�=��w=��=��J>3�>��>�C]>��>�l�>���Z���E?����|>�??��>��Ӽ
����ؼ��M�6=�O�gE�=\>��>76>V
U�<����?�ÿ^[�?,`D</���� ?^���^M7�Tj�>�ž>������4?#��<x�g>���>�.>��>�>{�>x���>ζ߾DM��+B�Rc[�֣;��>&��!���5�~���\�t���F�
�k�եz�?:����=��?����|�G 2��2�>��>K��>��5?޽r��伽�q>���>5��>P�z���~���dľE@�?vk�?a;c>��>S�W?$�?Œ1��3��uZ�߮u��(A�e�[�`��፿�����
� 
����_?��x?�xA?�J�<�9z> ��?��%��ӏ�C*�>g/�m';��A<=+�>�)����`�ծӾ�þ!9�vHF>^�o?%�?!Y?SV�"�`����>S�>�+?&Rr?�L^?a�C?TD���B?�d��ظ<?G�6>E.?l�1?!?E�>��>�hg>$���������e�����3���i���!�;������x�nV>�Ŝ�#��=��"��+=�j�A'�=A�P��8;pM>T�=m��>N�]?��>�҆>��7?
W��8�V���*L/?I�3=@
��Ɨ�������g�P�>k?��?aAZ?~�c>l�A��B�	Z>�.�>.'>�s[>��>t���jF�mτ=H>X>���=nM��끾��	��Q�����<�>o��>�5�>r��;�]>ܤо��Ͼ�)I>�I��躴��<	��K<�Qv1������>g�7?��	?y�?�Q��1<��So�� ?sM<?X�Z?��?�g�=����M�"�`yL�<y�]�W>��<�������_��U�C��y=��>؜���렾�1b>���/t޾��n� J�	�羭�L=+��d�U=����վ�:����=�)
>)����� ����qӪ�t/J?� j=C[���WU��s���>LØ>�Ϯ>�O:�_�v�_�@�8���)!�=!��>��:>ϊ������xG�9�t �>ӂE?;<_?[�?M ��h�s���D�H ��v����ږ�"	?q�>�?P:>l~�=�6��P`��e���D��A�>6Q�>MP��%H�?��������$�LK�>� ?A�>to?6T?1�?�:a?1�)?L�?Qג>i�ƽb����@&?舃?��=�Խ��T�j�8��F�D��>��)?w�B�Z��>�?.�?�&?��Q?ڱ?#�>ܯ ��@@����>�U�>�W��_���`>�J?���>�9Y?�Ӄ?��=>Q�5��袾�ߩ��]�=$>W�2?�5#?;�?���>;u(>��=�g�/HD>�d?L��?8�H?N�>cP?�oC���?%����%?��;?W?یk?x�U?7�.? K>��<��7��n�<Jx�������3=��=�V�=���=4+���ى�'�y�f4c<ZSټ���=��"=�C<Z���{]�1��>��t>�啾�]2>��ľ�Ɉ��@>����93��������9�Ș�=�\�>��?3��>3�#��)�=��>���>@�A(?�?G�?��;@�b��۾�K�8��>�rA?���=��l�_���iu�Z�c=	�m?�}^?�fX�+�����b?��]?�>�ڤ<���þq�a�e�F�O?��
?k�F�W�>�~?��q?v�>�de�X,n����L5b�)Xj��~�=翜>�:�^�d��5�>�k7?���>Bb>Ǟ�=�ܾd�w�0#��Z�?��?�?��?�*>��n��O�n��/����*h?�L�>ו��]+?:"�;��uhM�����jD��G����Ͼ�J����h�,B��m�(�-R��r�?��X?��z?��g?�����C��fg�S�n�� K����XY���/I��=�5�L���s��&�ǖ��ז�Ƃ]��%��N����9�?ܖ&?_��g?V�ɾv%�&���b�U=SC���� �jʽ�Ơ�B�8�D޵�F��ڙ��W"�+0/?���>�>{"D? #Y�*!��3j��<�rv�Y],>��>��@>5�?x��ON���l��Q���x����*�>�td?
�C??Wp?��罠�-����#�AE��q���"4>�^>�҇>DH����4"�N�<�1t�������-�Xn=-?��>Ԏ>���?6i?i��_��R�����1�x`:=�b�>��a?i��>!օ>SL���e(����>:�]?�"�>�Vq=΄��uE��(��]�����>
��>N?�^�>��r�<�>������8���f*��d���xb?��R�
$u�#��>^�&?٦��G�=Z)%?�,7�<F�����7 ��!KA��+?nG���B�W����X��o3�04���?�;?mc������5�>>B1?W}�>67�>��?h�+><����42��4?"4N?��Y?��U?ŭ�>?�<�UE�#|����7�=":L>:�(>-c�=�7P;���]H��������<��"��yý�L��[0<p�?;+�<7�Q=��=,mۿ�CK��پc�F�e>
��爾���yd�����c��Y��jYx���8�&�AV�5c�����Իl�5��??;�?�z���.������
���x���#��>�q�ف���������*�����ֿ�� d!�W�O��%i���e�P�'?�����ǿ򰡿�:ܾ2! ?�A ?6�y?��4�"���8�� >UC�<%-����뾭����οG�����^?���>��/��p��>٥�>�X>�Hq>����螾�1�<��?2�-?��>ʎr�1�ɿa���Y¤<���?/�@m�A?K�(�S��,�V=w��>0�	?��?>�Q1��6�P����L�>	5�?���?+�M=��W�}
��se?�2<��F����tE�=���=�@=���J>nO�>���OA�0ܽ2�4>Ӆ>��!�@���S^����<']>'aֽ�2��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=j���ƿQ_$������<��e��te�����3'��m{��`��S�l�*��6�=r!�=�|T>���>ѱO>�R>��W?��f?���>nK>���J��ɂʾ�����v���0�������������ݾ�$	������J ʾ+!=���=�6R�e���<� �K�b�]�F���.?ev$>x�ʾ��M��-<�pʾ￪�ڄ��ॽ�-̾�1�	"n�b͟?N�A?������V�[��W�'����W?HO�»��ꬾ���=l�����=�$�>8��=2�⾾ 3�u~S��p4?t~?y�ƾ;���S�>>�M	�V�g=^b*?=?�7=J�>��?.�3�qؽ'qK>N*>k�>���>�E >�ᮾ�˽k�?�eZ?��� ��9b�>�ľǁ]�%��=�>TA��o,<��|>=��<+�����P�Ѵ��xkS=�b?�f>-��@��!M�X���		>z�i?�i?��>��J?F3,?�1��׾�N���
�i�=��h?�Bv?�ѽ=�{�E������x?ſh?�Jc>	N��㸴��5���C⾻O?��z?�?�h=��:
��%���@?섌?��O�����tH���X<p�X>`R�>��*?�0�=x.=�9�>�Z?>Nm���hȿ[|,����?�@��@U/>�<�.�1<˩�>#?mO&�����N��W��aW>�t?[־f�|�zP�.>G�? "?c�>����p���Q�=�CӾ���?�f�?i�̾��=@�)�a]�����(Zɼs �=S1�d��V� �*�8�������a��'罏5�>��@����vb�>����w2ۿ�kȿ��~��}ҾX:8��
?�Z�>�c=z��=!n�����W_B���+�kAR��e�>�3>J��e����{���;�� ��A*�>u
�DY�>�xT�e��*��$+<$�>@K�>���>P鮽�R���љ?vE���[ο�ў�V���X?�f�?���?��??q:<iau��{���11G?�ls?#�Y?}E �s�\��=6���j?�S���"`��4��D�V�S>Z3?���>*�,���=�>۟�>�>�.��\Ŀ�������O�?$��?�o�	��>"y�?8,? ��>�������'�*���9��A?�2>n���� ���<����f%
?R
/?c��#a�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?���>�|?�S�=;�2?i�=Q �l�.�y �����=��=��?�XM?\'�>�i�=+��}!�=�E�V�J�E����"M� ;�>�a-?Y	?ȧ�>�#���. ����/��c<�`d���-�L�!�n[g=qb�=���>X�B>�٥��vi�j�?����Oؿ�җ���(��/2?(�>ђ?�:�@r�ɽ ���^?��>�S�OR������iR��o�?���?�i	?R�ؾ����@>���>���>�ս����1���20>t�B?��	�v���[Xp��6�>� �?��@u֮?w�h� �0?-���Ћ�n����i޾�>���;�>��?����r>���>�W�>4Zu�cX��䱀���>_�?.��?;�?ؗ_?�Rq��	;�
`�����>Ul�?x]�>��9=�Ȳ�������>%d������4�+��?��@��@��x?gl���ֿ�ޔ��־qϹ�l��<Q6�=��&>��.�^������_
c��R�=��>|��>T�f>�.B>o��=�b+=W����v!����A����{S��S&�������i+��Ν�˩���¾I9�z罬�<.GS��E~����"�$>-f?z?��?'?�3=c">�t��C�hS��ƽ�xz>�s>?c<P?LB&?>>���b�C��_���8���9���>�4>N��>K�>L��>ŉ$>��y>��$>廓>�>E�> ń=�t[>(k�>��>�<?���>�C<>��>Fϴ��1��k�h��
w�v̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��w�T�4:>9����j�5`>�+ �~l���)��%Q>wl?�f>!u>/�3�od8��P�{���j|>036?�綾*E9��u�<�H��_ݾwHM>�ž>0�C��j�E�����mui���{=x:?Y�?!4���᰾Ȱu��D���LR>X;\>�J=�`�=IWM>�cc�K�ƽ�H�Sj.=O��=��^>ט?��(>.��=�6�>�v��m�O�He�>i�A>��2>N#C?�#?������[Y��i�.�C�q>RZ�>@&�>��>�(L��4�='��>�m>fN-�t�`�I��r�C�z�Y>�Ca�1QY�Nj��?�=�ܙ��>`��=�U�I�X9=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ=v�>A��ػ��n���(ys���a���>��O?�p����Ƽ� 5�,t?H��>��򾎐��{�ƿ�j�sU�>���?�}�?��n��W��F����>m��?.�W?�@�>a�ھ�={� ��>VC?��O?��>�w�*��mO?'�?E��?��r>柋?e�[?��>!��\�E��ƿ���s�]=�=���>0��>ھt]8����`����`�23�O�>�ʜ=s��>���g��i� >LGr��ǆ��������>��8>��H>qj>@��>�	�>#4>�M����g<�o���K?Ѳ�?f��]
n�H:�<*��=�^�?�,4?M~[���ϾVԨ>|�\?C��?��Z?�[�>����:��x迿�����C�<H�K>�>�a�>�q���=K>��Ծ�rD��S�>���>/I��ھ=��]آ�YV�>�`!?��>�	�=B?CK3?F��>S�E>N|�碚��I��I:�>M>�>{�%?S�?6�G?������6��qz�HȤ��n��/#���q? �&?O��>�ԗ�q{��*W>xN��y����?
2<?L`��9?7��?���>�\?�w>��׽7��ま��>D�!?u���fA�h&����?iC?���>����Kֽ-Լ�1�P����?�D\?(~&?2���`��gþ��<,%�#C����;n�D���>�7>$����[�=N�>G�=9�n�g�7�ZPk<{�=E8�>�b�=s�5����|^@?�a�[���g �=�D��H=���>�*X>r���Lu?����k����7���Wy���w?a��?)�?�q=�[���3?�(�?"8?��>��r�R���ٹ��F���W<���y��=v��>��=�������3��*Ή����<b=��a�>?��>e?�	?���=J��>�[���^J��	о;��ޱQ�224�
D��D���s������=����`�I�>R㦽$��>�?`eP>re�>A�>�29=W�>Ip>�%v>Fۧ>�U>aP>��^>y��LR? �����'�V�辷����3B?-pd?�*�>��h�ʆ�������?B��?gq�?�?v>~h�-+�+l?�?�>���s
?\\:=7�N-�<bT������D��eT�G��>\:׽:��M��hf�8j
?/?V4��ɑ̾�s׽�蓾�MG�>b�?w|(?ޑo�CM(�����m�|���)�<H=6op��^��W;a���熿E/���!�������'1$?Ɗ�?��� ��	�N��-��P�>!��>o�>j{�>{�>+>��3��z& �K}�#�_�gqs>�D�?z8z>�N?t�?/U?�mR?�5�>��>��z�K��>0����>��>��A?(�&?T<?�$?�Q?��T>��D�'3��D�ܾ(��>��>�g?�H?r��>Z���0Ȼ�e<W�g#��;�'�'��<�O�++��(��W�=�M�>xO?�j�&�8�C���� k>�x7?;_�>���>����A(���
�<��>Z�
?@T�>�����lr��V��J�>���?O���[=�)>i��=l���DǺ�Z�=������=T���m;���<}n�= K�=��p����8�:-�;�(�<�� ?��?�ȇ>�2�>kh��N� �|��!�={�Z>`X>.�>�پDQ��z��v�g��#w>ݛ�?`״?uz=%<�=���=�Y���%��K���*����=V?]�#?��V?��?-"<?3�$?f >m&������ą��ʤ��{?�A,?�>�4���־%��ݔ7�6�?��>�Y�u������¾�2���2�=ћ<�
��<x��H�K�y�U=b�_=��e��?�r�?ma����-�?����^��eľ�E?X�>�|>���>�t.�,Vl�N�"-�=��?[�K?�>�>��O?��z?'e[?İS>��8��6��~���*6�di">MC@?���?�Î?��x?�/�>�>�)��ྦྷ"��D��Q�l΂���U=�IZ>�|�>�0�>,ĩ>Ľ�=t�ȽDr��h?�X��=Ub>��>v�>��>��w>��<c�G?+��>�\��ܕ�2䤾ݿ��A�<�$�u?Y��?ď+?D=˃���E��D���K�>�n�?d��?�3*?@�S�T��=��ּ�ݶ�`�q�#�>�ݹ>.�>���=ڄF=xq>F�>���>�-�\�n8��sM���?�F?���=��ƿ��s�5�{��Ԝ�ڌ<�/���j�]����m���R=$Ԝ�:��v��{�?��4��o���+M���W���.���,?,J=��>���=�P:�)��i��<��<��=3�=Ա����E=�iO�o�<}�x���ջ�H�<��-=p�k���˾��}?2I?Ě+?8�C?��y>�D>�X3���>�����=?�V>�&P��y���g;�囨�8����ؾ�y׾Bd��̟��9>2�I���>v63>oN�=}8�<+2�=��r=�ǎ=�RS�#=��={V�=�b�=��=�>�b>�6w?A�������4Q�7W�(�:?9�>�|�=�ƾZ@?��>>�2������yb�e-?5��?�T�?��?�ri�Xd�>���N⎽�v�=규�=2>��=��2����>��J>q��K��|���4�?p�@��??�ዿ��Ͽab/>�8>g>#�R�t1��]���c��\��y!?��:��˾b�>�=g�޾_=ƾ�-=}�4>D�`=6��!�[�oX�=�3|�#�:=�i=�܉>��C>��=$l��&��=�JG=׵�=��N>�P��^6�G0�H?1=���=W|b>B�%>Ey�>�?�F0?)Rd?�S�>�pm�k�ξs,��^E�>��=g*�>�M�=_�B>ۛ�>� 8?žD?��K?gq�>؄�='�>.��>x�,�f�m��C��|����<���?N��?Z��>�Y<g�A�!��eP>��1ĽGp?bA1?u?��>a{��˿'�6��B)���νUi˽q��s����9������4쑾Ca�g�F=�h�>m��>Vo�>�=���<�m�PK�>��=���=lB<�W<=��H=�����|��Ν�<L�.=������n>�5��c>/���Q#���S���|���<.+�=���>�P>S��>�z�= ���Z/>����L��r�=�N��oB�'.d�jD~�/��v6� hB>�*X>�Ń��0��|�?Y�Y>�?>�z�?'?u?}�>$2�^�վ?R���e��!S����=ޑ>2�<�7h;��W`���M�D�Ҿn�>	��>]�?�L�>t�(��HQ����>����x%>���8?�f;jn�<Nƍ���s�
˥�����܃��J=�.|?K�t�>��c?	Vq?�ҋ?�7�>�qνzݰ��@���F꾻���sF�����Lk�X��>ss!?F�j=ީ��:��Z��$=���>�1e�f�+�
���q־��=}	�|�>K:��l&��siW�wみ��eL:�5�^�z¤>Lb?�{�?�~\����ϓ���:�����9?���?�I?�Q�>e�9?q�<����p��P>;T-?�^�?�ʮ?L~7>ds�=^�Z�F�>S
?	�?��?�_j?G��dQ�>K��:[�5>
[���">�?(>�m�=	8 >�
?Ԥ?Ù ?���Q������9rj���<�*P=���>��>�uL>�>���=_��=��R>���>�ʜ>��h>V�> )�>���� C��?&"�߿�=��"?%Jg>>7������`~�O�D�n�{�2�>C�ؼ���={��<_9W�3�#�6�?��ʿ�U�?��>�	���(?�ɖ��Z���K�>�G`>�jt���>�ʻ>�}>�:>��C>��=��'>'�U<�Ӿ�>��0m!�9C�ՋR���ѾXz>s�����%�ml����mBI�xs���x��j��'���S=��C�<�:�?i���=�k���)�\��_�?��>k�5?�茾r��r3>��>��>[�����������gᾸ�?f��?�:c>��>@�W?��?��1��3��tZ�ޮu�]*A��e�Z�`�፿����Ř
������_?8�x?qxA?�o�<;z>���?��%�Yԏ��(�>�/�w&;�EL<=d,�>�'����`�Y�Ӿ�þH5�dIF>�o?�%�?�X?qTV������>�>��>9=?��?�Z)?`?�4�=��?.�>���>*��>�K?�%?ba?�ж>��7>�[]=؂��g̽������e�,��¼D�ռr��Z���V�s=
�<0��=V�㽛�==:��;�_&���2�K^=]��=�
>N��>|y]?���>S}�>A�7?j��7�
���.L/?P�;=���/⋾�᡾�r�t>�j?��?�3Z?�cc>�lA�TIB�H>;��>T�%>�9]>}Ұ>��տD��Q�=��> K>�ģ=m�I�JK��@�	�Z����6�<�Q>A��><p|>����(>Jh����y� �d>I6R�)���*�S���G�/�1��Cv��Q�>`�K?'�?!b�=Lp�ז��Df��.)?�F<?�-M?��?5��=;�۾��9��J�~w��ҟ>RB�<���n���%��~�:��L�:�{s>ߓ���q�]>H�ܾ�g�](��*oZ��	�]-p>������	��/���]��;�^>(h>�3꾔~*�����K���68?�2`�$�x��x����㚀=[d�>��>���������E��1˾p�>V�>j7>s�r;�����<F�wb�x�>v�H?�qh?>c?��y� 	���1��Ӿ (����>z.?��>�i�>���>;�<��4Q��#c�}�c��7�>��>Wk �
�O�W�ھ�&Ծ����ʸ>K�#?غ>��?�[?Ӂ$?��W?]GG?�?�h�>����TÝ��l/?��?��o=+RE��w��8�N��R��?���>�����>��?��?��J?��P?��?5��=���uoS�M�>��>�����M��']�=��c?��?*�J?W�~?� �=�"�2���1����e�4m>s�K?��#?�?���>v�>��]��	?��l?�i�?m�W?���=�O=?^�ƾ��>	��l�,?�$>�?��N?�y?��X?4?PG�<��<3��(��&�������K���γ�1^��U�νa`�=<��=��z�Wv(���ܼ�H�=�<�<�{G���>2x>���7�1>��������H9B>�-���K�������/����=0>�h?���>���=z��>t��>) ��'?�|?S�?�B���a��)۾�yF��ǲ>*OB?�<�=�3m�����u�xh=2n??H^?�{W�����_�n?�\?���j�p�_�4L���o�Ë`?��>�w5����>�Ef?�?��>��ݽ�r�$ ���`w�AAn�U� >��v>���"\J�(jb>/6�>kV�>-�>��;> ��8�5�����X.?T�?��?�ԛ?���>�~�\F��l	�`��<oT?��>Ω}�	?����g]�d���4����<��{���ܾqT�����[B����z�����="?Ձ?���?�U?"���T�X�4ec��s��Si��5���0����!sc�c�X�ŵy�7	X�������v�~��#u��9F���?�?Yx@�g��>��������8��`^>:VǾ �����ؽI�ۼ�M`�
�q�h�b��̾� ?&.�>��>e�7?�~U���;���,�M1�}���H>*@�>��>���>{'�����l���2�ž����νEVv>�yc?h�K?U�n?���\1��r���!��*7�k����nB>�U>w`�>#;V�j�iK&�A?>���r�^(�m�����	�eA�=�~2?d�>���>�)�? ?fe	�⮾^�v��0���<�n�>��h?�'�>%�>�nν�� ����>��l?���>��>떌�wZ!���{�ܧʽ &�>&�> ��>��o>B�,��#\��j��R����9�vu�=�h?���V�`�Y�>�R?�:_�G<�|�>~�v���!�����'�n�>]|?Ӗ�=`�;>�ž�$�v�{��7���})?��?~ɖ���'�+7�>xQ!?�L�>T��>x�?0��>8���~s�w�?��]?@�J?,�@?�g�>�WA=���}νPM%�,�4=k�>��[>�s=X,�=G1�F2Q�2��/�M=LJ�=`Sͼ5K��!'u<�����j6<#,=g�3>�ۿ�ZK�.�׾���C�
�K����-��s߇� s
��K���ř��+|�����C�ޢV�)�b������j�/!�?j�?ꏾ}���m@��1O�������>c�v�ϐ�������(�򭙾���ծ�$�@�P��j��e�c�'?O����ǿ簡��:ܾ! ?�A ?.�y?��!�"�|�8�O� >�B�<�+��s�뾍�����ο4�����^?x��>��0��{��>A��>͢X>Hq>����螾m-�<��?&�-?���>�r��ɿL������<���?$�@e�A?�j(�W���S=A��>L^	?�@>��0��Q�갾���>6&�?�֊?�M=vW��w��Se?�&<�F�u}��=y��=�e=���L>\��>�4��a@��ݽ�v6>eÅ>�� �~���1^��һ<5L\>0�н$���5Մ?({\��f���/��T��U>��T?+�>a:�=��,?S7H�`}Ͽ�\��*a?�0�?���?$�(?3ۿ��ؚ>��ܾ��M?bD6?���>�d&��t����=a6�P���y���&V�k��=Y��>\�>ʂ,�݋���O�J��N��=Z{���%¿�����$��<
ȼ����'��f4�+F��HJ���ܯ��$ད60=a~��Y>��s>$[>~`q>w�H?~e?��>)R�=��K����W���K��Q����G�6���ʩ����ҾV\���W��׏.��5��j�<�⩎=�,R������� ��b�ʜF�R/?�3$>��ʾs�M�f,</�ʾ�T���Ё� N���i̾3�1�%2n����?��A?w셿�V�������l����W?�M�����󬾨 �=㝬�y=��>�=�B�&3�1�S�KEA?�&9?L��5��<x�>KQ��>P%>�|?�X ?��=}=?��>����ے=���>���>)�D>-�?�p�=�9Ͼ��oj(?�(c?�ݽL[ ��$�=vIR�J>��J>%,>�ׯ�Hᔽʄ,>b�k="����=��=Lz�<��W?���>�+�E�������"�m�X=��w?�V?u_�>�$l?��B?��<|O���Q�N��I�}=ÆV?�:g?j>[����оB���g�7?W�f?W�D>~>l�(�徦
/�
|��f?��m?qC?'昼#L|���
�D56?��v?s^�ws�����=�V�m=�>�[�>���>��9��k�>�>?�#��G������xY4�%Þ?��@���?(�;<  �=��=�;?i\�>��O��>ƾ�z������I�q=�"�>���ev����R,�f�8?ܠ�?���>������:Z�=����%�?�x�?(a��]hG<F��Yl�����F��<qh�=��R;����c>9�8Ⱦ �
�w�����ļGr�>�(@��׽u�>�B;�q��=Ͽǅ�m�ѾĻp�y�?_έ>4�Խ>�����j�z�w���H�]�I����]�>��>:�M���{�֩=��k���>�,���>�K�	���;x��d�<�3�>���>�ŀ>��Ľj
þ䴙?���ο0i����ʢX?%�?��?�O!?��;��s��q���л�7D?o�t?��\?�����0Z�#�!�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?���>�?���=Po�><��=����U@�K�>�e�=��� �?]iK?��>�p�=4�=�΂/�h�E��jR��,
��rD�
��>�ab?�dL?fwi>������;��o �$�ܽ�Q'����G
7��A��eԽط,>�7>�>ڍ9���о��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*!rԿ����H�ܾH˾��>=k��=i]>�˽��%>=X��F署e�1̆>B�>n�>�{>ª�>[�>�Hr>�����(�*e���(��0�p���D�6BI�sѾ��%�}������Zl����K=�Ż�pr����Ic߽)�Ž�>�,X?7KY?
�`?��>�s@�5��=4����	�˺O��j=7j>D�?�W??�HO��S��L/d��@���dx���>�N>��>��>B#�>�Q�<�>��>ҁ�>��n>=c�;�\�=,�+:F�/>%z�>�� ?,�>ʣD>N�>v����K��.�i�9%��z6˽�y�?������I� ����O��%���~��=�i.?]3>�����
п����3G?]Ǖ�6$��!&�m >�/?��W?��>�����]�s�>���.�h��}�=�<��g�#�%�N>Z=?Z�>��>��%��N��'t�� ��Y'>�b?��1F�H�`�u|O�m�龄�>�Y�>庽\�$�ZM���V������4�=v];?&�?�N=�����ý�	�}��=�O�>�Q}�&S�=5\�>|��Y �.B��h�=���=!9>�f?�U>1?)=/`�>
%��*�A��*�>NL[>Z�O>[�>?�A3?����:���j�Q���M�>���>�ʏ>��=�Ga�g�=&�?j�>vi�^���C޽?�:��yi>����dx�򽧽j�s=k����/�=��=�݇�v6@��f=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾQh�>xx��Z�������u�p�#=R��>�8H?�V����O�e>��v
?�?�^�੤���ȿ5|v����>X�?���?g�m��A���@����>;��?�gY?soi>�g۾?`Z����>ѻ@?�R?�>�9�~�'���?�޶?֯�?�)I>~��?L�s?e]�>\zw��x/�c#��\���0yz=_�;nE�>�\>n���6F��ԓ��e����j����-�`>;,#=��>ס�|,��s�=�k���,����d����>�pq>�J>��>�� ?E��> ��>c={���j��������UL?à�?�'��Cn��<#��=hf[�ؾ?z3?Y�X��iξF�>x�[?l��?��Z?�Z�>�y�W��J����³�3�<�YH>v=�>�/�>�#2K>}�Ծ�E���>�7�>�~��p�پ� ����һ�)�>�J!?V_�>)1�=��+?��?��>�c=�aj��2����T���/>
�I>�4M?��B?�\)?��>�v��,���:��3/���(=�Z�?9-(?���>Y-��"����i=N����ŽM��?��9?I�־~�R?|T9?��>�i?I?'�&�`�׾au$���=�!?q����A�!a&���q?�:?�J�>N���3[ֽ��˼���a��X?E\?{&?&��@a�	Iþ���<?9(��^�;E<I�<��>/y>�+��ʴ=�>	��=��m���5�n�f<V��=r�>���=�u6���/=,?��G�}ۃ�2�=�r�5xD���>�IL>�����^?l=��{�����x���U��?���?Xk�?j��>�h��$=?�?b	?X"�>�J���}޾5�ྡPw�~x��w�H�>���>�l���F���˙���F��X�Žx�����>\��>��?%U ?�LK>���>�:����'��Y�Gz��9^�D�7�/�.�����٠���$�CA���¾-u{��ș>���� �>f�
?o�f>��{>���>S���K�>�pU>FF~>�
�>BW>��4>x�>�SA<?�Ͻ�LR?(���)�'�.��?����1B?qqd?�/�>Ui�C���)���?G��?�r�?=Cv>�{h�,+��o?#=�>b��Vp
?r[:=���3i�<vS��q��\-����殎>�5׽� :�UM�Jff��k
?�.?�;��ڃ̾�4׽HO�w�!��Զ?���>�n?�Y�C���9ɀ��u���>h=?��,�>(8y��������*������[���佦�=?Lx?u���R���"��DD��\��z2>/V�>�'?ْ�>�D�>�ӓ���<��~.�}a!�}���O�>��p?�e�>��^?Ҫ?�y�?�o@?�>n��>�v4��=?iWA=��>��>��?�d?A<?��?b/4?���> �T���������?�B?7�;?\�5?��?Ẏ�/�	��a���8L�����=�}��6��쮛��
<��<��m>�]?lS��8�8����&k>�x7?(��>���>���<���d�<h
�>��
?�L�>����Kcr��Y�Wd�>T��?�W�w�=O�)>,C�=���Cq˺���=g¼#��=:����:�G<<�}�=kG�=�7c��F����:
r�;:�< u�>6�?���>�C�>�@��-� �a��f�=�Y>;S>�>�Eپ�}���$��t�g��]y>�w�?�z�?׻f=��=��=}���U�����F������<�?@J#?(XT?`��?y�=?^j#?е>+�iM���^�������?nH2?��>���w�־���X L�̝�>"�?eMi��8̽
�3�m;[S���a>�I�(o��q���Z�mE���!����;R��?Jà?o(?>�%�n�Ͼ�E��R"��d`I?Õ�>�I�>�/�>3�v]u����T>:z?�|J?H!�>��O?�L{?*�[?�oT>��8�h�������M�8�">��??+��?�ǎ?�*y??��>��>�)�C�	���� �2	�T���_�U=�Y>���>���>?�>V��=��ƽP����e=��k�="c>~��>���>��>
�w>��<�T?Z}?���/���o��?
����= �r?�o?�K#?�m�=����7�~�ž<[�>ߠ?�a�?oa?m�k�Ë >�����۩:���>��?'�r>���<��<�<<�?��>��7���%��.4���4�F�?��]?t*+>��Ŀ'�r�_�_��ؚ���<:���Ӯs�����o1_�߳=�_���	�8ڭ�m�`��ޤ����볾)����}��@�>.@l=��>"�=t��<��Ap�< ==�T�<��=C�g�mT<�H�Ϗ���쉽�ӽ:b<��#=����b˾"�}?�!I?9�+?T�C?<+z>E�>DB0��ʖ>iH��J??�gU>+�O��g��$D;�-������h�ؾ�=׾y	d�N���1>�yK�&9>J^3>.�=��<$�=d�o=��=��G�s=@��=��=�Q�=p�=��>�C>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��><+F>�Ga��,�>���`�;s��#�?��:�kľg �>~�>�.ξ�������=�+^>�T�=Dh��fO�j�M=$=���� ��\�="��>�Q�>YV�8���>{�*��fn>�A>��y<��$x��kͤ<�Ԏ<aA�>��G>���>V�?4K0?4Jd?�>�>��m���ξ�4���Y�>���=�I�>��= �B>
��> �7?رD?��K?���>��=2�>���>��,�èm���Y���XS�<��?.ņ?�>6NT<��A����w_>�uLŽA�?�S1?�r?<�>���"�ۿg�/�T!��Jx�)@$��OL�����V�<������L��ԣ�#H>1K�>z;�>?,�>#I�>�>��>�S�>L>_��=�g>ܭ=���<#�I�a4�=�&�GU>�4=w��=�O7�= s�o�S�
��8�3R=��=e��=R��>�>>��>���=s	��~C/>⸖���L��ƿ=uG��,B��3d�{G~�3/�X6�ܵB>�7X>Ç��/4��U�?v�Y>eo?>{��?,Au?��>x!���վ�P���=e��QS�:Ƹ=��>@ =��z;�QY`�q�M��zҾL��>��>V�>��l>`�+��I?���v=�
�5�F�>���(>�o[�!�p�5��^��h��F�)D?E��Y|�=�*~?�I?;�?.��>����yؾ7/>.���R�=��Ӏq��R���?��&?��>#n뾴�D�_7̾F���>��>��I�s�O�m�����0��t'�k`����>x�����Ͼ�r3�?l�������B�ٟr�bc�>�SO?��?�Ac�*��cO�7��ި���8?4tg?՚�>�u?�*?����#=�j/��O�=ؐn?T��?�?x#
>rs�=r�=�s�>�6?�Z�?E]�?~@n?��B?�C�׽[>7)x�;/�>I.�<��>�>ut?"n?.�?�`ݽ�26���˾���Ɓ�� ���1�=��>�s�>�~>9���[+�$��<W*>tv�>�q>U	�=i=i�u>�ե����F�(?��=�w�>��1?��}>�Q= ·����<qmf�"�3�'!3�l����u�p<��ٻù<=�>�����>��ǿ>�?ojN>p�� �?�����y'��N>�V>�ݽ���>�VF>�:}>��>;�>^�>Ȉ>c#>�BӾF~>"��[c!��.C�{�R���Ѿ�pz>T���s�%����S��CII�~v���k�;j�/���<=���<�G�?���l�k���)�������?�]�>/6?�،�i�����>���>�ō>KI��6���Dȍ�kn���?1��?�;c>��>@�W?�?��1��3��uZ�+�u�d(A�/e�P�`��፿	�����
�s��0�_?�x?5yA?T�<":z>J��?��%�\ӏ��)�>�/�';�S@<=}+�>*��-�`���Ӿ��þ�7��HF>��o?9%�?nY?4TV�[.�X7@>H�!?{n;?xz?��:?<�H?	��4�+?�I��'�>D��>'B?�� ?��?�?>�>�2�==��=�E��ӟ���ս��ݽ�B���=��=���sJ_��H<�^ �X�O=>]W=ٰ�<�`���`<=7R�=�=���=q�>p+]?��>	�>�8?{!�7����(*/?�e$=��Չ�yN��\��6>Sk?���?�G[?�f>�A���B�C`>���>R�,>��e>}�><���VF�Q�=J>j�>�a�=�9^�A����F	�����5�<�I >���>q��>y�9�]�>s��f�����W>�LQ��D;�;�E}H��r0���k��$�>�A?�
?��C=!%���	�lSj��(?u�B?�-S?Յ�?ל�=xqؾ��@�((L�������>��G=����ך�:����;��<ך>鿏�U����*X>l�����N�y�P�C��k���2�����ۄ="���y׾_���sk�=+��=�
���,��+���⥿*%I?ފC=�⚾�);�󙾾��6>P��>��>`��Ec��7�<�nm���H�=zn�>֪9>���;���B/E��u�co�>ӂ2?�!k?��v?P��s�`�<+M�r������}$����?�{�>��>/w>PW�=���B��$t�v�/����>�\�>a��I-4�D�׾|�Q�=Q��0ܧ>R6?(߁>�n?�A+?'T)?�@w?FPB?J&?���>pH�d���V-?�?-��<�nU�<ʛ��6?����d�,?�f�>��� W�>�!?W?=�c?q8s?ʼ ?�%>Fw
�n�����c>y�>#�p�w��Jګ>GA?�Z�>o8?�ŋ?�V>U3�������h7*�X��>�V^?�?[�>�$�>�e�>�	�C��=#ѫ>GOY?�R�?A9�?���>�+?@�a?�et>�o'?a�?��.?�P?M[?�wS?]�?ᐦ=�潾k�=Y@�=�0�DaȽL)���=o⢼$5���]��67������͛��B�#���=gm=��i=��>�Br>^Q����1>f�þب�� �C>0m��~��|����9�Kٷ=!m�>�x?`4�>�"���=���>���>s����'?&?6F?�1��b�u�ھ�2M��>��B?r��=�]l��q���v��ok=VAn?��^?�kV�&���a?lU`?�Ǿ|�7�q@��̷����ھ��S?˺�>�'�̑�>p��?˱c?�?���c�l���Z�&`��m��="W�>�� ��ff�B�>Ǜ?���>Y�>O+�=`�о��c��̏���>�i�?���?9ǌ?�L)>�c[�P/�Z/�nJ���W_?��>zɾ~�?J] �:�޾hb���㒲�������������'��q���u��'�X�=T�)?3��?��?MH�?��(��s�Di`�-
��:�L���ž�3ݾÅG�<�\���M�<+��!�,�0OH�K�f�o=��p��)���?��T??�,��>����c%/�l�վsP�>L�}��]a���.<�"�1��k��=���/Ͼ�񛾥� ?Ӡ�>\�>K
>?q�W��u.�����(��Q�ց>��T>�a�>���>ɰ<W�s�pZ�*Ҿw6��_u@�A|>��U?�jI?��s?>��.��}���B�ǽ���x>:�>5K8>�\�ɵ/��)�5#E�= q�i|���ޅ���	��>W�-?�Nb>�\�>}N�?!��>ek
�۾�O�����Vǻ<��>xc?ӆ�>%lz>�A����k	?\o?D�ɻ�����K�=,\��6y�&�=�
�>�g;?Wc���ג�}��Atl�����F��1t=�R�>�3�?(_v�R\,��g�>�2?�"�9�.=KUi>�����о�呾*�='��>��>���=���>�>�������h��糾�Q)?��%?�_����>�"��>3�?�~0?��>t>�?]#�>�
��@��U�>�G?��Y?zlf?�%?\�t;�����7ݽ�kf��7���x>�>E�ļ��W>������E�����<�̅>�T�=^�U�����|�˽��=J�>P�3>*Qۿ,eK��ؾ�"��J�]�	��h��=���_ԇ�̿�+񴾷�� mx�w���m(��hU�,b�����l��g�?tI�?����+A��'Ě�ܐ��yJ���*�>��r�6}��򪾄���Z��,z�h%���!��P�d�i��2e�T�'?u����ǿ񰡿�:ܾ
! ?�A ?-�y?��(�"�Ȓ8�k� >1?�<�/��˝뾮����ο������^?���>���/��X��>⥂>)�X>�Hq>����螾6�<��?$�-? ��>��r��ɿY���k��<���?(�@�zA?v�(�P��M)V=���>�	?��?>�M1�E�S���T�>@;�?���?ϺM=q�W���	��}e?��<��F���ݻB�=�G�=
i=���v�J>S�>��(UA��'ܽn�4>�ۅ>�|"���*|^�վ<]>ɸս#��5Մ?*{\��f���/��T��U>��T? +�>^:�=��,?X7H�`}Ͽ�\��*a?�0�?���?&�(?8ۿ��ؚ>��ܾ��M?_D6?���>�d&��t���=r6�����|���&V����=[��>`�>Â,������O��I��V��=b����ǿ����0��ξ�/�=�𷽄�������,G�����M���?���=�P>'#�>�h�>jr>�9>�nW?bo?
�>̚7>@D.���Z���x�k��^����5�3��s,���Ѿ���B8����l%�w�5�u_���=�$G�=@4R�×���� �.�b�̚F���.?�h$>��ʾ��M�$�)<ŉʾŪ�jV��5��p0̾z�1�`n�Qȟ?�A?����%�V�b��;�������W?�+�t��Q���d�=,+��j=�+�>�y�=j��F3�VrS�e�.?l8?^"׾+Ϟ��V>f���J�>��(?}r?�`z����>��&?�3�Z3���r�>�e>�`�>5��>�!~=�����A��{?��[?��A���l�M>3�ɾQ푾�� �7��=ـ��I�D=4Fi>Z}=�N��)���O���H\�=|aW?���>�0)�ո�P?��E��vKW<��x?� ?�Ǔ>(
[?[�0?�����v�W��.���0=@�\?pak?|�>��V��1۾ ����G8?��Y?�:>�j��|׾�$��P
�"?ȹk?��? �۹X�w�k���_�|5?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?r�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������5R�=RY��#�?�ۆ?�����;,D�6�q��H���=^��=� ��?��������8���ž��V����䉼��>@ۻ��J�>������]�ȿ����iǾl�T���?���>S%Ƚ.Ǚ��Lg�D5r��WX�TfP��{���R�>3�>����Б���{�]j;�W������>�����>~~S�@,������@�4<�Ē>���>'��>�y���ս���?3E��3ο좞����0�X?�^�?�k�?�u?%r9<�$w�r�{����0G?ʅs?�Z?l�%��]�d�7���j?=S���U`�Ɛ4��AE��T>�3?�@�>Ð-�-}=�>�s�>5N>v$/�S�Ŀ�ٶ�T���5��?���?�l�)��>�~�?�p+? f��3��tS����*��M'�RAA?V2>ˇ��ݱ!��,=��ɒ�6�
?{0?!���*�Y�_? �a�N�p���-�B�ƽ�ۡ>��0��e\�M��I���Xe����@y����?J^�?g�?���� #�[6%?
�>}����8ǾL�<�>�(�>�)N>�H_���u>����:�'i	>���?�~�?Qj?���������U>�}?�[�>�&�?8|�=�>���=�派*֕�_)$>��=Vuy�t<?�[M?H��>hZ�=�-9�,1�g�E���Q�^;���A���>s�`?�I?�=`>CA��"-.��n��޽�V7����Y�6�2�K���w`<>W�8>�k>��L���Ծ��?Jp�8�ؿ j��p'��54?)��>�?����t�����;_?Hz�>�6� ,���%���B�`��?�G�?=�?��׾�R̼�><�>�I�><�Խ����Y�����7>/�B?Z��D��s�o�z�>���?	�@�ծ?gi��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*֧ٿ�棿����؊����=�<�=��/>�$n�>K>��B=el�����=��>�ň>�E>s�x>�+�>ب|>��C>�˂�.%�@Ԭ��b����L�۴�<������R��u���.� ���X*�[|�38ؽ�׺�<��a�t�\������=5�T?X�R?	�p?���>�l�S�>@��=P##����=�߆>1�1?��K?��)?{-�=�����ge�B��������d���J�>:XI>.��>��>��> 9��I>?>I9|>b>�3=V����=�P>t��>�x�>���>�C<>ّ>Cϴ��1��Z�h��
w�@̽1�?n���E�J��1���9��ɦ��Ji�=Rb.?.|>���?пg����2H?���|)� �+���>��0?�cW?�>�����T�8:>����j��_>�+ �%l���)��%Q>�l?g�f>7u>��3��d8���P��|��2l|>�36?�綾�H9�r�u��H��bݾ�HM>iž>~�C��j�����r� wi�o�{=+x:?�?�1���᰾'�u��C��.MR>U7\>�Q=�p�=�\M>{Yc�s�ƽ�H��\.=޹�=�^>}N?I�+>�f�=U�>�k��9P��W�>�A>T�+>�??%?�z��;���l��5�-��v>&��>װ�>�l>>-J���=z_�>��a>sG�P����k�F�?��*W>h�}�f`��t�ȡz=񱗽���=�}�=uJ ���<�6|%=�~?���(䈿��e���lD?T+?_ �=!�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��I��=}�>
׫>�ξ�L��?��Ž6Ǣ�Ȕ	�/)#�jS�?��?��/�Zʋ�<l��6>�^%?��Ӿ<i�>\t�nZ�����(�u���#=P��>v8H?�U��ļO�Q>�wt
?�?�_�۩����ȿ+|v����>3�?��?+�m�%A��*@�C��>ˢ�?igY?�ji>Of۾lWZ����>�@?�R?��>�8�ې'���?$޶?���?��a>���?�Za?]��>��*��Z9�Ĭ� �y���yϽs~>�!>q�۾ܧ3�pꉿ�=��+�d���$du>�A%=`\�>B�������&��=�Ip��ر� u��s�>_�>�T>�%�>��	?e:�>>��>��=�	�c��9����9J?~��?/��� n�rJ�=���=B��Q?�35?(�>=SC���n�>��J?���?�Zj?ʳ�>n]�H����轿󨬾��<��>��>?�>#^�=e��>+������Ж>4�>l��������@������>��'?Q<�>&2>b�&?�$?�[@>m�e>U!*�h��� H����>$�A>x�>\i`?y�>�N��>�3A���ޟ� 7�ZO�>B4t?��?Q�>p���� ���)�>I#��4�����?��?�f��t��=h�?-1�>lY?�]�>sg����!>�/�>�"?kw�dB�(�����m�?�??�}�>�H�c&����z����i����?�U^?N�)?����7m_�$[ʾߜ�<b-��0�fd;�����.>��,>U���T�=��>j��=��p�^T<�@.����=G�>� >})��&��6=,?U�G��ۃ���=`�r�SxD�	�>2JL>��|�^?�l=�$�{�����x���	U�� �?��?^k�??��#�h��$=?��?,	?�"�>K���}޾(��@Pw��}x��w���>���>�l�p�;���י���F����Ž������>�A�>jN?���>�N>��>���?]#�q ��M����Z�$���4��I-����~~����J�Uފ�C굾.+|�&��>_ށ���>?�>+{l>>�>U)�;�tg>btR>l;�>8��>�DK>c�?>��
>r#�;�|ԽU�Q?R\����'��羠��`�B?:5e?q%�>Za�����%�>?���?��?Y�w>	�g���*��S?���>��~�5�	?�[D=QH̻U�S<�������N����W�)��>c�ٽ��9��&M��g�ei
?p?Lt��˾��ҽ��>�)H�;�v�?>�N?Ɍ[������%��E��qӆ�S��@W	��?��,�3;���@��͵a�~q�05�pi}<!?Ȁ�?��;���(��3#=�!\�}�/��E�>���=�h�=�=?B2>z�1�}G�kU����g�P��=�%G?"Rp?w:�>#�4?kJ?-�;?�9U?A��>Y��>ё���?)�@�8��>K�?e6<?J(?]�<?�c$?/'?4�T>� '� �	�f2��1?v'?&W%?�/?wS�>�����%
��!&����b`�*��=��>)S�=�6������j�=췬>�?H�k�8�<4���p>��2?���>���>烎�V�n�͡J<c�>)�?�I�>� �P�s������>�?���%	=��,>�V�=
Fy�4m�;I�= Ӽ%)�=FUZ���-�<t<�1�=Ϋ�=Zܗ;��r�'�/;ߝ�"Ġ<�� ?q�?��>�"�>����S�n
���=�wT>%&J>t�>]�ۦ��B~��Kbi���d>Ca�?���?�L�=}v�=w��=gȥ������Z��?�����<��?'�#?_%U?���?A9?|.#?/V�=�A�E���~0��dC��]j?�!,?x��>~��7�ʾ𨿒�3�?�?�Z?�:a����x=)���¾gսͪ>�\/�90~�\���D��������ty����?���?uA�=�6�t�d���
Z���C?l!�>1X�>��>��)���g�y%�Z1;>���>�R?!H�>/>;?p�?%u?��<�?�B�����zʼ�/>8W:?�(k?��?�_?>R96>ӻ��e��:m����#���Z��AG=��t>ζ>�o�>R̞>�r�=CA��2uI�Y�,��l>u�W>l�>�d�>��>�}r>�G��QG?
��>�Ǿ���J�[p���`�s?���?8,?>TY=mX�w�B�x����>]��?K��?ϻ#?Yn����=��C跾�o�0�>�\�>���>��s=I�=[�>#��>���>���B���9��%�#0?�:E?4�=Ќſ�Lq�[�k�����X<̞���ze�q���Z�נ�=t-��J��hF���#\�
ՠ�u�������C���q{�Ȗ�>9l�=H)�=j2�=F��<���<l�K=���<4�=*{��p<�.1���ǻ�<����q<?I=?Z�m�¾�Zz?��F?��,?� B?bn`>��	>�5!�mӈ>Q࿽f?Y�`>�����Ķ�_4;��㳾�䙾�ھ; ξ?a������s>��K��D>.�2>��=<XQ<>�=�i)=��c=�<4)=��="��=L�=Q�=��=���=�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��8>fZ>��R�p�1�2[���d��\�ӛ!?�;��v̾ �>Ŗ�=�"ྰ�ƾC'=-4>}]=�a��|[��|�=Fy�66=��h=<�>�tC>3��=2���ܷ=P=���=��N>�be���9�)�(�2=1_�=d�a><&&>���>��?�`0?bUd?u3�>�n��Ͼ�9��PB�>��=.J�>B�=rpB>���>��7?��D?��K?C��>
��=�	�>W�>V�,�7�m�^g�wͧ��ͬ<���?�͆?�Ѹ>��Q<s�A�����a>�XŽ�w?7R1?�l?sܞ>.:��-�<k��%������Z<�P�I�l�s2>��Q���麼$��>�H�>A�>���>� ?�V�>}O�ݻ>��>>��U��.M�=�ֽ �z=S�����=�->-�����}p��ļq�M����3<?3&�9��=j��=���>;1>!��>���=n���!/>i����L�;��=�K��?-B�8d�(F~�
/��t6���B>_HX>fE��{0����?��Y>c?>Ձ�?�9u?Y�>�+�v�վ"N���Ve�]VS��и=þ>�<�9w;�Y`��M�uҾ���>�>,��>rl>��+��5?���t=���?C5��:�>������ �����3q��8��"����i�����m�D?s0�����=��}?��I?�̏?.��><L���ؾ�+0>e���'�=��ۃp�Ĺ���?�&?�a�>�śD�'�ʾ#��⢷>dH���O�>���`0�@�/f����>���v�о��3����ZX��
�B��q�oV�>�zO?穮?�]��_��]P���:q��:B?)*i?���>��?a;?�i�����M|���=�Bm?k(�?��?#�>�C�=��
�=�>�<?��?�b�?C�?��%�=�>�����G9>Q#J�>�W>��f>�*>��E>k�?)=?���>�,��V
�L ;q�����l����=�=h�\>%��>�f�>�R�=52�=��=#>�>�D�>��>r��>9��>�1�����:&&?d >���>��2?9�>�$@=9����'�<ѣ2�Z\;��$���:/ֽ�~�<�s��#6=�*Ӽ0�>D�ƿs�?XY>���լ?
���/C���R>�Y>�?��>�~H>�$z>���>���>>�>s]�>S/->�Ӿ�^>Š�m,!��>C�bdR�t�Ѿ�y>dƜ�T&����b���@JI�񋵾�~���i�#.��?@=�L��<�:�?�0��y�k���)�c���t?h�>�6?e+���X���>���>П�>��������Ѝ�Wᾝ�?���?��c>~<�>ОW?{i?v�1��3�vZ��hu�(0A��e��`��䍿7�����
��½Rb_?X�x?ݍA?w��<�\z>��?�%�}A��Ջ>�X/��P;���B=ɧ>����@kb�tIԾ	�þ�&���F>Ko?���?/|?)]U���l�j~>D6?�0?tu?�6?1�??���v%?�`>��?*
?@8?�1?�?V96>0��=����'=�ɉ�����'ȶ��Ұ��%7�� =��~=���ٽ�;,�P=_�t<� �(�W�]:�>M����<>&@=#�=��=�٦>��]?h��>WG�>�7?4#�,Z8�-����-/?Jy9=m���:���墾��>;�j?N�?;`Z?_Qd>��A�`C�t�><R�>�&>��[>�P�>6���~E���=�>|>Ey�=��M�������	�����)��<PS>��>�{>�⌽F(>t����y�w�d>F`R�#Ⱥ�=�S�<�G���1��Qv�5�>=�K?��?��=Z��k���3f��)?�:<?i3M?p�?4��=��۾��9���J��w���>
s�<���<���*����:�Q��:��s>�'���m��B�W>߹c��z��4����/��I��0`��g�ֺ�=o�{��fA�Eˁ���{=�������^�%����3����:?xyM��� ������_zn>pt�>C�>�H<s	V�܄W���N��}>��	?Q�>��;b��w�R������>��@?(o?�?d?���^��>'���,�����jp�=23?��>H-?mo>
y�=�ږ���U�A�J�V6�>�}�>�'�śN�w����s���-�v$�>�0�>��n>�?�>I��?��>r~.?��(?��>ʏ�>�:<A+���C&?���?��=��ԽP�T�Z�8��F���>2v)?��B�.��>D�?T�?;�&?bQ?թ?��>Y� �xB@�̓�>S^�>��W��^��J�_>��J?��>�3Y?Ӄ?��=>�x5�Ţ���ː�=<>��2?o1#?8�?���>�x�>V���B��>kxb?if�?��?t&�>*�j?���>GU;?��>���>��>h��>��l?a��?j��?ܞ?M=������>b�E���"���r>rc=?6���D�<7n�=�����떽~�н���F�]=֖S=%��<��='`�>��s>�	����0>��ľP��[�@>F����O���ڊ�:�:��߷=���>S�?髕>
W#���=嬼>1F�>5���5(?��?[?7";��b��ھ��K�r�>_	B?���=��l������u�|�g=��m?��^?k�W��#���`?B$X?���_�Y��������,���r?Ɇ>���=tj��4Qy?�["?H��>W۽�B`����:�4�a)����=��>�n>�_�6�>���>9$,?N�>�r>�33�q�b�����>fe�?�Ϊ?���?��=a�^wϿ���m6��dW?���>�yɾ��
?�p��+"׾�ƾ{o������׾����|��yy���V�k���u���g e=ж*? S�?�nt?�qe?�,��p���g��@��Ǘn��+�=	žb�\��oQ�|Z�����8!��:O���۾rB���o�:R2�-��? �)?C贾�}�>^�Ⱦ���0�y�->Ő��w�����=�3<O�V���<�2��𥚾�Ͼo{?%Ք>�]�>��J?��P���7�=0�n�+��%��#:�=ߦY>Ҁ>C��>��^=�D�d�!�s���愌��p��5s>�P^?_R?l?J"�4,��"��y"��������IvL>���=�ي>�D����h"��>?�L�t����᏾rK�Q�=`m3?�!�>@��>�|�?3�?����H|������+�.�e�<d]�>�)e?��>�e�>��ͽL�����>�r?j�=�� ��t����E��T��_�=˰m>	�?N�p��*>z����%������uǟ�$�7�`&�x0�?��,�L���5D�>F?533��[�>fϥ>(�=���F�d�ٽ󿾣/r>��?�I�>O	L>&NϾ(;-���C��þ+�)??"M��s�*��1}>ʋ!?ن�>O �>wǃ?ק�>:9þF4����?��^?g�J?�dA?qR�>��=�����	ɽ�&���2= ,�>�HW>]=��=~����[��L�4K=ꎹ=5iּ�v��MF�;y���E<���<E�3>��տ�D��ľ���BS�����_���i����������a{��"���iS`��ݽ�����6���*���\0_���?Z;�?�_ �_I;�Na��V������/j>ULǾ�O����'�����׾Zl��� ��!�$�y��zu�v�k�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >YC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾�1�<��?7�-?��>Ŏr�1�ɿc���q¤<���?0�@�xA?��(�ߋ��nV=��>��	?�?>�X1��R��Ѱ��$�>�9�?���?rM=!�W���
�Qpe?�<��F�ˢ޻��=�9�=5=����J>�S�>�P��8A�Uܽ��4>;ׅ>%,"�c��5^�'t�<m[]>�8ս�F��5Մ?+{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?:ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=�6�񉤻{���&V�{��=[��>b�>Â,������O��I��U��=����#��<`��)��Q���<�)@�Aϊ�6wʽ+�/�j咾��\�M�[���>�>	�D>W�>2My>�[>n,[?�x?U	�>|�=�����5�
\��\$�� ����;J�����?��Z��؂��𾸲�)���2�aM�-�5����=O�R��l��3����b�<QD�E�0?�1>�iþ�PO��h=a2ѾPU���8ǻշ����Ͼ�/�Hpn���??C?q����Q����l��%4�<�S?]����������E�=_
��nH<= �>v�=ڝ�ʔ6�kyS�-y0?	n?����kk��c&*>z� ��-=׮+?�r?dIR<�Ϊ>:%?r�*�!佡r[>0�3>罣>ER�>��>��A�۽1�?q�T?�����ΐ>������z���a=�<>��4���輢�[>�S�<����W�m���'��<��V?�l�>�O*��/�<ʍ�*�C��=.�x?*?N��>� i?N]A?f�U<͖���T��H�X[=��V?+Fj?�k>O���Ͼ�#��p�5?��e?�H>��h����--�X���Z?�.n?��?@�m��{�$ƒ�����4?��v?s^�ws�����H�V�g=�>�[�>���>��9��k�>�>?�#��G������xY4�%Þ?��@���?��;<��X��=�;?k\�>��O��>ƾ�z�������q=�"�>���~ev����	R,�f�8?ݠ�?���>������Q��=<l��� �?z��?�Ѳ��k	;P���k��c�i
<���=l聽"[��z�_:��ƾt������f���W�>��@u�̽��>��`���׼Ϳ���ھ"ag�̎?u�>�$ܽn����Tr���w�'MV�υM��o��ܲ>�
1>
ˌ�v��Cg���9���2}�>�YC��J�>���Il�6R��be=u$�>��>�YT>袽8!ɾnՔ?_�Ӿ$�Կ_�����*�<?"L�?}�t?�%?�����L���U��~ֽ$KO?$|?.p?
��u�����ܾj?�]��`U`�^�4��GE��U>T!3?�B�>ȓ-���|=9>���>,c>%/�n�Ŀ�ٶ�?������?ԉ�?(o꾺��>0��?�r+?hi��7���Z��=�*�7/��<A?�2>������!�	/=�Ғ���
?V~0?�}�M.�_�_?�a�X�p���-�_�ƽ�ۡ>��0��e\�pN��/���Xe����@y����?J^�?c�?��� #�V6%?�>G����8Ǿ��<���>�(�>*N>H_���u>����:��h	>���?�~�?Xj?������U>��}?Eѷ>b�?���=�>��=W��"���>���=�'Q��j?��L?���>���=N�3� �-�9�E�cR�~��?�C��n�>�8d?:�N?�Qc>z̿�q�>��!�Ƒν�m(�m���@�j�W5ݽK/>@�9>�>qQ?���ξ��?Lp�9�ؿ j�� p'��54?-��>�?����t�����;_?Oz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>D�Խ����\�����7>0�B?Y��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?pQo���i�B>��?"������L��f?�
@u@a�^?*�Cۿ���ו����ؾG�s= +�=2�c>E����=��=�(�<0�y�s>ya�>>ٍ>�q�>��$>�!>y�>(/���a*��v�������B��y���35��z�־�lǾ`�6��������]U�y�h��:޽�v%��d�5s��O>�O?5^j?V��?5��>���h�=>AV�d���Xν�cE>yl>N�:?�XE?�?��=����jlU���s���������^�?�9�>Tʉ>���>�5J>����Q7>w��>XLN>"�I>Sk�=��=�V~��ݠ=o5�>l��>��>`�G>�&>����꾰�́d��R}�<���0�?�霾O�I��̕��	��أ��q��=9�/?�>����8�οV��2�E?}j���*�d]���
>8?/?^�X?��!>�����͖���>��"��bL��c�=�hٽ�SZ���'���8>
�? �}>⢎>��#��k/�ۅS�l��u�u>Mo?�]ɾ3���,`�9sG��Ծ;n>���>�6?<� �q��e��J�k��}R<�A??Rt/�r����N��Qw���؈>��O>6*T<�b�=��V>�}F�=���E��P;��>�j�>-Q?��+>!�=�ڣ>7o��K
P��S�>T5B>4�+>+@?�%?}2������|���.�#�v>+�>��>�=>&6J����=�n�>b>O�8N��S�E�?�U�W>�1}��\_�y�t���x=(͗��;�=�ɓ=� ���<��g&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>�p��Y��|�� �u�w�#=���>U8H?�V��e�O�4>��u
?�?�d�3���|�ȿ�zv����>��?t��?��m�=?��]@�ր�>I��?�fY?�li>1k۾�_Z�U��>߻@?�	R?��>�7�\�'�p�?޶?k��?���>+��?ĀD?U�o>i|�=N�����\L���½㘨>>�ͽ%�e>��� v�Bŏ�0��H�Z�������>��X=�>�>\Q���3�5Z>	�C�h� ���>"�>>��s>�\>��?^n�>S��>L�&=nd��.�I��Ѵ�k*Z?땜?)o���o��(>�n=�K=�?�?�����پg�
>��2?�cY?Z�?�.�>���2��� Ŀr̜��û�>��>�L�>|;>R]W=�b>ª)�m���"=`��>y�<�����#��k���[�>q?�Dg>�C��?�7?��S=���>ǻ1��R��:�W����>��>A�>�#5?R��>�D��<p�<-�����J�]��}n>/�?�h? ��>U���`��=�?#:�vK��_�?�W?iv<��>�J?��X?�^�>�M>��=7%ؾinZ=k�>r�&?���/�O�`)�?�����>�?��>1�������b�����#���?�+b?��#?K���e� kؾ���<�!�<ތ޻D2�<��n:N>٣>�������=s��=1�=�P��<x����ٻ���=|��>
 �={P� 鲽0=,?{�G�}ۃ���=��r�>xD���>�IL>����^?yl=��{�����x��$	U�� �?���?Yk�?Y��>�h��$=?�?T	?l"�>�J���}޾7���Pw�~x��w�a�>���>��l���K���ٙ���F��b�Ž������>�n�>��?%��>ndD>�M�> �����3���ܾ�I�C�[�����v4���/�2�����8�L�)8d���mŃ��B�>ǳ＿͸>��?؂E>1�>؉�>ɔ*���k>FBn>�I�>�(�>}�w>�\>���=�}=+젽�LR?0�����'����9���/B?6pd?�6�>� i��������?p��?|r�?yGv>�{h�u-+�&j?H5�>���'s
?L":=3���n�<R��X���%�������>O0׽r$:�M��mf��l
?Z1?�	��Б̾@׽9!J�?`+=��y?�Ka?są��MC���n�HJa���!��|H���<��3np��.+�̕�.����e���ER���l���?x�?c�9��vB�y����c!վ�C>�T�>�?>q�>d��>Q.E���s���j���u��}��?�?�>�>�>F?�2g?��f?!�8?�q>q�>����^Y>���T�>ް/?��P?�^?�G#?��?�G?��=g{��1��6�\V%?�a?�=? ?AE�>gD�SO�K(ؽt�#=������=K�r>���.%����½�0p=�-m>W?1���j8�����1k>T7?6��>>��>8}���M���&�<KT�>�}
?�8�>�/ �<�r�JG�Z�>Q��?����T=��)>��=W�����U��/�=
��'T�=ܻn���9�"�)<s�= ��=�5�Vu׺��:^��;%��<�v�>"�?�>#:�>`.��ݟ �I���F�=,�X>�\S>�r>�پAw���'��`�g���x>�n�?�n�?�rg=u3�=�e�=:i��w?�����(ν�9]�<^�?#=#?�_T?u��?k�=?�h#?X�>���Q��`��7���m�?�E,?\k�>g*�ɾ�3����2���?�J�>�_����'�¤����ҽe�>��+���z��访d�D�����:�����r�?�֞?���k6�`�)l���諾gE?�d�>֤>�(�>��)�8�f�9	��]5>2��>N�R?���>��N?[�?�a?��<>�(�B�������j&���l>	e<?�B�?#9�?бj?���>0E>���O1Ծ��v�e��zǽ�G����;��|>Z�>K�>W��>a�<&��(
= ����=y�8>ȟ�>��>�%�>��`>1M_=��G?���>�^��\���椾����u�<��u?М�?V�+?��=����E�AC���J�>o�?���?�6*?E�S�k��=z�ּDᶾi�q��)�>Gڹ>�/�>iÓ=�EF=8\>�>���>63��a�7n8��*M��?�F?��=pſE�p��we��q����~;�q��vj��~����\�~�=aȘ���+>��}(V����tu������$퟾�x�U*�>�̂=���=���=/N�<�\���<3�B=��<Z3�<raz�{�n<�RG�P����x��=�ԻD�{<�J@=.��8�˾N�}?2>I?��+?��C?^�y>�9>� 4���>����@?�V>�nP�{����;�N����!��*�ؾmz׾T�c��ʟ�PQ>�@I���>_:3>�9�=�4�<��=Qs=���=��O�"=�3�=�A�=�V�=���=��>�S>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>s��=w�2�T��>��J>���K��B����4�?��@��??�ዿТϿ6a/>�h8>B<>��R��1�z1\���b��Y���!?�3;�d|̾qɅ>�ع=t�޾�(ƾ�2=��6>U$_=k��d\�6��=]6x���;=�Ml=��>�D>�J�=1䯽�=/F=�T�=d�N>J�<�Q9���'�V�6=	��=��a>�|%>8��>k�?5�6?`�e?B��>�*�0i��R�¾�z>���=2F�>Nǥ=�8n>T��>O�8?zB?i�F?[h�>�Z=MЭ>�x�>�m6��p�M�׾�����<�,�?eǊ?2��>	&����N�b�!��:�?��P?�K3?��?%Ӱ>|��܂ۿ���xpC�5�K����@�=��<f=b)��Iz�����[Jj>ԯ�>���>i��>�	�>;1�>~�o>��>�|>��N<�N�=v���{F�󼽕ϟ=�i��ũ��!�	<1 �<殣=�c=�c$�����=���=	u=���=��>=>���>z��=x���%/>b�����L���=�_���$B�,1d��L~�G/�z6��B>�*X>�X��0��
�?��Y>�?>���?mGu?I�>b.���վ�L��dSe�1S����=k�>��<�8;��T`�O�M�~Ҿi�>+ٓ>�%�>��Q>B&�<?�xi�<�J׾06�'��>�Ɯ�p�#��/��[u��d�������8e������#E?�j��~��=hM?�J?Չ�?��>�ޅ�YѾR�>����22v<�x�q�N�և�%?QH#?��>?�߾I��?̾���ٷ>DI��O����0�{��<̷�Ւ�>k ��<�о�&3��h��������B��Rr�q�>J�O?��?F4b��T��ySO���x��cp?�zg?��>mG?:?����o�Mj���~�=��n?ñ�?;�?"�
>���=�����9?t�? ��?9ܜ?Vf?�%�L7�> �
=�mR>|�2�f_�>?�>�/.>YD>>��	?6�	?�~�>Q��{*�Gn!��	������=���=���>���>�C�>}=y���e��M��{>��>v�>���>��>%��>Z�������P.?�4�=
�f>�p.?K�i>�j=A� ���<L�"���Y��_#�L��',��<*���H<<�Ra��.�>��Ŀ�'�?}*p>w����^?-���s׼���>��N>�=�x�>��F>��>Uͯ>���>I�>O:�>��9>%3Ӿr^>4��J;!�]IC��wR���Ѿ��y>����<J&�����%��[�I�"G���s�j�,.��N=�8V�<.?�?Z����k�n�)�Ė���?j�>��5?\����,��m>i��>Js�>�q��l���Hʍ��-��
�?���?7;c>N�>��W?E�?ܕ1�]3�"vZ���u�b(A��e��`��፿뜁�m�
������_?"�x?6xA?E�<�9z>��?��%��ҏ��)�>�/��&;�;<=!,�>�*����`��Ӿ�þ�7�yGF>֕o?&%�?3Y?�SV���a��Y>jy8?cg1?��u?�(5?[@<?�R�Ӎ#?�/->�`?
?4?X�.?��	?�A7>��=|��;��+=�ꔽ������߽2Ž��׼.�B=|ݜ=Ub�:��<
Y�<�1�<�������n����P�<�2=g�=��=�˦>H�]?�@�>w��>Թ7?����{8�$����.?�;=�+��MΊ�����O�A>��j?��?AZ?&�d>��A��C�c>q��>�k&>m�\>se�>O����E����=�>��>h��=��L�ċ��U�	�ї��%T�<O>�� ?lW�>R�սڧ$>>(���Y�|>� ��ۏ��@����8�7R#�>�^����>��M?V�?)5#=����<#���c�S�?�]?��i?E�{?�j�<g&�ҁK�kVB������>���<˓ھ����S���n%8�+������>�{V��s���Yj>^	��a��l�>�I�~�徣�=`���0=���N@Ҿj~���=��>^��:�!�eΖ�`��69H?9%o=�ר��MR�Jy���8>kƞ>|Q�>��8��N��@V@�q�����=�I�>8�D>F���s꾕�F�P<����>��D?~d?�J�?�}�0�p�EF�����f���8
��?ؗ�>WB?��">�$�=�꽾���
He�JC�_�>l)�>S���E�K(����񾸆�f��>�G?�1>��?<�L?:?yMb?A�'?�e?��>����'�þ�(?x��?݆'=5�%�8{J�l1C��'A�=n?�?�c*�Ĕ>j�&?�O?�*?�P?��?쐋=Uv�]�8�(�>ޏ�>�0\������ؐ>5�B?U��>�lR?�ׁ?���=�['�g���8���cy=ՆZ>�.?�c?m�?�4�>�^�>�ڪ��I�E9�=�	l?��?f��?h�O�Q�?���>�_k?�fm=�z7>��>#S:?�S?p�p?'��?�<*?�o�=W�l���R��o�==��h=Mf�=�d;�妏=�̯=��v= p���8���$�{G�=-><*��=U1�<X�>k�s>9	����0>�ľ�Q���@>�֢�(S���Ǌ�H�:��=�~�>~�?�>x.#�3h�=K��>:G�>����5(?��?�?f�!;Ԙb���ھ>�K��>�B?O�=��l�����x�u�)	h=��m?��^?��W�O���d?�ya?n��h7<�Pt�� f��r˾K�o?QpG>K�3�=�>!�l?�2?TA?�Q
�7Y��쌿�(f�����=y��>$T���W����>��$?��0?���>�s]=g���D����N�?��?��? .�?���=b�I��gڿ�d�a����H?|	?$�ʾ�*? :�Ѿ^�Y��>5��ݾ��Ѿ�/U����$ʾ���5�P�<OཹC>Պ?ف~?v`?��[?8��5�^��P��x�S��#��U�� A�IUV�H?��<_����.N̾\���ەb=>����Y��h�?�5F?� ���j?�W��
)�����ʖ>��������]�>��ν�ȽCQh>� ��1*�G�`���?�!�>�.�>�<?cpQ�i/�G1�K`0�¡��j�9>
��>"=E>89�>x�d��9��N��-������<d;� 5}>yQa?tzY?��_?:�ӽ�K.��ԅ�M�r)��X��&>�>>"f�>*X�����A�3�qR<��ns�� �*~���� �!�Y$(?��%>EF�>]��?�	?޹��J˻�L���V"0��/=���>��_?���>��>�����*�h��>�l?s�>���>����{x!��"|��/˽Q��>���>"4�>�'q>^.�	^\�H!������Y69����=�th?����L_a��]�>�R?��:ޣj<��>g�~�� ��q���$��7>�{?�ק=�?:>��ƾ��:�z��(���;)?�/?����*��`~>�."?s��>ݣ>i$�?e�>��¾ʠ����?�_?>[J?gLA?1W�>� =������ǽd�&��+=ˈ�>a�Z>|�n=��=���  \�N@�:�H=��=�ϼڨ���I<SP��	N<8\�<{^3>�dۿb:K�Z�پJ��F%�8
����4W��a��qD��O4���x������(���U�5�b�,����l� ��?�B�?�]���N������������๽>%�q�{c��6ǫ�W���n��f�ྸì��~!�1�O��	i�_�e�U�'?T����ǿ�����:ܾ�  ?�A ?H�y?��-�"���8�ծ >@�<�+��a�뾧���	�οI�����^?y��>��&0��7��>��>�X>�Hq>����螾�,�<��?�-?Ǡ�>�r��ɿJ���"��<���?!�@�|A?��(�����V=���>�	?#�?>�S1��I�]����R�>7<�?k��?�tM=��W��	��~e?�Z<��F�U�ݻ�=�=�=�K=��|�J>�T�>���PA��@ܽ��4>Lڅ>vv"���+�^�R}�<X�]> �ս�4��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�}��=[��>c�>,������O��I��U��=*q��㾿�IA�����V��;&D��h*O��\'���%>���=��ξk��ʸ<+�=Ny���^j>�s�>Z�^>:7&>�X?��0?ny�>�)�>������m���m=�� &�=Tޫ�z����-=X���f�x��	�Ǿ����$�����<�;��=
R�����| ���b�qF��)/?S�">��ʾĀM�I�U<�ʾ#���cz�ѳ����̾��1���m�:��?ҮA?+慿��V��s����/���pW?T��;
�ټ��;��=V��]
=���>lԣ=��)�2��<S���0?�?.ʾ�B횾�)2>A�����<,y.?K��>��6<�/�>}p(? �@�{T�o�c>b,>ۑ>�f�>��>�⮾DV�|O?�1S?���Qq��例>χ���~��Ǒs=�Z�=
A1�&�ټG)X>�I�<a���/���˽M�<N)W?�h�>��)�9l���0�*��:=y?��?��>�k?6�C?���<K��JS�PI��.k=�W?"�h?>è���о���x$6?�<e?!8O>�vg���辨�/������?�&n?��?������|�{)�� ��#6?��v?s^�xs�����N�V�g=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?��;<��[��=�;?l\�>��O��>ƾ�z������+�q=�"�>���ev����R,�f�8?ݠ�?���>������*�<xд�D7�??M�?J�޾w��=���<�d�N"о�>-u	>�[��1s��O��V���6�����Z���^i=�k�>��@�8��^2>��L�L�򿧈¿�X`���Gľ��;?��>y�	���ҾO�K���/�C�"/�:�׾(V�>/36>)!�<�"���Kr�K�7�����N�>@J���M>�A��@��Pz��z0{�-�>^��>�^>*Q
��z��ݙ�?��߾Cӿ:������݃L? ��?{�?j�?�b�1|������σ<�X?rIl?�l?q<��vn=���;�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?���>տ�?oj�=��>�
>Tƾ,Ɏ�m�G>�-�=��[�y��>9S?9s�>2&�=��DT+��Q���Q���,�@�j�y>L�e?�J?��_>�&�������� �����/��ɹ�0�2�M��R�׽ů6>9�I>�!>F����l˾��?Mp�9�ؿ j��"p'��54?/��>�?����t�����;_?Qz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>B�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*�mܿ_:�����}W׾�>>�J�=���=�J��j1M>�?>l]�=��߽�aD>W?�>5�>&p.>�!v>.2�>@/H>-������2���(��¥3���0��l�>4G��Z�����=&�@9ݾ�4��\�=P��2�����#� �ͩ�����=�uU?k�W?�bn?�&�>7l�	�E>�/��<o�����{;n)}>%�4?��<?q!?��<�ޛ���V��Z~������@�����>[G[>�c�>Tf�>Q?�>�[�O�N>YNa>�wQ>>\'>�#�=�z�<e.�t�>m�>��>���>�1>>�
>4������A.h�3y�3�ʽ� �?J��#�J�����<�������*�=N~.?��>�����Ͽ	Э�@�G?d����|�,�_z>>l0?oMW?��>���P�d�̯>:
���j�l% >r���j���)��7R>�?Bo�>���>��$�f�7��sG�ǔ˾��>�jE?���WBԾ�i�"=���Ӿ%�)>�? ?����*����T��	���g�9�)�<?��?��#E��И�ܺ��`>��+>K
����=��.>�W�fy��'N�ax>�&#>�^>r9?o<+>��=�>�h����O�b��>�NB>�4,>�@?O%?��/��n����-���w>�!�>��>u�>]�I���=�h�>Nb>��96��&����?�O�V>mU|�zr_�7�v�E�u=�m���%�=u%�=W���(�=��q&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>zx��Z�������u�p�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾>`Z����>һ@?�R?�>�9�~�'���?�޶?֯�?�FT>L�?��?�֣>��>�$�����@և��ͽ$1�Q->aA�>�&Ⱦ�er�9Bx��g��N'X���1��,�>��B=ǉ>-�ڽ����q_]<�=pt��( ҼZ�>�Ź=�9@>2Hb>��?K�>Q�t>�]T�cD?=Ya������9M??�?�9��e��7a��&t=���v�?�G?��# ܾ{�\>�(S?��v?f�`?�n�>�j�◘��+ȿ�]�����;��@>Ï�>���>�K��+;?>�������_>��>-B��/�Ѿ�+��#�:�z�>o#?\��>��=֣ ?a)?��>`4�>[:��ꚿxAL�<!�>Ӗ�>o(?��y?8�?����;��e��92����O��w>��W?��0?�6�>�Zu�Ѭ���=f܋�wN�T�?ܛ?��=T2�>~�?%�B?ݶ�?L��>��|�E��L����N>�q)?����qB�,�!�'�p�(��>��?�c?���_&��DZ���)�$;̾>d? �d?�k?#���f�0���j<e}n�0�M���;����0>�J=>�dl�=q� =eB�=`>���u.�P����.>�.�>���=v��˩��,=,?��G�ۃ���=��r�:xD���>�IL>����^?kl=��{�����x��)	U��?���?Xk�?H��<�h��$=?�?Q	?n"�> K���}޾5���Pw�~x��w�Y�>���>V�l���K���ؙ���F��l�Ž�1����>~��>�
?F�?|�A>3.�>���é'�̿�U+�_X������9���+����iC���2�]�弳¾��S��>ph�U�>3?ozP>5�c>m��>F��)>�nK>F��>��>�UG>b>w>���<ģ�ZLR?����Ž'�y��ƭ��_B?�gd?G�>ێi�\������T�?�~�?wq�?ARv> }h�c2+��b?�,�>����m
?Ӣ9=��ȝ�<dL�����K����#��>-׽_:��M�*}f�q
?�-?"V��s̾;?׽7*���=�K�?K�'?�(��*P��|p��vQ���M����~�E�뢾F�7�˂�b���K�����v�(�%�8�c=9�+?^��?�@ʾ�M��R-˾e�x�ձI�5b^>+�>��y>��>�Z�>��b�(�j�O���I��b�����>�yk?ꗎ>A�I???!�P?��D?;��>+�>�Y;m��>�1���ۅ>���>�9?Y�#?K*?��?| ?=R>��,�v�dwӾ�H!?"*?�&?���>�Y�>V㙾GA��ĭ6< +H�a;4�bf3��E�=���������l#V=w�>"�?P���8�G����3l>��4?��>y�>�����\����<ƫ�>th?�q�>8t��#0r� ��o�>���?�O�0��<�r)>ȁ�=Yi�#.ݺ#��=Xļ!�=xl��rx?��	�;�O�=I�=�mY�P��:iI�b�];��<�t�>=�?ד�>MD�>tC���� ����Bd�=/Y>S>�>7FپV~�� %���g��Zy>\w�?�z�?��f=<"�=���=�{���W��u���������<��?NI#?XT?�?��=?�i#?r�>^*��M��_��	��p�?&?�y�>^X���߾�����b@��Ծ>0]�>��p��aM���>�t!T��s��fU<Lp�]b�z"��{[�U���� �`��	��?��?4�0=�^׾���j��%�޽��*?�A�>%Vy>��?�N%�V&j�40��?�>���>.�h?>!�>��O?5G{?۞[?.�T>��8��0��oҙ�U+5��!>@? ��?��?�y?%k�>>$�)�G#�E�������k܂�]�V=��Y>&��>\�>��>7��=o	Ƚ@>����>��q�=�b>>��>��>�>��w>�V�<k�G?(��>]�����ꤾ�Ã���<��u?���?+?�d=����E��F��bK�>Co�?���?�4*?׹S���=��ּZᶾ��q��%�>@ڹ>2�>�˓=mF=�c>��>��>�(��`�3q8��PM�i�?eF?ƪ�=��ÿXȅ��W��O!���{��S�*�,��U	��a)��׃.>XԬ�}�>�V���.%���쾥	��1b����\�(��s?{��<6��="�t>dq��a�=	+�=�T=��@=պ_=�I-�e�a;\�����g�ǽWxw=�J�<u��<��=!���3�v?�ih?=�,?$F?�$D>�2<>&(��ӋH>��n����>60>�=#����NO�b���s�������־փd�-��(�>)۽5#>��>	D=�!5��4�=%�C>c� >���X:���s�=�sD<�0�=��<n�->��4>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>ĥ>\��>�N��{g�O���d��9�v�7�Q?�J�
����Ӂ>#��>��"�P���,>L.���¾=�V���2���=�����|=>�Y:��>`�>�ؓ=C���@��|����<�y�=������[X<�>50��T��=�B�=B��>
�?�b0?nVd?�6�>en��Ͼ]?���G�>��=�D�>��=�pB>R��>��7?��D?|�K?���><ĉ=	
�>a�>y�,�ĳm��o�̧�.Ҭ<#��?�͆?�и> �Q<�A����ze>��*Ž�w?�R1?�k?/��>�����F&���*��m��O�<�=�p��p2��ƞ��qz��>|��>w�>�ۤ>��x>�-5>'�P>�L�>�
>���<���=���� 0�<�����=��ż��=Z횼Ჳ�b/�;�%T������.<^H�;�Mq<�+<c��=���>?>��>\��=����C/>ǹ����L����=�H���+B��3d�I~��/��W6�ֵB>9X>����4��*�?�Y>[o?>���?
Au?��>�#���վ*Q���Ce��SS��ϸ=��>��<�#{;�Z`���M��xҾ ��>lƐ>�}�>�h>�p)���?��vN=�ྒD6�`��>萐�ĺ��Z�s�q��⣿������i���W�Q�C?㼇����=5�~?��J? /�?���>�\��ܾRx8>y+��p0*=@���j�١���^?ww"? y�>8�羽A�!�ɾ2X����>p�J���N�!E��h�1��2�H�g��>�V��f+ξ�!2��ʆ�QR����C���s��\�>G�N?Cn�?�h_��み��N����%t��f�?3�h?И�>na?�??[̨���]�w��=��o?,��?���?���=4O�=���ā�>IH	?@�?ᘑ?�8r?�A��v�>k\�;�� >F���<��=��>S)�=� �=��?��
?��
?b˘�ǭ	�a@ﾇ��D�_��=2��=�	�>�U�>��w>���=�R\=ٱ�=#�V>��>S�>��`>
�>�U�>m���Q�8��>ʦ�>eO:>:�2?O��a ;�ߪ>�ǖ=������;�~�=��+>u�ξ�d)>��<>Լ�j�=���>a���dz?�8>�޾n1?��R�2��<���,�> KY=#.
>��>�Ԁ>���>��>��8���=�]R>{,Ӿ��>|���^!��C���R�$�ѾYaz>������%�H��0���QrI�����\�cj�G.���I=� ��<s:�?������k���)�^w��Y�?�"�>N�5?��������>{��>8э>"W�������΍�����?^��?>6c>��>�W?��?�1��3��tZ���u�M&A��e�P�`��፿S���)�
�����_?��x?`wA?d��<e;z>9��?�%�ӏ��*�>�/��&;��5<=�&�>V+����`���ӾL�þ%9��GF>�o?�$�?�W?�WV��h���+>�b<?�1?�t?�l0?L�:?��d�"?�x'>?�j
?<C5?��-?�T	?��'>ӆ�=��*/=�唽�J���/˽��ϽX ڼ��.=��j=aG�N<�9=���<�������>K;Q�ż�Ο<�(=��=s��=���>��]?�P�>���>F�7?����t8��ˮ��(/?,�9=M�������Ģ��2�>��j?|��?IbZ?�[d>O�A�#
C�C%>�Y�>�|&>i\>`�>q��БE��=�I>�\>�ͥ=)ZM�*Ӂ���	��������<�7>���>ԛ�>�o��->�˦�9�w���y>��n�x��J���}C��0��g�	ֵ>ܯI?
)?uI�=\'ᾴ��}�d��?ѣE?4�S?/ւ?Uֳ=�ھ�TG�C18�͗��'�>1D�=dr��6�������s7���<6��>�UI�rZ��Ywg>��վ_���x�bJ����8Jw����Iah;�<��뾁氾6� >T�{=[վj�,�@�����o�B?����Yp�i�"��X���'>>�y�>�:�>��v��5%���J�Y�����=f��>�NT>���<��پq+H�
 �m"�>"BE?�m_?Y�?����J1s�
�B�	 ������ϼy[?�R�>�D?�eA>��=���|��;3e���F�eR�>a��>)8��lG�ԟ��I���#�5F�>׷?)� >Lq?>R?��
?�a?�7*?�-?�.�>�[��-8��3�!?䙋?Z:�=��F���ݽa�/�-�7�ǯ>�+!?�a��$�>Ԩ?�?tF?$�G?^� ?'~F>d���Q�d<�>�K>	k�G���;>F�?zL3?�C�?p�F?:�b>�Q0�������v��6S�� >U�?�PP?�f5?I�>
6�>q�ϾͲ˾oí>�l�?M�?F�i?V�>[9Q?nM�=���>��罿4�>66:?��?��?p?}?u,o?\�?�]&=�����<��=swʽ�W���L�����;W'�=$�;�^A>�>��<��-�w�;=�Y<�;�N�����\_�>��s>P����0>��ľBN����@>t���O��8ي��:�Hٷ=#��>��?(��>CW#����=^��>�I�>6���5(?�?�?�K";��b�M�ھ=�K��>�B?���=��l�I�����u���g=��m?�^?��W�R&����y?DC~?����b�"Ŭ�:������u?�*�>1�?=Dʕ=�o�?��=?E��>e?��&5x��R6�@f�G}�;��>v��D������>qV<?�=�>@ֻ>Ϟ�
w��;��z現�?9�?2j�?�g�?�->xl����T����6#S?1{�>Qj�����>*�y龅Y��D���h�&����&׾Q���r��G���?�v6��d��= S&?�+�?�4g?N?ZY�8o�Id��|���S�(�����g�C�	W�ѐ8��q~��6!��*������=.�A��|;����?��I?�_��rʹ>�(���U���	��=��ھ:������I�����}�=���6���B�5?��y>p�>a�8? ���$(��#�{��2�
���5>���>���>��?X�T�:}��ǽ���TQ��/{���#>.�D?0o?)�m?����^2��`n�0V�����1ɾ�l�>�!�i��^�����y6��yW�AD��{�<��1���&����>{�,?w��=aT�>ȍ�?�Z�>�{�#��ɟ������=(c�>`?��?���>��i�1eE�K��>Qfl?��>0i�>,e���"���|���w"�>��>/%?H�h>�U9�
\������t;����=sg?���R�^�˥�>�7Q?��8��r{<�3�>�~�gp!����%��$>�?�y�=��<>��ž�����}�{��,�?,��>��־�=9��F�>�oE?�h?V��>�o{?�ݭ>b�$��
?ґ;?��8?��J?m4�>z�>��!=pJ�t��gD?=��>|�>%9��ix<0s��9��ʽ�	X9���<�m�<�!�=ܲL���������CF=��0>�տSG�Sѿ���b𾌾�u���6����.���%��؋��e������l\@�z���3��l.�̇}��a��(�?���?B��O⋾��۪������>�>���Z����r�����V��V�վ������YMH�F�U���Y�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@u{A?�(�3�쾦BV=��>Ő	?��?>�Z1�?J������N�>�9�?���?̀M=-�W���	��}e?�.<�F�y]ݻ7�=�7�=�A=|����J>rY�>Rt�zVA�+ܽ�4>�Յ>uA"�����^�q:�<��]>��ս���1Մ?&{\��f���/��T��0U>��T?�*�>|:�=��,?R7H�_}Ͽ�\��*a?�0�?��?$�(?(ۿ��ؚ>��ܾ�M?bD6?���>�d&��t����=[7�m���v���&V�$��=V��>��>ق,�����O��I��5��=�O��.��������&O�z:���x��S#�,�ؽ Й�d��{�����Ž�
����=�P>K7�>	I>�'Q>��Q?��e?��>l�&>���!`��j��,�󋋾���_��K����ؾW����A�Y��������+OȾ��<��5�=�HR����Ĥ ���b�A�F�p!/?3i#>H~ʾ� N�	�><�jʾ.���mDs�������̾9�1�O9n�@��?��A?腿��V����G�������~W??����O ��)�= ����=rl�>샥=�⾋n3���S���-?�Y?B�žL!��O;>.���M�~=y�(??�S�<�+�>�t?]t�Q��u�_>m\@>R��>�E�>>N>=�������}?9sY?�uὈ���kʈ>n�þn�|��p=`�=<�H�V�����p>���;�	���:ټY���&�<�+W?g��>�)����^���[�S\<={�x?��??,�>�nk?Z�B?��<�����S�6��Nv=�W?�&i?��>jr��p%оË��X�5?Ϧe?��N>Xdh�,�龾�.��U�4?W�n?`o?F���f}�v������[6?��v?�r^�ts�����4�V�{=�>\�>���>��9��k�>�>?�#��G������oY4�#Þ?��@~��?��;< ����=�;?f\�>�O��>ƾ�z������
�q=�"�>���~ev�����Q,�a�8?נ�?���>������=��=���9�?���?L����ټ-h��Do�f�nt����= e��E�Ž�����<���˾�A
�Z,��0����>�R@�i��w��>>q�i�߿�˿�B����˾!M�� ?��>�?�W�� xt��J~��}[���N�྇�罣>�/>G�������Oz��C:�������>�}�'��>
GQ��M��������<�=�>Ú�>��>5.���#��P9�?����c/ο�������Z?�;�?A�?�?H�R<Cy�J!���n�0+E?Ör?!�X?8�<5U��J"�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�d�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�S�_?'�a�M�p���-�	�ƽ�ۡ>��0��e\�+M������Xe����@y����?B^�?b�?���� #�f6%?�>t����8Ǿ.	�<ƀ�>�(�>�)N>H_���u>����:�!i	>���?�~�?Hj?���������U>�}?�]�>�:�?M5�=%��>�J�=rڱ�J�k���!>Re�=J5N�@P?��M?!��>�H�=��6�Rj.��>F�o�R���D�C�ه>]ib?g[L?��d>�k��G�9�N$"���ýi�0�]�׼=��*��޽D�2>=>�>��B�*XѾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ya~����7����=��7?�0��z>���>��=�nv�ݻ��P�s����>�B�?�{�?	��>�l?��o�S�B�8�1=-M�>ٜk?�s?Fo���o�B>��?)������	L��f?�
@~u@f�^?"�aֿ$ě�5r��<_��Aۑ=�; :||4>!�6�HY >ѻB�xx=g�=9�2>���>}�r>��>��=}e\>�:[>H��q� �����蛒�O�C������F&�������n���Tm��� ~������W�����ま�s1��]���>��\?V�V?��c?-��>�u�8��<�����b=Ƹ{��;h=@T�>�.4?��??}%?�7�=`��>�k�+����!��C������>�_3>�6�> -�>��>0���q�j>��[>:9�>&�/>��[=5s:�����RxT>���>���>_��>��X>��F>(�����^Fa�h�u��������?�򮾝A�����`j�zr�����=*�8?/�>5�����ϿO��A??G��R�����?�=�J,?��U?o�>�f���Խ  >p�6�BV��2�=�ӽm+���gX
>H?�f�>vB�>��3��v>�I�H�����ԸT>Z,>?��̾�_c�@�v��;��Xľ�)>ފ�>�lZ=+��cԚ��섿�#}�S�g=��D?�?@�i�M��j��J���Q߆>��>�Z�=2]�=�n>��t��
�S�N!�=���=�AF>��?+0*>���=ڞ�>6Õ���D����>b:A>In.>��??��#?�5������聾��*�&Xy>�N�>�B�>�>ݡL��ٝ=�>�Fm>t�߼v��:�G�A��6T>�G��age��7���=Pރ����=CN�=�T���:��#=��~?���䈿��`���lD?Z+?= �=a�F<X�"�- ��I���?g�@�l�?_�	�{�V�L�?�@�?X��n��=}�>�׫>�ξДL���?�Ž�Ƣ��	�])#�lS�?��?'�/�ʋ�,l�76>�^%?@�Ӿ[j�>�r�5Z��0���u�I�#=���> 9H?�V���O��>�x
?2?a򾸩��y�ȿ0}v�)��>��?8��?��m��A��'@����>���?ggY?5mi>�c۾�cZ����>��@?N
R?�>�7�X�'�i�?�ݶ?®�?��F>�?��s?ӏ�>�ȴ���2��	��2|����4=wR���>���=^�оܐE��2��֡����o��e��Y>[�\=���>��˽\0��IST=I�]�"꛾��q��ۯ>��z>�$F>�q�>�! ?w��>B��>�Z	=�֛��ܓ��-���'S?���?��#���v=7�,�a�ľ��&?#��>��L����dY�>��G?��3?�B�?�q�>���E�����ÿ;ξ�~<��>)W+?���>�L@�_�=��)�Z�=�Z��Å�>�v���)=�w�`�V���S+�>B�!?y�>>I9=2�=?��<?,>y>�>�J:�M������ݵ?�?/>
bT?(U?��?<4�|
��'T���sĿG�����>�a�?�?�I�>|��,r��b>�R?>��'���o?.�P?Μ⾔��>�D�?)9??7?���>�������>�:=ױ@>��!?��
�	�A�,'����	?��?H�>�r��� ֽ�T�	������+�?#\?��&?�i�a`�m�¾t��<�pX�K����\<@E���>��>R2�����=��>@��=g�n�QQ3��r<�"�=B��>�^�=�U6�����!=,?[�G��ۃ�5�=N�r�xD��>�IL>�����^?Rl=��{�����x���U�� �?��?Rk�?���5�h��$=?�?�	?�"�>
K���}޾J���Pw�~x��w���>���>�l���I���Ι���F����ŽWV����>���>��?}*�>*�@>൪>����h,����v���[�����-���.�6��%᫾�cM����4���7��1�>�~"���>ar?�Tq>ew>߀�>��:Yg�>]|i>���>wS�>�I>>=A>%��=5>='濽KR??���`�'�M��Z����3B?�qd?�0�>i��������v?[��?�s�?@v>�}h�=++� o?@�>q��Cp
?�L:=0!�K:�<V��7��6��W�>��>�H׽� :�RM��of��j
?�/?�
����̾S>׽qӽ�=�3�?Ia?S�ql�dGP�Z�k�ˮ���G�=5�y�D.�^�6��]�
���T҂�� x���)�󋭽�7,?.{�?�2�����W�{�pz����?�[�>p	�>=e'?�#�>�G�=R@��m@�r^��R��zھ�Ⱥ>䗋?V��>J�H?��9?��M?wSL?�8�>�$�>*l��=��>i�<@̟>�
�>PG9?��,?��/?��?��+?!�d>��������ھcl?�u?c(?�� ?L�?n��⊽��$���⢼]z|�O_s�ߑ=�>�<��۽B����W=�T>��??���8�&����o>��7?��>9��>`����q�����<� �>Gi?Y�>�t����q�2S����>���?;���=Z<)>���=��L	�2q�=�U�� n�=�8��޶8��eT<�%�=�Q�=��ݹmd����;m�;�?�<�t�>I�?���>HC�>n@��� ����f�=ZY>�S>}>Fپ�}���$��C�g�^y>�w�?�z�?&�f=k�=���=�|��TU������������<ܣ?"J#?'XT?A��?<�=?\j#?�>�*�XM���^�������?m,?IԜ>ag��vʾ���� �3��?�*?�y_�z.��'�7ٻ� ���F>Q�&�Pzu�F���3LH��?"��bN����?Ê�?��i��$:�~��b.������ =?�>_��>.��>|�#��i�<���3>�`�>��R?��>��Z?h�z?a K?,o>P�?��ɯ�����Lo=��~=�A?Ҁ�?���?8�i?�r�>9[G>�.�֥��3����:��㽳����C��M'W>�d�>1?��>И=��2��D)��\N�fh:=�,M>7��>~��>�\�>B��>��J<�B?��?W.���f%��D}�"����=8s?�.�?�	?�=���O=���
���>��?I.�?�A?�
q����=�K�Pcվp���!E�>"
?J��>u�G>����A�@>�#�>�f>O5������$�$]���v?M.V?�JP>`�ɿ��|��w7�X�d�KC~������p>���� �A�>'ɹ��@X���S�fZ��tʧ�n������"Z�u佯�?yu�=Q��=Mؾ=�j���ǌ�~�E�E��<N��=Ej�=R�ռt�Ż���j�9�(�t%"=��=!N}=��<ǈ˾F�}?�;I?��+?m�C?�y>�7>_�3����>��x@?\V>˓P���;��������Ӷؾ�x׾��c�"ʟ�J>abI�3�>�83>TJ�=�/�<�=�!s=7Ŏ=��Q�#=�$�=PL�=Gh�=���=��>#V>�6w?U�������4Q��Z罧�:?�8�>v{�=��ƾn@?}�>>�2������zb��-?���?�T�?>�??ti��d�>R���㎽�q�=K����=2>v��=x�2�T��>��J>���K��*����4�?��@��??�ዿ͢Ͽ:a/>�E9>$m>6R��X2���Y��Z�Q�S�k�!?��:��c̾s��>�t�=]�޾y@Ⱦ��7=�9>��}=.V���[��[�=�F���C6=�	o=��>G>x��=�h���
�=�"X=y��=\K>U݄�U�,��:)�-&1=���=��d>�b(>���>QH?�00?"�c?�`�>�Xm�L�ξ���I0�>?e�=�^�>yJ�=�^B>3�>�7?��D?��K?���>{��=�ܺ>�`�>��,���m�#��Q��m�<�҈?n�?&ݸ>@@<o�C�S��}�>���Ľ�2?J�1?	�?�~�>���}�ſ��ܾCB���\�b(�Nn>|*[���=k,�=:F�- >w^�>mV�={0t>|j>�wc>*C>���>��>̵D>q $>��>z ��-�=2�Nh��$�N��L�=�&��ǲ�)������Od;+� =�@=����h���=B��>y*>��><��=x����R/>���@�L�ӿ=�H���/B�@/d�YB~��/��L6���B>�@X>wg���2��A�?-�Y>&�?>y��?�:u?��>� ���վ�P��Ue�XXS�ո=>�>�=�H|;�]Y`��M��xҾ���>���>^ߣ>��m>d,��	?�7�u=�⾃|5�Qp�>ػ���� �ړ���p��)��6ݟ�Ji�B�r���C?3$�����=�/~?H�I?8�?���>���OؾR�/>N����=إ��-p�N1����?�-'?QE�>��͹D�'P̾1��Y߷>�3I���O�����*�0��]��ͷ����>���о�$3��g�������B��<r��>l�O?��?�b�\T��CSO�Q���a��	g?/vg?}�>qH?H?	����p���d�=��n?���?I:�?��
>�>�S��wr�>I݌>��?���?7��?r\�.>�>TV<@��<�Ņ�Z?>$��=+C�=,g>/�?��?Mp�>�佖"�B���ļ�\��lef=R��=�h�>�1�>�|?>��<�	�=Ȩ�=ֹ�>,�|>��>ӊ�=!̲>���>/��Ԧ�&;?���=�ҕ>�t4?g�>T=������=�?���m�p��wl����;�=�U;��m=��{�_)�>��ſ�Z�?� �>"��o?���/�*�]�=>��1>�����>�R>Ӕ>��>���>�=�8�>��">�AӾ�t>����\!��.C���R�c�Ѿ�fz>����^&�ʡ��p���EI�i���i�Lj�<.���==��<�F�?6���]�k���)�{�����?V]�>�6?�݌���޹><��>w΍>�J��㏕�YǍ�_a�'�?"��?V;c>&�>��W?��?��1��3�fuZ���u��(A��e���`�8፿���Ȗ
�|��9�_?�x?�vA?��<�9z>\��?��%�я�-,�>@/�&;�)?<=�(�>�(��N�`�k�Ӿ+�þ�8��EF>A�o?�$�?+Z?eSV��rY��!>f8?��1? t?e�1?��:?���',&?Ѫ3>K
?��?��5?X�.?�#?��3>�=��q9�<=����)��;X̽�½uw���a-=Q�l=g������9�="y�<�ݤ�����P�:AX���b�<�4*=㞙=��=�>�^?���>> 67?���4�y��K-?f�)=����9@�� J�������>��j?�D�?�FY?7�`>� C�ThK�2�>�D�>�D#>|�a>2K�>	�EVC�SE�=ǹ	>v=>׌�=��7��F����]F��<}�<"�#>K��>vp�>.��\n>?ܚ��z��c57>xf=��%�������uC��;)���P��M�>}�N?ϩ?l�=o��K��κe���"?IH?T�S?��?
�<E��%�J� Y/���)��.�>6�O=������D�����;�F� ��Ђ>�-��v����_>��ľ���]ۀ�s 6�U�ؾ��ͼ/J�dZJ=�E��e@�񼥾��>��=������4�}���Y���JB<??z�<K^��FF��j���r�=!T�>�#�>�������\A�dq���p=���>l�>�3�;��OX5����?&�>��C?��a?��?H����_m��rA�����"������X?Si�>�?�A>��g=�H��WL�/�g��B�_M�>?u�>M����A�mӥ�)
߾��� �>t*?oz>U?C9I?(z?��^?�)(??֧�>�Ž����< ?�Ç?���=�n��}���h��]H;����>�y�>p���lR>t�?�,!?� ?�S?�?�
�>z0�L;Q���>ًa>��d����X\=\;?�U&?���?��s?
 ��Q5�y7�ݞ%��*}>�*�>��B?�� ?P��>+_>s��>�p�vyb���>��c?zߕ?��?� ;d�K?�M+=8?����ڽ�>�u(?�3?.�?���?4�b?�.�>�In<�0
��5ڽF�"���<A�.=72V;.�c=r`�U�H��=`
��\�Ὣ��=�Ɓ��܀=R�=�+�=�^>-��>o�y>����->�;��L��f�7>R��� ���ˇ��(F�T��=���>�' ?��>�&�
�=í�>�Y�>S��&(?{P?��?�e�;Na�p�ھN>P�F@�>sjB?���=B�k�����u��@t=�/l?m�^?]Y�����:�l?�P?R'���^�[rd�{B����	�~�V?���>�(a��+G=4{�?�bg?Jl�>����fz�����M8��>
���|�O(�>�o����4�|D�>�3?͚;>5`�=+�$��"�s�<�ģ⾹H?��?hu�?Q�?��=��l�5ֿ���-��rtW?���>�;���t?ǜ���޾�ʧ��狾:C���@��d����醾�K��]OZ�Co�$���%>�*?�ņ?Gˀ?��^?{@�hOr�jb�P%o��r�����'U�Y7:��\P��Ea�k���89�� �I��CV�=�u���=�u�?K�)?B�L�0��>̘��-Y���LӾ�z?>�C����!�g�h=7�f���=�sX=�{�C��#�� �?�g�>L-�>g9?�!W�'�<���.�T�3�q���%>�:�>��>E�>�lٷ�,���ڽZ˾瘀�^L޽�~>��M?��_?�P|?�込i��f�`l-�1��5�-�z��>#�	�W�>�2������#Q%��vT�+,��XP��=��e��>s?5 ��Dk?yU�?�>�Y�����$����_��#���>�d?d�$?o�=A$���>�D[�>�l?���>ͤ>�J���$�"�{�; ۽(��>��>�P?nPc>�6+��[�R%���z���E:�!��=��h?'z��Y�>��>(�R?�l�T�<4�>.�d�0� �Id�=�!���=��?N�=e'/>���I����z�
Ր��&?}�?\��qL0��y>�#?��>i�>M��?�ц>�/Ǿ�3����?{Y?Z8P?+A?�i�>+�7=�.�n��Յ?�B�t=�e�>�Q>��=�v�=��"���>��L�5�m=�7�=����;��g������K�����=:>��ѿ��C�V"ξG��D�a�	�ji�����+��"Z���ˍ�㓾�_)���� �q�A@���"�S�����;�?5A�?����W�.񧿕*���|���>�ӾP�ýbt��!愽bhʾ~"��'�S�O���F�x1o��n>�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >[C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾w1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@:rA?��(���쾍�T=���>pt	?�?>9{1�v3����y��>;�?��?�<K=Z�W�IJ�~oe?0a�;z�F��p�=���=�==���pJ>�,�>��\A��V۽\�4>�>71#���:^�]1�<^�]>z ֽ
��5Մ?+{\��f���/��T��U>��T? +�>U:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=}6Ἓ���z���&V�x��=Z��>b�>,������O��I��S��=fl���z¿�U&�M��#:w=$�;~S5���)��1/�)i��}Yk�T܂�?I�֏6>A�>��x>�a~>��Q>��m>E�]?e^t?���>�j>T<A�����&��پ�yf����0Ì�_��]��)+���!ؾۡ�i,�*��@Z��I=��E�=A3R����� ��b���F�B�.?�h$><�ʾ��M�] /<�aʾ翪��e���ϥ��̾k�1�r!n��ȟ?o�A?����b�V� �n%�L*���W?F�¿��R�=,籼�#=�7�>!��=��3�_�S�G/?�l!?�a��Ɨ��4>ҿ�����<�/)?�!�>�6�<�m�>4Z%?Nb��v��Q?c>�)>s
�>�A�>���=����{ѽ�� ?��Q?�������.�>�¾��p�o�=��>��;������M>QB�<?���䬻L���g,<1|o?��J>��I���1u������$��Zڒ?��/?X�?�!?�,k?H�<�|sR��0m��=�.LV=l�[?[|�?|��=[֗<峇���1���??4�W?u�=l��a%�Ļ���G���O?�.�?Fv?��ļ��O�刿8-)���>��v?s^�xs�����M�V�b=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�$Þ?��@���?��;<��R��=�;?j\�>��O��>ƾ�z������5�q=�"�>���}ev����R,�f�8?ܠ�?���>���������=�E��Iū?�=�?臬�j�c;���H�k�2p�<��<�ѳ=f����(���f�7�q=ʾ��	��v��F�h��@�>RE@@�˽�d�>|�E�����fο�&���}׾�>n��X?���>�.ٽ����T�n��{x�fK���I�������>
�+>z������p���3�p���K�>�fB�T't>r�P�Cm��G=��G�C�\�>!j�>`��>Şܽx]ƾo��?�����Qο���#'
�sV?���?_�?\ ?����8������2�μ�I?�x?��]?6V����q�&���@�j?�^���U`�S�4��GE��U>�!3?C�>'�-�#�|=x>��>mh>�#/�8�Ŀwٶ�x�����?���?�o����>��?�s+?bi��7���[����*�4�+�<A?�2>&���`�!�v/=�.В�4�
?~0?�|��.���_?��a���p�W�-���ƽbܡ>̿0��c\�'@����^Xe����e?y�s��?$^�?K�?'��c #�F5%?�>>����8Ǿn)�<���>�(�>�*N>�W_�Ĳu>U��:��i	>���?p~�?qi?���������U>2�}?��>a�?�0�<(+�>��>�@��-����ܮ=:a�=��>�l<�c?L�*?�0Q��f���&��c�qC��h��,O��Ю>�qv?$X5?V�>�ڼgg���7���B��oƼ{⼹�k�%U�<0eL�y��>�M><��>�֌�2����?Lp�9�ؿ�i�� p'��54?-��>�?��{�t�����;_?Jz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>>�>�I�>=�Խ����Y�����7>0�B?U��D��t�o�z�>���?
�@�ծ?hi��	?���P��Sa~����7�]��=��7?�0�'�z>���>��=�nv�޻��Y�s����>�B�?�{�?��>!�l?��o�R�B���1=;M�>ʜk?�s?*Oo���n�B>��? ������L��f?
�
@u@`�^?)�t޿+k��t����ő>�$�=,��>�\���=����?=��+��U1�>u��> �>ѭh>Hł>J`>��� �=?�������)�=v��V��g+�-�
�����[l�^M���ླ��qs�	v�"���y��L<�����=jiZ?�S?�_?@�?���W��=Pc�^�k<	�ҽt$�;���>��3?��6?�B$?�<=aٌ�u�c�t��)��7�{���>�@>���>���>@��>( �J�(>�5	>��>]g�=X�<IE{�AE=b�k>{�>���>ݏ�>zE<>B�>~δ�]2��4�h�]w�Q̽��?����J��1���8��'���ck�=ec.?ށ>���>п����,1H?B���0)�a�+�9�>��0?�eW?%�>�����T��4>���ĩj��d>! ��{l��)��'Q>3i?�Dg>E�y>��1���8���O�5����~>Y6?�r��qg?�PWu��PH��lܾ�M>v��>� �Jo�le��*7����k���l=M�:?	�?����
Ǯ��.o����1W>�\>|�=��=��J>��f��;ǽ��H��%=[�=��\>�?�R/>:��=ߧ�>䳜��M��E�>\�9>ؾ$>��??��"?���昽T��oX/�4s>�n�>Dv>�� >�DK�PR�=���>��]>�b�>������h�?�4~U>{M~�l�_���m�65a=���#�=ƨ�=9� ���;��=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾMk�>w�VZ�����	�u��#=K��>�9H?yS��T�O��>�Ez
?�?�a������ȿT{v���>��?`��?��m�1@���@�؂�>W��?�cY?9hi>�m۾geZ�r��>	�@?�R?l �>�7��'�1�?ݶ?���?�lP>3��?�?z?���>^U�@�$�H��Ҵ��I��;*7<���>W��=L̾o8��⏿��F o��� �t�/>FE=�>\������$��=�_���"���+�Գ>��:>��9>�7�>F��>a��>�7�>�J=����%6l��W��A�=?]��?>���W�����=��>���$?��?��6���� ��>>|N?|oe?F�p?��>�ڧ�s˔�A�ƿhKǾme�ٲ�>O�>�>�����$�>NK��4;D�Ӓ�>���>�D&�o�쾔�a� +�=O.x>�?� ?v�D�9�1?�2?���=,��>�7�uז�&�>�b�?R"?ђ0?z�a?R�?�>�C�K�P8������@H����>��?�`?�^S>����j֋�ʌ#>�k��?�����?gVu?h7.=�1?�j�?��=?I`?�p>�F5������-��ݡ>��!?�	��@A��p'�]���u?�?�P�>'Z��-�㽫=��`�~�����?��\?r�&?�����a���ž�h�<Q$�f���q'�;~���zr>\�!>��~��=�=x�>$��=��r�˃8��<,��=���>Ä�=�3��ϙ�3=,?��G��ۃ���=��r�ExD���>�IL>����^?dl=��{�����x��+	U�� �?���?[k�?'��;�h��$=?�?M	?s"�>K���}޾/�ྐྵPw�~x��w�q�>���>#�l���I���֙���F��Q�Ž"�ӽ--�>f6?�?���>�P>	��>V<���51�S���n��Ia��)���>1�Q��u��h}���׽����_��2�>�@x�
�>��>��0>���>Q��>wIȽ�Q>x�0> W>מ�>��'>Ҍ'>�-�=�^!=�ز��OR?Z�����'�������B?�Td?�=�>r`i��~�����?i��?xh�?�v>�h�"-+� g?y3�>8&���z
?�S:=��	��ǈ<�F��8��㋇�����>��ֽc+:���L��=f�{
?%<?+*��ۜ̾�׽�C��[�=�J�?LcB?/�X�x�9�L�Y���9���O��?(�ˏ�ܭ���6��5�Or���Ku�qX��$�(�_��=�7?��p?�|�����Xt��=��j���>M��>��	?���>ب>��X�M�P�g�Ӝ3�q�u��o!?*{?��r>�>?)0?�&?��;?���> ��>{D���?0�X��R>���>�4?�"?/�F?�� ?�w/?]��>P'��
�	��x'����>*SM?w(?�q�>�?�m��r-��̉<�v�=��0�QQ>I*
>���� �!�B�-�='Զ>�X?����8������k>8�7?��>h��>����,�����<��>.�
?�F�>@ �(~r��b�uV�>���?���W�=�)>���=������Һ.Y�=,����='6��+w;��\<v��=���=)t��B��8�:��;�h�<���>��?r��>���>Z0��{� �_���_�=�)Z>5NT>0>��ؾP����2����g��Px>Vd�?�?@1k=Q(�=f��=�����e��,��/`��R�<!�?�>#?AKT?�y�?Y�=?0�#?�>���3=���2���N��ץ?=!,?Ҋ�>���/�ʾ��#�3�ќ?uZ?4<a�=���;)�P�¾� ս��>�[/��.~�����D� @��C���~�����?S��?�A���6��x�-���vY����C?:!�>X�>�>�)���g�2%��1;>��>R?��>��Z?��~?M\@?M��>�(�ζ��@Ŝ���f�=i?>�)?zƀ?o��?�L?ȭ�>O�=?˽��VC���j�5C~���Gd,>�>���>eͷ>�RC=�U{�O�o=/�=���8=��]>��>���>
��>�1L>+�;�G?S�>�%�����4��t�7���u?���?��*?k�=)����E�8���W�>Y�?���?)*?N=V�k��=r߼�-��]�o�ʵ�>��><��>Jm�=��J=��>��>O��> �4?��X8�9�M�R�?�iF?ѻ=UĿ��o���a�H����c�����!d�����2b�=�=ҳ��{�
ꭾ�>T�����>��Մ��8��:��/�>T�=��=ص�=���<���:�<[=��<zL�<�+}���W<�;;��>ǻJ����}:�:1<.U=��L�Ǿ3+~?��I?��(?�wC?$gs>��>�i�č�>��[�vs?�T\>�*�޼��6�6�1��+���۾��پ�d��ٝ�4�>G�G��s>��5>ŭ�=H�><a]�=�X<=�W�=v����	=�I�=.�=���=H��=!	>��>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>s��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��7>!>�R��1�J\�5�a���Y���!?_;���̾��>v�=��޾5Yƾp�3=��6>@f='���\��~�=�o|��?=��n==z�>�D>�4�=�����L�=��J=�I�=��N>�9��d8��,���2=C�=�'d>��%>�*�>ǭ?��0?v�b?�i�>sl��Ѿ`�¾��>f��=Lװ>�a�=}�E>Ӷ�>>�7?��C?��K?ew�>��= �>�$�>�-�M1n����tI�����<�%�?�.�?o �>�h<�C�>u�J=�����B?�]1?�:?�3�>B��{�߿uxQ��n/����=��>Ϙ>�m��[��Ͻ��`>!����=W!�>o��>���>(Y>�P�>
�>�F�>��=���=㨙=�p�C�]+�ezo<dC���p`=�y|�Y�	>�;$>Ø�=�ǀ�/���W�<�ܡ�������=���>6A>{��>��=����>/>������L�pſ=J���*B�3d�6H~��/�7W6�"�B>23X>_����3����?G�Y>�j?>���?\?u?��>!�0�վ�P���Ce�aUS�eƸ=�>=�<��y;�pY`�5�M��|Ҿ�>"~�>㘢>�k>�+�^�>�[�n=���R<5�:�>�p���<�*��|�p���Dԟ��h��=�0D?(���*�=�~?zI?A��?���>�S����ؾ�H0>��� :=��NZp�5x���?Y'?���>"@�2�D������[��*Ҭ> 5�LM�1����*0�-�=:P�����>r
��þ�L�������H����8��>�gV?���?�V����V�@�?!����b����>pw?���>8&%?��>V�w=<�����K�=�NM?��?-��?��j>cy�=C�޽���>��?!6�?�U�?�^x?��]��F�>;�Ӽ<�>�D����	>I�#>���=p>�?ۖ?G�?5���e��Paﾚ]��v>�2X=8�=<��>R�>��u>��=	�:=*cR=�6]>P��>�>�>U2n>�*�>���>������)�%?p�=4��>4?�O�>H%p=]�������9Y�'�J�2��\O������@=��;�Ia=$Y�;-�>��ȿ��?;�r>���H ?���R���U>c
W>�_����>h�Z>�n�>m��>�ĥ>;>ڎ�>�_=>:6Ҿ��>���A ��C���Q�ҴѾQby>Ӑ��N�(��]�E���̕K�F��1�� �i�e���Y=��U�<r�?�-���k�א)�!��.?�r�>3�5?=r���Z��l>��>���>�X��d��'�������A�?���?`?c>��>n�W?:�?Ŷ1��3��rZ�A�u�g)A��e��`�K፿���ؐ
�^)��w�_? �x?�mA?���<8z>���?��%�?Ϗ��+�>�/�d&;��o<=�4�>R1��S�`��Ӿ#�þ�1��9F>܏o?"�?$Y?DV��7���>�2?��2?&�t?�7?[5D?�a;�W'?�>!� ?� ?DY9?��/?V?�VT>��
>���<}��<QH��dZ���o�
ޠ����;��2=�cL=�����P<[GZ=&%�<�r�D�|��(c<b�;�6%<�u=�N�=��$>���>)L`?�?�>�T>y�3?� �O-�8���ړ,?��<i���Њ�e�����C�/>��e?���?��R?��>oU���Y�5�4>�ל>�� >X�`>�Ը>���ڳ)�YL�=	-&>�>���=��V�v���z���R��})�=8�>���>�>������!>Hߟ���m�L@n>��G��	���_�4�G� �1��;m�p��>��L?v(?�ۧ=���(#��f�t�"?~�:?�P?��?S��=̱־��<�#�G�	`��.�>K��<qq����@���68�Qݻ2�t>�s���1f� �x>����v�9g��yi�>���O<><�߾�qx�]?���� }�-�=��>����-��/��}*����8?X=Mѧ�Ɂ��/��O�(>��>�:�>:DͽU�n�]:��޾`����>x�=7y	=:�����%�#��Ǉ>D?ֶ[?	V�?WO��&�w���B��c��׫��X���?t�>3�?�z&>w�=�I��1����f��N����>H�>Mg���J�{ُ�s���AJ&�a��>��?/]>� ?�L?�c?f�]?��*?&�?�>��ܽ�����(&??�?� 7=nB�G�T��%>�x�J�R��>��%?<�Y�Vݓ>ֽ?�?�G?��P?e{?Mr�=���oF����>_�>��W�ǲ����>@9H?�>B�[?�Q�?��%>�2�A闾<���Wq�=��&>�n1?-�?��?�J�>c��>�o.��n4>��>MZ?��r?�Ug??"-��
�>��>��>Hd~>[g�>\��>�0?�KY?v\O?b�=?.1�>O�i<xZ��S���pK��E��vʽ��F=>��=��=�ẽ��<\˼7�=Ա��	��=~��ҷ�Y��=j�=��>,q~>Uy����x>�)о����U8'>|a�<P��%�����^�Oc�<�GX>�9?���>�L�d0T=�X�>w�>#�I_%?v�
?�q?�s��sJ������|�Hn�>�=?Zh9=�a�� ��sfu�*�X���y?7�c?|�b�9p۾��b?#�]?j�=��þs�b�&�龂�O?_�
?��G���>Z�~?��q?���>q�e�9n�K��sDb���j��Ӷ=
t�>�X���d��E�>��7?�H�>�b>g6�=�w۾0�w�Po���?��?z�?m��?y(*>V�n�q2࿢������g`?��>9��,�#?T���>Ӿ�2���r�������΢��	Փ�����*-��<����ݽ␜=L?�cr?��o?�]^?f�zc�iZ�|:|�Q�x��k�OX@�;@��D�Ll�����J �sє���!=����me��>�?W0?Z���\�?w4о���h񶾘��=�R�������/�<����AH>{���к����H�W��l�$?���>���>ۨ4?�c�~F�д����z6��	E= ��rT�>�?�>d���G=���½�]0��E�y[c���>��]?�T!?>�p?��ֽ�PJ��������~/&=�^�����=Ѓ=�ni>�ff� �Ži�:��.A���{�;���u�����=V�E?���=?ɝ>:@�?O��>����ʋ��}��P�4\-����>aG?|�>��>��;=W&�s9�>�Ql?{i�>�x�>Aԍ�)2!�ik{�ӄ˽WF�>���>,��>?Mq>�a*�]s[�����pH��xT8�H�=x�h?����`����>P�Q?:�W:|+<Kw�>�+u��"�9񾙊$�1�>K�?xۭ=��9>�ž��
��z����jZ*?}�?!����B@�ob�>��?	�?���=�IG?��>�K���X>rz?�h?�5?tcc?«�>bi%>6!=a Ľ
��4��=�>P��=��=E�=�?��/������@=�@=y�z[���
�=��=<��=��r=���=�iڿ�rK���Ծ���M���a�	��`���g���_��"��	����A���/u����N�4�Y�p0o����Gt����?:��?7���ʄ��z���_���(��)�>K{�7j���֪��-�sȏ���ٲ��� ��1O�#_i�o6g�M�'?����۽ǿ�����9ܾ  ?�@ ?��y?��_�"���8�Ϯ >-B�<j?��L�뾥�����ο����g�^?0��>d��/��{��>)��>9�X>�Jq>q��q螾fI�<>�?W�-?ϟ�>&�r���ɿp����Ф<���?�@H�A?
�����	�b���>e�?�#v>uM���$�<~��s�>�>�?��?1>�"O�zj<a?�I�=�=#�xŒ�~�=�x=��n<����=>+�>�J�"A�D-�~K8>� �>/+�=�!̽��A�h�&>�@>c��rp��4Մ?){\��f���/��T��U>��T?�*�>t:�=��,?V7H�^}Ͽ	�\��*a?�0�?���?#�(?2ۿ��ؚ>��ܾ��M?]D6?���>�d&��t�Ӆ�=m6�q���z���&V����=_��>a�>Ђ,�ދ���O�J�����=�����̿/F��&���=�O�;�׍���=&,����G/��ͫ���,Ҿ8bX>�Im>���<{�Ӽ�4
�%96>PxI?��d?Q�?�ݣ>�����I��?�jK!�����#�g���j=�U>w��<�!<b��;��"W��0�a���G�� >��F��n���C�+��hRO��UE?x%����쾞�F�ʁ�|]�������˱<��սD���=I�||���v�?��^?�%��Tr��v<�`FǽR��qE|?����+���A�jҎ=M%K�!��<SB�>ʕ�=�]����4��$;�o�5?M ?�����ľ����}����<A�?S�8?���>y��>�"?ĶW��_��
�=[xA>8.�>�3?�/�>U�q������?W�A?C��_5���>2x��XB@�>k>�헽�UW�32e>%]A�g�@��=X�=ࠋ�9~R?�T�>s���0#��~���L�<�pN>�P?�k�>�>��X?��P?�L��c����N��l���2w>�k?��_?w�>�t׽-��H|���7?/�S?�5�>���3�N�%��O���(%?r�?1�.?���=i#�3�����/?��v?�r^�[s�����l�V��<�>�[�>���>��9��l�>T�>?�
#�wG��Ϻ���Y4�Þ?��@���?��;<�����=o;?X\�>M�O��>ƾ�y��1���&�q=="�>q���wev�����Q,�:�8?ߠ�?͔�>9���ש���=='��W�?:�?,�پ�k��B��Qg�(9��9
����k<g�\�$�û���c\,�LѾc!�Ø�1Y�x/�>Z�@�VC�l��>��~����_���Z2^�����ga��X?��o>f�0��(¾]�j�ON`�?F���M��9��$��>��$>�����fo��d/���<���>�d����>�l�����"���;��>#C�>�Δ>3`-�.������?�k���ο"8�������lU?1_�?�Lu?�	?��<��N�����p�=�vK?O�x?Z?A3�`��F���F�j?P����jV�|=2��lN��?>��)?l_�>�|���>��?>~]�>�C >�$��ſ�i��𾟧�?F��?FMݾ��>g�?�7-?Q��%��������%��{!��H?q�X>�竾�d��/����!t?��:?^d�����\�_?&�a�L�p���-�s�ƽ�ۡ>��0��e\�?N��	���Xe����@y����?K^�?g�?е�� #�i6%?�>b����8ǾV�<���>�(�>�)N>�H_���u>����:�i	>���?�~�?Mj?���������U>�}?($�>�?��=`�>��=B谾��+�`#>3*�=��>�
�?F�M?�S�>�N�=*9��/�eRF��AR�b�{�C���>i�a?~L?'Mb>�9��b=2��!�d[ͽ*d1�Q �:L@���,�5g߽w55>U�=>y>��D��Ӿw�?�d��ؿmb����'��4?��>�?���jt��L��A_?���>�$�B.��c��������?�B�?l�?w�׾�̼�)>��>3�>.�Խ�՟�T�����7>��B?R�B8����o�	��>���?�@F̮?xi�$	?��"N��m\~�3���7����=��7?.#�N{>B��>4K�=�ev�;�����s�p��>�B�?�{�?4��>�l?�~o�V�B���1=�P�>��k?u?�l���+�B>��?������iG�Lf?��
@jt@l�^?���!׿�	p��U�׵>�`>��h>�н��<���E����x�q�,���
>[�5>�f>��w>�o>vU7>����*�iá�����3�+��|��H�uF��s�(��6�#�O�v뾉_�,Q��<F�x��������仾�m-���=0�U?sR?=p?� ?)Yx���>�����r=��#����=7/�>�d2?��L?+�*?x��=�����d�%\���7��CŇ��{�>�nI>�x�>�K�>��>I�9Q�I>8I?> y�>�� >P'=<^��wM=��N>�G�>���>�u�>��>2��>�6���s��d����3�x�0�x��?��D�\V{�o����GC���F����\CD?0�˻���dҿڮ���?]f��,�����<[t�>�^?�1?%Ͽ=��!=���=��:�B~\��ž��N>W^8�5�Ӿ� �� ��=��^?�j>�L|>��4�t'7�vN������_g>�H9?���n�C���t�T�G���ھTcA>���>Lԃ��A �$K����/h�\�o=G�8?�,?�
��j���
s�ܝ�2�X>��]>��<��=��C>mhS��ŽksK��/<=R{�=�h>�?o�
>�<�>���S\a���>b6>��>'l?�9o?�1>��L>���z辂��>��?o3	?|��>����s�=�T�>�O�=�S�� �v��H���O��7t�=*�O���I���;�P>[�=*>���=4R=<B)��c���~?���(䈿��e���lD?T+?S �=��F<��"�D ���H��F�?r�@m�?��	�ޢV�@�?�@�?��N��=}�>	׫>�ξ�L��?��Ž3Ǣ�Ȕ	�/)#�iS�?��?��/�Yʋ�9l�~6>�^%?��ӾGl�>\���)������tu�<�&= �>�/H?zb��O^N���>�ad
?`f?�򾼌��F�ȿ��u�kR�>&��?h�?��m��U���n@�e`�>N{�?��Y?o�g>�ܾ�Y��Ό>kVA?�aR?7��>&���Q&���?�޶?Ҭ�?kI>ь�?��s?�l�>[x��W/��3������`o=�B\;uc�>nQ>5����eF�Aؓ��g��f�j������a>T�$=�>q9�v4���D�=F���+I����f�/��>M*q>"�I>�W�>�� ?�e�>h��>�P=�g������'����K?�Ï?u���m�8��<���=r*e�K�?�d4?�<����Ͼwi�>Jj\?��?�[?#Ǔ>��X�������<�.K>p��>���>R1��WfI>܂Ծ�?����>N�>����-1۾����q���>W!?��>2��=d� ?�A#?�j>�ٰ>~�E�������D�y�>���>�N?�\~?��?߂��!W2�+(��������Y�=�S>�y?�?H��>�9��᜿�V�MrN��1����?�e?�1۽ƥ?�Z�?��??i�A?=^e>�3�@,Ծ�H��}->q�!?G��?A�%*��P����?RT?Y�>�
��E�ý���A��E�s�?��X?�(?���I[��H��Z�<�ӏ�:����<�`?��>��>��;	�=P�>�,�=H2i�Q���_�<l��=��>R��=�8�F���%=,?��G�eۃ�m�=z�r�:xD���>�IL>
����^?m=��{�����x�� 
U�� �?��?1k�?4��;�h��$=?+�?,	?�"�>rJ���}޾a��.Qw��}x��w�	�>l��>��l���0���ə���F��_�Ž�ǽ��?�?(x&?�� ?f�:>'u�> L}�hs�A����.���y��7d��T2�Ôh�����m�a­���p�Uޤ�5dM���>�Xt���>\-?}UE>W&�>��>��=eֺ>+��>�`1>\��>"Ό>���w>(�>o�#��&R?p����'��&�����=B?/�d?A
�>ɉ���؄����5� ?��?{q�?��u>�4g�hF*�BD?Xl�>[�~�B
?1+7=!$&���<;r��l����������>�kֽ�9�S\J�ۧc�p�	?�C?�਼��;8kӽ�ɗ��B>=5ڄ?��4?*%D�Rk\�?Zl��nG���T�%7:�۩���X���\��{��i���� ��.6(���ӽ, 6?"��?�:���׾�c������0�J\�>��>��t>`��>�w�=r��&2�&2R�����n�Er�>��F??�>�<U?_BS?S+?�h?��>���>�!�ϐ�=�f�=Pϟ>?�)>? vF?7iK?� Y?!O?ڟ�>�� �iT뾱K���!?�2P?���>�V�>�f�>���'�=���/=>)���/U�Gv�d>���:�%4�;wᆽ(E>��?/4����/��?��>-�/?b�>ש�>����qa"�CVB=�??�+�>Cf�)�9�������>rf�?¼�3u=&>���=P���-���<�y��Y�
> =�:�ԕ���<�7>+m�=]�v���=�ة��O�5����:�>��?TÊ>�.�>'M��`������(��=H�W>}-S>��>�;پ��䗿]h�:u>q�?kG�?��h=U��=�!�=
������$��F���� =�1?s0"?AT?�~�?X�>?�#?Vx>���꒿�Ʉ�����?z,?�ȓ>͠�����6����9�Da
?su?hqX�_��Ԍ+��1Ѿ8��ms>�+��'������ƻD�K4����;g�����?�?��|��*�����n���|���@?қ�> ��>D�>�N*��}l�;|�X�U>��>M�R?�a�>#�O?{?At[?�S>��8�C��򹙿ԉ$��#>�P@?崁?��?K�x?ۗ�>��>^d(�% ߾r����n�6u�,�����W=�(Z>g_�>�)�>� �>î�=�,Ƚ,���?�9s�=P�b><7�>å>`H�>��v>�Ũ<�I?�7�>鍺�Z.��䵾Fㇾ�I�0�n?��?�5?mc�=���2;�0��K��>|��?�?�?��0?#�1�'��=��켝u��!�f��[�>�|�>0U�>���=���<M>7��>�e�>j���� 5�0��X?uA?��=�]ɿ�政��9��ԓ�H�삗��ܬ�����������������9���B��Q�Y���,����G�����I(��F��>F����;>���=��-�)�=���$dp=���=��>IQ�Tlڽ"�H�]Ve������A�Xh�=���=X��>�ʾ1:}?I?�+?V�C?�4z>p�>*3���>*I���V?��U>��K��@���;��L����ؾ��־<�c�䎟�=<>�L�8�>�;3>{�=SX�<���=��t=6q�=�m��{=���=a��=�z�=J!�=�>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�}8>�B>1�R���1��o\�5)b�W�Y�xY!?� ;�,�˾��>H�=��ݾ�kž�,=�V7>��f=���ֽ[�T��=�_x���;=r1i=��>�rC>	�=����i�=čI=��=�qP>�\Z���8��(���8=^��=�)b>~�%>���>j?�k1?��c?�Һ>�se�J�˾
Iľ	��>�`�=8�>k#�=JG>�I�>��7?U	E?�J?�t�>�:�=Lz�>4o�>lu-�D�m��徂)��}7�<�s�?���?���>$�]<�UE��N��:?����?`0?D�?tš>ga����/'�~e/��_��{qU:��%=�3q�o�X����IA�=򽜬�=�#�>l��>�۞>*u>A7>�oM>�L�>ng	>��<x��=:1F�G��<������=e�d�.T�<�aмaX��G��.,�����%W; ��9`�g<%$<%��=�g�>Դ$>-��>�6H=Pc��jyZ>g��V�C�r��=��վU�K�4wt����{�F�7���N@>�t�=]��֎����>��>�]>=F�?���?s�'>��I��P�wpg��(j�@=�Ì�=�2m���-��W�O�G�U�����>��>�Λ>�<�>~�,��@���=�^ܾ�_2��!�>������M�gw�i�n�VƤ��͞�_|f��m`���@?lɇ�r��=dn�?�]G?�"�?`�>�A���޾�x!>b|��8�<��SY��`���?��*?ݚ�>��,>�j�ƾΌ����>�=��I��ő��m*��~�;{?���>m�����Ӿ_�8��2��2z����E���Z���>L?��?�h�������Q�э���T��4?�md?+��>��?��?2��#K���r��=��i?u�?��?	�>��>��;SJ�>�E�>��?���?�+f?Z�H�`��>�vw=}�>s���G�=
�W=��$9=)�=D?y�?��?͟<���"��ɺ��W�o�=��>�w�>}�2>��B>�r>���=�v	>׷;>�2x>W�>�m�>B��>+��>�����)?��=h�s>�Q0?FYM>���<Q5�W��<�*̼��L�DI5�;����)��i���	�<��=��x��6�>����6�?.�N>?���?�������.Z`>�S>n*�<
�>�=>?�\>3ԭ>��>��=}M�>C�
>DӾ��>���:L!� C�,�R�Ҿ {>�]��ol&����O:��E5I�̏��@�Qj��-��X=�;��<t9�?PX���k���)�������?\��>��5?+Ì�������>�{�>t��> ��Ї��ȍ�f#��
�?=��?V;c>��>�W?#�?@�1�e3�!pZ�u�u�6&A�1e�ʼ`�N፿ �����
�14��I�_?��x??vA?�e�<S=z>a��?;�%�ۏ�4&�>�/��;��n<=�%�>:%��C�`���Ӿ �þ;/��ZF>�o?�%�?�b?�LV��=�{~>`�F?O�+?�rb?��?/
"?ce3�&)3?6c>�? �>�97?��?,��>�?>k��=n;��=��̼�3y�@mA���� ,�� j=�xV�$-�=!�_>�}�=��̽�����m��	p��>�=�W�=�B)�)�=���={G�>��[?�#�>���>��6?p_���2��	����,?s*\=Fby������ٙ����L[�=Pj?H��?��Z?��m>��A��.G�C�>�3�>��$>(&X>.h�>*ٽ`�M���x=Z�>��>��=��o������3m��B��<�>��>>��h��>F����0��2|>M~�����#�i�z�X���;��X��+�>�O?�E?�ҭ=;��@Z۽Gc��J$?H&`?�4?�}?�[�>5�=�ŷM�o|U����~.>=��(�;G���r������.]�=�Q�=\����S��J�\>Z
���߾�Ek��J��뾖#r=�>�|e/=���׾υ�y��=<�>�Ŀ�"�"�疿�֪�p?H?��=�`���?Y��G����>�>�*�>�4�h��d�>� a���=C{�>[@>�����3�0�E����px�>(3D?��a?��?PW��ܰq��2<�����\���X����5?^��>A�?�D>!u�=T�������b�p-F�ɇ�>���>y{���L�4���	_�R��1J�>�R?JC9>b�?��U?`/?��Z? �-?�
?f��>7�=�������$?+U�?�w=Π�n�S��o;�� G����>�M(?��M�s�>��?6?�#?��O?<?gI�=n�e�@�L��>�ȋ>��W�-����a>��J? �>��V?=��?�=>�i5��C���'�=�>61?�
"?��?��>4��>�j���w>���>_�d?�.�?�Kw?��=a��>��H>��>8�>ѩ>$x�>���>gZ?�d?O�9?qn�>�j>�n����	��ԧ<<%l���;�F��;�<>t,T=C���O�<L�=/�G=_�սA=��0�������畼^r<K��>Ƚq>������5>!X��{��N�F>�3�����NF��=k!����==Rx>�n�>���>0i)�B�=��>t�>��4�"?�I?��?	"+�zV[���Ͼ�8Y�j��>FJB?�o�=�l����Fr�C�,=Ҳj?�7[?;i����\�b?��]?�l�x=�0�þ0�b�"��	�O?�
?��G�i�>Z�~?�q?o��>j�e�}7n����D(b���j�ן�=�^�>�R���d��N�>}�7?R�>�b>?1�=Uc۾q�w������?5�?��?1��?�*>A�n�N*�l~���T��'�b?���>����� ?��L�ھ�ꎾߌ����⾒���ھ��O��u��4�"� 熾��텋=�W?�6w?k3i?��Y?���xk�w�^�(�t�n�T�����	��E��=B��B�Rr�?�]���8����<מ̾ss����?�UN?�㥾��?=��^�������>]L���1�6�w�<�/�>a��L�R�7���ݾ��4?���>�o>,�G??怿?�]�C�'��;(�pվP>>��7>��J>�B�>������A����������G�q>7�d?C/L?��m?���a�2���}���#�~��퉢��y:>+��=`��>��D��m0� ���:��[v�������s4��ƫ=�:4?�ޅ>�͢>�[�?�?\������-kx�L*���];-�>��f?��>e�>o宽������>p�k?R��>
6�>񑌾�� ��z�g�ѽb��>\>�>/k ?��r>��+���[����~��'8���=�mh?B�����_�p"�>:FP?���:�f\<�>�Ln��� ����k'���>|�?ר�=R�;>�ľl��{�8r��0)?	?� ���.���~>"$?�P�>O��>�W~?�ؓ>,|ľ=C8<!j?�b^?�p??��=?Z��>7t=�R����ؽv�"� �]=�\�>�c>x�T=��=��)��R�m�'��]S=��=��@��1���j;T8���d�<�#=� =>տ�
P�ǧ�����J���a��\���[�;<���s۽Noξ�+���hx�j��V���;�+	��N��YW���W�?+��?�-���9�����Ԋ������>.��"S0����-������^�վ]˾�C��W�D|�`Th�O�'?�����ǿ򰡿�:ܾ0! ?�A ?;�y?��*�"���8�>� >E�<0+����뾢�����ο0�����^?���>���/��S��>���>K�X>�Hq>����螾�.�<��?1�-?
��>��r�*�ɿa���FĤ<���?,�@�FC?���F����)�<H+�>�?�<>�fN����>�ƾ���>�W�?=�?� %�f�[���-wo?���=!�u���f=�B�<�U=$}H��e>��@>�{㽡�꽤�����=� �>w�9=j��W��@&=|�X>s�M��9�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=]x���տ�+;���%��e�=�-
�56z�����'>�̵>�7�O�k��N삾���>�ѳ>���=ɞQ>
N@>�{R? À?�?(�T>�{<��½�x��:�M�v�"z���2ӾЉ�W>������~��y3Z�'��wC&�a���$��=���Ҋx���U�ր�d�S�`�T?D�����6�q�ѕ���޾���jx
=����a���`������/�?/�y?�Ώ�؝g�4�A�v�,�z�<�y?��"� GD�;����rA>-���b[=I�f>�.Ĺ���������R��6?� ?Q�£/���>���h]���Y?�y?�a�����>Z�G?ON���)'�> 	=R�.>�a?�F�>}D��l�?�2?�zD?ü�Sl�Ee�>,6�PR{��]$>v�z=h轾�݊���>�>�Ĉ��"�2p�*\!<ҕU?H3�>�7�T)��O��y�E;� :�[?H��>J>�iW?��^?L�I>��پC���˻:>�g?��l?���=�8��j� ���~��W?�25?�����&<�XA�(�-�)/����>�f?ɳ
?�r>;$g�"`�8e��x�?��v?��[��������Z\�v��>A|�>,9�>�>9��>�>c�=?_�#������r5�I��?K@��?6N�<������=�	?��>�E��{žbԽ\W��!�=7��>�	��h�u����ҽ)�!�8?�>�?��?�@��t����=�1���?�Y�?�^¾���;����k����6|=)��=�PQ�3\7�K쾿1�O_¾S6�LQ�� FU��Β>j�@�Q��\�>��F��g��Ϳhz���о>n���4?���>�нП���,n���n�\�J��_P���� ��>��I>��9����T���4�ȱ�=���>:N"�k]�>��ý�D��٠`��<�=;K�>#?7)�>�ᑽ�s����?
C��QӿL������?Ea?�*�?���?��>ys���U������}	>QbN?�ar? �<?��?=�Bq���">\Yh?������\��:8�PN���>$B?;$�>P�(��% <h�@>
��>�O*=�^A���¿v���=�����?���?tuپ/��>��?>�?�a�΋�8F�(���|=2%?����߾�F��f',�m`���?�NK?��j�ڮ��_?<�a��p�n�-���ƽ9ۡ>�0�a\�ov��G���We�\���<y����?�]�?q�?��L #�B6%?+�>[����:Ǿ���<ف�>�*�>�+N>�<_���u>]	�^�:��i	>r��?A~�?�i?4���B����W>��}?�A�>�4�?�Y�=���>��=�V���`�%�>���=��?� �?RM?�i�>\D�=�.-�+0/���F�0,N�R��a�B���>�a?DCI?g�Y>A­�7��H!�r�׽��(����BFH��C5��/转q->JG@>�>��N�L�־9!?���ӿ ;���vV��H5?�~�>��>-5����2=K�Z?��^>mC�w���=H������UA�?���?� ?��¾���x=��>W�>w���,�3�'∾�}>��*?��H�������l�~�u>P�?a�@��?HLZ��+	?E��iD��J~������5���=�7?i9��y>���>��=�kv�忪��s�웵>T8�?Cj�?�6�>]l?;o�M�B��[,=�[�>�gk?:�
?�Na�X���A>!�?*������L5�Q�e?�
@�o@�^?nƢ���ٿ䇣�~(�N�ݾ	S>��> p>�&���>~>�%�=O�.�5m=�>���>e��>�G>�7>�J,>A9����%�8���q���y�1�����n�6��+���t2����þ*b߾�*�y
��顼m��7.2�`��O��=��_?��a?$}?�n�>V3U���)>~���w���Ͻ��z���=P??[|L?N��>�A>�f�����n�t����TxҾ�H�>���>���>C��>h��>��=OZp>�|�>�R>_�o>�ӽ�_����O>�A�>As�>�� ?W�>? >^p�>�*��ƌ����?��y����jݡ?<Ҿ<��r�C<��[���&�M�!(7>j�?�&=�ޝ�*�ƿ6����b?'.e���J	��z�<�?�'_?
��=񣏾�y=���>�T��Av��}�?�_ս��Ǿ�Y��ү�>ߢ�>S�@>�&�>�E0�~�3��&=��^5��(����l?Gl��6	��҂�"�D���þ�r>���>_t=���M�m������"bd� �@>	��>+��>G�=E&��UAW�������>��R>D݄=v�@=���>��L��?��W�:���=	MX<'��>?'�>�ņ=��?ό��^����>�8D���;>��A?��@?�O_=��IJ��_�x�S�<s�>�Vv>��#>Q�ν���=2)�>���=�X&�����#s���P�L�j>�%�=.�Խ�8�����=ս�EP<*.�=�)�T�����=�~?���(䈿��#e���lD?h+?s�=ՔF<��"�: ��gH��D�?n�@m�?�	���V�>�?�@�?��E��=�|�>�֫>~ξ��L�ڱ?��Ž"Ǣ�ٔ	��)#�^S�?��?��/�Xʋ�Al��6>�^%?ѰӾ���>�.�P���B�}���t���N=���>�:?��ﾈ�_�`�&�?�1�> ������;�ʿ�fh����>g�?�|�?'�a��P���5J�4��>���?��`?�>�������f>Ny5?DIA?R��>����%�c�?��??��?��I>�\�?�s?�9�>��|��}/��곿����!N�=#Ǟ;u�>D�>����ZRF�}ē��d��0ij�'���a>\U&=O�>��䯼����=����][����g�S�>PAp>wgI>��>X� ?0�>�D�>�=*<���V���)���K?���?S�K3n�.��<�ݕ=��_��?/>4?՘���(о���>E\?�!�? �Z?H�>Y��\$������)�����<�J>�h�>,�>=����aN>��Ծ�GF�ؚ�>�Ҙ>�K���پA|��ԡ޻k�>"�!?��>���=�v%?7�?�r�=�q�>�pA�H⃿�9&���D>6W�>��?���?sr$?M����*����"���$7��%6>X�l?s?<��>����D ����T�aUh<yJ���d{?�&F?�ك�'��>WJ{?�?9?:�L>mS��Ӿ.��9���>�J#?����X6�zQ�VjŽҟ?�?d��>��� ����d�;��v������>��\?��?uA�F�Y���沌<��	�]@
��O<x.��@XD>��O>$g����=b/.>��9=ǋ��=8�|r<�e$=8�>��=�[e��v���=,?�6G�H߃��ǘ=D�r��rD���>9BL>-���?�^?�p=���{�����x���U���?Q��?�k�?����h�[=?�?	?	0�>�G����޾'���2w�7�x�d���>���>Sl�W�9���ܔ���E��1ƽ�o�7f�>�U�>a'
?�[?��b>�T�>�!��)#�R�侣���^\\�@����8�6!'�*������W�$����
@��פּ�(�>��c�	��>��?0y>�7}>ܙ�>Y��;L{>��E>��r>���>� 6>BKF>C�>E����ܽKGR?�a���<(��k�Mǭ���A?��b?q��>��Z�
J���}�ZK ?mC�?�ƛ?��v>�g��H*��?2��>.^���d	?�:@=#[��-�<���v��J�������>xmڽ�?:�1M��-d�o�?i�?���m̾5�ӽA���LU=���?�3,?�+�_oP�2�k�s�V�xCR�a��P]a�矾��#���n�Q���9�������'��7�<�t+?�ʉ?j����H`���Kn�	{?�.al>F �>�,�>��>n�F>6
���0���]�˦%��|��]�>xw?JA�>291?:%;?&w'?1A_?ޝ�>>�?5p���>��;��f>2�?XI1?AaC?��>�UH?��G?sD�>E��!�pն��;)?��?KL
?�l�>ⴤ>f꒾��>�Ѱ=��=�s��z��l߽6^s=w�����h��}�<�=t=�9"?5푽��?�p�ġ>��=?M�>��>��1�c���{��-��>��&?u]h>,���rT�X�g��o?�Xk?݋��H�p<//9>	S�=ue=���=�2r<�˽D�4>s�.�3��'��	!=Y��=���>ͤ=�|�=��;�D�<�D?��?�i>�҅>mny�P��4���ñ;�i>� )>M>v?���ot�������h��K>6�?�ݯ?V��=���=���=�谾�q���}�V��,�<j�?��?��G?�=�?3�Y?z�?6�u=z}������>���z���$?c�?5�>]���ൾ�ҟ�egR����>���>C�_��"I��� ��!��eT=�>>��P����
l�WF׽w���)���?�I�?�8�=��Ŀ���������lX?} �>o��>M�)?x�<��񃿉R��jC�>p5u>{�[?>��>jO?�z?�m[?բU>��7����]����P6�EO">�@?vA�? N�?��w?���>' >"p+���޾����"�Ѷ�����Y�N=�`X>`Г>�>9u�>ߒ�=!s�������'B�io�=��_>7l�>���>8L�> |r>C�<	�G?���>К�����e���W��!6�}�u?�/�?�x+?�=|�OFE��#��� �>^�?�߫? *?k�R����=B%ؼ�Y��Zr����>�K�>G9�>�ɔ=�tD=��>m�>��>����Q8�ŚR��?FF?�q�=��Ϳ����>����x��҃�=nL���C�����Ը����M>橉������
��ʑ��(�CC|��\���G������L��>�л+�\>Ȟ�=5R����0=�)�=��Z=L��)=������<�/�<v>�=y �=���=��=���<�*˾�c}?�;I?��+?�C?�(z>��>O�4����>؁�;:?�&V>(TR�7���h;�v���q1���ؾ�׾��c��՟��y>�{H��:>�3>��=���<i:�=�r=�2�=�,�Lu=�%�=}�=�l�=��=��>,c>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>?9>��
>T�R�1>3��+Y�xh�{�Y�5�$?��:�d�Ͼ�|>�D�=R�׾þ��*=�g9>�K=
����Z� �=j���!=ˊ]=�G�>��I>���=3����=(3=C��=��N>9��9[�;�R�:�e{(=���=�0b>4..>:B�>�i?�<?�dl?��>�?���ڲ��4���
G> !>�8�>��=��@>�l�>A"?2L?@�@?�Ö>�g�<���>
m�>~=3� '~����#J�����=a$�?Pl�?�>%�>�����70�?Ƹ;��!?�|4?��?��>���ݿGb���0��0����=
�=�|�v�����<=����1����M��>g��>���>��c>�>��+>��>�<�=��=���=/#�7�=�=�,{==����$4=���}�,�(B"<�T�;���;��J=��M=�$a=�7=.��=y��>�>���>�)�=�U���/>�Ŗ�DkL��|�=�o����A��c�/^~�@/�W�7�d�D>��Y>�N��y�� l?��X>��?>b��?��t?�>,q�3kԾI3����g�o(S�M��=�>	>Ed<�;��_��M�rlӾ�	�>ڏ>�J�>|�f>V�+�@S=��z=���(^4����>l����M#��f�gq����bԟ��|e�c�;��D?����, �=$S|?TAI?�v�?к�>���F�ؾT6>�ۂ��s�<�%��xa��;���~?̅&?<c�>O��E��bžqn���g�>�XC��1P��t��w�+�Vb�������>�T���qɾ��2��y��>+��W�E�-j����>igP?��?��\��C��K�Q�Qm�#�E�_?c�g?t��>�� ?�?�묽�8ﾛ���կ=�l?���?q��?	6>�(/>8�����>�? ��?��?H@[?fO�o;�>~�<|�P>[�[�2>Ļ�<��=qm7=��>ݜ�>s�?�7�{�	�ڗо�n��r���%�<L�==v?>��,>N�q>d,�=��=��}y>�)�=�T�=��j>-_d>p�>gm����Y�-?�Z�=�l�>|�7?�S�>(6`<@�����=�/~� �Y���m�Y�w����d�<��r��%=nJѼ�.�>�ÿ&;�?���>Ez�}G?o�޾\��D�<>V>@\#����>�ml>Bl_>:�>)6�>���=�"�>ݳ�=^HѾ��>'���) �<2C��R�1Lо06w>�ٛ���$���γｄ�I�N������e�j�
�����<� �<�ԏ?9���Uk�7�*�����	?k�>�T6?����l��~>Ȇ�>߆�>����%��.���a)߾{b�?��?�Fc>'�>(�W?��?Q�1��	3�jmZ���u��$A�|e�w�`��ލ�ҙ��~�
�_:��+�_?��x?�yA?�˒<�5z>4��?`�%��Џ�56�>�/�0;��3<=�9�>�'��a�&�Ӿs�þ�+��XF>ǔo?�%�?�V?SmV�=�U�� 1>�C?Zy-?v?|7?��B?x���� ?]�>>;U?��
?$n3?��?*:?��q>L>�Q<!É=�½��a��������g�I=���=�!D=���<ۀ�<�_=�(���;D�2�U-���<ʅ<.Ί=�9�=�_�>�WJ?p�>t�A>aQ,?��F��D��ݾ_�H?�,���Ȋ�Y8~�lE9��Zؾ|<�J�K?H�?�]?���>~+F���9���$>X�_>o"�=k�=!��>�S۽/����_E=��>B�>z�S<AV�΀4�-�žYp޾�=Z#�>aT�>�T>�p��o�'>姣�x�|��d>��R������S�ϏG�b2���r��'�>,�J?�?�r�=�뾩	��_f��(?/�<?�M?z�?~��=�ھ]:�~IK��C���>?U�<�,�D��������9��WZ;�r>�q��Ƞ��ub>���L޾�n��J����vM=����pU=���վ~N��V�=h�	>����� �	��ت��$J?��j=nv��w}U��;���>V��>��>��:�Yw�w@������=g��>	�:>�Κ����`nG�$.�߂�>0C?�VF?��? /о�~��B�X�t׾o�ľS��^V?j�>i[�>5z
>�n��}��5�Wj�.j�.��>W�>��&���P�se�����4�>�>y��>sI���'?_?��>a�T?ܕ?vl�>��w>_��:��ϾOl&?3M�?9n=�w��\R��8��C�Ñ�>��&?�y?���>a?�??&'?<�Q?^�?m�>� ���?���>��>�iX�����<d>/�J?fǳ>5=W?q��?�<>ݍ4��s��������=�%>q3?�#?�? �>�
?�������!雽�N?<6�?�X?�>*��>G�>�>?�4���=o?�Mi?G]G?��K?�O?,JS?s���f��NЄ�����\靼��;�͂���+<M�ۼ�ڽ�MY��B�=B.�}
n����s⓽������:h1 =��>�}u>>S��1>���������D>�f��枾L3���8��7�=�>3�?�Ԗ>[�j��=�>ނ�>���Ʀ'?�>?�?N�;;��a��|۾ÁM��]�>��@?�}�=��k�����v�Ewd=��m?�^?-8U�͉��U�b?��]?�j�p=��þJ�b�)��5�O?��
?��G���>��~?l�q?���>�e��7n�Z�� Cb���j�3϶=�p�>1Z�.�d�FD�>˜7?rN�>��b>!�=�p۾��w�Kc��T?��?��?���?':*>��n�f.࿏�������+h?ë�>�仾�)&?�	P���þ��l��f��߾!楾Jf��@����������z��D�?/�=�?�(z?v]n?�H^? ��)rk���Z�:��^�]��3��	��#�F��X:��-C�ĭl���j]����[V=:n���<e���?o_3?N��1�?�򖾖���$�4����>�Z�������	>�(��⑽��>�U� \u=���I$?e�>)��>#�=?Ge��8��(�:E3�
!�K�> ��>RiS>���>�3߽��D�z�+�4���Dc������V�>~�a?�?a?���m�E�ΧZ�]�A�����ۿ�ye>r,8>��罩F���	W��T���7�1��������� �
�z�;=��8?�b�>Hݼ>��?�S?H,۾��$��m羫�a�+[���>�wZ?�\�>�a�> �=X���>��n?�'�>�ψ>Cd���K)��9��!��e��>��> t?.��>f�I��fb������m��Q<�b�=gU?�Ԃ�g�Lt>��S?��(�# �<8G�>�?�����+H�n�#��B�=��>�V|=T^E>C!Ǿ;���w�k�s����-?�?M��k�3�NN�>�?aY?j�>��0?���>�F��&�:=�?�L|?�P?�2@?pV�>!��;r*�;j�*��hMm=CA�>C"�>�G�=�An=�C��y6h�:&���B={!�=�=��.���W��A�=34�<i}=�EH>?mۿCK�p�پ�
�E��>
��爾ᥲ�pc��E��va������Ux����'�V��6c�2���J�l����?�=�?p���^0��.����������߶�>ߑq����}�=���*��t��b���Od!��O�&i���e�P�'?�����ǿ򰡿�:ܾ4! ?�A ?8�y?��7�"���8�� >XC�<-����뾭����οA�����^?���>��/��o��>ߥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���}¤<���?0�@��A?�&���X=��>�	?.F>�(5��_�RI����>��?ě�?M�l=Z�T�$�׼se?M��;�E�������=v��=J!=#����I>�H�>Ѡ!�=����(23>�L�>�H�V���K^�.g�<1a>z�ͽ��(Մ?�z\�]f���/��T���V>��T?+�>�9�=��,?�6H� }Ͽ�\��*a?�0�?Ħ�?�(?kڿ� ښ>p�ܾl�M?�C6?n��>cd&���t�(��=<�끤�����&V�Y��=6��>��>�,�0����O��L�����=i�����#�����O>e��=5�۽g�s� �X>�਽�F?�_=��W��>"g8�Iݽ/ѡ>x��>i��>�=��I?
K(?,��>��7>ֈ:������8�E >:Վ�w��.C�q�����K�|�܂ �fp¾I���ؾ�N��=��*�=*,R�G���N� �V�b���F�-�.?�G$>W�ʾǿM��c,<]ʾ2����ц��X���F̾�1�@0n�?ş?>�A?������V��������o�W?'j����滬���=�w���>=E�>��=\�⾜3���S�
�0?^�?�bʾsҒ��D>rR���=H�%?���>��:��>�/%?+��ϧ����k>S�D>�f�>�;�>�	>���[ٽ�?�)U?�|�����'�>Z�ž�2t�#&=fA>��%�o���F>�a;<LU��3�ǻ��{��ź<D&W?A�>��*�l��<���5���O=� y?�?'Y�>��j?�B?�s�<B��j�Q�p[
����=E�V?�th?�>5����$Ѿ���D6?��e?[�N>	�j���龆�.��P��S?�+p?��?6���|�{��g��UB�2�6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������-�=����rݵ?P��?��+��>�����Ļh�̾��>ކ<��E1��=J<�,`I�;���͊.����Ľ��Ga�>�-@�׷��e�>p U�`	�X"Ϳ�s�h^�d�վ�$�>��O>�ҽg۽j}B��i���6���֏����$a�>��c>٢�iA|��TL���0�	�>=�?
j��u�>@�(�A�Ҿ���Y><D�>�R�>$��>?=4�mV��R�?�����տ!�:�;\bS?s�?v�?<��>r�1=O����$�<kfw>��G?���?Wx?iwA>�PU�畠�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�h�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�VҒ�¼
?V~0?{�f.��_?Ta��&q��&.��dŽ�>�t.�0%Z�� �~����d�$����y���?�M�?��?}X�k�"���$?^��>7f��]�Ǿ*z�<`�>p��>�'N>xDd���t>���W�:��Y
>���?]N�?d?5��ק���s>�}?m�>4��?�	�=l:�>���=uʳ�FA����>�%�=.TQ��5?�cN?:�>MN�=�;��'0�F�F��FR�Ь���B�b�>s�`?�dK?�c>ը��*;&�\� �ʽ��0�Z(�}9=�t,��潐�2>�=>��>�WE���ξ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?oQo���i�B>��?"������L��f?�
@u@a�^?*u�п块������8;�ڰ=�>�=s:>�f7���=��;/��S#���>��k>��/>*l>�Uk>�3>)	#>����+�$����h��a�9����0�f�b�9��)l`�K��e�� ������Z"�a�	��`,�m��G+��6��=V�U?A�Q?�o?Թ ?g"x�Z >���`Q�<�7$�"�=�t�>�W2?��L?J�*?��=tE���d��?��iI��b���߹�>��I>�n�>j*�>�ԭ>	�����I>��>>U\�>Y>(=F|?���
=�+O>�i�>m��>Ra�>DF<>��>9ϴ��1��7�h�uw�{̽C�?����J�
1��
8��ۦ���p�=c.?&|>���s>п�����1H?����/*�־+���>��0?cW?�>����T��8>
��A�j��b>(' �>zl�6�)�3&Q>�l?��f>>u>ԛ3�LY8��P������+|>O26?����m9�êu�ϜH��`ݾ�MM>x��>w�G�qr��������si�w�{=�f:?�r?#��а���u�|<���\R>�\>��=+�=qZM>qJc��ƽ��G�O�.=��=f�^>�l?<�,>6�=�f�>�Ә��N��>�>�M@>��)>�??��$?K|�3���������+��2w>L�>9�>ъ>
�J�u{�=	��>vb>9��0��(E�[@��3X>ە{�p_�>u��z=�U�����=&D�=�	 ��<���&=�~?���)䈿���d���lD?U+?] �=/�F<��"�C ���H��E�?r�@m�?��	�ݢV�>�?�@�?��H��=}�>׫>�ξ�L��?��Ž7Ǣ�ʔ	�,)#�iS�?��?��/�Yʋ�9l�6>�^%?��ӾPh�>zx��Z�������u�t�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9�~�'���?�޶?֯�?y�>�P�?�� ?�Gl>R���Y h�}��Y�W���:�8��b�>���>���@��:��<ԏ�������5�Zh��f嘼V�>p������Sd>��=D���<�/]�>���> X>!E�>2�>��y>"�;>��j>k5>+���s>��K?0��?�F��n�_?�<�=�>\���?8I3?[>h��EϾ)
�>l�\?r�?d[?t�>R�F��Ƅ���o���#�<ML>���>���>ٞ���ZJ>ӏվ�ID��v�>�>+ޛ�xپ�u��f����>J!?Џ�>��=�� ?)�#?Bj>�>�AE�I���$F�J��>�/�>\�?�~?��?L ���:3����䡿��[�{�L>�Wx?�&?�͕>�{��Ǐ����)��<G�a���}�?�ig?�f���?%9�?�G??�rA?�af>�z��@׾����N�>B%?ګ�ūO�#�/��v��tY?��?�'�>�,����f\廻����ᾫ�?u9b?��$?A�ݾFV�����a�><���μ����<��~=�'<>��>S���p�=3��=7O�=D@�U���*:=��=��>:��=4���0=,?��G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>/�l���K���ڙ���F��]�Ž8]ڽ�S?)��>\8(?-S�>C'�=�A�>�'־e` ����:���%F�c.�s^G�J���7�Ѷ���^��=��Ϛ����o���>e���>���>⏂>�B`>d��><��<�2b>���=��p>��>��=��J>[u�=�Æ�k��<�KR?������'�c������.B?�ud?�"�>Xj�w�������?m��?�u�?�Xv>�mh� +�h?�>�>F���k
?�:=?
��<�N��`��B~��0�K��>96׽�:��M���f�Se
?F2?�����|̾l/׽C��� �=�U�?�+?��5��[��Fu��rO���S������W�v����&�j�Dc��-V������gf.��"�b�&?ܐ�?I�
��H���i����k�HdE��Ћ>���>�,W>�n�>�s>f����#��S��z-��傾���>m&e?��>�K?�Y(?jp6??�Z?;�>z	�>���d�5>Vb�F>�>p�?6�.?��6?��5?Q�:?WnN?n�X>�?��T��#��t�;?��
?��>�W�>���>	�Ž�>J>��~=[\d��"ɾ.�ҽ��<���=]�轟�\��'=�>�K?4e
��9��
�0~>�	=?��>��>�l�EYݽ�K�=���>!�>�D�>,Ѿ�Q]���x��>��?�^;��8=��>��=�'O��;��Un
>�V-��>I��=�����T9���=kݮ<,H罐ү���f�|��<�t�>6�?���>�C�>�@��0� �\���e�=�Y>S>a>�Eپ�}���$��o�g��]y>�w�?�z�?��f=��=��=�|���U�����D���:��<�?7J#?&XT?[��?q�=?^j#?е>+�eM���^�����Į?� ,?^��>���Ъʾ��3��?X?�;a�6���:)���¾sս=�>�Z/��1~�h��/D�J�����|~�����?Z��?K�@��6��t辊���vZ����C?��>�W�>,�>��)�q�g��#��,;>��>yR?�$�>��O?�8{?��[?ŏT>_�8�Z'��ҙ��q3��">S$@?U��?�ێ?�y? V�>Co>n�)��ྦ-���"��7�"ق���V=yZ>:��>� �>���>�>�=biǽ�l��T?�T��=Q�b>Xe�>۔�>d��>0Kw>O��<E�G?��>Q��=��+P�����ǒ1�9�u?��?��+?�= ��E�����Fj�>H/�?�Ы?��)?�SS���=��ּ�䷾3't����>v�>R^�>>A�==	@=�z>>��>BX�>f��g���{7�p9D��?��E?��=}�ƿ�u��0c��̙�~�;f����^��@�Ѧ@�ؠ�=JX��)6#������b�i���N�������������z����>�S=1F�=�%�=���;���:��<�;R=��,=��=L�|�9N�<u��2�㼱����N]�<Q_s=;y���b˾�}?JI?��+?X�C?�Cy>3&>߶5����>u&���?PBV>L�R�����f;������2����ؾY�׾6d�oǟ�ʊ>@�G���>FL3>��="N�<wc�=��r=�0�=~�Z�-�=�b�=e��=�%�=���=X�>��>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾr@?��>>�2������xb��-?���?�T�??�?=ti��d�>L���㎽�q�=K����=2>m��=v�2�S��>��J>���K��?����4�?��@��??�ዿϢϿ7a/>�Y>�(>�kY��78���;�oTo���)�Pw%?�1C�`����n�>u�>w�־&壾��=	I.>��=�/�"(R���=A�d�a�;�j�<֢>�g>O�=׸�;��=U
�<��='�m>�6�=����2�gв=Ȯ�=��`>v�K>|��>�?�Y0?@Ud?�C�>�	n���ξ�@���*�>@��=�8�>�ƅ=GB>7��>��7?��D?j�K?�m�>�=n��>� �>��,���m��a�_���!�<Ș�?�Ɇ? ͸>�R<�A���[>���ĽJ{?�X1?�o?"Ξ>[���ܿF�'��/��V#��\�<w#(=-�u��I&=H#l��욾Ս3�#�N>�:�>ί>Ϯ�>J)�>4K5>(LT>
Q�>kK�=d#�<'Tp=+=��=r:�Zf�<�Q�<�����&��3ڼ���=Y�q�3�%���m=�Z8=��=�����=!�>�?>��>�N�=1k��iG/>���L�L�1��=P����A�A~d��m~�~�.��`9��_A>PW>�����&z?��Z>A>iM�?�u?��!>���,*־����if���S�e޷=�>r�=��I;�%`��M��)Ѿh��>��>���>�Qm>��+��,?���w=�S��X5����>������ή��7q�"/������i�5�uyD?�8���a�=�~?ЕI?�ҏ?�y�>�֘��Oؾ^80>���\3=N�+(q��8����?'?z�>�)�1�D��̾�������>cVH���O�@���̂0�������}��> ���>Ѿ�T3��D���.�B��hr�u_�>X�O?Lۮ?7cb�}_��zO�ƨ��5����?��g?H՟>I?O?�����v���p	�=��n? ��?M;�?�|
>#�=
�_�&f?>?B��?�0�?��k?x��{+�>��=|/k>�8�&�=�d>�1�=Zv�={?Gk?1?U���P�	��>㾍6�"aI��<K�<��Y>4ؓ>䯖>ܓ=����(>�*�>�u>���>v�!>���>��u>-�ܽS��_9?jߢ=U�;7�<?�;>��>�N>q��p.M��Ջ�΁�=���*a��@>Y�|=�>�.ݽY;�>�����l�?J^�>	�6��?���d�&�е>�p�>[q��*�>m�>�v�5��~�>H�g>�Z=ށ�>�,�>8�Ҿ!)>���!��NC���R���Ҿ`{>���.?'�3S�1����I��Z��Z��MBj�P���3=��o�<��?���t�k���)�)��TZ?Қ�>�)6?Bf������)>�c�>4�>����d������ᾂ�?��?"<c>��>c�W?�?!�1��3��tZ�I�u��'A��e��`��፿x���Ж
�����_?X�x?gvA?a�<-:z>w��?V�%��Տ��*�>J/�%;��r<=V*�>1(���`���ӾջþB0�oJF>U�o?{%�?;Z?�UV�FNl��a'>H�:?~�1?�Wt?��1?��;?n@���$?��3>�M?(b?W95?�.?S�
?�F2>���=�W��Q�)=*���\튾æнKʽ�!����3=�<z=ۊK��e<�=Yy�<���׼��,;q��%��<�i9=���=��=Q�>+�]?�x�>ͯ�>�E8?�u��i7�� ����-?n�3=����ȉ��⡾2�D�>��j?�߫?�Z?F�e>�wB���B���>6*�>�-%>�\>�>I�!�B��ׇ=�>D~>8�=�R��;���R	�럐�N�<A�>�:�>�{}>Cᓽ��'>�*���&y��Jg>�WS��ݼ��V�B-G�T�0���t�I��>�L?7>?o]�=���2E��%�e�ݳ(?eu<?�;M?�f?��=M,ܾ:��J�ܮ���>���<�j��ޢ�-ơ�y�9�d�D;�t>/ў��f���rf>։�k�Jm�1]J�"V�l@d=x��}F:=Z��U]Ծ�ۀ��-�=��>�4���$!�n疿R����WI?3�t=����U�C���4>5�>dխ>O}7��>�@�5꨾!�=��>�8>t�`�̍�tjH��B�r�>��F?LW?vׇ?�uv�t�k�AC��<ġ�������?JE~>Ċ?�Y\>c��n�ؾ�b��'c�4;�Aq�>�%�>�"�l�Q�����x�=�����>w��>l�:>x?�;?A?w+[?�B?�.?�s>�]<����C&?m��? =�=vzս�fT��8��F��/�>�R)?��B�1�>�S?Ѡ?Z�&?v�Q?�?h�> �1!@�wt�>��>��W�F]���`>Z�J?]��>GY?n��?�=>�g5�����~��TK�=2o>��2?�T#?�?�ȸ>�?O�]��D����>�#�?�ށ?��x?��׼,�>.��>v�?���>z�>��'?H�+?G?
�~?yXF?ל"?�������u =A�ϼ$X�<�<Da�=���aY5<U�������=t>=h�߾9��>lT�W=_��s�>V�s>�0��Ҹ0>�fľ����_A>�v����������Q�9��Q�=cx�>�!?�ە>X##��'�=ɼ>Έ�>j���(?>�?7?�":;Ypb���ھ�L���>b�A?,��=ܹl�it����u�"h=��m?�g^?�W��
����b?^?����$=��þ)�b�p��?�O?��
?L$H�0ĳ>��~?��q?�~�>��e��#n�����Ab�:k�j¶=�}�>iH�6�d�$$�>N�7?�1�>D�b>M��=�l۾��w��;���)?T�?���?&��?M5*>��n��,࿫/������5e?� �>JL���#?�bc�0=Ӿ�ވ���}���ܾ}U��j���w��A���*�g����`̽ �q=��?#�v?��f?DZ?����j�c[��ew�p�V�������>D��E���@�,j�<	�����Ѩ��M=$��IkW�@v�?w�$?��ƾD�?�%���k���T^�>�'_����e�=�c�z8�=����ߜe�՘^�3{��ŭA?ȿ�>I��>��?��n���f�n�9����o龁�>/�>��E>�`>{y�,��+�=B��g�ھl q�@�w>Luc?P�J?�Xo?P� �]�0��Y��±!��x6�R*��{~G>y>���>IS���"�%�'�G>���r����T���9
�-k_=�/?Lŀ>h�>xؗ?ke?S
�	���;Yn���1�}xo<ɺ>|?k?���>g�>�Ȼ�3�=��>��l?��>�Y�>蕌�W!�W�{���˽j�>K׭>]��>��o>�t,�\�~������?9����=ɓh?Í��̤`��؅>��Q?M<�:�I<�;�>�Hw�P�!�'��y
'��>��?���=��;>�ž�,���{�o!���[)?S&?��&�*��$�>�4"?��>���>e��?D�>`����A;t?�%_?�PJ?��@?eK�>��#=�⫽��ʽ��&��/=�(�>b�\>�Is=J��=�M���[�] ��
9=�˽=ټ�a��(W<�����L<$�<�74>ۿ�aK�A�־BU�8��!}	�R��ҵ�Sl�������Q���;w����Qn$�$pW���e�ES��uo��k�?".�?#:��?����]���������-�>8Ct�X����"���k��疾[��?��A� ��P�egi��ue�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >ZC�<�,����뾭����οA�����^?���>��/��o��>ޥ�>�X>�Hq>����螾t1�<��?7�-?��>Îr�1�ɿc����¤<���?0�@ܢA?�$#�jw����4=5��>�t	?��F>G� ���!�b��s��>��?mڈ?��=1L�>Z+�x�g?�=�:�n���Sq�=3��=���<b�ͽ�o>�y�>�Y)�,>�H,���i>�>��c����f�S���<��v>D����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=v6�뉤�{���&V�|��=[��>c�>,������O��I��V��=����p�ƿ�b�	��t��=�s�=\^�����Hg�%�Q=�b��3`��Ou=^An:�M�=��;���D>���>0ل>��\?�d?{�?yR5>�ݽK�5e�Y��S������A����׽�"ľ37��V\ľ��#��;K�!��D�V�پ�>Gh�ː�ľo�o��g2�&�h?��>R�(�l%P�Tu]�W�*��(����=�Z6<|�	�؞��Z�̫x?&h_?[(`�t�5p�����D�� .(?�0>���@>ƾ�`�>��=ji�=���>��><�p��G��H�01?}�?`ξ�<����g>�o����=W#?Y�>���<O��>0/?�&��0�\�>��*>`�>���>yME>�F��>ڽ-�?R�M?�-���P���!�>�'Ͼ��r�v)=�X�=��^�d�T�]>���<�NT���*��UŽ�j*<T�U?�S�>V�5�ao�!XQ�v�9:���=7�n?�³>���>�{�?�B?#�q=�1��M�-�����.>�Z?��k?sh�=�I���ϾD��E�D?Jfx?�ew>�΀�[3ܾ3�2�/&���/?�$M?5�?Aj�:�)g��{n�ʻ�h&J?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������8�=wӖ���?~�?|�����<{����k�5���Eu�<�w�==w��N!������6�D�ƾ�j��ޜ������>u;@O������>��8� v��ο?����ZҾAv�+�?���>��̽���]Ij���s�./I�tI��ڋ�2�>>uF>�����,���[���,�*��u��>'#�rb�>t<�2���:\���=�D�>��>��@>o7V�Ó�̹�?'�R̿j ���ȿ�=�Q?�^�?��?,��>���<Y=���א�g���0M?I��?�ua?P	>w3r=b�=%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*�~�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?�$�>��?�l�=Ta�>�f�=�𰾇�,��k#>� �=j�>���?��M?�K�>.Y�=��8�B/��ZF��GR��#�;�C���>i�a?��L?�Kb>o��Y2��!��uͽ�c1��W��V@��,�	�߽=(5>��=>>��D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>B�Խ����\�����7>1�B?Y��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?]Qo���i�B>��?"������L��f?�
@u@a�^?*�hֿ����_N��P�����=���=׆2>	�ٽ*_�=��7=��8�A=�����=s�>��d>"q>;(O>�a;>��)>���Q�!�r��\���S�C�������Z�C��Xv�Xz��3�������?���3ýy���Q�2&�)?`���=\�U?MR?Yp?�� ?��x�k�>Z����8=E�#�̈́=�/�>�h2?�L?q�*?�ד=R���,�d��`��6B��ɇ�!��>�rI>��>�J�>�%�>5�M9��I>A1?>��>c� >�f'=��X`=�N>N�>���>D|�>���>᭬>@ԟ�M���<�Q����^�H�Kq�?oΞ�����]��1��;�G���� 2?8�>�Ȅ�C�̿C�����$?^n�t����<�o����>�Y?�*>&�=�>f;�ٽ�[�>}�Y����,��=2N?���>�O�>�(��L>�uL�o�����>�H?���g]��I����*����q��=#U�>�=T����ۋy�4c���q���0?��#?�b~������I��5���6e>`��>�(�L)n�_��>��k=M��o��m�<Z~�<�o�>{�?��,>xـ=ʻ�>N�����G�O_�>7�@>ӳ!>�_??�&?��ּ�ڒ��Yz�!&��uu>]Q�>�j�>>*>��N��e�=���>�_>8:м�l��
	��D���W>CӁ�Jif��=`�m�i=fY�����=��=�N����<�nr1=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ&l�>�k��Y�������u�է#=8��>u8H?>`���yO���=�Ro
?�?zK�X���k�ȿ�uv����>��?��?�m�|A���@����>\��??gY?jxi>n۾v_Z����>��@?jR?�$�>P/�x'�F�?�߶?���?�-V>ل�?c�m?;:?ω��n�)����Z���[�T=W<�7�>��t=���ҍ!�k���蠏���S���'�)u7>\0�<U"�>��
�Nվ��>����&˾Eؼ�{9>�R^>��>�[�>I�?���>?�>)��8�����9Z���K?�ŏ?D�7o��T�<(��=��`���?!75?>��m�Ѿ"R�>׍[?�l?E�Z?x2�>����S��n���� ���<�#M>L�>�8�>劋�WK>/�Ӿm,D�tD�>B�>Y�v�W-ھ.�������t�>�� ?�b�>f\�=� ?�6%?�!d>�^�>�b?�=���E�V��>���>�?`�?�?`��$$)�{���6��Y�Y���:>�s?�K?n��>)��n枿4�N-��
O�䴇? W?0Ʈ��E?�'�?��5?x�A?F	�>'�1�Ͼ^�ȼߊ�>e�!?��,�A��(�<,��?�%?]�>��|�~��t��de�����x1?߯[?�&?S����a��ž�f�<�9����85��;�=���^><�>㧇�T�=i�>���=b�c��4�f�f<=��=>��>=��=�f<��p��(=,?�G�Zۃ�q�=��r�<xD���>hIL>�����^?�l=��{�����x��
U�� �?��?;k�?{��Q�h��$=?�?U	?�"�>�J��5~޾���KQw��}x�Aw���>(��>u�l���Z���ș���F��;�ŽH��K�>$��>�`?[ ?%4O>0�>㧙�G'��B����1�^��=�88�,/��������1�#�{���K¾�^{��)�>���|C�>J�
?g>~{>p�>Ϩʻw��>�sR>�7�>_u�>."X>�3>>� >�c!<��Ͻ�CR? ���(�E��\ɮ�WKB?�_d?���>�1u�Y*�������?7�?���?ʽw>�%h���)�1�?�j�>�����
?}�<=���ߑ�<�ݵ�������2C�Yۍ>^�ݽO@9��M�{je��<
?$R?����y�̾��Խz���QL<��?��&?�J�-�:�}z��@���O���ѻ'gt�l���&�CQi��s���:i�uR��*�"��5�'�A?�{�?��:��P�^)��/��Ŏ̾�>-��>��»�!h>���9*���[�UNc��������9	�>�|�?�Ω>L�5?*`/?\'?��{?�?h��>�S
���>�f{>�i�>ն?�?D?��C?_`?��F??�w?�<�>|�>�-��(��,!?,K�>qa�>�#�>Pp>M�%����>>�Ž���]�'>��y��`�!�����=.�=�#>��?{��h9��r��Nyq>��7?@k�>>@�>����k�7�=��>�
?�!�>���S�q�=��/��>��?B=����<�*>�k�=���3�;=��=MA��C�=#2fd���u<<
�=PO�=(�!؉;�;��:2��<�t�>/�?���>�C�>�@��2� �P���f�=�Y>�S>@>$Fپ�}���$��o�g��]y>�w�?�z�?��f=��=З�=4}���U��}��n���&��<��?IJ#?XT?V��?p�=??j#?��>�*�fM���^�������?m8,?��>���W�ɾ�򨿏�3�?l?*`�KK�z�)���¾p3ٽg�>�#/��}��Я���D�����y�}ޜ�LC�?0�?�A�`�5��
�Ș����vC?��>��>ܫ�>��(��hh�����;>���>�!R?p&�>��O?�{?7\?�S>x~8�O��%䙿��8�E�!>�@?EX�?��?��x?��>c�>\	*���[������ ��7]��y�M=�kZ>���>`]�>���>�U�=D"ǽ℩��0?���=֭b>D��>��>y��>|iy>.�<��G?R��>e���G��p��0���"�<��u?��?a�+?�X ==y�=ZE�������>��?]��?�*?�R���=7)}���t���>Ѻ>���>�Ɣ=��?=N>G�>���>���G����7���F�R�?bF?9��=�3ÿ��x�:ԯ�/�~�>�=X��ꞑ�2W��"�����=���XE��%�t�l�o�i��<�۾O���{�q������!?t~�=��e>	->����޷=1�_�c��<�ټ�<籦=���<�m����P='�Ӽ�5<��=;�B=n+�0�˾��}?�;I?ޕ+?��C?)�y>);>��3�S��>�����@?qV>=�P� ���{�;�K���� ��S�ؾ!x׾�c�ʟ��H>�`I�%�>�83>�G�=�K�<1�=�s=�=��Q��=$�=�O�=og�=��=��>MU>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�<>��>��R�H�3�æX�ySk��_�	�"?�z6�i�о��>dW�=��߾�ɾăB=@�=>�'P=b� �<f\�ZՖ=����tJ=c�b=���>d�?>�ӻ=/k����=_�.=r��=�sZ>�¢�\o0��F(�"�F=���=]*X>�k>���>�??�/?id?��>�~m���ξ�,�����>���=���>��=�pC>3��>��7?D?%�K?�Ĳ>��=}�>C�>��,���m�u�7���J�<|�?4G�?�M�>F�k<M	=���'d=�la����?��1?�	?��>o������.�x�(����gZ.��uJ>fs�����5Ef=V�`�%�X����>�[ >yT�>zm�>�3N>C��>���>���>��A=�X	�v��=o;����T=2�T=��j;G�̼S�>�/����B�=`=����'�2������<�+���U�=�%> x�>��/>B�?e�"=Ds����1>AQ��h6�W�=�i����L��JX��5g��L��M��O>�a�=�<��w���H?J�l>��P>���?]4o?�=,�x��H���t���ד�r\���E>�Z>��n���V��T�*�=���þ���>�>��>Ifm>�,�� ?��x=+�LE5�^ �>:~��6���#�jq�FN�����h������D?*J����='~?>�I?��?��>x:����ؾ��/>1��h�=x���|p������?��&?�|�>W���D�4$��PV���)�>�G0��:P������J!�f5=�����c�>/s��Qj�]}:�v���d���*1�-�`�>��>?GE�?�.������R��Bپ�c	���?v?�R�>4u�>}��>(����������1�=tc?i��?Fm�?�V>�g�=w���Ǭ�>�O?���?�n�?�uq?*;����>�{�<ݶ6>�)�����=�U>L�=b��=��?��?��?K]���Y�X���G�S�N��;=F��=B<�>�ȇ>��l>���=I�=���=%\>xy�>Gl�>��s>�0�>䛍>��Ⱦ�Q��/<?�">�@W>B?]�2>�N����Ϗ=g�,<4+�ҥ���ՠ�!�����p�;�^�=�X�����>-ٓ?�a>�v"�>?�w�Ȑ(�9x�>W�~><6�ZM�>'	">�Wg>���>Ĩ�>�M>��>3�=��Ҿ��>�U�f� ��uC�.-R�jѾN{>�ޜ���&�ԣ��-���J����&���Di�X���<���<�J�?����l�� *����4S?Zu�>��6?����ň��R�>���>~�>uX���M��0T��n�����?���?R�c>)��>��U?+�?ܫ2��5�&�X���r��@�0e�(�`�ZL��
���*�5yƽ�=_?�*v?��@?���<47|>H�?�V'�s������>"0�~G:�y�W=�b�>�Y���.`��ӾȊƾP���gL>Яm?Ͻ�?��?;�R��Zm��#'>Q�:?J�1?�Tt?��1?��;?�����$?�t3>nI?�x?�I5?�.?0�
?!2>�6�=m'���M(=�e��}]xѽ�oʽ����3=�z{=P�4���
<��=|��<���?ټ�I;�$���߫<�:=�=��=Mɦ>�]?�q�>���>��7?,���58���!$/? +>=]�������䡾Y��R>k?�?�pZ?_�d>C���C��d>V�>[[&>��[>�0�>4���C�j��=O> �>�å=7�R�&����	��L�� �<4�>,/?='�>Pb+��G�>G1�@��C^�>*����нoh�iZ��=N��¦�W�>�m�>#E#?���<�<���ν����	?!2?o|?��s?�o>���οb��9��[���� ?B��u���tu�D���ВU�E��=z�>��:��Z���*�>����/�rk�T�M�����j�=�Z��=������ҾA���ѫ8=�$!>�����$�d���#��pE?�D�=���ޜu�Q��x
>5,�>��>O����z�}�E��]�����=��>pm1>ա
<@���m�K���
��u�>�-F??r?�4�?O���[t��fL�r��w���q���l[?&�>���>xP]>7�<��ɾH�xi��	E���>��>����K�G2���P׾>O�P�>���>R�!>�?j�P?i?�pN?��?_?y]�>S�c����0j&?VK�?�	�=�ӽ3�U���8�>D�[�>F#(?�?����>֪?��?�'?�P?eI?�>�����O?�x�>��>I�X�����\�f>�;K?:F�>��W?�P�?�N>>:4�8/������=]=>�[2?�_$?0U?��>��	?*f��k�<;�T>�8d?�Ao?��@?�#=�j�>��d>��?��>V��>Yr?S|?�l?�{v?�G?�?Nw<~1��B��<b��=���=��<h6��Q=|C���R뻺,�=A�>E=�h��V0�<6w�<�+�=��J�bk�<u��>st>�}��[0>LXľU ����A>S5��n����H���C9�쇷=A�>o?�<�>�#�盔=�ܼ>"v�>$���
(?��?|�?��;�$b���ھ.L����>��A?��=7�l�Bo���u�`
g=�m?g�^?^UW�����b?�H^?O4���=��ľ4we�����CP?ޔ
?ީM�G��>AI~?$�p?��>�b�0�m�������b�`�n��X�=���>���f9e� ��>0�6?u��>�z^>0��=_�ھO=x��ϝ�?�ˌ??
��?]�&>�o�l�]����Z���<c?�;�>q��}l#?��ĻBIپ�9[��UO��Q��X��Y��g��ت����ʄ�����A>��?~~?qbi?B�a?�@�L�z���Y�da��ww[�?�� <�Q{D�)�7��G�8w����k��D]�����[�����S���?&?�FH�Nc?����ٗ�ͮ��Q�p>��þ�=޽f�=��<(6�=R>LYX�O��]�T��=)?y��>���>�eA?�,a��eJ�K�+�OJ��=���l>��> �i>Ⱦ�>�X��N��B�#�a�=MB��y>���y>c?�S?ǆu?��ú3�ń��;#��p��tբ�0�.>\��==�>�@�	.��,� C��t�B��q狾�����=�T*?�Yl>DT�>�ؗ?��?i*	�����9�I���)����<���>�\_?̻�>
��>����/w��D�>9�k?z/�>�>ߕ��*�#��~}�nڽm��>2�>-��>�O>R-;�o�W��������[I;��&�=yc?5���	]����>�R?Ї�<� �;�f�>%:���5 �+��JT�eK>@�?J��=7�:>�JȾoL�^w�{g���)?�?�4����*�� �>�$?��>��>���?I��>Y����N=�m?E�\?�hK?��H?��>&�~=��k�_����%���X=F��>�?K>��S=M��=�
��h��=���ɋ=���=O�i��;���4O<��:K0�<ٹ�<�b?>�SڿоJ�_EվI�3����]
��<��)����C���� ��E������ov�f��K>A�ݝV�a�e�Ge���l�eK�?���?*��9U��G����΁��L��_��>�(x�dߋ�?����i|���=�D����!���O�a"j���g�X�'?`���޽ǿడ��:ܾ! ?�A ?�y?���"���8�ȭ >C�<+����뾚�����ο.�����^?t��>���0��$��>��>��X>�Hq>����螾>5�<��?&�-?3��>B�r��ɿO����ɤ<���?'�@��??���H)⾎�%=t�?�k	?�{>������7�ǙC��	?�#�?6,�?:d�=)7T��l�<e�o?v	>pm���x�D�=�)�=�����<f�>+��>ó2�v��G۽?G>�<�>�	�<s�T����2�;M	�>�<�Z��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=@����"ſS#�8�)���<�o=�*�,�ѽM~�g=D��1��XcY�顥�*(=7�=� E>���>�Nt>��d>�-O?m,^?Ĺ>uZ>�qԽ�W����Ӿ-�
�#t�.�p��6uB�@��� +ɾiq�����6���11��L�}pr>a�_��w�ە��\n��1�ϥh?k�*>c�3�<A>�m�"���"���"���=��.�#K���9�1}�t��?��I?��j�
<p��Ⱦsyz��'���0?~j㼠����:q�>)�<>ֆ=���>��">��8�a�"�w�M�0?M ?�=���ɐ��u0>������$=��)?���>j��<i��>>�$?��'��ؽ�"X>m�6>B��>�#�>[�>5﮾S�ؽ�R?��T?�M��暾a��>t����J��jI]=�K>#-0�,���Z>ȱ�<��������1��3ɶ<OW?�9�>W(*�/@��͐�,�;�w�=lr?��>Ɍ�>�k?�2=?#�%=T���FP�+�a��=�.V?��f?z]>L����\޾ϋ���q??�
i?ЏJ>Ytv��&�wD*�����/�?8Cq?�Y?R���qtw�����������7?��v?�r^�js�������V��=�>\�>���>��9��k�>%�>?g#��G�������Y4�Þ?��@���?��;<� �'��=�;?g\�>�O��>ƾ�z������g�q=�"�>���ev����R,�b�8?ؠ�?h��>�������z�=t����J�?�t�?��Ҿ�Z�����vl������>�?T<��&�����hԾC4A�����=%��!��R���G#�>a@J(�#�>���I��ſ�dh��x ��`��-�?rH>y�+�=�si�o�{�\I�I:]�{��O6�>{�G>�Ƚ�����9�B���=!?��ѽ�8h>������SbǾ�ꐽ��4>�1�>��>|x�������?�Ⱦ�,ֿ/p��q����M?�^�?���?�<?�� nŽO�S��Ѽ�?�3v?E�=?���=���D�<$�j?�_��xU`��4�dHE��U>�"3?�B�>V�-�ײ|=�>���>0g>�#/�w�Ŀ�ٶ�"���Y��?��?�o���>m��?qs+?�i�	8���[����*���+��<A?�2>���H�!�<0=�QҒ�ļ
?X~0?{�`.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>kH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�$�>��?�n�=Gb�>�a�=����,�|k#>� �=#�>�}�?�M?K�>�V�=�8��/�8[F��GR�q$�K�C���>��a?<�L?iLb>����#2��!��tͽrb1��S�?X@���,�a�߽h'5>�=>y>`�D��
Ӿ�U?���SyؿPh����&�V4?L\�>��?C��t�5��W_?�>��
'�����f� ���?H��?��?�e׾�ϼ�6>��>D\�>�ս2Y��q�����7>*UB?u��u&����o��j�>��?��@c��?2�h��	?���P��Wa~����7����=��7?�0��z>���>��=�nv�ۻ��Z�s����>�B�?�{�?��>�l?��o�M�B�_�1=7M�>ʜk?�s?TRo���f�B>��?#������L��f?	�
@~u@^�^?'HpͿ	��N����Gþ�Ķ=�#�=VvV>3vӽ��>ޞ�=��6=������=~P�>�^=>�E>>ё@>�iE>;�U>���)�&�����	����7>�u���� {�� ��_�5% �����z|���8���ｶs�UAF��b�h:��~��=H�U?7R?�p?�� ?s�x�O�>$����(=m~#�΄=�.�>Gh2?�L?��*?@Փ=	�����d�:`���A���ȇ���>qI>;��>
K�>�$�>�dJ9��I>�0?>���>�>1n'=�店\=]�N>:N�>���>|�>(��>ּ�>�&�����q[�*���þ�Y�?2�g��=���J���6J��e��1v;�5�!?R`>�Қ�5�οr_����&?�㤾;��2���"k���	?�[?���=vG�����=9�=�7�W�iC�>@c:��ւ�rU��S�>lm�>���>�Z�>s2��)�Bt\����<u>��7?��ʾ
�������>�<���>/�>��½��,��F���ˋ�1�|�0=_�56?��'?���&�n��+ý�����>9�>�I���5�֣^>��l<��1�^���l>Ϧ�=P��>:K?�!6>��,=Ա�>͂��?�Xش>��>AO�=�@?B+?ؼ��A�ae�Ō9�<{�>$w�>�>�B>ҚO��\�={��>�!^>��<g{���9�N�l�?>�:����P���<�{=�:��
x�=e�=vY���/��t:=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿԭ�>Ѡ����������t�#�=�,�>�F?����,�(�d�3�
 ?��?���u+��)�ƿL�s���><h�?!Y�?�m�~5���B�$�>[w�?A�W?G�]>Iھ\�U�%��>��@?�\T?�ڷ>�C���$���?�Ƕ?�ʅ?Z2Y>��?P��?ì?��~��=�������E�ѻ[
�<��>�C\ƾ5��E����������%�P�!>�'<��>�F:�����җ=�*.�L���9h���j>�3?>A͸>�έ>�?*�>�U>�l%>�ĽIt�Q�����K?���?���3n�A$�<ዜ=p�^�'?1H4?5:\�x�ϾuԨ>M�\?���?�[?^c�>���v>���迿�|����<��K>�3�>�D�>o#���MK>��Ծ�7D��r�>�Η>����@ھ(�������>�>�d!?R��>�Ү=� ?׈#?��i>s��>��E����ϨB��f�>׍�>��?��}?[?Ǻ�Jm2�����������Z�ML>x>w?��?�ד>�h��$������m5��������?e�f?�%�k�?9��?s�??�@?�k>f���Ҿ�֘�wO�>��!?ŀ�|�A��S&�s�sN?A)?&��>wb��k�ֽ�|ؼQ�������?\?/&?6��P-a��;þ��<LN%�6�U�0g <s�C�k�>k�>ӈ���=�V>L��=�2m��]6�Ôl<`�=�n�>�:�=��6��n��.=,?3�G��ۃ��=��r�CxD���>GJL>����^?�l=��{�����x��	U�� �?��?Lk�?���2�h��$=?�?>	?�"�>�J�� ~޾2��rPw�[~x��w���>���>!�l���C���љ���F����Ž�s�`_�>i3�>�K?���>�?>��>𧻓�<�%��Y���Oa��/���6���-�o��ꞥ�]�+��Z��ľ��v�Q��>ӣ���@�>�*? NU>r>F��>�QW��>YO>�H�>
p�>QFY>�,>f[�=}#<GVʽ�KR?����	�'����웰��!B?�{d?��>>j�w��7���r?��?
q�?|v>�nh�i+�dq?@D�>d���a
? �8=�r��K�<i	���������J�֠�>��ֽ�:�f�L��Mf��Y
?�*?=���j̾��ֽ�d��^�=7J?^3?uCD��T[�"t��&A��O�,b"=p�{�
�ʾU!��Sn�ا���V{��(��c+���ּB55?�?�}'�����픾��|����pO�>w��>>6�<���>nQ�,<��W�"�=��#���x)�>�F?�8�>|�C?\�9?�.M?sa?y��>fД>���0z�>o`�<=��>|!�>^4C?7b"?��-?�%'?��6?�>��� ���ξKI?�?\�
?ҽ�>���>Q�v�"Ɛ���[�����m�a�����*<=D�>@���kex��+=��=>9�?�Ó:�=��k(t>��5?>��>5��>bl���s��#(=��>�?���>�� ���n�`&���>�X�?>��1=X>#>��=h}<<�0<���=���
�=�����]`<�	�=�$�='uϻ�&<��<�O;4!�<�u�>
�?$��>�A�>�.��!� �����7�=�X>�*S>j(>3پaz���#����g�A]y>�x�?O{�?B�f=��=߈�=�u���U�����x齾�W�<ޢ?R#?~ST?蔒?�=?yj#?�>?,�[L��R^�����{�?]�-?�O�>�𾛿M��F��ǋ;�n+?��>/�T�Q|���4G�	n쾜�_��`�=?V/�#����Q�Yʽ����<���?DԨ?z�=�2#�~q	�Dٖ�%9b�K�@?�>�=>3H�>&{��bZ���8��
�=փ�>ei?'�>��O?�{?s�[?c�T>;i8�>,���Й�[D���!>��??�d�?�ʎ?��x?���>��>��*���߾����$o�q��i���4�S=�FX>qs�>%h�>�\�>@��=`(ȽBV���}>�x�=�b>�^�>|�>34�>xw>���<�+H? ��> ������/G��?ޅ�b�T��^p?gH�?#�,?F8T=����=�p���4�>k9�?�ߨ?�M)?QEG����=�jNƾ,�����>#�>D$�>
�[=M4=:^>���>3��>�߽,���3���=��G?
~H?���=7CƿZ~v����W����K�;-f��&8� �P�M�4����=��������ė���h� d���_�� ��2ㇾA1e�<m�>	x{=�m�=�"�=���;��̼��;�(=��;{I=Z����Uż�q�ץ޼�������<t�=c�Q=�h�0�˾��}?�;I?ޕ+?��C?(�y>*;>��3�R��>�����@?qV><�P� ���{�;�K���� ��R�ؾ x׾�c�ʟ��H>�`I�'�>�83>�G�=�K�</�=�s=�=y�Q��=$�=�O�=pg�=��=��>NU>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>b0;>wB	>sS���1��z\�=�f�4:^�1K!?�l:�P{ξ��>m�=<�޾l�Ǿ#�1=ʺ6>T`P=Ja�$�\�7�=��~�� 6=h�d=NM�>/ZD>'߼=ȭ�����=8P=[��=f�N>� ửm(�7�3��~7=���=��c>�1#>��>	�?xd0?0>d?> m�i�ξ���̥�>̷�==��>(��=�uC>Md�>V�7?��D?��K?��>ۨ�=��>슦>el,��m���侻O�����<!n�?ָ�?Y��>RS<�QA��7��&>���½gN?�@1?�i?K�>�>���̿V�%�xG���P<lڌ>"�->�O���Y�>	�<x���O�=�Sx>���>?? >�>�zU>��>�w�>��@=�U�=�բ=#�콦L�`_<��=>���=��=�6�l=����ߘ<��<��;�4���B��l�=��=�6�>J;>$#�>�҄=QV���G1>�N����J��=pk���F��cg�����-�V)C�~7>DHP>���K����j?�lS>N67>h�?mr?�>�p��;����NEb��$L�t�=0O>��/�-;���^�{K���Ҿk��>.�>�
�>~��>d~)���B�)��<��q*0��f�>ɔ��2࿽٧2�c�g��ҡ��!����j��)��%:?9Ç��m�=P��?��K?L�?)n�>[�l�!�'>�6���ȃ=$v��L�ۇ㼃?+`?���>����7�u}��I�b���>���0�Q�!񑿘��N�9<��ξ̰>������-�:�k�ZŔ�^|8��o��%+�>��4?���?��qՎ�c�b��������Z�.?��k?��>)�?� ?��1����JUs��s�=�-|?�{�?�l�?�oi>�r>�����?J<?N�?���?;	g?b��n1�>[Q;=!�>8η=�>��< �$���Q>��?��8?��?�#�c~��}��.n���es���
=}TX�(�m>��?)�=)���z����3>z�~>D?�>)u�=�&�>�ʕ>zbľ@k�E�?C��=m�k>��6?Iю>i>�/�<
ɒ=��L��V�)��2�?@�����=;��<�3
= dm=�:�>�6��Lړ?nc>�
���?��J̽G6>�H>>JG�:/�>e:B>b�>�s>���>e�=���>ޟY>x?Ӿ��>���a!�e-C�a�R�6�Ѿ_�z>���Y&�j�������BI��k���f�	j�[-��2:=���<�F�?"�����k���)�|���F�?i^�>�6?�،��
����>���>
ˍ>�F��ȍ���ƍ��\���?���?">c>��>��W?+�?�1��,3��uZ���u�G(A��e���`�㍿.���X�
�R*���_?��x?�qA?��<�Dz>&��?��%�'֏�0�>Z/�1;��==�*�>+C����`�
�Ӿx�þ�[��UF>?�o?�"�?V?B[V��&O�ȓ">
�:?@/?c1s?�u2?�a9?�
���$?��2>8?�?�5?��.?��?��<>��=�3;/iI=dP��nӊ�F|̽�9��P��(�'=^[�=�E�;z�;�&=F��<.����r;��
<<�l>=@�=
s�=_�>�U?�-�> ��>J�Z?٣ۼz�$��X�I��>�>������T��=E���㾏��<��e?�u�?�mf?�ߒ>�?n� ?E���h>�>>o�!>c��>�}�>��Ƚ��);�[\=Qt>��O>�>�S���� �UϘ���$>�%&>���>zm|>N-��"(>����Djz�D�d>��Q��ﺾɆS���G���1�ڛv�WG�>��K?g�?�]�=�i�݁���Df��)?8X<?-ZM?*�?-��=�ܾv�9�Y�J�9��z��>��<{��Ʀ�����)�:�\�:̸s>��栾�8b>��� s޾Q�n�hJ�����lM=�}��DV=r��־�I����=�'
>q����� �h��_ת��1J?��j=Zg���KU��h����>��>�ڮ>#�:���v���@�i�����=%��>��:>Fr��Q��wG��5���>t�D?f�^?Ճ?h郾�s�>�B�����褾����p?�g�>�?	+>>Λ�=ڂ�����t�e���E��i�>��>M,��G�y��\+�:�#��>/�?K�>@�?g&T?n?s�b?�S+?��?�Ǐ>o������0e&?��?��c=�;߽��M��T8��_D�p�>��'?l$C���>gD?-_?��&?Q?�?�7>���>.@�崓>hΌ>��W�a���\rj>��J?�5�>3X?s߃?FU>>�^7�����Z%�����=�>B�3?��"?�T?ᴷ>Q$�>E����<���>��I?�V?a�h?�͟=���>���=-+�>\P>���>�
�>�='?(�K?Xv?J?B��>��)���D��v���.弍v�=�)�&���y׮�>f�:2_�;P��=�l��(�M��ː=�r�=
�.>Q�~���>�d|>㧤�L�d>@����͑����>Y�!��pԾ�y���۸��g>>D�>�*?V��>%��I�>�>'��>2"�'?��?xq0?ȉ�ͯ]�!���u�Y��T�>��+?���=��n�����ǭo�Ȫ<��a?��l?	�����ܾ�Sg?qK?l|��?��ޟ��pǾKd��H3?R6�>2Aག�?Gdv?Rrg?4F�>ݡ;�S�I�������r���ž���=��>x�>��\���(?&�R?��>�R>��>�-�����*Rg�~A3?@�?��?-(�?RL�=�r@�\��v��0_��_q?I�>��Ҿ��;?D�Q�[��ݾ���ْ�+0
�#���ŵ���e��K�����B�vU��D��������-?��k?Ð?I�b?�/��35���j�k�|�;gB��(��3=��q�lJv�}%���E�.��T����������0���(a�8��?�?dJ���?�)���PR��FҾ��d>7"ھ�Q���s� �<�L���؅�=�ؾ�Ԓ��㚾��+?�,�>��M>f�/?4cp�>�V��M*�V�?��Z���>>e�>16>1�?��]�"����{=�^�������{=Ev>�Qc?�lK?5un?���R[1�W����~!�V�3�M���Z�B>�
>'��>ZY�����&�	,>��s�-��oN��G�	�T`�=A�2?�:�>$S�>DP�?:r?��	�R��#Vv�``1����<���>�;i?���>,��>�н�� ����>{�a?�o�>x��wξ�?�e������=��?0�?4�>��h�M鈿�쟿�����.>�/�#>Ī�?�Hb�����ǀi>�Fj?1<L����>���cgH��o����W=�]m>
��>2N�<���>f�+����ޛ���Ӿ��)?�
?��Ծ%)/���>C?�>��>L^n?�>6_þ���<:�?�U?_�??+�N?��>\_=��;�ý l��L�<~�>��">ߪD=�R->~�Bm����+���=ә>���tׁ�4<��H���5��0�=3yL>Q�ݿ�S���˾����^���F��/��R4�$m��L�������Ր�wec�����(��<O�Wa�hE��c�x�g��?�X�??�?���n�+���<�l�cx��*�>�zr��å�´¾H�+�*���ts�4��~�&��T��j�7�p�Q�'?�����ǿ񰡿�:ܾ3! ?�A ?3�y?��5�"���8�!� >�C�<�,����뾪����ο?�����^?���>��/��t��>ץ�>�X>�Hq>����螾G1�<��?7�-?��>��r�/�ɿc����¤<���?/�@"oC?f����6�s=s<?��>|�\>�eO�_�2�s���}7�>Ǜ?@2�?|�>p�>�5�����V?�J��a�N��f@�%��=�Q=>14*>$�k��>���>����Gi���mv>P�b>�%ӼH<�u\Y�Z�D�!��>���wO/�2Մ?%{\��f���/��T���T>��T?+�>o:�=��,?Q7H�\}Ͽ	�\��*a?�0�?���?)�(?-ۿ��ؚ>��ܾ~�M?XD6?���>�d&��t�ƅ�=�4� ���}���&V����=J��>C�>��,�����O��I�����=�V���˿j��݀(����:dh=Q��
5K<,�{����9����@��넽ۧ=���=o�a>:�}>v�s>z�1>b�e?��h?�B
?˨7>` ���ܽ�9��fb�f�t�h�(�oþ�&�Ʈ���d�@�Z� ��6�Ro�p =���=77R�d����� �g�b�j�F���.?{v$>�ʾg�M�I�-<�oʾ����ۄ��ޥ��-̾)�1�B"n�*͟?��A?������V���sM�W���ޮW?:N���	쬾���=����Z�=�%�>���=`��b 3��~S���3?+w?�辵 ����>��q=�6?�:�>�x<O�>��(?[���xѼ��l>�CE>K#�>u1�>^f-=�����
�<V'?|I`?U�� ��#�>`���G&��0<�sP>
�$��`׻��T>ZT�<ǩ��A�=������J=�T?<w�>�l,����t���w/Q��g�=2�|?|C?£>�h?��<?[rT<d��t7N�d���Q�=�U?j�m?��=`�̽��Ͼ����Os2?I�`?��@>��>����>/�o���L?�e?ޕ?�M[��F|�γ��}b�H�6?��v?s^�xs�����L�V�c=�>�[�>���>��9��k�>�>?�#��G������xY4�%Þ?��@���?M�;< �>��=�;?j\�>��O��>ƾ�z�������q=�"�>���}ev����R,�e�8?۠�?���>������.n�=����/(�?:�?�p�O�b=}���C����j�=��=��@��ޔ�i���D������(�?ǐ��k5=��>*�@�Qc����>�
�������̿RΆ�s�s��'?���>���׀ž�3��Pyj�16��=�7	߽�W�> �>�䔽���{�{�nv;�<�����>KQ��!�>�TS���Ŏ����5<���>���>�ǆ>�P���Ͻ�/��?;Z��a<ο���������X?�]�?�q�?�o?�]6<�v�O{�|��i,G?��s?h%Z?�&�;]�Ai8� �j?�_��oU`��4�uHE��U>�"3?�B�>T�-�Ʋ|=�>v��>�f>�#/�x�Ŀ�ٶ�7���O��?��?�o�	��>o��?ws+?�i�8��z[����*� ,��<A?�2>���>�!�40=�=Ғ���
?Q~0?8{�i.�]�_?*�a�N�p���-��ƽ�ۡ>��0�f\�N�����Xe����@y����?M^�?i�?Ե�� #�f6%?�>d����8Ǿ��<���>�(�>*N>iH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?/:�>Ȅ?���=q�>�Z�=Z���mP���\!><%�=hE��@?bWM?dH�>��=$�7�}.��+D��PR�����C�Dχ>��b?-�M?��^>������"��s!�4F���}2�'����C���2����HI3>B�?>>�I�<oѾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?lQo���i�B>��?"������L��f?�
@u@a�^?*m��C����ξX�˾9}�={N�=@>�ս�B{=�j�<ƚy<�W��ca�<[�u>z�O> ��>鍕>T �>ٟM>p=��K�)�8ޞ��ȋ�
�;����� �мk�@J
�RT��\�&�Aj̾2~���y����J���%ћ��6��`ߦ�!��=��N?3$I?�׃?)A?E=�y>�F�I��=�~�/i(<���>b�=?�P?��,?`V3=��2i��i��o��N�]�G��>�m�=uڪ>�T�>Y�>�Ǽ{��>�W<Hz7>!ԍ>ChU=�����=���=�Z>�C?��>�D<>��>Jϴ��1��L�h�'w�B̽� �?>����J��1��9��ޥ��{j�=%b.?S}>����>пr���B2H?t����)��+�:�>��0?qcW?͛>:��c�T��6>_���j�ra>�) ��}l�Z�)�1&Q>l?��f>!u>P�3��c8���P�z���d|>�-6?_.>9�&�u�ݫH�gWݾ�VM>�ľ>|@C��j�,�����ui�q{=x:?�?�V���ాb�u��B��\7R>�.\>أ=�v�=0[M>�9c���ƽ�H��.=f��=�^>{?:+>9Od=@��>\���{�U��>�>n�L>�q&>�[=?T%?�W�����N�}���$�,�>K��>��>> \M��Y�=�9�>�ma>������Pq�#]4���Q>�쐽�[\�)�u�^;X=o+�����=�S�=�����<�A?O=�~?���.䈿��#d���lD?J+?���=F�F<��"�; ��pH��@�?n�@
m�?��	�ܢV�6�?�@�? ����=}�>$׫>�ξ�L���?��Ž[Ǣ�ɔ	��(#�dS�?��?�/�Pʋ�Bl��6>�^%?�ӾPh�>gx��Z�������u�"�#=?��>�8H?�V��-�O�s>��v
?�?�^�⩤���ȿ6|v����>W�?���?_�m��A���@����>:��?�gY?`oi>�g۾'`Z����>ѻ@?�R?�>�9��'��?�޶?կ�?�Ha>���?��^?ܦt>œ��>��u��������=	Vm>�y>,iT���� aY�3��zk��k������>�}=,��>򻅽3�ξں>�w�vw�JHɽz�>U��>Ɛ�>!��>h$?��?/-�>�_E=����K�"���S?���?S<S�6�i�<[�>g�9=OǤ�LΣ>�g?8�><�h�f$�>:OZ?�s?A}E?��>�� �s����¿���<#��=�E�>9�>�<w=%�>���N7a�˸�>J_>dR6<�Փ�I�
�Q�<�s> �?ƀ�>���=Qd?�i?w�T>ђ >�(R�&�q�d���>��n>ʓP?~fl?'9�>����GQ��7��ؠ�>�Q�T�>>�.l?H?n]�>u����ʧ��h>��=9��K??�Ux?�^��e?�}�?��Z?�{?.D�>h��=A'��N�=�N=;#!?�w�}�B��<'�Q��"^?��?=4�>�i���н��¼���}��+�?*[?	�'?�L�x(^�uq��y��<eh���摻�7�;��E�Sj>�~>��m�Y�=)>��= �g�_7��<<�l�=YP�>u�=��3�Uօ�=,? �G�"܃�=�=/�r�(xD���>LL>^����^?�k=���{�w���x��xU��?��?4k�?�����h��#=?��?�?6"�>�J���}޾��ྐྵQw��~x�=w���>��>�l�A�0���Й��_F��I�ŽW� ��>/��>��?-2 ?4^Q>���>�9��'�;&����^�<��._8�F�.���]/���O"���	�C�����{��ʘ>b��x[�>Ԗ
?n�h>%6|>>��>3���� �>a�Q>�H> Ǧ>�V>�D5>>��,<W�ͽLR?3����'���辭����.B?apd?A'�>F�i�ۇ�����?���? s�?Bv>�yh��(+�fk?�.�>�� m
?`�:=y*�%l�<BW������'���C����>~׽�:�,M��kf�Dg
?�(?�ӌ�A�̾;+׽8�\��;_Fo?�L$?d��ni��2t����?�t���>�H�F����A� P���ס��h��������Jd>�??x��?yW��8�����e����x��>6~?�)�>Ly9>�\>'�+�I���t���)������?�Q[?�V�> �:?|� ?]|?9'A?��>�q�>�`��A�>�횽�G�>7o�>�d??d�6?7[#?��?W�:?�� ���[��/���ء�y�.?��?���>�v?�> 4�ޯ2>O%�~�%���+�ˏ����"=֬�=Ľ�uj���>�f/�>�L?����8�C�����j>�X7?��>�H�>���i�����<z��>��
?�+�>	����)r�:&�h\�>���?NU��� =ܩ)>Ų�=���Hʺ4��=#X��^��=�e��f9;�8"<%P�=]��=~Ig�������:��;Ip�<uL�>�@?�>�X�>����iS�N�� $�=��[>�Y>`>I۾(����W��ai�3w>ji�?۠�?��x=���=:��=О��P�¾�_�;;��fd�<�h?6L$?{T?��?֜=?�1#?>=��ޒ�8T��H�����?F,?��>����ʾU騿C�3���?rQ?	Ba���.)��¾�սW�>�Z/� 9~����7D��7��{��Ƨ����?¿�?�=A���6��C�'����u����C?�=�>�J�>S�>Я)���g�1(�aM;>�n�>��Q?��>��O?��z?��[?��T>;P8������♿�2�>X >J�??���?5��?�y?���>R5>�(�ϲ߾�����}��6���P=
jX>Ò>ζ�>��>�H�=4�ʽ컰�w�=��=�Ub>Do�>�G�>s��>.y>�{�<�|:?,�>�t߾(���a��Z:�����='�r?5��?�5*?gJb=��o�$��$þ���>b�?���?�&?����a�=��9���˾zY��J��>"Ɩ>Y��>�,�>�=��@>�
�>+ύ>������:���5�,���ϙ�>}�?G̈>,w�������>NqD�M��zz>ݕ���U�>�=b���<�"����y���'���ǋ�n������c醽%+ݾ���>�t� Jl=Q`<>�#@>Ba=�i�=�	F>;w;O`�=^z����)�K�v�����<�X��(�=���<8T>W�e>V�˾Ύ}?:I?G�+?�C?,�y>"H>��3�à�>�����=?\*V>TlP����@v;�-���h����ؾ�t׾(�c�Fǟ�SD>�vI���>�;3>-C�=�l�<�=�s=�Ǝ=�qQ��=l!�=O�=�a�=��=��>�P>�6w?X�������4Q��Z罤�:?�8�>p{�=��ƾq@?��>>�2������yb��-?���?�T�?>�?:ti��d�>O���㎽�q�=J����=2>o��=r�2�R��>��J>���K��F����4�?��@��??�ዿϢϿ8a/>^�8>[>79S�$�1��Y���b��lY��}!?�	;�6�˾���>曼=޾�fž�V2=��8>.�c=����[�D�=�R��`�<= �p=R׈>R�C>���=�_���+�=7�C=,��=�P>�銻x?4��*���+=TL�=�c>�&>zU�>�"?��?��6?�M�>n|��%G����ԇP>��A=� �>��>؅�>��>�A?�`?���?{��>vP�=�4�>Bq�>�o%�5�t�Cݾ����d=���?#
�?_/�>V&��}�߾�/�<-��̄�l?#?��;?��>��>|��l]�B�%��9���@��;E�=V�齇�N����z[������ '�=G˘>���>¯�>�k>�|>��X>�A�>��>-<�=$�j=����s9�=ֽsSH>� =��=b
�9I�=_x=&s��E�����O;�F
;fkD����I��=��>@<>���>}��=���C/>������L����=�G��Y,B��4d��I~�Q/�"W6���B>P:X>z|��%4����?��Y>�l?>���?#Au?E�>a!���վQ��UCe��US��˸=��>��<��z;��Z`�_�M�.|Ҿ�f�>0�>w��>	5i>B�+���@��M=Ļྐྵ6��>�����7�����r�� ������
g���n�$D?L��0��=(4}?�I?:�?Ğ�>����u�޾�n>6Ol��MN=���i��Op���?$?��>����D��Ⱦ�z���ݶ>g�F��R�ј����2��F��C����>[��Ph־b5�d}���J����A�@�w��ݽ>WP?�]�?��K�vŀ���R�Ѓ�-�����>Q>d?�Y�>$�?��?S���<�I7���y�=��k?��? �?N>:�=�%��<u�>��?i �?�ِ?:bs?s�@�}L�>w/(;޻">0쎽�d�=S>�|�=>�=m�?=�
?^�
?���a	�������`�_�<x7�=rp�>�Ň>�Ao>c�=n�g=�#�=��Y>���>�>��e>���>�>�ڧ����T�(?��=��>eV3?T��>��p=]��3��<�9d�89D�5z/������Ln�<���Z=%V���>?�ƿ�V�?0U>� ���?'*�ï��RR>��T>�ང��>��D>�x>7�>b?�>Vv>u��>��+>�FӾ�}>9���d!��,C�ςR��Ѿ�~z>����	&�'���z���CI��n���g�Uj�S.���;=��ƽ<H�?������k���)�����Q�?�[�>�6?ڌ��
��0�>���>�Ǎ>�J��h���ȍ�rgᾣ�?��?�Hc>w�>y�W?�?�)2��3���Z�r�u�,A��d���`��捿����ն
�$w����_?��x?�}A?�*�<�'z>ɯ�?��%�)��U�>y/�4E;���;=��>����EPa���Ӿʺþ~R�\F>J{o?(�?dk?*]V�=��=�H�>2�>]�^?'�D?�0/?�T?���"C?ӻ�1 �>nzS?�39?�>L?T�>?Ȅ�V��>���@�q=P�0���R�����<<�IV�;��k������>m/����*>�>RqX��o:��-Q;Ь=V=�ӭ=7��=v�~<c�>J]?+��>���>�7?4��9�6�/���Z`/?�*B=Oف�9�������>��3�>��k?��?�	Z?��g>��A���F�i>��>8�&>��Z>xǰ>݇�D�E�zo�=B>�F>���='ba�r,��f�	������1�</�">���>J|>�i��S1(>$	���bz�2ne>��Q��k��.�S��xG� �1�*qu����>t�K?��?Cc�=`� ����Cf�~ )?�<?=�M?�f?h��=�ھ]�9���J������>Y�<�����������:��&;��r>➾�ꟾ��c>!M�*�ݾ��m��I��o�c�E=vh��Z=x����Ծ��~��"�=*�
>/����#!�ꖿн��D�I?�l=�Q����T��K��̀>�ח>6��>��5�'x�>8@��p��#��=�h�>�!<>��������F�P�w\�>;�C?G�R?�e?����z5K��I�/J���;�3�='��>D}e>��!? !½�=��)���+��Zb���~�7~�>�_�>#�O�|P�p>���g�W����>Ic?c�o�~7?'�>��?!?��?7*?]�>h���Dy���%?m�?�K��χ�꽤���6�Mm�:R�>�)?���Mr�>�Q�>�!?:?�eP?�4?��<�{"���Q�e8�>	�>&k��󦿎Z?��M?d>��?�·?�=L>�EM��go�����5G�>�k�>�(�>��?We�>���>�A�>d���s�ǽ�>دm?ʆ�?��`?k�>��>g�>�4?x��>AW7?���>h?3d?>[�?R�o?�C?a
D=����k%��N(�?�]=1�E=�8.����=�5��PA���=7�/>Ȫ�=r�<�^y���
�$�=�l-;"�����> os>�f����3>Sa���Ȉ��8;>�Ѯ��ל�쉾[6��P�=´x>Zo?�@�>x�'�v4�=m��>D��>���4'?��?yw?�#��Cb�Tؾ�1K�]Q�>�{A?/�=�l�Ó��v�p�\=�4m?�o]?l�T��c����b?z�]?d�&=�w�þB�b����B�O?|�
?A�G����>y�~?�q?���>� f�8n�;��Bb�>k��ƶ=H~�>QW�G�d��W�>��7?jB�>��b>&��=ug۾v�w����D?���?��?���?9+*>�n�-��\��N���r�\?��>����� ?����:�ɾ�����ʉ��5�┣��~��~�����2p+��&���Ľ�d�=х?��v?9�o?3�a?9���e���^�4‿%U����k�3|E���B��oE�z�p�^<�m���:����="ǁ�R�5��w�?�?+q4�W��>��Z�6�̾*��5�>1ξ��=(�=�]<���=�Eռ�꽾@���lX���� ?�G�>+�>#H?L<g�;4�+�#��8��?�?Q>�R�>qb�>��>e����)�r��l�þ>���g�t��T|>k�]?�yQ?��q?����f�0u�!V-�V<�2¾pP>���=#�[>�yE����=))�$�@�~�j�@	�j͍�5�ެ�==�+?.%q>�c�>���?pC?w���,ŧ���*����g��>��m?��>a>����`�	!�>�mc?:��>��>�	������t�����]�>q}�>�D�>�X->�p=�jV��l������!u6�=�=��c?�#���fF����>��P?}-���a=��>v ����?��6xA��1=Q�?1��=t�">�=�����t�j���T���.?�$?ܦ��1~ ����>"�%?�v�>=�x>�z?���>�}Ѿ�BT<	��>o�r?�7O?��?.�>�@�������b����A���<�6�><Y>���=;��=�;�̡n���0���=�>b����K��+��k��>�=��=c=>vPѿ�qQ�ėȾ�����
g�¦f��}�����1k��nF̾�'E���x�h��~�3� {���<����<��LA�Fb�?��?9���ڴ�6���ш���� �o>vͅ��f;�gE��53�����V���辛��eYK��p���oq�s�'?X�����ǿ>����3ܾ:! ?�> ?�y?��4�"�x�8�ʬ >�.�<-͜�
�뾔�����οL�����^?���>y��3�����>���>A�X>�Kq>:���鞾3�<;�?Ї-?˝�>��r�[�ɿ>���ܤ<���?��@E?�\!������N�=Jk�>ǡ?G)>��4�Ӽ�j��-��>%t�?_?���=��L����Y�]?��l��yE���n��=���=BD�=��,�+ &>
c�>'c��V��ڽ�
G>Т�>b5w���/��q��f
=r3[>R���*��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�I���Mɿ�|�@���S�����k�4>�R(>ÿ���]��0Ⱦ�K�vz��>��UR�4�|>@s�>jl�>o�>~Q?H 4?g��>�>�8'=���湹��!->勾N8O��Ͼ1`G��ӾiU ��BQ�/1�m;���ȾT�þ�E�fpX<�$P�9>����L$c���7�q8?4 >�̾�U����.UҾ������a�%�ڽ�����!���_���?:(3?z>}���W������Y�<����Z?�T��� ��>þj�>�Aj��v�=}��>x�=���z7+���M���H?i)?���ZJƽכ�>��X0��8?cp�>�^���>E�D?�t�z��=	B>hR_��r�>�ڒ>|��H���eｮ)8?�Y?�^����þ���>�`����Ͼ��>�|>s����.�������b�+�7t�=��=H���V?ؗ�>��)����䓏��-��F=̵x?f�?��>�Ok?DfB?'+�<������S�{\
�8�=�W?4di?J�>> ����о?���y5?��e?Q`P>� g����R�.�?T�7�?9o?R�?�,��v;}�=������6?��v?s^�is�������V��=�>2\�>-��>��9��k�>"�>? #�tG���bY4�*Þ?��@t��?:�;<\ �^��=i;?\�>��O��>ƾ�|��z���o�q=�"�>����Bev����6Q,�n�8?à�?���>蓂�թ�i"�=�����?�_?�Vھ&o.��%��uC�� /�fu�=Cm�=B�}=UA���z��J�H<���o��7�ͽц�>�h@��
��I�>ї�����b{ܿ�ɒ�㈶�#'���4@?�MH>�����[վP�s��V�o�A��h���r�<+�>L�>+Δ�)��Z�{�dq;��-��@�>+��
��>J�S��2��͈��Y3<�̒>���>V��>�9��v�U��?�S���5ο�����x���X?T�?]i�?�X?�9<Hw��x{��$��9G?��s?:�Y?��%��6]��37�(�j?�_��qU`�׎4�cHE��U>�"3?�B�>^�-�ֲ|=>���>�f>�#/�q�Ŀ�ٶ����O��?Ӊ�?�o���>x��?xs+?�i�8��z[����*���+��<A?�2>)���1�!�K0=�VҒ���
?P~0?T{�F.���_?�ba��p���-�h�Ľ)ա>ϔ1�ty\��d�]��[e����(.y���?RV�?���?h���%#�W%?i߯>����QǾ��<d��>sc�>�bN>�za�ţu>���A�:�M�	>��?l{�?�Z?S����ݦ�N>;�}?�>�?��=�B�>xu�=�ʭ�C�IZ>l\�=����?��N?��>Ou�=~�6���.�^�F���P�� 	��tA���>�yc?��L?2�T>S�����$�ED!�~bս7�*��"���7�_!)����1�5>�7>ƃ>��F�QԾ/�?�z���ؿo����'��4?�у>(?q����t����#_?q�>AF��2��a�� �����?w>�?��?s�׾1:̼'>1��>�-�>#lԽ�ԟ�����8>ܑB?K�*A��@�o�R��>���?��@{ˮ?$i�	?8%��R��!g~�����17�y �=0�7?�0�=�z>���>��=�hv�������s�v��>"C�?�z�?8��>פl?~o�z�B�P�1=t6�>�k?�w?h�m�&�D�B>�?��.����F�pf?M�
@�r@&�^?w��Կ嫖������Ǧ���;���s>�9��XVU<٩?�\�=A�[�\ >�>O�V=��k>�ژ>,��>�G�>�����G���䂝��p���3��h޾v������u��6
������ξnK���������|���PG���>1a?:r;?�D?T�>��=�-W=�Y�)�>��C�M��=�)�=/�?�J?�q#?��z=a����#O��s�����wh�i��>��a>|�>��>ͽ�>��<�O�>x��>�#a>�"G>]ѩ>?�K�W�i=fZ�>��>V�>GN�>#l=>&�>�ô�H����ig�/zv�0�ҽ���?/���t9J�p��?����M��
��=��.?��>-摿�Dп�ʭ���G?E����I��4+�f	>�	1?5W?�>u[��N�P��>i����l�·>}���Oyo���(�C�O>v�?[�h>ePu>��3���7�SO��ȯ��~x>��5?nD��g+9�hRu�V�G��޾�jP>�6�>t�k�-+�
薿	�~�!�h�?5v=!3:?�?융��6��A~s�*~���PP>r�Z>��=��=��J>�e���ɽ�mG��l.=���=��\>�~?Q�*>�O�=W�>�c��@W�-:�>n�>PO�=8C?_-?k�N=���{�;�=+>$B�>t	G>c��=J��e}�=[�?ǳ�>~蹽�j5� �ǽ��愕>�c��@��	�Y�
>3'��?�=ne�=X�@��煾d(>�~?�x���刿���鵽`mD?!?�ΐ=�G<�{"�%���4?��7��?�@bl�?a�	�T�V�<�?=�?U������=�r�>E߫>xξ�L�J�?X ƽ�ɢ���	�v#��Q�?U�?��/� ɋ�Rl�m9>I`%?��Ӿ<O�>���MX������u�j#=���>3?H?�V����O��0>�q
?�?Y򾧨��9�ȿ�uv����>��?e��?��m��;���@����>��?�`Y?��i>��۾�[Z��u�>n�@?��Q?�.�>)-�E�'���?<۶?+��?}�3>#O�?��\?�2�>A�����E�2۲�1҄�^�������b�>t)>�$Ǿ�<�qN������'r�����=:�=X��>������e>m�=	���L3E����>H�B>M>�i;>{��>�X�>	��>���=f���|9J�����/M?��?��"��`���>>�3�=����A�>�z1?���<L�辊��>\D?���?��g?
oM>���ҡ�C����瘾
�HS�=[}�>���>!�=Մq>�%�1�W�>��V>F�=�6��S�Ž��T�ܿ>�c?L(�>��7>ؙ ?��#?��j>�(�><aE��9��^�E����>���>�H?�~?��?xԹ��Z3�����桿��[�;N>��x?V?�ʕ>`���생�MgE�BI�����N��?�tg?T�%?,2�?؉??\�A?�)f>��ؾ������>Cz(?����nTN�4��J��<�?�>~��>b5�©��=������Ƭ��=7(?��`?�| ?����ào������:=�M��༭^�=��-;�$>�4>����>Z=G�=_"�=���i��Y=m#=o)R>��=���F�<��A,??&G�`̓����=�r�ppD�`�>pL>:����^?W=�{�{�D���o���U�>�?���?�[�?���i�h�==?d&�??���>%6���c޾����v�]�x����r7>"��>�p����ꃤ�՚��I���Ľ��V=�c�>��-?x9W?EBY>�?���>����z��>�e��T#�4v�$�2��@��žE/�����o�ȭ2=�h��(�ǽ�j\>}���f>Pw?¬>�W>�d�>U�!�O��<�!	>BJ�=n�>�S�>|�q>k �=yd=�����R?���� )�'���A����A?a?n��>�qc��䄿�'���?��?̜?��x>
i�JR*��N?Y��>��}�[�?m3@=�#D�@�G<¹����
�u��s�@�>�VнJ�8�"�M�ʗi�u�?�(?{V��~Sƾ��.J���Hr=�?�s(?z*��eR�h�o��5W���S��I�F�f�o����$�ԃp����A\��J!��"�(�J� =�f*?�r�?)w����g���@/k���?��{b>!�>@b�>9 �>19G>Y�	�$�1���]�u�&�X ���>��y?�x>SdJ?3?��=?�BE?�$�>U]�>������>r��=[��>��>H=?a�&?��#?�Q?|
?�3>z��CB��a���� ?��7?���>���>�+?*l��V�ʶ=�]��U��. н��; )��������C�=�o>��?&���C����>R�9?�շ>懪>}8����j��D�;B�>K�>��>2�޾:�x����[.�>�Ay?����g8~�>�>c�Լ8��UU�=ԅ.8�#a=UEi�j̻y�,=�X+=J8d=�y�M�U��
���={�=n�>��?�>�=�>d���� �Q����=�_Y>=0S>K>vZپ�u���!���g�r�y>:{�?9v�?�h=���=R[�=�Ġ��|�����	�����<ڥ?�#?O9T?�~�?��=?�t#?�X>�I��F��AV��`ڢ���?~:,?�k�>����ʾ���}3�nR?�4?�Da������(�������׽�+>�E/�!'~��֯��C��1��A��#"��̜�?��?�9E��6���˳��+���S�C?g)�>�3�>3�>g�)�-�g�:��;>�/�>2R?h&�>W�Q?�Lw?3[V?!X>�6��w���g��Ӛ��21(>�y??~?�t�?lw?�{�>vt>Qe6�>w߾uT �#%�#�����1lU=
ha>���>"j�>-�>���=���MS���ED�o�=�Fh>���>��>���>��w>�G	=@@?:��>pύ�����BD��͵r�r	=�r?)��?�>)?���=�j�W(?��� ����>�j�?gc�?(.?_}�֦=1 ѽ��޾d����B�>f1�>z�>%-�=!ϼ��=��>��>�ֽ���]O�n���?��E?d�'>��տЖ���Ѿ1�󾲩�����2Ĩ;�ğ=U���3}9=bQO��{�wu��?ؾZ���5�9����8���]��&�>��<qC,>��)>���� B����=+=�;�EA=k�=�Rm�� f���뼵�*�jh/�=�=95Z<�P;`�N���ľ85{?�YK?,�.?�??�}�>N�>Uo��>~N���?��D>�L`��|����A�ҭ�߹���ؾ�оo'e��@��`>C�T�.	>C>���=�<'��=̔J=5%Z=�M���,�<4P�=�y�=2�=�F�=��>2
>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�??ti��d�>M���㎽�q�=K����=2>q��=w�2�T��>��J>���K��B����4�?��@��??�ዿТϿ6a/>/BL>�
>I�U�U{+�(I0���[�kw�[#?E�6�&�ɾ�7�>��=��^֮��^=U�>%WC=�"'���[��=#���+^c=���=�|>X1>/��=�Ȝ�}�=�(2=�J�=�GV>.ܜ�0�_�9?`�`|V=ˋ�=�2|>��>���>��+?!�U?ǶW?5��=���eqɽ�n����?���>�ϩ>��=9Y>�v>�d?"no?%�#?���>s�>�4j>8{�>���m\�����&n��^�Y=2��?��H?���>`�S>�����8�4��d���c4?A�T?6s ?"��>�N�`��&���.�$����=y�{kZ=wl���\�˸μ'����b��=�>�>���>��>��>%@>H�_>p%�>�>��=���=1��:���<\˻��<{=1Ƴ��~�<~ϼ�o;��·z2:���v�KM<��c���J<e"<�q>�H�>J�&>D��>疗=�j����>������H��/�=`���?��b���y��q,���H��=>��7>Z{d�f���DN?ܸ�> Y>ܝ�?s�q?T
&>s�-��殾�����#}��d�����=�:�=�p;�w�5��j�[�L��P����>��>
¦>`L�>�:$�#I<�v>=#J�Um3�@C�>B�}���!���+�.k�����?����^�L��n�=?�Ǉ�)��=�o�?M?[1�?<�>�}�h����>�q��h�
�&�hA�g���o?�0"?�i�>��ɂ.�eҾ�ͽ�>k�R���Q��>��3.���v��;�����>t���e�Ѿ92��Ն�kԐ��jA�L�h�X�>��O?��?Ŝd�����|uN�XZ�bQ���:?O�f?S��>aN?�U?]*��P4��:�r�=Ќl?��?�5�?�>�V>����Y�>C��>-��?���?މ�?�b�<��>�E=]�>>�=�H(I>O�Q�<B����>�!)?nP ?ӽ<?���Zx7�*����z?�Ӛ=n�F=D�>�ʢ=�> ?>\��=	,�>��n>-�>��>Eh>wN�>3��>	�վ�-�[?��l��>��?F%�>s>�b����V��(�Ž(�n���O<(���'�3�lF\��	>7� =��
?�����9�?�:E>�C꾙$"?�i־�ɼ>A���\>ϣ?���?nz&>v~�>���>�"v>%���ӯ>�>MQӾ�`>n���h!��)C�ÂR�ճѾ��z>����&�%��]���qPI�fj���h�Ej�K+���4=�g�<wH�?���a�k���)�������?�W�>O6?(��������>��>���>,1��T���Mȍ��u���?���?[c>�$�>`�W?t�?C�1��R2��RZ���u�"�@��%e���`����p���x
��d��p�_?q�x?�WA?��<pz>q��?9�%��ߏ�y�>�/�H;�K<=�*�>���`�`���Ӿroþ��L/F>��o?�&�?�A?nNV���m��('>��:?��1?It?��1?7�;?����$?�m3>!@?go?	I5?v�.?��
?:�1>���=�*��г'=Q1��늾�~ѽ�kʽ�w�F�3=�{{=�
�,�
<��=���<[��Xټg�;ۡ�F�<�&:=M�=1��=��>c]]?a �>�ƈ>�2?�� ���-�7���T4?��z=�a�X^���o��:'�A�>Qq?�0�?6WY?�tt>F�E��RQ����=��y>?>;Ak>�?�>Qk��)�H�p@=�>���=�\�=T���v����Q��{�"}-=2~/>���>�0|>�č�wl(>]��z���c>�PR�����u�S�P�G�ս1���v�U�>
�K?k�?���=B}�2T���+f���(?�~<?zeM?�j?�ݓ=W_۾6�9�j�J�������>\�<Q�����'	���:�w!�8�s>��\����Yf>��
�ǖݾ��l�)K������/=���ʗc=u��s�Ѿ�|�P��=�>����o:!�B���K���`I?�h=�M��ES��[��a>���>�s�>R�-���m�P�A�x���|�=F��>�?>)���N���G������>�D?[�??Ii?�q��Kف�bl�����ﾗQV=H�?���>Y�?:�=��=��V.���[�{�N�&.�>BF?w6�lVc��޽�E߾ױ2�}�B>�+?H>56�>��=?({�>�*W?�?jS?��>\W�U�޾ۈ'?�B�?6�2�0r[�{|'�<���Xo��U�>5?~(=��q>���>/�C?��?�x/?�?J�>�����U����>���>��^�9Ƽ���A>5�E?��>�;?�q�?wB%>g���|��=v]��bO>*��>��C?�3X?�A?жW>7��>lRž�Y_��M�=��m?qJn?`M?���>��>��>��>e���x/�>�
4>t�?��|?��o?��w?`�"?a��ȴ����y6����Ԃq==4�=�	>�a�=�|^�K����ƽ"2�;��:Ч:=m��F��m����<;��>-��>G���4S>(���!���zW>�̼j��ύ���x����=1Ce>??�@�>U�8���=�>���>(���?^�?T?�ѽ�Mb��ాBkR�l_�>r@?�o�=U�t�A���o��57=94c?�[?��2�Qg�^_?ʤ^?��v	;�����ݩx��{�4ZD?q� ?-�'�x.�>|�y?ӟs?���>P�{���j�t��Pqb�Ȗ�����=Q)�>S}���j��ʧ>�Z7?���>9IZ>S�!>�ξq�t��q����?�?�?��?�:�?�^>7*m��f޿��������d]?b&�>8���&�!?ٺ��;j���؎�Wd߾u���m*���И�k���?&��R���Eؽ#��=b]?�s?A
q?�>_?�L��R�`��K\���}�V�'��Q���E�DF�� D�&lm����l������#KR=�sx�W(����?��*?�tk�Ȍ?�{��ӻ��l!�:�> ���'ɇ��5i�;���p�ؽS�Ѿ!7侣�>�a'?�f>6��>A�%?�3h�����9��3���$��?�>��n>M>�U?�ɼoꭽcBL������;���A�R>2�b?�P/?{`8?Z�G=ߊ9��a��Uj8�Z�]�g��쉱�LA�>��>��4�Wf����).�$̘��V,�����Y%���>��[?�F�=�j�>��?���>Y/	�$߼��Ǿr��n=���>|�M?���>O|3>�F�#�d����>�Sl?n�>�{�>�B���� ��z��@Խۿ�>z �>���>��n>ȷ*���Y��;��e���t8����=\7g?~����^`�!a�>kwQ?���)�<���>3���r �����u.�Q�>b"?�=�=��;>�Jƾ�O���z�����-?�S8?ݧ��b����>kA?��>"�>�oZ?�>������ԓ�>KA?|�R?Jf+?�o�>|%�=��M���e��F��ϼ��>f��>�t�=-Z>V�\{�B$��7Z	<o�z>�"�� ��;�+��!jӽO&�N͂=܅S>bVۿ��K�зؾ�������
�V$��K���݅��}��b�������x���ڕ;�~�U��ba��挾)n��*�?��?K��fԈ�l晿?��g"�����>m/q�ά������_��ߏ�����%����!���O���g��d�D�'?����ͽǿְ���:ܾ6! ?�A ?�y?���"�ʒ8��� >�D�<�*����뾰����ο������^?���>���/��c��>֥�>6�X>4Hq>����螾k.�<��?1�-?H��>�r��ɿe���H��<���?&�@�`H?�K��D%)����Y?�?�a=�wH�(&�0|Ծ@�>�q�?7�?�>^G=����cH?�R��Q��"<�����=BV�>�q����`Չ>#����4����m��K>N��>��A=�\�=U���������<>���f��H�?e>Z�bxe��&0�S��A�>�U?=��>n�=�%?ĭB�/�ϿZ&Z�`?C��?{��?��-?�%��&��>�aվX]H?[7?;;�>B�+���r��w�=���TyJ<�˾��L�//�=}�>n�%>���w	���&�Q��;̄�=CD��?���x*
�*��H��|�a��xԽ�н���=kO_��~?��Ǥ��t=#Y½��(�+D>��Q>� =,�=H�O?.|r?g��>��>�7�=`�+�I:��v =���N�0�s����4��޿���C����ȷ޾1�����վX�<�GЎ=�R��u��� �D�b�r�F��.?C�#>Bʾ�}M��*<n�ɾ|�������<��`̾ۀ1��n����?/2B??����.W�"�����F`����W?lQ�n��2����!�=�S���h=��>���=`����2���S��5?>�?羑d^�/ړ>�(�P	{=ݮ?�+�>��#�^ʷ>�
)?��4st=��>��>���>|��>�=k.��^���,?x�d?r-���Wľء�>{���q`�n��=�>�����%���I>�^;�c��k<�#�d�0=�|S?�x�>X�"�l��80�F0�� o'>&�n?K��>�6�>�q?��?T�u5���$���ھ>H>�zV?
�i?�u�=� ���^ پ�&U?w�d?Ӵ6>� )��h���d8�e����)?Y%e?j�>z���w��㓿�+��(�*?r-r?�[�"������&"�酣>v`�>�4 ?q~2����>�:?��8�N��������C1�cޡ?�T@�R�?S�G=��:�B�=Jy ?���>�8;�Q<ľ:�����ҾD�.=���>�#��[k�_s�P���6?��?�?����}�����=7������?�s?����3���1�GwD��,���>��W=�����*�'�E��̾�(��b���>���>]~@V���#��>�bI�B<���˿_���	A��t�i�L?�d�>�\=�_�9�y�W�u���<��1�������>oc>�x>�E~�2y���<��!Y�`��>'�żb��>\����̾&0���A�<p�>��>��>5ġ�|g��ύ�?Ξ�Kο�'��&����U?"5�?���?�9?�Z�<e�g����P�]���L?��m?�I?ЏW��S:���a��j?�_���U`���4�2HE��U>�"3?=C�>5�-���|=�>-��>�g>�#/�e�Ŀ\ٶ�����e��?܉�?�o꾾��>^��?ps+?~i�8���[����*���+��<A?�2>܌���!�$0=�BҒ��
?V~0?�z�m.�W�_? �a�S�p���-���ƽ�ۡ>��0��e\�0M�����gXe����@y����?A^�?_�?w��� #�k6%?�>m����8Ǿ��<���>�(�>�)N>�G_���u>����:��i	>���?�~�?=j?핏������U>��}?�J�>���?&Q�=G��>�M�= ڱ�s��v�>��=7�U�p?tsL?�	�>���=c�9�V/�)�D�J�P����/�B�;��>ʦb?�L?�[>C���m�%�z5!��'���0��o�ϪA��V1��m��/6>7�;>	V>�,G��Ͼ��?Dp�2�ؿ�i��<o'��54?`��>D�?����t�����;_?�z�>�6��+���%��	B�n��?�G�?�?Ļ׾RS̼$>E�>�I�> ս����V�����7>�B?��fD��H�o�[�>���?��@�ծ?hi�Z	?���Q��ua~��w���6�h��=��7?�&��z>��>��=zbv�ʹ���s��ɶ>�@�?b|�?���>��l?��o��B�32=O�>��k?�i?6Cz�� �ψB>�?ƫ�6�HH��f?I�
@�r@��^?�좿tֿ������ξ�X����<h�=un�>	������==2�������<82=���>��>хE>�PF>	su>F�>0N��q%�Y���w��8mF�t��ԾȾ�� �پ�߸��m���־-w�ϗQ��/���	��精P}��ʋl<�/u>��A?��r?ދ�?��p>���=�EL>A�/�7'�>��P2U��0�>�Kv>��B?�aC?����ʾ;/5�T�U����<�-����>Z8>�#�>�}�>5>�m���L>��>:u�>��=>f&����yߋ>�N�>Gn�>.q�>�ƚ>�C<>��>Fϴ��1��i�h��
w�|̽0�?���Q�J��1���9��Ҧ���h�=Gb.?|>���?пf����2H?$���y)���+���>}�0?�cW?�> ��x�T�3:>8����j�6`>�+ �~l���)��%Q>wl?a�f>�"u>��3�2^8��P��|��Ic|>�*6?�춾�79���u�
�H��[ݾ{PM>4��>ަD��k�G�����;si�
S{=`z:?�?-S��Tװ�|�u��C��)?R>�D\>p1=�g�=OM>!c�v�ƽ�H��4.=x��=��^>�7?��R>H_�=4l�>H鍾�y��T�>���=��%>�U?�g?O�������Ĝ���b���>���>�-�>J�K=�{����=��?��>R~ٽ�C�<�t�u���W��>�f\��ɸ����=��bn�=�͖<����}~�*�=�~?Z��4䈿%�`���lD?+?S��=��F<��"� ���G���?`�@�l�?��	���V�$�?�@�?�
����=�|�>�׫>%ξ<�L���?��ŽEǢ��	��)#�S�?��?��/�Xʋ�Kl��6>�^%?��Ӿ0h�>�x�{Z�������u��#=R��>�8H?�V����O�U>��v
?�?�^�੤���ȿ2|v����>P�?���?V�m��A���@����>=��?�gY?�oi>�g۾X`Z����>û@?�R?��>�9���'�p�?�޶?կ�?��F>_3�?�jU?��>�޼5O�%Z��o猿ci�<֤�OZ�>�1I>5���ȸ?��U��`���i��*��?s=]�<��>�н�Ⱦ�rf>�H-=������:�>J�y>�c0<�f�>4��> s�>�>�	�=����߿��cj��=K?�;�?��akt���
=:u�=���.��>�'1?�q4=ǿ��;��>}o_?�hz?��V?�;�>`����R��{���U��G!P=�V7>���>�C�>/2���>�(ѾN�>��<|>zQ�>M�̼�1��4d�)m=?��>��!?���>�+>�?Rg"?t�l>���>�F@��Y��~�K����>�A�>�:?Mmt?�?�6���W3�1����ޡ�Jmc���@>��v?��?�=�>/�횠����:�_��X�&S�?r_n?��½�R?�d�?,K;?�:?�Q>`���w����`���G>L�?#�� F��3*����#?{ ?�;�>O�9����ρ��-�1U��~
?�xa?�h.?��ھs�M��L����<v��A|�<�Qͻ|��>/U>�3%��Q�=I'>�6�=DJb��yY�VV�=E?3>x}�>I�>slI�����1=,?��G�3ۃ�h�=c�r�@xD�V�>IL>���R�^?�k=���{����mx���	U�� �?��?8k�?���*�h��$=?&�?Q	? "�>FJ���}޾���Ow�ox��w���>���>+�l���5��������F����ŽN(𽻶�>b�>.�$?j��>�$�>e�>5���>оy�,�IK ��>� ���B���1���;��8Ͼ�-�d3��ؔ�nKA�Ҩ�>!�Q�Q�>�$?��e>���>�w}>=���|}=��B>�>'M>=��>2g=�!�;+]=q�3�o�R?*溾��(�)��1|����??��a?��>1�z�s�������!?�f�?aB�?�Cm>�Nh�Ň)��?�)�>��ؐ?2jb=�<n|C�m$���~������$�<^�>����;�a�M�^^�X�?�?O����ľ�νI u���=�Ax?Hc*?֣)���H���w��[� ����=	�z��j�+��-�]�~Ĉ�� ��\X���V4���;��'?��?��.����m��Gf��Gc��T(>�d�>��;>F��>/�>�Φ�7�'��R��������?�=?�-�>dF?��@?�	Z?��8?��>�k�>����4?�{����o>��>��)?yZ+?�j&?��?S�$?ɰR>ר�����[;�|?�?�0?|b?��>�U����q�|7��fk��^�;"#��2�<�9�<�*��iٽ����o@>�Q?W��:�6��;��N�g>��6?���>���>{y��NŅ�9|�<:��>��	?��>dR����r�U��E9�>́?q��� =�*>��=�3��Aʅ9���=�g����=�b��/R6���7<p"�=y˘=���:o�-������-�;�Q�<��>�?���>�O�>ޤ���V�G��M��=��\>�
V>@!>*uھ~6��N���SMg���>��?�ճ?�ta=���=��=j졾�_������&����=��?�� ?��T?:��?&;?��"?�~>h������􃿟����?+,?3��>���Iʾdר�.v3��?�?�Za����S)��¾?rԽ
%>�O/�� ~����� DD��������4��e��?V��?}�C�;�6�(����Cv��9uC?���>~J�>4�>a�)���g��<���:>Ǝ�>�R?��>ۈM?��}?lz^?`�8>�T/��̧�F|���<��>�.?ρ?���?Uu?��>���=T�0��O�u����`3�U�y���e=8oV>�֎>�g�>�I�>���=QŽ�$Ž`%����=��:>�0�>L�>���>"or>�r<ZZ;?�v�>p��a⾂�徫F��W�=v�}?�z}?n�2?/��>��C�
�!�����e9?�ڧ?�%�?��8?9|�=��={���L��.�����X>坁>�,;>�cA>숺�|��>�
�>�3�>�k�֞�y�3��#?v%Y?�k>�iο�u���ߌ�N����(�����u��U�(=�X��P�������B��8���Q���Tྡ����0��������#��6�>X�=���=�[�=�='=��$�p�;��>Ʀ=u^<��i��l���x��X?R�	ϗ���ڼ���F�r="���ƾzJ|?*�J?�-?8U@?��z>��>��_��^�>����?�0`>ae�Ș��M�/�VO��Փ���׾d�پ�`�wΞ�@x>�D���>��2>L��=�� <�d�=|�=�ۖ=e:r=���=\s�= )�=j��=�>#w
>�(w?���J���z2Q�d[�³:?�d�>��=&ZƾQ�??�>>�>��i����O�/?���?�L�?��?��h��R�>��<l��N%�=����
2>^{�=��2����>1�J>�d�>��h��N3�?��@z�??,Ƌ��Ͽ�/>�f8>lU>��R�*�1�H�Z���`�NPZ��S!?�;���˾�x�>g��=o�޾kƾy1=�6>a�d=ئ��\�Dۙ=�}�{|:=�En=�A�>;�C>���=�ί��=Z�C='��=īP>Dy���X4���-�eU1=���=Pb>,�%>�_�>ׇ?�]?M��?�,>L;�������Kþ��?��<�r>CM>����wA>h�`?L?:?	� ?��>t
 �'��>N�|>���Zx;�Gھ�Ӿa|�=��?�I?���>!�T>�)���j��f*��w��a2?ɌJ?8�?��\>�����F&��6<���z�-�"VH>�u�=5?5��c�k��<�gɽJ�=��>�ň>�څ>Jn�=t��>j�>���>
�*>��=t�G=�I�����Q0�Bl���U���?>s�>�8�>�#t>Q�ŻLF	>�8�=P`o<��м���=aG�>��> ��>lّ=m��<�3>B���J��M�=�Ч�VCA��yb�}ez� h/��@<��JD>7gU>!��y���^?C�a>�_@>V��?��u?�9>��y�Ͼ=$���gs��;Q�U��=�>�K<�=�;�j�a���M��Dξ���>
�>��>Δl>_�+��F?�i�s=CA��p5�e��>}_�����s��tq��=��u�^i�"��RD?53����=��}?��I?C�?���>��<�ؾ��0>]<����
=b���p�Cǒ��?� '?ր�>~N�$�D���˾�R��t��>jH�S[O��_���W1���4��c��ݷ�>���h о�1�sR���Տ�V�B�Nv�N
�>�LO?`��?8�]�^����P�R�Gᄽ=Q?|�g?��>�4?Bg?�����H���m��=�o?=��?[�?��>-�	>� ���@�>�f�>�/�?���?A6w?A������>��=1�E>@����=B��=�9�=w'$>�<?o�?�� ?��۽����
�V��Z���Y=�@�<���>���>#,>�	Z=��[=�:>��=�k>S��>�5>��>@�y>ʕ��&���*?�(
>Ŗ>��I?�ɑ>�>F���O�*��fܽ�Xj����U<x��"6��L��-�����=]� =��>�Ǿ�e�?M�U>�O�gv?�"�㽑=�?o=<��>��`���>��s>r>�D�>�ű>޼�=W�>>��>9F徥h�=� ������~6�$NE�?þ��{>닾�2�P|���=�l���ZԾs����g���y��}6�={_�?R�t���W���_��D?��>�5?�����L�喡=���>��N>چ��Ȉ����G���XՋ?fX�?�Fc>��>c�W??�?i�1��3�mZ�Ǭu��A��e���`��ٍ�����Y�
��ȿ���_?x�x?�uA?r$�<
3z>d��?n�%�Ϗ��!�>�/�� ;��<=;0�>� ��?�`���Ӿ�þ�P�X F>��o?�%�?xT?\fV� H�L'->i�<?�"4?i�n?��0?Y�9?s��X(?�>�%�>��?rC0?B-?|�?�*>��=������<�揽y��}�̽vGƽ] ���@5=�dm=N|��F��;p�2=*��<�ھ��@������0��¿�<Iu'=��=
��=0��>N�[?	��>�Ő>]u/?h!��G2�;t��a3?�+=p�|�4���䤾{��.>�jj?H��?I�V?0�U>y�;�̰D�{�>�V�>�%>��V>�ӱ>��ӲQ���=�>��>�s�=�P�y����������
F<��>��>We|>痍�hV(>�z��`z��d>�4R�,����&T���G�w�1�Ҕv�?��>��K?Ӷ?�9�=p0�˖�l:f��)?�v<?�HM?�?
ܔ=�۾��9�uJ�J��h��>LI�<C��϶��>��!�:�K<q:b+s>"����+���[>*���x߾?Uo���I�~�� *L=����L^=e�
�Ynؾ8Ł��y�=�}>]&���������L���I?��f=������U�V\����>���>�i�>l�=�_�l�Y�?�����r��=���>�.@>�f�� J��BG�̽��Ĉ>��C?˕[?��|?�0���u�XG�S��ܱ��/=x�?$>�>c!	?�>>�eH=�þ�T��ݪb� �9����>zV�>�i���K�Kh��/����%,�X�>s�?M*0>� ?ys\?x�?�\d?�v(?c?�^�>֓��课MC&?���?rڄ=.ս>�T�9�S!F���>ـ)?Y�B�̺�>&�?:�?��&?�{Q?;�?�>a� �D@����>>V�>C�W�9]����_>��J?,��>�8Y? ΃?��=>:5�<碾E�����=��>R�2?V6#?E�?ٌ�>��>A�h����=�?R�C?��?�6x?s$>���*?'��;�>ӣ	=a��>ݲ�>�f+?��i?��?5�C?ݷ�>.�w<#6�@��Z��~(��Ҋ���={�C>vYD�/�=�|��������?��acV��n]<c��x>��>d�>.�s>���1>�ľi;����@>]���O��!䊾�:�C�=ۊ�>�?���>Pd#���=v��>}@�>����/(?h�?�?��; �b���ھ��K��'�>��A?=��=;�l�~����u��g=��m?��^?��W�/���o?3�\?����a}O�퍟��ʾ
W��x?м'?Cx����>Nxv?�H�?*��>\.�~�=�D����/�e[Ҿ'>��>�e!���i���>D?B��>���>襋<tZ@��!������l�>�Ã?p[�?�Ms?g�>4�s��/�������­]?��>����!?��n;��ʾ�_���ď��p澾$���p���6��b#���_'��ˀ�(��9J�=��?��p?��s?T]`?Q����h]�kY���y�gV����"��lA�t%C���A���k���������ߛ�3�6=�3����K�/�?F?�~��?`���x��|���F6>���
x?�>([=0�1�v�G�K����C���|���x���D/?�л>@%�>�+'?״t�;mN�G�L�"*#����tʕ>y��>'�z>x?��Kc���U�����a��N)I�Vv>y�a?��K?�n?���C2�̑��{�"���Q�C����9>��>��>�#f��(&�D�(�b=�S)q��[��*����
��W�=w�3?��z>M�>�O�?{_?��
�����U���2���;�}�>��d?L��>���>��ֽ�����>n�X?�o�>Nnr>��ľ-l4�T_����;��>y�>%�>��>�ȭ��i^�5+���
��fI/��̓=�hG?^���W�ʾT��>ƚu?f$��#I���?$�����&���(����w8��M�>V�S���k)"�͡��`�E�	]�a8)?�B?Z��͚'�Ϗ�>��"?Yp�>k��>+��?
\�>'����9�?�_?�~J?}�A? ��>O<=:���2CȽ��%��L.=Å>Z>�l=�z�=d����[�^�߁;=j�=�pټ�;��b�I<=�Ƽ�:<]�	=�Q;>�lۿ�BK�X�پ�
�#�>
�$刾Ϧ���b�����lb��u��R[x�����'�vV��4c�ɟ����l�ކ�?/=�?,|��-��󱚿C���k�����>�q�͏�����P���)����������c!���O�&i�1�e���'?ӵ���ǿ���S2ܾx  ?�? ?	�y?r���"��8��� >~C�<�����ꘚ�e�ο^�����^?��>b�,����>���>@�X>�Lq>_��0Ꞿz�<��?ӆ-?��>\�r���ɿG����#�<(��?��@m�A?	(���[U=:�>3�	?��?>O/��c��Ǳ�)?�>y�?�Ê?+
X=�3W��=	���d?o�/</{G�����C��=6æ=K�=7Y��DK>�ٓ>���#�A�fٽ�5>� �>�� ���H�]����<m[_>�}ҽ�c��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=1��͏���#&���1��w=���=q_>�ȍ��I�=���<��E���}¾0�;�\>K��>WҪ>�6>Vq�>T�=?'�]?6�?�j=>΄�=�0�����u�<��Z�ŹM����؂0���о�d��B�?�̾7��:��YQ̾��O�
{@�[ `��B��Q44�p�_���.�'�)?�]1>󅶾��3�1���0�ZX��5=khʼ�ʦ��E�fa�Ί?�"?8����,W������B��H��^B?���7߾����k%�<�,����=6��>O>��޾�D��K��IC?|d?#�޾
�P�h��>�/�DSH=�8'?��y>Z���P>�$?Ilo��3>�k1>_L>czb>$'?N*�R`���8
�S?�V?��D�v�<�H��>�X �R���C>�$K>�Qټ���=$��>�S�=�pʾ���=�P�<��u>o(W?��>�)���_����U>==�x?��?�.�>M{k?a�B?9�<ne�� �S�v�(Ww=y�W?2(i?θ>\���{о�~����5?�e?@�N>:dh�p��m�.��T��#?8�n?$_?�����v}����<��mn6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>��������=������?�}?eò��/=D��AIP�,+����=ǒu=8>����=z��2A�ǥӾ����ؘ��1"���>,@��e��>�Zb�t�ӿ�̆���ɾ^�����(?��>��s<2����b�&Gq��X4�n�M���k��'�>hT>���n���M�|��X;��|{���>�/ �^I�>|N�o[��(���+�^<�0�>���>\*�>����d
��1=�?�k���οq���2�=�W?�?=��?�?c�|<�pr��4���Y^�9gF?O�t?^�Z?4�*�-d�5�:��j?=_���T`�i�4��HE��U>&"3?�A�>W�-�\�|=u>���>�f>2$/�b�Ŀ�ٶ�%�����?���?�o����>c��?�s+?�i��7��uY����*���-�d<A?2>^�����!��0=��Ғ���
?_~0?�{�.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>2�?�>�=�q�>ȱ�= ڷ��W�ɼ'>�f�=򭫼^�?Q?A��>@��=,WG�ro.�oqE��P�R���@��;{>?�_?CpL?[(I><g���}E��0��gʽF�:����0!J�x�/���佫u>@�*>��>h�6��ξ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*�̿�������+��mc
�*S=8�|>p��i%>��=w�= H�����;��>\�l>g؄>��>d��=��B>��I�%��F۔���z�_/�w7�U�X��
��
��uݾ���	�B��ZIC=B�<k�"���پ�'�w��=t�U?�Q?�Ip?� ?�Zt�g >�����=�($����=JV�>dh2?��L?ީ*?�̓=D��O�d��@���X���������>��I>���>~4�>d�>�Q��J>��>>0��>ġ >�+)=��,�\�=��O>^S�>���>)��>_�;>��>Ŵ�y.���fh�yw��˽��?Uߜ��J�� ��D���ꀷ��.�=�t.?��>1���(п������G?�Ԕ�e��H+�l�>�1?�8W?e�>G���W�Ee>�	��l��=>*���T�k���(�=�P>��?�bf>��t>��3�=o8���P��d����|>,6?eζ�F"9��u�I�H���ݾ�>M>D�>C�=�(\�x�����~�|gi�z{=�n:?��?�²�gŰ�&�u�HE���0R>�:\>��=[�=I-M>�7c�n�ƽ�G�(�.=>��=�^>u[?�_,>���=V��> :���}P����>�YB>-�+>5@?1%?���o���.A���.�v>��>���>�>qbJ�\�=.r�>�,b>C�i6�������?��_W>��~�yr_�V�v��|x=>���$
�=��=B �K�<�)�&=�~?���(䈿��e���lD?S+?_ �=��F<��"�D ���H��F�?r�@m�?��	�ߢV�A�?�@�?��I��=}�>
׫>�ξ�L��?��Ž6Ǣ�Ȕ	�,)#�jS�?��?��/�Yʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�k�#=Q��>�8H?�V����O�g>��v
?�?�^�੤���ȿ4|v����>X�?���?g�m��A���@����>:��?�gY?xoi>�g۾9`Z����>һ@?�R?�>�9�z�'���?�޶?֯�?�pa>u݇?�Wd?՛>�����G��X��/�|�\�J��
<>���>?��>y��!�E�X~��~��H�X�z���X>�=i=O�>�ë�����D�e=����N��g�N=�е>�k>�"�>2 j>�y�>�?�"1>ӀO=�f��`e>��0����[?���?�L��t��@>ɻb={ ���J.?��?���G��/�>��J?��b?�B?D��>����n��O�׿�����[�hZ>�~?W�?�^>s��>Y��?��H�u>��>�4_8j��3S�6�2���R>$<K?�u?�3�=j�?.�?��>B�>�<������M�ً�>�gJ>��I?�~b?5?V���}�:�d7���֑�?�O��8>��l?V%4?���>�󔿩r��g�Q>��c�S����$�?Q��?J�n��F)?Μ?��H?��N?R��>F`o>�8�(�7>Z�u=r�!?3(�S�A��Q&����}?�O?���>�"����սdּp��������?�+\?#E&?M���(a���¾��<��"���R�0 <v�B���>�>����q�=K>bӰ=Fm�IO6��g<v.�=u�>�+�= 7��M��/=,?ǿG�{ۃ���=��r�@xD���>�IL>����^?ql=��{�����x��!	U�� �?���?Yk�?\��?�h��$=?�?S	?k"�>�J���}޾7���Pw�~x��w�T�>���>7�l���K���ٙ���F��]�Ž�\/�
�>�v�>4i?f��>��+>O�>���4�*����Z��;�V�"q��3>�n�4��#��w��H-�۾ĻKO��`�s��-�>mƀ�ח�>o�	?�`>~��>��>f�}<��|>^8=>ݽ�>�8�>v�C>�\->CW�=3��
ߘ��NR?߬����'�s��PM���1B?�id?��>x�j�������(�?��?O|�?tZv>�mh�!+���?���>�$��2^
?�q;=[i	��X�<W*���s�\އ�Ҕ���>�׽:�
�L�z'f��t
?�?^a����̾�xֽ\V��ERm='��?�$?*e,��P�`m�C�N���c��=�<��e����d.�;�w�o��/l��5����(���Q=�,?�V�?���kw�*g���~�!�F��>>A��>���>�>-;�>��=��^O��!�y;|��0�>��u?���>o�??�H? 3p?n�f?W��>��>.*⾗��>��L�H7Q>�?��0?]j?37?���>��<?uD�>�������Վ1?��.?��>u��>J��>@ɾ3vq>�l��SM�<$Ux��0<q!���ĕ���<]l>�ε��m�>[�?�>��#8��y���|>2�6?qx�>h�>�ە�kN��U��<��>�*?.g�>������o�a�o�>΢~?���^��<ݔ/>h}�=��s�}Y�; ��=A{�׉=�>`�60�B}�<�D�=�<�=dU$<h�p�"�7<(����Z�<�t�>/�?œ�>�C�>�@��8� �`���e�=jY>WS>F>�Eپ�}���$��y�g�u]y>�w�?�z�?!�f=��=Ԗ�=�|���U�����B�����<��?4J#?*XT?\��?j�=?^j#?��>+�dM���^�������?�,?Ƈ�>u���ʾ=ِ3��s?�A?L6a�V��f8)��^¾m�Խy >Ub/�Q9~������D��_��-��EA����?sŝ?T�A���6�u辝�+~���zC?G��>�,�>���>��)� �g��E�nd;>7p�>�R?�U�>	P?��z?��Z?]�S>!�8�[��f��pa2��r$>2�@?�ׁ?�͎?J�x?��>YZ>�}*�#����1���`��Q>����W=�W>���>���>K��>�Y�=��ɽ�"���?�x��=�qc>���>�٤>���>��w>N�<~�G?F��>�_��a���⤾/����=��u?뙐?�+?0=v�|�E�/B���H�>n�?���?Q4*?��S����=��ּ�߶�T�q��(�>ܹ>=4�>��=�[F=zl>[�>3��>{+��[��r8��fM�~�?F?�ʻ=tIȿ����<��U�۾��B�Q�F�um=�J���s̽�5>$������{�$����R!<��=��S�0�������>%�=�U+>�.`=�]Q>t�$>����?=�{;��V=mW�F�9=f"��zн��>�W4=s2��T�=Vݦ=SK˾ɓ}?�&I?�U+?�C?2y>>>�2���>%���^?]�V>�7O�Qi��5�;�����\5��H�ؾ�s׾��c��П�]b>��H��<>c]3>v�=�؈<N=�=��q=��=�|a���=���=� �=��=��=��>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>mcB>V
>1AS��w0��D�9KY�s�X�Q#?��8��Ҿ[��>�w�=`Mܾ���7=U;>X�Q=��
��a�7Y�=����*D=��=��>��K>X5�=[�ҽT��=Շ=L<>�TT>�#��+��bbO��=g��=/t}>�y<>3��>�c?e�.?&Yf?*��>�\R��U¾��ϾЕ>G��=z��>���=G�O>Ҵ�>%�8?�G?�Q?f�>�F�==�>է>?T,�RSn�};���y=6o�?v-�?$�>��*<u�J����:�;�@���?T1?��?)�>�����Iv(���/�+���i��:K5F=��q�ǈB��Qͼ{��s��HD�=c۩>��>ۣ>G�y>��.>a�P>���>�u>B��<�}=�G;���<jӡ���=�;s�o�<���*|�_K޻#�B����M�;��V;�8�<�c><���=���>cj>��>�= ��#/>�Ӗ���L�
�=�b�� B��2d��U~��/��6��B>+X>�@��.��p�?Z>�?>Py�?-u?�H >U4�@�վG��*]e�}S�V�=x�>=���;�vI`���M�DnҾ��>2o�>�o�>�>sa4��G��x�:E����_9�"�>sS���%;��F"��D��jि�.^�Ѭ+�'�@?�����KA=m�|?�HP?��?Q�>�=�=�,�&��=W�w�f�}y��2��T轔�?b4?q�>9��T�5��ɾ�<��K��>V�@���P�����ވ/�{������"�>�ܬ�
pо��1��a������D�}�o�w�>��O?>�?��^�^�JO��l�?x��?Ȑi?삢>�? ?�r��Xt㾪�s��k�=�9p?f��?&��?L�>>!�=�Wh����>�?j�?��?Ls?�n����>h�ü�w/>�>��lM>�>��=[P>M�?�/
?61	?k��|I����i~��mRb��o�<�(�=1��>Q��>��n>x��=�=���=)SP>?	�>3(�>l>ُ�>���>l�ľ�F��:?���=�j�>��=?��>T��=����w�*�A���8I��Ql�����]:��d����񽊯o=�l=�'�>[Ⱦ���?ߦ/>T^
��?���-=�=b>�$�'i�>*	�>�FA>䠘>.�c>x�R={�>�>0BӾ��>���d!�w,C�*�R���Ѿ�zz>����?�%�?��V]���:I��o���h�;j��-��p:=�2۽<�E�?������k���)����[�?_�>�6?}܌�q����>���>TÍ>�S������Lɍ�=dᾴ�?^��?�;c>��>L�W?"�?�1�_3��uZ�.�u�v(A�e�U�`��፿����
�����_?�x?yA?�S�<7:z>M��?��%�eӏ��)�>�/� ';�A<=v+�>�)����`���Ӿ[�þ�7��HF>��o?5%�?wY?$TV�Yt]��He>��:?�CS?�vf?��B?��8?�Z��֯;?)�=!# ?�s?q�:?ۣ1?�u?�wx>��p>�U�;:ʞ=����2�I�|S��`��e˽F6@=�.�=@�z�c=�b�<	��=��J��m<�!ӽR;����>�A�=�i>FC�=�M�>�'^?\��>ӳ�>(�6?f���4�鱾X0?��&=�&���c���ß�I/�x->L�k?��?eUZ?��h>��@�1ZB�>�>1ƈ>>�'>Q�Z>�m�>�Q޽�VE�_�=�
>��>��=�\D����	�S����=�z'>���>�2|>�	��a�'>�{���3z���d>g�Q��̺���S���G�=�1��v��S�>��K?$�?Ց�=�[��9��OHf��+)?u]<?vQM?��?S
�=5�۾Y�9�@�J��>���>�:�<&�������#��0�:�)}�:��s>�,��
@��(ZR>�	��O㾪L`���8�X��op�=�|�S1=�����߾=Hm��a�=��=�ľc��j��g���H?�;E=�i����w��	���M>Af�>�ͬ>�6@�:gb��g=��հ��'�=���>�U>m<[5���D���ş�>��A?�qT?��q?�Z� t��M��o��{<Ѿ࠶=��>h�b>��>�8A=T�=۾�G��7o�!c/����>	?+�8�\�l�,���B���(���>�D?��ֻ:?XQ?e�>E�Y?�",?5��>�O�>g~6<�t��b'?p��?&�o=�
��*G���9�1%E��|�>�Y!?�M��ϔ>,M?��?�&#?kR?7x?^��=S�����?����>�5�>�[�,<��P�o>��G?훷>�U?�?",>�Y3�����6�½+>�+7>�V.?`�?J�?\�>l��>Hn���=�D�>@�W?f�?��n?^��=[�?�&>)X ?�!�=an�>�.�>��?� P?j�p?NJ?���>W�_<��޽��4ѩ�	�μ:�;J��;��=Q�ڼdH��/�J�<; a=X�5�qL���3��V��\�M�N����>
�>�bq���a>����qr��h'^>$@��\��eÆ�R�	����=�S>�K?�ĩ>"�ֽ�Q�=B�>X��>�� �3?��?#?��I�]�S�����9�N��>�4?�R�=�Dk��3����~� �x=�Px?t�O?Yu.��o�+�b?Ջ`?A�G����}�"����3J?n��>&�;���>��y?~_Z?k�>ƘF��l�����_�`�Cē��X�=�d�>[
 ��j�{��>�7?`��>��N>7M�=	I۾a�s����q�?$�?�q�?ш?��>�rT��H����$����I?I��>,W���9?%��<@���o��c&���c��"�y���'n��;9ž,6I�=�i�*8��hN=�3?A�t?��p?�9T?�྾q`���c�I�k���Z�(�� �zR��;K��!6��\��<����Yg��T��<n����H��<�?[�?ɥ��G?(̅�������Ѿ@Q>	�ݾ���> ӂ��ɺp��<�2��n$&����{�$?�g�>���>�h?��g�a�O�)�8�\O2�Cz��K�S>���>�k>���>BIZ<����ҽN��9��ʽ.2t>WU?4�&?ocP?R��S,+����;Q)�A-����R��>�7r>�[>����RH��'�-�I�^�h��t�g�������>�",?��>� ?�S�?�~�>*�)���7�Ծ)�/�E�����n>X�s?��>�`>�����������>��i?���>t��>P-��T��5z�����>9ǳ>T�>�;r>"-A��`�|���
Ǝ�n.;��H�=��d?HE��� i�(�>�,P?ݕM;��<���>>����&��X��W<��0 >� ?���=r_B>��ɾ#�
���.�n��7?F)?X���m��ה�>�Y?0��>LRu>�Rh?�~�><茶�S=w�>,�k?GKD?w*?�S�>/绬� ��Q���*�e=Vݘ>OxI>�S`=�R�=������� ���Α=���=58��@��V=js<.΢=�W���gc>�ڿ��K��־��ͣ��o�v����n��F����	���������q�����%?���W�6j�*���>q����?h�?�J���@���Z��Md�����l�>�jt��a������	��N���߾�9���o!��|S���j��2d�Q�'?�����ǿ򰡿�:ܾ4! ?�A ?6�y?��6�"���8�� >HC�<�,����뾬����ο?�����^?���>��/��q��>ߥ�>�X>�Hq>����螾�1�<��?6�-?��>��r�0�ɿa����¤<���?/�@�,A?В(�3��R[=f��>��
?SzI>��� �����-��>�?G��?�n^=��T�9M�ne?��<�@�������=p��=�= � CR>|̑>S�N�8��g���0>D��>�������Qo���<��e>թ齭R��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6��{���&V�}��=[��>c�>,������O��I��U��=�7��[~ѿ#UW�m7�J����=�
�>��̼���=m����������:}�=��(�Q篾��>�?(�>CDP>8E?F�E?�(�>���>�m>�x<񶩾�<��:g��z�X�P�q�\�b����o���a �t�
�F˾[;�Ҿ�$�=�>�F��:��#v�4�e��tP��'?k��=tJ���^B���<k�޾�����%�g�g�Ͼ�(7��o��j�?�Z@?�H���p�>�����J�3����=R?�ƭ�����<��8�5>�}�cf>:�>��=Ǿ6R��9q�Ā>?M�?�Ӿ��'s����>O�ڽš����?m��> +�=P(�>�?JӉ��	<>O�>��Q>��>`�t>���<h���Y�M�H�?"0(?�5h��>{�F�>:읾y���#�=�9�=U��j�=�tM>���;��t�7�=��b+�=pVT?���>��-�U�$��,����d��a�=[z�?Vh?��>[�o?K;?���=C>ܾ�D�38����=Pqc?��q?C>$%��w�$���f)?6Rd?Z9>��@��lѾ
m�k���{?�u?�G?Z���r�􈇿�
���&?��v?s^�ys�������V�d=�>\�>���>��9��k�>�>?�#��G�������Y4�"Þ?��@���?��;<��V��=�;?m\�>ޫO��>ƾ�z������>�q=�"�>����wev�����Q,�^�8?٠�?���>�������{�=������?��W?��ľ���U����:��)�Q��<h�ƽ���滂=��վA�B�G��f�7�󒯾�f�T/�>|?@x)�x��>����� ���nݿ� ��>a��	�μ]D?�p?t=�;s1ܾy`�N�o�[Ef��X�W�H��ԣ>�>����n��1{�I�;��������>���Ż>��Q�[��5^���=7<.G�>b�>]�>�߫��a��|�?�����)ο������ZX?n�?GL�?MP?��D<�Dw�$�z�5��@�F?��r?w�Y?b��T�Z�ֳF�$�j?�_��xU`��4�sHE��U>�"3?�B�>O�-�Z�|=�>���>.g>�#/�v�Ŀ�ٶ�7���Z��?��?�o���>o��?ps+?�i�8���[����*���+��<A?�2>���C�!�B0=�]Ғ���
?V~0?"{�f.�]�_?(�a�M�p���-���ƽ�ۡ> �0��e\� N�����Xe����@y����?M^�?h�?ֵ�� #�e6%?�>e����8Ǿ��<���>�(�>*N>\H_���u>����:�i	>���?�~�?Qj?���������U>
�}?J�>d��?{x�=�4�>�-�=%����4�5%">{��=\09�Yt?+�M?���>���=`*8�/��#F�8RR��
��C��ȇ>��a?�zL?�/a>�����,��!�:@ͽ=;1����T�?�z2.���߽��5>Ԕ=>�>�E��!Ҿz�?z��ؿFj����'��/4?3ȃ>��? ����t�	���:_?g~�>X9��,������ܘ�?�@�?��?�׾�̼�>��>�M�>q�ԽC,��9�����7>3�B?���<����o���>��?P�@YϮ?�	i�\	? ��P��_a~�o���7���=��7?a0�C�z>���>��=�nv�ջ���s����>�B�?�{�?���>�l?u�o�E�B���1=�L�>��k?�s?rxo����B>��?������L�Gf?��
@qu@$�^?-�0Ͽ;��wķ�����ޠ=V|�=��K>,�e�3�=�.�<�Hm:?��
�e=�v�>իg>��X>�z>��@>D�e>�@���=)��.��f��5�O��B��������wĄ��?�l���40ھ�O��-綠LK�/�[�N�-��+X��>j�R?^8J?p?e?��?%\P���>�5�����<�W޽ډ�=no�>UX(?�R?�^*?���=�S��bWa��z|�_ӫ����l�>Q|]>�=�> ��>�ƿ>>�k�Z>��,>ݬh>$�>�W=ࠩ��9@=�D>˫>��>aż>��>>�:>ٌ��qS���tg���w��(ҽޕ�?l7���J�{��:���θ�:ߞ=U_.?�p>�呿
�Ͽ4��{�G?�����-,��3	>�0?OoW?��>������S�l�>$l	��j��r>;��B�i�;h)�(�S>O�?ںl>�x>��3��99�R0M�������u>��3?�*���u5��u���G��{߾AR>���>��^�ɣ�qE�����gh�ѵZ=�9?�`?] ��r���>(p�î���xV>�z[>v�=׻�=EL>[=�M�ɽ�%C�0c0=p��=8�b>?�7>l��=
�>�*����[���>�/w>�+N>;�7?��#? �U���`�\�h������>�>�>ȄE>hU��>=��>�C@>���$?�����6�'~g>H��j�d�����F�=�A�Q��=�g=��>�,�1?8�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�i�>�|��Z�������u�9�#=��>�;H?�N���O�d�=��v
?%?X�覤���ȿ@vv�h��>��?��?J�m� A���@�Y{�>��?�dY?0vi>C`۾�JZ�^��>��@?9R?�>�=���'�;�?�ڶ?���?8`7>��}?�_?U�>�ꜽ5�4�����s���������>�me>r6->�Q����f��́�"S���N|�(�>�u%�>FW=i�>�b_�dݓ��?�=�k���ɾ��<���>Q�|>��B>d�O>���>+E�>�q>�=vY=a��7gJ�ȽM?,3�?�j�t�o�qd=�=�k�I�>
;,?�qú)=Ѿy�>�P?6�?nY?P�>�7��i���R���m�����]�G>��>nB�>�h���V>�wپ�)�f�>-[�>I��9�Ҿ-�\��NG����>�?ב�>�%�=/�?�7$?T�i>���>H�A��^���H����>/c�>^�?nz?3j?Cٺ���4��R��5���T�[�w�7>�s?�?U�>A"�������\�u���sc�?ӆg?�����?��?m�9?��A?��v>�	�^ξ����a�X>E�0?Y�<�{-C�1�*��M�=�J�>Dx�>t��>����ybC�gR��n�Y�bW?I�T?�H?���O�(t���d�;�ӽ/>�����=؅=�Z >��%>~�½R�*>��>D��=\JF��R���>�=�?�>�)�=w�Bs=/=,?G�G�rۃ���=��r�=xD���>�IL>����^?`l=��{�����x��	U��?���?Xk�?]��?�h��$=?�?R	?f"�>�J���}޾4�ྭPw�~x��w�X�>���>�l���H���ؙ���F��Y�Ž��f�A��><��>�d?�.?���>�D�>9�u�)�.���̾�� ��{k�����F>�2\6�u6�5�����6����-,]�>,�>w1½�ě>F|?[�k>��>X��>+����"=�'>1ռ>tz�>EQ�>1;Q>Q�������ʽ��Q?d>���n$��X�X9��A�<?I�e?��>�?D��B������?�n�?��?A�>(�e�j'�w�?�C?�}��$?w#=�/}�z��<|����-��Z��&�qj�>��佊);���I�Hp��?��?�d9�j�̾ �н�ȼ�=$op?�j?-�'��<e���|�'�Q���^����=Gn��O�����E�r�L���=-���+#2��MK;/&?�6�?���c�ɾ�Ί�W{��I`��[�=�%�>��>�?��>�X׾r>��A�`:���3�,��>S.y?O�>��B?�s?e�?��	?�9s>��>A���,?^f;���>j��>�x�>0^?�GF?��]?	�?���=������'F��^3?y?<@T>�o�>!�>Eˊ�#q�>��l�o�T='��Y���d˽A��=]6>A䘽JM>8ā>�6?�)�c�<��I���m>�%9?���>C��>������z���f=\|�>Q?Rđ>�����m�G��7�>Hp�?���)D�;S�>QE�=D�ȼ�T<�b�=�%Ļ��=��;��F�|$}<���=*��=`W�|!��|�<N�y����<u�>3�?���>�C�>�@��0� �R���f�=�Y>/S>�>�Eپ�}���$��k�g��]y>�w�?�z�?&�f=��=���=}���U�����8������<�?=J#?.XT?X��?k�=?[j#?��>+�hM���^�������?�,?n��>@��;�ʾ|먿�3�7�?�L?�Da����57)�+�¾�>ս�u>�V/��2~�m��7D�5��0�����??A�R�6��p�����j����C?��>�V�>�	�>�)���g�$$�0/;>)k�>&R?�!�>ZO?��w?�UY?;>W);�����*���Ư�y�E>��F?���?���?�h?��>!>�{<�Qv��6��N&���t#��w�2=�_>D�>�C�>��>�0�=d�ҽMc��
2�3�P=��f>���>���>Y��>z��>����TF?��>�l��E���죾7Ȍ��m<O�?2��?S�?�.�=�r�¢4���j�>F[�?�٨?A�8?�۶����=���/�žb�,�>���>w�>�3�=�+�=H|j>�m�>>T�>%w�F���xB�Ns���?hw7?��V=��ĿϚ��8(��2`��%7��>�(�Rg �~!=���:�f;=��G�?�i�����Ic���✾n�
�p�@��2���e ?�=�>�L%>[��=��A=����1z=��~�d=Y1޽�
���<cJ =�����R5����O��<�x���S˾ o}?2I?g�+?��C?F�y>��>�6����>����?�.V>G(T������A;�䨾�W��?پh2׾��c����n�>��H�Z�>X�2>���=P�<��=�0t=tٍ=��d�P=��=�͹=?��=^��=ak>r�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�z�>?R>��Q�b�A�����Z����zA ?1�ᷠ�_h.>Z-�=P6�R v����=u��=l*�n8��o�q�=�F�����g�>�S�>7�]>g>|t���/>�R=ټ�=$>q�:�>^�=������=��=*}>�U>Q�>
�"?O�3??�C?,�W>u�Ǿ��Ͻ�8���k�>nԠ�;5 ?'�C>2w�>Jk?��`?��-?��7?�3)?�L�>�+�>I�!>S�7���H�^���D���K�=�ۗ?�IL?zŖ>�!�(l��/#�ewR��.�>^�?�?�>�>9��c�5�47�Po9�B1ƼL��=SI�Q$=��g���	���>�ӡ>�n�>U��>�U�>�G_>�|}>z��>��C>��w1�<�-���z<q�E=�|��0�;���X���n7�=_�=��
��B�3>���=�`>Np6=J�=L��>�7>�`�>���=�_���r'>-���N�T��=Ԥ��'@��d�����-��};�O
9>�9O>q7��0ᑿ� ?'J_>4C>V��?�*u?/�,>���J�ھww��y�o�P9U��6�=��>��3�^ <�t�_�EHP�mt˾���>���>gϢ>�q>�{)��<���Y=�h�)�7�9o�>������S��c1s������ğ�=�i�lhd�JMB?U����*�=�_~?
I?�Î?Q��>��x�öپk>�V����<PN�||��Д��M?�"?��>�Y��>�?�˾l����ٷ>I7I�^�O�!���#�0�g�d��c��>������оZ3�lh���叿N�B���r��E�>��O?��?�;a��r��@�O�?��ㆽ�1?�g?@y�>��?><?{1��u�����.�=p�n?���?!/�?��>���=[���nC�>3��>��?0ˌ?�t?J��uE�>�UʼlY>fa|���'>V�">>��=S��=�?v�?��?�����P�������b_�Xׇ=K��=|�>�&�>�{�>��=f�f=uM>H�I>��g>AI�>�>ǩ�>��i>?*������?��>��>�_O??ǉ>5q>�ս���hL�����j��JZ���8*�Ҝ༚8;�=Q���wb�>dR���i�?��=H��>?e<羅�I=��(>�:/>)��]�>�_r>0��>	��>A�>l�w<��>�>FӾ	�>w��Md!�z,C�w�R���ѾEzz>W���&�����u��*AI��o���g��j��.���<=�!ɽ<�G�?;���Q�k�U�)�0���y�?Z�>�6?Uی���e�>���>aǍ>:K��ꏕ�ȍ��f���?1��?�;c>�>A�W?1�?ܑ1��3�vZ��u��(A��e��`�w፿؜��b�
������_?��x?�wA?�Y�<i;z>>��?o�%�.Տ��)�>/� ';��K<=F-�>r+����`�ǮӾ�þJ6�IF>��o?%�?�Y?�WV���ӧn>�`?��S?i2L?=�-?��;?\��.�G?��=�)?��?�r?[&?r�?-�>"h>q���M�=�$�����`�o�������Q=��T<-���of�<�߹;#�=����˿���>�Y<D:ʼn,�=�Q�=��=J�>��\?��>�Ɉ>��,?��@��$��҇�E0/?H���ZI��/q�(J��f�о�9>Ub?=��?��e?1��>�:��)Y����=K�}><%>!]>�v�>��x���6�d��=ۆ�=��=|�=|0���Д�	��7��@	�<�A3>*��>�p|>7����(>�a��hFz�}	e>�9R��V����S�[�G��1�w��c�>��K?�?V��=�F��ڕ�(Kf�G)?R�<?hM?`t?e^�=�r۾p�9�g\J���3	�>3l�<Y���͢�K���]:�ĭ�:K/t>V	������1La>��ľ�%� �V��^:��q��`���+����;���˗�$=V���>5*�=
�þ;/�Jě��{��I?T˟=4���^�9��7B�=V�x>��>D�"���7��Q���+:P�>�>�ༀ�Ծ!�C��M9�>@PE?<X_?ni�?� ��ds���B�<���/d��]3ȼ��?E{�>dg?�B>�=t���5	�%�d��G� �>���>*��m�G��<��|.��Z�$����>�4?��>��?��R?��
?��`?*?D?7'�>������B&?��?��=�Խ��T�� 9��F�� �>�)?��B�q��>��?W�?p�&?��Q?ɶ?��>�� ��B@����>qY�>��W�Xb����_>��J?q��>9<Y?�ԃ?5�=> �5��뢾�թ��Z�=>��2?75#?P�?x��>�.�>F,����=�?>/z?�=�?k�?U.J>I�#?�=f3�>�9�>n%?52?��1?1D?�;^?K?���>���<�K���Q���K���$ҼU�<^e�<j��=�V���E��o��� o��^N�`�s<�cź�yO�G&���������<�$�>މv>������;>��ƾ7/����I>}Ӽ�v���#����A�,�=�{>���>̔>�� ���=�K�>T�>`��'?�z?Q?�q�~�`��;׾�zT���>+�B?���=6hk�ٓ�aCv���T=�l?��]?5P�a����b?�]?�g�R=���þ��b�މ���O?��
?��G���>��~?�q?>��>k�e�c:n�@��Db�@�j�>Ͷ=�q�>9W���d�f?�>I�7?�O�>��b>�#�=�u۾��w�*p��o?�?��?���?�**>R�n�84����n����]?3��>1��o�!?#�;�8hҾxʇ����������醧�,����w����%�������k��=�Y?c�u?<r?[�]?����c�6a�}ـ��W����A'��A���E�$jB��in�k�����5����<����<��w�?��?���,��>��D� �4%־��F>" ��"n���=.�̼��<�ـ<`���9��eӾC!?���>u�>�"4??(X�QO6�D�:�&7�2%�ǫ&>^֣>9 �>_�>��h�`W��L��j�ʾ������νˇu>K�c?��J?�@m?�`�`Y.�+���Փ!�7��L���(J>�]>K��>��_�6�&��C(�!�@�}2s���桓�f2���=�/?�S�>��>�֘?x�?�
��㬾𿈾p,0�%��<$m�>�9f?���>���>Tɽ�$��T�>ԟ?&��=И�>n�C<���#��aނ�M�?q��>l�k?��=�����9�e|��x��S��� >�k�?��˾y�"����>�Y,?�;m>��=�#�>5�	x��Z<)�-��=)�>Ÿ>��]=:aP>B|��Y3������B�M�!?�a?C���/4�$Z�>�/??v�>a��?�ZU>�/�����<�c?ۑi?g�W?��D?L��>}�v=p�|���Ƚ�B&�A==8��>��d>�)/=�s�=K?��N�Z7	�"y="(�=/�5�)�Խ/$;���8,�<m�,=nG>�l׿��G��ȣ��"
��uȾ>��v���ɘ��B=��L�����~V�z�*��=����ϼ�Q��H��0o�������g�?y�?g��j�k��󖿿Ā�:>"�Z/>�q���Bֽ Ǯ����ް�u׾�ľ�k,�"�i��:��,Ń�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@̔A?��(����'�Z=R��>�t	?�E@>�{/�я�����G��>��??sH=T�W�)���e?	i<$]F��׻��=6�=Y�=X�OQJ>�^�>����>�q�ڽ�k5>�k�>�c�(��_��ղ<:I\>ڻҽ�o��85�?��M�c_j���1�]1�� ->��L?	��>LӾ=��?
C=���ѿ`�`��|b?���?Y�?a�'?�d¾�H�>�ؾ*�D?k0?o�>�N�_o��|�=#����.�����K�a�>�u�>�:�=W.K�o��;7�3�>m�=~( ��"ȿ+����?�=���=ћ<��
��n%<8C����Y�;��S
��5>LS.><(p>Dt>g�>_Q>AV?�Du?���>hD->��=�-K��A���
�Ͻ��`���۽�%���ս�ʬ�v8����o���#-�`6-��h�I!=��=
5R����p� ���b���F���.?v$>��ʾD�M���-<@oʾc����܄�㥽�/̾��1�N#n�?͟?�A?������V�x��^]�勹�ѭW?�U����Nꬾէ�=+ϱ�K�=
$�>���=���X!3��~S�+�0?VI?iXƾ������ >	!
�C�=�)+?2�>�p	�C��>��?�/1�o��:OZ>��7>�+�>-��>�>}����ؽ�b? �W?�2��%���>�<����|� ��=0��=vQ&��j����G>fu�;�}��c� �����|�V<�=_?���>G�=�-����6B��-��A�o?���>ؒ�>x�W?|A?9�Y=)�c�c�.g�L+>ީn?��_?�Ĕ=�k5>�ľ$�����I?�k!?�G��\��`�;���ߘ���6�>3�S?A?� ��n���,$���ھK,?��v?�p^�2r�������V�=�>�[�>���>u�9�tv�>x�>?]#�D�����,Y4���?��@-��?�<<a����==3?�L�>%�O��9ƾʠ��݁��fAr=��>�~��1bv�1���9,�+}8?}��?z��>Ł�����t|�=�ٕ�LZ�?��?���-Vg<y���l��j��"[�<���=o��(3"�C����7���ƾ�
�����(���j��>�Y@4轩'�>cO8��4�!TϿ���
bо�Tq���?q��>X�Ƚ����~�j��Ou��G�}�H�ୌ���>��2>�rѽ����v���h�U`�
. ?��e��Ĝ>���^t4��O�ս���>�
?Ր�>5č=�&z��C�?E�;wٿyh������`U?��?/&�?��>��6�� ��Gx���ڌ�Z�~?0G�?B��?�>�=��˅�=�j?8���[`���4��>E�aU>	3?�E�>��-��R~=�9>SZ�>n>�/�X�ĿCѶ����e��?&��?gl��>�t�?]+?�?��5������^�*�hH��3A?�2>����f�!��(=��Ȓ�K�
?�H0?��M��_?j�Y�xzs�zm0�҉��漚>2���E�q��?R7���_�bP���-���p�?�C�?��?���)�!��&?�>����ɾ}4�<E�>(}�>��H>�5��[[�>����2�V3�=���?���?��?�����|���E�=�D|?�w�>�i�?tw'>��>تe>�o��/4���\�=Yw|>H���?śP?���>�}3�7싾�A�f]�Q�X���׾� D���o>�"i?�+? ��>]N�j:>�9��29�1z�������6�f�Z=z$�p:>AD>�+>^z!�_F���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?z�%L��W~�C���E7�Q��=K�7?�)���z>��>�ߪ=0qv�#���d�s�Q��>�?�?�x�?ټ�>��l?�vo���B��Z1=�J�>��k?{?��`�(�xB>��?���F���;��,f?+�
@�u@ƚ^?�좿�ѿYf��Y��������>�=�= �N>n���>�G�=���:'=�Y:>Z�>�e�>C[n>�F7>�y9>��1>�����&��q���-���
2��g��N���^��v��hO��|������[����r�C�'��,���;��t���M<<H�=S?�uS?��k?ix ?y�f���>����D�<�	#���`=0�>?�0? K?M(?��=TF���jf�u4���o�����[��>*�E>k�>�W�>�p�>�L<�+C>�3E>�?w>��=�'=r�;2=g�K>}��>&p�>��>ND<>e�>Gϴ��1����h�/w��̽&�?"���|�J��1���:������Bl�=�b.?]~>����>п����2H?�����)��+�$�>��0?wcW?��>L����T�L;>����j��`>�* �!~l���)�q$Q>}l?p�f>u>�3�a\8�/�P�s��%E|>�!6?����oN9��u��H�fݾ�mM>+þ>��B��`������
��ai�ܜz=o:?d�?�޲��ΰ�T�u�;��
R>�q\>X�=na�=`BM>�c��*ǽ�%H��.=���=�^>�
?Pc7>�<J��>����pVO��R�>�>>��>w�B?i??��U��������W�ր^>�w�>���>ƕ>Q�K���>BX�>݋L>@��;D[��z7=�n�V��Sv>�N�U`B�?ѡ��'�=�͡��̾=�m�;�86��� ��m'=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾSh�>�x��Z�������u���#=R��>�8H?�V��y�O�g>��v
?�?�^�ߩ����ȿ/|v����>W�?���?h�m��A���@����>9��?�gY?�oi>�g۾+`Z����>ѻ@?�R?�>�9�|�'���?�޶?֯�?MI>���?s�s?>k�>ox��X/�05��~���`�=�RZ;e�>.\>"���QgF��ד��h��d�j���_�a>E�$=�>�7佸4���D�=�닽iC��\�f�.��>�+q>��I>FT�>�� ?�^�>���>({=�i���߀� �����K?���?.���2n��N�<Z��=)�^��&?�I4?fk[�{�Ͼ�ը>�\?k?�[?d�><��P>��F迿7~��<��<��K>,4�>�H�>�$���FK>��Ծ�4D�bp�>�ϗ>�����?ھ�,���S��EB�>�e!?���>�Ү=�� ?F�#?>Ej>��>jSE�^4��+�E�y��>+��>�V?(�~?g�?=���.X3�����塿w�[��xN>�x?�A?ؕ>ׄ��|z��+2?��I��I��ߓ�?�qg?�1�V	?N)�?}�??V�A?|7f>����4ؾ�������>�,'?/@3���Q���1��=�� (�>�~�>�{�>�����'a�y=<��B�"���f#?��t?��I?�ܾ��V�����Z7=��;�9�==�X�`��>4�>%2�F��=e��=}�>
䄾툽���8�=�>�>�0�=�L������,?���������=�r��7C�7�>
*K>֖���^?�%<���z��q��ty���\�sU�?���?N�?�|����f�y�=?
5�?�?P��>��S�߾\���m�	9q��.��q�=���>���P}�A���7,��c����Ƚ�z��_�>���>�E?�4�>�:>(m�>*����m%���� 	�\�.���I>�@]+�]���ꇾ?��T���缾Ċ���>S�Q�G&�>��?��I>%a>O}�>��|��	�>� T>��t>���>E>M�A>Ь	>�Bv=Z�н�GR?/���)�'����n��� 9B?�ud?�4�>�h��������τ?F��?4t�?TTv>Wxh��'+��o?�9�>���4n
?t]:=vl��[�< U��Ѽ�U"�����5��>�;׽�:��M�Wkf��i
?'-?~*����̾0׽����%���?[�?�	��D+������S���c�S=�=�K����j&�jca� s��˙��ׁ��j9�Ch<��/?�`�?,��,у����Wtp�bG�n�>-!?b�>�M�>��=#� ��ad�<?_��r�390�� ?B̊?O}�>t�I?*<?jP?xL?�܎>&t�>5-��~�>v�;H��>��>4�9?Y�-?�,0?�g?b+?�
c>&�����]�ؾ�?[�?�G?�?�?�Ʌ�;ýqc���h��y�N���8��=q�<�s׽��t��]U=��S>�S?���8�����a2k>��7?m��>��>�W0���)�<��>b�
?V^�>�����or�fW�b�>���?��O�=s�)>i��=�ۄ�I�ٺ�6�={���8�=Ŭ���X;�y�<�:�=��=�Gp��-����:6�;�T�<N`?�?�>�?	�߾�eھ�����4��e�<\Q�=V�=?�߾F���r�8�Z�hF�>Oo�?d��?�kM�)�>�SI�䡁����Y��{;�5��K�!? ؾ>��S?��?c];?{f@?�m->�i�i&m���f��9���,?�!,?���>����ʾ��b�3���?�T?Y;a����r>)�ԕ¾Zսl�>�W/��(~�� ��lD��Z��F��`������?=��?ZcA��6��i������\����C?3�>NW�>k�>x�)���g��$�c5;>}��>�R?�"�>�O?�<{?�[?�hT>М8�1���ә��X3�e�!>I@?��?��?�y?�s�> �>��)�.��U��t�������	W=�	Z>=��>)�>��>/��=��ǽ�^���>�e`�=>�b>��> ��>��>��w>%N�<�}M? �>�Pھ>!侖�ɾ�I<�}b%���?�U?+�7?R��<��Nl.����@��>��?<�?h�'?����݇�=l�(��{!��U�>Z��>��S>X�>�Q>��(>��>~�>ѭ^�H�ھ�@��`��[�>��J?�ӭ=�_���5K��@>q�ľ�(�=�M��j���L��&۾���=�������=J�~��T'�Z��� t��ʂ����%��Z�E<�>���3B>ϙj=y��=��=J=:��	>-���
m>�h�i�K�MO�M�<�	� ��K�=��<�!>�~ǾwLt? hN?=?b�J?��>J>½o�>�̨� {?P8�>���žw'N��ƾ�e���������]���Ⱦ) >�r�l�4>�n>��>��=�9�=���=�݀<:���̛=7C> �>���=Z�3>�>�=>eCt?T�k����]V��)�6"?dJ�>� >*¾��-'?��->�����������?`=�?-��?�4�>��?����>����V��qc<#�
�h��>���=i�g�;w�>���=���������ƿ����?}@�`K?�J���Y̿t�W>r�7>Q/>��R���1�z�\���b�MzZ��!?�A;�K̾�/�>2��=;5߾�uƾ8)/=V�6>��b=:w�~E\��ߙ=� {��;=oSl=��>�C>�V�=x)����=��I=7��=w�O>���#�7�[�,�Y3=���=��b>&>�.�>B3?=�/?w�d?��>�l��;�Q���>��=s�>ﴄ=m�A>J��>�c7?	�D?eIL? ��>�ˌ=mպ>&f�>�=-��}n�1�)ۦ���<9��?�e�?
Һ>�N<]�?�mB��=��Ľ�Y?M!1?�?)f�>0o�F��r��r6F��E >K�@>I��>�󉽴�7=C���N���CR=�Љ>��?�#?R&�>E�_>%��>ղ�>�B�>�->�e=Ig�=.�,��e����Q�=_�c=~�q����:��.h��xʤ��n�;���<�7�<!NҼi��=���>�>���><�=���5�.>�����L����=�'��~+B�d�B<~�i/���6���B>i�X>;僽0*����?4�Y>�G?>���?�u?*Z>�7��~վ�;��.�d��cS���=�~>�<��;��p`���M��OҾ���>��>Q��>��l>�,�� ?�v�w=8⾐Z5�%�>�q��������8q�?������wi���к�D?pE����=�!~?�I?��?(��>�����ؾ�60>�F����=c	��q��w����?	
'?K��>���D��F���0��&��>��ؽ?�T�O���c�M��F��e����?��ȾQ��\<��}��6����4�GC��F��>��Q?��?�災|V����%��=��0;%?�$�?w��>��>qƥ>̫ʾ�J��[B�\�>���?[��?b8�?;.�=�d�=n�%����>"t�>�9�?�"�?��w?����W?���U,�=4/��ήH>%�=�l�=�3<��><��>��>|��q��	6߾X⾣>9��Ա=:|>y�>�W�>�aT>��_=71=�}�>���>o��>9q�>r��>S��>:�q>ل��)5�B^'?3��=ɺ�>�t2?�>��N=
l���F�<��W�_a;���'��8�����U�<�
�u�==�K�����>�Cǿu1�?i�P>4�K=?5��K+��eT>��V>t���x�>�1L>�:�>CU�>���>Uu>�a�>�(>jKӾ�4>���.c!��C�nR��ѾHPz>�Ɯ��%���� 
���MI��K���j�?j��,��1N=�U��<oA�?#���2�k���)�������?!�>M6?�ӌ������>\��>���>�s��w���2���w[���?���?r>c�>�Q?{R&?�pV��/G��MG�5l�6�A���^���c�VԌ�}��i��Y�н�[?��|?nD?����Qr>+r??4��ς�v"t>���Γ<��g�<��>~����55��Už�#ž�-��+>�&l?G΀?�P?�DR�cH\�U�>Ku5?q*(?i�w?��9?�D@?XG��D(?h+#>ڡ?i�?;�<?��3?��?t9>*��=t�<3�!=7���<F��?uʽrmѽ��་�B=ц=��*<�*&�M�=ZQ�<��\�{�<�t����<;�Z=��=�;�=���>�*\?��>�"�>�/?J\&�ؕ/�{���)?�0*=�|��q㏾k⧾e������=��h?�0�?0�Z?�P>m)?��0L�2>�>�2>�k>�o�>B��(�F���|=;�>1�>�=ϱX��넾���T��|kB=.�>m?=9�>;��x��>DT�ubӾ+:�>�#.�h�ʾ���Z�#�(eK��ȾR�`>��4?�t*?��>��Ƅm��@�%b�>`�;?Y�?,�>?s���JF��%H� EG����=�>	���|>���#������%�P�mN7>V{�>i��J���
b>�y��D޾�tn���I���gXK=ay��X=�����վ�!�n��=ߟ	>����W� �k��cѪ�L?J?=6k=gM���8U�6���n�>�k�>J�>��;��#v���@�������=��>��:>�����	iG�#1�|?�>WNE?�T_?�k�?�+��>s���B�/���;h��k&ȼ��?6t�>j?%&B>�	�=���e�=�d�RG���>���>���y�G��6��~*����$�!��><6?У>A�?��R?��
?ǘ`?�*?�@? �>m��������A&?4��?D�=�Խ�T�� 9�UF�F��>��)?�B�x��>'�?��?��&?��Q?�?�>�� ��C@�锕>dY�>��W��b���_>ƬJ?���> =Y?�ԃ?��=>i�5�ꢾ�թ�'X�=�>��2?�5#?)�?��>�,�>�ͤ����=�#�>�+e?ק�?7Dq?>��=��?k�<>)(�>���=j�>F]�>�~?�O?e@t?NH?x��>R��<<䲽c<���R��#�j��s;"�;j�e=����Z�� ��j=��<�ۡ�\�D�l���B�L�s�X�<O��>b�>��վK݀>L��^S��jc=v�꽌���>@������U��H�>�?QX�>������=�x�>�?=��Yd?G?��'?��5��77�w���(Ͼ�)�>[�M?��&>�2N�oHr�u�[�U8�<1�a?&�^?�踾�A�`�b?��]?ah��=���þ��b�Z��j�O?�
?U�G���>��~?w�q?���>��e�V:n�!���Cb�t�j�Ѷ=r�>DX���d��?�>b�7?�N�>��b>�&�=u۾5�w��q��??}�?�?���?�**>_�n�'4���� ?��[8^?^!�>H���u�"?��G�Ͼp[��EՍ��3�q���F�b���wզ��o$�a&���ڽ�=�T?�r?�q?�v_?�� �  d�\*^�ğ���V�����`tE�
&E�H`C��n�b�5���С���PH=^e����?�;ò?PM)?1�K�.��>���������eվ.0H>��{���=��l�p]S=�M=|4j�)�*�� ���^"?4��>�&�>}�7?SGV�x�:�-�3���-��� �N16>x��>D	�>��>tT��2�L5
�D�о�hm���ܽ
7v>�xc?~�K?1�n?Mp��*1�����!��/��b��C�B>�h>���>ɯW����:&��X>�!�r�����w����	��~=��2?�'�>.��>�O�?�?r{	�qi��kix�4�1�飃<�/�>�i?@�>��>	нu� ����>��l?��>��>L���U!��{��ʽ�j�>]ح>���> @o>�>-�a-\�-g��Dr���9�'�=k�h?B����`���>��Q?�ؚ:��H<���>7Qv���!���B'�B>�e?�*�=�V;>O�ž3�`�{��E��n�(?�R?����{�(���q>�� ?L�>�ݝ>᥂?��>ԌľAlU��Q?qV_?��J?ԥ@?KZ�>J�)=&���X�ƽ��)�k�9=m{�>j�U>/Xj=���=���^Ra��]�I�M=�ǻ=<���{���#<��_z<٦=��1>�mۿCK�y�پR���:
�
戾¸���d��"���T���
��fVx����1O'�,V��Cc�������l�l��?r9�?!x���*��ᱚ����O������>P�q�;��﫾��K-������Ƭ�;c!�)�O�"!i��e���'?+�����ǿ谡�]<ܾq  ?X> ?�y??�e�"��8�d� >�c�<Ꜽ���Y���A�ο�����^?���>���)����>��>$�X>�Cq>V����)�<��?<�-?���>�r��ɿ������<���?��@ІL?��8�7!��˖B>�1�>�'�>���=ˊ�~�<��iﾵ��>%�?���?p>i�0��t�4�4?o�m><�C��a�=dS�=%�4�����*mc>&�k=Q@?�p�=iw��(%��,J�>kl�>&����Խ9u��5o�kX*>@�p��G��Ԅ?s\�5f�#�/�Q���s>��T?�3�>�E�=��,?*4H��{Ͽ��\�O)a?.�?T��?5�(?r迾�ؚ>��ܾ|�M?uC6?���>fc&�^�t�!��=d"�䇧����eV�{��=��>�P>ƃ,�����PO����7��=,;��nҿ�_��t��V8�=α�=�T����K6ʻ�Q=a%��:�]A���O<N
�=��>�Ȯ>�r->�yD>(�Y?E�?8m�>0�+>�
��|��+�߾�y��&ͨ�A���e��,�Gt���w�,7�D;�h�(�n���/羌=��K�=[*R�G���.� ��b���F�N�.?��$>��ʾ�M��-<�ʾѪ�hz������^̾��1��n�"͟?��A?������V�;�����-���l�W?�"�>�����`�=
����q=�K�>I0�=���3�dyS�e).?z+?ilɾ�4��1�=z����^8?]��>�{��5�>Np?h���p���ˀ>0�!>��>�\�>�e>�R�����z?M�c?���ɠ��1�>����r�����=��%>Q�����<o�8>�5�<W>����������G�<�kW?#�>	*�H*�xK��"�#��%A=�[x?��?�A�>VBk?�AD?���<�q� ]S�����Ao= YX?��g?�>}���оTƨ��~6?��d?!�Q>��d�ܜ��/��|���?��m?�n?�	�� }��Β�r�~�5?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�ٕ��Z�?��?~���|Dg<R���l��n��o�<�Ϋ=���E"������7���ƾ��
�����࿼ͥ�>EZ@�U�v*�>�C8�]6�TϿ)���[оSq���?M��>Q�Ƚ����A�j��Pu�b�G�2�H�ť���p>��>����/%��dw_�:�k��o��O�>+�>�6�>�;����������m�,Q>cX??6�ѽ-����?�+���sۿ�o��˾���?��?�5?C`?lS��'��-i���h=˫|?�?5��?�S�=KS�� �O�%�j?�_��xU`��4�uHE��U>�"3?�B�>T�-�Y�|=�>���>g>�#/�w�Ŀ�ٶ�=���Z��?��?�o���>r��?us+?�i�8���[����*���+��<A?�2>���H�!�C0=�TҒ�¼
?V~0?{�f.��D?����Ev���f��$S�Y��>�Ѿ'�־��=kvc�R���0����`����?���?ze�?TA�<d ��n>?H�>t���0��f�>JP�=�ҫ>�^>������3�P�"�o��>�Y>��?�D�?�k?�7��C���r��>���?�>3�??��=�_�>���=�簾�'��~#>���=֦>�?p�M?S�>I��=�9��/��\F��ER�� ���C���>��a?JzL?�eb>KƸ� �1��� � �ͽMA1���0@��,�8�߽	5>}�=>;�>�E�wӾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�v		?4��F��]X~�ρ�ۄ7��)�=��7?��{>���>]�=�tv�����l�s�\��>QD�?5q�?���>��l?ho�hC���0=�R�>m�k?�d?��t����:BB>{�?�������84�m1f?�
@�u@`�^?�碿�hֿ����_N��N�����=���=׆2>�ٽ-_�=��7=��8�[=�����=s�>��d>#q>>(O>�a;>��)>���P�!�r��\���R�C�������Z�B��Xv�Xz��3�������?���3ýy���Q�2&�#?`���=˫U?�R?:p?D� ?�wx���>����L=$|#��ф=�,�>/f2?n�L?��*?Vԓ=�����d�C`��iD��~̇�h��>�qI>�~�>L�>%�>A�B9O�I>S1?>%��>� >Uq'=�,亮c=��N>�M�>���>y�>�C<>��>Fϴ��1��k�h��
w�r̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��x�T�4:>9����j�6`>�+ �~l���)��%Q>wl?�f>	%u>N�3�d8��P�r��lm|>�36?ᶾpB9�F�u���H��aݾHM>[ƾ>�FC��e�E���$
�P�i���{=�x:?��?�?���䰾ßu��F���BR>�E\>)�=�n�=�KM>��c�d�ƽ�H�#�.=Ӫ�=��^>��>})>1�1=p��>�FѾ<�Z��>.<<З�=C%?�7?�Oܽ�E,���0�	����>��>��>��T>_
p��'i=+�?�xB>�{ǽ���&T��R6���S>�wx�fLS�c���ͻ�=�Gn����=�@"=�S,�����v�;%�s?��h{�cL��(����7?"˼>����
%�!��Mƛ��������?Se@��?�����E�8`/?���?ly�<$� ���>��>�&�'m!�
H�>t>���Ș��ӥ��:�?��?�H̽N4���{�O�N=��)?� ��j�>���ZY��
���u���#=���>O5H?�]����O��>��x
?�?�W����0�ȿ�zv����>��?x��?��m�A���@���>Z��?�hY?��i>ye۾]mZ�t��>��@?+R?��>�;���'�W�?�ݶ?2��?HI>���?�s?�k�>,0x��Z/��6��򖌿kq=�[;�d�>}W>}���|gF��ד��h��m�j������a>͗$=�>�D�P4��z9�=���H��ںf�0��>-q>I�I>W�>i� ?�a�>f��>�w=[o��hှ����B�K?��?��N2n��n�<�͜=h�^�c)?�G4?�Z[�M�ϾDɨ>�\?���?�[?�h�>B���>��o俿D�����<��K>�7�>A�>�4��qWK>��ԾBD�`w�>֗>�磼\Cھ�;��,ţ��@�>�k!?u��>p��=ՙ ?f�#?��j>{+�>�aE��8����E���>_��>�G?h�~?�?.Ϲ��X3�����桿�[�BN>C�x?�V?�Ǖ>F���t���h�D��FI��#��?�sg?�a�?�2�?�??��A?#f>L���ؾ����?�>��!?��w�A��;&�SI��v?�B?���>b���5�ս�׼R���]���?�+\?i=&?Ў��a���¾���<�#�V�N�� <xPF���>��>�����O�=H>'�=�Dm��$6��0f<�q�=,r�>^��=�7����s�+?�8�	���=�=��q���C���>�XL>H޿���]?Z�<�h|�Pି~P���fU�溍?�L�?<�?`���-$i���<?'^�?#�?�V�>����޾ٳ߾�r�_7x������>y�>����?�#.��@���Wǃ��V����&��z#?��>�6?��?O->&[�>�5:�{��+�ž��hT`�r9*�,AF��4��_�⬦����?�]�j��4�b�؟�>ї��D�>��>j`>>k>X��>���=�ȅ>!e>\6>XG\>�m�=�$�=iѼ����@Խ\�q?C���2M���������w(?�8?�+7?n\������4��+L?���?ך�?mө>=%��� +��D?3�>a�>�>�U۽}=t��ר�ᝡ;)'g��=w]>b$�>d,a���{���L�񸣽Q�?�u(?�ߚ<M���P>k���㼉6�?��?J����_�1�\���>��<o��0�>w����P�~)�Po�dz��Hfs�0E���W0����۝M?�{?$��ïɾǰ⾜U��1�U��Hx>��>��>�M�>�@>�q(�4�0�t�f�p?�Q$)���?K׀?���>�wI?J�;? ~P?�*L?>�9�>Qd��5&�>� �;���>ʷ�>��9?��-?�00?�j?vo+?8sc>����	��~ؾ�?H�?�?��?
�?�䅾�ý���Cg��y�EV��4=��<�׽]v�2�T=��S>�3?
��1�8��|����g>ǋ4?���>;��>쌓��=�����<���>�a?�l�>�����r�������>v��?�����<�b'>'��=�a�PA�:��==���� �=;��EH��$<4��=`��=(������}OC���;"J�<G�>�?2��>�F�>���֤ ����Fΰ=7�Y>��R>��>�qپi|��X!��J�g�gy>�d�?Qg�?ܒf=6��=���=0���iE��	������-�<Y�?�Q#?�RT?Ԁ�?~�=?w>#?tQ>i/�:?���_���0���?T,?%��>��,�ʾh騿�o3��4?%?�=a��+�
S)��v¾�ӽ>x>�/��~�گ���C�E	�I��?����~�?:۝?�B���6�q.�ؠ��M䬾�|C? U�>�m�>y�>$�)�^�g�E��:>���>Y�Q?�L�>�B?.gn?>/b?Å�=��2�"����o������,>0�2?uJr?d�?v�z?��>�>��	���ľ�$׾v�ؼ�%�%�n�}�N=�K\>�f�>��>�&�>y��=0��ʶ���E��a>V>�?�>���>z?�>,n�>(����G?	��>�`��З�F菉�Ã��==���u?��?��+?} =�����E�G?���M�>Gn�?���?�2*?ϧS���=
�ּ�޶���q�%!�>tֹ>'/�>�˓=�-F=�`>7�>���>��.`��o8��M���?�F?��=�"ͿMV���^=}9d��6e=�T���]�.�$��Ph��%e>���函d����I���;Ծ�����I�|F�c־n�#?W9�=;>�<�=l<��Z����kP>��ǽ���=�\O��d<<a��a�;=�νC&��:҈�Nl�<Ӑ���۾��?<�d?��?&j?�l~>�H?�>��?��=�?Ż5<ӗ����EԾ����X�[����
��վXB���>B�D��T�>���>�%>P�^���><U�=m�V>�h�=l$>_Lv=��w=~e�=���=�䚻�H�0�m?NYm��Ś�rD[������-?�fe>,�3=N;��=�9?�4�=�k��F~���+�
�z?H��?j��?/f�>@(g�D��>�V��6��'�M<����Ȣ�>�u�=�\����>���=��X����$�P��?
�@xX<?|����YʿkHR>S�7>��>�R��w1��\�<�b��jZ�S�!?�K;�<e̾�:�>gû=� ߾�rƾe�.=A6>b=��>P\���={�z�D�;=�ck=��>9�C>�غ=�ԯ��-�=��H=��=�O>�Ŗ��K7��,�8F3=5��=<�b>�&>\��>��?�I0?8hd?M��>Xn�J*Ͼ�����>y��=3�>�x�=[�B>���>�8?r�D?��K?���>���=u�>PϦ>��,�4�m��8�����w�<^��?���?���>�R<�"A�fp��V>�xŽ�G?&1?s?ꠞ>�w��ῠ %��U.��	�����;eb2=j�q���G�T�༄���:�Φ�=�K�>Ƣ�>�.�>�}>��8>R�N>p�>��>,�<�Y�=�K�����<����=����i"�<�������}��$8���ʼ��}:ew:�=<.c;�^�=s��>��>JX�>��=����@>1���sF����=S��2D�M�c��$}��{-���-�7I>�`>I���>���w�?/y>�*9>!:�?�l?��>���Y�þ�����vw�GM�~��=���=�&S��8�+a��H��Ǿ���>�ގ>-�>E�l>N,�G"?���w=���b5�E�>�}�����!��6q��=�������i��-Ϻ��D?F��8��=�!~?��I?���?ڋ�>� ��}�ؾ;0>E��o�=p�c&q��m����?p'?ȕ�>�쾆�D�>�پ�_a���>c�.�*K�ר��r<���)=������ ?���B���-D��≿ 4����3�fk���>�k<?ㄪ?�N�����41I����<�Jg�>��k?�f?w��>}
�>#cݽ�򾮏]�F>��|?��?g^�?�� >�ň=���;�>XT?t˘?ձ�?�w?^)�6[�>�d=u$W>�}m����=���={�=��=�j?��?�� ?t�����	�Q���h�wG]����<'Պ=T&�>!҂>��>�>%C�=)ů=]$]>F�>�:�>�^>K6�>�j�>����[��&?� �=hr�>�a1?wz�>��4=���Hs�<�9O��2@�H$�0׭�V�սTJ�<ZT"�:_=������>u+ǿ�z�?+�R>��?/������lO>!�R>�ܽ�"�>��J>�{>Y��>E�>͞>��>��">�^Ӿ�G>y��T!��#C��wR�p�Ѿ�Wz>����%����q0��D/I��o���i�^j�e.���<=�ç�<L�?�����k���)�,��Vv?�;�>"6?8��授�k�>���>2��>]@������vÍ��o�
�?B��?�0c>#�>��W?��?��1�}Z3��wZ��u�=A�`�d���`�5܍�ԗ��N�
�����_?j�x?�tA?��<�Nz>b��?m�%�uۏ�a(�>�/�*';��A<=;*�>?���$a�!�Ӿ֥þh��}F>��o?�#�?sS?lcV�P��|�=�H?�g)?f�?aA?��K?[ ���1?݆>zD-?�5?�?�
?��>ʧ[>%�H>� �jy-�����*�� �6��8-�="��<�����ɻ9��=k�=ݝ=#J�;mC�<
Dj<�|�<��,=��=<��=~@�>xW?���>V>�"?S�"��TA�n����?��A<]Ò��Ά�z���@Z;��1>�]?��?�W?p9�>s#7�f�f��u*>��>�>&p9>��>[���z�/��='�1>�h$>V�>�����r���[U���(�=yo>N�?E��>Dfl��v>�}d��
�����>��X阾�(��#�_>E���z�玐>$tB?�]?S��>O�㾆;߽�ֈ��-?�4M?_S?3T?�-�r9J�tn8��-�v'�,�>dպ<t����r����&��<��>�\��ކ�i�:>���7����o��;T��	�%<�;s�
���=����>��s�|�=`>!˩���*�1�������-G?V��=�h��4�i�*ٔ�7�C>>��>Q�>�(���4��PA�}T��{8I=���>�-(>�s�<"�쾥C��$���>/nD?�x^?su�?�#���ns�� C��
����U��Pn?n��>�?�>>nT�=�������JOe���E���>D�>��x�H�|J���^��sH%�DG�>��?/l$>)�?�AR?��	?t�_?��*? �?�ȍ>�������B&?3��?��=��Խ�T�� 9�IF�}��>y�)?�B�๗>R�?�?��&?�Q?�?q�>�� ��C@��>�Y�>��W��b��K�_>��J?ۚ�>p=Y?�ԃ?s�=>[�5��颾�֩��U�=�>��2? 6#?L�?�>��>Ί�a��=<��>�4d?���?@|u?�H(>ё?��H>��>�	Y=݅�>iv�>u=?ZJB?" m?+�Q?|��>ix�<�<���˷�^����}�ڽ��<Qǈ=�~$���`�ґ��A=�z�<��9�t�T����:��ʒ���&<w�>lJ�>Ԡ�����>����h���f��vb����Q=��8��6S�L5�>���>]��>���1V>d}�>��>�.�9�^?@�?Ar�>Ein<�~4�-����f�P �>1�
?�ۯ<X5���o��?�o�Ix>#,�?7a<?���1撾Ic?�\?�G����=���ľX�h�sh�IN?VX
?��@��O�>&&?mq?v��>M�c���l�~=���b�8ii���=	��>B�e�Fj�>�7?��>I�a>GC�=��۾A�w�9��H�?��?F^�?X �?��'> Fn���߿R
�:���d?�W�>��P
?Ž�<��Ⱦ	�o�v�����֣��~��M���񇓾ca&�?���&����=�b?�u?w?��W?�\��ha�ՖP�y��"�M�� ��+��@��[@���9�#�r������q���Ji��LJ��w-A�_I�?��%?0����>�������ɾ.E>P������_"�=X���-�:=G9H=�%q�]42�kf��gU ?w'�>���>>�:?��\�Kc>���1��Q7�����E
4>�P�>䇑>sP�>J��<J.����ʾ�����)нr7v>�xc?Z�K?��n?�o�+1�����+�!�B�/��c��I�B>,j>��>��W���c:&�mY>�(�r�d��w��@�	�ƣ~=]�2?�(�>g��>�O�?�?�{	�[k���kx�!�1�M��<=1�>� i?�@�>��>н(� ����>6�l?&��>�i�>a���`!���{�l�ɽ��>䍭>�N�>o>��,��<\��a��X���9��F�="�h?/�����`���>}�Q?�:yG<ۙ�>��t���!�Z���'�HZ>�c?�B�=�;>��ž]H���{��?���\!?wR?l����3� ��>n�%?I�>��>�.�?Q��>+������DG?o1X?�L?�8?�b�>ڕ�=~L����>�)�� =$Ɂ>,�J>v(C=��=�E��RX���ʊ2=���=LN�����W�;��ؼ�<|m= �.>�Jۿ=K�pؾ���\��	�����>��Cņ�U�7������c=z�6��_�&���V�0�e��㌾�El��T�?�?����-A��l�����N���RB�>/�p�*���ʫ�
������������Ue!���O���h��he�`�'?������ǿ氡�\;ܾ?  ?gA ?'�y?����"���8�� >uI�<������I�����ο�����^?���>B�4�����>צ�>�X>eHq>���qꞾ[�<��?Ƈ-?!��>��r�&�ɿD����Ϥ<���?��@��d?Gj���;X�Td�=𧖽8�k>��ӽ_��� |W��ĳ�V�R?3i�?
+�?
l�>�����>l�W?j׾q�q��$�{��=;�>JI�>�}.��l�>H�=F�>�d���B<%�2>%�n=j�K>�))�@G�Ң���5�>�(�MSK�5Մ?,{\��f���/��T��U>��T?�*�>R:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=r6�܉��{���&V�{��=Z��>b�>Â,������O��I��T��=����Jÿ�n�,��@z�=ն�=8	�;O�@�713���.�ʽ����Q���@�CK�=A�f>�|p>��@>�_>W�>I�N?"of?y�?�9>�ֽh���m��P��7�~��.�3��n�������Ѿ������!?�;�-��b��`{4�rPL= pR��Ñ�|�#�3�h�ïI���%?��!>�㲾�C���=�iǾ�~���-�!n��D�־�84���g�3F�?��>?UP����Y�"��M���F�i��U?`,���-�����=�2��q)=���>���=�澨�0�4]S���0?�?����g���d'>�����v=HO,?�t�>�(<|��>�j%?�O$��Qݽ]WQ>��6>A�>0��>�(>T�����ؽNn?=U?N��睾I:�>�]��y�{���y=n3>c6���̼GNX>>��<+k��e�9��	����<��W?���>Ć*��;�e%����2�{==3Zv?|�?�:�>ٍk?NiC?�9�<��r�R��0	�a[=�zU?Bh?�	>�w��4о�����6?}�f?d1S>^i�K��ߵ.�{R��?l�m?��?�����{��W��Yt��W5?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������u��=�ٕ��Z�?t�?�����>g<B���l�en�����<�Ϋ=���F"�����7���ƾ��
�����߿�ϥ�>2Z@�T�5*�>bD8�R6�TϿ���[о�Rq�u�?E��>�Ƚ��&�j��Pu�e�G��H�����z�>�I3<u��*�Ҿ����Od��q�:�>Ъ�<m��>�Y����M�t0��dy὎|�>IW�>��=uS+��b_�J�?�;پ�ѿ�r��N���A?���?�]?Z��>ݩ��\�����������V?/l?�^?[��)�$���_�#�j?�_��yU`���4��HE��U>�"3?�B�>\�-���|=T>���>�g>�#/�u�Ŀwٶ�����<��?ȉ�?�o����>i��?us+?�i�8���[����*��8+��<A?T2>ǌ��3�!�S0=�Ғ���
?5~0?�z�>.���M?ލJ�m�J�3�'������/> �x����LJ�V��Lz��E����� v�?��?��?0�X��k��0C?�S�>�X���%*����<�9�>*�3>�O>��<OfJ�@/��d%����>� �?�@���>�Ǒ�y������>�y~?s$�>��?�n�=b�>�c�=F�� -��k#>�!�=��>��?��M?$L�>�W�=��8��/�![F��GR�h$�<�C�"�>��a?�L?8Kb>���i 2��!��uͽEc1� T鼏W@���,�מ߽x(5>��=>�>�D��Ӿ��?Dp�3�ؿ�i��up'�Y54?��>�?4����t�V���;_?�z�>�6��+���%���B�a��?�G�?B�?��׾�V̼>H�>�I�>��Խ���{���^�7>f�B?���D��h�o��>���?
�@�ծ?�i��	?���P��Qa~����7�(��=��7?�0�#�z>���>��=�nv�ݻ��S�s����>�B�?�{�?��>%�l?��o�T�B���1=M�>ǜk?�s?Zo���l�B>��?%�������K��f?�
@~u@c�^?$�ֿwl��� ���T�l1>�;�>�h>�y2�[Q>��=͠��������=jg�>��>\5�>ػc>
ؘ>��>���ƀ'�����\ׅ���#��e�	n��.Y����,���� ��������7B��*���<�޹�U���z=���=��U?{R?�p?�� ?M�x��>9����E=��#��Ȅ=�-�>�g2?ڦL?բ*?�ϓ=ߨ����d�a`���A��ʇ�k��>\pI>��>�J�>+%�>�O9S�I>f2?>Q��>" >ih'=FK�lg=�N>�M�>t��>�|�>,�>>> ���yb��O�h��z��̽��?]���'�H�?v��mI��О����=�(.?��>xT���1п�{����G?ʧ��1M���+�ړ>��1?=�W?��>�����X���>%W�ׇj��� >/<��h�4)�#�O>�?��f>��t>|�3�m8��P������t|>6?]���d�8�T�u��H�aSݾ6'M>%��>��@��n��������ii���{=�p:?��?հ��?�����u��C���R>�\>W=)��=�kM>^oc���ƽ�H��-/= ��=��^>�?�?	>��<���>o�þ�,��a�|>�W{<p>`ZP?P�0?GŲ=h��<����bP�w�>�>g�>��>l�:����<��?s>H/��Q�s�>�bs���E�>�X�=όM�8WC�m��<�s����D>�h=��[��^I�� >��s?����у�9[ྉM���?r)�>%��;+?��y�'�����&��}l�?��@Ҍ�?��U%\��W9?�_�?�hT<�h�=1>��>2[���#��IB?9�=�N�(��V�=|��?�Q�?p�<I���y��M^>��?����>����w��͚��E@w��
��A�>N^B?9|���Ś�� L�	?�b?��Ѿ�-�� �ǿ�Fu��D�>"�?x�?Ck�ն����5����>> �?0X?i�>?c��|�F��>�'J?�T?Cg�>�C$��H4�	r?���?�+w?0I>t��?��s?�r�>Ǘx��]/��5�����pw=��d;(m�>rq>տ��HiF�֓��e����j������a>բ$=	�>@�yD���,�=
���P��h�f����>Fq>��I>�U�>�� ?�Z�>q��>*z=ʲ��#〾3�����K?��?���\3n�hD�<���=�^��%?�H4?�-[���Ͼ�֨>_�\?���?4[?�e�>���a>���翿�}�����<��K>�4�>�I�>h��kFK>��Ծ�7D��o�>�ϗ>b룼�>ھL-��ۃ��YB�>�e!?d��>Ү=��%?� ?�D>��>L:[�R�����_�Pk�=(Q�>��B?[��?ww0?+k��X?��#���Ԍ��>V�hE9=Pe{?d�?�
>�R��ߐ��Am5<=�0�"�G �?#2Y?��N
?Fl?��?;+-?���>�5��H�Z����w>�%?d�BXE���.�u�����>Ս?�u�>���7J�tl;V��*����#?��V?�,?q~��Je��ν���<��;������<�F=[�U>��)>�n��+�5=%�>�V�=9T�X�'�R�;甑=���>7�=%.�ꚽd+?�ߺ'i���V�=�;q�Z�C�3�~>��J>�����\?��@��}�����Lg��)hS�K�?�/�?�}�?hK���h���<?�>�?�\?���>@����nܾ�cݾ�	p�΀v����=�>���>�=��dc辙���U��������ɽS�.��U[?��>�:?�?Z��=d��>���M������#���|�A)�H�]��?$�/>��.���2*޽p�ɾqd�����>���&�?y?S?�>	6�>�M�>P����d>�6y>���=�`�>���=���<o��A����9�7yR?���xy(�T6�������{3?�G?���>��0���|�g�A^?�٘?N,�? Ƃ>CFz�&H���? ��>8X���O(?�3;I@=�H)��j(¾2���a�rCV>�v��k$A��5=�⍾S�?c�?lě���f����=�'��W��<yI�?(?w�!�:9F��TV���L���5��(�����L��8:���i�۞���酿b��0$(�� S=vI1?���?�,վB�ܾz����l�T!O���G>@��>�T�>�_�>U>ъ	��4�2T�LP�ZNP�Zg�>�1o?R��>;�I?�<?xP?3kL?h��>�b�>N3��6k�>���;���> �>.�9?i�-?D80?�z?mu+?E7c>f{�����K�ؾ�?��?
K?`?��?�܅��ký�a���g�U�y��d�=���<��׽�Iu��T=aT>�p?�����8�E���>Ik>_�7?<��>�>-:���K���$�<|��>��
?�y�>>	 �X]r������>�^�?+��}�=�)>J��=�����g�4Y�=�Xü�T�=bW��J(?��b<��=XO�=r�i��\ۺu;���;q��<��>�� ?MΊ>��>k���� �����_�=޵V>l�M>�9>�3ݾ�D��D'��x�f�G�u>�1�?Ka�?�h=֟�=���=�	��10��>��m��ǽ�<�?J�#?'8S?���?S>?|l!?���=������ ��������7?�6,?w<�>����ʾoਿL�3�s?9?�=a�}f��(������ ԽL�>�N/�m�}����4D�#ዻ������#v�?)��?Z�>��p6��X辶���Cv��~C?��>T��>x�>��)�{�g�#���;>Ȇ�>��Q?"�>`�N?-z?Vc[?"�M>�}9�;��Uw���v �M/*>��@?� �?Q�?�w?���>��>n�*�b��\r�����A	��Q]��`/=[�X>q׏>��>0�>-��=���Ĥ����>�H�=��`>M��>X�>D��>��u>8��<�H?o>�>�ݿ�?���줾ヾ|t=���t?0I�?��+?V�=��N�E� ���J��>�x�?���?p�)?؄S����=��Լ-���mp�*ָ>غ>�Ƙ>�G�=a�@=��>���>���>�E�
L��q8���L��D?y�E?K��=M/��;�c���9>�/��{�>iy4�R]=��G�N����Z�=8�˾�8��k�Թ�^#������X�#�.d��\,���?��5>���=\Ub�=.-��Ǹ�4�}<q�<R��<b7��*Id�����/�@��Խ�m�&������1��"����׾���?�N?��G?nBx?9 �>X�>�!>�H�>�n,�T�>ñ��9�h�����7�l��ĥ����ؾ�̾�~t�Y����=��$��2Z>�>}�K=�˾:��>nK9>'�,>�k�=�L�=9�2>va<>��=�>%�>~\k>�6w?W���
����4Q��Z罣�:?�8�>R{�=��ƾq@?w�>>�2������yb��-?���?�T�?>�?;ti��d�>M���㎽�q�=S����=2>r��={�2�O��>��J>���K��+����4�?��@��??�ዿ΢Ͽ<a/>~�f>=��=��W���8�o�g�Pm�ZV��O?�;��Ǧ��B�>39>��о]�Ⱦ��<��w>&�V<G�U��TU��P�=�S)�_p`=N�=��>��>��=PW���	�<t��<���=�hV>��t<��m�H��,�E=��>+^>��>��>��?L@0?}Wd?Թ>�gn�LSϾҠ��t+�>9D�= U�>ڞ�=��B>:K�>_�7?��D?.�K?�H�>���=�>�>�k,��m�S�X��5�<ㅈ?�̆?s�>i�S<��A�S���`>��6Ľ�p?%1?bV?���>h�	� �ؿW�쾏r0�XAt=��I>�>�)����=��<�#&�yX�\�����>1o?Je�>���>)��>�)�>���>���=�^�=���==���q?�	}�=�P �i��=�线��=�h���4��@����<h����#�TG=d_�=��>f�>'�>v۠=����e,>�/���~I�{\�=H����E���c����W-���=�iEG>[<i>���Hܐ��?��i>��C>�n�?έm?�%>#���C]ʾ�훿Ǿe�>�ϰ�=d1�=�eR���=�^�b��rL�΋Ҿ���>1ӎ>��>U�l>�,�I(?�c\w=�3�U^5��)�>�^�����<��9q��;��^퟿pi����D?�@���X�=�!~?��I?�ڏ?#s�>7N���ؾ�h0>�#��b�=V �n1q�Z����?	'?Hv�>�쾟�D�b_о��z
?�8x�	Z�����4����$�O��>�a˾^uܾ�OV�L􃿨E��+t=�~W�����>J�??�6�?G���Vw��k��}Q�:��8�>� ?�@�>ɬ?���>��O��料��P�z>%@�?��?���?�D?>�N��@�>��?ձ8>�k�?-��?��?��7>�gY?9�=v(O<�|�C�½f!=���>D�_�A��>��?`?u�O�� �t�žA��kQ��z�=z>�<�>��>�$�>�n�=:�>�=�A�>`�>R�>�΄>#�>态>0c���w���&?$�=#͍>�72?���>�,Y=����e��<��I��/?�{G+��d��s���.�<�����~P=߂˼	$�>R�ǿB-�?#�S>Μ���?�N��]�0���S>�bU>��޽��>��E>�3}>y�>{�>7>�w�>�4(>IXӾ	>>;���k!��C�jrR���ѾYAz>�w����%�I�����տI�Yn���^�Mj��7���;=�y�<NF�?����l�k���)�(7���v?��>�6?+��9����>_��>,��>^������-����h���?���?�`>��>y�X?��?k8�i�6�S�Z��yu�y�>�PVc���`��č�<쁿��
��ҽ�w�^?Z�w?�tA?�9�<L�>)�?4�&��\��?9�>�.�Nc:�a�=���>^T��/lf�.վ�X�����rP>��p?�F�?�?v�Q��e��f0>d+;?v)?(�u?D)4?H�??�I���*?L9>H1?5?��/?��+?*u?G�(>� �=��<ڨU=����G����ɽ�Pڽ*=/��~$=�ee=%�;I���(=���<����f4ռ"��;��B�<q�<�:F=|�=?1�=]�>0�f?���>��>�C4?���1��b�(?��<� ���e��;���4�����>)�`?۩?p�]?}d>��K���,���=>O�>�?>ע/>��>����A�T>�=�)>�%/>}W='}��V@��Ϡ��F��<^�<�2>ޝ�>���>��g�r>vB���}E���+> �I���Ǿ�����I�o�Q�3x�̪�>0�M?��?��E>���q�弱�]�ݕ5?2nP?�>M?��z?��J������������ݽ���>/]s�D2�Ą�U��df>��~���>�ߴ�TƠ��b>��kg޾Ιn�J�K���L=Tr���W=h ���վ�
��%�=y4
>����[� ����5Ū�1J?҉j=���ȌU��X���>Y˘>��>�[;�X�v��~@����u�=��>I;>��������oG��/��d�>�C?H]?R��?�����t��JC�b~������ԫ���@?*֪>Ա
?��M>s��=< ��e��a�`�;E��3�>�N�>�c�,BE��ݞ�I��j?%�jQ�>��?�>�i?CW?�?6�`?�(?1�?��>�ε�X����F&?ix�?Ԅ=�wԽ{'U��9��4F�#��>�w)?~B�P�>a�?Q�?8�&?X�Q?��?o>�� �&@���>=E�>X�W�Gb��o9`>��J?E��>�NY?�?�=>{5�q��Ge��d)�= L>��2?�#?��?˝�>8�>㕡���o=t�>f�b?�܃?Ҍo?���=>�?�n3>���>̉�=9��>L��>+c?l)O?��r?1�I?��>���<����n����t� I�q�;*;<��{=)�����/��:�<��<������Rs� L8��T����
<���>B��>-��j�>�Dg��G�����=��M=h�߾)@� ���7�hb�>�7?�	?�@�kL�>�>R�>Q�M���R?�?z
W>Җ:%
;�<5��˨���>��	?P[*�G
�����bZe��v�>�{?h$?�GZ�e>��b?ߧ]?&E�F�<�+Nľ�Wc��&�ƲO?Ѷ
?��E����>��~?��q?���>!e�'�m�R���?b���i�R��=K:�>���
e�؛�>��7?=��>{�c>��=.S۾��w�0Р�׿?�ӌ?S�?��?�[)>�n��'��א���a?wȡ>�C��r?mjx=�ʾ�X��{���T�7����������@Z����A�Z���P���;S�=�"?y�w?HSa?0&Y?d8���d�{�Y�ݵv�!f]������F���4�W
5�ROd�S��0{Ͼ����� �=]�b+3�M4�?���>����u�>�7m����i.�ZY�=��ؾ ����
�=��>���<�1i=E�[�fٖ=�D7��@A?�R?Ҽ"�P?a�|���N�R|���۴R��7L�`�>ux�>��O?�>�7�<e,��-l�������^v>�bc?�yK?��n? ���21������!��k/����nC>��>t��>��W��h�b!&�[>�� s����K}����	��A=�2?�>z�>�H�?��?�e	�&`���Cx�a�1��S�<�"�>�i?Z�>���>"н�� ���>Ҽl?���>O�>�����[!��{���ʽ�"�>a�>���>7p>4�,�m#\��f���~���9�/�=�h?������`�c�>�R?��w:=�E<�~�>�v���!����w�'�U�>�|?���=ܱ;>\�ž��*�{�6��=�)?�}?s���B�*��j~>��#? ��>��>ho�?6Ɯ>�����&�:\'?�:]?r}I?�DA?���>c=�̫���ɽ�h'���*=uņ>�f\>�Nw=���=���	z\���#�aF=S2�=�)���1���"�;}(�����<�e�<w�4>C�ڿ��I��þW6�d侉���%t���T�i�7�
�e���<��Q
��?�����]��q�L0��f#k��:�?.@�?:��y,���%��.O��<���\>�>�������笾B�����ھiʬ��6���O�Lf�Ǧd�;�'?i���Y�ǿ����q-ܾi5 ?�@ ?N�y?��Tw"��p8�8� >���<T���v�l�����ο����Q�^?���>��	{��n��>���>BY>�q>i[���ើ�A�<Z�?��-?��>�ir��ɿ}���f�<e��?��@(�I?Ҁ��8�S�b�=�½o�>��u�.˼�;A��XǾ��4?>F�?u��?���>���ѽ�>.�A?bMϾm�2���"�&8�=�UE��B�>�ܽ��=�;��M�=%s�=ߍ2>rr.><��>@�C��I=�_9 ���=&�>c���2��4Մ?#{\��f���/��T��=U>��T?�*�>:�=��,?L7H�Y}Ͽ �\��*a?�0�?��?!�(?Aۿ��ؚ>��ܾ��M?aD6?���>�d&�"�t�ƅ�=j4�W���o���&V�M��=W��>��>ς,�ۋ���O�qJ��-��=� �?(�����x��e>%b=uu�<蠼r��=���{s��Z��fX;��{�=�,E>�l,>4�X>45�>��H>��M?�ty?("�>�E>�w�[(ľE����uݽ퀅��~�������ӽ3���R`�uZ���u;C��!��E��*<�%]�=
�Q�����3!�t�c��F��0.?*�>j+̾'zM�~�1<�Tƾ[6��N�i�U���̾4@/��!m��ޟ?tA?}����lU����|N��޿��mV?a���6O����>.��V�"=5}�>9p�=*�ྙ�2��$T�[}2?�"?�uɾ� �����=���v�+�y�?K��>n��=�U�>@1?�G�����bK>�7q>��>�j�>2WB>�����ý��?�h?�J��X��ܘ>x�����O����=�C�=șS��
�-m/>LV�=[X��H���ν�p�<wr^?�e>�q5�I��/�����=�X�=1^?��>;�>��k?K�:?�uo<�P�8� ⾯d ��F<?[�a?�#!>G����ᾌ���GOR?�}?b��>����u�n�:����h�?�V?�f?I�����j�ϼz�x��T�)?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������*��=�ٕ�wY�?��?����*f<���gl��q��MS�<���=�:��#"�~�� �7���ƾ+�
��������M��>RY@Q�轚/�>�P8�@5�`UϿ����hо�`q�	�?S��>TȽ����i�j��Mu�۰G���H�����|�>k.|<I6&�)bn�����6�ۅ��`��>$�+�l�>81>=k8�w���>��]��>�>d����N۽`*�D�?�qԾ�^ҿ����y+A��3�?�p�?t�X?�?�>fe��XP������4?^=?��D?$.ż��&��@0���j?�٪��`���4���D�H�W>��2?d��>�.�7�=�>���>�>�X.��=Ŀ�g����?�>�?���i��>9a�?j�+?Վ��G��
��t�(��El�SA?1�1>������ ���;�*<��ޯ	?��0?������_?ܚa���p�y�-��ƽ�١>��0�9e\�y`��Ҥ��Xe����[>y����?�]�?'�?����"�d6%?�>l����:Ǿ7�<��>�'�>&N>�I_��u>	���:��m	>��?�~�?Yj?ԕ������IW>G�}?���>_��?���=~��>ul�=�9���;\�ȥ>jt�=S,���?��M?&M�>I�=��6�Q.��SF�7�R���M�C�;)�>G�a?��L? s`>�D��+�/��_!���ɽ��1���޼�A��?!���޽�B5>�S;>p>S�D���Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6��+���%���B�_��?�G�?>�?��׾�R̼�>>�>�I�>=�Խ����\�����7>1�B?U��D��t�o�w�>���?
�@�ծ?ii��	?���P��Va~����7�e��=��7?�0� �z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=9M�>Μk?�s?�Qo���g�B>��?"������L��f?�
@u@a�^?*Mܿ����������h�>���=�F>�if���>���<��F�!-����=�̛>�k�>��>w-t>ah>jX>����Y�@�����ut6�r��y*�3V�\�cN��1�
�ɨ���ƾ����uĽ������s�5�*�~:�����= �U?R?�p?ގ ?�x��>'����>=�}#��΄=�/�>�h2?{�L?O�*?�ד=Ǩ����d�P`�� B��]ɇ�"��>?rI>��>�I�>%�><�L9s�I>�0?>���>7� >-k'=U�_=�N>�M�>���>�{�>*
@>q>u���'߰��Lh�hGr���ɽ�t�?TD����H�_*��F�����a×=k�.?�c>6�� �Ͽ���HH?����ϊ.��h>�e2?'Y?7K> ����e�Ec>���l��!>����k�x(��mR>A�?y@g>��t>9�3�ab8��P�����V|>�6?q(����8��vu�ǂH�ݾ�OM>�|�>9>=�q]�������~�3�i�Y�z=�}:?��?&	��6����u�ï����Q>�4\>ҷ=���=m�M>F�_��tǽ�[H��>1=�=��]>�?Q�=Zd����>��� �����=�#`�u� >�l?*�5?�->�p���᩾Ȥ����>��q>爼�>�}i�z��<�m�>��>�5'��\s���������>�.;�
�����v>k%���1h>l��%K��L��n/<X�~?n��]؈���꾒V��� D?I�?e�=��7<�"������/��O�?��@�d�?�z	�D�V�y�?�2�?ԫ���z�=B��>8��>ξ5�L���?�^ƽ����	�1"�u�?:�?��-�w�s	l��j>�K%?��Ӿ�n�>~��W������u��P#='��>)/H?�l��A�O���=�Ys
?�?B�%�����ȿ6zv�f��>,��?���?v�m��D��R@���>`��?�cY?�4i>�r۾]�Z����>:�@?NR?�"�>h;�T�'���?�׶?���?BI>���?0�s?�p�>ox��]/��6������-z=P�_;3j�>�a>�����gF�@֓��f����j�&����a>�$=��>�:佲7���B�=P싽+K����f����>�*q>0�I>�T�>�� ?�]�>+��>'p=�p���ۀ�������K?���?.���2n��N�<g��='�^��&?�I4?�j[�z�Ͼ�ը>�\?j?�[?d�><��P>��F迿7~��p��<��K>*4�>�H�>�$���FK>��Ծ�4D�_p�>�ϗ>�����?ھ�,��PS��EB�>�e!?���>�Ү=� ?��!?�Rh>�>D�F��^��4�G�D>�>u�>�q?w�?0�?A����4�Þ���p��N�[���G>��x?FU?/ۓ>���㘝��	ܻD���P���<�?)�d?��㽙Z?��?�0=?��??�si>X�+ پ\4����>k(?�1��F��8(����=�?�L?�2�>o!���7����.<o�!��fS ?	�T?'?�v�>�\�����i�<[M���h1I�l5=$SC>#>s�Ͻ_�=�p�=�w�=��U�� �#�=��n=��>��>z�1��@b��,?u9(����g2�=�fr��cD�c�>S�K>N����O^?�=��
|�r��Ts��@zS�U΍?��?�y�?�9����h��=?�(�?�1?gt�>]B��#�ݾ#�྄v��fw�KD���>�;�>�兼���W�������c���*Ž<�I��J?�h?O#?&�$?=tv>T�?rT�/��?����$��r���A���g������H�C�%�H��=1�e=��վ����U��>Z�c����>��?�a~>mI�>r��>>)�����=b��>��>>�>�=׍,�WĽ�<G�����n9Q?Z)��o�*�߫Ҿg���14A?2�]?���>�����愿���?B5�?[�?M{u>ǎh�Q����?��>W-��X�?ߜ=�l�U�<1j��7��=RŽ�;�y�>Κ�P>�)�G��?o�l?m�?	 �s˶�{�������	�n=�L�?��(?��)���Q�u�o�w�W��S�jU�S)h��d����$��p�>돿]���$����(���*=��*?��?Q��J��f ���"k��?�5of>l��>�"�>
�>'jI>��	�B�1���]�-J'�����S�>-Y{?]��>ƏI?O�;?�xP?tiL?ӷ�>e�>z0��xd�>U<�;��>���>��9?j�-?=0?�v?zz+?�Kc>by������{ؾB?|�?PK??�?�߅�~LýCݗ���f��y������=�h�<d�׽�fu��U=�T>�&?�o��iA�`x� �s>�_T?���>�=f>~T����C����=��>���>m�B>g��&U��	�r`�>�?�[U��;w>��=���<b�J=]�=�8�)�M=��۽����k4�<I�>{�>.aO��X:kT�=�ԼC=Ul�>\�?���>S�>�4��� �ݭ�^I�=�Y>�S>��>�Rپ���%���g��Fy>Jw�?�{�?��f=���=��=Nq���Q��A��p����<��?�K#?}ST?��?L�=?nf#?h�>�-��L��9_�������?�,?�2�>�R��zƾ���m3�;�?�?�_�{v��(%�����m�н��>ۑ-�P�x�m���pE��i�;��D����?8�?}�u�Ζ7�Ϝ�]���N����9D?D��>�8�>�e�>)I)���a�~s�p�;>~I�>��O?�A�>j,?$sF?\kn?��ug�o���Ց���p)=��>c^?o�?��?��%?r�>��K>������}��浼�|?�l�&����tV�>0�>%�>���>�,�<�����Eq=U$e�2!�=�#�=9ٽ>��>o�>�E�>�SN<G5H?F��>k}��!��Ѥ�����b8���t?�	�?��+?��=���E�����no�>&J�?8�?"p)?0�Q�0C�=��ϼOG���ur�N[�>o��>�˚>��=Y}C=u�>���>���>�����8��M��^?>�E?P��=V��mi����>g��XZ�>�t��b'>���r>�ǩ=r侭�h��s�5��v�C�Z��O����N�� ���;?�ؐ�v=\=*������x����>�7�<7�	�=��������i�e��=���=L�e<"��=ͪ�=,�ξԨ�?�i?��?KBh?�>��>ՠ>?�^5��)>F] ����������(�T%��V������[����?a�y{оt�>���4�>�m?>�=pI8<�$>P��=���=�Î;^�=��4>dm�='w�=��l=��>1��=�6w?W�������4Q��Z罫�:?�8�>7{�=��ƾo@?��>>�2������yb��-?���?�T�?9�?,ti��d�>R���㎽�q�=h����=2>f��=Y�2�K��>��J>���K������4�?��@��??�ዿϢϿ6a/>X�:>��>�S���1�7�[��]� �X�; ?�;;��|ʾz�>���=V�޾�XǾ��/=�8>Z=� ��N[����=>By�9=y�h=}�>YaG>�b�=s/���׵=�[:=��=��P>`<��3�2��4��	2=��=��b>nY&>>��> �?�90?\Md?���>9�n�4�Ͼ?X���1�>�T�=ڬ�>��=fC>9�>9�7?��D??�K?�&�>S��=6�>Aܦ>a�,���m�)�)���լ<ʤ�?㫆?.��>� T<
B�����V>��Ľ�t?�1?ja?�ʞ>�X�7M�mo%��.�� ��[;��1=h"o��E����������=��>��>(�>�z>�4<>(]P>u�>8>��<���=xo��볝<kO���
�=�o��hY�<H̼�칗7����.�����:`l��Ա<<��`;]��=���>ӳ>E��>�ל=Ŋ�� 3>���n~K�|��=;T��,�B���d��~�v.�R@9��VE><�]>����??c[>�<>��?� u?�A#>cs
�@Ӿ�Ý�uRg�<	P���=��>�?�r�;�ݡ`���M�g�оL��>�Ŏ>Y�>�m>c,�P&?��Jv=%�gR5�G�>gJ��A���4q��-��⟿ui��&�٧D?B���c�=�~?:�I?�Ώ?�@�>֘�o�ؾZh0>�@���=�� �p�`[��N ?��&?���>�ƷD��Q˾�-罝@�>.[m��xK������$�c������<ܬ>AY��ڽ־�X5������Y����@��{��>2�M?�=�?1�5��p���wD��s�%tĽEy�>yc?��>.��>B]?��Խ�ؾ
�d��='�p?x7�?��?��>���=A��4�>2�?3ʔ?Wn�?s�q?'�S�1��>.]<��+>%󇽍��=/��=�ٓ=���=�S?��?��?6��q��&�쾃'�@e�e��<r��=Ft�>=�>m`>���=O�L=���=�Sw>���>�4�>c�g>e0�>W��>�ݥ�!3���$?>}�=[�>�
3?Tb�>�9=T}���t�<W�>��2<��i-������.��پ<�~Q�=I=]�ռE��>#ǿ-ϔ?<ON>%�1�?*��s����J>��R>�4ؽ!$�>��I>���>�F�>@G�>� >��>�+>�DӾ�Y>���k!��%C��}R��Ѿ�mz>���%�%�^��.����RI�We��f�j��.���4=��<6I�?����h�k���)�z ��ˎ?�X�>�6?E䌾�$��j�>)��>�č>�?��<���gÍ��V���?���?Ac>��>�W?a?��1�}3��DZ�3�u�sA���d���`��፿@���Lu
�#f��!�_?�x?�|A?�P�<5�z>���?	 &� t��e��>�4/��d;�P ==x��>>��s�`���Ӿm	þ<Z��F>�o?�$�?#j?�V���m�� '>ڱ:?͚1?�Ot?�1?b�;?b����$?o3>F?q?M5?8�.?��
?*2>��=�'��u�'=9����ѽ6~ʽ�����3=b[{=f˸=�
<��=��<��ټp};0��+�<u:=,�=��=��>� y?>��>jo�>6?�$>�������Y�?��<;z�����о�8�:���hS>B?�B�?��r?�L>|ρ�V�!���>��>Dy{>>Z>�Y�>u�&���0�=Y��=(>XU�<2qL�_5þ�,�������=�8?>[��>�W�>������W>o4��.&j�'Rq>�s�d<���㋾ŤG�_fK����\��>��o?H�?e9�><����r����i��&(?G2g?��N?g�u?�_��]��b�)���"��"�u�>����+�����ܚ�lq?�}d"�'��>U�D�����a>Y��u�޾.�n��J�!��"�L=�_��~W=�����վ��~�Q��={�	>�E���� ����黪�j(J?zNi=W]���;U�7[��N=>�ؘ>B�>O�:��t�Ol@�����ɫ�=�s�>�4;>�?����tG�����>f�B?�^?A�?$����v�n?�ٓ�П�Ӎ&��N?�u�>k�	?J�2>�}�=M���	9���d�`C��p�>��>����I�o���j����%�m�>��?�&>�s?>VQ?L�?��^?NI*?��?��>�w���w�� B&?4��?��=��Խ#�T�� 9�NF����>|�)? �B�ṗ>Q�?�?��&?�Q?�?��>�� ��C@��>|Y�>��W��b��7�_>��J?ښ�>s=Y?�ԃ?��=>Z�5��颾�֩��U�=�>��2?�5#?L�?���>9�>����{=��>�b?E�?,�o?:�=��?o13>*�>��=R˞>�M�>$�?pAO?�Ts?r�J?ٌ�>;Ў<>����W����t��LT��;�
;<��=oE��y�d �,�<&��;�����|�� ��SA�f܆���;1��>SU�>�5i>8�]�~�I����>�<8=�'ξ�ӾH�ɾ�K�<BN�>1Y	?��?⹋�D��>�a?�48>�!Y�&�k?��?�b�>�Ru��:#�$ھ�M߽���>qE$?R���꓿�3����a��v>'Bg?�mE?H���O�b?��]?�h�=�'�þL�b�@����O?�
?g�G���>d�~?��q?��>�e�9n�I��VDb�:�j�Tն=aq�>fX���d��@�>�7?�O�>��b>t$�=�u۾��w��q���?c�?��?>��?***>6�n��3�(1�m���>p?k��>&����+?�*Z�;����9��y��l���ɾ��ɾ�Ř�nϛ��\�w۝�d����:�=��%?qg?��i?)�V?���A6\��sg�u��J�F����j��F�;���=�!1���Z�����1�������s=,���)�?��?�p#?m�3�T��>W?��S<�D����BX>���l�����=v콯�T<"�e=Ng����'�ԑ��N(?- �>n��>��'?��g�*;A�
L8��t@���㾬�V>�>n��>�r�>Z,u<���p��������O��X��Zv>*Qc?wK?7�n?��'/1�Ɋ��;�!��*1�\���>C>i�>���>��W���|&�yL>�:�r����ϝ��_�	�Ҹ~=��2?�C�>px�>�\�?�?k�	�ޮ�3Sx�f�1�܆<?ҹ>�'i?O��>�Ԇ>�	н%� ���>��l?���>��>Ę��IZ!��{�<�ʽ�$�>��>��>��o>�,�O#\��j��V���Z9��m�=]�h?��`�6�>OR?���:��G<?�>�v���!�����'���>�|?z��=j�;>�ž�$�ͦ{��6��*? �
?i�����*��>h�!?���>k��>�u�?M��>�����;4?r]?��H?�A?�D�>�|=�6���Ž??$��d(=�[�><�Y>�xu=��=���i`��D%�T1=U �=OØ��U��#;�t��ǽ�<��=
50>YoۿJCK�>�پ������/
�9舾D[���N����wb������ax�֍���&��$V�5Fc�a�����l���?�8�?5e�����ǫ��я���������>��q�x�������.�����ɬ�^d!�q�O��,i�h�e�Β'?r�����ǿ~����@ܾ� ?#8 ?�y?P��"��8�� >!�<h��Ps뾆�����ο{���$�^?���>��F�����>MĂ>0�X>�$q>����p񞾡@�<N�?��-?C��>
^r���ɿ����Rp�<���?��@1@?+���,
�LV�=�;>dw>�ߘ�O|s=/!,�����9��>	V�?�6�?�F�>8~�f���g_?���<��z��ʭ���*��>�%>2x���t;58*>�����<M��=Q�>���>m0�=%�(��=��]���0��>�3o�Uƾ5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=s6�򉤻{���&V�}��=[��>c�>,������O��I��U��=Zh��$��M���c=����=�>�Կ��+,=Vޏ=O _�`;���7���:���=�3>; >��X>�g>#�>.�X?��c?#Z�>;�>��߼�X��1�D�$����E\:�72v�
�����.1���/���g,:��C2�8p�f�<�?��=S9R������� �F�b�^�F�F�.?�($>>�ʾ��M�3�2<a0ʾ�^���r���H��%̾|1���m�ğ?��A?�酿*�V�Z�����'�����W?�I���������=����=!��>\ʢ=ў�K3��yS�
�4?���>����P����&-=��ܽ����5�?�z�>J�G=��>�,?��)�;ӽ�'�<v6�>��>��>��=$1���۽p%?��s?}���>d��l��>d���k���w#>w$
>��f��J�=�ף=z�=5Ѧ�S	=h���\�82lW?�b�>j*��W��l�������>=�w??�o�>�jk?�
C?�A�<�k���S�I	
��Dj=�V?��h?l	>u�{���Ͼ�o���5?�Qe?�M>0�b�e�꾉/�Mk��?|�n?P?����R�|��e����ď5?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�ٕ��Z�?�?{����Bg<L���l��n����<�Ϋ=���E"������7���ƾ��
�����࿼Υ�>BZ@�U�h*�>�C8�]6�TϿ)���[оqSq���?L��>a�Ƚ����=�j��Pu�c�G�-�H��������>�樽'�g��k�	%v�֛q��M��)���)�=o7?���<3܅�yl�nxC��i�>�Q"?3Т���D���=Nl�?[���Կ����f=�Et?�Os?��9?D�>|r[�M=l�c����=�Dm?`�?;�3?G%��Ƹ|��L-=v�j?�_���U`��4��AE��'U>3?�8�>@�-��|=�/>!��>j>�/��ĿYӶ�L���f��?g��?�q꾷��>�?By+?�e�05���S����*��#��1A?>2>H���۱!��+=��Ԓ�2�
?J�0?G���-���<?��E��X���5��)��Z_t>�o��_\��w��*�]�#fk�3���ʡc��j�?�	�?�h�?�� �pb�i@8?&.�>����c-�'����&�>7�S>#�=
>̨|<�?�����Q�>���?3��?���>aC��#¨��g>�Co?g:�>���?���=�`�>e,�=���8=.���">��=
�;���?��M?���>>C�=�#9�8�.�u?F��VR�S����C���>��a?��L?��b>�&��6�,��!��>ͽ�1�3A�~;@�}+�3$�!5>Ѫ=>�+>g�D���Ҿ��?y\��ؿnl��Ҹ'�4?)[�>B�?����5u�:�5_?��>�����_��\�{��?;3�?&�?��׾F�˼��>ӭ>�;�>��ս�Π�Az���7>�B?G���-����o�-��>F��?�@��?*i��	?���P��Ra~����7�K��=��7?�0��z>���>��=�nv�ܻ��U�s����>�B�?�{�?��>%�l?��o�T�B�=�1=(M�>Ȝk?�s?�To���f�B>��?$�������K��f?�
@~u@_�^?'vhֿ����oN��Y���+��=��=ӆ2>�ٽ_�=U�7=�8�.<�����=r�>��d>*q>(O>pa;>��)>���I�!�r��Y���O�C�������Z�I��0Xv�Xz��3������p?��4ýy���Q��1&�5?`���=�U?ER?�p?�� ?y�O�>���'�=�N#�P�=C2�>*n2?��L?C�*?��=����5�d��[��_M��4Ň�U��>�gI>`��>p.�>N;�>�r�8#�I>=6?>y�>!	>zE'=N���9=��N>�=�>���>��>�P<>[}>�̴�H2��!�h��w��U̽ ��?�w��=�J�*��?*�����Au�=�Y.?T�>b���>п.�0H?g ��?#���+��>��0?�cW?b�>����6T�5;>���j��D>� �9sl�(�)�aQ>�k?�Pg>#�s>�i3�G�8��&Q�L����Fy>�*6?E����{8�R�t�H�$Uܾ�2M>���>����:�g���~���i�9y=�`:?��?�ֲ���Qs�����J�O>��_>��=��=�EN>3m���½�GH�.1)=Ep�=�E_>/��>W[^=�ߝ=-�>�`�����>{���=1�X�d?)�=?��>4�r>����yb���>��c>T���F]>>@��i�O����>���=�w>�}��3Q�='���z�>��=Q^�>�{<o+><�:��ԅ=�>�y��T��`�>��c?ʯ��0W��h�.@��?ٝ�>	�
>b���97��栿:������?��@�є?�����V�>$<?��?[�<�=�X�>��>�怾�p{���>�Z����˾��5��;��?��?ţ��vx����r���4>��&?���Y3�>-��KX���'����u��n=g�>)H?a��-^Y��>��w
?y{?���l����ȿ�Gv�� �>���?q�?�
n������?�\�>�H�?W�X?#Dg>aG۾M�Y��;�>��A??R?2ٵ>���F'�>�?�c�?��?]I>���?�s?�k�>�0x��Z/��6�� ���:p=��[;e�>�W>1����gF��ד�~h��v�j�����a>�$=��>JE佂4���9�=��I����f�Y��>-q>M�I>W�>e� ?�a�>}��>y=So��&ှp���l�K?2��?����2n��3�<ĝ�=0�^��&?2I4?�\[���Ͼ֨>��\?.?�[?Ge�>��V>���翿8~��餖<��K>5�>QH�>'��IK>j�Ծ(8D��r�>�ϗ>���q>ھ^.�����nA�>e!?X��>oԮ=[r ??*#?k>���>E�׌���[E�\	�>K��>-�?��~?&?����O�3�Xޒ��_����[�9�L>!y?3x?LU�>Q��������T�+"M�C���*�?3Mg?bx��?M��?��>?xA?�~g>T��eSؾ񫽤B�>1�;?DѤ�3W�|7���$�o��>��?I�]<�jT<�\>��Z>?Z���&��Խ>�S?��&?�?.���h��z����=���[+�ɐ�=A�,>��>�eT�/�=�::糽 z�<��<�N>`K
��B>��>]�m=�a*�,?U�*�{����,�=�{r�7JD���>3hL>Œ���L^?�>>�H�{����b��=NT�:̍?��?s�?}"����h�?=?�&�?4,?�>�>Z%��q޾�y�e]v��x�w2���>>�>����_k����k���%��(<Ž�Fk��Ta?� ?�2?�t$?�<|>�J?t (=�K��Q��'��n���C�diS�c�r�M��Ɉ����<�ܯ�?=���N�>z�@����>�E?=1�>�N�>c)�>����;>��3>��>��p>�>jP�<��R�;̈�e�߻��N?���U,�\󩾆ʓ�0?�`?��>s�������t�(?:A�?��?�0P>�q�Z�3�?z̨>eB¾RW3?�oͼ�ݬ��̔;'m���_#�ܾ὞��U5g>2�G���=�S�F�E4|�`w?��?� �����=,p��6Bj=�J�?�(?��)�/SR�s�n���W�khR�����|f�& ��1$�4�p��Ǐ��胿�!���(�IF1=�*?䝈?im��x�w��Yk��=?��'c>�i�>���>��>��H>��	��e1��I]�ɛ&�U�����>vE{?���>�J?22;?I�P?m�K?<�>U�>�������>_�p;���>�2�>� 8?L.-?��0?�i?�,?�;h>U��"����־%?�V?*?�_?i?兾xٻ�D����@��ez�|��@?i=f��<�}۽�tt��W=�S>d=?=�p�VON����k�>��6?b˳>��V>��̾n�x�Y�J>-�?w�>���>�1�� �����%�>5g?�F���8+>��5>�?�=�����ѯ=S�=�0���齲A���<20Z=���>��W=�U�u%�=C>�=��m=YX�<�g�>��?٘�>�W�>A3��4� ���o�=�Y>� S>5�>�RپJ~���#��:�g��7y>Xy�?�z�?�tf=`��=%��=dk��WK��:��ｾuV�<�?rJ#?�PT?Ȓ�?y�=?�a#?�>!,��L���_�����|�?�C+?�)�>֐
���Ǿt]��ʎ4���?�/ ?��a��#۽��A��r��!�=�!-���m��㫿>-H�i��,P��a�����?���?�Z����6�e���-����ƾ�WN?���>g��>�U�>��.�נX�|�\>3>w��>)O?U&�>k�O?�{?�k[?��S>İ8��'��ν���i0�;">�-@?8��?U�?��x?���>g�>K�)��X�f��8l�a��������V=�Y>�4�>)�>岩>���=��Ž���� ?�d�=Z�a>V��>���>W��>��w>��<��G?9�>�A��m�L������U��Ju?C�?�)+?=="=�8���D�U������>���?wd�?��(?gS����=p�ἍQ���2n�J�>��>�Z�>�i�=�6=Gs#>���>{��>9���2�^7�P�L���?kE?{H�=�0Ϳ�`��R�>u�|�l>��G>�����S=��:=�m�ACԾҦ���پ�ш���c��׾.��E���7b�+$?�3��m:?>�5�=-�Y���k��T=���<�B�<N°<W�
�ŀ�"3��R����X�1�� LM=�/>���<��޾Ou�?N_? %?�.g?e��>6E�>��>Q?�.��s�>�OZ�S�~�sؾ)<��-��3l�����ξ����ξ�l#>�x��K�	>d5?>R�*=7�<�La>���=}�>���;<<7=">�? >:&>�t�=�.�=?�=�6w?T���	����4Q�[�^�:?�8�>=y�=\�ƾ�@?
�>>�2������|b�.?t��?�T�?��?>si��d�>^��s䎽�q�=�����?2>���= �2�3��>��J>����J������u4�?��@p�??�ዿ��Ͽ�`/>+fS>��=XKR���5��i���S���v���?g*6��I��t�>Kv >��Ӿ���l�9`�W>ve5=��+��S���=��h��Qv=�=C�>j�>>��=U�����=��=]�=�9@>Yp�<pI��6#���f=eF�=K�Y>(,>�.�>�E?�M0?o�c?謹>�t�UB;6�¾�?�>P�=E��>�=[�E>߼�>�(7?E?t�J?Z�>�Ў=5k�>W��>�{,�P4n�H��	��p�<�χ?xʆ?���>mzv<{�@�����=�<��{Y?Y&0?�?7{�>�U�H��X&�ښ.�m����Jзf+=gr��8U�����~n�ò���={p�>��>-�>Sy>(�9>��N>w�>5�>TV�<z�=Ԙ��YƵ<o.����=������<�rżt≺�'���+�����Y�;J��;AJ]<98�;��=B�>�z>���>��=��� C1>z?���J��h�=�����B�qjd��)~�_�-��d:�~�J>�V^>JՉ�����x�?��]>�A>��?�0t?*!">c���Ҿl��Áb���O��J�=�� >�`@�W�;��`��,M��оy��>EW�>���>d)w>��0�A A�&�>=+��;����>�q��UҼ��ƽe�p����̘��-d��L%���@? s��,��=�y?plN?�Ґ?ڿ>����徠�>��X����<�+�	�_�a����u?� ?kc�>[r���<�RC㾇��'�>Q���V�'����6�Ȗ��r�D�>�ɾAl���<���}�&����7�7�w����>��N?\ʲ?�F��u����R���?�)>���>d�-?Y'}>�P?R��>h�0���ƾj\�q�K>��?��?���?"�4>ϟ�=�,���S�>��?ϫ�?��?�Ds?�?����>�6�;�� >����'��=�h
>ܘ�=ɕ�=(�?_%
?�
?`y����	��I���R]�[d�< _�=�#�>�>�"p>ٹ�= �g=�"�=�D]>Vȝ>=Z�>�d>`��>0��>,��^����&?���=���>�1?S��>ZUM=#���X��<s�B� �=�_u+��꽽J���H�<7�����H=�Y��E��>�&ǿ���?�Q>���s'?��[6���S>�<U>�ݽf�>��B>jY}>έ>2֣>T�>M�>��(>�CӾ�{>4���e!�R,C�3�R��Ѿxz>�����&�����u���>I��i���d�}j�H.��f:=���<�G�?�����k�9�)������?�W�>�6?܌���ױ>���>qʍ>�E������ȍ�+hᾃ�?J��?�^a>�`�>�X?�X?H�4�}U2��lZ�Ću�)M@���d���`�H�������_
�r/����_?i�x?��A?}�<�'}><��?�&�v֐��Ј>M:/�Y�:��4=���>�尾*�`��bԾMo¾p�X J>:hp?Q/�?%?�4U�k�m��'>��:?��1?�Ot?��1?Z�;?����$?3o3>kF?�q?N5?��.?$�
?�2>�	�=�
��o�'=7�� ���,�ѽw~ʽ�����3=�_{=�ɸ��
<��=���<���ơټ�;j%��I&�<�:=��=�=8�>�	v?#��>Ħ�>��1?/�Ih�އ��P�,?_J��n{���ӻ�W�¾;�����>�iE?�9�?��f?[�>�|���a�^2}>�צ>�v^>+�O>\��>�꽫W�Eg�=�J+>�>3{�3�7�<���t3�컩�j_�<��.>c{�>��>���<Y>#���[:���6>��:�:A̾M�!�\2��[,��-)��>D~F?�?�8>�cɾ�)ν�Do�.z!?��B?Y�`?�x?W3�;��w�p�=�c(6����p��>�~��������ᔿؒ2���<"[>�K�������\>}[ ��D;�p�+pD���龁E=���_P=���	��Aj�ά�=���=��þ-0�����ت��|H?3A=����I@�����_�,>~�>�%�>ܺ��J��\�8��H�����=m��>�:->,�E������G����À>J=F?��o?�i?�a˾�犿`*]�q����ʾ�����7?
��>�8?�r�=�$=��߾x;�GN��HZ�F�>�!?���FPt��$ž���S�H���=a�?�`�>ũ?a�o?6,?��?��&?��>rU>k⺽yK��e+?�Ɇ?�{���<�糃�YLJ���M�8$~>1�i?)�̽*�O>��?ω-?�^<?iQ?���>�s>�k	��[\�>ٗ>��2>��K���w��
s?I��>��?)�?�N�}�?���þ�I\�����cZ�=��?q�y?�x]?S`�>
w�>�^ؾX�O��?�i�?|ys??���>��=6�V�FM<ˑq=<��=�E�>#.-?`"?/C?�<.?�h�>׿�<�����'�8Z��������\=߇�<��>��=2�%���ݽ~�M=�x۽ᠪ������Y$���Խ�ܧ�)~�Ca�>��s>�����0>f�ľ'I��,�@>
.���N��K݊�\�:���=/~�>��?Z��>�V#����=���>C�>g���3(?��?w?�y!;ݚb�:�ھ��K�s�>^	B?u��=��l������u���g=�m?��^?�W��'��paX?�m?= Ͼ�.S��Ѿ�g���}�s��>@#�>�+�=��>t?(�?Ũ?��v��v�����ƤQ������s�=�>�i��3����>�5?�w�>�Ft>�� >� ���ʟ��Q�>��?���?�2�?V?>�jl��Xѿ�\�ੋ�0L?oü>^���q?*W��ݾ��������\.����ʾ>r����Ԑ۾���� ��Fd��ly_=F�'?�'�?��?��?���hum�|'p�����gRt�1ɾ���n<R��8��4�^��գ�܇���d����<�޼�}c�'��?�,3?6	ľ��>�զ�
�	�����=����u|Ͼ7���7�⽇��w��E_"�g3a���־��,?�G�>��?��O?��^�zq�A2�����=���>�?�>��6?�'u>h6��1��:0ؾv5����4Iu>!Tc?Z�K?��m?�����0�������"��5��_���E>�>�u�>{Q�� ��&�q'>��Ps�ĥ��H��:
�2ev=13?��>�:�>���?��?k��>ٰ���x�"�0��ͅ<&��>��h?���>�,�>�*ս	0 �ɹ�>��l?I��>%�>r����]!���{��V˽��>�
�>���> �o>�g,�<\��h��ن��Z"9��V�=��h?�|����`�8х>fR?�7�:@CJ<��>��v�M�!�����'���>|v?�̪=�;>Bzž[���{�U=��b&)?�?ē��b)����>�,"?}��>�b�>�7�?!-�>�����1K:��?�V^?1K?@?A��>�=V�Cǽ��&�B�"=���>�[>��c=��=��]�\����RN=�(�=?Fؼ�q��Ӯ�;�۸�V!c<��<3>�[ۿ�#K��+ؾA��_󾾖	��a���緽�>�����'����v��S��a����=�u�Y��^�[����l��3�?@m�?^���u߃�Z���O����� �^��>u�y��s��W���@�b���/���S�!���O��uh�W�d�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾x1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@nyA? �(�8����V=���>�	?�,@>2�0��6��	��83�>�5�?��?��M=b�W���	�Ime?�<��F� �ۻ�K�=	!�=�#=�%�4�J>�/�>�|��A��*۽S�4>I��>�h$����ݕ^�u�<G ]>}ս�P��5Մ?,{\��f���/��T��U>��T?�*�>U:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=r6�����{���&V�}��=[��>c�>,������O��I��W��=o��+�ÿ�=6���8�]���U62=�/�����1��
�������z$�S�m�h���=��%>���>B�r>oT">�cS?Q�o?���>�e>L%���Ӊ��Ͼ�lϽ\�˾��6��M ��5ؾ�
�%������|�����$!=��
�=7R�A����� ���b���F���.?w$>@�ʾ��M�w�-<Kqʾt����ބ�$ॽ�-̾��1��!n�͟?;�A?�����V�p��`U�T����W?)O��� 鬾m��=�����=�$�>.��=Q�⾣ 3�e~S��k5?��-?�C���h��ǿg>��[YG>>�"??�}>![>��F?k��P/��B�>��>�>��$?j??]����A��+?��7?�6ż!�p���>��˾�c��1wѽ��=���� 4=4�>�p	>*M���>�� ���P��[?��>�!/���$�^�����.�I'#�,J~?ip:?
�>�B?��?m�ݼ��!�v�+��1A�,<�vg?�?q��=`�y�Z�����?��]?��Z?�u�>#���%%�<�'�ڽ�u�F?�=H?��
?Ke��xA��	���,���P?��v?s^�xs�����O�V�d=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�%Þ?��@���?��;<��V��=�;?k\�>��O��>ƾ�z������3�q=�"�>���ev����R,�e�8?ݠ�?���>������sj�=wu��_v�?TΈ?�Ծ�ԟ�]��q7��m"�g{ĽKn�>-as�g3����� �S�K:�_p)�����&?���>^�@��=7L�>�E��Z������].����𾡊��-8?G�	?�L>����������X�+�Y��Y�Ͼ�?�>��>�7��@ݑ�X�{��f;�ܟ���>�g���>�S�4������\�6<Fƒ>���>െ>Zl��E�c��?j��B;οo���Ւ�	�X?�f�?<q�?�t?R�7<`�v�Z�{�<��s'G?�{s?�Z?�l%�P"]��7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�%�>��?Jl�=OU�>qY�=���z.�eE#>1!�=o>���?�M?�V�>N~�=��8��"/��\F��HR�U&���C��>��a?8�L?�\b>���N2�!�vaͽo1�����Z@�y�,�[�߽�<5>k�=>7$>��D�	Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?kQo���i�B>��?"������L��f?�
@u@a�^?*HiԿט��/���?i��?�=��>��G>�3����<&���@����,�a���X�>�B>��A>���=JK/>i]>z�����&�S���[��|U��@����j���ھ9��ʁ%���Ӿ�Ҿ��)�<b����P=�?�:����Eh��9�=JUU?�PR?Gp?� ?Hu���>����U�<�g#�A��=�>�2?��L?�	*?E7�=�|����d�ah���馾�M�����>K,J>���>���>*��>��;��J>�=>z��>�>^�%=���pG==3O>��>���>�ʺ>�C<>��>Fϴ��1��j�h��
w�j̽1�?����S�J��1���9��զ���h�=Hb.?|>���?пf����2H?%���z)���+���>}�0?�cW?�> ��k�T�6:>9����j�3`>�+ �}l���)��%Q>vl?��f>	u>��3��^8�;�P��q��q|>�26?j붾K9�M�u���H��iݾ�NM>︾>�D��k�����{�"ji���{=�s:?f�?1A���.�u��@��:R>�>\>��=�N�=�SM>�]c�H�ƽH�G.=m��=c�^>v?h*>%��=0N�>��L-N��g�> D>2z,>�Z??Վ$?��������S����+��v>��>�ځ>�l>}�I�$r�=X��>-<^>��#S{�ߨ���>��eW>�"r��{^�*wy�2q=˙���=kr�=����=�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>Tx�~Z�������u���#=6��>�8H?�V����O�&>��v
?�?�^�੤���ȿ9|v����>R�?���?a�m��A���@����>;��?�gY?=oi>�g۾`Z����>Ȼ@?�R?%�>�9���'���?߶?ԯ�?_�d>tϖ?Rbr?��=8��9�f��Ͼ��.���AD<���><?zѫ>z��>��(�����i����6��D�=QN�=�S�>O�L�U�辟�@>��=q쎾Z����v�>���>�uY>�U>�1?|�>7>i���>�;N��;dT(�9�K?�ݏ?�T���m��;�<��=��d��	?��3?$��!�̾s��>�]?D;�?s�Z?N��>6�vc������T?���ی<��I>e�>�g�>�q��2L>��Ѿ<�n��>��>���#=ھ�#��0?�:���>D�!?(�>��=�U?�
2?��>S�[>�L��%���Z���g>��>�=4?�h�?"�!?� J��-��c���6��:�i�E��=T�b?�_?���>Ft��;���Fg=���= �7�.O?8A\?�Y=��?�n?�3?�;Z?�,7>>�T��&��vt�=��>��?�pS��F�4�{�<c�?��?���>�a��N,��A3b;�b��'�Wz�>�Wd?��?����	:�ƾ���<��_ׁ�aߊ���4��S
>t�=�W2�E��=��H>o�>}O����M�����Oq$=B%�>�=�p7�,��o>,?�F��߃�{Ę=:�r�9zD�8�>}^L>����~�^?�o=���{�����y����T� �?���?�k�?$ᴽ��h��"=?��??,�>�F��Av޾L�ྦ[w�tx�u���>���>��l�Y徏���y����C��b�ŽS]{�-�>�� ?h=?t�t>:�>�(|>��m��0�;��1�۾qi�yR��o� �x�f�'D�Λ����h	������
���ʽ=+ϗ����>1�?���>5T�>p��>*��>z3>��Z>��}<��>�.>h->[��<��<*�e=t@R?}�����'��]辦5���'B?�rd??�>Ii�
~����k�?^�?�^�?ݸv>]Qh��
+��f?��>��>a
?�9=�u�R�<n��U������׀��>�ս-:�#M���f�Z
?��?�����g̾��ؽ���)p�=�_�?C*$?U/�7gW��*s��3U��S���.%A��x��)�e1o�{E��fm��gD����0�H�?<�T)?>��?~��k���勭�D�j�N@�8�L>�x�>�}�>OƼ>Y�_> ����g3���Z��"�ţ����>6z?��>�j6?�??��S?viJ?���>�˰>����ͩ>�F���b:>'A?%}2?�2?u"?��?�B?��>���=��\�O�?�8?�)?���>O�?lS~�&�������=ܤ�6����=j�=p�L���ѽd��X�<�=�	?�2?��B�m�[d�>�8:?A��>�E�>I�l�ir��a�;ߞ�>01�>�#f>��߾��T��	�'��>�q?g�Ǽπ.=�u!>K�T=��0���<f�=�r�;��=/��<�2[�B��<�ڱ=��m=����~=�|[��-���<�x�>4�?�>�9�>�D��Ϭ �T��ލ�=P1Y>�%S>g
>Nپ{|���%����g��y>�v�?�z�?@g=��={��=�z���P��r������?�<�?�C#?�UT?���?3�=?Fg#?�>�+�nL���a��f���?q!,?��>�����ʾ��މ3�ǝ?Z[?�<a�޸��;)�ː¾��Խ��>�[/�i/~����ED�U��������*��?⿝?�A�N�6��x�ݿ���[����C?"�>Y�>��>A�)�{�g�u%��1;>��>gR?[��>��r?
CG?�>_��=��>�������=P
?|I`?�z^?���?C̋??��>�sL�r(��i8��4���C;:��:��״^>x�>�~z>���>���>�>�<��%���(}^�GŻc�>=�?վ>���>�4�=�q��bO?�W?�߾��"��V꾃�ξ��H�=B}?��?:(%?�`Ƽ��>���+�6�!��+�>�|�?�o�?��;?s���M�=��X��2��ѪU�	��>/��>��O>W�>���<ru>�E�>ݏf>��k�4�,�H..���/>��h>��]?{�>�h���t�,��no0��pL��� �23(��Zv�Tya��k�@f��J��� ׾S�!�+��!���y���d��k�p�e��>��<T(Ѽ��;ȡ�<&��s˱=oj= ��;���=b'L=�	��
���ME<ۤ����B��^�����$�˾x�}?�;I?�+?:�C?M�y>_;>G�3�ߙ�>舂�t@?�V>�P�x���ԇ;�5���� ��[�ؾ�w׾��c�0ʟ�2G>�bI���>r83>�I�=kO�<��=Ms==� R�=�#�=NP�=gf�=s��=��>FU>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��A>�&�=��S��{-�`�C�ĜM�@�?��E!?�~7�4�ʾ��>b��=a��[���dv=�3>Y-K=1%�w�Y��g�=vr�Z�=�u:=Ƌ�>�pK>꿷=Kޛ�`�=%8�=���=&�<>D�`�$d��@p���a={�=9
]>�(%>'��>
.?��/?�c?�?�>�Lo�ncϾ����l�>�S�=Ӳ�>\��=�GC>�y�>=�7?��D?Y3L?C!�>I��=o�>Q��>�,�`�m��K�$���F`�<~݈?6ֆ?ao�>q�F<҈C������>�e�Ľ r?�1?�#	?~�>M���߿~�;�O�B���R��n�=
M�=C* �	퍼z{'�TQ_��p�B�9<�k:>���>�v�>�ͥ>�UK>��=��>�c|>L� ����Ӽ�fn�W�<�@����������� w>��}>2�<�w�<~/���ֽ1>��>)Q��t��=���>?A>���>���=����B/>:����L� ��=kG���,B�"4d�yH~�C/�.W6��B>58X>����3����?h�Y>�k?>x��?MAu?F�>����վ�Q���De�8TS�ø=J�>��<�9z;��Z`���M�`zҾ���>��>�>��l>^,�{%?�ӆw=�⾅a5���>�n��������6q�C@�������i��Eٺ��D?�D����=~?F�I?�?���>	���ؾ�=0>�=��,=���&q��8��)�?�'?	��>X��D��H̾�����>�;I�f�O������0�����ͷ�ێ�>I�����о$3�#g��=�����B�.Lr���>K�O?+�?�;b��W���TO����)#��?r?2}g?c�>�I?�??�!���{�,r���t�=��n?#��?=�?�>�>�=���I�>(H?ӣ�?^��?�%t?�!�{��>�� �E��=
`����=��>�6">��>eP?=V?�d�>����F�zp��� �'p�%s�;Y�m=B�y>���>>ٷC>��=@S=?:@>s��>�p>�@>��|>DJI>��q
�\�5?��C>�[U>��3?��b>u�,=c��	+<���Ev��l��Mw�۟B��Nm�hk��f��6vP���*�>�Ŀr��?Y\>�����?X�;v�=�|>��>����>��>��}>�Ƙ>�~�>�I�=q�>�oS>5ӾƱ>�vP!��>C�/�R�-�Ѿ|z>5���w�%�1p�F����H�z���|�#	j��0���S=����<;�?̓����k�_�)������?,^�>��5?����1��u�>��>���>8��񎕿����F��?i��?�:c>Z�>x�W?Z�?��1�3��uZ��u�j(A�/e�'�`��፿������
�����_?��x?�xA?dP�<:z>#��?�%�oӏ�%*�>�/��&;�SC<=�+�>m*����`�-�Ӿ�þ�7��HF>a�o?%�?hY?1SV�ت���;>b|)?�-?Lr?�/2?��=?j����?��>�x?:>?7�+?8�,?�S?�{.>ʦ�=񞵻a�<����芾�3�+�ֽm8�:j��<���=و2��e�����<�Ww=F_����B���<�d�����
^=�M�=}/�=��>J�]?}��>5e�>�;6?"� ��|7�^©�@�0?ۯB=.��~�;�������n�>ìl?��?o7[?g�p>m&B�l�C���>�ۋ>2/>A�]>���>�� }M�LQ�=9�>s>7�=͸G��[��R|	�&�ND�<�#>���>|><2��ѽ'>�j��'z���d>��Q�HϺ�k�S���G��1��v��^�>A�K?K�?���=iX��B��-Cf��))?�T<?NM?��?z�=%�۾9�9�4�J��9���>*��<"������$��Q�:����:B�s>�!��
M��?�]>����N޾5�l��zF����/=
L�&b=�	���־�����=l��=�F����"����'l����J?��u= ���TV��;��Fe!>�̐>>�>��0��dl�@�>�@����̵=7i�>�Q4>Ӈ��DD��@�u�>�K?�R?s�?�_x��t�/�4���)������@P?�ߥ>u��>|]]>.� >�2���*���a�s�U�\��>�d�>U�
�A�G�8���Jξz ����>-�>N�r>oz?ْB?p�?ӈ_?|�.?��>�c�>��h�����'�&?��?ʑ=�~�3����8��|9�u��>v�?�2/�U�>��??
�?�pf?��	?x�;>����L����>7`�>�QH����N=�J?�n:>1	t?y�R?<5�>����̾#�ǽ�;��<n>��,?�@?��:?U�>H��>T�%��;�=�2?���?�Hz?H�t?��u�]�K>�����u����J�>أ(?�n:?�$\?ԕw?�pC?Ҵ2?U�;�U�j�N��EX�����9�<�d=T�7>/g����=���=�W=z�`�c�nw$���F�F{|�w���&=�x�>7%t>#B��m�0>}�ľΒ��g(@>8���\뛾�݊�at:��D�=T��>)�?i��>��#�s�=�P�>8�>:���?(?s�?W)?�*%;�ib��0ھ1�K�$��>v�A?,J�=�m�"���`�u���e=n�m?h`^?KW�%J����r?+�N?`1�o���x&�L@��v?61g?:�t��5?���?;�b?+R?���-Az�Y0��3�r���e����=Y�d>Hf&�\-p�
y�>��?_�>P�s>���=]� ��^���x�x�?`�3?t�?|i?~�j>��h���ƿl����;��_�]?�n�>Ħ�k#?ߌ��]Ͼ��u����*��n��Ur��b��.��"&�2���ٽ�A�=�>?6Qs??�q?:�_?� ��Tc���^����EV����j��̬E�W�C�{�B�r�n���i���n���==Τ��RS�8߻?��>K��%?�©��^��g&����>��`���w��O�'����.�
=������N��
��&)?-K�>ô>%� ?��x���V���F��\E��j���H>'�>�>J>a�?��=m��� ��<}��{,�6����c�>%�l?��?n[l?]"���C���e����Ji=��޾��]=��0>��=�����5꽆D(��T�Pn�СD��Ϯ���ξ���>�r:?���>x߳>���?�.?���X;�t�]�O���0�Fk�>��R?�"?5C>%3<15*�q��>j�l?��>��>����M]!���{��ʽ�+�>ۭ>3��>^�o>�,��$\��f��'����9�'i�=P�h?Z�����`�N�>�R?��:S�I<���>�v�K�!�.���'�P�>Nt?��=d�;>xž�#�Ι{�4>����?�6�>�ƾ��3�'�V>K?�?���>��?'��>�$־u��
/+?�T?!?��$?�l�>�<%$�o���%�۽_�a=�E�>�i>���<���=��9��$W��H���h(�Ш�<�lL��Y���@�>W|<��u=/y<O�e>�hܿjI�W=̾SC����!��I|��t ��{�ƽ^◾BR��<O���x��͌��m-���.�������쁾��?��?��+��J�DÐ�l�Z����ق�>HQs�z�l���� 3��8�u��r�ྩ���J�{^�;o�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾{1�<��?7�-?��>Ŏr�1�ɿc���x¤<���?0�@#{A?��(���쾯YU=3��>U}	?V�?>�E1�1*��밾.R�>�:�?���?�xM=\�W��w
�<ke?
N <�F�e��g6�=$o�==���ˈJ>k�>=f�fA�ܽ�4>ï�>Ɓ"���i�^�G��</e]>y�սɵ��5Մ?*{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?6ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=�6�����|���&V�}��=\��>d�>��,�ߋ���O��I��W��=V?��Fǿpb;�y�`�y�$��&\=o3=:�z�kA\��k���3��0������ֱ���={���k�<<�9/=��H>WI?7�l?)m�>O`>�O��9�X�:�ྣ���ƻ�����q��9��=H���ξ�~�D4���3�k���m��$=���=9R�Ǖ��>� ���b��F���.?P�$>4�ʾY�M��0<�`ʾ ���Xy������2̾}�1�: n��ȟ?��A?����V�������t��"�W?0^�4��J��_�=�[��>=��>K��=!�⾥3��}S��2?�u8?Iy��T_��t3�=�������=G &?���>o4��l>W�>��R�����Am>���>
��>+�!?஗>�ǵ���L5?xY?��<,<[��k�>1:�O6W���s��2�L��N��=zG�>E>A+�f�>������<��[?$p�>S���k!�M���k�����T<�9�?��>H��>��s??�=ϽK��DH�c�ɾD��=�s?isu?W�=����̾��%��/C?]rc?�2�>�鮾�춾��Z�z��	?��W?2J?+8���_d�Mo��E���#?��v?�r^�vs�����X�V�a=�>�[�>���>��9��k�>�>?�#��G������yY4�$Þ?��@���?��;< �L��=�;?p\�>�O��>ƾ�z������D�q=�"�>���yev�����Q,�d�8?۠�?���>�������k�=lנ�0W�?��j?��߾1��**�ߜ?�PG6���O>e[>�D?��m>�ľ=�i�h۴����ҥ������Y�>�@�Ù��� ?���������ȿNÅ�;����˾úC?h��>�)�/�'�~�l������	
�-c�T����W�>�>:���T���{��o;�H����> �R�>N�S��"��*���Q-6<	 �>���>S��>/��ｾ���?W���8ο����ǡ�L�X?�\�? q�?�c?��;<��v���{�0��G?p�s?�Z?�|$�z�\��6�!�j?�_��yU`��4�nHE��U>�"3?�B�>P�-���|=�>���>g>�#/�u�Ŀ�ٶ�8���Y��?��?�o���>n��?is+?�i�8���[����*���+��<A?�2>
���D�!�;0=�_Ғ���
?O~0?{�k.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?&s�>���?���= 9�>u~�=4���s���>�	>KJ���?�Q?l,�>��=�/�:0��JF�x�S����O�C�N}�>Rb?0�K?�V_>@����) ��߽%�2����wEN��x:�����B�.>��:>H�>�?��'Ծ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ua~����7�c��=��7?�0��z>���>��=�nv�ݻ��W�s����>�B�?�{�?��> �l?��o�P�B���1=:M�>Μk?�s?�Ro���\�B>��?!������L��f?�
@~u@`�^?)&[ڿ��s^־_"�8��<˝�=��>o}/��5=Ѯ$����
C=V��>��=|�;[9>}Y>zd'>}
>�\����#�\���j���?��������ʧ���Q.��?�վ~̊��s��+�n�?-ýʨi�n�z�sD]�k��;�=��X?��G? �s?W�>5B�vt>���2�\=�-]�8=��>�G?H0C?\�)?4�=!���	c�G���X���ޥ���>��9> ��>s3�>ﴦ>`t�;��3>��Y>T�>�� >���=��=�Ҋ=0w>9��>���>Q��>�D<>�>Nϴ��1��V�h��w��̽� �?2���6�J��1��8������h�=Xb.?�z>���?пN���S2H?����)���+�R�>��0?�cW?��>��m�T��8>�����j�m^>�+ �ul���)��%Q>#l?��f>��t>J�3�!Z8��P��y���|>�86?����]9���u��H�*ݾ?�M> ��>~�C��U��햿,��Wi���{=�g:?~?��&߰��u�T2���R>��[>Q�=�'�=�aM>�Qc��ƽ�G�70=�\�=l�^>>?ʹ'>�s=�u�>:ۙ�W`K�Y�>E/P>�S1>va??ܟ#?��CY��CF|��<-�gUv>ƈ�>M��>��>}�I�wJ�=��>�Ae>��������	���?�Y�]>Z���jn���k�:	�=�<���W�=�
�=ĝ�F@��`=�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	�ߢV�@�?�@�?��I��=}�>׫>�ξ�L��?��Ž5Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l�6>�^%?��ӾPh�>|x��Z�������u�{�#=R��>�8H?�V����O�e>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?toi>�g۾:`Z����>һ@?�R?�>�9���'���?�޶?֯�?�I>N��?��s?x{�>x��^/��/��`����=8O;�X�>MW>x����^F��Γ��a��w�j�G��~�a>�$=��>J�f-���,�=2���@��n�f�@��>=:q>��I>S�>=� ?%}�>���>�=iՊ��ڀ�������S?Y��?B'�-�`�*���
؞������O�>V�P?�,�����cd?@�c?� d?|\?��)>��e���'��c����H�=���>��>��>(�|<��>��;�����Q[>f)+>��$���׾�඾�%7�	��>�?q*�>���<�N(?�"?�IR>`�?��i������m��L�=���>tz8?#C�?��T?]_������ē��}��]�4�G=v�P?��#?�K�>~X��Ǝ��G�=`t��Q��?*M?']�?Q]���ʑ>�^�?,z#?c�<? 3�>�Т=���3w<-��>��?�`-��tC�>D*�>]�5&?6�?!�>�������:������}�?:�R?��?�����W����>��<��j��ٹ��Q<;I��dR >(�>jJ_����=G>�h=��e��R�>S�;;ˤ=Ʒ�>�'�=�|D�?���@,?g*D��փ�ʐ�=��r�wuD�E�>�L>R����^?G2=���{�����|��z
U�  �?F��?�k�?~���P�h�#=?��?9?["�>�=���_޾ʟཱྀCw�݇x��p�}�>���>�$l��#�=���e���*=����Ž�^�d:�>�>�?RT�>R�H>��>N����%�q���c�3b]��\���7���,���Z��͹&�A�6�p����/{��K�>g?��WN�>X
?J�h>Ն|>���>����W4�>�xP>oG}>b�>�][>)Q=>�>�2<��ʽBR?b�����'�t��B����%B?�id?�4�>��g��}��$��wy?!��?�m�?�2v>nh��+��\?�0�>����f
?i2:=�?�h��<iK��/����e���>s�׽#:���L���f�b
?�)?�ٍ���̾�m׽S���D��=y*�?�89?
F�Xe�����G=P�:Ps���?=k=��������M������唿B�o� lB��Ȳ���0?��?^���G���5����t�G�H�S �=��?g9�>{h�>3A�>{4��$���:�{�F��h����?eۈ?.u�>�0M?.?c�[?�aK?�4�>��>K� �pd�>��������Cy>gj?��?? �9?�P?�T_?&z�>�>���u'��-�?�m&?�%L??���>��߾.������;���!��x缨�	=��>[@�;�u�@���t=G�?�򛾹�C�/���b>J+?��?7�?�ʽ^Q[�H�a=⇚>��?Q��>����O���Ѿ0��>�V?�o¼iG8=��>u��<~�B��|�w=o��=ө6>�=3/���s�<R�B>�=J�5�r����R=.���Y��P� ?� ?!ˉ>9D�>l,��Q� �E���l�=��U>�Z>ߓ!>��ھv���Ř�*�f�}�}><�?�X�?�}=���=���=����O������D����=��?>{"?��R?�?�|=?#?�>��Q풿C$��������?�#,?@��>���,�ʾ�憎x�3�͌?Q?'*a�����5)��n¾��Խ�>
T/��1~����CD��∻����9�����? ��?LA�V�6��A�躘�Mo����C?��>,�>��>��)���g�w �E;>���>��Q?�*�>��O?��z?��[?��S>[�8�p���P���D"�H >��??d��?U��?��x?b��>�>W�*�Eqྸ3���,��L�R��&�S={�X>�>���>ʳ�>�9�=_Žs��(�>�nU�=Y�c>D��>_��>Z�>�Gw>���<�S?4*?���D�#� L𾷭���6����?�b?kB?�bK>��'��X�7�$�}��>Y��?��?�y;?������=�˒=n���|��8f�>���>."�>9��=7v7=�;�>:�>Y9�>�d
���8���p��,�;ݱ�>A�[?��>�繿�6��kk>����,q�=S0���k��_>�b?��+x>j�,��t���v���z��\���������
���R'��<�>|!k�7�>��2>�0)>T�=#�=OYm;�J|���.>P�H���=��3�F�3s���y�'<��r=�ׇ=|�˾p�}?<I?	�+?��C? �y>D9>Cw3����>n���@?�V>��P�ň��4�;������#���ؾ�y׾��c��ʟ�)J>iQI�^�>�93>lI�=aO�<0�=�&s=�Ǝ=ݡQ�=�%�=�N�=Wg�=���=z�>'X>�6w?T���
����4Q��Z罣�:?�8�>{{�=��ƾn@?��>>�2������wb��-?���?�T�?B�?.ti��d�>O���㎽�q�=+����=2>���=��2�T��>��J>���K��4����4�?��@��??�ዿ͢Ͽ2a/>��7>�N>��R�HW1�%�[�ƅb�	dW�n�!?ص9���˾�>�y�=�kݾ�HžG-=��5>~�c=ʢ��4\��D�=jx���>=�l=���>C>�=�����!�=�D=q@�=pON>�䣻:�K�+�L�7=:��=��a>��&>o(�>3%?L%?^�V?�@�>zł�ݹϾe����Ou>���=�>��4=ah>Ŵ>�I?^�<?g�J?磣>a����0�> �>�&���`���o�� �x��]�?n�o?���>
�=�ׂ�����H��UW��o?�&<?Z�"?e��>DV���࿠\&���.�朙�����s:+=/{r��yU�D���6\�p�㽀��=Q�>t��>OΟ>�4y>��9>��N>��>��>)��<�X�=O�����<v�����=X��A��<��ļ�E���:��,����Ӯ�;$n�;\<7d�;+%�=@��>T�>) �>iT�=gݳ��.>��x�L�x�=<���WB�16d��~���.��n5��6C>^�Z> �����&{?�Y>��@>Zy�?�Eu?]�!>y�,վ6�����g��R�BJ�=��>�C;���:�8�_��}M�QҾ���>4�>�\>Bo>n-�}�K����L^�v�gd�>"��`N�=(����v��阿TH����i��P�� I%?��M�.>��?V�T?f�?pK�>~�/>�c���j/=v����\��n;�;��������>�!?1��>I���O�xV̾ ��_�>GHI���O�^���)�0����ط�Ӑ�>�몾L�о"3�0g�������B��qr��ߺ>��O?��?
-b��J��yQO�U��"ۅ�"d?��g?��>�H?�<??F��L[��W���X�=l�n?���?9�?G�
>�1�=G�@��\>3E�>�Ĝ?#ь?�l{?�U4��9�>�T��H��$7ǽ: y>��>���=��!>��?��?At2?����X��g����07��32	�#��=5�>��> �>�0o>w+"=,�=DQ�=m&E>��=�7��y�:>��>.������UV?~t�M�>v0>?��=AR5>��M��	>g�=%���Ʈ ������y�q<P���m}�\
K��?�>�T���<�?'4(>�y��W�?�%���W�>�>??{>�Yƽ���>��<>��>���>ڨ�>��=�h�>7�>IFӾj>����d!��,C�W�R�O�Ѿ�|z>����^	&����zt��]AI��n��Hg��j�N.���<=�z½<�G�?����[�k���)�����n�?R\�>�6?�ڌ�j����>���>zǍ>�J��K���(ȍ�hᾓ�?���?r<c>��>��W?z�?��1��3��tZ���u��'A��e���`�6፿����j�
�q ����_?]�x?�yA?�h�<�7z>���?��%�}я��+�>2/�n&;��2<=�*�>�)����`�k�Ӿ3�þ8�]JF>N�o?�$�?*X?KTV�ŋ^�si(>@�9?�#4?[�v?3?f�<?��$���!?�� >67�>��?��3?��/?��?�C>�?>��<�>R=�7�������ν,�Ƚ�z�e�=�m�=3�<O�Y;�V&=O��<�G� ��B3;<�����^|<A3=���= �=��>�?]?��>ԙ>��7?b�齴>#�$(��;�"?�F��
�������ؕ�#�ξ�/>v�t?w�?��`?N��>|�K���X�9,->'ܗ>p0a>�-|>�G�>��,���>���=%��=��%>h��=�0_�'Y��� ��q���e��N�>V�>P�|>����D�'>#ţ���{���b>��R�Ƕ��z*T�0�G��'1��>u�Hi�>c�K?�U?1�=��龀闽�[f��N)?��<?|M?K�?ࠖ=��پ�9�;K�Д��>;A�<R*	�i���g%��T�:�J�9:�t>r����ݸ�0(Q>e���ƾ��`�EA�)���%<����=�g���csH�Z�<5��=mD�u�����(����G?#��=��m��WD���ʾ��J>�v�>��>����Hʽ�4��]о�p�=�e�>��>��|=c���:pJ��0��ǐ�>�L>?��J?D`|?)���$j�̬4�6馾d_������?���>���>{�C=J�=��þw+���K�q�H��: ?�O�>�!�(�I�;�������7�Lv�>�ȫ>��>�%??/�u?n�??ۈ?{w?�v?�>O�><'��5;?��?r=����z���]K��#<���/?D�	?ǐ�M��>��)?��?�1?�F?z�?7��=Q���/<�H=g>��>��.�l:��B�>v6'?w�>;PT?h�n?��>�J��ԾdX�=��4>.��>�rJ?�Ʌ?�>?\��>��>�u���������>�?�0k?���?��ν�˻>��=k�C=�ё>
�J>�#?a�=?�Co?t�T?W�4?�%?���;QWa��D��i/��Ί�&z��Q#X<%[�>tu>a��;l���=�w3>�M�~���K��c�J�I�3�t��>�Rt>�蕾]�0>�ž����@>�6�����Ȋ���9����=1��>�?Hޕ>�"�#�=�Ѽ>��>C���((?�?K? �;xb�&�ھw�K�9��>��A?6`�=��l�z���u�%k=5�m?�^?�V�k���q�a?p�_?�N�u@��Ǿ0j����JM?\v	?�t1��)�>��~?�Ok?FL�>b�w�� o��l��"e���Q���=�!�>W���Dh�T��>�w:?9��>��N>v��=	|˾aw����
?u�?]a�?�`�?�s(>�ol�~ݿh	��⍿LG?���>����J?�<��6jؾT�f�a�o�xQ��-$��x��aþ�¾�둾��k�g\�5g0�G?K��?8��?�lc?f��N�K�v�[�@Vy�[�7
�P����S��
E��Q��*w�G.�wE��Tž�����B��W]��	�?q�"?�5x��?����C m�������>�<{�0-��2�� �w��,>�;⇙��F�r�ɾb�1?�n�>J�>h�?�){���_�G?� �H�xn���T>y>H�c>(�?���=z�_��2���:���6��L���ǒ>F>X?Q�?=UQ?P�~�l"!���g�)�1Q�=�3����>��>ڠ=�u�2�H�)���M��z�S� ��ڢ������=Ogj?�u�>.�>D��?��?�tľ�I��i���S�%fF��I> �m?,?5Q�>h=�N��}�>q�v?L�>1�=�Ǭ��q�\���|E��e�>��?h	?���>n늾�Zb�)C���!�F����fY?8Iv�2���Z5>�p?������	�r�>x�ս.�꾟k�T�l���>,_?Oj=;sh>����Ǿ`�:��ɾ7X(?���>x����+��U�>.V?R�?P�>�)�?��>'�ξ���=��?*�\?��E?�@?Z�>(Q>i'x�R�����h�׺R�y>� W>�=#-�=�A���K�!f����<0.�j佄xv�]�<�i]�Nw=��=S8>_Aۿ�J�`�ھ�S���߾$i	��B��L�ڽ�u���꽜nþ˭��^�K�VH@����_k��R���w�z����?�0�?��<�+R_������t�vH��h�>'���53�����:�0���eN�������&���\��bm���g�P�'?�����ǿ񰡿�:ܾ5! ?�A ?8�y?��8�"���8�� >NC�<-����뾭����οA�����^?���>��/��p��>ݥ�>�X>�Hq>����螾1�<��?7�-?��>Îr�1�ɿc���q¤<���?0�@�uA?��(�E��n�S=8��>^�	?�|@>6�0�t�����>�K�?��?!�N=��W�$��Ode?�<�F�f9ػ���=-פ=�=Z���J>A�>�m��A�[\ܽ,14>�Ӆ>�$�e�"�^�:)�<6]]>:�ӽ�q��Մ?�w\�f���/�~T��O>|�T?�+�>b7�=1�,?�4H�}Ͽ��\��*a?�0�?V��?��(?�Կ��ٚ>�ܾX�M?�C6?��>{`&���t����=���5֥�
��X'V����=��>؊>��,����}�O��*��d��=A��8Gǿ�"c��0� �>^� �pǽ ��(��=�$�<ۿ�Dg%��w�>Ǣ>�D=�#�=��>��>���<Q�T?�o?u+?�ϴ>�9����Q+�@��=�^6���l�#�Խ�ڽ��վ5��0�z+�!�#���k��D#=���=�2R������ �D�b���F���.?�t$>��ʾP�M���,<�fʾ�ʪ��_��4��.̾Ӕ1��%n�3̟?T�A?%�'�V����oy��Q�W?�O���?䬾vk�=����=�>,��=����!3�G{S���6?�s*?�&��Z���-^=�\M�X��<:�@?���>�T�;
y�>N?��}-���>΁>��>|��>`�>�.��M���H?E?:�(��*v�12�>�������|d=�|=�瑾�H��~�C>X`>�V`����<Zi=;D >%(W?`��>��)����a�����\==��x?��?�,�>�yk?F�B?�٤<c��5�S�g��ow=��W?�)i?Ѹ>#}���оꁧ�r�5?0�e?_�N>�kh������.��V��"?��n?q^?
h���t}�6�����am6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������"�=3���@U�?��~?�������?�6D���&���>�3>1���c�5��OȾ�aP�{B;N��BþG��Ƣ>��@/#R�ӿ�>W������bտ!F���|5�۾g��T?�?�>C<9�T�:�� ��ۆ��Z*�i-y��$-�^G�>F�>u���L�����{��n;��[����>(���>��S��,��ԓ����4<|�>,��>쳆>g(�����Ù?b���<ο����B����X?h�?�o�?�q?��9<��v���{�[��_.G?��s?$Z?L%�w3]���7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�e�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�\�_?�a�;�p���-���ƽ}ۡ>��0��e\��N�����Xe����@y����?K^�?f�?���� #�g6%?�>Z����8Ǿ�<݀�>�(�>R*N>�I_�C�u>����:�i	>���?�~�?Dj?񕏿�����U>�}?�;�>��?/9�=E��>UU�=������5���">��=j<��?�M?��>��=�%9��*/�/eF��_R�/�y�C�]ȇ>e�a?�L?�b>�p���/��� �FE̽��2���+8@�j*���߽�b5>�=>�6>c�C�FUӾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*�ֿg垿� )����2A>g�O>��:>�Eg���1=��=�Px���=���>]^s>�>��S>���>��>��=ZR��r]����eі��v��D����DT����� �����6�X�˾ ����L`=�@V�n(<�zֺ	�_�(9D�m��=@�U?�R?Gp?d� ?�&x�/�>4�����=L$���=D�>�R2?1�L?��*?e��=%���\�d�Zd��6��z���>pI>Br�>:�>b�>4l�9>�I>�?>���>  >�l'=�S�l�=��N>�=�>( �>st�>�C<>��>@ϴ��1��i�h��
w�q̽/�?w���^�J��1���9��ڦ���h�=Fb.?|>���?пg����2H?!���t)��+���>s�0?�cW?'�>%��E�T�>:>����j�A`>�+ ��l���)��%Q>wl?��h>�y>��-��60���O�����>u>5?`[��Gji�fnr���J��=��'>�w�>���Q���ɕ����S]���=u69?t?Պ���ٵ��=v�𺕾[�A>�^>�?=W:�=�6M>/,6����.yN�BG�<q�>��e>E(?I)3> ��=ۦ�>Ꜿ�sU�ӷ�>��L>�->�w>?{�%?f�&��>�������!�{�|>&��>���>s+>�K��<�=�N�>.�a>�׼Mz��$���H��jP>i�z��*b�Qz��~�b=�F��@�>�G�=$����&2�S�O=�~?���&䈿�뾐d���lD?g+?� �=��F<��"�> ��H��>�?g�@m�?o�	�ŢV�:�?�@�?�
�����=�|�>�֫>�ξF�L�ױ?��ŽǢ���	�w)#�]S�?��?�/�Pʋ�Dl�\6>_%?%�ӾQh�>px��Z�������u�N�#=I��>�8H?�V����O�Y>��v
?�?�^�੤���ȿ6|v����>X�?���?d�m��A���@����>;��?�gY?joi>�g۾,`Z����>ѻ@?�R?�>�9�w�'���?�޶?կ�?���>�ޘ?FI?K�/���<�dp��w����t���d��>�P�>pJ�>�A�/�J��Bz���_��e]�b�>M�A=�U�>����Jؾ>�=�2�"�X�p 2>�p�>Ql=PiL>B�>�Kd>�G�>�+�=	�p�ꝋ�M�Ⱦ��K?Ѳ�?:��?+n���<M?�=A�^� 7?G4?��[��Ͼ�Ҩ>~�\?z��?9[?p�>p���3��㿿�{��g�<\�K>&*�>�3�>���mbK>��Ծ<"D�`w�>���>�3��.>ھ�1��j��EG�>{u!?���>�4�=D�?�"*?�I�>��]>��c��,���t�z%�>�t�>!e�>�?__?z���'�}m������~�_�޽��?r?��>BӃ�G槿�5�>�Q>>@e�˝e?TM�?���;�y�>o�?�,?Q%?�ɑ> 9Z�̓վe+½���>7�!?d]��A��0&�ӵ��%?��?���>cՋ���ֽd��4&�������?��[?U0&?�.�H`�K�¾���<�n�A����{<bH�%">�Z>
���T�=��>ρ�=�o��6��b<�l�=�ґ>6��=j�5��5��9=,?`�G�9ۃ�b�=~�r�?xD�t�>cJL>���v�^?�k=��{�����x���U�� �?���?^k�?���"�h��$=?�?P	?�"�>�J��6}޾��ྔQw�~x��w���>���>:�l�Y�'���ř��gF����Ž1�[���>�$�>2�?J��>�Xr>�>p>�q����� ����|G|�^����S�ь)�2���@���wG��ڊ�"#��əf��{�>1gY���W>��?
X�>M��>D��>�A�C��>���=�!U>j��>��0>R�>��= p�=g�N<�2R?b����'��!龴���g�A?�d?Rm�>��]�Na��I���% ?�x�?�Q�?�jv>��g���*��x?��>�l�My
?B�7=%T�E]�<���� ������k��e�>��ؽ:��DM�Ve��
?�}?�ꋼ�ʾ�ڽ��z���=r��?ѣ(?̼I�*�}���}���J�������;��<�����.���W������vB��ѝ>���;�i,?��?2I��v�����9�c�x \���>�O�>��A>�r�>I��>�C!�KT*�Z�F� �2���ݾf2�>��?gK�>_[?>�,?p2D?�C2?��U>��>����#�<M����{>DC>�E?�U?P4T?�J?�FE?� ?��S><�ﾘ�پlb�>�y?��s?̫?% ?Y,�jb��� =�ͽ���mV�Y�w=1&����W=�x��Z��֫>:H?�Y���9������o>?65?��>gH�>֝��E��tt<���>��?��>������l�&2
����>S:�?�$��#=��">���=����d?)�ٚ�=WռƔ=)b���9U�7N7;�K�=*��=����e�q�]�z;��<���;�r�>��?F��>�Q�>�G��ʥ �(��f��=�Y>��R>J>�Mپ}���&��@�g��<y>m�?�q�?M�e=!B�=R��=�t���Q����7
����<��?�<#?�WT?h��?��=?�f#?��>�&��I���\���w�?+!,?h��>���o�ʾv��3�?�?d[?{;a�C��U;)�)�¾�ս_�>�Z/��.~����"D���������}�����?d��?�A���6��x�%���l\��:�C?\"�>�Z�>&�>3�)���g�n%��.;>܌�>LR?�%�>��O?`;{?��[?abT>��8��0��Oҙ��o3���!>�@?ⱁ?��?y?(u�>I�>�)�,྅S��l����7Ⴞ��V=�	Z>���>"(�>&�>@��=��ǽsW��P�>��i�=؏b>y��>���>"�>f�w>�L�<C&I?m\�>�)���8��
���%���L�}z?$��?�\&?�!}=~���?����"��>#�?Vū?hW-?�[M�}��=����px��*�e�u�>�w�>ye�>�=�=>\�>A~�>&�"��K��)��"$��]?��I?�>��ο� ��?�;�@¾�1�=�)v��=R�*#��/����=*�Ӿ�� ��+�����1��$����:x�����x6��OR�>��P=�>���=g��񲽵�i�!.�=�˨=t��<�̏���;�6�<Κ=����iʼ��J:���=�%̼�RȾ�C|?)AH?l*,?Nk@?[�{>�u>��'��,�>F���w?єG>��r�K�¾��7������@����۾��ܾ;ba�����fy>-NA�Q>�<1>
3�=G��<���=&�c=��=ɖ��f�=���=�j�=g��=��=�>�6>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=J����=2>s��=x�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>Me9>��>%lO���-���`�U.^�w[Y�L!?|P8��׾Β�>�֡=<eᾭ�̾
�;=A�0>�>=w���^�au�= ts���M=�Cj=�҆>�:>2'�=k�����=	�T=&.�=hkW>�>G�~�"���%�x=���=��o>J�)>��>�?1S0?�9d?��>�Un�)Ͼ����L�>2��=�b�>�х=�{B>?��> 8?Q�D?Y�K?���>�]�=Y�>��>�z,�c�m�=^�����b]�<���?.��?�ظ>E�O<�B���_>���ýEs?~m1?3�?��>H����J�-���1�S�~���k;�#+=勀�!�9����@0� ��N�>2��>���>�;�>�0�>��6>��A>C��>�R
>�&=W��=;z&�@<~ۼ���=^�F��<Sʼ��9v�	<���h>�0��:p%7���<�^;"��=W��>�<>���>���=����C/>������L�)��=�G���,B��4d�YI~��/��U6�#�B>�:X>%��4����?�Y>�m?>���?DAu?t�>U ���վ�Q��eDe�-WS��ʸ=l�>��<�|z;��Z`��M�-|Ҿ���>��>��>�Nl>=,�q?��iv=�-⾦J5���>iW���Y�WJ��>q��6��$��i�c	�$�D?u>�����=D~?s�I?`ԏ?�n�>iԗ�}vؾ�0>�Ƃ�;�=����p�͸��{?�	'?J��>�����D�Tf̾�0����>�I���O������0�K/�ܡ��/r�>����Ѿ�3��g�������B�[Pr�.�>��O?(�?[b�I���FO�����}��߆?�g?9�>BB?>? 0��1��>V���S�=��n?��?�6�?�\> ��=���F��>x'?$Q�?˒�?nx?�|d����>1W�;��>�Q��R�=z:>qw>�>��?M ?��?�㥽a
��<�$t��M�L�+=���=鎛>���> �l>�9�=\/�=G��=�lE>���>2�[>�mR>���>t>0��'��x6?ގe>?>��Q?a�>>�پ>P�1>A��ֽj�ﾥ�㽉������9��r�">_�I�S�>V����Y�?��C>���fD?hU��{�'>hB�=V�>��,>�O�>�65�d\k>X�>,�>�=vYO>�ۋ>EӾ��>���)#!��'C�dR���Ѿ�z>�j����'�d��(a��b�I�dԵ��D���i��.���1=�'�<�=�?,E��̗k��)��@���N?0�>	6?��������y2>jD�><ƍ>7����{��
����{���?���?S<c><�>��W?��?�1�!3��tZ�A�u��&A�c
e���`��፿����p�
�H��k�_?��x?YwA?��<�:z>���?��%��ҏ�8(�>/��&;�2I<=�(�> (��%�`�'�Ӿ��þ 4��GF>��o? $�?�Z?�OV�)���~�>a1?:�6?���?�=?a�N?�eڽ��$?��)>���>	�?.�7?�?�O	?�?#>��0>��d=��=˝w�/���'�螽u�X�2�����I=b'��=O�<�=�O=�3�mC�h7���t�X)1<j��;���=���=�p�>�$a?0��>�=�>��*?N8.�B!(�����{�?=��<�gc�߰���Ȟ��ƾ5�O>
Km?Z	�?c�a?�>˫H��:�;�>^+�>C�>��o>�>�>I��G���8=J0�=\�>���=�����~����g���g=N�G>��>b�|>�F����'>kb���@z���d>R��
���1T���G���1�9_v�*��>��K?��?�ƚ=T�辘����4f��)?�@<?�JM?��?���=�i۾:�Z�J��D��؟>���<������������:�"�:�us>7ߞ��v����W>y��Ͼ�Wn�&G��Z��=���� =Ŀ���}�|��6�=�9�=�'žf#"��Ֆ�}�����K?�}�=�ꋾ;I�˞ɾ�l>��>�д>6�ża<]�t5����b}5=��>��'>�s��N���G�������>�k@?��9?,mh?n�����}��uB�}n����込��˳?�U�>ǜ�>�Q>.A�=�UԾw�-�z�P�km^�H��>w?��ήb�Λ8�����X0��r�>���>)ҡ>�)?��#?��K?n�j?�!?b�?
f�>/ӽ��$��h;?�ӆ?W�������B��+� �U��=?.�?��}�>h�*?h&f?Lt-? �)?#�?���=����[N�3f[>�>Z�(�3ƕ�R�b>;�A?m��>�1Q?�Ғ?*�=W<��,4���'>�>>��H>�iI?��Y?��@?��>�>f�r��O�=4<?��?L�w?�?M�C�b	�>�B�<*R������j�=Գ?�F?��M?��w?Jn?��>�=w>��0�����.���C�R<CK˽e{��aH�\%��OM=�h�=&���Zΐ�̓�`RR=H=>&�zý���>y�t>� ��60>Ȼľ
Z���b@>;������^���:��=�,�>��?��>�g"����=L�>'D�>B��2(?�?�?X9;��b�w}ھ$�L�G�>�A?�9�='�l��|��T�u��
j=n?�m^?7W�?]����c?��_?0���>�>�ž�'}�����TN??� ?�n:����>f#z?�-t?׷�>)'k�;�k�Bz����b�u�y��&�=g��>D�9c�A�>v�3?���>+#a>�M	>�7پ�w�꫐���?�G�?�Ǭ?��?�7A>T�i�Y�ڿ����Za?É�>󇪾�G#?��V���ž�֘��Ó�q�;����%���
!���ү�f+�D���ac���gj=�?8t?�r?��\?��Se��|a��~���R��G�ԍ�F�B�d�8�tPp�S�����H��lZ7<�š���P���?Cn1?�Ke���	?=���n᤾�۾=��=�A��Z��0A=r_�<:ϵ���<��=��*u��J׾� ?&��>��>��?�~]���K��<�g�4�$߾.� >v��>�P>v�>���;�55��&޽��9,ɾ9�8��<�>�
Q?i�?\�L?�;��9]�}��]�xZ=���k�;��?�jl;�����H��>�Mj��Gj��aG��<��4i�(BO>�	??>6�>��~>2�?��&?5$�o�,���V��p�?�P�6�>U�`?Ħ?F>l�=ĮB���>c�t?���>SK�=k��$��%����X5����>�r?�t?�j�>�tܼ�Bw�/��ҕ�{T8�z�ŽyQ?�tT�Wߎ�t�n>��`?ͽ����[�>����N׾�H�dҽ�+G�>
��>��=N�>����D9�%B�:��h�-?9`?V١�:4���d>?�?dZ�>��>C�?��f>�j¾=�N=�s1?UDS?>�B?�!A?���>�Z�=��\��,�N����=!Z�>�_>X�2�݁(>��y�,�&k8��;ge�<:����;N�6��=��=&�~=A-�=��>��'L�B������[_쾶y���z��.~�d\ھ���jՃ�L��;�r�CU����������w�������J�?�J�?�E=ۜ?�ζ���f�KA�'c>bZ��ӻ$�cSϾ�6���c�M�J�����[,�v�j��*��-�z�-�'?�����ǿİ��99ܾ2! ?1B ?��y?P�6�"��8�� >�F�<���k��W�����ο?����^?���>��@4��w��>���>��X>vHq>���;螾!E�<�?��-?U��>y�r��ɿ3����Ƥ<@��?��@�RA?G�(��!�`rR=���>q�	?��@>�#2����!E�����>e�?��?g�I=gNW��%
�c e?��<��F�F�׻�#�=i$�=�=l���;H>R�>t�^?�s4۽Pj5>��>8�N����^���<JZ>��ڽ�>��2Մ?,{\��f���/��T��3U>��T?+�>�:�=��,?T7H�^}Ͽ�\��*a?�0�?��?�(?+ۿ��ؚ>��ܾ��M?_D6?���>�d&��t����=76�V���l���&V����=J��>M�>̂,�݋���O�*J��(��=����ʿ�!��	-��<�xP�)$��퇽�ý'��<7��9��m��X��o:�=�3>��>z�m>V�>��^?�?й?x��>��������Ⱦ����gy�~��|�"�l.��>������*侨�P8��\Ӿx�ž��<����=�DR�����C� �Bb��%F���.?��$>Mjʾ�M��Q8<<jʾCܪ�Z聼᥽�[̾]a1���m����?��A?�ㅿ�W�`_�t�������W?Ή�x���k�����=:S��/p=*�>��=
I�)a3��KS���3?ax3?�����)��6�>L�7����~6?h#?����=,u>͕?i&=����>���>M��>���>��:>7C��#ֽ,?�^Y?���<������>�D�	n��-5<=�G=��M�BC���=�Y�=�Tݽ?��>b�~�)>��V?���> *�������H�AGB=�Wx?��?�q�>IEk?��B?}4�<	O��uS���
��sr=��W?�i?��>����Uоݧ�D
5?��d?�FN>&"f�8Q��.�����?��n?�B?]���:A}����0"�S6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?r�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>��������==����:�?,H?�������0���UA�'�������3w>�)7��6I��x��L�^r⾁Wξ���p����>�n@�V���?�>ܹ�r1����ؿH<��_�K�cK?�R�>�16���ξ'�b�� ��6:M���;��wh��:�>l\>lk��*���G�{��;�������>n����>��S����������3<T�>=��>���>{������p��?^���+ο8���v���{X?�T�?r��?��?v"@<�v���z������F?_Us?C�Y?�@)�%4^�Д8�&�j?Q_��sU`���4�yHE��U>�"3?�B�>?�-���|=�>���>[g>�#/�v�Ŀ�ٶ�J���:��?Չ�?�o����>e��?�s+?�i�8���[����*�Cr+��<A?2>��>�!�40=��ђ���
?E~0?�z��.�8�_?�a�R�p���-���ƽ�ۡ>��0��e\�DI��R��EXe����|@y����? ^�?@�?��� #�`6%?"�>H����8Ǿ� �<��>�'�>!)N>4E_�\�u>v���:�i	>���?�~�?gj?ᕏ�����<U>��}?�'�>��?�]�=�Z�>0G�=v��*.�Cd#>�!�=��>�˟?��M?[K�>,,�=f�8��!/�G[F�8IR��$��C��>%�a?ȃL?�Bb>j4���2�/!��kͽ�o1�ȱ��K@�Λ,���߽�:5>��=>>��D�Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*�޿"4���վ��awk<ዏ�߁>K��B�p>��4>xz�\_���2M>b�!>I�2>J��>WJ!>��=%��=ۄ�y�"��ה�L��]H�� ��U��v2��M�^t#��������ھ�&��%Ž�큽7ɽ����VT ����=e�U?	R?~p?8� ?"�x��>�����=��#��=�2�>�a2?�L?�*?`��=ᮝ�^�d�_b���>���Ƈ����>�lI>	��>�J�>�"�>F�9̺I>[5?>��>�� >I�'=S�ٺ,w=��N>�M�>���>�|�>	D<>�>ϴ��1��O�h��w��̽
�?с����J��1���8��q����f�=�a.?�z>����>п����x2H?����)�H�+���>V�0?\cW?P�>�����T�c<>���Ťj�ob>�* ��~l�U�)�G&Q>ml?��f> u>�3�248� �P�����h|>e(6?<����:�آu��pH�ؘݾ�L>B��>�0K�u���햿$.�}(i���{=Yg:?]?`G���ư���u�ݧ���^Q>�|\>1H=B۩=E�M>�_��Ž��G���.=�Q�=v�^>j$?,8'>/�=Ϛ�>����J�{q�>�LB>)"/>��??��$?a�����c:��L�)��<v>���>l��>�>�XG�_Ʈ=��>�L]>%�%�����p�*\9���V>�j{���\�v�o�(��=O󎽶_�=*��=�3�� @�� 5=�~?���(䈿��e���lD?T+?_ �=�F<��"�C ���H��F�?q�@m�?��	��V�@�?�@�?��E��=	}�>	׫>�ξ�L��?��Ž5Ǣ�Ɣ	�.)#�iS�?��?��/�Zʋ�=l��6>�^%?��Ӿ`h�> x�|Z�������u���#=���>�8H?�V��3�O��>��v
?�?_�驤���ȿ6|v�|��>M�?���?F�m��A���@����>7��?gY?Yoi>�g۾`Z����>��@?�R?��>�9��'�h�?�޶?կ�?T�>Z�?��?fނ�������'5������Ƚ��>�^?�����*��7��Tɮ��C�����.Y����>��=8��>���$�����=��</+^��\���^�>p�[>i��=�tl>?�?s_�>�=�>�M�=r�k�6�q����L?��?L����n���<�̔=9k���
?��6?9,���ξ�/�>@6b?��?J�X? /�>�	��@���+��#.��{k�<�SM>5W�>���>��� Q>��о��.�fυ>�ܐ>�ǼiJӾ�>���u,:��>o�$?�W�>@��=-!?z\0?g>��O>�T�����a��-X>@��>O�0?τ?�7?�(��I�O�`���&K���9^��*����e?m�?���>��������d��=��9>մ3�4�]?dlr?�=<��>�P?� :?��?�J���"�0�վ�y_�]2�>C�?�Op�Ɵ]��7'�9 <��?��!?�L?ێ�=��:=�A���D�y���F?��_?�|?U1��8��U��=���;�W�<G��;��뼎�>3Q'>���-�>�Y>�ޘ=e���*�/�罓�_�8>n��>��>ۼ��D�.=,?r�G��ۃ���=�r�1xD���>�IL>����^?ll=�	�{�����x��	U�� �?���?Zk�?B��;�h��$=?�?I	?W"�>�J���}޾�ྡPw��}x��w�w�>���>�l���K���ݙ���F��y�Ž"�I��>Y�>'E?�`�>`�L>D?�>_���q'��8�޵���^��e�9d6���.��c������'���3�� ��`|��J�>z���-�>��
?�f>��> ��>�q�*��>qN>�dz>�ר>��[>��8>�L>��^<ίʽZ4R?��i�'�:���4��i%B?tmd?�'�>��f�MP��Ǒ���?�k�?�V�?N�v>6Ch�_ +��d?�j�>P��t=
?R�7=������<4��!d��o��R���Ў>�i׽�9��M��f�f'
?��?�C���Y̾��ս�厾b>�=��t?��%?��B�
�x�/tt�;�R���w��92�͒�<�܃���+�?W]�ˍ���8��N ~��c8�ؿ����3?eٗ?�w!�+^	�|����R���^�L�=pc�>|� ?���>X��>��Ⱦږ\�--B�l�3�JC���>k��?'�>1V?,@?��^?ى[?u��=_?�>�涾�r�>%֣��匾��?;J?p��>��>?��R?_�&?��>ą�> ���7����&?iC?T	?���>g8X?Q�����a�� >s�ڽ@�)��s&��Sh>��2���s���p���">ƞ>��?J���Qo�����d�>|�0?�5!?���>v��Ѐ�=�<=m*�>��>�>P��\�<��U����>�\�?�j��?�����]�=�W>��=��=��>�i�=0Z�=_��~÷�k9f�;��=�ס<H����s=�8�<���=q��>�?ᆂ>�?�>m�~�E��j����=3Y>��U>��>��Ծ����喿]Tc��y>�S�?*��?�@z=���=ƿ�=:У���ž0�������H=�?0%?�@T?T��? �?? %?J"�=.��t���`���n����?n!,?D��>r���ʾ��މ3�D�?>[?j<a����u;)�̏¾��Խۯ>�[/�d/~����CD��G��u��(����?���?�A��6�px�P����\��.�C?�"�>X�>��>{�)���g�%�i1;>;��>R?$�>��O?�:{?��[?�dT>�8�x0���ҙ�`�3���!>@?豁?�?�y?Is�>?�>4�)�#�X������ ߂� W=�Z>5��>�&�>��>h��= �ǽ�C��X ?�-g�= �b>���>���>
�>̆w>�_�<
H?�}�>�.���6��`�������J��Pv?��?g)?Ko=�;�B�V���g��>�U�?yݫ?un*?C�P�py�=N�Ҽވ��]�l�n�>Yٷ>���>+�z=C=J8>�t�>���>���Ɛ��M6�$*��g?�|E?{�=�9���*z�
���D=��]��,���\Y�lg=c�=�ghB=Ս+�[�o��Ѱ��Xͽճ��*ʌ��;���>��S࠾2�>z�;�>w��=/7�=Y��<�?=;��=,d����3���<�Տ;���?�3�'g���p�<�=I�=� <�˾l�}?�<I?��+?��C?��y>�9>��3�,��>&���A?%V>��P�L�����;��������q�ؾRy׾'�c�+˟�OI>�\I�R�>�93> I�=�X�<�=�s=m��=��Q��%=�#�=FN�=h�=?��=��>�U>�6w?T�������4Q�AZ罢�:?�8�>{�=��ƾe@?i�>>�2������lb��-?���?�T�?B�?%ti��d�>K���㎽�q�=t����=2>x��=b�2�V��>��J>���
K��x����4�?��@��??�ዿ̢Ͽ0a/>O�:>��>�VQ�=�.�J�_���f�M{\�30!?�-;���оz��>ax�=�F�ڳǾ�"*="�.>�1=����f^��v�=s+s�*XF=_I^=Q��>��D>�H�=��Н=�j]=:Y�=�PC>4kj;���֮��d7=�]�=��f>��(>N,�>L1?0?� e?��>�h��Ⱦƾ���>�ټ=O��> ?t=�8>rV�>��8?�*F?�3N?�L�>ʕ=���>���>��+�Km���澂���!x�<q�?���?e׺>��@<%�U���';��T��3�?��/?��?`��>������y'�x3��~����Y�4�=B�N��	(;�ص<si����k��=��j>�и>�>�I�>{�>C&>�X�>��>�@=��h=���<�y`=�;�1�=<٫�;ǻ@�=�KJ=�R�N𡽤Γ�10>��)�=ۻ==��<v��=��>B<>��>��=����C/>ø���L�ľ�=�G��,B��4d��I~�8/��V6���B>�:X>���*4����?w�Y>�l?>���?IAu?A�>j���վ�Q���Be��VS��˸=��>M�<��z;��Z`�K�M�<|Ҿw�>��>"��>�]>�M0��-C��N�<�;���*�Z��>r<���k5;����w�*&������ׁj�E��K;? +��Ⲫ=x�z?�&Q?͉?rG�>��*Ծ��4>���P{k�9-�N������#?� (?^�>�P־	wM��̾y\��?M�>7�H�nP�����Ȩ0�r���"��K�>�x���lѾ�13��7������v|B��r��m�>�CO?q�?�?b�0��K@O��dP���S?��g?���>QS?wj?_&�����.���ǹ=��n?��?�#�?N
>z��=h<��vr>S
?�-�?�6�?(�?���!�=)3|�c����c���:���>� �>���>x�*?��C?�:?�d���_�۾)��Q!�}�޾f�=4��<|��>X�>��>A�>�V= �>3{<qD�=%d�Z�z�[Wϼ���=M* �k�R�k?�r>���/�"?yt�=��5>p��X��<G�5>?P־����,>�@��Q��$P2=͔ս�֡�h��>ǿ����{?�O>##�� �!?\�}��iL>���>Ċ>��i����>_�{>-��>C'q>��>gc�>�>�Au>26Ӿ:�>���k`!��/C���R���Ѿ$fz>����u�%����fE��mQI�|���l�9j��.���>=��j�<�E�?�Z����k�4�)�P����?oD�>�6?QЌ�¡���>���>�ԍ>�N�����~Í�ok�V
�?��?�c>��>X�W?��?��.�y�1��Y���u�3�A��e��`�nэ������	��M���`?QYy?d�A?�
�<�z>rU�?��%�E��[5�>Ԩ.�Y�:�;?=�[�>���Pa��xվUDľ?��^G>Q�o?|�?��?$�U�- o��V'>�Q;?�4?��t?�1?�_<?\���#?x�2>�x?��	?�M4?�h/?�
?l6>q��=1q�;E�D=oÒ������Lؽ��Ƚ༭�J=�ـ=�P{�I<�C=.�<[e)� ���2W<p���<��?=$x�=��="��>q7^?�i�>�t�><D9?h~�K"*�Su��1�.?Լ ĝ�gRc�*qv�lI羭�4>,.s?��?��]?]��>�cG�iA�˴2>fٝ>�a>��[>n��>��e���z�A�M=�:>Z�>��=�Mp��s`����\~��|�l<RK>���>_,|>�����'>�u���(z�Q�d>��Q�zȺ���S�\�G���1��}v�WY�>��K?��?��=�W�����Gf�J-)?zZ<?�MM?+�?T�=��۾#�9�Y�J��7���>�m�<��������"��U�:��d�:�s>�-���o��)8]>�	��"ܾn��<J�-?��{i=N�YU=:�
�S�׾.{���=��>>꾾J� �*��������J?�w={ޥ��T��M���>b1�>�ߩ>%7K�w�~���?������J�=�H�>��8>����yA�}�F����24�>x�O?9K?S�c?�ܓ��̈́��GD��s���;�i��Sd�>�k7?k?C#���`�=󅮾_��>�R�(	r���>I��>Po����W��������uT�e`�=��>��<>�E?��5?9W?��?m�E?؉y>�}�>{q�=KT��r�:?5��?(ƛ��D�����-��l�H���r>{�?����8�>�B/?��|?KC?wuG?3��>�>��۾G$B��\>{�>�f�	��0�=>�3?i?X5Q?؜i?;>	����ɨ׽X�>�_>��b?h�\?ei1?%�?L}�>w���ճ��
)?U��?�:z?���?����iR>�`b>ې�<>�
=�W��ٴ?MtH?�?�Kn?�v?1�?�"<��J��?ཋ�����(��)V=�Ƨ=Ɛ=6���f�[������1=GGa<V���u'�=�:>�e<���~�h���u�>2Ot>����`0>S�ľ>����@>̀���
��B񊾡f:�mͷ=#��>��?��>��"����=E��>V,�>%���((?��?�
?��;�b�4�ھd�K�C0�>��A?x��=�l�����Q�u��g=��m?��^?��V�������b?��_?����o{:��%ɾ��t�(���D?J�?G�v^�>�x~?_�r?K�>|���j�������a����R��=a��>���b,O���>�$?m�>�wn>p�=m�۾@�v�_
��Np?;O�?�o�?��?��.>�X�	f߿����ʑ��3a?��>马��^?�?��T���H6���E��N�ؾ�2���-������\밾��"�Y����r�|=��?;;s?��j?�B\?$J��z_�g]��
��U�*��Ҏ�a�@���D��c?�W�n�7��+��i�����<�H��M�I��/�?	�?�ᅾe��>�;��٠e����K>�A�n�����=�����g�D=etV��f�J��7�,?`h�>��>`�(?��V�p9-�u-.�-�5�q��[>�l>=�o>f��>��<���0�M��i�j���g-W��ʢ>��g?d��>U�T?ħ?���b���v���
�Ԏ�>e׺���Q��>�C�>Qɾ)�����&L���i�!�+����N��S����M?!��>���⹪?�i�>pj1��ﾦ;��̾�~=�45>RFv?"9?�a>_����;��=�>�sm?� �>�s�>3я�TU!�k_|�c�彬5�>�3�>���>�?n>�34���^�}���+e��7!<���=T�e?
���3Y��S>8�O?��t;�1'<&ש>����!M ��󾣟)�,*>_�?��=��9>�t���P��gw�G����+?�?���2��F>&�?���>G��>�p�?�yi>X�Ѿ�ϼ&�?f�Q?�G?�L?�V?ko>�<��3ʽ��H��We=���>�/�>.U���V/>SI��e��lA���ʻä>Gnj��]�ϕ"����=�^=�I�;C�}>�����S�显Ly
�����M�ƾ�v���b<c앾���������U�^�l�K�L]���C������S��𫔾�?�]�?_�>]����R��(R�<��n2?C���^ݾ�]7��A����V��ڮ������7#�Bj�[���O�'?�����ǿ񰡿�:ܾ5! ?�A ?6�y?��5�"���8�� ><C�<�,����뾬����ο?�����^?���>��/��j��>إ�>�X>�Hq>����螾n1�<��?4�-?��>��r�0�ɿb���o¤<���?/�@QA?8!�����g=���>	�>��0>V�6�R(�� ��Z��>-ˡ?0��?��<�T�����^?ݎi�� K�֎��N�=ſ�=�Ƞ<D��\�_>�*�>��'�'B�V;ݽ8�N>��>�	 ��|���>�gi"<�wi>�|��/蛽3Մ?+{\��f���/��T��U>��T?�*�>k:�=��,?Y7H�^}Ͽ
�\��*a?�0�?��?�(?.ۿ��ؚ>��ܾ��M?YD6?���>�d&� �t����=�6����x���&V�U��=b��>��>Â,������O�I��a��=���)ƿ��!�.O&�����%;̢���& �-�Žr�	�!i�P�������;��=��9>�oU>�9>g�G>�!V?Ejn?m�?Ë[>�����!��о��+>	B����F�"����M��w,��"��*�r���i��b�r־�-<����=3]R�:8���� ��(c���F��H.?�#'>|^˾��M�#�d<0�Ⱦ�5��-�������J�̾`�1��5n�1i�?�zA?����U�q��UC��Ҹ��.W?-��5��p����=�왼+`=PR�>��=�r���1��T��e4?O!*?6e��[���lN>%�:��tz=�Z?R�?Jd/�Y�u>�?r����h�T6o>誵>��>� �>��B>c������R@?�j?G���9�� }�>��������M���2=�_��#���>
��;L�v���˽�����=�&W?랍>��)�L�2`���*�<B==1�x?U�?�!�>�rk?��B?�v�<vc����S�)�i_w=K�W?�i?N�>�w��z�Ͼ�~����5?��e?<�N>�]h����u�.�JM��?��n?	a?����"k}��������q6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=hz���_�?5pm?x�Ӿ��h���@��f �KȽ��>�	��=�[Q��C0L�����꾠ľ��F����>߂@�%��N�>�}�pxۿW<ɿ��������㿾6!?��?�5�����!�K�T����I�0�E��(�{O�>��>���������{��r;��v��Y�>�����>��S�J������-�4<X�>ר�>ֲ�>9��M콾�Ù?�]��"=ο��������X?Me�?El�?eo?�9<Q�v��{�p7��.G?��s?�Z?PU%�7]���7�%�j?�_��xU`��4�uHE��U>�"3?�B�>T�-�j�|=�>���>g>�#/�y�Ŀ�ٶ�A���Y��?��?�o���>r��?ts+?�i�8���[����*�w�+��<A?�2>���I�!�B0=�UҒ�¼
?V~0?{�f.���_?��a���p���-���ƽޡ>��0��]\����u��Xe����Ay���?A\�?N�?��7�"��6%?��>`���19Ǿ���<�s�>��>�N>r^_�U�u>�p�:��[	>���?�~�? h?T���S����b>�}?�η>��?w�= ��>;��=�z��~&<���!>
��=?EX��� ?B�N?O-�>��=��;�¼-���F��gR�(D	�^�B���>��`?�K?�hf>.����[)��� �� ���7��Iּ�O6��-�w潙r=>61@>��>�D�!}Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*N�`웿�ǾZD򾹝��n#=,� >�3~��=��>��y=q!>E>�R>�+>Wga>|LJ>��=Zk�=��g�#��瘿����UH���`7�"@���a�|MM��ʻ�����k�������e��r	��,���*��ۖ�}��=��U?9R?�p?ˊ ?ةx�؅>����D:=��#���=�<�>|k2?��L?ء*?B��=����b�d�Qa��|>��
Ç�a��>�]I>N~�>�P�>"�>:�A9��I>�??>p��>�� >��'=f�׺у=��N>�M�>���>
��>�E<>͕><ϴ��0��i�h�w�̽@ �?g����J��1��=4��ӣ���U�=�`.?}>����>пp����1H?U���(��+�o�>;�0?�aW?��>���?�T�>>ɷ�(�j�c^>�! ��}l��)�&Q>�j?Swg>�iv>o�3��7��sP�d`���s{>g�5?^����;���u��jG�2ܾ�nI>%
�>+�7����C떿I���h���{=�y:?�?^����֯��w������P>?�Y>��!=~�=�=M>�Xc�Le����G�e\3=[$�=V�\>R?��*><�=�f�>8百��O��>s/C>�=->�??�$?��A����'��V�,��w>��>�0�>��>��I��)�=M�>��a>P��M����(���>��W>��~��^��p��Hy=!h���O�=#Y�=� �� ?�Q�(=��~?<��3䈿7뾡]���kD?�,?�='�F<��"� ���I����?�@rl�?V�	�ޡV���?x@�?������=�z�>�ѫ>lξG�L� �?ƽ�Ƣ�-�	��,#�_R�?p�?!�/�ɋ�5l��7>�`%?��ӾYh�>#x�}Z�������u��#=��>�8H?�V����O�C>��v
?�?_�ߩ����ȿ?|v����>O�?���?T�m��A���@����>.��?�gY?�oi>�g۾E`Z����>Ȼ@?�R?�>�9�F�'���?�޶?į�?���>eҒ?2<?���a���[��.��-O��T�.m]>8H�>�&�<D�E�Q6��C���������g�N��>�k�=���>�H��0���=+�&>��<�'�o��>~B>}�=�sh>�*�>^��>�D>��]>�#��ˬ��p���K?��?��y�m��	�<-ܙ=�~_���?<V4?9Hi�_�Ͼaw�>��\?�~�?)�Z?6�>^�� ���ؿ��O�����<�iK>���>�?�>�|���YL>��Ծ��D��-�>Oz�>�p���پ�Á�~!��頝>�^!?F��>0��=��"?�g5?!��=��M=0�E��
~��`�F0>[��>Br?�\\?��?�㾦�T��,���b����q�A��%�b?��?pv>#��I�T���=�!߽���{�?|��?�d%�QB�>��t?#΃?�^3?"��=[0����%��>����W!?�����B�T�%�����?��?���>黄���ʽ�������g�?\?��$?-����]��������<��/�vb*�X��;񂃼->]�>�]~�Su�=�>u��=�&e��q2���6<���=�W�>�,�=n?��q��1=,?׾G�~ۃ���=��r�>xD���>�IL>����^?ol=��{�����x��	U��? ��?Yk�?O��>�h��$=?�?W	?r"�>�J���}޾3���Pw�"~x��w�c�>���>�l���H���ڙ���F��A�Ž���	�>p��>U?&s ?0UO>}D�>�3��� '�vw�����^�d�x8�V�.���㠾�B#�j��95¾~�{�RD�>�����>#�
?F�g>�{>���>>kлPX�>6NR>I>>f�>3X>�5>��>��<�н=DR?7�����'�ɴ�f���r)B?�ud?22�>f%h��{��J���x?�~�?-n�?�bv>Fqh�<$+��p?;@�>����f
?e`:=�
�ڃ�<7U��a�����a
����>*׽�:�6�L��Qf�bc
?�!?'k��Ϗ̾,׽_�n���>��^?w�
?�Y<�i����A��$7G��5x�$������<�D[��F9���w��V��m3��k킿��:�p(k� �"?p��?� �Z��Q�����I��q;� 4}��3?q�>��>�#G>z��Dk��$��`��i�3�k>��?C"�>�F?��)?�
v?�]I?X�<���>�r��0�?\Њ�&�K��aE>��.?�2f?�aD?��'?��1?y�>
��>O:�"K�:�?�?]Wm?�?�j�>��n�G6�6�>�(p<#���Ѥ�O��="O'>4�ؾ�7�R�(>6yy>��?�ꢾ4�S�=P�� �>�?u?�8�>�G�р��z�?�$��>��>���>��=�G�F�����[�>(�k?�D��J��<u�>@,���	���:�m�����+=��=@���F2���X>*L:>\��;<s�=N���_�=�)����5��t�>��?���>�D�>>>��� �%��Tc�=RY>8 S>�>�Eپ~��P$��S�g�]y>�w�?�z�?��f=[�=ے�=�}���U��������3��<{�?�J#?VXT?Ŗ�?x�=?xi#?��>�,�xM���^��d��4�?4!,?%��>�����ʾ�먿�3�n�?�R?�1a�����>)��Y¾��Խ[`>�V/�"~�3���D�YY��i���i��՘�?���?mpA�Y�6�M�����X��J�C?=:�>1m�>��><�)�t�g��%�N;>��>��Q?c�>�Q?Pw?bNW?{�I>�7��	���xyB�ť>��@?Uӂ?ֵ�??v?A�>ʫ>�s)�G�߾	���.��j�k����=��[>*��>z��>� �><�=0���u^��GO�2�=�s>��>(��>���>Q8p>��=�J?<h�>������⬾�8z�>�U��/k?���?��?��<7�ci1��⾈�>�v�?U��?J*?��M��=1r2�<L���n2��~�>?J�>7�>S�U=(H\=��>�]�>���>�'Q����W:��VU<� ?�G?�V>߰�EZ���x?�h-�̘�kG�=$�ƾ�?�$۾cU�>�٬>����PU���Ľ��.�������þ
�뾏�>�%�=O/�=1�=��=�H���=���<�ˌ��>������N��!j�;���=�=k�]���g++<��]=f�<�˾k�}?<I?��+?6�C?�y>Y:>��3�ؙ�>$���A?bV>��P�؈��"�;����� ��]�ؾNx׾��c�ʟ��H>A`I���>Y83>�H�=HM�<��=s=�=�(R�&=($�=,P�= g�=���=��>�U>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>r��=w�2�T��>��J>���K��B����4�?��@��??�ዿТϿ6a/>��J>)>�Y��V"���W��Σ�cZ�Q?w�1���D�E>h�+>Ə¾ {��m�<x�=>��<�:�PYb�j��=�'n�H��=��?=��>�P>��=1�׽�L+=�E��n>��>�Fݺ�d��a=�eD=݋�=,�a>%��=���>�	?�(0?�d?�8�>[vm���ξX��(x�>�\�=>�>l�=�C>eø>�8?ͳD?��K?`��>�<�=nƺ>쿦>Ny,��m���<����´<�x�?���?޸>u�S<�A�����_>���ƽ�g?��1?�?$��>�	���߿�&�672�i8��'�Q�U�<{y���6b�J��P4��s���C�=;��> Ľ>n+�>�}g>r0>�G>�A�>��>%��=�c�=Lj<��P=���}U>��߼r��;6����>�Wԏ9������8�Q�����	��#�:΁�;��=���>M9>Ŭ�>���=�	���B/>縖�{�L�=�H��:+B��3d��I~�P/�kV6�g�B>L8X>�����3����?��Y>l?>p��?�@u?�>�!���վ�Q���Be�SS�ɸ=h�>��<�z;�PZ`�8�M�|Ҿ�'�>G��>2��>�j>(,�?���n=m3�ؔ4����>�t���w�?^�Kqq�5��<џ��;i� 2���?D?�������=�e}?a�I?���?�T�>;7���\׾T2>�Ђ��Z=�h�m�6*���?y'?���>4q��CE�̾b���>�FI��P�q���.�0��Q��ڷ��s�>{ɪ�Ѿ1 3�Pa��� ���{B��Qr�]��>�~O?m�?�b�0���'O���+k���F?��g?�#�>K?';?����p>�7����=K�n?��?�.�?[O
>];>�A�:>ʉ(?�Q�?���?�f�?dFI���>ކW>�E��&�������>t��>�>��?�+?}�?�i���	�i�
�c����?M<3�=�l�><�>�>��>|"�<ظ�8ST=��ؽ�󊽂f��ok>��G>�"ྶ]�_GI?�>�=�.�=x2?#�>�_n>5	�$|�=2��=V@���c��Y��T���d=gȽ���/�E2�h��>~c¿�?�5>Ɏ込�?�����ۼiXV>�>c�(<���>/I>��>���>`q�>a�=�-�>��>>��Ҿq8>���!��0C���R��#Ҿfey>�����%�Rf��E��h�I����<���Dj�N9���d=�ֿ<0�?0���[�k�M$*�@a��'�?�x�>��5?�o��ꇽ�+>�]�>�D�>(K��(�������n��vҋ?���?�;c>��>B�W?-�?N�1��3��uZ��u��(A�e�J�`��፿������
����&�_?�x?*yA?�Q�<6:z>C��?��%�@ӏ��)�>�/�';��=<=,+�>?*��h�`�:�Ӿ��þ)8��HF>]�o?1%�?=Y?�TV���i�О&>�:?
�1?ܫt?��1?.�;?���g$?*4>G�?]b?j�4?L�.?�*?�N1>�$�=p���8=�|���
��H�ҽůͽ��(:;=u�=R��,<��=��<n&�o�c;T����I�<�A=�
�=//�=4m�>�b?�m�>���>�q&?�}[��{�5ۛ���.?\Z�yW���|x�{T�Zm���6>���?�w�?�W?@��>aTJ��-s�'>>�R�>s��>�)>��>c�����m���]���|=�5>?�i=`p�<B�t��,��%q��r?a=ygf>U��>p�|>Pn��n>,>�젾�"z�D%f>5,Q�5B����Q�{tH���1��kt�K��>D(L?�q?���=�羿���E�e� �'?
.;?��L?�,�?���=R*ھ"�9�tKK�8��͡>V�<�,	��Ƣ�z���e�:�9�,;��s>ٞ��짾�V<>�|���`��7�t�WPC�D���={���>� ��I���Z���s�;m>+ډ�k��K��_.����Q?���=VO;�������`>Qh�>H �>�T)������� �@ű�|�=8��>��>�gصv� �@q^�������>��W?QAI?�zc?��G�lE��S���Fm����?��>�
?SE>V�u<�r�-*�73`��X��>^k�>�f#�\�5��wk�s8�� �ۑ�>�F�>���=m@?��#?B��>�o?��-? �,?gڹ>؉�oᾣ�=?`�?�n}<�o+�������#�#*E�B~?��>�+���?WC�>�_?�-!?�:P?T@�>WБ=.����P��R>��>ϓD��� �>}H?2��>v�C?��|?���>'$2��.�+��Bo=�&�>`{S?�@?
,?���>�F�>���D��=U��>�?��l?��w?ZM>���>�\N�{Я>�Ɏ=��?�3?�~	?��L?�ut?��l?9��>��=�h�A���Xý?_���=�l�=yL�<!)���l=����ja���=�G=ܙ�=�l/>hcｦݘ=&?��]�>��s>�����0>��ľ9S����@>@����M���Ҋ��:���=؆�>@�?ު�>�a#����=ڭ�>~A�>���V5(?�?�?�";2�b���ھa�K���>eB??��=��l�9���N�u��g=��m?��^?ڡW�&��t�`?\�]?N~�I'3�͔þ�7}�fo��1oM? ��>�����>�7w?޸v?��>��m��}v������8[��f���=@K�>��
���]�7�>�s8?�?�>_�5>�= �۾�3x��m����?�6�?�?}�? a>"l��޿����qq���@\?U��>+���'�?wo��;����녾O���f��S��������������_��M��b�=`p?{�s?�{r?�_?Y!����_�D6[��~�V�W����M�oXE��LC�+4C�%�m�C��� �j좾��=��Y�p�>�S^�?/x3?Ʋy���>�"9�ݲپb�꾱�>�'���T���N!�c����;=F@W>������꾖��S%?:�z>k��>ku(?K��e���8=����#t�Z������>���>=��>R�>��U���;�%<��SF��OJ��8�>N�c??G?xf?�B	��w2����� �����~����Q>��>��>sM��	�+���3��pD�ؚj��q��G��,���Cc�=�A(?Z>-۪>�5�?�6�>c�2���s����Z4����<�>c�g?�>�<�>m2���*�F�
?8�y? ��>�3�>��⾢I��ߕ���>K��>菷>�?���>2���D��W⫿�]���_�� m=�>�?.c��(x�z��=�dA?�D�=�{P=}�>�w���K�c*)���ýf${��2??nr�=���>�Q������(�T��V���*?��?Vv��,�+��6�>�9?4��>�P�>���?r��>8���Q��;e�?m	]?p�J?s�A?p��>�`D=�����Ž�q"��,=wU�>��H>��^=z�=��%��5N�!��g�<��=d/��$ɽX_<<��Ӽ���<x�L=�SA>3�ֿxxN��4ؾ�T�3�
�ȭ��r��ƽ��1�ZΦ���Ծ�9���^���J(�k%׼l��#�����:v����?%�?%�g�}/T��L���8o��[��#��>E5�$r�=���=�ٗ������@2���o��VG���n�-�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >[C�<	-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾u1�<��?7�-?��>Ŏr�1�ɿc���}¤<���?0�@�??A'�	3��X�=�L?��?��[>����c$�i�澒�>��?p�?�=��P��ة�\�h?���=+X6��J�</�="~�=�f<�(:���y>7�>?�#��
k�ｾP>���>�/<Z��~%*�?Pp=�<5>�����֍�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�'鿭��_3��=sv�����?�>�D>���J^>���=F��	���>�=�>���>A��>�7�>e��>�'!?q�1? K�>�K�>aڝ�M����߾���=�Y���S����*,�������2о;���D4�j�{a;{ >���	=�J��M����.��a�5��*?��e>ك���Z��=J��t߾Eļ��#�V���ȭ�K�0���m����?3�J?p��@�3n��������O?|��I�x髾��t=9*�=1¼�,�>��=� ���G���\�w9=?�@?�٨��䥾��6>(�U��+v=E0?�:�>��=���>ՊE?� ڽ@����~�>$U;>�^�>��?�� >�⤾N ��j)?U\?T�x��d�����>������:�=Ǫ��2��<�~-��5�=|����Ͼ	�$>KRu=H �=yW?�s�>�)� ������5�\>=w�x?/_?-T�>�_k?P�B?C��<v���y�S����ky=��W?�-i?�	>.��.�Ͼ㈧� l5?ۭe?-O>Wh����.�
L��&?G�n?�z?|ޙ�!B}�������h\6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������>lέ����?+��?op���Q�;�Q��zR��W��Ow�/<>��
�3��^J̾-�1�ew��qT��P��Ž��>H/@���꽖>CA����iտ���鮾9����>R��>M �o���}��K��v�_��-�z��V��>7�>�Õ�����y+|�0r;��;���t�>����쀉>/�U�]����T����%<�֒>���>7h�>Rw�����պ�?����+�Ϳ'-��(��{^X??��?�z�?�w?s�}<�Tx��}��(�K$F?f&s?WZ?�R'��_��E?�'�j?_��:U`��4�xHE��U>�"3?�C�>��-�ر|=�>��>|f>�#/���Ŀ�ٶ�����F��?��?~o���>[��?ss+?�i��7��z[��z�*� �+��<A?g2>4���"�!�E0=�gҒ���
?w~0?q{�C.�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�#N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�O�>��?u�=��>��=s���u��n�%>X1�=<r�A�?)L?���>N��=]:�.�1���F�CQ����B�` �>F�`?�{J?QKh>ť�jI(�'""���ʽq�8�����F��G@�)5˽ �5>z?>5�&>Y�K��u־��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ua~����7�b��=��7?�0��z>���>��=�nv�ݻ��W�s����>�B�?�{�?��>"�l?��o�N�B���1=4M�>͜k?�s?�Oo���t�B>��?"������L��f?�
@~u@`�^?):��������0�a־4ug>=��>MX�>�u6��`��9>����3��=�>�>O�>�	�>��*>Yn|>M��>�^��D�I̿X԰�hO�����"۪�착�0�����!�������Z�=_>?�F{��6���f�=?�=��U?�R?,p?�� ?�{w�p�>����V�=o�#�CO�=-�>�d2?��L?��*?7��=ؓ����d�{b���3���Շ��_�>�6I>���>b(�>�"�>��#:��I>;�>>5|�>�� > (=(�˺��=� O>>3�>M��>R|�>�B<>$�>ϴ��1����h�3w�̽� �?”���J��1��[:��b���e�=b.?[}>���	?пq����2H?[����(�M�+��>��0?�cW?Y�>����T�U;>����j��_>�+ ��~l�a�)��"Q>�k?��d>is>��3��P8���P�l���|>�5?W�����9�"�u�-�H���ݾsM>���>#>����ޖ�8�~�0�h���z=s�:?)v?/=������fw�c���@R>>,[>�=��=��M>��e��Mɽ��G��.==��=�]>��?�1>?��=H;�>�P���R���>�?>b�)>m3@?r$?c���ܐ�?����w*�*�q>�n�>��>�5>�J���=P�>{�d>�q��FXu����{C���W>y�w�?�]�	�}���x=�ɕ�	�=���="���?��=�~?���$䈿�뾠d���lD?V+?� �=5�F<��"�@ ���H��H�?q�@m�?��	�ѢV�H�?�@�?�
��^��=}�>�֫>�ξ�L��?��Ž?Ǣ�Ĕ	�7)#�fS�?��?�/�Rʋ�-l�d6>�^%?��ӾWh�>Ux�~Z�������u���#=2��>�8H?�V����O�M>�w
?�?�^�䩤���ȿ;|v����>Y�?���?_�m��A���@����>6��?�gY?�oi>�g۾4`Z����>ϻ@?�R?��>�9���'���?�޶?կ�?��P>>�?�r?¡�>$v�A�.��,�����<�K=먆<̩�>�� >豾��F��	��U���i����*IS>��2=�*�>%f۽3����k�=T�A������ܟ�X>�>b7U>�=>���>X�>�t�>�>/�B=6r��և�A/���"L?Ώ?���yn�%K�<E�=)�_�UR?QW3?B�F�8;ZШ>d�\?Љ�?�[?m�>�x���������'���К<�6J>���>���>F����M>3վ�FA�[Q�>�3�>� v�@�پ|���8��B�>��!?���>Њ�=�\%?߄:?�(�>.a\>�";�-ї���z��+?oQ?��>�B}?^�3?(뾶dQ�pت�R6��uj��"�G>�D�?[�?���>�v�dԐ�����+�<߰%�w��?(��?f�y�y �>�2�?=Z?۔?��D��M0�b\
>�L�>��!?ae��A��H&���d?�(?���>�����ս�м���<����??$\?M:&?T���a�Y!þt4�<��!��S`��Z�;/D�q|>��>�u����=">F�=X�l��M6��6e<|Ҽ=$��>��=�6��_��1;,?��G��ڃ�4�=}�r�)xD���>�IL>k���Э^?�v=���{�����x��wU��?B��?�i�?����h��%=?b�?*
?�#�>�G��{z޾}��Ww��{x�`v���>���>�l�m���������G���ƽ�F��o�>�z�>�@?�e�>�OO>H�>#���''�s��x����^���bm8��R.����ؔ��qN'�{���{���s|�Eb�>s@����>N-?�xe>5�y>���>Gt�]�>{Q>��~>��>7�W>[P5>#��=��;��ѽ.5R?
����l'�����뮾��A?�sd?m�>�r�D䅿���*?[��?ᑜ?N�u>��g�@r*���?Dc�>4�~�ve
?'<=�����{<����1��懽-��}��>�mؽK�9��RL��=d��
?�n?����˾|j׽x�[�hK�=*_�?�?\Z�x�k���z���Q�+P�jf�B��H���܃(��!z������Jz�����}K���=�� ?�ԝ?d���7��z��~}��Mu���>��?Oɢ>K�>+2�>�h辨'O���v�iY��ž��4?���?���>(�I?��??��L?¢;?`��>
ٿ>2�W��>2�Y>��>�{/?q�7?(�>W�?^�>��??\E�>Fn��������u?��>?X�;?��8?��>oX���r�=������=�Ye��A=[X�=�"���"�s�=��J�'��=�Y?���$�8�y���C^k>�v7?���>���>17���m��y��<���>�
?Io�>L���Ohr��K�J|�>I��?�{���=]�)>Z��=Hˆ�f������=YJ¼���=���$�;��d < п=�I�=a#h��������:�\�;Y8�< u�>7�?���>�C�>�@��/� �b���e�=�Y>AS>}>�Eپ�}���$��u�g��]y>�w�?�z�?ܻf=��=��=}���U�����F������<�??J#?)XT?`��?z�=?_j#?͵>+�jM���^�������?l!,?��>~��z�ʾ��̉3�͝?e[?~<a�ո��;)���¾o�Խ[�>�[/�M/~����GD�����������0��?濝?rA�3�6��x�ο��\��\�C?$"�>�X�>��>6�)�i�g�j%�]1;>���>TR?�~�>�UP?�Zz?I_Z?��R>8��ԭ�����t��o`$>M??ж�?r�?qGv?��>�P>�,��aྻ���J4����9���sO=�,^>���>���>��>��=/�׽Sk��q�B��o�=ϥh>���>ѽ�>η�>�q>�q<lH?)^�>Y�����;!���郾��B��Yu?1�?ƅ+?�l=����D�������>�@�??{�?/*?�2T��'�=��Ӽ#���͎q�$@�>�>���>j��=x�M=	�>��>�$�>���bc�{�7���O��d?�~F?�'�=�~ſ��x�!���������������K�,�N�z���
(=,�Ⱦ�6w���ľQB;�ѝ�#H��s�&1��-k�vy�>\v=|:*>hu>Ob�\"�T��<��	<6�=���=��̽���<Yވ�o�������<���<�n�=B�2<ۈ˾t�}?�;I?`�+?��C?~�y>�<>�3�@��>ᅂ��@?4V>}�P����a�;�����[��3�ؾ�w׾��c��ʟ��H>�UI�{�>�;3>oH�=�B�<��=�s=���=1>R��=�'�=rN�=,g�=S��=�>�T>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��=>X�>��Q��n1��V��9c��^���!?Mo;��0ʾ��>���=�۾E\þE�C=.8>�^=P���6\�=�:t��k/=�Z=�}�>��?>08�=�u���:�=X�M=�=�jW>z�λ�*>�y���+C=���=�i>T?+>	��>�!?s'0?�d?�O�>0n��MϾ����1}�>t�=z��>B�=��B>7��>��7?e�D?l�K?'y�>k�=Sߺ>���>͎,�٢m���$ݧ���<Ň�?���?��>E'L<��@�Y���->��ý�?�71?W�?7�>H���տ�-3�=5���C��i�^~�<4��%'�<�B��A���BX��Q�;0v�>9��>m��>hΘ>>�>�ر>6v�=���=��>���5n.���k�ls}�φ<;=:�7��s�<��	<��½e/ӽJ�b<�P<b�L=;��<�9�=�(�>�
>�.�>bɐ=?ҳ���0>�ߖ�"L���=ܨ���B�+xd�k�~��.��3��A>�R>�ю��g����?�^>��A>wz�?.�u?��>�0���׾�H���``�S���=q!
>3�<�e�:�ټa�U�N�PZӾ���>���>���>NPl>�K*��?��<=��־��5���>dA��Ŵ�+��Ƀr������p����j�JN�P�??|Ӆ� 6�=E�z?��D?�p�?���>m�x�+߾Yd)>�ԅ�l�X<�.��i�5$K���?��$?�� ?9��;)H���;��Ž܎�>;�H��FP�_���H0���N��K�����>kث��[Ѿ�B3����t����A�(/o���>'�N?��?}C`�����N�?���+���w?�h?A֡>��? 	?fˤ�� ������Ӻ=�o?qK�?ɣ�?�b
>�x�=>��B��>��?���?]z�?�s?#|��:�>1�8>��\�F�D>Le>�W�=Oz�=x�?��?�Z?˜Z�^P�*��ٶ�QU���^�=��=���>V^S>��H>�G�=뽒=�q>~|�>W�>f�>q�*>�ĥ>v�z>�՘����;�.?xw9>AT>I�/?Ȩ�>f]=����{=��s��H��g�H�m�ӽ�������=*p���UݽÌ.�(}�>Q�Ŀ��?U>�Fپ� ?�����M��2�=�
>m=��>-�d>��>3�>�@�>��=3�U>v�M>QCӾJ�>����c!�b,C�@�R���ѾVyz>V���T&�M��Ur���EI��r���i�j�|/��P<=��<�G�?Š��U�k���)�I���-�?T�>�6?�Ҍ�����ȵ>���>Jō>�J�������ȍ��f�B�?R��?�;c>��>>�W?�?ؒ1�?3� vZ�#�u�f(A�e�J�`��፿ �����
�����_?��x?yA?"Q�<S:z>M��?��%�Kӏ��)�>�/�';�a?<=e+�>!*����`���Ӿ��þ�7��HF>��o?<%�?`Y?lTV��Z�<肺<��??cPn?���?�l?�2R?�T���m9?�m���>��>?lOH?��P?}��>�b�<���>����q��F�a ;�0Z���D�<�s�� �=�qK>��=�.���e���,�>1�M>���<}w>
6̼��J=�u�<�X�>�]?I�>�e�>�i7?T��Ģ7�����ȡ.?4�C=k����Έ�X���;��>9+j?�̫?�Z?b�d>Q�B�>�C���>�ً>�E&>|�]>��>9�w7D�#h�=��>9a>〉=�8Q��˂�~�	����gm�<*�>���>�|>�荽��'>Ä��-z�N�d>}�Q��Ǻ�D�S���G���1���v�}F�>��K?b�?ᄙ=�p龅��� <f��.)?�b<?UNM?��?�7�=��۾��9��J��T�%�>�4�<��W���� ���:��W|:�s>u5���ɒ�H%v>"X�7�о�Pq�jQ���㾏�=�g��c�=#�{O뾠����X�=A��=�!Ѿ9� �Ă���ǩ��}F?4P~=�����[�@���{0>#q�>���>a.}���,�:������
=��>҉<>.B�<p�ྣv@�U�䙙>�H?-W?��{?I2��‿�<���r�־���<�e�>��Z>��>�>���<=�ʾgK���o��X��(�>��>	\"�ʸP��y�_)ܾ'���Z�>��>#�=g�#?S�W?���>U�F??�*?�?<��>�u�<��پ�:?,�?_�o�����{��6F��)�~F?!��>���@��>9z�>��>|��>��H?��?�}>ミ��bm�7�a>���>2�L��۳�uY$?�u\?8<�>��}?o.�?�k>�C���V�I��=�0M>�,�>[M?��0?�A?J9?��>\��X����-7?�]{?��?-��?��8�ν�>D[���L�o����b>R��>�Y
?��o?ee?�[?�u�>�T�=Ƒ-�v����u;(ؤ��߰�*E	�)Һ`.�zL�<��G��=>]�S>=RS>�c�=�+��T��r��<�a�>x�s>^	��5�0>��ľ�L��>�@>�x��<H��&ӊ���:����=q~�>��?ᮕ>HL#���=Q��>|O�>����2(?��?�?��";A�b���ھ�K���>B?e��=8�l������u���g=�m?�^?&�W����I�b?�]?h��=�Y�þ&�b�ɉ�O�O?�
?d�G���>f�~?O�q?��>��e�D:n�#��Db��j� Ѷ=<r�>1X�$�d��?�>I�7?O�>��b>$�=nu۾�w��q��(?��?�?���?�+*>��n�N4�ed�Ň��܃~?Y�>	\����\?�&����q���F��=����վ/���^��y���Y��#��ǣ9��˄=*�?V?��?c�E?Ѿ~A,�z�B�G��C�Z�)�$��W��#��B���a���q�T���� �(\ƾ�Ĵ�����P:S�~��?�(?�a��b7?����o����鸾G`��k޽��_���<!���1��#+=@٧�����ݽ�# ?{W�>�6�>�3?�U�>:�~{.�[1E��f���[=��>�Ԝ>��>1�5�޲,�P*������D���Wi�a�>�Uc? bH?�h?E�M��%<�q�|�'���սR ��p�>�MM=�9�>|#u���H�f(5��=��|��x�{C������=��.?���>~e�>���?��>���^���0_����8��������>7f^?��>�q�>bT&�i4+����>p}?U��>7dq=m�<*��:����=^�?��?���>!6�>��*>�>��Dp��ݗ���j�1->�w?�k�!D��wp�>�S}?0P���e%?>�=Tlk�&kʾ��&��:�����>�3>>#�־Q����p��ȶ�ѱ.?g�?$���ց?�va�>��?6�>!M�>�t?[n�>����y^�=�?7nJ?w�P?&�A?��>�B�=LA���#꽻��>�5=j܂>�b�>���=�h�=�ds���2�����;{�=�����Y��C���<F�,q>mL�;���>lۿhDK�וپG�?�~9
�>舾&����Y������S��V��UGx�yu�$�&�!V�7c�D����l����?b9�?Uk���'���������h������>�q�~���﫾a�T,�����-Ĭ��]!�7�O��&i��e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >`C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���z¤<���?0�@�A?:�(��r���g=)��>�	?�(C>�2���&�����>��?��?HX=C�V�4cݼ��e?Ƈ(<(�E���û��=3z�=�
=���KI>�h�>3�~C@��uϽ��6>�R�>�i��j�,!`�H��<�>]>sν
:��5Մ?,{\��f���/��T��U>��T? +�>W:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=q6����y���&V�y��=Y��>c�>��,�����O��I��V��=����tDÿcY�M��d .<+��<��d�.�ƽ޷t�R���C�u��{l�@�N�3F>k�>��>ff{>�2s>\؊>�Y?�Z?�]�>�J>v�:�w?��c�~�h=�[�w�4��:b��}N�{��yѾ���U�, ���Ѿ��<�Ĵ�=*%R�P���&� ��b�I�F���.?��#>��ʾ�M�!)<��ʾHժ��8���@���*̾G�1��;n�9ş?<�A?{���XW�p��*��}N���W?3��������Q�=�_����=�M�>�ϣ=�~���2�{S�W�2?lDA?�}���*��@�>`ֽ�ݬ�<�	?\��>�K8>��>e�A?K���m˽A�>�5k>V+?%��>�ع>Qeʾ�A��9?�f?A���NN�ĩ�>6"��R��i�=��>�6�`2�q�=�
�g$e�C?>0#K�;	#>�%W?�O�>��)��h�-ϐ�<����3=Yqx?;?�͠>�1k?�jC?�5�<~T���:T��R�|4p=��W?�@i?��>=����Ͼ즾95?+le?U�O>pf�Mj�9�.��U��/?�n?*?K+��y}�%��Ɖ�(�6?��v? s^�ts������V�Z=�>\�>���>��9��k�>��>?�#��G������lY4�#Þ?��@���?]�;<��j��=�;?o\�>�O��>ƾ�z�������q=�"�>	���^ev�����Q,�h�8?ޠ�?{��>)���������=Y�����?q��?c�Ҿ�&>����.s����)z?�*>_>�Ll��q�v�ؾy�1�=W��������� c� �>��@v�(�Q��>����j��/ȿ7�l��"�$��sh�>��>
>�/��	LU��%n��3�c�M�2���	�>��+>����R���g}�dA�� ����>�����>�5/��7���Ϋ�*����>���>��>��ƽ.`ھ��?5�쾉�ͿQG�����ȂW?��?��?{t?�;�C�tIT���;�9@?�xx?��b?	�5<Y��J��j?�^��7U`��4��HE�pU>b"3?FC�>�-���|=>���>�h>$/�y�Ŀ�ٶ�����7��?ˉ�?�o�k��>W��?�s+?�i�8��NZ��m�*��|.��<A?]2>P���G�!��/=��ђ�a�
?�~0?k|��.��_?�a�7�p���-���ƽ/١>=�0��i\��G�����tZe���1>y���?7]�?��?����"�R4%?:�>n���d8Ǿ�	�<~�>$(�>J(N>}>_���u>w���:��q	>��?0~�?�i?��������+J>��}?�$�>��?$o�=�`�>Qf�=���-�-j#>�%�=��>�B�?˨M?xJ�>�U�=��8��/�ZF�DGR�D#�/�C�N�>��a?;�L?JKb>=��2��!��rͽ�b1�(4�=X@�r�,�g�߽8&5>��=>>��D�FӾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ta~����7�N��=��7?�0�'�z>���>��=�nv�ݻ��U�s����>�B�?�{�?���>�l?��o�S�B���1=EM�>͜k?�s?�Eo���`�B>��?������L��f?�
@~u@g�^?'d�ѿ!�������Ⱦ�]>��=}$7>~�ٽ��-������=a<�N=�����U�>���>n$F>dL>�>o�>]<��U� �c�������4k����� ��+����$n���#��(���qQ����R�!��Z����)b�����5��=i~U?�R?�1p?j� ?)^q��c >����ݧ=��#���=H��>M"2?��L?��*?�ݔ=p�����d��W���H��oB����>�WI>,]�>t��>H�>�Qy���I>�?>���>EW >��%=�	*�I�
=Q�M>�$�>�]�>�ȹ>�C<>>Bϴ��1��l�h�w�z̽.�?����K�J��1���9��ݦ���h�=Bb.?|>���?пh����2H?���~)��+���>|�0?�cW?D�>���T�T:> ����j�-`>�+ �Ql���)��%Q>ql?��f>�6u>�3�}X8���P�h���X|>"'6?����9���u�3�H�`kݾ�3M>ܪ�>&�G��k�S ����>`i���{=�l:?yz?�ܲ��ݰ��u�kI���.R>�\>�f=�i�=�M>��b��ƽ��G�y�.=���=ka^>�>?p=3>C�=I\�>{����M�>��>�68>��3>�@?5�&?nx�1Y�����(���{>��>�ր>��>�M�e��=>�>#l>�D�\���ܣ��,A�eyV>
jp�,mZ�p����=�t�����=��=�� �jv>�PY=�~?���(䈿���d���lD?T+?S �=ҝF<��"�E ���H��F�?q�@m�?��	�ܢV�?�?�@�?��@��=}�>׫>�ξ�L��?��Ž6Ǣ�Ĕ	�$)#�iS�?��?��/�Zʋ�<l��6>�^%?��Ӿ�h�>qu�:Z�������u��#=��>]8H?�S��1�O��>��w
?~?�`�(�����ȿ�|v����>A�?q��?�m�LA��#@���>��?�gY?�qi> g۾,`Z����>޻@?sR?:�>I9���'���?�޶?ޯ�?��Y>6��?�op?͉�>vӽf�8�o������ks.<VY=��T>Y�=�]ƾC�� ���R��z�h�"$��99>��G=Y�>P#���_��l��=�����X��-��`�>�X>iD>a>�>!{�>��>.��>*ʨ=��L�̄n����YL?��?���Aan�p��<Dk�=`�^�.�?d$4?�S��оy�><�\?K��?�[?(��>������7ο�)w��Cw�<��K>���>���>!ˇ�]�J>�վ�C��\�>y=�>ߞ�(ھ����{���o(�>�!?A��>��='� ?A�H?�w>/��e{T�m����È����=��?��E?��?��*?�� ��i�&�㙨�`��h7�=�CW?�|?�B�>۹��\᏿�.<x=9=�͋���n?�ڏ?
�=�η>c�?�s?��>]1�<��Ւ���G_>@��>v�?��h A�׳�<�彷'	?h�
?�Z�>ݯE�����ؼ���rU�y�?��^?2')?;�O�Z�?!��=��;7<�s�%���ؼҢ>{t(>�w����=@5>�C�=�"��W`�Y�i<��=�w>ܩ=�&�-�|�.=,?��G��ۃ�k�=f�r�6xD���>�IL>����^?�l=��{�����x���U�� �?���?\k�?���+�h��$=?�?R	?S"�>�J���}޾,�ྸPw�1~x��w���>���>��l���4���ԙ���F��K�Ž����>��>4?(  ?2�L>�,�>Fx��Yc'����9c��_�w�y18�L�.�̲�+����$�>��r����{����>ME���R�>e[
?��g>%�z>&T�>�K뻯B�>V�R>�~>
��>^X>�f7>)�>ʠ< Խ�KR?����8�'�j�辈���"3B?�qd?n1�>�i�������\�?n��?,s�?^?v>~h�X,+��n?{>�>���Mq
?S:=B�~4�<�U��S���2��i�r��>�B׽� :��M��lf��j
?/?d��m�̾�;׽�M�r7>Rm�?t��>��P���S�
�F�k�|�l���������M����N�3��c���D�������p�lO��O)?�O�?>>3�j�E�������n� l��J�M>���>B ?"&�>�d>�C�f5C�.Zh�gR�S�����?\�x?$��>��??�~H?$7C?�f^?�*�>�}�>��پ�?�=fŕ>�(?H��>X�>l2'?90?G?���=���<�_��;�\�
?�r3?��6?{�?��&?�f:��l'��Vz��0���a�L��*ْ>sp�=:��ڦj�{����н�Y?���8�<����k>�|7?߉�>���>@���'���v�<��>ų
?H�>c���	rr�Y��b�>l��?n��_�=��)>���=������Ժ�G�=�3¼p �=/y��!�;��d<g��=��=R.q��v�����:���;�y�<u�>�?���>�C�>T@��)� �:��Te�=�Y>�S>�>Fپ�}���$��S�g�^y>�w�?�z�?��f=��=��=}��^U�����M������<�?+J#?XT?N��?��=?dj#?�>�*�JM���^������?w!,?#��>�����ʾ���3�ŝ?^[?�<a�����;)��¾��Խ}�>�[/�y/~����OD��򅻴��Y��'��?保?5A�P�6��x�ٿ���[��^�C?�!�>�X�>8�>$�)�f�g�Y%�2;>���>;R?�#�>_�O?j<{?��[?hT>G�8�-1���ә�NB3���!>�@?᱁?��?"y?�t�>��>��)���9T�������Ⴞ�W=W	Z>b��>�(�>�>e��=-ȽZ����>��`�=g�b><��>���>C�>p�w>qC�<�I?	��>��ľFk�w�� ���E	g�*u�?{��?�b+?��ܻk��pe;����-�>(�?<P�?�.?2.V��$�=Y������%y�C.�>�e�>�t�>��H=���=�>$��>���>�����
��13���K���?-�B?�>�ƿ\�q��r�|����6_<V����d����Y�è�=�ߗ�Ӝ�����X�r���V��\���i��qy�8 �>�^�= q�=�=,��<�˳��̮<9M=�i�<-9=�(k��@Q<��:�ļ��1D��y����G<��F=E��+�˾A�}?�;I?[�+?D�C?ؾy>�=>B�3����>����@?�V>k�P�������;���������ؾtx׾��c��˟�jF>�\I�L�>�;3>�K�=lF�<��=�s=�Ǝ=��R�>=*�=}M�=:`�=$��=^�>HQ>@6w?񚁿Ҳ��<2Q��O�y�:?�:�>:t�=��ƾD@?u�>>c2������a��-?��?�T�?��?�ui��d�>I���厽�s�=���H<2>��=\�2�6��>��J>���I���w��"4�?<�@i�??�ዿ��Ͽb/>��:>R�>��R�-z2��Z�8b���Z��S#?8�:�y~ʾ�΂>0O�=�Hݾ�Vƾ�KA=��8>�|i=W����[�_��=[bw�08=	�d=T��>)F>FY�=����Gh�=��H=���=i�R>H�!�,���+�\�4=�A�=U�b>^�+>P��>T�?K0?YXd?�>�>�n�_�ξ;���/�>��=�(�>�=V�B>>��7?�D?��K?k��>V��=:�>{��>͘,���m��_徺ħ�s	�<ܓ�?�Ɔ?D�>�+U<�\A����yc>��0Ž�l?M1?lt?3��>r����ƿv#E�B��Ό��i̽��=|���+$@���뽆�V=^��l��>�?���>z�:�N>�Պ>q��>w�>��=�>+7�=.Y�����=&[��@�<U�;>��>�M=^˽��=�_�=�&�{��Ո�=1�>h��=���>�?>2��>�=I���D/>9����L�Hȿ=%H���+B��3d��H~��/��U6���B>�5X>�{���3��`�?��Y>p?>g��?q@u?��>� �R�վ�Q��Je�WS�Fĸ=q�>��<�ty;�AZ`�B�M�F~Ҿ�=�>Ȯ>-�>��n>YSG���R�G1d�=���=�>��?�D��q
	���w�Nj|�P���'����i�?ὰz/?��{�䞁=�t?��L? �?4��>�|><���5̴<����ſ뽥�:���¾��#>V�?/�?��?9G�C�S��魾�_4�(0�>�C�fU�*#���.���
�ھ�V�>�
���@޾�T8�C愿r���X?B�{{�4��>,<.?>{�?�D����iRZ�E��%�l9�>_]m?���> `�>��?򄡼W6��Ό�}�>u�z?(A�?���?`Է=���=���Ց�>`?D��?Æ?%d�?v�!����>þ�=��=x㗽���=YZ{>�,�=� �>��?��>0��>\1a�{�������{o��lv��.�
=���>��>ϐ>�ߤ=x\9��=���=Ƴ?>3[�>< �=��>�ƞ> /վD!�{�"?��$>6>%�F?}�=>a�&>�&=x��<�֮=�����>��Ⱦ�=���ܗJ�"�w��_O=@�^=�?^���A!�?��k>����??���=P=p$4>J~>q���1��>�
�=��}>D�@>�%�>�Р��y�==�O=�,Ӿ�>��Sm!��4C�̄R��Ѿ�5z>j���
�%���w���V�I�����w�0j�6��C=�S�<�C�?5����k�v�)�T��đ?x,�>T6?)���.���d�>���>[��>�H��A���\ƍ��TᾸ�?���?��c>
��>�OW?��?�0�43���Y��u�iA�[�d�(�`�䍿f���Ga
��g��v�_?��x?�A?���<�^z>҃�?I�%��X���Պ>X /���:��9=���>�f���)a��uҾ�þ�J��G>w�o?[�?R�?�~V�
W��.%>��<?�7?F�z?��:?z=?J�3�0"?,�>j:�>�?!U+?�,?W=?ª@>;> ���<����Ɯ�.��ф���ռɝ=��=�4����_<dn=�5=��D�f����=gZ�oi���5=W�s=Ai�=0Ϩ>�f^?Zx�>�>�`7?���#4�-���l0?�Mw=�5h�i}�+���ٻ�t|	>�	j?,�?}�V?�ay>�J���K�خ/>GC�>^�*>�wV>��>HK����>����=h>E	>sX�=�Ȁ������9��Ꮎ�}<?�>��>�1|>�����'>_w��E,z�{�d>k�Q�ZȺ���S���G���1�|�v�sY�>��K?��?1��=C[����Gf��.)?q]<?�MM?H�?��=��۾��9���J�S8��>+9�<���󿢿�"����:����:w�s>|.��������b>O}�}�ݾ��n�CJ���oBN=���`�T=�7��־�^~��b�=L�	>�J���� ��!��7��J?L�j=�,����T�PW���>��>��>��?���w�%@��:���D�= @�>�;>(כ��~��gG�iM��W�>ĆO?[?��?r���:��@���ľ+&�@���{�>8
>t�
?*O�=n��=c���lW���H���?��E��>��>����C�$"�S������<i�>���>@�D>W�-?qD|?޵�>Pq?|SC?��#?�>
�;k����V0?�V�?p8�=���`ؾIVX��!<���?���>��&�#�>�&?�G?H3�>hGQ?&?�J�>T}޾	V��{�>ü�>��t�����?M>p�/?](�>��H?�
�?7�*>e��Hz�m[���$>i\�>�
�?�7?�o?/?D��>�YѾ�ݾ���>(�z?m.*?�hu?Ee� XX>�5+>�A�>��h=�p�;���>�M?�=8?·[?L`?�j�>�~<٪ټ[+�����αt�nܽ!�-�a#,=��/�;8������;�=p�'>�L3��i�z��=�<�4�=�=�S�>C�s>A����0>��ľ4G����@>/u���M��+Њ�#o:�OǷ=Ą�>��?㩕>�L#�ʒ=���>�@�>����0(?V�?�?_�*;�b���ھC�K��#�>FB?���=A�l�联�1�u��+h=��m?g�^?�W�%��$�b?��^?���7p>�a�Ǿ��e�w��P~N?��?7�>����>���?[�q?Z��>��q�16n��圿}b��xc�G��=��>����_�D��>�4?�q�>^�d>Z��=�oݾ�2x�z��b�?>4�?[o�?���?/;>�o�Y࿢���ά���Nt?���>yό�Gx,?��K�d+g����E&��u����J��ⲙ�����?f/�P卾��
���=��?e(t?dw?<Y?; �?�i���b�|҃�G	P�a�������2�=H@�PT���f������d���� 4�£����P�n8�?.C?`O���
?l��-�Q���ž4F6=�r�����\Z�=
���W��(��<3�x�� W��w����*?���>� �>�K0?-8Z���K�f�:��4A�����
�=�G�>k%�>�5�>>^3�AC�(��7���y����K�+��>�l?�:?�P?�hǾ5�R�걎����}/#�K�j�j�|�5�^����>�-�nŞ�pJ�c�,�lu��5XM�R�������>c�^?hZ>f�;���?�N�>�b��[��0l���t��te���>l�~?5�>y�l>��C��Se�Z��>;�|?$�>+/g=�rܾyI��Ԏ�2ؽ%��>�G�>��>���>3_��v�e���h��4N��J�;��k?7�s�mŅ��ti>r�k?�Z�;9_��ܽ>� 1=�|�0��*����<8>B#?�b�=���>�x�b�8�'���(�վ0�(?`?A�����!�<-�>G� ?���>Az�>T��?��>$���G�p;���>�Y?�J?zB?�~�>-/�<,����ӽ5�I�<���>�}>��=���=��3�rV�~���<=Q0�=V�L��؊�Y˨���'�_�<R=��%>Ooۿ#HK�_�پ%
���M>
�6ވ�V���qo��I������T!��qx��Y�4�&��;V�O`c����l���?/6�?�U��Q��p���8���s���'��>�q���������;��r������!_!��O��i�*�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >`C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾s1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@�yA?��(�G��u+V=���>%�	?��?>�V1��H�`���[V�>�9�?���?�M=ɿW�Aw	��e?��<��F�|=޻	�=�f�=Ma=O��2|J>JC�>q|�v0A��Wܽs�4>.�>L1"�3��C�^�wԾ<�]>`�սP6�� Մ?{\�jf��/��T���V>��T?�)�>m:�=��,?�6H�\}ϿC�\�+a?�0�?��?>�(?fۿ�Nؚ>��ܾ1�M?D6?���>�d&���t����=�1�(������'V�b��=���>3�>F�,�Ћ�j�O��E�����=!��=���d�"�)X.��*��(���Q�<D2#;�R�;"��r> ���~��΄>�>�<0>���;wE��k��>�ؿ>�1K?^pe?V�?!��>�3>�.'�;�ľ�����F�/�?Gv����B[��tݾ&�����Y
����~�_=��=�(R������ �6�b��RF��.?�#>�O˾J�M��f:<��ɾ^��('��5�1̾�61���m�k��?Q�A?�Ӆ�s�V�>��=��}���
�W?"����۬��/�=V��g)=��>�f�=��⾊3�!US�Q�:?ͷ4?�����v��=Pv"��Ɏ=>�?�?��>�M�>XJ7?ޯ��+d���i�=��>��>�]�>�Q>1��K[���H'?��V?Vn!=1Y!�>J�>S@ƾ�	�Q`�>�A�><[��v��]�>��g�ؾiƁ���u�|x"�:BW?�>**�����ܐ�{K*��l:=Гx?��?�@�>�[j?�C?�8�<p�����R�����=�}W?��h?q\>Љ���ξ���*�5?A�e?D�P>jCj�J���.�y���?��n?r�?s6Ѽ��}������/�me6?��v?s^�ws������V�V=�> \�>���>��9��k�>�>?�#��G������mY4�Þ?��@���?��;< �[��=�;?j\�>�O��>ƾ{������_�q=�"�>���mev����3R,�\�8?ݠ�?���>������N>�=�G��3>�?C�|?�P����=?� ��~J�/k����m}<F.�;��G3��;��ݾ>���K��=�<��>m/@�p3�U��>S}���>�p�п=o��3���}+��"?�n�>���jþ¤i�O|���[��YE�9g���U�>�>'|��4摾��{��x;��蟼��>U��5�>�S�j��ي��]84<��>��>忆>��������?*N��;ο�������ĽX?c�?dm�?S~?��:<��v�45{�ݰ��+G?��s?d,Z?+�$�'�\��6�$�j?__��hU`��4�HE��U>�"3?�B�>A�-���|=�>���>"g>�#/�~�Ŀ�ٶ�b���L��?��?�o����>h��?s+?�i�8���[����*�ԍ+��<A?�2>݌��)�!�00=�!Ғ�Ǽ
?o~0?p{�n.���_?��a���p�I�-� �ƽ,ߡ>;�0��m\��5�����iVe�����Gy����?�]�?�?¯�� #�4%?�>M���29Ǿr��<�|�>�%�>�)N>g+_�\�u>���:�Nn	>T��?d}�?�g?��������[>��}?�$�>��?]o�=Za�>�a�=I񰾧-�lk#>�%�=�>�'�?��M?L�>=U�=�8�0/��ZF��GR�)$�1�C�G�>`�a?D�L?�Kb>2���2�~!��uͽ�b1��R�Z@��,�m�߽�*5>��=>�>��D��Ӿ��?Np�8�ؿ j��$p'��54?0��>�?����t�r���;_?Sz�>�6��+���%���B�`��?�G�?=�?��׾�R̼�>>�>�I�>>�Խ����[�����7>0�B?[��D��v�o�y�>���?	�@�ծ?ii��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*��ֿQ���Czɾ�=��ٽ�=��=��0>�s���Y�=��< �M��~<���=;i�>]�V>Rj`>�GJ>)v>vz�>����2"��W�������O�Jd�G��eQm�������7����L�ľ]��RZ��Rr��x۽���G\���»�1�=��U?�Q?7p?�� ?��u�& >U����=�i"�q�=(�>��1?�L?��*?`�=������d�nO���>��Fᇾ|8�>��I>	��>hf�>
�>յ���|I>�>>fY�>`� >.U'=�����=��N>`k�>���>S9�>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��w�T�4:>9����j�5`>�+ �~l���)��%Q>wl?��f>�u>�3��d8�8�P�'}���h|>�36?붾�E9��u�W�H��aݾFM>2ľ>�3D�l�q���<��ti��{=�x:?4�?+2��MⰾJ�u��B��	OR>�:\>�]=�i�=�UM>�Uc���ƽ�H�m.=u��=�^>�?*\:>B�=f�>)�`�E�����>r��=e�>E)Z?��E?zv8��m����7���D��Q�>1�>� >Ro>7_f�K��<���>Qt>���=�=��{�0\>j(ȼw��c,����ƽ�b��p>��r=w���eO�ͫ�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�g�>�x�xZ�������u���#=<��>�8H?�V����O��>�w
?�?�^�֩����ȿ2|v����>O�?���?I�m�A���@�{��>5��?�gY?�oi>�g۾Y`Z����>Ȼ@?�R?��>�9�I�'�}�?�޶?˯�?�^�>*�?,�a?J7=��}���%��ﳿ�N���q�=ͨR>u��>���=����.�j��F��P䎿J"���k�\��>`�=e1�>3�I���Ⱦ���<wD>=!՞��N=.z�>	N�>z\>.�>8C�>^��>f�>�����f���k��T���K?���?-���2n��N�<?��=#�^��&?�I4?�j[�w�Ͼ�ը>�\?h?�[?d�>4��L>��B迿7~��۩�<��K>+4�>�H�>�$���FK>��Ծ�4D�fp�>�ϗ>�����?ھ�,��SU��;B�>�e!?���>�Ү=+�?<2?�Ē>˜>��S������^�"Hm>/]�>\�?U(x?��?B੾B�F�KE��s����[�>J�y?�U?���>_���F���X��c%�<Z���h`?�:X?xG�=�%?f�l?O�E?�~ ?�?�=�k񽞩¾À�;�8�>[`?���T5��5���ٽ��?�e?@��>��v�ỹ�=[�����F�?N�_?i_%?�/��jc��j����<<���(��Xƅ<č0=۞4>��>_�Ͻn̲=��>辵=#
w���=����<A��=f�>���="+��j��@=,?4�G��ۃ�>�=l�r�?xD�P�>aJL>x��h�^?�l=���{�x���x���U��?���?@k�?H���h��$=?�?H	?�"�>9J��X}޾d��APw��}x�fw���>���>��l�O�G��������F����Ž�^����>���>sO?� ?�Q>⋲>m��T�&�����O���^������7��..��E�K�����#�������/J|�7J�>�쉽z��>��
?6�g>|z>A��>y�ӻ��>��P>�5~>4Y�>j�W>�55>=>�<��ҽ�KR?����'�'�z�辬���a3B?�qd?E1�>�i�6��������?���?Qs�?$=v>h��,+��n?�>�>G��Rq
?�T:=9�;�<V�����3����'��>E׽� :��M�jnf�rj
?�/?�����̾�;׽ƽW��+�=0�?��?Ǎ6�(�U�`��+aG��4�I�"�r����}�6��S�;���_��&�f8�CV���%?> �?A�A�0{��"������6H�]K���?�T?\?ayK>lo �����͂�4���/վ���>���?���>�B?ZO1?�L?�X@?�9�>��>cy��/<?�=���>е�>%�?wX)?&'+?��?*&?9H&>���� �&x߾�?�?}�?+F?\�?�:��q���*��<�U=�����g�u7�=l>U	˽v@Խ+OF���5>�?
4��9�I���Um>��6?�9�>���>����;��#�<XQ�>�=
?D��>������q�c����><Q�?�����=+>�Y�=I;��m���:v�=$k��+�= ���s_>�$�></6�=���=0H��Y�H:x�+;�%�;PR�<u�>8�?���>�C�>�@��0� �a��f�=�Y>:S>x>�Eپ�}���$��r�g��]y>�w�?�z�?�f=��=ؖ�=�|���U�����>���H��<�?=J#?(XT?_��?y�=?^j#?׵>+�jM���^�������?R!,?S��>_����ʾ���3�\�?6[?>a���<)�c�¾�Խ��>�[/�T0~�p��2D��-��V��%~�����?���?A���6��u�����^��0�C?�#�>�Y�>��>�)���g�1%��3;>u��>�
R?�%�>`�O?�5{?O�[?�kT>J�8��)��sҙ��2��">� @?���?��?y?�|�>��>S�)��"�N[�����"�傾7W=�&Z>���>B'�>)۩>���=NȽ�R��Z�>�b�=d�b>K��>+��>�>w�w>�<��L?M�?�t׾~� ��y��hg���D���px?ɸ�?l�?�ө<s��v-�pr�<��>��?a��?"�/?P�8�nm�=����Ⱦގ����>$��>:�>�(/<u��=�?>�S�>���>fO��#f�%�G��:&��F?u+)?�
:>6�ɿ�
s�@t��9�¾/J��}��6�;��yս���O%	��sپ*Q�������������!笾�tľ��6����-�>��=��">9��<%N�;$�o=�$�=�!>hϴ<��⼳���ӕ�=Ͻo=!�<���.	=��j=���<�껙E˾�s}?%$I?��+?r�C?�>z>8�>pk5���>���f{?��U>�cW�;D��+�:��d��^"����ؾ�A׾��c�<Ο���>q�H��W>�l3>>�==҃<�=��r=�ˎ=�Hf���=E�= ��=,��=�4�=SS>��>v6w?���ò���3Q��V�۶:?p9�>�v�=��ƾ�@?��>>�2��͗���a��-?@��?�T�?��?�ti��c�>����㎽�s�=����'?2>u��=�2�袹>��J>f���J��D���f4�?��@{�??�ዿ��Ͽ\`/>��7>%K>yS��	1��hY�(�b�oW��!?�;��$˾�d�>��=�z޾�wž)2=^T6>�Im=�����[�b;�=�z�asC=x�l=�̉>&�A>�=���.��=�YE=_�=�rQ>?�亓]J���0��x8=s��=_�c>s%>a��>��?�Q0?$[d?h2�>��m���ξ�A���F�>r�=�Y�>�ۅ=�B>ҙ�>��7?�D?��K?�[�>.0�=���>F��>�,���m�e�񼧾uì<���?^̆?�¸>,}P<�DA�ʓ��\>���Ľm?=C1?�{?��>Mw��Vؿ�k+��\=��4�����(x=3�i��`�
*�|���a����E>�e�>e��>�9>���=/�>Zɡ>���>��>:1c=�����P���%�<�p=/t >1��Y����߽�m�<bh>�&�<�q�������#�=M�<@J<���=���>�;>]��>���=��`/>�Ɩ�׷L��-�=5���*B�s<d��9~��.�I:6���B>X>X���1����?�Y>�?>L��?gBu?! >�=�¾վGL��+1e��gS� I�=�>��<��o;��Q`�=�M��yҾ���>�6�>��>��k>.,�$$?��r=���;5�b9�>�U�����zc�{Sq��F��"퟿�	i� ��D?W8�����=5~?��I?я?�(�>kĘ�9Kؾ� 0>Y���{*=��Jp��>���4?�'?1�>Dh�f�D��E̾���,�>rHI���O�}���0�0�xʷ�+��>������оn#3��g������d�B�
Xr�n�>P�O?��?P0b�X���VO����K��6r?�zg?��>M?�A?-��v�s��jh�=��n?i��?=�?

>�w>Ģ���G>	ZJ?�u�?��?�2�?���a�>�KE>���>2�����ɾ��>gt�>O�>?�x>�M>�� ��f�-E���C�������z���=�C�>�UA>92���a��]�=_��>��>J�=�$�=6�S>=�>'�i>�t�����N?��D>2��>�?\?m~>;��>^8^�q�1���J���3������=<�$��
�������d4z��h?,��[Ң?	�=Ɩ�f�(?��4��p�>�y|>�0>�.�=���>����y�=A�T=ě >u�>>*I�=�K>r#Ӿg�>ۮ��v!��7C�m�R�@�Ѿfz>�t��w�%�G�������;I�q������Sj��;���1=��g�< ;�?�B����k�H*�d%��-�?{q�>��5?���OV��qW>`��>��>�E��O�������k�c�?���?�;c>��>C�W? �?��1�3��uZ�.�u�k(A�'e�N�`��፿�����
�V��-�_?�x?/yA?�R�<&:z>N��?��%�Tӏ��)�>�/�$';��?<=k+�>)*��9�`���Ӿ��þ�7��HF>��o?<%�?tY?CTV�eKk���%>D�9?:�1?�Et?�2?$�;?�]��$?4A3>z?�K?hj4?��.? �
?hS1>7��=ʘ���",=�'������o�ӽpν�K�hR/=v+z=Mo�:W@�;�=f��<�����ۼ0��9nɣ��f�<��6=�
�=�%�=��>�c`?�U�>,k>.O0?�/'��J3��ݢ���0?�9=���4�v��Ś��쾚W>�ro?�ʫ?�4V?�*k>ʲD�ѓO���%>�/�>Se<>��s>�W�>�	��Z=���=��>��>�W�=:����$C��:�����;0%>	��> 0|>+���'>�v��3$z��d>��Q��ź�L�S��G�j�1���v�([�>��K?��?F��=�_�0���Gf��,)?2[<?�MM?��?��=x�۾9�9���J�\B�2�>�<�<������"��G�:��g�:οs>�1���x��~"a>����޾�n�L�I�>m�K�I=	���W=Z����վ�P~��Q�= k
>`���,� �����"����J?��j=�d��f�T��G��>�>g��>�@�>mT9���t�Gk@�[����&�=�K�>y�:>=��Q��L�G�-��"�>+�X?��U?�w?2m�낿�xK����Ο��6>��?�u�>B��>��s>
&��ھd���sb�x�O���>�` ?׿(��CL��e���̾%��c��=�m�>����o�G?��t?�y�>F;?ӄ?��?���>yJS=g��O)?�Q�?5��=>�����o7��m@��@�>��%?�&�f��>V
?�?P�?K�M?��?9>|���5����>h�>�uU�P���'>�hD?%ã>��c?��?]�N>y?%�8������P<4>	>�*A?��2?�"?���>���>	{U��<�'�>���?/lo?׎�?�q�>��a?�	u�2B�<���_ؽUh�>��?��2?���?�`?a�!?W�<w�D�c��m	���2
�=Q��=�>��Z<H��k��� ��*�n���y�<\ >�:=��Ƚ��`�>�s>��� �0>��ľBH��?�@>����yF���؊���:�:�=��>D�?ܪ�>s\#��Ғ=^��>BT�>����0(?��?�?_�";:�b���ھӪK�(�>JB?���=��l�9���u���g=X�m?W�^?�W�a)��k�b?��]?�f�|=���þ��b�����O?�
?��G���>��~?��q?���>�f��8n����lDb�]�j�XѶ=Zq�>FX�7�d�>�>՛7??N�>��b>9*�=u۾��w�r���?��?0�?���? .*>��n�{3��\�޺��ғO?���>|�����2?c�#��[��gt��Vݾ���/�о�΀��l|���ݐ�W ��N�Q�*=�$?�S?2��?x?���cr�Z�~��N��w+�'{1��h�",�qL(��YL��j�5�⾽v���	���<6�K�orM�'[�?��E?-j����E?د�D{��6ڕ�R�ľ��龢���d>X�D�c��쀽����!�����83?�H�>�1?��?��}�C���H�s�*����"�(>��(>(��>���>~��F�2H�kl`�z2�����>s�m?��:?/�l?���K�T�te�����~��|ܜ�=��h�@? ?½Ƚۜ�I5>��.��bi��(��g��C��� �>�&?|3�>k��>sH�?�?I|�y[%�Vվ"UE���
�=��>�+�?,E�=��+>a��=��߾��>��l?���>��>ޕ��nZ!�p�{�m�ʽ&�>��>}��>��o>+�,�#\��j��T���D9�Hv�=��h?7���,�`���>]R?]��:��G<B}�>ݧv���!�����'�[�>�{?���=��;>n�ž�$�p�{�y7��#U(?��?����z*�)��>]"?�l�>HV�>���?���>|ž��3�|�?��]?�J?=qA?9��>�A=y�������{ �g�$=`�>��]>�|i=��=S-�a;J������"=h4�=�)ҼC@�k�;Z:��O<-7�<(!>+fۿJK�щپ������%
�+܈��Ѳ�`��L���`���%��%x�d�p�&�
oV�6fc�h����l��~�?8)�?�"��'䉾ө��~������{��>3[q�D΀��������������Ӭ��V!���O�.<i�K�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >[C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾q1�<��?7�-?��>Ŏr�1�ɿc���v¤<���?0�@}A?u�(�\�쾤V=*��>��	?��?>`U1�oI������S�>�;�?���?_vM=t�W���	�x~e?k�<��F�D�ݻ�=�;�=�E=6��ȔJ>�U�>x���LA�Cܽ��4>�م>�|"�e���~^�5��<_�]>�ս2��/Մ?&{\��f���/��T��?U>��T?(+�>�;�=��,?Z7H�U}Ͽ�\��*a?�0�?��?1�(?ۿ��ؚ>u�ܾ��M?TD6?���>�d&��t����=�4�}��@���&V����=Q��>��>�,�����O��I�����=��������u!�1c�K�=���<�̞�E� ���߽����C ��pc��������=��	>_��='NE>��W>L(>+�N?�P?֌�>N�~>-ʧ���)�%�Ѿ��U�G�`���x��� .:�4��n�IY������h��e���"=�,��=h7R�b����� ���b�f�F�l�.?�o$>��ʾ-�M���-<slʾպ��G���8襽U+̾J�1�� n��̟?��A?R�����V�G��JX�	|���W?|L���� ꬾ���=!���M�='$�>���=p��/"3�*}S�_3?�P*?����+��I�>c;�=5<c>\d?��>Z��=���>b 5?Ǿ�ؾ�y�>#�I=k��>�'!?Au?��ľN-m�ǟ/?f)�?�D�:^Ն�o��>I��������g�=��Ӕ�]��=�(�>+���뭘����=�Á=Dȶ=��_?-��>��(��]F���o�ר;�:�=��?���>�h�>��[?F�@?���Ֆ;�����MѾYC>�]c?|g?�.�=a�!���B h�e�o?��j?�	x>��ƾ݀�D�����D�A?غJ?�?���=zmy�����m
�T�=?��v?s^�ws�����F�V�g=�>�[�>���>��9��k�>�>?�#��G�� ���xY4�$Þ?��@���?	�;< �L��=�;?o\�>��O��>ƾ�z������U�q=�"�>���~ev�����Q,�d�8?ܠ�?���>������z}>>l�g�a��?,��?��	��e�=���`�4.���ٽ�������=}����a	�Q�E����T�(��߄F��ę>��@I����>�@��V���2���$\i���9�>�?�S>���w�]䇿�{5�ds>���Z���K��T�>�>�������{�Iq;��^����>����>�S�� �������y5<8�>���>췆>c���⽾�?�Y���<οo���٢��X?yd�?�o�?s?�9<�v�;�{�c��G?,�s? Z?��$�.]���6� �j?y_��kU`��4�[HE��U>�"3?�B�>J�-��|=�>���>�f>�#/�l�Ŀ�ٶ����\��?��?�o����>q��?�s+?�i�8���[����*��D+��<A?�2>"���4�!�(0=�rҒ���
?Z~0?{�m.�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�$�>��?ro�=�a�>He�=P�_�,�:k#>�!�=��>���??�M?�K�>�V�=��8��/�[F�]GR�$��C���>V�a?��L?�Jb>����2��!��tͽ�d1��M�9V@�?�,���߽�(5>��=>c>�D�FӾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?LQo���i�B>��?"������L��f?�
@u@a�^?*wS˿)���Pr澶�뾵';<C���|�<ό���H�;ğ�=Q�6>�>�l>πm>d:0>ӫ%>׬�>X�`>�Rg=^`��T�"�e�������c�A�-�Z31��k;�k:�B�A���׾L���\��׌��(�������x� �L�l�\��~�=mV?�vQ?�?p?��>V瓽�>1���_��<Տ���h=��>�3?�@L?@})?��R=K
����c��w���P���I��Y��>��>>���>���>)�>�n)���D>�4>�σ>�a>Ma�<�G��"L=}Q>5P�>�>a�>�C<>��>Fϴ��1��j�h��
w�l̽0�?����R�J��1���9��Ҧ���h�=Hb.?|>���?пf����2H?%���y)��+���>}�0?�cW?�>!��s�T�2:><����j�5`>�+ �}l���)��%Q>wl?ֺf>u>ޛ3�&e8���P�|���j|>�26?�鶾�A9�8�u�H�H��aݾOLM>�ž>��C��k� ���R�\ti�?�{=7x:?��?J1���ా�u��B��QR>�8\>�J=d�=�UM>�fc��ƽ�H��V.=���=�^>�I?�,>y͏=x�>����*N�(ƪ>�B>\P.>�t??�T$?_������� -�:-u>-�>��>|>n�J��\�=���>�e>�y���3���$��>�"_>��~��m`�Ձ�ԣ�=&������=�ӑ=Z���e�<��=�~?���(䈿��e���lD?S+?^ �="�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>׫>�ξ�L��?��Ž6Ǣ�ɔ	�-)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?��r>�c�?.�k?�m�>藄��w>��k��Y㌿�����2=v�>^�F>����9����lk��XTh�0U!��6>`�]=�Ļ>^5-�g�����=�i��3�����F��>dFP>�5`>NȢ>K?bO�>�/�>K�:=};��xV��t��"�K?���? ���#n�&f�<�O�= �^��"?�B4?7�X�f�Ͼ޾�>��\?���?��Z?b@�>���;���濿�z����<��K>^�>k<�>��ZoK>��Ծ�7D�s^�>�ٗ>~@���Pھ�&��i��\D�>e`!?���>��=�� ?a�#?W�j>�,�>�]E�<���E�ϟ�>|z�>tL?��~?��?�ܹ��P3����I᡿}�[�o�M>��x?�T?ݕ>X���<����C���I�)D��Y��?�hg?�P�U?&3�?��??a�A?�e>u�1�׾�g���ހ>߄!?0s�L�B��r&��g��?�?��>�fm�IQٽ�j�����j����?�[?Q�&?x��
_�l���	��<�����U�p�<�I��)>X�>��ᗾ=��>��=��j�S�5��s;���=E��>���=&8���\=,?�G��ۃ���=Q�r��wD���>NL>d��s�^?�k=���{�����x��U�� �?Ԡ�?gk�?	���h�X$=?��?		?!$�>�I��x|޾ޔ��Qw��x�Cw�h�>���>?�l���>�������\F����Ž�<�T�>F��>6? � ?S�O>�Ҳ>��1�&�i�5����^��S�XS8�1~.�����Q� �����6¾#|�R��>�F���5�>k@
?!zg>gt{>ۮ�>õһl��>2/P>0�>#�>��V>YV4>W(>�m<��ҽ��Q?]a��	(�!��%���]�A?u�d?g�>k�R�-+��*Z�.�?�6�?L��?x>W�g���*���?^4�>�-�B�	?O0=LhN�y��<8r���f��=��b��G��>:�ѽ�9�̣L��>d�Ѓ
?I�?ﰄ���;;Rܽ=�w�(^�=[��?�-?��/�E9T�`Et�>zO�%5\� �<�������1�-�Uaa�����s�z�����O�=�� �0R'?ő?IT�C���`�GC����G��SK>'�>'c�>O?�RN>������$z����s��G��>�c?m$�>��H?�2;?'�P?B_M?�`�>I��>u���3K�>
��;���>U��>?�7?��+?�/?�O?i�+?b�l>��ܽ���ҋؾ�?��?K<?�8 ?�=?�0���7�����'(��<
����l�캓=[�<��ؽ�,f��P=8�K>�?���:�7��,���p>�*7?���>�6�>�Ċ��n��qq�<ѯ�>OZ
?�*�>S��eYr�U7��c�>7Â?��C�<Mm(>�b�=0No�����v�=s;Ƽz�=�Ē�5t;�E<$�=�ə=0V��8;���:�� ;��<�t�>�?���>KE�>�;��x� �U���f�=Y>�S>�>Eپ~}��2$����g�^Zy>�w�?�z�?��f=��=4��=:y���N�����O�����<t�?UN#?vVT?۔�?��=?�j#?h�>m+��L��>]������?w!,?��>�����ʾ��։3�ם?h[?�<a�	���;)���¾��Խб>�[/�i/~����<D�9���[��4��?쿝?5A�T�6��x�ٿ���[��z�C?�!�>Y�>��>Q�)�w�g�t%��1;>���>kR?�$�>�z]?1_h?��Q?��+>-N�D���������D6O>��M?S�?�.�?~_?m+>�\>J�T����U}��_�� �/φ�ep=��'>m��>��>l��>�U>��ӽ�2���v�&�>3�I>�??�%�>���>ր�>[��;ؓR?c1? p����-�.ᾏ��Hw��;�?L�?b�;?	u�="-��*U�Xo��x�>���?�w�?uS7?��m�:7�=��=��׾������>�W�>��>'��>� ����=S�>���>Q�彚K?�" �,�ͽ��>�
X?a1>;�ɿ��x�����?�þ�VO��^��'4o���c�U������=lN���?;Ŗ���<E��H~�C(��ä���?��_���,�>������
>��=�fͻ�=7�&>���=��)�u~s<�&���:�`�˻� �=�9�d�i���Ｆ����X=7}˾��}?�8I? �+?e�C?��y>W>Jt3�b��>�����5?��U>2P�v~���{;�۸������ؾ<X׾|�c��ȟ��H>"!I�f�>�:3>�B�=�B�<�#�=~�r=ۤ�=noT�s2=XJ�=�^�=�x�={��=>�>�;>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�g5>g	>4�R���1���\�'�b�rSY�.!?�>;�J�˾�>�Ż=_޾�Hžڣ2=��8>c=�|��<\��4�=$�x�o?>=�k=��>1)D>b�=����9��=�J=���=(PN>[b���{7���(�ڳ3=�=S�b>:&>�?(@#?�$?3�C?�L>vA��T�ƾ����E�>{��=��>�>�i>�Z�>n�1?��5?�>?��>ø�=���>u�>s�+�El������ԁ�������?�Ώ?rm�>x�=��y��-<�"8\������-=?
�[?V�!?T�?&�A����U�� 8�t����;�M>g���*ɏ�Q6>_�}>eUj=��>�w7?Bs�>߯
?؛v>�]��>���4�>�+>�X�=�[>��=ώ�=<L@��>�=t���א��g��;��<�6p=E:V����<=-;���������k��=���>
<>���>ɒ�=����F/>U�����L����=�G���+B�{4d��I~�r/��U6�-�B>�?X>�r���3����?�Y>�o?>���?h@u?��>��
�վiQ��DDe��US��ϸ=A�>:�<��z;��Y`���M��|Ҿ��>��>�>��l>,�@$?� �w=��a5�x�>�~��D�����6q�.?��:����i�L6Ժ}�D?�E��+��=!~?+�I?��?��>���ԃؾ�C0>ME����=���.q��Y���?'?%��>�쾃�D�|E̾�	��߷>BAI���O�f�^�0����˷�]��>+���F�о�$3�Eg��������B�dKr��>u�O?$�?�5b��W��mVO�����,��tp?�}g?��>�K?QA?�/���z�du��Bm�=W�n?��?c=�?>]�
>Ŧ�����>�?g��?�p�?h�~?�xϽ[+?�����>=�2S����<
2>'C>���=k�?�M%?��#?Mf����	�W$��xھЩ>�^>=�9�=?�|>僉>��0>^Ǥ=%�=Md�=���>�֐>w&�>9e2>��>B>̑���0��n&?Id�=+ƍ>�2?2��>b�U=恪���<�MQ��`B���(�."����߽X�<��
�YbM=g�ּ}J�>*�ƿ�ۗ?��Z>w{��?q����@)�m�T>wL>���;��>۰E>\�w>%��>�J�>v=>֢�>�C&>�FӾ�~>����d!��,C�F�R�}�ѾD}z>�����	&�ޟ��w��1BI�`n��cg��j�J.��B<=�Nʽ<%H�?������k���)�����X�?�[�>�6?ڌ�6��ѯ>���>�Ǎ>�J��e���_ȍ�hᾗ�?2��?�;c>��>*�W?)�?��1��3��uZ��u�(A��e�<�`�l፿�����
�N����_?�x?VyA?=^�<�9z>(��?��%��ҏ��)�>�/�';��@<=�,�>�)��]�`��Ӿ�þ�6��GF>K�o?2%�?QY?�TV�J�^�)>�:?B�2?�u?g1?� <?EC���'?K�->��?-�?#w4?�-.?*
?��'>1��=]��;m�V=o����䊾�fν-�½��ʼz�;=�`}=�B�D�;^`
=��<Vg�� Zټa�;EΉ��#�<�I7=Lם=���=��>��[?���>]Ë>�A:?-��Cr0�L���u�1?��+=�������Z�����ޟ>��d?/"�?3�\?q}>X�B���F�#�#>�w�>!�->�Q>+R�>��L����y=iU>�>V��=x�ృ����`��8��<o>��>�/|>!����'>�{��0z�f�d>��Q��˺���S���G���1���v��Y�>.�K?��?p��=�^龐+��KIf�0)?�]<?�NM?��?m�=U�۾d�9�p�J�>�b�>-U�<��������#����:��`�:Y�s>_2�����fc>���ij޾�n���I���羮�L=��zT=��q־��~�'�=�w
>u����� ����̪�`�I?asi=l���vU��蹾V�>�ۘ>H®>�(9���t�vg@�$T��䵗=H��>�;>����(��M/G�j�.Ԉ>N%F?Ɉ]?�'�?�h_q��bB�X����S��
�ټ�A?�t�>l[?C>�
�=<׹�#��S^d�� G��T�>[��>�Z���E��(��I��}#$��a�>�O?��(>\X?NyL?U�?m�`?�*?,�?i�>�Π�)���'?ar�?h[�<eE���jl,��G��4?�.?���.�>�m>h=	?o�'?�W_?���>dM>����Q�դ�>LȆ>�Q��3����>'�&?#�|>r~f?���?���>�n���ξ�'X�+>�.�>�}w?�R?]o:?��>ъ�>��Ѿ�[ʽ�5�>��n?�@}?�j?��2>�m�>,u�=0��>�U�=��>(�?�[�>~�B?��U?�)?2'�>�4���ƽ	|	��Ž��l=�z���e����=��-=�}����7>`+�;�W�I%��ͽ��.=�Zݽ��你��<2��>^Xm>u_���*.>�b��B,���B>��h�����̺����6�Ӱ=@��>� ?j�>���̕=˺>"��>���'?�?+?�%<�b���޾qlI�I�>�KB?�d�=@�k�rߔ��4v��^=��l?��[?�Z�������b?�^?S�c�<���þ=�c���龁�O?�
?3�F���>��~?��q?���>Ff�[+n�%��O1b�
�j����=ja�>�S���d����>3�7?�<�>�c>���=��۾��w��Ǡ��@?���?\�?�ˊ?�L+>Z�n�'����j꒿�m^?F<�>�ߦ��%%?^�S����\����[����ݾQ ��� ��H���f��9{&�R<���ٽ�ռ=Q�?�q?
v?�F`?�< �}a�_��I}�~�S�>��.��1�B��mA��l@���o�ȷ�rI��윾�a	=bЛ���_�t��?�NR?8�-��#?�Ǿ�wl�V���v(�l�x��S���o�Z>���L(=�H|1�Q���ٴ�*?��?3�$?iz/?�yJ��G���1� �Y�������=g�=!��>	?����a�uj�{þE��ݾ;��>�?z?my6?gP1?�a��3�?��耿1���0��X��>W��=�[>'XU����zk���.��l�}�-��P��ʧ���Da���?��I>@,�>�U�?���>8s$�@�о���ij�i�#>>�2m?��3>T�m>��X����4��>˩x?:�>]֒>x"���=��އ�����g?&��>%p?�զ>tH�ƛA��q���]���@=���=T"Q?�ц��4K���\>�SJ?Ӣ���[�=]�>^�b�\\�֘�XE����[<rv?f��=\f^>v�Q#���r������(?�t?ۯ���w(�{�~>m�?Ž�>8��>�?���>��ľ�G���\?��Y?�I?k&@?m
�>ޗ[=�����Rʽh�+��08=y�>��_>��S=���=A�"���P������P=�=��̼�ӽR:�e�<��;���<T�1>Umۿ�CK���پ��U�S>
�8刾X����e������Z��c���ax����PA'�[V�\<c�磌���l�'��?�:�?|u���'��{���c���$���g��>��q�͈������/��x�ྻ���xc!�_�O��$i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�4?��'�����&?E:
?�W<>��;�Q���a��B�?�"�?Dcv?l�Ͻ�8�<��=RUK?b�G�c��I�|<�>��*����\�ǽ;�R>��>��U���v���E�co>�>�½��H��> ����=��J>'�)��Yh<�҄?�#\�(�e�.�/��E����>��T?�r�>@I�=��,?4:H��mϿ�x\��a?h/�?���?�)?~S��lۚ>E�ܾ�:M??6?dR�>eD&�j�t�8��=�p»�㾊SV�8��=��>k�>�-����j�O����T��=������4]<��6��͉<�]c��Y�:)�f��S��)�oLo�|K���-�����'���]>΄R>f�+>�w>ڥR?ϰT?S'�>k]>id6�/�<�X¾[tK���5.���3%�����T�b ��E�����Z ���	��V��(#=���=�7R�'����� ��b���F���.?�x$>b�ʾϾM��`.<�wʾϪ��䄼7ӥ�03̾��1��n��˟?��A?���y�V�����������W?:J�d��u嬾O��=!'����=�4�>|��=u��3�5xS��^8?��?a���s+}�h��=���F>h)?2_	?�G>iހ<�~?���=���M><�=��>�9#?^zC>����I�Qx?xa?��8�0c���>T�̾��}��|��x�C<+綽�>��V>:1���Ǿ�cֽ7p�=}��=�V?���>��*�_�W���TG��b@=r�v?�F?N`�>rzm?��C?e��<����|�Q����=�n=��U?a�i?�c	>0-v��GҾ�,���b5?��d?�+N>'�k��꾗�/�j� �n=?5%l?��?LVa�kz��P���a��7?��v?s^�xs�����M�V�e=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�%Þ?��@���?w�;<��S��=�;?l\�>��O��>ƾ�z������8�q=�"�>���~ev����R,�e�8?ݠ�?���>������o��=+���޲?�ʋ?�q��d�=�.���h�@�@_���C8=2R&�I�L��Ӿ:8�����Z1���־C�Oߖ>�X@����>�����8�¿#����־�U��T�>o��>�T���۾�i�y!a��:I�=L�^���vU�>��>t���b�����{�ma;��f����>��c��>�iS�^A������5<��>m��>霆>�i���彾&��?�A���7ο����Ǒ���X?XU�?Wi�?f�?_<<n�v���{�����G?��s?�8Z?Q�#� �\��7��j?_��-U`���4�MHE�kU>#3?sB�>ѓ-���|=>֊�>�h>i#/�X�Ŀ�ٶ�r���k��?���?�o꾇��>]��?�s+?�i��7���[����*��,��<A?b2>v�����!��/=��ђ���
?�}0?�y��-�d�_?W�a��p���-��ƽۡ>	�0��c\��I�����zXe���0@y�m��?P^�?W�?��, #�-6%?��>螕�8Ǿ��<���>|(�>�-N>AM_�ίu>d�p�:�6k	>���?*~�?�i?��������rW>D�}?�(�>�?p�=^a�>�D�=6𰾄,��V#>F�=V�>�G�?��M?X�>:c�=�9�G#/�|QF��6R���G�C��
�>P�a?�L?�>b>����W<2��!�+�ͽ�f1����'w@�w,��߽�25>��=>>��D���Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��W�s����>�B�?�{�?��>!�l?��o�P�B�h�1=8M�>͜k?�s?'Ro���d�B>��? ������L��f?�
@u@_�^?)iο5;��-򵾪���gH=4�=�PY>:}���<����@������z>�	�>-l>�c>6�k>�`:>gR>�S��ƾ$�P������&�j����;��v�����l#��[�)�oٿ�Z���5Ӽ���i���^�~���VJ\�P'�=�U?M�Q?�no?Z��>g	z��>�/��Ş�<P$�8��=>��>U2?BL?ø*?���=_A���d�IS��{�Ğ����>oII>���>U��>A��><Ϥ:q�L>{1A>`�>Ca�=��%=�y":K=�Q>O��>7��>��>�C<>ё>?ϴ��1��h�h��
w��̽*�?����Q�J��1���9��Ʀ���h�=Gb.?�{>���?пd����2H?%���|)��+���>�0?�cW?�>���T�-:>u����j�M`>�+ �ml���)��%Q>tl?[�f>�Qu>;�3��]8�s�P��z��>|>�&6?���_9��u�f�H��Bݾ8M> ̾>�SM��m�����!��qi�hM{=�]:?�~?5���λ��y�u��3���zR>�a\>�c=�[�=�RM>�~b�29ƽ��G�AZ.=e�=$�^>��?�.>#v�=q̥>�t���(J��Ű>�*>>>E>?��?=����ڼ��~��0�kb]>��>ߴ�>�>C�T�짏=)��>"Q>L���n�[����X���Q>6����K��Y����S=e���K��=��~=����1�T�U=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?��>���?p_q?m�>�׽��H��������)��=�k>��>Y,{>0�Ae6�.3��D�z� ���8�͈z>Ɓ=���>�O$�4-����=������8�E����>��A>F�>>Y��>Pp?��>1[�>���l�e=�Q�
�����K?Ƴ�?`���n��x�<iI�=m�^�m?��3?�`�=�Ͼ7�>��\?���?�[?T�>����0���տ��[��5�<��J>��>td�>:S����J>׉Ծ��B��Ɋ>/˗>iL���3ھШ����8��>pm!?���>���=F�$?��4?ˋ�>@�|>)7M�p����_�m�>���>>9?�>y?|0?e����&����9#���Z�����=k
m??F?��>^������
�=&�� ��Mi?0�t?��o��?��?�i??G?���>X�1��¢��ڀ=6̓>	�?�'�:�R��;��Y(=?� ?#�>���m�"�7|/>"�����`��>)�\?�C?����]a�����6=�>�<������^\"���!>{�>��ӽ�#\=W��=z��=�=G�HB�=�900�=���>���=�P�b�@��=,?��G�ۃ���=��r��wD�K�>%IL>�����^?Jq=���{�r��fx��!U�� �?��?�k�?	��a�h�=#=?��?!	?*"�>*J���z޾��ྕLw�Ux�yw�W�>���>j�l�'���� ����E����Ž������>F�>��?�>5�N>5�>�D����'��(�_��^�|���B7�a-��h��y����#�P�o���! |��Җ>�ϊ����>�?�i>,[}>2L�>zEe��Ћ>f;H>��}>;�>f[>��7>�>�[><��Ͻ.R?3����'�Ή�Q��*0B?�nd?=+�>�i��{��m���X?d��?6i�?�v>.ah�K+�hg?�0�>T#��~L
?�':=`q���<:����pF�����㴎>��ս":��M�K~f�%G
?�$?*���̾��׽t$Q���>>ǒ?O�8?
E��<^���z�y^���W���k��c����<���<� v�
k���Q��Q��&�[�b�53?��?P��m�%���߾�.��QD���z>�z�>�?��>a��>��2�V-�W�^��+��f����?�|�?c��>8�/?`$?�j?�6?
��>� �>��a�>U�=��=�|�>>lL?�!?w{?l�>�s?�"�>���=H ���޾��>7??�<?"=?�?b�!����Pݽ��;�gľB���5�&>�>2ٶ�����8X9>Y�?3N�E�8�f���(�m>327?��>���>�厾s#���u�<���>��?�>7c��g�p���
�Ce�>�&�?�z�p* =�Q)>/�=C�l�L���
�=Oz��C��=@Qp��d&��j <��=��=����b��3�i�X��:>��<cx�>��?5��>�?�>�>���� �q���I�=�Y>�"S>��>�<پ4z���#����g�QYy>,x�?�z�?D�f=r�=C��=&|���R����������(�<��?�K#?TT?��?��=?j#?@�>e.�N���]��0��S�?x!,?��>�����ʾ��Ӊ3�ڝ?g[?�<a�����;)�ِ¾��Խб>�[/�g/~����0D��셻���s��1��?�?YA�P�6��x�ٿ���[��u�C?�!�>Y�>��>P�)�y�g�q%��1;>���>jR?W��>�5Q?Q2z?�PY?��N>��:��z��&��%���`->$�@?Á?��?�w?��> �>@�3��ྔ����C�}����j=K�V>P`�>S��>��>"�=�ؽ�m���2G���="Ad>A��>
��>$&�>�	u>�N<t�L?j�?L^þ�}'�V���(�����J\�?{��?�(C? 6 =v�D��
/�<9����%?���?tg�?��0?5��Y�=:���L���?��o�>�Е>%~�>*N�<�ʽ���I>��=6W?N�S<������:˼M?�\?�6�>�ɿ�Wr�����^ֱ�o�P<�a���IB�B��5i��-:=5D_�i�۽�Ⱦ�ٵ�����}��r�˾�$�����;?�"=0�S>~�/>��9���6=�/;5׈=O�=��<�@��<!#�'&y���=�"l�ÊT���6=�T=�˾}?�;I?�+?��C?��y>�;>��3�U��>7����@?V>@�P�����2�;����c ����ؾ�w׾-�c�Kʟ�BH>Y`I�'�>�83>�F�=�I�<��=Os=7Î=R��=�#�=�O�=�g�=���=T�>�T>�6w?W�������4Q�6Z罥�:?�8�>J{�=��ƾi@?��>>�2�������b��-?���?�T�?7�?!ti��d�>E���㎽vq�=D����=2>r��=��2�J��>��J>���K��Q����4�?��@��??�ዿ΢Ͽ>a/>�
6>���=�U�Z�2�c{$�(DN� �O�ۻ?��5�2�˾�3�>�W�=�ܾ��ѾXP=��V>ԍI=C�#��4R�iƜ=�P��X�<nE�<"�>A><�=�1ͽ_�=[�=��>�7^>t�мB����Ҽ�x=pM�=�K>kR1>|��>p8?��/?��c?.��>n�XmϾx���q�>%��= �>�m{=ɀB>yǸ>�8?��C?�hK?�>7v�=��>���>_�,�A�m��]�n����e�<枈?��?)��>H i<��C������=�G"��Ȓ?R�1?�?�
�>�n�P,ٿ��E���V�=.�ڹ�w39>(��z'���w3��p�d�A�f��=/	�>���>�$�>~��>�e�>��`>ͅ�>l>#>�����A=�UA>Ho'��i��Ge=2Sr��Y&>q)>�t�=`����1�9���V�=��=~�<^�޽{��=���>=?>z��>���=�����U/>TȖ���L��Ͽ=]N���'B�'d��>~���.�\o6�w�B>�XX>>��]2����?��Y>*h?>���?SDu?? >-���վ�O���:e�8kS�=��=��>�<��v;��W`�A�M��xҾ*��>��>��>w�l>@,�4 ?���w=��!a5�b�>E�������64q�*<��9����i��6Ϻy�D?�D�����=~?�I?w�?���>-����ؾ_C0>;B����=��e)q��I��R ?�'?5��>��ξD�|U̾_6���ҷ>�JI���O�X��� �0�P��Vȷ��>�몾��о)3��j��b�����B�Eer�8�>*�O?��?y?b��Q��,KO����p����l?�}g?� �>aF?=?~0���~�xe���ܸ=<�n?q��?�9�?>���=�{�@��>?�{�?�ސ?��y?sw�����>���f@>:P��fse>�B>%W�=8�=�=�>F�?��?H�潁������W��.T�d	�=#	�=)[�>�pU>.�%>>�W>K��=�r=��=?l�>���>�* >V�='I>�����9��o�>~)�=iW6>L1?��B>�5<>Az���{:�>�=�.l�5�۾���K#=$��=����f���':>�6?�S���?���>R���NA?���N�>�f*>���=�^5���=u^f>�?��>�to>.��>@R�>�KC;�FӾ%>����d!��,C�u�R�ɾѾ^{z>����&�l��xt���DI��o��h�j�v.��c<=�ѽ<H�?Ը����k���)�`���
�?�Z�>�6?_ٌ�z��t�>��>Jƍ><J������ȍ��hᾖ�?&��?�<c>��>��W?՚?I�1�A3��uZ���u�(A��e���`��፿����s�
�����_?t�x?�xA?
E�<:z>#��?�%��ӏ�C)�>�/�+';�sH<=f-�>�(��p�`���Ӿ3�þ�6�1JF>c�o?q%�?�Y?UV�:I;����=Vo?t78?.>�?dN?U�U? ��p�?+�i>i'�>���>b�M?�1+?��?��=�x>�� <��<�~ƽ�9��>�S��R����j���3J� `\�O�}�-g=_j�=��U= $�=��<"�!�eQ�=�	q=��<�j=���>�T?���>?R>-�?�zD����h���`�)?�>�Aɾk�:�19� ��06>��Q?��?��p?DV>M�L�dn��)
>��>NEU>��W>��>-ZO����ᚗ�6��=iS�>>�>N���ھ	c ��@��l�=d�=Y��>	�{>ݎ��C'>v��+�y�-�d>M�P�񚺾sS�?�G�w�1��u��5�>��K?��?X'�=���X`��rf���(?4@<?	ZM?Z�?��=�۾�9�p�J�C��g!�>iu�<����������v�:�TK/:ˆs>� ��x�V2W>�		��*ݾ:�l���H����@O=A�=*c=Z��!׾K-��)��=pm
>�ľ�#�؏�������lK?@i=(#���rZ�Tθ���>�
�>3��>n�m�:Q���@�"��s�=n��>�/5>ݓ�Z��b�H�	��5E�>�<?	hX?M�?�����X^���D�-ӾM>Ⱦ�9�mb?�(>O�#?u�g>W�b<���� �\ms�>_H��U�>B��>u���\��g��ܒܾB�뾏�q>�?u6v>X�?&EO?8
�>4|a?/:!?z?u��>�<&����(?�σ?&�*=Ei��tq���<�dy<��5 ?��#?����x�>��?9(?p>)?�M?�;?��(>��񾽳>���>#��>�\�	���HAg>�G7?څ�>��c?��?Un5>@|!����6�����=��n>�=?~h(?�#?�7�>E��>L���"	�gj�>L�?]m�?U|?Bf<3�?��z��q�>������=<�?s?8�_?�lY?OB?�� ?�A<�Y� ����04<������Y�Y����dG��3��r���$��Wr�R�/�	�W���<�1_=�.����=	>�b�>��s>|����0>��ľ�S����@>Ӣ�eH���Ҋ�Ew:���=|�>D ?ĭ�>�F#��ؒ=_��>�E�>9���2(?��?W?S�';��b���ھp�K�W�>*B?���=��l����u��ah=%�m?A�^?^�W�i��f�b?��]?4f��	=��þ�
c�;��D�O?_�
?BG��ҳ>T?]�q?�Y�>�Tf��%n����r<b�0�j�Hf�=ap�>�E���d��D�>ǟ7?�B�>��b>l�=Ev۾�w��8��� ?X�? ��?��?�v*>��n�a(�]���s��7`?l��>�Ʀ���$?pSZ�n�ξ<n������]��l&���������2����'��v����ڽ4{�=!�?�|s?E~m?��_?�.�}�c��0]�[�����U��x�<�BD��B���G�W�n���@��7⛾H�8=�d��p	T�f�?��?F� �$?����mӾ���fh6>���gx���">�[�WW[=���;K���[A/��}ھ�h3?��>�>��B?uTz��<4���%���O��uؾ>eY>�p
>�q>���>o��&%f��N�gM���`��E�ԽR�{>��[?#�B?�u?�r�}�+�p.���������Ǟ���>�gY=J�>�Mj��E��$,�� <���}�|�����]�
��B�=�a,?B�>�>���?�!?1��।��vx��j3���j=�]�>�#d?	�>��>a���a!����>stk?u��>�z�>�|��Nb#��ց��!����>�u�>�S�>���>�;���
e�>���K燿�E���=��V?��^�B�>ПK?�c����=�ͮ>"����M�x��>��p��=�} ?���=ç<>��ξ�׾X�b��ę�i>)?�)?�'���*�,>�<"?ػ�>E�>[,�?���>� þ�S���?+�^?�CJ?�VA?�C�>�I=���FȽ��&��*,=���>��Z>7�l=*7�=X	���\�g���.D=^R�=ַռ�S��/<d����L<#��<[4>�Aڿ U�����OX �B�ܾ�8��=��IX��14������_�޾N��@���󛿽�6�������9�����$�����?��?<4�﷚�~T��WW�11���>%������=��۾�`����+w���\R'��+]�t��~�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<	-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@1�A?P�(�n��t�U=���>�l	?�4?>m�1��B������1�>�M�?��?�K=��W���	��Be?n�<��F��5�w�=�l�=�v=M����J>�_�>�U��@A���ܽ��4>$م>�"��z�\T^�:��<�^>��Խ�ӕ�cԄ?�n\�bf��/��P���?>{�T?k4�>�]�=�,?*H��zϿJ�\��"a?�1�?��?��(?Jſ��ݚ>�ܾ��M?�>6?���>*d&�ƴt�j��=k��v���/��t"V�p�=ƫ�>��>�,������O��	��h(�=�a�e�ÿg�u ���=M�ש
� @g��j��`E�pȾ1��N�T�'�>� >�8>qײ>N��>�K>�L^?%�C?�Z�>�x>�20��q����-=Iʾ�`>(֠�������d��~���ӵ�l�+�Ӏ����/��7��=�|�=�'R������� ���b��F���.?|O$>F�ʾ��M�+-<�yʾW���0x��n	��,̾�1�!n�N̟?��A?Q�W����T�}����W?zV�K���׬�^��=KN��u-=�6�>7 �=c���3�H{S�w�/?��.?V��|�þ�M>�]��u>��'?��?����?��>B��f����>��+>���>á?��>��=��)=?̕j?�ھ����"	�>�	
�v77��n�=5�<&���ԉ>jt�>��o�R���T�(����BW>��V?��>�.�z3!��ۋ�� 5��~=�_y?�F?�S�>�m?�=?h��/F�4��.d�=�[?�h?۠�=�����ɾ���-/?N�h?�Ns>6�q�4g�s�.�g ��S?�3l?7�?«2�\Ɂ��L��`�x�7?��v?s^�xs�����L�V�d=�>�[�>���>��9��k�>�>?�#��G�� ���xY4�%Þ?��@���?x�;< �R��=�;?l\�>��O��>ƾ�z������6�q=�"�>���ev����R,�f�8?ݠ�?���>�������y�=Tﱾ��?S��?��(�=,i���p��� �-�k=|O���=�̃=�L�7w3�\پ!��������}�>�5@���"��>Ej྄2�#�ÿ�u���Y��5�|�?u0f>1y/��� ��}�[)v���Z��KP��d��NM�>ЏT>.���c墾Jy�E�7���J�>Yy9�Do�>|<6��r���쌾���=��>y&�>���>��߽�s̾"�?oo����̿:���9]�5�&?ա?��?]Y0?�y�=�1���a���X���;?k`�?�t?�e�=S�E�i׼'�j?t_��qU`��4�oHE��U>�"3?�B�>O�-��|=�>Ǌ�>^g>�#/�w�Ŀ�ٶ�`���P��?؉�?�o���>l��?ms+?�i�8���[����*�)�+��<A?�2>����<�!�40=�EҒ���
?a~0?�z�j.�J�_?�a���p�>�-���ƽ�ڡ>R�0��b\��;��l��"We���� Dy�(��?Z^�?U�?�����"��6%?��>枕�%8Ǿ��<j�>v*�>!/N>5O_��u>��e�:�;j	>1��?h~�?(i?Z��������U>�}?�b�>��?��=uG�>��=4ﰾ;>�+~">D�=U�9�4\?��M?���>$.�=T�9���.�WF��R����n�C����>J�a?ShL?��b>�D����1��� �|^ͽ2�/�sf@�h'��Uܽ;*5>��<>{>rD�Q Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ya~����7�k��=��7?�0�0�z>���>��=�nv�ٻ��R�s����>�B�?�{�?��> �l?��o�R�B���1=:M�>Ĝk?�s?:Ho���c�B>��?������L��f?�
@~u@e�^?'�hֿ����[N��C���J��=��=�2>.�ٽw_�=��7=6�8��=�����=w�>��d><q>F(O>}a;>�)>���P�!�	r��Z���O�C�������Z�B��Xv�Xz��3�������?���3ý�x���Q�2&�0?`�Z��=�SR? �P?�t?�F�>����� >-o�è�\>"�WwK=��[>B�:?oKI?U"?�=*֝���j�w����������έ�>�5>WN�> ��>��>�;���pY>L>3W�>k��=ե=H=?� =PbA>w��>���>	�>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?g�f>L u>A�3� T8�~�P��}��G|>p36?�����C9���u���H��AݾA2M>���>�F��k��������i��C{=x:?p�?����sⰾ�u��6���DR>7\>9 =�2�=HkM>��b��ƽ�H�m�.=��=͐^>�l?	1>�W�=���>>����K�8ȫ>d�?>��0>$#??2�%?��1���Cn��
j)���u>9�>�C�>Wa>�TR��L�=>+�>��h>�޼մ}�0Z��I��cV>(}�P�g�8Iq����=G�F�=���=%�v�=�J�/=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾUh�>mx��Z�������u�/�#=C��>�8H?�V��;�O�g>� w
?�?�^�੤���ȿ8|v����>T�?���?c�m��A���@����>:��?�gY?toi>�g۾@`Z����>һ@?�R?�>�9�~�'���?�޶?ӯ�?�|�>#ʋ?^@N?���>W� ���>�����°��E���A>:�s>c��>wm��S�\�����bx����y#���S>���<+��>����Ež�YH>���j�-�r��>�p>u_>���>he?���>�r�>���=L�\��W��������K?���?'���2n��M�<~��=��^��&?pI4?�`[�u�Ͼ֨>�\?N?�[?�c�>S��C>��8迿L~��e��<��K>4�>�H�> $���FK>��Ծ�4D�+p�>�ϗ>�����?ھ�,���M��"B�>�e!?ϓ�>�Ѯ=�
&?0�"?E;>P��>P�L������Q���>�ة>>�$?-�p?�?䮭�S�A��@���/��̺l�8��=�g?��?�4�>��aЙ��|�=&�ߏս-�{?��k?c�3�P�?�?�eG?6?��p>z.^���ξ.��W�>��!?7 �$�A��I&�P���?�S?���>�"���(ֽ��ռ`��P���� ?�(\?�B&?����%a���¾�F�<+�"�[�V���;�:D��>\x>杈��n�=b�>ǰ=R]m��_6�K�f<�w�=W��>��=�7�kV��F,?+�(�h�����=�Mr�1KD��t�>��M>9�	,^?��:��{�����A��Q�	��?Ո�?e~�?�ϱ�Ȇh�f�<?�?�6?�)�>*����Gܾ8���Sv�B<y�90�V�>���>��O���oŤ�����)	�������W��S�>�R�>� ?X��>&X;>���>先��N.�}��$0��c����>4�J.�����a��m�X�'^�:�;-
��jO�>|�~����>wG?�[R>��|>���>\&5;5?�>C8>��>���>��e>w�>�[>`�\;�����IR?3���C�'����ע���5B?_sd?�-�>7�h��������~?���?�r�?oEv>jyh��)+��n?C�>���o
?.A:=���Ud�<BU����,G��I�⣎>J׽�":�M��mf�Gk
?�/?m���P�̾�׽��(�g�w=�c?�*$?��g��j��y���p��]i�d�=�y��%���b�̉��9�������䒿 E�~Qy9?�L�?�/�����b��z�A�K��8>�>�>�6?=�%>�3�����W����wo��Rڥ>��z?�D�>=WM?�o ?ȹQ?6M?Ѿ�>�	?����?I$ý2��>f��>g�"?�FF?�?_0?Oe?���>%R>�^�����?L�"?9�?no�>~�>4/��c;3��5��K�n��i
�Fe����<�5���Ｙ�Y�(!=�H�=:Z?��W�8�����c�j>X{7?t�>��>���"�����<��>�
?�:�>� �ryr��f�kO�>%��?E���=�)>���=�=��κ$O�=������=�`��Ғ;�QP <T��=���=5�r�uts���:�h�;�B�<u�>7�?���>�C�>�@��.� �_��f�=�Y>7S>�>�Eپ�}���$��n�g��]y>�w�?�z�?��f=��=ۖ�=}���U�����=������<�?>J#?%XT?_��?{�=?^j#?۵>+�lM���^�������?�!,?���>���a�ʾ�𨿾�3���?\Y?<a�î��:)���¾��Խ@�>O\/��-~�z���D��2�����1�����?龝?�	A�v�6��v�����Z��Y�C?��>�V�>�>��)�c�g�\%��8;>k��>�R?�c�>��O?Զy?��Z?HPQ>��8�n:���k���j��(>�>?��?�5�?�<v?Bi�>�>R0����b����s*��2�����O=�\Y>�>P��>�T�>�k�=+MʽR���p�:��ا=�d>:�>^�>>��>�|>���<{N?��#?^��>e�^l`�˴���;�N�?/�?:�?�}�>����|�jw�� �@?�e�?ү?NF?��4��̌�>.��p@�Bi�[��>���>=��>F�����:>Ĝ�<��>�J/>S�:�iL�q��i�<���>a�=?��>��$�����=|9�����=�ȵ��`��r�=�@��a�=�@㾛�2��	��o��U]������=�������^վ>?����k|>C3/=f��<~�>1^���z?=!k>48Z��
0����=i@�=I�=83;�*e=��Mv�=�Z��d�˾H�}?98I?՜+?��C?��y>~e>��3�ϯ�>o���hC?V>�P�9�����;��������ؾ�d׾d�����7>��I���>4E3>�"�=���<�:�=S�s=���=��\�
=��=BV�=�s�=���=��>�@>�6w?ؚ�����?5Q��X罷�:?�8�>
��=��ƾ;@?��>>�2��ʗ��Rb��.?���?�T�?��?�si��c�>d���厽Vq�=`���'?2>���=�2�[��>�J>g���J�������3�?|�@?�??�ዿX�Ͽ�c/>#�8>��>>�R�n1�*�\��c���[�]-!?�5;�1˾��>&)�=�[޾=Ǿ:)=We6>&�Z=���e\�xݘ=WNy�t�<=�jj=H�>>�D>7H�=n����=Z?H=���=��P>eTn�T�6�Y*���3=Y��=f�c>�N%>��>�?	*?{�Z?��>�p��cʾɭ��{>�
>�~�>R�!=o�W>���>,�*?b�5?�J?ZF�>�=;:�>�>��4�WG��/��x����X�=yه?��?��>�:G=�����/��e2��D���?vR9?�?�Ҝ>�h�0�޿���(u2�jq��~^<Ƚ�=�����=�3L��x+��FI�Q��=fe�>0��>��Y>��3>��k>B{�>���> �#>��Z=xw�=KoG=��P������W=�R�wx��!N�����t.�����o��X�d<"��u��<@�=+�=)�>{9>d��>&��=���)>���2�M����=����z�B��``�e~���/�5�:�(�=>�1K>}0��&��� ?�X]>s�E>v��?��q?��>�8 �Z�׾Z읿��h�a��a�=�u>b�4�|�:�m^��O���Ҿ���>��>��m>�g�>�6�*r�G��/ܾp7?�͕�>�3~����=�Ӹ=ԁ~�ǡ�@,����b�k���?8
��f�����a?�U?�a?�U�>���=����O@��#��=�y���W��u$�z��=y�?���>��?��/3�)]˾�滽���>D^H���O�X����z0����鷾�Ա>ۇ��$Ѿ(S2���؏�
�B��}p�C��>��N?��?{�^�Ss���nP���J����Q? gg?x��>ν?�_?F����<����5�=�Xo?���?X�?�H>Qe�=Tˈ���>$�?�:�?��?])�?{�|�C?)03�^�>����'�=;�?>�{�<��]>�L?p�?1�?����/0�)d�
���J4�0�=f�?=@�>6e�>9:e>&A�=���<���=�"><[�>>z�@>n�S>��A>��¾b@���@?�$c=H=�>M�5?�A;>
��=S17���2=s����Y�Gf���ӽC_Ҽn�������^�.��>�����%�?��!>��z�?�5��	�i�i8�>��> �ļ_z�>ia>���>�0�>�U�>q�=�> �>IBӾ��>���c!�#.C���R�$�Ѿ?rz>柜�2�%�ʞ��t���BI��r��,i��j�/��u==�2��<�G�?������k�g�)�5�����?�W�>46?�֌�����5�>���>pɍ>7H��@���^ƍ�dg���?���?�;c>��>@�W?�?1�#3��uZ�&�u�i(A�0e�P�`��፿����
�q��.�_?�x?1yA?XS�<.:z>Q��?��%�`ӏ��)�>�/�"';�#@<=r+�>"*��+�`�~�Ӿ��þ�7��HF>��o?;%�?zY?2TV��)s�x��=[�+?CC6?�z?�=?z�H?T��6?���=t�?(?�,5?F�0?m�?��r>b0>����o��=�n��f"��������X�yU`=�a�=�&t=�Z*������ؼ^/="��<M��;E�A��u���C�<Be=��=��>F�]?M?�>|�>�^7?%���6��%���[/?��4=��홋��򤾱��{
>�Gk?��?��Z?��f>W�C��
E��>G|�>�z#>��`>�մ>���sC��9�=�>[�>��=�@�ϐ��KF��!��[��<��">m��>»|>D���vw'>kD���y��{e>>�Q��C����S�'�G�K�1���v�P��>.�K?��?`�=���垓�Gef���(?��<?cmM?��?x2�=a�۾�):���J�"'�gM�>��<|��Ґ��x����:�B3:Us>�㞾�T��Ӱc>�l�>
޾��n�@K�8��I(N=H���J=#�
�Ҿ�G�bI�=�Y>~��U�!��A������\pI?�o}=V�����\�Fa��b><(�>)B�>��(��+��]5@��|�����=�}�>q�@>x��0�G��U��0�>y6?�J?��}?:z���ˀ���T�t6Ǿ������q?�F�>���>ښ�=r���۾�y�Rv�|gP�KY�>��?�[%���a�q{��5h��\�>)�?�*Y=��?�S^?ӝ�>ʖF??F�"?�@�>3(n��t���q5?;�~?��
���v��ા�eT�%?���?9?�<"�_H�>Ͼ?y�?�L�>��@?��?h�r=����4H����>}��>��W��Q��vT�>��E?q�>�fY?xe�?`q>D�'��|���fD�����>e7?�#?��?Q��>{�>ږ������-��>z?o�m?L�n?�yd�-?�p�=W�>%�S�6�=%x?<�>4N)?�`?�'Q?�!?�`;jö�l>���������b��g�l��`�saB��8=�9B�u?,<:�������5co���=����f�<�*z�ws�>Dt>�7��-�0>��ľD���A>6衼/��.���z=:��-�=���>�?J��>��"����=,˼>>b�>I��k"(?�?�%?�N&; �b���ھI@L�1�>��A?��=�l��w��4�u�V�f=�m?q^?��W�=
����b?��]?*]�{�<�fBľ:d�q�龤�O?�s
?�G�I#�>�?�q?�9�>�g��n�^��WVb�/ l�B=�=%�>�c�43e�ˇ�>Ut7?�]�>l�c>9p�=z�۾�w������?٢�?c	�?���?��)>�n��߿}k��7Œ��_?yi�>w����"?+��o;����K���� �g�����������ਾ�8%�1Ȅ��(ѽ�E�="�?�q?n1s?�l^?=E���b��^���}���U�i@������B��C��UA�V�k��-�_������=�社��g��ؾ?0�	??A�1��>\J����hƾI&�>|!�P�%=Ȇ<:���nD�>���}0��	!�N'��R	B?��>jnR>`^?����9�m&O��V����}��>D��>n[�=:��>�-�m������Ѥ����db�>��^?a�0?\�U?��*�dp>��^���)��F�_���E>��I>�+�>ҿ������9�4mT�W�f��!������2�=I�>?��9>iS�>-A�?�� ?c,�9���3Ն�@b[�L�;��H�>�O?�:O>�p�>�N=��*����>[�l?���>z�>ѝ���f!��{��ʽJ�>��>���>�Cp>�J,�4:\��X�����;09��*�=��h?s����a�T�>R?X{:	tI<J|�>��u���!�e���'��Y>_?�
�=O�;>��ž����{��M���/?��?���@}7�}�S>Y�?U��>0��>�Q�?z\�>�i�����?A�Y?�TT?@&H?̄�>���=����3�R�-��'�<�܄>Bq>j��=��=_�3��Nb�f�&�zc=��=⥫�aȽ�%4�U��<��Q=��=�l>vۿ}�K�G�׾������ù	�ߌ��@X��^����������q���y��&��3/��$V���c�����l�v�?���?����ʉ�%Z���e��8��ʿ�>�dr��	�������
���H�߾Ư���� �3P���h��Df�P�'?�����ǿ򰡿�:ܾ3! ?�A ?7�y?��7�"���8�� >mC�<A-����뾬����οC�����^?���>��/��p��>ߥ�>�X>�Hq>����螾�1�<��?6�-?��>Ŏr�0�ɿc���m¤<���?0�@W�A?�(����E�T=:�>�	? �>>�K1��f���$s�>�F�?��?MbJ=7�W��-	�#e?�;�G�PWٻ'��=�L�=��=���j�J>�V�>Q��jl@�2�ݽ�=4>���>	�#��1�I.]�;�<�	]>=�ֽ&���hԄ?��[��If���/�bJ��w�>T�T?���>��=��,?�G�YϿ�\�va?v	�?ƴ�?=K)?׿��x�>�{ݾ�$M?Z6?�>[K&��t����=����v��p}㾑�U�ۓ�=3R�>,�>�.��.�?MO��������=����ʿyM�˰ �~@�=��=I�.<��Ž���m���f��ܙ��:�	%<����*�=�-P>�B�>��U>��q?BH?�f'?I%>f�c<��B��� ��Y�=J���Y��.���������^���k���徙F.��W�u��|�,�_�=�N�����R(��]p���L��K&?���=�;�k=���=�¾ǵ��P��k�����۾�)8��6w�t�?	hH?�j��+�d�GJ���,漡�����]?
������N����>�sN�Ȫt��U�>���=�bᾇ'6��t@�xM??�_*?s*��=��	<q1���<�*?+]�>���=x0�>^^�>^�<<�r�Q�>Oo�>Zl�>C��>�P[>���X�p{?7i?�r��A����>{��poS��ϻ=��=̎��m��=ן>�
�em�Ҽῴ��=^=�)W?{��>_�)���e����t�<=t�x?Ȍ?'�>�xk?*�B?�F�<�v��M�S���U�v=�W?� i?��>�{��Iо���"�5?
�e?K�N>�fh�7����.�U�?|�n?�R?ٜ��q}��������q6?��v?�r^�ys�����]�V�[=�>�[�>���>��9��k�>�>?�#��G������hY4�'Þ?��@���?S�;<� �A��=�;?s\�>�O��>ƾ�z������ �q=�"�>����}ev�����Q,�X�8?ܠ�?���>��������=nɰ�>p�?}��?'�ܾsм�./��dw����Tr>��X��~�<��Z=����&�be꾲##�I���r��r	�>��@�薾���>lF���n��̿�_z���
�:Ӈ��T?���>t��<�����=T�g�C��
@�����4�>�G>v!ս�>��X�}���I�&�]��	?©�3f�>V[,�X����w�/E�<ms>9��>!��>1�����K��?����ҿ����T"�$_;?�_�?��t??tI?L_�=��S�p���!b�=%�Q?���?�u?���=�:�=�nϽ%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�d�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�M�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>kH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?�q�>��?8}�=8��>�h�=hX���;G��#>��=�<��?{�M?Y��>1��=)8�p/��F��3R�o;���C����>o�a?��L?vb>d�����2�v� ��uν4=0���tWA���,�9B޽F5>��;>�>Q�C�$FӾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?hQo���i�B>��?"������L��f?�
@u@a�^?*�fֿ��5M��ޓ��D�=�=w�2>ڽao�=ѫ7=iA8��\�����=Y�>��d>q>d.O>]_;>m�)>��� �!�\q��y�����C������X�Z�e��4[v��x��3�������(���5ý����gQ��4&��M`����=g�U?�R?�p?�� ?)�x���>Ԩ���@=�#� ф=f.�>�i2?r�L?ɢ*?�ړ=����W�d��_���B��kȇ�#��>�rI>L��>�J�>�$�>{�Q9g�I>�,?>�~�>�>e'=�"溶e=��N>"M�>���>h|�>>�<>�
>_����*����h�e x���ͽ��?�����J�f
���y��Rw��ǻ�=�>.?�>���l=пB�H?x�����4f,���>�0?�-W?ϴ>�f���PT�\�>��� j���=���2Ql�=�)��Q>F�?Yi>�Ew>�Y/�Y�4�P��4��<�k>��9?�c���xI�g�s�2�I��q澻�2>p:�>�
�A!��l����|�ԣm�E�o=��:?�`?�@��燰�M�k������T>��X>�x=*B�=�P>Fn��J޽��8��A�=�[�=awo>f ?�H>�B=B�>Ԅ��&�C����>2�>�2L>S�@?'+?vܽL�$�
�D��&D�z��>F��>֏�>�>D��le�=�U?�>��
=�%��`�̽��]��H>;u���*D�b-���=�oc�Jj�=�|<9y7��P��s=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�u�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?roi>�g۾;`Z����>һ@?�R?�>�9�~�'���?�޶?֯�?_I>
��?2|s?�6�>��y�ZY/��/���b��rY{=0�5;sM�>kU>0���1�F�ܿ���_����j�v�Ua>_4$=��>��㽚7��~��="����%��q�e��޷>�Sq>��I>9`�>�� ?/k�>�|�>=n[��ɦ���?��w�K?��?����3n���<�t�=B�^��#?�E4?��Z���Ͼ�ߨ>�\?»�?)[?�`�>5���<���濿�����c�<��K>�8�>hE�>|���>K>z�Ծ<:D�[v�>W˗>���E<ھ�&�������.�>Tc!?���>��=�g ?�#?�7m>Բ>4GE����>,F�U��>���>v�?�k|?��?�P��@�2�I8���I����Y�b(8>du?X??L�>󧏿Gj��@c���慽��a�۪�?��h?�3ͽ��?,��?8�@?^LC?h�c>lq����ξ�z��q�z>��!?�	�c�A��J&���y?�J?���>+W����ս�Nּ	��,�����?�$\?�7&?\��I-a�@�¾��<K�"��|T��P�;e}D�C�>:�>�{�����=�>�߰=�=m��.6���h<H�="��>>C�=l7�;��G,?3|��jۇ�6�=�r�7�A�Uy�>�5E>9���/]^?�92�h7}�
ɪ�赙�ÜV�Կ�?�S�?��?�����j��j:?\��?��?>��>��ٸ־	�澡Yq�A�u�%�����=���>bR�Rx�I8������첃��IԽ��ֽ/��>Q�>�$?�E�>X>�p>�j���hD�#��$����f��6��TH�����54��ܲ���̾�ソ�þ*�l��7�>�*��6g�>���>n~>�v�>Kr�>���O��>��F>�>���>��=�Ճ>3�>��e�=�KR?����$�'���辽���b3B?�qd?Q1�>Bi�:��������?���?Rs�?#=v>h��,+��n?�>�>K��Tq
?vT:=9�`;�<V��w��$3����*��>E׽� :��M�Mnf�tj
?�/?�����̾�;׽�j��ǚ8=�]~?(�:?i7�i�\�/�}��Q^�q�]����=� 7��3v�Ӫ��?i�����d΁��!��u�'�~�^���3?N`�?����~��ĳ�<�����3��Б>=a�>c�)>���>l%�>�J�T�+���i�����z_���>`�U?��1>4�O?�&?i�a?�7?#T�>�h?�y��?i������>wJ>kn?�;C?f ?��)?�0?M�>%�R>,��䡾ǃ?���>�b;?̲?h��>R�3��}k<�~��L���7=S�սx\��){�=o��`i	���=ek>�t?&�!�	=�7�ޝ>��*?,n�>+բ>�]8���&����<)Ы>���>���>"���+n�����7��>�ۂ?��c�װ�<E (>�@�=끶�)ѯ�3��=���cU=E��:��[��K=�� >c��=�bA��ţ�L���b�<֓=�t�>1�?���>�C�>�@��-� �]���e�=�Y>LS>y>�Eپ�}���$��v�g��]y>�w�?�z�?�f=��=��=}���U�����J������<�?;J#?(XT?]��?y�=?_j#?ε>+�hM���^�������?V,?]��>��ǁʾ@ͨ�[3�.�?C�?Fba�܎�[)��v¾�
׽��>d�.�==~�����D��(���������n�?�?p/A���6����:i��5���hC?���>4Ȥ>j��>�)���g����ɘ<>i0�>��Q?�)�>��O?�5{?��[?�XT>��8�2��^љ���3�	�!>4@?���?��?�	y?Fs�>��>��)���zY��B����܂�&&W=Z>��>�"�>��>%��=8�ǽ�e���?��Z�=3�b>z��>��>��>̏w>��<��]?2?����GE��޾�j���6�<lf�?l��?�Z,?I�=2��\����DQ?� �?�ݪ?B�B?+�$�[�:v�%��Y����i����>���>�L>�P=��j=�Ƅ=+V�>�ӽ>��1��\��@��=�,?�??a`�>���雌�۵~>򻾮��=�
��Ja����z���i����5�;Kf>�۱�����s��w��$;ľ����n̾K�?�@�%~G>�3 =��)�y��:�O/��T=O$�=?x	>=���Fu>>#^�z�Ǽ��>�����Ҽ�NK���˾B�}?�1I?��+?%�C?}�y>�\>s4�I��>�Ă�6A?��U>�dQ�Yn��+x;���������ؾ�f׾��c��֟�c=>�0I�S�>&83>�X�=�m�<��=U]s=M{�=lQ���=P2�=�X�=0\�=u��=��>je>�6w?Q�������4Q��Z罝�:?�8�>�{�=��ƾn@?��>>�2������rb��-?���?�T�?C�?ti��d�>L��z㎽�q�=a����=2>���=��2�P��>��J>���K��=����4�?��@��??�ዿ̢ϿQa/>H�>v�W>�J��gA��=|������S����?ӑ3��Ǿ.�>�>eK��f��GA�=�(F>'��{d���-X�)�=�+�P�|=#�0=��>�s>���<b�Ƚ�`A>��>K"4=��>��=�����r=�hS�r�	�Qޢ>��Y>}�>��?�Y0?&^d?�@�>@�m�k�ξH��3]�>�9�=�>�>̅='�B>���>��7?�D?��K?+��>WL�=��>��>�,���m��K徣�����<m��?�І?䳸>�QN<XA�^���t>���Ľr?D1?Mj?u՞>C���4�q"��2�W�����<K�=$z�~�9���e���1�P�ֽ��=���>Wɘ>C��>��s>�xR>Z>��>;��=$Ð=�V=L��<�N�=_ޗ���=�q�E�=�f=�=/�0�9�ؼ�)D�)9��:�!�t}����=�J�>Ȝ>l��>4	�=�B��FH6>�E��%~I�z~�=������C���`�%�y�q�.��*���H>�Y>�Tv�# ��R� ?��f>))H>�C�?L�r?��%>�6�[�Ծޝ���`�#=P�^�=�B
>�=��a<�@�`���M�Q�о�b�>�Z�>U��>�I�>:�(�l�8��1��Z����P�j��>Ҭ��}�����w�����򉿼���[7r�+�"��X?k��
�~�m!w?2<?�t?a�
?���=U����y��=ԾY	]�PE�Pi�n�케�?d�?��?�\&���������ڂ�u̹>�T.��N�p��g�/��Q�=�Y̾�[�>=���Ѿd0�{L��uN��PC�,ed�U�>k�C?��?��B������|U�kd�*���T?^R?q��>��?�?��R�Ѹ���,6�=+iy?_��?;��?cǺ=a�1�<5|�Y�G>n?u�?���?-�s??߾�['?ѐY�躗>d�M��2K�1ĩ>qګ� ��<�f?+��>y$?Fs���C�N&��Į�}`!�|>�6�[=>�7=H�>�:*��(<��z=ˬD>e��={~<���=�{>P�>�����Yp)?O��=x�>%2?ؗ�>�TX=�{����<�ڇ�Ql1���.��a��n߽���<��&L=� ��}�>�#ƿ_�?f�Q>f��?hN����7�P�Q>�iY>c�^h�> 1E>�z>v��>��>�>���>>�;Ӿ �>���Uf!�--C�"�R���Ѿ7{z>����X&�o��M:��v<I��y��f��j�%/���?=��5�<�E�?E���)�k���)����)�?�V�>\6?�̌�F���>��>�ɍ>gY����� ƍ��lΆ�?p��?�;c>��>G�W?�?�1�B3�vZ��u�x(A�+e�J�`��፿�����
�����_?�x?yA?�R�<::z>L��?��%�^ӏ��)�>�/�';��?<=�+�>�)���`�\�ӾT�þy7��HF>��o??%�?�Y?TV��{����B>Q6?R�2?��s?`l6?�=?b�$�F�+?5��=TS?�u?�52?Wg-?��
?�pK>A*>.�<�|�=�S���O��aϽ
j�Y +�b=>�=�f��G�<��O=��==��᪽���6U���=�=U�=�b�=�>�]?���>�(�>R8?��.?7�%l���/?��.=�`����4������,>2k?Nū?�(Z?q�f>��B�mTE���>]��>(>	�\>rǰ>G����E�ـ�=mM>?>'n�=K4V�����G�	�ҹ����<d>��>œ>���3L">����Q��c�>�fe�ׂ��1����%�%�A�O9��"�>g;6?`Y4?r0>61��:eY�	Dy�T�?͌I?5S`?��}?z�=�<��	�N�=>3���
����>��}���揿Ǜ��D�>��ؽA�3>�᳾�Ӎ���r>PN	�[W�E{n�?N����CGw=���l&= e�2^��򨃾�L�=˅�=[ľ�]$�����͘���F?��y=�J��Mct�Eǯ�g�>0��>���>���\���A��~��X�=���>#�K>پ�����+�D�J������>�>?h2T?v�{?Y��&�}���R����?Wھr�
>J�%?�U�>	c?1�>
��䨾�[!�T�^�k[T���>#+?��1�Oy]�E�P�����F"�� �>���>��@=�?��U?��>f�\?��*?w��>5W�>Խ$|[4?R��? �H��ρ�����"M� �5���
?�?I���ܚ>)=
??�>q�?a�T?��	?��=����vF����>�ĥ>��Y��3��f�8>�cM?��?�M?�R�?T#9>�,+�罒��Y�<�p�=$��>og??�A#?��7?Lĺ>���>�󟾧d��O�>^�|?$�n?�)q?����(?�-��On�>�����>,?3 $?�Sk?�t?v?�n(?=<����6�<'���;�'>�?�|�>L��<J��=�Do�o��=p�h<��@����*��[V��f����˽��>e�w>"����`1>�,žƈ���C>>䱼f��7����8�6^�=�Ā>��?o��>e�!�a�=���>M��>� �٣&?�B?�L?46�; c���ݾ�'M�*H�>�LA?���=��l��C���Nt��e=8}m?2�^?eV�� ����f?o�Z?}N�
�<�:��v*���.���1?uޭ>�=ӽ9��>=J�?�ca?'&�>���&lQ�dL����`�ڔ׾pI�=䕯>14�q	}�{��>�N?�>��>ih>��%�u�3m�����>Bii?��?�O�?M�>��f���ۿj�d/��t�m?E0�>M�j���K?}7��SH�m��b%�n��B���lp�����;Ⱦ2�r����BW	���>�?�-]?���?ԼN?x��j�>�DZU��tS��?��.�����SE�t�W�y;a�Sk�/a�����͑��J�<�'��k�a�F��?��>2���?3�ؾ��m�2;����>
=���������=~����$�=�l�=o��N�H��w��Q�*?0H
?|ҋ>Ru?{~����r���D��un�Z������>/�)>�
�>�Z?��3�HRB:�= ����_����
�>ߕa?rI@?N/g?�&�_Q0�����o�JJʽΚ��#>��=�Lg>��i��z7��f-���E�NBv����L��>;��Ѡ=*B>?Ժv>ٖ>�	�?�p?J��,���������K�b0��S�>�-Q?���>���>L��������>&�j?��>l�>@����!��8{�9j���>�6�>˚�>��?>�`F���Y�ˎ�� ����>� ��=�`\?�}���b���>[FX?{����n<(j�>�K��. � >���>&�[�=!Q�>nڙ=��>f������,�v�g�y�p�4?�(? ���nD���=�+?�;?���>)dw?}��>2���w��Q�>�Z?��I?�F)?3g ?�i�=7)X��i����q��=�5�>��f>�n�=V?�=S��f�.�,|�qR=]�>Tɶ=K����1��8Q�c�I�)�=�P�>4mۿ
CK�ʘپ����>
��爾e���d��K��;b�����Wx�����'��V�7c�����l����?�=�?#���F0�� ������� �����>!�q�=�����b���)��B��p���Xd!���O��&i�k�e�2�'?۴��V�ǿc��� =ܾn ?	< ?ߧy?�� �"���8�T� >��<+���H��U���#�ο꫚���^?��>�
�(��k�>/��>��X>Wq>
���鞾��<��?�{-?���>W�r���ɿ���ۤ<���??�@�~A?D�(�����U=$��>(�	?p�?>>E1�/M�L����S�>�=�?���?�M=��W���	��qe?�� <��F���޻l�=�5�=͈=�����J>Z�>�k��PA�lTܽ�4>��>�"���҅^�Ѿ�<��]>��սR6Մ?�z\��f���/��T���T>��T?<+�>e:�=��,?;7H�R}Ͽ�\��*a?�0�?��?'�(?ۿ��ؚ>��ܾ��M?=D6?���>�d&���t�I��=@9ἃw������&V����=k��>B�>ׂ,�֋���O��F�����=W_���ǿ�-���l(�=�j�=��[�1�t�C�н��=n���7�#�� �<��=J��<:�>���>_�J>���>X�T?��@?�)?H.�=|����~��S߾��>�޽��Jҽ<-���*�#��-׾h��'	��$�EO��B;ў;���=��Q������!�X_c��MG�6.?�o>R
ʾC�L���<�%ɾ��������~M����;��1�$7o�TZ�?��A?�ȅ��WW����~����ۃW?�� �*C�Ո���h�=� ����=W;�>�^�=���
3�vS��J2?/?�6�g����Y�=X��o�>Zv?)�?�J��)�>7r?Y:��Z�<�[�>o03>l,�>0��>"� >Ssž}j'�
�6?Xdn?J�����G�=З̾���=�� >J�k�F��=i��>����`�c��[=c׿����Y/W?��>�*�.�荐��J���?=��x?p�?�(�>}kk?�B?1�<J#����S�O�ɟy=�W?l�h?Us>�L����Ͼ5/��g�5?��e?[#O>8$i��k龊�.��;��?{�n?W?�^��Vg}�'������6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������>�֜�q��?�R�?���m5��D'�wQ��|Y�'�H>������=�6>T�zg;����B!������2� �>� @�ۤ�
'�>V�ƾ!s⿝���^!��u"������>?5�>:��c���a���\on��H�t7��
��В�>^'U>D���,���Yw���N������}?��#�ں�>�� ������ ��cd�<_�S>c2�>�]>Jtl���Ҿ�T�?���˿���^6�=�1?�¯?�p?^�B?=�f>�yO��x#���K>.fn?���?=��?hho���B=g����j?L_��\U`���4�tHE�>U>�"3?C�>p�-�b�|=]>��>]f>�#/�w�Ŀ�ٶ�q���*��?���?�o����>f��?xs+?�i�8��j[���*���+��<A?2>H���r�!�M0=��Ғ�g�
?i~0?q{�a.�\�_?*�a�N�p���-�}�ƽ�ۡ>��0�f\�N�����Xe����@y����?N^�?i�?̵�� #�g6%?�>d����8Ǿ��<���>�(�>*N>mH_���u>����:�	i	>���?�~�?Rj?���������U>
�}?F,�>��?v1�=�N�>2�=-ﰾ��,�wb#>*�=�?��?D�M?%F�>�Y�=��8��/��VF�EAR��"��C��
�>��a?,�L?�Ub> $���d2�:!�-Iͽ�i1����h@�s,���߽c!5>��=>�>��D� Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*�[ҿXg���Sʾ�̻�ɯ>4�>\�x>���^�=� =��Լ�n����H=Kۗ>��M>�|a>�3>���=o�@>nR���U)� %��nᕿyeT�ى�����[����:E彈��8��S񖾥%.<(��a���z���?� �`�2��=�U?zR?p?ԑ ?5lx���>����t=g�#�ʄ=8*�>@e2?��L?��*?ؓ=<�����d�w^���@��Nʇ����>sI>P��>HK�>#%�>�Q9�I>z#?>E~�>H>
f'=|��k=��N>�G�>���>�z�> �}>�J>�㫿�����h�"㖾�eY�b��?0�����>�$ ��4����ǫ��q@(?2�>����̿He��9p0?�ӑ��=�:�g�m�>Z�3?�sZ?a<Y>V�������T��=cy����D�0>�/�:j��
��L�N>��5?J�l>�y>��2���7�r�P������m>c�6?�캾��:�?�s���E���ݾQB>���>�􊼞� �x��-�~�׆m��Ip=o�9?��?k���V���8h������L>V>��=��h=�B>mO���׽�W�s3=={2�=�_k>�W?{7>���=��>t����I����>�4>9E>G�:?��(?ZT�I5��}o��O%�[+x>݌�>���>3m>I�O�o��=J��>�vg>ǝ�z`i�S� �J���X>���MQx��`u�滇=o{��cV�=4
l=���F���<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>zx��Z�������u�u�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾:`Z����>һ@?�R?�>�9�}�'���?�޶?֯�?v�e>Iϋ?�Ua?X�>��Xr1�̃��̼^�������:э>��<W<���^�����ɕ��w�^��R6���>
9�=�<�>z�*��,{`=�!Ľ�U��� �N��>Z�w>�F^>Op�>m9�>��>^ �>�?�=cv�<�6��!n��!L?M��?9��zgn�FD�<�-�=&�`�(?Y�3?��]�`9ϾB�>�b\?bS�?��Z?o�>F7��>����������<�K>B��>��>er����K>��Ӿ�?D���>G]�>�A��]�ھ���R"���d�>�!!?�a�>7��=ͽ!?&�#?~�T>��>�ZH���2�H�<S�>���>x��>or?��?�����u<�O╿���ͲQ���=�"_??T?ĭ�>�x���
��q;@jͽ!q�9+t?)e?0�8���?�ψ?�w@?;�T?�r�>H�ܼ�¾f����v>��!?9)���A���&� ��J_?�T?F�>���{Qս�Լ,���y����?,\?�1&?�l��`�{þU��<����b��d<jD���>�>�̉�þ�=h>���=dm���5��zh<���==?�>��=��6�F���	=,?�G�Bۃ���=�r�	xD�U�>xIL>M��j�^?�j=��{�����x��	U�� �?��?Nk�?�
���h��$=?�?/	?�"�>mJ���}޾X�� Pw�S~x��w�c�>���>��l���E���ۙ���F���Ž����=�>u>�>1�?���>�H=>��>�!��,�'��s��M(��Gb����7p7�$�1��#�pg���}<��n �l���'|��ߚ>,�q�@��>N�?]`^>�
z>0E�>l�ԼsȈ>Q�E>�sS>^Ȕ>�D>�O>�T>��R�6���KR?j�����'�p��Q���3B?rd?"0�>i�����5���?B��?Fs�?�>v>4~h��++��n?�>�>���p
?ve:=P���M�<�V�����o6�������>�D׽� :�fM��kf��i
?X/?�����̾2=׽�+z��m�=ʭ~?D�0?��7��U�`�r�jM�ٲ_�G�<
I��]��ΰ�UEs��W��'���&焿O2���i�'?��?J�	���e;���dg���<��h�>W��>�p�>���>��s>V�7&�f�W�2�%��B�y$�>ηZ?�>&�C?��?T_j?�?~�=���>'2��X�#?��A��]&?q+l=�?P;N?�8?�+?��E?��>�S_=�r��F�?$l?q�.?�Υ>��>�^c���6cF9��<t�V���?�����c�j�]�X
��T�%h>�Y?���W�8�i�����j>݀7?��>��>6��h,��0<�<x�>'�
? J�>#���9{r��^��W�>���?%��y=��)>(�=\i��~dҺ�R�=.P¼�	�=Mu��=|;���<0��=��=h�t�7ك��R�:P"�;˯<�t�>6�?���>�C�>�@��,� �S��f�=�Y>1S>�>Fپ�}���$��l�g��]y>�w�?�z�?i�f=��=Ɩ�=�|���U�����*���Q��<�?AJ#?XT?V��?u�=?Sj#?��>+�jM���^�������?��,?I��>������������2����>�?"#j��--��	%��yɾ���C�=�a0��}�����1AM���2�*�����i>�?�u�?.8�(�EN���W���|��-s(?��>dx�=���>���N�m��':�e�f>1��>y�T?8'�>.�O?�0{?�[?�IT>��8��*���љ��C3���!> $@?M��?��?:y?��>V�>�)��FS�������%ۂ���V=EZ>�>�$�>0�>o��=��ǽ�A����>�e�=�\b>���>7��>��>!yw>y'�<��P?MI?�O���)3��Ⱦ#���뮆=���?��?.?|=%���F�3Ǿ���>G�?}��?�'?�=f���=�'?=þ"�k����>��?k��>e7�u�;>naZ=l-�>u�>�!W�=����/�c���n�%?qxH?d�'>bÿS�}��"�Tݍ���W==�2��^e�&���6^d�߼�=hc���k�.������DȾ�R��ќ��D����g>�;�?��=f�M>d��=��<������NQ=Ӑ�<0NF=9��Jb=3��U���{��P�<��l��p=��O�d�ľ�vs?G?ȗ7?��N?@��>�X@>�}ӽg�>�w�h�?��.>u�������(�{��~S���'Ҿ���f�[��
��Nu�=�T��N,>��R>�x�=�J�<3��=v�U�#=��<F�N=���=��=�F�=#֔=���=�2>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��>1l>.�C�OmR�#ݞ���ƾγ۾>i?��H�7T��>&w>>��>�,���i���=0/R>7y2�hB��yB����q=u�9��Ë<�&=īn>�~~>�a=�A-=��='�~��S4=���=p�Ľn���"�Þ{<e;=(�0>3\�>LS�>�*?�C/?=e?�>	`q�@�ɾ�g¾��>��=k3�>+�h=��>>���>�8?.�E?B�L?�G�>cC�=���>�!�>\�*�dk��bݾg����<���?��?�i�>�$�<U@�8� ��S>�kֽ�?�M1?��?89�>�t���ֿ���:"��U�<�B <�`�=vR�*h�=���<!�Ӿ����W�>��i>�V>3>��>x��>�[�>��>'��=e��=�M�=.�<���=������umJ���W>���=RH�=��=S��X��� ����<֌ͼU����=�(�>��>���>��=WT��7�1>[w����I�6��=��SB�H�c��{�4,.���7�|*A>{V>@2{�҅��*� ?`\>�MB>}��?��t?�; >����cԾ�����s�kQV�\�=^r>�=�,�<���`�%N�VҾ�W�>��>��>'r>V,��?���?=J�־��7�E��>%��F`�=�:qp�|�7��Zij�ﾫ��@?Z]���t�=
B|?��J?NM�?���>���v�Ѿ�K'>�셾�I=o�'0��3���u�?�?��>���kBA�̾
Z��!��>_7I��P�G�����0�V�����0@�>fݪ�Z�о�e3��m�����@�B��Dr��^�>�O?j�?��a�Z��0uO��������Ã?�Zg?�3�>�p?73?<��14�h���f�=P�n?���?-0�?
�
>J2A=Q���z>p�?���?�ߑ?�gz?��ľ5	�>�ಾ~��=˗N�>TG�>�9>W��>ߣ"?R�#?�-&?[ᚽ�$�A8�{%��-jB�Cp��]�<��>O�(>��=�m��j`�7
>��>��>`��>��?�"?҇�>ea��R�&�%?Yg�=��>�87?�Qt>av�=�ƽ*Z�=!��}�$�M��)���� �)�c:�#<M:=2_��> 5¿aR�?]C>�1��K�!?Ri���'�<]>PF>��9N�>�Y(>g�^>�Y�>d>�>dq�=�vj>;r>K3Ѿ�r>;��X�!��<C��R�(�Ӿ�$|>,읾0"&��'��[�I�\�������xi�m����=��]�<2��?������j��(�9K��|�?��>16?�%�������>��>)�>�4���������\ྫ��?��?�;c>��>.�W?�?L�1��3��uZ�.�u�U(A�;e�I�`��፿���ܗ
���-�_?�x?8yA?]U�<:z>@��?��%�aӏ��)�>�/�';�=?<=_+�>-*��O�`���Ӿs�þc7�TIF>��o?H%�?�Y?�SV��ڈ��#,>wV6?@*L?e�?f47?��A?�t��5?�|�<Ώ�>���>V+?��?�?9�>5�=��`>�=k����0����ǒ=lj�=�v�=���<F4��
�Ƚ���"=���<��－��:�B=�2ܼt�<�E�=v��>߮X?|�>�ѫ>�6?�!&�*1��Ч��6?t�3=C����9��8r��.˾q�>\-i?#��?�/]?l��>]^G���N��[>2B{>�ϋ>�˃>4)�>1V���� ��_,=���=�[>g&�<�v���y���V����ɚ$�j"!>�X�>�<~>em����&>�����z��&a>]�N�^���tT�xYG�v1��
w�d�>sK?��?b�=���r���Af�3(?�[<?yUN?�\?h��=�fپ�9�cvJ��S��}�>�%<����桿���T�;���^;��r>�М�����Fe>���ྼ�m��_J�{A�NTX=�W�`m^=C���о�u�����=>$>Ώ���&!��ꖿW���`I?�t=-���Z�C���s>�>�>���>��%�Hc��3?��J��}��=���>~=>>1���~=�0�D�����@�>�.C?��F?��z?�n��M~��W�L����ؾ��<�N?�>���>>�=H*�t������3s�@vZ��w�>�+?6�#��s���N��h�h�0��	�>�7 ?׃=���>�Kp?��>ɠ9?�,?�?뷌>�G��j�⾁�<?�9�?a-��q��?Pu��K���+�(B(?"N ?�|(��ѽ>~��>�ɭ>�)?C�f?�\ ?�u=�r��~ ^����>�>�> �[��7��||j=��F?���>��Z?2��?�;M>�e(�1�žC�d>>`Ţ>�P?�K0?=?�c�>��>����~*���Z�>9�?���?�<�?�$�<l/?�YI=���>�X>��>�?O�>a}J?�5h?S�S?.?@ܑ<�,�0�K�ǽ4M�3�E=�t=���=�@c�;������F>l�=�9o9�Q����;9r���	=��+=�h�>Lt>�"����0>t�ľON����@>[������ ��l�9����=V�>�?oٕ>>#���=�ϼ>�J�>����(?��?2 ?g#;{�b��ھ�L��>A�A?e��=��l��t��'�u�(�g=U�m?�z^?;pW����qd?�^?\���t0A���¾;t}�yP꾷�R?�5�>HvG�ɳ�>��|?��b?A�>#XZ��m�Tl���x^��@���;�=��>9���d�x�>�+-?
x�> %\>�	�=�9ȾDb�a`����? ��?��?=�?�a*>��`�^࿟E������g^?3��>劧�4L?[{>��/ϾQV��Zą��g㾔R���h��񚾡���fr*�$���<��`z�=?�p?��t?�_?\���I�Z�!�^��t��[�� �=��:�D�̋D�*qH���k�����������.=����fO��n�?O�?J��??�ù�����2*�"�>Eĸ�(�x��e>��E�Oim=� �=�V��S��{���?P�>��>�B?�	p�N�1�Ef8��`C��Z��2�/>/g>��{>1�>�o��@^�z��������>���w>]�c?��J?ىm?\��s>1�)���.x!�P�7��C���Q>>��>Ŗ�>��]��"���&��?�6�r�;)�`���x�	��|=��2?�z�>�˜>͘?�?�o	�Q����z�h62�5�<��>��h?���>}��>��н���G_�>NLp?��>�*>�S���?'�و�=��=�>!��>�q�>�9>�l�N%o��Z���n����Q����;��;?B���]�h��fu>h�U?�ǉ���f=#�?l ����B�
����R��ݯ>��[��k�=S��2���NM�<굼�3.?d�?뚲��32���Z> +?!�>s8�>Ie�?O1�>�|��[�k;��>z�`?�/O?�>?��>�ɱ=�>�����m�3�;"=�Ŗ>�ǁ>�I�=bO�=��M�ҳG���C�o��=��=:n0��#��O���ͅ뼆�=+I=4@H>xRۿp|K��qؾf��?E�O
�j���9������G���>��jj��-s�\��h�,�9V�q'b�p����k� G�?���?
���∾/6��3��T�� 5�>E�w�7�{��p����S����*������!�]2P�'i�^e��'?����C�ǿ󰡿a9ܾo ?q4 ?}�y?5��"���8�^� >�D�<K���T��;����οV�����^?O��>�����E��> ��>#�X>4Oq>E��!ߞ�&�<c�?Ax-?V��>�r�+�ɿe���Τ<���?��@�~A?-�(�n��HxT=#��>�m	?r=?>�<1��N��հ�o<�>�>�?P�?�K=��W��T
��Pe?���;�G���ۻ�L�=�)�=�>=�����J>:A�>I���A��V۽�4>՚�>��!�u���^��ʽ<2h]>l�Խc��/Մ?{\�xf�y�/��T���T>��T?�*�>;�=t�,?"7H�W}Ͽ
�\��*a?�0�?��?8�(?�ڿ��ؚ>��ܾx�M?yD6?���>�d&��t����=�6�T���C���&V���=]��>.�>҂,�ϋ���O��F�����=�z��B����g��� {��C������"��Z��[�K=�S��P�N�ҁ>["�=�O=��4>	Z�>���=��K>p\[?��T?�;?#Ch>Y+�-"�?�ﾣv>P��My��Ұ�����?"�g�'��V�n!�4�&��/�o�ȾM�/����=KBQ�p}���5��od�+�E�.2?��=C�Ⱦ��E�ա=��Ծ.3��Qh����ֽ6�ʾN�0�7�r��ɝ?A�C?#-���iZ��P��#m�Ƀɽ޼P?'��.A��Ƈ�'1>��༧��=���>1z>�L־�")���\�ܻ2?�/?������Rn>x\��ޏ�=�?/Q&?�����)?17�>u��>
��>��>F+?��?-�B>�ݾG&j�)�Y?��n?�k,��wq��A
>Δ#�a-	�Z6=k=<>A���?�=��=�Ä=C�񽃧g<�ȉ��L�=)W?���>��)�d�oa��w+�`.==��x?�?<+�>zk?��B??p�<�e���S�~��Yw=��W?_$i?+�>����4о�y����5?�e?�N>�yh���龩�.�MR�=?f�n?�\?�Ɲ��u}�|�����o6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?w�;<  �S��=�;?l\�>��O��>ƾ�z������4�q=�"�>���ev����R,�f�8?ݠ�?���>������� >�r����?���?P,�2)�;�%�l�]�R�	��5Y>�Ec;4$'�"�!>ob�Y��ޭ����/����;��/��>��@�gʾp?���rF𿤖¿������
RT�]D.?��>iZ�*ξ��w�q�k�B�B��`n�ЁY���>�7>��ܽ
��_%s�f�?��D+��:�>:汽%�w>��:�i���Ҵ�s�:�ɍ>�>�)v>a�̽�oܾAՖ?"ؾ.�ɿf�����kC?��?��|?6�?�=���a��<�Dy\?]�?�m?���e'�I��$�j?�_��vU`��4�rHE��U>�"3?�B�>T�-��|=�>���>g>�#/�x�Ŀ�ٶ�B���W��?��?�o���>o��?os+?�i�8���[����*���+��<A?�2>���E�!�=0=�MҒ�ļ
?Z~0?{�i.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�+�>%�?�Z�=E�>N�=0���%1�$Z#>���=�H>�Ι?֫M?{C�>���=�!9��/�bF�vKR�4*��C���>[�a?u|L?�,b>�฽��1��!�)Bͽ�/1��U�>�@�l",�,�߽��4>Ŷ=>>��D���Ҿ��?o�q�ؿXi���m'�i44?��>.�?(����t��Y�$:_?�v�>8��+���&��PF�u��?7G�?��?t�׾�h̼�>q�>aG�>-ս/���+�����7>��B?7�~C����o�e�>���?�@yծ?�i��	?���P��Ua~����7�C��=��7?�0���z>���>��=�nv�ܻ��S�s����>�B�?�{�?��>#�l?��o�Q�B���1=#M�>��k?�s?So��󾞲B>��?�������K��f?�
@}u@]�^?1��Ͽ�������n�ľ=u<><�a>��K�v��=���u+2����<�g7>���>��B>U;c>�Z>�e>�8?>������(�2V��Ǥ���Y�,^���������	�<�����Į��ۇ��Z<kw��p�<�y\�J�P������=3�U?�R?gp?�� ?e�x���>���1:=�#��˄=</�>�h2?�L?\�*?�֓=w���A�d��`���A��ɇ���>�rI>��>�J�>}%�>�rO9��I>1?>��>� >�d'=8�亖b=�N>�M�>���>)|�>c4=>�s>~���)1���vh�x��Qͽ1��?�+�J�����$���
��B7�=OA.?�>�����п����H?z���5��J,���>3|0?�:W?�x>,���wMQ��y>�	��`j�*H>-����j��k)�(AR>?�ni>�y>�3��9��P����� �q>}�4?@���ja2��u��vF��}ܾ��E>m@�>�h�������V���h��Vz=�:?��?;���j.���8s�5A����T>�a>݅=H��=s�P>z{_��н�M�r ,=���=cb>rp?:�D>6��=;��>.[����T���>6�&>�AY>��6?,4?��{�-���o��w �]��>/g�>�ϟ>In<>��M�K�=O��>7a>�3��쥼�� �-wg�߱X>�̌9�Rm�z�d���B=�ŽX��=P�=2��{�O��$C=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿi�>|e��V��8���u���#=��>�=H?Y��9�P��B>�El
?�?:q�򧤿S�ȿ}v����>>�?��?3�m��>���@��w�>��?]Y?�wi>/b۾V8Z����>4�@?�R?�-�>�+�ha'���?Zܶ?���?�ˇ>�G�?S�N?��x>�M���"C��ۻ�e�w�� [��=xQ{>�	�>��Ǿf2Z�6Ք���t�[$y�F!8����;x(=���>�;Ž}���.(�=�<<���Uw½*�>B�>H��=O�>}��>��>�sT>9���'�����T���K?���?y��X3n� C�<���=a�^�	'?vH4?]T[��Ͼ֨>o�\?���?	[?c�>+���=��5迿�}�����<��K>P3�>@G�>*"��HK>��Ծ�0D��p�>�ϗ>n���>ھ�*���*��B�>le!?4��>qծ=gM!?&a#?��P>��>W�=�C"����A�ms�>��>��?�l?}�?��Ǿ!38�-x���9���{X��Q8>�r?Y�!?1��>3$���➿Z8��n��]>ǽm{?�PY?�!���#?9��?�`=?VSN?킇>K�;�pҭ�_a��P8>��!?_d�G�A�o&��N�tU?�@?.9�>���Y�ս@�Լ��"���� ?�1\?Z6&?���[�`��)þ���<�{�J�l���;1�F���>��>'D��ꇵ=-�>Đ�=#m�@6�]�n<`�=z��>�x�=.�6�d%���<,?B�G��ڃ�G�=V�r�qwD���>tGL>������^?&f=���{�}���w��MU�� �?��?Vk�?E����h��#=?��?Z	?�$�>�H��m~޾���-Nw�|x��w�J�>���>[�l��}���B����F��Y�ŽMJ׽�e�>�Ѫ>T??���>�Q>�I�>��x�-�o}+��~4��xm�n�9��=Y�7�:��]\�2���w�u�>m
��Y2��BRs>/���G
�>P�? ��>궻>̿>����^>���>t�`>l�>�M�>T�=脈> ��=g���IR?����T�'�]�����47B?�td?�+�>n�h�Ɖ�����Ȃ?#��?�r�?�<v>6{h��)+��p?fC�>���p
?�Y:=�3�}�<�R��1���0�����ϩ�>�J׽[:��M��rf��i
?�/?�$��*�̾}
׽���=�=��{?��2?0+�s�V��7z��wU���\��N3=��:��z�qD��Zm��^��A�|�S���-8�����3�(?�`�?���)��h��`q��H��u>�i�>�Kl>���>�>b����0���e��`$�%�N��t�>��Y?�V�>��B?�E7?ŶY?sF?7��>wù>aľZ?�s<g��>,�>Ĩ?R�$?/c.?d'?b#9?�T�>4�ڼ;�&;ھ��?K�?ӑ?���> @?�?p�pt�<[$�����k��Y��R�<�қ�d �G�e=nRC>�G?����8������k>��7?���>���>����H��1*�<�[�>��
?aV�>I����Ar��>�A��>Ӷ�?gk�W�=��)>���=�+��y$Ǻh��=�w��N��=�灼�C<�� <���=[f�=�n���8H��:A��;��<�t�>8�?���>�C�>�@��/� �;���e�=Y>S>+>Fپ�}���$��G�g�"^y>�w�?�z�?��f=i�=��=�|��sU�����������<ԣ?.J#?-XT?Q��?h�=?@j#?r�>+�[M���^�������?�u,?���>���l&ϾT�����3�n$
?+�?ԗ`�+����(�c^���ѽZ� >9�1��I}�W��a�D��7{�L���V��d��?!��?��h��3�`7�=�������8�D?6ƽ>�W�>�*�>`�'���h�FV�^E:>�/�>8�R?<'�>��O?�7{?��[?c`T>��8��2��	ҙ���3�">�@?���?]��?�y?�d�>��>2�)�� ��Z�����	�݂���V=\�Y>��>�&�>`�>2��=��ǽ)y��V?��r�=ʅb>���>L��>p��>�w>���<0�W?x�?�~�<8� ɾ�A��ʨ�<�?3�?L?!j�=J|	�, P�/|���?���?Ql�?�=?U�^��/�=7� �&����S�X��>L�>���>� ��!>➷<5O�>*p�>?A/��8龾}-���P�	G?�;:?�H>d�����s�7:��e���:j��t�3hm���1�sԫ�>�>����d��J��E���������� ���Φ��y�Zh?9��=EN`>���=�k�<*I�=w�:�D>����q��=4t�������Y
���-����<�;�ϫ;Q:�=�2O���˾�}?�;I?�+?��C?�y>�M>;�3�'��>A���28?�V>��P�ҁ���;�_������l�ؾ4m׾j�c�<џ��9>�oI�b�>�:3>#Y�=
��<���=�$s=õ�=��R��R=S=�=[Z�=$?�=���=��>�T>�6w?R�������4Q��Z罡�:?�8�>n{�=z�ƾc@?��>>�2������qb��-?���?�T�?A�?1ti��d�>R��,㎽�q�=5����=2>0��=��2�T��>��J>���K������4�?��@��??�ዿ͢Ͽ3a/>.�R>/*>��N��~6��*]�O���r��do?�=�+j��m6�>�h(>����׾�a�;g�,>�]�;�QK�rd�(^�=|-�)R0=3�<iL�>NU>=�=�Խa��=	g�=WӲ=��>`G�<�����<�=�^�=�p�>�/>,��>��??0?�]d?͹>cn��zξ�!���ٌ>Q�=y�>���=.�A>�¸>%*8?��D?dL?-2�>�O�=��>ߦ>V,��Nm�}r��䧾"4�<�j�?��?�$�>�S<��A�ǀ��t>��gǽ-O?��0?u�?&�>C���KݿȖ���'�������5�i��=F�����e<E�ȼ�@���ߕ=y��>gd�>�e�>��>�:v>	<�=�h�=�|�>OqA>@F>b'�=�8��;h��Y�$Ƽ���;�.!>d� ��E�=}Z8>&b�����<�s��=�Wn��W�& �=b��>�>��>�}�=/����,>�ݕ�_�L���=�e��C�ʖd�����/��4=�f;>J�R>��t��䑿 j?M<X>�?A>"��?ku?�'>����*־ '��Q�i���T�~�=�y>��7���<�$�_�G^M��MϾ�d�>]��>���>	�I>b�(�|M>�μ\�Ⱦ�8���>_ož�fE��!v�kl��������A~���o�J?�����&<�\?�YI?<�?���>�A>�3�>}�=�_��,ȽQ���a��V��i'?c��>[�>��徏r�ۤ��W7�ra�>T,M�f�:��Ŏ��'�Z��=�ľQ>>�Dݾ�+Ͼ�N=����y����h�}���<L�>�(N?��?%��fw|�Z�Z��������X�>I�W?�A�>-�?@�,?�vT=M����୽��6>M�?�?|�?L!���x�=��^Y�>�7?f/�?�?���?�|�� ?���������	�=6"S>�H��{>Yo?>�?� ?[߁��4�9o��b:۾_��{�>K�7>g;�>h�=�y> =��=">�Fw>��>1��=�C> �>��>s���$� eS?u��=��
>Q�*?�C>�(1>?q��F�T>g��^)����m��*+g���
��P1<�b˼�X��g�>E5��-?�e=���۳1?����l�%=��>�R>fʽی4>x=X=��>�{�> D�>��=��>H:E<ʪľ%*>^|
�?%�&C@��1S�����h>���q��4�0���AD���V3��	h�����֭?�6!���o�?�����c��$�&?�0�	?��>�++?S���S�x��=D�>�y�>C�������ɶ��+"ܾG�?�t�?�;c>��>P�W?%�?��1�3��uZ�"�u�P(A�e�E�`��፿����
�G��)�_?�x?'yA?�S�<$:z>C��?��%�Uӏ��)�>�/�&';�@<=x+�>*��`�`�}�Ӿk�þ�7��HF>��o?0%�?ZY?hTV��?�>�48?�S=?@ �?��9?��A?�y��)?+9	>e��>gE�>�x.?�e,?0��>0)#>9��=�X<'ؠ=���������A��C�#���a=��=ڤj<�t��!�x=<�=�lݼ�?��GY�<�<iɘ���=?�=Nm�=�F�>�P?�P?�=�>��$?���rnԾf�̾VX?6[�=(� =��þ_����B��a�f>��y?���?@rf?��>^�J��VT�T�Q>�>Q��>�[�>�.�>����Q9�u�=*uj;��>��r=����8׾�����&8��-%>M��>�8|>Z���'>�z��e1z���d>��Q�ѿ����S���G�h�1���v�1]�>d�K?�?�ʙ=�Q�����Gf� ,)?�_<?�NM?��?�=��۾j�9�E�J��6���>�/�<%������o"��m�:��ޚ::�s>�+������6tb>��'-޾ �n�U
J�����L=%��4V=���6־�B���=��	>M���� ����7Ϊ��J?�0k=�^���U��#��1>$��>�>�M;��Yw�!~@��Ŭ���=^��>IO;>�����XG��B����>�RG?X]=?�e?�JD��:i���1��Oþ�@��� ��j?�	>���>��=��>�&ܾ�#�6M�8V:���>�$�>6�-��X���ּ'`�:�:�>u�?~�>hl3?R!w?9�?��j?��?h�?��>��<�ƾ�0?�!�?�&���V�=�.�K4���?)?������>)g?�f�>��?�Wi?b�>��>>O���_QC�5ˊ>��>
XJ������r>tY(?��>d?�"l?�r9>�y���u�ew���>(�>��G?<�-?��!?��>P �>`���G�
�J˦>5ǆ?Um�?���?��A>�s?�1>>
?��&>tі>�{�>K�?�(??V�t?�_k?w�'?	/=��y�1�~T8��2<���F{��{J�<e��v���M=HdV=��=jd�=i�����颳�B�z�S�<�_�>l�s>@
����0>,�ľ�O����@>�w��O��Tۊ���:�ݷ=5��>z�?ī�>�W#����=��>>H�>���e6(?Z�?�?\n";]�b��ھ2�K�%�>�B?X��=��l�F���f�u���g=�m?��^?��W�?%����b?C�]?�u��=���þ�b�А龈�O?	�
?_H�M�>"�~?��q?���> �e��-n�Y��4b��k�� �=t�>�_���d��i�>��7?,2�>Z�b>���=e\۾a�w����	?d��?���?���?.q*>�n�D+࿁S��M6���o^?<I�>����g`#?�p�Nоx����䎾������奄�a��X����!������ܽ�˺=�?ss?��p?(k_?��O�c���]��5����V�x����D�E�?RD�8C�{+o�o������R���3G=U��LO��v�?�K?c����Q6?6(��>�p�澓K=�P�Ӯ
>a`�>i4>1=vYe>������ݾ}S�?^.c>D�?��%?8�+�
���F��1�,�� ��S>�G�>� �>�>�D��d�Ѷ������i"ξ��⽅7�>�3[?I�1?Qc?I]�#�6���h�̼���N��	���'�<�gq� A[>��˾��@��<��[;��|n�����`������[=�#?G�r>߂�>Eԝ?��?����������!,N����>La�?��>�e�>k`,��8��C�>�jf? ��>�`{>U���>��{�N���\�>[�?xq�>խ>��$�Rsy���������T��B�=��g?�����p~��/(>H�F?��彩�=e��>�����Ͼd�3�sLȾb��{��>P}:�YK�>�FӾ��i�u�/�ʽ[c*?�?����g/���>z?�!�>�#�>�V�?�>�>���`M<�?�^?~�M?,�C?!�>�ԏ=}J��C`ͽ��)�L�==ȣ�>��K>}fp=lj�=�m���C�@H���2=Þ�=�A��O��Q6�Ւ�Π=�#K=!B>e�ؿ�jK���Ǿ3�������j�S�^Iս��Y��VM�T�ܾJ����D�m#w��t��pL��M��&{��V�C��?�x�?�XĽBm��䤿��p������>����uT�<a;�;�� ���W��	�������c��C��
u�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >[C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�{A?i�(�+��XV=���>��	?��?>�M1��E�����hW�>�;�?���?��M=��W��	�)~e?�<��F�.ݻ��=�7�=�3=�����J>�Q�>I��VA�f4ܽ�4>vۅ>�s"���P�^����<H�]>��ս�7��5Մ?){\��f���/��T��U>��T?+�>v:�=��,?W7H�`}Ͽ�\��*a?�0�?���?)�(?0ۿ��ؚ>��ܾ��M?_D6?���>�d&��t���=�6�2���~���&V�l��=Z��>i�>Ă,�ߋ���O��I��N��=I	�Ŀ3�!�Fs��|=���<�n7����|R]���ʽ����@|�9�ѽ�`�=5��=�A>V��>��l>c>��Z?��q?z��>�J>� X��9��)羿�
��燾�6	��ƨ���w�(�뾳Nľb��1T$��:(����T�<��.�=�1R�����9� ��b���F�\�.?m�$>�'˾��M��&<��ʾ����qʁ��z���̾Zw1�cn����?��A?���hW�D���/��Ǻ�#�W?��X��;\��N{�=�,����=�2�>�I�=�X⾩�2�i|S��53?�l*?+C߾�AȾ^o>��'���=qB?��'?� �3�> ?����u-�<��>��>�#?�z?�?>Px��:�L��+?�}f?�����^�"Ӱ>���}�����<�_ >]؈���8�Q�>)j`�屁���>S̆�HE= W?��>��)����������q==q�x?c�?���>Ytk?I�B?]�<�X��F�S���G{v=��W?[%i?��>����c�Ͼ�o���5?G�e?�N>�Eh�s��7�.�qO��?��n?_A? V���T}������v�6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?w�;<��T��=�;?l\�> �O��>ƾ�z������4�q=�"�>���ev����R,�f�8?ݠ�?���>��������=*3��p��?��?���M�>*/���������&>X��=��<k7�=����}eQ����E=�(�ھi�úuh�>��@㜦����>�fE��9�O���Ґ������m����?9M>q���^�ϕw��L��[�2���U/3��f�>cg>�P��<���{��j;�K���&�>Ь�_l�>�eS�����%/<M�>�)�>7v�>��.뽾��?����;ο�������X?�'�?uT�?�v?��9<Au�ɔy�u�"IG?�ds??Z?b|"��y\�7�9�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�g�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*��+��<A?�2>���I�!�C0=�TҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�$�>��?	o�=>a�>Nc�=V�2-��k#>��=�>��?�M?VK�>T�=��8�k/�o[F�CGR�8$���C��>�a?g�L?`Kb>���2�/!�OqͽWb1��c鼩V@�c�,��߽�&5>I�=>&>�D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�c��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B�}�1=9M�>Μk?�s?lQo���i�B>��?!������L��f?�
@u@a�^?*�vԿ6n��N�޾�뿾�U�=Oe�=��><)�v>��%=.]����;��>� �>U�.>��>�@�>�.>�Y�>�H��P�!������Β��dN����G'�`�_��i�Q��w������-����e��pὫX���}��GK�e8>��e�=�M?"�T?{�q?T:�>�&ü��>u��	�;�11��3-=��>(�9?��M?X&?z%�=I����d��͂��ݟ�!񎾔Y�>�jK>8�>4q�>���>�<��J>��1>ie�>�>��@=O���U�<��Z>#��>1(�>�4�>�C<>�>3ϴ��1��Z�h�w��̽&�?~���_�J��1��:��覷��g�=Fb.?:{>���?пY����2H?����q)�H�+�K�>u�0?�cW?@�>���T�T��:>޿���j��`>+ �l���)��%Q>fl?�f>��u>�M3�| 8���P�Z����}>�6?��@;�!v�@�I���ݾ\J>N��>��|��j�+얿��~�;Gi���}=s*:?��?��8���Yu�zz��w�R>j�Z>�J =wD�=L"L>��W��?��wJG�-U,=s�=��^>zg?(H->��=kM�>�1��d�R����>(�B><{*>T�@?[%%?4��������p�0� �u>3��>d�>�>�<J�r��=Z��>M�`>���ł�$q��>�6Y>��w��ra��
s�*+�=�ۚ��|�=���=���$`<���6=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>vx��Z�������u�l�#=Q��>�8H?�V����O�e>��v
?�?�^�ߩ����ȿ5|v����>W�?���?f�m��A���@����>:��?�gY?roi>�g۾;`Z����>Ի@?�R?�>�9�w�'���?�޶?կ�?|w�>Ek�?(�P?`�>M�R"J�vH��&or���	�lxd>���>�l$=��Ծ��F�ni���I����g�0��`��<�&�<��>,��U$�4E>��̽J����f>^]�>\��>l��9CF~>� ?z�>��>��=mk��,��X�+�s�K?���?����7n�+��<�h�=^�^�.*?gD4?�q^���Ͼ(ݨ>��\?��?K
[?e_�>4���5���俿�p����<x�K>��>�F�>{��XK>��Ծ�&D�}n�>�>Z'���=ھ�
��T,���R�>Ri!?��>BԮ=^f ?"�#?	�g>@|�>��C�Yґ���E�l��>���>҃?ԙ~?�?Bs���L3��𑿋���־Z�VAI>.u?�?XN�>Û��kŝ��� ;�k�)����E�?3�e?a	���?[݈?ä<?s�??�f>�ɓվMh��b�v>��!?y���A���&��
�"*?�?�F�>nAؽ�FμH�������?CV\?�&?S�l�`��>þ>��<%��s�8��;ΩB���>C+>���	��=�>�=�l���6��y<���=���>��=��5��.��0=,?ܾG��ۃ���=��r�<xD���>�IL>�����^?]l=��{�����x��	U��?��?\k�?L��?�h��$=?�?Z	?k"�>�J���}޾G�ྵPw�-~x��w�K�>���>�l���H���י���F��j�Ž5���~�?E�>T��>�c�>� >�ܽ>�[N�fs��E��K(�"������t�P�#����C�������}�����z��v�2���>�R�Z��>�#
?12;>���>��>\ý�>�	K>�)>u��>菱>~nA>^E�=ޣ�=�����KR?����3�'�}��y���x3B?(rd?�1�>;i����n����?���?As�?i=v>�~h�y,+��n?Z?�>��&q
?2U:=�7�#8�<V��7��\3������>�C׽� :�IM��lf�Fj
?�/?,����̾�;׽$f���=3k|?�5?d�1���N�'�v�Mnd�&M_�"	�=8��.픾u�M]e�!C��������y�q�&� ��<�"#?�"�?�[��"�\�������}D�[��>��>`�^>7=�>�e	>��(�	7A�-�5�V#1�$�����>�E??1��>H�I?4<?:wP?�kL?˼�>Nd�>#2��ho�>u�;l�>�>��9?��-?K80?B{?8v+?�8c>�{�������ؾ�
?h�?�J?�?!�?�����pý�����g���y�3|��M�= �<S�׽Du��T=O	T>�W?�����8�����8{>��8?���>+[�>���PK~�%x=��>�6
?���>{����p���	��U�>�܃?����h�<�e+>�a�=� ��:�K�b8�=�D׼灆=���='���<�w�=";�=ջ����8'@����:v�<�v�>�?���>�>�>�@��j� ����Fg�=��X>�GS>v">�Eپ�{��#����g��Hy>'q�?w�?�df=��=ڥ�=y���W����������<ݤ?�L#?�YT?#��?#�=?�l#?i�>�,��G��=_���	����?u!,?��>�����ʾ��؉3�ѝ?g[?�<a�����;)��¾�Խ��>�[/�j/~����:D�������B��/��?濝?�A�M�6��x�Կ���[��t�C?�!�>Y�>��>N�)�t�g�k%��1;>���>oR?9��>��N?Q�{?��[?2�R>R}7�������+�=�9!>�??T��?� �?��x?k��>�>q+*��K�}}���0�)A��@��I�U=��Y>\ӑ>$�>�R�>���=��Ž�ﭽ�s>���=G�a>��>=��>x��>F�u>Џ�<ɓK?1D?�#���E8��D�KL���<$��?)5�?KF�>�6�=�FԾW�\�ހ���p?�?�S�?@�P?�u���4"=���yf~�7���Zg>-�>@�>w�޼��\>g�*>�T�> `>3x;���˾�5��K�<A-4?9�G?�-D>;�ſ�q��m��d��1�Q<�K����e������}[�S�=�������,��XGZ�6~���U�� ���g�����|�T��>v{�=��=E��=u�<�ʼ���<7�N=�ܒ<��=o�k�ryo<-�=�4wջS�����%��E\<f�E=�Xͻ,�˾�}?�;I?ޕ+?��C?*�y>;>ڔ3�I��>�����@?uV>�P�������;�G���� ��S�ؾ%x׾��c�ʟ��H>�`I�)�>�83>�G�=oL�<?�=�s=�==�Q��=$�=�O�=�g�=���=��>VU>�6w?W�������4Q��Z罣�:?�8�>p{�=��ƾo@?��>>�2������vb��-?���?�T�?A�?;ti��d�>O���㎽�q�=G����=2>x��=��2�T��>��J>���K��:����4�?��@��??�ዿϢϿ2a/><H>�z>�S�?�4��1�&j���c�"?�4���Ӿ-��>F�=���/���?Ċ=b�2>8?s=��ƹ\��b�=��Y�E�<D��<Վ�>�WD>��=a�����=+`=���=(dn>� ������vP�Jc�=�8�=��f>;� >ܒ�>��?W0?Jd?�9�>�	n��ϾY+��wG�>��=RI�>���=z]B>�>e�7?-�D?!�K?l}�>�w�=�>?�>l�,�c�m�,=��ȧ�1e�<œ�?�ˆ?l͸>�U<X4A�x��2T>�RŽf�?OT1?�j?M֞>ԃ�bK���6�i�2��H���:fz>Ep��� ��>f��V;���=�kJ>ZX�>�z�>���>�]>���>\��>H�=�\V=d�>誳=��=��4=ˋ�=m{��+,�=����{绚O����!=�c��聽$��<!�<��=�-�><�>���>X��=aҴ�N0>
���[L���=;˪�D�C���c�#m��k.���=�R�?>(*S>j���eΑ��,?�!Z>�2=>V��?�yu?W%>|1	�:-־�^��u{g�
Y�c��=t�>32���;�n�^�ǈM�!�ӾR��>�Ɛ>q�>Kn>:�,�S&@���f=F��3����>z@���K�����t��Ǥ�ֶ���}i��?���tD?�Z��`"�=Nz?�{I?i��?{�>@\���վm�/>�����t<r��`�p�m���`?��!?��>p3ﾒ�F�D̾��ݷ>�<I���O�%���0����gͷ�F��>.���#�оn$3�@g��������B��Or�c�>g�O?z�?&1b�X���VO����_4���m?K|g?.�>wI?�B?����x�!o��Xx�=��n?��?u<�?��
>�'�=KF�����>�?;ۗ?��?lv?�W8�mQ�>!��;�'>����V��=�$>��=���=�(?8�?�?T���)�	���B��&^����<<9�=wؐ>.#�>+Qt>�Q�=;u=�}�=�a>���>s�>�&`>=ţ>I �>�g�����3�=?�|h>��@>�dM?�"'>�jl�%��P:�#��_{��4K=?��(�×B=�	���6��k�QN�>�9�����?��N>���4c?%��zЁ=�\�>(�J>&���A�>���=6F?>��>&��>]3/>��> �`>t9Ӿ��>����a!�H)C���R��ѾA{z>����b�%���ۄ���FI�Ar���m�;	j�_.��>6=��B�<-D�?ϣ���k���)�p�����?�[�>�6?�Ɍ��و���>���>�Ѝ>L��#������q���?=��?7Fc>G#�><�W?��?1��%3�NmZ�#�u�	A��e�#�`��䍿ӛ��~�
�ƿ�T�_?�x?�pA?k�<�Ez>i��?@�%��揾 T�>_/��.;��3<=;�>a$��Œ`��{Ӿ�þ��fAF>��o?�#�?�]?�[V�m�o���">��;?�2?8,s?��2?�:?��B$?;:2>��?��?ޯ5?��.?��
?�6>6q�=ʃ�5�!=�f���Ŋ�K
н
˽�}�-=��=��C:�<9� =�׭<�����S=;�x��=��<P8=��=���=�~�>�]?٩�>n.s>T�7?9���!-�����Q;?A=�p����)����[־e�>�n?�"�?e�b?��m>oIO�|$\��>=��>&>^md>��>�,/���2����<�~>L��=-��=�Ƽ5���ND�k���!��<C&>��>r0|>D����'>�|���0z�s�d>��Q�^̺���S���G���1�5�v��Y�><�K?��??��=4_龲,��gIf�.0)?�]<?�NM?��?�=��۾��9���J��>���>�X�<��������#����:��N�:��s> 2��-נ�d_b>��>l޾�n�J�����3M=�����U=��.־m<����=%
>������ � ��8Ԫ�-J?��j=2k���GU��i���>���>nخ>��:��
w���@���V�=ӱ�>	;>n������|G�;�[֧>�eU?,S4?�*�?�5Ⱦ�ڂ�w4c��1.��=8�D���c	?D��>a��>�I�8��{��/#���b�wp���>H��>�O���^�Q���O��� &@��R�>�4?��5�N�)?-.r?�g!?�q?��?ޚ?��>ÏϽ��վ/M-?N��?��#��y��]�� �:��c�z�>�C?<��((�>�+3?��?V>�>p�?j(?�>��S6j��^><�d>R>+��5����>�fD?b�?�pi?��n?TI�>�7�0����=?�w>g��>�KH?'�?��?lI�>�+�>嫶�'.���&>[�T?_bt? wf?<��>wT�>�ͧ>Z��<Õ�=��?�/?P�>0G6?��?�?%?d�>ب=�����⎽	ļ;�B>��������Y�1rN�䃉���I=y�=}�>1Y;��V�,d�����=��.�������>Mt>K��� 0>��žC҉�m�>> ��-Ϝ����Z8���=q�><�?Є�>�$��i�=`p�>�[�>f��?(?�?�?{�	;Vub��.۾w�L�].�>��A?w�=��l��9���v��&q=��m?b�^?]RW��{��H�d?~�[?3z�>�@㾤f��{����iP?U��>�Cp����>��p?�_?c��>8〾
\m�(���M@k��M�Eǘ=���>ګ���R���>��,?&8�>��f>!�=�n˾!q�+���T?���?��?�?~W>P�h����Ֆ��Eɖ�G*z?Ng�>+�h�xV$?(�G�q��l��)�h����|��ꜙ�����ם��{��1����O��<�I$?�Dl?�Gb?�=N?���Ra��y\��s�9\��.׾���@MJ��M]�IlG��(m��2���,��D���l�=�����O>��6�?� #?ˑ����>�,��r ľ�ݾ(.>������eݺ=�Y�{2N=Y��<�l�Ԭ-�������&?nl�>��>y;?
lG�H-<���)���1��_��h;>�$�>��>�6�>�=��I����V�[b����ѽ�)>޴d?��F?�n?
�
��2��d���) �bH!��泾��<>��	>���>?;n�K�$���#�$�<�;_t�l���F������=�*0?��>��>�2�?�[?�h�_穾	I���0*����<���>=�g?OW�>���>�T��f��q��>ok?���>f:�>�땾���)�x�2��#T�>�ʚ>L?kK> &k�H\�mN��m򑿾2D�x�=NHp?�wv�ds�A
h>��H?�ґ�xYc<++�>�X4�7�*��.�f��5�=8�?��=e�>���b�����Y탾@�?�F�>�\k�}����7>�?+>?��>;�?Ĝ�>���a����?��g?ְA?�7*?�@�>z�=�;�ͽ�U�r; L>�rO>!_}=�|A>+�*=��+�������:�,>��%k0�j"�<���=��#=�����M>�)ۿ3�J��9׾�5����*E������լ�?s�����>������	w�{*�M �T� �b�y���-Ap���?�?ꌾQ����*���C�!���y��>;y��=���Ҭ��}�n����۾�����"�"�P�[�i�[f�b�'?Z����ǿ����;ܾ! ?�A ?	�y?��H�"�v�8�{� >�9�<@0��O�뾺����ο�����^?���>��60��?��>~��>��X>*Hq>B��鞾,�<��?�-?W��>ˍr��ɿ5���Ƥ<���?�@�aA?��(�q��W=�n�>V�	?-@?>�~1���������)�>��?��?O�P=Y�W��
��e?N�
<y�F������=��=�=���j�I>JE�>�K��a?�^1ܽ�5>q4�>�!'���Z	_�pG�<[�]>>�Խ]���5Մ?,{\��f���/��T��U>��T?�*�>V:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?_D6?���>�d&��t���=T6�҉��}���&V����=Z��>a�>,�ߋ���O��I��U��=<r��S����nO����=�O=�Kl�^�A�R����-���p���J����佌tY=$�>c>��p>yP>�>�NW?�:z?�?��>���X�@�!,޾
�ս�}��b�8�^������r?��|ǰ���־�����.���$�k��z=���=w8R����w� ���b�D�F��.?|j$>��ʾP�M�2F-<Auʾ����t���
����3̾M�1��n�|˟?>�A?G����V����Dk�	����W?wT�~��款a��=b(���=�*�>t��=��⾥"3��}S��=0?/�!?&q�������X>W��ӄ�<�)?�h?�GŻ�;�>��+?'��_ͽ?�a>�YA> ��>�p�>m|�=)°��:ܽ�?7Q?l���B��A�>�a���x�_}�=!~>9G/���ʼ��k>�8="���'&�(9B=�>[?�#�>ū4�o�.��𷾀 Խ�e����Y?���>9�>��u?k�$?|8��:��p���>�R=K�c�L?� �?�a9>�����F�̾��"?ƀ?$Rg>�뜾��J�M�b���ύ>�pe?~�?Vt�&I��ڑ�܂,��p?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������f�=hꬾtа?���?9$��mc>�ڬ���W�����4=�7n=�=r��pj�>��@�6�G�ƾ�N����c����>�5@�L!����>+��}�R\˿�b���о��g��?,G�>B�Q��ڸ�1=q�hV�EKW�2�L�:]A�M�>��>k!���㑾��{��;��.��z��>��݉�>��T��Q��:���J< �>�Z�>���>O�������q��?����!ο����4���WX?a^�?���?�d?�<�Hw���z�A��>�F?�Ms?x Z?��$�`T^���7��"o?�Y��6%l��A�{TU���>�I?�>�>�B��O����>�>��=S!��:ǿjM��hw�Me�?��?}3޾�E�>��?q�)?�'����ټѾ���R�M�C`:?�6h>3!�������#��ۑ���?�=?�9��9,�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?*�>Z�?a]�=Z�>0�=-����2.��l#>0g�=LE?��?��M?9M�>mq�=^�8�/��UF��CR��%���C���>��a?��L?�_b>����1��	!�Ӆͽ-1�d*��`@��,���߽�H5>N�=>Q#>{�D�c�Ҿ��?Fp�9�ؿj��:p'��54?$��>�?����t�����;_?9z�>�6�,���%���B�W��?�G�?<�?��׾�R̼�>)�>�I�>k�Խ[���e�����7>4�B?Z��D��h�o���>���?	�@�ծ?gi��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?* \Ͽ$���O�¾
� �,�=�zE=ۋ>��2�Q߼���<-8h=e�<�ͩ=[�T>�tx>%p�>�>��e>y�>d���pk"�P���/.����I�v7�����7C���!��Hi�Xs�����۾Zqa��^��kյ�=�!��B;��=�O?�6S??�l?��?�xz���
>������:�T��w=���>�q/?�cP?p ?�j�=B��r�^���}��Ƙ����g��>�;>���>iC�>�v�>�#=�uC>�El>�g}>�F)>XՋ=��<w:=�>>3��>��?���>�C<>�>;ϴ��1��f�h�w�#̽,�?8���h�J��1��X9������[h�=8b.?B|>���?пh����2H?���`)��+���>v�0?�cW?)�>��E�T��9>���L�j��`>�* �)l���)��%Q>l?�eh>w�u>�3��%8��Q�vk����w>('6?�Ƿ�VG:�c�t��I�k�ݾq)L>�ƾ>w\�����6��ϔ~���j�o�=��:?	�?���ȑ��}u�֟�?lR>
x[>#=�?�=N>Xt�����>}F��3=���=x�W>6?�c*>PO�=��>�h���wK�vC�>�(?>&3>T�??WL"?uE��C�������.��St>"1�>��>t>OwI��z�=P��>$�]>OF��������+�9�QbZ>�.���^]�A_�%e=@ޡ����=���=���]�=��{%=�~?���(䈿��e���lD?S+?[ �=&�F<��"�E ���H��G�?r�@m�?��	�ߢV�@�?�@�?��H��=}�>׫>�ξ�L��?��Ž5Ǣ�ʔ	�/)#�jS�?��?��/�Zʋ�<l��6>�^%?��Ӿ��>�2��{��iG��a�u��9!=`�>��F?����j]�'�9���?r?sT�M>��=4ɿ��w��a�>1�?�x�?�m�����?�L"�>���?�X?j>�q޾ �`��3�>��>?��R?4��>�d�5g#�Qu?i��?%�?͙q>���?��X?4�?�ӽy�C��u��N'�'<����W�b>��_=��վ��e��t��;Y����d�����|F=��!=�Z�>���dkľ�w�=W3i�E.��J}�����>���=��_>0�>�1�>�}�>*g>D"�=&
/<F�I��4��G�I?�Ց?�y���X�	I����<�4w����>��L?f�ས������>��[?��p?~>T?��>�� �{H����������g$�;�x>�%�>��>�^=��Į>n}վ2�R��>ȍ�>�ev��m��'Ž�>��>�?> ?�^A>�|(?��/?�x�=�^H>�DU��ߜ�\-K����>m'�>5y�>x��?��? *�R9��Š�����H�y���(>��?� "?���>����C	������M�=x� �*�_?X�L?K0���?әf?��?Kw3?�yD>
����}����>p�!?'���A�~=&��/��~?Vy?e��>�đ�f
ս�~޼���8��0?U#\?]-&?g���`���¾���<R�(�
Rc�a��;MzD��>�>)����w�=��>�\�=)�l�!g6��g`<1��=ھ�>`%�=�X7�0=,?��G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>'�l���K���ڙ���F��_�ŽI���= ?d��>�>?�"�>X>	A�>d���P�-����2�A}e����Y�E��.�I����!)>����Z¾#jh���>��B����>8�?הs>WX>8��>A�漅7�>�|>{Qh>��>IJ->�2>l�>��=����=JR?8�����'�Y��}����0B?pd?i+�>��h��������z?K��?s�?�?v>d|h�S(+��k?<<�>���4l
?{8:=r��k�<�X�����8 ��y��I��>�X׽�:�M��uf��j
?b1?�Ս�_�̾6P׽;�����=��?!�$?vL.�%q�1n�/�,�0^e�_l�:�)�t�����6��pt����p����B���%��h�=K�7?�ݤ?w�5��˾���,|���=��P:>ӂ	?��u>�z?_�>cJ�a1�~e�O�_�Qw��<�>[��?�h�>}#P?�X?��c?5*?�s>ww�>cY����?|�O>^�>}V+?Ǹ7?R�?Pb_?YQD?|�%?<�>r������̾��?#?��0?v?�?����(Z����>�a��M ����7�>'�)>��_��q=Aj�>v�o>`%?�9��j7�T����p>�7?��>��>�ኾض~�]��<���>�?^�>Ѯ ��Rq�1�����>�ہ?��X�	=�i*>���=����l4�
�=9�ļ���=v���)-��cj<
	�=¬�=wػ�b��˜;f_�;7��< u�>2�?���>�C�>�@��)� �b���e�=�Y><S>e>�Eپ�}���$��w�g��]y>�w�?�z�?˻f=��=���=�|���U�����E�����<�??J#?#XT?_��?|�=?Vj#?��>+�iM���^�������?Z+2?�=�>l$�Q7Ҿ�2��Ix:��_�>�|?�Zk�x<�J��$۾������=��/�$��]���,uU���-=���i~�*}�?���?݀��m4�U��n���y��t�9?��>�ʇ>��?Pz+�&<�s���p>�>��"?���>eBP?�Vz?X^[?�+Q>�8��Z��\�������2U>�.@?���??��?��w?���>��>��)���wG�����I"��`��`LM=�I[>2�>��>z�>�]�=�ǽ<����7<�Ɵ�= �c>6e�>��>{l�>�jv>		�<_�G?���>RY��;���夾Ž����<��u?���?�+?��=$���E��9��$G�>Sl�?%��?�2*?�S����=u�ּ_඾��q���>չ>q/�>�=��F=�J>�	�>E��>�0��a��n8�7AM���?;F?���=�ǿ��s��z��m����<�R����X��ҩ�m�c����=� ���z!�x���H`�n|��oS��;���s�<r�Y��>Ղ=&n�=�h�=�o�<��|��=��2=�c�<2t =!�l���@<�5,�pӀ:�M� ��9��,<�6=�C��;�|?��I?(,?6D?�xx>�?>iz;���>�t��_ ?��X>�VC�8��M�;�����f蔾�cپJ(ؾ�`�p��M>k2L�w�
>=8>`�=lS�<��=XV�=Z��=��v;`�)=7 �=	�=bɧ=���=L�>4>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��7>_'>1�R�
�1���\��b���Z��!?[C;��J̾!2�>��=g%߾ϑƾ�_.=1�6>@�b= i�-U\��ߙ=��z�r�;=@�k=OՉ>��C>Jv�=)����=��I=���=��O>90����7� ,���3=���=�b>^&>)��>]�?Z�-?h\?���>�D�����g�о	=�>F->h�>֫�<)�R>FH�>4�7?~�9?s|J?�%�>�q�=�;�>�>�@.��	o�v��,	����C=v��?V^�?H�>�>O� �,����;�3t׽R!?7�+?�q�>�.�>ʆ
�KB޿�W���a��-Y=Bl>�,�>�yZ���(��n�=*��=�ʩ���<|u<���>e�>8=t*����>Yܱ>Q�
>�|�={�>���=��@�um;�
�>+�!>���.KC<O�#�6l�=Jzx=?���/<=�Vi><(�<*®<;��=�R�>˱>o�>E��=7��	�,>`���M�)�=�����B��4d���~��.��7�Y�@>��U>L����:�?�Z>,XA>:��?��t?Ob!>����Ծ.��s�f�4�P�}B�=f�>��>��%;�	�_�M�eӾ�f�>dП>�73>�~P>vtT�kL�6���Զ�G� [�>�����tS���X��f��&�������m� �X��?/?2����>䑀?��r?�4�?d�>Ɯ��}�`'>��v������n#�� ��Y"?��#?m ?N����t��B̾���׷>�II�9�O��e�0�w^��ҷ�s��>򪾯�о&3��f�� �����B�Xr���>K�O?e�?r<b��V���SO�K���8���n?�}g?g�>�I?`B?�$���r��l�����=��n?���?�:�?t�
>�# >,p�<��?<�?�1�?�"�?�ik?af�>��>{��>��}��\�d�h>��>��>���< ?�P?���>{q�|��+����jپ-��>ah�>r�>j�=>UE�2�y=V�I=;�K>��=�S>��=���=ɀz>,�ɾ<���yE?��9>W)�>�#=?�a>�� >Z?%�"%Լv��M���B%���<�;}�⽈���w<��='k̽�T�>п��?��d=su��`�?����>��)>��>��(k�>m�>���=g�>X5�>^E�=a�>�>�FӾ�>����d!��,C�e�R���Ѿ�}z>͜���	&�П��w���BI��n���g��j�U.��T<=��ν<+H�?���+�k��)�L���E�?�[�>�6?xڌ����3�>���>�Ǎ>�J��f���Xȍ�hᾘ�??��?>c>��>��W?ȝ?ߓ1�e!3�1vZ��u��)A�!e�J�`��፿���<�
�D���_?��x?+vA?��<D6z>͢�?a�%��Џ�B,�>H/�.%;��&<=#.�>�+����`�0�Ӿ��þ=��?F>8�o?�$�?�Y?FXV�����> 3?�*?�r?�Y/?u.2?9�>�+?�6>���>�?&O8?�~-?��>�� >ѥ3>��<*�/=yƋ�v��9���;HԽu=�"=���<t�:v��<=h=�(=��;[O��>�=���㒺��I=%u�=���=�ߦ>��Z?��>sh�>}q;?�Y�$�4�c��Ħ/?�p=�y��8ω��������>S�f?«?B)\?�[_>��>�qK>���>	m�>j� >k�\>�{�>'��D�8���=̂>�N>6 �=��U�p���6q��&�����<� >�d?���>&����w>�XҾ@�����=[�u���ھ�i��Z�<�NJ������$�>�<?9�?��%<]	��#�e���'?�jD?�gh?K�?�P=�����{J�2�?���+�P�!>@<`��²����G]/�"R,<�q�>�TԾ2���
�t>V��֭��4o��8=��f�"�=X���|U��S�	t޾䯃���V=�Y>U�ž�1#�Ȱ��\&���F?IQ�=⋥�=W�74���P>�>�f�>��m�pz˽o�<�!����5=/��>�u>u�[��wϾ$C:�+��wB�>QE?�H_?�i�?����r���B������`����ɼ��?�e�>Uc?��A>���=\������d�nG���>f��>$��J�G�.��/����$����>�0?�>��?ʻR?G�
?c�`?O*?�A?�5�>_ŷ����=&?(�?q��= ӽ��T�6�8���E�_�>�v)?�C��M�>S-?��?8�&?�xQ?�?��>� �;U@��h�>�4�>�W��\���`>��J?���>2fY?�Ń?'�=>Ά5�����ʩ�('�=�>�2?�9#?r�?�8�>���>�e¾�� =egl> �Y?ob?rIf?&�2>�O?�s�>E�>EX��ښ>x��>�U?�Y?�k?�C?���>���w��/���3~�
��;��0�Sd+���H9ڻ\�����;���=R� =�.�<� ��I�k�k~�e\�[�*<+W�>��s>u���0>y�ľY��i�@>����'��ڵ��ү:���=`��>�?��>4
#���=��>[C�>��q+(?�?��?q�;�b���ھ��K�s�>�B?�Y�=��l�)v����u���h=.�m?Յ^?`W�3��0�b??�]?����!9��pƾ�]��꾪yM?�	?/Q����>_|?,�o?GX�>�We�#�m�	Ȝ��{c��un����=��>���>�c��6�>(�8?ș�>�h>��=�zݾ�mv��N��^�?�Ћ?�-�?�V�? 2>�ul��A�^y����Wb?%�>ik^���*?��B�J������=R`��wξʏ�K����@w�[���aO�&d��h�F�bp�<�4?vz?��u?/t?��ӾUh���g�8�t��qX�D��}	��&Q���3�yUB�e�u��|0�<�+��Mܾ�@���L�F��~�?��?>2��3J?�꠾M��$��g4>9^��eq4��#,>�ڡ����;�<�o���E��]5þ��;?CЕ>���>��>?��E�i�5�444�9&�F1�ގ�=?��>(o�>%�>����؃�x6����-��/!�ڰ�>��Z?YF?>�w?��y�p��R<t���%���������1>�>#_><,���H�T�'��9I��������Sj�2x�	��<�d-?���>N�> ǈ?��	?���b�۾)�����]�����@%�>e�t?��>Wi�>+_�~@L�2?�>��g?�h�>�
�>�F���
&�����R�½��>;�>X@�>QS�>��g�}_��|���S���@�<�=
Gy?�f����k�8x>fR?k�<u�=wR�>(uؽ�#�?H��ҽ-�=�g?�yn=�P�>�0ƾK��KHr�Pꕾf��>��>���x�Z��b6��K�>�-?��"?gg�?�� ?e�������>g@k?Fc?�b?��	?f�>hҫ����ǜ�Ko�r>���=���<[=�����AǾ���6U�=���=)����h�I}ɻ�֟��"�;}*���cH>+�ۿ�CN�QG;�p���Ҿ}�����~��"�
���z��J��]��h=s�����~��J��y\��+����k����?�k�?�i`�ͷB�����r�~�ë
����>�!��U<�6����˽DI��1E۾颼�ʱ0��_�5t�$�e�n�'?G����ǿᰡ��:ܾ�  ?{A ?�y?��V�"��8�_� >6�< 3��V�뾷�����ο@���6�^?a��>��o0��d��>��>�X>�Hq>����螾*�<��?�-?y��>��r��ɿY������<���?�@i}A?g�(���쾼+V=[��>ӑ	?�?>I1�F�����R�>X7�?���?�&M=��W�m�	��{e?�� <=�F�[2໘�=�L�=C=O��2�J>B[�>�|��NA��ܽ5�4>�߅>.,"�={��t^�S�<<�]>��ս�!���?\�[�ݰd�c�0�4z����>کT?Mi�>"�=q�-?��H�0�ο��Z��,b?5a�?M`�?�=)?�㺾�1�>n۾O�L?��5?ĕ>��(�Q�t�f��=�BӼ��P�ɨྺsV��g�=A��>$5#>�O'��2�),K�a�f�e��=���"�ɿ:����*��>q�=٣[�۽A���ͽ�S��|釾g���L��E��=&�	>�|>RJ�>�b>�GP>�F_?6�s?�>p��>]�˽{і���Ѿg}�+e����q����p]�������l�� ��a8�s�+� +˾R=�KD�=�8R�j����� �O�b�<�F���.?�w$>.�ʾ�M�Ǧ*<zoʾ^Ҫ���������2̾O�1��!n�rǟ?��A?��e�V�.��t>�B{���W?UZ�\���ꬾ�1�=ű���=�E�>m��=��F3��S��1?n=1?~�;�1��WB>���=k�!?���>�*��T�>�?�}^�3j���\�>g;>e�>B�>�%�;P��ҭ��o"?�}"?0~�)���$�>�����C�]^<>Y�W>�=E`
>�K?��c=��"���=J�=IA>�a?dҧ>ƭ<���E��Ti[������hf?0?�,>�k?�5]?U�e����Pz���#�&��6�:?�/�?�@>���u/��N���u8?��m?׏O>/���Cl��/G��d��.?�s?�?��&=@��u䋿���G-?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������ɇ�=�B��Ư?��?B롾Fs�<3��n���U=���=�P�<�ȯ�'��G�6���ƾ%�l˯�T��v��>�@A��w��>N������̿���,�ξ�F���?Ҧ�>��N�EOȾ0�p����)V��=��-��x6�>	9>Ċ������z��M:�A����>�o��+:�>�h^�5���eO���ߜ<��>��>��>�ᖽ������?����gCͿ��cT
���V?��?d[�?�?`��<��y��y|��aC�QyE?}hr?�+Y?�.�AYY�d�4�i�j?3�(w`�J>4��ME���T>3�2?���>M`-�ۀw=��>���>��>TM/��Ŀ�涿"e���ɦ?���?��꾋��>�o�?�|+?���<陿�驾�+�|���>A?!�3>.���U!��=��͑��
?�N0?%^�'s���_?��a�9�p���-���ƽ١>ظ0�DZ\�������TXe����<y�r��?a]�?M�?7��V�"�?5%?��>����8Ǿ�
�<T~�>�&�>N>Uq_�ѧu>����:��f	>���?i}�?5i?s�������U>��}?Ii�>�@�?���<Z��>F&;���mя�>�=[��=#���.�?cGX?�i�>������a�\V5�ibM��e�S�ݾ�*I��*q>kkS?�F?0�>%_� X�=ݳ�{����@8�2�Z��mM�Y�3�Y��T>gŗ>�F;>򐍾����?Lp�9�ؿ j��"p'��54?,��>�?����t�8���;_?Lz�>�6� ,���%���B�_��?�G�?=�?��׾�R̼�>=�>�I�>@�Խ����]�����7>1�B?]��D��u�o�|�>���?	�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*lhֿ����N��T���,��=7��=��2>��ٽ�^�=��7=a�8�Q=�����=��>��d>Mq>L(O>�a;>ԓ)>���D�!��q��O���o�C�������Z�6��]Wv�^z��3������#?��4ý�x���Q��1&��>`�,S�=+�V?��K?�Ej?���>
�W��( >8���Ɂ�<R-0��Y�=?-�>%/4?�I?��)?�Ɩ=���
�c�N���ǭ�{Ä��0�>�?>(}�>M|�> ޭ>�{���	E>m�I>��>Qm#>�x=��I=�� =k0N>褬>�M�>���>wG<>�>ϴ�^0��@�h�fw�̽` �?䀝�h�J�s1��s;��ۦ��dZ�=�a.?x>����>пp����1H?�����(��+�$�>4�0?	cW?��>P��-�T��9>�����j�5_>f$ ��{l�ދ)��'Q>j?,oj>[7y>�3�K�6���O�������z>�5?���$@��\t���H�4#ܾ��D>��>�eL�R��ޖ�����l��a|=�:??����2���xn��z��ۊQ>n�_>[�$=�&�=�	Q>�>�޹ý�@�M�I=�u�=L?`>�B?.�>I�=�>g��01[����>J�G>�j7>�'B?q�?pJ��Ӆ���i������>�#�>݈>,�
>��E�3��=G8�>^R>^C���9���	���9�[X>_�V�^k�,���_|=�Z�,�>	�=�U��.�XN=�~?���(䈿��e���lD?S+?` �=/�F<��"�E ���H��G�?r�@m�?��	�ߢV�@�?�@�?��L��=}�>׫>�ξ�L��?��Ž5Ǣ�Ȕ	�0)#�iS�?��?��/�Zʋ�=l��6>�^%?��Ӿԕ�>
��fk���憿��u�=��>��G?�o����[���B��:?.?'�� ���ȿWyv�<��>hD�?{��?z�m����r�?�E��>��?��X?�1g>C+۾��]�s��>��@?T>R?�t�>�g�_�)��$?�1�?k�?QI>A��?��s?�m�>�Jx�Z/�6�������s=�Y;�c�> Z>����hF��ד�Mh����j����)�a>�$=��>�G�A1��gA�=e⋽�F���f�Ĥ�>H$q>��I>	P�>�� ?c_�>6��>��=�f�����#���p�K?r��?E��m�H�<�'�=0 ]���?�j3?�����j;�y�>2�\?��?��Z?�ԓ>���e����~��S��ɽ�<��M>W��>=V�>����)aM>=lԾ0#C����>�>�X���־HOx�$<o����>��!?���>&X�=�u)?�.?�
x=�̸>�>E����� h�W
�>b��>AM�>�Y?O�?�i3��D�
���u���uae��f>�Ɍ?��;?�5�>�#��=/���Ͻ�<�0��s?���?F��#p�=��?� ?�?Vz����k@�Z��<��>�<"?(���'B�c�#��}��A	?��?���>��������s��ԩ�)���?��[?;D$?b	�SKa��zƾ=[�<'���9�2���9���,>�>ko���=��>�F�=�l��#2�ݘo<���=���>��=M~0�����=,?D�G�eۃ�E�=��r�!xD�,�>�JL>�����^?�l=��{�����x��VU��?��?Wk�?o��0�h��$=?��?Q	?�"�>�J��J~޾��ྌQw�1~x�gw�W�>���>��l���A���ř���F����Ž���<�$?��$>��?"�>�m�>��p>tX�y���'���v _�p��
W���D��A鐾3��]����Ѿ!�7��ۖ>��X����>�;�>��>e��> ^�>1Vp=��>��F>���>�u�>��|>B��>62�>�.�=����KR?������'�������!3B?�qd?m1�>ei������ �?���?>s�?�=v>�~h��,+��n?d>�>=��0q
?T:=�E��0�<�U����P2��?�=��>�E׽� :�mM��mf�{j
?�/?��O�̾)<׽_x��=g��W�?��??�Y��j��mq�`5O��Vz�F�����<Vu�'>��=n�S8��-X��}���b����;��L?�K�?)TQ�ƾ���ZI���j�x��>�#?�O8>X�>��<�7U�N�F�qˁ�j�S�����6?y��?.k>I�J?��C?�=Q?.I?���=D?�'�o�>��1=�L?׍?�W?H�A?a�"??+(?xLK?���>��<�)�^�־/�!?�?+?ͥ>��?�̋��@�<R�>���ʾQ	�g�[>M=�=�A�=U�z==�9>#-@=�W?��M�8� ����j>�}7?^��>���>���&�����<��>��
?�J�>����yr��_��W�>���?�����=q�)>9��=����ɓպ�Y�=������=y ����;��B<��=1�=�Ds������:��;E^�< u�>6�?���>�C�>�@��/� �c��f�=�Y><S>{>�Eپ�}���$��v�g��]y>�w�?�z�?λf=��=��=}���U�����H������<�??J#?)XT?`��?{�=?_j#?ҵ>+�jM���^�������?u4,?�>�w�ʾ�ਿ��3��W?6L?va�Uk�{R)��¾^4ֽ% >/��K~�B��sD��f;�������?ǽ�?wA�0p6�vK辷��������zC?Br�>3��>ف�>Z�)���g��!� �:>Od�>4�Q?S$�>'�O?:{?U�[?bT>��8�10��ә��23���!>r@?J��?�?y?Zr�>g�>B�)�;��R��e�� �����W=�Z>.��>�)�>��>	��=�Ƚ
g��8?��R�=�b>��>ˡ�>/�>&�w>h�<BD7?��>Z���+�G췾�}h��(�=��?�?OT<?����+��2������c�>���?��?1,@?��]��=���\̾���8�6>�ȥ>&z�>��=�n=
	V>���>�P�>��&�Jl���$��c�<
M?B�*?�ͧ=|Ŀ��h�JMB��I���}=���p�7����}�)�~=t+����қ��TG��U��Ì���y��<����^����?x�j=�D>,��=�Y�:���v3o��=deڻ��C=UFj��0=M_��_(k8�a���J���=,��=#U���˾<v}?�KI?��+?��C?��y>��>��6�+�>$��G?%*V>sPO�R��S�;�����1��
�ؾ4�׾Lc��(�>0�H��J>W73>���=u��<�*�=h�s=P��=�1�G�=NF�=T�=TO�=���=�>�:>�6w?X�������4Q��Z罤�:?�8�>h{�=��ƾq@?|�>>�2������xb��-?���?�T�?>�??ti��d�>M���㎽�q�=U����=2>r��=v�2�T��>��J>���K��B����4�?��@��??�ዿϢϿ5a/>�:H>3h>��S��*�F�Y�WD�Lw[�?�?��7���ؾ=��>Y�=��ھ%�оlT=�I,>{_=��,���_��o=ȏh�-W=�=��>�<>�V�={���#�=��x=X��=��S>��&<�Ӽ�<�,��=	>Gqi>�%>U8�>.?`�:?]�T?��>�tT��6o���R�z*�>U/>MN>7�Y�0�_>���>A�??�3H?�@N?��>��<�c�>�1�>�0-��u��Hi�Ӳ���ݫ=Ef�?�͎?w��>�4 �~퀾�?�_�7��1��L ?�?��?��>)'�u�濇~(��.j���{>>a=O=����ؽ�B	>b!��	�L�g��==�>�7�>̶>�1�>Lu\>y��=��>	>D�=5��=�.c=/E>}8>dU=Qo��>�M�S��=
Լ�m����J����<G>�`U�P��!��=���=^��>�8>a��>�=����A/>����Y�L����=uH��,B�x4d��I~�/�*X6��B>�7X>~~���3��k�?3�Y>2l?>j��?�Au?�>����վ�Q���Be��WS��͸=ܵ>��<�Zz;��Y`���M��}Ҿ&e?H#�>����>K48�ΐ �5gd�p�޾�
���=�u�bR>�Q�sۀ�����M�����S(��dbo?�H���4�=��e?��F?
�K?o ?a�=�a�ft�<�w�l��>���S�=����H?��$?���>���c�f$̾ݜ���·>�H���O�Ε�/�0�l(��з�Ά�>F�����оo@3�%h������B� �r�3�>��O?4�?y�a��c���ZO�����V��TR?}�g?Iv�>�1??��b��t���w�=��n? ��?�3�?��>���=M戽�B�>��?Ic�?D��?Dz?�v����>[*1=Fa�=�� �3 >/�<>��=��>��?'�?���>�G���	�]%����� ӄ��OD=�9�=�5�>��>$n�>��=�Ab<��b=?lB>�Ğ>v��>��K>�Z�>⊌>t�о�'
��~:?hw> �>�7?cf>A�xÂ�6g�<�X���ޥ�~6D�8�м��սԭ�����\�=�������>��ο��?�'�=��'��?{�Ծ�B�=x�=�w�>��E��
�>�l>�#>ܯ�>3͓>ؐ+>L��>� !>�5Ӿ>�>����c!�t.C�{�R�%�Ѿ4z>A���S&����n2��vI�=v��~q��j��-���8=��Q�<�F�?8�����k�$�)�����L�?�X�>6?�ӌ��^��;�>���>9ʍ>�D��󍕿�Ǎ�|c�j�?��?BBc>��>��W?��?3�1�83�8uZ�v�u�x&A��	e���`�]፿i����
������_?�x?.tA?���<�:z>|��?�%�lԏ�!-�>r/�y%;��q<=�'�>v-��C�`�8�Ӿ�þ�6�1WF>��o?�%�?�Y?]cV�
m�C�>&r6?C�*?8�r?U.?X�:?���D�#?��C>��?�?�3?��.?��?9!E>���=�?;� 3=*��EH��o�˽� ѽ"7�*
=�7c=�k?���d<�=�D�<�Q��Q6���q�<�y�����<��1=�L�=���=<��>$q]?B��>v"�>��7?"���7�:��E�/?F�?=����4⋾ON��U��L>��j?��?b�Z?��c>�B��zC�c�>2ۈ>��#>��[>뀱>�n�h�C�=�=�>Zy>���=�'P��z���r	��a��\��<=9>l��>�vk>%ꌽ�>�]���cs���n>Ɍ@� n���+<�KuG���4���o����>eM?b??%��=#C߾RG���6e�
@$?��7?�L?R��?"%�=V��YN>���L��J$����>��<�b�+���:$��le:�B�s;kkm>6☾�]���yl>$N������p��]>�>��*�=Ld�o�;���;�Wv�	��=��>����;��QL���ا�b�G?���=jA���]�_𡾨lL>l}�>K��>(�����ǽ�B�ެ�~��=�>�>{%L>Y��<�;��L�����>0�C?��X?$?����Xat���A�!��f���z�ƭ?ys�>��?,�3>n��=���W�Cc�ظB���>6:�>����oC����=����$�iC�>��?�'>3d
?��J?t
?>._?��+?��?���>��5¾��x&?Sh�?f�=��нF*V�s�7��CF���>�c(?��E��
�>b"?e?�+&?�HQ?VH?}n>�����@�U��>Mv�>AW��'��D@c>>�J?�U�>1Y?(H�?��:>I�5������ƪ����=%�>��2?��#?��?O��>�u�>�&l����>��>�Ɓ?%�?'��?9꼁y=?�+�>K`1>����'�>�i�>�?��l?yC�?�FI?�k*>*��[�k>l���$�Y7 =ai=_w�=y63�p̎8���<�S^�S֚<-!�<��ս0v�ld�M��&��<9�<�a�>��s>T���1>�ľY����@>����MN����K:��+�=h}�>�?���>�t#�Â�=���>�N�>����/(?�?�?.�(;O�b�0�ھ��K���>wB?0�=��l��}����u�F5i=�m?�^?��W��=���_?��M?g��9������M��`�'F?e��>\���v�>#n_?�N?L�>�>�ta�(���GP��䀾gf2>%�>ۨ���Q�C��>��\?�Y>��>v�Q��j����r���Ѿ�8?q?���?�І?�҉>�v��޹߿�����ԕ���e?�w�>*����'?������;���\�d����Y���ī������������#t��6ᶽQ��=�"?ŝw?e~p?�g?�Z��yh���d�uz���a��g�G)��g+��|R�+�T��t�Q��+���������<�*����J�W%�?�?Vq����>.����D߾%�ɾ�F`>/����7��ޣ=8̼m��=,�=�k����!g����#?���>���>��=?N�V�*�4���3��v*��x��>	�>���>z�>Á��FE\�^S߽48��'���6�>I�`?A�A?�Wp?l,��>4����d:�c�=�+	��Fy>�O/>{|>udm�˽1�)�	=���j����B��x��%=`5.?^��>�B�>#b�?��>����/��cR��)�v�J<�Ķ>W�q?�*�>�P�>�>�D�)��?�S?8>�y�>|1⾹��v��8���~�{>"$��d�>�
�>�ɛ�M"[�a��椑��RY��Y�=Kq�?BMO��?�-َ>`�`?a�6�B:��>���=����
i>�W��F�?�>(�>>�d�Yh�V/9��G����&?`�
?{���Mz(��#�>'j#?��>�^�>�ކ?�O�>]�Ⱦ&m���?t�[?V�H?��C?t��>�ID=�𽽎YƽM[1��F�<	�~>�R>�t=�'�=�&�rlb�S��.�B=ϳ�=?���+�ʽ����`@����J<IU�<��:>�kۿqQK��?پH���$��/
�h׈�������y�@p��lg��'�w�.u�8=%��cV�$lc��K���)l�j�?�>�?%o��B@���o���T�������'�>�?r�7s����i<�	���9�ྃ�[<!�9P�-fi���e�~�'?j�����ǿ�����(ܾ� ?o) ?k�y?V�G�"��8�9� >�K�<d���[�뾛���J�ο3���3�^?���>���%��%�>��>�X>t#q>�쇾(ힾ��<�?z-?ϵ�>ir���ɿ�����<)��?��@�fB?d$�R�ﾏ�=%d�>4H?�p7>`�6�����9�>�͝?���?uW
=��S����F�d?����QI������6�=Le�=�K=/����D>]L�>���9�^&ѽ�a5>���>%U(��	��Y��v�<unj>�@���:��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=u6��{���&V�}��=[��>c�>,������O��I��U��=V�y5˿��)�I)��>�����]}<��+�;ἐ�=D��a��|C��ip�>�B>���=5�3>p�>'g�>�mN?��o? �?%��>%(�=�R��d���e�����m�P>��N�3̷��s�/Ӿwt�������@<ʾC�<�`T�=�JR�a=��y� �X%b�]�F�{/?��">˾�8M���(<B$ʾ�誾]̀�(a��3̾a92�Y0n�c��?7�A?�Ņ���V��J�=����ٹ���W?I�������]��=k����=�L�>��=�hᾍ=3�*�S�8?�B$?�%ξ����!�>;�;��ʼ=��R?~G�>[�,����>H�?&���+��l�>�@P>��>_�>9Vi����� �r���%?E�9?�`�<ٽ�)s�>�����c>D�`>�s]�\�`>�s?�!�=?F}��?�K��>�>��V?D�>so*��t�L#����/�:�=t�t?sE?h�>*�h?f	D?P
<����m�U�Vo�?�O=��U? j?[w>�>���о�h��ls5?7Re?��I>��c�ԯ��/���A%?v�o?�B?�%�:�z���m���6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������e��=Ű�):�?G�c?����+󃺓��^C��4��Z�=���;%$��߳�����Z$�s���u�9_���d���X�>K^@R.�CL?Rj]��6���ʿ���Uv�T��0<?'��>��xR��&�}��䐿��t�<�>�f�7���>O�>Rє�:֑���{��M;��Q��7��>�3�%��>��S��9���p���t9<5�>c��>���>�E���꽾ộ?�a���*ο
������s�X?#I�?�y�?�s?�2><��v���{����G?��s?bZ?D�#��v]�Ĭ9�N�j?|K��	2`��3��E���S>Ž1?��>ID-��8q=��>���>-�>A8/���Ŀ�Ѷ�����䗦?N��?���Q�>Zf�?�,?�����sA����)�j9)���??�5>l ��x� ��t<�q����q
?m�0?l��|�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\� N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>hH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?���>�ʄ?���=	�>^��=fb����^�}!">��=:U[��?&�M?N0�>^��=^�<�p�/�a*F�t0Q��l��,C�<�>�8`?��K?��d>����{3�h� ���ɽ��,��p���=�r�-�p�ܽ~�>>��>>�>�=G��|־��?;p�3�ؿ�i��1p'��54?���>�?����t����;_?,z�>�6�,���%���B�V��?�G�?8�?��׾�Q̼A>��>�I�>N�Խ���Y���~�7>3�B?���D��`�o�|�>���?�@�ծ?Ui��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*~QԿ}���]�	�}�*�M!��W�>��
�#��=�O���Tu�:��>�>[2l>�l>��C>qΉ>r�y>�����5w�����6�r���+���Ͼ^�8��|��#W���$#�y*��Ee�=�A=�_�D�ž���g׼�K�=o�U?TR?�p?� ?��w�*�>����/Q=��#�z��=p]�>]p2?I�L?�*?។=�W��g�d�\���H��ʹ�����>c\I>!��>��>�/�>����I>e�?>�^�>n� >��(=�p����=�WO>\D�>h��>���>χ=>S3><����ΰ���h�; u�~�ν�
�?;P����J�*╿�#��b����=uI.?�
>�ߑ�xoпV���#H?�|��b��#W,�;e	>N�0?"W?�r>����{�\��<>Χ���j�ڥ�=>�����j���(���O>�?<Mg>�fu>[�3�� 8�e�P�=쯾��{>�d6?h8���D:��u���H��[ݾi_L>V��>d�@��3����>$�5[i��|=f:?�s?�����۰�CYt����jR>0U\>M�=c��=|7M>A?a�~Nƽ��G�1=Z��=��^>�N?l
->#�=D5�>�����R�e��>,�@>�|+>��>?�%?D��KR��q僾��-��t>�>�>�>�E>�I��V�=���>�b>��������T�Q	?��7W>Ǫq��s^�1b}���~=PY��]�=�4�=ł �t�?�o�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�|�>h��W��C����u�؆"=�M�>
H?�/���zP��V>�T�
?��??��ն��\�ȿ]�v���>{�?��?��m��4��)�?��o�>`��?�?Y?��i>�j۾ְZ�\9�>��@?[R?�%�>�E�KT'�I�?4ɶ?ޫ�?#�e>�o�?�vQ?���>ю½�7����������v=�܈����>�i>�Ѿ�H��ɒ�Lሿ��j��C���>��`=��>�;#��|���*�=��������+�:�>]y>�f%>���>?�r�>:�>:f=�晽�|�� ���L?F��?��l�m�� �<�0�=_�Rq?7�3?�v��zϾ�ި>4q\?~|�?��Z?Yb�>`���\���迿�V��c�<�K>�
�>�`�>�7����L>?~Ծ��C��]�>~��>�����,ھ��4W��)b�>@�!?m��>Gʮ=��?��5?���=��E>Ʌ3�	,��� R��=l*�>ѯ?��u?�--?S�/�O��
��ꙩ�� q���O>��~?�~?�8�>�ޒ�#���?��=U+�=�蔽�CI?�W?�����a>h<�?�o=?�,?�k�������߾��0����>�"?���.B���#���(
?�f?[R�>ﯩ�i�:6��~n�����?w,[?U�$?����d�WǾ	��<���1̺Ӄ�;/t�I >�>:�z��_�=`3>/7�=��f���7�82�;��=걔>
��=�4����0=,?��G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>�l���K���ڙ���F��_�Ž�����>1��>b&?r ?bP>B�>%����4'����t����^��b��z8�7�.�̋�����n�#�_]��!¾O�{��<�>�
����>�
?��h>_�{>��>��»�R�>%R>�n>틧>�"X>�55>�>��%<�xн�KR?v���(�'������S3B?�qd?t1�>�i�A������y�?���?(s�?�<v>�~h��,+�)n?t>�>&��Hq
?�T:=�7�?�<�U����>2���ɪ�>�D׽� :�~M�hnf��j
?�/?��ɋ̾�=׽�ۋ�J2�=��?h?k`-��:p��x���K�R���p=r���,v���I���|�	Y��������������N=��(?�i�?m�&��ξ1錾P�u�T<.�9?�=c�?za>��>�S�>`(�$+���g�N�Z�ʹ��?f�?:��>��F?�vK?�V?�@4?�m�>���>G��<D�>W*�;�l�>W��>*oJ?Z�,?��6?�JH?�J?�F�>e����2徼:��tC,?˯>�
?�J�>�B�>����<԰=�j�>	B��/Ҿ:J�s)�=�V�=|�>I��=�c3=�p_>�H?,��9�[r���jk>2?3R�>�Ͼ>Ci���)���&�;�"�>�?��>�n��~s��:����>���?pnּ��<'(>_��=	w�ߝ�:e²=�?��i�~=�?ؼ?8I�k�;H(�=��=�H��&b�:��:�E<�k=u�>9�?���>�C�>�@��� �Q��@g�=DY>�S>�>�Eپ�}���$��U�g��]y>�w�?�z�?O�f=��=&��=�|��nU�����]������<ѣ?AJ#?+XT?Z��?p�=?hj#?��>�*�`M���^��J��Ȯ?�',?ߕ�>�����ʾ@騿ۄ3��m?\L?D-a���0D)��J¾؁սBL>�/�,7~����iD�54[�B��������?ŝ?;�C�Ӯ6��h�|����O���dC?JK�>��><A�>Ϩ)���g���k^;>,�>nR?)�>a�O?��z?�[?bsS>��8������Pu2��� >�V@??��??Ǝ?�x?�"�>��>�*���:���/���@�R$����W=�Y>���>��>aة>
�=�Ž������?�#��=��b>���>���>`��>pv>է<��G?-��>J���m��|���U��Ey;��u?��?�j+?�\=s���E�4P��iJ�>[f�?���?*?|8T�U��=�9ؼ�ⶾ��q�X�>�>R~�>0�=!�F=N�>	�>���>T��G7�2a8�h�L���?0'F?W|�=?DƿCXo���O�48��%�=W���I�]���
�<Tr�e��=J��-�/��𖾼f(������֖��#�����j��� ?���=5�#>.q�=a=y]k<9��<zrl=:מ<��<:���<N:=B��n���{��od�<1t^�r�G�|�&��}˾T�}?32I?�+?^�C?,�y>�)>N�3����>�����I?�5V>��P�������;�򴨾N%���ؾ�l׾��c��ȟ�])>�;I��>23>35�=�>�<?!�=��s=�͎=��V�--=T8�=A��=�q�=C��=�>31>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��>	�c>OlV���U���w=�~��dL?][��J!��uq>��>5�Ͼ� �Y��=�p9>���=���#nz�LG�=2Y���=r�{=���>�9>���> �<hV�=�=a;�Q�=iB><ٖ�΅����G� >?�>R��>�f�=�i�>:�?�0?�Md?���>��m��;ξ�g��>��=�	�>	��=�FC>ָ�>�	8?�D?�L?N��> ��=���>紦>�S,�7�m��|�����<q�? Ն?P�>�,@<��B��{�<A>�VŽ��?J[1?/?�
�>C��R��::��R�S��1�콁_%>�LL�'.>��Pe=]H�x:��E�Y>��>*��><��>�7>gc�>���>�ͬ>(^�=�"-=���=��9=z�/;��ս<��=Dj�;3��<X6󼘁���ul��" ����<�ӵ�ע���H=��-<H��=#��>H<>��>Ύ�=����C/>ʸ���L���=�G��R,B��4d��I~�I/��V6�W�B>�:X>�}��74����?B�Y>�l?>���?PAu?A�>| ���վ�Q���Ce�VS�@˸=�>N�<��z;��Z`�|�M�}|Ҿ���>�%�>7��>�Bw>�/�bH=�޸.=Yܾ/�3�S@�>G���g�ἦ\�\bp����WП��Hi�rba9��G?�,��,�=��|?z�J?bK�?n�>$-W�oSվƩ.>J����qr=Y��Jh� z���� ?D&&?��>c.�/�G�%E̾����۷>�@I���O�9�;�0�6���̷�c��>������о�$3��g��������B��Rr���>��O?��?::b��V��@RO�%���$���p?+}g?�>�H?kA?|1���u��p���z�=��n?��?~<�?�>���=���)L�>v�?�8�?��?
�w?��<�	?��y=���=hK��>�>mA�=��'>��?��?Q^�>/ǚ�D)��� ��~��^e\�5="۶=�x>:=�>�'y>,�=47h=1�=�"&>ǻ�>Ð>I�V>�T�>@2�>m���i(?Vvؽ5h�>/G?>t`>��>��>xzI>L��)�ʾ�q����=��=���=���ƒ;���E�?U���S>�?T=N�/����?Y�%��&�>L>=<�>v��7l�>Oŝ;8B@=R�>���>:,R>�ڮ>YN�=�Ӿ�>���c!��C�ӉR���Ѿ5�y>�����%�]���N��)�I���������j�u3��5)=����<f@�?e���>�k�*�)������?�;�><6?:Ȍ�蟉��o>A��>vٍ>���m�������}h��?���?�;c>��>I�W?�?ْ1�23�vZ�,�u�n(A�-e�V�`��፿�����
����.�_?�x?1yA?�R�<-:z>R��?��%�[ӏ��)�>�/�'';� @<=u+�>*��0�`���Ӿ��þ�7��HF>��o?<%�?wY?ATV��DX��+>�6@?�z0?j	w?ˁ2?�>?=��L�%?6�G>�?Q�?r�4?��/?GY?2I>M>yM<N��<[y��@����H�aн��B�Lh==��=E��;X�Z=m?J=�s;� *�L������k.��o�<��%=`�=���= �>2�\?���>�P�>��8?���
6����1?i�M=�I��.���p���;�U�>�hk?��?r(Z?v`>;�A�	2E�*M>��>�%>��[>���>	����A���=�>��>E:�=�[��0�����_��j�<��!>p��>�0|>�����'>�|���.z���d>��Q�[ͺ���S�-�G���1���v��X�>�K?p�?���=�`龸0���Hf�%0)?�]<?hNM?�?q�=7�۾'�9���J�@���>a`�<�������#��I�:��b�:��s>�2��-��&M�>����F��䈿��7�GE��*�G�����%��M�D�!���������,:< �쾩m�m�������?:?ᴺ<^㾉ξh̔��n�>AH�>��>˞ֺS`s�$�F��߾��<��>���>��Һ�j���J_�{)�
�>s�D?�m`?�t�?��{���p��TB��� �͵��ZԼ4m?��>��?��B>{�=|ΰ�M��s�e�O�G��0�>o)�>]T�'�F�}���>�C%��(�>�?l}">H?8Q?��
?u�a?Z�(?��?�(�>����kߵ�r�&?���?sXp=r�˽L�R�C5��"E����>.E(?\zS��F�>�~?�?��#?��O?�?�>q���NB��q�>�d�>
�U��ů�F�p>֮I?�m�>�1[?�z�?'Y9>��3�	r�� ��=��#>J5?��#?�I?�V�>ϒ�>��ž�W"<)�ý�[(?q��?'��?�'�>3~!?��>��>/�>�?H��>�+?uQ?hy?�W,?���>��=Sc��d���q�Yk�=�r����=�W�=����xZ�������=k��=`n=o"|�1�ܽ�
��"�=!d�=
��>��t>���1a3>X5ƾ���A�>>�1�� Μ�^��n+7�/�=��>Y�?i�>�P$��=X
�>x]�>���b(?�"?��??��;^gb�)�ھS�O����>�A?���=m�l�`"���v�ufc=�n?f _?��Y����d�b?(�]?�h�=���þ.�b�"����O?�
?�G���>��~?��q?���>��e�1:n�w���Eb�	�j�%Ҷ=Nq�>�X���d��A�>��7?dN�>��b>k'�=�v۾v�w��q���?d�?�?���?�.*>��n�(3࿖ ���?��"�t?�1�>ج6�5!?�Xd;����&�׾p�7�����y���u��`�nݒ��)���tj�}X>=ɬ%?y�v?$�x?/h?���fd��{A��2]�X���������1�>b�uX�e�u�v�7���$��z־�ʽ�}��[0����?9�=?�@��x��>�3�����
p��8>@���+<"��ˬ=Һ#�?�=~{&=Y����p��O'ƾc�)?\k�>n��>��??N�F���$���6��9�b��Zi
>�q�>b��>���>��6=��A�V)���\F���$��n�>�~g?�\B?䔅?_�O��==��΁��U>��諒C)��z;Y>�e�=6yy>@��i�y�y�'�o96�հs���j���	v����.=�!?xO>���>���?G�>"����C徭����E�M*��L�>+^?���>[̍>]T6��D��R�>��p?N�d>�&>Ԫ��N��v'������cծ>�s>ރ>�h�>#k侺~t�ʜ��.��Q�m��>��v?�EV�ؒ���}�>=1?0V!�X�=��>�(���xW�^Ӳ�)H�=Z�n�x?��=�2�>��"��@�r�����?���>��g�D57��[>�v!?y�$?G�>�?5�>,�־-$ڽ/b?�;P?��??�o:?U_	?��=�!l���_�� ��il�&]>���=T<o��=+ܚ�&;E��N���K>bm�>���;%C�u<.=3W���<Ԧ��D>��ڿ.K�N׾*1�����	�`�������=��(��g���������p����)��wP���a��Ҍ�Qk����?��?龈��|�*5��n�|�3��䣺>-wt�i���X���f�d��T߾�O�"�r�S��Pl��Cg�7�'?�����ǿⰡ�=Aܾ� ?�2 ?ǔy?����"��8�� >���<`���ײ�Н��/�ο������^?|��>B���t��>H��>w�X>Tpq>/��	����<�?�v-?���>�xr���ɿ����M�<���?�@�{A?��(�����U=���>Z�	?��?>1��>�����E�>�7�?V��?eM=��W��x	�]}e?2�<<�F�Jk޻
!�=n%�=i=߿�zJ>�h�>�_�sAA��+ܽ��4>�؅>rh"���a^�^q�<'�]>�Vս����3Մ?+{\��f���/��T��
U>��T?�*�>|:�=��,?\7H�b}Ͽ�\��*a?�0�?���?'�(?5ۿ��ؚ>��ܾ��M?\D6?���>�d&��t�υ�=56�;���w���&V����=Y��>a�>��,�ߋ���O�sJ��Q��=6l�������!�!�cug=;؝��:��(�|��{��2g��/�g��d�o�}=2��=��>�.�>�Du>c�]>��S?�T}?�^?�љ>eɽ�2������0Z;�4�����ē�ex�@e��$��`���kJ5��'3�TYؾ�=�I1�=�6R������ ��b�}�F�{�.?�p$>b�ʾ��M��m+< pʾOȪ�,������*̾ݞ1��&n��ʟ?�A?����O�V���m���q��+�W?zH�����鬾���=���p�=}-�>í�=���4 3�yS��0?<�3?ۉ���#���V>Dix�w)�=�OG?t^�>��3�h��>}$?�lڽ^
��݃>yx>��>R��>?7���̪���0?�T/?	�a�Tk�����>�"���Î�;e>]ۈ>��V=�>o��>/A�=��C����>�=G�=Y7Y?b"�>�1�F�T��`Ҫ�.�P���]?'�?-��>�@?kM?��ͽ���g����Ѽ�qO?s9r?��>H���־�~ľp6.?�+r?\+\>$�{��h�+�7r�E�?�f?��?V���e~s�ǻ��Y�����-?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������l�=)D��3��?_ك?�ϱ���»�n��KX����G���O=�87��i�.��I8�<�Ծ��/a��k�����>�D@�+����>�H���H�:�ο.����G��O�}���?i��>�u��I7���k��s5K��%6��e�5�>�O>�N��w��][|�ڙ:������>��	�?4�>�1V�~���������;V�>���>�=�>�Ż�tl��ff�?����~�Ϳ=���[��fY?��?#��?:?��	<�9w�Z{�Q���MG?��s??%Z?Qg��_���3�q(s?"�	��w_�D���x�}�=U �>F�>0�P���=w��>��>����3��������=�ej�?:��?�;Ѿ���>�̋?N�]?���&��.췾�IȾĤz���9?k/�>�´�l�*�h����o��=?gAm?���|D*�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>���?P>�=���>'c�=h5���*���>���=F0���?�	L?���>���=� A�+�.�h�E���Q�n��C����>�;b?��M?L�h>�E���*/��l%���½�7�^2���J��J5�����e0>�?>J�>h_L��ܾ��?�j�ŕؿ�h���'��24?ղ�>G�?W��#�t��;��9_?wl�>E9��*��!(��8e����?7G�?��?�׾�A̼�#>W�>�@�>\�ԽϽ�������7>��B?&��>��{�o�W�>o��?>�@Ӯ?�i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?mQo���i�B>��?"������L��f?�
@u@a�^?*Ȝҿjm���l�a�־�	>.c���q�=�cA��E�X=-��j� ��=�A�>{��>\�>w�>|�>t>E����"�Ý�E,���+���*���(�e�����㺾������$¾���=���=%<{���7l=:�ͼ�=�I?��i?���?gJ?�?<ϕ�=�����B�XV��޹�=vzw>
*?T:P?!]?�R�=�A��,�f� z��󁾗I��܉�>8Ł=�>���>ڧ}>9%��)V>
5�>&5f>�,�=��=8�>q�=�<x>}Y�>���>���>}c<>�>�˴��'��S�h�@�v�{2̽��?k|����J�&0���U�������=�Z.?�f>y��[Bп�����'H?����5#�b�+��W>�0?�dW?��>�����.U�R<>���Z�j�@q>{ ��!l��|)��<Q>rn?�Hl>�}>�I3��>6� <L�rɪ�9}>��7?�[��'�L��u��iH��ܾ@�C>�,�>�仑��J�������j���=:?�� ?��U���Ji�蘾c�S>:e>M�3=i��=�Q>�$K��H��r:��F=>��=��c>FJ?	�+>�ݎ=�N�>J/���O���>c�B>,�,>Q@?
%?h#��I���C���a-���w>2��>��>��>�J�8`�=�@�>��a>�h�2���t��H?�W>���g^���p��{=�����U�=.i�=� ���<��'=�~?���(䈿��	e���lD?V+?w �=R�F<��"�E ���H��F�?q�@m�?��	�ݢV�A�?�@�?��J��=}�>׫>�ξ�L��?��Ž4Ǣ�Ȕ	�6)#�hS�?��?��/�Yʋ�>l�}6>�^%?��ӾE��>Tw�P��.����u�Ag#=�:�>GKG?����Q��Y?�X�
?�?2������ɿw�I�>� �?H��?��m�}�?����>�c�?P�Y?�i>��ܾ��X��7�>;�??)�Q?�+�>�,��7)�=+?@��?�{�?��R>=��?��p?A�>2@���3�����E��j�Q=�|��[3�>�F�=������K�=m��������g�#��h�B>�-=���>�Q����ڔ=�f�kD��U\��}��>vI>J�->y<�>�L�>���>�ٛ>�h�<��z�2M��iL?�p�?�2��He��Ek=���=ĭO��@?�
3?�㮽��Ծ��>�oS?�	s?�V?�D�>�#����������D�<qU>Q�>��>i��i>ʔ��E)/����>1��>+ق<e�˾)�n��V<@��>�c"?˻�>�Q�=b+?$
5?�ƽ=��>�K�?����j�:�@>�}?��>i#J?��?[07���[�@���!0���o���o>/i�?d<?"��>����Ŕ��g=4W�=|�&�I�J?�e|?fT�D�>���?�?�h?��=�v���KϾ�V:B��><"?�� ��A�b�#�;��	?[�?���>�����u�b��oe�X%���
?Z3Z?�%?���$_b��-ɾ�/�<����';���:���>�%>0�^�g��=p%>ć�=*�Z�?'-�_��<{�=���>GC�=��#�@Wt�0=,?¿G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>$�l���K���ڙ���F��_�Ž��;BG?�e><�?f'�>��>bZ{>:cx�O����<��6�D-w����ź?���8��j�h������!g����Q����>|v6��(?�v?R3�>RU�>Ԙ�>�䝽�:�>'٩>3�S>�j�>f:�>Ǣ�>lƂ>ޣ>�\�<�DR?I����'����Q���C4B?��d?Ef�>3Wh�*���.��N�?��?�o�?:`v>bh�(	+��?�B�>�
���h
?v9=���V�<uT��'*�8#�������>Cؽ:%:�2M��;f�%a
?��?7����T̾�ֽ)�b��4�=�2�?=�,?�+:���r�02l�A�8���d��y��L�+f����@�e�}��4���v��d����!�y)�=�2?Ý?R�>��)Ծ Ϳ�j���;s}�qdw=E�3?
)�>��>�GH>�~O��U�����h"@�@�l�S�
?��?�<�><�U?�d?��(?1G:?	D�>�'�>b:Z�t��>��R�v��>��?i�1?��@?b�H?��:?��%?�%J>��������2۾�X&?���>��?���>�K�>{G���C1<9�>@s��G��cߦ�� B>��=�b=��ļ��>�hf>�?(��(�9����v�z>�8??�O�>��x�L�����1����>V�?=�>����g�<f��Q�>Y(�?�%켈^=��>R�=�4Ȼ�V���>�[��t��=�A���㿽�h	��ڐ=��=��E��F���޻նf<f3=u�>>�?���>�C�>�@��!� �^��f�=�Y>�S>>>�Eپ�}���$��q�g��]y>�w�?�z�?�f=��=̖�=�|���U�����8������<�? J#?.XT?c��?t�=?dj#?��>�*�aM���^�������?x,?��>�F���˾@�L�2��9?0�?�Na�V4��(��i�����:L	>��/�SM�����B���;�-��F��B��?���?��V�z+6��J�@����㮾�aC?Bn�>��>�a�>o�(��5e�yP���9>+��>�`Q?�ǻ>ɽO?O\{?��[?/�T>�C8�u��`ޙ���=��y">��??���?��?�y?��>��>�E*�TI�F2����X����ʂ��'P=�\Y>Y�>���>%�>8�=�ZŽ�հ���>����=��b>'U�>5��>�7�>�x>�9�<�G?r:�>J	��1�յ������ -��u?��?K�)?u	=y���D���|V�>M�?��?�5(?|W��P�=�uҼ﴾�r���>ȷ>M��>=,H=\i!>���>YJ�>u`�.���6�e�9���?�qF?��=?�ſx�q�w^p�1x��/}o<Cܒ�!e��%A[�!��=������e���\[�V���6f������b�����{�k��>�W�=�Q�="��=���<�Ǽ̘�</VJ={e�<U=
�o���m<nA8��ǻRՈ����$JZ<SI=j&�'�˾�}?�HI?��+?��C?�y>>�4�p�>ʍ���2?~�U>�`P��h��~�;�����7��~�ؾ�׾o�c������|>$�I�F�>�^3>i��=�|�<�#�=5�s=<�=D�M�ٯ=���=6,�=7��=x��=j�>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>9�C>~>��Q��P-�m�D�9M�1-Q��0%?;5��%޾E�z>^��=�ݾ�ʾ4==-<>@��=�m/� _�e��=��f�K�`=��==�7�>��4>��=�n����=V�=���={�b>ba�;>j�(���ъ=#�=�Hz>`1>̌�>v�?Pf0?Od?!A�>R�m��Ͼ�+���B�>���=pA�>�Ӆ={B>Ǘ�>��7?g�D?�K?~e�>�6�=��>!�>�,� �m�Y�̴�� �<��?xɆ?��>�Q<��A�2��	W>��Ž�{?�W1?�x?���>���8�Կ��@�.�9�(\>Wl�b+½�y��Rm=DQ�=�u!��j�4{>�?��?7�>eS�>�?�֗>B	�>�=�\e<Y�>G�$=W�;=
Q�j>f<)�<��>x=�>B��=qG��%5����<^h]�,p��ڕ����=��>�<>���>/n�=r���1/>lĖ���L���=!B��D,B��0d�cK~�%/��]6��B>�%X>1���l2����?Z�Y>�n?>���?|>u?"�>|5��վBR���Oe��gS�ٳ�=��>8�<�#x;��T`�9�M���Ҿ��>i��>y~>���>��L�?LJ�N@��:�ƾJ�8�f��>�[�װ�;%�˽d.i����	��W�b��1?��#9?����>���?Ee?�2�?r�>(3��~+���r>]��/��.�%�Z�!���i�G��>�H2?
�?M���.x��	̾0p��騷>wI�7P�[���0�0�4!�S偱>ʪ��о�>3�^j��i���p�B��s��>�O?��?|@b��K���'O�����s��x?Ћg?�ן>�H?wm?%ע�9%�M���z�=��n?��?�1�?��
>��=������>�?���?Y�?��j?4Y�׊�>���<
I>��'>=�)>^�=�M�=�[?qW?Rd?���32�g뾚��Z�^���T=Hu�=�y�>%<�>Lم>"�=s�g=���=��\>QӜ>�}�>�(u>�E�>B-�>�5��w]��T@?.�*>�G�>�kF?L�7>;*;���J>P�ǽN�.�0�9��3Y=A꽃�?=(��V����V<k��>�ʿ#�?�1�<Q���^�?��Ǿ٠(>` >�
[>�v��ػ>��>� >1��>�*<>�:2>�ur>" N>�CӾу>���Ge!�N,C�ނR�5�Ѿ�vz>ҙ��&�[��i��}KI�%q��5i�\j��.��;=���<�G�?0���>�k�:�)�{���;�?	]�>�6?�ތ����_�>	��>ȍ>�H��C���&ȍ�+k�E�?>��??c>y�>i�W?�?H�1�3�puZ� �u��'A��	e�>�`��፿������
�s����_?*�x?�uA?E�< 8z>���?>�%��ԏ��.�>e/�%;�Oa<=3,�>�*����`�r�Ӿйþ�4��KF>��o?0%�?�Y?8PV��2
�)iO>�?H?\�'?1�l?�-?hJ=?��Ƚ�g!?�qC>��?n�?�V2?ʓ4?�C?��~>b�>�2<�=��:���͒�������U�"�VA�=���=r����{=\�=,�;�y��08����;t���N�==�|�=K�=s�=`��>�]?O��>f{�>@�7?����8�\����-/?8�1=���=)��p���&��G>:�j?K�?o�Y?L�b>B�}�B���>��>��%>�F[>�>�� QE�r>�=2?>��>���=8�H��P��gn	�� ��T��<��>h��>�2|>r��B�'>�}��3z���d>Z�Q��̺���S�[�G���1���v�}W�>��K?��?u��=�_��.��+If�0)?�]<?OM?��?��=��۾��9���J��@���>�9�<���3����#���:�+��:E�s>q5��j����f>����޾�n�KvI�����X=���[=T�
�&_׾�m{���=X�>�B¾�� ��[��f;����H?�t=�آ��Z������>і>���>0�^�4����kC�����tۅ=ô�>�4>G��uI�V�H�I[�傆>�,G?:~W?�n�?g���ro�&�>�3�����S-�zA?8q�>�?��(>�u�=�ɼ��^�q�g���>�[��>7*�>
��dH�d(���Wվ|&�k��>��>�5R>`w?�`L?��?�-c?)5?g�>���>c�X�ׂ����&?TX�?�*(=载�Ys���8���D���>�(?�W6��=�>�?@w?�$?k�R?�8?���=>d �3;��Ô>�K�>�OV��]���Y>f`M?o��>.�[?�Q�?��L>w�-�����	���h
>Y�6>��,?	�)?/?��>���>N������'B�<���>�/�?�?��(�K�<��?9O1?�t���Y�>��+?T��>:�A?�e?WS?)-�>{������!����}v����v�<},l>>	>z������$kV��<�<)2��H��#T$��{�����=^���k�>-t>�)���0>žQ����@>%ˡ��9��XĊ��r:�΋�=��>.�?�͕>�q#�(i�=�z�>�,�>z��g3(?��?��?�TE;&�b���ھ��K��հ>;�A?�W�=g�l�=����u�9�f=��m?<�^?&�W��T��1sa?�q^?N���&(�����Z�����&�B?�?v��ӏ�>��c?wfi?^ �>�.Խ��p�rϗ�@ _�H9D��5�=o]�>�d�{0t��r�>~�B?���>+x�>��&=�þ�q�/��"<?7w�?��?7Qx?ڰ�>~Ur��Vܿ:3	��׃��{?�O�>�f��<3�>7��B<���������m���Ͼ��t��{x�"ƨ��E������K��U�c�-?%tw?[ߌ?2R�?_r̾�;�pp��҉���Z�Ӑ�	�$��K��:��:��g�������1�RF律�<,Q������?��:?��]�*�>|��5���󾦳�=5�Ⱦ.q�m-�=P�j�l�&��+��
��8���u=ξ��+?j�>�]�>��G?E�:�C*�x�L���H�Pe�v�)>��>^��>�9�>b�H=�!�m�C��m�������Ƚe}�>J:e?ݨ'?��r?�s�S�:��Jy�u�&�����cǾ���=k�=�|q>ǘ���0�(�&���U���x�F��������������<�?F��>�:�>(��?JE�>]���i��f�b)��u�='ڡ>W�}?o�>�̍>�$9���v6?�Ww?�Y!> �>2��ѡ:�����*��=��?�ڽ�ؤ>C�>^���L����Kg��<V����>���?�6�������p>�3W?�ʵ����=�?��"MT�<���e&L��D�>E5?$�<|��>O�ž�é�6�|���8�('? E�>�����.�	�>#*	?Q?�S�>xÍ?�;�>���|xb>��
?��+?�\b?�]P?�N�>PC>�j��_;���5�o��<Xӊ>�~v>)?P�)Ԡ<2��"�7T.��1�<5-E>q'�G��Ib=~���jĽg̻c>eۿZCK�h`پ� �[���4
�9�������.��8��ہ��M����w��.��d'�m&V���b�F�����l�m�?%7�?B����<��ٌ���s��������>N�q�����Q����Y&����ྩ/��uE!��P�!%i��e�Z�'?>����ǿⰡ��:ܾ�  ?�A ?O�y?��O�"���8�a� >b<�<�0���뾢����ο
���"�^?���>��/��C��>�>^�X>Iq>����螾q0�<��?K�-?	��>�r��ɿV�����<���?"�@�tA?,�(��~�éV=Z��>	�	?_@><�1�yU�ϰ��s�>�.�?4��?`�N=0�W�z��ہe?�!<W�F���|}�=�/�=�z=��|�J>�L�>����9A�)t۽��4>���>�|!��g�]�^��|�<�]>�~Խv����Ԅ?�y\�cf���/�#U�� V>�T?�.�>-I�=��,?�6H�~{Ͽ�\�4(a?�/�?-��?��(?�ֿ��ؚ>��ܾ�M?�B6?���>Yd&��t�ݎ�=-!�QU�����(V�	�=w��>|>�q,�b��͏O����c��=����������^,���<�x���^�^��#s��P��^���g��w�>ȼ=�Q�=�:.>.ɍ>�IM>H%>ƿS?ʬr?C��>%z>�Y���h���˾�%���O��ie��壵�n�[�斾����������M#�B���U����<� ڏ=�ZR�'v���� �R�b���F��.?��$>�{ʾ�qM�ݽ!<�ɾ����-p�����[L̾��1���m�\��?'�A?̸��>W�j&��,��h���iW?2����Q���j�='˿�	�=�K�>Cڠ=�T��r3���S��,/?{ ?�����.���>/6��W>�*@?o�?�J��Z*>t�I?I(��pg����>Y�>��>b�>�؀=1H������E�?ճ<?h������_0>@������Oy_=C�h>Q���<��>�z=K�����l��gE�<�Z?�_�>1�-����B9��xc��|����?�??	\�=��?:fW?a�V��U�H�h����E8�Z�V?�)�?T�>u볽�T¾r�����0?�P?8�>u/��[쾒@$��Z��g�(?�	P?��1?,XǼ�To��쉿f�Ѿ�;?��v?s^�ws�����U�V�f=�>�[�>���>��9��k�>�>?�#��G������vY4�&Þ?��@���?��;<��U��=�;?o\�>��O��>ƾ�z������m�q=�"�>
���yev����R,�h�8?ܠ�?���>���������=󬗾!��?��?�S���<���k�����Dd<��h=��L�{�0����d8��˾:���}��R���%�>��@{�� ��>��,���t�ο[���\�ξ�d�_L?�p�>����֧��qn��x�2H�
�G���z�>;�>�l��oC���~|��m;�m<�����> ���>��N�/��_Þ�0� <c�>�`�>_z�>�$��\����Q�?����¼Ϳ����r�Y?��?݂�?�?vz<W�q��!{��4ʻ�
H?�/t?�X?<	�ի[���=�7�j?-^��kU`�7�4��GE�nU>�!3?
D�>Y�-�;�|=�>���>�c>�#/���Ŀfٶ�����I��?��?�o����>A��?�s+?7j��7���Z��M�*���.��<A?�2>���t�!��/=��В�!�
?7~0?�{�I/�K�_?�a�/�p�p�-���ƽ�ۡ>��0��d\�3F������Xe����}@y�|��?5^�?y�?r��� #�T6%?�>A����8ǾF�<v��>�(�>M*N>]G_�U�u>��!�:��j	>���?g~�?�j?Е�������V>��}?�9�>��?�^�=Ӄ�>��=�"��^�0���">
�=O�@�z?ʅM?0)�>��=e�8�O/��{F�\R�a��C�t�>�a?[L?8�b>2븽'r0��� ���ͽ��0�`鼘~@���+���߽`�5>;>>�G>�6E��	Ӿ?�?�n���ؿ�i���l'�E44?���>�?���N�t����O<_?Pw�>�6�T,���%���G�O��?H�?��?,�׾M̼>u�>K�>��Խ����������7>I�B?��D��.�o���>"��?��@|ծ?�i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*n�Կ����j�Ӿ�N���R>ٰ�<�G=|[�S'�=r�#>@��)F��-�>Xe�>ڼk>�Ө=��O>4>V�>o����!��K��w���-�4�U4"�t,��������/�P��������#g�����b��#5��a.�r6�ٙ:���>�la?	�b?xPp?�k?�<�+>���J�;������X>7ܰ>В5?�]J?E�$?���=��^��b��׫��H�����>E,^>��>��>��>�E���=���>��>�B�>�A�>�M>���h�>� �>�b?^��>u�<>��>~̴��!��:�h��w��̽��?�x��l�J����;p��\����I�=�m.?_�>(���@п2뭿�H?�Ô�	���,��>��0?�EW?`t>�`��1lX���>�q	�Yk��� >z� ��l��c)�dPP>�?",g>��u>أ3�!K8��P��u��9�{>�6?j򶾁�9���u���H��fݾ��L>xؾ>ieO�h�$��V	�.ki�ݧ|= w:?X`?�T���t��{u��1���zQ>1-[>��=���=�zL>d�e��~ǽ��G�pr1=Q��=��]>�?��=[�=�Њ>ꌷ�Y/0���>��>X�>h7?P\
?o�<�4"��G��Ɉf�Ǹ>��>(.�>�&�=h? �j��=J��>.<|>j�̸�p����}����>�׽}��ɇ?= � =���7>=��c�XP2����=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿym�>�\��Y�����b�u�`U#=��>�<H?�B���P��>��w
?�?td�#���N�ȿ�v����>�	�?��?��m�p?��@�P��>ǡ�?�hY?fsi>�e۾�aZ���>��@?R?b$�>�7���'�?�?�ݶ?:��?��Y>`֐?��b?���>'e½�73�Sq�����}�=d����O�>[�=����TK�$ӎ��(���r��Q�6�b>(X==`�>�1���Խ����=�nD�C ��c;��p�>Е�>��p>��>g
�>]�>X�>�S=`���7�r�򀑾��K?���?�~���m�Ӧ<!�=�%`��7?(�3?�M�;~ξ���>�i\?fu�?�C[?š�>���ya������#��u��<rM>���>���>�!��ܖI>wԾ�H� >�1�>�1̼L�۾zM����H�>DJ!?�i�>T8�=�*?�M?;�b</��>E�#�	ޝ�W�����>ٸ?\��>��?�>�D;��k�K�������<cz��>'��?5�?AO�>f���О��n>
�f<_��DB�?%�?E".��4�>1	|?�7?��@?9q�=�S>�`����=�?C!?Q��q@�1�%��2�L??�?[��>	@����ʽDy��V�����?�[?y\(?�E���\�$���8<�<i���y���ޜW<�>���C>�i>Mz��_�='>K��=ճ`���4�e�;q�=t��>���=�5���y��9,?q�I��݃���=��r��bD�FO�>�GM>V���f�^?ѻ>��8{��欿Z{��8eS���?Ut�?r�?]Ӵ��gh��	=?���?��?>B�>6ӯ���޾�P��Xw��x�`�ȓ>�}�>�Rq�}�����"����A����Ž�8�<+?`t>�O�>ҕI?��4>"R�>t2.��:+��H�#�qq��3�M]��7�۟�+�_��M�2��������e�4�>�n�=ޫ>W�?�]�>�ȋ>(�>'g�A�?Mn�>q��>���>�fq>L��><*�>�n>)ӽ{KR?����b�'���辽˰�RB?�Yd?z=�>��h� ~�����o?Y�? g�?��v>Syh�v++��N?�>v�� p
?�:=Pq���<W7�����)��2��Ce�>)�ؽ�,:�wM���f�N
?w?���ɻ̾�/ؽ@M���a=�ɍ?zL?]G:�n'\��E��t�S�R�M�mpK�����)!Ѿ)�T��g��U����q��Ԕ��8�7�xf�=��8?���?��^�ɵ����Nt���l�C�u>�Y"?H[Q>��>F�b=ڼ\�b�J���x�ΑJ�l^u�rq�> ��?F�>/QA?�Q[?7�A?;�I?m�>h��>h1�|(�=I�>���>�o�>6�V?��=?�3?,7?7�6?7c�>&yD�>'ھ����.�>݌�>�\�>��0?-�?�C��v%��+�w>��<A�Ծ����>�*�Py+=�7�<�*D>���>�=?7���b8�z[��%?i>Y�6?��>��>儍�E������<]�>�j
?��>1���'p��z�o0�>�с?����O=��(>N�=���}`�����=�᡼R)�=ڴu��2�x$<��=d��=h�����%�e�(90��9HY�<u�>�?N��>�C�>�@��?� ����i�=�Y>�S><>pDپ�}���$����g��^y>�w�?�z�?�f=�=2��=}���U��V���������<�?�I#?�WT?A��?��=?j#?ʵ>�*�`M���^��/����?e",?ј�>�����ʾ�꨿�3��?YW?�<a�6���A)�ʢ¾0ս��>�U/��2~�m��C!D��ǉ����hW��B��?M��?@��6��c�۽��Sf��K�C?��>yP�>���>Y�)���g�"�P;>���>�R?6p�>C�O?WL|?J}[?t�X>�<5����ud��LE˼�g&>5�@?4m�?YP�?ox?�w�>�j#>����Gھ���y$��| �}l���1=s�T>��>̏�>w��>�r�=�	���w���UK��X�=[�d>�U�>1�>q��>�W�>���<�??���>2���_�ﾩ�ᾼ'K�� >�Q�?8N�?Z�?�ݽ�rľ�o�i����?4��?�ט?jh:? ����=��ؐ��B�o��@�>w)~>"��>��=%ߒ>}^>�s)>�F?�2���i�¿Ӿ!^g���>t;F?�=_,ǿ�#v�~G�� F��7�b������aX�0h�XN.��s�=�u��<Ͻª����J��0����������Q͡��烾��>r��=0�>?��=vUڻQ���w�<sj�=�)=���=�3���ȍ�-}�C�u�Xz��c���==O ="�`<�˾�Q}?��J?�i,?k&D?�|w>o>�:O�=M�>j��3?ߔT>7�C��G����<�t�������ھ�uؾ��`�rL��ل>u�P�څ>�M2>���=��<a��=�ix=J'�=��::�=�
�=?�=���=E>�=t>==>�6w?V���
����4Q��Z罣�:?�8�>�{�=��ƾn@?{�>>�2������xb��-?���?�T�?>�?:ti��d�>I���㎽�q�=\����=2>���=n�2�`��>��J>��� K��5����4�?��@��??�ዿ̢Ͽ?a/>��:>&�>"R��0�^�B�c�9�P�#?�8��M˾�W�>��=�=ݾ��Ǿc�O=)<>T[=���ιZ��r�=��t�{�4=#�l=���>�A>IU�=�����=��8=���=��Q>�����Y9�� �Q==��=fR]>�&>0e�>�?~�2?��c?s��>��b�}Cʾľ1�>{�=��>���=��P>=�>�i6?�F?�L?/^�>�t=�۷>F�>�0*���m�:�侅��&2�<���?�p�?��>Ё<�CQ�n��Y�:��۽��?�e2?��?b�>9��ё̿x��g����(���9'��!��z�X�>2{�>S�)G>Yu>~��>w�>�6>{�>e��=��(�Q�>��)>��=؍�=\A	��=B�7>��>>�׼-<���;q'!�4�M���=�o]���<��=�J,;�$�a��=|��>y�>`��>���=����.Z)>�����L�&��=����&�C�D�c���}�/�,��3?�!�<>�F>����Z���N?��_>o�<>���?�u?��$>?� *پ!&��)Bq��V�^��=M��=�F���:�e�\��?M��$վ���>X��>\��>�7p>��,�N`?�R�i=�_⾨k4�6Q�>c����� �=�z;q�-᤿�䟿��i�Ƥ��D?����X�=��|?�{H?@h�?�`�>�Q��=(ھj
+>�瀾Ц =D��9�l��z��k�?,*'?t��>a��X3E�I7̾�̾��̷>}I���O������0��7��Ʒ�v��>��@�о
 3��f�������B�=qr�8ߺ>��O?�?�:b�V���WO���܅��h?�}g?��>�R?M?~%��~g�<R���=��n?W��?�9�?>~0>�ý,\?*Z�>QM�?'�?�t?����X0>,1�>���>B�k�y\$>�I�>���=�ȱ>�b$?4T�>���>�3��m���,�ט뾷w0�)\>x�>2 P>��>*�T>��>y��<+��#�7>���>��L>�q�>�ɻ=W�v>�対@��SQ?�<_>��>��?ٺ>�TE��L�`$W�� �98��c󽵈N�����Y�����A�+���wٽ��>�?ѿ(�?Rei=_�.��|?:����=8�P>)�M>Z�ý4,�>ä�=`��=O�>���>��	>�I�>��y>SFӾ~>1���c!��,C��R���Ѿ�{z>C����&�ӟ�w���BI�|n��Ug�/j�7.��<=�B̽<H�?����Z�k� �)�
����?�Y�>�6?�ٌ�T	���>���>yƍ>:K�����ȍ��h�*�?���?�;c>��>=�W?�?m�1�'3��uZ��u�o(A�8e�V�`��፿����
�n���_?�x?yA?P�<:z>F��?��%�Jӏ��)�>�/�';�[@<=l+�>*����`�a�Ӿ|�þ�7��HF>��o??%�?}Y?0TV�=�j�'j%>{>:?�>1?��s?�M2?��;?v~�iQ$?�4>�R?�3?aG5?x/?��
?��1>�<�=[/Y�F(=sk��ء����н�_˽A�����/=�z=w	�9�|<k� =��<��01ټɰ�:����sI�<8�<=�`�=>
�=��>9]?c��>��>�37?����7�*A��Hb/?!�==����왈�d�����3> 9k?܏�?��Z?�<c>>.A�U�B�qh>��>
)'>1Z>c#�>���
E�~�=Ji>>�2�=y�G��H����	��j��格<��>��?�.�>h�U�IS�=���������=����`ž
���G�6�P��K��c}�>��H?�O�>/����o0�X�O�K�K��k,?]D?e�?��?(�4>�~����3�<�g��߾�D�����P*?��ͩ�(Υ�gG0�cG�=^�=���z��8�a>T��ܾ�?o�}�G��~���I=�l�Z?e=����Ӿ�\v�v��=$�>@�����������%J?�V=￣�m�V��=��Mu>|�>���>:�*�߸s�GB�����j�=��>�J=>@J��+C� �F��H��D�>�RE?�7_?5j�?p6���s���B�J���E<����Ǽ=�?���>�b?�B>Z8�=�����x�d���F�B4�>���>���1�G�]c�������$�!��>�I?,�>��?׿R?��
?ѥ`?�*?L?�k�>�׸����^f*?���?�B�W���^헾��'��+N�f"�>0,4?)��6>�>?�)?��)?!X?Ph?u\9>�	��01�~��>V~j>"sH�#s��4>��K?���>��9?��?Nga>cF�����H���>ݯ>>C"*?,'?,H?"Â>�>��+���=�}�>�i�?� v?&�?�p>���>�!�����>ݔ>�P�=Zg�>�<?�8?Y�k?ԍa??;�>���Q������ �e�}�d�K���g=�X�=W��< s^94Խ�$���</S-� �?����<�d�<mh����<�"�>�=Z>�Ԗ�q+;>do;Iޞ�D�>��<HŤ��U��뽡$�=-2|>�4?N��>u�
�>�=��>B�>Z �7(?�?l� ?Dk�$�`�3�ž�y����>a1?Z~=�n��ґ�Zs�6.�<�]?Fg[?�?������N?TIW?P���a���Ҿ&K�(��y=?,j"?X1=��=>SzX?���?k�>X~1��.����:Q�=����k>9D>W&��/�y�bJ�>�CV?<��=�����<)�����I����l�=?W®?Q��?��?[P�>E��Ք�ϑ�-��x{]?���>����rX(?��':����\¾=�n�L:������¾����2���Z4�c�j���5�!$>Ҏ?�}?D�?)1O?>L�"�`�2r�=Z���U��ʾ>���6�!�$D��G���l���(�޽�!Ϧ�ջ�:�����I��з?��?(S���>[����
�����O>�.���\���	=&+����;k6�D�x�*�P�FǤ��#?=k�>��>c�2?ЦU�#<�{6�:�0��=�o�:>̖>���>���>Z��;��8�_S��iξ�Dg���
��6v>�vc?k�K? �n?�Z�;'1�0�����!�0�/��j��4�B>�g>���>��W����9&��Q>��r���3x����	�4�~=w�2?�1�>���>SN�??{	��s���Yx�̄1�ւ<�&�>�!i?�:�>�߆>A�Ͻ�� �T��>��l?ݤ�>��>�����Z!���{�תʽr �>�֭>b��>�o>��,��!\��i��i���Z9�>�=��h?Ń��t�`���>)R?��:y`H<~�>�v��!����ս'��>kw?�v�=U�;>��ž�$���{�^0���?K?7�?H���W'�T$����>��=bs5>k$�?�h?R?	���N>�NQ?�D�?��H?��E?A6�>����˾^ ���qu�c,=$r}>�>��=���U>h[��N`��?�9��>�Et=w�B����x���`:=���͋+>�>�=�|ۿ�^K�1پ�������	�����w$��{釾[S��״�z��s�x�T��P�(��-V���b�Y�����k��|�?:�?j���n#��h��������]����>vr�6N{����q���Q�����p���8�!�NP��i���e�J�'?d�����ǿᰡ�:ܾ  ?`@ ?ިy?����"��8�#� >CT�<7 ��?�뾞����οQ���6�^?���>$��+�� �>O��>�X> Iq>*���Ꞿd,�<��?�-?6��>�r�T�ɿ����C��<u��?��@�IA?^�(��^�_�F=���>�F?�:>6!+��� Ȯ�DV�>z�?rÊ?�TU=n;V�����c?A�;-[F����N1�=08�=�0=˹�}F>�(�>�$�UbF��P޽�@9>��>0�0�<����\�*��<I�X>�2Ͻ𙍽5Մ?+{\��f���/��T��U>��T?�*�>\:�=��,?Y7H�`}Ͽ�\��*a?�0�?���?%�(?;ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���={6�#���y���&V����=Z��>f�>Ă,�ދ���O��I��R��=��#�ҿ�9��B�N�=���={8=R@V�͙S���R���~����R��L��=Ӿ�>޲>Dv>�Z�>\�Y?ӿ�?o�
?l�>?=�+����[���I��/�����b���9�F;�<��E��f�4�ޔ0��F(�ř����<�ύ=Q:R�h����� �ѻb�{�F��.?��$>��ʾ
�M���2<#(ʾB����[�����X>̾	�1��n����?��A?�ꅿ�V����#)�5i��	�W?��б��������=�c��aY=�-�>�ˢ=���f3�YYS���8?��?����d��D >A�����i<��"?
��>�	>���>5�A?�ѿ���>1�>U��>S1�>iަ>B��<ھ��D���$?]�g?'�W���ؾ��^>�E���ھ!����t>7�b�O]a��[=��������I��E�=�!W?bt�>\�)�+�2`��{X���;=I�x?�}?�:�>A�k?��B?�<^B��ٹS���
���t=i�W?Ni?h�>B���*�Ͼ;&����5?�~e?;�N>h�q����.�%.�0?=�n?*P?����"c}�b������p6?��v?s^�ws�����=�V�f=�>�[�>���>��9��k�>�>?�#��G������xY4�$Þ?��@���?m�;< �R��=�;?k\�>�O��>ƾ�z������@�q=�"�>���ev����R,�d�8?ܠ�?���>������>��=�ٕ��Z�?{�?|����Fg<O���l��n���~�<�Ϋ=��}F"������7���ƾ��
�	���oῼإ�>DZ@YV�q*�>,D8�]6�TϿ"���[оUSq���?I��>��Ƚ����E�j��Pu�Z�G��H��������>��/>����|7z�u�}�^18�$.1��;�>2
�<��>�$��ʜ�����<�d�>ݠ�>G�>�!Ƚ���5�?���ƿWD��"���xa?�%�?3?}?|('?��=?`���Qb��Ǧ=S?�t?�\?��=T���Vɽ#�j?�_��vU`��4�vHE��U>�"3?�B�>U�-�|�|=�>���>g>�#/�u�Ŀ�ٶ�C���X��?��?�o���>p��?zs+?�i�8���[����*�Y�+��<A?�2>���H�!�B0=�[Ғ���
?U~0?{�b.�`�_?�a�P�p�|�-���ƽ�ۡ>��0��e\�II������Xe����@y����?D^�?Z�?}��� #�R6%?6�>w����8Ǿ��<���>�(�>�)N>IJ_���u>����:��h	>���?�~�?Nj?땏������U>��}?Q7�>��?�H�=ZZ�>/��=�*��Ҷ'���">���=.N?��?�M?e�>�)�=m'9���.��F�r(R��)���C���>��a?V�L?Lb>4����2��� ���ͽB(2���뼨�@��.�6�;�4>�=>�>��D�ۣҾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>D�Խ����[�����7>1�B?Y��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?lQo���i�B>��?"������L��f?�
@u@a�^?*��ҿ����p���ꪾS��=���=�l>a��0{�=�"=NY@=);��>c͒>K�>���>Z#�>�"@>>�T>����%�i:��(<��_�O�%>�ߩ�7ک�����d��������֩���ѧ�7ƽ������,�^�Q�$���vi�=��U?�Q?u�o?� ?�?z���>k���9r=�#���=�7�>�?2?ÌL?hV*?v��=  ����d��R��>[��T������>��I>m��>�5�>�>)��8~AI>Q>>�T�>_ >��%=��"�+�
=�LN>�>���>(��>�T>���=M���a����Y��m��G�0�}i�?u���1��J���ZV��a��I"�=��/?�|E>ߏ��kPɿ�s��`=?i>��/Q��J|�Qs�=�?�P?�wp>]�׾���Ul>"�ݽV������=�Ƚ��F�Z�<���v>1�"?&i>^�r>��3�c�8�P�V���u>��6?�"��k4��xt���F�3�پKO>��>����{�����c~��Qh���l=��9?wX?�۳�����³r��~���jK>j&Z>v-=J&�=�qH>�.g��Ľ�E��)=w�=Eda>�s?��>d%=#ӟ>[���҉�zp�>�fZ>)Z�=w�0?�:)?�iH=c�:�m_����>ٽ�>��\>��=J�k�J��=�d�>[�>�_�����
����i���>?��/�U��3н{��<h�޽�j�=�j;�����s��x�=�~?���(䈿��e���lD?R+?^ �=I�F<��"�E ���H��G�?r�@m�?��	�ߢV�?�?�@�?��H��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�0)#�iS�?��?��/�Zʋ�=l�6>�^%?��Ӿ�^�>G�V��&��w�u��"=��>�>H?�+��-tO��>�-h
?$?�p򾪮����ȿ
�v����>~�?���?��m��>��@�
��>���?�TY?6i>(W۾�$Z�ou�>X�@?�R?l-�>X��*'��?}Ƕ?|��?�I>d��?��s?�m�>A4x�<[/��5��U���'l=6�Z;�c�>�U>����GgF�jד�{h��+�j�&����a>�$=�>=J�L4��4@�=w싽�H��6�f����>�/q>��I>X�>�� ?v`�>���>�w=�f��JှC���AS?�Kx?�&������ ���:>�?���>�_C?ځ>Rd;��>1qy?+{�?/@Y? �>F#��#{��@��K%���L�� �>>^��>͔�>zQ"�AYn>�.����=���>��>�S1>�￾�ϻ������>��?@(�>�Ă=)�>��2?N5�<�M�>��F������r�
?�?P��>��B?��>�Ҿ�Z=��c���e����j�M?�ٓ??<5?�ˢ>4������y�[=��$>���w�U?X�?�F>ߜ�>�X�?�ۃ?a1=?'`�>�8*>�ͼ���\��<Rq#?ʜ�4<C��+(�X&�F�?+w�>E��>^�n�p����w���D��37?
�]?O�(?|����_�Rjľ���<w�˼HQZ;��=)>ȼ	�>��%>�lC�<�M=�>{�=d�\���I�'J�<'/�=�>RK�=�&�Əa�(=,?��G�wۃ�W�=�r�PxD�P�>�IL>!����^?�k=���{�����x���U�� �?��?Lk�?1��A�h��$=?�?m	?("�>�J���}޾k�ྑPw��~x��w���>���>ݩl���J���Ǚ��F����ŽҮ��2�>ߝ�>k�(?�?h�>�a�>�u��N���B%�����<��q�7<��#����C�r׍��v�=<1����J�?>0�����>"�?��>��5>�>�býKi�>
G>�U�=�6�=k͆>q'�=3�<��>�L;nHR?����;�'����6���WB?Xd?�E�>$"i�d��$��_?9��?Um�?�bv>�gh��5+�d?B9�>���Df
?�g:= �
��
�<�Y��̋�;��������>�ֽ:��M��pf��e
?$?O���p̾��ֽ�B���<��?� ?�������R�-t_�+P���l���3$ ���J�������_I����=��O�>PRA?	��?���w�Ҿ,��5o��Q�1���>[?*��>u�>Y+>B��k8�5y��b3��b/���7?P|?�d�>��D?�m4?5�L?�hG?lgl>���>Iܰ�A��>jS��N�>EN�>h�+?/1)?h
!?M%?�I.?�[S>{�d���о�k?u�?�?�n�>�b�>�7x�b�Խ9y���X��nV��#Jƽ��;��<�+����<Z=��m>?�e�T8�A���o>&�3?�_�>��>�ҭ��*��;��>�??m��>�u� do�%����>��~?����L=�F.>�v�=�3�$��/f�=I�&���Y=��������<�=�P�=bu���:[*S<�W<c<fq�>��?Г�>pH�>7��� �I���m�=u
Y>�S>�> EپI~�� $����g��Zy>gw�?�z�?��f=��=��=-y��oU��M�����g-�<e�?�H#?�VT?���?��=?�k#?W�>�)��K��<^�������?[�+?S�a>���qľ1�����<��<�>�?g�b�|����󾻍���ܹ�W7>C����_��|����9�0�<a2�JPt����?(T�?���V�;��վ�_������~�-?H��>k;�>�o�>�q��Yd�iS��l\>c��>M�K?�#�>��O?�;{?�[?kiT>|�8��0��0ә�J3�I�!>g@?���?l�?uy?�s�>��>��)���!T����t�߂��W=<Z><��>�(�>�>!��=OȽ;S��j�>��X�=�b>x��>'��>� �>͆w>^U�<Q�G?���>����������Z����?���u?��?c�+?i(=�\��E�� ���h�>8g�?��?N*?��S����=\�ؼ�¶��kq�o
�>���>\%�>�ʓ=E=�T>T�>1��>�8�eO�UU8�2�L���?�F?-��=s�ǿ����ey�>F���1��=Fp`<����������=:ˈ����7dо������ܾa��X�Ҿ�䯾��Ѿ9��>���<
>:�>����x��=�6{=h�w>%M>3]N���]�[G����� �F=�����r,=f��d��=�ҽ�@���1w?ӗ=?B+?);F?�lp>�S;>;�t���>g�̽��	?�nc>�1������*R�B��	�g���Ǿ�d־o�a�pő�"@>!AZ�U�>l'>���=�L��3�=��=s��=B÷;��=�'�=�~�=���=8��=Q�>: �=�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��=>�_�=�CQ��-��JM��3j��@W��� ?�5���ľ�^�>J��=
-Ծ�����=[@>ԺV=��waW�(+�=��w�x
�=�_�=h��>7.>�=�᭽��D=-�M=�>�NX>y���#4�%4�~�/=���=zCj>2b$>ǈ�>X�?lY0?�Zd?�X�>��m��ξ�1��%2�>�Q�=�O�>� �=~B>�x�>��7?�D?;�K?���>�Ή=��>K�>�,��m��G�-����֭<���?�Ɇ?_��>��Q<J�A�9���b>�9Ž&t?�N1?�g?�ޞ>�U����9Y&���.�$���Oz4��+=�mr��QU�O���Hm�2�㽱�=�p�>���>��>:Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=(�����<�vż�����u&�:�+�2�����;w��;A�]<U��;�4�=}o�>��	>K��>�uR=�˾8>�F��lmB���@=�����v=���[��n���*���<��&5>{WG>�5�y���m�>!C">�mT>p��?��s?��Y>��쯾�ʝ������턾6u�=�M=��e��=�<�V�ȿ@������E�>(�>(�>��>��/���D�8~=�ھa�5�Qo�>=����H����4l�nq������!�m��<�<e*G?Il��a>�Bt?L�I?nc�?O	�>J���!۾?>����+0;��7�����ar?z�?�W�>��߾�:���Ͼe����Z�>,�>�(	X�����#!-���l<����pݮ>j:������-?�;X��cs��7aP��q�����>-}Z?��?�R��!��4hR�c���|���>�v?D�>eB?���>IF�Ѿ����o��<�8`?��??��?Q(4>��%=�=���>�~-?�ƥ?Ap�?�?�^=�" >1���A��=�3�j��h�ymi>aL�=W �>�Z:?��?�P��c��$������r%H�A�R>@�*>.�>�3�=�e>���=y�ļ�)@>�>��>p�M>��=��U>�g�>�ﶾ���F�1?й�=Hƍ>W4?c�g>u�;�L�ߨ�<��k�<jO���6�kG��?���܌�
��/�"=H^V�p��>��ƿ+�?ܳ[>Y����?��边-s�mc[>��%>����>� 9>E�s>��>�å>�z�=�؄>�Q>��Ѿ��>H���:���C�[�S�0�Ͼ�z>�؝���*�sp��j����I������z��i�+˂��:����<�?m�ܠk�o�'�� ��}?"�>44?(������7>٢�>�0�>O���.딿�ύ���⾭��?,J�?W;c>�>F�W?6�?��1��3�ltZ���u��'A�e�0�`�����������
������_?�x?]xA?I�<8z>ע�?%�%��я�+�>q/�t&;��=<=�(�>�*���`�p�Ӿ$�þ�9�]KF>@�o?U$�?wY?�QV���l�Q&>k8?��1?7u?� 7?i�@?�\��3?�>5?Ŗ?�<2?��(?�:
?#�'>���=<�<ݡh=*Z��3C��Y8����ν� �&v=��L=i ;ٷ ���#=���<9���<���I���`"�9�=<��X=��=�a�=���>[�Z?��>S�>E{;?�b�n�(��˭� j'?�5�;V��8c��{2��^��cx�=�Z`?.A�?�XV?�vR>�;D��5��]8>b�>��">B`]><ާ>Os���S�Ϟp=at
>7]�=cӘ=Z�y�
�n����cc����=U�$>�k�>3A>����C�>0�Ͼ���V>��ͽR(��awb��}�/�
��d\���>�~-?F?��9킿�d����q���?(�
?�a?��S?$��=;I���<E�׃��վv��������p��ٌ��uS�0�ݼ#�~>ҀսT���E�O>���&�dbm�ZF����w"=���n�u=�;���;�|��&�=���=�����!���BS��WK?@4A=�{���K�6����^ >d��>��>�8�ԂX�K�=�a���4O�=�3�>tK>�v-�y%辒�F�RQ��؃>��H?�P?���?��J���w��i>�.s��~R��3=��?ch�>�!�>�>jr�=8���r��f�[��s<�)"�>|X�>�h��H��ڵ����d&���s>^?��b>t�?SDW?��?^�e?�]0?
�
?�P�>%����Q��()?�?Io�;���lу�����V��L�>�e5?�D��7�>E�?4�)?r�8?+�^?]�?J-#>��o�4���>car>s&8��}���^L>�q\?�>�-R?b|o?�v>͟>��Z�����Z1P>��1>˻4?IF?�?��>˙�>B!���S >��>��n?G�x?5�o? ��=b�>�>���>��$=���>%c�>k?��Q?xou?HzJ?��>��F;rS �Y��P�p�~Ѭ<)��<7�;�Y^=>���J4��|#��s�=Q�	�����Nk�[�������Y���<��>1t>�k����K>>羾����
l>�A0����FO���(��&>��E>�P�>�@�><J�F`=+ٹ>NQ�>��$�?�|?�4?#)y��Y���پz8��|�>��;?S��=}\t������p��=�g?
Y?��o��u���L\?�\Q?�Q��-U��pǾ��L�����FB?̭ ?H�=:��>�y?�~?&?U:��;������^J��˒�:��>jr�=Ht��CV�p=m>=iE?���>r|N=���=]�y�BFP��Kd���?��?}��?��?�{>Z`���޿�5��E���_�\?���>�)��d*!?�(~Ծ�v���v����侟����f��� ��lH��4�,��d��2�۽�ӵ=0z?s?3�s?N�\?z
�b��^���|���V��K����WB���D�d9C�'Sm�������ݨ���=JA���X[�\�?��$?���Y��>�y��[�������]��=����З���!=��4�h�t����<_O=�b4�Q��X4?�1�>y�><�,?�h��k�w�F��(&�^F����L>UB�>b1�>�5?u��=ƞc��A��n�=eH��C���/v>�oc?�K?�n?{��&1��y��˖!�qk0�Qz��ßB>�X>@��>r�W�)��1&��<>�+�r�V���}����	���= �2?�5�>��>@J�?� ?	�	�f��"�x���1����<v�>�i?5I�>�߆>��Ͻ� �o��>Dcl?e��>�О>c�����_z���Խ�0�>��>��>�s>#�0�0X[�>h���ލ��9�1�=[ i?餄��a��K�>��R?�/�;,<��>M_��!�o0�-���>��?�?�=ȇ:>�wž��	�-Ez��|��f�B?s�
?�m־��E�ySz���$?��$>�2>;�r?`*'?��꽹8,>�o9?瓌?�Si?�L?>��>+������0���XG���d��X2>~�=�m�=/]�>a�?�i���W�0����=�q=>P�D�5��!�<��n<i��r��3�S>��ڿT[�������lM�7���UF����U��о��,�$��@&������j����!�k���wj�+����u�s(�?�7�?��)l���ۜ���k�G{���>볤����B�̾��n�9���~�W+���.��j�=�d���h��'?����,�ǿ����9ܾ7# ?�B ?̣y?���"�֎8�ѫ >g	�<�0��
�����K�οh���*�^?���>�
��'�����><��>4�X>'Fq>����枾���<z�?�-?���>�r��ɿ����I��<���?{�@�A?�I'������B=�>�@
?��B>	77����2����\�>~ �?���?�nO=��W������b?eߴ;`qD����b�=�?�=�.=��
�:�D>�><���7����.�,>��>��$��I�J&]��<�d>8Wѽ���5Մ?+{\��f���/��T��U>��T?�*�>T:�=��,?X7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=v6�	���{���&V�}��=Z��>b�>,������O��I��W��=�S�`�ֿI)����`�=�n�=zV=�ݾÁ�w].��6q�4Ծ�p�+X�w2�/�>�?
��>��>,b?�Pu?<��>&aa>6��'����ھ�R(ɾl���@��nC�;iZ�l�u?��#��4�6>�AľS�<��B�=k6R������ �c�b�G�F���.?LD%>��ɾ��M��D=<�ɾ������u;��E̾/�1��-n�+ȟ?�A?+텿бV�_���������eDW?���,x�q�����=C��>3="ڝ> Ǥ=��
D3��S��';?�?G���Q�H�5�>����#�w>*�?&J!??�,�G>�w?��žѵI��>,��<��/>�>!}�>d��&���; ?�{?(lJ����Da�>J�ּ�$�	ts�G��>�F-��2Խ�IU>'ϋ>�Lپ�P�=�~�=\�<=�-W?���>@�)�� ��y�� ����?=�?x?�i?u�>�k?��B?��<*��I�S�^�
��t=�W?
+i?0X>������Ͼ#�����5?��e?[O>iOh�C���.�R���?)}n?K?����0Y}������,�6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������h��=�ە��Z�?]�?ք��	9g<.���l�tl��Hk�<Լ�=U��E"���C�7�.�ƾ/�
��������ҧ�>Z@�M�%)�>xI8�n6�nSϿ���?[о�Qq���?U��>��ȽL���b�j�.Pu�+�G���H����R��>�Ȉ>ˍu�F���YYP�X7�k(�۹>�H+>���>ā#��s�9
�p-R=�W�>���>��Q>�/������ߛ�?J�W���%���]�;��Z�?�8T?f�??�A/?�۱>" �����u�>���?��?��z?|�@>�¾	�v�	�j?�Υ�ag_��w5��B��b>��3??��>X�,��D�=�t>!��>g+>�".�o�ÿᴿL����?���?n���]�>3ߜ?��+?84�G���qF��)�(� �<y�=?JI>I����� �h�:�p&����?W�1?_-���d�_?�a�\�p���-�b�ƽ�>��0��Y\���{r�Pe�0����y���?3]�?m�?!��� #�1%?i�>���L"Ǿ+�<���>j:�>WN>f_���u>���>�:��=	>��?�|�?h?,��������T>��}?	��>�o�?���=;��>S�=����G�z<��&>r`�=���Q4?�%P?��>Q��=��+��01�+�B�L�M�� ���F��t>#�d?��K?�EQ>(1���52�k)�ۅ��<����^W�L/*�hb�{�'>A8>�1>��G�L�Ҿ��?Hp�8�ؿ�i��p'��54?.��>�?����t�:���;_?Hz�>�6��+���%���B�^��?�G�?=�?��׾�R̼�>8�>�I�>M�Խ����S�����7>1�B?G��D��p�o�~�>���?	�@�ծ?ii��	?���P��Ta~����7�a��=��7?�0��z>���>��=�nv�޻��W�s����>�B�?�{�?��>"�l?��o�O�B�q�1=3M�>Μk?�s?�Ro���t�B>��? ������L��f?�
@u@`�^?*�hֿ����`N��R������=���=܆2>7�ٽ_�=��7=��8��=�����=n�>��d>&q>[(O>�a;> �)>���M�!�r��Z���Q�C�������Z�C��Xv�Vz��3�������?���3ý�x���Q��1&��>`���=0	E?�k?�l{?��>�>���t>=N��%ѽ�oz������Z=>$*"?G�*?X�?��=�E��eiZ�Ni��jg���6g��8�>1V$>���>�}�>$��>�V	=M��=ʅ.>�>m��=�?�=����^�=��>_�>�%?顡>�o<>��>5˴�3���h��w�T�̽���?S����J�.&��R	���l���C�=�\.?��>����6пE���:H?���*��b+���>��0?�cW?�e>C���QUT��Z>?��K�j�8�>�h��o8l�'p)���P>�P?�h>�Uu>�3�L{8��P��ݯ���z>�"6?羵�7��fu�u�G���۾[�N>��>�0�������i�~���j���=�:?�??p��������v��^����R>��Z>�=��=�wM>"�d�׿ǽHH��.1=���=�?^>ˮ�>�r�=�O>���>�ɡ���9����>!�M>RmL=_S?h�$?Rg������!1���ݽNQ>P�>�yм��>�ŀ�Vu$>K7?��I>��߽�ڦ���?�t���]�!>9e�?������->��,�@�<I��=C��=��:���O��~?���(䈿��e���lD?Q+?^ �=8�F<��"�E ���H��G�?r�@m�?��	�ߢV�?�?�@�?��I��=}�>׫>�ξ�L��?��Ž7Ǣ�ɔ	�.)#�iS�?��?��/�Zʋ�<l�~6>�^%?��Ӿ$g�>Rp�dY�����r�u�X#=���>|;H?�O����O�Q	>��u
?�?�_����X�ȿS}v�N��>!�?���?u�m��B���@���>0��?dY?0ci>�a۾�UZ����>�@?
R?��>�4��{'���?۶?���?c�B>̐�?�Gf?j��>�����T4�?��:���BH==,�!�>v��=V�˾�RI����E����l�U���hu>��?==��>U��u㻾jD�='�����*��9�>�È>�Xf>���>�� ?×�>�*�>�_=�=��Sq�ѳ���*S?u�u?�5���q�����5>��?��L?!��>TZ�^��>f��?���?��j?ڳ�>�������F]���C��X�=*C��J�>�">�U���>a7��M�>����x�>ԍ�=g�"ß�즔��� >�Ҵ>�[�>fPa>]�?A'(?��=@�%>��/��o��փG�߶?�i�>2<?�L?E�>t�ƾ��4���iw��W�n�;�?+�|?��5?2`�>>ɠ�8����:;;��=�O.���>?_7t?Fg�=��>%@�?��]?]�4?�Ǳ>�>>C����~��<=!�1?��|�y�D�n�F�DsM�S3?�8 ?M��=�`F��
�=t�>�߾kd� �?�M?�E0?�5���Y���Խ�n�R�m���J;��e�i��=���>��?>5M�1�Ѽ��Љ޼�F�������.��1*��>1ٽ-��t>/=,?��G�{ۃ���=��r�?xD���>�IL>����^?gl=�	�{�����x��	U�� �?���?Yk�?S��A�h��$=?�?S	?i"�>�J���}޾4���Pw�~x��w�M�>���>t�l���J���ٙ���F��c�Ž��1�>���>��?;h?�>��>��-�33����I�C�D�ٜ+�C�;��\���
��g�q�F�=��ľk�����>t6C<���>��>s� >%��>2��>-(>��T>�v=�Ne>Kt><�[>�>�7�>z�G=v�AR?�f����'�_<��c��!�A?�d?D��>�f�:��� ����?�)�?�M�?lv>�zh�*+��R?���>Y����	?i�>=*����c�<oW��·��~��:���,�>0�׽>:���L��Cf�0.
?Y�? z�̾�[׽����?¼nE�?��#?��.��Z��Lv�|�/���D��#�ra���������{�h��푿�x��Z���
l�Z��<�F?C��?�����'�Ǿ|_����,����>+c�>"�>\��>�݂>H�
���#�n�hK7�hޮ��"?(��?X�W>�o5?K�_?�@g?�
Q?�B>+'�>����x�>bV�{E�>��>̩/?M�	?�!?�%?8�I?�>y>7k=������Ծ���>O8?M]?(+�>���>��y�!H=n����=$jN��$���L�=�-�=S����:��P�=�J>��"?�����6��&���X>�9N?�� ?bDt>���JK����=�z�>���>�q>/��m�V��*���>�!�? zW����<%�W>�>(�=W����d=I����>㪛��\X�q]m=���=�T=��彩�6��tH=���<i�<�t�>8�?���>�C�>�@��1� �]���e�=�Y>!S>�>�Eپ�}���$��r�g��]y>�w�?�z�?�f=��=��=}���U�����D������<�?DJ#?*XT?^��?~�=?^j#?�>+�dM���^�������?�@,?d֑>����=˾򚨿��2�S�?�v?�a�M9���(��.¾v6ؽ�>Va/�Ԯ}�P��^�C��/�����d6���h�?���?1<���6�|��r������T�B?���>R�>ރ�>�`)�C�g�*
���<>QI�>O�Q?&�>��O?�7{?W�[?�GT>Ę8�Y*���ϙ�F.3�&�!>�@?���?��?�y?�m�>
�>N�)�� �Ub����j�Qӂ�ZKW=�Z>z��>�*�>��>7��=A Ƚ拰�s�>�_f�=rb>��>8��>� �>�w>�ͮ<��G?���>Vb�����o������f�<��u?G��?z�+?��= w�f�E��-���V�>�m�?���?7**?ӻS�I��=�G׼L綾;�q���>չ>E�>)��=�>F=UZ>&�>���>DK�M_�n8�@M���?�F?{ڻ=5��������e ��5u�T�E����qه��);��E�Y�;�+�*e����+������{����8��}΢��پF��>`B��d>E�>76O=�IP=���m�>��c>�)�<@��C��>6]��=�<��=Љ�=�2v=���l���o?�:[?�n7?��A? :]>�f>�=�zNF>0θ��%�>b�>h]�~#��_�%��k��i6��fľ�޾:T��<-��Ĉ�=�)@���'>��">���=s�=ȑ>� �=S�=�����D="��=e��=wF�=R>nP4>)>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>28>�8>D�R�C�1��\���b��Z�x!?/;���˾
W�>�+�=��޾��žAf/=��6>��`=���JL\��/�=�m{�؍:=/(n=���>O�C>���=dٯ��_�=�gI=��=��O>�*����6�|�)��3=���=Flb>��%>��>#�?l0?�[d?�=�>>n�v�ξ�3��p/�>��=]4�>s��=�B>�~�>@�7?��D?��K?V~�>J��=��>��>�,���m��X往ǧ�WI�<s��?�̆?k̸>?�S<x�A�k���Y>�WŽp?P1?k?Vݞ>F���B�$��.�� ���T=ͪ�=z��(爽�u@�ؕ��5�Q��=���>���>C��>8�>'m�>�Qb>��>�1)>r�:=֓�<YHͼW�=�0�_�@=�L�Ā�;4��������8����E�ּ���<"�.=1B=�z#=j��=[�>�?�<7d�>�*>0��$>ӵ���;���O��2���I@��0T�=����1��!���x�=
J>�l�<�]��8�>G>d�R>cb�?6�`?�[t>�?2��$�J@����
�����y��D���p���L�9�X���4�u��>��>^a�>l8�>�ۙ>����?�`Z@>oS������[>��b��p=����ςW�6c������*^�|��;�wU?���9,���<�?�B?�2}?�Z�>u���?w��hV=�A��t<]k4�L-D������>��?���>���x�:��yƾ�9���9�>�S@��Q��A����2�l�=����D�>����Q˾FR2�aF��N!����Q�ڍ����>{#S?�خ?���ˊ�x5_��{	�M����?�i?�|�>	?�g?e���M���z����;�V?���?_��?�JP>��=�����j�>V�?�ɖ?���?F t?�B���>���K&>E߫����=�8�=�
�=��>��?�?,�?4y���	���=�߾4N>�$�<�/�=���>/o�>�vb>m_�=�Μ=Ga�=lg`>�>�	�>��p>-p�>Es�>����p�rj'?�=���>��5?g�}>  �=�%��H�L;��Ž} ^�h�X���������:;��;��#�<nU�݆�>{�ÿ�R�?zb>I��(?| �wk<�^>�uR>6�.��>�QI>�2u>�'�>�t�>�UC>�E�>!{>r�Ӿ
��="Z��A��K�E��6]��r侙{�>3����,�������.B��4��{��o�
T��6�%�F4=�h�?S�<�\x�4�3����w��>��>N�7?����l���l>���>"�`>9��A���ļ��}���ڕ?���?L+c>G�>�W?&�?	�1��53��IZ�&�u�K%A��e�}�`�ԍ�}����
��Q����_?y?,AA?7��<"�y>���?��%����/6�>[/�P;��S;=��>�Q��ˋa��Ӿ�þ2���E>��o?U�?j?��V��%��'��=J ]?��\?Hb�?�?�F?SL���c
?���;�	?���>�?a��>�?]�>z�>��>��!��_齳�޾��X�|X���q�=�� >'�!<�ۇ�vF	=�7�=7{�<�n����eE�X:��ƩS�,2>�&2>���>F�\?���>`��>M�7?���5������p-?/=?#��V���a���z}�D>��j?��?�Y?o�_>�8D�J�C��<>�ω>py(>(1Z>�"�>F��=�@�掆=�>u�>�1�=�J�-������b��F��<z�>f��>��>U�<���C>`پ��žBT�=@�q�գX�.���M&��=��ٽ���>n6?v� ?�+=��0���?}�̾?J�%?�_?���?�-���`��PK�`�]�����n/D>���)�d���6���'U�����h��>���xǠ�pb>����p޾�sn��I�U��n�M=�d�~U=/�u�վ �~�+%�=[1
>ٹ���� ����Ȫ�>J?W"k=򍥾[�U��d����>|�>sĮ>\;���v��k@�`�����=��>^2;>���T��M�G�-�NI~>�A?^�6?��n?T�j�	7g�6*&� �ᾌ�d��^C���?�G�>e�
?^S�=�>|皾���\�x�&���>���>P�*��H�Hə�x��.A4��ij>�=?+M�>�?y�W?�%?�:k?�E(?U�?��>.�н��-?�?�L�X�{�Oؽ���+K��I�>�@G?�ؚ<�P�>�D?��H?�#?�L?]?
��>_����G�ed�>���>�+T����G8l>�cC?Ҋ>��+?	g`?��>��5��th��~�=��>�>b�.?}�\?CE�>��i,�>����P��=�}�>8Xw?���?��v?�5>��>P�>���>��J<z�>���>�$ ?biM?���?lGc?��?�?=5ս�׫�F	�3�%�=z1<�}�='�˽(GK�+_3��r�<	ˁ<b�7��ר<��K�%��D;�9H�@=Rj�>J@t>�T��3�4>�hž���h�E>����{��F��J�9��1�=7��>ö?w��>�^#���=�P�>�3�>c��+�'?L�?�3?��>;��a���پ�}K�Zg�>NA?0��=��k��䓿�&u��t=�6m?�']?�V�����X�[?!Jb?7%���S`���s�T�D�]�%VC?��?��=�t�>jt�?�on?s�?���'/I�㬄�E�?��6����O>uj>�+��4[���>�o%?�n>�[�=��b>�þ3&b��Q��J?y��?��?�/�?B�>�ʌ�E�E�������c?�]�>R����'?v�:俾΁�bw��5���n̾�F������$���B������ơ�=/?��|?��p?�%J?����x��DL��Zl��&H����#�͜8��j-�|83�h�g����,����
��E�B=���/4C����?N&%?R4:��.�>w���8뾁�Ⱦ�s*>Li���p.���\=*�Ƚ0�$=7�f=2y��8$��!����?$1�>���>8�6?�b�P�D�l�,�ZI3����T3>��>�H�>]��>��o;��4�����w˾�����н�
t>�b??�J?��m?������0�#�������������6>dB	>�Ԉ>U�[��!��&�?�<���o�1=��������T�f=� 1?r��>걟>"�?�w?��	�����O�y�Q�4����:
8�>�Ig?�.�>�h�>��ݽ���t�>�bk?�b�>���>����� ��{�lĽ�"�>>�>���>��o>D6&��y[��������d�7� �=��f?�u��f�`�-�>"P?���;�<�G�>�˄�/�!��|��K�-�<��=��?�r�=�9>��ž��` {�Ln���gV?�*4?cJ�w]�����*�>\��>x٣�?��?�.?6�����>��?S�?-?��n?�'D?�Ӿ^�����]�a�M��=�f�>����4�۠�>B&�ӤI�u5��1?9>ըl>W��j?1<O�=__`=\�O�]��1�>,Iۿ,yK��Y׾����A��	��i���������
��=��Nv��3nz��/�d@)��T��Te�܋�l���?��?!���_B��0 �������N�>6�p���|�;ȫ�=���씾��߾6���ԛ!���O��hh�B"e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >XC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾t1�<��?7�-?��>Ǝr�1�ɿc���t¤<���?0�@�"B?4�#���ﾹ��<��>�D?�+>��/�Wq������>���?胋?��=�XU�{���^.f?n�u9\�J�YT:"��=�đ=�(=y�mv?>���>U��6|:��⽏�0>�}�>����FT��KQ�Y%=@Of>߂�S0��5Մ?*{\��f���/��T�� U>��T?�*�>R:�=��,?U7H�_}Ͽ�\��*a?�0�?���?$�(?:ۿ��ؚ>��ܾ��M?aD6?���>�d&��t���=O6�����{���&V�s��=[��>Y�>��,������O��I��a��=����ƿyA"���\�=�N<s�\���꽸����ik�`��|�u�S�����?=Y�=�6R>���>�V>�#Y>OV?�+l?m��>�v>,9��r����˾:��b��e%�����*�������i�޾w�� u�o��g�ɾf�<�܁�=�lR��v��MT ��yb��qF�|�.?�^&>�ʾ]M�m5<<�Ⱦ�v���w�����|Y˾g�1���m����?�A?�����%W���`�Sz���CW?�#����:¬���=8K���F=�5�>t��=\�ྈ3���S���8?nk?[���6Q��<�+y��:H��+?Z� ?ˑ�=K��>4�P?4}l��+�=(3�>���>C1�>|��>I�=QԾ��K�/�!?7P|?��!��v��0��>�מּ�Ǧ���B�9;>�1��x�轆5�� O���ھpX����=�Ss>�$W?V��>�)��m[���7�'�<=��x?#�?�*�>`qk?��B?�z�<�c���S�`!��`w=��W?<%i?k�>J����оFt����5?��e?O>Awh�=���.��X�d?��n?O?���qx}�q������m6?��v?s^�xs�����L�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?z�;<��U��=�;?l\�> �O��>ƾ�z������0�q=�"�>���ev����R,�f�8?ݠ�?���>�������2�=B╾[�?��?*����h<%���l��j�����<���=���ռ"���1�7�{�ƾ��
�w���������>BY@�k轷$�>Vm8�<<��LϿ���Egо�>q���?>fsȽ���^�j�}Zu���G���H��������>�L>����̠����w�f:��e��_�>��y��@�>�
H�kH��:=��^\�;�f�>U8�>���>ڋ��	���"�?a%��Ϳ����>��W?�ʙ?w�?�x!?W�"=WEo�IMk��x<��J?��q?w�Y?(
���4_����j?_���T`�&�4�GHE�2U>"#3?�C�>�-��|=�>։�>�g>j#/�q�Ŀcٶ�����-��?���?wo����>L��?<s+?�i��7���Z��>�*���+��<A?i2>�����!��/=�/ђ���
?~0?{�4.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?���>3w?�ʊ>�?���<)���=���>��>���'��>x�8?���>z��=#
K�ׯ��1�ɒ4�B�辀�4�3�>t�?Z�B?��{>}
��d��_�;�P���;�c4,=�XI��~�	����>pp7>*��=|�[�kҾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�b��=��7?�0� �z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?�Qo���i�B>��?"������L��f?�
@u@a�^?*i=��<y��򣹾��\��l>л>�A+>������ ���Ӽ��=ccp<7��<��z>"��>W�{>z��=�;>�a>[zz�4#��Ƣ�mA���?���׾q.=�@��y8���U�-���-��3�;��m��-=F��Q�����#6����=&�T?�iU?��q?���>'����">{���=*r-���=�{�>L�/? 9J?k�(?�Č=�����b��W��^ॾ���{��>{&M>
F�>\��>,�>	w��C>��8>:�>X��=��<��»�=k
G>Y�>���>⩷>�A<>�>�δ�1��_�h�c
w��̽� �?�����J�.2���:������\�=�a.?6w>���>пI���1H?w��� *���+�P�>��0?SeW?��>����T�0>>�����j��^>H% ��wl���)��Q>0l?͈f>�]u>`�3��98���P��m����|>�6?�����9�]�u�>�H��#ݾq]L>rǾ>Y�G�@n�Z喿f�~���h�}=�:?�Q?Z ��ٰ�ct�t���sR>��\>D�=0�=��M>�a�M7Ľ�F��(.=�2�=�_>��?��6>�y>�6�>6���}��{+�>R��>��'>�?�?�&Ѽu|�*�V�[cc�F>�r�>ax�>��>�Q�e`�=��?�>duC�"V��%���J�ݝc>5�g����ᓼ�&=Eԉ�Q�]>�h�=����I�n�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿrd�>1i��W��u��d�u�t#=.��>�:H?gX����O�u�=�p
??#c�������ȿ�zv����>��?O��?��m��@��C@����>��?RbY?�li>�X۾*7Z����>	�@?�R?�"�>8�A�'���?�ܶ?���?8I>ċ�?��s?�q�>�0x��[/�m1������y=]1V;�T�>�L>
����dF�{ד�Ig��w�j�����a>ٗ$=*�>�<�<1���'�=R��D����f�y��>�-q>b�I>�T�>n� ?N`�>o��>p=e��n߀�׸���]T?A�?C�w�y��*=b��<�Ⱥ��?�3?��H>w.Ӿ���>��u?�z�?�(Q?)��>}	������DV������I���>g?�n�>V:I�%
O>쨾��M���2>��>��Z=�D� dY���)=��c>:�>̊�>��/>��?�G3?�V>w>��Y����;�?����>j0�>�|:?��r?�Z�>��߾�-������ش��cN�X�?�[�?79/?�X�>M֏��J��$+�>H�W>\�|�DD?3�?��T>���>��?d�U?>�l?���>`�)>�膾%�����缮� ?h��V�A�(�%����Z�?{�?���>s����{ݽf��5��Ȟ����?K�Z?�q$?�����`��N���4�<p�׻��&�Ҵ;�<����>��#>�7��P޽=��>$�=_e��1�<��<�F�=!Җ>�Q�=<��D��/=,?��G�gۃ���=O�r�IxD��>�IL>���x�^?�k=���{�����x��	U�� �?��?Gk�?.��7�h��$=?�?o	?�"�>�J��~޾͔�,Pw��~x��w���>��>\�l�-�G�������uF���Ž$��|�>{m�> .?�?5#ּT��>�����⾼�-���@�ǦJ�bWᾅ#���1����w�XI��D�=����K#��Z!>�X���=���>1�>��>�\U>�@=VLx>)��=�ab>2G>�H>��*>̏>�`-=Z��GR?�����'����󮰾�"B?%qd?9�>��h��������x?���?9m�?�v>|h��%+��l?�9�>��n
?�O:=,E��?�<�W���������[�0��>�ֽ�:�0
M��cf��j
?B*?�g����̾�A׽"Q־`�;��?��?B�S��K��$K��D2��wP�!����J�-�&h&������ ���P��X���8�׾�� >9?k2�?̃���ʾ�ʾ
ŕ�*�0�7�>^2V>Z��>��>�NP>��侪��F�y��lW�fV�X?�(�?�D�>�,F?��G?��U?u5@?xSb>O��>,[��`X�>����o�>D��>Na1?\�%?2�'?p?�#$?0�\>����e����о5?{�?qi?sE?�+�>j�����н�F��������-��ED=j�=���x,S�{�2=�D>��?�Z��/�L��.�_>��'?�'�>���>�������Tr�\��>�A
?�>��	��o�NG��{�>��~?�c���9=h>�h�=}bt��K����=kI�`�U=i�;�����<� �=��=�X<�HO�i��;��;�a;Ht�>Y�?P��>�M�>>���� �������=Y>�R>j�>`Gپ�x��� ��v�g�Ey>!t�?�w�?��f=q�=إ�=z���T�����V���KO�<u�?�B#?�UT?���?I�=?�g#?j�>_$��I���Z���
���?�-?�ӓ>cE���ƾ����f5��V?F�>�j^���[G��P��4��W\">�q&�4Ut��K��[�C��	<M���3�����?k�?x3)��7�rD⾡ѓ�����״<?�X�>�I�>�P�>s�/�|�c�Ö�*>W�>��S?�&�>,�O?W:{?�[?�mT>>�8��.���ϙ�n�1���!>�@?&��?1�?&y?^l�>��>��)���P_��|����ۂ�JW=�Z>���>^�>ݩ>���=�Ƚ�T����>��X�=��b>���>��>a�>�qw>ݮ<��G?��>�������o���������>��xu?���?��+?z�=�P��E�����Z�>^c�?7 �?��)?�T��B�=��Լp���0�q�X�>�ع>C�>��=�D=�s>}��>���>�.��#�^W8�=+L�%�?��E?T��=��ȿ�$��nݼ���.">�*�>�&L�F[ξ5O5������_�9�۾i���[�({�=�\���/��C��F0��>��6>I��>X [=P����@$��=��U>��\>�ټ%ҽPs��.���3�F�y�nY!=s$=(9>ù�<E���r�r?�`?��<?D?@{S>|�">$�O��>FC�9?!�>��˽s>��a�+��;������Vʾ"-;�CR����v>����{O>K{>%^�=;4=1re=at=�y�=�b��ԻcO0=�*�=�o�=:�>�A/>-�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��3>+?>3FR���/�сT�Ajb��%N�F� ?�s8���Ͼt|>��=qܾ��ɾ%D=�/>P�1=���h8X�B�=F�\�cw=�vW=��>�u>>���=,n��S��=:x=)�>1OR>���;����缁vt=��=ܖV> �)>v��>��?�I0?�Pd?�_�>�-n�[�ξ7����e�>���=�.�>�c�=�rB>"/�>|�7?��D?տK?�Y�>O��=� �>C��>w�,���m��/�`w���5�<���?Ɔ?�>��J<�'A��C�c)>���ŽA\?G�1?�c?Ё�>W/�����N%�8�-�V[�� M�;�#=~�w���z��'�6�"r�B�=S��>1�>�D�>�"s>�6>X�L>���>��>8e�<"��=+�ػ���<�o��w�="0��/W�<�ʼ:YT�x��j7�=üT�;�k�;,��<�<�>]'�>�}�=���>��6>��ž���=;;w�fT��'�8\5Ծ^�"���8��2i���(��΀�ֶ>�Tb>F�<V����V�>��>�L>���?�pj?�#�>�6�������㨿���]��Fk;����ܔ����<��(T���:��/��.l�>s�>�g�>K)m> '+���>��jk=V��x54�F��>0����i�ԥ�J�p�.ڤ�3՟�,[h�!~�(D?�7��a��=ϭ|?�@I?���?��>���m�ؾUa.>4��|��<cy��t����?|�%?���>�3쾥�C��T̾�ε�-?�>F�)�}�n��k��o]&��;=Om�Tt�>H�]��b��b�9��؊��朿��p��@����? g?���?xa�Wm��a��*�ӼS��>�h?�#�>$*0?�� ?��Խq�0!�囉��=H?3�?��?��F>�`�=V����?y%?tq�?��?N�s?d(��O�>���{IY>�s*���U=]�|=->���=�2%?��(?g�?$�V����=澦�۾��R�g8>�\�=���>a'(>��>=��=�w=�x�=b >r-�>Tn>���>4�>A�>�i������V(?qH�=JЎ>c*1?�̂>UgX=؎����<�-?�fA���-��`����߽Z��<�P^��R=J�ɼ}V�>ǿ+��?�S>:�e�?����'�.XQ>tU>�P߽�[�>'C>6�x>a˭>�_�>`b><�>ʋ'>LSӾ9j>����Y!�T6C�SR�\�Ѿ�vz>�����!&�&�������XI�񅵾wm��j��/��[*=��<�F�? �����k���)����q?>M�>�6?錾�ӈ��>&��>�>F>�����$̍�G_��?F��?�;c>�>��W?B�?�`1��3�jZ��u�k#A�Oe���`��ߍ�b���ՙ
�w��Ⱥ_?��x?�vA?�T�<�.z>6��?��%�>Տ�z0�>�/��;���<=�!�>�����`�K�ӾK�þ=V�f4F>�o?�$�?�[?KV�'�m�!'>۴:?W�1?NNt?+�1?
�;?�����$?�e3>KF?p?<L5?�.?��
?b2>
�=2���q�'=H6�������ѽiwʽ���n�3=N{=i���$�
<�=��<#��l�ټ�;�����<�:="�=~�=��>HW]?@:�>X�>�7?����7�;����/?4=����,抾������)� >Ԁj?���?Z?�ad>��A��{B��)><��>��$>��[>:�>��뽯�E��>�=�&>�>+��=�~N������	��.��/��<UQ>;�??V�>好@El>Px�����>˪m����5�H��!־����tv����>��@?o�?�}Q<X�;��U=MKb���>�EH??�w?ϑ?".�=K�׾�H�F������6�<"�B�=7������ُ��=C��jݼ�R�>��2��4��Vl>y�
���BBn��J�V�h^|='G�x��=J0�A"оf�d�2��=�Q>ꧽ�������d����H?�l=h£�(P�!�� �>���>Q�>��K�~�e�ܓ>��n��Z��=��>�5<>4��
��;�E�@��kl{>nGB?�bO?قk?Z̓���n��N+����,^^�~μ��>��>.\?�i>�??�xվ�� ��U�(�/�۽�>���>�~0��qU��@k��%��S1�U�z>R�,?��>�1
??�9?��?zmr?�y*?*�
?	��>���e׼�
R'?Վ�?-[�;J \��j�F�5��uO���>�#?�h�צO>�3?X�2?.�1?�J?0G?i�>�K�=L��ܩ>��>�"N�P+���dZ>�QQ?�/�>TTC?tvt?�>�)9��z��=�U<BKS>��+>`�4?�e2?α�>�\>2�>K����i1�i��>J��?��?�І?�j�>��?.�۽��?���=�?1>8�=R�?Aކ?v�j?xA�?�9?x�=p�Z����=�m�=�����;c�8�Y\�=Zm[=���=�K>�j>��=>	͋��H->��A�?����Hs��-J=�H�>L=�>>�&�i�>/7��5��s�@>Π%;�^^�H<������Ĝ�<�R>rq?�<>�di�(>���>��>c����#?/�>:H?�.&>��]�'��]���6�>/l,?>p����{��N��	j�T����\?(�p?��a�&�!��L?�]?Jq�k�X��ھ��;O6#�(MN?�!�>�7=C�G>�1q?֜p?���>M��;�R�����q�]� m��>܈>7��>tR!��.b�>
�<?��e>|�=\��>!+�<�r��Ύ��:I?*h�?
��?�Q�?��?Gփ�Q�翧�?���S?k*�>+���T&?�����ϾD��������A徭\ ��ٴ�n���- s�Γy��l���� �`�>>��?�T�?Pt�?�bP?`��s��Vn���z�5CZ��j�X�"�;�?��#��zT�����	�87
�l|ھ�lؼ z��dQA��m�?��'?�V/��~�>������C;%�A>@젾�7�0��=����07=��H=�k�f�/��Ӭ��I ?'�>�>�5<?\\�`\?� /2�~�7������4>���>_k�>-o�>��庛A4�q�ܾɾ����~ؽ�w>��b?1�K?#n?���1�Y���e ���8�����6>>�g
>;�>�tX�W���w&�hD=�a�q���j��H�����=�Y2?�{�>�x�>���?�?�������Dw��"0�k�7<��>�&e?*�>��>�gŽoL�D\�>3>i?�R�>D��>lĔ�M^ �?q��Z����>�6�>���>�`k>,l!��Q�ύ�IB��'�5����=~~l?�z��Epb��8�>��N?oݤ<u��<)��>P�s����;�Z�:�p��=.�?6�=((>T�ȾM����v�`��dD?'0?�Y��E�c���=�? F�>4%u=ߢw?*O?B�ξ+ֳ>���>=��?�()?�O?���>�ך�7�P���j�O2��q�6;��>��A<5n���>�*����������0>5l>����ц��U���=�@�d�=N�>GGۿ�qK���ؾX��xz�^	����ó��A�����񴾛����y�`�����pOW��e� W��%�i�*6�?�(�?�b��늉���������(���o �>`�r�E����L�����~"���ᾨi����!��/P��si�Re�N�'?�����ǿﰡ��:ܾ,! ?�A ?4�y?��7�"���8� � >�C�<P-����뾬����οE�����^?���>��/��v��>᥂>
�X>�Hq>����螾�0�<��?5�-?��>ώr�1�ɿb����¤<���?/�@�=A?�(�X�꾩R\=�n�>��	?��B>j1����7I�����>ݸ�?т�?`�C=��X�̊	��e?��<RyF�HN����=`��=5Q	=� �I�M>��> X�QCE�J�۽��1>%/�>ͺ��c��_�x�<�^\>��ͽ����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=r����ſ�5'��ʖ=�z>���	e���]��7��%|��+��S=��KmC=4�>�.><p>��>,��>��A?�e?�o?6I>x(5��D������*�>�����b?D��c��(s�w{վr����1#��-��P0�!�^��<�T��='R������� �G�b���F��.?~e%>�Nʾ��M��7<��ɾ�V���6��is����˾�1�[n��Ο?��A?!���5W������d!����W?���S@�)֬����=`ު��@=���>�5�="�73���S�)D?!?�����T����|��`2���=���>��>���=��
?�w`?����$Q<>��m>�ң>�9>>6G>oQ> ��!�D�??�`{??@e���羹H�>�a���ܾ�&�����>�i������>4��=�o��-�3��=2>w�->�W?���>�)����g�������A=�rx?Q{?H�>��j?��B?$��<���3T���
��|=P�W?��h?�8>�R���sоb茶��5?K�e?K%Q>H�g�b���.��_�v?[�n?�i?����[[}�D���n��6?R�v?�r^�Ds�������V�?�>�]�>���>��9��i�>��>?�#�MG��º���X4�JÞ?P�@~��?�<<��/��=�;?�\�>�O�<>ƾ�|�����*�q=�#�>劧��dv�U���Q,���8?���?Y��>����1�����=h◾>ث?�w�?	2��	��<��m��< ����<xjw=�{���k6�����A7�Wξ�7��6���w�(��>�@�
��v�>D�O��ݶο�Ʉ�9ؾZ�a���?���>���Bۨ��`p�v]v�g�F�m�H�z␾[��>:>gԘ�����z�UA;��T��Hf�><�Ѽ�<�>Q#T�HG���难�.G<�#�>3��>�I�>/{��ڼ�L�?����fVο�d��s��k<Y?���?7݄?ia ?���<�5u��}��ɺ��I?��t?��Z?�o��-He�g$a�!�j?k_��@U`�Ɏ4�yHE�yU>�"3?�B�>G�-�K�|=4>{��>g>�#/�k�Ŀ�ٶ�>���K��?��?�o����>q��?ws+?�i��7���[����*�C^+��<A?�2>5��� �!�I0=��Ғ���
?Y~0?�z�G.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}??H�>'A}?G�r>��?�t=�~��}!�<�Q>Kx�=Bb�O��>L�??�J�>f{�=S�R��?5��=�cC�	Ǿ�E:�\�g>Z�M?Q�D?���>�͗������/@�U�#�˘T�tND�g򴽰6���=[� >n�R>o9E�������?Mp�9�ؿ j�� p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��2a~�ӂ�� 7�4��=��7?�0��z>���>	�=�nv�л��Y�s�ֹ�>�B�?�{�?'��>�l?��o�W�B�d�1=�L�>��k?�s?3*o�B�ݲB>��?+�������K��f?�
@qu@v�^?B0ӿ9c��@��ݔ���yһ��=�^>2��d[>�$��&>�03�������=�j�>�H>�7M>���>� >�2���(�����H����|����+��Duɾ����V9����
5i���2=\���sP���
>��0�J4�=��T?@cQ?��l?7��>!���_� >�i��qb�<<1�B�F=�9�>�Z2?,qE?��&?_=b���b�b�\~�,���1����>�O>��>:*�>���>.�ܼ�\>�>:>\a{>�>{
=LM+�0�;;^:>bH�>ty�>�d�>\�<>"W>.���R3����h��w���ν
�?����&J�M*������r��>-�=�p.?��>���.п�����H?������Ԟ*�0>K�0?U+W?��>�`����W���>2	��j�� >n����cl���)��P>�g?�C�>:�>�(�KW=�S�U�{�ȾC�>��C?7��$Ľk|p�P�8�#���#�H>�H�>T�ϻ�/!�y	��2oWs����<�h7?�?C	���`��Wn1�=	��nQ?>"C�=�NK=��=�o>��� �F_�>��s&�=q�>!�
?�Q>��y>�C�> n���Ճ��O�>H��>��!>��?��2?�"μ@@��:�
�4�J���=8:�>tO> *�>#X����=$��>�$�>_G�=yo���[7�~A�`��>s������DyA�z�=���`/��u4���<�r&���&��~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ;h�>/x�jZ�������u�_�#=ߨ�> 9H?W����O�)>��v
?�?_�ᩤ���ȿb|v����>Q�?���?4�m��A���@����>��?|gY?�oi>�g۾`Z����>�@?�R?�>�9�ێ'�t�?�޶?���?��@>��?[�p?0��>�Ѯ�9e3�Y� ���'A?=#��$�o>۾>�t���F��ݑ�����<d�����Y>Ƹ=UM�>o���������=��"�#I�������#�>�$�>f�H>�2�>�U�>���>Iq�>��<�m��p�ᰎ��EM?�"�?�� ��P�� �'�� 	��I ���?���>.�?������>�q�?�y�?��E?Ì�>����������¿=c��/y<��n>r��>��G>��=��>����������=�d�>���<D�ݾY!��6f�=�%�>1��>|�c>/(>�?f  ?��>`4�>�L�BH���a��m?S�=}}?y(l?��?Kɾ�K�x��"t��>Y����5>�F�?yF+?�Ǻ>�ٕ������R=1`��������?μK?�Ć����>tW�?�\4?�JB?uM�>�6B=�����8�=��!?��b~A���&�t9��?��?cm�>Nz��z(ͽUr漼���f���|?��[?�8&?�;��oa�=�þ,��<q2�dLh��,< �_�~>��>�	��%�=�>峲=
pl��.7�Q%Z<��=WZ�>�	�=S�6�ƥ��0=,?o�G�yۃ���=��r�?xD���>�IL>����^?nl=��{�����x��*	U�� �? ��?Xk�?p��?�h��$=?�?S	?q"�>�J���}޾9�྽Pw�~x��w�R�>���>գl���I���ؙ���F��w�ŽE�eC�>&�
??V-?u�?��=�;>Ҫվp���$�'�p���Z�L���A��O��n�GaŽ[-F���I�����s|�!LT>���2A�>=1?���>B/>�#�>�r�:�H>g�W>O��=&>��#>��j>�>k$�=�k<�KR?������'�µ�²���2B?rqd?D1�>|i����S���?E��?"s�?�:v>�~h�H,+��m?�>�>*��	q
?PQ:=\&�mP�<V�����5�������>RF׽� :�HM��nf��i
?E/?' ����̾�?׽�㶾R=:'�?5�?%�.���N�3���s?���s�X�;�i`���羥���{��ύ����� ���0!�r >��@?���?�g�D�������䗿��:�%�?��=�Z�>���>���>�C��^�"�W\]���J�>���	�>�f?,{�>�DI?.�<?T�P?��J?c��>�>Cϭ�CA�>�xf; ��>O�>�9?�.?�/?!�?�?*?-b>��콩��GؾYc?��?�?��?'�?s���H˹��v���w����|��jt�%ls=���<�t㽂�f��/]=ƦU>bU?��á8�����8�j>u7?S~�>���>|���3���W�<��>��
?�:�>� ��~r��a�N�>���?J�!v=��)>���=;E��̺T�=Η¼�6�=����n;���<yu�=^��={��������:��;Y��<dh�>��?9�>mˉ>WV��� ��1����=!%Z>�O>��>��پ�X��l1���gh�̟y>O��?#+�?/ha=�q�=e��=N/�����K����!H=V�?}f"?��S?��?JT>?�#?�)>�S����'��u3��n�?{�/?�J�>��߾fģ�w2���B8�?b?�Y?H�]�����ʓ��� �_>v%�Ҫg����I;�L=����e��o
�?���?@h����*���ɾW̓��㌾�m?�8�>|M$>��
?]/�pk�A:9��]>�?DW?a~�>`�O?~l{?%\?-T>�8�����Z��5z	��>zd??���?���?b|x?���>�>�&��߾�����N �������[Z=��]>�ё>H��>�ڧ>J�=	�ɽ�����@����=��_>��>���>���>l�u>�	�<��G?���>+���/ �e���y@���:�!,u?b��?��*?��==����E����M��>LF�?���?�*?�YT�K��=lۼ�@��A\s�=u�>B��>s�>Ւ�=&[A=��>�4�>�_�>~��`!�ށ8���M���?TF?�ǽ=V�˿8D��������~��N&�/Tn��_��'�<o��=ћw��.�:`Ծ�x���=��|���螾� �	w����>K�E=tM3>�|>��@=���`9�<&y%9�c����=�ɚ�.�I=�*��s�;l罽c�|<�a<#VZ=�������~"w?'CS?�F/?�'3?��X>,%>����ߘ>R�ƽ��?��T>]J*�����xkV������ϖ��Ͼ�B����b��ǝ��s�=�����,>t�/>���=1!*<F��=-S�=ą�=������9�E�=֯=).�=��>���=�� >�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�??ti��d�>M���㎽�q�=L����=2>q��=v�2�T��>��J>���K��D����4�?��@��??�ዿТϿ6a/>�q8>>�;R���1�y^��d�Tc\���!?��;��xʾ���>䌼=8eܾҸž{ 3=��5>n�\=�S�Ԋ\���=�}���;=xDr=���>;�C>���=�����$�=�E=6��=�SN>����,?�,�z�0=h<�=`�b>�&>Q�>�?~61?�e?���>ojp��-;����`��>���=B`�>۰v=6_>>鎸>�.5?�&B?��K?G��>�M�=>�*�>��,�z#l��7޾�§��<ņ?s̆?���>-��;�I��V�!�=�׽�?7�2?V\?�/�>���ܿ�%]�Zq⾲U��@>֯&>y����
<�۸<�ٓ=�k�����[n>�?�I�>~H>�B�>;��=�B�>T8>��;�K~����>H�b>�O�X���	cŽ�	��(���@���N@6>�벽��m=�d��?uQ�o��=G�=�H�>yh>Z��>�w�=|���<,>4!��
�J��!�=���^�B��c�N}���0�yP8���H>�SU>�D��W���?<PZ>S�?>m�?��t?�>� ���־�/���Ld��R�㊭=N>��;�'�9��_���L��ӾƼ�>׏>z��>�s>�Q+�@?���~=�B߾�83� �>?����'����FSn�
���%�����f���x��D?%���u'�=�)|?0I?P�?�/�>{���4ھ/*7>ga��N��<"Y��i�靽t�?��$?v��>f��y'E�!"̾����>�;I�vP�#ԕ���0�>��V˸�!h�>ܖ����о�"3��v��E���C�)�t�`Һ>W�O?y�?�(a��k��.}O����d���D?��g?�>�(?+?�m���W�@��V�==�n?�t�?�?��
>�s�=������>��?�?uz�?AC�?�H��D�>�����/�B���)=���\Pw�6�d>�y4?�]"?-?�%��&��V���뾀t4� F�=+�k>��>Z�0>٦�><�>
�=�==�>�'?U8�>r>�?���>���=]�C'?���=���>\2?Q��>*�Z=6쩽�M�<�G�+?��+������Ὣ��<����ޞQ=�dļ���>%rǿC'�?5T>�p��?�>��~/�T>�T>+�ས��>�;F>H�|>���>)r�>�>�}�>d�(>nӾ?�>���h4!��0C��R�ʤѾMgz>�����&�C��S���@�H�쓵�wJ�&j�1��m-=�Au�<"�?=A��Æk���)���qj?r��>ݶ5?B\���I���j>��>�\�>�[������ȍ�uᾯ�?g��?]$s>��>��X?�?V��?P��S��p��s,�{�b��\�n񎿙�v�q
� $�n�N?��{?/%5?n�0��7i>��z?�["������>��+�j=�N�3����>�z������w+�t-��8�>�O� >l�i?Ï�?��?_ ��R�Q�=)>��=?C�2?��o?�-/?�:?1����$?D�(>�?[[
?h�3?*\.?z?�N&>;��=#���v#c=,ߔ��튾��ѽT�½�֭���4=��m=�۷ׂ<�6%=�<�[�?O��X:�㙼�?�<�lR=�]�=.��=]#�>g�N?��?F��>��M?a�8�l�!��Ѿ�:?�S����!���C��x^�Q?k�=?�U�?4s+?���GH�A�E����=@�>P��>6��>A��>�2׽���(����=}`>׾0=��,�}���?>þ�jg��J>�>���>�̘>5G<8�>(8��J����>%��	Nؾ��q�$C��`��PʽS�>��;??^�>�����- ���lc�� ?xF5?�YZ?OGx?Eu="�O��/Z�ֺ����gSR>��<>�km�������B���*=�c�>sN�=��v�b>A��Sb߾�n�N�I���辩[P="l���`=�<���վa}�b��=|
>�𿾨� �/��<�J?�aj=+��@V�E�����>���>ˮ>��8��t�8-@�ޅ��]�=��>�<>�F���l�c�G�%I�C#f>�1?}h?�A�?�����{�w��˹پ1���$?�מ?t��==C�>��}>|�c=(�ܻ侪dh��8����>ֹ�>�y���?��<y��+��p0��g>���>�>N�.?�"Q?w?��\?��C?�P?�u�>��#�K+ݾ_&?3t�?���=�4۽ϚU��8���F�c,�>�)?3�>�ɩ�>�b?�(?�J'?�LQ?�?��>� ���@�i��>,)�>ObW��K��'�^>YlJ?
��>gY?���?�u>><5����������s�=O� >�$3?S #?�?�ط>Ud�>oe��+>���>���?A�?��{?���>:>#?`�x>�c?:W��c�>�>?��E?��u?k��?:*{?�j�>�O=�T6���ݽ�z���~��Z��=^,L��8�>��L�%��#M.�>���3�=�3-=��=�~��̸4�;5�<�!=\h�>�+t>a�&1>�!ž4 ��):A>�:���қ�P��U�:�b��=`�>�?�s�>b�#�yX�=K�>aS�>X����'?��?�
?r��:m�b���ھ�J��Y�>��A?�t�=��l�	P����u�4.f=ښm?�e^?s�W�����X\?�JU?�
�G�Q�Ω˾�
��?��n"N?)��>ώ�=��>�_?��j?��>��~\�0K��v�W�#����w->!o>j��#u�����=��+?6��=�5�=��=h�+�vZ�m�� �@?��?21�?%�?��>�Ҁ�Q�忯R�����W?g��>�W��r?wR�:W־ᇾ^������!���Ӱ�Cך�$���u(�)ц�0v�����=�2?\Kj?��w?5�`?�m��Of�5*[���s�;6T�U�����5G���?�\SA�U�q���1s�ӎ���g=����4�B���?��'?�,�q��>����	�ϥѾ�2=>i˜�~7��+�=ű����R=�jk=�4\��]%�^*���, ?;�>��>c<?�;W�_<�e�/���6�������9>���>�H�>{�>�T1�.�1�����ž�U����߽�v>M�b?YK?,�n?�v���0��ⁿ�,!��b+�\ɩ��{@><>MT�>��X����&���=��[r�u��>ΐ���	�Oy}=�2?р>'��>tЗ?��?ۍ	��]��8u�t�1�N��<k��>YCh?��>�>q�ҽ�_ ���>�Gk?"x�>�
�>�x�u"��e}��
��6-�>��>�W�>�)0>ŗ#�u�d�1����{����8�4{�=��k?��P��W�>�N?���< +=�>����u�(3�}*��	�=j��>�F�=��>��ξ�P���k��Q[��5?�k?��э"�'�Z>�w4?~�?�8ܽ�މ?�>�>�L��{�>� Q>�:<?�<?��8?�$>�y�����;2���1�������>*�>���N�</y���Ҽ$k�
Wz=�!Z=k]�=�
����*=LCY�Y>K ���*>��пC�T�r�ܾ�~��(�����Uّ�����W�ξ����m~���T��<�^H`��hڼ�?����b����O��q�?��@r�v�o��Z��������S�>����֌<O�Ҿ��Ľ{�@	��ѿ�R�=�Bƀ���M�h,�O�'?R���۽ǿݰ���:ܾ! ?�A ?	�y?���"���8�L� >�F�<�.����뾏�����οY�����^?3��>��%/�����>\��>¡X>Iq>���f螾�$�<��?�-?���>ˏr�+�ɿ`������<���?.�@�~A?�(���쾑+S=U��>[�	?�N@>��1��"�E���l[�>0�?�Ȋ?ɫN=�W�H{��7e?�G�;��F�_�ٻ���=�`�=��=�+��LJ>t��>�w�}�A��`۽mB4>��>��%��9�X4^�OQ�<Փ\>�ֽx��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=n6����{���&V�{��=[��>b�>,������O��I��U��=U���ҿ�j��A¾�%Z>�@�_(
=��\�ǳ��潒��yC"�e�W>6_>\:�>u��>$�?��>�̩���e?YK1?!^M=��]>4�Q>lc�w�Ǿ?W���ξ˃�=�t,�?-�=�ѐ��T��u�����
��i3���پ�=�
g�=3R�א��@� ���b�7�F�(�.?�$>��ʾy�M�U2<oKʾ�몾w���?㦽�,̾-1��n��ǟ?��A?_����W����o�&*��.�W?�;�˖������=����Ϩ=��>��=���*3�8�S��2?�< ?/�Ͼ+��� >6_��>\|=�
?b�	?�� g�>�t*?2J]��l�Bxq>�v)>���>�Ū> �>�ᵾ��� ?|�R?�HG�E���w>E��O"���h<���=m������">�~B�>1��_?]��������<	�P?4��>5�+����H�~�l>~�=��[?�?�.>>� f?�\?����P�V�U�,��(o<<C?O�?�_+>F$������8���?<�?���>�^�������X���=վ��??�`#?�2?���<u$a���� s��S?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>��������=ڕ��Z�?m�?�����*g<��@l�
o��My�<Vϫ=$�+E"����7��ƾ)�
�����翼u��>;Z@gV�m)�>�D8�56��SϿ����Zо�Pq�9�?��>�Ƚӛ����j��Pu���G��H�ڤ���@�>��>�����⑾6�{��];�=��R�>����>�S��B�������2<��>�l�>���>��� �����?M���6ο��������X?'^�?�[�?_X?@<6jv�!;{�"��*7G?&}s?~Z?��#���]��89��j?T2���W`��4��:E�G�U>�*3?��>:�-��^|=?,>.��>�>%/���Ŀqն�4�����?��?�Y����>xu�?BZ+? n��5��7���*���Y��:A?��1>����s�!��#=�ȶ���
?�[0?L��2�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?·>C��?�z�=���>WP�=W����#��T>�u�=�[C�Il?K�M?�>�=�=W�6�Y�.�x=F�ޚR�Vm�ͥC�a�>r�a?�pL?Μ]>�¿���6�x��erս˨2��&�=`D�b�)��� �2>��:>jl>�D�m@Ҿ��?<p�4�ؿ�i��p'��54?0��>�?����t�����;_?8z�>�6��+���%���B�Y��?�G�?<�?��׾�S̼�>'�>�I�>��Խ����a�����7>'�B?1��D��`�o�x�>���?�@�ծ?gi��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?oQo���i�B>��?"������L��f?�
@u@a�^?*4�ӿ ����r���y����=0Y�=k�X>u�f��j�=,g`=yG�� q��(>kh�>�a�>6�>'Qx>�Kf>s�%>5�����$�h������GI����_��}@�����:�?��[�㺾U����;���\]�ȝ���3:���#��Xy��f~=�F/?;ځ?��g?s�>�׈�a�=f���A �=�b�?�>�pX>�@?X�E?�4?�D�=����K��Bx�h�����&�?\�@>��?�p�>�(>B���ў=lU9>�Ϝ>��I>G�f=��� ��=ULS>b�>?F�>{M<>��>+δ��2��]�h��w��K̽U �?�����J�a0���3��������=:a.?ߊ>��?п�����.H?����'��+���>ҿ0?wcW?��>s��"U�"@>f��Ԯj��S>�+ ��l��)��'Q>�o?``j>Zw>f�3��87�?Q��K���}>т2?�+����9�JLt�	zF��0߾�G>��>�TY�������|�|��l��[=?<?nY?�N��LF��	�t����2TI>��W>!S�<o�=DN>d�n��Խ�K��,=���=n�^>w�?	�6>��W=j�>�}���|?�#S�>+&>¼=>�;?�V#? �f�L���j���&���pt>���>�/h>m/>DP��D�=�F�>Z_j>H�U�Vͧ����;�-��2B>�r��?-i�<i����=֘���w�=�Jm=
��U�=�R�)=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>׊
��Ř�m(��4�s��C>=�վ>
RG?rw񾬺a��E9��o?%�?L��bx���ȿ�au�[|�>��?Gg�?"l��%���BA����>���?yB[?)f>w�پ��T�%�>�ZB?�O?�B�>ρ�~)�}?~?�?���?��H>�e�?@�s?���>�&z�+P/�c�L��R��=6�:�q�>�� >�����mF�ޓ�Ra��C�j�H]�
c>�b#=*�>50�xa��m�=a��wD��D�e�%b�>��p>S�K>�~�> ?Y��>��>��=����l������|xS?��?���摿BfC�̙��3�ZW?��>f-�>$�ܾ���>C|?#	�?�B?�$�>�޾Mգ��ʿÂ��ݝ�<(�2>��?R��>ey�.!x>w�ξwL�;�S=�t�>�U~=�L�n���|=��>V�>��>�܊>};?6'?���=ѻ�>9�������iF����>�1�>2z?P�P?}O?F����Z���%o���T�W��>S�s?nN#?Dh�>*N��Þ���r4���">�2��`?bP?�٫;`��>�"g?1j7?�.L?���=�0!�����Y��^E><4?���=�H���O��)F��=?V�"?��1��t����K�,��<m1���@��l�>�(?�?��=���Z�P�3��^<C.c�A�<���<��ȠO�& �=ց�A=>��B>��<3
���bS��7��l>L��>����4l ��i�-=,?K�G�qۃ��=��r�8xD���>�IL>����^?�l=��{�����x��*	U�� �?��?Mk�?��?�h��$=?#�?]	?Y"�>K���}޾��ྫPw�.~x��w�!�>���>͢l���G���Ι���F��*�Ž��c�>�r?�=A?K7>uJ��t�>�B	�?�Y���@��MJ��s�V�	��;8�,	d�!�7� 4���E-=U��>Qv��k�%o>���eJ�>f��>8�>���>*�>��{'?�����=�L�>�4b>(�=�:~>���<.�˽mTR?�����(�ٳ�qM��q F?Ue?��>�ec��r���#���?׎?H��?�j>:�h��+�ȼ?�� ?*${�In?�,=<��"�;�乾C�Ns����/����>W4߽V'8��XM�mib��<
?)�?@D��ξ����l��_�Z=��p?��#?��	��Y���l�^�:���W�hr�<!_M��,`�j<�ܙ���O���ā��|�u���U=6y9?�?��q������c�G?����>h�?M��>9�>�X>�c��-4��g�=�I��r̾n� ?R@�?�t>� 7?@_]?�S?T�;?�&O>��>X����n�>K��mR�>��>�%.?��?a�5?��?H<&?��X>�H0�J���n}۾�;?B�?��1?<�
?�e
?�캾�'+�?	�����n>s��~�%z��LH,��eĽ����]>�A>�� ?��ּ7�?�"�d@V>�[?�.?R��>`�x���}�7��=���>�7�>��>��U�r��;��o�>���?��_��a�<C��=��<$T���`w�T�5>�B7�#��< 61=*h���.U=2�����=3=a7�=�-ֽC�h��@a�{r�>��?l��>mG�>�4��� �����x�=� Y>D�R>�>(Zپ){��y%����g�1/y>�q�?Nx�?��g=�-�=���=����`������˽�]��<h�?�M#?�RT?W��?p�=?`#?�>?$��J���X��F
��G�?��*?1ʐ>nl
�0⹾�*���t.��E?���>�EW�@3���+�(��*��bv�=�)�hz�U��7F��,�<WJ�������?RF�?d����/<��x�����;���7?��>"��>���>d$���p����\?>Z��>SN?��>��O?�W{?��[?�AT>8��%���ř��4�)�!>�%@?���?��?%y?���>C�>��)�	྅`��CU�&K�Bǂ��W=dZ>c��>_'�>���>�*�=��ǽ5����>�Q�=" b>�x�>���>O��>�w>1�<��G?n��>!^��K���줾mŃ��=���u?���?Ց+?qT=ҁ���E�G��7J�>@o�?k��?�3*?y�S����=e�ּ<ⶾ��q��%�>�ڹ>W2�>�œ=�|F=`>��>h��>�)�3a��q8�yUM�9�?�F?���=�ƿ��q�Z�p�̭��);e<A����d�U���@S[�p�=�������������[� ����d������ef���{�%��>>H�=ES�=n;�=u��<��ɼ���<�,J=���<�=!So�aq<�08�u�һq�������^<rbI=v���Q\˾�"}?c�I?<�+?'pC?�Dx>�u>�2���>S�����?�U>�aO��k��L�9�?>��2���Tؾ��׾RQd��韾�'>F��5>�c4>L��=cTj<���={�q=�Y�=�b�sL=�+�=&�=.@�=�7�=�>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>4U<>�>�R��[2�w]�oiZ���S�%�?�:��Hʾ���>�9�=�m���ž6=o7>z68=C���Z�wm�=�w���;=Q�}=�=�>U�@>#~�=B��y�=M�I=��=��V>Be��h0���$���;=�s�=P�d>۪$>���>+�?	b0?RXd?�4�> n�Ͼ?���I�>F�=>F�>م=�pB>h��>j�7?>�D?��K?��>���=�>��>Ϛ,�=�m�(k�8ʧ�䢬<ז�?Ά?�Ѹ>R<f�A����f>��*Ž0v? S1?Sk?��>t�����3��u���ﴼ��=yG|��������{�����X<>��>9�?4��>5t�>"<�>B�>Ҽ�>�>!Yd=E�=t�����Pd�� s����n-�����=+�>��=�<���<)1�='$>cj�<�v�=�,�>��>1�>6�=���	$>�얾��K�"(�=E�����A�U�`�?���-��7��=>f�W>��~�ゑ��?9�V>��G>h	�?��s?I�*>��=�Ҿ����K�c�b	`�;g�=���=c�G���;��]�AZH��˾�m�>���>31�>w��>u/�{�:��i�=��	!���>�-ʾ)"��y+�rp��̡�������a��>�B�D?�:����*=��?.TT?�^�?�3�>==��Ճ�K`>�O������\�"�;��'{�*��>N?=�>�Y��%b'�	 ̾0������>M�H���O������0�z]��a����>6ߪ��aѾ,3��o��� ���B�/ur���>��O?�֮?��a�I�� [O�����h����?�Xg?�e�>�0?�O?Հ��I����~��=�n?a��?g�?�1>m,�={��$�>��?��?��?�Ju?=���>�>W?�<|_S>Yٗ�Gl>��>���=&$>--?I-?�
?/a���
�����X��d�l1=�u�=wM�>8܊>8ky>��=�}W=Q��=�b>���>�A�>�$s>5��>E�>5��e���7'?� >ׇ>1�.?�Q�>��:=Ƃ����<թx�Ko?��0-�q>ý,���K�< ���DD=Uu��4�>��ƿq#�?y_>�Z���?�� ����*R> ZL>t�����>K>�uy>�t�>�՟>O�>��>��'><̾�>G�
� �V�5�R~V��iؾ�J�>�ɤ����_x��/���IP���Ҿ�y���m��΀��2�˕ =2��?DIE�.�f�F�,���O�?���>I4??��g���4�<b�=��>�P�>,'���0��b��
𾆧�?+��?c>��>?�W?*�?2��a3�v<Z�ςu�
�@�$e�v�`��䍿D���Ǆ
�v���+�_?E�x?]A?�L�<��y>Ԓ�?!�%�������>�/��;��`;=f¦>m���m�_�M�Ӿ�yþ�����F> �o?<)�?�?y�V��Pn�G�&>��:?P�1?Qt?z�1?�V;?M
���$?(3>�v?BV?b85?T�.?�?kH2>=0�=H����2%=�u���	��Uн��ɽg��k7=&�{=���T�;�=ե<`F�vڼ��:����-�<:D9=M�=!�=��>�l]?��>���>^�7?pL��_8��Ʈ� �.?�7=����&��!���U6�c>�j?�۫?�:Z?~�c>{6B�6FC��w>�q�>7(>'�\>|ͱ>�2��E��І=�>��>w�=��P������	�_V����<0>X�?�՟>�45���>�>��o���I:�;�3|��g��s���74�a ���*�[>��?v2?��|�nm����˼+�b��Y�>R�@?�#?��?��,�)mx��8�i�"����*��=�삾�,�����������T�e~�����>�=�ᠾlSb>���ut޾'�n��J����HM=�~�>aV=��
�վ�0�?��=�!
>,����� �7��֪��0J?��j=�w���`U��p����>���>s߮>�:�t�v���@�c���J4�=���>,;>�=��%�}G�7�m>�>SQE?AW_?k�?"��\s�?�B�����mc���ȼG�?jx�>'h?�B>z��=K�������d��G���>���>h��J�G��;���0��N�$���>U9?�>��?]�R?��
?|�`?�*?HE?&'�>.������ B&?6��?��=��Խ�T�� 9�JF����>z�)?�B�ڹ�>O�?�?��&?�Q?�?��>� ��C@����>�Y�>��W��b��>�_>��J?ښ�>s=Y?�ԃ?z�=>\�5��颾�֩��U�=�>��2?6#?O�?���>��>������=��>W�b?8/�?Mp?���=#�?m2>���>}b�=��>���>��?�O?a�s?+�J?O��>��<�ܮ����Dvs�rO��T�;�0P<�U{=����q�G7���<���;���� |� �6<F�bQ���k�;tn ?$wU>+X��7�>G������g[�=�Y>iԜ�ֿ׾By��΅<;g>lw?���>z������=�Y�>>�?��"�%;1?��>@I?c�C>��z��������=�<?��==�B����w��ؐ�=	W�?��g? ���*1���f?[�?�W����Z��E^3>"���n/?��C?N)9���>o�?���?���>M���ˋ�p����c�կ\�g�N=�Û>���C�+�붸>��?.��>Ct�>K�>%0ž��~�q���d~"?�Ŋ?���?;��?I8�>�tb����M��/��K2v?��>�K����?-��9�����YU���5�k;��"����G��B���;~�L��]��k�=R�+?�?ajX?SgZ?��C�����n��d���p�Y&��!�c\r�2�d�G�8�r�c�?̯�ߪ���?����g�G-���A���?�'?P�/�P��>���ɽ�v̾DC>e���\H�r�=�ɋ��N?=N�[=h��.�h&��aO ?"��>��>��<?��[�>��w1���7������(3>ܴ�>�x�>���>��:��-�M�罝!ɾͣ����ӽa�s>�Ge?�LK?>Sm?!��j�-��̀��+!���(�V��*yG>��>.��>��Z���J &��<=���s���턒��+
��I�=�3?X�|>�c�>w�?iH?��	��Y��B3i�pI4��j�<���>J�f?���>�܉>��Ľi` �w��>�l?v��>��>'���;Z!���{�3�ʽ6&�>�>��>)�o>]�,��#\��j��<����9�s�=ǩh?U�����`��>�R?�0�:��G<}�>8�v��!����'��>S|?���=/�;>^�ž�$�'�{��7��hO)?"K?钾i�*�V2~>F$"?���>�.�>11�?�*�>�qþ�}F�!�?��^?�AJ?�SA?�I�>a�=K���:=Ƚ��&�Y�,=D��>;�Z>�m=g�=ۿ�6r\��w���D=�r�=�μ#Q����<es���K<F��<.�3>_mۿfCK�͝پh����:
�7���k���(i��ñ�Ja�����Sx����'�sV��Bc�������l����?L:�?�y���0��갚�v���U���S��>zq�_Y�����/ �$��~��Iì�	c!��O�� i�[�e�Q�'?�����ǿ񰡿�:ܾ4! ?�A ?5�y?��8�"���8�� >pC�<�,����뾬����ο@�����^?���>��/��o��>ڥ�>�X>�Hq>����螾�1�<��?6�-?��>r�0�ɿc���t¤<���?0�@}A?��(����LV==��>!�	?��?>�S1��I������T�>f<�?��?�zM=w�W�X�	��e?�v<�F���ݻ �=�;�=G=b����J>�U�>����SA��>ܽT�4>څ>b"�I����^�i��<��]>b�ս<��;Մ?3{\��f�{�/��T��T>��T?n)�>.:�=ű,?�7H�G}Ͽ��\��+a?�0�?���?��(?ۿ�ښ>�ܾ#�M?�C6?���>�d&�\�t���=�"ἄ�������&V����=��>2�>��,�V����O��=�����=����ſs%����d=���:\M��M�N���ZW�z�����s�\`�k_=]��=�>O>i�>j�Q>�5V>��V?\�i?�"�><[>�潍d���v˾E�#�+�z��5�;���gY��[����n���	��o�I�>�ǾS!=���=�6R�J���� �	�b��F���.?qw$>t�ʾ��M�Q�-<goʾz��������ߥ�E-̾��1��!n�4͟?>�A?������V�>��^[�?�����W?�N�z��묾���=���=�=�$�>���=p�⾁ 3�~S��o0?�m?h{���b���j*>$� �{=�+?:�?=�Z<�$�>�`%?e�*�T佣<[>��3>ʱ�>}�>G	>)���f۽\�?v�T?i����>8u��i�z���a=M>\>5���1w[>Dd�<? ��({R�'�����<,�`?}�>�Z(����%7=�V_)�����2i?}.3?6�?��?AkN?B�.�y���タ��h�l��UR?¥]?�|>��l>-ɾk�/�p�T?�I�?��<k�ƾ��;|�n�_"��B?�?�X ?R�V<��w��[��ZEm��VD?��v?s^�xs�����L�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?o�;<��U��=�;?l\�> �O��>ƾ�z������3�q=�"�>���ev����R,�f�8?ݠ�?���>�������m�=�����e�?��?�_��>�c<i���El������ƛ<棩=�F�%�E��"8�L$ƾ"A
��a����¼�)�>+_@꽨c�>�L8�R�OoϿ2��bjѾ��s�J?Z��>�gͽ����$�j�6�t��G�{�H����-f�>�>l���ѯ����{���;�JQ��Q�>4
���>��T�t�����fB6<1�>G@�>���>�Ӯ�>���+��?1k���<ο�������mX?�P�?�Q�?l2?5<��v��'{��n��VG?��s?Z?~Z)�$E]���5�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�^�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*��+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.��9b?M�_�{�V�� ���@�]�?�̟���L�c3�o#��t��P��J׮��е?��?@�?O}D�f���,G*?��>U�R�{*���1��#a>g= ?J�?�� =
��>�/����a�=}��?��?r�?�샿�䐿(��=gɊ?-Դ>��?F�}=��>F5�>0�z���(��&>[tJ>*���ؔ�>@U|?x��>�+=�+a�{��9.Q���t�-��۔I��dF>x]{?B�q?7�>�kƽ�4S>�s-�+e�4mV��8=-��cx��5I���>퐸=[�y>~޽��i���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*RjԿ(͔��d��v���fo�=x�>L>�� ��ɂ���=� !=��������Zk�>�Md>��h>�o>??=go�=$	���-�in���昿�0��	��8	��.�� H'�-�M�$i�@ԾfZӾ�����׼=0I=&M�P��Ǿ�����=i�^?'PQ?ĉi?0�?�ҼԐ+>���	=�� �	��=���>��3?�(<?X6?�=�3���?h�Ү������@��4��>!�p>�#�>|��>���>7�=��c>MXI>Xk�>,�=aM=����={�(>n�>�$�>��>�C<>��>Fϴ��1��j�h��
w�v̽1�?~���S�J��1���9��Ҧ���h�=Gb.?|>���?пf����2H?%���y)��+���>|�0?�cW?�>!��u�T�3:>8����j�5`>�+ �zl���)��%Q>wl?g�f>u>��3��e8�2�P��x���j|>�26?x㶾�79��u�۱H��Yݾ�>M>���>�D��j�R���'�]mi��{=�u:?��?�2��cⰾ�u�6B���TR>�9\> L=lz�=5YM>$fc���ƽt H�3�.=Ļ�=<�^>�W?^�+>髎=ߣ>vb��fEP����>��B>�,>@?�(%?Ĝ�%ܗ������-��w>�V�>��>�Z>�ZJ����=�l�>O�a>G��Ń�ٹ���?��xW>a�}� �_�3yu�y�x=I7����=��=؉ �� =�O�%=J��?F���������پ�i���g#?ɢ?�5=��*=g.9����A �ߐ�?=�@���? ��]R��(?͌�?/}��Y>t��>�	�>G�S:�r$�>Y��>,b{�ET���l���=�?��? T�� �y�6Zr���>�H6?{2��h�>�w�zZ�������u�\�#=Ԩ�>�8H?V���O�>� w
?�?_�驤���ȿg|v����>O�?���?��m�tA��@�;��>R��?DgY?�ni>�g۾]aZ�#��>ֻ@?	R?��>�9��'�8�?�޶?Ư�?aI>���?�s?�k�>�0x��Z/��6������!p=��[;�d�>�W>f���xgF��ד��h��u�j������a>��$=,�>QE�[4���9�=��I���f�<��>�,q>"�I>W�>v� ?�a�>}��>�x=�n��Jှ����
K?��?	��/���<�VK>gԸ���?k�K?E�%���TJ�>��r?��`?ӈ*?p�;>{!�ݝ��R\ſ�վ���=��o>���>[V�>�a� �>u��
p��/b>�~q>'ׅ=/��7o_�+{�=�u�>?�B�>7�>!?�#?�?f>��>f�F��Y���0F�$J�>��>�N?�[?
�?㸾l�3��h��������\�q)M>'y?�i?�Й>e�O���eº�w�)g���i�?�Hf?�M����?I7�?3�A?*�@?�vf>����x۾�IĽR��>��!?k%�m�A�M&���z?�P?\��>�2���ֽ��ּ���{���?�,\?\A&?���F)a���¾�S�<u#��qW��1�;IE�a�>��>�^����=>��=�Hm��26��g<d�=�p�>��=� 7��Z��)=,?A�G�kۃ���=F�r�bxD���>�IL>�����^?�l=��{�����x���U�� �?��?Mk�?Z���h��$=?�?	?9"�>�J��k}޾'�ྡPw��|x�lw���>���>	�l�:�E�������qF��	�Ž�/�&�>t��>_?	~ ?�O>kP�>�0��w('��_�"���^��c�s8�e�.�[�����z#�[�;¾��{� D�>���?�>��
?.$h>�{>�>��ʻ�M�>�
R>�y>?i�>��W>5>p�>��<"�нb�Y?$�����)�K�̾/�v�5?�fY?�?� :�"���0*����>�G�?�V�?s�>i/^�g!%�t�?�2?\���}
?ס6<q>0. =Vv־eBS��	K=����$ =>3Լ���P�U�����>�&?�{[=A�⾙.����9�n=N�?��(?�)���Q���o�θW�S�5���6h�Mj��Q�$� �p��쏿�^��%����(��r*=��*?j�?ь����!���&k��?��df>`�>`$�>-�>#uI>��	�s�1�h^�M'�K���hR�>[{?�L�>�XK?E�;? pO?y�M?��>���>�������>K�1< T�>���>��9?@[+?�-?��?�1)?��V>B��M����`پ��?.�?r�?*?&?����"sͽNh�Ic�R���~�H{=~��<�0�X�T���c=�~N>Wh?߲���8�l���c3j>#{7?Ƅ�>j�>�����P���e�<a��>I�
?���>����|r�)f���>���?sD���=��)>�{�=\ʆ���eB�=P㺼ܯ�=
Ճ���9�_�!<���=.�=����y���;O��;��<OB?��.?��
>��>�Ud��0�j���?�>4��=/�>Yi>k�پi����՝���q��),=���?j��?Ԥ%��Xu>>׽�뷾y���s��ۯ��S�f/?+��?�N?�ʼ?�uS?�9>7��>׮S��]��0w��W��(�?u!,?��>�����ʾ��ω3�Н?h[?�<a����;)���¾��Խб>�[/�a/~����BD�����M��4��?￝?�A�T�6��x�ٿ���[��x�C?"�>Y�>��>V�)�v�g�o%��1;>��>hR?�#�>��O?�<{?ͦ[?JhT>a�8�m1���ә�I3���!>/@?��?��?Sy?�t�>q�>ܹ)��ྞT�����o�����)W=	Z>���>)�>2�>���= Ƚ�Y��y�>��`�=��b>.��>h��>��>L�w>8K�<��G?r�>�$�����<���0����=��eu?�8�?��+?>�=�����E�������>�V�?��?-A*?O�S��m�=�Ѽ�ƶ�r����>U��>�~�>�s�=+J=e>nH�>ɇ�>���X�+�8��xQ��?a`F?�Ӻ=Q���[�D��j��(Dؾ�C���c�6�	���=�K����2>����ZG����7�y��c��A%l����������ߌ��;�>���=��>��
>�L��eґ��� ��M�=g�N>fc�= O��њ=N�=�-�l��r?�=�L >(��=X��=����Mh?���?�(?!�S?!D�>=��>Qm��@>�=��:?*x�> <�{��� )��㟾�Eo���۾� ��K��1ܾ�6~>%'<�x�=_&>K+>��=/��=��<Bgq=C�W�Y�|�"b�=[ >��>�>�3�>t�I>w?뎁��D��ԊP�6轒;9?�Q�>���=O;Ǿ{>?�g;>u?������W�5�~?��?�3�?��?�Oj����> Q���������=�򜽍�/>���=r�2��c�>�kI>9k�圿�,���6�?|�@ؑ??j����IϿ90>o(3>c>�qR��X1�6j\���a� Y��{!?�Y:�xʾ�	�>���=��ܾ"�ƾcb)=_�6>�pf=4���\��Q�=��|���7=:l=8ш>sWA>5?�=�b��*ܹ=`�M=J�=pQM>Y���'�9�q�(�g�@=�
�=4Qb>�&>3l�>&@?m�/?Εe?��>�kr���ξ8T���2�>���=Lj�>��p=p=B>`�>�&7?zsD?�M?���>C�=չ>y��>�+�@m�#N侘�����<�{�?���?�ݷ> �<�@�Ln��(>��ֽ�a?�0?�
?y�>'�Dڽ��/��p/�r�Y���[�>늾��[��ߥ<�P�����(:�=,R>M{�>��>t�=�����P�=��>�$>DG<lf="��.���솶�6�=e5�=����u����}��=Pg	�I��z�a���Ƚ�=�:K=���=B��>X<>ǭ�>���=?���B/>ʸ����L�w¿=pH��x,B�q4d��I~��/�YU6�\�B>*;X>�}��%4����?��Y>Ul?>���?/Au?�>� ���վ]Q��De�WS��˸=;�>��<��z;�ZZ`�	�M��|Ҿ���>�ߎ>��>��l>�,�#?���w=��b5�l�>S|��e���(��9q�$@������i���Һ�D?�F����=c"~?��I?o�?y��>`����ؾ�:0>'I����=O�%)q�i����?'?���>#쾉�D��H̾K���޷>�@I�.�O���Q�0�E��*ͷ�;��>������оc$3��g�������B��Lr�[��>�O?��?[:b��W��GUO����w(���q?�|g?4�>�J?�@?&��z�r���v�=�n?ʳ�?P=�?|>��=�#����>v3	?߳�?���?��s?�?��\�>���;U�!>�疽-��=te>\Y�=R�=*f?��
?��
?�a����	�C�����A�]�L��<g!�=~{�>�\�>��r>��=�:f=]С=�\>W˞>{�>*�d>C��>(A�>ĸվp�3��?�^,=�~c>�Z!?bG>;��=���=,�9=t5�ʵ��_r��Ƚn����=��<5$�=;���#?sLο�C�?l�">� ʾ:�"?�e��n'�ؘV>թ�=Z&���?�2�=se�>�T�>�h>?��=�@�>'�
>�FӾL>����d!��,C�X�R���Ѿ|}z>�����	&����w��RBI�n��ug��j�O.��X<=��˽<.H�?z����k��)����S�?�[�>�6?{ڌ�����>���>�Ǎ>�J��j���[ȍ�hᾥ�?C��?�
{>�G>OmW?��
?�0�zʾ	��A����B�8���(�p�$n��Ҕ��_������.�?�Ԅ?)�(?�'˽�̻>Z�r?��N��y����D>�wa��d�+`ȼ���<��g7��������a��:rS?{�w?`+N?���>��G�����[�=���?O-;?�Z??�N?���?�R����>�I�>�>L?�e>?t��>u^�>�[�>α>�1>��=��!��e��.�����8���r"��y%�=Bn�=:]Z=��U<q5�<��=����7%ƽv��<<.�<N��:���;�$9<*F�=��>�RY?�$�>"L�>ۨH?k|��@�3�N՞���>ceB>�Ⱦ�̾;�����G >[�c?��?�L?�%>��F���ʽd�*>^"&>.�#>->g>�z�>�G�޽Wg>}>K^=~%�=<zB�O����8��&�P�W>�AS==��>2�>ͤｸ��>#N��nϾv�f=��i]�؊X�ΛL���,�|��얇>i	\?��/?�	M>�.�����ɲa�].?�~L?��J?�g�?�(�;'Gվ�]Z��q�)5>B�$>A]νZ��顼�f[��� ��g>`G>(A���Ǣ��b>^m��O޾Um�p�H��'�ʏS=$j��!R=v�Y@վa4~�-p�=��>bQ���^ �(���8�����I?��p=�\���xP��]�� :>��>Aa�>��,���p���@�Oڬ�~S�=Z�>t�;>���x��T�G����w>�>>QE?:W_?k�?	"��^s�X�B������c��oȼ(�?6x�>h?�B>���=圱�����d��G���>���>y��-�G��;���0��I�$���>99?��>h�?g�R?��
?�`?)*?RE?�&�>���x����A&?6��?��=��Խ�T�| 9�MF�{��>{�)?�B�ڹ�>K�?�?��&?�Q?�?d�>�� ��C@����>{Y�>��W��b��B�_>��J?���>j=Y?�ԃ?l�=>W�5��颾�֩�V�=�>��2?�5#?R�?���>X��>����=���>�c?�0�?�o?L��=?�?�:2>`��>���=ћ�>3��>�?2XO?!�s?��J?ؑ�>Y��<�7��r8���Bs�y�O���;N{H<��y=9�� 3t�J���<���;Yf���H��t��{�D�������;u
?�T%>OӦ��>,��[��dy>��=����ҽ�� ������+�>��&?Qy�>{9	=�v�=�]>��?����I$?݋?��9?g���>Z�=�	�0��<�4c>d2?��m>a�(��Q��Vȉ�d�1=z�|?ou?$�ԾGj���]?�k?��Ͼ2;��@�g�Q�q>1���N?�"G?,k�=Y��>��?t#|?{8�>�@��A��y���mNa��۾M�$�k��>dh��Y��s�?q�u?�Ó>��F=�C��r�w��b�9G&?g\�?�	�?Kݐ?>��=ׁ�S����}v��� �?Z��>>��F;)?l=�=1���ƽ�y�&��g�	�*Y��3�Y��U�$|�&M�p���W.?U�?�i?��m?;�
�l·���l��ʗ�MXI�j��\!D�K�b��%Q�:.5�^oo��׾�w�������]r��Z�gDB����?N'?)|0��4�>c���?�L̾��B>�Ҟ�m���;�=4���^C=��]=�ih�U�/�jO���X ?��>�X�>��<?S�[��E>��>1��l8������2>��>+��>�1�>eb:��-��C齄ɾDQ��Y3ս
7v>�zc?�K?�n?|h�k%1�Ɔ����!�}�/��Y���B>fu>w��>̶W�Ŧ��8&�X>���r����jw��3�	�s�~=ֱ2?�,�>,��>UN�?2?)z	�7k���ex�J�1����<b)�>i?�=�>��>I�Ͻ�� �2��>a'l?��>	â>ց��F/"�}�|�τ��K��>�A�>�L?1�{>=-���\�'�H��1�8����=X�g?@����`��L�>��O?CɻSR�<�+�>�|�Iu ���2*(���
>�	?~�=�:>I�ƾO���|��c��LP)?M?XӒ�n�*���}>�"?�]�>�,�>�)�?��>eþ��O���?G�^?�0J?�:A?Z�>g�=T���5UȽF�&�9�,=���>� [>bYm=vx�=���\����*EE=��=�Lϼ���c<{+�� �S<��<�4>�jۿ�K���پ{�1q���	��D��
���K���w��"��0ᙾ�x�+���'�L�V���b��k��C7m��_�?M�?�ϓ�\��1t��\k�������> ep���}��=���H��0���P�Do���^!��EP�Z>i�A�e�T�'?�����ǿ갡��:ܾ ! ?�A ?�y?��?�"���8�٭ >$D�<*����뾣����ο"�����^?���>��/��c��>ƥ�>J�X>�Hq>����螾�2�<��?-�-?��>��r�)�ɿc������<���?*�@�|A??�(���쾦V=.��>/�	?�?>S1�GI������T�>L<�?���?�vM=u�W���	��e?�r<�F�2�ݻ��=9<�=�J=�����J>�U�>���SA�<@ܽ��4>qڅ>*{"����u�^���<.�]>��ս�7��6Մ?{\�qf�2�/��T��T>��T?+�>�9�=�,?l7H�@}Ͽ��\�+a?�0�?ئ�?��(?'ۿ�yٚ>`�ܾ{�M?=D6?g��>�d&��t�L��=�+�ƕ��1��q&V����=s��>��>��,�^��݅O�"V��"��=����=N��i+�;.�+��=$��=&�b=�����!-��J���T�&�/�UO��]=?9n=A��=��>v1�>�&�=K�K?z�j?O�?y�>���b�M��ϴ�=� ��K���騾�CV�jL���wȾ�쮾)�	��q5�F��lC��7#=�3�=�5R�����)� �R�b���F�Z�.?1p$>��ʾ��M�$�-<)nʾD����턼�쥽�*̾�1��!n�T̟?/�A?1���F�V�����C��o���W?�D������ڗ�=�ű��=t%�>���=���X"3�m|S�)\0?zp?����M��Nv*>R1 �G�=V�+?��?O`<�^�>]_%?B4*����t�Z>�Z3>���>K��>[�>k��#�۽��?�T?-���$��I�>g����z�^�`=�e>y�4�����[>Y��<ǰ��X�������<7*W?`��>��)�������1���H<=ڵx?��?�G�>Ńk?FC?��<�w��x�S��1�6�v=��W?�"i?{�>ˁ����Ͼ����h�5?��e?/�N>�kh�d����.�;T�N"?h�n?�b?�^���r}����o���K6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?p�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>��������=:��zj�?��?4Ī�\�h<����Al�K7����<�j�=[ �`&�����7�$�ƾ%�
�o���]����Ԇ>�`@)��*b�>	�7��D�MeϿ����оl r��?�
�>��Ƚ������j�Xu�ewG���H�̋��6O�>��>����.�����{�Cs;�窟���>�2�y�>t�S��*��!���2�5<�><��>%��>�.��U佾�ę?�a���?οH���L��W�X?Jf�?�m�?�m?�F9<��v�[�{� E�|/G?o�s?�Z?�%��@]�ɢ7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�
>Y?G�K��A�F?��Z}��תH��Ⱦ��*��~;�����w�F���1�&�?���?n��?^��t���A?-�>��q�Wj�u��v��=�:�>��>���=�s�>�I��R�{�+=���?<��?���>�m��<֗��>���?G��>d�?��>㞙>���=�s���6�A>�M>=��=��	?��C?`��>�D]=��r��$�XlF�d�X��@'�^\9���`>��T?�P?:2�>%����$;�� �<���1��~��mZ����:�+�wQN>�c>IG>w����^����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*k������7�48Ծ�x$>	�J>�`> �T��O�;���=�">�X)>ƢV>�P@>6g�=�K>�&�>be>0ᬽ�z�X.��x��@՟�`$�!Oྉ��.Ӝ�I��(����vоn�q� �J��Փ�h�/�-/"�M�Q�_�:�00�/�=k#W?a�Q?�l? ?=Q[�@_>�����N=�l�*��=�$�>�`2?�I?��'?�4�=C��	\d�甁�J&�����3��>w�P>��>��>���>)��ZG>x�9>)�>��>÷5=����=5M>b�>���>�0�>�C<>��>Eϴ��1��i�h��
w�h̽1�?���R�J��1���9��Ӧ���h�=Gb.?|>���?пf����2H?%���y)��+���>}�0?�cW?�>��o�T�1:>:����j�5`>�+ �|l���)��%Q>wl?o�f>'u>�3�d8�t�P��s���u|>D36?趾zC9�ּu�/�H�O^ݾ�DM>��>�D��i�����(��oi��{=�x:?�?���w۰���u��=��\ZR>�<\>%=R`�=�PM>1cc�.�ƽ#H��.=`��=��^>!J?_J,>uď=S�>h���2P��}�>@�B>��+>F@?��$?��'�������G.�Cw>���>'�>>XyJ���=�q�>a�a>�7�����X�s�?�zkW>�W~�*�_��Hv���w=�{��t�=��=5X �*T<�K�&=(	�?�Ǘ�Ǯ�r㳾FԎ��k�>��?3j½7�=� ;��쨿������?��@�`�?�3�)y���V?���?j4m9��x= ��>�ܓ>�&��ʒ=|W?i
�>^_:�ZN��Al'�甍?Qٓ?>X=��`�18g��^�<\�$?P���Ph�>{x��Z�������u�w�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?�I>���?�s?ve�>��x�V/�r6��#���|�=�oc;�p�>w>���5hF�ؓ�Bh��ʸj������a>��$=�>�7�s+��C;�=ŋ�rE����f�b��>� q>�I>�[�>�� ?�Z�>���>R=fI���݀�÷���E?���?��O�x���=<���=�v��G?�9?�)�=Y���z�>1�\?��l?�3>?T�x>j���Ŝ��@Ŀ����̡<��]>�]�>���>� ���nf>6�ܾ!�d���|>B}�>��u�꾱����I=��> ?���>v�=H]'?n]-?��>�Y�>
xX��ȏ���U�.;?S**?oK:?��?�EF?�kԾx�P�v%��������G�ﷻ>;|q?��%?C�/>�yp��w��2�׾g=f��!��`i?�"�?����?c\�?�V?� 1?��=�ߕ�ż������a=Y="?�&�/�A��o%��X��?��?'��>첒�f��L��)�
����0?h�\?�&?����_�?����|�<ڒ��({���4<��Y���>�>�p���1�=�#>�T�=*^j�O�9��� <p�=�ɔ>B �=t<�MI���,?7�:��(��s��=]0r��lD���>��L>\-¾V�^??�j�{�����wr���VU�r�?;��?�7�?߾��ӄh��=?	�?��?�X�>�ͮ�^�ݾ���4Kw��Gw����#>��>h���i��D���U=��Xσ�<�Ž�?2�zn�>�'�>��
?4v??"U>�U�>�񏾶�&���à�d\����9u6��p-��������3$��A8��q���jo�/��>\p�C��>�6
?T`r>^	}>���>
���>�F>`:y>�ؤ>�KR>F�%>���=t�(�9N��S�\?�;|�!�J���ס־��?��p?_��>�8��㉿��!�X��>�G�?���?Ͻ�>a�L�Q9<��U?>�?r�j�n#?�Ld;.�<�ݤ�����(o��=wq�Uj">�]~���#�G�d��nb
?��(?V�1>a�� $����:�n=N�?��(?�)���Q���o�θW�S�1���6h�Mj��Q�$� �p��쏿�^��%����(��r*=��*?j�?ь����!���&k��?��df>`�>`$�>-�>$uI>��	�s�1�h^�M'�K���hR�>[{?�>ϰI?)O<?��O?>ZL?���>�>hE���"�>��<�m�>CG�>��9?��,?[�.?�?�*?��b>h�������w�ؾ�5?�?*�?�� ?d"?�ӄ�	Mý����nO���x��·��e�=R��<�mֽq�y��*T=hU>��?nZ!���5�����J>{1?���>�a�>����Ð��-�n'�>�?�ɪ>z�辢�o��B��U�>*��?]���M�"=�$>�8�=�RS�J|;�m�=� '<	nt=���I`,���w<�v�=Zd=(�<���<2I�<�	���(���(�>��.?�5�>���>�m|<��#��Aľ�Ӂ>O�s�z$�>�?ټ�#
�����3����p��>�<���?'=�?��=�(=>�%�=�m߾�7ݾg/�׳���+�d�>��[?N?��?��r?�(�>�=ڡ��������ٽ�GV ?y!,?��>�����ʾ��։3�ڝ?i[?�<a�2���;)��¾��Խ�>�[/�]/~����;D�ꅻ���;��2��?�?ZA�U�6��x�Կ���[��y�C?"�>Y�>x�>Z�)�x�g�i%��1;>��>cR?V�>"P?�#{?�9[?��T>�(8�$.�������
%���">Y @?��?��?ޝx?��>w>3�)�X$�l������������O_[=��Z>��>��>��>��=j0ɽ+ʯ��=����==^a>/;�>"c�>]z�>�Dx>tE�<��G?��>���?�����⃾�;�6�u?J`�?��+?�8=����E��r����>&b�?X	�?�*?7�S����="/Լ`����r�eH�>G�>~Z�>-В=̛E=��>�e�>r+�>����x��8��\P�3?�:F?���=��ɿ�F������$�>�8>0`(>tݞ�yA��w�,<�FȻWF2=�|#���B�����m���l�%�����t�>B���E>m=��I�3���J<Sf�<�Z��'h�����(W(��tU�YüfU�=��=���!=o?(>�껾��t?�@?�>�PQ?/	 ?�.�=�X%>9>�>=�>�j%?���>_uc>2�Ӿ����A���ׂ�����^پfe�+�ɾa�D>'�2>��B>��=�Ü>,g�</j�=��F=���=k��=)���|>E�
>>�h=�fV=H�<>��>3w?����嫝��'Q�gN��:?��>3�=��ƾG@?B�>>3��Η���^��,?���?TQ�?��?�mi��k�>����C�����=(���%2>3��=��2����>4�J>X���@���'3�?��@ס???ዿ,�Ͽ{/>�+6>�>��R���1�ś[���a�6�Y�5~!?�4;��̾Qd�>
ջ=߽޾�zƾ��,=��5>>�b=jb�1X\�^ϙ=ęz��"==?Nm=��>�D>F�=���<Զ=O�H=Z��=�hO>�ܛ���7��.+���2=���=�b>0&>���>A�?2b0?`d?�<�>�n��
Ͼ.����>�`�=�#�>���=�MB>�u�>K�7?T�D?F�K?���>$��=e��>��>�,���m�X徟§��H�<V��?�Ȇ?�Ҹ>�6N<��A�5���i>�7�Ž&e?�R1?at?$ߞ>/���߿R (���/�[.��uF�;��<=Or��Am�p+�����ڽ~��=y��>ׯ�>�A�>��|>��:>�I>��>��>�$�<�ڃ=�~��w�<�ȅ��w�=D����	�<�hϼ��������v*��񚼑�/;���;%��<#�<6�=N�>�l>y=�> 
�=ۑ��8�0>�;����M���=j4����B�fd�F_~�L�.��z3��%J>ǊW>Ҕ�����V�?�u[>�<>d&�?]�t?EZ">�'��gվ�n��'+k�$�V�i��=G�>�F�<���^��K�&�Ѿw��>]ߎ>�>��l>�,�Q#?���w=��0b5���>�|�����)��9q�)@��	���oi�YҺ�D?�F�����=`"~?ذI?]�?��>W���ؾ	;0>�H����=k��)q�_h����?'?���>����D��H̾K���޷>�@I�2�O���U�0���2ͷ�7��>������оm$3��g�������B��Lr�\��>&�O?��?\:b��W��KUO����_(���q?�|g?/�>�J?�@?&��z�r���v�=�n?̳�?T=�?x>	�=)���o��>�a?3�?V�?��s?�n=�ՙ�>�d�;�T!>����n�=�$>�#�=�3�=N
?��	?��	?�����
�A��D���]� �=�^�=9�>�,�>�s>ȼ�=�li=�a�=�UZ>���>�~�>�xb>z��>���>�3��E�S?�0����>pIJ?���>����q���dF=Ό�=S57�<ߖ�m⭽7��<��>bM����Ϻ5�?�տ`?�?j�.>9)�M��>ҕ����t�;��>��>R���>�>Żhh]>���>�o�>�ql>�E>��:�FӾ8>����d!��,C�2�R�?�Ѿ-}z>�����	&�ޟ��w��BI�9n��Tg�yj�L.��><=�&ͽ<H�?ڻ���k��)�,���_�?�[�>�6?mڌ��
���>���>�Ǎ>�J��R���Oȍ�hᾢ�?1��?*:w>q�D>j�j?ge?$�X��T���:s�/T���(<��i�"`��i��xZ���������E�}?�q?�&?&�ռ�2�>z��?U~P��]ӽ�Z�>�p���i�藷<FDM=|O������E-ӽX������>�A�?�0d?�L�>��Y��d��|,>\A.?/�?"z?)<?3�@?�Uݽ�!?�1>�?��?�_2?�="?*p�>��=�O�=��)�<
������m꽱K�4p��`l=S =�X��M�8$|=fLK=�����l�4F<���<�9$=:K�<�^�=��>�à>��Y?��?��>�29?�N��H��Έ�~��>�+
>G�ɾ��N�����Qm*=G�[?��?a�N?�8>��R��q��8�8>�A4>:p=>��+>�Ϭ>��Ž$�t
�<#;=j�=�>;=�ڪ�9����M���t�T>I�%>So?��> ̬<:?륾�OȾ�_=>x�=����\#���@��y$�Kµ����>�I?�mA?a��>9��dE�=ba���'?�23?�%&?"1�?���=����M�9�
f�y��>ۏ�=����:���%��2r;��j�>}5�>z���࠾-Rb>j��|t޾ǚn��J��羜BM=.�bV=���վ�7�J��=�$
>������ ����b֪��1J?p�j=Xu��qaU��p���>���>ޮ>��:���v���@�*����2�=:��>��:> T���ﾄG�=7��>�>2QE?-W_?k�?�!��{s�N�B�!����c���ȼ�?x�>�g?�B>��=`�������d��G���>���>���>�G�`;���0��S�$�.��>39?Ȩ>K�?b�R?��
?��`?_*?dE?�&�>���i����A&?2��?��=��Խ��T�k 9�jF�]��>y�)?߷B����>F�?�?��&?�Q?ݵ?t�>!� ��C@�i��>�Y�>��W��b��@�_>ǬJ?��>B=Y?�ԃ?��=>Q�5�kꢾ�ש�W�=�>��2?�5#?.�?��>�,�>q.�����=*:�> "c?L,�?r�o?Dv�=��?��2>��>nZ�=�v�>���>��?� O?��s?��J?G�>�O�<]孽�Ƿ��fs��=B��B�;_V<!z=+~�~�s�|T��z�<�ݵ;�ܳ��y��y�\�D�9:��]Z�;���>G�]>�����L>Z�������'1>Â�=\첾��ʾe�n��#I<��v>C�?�<�>�[���;� �>��>#��sC&?n��>Ȯ3?���=3[a�(Fھ�����X�>�;?Ѣ�=��b��������&R=n?ĭl?�~���>�/�Y?�d?��
��6������=��=V?�B?1��=0��>�?r�w?�ƈ>Ҿk���v���I\���ҾO(��O�>GK����e?c�g?���>�I=���|�¾q�k�o�����>�Ō?Ƴ�?���?V�=H�u�u�Կ�us���o?d��>����e�/?�^i�����"j�D�]���˾uf��
�TD��I2��ex��mm�H}X��u�=�8?\
�?Xz?t�j?���҃���;������]���!���G�M�a��7:�ޯ,�V�2D��&{����E��9#=����A�#��?'�'?�/� 5�>M͘��񾔸̾qC>�'��"��1�=Z����@=��\=��h���/�0��)Y ?d��>�.�>l�<?U�[�F>�\H1���7������3>�ס>���>���>Tߧ:j�-�Z�N2ɾS���Ҷҽl5v>�xc?4�K?K�n?&m��)1����T�!�,�/��a����B>�n>鼉>�W����9&�X>��r���w��4�	�(�~=Ұ2?)�>5��>�O�?�?�{	�wk��oix�ć1��z�<�0�>� i?>A�>E�>��Ͻ�� �:��>rl?��>`ˡ>�Z��H�#���*������>���>� ?9�>�\&��L]�����䏿�+9���=��e?�}���Xd��B�>��N?��.�0��<qϞ>������U���$��I>2�?e�=W3;>�4ƾa���<}�����?)?de?�ے�"�*��q~>/"?C!�>�>�)�?>5�>xAþ�[�2�?N�^?�J?�+A?�9�>M�=bi���qȽ��&�a&.=㢇>�[>1en=j��=��Պ\����ªD=��=�3̼tA��n}<����Q<��<�&4>=mۿ�BK���پ��W?
��爾x����c�����ya��#���Xx���	'�>V�n7c�����l����?�=�?耔�a0�����&�������f��>T�q�H��������w)��ږ�R���Bd!���O��&i�a�e���'?ֺ����ǿ밡�;ܾ�  ?�A ?ݧy?M�o�"���8�\� >S�<z�����[�����ο=���\�^?]��>}�J/��I��>ͤ�>��X>�Hq>����瞾�5�<[�?�-?ס�>��r��ɿn�����<���?��@�{A?s�(�l��xV=b��>��	?T�?>nT1�	I�l���R�>?;�?)��?3eM=��W���	��e?�h<*�F�޻U�=fI�=�K=�����J>|W�>ҁ�qRA��Bܽѳ4>
م>�q"�_���^�b]�<Ό]>�ս3��SՄ?>z\��f�ߤ/�5T���K>��T?p'�>�6�=[�,?"8H�	}Ͽ��\��,a?�0�?J��?��(?�ڿ��ޚ>�ܾ��M?C6?K��>e&�}�t�\��=@�༢���E��&V�'��=Э�>�>��,�����O��昼���=����aƿ�T%��C��=of�9�kj����q�����E�u��٩m����N_=f=�=(�Q>0�>��U>�rT>W?��h?X��>��>{�I,���;i�;�v�����`��2�S����뾕�ݾ2������d�yǾ� =�;�=7R�m����� ���b���F���.?x$>4�ʾ��M�f�-<pʾi������᥽Y.̾&�1�8"n�͟?M�A?������V�����L�
�����W?�P����ꬾ)��=e�����=9%�>���=Q��� 3��}S��w/?,�?!����픾/>������<��*?h�?��<���>n`%?>�(���)�R>��/>�(�>JW�>�@>�"����ڽd�?�dT?� ��'d��7��>�澾-�{�!YL=�,>�03��˼�Y>ؗP<&v�������ˁ����<P(W?ߟ�>��)�:�sk���O���<=��x?��?�3�>}{k?��B?�
�<�m��l�S��%��1w=+�W?�%i?!�>�����о����w�5?�e?�N>�dh������.�S��#?3�n?�a?�j���t}�������wb6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?p�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������u��=Jە��Z�?f�?i����(g<���ll��n��8q�<]ȫ=C��a"�
��8�7���ƾݺ
�����忼H��>�Z@s]轀*�>�@8�7��SϿf���]о�[q�0�?�{�>��Ƚ����=�j�Mu���G��H�4���Ma�>ެ>���������{�;��Ť���>�
����>�ET��a���ߟ���5<�M�>Ki�>�ކ>X"���Ľ�-?����Dο2���V��lX?�>�?Qg�?OK?b](<�Mw��z�?��CG?��s?�*Z?՗(��]]���5�(�j?�_��xU`��4��HE��U>�"3?�B�>M�-�ϱ|=�>v��>Xg>�#/�o�Ŀ�ٶ�B���]��?��?�o���>m��?os+?�i�8���[����*��,��<A?�2> ���J�!�=0=�PҒ�¼
?O~0?*{�e.��e?|<��S�����X�=S� ��Ҧ
�g:J�?��qkw�t ��t�9����?OK@���?J�ݽ��8�!�>?��>������
)��>'s�>d��>���>M}�>C�ľ6(�"�<o��?z��?l@�>08��p���e>��}?Qܬ>y�?*��=L�>��9>D�q����-9>M�F>��=F� ?��H?	6�>~�=�*z��"�i B�$T�i���@��Ɔ>��`?u�??T��>��<>	�<.�#����@c���(BQ� Ƚpb��f��=��6>���>���������?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?qQo���i�B>��?"������L��f?�
@u@a�^?*��׿x����ߞ�r|��o]�M5\=�a�>E�G�O|�<{a7=?��=��h=X��=�v>q�>�7>�L>л<
��=�[���l�0���L	����J�ѐ��M���z��Ӿ
���o챾J2��c���y9�LΜ����v2K��>c=&��=��U?�R?	p?�� ?3�w�ɓ> ���o�=*=#�#�=�G�>�d2?��L?ц*?y��=����#�d�oZ���A���ʇ�k��>�I>���>�<�>m*�>���7��I>�?>℀>� >��&=�>�Q�=��N>ab�>���>�s�>�C<>(�>?ϴ��1��R�h��
w��̽*�?<���*�J��1��q9�������h�=(b.?�{>���?пf����2H?����_)�Z�+�g�>��0?�cW?М>@����T��9>����j�<`>f+ ��~l���)��%Q>ul?f�f>#&u>�3�bg8���P��w���\|>�26?r䶾5<9�վu���H��aݾOAM>x��>.D��k�������7yi�l�{=�x:?�?�#��Oݰ��u�tE��JR>"3\>nT=$e�=-TM>Vic�u�ƽzH��.=���=3�^>�J?�`,>�)�=��>����P��{�>�,B>��+>G	@?��$?�i�.�������yh.�h�v>V��>B��>s�>�pJ���=���>��a>�/�Q���/��z?��wW>u~� n_���u�Dx=�<�����=�+�=���� <�<�&=W&�?����yɁ�l��U_���?��?�/>Z+>�w>�[ˣ�wM��e�?�'	@�Ɣ?.����uj��.R?¨?g�0���=�d�>&��>��lv�'��>�K=��a��󮾶ZԽش�?Oג?#�ԼQÀ�/�o��.-=�>?�~��Ph�>zx��Z�������u�s�#=Q��>�8H?�V����O�e>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾;`Z����>һ@?�R?�>�9���'���?�޶?֯�?}0I>���?"�s?�h�>yUy�a/��:������~�=��i;Dv�>��>����lF��ړ��n����j����?�a><�$=��>
%佒9���=�=ͣ���?���g�Ζ�>�=q>`�I>�Q�>�� ?�y�>���>3L=K���������I?]��?����r��=
�=4�s�k?�5?��8��ȾP�>]Z?�z?I/T?�_�>��R{�����긾��<��V>K	�>���>�/4��7U>U�׾�DO�T��>| �>p��MᾺ������{�>�#?ѵ�>�P�=Q- ?|F7?^=���>V�L��e��)ug��r?}w?�?+x?�N6?&ξstP��O��:c��=�V����>K-p?�"?Sd">G�~�kc�vW��.���t9����s?�V�?�჻U,.? ��?g�o?}u)?"D�=J������gW�=��!?�!�|�A��R&����v?@P?���>�)��� ֽ Z׼8��Cp���?�,\?�@&?���$a�G�¾Zy�<w #��FT��q�;��E���>��>�D�����=C>��=�Jm��"6���g<�0�=yb�>\��=&�6��_��=,?ֱG�ۃ���=�r�CxD���>xHL>K��i�^?]n=�5�{�}���x���	U�� �?��?(k�? ���h��$=?�?�?o"�>J��}޾y���Ow�}x�jw���>J��>��l�D�B�������F����Ž#����>!��>G�?_��>�u>Ȇ�>�i���>���ؾ�m�:�h��b���9��32���h �W�FؽӴ���A����>L ݽ�ʳ>��?O��>E1�>=��>�]���`w>@�>c�4>�ܖ>j� >��=��%>;b>)~�W�`?�ɶ���.���^g.�2�?�H?,�?�R��匿$<!���>J��?Qͭ?e3�>�~G�b�C���4?�T<?�M��o�?��껶�X>�->W{ľe�1��V�=FIp���0<���!�$��e�.-]�6�?�r#?ƄZ����.�7����=�n=N�?��(?�)���Q���o�θW�S�3���6h�Mj��Q�$� �p��쏿�^��%����(��r*=��*?j�?ь����!���&k��?��df>`�>`$�>-�>#uI>��	�s�1�h^�M'�K���hR�>[{?<΃>�?I?B�D?.T?#K?R �>dI�>?+��(��>�<��>���>]�6?Q�#?,�'?O?��,?;)i>���D/��1�پ�?�q?��?|?�V?�\���'�LA�|�������������=��e=(���R��(k�=��A>��?�'���9�q���5>/G4?g�>;��>�a��@��rc=;���>Fs?���>=���_�p���)�>X�?���޼!=5�*>8#�=)����(��<�=*\��&�=wW����1��<��=�s�=���<�g�;�h`�0$&<Z>�>��1?�l>r�>{G �Ϭ�L՞�� >ǅw�tcZ>޸"�m��/o��Vǒ��i���<;ʙ?�W�?~ׁ<$x>F[_>��r��	1	��U��#���x'?��n??�N?h�?�9?�e�>+��w�����������t��??y!,?��>�����ʾ��ԉ3�՝?h[?�<a�F���;)��¾��Խ��>�[/�\/~����8D�ꅻ���*��/��??�A�T�6��x�ܿ���[��}�C?�!�>Y�>o�>c�)�{�g�k%��1;>ߊ�>SR?�!�>W�O?0<{?�[?QmT>g�8��0���ҙ���2�B�!>@?ձ�?H�?&y?>o�>��>ѳ)��྄T��1��"��݂�|#W=SZ>2��>�)�>&�>��=GȽ�X����>�b�=��b>��>3��>��>��w>�X�<2�G?��>%X��Ñ��社�ǃ���<��u?k��?j�+?3=q��#�E�qI��QB�>)m�?���?�2*?��S�G��=D�ּ�۶�P�q��%�>k۹>�4�>Qٓ=�F=._>�>���>2��_�<r8�.�M���?F?��=n�Ϳ��r��#������vgz>: ������w�=Ol�����>���=���m��F�l�c�^�42���mƾ�z���U;�^�>�kg��!�� ��:�@Ѻl��� �qE����c�9;+�j�=��A�z'��T����剨=�[�=�!;=�����z���;�?-1i?�>-C?�O?�
�=�$>�T�>T >�<?��?:�s>�� پ�.��0�&��w��<�о�e��]�����>�΢>���=�\�=��>�=|�x<��<��>�@{<�<��=�3a>0f�=^6>��>�h>u2w?��������"&Q�@�{�:?��>m��=N�ƾs@?�>>3��d����\�-3?���?�P�?Q�?�hi��s�>��@t���A�=MK���2>���=��2�.��>̊J>����?�����3�?��@-�??�⋿��Ͽv/>��6>S4>D�Q�T�2�'�U���[��~`�r� ?�9��Ⱦ��>��=��ݾ8Ǿȶ=3>-eb=���>\��w�=Yz��M=�
|=q�>ƩG>���=�z��H�=(f6=4M�=�O>��� �9�p?�|�(=ϙ�=#�g>��)>��>w�?`]0?sd?�5�>enn�W�ξ�b���m�>�>�=fz�>�|�=�4B><�>��7?��D?� L?���>�=6º>�(�>X,���m��徦����6�<ړ�?�Ć?���>vQ<�A�U��I>��pƽ�?�L1?��?���>"��tӿf�+�4�"��&ʻ"�<����<�w�����Z��=��=| �������$e>Q��>>���>��>B3�=��>]R�=�q����<���;��\=��2�� �=i��;�û�P�;E=i����f�T�e=)'�Z�p�X�l=R��=���>�J>���>&��=~���g/>KĖ��L��˿=&d��H3B��+d��G~�/��J6���B>�1X>�؄�#0����?�Z>�H?>��?�;u?P >~��H�վ�H��!Ke��cS����=��>�.=��~;�J`���M�ZoҾ���>���>��>��l>,��"?���w=C�`a5���>|�����&�f9q��?�������i�;�ӺПD?�F����="~?�I?��?H��>u��I�ؾx80>�I����=��S-q��h����?�'?��>���D�}H̾���޷>b@I�#�O���?�0���Rͷ�4��>������оh$3��g�������B�~Lr�]��>�O?��?<:b��W��HUO����>(���q?�|g?3�>�J?�@?-&�� z�r���v�= �n?Ƴ�?U=�?�>55�=�z��7�>uX	?3��?���?qs?1�>�3`�>�i�;m�!>�蕽�#�=��
>,�=V�=}�?\z
?�_
?vz��@�	��d��|��]�2d =h��=uz�>�>!r>���=��e=��=�P\>`�>E��>>rd>�ƣ>�̈>��ݾ4%:�9'	?1��<9�>fjA?" >�����s�웹=ا=t�ͽ�V�����B��F��=�
���"꽷�n�<s?h�˿c�?>~>�����#?�K���^;�XNU>fL >!����k�>���=s�7>��>��>�;=]��=��e>�FӾw>����d!��,C�U�R���Ѿ�}z>�����	&����w��VBI��n��xg��j�N.��X<=�L˽<+H�?�����k��)�����V�?�[�>�6?�ڌ�����>���>�Ǎ>�J��j���Zȍ��gᾦ�?E��?�kq>b�P>x�]?5?��F�H����2P�J�����F�g]b��7`��Z���Ί�Gp�-1�6��?.?�.?�M�M��>���?1�G�����~��>Mri���J��N��>����M�������y�_#
<�G?HV�?MkZ?.2�>��0����&>^Fw?~�W?�݁?n|f?5y|?.e�=q�?���>U�'?��?~'?���>�߽>�m<]�/>��!��D��]0� ��v�#��v��SE��U=��!>jG�=�l�}=�u=ϓ���^һ��X=d�<���7�= �l=%S_=�Ϧ>G_\?�	�>��>KR4?2^,���%�i�Փ?�^=򮞾�u��Z}�������=��^?sܮ?d%T?�+>��H�,0$��<2>��r>�(/>f>"��>�|����"�tZ=E->#��=�|=�&U�ʡ��Bt��\y�3�=��2>q?~>�K����>՜��_�Ⱦ
CU>g��"�+��ޢ�>]���I�_.��-e�>i9?\�?ץ{>r���* �yjU�b^/?!�a?yEF?"��?���<X>�R_���N���> 9�=]C,�ݡھ�Ŀ�鯿�&�0��>��E>wz(�ᠾ�Sb>V���s޾��n�fJ���羛KM=u�8]V=��^�վ�6����=�#
>����� ����l֪�\1J?}�j=�v��*]U�Em����> ��>�߮>��:�^�v�W�@�����H6�=���>��:>�o��g���G��8�z>�>;QE?2W_?k�?"��Zs�V�B�԰���c��ȼ�?@x�>h?�B>���=��������d��G���>���>���?�G��;���0��?�$�
��>59?��>�?N�R?��
?��`?)*?NE?�&�>I������B&?0��?��=��Խ�T�� 9�IF�d��>r�)?Z�B�͹�>@�?�?�&?�Q?�?e�>� ��C@�Ĕ�>zY�>��W��b��.�_>��J?ߚ�>t=Y?�ԃ?��=>X�5�ꢾV֩�/V�=�>|�2?�5#?T�?���>e(�>�ġ�=�S�>��b?�B�?�3p?s��=��?mJ3>.��>�=�;�>�9�>��?��N?��s?S�J?���>���<8X��x��!u��;X��P;�z6<hz=�a�qy�+��~�<S+�;#���wC������@�H��됼`B�;?�?�3>}�����<�`�ȏ��<>
ؽ<�_�����p(��M��i��=�3/?_�>�/;���=��>���>8c�D�-?i��>���>%�ǽ.z���rf�<R��>H�?��>dH7�]���;����=oe�?�8~?�u��a &�`[?Grm?�,ؾV��y�¾�h>6��P�D?x?��=���>��?��?��>���]��D�������7��]�0=�ȅ>/��>U�)c=�(?���=f�>/�>vgu���u�=櫾�V?��?�̣?�i�?�ۿ>2!Z��t��^h뾣ߠ�h5?Ќ�>�r��o*?����jP���$���E���	�!x��ɤҾ�����O���L罒$D���:�=[D? ȉ?��M?R�Z?��
�!v���u�y_���4J��N=�M�/��b!�0Q%��+4��D7��	p�����N'��s�H=@���B����?`�'?.5�J��> �����o�̾� A>/4��R&�mc�=/���>==�\=y|f�'�,��6���{!?���>ª�>��<?V�[�Q3?�O�2���9�������)>��>�m�>f��>]1�8�)*��Lٽ�ȾgB��j�ѽ��u>6tc?צK?]�n?zQ ���0��o��+r!�3�0�p)���=C>�B>���>V�W�g��k/&��I>��s�s�Γ���	�ۂ=��2?\�>C3�>L�?�?M	�Oͮ���w���1�+y<��>E�h?��>$D�>~ν� �!��>Do?=~�>5�L>_�Q�P<��;s�[��� ��>���>��	?�F�>בн�z\��a���ߒ�x1L�)A�=A�v?Hx���n�ς>��<?���;�H=��>U(ؽ�*�Y��7�����=�?�?�=��>o����	��}���/����)?2�?պ��B[*���}>�!?�q�>�٢>K�?�͚>b(ľ�P�Y�?��_?�J?�@?��>�$=����-Ƚ�X&��\)==i�>�SZ>!p=^��=1��̓[�|$���@=��=��
����<l沼�b<���<hn3>�mۿFK��پ&�,��2
��ӈ�$����_����PU��*��=fx�d����&��V�
6c�]���V�l����?:�?Yo���������W���q���趽>�~q�;�K���$���&����ྚĬ��d!��O�{1i�2�e�P�'?�����ǿ򰡿�:ܾ4! ?�A ?7�y?��8�"���8�� >tC�<�,����뾭����ο@�����^?���>��/��o��>ޥ�>�X>�Hq>����螾�1�<��?7�-?��>Îr�1�ɿc���q¤<���?0�@�|A?(�(���쾟V=���>�	?��?>&S1�ZI�����R�>�;�?���?tjM=��W�V�	�+e?zf<��F�
�ݻ#�=jC�=�E=4����J>W�>��'YA�u7ܽ,�4>�ׅ>7t"�é�!�^�Gr�<�]>F�ս�>��ݼ�?�[��f���/��f����>нS?��>��=�G+?RHH�|FϿ�^]��a?9�?���?w�(?ڿ�zY�>��ܾ$M?)�5?��>@�%�%�t���=�Ү��X�:��U���=�=�>3
>ܟ,�z���,J�z����n�=B$��:ÿ�C�B��mU�T�=�
=�X�ݖ���_�ICr���p�'��'=��=>�(>��j>]f>�3>�vO?jj?��>�^�>"��=ɶӽ՝���]�<��A�E�f�H9���6��c����ھ�o侧}�mI�9�<�{Mܾ�=�'�=�7R�7����� ���b�b�F�B�.?<x$>[�ʾ��M��n-<sʾ#���p����ե��+̾ؗ1��!n��̟?w�A?�����V�4���_�\���Y�W?�M�Ļ��鬾 ��=ٱ�)z=�#�>0��=��⾢ 3�S��k0?�B?�2���C��~�*>5����=��+?Z�?k�;<* �>��$?�-��6�j�[>�B6>��>��>�>�K��dzؽH�?��T?�2 �������>�۾��{��eb=X7>I�5�lLؼ?�Z>U0l<�<���"S�Bp�����<C�N? ��>��+���6���]�#T���e׼9e?��Z?B� ?t}�?�Gl?�\�=����n��?�|aD��cn?7��?�5>�����4��*��M3?� h?�h>r���Gn����5�^޾ʤ�>t�~?��?�3*��ox�ƕ��4�6���;?��v?s^�ws�����?�V�a=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?0�;< �R��=�;?j\�>��O��>ƾ�z��������q=�"�>����ev����R,�c�8?۠�?���>��������=˽�����?#�?�٬��[p<�%�m�����+�<4)�=$����.�]��j`7�Y0ž��	�d՛����'>�>�@[����>3q8��x� wϿR䆿ÈѾK�v���?�*�>s,˽HТ�Նh��;r���F�i�H�H���N�>��>ܪ���򑾖�{��r;��ß���>�K�� �>��S��)��~���V�5<��>���>з�>q6���佾ř?Y��TAο穞������X?(e�?m�?Xl?9<~�v�R�{�y��0G?�s?�Z?��%��E]�b�7��j?L\���T`���4��FE��U>K"3?B�>�-�ݼ|=�#>���>gl>�#/���Ŀ�ٶ�,���;��?���?<n�N��>���?qr+?�i��6��mY����*���/�K<A?2>،��V�!��.=��ђ���
?�~0?���.��Z?ي;���V�uVľ���� �������@�,FʾD�!�V�c����@ɽ��?j��?�X�?K��j���H?tY�>��l�6��!��Pޢ>}�>�#�>��=��>���y4ӾM;ƽ���?��?g;�>�ʋ�鷌��J�>��l?�r�>��?���=�\�>}h>�В��.�'�->�v�=..G<�N?��\?�~?8K�=�,��`���J�Gz�rm:��4?�,m>�+q?R�w?��>�~���<����`��ɳ���6<g�m����=��x >�1>��= 0｛�'���?Kp�8�ؿ j��p'��54?/��>�?����t�f���;_?Rz�>�6� ,���%���B�_��?�G�?>�?��׾�R̼�>:�>�I�>=�Խ����]�����7>0�B?[��D��s�o�x�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*׋ֿُ������Nި��ɼjԸ=��>�B��=���=.�l<�Z�,�=�i^>��C>��?>���>�)J>�`">~���[: �p9�����|aX���*��n���Q���������@Ͼ�sǾ�;�qٽ���<sl7�]MN���);y��=exT?e�a?V�g?�?Mu=90�=��ܾ�F&���罯�>�%�>�1?��,?�?�h������r�6V��%������h?\�x>g��>�?�>C;¼�L>��>�>�A�:uD��$��:�m=��=�Q�>��?�c�>�C<>��>Fϴ��1��k�h��
w�s̽1�?���S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW? �>!��x�T�4:>8����j�4`>�+ �}l���)��%Q>wl?��f>au>D�3�E^8�\�P�����#|>,26?�ζ�[j9�6�u�9�H�m�ݾ>;M>�ھ>@F?�WZ�a�����lwi���{=fp:?��?�Ͳ�ڰ�n�u�g��[R>&\>�k=c��=T4M>ؼd��ǽj�G���.=���=f�^>U?��+>��=\�>S9���iP����>�oB>��+>�@?%?�^��旽����� .��0w>�k�>e
�>�<>`^J���=Y��>��a>�������w���?��W>�I}���_��Ov��4y=�7���x�=|��=HL ��<�g�%=��?|���3,���Ǿ�,ؽJO)?X��>�S��<�L>�)���h���p��?
�@V�?��ᾭ�_�u�"?VB�?:�����=q��>؝l>}���-��o?0�#=�-<��松�u�?M�?4�<B+����f�x�=�%?n,��rh�>fw�mZ�����4�u�F�#=��>�8H?	V����O�>�*w
??_�驤���ȿ||v����>`�?���?N�m�gA���@�^��>��?�gY?yni>.h۾K`Z����>��@?�R?�>�9�K�'�Y�?�޶?���?�I>���?�s?�_�>s
x�X/��4��~���ˆ=1�\;�j�>�c>�����gF��ؓ�ti����j�����a>6�$=��>YA佱4���-�=拽�D��g�f�s��>;+q>��I>T�>�� ?�b�>���>	�=Le���耾캖��SE?�)�?�z��#z��ٻ"�2>���k?�B?%@�=
��?��>��s?dZn?��3?rM>�l� á��BɿX��E�Ѽ�B?> |?�j�>�h��B>+D뾉l�7�>���>�8�:F �b�A�'2">U�>d?���>z�;nO?�L'?��?>_��>c�<�9t���rB����>J��>�H?ڪ�?�[?`5��&�7����%����R�k,�>�"z??�U�>�l��uϞ��Η��<������ւ?/er?�s���?*�?�V@?s�<?��U>�:'��[�嘽�%�>]#?���C���$��Y���?�U?^��>R��1���$�w����?m�]?y^$?�@��[�ߓ��32�<�J��ku	�V���:���U>E�>�yc�_�=�#>�R�=�6h� J�Aw�;Zߺ=��>�#�=��:��{��.:,?��D�p����=��r�>vD��]>�iL>�����^?�=�3�{�����r��)�T��?���?[�?�V��<�h��)=?��?�?�/�>�D���޾���V�w��x��|�܏>��>�o�H\徘���X���5��1�Ž�����>#J�>��?'�?��8>�	�>N��26+��l��	�aLa�����i9��P/��Y�s���Z�!'������z�"��>.Q�����>r,?�k>
c|>�>�΀���> C>w�z>i0�>��F>}h>1>e�<��ƽD�V?����B�0����y���L�<?a`?`��> �ż�;������}?`��?wt�?���>�rX���.�F 	?x�
?�t����?��h<�z��1���vG�� 9 ���T������>�ٽ+�,��_�����"o?qO?���=M}׾	U����7�n=N�?��(?�)���Q���o�θW�S�6���6h�Mj��Q�$� �p��쏿�^��%����(��r*=��*?j�?ь����!���&k��?��df>`�>`$�>-�>#uI>��	�s�1�h^�M'�K���hR�>[{?�=�>G�I?J9<?orP?ŒL?� �>��>�毾h�>U��;
�>V,�>�9?0r-?.�/?��?V�*?�.`>G���������ؾ7�?S�?�?�c?Q?JÅ�-�½�5����d��5{�,�����=�s�<��ڽU�j�t5\=��S>&�?�8��1�� ��<�>�l.?���>.>�>�"M�s�B��>�h�>�(?��]>GJ�b~���63�v��>���?�Ё�^8E:~A>�jl=I?��k�Q=;B>U��fa���<�#X��Ņ����=��=@h��x�=��=A)�nႽ�~�>��1?1R�=���>��U>	�B��^����F>�i:�ۭU>l��=��Ͼ��r�j���w|p��i�=�ƛ?�~�?-u�=�/>:L>�I�V��%'�H�_�s_���?u?]x[?��?oy�?�Y�>Q��<g־PG��"���%W���O?t!,?��>�����ʾ��׉3�؝?c[?�<a����;)��¾�Խ��>�[/�X/~����9D��񅻿��;��5��?鿝?�A�V�6��x�ڿ���[����C?�!�>�X�>��>T�)���g�w%��1;>���>gR?�#�>T�O?�<{?��[?�hT>ʜ8�.1���ә�cR3��!>@?ٱ�?��?,y?�t�>��>��)�h��T�������"����W=
Z>>�)�>�>���==�ǽ�X����>�_�=/�b>Q��>���>��>m�w>�N�<^�G?_�>�K��dϾ�4��)���2?��y�t?ޫ�?��>4Խ�G�X���*�KN
?lU�?Ky�?j`�>)���n6=��4=Թ��O�=I�>�Ϻ>v��=V�l>�#�=g�=�޽>�#�>f�ڽCh8��CV�� =�i?�L&?[0=��ȿ�q�[aؽ�T�u�=�-���k�~V�<4�:�Ê�=�s���-�/���M�4��P2������E,��q󔾻M�>�м=��=�A>°>�&�7�%=�VN=�5�<9XZ=���7�<�S㼯�D�3�Ƚ�mK�ԧX=:T�<����!���h?��}?F::?.3?W!�>t�>�ᑼF-�>��*>V�!?*Q�>���v���_��X]Ⱦ;�[�����`���h�����h�@>��=^�}=I��=oz�>E�=���=�j9>1Z�='2=fB>��q=��>>���=��	>�v�>���=e6w? ��������3Q��_罃�:?76�>�n�=Ăƾ#@?��>>�2������b�
.?}��?�T�?��?Gsi��e�>��3����p�=ٰ��'92>���=��2�c��>$�J>���J���}���4�?ӆ@_�??�ዿ��Ͽ�a/>��7>�$>��R�/n1�'u\�y�b�a[���!?�#;�j̾�
�>���=�o߾G�ƾ��/=7>
�c=�z�LO\�l��=^z���;= n=���>�
D>%?�=Pޯ�G��=��H=���=��O>�6����8�M.���3=���=n�b> &>��>!�? `0?�Wd?=5�>�n��Ͼ�>���H�>��=@C�>Zׅ=lB>���>��7?�D?��K?J��>���=@�>��>��,�R�m�7k��̧��m�<藈?:Ά?%Ѹ>��Q<h�A�y���h>�3Ž�v?�S1?;k?��>�c�\�׿��ݾ�#���ޤn�?c�=�퀽�	ս�Ñ<c	�w�U�9+>�O�>Fs�>EƸ>�f�>��A>�ɳ>�?>�َ<�<�/<2n>���=�>=�[T�#��>@]=��Ҽ[SA�[�=;�<nE�|d����=����A�=Y!�>�v>��>"��=]k��0>/���^�L��K�=� ���EB�Jd�[N~��.�x5��D>[X>����b����?�_[>7?>�t�?/�t?T�!>!����־��f�`�T���=�4>7>���;� �_��pM��#Ҿh��>`ߎ>�>O�l>�,�F#?���w=��Wb5���>�|��s��
)��9q�&@������ti��gҺ��D?�F��^��=o"~?��I?Z�?��>���҆ؾ	;0>�H��W�=n�m*q��h����?'?��>�쾩�D��H̾N���޷>�@I�2�O���U�0���0ͷ�6��>������оm$3��g��������B��Lr�\��>&�O?��?^:b��W��KUO����a(���q?�|g?.�>�J?�@?
&��z�r���v�=�n?̳�?T=�?y>�
�=<(��v�>�m	?֤�?Ǒ?A�s?5�<���>�F�;~�!>�a���L�=�I>��=���=B4?�
?�
?�l��<�	�� ��o񾒘]�6�<�2�=��>Mc�>�Tq>���=yie=Mޠ=O�Z>T|�>�*�>��e>��>dw�>��徻r.��(?�6>N�F>�jE?kd�>��y=���>��r��=��˒���������"�c"�;|oJ>q�K�K/?�sѿ��?��4>V��?Nt����7ma>2�>z�&��>��>�`w>�s�>�1�>�>Bc>�A>�FӾ`>����d!��,C�]�R���Ѿ�}z>�����	&����w��ZBI��n��wg��j�P.��Z<=��˽</H�?����!�k��)����T�?�[�>�6?�ڌ������>���>�Ǎ>�J��k���\ȍ�	hᾦ�?H��?,u>��a>�JU?��?x9��hMs���n��3����K�>�o���o�M�������-.���u��p?�Ye?�� ?z��<�ֺ>\�?�Z^���o���>/PT�!cM�$K���>�׾��@�8�޾�飾��}<�?���?�S?َ�>���ٽ�C�<�cj?%!T?7V?��P?�p?��=w�?��>� 5?8�?��?�!?z��>C1^=�>Z�=�����O���T� ]���нd��:-�r=Wy=[��=��J=�"�<��˽��ǽB������ML=TQ=�<�=$C�=���>��W?2��>���>��_?�����O߾2��;3�>��=� ��G澴(��\��W��;E�a?NB�?ٯD?D}�=]�K�:>��Ǘ>abo>j�m>i6�=���>����L��Z��=.��=N_;��Ͳ=꺕��λ���%����c9.>�J#>t[�>��>ݾ{�th�>O�Qv����=����gr��Ԭ��-K�v�2�����\?@>�J)?��A?�ik>jtӾ��$�~�Z��2?�\G?� ;?��{?�K��f�^��eQ�3`m���=^Y =�l���7������r����F�W_�=��>�Ɏ��ݠ��Yb>E��"v޾��n�!J�����FM=<��dV=@�2�վ�3�9��=
"
>D����� �@���֪��0J?�j=Kw���_U�o��\�>t��>�ޮ>�:���v���@�e���[5�=h��>;>�S��1��9~G�t8�f>�>XQE?�V_?!k�?"!��~s���B�,����d���
ȼ��?3w�>�g?GB>4�=�����K�d�pG�~�>���>R���G�o;��Q0��g�$�F��>�9?��>��?��R?2�
?�`?^*?�D?('�>������� B&?6��?��=��Խ�T�� 9�JF����>|�)?�B�ܹ�>P�?�?��&?
�Q?�?��>� ��C@��>�Y�>��W��b��?�_>��J?ؚ�>r=Y?�ԃ?y�=>]�5��颾�֩��U�=�>��2?6#?O�?�>���>���ZV�=s�>vc?[A�?W%p?�S�=W�?W2>�E�>,��=��>���>f�?��N?X�s?z�J?��>�_�<,���Ÿ�)�p���I��x�;{�><��r=���-t�#���<=��;�滼`_{�?��s.G��H����;N��>ه5>�׾P��<��|S���%>?g�=Λ��<~Ӿ2ϗ�6�ɽ+c>��?I��>-��<�6�<���>lu�>`��V�?�k�>l?������r�&4�&wϽ9�(>��?�P>�</�_�����=D>o��? �v?#��~����R?�|?���}Ӂ�xb�����x�a!/?ۚ?x`5�A��>��?��V?��>���ƅ�H젿�_u���X��L`='�>�̾~�9�P��>��?��>+��=�]�=m��S?w�9˾�k?�b�?,	�?荑?\�>�S{�����w���tm?���>�⾚�)?�6��/L���@���Jw���E����b� �X�SH������T��#ҽ4J:<"[?�:o?��]?�	U?��;[��m{�;��LY�~ ��u+� G[��Hm�bp �b�#������Pž󍍾�� �^�/�A����?�'?�~0����>�䘾�*�<5; �B>����(��=�ߋ��@=�d[=�>h��q.�J\���7 ?��>���>�<?!�[��I>�~�1�'�7�X����2>���>�1�>�>�W�:��,�C���ɾׄ��Oӽ �s>kc?�K?O�m?�����c0��5��� ��!�����C>&.> ��>�2Y����}�%���=�e�r�.|��吾�?	��{�=j�2?a(}>���>��?�?�]�n�=gu�Hb2�?e<a�>K*h?_��>�N�>�|ɽ"���B�>�q?���>�J>Rrp�"c�!�y����z?�>_��>$�?gC�>��#�#�Y��[��3��$�J����=O,q?�߇�ڛ6�E)j>a�6?���<����->�>*%�A�#�k��g�3���>��?��=� >�/���%��ʇ��c���L)?�O?��*��X~>� "?8[�>9$�>e,�?f3�>�iþm�2��?��^?�3J?GA?\5�>��=n}���`Ƚ��&�:-=���>}[>s�l=�6�=����|\�����D=�=tμP�����<˩���lK<!��<(4>Bmۿ�MK�"�پ
����4
��刾Ծ���e������c����d]x�����&��V��1c�����Ƴl�ʈ�?0�?�b��+��-���u����������>_�q��Q��	�����5����j���a!���O��i��e���'?������ǿw���AAܾ8 ?? ? y?/��"�y�8�Y� >D��<�W����뾔���M�ο	���w�^?���>:	�KD�����>��>"�X>�Lq>���ޞ�y��<��?Y�-?��>r�r���ɿ����y�<&��?
�@�|A?��(����F�U=���>��	?�?>�R1��H�����4T�>H<�?���?�wM=��W���	�e?s=<R�F�N�ݻ��=�>�=gN=�����J>�T�>t���SA�[?ܽE�4>�؅>"z"�/��(�^�Ԓ�<��]>��ս	@����?�W���i�q`-����A��=~�H?۱�>�{=e�?��H���̿�&Y��R_?�m�?��?��$?��ž�3�>]׾�#J?��/?�>~s(�w�w�Gw=C_8��漌��1�L��y>��>Ř�= ����o��}=U��=v�� �ƿ\� ����B�<ۯ�;n�B�ő��!��#o����}fq�P���jb=b��=Y�P>-R�>WDP>�V>�Z?��\?���>Rp>�"�3�}�i�оzZ�Z/~��z�%��__�_���4���iྑ�	�<�nY�)nƾO=�	�=;8R������� ���b���F�U�.?)r$>@�ʾ �M� �,<�oʾ�����Y���¥�p,̾��1�mn��˟?��A?����V�� ����{���ɮW?�W�����款���=�
���K=�&�>?��=����!3�N}S�h?0?/k?�k��������+>�q ���
=�+?Jg?�>b<�>�G%?�)�R��̑Z>OB3>fg�>Y��>�>3��h۽q�?��T?|� ������>�ཾ�lz�j\=M�><�3������Y>���<����AO�����+W�<d;[?4^�>�d)���3�.����=��!�}q�?��7?�i?�Is?��Y?wd��R�C�h� sN�u��s�~?��y?�@�=��t=�Ѿ����m?�L?��->V=���e���F��&�� ?t�v?�?A��<с�筵�>�4�MuI?��v?s^�xs�����L�V�e=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?m�;<��V��=�;?l\�> �O��>ƾ�z������0�q=�"�>���ev����R,�e�8?ݠ�?���>��������=�����?���?�ά���e<?��m�U� ��b�<V��=U-�#�I�u��7�6��ľY%
�$�����Ӽ�A�>��@�6���n�>vY5�Y��ckϿ݆�a9Ҿ"&y�m?���>��̽�ۡ���f�*r�҇G�S%I��Ŋ�R�>Z�>�Δ�h�����{�@v;��r����>00���>��S�F.�����7<��>���>���>����ؽ�+ę?�]���?ο9��������X?�f�?
o�?Ys?G:<�v���{�����/G?Z�s?mZ?Б%�r"]���7�3�j?6F��V`���4��>E�U>�3?pE�>:�-��}=�/>H��>�b>�#/�'�Ŀ�ݶ��������?g��?cn�0��>6{�?�d+?�a��5���K��m�*���C�L.A?F�1>y���Ѳ!�,=��Ւ���
?u0?���i3��\Y?��S�fPn�����Y��Jv��V~�uA����&)��{�S����3%�0�?0o�?G��?@㟾��9 ??�9�>�V�#g�R�U��!">�+�=�w�>J��>=��>Z� ��-��9$=�?�2�?)��>9'���0��\��>�̕?���>)��?��)=46>Eu�>�-4�֜}�<�=d{6>�z�="T�>��T?0�?-n�<s`���4��e1��h���-��R5��>Svg?]Ht?r�>0%��y��rݾ7�����TT=�Y ��^>js`��'7>�V>��>��ʽBAU���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>B�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?* �뿔����(��FǾ�Z;��^�>�+�]�X=�[!=b�=߄C<a3>ph|>��>W,>���>.l>
��=�Ӏ�,� �����0>��g%2��E�s���[����eo����q��E��������Ľ.���tg�8�A�hֽ�J�=h�U?��N?�:[?�?�8�s�=�^Ѿ���=���=��>��M?m'?t?+=�ʑ��1a��܂�=p��c�h��?�p�>��>f�>2��>GA[=tpo>T>4A�>�I����WǼ���<+�>���>��>���>�C<>��>Eϴ��1��q�h�w��̽/�?����]�J��1���9��Ԧ��'i�=Vb.?b|>���
?пY����2H?���t)�x�+�e�>b�0?�cW?3�>-���T�>:>��ަj��_>�+ �;l���)�W%Q>nl?sao>`�o>>�5�46�6sS��f��Q m>��7?���B�N�QSu�+�H���ݾY�P>��>��Z<���m��!y���g���=�h8?T�	?�M���ж��v��Mݙ��4F>�S>�"=zz�=KS:>����������=���=���=��\>;U?g93>Oݎ=?H�>�m��OsZ�V��>� @>pc>\'>?�P?�_�����͉�&R4�eF�>$�>L{>J>q�F��E�=���>q�`>;y�(약�{�/3B��%P>+�e�n�Z��~�y��=r����=g�=>���01�%(=\v�?��?Ɠ�!��D�Ⱦ�O�>��>-?�Ja�=EF�V��y>��b�?z1@���?�� 0|��^?�0�?{���`�>,�>(C�>�C|���>�?-��>K�
,��p��H�?�K�?��=�IW�#ve�q~<�6?piξXh�>`x��Z�������u�S�#=@��>�8H?�V����O�[>��v
?�?�^�ީ����ȿ<|v����>Y�?���?\�m��A���@����>5��?�gY?]oi>�g۾E`Z����>̻@?�R?	�>�9���'�{�?�޶?ϯ�?nI>΍�?7�s?id�>x��X/�6��때�`z=c�\;@f�>^`>m���QgF�Eؓ�Ai���j������a>]�$=Q�>�A�n4��9�=l���F��d�f�_��>c'q>�I>VW�>`� ?�`�>���>h�=�g���怾}���
�E?�5�?���ˀ��P�=��=u׈�.��><I1?�G�=:������>�LV?Śm?%_9?uY>�~	��>���aſq8��prJ�Y�_>�?���>)��a�=�ھ��[�9X�>O�L>�����ϾPMN�4Բ=�l�>2>?p|�>��=e� ?��#?�j>@�>�^E��6����E�P��>���>�K?��~?��?�չ��Z3�n	��l衿>�[�GN>K�x?S?6˕>���Ã���E�CI�~璽���?�ng?�X��?C1�?�??�A?� f>p���ؾ1ۭ��>�"?�A��6B��Z&�]��j?"�?���>�Ҕ���߽�_��c�f���\?O�\?j�&?�<��`�������<+��������M<=ez��/>�>�3��|7�=u�>Z�=8Nh���:����;�?�=^h�>�[�=-';��ې��,?^A:��΃�ݟ�=;lr��rD��%�>�=L>#����q^?��>�|�k���x���+U�#��?e��?}(�?�i��`h��=?S�?p�?���>sT��xUݾ�ཱྀ�w��x����ds>�`�>�\w���S��w��l�����Ža����>�e�>n?�u�>�
">4ʾ>����E5�f�D���/e���bX=�:/�Cv
��~�M�&�����t����f�q;�>��|�8j�>�r�>�m>bIf>+��>7(<���>7qG>���>�Ü>l�>�I7>d��=��=shĽ'$^?^.ľ26�.�d�Ӿ��4?�	_?27�>z?�<���7Z!�8�>�Q�?^��?�e�>�:N��sC�8Q?-�$?�~����?���=|��.<�=뾾<ս��<�}���Ra>��~���&�� Q�z?Ծx�?��3?|&&>�l��C����<�n=N�?��(?�)���Q���o�θW�S�4���6h�Mj��Q�$� �p��쏿�^��%����(��r*=��*?j�?ь����!���&k��?��df>`�>`$�>-�>#uI>��	�s�1�h^�M'�K���hR�>[{?��>��I?i�<?��N?�5N?���>��><�����>^�,<���>E��>|,<?��)?��+?�d?~`)?��X>-�]�����վj�?�B?{?�m?��?�まoѷ�Y���bꄻL솾�)��#�~=;�<�ཁXb�gtp=�_X>L�?]�x�8�Ӄ���h>{i7?�h�>4��>�P��������<���>�,?�^�>�����fr�����_�>sƂ? �C�	=f�*>� �=�yj�؞9��0�=s.��Yx�=Q�����;���<&�=��=�iH��U�:��A;���:1��<�S?��5?M��=�i�>Ȁ��D�����d>�=P>*,�>z7�=�!��x���ϙ�1k��Y�z>ό�?���?��μ��]>%B	>�̾����7�p6ż� ����?�c�?�&g?+��?��z?�T�>�R>4�־�����8h��ˮ=�?�!,?y��>���8�ʾ򨿈�3�C�?�\?<a�����;)�#�¾ս�>]W/�O*~�6��~D�H�����=w����?���?�"A��6��z辌����\����C?A!�>d]�>��>��)�u�g��#�q=;>j��>!R?�!�>|�O?+;{?Ѥ[?�tT>��8�"1���ҙ��	3���!>z@?o��?��?�y?�p�>k�>j�)���W�������Zڂ�00W=�Z>⏒>H*�>?�>���=VȽ�V����>�vj�=��b>	��>���>��>5�w>�C�<�G?8��>
���fg�d4���6���;��3u?�s�?Gn*?��=!����E��i��Q�>�|�?��?H)?4@R����=B�ȼ����n�m�ȕ�>���>+��>�=��B=xC>I��>���>� �4��p�8��xJ��?W|E?M��=|�ȿN�t��g��@���6<?���n�Y�Μ���_��s�=�Z��Q�훥���V�6̙�=t������o噾+	t�@C?,��<0>cʻ=�3�;(��U��;�f=�(�<��p='ؾ�#�<b�L�;�Ǟ��J���$<l�#=���_��[?ANs?3`5?�3N?ȵ>���>y�d=>��>��r=�/?3�>��>jG��8\�帾�fH��鷾=���g?�c���� ;>���=c��<`�E>�Os>bˠ���=1��=�)=>���Q���$�>�,,>�x=�w�=p�L>�� >5w?˚������1Q�ds�^�:?�)�>�(�=!�ƾ#@?��>>O3������_�p/?���?@R�?x�?�si�i�>��1��v�=����&2>N��=~�2�S��>ҽJ>����I���]��)4�?�@_�??�ዿ��Ͽ�o/>_�7>��>FKR��0�³[�d5d�XX��?!?��;��˾JE�>N!�=Z=߾�hǾ��(='�8>�n=P���[����=0�w���A=��n=2�>үA>��=�u����=Y3L=t��=��N>?�5��\:�	�7��b6=���=5�c>�&>,~�>�?�;0?�td?�^�>9Zo�&ξ���(�>d�= ��>y(�='B>`��>�x7?�D?nL?bx�>� �=�	�>s�>�,��m�<�ধ����<���?��?���>%Hq<<n?�`���3>�v�ƽ�(?�61?��?z��>���wݿ���'��I~���<�rl=��x�j둽T���� �z�����=���>-��>�ơ>zLa>�+>��=>WS�>n��= >s=��=ٛ�*�*=LPͼ/<�=7'��| a=B�����s<5{��ü���^pF��8Իs��L�<;!/�=�>lr>]\�>И�=�G��h�/>�S���6M���=���lB�!Wd�&a~���.�Pw4�slE>�V>4#�����f�?Z|[>�?>7�?��t?�z">��r־	 ��;�f��UU�%��=�	>-�@��;�g)`�&M�FZҾ���>�ߎ>�>I�l>�,��"?�>�w==�b5���>>|��ƺ��(��9q�2@��#����i��uҺ�D?�F��>��=)"~?��I?B�?n��>���:�ؾz:0>,I��n�=9�	*q��h����? '?���>����D�tH̾����޷>Q@I��O���@�0�!��[ͷ�;��>������оg$3��g������ӍB�uLr�Z��>�O?��?::b��W��IUO����O(���q?�|g?i�>�J?�@?%��z�}r��qv�= �n?���?Q=�?b>�
�=[ص���>	H	?���?`?�s?.?�'n�>�;G�!>ؖ����=�>p�=BY�=`?ڒ
?��
?�̜���	���𾻊��]����<��=���>L�>=Ar>PG�=U�h=�:�=I�[>	Ǟ>܏>S�c>x
�>J�>d�Ծ3� �Am$?f��=-�w>�2?��z>q{0=K�½���<򛇽}�:��2-�������Ͻ�(�<O��S�#=^���y�?��˿���?N�>>�z��?�o�o���sG>J�w>)!S� ��>/�>��> t�>NÈ>˰>��>�>�DӾ�|>l��e!�6-C�Q�R���ѾXxz>ɜ���&�w��k~���>I�Rk��ef��
j�R.��N;=����<�G�?����2�k�6�)�\����?h\�>b6? ،�s��*�>��>Nȍ>�H��P����ȍ�8h�
�?��?v/k>��9>6�K?%Z?꩐�4hR�g�o�����.�Z���f�x�e� ���%���U��؛<��f?��_?�x?��N��>v��?�c��Q�Yˤ>��^��J��^��W:>$��;�Q�[H���"����>�!�?��T?'��>�a���Ԭ�����}?��S?�^?�h`?\�{?���<c ?K`�>�aT?'� ?���>�}r>�{�>BU�<G�>�T >V뀾�����������F��͕Խֵ�=Hy�=��~�2������������=w�ý���<+}�=纝=
�����=��>co�>��Y?|�>��>�)?Xwy�;��\Ϙ�E��>z�p=�}ʾ��־D��������#=�<q?���?=S8?�33>�%��c�J!\>��~>+R)>N��=���>z)��W�S��=u?�=���=�$2>Ԑ��:�о�U���_�=K�>,� ?B��>�������>�yƾ�Z�;�<4�<Z��ǯ���T�i�-��Z���1>�d?�eL?��>gC*����<�G��6?@�J?�wV?e�?k��=�Y�R�5��:P�㴋>+/�=t9��+��T�������Y+���|>�_U>��ʾg��;_>� �Gݾ+l�ˤH�˰���]=����T=���׾ʹ���=#>�Y���� ����������J?�9k=�����N�X���b�>��>�#�>Jx8�=L��ܒ?��̬���=���>��7>,`Ѽ�(�]�G�*�>c�>QlF?#�H?u?޼[�����äA������z��f�����/?��>��?��I>S�,>8�������k�=�_�oa�>���>Yo	��B5���w��~ƾ����,>���>�6>��?Dm?d?;�A?R�?�y.?���>��t<�`߾�%?#ل?&Y=�\	�n	��
G�j4� ��>)�?�r�Y��>cSa?�h@?��	?HKC?�� ?�;�=����wo��m�>���>4�C�
�ƿݶ��� �?��?�pp?��r?W�꼨�C�fՉ�oF=��Q>j�'��r?�_(?�1?�0?A�?$ 6�FDD�$G>��@?�c?^z^?�Q<>̝D?��>�G>��m�ut�>TZ?4�?�V?P�_?��H?�/?8=�=ZL=�� =>{�;V$�=��ż��$�z�=�e�P��<��< �=e��=��D=E#��r��<�\ļ���-G����>�Ct>R��\0>P�ľlD���:B>
[���C��ݤ��*�;��/�=2��>V�?� �>� #�R�=��>J��>����i'?2�?2E?m0I;c�a��gھ�L��n�>��A?Sp�=2�l��a���^u���d=L�m?x0^?��V�����kb?D3^?iW񾜩;��9ƾ�lh�����N?Hd
?� L�V}�>D�~?�q?t��>r�g���m��B��c���h��^�=�ך>s;��9d�׀�>^x6?�e�>6(f>���=��ھ��w�#���?ꐍ?���?r��?�\.>��o�`7�����o��P�2?fe?�5�C�?� �=���>Kj��;�� ���J;ɾ���f����h���
�����~�]�6��:�?/]b?;�X?�ql?b��n����v��Tv�Bq�č<�����@�+�Y�|����D�M�B�0����n]<�\M��1�ߤ�?>�-?�򯻅��>)�Q�����Ƥy��Qt>n̋���̽��i=��v���^=lo�= SN�eO3�����S�!?���>g�>�Q@?�A�1�=�h�%��M,�;k��Z9>�6�>�>=��>X)�=Np�tv;�����wHp��Ƈ�w��>I�g?�l3?��b?Lyžr�k�����m� �+��%߾���>�@h>+�>����^��� ���Z��8���F�9l��������/?���>]� >���?o?��,�3��Ã�.��R>�<��#?��?}�>�?Na�.\����>!�l?�+�> r�>�؍�b�!�jY|��̽�M�>��>���>�Vq>b�+�ӑ\�����z���9���=ٜh?|I����`����>F�Q?#" ;��8<6�>�dn��!�P��կ'�(�>�?Ԑ�=��>>��þE��*|����~7?l�?h��6��jM9>��4?gf?ɀ�>:Ly?���>)����o�j��>n�H?{�J?�,F?qX�>'b>4]���>��q�N��h�<\d>�.>�ү=Tw�=N6��)��Z��^s<�Ѽb��o"��DI�!=�l�=�f�=�U>Pۿ>K�tRپ���K�
������]��|.��w���*��@���qy�2��,&��U��Fc�9M��2�l��T�?g�?���"���%q���F��;M��S�>ـq�z���Pq����g1��A��қ���!��P�9i���e�Y�'?������ǿװ���:ܾA! ?B ?�y?���"���8��� >�I�<,��\��p�����ο����w�^?&��>l��0�����>.��>l�X>WHq>/��J瞾7�<��?��-?
��>I�r��ɿJ���ʿ�<���?��@��A?$r%�7�naH=���>C�	?ߙB>��)�[/�򋭾��>F.�?�R�?'~|=��T���"�c?#g1<��D��ˑ��=�ʤ=9�=���N�L>�S�>�L#�T�M�ecýg9>�v�>x+��m�cqY�vo�<(mW>��ٽPؕ� Մ?�z\�tf���/��T���U>��T?J+�>f>�=��,?P7H�=}Ͽѯ\��*a?�0�?ۦ�?;�(?.ڿ�8ٚ>4�ܾa�M?D6?u��>�d&���t����=�;�ߣ��`��|&V����=V��>%�>��,������O��E��U��=���.���.�vG%>Fx���	ὧ���{K���e'��2��ξ)��<��=���>�G�>d��>^�>[_8?5Cn?K�?��6>��<ՐM���h�y=v��ǀ}�x\��౾AZ�����E��O�����U�[S�qB+���=���=}&P�(��e����_�=E�#.?F�#>VR˾c�Q��1�\9ϾCB��tS��⤦��d̾�/��n��8�?�ZB?T�����S�ߢ�����F��q_Y?�O��z[�	6��Ȭ�=H���2��<D�>��=��ᾣe4�q�S���0?��?��ɾ.��i�=�����#>�:)?`��>�y�<�x>G�'?�򽱺��p�>�^->x�>��>{�=�u��F�W�[�?_�[?�l��2q��(�>w�Ӿ���;�=�vw=��W�O��<:h>����-ߚ�t�лi��=��=s�U?3U�>��$�-��꥾N ~�n�e=f�?hq�>��p>�$W?�O?5�=��þxoE�!��t�=׎M?�NU?��>٬���+پp&��W?�r?t�w>��h����6�}G����>��\?.4-?�̸�;��yD���@�ʂ8?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������f��=�\�]~�?}�?K���U�E�S8��2�aو��_(>JMH�I�߾��׾p� �*�v	(�Y�����[���>R|@==�>���>O���!Ͽ��Bp�����f&����?E+�>�=�����]���i��w��K��E���P�>��>����h����{�mo;��"��}�>���i��>ǶS�r��[�����5<��>0��>���>x/�����?�^���=ο�������6�X?Rh�?^o�?�m?��8<!�v��{��W��0G?�s? Z?rF%�(]�+A7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.���_?��a���p���-�<�ƽ�ܡ>�0��\\�h�������We�x���9y���?�\�?��?î���"�6%?n�>-����2Ǿ�3�<,��>�%�>�"N>�L_��u> �p�:��{	>M��?�}�?�i?{�������:U>��}?�;�> ڄ?���=u�>2,�=<`����f�ν">^�=G�F�n�?�rM?���>h�=� 1�>j/�-EF��S��	��rB����>��_?`L?A�o>9���%H)��� ��ڽn7)�Ke���3��;�H�ֽW:>��?>��>��9�jվ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*�[ҿ�Ƣ�����|�>=t��<�.!>�-����ͦ<u(_�n�%��=��n>��B>OH�>ߝ�>b�>��e>����,)��B���{���V,��R!�\~�u'���90��Q�����y� ������P����<F��=Y]���>.&�=��S?��M?x	o?��>�倽�$>e�����<* �+�=��>
/?��K?��+?*\�=������d��g�������ʈ�ț�>u�S>3��>�`�>���>���޼B>�J>���>�>��	=j��ew!=�bV>�ƭ>�=�>���>
I<>�>�ʹ��1��D�h��w��̽4�?*���w�J�40��K/������:v�=Qa.?N{>���<п)����0H?����x)��+�3�>��0?�cW?��>m��0�T��.>����j��g>�- ���l��)��)Q>�m?�mg>��v>�"3�F8�e�O�L+��KH>Lf6?}����9�|^u��.G���ܾicL>b�>�kA�ƴ�����~�k�h�y�k=x{9?�+? ÷�F����"s��Y����U>��]>d�=�L�=s�N>�m�vyʽ�KI�`+= �=~�^>��?�#>�y=��>c���&,+��²>��[>��Z>��B?�3?w+����ְw�/��g�>���>���>,C>R49����=�c�>lIx>��߻r�����PG�`(<>DG�:�w������=�]��0��=!�P=�|
�K�.�)݉=�~?���'䈿��e���lD?S+?a �=z�F<��"�D ���H��F�?q�@m�?��	�ۢV�A�?�@�?��P��=}�>
׫>�ξ�L��?��Ž:Ǣ�Ĕ	�$)#�hS�?��?��/�Zʋ�=l�y6>�^%?��Ӿgh�>�w�xZ�������u��#=E��>�8H?�V��~�O�q>�w
?	?�^�̩����ȿ|v����>9�?���?S�m��A���@�%��>=��?�gY?Aoi>	h۾�_Z�e��>��@?�R?^�>�9���'���?�޶?ԯ�?�GR>&�?�А?a?o5߾K�Y ˿FK�������O߼�ؿ>Ή=��Ծ���;;���1��@ۆ�Z����.>�X�=Z��>v�X�X��C2��A/6������9�=�	?��>#��>GZ�>��?�$�>{)�>�(>�P=��<R�7�J?r��?���a{��=�z>�N�_?�+�>_A����ľ��>[?歉?ޭT?�t8>����a����h������Q">���>�[�>'�v����>J�ȾI���ـ>$֤>J��u����x�\(>��>�r?(�e>�D=TI?0?�C�>Æ�>(�h��옿��j�e�m>r�>�P�>��?�;!?�s���XY�[⚿���<s��>Q�n?�{?i��>�䒿`3N.=]p����.=Z��?��N?�����{?(��?o�C?��J?���>�{=�S�k4���v�>�$?79K� i>�5#.��޽��?f?�a�>01����("��Y~۾��⾥�?�hc?X%?���O�\��tѾ+��;@�T��l�;4�=��C��53>I�[>�Aܼ���=�|>���=�g�wMv�ȴ��}>N�>�=����1�>=,?��G�9ۃ���=��r��wD��>�JL>�����^?�l=���{�q���x��FU�� �?��?=k�?
��ӝh��$=?�?n	?�"�>K��~޾ �ྱPw�}x�w�(�>b��>+�l�i�6���䙪�qF��e�Žj��5��>���>�+�>��?�0�>8ɮ>"����7��y���E��8v���=���L���%�~Q��[��!�=���%�γ��B�4��>�>#@>Ʃ�>#��>0�>���>���>".�=zn�>H��>��h>�U�>���=�&�=� >�uD�L����Q?�᣾I'������⧾�|@?�_?P �>
*��=���.!	�j�'?׶�?��?Qfu>:8f���"�� ?���>��y���>NF =��8<��=�ğ�a���ѽ�ǩ��a�>&(ѽm�4�Y|L���2�f�?�o?S�޻�Dھ�޽f�z��/>�v�?>�]?l�=�=�^���l��fz������M�����,*�����r���ᢿ�\��b�]����?f�_?�!̾(o
�iξ"*>���X���2��D?Aq�>L�>T�m>7Vj�5�\�1��h8�ԛf��x�><t?��>��8?�O%?�J?��G?H�>���>�e���|�>��<w��>�>u2!?�,3?N.5?��?�F?�:>�+�����A߾�0&?��?��?A
?� ?��5e��uB=�=A����rȽQ[W=�|�<˛7��/Q��׼���>�?r���q8�q���1g>�s7?���>�]�>�ԏ��n���ý<J=�>��
?]�>�����#q���
��8�>���?Y�����<�7&>���=�\5��s;d�=����"�=�`�mB����;l��=
�=9]��%||�77;�R�;�<�u�>�?���>}D�>]<��g� �p��8s�=<Y>S>�>�Dپ�|���#��N�g��ay>~w�?z�?�f=� �=.��=�x��MQ��c�����:��<%�?�H#?�WT?Y��?H�=?5k#?��>*��L��_��L��j�?x!,?g��>���ͳʾ��s�3���?{[?�<a�����;)���¾v�Խ
�>D[/�/~����&D�������;������?㿝?�A��6��x�˿��[��d�C? !�>�X�>��>p�)�g�g��%�L1;>��>DR?�B�>K�O?�y?y�[?��R>:�;��g��)����s���z>�A?��?�(�?C~w?���>�#>^�-�W�����[.�������@V=Q�]>�N�>�q�>t�>�G�=����ɩ��-��`�=�)_>{�><��>@��>Y�}>�V9<pI?�l�>���1��m���YN�Nƃ�x�p?8	�?U?9?��=���W>�	�����>���?�c�?��*?�E����=�2��򥱾J%r��>�6�>܈�>�Nu=2�=���=O�>�2�>������}�2�5�G��'?��B?f��=�<����j�4�U��އ��ʷ=\9v�M�5��
�:^�5���=*设��C��dȾ!B���֣�`�����K����ꊾ�m ?4=V�=�>3>W��<�b8�4Ѓ=���=��*<���<\�3<��=`=��Is\<�q���I�hT���JA�"'���˾܍}?6:I?M�+?_�C?Ӿy>�A>�w3�V��>�����>?_V>W�P�����;��������ݵؾqx׾�c�$͟�oC>=8I�"�>;43>7M�=PL�<��=�$s=6ώ=��Q��=�)�=I�=�c�=���=��>�U>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=J����=2>s��=w�2�T��>��J>���K��D����4�?��@��??�ዿТϿ6a/>$�T>
B,>!�N�W�4��S�2�/�����x$?�A�vQϾ�p|>�`>.�Ҿ�������=}'7>^#u=p�/���W�T��=��½�8$=\��=[~^>׼M>���=�0����>6�q=R:�=��(>�n?���˽k28��f=��=���>�y->V?��?¨.?^F?v��>����1�F'���(�>��>�
�>��=� �>}-�>b;?o�N?��B?["�>�0�=�Ұ>7®>fH��As�}��1y�*��kjh?�5}?N��>dx�<�����x3�F�F�Ǣ8��?�2?O:?�Q>M�Cu��q�"M�\��=����=ؼjR��V��������|�[�>m%\>:�K>���>�?���>�$?�H�>�H�=aڌ=���=��B==W<������=�+�=���=��^=
�x=W�=y�E=U�$�������<碷<e��=bz�=��>��>�@�>�G�=�����.>�����4L��Q�=�몾��B� �d���~��.�EA6���@>}LX>���M����-?y�Z>b�A>OB�?v�u?э!>|��j�Ӿ�.����e�x{T���=�>��?�
�;���_��WN�44Ӿt��>�ߎ>,�>ǻl> ,�`#?���w=��b5���>)|������(��9q�@�������i�ڳҺ��D?yF��9��=�!~?�I?\�?���>���P�ؾ�:0>�H��
�=2�3*q��e���?7'?՗�>@쾖�D��G̾�����>D=I���O���J�0� ��ͷ����>������о�$3�h��~�����B�Qr���>��O?9�?�:b��W���TO����z(���p?�|g?U�>�K?�@?�%���y�Nr���q�=~�n?���?I=�?c>��>���a��>t-?���?��?x?���ȱ?�>��=L^�\�=-&>���=�:>� ?��>zz�>�sĽ,�K�	����:���n�ག���r�>���>���>VKc=m�̽��=��*>�m>���>�t>b��>�%u>�����t� ?L4>՘�>}1?I�>;��=��n��^= y��(�D��N�����w��=T�<�96����<�l`�_�>��ÿ!U�?!��>�K ��?�9پ�� �~�F>�`>ф���>�&3>JG�>c΢>5��>A/�=��u>_J&>#JӾ�g>���V!�nC��xR�إѾ�z>팜�?�%��������nI�bu��Wf�{j��+���==�q�<DF�?�����k���)�B��� �?yS�>n6?@⌾�Y����>���>w��>"0������xˍ�mq�x
�?���?�;c>��>6�W?�?��1��3��uZ��u�E(A�e�p�`��፿�����
�d���_?��x?'yA?%Q�<+:z>H��?��%�Wӏ��)�>�/�';�:B<=�+�>*��1�`���Ӿ��þ&8��HF>o�o?2%�?_Y?\TV�k���5�>�4?l,3?A�n?0�B?��F?.�
���?sP>�?�o?�T$?��+?I�?��I>B�=ң���=da½�Ɨ�L�F�9N̽�=a�	�>=-{1=��p=�=f�=+5������眼o�5�|�`��=�R=O��=->I��>&n]?��>���>^n7?�L���7��u��7/?F�B=�M��X���衾Y��{>�$k?�ӫ?��Z?"=e>Q+A��LB��V>|�>�%>P�[>A�> �d�E�aτ=�?>z�>q�=�R�-�����	��]���B�<��>��>;�|>`��x�&>�a��p�x��e>_�P�ɿ��!�S�t�G�rK1�sdu���>��K?�?!�=������b�e��(?<?�nM?�L?+��=Ч۾M�9�XJ�'�0�>�̤<1������8����:�O+:��u>k���� ���d>��
�v-�/�m�7�I�����=����<K=y
��Ͼ8s���=Jr
>7W��-��Sߖ�lm���/I?��l=�ɤ�I?T�'ۺ��>K՗>�t�>5�ƀo���?�� ��YN�=�P�>�<>
����n�gD�����,!>q�>?�cl?�}U?��������,��I�
��!Ծ���W4F?u��>�n?�>��)�|;���bN�����R��>տ>kW9��<��G徨�侨���R�>���>!��=�*�>Е2?�r5?/т?�#?P:#>�y�>8Ð=գt��Q
?X_w?5es�q��낔��-��3���>`�?U�09�>�+?��(?�F,?��D?��>�b3>@��8S��ӥ>�Ne>q0b��g��^�(>��G?���>rӎ?��}?Xؽ=��.�L���|�����b
>~�?��?M�5?	)?>?�Bq����=��>��d?ܻx?J?�"i=IF?�&�>���>�ほ�6�>���>6�>��=?�Km?��?�?>�6�[���?O��h��t�7+=<b�`=Y[�=��꼨��$�8����<˞>�
ƻ�\���q��94�����ȟQ;�9�>��>3r����>J�ɾy¬��e)>\�|��W���ᇾ7�*����=�l�> ��>GE�>Z=�#�=���>��>���'�?� �>��?��=��O������\� h�>��I?���=Y�l��@��o8z�}�=b!s?._?�gY�s���b?�]?Qw�.#=��þ��b�/���O?e�
?�G�
Գ>	�~?m�q?T��>ûe��Jn�'朿��a��Ij�a�=ѝ�>Pr�He�1r�>UW7?�k�>.�b>�O�=�rھZmw�����c?�ǌ?D�?:�?Vn*>
}n��/ 9����%?Э?s����,?���=�����M�h��f��d��oC�+ ���ž��]�<�S��!>��>`o(?&gD?�O?G�?�Z���9���>����g9���C�(��R���63���i��U�� ��9<�7����r�=~���B����?��(?y�1�ќ�>�h���)�L�;��?>\ߠ�����a�=�Ǜ��1=�V=\ k�{t+�%�� ?Tf�>���>t;<?x�Z��>���1��7�����;�/>�-�>۴�>Ɲ�>��I:vn-����7̾#?��yҽ&�P>��Z?�,?�N?�ꜾG(I�2�	`��=��oԾ})�>��>�Q�>��ཕ<��"U�JE��Pn�P�������#���!�=�??��>�Ӌ>tv�?\��>" ��1��1��q�
����=�'�>Zf?�\�>�3�>����g~�4��>k�l?^��>	�>0���KZ!���{��ʽ%�>߭>?��>��o>/�,�z$\��j�� ���9�r�=Z�h?����U�`�uޅ>�R?؈:zH<�{�>�v��!�?��v�'�Y�>�{?U��=£;>�}ž|#��{�O6����$?�?�ؾ�:;�v�u>�i%?bR?���>m�r?�gu>�J��H�<�s�>��]?�_?��F?D��>�̹=������� D���=n��>�ȅ>�}=�D>D@ҽq�	��Nż.1���ǁ�1[�V�<T��5�[���ּ�	>6mۿCK�X�پ�
�4�7?
��爾�����c��>��b�����^Yx����'�yV��6c�y����l����?�=�?�����/�� ���,�������ѵ�>��q����󫾞���)��2��b���9d!���O��&i�S�e�\�'?����ѽǿ㰡��:ܾ4  ?_A ?�y?��\�"�C�8�߲ >G`�<Z	��ڙ�O���3�ο������^?���>��7����>���>��X>�Lq>Z��Y螾�-�<��?u�-?��>��r���ɿ����ۤ<^��?��@�A?X{(�3�쾀�R=B��>lm	?@>Ո0���`��b7�>f�?h�?�}P=<�W���
�.Xe?"�<�F��лM�=���=W�=$�(�I>f�>��9�A��rٽ�]5>�0�>�C����r�\�{��<��]>=	ֽ@]���҄?yr\��f��/��P���r>N�T?�4�>�F�=��,?$CH��xϿԪ\��-a?'2�?��?k�(??ӿ��>��ܾ��M?�H6?��>wY&���t�c��=#�#���_���#V��{�=g��>�>�,������O�.���&�=	���ʿ%7"� ����<�I<��2�Ő׽�"l���蒬�i��k �R�=���=0Es>�{�>Nr>�Za>z�W?�5[?��>.�Z>��.�R���_˾9����#����H�uՒ����$��=W���Rؾ����.���	��d����<�A��=�)R�v����� �b�b��dF���.?��$>�ʾ��M��0<�<ʾ�u��\'��fB��k�˾�R1��m�f��?��A?����yW�����@�%���|�W?h.��~�������=�����=AW�>z��=��⾠�2�&tS�q�??�#?_2��萠�=�<>Q���]�=ل1?S
?s��=��>��?ő;��מ��38>�~�>���>���>�?a>�˚��l��~z#?�gW?�u��*���[>�ٸ��y��`0���R�=�>o�X'�i��=��<���L2�=^z��ף=�AT?t2�>�e-�����>�������L=�{?��?"�>(f?�C?���<*v��N�@�J��=��V?��f?$�
>%ӑ��Ծ-T��Q�6?��f?O(Z>kS��5��,�1{�DI?%�i?�@?�7��p}�7���d �w8?��v?�r^�Ns��B����V�{<�>�[�>���>�9��k�>	�>?�#��G��ֺ��Y4�Þ?o�@���?�<<��V��=�;?�\�>2�O�>ƾ�y��9�����q=f#�>#���Qev����R,�J�8?Ԡ�?���>7���N��>Y�TξO�?�?#ാwn��S���{��d@��]��39<\K��i�=�&��;B�Kz���/�F��b¼蔑>��@�E�=��Q>D���r�����d�c��� �]��zC?�@?�$=�p̽lkb��X�jhK�^�x�5ؾ0(�>�>o���D��U�x��b8�Yc����>�߼��>��O��³�o���� �<�r�>K��>j��>����IP���ޘ?�/��Ϳ�4�����#LT?7�?:��?N�?���<��f���f�VS�:�9G?!t?Ky[?M��$W��a�'�j?|_��jU`��4�jHE��U>�"3?�B�>J�-���|=�>q��>!g>�#/�o�Ŀ�ٶ�!���[��?��?�o���>j��?zs+?�i�8��|[����*�,��<A?�2>���N�!�H0=�?Ғ�ü
?L~0?{�Y.��v_?xa��=q�@.��Ž���>n�-�9Z���]� �hf�W̛�j�x��?�o�?��?O���"��e$?�}�>I���b�ž���<��>��>�{N>��]���v>^��^�:���>�K�?N[�?�?h����ߦ��H>R�}?b�>�}?~P�=̙�>��=v`־�a�ػ�=�D��n����?X?�7?���=:�.��'�9�4�\�^�}����9��\m>�A[?[�2?���>��m<�Cc�
�:���ؽA�]��緼膾^l���k��Y(>̀>�>��I�m����?*p�&�ؿ�i���o'��54?@��>�?����t�����;_?Az�>�6��+���%��UB�_��?�G�?A�??�׾BW̼>�>�I�>�Խ!���M���E�7>>�B?���D��E�o���>���?��@�ծ?pi��	?{��P���`~�����7�y��=��7?0��z>s��>��=�nv�������s�O��>�B�?�{�?���>�l?�o�m�B��1=�L�>0�k?�s?&Xo����B>��?��������K��f?��
@Ku@9�^?���п������O�@Y���=>J�>�{:>��P:>>e�>�q�9қ�<��=��$>K�>�>�Le>z�=���=��������"r��hJ*�[U �p�Ԇ�Z̫�{�1����k�����:�0���n�̜���M��X��&��}Z�=�Q?�E?�HV?92�>����#�=^Q�кm�.���4�=��>�=?�yM?My%??Z=�0����e�����k���*{�>^�?>�v�>�6�>�>��5��~>��>>�,[>f�>�u<f;=C\\=W;>���>!�>�:�>]:<>��>�δ�A.����h���v�'Z˽d��?�J��-�J��,��i��Eq��=3�=�s.?�>����� пJꭿ�H?1�����rV+�9W>��0?WbW?LL>�ݰ��T�"�>K	�A�j�!G>�, �W�l�1x)�wdQ>ё?j7g>��y>��9��;8�L�F�����Œ�>8:?�����NM�
��LG���վ��>wc�>�߹���߯���V��$j��"D={A?"�?��6�^��pm���y-l>�>~>��`=���<��;>@�����w�su'=��=2�|>��?eE>�=��>A_�[,�g�>��Y>�j4>��G?�| ?N���9��u4�����>�X�>��>߈V>a0���)>ͨ�>Lm�>`�;=Q���:����+��u�=�-�H� ������H�=�d(�b>�">�@��3n~��]��Ӗ~?U��5䈿��9c���lD?�+?#�=Z�F<��"� ���H����?m�@Qm�?g�	���V�
�?z@�?������=�}�>ث>sξ:�L���?Q ƽ'Ƣ��	�7'#��R�?a�?�/�pʋ��l��6>�^%?��Ӿ�Z�>8�aU�������u���"=���>5H?�9����P��=�څ
?�?-,����`�ȿ�hv����>��?�?��m�?��T@����>'��?�mY?��i>bf۾��Y��T�>x�@?GR?���>�o'��?�ض?ƪ�?�V>]�?4�|?_.�>���O�9��G���ې�x[x<�Æ����>�:6>����շM������U��bg~���&�	S">g��=v�>V�������jI<sEƼ�����yļh��>�[G>��a>I�>b�
?� �>��>u�v<�5�������Y����K?V��?���-n����<WÜ=�^��?%4?�fa��	о�Ĩ>_�\?�ƀ? [?�C�>��.��࿿�r��N�<.[L>�X�>�}�>[K��dK>Vվ��C���>�ӗ>'����<ھ�遾T�����>Ab!?(j�>�ڮ=�"#?�?��^>z6�>>a2�yP��bZ/��D�>���>��?!9k?�?�߼�ݗ$��)��P���QE�I�>+|?^6?���>톕�r飿��?�+��	���}w?�OT?;"���!?i��?Z�S?��R?m��>�궝����,=>�?a�f�  m��I�����Ii?a�?�b?�3�o�$�]������mfо��?yS?ih(?���,�)�l�־� �<��-;�=��q=�=k�Q>O�>7>��d�=��=s٦��լ��,����=�h>
��>vH����j�X�W�8=,?[�G�yۃ�H�=t�r�ExD���>�IL>9����^?7l=��{�����x���U�� �?���?`k�?��1�h��$=?�?Y	?�"�>�J���}޾�ྷPw��}x�ow�C�>���>��l���;���˙���F����Ž������>�<�>s�
?�.?`�>>�d�>
惾>���Ӿ<���Yr��+���H��l;��+�-���Y��B�p<ٮ���t��Jt>5밽&��>p�	?�L>�7�>e�>��2$�>d��>G��>���>˽�>s&>��=��w=OBɽ�!M?�ε�/���c����=?��`?{�>?�m�dۃ��x	�_s"?@�?���?���>Wl� �"�0�?�K�>�+z��3?A=����$=���]��.���v<��ؐ>q	�d7��J��b�s�?�?<*�^	ȾF� �N�ž��W=�+�?�E*?��,��	r�JP����x��b�z�[��G��
)������}��ۑ��`i��혿c<I��f��s%?�x�?G𪾸���DbԾŪe�
�Y�>t>� ?��F>Hf?���>,%������D�qU��2���x>K�A?�̯>�O?P�=?a�T?�,V?Ό>�Z�>헐�L��>y�=d[�>���>2>?�B4?ϡ6??�,?Ss1>�½�����žk�?�?��?�i�>'s�>-
M�4pǼ6Z�ݢ�Րp��
ؽ���<*J㻻4ֽl���Ҧ�=G�I>X�?y]ǽ�dM��9�)R>�<1?�-�>���>��h���/�.��j�>��
?\��>�8Ⱦ�=w�Äܾy �>;et?�ݫ�]�(p�=b��=~�=:��=�� >Y�(�\Yf<x㹻��~՚��H=��=
��=��<2)�<K�=��R��v�>��?���>AA�>o=���� ����Li�=�Y>�!S>>�Eپ}��?#���g�Zy>1w�?{z�?�f='�=��=򀠾}X������������<��?WI#?5XT?E��?��=?�j#?}�>&)��K��]�����<�?�7+?��>�����ʾo����0�(�?�C?�3^�����+�4eþ8�ϽW>�[*�Ym}�������B�͡�w��$���e�?�͝?uX�+�4��(�JZ�������E?ģ�>�՟>z��>��)�ci�	����?>{�>S?`��>@�L? o?�*J?�P/>�?:�ϭ���0���-�:	>�=?���?j�?��x?���>b}�=�$����!M
�*	���f��N!6=6�N>��>���>���>�|>��-�8�&�{��=<f>sk�>��>�O�>�w�>�S�<�QI?vw�>���$��o���/����2�Ļq?{��?�,?�;=���~B�U󾪚�>�Ѧ?���?�C,?��;�B6�=���vt��"�z�c�>@��>/1�>Rk�=,�F=D">�6�>���>H��d�^r5���3�ͼ?��A?�X�=��ǿ-�t��9V������=@���rSM�������z�=�����)�G��bn��'���ِ��`���줾*ˀ� ��>i=D�==��=�2P<TLp��='[=��@=�B=��e����=6�g�w:ޛ���Q2��%<8է=��:��˾L�}??0I?�+?*�C?{�y>�)>} 5�W�>,C���??�?V>��O��j���y;�\���!���"�ؾɗ׾0�c��ɟ��_>!I��>]@3>���=��<���=�Ls=h��=s�N��=/��=�a�=�D�=���=>1>?6w?뚁�J���05Q�8Z�ض:?:�>>�=��ƾ�@?^�>>=2��M����a��.?c��?�T�?2�?!vi�Bd�>���b����u�=d����>2>%��=��2�W��>p�J>���K��|���C4�?n�@��??�ዿ{�Ͽ�^/>4�">�k'>��T��L<��g�f�q��mN���?_�1���;1�r>�(6>�"��Za����=+��=���=� ���W�e��=���5(�<�!=P��>i��>y��=����E�=>��=&0=	�,>���ES��-&C;;=NV>We�>^>7G�>{�?��,?�0_?�y�>d_n���ƾ����ډ>!�=ho�>]_=�@>�>/�4?��B?&MK?�_�>���="ع>�s�>�}.��k�ڶྃ#���9�<{q�?��?�S�>z��<+�/�{3�7b9�����?�b-?��?9�>�U����,Y&���.�������/�+=Omr��OU�����m�c�㽘�=ep�>y��>�>Ty>y�9>��N>��>��>�4�<r�=���轵<�����=i�����<�zż]���!�&���+�+��� �;겆;ϰ]<���;-��=��>A<>.��>���=���FD/>������L��¿=zG��T,B�I4d�!I~�/�U6��B>K;X>8{��4����?>�Y>�m?>���?,Au?q�>� ���վ�Q��SCe�:VS��˸=��>��<��z;��Z`���M��|ҾO'�>�ђ>,Ӓ>FzH>M1���E��l2=dپ׏6�:�>��ѿ�<�C����g�Pß��0��Ph�v��Z�:?�Ʌ��e�=JRw?t<?˔?՘�>�]���پ��>�YH��a<f���o�JݽB?�]/?��?<`��@�)�ʾI���]��>��I��	O�N��?�/��C�������>ý���KѾ�3�k ���ԏ���B��bp��3�>�P?���?��^�����z=P�������[?��f?�0�>$�?l?����g�:z�K��=�.o?���?P�?��>�:>55ݽ���>�P?�?C<�?]?��R��>�>��M>�I>R3����9�a>+7M=��&>��?�
??5���Tg�8S���V��Κ��F:=��<<�[>��>� >qj�=�p�=�_�=�C?>q�=>��b>�<>Wt>�zb>�
��/2��!?+Q�=���>Xz9?��>)
P>f9>��>����]������	�4��mx���H�>L/=�[1=H�*�]��>O���)�l?_�h>e8
�Yf�>�����͍�=/B��jzQ���>�0>t�u>;�>f��>�/>
��>��s>�kҾpj>�D�8�!��~C�x6R��oѾ��|>���\6(�(��}��j'E�g������i������<� U�<JΏ?�\���l�Du)��5���?>N�>�C7?��a���>ӟ�>s�>�q���Δ�,���Qj߾�8�?���?ILc>��>��W?��?��1��)3��qZ�ܪu��&A�� e���`�����������
��~�_?��x?�}A?
j�<�7z>��?�%��ˏ�]*�>�/��!;��1<=!�>	��>�`��Ӿ�þ�E�3KF>z�o?�#�?AW?�GV���t=��w>��<?�s5?�~?eY&?�c;?,_R�Լ?��>�?�D?�66?5�3?��?�8>e�>��ż�Ӂ=s���7��ꬂ��D��Lؼ0+���;=��f=t��=Z>=��������	ͽ>s9����{�+<��*H*>��=L��>��U?��>���>wm6?]j��j[�
���5W ?�A>j�$������!���fվ��M>Y�k?�R�?��r?*� ?���h��bs=:]�>L�d>݄�>V�>AR�b�%��*>�->��=)�t<��½�s���;X�>�fv8�`��=���>(�>�� ��=/�l�a��1��>񋾽�v��Op��g�Y<��.f��?�i?�Y?oV|=L�վh��;\���?Q-S?��^?au�?���=�ھ�B�$A(�5��=��>J����a�U{���&���OE�j�=)aV>�X�g��;_>� �Gݾ+l�ˤH�˰���]=����T=���׾ʹ���=#>�Y���� ����������J?�9k=�����N�X���b�>��>�#�>Jx8�=L��ܒ?��̬���=���>��7>,`Ѽ�(�]�G�*�>c�>QlF?#�H?u?޼[�����äA������z��f�����/?��>��?��I>S�,>8�������k�=�_�oa�>���>Yo	��B5���w��~ƾ����,>���>�6>��?Dm?d?;�A?R�?�y.?���>��t<�`߾�%?#ل?&Y=�\	�n	��
G�j4� ��>)�?�r�Y��>cSa?�h@?��	?HKC?�� ?�;�=����wo��m�>���>4�C�
�ƿݶ��� �?��?�pp?��r?W�꼨�C�fՉ�oF=��Q>j�'��r?�_(?�1?�0?A�?$ 6�FDD�$G>��@?�c?^z^?�Q<>̝D?��>�G>��m�ut�>TZ?4�?�V?P�_?��H?�/?8=�=ZL=�� =>{�;V$�=��ż��$�z�=�e�P��<��< �=e��=��D=E#��r��<�\ļ���-G����>�Ct>R��\0>P�ľlD���:B>
[���C��ݤ��*�;��/�=2��>V�?� �>� #�R�=��>J��>����i'?2�?2E?m0I;c�a��gھ�L��n�>��A?Sp�=2�l��a���^u���d=L�m?x0^?��V�����kb?D3^?iW񾜩;��9ƾ�lh�����N?Hd
?� L�V}�>D�~?�q?t��>r�g���m��B��c���h��^�=�ך>s;��9d�׀�>^x6?�e�>6(f>���=��ھ��w�#���?ꐍ?���?r��?�\.>��o�`7�����o��P�2?fe?�5�C�?� �=���>Kj��;�� ���J;ɾ���f����h���
�����~�]�6��:�?/]b?;�X?�ql?b��n����v��Tv�Bq�č<�����@�+�Y�|����D�M�B�0����n]<�\M��1�ߤ�?>�-?�򯻅��>)�Q�����Ƥy��Qt>n̋���̽��i=��v���^=lo�= SN�eO3�����S�!?���>g�>�Q@?�A�1�=�h�%��M,�;k��Z9>�6�>�>=��>X)�=Np�tv;�����wHp��Ƈ�w��>I�g?�l3?��b?Lyžr�k�����m� �+��%߾���>�@h>+�>����^��� ���Z��8���F�9l��������/?���>]� >���?o?��,�3��Ã�.��R>�<��#?��?}�>�?Na�.\����>!�l?�+�> r�>�؍�b�!�jY|��̽�M�>��>���>�Vq>b�+�ӑ\�����z���9���=ٜh?|I����`����>F�Q?#" ;��8<6�>�dn��!�P��կ'�(�>�?Ԑ�=��>>��þE��*|����~7?l�?h��6��jM9>��4?gf?ɀ�>:Ly?���>)����o�j��>n�H?{�J?�,F?qX�>'b>4]���>��q�N��h�<\d>�.>�ү=Tw�=N6��)��Z��^s<�Ѽb��o"��DI�!=�l�=�f�=�U>Pۿ>K�tRپ���K�
������]��|.��w���*��@���qy�2��,&��U��Fc�9M��2�l��T�?g�?���"���%q���F��;M��S�>ـq�z���Pq����g1��A��қ���!��P�9i���e�Y�'?������ǿװ���:ܾA! ?B ?�y?���"���8��� >�I�<,��\��p�����ο����w�^?&��>l��0�����>.��>l�X>WHq>/��J瞾7�<��?��-?
��>I�r��ɿJ���ʿ�<���?��@��A?$r%�7�naH=���>C�	?ߙB>��)�[/�򋭾��>F.�?�R�?'~|=��T���"�c?#g1<��D��ˑ��=�ʤ=9�=���N�L>�S�>�L#�T�M�ecýg9>�v�>x+��m�cqY�vo�<(mW>��ٽPؕ� Մ?�z\�tf���/��T���U>��T?J+�>f>�=��,?P7H�=}Ͽѯ\��*a?�0�?ۦ�?;�(?.ڿ�8ٚ>4�ܾa�M?D6?u��>�d&���t����=�;�ߣ��`��|&V����=V��>%�>��,������O��E��U��=���.���.�vG%>Fx���	ὧ���{K���e'��2��ξ)��<��=���>�G�>d��>^�>[_8?5Cn?K�?��6>��<ՐM���h�y=v��ǀ}�x\��౾AZ�����E��O�����U�[S�qB+���=���=}&P�(��e����_�=E�#.?F�#>VR˾c�Q��1�\9ϾCB��tS��⤦��d̾�/��n��8�?�ZB?T�����S�ߢ�����F��q_Y?�O��z[�	6��Ȭ�=H���2��<D�>��=��ᾣe4�q�S���0?��?��ɾ.��i�=�����#>�:)?`��>�y�<�x>G�'?�򽱺��p�>�^->x�>��>{�=�u��F�W�[�?_�[?�l��2q��(�>w�Ӿ���;�=�vw=��W�O��<:h>����-ߚ�t�лi��=��=s�U?3U�>��$�-��꥾N ~�n�e=f�?hq�>��p>�$W?�O?5�=��þxoE�!��t�=׎M?�NU?��>٬���+پp&��W?�r?t�w>��h����6�}G����>��\?.4-?�̸�;��yD���@�ʂ8?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������f��=�\�]~�?}�?K���U�E�S8��2�aو��_(>JMH�I�߾��׾p� �*�v	(�Y�����[���>R|@==�>���>O���!Ͽ��Bp�����f&����?E+�>�=�����]���i��w��K��E���P�>��>����h����{�mo;��"��}�>���i��>ǶS�r��[�����5<��>0��>���>x/�����?�^���=ο�������6�X?Rh�?^o�?�m?��8<!�v��{��W��0G?�s? Z?rF%�(]�+A7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.���_?��a���p���-�<�ƽ�ܡ>�0��\\�h�������We�x���9y���?�\�?��?î���"�6%?n�>-����2Ǿ�3�<,��>�%�>�"N>�L_��u> �p�:��{	>M��?�}�?�i?{�������:U>��}?�;�> ڄ?���=u�>2,�=<`����f�ν">^�=G�F�n�?�rM?���>h�=� 1�>j/�-EF��S��	��rB����>��_?`L?A�o>9���%H)��� ��ڽn7)�Ke���3��;�H�ֽW:>��?>��>��9�jվ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*�[ҿ�Ƣ�����|�>=t��<�.!>�-����ͦ<u(_�n�%��=��n>��B>OH�>ߝ�>b�>��e>����,)��B���{���V,��R!�\~�u'���90��Q�����y� ������P����<F��=Y]���>.&�=��S?��M?x	o?��>�倽�$>e�����<* �+�=��>
/?��K?��+?*\�=������d��g�������ʈ�ț�>u�S>3��>�`�>���>���޼B>�J>���>�>��	=j��ew!=�bV>�ƭ>�=�>���>
I<>�>�ʹ��1��D�h��w��̽4�?*���w�J�40��K/������:v�=Qa.?N{>���<п)����0H?����x)��+�3�>��0?�cW?��>m��0�T��.>����j��g>�- ���l��)��)Q>�m?�mg>��v>�"3�F8�e�O�L+��KH>Lf6?}����9�|^u��.G���ܾicL>b�>�kA�ƴ�����~�k�h�y�k=x{9?�+? ÷�F����"s��Y����U>��]>d�=�L�=s�N>�m�vyʽ�KI�`+= �=~�^>��?�#>�y=��>c���&,+��²>��[>��Z>��B?�3?w+����ְw�/��g�>���>���>,C>R49����=�c�>lIx>��߻r�����PG�`(<>DG�:�w������=�]��0��=!�P=�|
�K�.�)݉=�~?���'䈿��e���lD?S+?a �=z�F<��"�D ���H��F�?q�@m�?��	�ۢV�A�?�@�?��P��=}�>
׫>�ξ�L��?��Ž:Ǣ�Ĕ	�$)#�hS�?��?��/�Zʋ�=l�y6>�^%?��Ӿgh�>�w�xZ�������u��#=E��>�8H?�V��~�O�q>�w
?	?�^�̩����ȿ|v����>9�?���?S�m��A���@�%��>=��?�gY?Aoi>	h۾�_Z�e��>��@?�R?^�>�9���'���?�޶?ԯ�?�GR>&�?�А?a?o5߾K�Y ˿FK�������O߼�ؿ>Ή=��Ծ���;;���1��@ۆ�Z����.>�X�=Z��>v�X�X��C2��A/6������9�=�	?��>#��>GZ�>��?�$�>{)�>�(>�P=��<R�7�J?r��?���a{��=�z>�N�_?�+�>_A����ľ��>[?歉?ޭT?�t8>����a����h������Q">���>�[�>'�v����>J�ȾI���ـ>$֤>J��u����x�\(>��>�r?(�e>�D=TI?0?�C�>Æ�>(�h��옿��j�e�m>r�>�P�>��?�;!?�s���XY�[⚿���<s��>Q�n?�{?i��>�䒿`3N.=]p����.=Z��?��N?�����{?(��?o�C?��J?���>�{=�S�k4���v�>�$?79K� i>�5#.��޽��?f?�a�>01����("��Y~۾��⾥�?�hc?X%?���O�\��tѾ+��;@�T��l�;4�=��C��53>I�[>�Aܼ���=�|>���=�g�wMv�ȴ��}>N�>�=����1�>=,?��G�9ۃ���=��r��wD��>�JL>�����^?�l=���{�q���x��FU�� �?��?=k�?
��ӝh��$=?�?n	?�"�>K��~޾ �ྱPw�}x�w�(�>b��>+�l�i�6���䙪�qF��e�Žj��5��>���>�+�>��?�0�>8ɮ>"����7��y���E��8v���=���L���%�~Q��[��!�=���%�γ��B�4��>�>#@>Ʃ�>#��>0�>���>���>".�=zn�>H��>��h>�U�>���=�&�=� >�uD�L����Q?�᣾I'������⧾�|@?�_?P �>
*��=���.!	�j�'?׶�?��?Qfu>:8f���"�� ?���>��y���>NF =��8<��=�ğ�a���ѽ�ǩ��a�>&(ѽm�4�Y|L���2�f�?�o?S�޻�Dھ�޽f�z��/>�v�?>�]?l�=�=�^���l��fz������M�����,*�����r���ᢿ�\��b�]����?f�_?�!̾(o
�iξ"*>���X���2��D?Aq�>L�>T�m>7Vj�5�\�1��h8�ԛf��x�><t?��>��8?�O%?�J?��G?H�>���>�e���|�>��<w��>�>u2!?�,3?N.5?��?�F?�:>�+�����A߾�0&?��?��?A
?� ?��5e��uB=�=A����rȽQ[W=�|�<˛7��/Q��׼���>�?r���q8�q���1g>�s7?���>�]�>�ԏ��n���ý<J=�>��
?]�>�����#q���
��8�>���?Y�����<�7&>���=�\5��s;d�=����"�=�`�mB����;l��=
�=9]��%||�77;�R�;�<�u�>�?���>}D�>]<��g� �p��8s�=<Y>S>�>�Dپ�|���#��N�g��ay>~w�?z�?�f=� �=.��=�x��MQ��c�����:��<%�?�H#?�WT?Y��?H�=?5k#?��>*��L��_��L��j�?x!,?g��>���ͳʾ��s�3���?{[?�<a�����;)���¾v�Խ
�>D[/�/~����&D�������;������?㿝?�A��6��x�˿��[��d�C? !�>�X�>��>p�)�g�g��%�L1;>��>DR?�B�>K�O?�y?y�[?��R>:�;��g��)����s���z>�A?��?�(�?C~w?���>�#>^�-�W�����[.�������@V=Q�]>�N�>�q�>t�>�G�=����ɩ��-��`�=�)_>{�><��>@��>Y�}>�V9<pI?�l�>���1��m���YN�Nƃ�x�p?8	�?U?9?��=���W>�	�����>���?�c�?��*?�E����=�2��򥱾J%r��>�6�>܈�>�Nu=2�=���=O�>�2�>������}�2�5�G��'?��B?f��=�<����j�4�U��އ��ʷ=\9v�M�5��
�:^�5���=*设��C��dȾ!B���֣�`�����K����ꊾ�m ?4=V�=�>3>W��<�b8�4Ѓ=���=��*<���<\�3<��=`=��Is\<�q���I�hT���JA�"'���˾܍}?6:I?M�+?_�C?Ӿy>�A>�w3�V��>�����>?_V>W�P�����;��������ݵؾqx׾�c�$͟�oC>=8I�"�>;43>7M�=PL�<��=�$s=6ώ=��Q��=�)�=I�=�c�=���=��>�U>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=J����=2>s��=w�2�T��>��J>���K��D����4�?��@��??�ዿТϿ6a/>$�T>
B,>!�N�W�4��S�2�/�����x$?�A�vQϾ�p|>�`>.�Ҿ�������=}'7>^#u=p�/���W�T��=��½�8$=\��=[~^>׼M>���=�0����>6�q=R:�=��(>�n?���˽k28��f=��=���>�y->V?��?¨.?^F?v��>����1�F'���(�>��>�
�>��=� �>}-�>b;?o�N?��B?["�>�0�=�Ұ>7®>fH��As�}��1y�*��kjh?�5}?N��>dx�<�����x3�F�F�Ǣ8��?�2?O:?�Q>M�Cu��q�"M�\��=����=ؼjR��V��������|�[�>m%\>:�K>���>�?���>�$?�H�>�H�=aڌ=���=��B==W<������=�+�=���=��^=
�x=W�=y�E=U�$�������<碷<e��=bz�=��>��>�@�>�G�=�����.>�����4L��Q�=�몾��B� �d���~��.�EA6���@>}LX>���M����-?y�Z>b�A>OB�?v�u?э!>|��j�Ӿ�.����e�x{T���=�>��?�
�;���_��WN�44Ӿt��>�ߎ>,�>ǻl> ,�`#?���w=��b5���>)|������(��9q�@�������i�ڳҺ��D?yF��9��=�!~?�I?\�?���>���P�ؾ�:0>�H��
�=2�3*q��e���?7'?՗�>@쾖�D��G̾�����>D=I���O���J�0� ��ͷ����>������о�$3�h��~�����B�Qr���>��O?9�?�:b��W���TO����z(���p?�|g?U�>�K?�@?�%���y�Nr���q�=~�n?���?I=�?c>��>���a��>t-?���?��?x?���ȱ?�>��=L^�\�=-&>���=�:>� ?��>zz�>�sĽ,�K�	����:���n�ག���r�>���>���>VKc=m�̽��=��*>�m>���>�t>b��>�%u>�����t� ?L4>՘�>}1?I�>;��=��n��^= y��(�D��N�����w��=T�<�96����<�l`�_�>��ÿ!U�?!��>�K ��?�9پ�� �~�F>�`>ф���>�&3>JG�>c΢>5��>A/�=��u>_J&>#JӾ�g>���V!�nC��xR�إѾ�z>팜�?�%��������nI�bu��Wf�{j��+���==�q�<DF�?�����k���)�B��� �?yS�>n6?@⌾�Y����>���>w��>"0������xˍ�mq�x
�?���?�;c>��>6�W?�?��1��3��uZ��u�E(A�e�p�`��፿�����
�d���_?��x?'yA?%Q�<+:z>H��?��%�Wӏ��)�>�/�';�:B<=�+�>*��1�`���Ӿ��þ&8��HF>o�o?2%�?_Y?\TV�k���5�>�4?l,3?A�n?0�B?��F?.�
���?sP>�?�o?�T$?��+?I�?��I>B�=ң���=da½�Ɨ�L�F�9N̽�=a�	�>=-{1=��p=�=f�=+5������眼o�5�|�`��=�R=O��=->I��>&n]?��>���>^n7?�L���7��u��7/?F�B=�M��X���衾Y��{>�$k?�ӫ?��Z?"=e>Q+A��LB��V>|�>�%>P�[>A�> �d�E�aτ=�?>z�>q�=�R�-�����	��]���B�<��>��>;�|>`��x�&>�a��p�x��e>_�P�ɿ��!�S�t�G�rK1�sdu���>��K?�?!�=������b�e��(?<?�nM?�L?+��=Ч۾M�9�XJ�'�0�>�̤<1������8����:�O+:��u>k����B�����>��� �پ�1���`��������B�9�����N�ɾ�T���[�}M�=���=0�̾�W�=_���o��(.3?�@�=#�����������4�>���=�OP>�^�=��o�K.i�0��\*`>>!�>�1>�mH<����Z�Z����D�g>u�G?��N?�%m?[�h�a+n�@���@<�������?2��>>b?��U>�]�=DK���9���m�b�W��Q�>���>]��B�I��aþ{����9O�>��?+N�>�>��P?B ?�d?�D"?�n?�j�>97�����J?H?���;�y�� z�78�`w2��>;?���o�?>��/?�H>?v)?��G??( ?�i�=^����a�v�>fo�= �=���v��=�d?�?g[z?��d?���>����H���=��J>8O�>)P3?(� ?z	X?���>��? ѽk�>x�?!s?�|~?;�Y?�/>;?E$�=�F�>�@����>�?<��>�$J?��z?GEL?��?]v�D������$�M�(J�=(�����ݽ�!�ސ������V�����ϊ�� "=���<9�s<�1�=��<�)>sC�>�5h>�,��/(9>m�þW����pD>L�ۼ6�������1��r=p�r>�?Z�>�2�h1�=�N�>�v�>V���*?c?e?�<�a�I�Ҿ��O���>��??���=�Go��T��0�r��O�=E�p?@b?��=�$s��b?�]?���5t<�ϙľR�g�{T��O?��	?�I����>�?
q?2��>��d��Bn�����Aoa�N�k�0ִ=|�>!G�H^d�)�>(l7?\�>�J]>��=
�ؾ�+x��.���m?�D�?��?p�?$�'> �n�S/࿴X+������?��?���jc(?aG�=�	�O="u�����2~�V���T��߷����J�V7�����=��M>��%?��L?+�?$0�?>r�Z�b�tタaf���`�.�'�c��kO����Ya`�K-��5]��Y��m����|>D�o�sP=�"�?}�'?El��M�>�&��;/龟v��b�K>nƔ����܈�=gA,���c=!Qe=��^�f&��ಾ�$ ?28�>~�>�6?/QV��S5�4-�k4�����;|%>���>g�>���>q���D�H��,]ƾ�Hl�I)ֽ��t>�wc?�CJ?c�m? ����1�Up��P�!��_6�����(E><>���>�7W����R&�J>�)s��j�"���R�	�o�w=)2?�d�>s�>'{�?�R?�L	�����x�T�0�,�<VJ�>^�i?SF�>�G�>��ɽ�� �j��>�l?Bi�>���>�����}!���{��$ʽ��>�}�>4�>��p>�	-�/\�pf��\����9�5��=֐h?�e��׺`���>1R?�=�:��F<�ޢ>y�Y�!�X��#�'��>�u?|E�=��<>&Iž�)��{�?����!4?��?&�ľ��*�
#>͑�>-p?�*?�g?�[�>̓㾭.��\%?\vU?#53?W6/?	� ?`]u>=uF��U=�.t	��=t5�>|�>�	>���=�x�=�ч�$�Z<��X<?>��#Ľ���;�.ཫ+4��A=��1=1mۿ�BK�t�پ�<�h?
��爾[����c������a��.��[Xx����@'�ZV�S7c����Ÿl�Ň�?�=�?(���n0�����2����������>}�q�I�����9��d)����f���Yd!���O��&i�s�e�O�'?�����ǿ򰡿�:ܾ4! ?�A ?7�y?��5�"���8�#� >�C�<�,����뾬����ο<�����^?���>��/��n��>ݥ�>�X>�Hq>����螾�1�<��?6�-?��>��r�/�ɿc���m¤<���?0�@'`A?�(�7(�OAU=go�>|	?��?>^�0�v��5���'�>��?#ߊ?�|R={RW���	�E0e?��<@�F�߬�����=L�=3=����L><p�>E����B�P۽�:4>���>� &�k���^�m��<�]>�Tӽ6���H�?�;�Q�[����&�o��>vP? ��>h�����.?8�+�p�տ��F��U?p`�?.�?k�F?C�^�R�>�;��^?�.2?�4�>��[y���1>|=��=s1ܾ�P����=_j�>��	>����+hh�Go=$�x=���ƿ�^%�w���=qֈ�1i\�3�彛���Z���Ϥo��꽗�c=��=��Q>MS�>��V>��Y>�<W?��k?���>�>c�1��>;�2	�?E���)�������]�����쾆ྟ�	������qɾ� A�xi=�U�ܑ�1���9`��VG��W/?��>1Ѿ�zO�y�<��ξ����q{��i��q9;7�1��m��|�?yh=?����ӖV�����%��燴�~U?�g�������='�ü��=_R�>'��=�{޾�V2�<�S�o�1?�?�¾�ȉ�2�!>`n���a=��-?��>B7�<���>B?���.����ce>Q�M>c�>/��>�( >֐���ؽ��?�[S?��ʽk����=�>Y����vh�B{�=;�>a��@����LU>�6;<	��G:�Vs�l�v<�V?v�>�*�Sl�=Ɛ��I�I�A=R�x?Au?��>@�j?�C?�پ<p��S�<�
�%x=�X?�h?		>�c����ϾW2��\�5?��e?��O>��e�ݣ龱�-��<�|�?�n?'?����U}�����x��5?��v?�r^�us�����T�V�f=�>�[�>���>��9��k�>�>?>#��G��񺿿cY4�)Þ?��@|��?��;<* �蜎=�;?^\�>��O��>ƾ�z������x�q=�"�>����uev����R,�d�8?ڠ�?���>擂�����1=�l�����?JN�?߰�� =v����p�|S���6�j�=$��C%����W�D����*�s��Fi='��>��@1�;GX�>�,ܽP��ΰ׿ӆr�:?�䤒�"�?,�z>82+����[x��l���z\��3Y��KG���>�MC>x��������WsL��M��s�>mU���A>�M��a<4�LN��0�!��|>�F�>K�w>�k��d�� č?'+޾�u˿5��
�վ ]I?q��?��b?˙�>�_>�)t��'O���i=�Y?�'�??�T?�
ŽQ�$����%�j?�_��xU`��4�uHE��U>�"3?�B�>S�-�q�|=�>���>g>�#/�x�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*�"�+��<A?�2>���I�!�B0=�UҒ���
?U~0?{�f.�`�_?1�a�D�p���-���ƽ�ۡ>�0��e\�P������Xe����@y����?=^�?a�?���� #�^6%?�>`����8Ǿ��<���>�(�>*N>�H_�|�u>����:�i	>���?�~�?Ij?敏������U>�}?{��>{�?�k~=���>�A>Ǹ��6�yG�=���<��F��?n�S?l�>��=�S��=^-�s"D��Q��q�a];��>�^???�I�>l#��1�� �0�3�^79�$s��K�r�H�ؼ�M��>ȴ_>4
>����v����?Ap�4�ؿ j��Ap'��54?��>�?	����t�����;_?Mz�>�6��+���%���B�]��?�G�?@�?��׾�S̼>5�>�I�>��Խ����d�����7>8�B?0��D��f�o���>���?�@�ծ?ti��	?s��K���\~�{���M7�Y�=�7?��n�z>���>z��=�mv������s�픶>�;�?_r�?���>خl?�zo���B��2=�9�>V�k?́?�v��&󾙘B>��?�������4��2f?��
@�p@�^?���+̿JP��x�
���S�w>�>!�9=/ �=nO�n��!}=����$����b=��W>��>�`�=��	>�F�=�+�����~Ǫ��t���k2��������2��@��¾��;��,��]�㾛.E�=�{��'[='�c�ۭ~�M�=�`�=2�>?��6?M(4?nE�>b=�=��n>P�ErĽSeڽq��<�k�>W7?�-8?!N4?9=Z3����]�kat�K+����l���>�`�>���>���>���>D�^=�2>Q��=_}2>�:[��0���A�����_�>6@�>��?IG�>><>��>ϴ�2��L�h��w��̽� �?C�����J� 2���6��Y���Ai�=ib.?�z>G��]>п<����1H?*���+(��+�8�>��0?IcW?<�>4����T��;>�����j��^>�+ �
l���)��!Q>�k?��e>��x>��1�sV9�[O�}.���K�>�[6?���c,0��Wv��qB���վ�%S>��>uQ��a�%���s5��4h�ߍ�=7:?��?��������x�C��1N>��S>�TF=b��=�&I>����ǽ��B�:/=���=��X>��?�2n=�Ӆ<��>	3��bE���>0�=Ҝ�=�N?y�?6�!�
�/�(�!����>���>~Y{>M��=F�	��d�=��>�]>F-|��n��@�׽�r�dzU>J(�<��v�:­�1�|=e>� ��=���=�����[�,{�=�~?���䈿}뾚f���lD?A+?� �=j�F<)�"�? ��fH��"�?X�@�l�?U�	���V�K�?�@�?�
��Y��=}�>�׫>�ξ��L���?�Ž�Ƣ���	�G)#�8S�?d�?a�/�=ʋ�:l�~5>�^%?��Ӿo&�>��E�����Gv�+�=��>�EH?d���H�S��l<�{�
?z�?��������ȿ�Tv���>0��?n�?m�m�gJ��I�?�#.�>W��?��Y?��h>�۾j�Z��
�>,�@?��Q?3��>����_'���?/׶?�l�?�|>�k�?�Hp?ϒ�>�۩��:������B���0�=��[��A�>JO>���vZR�fЗ�ϊ�4�n�E�!�Co>��y=�8�>'��ѵþ��=����i����3�)��>�y>�Q@>�C�>��?��>��>���=�wܼ�̓������>?h�?`���|p���)::k>h7"����>��?�7=�����>��a?eP{?�h?��L>�
�������������<��k>���>���>A�(�U�>��U�4�#?>-��>[�=R�˾�h�����*�>�#?f.�>Ub�=�j?�!?�(@>d�>Ԇe�_U��+�Y��\�>|��>�3�>
�?�*?�(վakE�Gꔿ����xJ�RI>Vxk?�?? '�>җ���?��l	��C3K��п=�^?�F.?Ɇ½:?C �?�+?LX?��>b��q̾�cZ���=GK>?z/����4�nԾ��n�]�?��>z؜>=b]���>���$��վ�j?yZ9?&� ?�{˾� N���[����<�G�=����5*�<:�:�"�<T��=F�ս������=�>���-��Y =��^>m�
?ב>[�2�ߊ-�4@,?�|F��݃�a�= �r�ftD��>�IL>����Y�^?u=���{�U���q���T��?N��?�j�?�����h��#=?��?�?w"�>�J��s޾.��/-w�Tyx�Ot�� >���>GLl���X������ B��:ƽ�l��8�>�A�>�q?�P?��S>���>������$��G�����V^�a�?G6��Q+�)���-��H)�R���῾��s��>H���A�>ܕ	?wSf>��>�%�>L=��T�>�~O>I�|>�>x�S>O�5>��=%T<ޏ��]�J?d��/�%��Y��g黾IWA?"�c?� ?G½S�y���]'?&G�?M
�?^ɓ>#te��q%�tc?OH�>J�r�=?�-�=f_�;<�9=-Ŏ��2
�Nv|�PIp��׋>N��o�/��bO��u�a_?W��>��-�������������?#?�0��k�爜�S���!��¾�u���ھTK~��╿�຿����e����>�i�>?E��?JG��<9��񙾪ʎ�z�Q�9��>�;�>�-f>飋>�̇>� ��%=�Y�[�����w�ѽ�>�EH?���>{�>?i3?*�Q?U�d?�֢>��>�f�8��>$��=�\>ı>��-?Z_8?p{!?�?1q?���>�Q���5���9�8?$�?��?�&?�e�>9��	�D�{�X�s�[>`�\�D<>���=���F�ľ';��w�=��(=�p&?���[/��߾���=R.?���>���>����T��hҹ�M��>?���>��ľ�G�\e�����>U�o?<̻n=�5>��R>��^��=@�>�:���t=�r;�����/ �8�K<���=>_
��ü��h�A&��(�u=�v�>@�?2��>�;�>�A��#� �H���z�=wY>S>�>vGپ�{���"����g��dy>,x�?�z�?l�f=��=5��=����`�����������<��?�K#?ZT?l��?��=?jl#?��>*�VL��]��P����?= ,?`��>�����ʾ���3�ޝ?_[?=a�β�n<)�ׇ¾*�Խ�>�V/�/~����|D�p|�����az����?$��?� A���6�]x�L����Z��u�C?�$�>MZ�>_�>	�)���g�O#��*;>>��>.
R?Y,�>��N?�w?��T?�K>7��:��%���3��7Y%>=?#I�?��?��v?���>�f>�Y$��@��7��`����X�}��=�u=>V��>���> p�>H>�%���'���/��E�=nl>!�>ع�>���>���>�=��N?(f?h1�������f��>��=�x?�}�?b�?H^��[a"���#����U�>�զ?�x�?�j0?u�轙+�=s�e;wS��?���ɣ>Cv�>8i�>,n#>;�>tg>P�>��>���E���-�XnL�2&�>�r1?�>�;�-οc�~��.�գ���+�=��<�'�y�[n;XLF���r�J���Wd,���ھ����:���6o3��J������T���;�>���=��>�#�=�oH=�(=��>"Z_=q.&>��=^������4Ӽ�}@=vQ(�k�#�n��=�=���<����֥p?��@?}�-?0�I?��>0>�竽ud�>��E?G�7>��a����vX%�r/��#��q�߾��־��]�����H>]22�ʅ0>\�->Uu�=�0= ��=/�=��M=�B��s�D=�0�=���=�ʷ=d��=�>�>�6w?X��������4Q�oZ罜�:?�8�>�{�=��ƾ�@?^�>>�2������gb��-?f��?�T�?-�?ti��d�>]���㎽�p�=����$=2>@��=r�2����>�J>����J�����l4�?��@��??�ዿ��Ͽha/>�=>C	>O��35��Ko�3\E��Y>���#?�I<��̶�;�U>��>�ǿ������<�=�#>�<R=8��@[�RV�=Elr���m=�`�=���>:c>�+�=�a���\�=�zN=�Y�=�O>:5���]S�����ѣ<)ܠ=�/>��>e��>D|?iP4?�
@?�4�>��2��[���zо�T7>M�$=A��>��]=�u>M��>��+?'�6?��J?'�>�֑=�ʴ>���>4��ꁿIA��8���p�=��?C$�?L��>ip��������)�<�M�"��"�>�v%?3��>Ǝ�>�U�V���d&�e�.�>f���.�7��*=~Mr�NU�� �h�����<��=C\�>���>��>Ly>|�9>b�N>;�>Ӷ>���<���=싻�9�<������=X'����<��ļ�\��<%�r�+�臧���;y-�;�^<+��;�D�=���>�t>���>t,�=yR���`,>�雾(�O�ы�=�#��K0=�)b��.{�@/,�&,:�;�6>^Q>>���0����?_>��6>&�?v3v?'�>����Uؾ�"��F�y�i�i�wi�=*�>�<���6�b�]��Q�&:پ�0�>6�>�->��l>{�.��/]�`=Y�rxB��.�>�#��F�=Ȟ&�y�a��ޕ��Ɯ�wOh���<7(?�ƀ�8S">q|d?�9?w��? "�>��<��
��L=��/��v�*�����3�=�(?��4?���>��2�V��n��A�_=��>�a��p}i�l���aa~��m->z�,�yJT=��ؽbH�_�*�XT��g��Зb������M>�:m?�ݢ?�q:��Ά�5Z��/��*��>_�C?c)P>Ք�>`�=?�ς>�$ƾ��&����>[?\��??��?���>�I����>
?��?�Ն? �\?�M�z��>d>W�_>�'���.1=4�>��=�h�=��?j�?
d�>
��<9����J��":����=�i>=�ii>�W'>Y̵>��=t�L�Y��<6.�=6��>0,d>vL->���>�4�>,�B!����>2��=z��>y�4?�0�>E軺�^=]k=�[ۼٞ�*�v��˽de�=�d�=�ӣ=�僽D�>�zҿ�gc?%L�>VL���>������r�Mb>C>c�����>���=��>�߃>�?>�5>>�ڴ>#�>�Ҿ��>�r��!���B�@/R��Ѿ�Cz>3Z���l%�iB�������H�"Ǵ�XJ���i������<���<nC�?������k�R�)������?�W�>��5?(j������l�>���>�3�>����Ҍ��G΍��>�?/��?Q�f>��>1	V?��?�i2�80��?Y�C�t���A�%yc���_�JJ���f���	��h���l`?x�x?�:@?U|�<�bx>��?4^%��P��% �>�|/�i:��7=n��>�X�� �]�įվg¾����J>top?塄?<>?��T�kZ�;BW�=��Q?�5?�ud?*?�u?�z���,?���>���>�>�>�M?>&?�/�>��>���=v��l�ֽ=`�:���f銽
���ƛx�aѻs㕼"�2���V<���ox�=_�=q˽�������ۙ�<	<K%e=m�>�ݯ>_]?� �>'ڎ>��2?*�0;.�5i����-?��g=��� ��l������>:;p?Ғ�?9�Z?p�\>�J�5�?���2>Zݏ>v=>'�l>}��>?$��,�4-�=��*>�}9>Z��=��0������G���w3=�v>^�>1O|>�e��tS(>�A���	z��+e>W�P�3����R���G��1� �u�.��>��K?�
?���=����O��Mf�#�(?�=<?7M?i�?��=�۾��9��sJ����M�>	-�<u��򋢿(���]�:��A5:��s>�'�� Ͼ�	�>�����x���c�-D��x��_:���R��C��𪃾�� ��i��=�������x4�����UD?G\>��E�S�o�Cg���.�>��>ʐ=ǕP��x�=�><�%�Y����=��?�Ҕ>Y�l=���2$�¦����>7TF?hkX?�'�?��r�!�q��B����}������?�X�>h? H?>S��=5������Cji�9�L�=Z�>�G�>#��K�A�ਾ��ھ@� �^��>�W	?{�!>e@	?��P?�A	?u)h?��.?&�?���>hz��/:��>"?ؔ}??케�-��oz���$��x;�Hث>�(?^G���n>�I?�?��)?]�J?�?1=>V	���G�S�>�TU>�ph�䬿�ɤ==�k?qM�>�^?�o?Gӝ=ʙ�e�{�0F*���'>+r>��(?�v?��7?Jt�>�"&?�줾�>?`L?�V?�9a?ƭT?��	�
�>s��>���=������>�m?�?Ҙ!?�=.?,p?�m�>v0�=A#��YŽ�Ц�O�ǽ&��F)K�	�'<�<������\X)=�Q�=	�>a��g��8���3�~}>yʅ=��>W�>D���Z� >�.����j�3_>�(���t��O���;� (�=k[>a ?'=�>ɽK��=�:�>�U�>m����0?�?	?Ȟ=��\�I�˾� F�z)�>�3K?�">�s������t��p<=�s?��V?B�}�%U��N�b?��]?@h��=��þ{�b����g�O?=�
?4�G���>��~?f�q?T��>�e�+:n�*��Db���j�&Ѷ=\r�>LX�R�d��?�>o�7?�N�>-�b>$%�=hu۾�w��q��h?��?�?���?+*>��n�Z4�TN��Y��T?�?������?m��h���vu������E��jT��$Ӿ���$���;td�R콾��νI1%>4��=Z��>C/Y?�r?�!������ʄ�#|��5Q��?+�p��6��-q�M}u�.����05�[�+������R�=+�n��z@���?:�)?+H����>����k���ɾ�Q8>˄���j/����=��o��wQ=�Ж=9�����b��O�?(��>^x�>�XC?T�N��+8��.��5�����QE>���>�Ԙ>��>���<�*��z���aɾ�(���c��� v>�xc?��K?��n?�Q�R+1�����;�!��G0�>U��F�B>��>���>#�W�����4&��O>���r�	���b��L�	��}=��2?+	�>8Ԝ>�J�?l�?ei	��b��_cx�2}1��ك<�V�>(i?�=�>��>�Ͻ%� �<��>Z�l?���>�>�����]!�`�{�)hʽ�0�>9׭>"��>�p>*�,�$\��k��w����9�'o�=��h?���x�`�k؅>YR?eD�:8�F<x��>5w���!�����'�$�>�x?왪=E�;>ktžc(�ڥ{�,D���?3u?-S����8����>�W,?�@?���>#TV?R��>��Ǿ���K�>݃Z?��M?$ ;?��>1'�;K3�n�����P����=hb�>-�N>���=?�>�н%�
�{xM�+����U=��I�5:����<��׺�=�46=��>�lۿ6AK��پT
��A
�鈾���Ce����_��4��sUx����r'��V�
@c������l�|��?*=�?~|��M3��󰚿����)���8��>>�q�.������ ��'(�����ɼ��(a!�^�O�'i���e�J�'?�����ǿ򰡿�:ܾ5! ?�A ?)�y?��8�"���8�C� >}D�<�+����뾦�����ο?�����^?���>���/��M��>ҥ�>P�X>�Hq>����螾�0�<��?3�-?
��>��r�&�ɿZ����¤<���?.�@y�A?:�(��e��YV=n�>(�	?0�?>�1�%8��ư�R��>�"�?�?�P=_�W��	��[e?<�F��Q׻RF�=�l�=L�=���f�J>�-�>d]��lA�8�۽w4>���>��#�����^�a��<j�]>5cԽ1X��[Ԅ?�u\�3f��/��R��9^>��T?�)�>>�=��,?�2H�n}Ͽ]�\�%)a?�/�?���?t�(?߿�bҚ>��ܾ5�M?gE6?u��>�c&�w�t�]��=7Ἦ���7�㾇%V���=_��>h|>�,�	���O�3k��5��=`�8�ƿ�$��|��^=s�ݺ��[��}�������T�^#��"fo�e�轟�h=`��=�Q>$l�>%W>�3Z>gW?��k?�N�> �>@6�S���ξ�z�	H�����O���B��h��R��߾g�	���������ɾ�#H��於 �K��2��nl2��z�}�U���V?�R�>���R��ҡ4>A��G/�YG�q�~�w�۾ 2�5�5� ݋?Z�B?�v��M5�ȣ˾�ʹ�ȩp={?�ן�]%ƾ���ʪ=}]ֻ�*=�J�>'US>�$����0��hk�,$0?;K?5�����a�(>$����I=R+?� ?��\<>�>�&%?$F*��
޽�]>�3>���>[U�>��>�G���ڽCt?�"T?%���B����>~y��
�x�Y�d=��>��7�(D����[>���<��sb4��U���δ<�W?ia�>M�)���!���C��K);=��x?�?M�>{k?�C?x)�<C���a�S��;�C�w=m�W?�5i?��>���ZKо�E����5?�we?�+O>͞h���龎�.��<�+%?��n?�Y?a���R}�������!A6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?m�;<��V��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>��������=�ٕ��Z�?}�?}����Eg<G���l��n����<9Ϋ=���D"������7���ƾ��
�ݪ��!࿼Υ�>?Z@7V�W*�>�C8�S6�TϿ$���[о`Sq���?A��>~�Ƚ����=�j��Pu�V�G�#�H������E�>ۀ%>y�ν2�����t���5��+���>��&���>�-`�������7=���>Ң�>|�>E��.[ѾKc�?Lw����οK����o�s�f?j�?���?˸?�꼛S�H^�� �;��J?=�w?5QT?)�b�P�j<�j?�_��zU`�܎4��HE��U>�"3?ZC�>�-�w�|=(>��>_g>�#/�y�Ŀ�ٶ�%���E��?܉�?�o�7��>L��?�s+?ki�8��)[����*�[�,��<A?�2>���E�!�%0=��ђ�ټ
?~0?C{��.�[�_?)�a�G�p���-�o�ƽ�ۡ>��0�f\�N�����Xe����@y����?K^�?h�?µ�� #�f6%?�>b����8Ǿ�<���>�(�>*N>jH_���u>����:�i	>���?�~�?Qj?���������U>�}?�#�>��?�l�=Ha�>�c�=]�-��k#>R �=S�>���?��M?�K�>�V�=I�8�`/�5[F��GR�K$���C�5�>��a?��L?�Lb>k��42�{!��wͽ*c1��Y鼟X@���,�Ǟ߽�(5>��=>m>k�D��Ӿ;?F���Xؿ*A��ܜ+�M3?��>�$?�k�w����_?*�>r���G���Z���m�o<�?46�?��?��־��뼘�>M6�>�؂>�нf���2���!9>D�B?�`�����&?o�/؇>h��?�d@�z�?�Hi��	?���P��Ra~�!���7���=��7?�0���z>���>+�=�nv�ݻ��]�s����>�B�?�{�?!��>�l?��o�U�B���1=7M�>��k?�s?�Xo���x�B>��?������ L��f?	�
@zu@[�^?+ٸ�Q(���ݡ�C������=r\�=(F> .����=�֕=	W.=p����>^��>�=Y>M�e>.�E>'�E>�:>����TM!�����}�J�D�( �6N���]���	��Q��.��޼�~��n�$�Z�;�ǔ������D=����M�=r�U?��Q?�o?� ?S-z�2>���z =#�8x�=�X�>9b2?�L?փ*?椓=Ot��e�r��hা�݇����>��I>���>h��>`�>v��8S�J>�?>�f�>�7>E (=ϵI�="�N>~T�>~'�>��>�$<>�>!ɴ��+����h�;�v�W@̽�?���v�J�K#��V����m�����=�[.?q>n��S2п�6'H?3�H3�95,�@�>�0?�bW?�>�����U��P>u���fj��y>����s>l�r)�V�Q>q}?��e>�v>!�3�>w8�FUP�ؗ���|>@�5?|�� [9�ztu��iH��ݾ	L>&��>�Y>�?7�����J��lh��}=6u:?�A?���/!��!Eu�������Q>�\>��=ף�=M>eI_��ƽ�G�\�4=�=z]>�k	?,�">@r�=OB�>�Ғ�s<�yǨ>˟>ً >��>?U?��^�{����rq��#���u>ڣ�>H��>�g>�2<����=��>#f`>\����*]������K�u�L>[j�ӍO������q=Rn�����=��u=5d ��<>�^�c=�~?����㈿�뾟f���lD?/+?E��=F<�"�A ��jH��:�?P�@�l�?5�	�y�V���?�@�?�	����=N{�>cի>tξ��L�j�?v�Ž*Ǣ�^�	��)#�S�?N�?��/�Gʋ�9l��6>�^%?s�Ӿ��>��7��^��j󄿔-~�ͪ��?L�>��[?7[��B��8�(��j?1?�� �T�����ʿ�l�B'�>;��?��?�b�����g7�62�>�?GY?>�v>:�׾��H��՗>��D?\�P?l�>�/��I"�~y?���?4)|?aI>���?N�s?�h�>Kx�7[/�"6������J=k[;:b�>0Z>���]gF�pד��g���j�8��"�a>��$=l�>�D�2���3�=�����H����f����>�1q>��I>X�>,� ?Tg�>=��>�x=�b���߀�򸖾��K?���? ��<n�?��<�&�=�|^��?E-4?k.]�p�Ͼ�ۨ>Ҫ\?��?�[?u�>9��1���ݿ��d���җ<�K>��>~>�>pd��uK>n�Ծ�=D�_x�>ߗ>�g���Dھ�(��iP�>q[!?.��>zZ�=	� ?S�#?o�j>b%�>dE��9���E�e��>���>
E?��~? ?й��[3�p	���硿��[�Z8N>#�x?pU?Y˕>L��������E��cI�{䒽嚂?\qg?�F彬?2�?�??��A?�.f>W���ؾ媭�C�>�0?Po>:RU��N��<!�%?74(?˚�>��ѽ�k1>v ����9�0��[?I	n?+�N?�
�0�4�G����</�>��1>��
>�> u>[�>�܀���>i��>3S�>��Ѻ�8$ɽ�߷<���>?�=��Ǿ�_�(8,?h�I������=�=�r�!gD�{�>f4L>�����^?v�=���{�����o��5�T�: �?���?Wi�?����h��=?_#�?F!?:�>o>��Ww޾����:w��Ix�/f�->���>��i�m徿���t���D��pjŽ�����>��>v�?� ?�XN>Bٱ>ݐ��w4'�6��c���a^�
�� 8��T.����3D��B&$��1�f����fz�:$�>_�����>+?)�g>wx>���>��'��>k�S>w�>��>�Y>�*4> �>�!<$Pνj?R?����q�'����ذ�oB?tSd?��>f�h�w{��L��-~?��?�g�?�!v>jh��+�nu?�;�>����q
?��8=�����<0Q���z��������ů�>�׽�:��M�Uf��^
?*$?��^̾׽�k�_t���i?�5<?�Z2��\�-���Y�.#?��S�r�=�z��TU�~ً��Z���ሿR[��^����I>Sj?�]?t3��I�琢�tj��Mz���>�X?�gP>�#�>�ǯ>�e��$2(��0r�RR)���!��J�>�i?�/�>F?��=?Y}Q?��L?%ߐ>rª>����R�>�<C��>sy�>��6?�%-?&�.?�F?]&.?��f>7g������վ�?} ?�V?��?�?2���������l�ڻO�l��h��ӗ=2N�<9V޽=q��_3=��^>+�?2��j�=��	���C>u	:?���>�:�>[�����_���"
�>�6	?A�>�߾�Cc�����>�>��w?J��؇�<tC3>��=�cJ<��;�5�=�:;l��=�>;���GQ�+u=?�=X|e<Ԁd;��=��Z=�A=�s�>7�?���>�H�>O:��t� �����]�=�	Y>�S>��>ELپ}��F"����g��gy>y�?�y�?��f=�#�=���=�m���C�����������<��?�H#?�XT?���?��=?�i#?i�>�(��K���]��D��)�?s!,?��>�����ʾ��؉3�ם?l[?�<a����;)�Ր¾��ԽǱ>�[/�j/~����=D�텻���B��3��?�?A�X�6��x�ܿ���[��z�C? "�>Y�>��>S�)�x�g�n%��1;>��>eR?a"�>�O?'2{?˚[?kaT>t�8��'��8ә��5��">� @?���?��?�y?�n�>��>Z�)�	��_���W��1� ����V=C�Y>��>��>�ک>��=*�ǽ�����>��j�=��b>ϔ�>Ō�>��>��w>8�<C>D?�?�>URľ�d�CE��9\�pfm�wto?���?qH3?>��= � �D�N�˥�w=�>���?!
�?+�?�m�}4�=A�t�n���؞\��6�>^�>��>>��=>�=��=ϼ>�*�>=��A�h8��s0�Q+?�#??�:�=��ſIp���q�����Ղ<R~���f��a��6y_��=P���w��|����`�O۠��0���u��. ����~� ��>�R�=�B�=��=��<��Љ�<��<=��L<�A=��{���g<�3�G��m؆��Z_5�(�<?=HOG���˾Ώ}?�;I?��+?O�C?��y><;>��3�虖>k����@?�V>ʛP������;����_ ���ؾ�w׾��c�	ʟ��H>�`I��>�83>|G�=�L�<��=�s=���=�R�T=�#�=�O�=�g�=k��=L�>�U>c0w?����S����8Q�^罊�:?K�>���=,wƾ7!@?��>>�4��痹�oZ��/?���?+O�?��?/�i��\�>ۢ��|�����=V���92>���=�2����>�<K>cl��O���쳽f*�?'@�??�ً�a�Ͽ�N/>ot/>��8>�~\��G��u��=m߽Fn:���?JrA��sξ�?K>�[@>�ٜ���>��=�"1>�%�=���MI�1w�=q���G6=�;</Z�>I�>�<>�t���n=�ד=w�ߺ�R>�}"��̻Ko;�_\=��&>���>�[>���>�L?��1?.c?B�>��f���ʾ$�þ"��>�2�=7��>�~=��T>�>��6?�C?�QI?q��>�P�=ꋺ>�֧>��.��(o�=3�p|��h�r<S�?��?N��>p?<��B�0��Ue=�8Q׽!�?I�/?�?�פ>�U����:Y&���.�)���v!4��+=�mr��QU�U���Jm�'�㽵�=�p�>���>��>;Ty>�9>��N>�>��>�6�<{p�=�������<� �����=�����<wż@����v&�5�+������;��;��]<���;���=��>�6>���>}��=���>/>����~�L����=�E��*B��2d��I~�/�5Y6�5�B>3X>d���83����?��Y>\i?>C��?c?u?/�>�%�I�վ�P��kDe��`S�WƸ=��>>�<��u;�+Z`���M�x�Ҿ��P>�?>�J>|gp>+�B��oc������Ks�u�󾥈�>����>��:(t�_*�������p��}��"6?�6w���w>a�i?�VF?��?�&v>YI�=W*��2�#�N�L���R�5��E��-�ؽ�JH?��S?22\>Ə���o�>��N���<�>�D=�Ra\������0h��o>xW=�7k=U�����@�C*������"����l�B1��Un�>��r?���?C
��zs�?`����v苽�R�>q�?Q� ?AI�>hĖ>U��=h�ȽH��?��<�"?��?�'�?'O>�*�=d�Ὅ(�>�.?�f�?褎?y�n?68O�Z2�>	�<4��=|s��{H>�&->붸=d�=<�
?��?SC	?�i���t�9��|��o�Q�PH=�b�=��>L��>}�w>=�=��{=ܫ�=[�b>^E�>` t>KII>B;�>J�>������*?{>]��>�|2?@�>A=&=bݣ��q�<e��誁�O�D���豽�S�=�K�=�t�=�	����>���-ܚ?�
�>���>�?�h�'�t�Y�\>�lc>��� ��>��R>�g�>�ƣ>&۔>Uc�=�g>��b>|־�$	>��� �\�C�)�R�\~׾�m�>)R���/�&�x�潔�F�Y2������yk��Á��{;�\=�֏?���p�j��5+�r��F�?���> �9?�X��H�����>Zl�>�"�>����L���
�����پm��?���?Unc>/��>�X?�?�=/�K�0�JRY�su�l�@��d�'*a�I ���t���
��0��w�_?��y?ϑA?b�<��z>.A�?��#�'x����>w.��:�)�5=��>2i���]�n�Ѿv¾����\E>f�n?���?^?�mQ��o�={�>��P?�>?��a?�'?m�;?�i��?U(t>��?�=�>�-B?]<,?k�?,gs>��>���=C3/�Ć[�b5��޷)�$���t|�Y�����i�H��'E=�=S�4�k�V<� =E��:�:Ǽ8X8=>3=4x#>Y�=;��>�-Y?�~�>\>x�7?�z�j�3��4��&I,?�X?=Q����D��1D�QL>$zj?�T�?%!Z?7Hd>�@9���>���/>O��>@�5>��_>7
�>K]���1?�j��=�>�k>�ߨ=^���	�����q<�->���>�~}>�j��x�%>|���T�w��ff>��P�.[��*�R��G��2�x:x�e$�>}�K?#x?h��=�辄,����e�z�)?	�<?�MM?%�?�
�=f!۾�9��1J�?���\�>T֒<�[	�Xt���ء���9�U��:�?p>Zʞ�㠾:Rb>H���t޾R�n��
J����BCM=�~��?V=��� ־�3�-��=e&
>{����� �����ժ��0J?�j=Yv��f`U�Ym��+�>���>bۮ>
�:���v�t�@�������=m��>&�:>Ά��e �|G��9��%�>)QE?6b_?;o�?Q7��}s�*{B�����Ң���̼��?ah�>�8?�A>��=`���f+���d��F��>	��>Ք�1�G����������$���>X�?�- >%?B�R?ͥ
?�`?O�)?aN?��>�ⷽ�\���?&?���?s�=��Խ��T�u�8�+F� ��>e�)?ƥB����>�?Z�?w�&?v�Q?��?�>� ��E@����>FS�>{�W��`�� �_>i�J?a��>�9Y?�ԃ?��=>��5���ة��B�=e>�2?27#?�?N��>��?m���ibz���>�%?�cz?���?���>�d�>ܥ�>F(?3�z>
��>�,7?Y��>O�X?!��?ă�>22�>.���JH<�|.><��}=p��0=s�=쳼�]+��21�t��X�I=�}�;O�A>��<��߽�DJ��r`�6o�>��s>"+��(�0>��ľL0���A>���I?��񺊾�S:�60�=u��>]�?���>�?#���=k��>�=�>����.(?��?�?�~ ;�b���ھ��K����>;B?��=��l�x�����u��Sh=�m?��^?�W�
%���\?l�~?��辟go��}O���J�s>�:�B?anN?���=N��>�v�?��m?>P�>����#Y�,��Qֈ�EZ���%�=�R�>���mv��K�>k4?\��>l�0>��	��}�돿(?���D?N�?Y��?>�?�*�=#��j9�W�
��e��e�E?��>hL:�4Y�>r��=��˾T?��q���;�E�~�ңϾ�ѾW�~��v�_����=��*=�6?,B?2�k?�v?1��������e��^q�7�E��Rþ��o���h���n��]j��~(��@�����[S>�	~�n�@��?�_(?Ǎ.����>����'𾨿;y�=>&������=�施�xL={L=z3j�l�*�F֬�A�?�2�>��>UB<?*�Z���=���/�^}6��(��%Q8>VZ�>�#�>�K�>��\��1�����u�̾ ���j�̽�<v>xc?��K?�n?:u��;1��|����!���/�%���C>7�>��>{GW�B�B)&��N>�$�r���������	�g��=��2?��>1�>�C�?e�?�I	��V��;�x��1���<CV�>��h?g�>���>A|н�� ����>�l?���>-0�>�����N!��{��˽���>໭>���>�o>x�,��1\�2d������!9�� �=�h?S��Q�`��݅>8�Q?N�v:D1D<��>w�u�6�!���'x'��>Wu?�Ū=�>;>N�ž? ���{�S!���*?`�?g5��3V'��>��$?1��>ȁ�>��?"1�>���S�<�?�_?��H?|cB?�8�>��= ,���&Խ��!�U=���>�\X>>�P=��=V�&�vbT�^b���I=��=9o��乽	ef<����<b��<-�7>�hۿ)IK��|پ����e�I�	��y���ز�ş����
�Mx�����I]x��O�r$'���V�Zb� Ǎ���l�k3�?���?3哾4퉾�^��P`������~�>t�o�f�v�ƫ�BX�s͗����9����u!�� P�0�h�&�e�P�'?�����ǿ���:ܾ6! ?�A ?5�y?��3�"���8� � >�C�<3-����뾬����ο>�����^?���>���/��f��>ץ�>�X>�Hq>����螾2�<��?7�-?��>��r�0�ɿb���~¤<���?-�@��H?��(�|%�i�
=���> w?H�{>Y}�W�����7�>FY�?���?x;�=�\� �1���k?m��<��@���ڼu��=œ�=�e�=�����2>[��>�,:���_�7<����k><E�>L�����0�ѷ1��=�݌>#��<y��5Մ?,{\��f���/��T��
U>��T?+�>Y:�=��,?V7H�_}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�ޅ�=b6�3���y���&V�t��=[��>i�>��,������O��I��]��=]����E������
�w�!=ʉE=��E�=�ҽ����.���>���䪾��c�y��>C�=�(>���>#��}�D>L�J?�5g?��>$�>����핾-�w�}󶻽6����H(��V������ �c۱�ǿ)�Qf$��5�4��!=�A�=�6R�J���� ���b���F���.?�v$>��ʾt�M��-<pʾ����)ل�2᥽�-̾3�1��!n�Q͟?6�A?������V����>Z�g����W?�O�����ꬾ���=������=�$�>d��=���= 3�c~S�Kt0?�6?w��G�����)>/Z�kB=4�+?ɜ ?���<a�>?�%?�'��Y��]>�N3>4�>?%�>P�>�n����۽q�?םT?�-��iY��8�>����z�Ԗj=�	>��4�Ȭ߼��]>왆<�茾�mC�['�����<�)W?���>g�)����]���j���==��x?1�?�7�>Ѐk?8�B?�_�<L��'�S����x=��W?�&i?T�>�c����Ͼ&u��ù5?��e?�N>28h����0�.��X�?��n?9f?J����r}������p6?��v?p^��z�����C�V��j�>'n�>��>��9����>�>?Y�"�B8��ԧ��rZ4�z?��@;�?'�:<f���Z�=�C?�h�>��O��Gƾu����g��̾p= ��>c���Zv�I���N,���8?��?��>J������N��=\]���2�?���?�����C������j�/?���;��q=�վ��^�����V�8��Oξ�%Y��a�0����>n@`���tg�>�!��߿V�ѿz����ξ�d���?�g�>�P��֣��n��Nt���F�R�D��~u��y�>8x>����@���'d{��:�&͛��/�>���h(�>y�R���������8<�8�>2`�>~�>@����<���ә?M��=�οV����~�ƪX?O@�?}n�?�j?�=<��u��z����FG?��r?��Y?t�$�5[��B4�D�j?&l��#r`�φ4��8E���U>�23?�D�>�v-�C�~=ߐ>���>�y>�/��Ŀ�ö��{����?u�?o꾙��>�{�?Lu+?�_�y.��"Q��3�*���s�51A?�q2>9w���!��1=�����w�
?�0?�J��*�X�_?�a�@�p�}�-���ƽ�ۡ>�0��e\��N��Y���Xe����@y����?K^�?d�?Ƶ�� #�f6%?�>v����8Ǿ��<���>�(�>6*N>�G_���u>����:�.i	>���?�~�?Vj? �������U> �}?Y��>��?�?�=�A�>SF�=w2־[t$��I1>�3T=��<�?ϠS?���>�=�= �����*�Q�A���P����R�A���_>Sh?՟I?~Z>��սB)�PS#�+�G���нs�<�lJ��p�:���iS�=��2>�E5>8�/�����4?�[�9�⿴D������J?Mj�>ǳ	?K樾8�Ž��=�?d?���>W�ؾ-���k~��a<�E�?h��?�m
?�Z߾\����=��p>٘>84<�N��{��؋>�R?d|z��+���.V�hm>⢼?�@ �?�i�R	?���Q��5`~�*����6���=��7?#,�K�z>p��>�)�=zlv�
�����s�H��>�B�?Jz�?���>۬l?��o��B�D�1=YK�>ǚk?�r?�p���[�B>�?ð�����lL�If?��
@,u@��^?y�?ѿ\͖���پwp�y�=/2�=�%>�Y��zK>�r>�ս�:���>`y>�~>�g>�L�>U1>�>�_���^#�6�������N��)��B��a6����V�N��^���ľCԽY��_D���{T�
O	�?�C >h�R?\fT?�H?r��>5u�N��=��ʾ��=�� <�>��>4K?Z�I?W0?�*>dW����o���.d���▾?,?��>ɲ�>(�?�Ӽ>w�>���>��=��=x�J;|qY<<���W�����>��>H�>�9�>"^<>7�>�ɴ�?6����h��w�0&̽2��?�f����J��/��'������M��=�x.?gu>8���Bпr����%H?Z��/$��+��X>��0?�]W?G�>F'����U���>��6�j�p%> ��fl�@�)��aQ>�N?D�f>�^u>��3�DZ8�g�P�ʜ��h,|>716?���q9���u���H�'ݾ?M>���>�FD�q�c���k/���i�ýz=qv:?��?�M������ɬu�V\���R>4�\>�=���=OM>I�b�Iǽ+H�%m/=M\�=d_>e�?|>]�.=B�>*Ζ�>�8�z�>aJ>{�->�7B?[j)?2���9���Rq��:.� X�>���>Xa�>��	>�$Q�[�=2��>a^f>S��$�������7��wK>>H����b��͊���=}����>��=6���>��/K=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>��$����-��S�^�Y��=�>�\I?�Bξj����G�	�?̬?Y�о���u����qg��/�>E��?zʘ?�r�$��5SC�	�>�2�?cX?B�q>x)���lW�>o�=?�#F?���>����~5���?2d�?&yw?��#>�W�?��?./�>~6>z�?��Tÿ����7j�=ӄ�
8��R-7��%���X�z��\�,�g�ߗ�i��>��!=�f�>�!�m쾣�=��I>�yO�} C�tܣ>É>��=z�@<	 �>�z ?���>��=��L�nH�P��,�C?="�?�E�v4��3�C������.l�f?��?u��<�Ӿ�R�>��\?v(E?踍?�Ew>�2�Q7����Ὼ��{���"7>2�5?)&B?D�e��>�ʸ��NǾ��f>���>&W5=MϦ�L���w}۽��[>!E?B|$?$Z=�S?��;?	��>�s�>e�p�eޖ���!�*�>/
 ?�k�>Z�?�7?|챾h�@����ῴ��g�Q��>�"�?|�"?b��>�:��\��I���(����i����b?P��?O>!�!?��?�%B?@7?9ǭ=\�=�f���pǾ��&>V�!?z9���A�7&�1���?�w?��>s���&�Խi�Ѽʷ�(��d?�\?"K&?pa��
a���¾E��<Y�!�X�H�o+�;�"B���>h>�
���n�=J/>Ϫ�=m�D6�
 g<3�=ǃ�>-��=7�1q���<,?��G��ك�%��=��r��vD�1�>lHL>Z��֩^?%o=���{�g���x���U�{ �?_��?6k�?����h��"=?S�?�	?!�>)I���y޾Ò�6Pw��wx�qv���>���>l�l��琤�{���$F����ŽSܽ�s�>[�>�#?V�>��w>�t>�羈�*�6������fh��T%�oM�9����,��Dо�_�=g =�&����E� �U>�����n>��>b-�>w'�>�>�.�=���>}��>&�>�N>�uH=Q5��(g߻��=�b��$LR?������'�|��k����3B?�qd?�1�>�i�ˉ��:����?���?Ds�?3;v>�~h�=,+�Zn?q>�>����p
?<R:=�4�7�<�U��w���4���t��>�A׽f :�|M�nf�Sj
?�/?j���̾&=׽��~�T������?�.\?���f�s�}�T�8�G�O�d�,�������1�/GC�6^���!��X0��9T��"�����k>J�?��?(.���6˾mم��j�X]Z��<�=���>_��>���>`̏=���C��<n�}��Ƈ9�˂�>��v?��>�CI?kg=?؃M?=�I?+q�>4Ѧ>j׭���>�΁<��>�.�>y�;?�.?+0?z?S�)?�Q>1�	�A�����ؾxq?(D?�7?c(??j�N����мhj���~��(����T=��w<�(���H�<=~uV>pl?O����8��>���j>b�7?}��>�>�ۏ�m7��ˍ�<z�>V�
?`�>y�����q�i	�*��>ϙ�?!���=��*>��=sFz����U�=�ż�َ=8���~A���<��=���=�W���!ɹv{�:��;�ư<���>e�'?��>m�>�{���ܾ���=�Z�=#� ��x,=j���yz������FL�)��>;i�?փ�?�G�=��=�d]��ë�؆k��2��i��B%
>ي"?��"?�xH?�z�?`TN?�;?�n=l]ƾ,����叿/���w6	?�,?Bϑ>>��Lʾeʨ��y3��q?�K?�Ka����!)��¾ՖӽѦ>��.�R~�����Q�C��Ŷ���d2���v�?S��?��=�(�6�t4�h����|��˴C?���>a��>'�>��)��g��J�%;>ʧ�>xR?��>��O?�:{?[?aAT>L�8��%��Yƙ��1��:">A@?S��?���?�y?4��>��>��)�`7��w�����xP󽻞���yV=<Z>�Β>b+�>zҩ>�[�=,8ȽN᰽x4?�>]�=kpb>�]�>�ƥ>��>8w>�Y�<%�G?��>��������䤾����P�;�N�u?m��?��+?�d=�l���E��-���%�>+k�?���?�/*?��S�]��=*:׼�˶��q���>f̹>�)�>�|�=��E=�e>�"�>͚�>B�c�ta8�
?L��?�F?x�=mƿ�Zt��tm�2��2��<�|����O�>����X��>=������)��m���#I�cQ��y˄���������"��FK?�M	<��=A��=�=���9�=[�?={�e<p^�<e����[=��½�e����<��e�:��B�`��=q@�<�˾��}?�;I?ە+?��C?ɹy>;>v�3�0��>A����@?�V>p�P�����1�;�P���� ��Y�ؾ@x׾ �c�ʟ��H>`I��>k83>�G�=�J�<{�=Ks=�=�R�+=�$�=UO�=jg�=@��=��>�U>�6w?R�������4Q�RZ罷�:?9�>|�=I�ƾ�@?��>>w2������Bb��-?r��?�T�?2�?�si�Wd�>&���Ꮍ)r�=Y���.=2>��=��2�.��>��J>����J��`���z4�?��@}�??�ዿ��Ͽ�a/>��7>">��R��1���\���b��YZ�ۙ!?uB;��!̾�Q�>}�=�߾�ƾ��.=��6>=�b="k��Y\�Y��=`6{�N�<=��l=kى>h�C>y`�=i��Q��=�J=�M�=�O>�����7�N,�&4=�3�=�b>�-&>m��>��??j0?�Ld?Y:�>��m�@�ξ}%���?�>�N�=�C�>5 �=׆B>�y�>��7?u�D?_�K?'S�>Iډ=)&�>q̦>½,���m��O�)����2�<뗈?�Ć?��>0�S<�UA���4N>���Ž�O?�81?�w?P�>���'ۿq�%��QN���ə�= }ݽ�Hn�>�Ӽ��T��u��\��90>J��>�>~w�>B��>��<�,>p½>de�=��5>Uߢ>�X>���=4d��pؽE)��s}�
D5�X�Q>y��=a/�=QP���b=��=Ò<)��=^��=8��>�>�t�>-�=�H���/>o���ɻL�╺=�����%B��d��\~�	a.���6��B>7TY>����
��=S?�Y>��?>�4�?<u?��!>Ji���վΝ��	d�D�Q��s�=#�>9�<�&<�l�`�n�M�GҾ�M�>;��>a\�>� p>��*�g@���b=����35�r$�>�$��c* ��¶q� D���џ��i�s$�:��D?��+_�=j�}?w�H?w�?�i�>�Þ�.(ھ*�1>����9=�3���p�e��U�?@�&?%&�>W뾔�D��̾���3�>h�G���O��Ǖ���0� F����S%�>p٪�b�о�)3��i������<�B�s��:�>��O?BѮ?�a��6���QO���� Q���&?gg?8��>>G?>Z?y����p�y�����=,�n?���?n�?5W>R6�=�ֳ��Q�>�`	?��?���?�Os?��>���>(�=;��>�����=�7
>�=���=& ?�
?~�
?T蜽� 
�s�O�W�]����<�ۤ=v��>f��>�t>���=[m=1h�=�#Z>�>�ƍ>�a>��>^J�>��������#?;��=5�>5�/?v��>�DD=�孽�;�m���A���$�/���]=ҽ��=jͻ�4V=eI��~�>�vǿ9�?��T>.���	?�)�K����I>[�M>y�.�>�{>�O>쎭>:K�>���=E��>R�>>���nY
>'ݾt�	�k��Au,��ݧ��߉>����@�����P�6��q�᤾��JJ��<l�p�@�Wٟ=���?�돾����z�L�½��?V�>,TD?�cX�����vb,>��>��Y>/���)���^j��ŭݾVV�?b"�?�<>�.�>je?I�?���=t��o�e��S��U��%w�V兿�أ�>������Sq��)>?\�\?��`?��>�.;>�n?�WӾ\'P��˼���־S9��ˉ>b�B>�:��չ�L��%�c�uE>�ߑu>+h?%�?��>>�)��v<���=��?	?�wc?k�8?�3N?�I$�c�)?e�>;?�?�7?-�7?�##?�Ò>�H>b�����<yü��z�`����D�Z`�<�2%����=��>�fu=	�<�S=Y0�����@=�<?�;mL�=~�)>�Z�>A-]?Z��>�L�>�B.?ac���4�����>?�"y��ǔ�p;���ܲ�x���ח>ɝd?�?��[?Q�q>��;���u�-3�=�ߛ>�!>$Xh>�Y�>=�L���0�~��=�h&>J�P>c� >��ν�}@�-��c|���;<r�>���>�R|>ڌ���(>	b��9y�c�d>��Q������U�V�G�d�1���v�۟�>P�K?��?�R�=���F���9)f���(?U.<?D4M?�? A�= "۾��9���J��{��E�>.m�<����ɢ�����B;��"���s>7��ؠ��Rb>M���l޾��n��J����j�M=�}��tV=����վ)����=2
>������ �K��,Ϫ��-J?w�j=�v���yU��v����>�Ƙ>��>�:���v�F�@������\�=���>�:>�!�����N{G��4���>�D?��^?�H�?	Ã���r��<B�?r��Ӡ��I��Ae?r�>��??>��=�Z��|��t�d���D����>`��>Q�x3H��(������$�퟊>�Z?�R>#�?.�T?�
?g-`?Xx*?��?��>R�˽�j��">&?텃?�=4�սG�T�)�8�AF���>�)?c�B����>�?Ⱦ?��&?�pQ?ݩ?��>�� ��9@�%��>mO�>@�W��Z��K�_>��J?��>�?Y?Tԃ?��=>�}5��䢾����{��=H/>��2?5#?t�?���> �M?(^���q�>�i~?qӜ?{��?���>��>d�?��(?w��>H�>g�#?�?U�J?�??ˏ?YN9?�����=Z���W���c��=�\���B�43��4�=3b=|j=��8>�Ž����+��\�%�=]a�>L�s>�w�/>.IľI
����A>�y�������r����9�ײ�=�>H1?�u�>s*#�Iߒ=�5�>���>l��_�'?�w?��?��;��b��ھV�I�_�>��A?;'�=��l�B]��sv���k=�m?wb^?V�V�:���rW?S�Z?�Q���P���KѺ�ܘ�g�K?-J?��h�d�>��?Uf?i)�>�����kn��睿��������>Zѧ>�~%��w�ծe>��0?��>��q>R�=�پ~%��#H���?L�?!�?-?�?�~">��c�s��;�(�|S���S?5!?�K��q?-�,�wi�ੌ:	���ْ�z���
Ծ�࠾�𪾳k	���������<� >��'?�iu?�݁?V?�����v������/3���@��@4��H��;��Sf��oY�����]���>�f�6<=��=z���H�A�<S�?�'?��0��q�>�����$�7�ִ̾B>EJ�����E�=�A���d@=@jW=xCi��'.�o㭾��?�?�>�m�>:�<?L�[���=�mB1�#{7������3>e�>�ē>#��>?B�:��.�AH�%�ɾى��܅ѽB9v>�wc?��K?Ҭn?[^��(1�1�����!��0�<S��N�B>�}>Gȉ>��W��[:&��W>�v�r�����v���	��~=e�2?�.�>C��>L�?�?�r	�@]���ix��1��?�<O=�>�i?_>�>c�>"�Ͻ�� ���>�4i?r��>��>�V��`)"�v�|�+ʻ�&��>�>��>�eY>	[4�-�Z����������7��.>� f?釀��gg�_�}>×O?�ZR�G	�<�ݟ>�R4����!澁��ha>|x?���=^3>�8Ѿ����|�c��T%?�:?�E���'7�Lǉ>T#?�
?E��>0��?�N�>�%��Y �<��?�qb?��5?��1?�8�>��=���sRƽ��F�9�^<o��>�C�>1��=�v�<Y0�u�J������==�=��\<Ow���x�=	{,;.�<8�i=uc">Dmۿ�CK�r�پ�	�~�n>
��戾�����a������a�����gYx�7����&��V�N9c������l�Y��?�<�?.~���.��=��� ���������>��q�D��8󫾗���*��.��t¬�Xd!��O�(%i��e���'?ջ����ǿ����U9ܾ�! ?B ?s�y?L�m�"��8�� >�H�<O*�����*�����οꦚ���^?���>��-6�����>楂>�X>\Iq>:���瞾�>�<��?c�-? ��>��r��ɿ1���@¤<���?�@z�A?]Y)��q�<nZ=��>�|
?	�C>b�,��[�t��w �>~�?�Ί?< Y= �V�;� ���d?D<j�E�v�Żģ�=���=��=}%�K7J>(��>m���?�!�۽e4>i��>Ԃ��*��;`�R��<d�\>3Uѽ��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=s6�򉤻{���&V�}��=[��>c�>,������O��I��U��=#���ƿv�$����m�<Wk��,Y���꽿񨽭�T�w&�� o�uy�/�f=�"�=�Q>�>�V>!�Y>IW?�Uk?ֱ�>�|>] 软<����;���������F��ہ�{n��������}	����ۈ�tIɾ�=���=S5R������� �%�b���F���.?�$>�ʾ��M�e.<�mʾy���脼�/̾�1��n��̟?v�A?���,�V�� �ja�k���E�W?�E����묾���=x���c�=�*�>���=_��� 3��S�I�/?j�?����ɔ�Ő+>L� ��!=�v,?��?E-i<��>±$?.+%��ֽ�@Y> 2>r�>(	�>w�>lG���[�>+?��T?����������> ��Lx���]=ݥ
>��2���Ӽ��Z>���<�G��S�D��x��b��<M�W?%ы>q*�~~�Qǎ��7��C=��x?�?!#�>qwk?��B?m
�<����rS��G
���z=�~W?ui?�p	>=���`ѾJ���>�5?e�e?��O>��i�K�辆'.����gW?0�n?rf?t���=}��ݒ�)6��6?��v?s^�xs�����M�V�e=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?i�;<��W��=�;?k\�>��O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������Y��=(ٕ�.Z�?��?ۆ��,�f<����l��l���f�<�ɫ=��kZ"�l��?�7��ƾ��
����������>�Y@T轺#�>�A8��5⿟RϿ����[о�Zq�3�?Q��>�Ƚ������j��Mu�e�G���H������^�>(�\=�2彠yo���Y�� ��<Mf?��ƼYؗ>��"�(v���+��ή'=��>�S�>U��>�Ž�ӯ���?�[U׿m��]o����[?�6�?�w�?�z#?-�=��r�hB��^{��� ?�c?wwa?o���-�c�}�K�j?`���U`���4�HE��U>V#3?iC�>��-�ӵ|=�>���>�g>R#/�D�ĿYٶ�����?��?ۉ�?�o�K��>g��?	s+?yi�8��[��t�*��,�v<A?k2>���2�!�20=�PҒ���
?$~0?�{�A.�Č`?h�b���q��~,���F��>�\,��(U�g�ݼj���c�����[v��_�?���?�"�?���4"�)5%?��>9����ʾ�I�<m�>�Q�>;%P>��n�w>�S�d�9�u>Z�?���?D�	?�>���T���->�L~?���>��?��=�"�>�*�=F���ѓ��^�=ˀ`=%����	?�RQ?�c�>G`�="��m.�C�+�O������<�W�`>��\?�BO?{�>-Qͽ�ʚ��=���������Q�9�U����_�G�'>�m#>3>M6�����?Mp�9�ؿ j�� p'��54?0��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ha~���y7����=��7?�0�9�z>���>��=�nv�ֻ��B�s�˹�>�B�?�{�?��>%�l?��o�e�B���1=>M�>Ԝk?�s?Ro�t󾓲B>��?������	L��f?�
@{u@b�^?6�п+~��w���Mr��=; �=�9>�gU�p�=�=�D�c����=AA>͚>ν~>!�=R�=s͛=	n��� �L'��##e��j��Y��������;�ܾ6]���E�X0������@l����0K��ޡ�%E��[�VF
>�A?�}*?��9???�
��{��=K��;ɲ�.��<xi>�Ȣ>OA<?�W?��1?���᳾��M���}�4���1���E{�>�P�>��>x ?��>O�=�ك>yҀ>Rz>o��R���2i�<��o=Ϡ�>���>���>�>��<>#>����~D���h� �w���̽��?�✾ �J�<(���㌾|A��Z�=�.?�>	��=Fп� ���H?����j���+��>��0?%�W?N>7����:T�w�>׈	��Wj�V><�����k��c)�\dQ>t�?�f>�Pu>�3�j|8���P�Xv��Σ|>�:6?�϶��9���u�c�H��#ݾ�M>:��>�E��Z�U�F�4^i�L={=;b:?Zw?)�������u�����R>>\>N}=�D�=�RM>�Ud��Lƽ��G�^7/=�>�=�^>��?��.>���=�ݚ>�����cM�A��>8L>��,>��>?�$?$��������w�NH1��q>�)�>��{>
>�7G�s�=�-�>ϐ\>���5�����83���]>������_�T�x�@�z=���ť�=���=��i)6���=��~?����䈿#�]���mD?^,?i�=��F<�"�6���-F����?5�@�l�?��	� �V�8�?�@�?.��_��=~�>�ի>�ξ��L�$�?~�Ž�Ƣ�K�	�)#��R�?�?,�/�/ʋ�>l��3>f^%?ӯӾPh�>|x��Z�������u�|�#=R��>�8H?�V����O�e>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾;`Z����>һ@?�R?�>�9�~�'���?�޶?֯�?��">2P�?��p?��>rڡ�~11�$_��&����(�<s: <o�>&g�=�Ѵ�E�֯���#���m��:�'�y>f`�=���>1��c5ӾL�%=��.���'M��6��>1*k>��2>zI�>�?���>��q>ݦ�<S�Ž=̯���19?_�?�>
�ӏ��K�� ~���%� c�>��?�U��i䖾Ś�>2�[?��Z?�?i?]|�=("��Ş�#�ֿ����z�k=�.�>�]�>��,?K�=ߓ>����8�^ۺ>�r�>��(�	{�(�P�Is�Dq>��?ؖ?���?�"?��>�7�>ͽM�l���F�D���>6��>((�>i�d??I՘��l+�x������,j�G�<r u?�y"?T�>s��4��a���B_�ݕW��m?�?�]����>@!�?��9?��C?j�>Z;ü��Ⱦ6������=��!?�T��ZA�ݧ&����3Z?�?8@�>�Ð���ѽX�ȼ���U��<h?�[?I�%?�����`�����Ę�<&�% |���;T�E�bC>��>e;��� �=I�>�}�=��l�W5��GO<P^�=v�>]�=~�5������8,?��F��σ�iߘ=x�r��wD��>�;L>�	����^?z=�d�{����x��.U�� �?��?�k�?�����h�� =?j�?�
?��>QL���{޾���Jw��ox��q���>r��>��k�@征�������F����Ž��V��<�>o-�>��?t��>�=5�6>K`�Op%��F��C��]������4��4��:�ُ�������'g<&���84����s>9,�֒�>*m?+�r>�"�>�S�>	X�=ת>;�>	!�>Ux�>E+$>0�<z껽�sֽU)ν$�R?'�¾��(�tv�}ŭ��sC?��e?�=�>�\�II������?�C�?�[�?�u>�g��M*��D?H ?V����
?n�I=OzW�"w<�����]�=�MI�~0�>�ؽ��9��IL�\�f��X	?��?�����̾׽�������=�	�?�U&?�q#���P��Qi��?��N���м�-E��D�����i%l�0����ی�qr������;�=�%?N��?�$��V��2ᶾ��g��%���6>� �>1Β>��>EE�>�ھ��"���\�V����0b�>�o?�ˉ>bx=?�4?X�D?�NK?�I�>�4�>	���E��>�Y�=���>@��>�}:?<�4?K�4?�}?��?t<>���0 ���%پ��?�4?@?� ?&Q�>�/r�f</��t�a�R��C��������W��M�<B֙���f���-<��i>W?˄%��;:�����F>�&>?�?�t�>�р�-V��{=�F�>/�?�-�>	���D�f�=��4o�>>]�?���͍s=�(6>e�H=�S��@:e�m>�=c�;?|�=�6���R���ѻ芺=7Ck=�»2�|<�"�<ajл��<eO�>��(?V��>�V�>�
t��Y�����~X<���D=��<}�Wэ�����&W_�J�t>���?�ְ?Rb>���=�3̼�����@�����ľ��Z�L�?|�#?!UY?X%�?�W?� =?,��>S�?S��(����޾��>?!,?��>q��ɵʾb�U�3���?�Z?�<a�9��w:)��¾��Խ�>fZ/��.~�i��oD�� ��e���~�����?���?[ A�z�6�Ly�ƿ��H]��C?�$�>�Y�>��>��)�9�g�:%�=3;>���>�R?��>=�O?.
{?�f[?ňT>�8�t�����<;��J">%@?˫�?I�?�y?\��>�K>��)��$�����w�)��ڔ��f�Y=�cZ>��>�	�>��>�a�=�Uǽ�����?�+Ǥ=��b>r�>c��>~��>��w>�n�<��O?雳>"�־��6��p�D�D��fk?�I�?ތ0?|N=�� G8�zm�;��>彨?CӦ?z("?�<���">W���Ӥ���Z�腻>(�>��>��`=��=��O>��>���>���b��7��ܼ�?��H?W>�ǿ�ow��3e�:#s�|¼�����M�/ �9�9�'͠=����k�_]���Ed�ӿ������+������(q���>U�<�� >��>�/W�%�w���<���<��y=��;���,��<x§�� �;�,�r��c��Tu�=I��<�p˾;�}?S+I?�}+?p�C?�{y>>�N3�Bn�>�!��>C?<!V>z�O��Y��ca;��Ũ��-����ؾ�׾��c��՟��h>
�H���>[53>Hp�= _�<�T�=��s=觎=�EZ�]A=�T�=F�=׃�=r��=��>O�>�6w?Y�������4Q��Z罦�:?�8�>z{�=��ƾr@?��>>�2������xb��-?���?�T�?=�?<ti��d�>O���㎽�q�=E����=2>x��=z�2�V��>��J>���K��?����4�?��@��??�ዿ΢Ͽ=a/>$@8>s4>�/R��2���[��b���X��m!?G	;��G˾^��>���=�Zݾ�ž�.=��4>��_=Q���\���=�B~�S==x�p=l1�>�~A>�_�=b��޸=)�K=��=v�N>���:�6�D|(�At4=�4�=o�c>��&>i>�>�P?�F*?��b?z��>�gR��?������#�>f��=��>V��=�ZU>V��>��;?�(B?�F?z��>�L�=1U�>�\�>�*3���b����tV�=눊?�P�?�v�>u�F��D��C!���E�����Q?��-?W?���>�T����@&�F.��蚽���9�,=��s���R��a��o���E�}�=�-�>�#�>���>��x>�t9>L�N>��>B�
>���<)�=<м�X.�<2���Ի�=	:��u�<�}¼/ge��f� �*��9��lN�;`i�;�g<l��;%8�=h��>f�>���>Q{�=�$����.>����A�L��9�=�E��27B�4d�B~��/�Z�6�v�B>�wX>R��*&��ٳ?�yY>��?>�q�?�-u?��>&����վ�4���d��R���=n�>�=�ҩ;��`�|�M��|Ҿ.��>Tߎ>=�>��l>�,�P#?���w=��Xb5�d�>�|�����0)��9q�'@��
���ri��aҺ�D?�F�����=G"~?ְI?D�?���>�����ؾ�;0>�H��*�=1��)q��h����?�'?���>쾉�D�Q�ξS�ǽ���>��7�IQ��ȕ�W)1�2fm�a�����>Tv��1оB�4��Ն��}�A��}k��i�>�O?6�?mM����vO�d^��禽�(�>�xf?���>���>��?�$��������\۰=T�n?���?g��?��>m>�D���F�>���>�Ɣ?���?$�q?2%콏��>�li=��_>�༎w,>���>�C%=���=�H�>�<�>� ?n���羜��H��F��%�k���>9�>"s>e&2>�z�=@h=�C>�b�>Q)Z>��>�'x>�y�>�g>������t?~5>�œ>�2?rÈ>დ=�����,=@��1����&&��N|��7=΋���=�¼ ��>��ſA&�?�h>�l�Y4?i����`�m�e>�t_>8�>��>p(>`J>�S�>Bb�>\U>2��>�0>]GӾ�}>,��b^!�B*C��R��Ѿ�z>c����&�_��K����CI��p��/i�Ij�'.���7=���<|F�?į��2�k���)�I���	�?�_�>�6?�֌����Ǯ>���>�ύ>�G������Ǎ�l���?���?D����>��N?t!?����c�Ⱦ��p�$%z�&�2�!��N����x��:=��гC�����b�T?���?(ai?�<��h>v��?��� �� ��>=���;�gm���< >���?���(���뾓�n�K��=�\u?HI�?��.?�)��ʼ��>�>.?�f&?Eb|?*~4?l�+?�ӭ�B�?�Fv>��?�~?)�5?t�5?y?��>Cn�=��f�t)�<��,���Xv��b<J�<���=�x�=�W=���<�E<C�����P�ӽQ�޽�%�a�6=�A=�y<��	>D�q=
@l?A="?�z�=�?�`���E����#�>d��#��/�S��C8�{��?&
�?8X�?9�c>��ཚg��Ot�>�`2>m�1>`0S>K��>� �=�m����>'?�>����<>�v�b������"���>|�L��>t��>10|>�	���'>�z��(.z���d>U�Q�$̺���S��G���1�i�v��Z�>~�K?'�?K��=�_龄3���Hf�o/)?�]<?�NM?��?i�=��۾�9���J�E>�E�>�K�<4�� ���t#��#�:����:�s>�0���ڠ��a>{1��-ݾ�qn��I� ��;7K=ˊ��5]=q��׾+�~�h��=t�	>d:���!�?얿L�����I?�Hl=k룾�U�CY����>=,�>���>'3��to��E@��嫾T\�=!��>\c=>'����gﾭ�G�Q��r�h>��/?#9b?H�{?b����rq���8���Ͼ�U�I�E>L��>�ph>&#?^F�<O�Y>kk׾@*�p�i��4�J��>��?�)*�2�`��.;}���#)���>�*?�р=�,7?|;�?Gv?��i?r:?� ?a�>P���{��&?Ma�?�]u=E��Pa���9���F����>�+?Š<�nH�>K�?#?Jv%?(�R?}?T�>4��.>�!��>�!�>YY�ֳ����e>�vJ?���>�Z?�=�?o6>�1�NP��<���~�=�R&>��4?��#?�e?�s�>_ ?t4��>�;{�>�/w?���?0x�?�k�>�b?�=B>W?��:>X�>��?K��>B�^?�?��N?a��>ڹ�=��<��(�0�����	=g5�V�<��2��s�=�/�<s��y�q�+$� #
�?C�(� ��?�<��g3=�Y�>(�s>����0>5�ľ�L����@>�F���P��Wي��:����=�}�>��?��>�e#����=���>�O�>��s6(?��?,?!�$;�b���ھ�K�m�>�B?��=��l�{�����u�)3h=�m?�^?�W��+����Y?��f?�i�=�X���Cc��.~��_?ل*?n��P?ہ�?��q?��>'+=3�/�`B���p}�ogd��d>���>mT$�x���-�>��G?)f�>;��>�K=�*ݾ��P�ơX���?u.�?l��?�"�?2Nu>��a��k��&��랿�?E?���>a�{���?x�|=����c��������T��� �Ѿ��������T~��첾����3�=H�?��?�6u?D�I?�m;��{�iei��{���r��J��C����9��]W���s��k�Ǒ6��"�����,3>?Ɓ�/�3�/��?b�0?�^]��@�>ċ��zr�v־�G�>�Ǧ�������=M�/��v==�7�|1��06K����U�?�͸>�d�>�L+?�逿2:G����7�(�P�����w>�̎>t�>��>~��<ƌ��������ݾ.Jƾ�E���<v>�oc?��K?P�n?���%1��}��I�!�~�/�P��5�B>�M>���>͟W����3&�:Q>�~�r����u���	�}�=>�2?m1�>���>�N�??f	�)[���nx�ǃ1��t�<Z$�>"i?P)�>�>��Ͻ� �D�>fl?�3�>?~�>����"!��{�z�ʽ�$�>%׭>g�>�m>�,�B9\��W���{��l
9��~�=k_h?s��8�`�j�>��Q?F����@<���>��u�x!�.u�X'��=><�?~i�=��<>��ž�v�i	|��W��ɵ2?>P?@�þiX,����>�??50
?���>��?R"�>w�����=�w!?	]?>�G?E�R?��?C�=�1������$����<���>8Ro>���:7;�=B��!�R���[�=4)�=�qX�����Z�<|p�<�.<�,=Gh>vgۿ�@K�<�پi����<
��舾���l��C���e���&���Tx�ܬ�*0'��4V�VPc�������l�H��??7�?�^��0)������앀�X������>5wq���~��󫾑��K��|�ྜྷ���^d!�m�O��+i�Զe�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >ZC�<	-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾x1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@�B?�'��U�:=���>KT?53O>�e$����ێ����>_p�?؋?=g=u�T����$�i?�I�<_@C���j���=y�='�=�c���D>�4�>-j�9��QȽF�6>U��>K2�*~�,\Y�\q=i�X>�ҽ�
��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�4 �]�ҿ�	-����2x�<��|=9��<|;��Q;!������ܜ:��5��R>�'�=�P>��>�dw>��5>��c?�V?���>��'>����
���u赾ӝѽ\���dƍ�裾N�T�Ⱦ;!���������4�=��Z���=��"�=�5R�_����� �]�b�z�F���.?ˆ$>+�ʾ�M�ʑ.<iʾ}���Z���ե�j/̾��1��n�D̟?�A?����2W�����;�ˑ��c�W?�B�w��Iެ�<��=�'���=9)�>��=����!3��S�r�0?S�?繾�Ǒ�Q'>�S�a�={>+?�n?G�u<�*�>��%?��(�ߐܽ?�\>Ԓ4>E�>�	�>UB>�����ܽ��?�U?��$ٜ��Q�>�о�zDz�ؕ^=��>J4��Tм��Y>���<���F�fԊ��R�<�BW?��>��)�<������:8���@=c�x?��?s)�>Z�k?��B?�<7����S�%�
���y=��W?ui?L�>.���о�X���5?f�e?�qN>�h�]���.�b��?��n??��Xx}�������Kc6?��v?�q^�t����q�V�OE�>�_�>X��>��9�Tj�>�>?� #�\E��U����W4��Þ?��@��?r.<<�"��=�:?X[�>��O�3Aƾ���̂��h�q==%�>����_cv���YN,�ȇ8?r��?��>ܒ��_��vY�=�8��ZD�?&�?^[���a<K��W�k�M����<5Ϊ=���i%����7�dLǾ�
��i��&��_��>iQ@W�潆�>)p8��.⿧OϿL��σо�p�?�?XT�>n�ɽ�7��B�j��\u���G���H�����S�>.�>�͔�����2�{�zx;��8���"�>y����>�[S�����`{����4<��>l��>"��>4կ�Iν�L��?�/���?οJ���]��X�X?HY�?Sr�?�u?�6<�tv�{�
���>G?d�s?@*Z?l$�[q]�]�8�%�j?�_��xU`���4�tHE��U>�"3?�B�>T�-�d�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>���?Z�=V��>���=�	���w�~�!>�	�=_�7�ut?5�M?���><��=K6��.���E�5R�g���9C���>Gb?L-M?��`>VS���2�!��gϽ�1���༥�@���!���⽦�3>�=>�>�uB�� Ѿx�?m���ؿ�g���\'��44?X��>r�?���B�t�����2_?�k�>n6��+���&��G�љ�?sG�?��?��׾`[̼^>#��>�?�>uս����}��_�7>��B?��hC����o���>��?H�@�Ӯ?�i��	?���P��:a~����7���=��7?�0���z>���>��=ov�ֻ��Z�s�s��>�B�?�{�?G��>�l?t�o�4�B�y�1=JM�>��k?�s?mBo��󾏱B>Z�?������L��f?�
@|u@X�^?/��п����]c��֜�A�1>*�=|
U>{4=o�>��H>�>˜7=Yh->{��>�>ܽ{>��>kΆ>nD>�~��H#�����È�|�H�F�������&��z���Ǿ4E!�X~=���� ������E���A����� ���>�IJ?9Zp?s�d?��3>��O�=R>�C��� <����>&>v�>\W8?�mL?�2?��>Nc~���Y�����_����@��}H?���>�"�>7�?Tr�>�Tͼ�1:>�i�=��R>Gk2�?~h;�㶽�ڥ���=���>� �>i�?��<>�>�ɴ��<����h�fw�ǰ˽���?�l��X�J����g ��
j���ٟ=��.?��>�
���?пh����"H? ���[�n�+�
>4�0?wpW?|V>b@���T�\�>B���j��[>T� ��_l�F�)��9Q>�G?q�i>��x>S3��e9���P��F���}>^�5?�����5���t��G���۾L\Q>�Y�>u�sP�%��g��7h���q=��:?�-?����ͱ��u�1����4S>�A\>� =��=4UL>*4S�˽x�I�ؔ4=���=��\>�$?��+>`��=�3�>�c��~eP�[�>l�A>�!+>F@?��$?N�R>��7�-���u>���>!��>��>�J���=��>F�a>2
�0������|�?��dX>A�x��j_�W�t�05~=|�����=�2�=U����>��H&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�g�>�x�IZ��R��<�u���#=1��>$8H?�V���O��>�Yv
?Y?_�������ȿ|v�$��>Z�?y��?��m�vA���@����>H��?'gY?�li>[g۾�^Z����>+�@?�R?��>�9���'���?�޶?ݯ�?�F>�7�?~s? �>��s�ݝ.�5$�� ό���x=/�;r�>�.�=j����-F�u�
�����j������e>��%=�j�>s�Wq��q�=m߉�����p����>�o>�JH>@�>/l ?b��>q|�>eC=U������h��^R?G �?�u�{���=�H�;���? � ?�>�舾�?�>��C?�~?1Vt?�@�>���8塿�PĿ4�`�� ����>��?���>�)�Ռ>����2v��=`>�2�=��r�������vO��>L��>c-?� \�[ ?f�#?�lj>L�>�OF�42���F�8B�>���>Y�?�~?�?+��B!3����k��o�[�� I><�x?�i?&�>�ӏ�P���n�<���I�#ϙ�n�?F�g?Z=��g?�ω?b�??�bB?�nh>zo��gվ�Ŵ���>��!? 	�%�A��&�l��V?�O?<�>\��SսN׼@������?fC\?jX&?̝�jNa��kþR��<W'��0B�i�<��@��Q>��>�~���F�=�>zQ�=rem�a�6�G�j<�@�=�S�>���=t�6�#���=,?��G�ۃ�i�=g�r�3xD�+�>�IL>Z����^?�l=��{�����x��O	U�� �?��?Tk�?��.�h��$=?�?H	?:"�>�J���}޾��lPw�{}x�hw�4�>&��>H�l���I���ܙ���F����Ž�n�os�>므>�?��?�%g>�@=s�)�9�����V�\���I�%��A<���K��{C�.��>�?<;N>�����@�>8��Sn>}��>T؆>/��=���>N >��E>��=ѷ�>*ɼ>>�>���=�o=<y��Tj� LR?����>�'�d��거��3B?rd?�1�>�i�$���x����?���?>s�?�<v>�~h�6,+��n?�>�>��Eq
?SR:=o6��>�<
V������3�� �(��>uE׽� :��M��nf�!j
?�/?���΋̾�;׽�u̾�k���n?�r!?���yJD� �e��?J���Y�;@'�CM��{���-D�Q���'��jې������Nd>_?�9�?=Yݾa���ﺉ���#�Z)w�A�����>e��>�ٜ>�����߾$��%�_�=o�Mb½���>��?i��>�H?�t>?sQ?T�H?f��>�G�>�����)�>ٺ�;	�>���>�9?��-?�	/?,�?@*?w9[>@"�����ؾr�?|�?+F?h ?��?�c���e�����k�w��}��o���8y=U+�<Y�ڽ�_T��s=�g\>XW?���[�8������k>��7?2|�>)��>����*�����<�	�>�
?�E�>v �(r��b�bX�>:��?�����=��)>^��=�S���ӺQW�=}���i�=�Z����;��l<�{�=Z��=�r�j�n����:��;R�<8�>|�?�>c>Į�>�>$�����%+ �>�=^0��)V�:ȯ�<�������V���d��/P>k�?��?N�=�:�='�=���Oc�������v��h)=��?T�?�^?wۙ?E,%?yz=?��!>�E�����'���z�����>� ,?���>�����ʾW񨿍�3���?�Z?S<a�W��v;)���¾��Խ<�>@[/�/~�����D����4���}��%��?��?/8A���6��v�h���}Y����C?!�>�X�>��>��)�{�g�)%��-;>���>�R?)�>N�O?�>{?��[?:MT>�8��+���љ��.3��!>�@?Ѱ�?��?�y?dt�>�>#�)���\��\���!�9҂�"qW=�Z>"��>F*�>�>k��=2ȽW��;�>�y^�=�{b>���>ڙ�>��>��w>��<f�G?���>�v����ĭ��na��1;��u?A��?�+?��=`j���E��$��;�>�o�?� �?�:*?�S���=iRּ�ⶾ�q��&�>�¹>��>r�=6;G=�n>���>���>�o��c�/v8���M���?0F?��=�ƿV�q�Āq�򠗾��g<؈��1&e�w���Z��S�=�������h���ޅ[��頾rғ��������Ƌz����>�y�=���=�J�=%��<�vļ-��<�$H=�ɍ<Ȝ=�r��Dh<J+;��.������]��`<9bJ=�����˾��}?�;I?�+?��C?2�y>�;>,�3�i��>�����@?�V>�P�����g�;����W ��=�ؾx׾��c�"ʟ�|H>�aI���>�83>H�=�O�<��=^s=�=��Q��=>$�=�O�=�g�=���=��>�U>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>Z�7>ym>6�R���1���\���b��LZ�s�!???;��&̾�#�>�b�=�߾aƾ�b/=��6>�a=���e\���=\i{�(�<=�+m=�Љ>M�C>wS�=����`�=u�I=��=��O>=��e�6��-�#3=)��=Z�b>�%>w��>��?�0?�\d?Y�>�m���ξ�2���e�>f��=�/�>� �=��B>���>��7?ЫD?��K?1{�>\��=��>��>�,�-�m���r�����<���?jˆ?��>TS<TRA�|���J>���Ľ}?�P1?��?��>���3��e�6��|&�ke����(=k(�=�<�u��<I�%�����9c�9)�=)H�>t��>ީ�>�[�>	�S>�w;>�[�>Օ=�[�<��=�P8���f=ƹX<vYp=�m9�9:��쯫�7ɼU���Ʃ�A�����/3����;��ﻕ��=i��>~>2��>���=U ��t�.><���]�L���=�P���6B��8d�@R~��/�bw6��B>�eX>w.��b*���?�Y>�\?>Su�?I?u?�>,��P�վi6����d�fS����=I�>j�<���;��i`�y N���Ҿ_��>B��>�t�>`Yl>�S+��>�X$m=k�㾏N5���>>��ɿ'���1q��I�������h��\�9E?������=f�}?%4I?�Տ?j��>������ؾ�0>ھ����=���y%q�T㒽4?]9'?��>^!��D���о{�Ľ�>��;���I�4���	4��!!��躾�u�>�<��k#ھv�5�߅��%��aAG� �{���>�YT?*��?�M�"J����N�-�3����>�:Z?��>0�?o�?��ѽd~���]��0�= �h?7R�?�a�?ŝ>1��=�#�� �	??dM�?��?�R|?�f,�Z�>猤;�>j�7�}�>�l.>�8w=
u>y?eg?; ?�w������� �)� ����7�=+�>Ǻ�>��>3��>m�
>i*�=|��=9�r>��>&��>�}s>r�>v�>Sh���w���&?���=ݣ�>�2?�.�>YyX=L1��d*�<�SK�>I@�P+�!����nὖ˹<ҙ���O=��̼�>2nǿ�=�?o�S>���u�?R����0��nT>a�U>��޽���>Y^F>�E}>kѮ>��>gb>���>c�'>rIӾ�y>E��a!�>)C�>�R���Ѿ8hz>7���]&�N������PI�]r��_l�j��-��67=��w�<dF�?�����k� �)�3���)�?�T�>�6?�֌��舽�>[��>�Ǎ>U=������Ǎ��`���?d��?�6�=��>m
,?G?���=6�<��;p��ې���=�RSy��z�����4؏��N'�6�]��[+?�$f?ZXV?�M>��>�}U?9������j:>"�B�����>�`|=�Q�t���%	��/v������
�>�?�?NV�?�c?�xо�� ���#>��??�|.?��s?�1?��B?s�����)?�F>,?C?+C3?�0?wu?��E>�>4�:<r5J=����y�����;k���*�=�Cq=VѲ</��<�H�=Yא=[�-�Լ�a�<L�T<�NE=�=1�=��=8)�>��\?���> :�>��7?S���9�w䰾��+?�e=Ep������+S��������=��j?���?�$[?�f>Y?>���C��>�r�>�5 >�2Z>�Ұ>��սx2O�v�=)>�>!��=��X�!����3	����^�<E;>f��>/1|>s
���'>}���1z���d>��Q�K̺���S�)�G�F�1�*�v�=Z�>"�K?��?ڜ�=�_�M1��'If��/)?�]<?OM?p�?��=R�۾��9���J��>���>0R�<l�������#����:� ��:�s>1���ڠ��a>{1��-ݾ�qn��I� ��;7K=ˊ��5]=q��׾+�~�h��=t�	>d:���!�?얿L�����I?�Hl=k룾�U�CY����>=,�>���>'3��to��E@��嫾T\�=!��>\c=>'����gﾭ�G�Q��r�h>��/?#9b?H�{?b����rq���8���Ͼ�U�I�E>L��>�ph>&#?^F�<O�Y>kk׾@*�p�i��4�J��>��?�)*�2�`��.;}���#)���>�*?�р=�,7?|;�?Gv?��i?r:?� ?a�>P���{��&?Ma�?�]u=E��Pa���9���F����>�+?Š<�nH�>K�?#?Jv%?(�R?}?T�>4��.>�!��>�!�>YY�ֳ����e>�vJ?���>�Z?�=�?o6>�1�NP��<���~�=�R&>��4?��#?�e?�s�>_ ?t4��>�;{�>�/w?���?0x�?�k�>�b?�=B>W?��:>X�>��?K��>B�^?�?��N?a��>ڹ�=��<��(�0�����	=g5�V�<��2��s�=�/�<s��y�q�+$� #
�?C�(� ��?�<��g3=�Y�>(�s>����0>5�ľ�L����@>�F���P��Wي��:����=�}�>��?��>�e#����=���>�O�>��s6(?��?,?!�$;�b���ھ�K�m�>�B?��=��l�{�����u�)3h=�m?�^?�W��+����Y?��f?�i�=�X���Cc��.~��_?ل*?n��P?ہ�?��q?��>'+=3�/�`B���p}�ogd��d>���>mT$�x���-�>��G?)f�>;��>�K=�*ݾ��P�ơX���?u.�?l��?�"�?2Nu>��a��k��&��랿�?E?���>a�{���?x�|=����c��������T��� �Ѿ��������T~��첾����3�=H�?��?�6u?D�I?�m;��{�iei��{���r��J��C����9��]W���s��k�Ǒ6��"�����,3>?Ɓ�/�3�/��?b�0?�^]��@�>ċ��zr�v־�G�>�Ǧ�������=M�/��v==�7�|1��06K����U�?�͸>�d�>�L+?�逿2:G����7�(�P�����w>�̎>t�>��>~��<ƌ��������ݾ.Jƾ�E���<v>�oc?��K?P�n?���%1��}��I�!�~�/�P��5�B>�M>���>͟W����3&�:Q>�~�r����u���	�}�=>�2?m1�>���>�N�??f	�)[���nx�ǃ1��t�<Z$�>"i?P)�>�>��Ͻ� �D�>fl?�3�>?~�>����"!��{�z�ʽ�$�>%׭>g�>�m>�,�B9\��W���{��l
9��~�=k_h?s��8�`�j�>��Q?F����@<���>��u�x!�.u�X'��=><�?~i�=��<>��ž�v�i	|��W��ɵ2?>P?@�þiX,����>�??50
?���>��?R"�>w�����=�w!?	]?>�G?E�R?��?C�=�1������$����<���>8Ro>���:7;�=B��!�R���[�=4)�=�qX�����Z�<|p�<�.<�,=Gh>vgۿ�@K�<�پi����<
��舾���l��C���e���&���Tx�ܬ�*0'��4V�VPc�������l�H��??7�?�^��0)������앀�X������>5wq���~��󫾑��K��|�ྜྷ���^d!�m�O��+i�Զe�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >ZC�<	-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾x1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@�B?�'��U�:=���>KT?53O>�e$����ێ����>_p�?؋?=g=u�T����$�i?�I�<_@C���j���=y�='�=�c���D>�4�>-j�9��QȽF�6>U��>K2�*~�,\Y�\q=i�X>�ҽ�
��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�4 �]�ҿ�	-����2x�<��|=9��<|;��Q;!������ܜ:��5��R>�'�=�P>��>�dw>��5>��c?�V?���>��'>����
���u赾ӝѽ\���dƍ�裾N�T�Ⱦ;!���������4�=��Z���=��"�=�5R�_����� �]�b�z�F���.?ˆ$>+�ʾ�M�ʑ.<iʾ}���Z���ե�j/̾��1��n�D̟?�A?����2W�����;�ˑ��c�W?�B�w��Iެ�<��=�'���=9)�>��=����!3��S�r�0?S�?繾�Ǒ�Q'>�S�a�={>+?�n?G�u<�*�>��%?��(�ߐܽ?�\>Ԓ4>E�>�	�>UB>�����ܽ��?�U?��$ٜ��Q�>�о�zDz�ؕ^=��>J4��Tм��Y>���<���F�fԊ��R�<�BW?��>��)�<������:8���@=c�x?��?s)�>Z�k?��B?�<7����S�%�
���y=��W?ui?L�>.���о�X���5?f�e?�qN>�h�]���.�b��?��n??��Xx}�������Kc6?��v?�q^�t����q�V�OE�>�_�>X��>��9�Tj�>�>?� #�\E��U����W4��Þ?��@��?r.<<�"��=�:?X[�>��O�3Aƾ���̂��h�q==%�>����_cv���YN,�ȇ8?r��?��>ܒ��_��vY�=�8��ZD�?&�?^[���a<K��W�k�M����<5Ϊ=���i%����7�dLǾ�
��i��&��_��>iQ@W�潆�>)p8��.⿧OϿL��σо�p�?�?XT�>n�ɽ�7��B�j��\u���G���H�����S�>.�>�͔�����2�{�zx;��8���"�>y����>�[S�����`{����4<��>l��>"��>4կ�Iν�L��?�/���?οJ���]��X�X?HY�?Sr�?�u?�6<�tv�{�
���>G?d�s?@*Z?l$�[q]�]�8�%�j?�_��xU`���4�tHE��U>�"3?�B�>T�-�d�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>���?Z�=V��>���=�	���w�~�!>�	�=_�7�ut?5�M?���><��=K6��.���E�5R�g���9C���>Gb?L-M?��`>VS���2�!��gϽ�1���༥�@���!���⽦�3>�=>�>�uB�� Ѿx�?m���ؿ�g���\'��44?X��>r�?���B�t�����2_?�k�>n6��+���&��G�љ�?sG�?��?��׾`[̼^>#��>�?�>uս����}��_�7>��B?��hC����o���>��?H�@�Ӯ?�i��	?���P��:a~����7���=��7?�0���z>���>��=ov�ֻ��Z�s�s��>�B�?�{�?G��>�l?t�o�4�B�y�1=JM�>��k?�s?mBo��󾏱B>Z�?������L��f?�
@|u@X�^?/��п����]c��֜�A�1>*�=|
U>{4=o�>��H>�>˜7=Yh->{��>�>ܽ{>��>kΆ>nD>�~��H#�����È�|�H�F�������&��z���Ǿ4E!�X~=���� ������E���A����� ���>�IJ?9Zp?s�d?��3>��O�=R>�C��� <����>&>v�>\W8?�mL?�2?��>Nc~���Y�����_����@��}H?���>�"�>7�?Tr�>�Tͼ�1:>�i�=��R>Gk2�?~h;�㶽�ڥ���=���>� �>i�?��<>�>�ɴ��<����h�fw�ǰ˽���?�l��X�J����g ��
j���ٟ=��.?��>�
���?пh����"H? ���[�n�+�
>4�0?wpW?|V>b@���T�\�>B���j��[>T� ��_l�F�)��9Q>�G?q�i>��x>S3��e9���P��F���}>^�5?�����5���t��G���۾L\Q>�Y�>u�sP�%��g��7h���q=��:?�-?����ͱ��u�1����4S>�A\>� =��=4UL>*4S�˽x�I�ؔ4=���=��\>�$?��+>`��=�3�>�c��~eP�[�>l�A>�!+>F@?��$?N�R>��7�-���u>���>!��>��>�J���=��>F�a>2
�0������|�?��dX>A�x��j_�W�t�05~=|�����=�2�=U����>��H&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�g�>�x�IZ��R��<�u���#=1��>$8H?�V���O��>�Yv
?Y?_�������ȿ|v�$��>Z�?y��?��m�vA���@����>H��?'gY?�li>[g۾�^Z����>+�@?�R?��>�9���'���?�޶?ݯ�?�F>�7�?~s? �>��s�ݝ.�5$�� ό���x=/�;r�>�.�=j����-F�u�
�����j������e>��%=�j�>s�Wq��q�=m߉�����p����>�o>�JH>@�>/l ?b��>q|�>eC=U������h��^R?G �?�u�{���=�H�;���? � ?�>�舾�?�>��C?�~?1Vt?�@�>���8塿�PĿ4�`�� ����>��?���>�)�Ռ>����2v��=`>�2�=��r�������vO��>L��>c-?� \�[ ?f�#?�lj>L�>�OF�42���F�8B�>���>Y�?�~?�?+��B!3����k��o�[�� I><�x?�i?&�>�ӏ�P���n�<���I�#ϙ�n�?F�g?Z=��g?�ω?b�??�bB?�nh>zo��gվ�Ŵ���>��!? 	�%�A��&�l��V?�O?<�>\��SսN׼@������?fC\?jX&?̝�jNa��kþR��<W'��0B�i�<��@��Q>��>�~���F�=�>zQ�=rem�a�6�G�j<�@�=�S�>���=t�6�#���=,?��G�ۃ�i�=g�r�3xD�+�>�IL>Z����^?�l=��{�����x��O	U�� �?��?Tk�?��.�h��$=?�?H	?:"�>�J���}޾��lPw�{}x�hw�4�>&��>H�l���I���ܙ���F����Ž�n�os�>므>�?��?�%g>�@=s�)�9�����V�\���I�%��A<���K��{C�.��>�?<;N>�����@�>8��Sn>}��>T؆>/��=���>N >��E>��=ѷ�>*ɼ>>�>���=�o=<y��Tj� LR?����>�'�d��거��3B?rd?�1�>�i�$���x����?���?>s�?�<v>�~h�6,+��n?�>�>��Eq
?SR:=o6��>�<
V������3�� �(��>uE׽� :��M��nf�!j
?�/?���΋̾�;׽�u̾�k���n?�r!?���yJD� �e��?J���Y�;@'�CM��{���-D�Q���'��jې������Nd>_?�9�?=Yݾa���ﺉ���#�Z)w�A�����>e��>�ٜ>�����߾$��%�_�=o�Mb½���>��?i��>�H?�t>?sQ?T�H?f��>�G�>�����)�>ٺ�;	�>���>�9?��-?�	/?,�?@*?w9[>@"�����ؾr�?|�?+F?h ?��?�c���e�����k�w��}��o���8y=U+�<Y�ڽ�_T��s=�g\>XW?���[�8������k>��7?2|�>)��>����*�����<�	�>�
?�E�>v �(r��b�bX�>:��?�����=��)>^��=�S���ӺQW�=}���i�=�Z����;��l<�{�=Z��=�r�j�n����:��;R�<8�>|�?�>c>Į�>�>$�����%+ �>�=^0��)V�:ȯ�<�������V���d��/P>k�?��?N�=�:�='�=���Oc�������v��h)=��?T�?�^?wۙ?E,%?yz=?��!>�E�����'���z�����>� ,?���>�����ʾW񨿍�3���?�Z?S<a�W��v;)���¾��Խ<�>@[/�/~�����D����4���}��%��?��?/8A���6��v�h���}Y����C?!�>�X�>��>��)�{�g�)%��-;>���>�R?)�>N�O?�>{?��[?:MT>�8��+���љ��.3��!>�@?Ѱ�?��?�y?dt�>�>#�)���\��\���!�9҂�"qW=�Z>"��>F*�>�>k��=2ȽW��;�>�y^�=�{b>���>ڙ�>��>��w>��<f�G?���>�v����ĭ��na��1;��u?A��?�+?��=`j���E��$��;�>�o�?� �?�:*?�S���=iRּ�ⶾ�q��&�>�¹>��>r�=6;G=�n>���>���>�o��c�/v8���M���?0F?��=�ƿV�q�Āq�򠗾��g<؈��1&e�w���Z��S�=�������h���ޅ[��頾rғ��������Ƌz����>�y�=���=�J�=%��<�vļ-��<�$H=�ɍ<Ȝ=�r��Dh<J+;��.������]��`<9bJ=�����˾��}?�;I?�+?��C?2�y>�;>,�3�i��>�����@?�V>�P�����g�;����W ��=�ؾx׾��c�"ʟ�|H>�aI���>�83>H�=�O�<��=^s=�=��Q��=>$�=�O�=�g�=���=��>�U>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>Z�7>ym>6�R���1���\���b��LZ�s�!???;��&̾�#�>�b�=�߾aƾ�b/=��6>�a=���e\���=\i{�(�<=�+m=�Љ>M�C>wS�=����`�=u�I=��=��O>=��e�6��-�#3=)��=Z�b>�%>w��>��?�0?�\d?Y�>�m���ξ�2���e�>f��=�/�>� �=��B>���>��7?ЫD?��K?1{�>\��=��>��>�,�-�m���r�����<���?jˆ?��>TS<TRA�|���J>���Ľ}?�P1?��?��>���3��e�6��|&�ke����(=k(�=�<�u��<I�%�����9c�9)�=)H�>t��>ީ�>�[�>	�S>�w;>�[�>Օ=�[�<��=�P8���f=ƹX<vYp=�m9�9:��쯫�7ɼU���Ʃ�A�����/3����;��ﻕ��=i��>~>2��>���=U ��t�.><���]�L���=�P���6B��8d�@R~��/�bw6��B>�eX>w.��b*���?�Y>�\?>Su�?I?u?�>,��P�վi6����d�fS����=I�>j�<���;��i`�y N���Ҿ_��>B��>�t�>`Yl>�S+��>�X$m=k�㾏N5���>>��ɿ'���1q��I�������h��\�9E?������=f�}?%4I?�Տ?j��>������ؾ�0>ھ����=���y%q�T㒽4?]9'?��>^!��D���о{�Ľ�>��;���I�4���	4��!!��躾�u�>�<��k#ھv�5�߅��%��aAG� �{���>�YT?*��?�M�"J����N�-�3����>�:Z?��>0�?o�?��ѽd~���]��0�= �h?7R�?�a�?ŝ>1��=�#�� �	??dM�?��?�R|?�f,�Z�>猤;�>j�7�}�>�l.>�8w=
u>y?eg?; ?�w������� �)� ����7�=+�>Ǻ�>��>3��>m�
>i*�=|��=9�r>��>&��>�}s>r�>v�>Sh���w���&?���=ݣ�>�2?�.�>YyX=L1��d*�<�SK�>I@�P+�!����nὖ˹<ҙ���O=��̼�>2nǿ�=�?o�S>���u�?R����0��nT>a�U>��޽���>Y^F>�E}>kѮ>��>gb>���>c�'>rIӾ�y>E��a!�>)C�>�R���Ѿ8hz>7���]&�N������PI�]r��_l�j��-��67=��w�<dF�?�����k� �)�3���)�?�T�>�6?�֌��舽�>[��>�Ǎ>U=������Ǎ��`���?d��?�6�=��>m
,?G?���=6�<��;p��ې���=�RSy��z�����4؏��N'�6�]��[+?�$f?ZXV?�M>��>�}U?9������j:>"�B�����>�`|=�Q�t���%	��/v������
�>�?�?NV�?�c?�xо�� ���#>��??�|.?��s?�1?��B?s�����)?�F>,?C?+C3?�0?wu?��E>�>4�:<r5J=����y�����;k���*�=�Cq=VѲ</��<�H�=Yא=[�-�Լ�a�<L�T<�NE=�=1�=��=8)�>��\?���> :�>��7?S���9�w䰾��+?�e=Ep������+S��������=��j?���?�$[?�f>Y?>���C��>�r�>�5 >�2Z>�Ұ>��սx2O�v�=)>�>!��=��X�!����3	����^�<E;>f��>/1|>s
���'>}���1z���d>��Q�K̺���S�)�G�F�1�*�v�=Z�>"�K?��?ڜ�=�_�M1��'If��/)?�]<?OM?p�?��=R�۾��9���J��>���>0R�<l�������#����:� ��:�s>1��Aܠ��\b>:���q޾Śn�,J�����QM=~��1V=����վ4�'��=�
>Ѽ��g� �%���֪�b/J?��j=u��!dU��i���>���>ݮ>��:���v�؇@������B�=1��>!�:>�k��<���}G��:�(>�>��M?�F`?���?oQ,� 9����F�����n��[�>��'?}p�>�l�>�v� Ϥ<�þ^,:��_d�e�&�(h�>�<�>�L-���4��VϾ��!���8��%�>��?� >��?&fZ?m�?�i??��.?���>^Ѐ>��;WS&?�N�?�x�=xCս�U�D8���D�#��>�5*?з>�}?�>{l?6�?�&?��Q??U>���i@�<z�>W��>�	X�}���`>�J?���>p�X?�˃?/O=>]5�����;
�����=">z"3?ˉ"?��?��>�?�Ľ�뷼��>�?��?��?�}�>�O�>���>W�%?I�.>��>�?^�?rgr?Dx?e� ?���>�!�=g��;ƽ%�<	q��#��<)��=�U�=1����㼴���I�!�Dg�:�*�Ts콂]H���<�D2�����_�>k�s>���e�0>�ľjO����@>Q���N���܊�[�:��ַ=ƃ�>6�?f��>5]#����=Z��>tJ�>���*6(?�?y?�";u�b���ھ<�K��>�	B?���=��l�G�����u��h=?�m?��^?��W��#����e?o�s?�m�rj!��P���_�T��cK?�?��g���>�݀?z�W?��>g�ĽĢ[�ў�����aվ34>bu�>/E1�C������=N+V?�?Be=>�lQ^�v��ִ�DK?�?��?T=~?�X�>�N����0���'���6C?*)?�Պ�ͣ�>>� =a�оv�=���둻�G�ٽ;�󾟗�ݽ�QBf�;̚�T���T�=gN?�1v?��?��?I,0�W�F���n��D����I�τ��.�-%U�\w�9�w�QՒ�m���6�k���Nc+>[�~���A�΀�?�'?į/����>͎��Q��Љ̾nB>�c���7�{�=0ƌ��?=��Z=іh�*N.��5�� ?�ݹ>I��> �<?9�[��,>�ǌ1�,�7�~���(c3>�ߢ>��>���>�5^:�p-�[�齇�ɾ����Otҽ�Fv>�rc?�K?3�n?���-1��y���!�X�/�	����`B>�G>��>��W�Q�AC&��s>�h�r����ch��7�	�e�~=`�2?,�>`j�>�=�?&?�	������w�gT1�Mʅ<$��>�i?�4�>^��>5ѽ�� ����>�l?�	?%��>1���I$��+p��Ꜿ���>��>�<D>q�;G�¾K�R�0��W3��K�K�ڇ>0Wh?z�v��#��\p>8|)?�7ɽ�y��q�>�`�>��Z5��M>4e�>�.?��	=-�>a�:�p+U��Q����f�??��	?_-|�̱���@>��[?�*?�&�>��?�?��T��<�=�*? po?�"D?v�m?���>s;Ƚ��|�d������%���*>6؂>�w	>9�=R�(]�>=�Qb&���=�1=S��<*/�/\�<���=qb�=��p> ^ۿk?K��پT��I�;*
��������Q@��y���N��px��f�p�&�s�U�{�b�2{���l�nw�?�7�?h6���ȉ�����o�������W�>�Qq��Y������E�<���z��&(��t�!��P��#i� �e�O�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��8�"���8�� >ZC�<-����뾭����οA�����^?���>��/��o��>ۥ�>�X>�Hq>����螾x1�<��?8�-?��>Îr�0�ɿb����¤<���?0�@}A?@�(�"��@�U=���>��	?��?>zN1�I�i���$X�>i<�?���?'�M=	�W���	��~e?RQ<�F�h�ݻ��=H�=hm=��h�J>�S�>ф��OA�-/ܽ��4>�ۅ>�h"�I����^�<��<v�]>�սs*��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=���ǩ��:�%�d�$��uӽ�u�<���<\O������㚽-���	?�����(��=j}	>Eq>b�>:�n>N>��P?�(k?x�>E�E>�3D�	ٕ���>]q�a�<�0d9�A����)�1������8������"&��^�����=��=2R�ޓ��D� �7�b���F�I�.?��$>!�ʾ��M�s.<�hʾ����0ބ���T+̾�1��n��ɟ?I�A?u���r�V��	��W�����W?F���v���;�=5֯���=�>�>W�=���k3��nS�v�0?��?�&������g)>%����=m�+?�� ?lf}<�ܬ>]�%?�'�^K���]>�\5>���>�J�>Qv>\	���޽��?a�T?X���+3��[�>)��9x��Zp=0�>��3�e�׼-\>�U�<n����;� ٌ�0A�<�(W?��>Z�)����a��v���k==��x?��?�/�>�{k?c�B?2�<rf��}�S���Yiw=�W?�)i?ֺ>Ȇ���	оp���5�5?A�e?��N>\`h����{�.�ZU��#?��n?A_?�{���u}����g��Kn6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������_B�=�|�����? `�?󏦾.j<�R���l��*����9��=���Qqc����)�8���˾@w��)��%l�l�>�
@�=̽y��>}�.��߿mϿEV����ؾu�r���?i�>��ؽ�W��#�k�JOy�'�F�<B����"��>�N>�ɕ�i�����w�s]8��C���_�>ɛ���>�V�UI��H<��M�(<ђ�>T�>�ۃ>�<��%�����?=���/cο���	���S?Y�?;��?n� ?V�1<#�d��Di� $);
G?b$u?��[?���֯N� ��%�j?�_��vU`��4�tHE��U>�"3?�B�>T�-�V�|=�>���>g>�#/�y�Ŀ�ٶ�@���Z��?��?�o���>r��?ss+?�i�8���[����*�X�+��<A?�2>���I�!�B0=�UҒ�¼
?V~0?{�e.�O�_?��a���p�N�-���ƽݡ>%�0��b\�U �����We�����=y����?^�?r�?`��� #��5%?�>*����9ǾA �<���>i)�>�(N>vI_���u>����:�`h	>K��?�~�?j?g�������fW>C�}?���>��?mk�=�0�>2��=���E�+�>�#>"�=0<�<?�M?a��>
��=��6���.��F��*R�Ɗ��C�y*�>�b?��L?;�d>Ӵ�y�3�B� ��z˽�.�K�߼x�>��%��ݽ�5>�>>��>f�B�`�Ѿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?qQo���i�B>��?"������L��f?�
@u@a�^?*�̿<Ė�R�ھ$����H=,�=��">�r��<�K~=0�M�Y�f���f>j}�>��Z>pq>\NQ>w#x=��=����g!��㯿��0J�����*�����I�mԾ	�(��㾾{pv����������_�
����l<�˜���>%�U?�G?n�[?��>x�+]>˞��|^�Hͽfr>^�>��7?��C?��2?�"�=<u��%X_��'�����������>F	�>�W�>�P�>�X�>��¼-�u>
�{>�O�>p��=� �=�@=h.=t*a>	��>���>/�>�g>>��>Ӧ�����Y�h�z��̽���?˕���CJ�O핿���V���m;�=*�.?2q>)'��OIп�N����G?s㔾��ȹ0�_4>o�1?��W? �>a�� YO�C?>k�	�+Ni�3Q>���oj�+(�9:R>�B?��f>�u>w�3�Of8��P�/z��mn|>�36?T궾E?9��u��H�^ݾJM>ƾ>a�C�@i��������ti�ˈ{=�w:?��?,6���ܰ�_�u��A��HQR>Y6\>gd=�s�=�WM>s]c���ƽH��|.=���=�^>��?�,>Yd�=A�>�x��a�K����>y�D>�P.>�w@?�y%?����U��{����,��z>�g�>��>��>�EI�w�=���>h�a>����赀��R���>��X>��z��`��w�fz=.ᕽ�L�=R��=e� ��=�T�*=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾNh�>{x��Z�������u���#=R��>�8H?�V����O�f>��v
?�?�^�ߩ����ȿ4|v����>V�?���?i�m��A���@����>8��?�gY?qoi>�g۾:`Z����>Ի@?�R?�>�9�t�'���?�޶?֯�?�؉>0Ï?~c�?��?�>Uc��Ŀ����Y:I==1�=��4�MV���&�,I���� ���_�B���7���>Y��<v��>�#6�, ʾ9�-<�y�.v�f-����>`��>��=�%�>�Z�>��>�6">�^=���=k=���[[�c�O?�6�?�x�t/|�v���b�=2��]�>D�>ԭ@��D�#
�>�O?4X?Cte?x��>���xΗ�C�ȿ]	��tٽ�
�>?"�>?�(�>�
@>ľ���4ܷ>�G�>�]�=j�4}�aS�<���>/h:?��
?ˢV>�� ?a&?�0z>q0�>��>�σ����F�v��>�|�>�?B�?)B?@����6�Ȑ�9	5a�ڜ3>�`t?b�?���>_ߏ�����zY�?}���?ɽ옂?p�g?i�?��?��??��<?��s>˔�Z�Ҿ�����j>�V"?�_�WC@�e�%�F��i
?��?���> �}�R������7�X����N?��[?ߠ'?��!�`��k¾���<fA-���Ӏ�;�1���>�{>py���ٺ=.\>��=��l��2���<��=�ݓ>:�=+�5�wb���<,?}�G�ۃ���=J�r�/xD���>�IL>����^?m=���{�����x���
U�� �?Ǡ�?k�?���՝h��$=?-�?�	?B#�>+K��<~޾��<Qw�Dx��w���>���>ѵl���v��������F���Ž4 G����>V��>i?א0?�!a>5>�V��	�����!<�<�f�����A��8d��A��^�����l�s�*e��r���� 5>A��l_�>�.*?>v>�ј>���>,��<��>��t>~~>�J�>���>�Z�>s꙼v������KR?����'�'�|�辣���U3B?�qd?Z1�>$i�;��������?���?Js�?=v>�~h��,+�vn?�>�>"��+q
?MT:=3�M9�<BV��P���3��E�'��>|D׽� :��M�^nf�xj
?�/?���}�̾<;׽%�R�4�<&�?�J?D��IA��c�p4e�V�4��Fd�*U��8=����6�+���ߎ�����S���ྪm/>��?�_�?�B�� ��O\���E���f�l�>��\>\�>��>������������bW��8���5�7E'?�x?���>	;I?��4?��7?��S?2��>�J�>ky�����>�>�q�>]�	?ÎA?L#'?��=?�*?Cg?�>�U�4𾥛վ��?M�?�6?\=?
?�ꇾ��<�&=uD;�"���i���.>�)�<�܊�|�<<k5K=�|>-_?(v�j�8�q���:�j>��7?ϑ�>���>���p��O��<z�>f�
?H�>5����dr�BT�tN�>���?���١=T�)>�="���Һ�{�=�����=ɨ��_�;��5<s��=�=4�u��Z��7�:"�;"�<��?�	%?#9�>?y�>�Q���񾢩���׼ϨU>�x~>�n�=ܕ��6��q����7p���4>-ی?�G�?�U> O�=���=��þJn����9�u=��?�!?<�L?�Q�?��>?�^&?�>��{����\��]ӭ��?s!,?l��>|���ʾ�񨿁�3���?Z[?�<a���%;)��¾g�ԽQ�>s[/�/~����5D�#���������$��??�A���6��x辵����[����C?"�>KY�>��>�)�H�g�'%�@2;> ��>oR?$�>p�O?<{?��[?�jT>��8��0��ә�FL3�W�!>�@?&��?��?�y?pv�>��>�)�ྐྵU�������?߂�:W=�Z>���>6)�>��>���=��ǽ4X��a�>�O_�=ʍb>y��>���>��>4�w>Pc�<U�G?k��>I��%���餾-���6�;�W�u?۝�?��+?nq=1p���E�����X�>ho�?��?�*?��S����=�׼���Z�q��$�>��>]�>=�*G=\V>���>#��>n��U�pg8�]L���?�F?��=��ſ4r��u�6'��j͠;�y��ZD^������T`�|��=c����4�a����MW�8Н��B������)��lLz����>�l�=o��=l�=j��<{e�����<c-G=�c�<� =�[l��2�<��A�}��e��e1�0�}<��T=���˾��}?�;I?͕+?��C?f�y>2;>��3�@��>ᅂ��@?�V>�P�����
�;�%���� ��V�ؾ9x׾�c�ʟ��H>__I���>�83>�G�=>K�<��==s=�=gR�`=�$�=�O�=�g�=e��=��>sU>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�R>u��=Q�P��a4�v����%P��b,�#?Ӥ7���¾z̊>ֺ�=�̾.���2�y=��L>O�=��	�y Z����={Tg���A=a��=� �> TC>�R�=,�����=R\C<�d�=HS>��W��zM�`�d�v� =<�=��l>'�>���>��?;`0?Td?�4�>+�m��Ͼ�3���S�>�0�=uG�>��=7vB>ߐ�>&�7?t�D?��K?�z�>���=	�>��>Q�,���m�Yi��Ƨ���<2��?�Ά?Fθ>&�Q<��A����b>��Ž%z?�N1?]l?f�>d��r=��̟h���U�L�w�7��XX>�<�v�x��=��������>hx?$z?,b�>)�?�6(>��:>E��>���=�p�=P�⼃�L���5;E��=y�=��2>݁=�G�=�N�=WC����1��Ae<���<'�P=���= ��<YR�=���>3_9>^��>$ŧ=�꺾��>����G�`�<�举��B�.�a�v�����@������@>�('>�g��8䊿s��>(/�>*�m>��?9o?y��=tM ��lӾ__��SP���\p����=T��=JCv��A��W���S���龓��>SҎ>���>��o>+�N�>��k=��j
5���>�)���&�r��Rq��B�����05i�r%;��D?:󇿔��= �}?�H?(��?�d�>�Z����ؾb�->����=��<r�e��pg?�x&?�W�>����/D�N
̾񾽨
�>*�H�i�O�t�����0�׉"�ġ��k�>�
���о�*3�i`�����B���r�%�>��O?K׮?3�a�5Q���NO�#��$����.?G?g?F�>*T?�7?D��mG������=x�n?���?oE�?�_>�Ó=�ᨽԽ�>�r?9�? [�?}�h?�3�[?�>~�F�~��=󋤽���=�E�=��I=�ۜ=��>P��>�^�>�;X�E"�vf	��~�_����x׼ �>���>ʿ�>F_>EHH>lh>�6>C�>}��>��>�_>��>Է�>�N���T��V�>�z�=��>�+?�h�>GG>W��=[�UA�"���C�彘��c����=x�|�9�<G���� ?�rοـ?��>M��U"�>Sӣ��w�l��>e�&>���=�d?�=?>�\�=���>���>f��=">�>���>�FӾ7>����d!�m,C��R�_�Ѿ�}z>p���s
&���qw��vBI�un��qg�~j�D.��[<=�GȽ< H�?Լ��D�k�&�)�������? \�>�6?ڌ����2�>H��>;ȍ>fJ��&���ȍ��gᾰ�?.��?(ʊ>o�>�6o??�/?�5;���W
z�����Q22��cb��tb�Wf��mꋿմ�E�J�n�? \C?Ҭp?`k>>X�M>��?�W���9�>L��^��߰����><j�Ċ���`��������F�J>>kd?f��?��?F4��+ֻ�N>
�6?�%?1�?Z6B?��=?��(�?l3|>ͤ?��
?<7?�P4?�?~�Y>�>rN�V����	��96������FX���d���=
��=Ï�`(#=�Zs<�=iտ�4L�>B�=�Dּ�d�<^��=�٭=ڂ�=tޭ>ɭ`?�[�>¼�>TM<?��
���D��ݾ�)?梷=��������ƾ�+���6�=ӯS?]��?� f?�:�>*�<��~4���>��n>��>�~R>߸>�w߽�v.����=7:>)<2>�4�=��/��e��]Z�L�����;8
$>U��>�/|>�����'>�|��1z���d>��Q�
̺���S�g�G���1���v��X�>��K?�?��=_龘-���Hf�90)?,^<?:OM?��?��=:�۾��9���J��?���>�M�<������$��g�:�{��:��s>�1���-����T>R����澟�e�U�9���޾O}�<[�0�!=�k	���ѾN���"��=�; >4ȸ��$��I��]4���LL?�!�=�,���P�����u>>�>���>�����^L��*7�8���e\�=�2�>F%->	�\(��vF����C�>2KE?$V_?jk�?�)���s���B�����y��qȼ��?�^�>�g?P�A>�=����@�d��G��>J��>���X�G��5��1����$�8��>�<?t�>��?��R?�
?á`?�*?�5?u�>�6��S�1&?��?v�=�{ԽũT�H�8�8�E�|��>)?�B���>��?��?��&?�gQ?��?˭>w ��F@�!e�>'A�>ܛW��X��m�_>u�J?�B�>Y?ԃ?`�>>��5��䢾�|���3�=x�>��2?�)#?��?�Ը>?{�>XG�����=<��>T�b?g�?8p?)�=*)?�W2>�@�>n��=�7�>\��>l*?�>O?Xs?:�J?`��>���<5B����>q�\�I��VU;9�><�.w=���s����� �<���;�e��8�v�z�C������;�i�>&t>�����0>��ľ�P��o�@>!?��F��6����\:��V�=���>s?ާ�>�`#�蕒=g��>�C�>��&,(?��?$?C_+;��b���ھ��K���>@�A?Q�=��l�&�����u���g=��m?��^?5�W� !��Qq?;h?�\���f�����K�E��)b?ݝ?�]��5)�>�vS?҇??O�>�4��,�r�z���)�,<��j�=��>�3!��w�
ȝ>o�Y?ƥ�>�x�>ԋ=7�轐�y��
x���*??8�?z(�?�d�?.)>d�c�P��\ܾU��י5?��?K��Gy8?��y�W�v��P��Zt����޾��Ǿ����Z��^5������Z���߸a�J�Z��?@aM?6��?`<P?�"�}���Ixz�i1e���k�P�2�	����'�"�,��;O���t���!��_�;�d���>�O~��A��u�?'�'?�0��.�>@p��R��^�;5�B>@+��>��ﳞ=�ݎ�6|<=UDX=�!h�
�-�� ����?a�>��>�<?�[� !>���1���7������4>��>�(�>P'�>���:i.�I��{�ɾ�̄���ҽ��v>I�c?�dK?1�n?���"1�zU����!���,��w�� CD>\�>���>}�U�m8�/&�	!>��}r�M��ݐ�ܵ	�93�=��2?2�>!Ĝ>�6�??���꯾�kw���1�� p<���>��h?��>x��>Q�н� !�-��>ɤl?w��>�Q�>�Ԍ�!f!��{�xE˽��>�ǭ>��>�8o>Q#,�O:\��i���x���9����=�h?k����`��>e�Q?�kx:�0G<{V�>��v��!��s�K'�Su>'k?Ƃ�=-�:>�ž4�ۘ{��*��� )?ڜ?X��o�)�m}>)�!?��>�j�>xE�?hɜ>Ԫ����:�?�^?9�I?Է@?�I�>oP!=$���9 Ƚ��&���.=/��>#�Z>��n=Ž�=I���Z�?���D=�!�=L$��-�����;=M���_<��<M�5>T�ڿSXK��7ᾟ��S�W ������m�Ƚ�2�����p���Z������������?�F���q��q��C�d�J1�?���? ����������^�x!�lԨ>��}�PΓ����� ��LK�����3��0���X��lv��7l�
�'?玑�L�ǿ2����Mܾ� ?�0 ?��y?���z"�w�8��� >wQ�<a���w�ꗚ�|�ο������^?���>/�գ��'�>���>�WX>�eq>�O���۞�|(�<��?��-?�~�>.kr���ɿ8���S�<���?�@!~A?��(���쾺rV=Q��>\	?��?>�T1��P�����6�>2�?���?d�L=S�W�x$	���e?F�<�F��o޻���=�V�=�=:�NvJ>�{�>�o��]A�&�۽�y4>��>�"�ݿ��^���<zg]>@�ս� ���̈́?TA\�R�e�J&/����c�>�TT?��>	�=��+?>eH�6sϿ-H\�n�`?��?���?2-)?�<����>�ܾ�M?}6?Oə>�L'�h�t���=`׼��g��;�V����=z�>,�>{V.�%;�6P�Ę���.�=�� ��~ſ�l-��Q$�B��;����{����05���ƽ�����c�
�U�{�=��*>qDk>~kx>�3>��>N�_?��?0ס>Fd=E�����?]��{�Q�ߏO��M��_��}it�[���z��k�L�
�� 4��k8�2���G�F�X&=�	X�_א�g���b;��6�Ny?ŭ>
�Ͼ�E�Nm��2.��+V��h~�n�t��0��HH��>k�P�?��I? ��W�M�+)���>$+��#@?�kA�.��T���1	->k{Ƽ,���s>AȦ=]Q���@��
Z�ˮ5?2A)?%�־�ʛ�-��=5i����;�f?$��>��=��>u-?q��l��f�g>�>*��>���>5h)>w��@9��_.?0h?��׽�®�!�>p���.�[��>%��3>�x8��O)�X��>G9 �bVj���<ZF�����=�(W?e��>��)�<�Hb�����T==,�x?v�?�/�>={k?��B?�ޤ<Og����S���h]w=��W?�)i?7�>v���(о:����5?��e?�N>�fh����d�.��T��%?~�n?8_?K����v}������Co6?u�u?�7Z�$ꞿ����a>�:&�>O��>�P�>��8����>J�5?�
;�t���1���S�8��n�?�_@t��?� ����:��=??e]�>��8�mƾ�8ǽK���f=w��>_�����t�o�{}���8?�&�?G?1և���J�=4¦��ç?��?����q�<*���[_�`��XS���;�=Fh�+Q��ϳ���R:��yݾ
B��n����w'�>�b@ɒ����>��1��=��ο-����N%��ԗ
?��>|����B���>o���o�uB���;�Mc�Mr�>ߵ>���đ�ǋ{���;�������>�*
�'|�>�4T��u���h���,<�.�>@�>��>�����ƽ����?gz���'οz��P��<�X?Ҁ�? r�?�D?��@<�w�2�z����A�F?'Fs?�Y?�'�]�T�6���j?^^��OT`��4��HE�RU>�"3?�@�>0�-�~�|=�>h��>ai>n$/���Ŀ�ض������?g��?�o�*��>d��?s+?�i�b7��UZ����*���,��<A?2>،��<�!�
/=��Ԓ�!�
?�|0?�{��-���^?�)S�{�e��~&�;=�e�>6=������@ǽT2x�;Xa�����U��ܝ?���?��?����r�3V?V��>q����Ӿ�h�=w�7> K�>��>��K=jB>+]�FE5�6�.>���?H\�?y?�_��_a��=�=c�?J��>W�?��n=��>��]�P��1!ʼ�Ż���=�^�=ul?�a?z��>��H>]E�:#��j6��R-�\G�/H�	HZ>�G�?�f?y�>�9Ľ_�/=p&"������d�����=E�>��C�g.S=I5>9>��3>g�J�h����?Lp�9�ؿ j�� p'��54?.��>�?����t�����;_?Nz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>=�>�I�>D�Խ����[�����7>0�B?^��D��u�o�y�>���?
�@�ծ?ji�.	?�?������a~��M���7�g��=��5?kZ�u>6��>P�=k�v��䪿�Xt���>�?���?��>�$l?�n���B�U%=���>�{k?l�
?�S�����C>DI?��R����H��e? @��@�_?Iw���)ۿ�j��'j������l�<�d=-s,>���N�=��s���S�]�9��D=�>�>|Ze>�Ig>MH>��>o���'�#�����p����.�@c��g�%㎾o4��Ц�@���g▾�>���9=m2�<B>Q�RK1�k�ܽI{=��=P�W?4Q?��p?y��>��w��i#>�L �/KI=���L��=���>��.?T�O?�!)?w_�=L ��v�]�����w����悾k��>��:>?��>{��>�g�>v�<=+\>"�->P
t>
��=\�0=�����=�]O>� �>�w�>�/�>��'>6>u������lb��P��K½"l�?۟���;I�u���x}��Ok��`��=�*?�>V@��I�ѿ{z��̔I?�g��u�D!)�Z�>�95?�U?�>�����*�r�$>�|��!]���=c���e�qk(���G>�?~�V>H$j>�,8���6�#�I�>������>��4?�Ϻ�.�4�(o��G��0�<>5�>�3-����R햿Y����>]�-�G=*�:?��?iŽ�����z�����c>Z�V>�x�<h�j=��E>MrA��t��s�R�ߎT=���==hZ>o/?�)1>誘=�¤>Q]���xQ�W�>�<>M�,>��??��#?#�	�"���w����u/��{r> J�>(b�>��>�[K���=���>w�_>���������D?���X>��c�R]��e��K�=����ܧ�=��=_� ��b=���0=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾRh�>vx��Z�������u�f�#=M��>�8H?�V����O�b>��v
?�?�^�੤���ȿ6|v����>X�?���?f�m��A���@����>;��?�gY?woi>�g۾2`Z����>һ@?�R?�>�9�z�'���?�޶?կ�?^YI>at�?0�s?|��>�kz�On/���Y����oz=�^;{��>�M>�e���|F��ޓ��b��G�j�����a>؃$=��>�w��K��/��=L���C����e�Χ�>4q>�zJ>5�>� ?���>�V�>Nz=3Y�����Ŧ����`?��?��:�q����j�I5>���##?8�?U��>\����!y>�:q?��f?7�X?X�>�d'�&Z����ƿz%���X�<o�A>�N?��>᭽$ҷ>xP�-��>�x�>}��>�%�1uI��
;>�@�>��5?',?\Q>��/?�"?Æ	>�߄>fOc�`S��n�[�W��>G�>2Z�>�V?�Ҵ>?J���E1��+�������$g���=�U}?O�'?�`�>����,����m�@�>a�ɾ嵇?���?	�=~O?v&�?�]?�P?��>�-��R�_v��X�U>~!?)���HB��:&����>z	?~�?X��>����Eս��ͼ�������:?�{[?��%?����[a�88ľÝ�<!�,������<�P�.>f#>������=��>���=�p���6��u<|��=���>u��=K6����ly1?1^��b��9|>�8U��b���c> >����?hvܾ%�|����_��~*!���?�?{I�?�v#��9Q�d� ?���?�:?��
=𘆾�&۽� оĎ���N�=og*��JC>ꛯ>Ǘ<���#�,��Tݪ��]�q�/��Y����>���>r$?̝�>3��={��>B���C��W�"$���f�[���L�M�c�9��w��㒾h�ǽ��<�d���~Z��l�>s��N��>]��>4>I�t>}j�>�^�=@6�>��=̬e>5l�>m��=�%=�B�<R�0�ڽ�KR?����'�'����ֲ��]3B?�qd?B1�>9i�)��������?���?Os�?.=v>h��,+��n?�>�>Q��Nq
?U:=53�u;�<"V��H���3������>�D׽� :��M�
nf�fj
?�/?�����̾=;׽D�)�Zs�;O#s?W(5?��,Gc��V�V�.�\#}��P�uFѾ�޾D?�]���{���B���sg�����3�= ?#)�?�P��I���ڊ���|��h_�D>0��>i�=~L�>j�,>y�=��^�M�Yq��>���>-|?y��>��S?��6?H�T?q/?�.l>E��>��ѾH} ?���=o�>� ?f.?�<<?	�!?�}�>��?)mr>7�9�� �>L��T�'?��?�0%?Dp�>���>�-���@<J����\�7&���Ƚ(x�=� (=<p��k�H��~�<��>�W?T����8�����j>
�7?`��>���>g���*��U�<��>x�
?�D�>�  �K|r��b��S�>[��?��R�=%�)>���=���ҡҺ'Y�=4����=����t;�<J��=���=��t��1��cR�:h��;��<a=?[~?j*�>��>o���{���?����=��">�7?>ى�=9�߾jQ��N1���Of�|p>'�?�s�?D��=� �=,h�=�>���0��sF��R���.)=�%?l�?��Z?V��?��4?iS#?���=gs�N���'솿�i����?O�0?�u�>�.ھ�I���+�.;?I�>��X�#,x��J������^��5h>�� �*�z�Z��\�5�M�ݺ�Y�dџ����?���?�(���:��оa������92?��>���>j�>����g�!�?>U>���>o�Z?c�>3�O?n8{?8|[?0T>�j8�����N�������">�*@?��?��?Ny?bE�>�[>��)���߾Z:��H��5� w��#�T=��Y>`��>���>�˩>���=+�ƽ:g��73?�x��=,�a>n��>2U�>���>�7w>;�<FH?==�>�>������8�������o]��s?I��?�
&?���<�l��AC������>��?R-�?'�)?��P�N��=f!�K��9Pa��&�>.D�>��>���=��.={2%>�/�>�Y�>ߴ�#���9��e��V?C�D?I�=�$��t�N��="�Eؾܷ%>���>�;A���t븾�V=���~�����VP��?򢾬)'�:���$��=���?�w==�=��K>u�<%M<��>��P>%�Z�Pv>wy;�NԽ� ;��C�1�,���{����=գ1>RD&��VǾ�|?�<J?�6*?��@?�v>��>K�4����>��A�s?G�[>�������"�?�� ������pFԾ��Ѿ#\b��䠾�$>n)A�Z>�92>d�=�C�< T�=��r=�y�=����e*=��=NN�=e"�=���=�x	>p>��k?��C�Ft��"a���>|?X-����x����>#���&`������("���M?7r@�?&?1���>�~��/�V��$P>nH�;���=y��<�V�<�">�>&>�d�Mo��YM>�ɶ?c�
@Z�F?����ڜӿ�f�>(�>d��=�+_���0��!-��нf�ן?۟=�����~��>(�=�����iо���<��6>เ<РP�6�a�_
�=`�����=���=��|>��5>��=����p��=�q=���=>4\¼�|���Rl�<,��=,n>��>m��>8?�/?�c?0��>��s��о����S�>��=��>��l=vD>�>�8?F?2�L?�>u�=�'�>J	�>.�+�^�j�{�쾬8���V=#��?���?:4�>�{;��:�����W>��WнU�?�}/?��?E�>����c�`+����#g����׽�>�<��F��ۙ�0�뽧(��p(��J�=�m�>k�?P�>�.�>��m>
��>{/�>��9>�*����<n}�<��)<��;qW<���� =�KƼ��Q���'��m�ݽ/W=�V�<xr/���v=�[�=���>�$>��>�̊=]���H�0>pR���?N��)�=fi���B�� b�����/��S8�/�A>a�Y>��|������p?�Z>�`<>ov�?�s?�r>�-���Ծ������_��[V�X/�=�>"BA��^<�g�`�˲M��Ѿ%�>��>���>ʋm>�,,�o+?�4�x=<���5�i�>X⌾�T���'q��.���ٟ���h�:F���D?�+��`��=v~?�I?�?��>3����^ؾ�Q0>4���n=���ɟq�;֏���?֚&?
�>���D�@5ʾ������>�aG��N��ԕ�/:1��k������K�>r1���[ѾA�3�V���T���C�8wp�bĺ>jQ?o3�?�vV�����	P�UO�⿈�@ ?�c?��>|?�?7#�����x�����=a�o?��?Z��?G>b��=�����M�>�)	?ɳ�?���?��s?�.?�Z��>ϑ;�� >�-��I��=��>"{�=i�=Sb?��
?��
?P[��V�	���� �i^�.�<�ա=V��>|�>��r>��=��g=��=�&\>RȞ>��>��d>v�>MY�>J�����*��> �
>�R�>�iT?rn�>T4�=2��Z��<`ZL���w�P���<����ƽ����"��Wo���i��>#�ǿ6��?W+�>{	�7��>s��$]<��{>�#�=R�O��q�>T%>0Y_>���>��>��>>�߅>�4H>�iӾL>l��t!��	C��9R�֜Ѿ�z>몜��0&�ӓ�'W�� �I��~��b�*�i��0���e=�u&�<�H�?Q!����k���)��%��ߴ?O`�>z6?��������>��>�؍>u���G������ck�3��?���?���>FE�></&?v��>}� >�n��~%x����C�����v������tؔ�g�V�����`>?II�?F�?b��=xci>�Mh?K�`�Y?��ؾ�[8���Ǿ7a�>��i�|yԾ��>�ڡ����:<�>�؝?"�?�E?�s���=f-s>Axe?�?��>�ٞ>��<?K/�>�a?���>�66?6�B?��'?a�K?���>_N)=��}�I�߻Գ4>���c∾`�.�R̊��=!;�7<�"�=	>O�ü��
�71������� =i����?0=r�=�=<�<.L�=�&�>�rP?d�>�j>��V?��b���M���ξd?�ѽĄ��ػƾ�،�In��V>��?!��?.rV?�X=>���z�����=B�>��߼�t>b��>��<�Os��1�=���=$|S>ʵ>|�P�U~F����%�������kzZ>yU�>;t>c����i6>�i���0��hmV>��O��Kƾ8pm��FK���4�m�k��~�>�L?k!?i�=^p߾E�~b��$?9�:?��O?28l?6�z=Ԓ��U�3��I�9Q��}�>�u%=�-��S��N��K4C�q��t>Lf���ߠ��Tb>����q޾0�n��J�z��MFM=��iV=<�S�վ;,���=p&
>����� �����ժ��0J?!�j=�t���]U��s����>h>Pۮ>�:���v�G�@�����[?�=���>S�:>�i��?�~G��7��=�>oOE?yR_?�k�?�#��s���B����yo��LDǼ��?�b�>qj?��A>�ͭ=螱�X���d�G���>̝�>|��^�G�yC��h'��J�$�Ց�>Z>?%�>v�? �R?M�
?w�`?�*?m@?|�>j;��g� B&?6��?��=��Խ�T�� 9�JF����>|�)?�B�ܹ�>P�?�?��&?�Q?�?��>� ��C@��>�Y�>��W��b��>�_>��J?ٚ�>s=Y?�ԃ?y�=>]�5��颾�֩��U�=�>��2?6#?O�?���>5��>:�����=7��>|�b?>/�?��o?!$�=�	?�j2>���>ʸ�='��>���>d?8HO?P�s??�J?Zr�>���<����
���ws��FO�,��;!�H<��y=N��2�s�D��M>�<x�;O��0-��l�~D�m�����;���>-0t>�����5>�-þ�����B>#�ټĝ��/��\I=�ڥ�=Y�>���>(��>��%�	�=���>M��>M��J(?��?�?cBR�_c�Z׾�hM�%��>h�C?�A�=ߐm�f�ǅu��R=�m?YU\?�iW�����;�r?P�y?�s/�,@i�}e��BW�i��6`?((?֎�� ̳>3{?Ǻe?�?뱔�V^�����wIe��fM�/&>3��>v	8� a����>��^?d4f>-��>D�=0���Ḱ��N6�|� ?��?ٟ�?���?T�>�W~����<W�hs���7d?��>�2���Q ?q+�=�Q;�_Ǿ��J�P"������'���Ӕ�=������/.S��_=�;?Onf?�b?	G?g���b��H�;Qz��tX�����s��>�B�GC��uU��&z�������t���>FQ��pVB����?(B(?6f/���>(����b��ϾJ�?>񃟾�����=���(�I=�D=�{h�<31�2Э��� ?N�>��>�<?�I\���>��.�$�7������;>�H�>��>>�>ur��ɹ2����ʾ�]��j�Ͻ�9v>xc?��K?�n?\r��*1�K���$�!��/��a��4�B>Ql>���>��W����v9&��X>���r����w����	��~=��2?/)�>ﱜ>�O�??l{	��l��Iix���1�ҩ�<�1�>�i?T@�>1�>�н� ��H�>}Nl?��>o�>Gۋ��"��z�k�Խ�>�>�S�>���>�ti>��*�V�\�F���N���D8���=\�h?�񃾞�^�S�>`dQ?pZ"�<b<&g�>L�r�+}!�м���)�[>�?&r�=-6>��ľ����{�'+����)?U�?�i����)��Zy>��!?���>�Z�>p؃?[��>�&����{;�W?��_?�8J?>�@?r��>�=^ں�tʽ<�*���L=羉>6�]>Qi=�=�[�T&[���#�:�P='�=�d���=���x<�����H<�/=K%6>�yۿ
{K���ؾ������;
�v��C���Ƈ�b	�f>��	A���w��s��9%�q|V��c�B��'m�8q�?!��?���z؉�D���|��������>��r�<!}�Pӫ�=���ȕ�����Ҭ��m!���O��
i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾t1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@d|A?9�(�Q�쾸�U=I��>O�	?��?>�W1��F������M�>�9�?���?D�M=��W��l	��~e?�<M�F�2޻6��=)�=!�=���}J>�V�>�p��ZA��jܽ��4>��>rd"�Ś�[l^��	�<Sz]>�ս���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��={*�ªƿG#�T��L=m2�ۙU��.�r'��u�a�
��_�r��罧@g=�R�==6N>麄>��Q>�V>	1W?¬j?A�>۾>ʍ�o����k̾�ni�%(����t؉��{�D7������޾g	�П� �7ʾ� =�W�=7R�q���E� �_�b�U�F���.?5w$>R�ʾ��M�f�-<~pʾY����݄�᥽�-̾�1�"n�k͟?��A?������V�R��^V����f�W?P�ֻ��ꬾ���=_���u�=%�>���=���� 3��~S��h1?gN?�����Ȑ��0>N����+=k�(?D!?+��<J��>��%?�}�y���i�`>˵6>j�>���>'��=V设
���d"?|�V?�^�����_ޏ>zv����y��c=��>t� �����R�f>{�<����'�q��s��=)&W?���>y�)�� ��[���(��Y==I�x?-�?~#�>�wk?t�B?c6�<�n����S���.�w=��W?�)i?�>du���оDx��
�5?B�e?5�N>]vh�����.��S��?��n?\?�6��Rx}�������}p6?i�t?��\�����iY��wC�N¦>���>m��>�!:���>k�9?��%�\����G����5��џ?�@�g�?X��;s���z=�� ?n�>��X�ѺƾQ��������F=^��>Ff���+s�� ��1� :?:\�?���>��������=Pٕ�yZ�?��?烪��g<���#l��n���~�<+̫=��F"����}�7���ƾD�
�A���]տ����>"Z@gR轇*�>�D8�G6⿏SϿ���[о�Oq���?��>>�Ƚ��_�j�JPu���G���H�U����J�>��>����đ���{���;��4�����>���*�>��S��T��-m����.<
��>]��>"��>Yͮ�̥�����?H��M8ο2�����]�X?�^�?Zn�?�?cb:<�lv��,{�ׯ�=G?lms?OZ?I�&�H~]�E7�m�j?T^��'U`��4�EGE��U>�"3?�>�>��-��|=�>O��>Hf>�$/���ĿBٶ�h�����?���?�n꾋��>o��?Is+?�i�8��OX����*���,��>A?�2>X���s�!�0=�^Ԓ�B�
?e|0?/{��-�]�_?*�a�M�p���-���ƽ�ۡ>�0� f\�N�����Xe����@y����?M^�?h�?յ�� #�e6%?�>f����8Ǿ��<���>�(�>*N>bH_���u>����:�i	>���?�~�?Qj?���������U>
�}?�U�>Y�?{��=j/�>n"�=nҰ��.�z#>9q�=s�<�]�?�M?eu�>@��=?u8�7�.��HF�ER�?=�c�C����>b?��L?��b>[幽��1�G� ���ͽ1"2�O{�9P?�r�*��޽"#5>,�=>��>shD���Ҿ��?�o��ؿ
j���n'�t54?���>��?����t�����;_?Vy�>�6�
,���%���A�a��?�G�?7�?i�׾�[̼[>�>9J�> ս��������7>�B?c��D��<�o�G�>���?
�@�ծ?�i�d.?r��t\���v�
�����2��S�=V2?�Hml>�7�>4�=�Vx��ϩ��u����>R?�?��?w��>o�k?��n�VD��7=Eo�>��k?M�?��:��:aD>z�?�������hY��d?��
@ch@X_?+����տ!o��t_�t�����=*:5>t�>�=�D�=��HD���g����=�}�>Z��>smE>�>Vm�=�?>�*��`��.��k�z��-�nI����1Վ��������B,������о3�#�llG�����W��̉�.߫���h>��,?�??ԹZ?�Z�>{D��}�=\�-P�=e#���e5>�
�>E7K?�#p?'/2?P�>������\�!���૾�h? �>��>��>G�>@|>Əh>�8=��>dj>smw=o=p�M=�&>���>;��>ɖ�>�R<>w�>�д�f2����h���v�̽#�?Ry��ݶJ��0���3��͟���{�=�b.?U�>����>пy����/H?����((�(�+��>(�0?MbW?œ>���ȘT��,>���j��]>	 �eql���)�rQ>�e?��j>
_v>ϰ3�g28�|:Q��ܮ��z>S�4?A���2��6t��G��پ��R>%{�>�;�(���ɖ�����i�r�^=�l<?U�?i��0~��`Gt�����P>U>.�(=Gڷ=-�N>�J��ƽ՝G���-=��=��a>�P?�j2>*nb=8϶>)0���-���Y�>Y0>�M�=f�<?��?m4�������(�&�I�V>{��>ޘ�>-�!>�RB����=��>��d>�5~���ƽ!����o>�3.E>i�K<Q|��J˽��>'����0�=�֓=F*�e�<���K=�~?���(䈿��e���lD?R+?[ �=#�F<��"�D ���H��G�?r�@m�?��	��V�?�?�@�?��B��=}�>׫>�ξ�L��?��Ž6Ǣ�ʔ	�+)#�jS�?��?��/�Yʋ�<l�6>�^%?��ӾPh�>6x�zZ��~����u���#=���>�8H?�V��%�O�>��v
?�?�^�۩����ȿ0|v����>U�?���?F�m��A���@�[��>5��?rgY?�oi>]g۾=`Z�㋌>�@?�R?X�>�9���'�a�?�޶?ɯ�?'I>���?��s?�p�>8x�u^/��2��6���Q2=C^;�]�>�D>�����iF�Nד��g����j�����a>�$=�>�B��5���!�=5�B����f�ʦ�>�3q>*�I>*V�>g� ?bc�>��>�r=�����〾����
�e?���?oX�8������^�>*NP�T�?�U/?&�>�_��Bv�>u7[?:�y?��[?ݴ�>$��6ܟ���ǿ<����n�4
�>Z?C֩>"�(r2>�:������-P>Tx�>kl6��P���tf�K�p=��>i�#?g�>�$�<8G?0G%?Dm�=�d�>iyK��t��1Aо�x>$Y�>�P$?i�U?HJ�>�#B��2��a���ٝ���_���2>l�?TM)?~��>�痿* ���@	�~/o>I{���|�?���?MSB��>?��?�?
q�?�S>��9��� ������>��!?v���A�il&��l��?�=?
�>�7����Խ�,ؼ���N3��?'\?<&?̭�H@a��?þ/��<��#���X���<��H�>�>}�>���ؿ�=r>���=5�m��6��4f<��=(��>���=�n7�%ӏ�5�!?��C�z��%�*>�S���N�L�>\��=��޾�@?��Q��x�ʭ��ڞ�\����t?ٽ?�3�?��Իj�T��H@?>�?r'?���>��ݾ�z��=����R��I��C ��)���?��s����������C�|��31����}��>�Ʊ>�%?7��>>4h�%��>$�Ծc%<�{���<?�χv����?�S���)��������PU�F��=ఢ��lJ��x�>�vٽ�`E>��>�`�>E�>{�>}Y>uс>�c>ز>��>˛�="] >�a���L��s-��KR?�����'�w��˲��_3B?�qd?E1�>i�0��������?���?Us�?;=v>�~h��,+�qn?�>�>J��Dq
?�U:=%5�5<�<V��f���2������>�D׽� :��M�&nf�pj
?�/?����̾k;׽��о��5�kO�?�y?.n,���`���C�~W�?�j��A�o)��.ھ� ��t�=��Q���k}���(�85>�28?멠?F��t�G'&��G��0T�[G�=� ?��=��X>�'>ha5���&��
z����J���$?���?�Վ>�H?Vl;?��O?��J?N"�>z?�>�>���F�>�n<1ݡ>���>�.:?��.?Z0?@V?�i*?�\_>qk��n���[jپ�?)6?��?	�?W\?�k�����7���j:��jt�!m|�[c�=g �<�ؽ��s���Z='�U>�X?f��P�8�=����k>Ȁ7?_��>���>���G,����<��>�
?jF�> ��}r��b��V�>���?�����= �)>���=���f�Һ�\�=����V�=�1���{;�h^<���=��=]�t�5�����:8��;]s�<Y3�>��>�P�= B�>��1��>�����:< ���{���
;ˍ侖J��8���@�gB�>�Û?o�?�ޙ=��
>�w�=�Z��v��,������>�+�>�u�>P�I?z�?X�?�#?܃V=�c��Q��w[����׾�0?�,?w��>/��cEʾ�ը�t�3�J�?�?�:a�={�g>)��¾�Խ~�>�9/�k ~��诿{�C���t����g���&��?���?�WB���6�辰����V��U�C?���>���>=��>z�)���g����p:>�g�>��Q?�0�>I�O?�5{?�[?k<T>��8��(��iǙ�V�1���!>S@?ⵁ? ��?�#y?|��>b�>��)�� ྾_��\*��F󽽽����W=�$Z>���>0$�>A��>��=�(Ƚ����>��Q�=Jxb>,��>~��>���>ώw>d�<!�G?���>Jm��,��c6��N�����A��`u?/~�?�L+?��=���F�i��G��>}��?j�?�^*?�	T���=�ۼض�+q�cѷ>5��>M�>�j�=��C=7>��>���>>G��j�368��N���?��E?��=j+ҿ�Ł��9ʽ�-G���o<򕎾W�`�7�����}p9��]��/
s��ዾ�?�2n��X��K蹾!�þC���
Q	?�7@=f&?>5�!>�a��O-&��4�=QȽ�-��=�z��=g�L=�3��	�������'��[)�l�l��g˾�e}?8CI?ę+?�C?z>mR>T�1�U͖>�%���N?U�V>�WP�;c��5;�ͱ���3��^�ؾ6K׾B�c�����W>;�H��>�V3>hV�=ʈ<�,�=�Ir=C��=��k��Q=t[�=E��=�ì=��=V�>�7>b6w?=������4Q��V�s�:?\7�>�{�=3�ƾ�@?�>>�2��ԗ���b�q-?o��?U�?��?�ti��d�>����䎽Xu�=n���|<2>���=��2����>��J>���J��コ�34�?��@��??�ዿ��Ͽnb/>�7>d#>2�R�Љ1�?�\��b��~Z���!?�H;�J̾�6�>g�=,߾�ƾ��.=K�6>�nb=$g��V\���=��z���;=�l=�׉> �C>Xv�=,����=˜I=v��=0�O>�����7�a&,���3=d��=v�b>�&>���>�?O`0?]Yd?�5�>7n�Ͼ�B���D�> �=�A�>�ͅ=tB>���>��7?G�D?��K?���>Hʉ=d�>��>�,�p�m�
o徊ͧ��֬<薈?�͆?(׸>��Q<�A�N���f>�I?Žv?P1?yj?��>�����gQ �*��Ў��#9;�*=�e�J:l���7��-����H�=�	�>[��>���>�%p>re)>�F>�>�>��=mK�=D�	�HKr:B�˼�2=u�����<� Q�E���E>&<��G�����x!�J����M�e������=A��>��>K��>7�=�k����/>�����L��ڿ=$t��B@B��d�z^~���.� �6���B>x�X>;P�����0�?i\Z>5�?>�Y�?!�t?F� >tI��վe���e�1T�h1�=�_>��=��_;��l`���M�PIҾ)��>i�>{p�>�en>�+�{z?���{=��҂5���>��e�#����7qq�o����ߟ�z�h�]N��еD?��z>�=�1~?X�I?*��?{g�>锽��ؾ��/>PW����=eb��m�ꢔ�NK?��&?J�>���NfD�Z~Ӿam$�S��>��m���A��ܒ��2�_���,���VCb>�e���j߾ty<��˃�����J���o��l�>�Bd?]�?�ٽ]"���q]���˾��;d�>�J?%��>���>�C�>dG��h
�{�7�O+=�2}?!�?�O�?��>D��='��<�>�+	?���?ɸ�?��s?}x?�={�>ڢ�;h� >Y���0L�=V�>׋�=b*�="s?�
?��
?gj����	�������^����<�Ρ=���>�l�>��r>��=d�g=Xv�=l-\>ڞ>��>��d>l�>IP�>s륾	a��&?���=cO�>�2?�L�>{�W=+�����<�H���>��]*��ᵽ�߽'C�<�=���BN=��Ӽz��>Y�ǿ#Q�?5�T>�W��?�!��#�/��vS>XT>{Rݽ�S�>(�E>��}>�\�>T��>�>��>`�(>�MӾVX>A��VX!��,C���R��ѾWZz>䲜�c�%���������1I�fz���g�ij��,��;=�}-�<�G�?c���k���)�����b�?oR�>k6?�ь�*(���>���>ƴ�>�L��ꑕ��ƍ�Oiᾈ�?���?_��=��>1�#?�U>Jn>�F̽�y�FR��h$�5��+�v��3������zh��f�:[p?��?~�s?��'>[h�> �6?��@�8�v�$?b�����8�{\�=��>[�d����0���`���30��#>��? ��?��@?x�����=�q��ДG?��.?js?�"<?m��>֪�>�	R?'��>�he?��M?�?��7?݇2?�>i��w���V�|b�k$ӽ �=��ս�k=GS�����=�� <���<K'=�ʽ=?Jb��:�&���$=��<	J=]��=�g>,��>�1I?L8�>h8>�^?~c��_�^�_i���?�O����ƾ8���y7վIc	��>�V�?�r�?�7t?��=��������>޳>��<��>B�>R>�=M�����=��F>.gH>3mg;�����ѽ���8�a�i�����=z��>�E|>����l�)>pĢ�s�|�!xe>8�T�xa��CpS���G��2�$<v�	��>/�K?�B?P%�=�<�_w���e��.)?��<?�3M?� ?�؎=b*ھ�9�'�J��W��w�>���<;������� ���z:�����s>S����ߠ��Tb>����q޾0�n��J�z��MFM=��iV=<�S�վ;,���=p&
>����� �����ժ��0J?!�j=�t���]U��s����>h>Pۮ>�:���v�G�@�����[?�=���>S�:>�i��?�~G��7��=�>oOE?yR_?�k�?�#��s���B����yo��LDǼ��?�b�>qj?��A>�ͭ=螱�X���d�G���>̝�>|��^�G�yC��h'��J�$�Ց�>Z>?%�>v�? �R?M�
?w�`?�*?m@?|�>j;��g� B&?6��?��=��Խ�T�� 9�JF����>|�)?�B�ܹ�>P�?�?��&?�Q?�?��>� ��C@��>�Y�>��W��b��>�_>��J?ٚ�>s=Y?�ԃ?y�=>]�5��颾�֩��U�=�>��2?6#?O�?���>5��>:�����=7��>|�b?>/�?��o?!$�=�	?�j2>���>ʸ�='��>���>d?8HO?P�s??�J?Zr�>���<����
���ws��FO�,��;!�H<��y=N��2�s�D��M>�<x�;O��0-��l�~D�m�����;���>-0t>�����5>�-þ�����B>#�ټĝ��/��\I=�ڥ�=Y�>���>(��>��%�	�=���>M��>M��J(?��?�?cBR�_c�Z׾�hM�%��>h�C?�A�=ߐm�f�ǅu��R=�m?YU\?�iW�����;�r?P�y?�s/�,@i�}e��BW�i��6`?((?֎�� ̳>3{?Ǻe?�?뱔�V^�����wIe��fM�/&>3��>v	8� a����>��^?d4f>-��>D�=0���Ḱ��N6�|� ?��?ٟ�?���?T�>�W~����<W�hs���7d?��>�2���Q ?q+�=�Q;�_Ǿ��J�P"������'���Ӕ�=������/.S��_=�;?Onf?�b?	G?g���b��H�;Qz��tX�����s��>�B�GC��uU��&z�������t���>FQ��pVB����?(B(?6f/���>(����b��ϾJ�?>񃟾�����=���(�I=�D=�{h�<31�2Э��� ?N�>��>�<?�I\���>��.�$�7������;>�H�>��>>�>ur��ɹ2����ʾ�]��j�Ͻ�9v>xc?��K?�n?\r��*1�K���$�!��/��a��4�B>Ql>���>��W����v9&��X>���r����w����	��~=��2?/)�>ﱜ>�O�??l{	��l��Iix���1�ҩ�<�1�>�i?T@�>1�>�н� ��H�>}Nl?��>o�>Gۋ��"��z�k�Խ�>�>�S�>���>�ti>��*�V�\�F���N���D8���=\�h?�񃾞�^�S�>`dQ?pZ"�<b<&g�>L�r�+}!�м���)�[>�?&r�=-6>��ľ����{�'+����)?U�?�i����)��Zy>��!?���>�Z�>p؃?[��>�&����{;�W?��_?�8J?>�@?r��>�=^ں�tʽ<�*���L=羉>6�]>Qi=�=�[�T&[���#�:�P='�=�d���=���x<�����H<�/=K%6>�yۿ
{K���ؾ������;
�v��C���Ƈ�b	�f>��	A���w��s��9%�q|V��c�B��'m�8q�?!��?���z؉�D���|��������>��r�<!}�Pӫ�=���ȕ�����Ҭ��m!���O��
i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾t1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@d|A?9�(�Q�쾸�U=I��>O�	?��?>�W1��F������M�>�9�?���?D�M=��W��l	��~e?�<M�F�2޻6��=)�=!�=���}J>�V�>�p��ZA��jܽ��4>��>rd"�Ś�[l^��	�<Sz]>�ս���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��={*�ªƿG#�T��L=m2�ۙU��.�r'��u�a�
��_�r��罧@g=�R�==6N>麄>��Q>�V>	1W?¬j?A�>۾>ʍ�o����k̾�ni�%(����t؉��{�D7������޾g	�П� �7ʾ� =�W�=7R�q���E� �_�b�U�F���.?5w$>R�ʾ��M�f�-<~pʾY����݄�᥽�-̾�1�"n�k͟?��A?������V�R��^V����f�W?P�ֻ��ꬾ���=_���u�=%�>���=���� 3��~S��h1?gN?�����Ȑ��0>N����+=k�(?D!?+��<J��>��%?�}�y���i�`>˵6>j�>���>'��=V设
���d"?|�V?�^�����_ޏ>zv����y��c=��>t� �����R�f>{�<����'�q��s��=)&W?���>y�)�� ��[���(��Y==I�x?-�?~#�>�wk?t�B?c6�<�n����S���.�w=��W?�)i?�>du���оDx��
�5?B�e?5�N>]vh�����.��S��?��n?\?�6��Rx}�������}p6?i�t?��\�����iY��wC�N¦>���>m��>�!:���>k�9?��%�\����G����5��џ?�@�g�?X��;s���z=�� ?n�>��X�ѺƾQ��������F=^��>Ff���+s�� ��1� :?:\�?���>��������=Pٕ�yZ�?��?烪��g<���#l��n���~�<+̫=��F"����}�7���ƾD�
�A���]տ����>"Z@gR轇*�>�D8�G6⿏SϿ���[о�Oq���?��>>�Ƚ��_�j�JPu���G���H�U����J�>��>����đ���{���;��4�����>���*�>��S��T��-m����.<
��>]��>"��>Yͮ�̥�����?H��M8ο2�����]�X?�^�?Zn�?�?cb:<�lv��,{�ׯ�=G?lms?OZ?I�&�H~]�E7�m�j?T^��'U`��4�EGE��U>�"3?�>�>��-��|=�>O��>Hf>�$/���ĿBٶ�h�����?���?�n꾋��>o��?Is+?�i�8��OX����*���,��>A?�2>X���s�!�0=�^Ԓ�B�
?e|0?/{��-�]�_?*�a�M�p���-���ƽ�ۡ>�0� f\�N�����Xe����@y����?M^�?h�?յ�� #�e6%?�>f����8Ǿ��<���>�(�>*N>bH_���u>����:�i	>���?�~�?Qj?���������U>
�}?�U�>Y�?{��=j/�>n"�=nҰ��.�z#>9q�=s�<�]�?�M?eu�>@��=?u8�7�.��HF�ER�?=�c�C����>b?��L?��b>[幽��1�G� ���ͽ1"2�O{�9P?�r�*��޽"#5>,�=>��>shD���Ҿ��?�o��ؿ
j���n'�t54?���>��?����t�����;_?Vy�>�6�
,���%���A�a��?�G�?7�?i�׾�[̼[>�>9J�> ս��������7>�B?c��D��<�o�G�>���?
�@�ծ?�i�d.?r��t\���v�
�����2��S�=V2?�Hml>�7�>4�=�Vx��ϩ��u����>R?�?��?w��>o�k?��n�VD��7=Eo�>��k?M�?��:��:aD>z�?�������hY��d?��
@ch@X_?+����տ!o��t_�t�����=*:5>t�>�=�D�=��HD���g����=�}�>Z��>smE>�>Vm�=�?>�*��`��.��k�z��-�nI����1Վ��������B,������о3�#�llG�����W��̉�.߫���h>��,?�??ԹZ?�Z�>{D��}�=\�-P�=e#���e5>�
�>E7K?�#p?'/2?P�>������\�!���૾�h? �>��>��>G�>@|>Əh>�8=��>dj>smw=o=p�M=�&>���>;��>ɖ�>�R<>w�>�д�f2����h���v�̽#�?Ry��ݶJ��0���3��͟���{�=�b.?U�>����>пy����/H?����((�(�+��>(�0?MbW?œ>���ȘT��,>���j��]>	 �eql���)�rQ>�e?��j>
_v>ϰ3�g28�|:Q��ܮ��z>S�4?A���2��6t��G��پ��R>%{�>�;�(���ɖ�����i�r�^=�l<?U�?i��0~��`Gt�����P>U>.�(=Gڷ=-�N>�J��ƽ՝G���-=��=��a>�P?�j2>*nb=8϶>)0���-���Y�>Y0>�M�=f�<?��?m4�������(�&�I�V>{��>ޘ�>-�!>�RB����=��>��d>�5~���ƽ!����o>�3.E>i�K<Q|��J˽��>'����0�=�֓=F*�e�<���K=�~?���(䈿��e���lD?R+?[ �=#�F<��"�D ���H��G�?r�@m�?��	��V�?�?�@�?��B��=}�>׫>�ξ�L��?��Ž6Ǣ�ʔ	�+)#�jS�?��?��/�Yʋ�<l�6>�^%?��ӾPh�>6x�zZ��~����u���#=���>�8H?�V��%�O�>��v
?�?�^�۩����ȿ0|v����>U�?���?F�m��A���@�[��>5��?rgY?�oi>]g۾=`Z�㋌>�@?�R?X�>�9���'�a�?�޶?ɯ�?'I>���?��s?�p�>8x�u^/��2��6���Q2=C^;�]�>�D>�����iF�Nד��g����j�����a>�$=�>�B��5���!�=5�B����f�ʦ�>�3q>*�I>*V�>g� ?bc�>��>�r=�����〾����
�e?���?oX�8������^�>*NP�T�?�U/?&�>�_��Bv�>u7[?:�y?��[?ݴ�>$��6ܟ���ǿ<����n�4
�>Z?C֩>"�(r2>�:������-P>Tx�>kl6��P���tf�K�p=��>i�#?g�>�$�<8G?0G%?Dm�=�d�>iyK��t��1Aо�x>$Y�>�P$?i�U?HJ�>�#B��2��a���ٝ���_���2>l�?TM)?~��>�痿* ���@	�~/o>I{���|�?���?MSB��>?��?�?
q�?�S>��9��� ������>��!?v���A�il&��l��?�=?
�>�7����Խ�,ؼ���N3��?'\?<&?̭�H@a��?þ/��<��#���X���<��H�>�>}�>���ؿ�=r>���=5�m��6��4f<��=(��>���=�n7�%ӏ�5�!?��C�z��%�*>�S���N�L�>\��=��޾�@?��Q��x�ʭ��ڞ�\����t?ٽ?�3�?��Իj�T��H@?>�?r'?���>��ݾ�z��=����R��I��C ��)���?��s����������C�|��31����}��>�Ʊ>�%?7��>>4h�%��>$�Ծc%<�{���<?�χv����?�S���)��������PU�F��=ఢ��lJ��x�>�vٽ�`E>��>�`�>E�>{�>}Y>uс>�c>ز>��>˛�="] >�a���L��s-��KR?�����'�w��˲��_3B?�qd?E1�>i�0��������?���?Us�?;=v>�~h��,+�qn?�>�>J��Dq
?�U:=%5�5<�<V��f���2������>�D׽� :��M�&nf�pj
?�/?����̾k;׽��о��5�kO�?�y?.n,���`���C�~W�?�j��A�o)��.ھ� ��t�=��Q���k}���(�85>�28?멠?F��t�G'&��G��0T�[G�=� ?��=��X>�'>ha5���&��
z����J���$?���?�Վ>�H?Vl;?��O?��J?N"�>z?�>�>���F�>�n<1ݡ>���>�.:?��.?Z0?@V?�i*?�\_>qk��n���[jپ�?)6?��?	�?W\?�k�����7���j:��jt�!m|�[c�=g �<�ؽ��s���Z='�U>�X?f��P�8�=����k>Ȁ7?_��>���>���G,����<��>�
?jF�> ��}r��b��V�>���?�����= �)>���=���f�Һ�\�=����V�=�1���{;�h^<���=��=]�t�5�����:8��;]s�<Y3�>��>�P�= B�>��1��>�����:< ���{���
;ˍ侖J��8���@�gB�>�Û?o�?�ޙ=��
>�w�=�Z��v��,������>�+�>�u�>P�I?z�?X�?�#?܃V=�c��Q��w[����׾�0?�,?w��>/��cEʾ�ը�t�3�J�?�?�:a�={�g>)��¾�Խ~�>�9/�k ~��诿{�C���t����g���&��?���?�WB���6�辰����V��U�C?���>���>=��>z�)���g����p:>�g�>��Q?�0�>I�O?�5{?�[?k<T>��8��(��iǙ�V�1���!>S@?ⵁ? ��?�#y?|��>b�>��)�� ྾_��\*��F󽽽����W=�$Z>���>0$�>A��>��=�(Ƚ����>��Q�=Jxb>,��>~��>���>ώw>d�<!�G?���>Jm��,��c6��N�����A��`u?/~�?�L+?��=���F�i��G��>}��?j�?�^*?�	T���=�ۼض�+q�cѷ>5��>M�>�j�=��C=7>��>���>>G��j�368��N���?��E?��=j+ҿ�Ł��9ʽ�-G���o<򕎾W�`�7�����}p9��]��/
s��ዾ�?�2n��X��K蹾!�þC���
Q	?�7@=f&?>5�!>�a��O-&��4�=QȽ�-��=�z��=g�L=�3��	�������'��[)�l�l��g˾�e}?8CI?ę+?�C?z>mR>T�1�U͖>�%���N?U�V>�WP�;c��5;�ͱ���3��^�ؾ6K׾B�c�����W>;�H��>�V3>hV�=ʈ<�,�=�Ir=C��=��k��Q=t[�=E��=�ì=��=V�>�7>b6w?=������4Q��V�s�:?\7�>�{�=3�ƾ�@?�>>�2��ԗ���b�q-?o��?U�?��?�ti��d�>����䎽Xu�=n���|<2>���=��2����>��J>���J��コ�34�?��@��??�ዿ��Ͽnb/>�7>d#>2�R�Љ1�?�\��b��~Z���!?�H;�J̾�6�>g�=,߾�ƾ��.=K�6>�nb=$g��V\���=��z���;=�l=�׉> �C>Xv�=,����=˜I=v��=0�O>�����7�a&,���3=d��=v�b>�&>���>�?O`0?]Yd?�5�>7n�Ͼ�B���D�> �=�A�>�ͅ=tB>���>��7?G�D?��K?���>Hʉ=d�>��>�,�p�m�
o徊ͧ��֬<薈?�͆?(׸>��Q<�A�N���f>�I?Žv?P1?yj?��>�����gQ �*��Ў��#9;�*=�e�J:l���7��-����H�=�	�>[��>���>�%p>re)>�F>�>�>��=mK�=D�	�HKr:B�˼�2=u�����<� Q�E���E>&<��G�����x!�J����M�e������=A��>��>K��>7�=�k����/>�����L��ڿ=$t��B@B��d�z^~���.� �6���B>x�X>;P�����0�?i\Z>5�?>�Y�?!�t?F� >tI��վe���e�1T�h1�=�_>��=��_;��l`���M�PIҾ)��>i�>{p�>�en>�+�{z?���{=��҂5���>��e�#����7qq�o����ߟ�z�h�]N��еD?��z>�=�1~?X�I?*��?{g�>锽��ؾ��/>PW����=eb��m�ꢔ�NK?��&?J�>���NfD�Z~Ӿam$�S��>��m���A��ܒ��2�_���,���VCb>�e���j߾ty<��˃�����J���o��l�>�Bd?]�?�ٽ]"���q]���˾��;d�>�J?%��>���>�C�>dG��h
�{�7�O+=�2}?!�?�O�?��>D��='��<�>�+	?���?ɸ�?��s?}x?�={�>ڢ�;h� >Y���0L�=V�>׋�=b*�="s?�
?��
?gj����	�������^����<�Ρ=���>�l�>��r>��=d�g=Xv�=l-\>ڞ>��>��d>l�>IP�>s륾	a��&?���=cO�>�2?�L�>{�W=+�����<�H���>��]*��ᵽ�߽'C�<�=���BN=��Ӽz��>Y�ǿ#Q�?5�T>�W��?�!��#�/��vS>XT>{Rݽ�S�>(�E>��}>�\�>T��>�>��>`�(>�MӾVX>A��VX!��,C���R��ѾWZz>䲜�c�%���������1I�fz���g�ij��,��;=�}-�<�G�?c���k���)�����b�?oR�>k6?�ь�*(���>���>ƴ�>�L��ꑕ��ƍ�Oiᾈ�?���?_��=��>1�#?�U>Jn>�F̽�y�FR��h$�5��+�v��3������zh��f�:[p?��?~�s?��'>[h�> �6?��@�8�v�$?b�����8�{\�=��>[�d����0���`���30��#>��? ��?��@?x�����=�q��ДG?��.?js?�"<?m��>֪�>�	R?'��>�he?��M?�?��7?݇2?�>i��w���V�|b�k$ӽ �=��ս�k=GS�����=�� <���<K'=�ʽ=?Jb��:�&���$=��<	J=]��=�g>,��>�1I?L8�>h8>�^?~c��_�^�_i���?�O����ƾ8���y7վIc	��>�V�?�r�?�7t?��=��������>޳>��<��>B�>R>�=M�����=��F>.gH>3mg;�����ѽ���8�a�i�����=z��>�E|>����l�)>pĢ�s�|�!xe>8�T�xa��CpS���G��2�$<v�	��>/�K?�B?P%�=�<�_w���e��.)?��<?�3M?� ?�؎=b*ھ�9�'�J��W��w�>���<;������� ���z:�����s>S����ߠ��Tb>����q޾0�n��J�z��MFM=��iV=<�S�վ;,���=p&
>����� �����ժ��0J?!�j=�t���]U��s����>h>Pۮ>�:���v�G�@�����[?�=���>S�:>�i��?�~G��7��=�>oOE?yR_?�k�?�#��s���B����yo��LDǼ��?�b�>qj?��A>�ͭ=螱�X���d�G���>̝�>|��^�G�yC��h'��J�$�Ց�>Z>?%�>v�? �R?M�
?w�`?�*?m@?|�>j;��g� B&?6��?��=��Խ�T�� 9�JF����>|�)?�B�ܹ�>P�?�?��&?�Q?�?��>� ��C@��>�Y�>��W��b��>�_>��J?ٚ�>s=Y?�ԃ?y�=>]�5��颾�֩��U�=�>��2?6#?O�?���>5��>:�����=7��>|�b?>/�?��o?!$�=�	?�j2>���>ʸ�='��>���>d?8HO?P�s??�J?Zr�>���<����
���ws��FO�,��;!�H<��y=N��2�s�D��M>�<x�;O��0-��l�~D�m�����;���>-0t>�����5>�-þ�����B>#�ټĝ��/��\I=�ڥ�=Y�>���>(��>��%�	�=���>M��>M��J(?��?�?cBR�_c�Z׾�hM�%��>h�C?�A�=ߐm�f�ǅu��R=�m?YU\?�iW�����;�r?P�y?�s/�,@i�}e��BW�i��6`?((?֎�� ̳>3{?Ǻe?�?뱔�V^�����wIe��fM�/&>3��>v	8� a����>��^?d4f>-��>D�=0���Ḱ��N6�|� ?��?ٟ�?���?T�>�W~����<W�hs���7d?��>�2���Q ?q+�=�Q;�_Ǿ��J�P"������'���Ӕ�=������/.S��_=�;?Onf?�b?	G?g���b��H�;Qz��tX�����s��>�B�GC��uU��&z�������t���>FQ��pVB����?(B(?6f/���>(����b��ϾJ�?>񃟾�����=���(�I=�D=�{h�<31�2Э��� ?N�>��>�<?�I\���>��.�$�7������;>�H�>��>>�>ur��ɹ2����ʾ�]��j�Ͻ�9v>xc?��K?�n?\r��*1�K���$�!��/��a��4�B>Ql>���>��W����v9&��X>���r����w����	��~=��2?/)�>ﱜ>�O�??l{	��l��Iix���1�ҩ�<�1�>�i?T@�>1�>�н� ��H�>}Nl?��>o�>Gۋ��"��z�k�Խ�>�>�S�>���>�ti>��*�V�\�F���N���D8���=\�h?�񃾞�^�S�>`dQ?pZ"�<b<&g�>L�r�+}!�м���)�[>�?&r�=-6>��ľ����{�'+����)?U�?�i����)��Zy>��!?���>�Z�>p؃?[��>�&����{;�W?��_?�8J?>�@?r��>�=^ں�tʽ<�*���L=羉>6�]>Qi=�=�[�T&[���#�:�P='�=�d���=���x<�����H<�/=K%6>�yۿ
{K���ؾ������;
�v��C���Ƈ�b	�f>��	A���w��s��9%�q|V��c�B��'m�8q�?!��?���z؉�D���|��������>��r�<!}�Pӫ�=���ȕ�����Ҭ��m!���O��
i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾t1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@d|A?9�(�Q�쾸�U=I��>O�	?��?>�W1��F������M�>�9�?���?D�M=��W��l	��~e?�<M�F�2޻6��=)�=!�=���}J>�V�>�p��ZA��jܽ��4>��>rd"�Ś�[l^��	�<Sz]>�ս���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��={*�ªƿG#�T��L=m2�ۙU��.�r'��u�a�
��_�r��罧@g=�R�==6N>麄>��Q>�V>	1W?¬j?A�>۾>ʍ�o����k̾�ni�%(����t؉��{�D7������޾g	�П� �7ʾ� =�W�=7R�q���E� �_�b�U�F���.?5w$>R�ʾ��M�f�-<~pʾY����݄�᥽�-̾�1�"n�k͟?��A?������V�R��^V����f�W?P�ֻ��ꬾ���=_���u�=%�>���=���� 3��~S��h1?gN?�����Ȑ��0>N����+=k�(?D!?+��<J��>��%?�}�y���i�`>˵6>j�>���>'��=V设
���d"?|�V?�^�����_ޏ>zv����y��c=��>t� �����R�f>{�<����'�q��s��=)&W?���>y�)�� ��[���(��Y==I�x?-�?~#�>�wk?t�B?c6�<�n����S���.�w=��W?�)i?�>du���оDx��
�5?B�e?5�N>]vh�����.��S��?��n?\?�6��Rx}�������}p6?i�t?��\�����iY��wC�N¦>���>m��>�!:���>k�9?��%�\����G����5��џ?�@�g�?X��;s���z=�� ?n�>��X�ѺƾQ��������F=^��>Ff���+s�� ��1� :?:\�?���>��������=Pٕ�yZ�?��?烪��g<���#l��n���~�<+̫=��F"����}�7���ƾD�
�A���]տ����>"Z@gR轇*�>�D8�G6⿏SϿ���[о�Oq���?��>>�Ƚ��_�j�JPu���G���H�U����J�>��>����đ���{���;��4�����>���*�>��S��T��-m����.<
��>]��>"��>Yͮ�̥�����?H��M8ο2�����]�X?�^�?Zn�?�?cb:<�lv��,{�ׯ�=G?lms?OZ?I�&�H~]�E7�m�j?T^��'U`��4�EGE��U>�"3?�>�>��-��|=�>O��>Hf>�$/���ĿBٶ�h�����?���?�n꾋��>o��?Is+?�i�8��OX����*���,��>A?�2>X���s�!�0=�^Ԓ�B�
?e|0?/{��-�]�_?*�a�M�p���-���ƽ�ۡ>�0� f\�N�����Xe����@y����?M^�?h�?յ�� #�e6%?�>f����8Ǿ��<���>�(�>*N>bH_���u>����:�i	>���?�~�?Qj?���������U>
�}?�U�>Y�?{��=j/�>n"�=nҰ��.�z#>9q�=s�<�]�?�M?eu�>@��=?u8�7�.��HF�ER�?=�c�C����>b?��L?��b>[幽��1�G� ���ͽ1"2�O{�9P?�r�*��޽"#5>,�=>��>shD���Ҿ��?�o��ؿ
j���n'�t54?���>��?����t�����;_?Vy�>�6�
,���%���A�a��?�G�?7�?i�׾�[̼[>�>9J�> ս��������7>�B?c��D��<�o�G�>���?
�@�ծ?�i�d.?r��t\���v�
�����2��S�=V2?�Hml>�7�>4�=�Vx��ϩ��u����>R?�?��?w��>o�k?��n�VD��7=Eo�>��k?M�?��:��:aD>z�?�������hY��d?��
@ch@X_?+����տ!o��t_�t�����=*:5>t�>�=�D�=��HD���g����=�}�>Z��>smE>�>Vm�=�?>�*��`��.��k�z��-�nI����1Վ��������B,������о3�#�llG�����W��̉�.߫���h>��,?�??ԹZ?�Z�>{D��}�=\�-P�=e#���e5>�
�>E7K?�#p?'/2?P�>������\�!���૾�h? �>��>��>G�>@|>Əh>�8=��>dj>smw=o=p�M=�&>���>;��>ɖ�>�R<>w�>�д�f2����h���v�̽#�?Ry��ݶJ��0���3��͟���{�=�b.?U�>����>пy����/H?����((�(�+��>(�0?MbW?œ>���ȘT��,>���j��]>	 �eql���)�rQ>�e?��j>
_v>ϰ3�g28�|:Q��ܮ��z>S�4?A���2��6t��G��پ��R>%{�>�;�(���ɖ�����i�r�^=�l<?U�?i��0~��`Gt�����P>U>.�(=Gڷ=-�N>�J��ƽ՝G���-=��=��a>�P?�j2>*nb=8϶>)0���-���Y�>Y0>�M�=f�<?��?m4�������(�&�I�V>{��>ޘ�>-�!>�RB����=��>��d>�5~���ƽ!����o>�3.E>i�K<Q|��J˽��>'����0�=�֓=F*�e�<���K=�~?���(䈿��e���lD?R+?[ �=#�F<��"�D ���H��G�?r�@m�?��	��V�?�?�@�?��B��=}�>׫>�ξ�L��?��Ž6Ǣ�ʔ	�+)#�jS�?��?��/�Yʋ�<l�6>�^%?��ӾPh�>6x�zZ��~����u���#=���>�8H?�V��%�O�>��v
?�?�^�۩����ȿ0|v����>U�?���?F�m��A���@�[��>5��?rgY?�oi>]g۾=`Z�㋌>�@?�R?X�>�9���'�a�?�޶?ɯ�?'I>���?��s?�p�>8x�u^/��2��6���Q2=C^;�]�>�D>�����iF�Nד��g����j�����a>�$=�>�B��5���!�=5�B����f�ʦ�>�3q>*�I>*V�>g� ?bc�>��>�r=�����〾����
�e?���?oX�8������^�>*NP�T�?�U/?&�>�_��Bv�>u7[?:�y?��[?ݴ�>$��6ܟ���ǿ<����n�4
�>Z?C֩>"�(r2>�:������-P>Tx�>kl6��P���tf�K�p=��>i�#?g�>�$�<8G?0G%?Dm�=�d�>iyK��t��1Aо�x>$Y�>�P$?i�U?HJ�>�#B��2��a���ٝ���_���2>l�?TM)?~��>�痿* ���@	�~/o>I{���|�?���?MSB��>?��?�?
q�?�S>��9��� ������>��!?v���A�il&��l��?�=?
�>�7����Խ�,ؼ���N3��?'\?<&?̭�H@a��?þ/��<��#���X���<��H�>�>}�>���ؿ�=r>���=5�m��6��4f<��=(��>���=�n7�%ӏ�5�!?��C�z��%�*>�S���N�L�>\��=��޾�@?��Q��x�ʭ��ڞ�\����t?ٽ?�3�?��Իj�T��H@?>�?r'?���>��ݾ�z��=����R��I��C ��)���?��s����������C�|��31����}��>�Ʊ>�%?7��>>4h�%��>$�Ծc%<�{���<?�χv����?�S���)��������PU�F��=ఢ��lJ��x�>�vٽ�`E>��>�`�>E�>{�>}Y>uс>�c>ز>��>˛�="] >�a���L��s-��KR?�����'�w��˲��_3B?�qd?E1�>i�0��������?���?Us�?;=v>�~h��,+�qn?�>�>J��Dq
?�U:=%5�5<�<V��f���2������>�D׽� :��M�&nf�pj
?�/?����̾k;׽��о��5�kO�?�y?.n,���`���C�~W�?�j��A�o)��.ھ� ��t�=��Q���k}���(�85>�28?멠?F��t�G'&��G��0T�[G�=� ?��=��X>�'>ha5���&��
z����J���$?���?�Վ>�H?Vl;?��O?��J?N"�>z?�>�>���F�>�n<1ݡ>���>�.:?��.?Z0?@V?�i*?�\_>qk��n���[jپ�?)6?��?	�?W\?�k�����7���j:��jt�!m|�[c�=g �<�ؽ��s���Z='�U>�X?f��P�8�=����k>Ȁ7?_��>���>���G,����<��>�
?jF�> ��}r��b��V�>���?�����= �)>���=���f�Һ�\�=����V�=�1���{;�h^<���=��=]�t�5�����:8��;]s�<Y3�>��>�P�= B�>��1��>�����:< ���{���
;ˍ侖J��8���@�gB�>�Û?o�?�ޙ=��
>�w�=�Z��v��,������>�+�>�u�>P�I?z�?X�?�#?܃V=�c��Q��w[����׾�0?�,?w��>/��cEʾ�ը�t�3�J�?�?�:a�={�g>)��¾�Խ~�>�9/�k ~��诿{�C���t����g���&��?���?�WB���6�辰����V��U�C?���>���>=��>z�)���g����p:>�g�>��Q?�0�>I�O?�5{?�[?k<T>��8��(��iǙ�V�1���!>S@?ⵁ? ��?�#y?|��>b�>��)�� ྾_��\*��F󽽽����W=�$Z>���>0$�>A��>��=�(Ƚ����>��Q�=Jxb>,��>~��>���>ώw>d�<!�G?���>Jm��,��c6��N�����A��`u?/~�?�L+?��=���F�i��G��>}��?j�?�^*?�	T���=�ۼض�+q�cѷ>5��>M�>�j�=��C=7>��>���>>G��j�368��N���?��E?��=j+ҿ�Ł��9ʽ�-G���o<򕎾W�`�7�����}p9��]��/
s��ዾ�?�2n��X��K蹾!�þC���
Q	?�7@=f&?>5�!>�a��O-&��4�=QȽ�-��=�z��=g�L=�3��	�������'��[)�l�l��g˾�e}?8CI?ę+?�C?z>mR>T�1�U͖>�%���N?U�V>�WP�;c��5;�ͱ���3��^�ؾ6K׾B�c�����W>;�H��>�V3>hV�=ʈ<�,�=�Ir=C��=��k��Q=t[�=E��=�ì=��=V�>�7>b6w?=������4Q��V�s�:?\7�>�{�=3�ƾ�@?�>>�2��ԗ���b�q-?o��?U�?��?�ti��d�>����䎽Xu�=n���|<2>���=��2����>��J>���J��コ�34�?��@��??�ዿ��Ͽnb/>�7>d#>2�R�Љ1�?�\��b��~Z���!?�H;�J̾�6�>g�=,߾�ƾ��.=K�6>�nb=$g��V\���=��z���;=�l=�׉> �C>Xv�=,����=˜I=v��=0�O>�����7�a&,���3=d��=v�b>�&>���>�?O`0?]Yd?�5�>7n�Ͼ�B���D�> �=�A�>�ͅ=tB>���>��7?G�D?��K?���>Hʉ=d�>��>�,�p�m�
o徊ͧ��֬<薈?�͆?(׸>��Q<�A�N���f>�I?Žv?P1?yj?��>�����gQ �*��Ў��#9;�*=�e�J:l���7��-����H�=�	�>[��>���>�%p>re)>�F>�>�>��=mK�=D�	�HKr:B�˼�2=u�����<� Q�E���E>&<��G�����x!�J����M�e������=A��>��>K��>7�=�k����/>�����L��ڿ=$t��B@B��d�z^~���.� �6���B>x�X>;P�����0�?i\Z>5�?>�Y�?!�t?F� >tI��վe���e�1T�h1�=�_>��=��_;��l`���M�PIҾ)��>i�>{p�>�en>�+�{z?���{=��҂5���>��e�#����7qq�o����ߟ�z�h�]N��еD?��z>�=�1~?X�I?*��?{g�>锽��ؾ��/>PW����=eb��m�ꢔ�NK?��&?J�>���NfD�Z~Ӿam$�S��>��m���A��ܒ��2�_���,���VCb>�e���j߾ty<��˃�����J���o��l�>�Bd?]�?�ٽ]"���q]���˾��;d�>�J?%��>���>�C�>dG��h
�{�7�O+=�2}?!�?�O�?��>D��='��<�>�+	?���?ɸ�?��s?}x?�={�>ڢ�;h� >Y���0L�=V�>׋�=b*�="s?�
?��
?gj����	�������^����<�Ρ=���>�l�>��r>��=d�g=Xv�=l-\>ڞ>��>��d>l�>IP�>s륾	a��&?���=cO�>�2?�L�>{�W=+�����<�H���>��]*��ᵽ�߽'C�<�=���BN=��Ӽz��>Y�ǿ#Q�?5�T>�W��?�!��#�/��vS>XT>{Rݽ�S�>(�E>��}>�\�>T��>�>��>`�(>�MӾVX>A��VX!��,C���R��ѾWZz>䲜�c�%���������1I�fz���g�ij��,��;=�}-�<�G�?c���k���)�����b�?oR�>k6?�ь�*(���>���>ƴ�>�L��ꑕ��ƍ�Oiᾈ�?���?_��=��>1�#?�U>Jn>�F̽�y�FR��h$�5��+�v��3������zh��f�:[p?��?~�s?��'>[h�> �6?��@�8�v�$?b�����8�{\�=��>[�d����0���`���30��#>��? ��?��@?x�����=�q��ДG?��.?js?�"<?m��>֪�>�	R?'��>�he?��M?�?��7?݇2?�>i��w���V�|b�k$ӽ �=��ս�k=GS�����=�� <���<K'=�ʽ=?Jb��:�&���$=��<	J=]��=�g>,��>�1I?L8�>h8>�^?~c��_�^�_i���?�O����ƾ8���y7վIc	��>�V�?�r�?�7t?��=��������>޳>��<��>B�>R>�=M�����=��F>.gH>3mg;�����ѽ���8�a�i�����=z��>�E|>����l�)>pĢ�s�|�!xe>8�T�xa��CpS���G��2�$<v�	��>/�K?�B?P%�=�<�_w���e��.)?��<?�3M?� ?�؎=b*ھ�9�'�J��W��w�>���<;������� ���z:�����s>S����֠���a>�����ݾ�n�'J��_羺�L=��*X=T'�־��~�hi�=7�	>����� ���� ����)J??l=�v���oU�Ab���>���>��>�9�
v��_@��`��]��=d��>P;>������!�G�y5��ć>�E?��^?9W�?�����r���B�4���@ݡ�@����?Ϋ>=C?�]B>�H�=vo������d��G�	�>���>����H�𞾃���$���>Hh?
!>M�?��R?4 ?��`?�*?�O?H�>����?5��D�&?�Ã?Gw=\�׽�V��L8���E����>�)?6�>�e��>��?g?%'?��Q?��?�#>� �0�@�!^�>�b�>=�W�O��}a>uRK?(��>�}X?ʂ�?Qq=>�z5����楽���=��!>��2?��"?1�?��>��>�¾��=���>�e?}�}?��p?�>:>�?# >x��>���=j�>r8�>��?:bN?h�c?��8?#��>�Z�<2.w����C�h�nĽQ��n`$=yB�=�����I�b���7=�B<9��c�P�1&���.�;�f�<,�X;@t�>��s>�����0>�žlQ��C�@>a���J8�������W:��0�=^�>��?��>�M#�a��=���>�:�>���P(?!�? ?��%;H�b�P۾��K�9(�>#B?��=t�l��x��#�u�[h=_�m?��^?��W�r.���l?�~o?�L�X�3�U	��wH`�Y�zMI?�?O� <S^�>Z��?�g?�_?����uN��R����k��m����=��?�$"�aj�� �>��B?�Z�>ֲ�=�@>d���b�c�D��'%?���?�ê?���?
(>�dQ���ֿ��־'�|�}�m?�(�>���RP	?!�=�bɾ�����̩�Yi�j����	���Ό��멾�o.��)���;��`>p"�>^_N?�6Z?�p4?�h�eKs��`��3��P��K�P.�|QK�"kM��I�I{����0�9���ܗ�[K>Թ���AH�O�?�@>?�Xx�և�>V�e�������q�E>��Ǿ�7��@�=�����M��J6�GX�G
 �w�:���?���>���>P(Y?�"d�'_]�򆯾��4�C��&��>q�&>��w>�M+?2�~�pE���(�R��:�ܱ|=�7v>�xc?T�K?|�n?�o�+1�����K�!�(�/��c����B>�j>?��>��W�g��1:&�nY>�=�r�p��w��H�	��~=��2?�(�>,��>�O�??�{	�ok��lx�<�1�Ē�<.1�>� i?,A�>�>�н1� �G��>��l?w��>�>#����Z!���{�¨ʽ|%�>%�>���>��o>��,��#\��j��K����9�5v�=6�h?�����`�k�>�R?݈:طG<>}�>��v��!���@�'�A�>�|?���=��;>�ž%���{�07����=?<|,?r�
���(��b>��V?b�>�5>�z?�C�>ܼ1��K>F,?��o?�i?��V?7�>�Sp����]mؽ83�!6�>��j>!�|>B��<��=@��:b��I��.B}�||3> KH�ӽ�i뽅S!���f=s�?<��>�dۿDK���پ��r$�?
��舾bc���a��Ϩ�jV�����!`x�ٍ��&��V��6c�����ޱl���?y>�?���� 6��B���o�������h��>#mq��~�P⫾׻����˅� ���W[!�^�O��&i�D�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�A?%�(�`��(V=��>��	?��?>51��B���[�>�;�?��?ǦM=R�W��	�!ze?�e<��F�h�ܻM��=�%�=��=Z��ܕJ>4G�>ۋ�]4A�Iܽ	�4>��>H"���Iu^��޾<6�]>��ս�U��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=u6�򉤻{���&V�}��=[��>c�>,������O��I��U��=����ƿ�$�[|�_n=B
ݺ\�[��~�A����
U��$���lo�:��``h={��=��Q>�q�>�1W>�4Z>SfW?C�k?�M�>@�>%P�E���,ξ�A�kL������������裾^S�s�߾�	���������ɾP/�G=��U�ٲ���;0�+�[�ݣF��+<?ŘN>����@}0���=�ľ���m�8FW��i�;IS5��e�@�?�Hg?g˄��Bc����+,ϻ����==?����Ǿz����\>Ft=�o�=^�>F��=�Iվ��1���T�s0?�?~��L���#'>�O�=b�(?aZ?��m<�ԫ>�v&?�9"��ҽj<_>��7>>~?�>E>aگ��hὫ�?��S?�,��h֞����>���;{���C=d�>��5�0M�3�Z>5o<�� R��@����m�<],W?���>4�)��Hq����k==ϵx?�?�6�>:}k?�B?W��<]��(�S�2��3w=��W?%#i?6�>�뀽�о������5?8�e?��N>\vh����m�.��M�+?U�n?�`?i����m}�)������e6?f�v?�l^��i��`��ezV��:�>��>���>��9��M�>�v>?�T#�~L�������R4����?ȕ@ԑ�?:==<��FD�=�4?��>��O��@ƾ�-��;[��Ep=J�>�o��Uv����Յ,���8?i��?}�>����7��З�=�ە��Y�?��?e�����f<Q���l��s��!��<4��=�/�VC"����7�7�d�ƾ��
�+������C��>|Y@�L�d-�>H8�B6�6QϿ���B]оTHq���?|��>H�Ƚ�����j�<Ou�!�G�/�H�����R��>zWڽ������hJ���=��\�=��?W��	�>��H��z��;8����K>�T]>E>��1������؟?|���
ƿ�9���3�f)_?�G?�1�?�ee?���<��0>8�2>;�+��_z?�x?��b?�t2;�[q�O{��$�j?�_��wU`��4�uHE��U>�"3?�B�>U�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?us+?�i�8���[����*���+��<A?�2>���G�!�C0=�VҒ�¼
?T~0?{�e.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?/�>��?��=!6�>l+�='���@-,�$#>0J�=D�>���?��M?�a�>���=��8��/��BF��AR��$���C���>#�a?�|L?�b>:���%2��� ���ͽ��1�͸輪h@�!0-�;t߽Z5>��=>��>3�D�5Ӿ��?��fؿl�����#���3?Y�>��?�M�	^w�#kE���]?�M�>�-��2���狿�� ����?��?	?�׾��Ҽ�s>+�>s'�>�}׽����p���r;>�?B?�`�l����o����>��?��@7��?5Qi��g�>���cR��k����FǾ�s/��g�<��?_Iܾt8>��>�q�ƭ�����mw���>&ǯ?��?,��>��g?�Jl��:6�P��=K��>A�h?���>kZ
=Xt����>�r?h]�陉�|0�Mk?6�@�v@nMg?%���ެ�����hс�FН��t�=���='e>�$��:�=���<��N��A����=�G�>�u>&�>��C>��'>6�#>���y���Z���6��~�A�y#�M��D��b�
���������e��b�;с�a�,�+x&�9��K@���<�,�=<�T?�#Q?�,n?\�?��b�b|>շ���=��"�Z	�=}��>	/2?MJM?C�*?a^�=_���c��<������Zщ�n0�>�L>��>h�>���>��<��G>$l<>�2�>.�=��=9�K���=;P>Ǩ>��>fN�>fD<>�>Rϴ��1��f�h�[
w�
̽�?倝��J��1��=9��C���qj�=^b.?�|>����>пb����2H?�����)� �+�/�>��0?�cW?��>�����T��9>����j��`>�* ��~l�{�)�>&Q>&l?��f>	u>�3�e8���P��z���j|>�36?)趾�C9���u�s�H��aݾ)JM>3ž>	�C�&k�8������ui��{=�x:?��?�;���ⰾɮu��B���PR>�9\>�Y=[j�=�WM>�kc�s�ƽ�H��i.=���=¯^>�%?��+>RA�=�l�>)�����N�Q��>��B>��,>�??<;%?��
����:�����,�Ww>�t�>�j�>�>X\J�b�=j�>N�a>�r��[���B�/?��gW>ؾ~��^��(t���v=;-�����=�r�=�r ���<�(�(=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ^[�>���&U�����G�u� #=���>	2H?�h��YhO��!>��k
?�?�h�����ȿ�zv�}��>��?���?.�m�>@���@� t�>��?z]Y?�i>�H۾�vZ�\��>H�@?��Q?�5�>.�ؒ'�V�?~ض?F��?hI>���?�s?�k�>1x��Z/��6������9p=��[;�d�>�W>b���ugF��ד��h��t�j������a>��$=8�>aE�_4���9�=��	I��!�f�=��>�,q>�I>W�>y� ? b�>��>�x=�n��Kှ�����U?�|�?��6���h�T�M�-0%>�[�O��>��??�>㍍��7�>�/d?+��?�i?��>��1����^��,B���iS;��>��>���>+��=�3�>o+ӾR�@��t>�S>�3���y���y�W5�=ѵ>x�?05�>L��<7�!?�{!?�c>!�>*�F�-���X{E�C��>p/�>�D?��~?�C?�ܹ���1�V��I ��k�Z�("H>�5w?e?�x�>jo���ҝ���5���;��o��X��?��h?@�ѽ�\?�3�?�$??;DB?�i>M���־�벽
�z>�!?��A�7H&�F>�f�?�9?���>Df���ӽ��мX��A���L?KE\?�T&?"��a�^cþ���<�%��HX���;_�<�Z�>I>����=��>M�=JFm��5�`�l<�J�=ٖ�>_s�=qH6�BN��� )?f㪼rՂ��x�=��p�w�C�[bt>��G>[)Ǿ�a[?�
B�N�|�>嬿R��laU�d�?|=�?��?���q�e�T�:?�O�?�H?�.�>�v����оUy�{O���i�H��.B�=���>�����j�UQ��
���C��x���I����>yQ�>޹&?��>�_=��>f��XF�/+��u��f�+񾏯K�o^;���!�DAɾG�1�SЫ=�_��P�g�Í>2\F�ܯ�>�[?eG�>��>���>���;oȌ>�3t>�ċ>���>:�O>6��=U��=k�����ҽ�pR?����l�'�8a��@���A?1d?u��>�e��T��go�Θ?c�?�_�?NCv>Kh�Y!+�E ?���>/��?;@7=Q\%��s�<���V�������WE�>��ս�9��L�kxe��q
?9?1׍���̾��ؽH�Ծ��=Mz�?�|?2�%��f�B'R���^���Z�x���5��V��}4 �e�p�LZ��5���ᅍ�� ��QA>��?T�z?1�����yp���oY�(#2��>?f�>��n>Yʇ>�R>����C�%�� b�8�'�i�{�w��>k�y?�s�>RI@?<�?D'?��B?��>	_�>W����=�>�1<�>m	?I�:?^??�|3?�$&?��?1>�)O���g�����<?�?ĉ9?c��>��>����(ܽLߢ���E<�e��.��"�t=�q�<V����"���=Ա�=�X?x����8�l���^k>t�7?��>|��>y��-��I�<��>&�
?9G�> ��}r��b�KV�>k��?���J�=r�)>���=����iӺRZ�=������=�7��ay;�&g<��=E��=�ot�����-?�:���;cq�<p��>S�>��t>Kjv>1N�z��	a&���="�=��=��=�C ��=��s���KT��]>⅙?L��?c�=
�>���=$ފ���,�+�Ir�E.>�4 ?���>I\P?m�?.*?��3?���=���N��������о:s?n�+?��>�����ɾk꨿��3�?�?�?�ta��E�*S)���¾�Խuw>Kk/�~�����(�C�MHW�i�����g��?|��?;C���6���ֱ��}��g�C?���>�G�>>��>��)���g�����9>;��>�R?�#�>l�O?�<{?��[?.hT>J�8�i1���ә�B3���!>@@?��?��?�y?�t�>�>$�)��ྫྷT��_��������MW=�	Z>?��>�(�>x�>���=�ȽmZ��A�>��`�=��b>G��>���>��>�w>K�<O�G?���>^��?���뤾Ń�g=���u?���?��+?�S="�� �E�ZG��QJ�>7o�?���?34*?��S���=��ּⶾ��q��$�>۹>�1�>|ȓ=�uF=�b>��>Ҡ�>�(�a�q8��QM�n�?oF?{��='�ſ�q�h�m�����y\<�����a�����[�6g�=��ct�=���i�\��������#㵾�ٜ��{��h�>Z��=͢�=H��=6h�<��ż�U�<CG=W��<9�	=>�t�a-_<�F9�5z��т��p�8��O<<�A=��⻐̾#�w?g$J?cn)?r�@?B�{>">�[�^��>(ʄ��?�w`>�j?�����+�9�xM��Mѐ��,پ��پ�^��Ƣ����=�SD��>�2>;c�=<(<���=��?=C�y=,�仗��<��=��=�=,��=��>m[>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>X7>��>.�R��u1��+\��6b�O`Z���!?t&;��P̾�D�>1J�=�߾�sƾw�.=k�6>$ic=AW��M\�G�=oq{���;=N�l=?��>��C>��=1�����=d\I=j��=˓O>纗�8�JL+���3=�=4�b>&>y��>��?�a0?0Vd?l8�>�n��Ͼ�6��=J�>5�=I�>�=�xB>��>��7?�D?��K?���>楉=��>C�>_�,���m�t�ķ�`��<���?�͆?�Ѹ>�$R<J�A� ��i>�YDŽ8p?<S1?�i?��>�T�ɡ�V&�q�.�#��75÷�+=�cr�QAU�#"���d����.
�=�o�>���>k�>�Qy>�9>��N>s�>~�>���<us�=���L��<�������=z����<J�ż�ό�^i&���+��,��o�;	ӆ;(x]<���;���=]��>�E>��>��=��ZF/>_���M�L����=�J���+B��3d��H~��/��[6�O�B>t5X>Hj��[5����?��Y>�d?>Ѓ�?6=u?�>=(���վ�Q��Ne��ZS�r��=<�>R
=��|;�r[`�s�M�MtҾ��>ʵ�>��>B�o>m1,��?��*�=��⾤&6��s�>�����'��S�ښq�3?��П�{<i��˺i�D?����m�=��}?ѨI?���?��>�蒽�ؾ��/>o-���	=я�-�m�ָ���i?�y&?�8�>�:�D��~�����>{h����j�8�u8���ƥ�^�)=�����p<��6z�t���C/X��ϛ�=��>�,r?���?�N5�JJ����B�p����#>	�>>�D?e��>X~	?Bn?�d?��� ��&� Q3>*�j?[!�?���?R�|�*��=>Խ?;�>3�	?(ɖ?��?�1t?�4�E��>�w;̆">4���S��=��>�~�=3��=��
?XU	?
�?�7�������"���b�o��<��=��>:,�>:�k>ߣ�=,�j=2��=3LY>�7�>�>�ki>DA�>B��>B������&?�Q�=��>o2?��>��Y=�|��}b�<�I�E�>��+��r���ཅ$�<o�[��,R=�	м�>�hǿ��?�4T>!S���?����X0�8�R>��T>��޽�a�>�E>��|>ڮ>P�>�q>:Q�>�'>BV߾�*">�꾕]�?�<�PqV�XJƾ��P>���g1d����2��Ih��o�����"3m�*ц�p=�~�=��u?e���gk�ɽ2��}�0��>F4�>^d?j܆�����{=���>�Z>{��6��̒��"��k:�?�^�?��@>_B�>qR?��?D�� �+�ڳ`��!y���;�sc��c��o��&n��Z����뽏�Z?�?�L?�X=%ׁ>t?/1 ��G|�K\�>�D&���9�!�=2>�>�e��$P�;Ͼ&¾3A;��5e>�8i?�w�?�?�[j��"�pɜ�r >?ӷ?P?��?|�?vIh>JT?8�N=�"?�?��?ͩ?1&�>Mu>�3>�q�� �:X��3=���+���¼+yp� ������=�{<�5��!�D��h����~@Ž�޽x��k	���=u��<�>p9[>U�@?���>��>b�K?B�}V�K˾3�?L���᯾:ľl�����zؙ=�W?�y�?��?.u>� ��$8{��$>2B�>ݎ=��K>�_�>�BE<0���k�=��?>��>{��=��&���iC��Wf�k$=���=�&�>b�}>̆����'>����z�zwe>۾Q�
ɺ�a�T�P�G�S�1�7�v���>�oK?1�?gו=��龃����pg�;p(?<?�TL?�?�6�=�`ܾPD:�l�J��p��#�>��<XQ	�����W���;���к��r>���뚾[�[>����x���,h��:M�q�뾏!=s����)=<Q���ƾ�du� �=l�=�;�g"�����*��zjF?�8�=�����,I�S&��I>�Q�>�>�Җ�z�Z�֦5��̣����=��>��+>��"�eW�<LA�7�����>t<A?sH?e�?�����7�gL�پW;����Q�7	?��>4�>�G>*�x=n5�����Ycd��L����>}�>?��/[J�xO����)^"�Q�S>*
?�m�=U?a�R?)�?ɕ`?YL'?��?"��>��ý
C��z�*?�0�?�^��k�+v��b7�*zL����>�5'?H�d�lu�>?*.?�*?�$&?FR?k`?���=��֙F��Ӂ>+��>�yS�*8��H��>�dM?�S�> @?zR�?XdI>X3�Z�ʾ��V<��>�C�>�%O?&I/?�M
?�>]��>���Ie>��=(mv?vJ�?���?� �>���>��E<�x�>�p����>�?��?5Y#?cqK?�H? ��>۝�=i�"�c�P��K����=]~&>f�=:��=�N0����r�J�0�=��l=����K��Y����/&���=9�=wb�>�t>)��F�0>��ľQD����@>���u"���؊���:�eݷ=���>?Pŕ>k�"�6��=@��>�-�>1�� (?x�?N&?��*;��b�-�ھ�K����>Y�A?s��=��l�Ճ��4�u�TXh=$�m?ݖ^?ZMW�} ��3�d?e�]?�z�*���������fv�ʮA?���>�J3��_�>��?� T?~�>��4��Z�?��ѱj��k�����=���>���3�]���> �5?��>.s>'�>����]�����m/?�?��?��?e�~>��_�пO�
�����XH?N\�>�t���?%�~�2j⾆���1x��T��QB���?��(�ľ씥�c�;�bgr���J�L��=�d?�[z?��x?!�v?8,�&�S�<a�)H��j3U�$��hd#�4�V���+�@�#Wi���9��������zν�~�A.<���?2�%?^+�&�>�j��»�B����H>�D��c���p1=AW�'G���E�ꊾ��F�T����+?��>K��>=�6?��i�L`8���=�~�+��9��i�>��>�$�>���>�qM;@c�!��U��`�S�ڕ���>�a?ޙ=?Ao?<$�ؿ8��6�����A�J��{��C->>q�/>�8~>��n����r
(��?�Tft�:�P���Q����=e�0?؅>�e�>���?��?���v�ξz�����(�i�<Ɓ�>�3e?FO�>!V�>kL۽&�+����>.�r?�L>pߞ>�<;σ5��%t���|��^?��?x�?�E�>J���.6�ʂ������_UF���y<K�y?
��}��@�O>��`?�r�=�)� ԉ>QR>D�4�8?�xy��s�>��?b9>�)�>̮f��8۾q�`�=ݾx�(?FA?9꒾(�*����>k�#?�8�>RB�>���?D�>J��iv�=�?�^?��I?'�@?1��>c>+=�V���Ƚ>�'��l2=@��>��W>��_=w��=���XQZ�����E=p�=e&�9/��:0<v2���|s<l��<q*3>)�ڿ�K� �ؾ�S����	��V��:��ƈ��~�̝��������x���;�+��V�,
b��d��_@k����?���?[���}����䙿8��q ����>�t��k��9������*��|��3׭��n#��1Q�/k�hf�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���z¤<���?0�@�|A?h�(� ��IV=���>Ł	?8�?>� 1��J�&���E�>;�??��?�>M=��W��)
�'ne?�R<��F�5ܻ�/�=HU�=4�=j��_�J>D�>gw��XA�ܽ͜;�4>g�>,W"�ݗ��^��H�<�]>��ս`���5Մ?,{\��f���/��T��U>��T?�*�>U:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=s6����{���&V�|��=Z��>b�>,������O��I��V��=���(J¿�� ��"�D�<��a� V�,�ὦL̽����]��b�A�8���	u�<���=��t>���>��a>�q>�X?~Nn?���>��}>ɛ�!�v�����l%�8A���-.�^K��l�F�<Ǻ��j�<���4�e�)��4/��˾��<�n�=9R�w���� �,�b��F���.?��#>0�ʾ��M��2;<�~ʾ�֪��W��Z����T̾�1��n����?�A?܅��V�����O��v���W?ʼ�����⬾v�=���]=� �>+_�=Ҥ�z3�&�S��/?�L"?�3¾ڕ��=3>�C����<��%?l�?X![<�ǚ>�#"?�%��nѽP�{>m�a>Jϫ>��>y��=�鯾;�꽫�$?�S]?D%ͽ�5��݃�>�淾�ၾVb}<���=�B��JV�u�1>)��<�2=j!!�93=�&W?㘍>��)����Z�����ˈ==	�x?��?�-�>�yk?��B?w�<^c����S��^w=��W?�)i?��>�p��9	оr~���5?T�e?��N>�_h������.��U��$?��n? Z?�|��(u}�g�����#k6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>��������>�U��eH�?���?sô���r<�s���f���	���;=���=9��c�v�G+�c�;��o;~c�蓑�9켤�>��@��^��>�|��Q�п����,˾��Q��!?ߢ>tF ����1�j�+�u��:O�[�H�u�k��N�>\�>5���������{�rr;��T��k�>(!���>��S�@!��E����X5<��>���>���>�5��D齾�ę?:a���>ο�����żX?g�?Hn�?�p?&M9<=�v���{�/��.G?S�s?pZ?�b%��<]�!�7�&�j?�_��zU`��4�yHE��U>�"3?�B�>F�-�9�|=�>���>�f>�#/�z�Ŀ�ٶ�H���T��?��?�o���>k��?xs+?�i�8���[����*�H�+��<A?�2>����A�!�@0=�8Ғ���
?S~0?	{�h.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?|ڹ>�D�?��=���>��=)߹�[����L0>���=/RI��?�P?���>���=z�8��^/�=�F�D�R��.	���A����>��a?�I?��]>永��]������".A�V���J�3��� ��2̽��.>hqD>r3>�>A�#�׾��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*��Կ�졿3mܾ>\��B|=j.�=�Hf>^�0=�U�=�@�o�}���=*��>QB�>��%>�4�>��> ��>S�&>^��&�!�?���y���ߪF�V��K$�'\�8�ھ=o��ȳ���o��8��s���H��-��̽]�&�I���|��={bU?�$R?�p?�d ?x�z���>"V��R��<�#�u�=�N�>�h2?�2L?MI*?�ʐ="���t9e�(k���v��}i����>HaH>f��>�t�>�~�>�;��H>Js@>:u�>xM>R�%=�P���
=)�O>�Ī>K�>��>~D<>�>.ϴ��1��M�h�]w�E̽5�?���,�J��1��G8�����g�= b.?�z>����>пV���u2H?���)�/�+��>G�0?cW?�>����T��9>����j�a>, �~l�X�)��%Q>�k?�g>�au>��3���7�[�P�&�� �y>>�6?����F�9���u�/�G�v�ݾ<�K>�F�>��Z�b��:�������h�+z=Ʌ:?'#?Bг�U���y>w��ѝ�b+P>��X>�=G�=�xM>�%]��Ƚ8F�m�/=���=��[>]?P�+>���=|�>�R��ïP��T�>��B>��+>B�??q%?�`�N��胃���-���v>��>0݀>�>u:J�T��=�u�>°a>?R����_�M�?��W>7���y_��t�)�x=������=���=E\ ���<��$=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾRh�>sx��Z�������u�e�#=N��>�8H?�V��|�O�]>��v
?�?�^�ᩤ���ȿ5|v����>X�?���?f�m��A���@����>9��?�gY?toi>�g۾9`Z����>һ@?�R?�>�9���'���?�޶?կ�?�D_>T;�?~�h?t��>�fֽ/L/�����#�����=^'O=���>�b>�VѾ2]L��͖��e��n`l�0��0�>%I;=��>�������R�=Qǜ��Е�[�k�]��>F0t>�">sV�>p?K�>�Θ>�|=g<��Vm� ����I?�ޔ?�E*�zSl���7<5S5�����b��>��O?����9ᾑZ�>f1_?1�?,�k?`�>��ݾUÑ����������Q�<Ά>)O�>�0?<$�	��>M־�u׽��>�Z,>����
�YJ����=l��>iK?��?)>�3?��8?ǀ�=�;4>qEz�Rd���J]������?�8W?��?u7?z*�lph����EN���Vu�[���#�?��	?b��>h��ݎ���=:��� >	�K?�ք?���X�>{Ȁ?*�=?���>ãi>�L����l���R>��!?
/���A��Q&�׻��?��?�4�>(���6׽��м��-��U?�\?.&?f|�,�`���¾8��<ư*�oyG��V<�K�5�>o�>�E��b��=�>k�=��m�x�6�J�h<g�=�Ԓ>�p�=�7�;��0=,?��G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>#�l���K���ڙ���F��_�Ž0}2� ��>8��>`%?���>r�5>��>�䯾��-����d ��,_�u��7�5���*��^��慨(&a�rc���z����f��>�Э���>i!?�0J>��>�Y�>b.=��>��T>ĉm>k��>��M>��H>R��=�C0=a2�27R?����;�'���边*���XB?�d?�S�>l�h��ҟ�0`?{�?j�?W1v>~Th�?+�p?�*�> ���Z
?�g:=����</H��J�������v�딎>�׽:�`M��{f��]
?�/?ؚ���i̾�>׽u��m�,=/��?��"?��O�7�5�<��UZK��ń���]>ls=����K�HQp�*�������E���"�k�=È4?�ď?��FF�aK$���n��R��>�BL?���>�`2?��1>�61�#�A�)�_�A&��Y��ٟ4>��?���>EnO??�M?�w�?�C?���=���>	���7`?��_��w>�a�>n*�> Z)?��c?EO??�T?���>���C��/6��\hL?Ğ&?���>R�)?r�>?��ҽ�D
��|x�aiM>r�ƾ����te�=?Y�����Iʡ���>ר=��?U��8����l�x>z";?�|�>�e�>  ��I��'��<p��>G�
?*��>_v���~p�5C
�'��>�o�?U��Ю=S%>�+�=I���o��;��=J�j�r?�=� ��BBE�:�{<҈�=�U�=�t��S��\V/�)��:���<�t�>)�?Г�>�C�>�@��$� �e��$f�=`Y>LS>m>�Eپ�}���$��w�g��]y>�w�?�z�?k�f=1�=Ӗ�=�|��{U�����M������<�?2J#?,XT?c��?{�=?Nj#?��>+�hM���^�����î?�!,??��>����ʾi��3�C�?>\?�<a����|;)��¾��Խ�>T[/�6/~�����D�`��#�����՛�?6��?%A���6�z�2���]��6�C?� �>sZ�>�>��)��g�"$��1;>i��>i
R?�$�>B�O?h;{?Ҧ[?�dT>$�8�O1���ҙ�s3�P�!>]@?M��?<�?#y?�s�>^�>��)�ྻU��y����M�����V=�Z>D��>�'�>��>���=�ȽyV����>��i�=�b>D��>M��>	�>=�w>�?�<[�G?x��>����Y��,��g��n:?�R
u?v��?eJ+?0=�/��E������K�>痨?%�?��)?ET���=Tܼ�����im�v��>>�>��>��=��A=�m>ć�>��>K�����V8�G`K���?�KF?�`�=�AĿ��m��.^��5��l*`<����f�mý��l�ʢ=���!�"��ʡ��a�t���z��^���AY��h���UW ?lf�=h�>���=�
=�&�b<�{=^<t\={��)=i<_�1���;􁇽�\�;6c�;��f=���T�˾�}?�;I?�+?	�C?��y>�:>�3���>����.??@V>̑P�������;����� ����ؾ'y׾S�c�[ɟ��J>*hI���>"93>�B�=�b�<^�=�$s=�ʎ=��Q��=�(�=�N�=�j�=���=��>�T>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>WkQ>�P>|�R�H�"��\j�����a!~�$q'?��>���˾p�r>)�>�6�p�ʾ�3=��>�Ґ<ϟ6�%�]�9"�=��j�]�=�A"=��}>�HH>÷Z=������=�A@��$�=��m>�*V<��< M���=���=`^>���=,��>3�?m~0?}ld?.7�>-�m���ξ�"���_�>���=yK�>�=�LB>���> 8?M�D?J�K? ��>b��='�>Cͦ>�,��m�_�_���#��<7��?9Æ?�ո>0�R<�B�����`>�z�Žji?�?1?qL??۞>Z|�ؑ�LU(���R��7P�_1=�\�=V�a<�:
�G�v�Ȥ�5됾%�=��>Pَ>Gc�>B�>T.}>�,>�>͝>��=���=���;����sx<�أ<�f�� ә=ˊȽ��N��er�zLk�BT�=�Ż���9Ů��
���^��=!��>"<>��>���=����C/>�����L����=�G��@,B��4d��I~�A/��V6�.�B>�:X>�}��74����?��Y>�l?>���?9Au?��> ���վ�Q��!De�VS�]˸=��>��<��z;��Z`�r�M��|Ҿ���>�̓>��>��s>:-�'�A��H=����G0�i��>;ʆ�{?��T���rs�pW����_i�'�k�,E?�چ��W�=-�{?�xJ?a��?ï�>8��#Uľ��>�	��j�<�h�~a���O��?WT)?�G�>{��O	I�3G̾h����>-I���O�o���<�0�.$��淾L��>������о�3�kd������.�B�i_r��غ>b�O?��?#Sb��L���PO�,������`?�g?��>�L?	L?������p��F�=i�n?���?g@�?>U��=;�����>��>h��?{�?�}{?�̽no�>5���n8>�51�4�5>gk>��>f>�?�P?��>=v���X�'t�������j>���L�<$�p>mO>�Z>���=FX�=��=�U>��>p��>i*>���>�K�>-�������w7?��>ݏ�>�u'?j�E>z3;=�f�|�`=��߽y Z��,�k�����	�]���TCs��ֱ�YO��2�?�v���*�?��>7�}�$?3��#��=d�>��>�Z= �?�7�<�vX>��X>tX�>�7�=c3�>��Q>V6Ӿ
�>���� ��B�~�Q��Ѿ#;z>������$�+���`��zvI�2���(_��i�`���=�ı�<�W�?IV ���j���)��c ���?�>Ձ6?B>��o̅���>���>��>���������i��q���O�?B��?�;c>��>C�W?�?��1�A3��uZ�%�u�f(A�!e�V�`��፿�����
�8��-�_?�x?"yA?�Q�<0:z>I��?��%�Cӏ��)�>�/�';��@<=`+�>"*����`�r�Ӿ��þ8��HF>��o?:%�?�Y? TV��l��b�=I(=?�&?��r?q�A?+�H?��NR?�J>x��>ai�>~??�.?�!�>�+>��@>��M=
w�<NF����� ,:��-/�q��6l���㣼�S̽�戽Ov�=��=?�=κ鼎: =G���c׈8z�<�_�=��C>�l�>97^?���>ΐ�>ѫ7?]f#��]6��׭�Z�/?~=<&��=:������>�x�>~m?� �?��Y?�/\>��D�
G�#�0>��>�w*>l`>�Z�>�J�O�J��K=kL>�>�֛=�O�Ec���^
�����*{=��>b3�>=�>Z�Z�&>�����~�nEa>C�R�w,����R�.H���0��t�?��>��L? ?x�=A��ss����e���'?��=?L|O? �?��=�\ؾ�8�ɊJ�!�$�P��>���<��	�墿%��Kz9�h/H<�py>�����ޠ�Wb>н�	t޾�n�J���羺GM=���YV=����վ�4�S��=1$
>������ �"���֪�S1J?��j=�w���bU�1p��l�>ƿ�>�߮>��:�I�v��@������5�=���>��:>�a��I�~G�8��6�> JE?�S_?�h�?���|
s���B����7a���Qȼ��?o�>h?B>��=q�����]�d�G��>I��>-��V�G�!<��-����$�I��>�:?X�>��?��R?��
?]�`?*?�@?�"�>��������C&?�?�ل=��Խ��T�t�8�F�!��>�)?��B����>�?ɽ?��&?��Q?��?��>� �LF@�2��>\�>��W��a���`>��J?��>z;Y?�ԃ?+�=>΅5��좾n֩�"a�=�>[�2?_6#?S�?T��>���>
��G�=�ʡ>��g?wڃ?VWj?���="w�>��(>5?���=��>=��>%�?^?F?s�p?�@?B��>�}�<V���*���"Mz��v8=���=>��<� d=-��G���`?�-�{��SU=ڟ<���\&.�_�I��;���$;_�>��s>y���0>��ľ�P��W�@>1ӣ��O��E֊�v�:��߷=��>+�?���>aP#�互=��>	G�>����5(?�?�?��";��b��ھ��K���>zB?|��=:�l�������u�o�g= �m?ڋ^?ЕW�^#��_Lx?��>?��,��J�:~	�Dþ�F�N�?��>ù���z�>���?�B?�, ?�u�!{b�D����k��<�����=}��>�j�N9q����>�K?�M�>~�'=>-�` ��e�����>2?�׳?���?p��?���=�Y�������{�3����_?'�?�M���"?Q��=����B��J�,��,������jQ�f����g��/{
�P^�k�ޏ�<��5?7�w?��m?z\C?���`?��H�G6K��9�o��GU��2H,���F���H� ��R�

��ߎ��7v�	d��YQ8��8�?4�2?�AU��:?iH��|Ͼ<5���N�=�R˾��r���=�㽛��	�뼉�(�v�����۲;?.CU>}�M>�p;?�ԁ�w%/�k7L��_�;8�NLy>-�>_֣>S��>��=e���Q���������ɽ.7v>�xc?d�K?��n?o��*1�v����!�9�/��b����B>fh>���>��W�����9&�"Y>�X�r�����v��V�	���~=&�2?{(�>Ӳ�>�O�?�?�{	�k���jx��1��<-1�>E i?�@�>��>�н�� ��D�>9�d?и�>Vl�>Z"��m�,���~���;����>�w�>_&?���>#j^��Mb�mގ��Ӕ���9���=Ңq?1t���h��Ou>�B?O&��m�_��>e����$�5�پ0, ����=��?;>�R>ywƾ�y�]�x��ի��(?]#?�S��h'��6�>��?��>3�>L��?hש>�[��,�;V&?�*^?f�K?�cD?6N�>ah=Ebؽ��ؽ�M(��.�=h��>�m>�)=�Y�=���$sc���!�r�/=�B�=�^Q�]�ѽ��;�����<o1=/>iۿ�PK�\پ���?���1
�*�������3������ߛ��j��xx�9����'��V�Pc�����
�l��~�?�=�?�:�����ʤ��%��������˽>*Wq�Iʀ�a﫾B��3����i鬾�j!���O��i�\�e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >ZC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾w1�<��?7�-?��>Ŏr�1�ɿc���|¤<���?0�@ }A?��(����V=���>Ԑ	?��?>\S1��I�5����T�>[<�?���?�yM=��W���	�7�e?3�<��F���ݻ��=};�=;H=z��l�J>�U�>F���SA�,?ܽҷ4>�څ>�|"�]��,�^�l��<Ç]>��ս~;��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��=����*ο�=��i���.=�:�<'ꄼ�%� �?�~�?=�����3�1�2��Z�=�y�=�b>>]�>�4>��]>��a?8a?��>�>�[��E��뛾 �k�����Ծ��P�t���辪��J�]3����q�Ҿ!=���=7R�j���<� �c�b�O�F���.?�v$>m�ʾ��M���-<}pʾ_���}܄��ॽ�-̾�1�""n�g͟?��A?������V�P��4W�~���Y�W?�O�߻��ꬾ��=����D�=%�>�=���� 3��~S�/k0?+�?�<���L���*>����=�*?/�?³�<>�>Bs%?�+�S��/�\>+�5>,T�>�q�>�q>�>��ē۽b?G>U?ƕ���T��L:�>o���r�z�dI\=�&>�5��yܼ;�Y>NY�<�
����L�������<ڦh?w��>��K�����w˾�恾�C�����?�p?M�>N�?v
]?q]i���0���`��[�j�q>��^?�2�?J�>�꽲��� :>��43?�A0?��<8х��쎾Ԓ)����D�+?GjL?���>�h�=�k��Ҝ����/�� ?�Ww?!X�1O���)�p7j�7�>���>���>�7�ك�>�=B?�7%�,����4���07���?&^@�;�?��<�8�Y��=�W�><��>��M�nOž᣽����(z�=ʇ�>!�����k�r��5�/���9?Dă?
� ?Y�������=�ܕ�/Z�?��?+���T�g<B���l�'r��"V�<���=��iZ"�1���7���ƾE�
�5����ڿ����>�Y@#W轎&�>�I8�g6⿍TϿ����\о�Uq�Q�?R��>��Ƚ՜����j��Pu�ʴG���H�g���BN�>��>s�������E�{��q;��(����>	�f
�>[�S�'��ʛ��n5<��>���>$��>O#���潾�ę?�b���?ο�؝��X?(h�?�n�?�p?��9<��v���{��z��-G?��s?nZ?�e%�X=]��7���j?D��\Y`�b�4�%NE���T>3?�J�>B�-��t}=�L>u�>�>[*/�%�ĿSض�٤�����?��?�^����>�t�?lo+?�i�	1���5���*��{'�9A?Gf2>�o��ʧ!�0&=�����J�
?#�0?�x�k-�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�$�>h�?�b�= `�>Ni�=�-��_#>*�=��>�J�?ǨM?�I�>p]�=F�8��/�YF��FR��$���C���>��a?�L?�Pb>J"���2�9!��xͽf1��c�]W@�݉,�x�߽�'5>��=> >)�D�Ӿ�?}u�ؿ�r���-�$�1?(=�>��?s	�'�n��<黙�\?5ڂ>Q*��h���S��,g��^+�?��?Ql?��Ծ����r>e��>ك>��-ߖ�lB���V;>�GD?VU�ډ�ɦn����>���?��@(�?��h��C?��ھ�鈿l���h�zn���=�87?��ݾ��>g�?��=I0��������~���>a�?���?� ?`]^?��[���@�E��=,��>��W?�S?���=�پ֟U>�+'?S<��f�����h?��@�P
@mN?qә��
տݠ�m3��Ľ׾�@�=yA>�P>Jԟ�Ǳ�;�X�L�8=���=�=>J_m>��}>�^�>9T<>��,>p&>��|�s��꥓��^��-�H��_�W+�hs_�c%�Hh�N��ٛ�'�����~����wr�1iF�b�ٽ�B&�ۧ�=��A?<W?spw?�"?k�J�/ x>1ξ�;>J�*�д=�����C?m/M?ء-?%F�=@_m��l��_������H����>u8�=���>S��>�^�>�U�<m�c<��^>q��>#5>#��=s*�<�#J�@�>p.h>eG�>��>�G<>�>Aϴ�L2���h�q
w�\$̽s �?%���ϼJ��1��7�����~z�=<b.?x>���f?п����x1H?P����(�<�+�"�>��0?cW?d�>y��?�T��5>2���j�Rc>X$ ��wl�(�)�2'Q>l?Y�f>Ou>B�3��d8��P��|��dj|>�26?�鶾�C9���u��H�FbݾiIM>mž>|�C��k�Z����$vi���{=�w:?r�?�6��qⰾ��u��B��RR>�7\>X=Kp�=�WM>eoc��ƽ�H��i.=���=b�^>�.?!->Gf�=Cr�>�o��̀Q�y��><@>�`+>3@?��$?�.�*��1傾�-,�tax>�y�>Ā>O�>F�J�T֮=Ė�>[�c>�.�g���|��t>�8W>I����^��o�Z5y=M������=���=�{��"�<��Z(=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�k�>�r��Y��V��g�u�c#=���>�7H?�V���O��>�t
?�
?�b򾱪����ȿ�{v����>!�?��?/�m�B��&@����>֠�?�iY?�oi>�^۾5SZ����>&�@?	R?p�>l8��'���?�޶?﭅?�I>���?m�s?vk�>p3x��Z/��6�������t=�[;|e�>Y>�����gF��ד��h��q�j�b��h�a>&�$=��>E�e4��7�=���H��s�f�{��>P-q>��I>�V�>�� ?�b�>���>�w=�q���ှg����U?R��?�N?�֎�����݅9=/Ⱦ!Q
>qN-?�����Ҿ(�>Nz3?j��?^kb?�?��{���zn��R�Ͼ2Z>��h>f�?θ?��۽3�>j��\k��E�>'v�>m����/��`����T>���>O7?^i?�:c>Z�"?J!?��V>�k�>�F�m����DK���>8��>�?�{?�?�	ɾ��5�[���K��h�]�N^>|?�?y��>����^m����:�Fk�~Ya��u?�_e?���ĕ?��?��??2�>?��]>Н���ɾ����3�s>o�!?�%�u�A��<&�����j?�S?���>V���ս
�ռn��G^��L�?�!\?r?&?���*a�u�¾��<�'#��]��+�;�
G�x�>jD>qj��۴=U�>��=��l�ta6� ,a<�}�=|�>��=77�����P?,?G�n䃾�՘=�r�TzD�C�>+lL>S����^?�E=���{�]��Jy��eU����?��?�l�?>ഽq�h�> =?�?�
?�$�>@H��)޾���?w���x��s�*>���>�Em�h����ٗ��G����Ž󚤾#�>��?��?�a�>�j�>ì�>�� ���'hD�W�'�^�b��O��?�o>���#�S\W���T��V&�� ��Ґ��Џx>�wF�V�F>�$?,vW>1��>�<?���Z��><w=�K�<� �>`�\>z�=y�0>4Q>�Fɼ�KR?����$�'��������e3B?�qd?P1�>�i�<��������?���?Us�?!=v>h��,+�}n?�>�>H��Wq
?yT:=/9�G;�<V��y��3���.��>E׽� :��M�Anf�xj
?�/?�����̾�;׽�lB���ýN�o?�O.?��b���(�}��,{Q��2v���9��������5?Q��e��@��Fφ��������u>e�;?��?��f �ëS�����g���>�K�>~>')�>��V>g*>��2��́��r6�~c����?�Ȅ?�j>m?�.?)=t?.�U?OH>���>4'��= ?��r��~�<ˊB>d�<?�;0?��`?�>?�&?i�P>�:Ӿ��������S?0"?�D�>�?���>`$=6��<3�,10�AC���>�ܸ;_%��8���������0�=AM?!����8�����)k>�x7?���>���>���U(���r�<%�>߷
? :�>m����pr�8X�M�>���?��\=��)>���=�慼hӺ96�=D���-�=I���`
;� <�w�=/
�=u�6�Ź��:���;Ԏ�<-?k�?Agj> t>����.��T��`>�-S>�Kt>��H>�վ�T���s��)lk�}a>;�?�f�?|�=o��=��=�a��LT����;��=�Y?��!?r�M?ᦓ?�E?�^!?²�=���g�����~�Ģ���?w!,?	��>�����ʾ��։3�ڝ?h[?�<a����;)�ݐ¾�Խѱ>�[/�h/~����=D��텻���W��6��?�?HA�W�6��x�ۿ���[��z�C?"�>Y�>��>T�)�}�g�s%��1;>���>kR?�!�>,�O?�;{?1�[?�kT>��8��/���ҙ�323���!>�@?ð�?��?*y?v�>��>��)����R������XႾUW=�Z>E��>�'�>��>T��=� Ƚ[P����>�g�=;�b>;��>���>�>s�w>SM�<KaH?��>���������-$��*A��v?�̏?�,?��6=V���F��V��+,�>��?�R�?;~,?�WM� |�=��ۼ8�����k� ж>�	�>8��>5ե=nEM=�>��>Iw�>�(�u���5���2�6_?�PD?��=5�ſ�q��k��q���jx<a7����`������w[��=z������'k���	]��렾]���'ߴ��ܛ��~z����>�=�=Sm�=2�<kJ�����<B�K=Gl�<�!=��j��y<�Z=�����ȑ���M�#Lb<�$J=�g�m�˾D'}?�
I?�\+?��C?A�x>��>~�2��R�>�����E?ĳV>�M�؎���p:��.��yꔾ�ؾ�־��c�J����>�K��>"3>w��=�m�<<�=��s=|I�=����=���=���=E�=�?�=��>�!>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>ǽ5>WE>�Q�T�0��+Y�VDd�Z�W�~!?�:�JN̾��>Eؿ=^ݾ��ƾ�9=�)8>}b=����Z���=�[|�a�4=a=�>rVC>�v�=롪�H��=��K=l��=��T>Ӂ���C��#���-==��=��d>e�$>_q�>��?�a0?iUd?AH�>��m�~�ξU3���L�>E��=�3�><b�=ՎB>���>o�7?H�D?A�K?8R�>1��=I�>��>s�,���m��d�ǧ���<+��?�̆?�̸>/�V<UUA�����f>��@ŽXe?E1??U?�۞>�|���㿧��s\.���{���(=��8=�tk�U�ͽm�����AԀ�C�>�*�>���>��>��n>J.A>Q�X>]/�>�m�=��Y=i�>��`<��V�e&�;���<���=����ԍ��z=Z�t�Q?����=�"v�<�ȼ�{�;�a�=��>��>@��>i��=ﳾpd/>����p�L�@:�=d���$B��$d��F~��	/�	`6���B>'X>����-��T�?y�Y>UE?>h|�?/Iu?��>#��`�վY��e�%qS��;�=!�>�#=�ʁ;��M`��M�rgҾ���>Lߎ>t�>׺l>�,�g#?�^�w=�b5�N�>G|��-��*��9q�"@�����Ui��Һ�D?oF��՝�="~?��I?�?���>���݆ؾ�:0>�H����=a�_)q��f����?�'?���>����D�ֿC�J����U>ڷ����T������T�_G=5���+�>w瘾5ݾ3&`������o���_� ��-=?�yh?2��?u1ɼbS���V�1e;�?k�� -?��S?%�>v3?^?sq���E���4���>�=:�_?y��?
�?�֓=�ީ=2������>ap?@ŕ??A�?��q?�Q6�0��>N��;TN>�uսZ�=�>���=��=�K?�?��?�,��b�
�=��~T�QX���<�]�=�:�>x��>�Zx>\�>�X=�f�=hoX>��>�ކ>͘X>�K�>�T�>T���@����/?��>j��>?l??�S�>���=H�b��e~��KϽ�7t���<��&����	�4s��]>�<7��=�Y��|.�>��ÿk�?��n>m��?�=��_�g;>z�}>8���_��>��@>��>�q�>>� >�,f>g&>�ԾM�>1��S� ��iB��Q�:<оw�z>�{����(�P5	������G�N�C���i��灿v�<�K��<�?����j���)�����8	?�,�>��6?/W��=�����>�`�>ؾ�>���1���>׍�o���?O~�?�8c>��>��W?�?/�1�3��tZ�W�u��(A�le���`�=፿�����
����i�_?n�x?�xA?WI�<�9z>���?(�%��ӏ�t)�>~/��&;�IQ<=5-�>�,��
�`��Ӿ��þ69�(FF>8�o?�$�?�Y?�RV�~B%�(lN�Od?,(�>�s?.��>�RB?.mD��R�>�D>V?墾>K�8?���>�6?��f>�>�8��Br)>�?��rzf�ɔ�w�V�B
��Ұ7=k^����f;o�<����c�=�8>I�ս)j� 7G�\�i��Lu=	[@>r��>�4�>�w_?}��>��>��7?���U�2��޶�d�2?p��=���r����������}�>�[l?���?z�S?�gI>g�E�ޚL�ע)>��>�:3>Z�H>�3�>�ؽd�E�5&�=��>��>�$�=RI^��w��
�	��!����n<F�>m��>��}>�����N'>����U�z��ud>	�S�C5��_�Q�F�G��z1��v���>��K?�"?P�=������/f��(?L�<?��M?,�?�i�=�H۾B�9���J�Ǟ����>�ө<v��K���������:�$��:��s>T�����B�g>�#��۾@n���I���㾗�5=���T=vW��־w�{����=�> ���P���I���:��h�J?f�k=A���O������>�.�>�{�>ڲ0��EZ�Ea>�`����m�=��>1�7>/x��E�I�E�ږ�
>�>VQE?IW_?k�?-"��Ls��B�����yc���ȼ!�?(x�>h?�B>���=Q�������d��G���>���>g��#�G��;��0��P�$����>O9?+�>}�?A�R?{�
?c�`?�*?9E?'�>�������B&?ሃ?ׄ=l�Խ7�T�Q�8�.F����>	�)?��B����>.�?�?S�&?ۄQ?�?��>�� ��E@�䑕>_\�>��W�]a���`>�J?��>(:Y?�ԃ?��=>�5�,䢾f᩽+d�=^>��2?�7#?F�?쪸>���>�����`�=|��>�c?�0�?|�o?\��=��?"52>��>��=���>7��>�?VSO??�s?��J?s|�>���<�z��~.����s��>Q�Y��;m[I<��y=_}��1t��a���<} �;�������q��E�B(�����;�_�>��s>&��%�0>}�ľ�O��S�@>b����N��jي�z�:���=ކ�>��?a��>@V#��=��>UH�>8���6(?7�?x?��!;סb���ھ��K���>�B?���=�l�-�����u���g=/�m?��^?�W�"&��K0i?�1??v��k�>��+��9"�T�D�?��?�C����>v�?��N?�A?";��B�7��N���{�{H}�e*o=(�>؅��we����>�1?�>��.�g7>]�*�" �����=�?S�?{�?}@�?��">x��P�����1I��)�^?��>����}'?��L�Ǿ���Ì���ݾ����J����������.�N0��M4�t��=�?&�k?�m?l�Z?B���Cd�y�d��|��GW��I��D���=���F�6�C��q�����;�������A�=�d��Q�Җ�?t8$?��U��?㩾�Ҿ~���s�4>T���_o���=m+���8=��I<K݀�U�P��;���/?1͗>��>e�0?�j��<���I��H2�&���b>8�>	�>p�>#�>��|���W�޾R�.�Q�X��7v>�xc?U�K?��n?5p�+1�����Z�!���/��c����B>�j>:��>�W����F:&�gY>�A�r�n��w��>�	��~=��2?z(�>A��>�O�?�?�{	��k��lx�>�1�ڔ�<41�>� i?A�>$�>�н-� �E��>�cj?B��>^8�>e���H0"�̓{��w��G�>��>��>I3h>]5:��\�!Ď������29���=�fj?������_��Ɔ>zQ?&�.;G<�s�>�q��6J��%�-H&��;>�?�?�=U�8>A�ƾf���+|�Pȉ�u�&?��?�g���((��!�>lB?�+�>vS�>&*�?	�>�KѾ�E�=�?��_?��I?�`G?���>H�3=�Q��i޽;�"�
��=E׫>�
U>���<wL>��'�bjQ�����t=<�=1��;y �'�<�e#=�l�=+�,>-�߿r�D��R����	��V�(�T-N�y[V�W5��ś��~�Ծ�_���h����*lG:��n��8P��9��1�l�֑�?���?��	�(��y����w�tѾ$��>�b���v�<é��������+ھ��������>��H��d�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<	-����뾭����οA�����^?���>��/��p��>ݥ�>�X>�Hq>����螾|1�<��?7�-?��>Ŏr�1�ɿc���v¤<���?0�@}A?��(�����V=-��>�	?��?>T1��I�����yT�>{<�?���?~M=e�W���	��e?Lu<�F��ݻ|�=�;�=HF=>����J>�U�>%��OSA��?ܽ��4>Mڅ>W~"����W�^�]��<�]>��ս�;��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=k�Q�ƿP�$��s��� =����Z�M���諽��Z�v���o�
t� ~h=��=��P>�M�>2VV>��Y>_~W?A=l?�>\N>�T�i�����;>�	��v���/�Ú��h���Σ�1C��p߾Ox	�������Iʾ9!=�@�=b6R�/���+� �,�b��F�^�.?%v$>�ʾ��M�@�-<pʾ	���nԄ�V᥽�-̾�1�"n�]͟?<�A?������V����rN�ц����W?�O�~��Bꬾ���=}�����=�$�>�=-�⾋ 3�M~S���/?�W ?�6¾GT����->_D� =G�'?!
?���<j�>��'?q�(��ҽ.�_>�R=>�ߣ>��>(� >D:����ڽ��?!�W?����}��B�>���٩w�}<_=^	>�'@�06��ZtQ>�L�<�k���'��Hw��@�<K�Y?@�w>�#7��a�Ó����8ʲ���s?�N�>l�>:+i?��"?h���L�fpS�n�����=1�]?`Yu?�Q�=�m$��[����c�m%M?�+V?	>�=�����پ�y
����xm?�5]?#;+?Y��=t!���H���d���.?Ly?9aR����'	�LY���D>�a�>��?�<��͟>{fX?��W����+ƿ��I���?V@c%�? ��=����r�=���>�-�>�D��f���i���޾���=���>7ݹ��\�����?�hOI?�_?�m�>~;m�3����=�镾=Z�?8�?������h<���l��z��RƠ<�ݫ=����9"������7�D�ƾԿ
�>����������>�W@&\轐#�>�]8��6⿇TϿ����Vо,6q���?�}�>�ȽS���u�j�"Ou�>�G�1�H�����`I�>��>]�������~�{�0q;�L����>��
�>��S��'������}5<��>��>��>�+���罾ř?%d��j?ο&���ϛ���X?�f�?�o�?<p?\�9<��v���{�
r�-G?�s?#Z?sm%��<]�{�7�1�j?^���U`��4��EE���T>�3?�J�>�-�.$}=b0>�{�>�=>&/�όĿrڶ�������?~��?�f����>H}�?Ho+?Kh��4��@V����*�<
��7A?�2>g���ð!�)=��Ւ���
?(y0?
��u-�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?Z$�> �?�m�=�a�>�d�=R�%-��j#>A$�=��>�Р?ŨM?�K�>MX�=��8�1/�[F��GR�n$�3�C���>��a?0�L?uKb>����2��!��uͽd1�RN��X@��,���߽S(5>g�=>G>��D��Ӿ!H?e	��'ؿ^K��,�S
2?.�>�=?v�)Fq�V���]?�g�>.���~��)�4� ����?�3�?w�?�־�����4>o��>&��>~7ǽ�0�������1>h�B?�C�="���4p��օ>��?t�@��?jh�|B?0���.���\F|�K�����I �=��Y?w�����>�?�3�;F�>��e���{�>�5�?5��?�?�[?�lV��xJ�e��<�U�>�JE?%R?�=�~���<=�$
?C����������TS?7"@:@h?C?W����D˿����/���;��w/o=?��>�@�>��߽렒����<`�C><N>�>�>K3{>8'�>
U>
M'>$�i>�_y����c"��Ib���9a��-�C$�z�J�e
�)[7�4˾-���p鲾�U7�Y!����|�[�RAG�1�>�̣�=6W?=U?&�x?�R	?57�|I<>�3��)��=<d*��o&<[�`>�7?8M?�N1?��=����K]��U���r�����:��>`�)>�f�>�`�>�T�>s3=��=>Y>��[>��	>=z*<�o꼚�.=��F>���>���>�q�>�C<>��>Fϴ��1��j�h��
w�{̽0�?~���T�J��1���9��Ҧ���h�=Hb.?|>���?пf����2H?#���y)���+���>|�0?�cW?�>����T�(:>3����j�:`>�+ �vl���)��%Q>ul?�f>�u>ț3�ge8�\�P��|���i|>�36?O鶾�C9���u���H��cݾ;HM>�ľ>(D��k�m������ui�י{=Qx:?�?�6���ⰾA�u�fC���PR>�:\>�U=�h�=�XM>Ybc��ƽ8H�Ug.=<��=��^>��?��*>���=��>��E�R���>[&D> �)>�@?{@%?���"h��8����t/��Ip>f�>�ŀ>�P
>7"I��!�=1�>��a>�|
�'h��Xq�!J@�HB\>2�x�ؑ]�=)t����=
u���l�=ǔ=n���:?�[=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>�x�uZ��u����u�y�#=���>�8H?�V���O�>��v
?q?$_�੤���ȿ"|v����>O�?���?�m�yA���@���>���?�gY?\oi>�f۾�`Z�ዌ>��@?�R?��>�9�2�'�|�?�޶?���?D-I>���?��s?Cg�>c"x�^/�*4�������=��g;m�>P;>����1iF��Փ�m���j����b>T�$=A�>�#�x*��f�=�㋽�J����f�M��>75q>��I>lQ�>�� ?�k�>��>�w=䰋�������D?�W�?��(�{~�4��=�=}����O�>�AK?�����X)?xQ:?W��?e�M?�?�U�2^��l����l���r�=M�\>�?K��>P���>����s��r�>)��=D�`��=ʾ-Q��(��=
��>�Z:?f#?��>�
+?�/?���=e7�>�K9�����<�J����>���>��+?x��?I��>� ���8��ː�>���^�l�5>��?'?���>0@�ȥ��qOʽ_�<`����Q?���?�N�)j?>&�?^?hG?�B�=�1���� 2�\��=��!?��A�}M&�?��|?�N?���>g:���ս39ּ��8�����?l'\?J?&?����+a��¾r:�<��"�KtU���;!}D���>[�>����⚴=�>Ұ=pMm�
C6��/g<gj�=��>k��=17��z����/?����������U= Fs��I��Ke>�4y>����V?E���4�x��H���g���9|��!�?
��?�d�?+�+��`�۬8?L�?�?��?��00꾬$��scc�a_����� >u�>!K <������/�8������0e���>��>a�?p# ?��M>�ݱ>�˘�['�L�w���^�vk��R8�su.���񠾴#��a�L���|��>Z�����>��
?�cf>�}>4��>�x���j�>\�Q>�*�>���>s�V>��4>�� >G:<�ѽ�KR?����$�'��������g3B?�qd?R1�>li�<��������?���?Ts�?=v>
h��,+�n?�>�>H��Wq
?{T:=9�-;�<V��x��3���/��>E׽� :��M�Anf�xj
?�/?�����̾�;׽q�j�&s���-�?�?Ag=�*�-������:��i�Xa�=���'��}��nf�z�������i=��Q��g~=��5?x��?o�#����о1����=���h>�T?6�>iU�>@@�=��3�^<��Iv�4�(�ӿ���"?Q[�?x�->Ia?� ?�Q~?cP?�	>p�>�^��-?^�]�M��<���>��O?U�6?��C?1�+?��<?O._>�ƨ�)C���8���Q?P�.??/��>�y?��սZ�ӽ�;�Ud����
��*�=�>�<��=V�A�d��<L�M�n��=��?
����;�#�뾪�g>�d"?3��>D��>2�����7�f�W= �>�!�>��^>�� �T+��R�����>ܾ�?j�˼�F�<�l9>u��=�C��HC��\�=�G����=�v�<2&���%����=��=��Q��ܼ�Rt�0LY��J(<jw�>�?T��>�A�>�@��ū �Ӷ��v�=�Y>�"S>�>�Fپ�~���$��+�g��Jy>v�?�y�?��f=��=��=�y���P��U������D��</�?�J#?VWT?7��?}�=?Ej#?�>�(�)M��@_������?�!,?抑>���v�ʾ���3���?m[?�<a�+��r;)��¾��Խ
�>�[/��/~����D�Z̅����T����?ٿ�?3A�6�6��x�ɿ��`[��t�C?�!�>�X�>��>�)�c�g�i%��0;>r��>=R?�#�>��O?p<{?��[?hT>`�8�b1���ә�N83���!>�@?��?��?}y?�t�>D�>��)��ྷT�����-�����W= 	Z>&��>)�>�>���=�Ƚ3Z����>��a�=?�b>R��>c��>��>��w>[L�<�G?���>`�����𤾞ʃ��=���u?#��?Đ+?��=����E��K���B�>�n�?��?�5*?��S�3��=�ּ㶾(�q��%�>�ٹ>1�>I��=�F=�\>	�>}��>�+��a��n8�sCM�w�?xF?4��=�`ſ
C��Ӗ�Yw�תr�����Q���5 ��W���Q@=�/����L���RM���_�[/������͞�� ē�۩?�b�=յ=�h>+)m=�c�=������o>�1=f"	>�p��,�D<��8���"�����UZ��[6<�&�=��"��˾��}?>I?��+?��C?G�y>�F>��3�t��>�y���8?�V>1tP������o;�񩨾���W�ؾ�{׾V�c��͟��7>CPI���>yW3>�$�=붉<��=�As=1ӎ=��Q��"=��=52�=t]�=f��=
�>�S>�6w?X�������4Q��Z罥�:?�8�>g{�=��ƾq@?��>>�2������yb��-?���?�T�?>�??ti��d�>M���㎽�q�=H����=2>p��=x�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��7>�>_�R���1���\���b���Z�Ɲ!?IH;�/̾g@�>`ֺ=�=߾��ƾp(.=�F6>[�a=�`�QD\���=��z��;=�l=5̉>Q�C>.X�=D���Z�=��I=���=;�O>���>Q7�?u,���3=���=��b>��%>H��>��?�a0?�Xd?6�>�n��Ͼ�?���I�>H�=�E�>���=sB>0��>t�7?��D?��K?��>���=[	�>��>2�,��m�2m�[̧�/��<���?�Ά?_Ҹ>D�Q<ޏA�����g>�/Ž�v?<S1?�k?��>�U����9Y&���.�$���s|4��+=�mr��QU�M���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=$�����<�vż�����u&�:�+�2�����;r��;B�]<^��;���=c��>R>���>z��=���Z0/>�����L��ӿ=,<���*B�=9d��L~�|/�'v6��B>�JX>/7��,1��|�?=�Y>�x?>���?�<u?Z�>G2�o�վ�K��VTe��QS�Ը=��>S�<���;��a`���M�FsҾ��>6ڎ>���>P�l>�	,��$?�%�w=t�a5���>q��r���D��9q��>������#i�^wѺi�D??C��Θ�=�~?3�I?{ޏ?1��><&��s�ؾ[0>)C����=T	��q��;���?�'?��>�쾜�D�u��=����>Y�h�`�z���?��x�=��˾�z?As8����AC�N,���S��CtS�����^?h�c?h�?�Z��$[��7�P����Uݍ��i+?��z?R�>.�>p�
?�!��T�go��󸼽B�a?W�?c��?�3�>��=Y崽���>C	?ߖ?ɳ�?y�s?��>�A��>�|�;w^>hH�����=}0>B@�=&��=��?z3
?k_
?�T����	��y�m)�}^����<�ޢ=l�>�+�>�%r>���=�ai=G+�=> \>(�>�E�>��c>K��>Pۉ>�-ξ������+?�j>�	j><�8?�n>� >9�$���=�ս�u��-EὙח�ތ{�.�$�=�V�D����ި�E:?g�ʿ)�{?
U>C*����<?d�"��S�=�';� :>��kf�>��2>�Y>Gj>���>v��=� ]>��2>6WӾҌ>|���X!�(C��wR�}�Ѿ�sz>磜�A�%�h��~���^-I�%g��`[��j��(��g6=���<H�?>���k�K�)�;�����?6�>�&6?�ی��ވ�R�>���>;��>�>��o���n��`ᾓ
�?���?�;c>��>I�W?�?ْ1�33�vZ�,�u�n(A�-e�V�`��፿�����
����.�_?�x?2yA?�R�<.:z>R��?��%�[ӏ��)�>�/�'';�@<=u+�>*��/�`���Ӿ��þ�7��HF>��o?<%�?wY?@TV�2_���ۚ=�oZ?�=3?D��?k�I?��h?�Z��� "?�V�=�f�>�>�>w�H?��&?��*?ۍc>�.^>��
�_ŧ��㦽�tþ�=���y�-����R�=HH�=I)��N��e�=*N{>��<�84�鶟<y�����{���:�ꀔ>ө�>]�]?l�>��>��7?Z��"S8�b����?/?�i:=!낾Ȋ�l���߳�n>��j?��?OJZ?�c>�A��C�q�>ٚ�>p�&>��[>q��>*G��~E����=�9>�>��=�O�X���8�	��W��j�<>���>`3|>x���'>�{��E1z�7�d>��Q�|ʺ���S���G�}�1���v�FZ�>:�K?(�?���=W^�1��*If��/)?R^<?�OM?N�?�
�=��۾x�9�{�J�Y@���>L4�<�������i#����:��:��s>�1���	��cJt>���s�Ѿ/�h��V�+��E(�=���*��[_�%��$m��i�=t��=�����"�㵝�����aF?��$=�8���h��3���J6>wZ>a[�>23��D��g7��i��Q��=:��>�� >�=W�:+B�@���=�>hPE?}W_?�j�?+ ��ks���B����zc���ȼ��?{v�>h?�B>��=������d�UG���>��>���Z�G�;��K/����$�0��>�7?�>e�?$�R?��
?��`?Q*?yD?q%�>�� ���{�3?��?����9�)�~�v�$A:��WV�	f?��"?�����XL>��?3�?�.-?�Z<?��&?pI=N"���R���>�;�>��R�����K[u>@�X?o_�>��G?��?4�>��0����~�r���<>o�>�@?��+?��,?��>��>/�ھRU�<,@8�;4b?�d�?�Vt?I�[>� �>�j\=<��>�#<���>^?�E�>��>'�??xcX?c�?�*�<~��x4ѽ���F[<*=gD�=Ft=�a����>�*����?6�"a �b;½�a(=Zl���D��`g=ܕ#��5�>+
t>�ו�-0>�ľ�+����@>X���Λ�������9�j��=���>�?�P�>�,"��=�]�>��>����	(?�?��?��4;˥b���۾��L�-��>��A?��=��l�T[��"v���f=t�m?Ӕ^?'�U������;f?�F^?l�o��t��z�о{�8�E?��>��� @>�?`�U?�y�>�#X��Bb�#���Ƥ��%	žg�D=��H>���h|W���>(z'?�֣> @�>���=�)��?��h��&?��?U��?1V�?��>�r�;������䉿'4Z?a��>�ƾW�?������������bz���q���<��Lv��!���F{��VZ��|���%ｧ	�=p�,?ߙo?�m?� k?�.�~�b�n�h��x�TU�f�۾����B:�K":���7�Y�y�����v�Ⱦ����Ra���4����?�@5?�����>�O��ةþ��Ծb_>V��� �D��=���cC���%�Zo�4�V�Tz��\�@?w7>�>�iK?%ك��>L���S�H�V�����Z�>�1�>4�>�Z�>��<�5��9=�}��LK;?�:��[v>�xc?{sK?Z�n?Yy�91�߆��e�!��b0��S��o�B>��>t��>��W�2��/9&��Y>��s����w��1�	�N�~=;�2?�:�>V��>�G�?�?�s	�~�����x�&�1�:�<�]�>Pi?cu�>o��>qgнl� �	��>d�l?s[�>7�>_����z!��{�jͽ}��>+Q�>�>2.q>��-� S\��^�������U9�Y��=p�h?Oz���`�ˉ�>�Q?,_�:�C<^��>u�r�!����0�(���>$�?,Ī=�^<>�zž�����{�����F�(?5[?���&�*��n>D`"?��>�B�>�܃?��>����L��?��^?��I?�n@?TB�>�'=�f����ǽv�&�(=�Æ>�[>g�p=(��=���o�\�?���wI=�ּ=�Լ�����?<���%�M<
K�<H�2>�#ؿEF�Lƾ�����4������ł��A���8���ҾO����k�o��m��ߊo���c���u��S�X��?/�?p�F��)9�⓿��s��P��b��>uga�����+ǰ�;��hQ����ھ2�߾V"��tQ��m��Tc�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@�zA?t�(���/V=��>B�	?T�?>ZK1��I�����JX�>`;�?��?w�M=R�W�n�	�~e?��<��F�@�޻��=�9�=..=�����J>�J�>��nLA��aܽ�4>uڅ>ca"���֋^��<��]>޶սGA��5Մ?#{\��f���/��T���T>��T?�*�>�:�=��,?T7H�`}Ͽ�\��*a?�0�?���?(�(?2ۿ��ؚ>��ܾ��M?dD6?���>�d&��t���=6ἲ�������&V����=Z��>T�>��,�ߋ���O��I��g��=��������g���@�绿���
�	�$�����Dc׽�%ʾh�W���Ƚ�V�<o{>� >�̓>��>�ہ>,�]?�l�?���>��>q>۽)ʋ�j�˾o�u=>�����T�v����(�����ž��k����#�����վ	~;���= �R����ڛ ���c� G���/?�p >�u̾�5N���I<�gɾp&��ό��墽u;�3��Co��t�?bA?+���"FW�6�PU𼝇����W?N� �,��^B�����=rȟ�/Q+=���>���=W���2��S��x0?� ?�R��t����/>l�	��*�<��)?�O?=�a<���>�#?��/�)>�f>�B>^�>�q�>�	>�{��z�潴T!?SlW?+d������ۖ>�ٻ�����+;=�>�.�!޶�X>�x�<����B�g��刽���<{(W?A��>��)��Va��J��7Z==��x?��?C.�>v{k?��B?�פ<�g��d�S����`w= �W?>*i?��>뇁��	оP���R�5?ѣe?��N>�bh�(���.�AU��$?�n?_?�{��w}�d��p���n6?��v?s^�xs�����J�V�d=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�%Þ?��@���?<�;< �U��=�;?o\�>��O��>ƾ�z������+�q=�"�>���ev����
R,�g�8?ݠ�?���>������+H�=����ڬ�?	A�?,���Ed7<���G�l����s��<�m�=Dh���!���y:���ȾdK��H���[��R>�>z@���+�>��B�6�㿪pѿ5����TԾ��\���?˳�>�$����٨l���q���K�isH� ��Bf�>�>~b���ꑾ9�{���;�:���Y*�>����>@�S����y���1�4<�ג>G��>��>�;��:��f��?�]���3οu������S�X?dY�?s�?}p?x3<��v�%�{�ls�AG?�us?�2Z?<%�nH]�w�8�%�j?�_��xU`��4�wHE��U>�"3?�B�>U�-���|=�>���>
g>�#/�x�Ŀ�ٶ�E���Y��?��?�o���>p��?ss+?�i�8���[����*��+��<A?�2>���E�!�B0=�OҒ���
?W~0?{�g.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>��?��=	X�>���=x԰�t'���#>���=�?��?2�M?6g�>���=��8�</��GF�oFR��'�C�P�>k�a?alL?�Lb>�����3��!��4ͽ��1�o���@���+��;�~�4>� >>T$>$�D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?qQo���i�B>��?"������L��f?�
@u@a�^?*,Ϳ����5٪�8"��~>]��=��>>�Pν�*�=5�=����;o�>'��>��W>L^>�Lk>�78>�\>5����S#�R��ħ���sG�m�����0�]����g̃�K���<��0�þ=8ɽ��_��(����;�"�"�m¢�ne�=}�N?a�P?6k?�b?�+8�qKA>B���O<2���=��>�5?��O?�'?Ů�=�`��yd��|� ���������>�9>Ip�>G��>6w�>�H�vEG>�8>�nt>o}>��z=�?ּo��9)�_>�N�>�S�>�F�>�͚>g�T>O�������$c�3ݿ�e聾p#�?ݰ��d^�/֔�U�I�|����=�=K?�X>�ޑ��#ٿܷ��C?!�\��3�w����m�=7-I?:'?myD>�g��撽X;>\��Q����>s�����<- �,�o>,J?��f>Wu>��3��d8���P�c���c|>�46?�궾@I9��u�3�H��aݾHM>Jþ>��C�6l����3�.si���{=Pw:?߂?�:���߰��u��@��2SR>�3\>�T=e�=NZM>eEc���ƽ�H�_.=��={�^>�?-*>�	�=bg�>����FM�1t�>��C>�Z(>�??��%?	��5���c���F-�c�u>6�>��}>E�>��L�ܽ�=��>��^>�s�f���c��I�@�!�W>����W_�~�i�!��=�r��?>�=y�=�I���S9��!=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾMh�>ux��Z�������u���#=S��>�8H?�V����O�i>��v
?�?�^�੤���ȿ4|v����>W�?���?j�m��A���@����>:��?�gY?noi>�g۾6`Z����>л@?�R?�>�9�~�'���?�޶?կ�?%�K>���?:Zr?F�>v���m0�����&���q=��<Eʒ>�>�þE�G�Y���ǉ��l����dlf>#=H�>N3�ƻ�_�=ӓ��L���oa���>Wp>�E>Z=�>��?���>�?�>Es=!���`���i�[?�ϑ?ؒ9�vȂ��g,�C|�<c;]U"?��W?��<8�	���>`T?�[�?B!8?#�>���R��&y¿��;ԥ>��N>J��>5�?^����&;>� �|	>#0�>��>� ���uɈ���=hi�>�ya?~'5?x�=*9?�&-?�ߢ=�|�>Zr��윿S�g��J��>�6^?�ݖ?l�e? S�}�z�u؜�T|���y�� 	�N%�?��?��><ؖ�1"���&�=X(
���>v�G?pG?!Լ#�?���?;\+?���>�N?����8qо�g���>��!?�)�ʳA��O&�_����?UT?���>:/����սZ�ռ����r��F ?�"\?;8&?���a�j�¾�*�<b�"�sUV�ww�;ԓE��>��>+z��ވ�=�>8��=�]m�;^6���f<���=v�>Z�=�7��n��G?,?*~��ܚ���^�=�kq���D���|>��J>R���T�]?�>;��s{��Ԭ�fQ��ʏO��O�?-��?lM�?�\����h���;?ͳ�?hF?�6�>^�۾.j߾�:|�!{�6��>]��>��o�A�〤�p)��W����ký�-W�i:?�b?\s?���>
O>���>!�6��m�6n���C�H�c�;�ύJ���&� ������H�^����(G�ӛ�>��&��>�Z"?ª�>�n�>��>k缶��>M��>�9`>�>m>gRe>�*�=��>fU=8"��JR?����7�'��辻����3B?�qd?1�>Ji�����!���?\��?�r�?D<v>~h�R++��n?�?�>����p
?�Q:=�5��L�<�T��l���3����ɩ�>UE׽f:�FM��pf��i
?/?)
����̾�?׽>��+a=Q�{?��O?lo��O���|�m&d�ipm����=�Ɉ��%L��4/�^Ol�������z�OA��i�;�j
����=?�ԕ?�*�ö��W?�矅�sag���
=n'�>C��>�f?���>��M�q�H��<n�?��t��Ϩ>O�m?s{�>��Z?��M?⅋?�p>?�,%>Tf�>�̨�SV?���}+�>s[t>��?��>�Xi?�V%?�wG?mU�>.t�F��/z ��m\?�H�>0��>��B?�]?�����f����;a�&�29)���*>0�f>�����O����?�,@����^>�i?tab���!������>gOG?w�?���>X�B�g@�����=�h�>�?���>k�ξn�Z��h۾�H?<��?me���<�>x׋=b1w<	׆<��=�m���=�@<���b��=@��;��5���B�<+�p=-6��t�>8�?���>�C�>�@��,� �`�� f�=�Y>$S>l>�Eپ�}���$��u�g��]y>�w�?�z�?ػf=��=Җ�= }���U�����;���u��<�?;J#?$XT?_��?z�=?]j#?˵>	+�iM���^�������?x!,?
��>�����ʾ��׉3�ٝ?e[?�<a����;)�א¾�ԽƱ>�[/�j/~����>D��셻���R��4��?쿝?AA�W�6��x�ڿ���[��z�C?�!�>Y�>��>T�)�z�g�s%��1;>���>iR?�"�>{�O?%={?a�[?�iT>Ǜ8�0���ҙ��P3�A�!>k@?��?��?.y?[u�>(�>j�)�6�nR��h���q₾��V=�Z>���>M(�>��>��=��ǽIS��>�>��_�=�b>���>��>� �>�w>�I�<jVP?�8"?�J�$���<������h��39X?��?��J?�)һ���:-D���ľ���>��?t�?��/?����a�R��<�!P�0�>��?+�>Q~�>�� ��^=1��=�?h�">�}���AK�Ǿ�c�;-5/?z�@?(�5>��ſ[q�o)o�Wg��,m^<�o��7d��@����Z��ˠ=�����f�n���6w\�@��7����q�����G�z�W��>�#�=�z�=���=7H�<Y+¼���<4M=�R�</�=o�m�R��<1�8��仪���w�W�6)^<\�J=�,ػq�˾;b}?� J?�:+?�B?�z>�">�� �X�>'w����?~U>TL��7����?�V�������U׾=־ija����>�M� �>V�7>�n�=��<Z��=c�r=���=�Ϻ�f=�S�=��=�X�=G��=�>~l>�6w?W�������4Q��Z罤�:?�8�>c{�=��ƾq@?��>>�2������yb��-?���?�T�?>�?Bti��d�>M���㎽�q�=G����=2>w��=x�2�R��>��J>���K��D����4�?��@��??�ዿТϿ8a/>N�7><>F�R��1��o\��zb��ZZ�.�!?Y=;��5̾�=�>�=��޾�mƾ.=�r6>O�b=�o��P\��ٙ=k{�;=�ck=�É>�	D>�w�=}����=9TI=���=��O>jݘ�!�6��,�)�3=��=I�b>�%>�j�>��?�f0?[>d?�Y�>�m���ξ^��F�>��=-j�>s%�= C>ң�>c�7?��D?\�K?�^�>4��=Kֺ>��>	�,���m�z�ڧ�ĥ<4��?�͆?���>��M<9�A����gp>��Ž	?IF1?\t?ƞ>�	���ݿcv��w�]k��+� >ic>���Ch9���2������ 
�2�b���=��>��>�c�>E��>�Q�>���>W�>�B�<�������;��
N�}�(��><�л<��齄�=Ry�<Tɽ�f���;6��"=�>#��=]��>Q=>:��>ю�=����C/>w�����L����=JH��Q,B��4d�sI~�X/��V6�H�B>�:X>�}��4����?��Y>m?>r��?VAu?��>��.�վ�Q��XCe�'US��˸=��>��<��z;��Z`�<�M�&|Ҿ5��>�E�>9��=���>�bB�!�c�e���$�lC�L�$?0��!�> ���!9��� �������6��JY�C(@?��z�O\�=�X??��;?�5�?��>�z��a5����3>�ʾ����T,�[�=���=xT?�aC?�W6?�V��킿jJ̾�辽��>2I�Z�O�H����0����aŷ��{�>k �� �о!3�(g�������B�PPr�t��>��O?'�?�Fb��U���OO�t��V���q?#yg?��>I?EC?���yt�Xq��ކ�=N�n?��?�8�?T>��=�3����?2�?l�?�d�?�~k?����J�>ǖ�=�Qs>D����F>IU>Y>���=C�?r�>Y?�Fý�D����d�8Gk�*��;)�>]�>�G�=���>zpB>	��<I�8=II�>��v>9>�n>�4,>3{>����w�!3?�>EY>��4?.6�>�>>2f�n������P)��$�E����>�4d��34ʼJI�=��z<L0�>q�ʿ!��?�g�>����??���c��=�{>�U��N�>f�;>A�{>`)�>�#�>ƽ>&g:>�>�IӾ��>����Y!�Y*C�}R�Y�Ѿ2�z>4����,&�*��a���@I�
t���o�*j�&,��U7=����<�F�?uy��/�k�R�)�����=�?�_�>u6?�ǌ�
����>H��>�Í>oM������ō�Ba�,�?���?o;c>��>S�W?'�?�1�13��uZ�	�u�a(A�4e�f�`��፿�����
�����_?��x?yA?QR�<Z:z>Z��?��%�Lӏ��)�>�/�';�rA<=�+�>*����`�H�Ӿy�þ68��HF>t�o?/%�?lY?)TV��-��'�{��2?WIV>ʗZ?�	.?�5B?�ޘ��5�>��=��"?�0�>q6E?�*D?���>�*�=Iq�>I������;w
��/���aX��ZR�5MD�Ţ_=�S���<tCU=W����M��"�;���<���<+�w��<�<�;C�=��=h��>�`q?
U�>!�>�???�����1?�B����V?�g�=g�&�D��\Ⱦw� ����>8օ?�]�?\rW?g�>�񆾨���@[�>E�?�#�=�zQ>���>gȽ#*���z���>WQ>©>�d�4���]��A����}>=y�P>���>��|>MR���(>�E���hz�Ord>��Q�u���S���G�%�1���v�P4�>��K?�?�b�=L.�Lf���If��)?�}<?bM?�?9�=z�۾\�9���J����h�>�_�<�����������:�X,�:��s>���'L����b>��
��oݾ$�m�ӳI�#c�2=C=^a��T=�Q�J�վF�|�^�=�
>����B!�73��h����I?kv=�����V��+��y�>T
�>�ݮ>Qq2��^|��F@�wu���J�=���>[�9>���&N���F�'�����>NE?�o_?a�?ł�o�r�֬B�� ���Z��Òɼݞ?'V�>c�?e�A>���=(���s!��e�.G�r��>���>���/�G�����~��!e$���>�X?��>R�?��R?'�
?9O`?U�)?��?|Ґ>@綽ӷ��#B&?%��?<�=J�Խ��T�A 9�>F�>��>��)?:�B�X��>�?Խ?M�&?�Q?�?R�>�� �+D@���>�Y�>T�W�Yb��V�_>)�J?w��>�<Y?�ԃ?��=>��5��ꢾ�ש�sW�=>��2?�6#?Z�?��>��>�릾��=��>�,d?���?V�n?�U�=���>�>�O�>V&�=b�>���>s�?йM??�r?�I?�b�>���<:���Ͻp'f�v^<Lk5;K㻮zV=�%����]��lw���<��;B�¼����ȟ�^+��μ� <�G�>��s>���1>��ľUH����@>����9S���抾��:���=N��>X ?r��>�E#�B�=���>�J�>m��L<(?S�?2?�{/;P�b�	۾��K�6�>�B?Y�=�l��~��m�u�\�g=L�m?Ǉ^?դW����#-p?�H?���W�P��,׾�U������@?N� ?g�;ka�>�(v?a$F?y��>�	��+NA�朿��i��fy�E��<��>�%�"o�}4>>٩:?Sȥ>
�=��,>ڀ�����Oľ��1?ۤ?�?o��?C�->�݁�������)��<�T?p�?�G<��J ?�f�_e�����&⏾a�����Q{��;Jd�	'��@���]�`ֽz7�=�.?=	y?Jhc?�@?a���;W���g�mꁿ��F���;Yz��OA�=s0��C�$[�3q�2X�q�ʾ���Ȓ����0�0|�?�2?f6���>�P��kؾ���=I>���o�g�+��=c;U�a��>� ����ߵ2��i����4?�]�>wm�>��$?ʰj���I�T�<���>���	�{H>᠐>&Q�>��>gK�!䄾��=�����松����5v>�xc?��K?h�n?�n��*1�t�����!�κ/��c����B>ej>��>�W�>��G:&��Y>���r�s���v��_�	�X�~=̯2?1'�>T��>!P�??{	�l��lx�\�1�i��<30�>�i?�?�>O�>�н�� ���>@�i?�>oߞ>d�����#��{��G��2�>ֽ�>�r?m{>��B��X]��َ��4���c6���=��j?>��ZZ�cg�>�L?_�i��U�<?�>SU��u2 ����T�&�a�>�w?�3�=X.>�E��Z_��B{�ʷ����(?�?�1���2*�܀>w
"?4K�>Q��>z�?)��>��¾I����?j�^?��J?��A?o�>��=_и�o�̽�!)�պ+=�Y�>�[>�1m=W��=t��V`�s����O=п�=Oڼ͏���;a�ȼ��(<EU =��5>�ۿ+�J���׾�U��!�Jr	�����ﶽ뇾>��=붾�J����t�8��%�#�GnU�2b�؍�ʙl�U��?�W�?>���W��hq���9��0���0��>[�o���z�����������ᾶI��H�!��zP���i���e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >ZC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾t1�<��?7�-?��>Ŏr�1�ɿc���~¤<���?0�@m}A?9�(�n�쾙V=���>e�	?��?>BM1��H�J����W�>C<�?���?�gM=��W���	�[e?��<��F���ݻ"�=�=�=�@=I��r�J>�U�>z��TA��5ܽյ4>�م>h"���D�^�މ�<o�]>��ս�@��2Մ?{\��f���/��T���T>��T?�*�>;�=��,?L7H�Y}Ͽ
�\��*a?�0�?���?-�(?+ۿ��ؚ>��ܾ��M?_D6?���>�d&��t���=6�.���}���&V����=D��>!�>��,�Ӌ���O��G�����=�B ��%ſ;��
h��9�=�a<xI8�P��ʽ�Q������Y� I��u��=#��=x�R>:ȉ>LgS>%�^>�aS?G�n?���>T>G��D���>�ھPoͼ�v�Eg��I����*��ԟ��쾛Sپ���/��ֱ�H�ɾ	!=� �=�6R�^���&� �Z�b�P�F���.?�v$>R�ʾ��M���-<bpʾO���
܄�᥽�-̾�1�"n�`͟?��A?������V�Y���W����8�W?�O�ʻ��ꬾ��=.���3�=�$�>���=���� 3��~S�;J.?��%?-_ʾ����>�<>�?����� ?QI
?�Ϝ=���>"�?�P�����z>�C�>0�>��>��=~�������!?Sa?�*��ŝ���y�>jɬ�埧�TH<�[��=�`��u�<�>>�==�F��m�[��8�K��=>�b?�}>��J�q������S]���ֽ�?�?HV�<�[�?~F?����'
$��yU�$��v37>,�V?�Y�?��=6m!�.	��
T���5?=�@?d3>:8)�i��0��޾�� ?�:m?H?��W=��V�������"�Ұ?��x?�U�-�����Y����>�E�>
2�>cK'��̧>!/I?W	�������(�;��ƕ?�@[�?� �=K>-��W=/�>;1�>y!� :��:�ý���7�=���>�ˤ�u�g��m��T ��+A?�G�?K?{��I�����=<���88�?w�?.��5�j<���l��x��3ġ<� �=��z ��M�ɐ7�ޮƾë
�Ō��(GƼ���>}T@��^��>��9���!�ο��zϾ�q�z?/I�>�ƽ�4��yj�fdu���G���H�H+��N�>��>���r���C�{��q;��'����>���	�>#�S�f&��(���5<+�>���>	��>7*��R罾$ř?lc���?οQ���ޝ�o�X?&h�?�n�?q?Ɠ9<�v���{�Յ�O.G?��s?uZ?
q%�>]�.�7�e�j?�Y��AX`���4�gIE�9�T>�3?+M�>ȋ-�p|=�H><��>�0>D(/���ĿW׶��������?ȉ�?j���>-}�?�p+?zd��1���T��l�*��"�|:A?p
2>������!��'=�.ǒ���
?�{0?���,�]�_?*�a�M�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>aH_���u>����:�
i	>���?�~�?Qj?���� ����U>
�}?!$�>��?p�=�a�>�d�=D�"-�k#>E"�=`�>��?��M?&L�>W�=��8��/�N[F��GR�\$�*�C�_�>��a?��L?�Jb>���^2��!��tͽ�c1��Q�W@���,�@�߽�'5>'�=>}>��D��Ӿ��(?���JFԿ]c����}�f?n�(>%�?D⾭ꏾ���=8T?`��=u�,�+o���s���3��"B�?���?�! ?�׾�P�����=���>Cߣ>�_�W��n��w�7>��F?�k��%0��� P��ҍ>�%�?��@�?��L���?j����f���:~�zV��\�K6�=^#;?��ܾ�.e>s�?B�=�����tz��L�>���?��?֗?c9e?��k�&C@��3t=��>�am?OX	?X�"�@�׾��C>��	?��}����Gg?u�	@��@f-Y?e����Ϳ���ȴ�Hھ؊>��F>j�e>�ZB�n����T�=�L=Tʔ<h	>th�>�N|>�JZ>@�B>� >�8>�m������堿xe��o�F���	�@��05����t�w�'������ �¾Yz������2ս��A������d��g�=� T?�U?�j?�?=�dC;>Zv����<�$���-=:�b>8�5?�7I?�+?�F�=�՝�>h���~��ݣ��w��>�� > p�>���>��>E=�+L>��,>�Y�>�
#>��.=��ػ9�8ّ>k��>��>_¶>�C<>��>Fϴ��1��k�h��
w�s̽1�?���R�J��1���9��Ӧ���h�=Hb.?|>���?пf����2H?%���z)���+���>|�0?�cW?�>��v�T�3:><����j�8`>�+ �zl���)��%Q>vl?Q�f>yu>�3�_e8�`�P��{���h|>�26?�綾(B9�h�u�O�H�daݾ=JM>Fž>��C��k�����,��vi�O�{=Ix:?�?x8��Mⰾq�u��B��SR>-9\>@W=�j�=<WM>dfc�^�ƽ�H��k.=���=��^>�e?�,>1�=+��>^����P���>�B>�,>T@?�@%?�D��y��*���.�l%w>�v�>~:�>}�>��J�s�=�e�>�Cb>���}i��4F��?��V>X�~���_�$t�#�z=�㗽�T�=I@�=�� �w�<�;e&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ0x�>�d�QY��-��<�u��"=ԁ�>�BH?X����P�/�=�dn
?��?���׬����ȿVv���>��?�?��m��C���@���>U��?nfY?��i>�.۾=oZ����>�@?x�Q?��>39��B'���?ڶ?���? �H>��?�s?�m�>��w��V/��1��I����S=d;Y;�V�>�T>V���'cF��ӓ��f����j������a>�$=�$�>���C;��B��=8ً��*��!rf�᰷>�q>N�I>Zb�>�� ?CS�>,��>��=l����Ԁ�����ضO?N��?c�!��*��0^��M�<�{��N2�>��a?�C1>����mj5>F=@?+��?��Z?�y�>�D���᝿A�ȿ�<ھ9��=W�e>�&�>���>�F���=z��VC�� �>�ʢ>꽄1������=�	�>�D?t�?h%�=X&?�??l�/>�נ>�H� :��P
L����>�Ĺ>�H?]�}?R?2�;��C�󄕿����b�b�{>��}?�?�L�>����⟿c�:<X������Q�?j0k?��J�?8�z?U�%?43?_�#>	����}AK�wȌ>R�!?$�Z�A�9N&��
~?cP?���>r2��c�ս�8ּ����|��k ?�(\?�@&?���,a���¾b�<��"�;�U�w^�;�D���>M�>%���9��=>�=XNm�D6��Bg<7i�=��>��=�+7��}���?,?AdG�Cꃾ�ؘ=��r�yD��>ucL> �����^?�C=�,�{�����x���U�)��?	��?�k�?轴��h��=?��?G?.�>	G��Ix޾����]w��x�@u��>���>�ol����/���?����F��1�Ž��$� ��>^(�>�C?g1?#�L>@5�>~����&�l����O�\�����6���,��j�S椾�k3�����ӿ��}j����>�ל��c�>�
?�dy>h"�>@D�>�ၼX|�>�P\>-�>|��>��N>Dg%>�b�=}��<��ƽ�KR?����#�'���辿���f3B?�qd?S1�>zi�<��������?���?Ts�?=v>	h��,+��n?�>�>H��Xq
?lT:=�8�P;�<V��~��!3���1��>E׽� :��M�Dnf�vj
?�/?�����̾�;׽��N�f6�<���?+W6?�@K�5�M�3�x�(4P��j����<!䜾������4s�-(���� v���]��r=TN<?�0�?!�6�YH�xڙ�1쌿��:�~3�>Ik�>QkM>��?�O<=VE�q�a�
En�{>�&����1�>�ă?��J>hvb?�6?�%E?�0X?a��>��>6��X?�w��>]�=��(=�!=?4?��b?	8?�<?fk>�a�_t�@���7 ??\?��?�u$?�*7?h�V�|Q7�]�r�~�>�>.,:=}��=�c������#9ؽ"m?>:�?I��D9����2�j>��5?���>��>� ��띃�0�=�*�>��?Wd�>�8 �Yur�o�����>��?�L���=?�*>���=҂��ֺ�j�=�]Ƽ�0�=��K�9H7�"�<u�=�9�=~治�X����j;�8gT�<���>5�?7�>=�>91��� ����퓱=w"Y>vDR>�>�ؾE���B'����g���x>}o�?em�?fGi=���=0��=r\���6�����/ｾFs�<��?i(#?<GT?���?��=?<r#?��>J�*C���c���H����?x!,?��>�����ʾ��׉3�؝?k[?�<a����;)�ې¾�Խɱ>�[/�i/~����=D��셻���R��5��?뿝?\A�U�6��x�ڿ���[��}�C?"�>Y�>��>R�)�~�g�q%��1;>���>iR?�#�>��O?�<{?Ŧ[?hT>`�8�h1���ә��E3���!>@?���?�?ay?�t�>J�>l�)�&ྞT����� ������
W=�Z>i��>!)�>_�>���=yȽ�Z��f�>�a�={�b>��>?��>��>^�w>�M�<�^F?�m�>}Ǿ��)I��Vt������$�a?ꓕ?��??7�D=Rl���C��V۾1d�>��?���?��#?<����]�=u���l���g%�|B�>��>iV�>�f�=��9�
>�^�>]��>Yp,��l�8�.�gȌ�%,
?�pN?]>�
��aP�����~o}��/=��V<Y@��^ZѾ�3=��_�շ⽗����ӽ�b��Z�[���Ⱥ��HB���?@�;>��=�v>�>k>�=����?<>�t0=��|򽩕�=�Τ���q=w���[
_;#�\=���=fd�=ъ˾X�}?<I?��+?��C?��y>�;>��3�C��>c����??�V>��P�#���d�;�!���!��\�ؾx׾;�c��ǟ��I>�eI���>b83>�M�=bY�<��=s=ﾎ=OVQ��=| �=�K�=�`�=���=�>V>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�48>E&>��R�!q1�!�\��$c��Z�	�!?�;�3�̾-��>o�=D�߾��ƾZ,=w�5>�Qc=o�T�[����=��z�1N<=�l=%ى>��C>͚�=F3��灶=��J=���=�O>qڃ�S%6�,���3=ś�=l	b>}�%>��>��?`a0?�Wd?�6�>�n��Ͼ�?��5J�>#�=�E�>߅=crB>y��>e�7?εD?��K?���>���=j�> �>Ӛ,�E�m�l徟̧�@��<{��?@Ά?�Ѹ>��Q<R�A�ڠ��g>��/Ž�v?�R1?�k?c�>Q
������,��M>i�|�=�hx>�k����N���>��A��i4�E>q��>���>tN�>��a>���=@C>��>9׋<���=E�#>����V=G�,i��@W=���=��=mv�>�p�<f����N
���]�5���=T"=���=���>:>Ϭ�>g��=(���A/>����k�L�W��=�F���+B��4d�cI~�/�lV6���B>*<X>y��4����?R�Y>n?>���?�@u?�> ���վ�Q��2De��US�θ=Y�>N�<��z;��Z`���M��{Ҿ���>Oߎ>��>ںl>�,�d#?���w=�#b5�?�>�{��o��*��9q�%@������]i�E#Һ�D?}F��I��=9"~?��I?7�?!��>p���ؾf;0>LH���=D�~)q��f����?B'?���>�쾹�D�R����'��
��>G�e��W�a���<�Rs�=�Ǿ��>@�����Ǿ��=����幕�TQZ����ɼ�>%�Z?yݤ?(�6�"����>^��;��5���t3?Dwl?=��>cL�>��?�Ľ����Y���E�<�m?�R�?��?��T>0�O=F�#��-�>�X�>?�?*Ґ?��?�B���>'�����>J�R��>>�-[>�D>V�
>~�
?�>�>i��>�%ͽ�h�k��x� �u�;���K=���=e��>�D?>��|>-�D>%�>uU�=m�}>�5>#l,>>��>�dx>n���G�߾��B?z�=��>��<?�۪>��(>Z��<�Y�X�J���;ν�yн�G��ؽՊ��l�=�T�;�5 ?H:ɿt�??k>�].��} ?�[�R��={��=��T>��#��8�>�����]>�$7>�Ȃ>ܺ�=#x�>M/>IUԾ��>��	���z�@��/Q�'�Ͼ�r>ߛ���'�Z	�+��SA�����V��^�i�[:��.S>����<^��?��޺h�^*�͙�m}?ya�>4e6?���V䒽N�>3��>��>����7��ݍ�����?^��?�;c>��>D�W?)�?��1�3��uZ��u�n(A�-e�O�`�፿����
�u��(�_?�x?-yA?jS�<%:z>T��?��%�Pӏ��)�>�/�*';��?<=z+�>*��e�`���Ӿ~�þ�7��HF>��o?7%�?jY?6TV�����j >��:?ko%?��x?�v8?�uH?0�ὔ�?�)>��?ԫ�>P�9?��6?.+?W�1>���=Si�m�8<Z���`���V߽������2��<���<��<��:��,�=$�z=l��<�þ�r}�<�VԽ�͈���=�y>].�=?ק>HF_?6��>�qv>m�6?�&��8�`g��T2?�f�=��~��ي��
��zA�o�>�o?yƫ?�X?�K>��Q���<���'>�w�>�r2>X�O>�c�>�z۽n�a�)=�3>�$>�è=��{�A�v�5`�F���/�=�6>D��>�|>�����'>�T���`z��d>Z!R��T����R�(�G�L�1�V�v��m�>��K?/?���=4�D��\Lf�')?{]<?�eM?��?er�=��۾��9���J�^��q��>`�<P��¼��,����:�vu�:�/t>Qʞ����j��=��r��vX�%%g�-{ �����>��/��d�=PU���^ς��>o>Jۂ>�HܾUD���� ����H?	��;dv��ϰ��ݞ���>���=x��>M�������9�����=�=W1?���>U��=���p(��B��:�>�OE?�W_?�j�?�"��s��B�W����e���ȼ��?;s�>7h?"B>��=����=���d�/G���>��>B����G��:���)����$���>�8?�>�?��R?��
?�`?y*?}E?E*�>��������A&?r��?v�=��Խ6�T�� 9��F� �>�)?%�B�ǻ�>L�?�?�&?ĄQ?B�?#�>r� �)C@���>DW�>��W�$a����_>��J?嘳>�;Y?�Ӄ?��=>�5��梾�橽�9�=>��2?k4#?R�?��>m�>9斾6�c=a�>�5]?hxz?2[}?R�=�?tmu>���>E��=%�>2�>�6?�]Y?,�l?�O3?|e�>���;���`����ؼ�x =!�>=�}<	��<�2:s#!<O�C����:U�<<�p�=��<B�8<s�v�M吽�����}�>��t>|*��QT0>��ľ򚉾��@>�Ǣ�UF.��e:���=��>��?�(�>��#��ђ=iּ>�>�>��	(?0�?l-?�/n;Ղb���ھXVK�;��>�QA?���==�l�\s����u���h=n?�}^?�X��T��b�b?�(^?����<���þ�d���H'P?�y
?e
E��x�>��~?�q?�#�>��f��n�0ۜ�OTa���h����=h؜>׼�">d��=�>�7?b��>O�`>�p�=x_ܾtw����8�?�?��?u�?�F+>�n�,࿮%��|��{`?1�?�5���i.?6�<�㾭`��BU����Ͼ�Ŭ�����;k�_��2
3�>ⅾ���m,�<?�y?-�c?�mV?����8l�^+d�H��� M��������&C���G�ne<�ndo��c�����m���c�=�Ӿ�y���?g�a?�����3>?ݿY����UY� ؞=�28��|��
p�>��8>1�>y�Ϻ��`����������&?U��>�<�>(B?u�6�d!������F^־0G\=TTX>ϙ]>��>!�����4�!�00���]/�QP"�8v>�xc?U�K?��n?�k�+1�������!��/��c����B>�o>躉>�W�����9&��X>���r����w��2�	�.�~=�2?�*�>���>O�?g?�z	�l��2ox�3�1�B��<�-�>F i?�@�>��>*н�� �b2�>?m?���>%�>F����!�mw�6������>tE�>\��>`f>�
,���Z�����y��HQ8�+
>��i?�9��N�V��B�>��S?�R4<�,��K�>c�����&�C����-�=Ih?�J�=�l<>����ح�$Zy�˯��%1#?�.?3���m+�Y��>��!?��>s]�>�r�?�4�> Ҽ�<n<�?�"^?�>L?��D?�Q�>�y�<Oý{c̽��0��	=p�>`j>�6�=�F�=�"��W��#�'�=�$�=Q�4�'��o�<����;L��<��/>@῏EM�����r���辻�ؾٽ%�d������nI�|�������������� �������I���Ѿ�P��P��?
Y�?�ǯ<��;�6�68���D��r>H↾�)�IhD��,� {z���꾶����R.���f��n���^���'?7����ǿL����PܾU ?� ?��y?�����"��8�}=!>���<	������N���H�ο�����_?J��>f���X��u��>:��>$�X>�~q>�)��#瞾�$�<P�?-?
��>"�r�0xɿ����\K�<���?%�@`}A?_�(�$���U="��>�	?�?>I1�gH�v����X�><�?���?��M=��W�"�	�{}e?��<D�F�A?޻) �=�?�=]O=j����J>�T�>,��c^A��Lܽ �4>�څ>V�"����Fy^��\�<D�]>��սGO��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=}��cǿ��%�%&��fB=қo=�<=��6��?!�q�h�)���/�o�^6�����=��=WF>A�>�>b�+>�hM?��p?���>�i>$9�����M���B����ci(��4n�k �gܩ�����T"�%
�v3�H���6׾!=�W�=7R�h���7� �h�b�W�F���.?$w$>v�ʾ��M�\�-<�pʾr���݄��ॽ�-̾�1�
"n�e͟?��A?������V�D���W�����O�W?P�ʻ��ꬾB��=����Ơ=$%�>�=~�⾺ 3��~S��J-?�;3?���n���T>�>���X�=Z�:?��>�d=��
?��<?��གྷ���yCS>���=�k]>���>���=���Lvؽl{?��K?�����3w��)�>ۧ����c�6�W>=��㟣;j>�H�=��B�@=������`?�p�>��4�ZD2�ʠԾ��ѽ�y��L��?�x/?�	�>��8?F�B?Bji=���߂n��
2�aO?��?�J�=�.�=*���@���g0?gK=?���>�X��]���Ț��s?�?�?9�?K�=�����G��0��C?fb�?�O�e�����3�d�`�l>��>#?������>�>?T��=�������V�����?�	@��?~�ؼ���E�=׆?�e�>����������&��n@�=m9�>������P���'��h�I0?�o?S��>�˒����+��=/���NA�?�ˑ?�v��˾�=F���v�X$�\���T�=jBѽ �༪G���j2�Q�Ծ�B�N\��y:��:�>~i@�<�m�>R ��}�鿮>ʿZt����� �#�:�>B�^>��H��nþX�|����d�:���;�tJ���>�	>Z����D����p��1=���0��>�|����{>
sP�l0��޴�������>-^�>̌>�o��>��R��?�` ��ο�✿v�
�Y�W?vZ�?��?c?}>=��P�mr����f�E?��u?}X?�?E�9�,�9с��Hn?�p��y�7�R�p�R���=fX?1�>*�����>5�Y�{��>��=E�=��^��������Ģ?/�?��ɾ[p�>_�?d5?Y�����@��ڊY�9u7���?a�>��1���.��%
���Y���>�D?�t�^3?�\�_?+�a�M�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?ӵ�� #�f6%?�>d����8Ǿ��<���>�(�>*N>lH_���u>����:�	i	>���?�~�?Qj?���� ����U>	�}?֜�>N.�?�>Fפ>ق�=�zܾ���<
��>i-l=q1%���%?�K?�>Fa>���Ir)���,�n���QD�Qqy>��I?+?��>~���L�����JF�>t��Ʀʽ�
�Q5M��rM����>��X>Ы>�|��V�M_ ?R��ەؿ�Y��Y�/���0?��v>:?h���x�i� J���b?"�>���>⳿r���L����?N��?�K?�dҾ
��W�>?;�>ωz>̈́����ؽ�Ì��[8>4�=?��%�䦊��l��"�>��?�b@p��?oi�@c?`�ڸ����\��{ľ}B����<�F;?�EǾԲ*>k��>�=��{�$����O����>�ݱ?Gb�?���>��q?OSy�D1J��a�:'`>"�g?F?�=>��� ��>�=?,i������g쾂�e?�e@tg@�?������׿�Ǡ�PV⾨�׾X*�>g��>1N ?�s�w��p��=֐��/	��S�>�J�>�*�>��W>�Ԋ>V�=���=����c��������<JK�br�<g�ק��� &�m���h�����r�ƾ@~�	�j��%�B�D��?�������y�<^�7?!``?�0l?83�>I�#=�]�=���-���w���=��?>)�1?;xZ?��3?EM=bK��Awo�zn��+�������>�9:>\�>��?*��>�A�<�K>�� >��>g	(>���<��'=!�m<��N>u��>f�?\~�>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?e�f>�u>t�3�:e8�;�P�J|���i|>�36?L鶾+D9���u���H�$cݾ�HM>)ž>xD��k�i������ui�u�{=Qx:?��?<7��4ⰾ��u��B��)QR>q:\>Y=�i�=XM>Qbc�?�ƽuH�j.=��=!�^>,�?��7>&đ=Z4�>�����W�xS�>�J>s+>�Y=?`3'?��ż�T���!~��%��p>�c�>��>K�>�jN��Ű=B��>��\>Β＂�|�F����=���V>y���]�\���m�ƻZ=$���E�=�0�=�����K>�F�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�[�>n��R����և���w���=y�>�L?��׾DH��Da���?8�?��������ſ�uz�XB�>�G�?L��?Aed��ט�|A�L��>|)�?3�W?�n\>��Ͼ]N[�|`>��B?�P?BԮ>�c�4.7��z?��?L��?�I>���?Ϟs?�k�>+x��Z/��6��ؖ��pq=��Z;d�>oW>�����gF��ד�Oh��,�j�c��j�a>�$=��>]E��3��<�=��]I��+�f�Q��>�-q>p�I>�W�>d� ?a�>@��>�}=+n������b�����K?���?����0n��8�<=�=t�^��(?�<4?d�[��Ͼ�ߨ>�\?��?��Z?�P�>w���0���⿿����O�<
�K>�$�>BQ�>��W:K>�Ծ�*D�O�> ��>�+��/Uھ�U���Ĝ��M�>Z!?ē�>Cn�=�!?�q!?pl<'g`>��c�9ʌ�a�]��{�>z�>��?7\?p�>���	eJ��2���'���t�A��=@�?w�#?�W�>Y���C���;���)">P����0�?7�?�����>j��?��O?$?�d=s.�=ӖԾ��W<h��>s�!?/ �6�A�QL&�γ��w?f?���>듒��Bս�)Լc���L����?H)\?�J&?%��a���¾��<4�$�=�P��J�;�B�V�>�>�~�� �=�F>F��=�Qm��,6���l<���=���>��=�]7�齎�?iB?2���g��S�_=�	u���C�ִ>�ɿ>t�]��CB?�<�>�>�;Ǽ��Ƙ���O�A8�?���?w$�?B�����V���??�˅?��> ��>������ƾxi�%ӽ������\�
=�/�>��=��D��������W�����=%��|��>�b�>'K?��?�]?>�ԭ>����]�$��f�4����^�
����9��A/�Uu��B��Kr �m]Ѽ����ѯz�:��> �g�>�>�?��V>�w~>���>
%E�Z��>9`>l�|>rB�>J�g>bI>�>�M�;o*ɽLR?����ٿ'�-�込���G1B?�od?3�>��h���������?���?�q�?�4v>h�L-+��n?�A�>���p
?#X:=g:�TL�<�U�� ���B��?&����>�K׽� :��M��mf�/k
?�-?�􍼡�̾{H׽Wfz�Y1�UB}?B^A?Y�H���G�l�l�`i��O�lf=`Os�*�6e&��_�:����ŕ�~�w�@a&�i:d�,?�͗?D�:��+�䱾�Տ��OB�z��>fu?$��>��>��=�J0�q�a��1\�-V-�t����z?�ז?&v�>�E?ԭ*?�$;?��T?ԆB>4��>
���l�>�м�o�>U� ?;�$?ʇ?A�3?�?�?#�>^J��O�������n��>��?x!?eU	?���>�ž�.����#C�P"��c�<z��=��E=y#-�gَ�������>�?�����9�~���d>�k6?�R�>���>���s���s�<?��>�F
?�>�{��hr����i��>툃?�� �f�
=�g'>��=:P��8B���=���}��=�~�wZ�$N+<ܵ�=��=B�F;�ڻ��N;L�L<���<}�
?^t?��[>KU>������ %���">Y�>[c�>��>�Ⱦ�f��s���P�d�"i�>Zŋ?�1�?�ܺ=^F�=�q7>U�o��AѾf�������p��=�g�>��?�^?�ܑ?�%?��G?5J>������>����è�|j ?g",?���>��� �ʾ,�ψ3���?�[?6a���n@)���¾��Խ�>z]/�S0~�Z��D���� ���y��m��?���?,A�G�6�p辯���`���C?�!�>�K�>��>��)�c�g��$�W;;>���>QR?� �>\�O?C;{?�[?SjT>X�8�N/���љ��3���!>�@?���?^�?fy?w�>��>�)��ྫU������!����JW=>Z>ߕ�>�(�>��>���=�Ƚ�b��8�>�-\�=�b>���>���>=�>w>�v�<1EN?�N�>��ݾx���v��bޚ���ƽ�:z?}��?;�?��=��
�n�S�C~�'�>=S�?�I�?��??T�M�l�'>����㶾������a>���>���>��>C�5=/@P>=��>1�>��W��C�!2.��-�3X!?#�M?���<�Eſ��r���\�������m<�f���h�ޒ���ud���=���������o�I��w��L������6䠾nX�����>�Me=(��=�B�=Q��<[��=K�]=4R�<�W=�Pj�=��<R�3��	�:����
w:%e�<�l=F����|¾�;z?�D?gw ?�(A?��W>��*>÷����>��U�ۘ?�"W>�	<�tɷ��K�η��E-��+�ξ([оi8`�@���R�>�b����>��1>���=]�<t:>�i�=��C=��*�Jtc=�J�=;2�=��=xL�=�=��=�6w?X�������4Q��Z罤�:?�8�>p{�=��ƾp@?�>>�2������zb��-?���?�T�??�?@ti��d�>L���㎽�q�=Q����=2>q��=w�2�U��>��J>���K��B����4�?��@��??�ዿТϿ9a/>�A>X�8>��E��`1��^=��n{�?xB�.�#?ձ5�Q�ξw֙>�9>9<߾գ¾ꐍ=2,>d�=YQ̽�A[�)�6=���[&=��=&�>(=F>���=����)��=K�<ʟ�=ѣx>�lԼ�z�v[���
�=�~�=�a>��%>T�>K�?U1?��d?���> 5��]�°���>�0��4��>���=a��=Ā�>h�2?�]Q?udJ?��>$��=W�>h��>��5��a���得g��r3�h�?�A�?O��>nd�=V����02�[;	<݅?�9?�� ?gO�>�U����:Y&���.�������0�+=�mr��RU�y����m�>����=�p�>���>��>MTy>��9>��N>x�>�>9�<�p�=3ꌻd��<����=������<�użO���6}&���+������;竆;�]<R��;��	>��>O��=��>�V�=^þ��%>���O�B�Bڐ�zN���+J�!�g��{�A@5���*�ިP>�h]>޴!�,���E�>��z>��t>�"�?I�d?���=}%ڽh�ܾ�1������
+��=��=c��&�N�R���Q��̾���>;Ƹ>�->��2>_f3�� C�
�o=��޾D��o�y>���ig��v}� &e�e릿i[��\�I��=5�C?'���� �=�~?@qh?���?���>>D������%�<6��F�5=*���#���½�v?iN?�?�|��D�̾�o����>2�H���O��Õ���0�������C�>D���о&13��l��:폿�^B��
r�!��>p�O?��?�bb�?`��MO�`��nׅ��^?Ύg?t*�>Jp?�`?�����u�Ta�����=]�n?��?kE�?��
>;��=DJ��7M�><	?6��?���?j�r?�?�T)�>U��;J� >��;w�=�i>�Х=6��=�?�W	?!�	?�-��G
����ﾜQ[�,M�<�=�O�>��>R@q>>=�=f�c=�=l�Y>��>��>cd>���>��>,�޾��)��N?@�~>[~e>+J`?��=�ලA����B=~Ե=a�������H>ʇ�=���x�� ��P�BI�>������?�v�>q	���.%?+Ce��`=��>��>/o�,��>Xi:>��N>�k~>:v�>�a^>[�>8��>�?Ӿ��>���Ne!��.C�W�R���ѾL�z>����� &�����g���@I�Gq���k�E
j��.���:=� ~�<+G�?#����k���)�����ԕ?�[�>�6?Ҍ�5����>���>͍>�G�������ƍ��e���?���?�d�>3�>�3?? ?�o<X����V�mjW���!��?��)0v�
���Uk��R&�&���i?y�k?�0?N�=��b>O�[?Ǘ�p6#����>S� ��zI�߷�=���>k)q������f�����^=l����>_X�?�Ut?G?�D4��2��]�<>5g�>�->� s?���>Y?�V�^_)?��>��>�>r.?�?�V)?���>;�B>%�	��<~0��������ٽi�5�1�#��G>1>e>���=�_�=�����]F���=�)>�t�<���=<��=P�B�G��<�w�>h ^?���>Ĉ>��9?Y'�Gy8�r����7.?&W<���f����Ϧ��F��{��=@�k?���?N�X?7i>��?�HD���>�ӌ>3 5>�Y>��>�����>�p�=��>��">J��=�i��m���vЎ����<ٯ>���>%5|>v��~�'>�{��6z�ԣd>
�Q��ʺ��T���G���1�@�v��V�>\�K?��?.��=�\�p&��If�'/)?^<?�OM?��?R�=��۾��9���J��K�k�>�z�<������L"����:���:$�s>�1��ћ����>$ϫ�4\���΁��c.�A6����J�	�=�i�C����1����=&�:>�A>Y�㾧�%�4���4E���eK?�R=Nh��򦺇�Ѿ�k�>u�>���>d0�=��D�r39��j>������ƨ>џ�=��]=4�	���1�����>�>_QE?�V_?�j�?�!��s�k�B����9c��fȼ>�?�x�>�g?�B>M�=Z�����R�d��G���>��>���v�G��<��-0��(�$���>?9?A�>@�?��R?��
?8�`?*?�D?�%�>��������?&?���?�ل=��Խ[T��9�ZF�~
�>�p)?�B��ȗ>��?$�?l�&?�Q?��?M�>ݟ ��F@��w�>"K�>��W�FU���G`>c�J?���>�$Y?�҃?]�=>�z5�/ޢ�}��4�=�>E�2?TC#?q�?	Ը>�'�>����F��=B'�>�g?Nc~?��n?\\�=�� ?Z46>�V�>�B=�z�>F��>24?�|G?�o?%OK?&"�>З�;�[���K��+���H�E�]J7<4w�<I�\=�)��H\;�;⮼�P;<�<���@G�l�`����c�1�-YǼi��;�_�>��s>���~�0>�ľ#\��;�@>�����S���֊�z:���=���>��?W��>7K#���=���>�;�>���N2(?��?�?X<);7�b�w�ھ��K�&�>7B?#��=��l�y�����u���g=��m?��^?zW�����{j?9�Z?�R��4��Um���yؾ�V?��>v��<��?5�?Q�b?G~?�}��E��e���YJ�d}Z�.�o=��>k�־��T��R>;}?B�= {�>�ξ�mG���js��Ɲ��v?$�?�f�?/�?Z���2n��濫��ì���r?X�?�"˾"=?FP�=��������]��z@�8M��5ǁ�fR��jY��"]��U���Zb���l7?�ls?�A?�[J?F��u�]=Q��qo��CA�k���D��NkG�� B��NB�3p��:i!�|\�w��4$>`G����i��?�?�9C?\�1��)?o%����|�;��=\��{2��&>�Թ<�E�=��=����c˖�B��H�!?n�>��>�#$?|QR�B�1�q� ��G.��w��	�L=�&\>�UZ>���>2����~��D����¾���p?��7v>�xc?�K?A�n?Dn�Q+1�����ә!��/�hc��Q�B>dl>)��>��W�Ϛ��9&��Y>���r����Iw��%�	�å~=u�2?K)�>³�>P�?s?K{	�Gk���kx�݇1����<�0�>G i?3A�>��>Kнu� ���>��l?\V�>�>�?���W!���{���ʽ��>m�>Pa�>Žo>��,��>\��g���y����8�U��=�h?�o��s�`���>��Q?Aw:�L<���>|,w��!����`'��>�?��=a_;>��ž�(���{��	��k)?�N?�����*�a�>q�!?��>AM�>
�?zP�> ¾yz��*?i�^?�FJ?E�@?67�>�3#=�l��+�Ƚ��&�)�.=+�>�X>�m=xx�=���R�[����oF=_��=KbԼ޹��k;�;Q�ȼ�+L<sw�<��3>gF޿�xK�o�þ��bC���������D��K��8�ӽl~������ ���f���j�q���%�� ��)������?��?�c$�ç*��������^���Ձ>���wM(�Wɋ�Hν�;�x�־l���A,�'Y��Xt���n�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��o��>ݥ�>�X>�Hq>����螾�1�<��?7�-?��>r�1�ɿc���r¤<���?0�@�|A?�(�Z����V= �>�]	?ĩ@>9�1�m4��������>��?(ڊ?>�G="�W�ݓ��Ze?N�<�F�j:Ի��=U�=�d=���Z�J>(��>T�/aA�YRٽ�.6>U2�>]���b�sX^��a�< �\>;׽<G��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=3����Ŀ�<��� �dA<�;��>��%�������K�Qb����[��]�4Y�=8>��K>�(�>؁8>�A>�WT?9Hq?׃�>�#.>��6��量e�d����}��A
�f�g�SE����Kؾ��ܾ��'��W#���F!=�+�=�6R�>���m� �P�b�j�F� �.?�t$>�ʾ��M��-<Soʾƿ��0ڄ�#㥽�-̾6�1�4"n�b͟?��A?����^�V�j��U����%�W?P����ꬾ���=<���!�=�$�>Ɗ�=0��� 3��~S�.q2?K�?k� �ai��d�`>�S���5=�,?�+?�a���s�>�?󐆾�F��	>��x>Ő�>�2?
�`>8x������*?��Y?]<�g���æ�>7���L����罩ڵ�K9)�Cm����<�pڻ垾�t׽�Z�[�;���X?���>%e3��� �㋉�e@T����</�|?��?	�>q�m?tg<?X>]����!S��������=w?_?}m?�>����N�ξm���Q3?hW?w�b>5���) �b;�V\��9?"4e?�s?����ct�9�����#�,?��v?�<[���۫�BS�5��>#�>c.�>�6��s�>�x??�.�;����㿿64���?�@>%�?��<��'���=M� ?�m�>�_G�N�Ǿ

��;W����0=l��>�b���7t��F�9�8�լ7?x7�?�.�>�j��K�w��=E˛��d�?N�?Xܯ��}�<~�m������U�;F��=y�M��[��ʻ7��ɾ����a��Jۼ�ʈ>n�@����>&�9�H��e�ο����b�ξ��f�Q:?5��>Ւ�Y}��7�n��'v�kZF��G�o�}�tZ�>A�>=���������{��n;��䢼��>8���>�S�pY��!̟��3<6��>��>Kʆ>L̮�����z��? *��>?ο	��������X?"d�?�t�?S�?�9;<��v��{����$G?��s?�)Z?�R#���\���7�%�j?_���U`�َ4�&HE��U>�"3?�B�>�-���|=>m��>;f>$/�Z�ĿNٶ�����W��?ω�?�o����>V��?�s+?Wi��7��[����*�)�,�v<A?-2>ߌ���!�<0=�)Ғ�}�
?�}0?�{�d.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�0�>��?��=m(�>�=����>�8��O$>:�=J?>�D�?��M?"��>��=�f6�A�.��kF�:�Q��I�(�C��Ň>8�a?rL?�c>/��[�*�Z!���˽x81�Z�輦�?�da/�
ཊ�4>�*>>k�>u*C���Ѿ��?Mp�9�ؿ j��!p'��54?.��>�?����t�����;_?Oz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>A�Խ����\�����7>1�B?Y��D��u�o�y�>���?
�@�ծ?ji��	?~��P���`~�A���7�٩�=#�7?s(�8�z>s��>���=�pv������s����>�B�?�z�?	��>/�l?O}o�1�B�Û1=N�>Μk?ou?B�k�W�򾽵B>	�?��@����K��f?��
@+u@��^?�좿�@׿�}�������ľ�>V?>A��>j1!� 4=�A��E��껚�r>��>���>��>��>x�A>��L>n�~����=����<��$�^���(��/�gc��.n!�M�f��W��ʖ�1o����;��ӽ����1(�Kge�]��?Ӻ=�M?�M? �l?%�>|a��y^>h��5r}���5�H?J=t�>��/?��K?��-?�֔=����_������J���͑�a�>��T>]��>��>��>Yw��uf>YC>�(t>�Z>ǀ�;n��;DZ=��T>x��>q��>�>�C<>��>Eϴ��1��j�h��
w�x̽1�?����S�J��1���9��Ѧ���h�=Hb.?|>���?пf����2H?%���y)��+���>|�0?�cW?�>"����T�/:>@����j�5`>�+ �{l���)��%Q>ul?��f>(u>��3�pe8���P��}��*c|>�36?궾�E9���u��H��_ݾ~NM>�Ǿ>��C�Xm��������vi�>�{=�w:?��?�*��#㰾��u��A��yLR>97\>pH=�\�=�SM>�ic�L�ƽ�H��n.=��=�^>��?a�3>�~�=���>P��I�O����>��D>@ ->n�>?��'?ڧ,��K���o!��_>3��>�Ą>�Y�=��I�1}�=aL�>I�Z>?4;������~$@��kT>my���^���Q���z=}������=)	U=���g�F��]0=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�i�>Nq�Z������u�Z�#=���>h7H?�U��L�O�	>��v
??-`򾭩����ȿ�zv�p��>��?��?F�m��?��x@��{�>���?QfY?Twi>ne۾�NZ����>��@?rR?O#�>�7�ٓ'���?�ݶ?��?�I>���?̞s?k�>�)x�{Z/�-6�������p=އ[;ye�>W>����4gF��ד��h���j���a�a>՗$=��>C�$4��J7�=�񋽚H��)�f�ϥ�>�,q>��I>�W�>�� ?�a�>���>qs=yo���ှ�����3K?!�?޺ �x�]����=(�ؾ� ?���>GJk� ₾<��>�Q?���?�L�?���>��@�
ۉ�(���ҧǾ*��<p4^>�#?��%?W|,�Y�5>�k��w>^�h�Z>//o>�m�����)$��.�`>.��>^y!?�1?��l=*?wI*?n>��>z+�W���K�����>#3�>�?.a{?1�?�&��C)�F�������)L��*>>�\}?�?�_>��j������`6�@�����%9�?A�X?�w)>�PE?���?1~;?10|?�X�>���vL
�����¼#>|�!?n��d�A��N&�ݓ�`n?<T?,��>���c�սx�Ҽi��ڄ��1�?�'\?l#&?8���a��þft�<�p"���K����;�?I�ک>>�>�����=��>V��=`Hm� H6�,Tb<���=N<�>O��=P7�䂎�?.?��E<�䟾\��=ڗc�pEG�<�{>?�T>�6��O H?�?���p����xӡ��b��N�?J��?x�?�g��rc��9?�n�?Z5?+��>
3��Õƾ!]��T��J ��o #��c�=ܛ�>ĳB����������-����뽇�Ž�?�И>�H?	Q?.�#>�C�>�[��r�����}�nQ��o�˴H��v2�n>�	��@<����<�ū�^�H�>tش�!��>�a?�G�>h-j>:5�>���=CQ�>8	{>��>6F�>){3>��R=���=������R��KR?U����'�ҷ辥���!3B?�qd?�1�>�i�*��������?���?Ws�?�=v>�~h�-+�>n?>�>W��@q
?#U:=o0�n>�<&V�����2��1����>�F׽!:��M��mf��j
?�/?D����̾
>׽QЅ��DĽ�C�?I K?�K<�n2�2�Z�N<c�5<�H��������d��R(���_�W���cǋ�#m���A���=�+?	�?��:��� :|�8��r*d����>��>���>h��>5��=h�N�ݿ7�`{�7m �#&�#?���?��>^SH?��?�/?h�?9��=ք�>"�<�_��>����J9�>�N�>�_?w�3?��[?��$?;�?:G�>�Y*��
��o��T?[��>@-?�&?f�?�⧾à}=�o�;c�<J��e�2�ÿ<�Q
��/"�mW)>�>�)�>|]?�X
�E�5�/����s>#5?�P�>��>�~��o�{��e$=���>�=?r{�>M���φs��
��U�>��?Kq	��W=G�,>���=j+��<؄���=�qμ�׎=�֋���C��ʃ<^��=Zx�=�}y���%�;kv���wS�<�?x�"?�^>���>��M����~�����=p�H>�`>��=4�Ӿ�6�����V�h���N>4�?W��?��=�>mb�=��~�O�¾�T��-��7n=�?p$?f\?y��?vAA?�v'?j>8S��F��**��*魾��?w!,?*��>�����ʾ��ډ3�ѝ?`[?�<a�j���;)���¾��Խ��>�[/�W/~����&D��텻���D��,��?߿�?�A�:�6��x�Ϳ���[����C?+"�>/Y�>~�>$�)�f�g�x%��1;>��>lR?g0�>��O?�{?1�[?=�U>��8�u!��ǟ��A<�n�!>y @?ݷ�?֎??y?^�>7>�l*�Ƚ߾���-"!��G�З��+�X=\#[>mΒ>���> i�>A��=�ǽ�"��^�>�*�=d4b>YI�>��>x�>�ox>Թ<�W?o�?�j ��vI�����I.Y��z���щ?�4�?%t?\p�>�4��X����j���S�?�ɸ?�6j?�u>}}>z\��k����o��>Mە>Kͻ>t,D>�"	>�b�=���>J�?2@�='?���ƾ���=nm�>��/?�= ÿ��q��O3�m�m����G`���>�F����s�i�$=�C�����S�����1�X���r5��;Z����������D�>���<�x	>�)�=%q�<���<Zyg=�F=�)u=�=���c�<^
���U,�$_s��U�<w�4=%B= ?�������r?u�A?��?z3K?!�(>�|>��:p?�>�/7�g!? 5>\�ս뺥�����@��Z�������َþ��f��[����>�5<�\f�=*SD>�R�=�⸼d��=�l<��r��r>C8>�5[=E�;�=�s�=��;�08>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�-5>�>~P��Z1��ZQ�:hb�Y�Q��� ? �9�nɾ�$�>N@�=Υ�!ľ�B=@�,>y�b=8���e[�o��=�Yv�� I=)�b=��>�YA>E�=bN���N�=1�F=�=�HQ>�|���(Q�ێQ�9�=��=G�[>�&>��>.�?\0?fNd?�I�>�n��Ͼ*/��*E�>�!�=�N�>&��=BTB>㒸>0�7?۰D?��K?���>ܬ�=���>G
�>��,���m�[k�ݹ���{�<Z��?`͆?�Ѹ>��R<ҠA�M���e>�2fŽk?�T1?�j?$�>�U����+Y&���.����C/� +=�mr��RU�����n��㽮�=�p�>���>��>�Ty>�9>��N>��>p�>�7�< p�=v������<L��S��=覑� �<�uż:���V&�"�+�`����Ս;;��]<E��;5v >�F�>ڡ=7q�>�>�[ʾg�:>k����98�:b�1�ľ �6��c�9
��cA0�B� �	�_>���>D䊼w���t�?��>n>���?�n?�K>0ig�م�𼗿�����Jc���>^�>"�Z�Ѹ@�{�[���X�\þ���>�ߎ>c�>��l>s,�O#?�_�w=��,b5���>}������)�:q�@������"i��Һ�D?�F��֝�=v"~?�I?I�?��>����ؾl:0>�H��A�=H��)q�g����?�'?}��>"�u�D�L큾��M����>������I��9���Ye���l�x�p�D�>F���g �GVh�n��-<��@A�%�4�@�>j�d?�ˤ?ڷ�=����zj���8����x�N�>�%�?���>��?�x�>�^#�	��s4��PJ>�˅?ȷ�?��?��>F��=����~��>��?���?>Ѝ?��r?KP1���>�(P<�s<>�����=Y�>�N�=�/�=�d
?�?�?���4����*��эu���
=�_�=��>%�>8qs>�}�=�MB=a�=��>>�4�>��m>�0`>=��>rʅ>��D7���J?-�>n����|q?xZ�>�K6��Zs�@��7����߼��=;�>�HT<�A��,�%���R��!O�غ�>=�ſ�?���>��$�A�.?�ȏ�Х�=��>�=�>�u�Jl�=H��=S N>_�>�/�>J��=�ǒ>=Zk>�FӾM>���od!��,C�	�R��Ѿ�{z>���&����5w��LAI��n��sg��j�6.��T<=�Hʽ<H�?�����k���)�����R�?�[�>�6?�ٌ��	���>���>fǍ>�I��K���Gȍ�h�d�?��?Pnc>$�>	�W?��?��1��P3���Z�m�u���@�B�d���`�������
������_?��x?^tA?��<Xxz>���?P&��J��*H�>Z�.��;��z?=hy�>���h�`�3�Ӿ|�þ����F>3�o?i6�?�y?mCV�O�v�/>ܬ9?˲)?��t?�A,?M=?G.�V!?��4>�	?&�?0H-?H�*?�
?�>���=��9�x=\U��z{���k����˽B��({J=m3=6�����;b��<`[<�q��j,��K���L�y٦<G�/=��g=��=���>?K\?��>A�>i�;?A{$�g/�哦��,?K��<V�������������=a�d?�Ш?�"Z?�e>3jB���7�ê->^ �>�>O�c>�5�>
��/mK��À=#�>�>f�=�a@������������7���9>���>�:|>x��^�'>Wc���7z�-�d>2�Q�RǺ���S��G���1���v�lU�>a�K?��?m��=�M龿3���Ff��*)?}\<?HM?~�?*�=��۾�9���J�7�g�>��<��������"����:�J�:o�s>�+��{�$b>����R޾��n�"�I�2���UL=��z�U=��O�վ����=�9
>z��� � ����#֪�7J?�sj=�f��LU��m��D�>��>;ۮ>�a:���v��@������3�=��>��:>�ߚ�$���{G��5�h>�>TQE??W_?k�?
"��Xs�9�B�z���jc���ȼI�?lx�>&h?�B>���=H�������d��G���>���>e��H�G��;���0��L�$���>X9?�>~�?V�R?|�
?s�`?�*?@E?$'�>!�������A&?+��?�=��Խ"�T�q 9�pF����>��)?��B����>%�?��?��&?ۅQ?�?��>ȭ �tC@�۔�>RY�>��W��b��@�_>��J?ޚ�>z=Y?�ԃ?��=>K�5�iꢾ�֩�8V�=l>��2? 6#?��?���>٢�>L�����=��>fc?�/�?B�o?���=l�?"<2>���>W�=*��>*��>�?�UO?��s?~�J?ď�>Ob�<i@���8��Us��tP�<�;H<��y=�c��&t��d�B��<��;C����`��4�ֹD�Ӑ�!V�;t.�>�ut>�ѕ�ף0>x[ľ�E��CA>6Ѡ��M��������9��ɸ=���>x?��>�#����=�><�>�(?�?��?��;�b�5�ھ�`K��F�>��A?j��=��l�kz��Q�u�B#g=�m?�q^?�W�6��!�_?zj?'���m�����7���ھ�>7?=��>@SP����>�̉?�|s?d+?8�m�?�u��]���Jd�������m����>�n��ߤ*�=׷>���>+q�>F��>��<`}߾��R��UJ���?;��?9��?�f�?��=6�a�mv��j>�Î���!C?l��>ģ��a5?.�2>�6�p�I0Ծ�b�W���S콝6���cA�8�̼|QB�����=�2?D�c?�6x?(n\?6s���'U���z���m���_����%�6�}�T��h5� {�BwQ�����ݟ�Am��=Ŗ�7����͸?,el?�숾�g\?�Ɲ��H��/���/���׾��}=��>���=gԚ>���Eߗ���!�,��_?��>&^�>o�?�}����@��)޾�6�L�Z>���>�>�w�>b�r<x���M����wо/k���L��8v>2yc?V�K?L�n?Pn��+1�%�����!���/��b����B>Go>���>-�W�����9&�Z>��r����y����	��~=i�2?�)�>���>�O�?�?�{	��j���ix��1����<00�>6!i?|A�>��>��ϽN� ����>&�l?Ԁ�>�ؠ>�����P!�s�{�ڛʽ!�><�>���>�
p>_r,��\��k��3����$9��.�=S�h?�����`�y�>��Q?���:
0H<�h�>d>w�9�!�M����'�m>>��?���=��;>[už�:�j�{��4��@.)?_D?�ϒ�3�*�f�~>�%"?h��>�+�>�/�?6�>-þ5s��?}�^? BJ?5A?%%�>��=g\���Ƚ�'���+=�|�>��Z>on=���=�j�mr\��x�^�D=�"�=ij˼,���P< %����J<��<3'4>DvۿlK�/'پ0��h"��	������۵�����
��!��c
��|]w�W�N�#���U�˽b�-Ԍ�V�l�K��?P�?��������7���vm���0��O��>��p���}�㉫�,��3P���`྿?��Ew!�jP�
Mi�֬e�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >^C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾u1�<��?7�-?��>Ďr�1�ɿc���{¤<���?0�@}A?�(����LV=��>�	?�?>�S1��I������T�>q<�?���?u|M=��W���	��e?�}<��F�*�ݻr�=�;�=(E=M��ÔJ>pU�>��TA��?ܽ�4>gڅ>�}"�����^����<1�]>��սb;��5Մ?�z\��f�t�/��T��sS>��T?�+�>�;�=)�,?!7H�E}Ͽ)�\�_*a?�0�?���?Z�(?Aڿ��ؚ>��ܾU�M?]D6?���>d&�2�t���=�:Ἇz������&V�{��=��>�>��,�����O��B�����=K���ƿ�K����J<��z=��;	r\��33����pϾ�i��>���o=ȼ>�r>b�>+5> �G>�`?_ua?���>�G<>��
�������	�ܻ����)�p����l8��۫��־I�ɾ��u��e���V��!=���=7R�m���E� �e�b�b�F���.?w$>L�ʾ��M���-<�pʾx����܄��ॽ�-̾�1�"n�l͟?��A?������V�L���W�w���`�W?�O�˻��ꬾ���=����a�= %�>1��=q�⾽ 3��~S���/?f?�+¾�}��E�3>���=\�-?v}?skk����>�% ?:u8�t(�Y\>AUC>�0�>��>0�>�B���+ֽ��?7�T?�$ｱ8����>����/�m�E=���=�5�~����V>�ח<���r�~��|�<#�</�[?vի>�]6��2������§�y�y=�`?�>���>xp?<6?� �=��c�h���2�N�k�p�0?,�?�;`=�>`����K��."?��]?Y�i>󰾩@)��E,�Ώ	���2?�k�?ǜN?κ�<vl��#���/�1��_8?�y?k\P����`��M<���.�>���>A0?~�&�Ӥ>/71?��C�����ξ�J�3��x�?A@kR�?��<E��h �=���>;�>e��ݾdi��L܏���+=��>�8��"�_�������E?�}?���>�k��4�a��=^P���q�?~S�?~k���ԓ<��e�l�f�����<M�=��Y����[8���Ⱦ�
�`���`Vּ2!�>?:@���3K�>�Z>��*⿃eοJj���̾�Dl�jG?�b�>]Dս��{k��u���F��JG�������>�>�ꖽ4����{�M;��{��p�>�(��Z�>��T������`��
<�.�>���>60�>���GἾ���?�f���Qο���xM�~�X?�O�?�o�?�  ?C5S<�v��}�b���$G?1s?�DZ?�|�c�Y���=�%�j?/_��~U`��4�nHE��U>�"3?�B�>L�-�;�|=#>���>�g>�#/�q�Ŀ�ٶ�����4��?��?�o�U��>b��?)s+?^i��7���[����*��,�t<A?<2>p�����!��/=��ђ���
?�}0?�{�X.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?܅�>Q��?��=�t�>[�->&kپ둮<ÙQ>1N
=�}���?�|R?-!�>n�m>�І��/%�ϫN�VH������R���k>6�X?m�U?�L�>,����\T=0�����V?�]V��z~2��۽t����>^?H>1�<>��ӽRξ��?Kp�8�ؿ j��$p'��54?'��>�?���t�H���;_?Jz�>�6��+���%���B�`��?�G�?>�?��׾S̼�><�>�I�>8�Խ����S�����7>0�B?g��D��r�o�w�>���?
�@�ծ?ki�1c	?�:��6��w�~�
����7�V��=��7?�>�|>�}�>)��=��v�Xʪ�.�s�Ǘ�>u�?��?<�>Ðl?o��CD�8�%=�[�>8�j?,�?�� :�4�b(G>�?%&�hb��>� ��d?�
@yJ@� `?�⢿aֿ5蜿c9��ꕺ��i�=��=�2>��ٽ�t�=��7=��6���>��=��>�e>��p>�O>�`;> �)>��{�!�bj��x���� D�<��x���Z�I��=<v�"��0<�����������Yý���7Q�� &�{)`�s|�=�f?�G3?��D?b�9?I����+�>$3��?���`AS�3҇>���>h�*?�o?��/?	Y�=Yվ�3A�r�s��@�K������>��\>SQ�>G??mԴ>B��=�m>��&>��>��=#ּ;�4�ث���>]��>���>�E�>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?ſf>u>�3�@e8�$�P�\|���j|>�36?�趾(C9���u��H�ubݾIM>fž>QD�l����o�%xi�:�{=�w:?��?5:���㰾I�u�7C��BRR>�:\>K=+e�=�VM>Amc�_�ƽXH�cf.=8��=��^>/�?�).>5��=
�>}��g;P�ݩ>ٹC>�,>�??�'%?������A���Y�+�!�v>8W�>�I�>��>b�L�U~�=f��>��`>G@�WZ��>��g�?�w�Y>8f{���a��|��Gr=<���.�=CX�=�� �V;�}�%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>�w��Z�������u���#=7��>�8H?�V��.�O��>�w
?�?�^�ީ����ȿJ|v����>a�?~��?�m�hA���@����>��?\gY?�ni>^h۾BaZ�S��>��@?�R?��>x9�d�'��?�޶?���?aI>���?�s?�k�>�0x��Z/��6������ p=�[;�d�>�W>f���xgF��ד��h��u�j������a>��$=,�>QE�[4���9�=��I����f�<��>�,q>"�I>W�>v� ?�a�>}��>�x=�n��Jှ����H H?�?�Z��Pl��G(=��x�IV�E�??�?%J�S{��4,�>2�d?Ŭ�?1me?�w>7� �$�����@�ܾ��L<�k�>�a?;�?�9�+&�>�Ĭ��;{��fl>���>�;��R�۾e����=�J�>('"?%1�>;�H��� ?y�#?�{j>�>�`E��7����E�a��>p��>�I?/�~?��?�Ϲ��X3�	���桿��[��4N>G�x?�P?�ӕ>a���ڄ��\|E�%I����S��?�fg?vY��?�2�?|�??w�A?/$f>T��lؾ�I�>��!? �0�A��M&�y��~?�P?/��>�7��'�ս`Iּ��������?�(\?�A&?���),a���¾�8�<r�"���U����;��D���>��>�������=�>װ=�Om��F6�*�f<�j�=��>^�=�.7��u��2�:?�a<��澊>=$�6��`��;f>��>�����>�L��/w�r���Vѕ��u'�J֜?S3�?���?M@�i��j?��~?�;?\&?��ܾ�b��H������pľA��R��=� �>/�=���3&���B��[�9�� �*x�#L�>%��>��?�� ?�mO>���>u���*�&���b��q^��8�58�<n.�M��h����"�d ��¾� |���>$���t�>[P
?��g>,,{>�[�>[�����>�GQ>��~>ݷ�>_W>�V3>�T>D<�%н�KR?8���/�'������k.B?+nd?1�>�'i�ֈ�����;�?{��?�t�?�>v>�}h�V/+��i??<�>:���o
?ˇ:=H��l�<]]�� ��!��v�v��>q>׽ :�CM�C`f��o
?�1?�ލ�̾At׽+�����xƋ?�_N?>�C�����S��~m�4g'�iaؼq�.����[�wT��˒��݋���k�8�6�p�>55?�K�?� $������Ο����6�X�>`�>:��>���>�mo<�zW��]T�6-e�3���5�qc?n��?H\>��Q?�1?�5?$�d?�t�>���>.����u�>�N��Y�>o�?X�/?b6?O�2?]�??��M>zD�Y��>Rվ"/
?���>F�>�n�>�(�>�8���O=�Y�<,������Ͻ����t(c���%�1����=7�[>�X?���Ĭ8�����dk>k�7?��>y��>���#-����<y�>�
?G�>B �"~r�c��V�>���?����=��)>���=������ҺZ�=�����=�5��Zz;�Ae<���=@��=ANt��R���3�:���;�n�<q�?k?QY�=���>'L�����"� )Q>7<�>�\�=S<4>׾A:��OƖ��L�G�_>&k�?��?@$
>�W>���=�֓�����?���0�E">��>�>A�v?!�?�?9?B?�4�=Y2������X������?d!,?Ћ�>a����ʾf�#�3���?}[?�<a�5���:)���¾��Խ��>[/�/~����!D�,.����E�����?���?VA���6��w辘��� \���C?�!�>�X�>g�>Q�)�"�g�
%�l2;>w��>�R?�#�>��O?�<{?Ǧ[?�gT>r�8�z1���ә�E3���!>B@?��?�?y?�t�>��>�)��ྔT����;�8ႾlW=	Z>Z��>�(�>K�>��=�Ƚ�Z�� �>��`�=׊b>W��>���>��>4�w>TL�<l�[?���>��(�>]�������x���"�S?k��?'�?[3i�M���5�e��r���,�8�?)A�?q�_?����v�=	 �2�Ⱦj�ݽ��>��>M� ?h�3>*��9�<�K�>N�>�Ő�Q@�������(>'�?<N?+,@�C�Ŀ@ru��nL����K�;M*���Oh�?�ƽ?en��)�=O햾z[�����@L����^��o���妾����M?�W=���=G�=�G�<�Kм���<_�=��<0q�<7E����<e�S���;��'�q8+~[<J�L=�D���`
n?X�8?�s�>/7]?�AW>e$�>�=Tv�>q�=��?�pg>%�<�:��=["=�`۾������֥���I���:��)�=EV��y��=�n�>�<K>C=j̤=���=��=C;�9�=<R�����=�U�=W�=��=-�>T8w?a���`���\4Q�Μ��:?�C�>N��=Cmƾ�@?-�>>�0��ܖ��\k��?���?�T�?��?�^i�NR�>s���9׎���=����1>ÿ�=�2����>3�J>,w�nB��pw��-�?��@2�??3ߋ���Ͽ�D/>��7>O5>��R�ن1�6�\���b�siZ�{�!?�A;�jE̾E:�>��=,*߾s�ƾ��.=��6>�cb=�V�Q\����=��z��;=��k=�Ή>I�C>/k�=�3��G�=4�I=ݣ�=ĵO>�8���8�L4,��63=,��=��b>�&>�F�><
?�X0?�'d?Q��>y�m�_�ξ����h+�>�:�=锱>-��=�B>���>Y�7?��D?��K?/z�>�Y�=ގ�>}�>�q,��m�=������;�<���? ؆?aڸ>F~H<G<B���ގ>�O�Ž\?>81?�i?�О>�U����LX&�A�.�z����sⷭ+=�ur�/pU�����u���i�=?p�>���>!�>NUy>+�9>��N>� �>j�>�d�<�v�=�1��7Ƶ<�4��-��=g����
�<&�żw5���F'���+�ބ����;ă;�l]<���;���=���>7>���>V��=z
���B/>״��-�L���=�G��>,B��4d��H~�5/�cO6�C�B>�@X>���64��?�?J�Y>�r?>E��?@u?��>�%���վMQ��pHe�`TS�	Ƹ=��>��<� {;��Y`���M��zҾ=��>K�>R�>*�l>(,�("?��w=7��a5���>@x��F��� �[6q��?��q����i���Ժp�D?NF��?��=|!~?*�I?/�?��>����ؾ$.0>�L����=�	��q�I�� ?w'? ��>�%�D�bGb�;h.�y�>x�C��4\�/��TMo�Rj���n��P�>II⾥�վ��M�@|���D��	����嶘>�u?���?�<�ܥ�t��Q����k��f}>�G�?g6�>��>Yԏ>Q.��Z��W��)4>"/�?�I�?6��?����Fm=J���>�>�J�>jh�?(��?�@t?��'���>B��<�I>kM�r��=0>�G�=>�=t�?Q@?`?I�ν6��t�(�辙`[��s^=�EO=��T>�+�>�^d>��=.4�=A��=`'f>���>%�g>�FY>^Ɵ>��>}���
�W�%?݋�=r�>�4?���>K=�8��p��<c���y!/��^�A���j���
<S�B��6=�Mg�Ba�>�'ƿKȒ?W�R>�����?Wc��'ʭ�>CG>�.J>JbԽ��>[>I܇>�>�>�И>AL>*�>�,0>�FӾ�}>y��od!��,C��R�~�Ѿ!|z>�����	&�ٟ��v��'AI�,n��ug��j�?.��p<=�XĽ<'H�?�����k���)�������?�[�>�6?�ٌ��	��ϯ>��>5Ǎ>7K��v���Zȍ��gᾗ�?D��?�Dc>��>��W?�?�1� 3��|Z��u�2!A�% e��`��ߍ�ߝ���
��+��n�_?��x?kvA?FT�<�Nz>���?��%�f᏾J/�>�/�%;���<=�:�>���,�`���Ӿ;�þ�4��JF>�o?�&�?�a?�aV��~#�<IO>j�.?��>FՀ?�`-?lV?N���� ?nv>��?8�>��"?�?�?��=���<
u]�͑�=�Z �H��ӆ�n��v[���r�=��)=V���q�=S��;������۹u+=���<!����!̼�I�=��=Mo,>���>(UU??4�>���>��8?�Gl�8�:�����5?�&��᝾@�����ʾk��D��=�2j?o��?|�g?��\>bDU��H?��u4>_��>.�>���>R��>}@<�ΏE�t�=�>c{9>���=!*���_x�
���]���/<(A@>O��>�}>픍�**'>㔢���{�e>�rP�;P��t?T��G��L1�Gu��4�>�L?ߠ?W�=�龠����f�#�(?2:<?.qM?�
�?�[�=�ھ��9���J�G���ܟ>��<�C	���������x:�d;~�t>�Ş�y�����=���e聾{k����ި
�/O��"�T�t>T��f�񾊔Q��[W>�t>�g��uq#�����d����Q?�.=��@��ᶽ�Ѿʠ1>�G�>���>gp�=�+��XL*�C1���)>��>z�>>�4 >ͭ���^I�D���>�>LQE?�V_?�j�?�"��Vs�v�B�=����c��iȼ��?�x�>Wh?�B>���=��������d��G���>q��>�����G��;���0��8�$�!��>�8?��>v�?�R?O�
?i�`?8*?`E?�'�>��������A&?2��?l�=�Խ��T�b 9�1F����>x�)?D�B����>f�?�?��&?��Q?Ƶ?,�>ĭ �kC@����>rY�>��W��b����_>��J?�>7=Y?�ԃ?�=>i�5�ꢾ�֩��U�=�>��2?�5#?^�?���>
D�>�����=�(�>X�d?��?��q?D��=�� ?�=.>t�>��=���>о�>�G?��O?=fq?.5G?��>˟c<Rq��ו��8�y�s���>q;�O<�ve=r�������v��<�)�:��]Aϼ���,�����|�;��>�w>���(>��þ����O�?>yV��o횾f�����<��|�=V�>lr ?�ڑ>��#����=Wս>���>�@��'?�?�8?�sh;��b���ؾܡM����>��A? ��=9�l��(��G[u���t=Y�m?�:_?6Y������"d?�\?����*@�:�ž��s�H�����H?�<�>�DI����>J
�?�vs?Z��>'�p�̧k��{���Y�=Q��q�=D�>EM��ޱP�郄>��!?�Y�>v>B>7<����^9d�t	���?#��?M�?���?�@7>M�|��⿖��SF����E?&��>nt�V;?��o�Q��੧��a��F���u�MJ����4�J^W��s��읾(���7=��>��a?$!p?S;S?����jc��My�����(`�E?�$���4��d:���:���]�3�'�]P�RC��b=%���h�A�?�yS?D� �"2?��ʾH�-�O]��Ǜ�>���$�n�>G�>⨵>]sսy�Ҿ:"Ӿ�(��U� ?�`�>�#�>�,?�.��9�s.��Ҿ����ꮪ=�A�>�ԙ>��X>����,I�_���a���Qc����X:v>�xc?x�K?��n?�s�o+1�:�����!���/�Rb��A�B>Ep>���>��W���p9&�
Y>���r����`x��Z�	���~=��2?�(�>P��>O�?�?A|	�j���ix��1����<�0�>� i?�A�>c�>=
н%� �3J�>��l?���>��>��| �`�y��½f�>�>.��>m�p>E�&���Z��P�������"9���=�h?��� `�WW�>�^Q?�B��<W�>���W:#�����1$��H
>�;?��=��>>�ľ�o�Y|�mԋ�z>)?+G?Jɒ�d�*�h�~>0"?_��>r�>�"�?��>�Rþ!�D���?��^?�9J?\VA?�=�>�)=����[Ƚ�&�&,=�o�>)�Z>p%m=���=���T-\�4�\�D=�*�=��ϼH߹��N<T:��+3M<6��<U�3>=�ܿK%N��оT��A8뾇����r��֎��g����۽*���Q�����t�p��=�=����*�J���\�v�f=�?<��?}Yf�0�s�a]��끿�3 �!��>'�x��,�S6���Խ��z �p������J� Kh�^Ed�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >dC�<-����뾭����ο@�����^?���>��/��o��>ߥ�>�X>�Hq>����螾s1�<��?7�-?��>Ďr�1�ɿc���x¤<���?0�@�A?r�(����e�R=1��>PT	?�Z@>��0���������>	9�?��?��K=X�W����
Xe?�"<��F��:��Y�=6��=4�=�����I>�J�>��8B�z�ܽ�#5>��>v�"�+��E]��j�<�]>U�ֽɖ�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=Fe���ƿ��"����a�=b+�<䲖�� ��۽X�%�s���ꅾ�߽�L�=]�>\W'>��s>1�P>�tL>��T?(-m?��>o�>N�aH���Jؾr�(��&���@�7����g������M�,Y�- �!.�_�Ǿ� =��=7R�z����� �&�b�I�F���.?�w$>c�ʾ��M�}�-<�pʾ�����焼m᥽O-̾v�1��!n�F͟?s�A?������V����Z�i����W?TP�����鬾��=ﲱ��=%�>댢=|�⾱ 3��~S��/:?��#?� ��X��^D>��P�+X>i�,?(c?1�����>�m-?=T���;�玛=ۄ*>���>�h?��t>�t��,
)�N?S_?m�ؽ�߯�-�v>�����k��x���g%�=�����Ҽ��>�Z>�O��[䃽��B�����b?n�>�SC���1��-��(c���Ή=�q?\�?F� >��P?/�#?*ػ�_ﾼ.a�솺��k>z
O? �`?���='S�=V܂�l_۾U-1?a�]?��>U��o��J[���˾���>C]�?��-?�����势�쭿jDؾ ?rNr?�z/�g���v�̾�x���>��>K�>E��j�=l�8?:j�������%�����P�?�@#��?�&�=&3��|�����>j?�Iǽ|���?u\�\�¾}E�<i:T>� ��s��`5� ?�x8S?J�K?���>�0��>A�X�=.������?��?磾rcx<���дi�����c��<�)�<����<��A�̾�5!�N���1���z����ŽB��>´@go7��ķ>y�l�{m���ȿ.[w�|*Ծ\]�%�?pU>'�;��ؾ��x��t�4�B�zU9���K�$�>P�>߻���P���S{�1�;�k���=��>4> �>J�>�fS�v������'<��>��>��>㏩�f���B��?>�����ͿJ���C�O�X?�f�?|n�?�?�U<*$u��y���%��G?��r?k0Z?L�"��_�fC8���j?�A��n `��m5��cD��pS>l3?�p�>ԝ,�)u=��>�1�>�E>�L.��2Ŀ����9��W��?f��?��龩��>�M�?,a+?� ��������ք+�w.���@?4�4>�-���� ��O;��u����
?�/?&���8�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\� N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�p�>W�?a��=1+�>��%�ݾ_�=�?�=W澼�!��M&?|
V?�(?k�`>\��5�S�>��mQ���eEC��T�>7gj?�EP?A�?>X�p��J'�r5d��N���Ҹ<�d�Y�����>+Q�>,�q>V����6�7�"?�1��4ȿX��+�	�!�)?�\�=}J?Cw���r��N�U��3?G�>}�'��仿<�~�'#���?�~�?F��>m����c��'�=N�>�->uE�<`�V��þ�3>�,-?���8��1c�w�>y�?iM�?���?q\w��'?��۾�����F�����=��o�=;8?��ξz	k>U�>j�=��m�g���z�x��>
�?Ҥ�?c�>!`b?�zf���C�q2�=���>3gP?%�?���<�׾I6>/�$?���)Y��:� ��wg?=�@^�
@;�R?n���a�ѿ����q��-���C`�>�ܓ>��\>F�u���<��=��ý��P�n��=5J�>q�>�
L>3�>(F>��=馄�}K$��X��z����,C�
��D�J����'�_�<��������m��/J=�lj;K���_���t3��U����>�X?KA?�L??0��>�j��U�>��ھ�J\����1��>�>n�=?&B?;�'?1�=G�����P����/�ʾpS����>0b>F�?ѻ�>�ٵ>B�=X�>��;��=�+>D
����Yϐ=mDy>-o�>�d?���>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?�f>
 u>(�3�c8���P��v��<�|>0-6?�鶾`29�Ĵu���H��bݾB+M>"��>�.B�be�����g
�Dvi���{=Zw:?�?�y���߰��u��D��mR>�}\>�=KM�=�KM>��c���ƽ�H���.=F��=�^>+�>,+:>��=>��>d�w�e�H�;L�>/�/>��>86@?{(?���~-���ۓ�?#���>���>�SY>�8�=g�J����=��>Z�e>V�½nҎ�G �LK�%��>^�=�u=�凝���g=�Fƽ�H�=�*=��ؽj�4��8�;�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>rd��j���/J����{�+r�< {�>8�W?�Ǘ��}a�#Ea��	?�l?^�T����Q¿�q��0�>���?�v�?`bR����R�S�J;?�5�?�Z? �,>��߾ڈu���0>5�3??�Z?�M�>�5���C	?˫�?Y�p?{I>���?�s?�k�>�0x��Z/��6��򖌿�p=��[;�d�>�W>`���~gF��ד��h��d�j�w����a>��$=%�>�E�?4���9�=8��H��*�f�-��>�,q>^�I>W�>g� ?�a�>���>Dy='n��Eှ������K?�w�?����.m��c�<��=��W�}�?�1?��3�ـȾ��>�a]?�?�uZ?
��>�Y�����(Ϳ�ie����<�@P>� �>��>}�����I>V�Ծ��G�:̉>5+�>陗��SپQ���:O��>��!?�`�>Z�=aG?ϰ?0�@>p�p>c�w��y���g�u?�?�?@@R?�4?� �WJ�C=���Ҡ�	O���>�e�?I�#?���>�����-��0Tk;^�3>�f��2�?���?�B��>kn�?5�W?�s,?"]�<̜���T���0�>g��>rw!?�;A��3&���=a?��?�Q�>;����ֽ+�мz���`���|?��[?n&?�S���`��¾!��<k.'���<��b�;�!a��c>ud>Nˉ�C/�=��>��=;�m��C7�ч8<���=���>`��=�G7��؎���0?�]v�-���7�q=L�q���B����>�Vl>�Ա��O?�$��*r��O���䙿_*h��t�?���?���?-���7�b��@?���?��?P�>f`��6Ծ���&�|���J���
�aU�=]��>�q��]�G���V������6���U�>zx�>��
?P?�6O><�>귘���&��A���U�]�Y9�q{8��.�(3�햟�{#�Ơ�����k{�cA�>9؊�Q��>��	?dg>�zy>}C�>��:�(�>A�O>2�|>���>+�T>��3>�o>�u<%�ҽZtR?J��'�q��̢��4+A?-�d?V��>�Rm�6��Ev���?�{�?x#�?ʅs>�wh�rs+�[?�6�>�"����	?h�L=:ϻ)h<����R��������)�f-�>vҽ��8��9L��`�4,?{?N��qyϾ,\�Cc���3�^E�?�/?�9�&�_��z�f�E�y�;���<jHy�k{ھ;/-�V�]�Y!���}��,��L�9����=[�+?�?B2������s��2�<��L�>f��>a?�>�>+>��,���m����ŗ<�����X?��?|b�>�G?��7?�r<?�%X?��j>X��>g������>�7m�Y��>�V?V�8?��&?�=0?�6?�v?m,9>ތ(�����P��<�?�|?�b"?f�?���><|~��Y꼣!N� �z���W�����=�L�<?I0�3�5��v,=���>��?g�E�8� ����j>`�6?�>��>	����P��8��<�1�>'w
?3��>�+�,r������>0��?���L=*>)>���=��j��3�����=��Ἇ��=Rkl�]�/�
��;˼�=r�=����g�9w�w;��<;��<B]?Σ?��> Ä>�����
��R
��x�=�q_>�2@>Y >_վ��������g��}�>��?���?6�p=?��=\�>s�����ž���y���R=�?֪?��U?� �?�J;?�R&?W�>m������+ ���Ǫ�Hz?q#,?J��>J���ʾ,憎�3���?�Y?t:a�Q��1)�9�¾��Խļ>QZ/��.~����tD����|��u~�����?ξ�?acA���6��r�y���Am��ÓC?�%�>]�>��>O�)��g���x0;>6l�>�Q?D#�>o�O?�;{?&�[?�kT>��8�3/���ҙ���3�E�!>a@?���?��?�y?�u�>��>d�)�v� V�����=��߂��W=CZ>��>'�>M�>���=�Ƚ�g����>��X�=ׇb>�>���>��>�w>r��<�WW?���>���r��('$���Ͼ��8�?�~�?KB>�j>�ݾ7[p���S>���? �?ͭ]?���Ձ8>��*��Y%P�E��=�_�>M��>Y�U>כ=
#p>��(?�?��E��-���$�+�o>��?{3�>Z��=)�ÿk�v�0����B�*����:��������J����">�C���6<�V����7��Yc����g��WV������4�?H%�<q
*>R�>;��<�ꕻ~�= A�=�@6=��@<D/��X�%=q� ��w�</?��_J=���<�<+B�;����Wf?��H?�f?�/?W> �>���Q�>�L">ʨ?�'>�M����;7��M�V�,]��l޾X�ܾk�_��4��x��=P�����=ߢ'>���=>H�<ڱ2>	��=�t=��$��ܥ=�?>41	>@ '=.��=�v�=t��=�6w?<������y4Q�Y�W�:?�8�>|�=$�ƾ�@?;�>>�2�������b��-?j��?�T�?s�?�si��d�>k���⎽�q�=�����=2>+��=��2�C��>��J>����J�����v4�?��@��??�ዿ��Ͽ�`/>_�8>�=>.�R��1�)Y�3cb�wY��Y!?:�:��d̾�T�>�\�=KO߾ցǾ�'=d�6>]�i=����b[�8��=��|��:=
�p=��>��A>7�=�\��9t�=�kU=u��=sN>�5ջ�2@�~�)���9=I��=?aa>s*$>��>��?L*0?�Cd?���>Fcn�U�ξ����HZ�>��=W"�>{#�=�rA>�8�>��7?��D?l�K?�Ĳ>҉=��>q��>�j,�,�m���徣���2��<M��?���?� �>,&W<=]A���hG>���Žkq?3L1?�=?���>�U����8Y&���.�#���5S4��+=�mr��QU�F���Jm�2�㽵�=�p�>���>��>8Ty>�9>��N>��>��>�6�<{p�=�������<� �����=�����<�vż*����u&�8�+�.�����;[��;G�]<k��;���=~��>�3>ˬ�>?��=y	���B/>���-�L�ì�=F��,+B��4d��I~��/�S6���B>�AX>%w���3����?��Y>�r?>H��?�?u?��>�#��վR��Me�	_S��Ǹ=N�>��<�x{;��Y`�q�M��|Ҿv	�>[�>�֢>��k>�,��?���z=��ᾑ^5����>������1e���p��-���럿%i��^�يD?�8���p�=?7~?��I?鹏?
�>%��<�ؾ��.>������=i��+�p�0���&?	!'?���>���P�D��ʾ�����>
�G��Q�A���2�@h���|��T��>Zc����Ͼ��4�|���G����C�Vt�|G�>�XQ?%Z�?"'V� 偿�P��+�T���?�j?���>u?�n?�����a����L�=�l?���?O�?��>e��=Tǒ���>�c ?�1�?w��?ӳy?��=��r�>d����&>癈�Z�=���=���=:�>E�?R ?�O?�p���e�,X��T��x��C�<鑡=xI�>N>��>���=,�=_G=`�>�߆>�N�>/�o>|%�>>��>�ؾcV-�ݣA?);�>hq>\�J?�p>+��f@��V>#7��a�0WJ=�h�=���<?S==�as�an���L��P��>�Ӽ��چ?Z�\>����v?(o��"�<aw2>o�&=�.P�T��>�.i>���>tD�>]X�>���=��s>�(Z>�Ӿj�>/��C!��RC��R�Ҿ9�z>Sh��ʡ%��������J�b���b��j��&��<=��~�<�A�?������k��*�+���\~?��>�a6?���\a����>r�>���>�t��ʓ��e���j��?[��?;-e>{i�>RV?��?lf,���6��QZ�$�t��?��Vf�S`�O̍�����
��Q���A_?-�y?�xB?b��<�z>6�?ޞ$�����j��>"�.�;���C=��>�.��h)c��nԾ�ľ���H>��n?��?!?ihW��h��D	3>>5?}�?ʹz?3�?�cR?"��%M�>z+>Go�>��>�?�.?
�
?���>F��=.������e�ѽ�ϟ��b!����^�;��=@�=` ���x�=e�u=d����߽u~ӽўٽ���M~.=�e�=�(<4�>�ϳ>�SX?���>���>�>A?уZ�Ϧ7�=��MJ2?�����̈́�����m'��r��7 >d�b?ɮ?��h?;ii>�C�3f�.�D>�ڈ>fg>W>奟>Iև���)�文=1A�=��=m��<;�ƻ�QP�WW���${���<v��=���>m7|>I獽��'>�T���z���d>��Q��Һ���S��G�0�1���v�E�>��K?\�?n��=�`�B*���Bf�')?BX<?�CM?:�?��=�۾��9���J������>ޠ�<����¢��!����:�o@�:x�s>g/�����j��=��r��vX�%%g�-{ �����>��/��d�=PU���^ς��>o>Jۂ>�HܾUD���� ����H?	��;dv��ϰ��ݞ���>���=x��>M�������9�����=�=W1?���>U��=���p(��B��:�>�OE?�W_?�j�?�"��s��B�W����e���ȼ��?;s�>7h?"B>��=����=���d�/G���>��>B����G��:���)����$���>�8?�>�?��R?��
?�`?y*?}E?E*�>��������A&?r��?v�=��Խ6�T�� 9��F� �>�)?%�B�ǻ�>L�?�?�&?ĄQ?B�?#�>r� �)C@���>DW�>��W�$a����_>��J?嘳>�;Y?�Ӄ?��=>�5��梾�橽�9�=>��2?k4#?R�?��>m�>9斾6�c=a�>�5]?hxz?2[}?R�=�?tmu>���>E��=%�>2�>�6?�]Y?,�l?�O3?|e�>���;���`����ؼ�x =!�>=�}<	��<�2:s#!<O�C����:U�<<�p�=��<B�8<s�v�M吽�����}�>��t>|*��QT0>��ľ򚉾��@>�Ǣ�UF.��e:���=��>��?�(�>��#��ђ=iּ>�>�>��	(?0�?l-?�/n;Ղb���ھXVK�;��>�QA?���==�l�\s����u���h=n?�}^?�X��T��b�b?�(^?����<���þ�d���H'P?�y
?e
E��x�>��~?�q?�#�>��f��n�0ۜ�OTa���h����=h؜>׼�">d��=�>�7?b��>O�`>�p�=x_ܾtw����8�?�?��?u�?�F+>�n�,࿮%��|��{`?1�?�5���i.?6�<�㾭`��BU����Ͼ�Ŭ�����;k�_��2
3�>ⅾ���m,�<?�y?-�c?�mV?����8l�^+d�H��� M��������&C���G�ne<�ndo��c�����m���c�=�Ӿ�y���?g�a?�����3>?ݿY����UY� ؞=�28��|��
p�>��8>1�>y�Ϻ��`����������&?U��>�<�>(B?u�6�d!������F^־0G\=TTX>ϙ]>��>!�����4�!�00���]/�QP"�8v>�xc?U�K?��n?�k�+1�������!��/��c����B>�o>躉>�W�����9&��X>���r����w��2�	�.�~=�2?�*�>���>O�?g?�z	�l��2ox�3�1�B��<�-�>F i?�@�>��>*н�� �b2�>?m?���>%�>F����!�mw�6������>tE�>\��>`f>�
,���Z�����y��HQ8�+
>��i?�9��N�V��B�>��S?�R4<�,��K�>c�����&�C����-�=Ih?�J�=�l<>����ح�$Zy�˯��%1#?�.?3���m+�Y��>��!?��>s]�>�r�?�4�> Ҽ�<n<�?�"^?�>L?��D?�Q�>�y�<Oý{c̽��0��	=p�>`j>�6�=�F�=�"��W��#�'�=�$�=Q�4�'��o�<����;L��<��/>@῏EM�����r���辻�ؾٽ%�d������nI�|�������������� �������I���Ѿ�P��P��?
Y�?�ǯ<��;�6�68���D��r>H↾�)�IhD��,� {z���꾶����R.���f��n���^���'?7����ǿL����PܾU ?� ?��y?�����"��8�}=!>���<	������N���H�ο�����_?J��>f���X��u��>:��>$�X>�~q>�)��#瞾�$�<P�?-?
��>"�r�0xɿ����\K�<���?%�@`}A?_�(�$���U="��>�	?�?>I1�gH�v����X�><�?���?��M=��W�"�	�{}e?��<D�F�A?޻) �=�?�=]O=j����J>�T�>,��c^A��Lܽ �4>�څ>V�"����Fy^��\�<D�]>��սGO��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=}��cǿ��%�%&��fB=қo=�<=��6��?!�q�h�)���/�o�^6�����=��=WF>A�>�>b�+>�hM?��p?���>�i>$9�����M���B����ci(��4n�k �gܩ�����T"�%
�v3�H���6׾!=�W�=7R�h���7� �h�b�W�F���.?$w$>v�ʾ��M�\�-<�pʾr���݄��ॽ�-̾�1�
"n�e͟?��A?������V�D���W�����O�W?P�ʻ��ꬾB��=����Ơ=$%�>�=~�⾺ 3��~S��J-?�;3?���n���T>�>���X�=Z�:?��>�d=��
?��<?��གྷ���yCS>���=�k]>���>���=���Lvؽl{?��K?�����3w��)�>ۧ����c�6�W>=��㟣;j>�H�=��B�@=������`?�p�>��4�ZD2�ʠԾ��ѽ�y��L��?�x/?�	�>��8?F�B?Bji=���߂n��
2�aO?��?�J�=�.�=*���@���g0?gK=?���>�X��]���Ț��s?�?�?9�?K�=�����G��0��C?fb�?�O�e�����3�d�`�l>��>#?������>�>?T��=�������V�����?�	@��?~�ؼ���E�=׆?�e�>����������&��n@�=m9�>������P���'��h�I0?�o?S��>�˒����+��=/���NA�?�ˑ?�v��˾�=F���v�X$�\���T�=jBѽ �༪G���j2�Q�Ծ�B�N\��y:��:�>~i@�<�m�>R ��}�鿮>ʿZt����� �#�:�>B�^>��H��nþX�|����d�:���;�tJ���>�	>Z����D����p��1=���0��>�|����{>
sP�l0��޴�������>-^�>̌>�o��>��R��?�` ��ο�✿v�
�Y�W?vZ�?��?c?}>=��P�mr����f�E?��u?}X?�?E�9�,�9с��Hn?�p��y�7�R�p�R���=fX?1�>*�����>5�Y�{��>��=E�=��^��������Ģ?/�?��ɾ[p�>_�?d5?Y�����@��ڊY�9u7���?a�>��1���.��%
���Y���>�D?�t�^3?�\�_?+�a�M�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?ӵ�� #�f6%?�>d����8Ǿ��<���>�(�>*N>lH_���u>����:�	i	>���?�~�?Qj?���� ����U>	�}?֜�>N.�?�>Fפ>ق�=�zܾ���<
��>i-l=q1%���%?�K?�>Fa>���Ir)���,�n���QD�Qqy>��I?+?��>~���L�����JF�>t��Ʀʽ�
�Q5M��rM����>��X>Ы>�|��V�M_ ?R��ەؿ�Y��Y�/���0?��v>:?h���x�i� J���b?"�>���>⳿r���L����?N��?�K?�dҾ
��W�>?;�>ωz>̈́����ؽ�Ì��[8>4�=?��%�䦊��l��"�>��?�b@p��?oi�@c?`�ڸ����\��{ľ}B����<�F;?�EǾԲ*>k��>�=��{�$����O����>�ݱ?Gb�?���>��q?OSy�D1J��a�:'`>"�g?F?�=>��� ��>�=?,i������g쾂�e?�e@tg@�?������׿�Ǡ�PV⾨�׾X*�>g��>1N ?�s�w��p��=֐��/	��S�>�J�>�*�>��W>�Ԋ>V�=���=����c��������<JK�br�<g�ק��� &�m���h�����r�ƾ@~�	�j��%�B�D��?�������y�<^�7?!``?�0l?83�>I�#=�]�=���-���w���=��?>)�1?;xZ?��3?EM=bK��Awo�zn��+�������>�9:>\�>��?*��>�A�<�K>�� >��>g	(>���<��'=!�m<��N>u��>f�?\~�>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?e�f>�u>t�3�:e8�;�P�J|���i|>�36?L鶾+D9���u���H�$cݾ�HM>)ž>xD��k�i������ui�u�{=Qx:?��?<7��4ⰾ��u��B��)QR>q:\>Y=�i�=XM>Qbc�?�ƽuH�j.=��=!�^>,�?��7>&đ=Z4�>�����W�xS�>�J>s+>�Y=?`3'?��ż�T���!~��%��p>�c�>��>K�>�jN��Ű=B��>��\>Β＂�|�F����=���V>y���]�\���m�ƻZ=$���E�=�0�=�����K>�F�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�[�>n��R����և���w���=y�>�L?��׾DH��Da���?8�?��������ſ�uz�XB�>�G�?L��?Aed��ט�|A�L��>|)�?3�W?�n\>��Ͼ]N[�|`>��B?�P?BԮ>�c�4.7��z?��?L��?�I>���?Ϟs?�k�>+x��Z/��6��ؖ��pq=��Z;d�>oW>�����gF��ד�Oh��,�j�c��j�a>�$=��>]E��3��<�=��]I��+�f�Q��>�-q>p�I>�W�>d� ?a�>@��>�}=+n������b�����K?���?����0n��8�<=�=t�^��(?�<4?d�[��Ͼ�ߨ>�\?��?��Z?�P�>w���0���⿿����O�<
�K>�$�>BQ�>��W:K>�Ծ�*D�O�> ��>�+��/Uھ�U���Ĝ��M�>Z!?ē�>Cn�=�!?�q!?pl<'g`>��c�9ʌ�a�]��{�>z�>��?7\?p�>���	eJ��2���'���t�A��=@�?w�#?�W�>Y���C���;���)">P����0�?7�?�����>j��?��O?$?�d=s.�=ӖԾ��W<h��>s�!?/ �6�A�QL&�γ��w?f?���>듒��Bս�)Լc���L����?H)\?�J&?%��a���¾��<4�$�=�P��J�;�B�V�>�>�~�� �=�F>F��=�Qm��,6���l<���=���>��=�]7�齎�?iB?2���g��S�_=�	u���C�ִ>�ɿ>t�]��CB?�<�>�>�;Ǽ��Ƙ���O�A8�?���?w$�?B�����V���??�˅?��> ��>������ƾxi�%ӽ������\�
=�/�>��=��D��������W�����=%��|��>�b�>'K?��?�]?>�ԭ>����]�$��f�4����^�
����9��A/�Uu��B��Kr �m]Ѽ����ѯz�:��> �g�>�>�?��V>�w~>���>
%E�Z��>9`>l�|>rB�>J�g>bI>�>�M�;o*ɽLR?����ٿ'�-�込���G1B?�od?3�>��h���������?���?�q�?�4v>h�L-+��n?�A�>���p
?#X:=g:�TL�<�U�� ���B��?&����>�K׽� :��M��mf�/k
?�-?�􍼡�̾{H׽Wfz�Y1�UB}?B^A?Y�H���G�l�l�`i��O�lf=`Os�*�6e&��_�:����ŕ�~�w�@a&�i:d�,?�͗?D�:��+�䱾�Տ��OB�z��>fu?$��>��>��=�J0�q�a��1\�-V-�t����z?�ז?&v�>�E?ԭ*?�$;?��T?ԆB>4��>
���l�>�м�o�>U� ?;�$?ʇ?A�3?�?�?#�>^J��O�������n��>��?x!?eU	?���>�ž�.����#C�P"��c�<z��=��E=y#-�gَ�������>�?�����9�~���d>�k6?�R�>���>���s���s�<?��>�F
?�>�{��hr����i��>툃?�� �f�
=�g'>��=:P��8B���=���}��=�~�wZ�$N+<ܵ�=��=B�F;�ڻ��N;L�L<���<}�
?^t?��[>KU>������ %���">Y�>[c�>��>�Ⱦ�f��s���P�d�"i�>Zŋ?�1�?�ܺ=^F�=�q7>U�o��AѾf�������p��=�g�>��?�^?�ܑ?�%?��G?5J>������>����è�|j ?g",?���>��� �ʾ,�ψ3���?�[?6a���n@)���¾��Խ�>z]/�S0~�Z��D���� ���y��m��?���?,A�G�6�p辯���`���C?�!�>�K�>��>��)�c�g��$�W;;>���>QR?� �>\�O?C;{?�[?SjT>X�8�N/���љ��3���!>�@?���?^�?fy?w�>��>�)��ྫU������!����JW=>Z>ߕ�>�(�>��>���=�Ƚ�b��8�>�-\�=�b>���>���>=�>w>�v�<1EN?�N�>��ݾx���v��bޚ���ƽ�:z?}��?;�?��=��
�n�S�C~�'�>=S�?�I�?��??T�M�l�'>����㶾������a>���>���>��>C�5=/@P>=��>1�>��W��C�!2.��-�3X!?#�M?���<�Eſ��r���\�������m<�f���h�ޒ���ud���=���������o�I��w��L������6䠾nX�����>�Me=(��=�B�=Q��<[��=K�]=4R�<�W=�Pj�=��<R�3��	�:����
w:%e�<�l=F����|¾�;z?�D?gw ?�(A?��W>��*>÷����>��U�ۘ?�"W>�	<�tɷ��K�η��E-��+�ξ([оi8`�@���R�>�b����>��1>���=]�<t:>�i�=��C=��*�Jtc=�J�=;2�=��=xL�=�=��=�6w?X�������4Q��Z罤�:?�8�>p{�=��ƾp@?�>>�2������zb��-?���?�T�??�?@ti��d�>L���㎽�q�=Q����=2>q��=w�2�U��>��J>���K��B����4�?��@��??�ዿТϿ9a/>�A>X�8>��E��`1��^=��n{�?xB�.�#?ձ5�Q�ξw֙>�9>9<߾գ¾ꐍ=2,>d�=YQ̽�A[�)�6=���[&=��=&�>(=F>���=����)��=K�<ʟ�=ѣx>�lԼ�z�v[���
�=�~�=�a>��%>T�>K�?U1?��d?���> 5��]�°���>�0��4��>���=a��=Ā�>h�2?�]Q?udJ?��>$��=W�>h��>��5��a���得g��r3�h�?�A�?O��>nd�=V����02�[;	<݅?�9?�� ?gO�>�U����:Y&���.�������0�+=�mr��RU�y����m�>����=�p�>���>��>MTy>��9>��N>x�>�>9�<�p�=3ꌻd��<����=������<�użO���6}&���+������;竆;�]<R��;��	>��>O��=��>�V�=^þ��%>���O�B�Bڐ�zN���+J�!�g��{�A@5���*�ިP>�h]>޴!�,���E�>��z>��t>�"�?I�d?���=}%ڽh�ܾ�1������
+��=��=c��&�N�R���Q��̾���>;Ƹ>�->��2>_f3�� C�
�o=��޾D��o�y>���ig��v}� &e�e릿i[��\�I��=5�C?'���� �=�~?@qh?���?���>>D������%�<6��F�5=*���#���½�v?iN?�?�|��D�̾�o����>2�H���O��Õ���0�������C�>D���о&13��l��:폿�^B��
r�!��>p�O?��?�bb�?`��MO�`��nׅ��^?Ύg?t*�>Jp?�`?�����u�Ta�����=]�n?��?kE�?��
>;��=DJ��7M�><	?6��?���?j�r?�?�T)�>U��;J� >��;w�=�i>�Х=6��=�?�W	?!�	?�-��G
����ﾜQ[�,M�<�=�O�>��>R@q>>=�=f�c=�=l�Y>��>��>cd>���>��>,�޾��)��N?@�~>[~e>+J`?��=�ලA����B=~Ե=a�������H>ʇ�=���x�� ��P�BI�>������?�v�>q	���.%?+Ce��`=��>��>/o�,��>Xi:>��N>�k~>:v�>�a^>[�>8��>�?Ӿ��>���Ne!��.C�W�R���ѾL�z>����� &�����g���@I�Gq���k�E
j��.���:=� ~�<+G�?#����k���)�����ԕ?�[�>�6?Ҍ�5����>���>͍>�G�������ƍ��e���?���?�d�>3�>�3?? ?�o<X����V�mjW���!��?��)0v�
���Uk��R&�&���i?y�k?�0?N�=��b>O�[?Ǘ�p6#����>S� ��zI�߷�=���>k)q������f�����^=l����>_X�?�Ut?G?�D4��2��]�<>5g�>�->� s?���>Y?�V�^_)?��>��>�>r.?�?�V)?���>;�B>%�	��<~0��������ٽi�5�1�#��G>1>e>���=�_�=�����]F���=�)>�t�<���=<��=P�B�G��<�w�>h ^?���>Ĉ>��9?Y'�Gy8�r����7.?&W<���f����Ϧ��F��{��=@�k?���?N�X?7i>��?�HD���>�ӌ>3 5>�Y>��>�����>�p�=��>��">J��=�i��m���vЎ����<ٯ>���>%5|>v��~�'>�{��6z�ԣd>
�Q��ʺ��T���G���1�@�v��V�>\�K?��?.��=�\�p&��If�'/)?^<?�OM?��?R�=��۾��9���J��K�k�>�z�<������L"����:���:$�s>�1��
�	  �   zР��db>���j޾��n�J����qL=݁�E�U={�*�վ&'����=k:
>[����� ����Ī��#J?��j="\��n�U��n��9>kǘ>�خ>�`:�!Jv�W�@��Ƭ�yY�=.��>�
;>�������gG�Y)�m�>�-3?�BJ?��?W���Y�d�X�P��G��þ���� ?=j�>f��>��>�y7>��s������D�p�?��>���>\����=�Ȯ`�E����b<�H}>0:�>X>�P�>�(?�_?�Bi?�?���>�]>���貾��?"fv?{0
>��6���<��%0�I$8��>V��>���Y�0>ϕ�>��
?jM?>\?:�?�)��9�>�x�>	�>��K�iִ��U�=�GQ?U�?w�o?�9�?��>JHW��V����Rf>w�U>j�?Q� ?E� ?4��>���>Z���?�=��>�	c?�0�?�o?�~�=��?492>y��>D��=��>M��>�?�WO?*�s?��J?đ�>'��<�1���8��xBs��P���;��H<M�y=���4t��X�C��<���;mj��;�����S�D�K��U��;k��>$�@>{����>xk����MЧ=!�#>*��ƈȾ!ϔ<�K	>���=�?�%�>ʍ���[����>xȫ>
��*�Y?MR�>p�7?c��>�L��6�=������*}=��=?���>�(#�!~�یS��H�L�l?��M?Y������K�b?��]?4h��=��þs�b����b�O?9�
?(�G���>��~?_�q?d��>��e�%:n�'���Cb���j�)Ѷ=]r�>LX�O�d�p?�>r�7?�N�>&�b>z%�=^u۾�w��q��c?��?�?���?+*>��n�R4࿨���rˑ���]?�@�>�3���"?�|"�hrϾ�7��я���ᾴ���IЫ�:���B���#?$��y��!ԽH��=p8?�s?B�q?}�_?� ���c�)4^�65���'V��u�w��
�E��eD�0�C��,o��5���������G=hqy�y<�L��?TO(?%H8�f�>�ȓ��.��UҾ5�">-Ɣ�1��r=�=+儽�zV=��=lV�i&8������?gd�>J&�>5E6?�~T�ac@�^ 9�	�3��I뾟�>�>33�>J�>�T="��ĽHPɾ:�c��iн,(v>mbc?gK?i�n?j'�)<1�b����!�L2�cK����B>0a>���>�WW����53&�A=>���r�_���q����	�33�=��2?a�>�>m=�?4�?�k	�H쮾j�w��}1���<��>�h?=%�>X0�>�ҽ� �Os�>hpm?���>)!�>V炾��!�9�{��8ϽK��>e��>��>�?`>�80�|/[�*}�����p)6��>�g?5�����V����>��P?�D�;�<��>Z\��W3!�~���7'�Ċ>U@?;ʉ=�(>,ž�
��y�1��_?y?�YW� �9��q�jdA?�<?+BP���?���>{�[��
�_�>���?���?҇�>u���X�>w��>�Z<_���; T<�'�>�-��B�>'�Z>m��A�w>�B��}=&�C=$�����3Ƽy0[����O�x>3�!>���W�D�4���m����۾����7��Q�`��2����z���P5������9�3���ڛV���S;����@��K�?/��? <���訾Rʌ� Mw�A�����>Syu�K�H�� ���LM�l񨾢ھeƾ�>)��|V�c�X��qE�H�'?����ٽǿ��;ܾ'! ?�A ?1�y?��R�"�Œ8��� >wC�<�'��9�뾬�����οߦ����^?���>���/��l��>ǥ�>�X>�Hq>����螾�.�<��?4�-?;��>v�r��ɿY���V��<���?�@��G?sGr�ܦ ���>>U�>�@?�,�<�u8�u�$��D˼��i?�I�?pƒ?�:ݾ�"]����>F.�?��"�GC��A�=��0�r�,>В�=V��"�>k��>b�2��ڽ��ļ����Լp>y��~_�)S���������@�0*�=)Մ?�z\�Zf���/��T��{U>��T?�*�>�;�=��,?o7H�X}Ͽ�\��*a?�0�?Ѧ�?��(?�ڿ�ٚ>l�ܾv�M?-D6?���>�d&���t�ۅ�=�8ἐw��I���&V�S��=4��>2�>��,����O�`H�����=��-���j1��"�{�<}Z��Lٽ��+��8�<B<�`��#~F�Ih6�a��;]�>XvV>�\G>�q$>h�F>Sa?�r?��>�$�=ߌo����	�߾M:=��y��N��y����P��+��=7�|�ܾ��)C-�v��A��"K�-�=�U�A��k����ƃ�dHU���S?�9�>�E��B�R�������i��-=�< Yмh��`�-�-����?u�&?Jyk��b�BG��ɔ<x��W�A?;54�e���GǾ�>HT�=&�?>Tb�>�u>�%��$�(~.�vs0?�K?5f��@��3*>�� �Q�= �+?�y?)LY<�*�>/3%?+�*��+��[>�3>n��>���>�	>���hM۽K�?D�T?���j͜�3ސ>�F��i�z�BBa=n>FC5����.L[>��<����{U�*���ֺ<�'W?둍>��)�<��V{��e���">=�x?W�??�>Zkk?n�B?1P�<I����S��"��(w=��W?~#i?Ĳ>tʁ�:�Ͼdj��ִ5?W�e?��N>!h�a��o�.��O�<#?��n?�X?e���z}�]��p��-b6?��v?s^�ns�����5�V��=�>�[�>���>��9��k�>"�>?�#��G�������Y4�Þ?��@w��?%�;<��;��=�;?~\�>ޫO��>ƾ{z������/�q=�"�>����zev����R,�Y�8?͠�?���>�������[��=�����G�?f�?͍��.g<����Cl����k��<N8�=)���!�B����7�/�ƾ��
��������9��>DP@�W� ��>�7�p/�[Ͽ����R)оyQq���?�j�>�ǽ�
��Uyj�7&u���G��H��������>��>K+����\�W�M�q�ʽ�5?���<�R�=w����!��"/��P�b=��>���>Hٕ>G&������?�����ǿp����%:g?�\�?j�W??��>�'��s�j�<�� 	G>y�Q?��a?�`B?�IQ� _Q��⿽�j?e`��iU`�6�4��HE��U>`#3?I@�>M�-�?�|=�>Ƌ�>Rj>#/��Ŀ�ض�9������?X��?�o꾟��>��?-s+?�i��7��)Z����*�+��;A?02>�����!�0=��В�'�
?w}0?m{��-�r<X??�\���q��'<�	|���W�>f9�r(-�+P����I�q�i��J��`v��?�+�?��?M�a���'?sν>�`��~jԾ,=���>���>��\>ֽ_>>o����2��)>!�?�\�?_?W�cΥ���>�p?t�>.	�?*N�=��>���=Nޱ��Y�g#>ô�=B���?MM?��>5E�=ep9��/�1�E�)�Q�����C�U2�>�9b?*�L?��b>[h���3��d!�{DͽL-/�`(���?��*��x��S2>�h=>�W>�	F��Ӿ��?Op�9�ؿj�� p'��54?+��>�?����t�=���;_?az�>�6��+���%���B�]��?�G�?B�?��׾�S̼>=�>�I�>6�Խ����o�����7>=�B?;��D��x�o�Z�>���?
�@�ծ?vi��	?C�@O��Yn~��z�1B7�Gr�=��7?���z>���>��=qsv����c�s�x��>�>�?_v�?���>��l?�{o���B�-1==R�>Ŕk?�t?�Tc���򾉙B>{�? ����>�'f?��
@v@�^?_袿��ε��ϵ��ߥ��=�Y����A<���p��=c�3>�3:&�������6�C>J�|>��,> �=��!>��;>�����s"����̛�����z����(��xν�6�O �����!������q�̽�Hk�?Ƚ9���f@�������=l�U?�R?p?L� ?�Mx�ֱ>r���4E=��#��̈́=�'�>c]2?�L?P�*?q��=㝝���d�S]��/:������ʓ�>�aI>�o�>\A�>��>\Х8��I>]?>v��>�>�'=��Ժ@=��N>�K�>���>\m�>0<>�k>mʴ� N��uh���w�kr̽@�?�N����J�/9��"�������C�=�x.?��>7���п^˭�(KH?i���J�Ab+��B>��0?8aW?O6>\����V��>^��B�h��>~ �� m��)�$Q>�&?B�f>cu>��3�Z28�԰P�y~��N�|>��5?)@���.9�ȹu��H�.AݾSM>���>#@�@]��󖿂�~���i�'{=Gs:?e?�̳�tf����t��\��UR>{\>H�=:ũ=AAM>O�b��ǽ!=H�p%.=�q�=�`^>�?� #>&�w=Wh�>.ɛ�]�>�=�>�#>�Z>΁9?s�$?�1����������4���|>^�>�o>ȥ�=a E���=�>�>�_>�8	����%���XG�Ec>����~zT��a��Ȃ=+A���h
>E��=G���y�-�M�=uz?0���DS�k�޾	�I�N�J?�? ?���=TV>=���@��ҾJ�?��	@���?Zv��\�N�,?�j�?�֗��#W=�v�>a_�>�ž+/E�BM?^	P<+7��3����U9�?���?��߁�Ont�;u�=��!?:�Ծ���>ˌN�M���j����`��!0<�i�>N=>?P뾂5}��}��?�_?.8��e3��ެ��E�]�J��>7n�?^��?d@��������
���>i��?"�N?5��;����@E�]?��Q?���?w��>�I���P���&?�"�?�K&?�B>��?.%t?���>�Y%�1�+��l������S�I=�_O�*ԋ>���=��žR�G���o����h�I����\>Eu=��>�{�\��\X�=�hX�����6c����>�o>��A>#�>ƌ�>[~�>ڢ�>�=8��!�'��w�K?���?���2n�kL�<���=Ѳ^��&?~I4?(h[���ϾKը>κ\?u?�[?d�>>��;>��*迿~��A��<2�K>4�>4H�>�#���FK>��Ծ(4D�rp�>�ϗ>����?ھ�,���O��;B�>�e!?y��>Ӯ=љ ?��#?Ζj>3*�>�`E��9����E����>o��>�H?s�~?��?�ӹ��Y3�l���桿�[��:N>��x?V?�ɕ>9���փ��S|E�|8I�5���㛂?ftg?�Q�9?2�?A�??��A?�%f>r���ؾ������>�?�l��l0�9�-�}�G��	?.X
?r��>R���j��X�ɑ(�/v���%?��f?��?����qI�n?���#=^�;dk8��?;����d>I�>>��ʽ?�H>W<3><<�?���C!�C��<e��=�/�>d��=}U:�?2���<,?��G�ރ���="�r��xD���>�DL>����^?�l=���{����x��9U�� �?��?�i�?;����h��$=?��?�?!&�>{L���޾W��"Xw��xx�+x���>U��>^�l�N徨���"���F���Ž�0�?<2�>�?NT?�R#>D��>}�ؾ�M�	c��j徥�(�j��bE��e�d�˾��~���G�.� �ᘮ�m���O>˲�_�>g�&?���>��=#X>�O�=���>��g><�>H�m>T�W>��3>Ռ�=�*w��QzK?ؾJ>����H�S�F�7�@?[?ܖ?Bh�>������/�>��5?]�?��?p㓿��5���]?$f�>��6����>����d�=�7�>��Wq)��M�>�+���Hk���>���%hN������!?�6�>��&�ٽ�\=���""o=bN�?a�(?/�)�o�Q���o�r�W��S�:���4h��l����$�:�p��쏿�]���#����(�W�*=d�*?��?t��v����E#k��?��\f>���>�%�>�ݾ>/wI>��	���1��^�YL'������N�>CX{?��>B�I?ݯ<?�%P?a�L?ʕ�>�ե>!/���[�>�ݕ;�>B4�>��8?�-?#�.?��?�+?'Fe>:�����־�W?d?m(?%?LA?p���%½6mn�ui�@�w�q���֨k=��<�tٽؘj�(QP=��R>�f?z��K8�h���c>&�7?d��>�A�>Z����5���G�<�*�>��
?>�>q��j�q��`��G�>~��?���G�=j�)>F��=k���V�#�0Z�=|�̼� �=~���פ?���<�^�=S�=x85�l :9�9MC�;^,�<P�>� ?��>�N�>��� �S����=^�X>A�R>��>�Uپ;{���#����g�2y>�h�?�o�?E�g=���=���=���Y�����᣽�-.�<=�?�#?!@T?R��?��=?�H#?Z>11�"C���^�����֋?,?2��>[����ʾbᨿ��3�"�?^X?�/a�_���1)���¾cսY�>�U/�w ~�9���*�C����$������?���?�#@�2�6����Ę��d��!�C?��>�L�>+�>��)���g�"��L;>�v�>� R?�d�>`sI?MUq?T-m?�uE>��@�wt������j� �}b>�bM?�u?Yg�?�j}?�X�>L��=C���ξ����e�Y���m�5>�<1x1>]�>�G�>��y>���=	F��K�\J>��v/>�:>l�>'�>;��>�d�=9�I��"H?'��>c达ED��t��M���J��yu?)�?��*?�)=h�"=D�ǧ�����>�(�?;x�?�)?�JW��.�='q�e����s�F��>��>���>Q��=y�:=�>�l�>�g�>%=�b�^P8��H���?`;F?`��=�ǿ��q�(Ut��Ù�/�
<ҟ���mg��ᒽ
�R��K�=m���-#�·��S}]����9���>����G��u�u�# ?��=���=�:�=���<J�o�<~$s=:O�<uR=�i��	�<�D2�Dt�����Bf����<>�Q=�e�9��|��?�4�?��?��B?�s2=�L�=�ڽ��Y>�i-?\fh>�4��/����Q�u�J�~�¾]3Q�p����F�( ��i8�>�ʶ;�ڽ�$�a�-<N�'��-�>��*>K��<�E���̼0u�=p�>�%�<��j=AVn=�Č>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��N>22�=�M�H�-�/U�?06���p��_#?��9�,ƾ���>�Z�=��ɾ��̾�E8���E>|�=@=$���]�N��=���jm=c*l=G�>��X>��=�����C�=�}=���=�gH>ק�%;���WY���=�Y�=�y>��'>���>|?<-?zi?�>
�x����x���B��>�Q�=���>C�=fY>�:�>�W2?��8?��K?'T�>�ɩ<9'�>�y�>��,��Ru��O澺P��[I=K3�?&��?�޲>-�9<��B���v�@�����?��:?�Z�>�ύ>����ֿU<"��P1����S2��"��`S�#�<B�=1(�Vp���Z=g}�>f_�>
�>�$q>\_>�mb>���>"��=�r������;SRJ�UG�:�ZW>��=��W=��q��C�=�U�<�#;̰~<���;�ц=/=���x��=s �>�p=͍�>��=��̾��>�m��u9X���8=㾬�Q*�+�U�]�x�p,�"O�.�+>���=o��j���ޞ�>`_m>�%>`ֽ?�i?��:>���!��x������
��§u=��=��{�b@�h�^�p&G��m̾���>���>��>Wm>��+��0?�jWu=���/T5�s��>#X�����1�%q�O,��퟿��h��z���D?(>��bH�=�)~?�I?�ڏ?�m�>B���a�ؾ��/>A����4=2��sq��'����?��&?8��>G0��D�`��^y��E>A@ھ�/��롿��F��A>^�\���H>O���>Ӿ��M�Ɔ}��I��;'4��듾큩>WgP?��?���WK�c�m��־ۋϽg�?�n?���>b��>��>s־�P�ʾ�N��6<>�z?�?y+�?r�>D=�=ڭ����>A�?�j�?̳�?~�r?��=�r~�>r��;9�>5Օ�+8�=�>>���=3�=Y�?#R
?c�	?�4����	�ܸ��	�_�#��<�T�= .�>S��>:�n>~8�=��_=p�=��]>�8�>4)�>�a>Ť>���>�/��r�	�"?�>�|>�a1?ʃ�>i痼����.(�;����6�SO(�5FĽ��ｈF)= ��;s5�<�����>��i��?UK>���5e?�@딽n�|>�v>�#����>F�G>L�>h�>��>2@#><�>��>�8��>J��$�|�?�nV�2�۾߿�>QL���2�y,��t��}]��緾��|_h��ӂ�<�*�=<�?"UȽ-�g�FQ.�E���j?<��>��4?IL��4���n>���>��>�H�������r���޾.�?c�?p�]>N��>=T?b!?��9�D�*�DDU��=|��A���f���Y������}���[����`?��v?�v:?%N<�V>��?����a���u�>�2��A�ZmG=���>�P����[�(;)�����役�`>�m?��?5?�WQ�c�m�k-'>ճ:?�1?�Nt?��1?��;?����$?~3>�C?�n?\I5?t�.?R�
? 2>���= ����'=S8��(g�ѽf�ʽ���3=�[{=�M����<ܢ=��<����ټ�;���#�<	:=��=�$�= ė>aVa?^�?O�>�Q@?�^���A� a���h ?U�k<~�h������e��M��<-#S?�c�?��V?*%|>A�S�T����g>)ٓ>��/>���>��>3�$��@�P�=��=�/>�"=u+�<���,��D~�m/;�>h�>�@�>�	����)>��/�wh��O��=O�ͽ�ڭ������!���%�,��㾒>�w+?�?�vh=�疾�!!=h�n�p�@?��Q?��8?�1�?HW{�)/��&N���\��¯��+Z>�Eս+ט�봑��S���1�<>��K��Ϡ��b>�����޾3n���I����fJ=]p�6P=i��վX5�<�=[2
>�鿾#s ��䖿�����rJ?�j=�<��$�V�#y��&q>͔�>�>Ψ9��ez���@� o��x��=�_�>n7=>�㓼%��cG�՟��z�>=YD?'[?v��?�g����u��]@�ȃ�������&�U�?�ª>��?sQH>�'�=U������=�`�4C�U)�>��>���߄E����a����$�LR�>�?K>�?ՑQ?�
?�c?
V)?2� ? J�>�o��0��f;&?��??�=��Խ��T��9��F�,��>�p)?�RC�X��>��?�?��&?k~Q?��?-�> � ��#@�>'A�>ؼW�q_��q�_>īJ?���>]iY?�у?��=>�l5�좾�����=��>_�2?��"?�?�ڸ>j4�>���� ��=G��>�db?`;�?��o?� �=\�?�/>��>�;�=�X�>���>��?a,N? s?)K?F��>|R�<)櫽�ٶ�gfq���'���5;�H&<~�v=�����l�l0�/,�<��;���6���z�����B�	*����	<h��>[�=F}}�	��>�Խ���L��<E>��L>t����O���"{%> ܂>���>ѥ~>�\��=y�>j�S>� D�J?Z7�>H�?2~��RK�O����^�a��>�?]?�Y>\�Z��k�����t���d?k�5?:B���c��K�b?��]?h��=�#�þ-�b�t��g�O?0�
?��G���>��~?X�q?m��>��e�%:n�&���Cb���j�8Ѷ=r�>)X�K�d�Z?�>�7?�N�>,�b>�%�=7u۾!�w��q��a?x�?�?���?�**>s�n�Q4�g>���?��k
^?��>�Q��C#?������Ͼ�+��#����Q��.���6��&W��!�$��䃾��ֽ�3�=�?s?�Cq?;�_?�� �d�!*^���Q]V���t���E��E���C���n��R����w	����H=� p��l7�oA�?;|1?`X����>Z肾����#;�4�=2������x�=[���X8��t=*/Խ�W��K���*?<M�>5��>p?p�\��E��+�8�7�?%پ>��=�_�>��>&��>/,>6��W�;#S�7�r��ͼ<�iT>��k?(\P?7�i?�*�bk;��ن�}c����������b>\K=D�X>��m�,�5���$��m@��l�[��}��������<V�/?�_v>�#�>�?�l?c&���5��@�z�+#���<�?�>��i?0��>�ځ>�+�,&��ٖ>�b�?�n?fe�=z�;�O<�rMv��1��I>�^�>z�?��Ƚ�݃��Ee��T����zB%���I>��K?�.��2R1���>
�h?� =݁��(�=�ԛ�;��o־���n�=ZY�>���=��>୩�(��d�s�Q���)?>?�:��_�*�UyX>�%?���>�֠>���?�K�>�Ѿ�jW;��	?�NZ?`;L?�LB?�t�>���<�͒�5-��&�%�q��<���>�\>i�E=3\�=\8 �+�Y�c��"�^=	V�=�4��>�Ƚy�,<��'��g�<u�<��@>d��F�G���̾����.��d'��L-��Z�a�VEнaQ���K����t��&�+c���6M�-�7�T鋾��j��b�?y^�?����2h�pY��0�i�V|
��>���aF��OE��8oϽ+ш�����Ѣ�kl��z:�v�Z�1@W���&?������ȿb0���]ھ�?%�?Tq{?���ơ#�p�:��&>�=q����\㾴8����Ϳ����V�\?��>�[��T���74�>���>j�T>�u>%T��ﭢ�HM�<V�?{B1?
�?X�`�~hʿ��%�<�^�?-@�;?h ��V�}xJ>���>ذ> �=�n�1RR�Q��P>���?���?�� ?�[��X��@�?Uͽ�Q9���Ä���Y>#m>܌�<]��!�Y>���>����ؙ�(�`���B>�c�=Vq���:�6�����>O�>�������V�?��R��Z�1=/��8r���L>)>?�n�>+�$>+?}�=�c�ƿ޿]�X�;?��?k��?�D?r����д>��޾2�I?��;?;)�>Qe�̉_�O!>�\��i=B��aO�#l7>���>�?�=�?�61�7����=��="���sſ��"����
=���:��d��������=�����d�i�}��b?N=$��=��N>7Y�>�R>��U>�8Z?=�h?O��>�>��ֽ�1��f\Ѿ�-<}�v���&��Պ�׳�A}������޾%c�<�����+Ǿ��}�F+��* ���h���l��%��f�m�;��?n�>Ĩ�[��z�>�q�$���[�����=N=���y�7����?�?�n��@Ae���s7޽�u>��U?7Pu�[`��Ӿ�5��kN���<l��>��>Ʉ{��)߾%A�l�/?c�?@a������QO=��=��=�?�	@?�f�<G80>v�?��n�����v�>j|�>��=�Mk>�:�>آ־/��U�?��:?ן���7���&�><Ҿ+v����O=[��ͽ̳��Xs�>	�T�_����h=yQ>�a=T?��>�)�5!�� %ٽ��=�}p?$�>$9�>k?o~@?R.(<4���I��A��[O=lX?�h?E�>��߽��þ������0?=�g?`T>��@�����43����9?ˣm?F?���2��
��������)?��v?�r^��s����)�V�=�>+[�>���>��9�\k�>�>?�#��G��𺿿OY4�"Þ?��@j��?X�;<��ۜ�=�;?c[�>f�O��>ƾ{��ރ��͐q=W"�>�����ev����R,���8?砃?Z��>d������K��=���q�?�φ?�@���z�;���_�k��t��ݒ<���=&��xG+��쾝86��uľht
�Ὓ��/��^�>�,@�@����>��.���⿭kϿ���`Ӿ^.}���?V��>ľý�띾�Cj���u�J�F�[�F�o������>���=7��K̲��6i�ay3���J�73�>;񴽺�K���>�
Ej������i]>�Ƭ>\f?y�F>/ݼ�*�^�?�^�3���^��$��X�N?5��?O��?�Y?�H��[Ŋ��5��[p<R�=?>��?�l?�.��/:�n">�j?x_��iU`���4�dHE��U>�"3?�B�>T�-���|=�>b��>�f>�#/�s�Ŀ�ٶ�6���X��?��?�o�!��>q��?ks+?�i�8���[����*�
�+��<A?�2>���B�!�D0=�ZҒ���
?N~0??{�g.�KA?۟Y����vg�f�ڃ>�X����0=J��Q��#�}�O ��̋�����?��?��?~� �w���`?z?����CȾ�Қ>�K�>O��>f��>k�o��L�=Ѩ���K�%C�>,��?f� @_��>D뭿7U��Fq�>��b?�>��?���=�R�>+��=E���ڮ-��Z#>l��=0�>�ޢ?}�M?x@�>z0�=5�8��/�.WF�@R���C���>��a?"�L?�Ib>.��]2�C!�zͽm1����nN@�Q�,�'�߽�5>�=>�>��D��Ӿ��?Hp�>�ؿj��p'��54?���>2�?����t����;_?*z�>�6��+���%��LB�Z��?�G�?P�?d�׾gQ̼i>�>�I�>,�Խ����������7>�B?���D��t�o���>���?�@�ծ?\i����>,H�ܦ��D>��۰��o9��x�=��F?��F$c>z��>���=0�w�J����,n���>�s�?�C�?�v�>��q?�Y_�_�7��L��a��>�t^?�?�c��F��/>�e�>0��N�������g?`Y	@M�
@,[?����Fhֿ`���!M��ᗺ����=4��=��2>�ٽ�]�=d�7=�8��;�����=l�>:�d>iq>�'O>ra;>��)>S����!�=r��͢��L�C���-����Z�־�YXv� z�Q3�������<���2ýBw���Q��1&�q<`�P+�=-�U?R?��o?� ?����>�����z=o�!�*z�=��>�1?�@L?�Z*?��=������d�1^��B���{Ǉ����>�+I>)�>~��>��>
��:�I>�
>>t�>Z>�s)=� ��'=��N>w�>�8�>z�>�"<>�z>�Ӵ�">��0�h�=w���̽��?�~���J�\/��fJ��
���}+�=�j.?��>3��8п�뭿HH?�"��#-���+���>�0?�bW?,�>Y��~U��>����1j��>�p����l�T�)�pQ>wl?��q>��p>��.���7���M��m��d�s>\ 6?�x����0�ks�+D���߾��)>���>Y��<��!������v��s���=��;?{?N�޽L����W��֡���a>�9P>��<]��=9�Q>*�a�8�� �P�O%�<'>]�\>�?hp>���=	��>�ז�L̜��m�>��W>'��>*�6?
?-�-R�Gͧ��C��ơ>��>���=F�K>�^u���>�Q�>t�M>�ݬ�C�=��F_�0iM��^�>w�"���v���;��=U�B��=��=n;�8ҏ��+4=kln?7o���zվ�3��?���>s�u>��1���'��D���d����?�S@j#�?�$&�=N��G?�zo?�T>=p��N�
?@?�dt��L�e�>��t��s���̺�\�~��ϻ?��?���<eѪ�'��'mz>��%?���X��>����r����u�]�=���>�H?ӡ�� a��9:���
?��?��"��e�ȿ/�u�
7�>=~�?��?W�o��8����@����>�+�?EZ?�k>�C۾��[�J��>�A?)R?�e�>�Z�?�,��|?yg�?���? *4>��?��u?��>��<�28��������rޚ<0'�<!�>x�,=!�ɾ]?G��V�����z�g����0@U>�;x��>輽:ᒾ��=�䠽�>��o�&�>�O}>�22><�>��>	��>V�>S\2=�ɽR���"!����K?���?(���2n��N�<���=!�^��&?�I4?�j[���Ͼ�ը>ߺ\?e?�[?d�>A��P>��A迿=~��>��<��K>%4�>�H�>�$���FK>��Ծ�4D�ap�>�ϗ>e����?ھ�,��T��>B�>�e!?���>�Ү=��?}�#?��_>���>o�C�`z���CD�@ѽ>���>�j?�W~?�d?������-� #�������Y���W>)�x?��?��>E��YU����4�����8����?˽`?����?眈?��??�%B?H�Y>�J+�ܒԾ-����p>��9?�ʋ�ݡ�,��8���L?<�+?���>��?~�>������0�*�o��==��?g��?]o!�����UA>�q=�ߴ=ޖ��x<���>�g%=gW㾩$�;�4�=���=���>,�ľ��U�����^��=E��>\%g>׾�J�=�6,?DDB�������=��r��tD�H�>heL>����,�^?�(=���{�1	��bu��HU���?��?Jf�?B���h�6?=?.�?ܸ??��>�����޾�}�!x���x�J�>���>~�i�6;�V���(��5���Ž^�]��z?���>E!?�+?i򗽖�q>�^ξ�8�%�;�oƾ�b�dh���B3�+J��#�oD�id#�I!G��u�B����e�>Ru��3;>�V"?���=���>�y�>w]�@>��%>8��=�P`>�&{>+�e>I1>Q�Y�H�ýäL?2����;߽/����I� �H?Ѩ�?���>����b�o������?S�d?+��?���>�vT�bg>���?;Z�>;�L��ƙ>�f>lu5<�ܣ�_�ý/=��H���~>��?A�ҾO����!��&u��"�>���>7(���x����<���;o=�M�?��(?��)���Q���o���W��S����5h��j��P�$��p��쏿�^���$��J�(��r*=Q�*?9�?���\��!���&k��?�ef>'�>"$�>�߾>vtI>��	��1�^��L'�I���R�>�Z{?!��>�|I?��;?ZuP?�ZL?��>�U�>�<��FG�>��;H�>1��>#�9?:�-?i30?a`?j`+?�fc>��R�����ؾ5�?��?xI?g?r�?�����ýy�����d�>�y�a_����=S��<�ؽ�8u�s"U=��S>� ,?
�H����~7����K>��#?5��>�#>�-���X����<2(�>�*?���>����\�|�r�����>(r?�K��m'�:���=�0�=�y\=��սGM�<��O�	���-��=.�|�8*e���Y=���<�X=x�<uD��3�<JN=�t�>E�?���>�C�>�@��[� ����>f�=>Y>�!S>'>�Fپ�}��t$��V�g��]y>�v�?.z�?j�f=��=���=1}���V������������<P�?$H#?�VT?:��?�=?�i#?�>�+�RM���]�����=�?~*,?�A�>�N���ʾ�è�< 2�3z?�H?n_���DN)�ʓ���=׽w�
>G.�S�|�b��.TD��պ�������L�?g�?ՌQ���6������S��?C?�%�>���>P��>�)�P�g��4��I;>g�>�Q?��>jN?Y�v?��[?!�O>e`<��U���Ř�@e���>\J??�?(f�?�~y?���>}�>�3-�os׾���Z�XB��j��1G=�Y>ݸ�>�b�>���>z_�=a�۽D���Y�7�W٦=��g>|�>��>�]�>�>��9<�H?�%�>ѹ���x��b3j��=��*s?��?��*?���<F0�zCF����T�>��?�r�?�3?�7��;�=�����#��q�k�/��>I��>bŜ>�w�=H�M=�o>!5�>Yd�><�����5���p�?IrG?$��=s!�k4h�V����g���NC�����׋�-�>��$���>��OX�|���i���ب�yVK�#3���k������?�	�=�<b��<:�=j�%=�Ws=�=��6=��>=�b)<Bq�=i�k��Q1=�uJ������2=fǜ=EV�<,�&�pS�?<|>?�)$?�"�?��Ͻnf;�?��� �=�/?"{F?{+C��������0ľ�Nq��P۽[��p�!s���k�]�b=k��<a����>�H,>.����L#>I��=�h�=%@>"�=��W=��"=��=��F>;,=�c$>\�v?#r��]͝���Q�h�}k:?�(�>���=��ƾ(�??J�>>$&��ʓ��j~��?���?sN�?��?�wi��r�>dV�����'э=����%)2>���=ޥ3�2�>�I>��yE������v$�?�@T�??a�����Ͽ��/>�8>��>W�R�sn1�	�\�JDb�n�Z���!?|;�-*̾�.�>=(�=�3߾X�ƾuA1=�&7>�ya=G�z\�
��=Rhz��M>=ul= �>�5D>ӊ�=�>��ܷ=vJH=���=NNP>6��*18�3]+�U�2=)[�=f�b>ͧ%>h�>�?��/?Γc?���>�In��<;���
��>Zi�=�ԯ>��=��@>�q�>�7?�EC?޾I?Z�>s��=�>��>�H+�e�l�%�侧����<Ǻ�?s��?!ݸ>��n<�H?��?���=�q����?tc/?��?�ߞ>%���߿j8$�.�����\l��E=�w��J�E�ݼ@��	��3G�=�C�>1��>�m�>	Gy>��1>��F>���>�">�y�<`�g=���[��<=ZE�Ա�=�����=4T����K;�-�� )�Kk��+*�;��;5!l<+] <۫�=��	?|��=0ic>���>��9�>4n����I�;\'>�<&��O^��iD�b�j�F�:�{��r>�W�>�{�<oj��Ʌ? �>-8���?�`7?���=#(8�:,��y��a+��F���{�=�,Q�Ώ��z�G���6�E�+�ES����>q6�>+�>G�k>u�+��3?���u=%�Ep5���>X���!�7]�_q�%$��G埿��h�V�ˉD?�C��h�=[~?�I?�ˏ?B>�>�m��mDؾL�/> ��=��fPq�͓���?��&?�:�>�-���D���оY�ý�Q�>'�M��dN�ش��t!1�D�u9w=���C�>h���W�;\�2������p��W�@�l�k�HJ�>�HN?�U�?�\�� ��5�O�QK�����:?��g?iߜ>�
?8�?�x��,��}���L=�=��n?��?���?Uq
>h��=l���?��>ו?4�?Y�?�q?T�F����>�)�>� >,��Z��=O�>��=7�=�	?%:?��
?)��b	�m��+��K�T�x�<�b�=�o�>JŁ>�z>p�=�_=���=%V>��>���>|1`>� >�~�>�T�e>��	�>��K>�=�?W�>Ӆ�=',0�o����<;�k�hJҽ���<���@�ͽ��]=�->�O��X��>ȿ�˚?�=)��y3�D<N?T�+�gW;���>�7�=B_��v�>��[>�^�>N��>u�F>*��=x\{>���WҾ��>5��F �O�B�mwS��~Ѿ�y>ή��.�(��������I�Rʳ�-���i���I-<���<��?MN�|�j��)�1����	?4��>/o6?э�rǎ�P>�@�>�a�>ѭ��no��O��R�ྟ
�?v��?�N`>�"�>�V?�?wx4��2���X���v�0�@���e�!�_���������	�1&ɽ��^?�z?��@?��F<
�>�T�?�1#��Ր�tg�>,�/�c�:��$="ȧ>����A`���Ͼ�b¾�;���O>ȟp?"˂?<�?�3M�� =]0�=�>?aL*?=�\?2u6?�C.?�J��?F��=��?���> �??��??pJ ?&>�<��=��=��=mHA�l���"��F˽/�c=�~5��0��� 6��8Ƚf�=&�~���CH=�})�>2��{�<��=�=�g >���>�]?��>�1�>v	7?L!��8�L���,�.?q#0=����T��������Rs>�kj?�G�?��Y?�}f>RgA�,�C��>�|�>iL'>X[>4u�>e|��G��|=��>�V>�0�=�1@��#���
�"5��5.�<w�>31�>���>����Rd8>�&������>��.�5ȼ���<#1?� |���"��K��=�9=?�b'?A���X��-X]>s?e��"G?��>��%?�z�?�A�4"�����l3��_&þ֔?���̰���ڼ����Y���>��>�B|��d���S}>���avs��>N�Gap���ܾ��὎V$��\>r���Uھ��.���>E��=D����	�ꯞ��Q��1�-?-��=u��)�H�V���;V>�l�>�~g>4 	�SJ��y&�gu���t�=�\S>Õ>�0�����H_��6�!z>2�=?L*U?�T�?�r����t�ţ=�u\�m��Siu���?wc�>we?��g>�m�=���M��U_��G>�2��>���>���G�>�M���V&��$��ȇ>�N?Q��=&�?�D?���>XWi?&<)?h�?��~>�G��|k�b.&?�{�?�݄=#ӽ4U�9��F�Ho�>o)?v�C�ݢ�>�]?�?�
'?�wQ?��?	�>�� ���?��ݕ>vD�>�W��M��p�_>?�J?��>zY?�Ƀ?-e=>n5�K����&���[�=��>��2?E�"?��?F�>��>б��~�=ڠ�>� c?=1�?��o?���=��? 2>��>��=���>0��>$?�QO?��s?��J?D��>�ʍ<�A���l��J>s���N��Ё;��F<�Kz=7��s�t��+����<?d�;�ⷼL	�������D�u֐���;��?�(h>f]5�Vo�>g���N��2�>�^x>#�޽��/�}�w����=��=&r�>���>��(��������>w>6����Z?��>���>yS��"^�
�����ƾ�5�>-_3?vD�M�Q�2Ƈ�m�p�Y^���f�?�<I?t��Q쌾Z�b?��]?�g�=���þ��b�q�龐�O?��
?��G�\�>��~?E�q?^��>��e�d:n����Cb���j��ж=sr�>MX�@�d��?�>�7?�M�>P�b>C$�=.u۾��w��q��g?c�?��?���?+*>8�n�4��u������^?t��>3����"?��ɻ�eϾ�g���\��!�����#��6������#\#����Q�׽nX�=7q?EBs?}�p?�L_?�g ��d�^��
���AV���������E��(E��|C��~n����m�������I=U��-�6�9:�?�Y?�c־�v
?e R=ԍ��i��n�>�5���K-�j�:���=��T>}.6>�ʅ�xk\�-��t8?�u>�ș=�2?�� ��D.���H�P��>����Hٽ���>��<�K�>k�s=x��"�v=8����9��6E=�u>�uc?*�J?��n?� �ȭ1�68��s�!��A��ͧ��&C>̛>�2�>� W�����%��>�%=s�����ŏ�=
��=}.2?3�>pN�>hؗ?/%?S��������u���0�"\�<���>#�g?4��>��>��ӽQ� �s�>L��?<��>�d�>�ڸ�� ��w�}�O=�>��>R	?�W$=�mC��"Z��@��a ��>Y9��ld>j�W?������E��q>�DP?��9�	��;>Zs��~"����ۿ�_>��>t$/=;H>�uǾ���������̾2?9�G>ұ�>v���޾��R?U��? c�==B�?��M?��q��z>Ĝ?>E7?D5\?p?��G)h��7�=�N�����/	>,��=�;>:�=�+�<�f��2ǐ�丅:
q
=�%���Va="�=���c�>5E���5>ZjۿY>K���پ��_�8E
�n鈾Vǲ�-h��;��Fc������Nx����'��V�X+c������l����??;�?�{���,��@�������x�����>Ɩq��������#��`'��J��)����e!���O��*i�w�e���'?/���I�ǿ籡�6ܾ� ?y> ?�y?��h�"�˓8��� >4��<$"���� ���'�ο۝�� �^?��>��k��5�>$��>]�X>�Dq>�������<N�<#�?Ɇ-?���>cr���ɿΎ��X{�<���?�@�E4?j����e��m(>�<?u�?c��=��ɾ��(�8!@�̳�>3t�?�4�?�6�>yʂ�����KҜ?�s������̓=�{���j����>MS� �=��>�� �R\n��t���<>�Ҏ> ʷ�=�m�M�Vw
��b>fͽ�m�����?S�\�:�`���*�t���nB>(�S?<��>�a�=߈$?�IF�>jͿ<�X�O�[?�E�?:;�?�? ?�����>6\پl�H?h�.?9��>'"�xor�ef�=�J�;�����PQ�'��=\��>�>f�)��(
�J-S�+5u��d�=��6�ƿ��$�<����=��뺛�[��x�A�����T�����fo���v h=p�=YxQ>,e�>QW>u=Z>�dW?8�k?�O�>?�>�.�Rz��ξ�,@���������I���裾NN�w�߾��	�������-�ɾYUN��b�<�e�����/��9Jh���L��G1?��>+���U�+��Z���U�:*ݾ3���>вU��1���f���?,� ?�e^��]I�N�a�>8����aV?Ӭ��oܾTK۾��=����	j>hx?d&�>!ڿ��M�%H��C0?Z�!?v���m�mv/>(c"��<<�C(?��>n��@��>B�?8�,�� ��;�>��>za�>���>�&>�Т�:Ʋ�,�?�fX?���ߊ���b�>!���Sgw�bL_=N40>f�L���a���n>�
<O䈾�����ν�
=�W?>"�>�O&�ȉ��5����0?=�y?�g?���>��l?�FD?ə�<L���P���1�|=��W?��e?��>�)t���Ҿ�ҩ���6?�$a?m5>b�Z�KO뾟F-��x���?^n?�?h�k�6�{��������1�4?��v?s^�vs�����@�V�`=�>�[�>���>��9��k�>�>?�#��G������yY4�$Þ?��@���?��;< �g��=�;?f\�>�O��>ƾ{�������q=�"�>����ev����R,�d�8?ܠ�?���>��������">��Su�?沀?�f��Z꾼����^��-��?Ҡ�v4�=2�:��$=ݾc��Ϯ�<Q��|s�c=om>U�@��$�Pt?����D�i�п/Uv�O��w��n�C?�^�>*qr�PW��sG����#�/�Y~6��m����>�>{��:w��Iz�WE���X�:��>pIC>g����\�7������o�|>38�>c�G?7�=�"8�~�}<Xϒ?ˊ������B����� ~�?�G�?�h�?� D?��>�/��������ݶ�>)�|?{?T!��O25��̆=7�j?b_��U`�o�4�/HE��U>�"3?D�>8�-�հ|=?>`��>g>j#/�)�Ŀ�ٶ�$���b��?���?so�a��>x��?�s+?�i��7���Z����*��1)�=A?>2>Ԍ��T�!�_0=�CҒ��
?�}0?�|�6.���7?��S���d���Y�ߟ��>z�>�s��o���	>o�%���^�����!���ˢ?_�?1��?�C�]�
�t
?��?ܦ�1�Ѿ	�>�)>u*�>�d)>w=ӽ ���?� ���"��@�=��?��?L�?�T���#��O��>��i?�\�>�$�?���=c��>�v�=�F��i�M��"#>�w�=&�O��q?}VL?y��>�#�=m�1���.���E�LQ������B�N=�>ka?I�L?/od>:U��yu8��O ���ν\1��ļ�&B���%��ڽj3>�2=>%�>Z�H�VҾ��?p��ؿ2j��)n'��44?�>��?X��u�t�n��\;_?(y�>R7��+���%��iA�E��?HG�?W�?}�׾�Y̼v
>%�>�I�>r�Խ����:�����7>��B?��tD����o���>���?��@�ծ?gi�Ǜ�>M[�{%��fe��^���>�V���=�4?��־�t>S�>�G�=V�v��9��	jr���>&'�?w�?�"�>|nm?��i�r?A��T�<���>��h?C	?~�1=b��EH>�#?I
������n����e?H
@��@U?����h�ȿa]s��޾������>-m.�y�z=��SG<�=o�,==���<�]}=�#U=(�9>ڤ>r�T�D�o>�l��+���Ŀ������@�w���7��b��$��k)�/���E��A��\��ʮa��Ȕ�?D��y#H>_�=B�I?H�8?�t?���>A�?�>ܧ�y� ��L(�|�=�^>��*?"�??��?�6�=eH��� p��M��Nא��O�����>��]>R?�>Tu�>J
�>୞��M�>��=.�>��=��H=g�=�:�;��>�ڸ>U� ? y�>�,<>��>δ�6��K�h� w��5̽;��?Pg��۶J�I/��;�������X�=�a.?6�>���<п ����9H?����$���+��>��0?3dW?��>���iU�f>e���vj��>����?�l�Ě)��Q>�n?:�i>�Dh>��2��%5��XR�81��>Z�>(�2?����=���u��H��ھ�N>�<�>x�y�f�!�����|�B}m���=?�:?5�?m�ɽtŲ�mj��j��9cN>!�f>*�	=妯=�n>>�뀽��׽<w;��FU=&�=�`Y>9+ ?\�3>�͕=Y`�>�����Hn���>�U>���=�S:?i�?�K
�>�f���6�=����]>K��>a�>���=] S�d�>:_�>�o>��<1н<�����Y�rwm>t��<!pk��3E��o&=#\�7�t=��=�%�5愾�^�<��h?E����Z������i����B?���>�dO=(��!�����:��r��?�@;܏?�o�t�I��>%?$�w?8��< �p���?yH?��X��i/����>���)��������(���?�A�?� ��L����8t��d�>�D?m����o�>�t�8V��;����u�z�#=V��>�7H?�Z���P���=��w
??U򾠥����ȿ\xv����>��?��?��m��<���@�Rs�>��?�kY?qi>g^۾�bZ�m��>r�@?R?��>�@��'�;�?)ݶ?��?�G>H̑?Zs?P��>fl���.����������%w=�M�;�>R�=���B�F������5����j�����a>ڣ=k�>Q�佺X����=-�$���6m�mQ�>��p>��H>��>�� ?��>*f�>��=���lw��\�����K?���?���2n��M�<���=ݲ^��&?�I4?�h[�f�Ͼ�ը>к\?`?�[?d�>;��G>��<迿I~�����<x�K>�3�>�H�>�%���FK>��Ծ�4D�ap�>�ϗ>�����?ھ-���X��wB�>�e!?���>�Ү=k� ?�#?U�j>�M�>�TE�
/����E�J��>�_�>�#?$�~?1�?�����<3��Aۡ���[�49N>��x?UT?�K�>|������U�L���D�̑���?cg?]j��?�>�?��??��A?�=e>����׾������>	0?F��P&�����s��n�?n�?�� ?kǓ=Ĕ���f��_N��վ�>#l|?��H?Zz ���M�t�K�	>���r��K��;������R�ئ�=�)>Ҍ/��:�=[�>Y4�6q��F]�r؞����<UX>��Q=�Ľ�����#,?
GD��惾���=7�r�]�D��x>8�K>f����^?9[=���{�r����^��x�T�z��?v��?�\�? ��֕h��1=?B�?3?rn�>�n����޾:yྰnw��(x��W�K�>0��>�1l��	�U���댪�6?��*ƽ��0�̛?&�>�?��?�	�=��}>��h��~,���qԾ��b��W	���;�4�.�l9�����i��E�Q��5����c�o��>�J@�I�y>��?�8>��5>gB�>��/��ٍ>z`>+��>�~�>�K!>K�>�4�=�ѣ�ď��*O?Č����$��慨�ͥ�q�8?��/?���>��K�����¾6�?���?�C�?OX�>1�{�Z���>f��>Nl:�r�%?PU�=*�Ƚ����<���ݘ��֑=HX%>�Ӄ>����g��u�>����&?��&?t�`�Z̾k�ɼ0�����n=tM�?M�(?��)���Q���o���W��S�����5h��j��s�$� �p��쏿*^���$���(��c*=Y�*?��?������"���%k�y?��`f>��>E"�>�߾>�sI>h�	���1�^��K'�u���1S�>�[{?�
�>�
J?��:?�iQ?xK?���>	#�>�0��o�>O�=��Х>���>�7?�_.?D�2?��?��)?:�_>L}潠,��]�ؾQ+?��?j~?�s?�?���ƽ�Y�������z��np�v��=s�<��ս�w���>=kqR>"U5?��"��X��ᮈ�E
G>"�U?=�>�.?[Q�cg��б>{;?�S?���>Rˣ���V����?)�5?W����(=.ж=�=���=�N��k��;�7> &�;�n{=����R׽�%=�1a=>x�=���_K��>�=��>,�0?*��>���>un&�wp��%��G`!>f>��k>=8>� �s���s��ƺd�b�f>Y;�?v�?��=�L�=�b>�w��䩷� �Z��f��<��?�� ?�K?�D�?-�8?��%?��">ґ��ъ�9���k9���>?�,?Dq�>���c�ʾ ���o3�@�?�Z?Oa�)p�DO)��b¾�HսH�>�@/��~�;	��<D��҂�4������e��?ʯ�?�vA�M�6��V�����c��ԜC?���>�S�>��>F�)���g�\$�~C;>�x�>��Q?Q��>)QQ?�u?�^?�}U>�<�=��]{���#��f�=h[E?Gy?��?܄x?@�>�>��)���ܾ�f�iżJ`��Elk�!��=�vZ>��>���>�ë>t�=�Ǽ�j�q���D�r.�=��k>��>��>>i�>��^>���<�F?"��>�f����������*��gK@�Vt?_��?�(?s-=1��
E�d8�� �><�?���?-�+?��?�=+�=�(�������
s��	�>��>�>�>ǘ�=�J=��
>��>��>�W�yC�e�5�H�`��J?|�H?���=v4翓��{5�U>Q�4�>7�f7��w����+������%�)�%0���0�N	&�u���Ӿ�W��F�>�?��f���>ɺ�<B�T=��;��c<D����u>��<��9<P��ѳ���=���<��.=Wp�=?'�=��1�����<�?.?��?[?��D>���猽iͥ<��>�'?��-�#� �$u��H���r��]]��n#������Q��?����U= d�B��=�X>)�
>��*��#C>���=	��=���=�=7=}	>��=�j>ǣ�>��J��]$=��u?�J��$���E�R�7���9?���>e��=,�þ
�??�a=>3�����b�U�~?J��?�?�?0�?�pk����>M>��������=�w��B�5>��=�3��s�>�I>��������Z����?n�@[K??�P��\Ͽ�61>��2>�(>E�Q���,��IZ�01o�i Y�$m?ǭ=�0Nɾ[ �>�^�=�yھ@-ľ�"=1i2>�U=�L+���]�*w�=	���0F=	�y=�<�>��K>��=����]�=J�=1\�=�lO>����=���7�n�?=���=�rb>�Y >Q��>uA?�u*?SRb?�3�>�M���:̾�1Ծ�͂>�� =��>s�����> ��>��/?jNI?~�@?�ӫ>�M�=�D�>�;�>��#� d�X�ɾ�!����/���?DCi?"v>J;6=��f�:���m'����W?��?=\?�f�>�U����>Y&���.���K7�+=�mr�wQU�����:m�9��i�=�p�>}��>��>&Ty>
�9>��N>��>��>�6�<Xp�=�������<� ��z��=������<vż�����t&�-�+�����v�;㱆;%�]<���;���=���>��>��>�*�=�ҹ���(>%�����L�<��=9���KA���a�݉z��w,�y 0���F>�LW>�A�� ��[�?X>��E>M0�?��p?�{>�?�U$־'ל��;[���T�>��=H!	>�t;�� <�*�_���N���Ѿ8��>f�>�>��l>%,� ?��w=���K^5���> \��p���6�=+q��.��=�	i�vqº��D?	A��ZQ�=�~?D�I?�?e�>v���|ؾ
0>5V���A=6��q�����?� '?���>��$�D���	�_nѽLkN>wxƾ��!�����:�����;2_�İ�>����� Ǿ�:�Fc������7I0�	2���>��>?sO�?��l��yr��9Y�1����*��>�yl?Q��>��	?�"�>M�w��ھ��V�T8>Z�x?���?���?��-=	��=���4��>�\	?�Ǖ?>�?ws?r:�=t�>�j�r�%> h�����=;�>S^�=���=��?q�
?)�	?S'���(	� F�Ϙ��0Z����<&��=�>�
�>op>D�=L�\="�=��[>^��>g��>�]e>--�>�T�>�>׽�Ӿ�%?竊>�/��??�>���=�y�=�"�;RE6��O���=�������=��=(�J����;#�=��>J�ƿq��?��M�HA&��8?ꋄ��uw��z>�y�>󋌾��%?�v�=�l�=o�/=z��=p�=^��>��������>Ȼ%�+/�U0���\�`��@�x>�ܯ��fK�jx����kx�Կؾ����[g�C
}���>�y��=G�q?j�*�p�p�;a@�Z�ƽ���>�>�8?�2���wz>6��>��]>($��77������MӾrh�?��?��W>��>5!S?|?��"�WP�3-T��co��4�� Z�L��X���;z�i��ʽ�b?mz?Q�D?�Y=KWV>���?g �h���.�>�\,���A�)�=A��>�!ƾk�3��r�3jž����I>��c?�{?Zp)?M����(E�v">��:?��1?Cq?|4?u�;?��~�"?�]&>Z�?Y�?^;4?�.?Z^	?�>E��=�`
�e1=fĐ��y��)�ӽJ�˽�GӼAxA=��c=�B<L<�S=+x�<�	�������;�J���#<0;G=Qo�=�=/>ޞ�?���>���>��R?4>.�u/�����eY�>05�=[��<��M�۾�Y �a*=�\;?~�?�A�?�y�>ۇK��RH�e��=�l�>�{>a�?>5|>&���p���=�D=���=��=A!1��F���'��:��v�=��w=.��>���=�zq���J>�(��Z��t��>�lf��`{���ս:6�ִ��∾�7�>��A?��5?�*�=�������;�}_��5�?�'�>~@E?n4�?l�ξ�1��'��T�@x�=��	?�=�Oо��S������m��<�>��>l��zР��db>���j޾��n�J����qL=݁�E�U={�*�վ&'����=k:
>[����� ����Ī��#J?��j="\��n�U��n��9>kǘ>�خ>�`:�!Jv�W�@��Ƭ�yY�=.��>�
;>�������gG�Y)�m�>�-3?�BJ?��?W���Y�d�X�P��G��þ���� ?=j�>f��>��>�y7>��s������D�p�?��>���>\����=�Ȯ`�E����b<�H}>0:�>X>�P�>�(?�_?�Bi?�?���>�]>���貾��?"fv?{0
>��6���<��%0�I$8��>V��>���Y�0>ϕ�>��
?jM?>\?:�?�)��9�>�x�>	�>��K�iִ��U�=�GQ?U�?w�o?�9�?��>JHW��V����Rf>w�U>j�?Q� ?E� ?4��>���>Z���?�=��>�	c?�0�?�o?�~�=��?492>y��>D��=��>M��>�?�WO?*�s?��J?đ�>'��<�1���8��xBs��P���;��H<M�y=���4t��X�C��<���;mj��;�����S�D�K��U��;k��>$�@>{����>xk����MЧ=!�#>*��ƈȾ!ϔ<�K	>���=�?�%�>ʍ���[����>xȫ>
��*�Y?MR�>p�7?c��>�L��6�=������*}=��=?���>�(#�!~�یS��H�L�l?��M?Y������K�b?��]?4h��=��þs�b����b�O?9�
?(�G���>��~?_�q?d��>��e�%:n�'���Cb���j�)Ѷ=]r�>LX�O�d�p?�>r�7?�N�>&�b>z%�=^u۾�w��q��c?��?�?���?+*>��n�R4࿨���rˑ���]?�@�>�3���"?�|"�hrϾ�7��я���ᾴ���IЫ�:���B���#?$��y��!ԽH��=p8?�s?B�q?}�_?� ���c�)4^�65���'V��u�w��
�E��eD�0�C��,o��5���������G=hqy�y<�L��?TO(?%H8�f�>�ȓ��.��UҾ5�">-Ɣ�1��r=�=+儽�zV=��=lV�i&8������?gd�>J&�>5E6?�~T�ac@�^ 9�	�3��I뾟�>�>33�>J�>�T="��ĽHPɾ:�c��iн,(v>mbc?gK?i�n?j'�)<1�b����!�L2�cK����B>0a>���>�WW����53&�A=>���r�_���q����	�33�=��2?a�>�>m=�?4�?�k	�H쮾j�w��}1���<��>�h?=%�>X0�>�ҽ� �Os�>hpm?���>)!�>V炾��!�9�{��8ϽK��>e��>��>�?`>�80�|/[�*}�����p)6��>�g?5�����V����>��P?�D�;�<��>Z\��W3!�~���7'�Ċ>U@?;ʉ=�(>,ž�
��y�1��_?y?�YW� �9��q�jdA?�<?+BP���?���>{�[��
�_�>���?���?҇�>u���X�>w��>�Z<_���; T<�'�>�-��B�>'�Z>m��A�w>�B��}=&�C=$�����3Ƽy0[����O�x>3�!>���W�D�4���m����۾����7��Q�`��2����z���P5������9�3���ڛV���S;����@��K�?/��? <���訾Rʌ� Mw�A�����>Syu�K�H�� ���LM�l񨾢ھeƾ�>)��|V�c�X��qE�H�'?����ٽǿ��;ܾ'! ?�A ?1�y?��R�"�Œ8��� >wC�<�'��9�뾬�����οߦ����^?���>���/��l��>ǥ�>�X>�Hq>����螾�.�<��?4�-?;��>v�r��ɿY���V��<���?�@��G?sGr�ܦ ���>>U�>�@?�,�<�u8�u�$��D˼��i?�I�?pƒ?�:ݾ�"]����>F.�?��"�GC��A�=��0�r�,>В�=V��"�>k��>b�2��ڽ��ļ����Լp>y��~_�)S���������@�0*�=)Մ?�z\�Zf���/��T��{U>��T?�*�>�;�=��,?o7H�X}Ͽ�\��*a?�0�?Ѧ�?��(?�ڿ�ٚ>l�ܾv�M?-D6?���>�d&���t�ۅ�=�8ἐw��I���&V�S��=4��>2�>��,����O�`H�����=��-���j1��"�{�<}Z��Lٽ��+��8�<B<�`��#~F�Ih6�a��;]�>XvV>�\G>�q$>h�F>Sa?�r?��>�$�=ߌo����	�߾M:=��y��N��y����P��+��=7�|�ܾ��)C-�v��A��"K�-�=�U�A��k����ƃ�dHU���S?�9�>�E��B�R�������i��-=�< Yмh��`�-�-����?u�&?Jyk��b�BG��ɔ<x��W�A?;54�e���GǾ�>HT�=&�?>Tb�>�u>�%��$�(~.�vs0?�K?5f��@��3*>�� �Q�= �+?�y?)LY<�*�>/3%?+�*��+��[>�3>n��>���>�	>���hM۽K�?D�T?���j͜�3ސ>�F��i�z�BBa=n>FC5����.L[>��<����{U�*���ֺ<�'W?둍>��)�<��V{��e���">=�x?W�??�>Zkk?n�B?1P�<I����S��"��(w=��W?~#i?Ĳ>tʁ�:�Ͼdj��ִ5?W�e?��N>!h�a��o�.��O�<#?��n?�X?e���z}�]��p��-b6?��v?s^�ns�����5�V��=�>�[�>���>��9��k�>"�>?�#��G�������Y4�Þ?��@w��?%�;<��;��=�;?~\�>ޫO��>ƾ{z������/�q=�"�>����zev����R,�Y�8?͠�?���>�������[��=�����G�?f�?͍��.g<����Cl����k��<N8�=)���!�B����7�/�ƾ��
��������9��>DP@�W� ��>�7�p/�[Ͽ����R)оyQq���?�j�>�ǽ�
��Uyj�7&u���G��H��������>��>K+����\�W�M�q�ʽ�5?���<�R�=w����!��"/��P�b=��>���>Hٕ>G&������?�����ǿp����%:g?�\�?j�W??��>�'��s�j�<�� 	G>y�Q?��a?�`B?�IQ� _Q��⿽�j?e`��iU`�6�4��HE��U>`#3?I@�>M�-�?�|=�>Ƌ�>Rj>#/��Ŀ�ض�9������?X��?�o꾟��>��?-s+?�i��7��)Z����*�+��;A?02>�����!�0=��В�'�
?w}0?m{��-�r<X??�\���q��'<�	|���W�>f9�r(-�+P����I�q�i��J��`v��?�+�?��?M�a���'?sν>�`��~jԾ,=���>���>��\>ֽ_>>o����2��)>!�?�\�?_?W�cΥ���>�p?t�>.	�?*N�=��>���=Nޱ��Y�g#>ô�=B���?MM?��>5E�=ep9��/�1�E�)�Q�����C�U2�>�9b?*�L?��b>[h���3��d!�{DͽL-/�`(���?��*��x��S2>�h=>�W>�	F��Ӿ��?Op�9�ؿj�� p'��54?+��>�?����t�=���;_?az�>�6��+���%���B�]��?�G�?B�?��׾�S̼>=�>�I�>6�Խ����o�����7>=�B?;��D��x�o�Z�>���?
�@�ծ?vi��	?C�@O��Yn~��z�1B7�Gr�=��7?���z>���>��=qsv����c�s�x��>�>�?_v�?���>��l?�{o���B�-1==R�>Ŕk?�t?�Tc���򾉙B>{�? ����>�'f?��
@v@�^?_袿��ε��ϵ��ߥ��=�Y����A<���p��=c�3>�3:&�������6�C>J�|>��,> �=��!>��;>�����s"����̛�����z����(��xν�6�O �����!������q�̽�Hk�?Ƚ9���f@�������=l�U?�R?p?L� ?�Mx�ֱ>r���4E=��#��̈́=�'�>c]2?�L?P�*?q��=㝝���d�S]��/:������ʓ�>�aI>�o�>\A�>��>\Х8��I>]?>v��>�>�'=��Ժ@=��N>�K�>���>\m�>0<>�k>mʴ� N��uh���w�kr̽@�?�N����J�/9��"�������C�=�x.?��>7���п^˭�(KH?i���J�Ab+��B>��0?8aW?O6>\����V��>^��B�h��>~ �� m��)�$Q>�&?B�f>cu>��3�Z28�԰P�y~��N�|>��5?)@���.9�ȹu��H�.AݾSM>���>#@�@]��󖿂�~���i�'{=Gs:?e?�̳�tf����t��\��UR>{\>H�=:ũ=AAM>O�b��ǽ!=H�p%.=�q�=�`^>�?� #>&�w=Wh�>.ɛ�]�>�=�>�#>�Z>΁9?s�$?�1����������4���|>^�>�o>ȥ�=a E���=�>�>�_>�8	����%���XG�Ec>����~zT��a��Ȃ=+A���h
>E��=G���y�-�M�=uz?0���DS�k�޾	�I�N�J?�? ?���=TV>=���@��ҾJ�?��	@���?Zv��\�N�,?�j�?�֗��#W=�v�>a_�>�ž+/E�BM?^	P<+7��3����U9�?���?��߁�Ont�;u�=��!?:�Ծ���>ˌN�M���j����`��!0<�i�>N=>?P뾂5}��}��?�_?.8��e3��ެ��E�]�J��>7n�?^��?d@��������
���>i��?"�N?5��;����@E�]?��Q?���?w��>�I���P���&?�"�?�K&?�B>��?.%t?���>�Y%�1�+��l������S�I=�_O�*ԋ>���=��žR�G���o����h�I����\>Eu=��>�{�\��\X�=�hX�����6c����>�o>��A>#�>ƌ�>[~�>ڢ�>�=8��!�'��w�K?���?���2n�kL�<���=Ѳ^��&?~I4?(h[���ϾKը>κ\?u?�[?d�>>��;>��*迿~��A��<2�K>4�>4H�>�#���FK>��Ծ(4D�rp�>�ϗ>����?ھ�,���O��;B�>�e!?y��>Ӯ=љ ?��#?Ζj>3*�>�`E��9����E����>o��>�H?s�~?��?�ӹ��Y3�l���桿�[��:N>��x?V?�ɕ>9���փ��S|E�|8I�5���㛂?ftg?�Q�9?2�?A�??��A?�%f>r���ؾ������>�?�l��l0�9�-�}�G��	?.X
?r��>R���j��X�ɑ(�/v���%?��f?��?����qI�n?���#=^�;dk8��?;����d>I�>>��ʽ?�H>W<3><<�?���C!�C��<e��=�/�>d��=}U:�?2���<,?��G�ރ���="�r��xD���>�DL>����^?�l=���{����x��9U�� �?��?�i�?;����h��$=?��?�?!&�>{L���޾W��"Xw��xx�+x���>U��>^�l�N徨���"���F���Ž�0�?<2�>�?NT?�R#>D��>}�ؾ�M�	c��j徥�(�j��bE��e�d�˾��~���G�.� �ᘮ�m���O>˲�_�>g�&?���>��=#X>�O�=���>��g><�>H�m>T�W>��3>Ռ�=�*w��QzK?ؾJ>����H�S�F�7�@?[?ܖ?Bh�>������/�>��5?]�?��?p㓿��5���]?$f�>��6����>����d�=�7�>��Wq)��M�>�+���Hk���>���%hN������!?�6�>��&�ٽ�\=���""o=bN�?a�(?/�)�o�Q���o�r�W��S�:���4h��l����$�:�p��쏿�]���#����(�W�*=d�*?��?t��v����E#k��?��\f>���>�%�>�ݾ>/wI>��	���1��^�YL'������N�>CX{?��>B�I?ݯ<?�%P?a�L?ʕ�>�ե>!/���[�>�ݕ;�>B4�>��8?�-?#�.?��?�+?'Fe>:�����־�W?d?m(?%?LA?p���%½6mn�ui�@�w�q���֨k=��<�tٽؘj�(QP=��R>�f?z��K8�h���c>&�7?d��>�A�>Z����5���G�<�*�>��
?>�>q��j�q��`��G�>~��?���G�=j�)>F��=k���V�#�0Z�=|�̼� �=~���פ?���<�^�=S�=x85�l :9�9MC�;^,�<P�>� ?��>�N�>��� �S����=^�X>A�R>��>�Uپ;{���#����g�2y>�h�?�o�?E�g=���=���=���Y�����᣽�-.�<=�?�#?!@T?R��?��=?�H#?Z>11�"C���^�����֋?,?2��>[����ʾbᨿ��3�"�?^X?�/a�_���1)���¾cսY�>�U/�w ~�9���*�C����$������?���?�#@�2�6����Ę��d��!�C?��>�L�>+�>��)���g�"��L;>�v�>� R?�d�>`sI?MUq?T-m?�uE>��@�wt������j� �}b>�bM?�u?Yg�?�j}?�X�>L��=C���ξ����e�Y���m�5>�<1x1>]�>�G�>��y>���=	F��K�\J>��v/>�:>l�>'�>;��>�d�=9�I��"H?'��>c达ED��t��M���J��yu?)�?��*?�)=h�"=D�ǧ�����>�(�?;x�?�)?�JW��.�='q�e����s�F��>��>���>Q��=y�:=�>�l�>�g�>%=�b�^P8��H���?`;F?`��=�ǿ��q�(Ut��Ù�/�
<ҟ���mg��ᒽ
�R��K�=m���-#�·��S}]����9���>����G��u�u�# ?��=���=�:�=���<J�o�<~$s=:O�<uR=�i��	�<�D2�Dt�����Bf����<>�Q=�e�9��|��?�4�?��?��B?�s2=�L�=�ڽ��Y>�i-?\fh>�4��/����Q�u�J�~�¾]3Q�p����F�( ��i8�>�ʶ;�ڽ�$�a�-<N�'��-�>��*>K��<�E���̼0u�=p�>�%�<��j=AVn=�Č>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��N>22�=�M�H�-�/U�?06���p��_#?��9�,ƾ���>�Z�=��ɾ��̾�E8���E>|�=@=$���]�N��=���jm=c*l=G�>��X>��=�����C�=�}=���=�gH>ק�%;���WY���=�Y�=�y>��'>���>|?<-?zi?�>
�x����x���B��>�Q�=���>C�=fY>�:�>�W2?��8?��K?'T�>�ɩ<9'�>�y�>��,��Ru��O澺P��[I=K3�?&��?�޲>-�9<��B���v�@�����?��:?�Z�>�ύ>����ֿU<"��P1����S2��"��`S�#�<B�=1(�Vp���Z=g}�>f_�>
�>�$q>\_>�mb>���>"��=�r������;SRJ�UG�:�ZW>��=��W=��q��C�=�U�<�#;̰~<���;�ц=/=���x��=s �>�p=͍�>��=��̾��>�m��u9X���8=㾬�Q*�+�U�]�x�p,�"O�.�+>���=o��j���ޞ�>`_m>�%>`ֽ?�i?��:>���!��x������
��§u=��=��{�b@�h�^�p&G��m̾���>���>��>Wm>��+��0?�jWu=���/T5�s��>#X�����1�%q�O,��퟿��h��z���D?(>��bH�=�)~?�I?�ڏ?�m�>B���a�ؾ��/>A����4=2��sq��'����?��&?8��>G0��D�`��^y��E>A@ھ�/��롿��F��A>^�\���H>O���>Ӿ��M�Ɔ}��I��;'4��듾큩>WgP?��?���WK�c�m��־ۋϽg�?�n?���>b��>��>s־�P�ʾ�N��6<>�z?�?y+�?r�>D=�=ڭ����>A�?�j�?̳�?~�r?��=�r~�>r��;9�>5Օ�+8�=�>>���=3�=Y�?#R
?c�	?�4����	�ܸ��	�_�#��<�T�= .�>S��>:�n>~8�=��_=p�=��]>�8�>4)�>�a>Ť>���>�/��r�	�"?�>�|>�a1?ʃ�>i痼����.(�;����6�SO(�5FĽ��ｈF)= ��;s5�<�����>��i��?UK>���5e?�@딽n�|>�v>�#����>F�G>L�>h�>��>2@#><�>��>�8��>J��$�|�?�nV�2�۾߿�>QL���2�y,��t��}]��緾��|_h��ӂ�<�*�=<�?"UȽ-�g�FQ.�E���j?<��>��4?IL��4���n>���>��>�H�������r���޾.�?c�?p�]>N��>=T?b!?��9�D�*�DDU��=|��A���f���Y������}���[����`?��v?�v:?%N<�V>��?����a���u�>�2��A�ZmG=���>�P����[�(;)�����役�`>�m?��?5?�WQ�c�m�k-'>ճ:?�1?�Nt?��1?��;?����$?~3>�C?�n?\I5?t�.?R�
? 2>���= ����'=S8��(g�ѽf�ʽ���3=�[{=�M����<ܢ=��<����ټ�;���#�<	:=��=�$�= ė>aVa?^�?O�>�Q@?�^���A� a���h ?U�k<~�h������e��M��<-#S?�c�?��V?*%|>A�S�T����g>)ٓ>��/>���>��>3�$��@�P�=��=�/>�"=u+�<���,��D~�m/;�>h�>�@�>�	����)>��/�wh��O��=O�ͽ�ڭ������!���%�,��㾒>�w+?�?�vh=�疾�!!=h�n�p�@?��Q?��8?�1�?HW{�)/��&N���\��¯��+Z>�Eս+ט�봑��S���1�<>��K�zР��db>���j޾��n�J����qL=݁�E�U={�*�վ&'����=k:
>[����� ����Ī��#J?��j="\��n�U��n��9>kǘ>�خ>�`:�!Jv�W�@��Ƭ�yY�=.��>�
;>�������gG�Y)�m�>�-3?�BJ?��?W���Y�d�X�P��G��þ���� ?=j�>f��>��>�y7>��s������D�p�?��>���>\����=�Ȯ`�E����b<�H}>0:�>X>�P�>�(?�_?�Bi?�?���>�]>���貾��?"fv?{0
>��6���<��%0�I$8��>V��>���Y�0>ϕ�>��
?jM?>\?:�?�)��9�>�x�>	�>��K�iִ��U�=�GQ?U�?w�o?�9�?��>JHW��V����Rf>w�U>j�?Q� ?E� ?4��>���>Z���?�=��>�	c?�0�?�o?�~�=��?492>y��>D��=��>M��>�?�WO?*�s?��J?đ�>'��<�1���8��xBs��P���;��H<M�y=���4t��X�C��<���;mj��;�����S�D�K��U��;k��>$�@>{����>xk����MЧ=!�#>*��ƈȾ!ϔ<�K	>���=�?�%�>ʍ���[����>xȫ>
��*�Y?MR�>p�7?c��>�L��6�=������*}=��=?���>�(#�!~�یS��H�L�l?��M?Y������K�b?��]?4h��=��þs�b����b�O?9�
?(�G���>��~?_�q?d��>��e�%:n�'���Cb���j�)Ѷ=]r�>LX�O�d�p?�>r�7?�N�>&�b>z%�=^u۾�w��q��c?��?�?���?+*>��n�R4࿨���rˑ���]?�@�>�3���"?�|"�hrϾ�7��я���ᾴ���IЫ�:���B���#?$��y��!ԽH��=p8?�s?B�q?}�_?� ���c�)4^�65���'V��u�w��
�E��eD�0�C��,o��5���������G=hqy�y<�L��?TO(?%H8�f�>�ȓ��.��UҾ5�">-Ɣ�1��r=�=+儽�zV=��=lV�i&8������?gd�>J&�>5E6?�~T�ac@�^ 9�	�3��I뾟�>�>33�>J�>�T="��ĽHPɾ:�c��iн,(v>mbc?gK?i�n?j'�)<1�b����!�L2�cK����B>0a>���>�WW����53&�A=>���r�_���q����	�33�=��2?a�>�>m=�?4�?�k	�H쮾j�w��}1���<��>�h?=%�>X0�>�ҽ� �Os�>hpm?���>)!�>V炾��!�9�{��8ϽK��>e��>��>�?`>�80�|/[�*}�����p)6��>�g?5�����V����>��P?�D�;�<��>Z\��W3!�~���7'�Ċ>U@?;ʉ=�(>,ž�
��y�1��_?y?�YW� �9��q�jdA?�<?+BP���?���>{�[��
�_�>���?���?҇�>u���X�>w��>�Z<_���; T<�'�>�-��B�>'�Z>m��A�w>�B��}=&�C=$�����3Ƽy0[����O�x>3�!>���W�D�4���m����۾����7��Q�`��2����z���P5������9�3���ڛV���S;����@��K�?/��? <���訾Rʌ� Mw�A�����>Syu�K�H�� ���LM�l񨾢ھeƾ�>)��|V�c�X��qE�H�'?����ٽǿ��;ܾ'! ?�A ?1�y?��R�"�Œ8��� >wC�<�'��9�뾬�����οߦ����^?���>���/��l��>ǥ�>�X>�Hq>����螾�.�<��?4�-?;��>v�r��ɿY���V��<���?�@��G?sGr�ܦ ���>>U�>�@?�,�<�u8�u�$��D˼��i?�I�?pƒ?�:ݾ�"]����>F.�?��"�GC��A�=��0�r�,>В�=V��"�>k��>b�2��ڽ��ļ����Լp>y��~_�)S���������@�0*�=)Մ?�z\�Zf���/��T��{U>��T?�*�>�;�=��,?o7H�X}Ͽ�\��*a?�0�?Ѧ�?��(?�ڿ�ٚ>l�ܾv�M?-D6?���>�d&���t�ۅ�=�8ἐw��I���&V�S��=4��>2�>��,����O�`H�����=��-���j1��"�{�<}Z��Lٽ��+��8�<B<�`��#~F�Ih6�a��;]�>XvV>�\G>�q$>h�F>Sa?�r?��>�$�=ߌo����	�߾M:=��y��N��y����P��+��=7�|�ܾ��)C-�v��A��"K�-�=�U�A��k����ƃ�dHU���S?�9�>�E��B�R�������i��-=�< Yмh��`�-�-����?u�&?Jyk��b�BG��ɔ<x��W�A?;54�e���GǾ�>HT�=&�?>Tb�>�u>�%��$�(~.�vs0?�K?5f��@��3*>�� �Q�= �+?�y?)LY<�*�>/3%?+�*��+��[>�3>n��>���>�	>���hM۽K�?D�T?���j͜�3ސ>�F��i�z�BBa=n>FC5����.L[>��<����{U�*���ֺ<�'W?둍>��)�<��V{��e���">=�x?W�??�>Zkk?n�B?1P�<I����S��"��(w=��W?~#i?Ĳ>tʁ�:�Ͼdj��ִ5?W�e?��N>!h�a��o�.��O�<#?��n?�X?e���z}�]��p��-b6?��v?s^�ns�����5�V��=�>�[�>���>��9��k�>"�>?�#��G�������Y4�Þ?��@w��?%�;<��;��=�;?~\�>ޫO��>ƾ{z������/�q=�"�>����zev����R,�Y�8?͠�?���>�������[��=�����G�?f�?͍��.g<����Cl����k��<N8�=)���!�B����7�/�ƾ��
��������9��>DP@�W� ��>�7�p/�[Ͽ����R)оyQq���?�j�>�ǽ�
��Uyj�7&u���G��H��������>��>K+����\�W�M�q�ʽ�5?���<�R�=w����!��"/��P�b=��>���>Hٕ>G&������?�����ǿp����%:g?�\�?j�W??��>�'��s�j�<�� 	G>y�Q?��a?�`B?�IQ� _Q��⿽�j?e`��iU`�6�4��HE��U>`#3?I@�>M�-�?�|=�>Ƌ�>Rj>#/��Ŀ�ض�9������?X��?�o꾟��>��?-s+?�i��7��)Z����*�+��;A?02>�����!�0=��В�'�
?w}0?m{��-�r<X??�\���q��'<�	|���W�>f9�r(-�+P����I�q�i��J��`v��?�+�?��?M�a���'?sν>�`��~jԾ,=���>���>��\>ֽ_>>o����2��)>!�?�\�?_?W�cΥ���>�p?t�>.	�?*N�=��>���=Nޱ��Y�g#>ô�=B���?MM?��>5E�=ep9��/�1�E�)�Q�����C�U2�>�9b?*�L?��b>[h���3��d!�{DͽL-/�`(���?��*��x��S2>�h=>�W>�	F��Ӿ��?Op�9�ؿj�� p'��54?+��>�?����t�=���;_?az�>�6��+���%���B�]��?�G�?B�?��׾�S̼>=�>�I�>6�Խ����o�����7>=�B?;��D��x�o�Z�>���?
�@�ծ?vi��	?C�@O��Yn~��z�1B7�Gr�=��7?���z>���>��=qsv����c�s�x��>�>�?_v�?���>��l?�{o���B�-1==R�>Ŕk?�t?�Tc���򾉙B>{�? ����>�'f?��
@v@�^?_袿��ε��ϵ��ߥ��=�Y����A<���p��=c�3>�3:&�������6�C>J�|>��,> �=��!>��;>�����s"����̛�����z����(��xν�6�O �����!������q�̽�Hk�?Ƚ9���f@�������=l�U?�R?p?L� ?�Mx�ֱ>r���4E=��#��̈́=�'�>c]2?�L?P�*?q��=㝝���d�S]��/:������ʓ�>�aI>�o�>\A�>��>\Х8��I>]?>v��>�>�'=��Ժ@=��N>�K�>���>\m�>0<>�k>mʴ� N��uh���w�kr̽@�?�N����J�/9��"�������C�=�x.?��>7���п^˭�(KH?i���J�Ab+��B>��0?8aW?O6>\����V��>^��B�h��>~ �� m��)�$Q>�&?B�f>cu>��3�Z28�԰P�y~��N�|>��5?)@���.9�ȹu��H�.AݾSM>���>#@�@]��󖿂�~���i�'{=Gs:?e?�̳�tf����t��\��UR>{\>H�=:ũ=AAM>O�b��ǽ!=H�p%.=�q�=�`^>�?� #>&�w=Wh�>.ɛ�]�>�=�>�#>�Z>΁9?s�$?�1����������4���|>^�>�o>ȥ�=a E���=�>�>�_>�8	����%���XG�Ec>����~zT��a��Ȃ=+A���h
>E��=G���y�-�M�=uz?0���DS�k�޾	�I�N�J?�? ?���=TV>=���@��ҾJ�?��	@���?Zv��\�N�,?�j�?�֗��#W=�v�>a_�>�ž+/E�BM?^	P<+7��3����U9�?���?��߁�Ont�;u�=��!?:�Ծ���>ˌN�M���j����`��!0<�i�>N=>?P뾂5}��}��?�_?.8��e3��ެ��E�]�J��>7n�?^��?d@��������
���>i��?"�N?5��;����@E�]?��Q?���?w��>�I���P���&?�"�?�K&?�B>��?.%t?���>�Y%�1�+��l������S�I=�_O�*ԋ>���=��žR�G���o����h�I����\>Eu=��>�{�\��\X�=�hX�����6c����>�o>��A>#�>ƌ�>[~�>ڢ�>�=8��!�'��w�K?���?���2n�kL�<���=Ѳ^��&?~I4?(h[���ϾKը>κ\?u?�[?d�>>��;>��*迿~��A��<2�K>4�>4H�>�#���FK>��Ծ(4D�rp�>�ϗ>����?ھ�,���O��;B�>�e!?y��>Ӯ=љ ?��#?Ζj>3*�>�`E��9����E����>o��>�H?s�~?��?�ӹ��Y3�l���桿�[��:N>��x?V?�ɕ>9���փ��S|E�|8I�5���㛂?ftg?�Q�9?2�?A�??��A?�%f>r���ؾ������>�?�l��l0�9�-�}�G��	?.X
?r��>R���j��X�ɑ(�/v���%?��f?��?����qI�n?���#=^�;dk8��?;����d>I�>>��ʽ?�H>W<3><<�?���C!�C��<e��=�/�>d��=}U:�?2���<,?��G�ރ���="�r��xD���>�DL>����^?�l=���{����x��9U�� �?��?�i�?;����h��$=?��?�?!&�>{L���޾W��"Xw��xx�+x���>U��>^�l�N徨���"���F���Ž�0�?<2�>�?NT?�R#>D��>}�ؾ�M�	c��j徥�(�j��bE��e�d�˾��~���G�.� �ᘮ�m���O>˲�_�>g�&?���>��=#X>�O�=���>��g><�>H�m>T�W>��3>Ռ�=�*w��QzK?ؾJ>����H�S�F�7�@?[?ܖ?Bh�>������/�>��5?]�?��?p㓿��5���]?$f�>��6����>����d�=�7�>��Wq)��M�>�+���Hk���>���%hN������!?�6�>��&�ٽ�\=���""o=bN�?a�(?/�)�o�Q���o�r�W��S�:���4h��l����$�:�p��쏿�]���#����(�W�*=d�*?��?t��v����E#k��?��\f>���>�%�>�ݾ>/wI>��	���1��^�YL'������N�>CX{?��>B�I?ݯ<?�%P?a�L?ʕ�>�ե>!/���[�>�ݕ;�>B4�>��8?�-?#�.?��?�+?'Fe>:�����־�W?d?m(?%?LA?p���%½6mn�ui�@�w�q���֨k=��<�tٽؘj�(QP=��R>�f?z��K8�h���c>&�7?d��>�A�>Z����5���G�<�*�>��
?>�>q��j�q��`��G�>~��?���G�=j�)>F��=k���V�#�0Z�=|�̼� �=~���פ?���<�^�=S�=x85�l :9�9MC�;^,�<P�>� ?��>�N�>��� �S����=^�X>A�R>��>�Uپ;{���#����g�2y>�h�?�o�?E�g=���=���=���Y�����᣽�-.�<=�?�#?!@T?R��?��=?�H#?Z>11�"C���^�����֋?,?2��>[����ʾbᨿ��3�"�?^X?�/a�_���1)���¾cսY�>�U/�w ~�9���*�C����$������?���?�#@�2�6����Ę��d��!�C?��>�L�>+�>��)���g�"��L;>�v�>� R?�d�>`sI?MUq?T-m?�uE>��@�wt������j� �}b>�bM?�u?Yg�?�j}?�X�>L��=C���ξ����e�Y���m�5>�<1x1>]�>�G�>��y>���=	F��K�\J>��v/>�:>l�>'�>;��>�d�=9�I��"H?'��>c达ED��t��M���J��yu?)�?��*?�)=h�"=D�ǧ�����>�(�?;x�?�)?�JW��.�='q�e����s�F��>��>���>Q��=y�:=�>�l�>�g�>%=�b�^P8��H���?`;F?`��=�ǿ��q�(Ut��Ù�/�
<ҟ���mg��ᒽ
�R��K�=m���-#�·��S}]����9���>����G��u�u�# ?��=���=�:�=���<J�o�<~$s=:O�<uR=�i��	�<�D2�Dt�����Bf����<>�Q=�e�9��|��?�4�?��?��B?�s2=�L�=�ڽ��Y>�i-?\fh>�4��/����Q�u�J�~�¾]3Q�p����F�( ��i8�>�ʶ;�ڽ�$�a�-<N�'��-�>��*>K��<�E���̼0u�=p�>�%�<��j=AVn=�Č>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��N>22�=�M�H�-�/U�?06���p��_#?��9�,ƾ���>�Z�=��ɾ��̾�E8���E>|�=@=$���]�N��=���jm=c*l=G�>��X>��=�����C�=�}=���=�gH>ק�%;���WY���=�Y�=�y>��'>���>|?<-?zi?�>
�x����x���B��>�Q�=���>C�=fY>�:�>�W2?��8?��K?'T�>�ɩ<9'�>�y�>��,��Ru��O澺P��[I=K3�?&��?�޲>-�9<��B���v�@�����?��:?�Z�>�ύ>����ֿU<"��P1����S2��"��`S�#�<B�=1(�Vp���Z=g}�>f_�>
�>�$q>\_>�mb>���>"��=�r������;SRJ�UG�:�ZW>��=��W=��q��C�=�U�<�#;̰~<���;�ц=/=���x��=s �>�p=͍�>��=��̾��>�m��u9X���8=㾬�Q*�+�U�]�x�p,�"O�.�+>���=o��j���ޞ�>`_m>�%>`ֽ?�i?��:>���!��x������
��§u=��=��{�b@�h�^�p&G��m̾���>���>��>Wm>��+��0?�jWu=���/T5�s��>#X�����1�%q�O,��퟿��h��z���D?(>��bH�=�)~?�I?�ڏ?�m�>B���a�ؾ��/>A����4=2��sq��'����?��&?8��>G0��D�`��^y��E>A@ھ�/��롿��F��A>^�\���H>O���>Ӿ��M�Ɔ}��I��;'4��듾큩>WgP?��?���WK�c�m��־ۋϽg�?�n?���>b��>��>s־�P�ʾ�N��6<>�z?�?y+�?r�>D=�=ڭ����>A�?�j�?̳�?~�r?��=�r~�>r��;9�>5Օ�+8�=�>>���=3�=Y�?#R
?c�	?�4����	�ܸ��	�_�#��<�T�= .�>S��>:�n>~8�=��_=p�=��]>�8�>4)�>�a>Ť>���>�/��r�	�"?�>�|>�a1?ʃ�>i痼����.(�;����6�SO(�5FĽ��ｈF)= ��;s5�<�����>��i��?UK>���5e?�@딽n�|>�v>�#����>F�G>L�>h�>��>2@#><�>��>�8��>J��$�|�?�nV�2�۾߿�>QL���2�y,��t��}]��緾��|_h��ӂ�<�*�=<�?"UȽ-�g�FQ.�E���j?<��>��4?IL��4���n>���>��>�H�������r���޾.�?c�?p�]>N��>=T?b!?��9�D�*�DDU��=|��A���f���Y������}���[����`?��v?�v:?%N<�V>��?����a���u�>�2��A�ZmG=���>�P����[�(;)�����役�`>�m?��?5?�WQ�c�m�k-'>ճ:?�1?�Nt?��1?��;?����$?~3>�C?�n?\I5?t�.?R�
? 2>���= ����'=S8��(g�ѽf�ʽ���3=�[{=�M����<ܢ=��<����ټ�;���#�<	:=��=�$�= ė>aVa?^�?O�>�Q@?�^���A� a���h ?U�k<~�h������e��M��<-#S?�c�?��V?*%|>A�S�T����g>)ٓ>��/>���>��>3�$��@�P�=��=�/>�"=u+�<���,��D~�m/;�>h�>�@�>�	����)>��/�wh��O��=O�ͽ�ڭ������!���%�,��㾒>�w+?�?�vh=�疾�!!=h�n�p�@?��Q?��8?�1�?HW{�)/��&N���\��¯��+Z>�Eս+ט�봑��S���1�<>��K�p��ZΗ<�p�?���Z�\���C��8˅>�O9�\�|���#���۽��'�̱�>te�>�����1��0��V�¿�E?���=�g�����D�ZQ>���>�>��� ��U%/�� ���c�=��.>/�>7�5=�q����R�Rn�*��>�??�R?�8�?�B��c�Z��*��	{�r5">]7*?�9�>�1?���>Ƙ�=���!����Z�h�E�aK�>7;?Ry�,C@�J#�����*�@�p>�f ?�wL=%"?��j?,��>?�g?�q+?v�>6ڨ>q!��Swվ�#?��?!�=Z=�ɾd]-��U>�[ݾ>XGG?e����>w?2|#?�;?�"Z?6x(?�S�>$.���:�f��>X�>�gO������O�>��L?�߫>��e?��}?��=b�Z�̾Ј^��\�|>	�[?�?	��>m��>V��>����Bf!>"]?��q?>*z?�l|?���<�28?�cۼ�?�Ks��#>�J#?��?�`?�v?��-?��>:��<d���+�Kּ�R�<��<�V=uˌ=�P���&�pR.�L۠={D �P��D��1�����Y�=s0 =���>�et>a����70>[þ-����iA>*G��/����ɋ��h8�{ִ=]z�>u�?�x�>��#����=.��><�>#��	�'?�[?�?�h8�	b��۾�I���>��A?G��=h�k�0m���v��Re=W�m?E^?3�W�� ��F�b?��]?lh��=���þo�b����X�O?0�
?;�G���>��~?j�q?D��>:�e�+:n�%���Cb���j��ж=_r�>LX�5�d��?�>t�7?�N�>g�b>�$�=�u۾�w�r��n?��?�?���?�**>}�n�O4�P�Ͼ����'D?���>^����',?D�(�>^۾n��� �t��澝Jվ/u����R�;�4���	��P�7��k>P�?Mt�?�M�?$�k?����\�VGa�$ΐ��^A�%}���;���I�{�S�t!*�Lc�|���D�b���`O+=+}����A� b�?�A'?�/��K�>ʶ��&��t̾ �B>�0�����)0�=�D���8C=�Z=l�h�|R-�3����F ?K{�>Z��>��;?�1[���>���0�.m7�'����!0>�\�>r	�>���>�n;�-��&��ʾ�!���mؽ�e�>Un\?�Y? um?x�E��J�F����D���m.��x�>��>���>P����1��+���Vs��Z��#����%�׏,���e?Y��CD6>�?O�(?���{7M�!�&��E����>N�?6f�?X��>��> � �= ���>Z�l?!�>���>rc��v� �ր|�y�ҽ_c�>I��>2�>�p>�C-��d\������Q����8�f��=�Dh?Rb��gb����>�R?���:yC<��>�Gt�`�!����)y!�>{�?��=�hA>��ľ�W��;{�WL���e)?��?�����@ �"]L>�!!?q��>�z�>�;�?L/�>�ߎ���ۼ	!?�P?A�P?��T?���>��ɻ�����=ƽ�D�S �=�j>3�>�{>K�#>�c�CS��N#�0=g�2=,I5��q*�qr�;~h
<Ks�s[�<��d>��ڿNM��ξ~��v�X�3�� v��W���U���V���ّ����%������I���Y�����O{��4�?���?VW��+���>�����v� ���>@����(������T�g����ھjե���#���V�4c�K g�X�??��H�L���ᬿCɾ�.?p�5?�?��(����K8� i�>�<۽� 8=�Y��]����3ֿ���;�i?��?{�龧qϾ�'�>,?3��>��>��g��{L�'	��;B	?�z?E9?G�Ľ��ѿ��ǿ>�.>���?�Y@�UA?�(�+1��T=}�>U�	??�?>��0��C��8��6��>��?J��?w%I=��W�WM�P7e?�<,�F���׻�D�=���=W�=n��e�J>���>r�1�@��rڽ�4>� �>��$��R�k�^�q{�<]>'�ս>��5Մ?+{\��f���/��T��U>��T?�*�>V:�=��,?X7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=}6�ꉤ�z���&V�|��=[��>b�>,������O��I��V��=�P ��ſ�����Z;uqI�O%�c��:ۑԼwG������B_��1���=sy[>鷐>O��>��>��>ݜX?�,t?� �>�=s`���hҾj1�Ro=�#��3��=坷�J^n�z޸�.c޾9ٟ�����B�X8����� >���/=[�A�]����a�m"o��]F��p.?�T>ف̾�N��I=B�߾{���E[;?b���Ҿi�*��	w��&�?O�>?O���!
[���
��k���Q���O?�tO�Fy�#?����>�7�2=C��>oɆ=4��'�4�<�R�8'0?'?���y��8�(>����x=,�*?�?x�<{�>��"?�v&����^>Y�<>�6�>�&�>?�
>H=���Tݽ�4?��T?�e��桙����>|���D�x��|p=�U>�7��,��{�T>�ތ<�㌾�*�����W�<�W?G�>�Y*���` �������F=/�w?+?�l�>kAk?C?@��<�f���T��"��u=��W?Ui?`B>}��Ͼ����Z�5?�d?��K>k(i��辷/�-`���?n�n?Շ?g͚��_}��$��GS���5?��v?�r^��s�������V�=�>�\�>���>��9�sl�>�>?/#�vG������Y4��?m�@���?��;<,#����=�;?�\�>,�O��?ƾ{z��]���s�q=�"�>����Vev����TR,�,�8?Ҡ�?h��>���������>�+o����?���?������$=�����q�ZK��)¼TYC<yb轉�_��S��aA�+��,B��m��z�<���>:�@v�E���>�P�|ݿ��пɎ��X־�� v�1_�>KJ�>�Wp��1���:o�	�b���B��J�X���#C�>@�>S��������{��y;��p����>X�����>1�S�������6<x�>���>��>`������ę?Q���<οu�����%�X?Ug�?sl�?�a?+9< �v��u{����)G?�s?FZ?�	&�C5]�5@7���x?�-���#���FM��$6��;�>d?��>Hv9�l�>�`>͆?B�{>�sP�� ���Ş�����C��?	��?����?��?e�@?�:��S��nei�~c�c>��Q?��u>��Ⱦ�f)9�'>��y�?#?����]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�#�>��?xX�=a�>u�=Pﰾ��,��j#>?�=�?�!�?�M?gN�>�X�=��8��/�[F�FR�-"��C���>x�a?Z�L?�Ob>����(2�N!��{ͽ�h1��A��`@�[�,�9�߽�*5>��=>�>�D�Ӿ��5?(2��(ۿIM��D_����N?X'�>&?=��
	���[��;w?{��>���X2���h��� H����?�0�?@��>���B����>�S�>��X> ����������3��>OK?g�Z�gEX��끿h�=���?Q�	@��?��U��	?���P��Wa~����7�s��=��7?�0�"�z>���>��=�nv�޻��X�s����>�B�?�{�?��> �l?��o�N�B���1=2M�>˜k?�s?bTo���t�B>��?#������L��f?�
@u@_�^?*�׿�����I¾�u��@�>u�a>��8>�C��w�=�R&�^S{=4簽�$>�.�>�wi>�C�>I]�>��>$>>�����L%�e����ꊿ�<�7���-���;��!�H�޾̿�
���?���U�M����<��
�_��h��m�����>ذJ?D�K?��}?hf�>PS'>�q�@<�<'���Qd@=1�>20H?LDG?��"?���=��v�m\���t��'����s�	�>3�6>�ݼ>d�>K.�>r����`g>Y�2>�,�>8��=Ww�=�=�=�E=�	T>���>ר�>{m�>�!Q>Z��=T�䎯�Η���R���f����?]<��e9�I����cӽ�K�9魼��.?�*>� ��(ҿ� ��.T?@����1��b���o>��]?U?�p�>�n���= ~F>VϦ�$c)�̓�=̓�ё��&�@��ӣ>�Bk?��f>��t>t�3��h8��P��ư��c|>G66?��� �9�!�u���H�/�ݾ�qM>�Ѿ>��E�Tp�e����$��.i�z�{=�d:?�t?3߳�O���ڎu��-����Q>�?\>��=�J�=<bM>esd���ƽ"�G��-=	�=f�^>��?Z�> &=�@�>
������+�>šH>(�!>�=?�L%?������Ӽ����'L��lH>���>��>G�>f;6�@�w=��?P�>ˊ��Q%�H��<c����X>@ļ=�����ܽ��B=�O��g�=���<��%�]�+����<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿj��>�U��d���'��Wtu��c(=���>~H?������R��>�ظ
?T�?.��`��� ɿ��v�.��>��?��?��m��@��{�?����>`��?8Y?fjh>�P۾/Z�x�>J�@?\QR?�ö>���{�'�~??'�?���?69�>�V�?Ȁ?)�>%�a>1L쾭�����{#"=��>��D��r�3f ��nW�#q���A���d����y>��C=���>F+�=���W�=[נ�vE���'�R)P>Э�>O�>��?H�>ͺ�>��>QJ">1>�������D�K?���?@��A1n��'�<��=��^�.&?�J4?	[[�_�Ͼ�Ҩ>(�\?���?b[?7j�>����=���濿�|�����<��K>[/�>�J�>���zMK>=�Ծ,<D��p�>Η>�!��d?ھ1���U��hC�>#c!?���>��=�� ?��#?�j>(�>�`E�w9���E����>��>SI?��~?�?�Թ��Z3�����桿H�[��8N>W�x?�U?�ȕ>0������G�E�uDI�����E��?�sg? R�z?X2�?1�??1�A?40f>%���ؾ�����>��!?����A��2&��D��z?6?��>Lh��w�ս bϼC�����B�?�1\?eu&?M��a�+�¾��<�="��U8�W�;�9�Ӽ>V/>o��=ղ=�<>@��=�m��g6��V<�:�=�>l��=%7������-?J�B�V����t=nut��-C�0J�>�
;>��¾��c?��3���r��P��:���/�h���?qQ�?D��?�R����j�|>?��?��?�f�>�۴��������#c������b�9�>ɫ�>'v�;7G�l������h)��&�Ľ����a�>1Iw>��?�0?lQ]>NB�>�ތ���#�D���Xc�$���0(�|Z3�ю����2��`&=��ȾN�f��X�>khl��m�>Pp?r@=>� �>�^�>������>�K�=d�~>�>Grq>��<>�.�=}_7�v�޽�oQ?�!���g)�7������A?��c?" �>D%o�����z���c?�?A��?֥p>3�h��+�tt?���>*&���
?w9=%I组�<7^��2���u����^�>��ҽd�;���K��Ab��
?��?�����j̾��׽�T��e^�=b��?D>(?��&�CN���o��sY��P���;���t�����$��^s�e��������S��2�&�+�M=�,)?���?!��Y� 쥾�Jk��hB�<\Z>-��>�L�>�D�>��C>7��N-��^_�D$�N���%��>�,w?+�>�AW?�gJ?�U?�?D>�>~9�>���FV?��<f/�>Z�1>=+?���>
C?�<Q?oT?�����H�(���S��@0?�3?�?u�>���>v��Y��>sk��I����?V�c���� >�N�M����A�=��=�0�=��?��ܽ� K��G�r2�>dA4?�D�>C��>=���}䛾���=Q'�>q�?���>���Bn�)�
�`x�>z��?*�5��Q�<��Y>g�F=���b��<@ߍ=��O=�,=��^8�:�#<�ky=��}�BW�;��=�<䳆����9�t�>3�?���>�C�>�@��)� �Z���e�=�Y>BS>�>�Eپ�}���$��y�g��]y>�w�?�z�?e�f=��=���=�|��~U�����@������<�??J#?$XT?[��?z�=?Xj#?��>+�gM���^�������?�,?�W�>���D�ʾ�ݨ��Q3��?wV?�%a��Y�)��¾1'ԽG�>g/��1~�����S�C�v�	��`���ǟ�?���?�\B��6�mh辺Ϙ��A��2�C?�w�>��>��>N�)���g��3�m�:>rs�>n�Q?W&�>^0N?'y?�^?�(=>С6�*��˷��,[ �Cs9>~�=?�|?Z%�?Hlx?/��>v>ӽ�h��k��@�"���dg����L=�R>��>���>sH�>E��=/ɽP����?���=r\q>+�>g��>�_�>	�w>J�<��G?1�>��m7�vi��˹����=��
u?5��?:+?	� =�J�>�D������>��?��?�4)?�8S� �=ZԼ���^�s�C�>Ȼ>gn�> ��=��7=>�>���>�������7�0HD��
?dE?���=X���q�}|���s��S��<B��.־��=�0Q��cU>��;R���վ��$�A^�U�}�����l�a��ɾ�?k�>�]>܋=)�=�8���	=�X-=.f�,��hu��[�=��5�᷂=��1�(��9���	>��a��˾w�}?9;I?i�+?t�C?7�y>�;>��3�䙖>W~���@?�V>��P�{�����;�����A��#�ؾ�w׾	�c�(ɟ�CH>�cI�q�>W83>I�=oG�<o�=s=�Ɏ=�mQ�p=*�=XO�=�g�=��=��>VS>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>J7>wu>�S��_1�E1Z���a�^Y���!?u9;���̾��>��=,�ݾB�ƾ�'=�<5>�p^=_���y[����=q����bG=�b=�2�>rxD>��=�k���{�=�O=��=wSQ><ƻ5�H�� .��3=��=�a>d�$>���>��?�~.?��h?���>�t��̾�_Ⱦ%��>.P�=�s�>�=�d>ϲ�>��7?iz@?~/N?���>��=˺>�>u.�D�k�ɜ�(���j/�����?�?�C�>
�3<�7��x$�j�:�G���8?vR/?m ?b�>��x�*�Ʒ��pĽ�Y=o�=ܝF�"��@�j���V�S�t`>�ܼ>�R�>�o�>L��>��p>{c>[	�>V�Q>�9>�r9�����
�Ӽ�U>72g<� �=�e!����<��X����;�<fs=S��<��ӽTw���>W��>y4�:HҰ>\]�=�I����^>a�����C�y��=jƉ�"�1A�l�x��W:�R=c���>u�v>_=����.O?\	>���>��?��p?�P=�������mB���4M�)����&>��>������9���c�J�P���̾���>/�>�W4>/;>��#�-�7��*>��澉"0�l��>5Gg��p�<m���p��`��њ�ئ^���]=��M?�g��l�>�`?1V?��?�~�>4�꺾DhA>_������<n!�3 $�-["=nF?��?ú>d��w:�qH̾����޷>�@I��O���?�0����8ͷ��>������оD$3��g�������B��Lr�Q��>+�O?��?�:b��W��PUO�����'���q?�|g?7�>�J?�@?�$��z��r���v�=��n?���??=�?,>-	�=š���A�>	�?�h�?��?*�r?m�>�p�>��j�5�(>!�ν�W�=l>>(�=e��=}�?l?FV	?|��|:
�J������!j�K��<ŵ�=�>l�>�o>c<�=��|=�>l=��D>.��>⹌>z[k>���> ��>������澆&�>�B=�L�>̒,?��{>�r>J�r��u�>k.�/����њp�F1:��4t��X�=a��=���>s%��梠?���=���?���8�Y���>���>����>�]�=09��,8�>)w^>�QZ=��>���=��žS>�
�7T'��qH���N��Zž�f�>C����o۰��e��I���0��Qc��Ǆ���@��8<��?��׽�	s���+�h�Ƚ��?���>P9?(�v�F�D�!Y5>��>m��>f��,����;��`w�6��?5��?0=c>�>��W?��?�1��3�ZvZ���u�D&A��e�`�`��፿�����
��,��T�_?�x?GvA?f��<i:z>���?��%�Տ�-�>�/�d*;�<=�*�>!&��8�`�`�Ӿ��þ�+�}5F>a�o?#�?�T?�UV���$���>��9?�F?��z?��2?��A?"�˳-?`��=��?���>a�*?�,9?�D?�i>��4>[�#�:�=�'������g.���?*�;Hw�=5�=��ʼ���e5�8=I�<��/;�4μ������f=��e=o��=]��=���>�@^?E�>�Æ>?P6?�����6�A���;0?>cC=��{�UL��\U��X@��<
>`�l?v��?�`W?��c>��B��fC���#> �>76*>n�]>UI�>����q�B��p�=�>��>;g�=�Y������	�����¼<��>��>�3|>�����'>�{��B,z�B�d>��Q��ɺ�g�S���G���1�(�v��W�>��K?5�?���=0_�y(��tHf�n/)?Z^<?)NM?�?G�=��۾9�9�'�J��<���>�P�<�������9#����:��(�:J�s>�0���_̾5��=�'�I�Ѿ�.���Q������</-�����;4�$�g
�%�N���3>��>"���r��9z����I?��=�mo�#{u��ϑ� a!�3�>U��>0�$�`?���-Y�gHB�b�>  ?��n>˕�>Vھ�_>�ؐ
�W>�>r�6?r�g?I��?׸��[7���E�h���Ƒ��~AO>�?޵�=�? ?��T>�(�>����XS;�7`� �L��3�>~��>s� ��0L��.ʾAw(��c'��>K3?��=�m)?��?I��>�9�?�n$?�p#?�%�>��
<�'�J['?.�?���=B ý&��V{B��YZ��-?œG?�1�0n�>�d(?'?JX7?��e?�j;?d D>_c��(����>`�>�GS������>D�1?�_�>�Zo?�Z�?cxz��d5�+<��
�Ľ�8>Ӭ*<�1?�{?*?��>]a�>�ՙ�V�=z@�>zd?��?kqq?���=�?P>>}��>L�u=CB�>s��>#�?�XP?@Hs?u�E?���>
�< W��yE���8x�߷��;�;Y<�m=eN ���^�����}�<2!<����:���
�|�a�����s��<.X�>�t>�S��
�0>�ľ$����@>���:z��K	����9��9�=���>��?)R�>fk#���=o��>D�>���,(?��?�?�^;:�b��ھ1K��0�>��A?sx�=�l��t����u�^cg=��m?�~^?|�W����J�b?��]?Rh��=���þ/�b����Z�O? �
?-�G���>��~?c�q?/��>7�e�+:n�!���Cb���j��ж=ir�>_X�8�d��?�>q�7?�N�>U�b>%�=�u۾��w��q��j?{�?�?���?+*>��n�Y4�Y�վ��VS?j��>�^�d�)?�w=��E��������	$����ľ�>��󽾦4k��e�	
���C>?�|?2!�?X>?a�[:O��d��Ⴟ�GZ�k��m� �Vp1�	OE�-�>�w�l��h
���
�#����=B|���?�(:�?��(?��3����>_d������;9G>���~x ��;�=�G����T=�oK=�9g�3�.���@?�I�>W�>Đ<?��Z�y;>�91���6�^����[5>dt�>��>�j�>�<�-&����XȾ�J��F`ϽT�>o�^?�+X?��[?������Y��5�3�8���o�h�ő�=:M��~>zJ˾��콵�S� ;%���g�0E���ᄾ޽���^��tL?�.�̖�>F�?��?]˾8�r�y	r��8�z�?UiO>���?�`?���>	E����E���>��m?^��>��>�@���m!�ێ��ׄ���>�~�>a�>�u]>��T��Z�[�������\>��M�=2g?v���e�[��>tR?�K���<nޥ>Cb���'�8iﾺ��=Q>�?ݨ�=�aS>��ƾ���{y�y���()?��?Ag��O�&�TeY>�{?���>��>��?�
y>�1����$<�c?�b?�mL?� F?�I�>ّF=�䨽�۽� ��N=B�>;w�> 9�=��>�1�P���vJ%�Ry$=׃=��#��s���=]�����4��<�L=�y;>�;ۿQSK�e�ؾ����M��H
�	������3E��Ǽ����[���+y��
�e�'�$U��c�tt���o�s�?	��?(v���]��wә��x������5~�>ҍp��������T�i��4P޾���Q� ��P�^�i�}�e��'?]!�� %ƿ�䢿nOݾ�q?��?O{?��kt"�{e;�#>�s�<u���3l�򭛿z@пݐ��mG]?t��>ﾈ}����>H��>�Uk>m5z>��������ev<�d?6�0?|?�
����ʿz(��<�<`��?]�@�IA?	R(����V�W=�N�> �	?\)@>�0�Fv�Mg��d[�>۞?ӊ?�XI=F�W�i���We?�C<�F�������=�p�=�=�?���H>��>9���?�eܽ57>*/�>'b$����H�^����<�|]>S	׽�ړ�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��={|���A��T>�Ϟ��%1=��;cXڽ�)?��-��P�����̄������<��=F2>>
�>xe>��=�N?\�i?�b�>"�>�CR=#����߾i{�F#g��;9��n���&ּ����9�Ⱦ&\�����i$���"���߾�1��~��e�%������,侅���`�0�')>?�7>���0�k�>�=�ݾװ\���E=j�}*�+�;�����S�?S�S?�px�}O`���/������i�;?��Y��z���Z������a#��u �BW�>�|���	�|���B�Z^-?9`?��̾~��:>#� �kz@=
].?�}�>g�	<A��>��?I�x��
�.>�O*>@�>���>��	>�V�������?�Q?5��-g����>nH��"Sc�=/�=���=�H:��U/�`hP>J��<H���V{�����p2=.$W?;��>U�)�E��3������?=�ix?�C?�;�>�yk?e�B?n͢<�����T� 6�=�w=��W?�i?��>�U���Ͼ������5?>�e?
DM>?�h����.�ׂ���?\�n?O[?_P��B�}����J	��%6?U�?�YR�����d�%�#�[�↰>Ö6?��?� O���	> �K?�]�=�Y���Ͽ��6�V��?�v @l�@���=��f����<a
?N��>�9þ���!L���%����=/Y-?2j�C,����-�:O,�t?0�L?���>UO��%�u>�B}�"�?��?�j���$J=��� p��Y	�`��T�=�C�����6"����=�)�վ�����-<��>�@>�x��z�>�pG�T�ܿY�ѿ)������O��M?�p�>��򽝰���+p�<�n��0S�"�G�Fz}�#K�>B�>��������@�{��r;�~E��p�>x	���>D�S�("��t���7�5<��>@��>嶆>�8��o뽾�ę?`���>ο���q���X?Ng�?*o�?q?r\9<P�v�\�{�����-G?o�s?�Z?yq%��9]�J�7�j�j?La���S`��4�LE�=U>�*3?yB�>�-��}=B6>���>�3>)/���ĿdҶ�z���G��?���?�p����>���?mw+?/j�E7���l����*�0��JKA?��1>v���F�!�>=�{ܒ� �
?(o0?���'�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?E$�>5�?�K�=�a�>4y�=���,�]q#>��=H�>���?�M?K�>)I�== 9��/��VF��CR�5"���C���>��a?#�L?�Jb>���2�!��eͽ�V1�m=鼇V@�p�,�ס߽h&5>��=>�>��D��Ӿ۽;?���o�ɿ�o��#3���QD?�e�>f;?�������8i�{��?���>\�C����y�j�\*A�6Q�?],�?R?�����L"���M>(1�>ʫ>D��=p ���֍���=dt?I�o��C��6C��S��>���?��@	:�?<�B��T?���nR���Â�as���_��%@>�,C?����l�$>=W�>��1>��r�	Ͱ�r q��s�>���?��?�?�Ae?��n�5!?�g��=`:�>�3Z?�?�=⼧�����S>V?p�����b���a?
	@��@ �e?�I���.¿(Ǘ��O�e�(�Ez�=�^#>Q�7>�Y5��v>ۢ�=M��;��:\i>���>�hd>UŜ>�I=>2B�=cK�>�T~���&�����&��B#F�DR�ws �_6�KL���n��v8����?�V��H��Gi��Ϋ9S����1N�a�=]G>�M?��V?�Ov?�5�>5�	=���=D���m⏼���"�<�ln=�i@?+�1?  0?�$�<�V��?�f��ԅ��✾ny���m�>��{>`��>��>p��>2^���\>�5o>J�>Y��=��:< ��=���=GJO>�˞>X�>>L�>��9>��>�ײ�����g��W����̽c͢?�#���!M�|?���^������w�=�-?�W�=����?�Ͽ[��HiI?䋾����:�Ku�=��2?��T?��>޳�p�D�i2>1��[i��v�=@�
�: w��Z+�YW>[�?$�f>�t>̀3�iN8�־P��r��o:|>�&6?�涾d&9�k�u��H�)ݾK=M>�ξ>E�D�$a�����K��Li�^{=q:?�?Q!�������u�o���bR>J\>V�=�.�=KCM>�Jb��Fƽ��G��H.=о�=�^>5��>)sG>Zb�����>eнJ�#��>�o[>e��=�WK?]Q?������t��]ͨ�ny�=�>-<�>h!>!�����:�-$?R�`>�x<~W=���r�Ǿbd=�8�<�>���蕽�"��p��*h/>lX8�����oJ��`�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�H�>�pŽ���Fk��2�d�+B<~�>D8c?.��0}��6���?��?����1��_�οQ썿)�?���?�ݗ?'c�x�d�3�4�?=�?��d?F��>IA��_��{��><	g?G�^?V�>��4�x{��r?��?y͝?F�>�'�?9:}?�<>��>�2!���ƿ�����;~[=�j�=߆��p8���9��C�������S���1�줞>�� =R�>آ:�������C�|�����r�>��~>��=�`>�Ȇ>�>�E�>�f2�����V��"v����K?K��?i���.n����<��=߼^�-?�O4?�m]���Ͼ�ը>�\?�?�[?Tr�>���	9���⿿}��qҖ<��K>&4�>CY�>�؈�dK>��Ծ�ND�5f�>qȗ>�{���5ھ�%������L/�>�d!?
��>�=�� ?��#?$�j>h'�>�_E��8��Z�E����>���>�G?[�~?��?�ٹ��Z3����$硿q�[�97N>h�x?U?�ʕ>D������s�E��FI�^ �����?�sg?"M�S?1�?I�??�A?�)f>ʈ��ؾ�w�>��!?��~�A�[4&�r���?�I?���>"����ֽ��Ӽ����D��@�?!\?C.&?w��Oa�þ���<�#���P��<�7E�M�>��>.��3�=�?>f,�=�Sm��86�ǃh<���=}��>p��=�97�D]����??YPV�q;���1E����>�^��>�5>��о�Kx?&���f\��^���������?�H�?�3�?�8�<�za�(fB?�@�?�b+?~�>zj��`��X���n:�:�$=�$���j�?^�X>�<��G���n�������U�ٳ뽼A�>�U�>g"?��?��~>�d�>���o0��s�P�Ͼ*Ma����/�3��j7��G�a���ɡ�h���eϾ��G��m_>�������>� �>��>���>�>�Ľ��>AJe>�zg>�͜>G�I>�;t>b,>Yz��,��KR?I�����'����9���}3B?�pd?�0�>�%i������=?f��?�r�?a8v>�~h�?,+��n?P=�>���~q
?�?:=��1U�<�T��ټ�-������>U8׽' :��M�.mf�$j
?�/?-��H�̾�C׽ν��A�=Hփ?� ?����=���i���^�1�X�{ח�N�P��'��ӹ.��pp����� �������U �8��=�,#?�-�?��޾�K�(Ԩ�ٜm���T���>>���>���>m�>Ҁ>��	�g6$�PBd���"��[���H�>�Vp?3>Vp]?]C?GnU?CL*?���>���>�G��	�&?����AN�>Do�>7P:?�$@?�.M?{!?��<?,X�=�3��Ӄ���?�DF?�-/?D��>�?����V9L=��=�����2nǽ5a�ʭǽnz�E�ud�=�??�e���2=���'�w>�1?�j�>_�>j��!F���m�=�`�>�1	?��>X���Dm��|�A��>�+?�k鼸��<�1>W�=�#���h3���=�mt���=���<3�]��;n��=�Ά=��&���,�ת���;�8=lS�>��?@��>L�>����� ��f�E�=X>�!R>RL>(پ8M�����X	h��y>�b�?;U�?�e=���=+�=�(����F���+�����<�?<�#?(rT?���?�=?*'#?�K>V ��'���E��%�W�?u!,?��>�����ʾ��Ή3�ٝ?f[?�<a����;)��¾��Խ��>�[/�g/~����7D����l��5��?꿝?+A�N�6��x�ۿ���[��{�C?�!�>Y�>~�>M�)�r�g�s%��1;>��>gR?�!�>��O?*<{?S�[?��S>2i8�G$��]ʙ���7��">{�??���?��?B�x?,��>��>��)�8.ྴ���`��fQ�(ł�?X=��Y>dt�>��> �>�(�=�bǽLh��/?�8��=u�b>º�>㫥>l��>�Ow>QJ�<d�G?�>(?����v��.׃� P>��u?f��?�^+?��=,^� �E������n�>r�?�?�%*?�S�/��=(ռ[Ӷ��q��u�>��>�f�>
�=<�E=��>���>�a�>���J��n8�YN���?F?��=|Y��U�k��^
�/J����v>���yP��5?=���h,�=G�H��=oa�l�><@kU���@��ě��c޾�?��h5?�7�=��,>PK�;��q=媆����=�>�}�=�Հ<u����)=�û�S�<�H���<}�+�H��=S�t�o�ʾ�]}?��G?h`+?��C?��x>8*>g�+�l�>����41?G#U>^L�t����.>�G^��*����׾[N׾Άc�{���?�>(LE�i�>!
1>��=�)�<��=Ҷ|=!��=�m+�Yj=��=^�=�0�=ˑ�=i8>7!>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�@>3�9>�c����i�ٽ��F��(�a�!?k�=�4*�~��>��x=
�����;쫽��>+o�=��ҽB�R���V=�v@���Q=�ְ=)O>�Ь=#�>�Y�;��R>���=��y>�i>�e�^`x������-�=���=�4>�;a>���>��?Db0?]d?�ڸ>�`n�m�Ͼ�
���m�>S�=東>��=�XC>�۸>�08?�D?k�K?���>��=2(�>�e�>q�,��n�H\循h��r8�<?��?+�?�(�>[�V<�!?��}���=��oŽ��?�*1?#o?&�>;\����Y���!�¾�=u^�=�k���&�=���<��&�t�T�1�>I�>W]?���>�<�>;V�=	~t>�A�>��d>	�>��1�<Cn�<K ��N=Er)��U�=4�&�ɽ�jd���6�I[�����=Ȏ=M�;C0�lfb>"_�>�~�<! �>���=T�����1> ����~Z����>@֌�ğ9��:��o��D��7��h>�
�>!��<�吿��?�U���>�x�?o{?�������^���U+����!�e>F?>S��7�)�-�E�&�n������>ip�>�u�>xue>B�'��:�M~=��߾Y�7�4��>�ኾ�oE�I�	�w}o��=���џ� �e�̹<+�C?G�����>��p?�rK?���?�0�>jwŽ!�Ͼl�>袕�=����V���t�:?`"?�P�>.����RG��G̾8��~߷>N@I�
�O���Ű0����ͷ�+��>����	�о�$3��g������N�B�/Nr���>�O?`�?�:b��W���TO�=��W$��r?�|g?�>�J?�@?�$���x��r��H|�=��n?��?=�?�>B�=4���	�>!U	? ��?���?�ws?k ?�"��>,�;�!>��w�=�>,_�=v3�=��?�[
?��
?������	��J�ѥ���]����<gK�=2m�>Ox�>�r>�t�=�ih=TT�=��\>�c�>䨏>�xd>���>썉>O�;��?eq>%��>��/?��>i�_=jU��l�~=��O�}\N��N/�u�ν�u����:�|�;Ӛs=xR�����>KqĿ,��?�S>�� ��n?��掷�z�'>�XR>^�����>f�->4�s><��>��>��>��>5�&>����->KI��7J�I�<�{�p���þ���>�l���]��EC'�.����zJ���㾗�k����T8�:�;��ƕ?��;�9n�YD��;�&y4?9؟>�z-?1H��(D=S'�=���>���>���𔨿$������B�?Ȳ�?�<c><�>
�W?��?��1��3�6uZ�S�u��(A��e�L�`�=፿���>�
������_?7�x?�xA?~b�< :z>���?[�%��ԏ�|(�>�/��';�V4<=�*�>B+����`��Ӿ��þF8��DF>��o??$�?�X? RV�T��?P�>7�o?u_?�=z?WD?��K?4
��ke~?GP�>�R?�p�>�X2?�Q?�?b�>�;�>�����=����C7��B�;kHݽZ'<��p~=侉=)%}�2��=��=0>��
��n�>�>�<��f�$�R<KA7=>Y�>`�]?0��>�!�>�&7?���.@8������/?{0=����������a�ѕ>gk?"�?kZ?�c>�B���B�nh>^ˊ>W!)>�^>�<�>���X�G���=��>��>��="�J��΁��

��ː�t��< �>
��>�2|>�	���'>]s���#z���d>D�Q�κ�G�S�]�G���1�f�v��T�>��K?&�?)��=Y�D"���Ef��0)?ia<?�JM?b�?�$�=-�۾��9�h�J� R�~�>�w�<���Z����!����:�W�:F�s>K,���렾w8b>I���e޾�n��J�1�羻hM=V}��V=K���վR&���=�0
>	���2� �l���֪�+J?}�j=�d��pWU��k��g�>.Ø>ޮ>0�:��Fw��@����yR�=J��>��:>� ��&��VuG��5�Jen>�EC?|�]?*�?Y<��Z�U�a&���p��1����?_C�>�8?�Ԁ>C=M> +����	��Z���1��M�>jU?Hs �+/W��ͮ� ��W �k�U>X�>��=�T+?�~T?UV?ϴ\?��9?<?��>�f�;����BY%?���?1��=�Ͻ줾H,�#�9����>��?[�E�5ư>n�?&j@?�</?<`?P�	?��>pW�,7����>и�>�`K�멩�zu>u�]?R�>�G?�Iz?s�z>�=7���ؾ�X�=М[>�=�T+?o(?Kp ?�>IT�>�О��t�=�~�>��S?��?�Fv?͟|=� ?�#[>�X�>ST�=颧>e?a,'?�tS?|3e?A�>?%K?��4=�ƽ}�ѽ��D�?p˼+�<n>N<��n=�y ���ٻVh���9(%�rQ���<�fh���	��A�L�3�3_�>��s>s
����0> �ľ0O��A�@>s���wO���ڊ���:��ܷ=݆�>��?���>
Y#�E��=讼>3I�>	���6(?H�?�?1";��b�9�ھu�K���>;	B?���=��l�����`�u�X�g=\�m?0�^?��W�&��/�b?�]?�g�=�:�þp�b�߉���O?!�
?z�G�(�>��~?s�q?R��>��e��9n����Cb���j�3Ҷ=Zr�>VX�O�d�	?�>i�7?N�>t�b>�%�=�t۾��w��q���?i�?��?���?�+*>I�n�34�%k�n���c�F?%�>�N��vZ?P�������]O�� ����7뾵Q��/ז��;$gs��U=�2�꽡��=��?�Ǌ?��?�1B?ھ{Y�9AY������c���\�%�v�g�@�F�Y�P�Z�����&��1�<>8��A�%}�?��'?�0�8T�> %�����%�̾XB>W����ڛ=�׋�1 :=L�V=
�h���.�cd����?ﵻ>�j�>�[<?�`[��:>��1��8��G��:64>Tv�>��>\��>�=;�m-�@��ʾ�ׄ��νx�q>�
[?��K?	�g?�R�����s��&n����<L������MC=���>E��5D��bQ;���G���,8��0��uz �zxl=wM?Lb���>���?�h�>�����肾W��#>%8�>��s?���>?O�>�ڹ�Íd�m�>��m?e�>�:�>"��6����~���ͽA$�>><�>���>��j>�<)��l[�������/�:��V�=��i?ׂ��ke�b�>�NS?��ٻ�7d<�l�>:o��G �M���$�b6>M�?���=F�D>�þ��	��z��d���j*?b�?�3���&�G�o>tw&?��>RZ�>��?��>�Ⱥ��� ���?��c?��J?i�=?{�>��v<iMɽh����p(���\=�b�>x�~>�Z�=B>��#�Y�G����9=�ǃ=6;��m�����O�	�7���u}=��E>ݿ��P�Nݾ���4��c��d�~��9򼑋��O!�64ƾq�*���[�����)w������ǅ�����5�?�5�?��U��X���њ�Q�w����F�>��_�7;�������6�c�p�����:Mվ��/�NjM�![��|O�L�'?�����ǿ򰡿�:ܾ0! ?�A ?8�y?��7�"���8� � >2C�<-����뾭����ο@�����^?���>��/��m��>إ�>�X>�Hq>����螾U1�<��?5�-?��>Ўr�2�ɿc���g¤<���?0�@}A?�(���쾩V="��>'�	?��?>�S1��I������T�>n<�?��?�|M=u�W�8�	�-�e?}<��F���ݻ�=�;�=�E=\��"�J>�U�>����SA�)?ܽ!�4>,څ>k~"�!����^�a��<��]>2�ս;��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=����7ſ��%��e�C6=ku��$�g������������㿠��&]�p��[�V=��=�(->b��>	�W>�b<>�T?�+j?�K�>�>RV轏ł��*پg ����s�[��)~���wB��Μ��F��J�J���u���+���*�[���(���O�(��s��t��(4�Yw9?�*�=*(ƾ�/P�4�=���4���<=�듽�%ؾ��+��ju�o؍?�0"?�����MU�Z����߽��k��X?������û�|a">�M����<3?�>�J8=��徟�%��W�-v0?!]?����_��['*>�� ���=�+?E�?��Z<0'�>�L%?r�*��.�Ed[>Τ3>�ף> ��>�;	>E���U۽g�?��T?�������ܐ>c��r�z��a=�/>�<5����[>�o�<�󌾺V�K��^n�<�(W?s��>��)��|a��t��$Y==��x?��?!.�>n{k?��B?�դ<$h��~�S����aw=�W?2*i?��>����	о^���D�5?�e?��N>�bh���;�.�_U��$?�n?5_?n~��(w}����n���n6?��?��w������,��۸����>�:?ُ/?�2W����>؞u?~s*��奔\����_
���?�;	@��@I�����<�gE=�3�>�-?<���q���{�=�	�e
�>�o!?�3�a�m����Be5��?��C?��>m�~���*�=�턾-٪?U.�?�<���B</��g�i�����M��:p�)=j�����c���:�pjʾ���C��X.Q<��>�@���@u�>�.�H�ݿT˿;u��"�۾��R�?籓> �?ߋ�ރd�Ukj�¿O��tE���Q�SM�>3�>񲔽:�����{��q;��.����>��~�>l�S��$��њ��mT5<��>���>���>X(���潾Rř? c���?οy������
�X?h�?o�?p?�9<L�v�B�{�����,G?�s?�Z?�^%��:]��7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�#�>��?�t�=pb�>�b�=�&-��i#>2#�=�>��?�M?�L�>�V�=o�8��/�[F�
HR�$���C���>��a?��L?zJb>"���2�c!�vͽgc1�;�OT@���,���߽P*5>��=>B>��D�%Ӿi�?`p��ؿ�k����'�F14?c��>?��?�t�U���>_?�v�>�:�5,���$��WE�u��?F�?�?��׾�̼~�>]�>T�>��Խ�ԟ�:���_�7>$�B?���D���o�V�>��?.�@m֮?�i���?;��Z��%=��9"�����=y�{?��/�$�m=C�>�D�>���Ш���h��L?k��?s�?���>��u?�mZ�PUn��=��?�w?��/?|j�<x ����>ŵ\?�^�ϟ�������?-�	@aj@��?Vx��薴��ʇ�09c��Ϝ� ~>�l�yj>�<�O6<�,�=Kh���J�=�&s=�f�>T��>��>x\�=.!�=�ܘ=����E!�f���Q��.�/�b\a�p� �LK�=�89��݊�ls)��)��IR�H<��S�
��꽊B��(�3�����`��=ҫC?_TU?NBr?�m�>�o�<9�>�,�����<d���Î�cZ>��C?�5?d�"?|��������j��=���Z���H:���>R>f ?�'�>5�>x��p4>(��;�2�><�{>yN���T>J
(=�a>"��>s�>��>�B<>��>Aϴ��1��5�h��w��̽1�?����L�J��1��Q9������#i�=Kb.?�{>����>пi����2H?���o)��+���>a�0?�cW?�>����T�:>C����j��_>, ��l���)��%Q>il?0�f>�u>�3�gd8�9�P�i{��Fh|>@36?&궾�E9���u��H�`bݾuEM>�¾>�D�k������\vi�-�{==x:?2�?A3���᰾��u�B���QR>�6\>�Y=Nj�=XM>�Sc��ƽ�H��k.=���=x�^>�E?��+>9:�=�>�v��P�j�>pB>]Q,>t�??�"%?��&ʗ�m}�� .��v>,b�>��>UP>�+J���=[��>T�a>��l�������?�<�W>�}�?�_�k\v�9>x=}U��s��=�ړ=�� �S%=���%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ<��>�Z��c��5�����v����<S��>?I?������~��uH�qs?m�?������-�ȿh�v�м�>b�?
4�?fil����A�_0�>���?��X?�@r>�ݾp[�6Q�>��A?~_P?�>�>��6���?���?�Å?�>�"�? �?DeE>�m�=�뻿�����I�=�՗��:��MU����Ӿ, ��X�������	���"��1?,h�='4�>��d����!I>�̚��\�g��=���>b�;>�*>sG�>�?�q�=2X�>���BG�g��]Ge���K?ẏ?å���m���<��=��^�e�?m:4?�R��mϾ��>�#]?�΀?H[?�w�>9l�"�������� D�<Z�K>@��>���>+���OL>��Ծ92C����>�P�>�1��J�پa.��g���g8�>L!?�e�>Tۯ=ҙ ?Ŝ#?��j>�(�>,aE��9��e�E����>΢�>�H?��~?��?�Թ��Z3�����桿��[�:;N>��x?V?eʕ>[���胝�;hE�4BI�����b��?�tg?�S�)?<2�?�??H�A?q)f>���'ؾ������>��!?>���A��J&�G��?�I?z��>G��<�ս1+ּc���Y��&?|)\?�?&?���p*a���¾�g�<��"���T���;9kB�8�>�>i�����=k>���=�hm��=6���h<�>�=�>}��=$7��]��c�E?^D���	-��}��zM�sz�>��9>wȿ��f�? /3��F��ӣ�"���i��棋?��?�~�?f]P��r�1�E?�}?76?r��>���!��j=��_�цy��47�2䒼��?�Ax<�)�I������#֪�.��_�S�%��>��_>tW
?��>��U>���>@����4���f�Ǿ��i�6��z�=�/�>�&O��[t����0S�.�ʾ��\���>l�ֽ3C�>;�
?$�>疚>W}�>��ͽ���>��2>�Q�>���>�Z>��4>�>h)=�N���KR?����"�'��������h3B?�qd?M1�>Yi�:��������?���?Ts�?#=v>h��,+�~n?�>�>G��Uq
?�T:=�8�l;�<V��o��#3���1��>E׽� :��M�?nf�uj
?�/?'����̾�;׽?.���֘=��?Y/(?d�)��DO�Y8p��^W�3?P��@/��Ww�(���&�;�k�߮��vw��;E���j'��ʂ=��(?�v�?p;����������h�p�>��G>u��>�>��>@UB>B	�m4,�k[���#�Vv����>I�}?�a�>�R?�~3?iw;?��K?we?�b�>�9�u�?b־=�~�>�@�>�HO?SJ?�&=?��?��?Ճ�=�|z�/�徥gؾ I?��%?��)?��>D�>%-���ɶ=���=O��T ��,ʆ��
��_��9F��Wr�D^�=��q>�V?���ά8�����/�j>��7?X}�>%��>H��x0��"�<b�>�
?�E�>� ��}r��`��V�>���?8���{=��)>k��=����XѺ�U�=$������=��	�;��+<�{�=��=<t�f������:�!�;h�<�t�>6�?���>�C�>�@��/� �c��f�=�Y>:S>~>�Eپ�}���$��v�g��]y>�w�?�z�?һf=��=��=}���U�����H������<�?@J#?)XT?`��?{�=?^j#?ѵ>+�jM���^�������?w!,?��>�����ʾ��։3�۝?i[?�<a����;)�ߐ¾��Խұ>�[/�i/~����>D��텻���V��6��?�?LA�W�6��x�ۿ���[��{�C?"�>Y�>��>U�)�~�g�s%��1;>���>lR?~C�>N�O?�{?�k[?oxS>yT8���-����P-���!>�?? ��?��?�y?��>��>1)��>��\����3��pƂ�R�U=�Z>;+�>8�>��>s��=� ǽ�$���?�w�=�hc>_�>���>���>�kw>���<��G?=��>�]��6��U줾�Ń�F
=�'�u?䛐?ʑ+?�T=<���E��G���J�>ko�?���?4*?��S�C��=��ּ_ⶾ��q��%�>*۹>�1�>�Ǔ=�yF=�b>��>���>1)�a��q8�SQM���?�F?���=T�ſ
���ԨþJ�����=8l߾ϙ���=�0R����;1���T)=��پ�f�0�u�5����؛�R|X����yu�>�ׇ=&8>K��= ��=G^�4�3��ч<a�G>���<V�\��N�SZ7�ֺ��C��q;���3�Q=�����˾��}?�3I?��+?��C?ٿy>`2>B�3�@��>H����5?x�U>�
P������;�G���c����ؾ̅׾��c�Ծ���S>4�I���>�!3>�b�=S��<�2�=�Br=#�=*�G���=���=�Z�=q�=���=�>�x>�6w?a�������4Q��Y罐�:? 9�><}�=؁ƾq@?��>>�2��ȗ���b��-?���?U�?��?�ti��d�>8���㎽s�=)���%=2>q��=�2����>B�J>u���J��ǀ��w4�?��@v�??�ዿ��Ͽ�`/>�O�=�,�=��a�]�a�L���1��6~��?vKA������&�>�e��7ɾt�Ӿ�{����2><��=:��V�U� �X=Y]Խ. >���<�ƃ>V*>;D=�x���Q>��z>�4�>Ò����=�?<ܰ<s��=���>Ä>��>��?�`0?xUd?S*�>n��Ͼ�B���G�>��=:L�>��=��B>/��>X�7?��D? �K?A}�>ﰉ=��>(�>,��m�qk�hŧ���<D��?%͆?�Ѹ>�Q<(�A���Ka>��!Ž�w?T1?i?�ޞ>�B���7a&��^.�/ޚ�ng�8�+*=�/r��aS��@�N���㽉��=^B�>K��>;��>:�y>�!:>e�N>v%�>�<>��<���=�����<]ϕ��;�=z��n}�<T�μZ场Q�5��#-�fǥ��fx;��;�7X<��;�b�=�q�>��9��>,����V����>m$��Y�Y�J�=z��;B��8T��#��E��:1���U>��>>W�䥔�M?¨>a��>M4�?c��?-�`=mW�ܭ�=n��;�"�@ѻ�V!>+��=�^I�˷6� �Z��hU���Ǿ��>$ߎ>S�>��l>�,�"#?���w=��vb5�L�>�|��d��J)��9q�"@������ i���Һc�D?�F��P��="~?��I?B�?D��>��O�ؾ�90>�I���=���)q��h����?�'?n��>��u�D��ʾ�.����>-þdni������3���%>� پA�=@� �ߛ_��}&�p���ї���P����.�>�XH?���?�9E�����m�,�$�>�H?U�?&�>!��>�2?o��=A �y_����=d��?L��?]�?��j>螽=W˴�U�>�9	?���?��?�us?N�?����>�I�;� >�O��]��=�F>]�=��=bc?�r
?��
?�]��;�	�����!^�>�<�)�=��>�f�>@sr>��=��g=�:�=�\>Ӟ>cǏ>��d>`�>BT�>u��u}
�FG?�k>�"j>I�&?.L>燀=�۽����Z�j=(r]�}10�5;���O8�O-<�xS=d[�=I�k�w��>8���Z�?Z+d>��	�"�?Cbվ�1��̴>��?>m{�y9�>��>X��>!��>�h>a^
>dC�>[�Q>������9-�쾔",����<���TL��6�>1������P�'�-a<� y��k��d�
��ʇ�����Y$�X!����?nHZ<M�!�T�9�y�ھ��?���=84#?,Y��Z�?����<w��>
��>`cL��Ѭ�,!��������?���?>2c>��>]�W?L�?=�1�N3�cvZ��u��%A��e�=�`�䍿����~�
��+��%�_?i�x?hsA?=�<�:z>���?$�%� ֏�s(�>3/�1';�i�;=C�>� ��g�`���Ӿ̼þ$��@F>��o?��?�T?>1V�|��<c�>S4?O�K?��w?�K?�W?ؾnmz?8�>�8�>�b)>�S??�h?t�B?Ķ>�=$5��W�>�4
����z�ýs�ֻ����F��2�1>��G=�!�纽P�=\O=w:��O=G�= |Ȼ+��ؒ�<��=c��>�]?xL�>��>��7?����v8��Ǯ��+/?��9=*���(��QŢ����>1�j?���?�bZ?�`d>F�A�]C��>�Y�>�u&>O\>�d�>Qz�_�E�R�=PI>�S>h��=3WM�Wρ���	�V��� ��<�&>���>Y0|>(���'>�|���0z�7�d>o�Q��̺���S���G���1���v��Y�>�K?��?ӝ�=W_��,��mIf�F0)?�]<?�NM?��?&�=��۾��9���J��>���>^T�<��������#����:���:H�s> 2���ԡ��j`>j�� ߾��m���I�i���yQ=�E���M=H��Ӿ��}��K�=B�
>j����� ����ͪ��I?��q=�̤�~�V�X���C3>�N�>���>�<��:t���?��4���=E��>�8>�������F�?��J+�>�!?�Sf?J[�?:��C�@���*��q����)�>�X$?�`>9�?��>B��>�Q�B��J�_�A�^����>�$�>�+9��|B������Q 4�e�b>��?�|���u%?�-�?s�>��?&�3?"?N¬>OV=a�f��3?b�z?xm=�I!�ϐ���cJS�Q��>��?�VY��0�>()?d+?��2?��w? ^	?O�>�]�2f�o͘>���>z�S��~���8@>�`?��>�<2?eО?�W=��J��B���\�=��5>��z=Z�K?��?KK?���>���>㤡����=V��>
c?�0�?��o?�q�=��?_22>r��>��=-��>O��>w?�WO?[�s?q�J?��>F��<�<��1���<s���O��y�;�}H<��y=c���(t��M� ��<$��;Kp��a������D�����P�;;`�>�s>k	��e�0>p�ľ�D��>�@>����G��<݊���:�{�=T��>��?ޮ�>�O#���=9��>�I�>����4(?��?V?�L%;؟b�5�ھ$�K���>@B?��=��l�Ղ���u��g=��m?�^?ߙW�%��P�b?�]?!h��=�a�þ�b����W�O?E�
?W�G���>��~?u�q?`��>�e��9n����Cb�h�j��ж=kr�><X�+�d��?�>��7?-O�>z�b>�%�=Tu۾�w��q��|?m�?��?���?+*>b�n�84�_���P��t�N?���>��R��2?H�<��޾;�����V��uWǾ%rؾ�?���
��y@���lo������=�=�1?��o?,�~?�-?	�Ҿ|a+�z�_�}7���,k��!���>��M8� �A���T��O�����Z�4푾�,�=�{�[q?��?��)?#:�E�>�藾V���JѾ3eP>A����#�绬=�噽�pc=��=�l��8�sq��1?��>]i�>�;?�[[�0R>�@"/�ÿ5������->n)�>zJ�>�a�>��H<rD�hFཁ�ž) �������u>S%G?�w?�x�?�N��:j��Rfk���復�d��Lؼ���<�����>P��3sw�S/[�6sG���o�c���j���������=ޟ2?��<��>��?��>?i�O����n*�l�L���=}V�>�y�?�K�>���>�W��F��K�>��T?%�?�	�>˽Aq��������<o�r>hn>�
�>�1�=~��7K���N���f���F=���?�8�ح��0|�>�W?u@�	�="�a>��E>���g���ǝ�Y�>|�?j$��s�>������g�Q�'*ž��I?��J?F�оG�HZ̻GvL?�?C>N��?�o!>�=n���=�^)?�s?��N?e�E?J2�>}�	�����ŉ����̽�1��Y�>���>/A.>)b>F0V�Gy��|��D!2��IN=b�Ȼc��?,�����+˾<�P/�[SB>�nۿ��K���׾LS��d��A��I������kM����3淾>����v�j�W+�:�P�r�h�Lˎ���s��?ae�?Ǡ���^��^���<~��
���7�>�]t��bz�"T����� ���T���g����"��,P��Eg�]�b���'?�����ǿW���t;ܾL ?�@ ?�y?m��"��8�� >_N�<�F�����>�����οT�����^?l��>�	�+8�����>��>^�X>Lq>����랾�F�<��?v�-?��>�r�ەɿƊ���<��?�@o�A?��(�A�쾔�U=���>S�	?3,@>�z1��8�b����c�>�4�?���?
dN=�W������e?<�<��F���׻���=�Ĥ=m�=Q����J>V�>�\��PA��/ܽ�4>�څ>+�"������^�`�<�x]>�ս�,��5Մ?*{\��f���/��T��U>��T?�*�>[:�=��,?W7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?^D6?���>�d&��t����=_6�鉤�y���&V���=Z��>`�>Ă,������O��I��U��=����]ƿ�#�����=!��b������!�j�.蟾`i��{꽵�g=��=�P>1ۃ>��R>L�T>ujW?��j?���>#>W��υ�̾��/�A�����dS���g��"��Z�=�߾�
�Q-�P ��(Ǿ��W��"�b`��'��ש�x{p���L�J�<?O�:>�tž�m��#>L¾'C��S�C='���侜�8��w��nh?}	?k݂���R��- �V+����A�b?h����0پ�{޾t%E>Z�h��ZP��{�>m��=<澯�7��IU��|0?]v?≿�[<��ZB)>� ��=��+?ե?�nR<7��>�V%?t�)����-\>�3>9ˣ>���>ݙ	>!���۽Iy?��T?�	�����3�>襾��Bz��``=�>�^5�6V�Б[>�<ތ�`�S��v��4�<)W?'��>+�)����h������^==�x?R�?�)�>yk?��B?�L�<�_����S�C��jw=O�W?)i?8�>Jw���	о�����5?��e?%�N>�ih���龍�.�{U��"?f�n?0]?�����t}������]m6?�|�?�ބ�����B:���m�<߭>��?��,?�,>�;d�>��Y?�|p��.��������1�?�	@�M@��w��ɹ<�!��)�>f ?���C���<S ���C>���>���r��(���)=Y_,?Tn`?݄ ?�at�����|�=�͕��U�?k�?pT��"�i<���l�Ԩ��dÜ<!q�='i�s�#�-�h�7���ƾ��
������Y����>IV@ԗ����>�8��!�qWϿ���?о�Hq���?eQ�>(�Ƚ<�����j�'.u�4�G�\�H�
w���T�>e�W>@�Ͻ�7���
u������=��>��%=]8�>�s������ɍ�)}�=䠚>���>�ޘ>��fž��?���L�п/[��;I��"U?�=�?l6�?0�?Yׂ<Yyq�%h�ֳ2�5�1?#�b?�-Q?5hE��"b����%�j?�_��wU`���4�uHE��U>�"3?�B�>T�-�a�|=�>���>g>�#/�y�Ŀ�ٶ�@���Z��?��?�o���>r��?ts+?�i�8���[����*�m�+��<A?�2>���H�!�C0=�TҒ�¼
?V~0?{�f.�d�_?�a�N�p���-���ƽ�ۡ>q�0�6f\�K����sXe����@y����?D^�?i�?���� #�T6%?:�>,����8ǾF�<���>�(�>*N>�G_���u>����:�i	>���?�~�?@j?򕏿�����U>��}?�(�>��?��=�n�>��=����d�-�b`#>�%�==�>��?��M?�`�>&8�=��8� /�eWF��AR��7�C�� �>�a?Q�L?�>b>ȸ��81��!�F�ͽX1�P!鼲~@��.,�z�߽DF5>�=>�=>_E�Ӿ�X?����FϿV�����/�ex0?L">Ĥ
?C���ׂ������d?�o>l�#��0��%V�����⫪?~��?�?�s�w}����=1 �>��>]cm�F�}��	���Xl>f�J?1�f��c_�u]�>B�?�.	@�ɶ?�g�&?�i��1���~��;Bƾ������>��E?݅��Ĉ>���>g�>�1�������m����>���?���?-��>�l?��hJ��4>@��>AVW?F�?��h=�G��q�>�)?�]3��%��p?��@��@5��?t���!����$��Gh�������s�=/x=K�=>J$۽DZ�=�H<� J��>|=y��=���>
�l>��s>F� >|�	>��=��{��9�{������>xD�x$?��?����`�Qj��G<���;���˾�VM�a����L$�w���xz�1�u�'.�=��U?��Q?p?5s ?6�q�� >�����=��$�9��=�K�>R�2?��L?κ*?�h�=���w�d�������Q臾�>ZMJ>5L�>��>��>����I>K�>>t��>h >��#=�ï���=#:N>�4�>Y��>��>��3>�>�ʹ����ɸg��i|�6Iֽ�4�?�a����I�Ț��s����� �=�i.?9�>�֑�(	п�-���F?�������'��>\�/?H V?��>�i���tO���>?~�g��Y>Oq�wj���(�yUP>�?N6>�(H>+;���=��yK��qƾqB>�??����*�1����	�4���׾0�E>�2�>���<L��J��`���ꀾ=�	=�7?<?aV�`i��}���������c>l�^>�8=���=�S]>9�ܼ�(ҽ݀0�`BA=xY�=��R>ߚ?�*>R�=;a�>�,����P��;�>@�B>�`*>� @?�%?X��H���Q��5F/�{Gt>i�>�(�>�M>��H�	�=���>	�`>I���|��[��@�҃S>�V����`�\�m�v�o=�������=~{�=�� ��k=��3-=�~?���(䈿��e���lD?R+?^ �=E�F<��"�E ���H��G�?r�@m�?��	�ߢV�?�?�@�?��M��=}�>	׫>�ξ�L��?��Ž4Ǣ�ɔ	�/)#�iS�?��?��/�Zʋ�<l��6>�^%?��Ӿ&��>��!�غ��T⎿
q��==��>�J?���^l���ah�9?�q�>p� �A���>ʿ�'{�\�>܉�?�p�?}�d�#����C���>���?�nX?زl>���{�+��w�>R=<?Qx1?�E>z�3���a�%?��?�?�;4>ݮ�?�w?��>(�>Z�����C���3����s{`;���W���ޟ2��$����v���V�xD���?_i�=a��>��Ƚ3����y�=R���,Ģ�~<B�>�]�>!>>���>~�?P�>.l>��a�g�9
h��>@���K?X��?����n�D�<�J�=c^�� ?�^4?xud�,�Ͼ�>?�\?À?�[?�{�>����)��W���ˉ��䯖<��K>\F�>���>(���BL>d9վG�C�:F�>��>�C���ھ���6˲��,�>�S!?�[�>R��=T� ?q�#?��j>�(�>�^E��8��9�E����>)��>�G?=�~?��?�ӹ�Z3�����桿�[�V8N>^�x?LU?FǕ>'��� ���$�E�,@I�����ڜ�?�rg?�V彼?2�?�??��A?i/f>f���ؾ����Y�>�!?�t�Z�A�KQ&��&�ّ?ko?��>�Y��Y�սl Լ���^a��?�\?yK&?Q���!a���¾(K�<_!���`�1��;/DB���>�u>*��疴=	>k�=�*m�YP6��c<Q��=�e�>���=A*7�]���^;?�Jq������=�y��T�8#�>+��>Ev��8��?RC[=�rZ�
ɫ��N���E����?�'�?���?Y?���r�z�e?~�u?��?*�>h�۾P�H�C���T��Y#��4���=>Y;?�!=��:��࠿�.�� ������)`�h��>͎'>O�?���>��V=�7�>����\�%��`������|��?	�2�'��N��T��ԁ��������Q���҇�����>�]<x�>�,�>���=M�>b��>�'�<ZQ�>{#h>��2>{,�>�4�>h4�=�Л=U��=��-��LR?������'���辈����5B?xpd?s)�>ʾh�p���l����?Z��?0s�?�Nv>xh��(+�<k?�>�>M���p
?ID:=���$��<NJ��T��nN�������>�D׽�:��M�Tlf�6e
?W-?� ��
�̾9׽���G5s=J�?5~(?��(�s�P��zo�R�W��S���'�g�j��	���w%�[�p�.����"��S���'�W2=I+*?VH�?�}�������_j��!@��ac>�:�>�>���>��F>�	�I�0�}\]��@&�����w�>*�{?]�>��V?�>'?�]O?"2&?�s�>��>i��� �2?��+�=x�>���>_�Y?ͪE?m�<?H�?؎"?	�l=�k<�)��޾`�:?�H"?�O?��>^Z�>Ѯ����;M/�(�=V���NJ��	�="%�ɞ��f/<^�<�
�=�X?͔�"�8�����U k>Y�7?�~�> ��>���G-����<��>c�
?�G�>H  �}r��b�|U�>���?Z��~='�)>��=�v���.Ѻ`�=������=�>��Vw;�%p<��=��=ant�J������:��;}q�<�s�>��?@��>�B�>=���� �~��T�=rY>�S>�	>�Hپ~��A$��J�g��Yy>�v�?�y�?��f=]�=���=�{��U�����t���)��<��?�K#?�XT?M��?0�=?[j#?��>+��L��c^�������?m!,?��>[��E�ʾ�񨿪�3���?x[?�<a����;)�Ɛ¾}�Խ)�>�[/��/~����.D��ޅ����w��'��?�?�A��6�zx�ѿ��\����C?�!�>�X�>��>S�)��g�q%�2;>���>/R?3"�>��O?�?{?\�[?�MT>8��.��}Й��u4�"><@?U��?s�?�y?�x�>��>��)��ྙN����������DW=��Y>ꋒ>�*�>��>!��=��ǽ�6���?��]�=�b>��>_��>��>?}w>4�<�L?�3�>iɾZ{�����PJ�Q�=�)d?���?K&'?!�=d
���=�v�׾+�>�Q�?�r�?��"?��c��S>C��<�˾,������>IU�>�ř>��=R�4=P�>$�>�6�>�9"����^�7�"cT�?�	?�>?�վ=�տ����L¾�j���/�>۾2�O\�T� >y��,���;��!��>Z=�ٖ�dFO�cA��־�zԾ�{��]�>��#�xJ�>ց
>=��=O���z�=9�̽lc���$�7t=�4=��ܼ�7*;�R��, ��Ջ���=��=̺˾�$}?8�H?��+?��C?jx>�/>A3�"�>�����?�*T>�R�6L����<��ɨ�����:ؾ�t׾��c�+(��v�	>�I�o�>�3>��=��<���=�r=�=S���=a��=ϙ�=/�=���=�>��>�8w?�������� 5Q��7�`�:?)A�>���=��ƾ[@?{�>>�1��[����e�G)?8��?OW�?��?�wi��d�>��ڎ���=8�2>��=�2����>��J>k}��I��A����3�?��@V�??�ދ�˟Ͽ�`/>6�/>�>`S���.�(tU��g��jW�e�?f�:�=�Ǿ>Ή>��=��޾%�ž��=`72>k7e=���\��w�=5Ɉ�'IW=NFq=)�>�^D>�w�=9��K�=�O=���=��T>Õ��#�hX�ς=T��=^�c>W+>���>�:?M"?��R?� �>��½��9���/�>י�=�G�>G�;��d>�E?|4?T�O?�oR?
��>i��<���>��?H�N��F������q�Ҋ�=ن�?��g?���>eL=p�;��!�;��֯�nd?�� ?��>Y}2>�U�&�࿀p&�؉.�;��yJ�� 6= >q��P������`��"ܽ���=�+�>e��>��>��v>�7>�K>���>�>
>���<==�=J�d���<���~��=c��5��<>������˸ ��+�:R��K	d;b�d;�k<���;`��=�e�>���<x��>�)=-:Ͼ?�T>VоZ,M��bX>�ߡ�m�K���U�Xx���P�>:!���q>s�&>�x佧o��|4?���=��>Ju�?:nh?G�=ow]�Ygج�ÀA�[ɾ�c >/�'>�1U�A;�{�q���K��ؾ��>�> �>Xn>�,�j�>�3us=�`�ws5��s�>ٷ���V����^Kq������6 i�&�)�u�D?= ��@b�=6~?O�I?}�?���>-��I�ؾ��.>F����1=P��po���zd?��&?;��>�p���D�j�˾�����'�>��N���O��N��/*0��0߻�����>ֻ���ξ��2��e��A���@C�<u�0q�>�P?}��?0�b��_��`oO����+w���?�g?�>�N?�}?�������������=�,o?���?��?��>�J�=���l�>.	?���?4��?wts?St?�b`�>�4�;F!>UU��|�={�>���=���=�k?��
?T�
?�V����	��������]��M�<?��=���>�b�>��r>��=[�h=��=</\>���>ɏ>a�d>���>Wj�>{����L�qd?�L >���>*�?J�{>N�=Z-�y�=`6=�yr���S��1��C>��`	��-I<Y�=G(����>[���_�?��3>w����I?�t�ͯu�'��=�8�=ɹ�ڸ�>���=�#3>�e�>�%�>���=�ek>��P>�������<nھwC?��`1���\���Ӿeʟ>�K���ㆾ�P���<���_ۨ�K�
�;�m����y�+�l���b�?���;3N��JE�m솾��5?��>'c(?�o���X=�&!>�l�>4�`>{u(��1��ݝ��kž1�?Z��?2Q>���>dT[?�c?P9̽��j�V�`Gy�nsQ�Qk��$a������r��y��3G?�d?�4?�%R=H{>K0�?����V���9�>�%�'�T�����v�>_����䝾�b޾�3���׽u�->�h?�r?w|?9>н(f��9�>e�Z?�K?	M�?]�-?�M?�	��lCW?2�4����>tE�>�I?�EV?:�?pPH>5>;>�#���^$>l�ɽXe��?�<��ս�B㽤���s>�z7=�y5��b�=;��<��6��XY���=x��rS;=j{&<��w=+7>g��>6�]?RO�>[��>K�7?���x8�	Ѯ�t%/?s�9=L������͢����>e�j?*��?$`Z?E�d><�A�E	C��>�V�>lt&>&\>�a�>lc�ρE�� �=xQ>`>pߥ=�M��Ё���	�I���g��<�5>���>�9|>����'>Y~���z���d>T�Q�Qĺ���S�8�G���1��rv�]�>��K?��?��=�^�s���Hf��-)?V^<?tNM?��?�=#�۾��9���J�>=��>�+�<���]���H#����:���:��s>�1��~'��pZH>�3�T��[�S�0��R��=.�����<2�.���j����-�=J��=詿���#�+x���¬��?I?�p=�����!V��٤��k>�L�>��>�|3�@�f�%�:�^����e=���>��&>�������A�����7�>�Hc?|�Z?���?�H��4�����B�X�'��!��GC��@?��>O�	?;>֫�<Noܾ�$���q��0H��~�>h
?�CJ��G��Vپ�`�ML>���>�؎�G�A?�e�?z�'?e��?���>�l5?u
 ?��4<�k�� N&?��?eC=��L�GÀ��:�Q�I��=�>p�7?�H����>��T?�RI?3K*?�#?2�?IT>T$�&`��O�>\>J7l��ر�<�[>!�b?�k�>G�x?��?��>d����{�6ș>���>ю$>��-?�E?�I?�ΐ>I��>�b���A>8��>�88?��?�ц?>�<�?���=��?{��<�C�>W�+?D?�Z<?B_N?�5?�(?�Z�<;x��<P��|
3��2���x�<.�';)�\=<ˤ�	)�^1�O=ܗ�<�Η���!����<k�I���=��
=`�>�
t>@���0>��ľ7F����@>���;6���⊾6�:���=��>��?���>NT#����=G��>z?�>���/(?6�?� ?N�);��b�|�ھ)�K�f�><B?5�=�l�`�����u�wh= �m?0�^?Q�W�|����b?	^?uN��=���þ(�b����:�O?W�
?�H�e�>�?�q?{��>1f�,&n�w	��oEb��,k����=rj�>(e��e��P�>ң7?2@�>�Ec>���=�n۾�w�7J���3?���?y��?���?�h*>V�n�-*�I�������]?��>�[H"?U��g	ξ�J���{��"�㾿׭��Z���c��s��!Q%��_���ֽ��=�k?(�s?{Ts?��^?U���c�+ ]�.^~��qV�������#D��C�qQA�x.n�+�����V���yj`=�ww�Ö>����?t�%?�<�8��> ����2��ξ�B>Y��> �沌=I񤽎]=P�J=��`��,��(��)�?~�>�M�>�;?�o]�TL=�$�0���4������>�'�>�r�>�b�>���<�1�W�d�;c܀������h~>��d?�EC?p�z?�n��8���~�6q!��$W��ٻ���=k�<|��>�;��m(��@��aO�M�~�����-=���q�����=��8?r��>Z9�>�~�?d��>)¾d�٤=��7���A=��>��_?��?[�t>��(V3�;*�>��q?���>:�>�ؾ��վ�����=�꛼��>#X>���=�o1��	Z���xҧ��W�Pu𼷬�?�1o��iM��-�=��?�C-���ž��>��p=�D����/o5�I�2=9^�>]۽�,�>�]��������8B>��)?�?����,�uUW>k?�(�>��>#�?AZ�>�Ǿ�T=�i?�b?q�A?�-??$x�>���<3�����ҽx(�=
b�>��G>�9�=��	>M�5��1����<l�l=�y껉J��~�,<�!��:�U/=��X>5Zտ�O��`�����7�8�
�^�ɾ[�<ΐ������羚�`�=�j� �&�X�0�Ble��3q��Q�����Tw�?B8�?Q(g�s���n�e�;7����>6����佾~��t�q�/��v���h뾜T���[�>sz�F>{�"�'?����=�ǿ����3ܾ� ?�= ?D�y?Q���"�1�8��� >��<nh��`��N���h�ο����^?��>���&��x��>Y��>�X>�Dq>����垾ݕ<+�?C�-?Ѣ�>Z�r���ɿ���#פ<W��?t�@�vA?>�(�Y��,�T=C��>w�	?I�?>E1���r���$�> 9�?��?�pN=)�W��@	�Tme?#~ <*G�q�߻��=�q�=Ƣ=����J>v�>2���
A��Iܽ�\4>6��>&�!��x��[^��i�<�3]>P�ս�1���؄?�s\��%f���/�TC��<>�T?%;�>?�=��,?.H��}Ͽp�\�ba?�,�?��?��(?@���h��>#�ܾ!�M?�H6?��>p&��t���=�B�П����V����=���>�p>/�,�����O�峙�Ͷ�=5� �ߔƿ�m����L㎽�T�:�����_��!���Em�L���K����$p=Z>�yG>�ӂ>!IH>�4>��\?��t?Ͳ�>��=Oe��f���Ǣ��e=(M�����׶�t�n��e���m�������'t���� i���G?��n���7��獿+��}�z��1d���5?��I���ܾ��T���=�	Ѿ�Ӹ��P��r����3��RC�A�y���?g�+?~b�b}G��l��?��G��??��X�D��|��ox�>[����ｹ�V>>���/��.~�e0?��?2ο�ﰑ�"�'>XL ���=�a+?�(?>0<0�>ڬ%?]}%��]޽�,Z>�4>��>F��>s�>����۽7u?U?�� ��R���ʑ>P1��t�x��+`=��>q`7����2[>��<"-����k�����N�<�"W? ��>
�)�V�n��l����<=�x?z?��>p\k?��B?w�<zk��I�S���icw=��W?	i?a�>ob����Ͼ����D�5?�e?�N>Åh����3�.�BE�L?��n?�`?]��Xo}���"���o6?û�?�O�Y"���u�z<ik_>E?}�?�6�qq?�i#?�W�����~��I��)�?k�@H5�?�iI���(�I�m='��>E�?�tt��g��2���Ѿd�>Y׮>�����x���������3?0h?8��> ���;��V��=QⒾ�ܫ?g#�?|���+N<'����i�� ���<�Ɏ=D:��Y6��e�b9�!�ƾ�	��;���-ݼi܅>N@�Iҽ���>ţ?���noο\���CԾY��:?���>�Ž�D���j���s�sH�?GF�����wL�>D�>i���@�.�{��e;������>����$�>g�S��<��2�����0<,��>���>φ>��������?IH���;ο��������X?�S�?�m�?��?B;<�~v�{��i��G?y�s?�Z?��$�b]�^8�۾j?w]���T`��4��HE�YU>!3?bD�>��-�?�|=�>���>f>�#/�!�Ŀڶ��������?��?�o�"��>݀�?�t+?*j�s8���Z����*��,%��;A?�2>B�����!��/=�VВ�{�
?8}0?�~�t.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�j�>�X�?���=ӳ�>
[�=�~���#�r4 >���=�O��?p�M?�,�>���=]w8��o.���E�AR����W�C�9��>�db?/N?~f>�4����%��3!��-̽�\0��v˼tZD�HF��.�b8>d�<>��>��D�[�Ͼ��?>����׿\����^'�[*3?�i�>6?���m���p��<`?lB�>L�cD���2��(K�Q��?�2�?0�	?E�׾���w;>�F�>���>�½;���7e��u=>B�B?����E��L�p���>Ҋ�??�@�¯?g"h��?=�u���>ꗿS���g�7�M#>��?��j�?//�>�8�>���l���x��C�>�`�?O��?���>�0y?��u�s煿p�Z��	?�b?��&?�?�OMھe�>��?��P��8��+�Ծ�Gr?�F@6h@۔�?�謿�Oܿ������r&��V��=Kq=�_>���:J=��=���Ƽ4�+>s��>Z:�>u��>`a:>�>�>=���}-�-1��C���mq�5����G��	��ؔ-�Ă���辗�n�	,��K$����"o�;	�Ƚ�i'�_%�<D��=L>W?�W?�zs?'��>y���Z�>����.o�=]�5���=/�>��2?�M?�9-?�=�'��jha��{�2��獓���>:�@>�]�>���>�Τ>D,��0H>$v>0~>v��=y6м'�Ƽ�
=��?>`E�>W�>R9�>��6>�>p��r߰��Ee�+A����ݽ=��?Ś��fWK�╿���S��y�=7>,?�>�葿Nп���̂H?Y���s��+��H>�.?$X?]>���yT�P�>�L����g��{�=o����h���(�]�R>LM?Qzf>�vt>�|3�x8��5P��&��Q�{>26?>6���9�%�u�>H�$�ݾwHL>4�>uS�q��햿Y.���h��\}=<`:?L?����T�����u�u����R>�l\>[=<�=�QL>Ǧc�S�Ƚ�H���-=2I�=+�_>?��*>�k=:S�>$����	M��ئ>��C>��)>�@?�$?c!3�	[��Q��K@3�Uv>�.�>��>�=�=H�3k�=���>ŷ_>�%��������a @���O>'P���h���t�>��=����u��=q�=H�
�=�e�3=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�N�>R3�[3���@��wo�
k�<�Ȳ>��O?D���,����X��
?�H ?nT�������uɿ�u�#X�>��?��?*6h��嘿|IA���>J=�? �]?(j�>�9پ��6��j�>�,C?�O?kw�>=��
�Ç?�^�?�f�?��l>k��?7j?��>�S`��
�g����+�����Y�����=�˽���O>��H��'����s�L��o>��E<sԞ>��Ƚ'��z<>���;曔����y'�>-�>�-�>r�>RS?��>v[�>w��=#P�|��c�-G?���?V���f��ʛ�{��=�^��\�>[L?�s�ޗ۾�e�>ɛ�?6��?��>?tǔ>����ꑿi���%����u\<�Zg>�K?���>�z=N9�>�G��ý�r>91�>�����R�o���=&�d>j� ?9Y�>eky>:� ?�#?��j>R�>L8E�!ɑ��F����>E��>b?j~?��?ݧ���d3����W롿4�[��nM>�.y?�?
d�>�u���ל�Y�S���S��喽*�?��g?�� �?��?�q??��@?�g>x��&ؾ�̰�=��>��!?l����A��D&�t���w?R<?y��>����5ս�FԼy��H���<�?'�[?�=&?�z��a��1þn��<at&�MZ����;C>E���>�C>a��{��=�$>(_�=�]m�f86�/ug<��=>}�>2A�=n7�(]��QJ9?� R�b�(U!�7�!�`jP�S7�>`�T>5�˾՟v?5��,b��%����>Ι���|?Օ�?�Չ?�h���V�|&K?Q�?��3?��T�������߾l�־H�s#�~�E�PNq>@��>a0���Y�1���L8��GÃ�%��ۗ̽)�	?5F�>���>OX�>�h>��{>�̅��85��N﾿P�ei\��� �K7���@��0�W���|.ڽ`�M�����J�{qi>���z��> "?��>�!>�O�>��L=�
�>4:>�r>�إ>��A>�k>�Xm=�B�J�5�t-R?���V�'��n����B?�d?P/�>�\�������,�?�Ē?(v�?�u>h���*�o�?�}�>�R���
?X�B=�����/�<���ɵ���������t�>/�ӽ�g:��uM��kg�?�
?�?�L���C̾&�н�Ɲ���t=!D�?�5%?�='���Q��n��7T���S���*�r���8%��p������B������V(��&=<L)?�ʈ?y� ��쾻Ԯ���h��?��Bo>{��>�y�>☻>�	G>Ѵ��/��]���'��Ä�$�>�|?�ȓ>��d?N�6?E�V?�q,?N?�>g�>�žr�4?j�c�!��>V}�>�\?7�<?�)?s?�,�>x�=�����b�p?��1N?�J?-�*?)��>�(�>��T����p>�H8>Kþ��� "���;n>��f�	���R=�x?>�W?(q��8�������j>��7?k�>��>�.��,��`�<G��>�
?R<�>�	 �K|r��e�!R�>֠�?g���j=k�)>���=�\��RκXE�=�D����=����:�\�<7��=�͔=/�t����_��:�׃;��<���>�?��>�%�>��������L#��8�=I�O>|S>�^>�=ܾ��������i��~u>Ov�?��? �==B��=���=�-���¾k��v���L�<�J?B!?W�R?y��?%;?�z!? �>2~��ґ��&������e�?� ,?<��>����ʾ7��3��?�Z?;a����3=)��¾��ԽM�>�Z/�I6~�����D�[j��,��/��L��?>��?�=A��6�pj�a���XH����C?~�>xG�>��>e�)�]�g�$!�j$;>�|�>�R?#�>��O?B0{?*�[?�S>�h8���$Ù��I$��:!>�@?���?	�?�y?�Z�>��>��)�"ྎ,������B�dЂ��U=p�Y>	��>oQ�>�
�>H��=W�ǽܒ��%�>���=�+c>5x�>x��>.��>�+w>,/�<7�>?�5�>P� �Bb��yx���h�ե��0s?���?608?pP�=�#�֧S���
��{>A�?���?�@$?�ϡ�D�=��D��x���͢>���>ZdL>Ā�=]�=rx0>�G�>A��>�P��i�a������g?Y>?3�=ޙ��~�d���1��1о6��>�-	��	��?�뻁%��J׺n(澜�.>�"E��x�������������b?� �=c��<u�P=��
>q�
�
�>C��<��=^�>�E��SI���7н�3D=�P���V?�ݾ�;yz>Q�v=/˾�I}?AI?^�+?DhC?�z>}�>�=���>I���F?�mU>r�O�»��:�s��5ޔ��ؾ2,׾P�c�唠��>�2J��>*�2>=��=���<<&�=>i=2��=N�J�Z =��=�ݶ=Ɩ�=���=N.>�h>�C�?��m�=��$v���Z>I?H��>:�}>�ܾ݇?��=S��jž�=���)b?�� @hm�?��K?JB|��ؚ>��n�<�#���T>4����+~B>�-��(��>9�)=�l龛~����
�P��?�@s0?]b���ſ�5�=�>$4�=�,R���1��Ѣ<Ū�������K#?<�3��料��->�Y/>���C5��-��"�>���<�	@�19���c�=�4��}��<�F;ϕ>�V8>�F�=ю���=[��=�1�=`�>�Q��6b�|���-U�9��=�0h>��)>���>��?�_0?�Wd?(7�>�n��Ͼ�>��L�>��=�F�>؅=�lB>Ս�>2�7?��D?	�K?<��>ޯ�=��>��>ϛ,�}�m��m�>ɧ�,a�<ޖ�?�Ά?�Ҹ>� R<.�A����Jg>��-Ž�u?BS1?-k?�>ц��U����#������`=K߽�4�*8�t
���z��$��6�=P��>��>du�>��>۷�>Ci�>s<�>�Ձ>dG�=�|�ǄK�#>=R��=��L>b�F��ܡ���νV�E���.��/I��������#1]����lv���=>W��>F6t=(��>�9j=�A�����=HZ6�D_S��=r�����E�C�i�u�z��?_��� j>�Dl>V�H�,���V/?���=���=�N�?��?�������7����|��[hv�7�ӽBm�=��	>e���B4�X[�b�2�Ź��k��>�>=`�>IŐ>� 9�OAB�gB�;G�ؾ��1�,��>r���9����S�0q����R���O�q������F?�ʄ�,��=�x?zS?�܇?%��>̲��)��q{�>|qj���<�S"�W�R� ����?�M+?��> ���M5Q�%ơ�O����^�>�F��*88�����I4�S�>$˾.�>]��{<M��u+�*���H���+uT�w^��%�>?P_?z#�?XO�@�y�gW����Ƣ�=C,?�'w?�Tt>j#?y�?i�j<�d��Ѿe� >R��?���?��?7[>��=GT���>2T
?�y�?钑?��t?�@�n��>��9Ђ)>�R�����=��>�=�f�=�
?i_
?��
?�ܙ��	�|:�]��c��ɭ<��=�"�>y�>g�g>�=SV=���=��b>���>���>�Ap>�2�>�h�>Wp��S@����>>N�=�ʬ>�F*?#�(>+�=`ɽ�!>p8�<�ӛ�(w��p�U��F�63=ͱ�=�ұ=��4����>K�ƿ �?.�+>�>�$	?	�Ͼ�߽@^��>�D���w�>��>{.>��>� ^>��=SI>a�F>�����i�=J��<���о@r�����y�>�#;aƖ��L'�t�=={���
ھ[�&��J���d���X?�4�i�̻�?i=�"4��1(�����b ?Iy>�
V?�Q6�o^�>H�=���>#��>�A�5E���"������Ə�?���?#Gf>Y1�>��W?��?�]A��@3�GGY�cq��iA�&Fc���c�ō��<�����πܽi\?�w?o�??��]<h�w>��?x� �s���:��>�-��";�9J==Ǜ>ZA�� ai�Kj̾|���� ��<?>P�l?���?��?,�D��;�=s��=�$G?9�Y?.�l>9f?S�u?�J�bRT?^G����P?s6[> �.?�qm?��H?9ԩ=Mӽ-�O�(T�>������i���2Ľ�v����<��2>�6�<}
�E˂=_�a<[���>�`��<���Xj<l�u=��>���=N��>3U]?���>h_�>��7?W����8�q���;�.?9�Q=���ٍ��ܥ�N��d��=�Jj?��?��Y?�Z>Ѵ@�aI�	�>�C�>"&>�]> C�>��hL���=T
>��>T�=��Q��X}��O	����� &�<�>���>#^|>����Z�'>+����"z��~d>T�Q�tϺ��T���G�+�1�\�v�z:�>��K?��?p��=�J�P��=f��:)?�`<?�DM?1�?�Y�=��۾l�9���J������>4�<O������%���:���o:\�s> �������7�w>b�����
��*��`3�b���.=�Ჾ���=[|)����Q���lN>rk�=S�Ͼ�M���� p���G?�2*>޷�����!Ҿ˚:>O�m>��>�q�=����"�t������=�ø>�)�<������+�L�V��/<�>�dK?u�e?�px?�Ĉ�{�{�-CH�(!�`r���b=|�!?��?\�;?� >�Ȋ��b��/,�߅��U���>d0?�_㾫0�zvǾG:�>�:����=T�?��>�G?�W?7 
?X+�?�d<?�G�>j�w>��������+?2"�?/BY>U�>=~,�E����]�>DC?�l����>���>��?��.?zE?��?���=��ʾ��K�> ]�>�9X�����k�g=_�b?/t�>`y?S��?��h��]H�(���=�$�Ƭ>�Di>��L?O�>���>1��>	,�>�*S��?>S��>�#J?���?�x?)>L?�S>|��>�({=�|�>�>�A
?�-8?�l?7�A?^��>�w<�����']���;'�=�b��b]��3E;C����e���;>.�=?/�;Xi]�r���&�^��'�<h߃�(��=83�>�x>�0��׿5>�MľP���:LG>�Ԏ����l㈾W�5�}w�=��>�� ?�ɐ>l*��C�=���>d��>?}��A'?˱?gp?�w<��^��=ݾ�uQ�别>8�@?�$�=چl��f��?st����=�"m?�\?�S�������_?Ž^?���v=�۾�/W�z�Ͼ�HR?~�?��L����>�w?��t?8L�>�-���{l�������d�V�Y�D'=t��>���ٚc����>"�8?��>�pb>4��=ٚξAbn�A=���K?u�?�?���?�5>�m��Jڿ�G�Ɇ��	0?�= ?U����^&?,E뼁wȾ�X������Y�۾�(�����[������X�1
L�:^}<� .>�?�|?J��?c�r?,�ؾ��^��X����;x�����=��[G��F�c/7�`�[�Ӿ��w\�|&m�O�̽�U}�d-8�d��?9�?EƓ�3��>���3Q�r���pSY>w�ľE������=E<=��} >��=(�W�������G?*6�>��>��4?�J��?7��O.��Y5��j�<j�=L&�>ݪ>�:�>8�=�)O��X��оGl���fX��Fv>zc?�nK?�n?����0�g��9s!�"�.�./���C>�>~��>;OW����Q&&�K>�es����s��>�	�N�~=b�2?k��>z��>�=�?F�?�o	�������w��~1���t<U�>05i?ԁ�>aۆ>s�ϽU� ����>��l?0�>Ւ�>�J���7!���{�pj˽Q	�>b�>5�>7 p>�	,�"\�UW�����h�8�P�=ڀh?Gd��oT`��ۅ>L�Q?C}:�B<��>yJu�FU!�h�򾣴(���>�\?ט�=��;>�<ž;��i{�����$?��?I�����t�=�ZN?�P%?W��>�k�?m��>� ��\�����>�R_?I+D?
�7?K�>�R=I��Lս����^�?��=S�>�>W#�=��/��۔�a
��?��<�Ic>��=��z��>����a6>���=��=��ڿՕJ�*�ؾf`�*���	���5���1����k׷������u�7�*:�1GU�fc�eG��hn����?־�?wB���]���X������{�����>��k��뀽\-�����Q5��T�ݾ1����w"�E�O�O:i���f���=?���ϯѿʶ�����b ?��<?ȸ�?�jо�{)����Q�S>�(��_=�ڴ�ί���2俻u��zr,?آ�>����y~�?񜵽�~�,��>ܯp�������b*?��L?)j�>��ɽ�̿�˿������?�@8aA?51(�0���\=v��>̠	?�jA>k;1�$���7�����>b�?@ʊ?��K=jW�O��8e?ט<�F��Jֻ��=��=E�=�����I>�ړ>b��B���޽�3>#8�>�,�v���\��`�<o�\>��ν��3Մ?){\��f���/��T��U>��T? +�>g:�=��,?Z7H�`}Ͽ�\��*a?�0�?���?#�(?7ۿ��ؚ>��ܾ��M?\D6?���>�d&��t�Ʌ�=]6����y���&V����=^��>h�>��,������O��I��?��=+h㿡�ǿ3�F��������s�����K	M<�7�����8��ˉ��䉾p�q>�>�^�>�Y>�9�>�<?��??��!?-�>]�)>�f�FN�ͷѾ,k��r�"��^�����Ll�ќڽ�P���Ѿ>�򾷣
����'۠�#_德q>�r=�ş���R��F)�\_m���#?}�?9l��S9c��P�<�1Y��_F�
����>���˾�fJ������ԕ?N>?߾����8�Ɋ��f��m���1_?S�>Ɣ����5=�>���Ϸ����=�=h]˾:W9�W�1�U0?��?�����)����3>^lͽ B�=l�'?u��>��< V�>��%?��#��۽�u^>�V>BH�>�)�>��>~���+�ν�%?7oX?~J �6$�����>ȾΔ��΃�=*	>X8��,K�ܭ6>�J;�싾0��:�ȏ�L�<'W? ��>b�)�� ��[��!��H�==O�x?ܐ?�2�>�zk?��B?�Ĥ<Fb����S���pqw=��W?
'i?C�>r����оhn����5?��e?�N>]ah����p�.��U��!?D�n?!Z?՝�du}�L��y��n6?��v?s^�ts�����M�V�_=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�"Þ?��@���?��;<�����=�;?f\�>	�O��>ƾ�z�������q=�"�>���|ev����
R,�f�8?ܠ�?���>������X>��`�#(�?t~?�|�C �tk澄T�p:پ[&
<y�>*�c>�G7>U1���C��<ھ ��~��Gc�N@>�j@��T��b�>'�?�GRֿðܿ΍��﻾�S����?i��>@S�>;��������K�nA�u)��g�¾�X�>g>�s�tY��Mt�*M6���H�
��>�2��M�>�V��S��CC��_Q[<�B�>%;�>�j�>l����[���,�?~�
cͿ�#��/��t�X?l�?��?��"?��<��|�2T���`��)H?��s?M�Y?XS�bNk�v����j?�O��aQ`�φ4�vSE��U>�%3?�F�>��-�P|=,>��>�Z>�/��ĿLܶ��������?���?�y����>�?�x+?�a��2�� f��H�*�JJ&��9A?�1>�����!�^.=��ג�I�
?��0?t���%��N_?�_a�x�p���-��PýB��>�:1�l�[���� �c�e�,���y����?�L�?"�?N�:�"�L5%?w�>;3���Ǿ�,�<���>馶>"�L>!�_�wRt>����;�Ko
>��?T�?fu? ���Dߦ��>�F}?�o�>�σ?�=	��>�Z���Δ�ٰ=�^>�>
>2��Iq ?HZA?� ?�y>�fl�;`*��PB���]��1�(�@���o>��T?ȩ7?�b�>>6;KI���o�ϒ��ꋽ�ug=�g=�[��c���c�>�w�>�N%>f�	(���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Pa~����7�^��=��7?�0��z>���>��=�nv�߻��X�s����>�B�?�{�?��>!�l?��o�L�B�`�1=5M�>ʜk?�s?�Ro���g�B>��?������L��f?
�
@~u@_�^?(B�׿F|���dϾX���;<�"4��w�=�ѿ����J�1�&����#�>���>ư�>*��>;4i>z�g>��>�����#�t���κ��F���J�F�.���Ͼ�J���� $�z��� �����=��=4E�=����g,��������="BU?o�Q?��n?s  ?�<i��#>�>����=� ���=vA�>��1?RL?'�*?,��=���Oe����;妾���#e�>�J>(��>��>{�>̄��H>��?>�r�>�>z�!=}�n�Q�=c�N>��>���>g%�>A��>���>@������'�G��m�G�����?�M]=V��˴��Rz��c��\E��r?}�<�"��N#ֿ���D?"|y��p9��WT���3?���?u�>N*��*ˀ��>=>i;��h�0�]>n�=>㵾Ҍv�j�o>��?��e>��t>�E3��e8��#P��(����{>��5?l����8���u��H��_ݾ5�L>�K�>	�+�'�����-}~�M�h��z=�X:?�1?짯�㱰�\Ev���(�Q>��[>�=�Q�=�M>�Ga�X"Ž�H�?�*=j�=��\>�`?L�X>�k�>�[?Q�@������>�Ѓ=�=�O?�f<?�>IBg<ޜ��|���L���>���>�>NB��U)>��>�W�>�JK=��|�k���p�q>�"���ľ2�=����=��9v��{��<H��f�T�Ӽl<�~?���'䈿���d���lD?Q+?X �=�F<��"�E ���H��F�?q�@m�?��	�ߢV�?�?�@�?��Q��=}�>׫>�ξ�L��?��Ž3Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�?l�z6>�^%?�ӾPh�>dx��Z�������u�}�#=Y��>�8H?�V����O�i>��v
?�?�^�੤���ȿ3|v����>T�?���?_�m��A���@����>8��?�gY?toi>�g۾/`Z����>λ@?�R?�>�9�^�'���?�޶?ӯ�?��J>W�?�s?|�>�}��a0�넳������Tz=��<�:�>*D>:���cE�����݈���j�{��>wV>�!=J�>�ս3ֺ�Qܠ=d搽� ��`����9�>ԏ|>��O>���>� ?��>+e�>�a=[Y��e����T���J?�E�?�B�?Dm�I�j<.۱=��M�'�?ٙ2?>�"���ƾ�_�>b�Z???r�W?���>i�Rԛ��9��/6���0<��L>_��>w�>�'G�zH>u�׾1jC�̣�>�_�>��μ²��^��.3f<%Y�>T�?���>e��=� ?�#?8Xl>l�>��D�*����E�a�>���>��?��~?#�?!���43�Ւ�Wס�0)[���N>m�x?�)?��>�m���f����K��H�W1�����?�g?� ?(��?V??��A?v�f>�
�3�ؾ.����> Q?�f��W�8���%�����?ڊ?���>��>��g�p��<����G���?�gW?j�%?���|h�m(��{��< c�>y�<R	=��=��G>S�>�>���u�=�G>{S�=On���U��J���>�C�>㞪=�\'�aKڽw5,?k1H�5ۃ�G�=��r��zD�Z�>�'L>^����^?i�=���{�}��w����T�R �?Ȟ�?Mj�?X��Ęh�^=?�?
�?�%�>S?���u޾n�ྱ&w�nx�4p���>L��>�l�j	�X���:����D��ƽ�ߩ>B�>+��>���>Q'/=:�>>�\��"K1���!� �%�k�@z(�pP\����&���(�.f�=I��;f����C3�͏�>?������>t ?�R�>>>D>y�>a>���>�Ω>]�d>��p>�2+>UD>�3�=�G9����#$M?����I�%������Ѿe�:?��g?�B�>%p&��Ă�ɳ �j�?�3�?�J�?K�>>�e��
*�I�>���>/��/�?W�]=>�ݼ@P�=�q��w�#�����⪛��q�>.����2���L���X���?�?���;g�Ҿ.�������o=eL�?�(?�)��Q���o�)�W�PS��x��Eh��i����$�Ԙp��쏿�^���#����(��>*=�*?2�?E��V��^"���$k��?�"lf>��>$�>W�>�nI>��	��1��^��I'�[���6L�>~X{?1��>]1E?Ϲ<?�M?PE?{ �>��>삢���>�EY=�`�>���>	�/?�a%?�(?��?�y+?�g>�2½@O�i�پ?d� ?;�?�B�>��>�}��)3�����X;�O��� b�EB=d��:�R�~G�⤖=��u>A_?���_8�-��Tk>F�7?'��>X��>�ݏ������<L��>�
?qˎ>����cr�%��R�>���?&8���=�*>$�=�툼c� ���=�"ü�Đ=�灼�k<�Je<�G�=���=����D����!;N�;�J�<�K�> �?}��>_��>*����� �rw����=}�V>>�P>��>m�پ|x��]R��y�g���y>�o�?�Y�?k�h=jV�=)�=a���7����Nܼ���<X�?�#?�DT?ll�?��=?v#?�>n�����#������y?��E?�W�>s,�����ɿ�{6�G�4?d�1?U����#1ھW�%���D�r�l>�c�Z����/ӿz���p���@���?��?���f7��&���C��dU<���9?SW�>d(D>ly+?��!�G�����پ���>G�>!�S?+{�>�/]?rq�?�e?��>H�6�!��ƍ���C�=���>�-V?@]�?��?�_�?���<cO��m�'�B�<��i��y<����ES�=z��>}�>��?��>37>r?|�2�@������̀��Т=z·>��>�E ?� 
?�&=��G?���>v���sz�c̤�{J���{5�}�u?o��?ɢ+?�-=�r��E�����H�>�H�?޺�?��)?ʒS�j�=A]ռp��E�q��L�>��>�~�>��='3A=��>�|�>4�>�5�^��58��LQ��6?aF?d��=-���*���׾��o��� �gξ�ɵ���n���Eѱ�M郾M�E�|�ɾ�;=�M;����	O��X�6�_����>���=��=)��=�"�|�z=��|=L0b=+��7֓�
H��-�?=�~`<��L��u�E��;xI'�7�<�ɽ�*��>�z?��>?�� ?I�@?��>{	J>��t˕>$m�97?1�E>�d��U����	��1�����о�]��>���#>�ü�-4>76>���=�
���=�˨=��=t^���=���=��=��==P�=��>���=�/w?Й������B6Q�>*��:?�5�>�s�=Owƾb@?��>>2��2���Jb��,?���?@R�?��?�ci�De�>(�������\�=z���~62>~��=��2���>�J>���II��낳��1�?�@�??iዿġϿd/>ls>X��=��N��m-���\�
�o��Pi���?�:�_QҾj�P>u-�<
��,����{�=�ZB>v�=�_��hFS�e��=s�����=��=��>1;F>�Ȥ=Q������=@�='i>�eZ>��;p�����<>L�=�KJ>6�>?��>�?5�7?f�f?��>�4�$����E����>[Ql>|�>,�>�s�>͟>d�?�06?vzG?譧>������>�T�>��-��j���ʾ{&P���?>&4�?��x?��>p<n�t���C��R�0�[=��?�/?,!?�M�>����p޿��B��'�@Jӽ36���pt�f}��e��I57��<�`P<�b7�TT�>�s?�,�>:�>fA�>(��>�F�>b�л�I�����=�����=|�<��u>*U�=U(:=,�>xM��Ccн�U8��	��,�F�~>�T�==83%>�s�=�E�>�B>r��>XT�=�����->ӗ�M��Ҹ=�ը���B��$d��~��[.�]`4�64E>��Z>@���Ƒ�/�?)�X>|�;>�-�?='u?)�>�t�}ӾQ���Kc�(�S�
}�=��>F�;��];���_���M�77Ҿ�%�>4t�>�C>)�>0k�M,��^T>�&�����+��>�X>�Pu?�{�����K�����-��E"|�M۽�3?�����$>N�x?&?��?�^�>������ξRRH=#�'���@���'=}�v��o'?��M?��G?h��F̾�����>z;I���O�p���d�0�	�ͷ�;��>�����о�#3�h������:�B�[Dr�:��>3�O?C�?�2b��V���UO�R���#��Uq?h{g?�>�K?�??k��8y��q��u�=��n?���?�;�?.>u�J>W�<�o
?��?��?I�?�?H?.����x>��<��=��`��д� �h�]�=hl#>ܩ?��?��?�i���ѾX�$��.�Ό ���=�&5>!p�>���>+_�>01�=�*�<�Z�;J�)>e�>bZ->������=9�>�fd��޾�%?�=��i>�2?_߸>�#�mM9�J!>�ʳ=�B��������<��K=�������ʒ��4�>44Կ䓣?!�g>ɔ����>�X׾/���[�>�&�>��ݽK #?��,>�4�>��>��=�Z>F#�>De=�WҾe�>�n��w"��A���Q��9Ӿ�y>0�i8"���	�+��mmE��ϳ�l��Cj���lX=��o�<�2�?	%���l���*�Ce��DL?O��>�~6?S���#��L>UC�>�>�r������3����c;�?`2�?���=_y>��?�30?��s��ϾZ�E�Fv���2���	��4����q݀��?�����bYC?�&|?;tb?��=S!;><�L?�r!�s,۾+�D>(�1��Eپm��4T>4]T�����E���_\��G�K�M_p>+�F?��A?CW�>��q�n��=��s>"�@?��?VMI?&�S?<�W?��;��?�>�'?�?{4?�+?�W	?�$=��V>)�=��D=�nK��4qu����=��)���=L���3m��r�c=o�X>>({=�(��؇S�����㏽�V=��{<O�N>��>.�R?���>Ʋ�>l =?��ս�l%��S��Ms?D�<s
���N������[����>A�e?�D�?��T?ă> �#��+T >w�S>̫;>�x>��>1�޽�yE�L^�=��>�za>���=m�A�L�C��m�d����{�Q>���>��z>�ҋ�J%>u%���z���b>�!R�����zR�`LH��U1�K�u����>?L?��?�B�=%;��s��3Ye��(?J�;?��L?؋?��=3�۾�9��.J�De�%�>���< �����H㡿�?;�����r>���?��TNa>h���~޾bXm�h&J�����YQ=r��<�Y=E`�]�վN��f��=�|>X����S ����^���f�J?.xo=ä�/rS�xg��0�>�ޖ>(b�>�:2�Q�w��@����D�=�'�>��9>�z��q;�`_G���h^�>��C?h�i?�9�?
ګ�$6f��L�8S�����T�,?j�>M8?փ>W>~h�� )�h����,M�ղ�>��?ٴ��Ug=�P�8������5�k��� �>e�>�T%?npp?v?l�f?j?�>X_>��n�8\ɾ3&-?s݅?�~->�]9�o�D�ӽ �),��|�>t�)?������h>b�
?eL9?c�/?*w<?�#?�6r>�`��r*�@��>�8�>H�y����9%�>��a?�?
Yu?P�{?ru(=�'B�?ܾ���>��=߼T>�s0?z� ?���>��>��?Y���>	�>�/}?x�?��b?�b���>�>7��>�+=m{A>f�>��.?YF?��o?|�P?��>���<2٨��U���c���ݼ��.��V�*&�=��:��(=>���<��<����0���=�S�7�A<X��=�t���d�>��k>,��ÌC>_����?�(�>>��Ӛ�n��;.+�é�=�G�>�*?gē>	��$�=K�>���>�w�s-%?^ ?ҝ?���;8R^��Ӿ�'E��"�>�@?�K�=�k�����v���N=�o?�_?�D����I�b?��]?h��=���þJ�b����\�O?M�
?�G���>��~?c�q?N��>��e�:n� ���Cb���j�/Ѷ=cr�>RX�P�d��?�>a�7?�N�>'�b>=%�=fu۾�w��q��i?}�?�?���?�**>��n�Q4�o9�t���"\?Ѕ�>\Y��O�?oF�;�̾�,x��[��3�����������(���)���}�ͽ���=��?VSt?��m?�]?Ο��Le�"U_������pZ��T��Y�RD�w@���@���k��
�����ƣ�-'�<GmG�n�6� ��?� )?O>�.��>�'t���꾮6��d>������
? >1$�� 
�=L��<@����-�����?E��>RȽ>��5?*`�A�"9�<�K����y��=U�>��>7�>?��;1�A�㽑�վ=���jE�mx>n�b?A�K?�Jn?�����0�TN��r�!��y<�2N����C>h\>��>2&R���Kl&��~>�^^s����KD����
���}=�b3?,w�>%۟>L�?&�?"���宾R?v��}0�PNt<���>{�g?���>};�>>�Ƚ&��A��>E�l?٨�>L�>ܓ��Z!���{��ʽ!�>�ޭ>��>$�o>��,�"\�Qh��c����9��u�=x�h?₄�7�`���>UR?���:��G<Xt�>Ow�0�!�����'��>�}?���=��;>Q|ž�"�}�{�#9��?-?��!?ʛ^�x�����>E�I?��?�Y�>.�{?"��=>�¾�ԓ�!�?Gi?��A?rLZ?���>���;�������%�Ā���R>�Ҍ><��<��=��,���S��
��?�=��=<���k����=3U<)�ú�
�=bE>��ڿ%�J��پ��Q�f�������C���'����c������9{������Z�vV���Y��6��[o�\��?z��?�ґ����aט�������f�>��d��u���������x��ku۾������p�Q�>�i���g�B�'?�����ǿ����:ܾ�  ?�A ?�y?����"�Β8��� >.1�<9���뾭�����ο�����^?���>��,�����>'��>��X>kKq>���{鞾�!�<�?W�-?���>�r��ɿR������<���?��@�[D?�#�Vž�=��>b�	?H;>��N�R* �Fϼ��l�>��?���?���=��N�c*s���U?\��>�.aL��sy=�׮=�7�=f�4��>�Ы>c��{L�~�ڽ��0>h~>�ՠ�BFG�T�j����=goy>��i�IjZ�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=o6�􉤻z���&V�|��=[��>b�>,������O��I��V��=��￡չ�z�J��l<��P���g�<���0�>�ч<�==yž��瑘��9�%��>�ʒ>�g>��S>pΛ>��"?�=E?���>R
a>(�{=����A����(�z��53 <#����㭽[�A�R_پ�:��4-�W����f8�%���@`�=WX�h��2I��AT��)�����?'9!?�����������s�;�#��~��ۼ֧�'4;��F��(:�?��X?�����.n����Gu��Mܽ�?�Lҽv��y���z�4>�Z���<U�#��>o�u0!�ZT��cRt���0?T�?"��BS��F@3>0Y �z0=�Z+?�p�>���<u��>�`&?'�(�����T[>2.>
��>j��>��>����w�ܽ�?d\S?}��ۃ��Î>�K���{���n=�_>��6��dܼ85Z>���<����������<V�V?ҳ�>(�	.��9����"��v�=F�w?X�?�1�>��i?q\D?�&�<�b��QR�k���O�=!1Y?/j? �>�Ɔ�u;<���X�5?�c?�Q>�ab�:��c,��B��q?��n?�
?K4��{�{�Vے����=_5?��v?s^�ws�����;�V�c=�>�[�>���>��9��k�>�>?�#��G�� ���xY4�"Þ?��@���?4�;<��K��=�;?l\�>��O��>ƾ�z�������q=�"�>���|ev����R,�e�8?ܠ�?���>������A]>�v��ds�?�?��ʾ�{��*G�(�j���ܾ!�=���<	�.���=���=L�9�Ծ9���˦�������n>��@eᱼ%�>�u�>ӿ�Ͽ�9��J�_ح���3?c��>M���u�(�_��Ic�q+B�__�, ���o�>�T> ��������{�K2;��ូ���>b�e��>T�y ���B����7<Կ�>���>2��>*��=轾^��?�"���7ο�����	�X?�u�?<o�?]?��-<V�v�l	|���1&G?qs?� Z?��&��5]�Y�6��j?�[��oU`�8�4�DE��U>�$3?>D�>Ɣ-�+�|=� >���>Vh>�&/� �ĿFٶ��������?E��?�l�&��>���?r+?cg��6��nZ����*���7�z<A?12>y�����!��.=��Β��
?�|0?�~�$,�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>bH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?pP�>-�?7��=x$�>�k�=�԰�o�7�s!>���=pR@�W�?�zM?c�>x�=Z�8��/��5F�	
R����C�}��>��a?ML?��a>v���e�6�j!��EнW1����?�1�&�'�ݽ �4>�>>Va>��E��dӾ$�?�j���ؿ\h��hV'�K14?.ă>��?���T�t����B_?4z�>s=��+���%��'=�j��?�E�?-�? �׾�&̼<	>��>8H�>�Խ����ێ��p�7>��B?� B��w�o���>b��?��@�Ѯ?��h��	?���P��Va~����7�g��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?uQo���i�B>��?"������L��f?�
@u@a�^?*A�ҿ�Y��KM��rԾY����:=�qQ>�Փ=uF�<,[�=���=i��<�	>.��>J�>�N�>zn�>�E�=K�]>Ԕ��<b&�2c���Š��!Y��վ V!�D�s������B޾92���B�X=�7���{>���4	����?�8^>rN?�eU?��r?51�>Z��U> �1~�<t�1� �=�H�>N�4?�eK?-�%?A�=��;0d�h�z��S��Y͋���>�Np>Ň�>L>�>ё�>W�U<��h>L3A>�΄>	H�=�}!�J��e��<�Yp>���>���>���>��Y>�l>5�����r�K��ܬ�۟=��f�?t�z�>�Y�q���p�n��Y�C>��� ?��C<�C��m���ֹ�M-A?�m���"�	qݽ<R���K?
j�?��=����sM��ɽ�>U�����ƾ�P�><�H�M�����U>���>"�e>_;w>0i2�SZ7��Q�.R��j�|>5?+崾
�:�!4u��DI�4&ܾ@4L>�	�>^�"Q��,����~�.�n��Wq=�l9?�?�\������3�s�5F����R>��^>OA'="��=3}S>x�w�1�½;3F��\=Ͷ�=_�e>V�>)k�=�5%>?��>ǽ��������>{kJ>\�>`�H?.?�W������r���ֽ�
 >"3�>$��>j�4>�!��E>� �>�L&>�ؑ�±Z�����F\���{>�g��r���'�=b b>�_D�pFR>�1>2K*�t��<I��~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾQh�>rx��Z�������u�[�#=P��>�8H?�V����O�\>��v
?�?�^�੤���ȿ0|v����>Q�?���?f�m��A���@����>9��?�gY?loi>�g۾>`Z����>̻@?�R?�>�9���'���?�޶?ԯ�?_�I>t�?X�s?�5�>�Uz��@/�� ���㌿�x=~i;�g�>�r>���ʼE��v��%8����j�+"���_>m�$=ʏ�>���ռ�8�=_��3����An����>��q>R.J>��> ?>��>i�>;=�4���-���薾t�K?ӳ�?����/n�҂�<sʜ=ء^��%?I4?[i\���Ͼ�Ϩ>޺\?�?�[?�k�>����<���忿�~��{��<ƾK>1�>PJ�>C-��CK>O�Ծ�3D�xs�>�ї>�%��|Cھ�*���9��/B�>Hd!?���>�׮=� ?:w#?��j>7�>�TE������E�~��>��>(J?��~?b�?6乾�[3������䡿��[�A�N>+�x?]E? ˕>�����q��G	F��
K��󑽇��?-�g?佷�?gC�?X�??ܥA?	�f>�	��׾�0���ހ>7�!?���i�A�2B&�����?w^?e��>ْ�cֽ�׼L���X��~?9"\?�K&?2���"a���¾^��<:�"�g_c�v��;ψB��>��>����.|�=s>��=5im�<m6��g<Ҭ�=q��>���=7�Y��-=,?��G�ۃ�)�=��r�xD�+�>�IL>����^?5l=���{�����x��.U�� �?��?Zk�?�	���h��$=?��?G	?�"�>�J��I}޾���(Pw��}x�ew���>C��>ڙl�%�O���Й���F����ŽF����p�>���>�b�>Xf�>�Z!>ɝ�>��۽�� ܾ�{��wAv��?��O9���?�d.��O�� �Z���=�ri�������l>��<���>y?V��>��>�\�>��=݀o>�]�>@��>e7+>�Dg>I��=�܇>s&*>&��=0LR?]���#�'����#����/B?Vhd?`�>Di�d��������?凒?�p�?h;v>�yh��++�bc?�4�>[���e
?�E:=���~�<<���� ��O�����>�3׽K:��M�đf�#b
?�7?�����{̾�ֽK���L�n=sM�?x�(?9�)�r�Q���o�Q�W�S���1,h� p��$�$�q�p�%폿�^���#����(�Js*=?�*?��?(��������!k��?�sdf>J�>�$�>�>�sI>��	��1�� ^�(M'�񹃾�V�>,[{?�M�>^ZI?٣9?�M?ͽJ?�M�>z#�>8޺��7�>�ǳ��r�>���>ˈ2?Y6?�,?D�*?
�(?�w_>zHI�����0˾(��>��?<�?���>���>�ݤ��͛��U�=9�s=�]k��CX��[���3�=��٭;zL6>��G>#>,?m�c��k;�l�پu?�- ?M-?9 ?���t�F���&>��K?��?wབྷY��dȀ��پ�9$?��?�E�o�!�N>8�>��w=�Y!���k�����k�{>��9<;@�!K�=��>6kY>3%�<�,�<2�6�%>}�>��?<��>�|�>����0� �f�B�=��X>�T>(>�Iپ<d��'����g�A�x>���?�o�?��j=��=��=�i��e����벽��#�<ٟ?�F#?*4T?o�?%>?��#?�.>�3��J���a���<����?��$?>H�>D��|�	��Ǿ�1�C�Ք?h��>G�P�����)0�͵&������=�pc�'�C(��,)1�����R\۽��?���?�uT��.������d��P:�\�5?��>�|�=�~ ?CӢ�y� �����b�=���=-�b?)&�>�9?���?:d^?��>El�qi��Fܫ��7�� z�;3V?���?H��?J��?�=�>����s����@�d��
Ѽ=��q��p�gz_= 9>W�>Z��>� ?��
>%^����2������=��4>sn=>D��>B:�>���>�(>I�G?���>w���'������5���9��u?�M�?V�+?��=��w�E����L��>�J�?��?<�*?\�Q�0��=�8ڼw���PXp�q�>@��>D̘>(�=j)F=��>�N�> ��>�[�f���8�d�L�̔?F�E?:̿=zſ�q��w��b��D��<K|����f�B`���T���=�����c��.�^�x奾��������ʞ�8"y�LB ?�F�=l�>��=I�=�C�=��;�1!=��<�P	=%jr����;�G%�8.�;,Ө�7�;�:I<h�=�Q���y˾(~}?�)I?<�+?3�C?�ny>�z>1)3�!��>M��e-?s�U>HP�������;��������t�ؾ�p׾e�c�V�Gi>7J���>Z�3>�&�=J��<�/�=?r=��=�^�`z=��=�j�=�~�=J��=��>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>έ7>�>�hR��E1�37\���a�m�Y�ȱ!?�W;��X̾�z�>`��=�j߾^Ǿ�y'=��4>W6b=���l�[��3�=�C~���<=�n=w҉>��D>W.�=I����u�=,sK= #�=�O>dx���09��*�vV1=k�=v�c>}�&>~W�>��?Q B?	p?�ӫ>����\�ǾL.龞�{>�[=�F�>f)�=�>���>��%?�G??�P?R0�>�T}=%_�>��>�-���p��~��r�{�=d�?Q��?��x>��۽�%j����Dw4�Q%��n1?Ǌ,?���>,��>�3���ۿ�>a��9�G��9�=F�E����<�$R��=,�ne�=�T'���b�X��>M��>���> {�>�4�>���>Rk�>a�>ӂ=!��,"�=�����a��b=�e�<H,��������<�=��O���W >n� >�>+�X>�m&>t��=���>#@>��>Ŏ�=����M/>����V�L�ҿ=�F��$,B�V.d�pF~��/��]6�.�B>_'X>D���R3����?��Y>�n?>��?�Au?��>��d�վN��u3e��8S���=̨>� =�Nx;�P`�q�M�gnҾ��>'W�>[��>dWk>�k-���B���=���/�#��>�o�q�T���
m����:ݝ�L�j�ls�W;=?�눿2��=T�x?.�I?�4�?���>gr���Rо�82>�vr���@=)��/'R�#}���?B�$? !?�;�:��B̾�����>C:I���O�ٺ����0����з��r�>o媾x�о�!3�e��������B�<r��к>ӧO?��?��b��J��_KO��������Uf?�{g?J��>�D?�J?�:������i��&J�=��n?B��?�:�?m0>�oR>�:�:�8�>��?���?C�?�p?L�/����>�%>P�>�(꼬I�=E��=���=�5�=�R
??G�?��U���ھ�_پ̢Ծ$_����8@�=�cy>���>ŕ�>cc����=���=~WZ>R!�>���>��x>��>O/0>���E��U�#?�h�=">I�?��>DG>��[��B�����=Mež׏���1�㰤���|����<�kV��#��jG�>�EȿV�?�_>_`ž'u6?�6�z=��=��h>+�=�ߣ>�{��L�A>/E�>Q#>���=ӆ�>��>�Ӿ��>����W!�LC�AqR���ѾRjz>�Ɯ���&��y����z(I��[��R~�lj����4J=����<�:�?b ��rk�չ)��?����?�R�>P+6?����&��"m>y��>N6�>����������Q��?��?�=c>��>O�W?��?��1��3��tZ���u��'A�!e���`�፿����^�
�O�����_?*�x?�yA?�f�<z8z>뢀?��%��ҏ��'�>�/�V&;��?<=�*�>�(��%�`���Ӿ�þF9�9FF>��o?m%�?�X?bQV�s�=�>d8H?PX?u�j?��1?��?
7M�^�$?�z�=�P ?�^?%�?U�0?��>{�.>Hz>)Dh=��=:᣽f�'��L��Ҍ���*�����9�T�ṳ�*��m��=�,�<*���R���=[*2� �F�=��>�=1��>��d?��>�,�>�#U?����_�M��L�	?3\�>�B@�����丘��n
�q��>��U?�ϻ?Z�v?�>�^9��&S��!�=}��>L�g>�o�=i��>��=f�� ��=��=T8�>�U>�'���=%���@��G�����>*��>]|>!9���1(>n���x|�
e>58R��˹�:eS�z�G���1�u����>jwK?{_?F��=���o0��h)f��)?P<?�JM?��?c�=�ܾ��9���J������>h��<ZB�ۋ���ء�dz:���H;�qq>�����Ƞ���a>]u��9޾�{n� +J��O�
IL=̗�]�V=�"�i�վ��}����=�	>����� �^���֪��J?�^n=􉥾n�U����D�>�o�>̟�>p�8�%w�v@��}�����=���>�};>H������G��4��ɘ>И+?o�n?ص�?U-���h{�+�]�g���H辀<1=(:?9;�>y�&?�=h>���<􈮾VY��ke��~E��$�>k� ?׵�m�L����5��W ��g�=Dx�>Z~�=Ӝ�>'�@?�z?�0k?$?Bz�>�5S>��ٷ���/&?Ms�?���=�m���,E��!��@6�ŧ�>c�&?�U;����>>^?�(?�/?B[L?k?�Y>��f�3�Ab�>}��>�aN�ah��i 0>�1R?���>qr_?�ل?���=�7��@ʾ�����=� >��,?G�)?��?�`�>�S ?_a���I;=�L?�|'?/U|?�-q?tP׼���>� �>�>5��=�p>7��>n��>k�i?I�{?�Nc?%b?������ �+<�e����ϼ����ח�=����M+K�Pק>I��="ol�3�	��l���>��Xʎ=��=T�>�du>������6>ʦ��S��qJ>�t���xN��24����=#̀>�R�>R�>Y���(�=�w�>�\�>�J�֠*?�a?��?(��90b�I�Ӿl4A���>�M=?P�=Q�m������w��\=�j?��[?�)\����i�b?��]?�g�=���þŸb������O?�
?��G�u�>�~?:�q?��>��e�#:n�8��Cb���j��ж=�q�>�W� �d��>�>�7?WO�>�b>a&�=�t۾��w�Vp��s? �?��?���?R+*>��n��3��7پ�x���_?X)�>88׾�'?ʏ�=�Pھ�L����R��˟�>�I�0���t���I��҄�Hj���^��6h>R�"?�[P?&�f?6�Q?cޝ��>��m�2�\�`�~�^��aY��LF�3�@��p8�=]]���1�:�ʾQ}d���½Þi���G�<��?��&?!@?�`m�>����':򾴧޾��M>D�����޽�S�="����B='o<�k���0�����e?��>�B�>��9?Q�L��:;� �;�%2��?��#>��>�։>���>�^<�A��� �8*ž-���|���-w>|c?H�K?�n?	���Y1�����Ѓ!�b�8���}B>x�>^ʊ>��S�!F���%�J>���r�S�������	�Ŵw=��2?Zm�>"G�>���?��?I��H\����v��1�~;"<z��>�'i?6$�>��>�LȽ�j�qr�>r5k?x>�>���>�^C�m "�\Ke�*����[�>�+�>U�	?�C>��6�=�O�F����֒�B� ��>�el?�oY�6���a@�=��Z?��?����|��>J&z�i�������䫽�+>8?��>f�G>�pܾ���>}k����i(?��=?h������]>>�??�X?N�>��w?�4>�׾7<��=)?UO?� U?� e?�h?\>㗣��	%�էw��h��9�#>C�`>�GӼ���=$������1ؽj�=����; ��S�/�:�S�<oO>�%>9t>!�ؿ�uJ�a[۾b��Rؾ�8�k̙��̈́��+W�'�<�Ⱦ���f����K�����ڎs��D����Ne��S[�?��?gń�����'X���4������)�>��R�4�z��i�����r��<۾<P��yh�1�=���l��6m���)?W_��Dʿ�3��`*�>�	?.�?뺑?7�þQ�c�4���u2>��-��A>�晾R���r��֊�y�?��>z[꾁Í��B�>�%f=���=)�>�.K��:��Vh�ڜ?��/?�~?ް�;�.˿Ɋ��ԟ�=	�?�/@�;A?�6(��3�Ti=qI�>��	?��@>�3�O��qD��JF�>�4�?�Ԋ?$�I=K3X����Ƈe?��8<��E�=.л#N�=���=4J=�I���K>�̓>����L@���ٽ��1>�C�>�:�'��G^��<1Z>��۽�J��4Մ?&{\��f���/��T��U>��T?�*�>Y:�=��,?V7H�`}Ͽ�\��*a?�0�?���?#�(?6ۿ��ؚ>��ܾ��M?]D6?���>�d&��t�ǅ�=�6�􊤻~���&V����=`��>k�>Â,�݋���O��I��N��=������� Ed���O�b�i;��ӽ�a�zV!<o%;�?���'��\Ծ�T��A�=p���B>c �>��>���>��W?TR+?�C�<F��c�r�0�$�h�'>�}�e�Խ?&ʾ*7������Ⱦ���Ov�n������޾|m;�y�=��R��O�����zw�H�b�P�:?���>9��3�(��l׾y��3�ؽݽ	�?����G��b���~�?��a?_A��1�b��r�$ŽÚ�r^g?=�K�w�"�S��j>�`�z�< 2�>I�{>��;��1f��"F��w1?]s?U%��t���4>���+>$=�(?�c?p��<tb�>@H?Ķ(��]�:�K>O�>�z�>4q�>��>\�,����?S?W����������>R���!�w��L|=k>>���p��VY>\s�<��$��S�� \7<](W?9ҍ>�)�u��������==��x?�?�G�>�tk?m�B?�ǣ<�x��`�S��.�ʸx=�W?:5i?��>�ف�TDо>D��/�5?k>e?rN>��g����v�.��!�9?��n?9X?p���(g}� �������)6?��v?s^�vs�����G�V�g=�>�[�>���>��9��k�>�>?�#��G������yY4�%Þ?��@���?�;< �Q��=�;?o\�>��O��>ƾ�z������>�q=�"�>���{ev����	R,�b�8?۠�?���>������@*>U�֮?i�?$���K{=��>�J�U�j�W��c=�w>>�H>_C������8���#�D>�������e�U��>~&	@�t�=%�?V.���ҿ$�ݿN�`�����P��٘>���>�i�>�7�1���4d1�>�.��R^�|���*,�>�L>u>������o�z��R8��x��q��>����=�>��Q��=��x��Jl<⤖>/�>S�>Rv���������?����Ϳܾ��@�k�V?#ٞ?ꋅ?��?@�m<�n��rt�g���G?�]t?��[?,���#W��!��j?3_��EU`���4�UHE�lU>
#3?�B�>(�-�`�|=�>��>�f>�#/�n�Ŀoٶ� ���D��?ى�?�o�Y��>h��?Hs+?�i��7��g[����*��K,��<A?�2>!���m�!�Z0=�{Ғ���
?7~0?�{�\.� �_?p�a���p���-���ƽ~ۡ>&�0��f\��O�����Xe����Ay�v��?6^�?Y�?!��� #�c6%?��>Ý���8Ǿk��<g��>Z(�>V(N>N_�G�u>����:�k	>���?�~�?$j?��������9V>��}?()�>�?π�=I`�>�`�=P찾,�{h#>�-�=�>�f�?�M?m>�>�<�=Z�8�e /�VF�ZBR���x�C���>��a?�L?�Nb>�	��_2��!�jcͽ�W1��	鼏P@��=,���߽85>��=>�>�D���Ҿ��?Mp�9�ؿ�i��p'��54?/��>�?����t�$���;_?Pz�>�6� ,���%���B�_��?�G�?=�?��׾�R̼�>>�>�I�>>�Խ����Y�����7>.�B?Q��D��v�o�x�>���?	�@�ծ?ki��	?���P��Va~����7�d��=��7?�0� �z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?TQo���i�B>��?"������L��f?�
@u@a�^?*z�Ͽ����=��M���ٖ=���@>�o��@`=k�=�����1���>��>�.o>�A>#S2>ٽT>S$>�j��e�#�u��`���7@���'�Q�S��������b�������ٷ��"!���眻:_���(`��r�㷖��s�=ƟT?nR?��o?�� ?���|	>_Z��n��<���ԅ=6p�>�02?�~M?�#+?[��=uМ�TMc��΀��s��'G��s
�>#�H>;6�>ݸ�>��>3(X<�^Z>4H>��~>���=�<�_"��� =�RJ>�Y�>H�>��>6K>lw>T���@����)^��4���yE�v�??Q��8�����Ғ�p�(�F���h�J?W�>�}����ӿ\����Y?�B��$������=J�1?/�p?Ggo>�)��	�ܾKi�>.�<r��z �>3��=U"��G=��߈�>(�>�xR>qto>2�2�JE8�ѫK�^Ĝ�Kf�>[�4?�$���6���j��HH�;�ھ�W>���>��%<��헿.fx��>r���=հ4?D��>�1���B����s�ٕ�ZnY>L�x>�=J�=��M>
�w�N롽e�"�u�a=\�>�lq>�4?�.�>-�>���>ψv�P�~�>��=b��>��6?*7?�幽�����P����d��|0>��>��>	�>�'Ž�ƪ>vm�>%]w�v��;1Tc�ke��䂛���>�j���8��/�3Y�=��U��Q>h�>&L�Rރ��k�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>zx��Z�������u�p�#=R��>�8H?�V����O�d>��v
?�?�^�੤���ȿ4|v����>X�?���?h�m��A���@����>:��?�gY?soi>�g۾;`Z����>һ@?�R?�>�9�~�'���?�޶?֯�?�K>�Đ?ht? j�>�H��W�/��6���R���f^=�k�;B_�>�P>(,���;E��˓�9���j�c6�L�\>'�#=��>;�罄i���հ=����m���	w���>}Rq>��H>J��>WV?D��>Ap�>�"=M��)�������b�K?���?���o1n�7Q�<���= �^�%&?HI4?�~[���Ͼ�Ө>	�\?\?�[?Me�>(���=���翿~��u��<��K>[2�>�G�>���KK>k�Ծ�0D�p�>�Η>�(��TAھ�-�����BB�>Uf!?��>^Ԯ=�@!?�&$?�h>�#�>!B�@����)D�� �>��>�?�~??/[��	{2�t���_&���X�A�N>�:y?6l??�>���͚��ϭW�
<��R����K�?�qd?c�ս�V?��?��??��A?��f>(��?BӾ].��g�v>hg?#0�-@A�bG&�4���	?}?b �>�c����ѽ6���xr�	V�� �?�^?('?-w���a�f���{�<�����J�f�;'W]�-�>�>-��G�=��$>��=ʼ]�}�4��<#ɿ=���>�5�=~+���~�=,?�F�;ԃ���=�r�_vD��>�ML>����^?�f=�<�{�t���y��eU����?@��?Di�?lᴽ�h�(=?@�?"?I�>�C���u޾��)[w�уx��u���>���>zn�������MF��ƽlp�;�?j�>�\�>*��>�w�>�1�>�����0�Ͼo���j3x�� =���H�l��'.����P��%�&=��Ѿz\��J�F>�߅��1�>Q?)I�=��>U3\>��=e;�>z9>�0>��>�̽>|T6>K��=%��<& E�3KR?X���B�'�.�辫���41B?�qd?�/�>[�h�䈅�V���~?��?�q�?]:v>~{h��*+��n?c@�>'���s
?�i:=�T��<�<�Y��8������Ѣ�>]׽#:��M��wf�kj
?I.?9#����̾{,׽^��x�m=;Y�?V)?p�)���Q�z�o��W��CS�g���#h�����$�ƅp�3���_^��R����(���'=gw*?*�?�{�8�?���?k��?�f>���>��>�>��I>1�	��1�Z�]��'��僾b��>�:{?���>�P?Ǯ1?b^D?�>?#�>/2�>���)I�>֖<	�>v�>�k&??y�0?�*?d];?�0�>\?��Z1����ݾ�d�>��?��
?0�>��>���@齅k`�A�f=�ͽT�����q�uE���Ž�y����=�˓>�k?���]�7��4��)gn>�2?�	�>���>�o���v�OG%= �>VR
?��>� ��>s�������>>�?����#r�<*�">އ�=
z����;p�=���;V�=��~���!���y<���=A0�=�#/;��H<sv<�~8;�;a<��?�/"?�"�>oˆ>��p�Ϭ�	�ev�=�k>J�S>s)">'j۾���������[g���_>�Ѝ?oy�?4,�=~D�=��=I1��	$�����b;��;�R?mA?��R?K��?f�;?��?M�>�a��$��O���<���?)h+?|1�>d�%��
��7οS�W���?tW??O\ܾCv��h	�O�R�r�>�+)�ou��N����������B!���L�5s�?D7�?EE�����s¾
c��$���=�w?ݲM>8��>�%?�<���s���
��O�>��m>�i?m��>U�?��?�F?3��=��]��A���ء��}��A>b� ?k�?�;�?ƥ�?��u>��<�앾O1��2����mJ>ߎ��͙���>��>y�?-�>O��>N�l��p�j�ż���>�)�>���>�#�>h)�>�9=��G?���>Ϣ�������������'��u?�R�?��*?�
=2N���D��y����>a�?8ի?�&*?2R�tn�=Oܼ-��h�q�yη>Pk�>�)�>֑=��:=�x>L��>�W�>+T�<�nJ8��N� ?�kE?pǿ=��E����u�ȣ�>�!ľ�Ń�KD>��P>��,�����p�2a��"���jj��L[S��	=���x����>2>�>Y7C=�|=>iK7����aϊ���r>F�>������O?����缴�K�Mh��Ž��=j��� ��<~?�mH?g�%?1 9?`K�>M:>%�A�sZ�>ΰA��?�!%>M���Ǿ�!:�x���b��LHʾ�|��Ik�[?����>��.���&>��<>6�=��;�m>ы�=�P�="��::��=�f�=���=��=���=��!>Zc7>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>4 .>\{ >�7R�e�1�
�X��@V�A�Q�L!?ͬ;�ΞǾ��>�e�=>�ݾ�`¾�ǋ=��A>D�K=i#��Y�}J�=������L=��x=��>��1>dl�=CI���=x��=�_>��a>YB̻[~]�0�3��lN=��=��m>�*>3�>IB?<7?ci`?u�>�+�-����\���9�>7�>r�>+�:=�q>���>�l8?�W&?%[/?Aʖ>��Q=D��>�>R����Y�%ҾG�ս��>rӊ?4B�?&f�>� W����-9�T�E�#�+����>��;?��?7��>���sD߿zh1���9�jp��w����,��O�n����iܽ��<�p�.������k�>���>"[�>�x�>�p�>��s>�L�>z*�=b��=���<Q&T=w��=n漛�>N���μ�`�:5dz<�s���d��)Y��t=k����=�Q	>���=G`�>�0>u��>4��=C���w�4>�����K��=���LC��c�Vq~��-��)=��2:>�;I>�g������n�?-�X>\f8>�V�?�lv?��>�����ܾ����$a�.b�կ=��>�0��7�<�\�	�N���о�®>t��>�y>,/>-�M�</���=����� #�>I��~K���s��W��א�~���Pw�ٴA���?�U����=�~x?k%Z?:��?�~:?��Ƚԧ�O�p�� $=�qZ=<�W��t���0y���A?�)?Q?�*���%��J̾*���ܷ>+BI���O�m�g�0����˷����>������оI$3�#g��k���A�B�Jr����>��O?b�?�8b�SX��YTO�k���*���p?�{g?��>�J?G@?&��Cw��o���o�=��n?V��?<�?�>ʭ(>�F�WT�>��*?Y�?M�?�e?h
��#_�>�5>H��=]�b=��+>$�T>OO;��Pp>�?,��>[�?��4�0�9���%��4���þ�n���c>)�v>O��>l��>-P�`�:1��ǉ�>/��>�U�>�`$>�Mh>�\>��žVX�
�?(�=�}p=�?wޝ>��o<e�k4@>�О>�����G�����e[>��A>����M�}=� �>�ӿ��?��>D�"�8��>�᜾�0P�M�>XT>q�$���?
T>a#z=�[�=�5K<g�/>� �>�M>�FӾ�}>����d!��,C�2�R�!�Ѿ}z>]���J	&�����u���BI�yn��7g�^j�?.��0<=�HϽ</H�?Ⱦ����k���)����1�?�[�>�6?bڌ�����>���>�Ǎ>�J��Y���sȍ��gᾢ�?��?��c>�j�>�W?l�? Y0��93�6Z��fu�w�@�0Kd�VT`��؍�ك���x
�@}����_?��x?T;A?;&�<��y>ɠ�?A�%��揾b%�>�/��Y;�P�3=\p�>�a��^�`��Ӿ3�¾����F>��o?{݃??��U��	&���0>�<?N�2?�;p?2?��:?����$?	N>�?"�?�Y-?�2+?��?�{">� �=��9�\=9������Qn��4�Ľ{`��LB=���=����<f�X=EN�<��]�P����:3b�3�e=�cA=>ݨ=��>��>",O?�<�>�m�>��H?Js,=i���ξT,?�G�=�=����Ed��F��d=�dt?�ʪ?��}?�S�>1 R�,���rR>�&?���>`C>>W�D>;��D]�:��=C��=�;�>�CF>�N;�c~��j�~���a$I=Ӎ2=���>��>�P���.>]t����~��)t>?�H�������U��mE���2�tTs�p�>bcG?N�?[@�=��4�v��Cb�{�+?x<?�gI?U�{?���=�վE(8���J�t�"�L �>�1<�!�_���w��{�:� X*�?�d>fQ���Ŵ��5>q���.꾣�i��XJ�sz�]�X=R]�3Z�<��Oþ�dS���=��=p������tΐ�MЪ���H?��=ɜ���(O�ᡵ���>��>ٺ>���;����D�>�����&=���> xj>�R�<������?���	�T��>��G?�e?�x�?U.F�>�j��S��X��̧�1�T�{�?���>���>yM>� �="�վ����9g�P>��K�>)M?=(Ծ4�:��Y���U߾VY=�LD>��>�4c>��?ŕQ?Y-?��q?Ӑ4?^��>��>�Gսk��f(?N@�?�1�=�p���'���4� `A�c/�>-�!?�3��E�>?�F?�}&?��Y?K0?�>����r5�*��>d�>$�P��i���^>f�E?/�>nIQ?9�?�H>�;4����������>{��=�4*?Q#?_D?�q�>,�?Q��;wZ�>ri�>��?Gʎ?�_s?m=9b�>w�?��?٨�=���>"��=sf�>�_?n�q?\ZL?j�;?!mT�vؽ;��)5��񿶽���^�;��&=��ʽ1q=:�޽6 >�Q>�Ql��	��=��Y��}����=��>A�s>O����2>��ľɕ����?>���S��������9����=��>,?���>X�#����=��>���>����'?{\?Uq?x}D;�:b�7ھ:nJ���>��A?.y�=N�l��y��%v���f=�0n?��^?^ W�����O�b?��]??h��=��þz�b����f�O?=�
?3�G���>��~?f�q?U��>�e�+:n�*��Db���j�%Ѷ=]r�>LX�S�d��?�>o�7?�N�>.�b>$%�=hu۾�w��q��h?��?�?���?+*>��n�Z4�i.辊�L\?WB�>G���S�?�;m< ⾓ှbz��I�ھ����	���������@�#���n�������=�?ݏx?��f?G�\?"� �7�Y���^��rs��W�a��+���=��j>�	{B�~�g�(C�g��(#����8=*.Z���F����?��,?m��A�>b'z�����ߴ��-X>�{���D��p=C��Ӻ�<>�N=�D�c`ֽ%K��g?�W�>��>��B?�rJ��%8��*.��6���k�>@�>�ޑ>���>[C�:�7�fS��<��A̅��U�(\v>�oc?��K?{n?/� �D�0�lP���!��9�! ����C>��	>c7�>�U��Y�Q�&�/>�Y2s�{���� �	�1�v=��2?H��>k��>,͗?7�?��	�����Lx��{1��b�<(#�>o�h?��>���>'wν�m ����>��l?���>J�>����pZ!��{��ʽ�$�>�ޭ>���>�o>��,��"\�fj��<���%9�>n�=ڨh?���H�`���>KR?Xw�:��G<�x�>�v�#�!����+�'�6�>�|?���=Ơ;>X�žq%��{��9����,?(9?#j~��G�N��>�< ?x.?@�>e)~?Y��>�趾$FX�A`?��X?�GM?)�F?<G�>�@�=����rj��#���=��E>F�L>�q<�7%>��ӽ��v�':-�>�<=�>�Ɔ�Ž�8�4���r��<�S=d9>0�ڿ��J�KNپ�W��5񾲣	�{ۉ��q�����	�@�������Z6v����9��U��a�����as����?T��?YՓ�����@��(��V���đ�>�bf��y���h��Eu�g���U�޾�7��� ���O��h��f�ѐ,?��@��п�~��ω侼q�>H� ?6މ?� ��B�V��a$����=L�r�mi	>c�ξӟ���޿��.�"?���>���5P;��>���-d>=mY�>HA�4�|�� |��_O?� ?5?J���п�����;��`��?M @�sA?��(����G+[=B��>hL	?��@>y�2�����1�����>�?L��?��J=�W����ke?r<FF��XԻFg�=���=;�=�����I>��>����pA�M�ܽ��3>�d�>/� �Ri�6$_�!i�<�#]>zAֽO���0Մ?�z\�f�#�/��T��V>8�T?�+�>�;�=i�,?
7H�K}Ͽ��\��*a?�0�?Ϧ�??�(?Fڿ��ؚ>��ܾ �M? D6?���>�d&�4�t����=�$�I�����㾗&V�6��=H��>�>%�,�k����O�VD�����=5��Izȿ_�A��n)�jҽk���7��% �:�˾��>����g�@��VE=��y��.��fV>��>��>�X=��4?}�??��>�V>���=ڙ��͹�8XŽ�[��5�y�=��:kv���������ٟ�=1Ѿ:p���׻�еK���*��VS����ީ���H�޳g���?|)�>c�+J�A�=k
+��ľ'ڤ�k�o,��a&������z?��.?3�g�M�L�� ��^����%Q�~Z?��>+:���޾"y���(����!>��>���=+��>�7�5�0�T�0?�?wܼ������a.>=	����,=@�+?e� ?��<��>"V$?�?(����`>�;>��>���>�E>����νS�?�R?����V[��nڌ>b���>{���c=�{>�G1�8��t�Z>�f<5e����r�[/����<�(W?���>��)�� ��]��r��C�==��x?��?1�>'|k?��B?Z	�<{h����S�����w=m�W?z+i?��>r���
о��5?�e?��N>�[h����Q�.�fV��!?��n?�\?Ý�u}����|��wl6?��v?�r^�"s�������V��=�>^\�>���>p�9��l�>8�>?n#�KG��ߺ��}Y4�Þ?n�@i��?�<<#�Z��=E;?5\�>W�O�?ƾ�y������
�q=i#�>�����ev����R,��8?���?��>��������>���� V�?�d�? �X��@p����Y�p�L���^Լ=+�=|� =�m轋J�]�2���ʾ�Z�U6����;��?>�x@�a����>�A���iȿW�ԿA�_�pV�\����?q��>"���V�6>C�rr��@F���b��S��QR�>��>C���W㑾��{�g;������>F����>)�S��+��X����7<�>��>߾�>r$���὾g��?�h��c8ο�����űX?�i�?�o�?m?@8<��v�\�{�V��G?}�s?/Z?H%��$]��M8�$�j?�_��eU`��4�HE��U>�"3?�B�>B�-���|=>���>2g>�#/�s�Ŀ�ٶ�+���X��?��?�o���>j��?us+?�i�8���[����*�'�+��<A?p2>���D�!�C0=�XҒ���
?P~0?0{�`.���_?�a�N�p�"�-���ƽ%ۡ>8�0�|`\�"������*Re������@y���?e_�?��?6��1#�	6%?��>�����6Ǿ���<���>��>�%N>u_��u>]�F�:��i	>-��?�}�?Ef?,��������]>�}?"�> �??��=˃�>��=G�� ::�p�">4a�=��>�ͻ?g�M?�9�>���=��8��,/��LF�~DR�;,���C��<�>��a?znL?�*b>����{3��!��Gν˳0���弄@��#*�Z޽h�5>�=>�l>��D��.Ӿ�?���+�ؿi���1)��!3?-�>0�?�����u�O�	�*�_?��>"��1L��.��(��	X�?���?C�?��׾	C¼s>�R�>� �>�ҽ����=��2/7>��B?��w>��&po�\�>v�?�v@��?��h��	?���P��Ra~����7�m��=��7?�0�&�z>���>��=�nv�ݻ��V�s����>�B�?�{�?��>!�l?��o�M�B���1=8M�>ɜk?�s?�Ro���a�B>��?������L��f?
�
@~u@`�^?(��Ϳ�:���h߾a�˾v�#<�[���>,��4��i>	<�����">{Ω>���>s��=���=�XJ>�/>7�>�����u%�����2����~R�WPE�<�&������'��9ԾN�
���(�Ƚ�I=V��B2��	�?��76�ͷƽ��=�2U?V�P?n�r?x?§��]�>�����<{���ю=�s�>�-0?K,K?��/?j��=b⚾�d�m�}��Q���ր����>��A>0��>�\�>�>�ុ�H>�?>�Mv>.��=T�;=�tL<���<��J>«>�V�>%5�>��q>��>�n��q���Z�5�-�N����%&�?[i�=�m��^����ʾ�/C��SJ=,+? ���;צ��7Կ����~lP?����6<��
q���=�=�>�B�?1ɀ>w/k�M������>��.�ɾ���>���t?ҾH�i�8��>Qp?`�e>�qu>.f3�u�7�V�O��9���Y}>.�5?�q����7��uu�ϦI���ܾ[tK>J׾>IQ%����薿�}}�xh��q=��:?;�?���f鱾"�t������R>Z>��=�ı=	�L>�+a�k�˽��I�pa9=n�=�]>�?�J�=u�%>�J�>y�򽍶E���>��=βS>��<?��?�;��׽-��|%�����>Q�>�Z�>��P>�p#��2>] >iE�>��s<*���"�n���H�=�r�h�`����e��<�D��|&>k\7=��"��'X���E=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾNh�>}x��Z�������u�h�#=Q��>�8H?�V����O�e>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>:��?�gY?soi>�g۾=`Z����>ѻ@?�R?�>�9�}�'���?�޶?֯�?��N>e��?�w?m��>i�7��	/�i?��͘���'=�tn��S�>t�I>q˷�)78������f$c��h�F:>���<���>�(N�̬����=#���O��>]Խ\��>��>��m>��>�l?֝�>w"�>T��<|��9�z�}᪾��K?���? ���2n�XS�<䟜=%�^��&?OI4?Gg[�?�Ͼ�ը>̺\?c?�[?'d�>$��G>��"迿�}��T��<+�K>4�>�H�>c%���FK>��Ծ�4D�gp�>�ϗ>
����?ھ�,��oe��,B�>�e!?ɓ�>UӮ=Ι ?��#?�j>2)�>�`E��9��8�E���>���>�H?��~?��?�Թ��Z3�����桿\�[��:N>��x?�U?c˕>.���䃝�iwE��BI�����D��?7tg?T�@?A2�?�??w�A?�)f>���bؾV����>К?�ս�=��u�lԽT?��?d��>B�ͽ�bo�63���1��2���u�>HR^?��*?&m�U�f�<.���Ē<�ɼ]���8D< ��<M{�=m�>�4���=A�#>#�=g�k�C�7(=ż�=Տ�>�7!>9J��i+��:,?PK�\�����=o�r�tuD���>��K>(���؝^?�^=�n�{�����u��b#U����?.��?sg�?ʹ��h�9=?A�?"?$��>�6���޾yq�ňw�j�x�j�0�>���>�n����"��������I���ƽ����� ?bߪ>���>���>D��>���>U򨾬v*���¾}��T���� ��b=�oB����GS¾\�����=��Ⱦ���}�E>�b��K?���>�OC>�xa>;n> �	>�>	#�=L��>��>�i�>�h�>4i]>�c*=�\j��KR?����^�'�o�辱���72B?Srd?�2�>�h�H�������?���?Rs�?1;v>Nh�g-+�n?�>�>����p
?4d:=����S�<�R�����@D���&�u��>�E׽L :�M��tf��i
?/?L����̾�6׽݉����n=M�?��(?�)��Q���o���W��S�����4h�Jf����$���p�=쏿�]��#��H�(�C^*=��*?E�?�����@#���$k��?��hf>��>��>+޾>�vI>��	�\�1���]��L'�S����H�>�T{?�r�>y	L?.4?��F?=FI?�h�>+��>)≾���>�Ć=��>���>�J(?��?#�*?CP?3?'j�>�W�����@�¾:B?3n ?g�?Ն?���> �¾����oo�=h�߹yTd�Ɩѽ�W7<^���� ��ý�ҡ=Z�}>�X?g���8����� k>q�7?,��>���>������3�<��>��
?Z>�>����0vr�^�-W�>��?I����=��)>���=Ea���`ֺV�=0������=#ׁ�.�;��<�y�=���=as��0���:���;�4�<v�>��?Ꝋ>�^�>
 ��̪ �ܧ��կ=�Y>bS>O>s9پ�{��c"����g�nMy>�s�?xv�?�
g=���=�D�=�x��@H�����5콾A�<;�?�5#?�=T?s��?�=?(c#?��>.$�.J���Z��t+��ڣ?]11?㐻>�r��	���ӿ�;O���??B*\?���h���+���./-�)�>v<!�����u6ǿ}���F6=�Y���V��|�?��?2V��m%�MB��j���ھ�_?��>�>�?�P.��S�S��-��>(Y�>$��?���>T�j?B�?��k?>KI>��8��y��0��Ug��}�>:<=?�Fu?��?do�?{�?��w렾Gj$��p���:�=zZ)��l���ٖ=:+
>�> ��>��>���=��=��O��R���">^h�>a��>�6�> 2�>� >�U >r[H?���>�l�����ϟ��|��2�t?+��?+?�-=���B��@���M�>��?_«?u*?ۡD��.�=�몵��v�V��>�8�>�L�>6��=61=�>{T�>�>�d����(�5��'�t%?�(D?�v�=���v�v��,þ�۾�Ǔ; y��\j̾��'�)�k�=H!��+��=kT��t+ƾ��-�&���O�!-7�������>_P,>BgS>�FC;A[=����`�����h�e>��=�
�<|Ob<�	ҽ�v۽���<j�.>S=�<��==,c��5~˾��}?#;I?Z�+?��C?��y>�J>��3����>tH��JB?>V>��P������{;�X���A��9�ؾ)i׾��c��̟�BL>�=I�h�>IS3> @�=�؇<��=!)s=���=N�Q���=v�=�S�=�o�=���=��>�U>�6w?W�������4Q��Z罤�:?�8�>h{�=��ƾq@?��>>�2������yb��-?���?�T�?<�?=ti��d�>J���㎽�q�=B����=2>u��=u�2�R��>��J>���K��G����4�?��@��??�ዿϢϿ:a/>ȩ>T�=�
P�V1�#nK�0JI���l���?�h=�r�¾��>
��=��վ��Ͼ��<;�~1>6~w=!� ���]�?W�=��A��׆=g'<=eZ�>@?>���=�Ž�|�=9�A=r�=�5T>㱊��I��Ƞ�G*�=��=>+m>��>��?o?}�$?�U�?���>|(�]��@ŗ��$>���>P��>z(��T>��>�a?U09?��:?E�>�F>��>�W�=1Q�ю<�������6�ۧ_>��n?#�z?��>��\;�x��'��A1�I�����?׉6?~�?C�>�n
�h&���7��/���~g�=86���?[�T�W��9q��t~���]�E>��>�P�>�F�>m!�>���>X�=�F�>�M�=��<��=��<-��=6�:b�N=�S	=�g�<A~;��<�S�q����0�ԭ��V>_t�<;5�=E�=1'�>t>��>�O�=}���:O2>���P�J����=2ץ��@���c��	~���.��O6��D>kE[>�Cz��^����?XfW>"�>>?B�?��s?1�>?��8ؾ�d���wa��SM��Z�=�\>�;��I;�|�_��;O�"7Ҿ	��> �>�^�>>>�>X��F�a�>*�ԾϹ��D�>��)���[�TcZ��n�����t�Ԉ$��E?������=�/]?��]?��?s?�9�0F��\��=;���6�����걾�v?}�+?y�?����7,��N̾#M���ٷ>�?I���O�俕���0�����׷����>����о"3��f��L�����B�e7r�E��>״O?��?�Jb��P��LO�����\��gj?�rg?�0�>�N?>?�͡��y��n��(j�=��n?���?:�?��
>m,>&�Ӽ��>-8?�q�?�_�?�#l?����>�l�=��&>~?��;�=�s>J�1>3eB>-s?�?0]?Ax��/����z���f��nV<$�`>�>��g>u�&>Z!�=���=��=$�H>��>��>p�^>�>ΦO>�L���|�i-$?��6>�;�>�
?�W�>����V齈B�=N2��E����^�	6�C��:�A=JS*=���=[ >��>9˿P͟?o��>���u_U>:f��l&F�}��>�,>�o;�$<?S�j=�G�>��=�G&>g�>}�?P����Ӿ�;>O��!�.>C�g�R�n�Ѿ�^z>�ǜ���&�����	��RG��մ�޹��9j�H��!=���<���?�$ ���k���)�N���{<?�&�>�5?쨌�禊�}�>���>э>(�������Ե��0R����?���?�Qc>���>��W?	�?�1�V=3��RZ�L�u��A���d��`��ԍ�������
��d���_?X�x?�uA?�0�<^z>W��?��%�c���x��>�/��.;��==���>"Z��2�`���Ӿ�þ�Y��1F>�po?��?�-?�ZV���7�r�&>Q�:?��0?�4s?;�0?�;?��G�%?O}E>bi?�P
?֩0?3i*?u]
?�9>�=�=?��;hgb=���㊾�}ͽ
���S��f=a�p=$����;�=]�D<e�̼1�BO����~�9�<OG+=gi�=��=b!�>%cV?���>���>%�:?�m�x�+��Ɯ��{$?���=M+S�3�k��������U�o>q?G�?fF?�/{>�9�H���>�c>�o2>�VS>�l�>�0����j��/�<D�>��1>�k�=4b����d��� �����,=B�0>�,�>=}>�)��<�(>T����u�>-g>A�P��ݻ�P�t3G���3�IVu����>��K?0?�0�=�g�BÃ�f�d�~�&?><=?3]M?@�}?�L�=�ھ	�8�I���h$�> �<;E�)���q�,;��.�;�l{>ؘ��"���b>�����޾�|n��J�|�w�N=[�B�V=B2���վ�"����=�T
>���� �����ͪ�i7J?s!n=ǒ����U�����A>5o�>��>vq:�k/x��~@������Y�=Q��>7X;>[���I���G�iM�l�>�xL?~�h?0`�?=a9�AJf��P�����Ѿ��+=�� ?�[�>DD?�>�>��=j�侥R���g���?�$0�><�>mC��RQ�"p��i���3��d�>�6?�f>b?/�C?[]?�|k?s�0?u�?e/�>w���Υ��r+?�?q�>]��<��0�12��](��<�>�;?T���)�>�?Z?3?eJL?8?��*>'��:��5͎>�=�>�[�sB���NC> �N?:0�>��q?$jt?�\�<d[I�Q�Ǿ���rU6>k�]>n�*?T�?��?�p�>��/?u���H=5�>p�'?ߖ?��h?Ao>�ʽ>��>���>|p�=�_�>(��>���>�F?�W?MS?K�?(��=<����j��`Q��.�T�Dʖ��ӽ���=\;��E4�<5vR=ty�<V=X>�=IC�<W�>?�2�7	z�#̍=Je�>��s>�����0>��ľ�6��rA>�A���Q��yĊ�zO:�P��=(~�>��?���>�
#���=���>�S�>|��#(?��?a ?�"";E�b���ھ��K���>ZB?G(�=��l�|��J�u��h=��m?�^?gIW����M�b?&�]?ng�@=�Y�þ��b�Ĉ龏�O?�
?<�G���>:�~?-�q?���>�e�V9n����^Cb���j�aж=�q�>/X��d��?�>��7?�N�>��b>f!�=�u۾s�w�>r��?��?0�?���?�**>d�n��3࿕��蒿�@^?q2�>啞���?i�s;�2Ͼ
����'����Ծ�ʗ�����1w������3�&��ˁ�󾸽O�=?�?t?��p?t	c?�"��eg��o\�!���<T�d5�&�е>��2C���@�'�p�p��*]�����:�&=c�b���J��1�?,�,?�G��(�>R쁾x.��¾�P>�]�=��f��=|K����=���=��@�)�4l���I?7�>��>�:M?��D��(X�b+�\N8���پe[>�}>�a�>��>��;E*�G@�5���mo�'�½�v>�wc?��K?=�n?���1�i���!���5�^_���B>�z>��>�vW�����5&��\>�*
s����M���"�	���~=��2?D��>��>�6�??B{	����w�N51���<Y��>hi?/D�>�<�>��νʆ �}��>��l?T��>h�>i����Q!�c�{��ʽ�#�>��>θ�>z�o>�,��!\�Oj�������9�ȍ�=g�h?*����`���>DR?7%�:(�G<䀢>��v��!����	�'��>
x?\��=u�;>}�ž�%�9�{�k>���*?�E?f{��У"�_v�>�. ?5��>!�>_�?�^�>�����t���?��^?�iN?M�C? ��>�VI=�냽|;˽B0+�R =��z>b>��=I/�=�&��m�Q��a =z0�=������<�=,�����<,��<N0>�ֿ��M�c�����~�վTk�񇥾�W4��P���۽��;HA��DS�(нߍ!�#�t���I�O�����o�s��?J�?�����đ��Û���i��A�ov�>��4!ƽu왾���ϯ���Ѿ�\~�B_�T�g��f}�=s�A�'?|���ܽǿ鰡��:ܾ(! ?�A ?&�y?��7�"���8�� >�C�<&.��뾧��� �οj�����^?i��>��x/��s��>$��>��X>�Hq>����螾i4�<��?E�-?���>L�r��ɿR����Ť<���?/�@u�A?��(�����V=���>0�	?L@>D'1��1������n�>��?1�?��L=r�W���	��{e?x�<�F�`�ٻ�`�=�_�==0���SJ>gc�>G��V�A��ܽ��4>�>��#����w[^�J\�<��\>!׽����5Մ?+{\��f���/��T��U>��T?�*�>R:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�ޅ�=�6����z���&V�~��=Z��>a�>,������O��I��T��=+��s�Ŀ�)�'I#�x�9>K��n�3�t��7h=��M=��꾼�e�Rqe��� =%z<4��=)�>�}�>܀>��G?#Wa?���>[>��:��J��A{پ1��;�a�6u)�^J9���ý�=���s������޾Hl+�f�(����Q|2���;=/]�}*������.X�+��A?��>�ۙ��ss��C����e-?��j�=����$徂?��d��r�?��j?�8��=�}��z�I1�=
'E�BO?�=��+�d���p��=�o˾�U��q�>��></	�+�M���R� �1?�X?F���L���R'>ㆳ�<B=�1)?�=�>@�<zL�>��?�,�
��dTP>�4>�X�>���>��>cM���>�/g#?��T?�j����+K�>����D؂��=�>4�%�gK���J>^p�;̧������ƽ�R;EsW?���>��)�q.�D���ץ輯�=l;u?��
?��>��l?i:?@���e��|�S�]��غ=�[?��l?�8>N�\�ad¾����C7?�Pe?[>8�\�d�ܾ��)���
��'?�i?}?�I;�{�|�����*���d3?��v?�S^�el������V���>���>��>3�9���>Ǖ>?cZ#�NB��̫��$N4����?��@Z��?e=H<!�,��=�:?�3�>I�O���žtŲ�%i���#r=})�>|t��Iv�2��u{,�=o8?N��?�q�>�������->Ǥ���y�?]��?/���w�!�߾s�u�_��^�뼈�>�k�>H�<�p�W�����A�:���h0Y��KJ>��@�c�=Pt�>ʢ,�Ԧ��[#ӿ����v\'� }�{	�>���>��>�h��-k��׊�1�_��j�eǳ��I�>V�>ؔ�_���=�{�bo;��៼B�>�a�7��>��S��#��R���z�5<�>>��>�>�0��佾Ù?#W���>οC�������X?�d�?�o�?�p?a�6<�v�y�{�X��5*G?T�s?�Z?�C%�n?]�]�7�f�j? ,���`�ub4��E���V>"3?^�>q-�@=?u>Ƕ�>�>&/��pĿw���	$��B�?G{�?�1�-w�>2��?D�+?�u����H���7�*��,ź?A?H�2>n��S�!�>5=���"b
?�0?���qT�]�_?*�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>`H_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?f��>_�?~�=�%�>#�=�Ұ�5'�ze#>M��=�1@�0�?"�M?D9�>ޜ�=h9��/�IYF��VR�K,���C�VƇ>I�a?�tL?�;c>7O��f2�� �
ν��0���伀�?�la,�=ύ�5>�	>><�>UD��aҾH�?Z��#�ؿ g��w7&��4?�d�> ? ���t��&��
_?LU�>>G��+���)����ܘ�?�-�?��?Й׾��ͼ @>�>��>Fֽ�3���\����7>�hB?�������o�.�>:��?G�@�?��h�	?� ��P��ia~�`��%7�=��=	�7?O.��z>e��>��=vnv�Ż����s���>�B�?i{�?A��>��l?�o��B� �1=�M�>ٛk?�r?gfo�t��B>w�?t�������J�of?��
@=u@�^?u�����ڒ�]2��6������$<>���>J;���
н �=Gr�$P<�W�=�<�<*+��OO>�i0>cD�=k�c>7���H �������z��)M��O�������k*�޽����6��)ξ@(���`���	˾�u>��@�[�q��16����=�T?'WR?�m?�$?i!��>x5�Cz�;�k���=`�>r4?�`O?�^-?�ޝ=Ã���8^�O}��Ф�G���ㄺ>'oI>*��>KU�>��>���<ȦY>{�;>��z>}��=5G�:�� ��Qu=ACV>p��>���>"b�>�_n>p;�>	¿�Oȿ��B�<�z�&D�%�?f�=qɑ�w�����(�;!�t
>��?[}?�p����Ϳ^ݹ���=?1C|��Q��![���$���?�-z?�+�=���<Ԭ��h�>Aݽ�P�\����>o/��)M���=��h>wH~=��e>�Rv>13�b&8��Q�����c}>,�5?2���g:�&u�:H�q�ܾR�K>7�>�]�9�����4���j��s=L:?�~?㑨��]��]^u�A����O>z�^>-<"=�ϱ=��L>�u����,�F��;=T��=��b>RY?�g�=Њ�=7.�>���k�=,J�>}=3>�o,>�+I?wq0?F*�+��œ���X�$}]>O��>kY�>ڶt>I9���68B�?kУ>U ���~��i�:�M!�u	>Ų����?�A�=�B����Խ��>oȷ����Q��Z����~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�\�>x���Y������u�r�#=r��>�9H?�L����O�J>� t
?�?�d�����+�ȿ�tv�!��>��?���?��m��@��X@����>���?�`Y?N{i>`۾�[Z��{�>A�@?#
R?��>�:���'���?>ݶ?�?��H>۱�?��t?T&�>�G\�p\.�����J���[�P=mA&<H�>a$
>鹹�<VC�򒿬D��c�j��y���_>�s$=HJ�>3��>;���k�=����	��:Tf����>�x>Q[S>e��>��?���>U�>�=*=
܁�Ʒ��~┾^�K?���?���2n��I�<N��=��^��&?I4?�p[�R�Ͼyը>ɺ\?N?�[?�c�>D��O>��9迿Z~��-��<r�K>(4�>#I�>�"��uFK>��ԾP5D��p�>'З>�󣼤?ھ�-��xA��FB�>�e!?œ�>?ծ=ۙ ?��#?��j>�(�>AaE��9��W�E����>آ�>�H?�~?��?�Թ��Z3�����桿��[�t;N>��x?V?uʕ>a���񃝿|kE�%BI�F���]��?�tg?qS�/?;2�?�??a�A?z)f>؇�(ؾq�����>�l ?>����@��%������?�?�\�>ؠ���ֽ�h��m�����ZV?��[?1�%?����`������<��V�����5�;R��0�>A>ڣ�����=)�>(|�=��i���5�i�J<��=�Ӕ>�m�=��4������,?3�(�vA��mM�=�Wr�N�A�
�>cKM>������_?�H2��{�#���z	���Y�<1�?	��?+ϖ?���g�f��I<?���?�5?��>����*=پ��ݾ2�o��s�:���0>G,�>B�h���X#��I���{��Rý�� �S`�>ʇ�>X �>F~�>��S>y4�>���&A�21�g���;F�N���:9�&�6����L��*nq�؆�ξZ~��ŗ>�����>��?�!A>��s>I��>0��=���>\��>�x>=bs>�C�>n�N>B�a>մ�=&]�=�LR?������'��� ���x7B?�qd?\.�>�&i�����5��?h��?*r�?�Cv>+h��)+��n?�?�>���Bq
?�=:=��O]�<Y�����R/����	��>�I׽) :�'M�2gf�di
?0?g����̾*׽�����n=[K�?N�(?��)� �Q�]�o��W�S�fq�9h��p��'�$�!�p��돿�^���"��Ǜ(�Pz*=R�*?��?������}!k��?�ˁf>��>�%�>zپ>�I>v�	�"�1��^�LO'�V���Z�>�X{?�͢>��M?D?��T?_OW?VP�>��>~M���|�>��;lӃ>���>��,?z�8?��[?E?vA%?q�>�����߾��ݾe��>�?xg?��?���>��6�	T"�K�N�:��;pUA��a���ҽ�Q�=����!a=�/�=�k�>��?'h��'3��^�\m>��=?���>��>|_��d�|�/@=R�>�?6=�>���mjr����,N�>b��?}��$� =	>/��=)b��ym��ʥ=ۮɼ���=݃���?:��O;;ч�=c@�=���:�Oi<8;	� <�
=5��>r�?6#�>(�>QU��! ������=��Y>t7T>�>^�پ.k�������g�M�y>(��?���?� n=��=a�=�_��;�����>^��\��<�?4#?_>T?�V�?�=?�#?��>��=D��"\��o����Z?A?��>a;�2	�"�ɿ�<��?w�?t�7���[:"�i�M�]轐��>8\�f�n�V��E+T�a���=���Ҽ��?��?~*н����Έ��e��^�j?#��>�6�>�@?"4�,�E�K*���>r3�>Nw�?E1�>�t?�?�yS?���>��E������)��wp����>��m?0��?� �?S��?L�?~��)����+�W��l2M;|9����:��¿=�J�=�>z�?�2�>G}>�H���O��߂�����=`>k��>��>#{�>�ʞ>E˽�L?zp�>�����K����*��iW�=�\?펋?�%?1}>+��n=�8n澙��>�G�?nu�?��N?b�u����=j'%�`��:�ǾNq?>�>1L�>Y��=z>�B>���>�m�>\����F&��� ��A�q�'?#^U?AU>�ҿ政�᱾����ᙜ�����]�I2<�ђʽ��">�+�Ш�����;8&������о����A
�(����]�>�̀=���=�ܙ��ܟ>��"�[� ���==%>q>��O��!�oщ<aɺ=U��=}�=<S�= �a>/��<�\˾_�{?ϹG?9D*?'�A?�ox>K�>&�3�6��>g���ͭ?Z�V>��C�Eܺ�&�7����n��ԓپ�Ծ�Oc�k砾Kq>Q^I�J�>�4> ��=ЇS<#�=R�x=�0�=���d�=��=/<�=���=Q��=w�>*�>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?��>>�2������yb��-?���?�T�??�?;ti��d�>L���㎽�q�=E����=2>v��=v�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>���=�[�=i=�_�!���v��*�t��P?1�P������>>�ѭ�q���.��={Q>�{�=C�X�-�7�~��=�^߽ChO=��=&��>�'�>�&�=���R\�=~ė=�M>��b>+���,���W<#+0>�"k>��k>�?*>CZ�>v�$? �;?Уx?���>P����~�������>�q�=H��>�C>d>:��>�H4?\OC?fb9?R��>��>7)�>3ݮ>�m4��b�o����׾du0<}��?�[�?F7*>�bQ��څ�Wh�L�)�_�o�+^
?z�6?ߧ?\Q�>S2��w࿠&��*��Ҷ�����=��}���a���Ƽ��,����{��=��>p��>w4�>>�j>�*3>�O>�3�>f_>�$=��q=e�<=�;�{�����=^��;�={䡼�3��G���}�6���⻆�<��!� ��<P�'�h��=���>�@>i��>���=k ��L/>(���Z�L��Ŀ=C��_*B�N3d�3H~�f/�-Z6���B>�7X>]��*3��=�?��Y>zo?>߄�?HAu?0�>! � �վ�O��J?e��ES�Ÿ=f�>��<�Oz;�MX`���M�xxҾo��><�>G�>�b>�.��I<�x>�=��ݾ�H;��#�>�g��,F#�����n��ˤ�𺞿(i���ϼ6�<?}������=A�z?�wH?�%�?&�>/��[rӾ�j>�g�J5P=��
�� l�9\ݽ��?�%?���>]m��s8�# ��T/V��'�>	�~���-������#��z�<
_��e��>����0޾�;9��ꈿጿ�6P�P�#����>cB?��?��i��b~���]��F��v�i�i:�>�N�?nY�>(��>,2�>��;�}��IN�����%F?��?@��?�j>�&#>�q���H�>o�
?���?5�?=Kp?�*����>� 	=�`/>����=s>�=��=��	?2�?�?��p��)��(� �͠�I;<�e���^�$=�
�>��>��>�=MX</��=@#n>3��>!�>��Y>Ҕ�>�|�>����c?�>ſ{>�@6?��>�ق=����=_�>+�ѽ�Zƽ��Q�ɦ�<o>�>�-�=��;(��>
j��)��?�J�>gZ���p�>�7Ѿ)���Y�>���>�U��^8�>�T>.ɓ>���>d�P>�=�P�>�7�=ƥӾʧ>��7V!��C��RR�S_Ѿu�y>�֜���%�Պ�������I��̵��z��j����y�<��Ȼ<7#�?i@����k�w�)����S�?P�>0V6?[����i�� [>JH�>q�>B��Qi�����pcཱྀ�?���?Y<c>��>��W?�?G�1��3��uZ��u�@(A��e��`�o፿뜁�
�I��4�_?�x?6yA?�X�<:z>.��?�%��ӏ��)�>/�';��@<=�+�>�)����`���Ӿ��þ�7��HF>��o?/%�?�Y?TV�	����^>?�F?��@?��~?�>;?��3?)'�&�?��1>@�?��?��?"?�+?�8X>ݑ�=��d<��=w���R�A�ǽ[��ϑS�;m����=P��������<)�=)�<=H=_������������A=Te�=p�=�x�>|o\?AQ�>t!�>��9?ά���'������E#?V�<�(������]d��|ӾMs>��l?�b�?ޠW?��>�;���P�a�%>C��>\�0>���>uR�>�,��DT����=�~K>�JA>4@n=�����
�GQx��R=;X>��>d�}>Ś����(>?��0�y�Ve>�'P�N׺��tT�ŒG���1��%v���>��L?�?�L�=�~��<����e��(?��;?Y M?�?��=:�۾E2:�F�J��<��:�>#ż<���Ң�V�e�:�xcM;G�t>�m���Eݾ	)q>������R�s��O���C���>sG#���È2�El��Do��Q>�6>c󾡁<�d�������N6?dzK=�]X��PY=q���^y[=`�>=1�>���<����J6��Ȣ���	>
��>�0�=�
�K���;S�+
�^��>J�X?-nj?�J?����o�'�N�'��@���!<)/?��>P>?7'E>�=ە��R_
�#i^�o:G����>g��>S���C����������^>k�?R�^>+��>��I?G�?�y|?K�'?���>�ǰ>��L��$ξ�T&?Kd�?h�=s�̽�ZR�f8���E��9�>;)?�C�8��>��?��?#V'?��Q?��?��>�� �m�@�52�>�>��W�����4`>�QJ?sV�>sY?ݯ�?A�=>��4�x������K0�=�>�O2?v#?F�?�?�>��>'�����7>$��>*'s?���?�o?$���A)?��z>�)�>�-<I�>��?Lm$?(Gl?w�i?��2?�}�>��<�@�N:����Pn{��z�=�O�m=�������-�3l��Ig<�e�����yڵ����	r=�b<Z�>�t>Oߕ��U1>��ľ]3��K�@>�6���D���Ҋ��>:�9q�=��>F
?�Օ>�#�]��=E��>�!�>H���%(?E�?	?��;��b��+۾u�K�v9�>5�A?K �=7�l�f���iv�i=��m?z^?YW������%a?pc?��ܾ7�^�þ�
m�^��D?��	?���<��>��?]�m?���>��K��p�}>���[��D��=�>�^�ؖX�)u�>v�5?QV�>}�Y>�=;F��4�f�	��m�$?�?�?�Ͷ?��?�m/>b�e��ٿ�~���K���^?���>@��� #?����n�Ͼ�O���(��=�W�����=C���x��̲$�;ރ�q׽l�=[�?)s?J\q?��_?ӳ ��d�2^�H
���kV�)��%���E��'E��C���n��b�|0����e�G=��T��HE�Qc�?�O?Qy=�v �>��Y�2���"J��aۊ>� ����=�>Wo��\�CF�=�Y>�7�ݽ�ʨ���?���>$��>�>B?s�e���L���A�Sg�����{��>r8�>}�>�\�>E�=L0v�T�޽��Ͼö`�p��W�>�}p?�LA?��o?>���U4�L��(��	4<�$��f�J>*ď=��>i�<�<��=�;�p�r��>7��g�Yh�(�J�n�`?)�?<Ȼ>���?	?�\��5����PC�ˊ��|�>Qgk?���>���=�T��""�{��>�]m?֏�>���>�f��\�!����}˽��>|�>��?v>��3���Y�ۍ�䏎���:����=Z�h?������S��t~>%oK?��;Ղ�<���>���,$�������q>��?߮=��a>@Xþ^���Oz�(ݍ�Ԡ(?e=?y����{(�SC�>�-"?�c�>���>7�?��>'?���`";RU?L�_?Y�J?J^B?�I�>��=�!���RȽKC$�$26=�Y�>�[> �q=L�=�Q��\�b�>>=W�=�μ���}��;_˼k�1<z�=<s7>ʢ޿��W� ��2�������;j���=>}�ľi�'����o�0�{���c�#��=W}�[���������~H�?9��?�!��^R۾�8��pۑ�`O��L%?��Ǿ��X��N����P��������Ǚ��p��\��b���?p�ށ#?����9qƿ�ꞿm�#|?�;?rE�?W���U$��=�v�#>��=9 <�'��X�����Ͽל��g?�U�>z�����>
L>ꠃ>(�s>:��g��9:!=�# ?��/?��>0o���˿�y���ko<ł�?	@y�A?��(�f��^=��>L�	?%X?>d1��+��E���Q�>�8�?V�?��S=HW��e�Ke?���; ,G�ڤỏ�=L�=��=/g�tJ>d��>]��r�@��v۽�?5>�c�>��!�5*�;^���<��]>�ҽ\���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=��E̿�|�U`!�:A6=V);i(�|����ϝ�O�ؼ|����<�"�����=q4
>��?>!�>��I>�>�3^?��r?Ǟ>Z<�=��L�x|���˹����=NA�����/2�����x��V]�o�ȾR��~�e�����2A��M�=KpP����K %�,�k���E��1>?�2�=��Ͼe2O��<ݏ׾�H���/p;,�Ž�2Ѿ�$6��h��6�?HBI?l=~��;O��U����{���#W?۫��C��������=4�׼� J=F�>C�d=����C��O��r0?Fs?�Ϳ��現�U+>�0 ��U=Om+?�3?�M<�s�>Du%?-{)��߽3O\>C�3>]�>��>��>"&��-�ٽ�?-�S?�� �搜��p�>�����({���^=RV>�5�%�nM[>���<=���B`�A�r�<�$W?檍>:�)�� �,e��x���<=��x?&�?YN�>�sk?|�B?���<o����S��"�;w=
�W?]!i?�>�m��оV�����5?j�e?��N>�Wh�%����.��L��*?��n??Z?D֚��m}����
���d6?�ׅ?g�p�)���fu0���ʾ�?.}?�e�>i$7����>�:E?*�0�����ե��#vK�tǆ?�@�m�?t>�K��,u�>�?dc5?��n�G�D�����яL=����2`?��7�f���a���K�Lf�>���?�6?�C��/ ���"> F��"[�?~V|?h����������W�����cj>dN�=Tޜ�l��K۾V<�������D=���n=�Ǘ>��@� ���?@犾z�IܿDX�i�ռ�ཋ�-?wZ�>so��]{m���A��W��ܟA���A�@�ɽ�N�>��>)���~�����{��q;��U����>��z�>�S��&��5�����5<"�>ݭ�>��>^5���뽾�ę?�c��@οF������.�X?�g�?�n�?�o?9<��v���{�����-G?ʉs?Z?�}%��>]�z�7���j?p���x`��4��PE�k�U>93?�>��-�.Q{=iG>���>��>�-/��Ŀ]Ŷ�{5��j�?	��?�U��>`s�?W�+?�I� =���|��l�*�M����A?�[2>����!��=�N���'�
?��0?\-�x1�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?Y �>�ݏ?Yy>,�?� �=�V�������E�=��o;t�:? I?��1?�|<I��l�.�bE�
z5��پ0���>j~l?��J?���>�1�kE�<����o��6q�I`�<���	0��s�d�L�<.�T>N�>��ҽli�b�@?;�J��p�������9�p?�
�>Y(}>H��k0�AC��Jw?*�>5�R�K���8���7=!�?�<�?��?�F���~�/p�<ԅ�>BA�>�;>�K��_���I�='^?�ռ��|�I��{!l>��?�4@pب?��t��l	?&������ �~�����F3����=R7?���ow>�v�>���=�*v�@˪��s�Sݵ>u6�??p�?�p�>�sl?�o���B�GD0=6��>�k?��?U���9��A>�	?�P�����կ���e?X�
@�x@k�^?�ߢ�VZ߿����琾شž0�.>Y@	>m�=NC�>	Rr�V��;���=�Y�=��>6>>2�I>��%>6 >	��=�,���#�����6����'�n��d�&!s�O3��k���r ��Y�8����'ͽ,�½ߧ�2C@���0�����>�B?�\�>���?7{+?Bަ<�C�:�zȾ�.��ﶾ�p>T]�>J?�sv?�N?|��>�ׅ�̒_��{�������u��	�.>���=���>��>�1�>�3���*>:�>f��>��>�$��:E��}g�=(65>d%�>y�?��>�mg=���=����֜�8�_��.龅�O��ި?���xp[��`���7��uƾ ��=B�"?�%�=AE���Wٿ�ڮ�7�D?���h��-�b��\>��<?$pZ?�	��v����Ϸ��z>_��I���/{ֽ�+(���������I>�p?�	>��{>r�(�� ?�
 U�������
>e�X?�;5Mz�����'(>���;�(�>���>c}ƽs-��3��f�t�{�N����<��1?�]?>uP�mԱ��
��bP��sAk>��$>�S����|='�m>�x��fkϽ��?����;�g�=w�>��?
�.>�ۄ=u͡>����*$L���>|�A>�Z(>��@?Y�#?x�=�%���t����6�ogs>�>�т>��>�K�!�=��>}�`>ʷ�`���P��Q>�Q�T> ����_��f��ь=�<�����=~ӑ=�����=��0=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>�1ܽcҠ�,����т��=���>�e?���f,��巾?���>ė��_��j�{���<�>N�?��?<�d�?��;yj�
b>h��?kd?�੽K����;�8��>�D? �0?;�=laN�v�5��,?���?*�?��i>ּ�?t�u?Y��>�}��E)/�5G��?$���==�m;=P˼><E+>�����>�����Ē��Ϲm�����~[>��<~(�>b���¾�J�=XUZ��!R��q�>ךJ>cCC>���>��?s��>��>Ӑg=մf����㧪�sL?�E�?J�	�i�/��<ǖ�=�a�RM?i�2?�o���ξ�v�>��[?w�?[S[?5a�>}r�����$���T��k�<q]B>�y�>��>[�}��}O>>WԾ�E����>��>��4�wؾ�ŀ�ϲ��jŝ>�=!?���>N�=g�(?�*?֫�>Έ�>*@�����$\��d�>�8?�oP?dKz?&�>������-��㠜���G��M?>ٳ�?�
?�}�>=щ�ⴑ��k�=}��Ŀ���T?rSF?<�x��?��?s�(?�?��>����U��|��$!(>��!?"�;�A�k7&�7��2|?]J?P��>V2�� ֽ��ռc��'m���?*\?E&?:���)a��þ���<� "��.T�Ey�;�C�t�>��>_g��k��= >��=m.m�~B6�ŵg<�c�=p�><��=
�6�M��C54?sҺ�0�����=5鄿E��ޏ>��>f�ҾYh?����w�����F'�����9A�?���?ꇞ?��Fc�5�A?e�k?��?�?ۏ���Q��^;�Ӣ-�k~C���E�_�a����=ױȼ]v����ԥ�ׄs�����,���[?T<�>���>�f�>��s>��>���%h#��5��2���=~�ߐ2�NF�S&L��!��S��KM������Tþ�����j�>�@c���>Kh?G�e>�Z>��> ��M>�>�H�>�>b�>>>�Ҩ=����O��KR?W���/�'�������P3B?�qd?1�>�i�5��������?���?_s�?�=v>�~h��,+�Qn?>�>b��Kq
?�Y:="B��=�<�U������2��v�.��>�D׽� :��M� nf�}j
?c/?R��G�̾�9׽E���D�o=�]�?P�(?�*���Q�&Vo��2W�YR�Ø��f�����{�$��p��ۏ�����Ƀ��'��4=�}*?�Q�?|����쾙e��t�k��"@�]�g>c�>_�>� �>]lI>��
�X61�-T]��(����[��> �{?�p�>m<?[M?��l?��f?�Ņ><��> !��t�>kd ����>��?��
?|n3?lHT?�e?�z�>-#>>���	�ë���N0?�s�>'?V�>�V�>,���3����\<�=����zE�/�9�]��:[��	��5`1>]a�>�W?{��e�8�p�����j>{�7?��>��>���3"��B��<Z��>��
?�>�>� ��{r��^��X�>���?��Lr=��)>\��=\5��JҺ]�=������=���Ă;���<��=V��=�q�,?����:F�;���<�b�>Y�?�ok>_�w>�J�����E�����=j�/>���>2��=������Њ��GHw�S�\>�>�?:��?���<%��=�$>�/��O�ľ��6��R� �Gs
?��"?��L?p�?[8?�K?��>a���|��ON��9򭾼K?:!,?��>���ܳʾ����3���?�[?�<a�c���;)��¾B�Խ��>�[/�i/~����]D��򅻥�����#��?�?_A�H�6��x������[��?�C?�!�>�X�>��>�)�b�g�g%�71;>���>3R?���>I�l?�7|?�G?���=��8��������9F�XeR>hI_?�W~?&��?��`?f��>`pb=�V�����\ ��(輻- �Ǎ�Vd�=�O>�q\>���>� �>��>=���&���\�r>z`�>h@?+"�>���>���=O߽P�G?���>>d�����M񤾎�����<��u?���?��+?��=���U F�V��~$�>�i�?"��?7*?��S�H��=�Uּ�ᶾ��q��0�>:չ>Q+�>��=�zF=�e>��>&��>��BY��m8���M�s�?-F?=��=� ƿڢq���p�hŗ�h�d<4��:e��o���Z��-�=�ʘ����ȩ�%�[�!���˂�����{���l�{����>�r�=��=P�=�q�<̗ȼ��<m�J=��<Lz=�Np��hl<�-9�ӻ@�������[<��I=%?�m;ɾ�x?�rJ?&+?TWG?��z>� &>E��F1�>J���ۜ?��;>��r����t�'�����쓾3�վX ԾVR]�ܙ��O
>pw?� >�]A>sx>���< �=zu=/^=NE��L��<��=�Ĕ=��=��=n>l>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>!g8>��	>S���0�J�^�P�\���S�x ?N�:�5dþ���>n#�=�z澉6ʾ���<a�1>�{=����\��=�zy�}s:=<_=D~�>a�A>��=Τ���/�=�c1=�'�=h�R>\�;�p,�aZ��$=���=gH]>C9)>5��>��?$}0?p0d?���>�qm�k�ξ����Ë>��=�.�>Ʌ=m�B> E�>z7?a�D?×K?Ͳ>�z�=k��>ۧ>�L,�A�l���3ᨾ]s�<���?x7�?�z�>�|<�%A��%��=��½��?@�0?�;?:�>ݪ�(�9�k�)��L$����<��<9��֒K���Ҽ��M����ڌ%>g��>@x�>�>+	i>��*>Cej>�s�>�8�=NK���r<^=ݽt1мH��=��X>`�_�=��=��@�����{�u=�'�:E��=%�3���u=��<�:>��>b��>�	�=l:�>}i�<rF���FT>v����|H���@>�v���`�Xy�XW���PF�4�6�`wy>J��>wŽ������>
�k>�>�R�?�*i?��&>
���w־�����DN��$��Y>��>�>4�U�8�?KX�}6H��hž`��>��>}��>��l>=
,�z?�x=�	��a5�&�>������=�<q�-A��X�^i��Ǻ��D?�C��)Y�=t(~?�I?���?Ў�>O��ؾ~0>uV���v=��m�p��O����?'?���>�׽D�]H̾����޷>�@I�6�O���=�0�J��9ͷ�^��>������оV$3��g�������B��Lr�s��>.�O?��?:b��W��+UO�����(���q?�|g?��>�J?�@?�%��>z�jr��w�=��n?���?E=�?�>��=p˫��D�>Bu?V��?Ү�?LXt?{e�U7�>;+�;,R7>�혽�+�=�>���=��>Hp?Q!?�<?����'�p2�Wc��H�Q�yaS=���=LM�>�n�>���>��=�J�=#��=M�>0H�>��>~�f>�P�>6�>�?���E��?�V=�U>�s=?��>h?�Q%��"��=B<�����)*��I�e�m�����<���=Q>���d+�>�¿�v�?��N>|ﾘ-?AΥ�_�!��~�<X�t>?�>��?�)�>L��>Y��>[f�>�@�=b^><]">�̾���=��}���(<���`���־��>�ο��Y�����<��+�l�k�ľ ��6N_�Dk��:�V�&:A=�X�?�Bp�UXs���-�t���A&?ˬ>�r9?g$��UL�<��=h� ?K��>E���s���c���׾�L�?��@<c>m�>\�W?�?f�1��3��uZ��u�Q(A�^e��`�s፿朁�ݗ
��	��	�_?��x?7yA?�V�<�:z>^��?��%�ҏ�)�>!/��';�D<=�,�>L)��.�`�)�Ӿ>�þ7��IF>�o?%�?0Y?iRV��q?��F=�LJ?6?6�?�?�wJ?QH⾺@�?y��=�'�>=�D>2��>,	?�{?h�>{_>�틻�ǡ<��w�5Ny�#���#����Y�=�8�=㣇�ӵ>��">7нH��t�&>��>Q�3���>�z>�F@�*%�<K��>�\?A��>8N�>�8?���c7��ݮ�s.?h9=�:�Tщ�����!+򾹤>�i?g�?�Y?�Vd>
|C���B���>9 �>�y)>�\>�>���l�B���=`]>��>S��=u�O�҅���8	��ے�s��<�">{��>�K|> 䍽(>S��(z�;qd>�Q��ú�4T���G���1�G~v��k�>-�K?�?�`�=~g�㾖��?f��)?�F<?KM?B�?E�=G�۾s�9���J�"E���>�L�<���"�������:�]�:��s>l�����JL>0��7?�(*P�Zoo����>@�.�+��=x�*�qE�&���u�>Jk$>,;ؾ�=��ϖ��r��h�]?�kX=����B��E��E,>v�e>�M�> ���ԣ4�����C�J�>�g�>�R>�8=!� ��iW��?/�i�>�0E?u=_?�k�?肾��r��
C��@��mw���ٽ�AC?��>��?X A>R�=)F��4����d���F�6#�>(��>E��h�G�`�������$�E�>M�?��>��?e�R?�?JO`?g�)?�]?�>����KḾ-B&?,��?P�=��Խ��T���8�7F�1 �>��)?%�B�>�?��?��&?��Q?��?��>Z� �<D@�d��>�X�>��W��a����_>ثJ?뛳>"=Y?Ճ?��=>��5��颾�ԩ�[�=�>^�2?6#?�?���>V��>�����=_`�>Z�c?�Ђ?kzo?
�=Q?��,>���>��=q��>�V�>��?[UO?��s?�J?���>7�<>i��kV��W$t��HZ�^ϑ:�6F<��d=.K�}�j���j��<e�|;PԢ�˿7��zݼb�6�!S��v�;2^�>t>�����0>�ľQ����@>eL���I��Y̊��s:��Ƿ=U��>m�?5��>SY#����= ��>�;�>#���1(?��?�?*�&;?�b��ھ=�K���>�B? ��=}�l�$}��b�u�aNh=��m?��^?]�W�_��Zc?"�_?�Ǿ�AX�Z�þ���I[��Z�Q?�
�>����+�>�DV?��|?�h�>f�=	Q?�f.���K�q���3w=�ҽ>���75S�<�e>��1?�y#?���>�E<>ߦ��|��\wþ��J?Δ?y��?���?f˻��e�����^�� n��$�^?D��>p���"?����kϾ3G��I���K%������媾k啾�l���b#��%��(`Խ�X�=�$?=r?�p?ߠ_?��Y�d�v�^�5���U�e{�I ��F� �D�׍C��dn��7�����
显��L=;WK�ظQ�l��?�}*?��&�kP�>�1���ᾂ�羯IZ>�Q��X�����=�I���g%��=�:�q2���[��6%?�(�>4v�>+8?B�}�σU�ILF��?�\Y��[E�>x��>��
>HP�>i�Q�w�=�������ھ~��s1Z��`�>0_?*�E?�oo?��ؽL�/�{~���;�ݖ����\�(�b>�.k=E'>�k�+���8��t;�/�k�u������&��NY�=X�5?�Q�>�}�>��?x?�������4*�[52���1��L�>��p?���>�͇>z�F����-�>�eQ?���>��>�c���-�s���X]����>�t�>G?�8!>pk��L�J��H��􆡿[I��<�Sn?����|���e�>.�5?��->�Q�=oh�=#�ｴ�3�C���#z���
=J��>�=�Ο>f���-u龫�^����$?J�?�[���])�H)�>+!?�m�>���>���?�G�>��ƾ��}�P�?m_?�L?Oz@?7�>�G/='l���-ֽ�&��C=z%�>�we>�W|=EU�=�*��0[��#�x7=�M�=
�ؼ��½�M�;�gؼ��X<=�=��2>f�޿��\��"�Vf=�ri��a.��@˾���<D�ľʯ">=�ǾS-Ѿ�I�������;KD;�l�g��N��\��Ԡ�?*��?�>6�����ȉ��|���!����>إľ�j0�Ar�7	��H�۾b��u��2#��Y�^6�/�:�*�'?M���ǿxG���޾��? �?5Wy?W���.#���9��*>\"�<����?�"��ϿU��a�]?*��>
��81��^o�>B+x>U
i>��>�m���Ej<L�?Ql.?r�?�#}�G0ʿ諻���<��?ʎ@}A?�(�����V=���>�	?��?>�S1��I������T�>i<�?���?�{M=�W��	��e?�}<��F���ݻ��=j;�=�D=j��ÔJ>vU�>+���SA��>ܽd�4><څ>.~"�����^����<��]>�ս�:��5Մ?){\��f���/��T��U>��T?+�>f:�=��,?Z7H�`}Ͽ�\��*a?�0�?���?#�(?>ۿ��ؚ>��ܾ��M?^D6?���>�d&��t�Ņ�=u6�h���|���&V�r��=T��>c�>˂,�����O��I��Y��=��{LͿ��&���.�S)-=�:߻�l7�t½TϽI��:Z땾1ya��:۽�=�='��=KO>�#�>s�->w K>!�b?"Or?��>�ȴ=�W�jA��^�侈s}=�)�������]�1Y%����������;K����<m�*.��y;?��	�="
I�t������})w���S�>+?�۷<�Й���]��DȽ�Y뾶y��#*��%�d{�.1���c��d�?�`<?ީ~���E�v@���m�ӽ#1N?_}�����_>G��<���=k;�>�n=� ��2?��2h��k.?��"?�¾	��&$3>+���%=w9-?�e�>�r<a��>�� ?qI�&���e1g>{�E>|��>p��>o�=����ɽ�?�L?�(�m��iy�>���
ԅ�[ۼ=��>x?$�U�W�GR]>NC�<Gm��&�8<��S���=��]?��e>c�=��Y侸����j�9E<TW?�s?/�>� �?�D?o�޽�"�<�k�)U&�j���0?�*x?���=�W	�\پ1�߾�1?��J?Ռ�=������M%�Q��[1�>�K?#Z#?ʹF=�1������z�
�H"?��?��i�J�����;��>h? �>��.�gB�>��C?7�ݽA&���Ŀ��5�Pŕ?��@AC@覯=��ʽGV$>�+?p)?�����N ���\�d��c��;�U5?�g�wm���z3��4�� J+?W��?-?(�5�����	>�P��	�?ɇ?ӵ���;�R�Z�d�~W��=�D�=����x�s���=��̵��2�7����q�H��>Z�@G�U<�>���²��̿�7�����i���C?��t>g��e���td���o�d,L���?�]Sf�VQ�>7�>���������{��o;�m��`�>���1�>F�S��%��	����{5<��>C��>���>:;���齾�Ù?b��P?ο���B���X?
h�?{m�?�t?.49<�v�c�{���P.G?��s?�Z?�\%��K]�Y�7�ZYn?ˬþ�e��$?�ΔJ�VD�>�<?hB�>�/(��F�;�|#>��?���=5�3�q���\J���tؾ�7�? |�?KY㾓`?ꝛ?�?0?����u��|p��S���8����P?(>V>�W��2�nN� ed��
?�0A?� b��)�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?Xݷ>Ԅ?���=��>hf�=g���X���\s>��=��&���?TL?T��>.��=i�8�\�/�6xE�S�Q���xoD�k��>X�b?ҴK?gDe>����~7�����+ֽw�'��� �� A�t�#���ݽ�9>Ѧ;>�>~�C��YѾrF9?�Z���ؿ䞨�kO��W�u?2��>��u>ү�@��b�f�9�?GI�>���l7��E����Z��j��?�V�?��>�ھ�L�d=��=#�l>�hr>ޣr=�L�+����>2�O?���`��t)?��P�>>�??�@��?�gd�YC	?'Y��X����~�����d5��_�=�c7?��C�y>��>���=�Xv�&���1�s���>�C�?(��?�>5jl?f	o��B���6=��>��j?�
?���\���D>��?������(,f?��
@s@v�^?����!dֿ�휿KM������r�=��=��2>&�ٽ�\�=8=1�7�IO�����=���>��d>?q>19O>�R;>|)>R��b�!��j�����}�C���:y�.�Z�*���Lv��|�k7������,���ýp���kQ��&&��_���=�^?�?B?#e?Cl?j\���(%>b�پ��	=��/�=òu><d2?��O?�-?�V�=��z���]�5R��h�̾�+��7��>^�>�7�>���>c�>��m;R+>>i(h>�3p>ȣ�=�c�=}F�<�wd=�4!>���>W0�>K�>e�#>���=8���覿��J��Cھ޴��Ba�?]�ݾx+@�	����m���¾���=�?W >������ҿb���7P?��������X���f=�b2?Z;?��>� ����,��->� 1���C��9�N2��3�������i>N%?�f>[_u>ҙ3�9W8�t�P�L���l�{>f=6?�궾jF9�ۨu���H�L?ݾ��M>�׾>�?�ae������#���i�n{=�^:?�w?�鲽ܻ���vu�N#��jR>�\>�$= ��=�UM>��d��2ǽ��G���.=t��=l�^>~?�7>+9�=b%�>?!��9/R�w6�>'�E>�)>��??:&?w�����~�|��A&���s>�:�>�cz>ˆ�=��X�;S�=���>�Y>�����@���{�KG<�5�U>2�V���_���w�1͆=V׏�;� >���=�����8���8=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ$@�>�h��r������=�}����=��>Y�6?����j��&���Jc4?Am?�8!�����;���4ށ��	�>qJ�?&��?����V4���"[�H��>�_�?hǇ?��X��v������z�>��G?�Ye?��>/ @�SbZ��(?]C�?%S�?��_>�ۋ?��k?��><w��K*������|������=N��>E��<��!�D�����𐿨�c�����>0x@=r�>I=�@z��|2d=��^�%_��A�v���>4�U>`,�>���>�/�>o��>���>bo�=��(���[�0<��TR?س�?]���7�ϣ��~ޘ=��n=7$?j)R?�ѽK���wS>t��?N'�?���?�$$? ��:T���Qɿ�þ����[l�x}!?�?�> �$���l=�4���/�Ƞ�=�8>�=ŽŢ	�W&G�.%�츜>Z�3?�"u>8�}=��.?� �>�8>��>S�B�u����>Q�>;�>iF?b��?��?܋�?��~�@Ǖ�`�3��(	>}�p?�?��n>4ɣ�ؒ��(�7�t+_��/>��T?�yn?B�ҽ��>㝗?��O?|5?��=������ʾ=�M��YF>!�!?����A�VF&��'��y?Ab?4��>葒��ֽ/(ؼ����"���?�<\?�Z&?Ω�E7a�7þ���<��$���i��P<{�F���>[�>�g��&��=^�>W4�=�Hm�\I6�I�l<�l�=���>o�=��7����T6?�dĽwꜾ�==xH��V�3�|��>��N>�7׾��a?XMʽ��n�����70������Ƅ?���?歩?� ������.O]?��?�A*?D�?�j�?��5�ľ��ܾ���f�7����=�d�>�$�9���
=��_���xd��˞��x�"G?���>ڕ?�?�̙>��>��A��G�0-��.���?!P��'�
�D�y�7�\_"�������T�>��<�Ծ�f��@��>	�:<�o?Qr�>�1%>�4�>�{�>�­��>�y>�kx>:�>x�>��n>��=�a�<M����KR?u����'����ײ��L3B?�qd?f1�>yi�+������i�?���?Bs�?�=v>�~h��,+�Bn?'>�>=��5q
?S:=T)�!:�< V����3�������>UF׽� :��M��mf�~j
?�/?K���̾�<׽�WV�7b��L�?�Y;?��:�^VS�J�r�yTK�blB�*��=��|�� ����u�h����l�G
x�O���T�=��+?(P�?s�E�x���%޾�{�I�)�z�{>u2?�c�>��>�4d>ҥ(�U�&��UR��)����\��>˫t?f�>��b?w�?�� ?n�??k�W>�E�>�S1����>ۺT=`lt>�nl>�bB?D?��I?��?>5,?�>�c�1O5���ؾ�)?��>WW?)z�>N?Ow����<��<���I�!��:h����;�R�=H7����@>��>9`?/{�p�8�����Ϟj>�W7?�5�>��>�������WS�<���><�
?h&�>Q �;�r��s��-�>���?t��R�=8*>��=�c��6��<L�=/tļ�"�=�ǀ�J�<��p<�>�=���=e�^�.{�����:r��;^��<��>[�?�p�>�\�>�j��й ����K��=O8Y>�kS>%�>qپ5���"����g��	y>�i�? l�?th=�F�=�h�=/٠�*f������󽾽�<�?�X#?>T?K��?O�=?�]#?w�>w'�}I���S��$���?�#,?ى�>
��ήʾ9��3���?�K?]1a����c,)�ً¾:^ս~�>�]/�g:~�����D�F+��	��
d�����?��?�_@�*�6����t����j��R�C?��>�J�>��>�)�`�g���w:;>�z�>�Q?�#�>T�O?Y<{?��[?`hT>C�8��1��Bә��r3���!>�@?%��?��?Ny?Rt�>n�>2�)�QྡR�����������W=�Z>H��>e(�>p�>��=Ƚ"R����>��^�=�b>��>���>��>�w>�F�<��G?��>b_�����社pă��=�W�u?���?̎+? f=�����E��@��vL�>)o�?���?41*?��S�Ǳ�=��ּ�޶���q��&�>�ع>�2�>h��=Q@F=�r>��>`��>r"�o_��p8��uM���?fF?���=�ƿ%�q�B�p�������b<�E��\de�1v���x[� A�=�����'�������[� ���Ӎ��	��ѥ����{���>�M�=�q�=���=_��<�rʼ��<F�K=l��<w�=P�p�Q�l<U9�#"̻�툽I�+��IU<L�G=�2 �̾�c}?baI?X�+?��C?q�z>�,>I�;�Z��>/-��^?��V>�'L��$���,:��姾�k��Kؾ�&׾�id�����>�C��G>8�3>��=��j<�=�Nq=pю=�=5��r=?�=)��=�'�=��=� >��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?��>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=v�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�t7>�>��R���1��G\�2hd�\���!?3i;��S̾���><7�=t+߾iƾ�Z/=g�6>�_Z=Pr�+�\�qЛ=}��88=wo=�|�>��D>$N�=���$&�=�D=���=!~P>����FB�Ի2�N7=m_�=]�a>��&>V��>��?�`0?�Yd?g5�>an�o*Ͼg5���>�>�G�=�W�>���=k?B>���>��7?n�D?��K?w��>�؉=��>��>�,���m�Qq�Yɧ��ܬ<_��?І?�и>�bS<RnA�|���e>�4'Ž�w?Q1?3h?�ޞ>Ϸ����S����:�S�.�ʧ
����=G�|�]���.><��`q�c}�:*�=㒽>�>@ّ>ԐY>θ�=S�=G�>B,&>\��ˉ��p���|��"�*Vx>�ޙ��a>��=�$��e�����H����N<�'=��J��Ё=�H>�+�>��=W��>�������>���HUq��q�<�N׾�5�N�V��n���aD�>�j�7L>��>��26��)}?��>�ė>?/�?$?�f>�Ii�<���|���Sb��8�"�8JM>��;>7�P�}QD���v�ti\�H�¾J*�>쥔>wh~>�+q>�� ��>�B��3 �~�$�m�
?�:�6몽x�����c�廛�`F���Mg��n��L G?_����>�@�?��Q??��>�����2:����n<k����K�½�-?�W?9��>A�ɾ�R2�l�˾�X��y#�>��G��%P������0�1� �b����.�>�n��4KѾ�3��j��* ��}]B���r�0�>��O?�ڮ?H�`�籁��NO�������\q?�sg?��>�?�_?�잽rQ��_�=q[n?�~�?���?n�>$��=�禽0�>UU?^��?+M�?r?P�ٸ�>G�U�a�>����&�=�� >�J�=y�=it?�U?��?�[��E�������h�U�EA�<7��=�5�>AG�>O�w>�q�=8��<���=u�a>�3�>L�>��U>頥>�`�>!@��i
�26?NA�>S.�>��K?[�>ԛ>���X5���@�"Wu��'罐�A��ڀ��=�
=%>Y��� �>��׿'�?V��=���E�>*��o����>%A�>�s����>��>#��>>�>p��>�?9>��$>�>�����H�=�,$�_0�n<�`zT�ں����>��ƾ$�a�m
�����k�b�ؾ{�R�S�E����DR�	~t����?N�A��l�7�(������=#?J��>�T?o�!����z�=^�?c��>;5��D���D��B�žf5�?�B @�;c>��>S�W?2�?L�1��3�vZ��u�\(A��e�/�`��፿���	�
�r���_?��x?+yA?qU�<^:z>X��?6�%�_ӏ��)�>�/�';��@<=�+�>*����`�I�Ӿͺþ 8��HF>d�o?*%�?aY?�SV������S�>��y?s�4?ج�?�� ?��!?��l�W?����m}>j�>΄3?z i?+$?��>�,?��=8�ѽOi����>DJ;5m�<�'d��IY=������]�e9��;�j=�>��o�b�7��*罇Q�=E�=��8<�U=�D�>T�]?q�>i��>��7?Y���#8�A����//?Ƭ8=E؂��q��U���b���>&�j?��?^IZ?%�c>�B�f
C��D>X�>м&>t�[>�C�>����E����=��>�l>���=��M�����ϲ	��8��o��<�>>ã?�׿>JM&���W>�Z����e��C3>��ܼ~EK�iۦ��$=���7���*����>�rS?��9?�Hr=����#��
s���$?��$?g&?P<�?Pr=k"���+'��!h�k|�OX�>?�n=���ې��ڣ��W�K��d_>X�>�UF�=���d>����)޾�Ln��J��8��S=Zn��CQ=r���־��}����=��>&>��rG!��+�����L�I?�d=b榾�T�����I>��>��>u�9�5r~��!@�A���}�=?�>��9>bƎ�٠��F�X^��>��S?K`Y?�1�?$���Ir��(Q��������ru�=B�?��>5J�>��>;H>�⾊r+��l�cM�|�>%�>lM.�X��֓���ھc��=_�>S.�>�U�+0?d�G?��>�l?H�7?�b?�Ke>:���־B&?晃?��=�Խz�T�F�8��"F�A�>�@)?�C�C��>oS?з?��&?��Q?á?kK>�� �Ԟ@�ox�>[�>jX��1��A6`>B�J?[��>8]Y?p��?ro<>�J5��������9�=C�>��2?U#?ߗ? �>��>&���ӎ=��>Dc?"�?`�p?��=�?k�/>���>}֐=�>f��>t�?��N?��r?z�I?I��>f<�<Mf�������s���L�{&�;3�c<��|=t0��G�u��(��U�<�F�;�b���kw�ڴּ��@��R��� �;He�>�t>�񕾲1>��ľ�N����@>�����K�������N:��p�=ӕ�>:?�Ǖ>{�#�`P�=�z�>.E�>=���.(?S�?�?��$;?�b���ھ�K�;�>>B?Mr�=X�l�xy����u�g=%�m?|�^?fuW�61��I~^?�u?�e���%�4����]��ԓ?oL�>�>=ϣ�>|�x?A�`?�R�>��^��+�������R��3qX���0={�>�N��J�X�D��>�..?�Z>�]�>��� ���<�r�]�!#�>�ә?g��?S�x?�*>��s�2'ƿ���������!Y?��>.����V?f������|����=���\������W�������1%��耾�^ֽ8��=-�?� r?�fp?��^?}C��Zb�a����O�>����cG�eC�fG���q�P��������S�2=ر{���@��\�?½&?�00����>��)�*�о54@>y&�����w�=�J���]>=@�h=�0f�Ep)�
ĭ�J ?ض>6B�>;?��[��$?��G0�^�6�Z�����6>���>ʕ>�.�>Q;��[{-�J���̾W����-˽�D�>af?=%O?0�r?��
��m0�����z�1�l0Z�a�*�C>�	">o��>�ZV�ŀ���s1�Tv?��x���r�����o��=A2?�?�>U�> �?���>���]���F���=����;槌>PQ?S��>S(m>F���X�(���>j�l?#��>K^�>|����^!��|��Eͽ���>�s�>4��>q�o>,��\��S�������&9�5��=[uh?ٍ���z`�ǅ>��Q?_��:
/E<�P�>4�w�J�!����7j(���>�R?�ب=�;>)vžl=��p{�p��y�(?�B?�5��?*���>� "?��>�>X�?��>;4þ:	���?xC_?� J?�!A?I��>��=�<��L8ʽ1�%�|7=�ׇ>��Y>�m=ގ�=��ןZ��B �Y�6=���=�s��{̾�U�;� ��D<���<�k5>�ٿv+O���޾7���P���O����1������) �9-��-1������� ��.����T�&N��̈��_����?p�?.7��.�q�yo��퀿T��\{�>
\n�
��C1�����e��ؒ�������!���I���`�fZ�Y�'?�����ǿ򰡿�:ܾ@! ?�A ?,�y?��H�"���8��� >RE�<�.��ԝ뾩�����ο�����^?���>��/��d��>�>T�X>�Hq>����螾a,�<��?4�-?/��>��r�$�ɿU���¤<���?.�@|A?��(���ԭV=���>��	?{�?>i[1�NN�-���L�>�6�?
��?��M=�W�|�	��re?�\<��F�v�ݻ���=\�=�H=��ŢJ>�\�>���!SA��(ܽ��4>��>:�"�4��T^����<�x]>�uս����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=h������O�"�b��5J;�0J�����6,�>�~�O������xH�G����{�=��R>�(">_�>oa%>�mV>#Z?�o?qL�>�$�>��i��hվ� ��B>G+[�� R�������U�[������H	�\���u��!v��\��+�:��w�;�V��ҍ����HDn�zKQ�:K2?zN.>�����QV�L=�<19Ⱦ����<^Ƚ�'����ľyw)�	;X��8�?�R@?�����H_���0�< �޽]=3?�IW�c��B	���p%>�⻉��<�T�>d�=����L2���:�/L0?܏?���}����,>�b���/=�}+?zv?�q]<�ܫ>�a%?��)��޽�\>�54>��>��>r�>2����R۽n?��S?���휾t�>������w��~i=�@>N�4��.\>��<�~���E�ԯ��2��<�$Y?Vَ>��&���s鷾;��u=�!y?�?�Ӵ>�s?�#I?�<=����^�o��{J<�E?J(l?rp�=g�Ϻ�����^��K�9?�i?�>�����龛��kE�?� u?�j%?#N�=Z���ϑ���2?�+�?�n�󀜿��>���ܾ��
?�\?n˰>�JA�&�����@?给�8̤��8��(�?��?$�@�@�❺�up��iI>�=�>ԁ?�H��9�&y���	���=��:?h��z��BnJ�t��bA?�s�?<�>n�ѽ� 1�|��=7���~R�?:�?����J�]<U����k��������<�٬=o��.#��(���7�ͼƾ��
�vV��R���X͆>�D@��꽔i�>��9��F��?Ͽ�D�ξ��o��?헪>��Ƚ�N��C�j���u�'�G��I� P��՝�>&>�Ι��璾I�{��;�㪼2e�>,�����>!�U�;��K���+�<^ӑ>���>i��>񷭽 ǽ�<��?J~��-�ͿRc�����KY?+��?{5�?�D?kZ<�\s��w�VS˻��F?m�r?�0Y?W"�T-Z�kb3�5�j?�_���U`�.�4�nHE�*U>�"3?:C�>Z�-� �|=�>ʊ�>�f>�#/�e�Ŀbٶ�N���g��?��?�o����>[��?Ns+?�i��7���[����*�
z+��<A?�2>x�����!�80=��ђ�ݼ
?�~0?�y��.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�b�>�S�?v'G>c~�>�E�<߆ľ��&�țw=U�=��M>��?�Cn?,��>�`?>]_Z=IPa�(�O�"*p�f��_8���|>�a?��n?���>�祽���i>�v�3o��<딽��w����,�P�_�!>���>	�H>�9�����V:?ҏ3�D$ҿ�ڠ��VP��g?E�>��&?���&��d?>@ |?O��>���`���!,j��=�Q�?1��? ��>������<ߡ���2�>�I�>".M��y�<<��~� >��P?V����r��|�B���>i^�?,@A��?�.`���?���]���:������)��> �9?(�]\>(g ?�K�="�u�Ԭ����r���>Vб?J��?2��>��i?Lm���?��h-=c5�>Mg?�:	?����k�G[W>�;?{D��9��V���e?�
@��@Ob?���ҿ>���W��tR־a$�=�)�=9��=�KO����=�> l<L����l>�Ӛ>Q�>���>U>�f2>��>����Q�+��X��V\���?�����+��}?�^ʿ�7}~�]��c���M��b�+r��潤�e��NC�.{̽^LA>�a?��>k�v?�zE?ܾ�=�	=�3��."-��Y\�dPp>2��>�d?��g?��(?!�=\����0K�ly�&�̾Xn��?�n<Ӻ�>�,�>C[?d��=5˵>��>��>5c> n��c3G=���=}�o>ط�>��>��?�QB>~e,>���94���"g���|�i�߽9��?�i��� K�����ֺ����q��=RH1?�W>钿F�п4����E?���+��J��>q0?��T?R�&>�v������[u>d0��[��(>����]���"��QU>0�?I�f>��t>$�3��^8�	�P�����B|>�:6?�涾�<9��u��H�#uݾ9:M>���>V/D��f�(�����hi�e�{=�v:?j�?경�ా��u�HM���mR>�\>�=�=�PM>�0d��5ǽ��G�#.=��=��^>�<?v%,>G��=cɣ>~	���O�̢�>�|B>�V,>�??(%?"��)��R���o-��6w>���>��>>�>2J�&�=���>0�a>���8Ѓ�����@�^�W>B*~���_�Lv��ry=Q9�� T�=]�=-� �W-=�uc'=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�� ?�nJ�8g���
���W���Y>���>�p$??�侇�h�%�]��QB?h��>�$�^
���u>4��q?}��?�F�?�t�������W6�>k+�?���?w��>z�:Z�?	?-jX?�w}?al�>!0�13N����>���?-��?t.u>�8�?��w?iK?[���^6�c%��n����Nܼ��v>��.>�k�=�Q��%UG��w}�Lj��w.�ނ,��=��<�?�>,^�.y�e�=.�Ž�n��G�<�H�>�y=��>=�M>�	�>��>^ѓ>���=�pe��S�n!��@F?��?Gz'��(�.��=C��;B���>W"�>��#�a���ިH>=X?t�?��`?���>��#��흿�*ڿ ����4��M�X�'?��)?;Y�=��>�
���V;���,>1�>S#]=����i߮�P�2����>��:?�&?�>=�/?�|?$�F>Y:�>�X{�)E��b�-�C��>���>��!?�y�?�!?���S�%�-��؟��T� ��=n?�?yS�>�&���"u���L���� ^?̏?��Z=Kl?'��?y�E?<g?��>�pݾ���̭� �>"�!?���1�A��J&�,��y?�K?��>�>��5 ֽּ����v���?�*\?�?&?����.a��þ#�<��#�l$\��, <��C���>Ɋ>�x�����=5�>�ư=Ym�L16�O�h<�O�=�>b)�=�$7�"���F�<?`�ƽx��|=d=9C��>qL�%3F>�T�=tC־iG?��5�G�����ĿI���H���3Z�?K��?�n�?�+����h���Y?B�`?2O?�?��є�����%2��)����&��o_>�C�>@Y=���8����ʿ;F��|�i��v;?T�\>{�?�?�P�>��r>�o��T�V�/:����Q�Yx�/񾜖E�n�R������]�E���?��)gþ����t�>�'K�՝�>�?��I>*X>_�>EY�<Xp>Q�>l#�>H[�>}�>�y>�#�>��>>�T/��KR?������'�w�辣���q3B?�pd?�/�>2i�����
���?d��?#s�?�=v>�}h��,+��m?�=�>2���p
?k:=H���E�<�T��Y��J*����*��>z<׽,:�`M��if��j
?�/?���;�̾�.׽����p=<J�?GL(?�*�?�Q� o��V�oS�<f�?�d������$�2�p��Ə�6�����ѩ'�v�(=�r*?��?�r���ů�%nl��(?��af>���>��>��>�J>nd	� �0���^��q(�����ջ�>?�z?��>��P?�5'?s�G?b�a?�>�Ϩ>�O���?2Mb=X&�>�r�>�4"?�K?��3?�?��?0}>�D�Y=�D侢30?�a�>Fl�>(F�>��?��5��l�<B�=^pp��b��V$���=��Y;�5��F����=üY>�X?��v�8�e����k>d�7?7��>f��>j��-����<�>�
?�G�> ��}r�c�gV�>���?	 ���=}�)>K��=3�����ҺY�=c����=�8���~;�Y<ق�=���=�[t�������:M��;}s�<��?�E?uS�>��2>����=Y޾�⾩$)>�G�²'>���=_0����{��]����U����>#o?e]�?�=J�N>��=X�������n,�"����9�>חG?6�c?�h�?�jG?Ls�>^η=�c)��k��"�����˶?�%,?近>���yʾ�娿��3��b?�/?}*a�ʟ�n	)�v¾�1Խ��>/��T~�����7D��u�!��`M��Ȏ�?�ʝ?�@�?�6�ݖ��Ș�cZ����C?��>��>��>H�)���g����Y;>Nt�>�Q?@f�>��W?׺~?�if?�� >�06����]W��/���ŷ>gL6?��?�4�?�a?�r�>C풼�d�.h�:���	���۴�?�N��^�=Q�\>�y>tq�>gZ9>_�y=y��~�E� c���y=e��<���>yn�>`�>t�>6@ҽ��G?$��>�]��'��?줾jŃ� 
=�+�u?�?��+?.R=C��!�E��G��XJ�>ho�?���?&4*?��S����=��ּ�ᶾR�q�d%�>�ڹ>2�>ȓ=|xF=~b>��>��>�)�!a��q8��PM�a�?�F?ת�=������o��В�W�y���>#�	�O	־1GY>𼵽��{���q�L����w��_�߾��Y��ᔾ����?T�Fe?G��=mA�Ո�
�	>*�@�bs���|�����=����	� ��=�q>)�+��YC��@=�[�H �<f8j��˾�N}?�}I?�+?=�C?�z>>	�8�.Q�>���� ?��T>[�L�LA���Z:��X������2xؾ0�־��c������>] G���>�?3>�l�=�j�<��=H�q=V�=��8��|=?��=¬�=��=j%�=��>��>�6w?W���	����4Q��[罖�:?�8�>�z�=��ƾS@?b�>>�2��×���b��-?���?�T�?h�?jti��d�>��-㎽{r�=븜�=2>���=s�2�[��>2�J>���K������v4�?��@��??�ዿ΢ϿKa/>7>x�>��R�dd1�@>\�k1c��	[���!?V2;�*C̾�>�=�r߾�ƾ�-=�o6>dTb=0f�:\��=�kz�e<==(l=��>��C>+��=vͰ�-�=�=H=%3�=�sO>˖��9�9��.�r�4=GU�=��b>��%>��>1�?Q_0?�Wd?�:�>n��Ͼ�=��F�>B�=�E�>��=ytB>��>��7?��D?M�K?���>ܷ�=��>��>�,�J�m��m�<̧��ڬ<S��?�Ά?ո>�0R<4�A�a��-e>��$Žw? R1?/j?��>�5�F������Np���H��	;��i<�e7�(wN>�ts=�_��7�ϐ=�*f>+��>/��>��->�s�<R�S=L��>K��=�|����=�`;�?#�\�>p�P>�l^�>	�=���
��=
c���D=�5}�Η=V��;u�<܅�<�@0>v��>r; ;-f?�3=���ο=�X�Ao�	=�\��#7a�4{�4#����P��'���>��n>񫴽̒��g(?�>$�y>�=�?�+�?���=Ԭ����
�՘����޾�-#���>��>o�����Z�C-b�F�����=�>箏>
t�>_^n>� ,�]?��hk=)�⾇	5����>���*��0��R�p�H����!���	i��T��aD?\��<u�=��}?�I?ؼ�?bh�>������پ��.>���}=�\�Q�o��Y���h?#�&?���>bB�kE�@z��3��D�>
᡾�V,�cY���LC��� <$q�� �>VV�ͬ��7�V"��K7��jn"�������>/>?�?zD��Út���H�3O@���>��,?�7?S�V>}l�>�P�>l�c<��׾����2�%=�2??�i�?� �?�%>H��=r>��0%�>��	?1�?�{�?�u?�|=����>)�8f >�O�����=��>]��=F�=<�
?�/?��
?����f���꾲��VdY��b=���=W��>@�>��m>a�=s+i=lţ=�[>3.�>���>�e>V��>�!�>(�|��<�_�?��>R�>O 9?�C>P��=쿅�2���G�������*�� ����=�|�=juL>�]���l�>��ʿjצ?ݻ=���l�>׮�|H�=O?�=�9A>�=��?Z�=�?>i��>}��>���= !p>���>�оF>94�f"���B�ZvQ��:Ҿ�y>����$�"
��S��M�+︾��׬h�߶����:�E��<*S�?�����j��)�r�??j��>I4?7b��޺����>��>˸�>W���*���ҍ�DB߾�=�?�?�@c>�$�>�W?��?�q1�1�2�XnZ�ɞu��5A��d���`��፿����!�
�z��Ի_?��x?�A?�E�<�<z>���?7�%�[���>s/�;��==��>����`��xӾ6�þ=��F>�o?S�?WZ?��U���r��՜>�j�?]K,??
e?�Q.?�Xt?�馾bZg?L!=��>��>{�)?xJ?��?Nn|>/=n!��N~t>��ٽ����K��=�R�Gz��l51=��=Bd��Lg�<B�߼�ğ���Ƚ��=
���<�+='��=A=�?�=���>��]?J�>g��>��7?r��u8��Ů��&/?�9=������MŢ�(��>��j?��?�bZ?lTd>��A�Y	C�/>�S�>1j&>=\>6a�>T{�	�E�<�=�M>�_>�ϥ=�`M�ǁ�&�	������#�<g->���> ^|>C��)�'>CZ���z�Rid>WR�}ƺ���S��G�n�1�.^v��s�>�K?�?>�=k�β���>f��!)?�S<?�TM?��?T�=��۾��9��J�0���>���<'��ҽ��� ����:�q��:�s>���!����h>
��{�q�n�ߧI�	^���`=q�]5=lI��Ծ� |���=��>과��"�� ��^���J?6!e=���oX�� ���^>f�>{Ͱ>�,�� ��|�@�������=gB�>n+>>�9:�x��,�G�5��i׈>7F?b7^?�N�?[���yt�9�D�<� �����9����?G�>��?f�5>�5�=��0���Xc���F��b�>���>���fH�����Hﾸ�!�V��>-?C�>H	?6YP?�?�7a?�#)?s(?h��>s�Ľ�C��ʅ&?���?�8�=%�Խ�[X�[8��9E�q/�>�(??�9˕>��?�	?��&?s�Q?��?�+	>�����A����>�/�>F2X����B�[>̱J?�S�>�?Y?��?��:>�j5�jġ��b��j[�=ӥ#>N4?w�"?�9?2e�>Do>��=���>7{?۲\?Ƥl?�\i?�<� ?��>�8�>s��=�}�	 ?ލ?m�R?���?�?�R<>;i�y�Y���,<���=�"˻�pT� @�=FLu>;~�>�O��"�=���=K�ϼ�=��~���n���Je=Xџ���<�V�>2�s>���0>r�ľV4��� A>����g��vŊ�Y�:��F�=5c�>2
?��>9+#�a�=⪼>�4�>a��,(?+�?s?�^;��b���ھ]�K�=�>p�A?qt�=��l��|����u�<<g=�m?��^?J�W����D�b?�nm?�{̾г#�1BľW���v�� ?D�?/���~Ҝ>[�P?uwc?
��>V"Z�g]��ē��d^�D������=s�>��_~�|ҍ=�GM?>�?զ�>��<�ɾ{Å���Ѿײ+?a�?�2�?Jޠ?�~\>�4}�}�ῸU��%G��^?�z�>$9��a�"?�����Ͼ����c��3⾏;�������T��h���e�$�c����Xֽ�\�=3?t�r?KWq?��_?C� ��.d�56^�Q���CV�������E��E�;�C��n��8�:��(��.1G=	�V�u�D��x�?�#?�4��c�>a�~�,Q�Tx�*a>ώ����R�d_�=~(�#
����=5a��M���ۓ�-4*?^r�>��>4�?*Kh��i_�4�6��fP���ɾc1�>�#�>�I�>�L�>�dG��{j��������e�Vx��}>G�d?�fK?�l?�x��3������#��)�䴝��nN>��>��>1�h����Q'�bB?��o�~��Ώ���k�=Sq2?�ނ>���>ܔ�?�d?�������$��UB1��M<�\�>,hg?+��>L��>.�Ž��!��;�>��w?�,�>i8>k`����-��z{���T�Q�>�X�>*?X�>�rf���O��������_�;���<I�m?�׎�.<��rb�>N�8?��=G
<�7>5���.�>T��`�E��K9?]�=� �>e6��C��XwX�ɪ��'$?�?gަ��>�Eج>�!?���>*�>��k?�Q�>������=\:�>�A`?$OM?L3K?h\�>:�c=(�%��Q�0���%=��R>��4>T��<K >�*G��,�x|P����=�=����MϽ5q=V�z�ע�=��=�3>�0ͿnB�����/���:�3���×����<�S���O�����k"K������D��
a&�dh[�^65����dt�u,�?��?�Ѿ�b���(��O���ָ��|�>��ž�;�����m�0��ѻ��G�Sg��I<��V��T����R|���7?�ʛ��տ����Kt@���?�R5?1c�?�����4��2��,�ҘL>i;�:�*����ߜƿ�����7?���>�`ξ	@J>%g�>��=#�6>�?⁩�#���6d�><�>���>�?U�{������Ϳ9�=���?�V@�}A?o�%�&��ĉi={ �>~�
?��;> �9�����A�����>���?_&�?YM=�
V��rڼ��c?��<�H�3����=3)�=�(=W����I>>�>�1��?�Qٽx�:>�>YE�����W�>�<h�]>�Qǽ�l��0Մ?{\�~f���/��T��U>��T?�*�>	:�=��,?R7H�^}Ͽ�\��*a?�0�?��?&�(?(ۿ��ؚ>��ܾy�M?oD6?���>�d&��t����=�6�Ȍ��m���&V����=M��>��>ׂ,������O�^J��v��=�=��3ÿ�]�\(2����<�=d5��EI\�i�<^�]�������2�}��=��>@�!>��>�bz>o�>��m?�o?��b>��\>��Ὕ�x�����F�=�����ӽ8��l<�M�޾���
T�a[����JV	����"�Wx>�ts�����p ��i]�XCk���4?�C�<b���T�x��=�S辪��۠!�i�"0��o��=j�⫩?!T?�z���X����qQҽ��F�K?�ح�:'����e�=rEA<����J�>.�(>;�9�W�_��a����-?I�)?� ޾.����>��d�M6�=�?�h�>���<���>��(?D7k�M�^�=Y�>&�>U!�>m��>�OV=s�����{$?�:?�!�݀��K�>�������t��<+��=���Ď�;�"L>��������ء=˙�K3�=B^?�r�>� �A��~ؾ=R��c�<bN`?b�?���>�K�?\]W?J�J�cY�/�w�k��"Q=�A?Q�v?]��=y�>�ˣ�[eо�EF?i|?�>��������O���fо�f?C/p? �K?��	>6S�3���|��ݢ9?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�(���d�?��?�����NX<����l������ȭ<�Y�=en��E ����v8�G�ƾ�
�D���ۻ�A �>�>@��a�>� :�m⿒GϿg���:ϾGo��?6��>��ɽ?��J�j�p�t��.G��H�E���|�>|>e>�1v�?`����}��z4����H(�>*\5�5��>4w�zaؾ�2e�t|�;^�>���>�QZ>��2�co����?w�Գȿ�Ǣ��� �n�b?���?�/�?"	?򧘼�Ξ�
�����=�y\?8w�?}?~�1$����#���j?�}����\�LH�<:R��4�=��!?�-?]@#���i>��=IT�>���=�J.�mÿ]ƿ�2�$�?���?T@�P1?�Ϧ?-�E?�3¾x՘����̟#��ȟ�d�]?�Z�>K�Ⱦf)C�
6�mO����?0�?�~̼R8ݾ]�_?*�a�N�p���-���ƽ�ۡ>��0��e\�!N�����Xe����@y����?N^�?i�?յ�� #�e6%?�>e����8Ǿ��<���>�(�>*N>dH_���u>����:�i	>���?�~�?Qj?���� ����U>	�}?���>g�?��<>G�>��";]�׾A��{q�<�E{=��>�|?�4?��?�M�;�aC��(3�`lG���L�ܾ��<�Ji�>�k?��\?{L�>�����-�����R
��_U�Y����a*V�@#m���>�>+>}-M=zg��������?Jp�7�ؿj��Ep'��54?;��>�?��r�t�����;_?Tz�>�6� ,���%���B�a��?�G�?9�?��׾GQ̼�>I�>�I�>��Խ����[����7>=�B?D��D��s�o�q�>���?�@�ծ?Xi��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?oQo���i�B>��?"������L��f?�
@u@a�^?*��ܿK�����Q��о��=e��hg>r����%�=��<6�߻1+g=���>�V�>��e>nSh>� >�U>�>�����(��x���/��+IJ��v'�����hf�����{�.�4��� ̨�M��9�����}�|~ƾ�5�'>��>��X?$�C?��n?��
?�����">���"�g�h���lL= �>��+?I�F?GH'?}��=����<\�Z���i����_���M�>L^>���>�T�>)��>�e<=2G>w�=>ջ�>W-'>�W����j<[�f=9A>��>D��>��>"}>Z�7>O�ǿV���c�g(��j����u�?�k���{c�囿�
V�ӚǾ���<��?�&>v���'w忾ï�V�P?XZ�ہ�4��m� <Ek1?^�m?�d�>Ğ��BQT�x~q=�}��P �h�1>�������;�'��Ц>�8?öf>�!u>g�3��S8�>�P�R����|>x$6?����u)9���u���H�xݾ��M>þ>{Y@��P����d�i�zoz=q|:?�s?�]���Ұ��u��/��1>R>"\>��=O��=�.M>�%c�ǽ��G���.=5j�=˘^>�?��0>�[�=�Ƞ>�'��a�<��w�>D=>�>�R<?�+?�vU�-NͽS_`�v� �d��>���>�w>/,�=�S����=i5�>��b>]�����E���1��]>\b��F�a�f]h��Z=R��B`�=��=�=��%@���&=�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>�x��Z�������u�2�#=A��>#9H?�V����O��	>��v
??�^�੤���ȿS|v����>L�?l��?��m�A���@�.��>���?�fY?ni>�g۾8\Z�t��>��@?�R?=�>�9�ΐ'�!�?&߶?��?�q�>�P�?�hm?ec�>�kf<�c�H�ȿ���2��=�>�=�>�b�=p���z���Lt��K��������ξ(J>��=��>�)���N�{��=�3��r���X y��[�>!>�W%�o�>�\�>���>P^D>�G�=���8�q�)1����N?��?3_���R�/����>*B'��`�>��?f�L=�./>��o?�+x?Hc?�I�>ŧ�90���Կ�����#;ґ<M�?�7?)0�=��=^��
���Xx>tA�>$>�[��k�y#��Ǩ>�[?��?Y�>y�+?�?�`;>�$�>*}h��ħ���;��d�>p�>Bw.?=�?'z	?Xؾ��q��P���`����>���>9�p?�M?_��>�ԙ�j:���Ln�,V(�kU�H��?�:�?h���HII?��?u|)?r�^?�>˜w��Z��$�n�>R"?�3���~A�u�$�6�?M.?gJ�>;����_Ƚ[��>�����ח?��]?B4(??��5ua���;���<g�U��mz��d:�@F���>S�>Y�l��d�=�{>[%�=�b�,;3��K�<���=$��>���=��4�%푽,=,?�G��ۃ���=y�r�2xD���>�IL>����^?`l=��{�����x���U�� �?���?Vk�?j��@�h��$=?�?L	?V"�>�J���}޾3���Pw�~x��w��>���>v�l���H���ՙ���F��&�Ž�Kݽ�Q�>�|�>j�?1�>SB?�v�>a�>�t���<��g�c�i��xd�m�߾��N�;�@�BҾ��r��vW=�b���A���2n>�
=���>��>�k>��=�<>~ԁ�L�>}�>�x>�x�>��>�Ă>�?�=d�$<ǧ���KR?����վ'�l��_����3B?�qd?[2�>�'i�5������?Ӆ�?s�? :v>5h��,+��n?�>�>���p
?�X:=?)�8K�<bV����V5������>�@׽  :�%M�Fmf��j
?t/?5��#�̾s6׽�IR���T�a��?�?N2���b��a�<@R�AV�\
>�Ս�b�Ӿ[��c��������n��j}�����5,�=�G4?��?"��U�w��m����E�]�J>�?��>��?���>H��K_Z���w�O9����j��>��c?�`�>�nF? �?��=?�UN?=�>l`�>�(��{*�>���<bӌ>���>	U	?^(9?�N0?m?7r.?�G|>����T��.�&�5?ύ�>�2�>���>��>@�{�V^��#�8$��<��?͎��O>��L��% �����]h�<Vp~>�?���u�6������h>��9?��>�0�> G��[���k�<�#�>$?���>Ϗ�6s�����9�>Ɓ?�5�C��<�;(>�r�=/����?��=0��N/�=*�5v/��D<��=Aa�=��<�R�;k�:��;&�<x�>�?
��>A�>TK�� � �"��Bn�=Y>�,S>,>�Cپ�}���'��%�g� Wy>Fv�?`z�?��f=f$�=>��=����HT��]��q���v�<��?O#?�UT?<��?��=?Wg#?=�>G,�AM���[��y����?D(-?��>Z��m�ҾKѩ�Ec0�E�?w�?k�_���
�W-�^���n ����>5�1�����⯿2�;��ӎ<�-��p}�0��?Sd�?qL޼�8�����藿Ϋ�AJ?���>�֫>���>-*���e����0>�� ?�YW?nD�>�4Q?��v?�F[?��a>/K5��v�����͛��|q*>�z>?���?vf�?�Eu?���>�>��,��۾����J�&� ��a9����m=w�[>N��>G�>���>���=E�ɽuP����1��V�=�f>��>!�>���>E'}>\��<��G?���>a��+��o���+����b<�J�u?I��?E�+?h=[i���E�T��(R�>�m�?m��?**?��S�Λ�=t�ּdӶ���q���>ǹ>�2�>�=mG=�7>��>Þ�>-)�o[�.b8�^JM�e�?<F?=ɻ=��ʿ��~� -e���� ���.�����k�P�˽�-G�T�=���2���,��J�P�����e���˸����e�\���>�E
==qUx=�"=��ջ�~<H��=r=?=����M3R�`�����D}������A�<�GM=��Sx˾to}?�8I?��+?t�C?N�y>�>}�2�1��>�ڂ�3B?�V>�Q��c���V;�hi���ڔ���ؾRb׾h�c�򷟾p�>>�G���>s�2>���=� �<q��=�q=B�=��B�ma="�= ��=ӈ�=}�=��> >�6w?X�������4Q��Z罥�:?�8�>d{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��:>�c>}�R� C/�zeP�Z�aZU��?4T;�_$ɾ���>�k�=nm��$¾�E=��=>_�m=k����\�$ʒ=��}�?�A=��_=UV�>��A>�=�t��A�=Ö<=f��=�dM>�Y̻�p9�"{*���/=E��=�Ib>�(>�C�>��?IX-?�d?���>u_e�QZ;��¾���>'��=�u�>��=u�;>y/�>9[8?�@E?ӒJ?i�>*Tw=-�>��>��+�K�l��J��x���_�<�1�?е�?)��>i�<��7�����;�����?{1??S��>�:��|��ܾ�f�d�o��K�ɔ����e;:>kNN�y��@�G>���>Q#�>���>��n>��>�@0>Xy�>o��>E�M>ˠ��tPP<B`��$e>�X�x>뻣=���ʽD�=��༻��<��=�vh=M>>��q<d�=�� >���>i�0>���>?�=�薾�$>r�.���U���=�;��X�1�o��x���8����X�>�q>���<�����>XX>��R>�E�?��?/�_>O���������䤀�?�1����<��;>��9���/���M�uKU�?�����>Jݔ>T�>�SO>E0��M>�'q��Ԁ���.���	?8���2c��
�k��o��|�������2o�
8>h�_?qp���U'>�?Ѿp?Mԅ?;c?�]��w��W�<�
�9&� .��\����)�X9?D�/?��>�]�P�`��&��s�Ͻ� �>�G�2�R�IS���,0��~Ǽ���#��>�p��|n۾�0��v���ޑ�N>>��x���>��M?���?W.=������N�0y���)��>�Nf?���>�O?�3?5G�����ŧ���u(=��g?8a�?[�?�>�Q>�㗻�x�>e�
?�Y�?��?2a?Lsn�X�>�_�=��>��9lAc<�1S>�>n�P>��?z�?���>�붽�� �ھ�M��b�g�`�P�>���>�;�>��A>vo6>f�,>�-����>T��>h�>iс>��>9ˑ>(^��W� ���%?k1>��>2#<?�u�>�A>qy���M�,�,�=����l�� �;�
��� �Z��1��=H�U=`��>�ǿFY�?Yj|=�����>��޾߀�pgq>���>`�8�9��>?�>��<X1�>���>c��=�΃>	�>�2ӾCs>���Bk!��0C��}R�T�Ѿp�z>�����7&��������bKI��f��kd�j�[1��"F=�.�<	F�?���U�k�W�)�='����?Ʉ�>K6?#֌��툽��>@��>�܍>?9������&͍�lR�I�? ��?�7c>	�>��W?��?��1��3��nZ���u��*A�e��`���������l�
�������_?��x?vA?�<.z>`��?:�%�#Տ��#�>[/�[#;�[b<==-�>�&����`�ܡӾ-�þ?��5F>�o?�%�?T?�SV�$����â���J?��?k�i?� ?��3?�����@.?�g�_z-?h��>i� ?(�?��4?�6�>� ?4�J���hq]�=�>�	�	�s��������=Z^=@������ >�.a=��%�D�>>,?�=��>��;��=2��=���=5��>�4^?���>��>=�;?��_-5�x����i%?wl=�ʃ�6����E���꾜�>xl?C�?�^U?__C>�=C��&F��b>��>BJ7>ǪZ>.ծ>���?����=x%>�/->y�n=��C�uu�޺�����1'=��/>4?�A�>����� >�$~��]-��g<>����J2Ͼ��53I��)�%j.�`��>��E?�C)?�W=���7`���Z��m?��-?ܳ_?w��?��>C��aQ��{Z�*�ǽP�>��=4���e���n��)�5���9=篩>V���ݾ�=�$���r�E��"z�� ��+>�~(��~��7^%�m���6���?O>3�Z>�`��_���m��@k���?_?���=􄃾���`H\�B�>�9�>��>>�.�<yW�]uB�O���\�B=r��>Q/�=CD=�����N�ho�F��>J�N?9�c?f6�?cQs�~he�D�H�In�����|��=�e	?�w�>Ny?��,>M5�=L�ȾEJ��a���=�<?�>��>�C$��5�̑���U�:���j>J�?;��=}�>�vC?��
?�g?��$?�0?���>���$�Ӿ��&?��?	(�<��<���a��0�h=�5��>��&?�Z�1�q>��?^�?r.?��T?2�?!�=ݱ�^�D��3>��>?�j�G��puf>U�;?ru�>M�i?1Tz?���=D�/��оD���/n>|M>�Y7?��?�+?	0�>qj�>wϡ�q=؅�> �b?H�?�ip?!D�=�?+�0>�y�>J��=��>t��> �?&P?��r?��I?�>v��<5���!����w��'���s;^�I<�l=}N�Tp��w$�S�<��)<����L�v���ϼѕC��x���T <hb�>�s>�啾d�0>��ľJ����@>1���U������Μ:��׷=gn�>��?6��>�:#����=6��>�K�>'���2(?-�??ʏ;g�b�d�ھ|K��/�>�
B?���=_�l�R~��|�u�Q�g=e�m?��^?d�W����@Ka?��^?�k�T?+��Rɾ�3e���Fr@?�X?��2�?F�>�Js?~�X?�+?�{A��4w�mɜ�Hb���5��iK=�a�>���Z��a�>��,?p��>є�>�Di=M�о��d��1����?�ڍ?T�?�ۉ?�� >�&l�a�ԿHs��}J���^?���>�=��1�"?���I�Ͼ�]������ ⾚������M���}��`�$�"ۃ���ֽj�=��?�s?O\q?-�_?(� �
d��-^����\V�����*�E��&E�U�C�S�n�KY��1������H=�k�{cA�'�?s�"?r�0����>�ɑ�����xؾ�W>5󬾓,���a=�]ýћ�<!J[=^�c�,i����-#?W/�> �>=�.?�Ub� D��B.�)4��kݾ��Z>	�>�>���>�QӼ�b+��]���&˾���/���4�>��n?��>?�Zr?���"�����.�D�<���.�>��<>��>ޚ�:���((���>��l�~p��w�� ���ft?�/>�>C��?>E6?z���� ��w|�|�K�D�����>�tg?V�>��R>��������O�>��l?k�>t��>�䌾� �I|��ѽhC�>7y�>���>0Lr>�/�x[��Ď������9����=�Xi?������Z�>߆>�Q?�3�;\�Y<3�>WM���R!�y�ﾨ�&�X[>B�?'T�=j�@>�þB�
�2{�����@)?��?c|���*���~>:"?>��>;L�>�5�?�8�>;�þ�c,�M�?�%_?�mJ?�2A?��>1�=���;�ɽ�@&��W*=���>h�\>�Lq=U��=���%[��@ �$�F=��=��μ$ø���<�8����Q<@��<�Y4>���K�Y��MȾ��D�\u��Љ'���о��=ZA�������#u�YP�4`��L��3=�&���轟���d�I�a��?Bv�?� 㾴;�,O��QS���!���>�ξ�~^��Z��I!�����8����f��y�(�uO@���c��n'?�T���ƿZ,��U�ھ~;?�?��?�B���!���8�d�.>4iG=%��g쾴0����Ϳ�痾� \?��>L�����нh�>c�Y>��>$��>
���퓾����:?�C0?&�>Tj���_˿����$�=[��?]X	@l}A?�(��쾙V=e��>�	?�?>K1��G������W�>+;�?Y��?�AM=q�W���	�'e?+�<%�F�L�ݻ��=7&�=�Y=����J>8U�>7s��FA��6ܽ��4>�؅>hq"����-�^�➾<@�]>��ս�?��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�}��=[��>c�>,������O��I��U��=8����ƿ�� �d�$����<n��S&��sI������I������'i��˽�q=���=5�V>�Ѕ>��H>�8^>�5Z?�j?FY�>P|>����琾I;�-<�t��?@#������v������Y��ܾ8��XO�ܺ��5Ⱦ�zN��i��$R�����2�g���he���7?�&=$j��J�4�^k�=�U��
Dq�O!o=㐻���/�2��9m��?"�>?%�~�\x/���ݾM�0�n �H�??W�P���A۾��<hU����=$�>"�>=f����-J�b�b�?v0?V]?J����\��]$*>�� �s�=�+?��?��Z<>*�>mM%?��*�>*�gb[>��3>+У>���>�H	>����D۽��?x�T?���(���ې>U`����z�p.a=�5>/65�m�鼞�[>[ے<1��U��S��;$�<f�[?��=P��X��#�����,{�:��h?N�?݉�>8 �?��?�Jн��ξe���� �؎Ƚ�<#?��p?���=ʻA>���ܱ���F?g+j?j�)U�A¾��5��0���?�w9?��J?�uh>�������z���P?x��?�9������L"���ž#C�>~�$? �?�Y�3\�=�R?�L������pʿ���Nأ?r@7� @j�I=oj�__�>�Z"?�9?Pj��6�%���-0��/�=�"?Ǆ��c����A=��6*��$?:��?g��>ہ
=�t'�L��=Rڕ��Z�?�? ����9g<����l��o���Ԡ<E��=M�_"�P����7���ƾŻ
�f���7���;��>�Y@&Y�]%�>;R8��6⿲RϿ����Rо
Iq��?��>��Ƚ������j�CLu���G���H������>V�>bD��<���	�{��s;�Zi��a��>.��~�>�S��ȵ�N���f<[C�>?��>���>�-���W��ē�?$"��8ο�e�����r�W?�>�?�?ޚ?*�2<Zvs���{��w�CG?��r?� Z?�"��+^�>X8�?�j?WY���S`���4��HE��U><3?09�>t�-�E�|=�%>��>'S>{/�x�Ŀ�۶�����/��?���?4p����>��?�p+?a��4���Z���*��y>��;A?�2>փ��:�!��*=�X���C�
?^{0?,���,�]�_?)�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?h�?׵�� #�e6%?�>c����8Ǿ��<���>�(�>*N>ZH_���u>����:�i	>���?�~�?Qj?���������U>	�}?4g�> ܄?x=>ō�>:�=�7���nf��9�<��p�vM>�?�\D?ny�>#�>�=�^L�Df��Z��JU�W�V�n9�>p[?@&:?ݻ�>�=\�j�?��h��O͝�%�A��+�s�N��>{���;n>݉>v9->�K�#��@�6?q�D�8.ؿ�՝�p9��dY_?$��>���>�.澀�⾥ �=Y[�?Y�>��+����z��j=���?6 �?6u?�1���:�z�=)��>�	�>�� >�Ϫ��X����,>V�J?�q��̛�(�p��Ӫ>v��?��	@Å�?/^���?�Q��㉿���/���&�2(>y�5?�a�e5R>���>P�>�+s�ͪ�Vt���>��?���?�I�>��g?V�q�
h;�֞5=���>�ic?k?���<���#M>4E	?6J�В�<�
�i?x�	@��@��a?jL���dֿ�FE�������%�= �=�2>�ڽ�f�=W�7=-�7������=� �>{e>aq>�O>ZU;>{�)>���!�!�Xk��!�����C��X{�4�Z�@���1v�Zv�a6�������V���Zý�q��Q�2&��_��̾=¡t?Z�
?�u?k"?���=��>~ �t�v>���=��>p�4?@o?�P?N�=�'���I�)d�A7��V����>�B=(8�>�}�>$�>�W�U>��G>~V�>v=x>��=�>�n�ԼJ>>��>���>��>'��=���=��[4���}E���Ѿ�D.�ǎ�?>i��,hN��=��#���ᨾ���=}%?D�>( ���WϿ6q��:A_?�|i�>�ک���">|�4?�A?��_>lА��o<��">�ν�"��vmo=16�H"O���?��>%{?6f>l�t>�3�k8���P��񰾟�{>6?������9��u���H�=[ݾO�M>8;>�C��|����%L�݆h��|=�O:?[�?ld�������t��M���R>��[>��=�6�=�M>�d���ƽ9�G��,=Bt�=	�^>n?8B+>Ż�=��>���&Q�\~�>��B>��+>PD@?3>%?!P�L���$&/�8�w>�1�>��>��>_�I��5�=��>��a>����K��Ѫ��v>���X>eJ{�y]�*gu�3�y=qҖ�?E�=�~�=ds ���=�h�%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾX��>oW?��Ϟ�P��=�l��>�3�>�Bc?=�6>�w�R�+�%?c�?�� �+���˿ݵo����>���?�@�?����%;��AB�a�m>ks�?�֌?�pc�o&���ح�.F�>��S?�'?.o�=`�<�u� =?�ս?_��?�GR>��?1j�?��>��D��d�gF���ۋ���S��M>��>�	j>�}��;�?��~�7󌿘�i��.�`F�>t�=�g�>b[���[P�G�=:샽琢��l�F��>j!�>ۭ�=���>��?)��>�>@=�u6=�U�?@��l�B?�ޗ?�)�"[-�?Q�=7}�=d�{�??�LA?M���ᾄ�=u�\?�5�?MGk?fO�>F��wi��|[��xʾI��=�=pk	?�?�Ԑ=t��=/���v��_G�=��>�Q̽�þ�;��	5=آ>��?�\�>p	>}�!?�!?2a>6�>�F��0���F��>#L�>��?��|?�|?Wͼ��0����o���h]�*3F>r�{?־?ŵ�>��a��-6�;����ͨ�Ƽ~?OLb?���}�?��?�l;?�=A?�S�>�S��Jھe�ǽ���>E�!?����A��?&���u?�G?��>�蒽� ֽbh׼���D\��I?'-\?N<&?W���-a�þ�]�<��!��4e�[ �;Ż@���>!|>^���Vִ=�>�Ȱ=��m��6�Lj<���=���>T��=�27�!b���;?��=�iS���;>�І���F�|��>pS�>����֔g?��<t���Z����ۚ������ʟ?�-�?w��?~{���v�MV?L ;?�Uc?���>xс�!^��jj¾��4������(�� >o[�>�i!>P]#�{�������c��G&����\�>Ax�>�
?�F?��s>�V�>'o~���9��-��X"�)h����;���@�y��K���c���_��TE������B��>�z�:�>�?�"w>u;D>.R�>p���(�>�$�>���>���>{��>6>�>�l�4�ýOMR?l���ƽ'�۰�1���(B?�^d?��>q�h�߂������?�{�?�n�?�v>r�h�C6+�eb?�]�>��� }
?J}:=���I�<TA������Y�����>/.׽$:�M��Kf�~
?�(?nh��Z�̾�$׽�4��31	=�e�?�� ?G�&��H�>ke���W�زV��;W���������&��Xs�wq��e�~���Hw��9R=2.?@D�?/&��"` ��Uɾ�r�:�"*`>o�>�>��>,�J>��	�-�5�Y�W�B�������>�{?Z>�b?k?>�Z?�y`?Y!�>��>��ž��	?�7L�+�>L��>!�Z?.R?�RO?��?��
?�P&>e�/�#� �7��;Z0?z�>T(�>���>��?��e��8g��K>��!=����q(��l�=�!<����4R�]T\=��*>Y?ј���8�X����k>�7?�>���>;���,����<��>��
?G�>R ��~r�ac��U�>ˢ�?��=*�)>���=}����ҺY�=!�����=1��jw;��w<@��=���=�us�^���'�:|k�;Bm�<0�?�t�>��>,Z>Q�E
�`�о�a>>E�@> Ǳ>��>�꯾�����i�t�o�>��?9��?Ѡ>4�=J֦���ھ�Sx�Z`4���ri=�)?��;?v#B?��?�`?��?�a\>�7�o�W�Z���ξڬ�>z!,?j��>W��Q�ʾ�񨿥�3�5�?�Z?P<a����;)��¾��Խ�>�[/��/~����GD�o������|����?���?�A���6��x辧���e\��h�C?�!�>Y�>��>5�)���g�%��1;>>��>�R?RB�>�Z?��{?,�a?�L>w--�o��������<�[�>�*-?r/�?�?h�f?���>�ƍ=�eE�y辄T��"�$;-н�.���9l=�M1>i��>�o�>�p�>�.<>GrT���Ži�g�(-�=-И>L��>�`�>UV�>zf>�N|�RH?��>�:��#I�J��������%�=^u?��?i�,?��F=#���F�XW �3�>p��?��?Wk)?%qH���=��������e�8�>ͅ�>[��>�=��}=V�>�W�>�[�>��Mf���;���3���?}�@?���=4Ŀ�-o�#Aw��P��U��<͠�X�l�m����a�(Op=��������{����P�����3���B�����R���]?�ފ=���=�+�=^�=���F�=�J=[�<�%=��N�H�w<���7������3�;C��;��=�����`ξ�R|?��J?7*?�D?�{>l>=�N�(�>[�g�Mz?)H>|i(�������0���D����վ�Ҿ�5i�it����>;FX��(>�;*>P��=K>�< ��=\��=��=lȅ;h�=��=�s�=��=��=>�>�6w?Z�������4Q�[罖�:?�8�>�{�=��ƾn@?��>>�2�������b��-?���?�T�?Y�?Qti��d�>+��;㎽�r�=�����=2> ��=p�2�x��>�J>���K��π���4�?��@��??�ዿ΢Ͽ1a/>f�6>;�>��R�ޘ1��E\��5d�b�Z�$m!?rC;��̾���>κ=#߾�1ƾ��/=%�6>��]=	����\����=z�TC:=�m=���>"D>�{�=���ׁ�=��J=J_�=̔O>V>q��9���,��N5=���=�uc>�>&>/�>�0?�2?��[?��>m�p���ƾ�&ľ���>~
>(��>��}=h�$>#(�>@L.?��C?U�F?���>�=���>��>��-�
�i�ε��1����t�<���?	4�?��>+K�=3�4��vN>�:@ڽ�^?R0?!� ?4��>��#߿z���I�C���i��n8�^ә�n`�<=�@<������`�,>�;�>���>_M�>t?g>T��=O�h>��>c">l])�BN ��-�=��52����>�~�����hA<�>=�H(<����W<�p<'A=�_��߽<c�>�d�>c��MR?���=~�|�b��=�>�Y�_�EW�<s��c�d�`'���w����`�D��nk>ᗵ>Sq��<��Rt?�;>c}>�?�?��t?M"[=���3�(����ؾ,��#�U>�>]�����S�:�l��N�	��h��>�}�>WΆ>�rQ>�	.�Ŭ6��(9��S�0���=�>f�M��<G�U�M�X��՝�!����Ou��]o��H[?}���4�W>v?@<?ֻ�?'��>����Ҿv^�=V�J�	ω=�?��w0J�%4ۼ�m;?�%?<s�>b���g;�e֫�~!ݽ��>~�U���N�>���c*#�K�(��I��`U�>h���ƾ�{7��d��R���3j.���b���>��M?�i�?��0�c��/I��%��~,�=��>Tni?�B�>ԟ?�t?Q�i�i��k���b=G)t?�n�?j��?6�'>@q�=;��;�>�d?�<�?���?�qt?�UJ���>�$;>q���\��=�>v�=1�=�M?�?A	?�R�������3w��Lp�y�<
�=ϑ�>^W�>b o>��=�Ix=vC�=�\Q>��>2&�>�}q>걟>R��>"&��O���?X=\>bڡ>@m:?:��>���<�Ҿ�y����4��f�R�5rk�j�M�U�`�2�Z��="
!>m.����?�¿���?�.��=!��q�>����S#�O�c>k��>�s���K�>�x>��>o�>�7�>m:�=�j}>�~>�2���z�=�����&�k���^N��P���{�>m��D_2�)�����x�������Bܾ�]T�Ve���H?�����=�?
H�� na��!$��lq�Am3?֊>��I?��r�N�H��O&>1�?k��>�f����G����ƾ��?���?Kd>n��>E�W?0?S2��&3�Z��u��A�jd�^�`�S���˗��*�
�=J½��_?��x?M�A?\�<r){>X��?�%�����A�>�/���:�ŅA=�n�>�/��A%]��Ӿ�þ[�VKE>�o?f��?�?(�T��,����(>�)�?��>�U�?�0?Ca^?��׾��T?��>e��>��=jd1?�#?^�?�:�>��>O�?=b)>8��E���Г=����P�м��=iI>=��=%�=�=��Gq<��ŽN�����V)=��>�z�=/��=]��><�]?_L�>���><�7?#��Hw8� Ǯ�F,/?�9=f������Ǣ����>#�j?���?�cZ?0bd>;�A�QC�(>�W�>zs&>2\>�d�>�{�x�E���=`M>\>�ȥ=�eM�{΁���	�㇑����<�&>���>��|>�B���W(>�,����y��/d>��Q�)T���T�'�G�2��-v����>��K?0�?���=�z龝ږ��Ef��)?J<?gWM?��?�=��۾�:�t�J�m���2�>}�<������K����:����:**t>�ʕ���xG>з�W�Ծ|��kQ���޾L�<v��Us=Q!��b־�Cu�� �=�> R��l���#������h�J?�-=7��������M���:Y>�>��>;p<���ʽ�B��
�����=l��>#c>O�A�"�.@A�0��E.�>�B?N_?��?�퀾�Gp�nk?�٫���w��@�ż~?kF�>�?�bJ>z�=�x��Ē�Vb��B��Q�>z$�>q����H�Xԗ����8I"��X�>9}?� >s?�gO?ZK?�Z`?[�)?��>$�>q7��� ���D&?�M�?8ن={?ͽ�S�T�8�]tE���>�(?�{C����>�T?��?�3'?S|Q?�?q�	>@. ���?��֔>�X�>�!X�՛��%n`>K�J?��>��Y?���?W�8>~>5����������t�=,�>V�1?��"?�C?�p�>���>"���� d=��>("a?���?��l?l�=E?¾)>9:�>��=��>U��>��?#HL?�u?|?J?P}�>�*%<����Cp����o��㻂W��{�/;톁=���q�ٹ���<�7;Q*����`��~�������9�4'<���>��x>����5�=Wñ�n/���aP>� �;hN6������0N��!}�DH>Ʒ?�>=���7�@�Ue�>C��>z����?�Ȝ>��?��=��n��t��G��y>l�C?��>pI�!���2���|�=/`�? %O?�̰�ީ��%�b?��]?�g��=���þ�b�b�龄�O?��
?(�G���>4�~?	�q?~��>�e�Y:n�G���Bb���j�C̶=�q�>�X���d�u>�>��7?O�>��b>�)�=�w۾�w��q���?e�?��?��?+*>�n��3�����؏�)_??�>V*��\-?����;D���x���|ھ��&��V������c/�����9Ͻ�A�=j�?��r?�Bp?�1_?IG ��c�0�[��@|��MV��Q�5=�i�C�ǷD���C�ȍo��B����/Ĕ�s	^=�	D�.�W\�?r$F?�9����;>:���3��gh�^��=a���U�=1R>�:}����=y�?>������<�eؾi��>U�>X�(?�=?�S��`�zz�a�u������݁>$ߛ>L�
?�5?�a�<Jm���̼��.�.t��eھ*9v>*vc?��K?�n?�p�*1�����c�!��/�+c����B>�p>~��>�W�A�� 9&��Y>���r����ju��I�	�u�~=(�2?^)�>	��>�O�?�?�z	�bm��Ihx�%�1�5a�<^2�>Fi?<�>�>l�Ͻ� ���>��l?|��>녠>���!��o{�|7ɽi��>�^�>���>�un>GE.�vE\�
H��dj���9���=��h?�Ƅ��5`����>u�Q?_C�:��H<��>�w���!������(��>�U?^�=2;>��žD3�l{�4B��'�(?:i?Ç��v�)��w>�"?ҍ�>�	�>��?�3�>5�þ-��9R)?9�]?j�H?��@?T$�>��"=w鳽S�̽�N%��-=_	�>�\>��e=���=~*��[�M�E�==yi�=�Ѽ������	<����`h<�i =�;3>� ����%�E�}��W�� m�Z��;�����#�ɼD�:�����Y�x��d!��k�ت����@�F��ĩc�7�?;�?�:ǽ�$�����1������>�¾{���u��o"��q���`�_Ǿ[;'���4�,G�u�?�M�'?@�����ǿ����<ܾ  ?�@ ?�y?`� �"�!�8��� >�]�<����R�뾪�����οA��� �^?���>q�-�����>���>ЩX>5Eq>���垾L-�<��?ч-?���>P�r�@�ɿ5�����<��?T�@��#?O�r�lѾ-Du>G*?��(?ʔ= �p�㻂=�ʶ���H�mQ�?��?�WN>�����V�?�1�>PDW� �ؽx�Z=�k���<	���Kb>&�>�����S�����L+�>�c�>��8��O��[<$��⻆�^>=�W�[����?��S���e�^j1���z�qu>�lV?m��>���=�2?j#:�Wο!)`�eU?��?��?d5*?"Tо��>fSھx�O?С9?��>�)�{�r���=r$P�N�<\ξU�O�l�=^m�>�K>�hH�{[�3�B��=< ]�=�4���ƿq�$�~��� =:z�p�\�bC轵é�$R�#b���o�e��:vg=�X�=��P>�C�>0�U>7�Y>tW?I�k?���>>W>�o������;S
��Ȃ�A��薋�a ��c���	�(߾W�	�n��Q���ɾ~;�C�=�oQ�gǏ���"��Uc��iE��3-?ʥ>��ʾ��L�e��;iɾG,��U�r�ؼ�� �ȾY31�PWl��s�?��??�˅���W��Z���ļ�鼽�V?~z�s�3����_�=N����0=��>E��=b��M2���Q�X:.?�&?c�¾Ԝ��!k$>�q�6�i=��(?a?�W=3α>�x?�4A�_B��YO>��:>�b�>�@�>Η>"��zЙ��\?u�Q?�L ��ڠ�T�y>�����z�:=1�>�� �����c>+�c<�1��D��`1�=� =�_U?v]�>�J)���Ƃ����5��[�=Dv?��?�>�l?�9?�W�ʄ��B�N�N���n=c+K?0Yi?p`�=G,3�#ξbZ����4?Uc?`�=>��]���X�0��_���?�rk?��?G���Bm��ؒ��Z�� �4?]�v?�r^��r�����Z�V�X>�>�Y�>!��>e�9��h�>�>?"#�^F��ع���X4�?>�@H��?��;<4)�\��=;>?_�>@�O��Cƾ8���W���o�q=O!�>�����bv�M��%I,��8?ޠ�?���>��������=�(����?@�?�ߨ���<7��Am�e����s�<_�=IT�*���_�j6���¾S�7'��Q�׼	�>�@wɽ��>��<�.��9п�S����; m��?"��>������{h��r��rI�8�G�����0��>��=���!⃾��|���8�Y�;�)�>�����(>K]0��(˾�p��0ˌ<�Ӱ>?�>�$X>?�
���z��\�?ށ��Cǿi��f�ӾKOF?þ~?��t?��?�@��xu��
�����`�-?��_?s�R?�ȟ��U�������j?`��5U`���4��GE��U>�"3?B�>��-��|=�>���>-g>�#/�"�Ŀ&ٶ����#��?S��?�o�t��>���?�s+?}i�/8��-]����*�i�,�}<A?>2>W�����!�M/=��В��
?�}0?Dy��-�O�X?0\��"t���4�^;=�]��>��#�O��~;��Nv���r�`��oA�&�?RB�?�h�?Qj�������?�ӭ>=�Ծ��ɾg�S<�V�>�H�>�6>�P�<��j>X,��CF�сT>�r�?���?@�?�ˍ��@����>�dg?��>��?���=D"�>
��=�̰�(�e�#>���=6i<���?�vM?O��>$5�=��8�&/��OF�8<R�����C�� �>��a?olL?)�b>�g��<3�s� �Lν��1�pS��@���-�s߽o5>�=>��>.�D��Ҿ��?Mp�9�ؿ j��p'��54?/��>�?����t����;_?Pz�>�6� ,���%���B�`��?�G�?=�?��׾�R̼�>;�>�I�>H�Խ����\�����7>2�B?Y��D��t�o�z�>���?
�@�ծ?hi�z	?���P���`~�z��!7�&��=��7?s1��z>���>!�=�nv�λ��M�s�d��>�B�?X{�?���>��l?��o��B���1=bL�>}�k?�s?�o��󾊲B>o�?������nK�  f?��
@cu@�^?-hֿ�����N��䗺����=L��=��2>l�ٽ`�=��7=��8�89��!��=7�>w�d>�q>.*O>Tb;>Ē)>���'�!��q��C�����C�������Z����Wv�zz��3������A��u4ý�y���Q�?2&�O@`�'�=��T?_R?�p?�0 ?m�u�FH >$������<kR"��2�=�C�>�f2?�L?sq*?��=�Ǟ��xd�~瀿���J�����>�tJ>��>�^�>�p�>�h>;��J>�>>���>�j�=�=�N�p�=*�L>?��>�D�>U+�>u�<>n�>Eʴ��/��,Qh�5dv���˽��?�L����J�6��������4��=�.?J�>�
���Cпr�����G?"i���w���+��u>�M0?v;W?z>�`�� mR�3>���T�k���=�� ��j��)��(O>�?X�f>��v>��3�HS8��.P�����T�|>�6?=궾��7��eu�?�H�m޾W�J>�[�>Y�E�?C�5𖿈c~�t�i�mr{=�::?�R?CL���ְ���u��ʝ��0R>�[>�$=
�=�M>Ga��Ž0H�N,=#�=�+^>2@?�>FF���h> ���w�Y]�>?t>s>c8?d�?%>u�K��(���B�ˁu>�"?U�5>�>=����KO>۔�>��d>�1X<���Ű����5���>PN���9u��X����=h3~<6R�=c���;g��A�B���=r t?*,��]l�����@I�pL<?'�>66�=pp��/ 0�7����뒾E\�?v@ ܌?�N��I;� %.?��{?s[ ���ٽL�?�O�>������>bj����<4���=�xv�?�?@-=����Qj���>??����h�>�x��Y�����=�u���#=���>�8H?�W��	�O�;>�yv
?�?}Z򾹨��.�ȿB|v�J��>��?���?`�m�UA��n@�Ɓ�>���?gY?�vi>fd۾�gZ�ۈ�>>�@?�R?��>L9�[�'���?#߶? ��?I>���?&�s?�]�>�w�yR/�0��ۑ��=Q[a;{[�>1>+���lF��ԓ�wf���j����a>eZ$=��>tA佹-���'�=����E����f�+��>vq>G�I>KU�>_� ?�Y�>F��>�<=����+뀾�����K?���?0���2n�DO�<���=�^��&?�I4?�j[�z�Ͼ�ը>غ\?h?�[?0d�>B��Q>��>迿2~��K��<@�K>4�>�H�>J%���FK>��Ծ�4D�jp�>З>�����?ھ-���U��^B�>�e!?���>uҮ=�� ?5�!?�m>��>�h?�D���&�@�<&�>J�>� ?Щ?�?���T�+�J���gb��|H^�A�W>G_x?Α?_5�>�D���A���v1�=���끽 C�?>&g?�H���?�7�?�;?��A?F�a>��'�Y�վ��i��~~>��!?캡��bb�BP@�"
�}>?CK?�?{���t��^ފ=5D$����q�>��{?�io?���8��J`�L��;`M�)�����<BN��B�<� l>����\�'�>���>��������'xN��(��tڇ>��>��{���*�t?,?��3����͠�=��r�>ED��n�>�L>/;���_?e%;�c�{�������kT��	�?�y�?��?���{h��9=?��?��?0b�>DJ��-R޾��,�u���w��n�޿>��>��k�σ�I�������샿W�ýL�ֽB~=?�O�=怙>y�?��m>�>�w�4���d
�����_���F�h
Y�	�����O��侾�V>P��v��D�F>w����}>�Y�>0�>>�>}(�>�/<�^�>��|>�T�>��>\�r>L�">v�=��a��5̽FI-?U�����ᾅ��#S��3j?�x{?%>)?�5.>�����pҾ/�>N�W?��?���>��}��xD���'?��?D˅��?Y"�=^>���f�ٽ�p��*���6>�ܶ> ̎�����I� z罏�#?�?s�=j�	��(�<�����=˅?F�&?�~+��WS���n���U�p�S��/�.�_�#���q$�y%p�@���䑄�\���-'�$(+=\�,?1|�?0�$�����Ͻj�F=��Tg>%��>7Ő>�ݻ>�I>�	��2�mw_�4g'�S����P�>�z?��>A�H?��;?��P?�$L?iΎ>��>cs����>���;��>=��>֔9?%�-?��/?�O?Ue+?��c>����5�����׾�P?d^?�? ?Ғ?a���J����E��� ~��z����$o�=��<ٽ�t�W�W=��S>(u?���	�9��8���{>�7?-��>���>�����(x���;�[�>�?�H}>�� ��Zo�]S��>�>�~?dt;��!=_�.>W �=͡������⵫=�^�����=�ލ��g���;��=I��=@��;���;q��+z&���<~~�>��?4s�>7�>�L��� �ԑ�P��=wRY>7�S>�>*Xپ����f'����g�c�y>`q�?�]�?��g=���=^)�=�_��q8����������|�<o�?.M#?HT?��?o�=?k#?�>�7�7X��y_��DԢ���?v!,?��>����ʾu񨿁�3��?�[?L<a����;)��¾R�Խ��>S[/��.~�s��mD�@܅����l}�� ��?п�?�A�0�6��x�ǿ��[����C?+"�>�X�>~�>:�)���g��%��2;>K��>�R?���>��>^�?i\�?6<ֽGcG����4�*o�e��=�3C?A��?���?MoE?�H>I�J>+�˾^��(O��="����qf�
A�=��&>Hn�>"�5?�t?5�=�����̳�=P�ž^��.�>ǜ�>���=�@>���=��>@�E?+�>���z��Y���N]����=U�r?{?d�J?�tt>�E&�8	]���~��>��?-�?69�>����=dw�=t>�K�#�Q�D>�[v>�ٙ>^�/�K�>�>�}�>U�>�Q���9���M��Q���?B�J?Dװ=U�ҿ'qd�lO��I��@�Ǽ����O�g�����0=D��l�=2_n�ŗ �b���^�[�g����̔�y���B����t��o?_v�=��>fg>� Լ)���D<���=�u����<�,���b;A�A��m_;���$ݾ��	"=�>�+�; U;/��?d��>'��>��W?,U>l�>C{>�_�>�x>�.�>�1r�;��oT�M��W=C��T���-�����ٕ���0��>>>�<F>�W�=`��=��=L��=�>=�~���\=��@�<5��=cl�=� �=�Z�=X��=$o>�6w?V���	����4Q��Z罙�:?�8�>P{�=��ƾi@?y�>>�2������vb��-?���?�T�?8�?8ti��d�>N���㎽rq�=)���	>2>^��=l�2�K��>��J>���K������4�?��@��??�ዿˢϿ6a/>;>���=�O���+�}���7Ir���O�1�?�C8� kʾDi>���=]־-�þ�l=�u>>fZ�=��"�tNP��=�w��7e�<���;�*�>q@k>e}�=������=٪X<�L�=RNK>��)<��;&]���`S=���=��R>�+,>��>r%	?c*2?�w?��>E�M�����CA���?T>^ơ=��>��=N>x2�>R�7?W�1?�x(?��>���=��>%|�>=�8���w�Έ��ar���U0=bw�?ԃ�?X�]>Ć�<lE��>���%����I��>"� ?��?/m�>�U�r���X&�ǚ.�Ή����:�!+=�mr��OU�����*l������=Vp�>^��>��>�Sy>��9>~�N>��>o�>j>�<r�=���߶�<?�����=妑�6�<�wżb���N&���+�����\ڍ;1Ć;o�]<���;��>ё?@=�݌>���=������q>��'�*�<�.��>s(^�^@B��p��,�����^g��3�=2E>
��=�Ď�3I?�j2>�]9>���?�)n?D�-=L�%����f���JW���U��a+_<d >mc*��4��WY�W&��¾���>}ێ>���>�l>��+��?�
�w=,��U5��>�������� ��,q��:��5�i�(�ĺ��D?OF���o�=�~?z�I?�?���>um��]�ؾ�R0>�@��0-=f�\q�Xn���?�'?ѐ�>L�q�D�%��2�����>=�8�l� �����LD����P�e>��g�u�ܾ��'�q���� ��պN�0 �d%�>�4?2��?���<��"���t�}[½��>��?�r�>���>�d�>y�ԑ��E8�U>��r?���?@d�?�š=7?>3�+����>��?N��?ࢌ?�d^?xA\�'�>��i��2C<����>ԭ�=��Լ�=zM?@q
?��>�@���	4�1����.�QI�<�7�=5��>��>]�+>5�>�%/=jV��p�/>؜�>��Y>r
&>r��>���>q�������?B��=���>w�1?�j>��e=�v��;i<Sȷ�T[.���	�sB���, ���<<��<��=��+��>�BĿ�!�?��c>�q�o?9����Y�e�z>�f>�Aнr�>y�P>`F|>F�>zӣ>�.#>��>��>�
	��1@>����*"�}BM�/]�v�ϾP�|>wƶ��'����yoS�r꽾(L	��o�pZy�`1����<`9�?KG�#�]�~T�*������>͆�>R�0?�L�����A�=<��>�Zp>�������ڊ��۾���?���?Dc>��>ױW?��?��1�.3�WgZ�7�u��A���d�ɩ`�>ԍ�����}�
����ջ_?��x?GmA?�ݑ<�4z>Ӛ�?��%��Ϗ��%�>/�j.;�w�;=��>�*����`�^�Ӿ��þ���ArF>:�o?��?�P?\BV�TCl�q�&>+�:?r�1?�*t?r�1?U�;?M���$?�x3>�I?�m?oL5?��.?a�
?�$2>��=Av���(=����ߘ��5Xҽ��ɽ����Y4=9�{=?"�9�<��=�f�<=���ݼB+;ܼ��{��<��8=��=���=��>��\?�>�c�>o7?���M�7������/?��;=�т�𮊾2]��H��5>�j?L�?CZ?Kc>�^C���B��>��>�'>�"\>5�>�p�ND���=��
>=B>?Q�=�>R�2w����	�<�����<�P>�e�>�|>⁛���>~���$�p�.�c>m�I�}�����P��F�?�2��A{�*��>wmN?�� ?�h�=md������d��=%?Z�6?��J?)A?�r=�U۾��6��CJ����HM�>��=:Z�=C�����]�5�4�;��`>a���[H���2>W���4�P���%e�&�52�<�O �U��<���"'ӾF�|����=hp>74����r$�������)S?���;�ʾ�픾K`��:'�>)q?>�Ց>�;��x���,G���Ѿ��=�$�>2��>gL=����-u>�e��`
�>`%?�-�?��?ǎ�񶀿�^�HB�:����I=w�0?\��>�n
?��>����K�O��2Yv��<�Ή�>	�>)�7�N�TS˾@��"C��>Q	?�p(�>�?W�a?l��>�Od?L�?v��>�>�HX�����;&?ŀ�?�i�=^�Խ��T��	9�
(F�d��>})?ӷB��ܗ>��?�?��&?VrQ?�?!�>m� ��@@�5��>�A�>`�W��b��f`>6�J?�³>eEY?�ǃ?��=>��5����������6�=�>��2?`,#?r�?Ŕ�>w��>�=��x�=��>a?�T�?��k?L�=)^�>�0>,��>g��=�N�>���>ړ?b@P?Ȯz?�<@?���><��O'���"��:��]1�}h2<z�<Ha�=��Ǽ��o��v� w�<�#�:[��5\�=5-���s��D��I;h$�>u�w>�r���*>s��Ө����H>lA��r��P8����A�(��=��o><?�>9=����=���>���>����'?�l?�8?�#e�f2`��־Y����>� E?ni�=mGj��ē�hKx��.==�p?U�_?�]W������b?��]?�Z��=��þ��b�G�龑�O?D�
?Y�G�8�>��~?��q?6��>��e�>'n�����Jb���j�d�=c�>�]�>�d��V�>��7?�f�>��b>��=}u۾j�w�kr���?I�?��?9��?*>q�n��/�%���D���]?��>�^����"?���Y�Ͼ㵋�����	��e��jT���}���a$�����q/׽�E�=|8?�$s?5q?��_?v� �pd�j ^�����SV�q�����E��E�[qC���n�D@�����\٘�6 I=�J@�+3���?�0?�@�`|�>��ľz��O���ڈ>����v��g>��н󦨻�E>�+P��6������0�>E=�>>4?^�6?��h�y[���Q��n!��B��G >
��>�'�>�_|>f"=�� !���ؾ]����1K��Yy>@U\?<I?�0l?���:22�0���E &��(¼�\����x>��3>��{>˗m���>;��3B��bw�v��ܓ���
�>�<�s*?5��>�:�>��?(�>���j����~��/���=e8�>vc?���>L�>�4�.� ����>hm?���>c�>e0���� ���z�f�ǽ�O�>�V�>9�>�Bm>��.�/�[�I⎿U����8��@�=��h?�����1_��2�>��Q?+�;]�K<-M�>�u��	"���'�*�>�_?w#�=rz:>�ažE���{��ꈾ)I'?��?񀓾^�)�r��>��?���>벨>h!�?�X�>��þ���	5?]?<�I?�g<?��>
>=�H��'�ս�(���-=^�>�;S>�Pc=��=UL�u�W�f���@=���=e�ټD��� Q�;:�ͼ�R<��=�6>�� RF��,��7���r��2�����'���������M����ݬ���Ⱦ}�d��t���)�f�=-��Ý���@"��?��Ǿe�`< ��7���gા(�>hz�!���t����&��@|�w����9�6���=��v�<�'?޺���ǿ����:ܾF! ?�A ?!�y?��c�"�ʒ8�d� >�I�<."��;�뾧�����ο������^?Z��>v�0��l��>S��>�X>fHq>P��=螾�)�<q�?�-?���>n�r���ɿp������<���?"�@�]&?�\`�=�"��_g>'1??�?io><(��p�%�q������>)�?~��?�E=Ad��\I�=ZB�?�e��b���Y�Ba�>�9�>y��<#5e����>���>j�Ǿ������i>�?�>ف>H��g�f���&�>�O�>uܴ��81�я�?�SX���b�?.��{~�!E>xU?"e�>��=��-?� H�MϿE�]�m�^?���?���?r(?����aM�>�ܾC�M?��6?��>Z�(�Ls�΅�=�a,��U;d�ھ��R����=�.�>sW>�:9�v	�&M>��V!��з=����pƿ��#��!�HC�<�#9U�[�C�l̥��jQ�=��Ύp�ŏ�WP_=���=XuO>��>�V>�U>f}X?G{j?���>�>M\��C���~ξ@������HV�|����������^�-Jݾ��������p$ʾ��=��1=�O�뵋�;^A��z��a6�O�?�M�=k���B�I��p�}�ɾ~���d�ͼ|�4�48��J��b-X�	�?k�4?�����W�� �I:������Q?I��~x���������=��=朮=l/�>�z�=�u�	4�v�D��.?�@<?	���쫌�2R>�˽Y�9>��=?�?�U=�P>��>�e�� ��Ȁ>I;A��>y��>�n�>]�¾�[R�^?5,S?R�½_}��[�>8�������=%i�=��P�J���k4=ē���7j����KH�S�==M?Uqq>ʵ ��]4�O���(�w=;6>pt?�q�>D�>��S?��:?:N�=kƾCS[�� ��]�=n�N?c@??�I�=�.V��޾^&˾C�&?�L�?��>uK��R꾳�N����m��>�j?�)$?���=*����m��Ek����0?��v?s^�xs�����L�V�g=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?P�;< �W��=�;?k\�> �O��>ƾ�z������2�q=�"�>���~ev����R,�f�8?ݠ�?���>������8)�=ᴖ��l�?�و?TP�������!Kn��+��˩E=��=�f���钼wN��6����{�#��x
�	�n>�2@�M����>��L���߿(пJs��ї��Ä�K�?a�>��֍��lb��v�'�>�?�B��!���ʗ>���=r��������D��!�N�Q$����>"нG�>;����ȕJ���<���=1�>�]X>`�:���Ծ?�?F��ؿ7^��뢟�0��?	{�?�O�?7��>��G�����z�:=T.?`�L?�D?�6R��@�������j?�_��mU`��4�sHE�U>�"3?�B�>X�-���|=
>���>5g>�#/�t�Ŀ|ٶ�/���I��?։�?�o�*��>n��?ps+?�i�8���[����*��c+��<A?�2>���D�!�/0=�+Ғ���
?4~0?�z�Q.�K�B?��\�f���j�l���T�<�>V�����O��?����d�~�`���,&�!i�?#_�?��?{�Q�T߾[A=?�L�>J,6��߾eм'�?�j�><��=Z��=��>p����1�x��<=��?8V�?�?���Dj����>���?���>`.�?�|�=���>P��=΁�����7�%>.K�=(�=�??��L?���>�c�=r�7�8/���E�{JQ��%���C���>&�a?˩L?Lb>pe��7k-�`� �<HϽ�0�r �LyA�ئ3����ߣ4>0�=>U>
�D��@Ҿ��?Op�9�ؿ j��p'��54?.��>�?����t�����;_?Tz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>;�>�I�><�Խ����\�����7>2�B?P��D��v�o�r�>���?
�@�ծ?mi��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?jQo���i�B>��?"������L��f?�
@u@a�^?*�gֿx�
J��������=t�=�2>k�ٽ�u�= �7=b_9��Ŕ�'��= �>n�d>�q>� O>pe;>~�)>����!�
q��������C�e����Z�����Rv�u��&���������"ý%z���P��2&��H`� ��=��U?uR?�p?B� ?$Ox�6w>ӻ���^=qU#�%r�=fI�>�`2?t�L?�*? `�=������d�Y��P?��Z͇����>�vI>0y�>jB�>��>"�t9K�I>IA?>}`�>�� >�e(=c��
=u�N>5L�>M��>�h�>;>��>�ִ��$����i�d�y�&3ѽ��? ����HJ�-3��pY��mw��]�=B:.?�>���4�Ͽ�8���PH?%��.����1���>�2?�V?]{>�V��BMa���>����g��>71��$�l��a)��3S>K�?c-g>7u>n3�LA8�j�P��쯾�|>�%6?�|���U8�6�u���H�L�ݾYOM>e�>V�6��7�"�r�~�P�i�{�}=Ɩ:?Jt?쨵�1��l�u�3���}�R>AH]>�=ʫ=��L>�,h��ǽ�F���0=��=A#^>�F?se���2>:��>�j?�h<s5>�窾�I=rdK?.\K?�Ǚ>iM>�	��󧾕�?��>�h�~��<�����s�=m�.?�E�>d^�ï��ڣ��,���?yV>��=�֖���|�q>��=�E=���<f���Nƽ��q�Ł\?�
��iw��J�H~�=#N?��>���=��r���C��'��}�ʾ z�?s�@��?y�1���}��uE?�ڢ?����H���ަ>��?3�U�������?q��<z����}�=��?�8�?�~�M��)�d�a�k>2G�>�
!��h�>8���K��� ����u��g%=I��>�:H?����R���=��s
?P ?M������ȿ�Lv����>1��?��?S�m�P>���#@�,_�> ��?gyY?nqi>�q۾�[[�X�>�@?�R?`>�>��v}(���?U�?@��?�G>8+�?�u?���>�A����2�����苿�|�=��<��>�u>�¾��E��j��t���>�j����إd>bd=.�>�彻P�����=�ڑ��X��;�}���>�dn>��Y>�Z�>��>�/�>B��>�5$=Ȫ��E������K?T��?���N2n��P�<���=ݮ^�4'?�I4?�7[�@�ϾҨ>��\?+?�[?Fe�>���6>��a翿�}��O<��K>�3�>E�>-&��:GK>X�Ծ�2D�Ls�>1З>����
@ھj0���ࣻ�D�>zf!?3��>�ͮ=�A ?S�"?x;m>���>.�E�kz��'�F�}��>���>�W?��?��?�����\3��y���$����[�ɥI>��x?�?P��>C���~C�����=�8�X1���ā?P^f?����?m�?o�>?$[@?uff>��=ؾ�ı�F�>�O&?nK����&�Tk���Q���?K�?P�?�t�=� ����ܽ�1����m>?�ˀ?�?�%�sb� k���*�<j}*=C�=7)=%(�@�&>�G8>�,V���s=P��>w��=�s����[�L�1ɳ�(?_ӈ>+�������+?5Ҫ;�=u�f}�=.�s��-@��i�>S�S>�+�� �_?�C���|��y��.,��XwK�Sw�?;
�?�4�?-��jg��=?t�?(?hs�>��a߾�=�CT}��(|�v7�0->Ĺ�>x�A������ �����~�����ҽ�[0?�۽>F?$U?M�b>;/�>T"�ßھ����;�sHf�p0�B�/�j���q$��Y��<]�0>$x龬[��_<>�����>���>��%>$E4>��>�;�a^>���=���>2��>f>(>�>�=��ܽ���??�gQ��6׾��.�����W?|�=?�`2?O�����
L"�2�>�uy?���?��?Q
���iF��9J?�P�>�N#���?w��=�#>Eet>	������6�>��>8b�>:�%�eNf��'~�3���V?��?� ;���˾��=�圾�Y`=�a�?��)?��+�NV�Eu��jV�BL���̼�}I�����"�m����V��� ��� M*�5w=m %?��?l��ع�������m���B��_>��>7�>+��>ӕc>����0���V�v�$��f���Q�>s?4|�>��I?��;?H4P?:PL?,��>L�>�ܮ�0��>�<,��>>E�>�c8?e-?��/?ؖ?x�*?[Re>5���Ю׾U�?m�?��?��?�l?�酾r�Ƚ�̛���k�[�y�u�}��J�=�һ<��׽��|���P=@�T> �?�3 ��86�����Od>�7?y��>GG�>ދ��E����<��>�R	?�z�>	�����t�{	�9T�>�?�f%���=� 1>D	�=�U��p�;���=����pW�=�m����{�V�;�2�=F�=Ia:<��D�e�Ż���<�8�<[~ ?��#?�6�>ڑ�>Y����x��tx����=���>��l>`�>�y㾳9���p����]���t>܍�?�A�?�M=���=+�>�����m������������<<��>�?A�I?�=�?K�>?Ф$?�K>��������k���[����?Z ,?��>�����ʾT憎r�3���?�U?�7a����3)�<�¾��Խ
�>�Y/��%~�m��zD��\�����
������??XA�>�6�{�5���+V����C?��>yW�>��>ȿ)���g��!�*;>Q��>�
R?UR�>i/�>^�?��U?�Y��
�Z�A�������
K
>#7y>(�}?���?�_T?)?7�>)�>ӵo�OY �V��LG����Խ��ƾ����ވ>O��>@�>�ۥ>�:���-��,��7���=�d�=;hm>�8�>G��>*V>t]}�tHF?��?XqY��I �m�ʾ����k>�l?�m�?�MB?xH��l�5���b�c��#��>�E�?y��?�3?>�A�W <�4>b�6�sF�ݱ->�a>W'n>�E#��L!>��2>*��>@��>ډ.�J1��N�����?��g?5,�<�Aſ�o��gu�����l��[F����`��ћ��c�)0�=$���i��(���]�?򟾨1�����	��e�v��R?���=�i�=��=t`<��ϼ, `<Jo=IHw<��=2�|�n�i< �L�;��`�k/�;�Ǎ;��=�!�0vҾ3�?��>]D?C�W?�*|>���>ӑ>p-�>�!'>bD!>��#�갥�֯����<N����^�*^���\�;Hоul����h��zM���=�0>��<s��=)y&>Y?���I=�s=g��=���=�5�<W�����o=�J�=��5��6w?W�������4Q��Z罣�:?�8�>\{�=��ƾo@?x�>>�2������xb��-?���?�T�?=�??ti��d�>P���㎽�q�==����=2>k��=y�2�R��>��J>���K��>����4�?��@��??�ዿ΢Ͽ:a/>G�:>�e�=�R���.��
T�aYW��!U�S�?6�:��3ɾV��>=��=�ھ�]Ⱦ��=��>>;�=����{[�

�=~Ou��T?= �Y=s��>��F>��=1<��j��=�gH=�=��L>9�7��h+��C*=�=��[>�!>���>��?�L0?�Fd?��>��m��Ͼ�a��-G�>%�=�C�>���=�NB>qR�>q�7?C�D?u�K?�G�>���=���>D�>��,��m��S�𙧾�ư<A~�?E��?��>umQ<>\A�Ι�fd>���Ž	k?�_1?�i?��>�U����8Y&���.�F����<5��+=�mr��QU�E���Lm�6�㽤�=�p�>���>��>;Ty>�9>��N>��>��>T6�<{p�=L⌻���<� �����=������<�vż0���\u&�&�+�䏦�V�;��;��]<Ѡ�;�u�=���>�>���>N�=���Ҩ2>�l��hJ�?"�=W%���1B�T^d���}��J-�t�8��;@>� ^>��n�r���֛?�V>��B>�U�?��s?6�>��xlؾ������c�ڌR�N��=��>�E=���:���`��L���ξ���>�ߎ>�	�>3�l>�
,��"?�C�w=��^5���>�u��Ԥ�j)��7q��=��(�Ii��Tպ#�D?�E�����=�#~?�I?�ޏ?g��>�6���ؾ�@0>[F��� =_	�'5q��h���?2'?���>���D�WϾ�����J�>f}G�0�P�0�����/���P�ve���{�>�Q��G�оwX3����m���W�A�Mk�J:�>��N?Bѯ?�^��+���O�@��h!��<�?�e?���>"?P?���뾧����=�n?���?�~�?F�>2��=b\0=B�>Z�>K�?� �?�?g?Я�-	�>�N<� �=/��F�=M�	>�\�=�
+=�m�>(�	?��
?������ �'f�c�f�m?�ÙY=��>ى�>K!U>Z��=�>U�>�)�>���>��t>4�w>Dp�>�v>����_,���&?���=���>��1?g�>�3H=�����|�<�2�7�9�o�)�L=�����y$�<�k��[9=��ռ>�>��ƿ�x�?��T>f����?�x���u+��S>��W>�3�ٝ�>őH><�|>\2�>���>��>�>��'>�2Ӿ�g>=��[j!��.C���R��Ѿ��z>���`.&����\%���
I�*Y���o�k�i��#��95=�A��<�A�?������k���)�����_�?]��>� 6? 􌾠����6>ߝ�>�Ǎ>�,�������͍��\ᾆ�?���?<c>��>�W?��?I�1��3��uZ���u�(A��e�&�`�o፿�����
����.�_?�x?�xA?�O�<�9z>:��?��%�lӏ��)�>�/��&;�r><=+�>*��S�`�R�Ӿa�þ<8� HF>H�o?1%�?|Y?ETV��Ln�m70>V8?�2/?X�s?�C0?J�:?.���%?�y3>2s?C	?T�2?2s.?l�
?z�)>\�=p�����==��Ƌ�ˎѽHXϽ��/�,=Eu�=d�;	�D<��=���<,۶�͸ۼ��P��������<c<=<k�=0��=<7�>��h?��>)�>� ?��ܽM�ć����A?t�>	璾����2�о�B ��!>��K?�H�?)a?s�o><*Z��5𽁫�=�>
Z�>�e8>Wv�>���HJ��E(<X�=� @>�>��0��؂��������h&=�o>���>:ׂ>��{�c[ >�x���[��w>�<�����e�6���G��&6�d��9�>`�O?� ?F1�=���r}��3�c�[�*?ވ=?GtI?ɗr?�|=�ԾV^=�6B������>��<v@	�̤�J��	2��h�<N�>꒢�w���67b>���k޾��n�J�n�羥M=|�$"V=t��վr���=[
>����� �7���Ϊ��/J?��i=�s���IU��~��|�>�Ø>��>��:��nv�	|@������=�=���>h�:>4ș���rG��.�aE�>�?E?.a_?^l�?�*����r�s�B������w��=�ʼ�?�X�>ph?PwB>�v�=����A� �d���F���>Ԍ�>X����G��2���/��@�$��z�>T0?Y>��?��R?��
?�`?k*?�8?��>����ܸ�d6&?��?
)x=Z�½�um���9���6��?��-?hT�	Ą>1?�^?8`$?�oR?�?_��=j����;��{�>T��>4�Z��p����[>rL?���>�jX?�Q�?R�\>x6�/[���1��`Y=f�>;�0? ?�??�e�>T��>ٟ��w�={��>*�b?n;�?e�o?���=i�?�M2>w��>���=�>�)�>`?.JO?N�s?��J?T�>�̊<��Ht���Iv�HVM�?��;��E<t�y=����Xs�x��y.�<�+�;����x���}���E����o�;`��>Ixn>K���R>>�nž�z��LB>>�8��U����Q��d�>��R�=�ڂ>*�?��>)� �~=P�>��>�$���&?9�?R�?z�;�b�@eվa�@��R�>��??&h�=ugj�//��֯v�{�p=3m?V,^?}\����Z�b?�2^?���U�<���þS9c����S�O?a?SvD�bH�>p8?r?�u�>�"h�	bn��)"b��j��в=���>�1��hd��G�>�7?BN�>�3b>�!�=�Dܾ��w�ɠ��?���?C�?��?y*>x�n�<࿫'����� �\?��>fa����?�}���A;p���Xc��B�⾪���bѬ�UZ���q�.�C��EH��6A�=�+?b�v?=s?�ZW?���Bce��/^��~��VP����DQ���@���=���7���a�~��Xx�Q��Ak�=\ ��3�x��?�"?q�v��j�>siƾ��i�޾��<�����Ya�Tb2=��=^)>2�=�V������$�
?��>_{�>�@7?8�Z�J�֏T�f�6��� ��K���I>���>��?�ɀ>昴�HY����ƾ�$z�Ut���Pv>{]c?ڣK?��n?ȝ�01�ׄ����!���0�{���"�B>,>4�>f�V��E�&�!a>�V�r����v��d�	�,~=C�2?��>f��>0H�?�?h	��f��wx��1��ǁ<h�>�
i?�R�>5�>�ϽV� ����>q�m?$��>�7�>Z�����!��gb��⟽��>)s�>E�?�/�>�vнC�^��̓�������4�W��=ie?[퐾���#�>��R?��<4iI��W>� ��
��+޾2@G��;�=r�?�۫=)6:>�&����~���`l��hM)?�I?I���3$+�Ĥ>�#?���>�[�>`:�?��>����Zwѻ�>?F(]?��I?tyB?P��>��=�Ĵ���ʽ�$�f�5=/��>ҌZ>Y�=U��=���q�a�O��S�Y=ur�=���� ׾�ɚ�;�BҼ�
�<�=-m2>p�ۿz�G�=�˾��������������X��5��G/��P�����r���	���B�lOZ���a�)��H�^��2�?`��?ͤ���"������#�������>{e��Fu����i������L	��9��3AG�&�c�8^�O�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��5�"���8�� >vC�< -����뾭����οA�����^?���>��/��o��>ܥ�>�X>�Hq>����螾�1�<��?6�-?��>Ŏr�0�ɿb���V¤<���?0�@1A?ͧ�E����\8�ts�>U�?��B>ѭ˽�<��2��B��>�H�?]��?2/��/_��O�^s?_��=hP�������>�L�=�=s�;�/>��>��	�L�by���6>#�>K��-����TϽ�U>� ����;Z��?s�b�t�_��0.�Wro�zB>�ND?_��>�,~=@Y?�Hc�P ̿�J_��jZ?er�?��?y��>E!߾�֖>Ǎ¾�]]?�w2?���>�{a���}��m�=nd׽QƖ=���3Gp�j�{>ʆ�>��=w�4�3�+������M>�[�>�2}ƿ�a$��@��/=?$g���`������	�]��B���n����Ti=��=��N>ev�>g�V>�5X>�BW?�"l?�e�>�>�o�ML����ξ�!�xB���2���������� �J'߾H!	�kB���" ɾ�=��K�=FR����<� �	�b��uF���.?��#>�ʾ��M�)<�Lʾ������j���O�˾;�1���m���?&�A?����W������������W?���6�������
�=8ٱ��F=�ɜ>P͡=}J⾩�2�2�S�+B*?�Y%?k���f��9�I>�2��/�W=A-?,�?<z=���>�],?+Z�t����/>�5>���>���>j.�='���$�ֽJ�?�M?B���Ǟ��w�>~���;`�
_i=�>YL&��X���U>>�<+K���_�����K5=��U?�R�>v�(�s�$��׃�x	��n�=%|?�?@I�>�m?x*J?h�<,Q��[�FM���=��b?"[?k��=>��塹�j���� ?f�J?H�n>�zn��X۾\����a?T�p?�?�F� ������
&�b�=?�p?}|e�訿���f�/m�>�o�>��>��<��2�>7�E?ǰ%��T��鴻��u6�lh�?Z8@�=�?_�����g���}�
?R�>��QŶ�]��;��1=��>\虾2`i�=�:�� ޽�O?���?���>Dꖾ8m�\>�=L)��w�?F��?������;%�!�m���@[:�.=�<��qP�h�/�HU��G�
�iV����<��>��@ ��4�>g1��,࿑�ѿ$φ���׾��}�?�?�>�}��ǃ�W_�7�m�qE���G���~���{>��m=��&���A������H�og�<���>|���&�>lE_�:���=��}�=�+Ғ><�>���>���������?��&��㿈���Q������?�?A w?$ٿ>��>JM�჈�Zz��?D�H?ʎ2?��=�$��13��e?�c_�B�O�'9��o@��W>�hT?;S�>����a>��>N�?��d>s;�nƿ)����iҾyǦ?D��?_y�а?պ�?,
3?�5�����������?��!�=��b?:>�ԗ�����$�	כ��>�w�>/=����|U?��Y�xC�b@���6�j��>m����3��R ���M�*Tq��֔��߀��n�?m.�?N�?~�|��.���?�&�>m2��������=ƬO>�[�>�x=H1 �J�>�n(�n�6�45W>H��?6Z�?��?\�����iX/>��?1Γ>�+�?	B(<y�>�x�>�|�>�l>?�g>��E>-�>?�Vu?��?k�(�-XӾ��=�~��65�u0þT���>� ?��!?J��>CH�<��&�Ck���Ϝ���K��J�k�6�M��A�Ъ�>폱>��>��2�����h�?����ؿ�:�,���3?J)�>�?����m���/]?�c�>���'⳿����4��t.�?N��?�x	?�Iھ�W뼏!>��>���>f�սz��������X0>,C?��=��_�o�G��>�%�?Sr@6W�?l�g�'? �����,�m�5������>Jp6?�����>��
?̚b<��`�t錄�[w����>67�?M��?�r�>P	i?񀿧�6���<�?��a?���>x��=�#��7C�<�?�|��P����� ??��@�9@��n?-/��^hֿ����SN��$������=���=�2>5�ٽk_�=j�7=��8�G:��o��=-�>��d>�q>
(O>a;>�)>���9�!��q��W���?�C�������Z�8��$Xv�Cz��3������ ?���3ý�y���Q��1&�@`�^H�=��U?�%R?�p?d ?��v��>\���E=$��B�=�ۆ>jv2?��L?��*?���=�ĝ���d��2��L���򇾎`�>�I>W%�>��>��>��_:J>��>>@�>^� >Yy$=�R˺/�
=�:O>r>�>���>�0�>�N<>[�>�̴��/��ٛh�w�D�˽V�?f��[�J��2���<��B����Y�=�b.?q�>7��#>п~�.H?Z����+���+��
>�0?aTW?�>�����JT��E>���j��<>w9 ��ql�v�)��*Q>�b?x�f>��t>q�3�]g8���P��`���t|>6E6?�Z��G*9���u���H�H�ݾ8M>vѾ>��8�cb�c�����4ci���{=|[:?i\?(ܱ�K|��Pv��Z��9|R>�s\>D=�B�=5�L>[�d��.ǽ?�G�e[0=���=@6^>?�	> n�=�b�>ݏ�X"�A�>��>l�(>�<?�'?Z𼙘�.b��N����>>�g�>=Q�>��>��N�Hr�=j" ?��>��A�2�Ž$&L��,��DJ>��彅o�3a��1��=�f�]��=���=$9�6G�~�h=��~?6��㈿x��h���kD?%)?��=oF<W�"�K ���H����?N�@m�?�	�'�V���?
A�?.��F��=a}�>r׫>lξ$�L��?Iƽ�Ƣ��	�d&#�S�?��?��/��ɋ�4l�4>"_%?ޮӾH2�>%"�������)Xv�6h$=��>��G?�����B�T�<��	?��?1�W���ȿ�t��&�>T�?��?�n�Ze���?�DP�>��?�
Y?ΰm><�ھ,WZ��ɍ>@?�7Q?��>t�) )�4�?~�?�,�?FI>(��?��s?�l�>1x�|Z/�!7��]����b=�>Z;b�>%X>%���veF��֓�Eh����j������a>.�$=��>�>佢2��U;�=��J����f���>(q>d�I>�W�>�� ?�d�>���>g=�u��$���͵���K?M��?E��e2n�nt�<V��=Ԯ^�Z*?�P4?e0[���Ͼ�Ϩ>%�\?P��?R[?�o�>����=��+翿 |����<-�K>-,�>�Q�>Y鈽I-K>9�Ծ>2D�5r�> �>�G��AھM.��0��IA�>i!?o��>Ϸ�=� ?��#?�j>3#�>�aE�9����E�Գ�>'��>�M?��~?E?�˹��[3��	��B硿Đ[�>N>P�x?]R?�Е>̌�������mE�A\I����q��?yrg?�8彠?�0�?U�??��A?�%f>���ؾbҭ���>i"?d��$hA���&��	�P�?-�?�;�>��?�:�Ͻ'���������C?q/[?�3)?Š�nsa��ƾ�=�<�3�c�G:�&�;
��:��+>+T>b����=�=�>wA�=h�q�T�8���-<5�=L.�>u]�=6;0�����<,?�G�܃�rޘ=%�r��rD���>$OL>.���ܪ^?}a=�y�{�����w���U����?(��?^l�?������h��#=?��?�	?D�>P���q޾]���>w��Yx��r��>��>7�l�&�+�������E����Žs��>H~�>t1?��>���>A�>B��������5��M��:0��-�H������z����o������վ�)l����>��:��>!�?X�S>�er>E�>]|=7Ί>���>���> Z�>��>g�<��=�7!=U"���ER?F���R�'����ﳰ�2B?�fd?h�>%<i����D���r?d}�?=m�?�Iv>wh��-+��l?2?�>_��lp
?~=;=��X�<Ce��������Y����>�׽:�M��-f��g
?13?ԍ���̾<׽��Pvn=II�?�(?J�)�� R��o�\�W��S���O�g�!a���$�b}p��⏿oX��#����(�j�*=͚*?��?3q��h�Z&���k��
?���e>���>B'�>�ɾ>OI>H�	���1�V�]��+'�P���E>�>fK{?�j�>m�I?��;?pOP?�{L?���>n�>鯾�a�>
L�;��>�E�>��9?��-?��/?!H?}l+?[�b>�����*����ؾC�?҄?M1?�	?Ŧ??Å�#XýGF��b`b��gy�h����Z�=���<>�׽S�t���T=��S>T?7���7��,���i>��7?�?�>�\�>�k��@z�} �<�+�>�x?�>I�����q�!��[��>Cu�?�l��=��2>���=Z���Ļ�d�=������=�?��`I��m�;�G�=���=�݇�N.�Y溾��:%��<�+?�?R�6>��=�,H�����0ľ=�_>���>6R>���>�*l� �w�"����(v�{��=�x�?�Y�?v(<4��=��O>��U��F��=���B�$�G>r��>?�?|U?��?�$D?��4?�� >���<��ඇ����� <?�!,?톑>��?�ʾ#򨿒�3�ќ?�X?�:a�L���=)�9�¾Mսܴ>yW/�,~����D��1�����t��q��?���?9:A�-�6�7y�%����]��T�C?��>�[�>,�>*�)���g��&�[4;>3��>�
R?=��>���>�̦?�m�?p\4��!������	5���ξ�,ݾ=[�>N�>,�?Gų?�c#?%�L>��/����4�>k讽������"��)->��q=e&>a�?E��>�=*��ש<�5ʾ�X|=��!>�:_>S��>�l>!3�=�?3�0�@?��>��ƾb�5�ʐ*�5�}>�=0��?�w�?��>c>�����\� ��m�>���?W=�?��s>"�뾖�v<L,0�B맾ѭ�b5�>��?������wT=a�v>s?i�?�c��O(�~�Z�z��?/?)
F??���H�d�Y���>��a��:\�v��\�����L�#j��{n�^Aֽ!�?���Ҿ�N�0���F��jо7�?ۯ�=���=$�L>%+�KV��]xd��8>��𼑪B>�=ݐ��<�&�=�:��=���<�R�=b�>�)���?H��>I6�>�bm?�)==�>9)�>��>��>m�?��3?�q>����	�羴�����=���%~x�ۨ��,����=���=7.�=���=�y(<���=v/޼��=yg,��Q�R��=�,>�]�;�Ԟ=���=I��= �f?�����˜�dCc���x>��H?*�Y>8;�;8���.?\Τ>鄿��ǿk�쾬=s?-�?
]�?���>@���x>�7��ܖP>�?�<?���-cf>�\=����X�>�$�>��9�*����?�j��?}�@7YX?����;7��r�<��6>��>1�R��}1�(�X�2p`��W�5�!?�2:���ʾ��>w�=��ݾ�Ǿ�#=Ȣ3>�~i=��! \���=�	w��==:�f=dш>�
E>�ؿ=v���:Z�=��H=���=s5P>����E�8�%�)�i:2=���=��a>��(>"��>���>��/?2��?F�G>!{þ��K�:_���)>ӷ!�д>�)�Qv>.�?��I?rc?�,�>H�=�|�=غ�>���>ؘW��{�aS־�r����>���?�<�?双>� (��ʽt�M��>n�מ�����>}~6?\l>DG>v�U��%���-�w���K:��!=�kr�W<V����c����#��=Vv�>���>	��>d�s>֢8>�G>��>��>�f�< S�=P辻9#�<4y��:*�=Sx��$m =-�ѼZ@��V�:h��),���>�;c�;s�^<�}
<(��=u��>:�>��>��=G|��l0>O斾�qL���= v��b�A�=d��~��.�>�6���A>�>X>F���>6��9�?��X>��?>3{�?Lu?< >�p��qվ,	��Qe�_�R��ҹ=�>��<��L;��`��jM��PҾr��>�D�>J�>XX>=y&��<��r�=W�Ҿal�[s?�Bb���8=4ќ��Xs��,���e��G�c�1�ټ(6;?����6f:><o?{�E?^}�?���>l�3NԾY��=a��j�ͼ����f�9�?�4)?���>�����H��q�;��t�|>S�]$n�㱛�>o��b���7�>/ t�UDо���e�k�'�{�o�*��਽���>�6?���?!j���;����3�(f�K�>a� ?�b8?=�G>G
?���>��ؽ7I־i�L�?<q�H?�T�?L-�?�s�=J�=����w(�>�?uX�?D��?`�s?
?O�'��>���<��	>A��cx�=
v�=y<�=ƻ=6T?��?o�?$k��S{����ү���,X���=F��=���>u��>�2p>��=�ه=��=��T>ݖ>�k�>��I>���> K�>�A����� v&?߷�=!�>�[2?^-�>��1=1۫�#��<Y�s�FA�Ga/��>���ս'�<z=���c=�Ĭ�c]�>�(ſ�>�?�F>�v��r?"u��5�&���O>�F>P�꽘��>g�I>��>�z�>`��>�>�/�>�Z)>�IӾP>����b!�:C��}R���ѾQRz>������%���������+I�dn��7a�cj�#���1=��@�<N�?c��[�k���)������?N`�>p$6?�ꌾ���1�>��>_��>�P������kÍ��5���?Z��?��d>?՘>!�W?�9?� 5�ef.��)X��Qu��?��ec��Dc�,ƌ�����\�	Y���/\?G�s?�e@?�5�<��w>�?��ꌾ(X�>\G1�[@���=Z�>s���i�nӾ��������+Q>�np?��?N?�J���n��
(>A�:?+~1?hIt?,�1?��;?�X��$?��3>SQ?��?L5?]�.?$�
?�1>�G�=7���8U*=�Ӓ�������н�ɽL_�)2=�0y=�&�m)<?G=!��<���'�ټ�);���o�<}b;=���=�0�=���>�M]?�=�>v�>ƭ7?���*S7��ԫ��/?�9=��|�^Q���դ��p�u>Zzk?8׫?Q�X?ñ`>¤B���@���>N��>�%>�A^>|"�>Xｇ�I���=(#>�$>Á�=W~Y����q
�`��v��<��>�?��*=���2^/>���p�3���U>u�Ⱦ��Ӿ?���t�%9�8������>F|`?s�?��=@ ���
,�:�z�FI	? �0??ot?x�m?S��=򾒾�`1��v8�ᲽQ��>�'>>{��/����d�=�qvZ=��>Y���
����\>�?�׾�$�n�/�L�����~B=W���^=�[��Ҿ�������=9J>E�����b������w�J?n R=	¥���^��Ч> ��>Zg�>��*�<x�Ԁ@��謾-ʑ=DR�>��J>�?����F�y�N�>ELE?r�`?棄?m���B�q�k�C��8��S����ڼ��?��>�?r6?>�:�=����d5�|rc�=�F���>|D�>���ڃH��ힾZr�c#�f �>�?�*&>9�?��P?Q�	?S=^?�7(?� ?���>���³��#7&?Ej�?V�=]�Խ�!U���8��E�d��>�)?��B��u�>�^?�?"�&?�}Q?��?�G>Z� �%@�졕>=r�>�W��a����_>��J?e��>�Y?�?�>>rK5�k���	����=�>a�2??#?O\?)�>ԣ�>P�����}=0�>��a?���?Myo?���=0i?��+>���>���=�j�>J�>R?�xM?5(s?`�K?�.�>m�<8٭��:���k��%�x;��.<��=m��~�d�G�
��p�<�Q���̼��ҹ��1G�wz��8�;�x�>4dl>���� I5>yþ~���V�;>�򷼚���^Ռ��S>�pI�=�N�>0�?��>\�%�C��=ۢ�>���>��'�&?:�?>w?��:IIc�+Zݾ�cN�F�>@�@?CV�=cfk��G��UVt��!g=�n?�s\?��W�'��0�b?��]?�0�,�<���þ�Vb�U��O?��
?^LH�d��>��~?��q?J��>xe��n�����Gb���j�^*�=4��>i��d��e�>��7?F��>��c> ��=&۾�w�v���z�?��?�?���?�*>��n��-�L/��Ҫ��U=^?2��>��C�!?<Q� �о��������n�ᾤ��;����O��l��w^"��\���kӽp�=b?2�r?�q?܋_?UK �dXd��]�=���JW�)�����|;D���C���A�2�m��C����ބ��@=�20���6�!ũ?
�H?4�'�`�>������\ؾ D=�5������>b,=���=riL=8y��L켇��`G?��>Mk?�#5?�C��D�l�I��R��%�<B1<$��>8��>�A?�x=� Ľ(d�<"!۾���=w�9yk>'Vj?�H?B�s?���+�'��U������ǽ1"����Y>��!>[�j>�����Q�ǈ'�d�;���m�M������xb�A�=@�6?_��>V�>I��?w��>�F�9��������)����<V��>�nq?���>�%�>������þ>װm?�#?�X>��Ⱦ�n*��C[���
r�>*�?�2?i�>�&��	rq�����2��Q��)�=-�(?{���a��3�>��]?�7N=9�<�->�üO��W�Gű�=�Ⱥ>z>WӲ=;���@.��Kt���Y)?;�
?�M����&��)�>^(#?��>ؤ>JÃ?b��>n迾)H��I�?A�^?e�J?"�B?��>�C�<r���*ɽ��(�!=Nу>�T>N�`=��=����^�����,?=��=��２����6<�6\� (s<H�=�=<>�{࿤�A�r�������Y�h�
�Ǭ��H�ݽҼ�����S-�����g�|�gn��-��iK:���<�!�����t�j��?̳�?�����z��>���4����辭ͯ>�����Av�M����̖��Yþ�8��9��i�7�a�V���^�։'?����8*ȿnȡ���Ѿ��!? 1?�Sz?�v�T ���8��.>�W=�_��Jw��T����Ͽ?𙾀�`?���>P��;���4�>�X�>c c>��l>q񄾚����<,�?�8,?�U?�j�(�ɿ�X��0���|��?�@FqA?�(�t����U=���>܍	?yj@>�0����Ͱ��Y�>G-�?uӊ?��K=��W��S��ve?��<�F�b�����=�	�=�=���{J>S��>�C��%A��s۽}B4>��>��^��e_���<�A^>K�ֽ[.���?-U��ta�K�8��Kt��'�=�.?���> Y�=�Z?�A�vLӿ�>N���W?���?s1�?n?��澷v�>b۾G�8?^�0?j  >��8��:���N�=�~:ǥ���q����`���=���>Dr�5����
�1�n�<ӥ>^��ſo�"��j��b=J�U�r��N���O�� ��o�l�[�齅�`=�i�=��R>;`�>��S>^<X>+�W?��k?��>
>�������p̾5�#�iK��S5����#�����4a�w�޾%��f���{�;�ʾ}U;��_�=4�R��#���[!���d��C�ҩ,?�.>��ƾ)7L�i�:<9mʾ�=����i�E �� gƾ�p/�5k��ܟ?�@?钅�f�W��d����&~���V?M���b�6���� �=����B0=�!�>�c�=a��/�2�(P�N<0?�'?B����푾��'>���;�=�A+?O�?���<�>��%?�!*�E��%�X>�1>��>���>�5	>�箾m�ٽ��?.KT?���#����o�>6-��7uy�uEf=l4	>�m4���ռ{]>�<�'���?��g�����<WW?ᦍ>'�)�m�_Y���H��J?=Ɯx?2�?�b�>Ɍk?BC?�͟<G���l�S���
P{=O�W?��h?k�>�����Ͼ!�����5?��e?UtN>�h���龎�.��P��!?��n?%?)/��R~}����6���e6?��v?��]��A��@�
�U���>���>��>i9�~��>�??E ��l�����C�4����?)�@Y��?��!<�! ��=�?R	�>�Q���ž\��������q=��>`����~u�����*0�bF7?$��?� ?-Ⴞ���<k�=�ە�#D�?9�?T���"Z<���t�l��x��y�<Fn�=��\����쾃17��5ƾf�
�!|������K�>�@�:߽�e�>8�'���/Ͽ'2����о��s�)p?�0�>�ýS�����i��Lt���G���H��ʍ��v>>�=�ʽ[W���'m�UpJ�La=Lu�>Ms��>>��u����B��:l=wх>���>�ԩ>œS��3��r��?�E�Hο����-�޾�_6?���?�z?8�$?�W>��v�����Ȃ�C�>?�Ԇ?�.J?&�ݽ��8��<L�j?�L��I`��4�wKE� �T>�!3?�2�>��-��~=yH>��>�p>�+/�U�Ŀ�ֶ�������?:��?�k�Q��>���?q+?�j�L9���h���*��"��>A?�E2>���آ!�=�wӒ�ԭ
?�`0?���0���T?�z�g��g�J�@[8>4�>��3�5�Fۖ���ǼW�x��~��8�k���?�G�?�1�?ۘ(�4�R��O?��>�ܾ0p��<t?��?}��9�9�=7/�>w�̾c��;�ƽ��?b?�?%a�>=M���ٷ��`>��?D �>!w�?,��=���>r��=�c��'OI��">k��=�3��;?�M?#�>���=�@��]/�%�E���Q���]C��>~�`?`#M?	�f>�.���)�X� ��۽�4����?���/���߽�:>L�@>>"B��oо��?Mp�9�ؿ j��p'��54?/��>�?����t�����;_?Qz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>A�Խ����\�����7>1�B?Y��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�f��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?kQo���i�B>��?"������L��f?�
@u@a�^?*ٲ�5����Nؾ�ʾO魼�f�6@>)*��z�=?U��b�<�	w=;�>�x�>{��='~>խm>�,{=���G)���)�����CL���^4���R����9��Ⱦ�:�����x��������I#�FMI��<;p �A�/X2����=3T?�7U?��q?��>� |��q>6l�
��<�E+��5V=�D�>�0?v�J?n*?���=-���b�	����%���E��0��>]�G>rK�>Ze�>�O�>`�p��=>'�<>J��>b��=�#4=ϼܺ��<A�H>�X�>ͧ�>
�>P<>�{>�ʴ�/����h�Yw��˽O��?.���o�J�P0��zA��n���	��=�c.?ѝ>b��<п�ﭿ�-H?_���(���+��>�0?�^W?S�>����ZT�� >����j��\> ��^l���)���P>�j?�i�>)�>����"O���Y�ܽž2�O>��9?�Gv��!b���d�W�u�^ѽ��*->�� ?/�g>���i𓿠I�g\���>2�=?mm�>�M��٨�|｟���h�P>���>���)�+>��&>�Q�y���qu�#	�=J>J�!>K�?��>��c=�>��D<`��G�>��0>8%>h�=?�?t����Ŗ�i�~��(�V�d>��>7X�>��>��@�H��=N(�>�e>l�t����C/���F�$VE>L
���wS�n�Y��=��H���=Qɰ=� ��8L���<i�b?�S��:z���u޾�o%?U)�?$��>�~�>��`>nu���Ŕ����p�?7'�?ο|?g�X�J�����I?��?$x�̼>��>Y?�Ҿ5� �P��>W&y�t2����)�E��?TN�?���-)��ob��g.>Rk2?���Ph�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?�M@>�M�?�Iv?���>��v��-�s���TK��z�=݆:;ٌ>cg>�|��G/E��{���o���d�a����K>-	=�>�d�E��N��=[⎽pc��-mC�^�>�ot>�b_>���>��>
��>P�>�]�<ؑ�����c픾��K?y��?<��� n����<ߙ�=b�]��&?�Z4?�!c��Ͼ{��>�\?���?t[?���>n���H��3ܿ�W_��f�<PkK>�'�>vU�>����3�J>s�Ծ�AD�i�>`�>=���TGھ����4��'��>T!?�H�>�2�=˘ ?�#?��j>"�>�bE��9����E�[��>��>O?��~?� ?:й��\3��	���桿Q�[��8N>~�x?wS?�Ε>Ì��퀝�-dE�LI�b
��a��?Nrg?vg�f?�/�?��??~�A?�f>���*ؾ����R�>�'?pP�����:���&q=c}%?@�.?U��>�T>щ��%�<;G�;k��L�%?��Z?�/Q?����͐� B쾠�<�Ľi��F��8%"<�0�=ٖ���=;R����=��K>�����?!D���
>���>}N�=��6���;�*?��;��{���$='?t�9,C�]_�>h@>�����?l?���j�\����$����|���?8_�?��?h���yd�L�:?I|�?�H?w��>P��bᾞa۾4Z_�:N������>3S�>�?F<���c�����{r����	6�L�3?�c�>��:?��>R'*>� �>��w���Y�6Ҩ��]������	��Z��E�օ�B\����5
��Fʾ��D��|�>il����>p��>�g@>a��>��>�@?����=�Y>�T�>H��>���>�=>���><Oc=����P�H?_��j�¾������>�o?�k=?��>|�K>~Ǉ��w=�]?l�?#�?���>b9l��-����>`�?US���?�E,>��E�V
l��|O��Ŏ��νL�1���%=��g�� �YW������>�(?",�>zS��R��=����_o=XN�?��(?��)���Q�D�o�$�W�AS�_`��h�=b����$�m�p��쏿�\��+"��5�(��*=̈́*?v�?���������8k��?�nf>��>o�>�߾>�aI>��	�ý1�� ^�cI'�徃�I�>�V{?�a�>NKI? �<?��P?��K?{�>ԧ>X'��d>�>��;�M�>���>}%9?��-?0/0?��?4�*?��b>�(�������׾-&?�?Kk?��?1�?�����1ǽ�l����M���x��!�K��=�H�<)�ؽ��x�NU=�R>��?�C����#�cs���6>6�U?���>_v�>S�HYʾy��e�>�?�A�>��#r��;�?�l�?�����Ƽ?��=�#>�̙=�B�y����H�<��=i�	>���=v)<�xu���<�������<�^���� =�C�O�>@G?j�>�K�;S"��2-Ծ�
�����=&s>�V�>5��>-}�$������3�����	>�	�?"�?z��9=V�G>Mv�5���.��
پ��\��"�>�&?��?+b?�3? �p?��<�4#�;b��΁b�����8?N!,?-��>`��f�ʾ�񨿒�3�\�?=[?�;a�`���;)���¾s�Խ�>[/��.~�c���D�⺅����|����?ҿ�?�A�F�6�y�ɿ���[��>�C?s!�>�Y�>q�>�)�$�g��$��0;>���>�R?���>S�$??�Ny?U>*�.�JĿ���ݤ��ڥ��د?�&u?��?'o?p��>�>|�a�ﰾ`���t.B��B��O�]����>z��>��?��>�1d>Q��$���q�/�l��=�K>P��>�R�>�͢>�n= �>��C1?�=�>K��x��f�G楾l�>FB�?��?R�-?��>�(��D��^��C>`��?:֐?��H?���9�>`��>��Ј:����> ՟>A*�>��=bR:�	�e<�?��/?�gw�D8�5�_�Ӫ�=7?m�^?Q�=�Iؿ��a�$�2�1D����B�nȡ��ґ�@D׽%Դ�ND�=�膾�e��:ᢾ�HU�5=��jvF�rN��rݤ���~��?y��=	�>��=�C<}޼x%�<Z=��ֽ�G=Y�
��<~6���4=;�"��,<���=:j�=1����1��p�?Z
�>>R?��$?Z<W��=,�C>�)Ҽ�V�=|�@?Ŗ�>M'�����rپC�ӳ�zǜ�:��ta��0�6+(=�t��">�4�>ʁ9>�=����<���W�c>�7!=��=�i�>�L)>�Ei=��&e�=;�*>gn?����K����Z�dr
�	g#?��>L��=������/?�m�=�"{��������H^�?��?�>�?D��>�c'�׭�>=�$-�o��=:�{=�&�>�á=`{���>KJ�>K��75��h���z��?0�@�R7?�8����ο�o>K->���=�XQ��]E��k��&Ͼ����@?fM>� z���NA>�F�=��wW����=9s>>>�=���t�.�o� >���a�=�.��޿g>�"v>N��=�i����<{��������>�&Ⱥ0�9|�^=��=>��<��>��->Q[�>ON?ίA?<�H?a:><Z]��qѾ�#�H:�>84�=?�>��ü��.>F*�>_�(?�"B?S�?�f>�(�9m�>뿂>͏B� ���b�jW��~�>�G�?��?��?Hdm>����+A���V���+��H�>�?>��>M�>���lI߿��)��/������#��
#=j�q�oUü��@�J}�;�½t�=���>�S�>��>��|>�!>�R0>7��>���=u=�\=<A<�~�=6J �뮒=ij�;�:q<1� ������T�"�[���FqC<u��il�;��<���=X�
?^�Q>?�>6N)�]�����=|�|�}7���W>L9����#]��q��7�U��A��Ϣ>�>6�+��x��jP!?��>��>�<�?t�?y��=Q��0W�57��a��兾�4��X�=~��!���5]���<�/���ry�>��>�ש>�Sr>�J,�ː:�V(=��־m�/��>0O��G����$�l�v�i��)0��?^b��"����3?e��&>Ԡq?��R?a��?o��>�@��
�Ӿ�2�=���Dk�Ա�-��������?��%?ʮ�>��例�4����S.�����>��<�k�E�tC����2�L��������>(��F��cd*�O5r����ƙ �^-��f2�>��2?K.�?`!W�|�U�'�{���9�W?P�N?�>xu�>��>zP���9־����65>5X?g��?�?��?>���=yeȽؐ�>�
?��?��?�,p?��>���>��Q��8>V������=�>N��=��=��
?�D?��?Hl���	����V�쾢�U��8f<vz=̙�>�φ>I�y>k��=!iR=��=)�S>��>��>^1]>E�><�>;����5
��?�H=RR>W?�ڄ>n�=�������.o׽
�;�;��͍�^���f�=���<��*=�q�;���>��ʿ���?@L>�n�o�?��߾�)V��->_�X>B�V��>FC>�,�>���>��>�>AU>[)>�FӾ�>����d!��,C�`�R���Ѿ�}z>����u	&�Ο�.w���BI��n���g��j�B.��L<=��ɽ<(H�?����"�k��)����F�?�[�>�6?�ڌ������>���>�Ǎ>�J��Z���Rȍ�hᾚ�?5��?-�b>W~�>^�Y?�M?44���3�*�Z�6?y�Ұ@��ud���`����5����E	��ϴ�6+`?þv?|@?�h<a�u>�>�?0^#�0����Ì>��-�F�:��=�5�> �����X�~-Ѿ����'���=>�m?]��?�5?�Y�8�m��'>_�:?ӝ1?�Jt?��1?J�;?��y�$?�W3>�??�m?ZK5?j�.?1�
?��1>
�=#���W(=�<������Q�ѽ�jʽ6��f3=��z=,����
<
�=ds�<�����ټy�;Ua��]n�<��9=1�=G�=R��>�/]?0B�>�%�>!�5?^D���8������,?�'=�m���슾���V���\>��j?��?<�X?2�]>��B�8�=���>}�>')>�4Y>sѭ>t��{F�3q�=N�>��>���=E�I�����s	�&����<q�>R��>W b>���=cum>��羾Hf�ۢ>�ϥ�rꅾ&K��*F��5���`�A9�>J?L6?�=KPԾ�����3H��B:?JmT?t&p? i?���=���J x�`>��h���;>T�\>Vؾ ?{������9�G���E�>�e���6<>���w����z�!�N�K�2����J�n��=���GHϾ2����=>7>\9���|
��%������~cQ?�w�=|����i�1P���v<>4 �>�J�>�3���Jh�>��ľ'��<���>��@>ؼ�;��ʾL:�4���W�>L�)?��h?V�?�◾A��
r�C)�Z��m�W��09?�O ?�?�2>;D�W�����׾h�v�d�D��>O=�>|:��Q�>�?þ� �
9��3>�K�>�,>�"8?Ũg?Z	?:7?�?�Y�>�TD>��P�ޤ��oB&?0��?���=��Խp�T�`�8�GF�Y��>��)?#�B�ͷ�>1�?��?��&?�Q?��?��>c� ��A@����>�W�>��W��b��4�_>m�J?���>	<Y?mӃ?�=>n�5�2��ܩ��=�=O>�2?�6#?ԭ?I��>���>"�����e=�O�>u�_?�o�?�{m?�;�=2�?��;> �>&t�=g��>I��>��?�
M?�bp?K?Q��>�h-<H����괽���"}�A��;��<�}h=D��4D`�#���=?&h<�����r����	���J��:Z���:���>��l>��Kt0>)l���v��UF>�<<x����sYW���[=�sV>=�?�˫>A��J�<�?�>N��>J��?#?[P?�?�Ҹ���a�?ؾ�6O�쪳>ޘ??!��=�:k� ����y�f��< ry?�]?	ڂ����)�b?n�]?g�=��þS�b�t��D�O? �
?��G���>Y�~?^�q?ݶ�>#�e��9n����hDb�P�j��Ѷ=q�>
Y���d��?�>��7?�O�>��b>��=ov۾g�w�&q���?�?a�?y��?1,*>�n�l4࿧$��sݑ�. ^?/]�>FJ��ݰ"?���<�Ͼp���ѯ��2^��ͪ�D��Q���tC����#�y��
�׽:��=9�?�*s?t�q?T�_?!r ���c�ؿ]�>	���EV�h*�6��wE���D�JC�3�n�y��O���b����C=y�q�j�>�&��?�I(?0n�'��>坾���~XȾ�d7>]2�������V�=7���G� =��J=�_D�L�-��·��?	�>���>��<?�a^�uuJ�T1;�Z 9��3��qH>��>6Х>��>�n׺�����ս9�Ͼ�8��������v>./c?��K?�n?q���p1�*Ȃ���!��i/�!=����D>�>L�>�4X��Y�&���=�u&s�r �X/�� �	���v=o�1?�T�>�a�>&M�?�?��	������w�D1���<���>C�h?�	�>B�>Q�Ͻb:!���>7�l?&\�>/'�>����6!���{���ɽ�^�>�1�>	|�>�.o>'X-�+\�Q���`��b
9��z�=��h?����k`��υ>p�Q?�D�:��K<�w�>�w�<�!���򾊳'�a>�?��=0b;>Qpž����{��U��J�#?!�?�e����'�'rl>t[?84�>y��>�=�?��>ɷƾ8R߼��?{Q?IDE?։=?���>nR�=xUf�O�޽\�!�[=�S�>zJ>@XL=���=��a O��3�g=��=B飼�T����9<-b��h��<�K�<iX/>
&ݿO?r����ֶ̾�8:�
�k�����K�����?񗼳׋�����q�֏ �pe���	�Sj�ۋ�-�F�]�?ް�?]1�,엾؈q���:�`��.�>���j[$� :�������������ߴ�x�J����(��B'�L�'?�����ǿ��:ܾ(! ?�A ?1�y?���"���8��� >�@�<�-��y�뾛����ο���^?f��>��0��5��>���>��X>�Hq>z���螾f/�<��?3�-?*��>[�r��ɿS������<���?$�@5�+?@�B��#Ⱦ�F���~�>I�>`��;6־Y�E���A�ZP�>bT�?Yc�?�.>�5���ľ鴍?*i+�v���;.�E>�O>3�5>�j�[��=���>]i�T����=F��=|G,=cS�ì_�*�����E>��d>����6 g��x�?`�U��[��/�3�~�e>>Y�R?��>�{�=�!)?��I�iiп��_�_�V?���?J��?nT"?��׾��>
hھ�+J?T*7?g��>Z2��t�nY>�A��B$��r¾o�J�⇹=!��>*n�=�9;��M��E�/�<��=����ƿD�$��V�Q��<g4M���\�E�齕ҫ��kS�4���o����>h=i��=ӴQ>>GV>[Z>�W?;�k?zҾ>"|>N%��t���ξsu�>c���1���������ߣ����J߾�`	�1�����ɾ~6���;�Q[�b����%:� �q�ۈH���?�T�<h����yG��ȉ<�u¾zޥ���<�`0�)����2���Y���?�0M?������f�c����%=�Z���N?f�;��x��Wþh=9r��(�;���>�{=���ݎ ���5��?��?оx$��#�]=��X��=��M?�?�?>��i>���>�V����R��L�>���>���=:+?�ǉ>R]��4c3��Y?�!R?��(����5>aР���ݽ���=��=�6\�������=��/��=?�1��=�0���ڊ=Y6R?���>�����6m��V�
��[���l?�f?\��>S|=?��?,�A�$G��������� ���_?^^?j��<�� ��a?��5��ʥB?`�N?���<�w$�F4��UF�+u��~�>�v?3�C?u��.�{����RX����)?��v?s^�rs�������V��=�>�[�>���>��9��k�>��>?�#��G������{Y4�Þ?��@z��?d�;<V �c��=�;?z\�>�O�?ƾ�{������4�q=�"�>Ԍ��]ev����R,�`�8?ՠ�?m��>.������i�>4��� ?D��?sp���4���Q:�vr���ؾ~V"<Cd�=�
�=4�=i"ܾ�6,�-��=ض�������9�q>��
@�,�=���>����Dq��h8߿�#���􎾤謽�`?��	?�����&���aE��W� Z�ssh�y������>UHC=�.=f�-�.a�O�@��M\=`T�>q���=h�.��b��e���3>�,�>���>��E>��j=��ɾg5�?l@۾��ƿ;ȯ�w���;b?�g�?���?��!? @O�'$
�>~���x��?\ď?:?��A��I\=ʉ�>$�j?�_��wU`��4�qHE��U>�"3?�B�>S�-�K�|=�>���>g>�#/�x�Ŀ�ٶ�7���Y��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>	���H�!�B0=�SҒ���
?T~0?"{�e.�t�N?��_�������M�t���-�>�(��!�Y᜾��K�l^m�WR���6��}��?T��?k�?�E޻B� _)?kӞ>����F��֚�c~
?2�?!�k=�#�>k�>�#!�-�+�\��=���?H� @�|?������7\>��g?�S�>��?F��==�>���=)���8�"��p">���=��=���? iM?��>���=X9� �.��6F��R�`��oxC�ٰ�>LHb?�`L?��a>n4����2��5!�'ν��1���+*?�)�+��P߽%64>.�=>΂>s�E��@Ӿ��?Up�9�ؿ�i���o'��54?,��>�?����t�����;_?]z�>�6��+���%��}B�`��?�G�?;�?��׾�R̼�>1�>�I�>$�Խ����b�����7>0�B?>��D��x�o�J�>���?�@�ծ?wi��	?���P��^a~�%���7�F��=��7?�0� �z>���>��=�nv�׻��C�s����>�B�?�{�?��>!�l?��o�Q�B���1=PM�>ʜk?�s?�=o���>�B>��?+�������K��f?�
@yu@V�^?c��������x�ܯ�rF_����EB�;1F�1h�=�2�=7s;�03=�T�=��M>�(�=}�S>�D>���<�n�=wځ���/�/���Z����a�lIK�qI�ؤ¾��aN˽�#�� ���:q�}�/�\( �]�%��Y�,�J���Y����=r�U?�R?gp?� ?�2y���>L���"S=
�#�Rޅ=>�>�c2?{�L?�s*?"��=n�����d�[[���4��������>��I>5L�>�/�>D�>�m�8�I> ?>�e�>G>�D'=^�Ϻ�D=��N>J�>´�>�i�>�D<>�>0д�2��I�h��w�p̽ ��?������J�x1���:��c����b�=�a.?Ƃ>����=п����2H?����(�ڷ+�c�>��0?<cW?p�> ����T��4>���W�j��i>�( ��ul�Ƌ)�q%Q>�l?L;g>��t>��3��r8���P�����؝|>� 6?�඾��8�:�u�y�H��ݾY�L>��>�s!�t*�W�R�~�Fi�E
z=V:?�H?�г�����t�O�����Q>kY\>��=~��=��L>olf�"oǽ��F��4=m�=��^>?��>	�u>�a�<gϩ>�ӗ��+R���>�u�>�k�>0F?\3?����D����)@�l�>$\�>:�>}�h>w�a�1��=��>���> s�]Ć�H%g�O�{���`>�� �'�/�a	�"U1=������V=�_=�����KQ���=�Jh?U���Gҏ��("�D�Y>�G?_��>jqv>K�&�I�@����ܧ��ʩ�?eQ@���?àS���@���"?��~?p񼽿�W���>�{�>{�J����h�>��F�v� =�C�\i��ߧ�?<V�?�o��h���̍�bk�>s6:?~�'�\h�>�x�rZ�������u�d�#=q��>�8H?�V���O�X>��v
?�?�^�ǩ����ȿ2|v���>I�?���?I�m��A���@����>8��?�gY?�oi>�g۾R`Z�'��>��@?�R?�>�9�'�c�?�޶?寅?��I>�V�?;�s?���>��z�{�/�Ϡ������4��=�};���>7�>N���aF�'����8��+Aj��;�	�`>�t&=͸>�G��!��H^�=]���2��1h����>�p>��L>��>�	?Bq�>
��>\�=����@C���閾��K?���?+���2n��M�<���=,�^��&?vI4?io[���Ͼ�ը>�\?d?�[?d�>+��J>��E迿-~��0��<o�K>;4�>�H�>�$���FK>��Ծ�4D�mp�>�ϗ>����?ھ�,��M��VB�>�e!?���>�Ү=� ?k�#?��j>
��>XE�O5��O	F����>װ�>�I?#�~?��?%ڹ��c3���Qǡ��w[���M>4�x?;?p��>5��������:���F��[�����?�g?y��I�?P#�?͏??��A?�e>��!ؾ����,��>��-?-����X������<R ?'��>�`?��>ƍ��Tm�q�1�*��x�?ϣ?�,?�<���K�Wa���A�<�.�<�w�=k�{�\5B�B;���=����~��=]�0>׮=�����G�#�������*�4?��>N��<6�'D,?�\B�ac���5�=��r��`D��&�>��L>�y����^?�A=���{����փ��`�T��?���?gb�?/��?�h�`=?�?l?�m�>����޾"m�BFw�~px��R�lg>���>e/`�	
�Д��ן����ѯŽE.6�3k	?46�>�Q?�o?��]>��>�j�����BԾW4��TBX����u�9�O�%���[���z|�I/�����3�G����>̼���m�>��
?Hx>�OX>�y�>���kp>[FK>:�>â>"�9>^�">��>��N��M�2S?�����B׾�뾟t��@?�U?N�?��������?K"�PV�>�:?�h�?x�0?}m���:a��??g�?���F��>��L��_<��>���r6L��ܑ��{i>J�?Ow��)�U�"�B�q���7)?�=?�N�C��]�Y>2����n=O�?N�(?��)���Q���o���W��S��x��g��@��g�$���p��菿;Z�������(�4*=�*?t�?S������/��/k�'&?�NNf>8�>�'�>o�>θI>x�	�2�1�>�]��F'�[ʃ��.�>�Z{?,}�>�I?��;?�nP?dL?�ώ>�`�>����k�>���;�>���>@�9?�-?�(0?�s?�o+?DRc>b�������zؾ{?�?�E?�?n�?ׅ�DCý)藼	�f�.�y�Ed����=���<��׽c2u��T=a�S>-v?�ֽg=��?�D>�-?b��>��>}�K��5/��A�%�>R��>_�}>�>��%S���z=?u|?�ソ;��<Ш>�=ꂺ�Mҷ�M]2>~b�=�7�=00�;���DQo=TԎ=U"�=l�'=Y�-=Ơ�<`�����<�h?ּ?�G�>{z>�9��b{���c �n��=6ǀ>��>2�>:��\Z��֮���]�U"�>�؋?E��?���=�r�=[�>�F��cY���E��H����ż��?B�?b�M?�V�?ES@?�8? -(>A��Ӕ�t����b����?H&,?Ѓ�>��P�ʾg쨿��3�M�?$[?�a�>��
B)���¾N�ս�m>C;/���}�o����0D�j���y��<����?˪�?'�C���6�@8�¶��N��X�C?4�>=L�>���>7�)�z�g�2���;>��>H�Q?�d�>�~?~X�?��o?�ݢ�]Y[�d���㛿��X�EX'=J�?��?Fٍ?�[x?��O=��M=�jG<��&��E'��Q��]�T�d�^E7<�">�ߢ>���>��>(7�<�A���A6������P�&>�5�>Y:A>�]/>�:�>��v�SK?���>������y
�5@����.>be?�a�?r�B?�e���?���c��36�C��>�%�?��?���>��G�=���=k7���V��XJ>�ޓ>8/�>)П=�(>�R�>��?�� ?�jL���.��m.�n�d�� ?�6?m��=0�п�t}���������)�����վg�v��K��6���	�=�芾��������[��?��Z�j�َ�.���Nm�0�?��J<1}E=>�&>��;LPQ�#m�=��9f��s`'=�Ǆ��g�P�м�Y�<��A�U0=Ix{=�	@=$K;q��y"�?yM?��e?+x&?ɬ?��>l�&>� #?���>���>��d��ߊ�5���s¼c�j;���LW=QM>��Q������>L�=�X >]�>�*�=���ז;�˙��b0=�Q�=���=�	�=�٧<���:��J=\�en"�w?2���1ם�oZQ�����9:?�.�>�׫=�iǾ��??Y=>%���s��7#��?��?B�?yr?s�h��m�>����!E��g�=�嘽e�3>�u�=��/�J5�>2@I>5n�A:���i���G�?b@o`??�Ƌ�SϿ�c0>�bL><֤=�j�S�=�(���c�w�D�a� ?m^D��x��>5=��޾Kܺ��ʑ=W�]>h@>����:C����=��ҽ�Z�<�i�=���>��k>�>�8T=�=T���H�=Z�=���F%)=�I�����=Ѧ�=��b>�AN>���>�x?�>1?�jd?⦸>�p�`;u����Ɋ>���=*�>�ʃ=�w@>�>f�6?}D?�yI?�a�>�=��>l�>C�+��=n����Z���(�<��?>�?�#�>5��;.�H��n ��J?�s����0?��/?X	?RU�>�U����3Y&���.����z�>��+=nr��RU�����:m��㽳�=�p�>v��>��>UTy>��9>��N>��>��>\4�<�p�=�⌻+��<� ��;��=#�����<�vżꛉ�u&���+�%����;���;�]<��;U��=qo�>�T>� �>���=�t����->�Ȕ��J�_�=4���\UB���d�R�~�-�-���1���>>�[>��{�͑��B?�VN>�B>>p�?�t?Q9>��+R׾�S��D
f��Q���=��>�j=���;�+"a��jL���Ѿ���>�ގ>�>,�l>�,�d#?���w=��gb5���>`{��ܼ��'�9q�!@�������i���ҺS�D?pF��W��= "~?�I?	�?��>���̆ؾ�;0>�H����=��*q�&g����?�'?g��>��9�D�m#̾���1ն>[�J��IP�fȕ���0���5��}��Ej�>	-��(�о*3��L��$Ə�AB��9q��Z�>ȇO?c��?��`�c���iO��������*�?/bg?���><?��?�Y��/���h��;�=Z�n?��?��?�>!/�=���xR�>��?ؑ�?]w�?h�n?�3���>��`;�L>�T����=�a
>U��=��=��
?N?��?R���T���龞6뾶�Y�^}�<[2�=���>�P�>��w>���=��l=�ǟ=��K>�Ӗ>�+�>;9]>xȜ>�J�>�@���%��|&?�8�=���>�2?���>�X=3~��#C�<`L�̍?���+��긽��ོ9�<�#s�aQ=��ȼ���>Pǿ��?àS>�M��
?���{�.��vS>ǘT>�߽I~�>F>L�}>��>V�>f>8�>=(>v<Ӿ�h>#���g!��/C�Q�R�k�Ѿ�dz>�����&�ԝ�	j��0KI�Xf���\�4j��)��32=�.�<hG�?�p����k���)������?h_�>M6?b⌾���)m>u��>뺍>�@������Gō��`���?w��?�Bc>��>�W?H�?�1�3��rZ�\�u��$A��e�w�`��፿�����
�����_?��x?KrA?���<7z>���?��%��֏�("�>/��#;��:<=�$�>�%����`�2�Ӿ>�þ�D��=F>O�o?�%�?JV?�WV�1��}�8>�7?]�1?j�p?º1?i ;??w�c�%?��>>al?\2?nd0?�=)?/	?ӆ3>/%�=�r�;tT=� ���Q�� �νj�Ľ:�ۼ�M6=�=��+�s/<*=���<V�м�I���,�: ����+�<k�0=0r�=���=ۈ�>��[?Z<�>��>c�&?�]�n�2�_�p��<?�>`m~��`��5Mɾ����)	>5tg?�?R�^?/+�>�]L�^Y�+S
>ـ>=)>T�m>�>����:Y���==�>&->��=�z�v����0���l��c��>���>^[x>�[���>(��F�v�g>I>�P*��]N��I��k9��R��w��>�9M?[]*?8n=�Z ���`��b���%?��:?p�??Yi?N�6=�Kɾ*�8�J�I�.Vݽ��>Y�;ʜ	���������;�/��"~=��t>ի��ݠ��Yb>P��8r޾ǚn�4J�/���2M=)�:LV=�\�վd9�M��=N!
>����J� �F��Zժ�80J?űj=|t��dbU��p��r�>m��>3�>��:�w�n�@������6�=���>��:>�t��e�~G�8��/�>c3J?vl?h�}?*�~��pd�8�=�فо�B�����?�ҩ>w�>̿>R�=�ݽ�x,��o\�k3����>�w�>{c�Z N�����������&�ޙ�>��?�m�>�?d�1?l?_n^?��!?�?0��>�SE�Oڤ�)d&?�0�?�+�=K/��h���4�g-E����>��)?}�*���>�?�q?�&%?"xK?G?d�= K��w�7��g�>}:�>��_��ӳ��5M>،M?�޺>,�Q?���?�Ev>��4��;��<�e�>�x>+p/?d� ?L?|��>���>Ң��{�=<o�>{�c?(��?Dn?��=7�?F�4>�A�>�=�=0�>�}�>�s?aO?�#s?^�I?���>���<vk��(���Eq��Ɂ�;$);a,<F~=�}�~g����^�<�<N����S�yռL^=����Y� <4s�>My�>��s�Bx>�����,>�t�)Tt�m���򽾠;=�HV>^-?���>�c�tJ<�Oq>���>aD���?Gk?Ԧ$?���=�l�LG���
\�>�;?~��= ��hᎿ�z�܂�={f?�>?�է����I�b?��]?�d��=��þ�wb�\y龖�O?��
?g�G��۳>��~?i�q?R��>�f�H:n�e��4b�C�j�۶=�w�>�[��d�N�>5�7?#G�>\�b>J��=u۾��w�.s���?���?��?��?6-*>��n��+࿷���V��O�^?��>h����� ?N��h�̾�$��'h������䬾Ԍ��a ��I���8� �������ֽ�=\?+�p?�5r?�u`?#�ܲd��Y�旁�`�W�X���P�C���D�qYC���k�N�������ԛ�^R=,�N��.I��=�?�g0?��9�2A�>�MǾ��ɾ���i��>��ľ��P��7�<]1)������=�4�J�!�]p��$?�(�>�9�>�G?��y�~�H�Nw�
:`����%L>���>��>���>����p��ⴣ�� �����Y/�C�>��\?��M?/4c?�J����~�(�*��Z�hͻ���=Go8=�"O>q/��� �;@'���<�{e{����F���(�����#>9-?%�q>p d>+��?��?�����ʲ���'�Q��H�9<�5@>��U?��>1��>LϽ/�I^�>�Gh?w��>���>�{��n)�ױw�H���⨴>>��>�?n�>N�V���K��挿�[���8C�3q%=ϯm?�tw��{]�!�c>�EN?y�<��k<�D�>d��R�d�s�6�4��={R?���=ME>b�Ⱦ�X��e�n}}���-?�^?�j����3�Qo�>aj7?p�?��}>��?��>`Ͼa9�<Y"?R�a?��>?F�2?��>��=��9�toҽ!b-����<�@�>�v^>{�^=�2�=kW8�/�V���K�!V
<�">��A����鲕��m����=�j	�!�'>�Ͽ�5F�ܖ�����Ѿ
�!�~0��5r�=3�����Ƚa����9߾'�����t�f),��6a��ゾv���:�8��?�?��@�$I�HC��F���p��.C��S��>��̾�P���zҾ-��S����}ݾ��0�O�zub�����>�<r'?%Z��1�ǿ/����^ܾ ?�S ?n�y?�8���"�=�8�# > �<����`�����3�ο�К�v_?�>n��c��>��>'��>r�Y>Iq>Մ���j��W�<K�?��-?���>Ԥr���ɿ�h���.�<��?w�@�A?��(�_��n�T=7��>֨	?n@>�1�r;�2)�> 8�?A�?�LN=_�W�aI
��qe?�u<��F��&�y��=�<�=k�=	��qxJ>JR�>%��jfA�z�ܽ˅4>�څ>@7#�-����^��
�<*�]>~�ս�Q��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=G ��Yʿ8s*�����zv=.鎼��.���ӽw ��\��=	�[��.������Nɴ<��(>�Jz>版>�d>� [>�_?׼q?�f�>��Z>���}���]���<=�Jپ���` g�Ļ��m���3/ �*���!��_��J�߽���@=�|�=��Q�5A���~ ��c�F�qF0?�>��̾��L�Qہ;�̾wC���#��p����];�3���l���?ÊE?�L��T?Y�	s�J3�s���(W?_�yG�y$���,�=�_��}5=���>�Ȋ=;�侫@4�~�P��u0?f\?k����\���%*>K� ���=E�+?��?�GZ<�&�>SM%?>�*�Q1��_[>*�3>�ԣ>���>�@	>���WV۽͊?+�T?)������ې>�a����z�ba=�.>�95�Z����[>3��<�󌾵�U� G���B�<��Z?���>6`���;������=��">mfS?� ?���>��8?cm?:~>T�����R����se��e4Z?�{?�l,>��<�u	�E�徦�C?w+�?��v>
�þ(��K���G��>�y?� *?}�ཱུ�g�c[��)����??x.v?��+�hI�����mZ����>�?,? �?̎i���V>�+t?���f�����˿JB�C��?��
@`�@��/��j��h����?e�!?0A�Q�뾗fn<��ľۃ˽�&?�U㾁?���W��#���?U�y?X�>1�ؾ��Ѿ�>/@���!�?��?A�̾6�x�9A�-ᄿ���k>#xL=�J}��r�{o�ee=�LȾ�B򾖦��O�ѽ"9�>�@P��2�>�o��'�ӿ���a���9I��J֎�4:/?���>�j�
?a���c�8����D�Q=I�U�����>�y>��q������{�,9��_��i��>/���!�>�[G�Y����Ӄ�<���>m��>:}>�?���1���?�����Ͽw��A��9Z?��?j߂?�i#?z�F=��{����o��<ML?�l?فW?���2J�N��/�j?����H`��4�!E�$(V>tD3?���>�x-��3{=A>��>B�>-�.�-�Ŀ�Ѷ�:�����?���?<��m��>�|�?w�+?�[�b<���M����*��ȍ���@?��1>���z�!�r	=�������
?_0?���.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?���>��z?��o>�)?k������Y��,# >��>/�� �>��J?x}�>��=TQ�Ěb���q�*���v�5�X3�>�^?�C!?d�>&dؽ���=)3��{T�u�C������;�����rÂ��J�>\`>b�=}X�<(<��^?i��h�࿃A��@�C�w�6?��K>�>�徵�ƾ�&o��HU?�ĥ>�(�=#������1���.�?7+�?4�?�˾���T6/>�T�>��>�h[�c��Y: ���>dFp?��׹������U��>5��?�R	@L��?q�����?=��n]��8>��<�߾j,|�5��=�z6?�&�~b�;&$?a=�[�^}���'e�Sy�>���?:O�?�ٻ>:b?�	b�.(!�׳]> �>�m:?-u"?ZJ>&�/�_�>�Q=?cc>�M摿`4���x?tG	@�(@\�s?�zÿf
ٿx����Ų��d��=�XP=
M�=����k=�ռSP=�C�=��>�1�> ��>��x>�LL>B�=Y��=8o���!�/T�����?��K�3�	��Y[����~��@���žCq���4�x�2~�� N�u*(����6�>L =?\^?��d?]� ?k��t�<g����҅>ip9��2B<�#�>��?�6%?.�!?t�>w;����o�}w�S��(Lʾ	�h>�1c>���>��>�s�>rS�=�Q�>�s�>���>1�>y>�x�=1�>�>r��>X��>r��> C<>��>2ϴ��1��e�h��w��̽7�?݁��y�J��1���9��򦷾�g�=	b.?E{>���?п@����2H?M����)�T�+���>��0?�cW?��>Z��O�T�9>ҿ���j��`>L- �G�l���)��%Q>�l?��f>�/u>Y�3�GV8���P��f���,|>6?.׶��Q9�m�u�[�H�$cݾ�fM>¶�>�F�Sk�����O�x�i��q{=��:?H�?� ��i1�u�f���8R>�\>n�=�.�=";M>��d��ƽ��G��|.=zx�=�K^>�M?��+>iA�=��>�/���>P��f�>CMB>9I,>�@?=%?7���ȗ�1g���-��"w>]:�>���>� >KJ����=a�> �a>%�맃�4"��x?�.�W>}�6,_�U�t��my=.��C*�=D��=�N ���<�D�%=��~?�x�� ㈿뾦M��"vD?0?鮐=�>G<."�� ���@����?�@:h�?Ճ	�1�V�d�?SB�?i��/��={�>ޫ>xξƜL�ӯ?"ƽR͢���	�w6#��O�?�?%�/��ȋ� l��6>AX%?��Ӿ�q�>ү��7��ϓ�  q�u�w=���>�<6?��	�hp0��g�����>=�?����;���`ÿ+wz�Wy�>Z�?�ٕ?+�K��.��P=��{�>���?�/?h[�<��0�Ŕ-���l>��N?�|Z?X.W>O��%R$��O?p��?�7�?���>���?�Rp?�0�>��Ѿ��M�����B�V�w�~�|�F����>9�>>����$��J��J~��h5���>�Z=iń>��
����:�;=�W��ϯ��G>�L�>	Z�=��=�o>8h?Ӑ�>x�w>�����P��RU��૽��K?�?���>+n���<���=�^�G?sG4?
�[���Ͼè>5�\?���?A�Z?�Y�>?���>��W㿿���#��<��K>�6�>�F�>�K���.K>�Ծ�3D��j�>oΗ>G���?ھ<��A7��D�>�a!?��>���=i�?¤+?;��>��>��T�1���si<��<�>���>Ls
?�w?���>p\־���%��[癿�ZU�)�>
ug?�B?�Ņ>.�+��0�7�,=\��q?5�u?;��=��>�Hd?�mQ?6�^?�>�� ���վ��	��ӿ>��!?��A�M&��?�O?���>}/����սwJּ6���|��^ ?�(\?A&?n���*a���¾�:�<��"��)V�f��;�qD���>ً>R���X��=�>�ڰ=nLm�E6�b�f<*l�=F��>��=�-7�Jt��L0?�{=n����>���nyD�Bj�>��0>�.��({?�a2��᡿�����ܬ�]d���a�?&|�?���?6v9��t��J1?|7�?�Z?O(�>��� �����A��Z�5�E���:>���>B�
>�
�М��[����ܜ��e��na̽rd?���>�'?S~ ?Ą�=��?�����d�������kH�k�,���2�_�<��输l{��ሾ:�D�]`־�2���>�>�����_�>��	?�C>�D�>�(?)�y=Ǜ>���>`��>C>9s�=V�>`!�>��i=gZ���W?P,Žd0�����H�o�?g��?L��5wi��_t�$�I��V? �?�ɟ?�	o=�il��*�"��>�0?���(8�>;�d>a��>�5�<�����\�Q���!�ˆ�=��%��!,��'r���"���>r��>�%Q��^�5{d��c��}��=p�?�6?��7��tQ�hmO��u�XWX�s�<��.������M<�A�i����B-��t�q�{D-�˯�<�?�z�?h)�����{���F`��:���n>�� ?\�0>�-�>��>�\���	~I��N3��������>E�?OW�>uB?��<?�P?�S?
`�>���>2m��Yo?#�<S��>�S�>ȶ8?��*?��3?��?��%?w�F>�	�|�������T
?a�?|?l�?h�>_��15Ž�<-�:��t�P���㹸=���=�X�d�<��L�=�'P>2
3?<=>�1��`?��<m>N'�?�p?Md�=���}{�;,��Z�>�][?\��>�� �Ubm�J}��?��?�߫���/=���<AF�=B�>
>7>3e4>�>�6C-=���ܐ��Y,>*`�=��
=�ۜ=���<]@�=Z�P���C=�t�>�?m��>�F�>�C���� ����L�=�Y>�S>9>6Dپ�~��+$��m�g��Wy>�v�?;y�?%�f=w�=$��=�}���V�����y������<ˤ?BK#?&UT?���?��=?h#?�>�)�fM���^����^�?q!,?z��>��|�ʾ��|�3�Z�?�Z?D<a�����;)��¾��Խ3�>�[/��/~����&D�S����������?῝?A�y�6��x辅����[��ΓC?!�>MX�>��>V�)���g�%��0;>Պ�>KR?8�>/;L?K�z?��[?�'Z>h�6������ڗ��[<9-6&>sGA?��?�0�?|ix?�$�>~�$>V "��<޾-���.��F��銃�A=�
W>���>i~�>J~�>��=a�ȽM��lP0��J�=0�b>���>px�>�p�>��v>���<i�G?���>8T�����D⤾*����`=�u�u?P��?�+?��="|�P�E�3=��W�>mo�?7��?1*?��S�5��=��ּ�ⶾ��q�<!�>�ҹ>�+�>�=�vF=U^>��>z��>�%�N^�+p8�	M���?(F?&��=ƿ�q��Mq��旾��^<H%��j�e�:e��t�Z���="����e�Ω��i[�-4���L���ᵾ?v����{�_��>k�=x
�=��=�1�<a�żDf�<naJ=�J�<[�=��o���i<K�9���ӻ�����h�ϴ[<�-I=6��3l����~?��N?��+?��;?�U>�l>�2�5��>G���S?&h>� ��D麾F9�1�����=BԾ xʾ\�J����>�����+>+�[><��=�"=�4�=XY�=tx�=m��(�=j��=�ü=K�=�>���=��>�6w?���5���4Q�Z\�j�:?;:�>�}�=��ƾ@?�>>�2������c��-?���?+U�?��?vui�Ud�>\��Yގ�Dw�=����};2>���=��2�֢�>��J>D��#K��x��*4�?[�@s�??�ዿ�Ͽb/>��7>�$>5�R�+�1�ʚ\�x�b��oZ���!?�H;��H̾�5�>,�=!.߾��ƾ�c.=��6>�sb=�i��V\��ߙ=9{���;=~l=�ى>�C>�l�=�2�����=G�I=���=	�O>#����7�<3,�D�3=���=�b>a&>3#�>���>Ʊ2?EDk?���>6�O���ؾq��㤦>I�>���>�ǐ=/b^>x��>)I?��H?��H?5�>,�<\1�>�&�>�T(��,b��1��W���P�?�S�?��>vھ=�$�H���:�/�X�}p?��-?�?c`�>���H��z�'�'�)�p�;���O� a]����=�>�OE=����G�ļ��7>�4�>.`+?�t�>�S2>Rs%>�� ;^��>D� >N}�Id=f.;B��<���s�=��B=ޥJ>�����L:��W��mt�#�:�?�=O'�;��=^<�="h�=���>B�==��>�̻�)پ��>���g�'�=�꺾n�^���z�4섿��9�5�����>�6 >��(�04���Y�>L��>V->�@�?Sq?��>�P�����󋤿�4c��x:f ��x>[>�󩾶9B�G�q���F�$�־6
�>�ԏ>c��>��o>%+�f1?�M�p=���/�4�z��>���R��-����o����5���zi���&�+ZD?���k_�=�F~?4�H?�я?8�>�"��G�׾�G0>Z偾7�=�6�t	r�
����?��&?�H�>����D�o8̾�¾��>>1I�?�O������0����÷���>�窾�о�"3�c������0�B��dr���>�O?E�?�Ab�C[��-aO����ㅽ�j?zg?�9�>^?�>?y��0Z�P���h�=��n?���?]:�?>@��=���$Z�>�P?w]�?�΍?�tk?:�/����>P�<b�">9Ǌ��C�=ݹ(>�>��>V?y?���>X�����	���ԇ�D1u��Д<����v�>2�>��>�*1>�uF=p��=1D>�^�>V�>R
u>���>� �>b'����h ?�2*>F�>̋?I/�>s��<�{�
��=M3�0�C�5�6�Hk:�D\���%3>�4>�=�@b���>p%Ϳգ�?��|>M��Z?&�F�9b�=�7 >ʚ�>�]
�N��>�o>�Ҟ>��?��?>`��=Ꝅ>�-�=Ҏ׾,R>A���#9��E�+X��5�����>�g�pw���3	��P�5�^���������o������CW���=�#�?�Ə=��|�ʰK��8��+?.�>��?�8�����R�����>���>Ɔ��)r������'���?��?s<c>E�>Z�W?�?V�1�u3��uZ�/�u�v'A��e��`�b፿Ü���
������_?��x?(wA?�C�<7z>���?4�%��я�;)�>�/��&;�V<=�+�>�)���`��Ӿ��þ=�iIF>m�o?�$�?�X?�WV���]=Q�y���5?O�4?VB�?��?��={,R>��o?�ۺ>��(?khR?g�?1&-?�j?�>�>q�>�Y���B��X:�r�m��F��U�k+ҽ
�ǼZ�&>nY��!M���S�Z<<+>O�l3>�����<�q�=�׶=2�=��>��]?hI�>Р�>�7?���k8��Ǯ��(/?�:=��������Ţ�>��>��j?���?�ZZ?�2d>��A�j"C� >�R�>�u&>�\>|J�>�N��yE��=`M>�p>���=��L�����	�mz���e�<�>0��>V�>#>^���*>	��4�h���I>!0{��L���JU��PO���5��#z�_6�>�F?1�?s=����卽��d���$?��A?�WL?�{?��Q=U�޾��.��>H�e�!���>�Ǻ�p�����oŞ���4���}:�r^>{H��:裾F[>�^	�m�׾�vl�6�J���߾�7=�	��ju=?����۾�s�i��=^:>2���4�"��i��PZ��ЧI?ʘ�=Ӣ���X�D5���>��>���>�?���u���<�.������=U��>�{8>,/���kﾥD�� ����>g�0?��_?ƺ�?�N��,G���%���о"�ľq�>X��>�.�=:�?&�m>��z<#>ž� ��U��z1�`_�>���>tU�~�L��< �D��t-���>I?9?*b`>�*?��<?��>�e?�f?ܙ?��>"�ün o��*?^ց?H��=��1����>�q@���?&�2?���l��>K�?J�?m8$?qF?��?��>S���9�5�O�>5��>7�^�)���Z�m>�S?y��>��U?4��?[��=��.����s�[�(�x=��>S�6?�%?H�?���>��>Q ���=` �>��b?4E�?��o?�Q�=�?_`2>+��>r��=�>z��>V�?�/O?9�s?��J?���>���<	���I���q�W�@���;z(L<#�t=�����p��+�|��<ׇ�;�����<z�f���^E��񍼧��;h��>�`z>5>����=>:7����N�2nR>K3��%Yj�"�_�񺛾&�4=Q��>�	?i��>��:��"+=܍�>��>����-?$�?�L?�ݼ�n��پ���"%�>?D-?��	>k�h������8��le�<��e?�yM?!�k����l�b?�]?>h��=�@�þ��b�[��h�O?f�
?:�G�A�>��~?[�q?I��>&�e��9n�����Cb���j�>Ѷ=Hr�>[X�c�d�)@�>��7?�N�>s�b>o$�=fu۾�w��q��s?��?�?���?�**>.�n� 4�"?��V��f?��>���Y ?{ʽ�W¾�ޛ��5���޾�a��l��S����ƍ�s���ݐk���»=]�?��n?/dh?h�f?	��jj�BY�	�E	P�2��l���E��@�b�6��zp��+"�P��cXP�<6���_}`�䇵?l9?�𽿶�>_����+վݾ(�?>�/��F��"�<Y����=���=�t/��$����T ?�5�>\e�>$FB?��`�P�C�K�,���9�/󾞣c>��>*I>��>��<��I���W���6���� ���j>�PI?w�O?�؍?��=��9G�U�L��LS�t��2��2�>�f>�{8>0?��{����N��PG�a}`�2�^"M��@�8[9�7Y6?��>y�E>�W�?�?lI��K��už8�V�t^>�&j>�/y?4�>0Y�=m��<� �ˆ�>z�l?p#�>�ǡ>ꃌ��s!��$|���ν�f�>��>�'�>-�q>�-���[����q����9�)S�=cNh?0<��]a��T�>&-R?��)9|-E<N]�> w�0�!����A(��@>�s?���=t=>Mlž��{��,����M?!�)?y����;����>|�g?��?�
=^�?���>D���D��=I�,?��?'H+?�x?���>E>>��[>O�����?��1W=��>x%�>4t�=Tܾ= ���#��K<�V�����1��=Y�>Cۏ=���_0��/ż�S�>g�޿��P���ݾ���M�U"��ɞ�ZϽ�O��y�	��<߾���Vn?�-󽃭�;J=��y�D?���;��<�?^��?�O�����&����y��U��~�>�k��3��䓒�W�����#���㷾�!���S���b��sX��L?�}�7Oſ@���־�m?"?��u?�-�H{�v�1����=Ω5=����9c�\b���ο쪒�M�^?1��>I�߾�0�����>�9�>���>�^�>�2���D���4=5p ?�>/?��
?
�p�(ƿ����4=�2�?��@�A?��(������U=r��>7�	?��?>+Z1�LB�^���IP�>g;�?��?&�M=��W���	��}e?��<�F�"޻L�=�<�=�W=����J>7V�>#���TA��+ܽ�4>�Ӆ>2g"�~��ot^��+�<�]>��ս(7��2Մ?%{\��f���/��T�� U>��T?+�>�9�=��,?P7H�\}Ͽ�\��*a?�0�?���?7�(?ۿ��ؚ>��ܾ��M?oD6?���>�d&��t�|��=�6ἷ���\���&V����=Y��>a�>ق,�ڋ�ˇO��L��]��=J��m!ɿ��"�E$���<@�v^��h��y�㽪�g�C�̾�`���a�x�=a->�df>ѳl>��>���=i�Q?�7y?�\�>#צ=��%���������:S�+a���14��+����1����+����(�;6�K:��8־�lD���W=�.Q��Ɛ������`�&H�_)?%>({Ⱦ"�P�p���Չ���ɥ�%x�ű��L3Ӿ_;6�Ys�j�?<�F?u@���,U���e���C��t�W?w������=��~�=��:�>+�<-	�>=/}=6뾵�,��G�3�0?o?ċ�����_*>����\�=ك+?ή?�\<(��>�A%?��)����?H[>�3>Fޣ>��>Y
>��$۽�m?�[T?�� �=���Wܐ> Ͼ�ފz���c=�V>v�5��n鼈�\>��<g���3W����<#|r?5�>\c��'�n,��o=� �=�%�?b*/?��W>3�v?�uO?��>k�����C����!>u63?)h?��>S\��mF�	�	�m�k?�^�?���>���q�ᾊ@8�~?
���?�l?
3?4��=z�Y���h��1���w$?��d?�pD��/��e�
�U�.�_��>F8?��?�cI�GS>3?I��=C����%¿�-��h�?�@I@+	��3��\؁<�M'?���>_%ʾ \��3@P�@M��������>�����}��P�z�B���J?l2�?�
?剾���Ū=iF˾m�?�ڂ?Ի�����)���]����"@��q�=<i\�r������3��1�3��f�ž~j�|�~>s@E�7�@�?�q���ݿ�Ŀ��}�x�/b���(0?��>�_@�a�I�{{��+~��M���T��,�%��>��>}�m���&���պ>��4)��x�><Q��� �>��<����	��f~�<�؎>��>�r�>���s����?����Ϳ}��<	���W?�ƚ?���?r�#?��<;a�%?g�Ԥ<�9�B?��o?�S[?g주��S�ly�,�j?S_��XU`�ʎ4�'HE�vU>�"3?[B�>�-��|==>P��>h>j#/�N�Ŀ}ٶ�1���3��?��?�o����>{��?�s+?�i�8���[��_�*��V,��<A?�2>.���?�!�r0=�<Ғ���
?*~0?�{��.�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>iH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�M�>J �?&��=�V�>��=����$(�3s">Se�=�>��?	&M?si�>%�=��8�j�.�i6F��+R�����C�� �>�	b?�+L?d�b>�H���t5��� ��ͽl@1�U�
�?�y�1������3>�=>=�>D�x�ӾY�?U: �6�ڿRE��kn�ɘA?Q�>�%�>h�ؾY�M�|T5��O?�	�>�\��m���������I�?��?�?侍�2�'3>Fr�>Z�>Z=�J�f�5�2�(�=�K;?M�=Ӭ�����!a�>���?�@Э�?]�Z�O�?'辺E��FQ|��Ҿ<��.�=��<?�Ѿʎ->�(�>�Ci>HoR�Yo��ԫF����>N�?��?��?��g?<�h���1����=q�>�/D?>�?�S�=�	��r�=�?:sž{�������5{?��@q�@mju?�#����ؿ�	���������b&>�
�=��C>�_�;Ǎ�=�>b)��w\x�\��>��>jl�>���>�CU>|��=D����\�����1ʘ�dLH������������6[���x@��վ���v=���=����ylu�a���$;��
>ZIP?�uS?�yi?��?ՐW�7$ >�����j=4����f;�!X>��0?�GF?��?G]=W���^��'v����������>�E/>��>���>��>�	=U�E>2�4>#�>�c�=۞K:�ὼ�x]<�cN>�a�>c��>�ߘ>F�>��>����e��|e�
=� j�f�?4���=SH��L��eb��� �����=��,?���=Ȋ��O�ο�a���LI?𓀾v5�:!4��>��/?p�Y?}3>�5���R��V8>�`�n����=Z ���YA+���f>=s?կf>u>Ϙ3��c8���P��|��Da|>�/6?1趾%B9� �u�W�H�E\ݾCFM>4þ>�D�>m�������ji��{=�u:?��?_1��Mా�u�8���IR>`3\>A�=Q[�=fFM>��c�g�ƽfH��6.=���=G�^>AD?,>�M�=�p�>�ę�k�Q�r&�>�@>��(>P @?�$?���ھ������a.�yt>8B�>�>��>j�I��_�=���>�{`>)�������>;�)W>f
}�ޥ^�&}�d�u=+U�����=�w�=�5 ��<�� =2�~?�[��{؈����h��D?�1?C�=U�S<NQ"��
�������?��@�[�?׆	�X�V���?.V�?P~��ڱ�=7��>�.�>�ξ�OM���?�!Ž`⢾e�	��#��.�?J��?�q3�Ұ���k�W�>`%?S�Ӿ���>[���o��r���e��ѻ=�Y�>"L=?6L���Y{�pDJ�>��>�?H�ņ����ǿ��z�@Y�>Ap�?X�?�`����*�'�w(�>�H�?��E?V�>>�ۥ�S�>�pu>��O?t�Z?D��>6�JF���V#??G0�?9>Ot�?Er�?wc?��:�L��pȿ���r�V>�N�5�?A>�>���Z������҇��\�&A��))>5�=��>*�Ͻ/!T���J=St;�)�v�r�L�+j�>R|E>�	>�`�>h?-��>D��=�%�����-��}�H���K?���?����.n����<���=z�^�i#?*I4?�O[���Ͼ8Ϩ>R�\?���?�[?a�>���<=���忿���e��<j�K>`0�>+I�>�2��W<K>�Ծ�4D��m�>Yӗ>����gCھ�1������FA�>Uc!?=��>���=�&?V�?\��>���>O�j�.Η��{*�w��>���>� 3?Y��?���>�R��Q9�}��Xӓ���I��I>/\k?Ҕ?5Y�>��������ݱ�w��;9�5�?R[y?-����?�Ɗ?��-?�W%?5�K>M��%��:�-�4�>��!?���A�QN&����?�Q?���>�*����սSAּI���z��8?�'\?\@&?����)a�g�¾�0�<��"�v�U��#�;lD���>̏>4������=�>�Ȱ=�Rm�D6���g<�p�=�|�>8 �=*7��p��o�?�pV�m~��bm;f�~�̃/���L>j��>H�
�^P?�m[�����ڲ������ת=�d�?���?�X�?���=zg��%?_��?��?�)�>��`���þ����{�y|���*�� �>
�3=�/�
��x�����
���>L��F�>���>93?��?�E�=�>�>�5�!�&�e:�������C��&��S@��%���j���Ͻ���r罾�{��ܩ>GR5����>��>���> ��>!��>���4�>�Z�> �>aq�>vq�>�~>#��=L��8���Ԧ[?�G��a!� "־��K���V?4�_?��>��=F�^���*�p�?���?��?>�a��v �=h�>0�*?X�����>Ø)>F">�U��Ͼ���*�,�d<3ս��c>e;5��b7��7�Bp��-�?��?����5����"�ΐ��9�y=�3�?��-?��$���R�Mpt�Y�S��YQ�����^"�}��I�,���h��ŏ��Z��o�����/���<�"?�G�?���++Ծ������m��B��nN>G��>�1�>K0�>�Xl>���K���m[� ���(����>�|?��>��H?��<?/'O?��L?<W�>է>r;����>W�<�>��>R:9?�!-?��-?D?V�(?\\>v����r���!־�4?eL?�?�o�>�8�>����]п�Yz�������u�0���^�g=���<�ҽ(�t�ktg=TpF>��?�����8�2%����m>�8?�5�>���>�?���5�4�<���>SD?��>l���=r������>��?���[��<�}*>0��=��v�db4����=YKϼs�="hw�J�N��<���='Ŕ=�nD�b�Ⱥ�B���W�:'K�< u�>6�?���>�C�>�@��0� �b��f�=�Y>BS>�>�Eپ�}���$��u�g��]y>�w�?�z�?ӻf=��=��=}���U�����F������<��?@J#?(XT?`��?{�=?^j#?͵>+�iM���^�������?�!,?��>m��1�ʾg�I�3�۝?�Z?�;a���<)�ؐ¾��Խ4�>y[/�C/~����+D�y���������9��?⿝?�A���6��x�z���+\���C?�!�>eX�>��>��)�;�g�%�+1;>��>�R?ܱ�>:�O?z^{?0�[?ͱS>�8�7T���+���>�b@?��?�5�?��x?�>y�>��*���w������<��!7���we=�W>��>���>��>/�=��½�౽��>��=7Xa>?��>�e�>���>��x>��<u�J?&]�>e��LN	�A�ƾu?��W�K�ږ~?�Ӓ?��2?-Ϭ=���CA�F���ɶ>�̥?L��?Vj&?��?���>;�d�ɾ듛�hI�>�f�>�j�>���=�y=S`�=S�>��>���x�5����={?i1??���=�Vǿ�k�}J�� l���+6�����W�������;�k�ky�=��O��m���qP��U���熾�rž\:��#
��F�?��	>���='T�=�o!<v`ؼy2;=7�=ʳ<�T�<��<�T���ɴ��)���\���(��-u=s.=�����o?�eP?��?��Z?��r>��=g�ʽ)۰>��p��0�>��=�X�:����H�e��=��Vġ���ξ��ľ~ {����6>�1ͽ���>�10>��<�x=lv.>��=x(>�H�<T�;(>���=��=|�=�xI>�:�=�,w?j������Z1Q����)�:?�M�>?��=ѱƾ�@?��>>�'�����z�9G?g��?�]�?I�?�i�PF�>����b������=e�����1>�S�=��2���>�K>r���T�������#�?�|@�?? ދ���Ͽ	R/>��5>�>�?R��61��Z�N7b�V	Y��!?8�:�hξ4�>m7�=R�߾�pǾ��,=�6>1e=)5�U\�R�=f�� �@=�m=�.�>M�D>��={�����=Y�J=j��=�Q>^�+�ͬ.���"�<�;=P��=��a>��%>Ȉ�>j?��0?Eg?]h�>�X���Ѿ�⚰���>�A>Ⱥ>w�$=D�9>�4�>��2?Pf??&)E?$��>���=և�>�Z�>
�.���s����d��:�]�<j�?e�?\ú>w�`=��$����b:�L���X�?��6?0�	?/�>�U����8Y&���.�C����16��+=�mr�RU������m������=�p�>���>��>Ty>��9>l�N>��>��>�5�< p�=�䌻;��<� �����=������<�uż=�����&��+�#���,�;Ч�;#�]<P��;&�|=R��>��>���>y �=�<��
��=��G�I��k뼃񼾱8B�Ȱg�m?����-��k'�~�d>��f>B����ϐ�W�>��>4DA>�N�?`?g?<�W> s˽6F���̭�c(�Z���;��=��>B����qH�ǜc��OD��Ӿ���>%ڎ>
�>5m>� ,�	!?�ZWy=Z�rf5��(�>�����d�����%q�C7��i�i���ߺ�D?r>��h�=�~?��I?@׏?qj�>T����Aؾ��/>�;��--=��}�p�s�����?�'?܀�>���D�$�˾�k��K�>��G��PP�ӕ�e80����.i���g�>P���BѾ�2��*��Xߏ�mB�n�r����>ߏO?�ܮ?��a��U��E�O�+�.��>�?h�g?,�>OV?�?������;��#��=!�n?ó�?�$�?i>��=V����>�z?I9�?�<�?�q?�@����>�۞;�t>�ӛ�/�=��>���=��=ts?��	?�
?%+��n&
�_�ﾱn�b�X��d=�M�=
�>-��>\}r>�O�=��l=� �=��`>��>w�>��e>���>\ǈ>�XҾ�!�S�%?Gy�=�.�>m3.?��[>^`>,(�?Uo��2=/�=��D��nE�D����F>й>Ct�=}$�U��>�Ͽz�?Of>!=���?%��2���5�=���>rн�֦>j]|>�>��>�X�>�->�� >>b{�&�)>�@���;�(�4��I=������0�>��a=����=ޘ�z�6������ξ��e��-����;��h����?�D�;�f��@���n ?��>E*?y.���J;U>eT�>ϲ>��ӾԳ������,�վs�?���?�;c>��>I�W?�?Ғ1�23�vZ�+�u�k(A�*e�V�`��፿�����
����+�_?�x?/yA?�R�<':z>Q��?��%�[ӏ��)�>�/�'';�@<=t+�>*��%�`���Ӿ��þ�7��HF>��o?;%�?wY?FTV��2��,>G�<?>,?ˬ}?�V.?x7/?kj�P�(?�?>��>S� ?!3?�
-?�d?��>�z�=����!=/M���j��MȽ��߽��;�S==H=|��<�=&%=(fV=b��`z��
�=�q<ڬ
=�f=�b�=��==��>`�]?�H�>I��>��7?����o8��Ʈ�f,/?Џ9=^�����
�����t�>��j?���?�_Z?�dd>�A�C�K&>dY�>r�&>+\>�]�>�{���E����=�L>�^>%ϥ=� M��Á�@�	�����>��<�!>�K ?��>�2���5>񴉾	�Y�2�m>`�i��C���<��FR�<03�g~5����>O�C?�?fA]=�$�"+��d���!?JcJ?��E?Qq?��;�U߾Ts&�.�F�X$*�a��>
��:�0�����	`��e�,������i>�ξݠ��Yb>P��8r޾ǚn�4J�/���2M=)�:LV=�\�վd9�M��=N!
>����J� �F��Zժ�80J?űj=|t��dbU��p��r�>m��>3�>��:�w�n�@������6�=���>��:>�t��e�~G�8��/�>c3J?vl?h�}?*�~��pd�8�=�فо�B�����?�ҩ>w�>̿>R�=�ݽ�x,��o\�k3����>�w�>{c�Z N�����������&�ޙ�>��?�m�>�?d�1?l?_n^?��!?�?0��>�SE�Oڤ�)d&?�0�?�+�=K/��h���4�g-E����>��)?}�*���>�?�q?�&%?"xK?G?d�= K��w�7��g�>}:�>��_��ӳ��5M>،M?�޺>,�Q?���?�Ev>��4��;��<�e�>�x>+p/?d� ?L?|��>���>Ң��{�=<o�>{�c?(��?Dn?��=7�?F�4>�A�>�=�=0�>�}�>�s?aO?�#s?^�I?���>���<vk��(���Eq��Ɂ�;$);a,<F~=�}�~g����^�<�<N����S�yռL^=����Y� <4s�>My�>��s�Bx>�����,>�t�)Tt�m���򽾠;=�HV>^-?���>�c�tJ<�Oq>���>aD���?Gk?Ԧ$?���=�l�LG���
\�>�;?~��= ��hᎿ�z�܂�={f?�>?�է����I�b?��]?�d��=��þ�wb�\y龖�O?��
?g�G��۳>��~?i�q?R��>�f�H:n�e��4b�C�j�۶=�w�>�[��d�N�>5�7?#G�>\�b>J��=u۾��w�.s���?���?��?��?6-*>��n��+࿷���V��O�^?��>h����� ?N��h�̾�$��'h������䬾Ԍ��a ��I���8� �������ֽ�=\?+�p?�5r?�u`?#�ܲd��Y�旁�`�W�X���P�C���D�qYC���k�N�������ԛ�^R=,�N��.I��=�?�g0?��9�2A�>�MǾ��ɾ���i��>��ľ��P��7�<]1)������=�4�J�!�]p��$?�(�>�9�>�G?��y�~�H�Nw�
:`����%L>���>��>���>����p��ⴣ�� �����Y/�C�>��\?��M?/4c?�J����~�(�*��Z�hͻ���=Go8=�"O>q/��� �;@'���<�{e{����F���(�����#>9-?%�q>p d>+��?��?�����ʲ���'�Q��H�9<�5@>��U?��>1��>LϽ/�I^�>�Gh?w��>���>�{��n)�ױw�H���⨴>>��>�?n�>N�V���K��挿�[���8C�3q%=ϯm?�tw��{]�!�c>�EN?y�<��k<�D�>d��R�d�s�6�4��={R?���=ME>b�Ⱦ�X��e�n}}���-?�^?�j����3�Qo�>aj7?p�?��}>��?��>`Ͼa9�<Y"?R�a?��>?F�2?��>��=��9�toҽ!b-����<�@�>�v^>{�^=�2�=kW8�/�V���K�!V
<�">��A����鲕��m����=�j	�!�'>�Ͽ�5F�ܖ�����Ѿ
�!�~0��5r�=3�����Ƚa����9߾'�����t�f),��6a��ゾv���:�8��?�?��@�$I�HC��F���p��.C��S��>��̾�P���zҾ-��S����}ݾ��0�O�zub�����>�<r'?%Z��1�ǿ/����^ܾ ?�S ?n�y?�8���"�=�8�# > �<����`�����3�ο�К�v_?�>n��c��>��>'��>r�Y>Iq>Մ���j��W�<K�?��-?���>Ԥr���ɿ�h���.�<��?w�@�A?��(�_��n�T=7��>֨	?n@>�1�r;�2)�> 8�?A�?�LN=_�W�aI
��qe?�u<��F��&�y��=�<�=k�=	��qxJ>JR�>%��jfA�z�ܽ˅4>�څ>@7#�-����^��
�<*�]>~�ս�Q��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=G ��Yʿ8s*�����zv=.鎼��.���ӽw ��\��=	�[��.������Nɴ<��(>�Jz>版>�d>� [>�_?׼q?�f�>��Z>���}���]���<=�Jپ���` g�Ļ��m���3/ �*���!��_��J�߽���@=�|�=��Q�5A���~ ��c�F�qF0?�>��̾��L�Qہ;�̾wC���#��p����];�3���l���?ÊE?�L��T?Y�	s�J3�s���(W?_�yG�y$���,�=�_��}5=���>�Ȋ=;�侫@4�~�P��u0?f\?k����\���%*>K� ���=E�+?��?�GZ<�&�>SM%?>�*�Q1��_[>*�3>�ԣ>���>�@	>���WV۽͊?+�T?)������ې>�a����z�ba=�.>�95�Z����[>3��<�󌾵�U� G���B�<��Z?���>6`���;������=��">mfS?� ?���>��8?cm?:~>T�����R����se��e4Z?�{?�l,>��<�u	�E�徦�C?w+�?��v>
�þ(��K���G��>�y?� *?}�ཱུ�g�c[��)����??x.v?��+�hI�����mZ����>�?,? �?̎i���V>�+t?���f�����˿JB�C��?��
@`�@��/��j��h����?e�!?0A�Q�뾗fn<��ľۃ˽�&?�U㾁?���W��#���?U�y?X�>1�ؾ��Ѿ�>/@���!�?��?A�̾6�x�9A�-ᄿ���k>#xL=�J}��r�{o�ee=�LȾ�B򾖦��O�ѽ"9�>�@P��2�>�o��'�ӿ���a���9I��J֎�4:/?���>�j�
?a���c�8����D�Q=I�U�����>�y>��q������{�,9��_��i��>/���!�>�[G�Y����Ӄ�<���>m��>:}>�?���1���?�����Ͽw��A��9Z?��?j߂?�i#?z�F=��{����o��<ML?�l?فW?���2J�N��/�j?����H`��4�!E�$(V>tD3?���>�x-��3{=A>��>B�>-�.�-�Ŀ�Ѷ�:�����?���?<��m��>�|�?w�+?�[�b<���M����*��ȍ���@?��1>���z�!�r	=�������
?_0?���.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?���>��z?��o>�)?k������Y��,# >��>/�� �>��J?x}�>��=TQ�Ěb���q�*���v�5�X3�>�^?�C!?d�>&dؽ���=)3��{T�u�C������;�����rÂ��J�>\`>b�=}X�<(<��^?i��h�࿃A��@�C�w�6?��K>�>�徵�ƾ�&o��HU?�ĥ>�(�=#������1���.�?7+�?4�?�˾���T6/>�T�>��>�h[�c��Y: ���>dFp?��׹������U��>5��?�R	@L��?q�����?=��n]��8>��<�߾j,|�5��=�z6?�&�~b�;&$?a=�[�^}���'e�Sy�>���?:O�?�ٻ>:b?�	b�.(!�׳]> �>�m:?-u"?ZJ>&�/�_�>�Q=?cc>�M摿`4���x?tG	@�(@\�s?�zÿf
ٿx����Ų��d��=�XP=
M�=����k=�ռSP=�C�=��>�1�> ��>��x>�LL>B�=Y��=8o���!�/T�����?��K�3�	��Y[����~��@���žCq���4�x�2~�� N�u*(����6�>L =?\^?��d?]� ?k��t�<g����҅>ip9��2B<�#�>��?�6%?.�!?t�>w;����o�}w�S��(Lʾ	�h>�1c>���>��>�s�>rS�=�Q�>�s�>���>1�>y>�x�=1�>�>r��>X��>r��> C<>��>2ϴ��1��e�h��w��̽7�?݁��y�J��1���9��򦷾�g�=	b.?E{>���?п@����2H?M����)�T�+���>��0?�cW?��>Z��O�T�9>ҿ���j��`>L- �G�l���)��%Q>�l?��f>�/u>Y�3�GV8���P��f���,|>6?.׶��Q9�m�u�[�H�$cݾ�fM>¶�>�F�Sk�����O�x�i��q{=��:?H�?� ��i1�u�f���8R>�\>n�=�.�=";M>��d��ƽ��G��|.=zx�=�K^>�M?��+>iA�=��>�/���>P��f�>CMB>9I,>�@?=%?7���ȗ�1g���-��"w>]:�>���>� >KJ����=a�> �a>%�맃�4"��x?�.�W>}�6,_�U�t��my=.��C*�=D��=�N ���<�D�%=��~?�x�� ㈿뾦M��"vD?0?鮐=�>G<."�� ���@����?�@:h�?Ճ	�1�V�d�?SB�?i��/��={�>ޫ>xξƜL�ӯ?"ƽR͢���	�w6#��O�?�?%�/��ȋ� l��6>AX%?��Ӿ�q�>ү��7��ϓ�  q�u�w=���>�<6?��	�hp0��g�����>=�?����;���`ÿ+wz�Wy�>Z�?�ٕ?+�K��.��P=��{�>���?�/?h[�<��0�Ŕ-���l>��N?�|Z?X.W>O��%R$��O?p��?�7�?���>���?�Rp?�0�>��Ѿ��M�����B�V�w�~�|�F����>9�>>����$��J��J~��h5���>�Z=iń>��
����:�;=�W��ϯ��G>�L�>	Z�=��=�o>8h?Ӑ�>x�w>�����P��RU��૽��K?�?���>+n���<���=�^�G?sG4?
�[���Ͼè>5�\?���?A�Z?�Y�>?���>��W㿿���#��<��K>�6�>�F�>�K���.K>�Ծ�3D��j�>oΗ>G���?ھ<��A7��D�>�a!?��>���=i�?¤+?;��>��>��T�1���si<��<�>���>Ls
?�w?���>p\־���%��[癿�ZU�)�>
ug?�B?�Ņ>.�+��0�7�,=\��q?5�u?;��=��>�Hd?�mQ?6�^?�>�� ���վ��	��ӿ>��!?��A�M&��?�O?���>}/����սwJּ6���|��^ ?�(\?A&?n���*a���¾�:�<��"��)V�f��;�qD���>ً>R���X��=�>�ڰ=nLm�E6�b�f<*l�=F��>��=�-7�Jt��L0?�{=n����>���nyD�Bj�>��0>�.��({?�a2��᡿�����ܬ�]d���a�?&|�?���?6v9��t��J1?|7�?�Z?O(�>��� �����A��Z�5�E���:>���>B�
>�
�М��[����ܜ��e��na̽rd?���>�'?S~ ?Ą�=��?�����d�������kH�k�,���2�_�<��输l{��ሾ:�D�]`־�2���>�>�����_�>��	?�C>�D�>�(?)�y=Ǜ>���>`��>C>9s�=V�>`!�>��i=gZ���W?P,Žd0�����H�o�?g��?L��5wi��_t�$�I��V? �?�ɟ?�	o=�il��*�"��>�0?���(8�>;�d>a��>�5�<�����\�Q���!�ˆ�=��%��!,��'r���"���>r��>�%Q��^�5{d��c��}��=p�?�6?��7��tQ�hmO��u�XWX�s�<��.������M<�A�i����B-��t�q�{D-�˯�<�?�z�?h)�����{���F`��:���n>�� ?\�0>�-�>��>�\���	~I��N3��������>E�?OW�>uB?��<?�P?�S?
`�>���>2m��Yo?#�<S��>�S�>ȶ8?��*?��3?��?��%?w�F>�	�|�������T
?a�?|?l�?h�>_��15Ž�<-�:��t�P���㹸=���=�X�d�<��L�=�'P>2
3?<=>�1��`?��<m>N'�?�p?Md�=���}{�;,��Z�>�][?\��>�� �Ubm�J}��?��?�߫���/=���<AF�=B�>
>7>3e4>�>�6C-=���ܐ��Y,>*`�=��
=�ۜ=���<]@�=Z�P���C=�t�>�?m��>�F�>�C���� ����L�=�Y>�S>9>6Dپ�~��+$��m�g��Wy>�v�?;y�?%�f=w�=$��=�}���V�����y������<ˤ?BK#?&UT?���?��=?h#?�>�)�fM���^����^�?q!,?z��>��|�ʾ��|�3�Z�?�Z?D<a�����;)��¾��Խ3�>�[/��/~����&D�S����������?῝?A�y�6��x辅����[��ΓC?!�>MX�>��>V�)���g�%��0;>Պ�>KR?8�>/;L?K�z?��[?�'Z>h�6������ڗ��[<9-6&>sGA?��?�0�?|ix?�$�>~�$>V "��<޾-���.��F��銃�A=�
W>���>i~�>J~�>��=a�ȽM��lP0��J�=0�b>���>px�>�p�>��v>���<i�G?���>8T�����D⤾*����`=�u�u?P��?�+?��="|�P�E�3=��W�>mo�?7��?1*?��S�5��=��ּ�ⶾ��q�<!�>�ҹ>�+�>�=�vF=U^>��>z��>�%�N^�+p8�	M���?(F?&��=ƿ�q��Mq��旾��^<H%��j�e�:e��t�Z���="����e�Ω��i[�-4���L���ᵾ?v����{�_��>k�=x
�=��=�1�<a�żDf�<naJ=�J�<[�=��o���i<K�9���ӻ�����h�ϴ[<�-I=6��3l����~?��N?��+?��;?�U>�l>�2�5��>G���S?&h>� ��D麾F9�1�����=BԾ xʾ\�J����>�����+>+�[><��=�"=�4�=XY�=tx�=m��(�=j��=�ü=K�=�>���=��>�6w?���5���4Q�Z\�j�:?;:�>�}�=��ƾ@?�>>�2������c��-?���?+U�?��?vui�Ud�>\��Yގ�Dw�=����};2>���=��2�֢�>��J>D��#K��x��*4�?[�@s�??�ዿ�Ͽb/>��7>�$>5�R�+�1�ʚ\�x�b��oZ���!?�H;��H̾�5�>,�=!.߾��ƾ�c.=��6>�sb=�i��V\��ߙ=9{���;=~l=�ى>�C>�l�=�2�����=G�I=���=	�O>#����7�<3,�D�3=���=�b>a&>3#�>���>Ʊ2?EDk?���>6�O���ؾq��㤦>I�>���>�ǐ=/b^>x��>)I?��H?��H?5�>,�<\1�>�&�>�T(��,b��1��W���P�?�S�?��>vھ=�$�H���:�/�X�}p?��-?�?c`�>���H��z�'�'�)�p�;���O� a]����=�>�OE=����G�ļ��7>�4�>.`+?�t�>�S2>Rs%>�� ;^��>D� >N}�Id=f.;B��<���s�=��B=ޥJ>�����L:��W��mt�#�:�?�=O'�;��=^<�="h�=���>B�==��>�̻�)پ��>���g�'�=�꺾n�^���z�4섿��9�5�����>�6 >��(�04���Y�>L��>V->�@�?Sq?��>�P�����󋤿�4c��x:f ��x>[>�󩾶9B�G�q���F�$�־6
�>�ԏ>c��>��o>%+�f1?�M�p=���/�4�z��>���R��-����o����5���zi���&�+ZD?���k_�=�F~?4�H?�я?8�>�"��G�׾�G0>Z偾7�=�6�t	r�
����?��&?�H�>����D�o8̾�¾��>>1I�?�O������0����÷���>�窾�о�"3�c������0�B��dr���>�O?E�?�Ab�C[��-aO����ㅽ�j?zg?�9�>^?�>?y��0Z�P���h�=��n?���?]:�?>@��=���$Z�>�P?w]�?�΍?�tk?:�/����>P�<b�">9Ǌ��C�=ݹ(>�>��>V?y?���>X�����	���ԇ�D1u��Д<����v�>2�>��>�*1>�uF=p��=1D>�^�>V�>R
u>���>� �>b'����h ?�2*>F�>̋?I/�>s��<�{�
��=M3�0�C�5�6�Hk:�D\���%3>�4>�=�@b���>p%Ϳգ�?��|>M��Z?&�F�9b�=�7 >ʚ�>�]
�N��>�o>�Ҟ>��?��?>`��=Ꝅ>�-�=Ҏ׾,R>A���#9��E�+X��5�����>�g�pw���3	��P�5�^���������o������CW���=�#�?�Ə=��|�ʰK��8��+?.�>��?�8�����R�����>���>Ɔ��)r������'���?��?s<c>E�>Z�W?�?V�1�u3��uZ�/�u�v'A��e��`�b፿Ü���
������_?��x?(wA?�C�<7z>���?4�%��я�;)�>�/��&;�V<=�+�>�)���`��Ӿ��þ=�iIF>m�o?�$�?�X?�WV���]=Q�y���5?O�4?VB�?��?��={,R>��o?�ۺ>��(?khR?g�?1&-?�j?�>�>q�>�Y���B��X:�r�m��F��U�k+ҽ
�ǼZ�&>nY��!M���S�Z<<+>O�l3>�����<�q�=�׶=2�=��>��]?hI�>Р�>�7?���k8��Ǯ��(/?�:=��������Ţ�>��>��j?���?�ZZ?�2d>��A�j"C� >�R�>�u&>�\>|J�>�N��yE��=`M>�p>���=��L�����	�mz���e�<�>0��>V�>#>^���*>	��4�h���I>!0{��L���JU��PO���5��#z�_6�>�F?1�?s=����卽��d���$?��A?�WL?�{?��Q=U�޾��.��>H�e�!���>�Ǻ�p�����oŞ���4���}:�r^>{H��1c߾�~>w����u?v��d�)6����d<8����;c6��!���!�3�=(�F>�В�X)�!���j=���JX?�!M>$4��5I��0྽�<�N�>��>����Gv��B^S��l�p��=��u>Î)>sd������g�S�_oƾ� �>�B?K�^?�Ǆ?ą�]zp��+;�48��\Т�0�a�/?X�>� ? �=>���=챲�h�u�d���C�߭�>;(�>{S�߹E�E����?��J����>�?�r4>d�?'�S?"N?7Y?�(?�?�)�>�^���^���B&?���?��=��Խ��T��8�5F� ��>�)?g�B����>��?w�?��&?e�Q?��?��>�� �i?@�۔�>pZ�>�W�d���`>��J?���>8Y?�ԃ?��=>��5�M梾4����v�=��>m�2?�5#?��?ׯ�>���>��@M�=h��>�Â?BP|?�Y?�X�>�?�?>"T�>�6z>�S�>��
?ݗI?ptv?�ˁ?��=?��i>63�<����&��N��=XK�=���<?��=���;R3��&�ם<=G��
�<�ep=Ha*=�=z>�;��`��>�_�>%a
�X~A>�z�p䑽&+�=w]��tb�'k9�Q��)�H�&��>�E!?��a>.d��a�ɻ�?�>��>s����>��?�@?j�/=����ʡ�kH~=-�>�X	?���=co��6���7j�9>�P?"1?Y7��f����b?^?A��6H=���þP}a�B�sO?��
?D�F��h�>b�~?� r?��>��f��Gn�h��b�a�>�i�悶=(Y�>)v�j�d�p��>��7?�<�>�sa>m��=��۾s�w�`���
?�܌?��?�ފ?*>#�n�x࿢o۾���|�Z?���>�Q���?$��{þ��Ծ�釾�������!ߠ��F��z�+��<?�������<�?!C^?\�v?o�i?���w'i��t^��dw���U��q�����yS�b�8�:Z,�-���~�.�*, �M軾u�<�!u���B�V��?n-(?E\����>�̖��例��,Z1>^���N|��l=V����U =.�i=�?��1�Sv��*|!?�;�>W��>��>?�hd�-=<�%l,���;���H?U>HM�>��p>	�>k�=O�I����LҾ�����ԁ�> fS??�W?��f?>�����!�� �����NŽ6UA�f�*��5l�Q�=JZ�H\ܽ�H,��Z�*rt���>������v +���-?�Mg>U�#>�t�?'?���CF�jՃ��]�f��=D�=�T?�<-?�@�>�E�ƽ+�ғ�>��l?Ҙ�>�ܠ>8Ì�%;!��}�7�Ͻz��>mL�>���>c�m>�X/��[��<��à����9����=Qph?�Y����a��҄>�4R?�#;L�@< y�>?�x�}1"������*��>�?S¤=j�;>�þ��2�z��Ŋ�c7*?�$?���[�-�W�>�O&?d�>Ճ�>�߃?�ȝ>�fȾ/ѻ�i?#�_?�GE?Ve<?���>��G=����hʽ�d&�)=�t�>��a>C��=�.�=�� �H�]�Yw&���/=��=����V��p[v<_����{<o�<o�2>�ڿ�T@��]Ѿv����龟��d���E��]��gS��蠾��о^�S������I=k���y�⊽�}���	K�?1|�?��� Fy�0㗿�uu�����"y>���W̄�>����!��Rs���H�q��U�7��F]�� ���_|�?�X�����@	���T���k?7�+?��m?:��=,.�ڊ1����=�:<���� ����9�˿Yۢ�p�a?D,�>4Ծ���	��>-�f>1J�>IŇ>�𧾝H����<h�?�g7?h� ?|�[�6̿<���煑=���?��	@[�A?��(����ohT=V��>"�	?��?>��1�H4��ذ��!�>H.�?3 �?E�N=Z�W�^�
�^oe?�<C�F�"�߻J��=�A�=+n=���J>X�>Ʀ�ulA�wܽ,�4>�օ>?9"�g��`b^�x��<[�]>\�սe@��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=?��A�ſ�N+��h+�E�;���������쳽e�`��XF�|���R^�p\м��>Q�g>���>��>�R>�)">��_?�΂?�U�>��>S%A�Z��g�۾�����М*�`,J�-�����Y��f�徘���1�o�5���7t=���=ĝQ�����OK!��oc��tE��.?�K >��ʾ�N� �;��Ⱦ���d�~x��� ;g3�/o�X��?B?����V6V��#����x]��hX?�P�E������.��=Y���=e��>6F�=^
�__3��+R�A0?�L?�m��h$����*>ǀ �B=�+?�1?H:<{.�>�f%?�/,�,��ƤZ>��3>N��>���>;p>e>��pkܽ'�?![T?�W�����Ŏ�>����~y�K�c=�v>�b4�[�)5]>ʙ<(���}�J��Џ����<$�a?V+�>CD�w�D���ž�
>7!3=s�,?$)?J?�D.?ny?l�v>U�Ӡk�L�!��|���~d?�u|?� >뮈<6����Y�f?l�?WcV>����ھ?B���0��V�>r]Z?c�B?bc<�q*`��Gt�]H־��?p[z?�I+��}�����������>�d?�?lxG�Ac>=C?e
>ԉ��hͿ�J ��x�?�*@���?gc�����)=��.?p
?l����m�$��=��q��z��< ?�O���i_���оW-��&�.?)[?5��>�v��R��)�>5+���z�?+�?린�梻"��Sz^����������=�79�����b��2�G��ھ.�_���5���̀>�@�/���>΍��x޿P�˿��s����Q\��1�,?�Ƃ>��h�㦚�0�m����[o���@�3	!��Q�>b�>ީ�������{��r;��b�����>4j��A�>��S�/���M���w�/<�J�>���>���>�3��2���磙?�����οs������A&X?uY�?1L�?^{?�Z<��s�DPz�1�#���F?Rs?&�Y?	%�48Z���/���j?Es��r�_�z:5�LD��"`>'3?@�>�+�;�=*V>T=�>vE>,�,�K�ÿ&ö�L�����?*j�?��v�>�?]�,?�\�|���1����(�oZ�B�@?F�/>*�����!�<�S����
?�v/? ��u�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?c$�>��?lo�=�a�>Jd�='�4-�[k#>�"�=}�>���?z�M?�K�>�W�=��8��/�;[F��GR�M$�<�C��>�a?�L?�Kb>���8 2��!��uͽ�c1��O鼡W@�=�,��߽U(5>��=>�>n�D��Ӿ�W%?�Ǿl��v��������MO?���>@B�>"���`H��Q=�P�?,�>,$��1���Fn�H�`����?A�?iO?�^��b�[	>ǣ�>x�<>v0���ƕ=�3���C�=�<5? �<�b��3:����>��?���?,ȱ?6l�� ?N!ھ����y{����}��	O�=��-?N�ܾ���=M?k�s>��s��Ű�ƪr���>̮?/Y�?��>ж\?��b��:+���=���>��3?�
?>L��oz1>'�?�>��������&u?þ@�9@(�o?Ϧ��P}��į����h���U�=��m�Y�8=9v��n�=Q%+=D}<��$;=G>�E�>�|>�:�>��>���>Rs�=!���;�!�����U}���@�]��u
����F&��MM�^��Y྅x���G�ކ���y��\��]6��l�����=XE?z=[?_`?(?ưm��
>�BԾ��[=�\����=#�X>?K�8?	?J�>:]}��Wa�V|�0ɲ�����ۚ>� >:_�>��>�i�>d̦<�s>�5>�A�>yd�>1�=Z�
��є��B�>�G�>5a�>�F�>X�=��_>����������o�S�ܾ���<ׂ�?墫��R��G��A���K���?=|P,?�[�=G���k׿;��4E?y�Q�pJ�!�6��z�=�/?��I?�L>>��T�>�>�">vP���搾dN�=®J��x��'�%�@��>{<?�hd>Xv>\�2��[7��P�m����>�6?V�����:�=&v��	I���ܾ��K>Jx�>m�P�����J����~�Lte��I�=��8?��?�ζ����	�o�M����S>�S[>5
%=�q�=�G>�"h���ýpJ���$=��=Md>U1?��+>�#�=��>�䙾buP���>`>B>A�)>f�??�M$?�b�gF������,��Fu>d��>|�~>IZ>��I���=FA�>�a> [��[����
��>��X>�t���[�d|q��Zl=X?��+Y�=�!�=x� ���9�4�,=J�~?�w���∿�#뾘I���zD?*?8v�=M�G<�{"�� ��XK��L�?��@�f�?�	���V���?AB�?_��ì�=؉�>?߫>ξ-�L���?j�Ž�Ƣ�ԍ	��,#��N�?��?��/�ŋ�+l��5>�W%?�ӾE�>�v�;2᛿ڇ�Bc���>�?�(?nVϾ�]+����O�>�j?$mվ�8���Nſ&�k��=�>���?e�?�IN�3���q�%���>c��?N7E?�e�<��}�����ӛ>�z?t�O?Ā[>^�6�z�L��F1?ҽ�?^ݎ?��X>ߎ�?��?���>9����3�{�ƿ�Or�ۛ+���X���?�=�gQ�,���5��]ԑ�A��Y�5�Q��>��<;��>�j���E ��7}>�]c��U���NY���?ĉ�>��A<	~�=��?�	�>��>�ꔻ��d���W�#Y��b�K?ײ�?8���/n���<���=5�^�L%?|I4?K[��Ͼ�Ϩ>(�\?���?�[?�b�>'���=��i翿g�����<��K>m/�>�H�>�#���OK>��Ծ�7D�;p�>�ؗ>�P��};ھ�/��գ�)K�> g!?ޑ�>5Ǯ=� '?%�&?�,i>�o�>[^����E/�Q��>)��>'�Q?*2�?���>�D������km�2ݜ��X��Ҏ>��x?9&?L��>$�������  U�h��=�䛾'�V?r��?8��=���>x�x?uj?��^?ߊ��i'���C��_0>x��>��!?���ݕA�&��
e?�Z?���>�ϓ���ս��ؼ7��������?##\?�"&?_���0a��¾���<܁!���b����;��I�Di>�>^��\ȴ=�a>�ʱ=bm��6�V�d<�8�=s\�>���=x�6������0?�=�H�����=8����$L����>f��>I�ߞd?X6W��E6�O␿Z�������W�?���? ��?B���)q��U?�+�?ݔ?���>�ۥ���J-��/��G�ҽU��&����?�>��>��$	�❿$���n���� �b���J��>�K�>��?'?�(2>��>�%�b�����\��L�П+�a�0�}<�h{�`D��c+=��۽��Ⱦ�}�&��>��*�>5��>���>)�+>��>�y1=i��>��>f�>y��>���>�i�>PB>��6=W��wX?�:#�Ϛ�<�X�w�pz�?��S?�5�<49�=��>�E�0�d*�>�Ρ?S��?�@�=�[v�&����?np"?m�����>�t�>p�o>�1��k�W�潁1�<Ko�6y>����/�0�A��F&�Ŝ?���>,b��i����B�Lt�'L�=�?�?h�F?�6���S�Ls��66� o����d�z����E�hd��C�����j����,��=ѫ?��?��־n���>����g�	�-�+"]>�T?#qq>��?��f>#�0��|��.+��K(����N��>��?�!�>�RD?{�>?#�L?/tO?^S�>��>�'��p�>e��<��>���>s�2?�+?��*?bc?h�)?�N>D��ů���ᾮ�
?'z?C�?%��>tG�>�����p��`ț<��W�Xd"����=�<Щ��i�뉔=k[T>Y�-?,WU=�D�.}<�4��>fl~?���><��+�߽�29��6R��}>� ;?�A�>Wv�6y�=�����?���?�q|�M}�W0O>~0	>1��=];>.��=Z[����7=,@�+���_�<�E>ܛ�<1>�q�;�ŗ=!�"��p=�t�>��?Ⓤ>F�>9A���� ����g�=
Y>�S>R>�Fپ�}��H$����g��Yy>�v�?z�?�f= �=	��=�}��	W�����	������<��?K#?4YT?���? �=?�i#?��>�*�PM��"^�������?�!,?���>�����ʾ&��3�˝?�Y?�;a����c<)�͑¾�Խ״>~[/�/~�Q���D�c������׀����?"��?�A��6��x�򾘿\���C?m!�>ZW�>��>��)�Q�g��$��/;>���>0R?���>�PO?�-{?�V[?�W>�&8���������_ ���#>�%@?m�?��?�x?�|�>�P>��(���߾%����$"������(��`�T=UZ>.!�>��>*��>W��=e�½:p����>���=#�b>2��>V�>���>^3x>T��<�G?���>�ܾ�u�*���>���*�=�Szu?v��?ː+?��='y���E�t��YP�>r^�?�?Q�)?�0T�n��=�Nټuȶ��r��C�>�ֹ>R��>��=�D=�Z>��>�k�>
s��_��w8���F��?	
F?<�=�ſf�q���p�s����'b<���)�d�����/@[�끤=�͘�����ʩ��[�������]
���Μ�I�{����>i��=�E�=��=�b�<��ʼ�=�<.�K=�e�<HX=�Ho�kyn<<�9��lѻ�*��:�"�J�Z<�dJ=I�껶�ɾ��{?V�I?��*?ǣD?�x>>��0�x�>�sw��?SC[>%�T�b!���;�祢�?���X�ؾ�3پx�f����>��C�&�>��1>�=p�G<�S�=�ex=E�=��g;�`/=@F�=س�=�.�=���=��>LP>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>"�1>	�>9�P���.�?}M�(�[�D�R��$?e.<��&ؾW�>s��=�Y�y-;m�=��5>�{w=h���\���= 쌽��V=��g=&s�>�fI>�ٯ=~ؽ�c�=&1g=҂�=�W>8����Ŝ�!`뼪:P=��=�d>�P+>O��>�?��0?��d?d�>��q��Ⱦ7�����>�N�=��>��O=�|3>a�>
�7?�@?֑F?k��>cN�=��>#�>9S+�Dl�!�b����
=|V�??|�?��>=&=xH,����'=��v���Z?O�0?X
?�y�>���P��6&�M(5�M����м�u=�$c��Xʻ��>;f��i�m}*>)ٿ>�+�>���>�j�>��_>�F>���>�>�����%V��o	��i�=���=i)��iG=U�=@�ż�P='�<G��=2A7�@�,=��[=��=If�>>7�=��>ŗb=ǃ��j�2>��=��|�%=��q��l�J�S�Uᗿ�>���s�d>�}|>qY(�����
��>�}�>gi�=��?:"|?z2u=MU��6P��k��0g]�y
ֽ�!!�*Y�>�U���5��oa�
L�-����-�>h��>��>��k>��'���8�t=���9 2��g�>����U�r�|��ui�U�������f����QnC?s���6k�=�?�N?���?C��>!v����ʾ�~&>&����=N������ɉ����?%%?��>Ѕ�k+F��̾~�����>�MH���O������X0�<.����?��>CΪ��Ѿ03��Z��(؏�l�B���r�º>��O?<�?�a�_T��	`O��|����]?hg?)o�>�y?�p?����b�I��+�=k�n?��?J�?��>�1�=o]�����>� 	?sɖ?��?Yr?��;�h��>�#�;�k%>�m���=�@>�Y�=2�=��?�V	?�?"���0
�ο�����GY��y�<c�=��>�e�>�or>�n�=~u=c��=�^>F-�>���>�we>
ߤ>"��>ء����O?�>1��>�.?s'F>�A>�rU�L����:jLz��G��d�W�����~i=ĉ�=f��=f�����>�cͿ.��?n��>d���9?����t5��z.�=%��>25)��N�>�U�>($�>�k�>��>2|4>g�=d/8>9.Ⱦ'�W>�O
���"�0�N��R�>	R�S܍>����f��4	��Fg�#Re��|���C�\!`�s����pC�Ф%=>g�?��I�A&e����q�K���?uW�>�%?ޕ-�b�+����>A�>Kk_>��վ�]������$>����?/��?�Mc>H"�>~�W?R�?=Z1�<3��Z���u�KA���d���`�!鍿\���$~
�����_?p�x?f]A?��<��y>w��?Z�%�Ώ�� �>�!/�u$;��==�C�>,���`��Ӿ��þ���_fF>��o?h�?|B?��V���c���ž�D<?@?��?���>��>W1>/3_?Uf�>v�?y|?��?�)"?ŒU?�'?���>g��<&������t���>(S���мj�=�е=��=���=�X;��='.�ŉ��7��=kS>
�>w,���wo=~�>>�	�=��>�]?�L�>}��>V�7?����o8�T���$/?�h9=L������Т�$��>��j?���?�VZ?}3d>;�A�&C��>RL�>}�&>F\>�[�>��@jE��=�r>@�>B�=��L�a�����	��l��	h�<$>+�>a}>�C��D�(>oɡ��v�vtb>��T�<˹�~;R�"�H���2�/]t����>5K?p?i��=�R�h֔��f��,(?P~<?$�M?�D?��=�ܾq 8�v6J����ݲ�>�<r
�9t���.����9����5p>�e���Ӡ��b>J���l޾?�n��J���� cM=���hT=R�4־���=�
>{���!����̪�a/J?�l=o��h}U��t��!�>w��>��>�;�#�v��l@����|"�=>|�>C}:>!̛��ﾰjG�]���>C?;_?_�?����Ir��XJ��u��ܤ�j�e��>?`�>C��>�9>�X�=���А���f�U�B���>a��>���A��j�� ����#�0>�>T�?��*>��?'Q?s?<jX?�w(?1��>щ�>�_{������A&?5��?��=��Խ�T�� 9�KF����>x�)?+�B�׹�>G�?߽?��&?�Q?޵?b�>� ��C@����>~Y�>��W��b��7�_>��J?Ӛ�>o=Y?�ԃ?��=>V�5��颾b֩�V�=�>��2? 6#?P�?���>��>e��1>��?_yx?�r?�`s?l�,>a#?�>QF?�<�>>m�>kj?�D?� p?��j?�6 ?P�?>��<W?}���&�"q��@��;j=�N�=�>(�2=d��=�k����=��=z4=��=��-=}>A;���e����>�>ݔ���y;>y	���F���T>�6?=�5��IA���]~���0=pه>*�>-��>,�;�4Z�<\a�>:�>�l�$�!?}�?:+?!�=��c�>��Y����u�>,?�V�=&$n��3����k��H��h?�9X?~�m����u�b?�B^?�����=��þ�B_�8��O?&.?�WE���>7�~?!r?JK�>|vg��n���T�`�r�e����=%��>zc��d�ז�>N�8?��>��_>0��=F۾@�w�ĥ����?#��?���?��?�P*>�n���߿Z�Ѿ���t T?@��>Ej��a[?�I���Ǿ�̾ꖾ�լ��������������a�� &��e*�+Ͻy��=�)?R?(�w?��^?���k���M������`� ��D��7N<�E�6���"�n�k�f�5������ʾ=%=�X|��xA���?\'?��/��r�>�R��W�rCо�>>֛����{��=G왽�-=b�Z=�b�=�,�;B���r ?v��>w.�>h�<?�\�J>� 1�C9�������4>ٽ�>�6�>s��>>��;M2.�����	�̾솾�ѽ��}>�`?6M?��Z?038�yz=��_���@��t�YT����=�|�����<�hF��P��\ ,�
�O��z����=���_"���{*?))�>$�u>��t?:l)?���,��x�ӽ!.$��Mo=`v|>vH?���>|~>���,�����>�l?V��>�Q�>#싾 V!��{���ʽ��>���>y��>}m>iD-���[�HJ���d���39�K��=�Xh?����`����>��Q?���:`><$f�>{[}��� �$�)�W�>3�?
��=�|:>��ľn���a{��	���Q)?E?{뒾��*���~>�f"?��>���>�5�?#��>�Oþ8�M9��?�^?�J?hA?4�>Ӡ =�����/Ƚ��&��,=ד�>][>*^l=��=&l�]�\������C=���=4�̼;���<Po����F<%��<��3>�5ʿ`�2�5aپ�0�'��E/<�/ę��S��D���5� � �޾[��݊h��A=2>��p�����a���� ��m��?D5@nWt�$
�����%!��>_��?�>�k���|���c�����?u�wMM�'�$<�DZ��%�g�^�;���&?Q����'ǿ]⡿9�߾s?��?�w?h��<�"���8���>,��<�ļ'
������ο
H��	2_?We�>ڶ�2a��n{�>��>�f>�fs>�������K��<�C?hq+?�= ?z�p��ʿ⻿c��<���?��@
~A?/�(����D�U=3��>D�	??�?>�Z1��C�����rJ�>J;�?���?ŵM=��W��
��ye?N�<q�F�s�ݻ��=W8�=�m=���J>~S�>�v��dA��Vܽ�4>�؅>�"���:u^��<N�]>R�ս�E��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�}��=[��>c�>,������O��I��U��=F� �8�ĿH�"��N!��
;%����'i������'ͽ�W
��Ǜ��~�������=P�%>ouX>�q�>geG>��4>��\?��r?k�>��>	)�,_��Fž��4</<���S�Q5��-3��pܥ�����þ������e���žQ�<����=xFQ��T��� "�0�e�ڵF���,?j3>�*;pN����;>�˾HV��'$�UJ��qѾi82��|m���?�qF?,����/W�U�)U�跽��U?�Y����c�����=�<��݁�<P$�>���=��边�3��+Q��0?7p?>��1ꐾ�J*>P� ���=F�+?�I?!o7< ԩ>%�$?�V*�FW�F[>��2>Z�>*��>�	>+����ڽ��?��T?��mA���>w�����x�[�]=>>:6�h���[>yl�<�t��܂M�ڑ��׶<5�Z?�>�)1�3�<�G������<bs�=S"\?ʥ?�޿>OR?ʗA?Fq>x�����T�^�*�e8o���a?��?��>Jc����a!ȾL?Ħ�?��y>6M��p/���&"����c?��_?�u4?F���c�pჿF���T2?��x?,�$������ھ榵����>�� ?ք?�U����>��^?���� ���Ϳ��Χ�?Y@�@����!IG�<���[|?ݷ$?�jԾ���ϨS�����_Q��
?/�A�����	�@H��L%?�#f?�=�>)�h��G&�/>�������?��?�'ƾK���(n�U�w�I%�����}��=�A`�a;]�6}��GM���޾������22�9o>S�@���r2�>����!߿}�����rž�����E�>[�>�o>�ӑy���z��H���m�T�U�ZN�aN�>��>�������Q�{��r;��[��g�>���>^�S�(��˚��pu5<@�>���>O��>�)���彾
ř? a���?οm������X?Gh�?�n�?�q?C�9<p�v�o�{�1)��-G?��s?'Z?|f%��5]��7���j?�Q���V`�ђ4�qBE��/U>�$3?�;�>�-�U�|=�>��>��>/�X�Ŀ'ٶ��������?T��?�m���>w�?<v+?�g�G8���[��D�*���P��3A?�2>q���|�!�Y4=��ǒ��
?	z0?���/�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?i�>��?���=�j�>a[�=찾:/�3�#> ��=��H��?�M?�>��=C9�
/��[F�MXR����̩C� �>�b?#~L?�}b>!&��k�6��W!�ʽ�T1�Tq��}2A�;�2��B�24>xQ>>�>��E��Ӿi� ?�d׾Rh⿯N�����KBR?tU�=��>ܶ��`��Oڽ��;?U��>�7�t|���|���(ǽ,ץ?V�?P�?d;0.�1�`>¸�>}z�>b��E>��]�=�?>��Y?z-Z>?#��3͊�o]�>+d�?@G��?�E���?������}��QR���F�c">�B=?u��-6=>�L�>�>�r��>��ȴm�rA�>��?���?k�>Z?�S��0�k2�>a��>�*?	�I?��=����8>�$?"�ɾ������udy?��@~"@"�?���A�ܿl���������㾃L�=Ϲ=��>C1�N��=Ȑ`=�,��o�Z���W>��>C"�>Zn>`�m>�&>�Z���������`^�:�!�!�H�����[�����������1׾�������z?�J�½A�Q�{T�������1>�oD?��f?�b?��?�5�=-�=)羱q_>��]�n鼔\�>��
?��9?G�?.>�b'��k��d�}��(觾{�>�� >�X�>xͪ>�p�>� �#�>�Ԁ>��>���>������=�6>F��>#��>��?t�h>}:<>�>ʹ�X1��"�h�b.w��,̽m��?������J��0��A;������?�=t_.?�n>a��>п����M4H?�ꔾt)�J�+���>��0?�dW?��>9����T�m6>���j� T>{X ��l��)�q$Q>�p?��q>-�~>��0���3�#M�ϫ��)�>}+9?@����Q��x��I���Ծ�wM>o�>uϿ���F��x�x�P
m�[�v=�H??��?�ޡ�����l=���E��*�_>eH>I�<�=	%5>J�h���ؽ*�:��9A=���=�P>�P?��+>��=�ߣ>�C��XP��d�>jyB>��+>��??z%?�p�z���U���].�?w>"P�>-�>�G>O!J�,*�=��>�a>�E��&���(@�;W>�$}��_�]�u���w=|җ����=ry�=� ��=�@�%=!�~?Z��+䈿g��c��2mD?}+?���=ŬF<F�"�< ��H��P�?e�@�l�?��	��V�i�?A�??��v��=�|�>J׫>[ξ��L�±?��Ž�Ǣ�ڔ	��)#�SS�?��?�/�)ʋ��l��5>�^%?�Ӿq6�>�ֺ=���T���l߄�d�=���>�&?'�ɾ�Q������>�~?@��g��:п:|v�F!�>ؖ�?��?�+D�)߮�6�`��?��?B�)?���nv&�&�����=�:?TU^?��>\^*��7<��2-?�?`��?��^>�B�? ~?Ͽv>������&�.Ɀ�������k���I>r8B�TA����6����؉�峌�y&R�O�K>�3�<#ֻ>��<
����~�=��.;=���b?���>�>[�e>���=L�=�~�>:k�>j��>���="��~:�'����K?b��?s��Nn��Q�<���=0x^��1?�54?ڍ`�S�Ͼ"��>D�\? ��?��Z?�I�>{��(<���ؿ�$���S_�<�3L>�G�>�E�>{����K>��Ծ��C�SQ�>ϗ>󯤼�Pھ6"��||���P�><e!?�u�>�a�=%'?%+?��u>k�>}�i��i��|\X�BYN?�>�V�>G	�?8˝>n0����#���~�����0h�-�v>L�n?�i&?r��>�y��
#��z0g��M��G�>��J?�1�?���>���>֎?�{?BB?���=�,���u�DBb>[C�>}�!?s���A��H&����z?�L?���>�1���ֽ<׼���C��&�?$\?3=&?՝��-a���¾��<r#���R��f�;��D�)�>.�>����	��=�>˰=\Nm�%E6�#�f<!m�=���>Y�=�27�z��h�3?��<=��Ծ&M>�b���[�P)�>ʊ>σ!�]�p?�ܼP*����򤳿�-���a�?�;�?� ?����Z�u�"�?C��?(�?e$?K�����Ѿey��U�x2|��W��;��5�?���=�L#���������,�����r4��?%��>��?�J�>bʲ=���>ʹ����
�&�.��M�s_o������+�� 8����-	���E�������Ⱦ�H�����>O+��d�>��>�o�=�9>�J ?�>�\�>9��>�e�=!��>)�>a��>���>N���v�m��^?�@��>�W��TR�^?��r?y�?�]ǽ�fT�r�4�R?U��?�?�O>��s��=�>��>�@?�R~���w>͍h>�6�>Ɍ�x�	�V<���>����C�9"�<F�}6Y�����j�.?�?�H�B�-�LؾԨy�R|�=�?-�(?B�)��^������A���a��_�\!��p��rP6��3g��ϐ�|��V����5�� +=�?v�?_��&@�	C����`���8�{J�>� ?�ve>�$�>M/>��Ⱦ�;��gE�@3��{�����>@P|?H��>W>?��G?�bM?�UO?��f>��>ξ���?�;��>D�?e�,?��-?=*0?��?~�$?�).>���'����꾀�?T�?�?d� ?4��>򈂾���"Y=]�˼��k���<Ca�=|�=����7��Y�=:]Y>9�1?�#>�N�p�G��[>'�?MR?b�>�a�;��Qp�f��>w�B?�_�>*'�@�������?wC�?����`U=ޟ�=F*>x�J>D7�=S%>����I�^�(�����E=�=X>c_�=�k{=)�>J�˼��ȼ���=�d�>}�?���>BC�>�0��� �ٮ�	��=��X>��R>@2>�8پ�����%��*�g�hy>�u�?�q�?�if=�E�=Q��=We���R������콾sR�<1�?�<#? UT?ȗ�?��=?VW#?)�>���H��;X��A����?W�,?���>Y7���ǾĚ��!�1�%?��?ya�YL�{�*���ľ�jƽ��>�-�Q{}������)D��o)�w��ʙ���#�?�?�����7��n�"瘿褣�9??ذ�>!��>���>�k(�Ki�����<>Z �>'�O?�>�HO?�t{?�[?�V>�<8�]ƭ�A��������!>�??<ف?ˋ�?��x?K��>�k>/(�A�~,����"�����(���Z=�<[>Ò>���>op�>�z�==½���?�>�B�=�b>�q�>0ۥ>�+�>�w>��<o�G?(��>�]������뤾�Ń��=��u?���?q�+?T=��/�E��G���I�>Uo�?���?�3*?ɼS����=��ּ�ᶾ�q�L%�>�ڹ>�1�>.ȓ=>zF=�b>��>[��>�)��`�Qq8��NM���?�F?'��=ƿ�q���p��З���c<����;Le�"�����Z�Ƥ=������ꭩ���[�dx���Z���ᵾ֤����{����>�Ɔ=N{�=���=���<��ʼ�V�<
�K=��<��=�*p��)n<�8��!ѻ����u'��"Z<pmI=���<�ɾ��|?ЮI?wr+?qC?�ft>�'>�8�Z�>x���?�U>y�`��#���+<�B֧�ve���7ھ5ؾ�
d�ު����>�nI�w>�3>D��=*��<��=�`z=���=f߹u=�'�=��=���=)��=�>W�>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>r��=w�2�T��>��J>���K��B����4�?��@��??�ዿТϿ6a/>s7>�V>�mR�7%1��v[�"wb���Y���!?�R;�!�̾!8�>��=,�߾�\Ǿ�&=1�6>��e=_��=\�	˙=�d���B==ݟg=�L�>R�C>d�=�D���Ʒ=,�J=��=��Q>�h»-4���#���5=
��=�c>n'>��>��?�c0?�Wd?:�>�n�vϾ�9���O�>��=8�>_ׅ=!sB>`��>��7?�D?k�K?Zr�>���=8 �>��>��,��m�i徿ʧ�D$�<��?n̆?�Ը>*iU<nMA�����^>��"Ž�v?jU1?�l?�ڞ>C�^+ٿ�o�.����+=Σ����g��v����K>F�>�z.�'���2x>졽>ё�>^�>On>���=O�û���>I>�-�;g��;+\$�YΪ�v'�$�����G�%W>��N���ԼEl�={���%=����^�ܻ˼���<[�=��>�B�=S��>{P=���fJ�>Rg�_e��V=��!�Y��\�ו��UK�9���,�>��?>�8?�)�����>݂�>�O�=�"�?$*�?}��=�#�'�{��Q��5/��"����A�XR�>�f���^9�gk���]�9z��"T�>Fя>�%�>X�m>O!+���>��=s=�-�*�4����>�뎾��(�w	��fp�X���L�����h� ]���rD?���zb�=|u~?�I?ڨ�?)[�>🞽Y�ھ��3>灾���<(�g=t�]����?0�&?	��>>f�mD��J˾�1���^�>d�F���O�0Օ��1�w��c"��pد>�����Ѿ:3��/��}����B�(�t���>�WO?�֮?X`��D���$O����������?W�g?'r�>��?�?�ɞ�ޖ�S����=�rm?�_�?`a�?�&>��=�����>�G?���?�Ύ?X�g?��8�w�>�s�=�$�>�8���>cP<>^H>:,>��
?��?t��>"������D��پ�D^���<�cM>�Y�>�Gx>�0~>j�D>O'�=V/<>xٓ>/�>LԶ>�P�>�I�>�Iy>	�����e0?38�=\��>�!&?#wh>�$>m�8�&h��=E:�p8���vq�}zS�#��=Ϲ�=p�=� ?���>�vɿ�? �$>�����?��<���y�=��>��<�m�>���=t�>&�>A�M>���=�>6�q>�/���<�>�
�["4�.`�Du�2Ӿ�em>����%������hq�C���ys�y�����f�+����F�Ǳ�<�z�?�"=mBq�)|8�5EK���,?���>�?� [��%�����=%<�>I��>��)ǫ��䕿�����?��?�Bc>��>��W?8�?��1�M3�PtZ�:�u�[$A��e���`�v፿����n�
���0�_?�x?wqA?Y��</z>���?�%��͏��)�>�/��';�W�;=�2�>�$����`�+�Ӿ��þ�;��<F>��o?$�?mT?�SV�S;�=��$�@?�W?���?�'?��?�q����K?y�%?h?�_?�+?�[H?čO?Ns ?��>ζ�:�ߊ��=��kf�Ԋ��2缠H�<Ӌ�=� =����9w5�m��=��#=��!�_{��({0����;��<��<�!�=�K�<���>ߡ]?�T�>��>��7?g���r8��Ů�B*/?x:9=����
���ʢ�	�4�>�j?���?VZ?�Rd>��A��C��'>�R�>Lu&>�\>�X�>A��	{E�M�=�V>�l>䫥=Z6M�򿁾�	����9�<�!>��?U�>��g���D>����_�z��lp>�B���d��W,��<iV��j7�Q�6�M�>:�;?rf?�e������!⼮*^�\�!?�>X?ǠO?��?z�Ѽ1��
�R�V���f��HZ>�&U���!�[���3s��\�#�4�=�+>蠗��e��)s�>�4�G?���)�u����0� >���
<}>���9� ���˾�=y݈> f�����)̏�Rծ�4�R?L���a޾����	v�,]�>��>.��>!֥�ܞ��}�R��ڈ�Z�>F�>tG=��̽ҿӾ��R����DU�>NkE?�x_?Oc�?ơ��Ss�RC����̃��Ufż�?�X�>�{?fB>�}�=�����nfd���F����>'K�>���l�G�|&������$�"��>�@?b�>��?�_R?��
?�p`?A�)?$7?�Ӑ>?�������<&? ��?ʀ�=3�ӽ<`U�^(9��F��3�>��)?S�B���>�?ҹ?Q�&?�[Q?�?$#>o ��@����>�>��W��O��.�`>�J?��>5;Y?%Ń?#�=>TE5��x�����f�=M�>��2?�#?Hz?��>��>���<�=��>�
c?s0�?��o?a��=�?U32>���>_��=��>Q��>~?XO?�s?��J?Ȑ�>�<m4���6��^?s�x�O��ł;��H<˿y=����'t�^S�n��<H>�;�`��KT��!�񼩹D�2��0��;B�>y>���k�4>�gþ(����6>�}��2u��j͊�g�&�0��=^b�>e�?En�>h�(�W6�=}�>���>D�(?E�?��?�!�ܬc���߾WW���>�QA?���=��h�����,v���M=�l?�Z\?btL�o���a?J�N?}!��7��5����;�F�߾�V?b�?G,��
�> �?�m?��>Fi����w�\���s�G�=��uC�=kI{>G���`�]V�>�}1?ݥ>�͏>�D�����J�N���S���?oЖ?���?t��?Z>{3^��ҿ����D��Aw^?R��>�>��J�"?E�̻�aѾ�8���Ɏ��?侮L��^ʬ��C���a��f]$�"҄�~�۽�<�=��?,r?Z�p?,�_?�+�,d��r]�_��W�T�U������E��TE��IC���n������������K=Y�w��@���?"�+?��$�F��>���NK���!ʾ~>>N����
�s�j=�M�����<W�L=��x��D>�e����`?ﴲ>eF�>7U<?��]�C�@�'�,�}�6�9���.>���>�>��>g
�GeE�3q��[;���󽽏Qv>�c?F�K?7�n?j3�d1�4����^!�),�';���JC>*�>���>�&W�S���Q&� _>���r�*��29��W�	� �|=�2?+L�>xϜ>�R�?=?�C	��?��ӷw��1���~<�w�>i?���>�؆>�kн� ����>��o?�i�>ל�>����p0�%
���O����>Q�>m�?⯢>�4�={P�z�S����;�|".>�]?rň��L��>;�D?����Ͻ�|�>�4��"����K=D��m>"<?�:�=���=�iʾ����Fg�Il���,?VA?��f�d ��2>2?9E?�=�>���?��=N.���G����?N�e?d�W?e=8?�]�>K��=���VBֽSpܽ�~�=IÌ>G� >�g=3W >�M���%�����RqD�JED=�{'=�Bm���Ҽ3�=M{�=`hN��1�=��ֿ��<����u���{̾���IE��;a�'vZ�d�\L���Ź�"���]@1�Re�<�q�����yc������?U�?߱��D����x���%{���ܿ�>��-�u-�=~1t��2��n���*ݾ��<�¨�VQB��Kc��H`��%?��˾awο����	_>_\?�Ĵ>Г>?��]J���:�֎8>D��=�z��龋ۉ�I����쾓b?/:�>�����=Yq?bʥ>.YV�f�>��^�9��������/?�]7?[��>�ʕ�����U��'2w����?�4@tcA?e�(���P=i��>>	
?"�>>��1�Q��5���V,�>���?ߊ?�mK=�W��	��2e?ٯ;o�F�OZ»��=�~�=�#=�^���J>���>D���BA���ܽͣ5>�F�>@�!�"����_��b�<G�\>jBӽ�[���Ԅ?�v\��f�ٟ/�)U���U>��T?K-�>0�=p�,?�2H��}ϿI�\��-a?Q0�?8��?��(?4࿾DϚ>�ܾj�M?PC6?���>.c&���t��g�=~��R
��k���$V����=O��>��>�,�`���O�P��}��=Ɏ��F^��w.��n$����=�=����3�������������-�d�ǽYK�<�U�=T|>]�>�^p>�\7>2�_?��?Q��>a=Nt�ٻ��AA��Y�%��&�?���Y�V��Ĉ̾��	��d��G��������gǾ��<��v0>u�R��T��bV�j A���k�+�?�K7>�J���G4���ؽdq�#Ϧ�^�(>EK�ht��)"�dk����?V`C?��|���Z�6���9=�$V��\?�C��0־n������=g����p�=UЈ>/�&�)�پ��/��G��3?�M?៰�"o���+>��5���0��'??w�?�Y��>�>T6?�J��� <��>���<� m>���>i�>�����,9���)?e+j?��5�<۾jR>[@����h���<լ.>�q�g1���dI>��3>�D��1�=s
y��hƽ.wW?�$�>P�'�������+�%�yώ=��}?�?�Ń>�m?�:?��H<#�ᾡoF�7���;�<R�W?�lb?�>�$���}Ӿ�β��j1?e�h?�~�>�P����T:�/��D�?��k?֨?6�=�x��ꐿg���7/?L�n?�n<��Α��5۾"ł�hy�>pc ?w5�>WOG�!-�>��?�!��6����º��I�[�?��@B��?�5�==Ѿ� �
>3?1��>����쾖�V�� ��X�=*p1?0t����мB�/弾&`/?�S�?�.?��b��I����=aו��[�?T�?������a<����(l��;�����<��=G���#����,�7�g�ƾ��
�趜�n�����>`I@��*�>�9�~3⿪;Ͽ����о0'q�d�?k�>�]ɽt���x�j��Ou�`�G�>�H�_x��v�>ìV>��<�lA���g��lH��$a���?�l@>sS>#�=5i��Z����0>�,�>t�>hQ�==�=v����8�?���ؿ�ͣ��M���d?/�?� �?W��>:�c�L�=�wl�r���:?uw�?�uN?ܐѽǓ]�Ĳ���i?�U����_���"���,�T��>�a*?��>!�;��Z;���>��>6(�=�W0���ÿ�_��|:㾾ߩ?͡�?�}�C�	?�̛?�? ?{j:��F��2L�o:1��h<�M?Mf>�<��D�3�VRJ�;���"�/??[c?�9����2�\�_?&�a�M�p���-�w�ƽ�ۡ>��0��e\��M��'���Xe����@y����?K^�?d�?��� #�a6%?�>h����8Ǿ��<���>�(�>&*N>^H_���u>����:��h	>���?�~�?Sj?���������U>�}?�5�>}��?^D">�v? xt=���y,���i>�yM>�Щ��!?&�d?���>,>XG����5�#�6�2},�����C���>��y?b2P?~�e=6nj�5[/��3-��o�� ��x������*�p��fw�S��<.�=̫=h�&�N@ɾm�$?��%��Sҿ�K���;=i�9?(�?>+�?9��;＾.?߼�lZ?S��>���I�������x��`V�?!�?"��>�P����=�oc>�fE=�A>?��<ߦ��cz�V��=�o9?��ӽ�*��Ƒc��	�=�t�?�@��?�YT�|	?E��~����|�&����2�4,�=927?(����s>j��>0�=�1v��y��Y�t���>�5�?�v�?���>v�j?�l��F@���+=cW�>��h?�h?*K��!��O>��?X�߉���	�ge?�@3�@a�]?�����Yؿ8���Ԝ��B���>&��=(�_>�q����=�}�=��R=a4e;)$;>��>::K>/�e>��>M@>9� >-���%�%��뤿�i���==�x�����]����Ɋ��RܾC�ؽ2�~�b\Լ��B�-۽.��:�ҙ#���=}q?��U?�~y?04�>��<��f>bD澲��𸁾�{�= N�=�2?:j?p�:?:�>r⍾�l�ZV�������[���>h7>���>��>E��>�S����->Tǫ=��=��d>��x�/┽�d�<է{=���>��>��>x:>@^=>ް��g�����!�V۲<�ւ�yE�?@�|��� �����2��𓦾�iR=��%?��='Lr��Nٿ�����L?A־�-�X��;�c>k�<?��_?�Y"��2��N�|=�[=+���	n��J<�V������f�+�N=�.?q�f>�ru>�3��v8�gP�Qx��A�{>@6?���8��u���H�<�ܾƫM>��>Ɋ:��%����&B���h��x= 3:?�?iP���9����t�͞�%�R>Y�\>��=	0�=��M>�e���ȽTG�ۧ.=z�=��_>`-?0?>���=%6�>�>��y�n�ɓ>ukF>�>>l>?l)?;e�;��u���{�f!�d�[>eq�>��>t��=�W���=��>�KY>�u��s����{�L�
�[>�oq��`u���.��=�7Ƚx��=a�F=/t��\�M�0=�~?���(䈿��e���lD?S+?a �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��L��=}�>	׫>�ξ�L��?��Ž5Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>x�mZ��p��+�u���#=��>�8H?V����O��>�w
?�?�^�ݩ����ȿW|v����>]�?���?"�m�sA���@�Z��>)��?agY?�oi>�g۾`Z����>�@?�R?p�>�9�A�'�j�?�޶?���?��O>c��?��y?�+�>!y��'�>����R��CN�=�w���>�K]>�ힾH�:�����0荿��k��P���^>џ=1�>N����ϴ�a�=H஽�\��NB��K�>�>a>��7>��>u��>���>�sx>��=vd��w/i��끾�dG?�?^9Ѿ!�1�ʿ7����=��=�?��?*��9�S�z�!Ep?η�?Xu?��?�(�!뗿L���u�¾]��=	��=��?���>�)s����|%��H�>ޟ>C��&y��Ś�;��l����>��+?b1>5���Y| ?T�?�̺>D��>�U��9��{$�SP�>��*?g1�>�Ui?��>����h%�^������©N�ۢ�>N�o??_at>#��˨��>w��>D� �/��?�[?}�Z�j�9?��?�q?]o?�)�>a&�ʁپ㥿����>�'?Q��6#�o��`�A��� ?f�(?�W?BJ�=�����=�4&�����m� ?
�p?TZ? ���7��`��/�#;َ7=��`=`&0=�����*'>�;]>+�罋b>�p">���<s���GnP��'j=K��=�]�>T,>fz�2�~K'?,�I��^(�7>�fg�O�3��f�>�?�W����U?Ab����n��G���}��컬�m�?p��?v��?�|%=�G^�1�?�׏?1�5?>V�>6о0c��r���֐f�e.���"����>�T�>��;�p����|�������R��h�ʏ̽� �>�>?Ӹ/?���>�>���>j����1������D�DX�T��ׁN���,�s�������O����J=��ɾDڅ��R�>ƈ����>�^?�	>�4>2��>7ƃ<6j>�(�=p�,>��>U�>���=Β���r���'�A�R?z���7��@澭�9?O5l?@M	?ΖK��d��.�޾�}?Qw�?�~�?GΟ>�v_���4���?�u�>��w��?yo�=�-�4���V蛾�����c��ׂ��T*c>J���9�1�3�%!J��?c�?�eP;��ʾMU����`��듼B��?P�U?C�2���Z��.)�,怿)��29��y�i�<�J��s}������v�=J� �R�=RU%?b�?c,ھ�VȾ��H�Q�,���>�
?��> �9?Q== �#������W�y�3�����r
?�XX?���>�I?U�;?Q�P?��K?�ǎ>�t�>^対t��>�R�;T9�>��>6�9?7.?fX0?��?�J+?:�a>S:���4���ؾ�"? �?.?~?��?4O��deĽk��f0}�X�x��Q��}F�=u�<��ٽ��v��.V=�tT>SW?��Up5�@�����f>�3?��>���>�T���젾@h=M�>��?�Ƙ>����o�&0����>Q�~?3a�s&=��;>e�=K��'E�<JZ>����v٪=��n���)�t��*l�=��=]f�<�ʍ<(�6<ٌ/<�4�<�s�>x�?Ҩ�>�Y�>EZ��� �_�����=�Y>�S>f�>�Dپۂ���%��R�g�?7y>ur�?~u�?�g=.�=���=a���e`��K��/����<�?nL#?�JT?���?��=?�h#?��>�%��N��cZ��������?J,?��>����ɾ�٨���3��?�U?�`�X)���(��h��˽ӽ@�>�/��)~��寿6�C�۷��*���
��X��?���?W�F�z�6�ݳ�}���9� pC?W�>��>7&�>��)��,h��5��(:>��>��Q?��>�V?��?�%Y?O��=p=Q��n��ϫ��x��=Z8>�DC?.�? �?2$q?��>`'=K�`����
�ܾ��u��������vb=e�b>> �>���>I��>@�>Sҥ��=��퀾��=U��>���>b��>R��>�JU>�E=��G?i��>�i������ޤ������7=���u?���?e�+?��=8��R�E�zD���H�>�l�?^��?e'*?&�S����=�r׼$඾�q�x,�>�ܹ>�7�>��=��F=�d>��>���>��Fb��s8�EM�u�?nF?��=VVſ��p��:m��p���y<7����d�����Z�dv�=(����N�˔��(^�e�����)����e���~{��U�>�K�=�v�=���=�K�<؞μNڵ<�1J=[��<�=݇k��.o<��D�&.ǻ�7��G����v4<��D=1����[ʾ��{?�I?�,,?{lC?�Ay>W>[|O���>ހ�W?V>�ST��<���=��ɧ�,j��&qپ��վ�d�%��҈>"GK��>D�3>b��=N�v<�R�=� t=Ex�=�ʻ
�	=�C�=��=߫=��=x�>k�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�C6>A�>��R��2�إ[��Ba�ڹ]�!�!?��:��{ʾ	��>BǶ=�߾@ƾH�:=�"6>�,d=��!c\��=4Px�[s4=��`=�߉>�F>fɺ=	���Ρ�=]YD=�\�=]�N>��}�^4�?r/��\,=��=g�`>�2$>D��>��?1e0?Xd?��>Bn�$.ϾP-��,[�>}+�=�W�>�K�=�~B>���>��7?��D?K�K?`��>F��=���>{	�>��,�Y�m�/j徴ǧ����<U��?�ˆ?˸>r�P<��A�{���c>�TdŽ�q?dH1?'k?�ߞ>@
�Q����0���=���=�Q0>�}�����J�=�c���2>��>���>[%T>�\�>�b
?HP>�ץ<�۷>FJ->�+�;el(���=k=���V�=�j=�=!=��]����D�{��7����;X��=$tg=CA�=ڋ��\>7N�>�\>���>�IE= U¾�\>�Ȼ�ҜT�ߧ=�u;BM#��_�y����-4��?�x�D>�0/>�W;ד����>Z��>�:U>���?�i?39>�(��p���/�����s��޾���i>��d>u���uJ�}r��X� �̾��>e��>�7�>oEm>��+� ?�y=[;⾯n5����>ں�����)��Iq��8��y柿�h����S�D?�A��~X�=�~?��I?��?���>�E���uؾ2W0>�:����=����zp��⑽e�?��&?9�>�(�[�D�aȾ�۸�<�>��7��{R�1Ö�h�-�k�ż,F��[а>�i���=Ѿ��6�顆�����C.C��ir��a�>��N?��?�7T�0H��K�P��� ���%��>��j?���>��?�
?�����8�iu�ϟ�=�Qi?���?M�?K
>G��=8���Q�>�2	?ƺ�?���?s?N�?��a�>���;�N >����U�=Ԋ>=E�=]�=c?��
?��
?�|����	�8����E^��q�<�ɡ=t�>���>-�r>���=�1g=��=~0\>Z��>�ݏ>չd>f��>�C�>@���z�w�&?@w�=���>RB2?@`�>-aV=��e��<��N�i/?��J+��︽�Ͼ<����L=/�μ��>b�ǿ��?'BT>_��}�?���ώ2�hT>�CU>��ݽ���>�AE>�|>���>���>J�>{O�>̟(>��ɾ�0>���5�$���5�nA��]վ/�f>�#����&	����Ї=�wu��jA��Ed�ù}��F��� <77�?���nf�[���?��ml?1�>��/?�����晽ߞ&>4��>�7�>Ϧ �C�������W�徟��??��?<c>��>��W?��?Õ1��3�auZ�`�u��'A��e���`�[፿S���Q�
����C�_?y�x?�xA?{Y�<;z>M��?�%�rԏ�))�>/�.';�|P<=/,�>�)��0�`�ӯӾ��þ�5��GF>��o?%�?�Y?�SV�q�m�j'>8�:?H�1?9Lt?��1?X�;?p����$?j3>K7?�n?�G5?��.?Z�
?�2>���=!V����'=YB����>�ѽBuʽ���3=nN{='^
�t�<��=��<���Pڼr�;����4�<S�9=�ݢ=]�=���>�]?�P�>���>��7?C���y8�Qî�+/?}�9=�������YĢ�?�2�>��j?���?�cZ?1\d>U�A�� C��/>/U�>_&>��[>�]�>ɏ��E���=S7>m_>9ӥ=ΚM�'ہ�(�	�����#G�<�'>2q�>���>��9����>�V־�. �]F�>�
�_r�&^_�pb�%�T��B`�	�?��[?��9?���=�����k�R�g�80(?Mr=?��D?#:j?ٌ�=D��ԜN��=S��2�|�
>c��=�0�.����˓��=H�/L<�n�|>6���e��)s�>�4�G?���)�u����0� >���
<}>���9� ���˾�=y݈> f�����)̏�Rծ�4�R?L���a޾����	v�,]�>��>.��>!֥�ܞ��}�R��ڈ�Z�>F�>tG=��̽ҿӾ��R����DU�>NkE?�x_?Oc�?ơ��Ss�RC����̃��Ufż�?�X�>�{?fB>�}�=�����nfd���F����>'K�>���l�G�|&������$�"��>�@?b�>��?�_R?��
?�p`?A�)?$7?�Ӑ>?�������<&? ��?ʀ�=3�ӽ<`U�^(9��F��3�>��)?S�B���>�?ҹ?Q�&?�[Q?�?$#>o ��@����>�>��W��O��.�`>�J?��>5;Y?%Ń?#�=>TE5��x�����f�=M�>��2?�#?Hz?��>��>���<�=��>�
c?s0�?��o?a��=�?U32>���>_��=��>Q��>~?XO?�s?��J?Ȑ�>�<m4���6��^?s�x�O��ł;��H<˿y=����'t�^S�n��<H>�;�`��KT��!�񼩹D�2��0��;B�>y>���k�4>�gþ(����6>�}��2u��j͊�g�&�0��=^b�>e�?En�>h�(�W6�=}�>���>D�(?E�?��?�!�ܬc���߾WW���>�QA?���=��h�����,v���M=�l?�Z\?btL�o���a?J�N?}!��7��5����;�F�߾�V?b�?G,��
�> �?�m?��>Fi����w�\���s�G�=��uC�=kI{>G���`�]V�>�}1?ݥ>�͏>�D�����J�N���S���?oЖ?���?t��?Z>{3^��ҿ����D��Aw^?R��>�>��J�"?E�̻�aѾ�8���Ɏ��?侮L��^ʬ��C���a��f]$�"҄�~�۽�<�=��?,r?Z�p?,�_?�+�,d��r]�_��W�T�U������E��TE��IC���n������������K=Y�w��@���?"�+?��$�F��>���NK���!ʾ~>>N����
�s�j=�M�����<W�L=��x��D>�e����`?ﴲ>eF�>7U<?��]�C�@�'�,�}�6�9���.>���>�>��>g
�GeE�3q��[;���󽽏Qv>�c?F�K?7�n?j3�d1�4����^!�),�';���JC>*�>���>�&W�S���Q&� _>���r�*��29��W�	� �|=�2?+L�>xϜ>�R�?=?�C	��?��ӷw��1���~<�w�>i?���>�؆>�kн� ����>��o?�i�>ל�>����p0�%
���O����>Q�>m�?⯢>�4�={P�z�S����;�|".>�]?rň��L��>;�D?����Ͻ�|�>�4��"����K=D��m>"<?�:�=���=�iʾ����Fg�Il���,?VA?��f�d ��2>2?9E?�=�>���?��=N.���G����?N�e?d�W?e=8?�]�>K��=���VBֽSpܽ�~�=IÌ>G� >�g=3W >�M���%�����RqD�JED=�{'=�Bm���Ҽ3�=M{�=`hN��1�=��ֿ��<����u���{̾���IE��;a�'vZ�d�\L���Ź�"���]@1�Re�<�q�����yc������?U�?߱��D����x���%{���ܿ�>��-�u-�=~1t��2��n���*ݾ��<�¨�VQB��Kc��H`��%?��˾awο����	_>_\?�Ĵ>Г>?��]J���:�֎8>D��=�z��龋ۉ�I����쾓b?/:�>�����=Yq?bʥ>.YV�f�>��^�9��������/?�]7?[��>�ʕ�����U��'2w����?�4@tcA?e�(���P=i��>>	
?"�>>��1�Q��5���V,�>���?ߊ?�mK=�W��	��2e?ٯ;o�F�OZ»��=�~�=�#=�^���J>���>D���BA���ܽͣ5>�F�>@�!�"����_��b�<G�\>jBӽ�[���Ԅ?�v\��f�ٟ/�)U���U>��T?K-�>0�=p�,?�2H��}ϿI�\��-a?Q0�?8��?��(?4࿾DϚ>�ܾj�M?PC6?���>.c&���t��g�=~��R
��k���$V����=O��>��>�,�`���O�P��}��=Ɏ��F^��w.��n$����=�=����3�������������-�d�ǽYK�<�U�=T|>]�>�^p>�\7>2�_?��?Q��>a=Nt�ٻ��AA��Y�%��&�?���Y�V��Ĉ̾��	��d��G��������gǾ��<��v0>u�R��T��bV�j A���k�+�?�K7>�J���G4���ؽdq�#Ϧ�^�(>EK�ht��)"�dk����?V`C?��|���Z�6���9=�$V��\?�C��0־n������=g����p�=UЈ>/�&�)�پ��/��G��3?�M?៰�"o���+>��5���0��'??w�?�Y��>�>T6?�J��� <��>���<� m>���>i�>�����,9���)?e+j?��5�<۾jR>[@����h���<լ.>�q�g1���dI>��3>�D��1�=s
y��hƽ.wW?�$�>P�'�������+�%�yώ=��}?�?�Ń>�m?�:?��H<#�ᾡoF�7���;�<R�W?�lb?�>�$���}Ӿ�β��j1?e�h?�~�>�P����T:�/��D�?��k?֨?6�=�x��ꐿg���7/?L�n?�n<��Α��5۾"ł�hy�>pc ?w5�>WOG�!-�>��?�!��6����º��I�[�?��@B��?�5�==Ѿ� �
>3?1��>����쾖�V�� ��X�=*p1?0t����мB�/弾&`/?�S�?�.?��b��I����=aו��[�?T�?������a<����(l��;�����<��=G���#����,�7�g�ƾ��
�趜�n�����>`I@��*�>�9�~3⿪;Ͽ����о0'q�d�?k�>�]ɽt���x�j��Ou�`�G�>�H�_x��v�>ìV>��<�lA���g��lH��$a���?�l@>sS>#�=5i��Z����0>�,�>t�>hQ�==�=v����8�?���ؿ�ͣ��M���d?/�?� �?W��>:�c�L�=�wl�r���:?uw�?�uN?ܐѽǓ]�Ĳ���i?�U����_���"���,�T��>�a*?��>!�;��Z;���>��>6(�=�W0���ÿ�_��|:㾾ߩ?͡�?�}�C�	?�̛?�? ?{j:��F��2L�o:1��h<�M?Mf>�<��D�3�VRJ�;���"�/??[c?�9����2�\�_?&�a�M�p���-�w�ƽ�ۡ>��0��e\��M��'���Xe����@y����?K^�?d�?��� #�a6%?�>h����8Ǿ��<���>�(�>&*N>^H_���u>����:��h	>���?�~�?Sj?���������U>�}?�5�>}��?^D">�v? xt=���y,���i>�yM>�Щ��!?&�d?���>,>XG����5�#�6�2},�����C���>��y?b2P?~�e=6nj�5[/��3-��o�� ��x������*�p��fw�S��<.�=̫=h�&�N@ɾm�$?��%��Sҿ�K���;=i�9?(�?>+�?9��;＾.?߼�lZ?S��>���I�������x��`V�?!�?"��>�P����=�oc>�fE=�A>?��<ߦ��cz�V��=�o9?��ӽ�*��Ƒc��	�=�t�?�@��?�YT�|	?E��~����|�&����2�4,�=927?(����s>j��>0�=�1v��y��Y�t���>�5�?�v�?���>v�j?�l��F@���+=cW�>��h?�h?*K��!��O>��?X�߉���	�ge?�@3�@a�]?�����Yؿ8���Ԝ��B���>&��=(�_>�q����=�}�=��R=a4e;)$;>��>::K>/�e>��>M@>9� >-���%�%��뤿�i���==�x�����]����Ɋ��RܾC�ؽ2�~�b\Լ��B�-۽.��:�ҙ#���=}q?��U?�~y?04�>��<��f>bD澲��𸁾�{�= N�=�2?:j?p�:?:�>r⍾�l�ZV�������[���>h7>���>��>E��>�S����->Tǫ=��=��d>��x�/┽�d�<է{=���>��>��>x:>@^=>ް��g�����!�V۲<�ւ�yE�?@�|��� �����2��𓦾�iR=��%?��='Lr��Nٿ�����L?A־�-�X��;�c>k�<?��_?�Y"��2��N�|=�[=+���	n��J<�V������f�+�N=�.?q�f>�ru>�3��v8�gP�Qx��A�{>@6?���8��u���H�<�ܾƫM>��>Ɋ:��%����&B���h��x= 3:?�?iP���9����t�͞�%�R>Y�\>��=	0�=��M>�e���ȽTG�ۧ.=z�=��_>`-?0?>���=%6�>�>��y�n�ɓ>ukF>�>>l>?l)?;e�;��u���{�f!�d�[>eq�>��>t��=�W���=��>�KY>�u��s����{�L�
�[>�oq��`u���.��=�7Ƚx��=a�F=/t��\�M�0=�~?���(䈿��e���lD?S+?a �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��L��=}�>	׫>�ξ�L��?��Ž5Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>x�mZ��p��+�u���#=��>�8H?V����O��>�w
?�?�^�ݩ����ȿW|v����>]�?���?"�m�sA���@�Z��>)��?agY?�oi>�g۾`Z����>�@?�R?p�>�9�A�'�j�?�޶?���?��O>c��?��y?�+�>!y��'�>����R��CN�=�w���>�K]>�ힾH�:�����0荿��k��P���^>џ=1�>N����ϴ�a�=H஽�\��NB��K�>�>a>��7>��>u��>���>�sx>��=vd��w/i��끾�dG?�?^9Ѿ!�1�ʿ7����=��=�?��?*��9�S�z�!Ep?η�?Xu?��?�(�!뗿L���u�¾]��=	��=��?���>�)s����|%��H�>ޟ>C��&y��Ś�;��l����>��+?b1>5���Y| ?T�?�̺>D��>�U��9��{$�SP�>��*?g1�>�Ui?��>����h%�^������©N�ۢ�>N�o??_at>#��˨��>w��>D� �/��?�[?}�Z�j�9?��?�q?]o?�)�>a&�ʁپ㥿����>�'?Q��6#�o��`�A��� ?f�(?�W?BJ�=�����=�4&�����m� ?
�p?TZ? ���7��`��/�#;َ7=��`=`&0=�����*'>�;]>+�罋b>�p">���<s���GnP��'j=K��=�]�>T,>fz�2�~K'?,�I��^(�7>�fg�O�3��f�>�?�W����U?Ab����n��G���}��컬�m�?p��?v��?�|%=�G^�1�?�׏?1�5?>V�>6о0c��r���֐f�e.���"����>�T�>��;�p����|�������R��h�ʏ̽� �>�>?Ӹ/?���>�>���>j����1������D�DX�T��ׁN���,�s�������O����J=��ɾDڅ��R�>ƈ����>�^?�	>�4>2��>7ƃ<6j>�(�=p�,>��>U�>���=Β���r���'�A�R?z���7��@澭�9?O5l?@M	?ΖK��d��.�޾�}?Qw�?�~�?GΟ>�v_���4���?�u�>��w��?yo�=�-�4���V蛾�����c��ׂ��T*c>J���9�1�3�%!J��?c�?�eP;��ʾMU����`��듼B��?P�U?C�2���Z��.)�,怿)��29��y�i�<�J��s}������v�=J� �R�=RU%?b�?c,ھ�VȾ��H�Q�,���>�
?��> �9?Q== �#������W�y�3�����r
?�XX?���>�I?U�;?Q�P?��K?�ǎ>�t�>^対t��>�R�;T9�>��>6�9?7.?fX0?��?�J+?:�a>S:���4���ؾ�"? �?.?~?��?4O��deĽk��f0}�X�x��Q��}F�=u�<��ٽ��v��.V=�tT>SW?��Up5�@�����f>�3?��>���>�T���젾@h=M�>��?�Ƙ>����o�&0����>Q�~?3a�s&=��;>e�=K��'E�<JZ>����v٪=��n���)�t��*l�=��=]f�<�ʍ<(�6<ٌ/<�4�<�s�>x�?Ҩ�>�Y�>EZ��� �_�����=�Y>�S>f�>�Dپۂ���%��R�g�?7y>ur�?~u�?�g=.�=���=a���e`��K��/����<�?nL#?�JT?���?��=?�h#?��>�%��N��cZ��������?J,?��>����ɾ�٨���3��?�U?�`�X)���(��h��˽ӽ@�>�/��)~��寿6�C�۷��*���
��X��?���?W�F�z�6�ݳ�}���9� pC?W�>��>7&�>��)��,h��5��(:>��>��Q?��>�V?��?�%Y?O��=p=Q��n��ϫ��x��=Z8>�DC?.�? �?2$q?��>`'=K�`����
�ܾ��u��������vb=e�b>> �>���>I��>@�>Sҥ��=��퀾��=U��>���>b��>R��>�JU>�E=��G?i��>�i������ޤ������7=���u?���?e�+?��=8��R�E�zD���H�>�l�?^��?e'*?&�S����=�r׼$඾�q�x,�>�ܹ>�7�>��=��F=�d>��>���>��Fb��s8�EM�u�?nF?��=VVſ��p��:m��p���y<7����d�����Z�dv�=(����N�˔��(^�e�����)����e���~{��U�>�K�=�v�=���=�K�<؞μNڵ<�1J=[��<�=݇k��.o<��D�&.ǻ�7��G����v4<��D=1����[ʾ��{?�I?�,,?{lC?�Ay>W>[|O���>ހ�W?V>�ST��<���=��ɧ�,j��&qپ��վ�d�%��҈>"GK��>D�3>b��=N�v<�R�=� t=Ex�=�ʻ
�	=�C�=��=߫=��=x�>k�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�C6>A�>��R��2�إ[��Ba�ڹ]�!�!?��:��{ʾ	��>BǶ=�߾@ƾH�:=�"6>�,d=��!c\��=4Px�[s4=��`=�߉>�F>fɺ=	���Ρ�=]YD=�\�=]�N>��}�^4�?r/��\,=��=g�`>�2$>D��>��?1e0?Xd?��>Bn�$.ϾP-��,[�>}+�=�W�>�K�=�~B>���>��7?��D?K�K?`��>F��=���>{	�>��,�Y�m�/j徴ǧ����<U��?�ˆ?˸>r�P<��A�{���c>�TdŽ�q?dH1?'k?�ߞ>@
�Q����0���=���=�Q0>�}�����J�=�c���2>��>���>[%T>�\�>�b
?HP>�ץ<�۷>FJ->�+�;el(���=k=���V�=�j=�=!=��]����D�{��7����;X��=$tg=CA�=ڋ��\>7N�>�\>���>�IE= U¾�\>�Ȼ�ҜT�ߧ=�u;BM#��_�y����-4��?�x�D>�0/>�W;ד����>Z��>�:U>���?�i?39>�(��p���/�����s��޾���i>��d>u���uJ�}r��X� �̾��>e��>�7�>oEm>��+� ?�y=[;⾯n5����>ں�����)��Iq��8��y柿�h����S�D?�A��~X�=�~?��I?��?���>�E���uؾ2W0>�:����=����zp��⑽e�?��&?9�>�(�[�D�aȾ�۸�<�>��7��{R�1Ö�h�-�k�ż,F��[а>�i���=Ѿ��6�顆�����C.C��ir��a�>��N?��?�7T�0H��K�P��� ���%��>��j?���>��?�
?�����8�iu�ϟ�=�Qi?���?M�?K
>G��=8���Q�>�2	?ƺ�?���?s?N�?��a�>���;�N >����U�=Ԋ>=E�=]�=c?��
?��
?�|����	�8����E^��q�<�ɡ=t�>���>-�r>���=�1g=��=~0\>Z��>�ݏ>չd>f��>�C�>@���z�w�&?@w�=���>RB2?@`�>-aV=��e��<��N�i/?��J+��︽�Ͼ<����L=/�μ��>b�ǿ��?'BT>_��}�?���ώ2�hT>�CU>��ݽ���>�AE>�|>���>���>J�>{O�>̟(>��ɾ�0>���5�$���5�nA��]վ/�f>�#����&	����Ї=�wu��jA��Ed�ù}��F��� <77�?���nf�[���?��ml?1�>��/?�����晽ߞ&>4��>�7�>Ϧ �C�������W�徟��??��?<c>��>��W?��?Õ1��3�auZ�`�u��'A��e���`�[፿S���Q�
����C�_?y�x?�xA?{Y�<;z>M��?�%�rԏ�))�>/�.';�|P<=/,�>�)��0�`�ӯӾ��þ�5��GF>��o?%�?�Y?�SV�q�m�j'>8�:?H�1?9Lt?��1?X�;?p����$?j3>K7?�n?�G5?��.?Z�
?�2>���=!V����'=YB����>�ѽBuʽ���3=nN{='^
�t�<��=��<���Pڼr�;����4�<S�9=�ݢ=]�=���>�]?�P�>���>��7?C���y8�Qî�+/?}�9=�������YĢ�?�2�>��j?���?�cZ?1\d>U�A�� C��/>/U�>_&>��[>�]�>ɏ��E���=S7>m_>9ӥ=ΚM�'ہ�(�	�����#G�<�'>2q�>���>��9����>�V־�. �]F�>�
�_r�&^_�pb�%�T��B`�	�?��[?��9?���=�����k�R�g�80(?Mr=?��D?#:j?ٌ�=D��ԜN��=S��2�|�
>c��=�0�.����˓��=H�/L<�n�|>6��7������>;LD��;�Ω��C��g#
�(������A%�>".����F!����*=�L�=_�\�S�ҾUژ�Eg��;d?�bm�>�ؾ�0ｰ���.<V>kK�>�>u>���X�G���\�v�8>�>�U��R"����Ae��p�JI�>��D?��^?S��?�%���r�i�C������ǝ��*��Sh?�5�>��?�%A>���=w�����nd�lZF����>o��>'^��G��B����_$��F�>�s?I� >PN?BGR?�#?:n`?o4*?��?�А>�8�������&?u\�?�
�=_�2(N���8�V�I�>�>00?&�9��J�>U�?
O?1/$?3K?:�?�% >9���=����>���>&.U�eX��k>��J?��>,�U?>Ƃ?U�K>Ʌ6���� D#�Ë�=�(>�01?�l#?$?���>���>U틾�3�=&U�>�xa?�$�?'t?#�>T�>E��=@�>FɊ=�_�>�3 ?�'!?�`S?D{?�4J?���>av��z���k��r�8��]<ۋG��t<8�A=��;����M<��0=���;H��������� ��*̻��M�<�v�>F�q>-a���->�!ľ,%����H>%��95���*��/�\�=��>H�?���>Nl��p=��>�}�>����&?)w?}?	\�z`�ćپ�U�é�>RA?�Y�=�m��l��A�r���p=��o?O�]?q�b������Y`?�P?��ھ��8��bފ�����<?} ?T9�P2�>�8n?��a?���>��k�V@c�<N��^�\��fr��d�=ݶ�> Z��F`��>�:?���>�dF>�i(>䇻����E��H�1?Y��?��?⑇?�F>m�p�X�ҿ7��vq��"�^?���>�Ǩ�Y ?~�%��hҾ���=X��31�T������}{��x]��9t!��ˆ������=�8?��q?n"p?�D`?�c�c�(R\����� T�:�����F�d�B�o�B��m�k�������ꖾ��\=�q�BE>�!P�?y7??�g���>����ԍ�MV��Q�!>Ƹ� ���i��6��I	��N�=�ݕ���w�;���e?��>%S�>��B?��\��!<�"B��(D����AK>y�>�g>�|�>4޼(,Q���P���þ�x�K���v>�-c?�]K?�;n?�=��#1�����bq!��O%�e���Y�A>>��>O_W�����&�*3>��r����'?��`�	��}=ai2?tX�>?��>��?;�?(	�����(�x��)1�Vm�<�t�>�i?CL�>C�>+!ѽ5� ��>�l?�M�>�Q�>og���2�0���x�M��y�>"}�>>F?��v>Ǽ���Y�s���H��i�=��b>��]?����҂E��Wm>u�>?�d����=x��>�~ٻ���-�ླ{#��v�=���>�.@=�F�=��Ǿ)���z?h��W[��9,?��?xՂ��'���|>��?�g�>�d�>��?� �>ut��q�0=�n#?h�X?�Z??.�2?D��>�r����Žh'��=@��>��;>GV�=���=U��d� N齝�$>I�=�Y�;�%�1,	>�&=J�=�?=�.(>;��F�����[� ��n޾cw�K���(UW��x���=�F���fӾ�5~���㽊Y�=�V ���罜؇��3�����?���?Pi���J��:���I�~P���>����������ĳǽ��}����ź����#=!���`���f��)?VY��п9���<v��GF?���>�'4?%!��/,���e�M��>j߫=�@3�G�*�����ڿV�ƾ�~z?��?@>?����=Z��>U7�>���=Į>��׻���ؾ���>Z�i?�s?ǶH�?����aR��\�?�9@�B?�+�X�xS:=���>	8?4GF>��/�f��6F���>i��?��?g�'=X��&�/eb?��<�@�5~����=�S�=��=~�$�G�D>�y�>�m��Z=���ͽ;lI>���>�&�uk
�Ca���`<�.p>�1ܽڶ���Ԅ?"v\�f�8�/��T���N>3�T?�/�>�5�=!�,?C3H�}Ͽ��\�.a?}0�?���?��(?�޿�L͚>Z�ܾB�M?D6?� �>�a&���t��k�=��*�����㾕$V����=Ц�>(�>p,�g��ʁO�>/��h��=�������(�D��]��<� ��.�Ľ���mϼ�C>�D���`þ���ͪ=?^u>�̇>胔>)�7>��
>�k?�L�?�wy>�(��O����ĽhyϾ6�Z=�������s�K��/��������v���?�����w��3ܾnvK���=��b��ۜ�R���;&��Q���?�+�=V.���G�c~�������4ؖ<�]1��_��/��`m�-g�?J8?�i���EH��ם�Z�>��ս�S?
��jm�:þ�B>�ֹ�#��<�>�~=�g�]%!�$+?��4?��?BP��ь��qo>�����ý �&?��?�|�=���>��?�ج��k���Њ>�E>?�>d��>���=�����ƚ��?o�c?,�S�󝕾D�1>���Ym����S<��>R'm��-�H
$>�u�=��M������Ԛ<!��aY?M��>����W�k#>�:�h��=v�?FZ�>L�x>�1�?��4?�m��5୾ӹ8����cB�{1]?�_]?lm>uE��J�f�ľ�A?r�S?��>X���*�\:�A侅�?cEa?o�=?༢=uG\�v���;ݾ��%?��v?�r^�(s��N����V��;�>[�>���>��9��k�>}�>??#��G������Y4��?Z�@J��?��;<}%�Ҝ�=�;?�\�>��O�0?ƾ�y������M�q=� �>j���{dv���dU,���8?Ƞ�?Γ�>{������Z��=#��m`�?�2�?�,���L<?��7ml�G�� �<=�=p���?'�p��7�g�ƾ�
��R��������>�@��Θ�>��:������ο~��c�о�'p�"_?��>��ý�ģ���j��u�JUG��9H��,�����>��> 
��y���{�~r;��]��I{�>gB���>��L�]ݵ�"נ�}]5<sݑ>1��>��>�	��bƼ�N|�?����e/ο�۞�$`�?�W?)��?Z��?T�?�s<]bt���w�Y�pH?�bs?>�Y?߈-��,]���6�X8j?~�
��5@�q���#�
�{>־??ª�>��g�a� ��=�?�E>9�.��6���˲��n�P��?���?�l�0,?	��?W�.?;�S��ǿ��ax
�=�q?�<>C!�#H���4��G���h�>Fo*?U�Z�F�#�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?4�>��?Ȓ�=�C�>�P�=A����4��[#>j8�=�<>���?��M?d�>�=�8��/�QLF�HR����C���>��a?��L?5!b>w鸽��2�D� �<|ͽ�>1�j��^@���,�/p߽�j5>��=>��>��D���Ҿ�_,?�a���пu���'�+>˻Q?2�>a'�>�j/�@�
�v��v*�?���>u ��ି�Â�"�ľ�r�?\J @m��>��t��=N>���=��>�Պ>�߁=#.�T���2�>t]?GT�o�a�MV��D�>P�?�7@唩?Q��	?���P��Ua~����7�_��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>!�l?��o�O�B���1=8M�>͜k?�s?�Qo���d�B>��?!������L��f?�
@u@`�^?*�տ͗��
���>��f�	>A��=uQ>|k���=밳=�h���)��Y>}-�>
~>�>)�>��#>8�>����=&�	���k.��.�D�`@���*WG�o
��[�����ʾo���׽3�Y��DF�f$�OB��Zs���=�t?~)W?��s?5D�>���;$RB>`��l-���Nb� ����<��&?/�a?��??N��>�*��sI��ځ�'	辐�����>W�=���>v��>��>���;�^>��9N$Y=˰6>���<�t<�ȗ��C�>�|�>/��>�Q�>�?:>ߪ>M"�������e���k�Uҽ%١?����SH�$y��e؍�t����͛=��,?͎>���E�п��SI?3������&��>��/?�V?�>�e��5HV�͝> ���,f���=r�o���)���H>�?�<h>c�u>�.3�~8��P�e����~>��6?#g���49��t�l�H���ھoP>\�>v�p�yܖ���~���i�*m=��9?�?�Y���Y���-u�z��MS>�*]>��=S�=H<O>d[�㿽0�E��<=^A�=�Z>�[?	 >��=ﮟ>Tў��]m��Ũ>l`>��>��/?�?�䀼vD��{���3�?�v>���>�y>q��=�IS��S�=�`�>0l>݉���n� I�W_��>=���v�]{ѽ>��=E�����>�K�=�ڽ��_�X�;�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�j�>����[��%����u���#=w��>f5H?R[��D�O��>��x
?�?�a򾡩���ȿ��v����>��?���?p�m��=��@���>ٟ�?.hY?�~i>on۾�}Z���>׿@?KR?��>�8�n�'���?��?<��?�D`>�a�?��i?g��>��ݽ��)��6����|�0�%>0<��>m�>EȾ��>�B匿6 ���Hj�S�����\>V�2=8��>����¾�U�=�=%�Bf��S�+���>��>��(>pL�>�?O �>׌t>��Y=�H��m ��w ��T~J?��?�� �krP�ҧ�
;? ��5p?��#?�)�:c����>~�?�9�?��b?�s�>K�þ*���X����ľ]��=ɱ?>��?��>B�ʼ�U�=wH���Z��z�>e,�>1ә��I���N���t>�=�>{�.?k/�>󡴽t�?�p(?�k�>y��>�`U���.N�t��>q�?v��>��?�;�>�������|�K����(�z��>�?L?�?��=j͝�Ά�����>b�ʽ$`���߃?�H6?�ν��>�CF?eO?��d?�"�>�I�=�Ǌ���:�˭�<>�-?f�y��� ����sU`�SK�>��?�6?oo��_$�X��=�@(�}�\���3?\lI?�$3?B��YC�	�6©�� �<����w�==P;I�� �=�	>�l���`>��\>10н�Ԯ����=J.�=��E>q��>e;�>�㵾V�����+?pX��������=m�r�\I���p>�I>��Ǿ�[?��E�v�>í��w���Ui�a�?:=�?*��?�����.h�B�:?.��?�?�m�>�V����վ(V�{j������;��g>e�>�;H��㾏f���k���������+���#�>�*�>n?w��>��(>wӵ>d���/� ��.����	���@����<)=�r�1�פ�6ߧ��?)��P���ž_1}��ߩ>��M�j��>B�	?`�B>)yU>���>��<��>;Q >,�r>��>{Ov>��P>jR�=��[�W��e�R?P���%��%�m����^<?0/e?ܱ ?=���������#8?K�?_l�?S�x>��c�:k.�t/?}\�>�Z}�cK?��M=����fF�=����8ե�H����>a����<��C��h]�S~?��?,��wӾ (��y���<y$�?c�L?� P��[�o�E�Jpt����[!!����IHG�� �[�v�<�������q��������=��!?�%�?�{�m�׾����CX��+�'A�>/G�>��>��?���x�G��i���Q�_����
?qz?f�>HgM?`)F?}�I?8�:?���>3��>������>����v>G��>��B?�_B?��D?Y6?rlJ?{V�>�~/��&��0�V�>Q�>F�?���>
M?��)����<���s(�=�|��nQ�6�λ�<<=��+��4��.T�=5��>��?/꽆//����2��>��!?H��>�?�ǥ����u>?��>B��>X?�>|��c9i�f���N�>x�y?����{3<Rt*>���=4���tR�<ڶ>����x�G�A$߽�r���].>���=�ȭ<�=���Ԅ����!���>��?�V�>�[�>��� �}1�x3�=�a>��Q>4&>��վ!����'��Me�6�j>��?䌴?[]a=ۀ�=�
�=h��sO���������
=E�? "?NqQ?�S�?/t;?��?Y��=��L��������3��FP?I ,?̇�>����ʾ��N�3�%�?`Y?R;a�����8)�́¾�ս>}\/�n.~����|D��4������y����?0��?9A���6�"l�i���lV���C?�>o_�>\�>��)�y�g��$�c";>���>;R?I��>�I?�q?o-J?�X>��5����ï��Vų=`�7>1?��}?��?��p?��>h�>y3 ���������X��-~���{=8Z>L��>�9�>¬>��=ӍZ��[�?8�� >�~>��>B˫>/��>~�`>�h='�G?���>7Y��9���줾fǃ��N=�6�u?/��?��+?[|=����E�C���I�>�l�?��?2*?s�S�w��=�ּ�߶�'�q� !�>�ٹ>�0�>�ѓ=�iF=�_>��>���>�/�,`��o8��mM�M�?~F?��=J=��ܚI�d���.�~�.=�#�-o��'��&�=���}>�-��MM��OȾ�}�@M���$M���Y�F��Ƥ���?���=���<��=>�9�=����Ⱥ=�j8=@�.<_���1=���C���2w3�_v����)�;<�="�?˾��|?�rI?�+?2.C?(Sx>�	>�7:��>|���?��W>w�X����C><�X��i����ؾ�V׾Md��y��C�	>L�B�Q`>Y�2>��=��x<�U�=��w=D,�=��Ļ��=I��=q��=R�=�h�=��>A=>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�5>ȥ>��R��Q2��#Y�p`�?h[���!?5�:��ɾ�%�>���=>�޾xtľ�1= K6>P6a=���Z�[��Y�=O�w��.=,�j=-Ή>�ZG>�ֻ=a����l�=�E=EF�=�M>�� �8�/�u6��y<=���=:�^>��#>���>v??X0?�ud?�?�>��n�-[оĦ��K��>��=�>.9�=@>D �>k�7?n�C?s*K?�K�>�=�R�>�<�>D,��m����/��zU�<��?̖�?�;�>G�D<'wA����ѕ>��˽
e?��0?��?�E�>XK�Û�^(&�0X���6�	�<��=J����@=�E>d;�p5��-=g��>���>j�>��>���=�7>d��>���=@�3=��u=.�5�~��=k)�����,�=&�>G7�<�J��#�x�!= ��;�=텽�?k����<�>�%�>��)>SP�>	�Ƽ���S�/>�X���LS�� !;�n��\��ńv�����A�J`��H>F�x>(|9�������>%R�>0�b>NQ�?*�l?,��>�UW�'���ݣ��w��a=�v�=S��=_�K��8��]��O���޾��>��>4�>|�>��9�DYK��9>߹�=���H>�Tƾ��>c֖��R��դ�񖑿k�M����8�/?Q�}�J��<?6�?��+?��u?��>ŧ����jB�>)1.�t	0�=<Ͼ*&�#�=e?(�1?^��>f:��ԟA��Ⱦ����L|�>��3�w2T�޴��H�-�CּWv���u�>�Ȣ�uvξj�2��\�������E�$v�+�>�7P?D��?�FM�V����P��%��������>�l?�֠>��?H?S���FJ�hDm�.��=O�h?�D�?��?�>0��=l�����>5	?	��?�̐?^u?�3���>v!���>[}���M>+#>x�=�>9�?X?�?G��r�r���i�HMF�1�=��=lܖ>^�>-�m>D�>O �=���=�UN>&�>l}�>۰d>We�>� �>�#���y�)W)?�,>��>�:+?ڪ�>��=k���h�H<���Dw�s�=��(߽es���<"C����-=��݄�>$Ŀ�?j�W>B���.?%�����[�6F|>�`>pؽ���>ct8>�3�>J�>-�>72
>آ�>�>�%��T��=��1��5.����e��U辡��=FoX���%�y��l���J���¾	��	W�;Lp�"�j�x�p��ϐ?Sy��1W^�C<�o]���>�3�>�b?�
��cjH��b�=L�?�|�>���HI��/
��>���?���?I<c>$�>�W?�?��1�3��uZ���u�_(A��e��`�2፿/�����
������_?��x?'yA?J^�<�8z>"��?T�%��ҏ��)�>�/��&;��=<=�+�>	+����`�A�Ӿ&�þ1:��HF>T�o?�$�?�X?~UV��1��}��>P�M?��4?vZl?jq"?��_?�a)�b�
?i�=�y ?m�>q+?�[1?=(?*j�>�w�>M!�=Ձ��c��]�U��c3���Ƚ^Tܻ�3��0��<i��(e =%1>��b=t��f鵽AM������ ���ֿ��sc<��U=2g�>��]?�	�>���>�6?v)�W�7��-��3�.?��-=�?��x���})��k���P>�bj?p��?+cZ?�*b>P�C���B�%G>�+�>2O&>��\>���>��x	B��Ї=9�>(>͢= Z�Uf�� �
�~2�����<�|!>�}�>#��>�u<<M.�>���Ɓ��t=�=��y�����ֽ��̾G6��m�;)�?*�s?�.(?ϐ>��侨�����r��{)?R�T?�o?�@?2e>%_���M�cJI��,M��(E>�)=�7N�2Y��>���v�K��,P�U�>O$��|پ8��>ˡD���T�1+��<����8����<�b��}�>��#���6�]���A�^���=��L��}��褿�EO?=0�� ,3�����s��d�>P��>)!D>�7轴�л�/�O����=LF�>�>!����߾KF��
��j�>�rE?�2_?��??ʃ�@�r��PC�,���<���H����?��>\;?PC>!֩=�Q���c�#,d�g�E�mg�>��>���)H��"��@�"�eB�>Fp?@I!>C�?��P?"
?nl`?P*?\"?=�>R蹽�N��_�%?�g�?O|�=�����W�	a9��
G�|��>z~+?Dd=�3�>X?J�?;�&?��N?O�?��>�'��2`=�m��>�9�>�>W��Z��D�c>��H?��>g\?k�?�VA>�|3��G���c��Ҍ�=��&>��4?��!?{.?�z�>��>8��E�=6��>|c?�)�?��o?�}�=��?��1>��>]��=y��>>q�>r?�oO?��s?v�J?�2�>��<�������v��V�c�;w�P<0�z=42�y�s�2��2��<>%�;絳��҃����QD��拼M��;*��>�]t>r�����>4�Ҿ�6��珆>�(c=�b��Z���d�.�y=���>��?+J�>�z��{<���>���>���!"?�V�>\ ?KE.<��[�$�̾�\�Y~�>��G?��	=f�i��,����b��[=�r?O�j?W������Mb?9�U?@v��9�^˾��u��ž��T?۹ ?��U��ܺ>߈r?��t?N��>H�<�(�^������S��\�֊�=��>��w�[�Z�>xm0?߀�>��M>���=�����|�sf��.�?uN�?�Ī?���?Fk>[�w��޿Kb��SG���"^?��>E��e�"?|F����Ͼ}���D���C�UǪ�1������\���E�$����5;׽>�=��?�s?�>q?ۼ_?&� �*�c��^��	�� OV��&�����E�yE��rC�n�n��b�����> ��Y�H=c)a� I���?��7?{`2�e�>�(B��.��2�'��>�%�D8=�<Q����?1��'�=Ÿ��W�H3��s?�I�>���>�93?��u��7���-�L�l{Ǿv��=�?@��>�N�>��<~��л5�%Z��W�uaA<��v>@�c?�JK?zp?Q�+\1�%D��p5 ���׼{L����S>��>	j�>5�O��!�(�%�$K<���o�
��"��	��ur=./?�X�>���>	�?~�?;m������m�g#4���<.��>8�f?���>�^�>�4⽞t�_8�>�l?׎�>TQ�>�r���"�x��g�޽C�>�!�>Cf?�*�>�6�R5R�B����卿��6���>�<e?�5���M����>WN?c8k�[�<�Y�>��B���j��Ï�ƒ�=��>2��=#>��\���z�i4t�T)?}3?K����*��S}>��!?�>�Ф>5�?���>��¾ȉO���?��^?1sJ?�FA?���>=0���{ɽ��&�f-=�M�>�:Z>��k=4�=����\�n���C=�8�=˼���O=<{���Q<���<�?3>l 翕�?���p"�XǾt.⾯s��wP潜@��~�ɽ V��L ���
�e� ��Xl��q����,c���Ԇ��?�%@�u�I�ʋ���B��&@���>�,(���=�X��.��Ty��o��_V��e �H"5�ۀC��V��x+?�o�K�ÿ%Ð��2�=v�e?h��>L�=?��F���B����> (>^����rܐ�#�������ۇ?ԋ�>i��N��=2��>��>6�h<Kmy>5��8�6��b;̆?pU?σ�>�&��?���uſ���4��?r|@{"A?o�(���J=�)�>��
?p>>9�4�/	��|��4�>yǞ?6Ί?A�I="�W���	�G�d?��/;�{F�l�p�C��=.P�== =v���$K>Ǳ�>���1B�c��s4>-�>'����n`��9�<tKY>��Ͻ,X���҄?�m\��f��/�&T��o#>��T?�A�>�=Ȯ,?�-H�dyϿ�\��1a?�.�?���?;�(?n(��>G�ܾņM?9B6?n��>6\&��t����=5�ἆ᩻���AV���=ߕ�>F�>0�,�m��8+O��U����=Q��;ɿ�(&�wh�&@={k����Ƽ]�,���?��󊽃����c�9��[�U=a��=�ht>�ێ>�19>��D>e�c?%�v?u��>Wd�=�r���{���Ӿ���=�K��/"�����ٱ7�>@��&�ھ���R`
�^���J�v���ULI��A>�g��8���f��F��Z��c!?��[>�?����G��ǽ�쳾3���yżT.*�j����)�S�k���?d�P?�_~�b}^�'�	��K�=UL�<G?��K�Q˾^����	������U���#�>�;=�=Ծ� ��I���2?�?�ѭ��/����>,3�=�5<�|/?�o�>w���)|�>EG0?v�<�p{;��΂>H�>��t>���>�B>�߼���c�q3?�Y?#, ������+t>�ʾ�b9�uݫ<<�>V��Y�<xDH>f�i=�Rp��E�<3�k���z;�]Z?E�|>����h���������	>y��?\�>5F>��u?�H?gA��󳫾�*��d��@����Z?�VZ?��>���۾�Ѿe?l�e?Bo�>�(�V}��[C�x���|	?w_?~E?��>@Pu������ZҾ �?��v?�p^��o��q����V��-�>�W�>���>A�9�Wn�>��>?#��F�������^4�1��?�@w��?��<<s�4��=�@?w^�>��O�:ƾ]l��������q=�2�>�����^v�����t,���8?��?.��>����3���E�=�6���N�?���?�Y��$�Q�����"q���]�<�io=��";$�3������;��|ľ�"��W��޶��>�>��@�i��h�>��]���߿��ɿ ���bȾFǁ�>�!?_ܕ>��ͽ&���_1o��+v��K?�}�<��~n����>o�?>�z�C11�;�`�Z�:�WG/<[`?
2�=�҆>�Y=ԅs���̾Ѥ
>��>w�> �<>�Vn��U��(�?�?�3ſ�뫿^�پ�Z?k�?,ʔ?�՚>��'����1;�8��-�P?��?��A?�sn�M�;��
�� lg?�v��[S�$�������i>�?߻}>��g�����p�=ን>ϧ<=:���g˿A�ȿ�9�qM�?03�?�,��dO?�ۛ?��(?��{��h��d�T�Q�C�h��YsH?lkp>��S4�(X��I;K?�uA?y;#=�G�]�_?"�a�G�p���-���ƽ�ۡ>��0��e\��N��6���Xe���Ay����?K^�?c�?���� #�b6%?�>o����8Ǿ��<���>�(�>6*N>WH_�m�u>����:�i	>���?�~�?Yj?�������V> �}?*��>�6j?�t>�?��_=&y��KhW�7C*>ue>�F���+?��w?m�>7�@>��J���'�1�2��W��⾻iL�}��>�a_?�`z?O�=�ή��#��(0����=�:��H=2�����B�� �v�=��>B�$>s4-�씟���?ٜ�|�ؿ�T��q�%�<_4?o��>~�?'��+�u�E[��9_?Ǎ�>� ��#���A���+�u��?�W�?;�?�w׾�;Ǽ->��>�{�>�ӽ�#��%����7>��B?|��A���_o�_�>T��?�@�?	�h��	?���P��Qa~����7�c��=��7?�0�$�z>���>��=�nv�߻��[�s����>�B�?�{�?��>�l?��o�H�B���1=7M�>˜k?�s?�So��󾂲B>��?������	L��f?
�
@}u@]�^?(�hֿ����AN�����H��=T��=2>N�ٽ8_�=?�7=k�8��?�����=^�>7�d>�q>�(O>�`;>��)>���=�!�r��^���D�C�����f�Z���Xv�cz��3�������?���4ý�y���Q��1&��>`��=Zn?��W?r�p?��>���<|9d>Rĭ��B������$󯼤#>G�a?�i?�&?;�>�]:��N�����⾻iH�ڃ�>�U>$�>�>�>���>L�׽ɑ�>f/�=!�v>^�"> ��<h�/��<��G>���>ƭ�>]�>>�>Q9>PC������K�����%����?����'������$��_q���N�==%?��=x��0�п[��^2L?m�������Y����P>�3?·Y?�e|=�.e�Y�L<�f>�.
�wG>4�|CW�a�!u>��?ئi>dx>�0�j�8�XO�ߨ���ކ>Ǆ7??O��1+��Tr�T�I�%�˾��]>{H�>��#<J���ܖ����~�l��wy=[8?��?uK��款ɔ��ј��x�H>��f>v�=s*�=�G>���MŽ�B�}ؗ=)�=�gJ>-(?�L>�c�=IĦ>�Ġ���m�or�>*�/>�l%> 8?Զ#?�c���۵��䄾��,�%�V>w�>sX�>$
>Λe��<�=�g�>SIy>��*oc����jB��Ss>��5��(j��iG��@�=<������=��=�ֽl)I���=�~?���(䈿���d���lD?R+?c �=��F<��"�D ���H��F�?q�@m�?��	��V�A�?�@�?��L��=}�>׫>�ξ�L��?��Ž7Ǣ�ɔ	�&)#�gS�?��?|�/�Zʋ�=l��6>�^%?��Ӿ�i�>h{��Y�����u��#=��>�7H?�T����O�� >��w
??�]�v���m�ȿ�|v�u��>��?��?p�m�QA���@���>Ѣ�?fY?�ri>�j۾�_Z���>Q�@?�R?f�>�7�#�'���?&޶?���?TL>���?�;q?8��>&���[/������g�=��ֻ6,�>Y�/>�Lž%�<�[O��ƈ���e�\�9`m>U=Oɶ>��ս�&���u�=7~�����^�����>/�|>S�Y>k�}>]��>���>Z�>�l=��<�1ٍ��	��*�I?rP�?/h ���b��6�I<̭J�8?!I"?X;"�����p>�Xo?r@�?)si?��>��E������gƾc�=��`>^��>/P�>������=��о�nf�}��>���>B���ݾ�x#�}�:(�>�d>?>�>�����7$?�L?���>XN�>G��H����'���5>�?���>H�v?o�?���9�-�B��~���N?�S��>�o?�?���=W���\��D�M>��<��=����?R�?�L���I?�vu?8�>\�c?�;�>�\e�� #�aB(����=b�$?Ӭ���/�_]!�TvJ���>��"?H�?�3���Q��]��_r��V��6�?��f?	U.?�f
�/�N�b�ɾU�*��'r�_+<V,<ɔ��q�=��>.�ʽ���=��X>"	;鼂�+����a�=���=Dp�>��>[ߚ�KdK�nh+?�/��\y��3o�=/t�!�D���>�[7>��Ǿ;�^?�P?��{�H���ɝ��de��T�?GN�?\V�?Rǟ�Qi��8?��?�?�}�>L���Hؾ� ߾p�g�	Qf����g�>��>�ؓ�$�ؾ�\���먿�郿UV�������)>"��>�#?O�>c*�=��>aܾ�!�Չ��2q+�#S!��	6��[f���#�8<��S���ҷ��lE= �8����x�>"*~�/x�>�F�>c�>��>4?:4!��w+�V��>X�h>6��>���>!��>G��=?5� R��_T?�	��o�����iK���?�$�?��5?�\\��H��]y���?Jp?���?T �>U6B���c��>/?A��>=���.�>��,=f<� ����Ҿ� ��
�gټ�R�>�p`�XwH�����2H���6�>��?�T�;Ů־���ݨ���B&=�ч?��.?�{3��zT�`��Pb��\7���u��s������u��>�����=?q�0 ���=
,?�R�?������nd��A�o��L:��S>�I�>�L~>�}�>wl�=-�	����Ga���*�u�~�k��>Į{?��S=�Xt?�(N?9D_?��8?��>���>�:��J�x>ё��O�>�0�>5BF?ЯC?�WG?y�H?��o?q��:���/
��羺t�>�:?�A?�L�>�Cj>�ǽ���:��=��(>0hR�e�$�s��U>)�=�o׽�gؽ�׆>�"?0�6�X])������>[>��?�&�>O��>0敾 �a�i">"�?̊�>��>���/'q��X�VH�>�r?�fX�:_D=�� >���=�n<o���xv=��=h�<Q�������=v�/>a.>�>J�Y=&b=n���g�� ��>w�?,A�>F�>Tә�������
(=��|>�I>�,>�>Ѿn釿�����mm�؟b>q.�?a�?�/�=ѕ>��>����;י�.ʾ��-<��?��?��M?��?A�-?��?�y >$��q��ӄ���j?�q,?i\�>e����ʾ�Ѩ�3�~�?^x?��a���>&�h���׽{�>[�+���|�ɞ���;@�K$)���pL��bZ�?D��?ZN�Y@7�k��"���2���oC?�#�>�D�>��>*��Ig�����:>���>��P?<˹>��Q?��v?�e?q�>��8�����#���L�=V
>tDM?���?'��?�q?3h�>���=�J)��)Ǿ��ھA�;C�C�w���=\�Z>ݡ�>S$�>�7�>v��=xY��*�cǇ���=^g>� �>$�>��>�v1>?�B=��G?p��>�b�����j䤾���=�:�u?��?��+?�1=c���E��B��>I�>�m�?]��?-*?r�S���=�A׼�㶾d�q�)�>ݹ>�4�>m��=�F=5h>��>��>�!��_��q8��DM�4�?�F?M��=�@����h���_�)e��mt�<�E������� &*����=p���vf/�K������e���;���T���|����{���1�>1�g=�f,>��=3��<`�&���5=߉X=圃<!Mu=�a�����<i�u�A��;����~��<�<�۔��*ܼKp̾J�}?��H?�+?pD? �z>>s>��2���>ah����?h�S>ޒP�e�hr9��ʦ��o����ؾg�׾�0d�1Y���=>��S�#>q�2>���=���<���=�Us=�*�=�_�Q� ='6�=�^�=�̪=�=�>)�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�>4>��	>;zR���5��gU�<O�qQd�� ?~�:�Q%ľgE�>7֣=D�߾�濾�G=�g,>F==;��[�tͩ=�@��,%=�l=B�>�kC>�v�=Q뱽��=x�J=�}�=[DW>�ڪ<#��	l����4=Uw�=�N>�>�Z�>-�?�n0?�i?Z��>���Vᾍ,���ۧ>N��=���>t��=�>�w�>�+?�*=?��F?>�>"z�=��>�g�>\�+���q���ξe���LL�=B�?:�|?�>?��<_�h����E;/�V�T�k�?��)?�?k��>۩�
��48$�׍��>5�Z��;�S�=�*��0
a��炼L�����ѻ�=*j�>�P�>��>��>җ>��J>���>��>6=�<=vm���=��̼v�T=|4�<� <T�U<+�=ert<LDk�`S�<֓�=|�K�k�1=�w<O>蒯>�U8>���>+�!<�i��fwD>k򽾁�O��$>x*����;��d�$Ѕ���6��Tc�_/>(f�>V3<�_����>>Ś>��F>_��?Yq?��>����㒾򲒿8���c��@p=F�>�����6��i[�2S��fþ�9�><}S>l��>���>��8�X(B�'(�=�f��[?�i��>?���UNʽ2�U��5��њ�������dR��>C�A?�����J�=_�?�B?�g�?���>ēU�lZվ�q>�b��'u�.n�x�q�U��?�)?��#?���>=��B7��ɾ�s���)�>�A��Q�t���Q/��������#9�>�%��OX;{[2�Ә��)X��w�A��uk�,��>[�O?*l�?��Y�o쁿�O�%�ZM����?80f?ȟ>��?��?44��Y?��x����=��k?�#�?���?i>
���u�;�]�>�'?]�?R��?�MY?��?����>��üF�>���d=K�=��*>��u>}?���>p��>�3�^�y��p��zi�y�g=M,>㎟>�L�>�P>K�Ի?F�<_8>]~/>��@>J�C>��.>�>k�}>�P��M� ����>
< ��>?!G?� ;>�V�@|�<�%_>� ��:R�T[���I޽��(="s="P�I�����>p�ǿ랃?Y��>�Ǿ�u?���������>��[>}|���?WQV>	�8>"~`>�>|D�=�_>��>����Ⱥ=�p$�NZ%����M���Ͼ��=&U�}л!���⽽��
��u������U�%�r�fR�}�:��?cċ��X�8`�����S?J�>N2?�盾os$��>Q]?��e>k:��x��ȇ��I��S�?ۤ�?6@c>��>��W?�?��1��53�nZ�زu��A�re��`��܍�����1�
��X��ѽ_?��x?uA?��<QBz>���?4�%��ߏ�7$�>/"/�k%;���<=X*�>'��^�`���Ӿ�þ!��:F> �o?�?(Z?�=V����a>;�.?�,?+,x?�f2?�Y5?�J��[+%?��>G�>�Q�>��)?^�&?|�?߽�>��E>^��U	�� ����z��'	�5!�a����=X�=ݷ�<g"t=�0=���+�Ҽ�L�<үA=Z2p�n<��k=7>�q�=r>��^?�D�>u�>�DD?(_��3�9H��� ?tg=��b�����^�����Y�@>�yu?Pѫ?Ä=?3�<>d;Z���g�%�|=�uX>mC/>h�c>��>9⼽�
��M=	�=���=�='k佨�������M���7&=��+>k3�>��>e�=��/>34ξ�!��I��>���;M�5����&�(>����=ǌ?�z[?g�5?�>������o����7?w>?�La?:KV?���>�����5�X�G��{��d�=�x�=d�ľ���*��yqE�ô=b��>s8���f�0��>;D�T�g�b���;��<���
�f�8�h<�>��%��"�?p����>�z�>�3����;�x��ٯ��t?��½����X�R����>���>�~>`�l=\8��I_H�W�����&>Ǽg>���=\
�վ.�L����,��>�lH?�_?� �?Ԭ��zp���;�l���)��x5���?���>,5?�{N>���=�Ҭ�����me�)H���>	�>�)�H�A�1��>���Q)$����>�?y�;>?�P?*!
?vU]?��+?)c
?��>W��Oo���D&?��?���=�սk�T�D�8��"F����>X�)?��B����>�?e�?/�&?ScQ?)�?��>�� ��.@�ҕ�>�?�>��W�2a���'`>V�J?��>8Y?tɃ?>>�v5�A䢾�;���x�=�N>��2?�:#?�?���>p:>wȁ����=	I�>�'�?��a?&d�?�*�1�?��>�W?�6>�^N>��>�9?�~?V�?X�7?�n[>	�<�v�{�����*�<��=5Ƭ<w�)�hX�< -�<��=JQ�;��-����W'�<�)�=�<���rk��Ǽ���>�ʀ> &���� >D�ɾM���l��>�MW>"���*���y\���=�!�>?C�> � �ʪ3�CG�>=��>�C��]%?�"?[m!?xwԼW�W���p	����>e�T?�w'<\q��/p�;�U��f=��u?Tǃ?D�����&�kPd?}]N?�z���Y>�0����#G�#����B?�G&?�CV�>PC�?��?�O�>�~��ҷj��}���e�����G�=�v>�� k�y��>��M?w��>=E�>��=,¾�D_�����?�͊?&v�?2ip?��l>�~h��B̿���� ��l�]?���>�S��w�"?�Y���Ͼp�����$�t����[��՗����$��	��`c׽Nl�=��?ts?Gq?��_?����c��]����W)V�B�S��o�E�{E��zC���n�v�m����Ƙ�Z#J=�K��PJ��9�?��4?1>`��B�>�d�����ӥ��+>�Cɾ�b�6��ql�ث�;*��5[R�c㗾Qy?�^�>��>[O?��c�E�8�;)������о&��=�&�>��>�X�>NrA:��'����oi���<C������@v>�c?�K?G�n?���� 1�
t���s!�H�1�-����qB>�g>���>�[W���W5&��U>�t�r��������r�	��,=Ԙ2?!�>���>?�?��?�J	��C��qJx��g1����<Z�>�h?F9�>W��>�н�� ���>��j?B��>gT�>C�����4�^���AS��&�?2>#>�f�>���>��F�N��ᑿ���Rg7���>�a?�k��Ā4��y>��6?yͽv�=�u�>�����
W��!�41M=�|>��<�>�����|�1�P���$���(?�?�����*�ǯ�>��!?���>/g�>mb�?��>zN���G<.�?��]?��H?�@?J��>^!�<�>���hƽ�7&�ȶ-=���>%}\>̭p=q��=_R�xrb�����uG=��=ਿ�n	��3F~<>:���Ed<J��<�3>��ؿ��D�Y㾝��1Oݾ^���Ry��۽�W��A*���/�������x�hx��f켛|<�y�M�ӭ����s�.T�?��?2͂�"���y���rg��\���>���Zg�m����� �-J���۾���D���N�d8j���d�F??ڿ뾬ǿ�$��Eݼ;�vj?�]�>'N�?�����1:�qRC���c>��<ɊZ��긾���#ο9���V?�b�>Q���B�>��)?=�C>�&���?��I<	��ώ�<T�I?��?K��>%j�=_Ļ��1̿�+= ��?#@�A?u6(�x��1=L=�P�>�^	?�U:>��.�Ϣ�Ψ��3q�>�S�?N�?��N=��W�j��l�d?Q�;��E�š���=���=�4=
/��I>呑>FD�R�C��~ٽ��4>>�>�( �>����Z��[�<�Z]>+8ӽ����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=u6�󉤻{���&V�}��=[��>c�>,������O��I��U��=g��0����O�{X���y>i�$>\em�.�<�FiU=?��>��þU���f5�Cp�<�&�>$Z�>
5?��>{>R��?�1�?l�2>-�5��p=�Ȏ=�[��ɼܾ��U��욾 ��>;�#��ٛҾ���s���$�_�˾�G:�q�=�7T�������G�F$S�� ?{�=�~���PL�@?ռ��;�ᚾ���<Gbv��Ѷ��0�GIl�t@�?��:?E�y��IS��f�/��b��OR?x�7������}���4�=��ļ��=�>��e<�x���!��)P�8?�?�Щ��u��^Y>U,�g�w�s�(?�&?�p�<�>�XC?���=x�ν-�=���=�g{>Vn�>S2(>�oǾ�=;B�3?v"{?z�����T�y>7렾����!��"��=0��t}1�W�>�f��nf��ܯ�2!�=��9L_?�ΐ>�*"�߳�ں~������>l�s?,\
?��>u�y?�wA?M!�=�ʾ�5X������(�x�1?C[}?�!>���w&�~ľ�}1?�b?���>6��<�4.��h-��f�*p�>)�G?�??w>�g�)r��}���7?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?r�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=ߺ���h�?aW�?�@��|�;<��hrl�P���r~�<��=�.�N�*�9^8��]Ǿ��
�딜�Կ���*�>�7@�}�
��>�n=�h��;�ο+/��
"о�;q��9?&�>�)����,hj�.�t�N)F���G��S��K�>T�>^���ȓ��{�6":��t��#�>YF��t�>�\T��E������&�A<
�>��>�&�>Ŷ��9h���ə?F����Ϳ�u��W>��X?�J�?5'�?ڐ?�7:<$pu���|��j��GG?bs?��X?��'��f[�x�;��s?O�V	O�l�ξa����=4?���>��=�sG/>�b�>��><�>Y��K༿W�ǿW9��a�?���?^����?)��?�4?]bR�xլ��.žZ�k�:�@=e�|?�/G>~=����2kq���׾�*?%�+?o�v�0s�6�_?�a�K�p���-��ƽ�ۡ>��0�
f\�IR�����Xe���Ay����?=^�?O�?���� #�56%?f�>Q����8Ǿ(�<���>-)�>7*N>�G_��u>����:��h	>���?�~�?Rj?��������V>��}?zz�>�?�b�=�7�>[
>�)��<���:>��!>U,��?hU?=M	?5}�=i�D��!�P�>���M�2���YE����>�tk?<�b?�n�=C�O�K��$��}ͽ�D�G��l��������>*e>�{�=e+ؽ�z̾��?Rp�6�ؿ�i���o'��54?5��>�?����t�����;_?Hz�>�6��+���%���B�a��?�G�?9�?��׾�Q̼> �>�I�>��Խ����f�����7>5�B?Y��D��c�o�R�>���?	�@�ծ?Xi��	?���P��Va~����7�a��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B�}�1=8M�>Μk?�s?|Qo���j�B>��?"������L��f?�
@u@a�^?*��ٿ}����|���ǾU	<=�V�=�D>�`
�*;>�=��7=yB���W=F�>�f>8k{>�>�`>P�	>Q܆�Y\*� ���.�����I��������7�����E]D�]��
¾��ھ'� ���a��=�<����p1��Y-�=��|?��X?�v?�G>Sh�
'c>Y���fx��^�SW�b��=�z? vX?g�6?dS>Ѷf���Q������yѾ����S�>�$\>m��>t��>��0>J�t���>�U�>�{k>+�=��!>1G9=�E�>��>� 
?6N�>��>|x> w=/���	���ë=�	~<Jgf��Ɋ?9�l��H������/����|��!?�">ˈ���]6����O?U�1��+��6Mr>��?�|F?ra�>EXO��;8��#>�i��X�%wV;�#M�;+��6C�� >��<?�ie>0��>{+���.���Q�{���%��>�_4?/�ξ\��*u��LI�`�ؾ1�\>���>�Rټ
������Y����t�0��=�8?�?%&�빲�]�PM����X>�9T>"��<Z �=i�2>1kt������Z<���=LS�=,Uc>d?�y+>���=��>���{S��~�>�<>��+>�g??z?$?����N��X�0�3#u>4G�>�G>�g>͸M��=&��>��c>�
��/��6�
��">�o�W>�c����_�Pwj���m=h<��w�=�ƍ=Y%��;�a�=.�~?���"䈿G�B`��
mD?]+?��=�F<�"�  ���E����?Q�@�l�?��	��V���?A�?�
�����=�}�>ث>�ξ�L�9�? ƽ�Ǣ��	��&#�S�?q�?��/��ʋ�~l�]9>'_%?c�Ӿ9�>�O�zR������u���"={��>�7H?����+P�7�=��t
?	?�^򾯧����ȿ%xv����>H �?��?S�m��=���@���>���?Y?2�i>�~۾KRZ�Σ�>|�@?z
R?t3�>@�ە'���?�Ѷ?���?͗]>�N�?+l?Њ�>H���d/�����QC���.>Л���E�>>wG>�ʾY0C�-L���`���n�����>��d=t��>U&�Cؾ	6�=o"��䞾-�c��ƣ>*�p>�E?>��Y>�	�>N�>8��>�w�=OR���2{����R�K?$��?���)n�ڣ�<���=R�^��*?SC4?��[���Ͼ�ۨ>M�\?׾�?Q�Z?�W�>����<���޿�/���!F�<f�K>�F�>�:�>�F��@K>�Ծ�PD�:w�>:ė>'����6ھ�)��כ��N�>�b!?y��>:��=Sh*?\� ?��y>��>NV����� v?� ��>��?�h>	mL?��	?Y���_������:w�?t7��a>-e?q�?�q�=��������[2�>׈�=:C���L?�1c?��=��?��N?~|P?:�F?�{o>�ԧ�n��6K$�P7�=P�!?#��^�A�MC&���o?�[?'G�>�����׽�ͼC���m��l?�\?o�%?�����`�a�¾2��<$�#�	�O���<,�H�iQ>ѿ>�ǆ�P"�=b�>Հ�=�-m��6�t~j<Mo�=9��>@��=��6�S���N<,?�H�ݥ��r��=��r��zD�!�><oK>���N�^? �=���{���̇��J\U�	�?!��?�^�?해���h��=?: �?9?C7�>����b޾���W!w�wrx�Kg��>���>�hp���侙{��P���">����ƽ-p`���>��?e?��x>�F=�n�>
�t���Y�����^�H��H�]f�RZ4����;����!r�[ 8�"�վ�̾��>��D�N�>��>�Џ>�W>�"�>,����=��j>��>~?�(�=�/B=1� �
�����
�%wX?`ݔ��<$�{������A�$?�:i?��<?ahI�h�����F��?�B}?Vr�?���>�%h���^�|?��?�:��<N�>��=KƜ=i�d���߾�Ž@!�=%�"r�>$�0��f'�ͫ�	k�.H?�j?*[{=r���Md��
�Y���ʼ�k�?�yK?`�N�iNU�t�C��c�h�,������B���Nu��= ��s��K��&�|��Av����X>n~&?���?��˾w� ��Qa��C9���>J��>݀�>M�>S�>A����I��S�A���P^�y��>���?���=��e?�FN?	�E?��?wDS>QY�>0`2�go~>�_Z�x1�=#g�>�SY?��;?��6?�O?�2?	5�>|�,�K^���\װ>�)�>�?���>�K�>����G�������u�Zw�`���F�u��7��1Z��=S�Պ�=��>�r!?�/��3�6���d;�>�2?uƺ>
��>�?R�s_��7�=���>??#��>�$��$r�}��(3�>f��?���9Ҥ<�.,>s>>N�W;�!A�I�9=n
�=�5�����;�;��� �=O�=s�>��$= _�<�y =�;��lx�>��?_��>�O�>Cj��� �v��Xy�=�Y>B
S>8>�>پyz��?*����g��]y>tt�? s�?�g=�0�=U��=]����z��Q��5���:�<�?�O#?bLT?���?C�=?a#?��>�%��D���[������?�',?	t�>s��:�ʾ�ڨ�t3�X�?�v?{6a����)��(¾�nԽx> F/��5~����i�C��Ix����JG�����?x��?z`C���6�t<�9���DN��N�C?|�>FB�>���>3�)��g�^#���;>w|�>��Q?n&�>��O?q2{?Ҝ[?�LT>��8�F,���ș���0���!>�@?@��?��?`y?+a�>"�>$�)� ྲF�����݂�ްV=GZ>c��>7
�>�>)��=��ǽP����>�䉥=h�b>`��>c��>{�>w|w>��<��G?S��>a]������줾�Ń�J
=��u?̛�?��+?�T=���E��G���I�>Ko�?���?�3*?��S����=I�ּ�ⶾD�q��%�>�ڹ>�1�>�ɓ=rzF=Jb>��>���>�(�a��q8��PM�Q�?�F?��=�����h��y��5����=���,��X��V�I#>�T���0�ۇ��.�[�a}���惾������a��>-?��=�i>ܵ�=��f�1�:�yU�V�t=�ny��=����W=�]D�(Q<$e���ڼg� 
=iq���"޾��z?��N?γ(?A?�(�>ل>l%Y��H!>�C��H�>Qe>�*:')���:����{��6�������@Ѿ9̎�]���cC>|41����=j�>��U>�%C�
�>U�'>fI>�b1�.�<�)�=��>k<�=��5>;/�=0í=�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�i7>�r>̵R��1��I\�g�a���Z��x!?�P;���˾^�>�T�=�߾�;ƾ�J0==d6>�9b=͋�KO\���=�Ez���;=-�j=���>M9D>0�=Zկ�v��=��I=��=A�O>>����5��l*��1=:L�=i�b>��%>.&�>�5?�0?.\d?:�>Yn�Αξ�����ϋ>a�=�{�>���=cpC>�m�>3�7?�D?��K?ky�>|Ή=To�>�̦>��,���m���侳����O�<U��?���?� �>;tB<@��/��L>�D�ɽ?�?W�0?:s?�_�>������#M4���?��F�^7j�����#i���>Ѹ_>�#0��P�ox���>dH�>�v�>�
?���>��=:C�>��+>x8��ސ&=X:�=Y!
=:�]������<m��-���_ ���>􋔽*�=N{�ݿ��\�a=��R=ҫ>T�>NN>3��>w�;�1��Z�.>by̾^F�I>}\���?G�8Xw����+3��+�];4>�vG>��$��'�����>���>GD<>��?S�o?�">�� �xHþ����<J��y%���=��= I�g�.�h�]���H��⾻U�>�Q:>{Z�>ߥ>��M���P���=3��?�+��!�>���
Ie�W �����)1�����)C��x<�NW?�慿	L3>?ό?C$*?��Z?;��>�A߽���qk`>��@���������Y蘾�?�=? #�>��ܾc�o�?���d�����>������l��o��V� �xQ9�
M��l��>{q��}�̾.�(��W������:��UO�|e�>VW?1��?���� ���<�\�
{�O.ڽ^��>n�y?��>�8 ?Dz	?w!ν8ھ\��c�|=��o?e$�?��?J�)>�������;�_
?4"?�3�?�Cp?�C�?��#��~�>�FT<0 y>k+���1�>�dG>b�4>9>
�?�c?��> �ݽ����� ����,��w:�,D�=j8(>�&�>�(�>�w>�*>��>�)�>�0�>���>�d�>ٞ�>+��>ގ��Ź
�^P(?�i�=�[�>SV0?��>�jO=����DM�<�%J�
A�:>%�t.��fݽ.e�<��r�S=�Rټ��>8�ƿt��?��P>�%�+?���>5��YW>A�Y>��Խ�p�>�
K>�d�>HĮ>T��>e� >�ω>�`(>@Ӿ6�>����^!�FC��oR��Ѿ{z>x���&�����P��� I��k���c�Lj��(��V<=�l�<�?�?�����k���)�#���D�?�{�>6?،�ł���>���>p��>�/������ɍ��w���?���?N�f>pZ�>v�X?Tc?RJH�� ;���W�_Tt�4e?��/c��\_�1 ������~����ڽ�]?B�w?�5??
��<x�z>:��?Nh'�����Ժ�>Pm/�#�;���=3<�>�����0X��YҾ�þ�!��WB>��o?��?�|?��Q��ꍾ�>��#? q?G��? _?�i?�:��h�?�9>U_(?*?� ?�?ev6?<�?�"�>�0=�K���]�nwu�89:�r���[�.=���=?~>�����=ڭ�=ͽ=�\=77�?�@���(=�>	F�<��+�L-�=��>fse?��?�>9)?�B���%��B���:?,w��O{���GY���X�F�þ��.>��g?���?��W? M>S/Z�Q�^����=�e;>�n/>��Y>-�>{�0���:�=}�=�i#>�y�=����ž�؀�L����Jm=J�R>��>�<�>��<�mm>鄧��,��t�:>�˼D��&���f��?�!j6�|L?FH?;f?�X=��ھ���/�|��[-?��??�M?)�@?��_>[ž�I��\f��M�����"�Žpb$�����ٝ�ͷA�c"���>U��k����©>
� ��E���0��:��'�����F>�.Y�=0���־EZƾXy�� W�=���B�.�� ��g~��m/K?�0����^�{�] ��H\>�>�s�>�=c��=Y�M���ϞK��W�>ȥ*=��=q;h�5����u>`R?��[?���?�^E�a�{�#�7�'��z��{�����6?�	?=�?҇>���Ӿ��+�1�aqF���>)��>L�K+O�6s0����A=3��LS>�l?M�=��?��[?�k>?&�C?�m%?h4?A�>GFq�Se��A&?"��?!�=��Խ<�T�� 9��F����>-�)?��B�\��>��?�?��&?��Q?u�?��>� ��C@�A��>#Y�>)�W�b��>�_>g�J?���>�;Y?8ԃ?��=>��5��ꢾ�ԩ�S�=�>x�2?35#?#�?���>��>.�����=L��>�c?a0�?b�o?��=��?g82>;��>���=\��>���>�?�WO?q�s?��J?��>r��<;��61���?s�S�O�걂;dH<��y=���8t�K���<�&�;it��)H��H���D�:������;���>��u>�����,>}_���^��;�9>^�ڼ7��v����<��3�={�{>}� ?UΒ>�-$�F�=��>N��>F��]�'?8[?�c?�����c���پ�G���>�)A?���=w�l�_A��� u��:g=�l?�@^?i�R� �����b?Y�]?Ba��=���þ.�b�r��#�O?p�
?��G����>g�~?��q?M��>$f��:n�0���<b���j�6ö=�p�>�S�g�d��?�>h�7?�F�>�b>(�=�m۾��w�sk��?��?��?��?=+*>t�n��3��4������ƻY?���>W]���"?;�>ؾ:��Ẏ�����,��R��8���੾��%���_׽E�=g�?��r?&*p?�[?t �Duf�D"\��w~���S�������E���C��C�V�k��5��^��͔��x�=�.O���6�C�?ax-?s�IG�>�P,�O��������o=~Р�#���V.>�%��3=ȫW=��~�^8w��G���K?�H�>�}�>��1?<�s���O�w�6��<��?��sV>�ݟ>�X�>�>T30�C�+��6��Ц�ߪ����<4�u>d�c?\dK?Pn?�x���+1�'N����!���3��x����D>(>��><XW�5m��%��>��Hr�4*� ���~:	��=�=i<2?�"�>	�>��?�?&��׍���x�.n1���g<y�>th?�b�>G��>�Ͻ�q �Ut�>t}`?!��>5S�>T���R�(�uJ\�zɎ<�hS>U��>x�?_ͯ>�L��O[��q��Ֆ���T�\�>6g?�鍾��6����>pC?8w�<��;�[o>UL,�rE%��@��h鋾�]:>�?���=p�>�;�����~��<��(9)?�A?M���+�*�$�~>5"?��>��>4�?���>ņþ98�g�?��^?�J?<A?��>�==�Ĳ�TȽ�}&��.=���>�[>�h=��=�Y���[����+ME=��=pͼ�乽r <�����M<��< �4>rҿ%3*� P�� �*��k���Y����o��3p���d�7��`����tz�xA9�#�N�sC���p~�"���B=�Ln�?%�?/�x�������qJ����W�>�~�l��;闾;�Ѿ8��H��f ,�::I��Qs�E���'?������ǿ����w8ܾ�! ?k@ ?��y?��О"��8�N� >�&�<<�����o�����ο���N�^?���>���0�����>9��>�X>�Hq>����瞾�%�<�?��-?���>��r���ɿc����¤<���?��@mA?��(�_�쾌�T=���>L�	?�P?>��1��>�K���%�>�0�?��?��L=�W�[�	�ee?�<��F�	�ܻ3Q�=x��=O�=B��d�I>o3�>��uA��hܽN�4>`Ӆ>lF"�i����^�9��<�]>�kս�0���ʆ?��c���h�c�*�:���E(>��h?A��>�c�=dN�>��J��ǿ�?��I�?;��?CE�?g�#?I��E�>�FҾ��G? �@?�٭>W��t����=bc�q"��멾j�E�ɈP=(?�:>ZF�>�������f���>.� �1��2��-n��ɜ=l#�=�x��3�RK5��:�<Ï����=�6
��o��=���=-p">je>aW'>��$>R�`?6;~?8�>5��<��㽬���LϾ�d��͊��/�ֽ��~��9i�U�˾�u�i�оy��@�/`�����=�1+�=�Q�xÐ�6� �-b���F��J.?~"">�Vʾp�M���$<�ʾ}���ーډ���{̾�1���m��ǟ?��A?�ᅿ�W�����5�������W?������������=���=]��>tѡ=!�⾰S3���S���/??\??۾�"���->I8�W��<��)?l� ?Q�?<ޠ�>!�$?5-����z0W>B�1>�آ>�2�>�Q	>P��Wٽ��?v�T?ʉ�Fy��uq�>oѼ��z�O_=?�>��7��G���aZ>E��<c���Ϳ3�����3�<jX?���>S��ռ�(涾��GY�=ċ�?���>24�>�ˆ?fD?Q!�����Kk�vX'�z�=jv?/hk?���=v�������g���	-?4_?� �=I:`�a����D�b��S?~^j?�#?4�D��S������	��f>?��v?�r^�@s�������V��<�>�Z�>���>|�9�{k�>��>?�#��G������tY4�Þ?��@q��?��;<�����= ;?\�>�O��>ƾ�v�������q=�"�>M����ev�����Q,���8?��?Q��>�������R�=SÕ��t�?��?�����^<�����k�y��D�<�ڪ=���d����}�7�g�ƾ|�
��՜�U���5�>D@���k�>X<:��;⿷2Ͽ�����Ͼ:�n�#�?�>˽�����j��:u��7G��&H������l�>�/>������Mq���@�����Ň�>�V�=�OV>/����,�j�۾ӛ��*i}>q'?1i?r��=3���,�?����ʿ�Ձ��M��I?��?���?�T/?zN�:p�D�/}Ǿx���`?{3�?ང?p�<yㅾ���=z�j?G쩾�`�DN4�\IE��T>8�2?"��>��-�:�=ZX>���>�&>51/�Ŀ�ݶ�i��k�?~q�?�s�B��>�r�?�s+?�B�2��m����*�/���A?
41>�$����!���<�������
?�U0?���Y��es?��m�#E��pF�?�ܾ$L�>*�>���mk�>�	��Z����*9ƾvZ�?�A@���?u?�����bUR?��>qq����Ǿѥ�f[_> ��>�E>�6��M��=L�F�
r#�g��>�.�?��?D	?㣇�SJ��_�">I�i?p��>_z?Re>�T?f�Av���^���� >�!�>��=l
&?ؒZ?�%�>�6�<7,{�}X;��M��%�k�%�D�%w>�g?L�r?H\x>3�	�.O{��6�PO�=�gV�E_[���?�����!�lE>;w>��L>��z�N�ܾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji���?TX�}y��T�|�o���<�g�=�6?��@�w>�-�>x=V7w�ݪ�>s��%�>7�?��?��>	ul?C�n�?/D��&=�>�i?>�?�ZA<���ǲB>�?�k�Ԅ���H��g?�
@\I@�y\?����Y�ʿ�˞����g��o*j>[��>x�o>Y�#=j�V>7�=L����q=���>QNG>@'k>c�>~[>��#>���=G�z�������󚿪#���;|�ڽ+��;޼��+�SҢ��5�������e������]�/�F��,׽'">8/F?LO?��a?�U	?�8����>���l�$�f����<��Q=��)?vC?��?�>����x��f�㒰��\��n��>��`>2��>�C�>���>��=��>ga#>Ij0>���=�ڷ=U�=�<�C{�=-��>�?�]�>E�9>��>����P����f�c1n��ֽ��?&-����I���η�����)�=�-?���=0��\п�⭿�.H?�Z���l�F�#�-�	>�90?�V?�>�����]�u�>�	�J�h�D9>K��^�f�q�(��\U>"%?WLc>x�u>|;3�+�9�;H�@���u7g>
/?�ܸ��`;���t�-�E��p߾�hG>��>cG����奕�\k~��pc�2��=�?9?D�?�@��{����+v�f~���=\>��R>i�%=���=YN>�oo��q۽;�?�k�==���=�Fi>@?g�->��=%��>�B���Q���>��>>(o'>��>?�e$?<��dF��B���ч0���s>mZ�>.�>��>k�J���=���>W'd>���o����S��?��GX>0瀽��^�U�}���o=m��=uO�=�Y��-�;���"=ތ�?&]��*U����߅��O6:?�3?��7=S�a=Z�<��k��2�̾��?�,@$��?n���3�u8?I��?u�����*>D`?�5�>��}�HD�����>h�������X���{���,�?�*�?��P:�{���u�G%2>w$ ?$��Ph�>{x��Z�������u�y�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?�	:>T�?p�l?�&�>���"1�t���Ɔ�%�=�1~�>[;�>���A�:�:G���섿��d��}��ȏ->�P=^:�>�{潮������=%[��)
���2ٻү�>�*>�K>�-�>�??��>&U�>�_p=L7���7�bH��v�K?䲏?���a0n�4��<=�^��&?�D4?�[��Ͼ3Ш>#�\?���?'[?5e�>����>���濿[�����<�K>�0�>�I�>��&LK>/�Ծ�.D��m�>iΗ>q(���>ھ,���G��8@�>Mc!?���>�Į=� ?ۤ#?fk>2i�>tbE��<���E�1��>���>Ea?o�~?��?ҹ�.j3�����ء�6W[���N>k�x?�O?�ە>��x��i�F���I���N��?�ag?G�㽘T?�,�?~X??x~A?�_e>����׾�������>�x!?���AdA��1&�b��?��?��>����+�׽ؕ�a���a��C�?�f[?�%?%��!Ra��cþ� �<� �V�7��� <,5%�0�>1�>uQ��K*�=��>��=�9l��5���h<�ܷ=���>Ģ�=]�4�g���2=,??�G�{ۃ���=��r�BxD���>JL>����^?l=���{�����x��N	U�� �?���?^k�?7��6�h��$=?�?H	?k"�>�J���}޾'���Pw�&~x�zw���>���>̡l���O���ޙ���F���Žsm���>U��>���>�?[�?>�<�>����+�A��e�'zZ�q���U+�H"(�C������
X���T㼾HAj�oK�>�=�0�>���>V{>�>�|�>ƌ�����>��>�HV>�H�> O+>��$>�|�=�<=�体WR?����'�S������N"B?݉d?�
�>,pi�^������/V?ی�?���?�w>�Jh��+��h?է�>0���
?]l==ik���<�����N�|���ZU�B��>�ֽN%:�x�L��f�L=
?�?�����̾�\ֽ|c���{=쮉?�(+?�%�'P��_���E�f�D���y�=o�M�������l�:����?}��W~�#�"��=��*?���?���HX߾�rҾ��{���:���I>b��>,��>��>[�P>�6��B���]�^ &�F�2���	??M~?6`�>]NI?�7<?'hP?�`L?��>c.�>}��s��>���;���>�V�>�9?��-?Ю/?�O?s�*?G5_>	���_�����ؾ�x?�r?C�?,'?(�?�����뾽�ї��u�ߐw��s����=v��<�ٽ��p�^Z=W�R>�?����n8�
���xgo>�a7?	6�>�A�>�ۏ�/������<�m�>��	?��>\q ��q��:�qY�>6	�?����R=��+>{8�=�����0����=��̼�֒=
Q���+9��<VϽ=�=#��㯺/7;v>�;&'�<�
?�#?��>�P�>ӻ��_���nоZ}>p�>&��>�r�>�Ʃ����j���K�s��#>�?�C�?��=:P">��=4�꾹`۾���ņ��X��?�H?��H?P3�?�yI?QU�>s*">�X,�Yw��`�}��>*�ҍ?�!,?F��>V��H�ʾ=񨿚�3�ٝ?Z?�;a�����;)���¾ �Խ��>�Y/��-~�����D�~��I���u�����?���?��@�n�6�Bz����]��ԓC?�!�>�V�>V�>��)��g�4%��1;>���>TR?�ʢ>0�l?+�k?7L^?�H�>�mF��	���͡��}�=�l>j?��?� �?�pG?��>w��=3SF�b\���XK�j����Խ���u�<��|>�[�>|��>}�o��e�L��=��*�n��G�<�~j>0�>��>���>U=�=fqa���G?��>)Ͼ��L��D��K���;���u?��?-�+?,�= b�]�E�W���4��>�B�?���?%g*?�"S����=��Ӽ�Zr� ��>p��>d-�>���=SH=�!>�l�>���>�p��R��8���N�0/?�]F?Oݺ=�d����F����[ʾ��6>	���¹�_B~���f�Z��<W���r�
�sNþ�9}��þ������c���)��0�>�T�=�(>�->�c�<2^��G#<CY�<%�\=�8��TK��BѼH�K�DKq�HjŽ��!� =��>�) >v����z?�)Q?��>?e1?�'>�>������> ��Cs?��>׹�O���`��྾�'��.}ž̾��u����ù>O��7F>��R>
�>���<Jq>:�,�p=�E=���=YR�=0�=B��=���=��>U>I�x?��w�7y��4[8� ��� K?��>�E>T�M���*?n�=Is���w�����G��?���?e?�?�?uf�R�>b����6��=g�H�:.�>�Ǣ>�ꊽ���>��=�`㾼���s�ǽx��?�

@U�R?o��l6ǿ�|�>Y�>`[>[1V��E�"o�<m��=ޑ��E�>EA�i[�W=u��<�������_Mt�%��=�ɱ��ㄾ!�c�T >낽G	�=qb >悱>vO7=�DE=%��N<>1���y�>"F�>�Mh=W �<,���Q>�Y>�>{�e>��>&v?��1?��b?��>�Du��Aо�c��\-�>/��=��>��v=f;>G)�>%k4?s�B?|�K?*%�>���=�>�>�ǧ>��-�J)k�~x�U���OM�<��?N �?7�>��<��E��Y�:�?��ý�?�,4?��
?�>A�����_�02�H >�ͬ>"����s�u�j=m�F>��k���a���>ϟ�>J�>��R>4��>�Y�<��T=xr�>�U>�;�=қ	=�����`t=�/=��ѽ�%�	ؼ�1�<����yϽ<)�=�X��@�ȽRb?=� ;F/K=Ʊ�=���>(>��>ꁗ=����{/>s䕾�M���=�<��%:B���c�a�}�|�.��Q5���A>#�U>���n(��,�?�Y>�>>Ti�?�1u?�� >UP��lվ�,���e�N	T�i��=�>w">�{P;�\`�t�M�;Ӿ[/�>̆�>xj�>1�o>p�,���?���c=S�پm�8�4�>/~��䕼� �I_p�+!���퟿�(k�'��;.�B?�q���2�="~?1�K?q~�?���>g������@7>�^~���<t*���p��s�|1?X�)?YH�>N:��>G�#���̍�Y��>�b��>BU��������7Z�=�������>����}����%�9���aC����6�$(�>�>ZHN?�ѧ?K"ʽ�B���;G����B�-����>��b?�g�>- C?F�G?��&��%�Yƪ�������M?Ld�?�?(8>���=��4^�>�	?���?���?�qs?�#?��H�>�k�;Bh >�3��vx�=��>�=�8�=hW?�n
?A�
?�H���	�m�M���<^�u��<$n�=�e�>���>�Nr>���=��i=���=��[>u��>��>�d>O�>�g�>�W��x�_�<?<�)>�C�>��%?r#�>�3>��޽���������u�s-ƽ?Y��߽H,=���nJ����,�>����Ț?�fa>y����?�a�,
�`�|>�>��ֽ�t?��^>�BB>��>iw>�x>X��>r(>q.ӾQ�>���xv!��B��HR� �Ѿ̏y>�_'&����p[��+�I��~���r�w�i��%���8=��M�<R:�?F���h�k�c�)������L?�9�>��5?0���Y����>h��>���>5��؂��W����?���?���?�`>�}�> �E?�~�>T2
=y���8��,k�����H��+Y�zD��d��{)�S���O/?��q?:�N?ը�o�>��>?ɹ ������<�!�/�
��ܶ>2�>��m������u�q���ۉ�R[v>)�?f֍?�"?"񄾊�l�U�&>�$;?�1?�2t?�1?��;?n;��x$?�92>��?4?z`5?1�.?��
?2>���=̻́B,%=&���[E���Hͽ�ɽD;��v!2=7�x=֎��<>= ��<4�ռ� ռ �:����&�<#�:=���=m��=L�>�1]?K��>u�>)�8?����9�R��M�-?�)=
 ��9���_夾���lj�=��h?���?e5Y?��c>�~?��N@��Y!>��>�W!>#�N>�.�>��PD���=|>�>[�=X�T�������V�����<=�!>��?�A>�'�=V8�><d������.�>��k���	�����(�5���B��i8=�D?��\?" (?5�=����~>$Ci�GbF?��L?Z$;?�3�?�䟼�������G�J��*V�>�w/���&�:ͳ��­�=�!��<���<�H��j:�>��8�+��%B�Z���/��rr�����]>uP�2��x���mi=��=�*�x(�C����ि��??P�<y0��T��.n��+q>	�>b��>���6i#�I����+׫=�N�>��=݀T=
�Ⱦ��C�L�.���>h$@?�]T?i+�?�3��i\����D�W���6wG��h>=Qn1?E��>�Q�>;>����d~���_�ԍG��L9�BX�>G�>&�,Tt��T��j���T[��t>4P�>}C>��>9G?��4?�O?) 9?	<?���>*3P��?�K+&?���?Ef�=/�ҽ�cT��&9��wF����>B:)?�A��9�>;�?K#?g�&?\MQ?�}?Q/>�� �ϋ@���>���>6�W�UU��*
b>��J?��>c�X?ݝ�?�n=>��5�����N���>W�=_� >��2?�O#?E?K��>И�>뭡�~!�=���>�c?N0�?J�o?Zg�= ?�%2>���>��='��>���>?�UO?�s?��J?l��>;��<�E���:���@s���O�<�;<�H<g�y=���Y,t����؜�<9��;i���J���񼰡D��������;d�>c�s>���0>��ľ�n��7�@>]��W���͊��y:�K�=6��>]�?؊�>��#��9�=(��>]c�>����3(?��?�!?��;�b���ھ�K�]��>��A?I��=4�l��}����u���g=a�m?}^?֔W�+����\?�`?VM߾*�\a��r9��[�2JG?8�?<�����>m��?�,y?T�>êV��Tb�˗�@�^����N�=�t�>�!���k����>��:?�W�>;�&>Ts�=xYԾѻ~�&m��Ѡ?U�?"��?�#�?2oO>`�l���޿8N�rw��+&m?_��>]���Ĩ?�/I=�y;����6�������㧾���� �����q��U��c5�=V�?*�n?>�c?�mU?��"�%?e���V��jp�X�B�`8׾����H�i�9��fE��m���
�3���C�A�]�=��n�ڎG�u��?��&?�N$�7��>��r�4#꾵;۾��>�7��_��9e=���f��=�|=�[y��o:�W�����?/j�>|��>��6?V�l�q�=�<(.�>2�l!�+}V>�#�>Fr�>�{�>z�:��F�[��Ij��bJ��+h��dv>�c?5K?|vn??) �]V1�C��Y!���0������UD>k�>��>#4V�[���%���=�G�r��������/	�_�~=�1?� �>Z�>0�?��?����'����{�M{1�7��<�]�>�'i?l
�>��>yѽ�!�qL�>�Ld?���>? �>*��"�5��1W��t�=h<�>�@�>wc?]�>�M�%�J�[���5���4�9t=>�PY?wa���vV�H��>i�O?[�b<�l%��;i>���N�I`����6���>�w�>}�P=�
7>`3���x�S�v��m��O)?K?�撾�*�5~>($"?݁�>�-�>�0�?")�>qþ�G�Z�?��^?!BJ?_TA?XH�>��=N��v?Ƚ��&��,=,��>�Z>�"m=�}�=���q\�v���D=ny�=��μ�P����<������J<���<��3>g��6a8�o�����=�BzǾ�t����;&gv���U���.Gξ={̾����_����t���f�����Ͻ��?@��?�<�{}��Y胿��d�+&���>�.Ӿ9R�<` þ�˽� ���� ����z7�N}W����`�O%?�}����ƿ)q�� ׾�}?��?)4y?F4�B"#�p!9�l+>���<.'����A��ԫο<C��9a`?'x�>�,辙�����>A�{>�F>~v>���Tg���R<�`?�/?0��>	�t�.�ǿt���E~�<�t�?I�@�|A?Q�(�c��FV=���>��	?*�?>hR1�iI�U����T�>x<�?��?�zM=_�W�#�	��e?�<��F���ݻ��=�;�=ED=#����J>U�>t��LSA��?ܽ��4>څ>{"���p�^����<�]>��սW;��
\�?�n^�
�f�~.�����Z�>N�U?��>b�=*�'?C�H��Ͽ��X�Je?x��?�M�?/�'?����렟>�cܾ.QL?�\8?��>+�&�\Ou���=�+�ߓ�8�۾�U����=`�>�� >�k0�(����M��c���=<v���ɿ̛*�)���=S֊=N_��"�R%t�9ܿ��E��4����"ν=@��=�M>�>DTM>@�l>��d?�-�?]�>�O�<�D�K��������3�q�t���ް��I����������ྠ�����yG����2�>�ҕ=R�����-���^�)+H���*?k{>[�ľ{M���;�˾�T��_琼㷽%�;��2�l�k�՟?��B?}t�� W����?E��⻽#�V?�X��K�@i���C�=(�����=�W�>�ɜ=9-侂�5�)�U�_3?�H?]���a���>B+��}=�~7?���>I��=[N�>��%?l�(��e��Q�,>�c>jC�>Z�>�>T&���6�@�"?��[?�����/��|l>����-��1ƍ<��>UT�����K�B>L�,=,���)eA�.���~)=�`?��>��!�N��T�ƾ�.��F;>Ʃ�?Z��>DP?��w?N)?��W�ƾ�Fa��P��K>��{?SVE?�̾=t�-�&���^���}@?��H?	�>�J����U�!���׾�[3?o?i�2?Xg'������ ��� ���%?��v?=o^��s�������V��K�>�O�>]��>j�9��p�>��>?3#��F��N����W4�/Ğ?��@ۍ�?!,;<������=1?�W�>��O�� ƾ���~��[\q=� �>;����iv�Y���3,�]�8?1��?a��>����ެ����=vڕ��Z�?e�?�����8g<����l��n��z�<˫=��F"�Q��]�7��ƾ��
�ڪ��Sݿ�8��>Z@\V�1*�>)I8�26��SϿ���@[о�Pq���?��>��Ƚ���C�j�1Pu�8�G���H��������>,�>����rm��3(|�N�;�܄���^�>GG� ��>��S������8����<�n�>���>)��>�������S��?~���oοY�����[>X?JC�?�|�?s�?[<1Ar��{���'�e�F?��r? �Y?����[�xC9�-�j?7M��6P`�.�4��DE���T>�3?�W�>S�-�;�|= %>���>_f>N /��Ŀٶ�f������?ӆ�?uk����>��?x+?\h�y6��La��U�*�|!9��1A?w2>�{��J�!�*/=��Œ���
?/w0?ނ��#��{?׆�����%�\f;��K�>�J��ݹ:��D��	��Q_��ã�9���\��?0�@�c�?'n��i��h5?b¨>���X{�*A+>�֊> �(>�>of�=�`:��#��I@���=��?�g @��?t���џ�g��<�b}?���>Qw{?AVa>�?OZ���!����>@!=�2=%?t�\?�S�>��C=��u�8�7�!8���:��&�I���p>if?�#g?��E> �P�e���V1��v.��<��x���������n3�8�1>	=C>�y/>�ʔ�lk��e�
?�s���ʿ%n���6ؽv�?~ �==�?�0��s��d%̽n?��u>�\-�F��$1���n��?Y)�?��??<��/%��i&�=*O0>n��>���D�7�]�˽a�>E?׃��̓����W�0c�>n�?M� @�~�?9�V�G�?ē��R���.vt�$��@*���3�/O	?���8��>�7�>v�b=�Sr�@����co�*��>�*�?e�?�>��w?j�����=�M�<>�
=��?��?n�i�x�[���e>���>o�H�����kBо�q?��@��@ND?t߱�.Կ�����'��gJ����=}�=��M>����4�=�	o=��{�r����A)>U��>R�\>Se>
q_>ǎ$>�"">����-#��﬿�ʚ�m@��c�=�m��`���:�_���ٶ�e����Mk�&	½xŗ�z�7�ط:�����^O�=Ph_?��G?n5X?��?��ý��0�uU�O$�<�ؽYT>2l�>��T?�#E?t�$?s�=�8��L�O���۾$8��<��>�UF>�� ?�?�Q�>��!�*�s>�Z:>Gx�>rE�=U�սԞ�=��=n�3>���>vJ�>���>^9>۩>̣��~J��u�g�ts���νަ�?+ ��pMJ�~3���ꍾ�ķ���=��-?\> �EJп���A�G?����� �BW)�a�>��0?�6W?8c>𨰾��Z��>,�	���j��#>� �g�k��3)��5R>?Pc>�r>�Q3��s8�:O�0ݭ���y>`f5?Y���c�:���u�<�H�B޾��K>Ґ�>�[�v�� ���i�~� 1h�~�v=��9?�?R&���	��ӆv�W���OQS>�6[>Y/=n�={�K>�g��
ȽhbH�X�,=�1�=��_>�?߅G>�l�=Z˴>A:���̇���>A��>(�&>��D?��.?�=%<Ǫ����o�ѐ`���)>)��>��>�>AMa���=��>�ہ>�A��6����Z-�"�A���H>@�ʽ��a�Ңo���=�㛽�Z>��n=�?+�Nf�EuZ=,�?��.$���˾���(?��/?ۄ�=����D�z�������?0�@b[�?p=����2�|�?n��?��-:> �,?���>(�Ⱦ�%ҾP?jc�{,	���,��d����?M��?��*��8����j�G>�� ?�(����>�E�
���
��/t��=C^�>g�H?���c�$\A���?#?�+���ä�?�ȿ}�v��|�>^+�?S��?�kk�����!U?�K��>O��?l�X?�}l>�|پsMY�.�>hI@?��P?l�>As�̺$�=�?�ö?��?^	F>!�?��s?ޢ�>�(��c7�
o���ր�1]�=��;~S�>��.>*��92@���������{j����5f>�=Z��>����X־��=k���W����hݽ�ɹ>_�y>X�,>�E�>ӌ?���>s�>��x=�\��PZ��N�����K?���?����n�S]�<{�=�&_�*?�94?�Z��Ͼ���>��\?���?��Z?�X�>v���:��o쿿����%ٗ<�K>N�>�z�>[���8K>�վ�D�{a�>���>����}ھ��������?�>n!?|�>�F�=Í?�$?�vf>�(�>9�B����� �D�E��>���>-�?�;{?:{?,���4�S:����N�\�<R>�-z?��?i��>V���e���
�}��Hr��Ֆ��z�?��e?�Y߽�?)&�?��=?�7??bie>�"�ђԾ������>��!?�4���A��1&�����j?�e?���>�j����ֽ��ؼ^���l����?�\?�@&?����"a�]�¾��<��%� 
R��N<�|@�J�>�h>/r��ϴ=�%>�n�=H�l�t6�Kf<9v�=-d�>U�=I�6�$���G,?�&D�g郾
A�=��r��~D��>��L>������^?��<� �{�+��do��7VU����?��?Js�?���+�h��=?N�?�?�E�>)���f޾`w�Yw��kx�|Z�Pj>�>n�b���T���͟��d:��J�Ž��⽖н> ��>
3?��> �>�p�>�0n�F�C������ĺe�4�a.�-2��.㾨��}�e�g��cؾt�^���>�w����>)�?�GH>�>5��>c������> ��>���=c�>��7>?�>=�=}==�Z�=KR?�����'�"�辸���;2B?�pd?u2�>�i�9���2��)�?k��?kr�?Y8v>Oh�Q-+��n?BA�>+���q
?�T:=�8��+�<�W�����H/�����>A׽�:�	M�Kof��i
?x/?Q��0�̾5׽��bFn=/ȃ?l�%?c&��O�Pp�YpV��Q��c#��/n�@���i�$��Wp�mҏ��v���1����(�[�3=~J*?�ۈ?m\��5�qկ�Nk���=�bqh>���>���>1t�>�eS>tq��.1���]�H'������>�|?��h>^Q?��<?+�M?��U?�ދ>ڈ>E�ݾ�>m�=_�>c�?�C?�G6?ʶ-?�?6�,?��G>-�M�����վ�<?�S?|?�?jS?)
}��gS�|֡�Ҙ�=�8p�ܮ��/ۑ=��;͋��"��`��=TN{>�-?���+R8��l ���o>� 1?G��>�>�?��﯊���<�b�>Ĉ
?�]}>T:���u�0��A��>oE�?b���a�f=�� >\(�=>�����AN�=a�̻T�=�$]���	���n<��=�ɂ=Iɺ3%<Z@=<���<��)=�?T�?��:>��>*���"��Y��D��>"�[>J�>�p>�9��U��֦����b��/w>5ե?��?�3�<�3R>�K>>ڡ
�H�¾p@�������Ё=r�?$�3?��Y?/۶?-�??�\
?�܁>q�=/��d�k�t2�P��>�|,?�ُ>����'ʾc��3��?��?�a�Ui��J)�(�¾��̽�w>�?.�a}�u�����C���k���Uʗ����?���?B�;��f7��辭�������C?af�>A��>��>�'*��h�����:>t��>��Q?au�>��R?�rv?TxY?�	X>0:�;}��W���9l��x&>5v@?��?S��?�u?���>�n>6�(����`��e�WIϽ��}��=[�>.��>S;�>��>���=�ʽ����b�I����=(�i>���>�U�>W�>�h>׈��G?�n�>e�������������nv+�W�u?�͏?�,?��=�I���F�������>Pާ?���?�|+?�QS����=q?������w�q���>6H�>H�>�-�=�e=��#>O�>s��>�8��a�m�8���P�n?^kF?ߜ�= [����B���Ǿ���=v�>�M>+�˾R�⽩;���a�k���곾q����k��ཾ�Y;�����i��w��	�>Ҍ����=��>�-->bY��䓰��O<Z1�=��<���D����=@.��G�����&�ô����d%)>��`>��¾\�v?V�L?\51?S9?��P>
�*>�5`�qސ><���?�a>���p�����E��ɩ�O*��-�ξkϾ-�l��렾��=�lx���>�e2>���=@�6��>�%v=T�[=6{�;�=�Q�=ă�=I�=���=^>
��=hi�?'L��ⵥ�kJ������AO?@R�>K4�;��齵N?	��=G��#��(�0�?}�@-'�?V?o\O����>����%B��W<������=�̴=�f=�����U�ZU����(c3�{~�?��@x�_?U.���Eڿ�s�>��4>q�>��R���1�-�Y��_�Ig[�)-!?�W;�'̾啄>˛�=�n߾�Uƾ�+*=��4>��Y=O�sr\��Ú=��~��K:=	bs=4N�>�C>���=<���̷=�,F=dX�=־O>TH���S9��.��1=?2�=�c>N�&>V��>��?G�0?�Kd?3m�>�rn��ξ�����>���=棰>ݑ�=%�A>:շ>��7?a�D?��K?֨�>��=�:�>^��>��,��ym�6m澎Q����<X��?���?{�>�_<�B�h���c>��ǽ�^?H�1?��?˹�>�U����9Y&���.�#����y4��+=�mr��QU�O���Hm�2�㽰�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�='ጻ���<� �����="�����<�vż�����u&�;�+�2�����;x��;C�]<i��;B �=6\�>!%4>V��>*N�=:�����G>\.��U}S�bЈ="氾NE�`�\�NPy���'��Z#��Y*>�&A>��V�4/��m�?��V>�&*>K��?� y?Yr)>��ŽB(ƾz��8�O��X\���X=?,�=X�L��8���a���J��`ݾ-�>� �>��>��m>,�wO?���x=W���H5��G�>k���e��X�]�p�9-����i�F�<�?�D?�>��;�=g<~?J?4��?9�>�����nؾ{�/>Թ��M2=R��cyq������?m�&?�O�> s�yD��A��^�ֽ��>��ֽ��c�R֐�^~	��Cd<��Ͼ=�>��Ⱦ:�徜:/�����39��$(��ؽ~J�>��=?�?�Xb�����P�8�X�:��;V��y�>�Qs?`�>&$+?O�*?~�]��������۬�^[?Z��?�E�?�1�=Ɏ�=E����^�>u*	?���?֫�?�s?�`?�.2�>�;4� >�阽O��=��>�՜=�b�=�T?~
?��
?<k��G�	�f��e��,^�uj�<���=xh�>t�>,�r>r��=�h=�O�=��[>XǞ>Wɏ>�e>�>!N�>M����[��X3?�T>���>\�$?@�>�Wh='�(�����~��]A�"�D�YȽ3L����E=�Lp�m6�<ы{�?x�>V4��ї�?�S`>V���?�C�	���Yh>�c~>����%(�>~�7>��,>��>X�>�f=>	�>��A>2�޾a<>Ƀ�f;��߾�l�����Q>8A^��b�@�	w^<�KQ��e���(�'������:�(��n)>��?>��=%�D���fq����:>�$�>}J?u}���Q�R-�=b�:?|�>&��)D����z˾ݑ�?���?9�d>ph�>+�Y?��?�x;��%7���V�:�s�'hA��c�Ca�HT��〿��7����@^?��w?k/A?i�<4�~>��?�=(�h����|>��0���9��a=>_�>^ɧ��V���ؾƾ��C�:>}�m?��?�?f�T��^����`>U�F?��7?��?R�<?��C?2�޾ncc?�"
>�H?�)?�7?G?F��>R�>��i>w���h;��2��x0��N�"��e �w��-T>,h�>l�>Q�>�\��}	��~��<Żl6�S�Ļ���<RL<<\�=q[>���> �]?�L�>皆>��7?d���w8�Ʈ�v+/?��9=������iɢ�����>C�j?h �?�dZ?xad>B�A��	C�h>\X�>.s&>�\>	e�>A|ｎ�E���=�L>�Y>�ĥ=�_M�ρ�#�	������<('>��?yԊ���=�R>�N��u�Ծb��>�ؼ�׹(��a�a�X�4\;��Xx=���>�%X?O�(?ˣ�<�i�,�:>��z�v�4?m{]?01?o��?,&=�Ծ8��/���'�	ʈ>@�����8�e̶��?��=�-����rc�=�4��؟��;e>���P徬pi��F�`��r�1=/���8\=K��?׾�O���H�=���=�Ǿ��"�hȖ�@-��`2I?u�==�E���K?��W���<>c.�>]��>^�<�Ǚ�Jw?�E��H[�=`��>�4>YO+��*�v�F������|>�MR?v|a?�i�?�M�
���87�D پ��T����H?J�?�v�>�N>O��d�־����oS�e8����>if�>�>�'m���؎��T��+��R�?WS�>��1?љ|?NI?��O??@p�>�o�>N�M�
L���A&?D��?,�=@�Խ��T�� 9��F�{��>��)?��B� ��>|�?ڽ?g�&?��Q?�?n�>� �D@�W��>oY�>M�W��b����_>��J?��>�;Y?Qԃ?,�=>��5��颾3ϩ�hW�=�>U�2?%6#?ί?���>|��>L�����=ƞ�>�c?�0�?"�o?���=<�?�:2>M��>&��=���>c��>�?SXO?=�s?��J?��>T��<�7���8��"Ds���O��ǂ;iuH<��y=��3t��J�>��<��;�g��;I������D�-������;��>J�I>dy^�i�0>�;M|��&`>�����ؾBq����\�DW�=t��>T?v�>��ӽ\�<��>t1�>4$!� `%?�� ?�S?Ы�;Id�gj��3�9��>�:?��\=:Gp�Ŭ������pɪ;̖`?�O?�;X�1V��b?�]?�g��=�^�þ϶b�N����O?(�
?�G�3�>��~?3�q?��>o�e�0:n���Db�k�j�Ѷ=r�>EX�4�d��?�>w�7?�N�>g�b>$�=u۾��w��q���?{�?��?���?*+*>f�n�[4���Iō��g?�g�>-��	"?���<c�ľI����T����侌⡾�R���ژ�M7�����"�� Kｻ��=��?ft?�Hm?��[?�����e�#�W�<�}���J��Y�l��@��I���H�K�k�+#	�mZ˾QN��u�=�`���8�;�?!�'?�f����>,�\���վV�վ0�>�p��X������=X����=c!�=��C|_��۞�A�?��>���>5�6?Nm��?��Q#�<	;���ؾ��d>ނ�>(��>f��>�[����2��VŽ�c���޽�^��yt>�d?]8L?g�m?�-�g�0�	ꁿ<�#�V3#�ᜢ��$O>ϊ>�ً>�R�(��&�|m<�M�r��������Vy	����=�2?�>N��>U�?�?Œ	�<���|~��2��;E<쀺> �g?���>���>Σͽ����ע>� e?|ߟ>_"��F0��������N�ؽ�Fk>���>fʊ>�P�=<e����h��|��)E���9�fn�=:p?#&�2|��r��=:�]?H�=o�=*�>#��:�A�+��o{��j:>�)�>in%>�Á=@⓾U;�<��_��O)?NK?�璾(�*��6~>�$"?���>�-�>�0�?L*�>�qþ��E���?��^?�AJ?!TA?�H�>?�="��0=Ƚ��&�+�,=X��>^�Z>�m=,��=m��Qq\�Nx���D=�v�=�μ�P����<փ��h�J<O��<��3>�TԿ��A�	�Ӿ���L�[��s����B�n�D���"�������!h���ݽ��"<���4�O��C�}������?�5�?�/P��|�D�����r���-����>c�e��\�=%�ܾ�z�4%�����|�׾Ρ7��R�GkO�����'?$���˽ǿ�L9ܾJ! ?A ?;�y?����"��8�9� >K9�<"1��Z�뾫�����οq���x�^?c��>���-�����> ��> �X>Iq>����瞾�*�<Z�?M�-?��>��r�ٕɿʊ��ۿ�<���?��@|A?7�(����V=o��>K�	?��?>�P1�DJ�*���O�>);�?l��?|M=>�W�8�	�R{e?^'<�F���ݻ
#�=I�=XU=����J>�S�>A���OA��2ܽ��4>[م>_�"����A�^�Ԙ�<��]>��ս]1�� ݄?}k\��f��/��C���^>��T?�j�>�T�=�G,?�"H��uϿ`\�!]a?e:�?��?|�(?���uH�>��ܾcM?�D6?.�>$v&���t��Y�=��༩�Ի؋�\V�ӽ�=�C�>��>.-�p��.iO�E���/��=[ � �Ŀ�r%����ռe=\����1�Xm#���C�\���;BF������=>�>Zt/>Ba�>~.�>=�K>�>^?�|?��>��<z���1ɓ��M��~�x�]���w���_��:������\;�a��'�6����m�� =���=0/R�b����q ��b�l�F���.?�}#>z�ʾw�M�FS%<O�ʾn���ZK���7���v̾o�1�8�m�\��?E�A?�󅿥�V�����������W?Z�����\𬾡��=$����=�Μ>C�=M��~3�͙S��\0?ur?�W��Ӿ���W>W[�l��<9&.?��?ä�<�>
�%?��5�P���dF>�->��>��>�>�:��?ܽ�9 ?�'T?�����G�����>�F���(����<�}�=��0����m�Y>�Ó<IN��%G������s<�(W?��>1�)����ꐾb:%��<=h�x?��?e/�>ϻk?A�B?��<����R�S�
 �lx{=�3X?��h?]`>�`���ϾY����N5?�e?��M>�1h�̺龂2/����e?��n?�.?��r[}�p"��D.��56?��v?s^�ws�����O�V�d=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?p�;<��Q��=�;?k\�>�O��>ƾ�z������:�q=�"�>���ev����R,�f�8?ݠ�?���>���������=�ؕ�[�?~�?n����Cg<����l�cn��2y�<}̫=��1G"����7���ƾ��
�����ٿ��>�Y@T�1*�>�H8��5�uSϿ��ZоWNq��?���>��Ƚٜ����j��Ou�}�G���H������R�>��)>���m0��Tz��?�c�<q�?�IX�ؠ�>JN�4پd����3���>1��>���>�y�<����^��?m���ӿ�ʕ��.�X5c?���?!C�?3�,?1�=�f���Ь�)#X�>lN?l�?�̂?��?=�sx�gt�&�j?�_��tU`��4�uHE��U>�"3?�B�>W�-�I�|=�>���>7g>�#/�u�Ŀ�ٶ�>���X��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�F0=�YҒ���
?R~0?{�g.�cSz?0�L�܃��.9��M��?.���=I�R>d���^H��i���YE��`�?k�@�4�?'̽f�2�'xA?9�>Lj��c��+�<�!�>��>A��=6dv�����Q*����!>�r�?���?�_?�*��ᩘ����=+�r?�˷>,��?���=��>S��=.|��G/���D7>��>��L�@k?=M?f��>�ا=T5H� �,��{?��fK���t	E�F�>�:e?�M?��h>�����%���������J���9���K���Z�vc׽�Z7>��<>=�!>y�S�e�Ծ��?Hp�6�ؿ�i��p'��54?%��>�?����t�����;_?Iz�>�6��+���%���B�]��?�G�?>�?��׾�R̼�>8�>�I�>1�Խx���W�����7>1�B?[��D��q�o�{�>���?	�@�ծ?gi�'�?��޾�؃�a)w�؉�/.{�ޗ�=��??�Y�<-Y>�6�>�7=Ox�g憎a�l��>z��?q|�?l��>�Oq?EXm��X�>��<�(>�rf?^c?���=�wþM�~>f�>,�#����a�߾ɫ}?�@C
@�^_?0���7�ƿ��ն���Q���=��>��U>ʽݴ=�:�^�n=}k>�^>'g�>Xk>��>�K>��->��ļK{{�k�#��E��)N���C�ϒݾ>%�������Ͼr3��v������g������c�"b��?9��#�_��^��=r	B?vp?��a?#?�%=zt5>x$�"X�����K>�$�>��+?:�8? �?��<nľE'���������Љ���?�W�>0k>K�?zv�>%z�=8Up>���=H �=��="�J�"uX��ӓ= m>>I=�>OY�>s��>:@<>P�>�δ�j2���h��w��5̽��?V�����J�,2���;������V�=�].?i>��>п�󭿛1H?1 �� *���+���>��0?�cW?��>���	U��4>\��I�j��m>�/ ��sl���)��Q>�e?tXn>Ėb>��'��1�B�A�#ʩ��ۊ>��*?a�_7��t���Q��P˾EA5>��>�X,<%�*�p�@�p��{�֦C=�?9?g�?�{伅���ai��kz��E|>xU>��A=~��= �>�����Y⽹QI�3�<kh�=�@4>�?>�}>�N>c��>(�ξp��q��>�ݤ>�L�>��*?��??Ś=�7�Ԥ�鲇���L>�[�>>��>(M=e^��og=i/?gZ�>���<4է���佛/+��I�=�l�􄎾�vֽ/d��V�2�{�>sR=�Y��5&��[ o��)�?v��*6z�j�����}���T?�L?��M>�Q�$�C�!;�������F�?V�@��?�+���b3�~�>���?�4��ߏ=P�?��>��ܾ�M��G�>�߰�R.������M�f�?��?E��=z0����j��h= �-?� ƾK9�>����L��.����u��#=��>RH?�J����L�S�>��?
?��?���柤���ȿ�yv����>g�?Z�?عm�V6����?����>���?�QY?��i>ՠ۾��Z���>h�@?�Q?��>+G���'��?ɷ�?h��?
'5>$�?y>g?y�>S��=�92�����H����uq=	P�\S>
|7>Q$��~�E��"���(��w�c�{�ǢV>��\=\��>N�������q�����J���s<���>��@>4�]>]��>��>'��>��n>7�Z=н;�Z]��T�{�K?���?���2n��O�<.��=��^��&?ZI4?Gk[��Ͼlը>�\?a?�[?d�>H��Q>��:迿@~��R��<��K>&4�>�H�>�$���FK>��Ծ�4D�bp�>�ϗ>�����?ھ-���V��2B�>�e!?}��>hҮ=h�?k�$?c�x>�½>}!C��K��vCA�%L�>ʏ�>j�?��?;�?D���l2�����0����Y��K>�u?/�?�b�>1��o朿4D�\$&��Ƿ��|?b�h? �н�R?*1�?�C?c@?M�h>�9�Q�۾%-ý7�~>i!?Y���@�z�%����c�?ԩ?DU�>�S���ؽ�
�9�N��u�?+[?��%?n���"b������7�<����u�Zr@<X�(��>>�~����= x>y�=To��q@�(��:'T�=���>��=_`>�\��,?l��������=��r��E�3�~>��O>����]?<8���z�7���O��ZbW���?�r�?�N�?�}���h�Om<?��?A]?��>���zݾ�D྘y��e{�"y���>%��>��^�j�%.��{��z9����ƽ�rϽlm�>k�>�u�>��?!�R>�Y>ֻ���A?���־���P�}I�9%��&����W��j��y�-�}���v���ө>�2f>]�>d�?6ik>��>O��>�Ž�V�>��>.�k>Y��>>:4Z>-v�=#�=5�=�ܥU?b�¾�;��B�u����;?��b?#��>8*������3�.	?�Қ?Ʀ�?���>�hY�c.*�B&?L?���$?�.�=v�<�>=�wɾW.L������̄��f�>���Ou9�\zO��ϖ��f�>ƙ?(�
���;\X�'�����=���?��!?�^'���O��6r���W��	P�F�¼޻m�����p$��Cp�4������E]���$��n=`,?堉?xp��Y��mz��E\i��>?��o>x��>8d�>�R�>��>>
�^�3�� _�,�'�Ǻ��y��>��{?�=�>�qJ?i=?xMP?sfL?�(�>5Ϧ>r���Nl�>0�q<H��>���>�9?�G-?�-?��?�{*?V?Z>Y�	�r_���\ؾq?�?�?{�?'?�����Iʽ�2���6�������ש�=Y.�<g�ԽKS~��S=$UV>�8 ?����L�2� �����>ae+?K�\>D�E>�Φ�x�s� TC��$�>���>�D>���
q��h)�S��>�`?��;�y��=�q>�uR>o��=�����=�y�=�{>�ى���==��=��==���-΀<��=��=M�=�@��?uA0?'��>��>��ž�H6��ꗾNR�>S��> _�>G��>,þ�-��j�����X��%_>^��?r$�?��m��7>.	>����.���`�������2�>�	)?0$?�Э?��N?��?H=(>�
�����Pօ��K��P��>\d,?Sِ>���|�ʾ�Ԩ��3���?�?��a�-��E%)�����H�ʽGd>L�.�Gz}��ѯ�רC�"�废��f򘽃��?��?F>�d7��a��ʘ�2/���vC?p�>�Z�>��> *�<h����:>2e�>�9Q?�1�>_\b?u?>�M?. �>Y�=�����~��]@�=O*�>�q?}.�?R�?�`]?��>�t=�!ؽe#�S$/�_���	�ڽЪ �>�l�&H�>�|�>د?�R�=�l�|FH���<��{�-�>t�>��>�>���>mM>F����F?��>�ޱ�P	�+���R䆾l��xv?��?�/?)=î��G�� ��E�>t�?��?�.1?�zT�z�=�R}��þ�w��Ӵ>)=�>��>�;�=r^�=��*>���>Ǒ�>�	�"f��(9���J��6?�7I?/z�=��ǿ�!��O���3~9�:�Z<v� ��W��+7� ���]Ǽ�f���
߽�.��}�䊾c������D���S�ھ4��>��/=29F=3~�<84Ļ�彭k`�O =�@�=��>do��?j��j2���</ט�- �<�R�<е�<c�=|q��˛q?$2?��?��l?V�%>�`;��
���x>�a�`�>$m>t�Խ�ؾ(ڗ�������跾�*оG���u��M{>A{o��M^=�p=$2�=7?�;��>*�;BC�=9����3k<)I=��C=��=�"�=?�>��B>$�~?�j�#���J��K;�� ?�?��>��*���.?�>�=t���P������z�?�&@���?��>�(��TM�>�:��c9(�+�����t	?ѱ>`�Z��9 ?j���	{�����F����?`@�hn?&���O�Կ��>h5>�>!�Q���2�D@��7V��e�Զ?a<�X˾p�m>=<�=�r޾�Aƾ�P�<!">Ƚ�<�o�T0X�@n�=�����SW=�$�=yY�>}�=>�C�=Nᬽ4��=|�/=Q-�=�\T>԰t�v-*��6��)`=�.�=��g>)�>(�>�?�C?i�c?Ǿ�>��\��l��1���Qn>Ǡ>�@�>*�S=+�>g�>�+?r�A?1�K?���>�ѣ=�^�>��>�c1���^�$k�O�ξ�Y����?ݾ�?}-�>|��=��c��-�xN@�!���\?��U?�--?Ӿ�>͆����ceP�W��֮m�+hw>t�[={ Ծ�CQ>脿=ŵ��"M�x^><�>g�>�
>�\>���=�UP�-�>\`>�M�`L�M+ϼ�/���{�=�l5=�hO��dN=�_�`a=04�|r��s=9�==8f=���=P>bc�=e&�>HN>]Y�>!`=m+Ͼ�{">ɰb���;��x=�O���d8���h�Y�{��J1��0��,v>QLb>�qϽ�����L�>�V�>��n>bb�?�i?
�2>����6������ǃ��ہ���M=0~>&�!�(�6�mP�JRK��;���>�-�>d.�>�m>o,��E?�I6u=v&�5�ȟ�>�ŋ�����.��0q�h2��<џ���h�>颺YAD?�<��_�=�*~?��I?ӏ?�Y�>��JؾP3/>����	=]���q��3����?��&?��>]쾚�D�d�����;r��>�7_�i�#������	*���P=������\>r�������t+��*���ې��r3���X�g��>��I?$�?��3�pɅ��e5����R�Ὢ��>Ϣ�?7�>K�?��?��]����tz�{�u>�P?L[�?/B�?�T>l��=����'N�>U$	?*��?��??ys?@_?��X�>���;K� >#����Z�=�>^B�=�=[?(
?��
?]+��R�	���'��7`^����<Y�=���>cl�>6�r>��=k�g=�[�=9�[>�О>y�>�e>��>�_�>���P�%�'?H��=�.�>6K2?
��>�!c=�����٭<O�W��L?��'�.���}ݽ���<�/5��0=?�ּۜ�>�RƿV:�?�GU>]t��8?��6���V>`�T>��޽�B�>KD>��x>X�>X��>��>ܢ�>�2+>�ؾ��O>�^�S��o)�V�8���� H�=�nj�$c]=�,�r*]��=|��վ����_�x��fu��!��Xv>ͩ�?R��=��S��
J�+Գ<J��>�>>\:?^(��J�8#��2�>�>&>U` ��Ś�4o��.O��I�r?>��?qq>�a�>��g?�?��c�M�(�T>�<�c�=k:���D��E\�����p|��h��絽Q�[?˓y?�J?8�=��>�ց?o�.�'؊���V>ȍ=��`7���>	��>IHf�:���㾸i��C����=�fh?�ʕ?��;?+q�>�m�V9'>+�:?��1?�Qt?�1?͆;?���h�$?Ј3>lK?Qv?�K5?��.?C�
?��1>V��=:����&=tC����o?ѽ�Cʽ�J򼀰4=/�{=7�a���<�p=�t�<_��/vڼaX;xš�e�<��9=�=LA�=7�>��[?�?�2�>h�&?S��1&���r���'?k�*;@��2_���Ҿi����n=T?!Ŭ?rP?>��M�W�1��+!>sթ>�f>�5>���>ٟ)�{�x�͓X=�r�=GF�=��9=�e��ƄU����)���X�<|�A>k7?4V+>q�ؼkk�=�̦�ѯw����>/N�c�,�`���H�h�;��9<��>��E?�0?kŽn;�#���f��?�|?�@$?��u?�&=�췾����6#��ڜ��L>6�@�`�?���������"�ˢʽ|��<+���٠��\b>����o޾�n��J�H���M=����U=k�־9���=#1
>(���5� �T���ժ��$J?whj=us��+[U��i����>ƫ�>�֮>}:���v���@�.����=��>��:>I������(xG�4�Oa�>�IE?�p_?dń?�ׂ�D�r�:QB�k��w+���	�^�?Z*�>�t?��>>�U�=૱�ϴ�X'd��rE����>9��>	���G�����A����I&�8�>>Z?b�&>��?+/T?,�
?_R_?�)?��?��>ϖ�������J&?�w�?���=�Խ tU��9���E��q�>J0)?��B�Y�>X8?�`?Q�&?ʇQ?��?&b>Pb �oR@�Z��>Y��>�X��Z��$�`>��J?䜳>�mY?���?"�<>�75��t���������=�J>��2?�v#?7�?��>/��>������=ڥ�>	c?�.�?j�o?���=��?�*2>���>,�=8��>v��>�
?TUO?|�s?��J?/��>t��<�1���+��PBs�Q!O����;5.H<��y=̌��4t��W���<U�;8T���N�����r�D�)7�����;o_�>W�s>q����0>!�ľ,P����@>���PQ���ۊ�o�:�jַ=م�>��?u��>�V#����=���>�H�>v���6(?T�?�?=�!;��b�{�ھq�K���>XB?���=��l�$���L�u�w�g=��m?�^?X�W��$��#ca?�`?���e7��k�� �o��$���lJ?2t?���&/�>�?�?��u?N�>$u�x^p�Yx��:
d�k�`� 7�=ve�>���d���>��9?j��>/>�=J�ؾ]�r������?�7�?�a�?�l�?7>�Ao���g���ɔ��\<?Jۮ>(�U�"?~�����`~����t� ����4(���+O�8����A��A��w�սdy�=hL?9J�?vl?#EM?����Zv�)^�Tr�_�B����L�&��D��K�x�K�I{�������:B.��4�=OkW��^E��t�?��?�h�S� ?|M�@
�q���>;V�_�XT_=�ް�2�=�-�= :Q��/�2�վ:~)?��>-��>�2P?.I��	�C��M�+�.��8>�_�>&�:>N��>+�?<'�4��=a4���5���.���Mp>�o?/�E?�`?�J�<��&��ώ�;�@��D=D�;���>�o�>/�?`���Ps�F�9��<��兿����u�����_��=ʥ-?��[>�>"��?�|�>�B!�j��F+�P��5�����>kjY?P�>�|>iʮ��G,���>�+s?K�>�d�>��c���-�u��2P`��Z?v��>��??��>3����Z��q���猿35�� =Bb?�*���w6�q�s>b^.?���=sc�=��>������1��Ⱦ��8��%>S�.?��0>�P>��Ǿk����~��b��P)?�K?�蒾h�*�u4~>p$"?���>S.�>W1�?z*�>qþ�ME���? �^?3BJ?yTA?�J�>��=S��N=Ƚ�&��,=쇇>}�Z>�m=�=K���r\��w���D=�t�=8�μ�P��^�<ʈ����J<��<��3>�Uٿ�wK��ܾS��R+Ѿ��y������Ω��P��xǾ&�������D ��g�m��k��~�Jք��*[��+�?��?Ppi�֧��d���#*��0��K�>�e��æ�����z�������#�þ2)��M�<U��{O�M�'?�����ǿ򰡿�:ܾ2! ?�A ?5�y?��6�"���8�� >5C�<-����뾭����ο=�����^?���>��/��l��>ץ�>�X>�Hq>����螾l1�<��?8�-?��>̎r�0�ɿb����¤<���?0�@}A?��(����9V=s��>�	?g�?>�R1�nI������T�>6<�?���?tM=l�W���	�J�e?�<��F�s�ݻ��=.=�=JL=��:�J>�U�>Ӄ��SA��@ܽ��4>�م>]|"����с^�·�<"�]>�ս�:��Q�?�K`�`T���yL����<��x?%�>`��=��?�:R���ѿ��H��=�?�@ru�??6Rھk�>N�ľ�W2?|�L?���>;y���q��c	=����)������\�_�(%>[?=��>j�ֽ�����^r�uș>�� ���Ϳ�<?���(��[�>/�*>������=�T}ν�Q= 0��qkL���� �N>#�	>�	>�>E�>��J>��[?�9f?pz�>̹Z>�2��Fɾ�N�~u��a�[�l?v����PUc��վ}������	�����9׾�M��� =���=�6R������� ��b�Z�F�}�.?�v$>��ʾ��M�1�-<�pʾ����X넼�㥽�-̾r�1�G!n�`͟?~�A?������V���YR�\���%�W?yO�K��ꬾ���=������=�$�>X��==��I 3�q~S�00?�d?	]����p�ݜ�=�� �b��<�6?/��>�C����>�q?Om=�(�!�b8>(�5>�4�>%:�>O�=�r�����o� ?�Cc?�M����� �>+]Ծ啈�8`/=1�=��H���E=�JU>��<����j�,�CN��v�=�%W?ݣ�>��)�����w������4==>�x?!�?��>�}k?�B?�_�<�y����S��A!x=(�W?�i?#�>���\�Ͼ�F����5?��e?��N>(�h�6���.��^��?@�n?�[?�����s}�������v6?��x?H]O�������Ġ_����>\X�>vI�>�Y-����>�:-?��ҽT���9�ÿ0�&���?�*@���?�����1'<Ϫ3<l�?'��>����f��Oh=����|�=���>��]��4��no��7���dS?�Y�?�?������[��=̅��Q�?�'�?�i��>>_<���o�k��3����<J�=�#�=�#�5����7���ƾ��
������#��,��>vG@ܦ�O��>8��YϿ�텿�Ͼ�p�S�?C#�>zYȽ����9�j�F*u���G���H�5���lp�>��>ض��︑�e�{�v;�����F�>[Q
���>�T�J`��cƟ��D6<�>���>Yǆ>g��������?q����Iο����]�7�X?�M�?���?��?\2<�Jv�{�*u(�VG?yQs?��Y?N�!�\���7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�b�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.��_`?��a�@Lp�\�,�,��>%��X/T���̼�	��te������{��ɭ?���?��?�����"��
%?I$�>l����w��h+=��>��>v�K>�u�t�d>��7X<�U�>��?=�?D�?�F���Ǧ�[>g�?���>��?��=.��>��=h�J->���!>[��=q8�^�?��M?�"�>U��=�}9�>3/��XF�QnR�5���C�ب�>Эa?*qL?k#b>ۖ���<*��	!��ν�	2�m���i@��u.��^޽�5>�[>>h�>�+D���Ҿ�8?G>��4�ѿ�ힿ̰	��/?4"'>H��>_待��cE��4O?��Y>������[���CsĽ5ު?�X�?�?ǻܾ��"� >���>�'�>?�������&\��j>>z3?g��Ӻ����i�>�>���?�@��?�k�`5?g����R����Ab���=���z?�Q��O-�>[J�>8^>/.j������g��;�>)u�?C��?�O�>	
n?�j|���-��\>
�6>��}?} ?X<�=�1꾥�&�f��>������{����w?M�@=�@'zC?�N���޿����W���K���E>稣=�O>�T�s�=$�;L0��1�=qp�>V�>��<>�0>�i>��=FA�=��V}�j��CB����5�̘�-%����߾KG-� ��T)����|��`Ӻc��YY��)��Lq����ߝ=j�G? R?T�]?���>�ʽ��=@��������6�=�f�>�,?��6?5�?¸�<*���on��7�����į��f�>��R>���>4�>sL�>F���DKa>lo>>wKK>���=��l��e<%�I=�9*>=�>n� ?b۳>�C<>��>Fϴ��1��k�h��
w�p̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��t�T�4:>9����j�5`>�+ �~l���)��%Q>wl?�[>���>g1���1���D�0O���Cy>��*?�^ݾ>h���w�~gM�'�ھh�<>���>�נ;N���ї�|ŀ�r����"=O/?>v�>{���y���Z���������b>a]>W�<�=��">��G��� �j�a�{:1=���=��O>7�?\�?>]'�=A�>���Нr����>��c>W�>�}#?��%?���:�����J�Gf>^��>��>j�$>�\���='`�>='�>Q��<�=��׽@o��T�?>|�ν#���΂|�	3�=i�&���=��<3v%���q�I{�=V�~?J��Z㈿$��n���jD?�+?� �=�3F<Ӄ"�+ ���J��1�?��@�m�?�	���V�_�?A�?���ʾ�=��>.ث>�ξ7�L�9�?"ƽ�ˢ��	��(#�CS�?i�?��/�zʋ�l�7>�]%?��Ӿ��>\�s<��"��8�u�1�!==+�>�H?v��u�O��d>��j
?��?|򾌱��R�ȿ�qv�:�>|�?i�?��m�%5��@,@�)�>^��?�-Y?��i>�#۾�.Y���>�@?�Q?��>��o�&� !?S¶?��?�O>�O�?�<r?m/�>O�[���1�����ψ��=_��<
��>u>+��QF��S���(����i�ǩ��\t>�S=a�>�)ὧ�¾�c�=
wf�����F!��?3�>r�>�
L>͚�>�;?���>Nn�>��<.����s��g���o�K?���?���2n��O�<���=�^��&?HI4?t[���Ͼ\ը>̺\?[?�[?d�>B��Q>��B迿O~��ҩ�<[�K>4�>�H�>G%��<FK>��Ծ�4D�Op�>�ϗ>l����?ھ�,���\��B�>�e!?���>YҮ=�?M�4?�ز>^�?�~.��ؙ���c����>�'?k?<Ԃ?d�)?�)��(�A�����S���f�L�=Ѓ?�?��>��x��v��ܼ�=M��tɾ�p?�Ɂ?
d�>ڰ ?.~�?��n?��?���=?���}���-���IZ>��!?�I�A��K&��rz?O?
��>p���ֽU�ּ���~��N�?9'\?�?&?����-a�aþ���<�_#��U�d��;bD��>�>����ݛ�=Z>�ʰ=�Lm�!M6���f<2U�=Ox�>��=�+7��s����,?��!=��q�Ժ�=|u�Y�G��d>�0�>(���i�>?�C���Mp�Ǫ��"���Ps�U��?�R�? �?� ���`�2�*?�t�?#�1?��>�ᒾ>Ҿ%J�����υe�K��@�=g�?��Ἃ�ݾg����\������ML��r�
�b��>�r�>B?��>�
>���>CQ��#x*�N�����8�]����-��p�W�x����R?�]"�)R���A
�>���U��>	?�'>��#>:��>��=.&l>���>�9>,��>;�/>�3�=�/Y=hͺ������KR?����$�'����²��g3B?�qd?S1�>wi�<��������?���?Ts�?=v>h��,+��n?�>�>H��Wq
?yT:=9�;�<V��y��3���1��>E׽� :��M�Enf�wj
?�/?����̾�;׽8ż�0>�=�!s?��?�q�-P�(bo�ɺU�*�@�ߥi�2���s��$��>_�Ո������:!����
��F>+..?�ה? �˾����羇�j�s�(�:��>1��>��{>P�>�{�>�����=��Df�60�C}v��J�>��?���>�:I?\�;?�QQ?4=K?��><��>(�����>��%;4P�>c!�>|�8?�,?�#/?f�??�+?��c>�Y����	ؾn?;�?V�?q�?_�?�և���½�y������x�E����?�=�A�<�]۽L��,�J=�MV>�T?���8�����4k>U7?և�>���>/��&,��z��<��>{�
?QJ�>@ �q~r��c�IQ�>���?E ��u=�)>:��=][����кMd�=�����ܐ==B��h�;��<�y�=���=��t�����S�:,��; ��<IH?~?��}>��>�뎾�����微م>�>@P�<�{�>�Kɾ�I��V���:\Y��:{> (�?ra�?LEh<���=�{>��=�+˅����!q������m�>�T?|�U?��?�:?�f1?D�;����u��i�����˾m�?�!,?̊�>|��q�ʾ��ۉ3��?^[?�<a�����;)��¾��Խ�>q[/�
/~����;D��م�����~��7��?濝?�A�*�6��x�ο��F\��G�C?�!�>@Y�>��>@�)���g��%��1;>���>>R?6��>UQ?�y?�Z[?�Ad>�c5��T������z�":U�G>�E?uA�?��?�t?�=�>��=`�<����DU���U����H�}�x�=T>�ϕ>�'�>@�>���=�������g@�܄�=�?g><�>ΐ�>���>��>�f<'�M?�1�>Xٲ�Y\Ծ�ľ� ��%=�/�?���?�R�>�6f�3��H�q�=�׾^X�>8��?���?^�Y?ڶ��U1�=zf=�[������>	�>�9�>��C>®�>_y�:�,?r��>ᮞ�Y���K�'#��I02?�q^?�@�=!�̿�?����ž'Vɾב>��j�xG(��
���kl��T>�`������	��ɶ]�:������ѳ��$�� /?>cV=_��=^�=1��=_��<n�X�R#^=wlû_�=��н��u�Vg����=fR&���LR6�e��=١�=���P�o?��G?��*?��:?oKE>�>?��:u>&i⼼?�r�>��)=����z'1�خ���������D澃�m������=������=q�=>Ve >��H<K�>�A$=�2=����-��=���=a4u= 6�=�-_>�}3>Ֆ�?q������M��Δ���R?���>�n>�`[���?�>3��쵯�����W�?���?Ƚ�?�?;�j��>o�˾@�%=6�m>þt�5����>���0�>��<>�.�M���t�����?2�@0`?�0��pڿB�>�7>�a>zmR��l1��]\��b��3Z�8u!?�y;���̾��>���=�+߾�qƾ��/=r�6>`L`=�H�ne\�a=s�|��;= �k=�ŉ>�C>��=[?��A��=I�J=�1�=h�O>�����C7�y�-��1=���=L�b>C�%>���>7�?J�1?�	b?E��>�ʁ���ɾX��h:]>���=��>m�<� >�T�>�-:?�_I?�H?6�>=S̼>���>P�8�$^n��~˾�����s<{�?U��?8��>J�=��)�/)�fx9�=�۽V�?�C7?�I?�ܘ>Z�`[�H`H�C�>����=�dX>׹�=&����M����<=�"��m��&�">���>���>�V�>IB>I��=�ѯ=3��>��>�0��l땼&�=�>�3Y�M��=�M��s��= �Ӽo��2�o�M=��M=�t���|"�7�%�o��=�m�=�l�>�l,>w��>�o=2c����:>����zD�LC�<a���7sB�"$\�ҳ{���-�)P4���g>�9e>�Cʼw5��@F�>\p>.�c>B�?	sl?gd+>c�N�{�̾u���A��RqB�N
�=u�>e�/��:�1�_��qN�#Ͳ����>���>��>��l>u,�f#?�"�w=1⾫`5���>Hy��$���%��9q��?��[���Ji�LLҺ��D?+F��t��=�!~?�I??�?��>(��d�ؾ60>J��@�=|��$q��^��J�?e'?���>v��D���о���=�݋>=c׾,�1��9��xT4���h<Ss��W?�> ����Ǔ���(��|�mc��)�^�+���(�>�/�?!4�?AÛ���{��Ab����.��=%(�>s�S?�a�>�?%?��?�Ύ���ľ����Œ�=�=r?���?���?�HN���=���83�>1	?Լ�?���?��s?��?�y�>{9�;�� >�s��<��=^�>�J�=���=�d?��
?��
?�a����	�$��"�^��y�<ڡ=�q�>Ri�>��r>���=ѻg=�V�=\!\>�ɞ>�ۏ>R�d> �>0I�>�៾�<���8?r(�=�b�>@�3?�Y>p�*�;�[�:�μ��!�Z�s��UW��쬽 ���ҏ<�0M��������k�>_����?�jl>�	
��&?Nx��D�4@>P
�>����h�>�*_>@�@><ˤ>�p�>U�0>vl�>�>vA�j�>� ��|%�qg1�YP��:޾�I>�@��E�(��Z�/���u[��)��jh���n���p.���=#ώ?���%�W�'�(�.
B�W$�>j7�>��:?�΁�vأ�^�+>2�>���>�o���������۾+�?���?�d�>
7�>r�k?Ώ?r����Y�#J6��R��a��]J��mb�����{,m��羡x=,em?�`? �,?ڬ޽���>�8�?��G�G��4�m>�A��7����>)�>�=��1>��(�������ս�w^>��o?�?IF*?V�8�����>�?�)4?'�^?�,?�Y\?Q6�.� ?�A>A�C?��2?�~`?�2?6چ>r�!�,���v���>��[���PS5��X��¶���	�=��<>��<��<��-�2��uʽc3׽\o�<�h�s�d��=t>=�>��>��[?\�>T�>�u3?��#�z4�<����,?+��<;�{��h��*��������=��f?�-�?�Y?3�n>�C��4?�#X#>���>��4>��Z>�O�>`O��@���r=�0>�_ >���=b�5�W��@�	��ԗ��QK<e%>�?85*>�F>]<.>?����6�����>�D���*���ʾ�Z���B�NB0��G?unp?:7?��9=M��v�cn�%�=?!r<?�;?m�?[,>D��J���jG� 鉾�Ln>E�s=�|����|.��-�\��l����=.��8�վ#k>'���"��8��U��n�J�C��Y�A�=����fھ����<}�=�1�t�7O,�C◿�蟿ԢK?����:������9RC����=[	`>�c�>�c�<����G7��v��<���>�!>�=��徐l<�t�1��E�>�XE?�K_?Mj�?L,��� s��B�qt�����?Ƽ�?6��>�E?&�A>pJ�=ſ�������d��G���>���>��v�G��"��d���$�ʰ�>�;?�& >?�?�R?)�
?X�`?"�)?�)?�ؐ>�m��ȸ��A&?8��?��=��Խ�T�� 9�YF����>��)?��B����>b�?߽?��&?�Q?͵?M�>�� ��C@����>�Y�>��W��b����_>��J?���>T=Y?�ԃ?��=>Q�5��颾`թ�VV�=�>�2?�5#?8�?կ�>k��>������=-��>dc?�0�?��o?���=0�?�92>���>��=���>y��>�?#WO?��s?��J?O��>���<3<���:��@s�L�O�o�;��H<��y=����8t��R����<G!�;�]��#C������D�% ��:��;�}�> �m>@2��m�2>i;žV5���C>��ּ�R��"���>����=y�>6?��>���=7W�>�^�>c���'?�?�S?��;�Rb�_gܾLM���>g�A?�K�=��l�������v��V=vm?1*]?��Z�V����[?�q?�Sվ�y3�g���p��({$�%ND?k�?���<T��>3�?��n?���>�a��6�t�����	�e�y(f���G;M�>�F��Eh�ǅ�>��U?^es>�־�*������Z�d�fn���4?+D�?��?k�w?/>Y|c��ۿT��CN���_?U��>Q�����?iA�;�ɾ���Iؚ�G���<������"���͙��I-�͋��>D���B�=�?�Yi?�s?k_V?`�@Q�]�Z�n�p���P�j-�����LB�o�D��I�"Ph����f����6� |d=�N|���A����?Ε(?�W/��I�>k�����{ξ��;>���!�����=�9���ZG=մN=V}o��3��ͮ��?E@�>M�>^�;?z�]��;���1���5�|����92>쯠>��>�S�>u� ��l-�J��P�¾�U{�%�ѽv>�}c?�K?.�n?�� �+1�g~��!�!��#/�Ȳ��*C>�X>��>R�V��L�h6&��I>���r�>�����9�	�4�=��2?��>^~�>tF�?��?LW	�tC���x��R1�\|<�>R�h?�5�>�>)�Ͻ!�:��>��l?���>�T�>J���du!�M�{���ɽ=Y�>#,�>���>�Hp>��,�7\�V^��,u����8�g;�=9ch?����A`����>��Q?�_;^RO<�Ρ>�`z�ث!�F��*g(�@>�?���=_�;>��ž� �d�{��O���O)?jK?*蒾6�*��4~>s$"?���>�-�>A1�?�*�>+qþw�E�ı?��^?2BJ?FTA?�I�>_�=*���=Ƚ��&�"�,=��>�Z>Gm=[~�=>��;s\�/x���D=�t�=/�μvQ��}�<Ɖ����J<���<��3>y�ܿOt;���/�P��U���،�����M;�G־��ú�ž "��b>]��
��/��fd�� a�V斾��9����?q� @�>p��þ�&��*fZ�	�򾊳�>o���A}��-��� F�L~����< ��Z=�\��q�t�H�;�'?�����ǿﰡ��:ܾ%! ?�A ?�y?��9�"���8�� >B�<�.����뾪����οL�����^?���>��/��g��>Х�>��X>pHq>����螾�0�<��?=�-? ��>֎r�'�ɿX����¤<���?-�@}A?��(����IV=��>�	?-�?>�S1��I������T�>g<�?���?R{M=��W���	�(�e?��<��F���ݻ!�=�;�=�F=v��ՔJ>`U�>E���SA��?ܽ��4>"څ>)"�^����^�邾<��]>��ս];��y�?��\�(Lf��/�O���[>��T?�@�>VÞ=k+?�+H�LcϿ�[�кa?�H�?��?(~(?�鿾-ۛ>��ܾ|M?Q6?۾�>I�&�}�t����=�1��'����UV�c;�=���>Q>{�-�r��}�O�n����=#k�_Z̿�B0�!0��\�=A��=jWý�?���=�ۇ�ܡX�������=���=p+>4��>�5J>�|:>�'p?�?��>ih<b����2��o�z���e��g�V��D���$2�a��Aj���@ʾF��ϑ
�|=�X��iQ>�M;�=�	R����e��^�ϐF���+?C�>�jǾJ4N���<�ʾ?��I�¼�i��ξ�_2��Sl���?B?-���S�-$�/�������U?@���l���P�����='�ּj�=ć�>H��=���Ư3��hT�
x0?cw?*���ې���(>����-=��+?ң?}!n<�ѫ>�8%?�H+�_$�GjZ>]�3>9�>0�>��>d5��2gڽ�~?�T?�������>�ξ�	�z�Fc_=�>. 5�U��\>�]�<�)��Z�a�'���u�<X$W?�> �)�^��`Ȑ��A!���>=��x?��?m��>��k?��B?�E�<Á���S��
��.z=��W?��h?�W>�x����Ͼ\"���5?)ye?VtN>�i�6��{�.�$h�)?b�n?Rr?����7n}������T6?��v?�r^�cs�������V�K=�>\�>��>��9��k�>!�>?�#��G������wY4� Þ?��@���?��;<0 �ɜ�=�;?Z\�>��O��>ƾ�z������˔q=�"�>댧�Wev�����Q,�Q�8?ʠ�?u��> ���������=�ٕ��Z�?}�?p���!Cg<U���l��n���<�Ϋ=��
F"������7���ƾ��
�����࿼Υ�>CZ@�U�q*�>D8�\6�TϿ&���[оwSq���?P��>Y�Ƚ����?�j��Pu�\�G�-�H�����UG�>�>0�gi���y�{I2�q��LU�>$�j���>QBe�v���K|���;:�
�>=��>�x�>�������?��
�mͿi]��@��e�e?k��?2a�?Vl1?�#���j��#������[R?�?G;k?TNۼ깉�	���%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�d�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�G�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�=2�?��w�9剿�^�8Q���	?0���7�l>���=����1�M����y�X��Ϫ?��@8��?����&��3?��>#��6󐾊_��Ȑ>~R6>[H >�(�;w�#�E�Qn&�Gws=|�?}��?��	?�_��A���Cܭ=�?눪>��?k�@>���>�:>?�������<�`>�R>��?�;y?��?�<5>.��6�ڍ/���\�t�.���a����=v�?euj?m79>k����SN>�-�aU�F��B̧��O��j߽��n<��y>"��>Us>:�S���?Lp�8�ؿ j��p'��54?,��>�?����t�����;_?Nz�>�6� ,���%���B�`��?�G�??�?��׾�R̼�>:�>�I�>9�Խ����\�����7>1�B?_��D��t�o�{�>���?
�@�ծ?ji��?�þ� �������ݾ�u��,�<��=?j�:��>rݸ>�}G=�z�B��U:e����>�J�?C�?���>��?)�w��U{�w>r&�=�Ӆ?�!9?y��=`��l�b>��>�$6�R~�O��
+�?��@�@�N?+H���hֿ����^N��P�����=���=ӆ2>�ٽ0_�=��7=��8�!=�����=u�>��d>q><(O>}a;>��)>���P�!�r��\���R�C�������Z�C��Xv�Wz��3�������?���3ýy���Q�2&�?`��΄=�YY?Wi?WX}?\P?� h�f(z=o�n��=s��=k$I>�y�>�*?&�9?Z�?��<DY��F^��H��C�徺@����>�t>&�>b��>۸�>/+X�z.k>E��=��>>�C;����ӏ��電+�d>�ٰ>��>���>��;>��>�ϴ��2��lyh��v�Ζ̽��?0���0�J��1���I�������[�=nH.?�&>-���;п�����,H?y���2�&9+��T>��0?�UW?G�>N�nU��*>���ެj��w>� �)l�2�)��Q>�C?�qe>aEs>+3�-�7���O�Q1���D|>Li5?�4���2:�ܜu���H�w�ܾi�L>��>pCQ�����䖿E�~���i��}u=q:?ӡ?vV���簾��u������R>qrZ>�={Ӯ=Q�K>�m�Fƽ\�H�)B-=L�=��[>�?���>��=���>߼Ǿ�7���B�>��>��k>H
I?15?�E�$��3���߯g�)bZ>-��>�t�>�ݫ=�熾Յ�=Nu�>К�>п�=�웽��<�7Ƭ��N>S�6��8����J�;,���:>-���H8�)�3�קl;��?���yꈿ�ѾQʡ��t1?{�9?�(>>�x�[Ah�`m��8������?>�@��?.Yy�V#F�9��>jv�?xe�t'>^�?�&�>�B���V׾Dd?��	�e �S���]U��O�?�8�?�����m��F�Y���9=��?��\�Oh�>xx��Z�������u�`�#=O��>�8H?�V����O�h>��v
?�?�^�੤���ȿ4|v����>X�?���?g�m��A���@����>;��?�gY?voi>�g۾8`Z����>л@?�R?�>�9�z�'���?�޶?կ�?�F>��?��r?� �>�	a�n�0�2V���F���=�`�:0��>��>;i����F�p哿nN��qAj��G��Ic>B�*=NG�>[�޽B����R�=�����T��c5Z���>�q>`iK>q͜>�1 ?B��>���>c�=�̓�`	}�.���q�K?_��?=���1n�>��<���=D�^��#?�H4?{pZ���Ͼqݨ>^�\?���?�[?c]�>���9>���翿����W��<��K>V6�>bH�>	���OK>A�ԾB;D�(m�>�͗>u��.<ھ�$��|����C�>�e!?���>5��=�?��4?�ހ>ô�>�_=�Ƣ��rvK���>��?�q?��}?:3?��ʾle/��?����wI���=.�R?A$?�>��������wA=^�t=N��|u?`Q?Ҍ >�? ?��?<g?�(?U*�=�5��I��,����>��!?p8��A��-&����kl?�P?}��>fu���<ֽu׼����m���?\?p2&?���a2a�Yþ\��<T '���J��e <&FG���>N>7����T�=��>���=�m�A^6���a<K��=�e�>��=�%7���a�,?m�=�#O�u�>$6z���K�{ۜ>T�>I䑾\fg?S:G��f����Rq��
΂�oK�?���?^Қ?�н�*d�]�4?{�?ff?�L�>'����eھ�����{��(��'�)����=�1�>���<@ٽ�����;��R�v������(	�QM�>�n�>,,?�Q�>�>��>����"������.���f��u��#��o�)4��
׾As������ʾr`���>aԢ<Q�>U��>�w>s%e>�+�>T>2���>YW�>�~8>��R>�)f>��=z��=�e���~���R?~;¾u�'�$�Zf����@?��d?���>�}��?R�� �Rh?�I�?|ќ?�;z>�f�eK+��?n� ?t%
?�6H=a��oM�<�8��^v�������Y�>�bٽ�9���L��Ck�	?�.?똜��1;��ҽ�����f=�~w?c�?l<����b�É|�|�U���=������������C&�E�t�U����避���O, �ߢ�=^�%?�H�?��Ǿqe��aݾ)�n���8��@�>^j�>l�>-��>�?c>-��%�~�S�$;�?�/��4�>D�{?86�>�J?f�>?��Q?��K?�_�>7_�>�d�����>ep�<)��>���>h�8?*�,?�-?�b?�A*?�(Y>>	�"� �?�ھ��?��?_�?�3?{�?�L���k�����iE���#���{�S�x=��<Ofν$�]��1m=��a>�X?ڙ���8�����k>5�7?��>0��>���L-���<�> �
?�F�>( �~r�)c� V�>|��?��ρ=�)>@��=������ҺY�=������=�7��!z;�m<���=���=,=t�����?�:]��;�h�<@z	?�1?��>��>��	���	���G���>��>Շ>Os�>�����5��~����wQ�x�>!��?��?�+�:�=Z��=28��s��4�Ҿ�����B?�|1?(Oa?W�? |?.�?"�8>�d��B��ڞd�^���d?�1?��b>3���R���]���5��\?���>6 o��e"���+�0wʾӴ�<�lh>�V�P*f�kˬ�	�9��6�=9�GQ���i�?�	�?;vA�e_���㛿pT��>vK?gX�>�X�>8��>�4�j:j�5���7>Mr�>}�Q?��>s�O?>{?ǧ[?LmT>P�8��/��ԙ���2���!>o@?0��?!�?�y?r�>��>'�)�IྟV��L����߂��V=�Z>��>�)�>��>��=yȽ@c��`�>��c�=�b>���>R��>@�>
�w>	��<^�F?{0�>�ȯ�*��ۮ���D`��]˼ ?r?A��?�!? B=3��#,J�?A�(Ⱥ>ZR�?Y0�?�q7?��m�Q��=���;��ʾ������>� �>��>?��=(Ĩ=�u7>8 �>כ�>�I����3�8��e]�Ϳ?��C?*��=$�����8��X�n���#?�%�o��m�������&�{I�p�M���۾�T����b��%��Z���Q���.�>��9L��>[�%>�&�=Z�Ⱦ�ϽV�= �0>����`���++}>ъ���bf�m�˽m�E=r�G=NH:>8p>q�Ծ,vh?q�o?�o?c�)?-�>��>���U��>�2軗�,?���>}O0=?���n2��ľ�]c�愸�Fg���8���ľ�{[=8&��r|$>�
�>hL�>��R<V-=�a��OC�=��"��9x�䙄=`��=&��<z�=�� >�x>W~?vn�D)���/���~���D?0�>QA�>?ཥ ?���=����7��ZI���?�K�?���?�`?�r�C7�>Q��+ ۽�y/>�F0��ռ>+2>�zi�>��>�躼!1򾧷����üĝ�?�w@�8d?�r����ڿ1>1�3>9O>�$S�6�1��U��4_��e\�\ ?B2;��*̾+��>���=ʊ߾Fxƾ=0!=�l3>~�R=��u]��ۚ=qg��8F=�bo=�y�>��?>ֹ=f���*�=�X@=���=،Q>&���7PG���-�Z�5=c^�=;]c>'>���>W�?�c0?�Ld?�i�>��k�vTξ�����ŋ>g��=�ɰ>b��=�@>p�>�7?iE?}YL?B��>PW�=l�>�	�>�-���m�+�������< ��?�ц?�>�`{<B�?�ɦ�:>�7�ƽ��?b�1?w�?��>���L��	R4�Y7���ۼ2W=�(�=pQ���/��H��Pk�f����%>"�>�>�m>��Y>=>P@�=�S�>�[>`F�����
6=R��=~��P�$$��2>��B<BV�;�2�<��<��2<�=<�D[=�@=��;=y�>;?�y6>���>>.�;3оQd>Bo��s3���>:\����8�վe�jw���*��,�a�>d�>;���9�����>��G>B�p>~��?�w`?6Π= d}�M�׾]z���Ǿ�8���հ</B�=�-��ɲ8��mU�څD��9ؾC��>�׎>�>0m>�+��!?��}y=��ᾗS5�F��>�s��Ԑ�	�7q�/���⟿�	i��AӺ��D?�D���a�=N~?��I?,ߏ?�e�>�2���ؾ^Z0>Cd���=3��7Nq�*Γ�:�?~�&?d�>A��D����<<'2�>tm����8����P�$W<2K��ӒF>hM۾�����=��������yy>���\����>KT?�ʦ?.�w�h?��C!<�� 4��R�=��?
 p?r�@>��?[
?qht�p��ɑX���7>(ns?��?*�?�>rϻ=���*�>�D	?Ģ�?���?�:s?k�@����>�x�;��!>���2�=�>Y��="8�=�q?�>
?7p
?2����	�ļ�k��VM_�v��<�0�=gv�>��>��o>�|�=?�e=	~�=��[>��>@��>��d>c	�>��>���� ���#'?X�9>�f�>`C#?��>]=u���e߼����s�l(�,�ս����6���醷��Cϼ�s��e��>57��H>�?��J>Ly��G?
����ܼ�>j A>�h��6�>��>Y�>�՟>sQ�>��\>p�>Z�>f^ӾNM>}��"!���A���R�y�Ҿ��x>M;��v'����V�AJ�`0�����j����.=�ke�<� �?�����j�6�)�n1�F�?���>+ 6?�����C���>��>�3�>�����Z�������N྅��?w��?��>��k>�d?��-?�ƾQZ �1M-�لI��>� xX��,O�C�����y��`$�����`?�$x?�[?�}��f"�>ޜ�?ٻ2��4��d�v=�9����=C��>q�w�fů��̝����#j����=��?�[�?1�V?v��U�e���=��R?� ?l�D?��F?QlO?K��@T2?Ӛ>�:7?�r>?�70?v�!?���>LA��-^=[�r���Q>�G��x���Q��X��f
=�vg=	>uc>�2^�3�ٽ����n��|��<ɜ4=<g�<2lx<geo�� �=��=�Ѧ>ٴ]?�[�>�|�>�l7?���8������/??:=�t���*���F���4�}q>�j?`��?՝Z?imc>��B�4�C���>�<�>��&>�K[>��>)��D:E�}�=O%>��>���=TDM�����y�	�N���Z�<>�>�<?H���=���t@>������=5�>�۾��;�t���cS�ؐV��i>>�?
<F?4�-?�=z�bF����>�Ǉ���!?�[>?�\?R f?m��=��þf��EQ��P���ɂ�>��5���\�I���������<�^f��`=`�
�8G��[�b>Ԧ��S޾v\n���I�~_�͊P="��p�Q=aG�x�վ��~�ڞ�=l�
>���0� �t䖿㰪���I?5�j=���4NT�.0����>�Ә>ޮ>�A7���s��@�x����5�=l�>=X:>+d��V��ˇG��C��z�>�bC?~hb?4߅?.��@c���?������s���?Y�>�a�>*�>h�P<fR����G\g��*=����>�N�>u�!���F�߂������1"��E�>��?/��=�N?�L?��?��g?*�?��>.�`>�?��<���&?���?w�~=ܠнn6R��r8�4F��	�>��(?�rJ�(}�>�?�M?z@&?��P?�i?>� ��?�J)�> �>��X��W����h>RI?4��>�JY?i��?��7>�N6��������S��=��&>��0?�!?Y�?"��>'��>�]��B<">o>�>3�H?m�?옃?�iF�@�?(��>G�>���=AD�>�8?ԅ?��F?�\?EN3?��>�<$���G�������.�ռ= �<��=y>�z�����hm��&a��Ԟ��c=o�<�;z=�:��
8n�U~����>rr>핾�//>�ž�]����B>{{��`A���-��7M;�\.�=�R~>��?�q�><�!��9�=�B�>�w�>�>�9#(?|�?��?�Qe;
Jc��ھ�
I�$|�>�LB?(�=�Sl��P���u�ٲU=��l?��]?=7Z�rY��$`?��g?���	�������~�ݎ�D�b?�?����4#[>:s?��\?���>�t-��馠��eS��ul�m��=�{�>i�4�k>w��}�>��?�>��>��;o���ޖ�n��F�>��g?�e�?��W?���=�pH��	ɿx���|P����[?�j�>N��i�!?d�ع�˾y���W����2㾩د�T���Ǖ�@Q��H����~�I�ڽjx�=7? "t?�.r?"5c?�=���h�)>`��/}�i�N��G���@�C���D��uD���q�qx������1#@=r~�u A�&A�?U�'?��1�\��>������'�;�tC>]"�����zJ�=6^���?=i\=�1g��/�±��8�?o��>���>�k=?�Z���>�U�1��h7�����OX4>/��>�t�>Qu�>�6�:k`/�ݐ��@ɾ'a���ӽ'l�>��H?0�P?�_?y�����z"������<~g�8�@�4��=���>�����Ļ�.@���J� w���辭���^��kCw>� ?�*>�e?Ғ?x>�P���|0��a+��� �8��	L�='�^?� ?K��>P���N��+�>?�i?� �>悺>����O�M����<y��>E�p>O?�>X���<�����������Y��Y�=��r?�D�����ت>�O?�V���>
<=6r1��I���ԾT;�����%?I&>��>}xG�Ԑ���Cz��8)?S�?�H���!*�V#~>_"?4�>���>�&�?��>�/þ:��!�?[�^?SJ?BA?��>n�=�����Ƚ��&��m+=�i�>�'[>��k=Mn�=�j��|[�u���nF=�}�=|м㚸�п<Xⰼ̻Q<h��<�83>�5׿�_K�=�$	���Ҿ���;�q��F����j��$�BI��v#�� �A�,Խ���?L��IS�)mo���Z��e�?D>�?Aʾ:����D|�rix�c��E�>��!�z��j¾F<�����M��#��y�3�UZ���T�8^E��'?B���L�ǿ𹡿��۾R ?e" ?��y?%����"�D�8�U� >���<C���������m�ο�x��_?7�>���r4��;��>���>�UX>3�p>BH	����<��?*�-?M2�>P�r�ŏɿxw����<���?	�@�|A?��(���쾢V=���>1�	?A�?>fU1�DI������S�>7<�?���?&{M=�W�Y�	�ve?�}<j�F���ݻ��=v;�=XJ=+��^�J>�U�>Ղ�SA�1@ܽ5�4>�م>:~"�@����^�_��<�]>��ս�:���҄?�j\�cf��/�J��=	>*�T?�G�>/Ǡ=��,? 4H���Ͽ��\��#a?g*�?���?5�(?~���8��>��ܾ8�M?
R6?� �>�}&��t�]\�=��ꡥ�����(V�j��=9��>wc>�k,����O�屚�.8�=xa ��Ŀg�"����x=�;x&H�U�
�Ԡ��oB�E,���\�-���h��=m�
>�!R>C��>K6Y>&=>�_?k~?Q�>���=v޺a!����ƾ���=��O�ȍ�a�����:��(���X�p��1���A�����=�2�=�1R�g����� �R�b�k�F��.?��$>�˾N�M�U/<�Dʾ����ὄ��o��W?̾��1�Wn��̟?�B?r���W�x��̕�������W?�1����'��{z�=�K�� =k�>��=����	3�^S��0?1�?����X3���+>O��=|,?�(?Is.<�m�>�"%?&�)�=��q�[>��0>L9�>���>�*>DƮ�,1ڽ�_?RT?�m�q˜��d�>�A��=`z���d=.�>J5�����[>,N�<����ݱP�|���}�<�W?>�s)��P�)8��H{6�iJ0=6�x?~�?h0�>��k?�C?Gd�< ���D�T�6a��\e=�>W?�mi?�>����7yо1া��5?�se?t�L>[g����ȍ.�#���?�/o?��?4`���}�<1��\2�h:6?�vn?ID��ݬ��Q*�/N=�Z>dm�>�?�4#�KbA>��_?oX(�#��jԻ�W��5��?7@��@,�T��m��=6� ?tN�>鑰�C�޾O�+��Ũ�v�E���?5(��擿2����)��G?��??��[(��	>UD_��I�?�8?�ξJT�/I�0�G�5�߾�t�=k�=��+����!Y	��oP�V��4׾����Qѽ겟>�h@k�=�7? \P�S����Cܿ7Ay�3��A	w���?�4�>����U�־j+��`����F�#C�4t��O�>��>����������{��o;�I���!�>�g�>ؽS�]!��r���v�5<��>��>j��>0���彾�Ù?d\���?ο7���M��P�X?if�?p�?�m?t�8<w�v�-�{�;p�T,G?��s?�Z?�%��8]���7�$�j?�_��vU`��4�uHE��U>�"3?�B�>R�-�X�|=�>���>g>�#/�y�Ŀ�ٶ�C���Y��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���F�!�A0=�QҒ�ü
?U~0?#{�f.�\�_?*�a�M�p���-���ƽ�ۡ>�0��e\�bN�����Xe����@y����?M^�?i�?ѵ�� #�f6%?�>e����8Ǿ��<���>�(�>*N>XH_���u>����:�i	>���?�~�?Pj?���������U>
�}?�ζ>��?��>�X�> #�=���%J�NV�=O��=�;����>]�G?`�>�[�=�H>���0��ID�]jR�����~>��7�>o�]?
�O?��>V��`k?�.#��� ��;��o��3�(����ҽ�,I>H�:>#�>��L�x�վ�g?����߿�3����1>$�?�B>��?�3� 4����Sv?��6>)�5��������<�
����?��@)?Fо�����=N=�>:�=�w�D��M��=�;>t}a?ˇ��ˬ� �c�W��>��?��@b�?C=w�S%?H�ξj/��h���C� ��ʀ��ӓ=��Q?(ξꃉ�g�?-�V>���������k���>V �?O�?#��>nFa?�v��.�2�=�!g>�Z(?;y�>6��=��о���>�.?��-�N���^�Ǿh�?$@^@�]l?Y�ʿ��ܿ��|����Z���3=`0z=7�>�7�P �=b��=K�潹-ҽS/>��>l�>�8�>ľ6>C*>���=�����&�\꠿����3�˸	�i���Lp�0T�91S��`�qh��I���ꍼ��������;z0���)�w�>8�H?2�V?�g?b��>ܓ:a��=�+ݾ~�%>�����=��>ME ?�'>?\0?�>$�����q��ur�O�¾ۼ˾Ք�>�(a>��>3��>��>�S½���<bg�>d��>�l9>��Q=��=�]���0>Dg�>�?�8�>�H<>��>Xδ�v0����h�jw�� ̽h�?�����J�
2��G6��H����i�=b.?�n>���=п����!1H?�����)���+��>=�0?�bW?�>S��#�T�50>��9�j��\>$% ��}l��)��!Q>Vj?��k>o>�s.�0k3�j.M�ޣ����>�%4?�ʾ�>:�&#w�*vH���۾r�D>C`�>�<$�zF��:��u�}���V�~k�=�9?> ?�Χ�j�ľ5�x�[U��<=�>��{>��q<��=n�.>����$�	��/>�"�=EK=�k;>�?�>#��=)J�> 񡾄�<��t�>�:>#��=�1<?�o ?��m�,��'䄾�� ���~>�g�>Aʀ>Bn�=/?��=�=^b�>�Qw>k!�>��`���+,���r>�D�c�`�����8f=�{��6�=x/q=�����H�g�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>��G9���䍿�WL�M�=���>ML?�׾�@>�8�^�n?� ?#��瀧��ƿaw����>��?�M�?�L��g����M���?�U�?�D?��v>���"��q��>uOO?YY,?�s�>� ��\?�ȸ?闋?��T>�_�?�f|?b�?�F�G�Q���)>����<r`@<��>�$>�6����L�p%���+�� Y��*����=Li_=��>�����7>���䑑��n���>S�">u�c>P��>~Y�>���>�&> ԇ;�G��&v�=�m���K?�4�?�0�.6)�pU�=�H0�sD����?�n1?񐁾�U����>�i@?p�L?�?R??��=g�/�̈���f���1ľ�ߦ����>�?�T>P)�<���=z>�=sR�>'�>,Aн�ľ�:S���=��?��	?���=��Q=�!?�9?E�>���>�[W�`ᠿ�F\��[�>��>���>(;q?�-?�_����3��f���ۨ�v�R��=Z9]?Yp?��>
ܚ�+���z��=#y��{Q��r��?ID9?}嫾��>�R�?�Q?!�W?��>��D><���>(�>�?�
�iL>�2+%��-�� ?�@?��>�3���꽊����0���o?�Y?�L#?�� ��{Z�)Vþ�c=�v���?J;;�<s[��`7	>6�+>�D\��]�=�%'>�=�$p�ĉ7���<���=)��>	��=��F�XŶ��a?8��=�־[�c���E�3 O�*v>�9�>es�%�C?��d�ի�����ӏ�������?���?�j�?��¾;l��C?R�?�)?��=`N�<����o6)�-4վ:u�]�߾6"f>���>~~��մԾ#���Vٸ��~��q�=F��a:�>��>��?�z�>�Z>fG�>y����:�}��;� ��}]�2�I�=�>�#�i��V��O}�RP��þ����q��>�"X�֬>��	?Գa>��k>M �>!a`��!�>�uk>��>y��>{9a>�_&>f>��-<�Q��3MR?__��4�'�h���h���B?6=d?�o�>,�h�͍����{?w�?�`�?m\v>;�h��C+��??9��>����g
?��:=�P��\�< 9��>���9�������>^Eؽ�:���L�yhf�3g
?�4?Ht��:�̾s}׽W��d��=Ǆ?�v,?T=0��%c�96t��rM���?��5���B������'���v�0G���g��Фv��{)���=o�*?��?��j�9W����y���D�YLd>g��>�h>F��>G��>p����-�9�f��I:�Z㘾�3�>,�}?z{�>w:E?y??�8R?ghG?���>�;�>���߸�>/S�<m��>���>�<?0�3?Q�1?|�?�i%?��T>�>׽����&)޾u�?��?c�?[ ?;?oV���
ƽC6+�Hh���|�Ζ�Tw`=^�<"i�O�T�㕅=�bR>l2#?�i�<��4�Q6�Uo�>a<?���>�P?%�`���;p�M���>�?O��>6Wþ�r����#�V�>H�L?���51=A�>�E=/�2<��ּAJ�=����}�<f5==o�H�?ݺ5��=�3�=W2�Xݐ=��<��/��4�k�>��?^��>�N�>�}��i� ����\<�=F�X>IS>�.>'LپMz��p'���h��y>8h�?�X�?��f=��=|m�=q��A������6�����<��?�A#?U T?���?��=?�e#?B�>�:��Y���\�����?N!,?P��>D����ʾq�h�3�y�?�[?6<a�^��F<)��¾c�Խ�>E[/��.~�[��;D��@��X���{�� ��?���?}A���6��y�~���Y��?�C?�!�>fX�>V�>]�)�T�g��$��0;>���>�R?Zd�>�$@?��?z^?�7#>�#��P������/�<g=^>nBT?��?���?�9�?��>m9>1�B�U{ݾ�����:���0���^���5>��Y>�@�>3�>�f>���=��>��Z̽j��3�&>�>�>���>�/i>d�>���>Qs>��G?g��>P[���������5����+<�k�u?���?؊+?�=p����E�y<���F�>Hj�?G��?.*?��S���=�ּ'ɶ�7kq�1 �>���>"(�>��=i/H=?�>3��>���>�=��\��{8���M���? F?qZ�=8�Ŀs�p�pRp�������;����b�����mf�G�=�8�����S����\��I������F精�����z����>Ci=�,�=���=�Į<i�ټB/�<��S=kН<��=��p�%�B<�s8����Ƃ������K<�4<=�E���V�w?/XO?��3?5�0?�Sx>�=�V�Hi�>|�r��??Y>!~��6Ⱦ5
7�� ��DW��È���(|V��ꊾ}>�U��]�;>�>ߩ�=���;��=֣D={��=���<\��<���=��d=�N�=��=���=�L>�Hm?v�V��ƫ�J�s���=��>�Ό>�>o?߾4f?Ks>zA��"�ȿ�t���p?}��?#��?��*?B�{�~>�HW��T�=H�>�5��i>>�Y]>��W��>:��>�}F�NG��|�0�l��?t�?��O?^�y�c�ֿi�3>Ў�=<E�=��2�/�4�K׊�"bz��e�j��>O��1E��x�K>�	��&�T3�ed_>a�>�n>�0a<�=0��x=t+R�O��=��>�W�;��#>��>�>=��k>*ج<U�=`�>Z9>��*>�f��zl���=|��=_%>���>6�?ta0?_Wd?Q0�>:�m��Ͼ�E���A�>�0�=�E�>nޅ=2rB>���>g�7?�D?P�K?y��>9��=i�>�
�>��,���m��m��̧�]��<s��?<͆?YԸ>LQ<��A�����f>��MŽ�r?�N1?�f?��>�p����������/�$~	����=���>d��!�<���=��9�V|ӽK�L>V?YU?��>!�>_�m>�.�>j��>��6>��潣��;�jջPݍ<�T=�Nj=#��;��j��d=�ͼ=l}<K�w��hf��x�x�K=؊/>���<H�=Qs�>XQ�=�<�>D'�=��>�>�B���l�f�=SԚ���O��No�?1��J���ܽĒ\>&Ph>"���F���-�>�o>��h>�s�?���? � >俈���>����EA�[o�d�&>��>f� �K<�X,_�&qB�����ɷ�>�*�>֡�>o>�$-�7>�"d=���0;4���>�.�S{��'q�����ş��h�m��_�C?�ׇ���=��}?�I?Cm�?l�>\����ھ;�+>�䁾}�=y�EVt����$o?g�&?�=�>B��,D�E̾�徽UƷ>�kI�Q�O�4���۰0�������m�>7�����о3��h������.�B�h_r�g��>�O?>�?�b�8Y���ZO�����A���j?Lzg?��>0??[B?y͡����%���D�=t�n?��?�=�?�->--�=B��E��>�2?���?�$�?-�t?G3���B�>�X�=��%>��c��^&>�#>6��=�<�=�z?��?�?��� A��!�fM龋"M�~w=��
>��>� >�w<>���=���;.΀=�)�>���>���>V#q>�e�>=�>�Y���	��B!?]��=�$�>��1?��|>��B=����ֽ<_�\� 8K���9���Q���ȇ-=<�x<�^w=a������>��Ŀ.F�?�%Z>r���?�y�Jڼ�Cm>|/D>�[ͽ�I�>�Z]>���>���>�B�>c>Y�>��->���>�&�Hu8�����>9�.ƾ�Ҥ>��7�$Ұ���� �˽D���Ǿ�5�ӿh��iz��̿>:�?�Ck>�̓�"i��< >!��>��.>�D?�tg��������=��?��>1.��袿\Y���[�K�?5��?��b>���>h}W?pN?�X2�rr2�"Z��\u��qA�o�d��`�[䍿1�����
�ZM��Ȱ_?.�x?rOA?�׋<�Cz>���?��%��ю���>b/��;�vJ?=� �>ń��+a��Ӿ+�þ�e��yD>"o?B��?8�?DoV�1z >���BAI?�@?�>�>�gk?�q?����?�0?�v?g��>�M?~�9?��>�/�>�q=������~>$��{�z����}
�Q8�=� =��K���=X4>��n�U��Cš<1c�8�!���(=��=S\�=F=���>��[?n��>l�>BK6? ���6�T����%?��5=����]l���Ƨ��Y���}	>~k?�@�?��Y?^\>ڜD��H�~�>��>�">�1^>�l�>��0�B���=t>*5 >�ʹ=e�,��h|��	�����f��<�1&>���>��`>vP���`>�w����h��h�>_�/�$J̾��6�3�E���9�\���U��>Et@?_?�O�=�4㾫�齗�W�fl/?DA?n/]?ڵx?��N� ��	�-��&��཰ݔ>���<�
	�1A������=��g���)5>�d�����gb>"��ϙ޾�kn���I�:�羃UP={A�i�R=�]��	־h\�ߘ�=�	>w����� ����Ҫ��-J?7Cn=�5��6�U�N���)�>���>��>M�<�[x��u@�ٗ��f&�=���>�q:>�򜼜�(uG�+��p>KC?�_g?C�?죡�ZJ��mI�݉B��/����J=�?�R�>���>�vN>�N��VžW>�&r��?�K�> =�>t:E� ]��ֽ�@���T�����>��?��6�?BoY?���>�&l?��'?~?�>��h>z׉�

��kA&?؏�?lx�=!�Խ-�T��9�'F�M�>*�)?hRC��×>q�?o�?��&?VeQ?�}?O$>² ��<@����>�i�>��W�f����`>��J?�y�>�~Y?��?O:=>h{5�1ɢ�w�����=mH>T�2?d#?$�?�׸>��	?Yۓ�;;o>=��>B� ?���?��l?��]=��>+]�>rɆ>��`=���>�!??W==?��<?��?O��>	߼'�=���?��1�<�܏�b<򼾼�<L��<��ὦlҽ/�����;;�D�IWl�u0�<���=�K�Q`����>+t>���gn2>�aľh܇��A>P���U��ˈ���7��\�=N��>o?[Q�>� �_�=���>�(�>���:J'?�)?�J?I����a�,4޾��P�8�>B?�B�=il�+����v�-�b=<)m?Y�\?��[��:���R?�Pt?� ��������mھ�O��k<?��>ۅ��@�>�?��S?�W�>{SܾJ���Z����NW���5�-N`=���><���.&�|Ў>�8?���>���=��8=W�̾=;k����sp�>�Ē?{߻?�R�?���=�r����N^�M���ö_?>E�>�⨾�W#?u���a�Ǿ�Ԋ��\��܌ܾ<X��д���u���؞�����i~�5g���i�=*j?�q?\lp?=�]?����-�c��5\��A|��V��!�z}��gF��wD���B�b0m��4��t��q�����B=-J���;���?h�!?�I�w��>����ܾ�O����[>ˇ��O$�{R�=�xü'ѳ=$��=��$��z���h���P?�t�>���>Lr8?6�V��sD��<�$�0��`�A�I>웰>�Л>�c�>�	���_�E3�N�Ͼzt��䪽grh>/�x?��A?ɕX?�Ͼ$T���n����׭�iE����n>�����2p>»#����%:�nGR�����w5�����z��E0�>��?iv�>�8�>��?JO�>^�����臐�R�B��(ϼ5YJ>v�\?o$?��>_��V$���>��l?���>��>xl��7d!�+�{�q�ʽ���>��>o�>b#p>VS,� \��h��׍���+9�3�=u�h?�u���a��Ʌ>c�Q?��:m�L<�h�>7!y�j�!��򾎭'�>#>x?��=��:>q?ž �/q{��剾s�<?,��>H5�b��(�>lO6?�>�C�>�t?ԋ�>��}�f�>��?lrk?c�O?IK?�&�>��>�[7�	ĽV�'��p�=<Қ>G�>>����o�:>�E�y s�>k��]�=�w�=	�s=���uȽ;��i�_+�=��=õ�=�Yۿ0K��Zھ�q�Ӛ��	����ߘ���ᄾD���#���V���Sx��@�@%)���U��"c������n��)�?��?$����ϊ��/�����������¼>zp�ˬ��d���������K�ྭ\��o�!�h�O�Җh��#e��E+?��c��A�������_����>%��>��?�^���D�QK/����>��=�μ���������uʿ3Z��;�p?w��>8D�E����>�1�>��>���>e���ξ;!�=bf�>'M0?�w?۴������ڳ���=���?�;@��A?d�(����i�Y=�F�>�	?��>>�0��T�x���J�>�#�?�׊?��Q=oWW�����/e?8�	<�F��7�Q��=d��=!�=�g���J>He�>���A�YܽN4>�<�>� ����^��ͻ<D�\>ڷս�A��zք?�z\��e���/�"S���i>��T?�5�>��=ȱ,?�.H�yϿħ\�<+a?,�?<��?��(?ȿ�D͚>a�ܾw�M?D6?���>-\&�s�t��g�=�!���h��}(V���=�>�r>��,����эO�	�����=����ſJ�6���%�1M>�J�8�b��q=pP>A�,����n�C�y�rۮ=�P>�*(>�"I>��R>(=�=��Y?��p?��>���=[�=#۾�?���>�51��9ᾑ	���ƽ˃���/�/M�H����������ξ�Pe�"͚�7f�_}������^<���(�%cc?��?I)<��U��	����̾����k���ڽ�f���U$���o����?��|?�;:��yW�X�����M뢽��?�/�����NY¾1k�=)B��tS ��H�h��h��q$��'&��t0?��?
���"Ȑ��()>4����=a+?D%?��h<ϻ�>�%?�R)�;� �[>�-4>��>ڂ�>�!	>�Ů�F�ٽ_?LT?߸ �c��ӏ>�f����y�:.`=��>�4�<6�`.[>3+�<ء���wW�y����G�<� W? d�>�@+����T눾nE9��p=��z?�Y?��>�h?<�D?:�<E��f]S����4=ȪT?�j?ҧ>;��h�Ѿ�/���6?gb?PU>؊a���^+�)���?�To?^�?�#�Z�}�����~��FY9?�cj?kQK�H̪���$�G��w��=Η>�!?��>�햏>rQ?���ݬ������/��?"
@X�@]!:���&�_��=f�?q�?�پ��f����������>7R?�\���.��
�����c�Z?�P�?�'?A¹���
�y��=p!c�^��?S�y?F ���V�f�9��T��]��y�A=]eX>R��E>��.��oO�V׾�*�m�U��RܽL٢>׊@&	+��B?ٽ������ڿ1�^��������IG?j?����վ&������+ׁ��a���Ҽ���>eA>A���f����z��9���Ⱦ�>oKݼ\N�>�P�Ca�������+<���>|]�>�ʄ>�?��5���
�?�����˿��������Y?儞?��?��?)<�Z����{��!ռ�]F?.Tr?Y?݅K�~UU�^�0�ôj?����q`���4���D�P�S>B
3?n��>>�-�7z=��>xS�>�'>h�.�-�Ŀ�춿�_��]Ϧ?���?�E꾥��>�_�?�+?�[�0 �������*�����"A?I�2>~�����!�D�<� ����
?�80?����`�_�_?)�a�=�p���-���ƽ�ۡ>�0��e\��N�����Xe����@y����?I^�?g�?е�� #�d6%?�>^����8Ǿf�<���>�(�>�)N>wH_���u>����:�%i	>���?�~�?Lj?���������U>�}?7��>�:�?�\x=F�>���=.����;.<Y2>���=�񽢤�>��6?���>`�>_L��42��+[�TVT��e �h�B��_H>�F�?4�a?�[%>~��<+5t�M�?�����Y�ֽ����_��|2��Z��h��>���>��@>�1��0���O?`0߾l�ۿ ��:��=G�>�1�=��
?u�ؾ���[�Y���c?J>�6�U7��&l����k�7�?���?�F?� ӾX��kb=��?�/B;X�V}�����k>�`y?V�h��"��^id��YD>�
�?ª@���?��A�I��>�g��AH��W�����=�F ����V?����-���[�>�pm>Q࠿"���~�����>k�?x\�?�`�>'�i??]��M5�:>��g>f�1?��>zpx>���?�?�uT?���C���	���}?�9@h@N��?�+Ŀ$�߿�}���Q�{\̾M �=Mw�=��v>�R!���=>v��=h,=��=�Fz>$(�>o�>�a>�v>b3>Ф�=�r����/�]U���؝�{@E��4�xڸ���W��鱾��:�s=	�h�ؾ.�p�F*�<RM'����:�3�w��+<��[��=pC?;�f?H`t?���>����=��B��g���M�<רo=�� >��6?7?��>ڢ���������Y�����bʾ)�>d�>1��>U��>��y>#9�*�>���>���>�L`>��>�������6>�Ң>9��>xt�>v<>��>r˴�,.��*�h��w��c̽��?[���J�^4��q2������^-�=�N.?�=>���6п���1H?z͔�S(���+��>��0?SW?r�>u.��>yU��>���H�j�^E>vE �ַl���)�!Q>n?d�f>s;v>E13���7��P�V^���~|>��5?���̧9���u� �H�l�ܾ�PM>�־>�G����r���<�~��\j��Jw=�A;?��? r��d$��'�u��`��I�P>(�]>J=z�=׌M>�c�90ƽ�F��2=�=	h]>��'?L��5p�>�E�>�$����L=1�>��p>P�="�=?!�?㧮;��<NO���\=q��>�z�>�B�>�%�=GnC�u">�[�>��P>k13=nY!��3U���2�k��գd��ؒ���阅�J�.��[<絼:�3��Y�����;�~?���(䈿��e���lD?S+?_ �=;�F<��"�E ���H��G�?r�@m�?��	�ߢV�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž5Ǣ�ɔ	�+)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ %�>���eY����V�s�3z=b�>��H?�"��!�d���?�h�?�<?x��@���Ɋɿ/�v�`��>0�?�a�?�vm�yϚ��4@�w��>:��?}�Y?��f>�۾�U��Z�>�@?�tR?�ܵ>Q���Z'���?i�?҅?��8>��?�en?�>�>��'��E;�㬲����%`�=�r�<�ߴ>3�>����NC�B���y����n�1� �2VP>_0�={I�>�u�V%���z�=���:�&��ѓ��>*&>�;3>���>��?m[�>
��>;5<����JI������7�K?s��?���4'n�S�<9��=^�^��!?�>4?��\���ϾŨ>q�\?࿀?� [?�Y�>X���>��2忿������<}*L>�I�>>=�>�戽5K>\վvDD�H~�>���>5����4ھ�)���H���Q�>�f!?�w�>Y��=ҹ?�A?��P>�+�>�Sj�E���\m���>��?�p�>B��?��?���x����*X��ife��/=��N?��%?H�>
���4��ppD=��>��)Ͻ�k�?��7?ղ�i��>��?�;<?�A?px>��������h��>x�!?�����@�l�%�7��*�?��?���>1���ӽ��ἒT�@���?c�[?^&?���l`��%þ��<�W�u� �1�<�����>9>,����8�=�>l­=�l���4�}�<u�=}�>e;�=��9�}򓽪t?k�=\R��dr���+rD�+M{=��>�ֳ�~�?�ؽ�5��4o��VP����ϽL�?ό�?uޖ?I���}Jo�X� ?d�?��K?ݷB>�_�V�LT/�����;�I,��$R>��>Y���e�������+�����(>�j5�Sl�>ˤ�>�w?���>f>�X�>�����=���̾����Q]��%�M�Z�� "�����3i�n�������̾GC��5�>�N��%�>j�?�<�>�MT>#�>vV�<j4�>�-�>��>��b>��w> g;>T]+>��=�Eƽ>CR?g!���(����2į��\A?�&d?���>��m�re��{k�N ?fd�?:�?h�s>��h�'�+��*?�y�>���>
?;C@=��»�؃<�S��>��Ỷ�ת
���>"Sս�b:�J3M��d�w�
?9�?�%���̾��޽֢��"�=_�?��)?E�*��lR���p��
X��?Q�Ϻ��^�L��ѷ$���p�k���0����ヿ|t(�s�$=��*?˥�?���A�l����j��M@���d>���>ܐ>E��>��Q>(�l0�<6_�f�)������>�p{?oQ�>�t7?�
>?�S?�XB?��>�/�>ɱ��ts�>6)d=�+�>t`�>�5=?��!?��$?�?Q?�[9>��#�D�ﾂ�׾$�?��#?KG*?O�>���>��f�?����D��#�۷k�^��z����M�<4.����=n�K>h�!?r0�=�4O�6�Ƨ>y)�>4��>�?+;Ra��Sڕ�2�1?�F?s-]>//-�<˙�V�0��><�?�hL�M���m��=k�=���"�'��>-�ƽ��=6�>d�E=9m�<��=l>Gt;&5>z?p��T=�)��~��>��?�N�>r��>矇�V� �v=� O�=S�X>'`S>�N>�TܾIn��梗��ff�{j|>�z�?�5�?[/Q=]�=���=�����������¾��<Iu?�$?BrT?F�?H+=?��"?�K>���C���w������2�?��+?ά�>���'�ƾ ���d�2��?z�?)�`�ձ��*�*�ľ��ν�>$)-���|�|߯��oE��X$�;���V�����?tn�?A�E���3����\���2c����D?���>4��>M��><�(��.f��y�@�@>Wu�>�O?�8�>�n??5w?��Y?��%>���iP���Q���1���C>@?߬~?g��?��|?��>Z�>�e���HU۾o�3����� ����<��D>�a�>G��>�>�;>����:��C����>&>���>��>�>�n�>�ߧ=��G?���>���e�J菉�X��y;��su?��?ʛ+?��=�Q�'�E�D���	v�>�b�?��?m)*?�mS�C$�=4�ռ奶��mq����>&9�>(:�>���=�D=��>��>V��>���i��h8�v}M���?Z�E?]t�=5�ſ�Bq�p�t�������<U����wd�����nR���=�$�����rX��-Z`��栾�����7��FꜾ�-���>�ĕ=�?�=�[�=CI�<�[ļw�<�:H=<�B<m|�<��w�J�c<�Y@�p������@-a��3F<n�:=���j궾S,q?��Q?i3?o+?0>&>ΑL�Ve>���=��?7>DQ�/L��	V�����XX��\) ��S����_�Ø���b�=M�=ѡ~>�_�>�b_=����$�=}d�<��s=l)=�.p;æ�<��:=���=Z��=^�=A#>OPk?wHh�Y���Y�c�T�!�U�?��>���>;|���(?�o�>�ޏ�VNȿ"��Utt?�c�?w�?�8?�2ѾHY�>֜e�jc=B�'>x3ƾ>[>�b��V��>��<>Ȇ����s�=��?� @j3:?����NٿpR4>}/�1�,>��;�L�.�Sw~�a@��ԡ�P��>�7e�&�ھ&M�>����D.*�H�O��{v>�F�>�á>�]�<=��c=Jͽ��>Y���8��>�@�>4x�<݁ݽ���=��x�>o,>�o�=��S>���=֕>p��=%t> ��=E��>8?yN*?��\?#)�>5�:��w���Y¾�8�>�23>���>_��=���>ܾ�>�5?��B?M�J?@Y�>��=���>�|�>vW���\�p(��$��^�轋�}?��c?���>~җ=�J ��W+��oK��� ��h?�p?l�>���>0t�i�����=��+������Ӗ=� �>�v	���`>��=8�轂sľ���=b�}>>��>�L�>�9�>6p>�o�>��>�l�>NL >��=���=��=�[���.>�<��<��m��fO�񸲽��<��¼}�%���E�=�����O�=��>n��=��>���< 9þ�>s���V\�� �=%���"M�U�p��z���(����+�U>*R>ӿ*�t��t�>��>�`�>�*�?V�j?LP>��:��=����f������j>~��=�<�<��n^�x�P��է�%l�>(��>T�>��l>�{&�D=�A$�=��ؾ�U3��8�>V���dZ������e�Ӟ��Ԝ���m��T'�j�8?������=D��?:�P?�?P��>�Y��t��;a>��]�'�ƻ-�zj�B5����?�'.?�0�>�2����G��F̾�뽽�I�>ۃJ���O��ȕ���0�c%����ζ�>!�����оi!3��p����/�B�Q�r���>
�O?��?�b�"Y���WO�9{�{i��Q?�_g?9��>H=?�|?�����������=�n?���?�N�?��>��>��򽑟�>>�?7*�?���?�Ќ?,��GP}>�=�=�>��,��>W>%�a> �x>�I�=�(�>�>t?��_��`����)�$����=�(=�ih>s��>�<�>��s>���=�,�� �=��>?� ?%�>�y>���>y=j=�K��<� �qA'?]�=�C�=��3?Q�2>4">$r�a@D>];�O!+��Tk��`)�K��=�_>�8�< �>�;�=��?,~���`�?��C>�� �q#?z.оaTN>�r(>��>���)�>���;��>M�>���>^�=��>�:@=�޿�V�>o�,��O��o��&�O�}����>�T��`��G���(��=E��о9�!��\�����'b*�Ψ"�e�?	z�=������J�X$�>ơ.>"��=��2?�;*g��>�7?�P(>_���#��Ls��������?���?�J>u��>��Q?��	?�6���0�8FQ��zq�d�D���^��W��򎿠X���
�%�a�_?b?��}?�kB?�h���Y}>�Wj?l����p��Ve>z4:��b9���.=B��>w��$�l�vؾ�ƶ��н7�>��a?��|?��?؞t�\�>�*�F"0?�"?0?�0`? 4J?�u����>O��>:w�>�~�>x�+?��+?S�?�*�>�#->��`��=�^����c������=��J�;f�>l$.���M>g��=�f<�W=���= D<<��x<��I�7�=��=�|�=I��>�{\?���>�F�>D�6?����8�����h�,?�b6=�߁��f������.�@7>��j?栫? �Y?��b>��A���B��\>e��>��%>Nr[>�Ұ>W8�@�C�U͆=��>��>ta�=�[C�~��bA	������c�<��>�A�>:��>��,�@�;>1ҟ��9r�ѡa>S��D��M�R��H���2��b����>:�I?��?�K8=C������7�e� �?�XK?�T?�wv?�Z�=�~޾�A�H\M���/ӕ>�1�8��I��'�����0��ȼ<K�Z>Q���8G��[�b>Ԧ��S޾v\n���I�~_�͊P="��p�Q=aG�x�վ��~�ڞ�=l�
>���0� �t䖿㰪���I?5�j=���4NT�.0����>�Ә>ޮ>�A7���s��@�x����5�=l�>=X:>+d��V��ˇG��C��z�>�bC?~hb?4߅?.��@c���?������s���?Y�>�a�>*�>h�P<fR����G\g��*=����>�N�>u�!���F�߂������1"��E�>��?/��=�N?�L?��?��g?*�?��>.�`>�?��<���&?���?w�~=ܠнn6R��r8�4F��	�>��(?�rJ�(}�>�?�M?z@&?��P?�i?>� ��?�J)�> �>��X��W����h>RI?4��>�JY?i��?��7>�N6��������S��=��&>��0?�!?Y�?"��>'��>�]��B<">o>�>3�H?m�?옃?�iF�@�?(��>G�>���=AD�>�8?ԅ?��F?�\?EN3?��>�<$���G�������.�ռ= �<��=y>�z�����hm��&a��Ԟ��c=o�<�;z=�:��
8n�U~����>rr>핾�//>�ž�]����B>{{��`A���-��7M;�\.�=�R~>��?�q�><�!��9�=�B�>�w�>�>�9#(?|�?��?�Qe;
Jc��ھ�
I�$|�>�LB?(�=�Sl��P���u�ٲU=��l?��]?=7Z�rY��$`?��g?���	�������~�ݎ�D�b?�?����4#[>:s?��\?���>�t-��馠��eS��ul�m��=�{�>i�4�k>w��}�>��?�>��>��;o���ޖ�n��F�>��g?�e�?��W?���=�pH��	ɿx���|P����[?�j�>N��i�!?d�ع�˾y���W����2㾩د�T���Ǖ�@Q��H����~�I�ڽjx�=7? "t?�.r?"5c?�=���h�)>`��/}�i�N��G���@�C���D��uD���q�qx������1#@=r~�u A�&A�?U�'?��1�\��>������'�;�tC>]"�����zJ�=6^���?=i\=�1g��/�±��8�?o��>���>�k=?�Z���>�U�1��h7�����OX4>/��>�t�>Qu�>�6�:k`/�ݐ��@ɾ'a���ӽ'l�>��H?0�P?�_?y�����z"������<~g�8�@�4��=���>�����Ļ�.@���J� w���辭���^��kCw>� ?�*>�e?Ғ?x>�P���|0��a+��� �8��	L�='�^?� ?K��>P���N��+�>?�i?� �>悺>����O�M����<y��>E�p>O?�>X���<�����������Y��Y�=��r?�D�����ت>�O?�V���>
<=6r1��I���ԾT;�����%?I&>��>}xG�Ԑ���Cz��8)?S�?�H���!*�V#~>_"?4�>���>�&�?��>�/þ:��!�?[�^?SJ?BA?��>n�=�����Ƚ��&��m+=�i�>�'[>��k=Mn�=�j��|[�u���nF=�}�=|м㚸�п<Xⰼ̻Q<h��<�83>�5׿�_K�=�$	���Ҿ���;�q��F����j��$�BI��v#�� �A�,Խ���?L��IS�)mo���Z��e�?D>�?Aʾ:����D|�rix�c��E�>��!�z��j¾F<�����M��#��y�3�UZ���T�8^E��'?B���L�ǿ𹡿��۾R ?e" ?��y?%����"�D�8�U� >���<C���������m�ο�x��_?7�>���r4��;��>���>�UX>3�p>BH	����<��?*�-?M2�>P�r�ŏɿxw����<���?	�@�|A?��(���쾢V=���>1�	?A�?>fU1�DI������S�>7<�?���?&{M=�W�Y�	�ve?�}<j�F���ݻ��=v;�=XJ=+��^�J>�U�>Ղ�SA�1@ܽ5�4>�م>:~"�@����^�_��<�]>��ս�:���҄?�j\�cf��/�J��=	>*�T?�G�>/Ǡ=��,? 4H���Ͽ��\��#a?g*�?���?5�(?~���8��>��ܾ8�M?
R6?� �>�}&��t�]\�=��ꡥ�����(V�j��=9��>wc>�k,����O�屚�.8�=xa ��Ŀg�"����x=�;x&H�U�
�Ԡ��oB�E,���\�-���h��=m�
>�!R>C��>K6Y>&=>�_?k~?Q�>���=v޺a!����ƾ���=��O�ȍ�a�����:��(���X�p��1���A�����=�2�=�1R�g����� �R�b�k�F��.?��$>�˾N�M�U/<�Dʾ����ὄ��o��W?̾��1�Wn��̟?�B?r���W�x��̕�������W?�1����'��{z�=�K�� =k�>��=����	3�^S��0?1�?����X3���+>O��=|,?�(?Is.<�m�>�"%?&�)�=��q�[>��0>L9�>���>�*>DƮ�,1ڽ�_?RT?�m�q˜��d�>�A��=`z���d=.�>J5�����[>,N�<����ݱP�|���}�<�W?>�s)��P�)8��H{6�iJ0=6�x?~�?h0�>��k?�C?Gd�< ���D�T�6a��\e=�>W?�mi?�>����7yо1া��5?�se?t�L>[g����ȍ.�#���?�/o?��?4`���}�<1��\2�h:6?�vn?ID��ݬ��Q*�/N=�Z>dm�>�?�4#�KbA>��_?oX(�#��jԻ�W��5��?7@��@,�T��m��=6� ?tN�>鑰�C�޾O�+��Ũ�v�E���?5(��擿2����)��G?��??��[(��	>UD_��I�?�8?�ξJT�/I�0�G�5�߾�t�=k�=��+����!Y	��oP�V��4׾����Qѽ겟>�h@k�=�7? \P�S����Cܿ7Ay�3��A	w���?�4�>����U�־j+��`����F�#C�4t��O�>��>����������{��o;�I���!�>�g�>ؽS�]!��r���v�5<��>��>j��>0���彾�Ù?d\���?ο7���M��P�X?if�?p�?�m?t�8<w�v�-�{�;p�T,G?��s?�Z?�%��8]���7�$�j?�_��vU`��4�uHE��U>�"3?�B�>R�-�X�|=�>���>g>�#/�y�Ŀ�ٶ�C���Y��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���F�!�A0=�QҒ�ü
?U~0?#{�f.�\�_?*�a�M�p���-���ƽ�ۡ>�0��e\�bN�����Xe����@y����?M^�?i�?ѵ�� #�f6%?�>e����8Ǿ��<���>�(�>*N>XH_���u>����:�i	>���?�~�?Pj?���������U>
�}?�ζ>��?��>�X�> #�=���%J�NV�=O��=�;����>]�G?`�>�[�=�H>���0��ID�]jR�����~>��7�>o�]?
�O?��>V��`k?�.#��� ��;��o��3�(����ҽ�,I>H�:>#�>��L�x�վ�g?����߿�3����1>$�?�B>��?�3� 4����Sv?��6>)�5��������<�
����?��@)?Fо�����=N=�>:�=�w�D��M��=�;>t}a?ˇ��ˬ� �c�W��>��?��@b�?C=w�S%?H�ξj/��h���C� ��ʀ��ӓ=��Q?(ξꃉ�g�?-�V>���������k���>V �?O�?#��>nFa?�v��.�2�=�!g>�Z(?;y�>6��=��о���>�.?��-�N���^�Ǿh�?$@^@�]l?Y�ʿ��ܿ��|����Z���3=`0z=7�>�7�P �=b��=K�潹-ҽS/>��>l�>�8�>ľ6>C*>���=�����&�\꠿����3�˸	�i���Lp�0T�91S��`�qh��I���ꍼ��������;z0���)�w�>8�H?2�V?�g?b��>ܓ:a��=�+ݾ~�%>�����=��>ME ?�'>?\0?�>$�����q��ur�O�¾ۼ˾Ք�>�(a>��>3��>��>�S½���<bg�>d��>�l9>��Q=��=�]���0>Dg�>�?�8�>�H<>��>Xδ�v0����h�jw�� ̽h�?�����J�
2��G6��H����i�=b.?�n>���=п����!1H?�����)���+��>=�0?�bW?�>S��#�T�50>��9�j��\>$% ��}l��)��!Q>Vj?��k>o>�s.�0k3�j.M�ޣ����>�%4?�ʾ�>:�&#w�*vH���۾r�D>C`�>�<$�zF��:��u�}���V�~k�=�9?> ?�Χ�j�ľ5�x�[U��<=�>��{>��q<��=n�.>����$�	��/>�"�=EK=�k;>�?�>#��=)J�> 񡾄�<��t�>�:>#��=�1<?�o ?��m�,��'䄾�� ���~>�g�>Aʀ>Bn�=/?��=�=^b�>�Qw>k!�>��`���+,���r>�D�c�`�����8f=�{��6�=x/q=�����H�g�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>��G9���䍿�WL�M�=���>ML?�׾�@>�8�^�n?� ?#��瀧��ƿaw����>��?�M�?�L��g����M���?�U�?�D?��v>���"��q��>uOO?YY,?�s�>� ��\?�ȸ?闋?��T>�_�?�f|?b�?�F�G�Q���)>����<r`@<��>�$>�6����L�p%���+�� Y��*����=Li_=��>�����7>���䑑��n���>S�">u�c>P��>~Y�>���>�&> ԇ;�G��&v�=�m���K?�4�?�0�.6)�pU�=�H0�sD����?�n1?񐁾�U����>�i@?p�L?�?R??��=g�/�̈���f���1ľ�ߦ����>�?�T>P)�<���=z>�=sR�>'�>,Aн�ľ�:S���=��?��	?���=��Q=�!?�9?E�>���>�[W�`ᠿ�F\��[�>��>���>(;q?�-?�_����3��f���ۨ�v�R��=Z9]?Yp?��>
ܚ�+���z��=#y��{Q��r��?ID9?}嫾��>�R�?�Q?!�W?��>��D><���>(�>�?�
�iL>�2+%��-�� ?�@?��>�3���꽊����0���o?�Y?�L#?�� ��{Z�)Vþ�c=�v���?J;;�<s[��`7	>6�+>�D\��]�=�%'>�=�$p�ĉ7���<���=)��>	��=��F�XŶ��a?8��=�־[�c���E�3 O�*v>�9�>es�%�C?��d�ի�����ӏ�������?���?�j�?��¾;l��C?R�?�)?��=`N�<����o6)�-4վ:u�]�߾6"f>���>~~��մԾ#���Vٸ��~��q�=F��a:�>��>��?�z�>�Z>fG�>y����:�}��;� ��}]�2�I�=�>�#�i��V��O}�RP��þ����q��>�"X�֬>��	?Գa>��k>M �>!a`��!�>�uk>��>y��>{9a>�_&>f>��-<�Q��3MR?__��4�'�h���h���B?6=d?�o�>,�h�͍����{?w�?�`�?m\v>;�h��C+��??9��>����g
?��:=�P��\�< 9��>���9�������>^Eؽ�:���L�yhf�3g
?�4?Ht��:�̾s}׽W��d��=Ǆ?�v,?T=0��%c�96t��rM���?��5���B������'���v�0G���g��Фv��{)���=o�*?��?��j�9W����y���D�YLd>g��>�h>F��>G��>p����-�9�f��I:�Z㘾�3�>,�}?z{�>w:E?y??�8R?ghG?���>�;�>���߸�>/S�<m��>���>�<?0�3?Q�1?|�?�i%?��T>�>׽����&)޾u�?��?c�?[ ?;?oV���
ƽC6+�Hh���|�Ζ�Tw`=^�<"i�O�T�㕅=�bR>l2#?�i�<��4�Q6�Uo�>a<?���>�P?%�`���;p�M���>�?O��>6Wþ�r����#�V�>H�L?���51=A�>�E=/�2<��ּAJ�=����}�<f5==o�H�?ݺ5��=�3�=W2�Xݐ=��<��/��4�k�>��?^��>�N�>�}��i� ����\<�=F�X>IS>�.>'LپMz��p'���h��y>8h�?�X�?��f=��=|m�=q��A������6�����<��?�A#?U T?���?��=?�e#?B�>�:��Y���\�����?N!,?P��>D����ʾq�h�3�y�?�[?6<a�^��F<)��¾c�Խ�>E[/��.~�[��;D��@��X���{�� ��?���?}A���6��y�~���Y��?�C?�!�>fX�>V�>]�)�T�g��$��0;>���>�R?Zd�>�$@?��?z^?�7#>�#��P������/�<g=^>nBT?��?���?�9�?��>m9>1�B�U{ݾ�����:���0���^���5>��Y>�@�>3�>�f>���=��>��Z̽j��3�&>�>�>���>�/i>d�>���>Qs>��G?g��>P[���������5����+<�k�u?���?؊+?�=p����E�y<���F�>Hj�?G��?.*?��S���=�ּ'ɶ�7kq�1 �>���>"(�>��=i/H=?�>3��>���>�=��\��{8���M���? F?qZ�=8�Ŀs�p�pRp�������;����b�����mf�G�=�8�����S����\��I������F精�����z����>Ci=�,�=���=�Į<i�ټB/�<��S=kН<��=��p�%�B<�s8����Ƃ������K<�4<=�E���V�w?/XO?��3?5�0?�Sx>�=�V�Hi�>|�r��??Y>!~��6Ⱦ5
7�� ��DW��È���(|V��ꊾ}>�U��]�;>�>ߩ�=���;��=֣D={��=���<\��<���=��d=�N�=��=���=�L>�Hm?v�V��ƫ�J�s���=��>�Ό>�>o?߾4f?Ks>zA��"�ȿ�t���p?}��?#��?��*?B�{�~>�HW��T�=H�>�5��i>>�Y]>��W��>:��>�}F�NG��|�0�l��?t�?��O?^�y�c�ֿi�3>Ў�=<E�=��2�/�4�K׊�"bz��e�j��>O��1E��x�K>�	��&�T3�ed_>a�>�n>�0a<�=0��x=t+R�O��=��>�W�;��#>��>�>=��k>*ج<U�=`�>Z9>��*>�f��zl���=|��=_%>���>6�?ta0?_Wd?Q0�>:�m��Ͼ�E���A�>�0�=�E�>nޅ=2rB>���>g�7?�D?P�K?y��>9��=i�>�
�>��,���m��m��̧�]��<s��?<͆?YԸ>LQ<��A�����f>��MŽ�r?�N1?�f?��>�p����������/�$~	����=���>d��!�<���=��9�V|ӽK�L>V?YU?��>!�>_�m>�.�>j��>��6>��潣��;�jջPݍ<�T=�Nj=#��;��j��d=�ͼ=l}<K�w��hf��x�x�K=؊/>���<H�=Qs�>XQ�=�<�>D'�=��>�>�B���l�f�=SԚ���O��No�?1��J���ܽĒ\>&Ph>"���F���-�>�o>��h>�s�?���? � >俈���>����EA�[o�d�&>��>f� �K<�X,_�&qB�����ɷ�>�*�>֡�>o>�$-�7>�"d=���0;4���>�.�S{��'q�����ş��h�m��_�C?�ׇ���=��}?�I?Cm�?l�>\����ھ;�+>�䁾}�=y�EVt����$o?g�&?�=�>B��,D�E̾�徽UƷ>�kI�Q�O�4���۰0�������m�>7�����о3��h������.�B�h_r�g��>�O?>�?�b�8Y���ZO�����A���j?Lzg?��>0??[B?y͡����%���D�=t�n?��?�=�?�->--�=B��E��>�2?���?�$�?-�t?G3���B�>�X�=��%>��c��^&>�#>6��=�<�=�z?��?�?��� A��!�fM龋"M�~w=��
>��>� >�w<>���=���;.΀=�)�>���>���>V#q>�e�>=�>�Y���	��B!?]��=�$�>��1?��|>��B=����ֽ<_�\� 8K���9���Q���ȇ-=<�x<�^w=a������>��Ŀ.F�?�%Z>r���?�y�Jڼ�Cm>|/D>�[ͽ�I�>�Z]>���>���>�B�>c>Y�>��->���>�&�Hu8�����>9�.ƾ�Ҥ>��7�$Ұ���� �˽D���Ǿ�5�ӿh��iz��̿>:�?�Ck>�̓�"i��< >!��>��.>�D?�tg��������=��?��>1.��袿\Y���[�K�?5��?��b>���>h}W?pN?�X2�rr2�"Z��\u��qA�o�d��`�[䍿1�����
�ZM��Ȱ_?.�x?rOA?�׋<�Cz>���?��%��ю���>b/��;�vJ?=� �>ń��+a��Ӿ+�þ�e��yD>"o?B��?8�?DoV�1z >���BAI?�@?�>�>�gk?�q?����?�0?�v?g��>�M?~�9?��>�/�>�q=������~>$��{�z����}
�Q8�=� =��K���=X4>��n�U��Cš<1c�8�!���(=��=S\�=F=���>��[?n��>l�>BK6? ���6�T����%?��5=����]l���Ƨ��Y���}	>~k?�@�?��Y?^\>ڜD��H�~�>��>�">�1^>�l�>��0�B���=t>*5 >�ʹ=e�,��h|��	�����f��<�1&>���>��`>vP���`>�w����h��h�>_�/�$J̾��6�3�E���9�\���U��>Et@?_?�O�=�4㾫�齗�W�fl/?DA?n/]?ڵx?��N� ��	�-��&��཰ݔ>���<�
	�1A������=��g���)5>�d�����gb>"��ϙ޾�kn���I�:�羃UP={A�i�R=�]��	־h\�ߘ�=�	>w����� ����Ҫ��-J?7Cn=�5��6�U�N���)�>���>��>M�<�[x��u@�ٗ��f&�=���>�q:>�򜼜�(uG�+��p>KC?�_g?C�?죡�ZJ��mI�݉B��/����J=�?�R�>���>�vN>�N��VžW>�&r��?�K�> =�>t:E� ]��ֽ�@���T�����>��?��6�?BoY?���>�&l?��'?~?�>��h>z׉�

��kA&?؏�?lx�=!�Խ-�T��9�'F�M�>*�)?hRC��×>q�?o�?��&?VeQ?�}?O$>² ��<@����>�i�>��W�f����`>��J?�y�>�~Y?��?O:=>h{5�1ɢ�w�����=mH>T�2?d#?$�?�׸>��	?Yۓ�;;o>=��>B� ?���?��l?��]=��>+]�>rɆ>��`=���>�!??W==?��<?��?O��>	߼'�=���?��1�<�܏�b<򼾼�<L��<��ὦlҽ/�����;;�D�IWl�u0�<���=�K�Q`����>+t>���gn2>�aľh܇��A>P���U��ˈ���7��\�=N��>o?[Q�>� �_�=���>�(�>���:J'?�)?�J?I����a�,4޾��P�8�>B?�B�=il�+����v�-�b=<)m?Y�\?��[��:���R?�Pt?� ��������mھ�O��k<?��>ۅ��@�>�?��S?�W�>{SܾJ���Z����NW���5�-N`=���><���.&�|Ў>�8?���>���=��8=W�̾=;k����sp�>�Ē?{߻?�R�?���=�r����N^�M���ö_?>E�>�⨾�W#?u���a�Ǿ�Ԋ��\��܌ܾ<X��д���u���؞�����i~�5g���i�=*j?�q?\lp?=�]?����-�c��5\��A|��V��!�z}��gF��wD���B�b0m��4��t��q�����B=-J���;���?h�!?�I�w��>����ܾ�O����[>ˇ��O$�{R�=�xü'ѳ=$��=��$��z���h���P?�t�>���>Lr8?6�V��sD��<�$�0��`�A�I>웰>�Л>�c�>�	���_�E3�N�Ͼzt��䪽grh>/�x?��A?ɕX?�Ͼ$T���n����׭�iE����n>�����2p>»#����%:�nGR�����w5�����z��E0�>��?iv�>�8�>��?JO�>^�����臐�R�B��(ϼ5YJ>v�\?o$?��>_��V$���>��l?���>��>xl��7d!�+�{�q�ʽ���>��>o�>b#p>VS,� \��h��׍���+9�3�=u�h?�u���a��Ʌ>c�Q?��:m�L<�h�>7!y�j�!��򾎭'�>#>x?��=��:>q?ž �/q{��剾s�<?,��>H5�b��(�>lO6?�>�C�>�t?ԋ�>��}�f�>��?lrk?c�O?IK?�&�>��>�[7�	ĽV�'��p�=<Қ>G�>>����o�:>�E�y s�>k��]�=�w�=	�s=���uȽ;��i�_+�=��=õ�=�Yۿ0K��Zھ�q�Ӛ��	����ߘ���ᄾD���#���V���Sx��@�@%)���U��"c������n��)�?��?$����ϊ��/�����������¼>zp�ˬ��d���������K�ྭ\��o�!�h�O�Җh��#e��E+?��c��A�������_����>%��>��?�^���D�QK/����>��=�μ���������uʿ3Z��;�p?w��>8D�E����>�1�>��>���>e���ξ;!�=bf�>'M0?�w?۴������ڳ���=���?�;@��A?d�(����i�Y=�F�>�	?��>>�0��T�x���J�>�#�?�׊?��Q=oWW�����/e?8�	<�F��7�Q��=d��=!�=�g���J>He�>���A�YܽN4>�<�>� ����^��ͻ<D�\>ڷս�A��zք?�z\��e���/�"S���i>��T?�5�>��=ȱ,?�.H�yϿħ\�<+a?,�?<��?��(?ȿ�D͚>a�ܾw�M?D6?���>-\&�s�t��g�=�!���h��}(V���=�>�r>��,����эO�	�����=����ſJ�6���%�1M>�J�8�b��q=pP>A�,����n�C�y�rۮ=�P>�*(>�"I>��R>(=�=��Y?��p?��>���=[�=#۾�?���>�51��9ᾑ	���ƽ˃���/�/M�H����������ξ�Pe�"͚�7f�_}������^<���(�%cc?��?I)<��U��	����̾����k���ڽ�f���U$���o����?��|?�;:��yW�X�����M뢽��?�/�����NY¾1k�=)B��tS ��H�h��h��q$��'&��t0?��?
���"Ȑ��()>4����=a+?D%?��h<ϻ�>�%?�R)�;� �[>�-4>��>ڂ�>�!	>�Ů�F�ٽ_?LT?߸ �c��ӏ>�f����y�:.`=��>�4�<6�`.[>3+�<ء���wW�y����G�<� W? d�>�@+����T눾nE9��p=��z?�Y?��>�h?<�D?:�<E��f]S����4=ȪT?�j?ҧ>;��h�Ѿ�/���6?gb?PU>؊a���^+�)���?�To?^�?�#�Z�}�����~��FY9?�cj?kQK�H̪���$�G��w��=Η>�!?��>�햏>rQ?���ݬ������/��?"
@X�@]!:���&�_��=f�?q�?�پ��f����������>7R?�\���.��
�����c�Z?�P�?�'?A¹���
�y��=p!c�^��?S�y?F ���V�f�9��T��]��y�A=]eX>R��E>��.��oO�V׾�*�m�U��RܽL٢>׊@&	+��B?ٽ������ڿ1�^��������IG?j?����վ&������+ׁ��a���Ҽ���>eA>A���f����z��9���Ⱦ�>oKݼ\N�>�P�Ca�������+<���>|]�>�ʄ>�?��5���
�?�����˿��������Y?儞?��?��?)<�Z����{��!ռ�]F?.Tr?Y?݅K�~UU�^�0�ôj?����q`���4���D�P�S>B
3?n��>>�-�7z=��>xS�>�'>h�.�-�Ŀ�춿�_��]Ϧ?���?�E꾥��>�_�?�+?�[�0 �������*�����"A?I�2>~�����!�D�<� ����
?�80?����`�_�_?)�a�=�p���-���ƽ�ۡ>�0��e\��N�����Xe����@y����?I^�?g�?е�� #�d6%?�>^����8Ǿf�<���>�(�>�)N>wH_���u>����:�%i	>���?�~�?Lj?���������U>�}?7��>�:�?�\x=F�>���=.����;.<Y2>���=�񽢤�>��6?���>`�>_L��42��+[�TVT��e �h�B��_H>�F�?4�a?�[%>~��<+5t�M�?�����Y�ֽ����_��|2��Z��h��>���>��@>�1��0���O?`0߾l�ۿ ��:��=G�>�1�=��
?u�ؾ���[�Y���c?J>�6�U7��&l����k�7�?���?�F?� ӾX��kb=��?�/B;X�V}�����k>�`y?V�h��"��^id��YD>�
�?ª@���?��A�I��>�g��AH��W�����=�F ����V?����-���[�>�pm>Q࠿"���~�����>k�?x\�?�`�>'�i??]��M5�:>��g>f�1?��>zpx>���?�?�uT?���C���	���}?�9@h@N��?�+Ŀ$�߿�}���Q�{\̾M �=Mw�=��v>�R!���=>v��=h,=��=�Fz>$(�>o�>�a>�v>b3>Ф�=�r����/�]U���؝�{@E��4�xڸ���W��鱾��:�s=	�h�ؾ.�p�F*�<RM'����:�3�w��+<��[��=pC?;�f?H`t?���>����=��B��g���M�<רo=�� >��6?7?��>ڢ���������Y�����bʾ)�>d�>1��>U��>��y>#9�*�>���>���>�L`>��>�������6>�Ң>9��>xt�>v<>��>r˴�,.��*�h��w��c̽��?[���J�^4��q2������^-�=�N.?�=>���6п���1H?z͔�S(���+��>��0?SW?r�>u.��>yU��>���H�j�^E>vE �ַl���)�!Q>n?d�f>s;v>E13���7��P�V^���~|>��5?���̧9���u� �H�l�ܾ�PM>�־>�G����r���<�~��\j��Jw=�A;?��? r��d$��'�u��`��I�P>(�]>J=z�=׌M>�c�90ƽ�F��2=�=	h]>��'?L��5p�>�E�>�$����L=1�>��p>P�="�=?!�?㧮;��<NO���\=q��>�z�>�B�>�%�=GnC�u">�[�>��P>k13=nY!��3U���2�k��գd��ؒ���阅�J�.��[<絼:�3��Y�����;�~?���(䈿��e���lD?S+?_ �=;�F<��"�E ���H��G�?r�@m�?��	�ߢV�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž5Ǣ�ɔ	�+)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ %�>���eY����V�s�3z=b�>��H?�"��!�d���?�h�?�<?x��@���Ɋɿ/�v�`��>0�?�a�?�vm�yϚ��4@�w��>:��?}�Y?��f>�۾�U��Z�>�@?�tR?�ܵ>Q���Z'���?i�?҅?��8>��?�en?�>�>��'��E;�㬲����%`�=�r�<�ߴ>3�>����NC�B���y����n�1� �2VP>_0�={I�>�u�V%���z�=���:�&��ѓ��>*&>�;3>���>��?m[�>
��>;5<����JI������7�K?s��?���4'n�S�<9��=^�^��!?�>4?��\���ϾŨ>q�\?࿀?� [?�Y�>X���>��2忿������<}*L>�I�>>=�>�戽5K>\վvDD�H~�>���>5����4ھ�)���H���Q�>�f!?�w�>Y��=ҹ?�A?��P>�+�>�Sj�E���\m���>��?�p�>B��?��?���x����*X��ife��/=��N?��%?H�>
���4��ppD=��>��)Ͻ�k�?��7?ղ�i��>��?�;<?�A?px>��������h��>x�!?�����@�l�%�7��*�?��?���>1���ӽ��ἒT�@���?c�[?^&?���l`��%þ��<�W�u� �1�<�����>9>,����8�=�>l­=�l���4�}�<u�=}�>e;�=��9�}򓽪t?k�=\R��dr���+rD�+M{=��>�ֳ�~�?�ؽ�5��4o��VP����ϽL�?ό�?uޖ?I���}Jo�X� ?d�?��K?ݷB>�_�V�LT/�����;�I,��$R>��>Y���e�������+�����(>�j5�Sl�>ˤ�>�w?���>f>�X�>�����=���̾����Q]��%�M�Z�� "�����3i�n�������̾GC��5�>�N��%�>j�?�<�>�MT>#�>vV�<j4�>�-�>��>��b>��w> g;>T]+>��=�Eƽ>CR?g!���(����2į��\A?�&d?���>��m�re��{k�N ?fd�?:�?h�s>��h�'�+��*?�y�>���>
?;C@=��»�؃<�S��>��Ỷ�ת
���>"Sս�b:�J3M��d�w�
?9�?�%���̾��޽֢��"�=_�?��)?E�*��lR���p��
X��?Q�Ϻ��^�L��ѷ$���p�k���0����ヿ|t(�s�$=��*?˥�?���A�l����j��M@���d>���>ܐ>E��>��Q>(�l0�<6_�f�)������>�p{?oQ�>�t7?�
>?�S?�XB?��>�/�>ɱ��ts�>6)d=�+�>t`�>�5=?��!?��$?�?Q?�[9>��#�D�ﾂ�׾$�?��#?KG*?O�>���>��f�?����D��#�۷k�^��z����M�<4.����=n�K>h�!?r0�=�4O�6�Ƨ>y)�>4��>�?+;Ra��Sڕ�2�1?�F?s-]>//-�<˙�V�0��><�?�hL�M���m��=k�=���"�'��>-�ƽ��=6�>d�E=9m�<��=l>Gt;&5>z?p��T=�)��~��>��?�N�>r��>矇�V� �v=� O�=S�X>'`S>�N>�TܾIn��梗��ff�{j|>�z�?�5�?[/Q=]�=���=�����������¾��<Iu?�$?BrT?F�?H+=?��"?�K>���C���w������2�?��+?ά�>���'�ƾ ���d�2��?z�?)�`�ձ��*�*�ľ��ν�>$)-���|�|߯��oE��X$�;���V�����?tn�?A�E���3����\���2c����D?���>4��>M��><�(��.f��y�@�@>Wu�>�O?�8�>�n??5w?��Y?��%>���iP���Q���1���C>@?߬~?g��?��|?��>Z�>�e���HU۾o�3����� ����<��D>�a�>G��>�>�;>����:��C����>&>���>��>�>�n�>�ߧ=��G?���>���e�J菉�X��y;��su?��?ʛ+?��=�Q�'�E�D���	v�>�b�?��?m)*?�mS�C$�=4�ռ奶��mq����>&9�>(:�>���=�D=��>��>V��>���i��h8�v}M���?Z�E?]t�=5�ſ�Bq�p�t�������<U����wd�����nR���=�$�����rX��-Z`��栾�����7��FꜾ�-���>�ĕ=�?�=�[�=CI�<�[ļw�<�:H=<�B<m|�<��w�J�c<�Y@�p������@-a��3F<n�:=���j궾S,q?��Q?i3?o+?0>&>ΑL�Ve>���=��?7>DQ�/L��	V�����XX��\) ��S����_�Ø���b�=M�=ѡ~>�_�>�b_=����$�=}d�<��s=l)=�.p;æ�<��:=���=Z��=^�=A#>OPk?wHh�Y���Y�c�T�!�U�?��>���>;|���(?�o�>�ޏ�VNȿ"��Utt?�c�?w�?�8?�2ѾHY�>֜e�jc=B�'>x3ƾ>[>�b��V��>��<>Ȇ����s�=��?� @j3:?����NٿpR4>}/�1�,>��;�L�.�Sw~�a@��ԡ�P��>�7e�&�ھ&M�>����D.*�H�O��{v>�F�>�á>�]�<=��c=Jͽ��>Y���8��>�@�>4x�<݁ݽ���=��x�>o,>�o�=��S>���=֕>p��=%t> ��=E��>8?yN*?��\?#)�>5�:��w���Y¾�8�>�23>���>_��=���>ܾ�>�5?��B?M�J?@Y�>��=���>�|�>vW���\�p(��$��^�轋�}?��c?���>~җ=�J ��W+��oK��� ��h?�p?l�>���>0t�i�����=��+������Ӗ=� �>�v	���`>��=8�轂sľ���=b�}>>��>�L�>�9�>6p>�o�>��>�l�>NL >��=���=��=�[���.>�<��<��m��fO�񸲽��<��¼}�%���E�=�����O�=��>n��=��>���< 9þ�>s���V\�� �=%���"M�U�p��z���(����+�U>*R>ӿ*�t��t�>��>�`�>�*�?V�j?LP>��:��=����f������j>~��=�<�<��n^�x�P��է�%l�>(��>T�>��l>�{&�D=�A$�=��ؾ�U3��8�>V���dZ������e�Ӟ��Ԝ���m��T'�j�8?������=D��?:�P?�?P��>�Y��t��;a>��]�'�ƻ-�zj�B5����?�'.?�0�>�2����G��F̾�뽽�I�>ۃJ���O��ȕ���0�c%����ζ�>!�����оi!3��p����/�B�Q�r���>
�O?��?�b�"Y���WO�9{�{i��Q?�_g?9��>H=?�|?�����������=�n?���?�N�?��>��>��򽑟�>>�?7*�?���?�Ќ?,��GP}>�=�=�>��,��>W>%�a> �x>�I�=�(�>�>t?��_��`����)�$����=�(=�ih>s��>�<�>��s>���=�,�� �=��>?� ?%�>�y>���>y=j=�K��<� �qA'?]�=�C�=��3?Q�2>4">$r�a@D>];�O!+��Tk��`)�K��=�_>�8�< �>�;�=��?,~���`�?��C>�� �q#?z.оaTN>�r(>��>���)�>���;��>M�>���>^�=��>�:@=�޿�V�>o�,��O��o��&�O�}����>�T��`��G���(��=E��о9�!��\�����'b*�Ψ"�e�?	z�=������J�X$�>ơ.>"��=��2?�;*g��>�7?�P(>_���#��Ls��������?���?�J>u��>��Q?��	?�6���0�8FQ��zq�d�D���^��W��򎿠X���
�%�a�_?b?��}?�kB?�h���Y}>�Wj?l����p��Ve>z4:��b9���.=B��>w��$�l�vؾ�ƶ��н7�>��a?��|?��?؞t�\�>�*�F"0?�"?0?�0`? 4J?�u����>O��>:w�>�~�>x�+?��+?S�?�*�>�#->��`��=�^����c������=��J�;f�>l$.���M>g��=�f<�W=���= D<<��x<��I�7�=��=�|�=I��>�{\?���>�F�>D�6?����8�����h�,?�b6=�߁��f������.�@7>��j?栫? �Y?��b>��A���B��\>e��>��%>Nr[>�Ұ>W8�@�C�U͆=��>��>ta�=�[C�~��bA	������c�<��>�A�>:��>��,�@�;>1ҟ��9r�ѡa>S��D��M�R��H���2��b����>:�I?��?�K8=C������7�e� �?�XK?�T?�wv?�Z�=�~޾�A�H\M���/ӕ>�1�8��I��'�����0��ȼ<K�Z>Q���jˠ��bb>����M޾��n�+J���羆�L=6w�8pU=���վ����=
>����� �?��ժ��(J?�k=Ym���GU�Z]����>���>�ή>�Z;�<]w��@�F����^�=~��>��:>�������oG�P.��2�>ZD?�>]?��?f<���Sp���>���5����s�= ?"��>��?��M>,'�=F���Q���d��FG�NX�>@�>�B��DC��閾i����M%����>N�>�7>�V?FOU?�?��R?�^ ?�r�>N��>�z������F&?ى�?a߄=��Խ|�T���8��!F�r�>y�)?��B�Rח>j�?��?�&??rQ?|�?v�>e� �4)@����>�^�>1�W�d���`>�J?+��>b>Y?Ӄ?�->>5�Mܢ��m�����=	>��2?{7#?��?ⷸ>ߡ>k��?q>~��>�?Fk�?j�?��_��Ҡ>Y��>t�>��0��%�>���>ɤ?5�D?X�n?�??�A�>B1C=�]����'�=��ug==�<���:��@=�G��Q;���.��@�=7��j�8��P�����O�ν�@漝~�<7��>�it>#����1>�uľ��<@>.0���E��!ߊ���:���=��>V�?ᨕ>�#��=;�>�'�>����&(?2 ?�Q?��;�rb�&]ھ�,L���>��A?�L�=
�l�����^�u��bj=Mn?�?^?q�W�td��s�l?C7[?�J��v*�ۃ�]r�����[?��?����h �>�?�%�?��>����\�y�6��YK��=���=�Jx>
P�!C����>��4?iS�>�t�=��=�ɪ�Cb��Nܾ+��>�?�ˬ?V9�?ܘ�=��Y�^��p��^����[?B��>/0��[}#?H�^< <Ҿ:�������9e׾s驾*ﭾGD���?��%2�|x�nsν��=�?	h{?I�n?S]?�#�E/l���^�#���x�L�����
��eC�E���H���n��%�����ǫ�J�=��8B�.�?��&?��.����>����̍�;�C>���a��ۚ=x����XL=s#h=�Nd���+��r����?�ͽ>h�>ױ;?wH[���>��1�n8��<��`�7>� �>��>���>��λ��/��)��;;�釾�zн�X�>�[g?*a=?��c?�����?�#k�pR��KA������">x8<>)ӌ>9�L���.�ކa�o�m������q����F�)>�*&?-)>��?���?�G�>y���O��t���H;�hp�= C�>`�P?��?B��>e�۽{�2����>�+n?l��>�)�>�V���� �O��T]��SJ�>�>( ?Q1�>�$�s^����Bw����7�lU�=Qn?H�|�Ff��g{>ĩH?��;<�	=�ţ>e�c�x"�=y���kN����=�
?V�>މJ>͹�ˤ���u�3���%?Hz
?�'���p)��l>�!?y-�>줟>�X�?���>��¾��y��?��]?��K?ϓB?�-�>8!9=�D����Ƚo�*��v5=>3�>3�c>Z}�=��=��p�O���ՙB=�G�=��������Y�;�м
��<qb	=��3>��ۿ(eI���ӿ��T�2��Y�y�mn$�ДB�
�N���־p���-�o��hܽjQ`��8G�Ouu�}^���.|�Lx�?�[�?�ӑ�Mg��=�����	�#��>ҩq����ϾX?��+�����fɾ;�*��cT��c�a���!?l7��تǿ�d���Ѿ��?pB?�w?��	��e(��;���>y�<��l��ԙ�tο����ێ\?���>-T��ج�1��>�H�>� J>_>՚��5���v�<�(
?N�,?�>�u{���ǿ
������<V�?��@��A?��(����IV=���> �	?q�?>�01�<��ⰾ'P�>�9�?��?��L=��W�y�
��me?�<�F��޻�=D]�=S�=���P�J>;h�>���wA�#�ܽ�4>(��>e�#��}B^����<�[]>��ս����M�m?}B��l��A�Ex��ռ��Q?V�)?�X��79?_�V��(Ύ��	�h?��@�0�?VN?������>׻۾�:?3�=?���>gK\��W9���%>@v���;��9Ӿ�O$�q��<�p�>8b�>��<��'���W����1q>�a ���ȿ�/�2j1�[�=��=��u=���<��=�G�dyľR�,�����>�2>���>�c>�8'>�K>ob?�ƒ?�$�>l�=�G��HR��6�辖�'�*�U������Vھ�Δ�<���)��,<����Ǥ4�'��1�ľ_wH� �=	�X�'x���9�|�U��(<�~�4?�r>�b��]Hf��������)��=���෽�nپ��0�ͼl��Z�?m<R?=����dS�r��[�����4���D?�O,�̰��ٸ����=�h/�*�f�@�T>��]�?W�9�$�D	E�d�<?N�&?Q����vs�^9�>��s��5��+�,?��>w�ݺ,��>�'?����~.��>>��="Z�>�'�>Z�>R��'�b���$?K3k?fT��aǆ���>xGھ�㠾H�ྲྀJ�=����(|��UU>��>{��h�����Ͻ2��(h?�=�>�q�����0�5���ۼ=}z��?W�6?���>9[?��k?t�d>��L���b��-�؃=�<?BՖ?q;>�6ɽ�D̾1�־��:?"d?�(�=n���ɾ�`I��V�/�B��>�Aw?y6�>��N;xW���h�w�đ?�!j?�%W�����%�� ���>�B�>���>��)�9�>�/?��/�T����u��˛-��b�?�x@0��?��B������;=d��>(v�># ���㷾E*��T��jj|=�� ?���D2q��(�9ڽ�+E?��?00?������p}�=�	�3�?�Fu?�����3�g#���r���о҃
>�D8>ì��� ������'��4��w������\錽s��>�q@�1��
?5������/�ֿ��~��(�������1?�`�>Ӣ�<�Ծ]���������b��C��k��:�>ĺ>먕��*��P�{��y;����C'�>VY�J��>��S��.��՟��42<��>K��>� �>1���N	�����?�b��/ο2��������X?[f�?�g�?xg?�=<��v��{��1��5G? �s?J0Z?�1$���]��P9�,�j?a_��lU`���4�MHE��U>�"3?�B�>;�-���|=�>���>vg>�#/�l�Ŀ�ٶ�4���K��?ۉ�?�o���>k��?�s+?�i�8��V[����*�[&,��<A?�2>O���o�!�)0=�Ғ�μ
?5~0?+{�~.��_?
�a���p���-�s1ǽ(ɡ>��0�N&\�������?Ze�����ty���?j`�?��?@��#�O1%?^گ>ܖ��E"Ǿ�l�<7f�>/4�>=0N>��_���u>�j�:�td	>Y��?�z�?b?��������"T>�}?M��>*�?I=
>�?�>ᬛ��SѽuT>�=�P��1�>��>? �>�]�<�$�(,�-�J��AL�: �)�7�<�h>&�u?�Z?q\�=]���M�=�@*�z�4�h�^�,����n��G���;���^H>���>���=$�^�q)����>1�𾐼տ�*��	�>��>c,�=%]�>LGž���� <%��0?A\>��!�M{���0��q*I���?q�?��?��ƾ�Mҽ�G7>���>I��=҄"����Ŀ��=��>��P?&6	��V����_�R�>s��?l�@V��?��>����>n�ݾc�����Vc��ߤ�]���+8?`[�����=-�>���m����n��^�i���>�߲?s#�?��>wg?��d��t<�	�Z���K>�=?a?�a�=���Sî>jz�>C��ݝ�S@žtgw?f1
@f@� K?�M����ܿ����_Ǿ�m־cr�=;e>C.�>Qc��4�!>(�8=��,�ڻ!=W$y>a�>�1>��s>&�5>.+>`�?>�݃���!�_Dɿ,����'��s
��+�r��'z�Drf�|��q���ž�@ϼ �����Q�u�<�u�7���὘�v>:�*?�Q?�/n?�d>`�=GC�=�J%��w4��j�WX1>9�7>0 ?�R8?N�?��|���־tp��������.�����>���=ۨ�>.e�>@�>�b��7=J8K>�T�>hu>�g>\Ŷ<7�ż��>�K�>B��>+��>5�;>��>gϴ��4��nh�Rw��8̽g��?�;����J��B���S�����/'�=+3.?9>E��e/п�P6H?ӭ��^-�B�+��o>I�0?�$W?�B>�3����U�TM>T����j�O� >z� ���l��)�5yQ>x?�KX>�n>��0�B�6���R�?ի��l�>��.?g���֕,���t��J���߾ѱX>�j�>V^�;���D듿��{��(p���R=�\;?�j?֒�f׫�B�V�=���ǒ^>��c>�.G=�S�=!�Y>����(̽��F�e�)=��=?�b>�?�)>/��=�?�>����K�#s�>kU<>��$>X@?�O$?����%́��7(���z>���>�Ѐ>I�>�J�](�=���>sa>���	���u�;�p�[>�Vs��a\���e�A�|=X����=�f�=Ӵ��A9��.=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿi�>�s�.Z��-��#�u�ĵ#=���>X9H?&S���O�[>��w
?{?�a�ܩ����ȿ�{v����>��?+��?��m�"A���@�o��>���?�fY?(ni>h۾^Z�)��>�@?�R?F�> 9�H�'�d�?c޶?F��?��R>>?�?"�c?#E�>����I������?��<C�=P.�;��>��I>:����98�J\��݁����s��0��Ze>��=h��>h�)�̻����=q'���P���$�<� �>
a�=�ɛ=�V�>�
?�?G�>�?=�ǽ�����T����K?}��?����+n�)�<8��=��^�"?�E4?�\�[�ϾoӨ>��\?���?R[?�^�>����=���翿�{���ɖ<��K>A0�>�F�>�)���JK>��Ծ<=D��n�>�ϗ>M����;ھu-���E���?�>�b!?���>��=�0,?�=?� g>"B�>�3��*��6�f��>1?}�>�#�?P-F?>O���6��.��T¦�ĉV�2�_>vĉ?)�
?4�>7����}��=p�=�{n���?8��?Le=��>DƁ?�>D?lY�>V=��4��;�4�<!��>vZ!?�]��]A��&�Q��[?8�?��>��Yӽ{eؼ��8����?F\?|c&?�/�"�`�Q�¾4-�<R�+�{M;��4<i�5��>�$>�D��M �=).>���=TKl�F{5��d[<0��=C,�>X��=�a6��(��5,?��G�T탾P��=@�r�XxD�-�>,�L>�5����^?ޓ=��{�C���e��TuT�?�?-��?\�?9���%�h� =?��??�
�>���eu޾���TZw��x��i��#>��>u�j�12�J��������8��49ƽ�^%����>p �>PW	?���>��P>QT�>XC���)�?����_�1���3�U'��������|�����r�¾Vs����>-B���>L	?ox>D >W	�>�q�;��>M�X>p��>�B�>z�R>�`1>�>�i�<Z伽�\R?�z��&�'���89��J.B?�d?�J�>7�g��r��ݱ���?���?{K�?��u>�h��+��T?XA�>����n
?��;=[���]�<�#�����X�������>�׽WR:��]M��f�x�
?LI?s�����̾�Qٽ�N���3>��}?5�1?��(��[��cd��^Z�H�A�>�$�s24��:I��O�]��d������%����!�s}2=�#?҅�?�/���ľ�g����w��`���>H��>nA>Y��>-z�>v �-g,�G"\�z;� Y��?��> �?@֑>�I?��<?1Q?��J?p2�>沤>f�9�>5�߻���>�n�>�8?�(?Ԃ.?�V?�*&?�	O>7�Zp �pݾ�:?�r?l]?��?�k?�������
��罆9��o�`dJ�[�=b��<�籽�?Q��==�0O>�m?�� �8�Ʈ���&k>�q7?���>h�>ʷ���Ԁ��V�<�Z�>�
?���>� ��r��R�:�>ං?���	=��)>�y�=J����¦����=8Wü��=Ƀ�Ol<�h�<H$�=)��=�c��;:��$�:~h�;���<t�>u�?��>E�>�A���� ����4[�=�Y>S>�>CDپ�}���$���g�Xy>�v�?�y�??�f=�=���=�~���T��%��E�����<�?lI#?kVT?T��?��=?j#?a�>�+��M���^�����Ѯ?�,?p��>���øʾ!���3�3���?�[?�Ha�����=)���¾�pս��>^@/�I~�����1D������}����?��?;�@���6�+d�tǘ�PS��w�C?d#�> n�>s-�>һ)���g��*��;>`��>^ R?y�>�N?�z?�[?v�H>�d7�Ҭ���*��g�[g>Z	??@6�?(�?�+y?�	�>v>�Y2�(�㾠����i����)=���[=��X>e%�>�7�>[d�>@��=U�ɽJ����<�"Ҧ=$ a>\B�>ӈ�>��>?Lt>�<��G?���>Y����q�������I�<���u?�?�+?;=�����E�R>���R�>2o�?���?�3*?��S����=#׼&ܶ���q�U)�>f۹>40�>~ݓ=ԹF=�a>��>���>� �T`�0o8��`M�4�?�F?1��=^�ſ�q�xn�2<��.<1<�n��:�^�鼖��j]�ɤ�=�(������-��rFY������6���J���g{�:��>�D�=��=a��=�2�<X��Qg�<��S=���<�W=�Ge�ٔ<��.�M��#���RAm�9�_< _L=&�λ�w����w?-N?�+?�C??��>�$>֛�\1�>��+��?�ja>����ͺ�>�9�:���cb��5ݾ��о�`����8�>��W�{��=��>o�=}i�<V�>�O�=���=<�2=q'�=��=�O�=�b�=��>� >�L?�[�xp���������;��>��b>-�> 
���3&?_�������!Ͽ��ھ�h�?Mn�?�H�?�t?�o�>�Ѓ����=�>KF���&>(%�>_��=X>=��>7P�������ý
e�?Ɉ@h�b?Q􀿳�A��>oj>'z�=k�I�y�-�����T�����?�?�w��Ϧw>w�2=�<�*W��惫=�BZ>E��=v����U�=%ՙ���k=�z=��>��D>���=.ji����=��z=�)>0dZ>�<����FP0��5=w��=�k>��.>��>��?�p0?Ud?>�>ĳm�[�ξ�d����>���=d�>�U�=��B>Fy�>��7?5�D?�K?�P�>,��=B��>��>=�,���m�Vj��⧾���<��?#І?0�>*V<WA�Ï��^>�oŽ�]?�D1?.p?��>A&�Vh��m>��`>�����7�=z��=`����=>�X�&�'�R��O�>��>H�>p�>�Bz> >�!>��>>*>]f�y��;�6�=K�.��;>�؂<��߽sSq����vͽ�h��V�=+Y<=Ы���d<%��(��=���>�;>B��>h��=���aH/>������L��Ŀ=�H��-B�s4d�'G~��/��O6���B>�;X>P���3��U�?��Y>_o?>O��?�@u?�>."���վ�P��>@e��PS��Ӹ=�>l�<�'z;�Z`�k�M��zҾ��>��>ߢ>s�l>��+�"�>��u=���<5����>�f����	��3q��+����!�h�p�ݺ��D?7��g��=�~?c�I?�Ώ?݂�>練�j�ؾr�/>�����=z9��^r�s
��(?U''?9�>���D���̾I1����>_xJ��vO�5����0�t��x���v�>fh��H�о�3��`��O��k�B�
s��-�>��O?�ܮ?#	b�E���O��h������#?�,g?�ԟ>?[?�v?�������򌀾 ]�=ͷn?/��?�S�?�P>A'�=e��|��>:�?��?8�?:5�?E)���x�>���=H�*>X�&��";>��;>Ǯ=P(�=��?�?\��>D��n0��}��f	���s��a5=_.�=�͙>x)�>�*�>��B>p��=xz>G9�>��>��>��>_�>�
�>Z������d?h�=~82>�/?O�>Z�w<��!��*�=��\y���Yh���}��=t�>T�>�K>;�8t�>�¿�1�?��>�l��W�?E%�G�=�x>���=HM	��?�!�>&Y(>�NT>�kJ>.-�=���>P��=.`��ؔ+>�.%���;����lD�9WҾ���>z�T���̾��1���2�z�;���������b����.�~�ü�	�?��4��b�p$ ��b2=f��>z�">��?3����7���o>�!�>i�I>$�C/��a����R־2�?X��?�6c>��>h�W?�?]�1�3�sZ�r�u�m(A��e���`��፿ۜ����
�g�����_?a�x?yA?�S�<�8z>2��?��%�xя�K,�>G/��';�L<=_,�>V*����`���Ӿ͸þ38�FF>˔o?�$�?Y?�SV���>��u���f?�_D?��E?��d?P�Z?3�־��>���>��	?�#?|H>?�
?W%�>O�Q>���=!�<U6�=qs\������M�>��?����Ή=v�0=�1i>�.�=��=��=�o
=�<�=�)����%�=�Q>9[>���>�7]?}�>G>�>l7?e���7���Hy.?�b>=͂��Ћ��
��T�d�>4k?e�?XDZ?H�c>~(B�D�C�y�>>V�>Z'>	\>�ȱ>���`�C���=��>� >[&�=�Q�񶁾
�	�����G�<��>2�>��W>B���-:=o���Z�I5�>+@�(� �-���L�B�e��mվ2�?��n?��=?E�}>u�ݾZ� il�V{?�^?!�[?�
z?l3�>M�N�_��������Z�>���>�i3�nX��y���>��5�jg�><��`��~dR>�����ھH�j�mL���侩q�=Cv��{=�i	�ъ׾Oǃ��;�=�:>D-���0�����㩿:�J?T�j= M���^��*��� >��>�D�>��;��Ő��<�ʖ��]��=��>��3>��0�.龗H�B�g��>h+?��u?�I�?~��V`��h8��<��ހ���=*�?�^F>��?r�5>�f�<�ƫ�1)�i~����O��>�v�>,���5V��d��<W߾� ��N�>�?U�=�	?�J?cd�>W�]?L#?	��>��X>��;ɚ��.13?�<y?�ռ^�������"�"�"��a�>'�J?�o���8+>���>�	#?�3?�M�?f?����;�뾢�B�KW�>��>��k��[��Uk�>�X?�N�>�*?�]�?��I>C�H���M�tو���>�8>�fL?Tb?�=?x��>4�>������=��>�`c?�Ӆ?B n?R�=�&?��1>��>e�=�ʜ>̱�>;�?ðM?�s?�yM?-��>NQ%<�K�������!��t<�8<J�9<{�=P.���$�,J�gd�<��;/\ּe��QS�H5��*�=v6�>\�s>�����1>j*ž�3��T!A>����uq��yq����:�q$�=���>6�?�|�>9K#��P�=XE�>���>���8(?��?S+?D$b;FSb�ɷھ�K�MͰ>fB?�j�=�l��w��#�u�g�g=��m?y^?<�V�x���=�d?�bX?\��j8�1��}-b�y߾��O?kp?��_�g�>��q?�sn?�k?g��̌c�����7Z�Gx�����="v�>��� �a�"'�>�T7?c�>9L>�>>�}߾�q}�P���~??b{�?��?B��?q>�e���ۿ����g ��_w_?���>��*�#?���ٵξB늾s�����'���������h񥾬�'��~���Խ'з=R�?S�p?�9q?@`?����ee�Ҳ`��&����U�B,��H��B��D���B��^n�M������`����.=�_�,�5��n�?y�Q?��O�v
�>�x��C;��I���HE�>|7־�}���7>��ོ�=��C���KT��M���8?.o0>���>0e.?c�S��N�%^:�ʒ(�X ��=�>��>.��>tR�>0�<���j۽���(>ɾ��D�@��>��U?��@?��{?�&�)X������'����a���\\f>^��=��>RӉ��e��C-���2���M�F�������(�+��>��c?M �Ȝ�>�!�?��E?K�:��~�������r����<��a>1 [?9p�>���>g�Ǿ=X3���>��z?r�>UU�>�h�R�7�����5@m��`�>Y�>pv?�m�>/G�̳S�k1��Q,��1�n>>8q?�^�������>��L?�佫��=/;�>��>2�����S��9>d��>e
>�}>�!������x����EH?��?&?�Z�2�L�>y�Q?ڳ?���=�Y�?��@>[i*�,cD>�>5ш?��+?:σ?�T�=�e�=`�&=��Ͻ�hL�$@�=c�=V5�= �=�Hٽv�"�sϖ�ZGT��q�='��>�P�?�D�Uy�ɯ���<�`u=* >�Eۿ\TN�ZӾ����I��I	��>���3=0��n^�������MR���>W��F�,�Q���N�8�t�[W��Y�?��?�5����i��畿��n�i��Gm�>��&�Z�>9y���: H�`�Ⱦ��t������4�gz_��rt�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >KC�<-����뾭����οB�����^?���>��/��p��>ޥ�>�X>�Hq>����螾�1�<��?6�-?��>Ďr�1�ɿc���w¤<���?0�@�V;?
q�y�� ��=S3�>e?�b>;0u�P����;�?û�?��z?�+w�BP��@ڽY�?�>�{8�������=�2>!�=( �d�p>�>!L��?���$��q]>��<>e�= ǰ��|���/�<�>�Ļ=����)Մ?,{\�tf�ϣ/�	U���U>C�T?�*�>�5�=��,?*7H�r}ϿQ�\��*a?]0�?ͦ�?��(?dܿ��ך>s�ܾs�M?�D6?��>1e&���t���=�DἏL��/��('V���=��>��>(�,���P�O��G�����=����ͿdB���2���	=�"�12�1�<.�%��	��bξq�N�z？)�=&zp>��L>�%�>��>�ˏ>�k?=s?���>cb>���5��5�ھ�I�<K���S��\>���3��,�S
��:���:��_#���!�h��T�-�7 E<|Q�Ĉ�b?�$e��2��"9?���=�*��7�8�(�y�)�Ⱦ>��^���~�*͕�vL(��n�I��?��7?x�y�B`�2o#�"w�=3�ͼL�V?�ܽ;#��Ƃ�aY�=-����;,��>� 1>�Lɾ�>�u�E��t>?e�?�л��g����=>)1~=�� =��?�?�08���>��X?�����e!�]c�>~�>���>kĺ>�B�=��ž�K�C8C?Z�]?��ٽ�ݘ��R>kl�������%<LI?؋��;"=�kȽ_|@;,E�H��>w�=�s��'W?ڝ�>z�)���-]��T�A==L�x?��?�,�>�{k?	�B?��<`j����S�� ��Vw=t�W?*i?�>����G	оM���(�5?Тe?P�N>Zbh����i�.�$U��#?��n?^?7x���t}�������o6?��v?�r^�`s������V��=�>�[�>���>��9�wk�>2�>?9#��G������Y4�Þ?��@���?��;<� �q��=�;?p\�>�O��>ƾ�z������̔q=�"�>����uev�����Q,�K�8?ڠ�?R��>ϓ�������=�����S�?���?�a����9;���Ol�/t��D-�=&�z="�JO��Vg꾀�:��=⾦�������C�����>0�@��/���>�tT����|Ϳ&�������圾o�C?d�>!Y^�S����l��lt��bS�51��dk�O��>�Ww="��������f���+���b�?�Ķ���S>��ýҾ�읾�M�=1�>���>%5>K������?����Doɿ�ꟿzݾ/L?�,�?��^?(L?6h���}|���?��g��2?y^�?�f? bV�Hz� ���j?J_��U`���4�5HE��U>�"3?zB�>I�-�ǭ|=�>��>�f>�#/�R�Ŀlٶ�����=��?���?�o����>u��?�s+?vi��7��Z[����*�U�+��<A?�2>(�����!�40=��Ғ�e�
?/~0?�x�F.���_?6�a�R�p���-��ƽҡ>l�0��/\������Ve������y���?�d�?5�?��n�"��%?��>{���_Ǿ�U�<j��>>�>�zN>��_��,v>m�� ;��z	>��?pr�?Or?M�����pF>z�}?f�>�F�?}H�=DY�>\��=�0�����D>E�=����>��>ЊJ?�,�>0 �=�9<��,��fG���Q�T3	�c�F��>��a?��M?X�x>�I��O�6�����ҽc/(����d7�%]�R��Ϣ4>_�<>�>�-���ɾ��?Lp�9�ؿ j��p'��54?.��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>;�>�I�>C�Խ����\�����7>1�B?Y��D��t�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�b��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?TQo���h�B>��?"������L��f?�
@u@a�^?*�7����:ϥ��7��A>�0=��`>�k{����=�B=,T�;[���Ay>q��>�ӛ>w�>���>���>o��>�&�� ��ᗿ�z��g�L���!������N��h�+��b�!��ꐾ�LK�i�f=���3��[���������=�`T?�8R?��p?���>0Gp��S#>X���=��<@����v=K��>�1?��I?�(?0Ȑ=Fj��@d����Ϫ��ރ�J�>��L>Ԟ�>��>���>k� ;Z�J>�4@>灀>cT�=@B=����j=�M>N�>+��>Ƽ>�g>��j=�_��)���/r�+�p���ż�?�x����n�+~�vM����!+�=��?��Y>h�y�P�ο)5��;�E?�6��F����S�K~�=i�0?��[?���=�5���?b��+>��P��u��=m0B��rZ����;�=ڤ�>�r�>M��;�5-�"H����|VQ�T�?t�?f���:=[c��Oz���`>�~>�>�@
�툤�0��,��	">�9M?4�?����@ʾk���.�0�>y��>��B��Xc>_�>�`߽�t=�ל���D�@�->�u>�L?PJ>R$>LK�>D:���J�H�>�#S>�(�=ɰ??��"? ���oq�V��7j<�omb>�6�>:@:>�">b-=��9�=�'�>��8>`�����v���0�N�Y>.�*�ôF�*�:�%wd=������=p��=dk��9�L�=p�~?�}���䈿��\Z��mD?w,?c �=�G<��"�y ���F����?/�@�m�?�~	���V�
�?@�?w	��^��=)x�>�ӫ>Qξ(�L�m�?lƽmŢ�;�	�,#��S�?K	�?��/�6ˋ�l�`9>�^%?��ӾPh�>{x��Z�������u�v�#=R��>�8H?�V����O�e>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9�~�'���?�޶?֯�?YhW>��?�	?��>���>jUI�c<��	����>�-
=�?�K�>��=���<Ԓ�歠�d҂�^?�����>�=޳�>�C��G\����>�A�����U�<�Bz>nh>�6>���=ߑ?a��>U��>��>���c=�@��WX`��zO?%�?�����f��7=�]�=�v0�+0?��D?�����+j�>kW[?tց?�m?W�>��yu��:��]����#-=}n>Һ�>���>Ln
:��v>���'&��Ù>�z�>�5=���<Y�snl��5�>�#?�V�>��>k�?s$?ԉ>@�>]<6�K�����K�>��>�վ>�v?N�?�?����^�4��+���N���WU���+>`As?n?�a�>�����L0>N�S���̽�n^?��x?\N�n�?��?��F?��?��}>�@��h��&=b��><&+?E��к_���=�|���4��>8&?Ӹ�>�X>�g���c�1=��1� 8���>|*?�;/?=���b�|��!�9#=Oy��2a<<ec<�E<��U>F�>��D����!�>7�I����=�۴<�Fλ�D�>`;=Y/�X_l=�<,?o�G�\ۃ�
�=H�r��wD���>	JL>��N�^?Rk=���{�����x��q	U�� �?���?Ck�?S��"�h��$=?�?�	?r"�>�J���}޾��ྖPw��}x�w��>���>O�l�W�*�������FF����Ž4�@��>�I�>=�&?h��>��_>&�>>0��x�&�����Ԟ����U���xx1�����	�c����R�?��*IھK�.�๖>�C\����>U�?f�r>��>���>�p8� �>�@,>�	>���>�6>�">dm>Ɍ�=��<l]R?��� �'�5��pg���B?-Zd?nD�>}�b�Ɗ������9?}�?�p�?��x>� h�~`+��N?n��>w��V�
?�4=1,�6s�<�����E��f��D��Փ�>D�ٽA�9���L���e��}
?Qh?���	z̾�qֽ�>��Ͱ=��?7?kM)��zS�Kt�tj`���C�\Ӽ�ݽ�W���9���h�����n������Z��	��<͟#?���?��"��� �9�Q�-y��@�*��=S� ?�&/>u�>3�>�����nE��RW�;}��َ�^�>�u�?��~>'lX?'UE?R�2?��6?��?֠�>:c⾍�?�r����>�1?T� ?$1T?o%)?��?=�$?��>@9�<2��D%��{ ?Dc�>R#?�A?[ ?&z7�p2)���>����㟾��̽*b2>,3>\�"�-b��� ���>�X?�z�7�8�*���Rk>H{7?�r�>���>Y���)��,8�<m�>}�
?�B�>� ��}r�#d��Y�>G��?����X=A�)>���=���Cnغ�G�=B0���ؐ=S>��Q};�� <�}�=3��=e�s���|���:g�;���<gu�>��?���>F�>�:��	� �����?�=<Y>^�R>�;>W/پ�z���$���g��Ey>Q{�?�z�?ޡf=���=��=�n��JH�����>����<ǘ?'H#?URT?锒?��=?�l#?ʶ>�-��J���\������ө?�R+?���>2
�-�ǾH}���/�,?]?�>Ɩ[��8��`-�T"Ⱦ�ڈ�w� >�V-���v�5���H�K-��i���[��?�?�v�?�}ü�+7�d����񗿄���#@>?��>̽�>wl�>fv(��)b�WL�F(>���>��N?܇�>�O?�{?�$[?X�T>	I3�Y���%���N�M�{>uNA??�?�*�?o�v?���>v�>�`���׾���P+)����+��8�.=��S>ג>���>p�>UO�=���Ӈ��>=�,�=�L}>�g�>+J�>�M�>�k>��=%�H?v��>��þ
'�����A�~��*��s?���?��)?�>�<���e�D�wm�K��>���?�%�?�|(?��Q�F��=�ȼ����X�t���>�k�>g�>+$v=��D=��!>���>^��>ȸ�(��e�:��2$���?��E?��=�/����d�Mz��[(<��E�=�<*��o���#z>�А��˰>2����:���)��G��˅���M���T���A,���?���-R��q�5>��=��=�߇>�;O�5<��=�A�=n�v���-=��=4m&��0����=�㙼�j�\!߾4Rt?{I?��0?�.?1&�>�+q>�a�����>:��l�>M,>�P���ľ��$�����jh����4��v>m��߰�5N�=&d��5�?>:P>w��=S��=��>�R����<=�N�NF<ٶ�=�l�=<r��>T�5>6H>S6w?����~����6Q�uq���:?xD�>���=��ƾ�@?��>>�3��w���`��#?���?(S�?��?$|i��a�>m�������(s�=����B2>K��=0�2�,��>� K>����J���-��1�?��@M�??{ዿl�Ͽ@i/>�)>y��<|![�ޗ<����}^p�˓9���0?1�6������u>P���W�þ�҇�ǲd>�>{cL�e�_��M�=쿽��W=�>�$�>M>�W�=�����0=�d�=ܱ>C,>��z<@��;���/�D=�g�=��S>1iy>�_�>�?>�1?�d?\'�>�gl�a�ξgɽ�Ǉ>�*�=��>�!x=��D>���>�A6?+PC?A5K?��>ؘ=���>d]�>�5-�5zn�9�����<��?���?4{�>)�c<^�=����<�k����?O/?ǒ	?v�>S��pp��!�v�?�M1�����pa=(�5;��b:�=�*YɽE�:>
%�>l��>r��>���>T�g>`B�>���>���=���<�+�=	���η;q�-����=�p��(�=&���G<=�ʼ�fA�;�-��-�O�������D� 2�=���>o�>N�>��=�U���1>ʫ��۪L�|�=E���-�A�.;c���}�#�.��h5���>>�JV>���Y���K?��Z>A>���?	�u?�X >\�fiԾ�Ý�)9c�DS����=N>"~;�q�:��+_��	L��Aо0��>�Ë>�*�>���>g�/�T8�j!�=���l�4�e1�>�[����9��@��6m������K��.�j��<����7?����3�>�z?��J?*��?V8�>ㇽ�!Ͼ��.><�k���_=���̈�9����?�%!?��>����&z2��f̾
^���>��I�Z�O�����ϱ0�G;�x췾qǱ>7����о�3��[�������bB���q����>�pO?��?ўa�0M���1O�w��񻆽s$?e`g?�Y�>l+?EA?6ۡ�����4����=нn?6��?V2�??>�;�=��R=J ?i��>� �?*�?�9b?������>�un�=�~>6ߜ=hH�=)�i>��=`>�2?s�'?<�?A�8 �FxȾoz�����L�=�	�=�0�>��>$��><㯻�\����=iC�>��>l"�>F\>��>7��>�ں����+?�|">�&�>Ma5?{Ý>�	N=�k��/�=�C�W�T��s/��=���Ͻ!���=��=^�&:���>e�ʿ�8�?~�F>��D ?���˺V<I	>��}>�PA�ĺ�>Ǽ[>�>�>F@�>כ�>$	>M�X>��>�EӾ�{>��?c!�,C���R���Ѿc~z>����&�@���|��cAI��m��g��
j�t-��<=�4��<�G�?����k�I�)�P����?�Z�>u6?�،�����>���>�Ǎ>�J��ޏ���Ǎ��e�B�?��?�<c>n�>�W?ԛ?��1�c3��uZ���u�)A��e���`�e፿!�����
������_?3�x?>vA?݄�<�<z>���?��%��֏�*�>/�n&;�g@<=�-�>+����`��Ӿ�þ3�%KF>W�o?�#�?[?<WV��yt���)>=�:?�A1?�s?=�2?�;?%R�=�$?C`3>9�?>?2{4?��.?��
?j�1>���=��hr1=ea���ԋ��Qν��ͽF�ڼ��5=HRw=
a,;%��;v =p�<�	��~BռN}\;1y���a�<�%H=첢=M�=jƦ>D�\?���>�Z�>�f6?�ԽΓ3��1����)?�\\<��G��`�yϙ�L��{�=z�_?Ģ�?;p`?D�b>#�O��7��"*>u�>Q�'>�b>�>���i�4��ɂ=��>l�>���=���t�����������o=#4>�z�>c_P>! �>[4>:྘�x�iO�>q���߷��:�ǓI�NK'�����>v3?�3?*�p�X���3_���q�!m0?�{@?,f[?�b�?�X�=���ǳ7�LC�[0�n��>�@�=$D�癿����V0�=�;j�>��a�`��~dR>�����ھH�j�mL���侩q�=Cv��{=�i	�ъ׾Oǃ��;�=�:>D-���0�����㩿:�J?T�j= M���^��*��� >��>�D�>��;��Ő��<�ʖ��]��=��>��3>��0�.龗H�B�g��>h+?��u?�I�?~��V`��h8��<��ހ���=*�?�^F>��?r�5>�f�<�ƫ�1)�i~����O��>�v�>,���5V��d��<W߾� ��N�>�?U�=�	?�J?cd�>W�]?L#?	��>��X>��;ɚ��.13?�<y?�ռ^�������"�"�"��a�>'�J?�o���8+>���>�	#?�3?�M�?f?����;�뾢�B�KW�>��>��k��[��Uk�>�X?�N�>�*?�]�?��I>C�H���M�tو���>�8>�fL?Tb?�=?x��>4�>������=��>�`c?�Ӆ?B n?R�=�&?��1>��>e�=�ʜ>̱�>;�?ðM?�s?�yM?-��>NQ%<�K�������!��t<�8<J�9<{�=P.���$�,J�gd�<��;/\ּe��QS�H5��*�=v6�>\�s>�����1>j*ž�3��T!A>����uq��yq����:�q$�=���>6�?�|�>9K#��P�=XE�>���>���8(?��?S+?D$b;FSb�ɷھ�K�MͰ>fB?�j�=�l��w��#�u�g�g=��m?y^?<�V�x���=�d?�bX?\��j8�1��}-b�y߾��O?kp?��_�g�>��q?�sn?�k?g��̌c�����7Z�Gx�����="v�>��� �a�"'�>�T7?c�>9L>�>>�}߾�q}�P���~??b{�?��?B��?q>�e���ۿ����g ��_w_?���>��*�#?���ٵξB늾s�����'���������h񥾬�'��~���Խ'з=R�?S�p?�9q?@`?����ee�Ҳ`��&����U�B,��H��B��D���B��^n�M������`����.=�_�,�5��n�?y�Q?��O�v
�>�x��C;��I���HE�>|7־�}���7>��ོ�=��C���KT��M���8?.o0>���>0e.?c�S��N�%^:�ʒ(�X ��=�>��>.��>tR�>0�<���j۽���(>ɾ��D�@��>��U?��@?��{?�&�)X������'����a���\\f>^��=��>RӉ��e��C-���2���M�F�������(�+��>��c?M �Ȝ�>�!�?��E?K�:��~�������r����<��a>1 [?9p�>���>g�Ǿ=X3���>��z?r�>UU�>�h�R�7�����5@m��`�>Y�>pv?�m�>/G�̳S�k1��Q,��1�n>>8q?�^�������>��L?�佫��=/;�>��>2�����S��9>d��>e
>�}>�!������x����EH?��?&?�Z�2�L�>y�Q?ڳ?���=�Y�?��@>[i*�,cD>�>5ш?��+?:σ?�T�=�e�=`�&=��Ͻ�hL�$@�=c�=V5�= �=�Hٽv�"�sϖ�ZGT��q�='��>�P�?�D�Uy�ɯ���<�`u=* >�Eۿ\TN�ZӾ����I��I	��>���3=0��n^�������MR���>W��F�,�Q���N�8�t�[W��Y�?��?�5����i��畿��n�i��Gm�>��&�Z�>9y���: H�`�Ⱦ��t������4�gz_��rt�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >KC�<-����뾭����οB�����^?���>��/��p��>ޥ�>�X>�Hq>����螾�1�<��?6�-?��>Ďr�1�ɿc���w¤<���?0�@�V;?
q�y�� ��=S3�>e?�b>;0u�P����;�?û�?��z?�+w�BP��@ڽY�?�>�{8�������=�2>!�=( �d�p>�>!L��?���$��q]>��<>e�= ǰ��|���/�<�>�Ļ=����)Մ?,{\�tf�ϣ/�	U���U>C�T?�*�>�5�=��,?*7H�r}ϿQ�\��*a?]0�?ͦ�?��(?dܿ��ך>s�ܾs�M?�D6?��>1e&���t���=�DἏL��/��('V���=��>��>(�,���P�O��G�����=����ͿdB���2���	=�"�12�1�<.�%��	��bξq�N�z？)�=&zp>��L>�%�>��>�ˏ>�k?=s?���>cb>���5��5�ھ�I�<K���S��\>���3��,�S
��:���:��_#���!�h��T�-�7 E<|Q�Ĉ�b?�$e��2��"9?���=�*��7�8�(�y�)�Ⱦ>��^���~�*͕�vL(��n�I��?��7?x�y�B`�2o#�"w�=3�ͼL�V?�ܽ;#��Ƃ�aY�=-����;,��>� 1>�Lɾ�>�u�E��t>?e�?�л��g����=>)1~=�� =��?�?�08���>��X?�����e!�]c�>~�>���>kĺ>�B�=��ž�K�C8C?Z�]?��ٽ�ݘ��R>kl�������%<LI?؋��;"=�kȽ_|@;,E�H��>w�=�s��'W?ڝ�>z�)���-]��T�A==L�x?��?�,�>�{k?	�B?��<`j����S�� ��Vw=t�W?*i?�>����G	оM���(�5?Тe?P�N>Zbh����i�.�$U��#?��n?^?7x���t}�������o6?��v?�r^�`s������V��=�>�[�>���>��9�wk�>2�>?9#��G������Y4�Þ?��@���?��;<� �q��=�;?p\�>�O��>ƾ�z������̔q=�"�>����uev�����Q,�K�8?ڠ�?R��>ϓ�������=�����S�?���?�a����9;���Ol�/t��D-�=&�z="�JO��Vg꾀�:��=⾦�������C�����>0�@��/���>�tT����|Ϳ&�������圾o�C?d�>!Y^�S����l��lt��bS�51��dk�O��>�Ww="��������f���+���b�?�Ķ���S>��ýҾ�읾�M�=1�>���>%5>K������?����Doɿ�ꟿzݾ/L?�,�?��^?(L?6h���}|���?��g��2?y^�?�f? bV�Hz� ���j?J_��U`���4�5HE��U>�"3?zB�>I�-�ǭ|=�>��>�f>�#/�R�Ŀlٶ�����=��?���?�o����>u��?�s+?vi��7��Z[����*�U�+��<A?�2>(�����!�40=��Ғ�e�
?/~0?�x�F.���_?6�a�R�p���-��ƽҡ>l�0��/\������Ve������y���?�d�?5�?��n�"��%?��>{���_Ǿ�U�<j��>>�>�zN>��_��,v>m�� ;��z	>��?pr�?Or?M�����pF>z�}?f�>�F�?}H�=DY�>\��=�0�����D>E�=����>��>ЊJ?�,�>0 �=�9<��,��fG���Q�T3	�c�F��>��a?��M?X�x>�I��O�6�����ҽc/(����d7�%]�R��Ϣ4>_�<>�>�-���ɾ��?Lp�9�ؿ j��p'��54?.��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>;�>�I�>C�Խ����\�����7>1�B?Y��D��t�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�b��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?TQo���h�B>��?"������L��f?�
@u@a�^?*�7����:ϥ��7��A>�0=��`>�k{����=�B=,T�;[���Ay>q��>�ӛ>w�>���>���>o��>�&�� ��ᗿ�z��g�L���!������N��h�+��b�!��ꐾ�LK�i�f=���3��[���������=�`T?�8R?��p?���>0Gp��S#>X���=��<@����v=K��>�1?��I?�(?0Ȑ=Fj��@d����Ϫ��ރ�J�>��L>Ԟ�>��>���>k� ;Z�J>�4@>灀>cT�=@B=����j=�M>N�>+��>Ƽ>�g>��j=�_��)���/r�+�p���ż�?�x����n�+~�vM����!+�=��?��Y>h�y�P�ο)5��;�E?�6��F����S�K~�=i�0?��[?���=�5���?b��+>��P��u��=m0B��rZ����;�=ڤ�>�r�>M��;�5-�"H����|VQ�T�?t�?f���:=[c��Oz���`>�~>�>�@
�툤�0��,��	">�9M?4�?����@ʾk���.�0�>y��>��B��Xc>_�>�`߽�t=�ל���D�@�->�u>�L?PJ>R$>LK�>D:���J�H�>�#S>�(�=ɰ??��"? ���oq�V��7j<�omb>�6�>:@:>�">b-=��9�=�'�>��8>`�����v���0�N�Y>.�*�ôF�*�:�%wd=������=p��=dk��9�L�=p�~?�}���䈿��\Z��mD?w,?c �=�G<��"�y ���F����?/�@�m�?�~	���V�
�?@�?w	��^��=)x�>�ӫ>Qξ(�L�m�?lƽmŢ�;�	�,#��S�?K	�?��/�6ˋ�l�`9>�^%?��ӾPh�>{x��Z�������u�v�#=R��>�8H?�V����O�e>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9�~�'���?�޶?֯�?YhW>��?�	?��>���>jUI�c<��	����>�-
=�?�K�>��=���<Ԓ�歠�d҂�^?�����>�=޳�>�C��G\����>�A�����U�<�Bz>nh>�6>���=ߑ?a��>U��>��>���c=�@��WX`��zO?%�?�����f��7=�]�=�v0�+0?��D?�����+j�>kW[?tց?�m?W�>��yu��:��]����#-=}n>Һ�>���>Ln
:��v>���'&��Ù>�z�>�5=���<Y�snl��5�>�#?�V�>��>k�?s$?ԉ>@�>]<6�K�����K�>��>�վ>�v?N�?�?����^�4��+���N���WU���+>`As?n?�a�>�����L0>N�S���̽�n^?��x?\N�n�?��?��F?��?��}>�@��h��&=b��><&+?E��к_���=�|���4��>8&?Ӹ�>�X>�g���c�1=��1� 8���>|*?�;/?=���b�|��!�9#=Oy��2a<<ec<�E<��U>F�>��D����!�>7�I����=�۴<�Fλ�D�>`;=Y/�X_l=�<,?o�G�\ۃ�
�=H�r��wD���>	JL>��N�^?Rk=���{�����x��q	U�� �?���?Ck�?S��"�h��$=?�?�	?r"�>�J���}޾��ྖPw��}x�w��>���>O�l�W�*�������FF����Ž4�@��>�I�>=�&?h��>��_>&�>>0��x�&�����Ԟ����U���xx1�����	�c����R�?��*IھK�.�๖>�C\����>U�?f�r>��>���>�p8� �>�@,>�	>���>�6>�">dm>Ɍ�=��<l]R?��� �'�5��pg���B?-Zd?nD�>}�b�Ɗ������9?}�?�p�?��x>� h�~`+��N?n��>w��V�
?�4=1,�6s�<�����E��f��D��Փ�>D�ٽA�9���L���e��}
?Qh?���	z̾�qֽ�>��Ͱ=��?7?kM)��zS�Kt�tj`���C�\Ӽ�ݽ�W���9���h�����n������Z��	��<͟#?���?��"��� �9�Q�-y��@�*��=S� ?�&/>u�>3�>�����nE��RW�;}��َ�^�>�u�?��~>'lX?'UE?R�2?��6?��?֠�>:c⾍�?�r����>�1?T� ?$1T?o%)?��?=�$?��>@9�<2��D%��{ ?Dc�>R#?�A?[ ?&z7�p2)���>����㟾��̽*b2>,3>\�"�-b��� ���>�X?�z�7�8�*���Rk>H{7?�r�>���>Y���)��,8�<m�>}�
?�B�>� ��}r�#d��Y�>G��?����X=A�)>���=���Cnغ�G�=B0���ؐ=S>��Q};�� <�}�=3��=e�s���|���:g�;���<gu�>��?���>F�>�:��	� �����?�=<Y>^�R>�;>W/پ�z���$���g��Ey>Q{�?�z�?ޡf=���=��=�n��JH�����>����<ǘ?'H#?URT?锒?��=?�l#?ʶ>�-��J���\������ө?�R+?���>2
�-�ǾH}���/�,?]?�>Ɩ[��8��`-�T"Ⱦ�ڈ�w� >�V-���v�5���H�K-��i���[��?�?�v�?�}ü�+7�d����񗿄���#@>?��>̽�>wl�>fv(��)b�WL�F(>���>��N?܇�>�O?�{?�$[?X�T>	I3�Y���%���N�M�{>uNA??�?�*�?o�v?���>v�>�`���׾���P+)����+��8�.=��S>ג>���>p�>UO�=���Ӈ��>=�,�=�L}>�g�>+J�>�M�>�k>��=%�H?v��>��þ
'�����A�~��*��s?���?��)?�>�<���e�D�wm�K��>���?�%�?�|(?��Q�F��=�ȼ����X�t���>�k�>g�>+$v=��D=��!>���>^��>ȸ�(��e�:��2$���?��E?��=�/����d�Mz��[(<��E�=�<*��o���#z>�А��˰>2����:���)��G��˅���M���T���A,���?���-R��q�5>��=��=�߇>�;O�5<��=�A�=n�v���-=��=4m&��0����=�㙼�j�\!߾4Rt?{I?��0?�.?1&�>�+q>�a�����>:��l�>M,>�P���ľ��$�����jh����4��v>m��߰�5N�=&d��5�?>:P>w��=S��=��>�R����<=�N�NF<ٶ�=�l�=<r��>T�5>6H>S6w?����~����6Q�uq���:?xD�>���=��ƾ�@?��>>�3��w���`��#?���?(S�?��?$|i��a�>m�������(s�=����B2>K��=0�2�,��>� K>����J���-��1�?��@M�??{ዿl�Ͽ@i/>�)>y��<|![�ޗ<����}^p�˓9���0?1�6������u>P���W�þ�҇�ǲd>�>{cL�e�_��M�=쿽��W=�>�$�>M>�W�=�����0=�d�=ܱ>C,>��z<@��;���/�D=�g�=��S>1iy>�_�>�?>�1?�d?\'�>�gl�a�ξgɽ�Ǉ>�*�=��>�!x=��D>���>�A6?+PC?A5K?��>ؘ=���>d]�>�5-�5zn�9�����<��?���?4{�>)�c<^�=����<�k����?O/?ǒ	?v�>S��pp��!�v�?�M1�����pa=(�5;��b:�=�*YɽE�:>
%�>l��>r��>���>T�g>`B�>���>���=���<�+�=	���η;q�-����=�p��(�=&���G<=�ʼ�fA�;�-��-�O�������D� 2�=���>o�>N�>��=�U���1>ʫ��۪L�|�=E���-�A�.;c���}�#�.��h5���>>�JV>���Y���K?��Z>A>���?	�u?�X >\�fiԾ�Ý�)9c�DS����=N>"~;�q�:��+_��	L��Aо0��>�Ë>�*�>���>g�/�T8�j!�=���l�4�e1�>�[����9��@��6m������K��.�j��<����7?����3�>�z?��J?*��?V8�>ㇽ�!Ͼ��.><�k���_=���̈�9����?�%!?��>����&z2��f̾
^���>��I�Z�O�����ϱ0�G;�x췾qǱ>7����о�3��[�������bB���q����>�pO?��?ўa�0M���1O�w��񻆽s$?e`g?�Y�>l+?EA?6ۡ�����4����=нn?6��?V2�??>�;�=��R=J ?i��>� �?*�?�9b?������>�un�=�~>6ߜ=hH�=)�i>��=`>�2?s�'?<�?A�8 �FxȾoz�����L�=�	�=�0�>��>$��><㯻�\����=iC�>��>l"�>F\>��>7��>�ں����+?�|">�&�>Ma5?{Ý>�	N=�k��/�=�C�W�T��s/��=���Ͻ!���=��=^�&:���>e�ʿ�8�?~�F>��D ?���˺V<I	>��}>�PA�ĺ�>Ǽ[>�>�>F@�>כ�>$	>M�X>��>�EӾ�{>��?c!�,C���R���Ѿc~z>����&�@���|��cAI��m��g��
j�t-��<=�4��<�G�?����k�I�)�P����?�Z�>u6?�،�����>���>�Ǎ>�J��ޏ���Ǎ��e�B�?��?�<c>n�>�W?ԛ?��1�c3��uZ���u�)A��e���`�e፿!�����
������_?3�x?>vA?݄�<�<z>���?��%��֏�*�>/�n&;�g@<=�-�>+����`��Ӿ�þ3�%KF>W�o?�#�?[?<WV��yt���)>=�:?�A1?�s?=�2?�;?%R�=�$?C`3>9�?>?2{4?��.?��
?j�1>���=��hr1=ea���ԋ��Qν��ͽF�ڼ��5=HRw=
a,;%��;v =p�<�	��~BռN}\;1y���a�<�%H=첢=M�=jƦ>D�\?���>�Z�>�f6?�ԽΓ3��1����)?�\\<��G��`�yϙ�L��{�=z�_?Ģ�?;p`?D�b>#�O��7��"*>u�>Q�'>�b>�>���i�4��ɂ=��>l�>���=���t�����������o=#4>�z�>c_P>! �>[4>:྘�x�iO�>q���߷��:�ǓI�NK'�����>v3?�3?*�p�X���3_���q�!m0?�{@?,f[?�b�?�X�=���ǳ7�LC�[0�n��>�@�=$D�癿����V0�=�;j�>��a�rJ���I>�B�yQھ�h�3�R�_���=g��Pl==��2ݾ��ć>6\0>�1ʾ#�)�����mܩ��V?�,�=����/}��H˾��8>��>b��>B������8�˩ƾ3��=��>��|> 4m��0�֫S���9��>�Z=?��a?^��?\��a,w��W;��P� ܦ��V�rA?��>y�?�3+>ڗ߼;n��y�����h��5�U��>G��>U����X�d��*(�8��d�><u?$��=y�?Z�N?��>�nU?8�?8�>6�q>=��kО��(?��?I~u=���En��$8�SL:��E?"p-?�yx��Ջ>�?�o?��"?p{U?%�?�i�=�� �]�?���>���>�BY�[����r>��N?��>C:V?0��?h;>�'@�L���ي�P=�4>>D�7?³?�?�Q�>�p�>�W���`;ሜ>�g?ԅ?��r?�>�?
?��>\/�>��=��>lh�>��?�^Z?��m?m	O?SM�>5�<����������'�;9�Z���C�11�<+Z��v������wO=�I��{��_�s���|z������ݸ�>>1v>r����-7>fľ�ۇ���=>;й�l-��y����4���=���>�v?���>��&�kޙ=�4�>�P�>O�B�'?�,?�?�o�:��a���׾��G�i��>1A?H��=S�k�=���Ku�
�b=�6m?E'^?IY�������b?#]?�&�T<��*ž��e��s��O?�R
?��L��G�>�}?c�p?�o�>Ʉh�8{l�c���y�a�Q�i���=U��>^����e�*��>�77?>,�>}�h>P�=�r޾w]w��Y����?�n�?)��?!H�?��!>��m�<�KA���%���e^?���>�~����%?2�^���ʾ���󀌾C�*$���_���N֪��-�u{~��ѽG�=�?-n?�wr?�(_?�d��fb�x�a�*�~��eP�~��Y_�]�<�<H��A�&�m�RX������Ԍ����=P��@>�=��?��(?4�Q�ճ?늾�c޾�Uþ��2>�F���F_�?�N��O%�n���_��::pO��T����f�%?��>�I�>} ??gMj��@D���J�?1=���ľ��=f]�>V�>��>U��96�V�������@8$������>yAH?��8?]�h?��)��v���*�?���@���鹿>$ō>���>�/�<���_�e-��%R��n�I��՛���t>'c?�����c>�?�j&?A�3� ;��3�t�D�)�3��f�>�I?��p>(�>ȸT����V��>�<m?2I�>�J�>����3"�+}��_ܽq��>R�>2�>�u>�w#��[�����c��xi:��c�=�Ni?b䄾�j]��Ȁ>n=P?��<w.<rk�>o����T ����]�+�t
>b�
?à=�,B>Y���mJ���z�:����G/?��?V`���p8����>(.?��?�4�>�c�?ip>�ھn3���?E<?�G?tQ?�D�>G��=%n��W�Ͻ� ���9=ϸw>�bi>D-<=�N<o�:�����7z3�K$O=0%�=(��N�ֽ08�|���_��Kw:�]>Mп�]X��{˾Y��+�C�(��ř�rN=Qf��J�Ͻ1�ƾ7���Ҿ�&��N���7��Y˖�hxT�f��̬�?���?�~�(Ԑ��i��"�u�ls ��S�>)�5���p�;%¾t�*#~�s����}�Œ)�YJ�0��bЃ�Z�'?�����ǿ밡��:ܾA! ?B ?*�y?���"�o�8��� >C�<�&��)�뾎�����ο����R�^?���>���/��K��>���>��X>mIq>X���螾�A�<��?�-?Р�>.�r�8�ɿ(����Ǥ<���?�@6<@?b�$���Å=��>�M	?t�=>�6�������_+�>���?��?w[D=o�W���:�lDg?ޕ<��D���f�\�=��=55=
c��YI>�W�>�X#���=�ٯ׽�5>{�>���x	�]��V�<?�Z>��Խ!����ф?��\�_of�)X0�����;4>F�U?���>ژ=�-?@�F�WϿT[��`?38�?\�?��'?`f¾��>Ŕܾ@<M?�6?V��>�P'�`�s�2�=P��ļ�%C���W����=�s�>|�>�H+�WA��Q�������=�E��T˿����.��h�=�ӊ�������!���;�qL��?r��c��,r='z�=�!A>b�>���>&I�>�h?4�g?�G�>6�*>g�H�g���_<ž��@>����x<����xQ�w��|b̾p�Ҿ�6.�uJ��������d4��=�F�wq��3��d�r��3?��;?s6�=�~ľ$jM�J�弸Gݾ�d���$=���	��;��Il��&�?��<?����V���x�<6�__?D:��d����!�-=r�z�?3�>*�U<��Ӿ�zI�z+t�R�@?m� ?7�k��(�>]1;=O�{=��(?#?�ry�]�=f�
?%�s�l2���q�>xY|>E�>i�>���=x���]2�*�1?&�y?��d�r�����<����\���;�=@�>�)���Ľm�>I������>�Cd�e�i<|FW?�F�>�c*����쎾��8D=_wx?J�?fў>~j?��B?���<����;S��
�[<x=��W?[�h?>�_���]Ͼ� ���5?��d?�K>��h�LM�4�.���'?Pn?U!?�����}��󒿽���5?�v?Y^�Bz��!��U�ڑ�>ǆ�>e��>_�9�k�>5L>?�#�9�������,4��̞?��@&��?ͨ=<)~����=m3?�?�>Q_O�kEƾEL��f���Fo=���>Lp���/v���G,�gf8?Yw�?�U�>.���������=@���#��?���?����B�<5��6�j��q��	�<�A�=(��h����K;�:>ʾ\��i��5L��F�>��@�����>?<�j[㿬�Ͽ��H�žy�q��k?���>ﵽQ9���Aj�[Gr��J�B�D�ꋂ���>�� >�R�r��6��+A�%(B=9�?��=����̰��\��������m6>�D\>P�	?��=���H��=3�?-����T���Ѥ�a�~�N?�w�?br�?�+F?K*j�׻׾�f��6Ui�Z?=3�?>�|?�܃�֗�k�x�޹j?D��nC`�)v4�n>E�)U>.3?s4�>z�-��f|=Y>���>>t%/�k�Ŀ�ڶ��������?��?�����>Ǆ�?�t+?o��)���F��Q�*��8u��4A?�E2>�b���!��6=��ߒ�Z�
?m�0?$M�$.�t�_?	�a�J�p���-�f�ƽ�١>;�0��Z\�� ������Xe�����?y���?^�?��?3��� #��4%?6�>����x;Ǿ���<ƃ�>�,�>�0N>�F_�ʽu>���:�)i	>ˮ�?�{�?�j?W�������\>C�}?�B�>��?�-�=�-�>���= &��:Nk�FZ>���=��:�@e? N?M)�>���=8�-`.�S,F�S�Q�~���C��`�>� b?�YL?{_>�V����6�� ��0Խ%�4���ܼ�vA��}9��A۽j�2>ŉ;>A�>7C�/Ծ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�o	?D�NP��2a~�U���7����=V�7?�0��z>���>a�=�nv�i�����s�㸶>xB�?{{�?V��>®l?��o�
�B���1=<L�>�k?�s?o�����B>~�?�������K�# f?��
@?u@H�^?����n��S(ľ�pվ�>ce�=�>�g��A=�8���9��	b=j�&>��y>}s.>L|w>�6�>�Io>9�8>e1~����
��v-��CE3����_���z�����b�{��f��ה��������̽>�5��|��b.��_���m�=�U?�IR?8p?S��>|�d���>���� ��<R��bC�=���>S1?�_L?x�)?���=�(��_$d����	��Y��� ��>D�G>��>}��>���>wB�;�H>/U?>w�{>ͦ�=��(=��޻��=�PR>�\�>��> ��>H�>q/�*ױ��4��,�d�ju]��UZ=�K�?�Ӳ�.%A��0y�4J����4$@>)$]?Ũ��Q����޿[+ƿq�`?��޾ǘ&�6p� � >�y?�|�?	������� A>:J�>*�����AB>��S��0��:����z>PU�>
w�>��~=�9�-�N��l���(��p�>��?�;��Q/�=O�}�GKv��a�T��<"v�>��<�g�]����.������\��=h�J?��?�m5�등����|������>j�%>��s�p�T>q��>7�K������|��=6�>�,�>�|?��L>�J�=�i�>�L��n�'��^�>�J#>��=��2?6*-?lF�8�½͇����N�B(>� �>=7�>�v>(�s�1�=���>@cU>��	\�A����Ck�7cE>�����B�{}���=:���{��=��I=�ٽ�-��"�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾOh�>|x��Z�������u�s�#=R��>�8H?�V����O�e>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>:��?�gY?roi>�g۾;`Z����>ѻ@?�R?�>�9��'���?�޶?֯�?�.f>*��?�wH?�Z�>��U�[�B��Y������o$�>���<���>��>��ؽ�=��Ê�(~]�𯄿�g���7�>�����]�>w���bܽ��>��g�����+)�>�|�>�d�=C'�>m�R?J��>s��>y� >Q��3ɝ�����K?W��?��F,n���<}p�=��^��?�L4?�+[���Ͼo�>d�\?o��?�[?Wi�>���;���࿿�z���N�<��K>&0�>�.�>%���K,K>f�Ծ�TD�<R�>Fї>����3Jھ���̝���2�>Ec!?j��>�c�=;4?~.? v�>��>U_R������J�{Ԅ>�R�>n��>>n?h�?u�����!��O��8��ϸX��;_>�5~?�e!?��><Ú�ҟ��~<>��v����	8Y?�h?�B��?5q?i�D?�TN?��>�0ϼ����4v��:�`>Q�6?�����c���>�����q�?�?>?B�>��Y���^>(�A>�GM��'־�?�8?�?��ؾ�vu��5/���<?D��= =��Z�I�Y�վ�=�z>?m�����<�,�>=R7��6�&�P�A�V�m�/�0�>.g�N���hB�=ر+?(f�T?~����=�(p��v@����>4�G>�\ȾO[?E�+�@�w��������[�+�?}?�?X�?X�� <j��>?��?�?b^�>re��C�پh�	w����u�ѯ��>���>u�ݼ���n1���3��ځ�V�ҽ4E����>���>V�?ӎ�>ـ�>q0�>h`b�pZ"� jD�_d����d��V۾��0��,,�ä�_����)�Fz&�����⒉��#h>�O�z�>��??Dk>�w>4�>Ԩ��f�=�0���>�@;>
�=1�=#^>f׍��'��KR?����n�'���±��[2B?[pd?d/�>ki�����{�?D��?-s�?�=v>�}h��,+��m?l=�>��p
?rZ:=DC�]%�<RT����-���ƨ�>�D׽!:��M��kf��j
?[/?6����̾�C׽��X9<��?�~:?��@�%)�>�h��K�/2���5�q���ת��2.;�����˕��y����}�̓���=�@?�Ɉ?1��>��O]Ͼ�#c�n��=�{?(`o>v��>���>�#꾝�
��^����p�׾Z��>Jd�?J�G>$Tt? X?��C?�oQ?�>��>����P�>û=�?���>Y?.U?4A?���>qRA?��>����������?M�>dX!?���>s'�>B�(�����W�=�}&��n����׽v�>lY>��>{��ε<GJ�>�k?����8�h1��p�k>�7?X��>���>	����u�����<#��>��
?>��>J����r�?I�w��>Ò�?�w�a=��)>��=)C���5����=k�üB��=R���%;�\�$<(�=��=bu{��>��0/�:K�m;��<]d�>��?�Ɋ>��>3���j ����蔯=װW>��R>�>N�ؾ�x��-#����g��x>U��?�n�?4�f=�:�=B��=3��s8�����ꏽ��K�<�E?�%#?�*T?u��?_�=?ً#?V�>s��A���?���㢾z}?�5.?zor>+	���Ͼ����=&��?���>�P�BE��vf4�_7;�{"����=ս(��dq�
)���CJ���@��x�U.\�4q�?�W�?��;�4��B��0��0���@�6?L��>��>��>�< ��Ge��C���@>�?�zU?��>)�^?�� ?GR?�ǧ>��C����Ջ���h�>I˽>�z#?�?M%�?�2?>ؔ>�XB>4
����۾�,�<���e�E����'�=;��=�J>���>�*�>��\���8�@�4�$��''�[Ix>���>8��>_�>�^�=���W?��>�T��79���<�Ui���Ş>��?!�?F�S>󮡾�$�AW����??�9�?2�?w�1?�U��?�=��w�������=�(?�� ?�ƌ>����bI<��>��t>���>Ӿ�f1�n7.�U�M�)?T\?b�T>=P���o������N�Z�E>�~�h�x�ހG>�5����O���H�_�A�����]����O�h���Q]c=����?����ì�?3`>�p���������=$�d��Q������?��
��y�P�}_�=�B���B=<���0�*�e��=��˾�g}?	,I?�+?׃C?*�y>�|>��2��s�>����?�U>��O�������;��������O�ؾo�׾ed��柾N�>��I��>G�3>���=�d�<��=�,s=��=����:=U��=A�=N٫=��=E�>_8>�6w?>�������4Q��W�Ѷ:?9�>|�=�ƾ @?+�>>�2�������b��-?~��?�T�?^�?�si�d�>,���⎽�q�=ȷ��=2>���=��2����>��J>u���J������`4�?�@ �??�ዿ��Ͽ�`/>k��=N� >٢G�VB1��>�څ���z�g�'?&�2��_����b>:��=����ǿ�i�=#Q4>���=�s��m�X�W��=�D��:G�<D{�=?{�>OO>�1�=�����$>���E�
>�E>B��i4�=;ء�=��=�P[>zm&>��>|?r�1?��h?�5�>a�v��5ϾϾ�>Ն>�$�={u�>W�=�dF>���>X�1?�:B?L?m|�>���=6��>���>��*��"m������M�=$Ç?Œ�?,��>,�><68�;���Z>��dֽ��?�8/?Ģ?"��>���+�Ήc(�p28��f_�����ah<�\��2��+@w�����=u�LY>k��>>�>﷩>�k�>�c>��Q>���>~n�=�=y�?='ܺ���\��O]�:��=s�ƽ���=�i?�!O�O�n��o˻�DG<F��;}��<k�&�70�;�$>��>�S�>�?IU	�%C1�L`A>X���J�K��@>h&F����Z�T�mZp��n&�W���5�>��w>@�� ��$�?о�>հH>���?��a?ڃ#>���f徙�����󓂾��=s�$>�v4��x&�2��|,�^ľ``�>���>`�>�Iy>�5-��9��v}=���c�1��8�>{���\���-���mp����#֝�k�d����;w�=?����� >&�}?$�K?f�?�W�>�ⲽ��ξ+%>�i���Z=o�ć�ۍz��~?��!?-�>4 ޾�Z@�U��Ử���>a��g�*��T��c9����=����>�¾a���8��}��n2��"�I�dM�?�>#�2?5��?v���Zil���7�g� ���(5�>\�e?M��>�o�>���>ظý]�̾�>���>E�u?tU�?�Լ?�R�������>�D9?�?i��?���?��[?M�� �k>�?>��>�=*�>�)�>k�>��=��0?j?&2?|�s����Y󚾝��j��ۼ&�=�Y�>�>�k�>����8�=YI->`Z^>s$�>���>���=<'�>��>S��&"?��>N��>�83?L��>o��=�ʽz1�<���[��%�e�Xx$��5�>��8�3=kM�=�&���>3����u�?-�f>պ�?����M�����e>Sg�=,1�����>�~=�hJ>���>]1�>�\�=�t�>��z>�Ծ�>����*!�ԊB��VR�	oѾ��{>�]���'�R_�s����JJ������5�R�i��
��ä<���<I�?b��N�k��C)�t���;P?Z��>��5?�V��-���>�\�>���>2�����������%�?���?I:c>��>1�W?�?~�1��3��uZ���u�N(A��e�W�`�i፿�����
������_? �x?*yA?�M�<Z:z> ��?��%�	ӏ�F)�>�/��&;�*@<=4,�>�*��v�`��ӾǺþ{7�_IF>��o?%�?�Y?�SV��b���I@>ivG?�*?h$~?�V5?N�;?����E?flU>ݜ?;�?S�2?�4?ܕ?c�H>1Z>�c=$��=nƟ�X���D�ƽ���5���/2=��b=��,=���<�L=C�����6��~��G���$@���j#<� �<���=�>끟>=`[?f�>sǂ>�7?�l#��8�������-?��2=����?n��S��8-�0�>�8i?r7�?�[?v�^>��C�1�I�U'>���>n�&>�b>M[�> `���:�߽7=
�>��>�w�=a'��z��L��K����<u�">�?%�N>��b��Ia>�졾o� �	�j>i�=�
8��s��^�&�b�U�`����>�K?p�>o9E>R�¾�b���i���2?�Mj?a5}?�J?�l�=Gaݾ�Y<�͈h�<�b��?��N>d���~���H����P��g>���>�OI�D�����=�������=3�����q��>*�8���3<E�1��r޾���� >7�u>�"��`)����������KU?�� =�ľw�������<��=�M�>�<ʽ��R�����?���p=�8�>p�>��1�aԳ���h�^�-��S�>D�D?3�^?D��?W@��Ɂr�yAD��p ��=���ϼ\?79�>�&?��<>��=椰�P���b��E���>c��>�m�_$I�[㜾�h���C$�t�>R?�>�>?:#O?��	?�b_?4^)?+�?G�>
����x���.?Yrx?ވ=�wս��5�)�4���4��� ?��5?������T>�~?�"?g�*?a#]?HE ?۽�= ��ъN��>���>K`�#ܩ�+8z>�=A?&�>�J?���?T�Q>�Q�.ִ��W��l��=�V)>7z7?�?�q�>�.�>=�>gP���~�=;)�>��d?�/o?7�w?36�=k��>ĚS>2L?�E >!�>հ�>'�?�xP?@wv???}w?�t�DG��l �{;#A�������%ϼz��<o;Va��S<$;<���Y#�A<+��9`=������ ��<!]�>��s>s镾�1>O�ľ�3��;�@>棼�Q��>Ί�Yn:�n�=I��>��?���>�V#���=䪼>Z1�>���S-(?P�?�?%;@�b���ھ��K�s�>vB?}��=��l�|y��&�u�h�g=��m?c�^?t�W�c���5j?} C?_��ا,�]-���Yv�ھE�H?�?3����n�>#�u?l�j?�K?��n�H�����d�+��ٷ���>���>�!�2Wk��I�>7K ?�?|�>�y�>���\(��z!��{��>���?DN�?���?0��=��o�����}���ݑ���^?�v�>ϧ���"?w����ξ,!���8���$��g��5����B��(���[F"��p���&ؽ�=w�?S�q?�&q?o�_?����X�b��H]�/����U�q�����E��+D���C��o�J�����?���-gG=
���e,��͹?+*O?�=��>�`�������a�z>���Z�=i>�6��7�2J�=����}���6�"*?��>�|�>�M?�82�G�<�\,Z��+G�
����>��>|D�>�'�>���T�� n�sʾ�a���)��>�NL?��>?,aa?}�(�f�3�<���v��!gJ=�С�$�>Fu�>�!�>�р��E��v����(���_���[a�$U-��>'wO?�a�=��>͔�?��8?��I�K�W������%�4��:�>q�K?��>0��><:*�or)����>NHm?ؿ�>[;�>񑅾��%�����$��O�>MK�>B��>���>��ڽ�I\�CZ��,ㆿsw7�;�=�b?�vy�A��{��>(eU?��G���<�N�>��������b۾8�>���2>GN�>s�=f�X>0-��5�?�z� �z�$N?��>(�(��9�G�>|%?+� ?�i�=�T�?pS�<BK�d�Q>0U�>zI�?.5"?��y?F�p>58u=�ED�Q�qB�����<uq>�T�>��G>�`��ˁ�*!��B��A>�ȏ>�w��&�<�����F��k=,,>�T�>¨׿��C�Qs߾&3�h0�����+d����=�ʾK(J;jl̾"v �&��9�߽I8�<�����H��6B�t����?��?֖m=�������X������:"?�n��h%�R����'�L�3�q񾾌q�����/w�d���|�w}(?�e���ǿ����z'�RI!?m"?Lx?O��� �fX5�k>��<!�̼��Ŗ��ߪο�֝� r^?�r�>��쾀܋����>b�q>��N>�Gu>�X��`՛��t<�^ ?�U+?�?��z�,�ɿ-������<���?U�@Is4?Z��������t�>|d?�?ifK=�40�evA��v���-&?>��?�|d?�䜼RG�C�����?�Z>��"�.�:�o�b>�ɕ>D�?>�����]}>�Я>�R��Ӹe��Z�< �>��7��m>ʣ=�Wk����i��>�E#=�,$���?�t`�lGn�X;��b~���I>OY?Ő�>È�<i,?P�,��?տdfc��sP?}��?�6�?T�?��־�>|MӾ+D?�F5?�ܖ>��4���q�Z�>��¼^������jb�R�.�W��>�><���W���p0�	�<m:�=4��_&翐(D��M��G�=�ҽ=m*&��e2�L�'�B��>�.����U���
>���>L	��}�>ɉ�>��>��F?J�[?1�`>�pt<���]5}��XJ��"=,Mо����L��;�n�e$����%t~��0���ؾ$>ھw�¾2�1�9ҭ<�=�g����'��.u�&�N�Y�H?p==/��1N�2�<��ž�|�� d*=~�Խ�ھ+�?���x���?Q�/?�G��G;�d"�K��'�ֽ��N??��3��9��G�=��<���>��3=�7���=6� �T���8?��?�{�ܗ����>h6;��n��4P'?��?;����Y>(cD?Rv���y<��>;�b>q{�>#��>Q�>[i��!����/?��a?�o����9�:>Jl�8��-N�=P�>��.�Z�,��m#<-�Ä���$�>�����?w�}(W?���>y�)���a�����MV==%�x?��?�-�>[{k?��B?�ۤ<h��v�S���ew=��W?�)i?�>y���=	о����ڿ5?��e?Y�N>�bh������.�=U�k$?�n?\_?Uz���v}�^��C���n6?��v?s^�xs�����L�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��V��=�;?l\�> �O��>ƾ�z������1�q=�"�>���ev����R,�f�8?ݠ�?���>�������i">9�|��D�?�Y�?G)��k����,��l�NI˾�*�=b��=�>>��j���GW��#��~����=�֊��_�>��@���qס>`�Ӽ���8�̿����	��[_���g%?{܋>�=�fm��p�!^e�P�O���@���Ǿ�{�>��>� ��VQ���(w��9��<� �>�������>�Q�LP��l6��L�d<�d�>�>�}>
j���{�����?>J�D3Ϳx���a�W�R?L�?פ�?h\"?��k@m��x��ˍ�v�L?�V}?��Z?�g�PqB��|ѽ:>j?�R���eX�x�,�#R�3�i>	6?��>>�*����=�(�=���>E�<>��?���ÿ鄳��
�p~�?���?������?H;�?��<?�	�y���T�ϾI�<�3�p;ҲG?xr">ኾ�q*���=��㘾�M?�$&?н�{�n�_?��a�Q�p���-���ƽsۡ>_�0�Ze\�xD������Xe����]@y����?7^�?l�??��� #�
6%?��>A��� 9Ǿ��<ڀ�>�(�>1*N>�I_���u>_��:��h	>h��?�~�?&j?ϕ������U>��}?'�>��?T��=�[�>qb�=����(/��=#>�R�=�@?��??�M?�U�>��=�9�(/�@WF�EBR�� �)�C�c�>��a?�L?/b>�����2�Y� ��ͽL1�k��dB@��,���߽,5>��=>�>�D�9 Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?qQo���i�B>��?"������L��f?�
@u@a�^?*e޿�=���ھ�Y���q.>��=� +=��ǽ��=��i>_�=r����>s��>,I'>0�8=e��>�x]>���>����E�'�-���v���LG]�@ؾ�Y��<�8�;��A0 �H2���~��nO�<�F��4��"Ꞿ7*���`����=��O?�U?�?r?���>&v��>����)<c�!�d�m=��>�/?"�D?q'$?��=H#����b��c������+/��Zz�>řQ>X��>f�>�e�>*���a.>�H>��o>�~�=i�-=㦱�W1(<V�O>�}�>�?�>匵>� �>󇜽���Ks�����X���<��3S�?���zv���{n�aJ��A�徂[L�2)?C��<$Ӊ�� ׿/���O�M?����n7�=f�_S'>�)�?(�}?,6ѽ����_�>5!�>!9 �����ݗ=i�>�{=�B��E�=�-?>A=)�O>t�K�H��S�C��1]���W?�)��b�*�~��K/���-�xN�>i�>o����*��:��t=����8��Q��{,?��>x�=�kD�،+��s��j�{>�S#=���=�D>��2=ٔ>��C½�b��h�<��L>�У>��?�>w�j>R*�>�����'�d�>�H�=�Y�=�5?C�?�u"��۶�a���k��n�y>��>�>>#��=��/��J�=Ĩ�>YQn>���;�^ ��8�����`�f>��<��w���z�Py�=L�ؽ���<���=ʑܽ�;!��8�=�~?���)䈿���d���lD?P+?M �=?�F<��"�F ���H��@�?q�@m�?��	�ݢV�?�?�@�?%��X��=}�>׫>�ξ�L�ٱ?��Ž8Ǣ�Ȕ	�)#�hS�?��?��/�Vʋ�<l��6>�^%?�ӾQh�>|x��Z�������u�u�#=P��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?g�m��A���@����>:��?�gY?voi>�g۾A`Z����>ѻ@?�R?�>�9�~�'���?�޶?կ�??��>?��?k�-?��>ȶ=�gW���6
���g�>�������>H1X>�%z�i�O��=���7�<&N����MZ�<�e=|�>x�U��!���>ν��;����a�>���=�7�=삻=�?O[>�Ġ>4�$=RE��T��"�	��N?�?�k��j�'�=$�=��I�?�??�9?�����a��>��[?o��?�(]?�٤>�=�`���KG��������V<�>O(�>h��>�)�(�[>�{߾�y@�ۑ�>a�}>�8ϼv��	1y�����^C�>ic!?���>���=��'?X?v+�>JN�>,��	��@W�j�x>?��>�?aO?#?��1���1��͚�Ԕ��DD�V>��x?�D?p�>~,��9��������7���U���v�?ԡb?�:����?e�m?�
?��f?���>c��d(�Ѧ6>��<��>?l ���7z���S�ܓ.���.?�X?�f�>��	��	-=	[+>��"�dW8�iW�>e}?��J?��1���|�q�h�G��< c<���:��a+a=�>��>;�^��t/=R�>�&>(��o�F�^�<L�w�h>�Z�<��<bp�=+=,?��G�Vۃ�'�==�r�xD��>�IL>v��{�^?Wk=���{�����x��^	U�� �?��?Yk�?6��C�h��$=? �?j	?"�>�J���}޾{��	Qw��}x�2w�y�><��>r�l���O�������nF����ŽD����?yX�>3d?�}>#	�>���>!������7���֨�9~�X�!�?���(�^�癆�	Q���7<e�ݾ.����ð>5<Й�>k�>v��>�x�>�?�����#>�U>=C�>@�>�J�=pc=���>5 �>��=�VR?����A�'���"����B?h_d?�G�>�9f�5���y��w?h��?Po�?@�v>�:h��++�Jd?<��>����c
?!�7=���냋<�8��?����> ����>�;ٽ�!:���L�'f��i
?C;?"Ǎ���̾�;׽[8���3=	��?ð5?V�"���H��p�؁Y�Z�O�rL;P���&���r���t�������}�� z�'�;��=s�&?���?	�����v��|�f��B�$�k>eP�>3>���>eFB>�^ �!j!��GT��H)������>�'y?�!>\q�?�H?��P?��W?��?~$?���㵪>`�=&��>Bi�>4�C?Oh?ʹ&?�ݹ>��|?�V	?g���}�b��9?�V�>נ9?��>ܛ?�T7�`[2=��߼��n���6��b �0y轒=>E_ >�ͽ�R=J��>zW?���8�G���Hk>|7?rz�>���>@��Y0���'�<�>e�
?�@�>� ��yr�Xa�+V�>]��?#��"w=D�)>���=\���H2ѺxS�=v���2�=Q(��݋;�K�<I��=y��=��s�&
~��x�:���;���<�|�>��?�>*��>�3��k� ����=��X>JS>0�>�پ�h��z&��h��Sy>o�?;d�?"Ig=9$�=���=l���I5�����"�����<,�?�>#?�KT?���?m�=? d#?��>�#��H��&Y��`�յ?w�:?�='n����EⱿ0��p;?�-�> �W����4j��[8�&$�<����p�0�$6[�%���q�3���=S��'�6<x��?��?^�f��w6�X^�\���Ց`��^>?]i?=�f�>��.?�GI��={�;3�gE>6�8?�??�^�>SQ?a>v?�w[?p�S>��.����95��zg�]�>��>?�?{?
J�?��p?^�>�=�=�s�dG;ja���E�6�ܽj%��~\=TH7><�>`
�>�j�>l��=�T��%�۽io4��X�=�>��>�u�>j��>֏l>��<��H?,�>�$þ3)��̡�]����$�$�s?��?T�)?���<�c���D�L���+�>���?��?�A(?��Y���=�2ۼ�����w�
��>hҽ>5�>�8x=�y6=\�>���>���>��0@�V�9�p�N���?�E?���=�;���.f����~ž��M�O�Ǿ�����F(=�U$=�鴾�F�D�ؾj��p��������&Ⱦub��*闾�-?^h�;�.�=���=��.<�h�c)�<��=2s=���<��
��<�v�=��:���~�}�<��<�?�={Ȥ<�.Ⱦ�e}?��G?*?��@?~�q>S%>�W�5��>�ݢ�v�?3E>	��Yڿ�v O��u�����-�̾�AϾ��a��=��M�>#�O���>�4>q��=o'�<���=4BN=%?y=���<��=]��=.�=t�=$�=��>�v>�6w?X�������4Q��[罩�:?9�>k|�=��ƾ2@?��>>�2������zb�.?w��?�T�?��?Vti��d�>H���㎽�p�=����I?2>0��=��2�D��>c�J>[���J��5���k4�?��@��??�ዿ��Ͽb/>��!><� >�K��Y4�@6h��%����o���%?�=���ξ�<n>��=��`���'�h=?�$>G�=�<�XAa���=�$��_Ic=��==�>��L>s��=*����=�)#=�O�=g{T>GA��&!�l<��3=	�=R%w>��=>�Z�>N2?�e0?�kd?��>�Xl���ξ ���?ۋ>���=���>jr�=s�C>;{�>��7?_#D?b!L? �>���=C]�>TF�>V,���m�J��m�����<qc�?4��?v�>�E<�IA��f��=�
xý��?�1?Xm?8�>;{�5�ῃg'�G-�����`7�;Z�=f%t�;�^�?*�"!�D��{Z�=С�>�F�>��>�5z>#=>�%R>��>G�
>~�<�Ԁ=ۭ�:~ɼ<E�n�m��=lݼ��<�gż���]��H��|W�(�q<� �;T�c<@�:��=���>�|>A��>x=���5[3>�k��#�K�7>gC����G�P�k�Uɂ�3�.��b�!.	>�<>� �������?N�X>��'>c��?<Zi?��=>4Q���Ӿ����;9E��D���f=�A>v� ��..�Y�G���I��ݾk��>��I>�i�>�*�>��E�;���/�=$j��I-�3k?���P���^.�i���߃��w����&{����<_h>?�*�����>��n?�KK?���?���>�;�oO�����=��4��s=�������j�<YP?)].?H�>g5�>\�EB̾,����>0*I�	�O����ű0�3D�
η�ܓ�>������о�3��g��������B�PIr���>ѶO?R�?�7b�2X��}UO�:��4��o?�|g?d�>FH?�A?�$��Iv�i��e��=��n?��?s=�?�>�"��_y">�)?��>��?oq�?9��?E�����>��=�P�>�=Y�>��><�>���;�F?\.?��?j�����)\����'.��R˽���=��f>?�=>-�s>�N�=ډ=��>��m>��>�K�>Tz�=(�&=(l�>�3�����NP5?�GR>��@>��0?��>��=�i=�D\�B�ǽ�@�#Gн#����E1�aQ=�=�>�G�=�*�>n�ÿn��?*�k>���.?)N�U����|>_�>����w?w]�=/e�>�&�>��>� >�rS>��>=�ӾS>4]���!�8'C��R��eҾQ�|>�\���+'���������M�lx����� �i��'���=��R�<��?FW��D'k���)�����
�?i��>г5?�/���Z���>A��>���>2���A`��������H�?A��?{Cc>U�>M�W?D�?�1�)3�vpZ���u�+(A���d�o�`��ݍ������
�[G��S�_?�x?�pA?�:�<s1z>&��? �%��ˏ��,�>�/��";�V<=,�>!��d�`�O�Ӿ4�þ48��0F>�o?�"�?W?U:V�������>��0?N� ?�p�?�7?�6[?dNc��O(?��g><�'?��?�@??�?��? ԭ>2/�>P9>!�>��������wC��;�	�<X�r��8i=�!�1�<�E�:��W����=A�h<Ա���"���'�8[��}=>l9e>ђ�>��[?o��>l��>��6?Z]���6�;~��e-?�C=�C��ƶ���m�����f��=G�i?���? X? Ke>��?�i�B��z>6��>��'>/�Y>3�>����7@�UԌ=_	>u@>c�=�&U��^�������c��<�%>;v?��> �ٽ��,>4�l���K�e17>���1����K�=�����������>�ME?��?�i>�fҾ�~��d���"?K�J?
�Z?��m?�Õ=�Oپ��1��\r��ڵ�!^�>D����y���g�����t�Z�#�4>)�>�x��⺖��D>3����澗�l��%C���ھ�R=���jq=k�z��Á����=3*>���s�����,
��$�F?D}Q=X���RK�Gɾ��>U*�>��>Ѥ+��f�nA�]���I�=�
�>5>E��*���:�L�2;���S�>�2D?+eZ?���?�0����u�ĘG�4���3ę���E�?"��>"�?q�->V�V=�r������`�T�A���>q6�>��uJ���������j���{>`?�>3)?�~N?�y
?�(Y?�&?��?�j�>�@ཱི϶��5/?�Kz?�6�<G۽@�M�� 4�%�*�;h ?��<?ISn��N$>{�?t?�i0?��b?�#?�t�=���t4�[�>�\�>ߝV�,n���!�>#%[?��>y J?2��?��>cB�����ov���>�9>�.H?�%?IT?�~�>9p�>!���\�&=��>�s?��~?ܝt?mg�=��>^�^>�?I�>ܧ�>_D�>k?BCB?)\?�,X?�o?G��<��2�� �SF�!q�<Eu<8oS=�"=A��R7��7rU<<��=T�~�ս���(<|�ټ�q"�,r���/�>�u>ۤ����5>�ž�9���A>؊Ҽ�����_��@J7�i��=a�|>g7?���> �%����=_κ>��>M��&)?��?�?���;ea��ؾ��K��>�OA?�m�=Z]l�L[���t���}=��m?�!]?Z�U�N��	d?�Z?�/���9�a{ž�m�'���P?A�?�\���>G�x?�wk?j�?�"K���j�n���`��
n�L�=���>+���d���>��6?���>�i>��>��پ��=����?�?�(�?���?a�>IBr�Maܿ���梑��
]?�2�>㰾�� ?Xѫ:D�Ҿ�ώ��m��H���߭�k�ʩ��������-����������=��?Wr?��q?OT`?�E����a��o_�C����S��f�����@�I�G���@���k�%�#�{m��I;�<�ri�*�F�eλ?�D?^���B?!ڶ����Լ�!V�>�a���o���S��������=Ŷּ��0���W��(���9?�'w>��>�8?l�k�g�R�;\�u�<�#W��ݺ���>",�>7�?�ۼDe����9^��t��Jмǳy>b�R?�=J?��o?�L��:�o��3޾��u��#Y���V>��4�5�>w,��ȱ�������_��/`�)�B�6 z�9�&�㼻>WZO?C�<��>��?*�6?Γ]���T�P��2���Y��>��>`�/?��=���>v���6����>��`?�?���>9o��
�!�,,v��Ǎ�O0�>䗭>���>v�=�E��O��j��o9���w=�Y�&=�7b?4C|���b���>?�L?�R�����<��>����"���վK"j�8��=.M�>�����\*>��Ծ8���k|�8�����a?�'�>FF�L�C�?�>�BI?�}?��>6 �?��6>bB�������?���?��g?�P^?��>����[�.�z��吼���5=�J>��=�ڰ<?�f�R��C�e��AI��
>�P">�W�=Y=��>=�k��N>�[=�> \޿��O�o�ǾO������L�����uX������ƾ����B�e����-CR�j�M�_�M��<n����!�?A��?���������g���\q�,X�r�>��m�-z������XT"������޾C����*�S*A�v	U�*�a��'?`Ñ���ǿ0����Dܾ�  ?G ?��y?.�"�ɒ8�J� >
W�<
Y�����;���l�οF���S�^?���>������>��>n�X>�Jq>w��Nߞ�Za�<��?i�-??��>)�r��ɿ����5=�<���?��@�.?#Ϯ�RA���>���>�0?�u�=`�����)��o
�\e?7�?N:h?�#<A�k�6�2�@]w?[$>�vD�P�3��{�>?�W>R�=95���X>�n�>��������K��e�>?�Y>dC=�H����5��⼋�g>���y`���Ԅ?\�pf�5�/�_S��o>d�T?�!�>| �=e�,?P+H��~Ͽ��\��'a?�(�?U��?��(?�쿾0��> �ܾŃM?#C6?���><s&�+�t����=��ִ����㾿-V����=��>Eh>�,�E��Z�O����w�=�;��sƿ�Z"�Y�� ��<؛Y��b����Ͻb9��f�K��F���_j�'�B!j=2��=�<Q>5��>v�\>��P>��X?�bj?��>�V>���������˾�}ແ���7X������� �ɟ�n�쾦پ����
�J�cuʾv�%��Y�ON��ו�j1��a�ĈG�~�w?e6=V���X6�n��=�3;���(ኽ�s���½`�%���x����?W�?5����C9�4�̾z%z>���<X�?����)�)Rg���=|4���wW�r/�>+��=G����?�2�<�K�2?�?:ƾO��c�.>iv�|=�*?�?�;��>��#?K�����w>j->��>:�>��>p���]�Ž�7?t�V?$/�;��f�>�ܺ��L����<W�
>�3�Q!0�Q�H>K%�<���?N������`/=�$W?���>f�)���d��J��!==��x?ɍ?��>1vk?B�B?�M�<q����S�����w=l�W?�i?9�>t���о������5?F�e?��N>5nh�U��/�.��Q�?��n?Y?�朼�q}������Uh6?q�v?Br^��r��<����V��:�>�Y�>3��>9�9��h�>�>?4#�mE��h����X4����?�@���?��;<���0��=37?AZ�>��O�o4ƾ6k��r���<�q= �>���cv�����`,�]�8?���?L��>���� ��
�!>Pԡ��q�?>��?����u_��M9��{e�_/����w=K�<	�=Č�<����;������(�Ryz���U��[�>�a@Qd��{*p>Et��|����}Xa�sd��3¾��?i�S>�2>A��U�z���G�Ywy�� �>�����>���=�RݽI+f�|�n�"D=�޳<D9�>��C=���=Z3h��M��7�ݾ��>u��>*4�>�~�=O�ν[|��M�?�ľN�ǿ�~���ƾ�o??Z�?8c�?ٻ^?�v�����0q>�ޝD>0T?ca�??n�?���{M��P�����j?e���R`���4�LE�&U>�%3?�=�>��-���|=�>Q��>Zg>8$/�2�Ŀ�׶�������?\��?�p꾴��>���?�w+?Og�#7��	e��=�*�'�(�V8A?Z2>�}��[�!�.=��ђ���
?�~0?�s�j.�E~`?1}_�QSp���,���Ƚ�X�>Z'�kR�F q���'���g�k3��Dcu�ح?bU�?{��?1�%�x�#���#?.$�>�}��y�Ⱦݍ�<>s�>v�Y>��_�~�>u����=���>G�?�J�?U?Y狿���Qt>�~??�>k�?���=���>���=�벾�Ƚ���>f��=m�d�I�?��N?te�>�K�=8�H�G-�;�E��WO����wWC�ڪ�>g�_?�H?��b>�㸽�;���3#���½:��k����7�����L�:z9>^�<>�b>��J��hξ>�?�n�ؿj��Z'�54?ƾ�>��?����t�!��|=_?#w�>�5��*��U$���0�˚�?G�?�?��׾d�̼">��>vI�>��Խ����������7>;�B?���C����o�S�>��?��@�Ӯ?�i�j	?f �qP���b~�p���7�}��=F�7?�0���z>��>,%�=�iv�|�����s����> B�?{�?o��>Ѯl?�}o�J�B���1=nL�>t�k?�s?��q���ƲB>h�? �������O��f?O�
@�s@T�^?7�}�޿RM���'�Җƾ��#>#�8��B=��x���d=-�=l9��8�=ح�Ԯ�>�Z�����>e
:>�ӆ>ò>���8f#�4@}����P�-��JI�� J�$���|��)&�,.:��wx�-��~�	��I�~�kɊ��6��r��{��=��U?�R?�p?u� ?�<x���>ȭ��1=��#����=c1�>a2?P�L?X�*?e�=.�����d�D]��F��;Ç���>ZcI>A��>FG�>1&�>��H9��I>�E?>=�>}� >E6'=�&�K�=��N>�I�>���>r}�>�[>�<�=�޷�����<�_��?H��Ͻ��?3̤�P�N�����叾�о�2�Ҽ1D.?ت�=U���n�Ŀ!��ڗH?A���Ly�\��b[>�3?5W?ø�=e����{7�#R,>������8DE>�᾽��s��-��>�H?�ޔ>�f_=^�>��}>��Ae�>z�g��>�- ?sA۾4��7[d��Uu���Ǿ��$>(ސ>o&�Zx*��-����p�g�<��='J?.�?���uľ��'��O��e�>��d>��!��W�=��>I�0�ZϮ���9�>ν J~=Y��>��?��1>@�=6m�>������K�]�>ϲ<>�'>]�=?�d%?#���Ȕ�A	��a2���p>���>�>os>d�M�b�=F�>h�^>\��]2���}��~A��-Y>
?�ٍ]��Q|�1�v=�y�����=��=02���<�X�2=/�~?g��*䈿�뾐c���lD?&+?\�=]�F<��"�5 ��2H���?[�@0m�?Z�	���V���?�@�?��p��=!}�>�׫>tξv�L�t�?	�Ž�Ǣ��	�((#�`S�?`�?*�/�9ʋ��l�h5>�^%?J�ӾOh�>~x��Z�������u�f�#=O��>�8H?�V����O�g>��v
?�?�^�੤���ȿ3|v����>W�?���?f�m��A���@����>;��?�gY?qoi>�g۾=`Z����>ѻ@?�R?�>�9�~�'���?�޶?կ�?�E>�@�?�Q#?�>p/��B;a��������F�>b�5����>���>���>����}]���%�ɮ��\P#��ޮ>�e�;U��>�ҽ�_����>�
�n��j�'��]�>��>F,.>6�>@��>�h>��>�ӭ=XN<�W����Ӻ�L?]��?Y���n����<�ڜ=��]�#.?4?�_��1о���>�\?-ɀ?�0[?���>��l7������\W�����<~K>"�>ǀ�>+z���eK>X�Ծ�D�ܘ�>y��>�^��jHھ����a���m�>�h!?���>�ȯ=��!?�G?D��>J�>Ő@��@����I�}r�>��>��?Qc?Q��>?׾��"�:���٭�;�X��=>F)o?��$?9��>o���[}����t�����P�l=n�~?W�k?B`����?)�?Oq?w6R?��>��!�Z�Ͼx�0<t��=��F?�H��X�m�(�D��(�<z�?et3?:��>6޼��k�u��$2�N��j?��I?�&?�ɾ��R�l=�� 5=�,���i5=L����R�}K�>b�>��i�r��=�ͪ>y>d�龚�n�@�>V۴��B�>Ⰰ=�c���;=<$=,?��G��ۃ���=W�r��wD�#�>IIL>N��I�^?�k=���{�����x���	U�� �?���?Wk�?=��J�h��$=?�?\	?'"�>�J���}޾g���Pw��}x�Xw�v�>���>ޟl���?�������nF��6�Ž:�^��>���>t?��>cs>���>�nܾ�'������^�T�B�N��9��^�:C��8��/����)ƽ�g��ev(�k�>���!��>F�?-c�=w�>�Ӕ>���> �%>�8>	R>��y>`@�>1p�=+q�>�b>:�g��R?W���P�'��
� x���MB?��c?>��>N
a�w������h?/�?�B�?cx>�h��)�J�?���>����ɕ
?@�E=Vi���u<�귾��$��+-���>��սu�9���L���d�#?�?�L����̾rO˽��a�.�-=�F�?�T?�,�r
J���l���8��[����=X޶�I�������f�"ܓ�����L�����6���>ׂ ?��g?�m�sӾ�;2���P�.�5�f�=~��>zb>[�>���>���A�N[B��;4�EO��,?��]?1�=���?��7?7�;?yFF?&�>AT�>���
͆>	Z����/?^]?f��>m*?�6B?*y+?l�)?,}�>M%�<z���wҾY9)?:X�>d�?0i�>S�>݉�G���U<i>_�v���;P½�=/В=�j�=&��_�=�?�>�W?��I�8����k>�7?��>0��>}���,��=�<��>:�
?!D�> �x|r�qa�{V�>���?���E�=]�)>���=���QsҺ-]�=q�����=9��}p;�i�<��=9�=��u��z����:�o�;���<.t�>��?���>�H�>g>��"� �n��X�=cY>�S>�>�<پ}���#���g�Ty>x�?�z�?'�f=�=��=�x���R��f��������<U�?hI#?fVT?ٕ�?)�=?�j#?��>�)��L��h]�����~�?�?/?��=E��A־��Ұ�����l6?"��>COZ��4��&+��$���v��8=̼"��)f�E��Z�]��>>=����e <��?�ũ?����.�4�����c��4=t���)?QU�>�A�>��>��'���K��;�w�(>J��>��O?���>]?$Z?�G?��.>Y�>�"���#���Qp>xm�=��=?��?J��?O�D?3�>̅>r������]����u�B^�&�=_S#>�o>��>#T�>���=�}���H�[͇���=S��>%
�>(ǿ>�7�>�z>
��=�I?ҳ�>,����v�"S���퀾�{�K$u?횑?�_*?TB�<�����D��U��v�>��?�T�?�i'?:�N� �=]�ռ�ӷ��zu��>r��>|	�>Z�=\�N=��">]�>�)�>NW�����7�Y�9��<?t�E?A;�=�~ο����$"��콾L�(2����%��>�)K��ϓ=�Z��ؗ�Yhz���$��۞��c���)���=$Dɾ�2?g~=~�B?�<�XR�n��<�3F<�\4>���_흽�z=?OC���h=."Ƚ�K.=%;��7G�=dk>WU����˾��}?d1I?��+?t�C?p�y>(>�e5����>^����H?�5V>�O�-����;�|������\�ؾ�I׾g�c�"ß��K>�hI���>�93>�!�=5��<�=0t=Ǥ�=�T�T%=�;�=HR�=�Q�=��=��>��>E6w?ޞ��~���w;Q��d罩�:?�R�>�c�=��ƾ�@??>�7��;���V�&?+��?�J�?�?.�i��Y�>"	������"��=Н�;(2>)5�=�2�b��>�J>��.O��m_��n+�?]~@ߘ??�㋿i�Ͽ#�/>�\Q>H竽@�m��<W���r��gT�@{��F?�9��
�XmQ>b7�={ž<J�^3�=�h>���=nռ<�*{�kFa>[��D߿�Z?=�(�>*h�>j�o>��P�����r�
>�P>���=�z�ܯ=�9��/<S� =S,�<ɤ=���>�?�/?&pd?�&�>w�j��UξY�����>���=��>��=C>�>>r7?_�C?SL?�>�>}�=���>H�>��+��m����jҧ�UE�<2�?Æ?=�>Xe<S�C���)=�9���}�?)0?��?J2�>hU�F���T&�(�.����������*=Or�WU�=����~����R�=Im�>���>��>qYy>��9>Y�N>�*�>�>D��<ma�=Y㏻O޵<����=ں�����<�ż�����0&���+��/��;��;��;�3_<[ �;�$�=ap�>a�>Ie�>2�=����(2>N1��}SL����=ԧ�0�@�{e��}���.���9���<>�\K>@2������U�?wYZ>�>>���?�s?{>lz�8�Ӿ����W�b��GT��ҟ=�}>7��68�(]�K��Ҿ���>�e->Q��>���>�@��K*�s�=���)�2�1l�>Gh��*/��߻L���e�+g��p��^e���=*?w�����I>ޫw?�G?�|�?�9�>D�6��Y龔�>�툾���<9=������|)f���
?�`?���>Qɾ�R����"a����>e�	��L��Ӓ���3��Cf��¾�¸>�ű���ܾ:�3�����ͮ���UU���|���>��P?���?usY�bu���pT�C7������?�c?��>���>_S?C6����1�G���=NOc?i��?6�?���=hڰ�y�,>"��>��>���?f�{?�t?�0��v`>��g>k��>U�_=D��{��>'£>sS�� Q?�1?�N?�����%"����LT�����1����>���>>�G�>��/=~�=���<V��=[o@>�>�LZ>'o�>Iz>����+���7?�@[>�Vg>��7?M�w>���<�:C�n�>�65� �)�����C�z�����g��=Gu[�.ḽ�-�>�������?#{�>�����?.����=�k>�>Ҥ�� ?xZ>A9�>F��>�Nq>��>M��>iΥ=jEӾ�x>����c!�A-C���R�C�ѾO}z>)����&���;���}?I�@n���g�j�
.��W<=�O��<�G�?�����k���)�Z�����?�Z�>w6??،�c
��3�>���>�Ǎ>�K��x����Ǎ�Fh���?���?�;c>��>D�W?%�?�1�3��uZ�,�u�l(A�e�O�`��፿�����
�����_?��x?yA?�Q�<�9z>Q��?��%�Sӏ��)�>�/�';�K@<=g+�>�)��%�`�w�Ӿ��þ�7��HF>��o?9%�?wY?6TV�+-��-]><�??�G-?s�?�9?);?9���D? >)>�C?5J�>�1$?��C?s^?Ʋ�=ΫN>�<8<S�=5ս�)����(��=�ߟ�5ܰ=x���P�V<q�>�����8�<������.��&�a�8�<詻%
<�[>�{�>�	]?���>���>P�:?���SD3�v񰾓J+?�@=2=o����z ����K>��i?� �?\?�?n>�A��=�`Y>X�>�@,>0�[>eI�>?$�QcF�tP�=%>S�>w˟=On�{\������<��4��<E�>�?/u>�>���%>�jr��2��!>~�%��|k�����#�Gkݾ�iB��F�>��K?��>k�=�o�i{,�s�f�p�@?s�D?�Y�?�T?���=Y���bD������C���U?W��><p!�Cn����Ġ)���=���>�w��ק��0->)��9��Qk�G����39�=���p��<�*���޾nȀ����=c�>aj��� �֋��z�����L?hI�=����LI�#��B�$>�>F��>�n8�#���F�Q���q0�=��>ص4>��켜��~�B��k�`	�>�i<?��7?���?(+��8 k��_R����Poþi=��Q?j�(=8��>���=�'�>*��o�����[��	k�9�?�l�>�E�8�E�$vD�g�1�ۛ*����=�)?5�>z	?ĭ�?��?�_�?l�P?��?�>&���? �+x5?�=}?B��=��f��J�T���X��?E ?�c�LY>�)?�#?<�/?�)n?�Z"?��>V�
��}���y>>{$>>ZS�{��"z�>�B?t� ?�SE?��z?��s>!C���)���;���=��u>wOK?�q?"�?�Z_>Ļ?༰���ν���>�ɘ?��?k�l?HZ>6y#?+�>���>~h�=���>� -?P?}OQ?��e?��J?� �>R�Y�%J�_`R�����g�'�<9�=	�t=:k�B�i���#��?&=6��W8��o;B�>+�����u�Z��<�Y�>��s>镾�0>žN���nFA>o#��`��sf��v:�q?�=�g�>�?�;�>�&$����=bѼ>΃�>��iA(?��?�?��>;0�b��#۾�pK���>vB?K<�=)�l��y��r�u�i=��m?��^?�-X�f)����b?x ^?����<�[lľ�3d�5,꾱�O?ں
?��G�D��>�~?��q?(��>CSd�R�m�Cޜ�[Gb���l��A�=�:�>�O��Xe�8P�>��7?7g�>�,d>Е�=Ö۾Kx��ğ�6?���?��?��?%�)>Ƅn��'� �������v?�>���_�#?��=�^Ѿ�9�-V�̾�T�P�ʾ
����ƾ5A���o��|��qn>P'?�kv?��d?��x?��
�N�W�nk[��s��g�Z�&��\k�~�6�Qg��H���b��^�z��@Ǿw�;��~��~A����?P�'?�0�ٿ�>����S�̾B>-=��6�Ǚ�=U����=?=Z�Y=b:h���.��H��F ?m�>,?�>d�<?��[�V2>�U�1��7�I���̄3>b٢>��> ��>��:��,����*ɾ������Խl�v>ňi?�?`?du?��2��������p�F��G
���7>�c���G���������&�d�!�	s��� ����]��z�e�s�?t��>-��>P��?��^?��� ���V%1��O�s�>���>�ؐ?]V�>5�>�/����L��7�>F�d?�U�>T��>���� �C�h��(�����>�f�> �?�]>A��g)]�{~��������6�?�=oMk?����)v�nq�>�qK?�{�<M =ȇ�>��)�����T��m� �Y�|>��>:�	>IT>>]����vYv����|�-?.?����:S>�r�>�&�>���>��?z�>����a>�+,?�\?8�Q?kPM?!(?,��=8j�����!�	��:�E�>�O>�I=�k>��W����ED�j1?>�GM>��N=kѽ�5��k'�;]F�<�#>6�>��ڿ�OP��徠L��+��
�Ȝ��/�T�|���?J�QJ������v��f��r��8��X�w����n���?�c�?"�z�#����蚿w�{�;���3C�>�w�($�ᇡ�q�ɽ�������]��M�SAj���`�+?�d��뭴��b���Z���?H�?�D�?ǁX�5;
�f�x�,�L�l�i<��Ӿ� ����ݿ�]@�Luf?'#?,Ͼ0=O�>`K
>�}�> { ?G�����ʾBsL>��?(|?Q�(?�2">�׿�ֿ�hM>�@�
@|A?��(�M�쾝IV=w��>Ŕ	?i�?>�R1��>��찾O�>h9�?���?�:N=��W���	�ʃe?N�<E�F�)�ݻ���=;�=�=���\�J>Q`�>�d�ngA�C-ܽ��4>�>#�׵�Jx^����<c]>/�ս��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�����ſ�u=�Б8���G�&��������K{�ļӽ����+������`�f�>�.�>���>�s�=*dE>+�`?w�m?+��>S�>�T��ɨ���վ�3>ٸ���(7��{:�J��A5���׾�a��9�����p',�����8;�
58��CQ�3N��c= �x�[��-H�1e=?S�>[ӾfvU���P��/Ⱦh`�����<*��۵־އ-�vt��Ξ?��A?�x�-�E�%��s<a�׽i�f?>����� ��hоt�3=Ò�Q�M;�v�>��H=�����-�j�D�2v6?��?�n¾����St�=����c=��?���>{��=kS>j�W?*�b�����P٩>,>�!�>��>�j���8���y��5G0?7jl?��D����d�><���;���U�}=y>�xܽ�m^�s&l>�=ZŒ�b�ӽ.Ż�>e W?���>`�)����`���9���==i�x?ג?E@�>e�k?��B?`�<�m����S���� w=��W?�+i?ش>ª��n�ϾHx����5?��e?��N>�Th�E�龏�.��R�x0?j�n?�b?6F��q}��������i6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������(*�= tR�h>�?q�?����d&= 	 �}/z�2F��[M��#D�=N:=P�����	���I��+;@��H-�5�=��>#K@L�O��m�>Q�1=D�ȿ5�ʿ�W��O ����O?�I5>|�Z��~���op���O��[C�xY�
[̽�L�>�>�����鑾��{��k;�𯟼_�>�v�[��>��S��;��嘟��84<��>Z��>���>S`��M����?�b��Q>ο���՟��X?�e�?k�?�o?cs<<��v���{�T���6G?�s?Z?a�$��"]���8���m?�1־��5���A��n��'�>
щ?	�>=5O�e">'�>!KK>��>�e����Ŀ>�Ͽ��,�'��?��?҉徻�?P�?l�Q?և
�d.ÿ!ߠ�;TG��>�q=?��=^��H`�8G�k��i�?�)?�bO�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?#�>��?1o�=0a�>
b�=��O�,�Jk#>�%�=�>���?O�M?~K�>4R�=�8�3/�[F�FGR�9#���C���>�a?��L?�Kb>���c2�/!�jͽ�i1��S�R@�G�,���߽�(5>��=>`>%�D�Ӿ��?Kp�6�ؿ�i��,p'��54?9��>�?��e�t�����;_?Pz�>�6� ,���%���B�`��?�G�?9�?��׾�R̼�>;�>�I�>-�Խ����L�����7>2�B?Y��D��t�o�q�>���?	�@�ծ?ei��	?���P��Va~����7�e��=��7?�0�!�z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?pQo���i�B>��?"������L��f?�
@u@a�^?*�$޿��	��j򾎼>2l�=I�9>����k�4�%]�ϪܼwO�=���=u�>WH>9�>���>ޜy>A>�+��?�&�>2��O���.�B��������J����2�����s �D�f�c���1P�.��\։=<w'=�n9�s����=-�U?7
R?`p?K� ?t3{�K� >]�����=�x#�Q�=�>�>�{2?��L?��*?�R�=UQ�d��X��S5���[�����>*xI>���>~��>麮>9��'�I>�Y?>���>z; >�X+=���=J�M>���>P��>�>m>kG\<����D��1b��A�KR�T�?Ⱥ���WL�;���nԾȾ���;�\%?�2x=С����������ѯ\?������X�M�<�WS?9D?l�O>.꾿vw��D'>�'�(6��倁=
GR��;��m�j&2>�U?�f> u>�3��f8���P�<���)V|>�56?鶾|C9�+�u���H��_ݾi@M>bǾ>��C�ii�}�����Cai�G�{=#t:?�?"2���۰���u�7���NR>4\>�==B�=NUM>nQc��ƽ�H�..=X��=��^>�D�>��/>�o=�5�>�	��|�Z�^�>u�=>��'>@�J?-�,?�n�5���x菾��M���c>���>�R~>�$><M�c��=���>�c>s_2��Vc�H��.�4����>y����J��:�v=����0��=\a�=M����M��,=%�~?~���㈿D뾭j���mD?�,?9�=#QF<�"������H����?A�@1l�? �	�:�V���?3A�?�	�����=N}�>=ث>ξ��L�4�?5ƽGŢ�r�	��'#��R�?�?��/��ʋ�'l�r9>�_%?\�Ӿ��>Ҧ�hU������u�?'=	��>mDH?����TWO�>�W\
?5�?�/򾲢��.ɿ�v�R�>�?�?��m�-����?�b�>��?��Y?4�h>D۾�Z����>�@?�4R?�]�>me���'�T
?��?���?8IB>���?�Ћ?��?�H\�$����G��P��� w�h��*m�>`Ͼ�M�O�M$���y����:�[���M�rL�>фh=�O�>�Dv<�����v�Φ�c!�����<��p>�M�>���=���=mܢ>�#�>�>L��;L(ѽ[#��'��%�N?���?����i��-�#~�;�`��?%�3?�݌=����>�(Z?!�v?ٲg?���>�L�鑿�XÿAת�N�0���=��>��>�(����>�7ؾs�@����>�b`>�1=*��)����/]����>�\4?��>��1>�� ?�#?i�j>t#�>�^E�k8����E���>��>kO?��~?M�?�Ϲ�	\3�	���䡿ސ[��6N>n�x?2R?X>$��������D��I�����~��?{g?��彯?�5�?��??-�A?�(f>��_ؾ����6�>��!?I�ӷA��K&����t?�J?#��>��x�ս��׼��k��"�?&,\?�D&?��'a�þM,�<s#�\k_�q��;�;D���>_�>����x�=�>�Ѱ=t*m�8,6�E�e<�E�=���>�`�=�7�_@��0=,?��G�~ۃ���=��r�?xD���>�IL>����^?hl=��{�����x��	U� �?���?Zk�?^��@�h��$=?�?S	?m"�>�J���}޾5�ྺPw�~x��w�^�>���>�l���K���ڙ���F��]�Ž�)�t��>G��>Q; ?B��>I�>���>����=�J@��񐻾ٖc�W�{�?�j�5�Ku�b���/�q�$=@վ�\�r��y�>,9��ƽ>p�?��<>�t>A?19R��љ>���>j|{>���>��X>�3�>Ő>x���9��KR?�����'�}��{���x3B?�qd?<1�>xi�������h�?���?Ss�?�<v>h��,+��n?�>�>B��,q
?�T:=�7�8�<<V������2����B��>!D׽� :��M��nf�Oj
?�/?����̾�;׽͇�����=�#�?�0?`$�N�H���k�pm^�`O�)ʽdrN���I0���t��'�������;���M0�K�=է&?ac�?3 �ʤ����c�b�w�A�#Q>+��>j͘>���>�x)>���l�8� �`�h+��������>Uz?���>auB?a�:?�g?�Z?}m���C?A����P?!>���;]�H?��d?�O?�)S?��3?�[?��>�?����¾�L���Y�>�}?-4?L�?�~�>z⫾�A>P��=Pͱ�p����x�:��>f����z��р>4}�=eɄ>BW?���)�8������k>�7?��>���>���$��Sc�<	�>��
?�B�>� ��{r�Ab�]U�>Y��?����=N�)>L��=Ym��i�Ѻ<R�=������=�q���i;��B <��=�=Ut�8a_�dD�:W��;�k�<�t�>1�?���>�C�>�@��1� �S���e�=�Y>�S>�>�Eپ�}���$��{�g��]y>�w�?�z�?Ҽf=��=Ȗ�=�|��wU�����7���-��<�?XJ#?XT?Z��?��=?Vj#?�>+�]M���^�������?}",?y��>�����ʾa�{�3�n�?�[?�>a�׳��9)�=�¾��Խ��>C]/�4~����VD�7�����넙����?Ͽ�?ONA�#�6�Li�L���*T���C?"�>�U�>�"�>N�)���g�"��<;>��>R?�7�>��O?O#{?��[?�oU>vo8�/��jٙ��S��">2x??���?=��?:y?x|�>�9>��'���߾�O���]�'E�7��T=Z>�Ӓ>\C�>8�>���=�=Ƚ�4��S�?��.�=�b>�y�>�O�>��>��w>���<�H?�8�>﮿�=��"����!@>�$u?9]�?,?ۦ�<�3��-D�tT��ə�>�c�?���?@9)?fFZ���=�߼4N����o��?�>��>�K�>��=\�>=�>@��>���>/b������8�w�@��?QF?���=Ԯ��򮂿#[žK��J8�E�׾�ܠ��m/>����"�F=��M��.������A�w��b��,�C曾�hܾ�����R
?#�D=���=���=ڃ�<X�今�@�6�>�:s=�����ӽ�Sv�K��=�V���,�WO.�CK�=�d^�5�˾<�}?v<I?	�+?��C?�y>n->� 4�Γ�>@���g>?pV>�P�`����;������$��X�ؾ�j׾�c� Ɵ�)U>+fI�H�>K*3>�8�=H!�<!�=�5s='َ=I3T�^�=^*�=O�=�h�=-��=�>)K>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�96>e�>9�R�ww1��P]�w/d�V�Z���!?n�:�Y%˾gN�>�u�=�r޾�\ƾw4=��7>��c=4-�/\����=�8|��;=-us=�:�>=gC>s��=}��M��=�HH=���=�&O>�a���I3���/�S30=.�=B�c>zN%>d5�>2�?Es/?xj?���>gcg��ɾ�Ѿ>è>�	>2d�>&Հ=Bm>���>)�6?nC?��U?+��>+|E=���>�Ŝ>�Q/���j��R۾r͖�{����?���?e��>����\�uy�}n2�������	?�],?��?�;�>+���߿�pn�Z;V������퀽�(�F��~�C������ �CT�a�6=��3>�@�>�r�>�I�>���=N8>W=�>3>�I>�,�=E�g��>�A�B�4�>z��=8�<.Tx���K���f������a<XE���A��Xd�DO��/�=���>@�> z�>���=f���~/>����آL�X��=Ǘ��^*B��d� L~��/�܁6��4B>a$X>`Ȃ�e ��A�?%XZ>�x?>tq�?�!u?�>���n�Ծ�P��Y�d��Q����=%�>��<�2;��(`���M��[Ҿ�;�>˪y>� �>�~�=#B<��7M��ku>f���\LH��R6?��$��^R�&�>_P�Ө�e'����h�Aj>��_?q����S>(�?V�)?��?��>r�Y�ꇾw
�>?��fJt>;�Y6/�d[����?-h??�B�ަ1�WH̾Q���ݷ>�@I��O�n�U�0�W���ͷ�Ԓ�>����e�о�#3��g�������B� Nr�V��>g�O?��?9b��W���TO����%���p?J|g?-�>�J?BA?�$���x��s���x�=�n?���?�<�?_>�>^B��K�>�<?P�?G��?7f?A�����>��>��_>����eM>��>a��=z>L$? �?�\?�\~����3�vx��t��I�=�c>�'�>\_P>�	�>ʩ<>5�=�����<(6�>��>���=Ղ>�X;>ڦ�R=��x+?Fa�=�:A>�?�٥>�ii=�>���<�&>���#c�K���"���(|�����.!u<mT>*s�>qVſdS�?�G�>��K2/?㉰����P�>�$��<冾�F�>I�����>E�>2k�>��s>��I>�7��[9Ѿg}>'���X"��QC�G]P�J�Ҿ;��>�h����*���
��� ��9M�Ƹ��[�gni�E��~�=�N�<�]�?����k� �*����TE?���>RU4?k���[��,?>qN�>���>!!������쏎�\l���?���?[;c>b�>#�W?��?Ӑ1��3��uZ�p�u�o(A��e�G�`��፿	���v�
�)	��>�_?0�x?�wA?wM�<,:z>��?C�%�'ӏ��)�>|/��&;�??<=.*�>�'��a�`�=�Ӿ{�þu5��IF>�o?�$�?\Y?kVV�߁Q�� >��6?p�/?��u?��4?2w<?�^�4�$?�50>�.?)�
?�5?R(/?�"?��<>�c�=����$=�e���	��A�Ͻ2�̽NB��8@=r�z=0�|�ʰ�;�
=+��<	�޼*���$9G8dA����<Yf7=0��=���=�H�>��Q?���>j<�>ߗW?L=/��1��۾��^?&0>�r���[��������D>o]?��?�d?&>�3���.�6go=m��=Kw>F>�>��>�]I=����՚<��v>���=�M�=pT�;踐�������~>3�s>'��>�0|>'��ȷ'>�|��N1z�;�d>,�Q�-̺�Q�S���G�y�1�G�v��Y�>G�K?��?О�=1_�X.��PIf�(0)?�]<?�NM?��?��=x�۾��9���J��>���>	Z�<��������#����:�l^�:��s>�1��(���a>a���޾&�n��J�����N='\�"�S=���/־'(��Q�=D
>Ѥ���� �x��zʪ�;9J?_Dl=�W��,�U�:k���@>}��>�>�=�f�w�Ey@��t��zn�=߂�>�;>����P�F�G�(b���>1�:?/�L?9��?�<���S�gZ�e���'���>6�$?;��=��6?��p=?sؼ�|L��}ξ�"��{� ���>s�>�}޾��L��/о8u�� �4i�>侵>(�>�t�>���>Q�?Z�?]�>?b��>|Fn>Ⱥ�����V":?��n?<-P����|��JH8���F���?��?�C9�@��> [�>�7?��K?g�k?D�"?P�>EԾ՛���Y�>ZeT>��e�����>�>�"?u�>�r?]n?��#=w�)���ƽ����!�=��>�>L?U?��L?\�]>��>�?Ӽ.lV>̶�>5�?_ �?V�q?�ܿ=+�?��=���>[0�>���>���>)�?:|X?�?;�_?���>y�S�j�)��/�o�2���'��=�{2>��=j�����Z�=j�6=g�'��b(�T˅�V�ý� ��"�qÙ=�`�>&�s>�
����0>��ľ"T����@>v���!O��֊��:��ַ=���>,�?N��>]#�W��=���>J�>���z6(?,�?V?�c$;�b�{�ھ��K�\�>	
B?��=,�l�������u��h=��m?�^?�W�^$��`�b?��]?��򾷱<��vľa�b�}��~�O?�
?�VF��/�>�`~?"r?���>6�e��m�e᜿�`b�u�k����=4�>[��,!e�jH�>�`7?�a�>8e>���=�ܾC�w��X��5�?��?�#�?5�?x�)>Wn��W�Pw�A�1�{?`��>E ̾@xP?j��<Q�Ѿ�r�4����,�柾�b��`1W��1���k5��&��߿E��y�=�z?h\�?E}l?Z��?T1(�ߊ@�6�[��ۊ���=��m0��� ��A�[�JLd�םO�������y˹�w�$�(���3C��?�,&?o4��n�>Մ����c}˾S�=>����4m��ƣ=%�����2=�*Q=?�j��=3�:n����?y�>�d�>e'@?��]�\4;�k�1��=9�ֳ��R~!>���>��>O�>���^(���eʾ4���&ݽ���>�_`?�)E?�Qx?�? ��4(�{���T*��6�}��9s>66">n�>4<��ΰA�s���:2��Wq���������u�8��<�-?��e>ٓ>���?�?�޾$�������P/��S�=fX�>�`e?��>뫏>ֿ����>Pcj?���>��>�ʡ�3n�������E�>���>o�"?��>�)�5M�����s�}�F�!��3�=�n_?�a�(k��J4 >��l?��@�<f��>B���+Ŭ����[���m=\80?+��=�>봣��4��}Ձ����k�1?{�?͹����:Q�>���>���>O	�>}�?e�>6(���o�=�5?��U?��[?џM?� �>�n>��X��*½� ��>=�o�>���>�1=n��=�&1��=`��K`=�~	>��2�-����<@ɵ��a�=�N&=��r>�wۿ1dM��޾Z��G��d�∾$���F���ڑ�����7����<��'
�GdZ���i��Ê�|�s�F[�?��?�s��o���5f��B{�)����>�>x����G����S�����&���z?��>R��$m��hg���?�b������
묿jo�L�*?5�?�u�?�a���`�#��v!>^�{�Ț8��þ'̥�Hn̿`��_a?i�?��Ѿ��ҽ(��>Z>~Sw>�D
?�抾��ƾ�$==��>���>�5"?�g��b��U�ѿ�>=n��?�@�|A?T�(����00V=1��>��	?��?>�U1��F�����T�>�;�?���?kM=Z�W��	��e?~�<��F�p�ݻe�=�;�=�?=���ߒJ>tU�>~���LA��:ܽ�4>m؅>sg"����1�^�钾<؈]>��ս�;��5Մ?*{\��f���/��T���T>��T?+�>\:�=��,?W7H�`}Ͽ�\��*a?�0�?���?$�(?3ۿ��ؚ>��ܾ��M?_D6?���>�d&��t���=�6ἶ���v���&V����=Y��>X�>��,�݋���O��I��\��=����Aȿs8���1�,�;�R������c?�S8[�"E�����O���G�C�h�=b�7>��>G�.>>�>`�)>�GT?��f?�ҷ>J�m=�5�4����Q--=�;f�њ!�$���'S!������Q��'4�Ur��O''�ZJ��f ��O�)�Z�R�[��c��
���^�'];�j8?ak>R����Z��ru���㾈���0�<�ͽ���؈3�{Yr��?ӎG??�q���J�������=񒋽�1T?Z2x�w��WG���?>0���
Ո�6��>#>.,��B\��QP�"�H?.�"?���=�+���h>4�ƾ�>!�uf5?a�6?7�>s@[>�	L?�X���=���(?�x�>0�>��?86��G�����:��?��b?�Z�=�b}����>��Ծ��w�0����=G�#��3���>�}޽$����Xf>!<�f/H>?(W?���>��)���mb����t==D�x?Ҏ?�*�>hyk?Z�B?���<>e��m�S��!�kDw=��W?-*i?I�>ߋ��	оH��ý5?��e?��N>fh����r�.��U�� ?��n?^?�����u}��������n6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?p�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������̦=ي��	�?l��?բ��Z�I>{����}�Ԑ߾Ӻ:��j�8�u=�M<��P�5<�Zq���a�q#�O�{<�:�>�@�I���	?�%νx/��U˿y�����о� �B8?��>��������~�w�H���w�?�ڔI��n�>z�&>��0��Lg�;x��l�7�,@׽`��>wv����>��;پ#�=��ک=_��>���>��>.z(�|f��?���Ϳ9��������F?���?���?d�?�T�>���b� }��*_?ہ�?
W?�왽�����g��b?h�ξr7l�<�S�I�^���b>g+c?6�>@L��B�8'���I>`�@>�u�Ӳ��w���Y8�ݶ�?�%�?��;0�>b��?�-3?#�1�?���a�� O���Y>WE?�)�E�޾�H��P�1�ƾ�/?��$?�����V�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�$�>��?�n�=�c�>^^�=�𰾠0-��f#>�&�=.�>�%�?%�M?M�>SN�=[�8��/�^ZF�AHR��#�j�C�L�>��a?��L?3Hb>M��� 2�!��mͽ�a1�>\��[@�X�,�Ó߽)5>q�=>>r�D�yӾ�?�p�'�ؿ�j���u'�"64?@��>�?"����t�1�P8_?�x�> 5�S+���&���K���?5G�?B�?U�׾�=̼b>(�>�E�>q�Խ��_{��^�7>��B?x.�gA��W�o�.�>���?}�@�Ӯ?ti��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*�	޿�	��^��c!��%s@>��3=�rA>���Lo�<��N� U�̽��=�t�>-J�>�m�>�>�U>l�?>�-��^�%�ș������ =�p�=��������
_߾7%����������$�H2N��<����p�D`	�iB�=\�U?g'R?*p?�� ?9�x�M�>�����%=�#��΄=�D�>�}2?��L?��*?v7�=�>����d�Pb��R=��jև��y�>�9I>�[�>�I�>���>���7�
J>�2?>@�>�$ >s�(=�[��+G="O>�k�>��>Gf�>կr=T��<�ʲ�j���[���X�~ҽX/�?��¾"E^��f����i�!�QEP�]<+?#��=eW��&iֿ�Ϥ�^_? ������1C��֨=ԑ>?�M?In>�K��2�=j�x>�J;�_��/��=����%Q��).>"??3d>�#t>�3��Q8��*P�;ˮ��G~>��5?����6��u�?I��Oݾn�N>���>�jn�Fe��˖��~���h���v=�+:?�-?����1#��t7t��x���T>�]>+{$=룱=��M>O�\�*�̽�(H��,=M��=?�_>�R?��2>���=�߫>l��H�N�ϲ�>vF,>?]7>��@?&�$?���a�b�o���'4��y>0��>�h>��>R�B�aB�=�e�>�aU>I�;�Dލ�=F�%�<�W+`>�kR�ۀ^�E��슙=�3T�p�=��=E��W�C����<�~?���-䈿�뾙e���lD?i+?�=��F<��"�= ���H��4�?i�@�l�?��	��V�G�?�@�?�
����=}�>׫>�ξN�L��?_�Ž�Ƣ���	�~)#�GS�?��?�/�Zʋ�l��6>�^%?ӰӾ}��>�������҈�^t��n=���>P0K?��=T����>���?�o�>��龃Ϣ���ʿ��x���>H>�?XW�?��k�J���<��_�>K�?�`?$�X>#�;�\�".�>�4?'�X?m\�>����,�OL?N�?n�?J>�Ў?#n?�A�>�rL��L�G��䑿�U8���=9QK?ZX�>��6����VW���C���:��Cؾ�v�>�f�=�D�>aJ
�p���Uh�=ZJ�Z\����Y�$>�t�>-:S>�> �?4`Q>���>���=e R=!P�<�^�B!L?ԇ�?��:�m�cc�<��=�M_���?�A4?�4_���ξ��>eY\?�ր?�^[?<h�>�o��������&>��:�<��J>h(�>���>ۊ���-L>�Ծ$�B�/Ǌ> �>�]����ھ9����YS�>�}!?!��>�߰=�� ?��#?�j>�B�>�_E��3����E�L��>
��>�N?��~?Q�?�Ź��g3����[ࡿ.�[�N>^�x?|O?`��>����y���DF��9I�������?vzg?_t��?�)�?Y�??��A?�:f>:f�f�׾�����>�"?��~�A�&�[o��?��?���>@[��jgսM7Ѽ�������K?Kv\?ߞ&?�<�VD`�w{ľ-�<	�#��#`���;J�-�';>N
>O�����=a_>>��=��i��6��A<�A�=�K�>D��=:�4�-֋�2=,?z�G��ۃ���=��r�AxD���>�IL>����^?gl=��{�����x���U��?���?Yk�?~��=�h��$=?�?X	?u"�>�J���}޾<���Pw�#~x��w�]�>���>�l���J���ҙ���F��R�Ž��7�>jj>_�>��>.�>[e�>1f��-�8��ښ�٭�f���V��H�b��q/�F���o�Qߤ=��Ⱦڐ|�#�^>�����>؞?���>V��>�>��3<���>;�>�[>���>��)>t�>�tD>��=��k��Q?=2ľ�+�MS�������B?�g?L��>LU���h��3��Θ?%_�?- �?�#i>�m�q-���?CE?��u��s?ԝL=F�׺Qe��A���,{��z�Q�,�>D�����>��@B�ԕh���?�O?	6����Ѿ�½���"�=�҇?g1?5�,�(/E��Ck��d��oG�E߽<�!��h�l�?�A؀�(��Ds��|�I�?����=ٴ?֎?��0>�2�,�aJ���V�U_o>��>ڮ>~�?��4>d
���1�*�]�� !��6�=3�>L6k?(/�>��R?�<?Dwj?a�~?w�V>�C�>3x���'?jPy�![>��?�*R?�#?S?ZX,?Gt?eE�>�6������`��0<-?8s�>(?#R	?�L�> ��c����|u�6E���.`���=ƅ>�⦽�}N�8�ڼ��<�9>X?g����8�)����k>ρ7?M��>[��>���,��}��<3�>v�
?�G�>�  ��~r�+c��U�>���?����}=��)>t��=������Ӻ�`�=������=�*���r;��v<�=���=�iu�������:p��;�~�<�l�>?i��>oV�>@��(� ���ϊ�=N=X>��S>7$>��ؾ�|��j4��_�g�Gy>K]�?#l�?s�f='2�=���=?���Ǿ�f	��ν� Z�<�?�l#?YT?Pr�?l�=?,�#?Թ>����@��\<��t0����?�l+?-SY>T0�B��٭�pq/�M:,?�(?��c�����3��辤]5�Y7>'�9�Ņ�5���.>�"F�=�S��VO���?��?�禽qH�0`�q����R}��tR?=�>�$�>V�>��$���d��,	�\�>4��>;rK?��>��N?V�u?�4b?(c>>�p2�I���n��S9�;�<8>��??V�~?~�?LDf?-ȹ>��>h����,
龴8�9���q���'&=~�D>
��>���>r��>%�>1�ͽlx�B�Y���=^��>��>�9�>��>QU> �|�N?;��>�׾���h���枾�B�����?:�?�|$?��G=�x��2-0�%c��l��>P�?�7�?��8?����@�=A���<͛���k�*��>f�>�ђ>�Й<�w�="�P>`��>}� ?!���0%�u�'�>쪼�M ?�B?��
>�9ǿ��u��憾� ����^<����0�^��\��Y��\= 坾8�'��'��QK�е��M���3긾%.��}4m����>�t�=)H�=�=��|<���<�#�=�=ȳ=3�s���q<U����_<����H��|��_=����q�˾�}?�;I?�+?A�C?�y>H3>��3�7��>�����A?�V> �P������;�����!��B�ؾ�t׾��c��ȟ��G>RuI���>273>=B�=�V�<~�=�"s=���=�XR�m%=n"�=�R�=�i�=^��=��>;S>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>JS>�%>mAS��.��+^�&v�8|a�uC(?�D0�������>��=�վ�=��(�=�O`>QÉ=��׽�?d���=�l�ׯJ=�JL=���>��5>@ڽ=�>ǽ}w�=�	�=�^�=#�>�l}����F����M=�>B�q>�\3>"o�>� ?cq8?y�l?1��>9�S�,*þ�ľ���>R��=�`>���<oh�>B��>K7?jAH?�e?\��>�r�9�>>N?�
s�a��tv���Z�4s?r�w?���>��ӽ�܋�����5��0��� ?��0?uw?��><p��s翳�T�)�1�Br��i��k���h���9���L���s�����G��f��[�>�Y�>�SB>`Ŵ=�?0>wX+>��>*�#>�G�6?�X��n���0̽}�=?��=v!4��(+7���.�����-(=uP%��{��.�=��»/S�=~L�>��>��>ob�=<!��W0>�����M�y��=Gg��F�B���c���}��.��L8���@>��U>{N���C���?��W>aZ@>��?��u?D$>��	���վp����b���T��h�=w~
>�8���:� _��M�ȺҾ���>�S>�D�>��y<2�>���8��׏>����G��	?s��t��g,���F�p9��n����u�� ӽ��c?f����V>�A?�@?xP�?�?u���?���>�=�蜽�B=+j-��˾��:s�U?Mm*?,(?���zIS��H̾.���޷>�@I��O���/�0�e��=ͷ�\��>������оi$3��g��������B�)Mr�'��>-�O?��?�:b��W��EUO����:)���q?�|g?,�>�J?�@?�$���y�wr��_u�=�n?���??=�?a>�+�=ڟ����>�9?�D�?�z�?Gs?V�9�Xl�>0�<0t>2���ԯ�=�>�ר=���=3�?F	?�?�ᚽZ
���ﾋN����`�+�<0��=�>2�><az>�a�=^a�=�Н=��W>�f�>�Ό>�Q>
��>	�>��վ�K5�"[?�1 �+ �>!�(?%��>:��=h�Ͻ��>ǁ½-tN�#��7P?>�!���?�HL7��yn�;�q>,�>O������?7O>k��%�?K������"�>�Ž)t/�N{�>�"�>��6>�0{>��?���=j}>:^�-sܾ��>b3�٤"�	;��rB�����ʁ>C������4��/ ��4R����a �?bm��%��ҩ:��s=q\�?����a�o�(������>��>�86?uIr��c��;>>(q?(Ғ>�S澎���+G��\��?��?�;c>��>K�W?!�?ג1�/3�vZ�-�u�g(A�+e�R�`��፿�����
����+�_?�x?)yA?�R�<(:z>Q��?��%�^ӏ��)�>�/�*';��?<=o+�>*���`���Ӿ��þ8��HF>��o?;%�?xY?2TV�G�ں�CY>~i8?�?qZ~?K�E?��L?�lٽ)$?B�>�?S�>oU)?��1?�O?��>��Y>��@=���<�J��-������T	���@ѽ��<[�m=�-���m�zp=l��=�Y'��^�R2=^�Om����a=��|=�`�=
S�>R�Z?���>�i�>m�??�� ���*�����29?y�G=����^r��s`�Alʾ%�?>$r?Qv�?!�`?��>4{E�+O��7>9�x>�~>> �u>�&�>|�E�r����=�3l>?L>�)�<����(������e夾�?j=��^><��>��|>�h���(>�+��Оz���d>��Q�m\���S�U�G���1��Lv��K�>��K?��?�Ϛ=��#���u;f��%)?'v<?�cM?v�?�֔=
�۾��9�_�J�����'�>	��<���ӫ��K.���:����:�Fs>����ק��0->)��9��Qk�G����39�=���p��<�*���޾nȀ����=c�>aj��� �֋��z�����L?hI�=����LI�#��B�$>�>F��>�n8�#���F�Q���q0�=��>ص4>��켜��~�B��k�`	�>�i<?��7?���?(+��8 k��_R����Poþi=��Q?j�(=8��>���=�'�>*��o�����[��	k�9�?�l�>�E�8�E�$vD�g�1�ۛ*����=�)?5�>z	?ĭ�?��?�_�?l�P?��?�>&���? �+x5?�=}?B��=��f��J�T���X��?E ?�c�LY>�)?�#?<�/?�)n?�Z"?��>V�
��}���y>>{$>>ZS�{��"z�>�B?t� ?�SE?��z?��s>!C���)���;���=��u>wOK?�q?"�?�Z_>Ļ?༰���ν���>�ɘ?��?k�l?HZ>6y#?+�>���>~h�=���>� -?P?}OQ?��e?��J?� �>R�Y�%J�_`R�����g�'�<9�=	�t=:k�B�i���#��?&=6��W8��o;B�>+�����u�Z��<�Y�>��s>镾�0>žN���nFA>o#��`��sf��v:�q?�=�g�>�?�;�>�&$����=bѼ>΃�>��iA(?��?�?��>;0�b��#۾�pK���>vB?K<�=)�l��y��r�u�i=��m?��^?�-X�f)����b?x ^?����<�[lľ�3d�5,꾱�O?ں
?��G�D��>�~?��q?(��>CSd�R�m�Cޜ�[Gb���l��A�=�:�>�O��Xe�8P�>��7?7g�>�,d>Е�=Ö۾Kx��ğ�6?���?��?��?%�)>Ƅn��'� �������v?�>���_�#?��=�^Ѿ�9�-V�̾�T�P�ʾ
����ƾ5A���o��|��qn>P'?�kv?��d?��x?��
�N�W�nk[��s��g�Z�&��\k�~�6�Qg��H���b��^�z��@Ǿw�;��~��~A����?P�'?�0�ٿ�>����S�̾B>-=��6�Ǚ�=U����=?=Z�Y=b:h���.��H��F ?m�>,?�>d�<?��[�V2>�U�1��7�I���̄3>b٢>��> ��>��:��,����*ɾ������Խl�v>ňi?�?`?du?��2��������p�F��G
���7>�c���G���������&�d�!�	s��� ����]��z�e�s�?t��>-��>P��?��^?��� ���V%1��O�s�>���>�ؐ?]V�>5�>�/����L��7�>F�d?�U�>T��>���� �C�h��(�����>�f�> �?�]>A��g)]�{~��������6�?�=oMk?����)v�nq�>�qK?�{�<M =ȇ�>��)�����T��m� �Y�|>��>:�	>IT>>]����vYv����|�-?.?����:S>�r�>�&�>���>��?z�>����a>�+,?�\?8�Q?kPM?!(?,��=8j�����!�	��:�E�>�O>�I=�k>��W����ED�j1?>�GM>��N=kѽ�5��k'�;]F�<�#>6�>��ڿ�OP��徠L��+��
�Ȝ��/�T�|���?J�QJ������v��f��r��8��X�w����n���?�c�?"�z�#����蚿w�{�;���3C�>�w�($�ᇡ�q�ɽ�������]��M�SAj���`�+?�d��뭴��b���Z���?H�?�D�?ǁX�5;
�f�x�,�L�l�i<��Ӿ� ����ݿ�]@�Luf?'#?,Ͼ0=O�>`K
>�}�> { ?G�����ʾBsL>��?(|?Q�(?�2">�׿�ֿ�hM>�@�
@|A?��(�M�쾝IV=w��>Ŕ	?i�?>�R1��>��찾O�>h9�?���?�:N=��W���	�ʃe?N�<E�F�)�ݻ���=;�=�=���\�J>Q`�>�d�ngA�C-ܽ��4>�>#�׵�Jx^����<c]>/�ս��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�����ſ�u=�Б8���G�&��������K{�ļӽ����+������`�f�>�.�>���>�s�=*dE>+�`?w�m?+��>S�>�T��ɨ���վ�3>ٸ���(7��{:�J��A5���׾�a��9�����p',�����8;�
58��CQ�3N��c= �x�[��-H�1e=?S�>[ӾfvU���P��/Ⱦh`�����<*��۵־އ-�vt��Ξ?��A?�x�-�E�%��s<a�׽i�f?>����� ��hоt�3=Ò�Q�M;�v�>��H=�����-�j�D�2v6?��?�n¾����St�=����c=��?���>{��=kS>j�W?*�b�����P٩>,>�!�>��>�j���8���y��5G0?7jl?��D����d�><���;���U�}=y>�xܽ�m^�s&l>�=ZŒ�b�ӽ.Ż�>e W?���>`�)����`���9���==i�x?ג?E@�>e�k?��B?`�<�m����S���� w=��W?�+i?ش>ª��n�ϾHx����5?��e?��N>�Th�E�龏�.��R�x0?j�n?�b?6F��q}��������i6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������(*�= tR�h>�?q�?����d&= 	 �}/z�2F��[M��#D�=N:=P�����	���I��+;@��H-�5�=��>#K@L�O��m�>Q�1=D�ȿ5�ʿ�W��O ����O?�I5>|�Z��~���op���O��[C�xY�
[̽�L�>�>�����鑾��{��k;�𯟼_�>�v�[��>��S��;��嘟��84<��>Z��>���>S`��M����?�b��Q>ο���՟��X?�e�?k�?�o?cs<<��v���{�T���6G?�s?Z?a�$��"]���8���m?�1־��5���A��n��'�>
щ?	�>=5O�e">'�>!KK>��>�e����Ŀ>�Ͽ��,�'��?��?҉徻�?P�?l�Q?և
�d.ÿ!ߠ�;TG��>�q=?��=^��H`�8G�k��i�?�)?�bO�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?#�>��?1o�=0a�>
b�=��O�,�Jk#>�%�=�>���?O�M?~K�>4R�=�8�3/�[F�FGR�9#���C���>�a?��L?�Kb>���c2�/!�jͽ�i1��S�R@�G�,���߽�(5>��=>`>%�D�Ӿ��?Kp�6�ؿ�i��,p'��54?9��>�?��e�t�����;_?Pz�>�6� ,���%���B�`��?�G�?9�?��׾�R̼�>;�>�I�>-�Խ����L�����7>2�B?Y��D��t�o�q�>���?	�@�ծ?ei��	?���P��Va~����7�e��=��7?�0�!�z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?pQo���i�B>��?"������L��f?�
@u@a�^?*�$޿��	��j򾎼>2l�=I�9>����k�4�%]�ϪܼwO�=���=u�>WH>9�>���>ޜy>A>�+��?�&�>2��O���.�B��������J����2�����s �D�f�c���1P�.��\։=<w'=�n9�s����=-�U?7
R?`p?K� ?t3{�K� >]�����=�x#�Q�=�>�>�{2?��L?��*?�R�=UQ�d��X��S5���[�����>*xI>���>~��>麮>9��'�I>�Y?>���>z; >�X+=���=J�M>���>P��>�>m>kG\<����D��1b��A�KR�T�?Ⱥ���WL�;���nԾȾ���;�\%?�2x=С����������ѯ\?������X�M�<�WS?9D?l�O>.꾿vw��D'>�'�(6��倁=
GR��;��m�j&2>�U?�f> u>�3��f8���P�<���)V|>�56?鶾|C9�+�u���H��_ݾi@M>bǾ>��C�ii�}�����Cai�G�{=#t:?�?"2���۰���u�7���NR>4\>�==B�=NUM>nQc��ƽ�H�..=X��=��^>�D�>��/>�o=�5�>�	��|�Z�^�>u�=>��'>@�J?-�,?�n�5���x菾��M���c>���>�R~>�$><M�c��=���>�c>s_2��Vc�H��.�4����>y����J��:�v=����0��=\a�=M����M��,=%�~?~���㈿D뾭j���mD?�,?9�=#QF<�"������H����?A�@1l�? �	�:�V���?3A�?�	�����=N}�>=ث>ξ��L�4�?5ƽGŢ�r�	��'#��R�?�?��/��ʋ�'l�r9>�_%?\�Ӿ��>Ҧ�hU������u�?'=	��>mDH?����TWO�>�W\
?5�?�/򾲢��.ɿ�v�R�>�?�?��m�-����?�b�>��?��Y?4�h>D۾�Z����>�@?�4R?�]�>me���'�T
?��?���?8IB>���?�Ћ?��?�H\�$����G��P��� w�h��*m�>`Ͼ�M�O�M$���y����:�[���M�rL�>фh=�O�>�Dv<�����v�Φ�c!�����<��p>�M�>���=���=mܢ>�#�>�>L��;L(ѽ[#��'��%�N?���?����i��-�#~�;�`��?%�3?�݌=����>�(Z?!�v?ٲg?���>�L�鑿�XÿAת�N�0���=��>��>�(����>�7ؾs�@����>�b`>�1=*��)����/]����>�\4?��>��1>�� ?�#?i�j>t#�>�^E�k8����E���>��>kO?��~?M�?�Ϲ�	\3�	���䡿ސ[��6N>n�x?2R?X>$��������D��I�����~��?{g?��彯?�5�?��??-�A?�(f>��_ؾ����6�>��!?I�ӷA��K&����t?�J?#��>��x�ս��׼��k��"�?&,\?�D&?��'a�þM,�<s#�\k_�q��;�;D���>_�>����x�=�>�Ѱ=t*m�8,6�E�e<�E�=���>�`�=�7�_@��0=,?��G�~ۃ���=��r�?xD���>�IL>����^?hl=��{�����x��	U� �?���?Zk�?^��@�h��$=?�?S	?m"�>�J���}޾5�ྺPw�~x��w�^�>���>�l���K���ڙ���F��]�Ž�)�t��>G��>Q; ?B��>I�>���>����=�J@��񐻾ٖc�W�{�?�j�5�Ku�b���/�q�$=@վ�\�r��y�>,9��ƽ>p�?��<>�t>A?19R��љ>���>j|{>���>��X>�3�>Ő>x���9��KR?�����'�}��{���x3B?�qd?<1�>xi�������h�?���?Ss�?�<v>h��,+��n?�>�>B��,q
?�T:=�7�8�<<V������2����B��>!D׽� :��M��nf�Oj
?�/?����̾�;׽͇�����=�#�?�0?`$�N�H���k�pm^�`O�)ʽdrN���I0���t��'�������;���M0�K�=է&?ac�?3 �ʤ����c�b�w�A�#Q>+��>j͘>���>�x)>���l�8� �`�h+��������>Uz?���>auB?a�:?�g?�Z?}m���C?A����P?!>���;]�H?��d?�O?�)S?��3?�[?��>�?����¾�L���Y�>�}?-4?L�?�~�>z⫾�A>P��=Pͱ�p����x�:��>f����z��р>4}�=eɄ>BW?���)�8������k>�7?��>���>���$��Sc�<	�>��
?�B�>� ��{r�Ab�]U�>Y��?����=N�)>L��=Ym��i�Ѻ<R�=������=�q���i;��B <��=�=Ut�8a_�dD�:W��;�k�<�t�>1�?���>�C�>�@��1� �S���e�=�Y>�S>�>�Eپ�}���$��{�g��]y>�w�?�z�?Ҽf=��=Ȗ�=�|��wU�����7���-��<�?XJ#?XT?Z��?��=?Vj#?�>+�]M���^�������?}",?y��>�����ʾa�{�3�n�?�[?�>a�׳��9)�=�¾��Խ��>C]/�4~����VD�7�����넙����?Ͽ�?ONA�#�6�Li�L���*T���C?"�>�U�>�"�>N�)���g�"��<;>��>R?�7�>��O?O#{?��[?�oU>vo8�/��jٙ��S��">2x??���?=��?:y?x|�>�9>��'���߾�O���]�'E�7��T=Z>�Ӓ>\C�>8�>���=�=Ƚ�4��S�?��.�=�b>�y�>�O�>��>��w>���<�H?�8�>﮿�=��"����!@>�$u?9]�?,?ۦ�<�3��-D�tT��ə�>�c�?���?@9)?fFZ���=�߼4N����o��?�>��>�K�>��=\�>=�>@��>���>/b������8�w�@��?QF?���=Ԯ��򮂿#[žK��J8�E�׾�ܠ��m/>����"�F=��M��.������A�w��b��,�C曾�hܾ�����R
?#�D=���=���=ڃ�<X�今�@�6�>�:s=�����ӽ�Sv�K��=�V���,�WO.�CK�=�d^�5�˾<�}?v<I?	�+?��C?�y>n->� 4�Γ�>@���g>?pV>�P�`����;������$��X�ؾ�j׾�c� Ɵ�)U>+fI�H�>K*3>�8�=H!�<!�=�5s='َ=I3T�^�=^*�=O�=�h�=-��=�>)K>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�96>e�>9�R�ww1��P]�w/d�V�Z���!?n�:�Y%˾gN�>�u�=�r޾�\ƾw4=��7>��c=4-�/\����=�8|��;=-us=�:�>=gC>s��=}��M��=�HH=���=�&O>�a���I3���/�S30=.�=B�c>zN%>d5�>2�?Es/?xj?���>gcg��ɾ�Ѿ>è>�	>2d�>&Հ=Bm>���>)�6?nC?��U?+��>+|E=���>�Ŝ>�Q/���j��R۾r͖�{����?���?e��>����\�uy�}n2�������	?�],?��?�;�>+���߿�pn�Z;V������퀽�(�F��~�C������ �CT�a�6=��3>�@�>�r�>�I�>���=N8>W=�>3>�I>�,�=E�g��>�A�B�4�>z��=8�<.Tx���K���f������a<XE���A��Xd�DO��/�=���>@�> z�>���=f���~/>����آL�X��=Ǘ��^*B��d� L~��/�܁6��4B>a$X>`Ȃ�e ��A�?%XZ>�x?>tq�?�!u?�>���n�Ծ�P��Y�d��Q����=%�>��<�2;��(`���M��[Ҿ�;�>˪y>� �>�~�=#B<��7M��ku>f���\LH��R6?��$��^R�&�>_P�Ө�e'����h�Aj>��_?q����S>(�?V�)?��?��>r�Y�ꇾw
�>?��fJt>;�Y6/�d[����?-h??�B�ަ1�WH̾Q���ݷ>�@I��O�n�U�0�W���ͷ�Ԓ�>����e�о�#3��g�������B� Nr�V��>g�O?��?9b��W���TO����%���p?J|g?-�>�J?BA?�$���x��s���x�=�n?���?�<�?_>�>^B��K�>�<?P�?G��?7f?A�����>��>��_>����eM>��>a��=z>L$? �?�\?�\~����3�vx��t��I�=�c>�'�>\_P>�	�>ʩ<>5�=�����<(6�>��>���=Ղ>�X;>ڦ�R=��x+?Fa�=�:A>�?�٥>�ii=�>���<�&>���#c�K���"���(|�����.!u<mT>*s�>qVſdS�?�G�>��K2/?㉰����P�>�$��<冾�F�>I�����>E�>2k�>��s>��I>�7��[9Ѿg}>'���X"��QC�G]P�J�Ҿ;��>�h����*���
��� ��9M�Ƹ��[�gni�E��~�=�N�<�]�?����k� �*����TE?���>RU4?k���[��,?>qN�>���>!!������쏎�\l���?���?[;c>b�>#�W?��?Ӑ1��3��uZ�p�u�o(A��e�G�`��፿	���v�
�)	��>�_?0�x?�wA?wM�<,:z>��?C�%�'ӏ��)�>|/��&;�??<=.*�>�'��a�`�=�Ӿ{�þu5��IF>�o?�$�?\Y?kVV�߁Q�� >��6?p�/?��u?��4?2w<?�^�4�$?�50>�.?)�
?�5?R(/?�"?��<>�c�=����$=�e���	��A�Ͻ2�̽NB��8@=r�z=0�|�ʰ�;�
=+��<	�޼*���$9G8dA����<Yf7=0��=���=�H�>��Q?���>j<�>ߗW?L=/��1��۾��^?&0>�r���[��������D>o]?��?�d?&>�3���.�6go=m��=Kw>F>�>��>�]I=����՚<��v>���=�M�=pT�;踐�������~>3�s>'��>�0|>'��ȷ'>�|��N1z�;�d>,�Q�-̺�Q�S���G�y�1�G�v��Y�>G�K?��?О�=1_�X.��PIf�(0)?�]<?�NM?��?��=x�۾��9���J��>���>	Z�<��������#����:�l^�:��s>�1���h���'U>8��+���k�I�I���辩�g=R�
�<�6=��8�ҾFx��W��=��>�D��<� �Mz��۩�K?��^=����e\�P�I�>y��>S&�>{�*�M����C�Ö��܎=��>V+>A�м
��c�D��� ��2�>��@??�E?U�?�f��:+~�)����e~��"�>�N,?"v>0�?��=+(<>A��7@��[�ǡL���>���>	�-���'���4��1�7��hճ>�01?�b�ݷ?|�s?[��>� �?Χ2?s��>��?{��4����V9?#�|?Qg7��غ�:㾸�K�P�<� �@?�?t�n��>׍�>=�?��c?Qt?r�?F�>J�-��l���>��>]�H��������>I�8?�@�>�cy?`<h?-�u>�_?��[���{�=��<� �>�ч?�-?��?�˙>�,�>�n��9a�Y�>���?�2�?S�a?�"4>G�"?/\K=�0
?DS>?h��>�C?�DX?���?�N?ø�>'�=w���v�����;�Q<i���R�?=�B�=�V��<K�衜;�׆��~%��4Խ_5Ľ�>��ݽdm�<B:�����>q>*����/>�ƾ_܋��H>��ϼh*��H㋾X:��m�=�~>��?�ԑ>�b'��Q�="�>��>�-�Uo(?�Q?�l?㜫;b��ݾ�M�Ze�>/�B?R�=J�l��8��T�v�kyl=�dn?�]?�[�ã��r�b?�]?Q��<�\2ľ�/c���龤�O?�
?"H�L(�>r�~?��q?I��>!xe�`#n������Kb��Vk�?�=�u�>O\��e�Y-�>��7?^�>�c>F5�=�۾~�w������?���?��?X �?�?*>��n��*࿷ ޾�A��_�n?
�>�����S?�=l��m�"���!ܾ�()�l/��+z��[a��}^� I:���f�B�>��
?�L�?	�Y?�ہ?�)���:�ux%�恿F{b�#��FH�|8>��cS�lI�8�l���!��I}��h�>=�~�Z�A�~i�?p�'?0�3��k�>U���𾃶ɾ$D><l�����!ՙ=���4�:=>�R=[�f�S�*�y���?Ƃ�>���>b�=?��[��J<��.��l8�����D,>���>�֓>t�>�� ;n,��T��ƾ�⇾ѯӽ,m]>1��?��l?�x?�Y¼l��J��z#��ǹ�Oٿ��D�>����k���e�Cjc��X��D�w�d�m��.�s�5��̽e9?�@>��>�
�?��?���K*K���]���s��>L�1>јv?��?�s�=��=��/����>�l?���>/�>򞌾�F!���{�&G˽���>�֭>R��> �o>�-�/\�]i���~���9��I�=p�h?oy����`��م>Z�Q?���:;%E<�l�>�Fv�w�!�@��I�'�:�>�t?Fv�=K�;>�kžr���{��9��\�.?o?����%'��m>g�?���>1>�>x?�ݩ>z=����i=�?JMX?7�P?fQ?+� ?��W=d2'�W,ӽ�����=�҅>Ӊ> �K=��=7R� ��`�8�U�b=l?$>�i�~�ֽ�����������8�=m�>�pۿo�K��k۾���@�f�
�ĺ���K�� n����	�p|��c�����x���� o$�(�T��[c�4���]n��-�?�a�?d���QF��n��d��t���[��>��n��3��\��y���[��/\޾�쭾-z!�J=P��h��Md�g
?����%���)�����H�U?=?�@j?WF3�6�:�#ၿC�!>�>�.�=l�!��m��T�пWMҽ)�j?�E�>O���p;\g�>��>�z�>}�?,�待s	�kb>7�/?�?�?�k���į��3ƿ����?�c@e}A?��(����#�U=���>��	?O�?>�&1��J������X�>?�?��?��M=�W�����e?�<��F���޻�&�=�=7q=-��_�J>^�>����KA���ܽ;�4>�>�U"�r���\^�qV�<�x]>�ֽ����5Մ?+{\��f���/��T��U>��T? +�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=|6� ���z���&V����=[��>b�>Â,������O��I��U��=�����ÿF�K��$(����<� ���S���
���g=-��;?	��C��-����<V�>�ƀ>�	�>��
>�D�=;;Z?'�s?|~�>�~}=^l�_�D�j�Ѿ������x���9�:���=�:������|������Lk
�*E̾�N�:�����e�����Y�
�5�Y���B�r�7?�R�>~E侢�i�/8�=�ܾ��0��0��늽Io޾�/���]�rϟ?�%?�\��9U��9	���=��m�k�n?�Nͽ�}�E��NZ>.���r�=��=��4��b�O���Bp:?�z+?WY��hȇ�!$N>h���F��=;?�Z�>��<	��>�K?t��<��U<�f�>���>��>�d�>i���פ��{��2�>�]a?�um=k�|�/�>b/�_����潊?
>+ܐ<�NQ<�Zd>���=����d���y ��=�(W?���>�)����]��$#��O==Z�x?ڎ?-�>�zk?��B?c!�<�b���S�����w=��W?�#i?��>����оFy����5?��e?R�N>:ih� ��k�.��S��%??�n?_?�@��hv}��������m6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?r�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=9!��ۭ?Kt�?&s޾��=����'v��z྽5��6��9#c���E#�|-��<��XϾ�;�[��jL=�O�>��@�ԗ��0�>�d���)���̿n�t����3p�]?��>��{�
?���Ej���a�O�W�=�7�9�`����>tU>�����h��|�,�;��	���>޳�%��>acR�Eᵾ郟�p�H<�%�>�o�>��>ҥ��;C����?�	��)οa�����O�X?$�?:��?��?��<�v���{�����bG?`�s?)*Z?it#�;�]�|
;�%_?�پ2�-�>�C�S�N�k�=���?��E>?f ��$Z�(#��I�>L�>qVX�S.Ŀ�2Ŀ���ܾ?p��?�w��O�>!��?�%e?�`1�e:��,tG��iB���>h?D��>�>�&7� �3�=Y��)?$ ?i@l�G`'�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?Y%�>��?7k�=b�>�i�=u�� -�Am#>��=I?��?#�M?&M�>�^�=��8��/�IYF�iGR��$���C�F�>D�a?ۃL? Mb>2��&2��!�>nͽPh1�B鼊V@��,���߽q%5>?�=>P>G�D��Ӿ�?Rr���ؿ	m���m'��=4?�ԃ>��?���Էt�=��8_?x�>�&�i+���)��Qs���?�H�?��?P�׾��˼/>6֭>1'�>3dԽ����n����7>��B?�� ;����o���>7��?$�@>ծ?g�h�[	?�$�[I��s[~�`��Y�6��z�=�7?3�� {>���>�/�=,iv����ȿs����>�<�?�{�?���>�l?��o��B���2=�8�>�k?Sq?��w����B>G�?�������C��$f? �
@v@�^?�4�ݿSC���U��O0ȾS�>}yg�̏�=�y�!_�>jɩ>E�x�T�m>�ۙ>O�N>=�>d��>�'>�D�=i����%������8��<,F�p)+�$/.��[���=�a��Vv��qܾxG۾,�9WI��6�=ﮄ�/��w��.��=�V?�P?e�o?23?Ȇ�SU">y���=�A/�e�=���>�%4?#DL?4�+?�ܬ=�ޒ��|c�J ���/��	���x�>N>���>��>��>�ڻY�P>oU>>¦{>8��=^�<=����V�<��L>���>��>k(�>��=7!�<�p���E���N��QA�EM��?�Y�HY�1*���|&���оԽ%>�?;W�=�+���ſ���&	X?�oj�ߢپ��L�E%�=� B?8TI?�!5>��ɾ���$+=��������2=�v��n��zv&���0>3?ֻf>�u>��3��f8���P��z��md|>p56?%涾�J9���u�-�H��cݾLM>J¾>�D�/l�$��� ��ki���{=px:?��?y7���ݰ��u�A��]KR>:6\>O8=mh�=;\M>�oc�M�ƽ�H�sU.=���=��^>�V?e�+>$p�=�d�>�M���[P��٨>C>�f,>`�??�$%?�y
��약�#����,�ex>L��>�[�>��>�)J��4�=-D�>�b>����ށ�$��(A�l|V>�	��Z�_��:n�p�w=0���}��=�6�=f �o=��Z$=��~?���䈿��ve��mD?�+?� �=*tF<��"�3 ���G���?_�@�l�?�	���V���?A�?
��5��=�|�>�׫>nξƗL�V�? ƽ�Ţ���	��'#�1S�?��?f�/�:ʋ��l��9>_%?��Ӿ�w�>���I��b,���u�Lp)=M��>�H?'���@�P�0�>�`
?M�?���#����ɿ8�v��h�>�
�?Hߔ?�m�����?��>�h�?3�Y?�h>uN۾��Y�j�>��@?R?*��>�(��(��?g�?Ʌ?�.V>R�?��?��(?���iʾ�Ě�΀����H�k>��>UB=9�l��"l�iO���_�+�S�g�!�&�>H_�<���>�	ͽ�pľ���>�ݽg��.4��5x->>\�>ֿ>����A�>�۹>�>r��=	�=��l���l4L??Ⱦ�*�l����<q��=�^��o?|�2?�\I��;�+�>��\?H��?��[?S��>=������������J,�<�
L>I��>�U�>?䆽�J>��վO�A�>�>�>��t��nؾO���p����ӛ>�]!?�X�>H�=�� ?��#?�j>�(�><aE��9��6�E�<��>S��>�H?��~?��?�Թ��Z3�����桿��[��;N>��x?�U?oʕ>B���ރ��jE��AI�����V��?{tg?�R�<?"2�?��??[�A?�)f>����ؾ�����>��!?���A��L&�C�u{?1O?
��>�5��'�ս�ּ���x����?*\?�C&?����)a��þ�)�<��"�I�U��j�;��C�,�>��>x������=�	>c԰=rCm�D6��f<"a�=q|�>��=�)7��l��0=,?��G�}ۃ���=��r�?xD���>�IL>����^?il=��{�����x��	U� �? ��?Zk�?h��?�h��$=?�?S	?n"�>�J���}޾7���Pw�~x��w�\�>���>*�l���K���ڙ���F��a�ŽG�C�W��>ԭ�>���>��>�`$>s`�>o����%������޾J���29N��1>�d+��Jվ�)m<�'c=�5��1]��1�>��I��u�>]�?��=���>u�>��=x��>2�Z>�ö>���>��w>� >�(q=}!�=U}��@R?l��C�'��辎
���A?l�d?�|�>*�j�)�������Y?u[�?d�?�(t>Y�h��8+�u�?E �>,���u
?VT;=�����<%ҷ�h	��و���#��>0ֽ{:�K�L� g��;
?#>?F����̾��ؽ!#�����=�z�?��/?�(/�&�D��n�1l[�P<K�4h�_x��J��r�.��u�����V��	��2�$�ԁ�=h'?H��?�W����޾>��� p��@�NSd>��>:�>d��>��V>7���8/��]�N!�/V����>�Hs?Ǜ�>Ĵ_?�(*?P\P?�:Z?1�=���>���~��>��[����>X6?�`?]9+?�zC?��7?K�W?�B=wS��߾g,��Q+??R� ?h|�>���>S��}5�=��x=.����g�%8�=>�^<�cB�i.%����<Şy=��>�R?���}�8�&���w�j>�7?��>���>s��8�����<_��>˲
?[9�> �?�r��h��h�>O��?���6=�)>���=?#����κ�C�=1���$�=����0;��!<}��=��=��r�������:��;YC�<�t�>,�?���>�C�>�@��� �K���e�=2Y>�S>_>XFپ�}���$����g��\y>�w�?�z�?��f=5�=z��=�|���U������������<�?6J#?!XT?Q��?j�=?gj#?��>�*�PM���^��k����?r!,?d��>��3�ʾ��w�3�U�?([?�<a�����;)�m�¾��Խ޲>\/��/~����`D��������}�����?鿝?�A���6�2x�����#[��U�C?6"�>�X�>y�>	�)�C�g�)%�3;>Ί�>6R?'3�>Q P?H1{?�[?��T>u�8��������K<��">�@?.��?�܎?7�x?M��>�l>[)���kc���d�*��؂��QX=�Z>zb�>L"�>�>��=�Ƚmj���h?�I��=�1b>3��>b��>��>��w>��<��L?�S�>��¾/��,��(���}yq�8B�?��?g�1?g�=�
�#�)�j�;��>4*�?��?t??>"��\�=�c���ߐ�߱���.�>���>S�>�U<f��<�>>��>�H�>'s�����o=�����:�?��T?N6�=Z�ʿVro��Wɾ��¾�hB=�9��ƞ�n9Ľ��� �==V엾9u+�'���g�+���q��^�R:��?Jƾj��)�?ꚉ=X4�=J��;�a�<�e��*7�=�>X#=�΁�����=�i�2!B="���(E��qĽ7�=�i=(�˾ӏ}?!<I?-�+?��C?�y>8>��3�Ř�>����G@?fV>3�P�����ǉ;�����v!�� �ؾv׾h�c�[ȟ�QH>AfI���>�63>NE�=�P�<q�=s=9Ǝ=��R�n=�#�=^Q�=.g�=���=��>nS>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>=> �	>-iQ�m�0��gX���g�nZ��C"?M;� .ʾ5��>k��=PEھ?þ�JP=�x?>��=�Q�Da]���=u�-�+=���=Dh�>��B>W�=�һ�	��=l2=�l�=�V>��7���)�O��.=ƣ�=F]>��&>��>L�?�0?�Fd?�ػ>��m�c̾����J$�>���=H�>�ń=G�J>�Ҹ>��7??]E?�vL?��>�:�=Ś�>%V�>Ή+���l�E��a��#�<S��?뻆?0|�>� �;��K�����L=�qX���^?�1?N�?��>����ؿ��J�X3� 7@�ݘ꽗���
�����k=e�p=[SE�
�6����=B��>K��>��>ሇ>+j�=��;=K��>(X>���<��H<nD�<��3=	^Ƽҹ=�f��/��׆%=1�V<2��VK ��:��	��f�T������L�=Ϥ�>�.>@N�>��{=�|���4>׏��t~L��d�=&���S�I��i_�0��><3���Q�.�!>�+n>��G����R?�5>=j>��?�fy?��=���Ҿ/ė���Y�ֽg���=w��=!�$�A�7�=�[�GJC���ϾN��>�Z>_��>6pL>@�4���Q��/q>���Y$��y�>AӀ�� �j3���_��ݩ��ĝ���k��n�=9=J?/���y>�#=?�~3?E]�?��>���Y���/==.����<S�'�j�;�>���
%?�#?V�>�@侩{[�HH̾!����ȷ>�VI�u�O������0��T��Ʒ����>8䪾Ѿ�3��h��������B�r�r�3%�>ĴO?iݮ?�nb��E���LO���[S��H?�}g?�8�>�H?kA?(���T�`����=8�n?��?�2�?:�
>^�=� ����>)f?�e�?�U�?�Fq?<5���>\���$>dw���4>(�>/0�=l=>�?�
?%�
?5H����
�6����B��=�H��+M=�ّ=?��>���>w}>�p�=Q�=5��=.�]>�>A�>�M>k�>z�>M���N��c$?���<ۼi=��+?'=E��=��>c	�>�=T�*�b��bZ����d,�К	�NZ�>f6�=Qm�>��ɿ5�?U�>r�$��q3?���[�0��`�>(18=H��}E7?ʿ��ڥ>��
?TH�>+��>b
�=��<s׾6�=L���t'���=���L�?MӾJ؋>�A��q�?�`���ؽ �S�c[����d�������=�"Q/<iH�?����`�\*�X�?��>�v4?�Z������{��=>:�>�ڑ>�0��I������D�3��?&Q�?�;c>�>y�W?R�?N�1��3�vZ�;�u�`(A��e��`�j፿'���B�
������_?��x?�xA?�W�<�9z>B��?��%�ӏ�(*�>�/� ';��A<=�*�>�)��8�`�U�Ӿ_�þT8�.IF>_�o?�$�?jY?nTV�ci6�j�6>SN;?L2?,pv?k�.?r�;?:S��$?@�.>��?N�
?�9?H�,?�?�I>޷>���%H�<P�������J���hս}�!��w#=p�s=T�u<���<'�@=�n�����[Լz��;ro��@��<<=Ʉ�=�^�=���>��]?	�>�P�>).5?� +���6�� ��D�)?��K=��t�@fx�Ø������>"�m?�ɫ?`X?tB>��A��>���>�!�>h�8>��V>�~�>P8
��T�BO=s�>�x+>��=Ip9��Vw�,�
�����2��<�>���>3|>���}�'>|��x3z�A�d>D�Q�e˺���S�]�G�d�1���v�Z�>��K?��?*��=^�5���Hf��/)?�]<?,NM?��?��=N�۾��9���J�l?���>Av�< ������p#����:�M�:��s>(2���1��p7>�C�����i�s�K��H��6��=2����=�G�,�޾�vp���=��>�������9�������K?��5=wD���[��ߵ��O(>L|�>�t�>$���u>���D�&���nfq=���>6�?>ā��('��d?�E�W��>�&?�QR?Q��?�)򾳩L��v!���׾��j�N�=(�D?��=V�>��>k�->h�����׾�9��J���?��>���I��x����.���/��>ȋ$?(ظ>�|?z̈?��?7M�?��u?I7�>���>�]��֓�;@?�Dl?�r�"���d��`�6�Eh:�õ�>�A1?,m��d�>�I"?S($?� K?�ci?��?�!t>�Ӹ�~�b�Iz�>��[>�2|�W?¿m�>��3?
��>ڧV?g@W?=h7=2fR�#�g�����$��|�=�m?m?�c?h�Y> ?����6ku<�E�>B�?�aj?Ɋ?�|�<X9?w߭>��?�r^>O_#?�H#?�&?��h?L��?��4?(�?�+<������2�������
�=���<s�i=�m��B���f��T0=%�)>����!��.X=�A�^����3>�h�>��s>(��c�0>�ľ�[����@>�E��UK���͊�
�:�b�=���>v ?S��>	?#��ϒ=��>E;�>u���4(?��?�?°);#�b���ھi�K�c�>FB?���=��l�<�����u�x�g=��m?��^?G�W�W����b?d�]?Xf��=���þQ�b��龤�O?r�
?��G�t�>��~?[�q?A��>��e�r9n�(���Bb�C�j��ض=vr�>�Y�W�d� =�>Ǜ7?JM�>��b>t+�=Yw۾r�w��l��A?,�?�?���?�.*>:�n��3�{� �ݳ���^?�?�d����V?�>`5辿��n������L����پ�Ⱦq<��dZ7�g���}\�0��=�?�d�?z�u?��w?s��F�H�[�X���t'�޾�; �D�h�c'��rZD��_p��D!��&�O5��LG�>��~�ן@���?�(?K2����>�B��$7�ޣ̾�n?>���>�S��=hy���==,-O=Лg���.�����J  ?HR�>IQ�>�<?�u\���>���1�'g6������;>��>�$�>��>�h<��!�_���rɾ栄���ս�h\>��h?�V?�\g?�WG�1���u���4���l�۾ʲ'>lz�=q�=�c˾E����A/��&1��
c��~Ѿsu��K��V��R�2?e�e>�>O^�?UO?s�"�ͧ�Ȇ��i;�e(�>�M�>I�`?�2�>��>�;����C�؅�>��p?M1�>\{�>�䐾����V����7�>s��>J-�>�h`>�%n�h�e��뒿E	����6�%S�=�"n?�Pr�:�i�c2Z>�aL?}��
��=p�>�r���)��F�}6K�]e�=��?;T�={pT>Va�����xk�ԙ�e�M?�$�>ԫ����{�>�N>��>!�>~gl?'�?��پ���>��#?�`m?p`P?@�X?u�	?�Z�>���昄�P�-�%Km=���>�G�>Gy0=��=Y�Y���;��3#�<�>��>����Y߼��$�=����K#��t���>v�ۿg�L�Jh߾���x��K�
��6���Ȭ�,������t���5�����q�'�� !��<Q�Of_��ϐ��p����?0�?-_��	��?_��+��y��J�>�5h�+1T�����Q��󯖾��ھ����s�#�YmM���f��e��?��Ѿ.���N�����?zo	?@�?k�4��1��@��7>ջ��m�;�hƾ;���aܿ��k��D?	��>�-���%>3��>O�<���=bA�>�o��oܾ��~=�A5?3*?��>ߞ��(�ȿe:ǿ��t����?�$@��A?�(����`�R=Y��>�#	?Ƴ?>L�0����N�����>�G�?p��?ɈP=�rW����8�e?- <*G�&ڻz��=K�=��=�+���I>�s�>$���6A��ڽ��3>O�>��!����.�^�}��<��]>սO唽5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�}��=[��>c�>,������O��I��U��=i��xGƿw�?�6Y3�=�<�U����2����uM���=%ۥ�J�����]��j8=�W�=.zq>��>/%�==>�0W?[mQ?Ϡ�>��>�)��˺������ܥ=��<��캼�w��e^�������Tľ/�%��������{�྅�K�����)�h�P�������~W���_��fD?5�>���A�e��ǽ������v�ё�<e����Ͼg�2���m�{��?B�?�q��I��r��_��=�����d?��0�H$���a>�R�j���Ԓ>Ǧ�=9�De��OE��OE?��?��ʾ_'����`>;��#x+=K9!?J��>?
>��>>K?^{�齺��4�>�b�>-��>hB?.�x��j���d�50?��`?���<��[��w�>��ܾ��l�j�V<�H>M�:����o��=�{;=����r�Һ�烽Qb�=H+W?i��>�)����Y��C��>d==گx?`�?�:�>}tk?��B?�_�<�W����S�a�7�w=��W?" i?c�>p��"оt����5?Q�e?E�N>�gh������.�O�X"?��n?�Z?sG���s}�������Jo6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?j�;<��U��=�;?l\�>��O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������R^�=F3��il�?H1�?�`ľ���=҅�ȴt��Ѿ>S��k�=W����q-����}9�A-ھL+
�B|���=]��>�@��v��)�>�/#�v�ݿ��пف�w྄�$��$?��>}�6�6��۝���H|��<���6��.F��>f>�*���t��?|���;�<%�����>$y��N�>u�Q�����G����M< c�>�^�>�ӆ>�G���^�����?���X>ο�������+�X?�<�?�l�?mr?�;*<�!w���y�,���G?֏s?�CZ?��!���\�]�:��b?eڴ���R�S6�?4N�	N.>�$.?'y�>z}=��^9=��>9�>�ұ=�.��¿�ܹ�����n�?
v�?�Dﾈ��>풠?��7?�z�|������K<<�<ǉ<��C?�>P����j�lE�_=��n��>"�7?�b����]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?a$�>��?�n�=�a�>Ed�=W��-��k#>�"�=��>��?��M?L�>kW�=��8��/�;[F��GR�Z$�>�C��>��a?�L?�Kb>����2��!��uͽ�c1�P鼵W@�j�,�՞߽>(5>��=>�>^�D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?kQo���i�B>��?"������L��f?�
@u@a�^?*[Qſ�d��5���Ǖ��nU>�0>�Ӧ>�_��^t�F�=�ݽ��X��|`>�S]>�R>g��>+�(>��=��>n�~�%J�pݼ��	��[�H�#���/� @b���:����T��ƾ�顾7%:�:Rν1L�+����j�l �g��=j�U?R?�p?Ï ?��x���>����3=/�#�z̈́=�.�>�h2?g�L?[�*?ԓ=[���W�d��_��V@���ʇ���>HrI>}�>�L�>%�>�I9��I>�.?>9��>'>�r'=�$�k_=��N>�N�>���>�w�>Rd=��s�,��:����8���w]ľ��?j���B�w������A����R�=�0?r�=͜���Ŀģ��iV?ݭ���쿾���}b=��&?s^a?�2�>j;��x�����5>���<eؾx��<YD�����qxk���C>��
?B�f>nu>\�3��c8���P��{���l|>?46?궾I9�ؿu���H�q_ݾ3IM>n¾>,CD��j�{���U��pi�,v{=�w:?4�?�0���۰��u��B��oSR>x7\>�`=)t�=<]M>�Kc���ƽ[H��u.=���=�^>2�?;,>h��=�^�>.���y�R��e�>Y�B>=�,>ld@?9�$?P��5���G��Ǽ+���x>���>�>n#>��I�TX�=�.�>�Vc>ȏ���^���h��y@���V>�0��U�]�@u��Uu=f����_�=�9�=� �4�<�2�*=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾOh�>{x��Z�������u�v�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?toi>�g۾=`Z����>һ@?�R?�>�9�}�'���?�޶?֯�?2K=N�?���?Q�>��Ѽu&����_����4�>�&v�τ�>ų!�%-G�8�t��󱿘B�=��C6�8�?�G�=�[�>��D�{��c�>�k�����������=P>_�*>;��>���>�5>?��=�K==��=��]��K?���?���1n�
��<ss�=��^�='?QH4?�Z�b�ϾAި>��\?w?�[?Fm�>����8�� 迿�y��ʒ�<�K>,�>'V�>�/���HK>]�Ծt;D�[t�>fƗ>�ģ��;ھ�1��ꃤ��G�>�c!?!��>�ή=]� ?'�#?��j>�(�>aE�e9����E�X��>ߡ�>7H?��~?Q�?tֹ�3[3�����桿_�[�X9N>�x?�U?�ɕ>J���p���r�E��4I��쒽5��?sg?�Z� ?�1�?3�??��A?+f>��xؾJ���Q�>��!?"��A�qM&�f��}?GQ?���>Y6���սj4ּ`��V|��p ?�(\?&B&?;��+a��¾�:�<�"�J�U�E��;�jD�{�>��>����"��=�>�հ=<Mm�@B6�8�f<e�=8��>��=0.7�r��1=,?��G�ۃ���=��r�@xD���>�IL>����^?nl=��{�����x��	U� �? ��?Zk�?r��?�h��$=?�?S	?p"�>�J���}޾6�྽Pw�~x��w�_�>���>�l���J���ٙ���F��[�ŽD��E��>��>��?�;�>A�>}�>5h��N�~�-�|����g��F�L���1�N2'�[����,�1=�<Z���]���$H=�*X�z|�>�3�>��>�w�>~_�>������>���;�>?��;?�|�>Á�>^ư>��t��k��LR?����(�'����Ĳ��-3B?�qd?U1�>i���������?���?Rs�?�=v>�~h��,+��n?8>�>1��Cq
?T:=�:��A�<V��E��E3����>��>pE׽� :��M��nf�Yj
?�/?��c�̾�;׽� ���_�=���?2?�.���-��}h��d�k]7��Cཔ?M��þͅA���w�$]��N�����|���+��L#>�"?`��?�x辡	��n����y���P�&W>�%�>w٪>.�>ׂ8>� ���*���t�U�)�ǝq�}��>�Kd?�.�>�3A?.�?�A[?#�m?�n�=Q�>%׾l�>��>-�>?O36?α$?J�M?�'!?�IC?�@�>H;�sH ��%����.?�� ?��?ϸ?�
?�����<"��u��=�2޾u��<`��=���RKw�$|<Bo�<��L>�?���^8�,���R]p>�l8?T$�>��>�y���z�7�<�>�N?���>eF���r�n����>5ׂ?s���<P&)>���=�4���w��A�="(Ӽ�~�=�D��g�9�<84�=ݕ=�7��ۅ9&[�;�D�;.޹<�t�>6�?���>�C�>�@��-� �b���e�=�Y>7S>>�Eپ�}���$��v�g��]y>�w�?�z�?ǻf=��=��=}���U�����H������<�?@J#?*XT?`��?z�=?^j#?޵>+�iM���^�������?lh#?#�H>���!{�k詿��'�B�?΀?ۢx���8�iz������H����=��1�[Ά��8��"�=�x
����c��?���?����
fD��⾲��������H?��>�0�>��>x:�:�y�f�-�PS>��?�Z?x(�>��O?o9{?c�[?�T>p�8�d,��&љ��2�{�!>�@?ٱ�?*�?�y??y�>��>+�)���EK��{����傾�V=aZ>���>a"�>��>���="ȽX~����>�CX�=:}b>���>��>2�>�w>�ү<�V?8c�>٥ྠ�dyžo�������)p?��?�-?A;D�Ѿ�������&��>Fé?���?,�<?}@���i�=+������W��E�?�9>Fҩ>��]=��0�$��>�IK>i�>����X�p|9���+=��?�R?M�4=��ɿ����Dо|ܾ��<OIƾ�2����=�ޑ�Q�c>�6��Ã��l��A��~�ހz��?����ܾ8���ϥ?]��<�>�v=~��<#�߼���ZvN>;�">�?�=/��q�ż�>��!��=I����p��<n��~��=jϠ�x�˾pQ}?e�H?=}+?��C?�y>@�>�00��>�>Ju���$?�U>gN�o8��1�;�0������}پ�׾�tc�g+��>�> H���>H�4>x��=�?�<K��=�Br=ŏ=l �m=`��=��=�&�=���=و>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/> <>>d�>��R�B�1�>`\���j��X�
�!?��9�$Ǿ��>�=�JھL���.�A=�A>>�?y=��J�]�J�=���SM=��v=g�>;�<>���=j~���C�=K+k=$(�=�ZX>�&�,1��2�`�6=��=��b>�Z$>��>�? �+?f6g?x��>��T��鯾_ܺ�d9�>�#�=6��>���= �j>�ý>4�:?�2L?��Q?hد>Zg�=u~�>�;�>|�-���t�ھ����_��{x�?k�|?g�>��d��s�ש�p�:���̽�p!?Q�2?��?��>�R�B��I0'�0/�䙽T%��� =:�p�S�c��G���#��p�=S��>��>��>�x>�&5>�L>'��>{�
>��<ڤ�=���:��<�o��g'�=|`|���<��ʼ6QI��j�k!�^���$���f2�;j�g<ߘ;9?�=ɿ�>g8>"��>�S�=&	��'/>Ή����L���=�`��?+B��-d��P~���.��C7��A>*�X>+����0��+�?�X>�?>i�?�6u?�� >x��4`վPN����d�}T��=�Q	>��;�A;�8�_�I'N��vҾ$̋>�&>ӷ>�V >0�2�>-F�0&�<�ھ��U�0��>������غ�}�Ձw�����婿���i@A>s�N?�ً��R{>�I?��P?P�?���>i<��e��9g�>p_{��%s��B:��s��� �͓(?�;(?,�A?(D�X2U��I̾R���޷>�?I�R�O����0�����η���>'�����о�$3��g��������B�UPr�[��>�O?H�?�5b��W���SO���� ���r?�}g?@�>�H?�@?�.��8v��o��Q��=a�n?��?E;�?>u>d�H���>�w?�M�?�#�?��k?^�P����>
��=�S)>؄�f�,>��L>I4�=˦>�?�?_�?�7��Sp�ي��<����b�B�=Y՗=r>�n�>�L>��=SRi= }�=Z�W>�*�>�v�>��>�W�>U�>׬پw7���?(�>ݓ~>&�G?��>֖	>�Fнc�E���5=��(q������˼�������yν��>��Ŀ%!�?z�}>�E�"�8?�>��t:A�7'�>ܠ>o�	�>��>T�W���=9k�>�o�>"H�=��>Ŷ��@Ӿ2W>;��dl!��)C��zR���Ѿ��z>̩��.&�æ��v���QI�Wg���a�j�L1���;=�hJ�<G�?j���!�k�-�)�-����?s�>w6?�쌾_����>a��>հ�>�B�����1ʍ�C����?��?=;c>$�>]�W?;�?X�1��3��uZ�:�u�y(A�Ue���`�፿���\�
� ����_?��x?�xA?1V�<�9z>$��?��%�-ӏ�*�>�/��&;��C<=�*�>�)��e�`��ӾM�þ7�IF>`�o?-%�?dY?�UV�~�����@>��8?t(7?C{?"+?��??��!�y4%?�F>DE?��
?�V9?��/?F|?xA>A�!>M�=A��<e�����o�Nǽ�VĽ�g��eZ�=�̂=��=�s�;D�<����a�V�>����f;���U�/=\A=�t3=X�>�ߩ>�R]?�^�>L��>�8?2!��6�~���a�.?M=�T���˃�9����H��	>�.l?6�?[?�`>A��gC�3Y>n��>�(>��[>ӱ>�0�U�B�8��=ʧ>�C>�i�=S#L�{�'��ȏ����<d!>��>�0|>���:�'>�{��3z�ݤd>7�Q��˺���S� �G���1��v�3Z�>a�K?�?�=�]龚0��If��/)?�]<?�NM?
�?+�=!�۾��9���J��>��>�P�<��������#���:���:�s>{1�������a>���G�޾Gyn��5J�x9�#I=����V=d��!�վq����=S>�
���� ��͖��Q���J?��_=�_��ogT�Mߺ�`�>#�>H�>��<���k��o?�6j��7��=J�>G>>�`������	G�����G�>��X?��@?Cȅ?Z�V�nm�ٸ2��꾊���(dֽ{M?���>5��>�Z�>#�.>ލ�U�����QO\����>6�>q���+N���˾v���H����\>i�>��4>���>�Q?�S(?6>P?|�?��?�!�>�!ͽ ���'�?�7�?(^�����Bz��P���ھ�!�>�v�>�(��Sx>��O?W�P?�O?��d?O#K?�C>��W�������z>z�v>m36��ꢿ�'�=�1?�M�>�B? Af?C!;>a<6�������Cp>D�>@e'?���>�?iI�>��>�������=���>��d?�ރ? �p?�|�=��?�j,>���>�Ζ=�;�>h4�>�0?��O?@s?��I?hV�>�c�<�+���f����l�ANv�^
�;�?<�#t=;M��j������<-J�;
�j�VS�����Q�E祿)�X<��>
{>������->vþp?����<>�i��n��l��}�*��`�=�
�>ͧ?�ϛ>�>%�D�x=���>C�>�q���'?��?�?��H<�Sc�)�׾�!d��K�>U�F?&+�=��i��ߒ�8zu�:`h=$?n?*%^?�ym�D��ɍg?�O?ˀ'��Z���籾)��
��L<�?j/�>��A�`�?���?g��?A�?kż�(��ߩ�O��2*�_Ղ=�\�>������j@:>�2?�'>�U{>�k�=�3���'�W(\�4�!?�	�?�E�?�҆?y�>�g�=ɿ���L��/x[?�H�>XK��>� ?i����Ѿ�����ё���pê��Э�$5��tԨ�\n&�����X�ѽ���=��?��u?��o?�]?� ���c��M^�tE|���U�����>�zE�x�E��F�/�p����'<������9m=�1V�O�,��?>�%?��H���	?���]\ �y�����n>hq��4����p��j]��������<����j�K!F���?��>�7g>�1g?3�W��� �j�H����ս�� >� ?�pe>�h?���=
E�dU%�͆��D����Y>Q_v>��c?�&K?��n?����&1�vf���^!�ä1����-�C>o>�a�>��U�����%�M�=�	ms���62����	��=-;2?�~>�j�>�
�?��?�	�����+�w�001�sS�< *�>�h?�e�>C$�> �ѽ�W!�[|�>�vl?e�>�̟>͹��7�!�^|���˽1,�>�)�>̏�>8�n>��-� U\�4m���s��uF9�;��=�h?���`3a��ۅ>��Q?��ǹA:<v�>�]t�:l!���v�%��[>�o?�=��=>ž���@�{�A��O)?�`?�1���*��!>�"?��>�w�>v!�?\��>�fþ+ű9W�?��^?�PJ?k�A?ou�>΁=�T��k�Ƚ�#'���,=�{�>	�[>y�m=�k�=X���Z�y��("E=���=�zм���߲<�b��Ȫ?<��<�v4>�7׿=D�\�ؾ3�����ZI�:R��U�%�&�:�BE�����>��犊��)E�H�½��I��M$��r��P��W�?��?�[���ۖ�S���ݢv�Y	��:�>no���ý�R����,��q��3��d���08�X�{AO�X�5�@#?	����Ͽ�ed���ѧ�#,%?�E�>�fy?�����-Y\�D�>�q��$�Q����<�� vп ���l?t�?��ݾ4���&�>�S�>w�z>��5>�v�_����u`=�e�>�2?���>���-ϿV����M�����?�r@O{A?t�(�����GV=���>�	?��?>uR1��H�����;U�>�<�?e��?�M=��W��u	�}e?�l�;��F�_�ݻ\�=B2�=V�=��y�J>W�>��HKA��*ܽ٪4>N݅>!"�����y^�|b�<��]>��սQc��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=w6�Չ��{���&V�|��=[��>c�>,������O��I��U��=����&��8P�tD$��^=tK�aq��W���2<{��
n����H������;ďs=��a>nܙ>��E>T�m>�l^?Oa�?x��>,ټ��_���ns��� <(G�'�6�?㮾Y�������^�e����� ��nh�P7=��I�=gQ����&j!�8�b��'H�P�,?��&>_zǾ0�J���'<s�˾՝��zD���Z��t�̾y�/��k����?L�=?iY��T	U�*��F�ҼY����X?sJ	����Z$��N��=
����&=L\�>_U�=u����/��,R���0?�?w���M���L)>�}�2S=J�,?�� ?*S(<K:�>G�%?}�"�G�ٽ�.`>�I1>z3�>���>��>�1���e׽:�?��T?����%˞�yX�>�¾�4}���=�7>
�3��/㼈�W>Bi�<�/���_%�k󠽨#�<<2W?ͩ�>��)�tH�x#��S*'���B=T
y?�@?���>\pk?�"C?.?�<T��ΔS����u�j=��W?�*i?��>�R��j�оާ���5?>�e?w?P>��d�3��Z�/��/�!s?��o?:�?����!}�����&�5?OP?F_^�ӑ��ҾJx��l�s>J�?��>Xx"�M?��??�������Բ�wK�� �?֭�?)��?�Ѿ=㞽��=1�!?5��>o;�����нJJ��?55>�R�>���}a�������Kо�'?gt?��>tߧ�
�/����=�ؕ��^�?c�?=�����m<���Gl�Ǖ���Q�<�ګ=���u"�v�7�6�ƾ
�
���������Ȇ>�L@N���k�>Q�8�P+��VϿ�񅿋4о�%q�O�?Kj�>�ǽb���şj�Mu��G��H��i��aj�>_�>	*���N���{�iy;�P%�����>r��1G�>��Q�Ǭ���ȟ�0H<���>���>8�>2(��`���ؙ?�����ο
x���C���X?K�?��?�?eU9<��w�h�y���!�tG?�'s?6�Y?+�%�C�Z��5�isr?�Fƾ��d��+��F����>�F6?�u�>�b1���G>Ô�=��>l㸼�#%�ƿ��즿�ԍ�x<�?��?�=վ�;�>���?�&?�C��*���~��..����=C+??=z�>��F��һ>�CRk���?{4?�.��M6�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�W�>�6�?)'���?D/�>���u ;��P>�f���<��
?��c?��?4��>X�0>� �j:$��-��xr���#0����>�Y?�aC?_�>V�h<w�Q K������MD� ���M�P���Ծ��^걼 �4>�Μ>w��֥��)7?]�)��տ����٤I��z`?�^9>ޕ?e�B�6J�����SJ?��F��;ػ�|���(�6��?�	�?}�
?8ž
�<��>�dҹ�(�>RKX>�:Ƽ(�J>|wZ?��7=�f��-U���>���?iF@��~?��=��	?J$��P��VY~�H����6�R�=��7?%;�"{>���>.V�=�tv�"�����s�̨�>�C�?Iw�?\��>P�l?Suo���B��S2=�:�>�|k?�r?Hx�z����B>-�?c��[����O�3f?��
@]q@=�^?u��ֿ�؝����_��x �;K�>��>7_��ɚ=۝�����<?�Z=��!>��>
�_>E�9>�X>->.Ű=[A��]�(��O��r���~�W���,�S�H�(`������fg��eվv���K�9d�F尿c�9���c��=нe_�=�sX?��M?\�o?U�?�����>������<�S!�]/�=Ȭ�>�2?M?�,?���=󠙾g�h�(b��Bp��o����k�>��F>���>��>��>����FP>1>�B{>�)�=�5�<v` ����<�eR>#��>���>"G�>C<>h�>/ϴ��1��j�h�Jw�W̽�?G����J��1��[9��Ŧ��h�=0b.?�{>����>пO����2H?N����)�E�+���>��0?�cW?Y�>G����T�:9>п�"�j�v`>�+ ��l���)��&Q>�l?ޖf>	2u>��3��g8��P�T���m|>:&6?ȶ�JE9�-�u���H�7aݾb.M>���>[�D�@l������ �shi��'{=�t:?�?t��.ాX�u�g?���tR>%o\>�=hN�=�UM>`�b��Bƽ4�G�؂.=ܟ�=�m^>��?(�)>ݵ�=�W�>U���82R�^۩>�B>�,>]D@?��%?�Q�\ޛ��!��=�/�^'x>��>��>�>�5K�*��=[��>Ib>�p�%冽�W��>���X>q�u��^�jv���{=F��c��=��=�7 ��=��."=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ_��>��4�uX��Jz���T��x�=[�m>��I?˵�Q<�X�����>���>��⾛���o�ʿ7~���?D��?��?fc�Bb��:�_��>���?;9U?~+F>d뾔�D�/�f>f1?.7@?���>�(��CF���	?F��?���?�X>]&�?g@d?+��>,��]l4�9շ����;��=�ӕ���m>���=��̾��L��ғ���5(m�5,� <�>L�R=˞�>0½��щ7=�ѱ�����-�(�+|�>��>�r>��>���>A�>���>o�*=�v��!��=���=�8?B��?l���mQ�"h�J������>�X?4�����!��>�De?~��?"��?�9�>$r;�\���#��"���GN=���>���>��>;� ���M;w��1�~>?y�>>>����5r�(NƾTl񼱍�>��?52�>��D>��*?7^?K�,>,?{�>�η��|!@��s
?�Ʀ>͎�>��?���>|�Ⱦ�z0��Xv� ��8��4�b>tWx?o?jW�>S���A���M/>%G��*�>Ƥ?nyE?���/�>!ó?WXX?g?�\�>�ɾ���^<�=��=�!?�&���A�g<&����M?tP?��>1��?ֽsּQ������!?;\?�P&?W��	Ha�+bþ:��<��>�Z���;"I�|�>�Z>�������=#>�C�=�m�k6�upj<�A�=�p�>��=a�6������3?!�Ͻe%��0R>5���F���>�l>�߈�'w�?`BZ=�̆�"���?���!뎾2Ju?�%�?wl�?�6n��wi��LE?�(�?l�>SG?$�)�F�ܾ.�qѕ�~��0�6�w�%=���>�=�<����̩�^A��4ǂ�p�<�k���>��#?��>�4�>cB�>u;�>�:������mg��4D�"����B5��i�b>����&�A�=����YN��¾J�`��u�>lO�u��>]��>�X@>�>[�>&�߽s��>f&o>���= �>yU�<E��>�I#>_��#�\��QS?j���/�%쾃ͯ�D�7?Va[?m-?�|e�����p�T$?��?�z�?CF�> Vg��^0�'U?�k�>_2�9�?Zn[=��ۻ��<ݙþd������;���>����3�x�@��g���?![?�"�;�㾼4Ͻ}����]=k��?��1?��.�˒*������D�#>I������}:�V���r��:|�5E��[9x�Uփ����5Dd>�2?6��?������1����
}��dU��!�>�t�>�p�>�[�>�O>!�����!��4�*3��.��y��>bZ? XI>y49?8b?��?��d?Q.�>\�>#�����(?�P)�}D>��>]c+?H�?9&?�<<?�=??	�e>�����-쾮��On?��?J0?o�?�2?׿������`�/�R��;vw��s|׸��A=�G���A��䛽@ؤ=�P�>�Z?��R�8�4���>�j>�}7?�z�>���>K��B;�����<��>��
?EN�>�����}r��e�T�>)��?Y��=��)>���=�o��WEۺ�M�=�s¼V�=�����k;��q<j��=�=dp�n-�Ҹ�:s��;L�<9�>��?X�>��>�:���b ����7�=c�X>�[S>��>��پ`����&����g��,y>�\�?�^�?�Lf=CP�=Ӵ�=E��Y���!�������`�<?��"?�T?&��?o�=?�{#?1g>�
�M,���k��ue����?�),?P��>{�:�ʾڨ�C�3�M�?l�?"a�
����(��¾�ҽK>/��~�o���9D�R������阽��?���?��>���6��N�Z֘�����1�C?��>*R�>m��>&�)�	�g������;>R��>N�Q?��>s{T?�3p?P�Y?{V>�n<�������������>�R>?�-�?v��?0ey?���>��6>�K��?�����)������������<5�L>gx�>�q�>d�>
��=��$ȽҀ��>�m>��>$ط>��>Yut>�	����G?���>�J��^M��O�������<�g�t?���? +?=d��vyE�a���$��>I��?�߫?��)?V�U����=�M뼍��1Aq�w��>9�>��>��=��7=�,>G��>��>X�:�|�8�sHN��=?i�F?H��=������]�%�r�H{��'m.����ǉ��_-ý$J"���=n����V績2���W���Ң��þ�ᓾ�*?�6<?�0'<�=��=�e��"��O3=���=J˱�&#�=6s�� �n=�x�e�<�?<+G�<�L�;�e
=�7��R�˾3�}?r;I?Δ+?z�C?<�y>�>>x�3�^��>���@>?�"V>�P�^��Au;�ӣ�����M�ؾ}|׾~�c�V͟�H>�VI�ϵ>93>*I�=��<� �=��r=�Ŏ=0�Q�{=Z;�=�G�=�h�=:��=�>dE>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>X`7>�j>_�R�h�1�^�\�1c�}�Z��!?%-;��D̾��>�N�=�߾��ƾ��-=�i6>
a=���=\�p�=�V{���;=͈k=��>̫C>o�=ׯ���=��K=(�=��O>O���m6��[*�ϻ4=���=	\b>3l%>���>��?^0?4Zd?�8�>�n�LϾ+=��`F�>���=�G�>���=�nB>���>��7?�D?��K?q�>ᓉ=��>L�>D�,���m�|w�.ɧ����<���?9͆?�ȸ>��Q<w�A����c>��4Žw?mR1?�g?՞>H��8�߿a���?���i�=v8�<�9-��D�� e�� 1�����^	��z�=�K�>���>5��>���>-�=��=�@�>�5P>�
�ۣ�=�<1>�[���=.f�=ć�=w���Q��9`�{�޽��0�q"��S�=7a==��=���=:�>A�>�Æ>Ζ�>x�������>�k��AM�Ad�>�ྗe�zDY�O�����(����<
>�r�>�(�<}я�J�?�,�>�q�=���?�{?~U�=/lv����0鞿yH���nn��P=��X='3U��"?��c��b�g潾���>�Ď>�[�>Xl>��+���>��gw=��k5�JG�>���n:"�!��q[q�0��*��h��O���D?�?����=~?�qI?KЏ?T��>䪘�ޔؾ/e0>������=\��P�q��F��|�?�'?���>�:�f�D��*㾧������>44q��BQ�U����B���;�x��"$�>uh��C�žF!2�����|w��K?������>˝A?���?͔��2Nt��7����>�F}?�Cc?\��>Z|?U?@�U�|Ⱦ�96��Yd>dEg?�*�?
S�?���:�$�=���PQ�>��?^�?q�?YXt?�I��)�>�铻��>�����=��>��=Z+�=��?�	?�?쟽c�����(�ﾺ�P��=���=��>�I�>�q>��=�8i=Uj�=	�d>�J�>�k�>�R[>�H�>܋>���J�
�})(?��=���>> 2?�8�>�@=3"����<�PY�9�?�\�+�����8��G��<Ҫ:�1W=���,��>8kǿ��?uQ>��f�?�D�#�.�Q=H>VaR>�׽���>	oG>W>J�>�z�>>�ш>
�)>mؾ��J�<���0��r;��2�sn��,��>����Y��� � ��W���վ#g��zZ�5fv����`L�=��?/��~La��&/�g��=�g/?*#v>�GX?���ʋa���j���>`x�=/���JF�����U~�&�?���?�5c>��>��W?��?ԕ1�� 3�IoZ���u�%A���d�'�`�V㍿����j�
��5���_?��x?�wA?��<�-z>ݟ�?�%��ˏ��&�>�/��#;�$<=�'�>X,����`���Ӿ/�þF&��3F>A�o?�!�?\S?�RV�' �m5a=�Y?kU?�ǜ?pgv?8b�?]����9?4_�=�1?�ę>s�=?>�5?�C?>Z�>F`j>�K_<Tz���K��]���tE`�-�=p�X�<�b=�q�=|����:B�>��=~8�3�H<��o>Wu�=���6�X��6=.9�>K��>q�]?���>��>�M7?Y|���5�񄱾<i2?��"=�ǂ�G���:8��h ��>�ol?}��?��X?�1W>/C�l�Q�6W(>���>�a->	zj>}��>iD���\Y��g=�>Z">��=pD���冾��	�����=h#>ڗ�>��>�C����>1������o�=>$x������2J��$:�zm1�2�:��v�>��R?U9?uo >2a��=A�:'^����>p�U?��D?��|?/^3>����!<�X�S�]#c��{�>Y�=Ip ����������a$����=���>Y(�������a>���G�޾Gyn��5J�x9�#I=����V=d��!�վq����=S>�
���� ��͖��Q���J?��_=�_��ogT�Mߺ�`�>#�>H�>��<���k��o?�6j��7��=J�>G>>�`������	G�����G�>��X?��@?Cȅ?Z�V�nm�ٸ2��꾊���(dֽ{M?���>5��>�Z�>#�.>ލ�U�����QO\����>6�>q���+N���˾v���H����\>i�>��4>���>�Q?�S(?6>P?|�?��?�!�>�!ͽ ���'�?�7�?(^�����Bz��P���ھ�!�>�v�>�(��Sx>��O?W�P?�O?��d?O#K?�C>��W�������z>z�v>m36��ꢿ�'�=�1?�M�>�B? Af?C!;>a<6�������Cp>D�>@e'?���>�?iI�>��>�������=���>��d?�ރ? �p?�|�=��?�j,>���>�Ζ=�;�>h4�>�0?��O?@s?��I?hV�>�c�<�+���f����l�ANv�^
�;�?<�#t=;M��j������<-J�;
�j�VS�����Q�E祿)�X<��>
{>������->vþp?����<>�i��n��l��}�*��`�=�
�>ͧ?�ϛ>�>%�D�x=���>C�>�q���'?��?�?��H<�Sc�)�׾�!d��K�>U�F?&+�=��i��ߒ�8zu�:`h=$?n?*%^?�ym�D��ɍg?�O?ˀ'��Z���籾)��
��L<�?j/�>��A�`�?���?g��?A�?kż�(��ߩ�O��2*�_Ղ=�\�>������j@:>�2?�'>�U{>�k�=�3���'�W(\�4�!?�	�?�E�?�҆?y�>�g�=ɿ���L��/x[?�H�>XK��>� ?i����Ѿ�����ё���pê��Э�$5��tԨ�\n&�����X�ѽ���=��?��u?��o?�]?� ���c��M^�tE|���U�����>�zE�x�E��F�/�p����'<������9m=�1V�O�,��?>�%?��H���	?���]\ �y�����n>hq��4����p��j]��������<����j�K!F���?��>�7g>�1g?3�W��� �j�H����ս�� >� ?�pe>�h?���=
E�dU%�͆��D����Y>Q_v>��c?�&K?��n?����&1�vf���^!�ä1����-�C>o>�a�>��U�����%�M�=�	ms���62����	��=-;2?�~>�j�>�
�?��?�	�����+�w�001�sS�< *�>�h?�e�>C$�> �ѽ�W!�[|�>�vl?e�>�̟>͹��7�!�^|���˽1,�>�)�>̏�>8�n>��-� U\�4m���s��uF9�;��=�h?���`3a��ۅ>��Q?��ǹA:<v�>�]t�:l!���v�%��[>�o?�=��=>ž���@�{�A��O)?�`?�1���*��!>�"?��>�w�>v!�?\��>�fþ+ű9W�?��^?�PJ?k�A?ou�>΁=�T��k�Ƚ�#'���,=�{�>	�[>y�m=�k�=X���Z�y��("E=���=�zм���߲<�b��Ȫ?<��<�v4>�7׿=D�\�ؾ3�����ZI�:R��U�%�&�:�BE�����>��犊��)E�H�½��I��M$��r��P��W�?��?�[���ۖ�S���ݢv�Y	��:�>no���ý�R����,��q��3��d���08�X�{AO�X�5�@#?	����Ͽ�ed���ѧ�#,%?�E�>�fy?�����-Y\�D�>�q��$�Q����<�� vп ���l?t�?��ݾ4���&�>�S�>w�z>��5>�v�_����u`=�e�>�2?���>���-ϿV����M�����?�r@O{A?t�(�����GV=���>�	?��?>uR1��H�����;U�>�<�?e��?�M=��W��u	�}e?�l�;��F�_�ݻ\�=B2�=V�=��y�J>W�>��HKA��*ܽ٪4>N݅>!"�����y^�|b�<��]>��սQc��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=w6�Չ��{���&V�|��=[��>c�>,������O��I��U��=����&��8P�tD$��^=tK�aq��W���2<{��
n����H������;ďs=��a>nܙ>��E>T�m>�l^?Oa�?x��>,ټ��_���ns��� <(G�'�6�?㮾Y�������^�e����� ��nh�P7=��I�=gQ����&j!�8�b��'H�P�,?��&>_zǾ0�J���'<s�˾՝��zD���Z��t�̾y�/��k����?L�=?iY��T	U�*��F�ҼY����X?sJ	����Z$��N��=
����&=L\�>_U�=u����/��,R���0?�?w���M���L)>�}�2S=J�,?�� ?*S(<K:�>G�%?}�"�G�ٽ�.`>�I1>z3�>���>��>�1���e׽:�?��T?����%˞�yX�>�¾�4}���=�7>
�3��/㼈�W>Bi�<�/���_%�k󠽨#�<<2W?ͩ�>��)�tH�x#��S*'���B=T
y?�@?���>\pk?�"C?.?�<T��ΔS����u�j=��W?�*i?��>�R��j�оާ���5?>�e?w?P>��d�3��Z�/��/�!s?��o?:�?����!}�����&�5?OP?F_^�ӑ��ҾJx��l�s>J�?��>Xx"�M?��??�������Բ�wK�� �?֭�?)��?�Ѿ=㞽��=1�!?5��>o;�����нJJ��?55>�R�>���}a�������Kо�'?gt?��>tߧ�
�/����=�ؕ��^�?c�?=�����m<���Gl�Ǖ���Q�<�ګ=���u"�v�7�6�ƾ
�
���������Ȇ>�L@N���k�>Q�8�P+��VϿ�񅿋4о�%q�O�?Kj�>�ǽb���şj�Mu��G��H��i��aj�>_�>	*���N���{�iy;�P%�����>r��1G�>��Q�Ǭ���ȟ�0H<���>���>8�>2(��`���ؙ?�����ο
x���C���X?K�?��?�?eU9<��w�h�y���!�tG?�'s?6�Y?+�%�C�Z��5�isr?�Fƾ��d��+��F����>�F6?�u�>�b1���G>Ô�=��>l㸼�#%�ƿ��즿�ԍ�x<�?��?�=վ�;�>���?�&?�C��*���~��..����=C+??=z�>��F��һ>�CRk���?{4?�.��M6�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�W�>�6�?)'���?D/�>���u ;��P>�f���<��
?��c?��?4��>X�0>� �j:$��-��xr���#0����>�Y?�aC?_�>V�h<w�Q K������MD� ���M�P���Ծ��^걼 �4>�Μ>w��֥��)7?]�)��տ����٤I��z`?�^9>ޕ?e�B�6J�����SJ?��F��;ػ�|���(�6��?�	�?}�
?8ž
�<��>�dҹ�(�>RKX>�:Ƽ(�J>|wZ?��7=�f��-U���>���?iF@��~?��=��	?J$��P��VY~�H����6�R�=��7?%;�"{>���>.V�=�tv�"�����s�̨�>�C�?Iw�?\��>P�l?Suo���B��S2=�:�>�|k?�r?Hx�z����B>-�?c��[����O�3f?��
@]q@=�^?u��ֿ�؝����_��x �;K�>��>7_��ɚ=۝�����<?�Z=��!>��>
�_>E�9>�X>->.Ű=[A��]�(��O��r���~�W���,�S�H�(`������fg��eվv���K�9d�F尿c�9���c��=нe_�=�sX?��M?\�o?U�?�����>������<�S!�]/�=Ȭ�>�2?M?�,?���=󠙾g�h�(b��Bp��o����k�>��F>���>��>��>����FP>1>�B{>�)�=�5�<v` ����<�eR>#��>���>"G�>C<>h�>/ϴ��1��j�h�Jw�W̽�?G����J��1��[9��Ŧ��h�=0b.?�{>����>пO����2H?N����)�E�+���>��0?�cW?Y�>G����T�:9>п�"�j�v`>�+ ��l���)��&Q>�l?ޖf>	2u>��3��g8��P�T���m|>:&6?ȶ�JE9�-�u���H�7aݾb.M>���>[�D�@l������ �shi��'{=�t:?�?t��.ాX�u�g?���tR>%o\>�=hN�=�UM>`�b��Bƽ4�G�؂.=ܟ�=�m^>��?(�)>ݵ�=�W�>U���82R�^۩>�B>�,>]D@?��%?�Q�\ޛ��!��=�/�^'x>��>��>�>�5K�*��=[��>Ib>�p�%冽�W��>���X>q�u��^�jv���{=F��c��=��=�7 ��=��."=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ_��>��4�uX��Jz���T��x�=[�m>��I?˵�Q<�X�����>���>��⾛���o�ʿ7~���?D��?��?fc�Bb��:�_��>���?;9U?~+F>d뾔�D�/�f>f1?.7@?���>�(��CF���	?F��?���?�X>]&�?g@d?+��>,��]l4�9շ����;��=�ӕ���m>���=��̾��L��ғ���5(m�5,� <�>L�R=˞�>0½��щ7=�ѱ�����-�(�+|�>��>�r>��>���>A�>���>o�*=�v��!��=���=�8?B��?l���mQ�"h�J������>�X?4�����!��>�De?~��?"��?�9�>$r;�\���#��"���GN=���>���>��>;� ���M;w��1�~>?y�>>>����5r�(NƾTl񼱍�>��?52�>��D>��*?7^?K�,>,?{�>�η��|!@��s
?�Ʀ>͎�>��?���>|�Ⱦ�z0��Xv� ��8��4�b>tWx?o?jW�>S���A���M/>%G��*�>Ƥ?nyE?���/�>!ó?WXX?g?�\�>�ɾ���^<�=��=�!?�&���A�g<&����M?tP?��>1��?ֽsּQ������!?;\?�P&?W��	Ha�+bþ:��<��>�Z���;"I�|�>�Z>�������=#>�C�=�m�k6�upj<�A�=�p�>��=a�6������3?!�Ͻe%��0R>5���F���>�l>�߈�'w�?`BZ=�̆�"���?���!뎾2Ju?�%�?wl�?�6n��wi��LE?�(�?l�>SG?$�)�F�ܾ.�qѕ�~��0�6�w�%=���>�=�<����̩�^A��4ǂ�p�<�k���>��#?��>�4�>cB�>u;�>�:������mg��4D�"����B5��i�b>����&�A�=����YN��¾J�`��u�>lO�u��>]��>�X@>�>[�>&�߽s��>f&o>���= �>yU�<E��>�I#>_��#�\��QS?j���/�%쾃ͯ�D�7?Va[?m-?�|e�����p�T$?��?�z�?CF�> Vg��^0�'U?�k�>_2�9�?Zn[=��ۻ��<ݙþd������;���>����3�x�@��g���?![?�"�;�㾼4Ͻ}����]=k��?��1?��.�˒*������D�#>I������}:�V���r��:|�5E��[9x�Uփ����5Dd>�2?6��?������1����
}��dU��!�>�t�>�p�>�[�>�O>!�����!��4�*3��.��y��>bZ? XI>y49?8b?��?��d?Q.�>\�>#�����(?�P)�}D>��>]c+?H�?9&?�<<?�=??	�e>�����-쾮��On?��?J0?o�?�2?׿������`�/�R��;vw��s|׸��A=�G���A��䛽@ؤ=�P�>�Z?��R�8�4���>�j>�}7?�z�>���>K��B;�����<��>��
?EN�>�����}r��e�T�>)��?Y��=��)>���=�o��WEۺ�M�=�s¼V�=�����k;��q<j��=�=dp�n-�Ҹ�:s��;L�<9�>��?X�>��>�:���b ����7�=c�X>�[S>��>��پ`����&����g��,y>�\�?�^�?�Lf=CP�=Ӵ�=E��Y���!�������`�<?��"?�T?&��?o�=?�{#?1g>�
�M,���k��ue����?�),?P��>{�:�ʾڨ�C�3�M�?l�?"a�
����(��¾�ҽK>/��~�o���9D�R������阽��?���?��>���6��N�Z֘�����1�C?��>*R�>m��>&�)�	�g������;>R��>N�Q?��>s{T?�3p?P�Y?{V>�n<�������������>�R>?�-�?v��?0ey?���>��6>�K��?�����)������������<5�L>gx�>�q�>d�>
��=��$ȽҀ��>�m>��>$ط>��>Yut>�	����G?���>�J��^M��O�������<�g�t?���? +?=d��vyE�a���$��>I��?�߫?��)?V�U����=�M뼍��1Aq�w��>9�>��>��=��7=�,>G��>��>X�:�|�8�sHN��=?i�F?H��=������]�%�r�H{��'m.����ǉ��_-ý$J"���=n����V績2���W���Ң��þ�ᓾ�*?�6<?�0'<�=��=�e��"��O3=���=J˱�&#�=6s�� �n=�x�e�<�?<+G�<�L�;�e
=�7��R�˾3�}?r;I?Δ+?z�C?<�y>�>>x�3�^��>���@>?�"V>�P�^��Au;�ӣ�����M�ؾ}|׾~�c�V͟�H>�VI�ϵ>93>*I�=��<� �=��r=�Ŏ=0�Q�{=Z;�=�G�=�h�=:��=�>dE>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>X`7>�j>_�R�h�1�^�\�1c�}�Z��!?%-;��D̾��>�N�=�߾��ƾ��-=�i6>
a=���=\�p�=�V{���;=͈k=��>̫C>o�=ׯ���=��K=(�=��O>O���m6��[*�ϻ4=���=	\b>3l%>���>��?^0?4Zd?�8�>�n�LϾ+=��`F�>���=�G�>���=�nB>���>��7?�D?��K?q�>ᓉ=��>L�>D�,���m�|w�.ɧ����<���?9͆?�ȸ>��Q<w�A����c>��4Žw?mR1?�g?՞>H��8�߿a���?���i�=v8�<�9-��D�� e�� 1�����^	��z�=�K�>���>5��>���>-�=��=�@�>�5P>�
�ۣ�=�<1>�[���=.f�=ć�=w���Q��9`�{�޽��0�q"��S�=7a==��=���=:�>A�>�Æ>Ζ�>x�������>�k��AM�Ad�>�ྗe�zDY�O�����(����<
>�r�>�(�<}я�J�?�,�>�q�=���?�{?~U�=/lv����0鞿yH���nn��P=��X='3U��"?��c��b�g潾���>�Ď>�[�>Xl>��+���>��gw=��k5�JG�>���n:"�!��q[q�0��*��h��O���D?�?����=~?�qI?KЏ?T��>䪘�ޔؾ/e0>������=\��P�q��F��|�?�'?���>�:�f�D��*㾧������>44q��BQ�U����B���;�x��"$�>uh��C�žF!2�����|w��K?������>˝A?���?͔��2Nt��7����>�F}?�Cc?\��>Z|?U?@�U�|Ⱦ�96��Yd>dEg?�*�?
S�?���:�$�=���PQ�>��?^�?q�?YXt?�I��)�>�铻��>�����=��>��=Z+�=��?�	?�?쟽c�����(�ﾺ�P��=���=��>�I�>�q>��=�8i=Uj�=	�d>�J�>�k�>�R[>�H�>܋>���J�
�})(?��=���>> 2?�8�>�@=3"����<�PY�9�?�\�+�����8��G��<Ҫ:�1W=���,��>8kǿ��?uQ>��f�?�D�#�.�Q=H>VaR>�׽���>	oG>W>J�>�z�>>�ш>
�)>mؾ��J�<���0��r;��2�sn��,��>����Y��� � ��W���վ#g��zZ�5fv����`L�=��?/��~La��&/�g��=�g/?*#v>�GX?���ʋa���j���>`x�=/���JF�����U~�&�?���?�5c>��>��W?��?ԕ1�� 3�IoZ���u�%A���d�'�`�V㍿����j�
��5���_?��x?�wA?��<�-z>ݟ�?�%��ˏ��&�>�/��#;�$<=�'�>X,����`���Ӿ/�þF&��3F>A�o?�!�?\S?�RV�' �m5a=�Y?kU?�ǜ?pgv?8b�?]����9?4_�=�1?�ę>s�=?>�5?�C?>Z�>F`j>�K_<Tz���K��]���tE`�-�=p�X�<�b=�q�=|����:B�>��=~8�3�H<��o>Wu�=���6�X��6=.9�>K��>q�]?���>��>�M7?Y|���5�񄱾<i2?��"=�ǂ�G���:8��h ��>�ol?}��?��X?�1W>/C�l�Q�6W(>���>�a->	zj>}��>iD���\Y��g=�>Z">��=pD���冾��	�����=h#>ڗ�>��>�C����>1������o�=>$x������2J��$:�zm1�2�:��v�>��R?U9?uo >2a��=A�:'^����>p�U?��D?��|?/^3>����!<�X�S�]#c��{�>Y�=Ip ����������a$����=���>Y(��Qh���4g>-���޾�Pl�U�H�I��<=�W��N=�����վC7|����=�5>Ţ��R� �B���r����I?D�f=d���V�W�珺�ժ>}��>I��>gP/��|��@��)���^�=Ho�>��:>�������o�G�������>��D?Z�^?켃?�I���qr���A����v�����U;?��>�-?X�7>|�=B���c�޿d���C��1�>)f�>�X��H��N���W뾖f ��>�)?1�>7�?n�Q?��?�]_?��&?Κ?�m�>錧�D���q&?��?0�=�Խ{�S���8�e�E��W�>�)?ȓB�)C�>�g?��?�'?p�Q?��?�:>B� �i9@���>\��>��W�hW���_>�J?(³>�Y?5̓?�
=>��5����ı�����=��>��2?�-#?�U?�I�>W��>Ʈ��\�==��>�	c?r1�?=�o?��=j�?�22>���>S
�=���>��>�?�VO?�s?c�J?���>���<	:���>���Qs���O�M7�;7�H<�y=Ԝ�:t�V�غ�<���;dQ���B�����k�D����D��;K�>�@|>�����@$>!��������V4>Pp��ޢ�a�����)�9��=ь�>��?H�>g� �`UM=BX�>|/�>�� �z$-?��?PB?��<0{b�BY�$`y�ڰ>#@G?a'�=��h�=g��y�r��S�=��s?G�\?^U_����B�b?ߧ]?����<������la�{����O?�Y	?��I�F�>|�~?c�q?� ?8�\���m����s�b��-n�Lr�=�>�M��Yd�Ɵ>D�5?[3�>fRY>C�=� ׾�v�g���?�y�?\$�?��?V�*>p�n�I��͙�������]?Ҍ�>�����"?c�
�1Hо=��ڞ��ޅ�nH��/���q��d���F$�����X׽e��=xe? �r?�yq?�A_? ��Nc��^�����lV�k,�0��E�s.E�~�C���n�3N�i9���,��&�D=k�r�R<�^��?*�6?��2�ru�>�.�~:��$��W�}>@w�B4¾؇�<7U����=�{^�ܯL�~���9�?{��>W�8>�YR?:�Q��$F�%�ep����ݾ�ku>�^�>�^�>u�?�)>q���`����8|2�o��=���>U*a?pJ?�ij?�%!�X�.�J�}�'���̋��ȡ���C>P�>�r�>"gc�ƛ#��2&�>�7��Sp���
����#L�혁=��&?��d>k��>���?b��>����+���SL���(�5-�<�)�>�@_?M�>�_�>����!*����>�iq?�X�>�߳>�x��OM&��(n�� �49�>\�>H��>A�>�J�o�S�"���"m���1.���c=\tx?a�r�?�y��'�>Ѓ??������9���>���bP����\\G����=̈́�>�T<-�.>�F��"����Si��镾ց?W�"?���;8$���>��-?�o�>(~$>R3�?�x>{����[?�mz?�o_?=�7?���>f�佨b0�j&���I��/v=�4>�I)>��=�I�=,m�QE3�þR��v�X�^=-P��|�н�W=a=P<=���1	>DNۿI7J�g�ھ>���d�[�
�e牾J��`�����0\��? ������8�0���P��v]� ۍ��!o� ��?���?����D��� 䙿r*��g@ �+v�>B�k�v�v���������,����侵��з ��hP�E�i���c�rz'?:�����ǿƬ��ܾ� ?M ?n�y?�͡"���8�h!>���<������뾆�����ο z���^?E��>P?�������>+^�>w�X>�-q>�����Mԓ<��?�~-?|��>��r�C�ɿ�s��/I�<W��?��@E�W?���GhY�fz�=��=hG?�}(?:��=�@�D���?ݟ?�@�?��>�z:�L5J�x9j?f^�=��g���h=� ��:���\l���T=|g�>�?5��0������@�P>a��>��>�4>��Ԣ�;�<0>�Ǉ=|M�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=4��E����`�
h�r��:ur�=H��L]j=����z���̾DQȾ0K�=h)e>,/?-��>����b<��P?%Lz?L�>�-J>��=qԾ��޾(�=�H&�|t�7���{��Sa�?���s��Eh�����`����O�af�={R�$r����e�d��OI�Xy+?�Af><��tgo�O��JHľ�ؽ�qu<s����<�!CX���?R4H?��n��qZ�XZ���5���#�W�P?|��O�;��d�� >�����q1J>	+	= [��7��%��`0?�N?=V���I��6� >����	=�`+?C?�6�<:��>�w%?Be%��(彚�U>VJ,>1=�> -�>�>�!��r`ٽT�?��R?F����EA�>_h��D�|��(e=��>+u5�iO��+�Z>=��<���n0�e�����<�\S?�Ȯ>�L��®����=5����=T�|?ħ.?4��>Z��?��E?��>���Z�k�l�S�<߳?�O|?R�=T�`=ȩ��e���U�>%�R?)�>�:��ܕ�\��ȥ��-?W =?�\B?��D��B������o��5?�l?+�p��ꑿD���图4�>=��>]2z>����-�>B�`?Gj�pvs�r��c�(��e�?�1�?i��?� ������Cx�=V�5?�o8?k����]��(����V�>��>?�S��Ch����6����P~"?��z?�?��[�t����=ڕ�![�?��?�����Ig<����l�po��Q��<gΫ=p"�uD"������7���ƾ �
�9���Wؿ�Ӧ�>�Y@2c轧,�>,E8�x6��RϿ���c[о�Nq���??��>��Ƚ����g�j�!Ou�S�G�D�H����P��>nF>�C�怈��C���5���G�>5H�lT�>�8��������n��؅>Q��>� �>i���9��lt�?#���
ǿ@���&��/5a?�
�?��?G?���4�8���T���`<uML?�Ug?QR?J�3���+�ySٽ�Yj?|Ӳ��b�NS2�J*E��\`>��/?#��>fD.�T�\=A >���>�\>��0��ÿ��������Ae�?��?5��&��>r��?�U-?p���Y�������)�TA�;#�D?�C>o�Ǿp�!�59�򱇾	?�m7?z��e��]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�N�>mǊ?B@I=��?�8<5:ؾ[��>�om>��}>�?_�G?��>Y��=Co�4�m5���Q��'���,�b �>{Ic?�G-?���>K+ս�
��3��S4�#Hn���6��Mr�qʎ<��^��u�>�C�=CP>O��@���$?��8��,ֿ�^���U���@?�**>���> �٤��E�<�~Q?n��>!)�(t��87��(Y�B��?��?�?v�վ!>߽`�>H�>��k>n;=q�~�]�]����>��T?,����j��S����>���?�e@͗?��B�5-	?�c��b���~����I�5� 3�=�y7?�n�w�y>J��>�#�=�v�I���/�s��=�>��?#r�?���>6dl?�6o��{B�X\7=�h�>�k?��?���ۅ�^D>,�?���Y掿 ��,f?��
@Xx@�]^?ز����տ㯝� wϾ�MȾ�=#\�=�=p>�g�Y>.�Z:�������>�j�>�5i>i��>G�P>�>I�=7L���(��~����]{b��z��� ���r�5X�4���r�	��8��gί��F��(�+��
:j�7�%�n�ָ��S�=�G�?��#?B�$?��k?��=���<4>���=��
�6�2�mӚ>�1c?eR�?~�t?��o����K��7���(Ͼ�6��^>��[>nZ�>���>��>��{�>٧�=^�<BeV��[<=�m�=�n%�R�>:�>O0�>�R�>�97>?&>����}I��lg�Qhy�@~ҽ��?ɚ�f�J�hp��y&��`��-��=A6-?�>����п�:��2H?9풾�����+���>� 0?1�V?T>����l�J�ӹ>7b�h��Z>�Q�΃m���)�<�P>��?��V>��~>�b4��:��%L�!s���{m>ȿ5?�'���?�8�w��F��㾑D>��>����O�b���Q�y�2R]�l7=G9?��?��������r�Lc��Q�M>��b>�(=!{�=	dQ>5�3��~ڽ[�L��=j\�=3�g>[?��c>���=�پ>~���~��"�>��|>��R>�G?
t?�#:ZC�����"�1���#>m��>O�E>Ͻk>F*� }<���>��'>�MýB�N�u��[_8��]l>/���?�B|� �<��+��=}�=�A���F#�W���~?���(䈿��e���lD?S+?^ �=
�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�ú>�Tq�ۊ�47���>[��u�=���=��`?ow���W�	Ï��s$?1��>��+f���0���G���?�C�?u8�?1䇿���������=j��?��d?:p�<Ɋ��9�B�̵�>��?�,]?�?�>���CnX��M?��?4Z??�I>���?Dns?`��>�|��q/����aA���&�=ab�;�%�>��>]K���SF�D����\���vj����/zc>}E%=�c�>i.�v_���״=���	���Ah�A��>�ro>ܺI>1#�> l ?���>�R�>'=8�������2����E?*�?m��l�d�~��=5��=�A��~J�>�?��������5��>�r`?{M�?��?+-�>����T��,ƿ+ྤ�>�Mu>s�>�?� ��6c�=�������a�>�f>�Kͼ����(��sf"<�+�>�R?�>B���c"?��#?8U|>o׶>�9L�褎��|=�>��>\��>`u?Rp?��?׫�a�3�<����{���N���>�t?�O?�h>�҇�(Ҝ�_�x����<bûf%f?��X?σ;�Ȼ?R�?��*?��??��7>�������&���=>�| ?���ͷ@���%����Y	?��?���>��|�n6ٽb��b���Q���K?�_]?�%?���G@b���ľ��<~�X�r�����:�Qm���>|>?A���`�=_|>�=�Qn��k9��gN<ib�=˪�>M��=��>��ꐽQ&?XYݽa�.��Z�>�5^��hT��a_>�9j=H�^��8t?��;J� %���Q��kq�B��? ��?X��?ނ"�`�l�Y2?70�?�?�s?�����侖PѾ�/s�6��#{@� �<��'>Ei<����Sj�������F��R09��h>�Ί�>.�/?�Y?��?ӯN>��=x��z �~�z�we����^H��'B�1������������ɽ�E#�?ݵ��I�����>��n��>�U?�dQ=��>d%2>ܭ����>i�b>$�>/e�>I@">.>��,>�#�=�vA��_?Rޢ�x���̾�uf���q?��?�n?���˰��(0��ZDJ?�&�?,�?�M�>�W���b6���>*U?8ߝ�0?�GJ��h���B�>�p�׿��3��Њ=���>��ڽ���+�T�P=��n?}�?:�f�\���0������n=WR�?��(?g�)�|�Q���o�!�W�� S�R��`h�擡���$�Sup��׏�QR������u(��',=��*?��?~�����+���1k���>�+_g>	��>H*�>þ>��I>��	�/�1�Z�]�'��p��\N�>�={?$��>�J?��;?�O?8*M?��>,��>=b��r$�>d��; W�>C��>e:?ɳ.?��0?��?��*?�a>8���1��kؾQ�?��? ?H?o�?�����ڼ�$"����x�v|����� �=J�<Z�׽�s��T=۶T>�R ?�:#�!l1���w*J>�6H?'?DT�>칮���@p=���>p�?/@�>Ea���r��z����>��{?�
(��=�>��=��3 �G'�=����}{=�/���o��;����=!n�=x=s#g�u^)�L6<���=��?�Y??(�>>�>،��u
�:����=�>>*�T>��վ}������g@^�5m�>Z
�?���?�K�=��=�d�=����ξV��4ˢ��{:=�Q
?�*?�i8?0�?yM?+?ײ�=CE!�J͉���� Q���?2!,?���>x��۳ʾW�É3�I�?X[?*<a�Ҹ��;)�܏¾��Խ��>K[/��.~����WD�����z}�� ��?���?�A��6��y达����[��h�C?�!�>TY�>��>i�)��g��$�1;>���>�R?o�>��V?�t?�U?��>Jh/��թ�r��{�<g>�h7?�$|?&_�?�Ȁ?�d�>dc>kN@���Ot��Ɨ)����嗂� nH=�>>5�>��>���>��>��ѽ
����X�]ݓ=�W>�>>�*�>]�K>�g�<�F?z�>rȨ�Vj��E���[��>��\�r?���?Ep8?_��=r>�_z9��>�k0�>M��?p��?F+?�*���=�Z�N�������N�p>{\�>3Q�>�~�=���=�q=}��>�B�> 2���,�zDE�z�9��K�>81?C;�=����A�/�1¤�E�����=3����雾�,�<\F<��U�Q���,��%���Du�m⿾'~c�;ƾB]ɾ_��2�?�l�=+>���=���=u��z�d�=&�����=W��i#>���<͖N=�@*�
�k�y���L�>�j�=x˾!}?Z�I?Ĝ+?"�C?
fy>��>#F<� �>%��~�?VS>��Y�����}�;�8����*��sؾ�w׾�1d�������	>�>M�h�>24>'��=�X�<���=��p=���=��9��=}P�=�/�=��=N�=vw>0�>�6w?X�������4Q��Z罤�:?�8�>_{�=��ƾr@?��>>�2������yb��-?���?�T�??�?Bti��d�>L���㎽�q�=H����=2>p��=w�2�T��>��J>���K��K����4�?��@��??�ዿТϿ5a/>�T
># %>1�S��'9�.?���~��2s�9!?��(�J�о��A>)��=�Z��Ǿ��<�6> ��<��:�uN�)��=�a_�W�y=��=��>1�9>��=���=�Q�=Z�=��j>�ƀ<��?�� ��EH�<vs�=B�v>�tB>/��>�h�>b8?�!�?�J�>wL��A���_�1�>B��>3�>��F�>��?>�w"?J�.?�th?��>�O>�a�>�A�>i\J��C��
������*>�͂?�j�?V��>��t>���=�g�(�i�"����J?WW/?��>Rx�>�9��}�~q2��a;����v�H=�P�= C��:B��鹽?�|B�G�='��>u�>�f�>j�>P֛=f]'>L�>�>@T���*�=���*�=�5|���I>��';�ZĺчX��dk���Ƿ��R��<ul�<�C(=sϿ��V�<�f�=�A�>p�>��?���=!�Ǿ #�=FȾJ+���G>��_\�Tt���q�*����+��k">m�g>��3�p��pa�>ʎ�>JL==
��?BSx?��5=�aD�u*������K����u��:��p^&��i��e8���u�	k�^)��j��>z��>��>��l>�,�"?�	�w=��ᾼC5��+�>�b���
�q�*q��6���li�=��|�D?g<����=�~?��I?�܏?Ձ�>e"��S�ؾr0>9���=���6q��S����?��&?׊�>f쾵�D�w�Ⱦ�U�����>�bL�[�L��g����2���;hǶ�Ա�>�'����ɾn�1��<��L����@�Et��
�>X'O?���?BNr�K����OK����ɝ`�ι?��d?(�>�?(?©��k�往������=�k?S��?z��?A\�=}r�=�,��5�>,�?��?H��?��r?��E���>.��;Y">�!���D�=3�>Z[�=CT�=�?+	?5_	?�雽��	���߀�]�`�y�=�;�=�#�>� �>{�n>�q�=�Z=R��= �Y>3��>P��>��e>6��>�W�>UD��Ħ
��+?�o�=*J�>r�/?1j>�V=�������<�b�VL���8�E�ͽw�뽕.�<,�����U=mZ��K�>>�ſm��?jzR>��%)?Mo�t���E>vDF>�\ý7R�>�]>�>e̫>�u�>ֲ>q�>�&>R�۾8�\>e��,�8� ���P�}���_�>9\>��m�h-+��+B<𺡾�ھ�(��@��2���.�؆X>\X�?�����3�����/r9���?�>�:;?tLҾz�$�ioV>1>?"��>t+��7��z�l����ދ?��?��`>���>�[?7U?�$��E4�ݮY���s��B���]�OA]�␎�f�~�Ӧ�3���BkY?� v?>�@?U �<r��>l�?|�+�������>Ѝ5���3�ۛ�=�z�>�$��U�_�̾�������&�@>�qo?Ma�?J�?��L���n��3)>�v:?Ka1?{�t?G�1?D;?@\��$?�43>f?�Q?��5?�e/?�=?^�0>�4�=���#=2������g�ҽ��Ƚ;g��`5=��}=����.<,=Fɞ<i����ؼhG3;�t���<Ŀ:=�ܠ=f�=o¦>��]?�W�>/��>J�7?$��n8�O����1/?�;=싂�J�����h!��>��j?��?�XZ?�yd>8�A�e	C��#>4�>f &>X6\>�]�>���\E�k�=�{>ұ>Z1�=��M�����	�������<= >=�>?A�>p����r">R�����w���Y>�X��Z��X+Q���E�>�-�[�h����>6�O?ZW?ˆ=�9������g�l)+?�;?�L?L�?H��=�۾͈<�E�G�,��}��>|ߓ<�:��q��������9���U;��|>��������a>���G�޾Gyn��5J�x9�#I=����V=d��!�վq����=S>�
���� ��͖��Q���J?��_=�_��ogT�Mߺ�`�>#�>H�>��<���k��o?�6j��7��=J�>G>>�`������	G�����G�>��X?��@?Cȅ?Z�V�nm�ٸ2��꾊���(dֽ{M?���>5��>�Z�>#�.>ލ�U�����QO\����>6�>q���+N���˾v���H����\>i�>��4>���>�Q?�S(?6>P?|�?��?�!�>�!ͽ ���'�?�7�?(^�����Bz��P���ھ�!�>�v�>�(��Sx>��O?W�P?�O?��d?O#K?�C>��W�������z>z�v>m36��ꢿ�'�=�1?�M�>�B? Af?C!;>a<6�������Cp>D�>@e'?���>�?iI�>��>�������=���>��d?�ރ? �p?�|�=��?�j,>���>�Ζ=�;�>h4�>�0?��O?@s?��I?hV�>�c�<�+���f����l�ANv�^
�;�?<�#t=;M��j������<-J�;
�j�VS�����Q�E祿)�X<��>
{>������->vþp?����<>�i��n��l��}�*��`�=�
�>ͧ?�ϛ>�>%�D�x=���>C�>�q���'?��?�?��H<�Sc�)�׾�!d��K�>U�F?&+�=��i��ߒ�8zu�:`h=$?n?*%^?�ym�D��ɍg?�O?ˀ'��Z���籾)��
��L<�?j/�>��A�`�?���?g��?A�?kż�(��ߩ�O��2*�_Ղ=�\�>������j@:>�2?�'>�U{>�k�=�3���'�W(\�4�!?�	�?�E�?�҆?y�>�g�=ɿ���L��/x[?�H�>XK��>� ?i����Ѿ�����ё���pê��Э�$5��tԨ�\n&�����X�ѽ���=��?��u?��o?�]?� ���c��M^�tE|���U�����>�zE�x�E��F�/�p����'<������9m=�1V�O�,��?>�%?��H���	?���]\ �y�����n>hq��4����p��j]��������<����j�K!F���?��>�7g>�1g?3�W��� �j�H����ս�� >� ?�pe>�h?���=
E�dU%�͆��D����Y>Q_v>��c?�&K?��n?����&1�vf���^!�ä1����-�C>o>�a�>��U�����%�M�=�	ms���62����	��=-;2?�~>�j�>�
�?��?�	�����+�w�001�sS�< *�>�h?�e�>C$�> �ѽ�W!�[|�>�vl?e�>�̟>͹��7�!�^|���˽1,�>�)�>̏�>8�n>��-� U\�4m���s��uF9�;��=�h?���`3a��ۅ>��Q?��ǹA:<v�>�]t�:l!���v�%��[>�o?�=��=>ž���@�{�A��O)?�`?�1���*��!>�"?��>�w�>v!�?\��>�fþ+ű9W�?��^?�PJ?k�A?ou�>΁=�T��k�Ƚ�#'���,=�{�>	�[>y�m=�k�=X���Z�y��("E=���=�zм���߲<�b��Ȫ?<��<�v4>�7׿=D�\�ؾ3�����ZI�:R��U�%�&�:�BE�����>��犊��)E�H�½��I��M$��r��P��W�?��?�[���ۖ�S���ݢv�Y	��:�>no���ý�R����,��q��3��d���08�X�{AO�X�5�@#?	����Ͽ�ed���ѧ�#,%?�E�>�fy?�����-Y\�D�>�q��$�Q����<�� vп ���l?t�?��ݾ4���&�>�S�>w�z>��5>�v�_����u`=�e�>�2?���>���-ϿV����M�����?�r@O{A?t�(�����GV=���>�	?��?>uR1��H�����;U�>�<�?e��?�M=��W��u	�}e?�l�;��F�_�ݻ\�=B2�=V�=��y�J>W�>��HKA��*ܽ٪4>N݅>!"�����y^�|b�<��]>��սQc��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=w6�Չ��{���&V�|��=[��>c�>,������O��I��U��=����&��8P�tD$��^=tK�aq��W���2<{��
n����H������;ďs=��a>nܙ>��E>T�m>�l^?Oa�?x��>,ټ��_���ns��� <(G�'�6�?㮾Y�������^�e����� ��nh�P7=��I�=gQ����&j!�8�b��'H�P�,?��&>_zǾ0�J���'<s�˾՝��zD���Z��t�̾y�/��k����?L�=?iY��T	U�*��F�ҼY����X?sJ	����Z$��N��=
����&=L\�>_U�=u����/��,R���0?�?w���M���L)>�}�2S=J�,?�� ?*S(<K:�>G�%?}�"�G�ٽ�.`>�I1>z3�>���>��>�1���e׽:�?��T?����%˞�yX�>�¾�4}���=�7>
�3��/㼈�W>Bi�<�/���_%�k󠽨#�<<2W?ͩ�>��)�tH�x#��S*'���B=T
y?�@?���>\pk?�"C?.?�<T��ΔS����u�j=��W?�*i?��>�R��j�оާ���5?>�e?w?P>��d�3��Z�/��/�!s?��o?:�?����!}�����&�5?OP?F_^�ӑ��ҾJx��l�s>J�?��>Xx"�M?��??�������Բ�wK�� �?֭�?)��?�Ѿ=㞽��=1�!?5��>o;�����нJJ��?55>�R�>���}a�������Kо�'?gt?��>tߧ�
�/����=�ؕ��^�?c�?=�����m<���Gl�Ǖ���Q�<�ګ=���u"�v�7�6�ƾ
�
���������Ȇ>�L@N���k�>Q�8�P+��VϿ�񅿋4о�%q�O�?Kj�>�ǽb���şj�Mu��G��H��i��aj�>_�>	*���N���{�iy;�P%�����>r��1G�>��Q�Ǭ���ȟ�0H<���>���>8�>2(��`���ؙ?�����ο
x���C���X?K�?��?�?eU9<��w�h�y���!�tG?�'s?6�Y?+�%�C�Z��5�isr?�Fƾ��d��+��F����>�F6?�u�>�b1���G>Ô�=��>l㸼�#%�ƿ��즿�ԍ�x<�?��?�=վ�;�>���?�&?�C��*���~��..����=C+??=z�>��F��һ>�CRk���?{4?�.��M6�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�W�>�6�?)'���?D/�>���u ;��P>�f���<��
?��c?��?4��>X�0>� �j:$��-��xr���#0����>�Y?�aC?_�>V�h<w�Q K������MD� ���M�P���Ծ��^걼 �4>�Μ>w��֥��)7?]�)��տ����٤I��z`?�^9>ޕ?e�B�6J�����SJ?��F��;ػ�|���(�6��?�	�?}�
?8ž
�<��>�dҹ�(�>RKX>�:Ƽ(�J>|wZ?��7=�f��-U���>���?iF@��~?��=��	?J$��P��VY~�H����6�R�=��7?%;�"{>���>.V�=�tv�"�����s�̨�>�C�?Iw�?\��>P�l?Suo���B��S2=�:�>�|k?�r?Hx�z����B>-�?c��[����O�3f?��
@]q@=�^?u��ֿ�؝����_��x �;K�>��>7_��ɚ=۝�����<?�Z=��!>��>
�_>E�9>�X>->.Ű=[A��]�(��O��r���~�W���,�S�H�(`������fg��eվv���K�9d�F尿c�9���c��=нe_�=�sX?��M?\�o?U�?�����>������<�S!�]/�=Ȭ�>�2?M?�,?���=󠙾g�h�(b��Bp��o����k�>��F>���>��>��>����FP>1>�B{>�)�=�5�<v` ����<�eR>#��>���>"G�>C<>h�>/ϴ��1��j�h�Jw�W̽�?G����J��1��[9��Ŧ��h�=0b.?�{>����>пO����2H?N����)�E�+���>��0?�cW?Y�>G����T�:9>п�"�j�v`>�+ ��l���)��&Q>�l?ޖf>	2u>��3��g8��P�T���m|>:&6?ȶ�JE9�-�u���H�7aݾb.M>���>[�D�@l������ �shi��'{=�t:?�?t��.ాX�u�g?���tR>%o\>�=hN�=�UM>`�b��Bƽ4�G�؂.=ܟ�=�m^>��?(�)>ݵ�=�W�>U���82R�^۩>�B>�,>]D@?��%?�Q�\ޛ��!��=�/�^'x>��>��>�>�5K�*��=[��>Ib>�p�%冽�W��>���X>q�u��^�jv���{=F��c��=��=�7 ��=��."=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ_��>��4�uX��Jz���T��x�=[�m>��I?˵�Q<�X�����>���>��⾛���o�ʿ7~���?D��?��?fc�Bb��:�_��>���?;9U?~+F>d뾔�D�/�f>f1?.7@?���>�(��CF���	?F��?���?�X>]&�?g@d?+��>,��]l4�9շ����;��=�ӕ���m>���=��̾��L��ғ���5(m�5,� <�>L�R=˞�>0½��щ7=�ѱ�����-�(�+|�>��>�r>��>���>A�>���>o�*=�v��!��=���=�8?B��?l���mQ�"h�J������>�X?4�����!��>�De?~��?"��?�9�>$r;�\���#��"���GN=���>���>��>;� ���M;w��1�~>?y�>>>����5r�(NƾTl񼱍�>��?52�>��D>��*?7^?K�,>,?{�>�η��|!@��s
?�Ʀ>͎�>��?���>|�Ⱦ�z0��Xv� ��8��4�b>tWx?o?jW�>S���A���M/>%G��*�>Ƥ?nyE?���/�>!ó?WXX?g?�\�>�ɾ���^<�=��=�!?�&���A�g<&����M?tP?��>1��?ֽsּQ������!?;\?�P&?W��	Ha�+bþ:��<��>�Z���;"I�|�>�Z>�������=#>�C�=�m�k6�upj<�A�=�p�>��=a�6������3?!�Ͻe%��0R>5���F���>�l>�߈�'w�?`BZ=�̆�"���?���!뎾2Ju?�%�?wl�?�6n��wi��LE?�(�?l�>SG?$�)�F�ܾ.�qѕ�~��0�6�w�%=���>�=�<����̩�^A��4ǂ�p�<�k���>��#?��>�4�>cB�>u;�>�:������mg��4D�"����B5��i�b>����&�A�=����YN��¾J�`��u�>lO�u��>]��>�X@>�>[�>&�߽s��>f&o>���= �>yU�<E��>�I#>_��#�\��QS?j���/�%쾃ͯ�D�7?Va[?m-?�|e�����p�T$?��?�z�?CF�> Vg��^0�'U?�k�>_2�9�?Zn[=��ۻ��<ݙþd������;���>����3�x�@��g���?![?�"�;�㾼4Ͻ}����]=k��?��1?��.�˒*������D�#>I������}:�V���r��:|�5E��[9x�Uփ����5Dd>�2?6��?������1����
}��dU��!�>�t�>�p�>�[�>�O>!�����!��4�*3��.��y��>bZ? XI>y49?8b?��?��d?Q.�>\�>#�����(?�P)�}D>��>]c+?H�?9&?�<<?�=??	�e>�����-쾮��On?��?J0?o�?�2?׿������`�/�R��;vw��s|׸��A=�G���A��䛽@ؤ=�P�>�Z?��R�8�4���>�j>�}7?�z�>���>K��B;�����<��>��
?EN�>�����}r��e�T�>)��?Y��=��)>���=�o��WEۺ�M�=�s¼V�=�����k;��q<j��=�=dp�n-�Ҹ�:s��;L�<9�>��?X�>��>�:���b ����7�=c�X>�[S>��>��پ`����&����g��,y>�\�?�^�?�Lf=CP�=Ӵ�=E��Y���!�������`�<?��"?�T?&��?o�=?�{#?1g>�
�M,���k��ue����?�),?P��>{�:�ʾڨ�C�3�M�?l�?"a�
����(��¾�ҽK>/��~�o���9D�R������阽��?���?��>���6��N�Z֘�����1�C?��>*R�>m��>&�)�	�g������;>R��>N�Q?��>s{T?�3p?P�Y?{V>�n<�������������>�R>?�-�?v��?0ey?���>��6>�K��?�����)������������<5�L>gx�>�q�>d�>
��=��$ȽҀ��>�m>��>$ط>��>Yut>�	����G?���>�J��^M��O�������<�g�t?���? +?=d��vyE�a���$��>I��?�߫?��)?V�U����=�M뼍��1Aq�w��>9�>��>��=��7=�,>G��>��>X�:�|�8�sHN��=?i�F?H��=������]�%�r�H{��'m.����ǉ��_-ý$J"���=n����V績2���W���Ң��þ�ᓾ�*?�6<?�0'<�=��=�e��"��O3=���=J˱�&#�=6s�� �n=�x�e�<�?<+G�<�L�;�e
=�7��R�˾3�}?r;I?Δ+?z�C?<�y>�>>x�3�^��>���@>?�"V>�P�^��Au;�ӣ�����M�ؾ}|׾~�c�V͟�H>�VI�ϵ>93>*I�=��<� �=��r=�Ŏ=0�Q�{=Z;�=�G�=�h�=:��=�>dE>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>X`7>�j>_�R�h�1�^�\�1c�}�Z��!?%-;��D̾��>�N�=�߾��ƾ��-=�i6>
a=���=\�p�=�V{���;=͈k=��>̫C>o�=ׯ���=��K=(�=��O>O���m6��[*�ϻ4=���=	\b>3l%>���>��?^0?4Zd?�8�>�n�LϾ+=��`F�>���=�G�>���=�nB>���>��7?�D?��K?q�>ᓉ=��>L�>D�,���m�|w�.ɧ����<���?9͆?�ȸ>��Q<w�A����c>��4Žw?mR1?�g?՞>H��8�߿a���?���i�=v8�<�9-��D�� e�� 1�����^	��z�=�K�>���>5��>���>-�=��=�@�>�5P>�
�ۣ�=�<1>�[���=.f�=ć�=w���Q��9`�{�޽��0�q"��S�=7a==��=���=:�>A�>�Æ>Ζ�>x�������>�k��AM�Ad�>�ྗe�zDY�O�����(����<
>�r�>�(�<}я�J�?�,�>�q�=���?�{?~U�=/lv����0鞿yH���nn��P=��X='3U��"?��c��b�g潾���>�Ď>�[�>Xl>��+���>��gw=��k5�JG�>���n:"�!��q[q�0��*��h��O���D?�?����=~?�qI?KЏ?T��>䪘�ޔؾ/e0>������=\��P�q��F��|�?�'?���>�:�f�D��*㾧������>44q��BQ�U����B���;�x��"$�>uh��C�žF!2�����|w��K?������>˝A?���?͔��2Nt��7����>�F}?�Cc?\��>Z|?U?@�U�|Ⱦ�96��Yd>dEg?�*�?
S�?���:�$�=���PQ�>��?^�?q�?YXt?�I��)�>�铻��>�����=��>��=Z+�=��?�	?�?쟽c�����(�ﾺ�P��=���=��>�I�>�q>��=�8i=Uj�=	�d>�J�>�k�>�R[>�H�>܋>���J�
�})(?��=���>> 2?�8�>�@=3"����<�PY�9�?�\�+�����8��G��<Ҫ:�1W=���,��>8kǿ��?uQ>��f�?�D�#�.�Q=H>VaR>�׽���>	oG>W>J�>�z�>>�ш>
�)>mؾ��J�<���0��r;��2�sn��,��>����Y��� � ��W���վ#g��zZ�5fv����`L�=��?/��~La��&/�g��=�g/?*#v>�GX?���ʋa���j���>`x�=/���JF�����U~�&�?���?�5c>��>��W?��?ԕ1�� 3�IoZ���u�%A���d�'�`�V㍿����j�
��5���_?��x?�wA?��<�-z>ݟ�?�%��ˏ��&�>�/��#;�$<=�'�>X,����`���Ӿ/�þF&��3F>A�o?�!�?\S?�RV�' �m5a=�Y?kU?�ǜ?pgv?8b�?]����9?4_�=�1?�ę>s�=?>�5?�C?>Z�>F`j>�K_<Tz���K��]���tE`�-�=p�X�<�b=�q�=|����:B�>��=~8�3�H<��o>Wu�=���6�X��6=.9�>K��>q�]?���>��>�M7?Y|���5�񄱾<i2?��"=�ǂ�G���:8��h ��>�ol?}��?��X?�1W>/C�l�Q�6W(>���>�a->	zj>}��>iD���\Y��g=�>Z">��=pD���冾��	�����=h#>ڗ�>��>�C����>1������o�=>$x������2J��$:�zm1�2�:��v�>��R?U9?uo >2a��=A�:'^����>p�U?��D?��|?/^3>����!<�X�S�]#c��{�>Y�=Ip ����������a$����=���>Y(��߮���O7>����ؾ��l�o2D�]�پ�=�����=� �
�[���k�>ў8>쐡���06���X��8�L?�t�=�&����_��ߪ�^��=s��>�>M[��3a���:��$����x=���>��O>���t]�mF���My>�J?B`?2��?68m�Ps���;�%w��L��]���B?�h�>�?1@>�kN=��ľ�����e��7J��=�>0z�>����G�搣���a��^��>@8?�>�M?.M?��
?�"c?̖,?0�?��>�����о�%?�.�?�x=P�Խ�M�1�7�-�H����>ڠ'?R,B��>q�?��?ft&?�R?I,?�>-��ո>�_ϖ>5�>Z�W������_>��I?Ub�>|X?㷃?Ə6>rH5�Ş�������=�9>�1?��!?��?��>��>������=��>�c?	1�?Q�o? ~�=�?�A2>��>  �=ϐ�>[��>�?6VO?"�s?*�J?���>�<���]2��Ss�(�O��ˀ;	tH<��y=f��h�s��@�Z��<9?�;���Y���D��p��~v�;�f	?X�I>�����'>*@ξ�|��wUG>~�`���ٽ������Ք�=!>>���>@��>�^���=ʧp>N,�>�B��? ��>��!?��=�[�t���#.���=>q�X?��z>��T�G���笃���껯Zn?�c?x�4�O�b?��]?Nh��=���þK�b����r�O?B�
?d�G���>��~?k�q?k��>��e� :n�'��Db���j�vѶ=<r�>LX�J�d�n?�>x�7?�N�>	�b>�%�=ou۾�w��q��n?��?�?���?�**>k�n�N4࿋U��V�����]?X��>���(�"?*��r�Ͼq����`����ᾟ���©���9���%���f$��߂�B�׽�n�=,^?:�r?�p?��_?KV ��:d���]�r��h�V�J��-�H�E���D���C���n�k,�����������F=������H�ew�?��?��c���>GC��}�����꾮dT>W`����j�3��<H�����=,��=�k_���������+?�`�>$S�>�,?ͧM��l;�SV�3q/��qݾ.H>s �>�Ji>�p�>�i =���I�T��jӾ�!���+��q>��d?�K?Gp?�c����1�ד��/%#��*�����K>�>�V�>�vU���"�4�'��?���r�+�d$���s�m��=:�0?f�}>�>�}�?kE?�`�*���~v���0��J�<�&�>�"i?j��>�K�>8ν�"�P�>>�?;e�>��?o�h=7uF�A�/$��[��>ͥ>��>	�>_���V����mږ��I�״=)�7?����Ƶ$��^{>"�D?�ʫ�,���C�>����F$Ӿ+־k��=vw}>�&?gn=T����1�?�F~s�Vh����?!�?(R����(�!�>�z?�u>���>�p_?���>�)۾g������>Q�C?�;N?�2P?�0�>T)��\�ν�OȽ�c=iV�>�ɬ>m��=㔽zC�a���9n�a��=Fm+>a�=�:��m�6=��q���;=����6�_>kۿ�CK�:�پ=
��3?
��∾����Yh��Q��F\��5��1`x�����&��V�6c�d�����l�n��?J<�?����r2��鰚���������%��>��q�|�������)��������Ib!�K�O�c%i���e�I�'?$�����ǿ�����۾�. ?
 ?V�y?���[�"��8��� >���<���MA�܄��v�ο�����_?=��>�G�]夽���> E�>�\Y>͚r>�B��GI���E�<��?��-?���>�q�ۂɿT���f�<:��?��@nA?��(�P�쾔8V=r��>ߒ	?��?>�R1��?�6���fO�>�9�?���?L�M=��W�V�	�n|e?y<��F��M޻�9�= Q�=ڤ=;��]rJ>"X�>�}�YfA�Uܽ[�4>Hم>֯"������^��c�<|]>��ս�g��c̈́?�l\�If���/�!Q��>*>V�T?c5�>���=p�,?$0H��xϿ@�\��a?%�?'��?K�(?"¿�?��>-�ܾ �M?56?=ؘ>�N&��t����=w[޼mɡ���p2V�sN�=���>�4>Y�,��s�kO�����ca�=L��ƿ͇$�և�Rl�<\c�J|_�B1潒ݬ��R�2���p���꽼�]=���=�eP>�C�>�YY>�X>��V?�bk?�ӿ>f>��ὣĈ��;��$����h�V����_�/d��+;�%߾�~	����Ȟ�\�ɾ�==�D�=$�Q�Dk��� �s�b���F���.?.� >ɾ�jM��<�yʾ~���"���̣�ͥɾޅ0��m����?�A?�����V��U�c���켽��V?l�����!���2��=X��K�=��>军=�⾢�2���R�~r3?�?U����n/>Oҥ���<�&?�?X�(=m�>�?O9B���ٽ�xf>�8>�)�>�H�>��>e���݇��A?�JV?�R��^ۮ��Q�>`5������s�=
�>��$�g�a`2>�����ċ��`
��'�8��;%W?̝�>��)���G=��܊� <=�x?e�?��>�dk?r�B?V�<�I����S���]#w=��W?;)i?V�>ꯁ��оSx��'�5?��e?k�N>�Yh���龹�.��T��*?v�n?�a?�����s}�9������r6?U�\?��d��	��a,�;ڒ�g"Z>E��>���>�05�FM�>VB?|�!�Z���qg¿l�3� L�?�+@���?V�<�U��"�=�w?,�>,(����uo���'���S<7�?�A۾���&��u�1�a9(?eu?~?`����꾺��=[����H�?��?����I S<�����k�\i��V�<d�=\���"�#��8��9Ǿ��
��\������^�>];@Š潪!�>*�7�|8���οl����Ͼ�_r���?�s�>ڌƽ䊣���j�2vu��G���H�*?���>C���S>��:�!`x�����~|����>��#��>(���}��̾R�u=^,�>��?��>�3�=I�Ⱦ�O�?' ��\���Ζ�A'��80?iB�?gqE?�a
?�hG>(s0�	)��$8 �#�n?쑛?�Wn?�V��
ξ�+$< �j?l_��pU`�܎4�aHE��U>�"3?�B�>K�-�ٲ|=�>���>�f>�#/�n�Ŀ�ٶ����P��?މ�?�o�-��>t��?vs+?zi�8���[����*�b�+��<A?�2>����8�!�=0=�sҒ���
?C~0?�z�`.�t�Q?��� �y��M��fY>���> �	��_I>���s(���g�7�f����<�o�?7�?��?1�:�rX�qbB?���>us�����=�:�4^>g��>�?��t9?
r1�)�/z�>���?�_�?���>����y򗿡��=a��?R��>�L�?��[>��?#>S2˾���<�伱�>t���0�?��\?"m?%=�=�C���/K���Z���T�J#�O�<�=J�>�#\?�>&?�Z$>�zw��ǀ��$�.ve��&���\��@7��ds<4$ּ�Oh>ƌ^>�>���������?Mp�9�ؿ j��#p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>D�Խ����\�����7>1�B?[��D��u�o�y�>���?
�@�ծ?ji����>x	��ۂ�"Xx��b��AX��->��.?� �uub>�k?c/�=��r�_����l�Wd�>�X�?�Q�?���>��?}����P��}^��$>3�?���>e�=X��#��>��>�3�l���T$�rSE?T�@6B@�@l?	���������o3��e*��u��=���=#G>
��]U�=� 
=�l�=�b=�7'>P�> �3>��L>�'6>CU>)�>�T|��p ����tY��;�R���"�Ѳ �7��M0���e�������Ⱦ���JW���t��;�a˽����;��M�=\�Z? �T?C'r?  ?kљ�Ʊ>\��O�=Kc)��[�=�Ƒ>�5?�K?��"?�K$=,|����d�x��u<���a�����>�(<>u�>t��>p��>;޻'N>	L>��j>��=�U=��:N=�MU>�"�>���>Ȋ�>�O=>��>l����,�d�:s�����^�?��J��앿?.���f����=�\/?�>�*��@*п��'�H?笔�G����+�ֽ>�0?<yW?e>:᪾C|��>����4Xe�8>�4����q��M)�h�J>ʆ?_3h>1]|>^/3��%=�LIC���=�*>�<?8v���%���3x�>)K�K)ؾ7w9>k!�>,N�=�������a�t���g����=�)?�m?U��:C��{���ap��'0>�^(>��1=nX�=5�>I�y�д��51@��c_=�~Z=�y>E?��0>�1=	��>%����]J��Ƨ>�C>
($>a9A?��?`�*����%.��r�$�D�z>���>��}>
�>�N����=�F�>P9f>MC�4蓽��jo5���K>����a�i�V�H	�=�l���$�=�L�=4�s4��)=7΂?�����~����ZB��|�]?�B? �`>"Ac>I�I�ʨ�X�P�}��?x�	@��?���c�`����>9ڕ?&��F�@E�>��>��'���k�2?�Ⱦ�Ͻ�Z��z�����?���?� ;�Jx���Q���=æN?�%��yh�>Ux��Z�����e�u�[�#=)��>9H?AV��R�O��>��v
??`^�������ȿ0|v�l��>W�?���?v�m��A���@�.��>:��?�gY?�ni>Ig۾q`Z�t��>л@?�R?5�>�9���'�X�? ߶?ͯ�?ҧ�=�<�?5j?1+/?�>M�D�`��5��{=U/�<���>���>��3��"8��������j��{�=�k�����>�*��[)��X��`��<So����Ou�>Y��>SG�>���>gT?c��>O�>�v�<Qbl�!i��w�۾O�K?O��?���&n����<P�=�g_�*@?�'4?�"S���Ͼz��>�\?���?[[?ԟ�>7��S4��տ��o�����<i�K>BV�>Հ�>h�5�J>ˢԾ8�D�L�>�>����پ<��z��U�>�\!?�=�>�>�=�� ?��#?��j>D)�>�`E��9����E���>x��>�H?��~?��?\Թ��Z3�����桿��[�4;N>g�x?�U?Fʕ>A��������pE�cCI�������?}tg?�S�t?+2�?ۉ??�A?#(f>z��ؾy���1�>�&?����v2��@=�#Y�֑�>SC�>��>ʽ��>W��X�3��`�|��>��`?W_B?�ھ�9��;⾀�<ȗ>2y�	c�p�G=���>S�r�Y��=�&�=y�D>�"ｂ�̽�gd��8��]���Л>��=|�F�'Ԝ=�R ?����qu���<�Ls��V�Y�g>�Nz>-�վR�a?�l�C�o������9��~ю�g��?�F�?���?ac����n�;b3?��?O�>z�>H�����>�˾C쏾� H�W�-��a��&�>��a��/椿xY��
Oz�6����2��>E�>D�?~(?�6>���>X����&�ډ�q}�ٱX�Y���<9���0�^��Fw�����'�F�¾��q���>�k��y�>7h?�+h>B�c>��>ix����>.�T>���>N�>7@>�W>2��=�u:LJ��p?9_��x_���4������x?$�S?o�b>�,�>Kɟ��@��?�߉?��?
�>i35��.���>*,^?j�Ž	S�>�'>~�"�|=��8����Z� ������>��)>��D��q��W��ZK�>���>�Η>9�ھKx�a����io=	M�?��(?p�)��Q�A�o���W�FS�j���-h�vb����$�[�p�f폿�_��!%��[�(�i_*=��*?��?�����!���$k�v?�Hf>2�>g�>D�>�{I>��	�>�1��^�"Q'�;ʃ��E�>R{?���>��I?��;?�sP?�xL?��>�H�>���6�>�g�;�Ԡ>���>��9?0�-? 0?#e?Wj+?-c>y�������Yؾ�!?�?�[?��?��?�ᅾb�ý�����5c��oy������-�=�8�<�ؽ,hv��=T=��S>�X?�����8�t���@k>W�7?"~�>@��>���<,����<��>�
?�F�>�  �5}r��b��U�>Z��?���ք=0�)>���=ǁ����Һ�U�=r�����=�>��\x;�v{<f��=
��=�-t����R�:�n�;�y�<�p�>+�?���>YO�>�)��;� �\��'K�=�X>-S>z>�:پ={���"����g�>y>�s�?Vw�?��f=u�=���=�j���I��S�����h��<�?�H#?oJT?���?K�=?&l#? �>w0�fN���`��;���?S!,?���>b��P�ʾ*�}�3���?
[?\<a�����;)��¾��Խ�>�[/�-/~�K���D�~������]{��C��?Ͽ�?5
A���6��w辗����[����C?�!�>Y�>��>��)���g��%��/;>���>�R?q��>T�P?CW{?�C\?�mU>��8����������)���">�@?�ׁ?:��?)�x?�>�>I!>��-���ྶ���$���0���(L='X>ㅒ>	Q�>Y�>��=}νtE���?����=Skd>y)�>&��><��>Ww>��<MB?��>IC��t��Φ���Ӆ���;�h?9t�?��3?o��<�`$�a�P�c�Ҿ���>f�?Ξ?�
?`F��V�=�I0=;پZ�����>��>Sf>��(>^e�=�AE>]��>:��>&�
�:��d�7�@�強�
?3;?n��=�ҿ�bp�����w��Q�ǽ"/ؾ~����g������=U\��Wn���Vо�~�� �CZ����܍�=p���I�>6%Ƽ�a�>d[�>4>",>��G=1%������@�i�L׼EE<=�2>��=�BW=����J3=�ܼ@>־W�?KmQ?|n4?1�>?Z�A>��>4�k�>/g��� ?�{�>��<1n��\�e�&>˾���ʶ�k����+n����a�>�؏�Yv
>��*>.�=X㒻.j�=�����<H���.�=N��=	n�=t�=�H�=�� >�W
>U"w?����;���2(Q�e��¬:?�5�>p6�=֢ƾ4@?h�>>&7�������K�X.?���?�H�?��?�~i�Ґ�>f��������=r眽%2>�j�=�3����>�	K>\j�iN���ĳ�#6�?��@آ??_狿�Ͽ?/>�2.>&�*>��J�.�$��_��o�g.�>'=?�;��f���3>��;�믾>����,>�2�>w��=	�p�vqD�9��=�
���,�����=Ԭ�>��1>���dF���=^������=�b�>D�=�X:��V <�A�����=DΗ=��>�S�>��>�-?�E?.��>�{������?���(C> z)>���>�����=Y�>1H?9vP?|O4?�k�>s
��{�>(�>:*E��r�nx���K���d�<��?�K�?J��>(좽��׽^#�[>�_�ɽ�??R0?w7 ?��y>�U����Y&���.�扙��>��+=`mr��RU�����{m�5��x�=p�>��>��>�Ty>��9>]�N>-�>�>�;�<�q�=!Ռ��µ<C���C��=e�����<wż����	k&���+�ō����;?��;o�]<w��;��=���>+ >n�>���=v���v�> �n��J��80>lt���'���\��:���+2��/[���>���>)���P��P^?��>�ZH>�?F�8?�u>�?&�&6Ǿ	J��n/h�P�J���">f�=�M��+`P��\��G&��8߾���>�0�>	�>MJm>N�+�;?��x=�⾑Z5�R��>?���8[�V��-q�25���퟿��h�G�Z�D?=�� A�=�A~?J�I?��?���>�!��W�ؾ%0>\���KL=����dp�~��ĳ?a�&?M!�>B�뾡�D��۾v���T�>�."���I��я�eC,�@_O�G�ƾy��>�����оL�,��'����[o8���<�3D�>�>?[A�?Ѕ����� L�R��0�d�Z��>��h?3��>��?]v?��k����y��w>�|?x��?w-�?* >�C=d
��� �>(�?*{�?�+�?k�t?��_����>/�p��W>� ;;�1>�j->�E==��=��?�?t�?�G��/	���羝� ��'U�xm�=��=�>�ח>:Ə>ӯ�=���=,T�=�H>��>\�>Uo>��>�u|>�%�}�
�T@?�+>�[�>>�)?Ͱ|>R荼Z7��S9�A/=�#����@��g����<�m̼
�=B>�ͽ~�?lU��v��?<f&>�O���% ?�	羵��=Ü5>��>��R��>�7>��_>Q(�>���>X�N>6'�>��	>|?Ӿx�>���!c!�+%C��~R���Ѿ��z>���?&�B���k��r1I�7f���a�Gj��,��l?=�hL�<�G�?����Z�k��)�C���.�?Ff�>t6?9ˌ�+��̧>���>8ˍ>J>������bȍ��iι�?B��?bSc>X��>~�W?�g?$2� 3�hZ��u��'A��d�Xd`�����~���IO
��g��*�_?B�x?PA?q1�<��z>?�$&�x#��|J�>�/���:�U�@=��>�a�'<Ӿ�þp��!F>|bo?��?�<?��V������9*>�F?&Z%?�8t?)K=?�8?Ur��;1?�B1>�V?%o&?*BF?>`1?�?�>"H�=�M�=� �<��<gH��%���Y�Y�G%���H���=[�<�5�<Q�:�я=���;T�<0�|������7ɧ�תa=�I�=O8�=�m�>i�\?Ks�>0ȃ>��8?���?�;������y+?2yW=j���Ҍ�-I��tﾴ>wk?�i�?�U?n�_>�a?���A�Fp>���>d]0>��X>i�>�޽��L��'\=1�>@U >ǵ=2�<���{�&�	�TN��$zM<�h&>PH?�J�>��<�l�R>Oa�� +ͽ$�x>ɾM��u�(s���%�����ľ�z>v'?c�>�^?>�S�r�m=�l��X@?� ?J�:?�_o?�HJ�����k�J��Ƌ��n�=���ܾЯ���ӧ�8�9��	Ǽ� ?�ZM��J\�E�$>��
����0����_��[Ҿd��=q	��/I�!3�����s]�y�>�$>e-��Թ��ꊿ��	H9?^�<�8ɾ�ߥ������s>�Խ>FO�>�-��Q9,�pSK�g�;��0>���>�yf>$�S��>�;�@�Ѵ�����>��D?��^?�E�?`��mzs��B�����k���pӼ��?�ѫ>�?��A>Ԃ�=����i����d���F��P�>�>�>ۃ�� H��Y��w��'($��g�>��?�>nL?��Q?��
?I^`?*?�>?�o�>����5���C&?g�?�T�=1�ս�W���9���E����>p)?�SD�팖>�#??�?�b&?Y�P?�r?)�>�0 �A�?�%v�>�,�>"�W�Qb��[�[>�kJ?� �>ĽX?Gg�?v�>>"�5�|飾G�����=Pk!>=�2?
�"?Y�?6��>@��>�������=z��>�c?t0�?��o?�v�=.�?m62>>��>H��=q��>Y��>�?�VO?F�s?��J?N��>U��<�3��11��Rs�;�O�ó�;դH<��y=���0t��F����<2U�;�@��/H��G����D�� ��--�;]��>8�>>c�n����=�g׾�Ո���>���¾�۴���l�U��=�y�>h?�P�>��=��ʠ<�>���>no�_|?).?�/	?���;�FI�rCX��^�>G�H?�u�=��v�����:���|���w?�Z_?y����Y�(�b?U�\?]�̮<��~ž�i�0u�
�O?�>
?{zJ�?
�>fj~?��p?f�>�De��Wm�l����aa�i�8e�=$�>�{���e���>��7?���>��a>m9�=M�ھ�(x�?ϡ��?�?��?'ӊ?a:+>�3n�A�߿0���~9��K;]?HF�>~b��5. ?���&̾�j��"����h�_Z��n���x��pu��^�'�섾+Dٽ>&�=G?ep?}�q?io_?P ����a���Z�۵}�Y�S����ҿ��rB�v
E��D��m�)�����+���hD=d�}�6s@�˖�?Az'?�..�C�>F�����e�;l @>���%���H�=����i�(=ͧF='�j��.�ū��i?�;�>N��>��;?�Q[���=��0�4�6�����3>�u�>��>���>��9��-��齣�Ⱦ?Մ�o�ӽh�u>,�c?��K?��n?�^���0�s3��i�!��4��2���nD>ʒ>貉>]�W��G�xj&�]y>�]�r���������	�3�=��2?�'�>���>./�?��?�	�����y�v�B.1��7u<l�>��h?T��>Ɇ>��ν
!�/��>�kv?�f�>�ϫ>C>�������e��J꽖 �>%�>���>�U�>��
��Z��}�������<�@}�=Csh?ł���-����>˛=?�xp��볻�:�>���O
��Ծ�H<�y>�=�r?�O�=��>U�;�F�c��IᄾO�)?�5?񘛾t�3�g�2>ǅ?�k�>���>��?��>�^���b���Z?o�c?N�V?R*B?���>+ݼ������M���?&=�?�>!6�>�{�=?�;=N���A��QA��|^=R�>CZ<�-����r��ʹ�7;�;�vC=�5I>�տuOG��������vL��"�E���{Y�S
�Q<ֽ������뽵�9����f����*�m�R��	o��.����?N��?��	�ϐ���N��2[��S�˾�mX>sS���x��B�r�G��)��Ĺؾ�������=#4��%8��*8�ޖ'?�̑���ǿ�����Cܾ� ?> ?t�y?����"�[�8��{ >���<�����p�̑��o�ο����k�^?F��>��K����>e�>��X>�q>������U�<��?y-?-��>z>r�&~ɿ}��ې�<���?��@Xt.?��Mn��{p>�?\h(?c$�>�餾H�H�*⾋�?���?c f?�
�erG�D;ֽ�+I?@��=#+8�@��"�>G�=��e=I3
��g>M�>�2��J�)��Y�k�>
{>�)�<=�(�i����x��J@>�,7�ٵ<�3�?B�K���^���@��N����=��M?�_�>,~>�"?F2(��ο��]�&�d?���?�?�v?&��P��>��̾6~>?�#?Q"�>=��)f����q*�'j�����O�YD>j��>�N�=�9�.��tU��饼��>[.��fſ̎0�r� �}
�=�0\���FM���G����<�0���XR�ԅ����=��= 3>�Hn>�H>!�Z>�8\?t�g?�^�>�g;>�v�����o��M61��&���_�K͌�Y���>������о��򾺎�3���þ�J>�1��<VCV��ą���xm���Y���+?�=>�qľ��E��_�=�>��`���.D����#���K"�\�U���?_�;?#�m�N�5�Ib�{!��`���-;?$���v�9���#V>��μ+q�<`�>���=��Ѿ��j�;�bu0?�9?�x��NX��5�)>�����=��+?��?%]T<�(�>�=%?�+�)���m[>��3>5��> ��>�e	>e⮾�۽�j?�BT?w]��Ҝ��>�I����z��`=��>�j5���[�[>���<ߴ���cR��k����<5�V?���>��)��&�.�����M��LH=�_w?_�?���>�f?˰@?���<���qQ��r	�ecn=M�T?g?X�>����D�Ӿ��4?pif?��S>��h�>���,�K���s?�p?��?sN�:�{�qǒ�����15?��v?�p^��r�������V��>�>lZ�>���>��9�Zg�>�>?
#�H��麿��Y4�C?#�@s��?��;<�B��=f:?X�>٪O�s@ƾ���󁵾)�q=T"�>�����ev����xO,���8?Ġ�?��>Ԕ��W��T�=[�C�"O�?'j�?PU�����=����OCh�7����#��=�0=>}˼�����B����
�`����<z�l>�x@Ǻ�����>ȁ�IڿV�ȿQ�r��ĕ�?;��;�>(Zq>K��<�����p�K�w�=�W���Y���i�7��>)P5>q=��X<����e�UL<�Pn<"I�>PS�=J�>�߮�n�ھ� ׾ݎL��k�> *?�c�>{������?�߼��4�����������1?w#�?��?��"?�!�>�Rq��pt��oἙE�?@��?�'F?�t�w=���@>��j?�]��4Q`�
�4��GE��U>� 3??�>^�-�]g|=�>��>}>	/���Ŀ�ض��������?���?n꾋��>���?q+?hh��6��\a����*���4�A=A?2>�����!�63=��Ԓ�Ŀ
?�}0?����+�6�]?��_��.u�WR9�^��>����E�^4I�aoC��sn�Η�(�2��?�?���?
f�?`�@��!��a$?Ǫ>�H��Ye˾?A5=���>��>q 2>����1�>��]n0����=J�?z
�?pG?�*���⨿M+>���?�*r>]�?��>��	?��J��q��p�$>ml
>IQ�==�M?jtI?x�?��,=d5��&[��Ej���q�o�b�8��>Ktu?�6?+=�b_���޽�׾�z���ʜ=�D=D�a��27��=�O�>;�>>�JP=µ�������?Mp�9�ؿ j��!p'��54?.��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>;�>�I�>A�Խ����\�����7>1�B?[��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ha~����7�K��=��7?�0���z>���>��=�nv�ۻ��W�s����>�B�?�{�?��>�l?��o�Z�B�!�1=.M�>��k?�s?�]o���_�B>��?%������ L��f?�
@~u@W�^?(�ѿ�˾�P����>�%��Z�=@H�u�1>�q�>G>J 0=�"�>�B�>�V�='Nv=3�=���>�I�<��w�kl.���Ƀ�|pE�w9�L�,�Fӽ�G���@����Mkɾԧ��,A̽}�齑�ս9;)���j<��ӽ�h�=3�U?��Q?��p?�p?6ih���">/���M=�<�@&���=`E�>|U1?e�K?9i*?=����c��I���d���-���)�>��L>��>�k�>`��>��й�`F>��<>�>��>!=<SR��=M>k�>w~�>��>��V>7��=��������S$q����ɀ����?�����K����F�������=��*?�h�=򰍿2&ʿ\줿��??�����@�^�=��>E>�w8?7O?im�=���`��m�= 7����]B>E��u�v�9�3���I>��?��j>�o>��3�f':��+R�	�����}>�5?/մ�ڈ<��t���H�J�ھ&�S>��>%}������V�{�\�f�|�n=��7?��?>����,��
�w�u鞾JR>W>��=�=WU>�'P�m���fhG�9�=���=d�c>N?sv>`�=�K�>㟾���L��>�'J>��#>Ax3?1w#?����i]������/�r�j>���>ن|>�c>��5��w�=��>�z5>-F��tGo�p3ؽJ�:�]}I>O�e��u��%��H_k=zb����>pS�=��Խ��9�i��<�#u?�/����s�M��,�;Ha?�?PL	>���=�}��/����z����?I@�w�?��%���V���?�˂?1^彎o�=X��>u?>#��(��?��=�ά��t��t:�Z��?w��?
D�=������"�>5%?��ʾuh�>�x�}Z�������u��#=Q��>�8H?�V��h�O��>��v
?�?4^򾧩��w�ȿ|v�T��>#�?���?\�m�A���@���>'��?kgY?�ni>ug۾�_Z�I��>v�@?�R?��>V9���'���?�޶?ί�?w�G>y�?�s?8��>Y�x��q-����]F���Hv=a9�:���>��>]���3?F�4�������j����CRc>vv=P��>]ܽݼ���=����6��Z�]���>�Mt>a�H>�;�>i�?��>� �>g_=�-��֟��L%����K?���?,���2n��K�<��=�^��&?�I4?�m[�H�Ͼhը>ź\?j?�[?5d�>3��R>��,迿(~���<�K>34�>�H�>�$��FK>��Ծ�4D�p�>�ϗ>p󣼉?ھ-���X��9B�>�e!?���>(Ӯ=@� ?�|#?��j>pb�>�&E�t/���E����>��>��?��~?�%?:���o=3������Ρ��d[��@N>��x?C?�ە>T�������h��!J�$���}�?�Pg?��{�?�͈?�{?? �A?u�e>�����׾E@�����>a�%?G��p8%���D����>{>1�8?`�?b>��K>$'>
�f�ǰ!�g7?Ӑ?��E?�ȹ��w�����^f.<oO&�$�-UT�bC����=���Po���=�\���>�󀾞�<�)>x�>'_S>#���y"���I>�7,?��D�nǃ�gp�=^�r�
jD��>�K>*���e�^?E�=���{��
���{���cU����?3��?Fk�?s���`�h�w=?��?4�?�>_!��wg޾"��#�w�5�x��Z�/�>��>�i�;��G���P���[G��d~Ž�Z��:@�>��0?��>�?�>X��>�9�>`��XC�Y�7��Z�4_����4�ҺS�q.������l!�p`�=Ɨ��dN,�|�>[�e�P��>r��>?E#>�$>�ô>�=<!�>Z��=���= s>���=w��=�]=My�S���K?Ӿ�.��6�7����N%?��[?jD�>+���98��p?�w?�I�?�D�?��>=�u��\5�d
?Z�?3A^���>6�>@��=?�|=���,��J�[�G��j>	����n1��4�3�,;�>$8*?�j��6ԫ�ǽ�=�ğ��$}=�p�?&)?��(���O���m��<W�HS�Ԩ#��e�~̞��$�ocp�������Z샿z�'���7=e�)?i��?������)����j�N�>��7g>���><f�>��>S1D> =�/�0���]��E'�����>��z?���>&xK?��:?��S?��P?)�>��>���Z�>��W��z�>h��>�2?��(?n�.?��?��'?�k>_G�������Ҿ		?��?�?��?M3?���Ź�! ��*�P<�a��R��c
W=/�<���rsV�Ј�=LPU>��!?^R�BO:�@����>�0?���>$_�>ZT ��U}��o����>��?�>�>�7��_�W�p�$��y�>���?�X��ߍ�=G�q>Z�=��b=��!>%��=V;z>nr�<$Je=ޣ=.�	>�+	>ݙ���K����.=E�3=���nW�>GX&?{|�>��>�K��9Ѿ����I[<�u>~b%>f{'>aⲾG+���w�� �o���_>B�?���?_K_<�+�=GZ>J���ZZؾ������/�<5Z�>�E?&�>?�p�?�>*?�Q?̋>����+���������?�,?u�>&����ʾ*꨿�t3�Ȓ?~Q?m=a���s>)�f�¾��Խ�>QT/�%~�����zD�G|����F���̝�?l��?x�?���6�'r�ʹ���@���C?��>FS�>���>K�)���g�$���:>t�>��Q?#��>w�O?�{?6�[?��U>�
8��ƭ�Qܙ��_���>V�@?>с?���?[�x?^9�>/�>/�)�8:߾�5��sf��2�F���Z=%�Y>��>���>$ɩ>��=ԴȽ�C��>�b��=!�a>���>KO�>!�>Y�x>^�<��C?n�>d��b����L������m��_e?C"�?�+?_���C2��TB�V���5�> &�?�!�?jy-?u���FD�=�r�I���csF����>p`�>!��>}
>ͨ�=�)>m]�>���>�+�{���g=��ж���?��U?\�a=�mƿ�*�������|���/>q����u�>�;=�K�>��ټQL<�c�&���[��������s��1�=<�?���=�M>A�<��<����<�&��x>�~��2l�FÞ��\�=ӈ��=Gd��l�<=�=-�3=G�;�I�<A�ƾ��}?�IL?��1?��E?9W�>6>f%���Co>���8?�l|>���m�����A�D簾�n��
0ξ3վߞc�B_�>���D�>8�3>�-�=nS�<��=y{l=Ɛ�=�Y<J�=��=���=VB�=;��=N�>F�>hSv?��}�R���̻N�4��T�7?���>R`�=���B?�d<>����wt���H	�T;�?�n�?I�?�r?C�t��)�>U���[M=ҩ��.>zz�='� ���>k�T>����d��N��@�?�W@��>?8����Ͽ��J>/^G>���='O��R/�C~������\��� ?b97��վ]{>d��=�iپ�b��n)=6�2>�WO=2��s�S�Oգ=�~��ٵ<�w<��s>"�U>z��=f#��]d�=��P=$r�=+�)>�Ir<\���iα�B�^=!�=�0S>�~><�>�0?��-?Q.c?2��>��n��Zо�ȾV�>OK�=���>K=�6/>���>(R4?d�H?��M?B�>&� =6$�>i�>'M)�~�e�Dy�\T��;�=��?�?T��>9�7��@�:1�%?����fK
?��7?+�?픋>����A��1-�/>�c9������<$���C(}�x�=��d�%����P>"�>+�>�_�>�E>��c>��V>uc�>� >�n��.�=OA=*|>��j�#� >��ջm��<�"�����L;F��+1�<2�=%���������="p�=�,�>P�">9O�>���=-R����*>�L;�`V���,=��q��3'��$d����2��/��q>7�}>�
��R��x��>��>ɪ=>��?�y?��i>c�e�������z�e@���8���	>��
�7�@�'�e��9�@
�����>��>O��>sn>�+�)�<���=<�M�5���>*ӊ��L������p�y4��u����i�At�lVD?ᇿS��=A�}?�H?i�?ڞ�>fז��U׾.1>:��<$=��=(p�%쒽�?�%?y�>_�U�D�  Ǿ��ʽP�>]�B�^L�銒��.�t8��E�>���$|̾܉1�U����%��QC��kw��v�>��O?�/�?�4O�l񀿞�L��V�l̍�$?6�`?�f�>��?��?s����0����=�Co?6I�?|J�?0 >{�=|,,<r1�>L�'?%�?�c�?�5�?|���M�`>�>ǽh��>? �=dI-=�z=fJ=��S=Tv ?�M?���>����F���ھN��_�{�Ƒ�<�8�=� �>ul�>��l>f�5<O��<>�&>Y1>�J/> �\>t>]>ҧ�>Z��>���31�"�)?�}�=D�>;>2?6u�>K�S=�ẽ+��<��b��@���'������t�E��<�&�T�<=�+��yL�>�Gƿ��?��V>6W��{?$�1�+��V>,�Y>�5Խz��>��<>�?n>m[�>�:�>f�>1��>��#>1�Ҿן>��6�I�4���X�˛��C>�����9���,$��j�<��������S;b���~�~�5�*=��?�n�__��s"���{��>��>62?�X���Ƚ�o">x3�>)i�>���+���~��ɕ���?��?�!o>�c�>,G?���>d*J���k9������8�V�#��=D�*�w�����s.�Ur�aif?��j?2��>�8a��;n>~[?��U�:�P��C> D@�����)=(�?GUj=�{�iL	�&�a����>���?�)�? ��>�8�r�m�y'>n�:?��1?"Nt?U�1?��;?�����$?�l3>�C?�o?M5?��.?^�
?,�1>2��=+b���(=�:��튾)�ѽ=tʽ�����3=9`{=	4׸U#<h�=�4�<Sz���ټ�K;C>����<�!:=��=��=y4�>�ZN?]�>?�	?^��K�CY����,?^��=���ؗ������7Y��M��n?9B�?�Y�?�ƾ���b��I�=GS>\S>r�e>�Є>V�#��ၾ�_\�6	�>e-Z>��$;���)t˾���3"#�Tt=���>���>�>�[B=tN�;���������=��Z�h����������+̾�<�>��>Wh;?��?��d�Uf>�)I�n:2?��W?fԁ?��?c2�>;B:�p%d��la�$���˲>��>������t���H�.��k(�>����؛��{`>�����߾��m�Y�K�7澥8a=����kI=���zgҾ�x�{�=� >k���~W�G��CF�� aH?�1K=����|+]�v��m>SF�>�ӯ>$2&�"u����@�(��F)�={	�>9q>>vJ��_�+�F�����{>.AM?�f?�-�?�n�֓p��r>�������� ���?��>YT
?v9>b�=��ux�R�o��F��+�>���>(l���K�������%�J��>:� ?��3>��?c�H?�l?��\?g/??�?�L�>�֒��U&?�g�?���=f_ս�T��O9�F�0�>�q)?C�B���>��?��?)�&?YWQ?��?>� �6	@�Jk�>ڊ>��W��W��cz^>��J?v'�>�Y?ν�?�D=>ܓ5�'������zB�=��>�2?W�"?�f?S��>}��>B�����=ƞ�>�c?�0�?�o?���=1�?s:2>=��>���=���>H��>�?LXO?<�s?��J?��>Q��<�7���8���Cs���O�^ɂ;�tH<��y=����2t��J�E��<S�;�f���H�����D� �����;�J�>�WF>�������=��;�u����A>��R�����~������14~=�X�>](?���>G;��=T��>�?����{/?f	?��"?7˯=�8c�L���3��4Ì>r�:?�n3>�c�k'��t����L���l?Ot\?�׈�#c����b?��]?���9*=��Lľ��d����^�O?t�
?�aH���>�~?L�q?F]�>7�d��m�fȜ�^�a�W_j��ܵ=i�>�F��e�X�>��7?ɐ�>��c>���="fܾ��w�D����A?��?�ӯ?6��?i&(>Ñn� �߿	񾎍��U�`?�H�>1;���R'?SS�+Ӿ����"���n��ӫ��騾f��D䦾�e-�t��M�ݽn�=�u?��q?0h?O�a?�l���G`�^e]��F��JIT��o7�a3F� �C���B��0i�H���������J=3J`�r=�;�?Jq'?�h"��r?�t����X���=�$>�y��P�g��=o�Q��J�<�Y�<�z��2�\V���?*L�>֨>�<C?E'V���3�˵0�/�?������:>,�>U5{>���>����@�V��g��G����ʽ}�B>�bv?��b?�q?���,31�v�u����g3�<(���,�s>���=`?�>� U���� �(���J��l��߹��Τ��i�~��=Ƽ?�~l>'nA>�g�?�C?V�����9��W.���"�hr�>Ko?�'?yv\>>�3����>�>y1p?���>��>0z_�7O�P9s�5�ݽ?�>�/�>�3�>*%�>u��Z�����o��K8��2>�2c?����zC��f�>RZL?f��sZ�<}p�>J�������xV+��=��?�J�=J3>#�Ⱦk��{l}�a,t��#?��>&����8���ļ�?_OB?��>DE�? a?;�۾�׉����>xdg?f?��?��>$�t<��%���6�<me>�Z>�Ţ=��=�檽��׽��A���.���> H=_ڽN�ֻ%� �E�U��	2=���>Q�ݿx�8�;;�#�x��1�������_��<O���1�ڽF��g�r�\��a�x�L�~�j��J��W���3�k��?*]�?/���� ���Q��Ӓ}�����)�>3�@��I�ٟ����<l��޾D ����$v7�R�R���P�'?����ǿ����	Qܾ% ?A< ? �y?����"��8��D!>b��<Pᖼ� 뾀{���οɜ���^?z��><�)�����>9��>kZY>�Nq>�)������Q�<��?�,?�>��p��Pɿ}t���U�<̰�?N�@�@?� �>��x]�=/*�>b�	?@O8>�C?�J �������>Ke�?��?�w=��X�(L�`?��<�D���c�.��=�[�=��B=J=�� ]>�N�>�2�}�J���v;.>;S�>p7��]��g9q�C��`>Sh���G��q��?.PN��T��&6��#��!��=�@^?te�>��>�6?��0���ѿ��j��d?L�?{��?R?�վV��>�Ҿ.z5?Ť9?u�{>gI&�M_Z�Qs>����iI=�I��5�d���/>8�?�N@>R"�:��	�� ;��R>�{�P���%m����"��=y<P聽qk���LW��>{���*�����q�=��=S� >��}>�TJ>	^>�}Z?W�r?�R�>�37=Ð$��7��}�վ�6�9h�k��85�����F����žc���ݾuo�U���&��@�,��>��[�8�|.�+;`�^�[��3?_#�=�^��6PR�&�>�mʾ�B�������뽉Ϭ������E�Ͼ?��5?����DQ'�����O��	��b�5?u�k=;H�9����29>g='=�;=�XR>]y)=�Ѿm:�b1�l88?zQ?B�	����EMM>�Ҿ�3��&?�E?�O���~>aK?$�B�����=`@>�>���>���=�O�[�Ժ?��D?N��U8;mΤ>�t��2�y���U=s�X>u���<��4�>�ɼ=b�n�=V��ҿ*���W?�?R>�n@��O+��w��p0�(A�=[�v?I�?^K.>}9?��>?���=�3þ!�&�V��!�)=�0?�HM?�#�=~V"�A<¾��Ǿ��?h~u?��>�����K��͙@��j��y�> vp?��,?��=fDe�9l��m,�(4?��v?�b^�l�����T�V��<�>�=�>ё�>J�9�iW�>Y�>?L>#��H�������a4�n?��@@��?�9<��␎=�1?OG�>éO��>ƾ����w����q=�>S���?`v�z���-,�܅8?|��?�~�>˨��ڝ�8��=���b\�?��?�e��	�o<F���l� A�����<,ū=pf���!����\�7�h�ƾR�
�\����\�����>S@�8�n<�>Q>8�w,��IϿ����\о�-q�Y�??P�>�ɽ�����j��u��G��H�����-��>>�F��6"��m�d�p�=���=��>T>���>��&���������Z�<i��>�<�>D&�>0v�������z?"���㩿�����2���?梚?�Ē?�'?su�=7#=mYt���,���f?�^�?c6?4ʗ�YF��Qs�=�j?`���S`��4�)GE���T>�3?�7�>$�-��4|=��>��>�s>�/���Ŀ�ֶ�9���_��?���?sf꾵��>���?&x+?]�6���i��H�*�4�3��:A?*2>+�����!��==�e䒾�
?�{0?K���0���V?�N���U���>�8���*�|>�jv=v	Ž���=�O���O������Ȉ�BH�?���?cv�?W�M���#��f#?�=�>�ы���K��B<��>?��>�i�>��s�JW�>"¾G J���I>�,�?�h�?V ?�9������ H>�҄?�>���?x��>��?�J�>��ڽ`��<�7�=[%*>��,��?��>?O*
?��=�����T���Q�%6]�-JԾ�+G�kܩ>	m^?Q�(?1Y�=IJ�����>��2�=�wf�L#=5���c荼�S��܅�>�F�>h�b��������	�?i�Q�ؿf���['�7&4?��>2�?f��`�t����E_?8��>Q2�<(���"��iD�c��?�?�?��?��׾�̼D>��>�/�>��Խ�'��5z����7>F�B?u/��:���o�p�>b��?��@�Ѯ?� i��	?���P��Ua~����7�\��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�O�B���1=7M�>̜k?�s?�Qo���i�B>��?"������L��f?�
@u@a�^?*��ʿ�L������*���)�<��6WD>lI���4�=)>�>���=5��>�>5[#>���=���=�-�>���=��u�JI*�:Đ�8j��L�x�d��|�ƾ��@�V���"��K������`嗾|2���+ҽK��K;��yZ�sF���=�zV?S?�o?�� ?{�����>���P�=�"$�A��=l^�>QA2?��K?�5*?���=�柾�f��2������BY�����>y�C>��>�;�>Ĝ�>WK�;i�E>LB>��|>M� >6:=��0��=iS>r	�>���>x/�>��H>"�>@���3���Si�c|�����fϢ?�Ր��L�ﴔ�����/��`@�=T�-?�Y>�菿K5ͿB����7C?�ɘ����03��y>I�5?H�X?�O'>�}��݊����>t+�/�O���>h�߽[o�&�,� P>��?شh>*�r>�2���8�	R�]����
�>�6?�a���H0�=�t���H�E޾.�Q>zD�>�+2���᜖��}�;�h�0v=/s:?�x?9o����l����pT>�f_>=� =F��=��S>�;Z��sŽ6CK��@=�p�=��b>&�?=�(>?�+=�֚>�x��B�z���>q�L>��5>��9?�O ?�����ֆ��?'�t�t>���>�^~>�>z�A�*��=���>ΘI>��h���P��j۽,*:��KY>3А��	i�c���H�= ����>@�=�2 �"B��EB=l?GΗ�翁���%�k��X?eh@?�ql>�/>�7N�
���ޙ�<	�?Q�@�m�?6  ��3k�ߥ$?|��?�2ؽn�	����>2@�>kc���5!�C�?�h��������o���D�?c��?�	^>�Q�`[j�U�r=0QF?����8��>9�h���+.��Mt�=C	�>�vH?"D�L�T��A�8�?�h?���y+��N*ȿ=u��M�>��?�r�?$�m�5�����;��E�>�9�?KwX?~�e>��־nZ�t�>>J??�5S?���>Z^��('���?�'�?��?II>գ�?o�s?Y��>]�_�Բ-����YZ��dq=4�2���>j�>uB���eF��������3Jj������`>z�=���>��ڽ����tv�=4L��t2���X�0�>_�q>IG>�ś>�^?i��>`И>b^=~���:���������K?H��?���x2n��R�<���=´^��&?�I4?�y[�;�Ͼ�֨>��\??#[?�c�>����=���翿�}����<��K>4�>�G�>�(��yGK>J�Ծr5D�p�>�З>C��}?ھ�,���0���B�>�e!?���>WЮ=�� ?��#?E�h>�u�>\E�%���F��>��>�	?�d~?fd?"i��F!3����ɡ�`[���M>m�x?1�?L�>�m��@����9�>GK�ڙ��nc�?�lg?g��P?��?��??�aA?��e>�>���׾P����>�r"?HC	��8�n�.��,��E��>�|?���>.Ի�I����<�,�]�Pf?��l?no%?�P�O�^�,�ƾ���<օ��4�����j�e���K^,>��t>�\:���=J�0><�g=\ǃ�Iq��e�=�#>�ˉ>D ��V67����=�;,?�F��ڃ�R�=:�r�tD��>fL>���:�^?v=���{�4��2y���U�� �?���?�h�?qQ����h�M=?]�?� ?A	�>�S��Po޾s�� w�j_x�^q���>��>�i�X�侸���L���+F���/ƽb��;l�?
�?��?Q+?U�>� >�P��]�#����9�����^�ؾ�|%�/5=���F�!�ξ�&�BwW=ꙹ�ؿ����?��@=�݇>?G3?�GJ>'p�>��	?��=�3G>䰛=!0�>Gי>���=ć�c%X�����п��J?ʙ۾n:0��Y�/#��D2?��t?0��>	`�G֋��10��?�]�?��?}��>1�k�܏2��k?��0?��<���?��<���<y�T=<=������8��	�_���>�|ݽ��C�d�V�z鐾�ì>��?q��=�ؿ� ��=������n=�M�?�(?��)���Q���o�V�W��S����7h�Ui����$��p��쏿�^���$��۠(���*=��*?��?Q��ߓ��$k�?��ef>��>�$�>0�>vvI>��	���1�^�M'�p����O�>�X{?ܗ�>;�I?Q<?܄P?��L?#�>�?�>En�����>魿;��>:�>��9?�-?��/?(?2E+?�c>���'����1ؾ?$�?zB?�7?m�?��Hký_w���i�bky�3�����=R8�<^ٽ t�PW=��S>߿?_��9����Id>\�5?�d�>��>�:��ꁅ��<y��>��?jÒ>������p�0��,��>�͂?6���j�<).>��=I������;��=�ἡS�=n����YH��':�:x�=�5�=g�K;Ҍ�����uV<܀�<E��>z�?��f>��>�e�X�����]�1��=��#>�;�=���`���F��f�i����>wҘ??��?��}�>kJ�=�ؐ�}ž���!վ`_=:?��-?��N? /�?��'?�9?^��>�ﺾ����z��������>g ,?�s�>B��1�ʾ��3�,�?O?#a�[��>)���¾$սX>!6/��~�L����	D���o�������U��?¸�?s]@���6��J�����;��(�C?8�>�{�>{��>��)���g��*�A�:>�k�>>�Q?�N�>��O?,�{?F�[?��T>O�7�h쭿����qv'�u: >r�??�g�?���?��x?X��>��>��*���߾��������~�lF��
�_=�GY>�̒>IH�>CW�>$��=�Nƽ��#C@� �=��a>jb�>~z�>�(�>�v>I[�<k	C?@��>����f��S��0���y��<�~g?��?�[1?�㬼ރ���D��h�`�>�?_E�?R?��!��� >Sݱ���ξ��W���>Ė>��3>D�=��=igZ<�W�>dy�>�p�����
8�7�<&�?0R@?�q�=l�ѿ�e������j�>4Y��<>L�F���>y����!?v��>ٓ�=���=�i���y��ž@�a�Ʋa�o�T�K��>��>" =�8��=�n�>�y>��F�U>�C^�rF��6�=��J>�:P���R<�r'=̥�=������=�޾W��?�~?%�?��N?�*>�ͩ=M�k=�B�> ��`�
?�:>����f�����_�9�Ծ�%*��ξn���뭾��4>��m�P>)Pl>-��=���= i�<'�>D^��k�<|�`�XR�="˿=sE>� >�19>�NP>)?v?t������|O���뽬.7?�T�>:\�=$�¾�W??�@>΄�[��Q��~?�8�?���?��?�Au����>tԤ�����Ubr=����!->�r�=_���ܻ>�XU>QR�uu��"꾽���?Rh@�v=?I�����ο,3>�ȁ>r�> �[��;#���+���̾¼��x�!?�a���ľ�7z>��S>S?������=<e7>�V�=�ϽSnG��j�=2���E�F=�FL=��>>v�>f[*>z�����=ޭc=v�=�x={�-;���O��<v:q=���=�N>��(>���>Y�?M9/?�dc?jZ�>��n��ξ^8¾�ߋ>T��={ �>qw=�b;>��>��7?WaE?�TK?�>Nq�=f6�>ek�>U�,���l�����T��@׏<	>�?���?F%�>�>d<�]A�4���a=�i��-�?z�/?u�?� �>�����r���q�}@���<��=�dI�?Ľ]љ=F�5������>��>]G�>++�>Ib>��O><�">���>	r>��<G��=g�)=I;�=����a�=�Ik����=�<�;������	�@3�+����;Ӕ8=�W=b W=T	�=���>�?>��>�[�=Wl���*>\z����O���=.���C9��5`�%}��z/�4>���9>��Y>n��������?�Uf>:AN>+c�?��x?Zb>�d3�-�����!c�� 1�
2�=�+�=�s\�~B��X���@��
׾O�>�܎>��>�yl>��*�O>�/�t=70��4�+L�>
����x�}���p�sȤ�������h��d4�I�D?�����=tg?
�I?��?���>s�����־�4>���'�=����
s��t��ڦ?ʪ%?ߥ�>�쾋mE��B̾���lѷ>�QI��O�g����0����ŷ����>����O�о�!3��e�� �����B�^Kr���>�O?��?lAb�W���JO����9)���p?@xg?T"�>H?A?`'��jk�jp���q�=�n?Y��?T;�?8>�3�=3r����>�	?�P�?���?��o?��D���>���>�<����=��>��=���=��?,�?�
?yV��'I��s�/:徔8_�$b'=oS�=[�>��>�hu>ua�=��1=�~�=VLZ>u؞>a=�>��w>4��>Lφ>n���qk
�nG(?�^�=h��>V�2?�#z>�XZ=M:���b<h���2�!}%��R��J���;j����A=��]�e`�>��Ŀ��?&�i>�I���?O9�i�c�5�^>?_W>/Ƚ���>eS>*7~>]��>a��>(�>�(�>o�>%�ɾu,>O���'�
�>�R�P�V۾c��>�2��9(��g
�#C����G�	��T]�*ug�[t~�z�8����<^��?�j���j�Ik����xc?��>��/?ɣp�`��Q�>z��>l#�>h��s ���򊿱e߾S�?c��?KB�>f��>]�?݁:?R#�=�S�<��g�;��@�4�1�(��~?������o��&��f/�窏?�"d?�r�>��e��c�=�P_?Y3���n��7F>��������4��wO>�ቼ�<���?�7�����]=�Ex?Z�?���>����{^���$>oL<?��0?�s?E�2?K�:?���$?��.>��?P�
?�|4?=o.?��	?�*>���=��Ļ��4=�s��Ί���̽����@S=8Au=�E���tN<Ă%=��<�R��'�����;b���[>�<ځN=@Z�=���= v�>@H?�P�>T;�>5;K?���=hK7���D�B�>|�b<q������	��l�0Ծ�?�7�?�9�?�ؾQĽ)�m�'��=</->��B>L�_=퉑>�z��3R��,�Ͻd��>
�>ߔ��Hɜ��_9�����f>����=�AS>0+
?+�>�즽\Ct=�d��ھd�b>4:ƽ��4�������U�쾟ߦ��|�>�62?��?I���t�Q�a>D#�wiP?��<?�A�?�]�?%N`>�m �YIZ���p���lX?AE�>��Ծ�/��c_����J�� �=�t�>_�������za>u��B�ݾkn� !J�y��}+Q=T���IQ=Q����Ծ�%}�K��=�s
>�O���X �i����`�� �I?2e=�[���U��
��]8>�ș>Ү><�:��hw���?�����#�=�u�>��>>8K���G��tG�������>X�A?�Z?�߁?���xw���A����u����?��>�u?��=>F�=u���(�E�a� >�yl�>`��>_W�!tE�
��L%��"�!�rm�>'?0��=G� ?��M?�? s`?h�.?�.
?0і>X���.#���%?Uw?�&:=+����߆���H���8����>��?K_��ܺ[>�?G?d�&?k�M??�c>��W�'���>z�l>�R�Ff���a�>P?��>GE\?ppr?�I>4=�(���@�=N�R>�̜>�??�|
?�?-�>;��>gǡ�e�=i��>�b?��?q�o?�R�=w�?(2>8��>NǗ=���>w�>�?6O?U�s?��J?Y�>�ɏ<b���I��#]s��sK�Wwz;CQ<�y=���&at��k����<=m�;�����c������,D��Ԑ���;���>G�K>-�J��7=}Ϥ�'����Y�=��	��������"g��T�<;��>�U?��>a�U���;P��>�"�>S�
�~�"?��?W?���=��p����@�y�j>��=?^�W>��`�Ʊ������⽨�w?ԧj?RB��� ���a?=�[?#�:�BTǾ+qt����K�N?#�?*�R����>k&{?קo?:��>{Z��i����f_��3b�t޲=��>�m��Td�I<�>[�8?P��>Q�m>P��={l۾x�𠾬�?1V�?���?&Q�?�e!>�!l���ݿ����8Ƒ�	�\?��>�¥�b]!?/h㻖�;�_��Ꮎ��߾���rR���U�������8'�4����Vؽ~º=�Z?�s?��q?�Y^?�� �}bc���]� ����U�) �����E�ǭD��C�5n��������U=�z��;���?�*?�r��s�>ə��h����Ӿ��7>��1�=e�=Ƚ��l=�=�qg���"��ի���?õ�>�5�>�8?�E]��T=�s�/��2�`��<�C>`{�>-�>G��>��<#�6�rB��� ʾ:���w�̽2�|>��`?F�H?��k?4���e5�⌁��T���4�W�����6>�a>���>�YO������#��f:�|eo�B$����������P=XR.?��~>7�>�B�?M?u�r^��
}E0��7�<���>�l?�>c�>���OR�\��>�m?83�>�|�>�+���F���x�8ҽ3��>�ר>���>�Ht>��(��Z�ߒ���f����7�U��=g?!V���)V�E��>RN?#E,���!<<K�>o�C�|����10�5�=��?��=�#0>�OǾ��� �|������'?l��>����7�����>k�1?���>Q�?ہ�>kMZ�jel�^�>"R?\�q?sD?��u>�]b�(���������PƽX>>a<>Z�;�Ӗ"��k�X��� ����+�:ܘ�=��=���O5ļ꯽�7ݼX�=�k>��ۿ��L���۾l��w��a���*�������w�����1���'���\`�˓���P��uZ�p�m�&���ʩ^�5��?��?�r��,ˉ�Ȳ��0�������x}�>0�d�9������X��Sܖ��g۾૾�	��K���c�H_�X�'?�ȑ�o�ǿ0ơ���ܾ�5 ?W� ?>�y?w��P�"�0�8�"� >�.�<D���P��L���E�ο�b���^?nZ�>|P𾮘��R�>Q�>(aY>}q>^��鉞�4c�<�?uX-?d��>�p�jɿw���"�<���?��@�$?LE�������>ȎT?�e?w�y>nq��).���	�z�%?��?C	D?	޽6H�[
��A�-?�4�>ڤ+��.2�2)>�P>G`�=��T���g>t>�>��
<vc��X�<NN=R�'>u&�=���o^�:g/�͞�>����k;Z=��?�bW�M^��D1�����!>�X?w)�>���=o�0?*A�3=Ϳw�_��d`?NO�?J��?�m"?�Ͼ�Ǟ>��ؾwG?MT7?0�>�%�:m���	>먼�S';��о�oP����=�`�>ַ>u��9�
�c���
�J��=�����ƿڙ.�W��`/4=ճ�<]YŽ-�x����g���V֑�*"M���y���)=��=4>(m>��G>�-]>�4E?�o?Ɖ�>>7�=xw��w����Ѿ�A���Q��+�1UP�����S��ھ����\����W¾�G���ܽΪY��������(s�/�I���I?�ߗ>�m��x2���>��6��8��Hv��U��2��se.�5�0��a�?��&?󷃿S�"�_����7�E[��G?�л�W9�y�����<>Ck���J
=��>Y 
>�z�����B6�(d0??U��ѽ����&>��7=��+?�6?�K<�G�>"�$?܎*��%߽i\>�k3>���>�{�>�]
>8����}ҽg!?�S?K �H����!�>'���3{���R=F>�7�,�༺�\>�y�<�����D�����6�<�W?�p�>�)�y�󄐾�?���B=j�x?S`?(Y�>O�j?��B?�k�<�9���R�R�
�jt=�0W?\�h?�a>h΃�iо�R��x5?��e?��P>�ug���辆�.����>1?Q�n?�v?���Z,}�%*������46?��v?�r^�ts�����;�V�^=�>�[�>���>��9��k�>�>?�#��G�����Y4�$Þ?��@���?(�;<��9��=�;?c\�> �O��>ƾ�z������#�q=�"�>���wev�����Q,�c�8?ؠ�?���>������.��=1
���d�?��?Kڛ���J=sB�nIk�9�u�;���=��o�R��+��:���Ҿ���l1��;S���Ă>�@�6�����>�Q�O�߿��˿EN���Ƹ��0L���?��>!ό���� Gk��Yu��G� N��;���߾>��^>"�^ժ�b1d��C����N�>A�<'`\>�UO�����F|�w�z<��>��?c�>%훾e����.�?5���X��@�����%?2<�?���?~m$?1�=��C>SL�z9D����? Ԙ?�G?�As������ �>�j?w_��UU`�ގ4�_HE��U>�"3?�B�>W�-���|=�>}��>*g>�#/�m�Ŀ�ٶ�6���Q��?܉�?�o�(��>o��?ds+?�i�8���[����*�ȥ+��<A?�2>���L�!�D0=�bҒ���
?T~0?E{�].�dlX?�LF�� ^�S	3����֪�>��F:"<��"���LFt�iq�N���W��Fx�?�D�?�\�?�N��$���?�ь>j�ľBaž�.���[>Wt ?Ȋ�>ԋ1�iD�>d����?��OM>}�?�?f?�ꋿ5򫿞� >?�i?/��>�v�?��=\O�>��=DP���r>� �">_�=��?��!??�L?�8�>��=#w:�A�/�U�E�z�Q����f�B���>�fa?WvJ?LZ>����p�D�՘ ��ɽUG3��E�J�>�e�+�=ܽC7>/?>؆>%D�u]Ͼ��?fp�3�ؿ�i��Ap'��44?p��>G�?���;�t�n��?<_?�z�>�6��+���%�� C���?gG�?��?.�׾�U̼�>��>J�>�ԽA���o�����7>M�B?Q ��D���o���>���?�@�ծ?�i��	?s��E���U~��y���6�-��=��7?W1��z>���>��=dmv�����?�s�t��>�?�?x�?���>#�l?�so��B���1==T�>��k?�n?��z�}󾦤B>�?���!����V��f?R�
@hv@��^?��A�ӿ���������P���l�=�Ǎ=q�9>�SE=��=��>�&j>+`=օ>�2�>M3>���=�J=m��=YŐ>A�v�^�,�rD��Y���%�a�qp$�2���sC��$�_�>;�¾�t�=���,쬽��I�G�ԽP@����<��;���=٩U?�R?cp?�� ?<�x�x�>����8=,�#��҄=*0�>6g2?|�L?�*?Г=������d�Q_���?���Ň�_��>gpI>)�>|I�>5'�>=}P9H�I>�*?>D}�>�� >xc'=Y��nn=��N>(M�>c��>�z�>�D>>ǋ>c3�����0h��=t�u���Ϣ?S-����J��R��4܋��3�� ʨ=0/?��>Jӑ�<�Ͽ���"�F?����S��3���>j�1?�W?��>�n���,i��A>_�
g�SM>����Zbq�l�*��XS>�O?�k>�s>��0�Rz9���R���$g�>��5?�d��?`*�l�q���I�xݾ��Q>���>�f7�N;��2���qz�2�f�f�z=p�5?�� ?G����!��Փ�𷛾�N>KoM>��=2��=�gO>��a��Iǽ��@�iL=��=>�j>�8?�si=sy#�VS�>C�v������q�>=��>^�=&L?�a?bD�<�"��0���=�B=ik�>/��=Bж=-��>�>f�?��J=�L���M�r[S�a@��z��=�,��u��UK��3��4���>��=� ��[ ���T>�Wa?�F�v�D�H��}���R\?��N?Q��=�U�=��T��9���pp�1�?�[
@�w�?8� �"g��2?Y7�?����!<|�>�_2>��;���>�6�I�c�EwӾs\�;D�?Q��?�A;>�oj��2���m2<D-?���h�>5y��Z��z��y�u�h�#=ƨ�>9H?�U����O��>�Qw
??�^�ũ����ȿ|v�j��>0�?���?$�m�zA��N@����>��?pgY?�ni>�g۾6`Z��>��@?{R?��>{9��'���?�޶?���?��L>*��?��x?;�>��B�5�(�'ձ��f���?W=;K/�*)�>�c�=l����sB� ����ފ�/i�t��F�i>x,=(^�>	�ɽ�ϸ����=�̈́����>�O�2��>q�t>�5=>��>���>��>.��>I�=@������V�� �K?��?`���3n�3��<	��=��^��&?JJ4?�Z���Ͼ�̨>�\?���?�[?�f�>���Y>���俿�{��l��<(�K>�/�>�K�>�/���-K>��Ծ�5D��d�>7̗>�`��?=ھ�+���裻�E�>�c!?��> ��= � ?<�#?P�j>�%�>jdE�>���E���>���>�/?�~?��?<Ź�\H3������ޡ�|[�!�M>��x?R??��>D����y����J� HJ��2���?�_g?]O���?�%�?Ay??�A?��f>��@�׾.+�����>�$?�	��Z����B���پZ��>_w0?��?➤>YbV>;��=F3��"�3?��?��V??���0����	���<��_�f�u=|FW<�K��t�->�y>�%=P�>�I>-��=��n��=�=�>S��>@��p��})	>�<,?vG�=ۃ���=<�r�XwD�2�>�BL>}����^?ir=���{�Z���x��ZU�� �?��?k�?���h�2#=?��?�?g �>\K���|޾̓�=Qw��{x�v�I�>��>3Tl�
徆���ڙ��G����Ž��̼T�?�0@?Щ?ŉ?�a�>�[>]Ȏ�#�"�����¾�^B�#"����w�;�eC��޵�����?>�<��q�����>�5;��y>��	?ag>%�v>C��>U*�=�f>-�>w�->�O>��:��~�=�^">��'�E"�VWG?������3:�о�\U?�bu?z�>7�߼�چ���*��{?X�?�_�?���>�J����?��V?��'?%�6	?�>��
>�R>���r�Ծ�
��A�K�~B�>�U�<	�>�ݴ=�c�����>j?��=2$����m�A
���q=�a�?��(?�w)��uQ���o�J�W�rS��/�[�g�Z<����$��`p�/܏�Xb�����.G(��M,=rA*?��?�/�)5����j�9�>���f>tz�>���>s��>�LH>ѡ	�H�1��%^�dl'�m���g��>�{?���>�~I?��;?jhP?�`L?���>�T�>�!��	�>�s�;Q�>2��>"�9?1�-?30?�h?2Z+?)c>"A��t���ؾ~�?��?L?�4?�?���CDý�s���#h�vy����G#�=Xt�<  ؽz�v�|�T=#�S>�?�'`8� ��8�a>�6?���>�
�>"ь�Et��
}�<FU�>�?��>����(Fr����m�>�ā?�-��=u	1>7�=Y�d��/��=�Qּ��=�9�^�J�1A�:;[�=�=�=+���l����:A��;��<�#�>U�&?�>�b�>�D�w��8�kB�e|.>kq&>C��=�}˾����pϙ���m��u>��?'�?�O>���=���=(ᄾ�ɾ��
�O:Ⱦ��< �?�(?��P?���?�T-?u1 ?�z3>�'"������%q�� '?K!,?L��>Y��g�ʾ��%�3��?�Z?�;a����n;)���¾O�Խ��>(Z/��.~�4���D��H�����Rx�����?ֿ�?�A�`�6�y�ھ��[��,�C?�#�>�W�>��>_�)���g��%��.;>��>FR?�>�[M?�'w?��X?#�=>><�����蹖��u��e�>C:?��?�ϋ?4�t?�1�>�>m_#��۾�5�!�+���ᅾ��?=�zS>��>��>��>���=n	��J7׽��@�	$�={v>*��>9�>GH�>�~>u��<,�G?n��>���������α��=�"���t?i��?)�+?�<=UQ�uE�ZZ��ZI�>�'�?B5�?XF&?�@L��=��ɼ�A����o�M�>�P�>*M�>��=?<C=�>Z��> ��>8���N�2�7���2�N�?J�D?���=��Ŀv3��Ն3�X7/��𼋎��8B~���>�'���)�>��=r�`>B�>/����������;�����B�����>�e>>ͭ=v��=��+>ky`=D�~���J=��=� ���}�[I�=��;���Aչ� �=���=K�����jr�� �x?b�P?x{*?bgC?�8x>���=�|;�Of�>u���Rf?��7>U�a�>���u�N�ǈ�������(̾��žrd�7X���>�i���>\9>��=�Y<c��=�/�=���=P�s;Â=�&�=cّ=N�=%�>2�>��">Ns?O~u��w��,�K�	+�?L3?�N{>�.=�ܽ��K;?�>�N���ַ��e�H�t?�r�?�C�?�) ?����Ǡ>������h=��ý�>��=��
�MF�>${I>�R�����]���!�?t@5N:?!����ӿ&O>�G>��=��W�A�H�M���t�P�]�~o%?��(������}�>��%><�ľ�-���~
=>$>��/=x$�m�T���=ut���=�1�=V�>��S>�J >Vi���~0=̇=o��=�B�=��8�⿼�ܼ?j�<�=>D�]>�y>nc�>m#?��0?�d?	f�>x�i��qξ"¾��>���=�ϱ>j �=��@>�W�>�7?��C?�ZK?f�>��=�a�>h��>#�+�hm�0�������<��?
ʆ?��>�)<_�A�����=��;Ƚo6?�w1?��?|�>��Cs���0��8�F�
�x�輳f�=����Ϸ�$�<>�X	��෽�V/>���>^ƨ>Y�H>V�>�?>�ZY>%��>M��=�J����=oA�<վE=�'�F}�=��ټݦ8��h���4=GW�=fl���u��y�<��*=�퉼��;�L��=µ�>S�>�F�>�=ꝱ�0�.>�.����M�^ӷ==����@���c�Ա}�u~.���7��/@>�3X>&6��}�����?@E\>�F>]��?�Av?$� >:��Lؾ�]���j_��WN���=F�>2@@��1<�1�_�ڦK�Ӿ���>�֐>��>�rp>�:)���<��^y=���6��v�>�m��;��\��wp�⭤���)ih���Ը��C?����\�=�}?9aJ?���?Ҟ�>@Փ�!�۾�]'>qƄ�u=���#ss�e8��S�?d�%?E��>�f�.�D���˾>���ݼ�>eH��O�=�����0�)��%���%"�>㪾�оM3��G��w���c�B��
r���>l�O?8��?��`�|F��a'O����L���En?Ug?>��?�?���K���E��C.�=�5o?���?��?^�	>�9�=*��Z��>�F
?z�?`C�?��r?��B����>��g8�$>n�����=�>6��=���=k?%�
?Z
?����@Z�2l�C��b���<���=�I�>�A�>��v>�$�=5�W=Mh�=��\>�>�
�>��c>�>��>�=��Id���&?wA�=�ߍ>Y<2?�k�>�Y=4ઽ�x�<�kH�q�>���*� -�������<X%����P=�̼^�>Zoǿ>-�?(�S>_��P?���r�/��T>�|U>��޽ ��>��E>�[}>yC�>��>�>�:�>��'>��Ծ�>��`k!�etB���R�SҾ<�{>�T����$��'�#3�x�F�	��+p�9�i��!���8=�&��<ː??:���k���)��" ��?���>UG6?���G���>@��>(�>i���NZ���p��S�ྎ�?[��?��p>�Y�>GX?Bj�>0.>5C,=�P�桉�I�;���B�1ND��t��B����3��w���l_?���?J�-?�{Խ3�=VXX?�{`��_��'.i>cW�!W�
���ȳ�>���&�;������;�=�'�?�B�?���>Qx���i��%>�:?��1?�"t?��1?_e;?B���$?.�2>�|?B�?�!5?�.?��
?nV1>`��=Q���3F%=�~���/����ν��ʽ	���1=���=�����;N�=ט�<>���@/;Rv�����<�2;=���=�#�=�ߙ>(Ns?�^>��
?ή?��4��b�rl6�om?0pa��[)�����Fa�w�q��As?,��?���?�!!��8��MH��"]=u`>�T���s=�G>Q!?=���p�=��=x�>n�e=�s�=��<�žS�ѾX��Ak���y?���>��=5^=ص̽��W����=��:�C�ݾ�m���ݾ��Ѿ�#{�|[�>�9?��?����w����p�= �D���8?�'X?��?\ʠ?���>�ϣ��w�����]���?��>CM�\����\��i \�o�i<z��>���D���~d>�
�~ݾ`�l�O�K�a���cG=s�
�'R=!�O�Ӿ��u���=Fg>bþ�!����aϨ��UH?�!c=3���T<Y�S��Q�>*�>>y�>\�9���w��@����=&��>r�I>�v�K$�6�G�� �r�y>�VM?�Pc?���?�G��G�s�bU?��J��]C�����>�?�'�>k
?<7>sj�=��������In�9I�p�>�:�>���F����M�������>��?P�.>*)?fN?q�?��]?�71?#�?��>�Z�Q����G&?Ss�?1�=��ս�T�C)9�N$F���>��)?Q�B�!~�>[z?�?-�&?gQ?�?ҧ>ٕ �@����>��>�W��W��><_>ŪJ?�ͳ>�Y?췃?��=>�5��𢾔���C��=u�>�2?/#?3�?"�>���>�롾_cz=M��>��b?�;�?L�o?���=y�?��0>�F�>n��=���>���>�"?RCO?6]s?S�J?���>_�<�]��?����r�~�M�?*�;��R<0�=�����s�U&�W�<?��;䎹�Ϯ~�ʾ�`�D�?ؐ����;^�>K	>�^����=�aþ����Ӎ>:z��������ϐ���8α>i!?��>�-.�Q<� �>E?W���?�'?S�?�=R=[~^�����d��2}�>Y�<?�@�=O�b�i���ڕ��ܸ�� ��?��t?��#�п'���b?��]?���=���þ�bc��� �O?^�
?��G��s�>��~?l�q?x��>Հe��+n�d��Kb�Gj�ٶ=B�>�c�1�d���>��7?�x�>��b>�p�=i�۾�w�Sy���?���?d�?��?�)>f�n�o�߿�`�ڨ����N?���>ib��y�?�&��7ʾ�6a���cr�(����������̫�{�'���k<Žʳ�=�?��p?�r?$�c?ۏ���Wd��K]�~Z}��
V�w�	�v��~�E�nF�>AB�ށi�.a�^��h莾�@=b�s�ه9�ܳ�?�+)?ӭ�/��>B���������ؾ��">�͓�� ���=' ��ܻ�<H�=�^�u�!���.�?~s�>��>��<?�]�ƻ;��{.�(~/�s��D?>�e�>5��>���>aT��DH�JB��Ͼɋ����߽q�H>٠s?R�T?)eq?]x�q]5�I�x�`p��k���6���n_>y��=���>xQZ�Z(8��1�\UQ�Q⃿|=�\#��? �k�F=��!?���>���>Y��?��?���r�^�WE"��]����>I�t??}�d>��)�e���l�>!�l?�l�>�ţ>刾����U{�ѓ�iK�>	Ȩ>��>��k>��2���]��+��s�4�~+>�(b?����Y��>��P?���;e��<n�>^e���#���������;>$l?�#�=�j>>4�¾��}�y����"�'?���>��{�O+����=�%?^?7Q�>�+�?2��>�ʾ�`
��0�>�b?�]?�zM?~Խ>r��fy������ݽ���<OƓ>�<�>ƿ�=�K�=R���9���@�_=ۭ@>2�;�qM��'�;�����lǼ�S��G�3>��ԿGPH�i���(�������I����B�t|��ό��B�o�)G�r/���}�E�X��Gk�������P�:{�?��?G^���9�֪��T���5�Uܪ>�O>������鬾=��������ھG1��7���D��_^�P�_�w�'?=����ǿ����+;ܾe! ?�A ?Ψy?4�П"���8�ԫ >��<s���C�뾇�����ο������^?���>
�!�����>&��>��X>.Gq>b���螾|�<��?ӄ-?���>��r���ɿ����K��<���?��@<?}��Gmݾ��=� ?(�?1�>>�#_�~�&��ƾ�d�>Y��?-��?|~�<>�Z���z��{b?���<�E���'����=��=2bO=��;��]8>�>�r��F���½;>�vj>&�<F�F�z�����[�H>��H����m?��K�<u�J�1�����&��t��?r��>��>��b?�&1�9�ۿ=1_��!U?j��?`�?z�?����ۜ>���	�'?>�%?�-�>њ�˫*���=����
\=?랾)�E�ė�=���>|!�>�����޾��o�dF*����=v=��WĿ��(�˹%��#=�<<r��G���.o�C����☾��E�ۿ�����=��=x�A>�+z>qHO>wS>��\?�f?�L�>���=��彨򃾵�ʾ�v��dy���֙�iZ��s�� �侼>۾RY�������þ��6����ߵg�j���B�A�Q���D��)?).�>#=v�k�7�:>B�u�d�x�#����UνW�ʾ.���7J�j�?�	1?�l��(���
�������G�2?��%������þ���=={�T<j��>��=c���4��kC�4�/?��?��ɾ�3���4#>1�R��4뼉7!?>?���;VÎ>��$?0i�ekν�:6>��>g�>�j�>�r>�>���c���2"?2�F?�8�0י��Z�>��������ƽ<h>�X��J��D�[>��k=�%�������a�� �8=��V?��v>��*��� �������ᓼ��c?�	?��>3RE?�t7?-4
=4�̾�v:����C�<�G?*�g?N�>1��|�F���Ū?�Mj?�J�>��[�My�ȁ,�B��%��>%�f?9-?�|�=�Ok�d����s�fG?p�v?@H^��]�����7V�i��> 4�>��>S:��>\�>?�"�$N��T����]4�c��?�@���?�1<5��Pb�=�(?�#�>��O��Bƾ�1���:���r=�
�>�d��b[v������+���8?&��?���>Y�������=ހ�3��?^V�?t�S��>t��e=x�����g>z![<�z�=�@��&�X�Ժ�j� �!z������>�		@�O=��>4��s��s��;�J���ʽ�����>)�;�!>a�d�w�T�zp��Z�~�ʾ|��)����>#T>mƽ���/�q���6�N�=��>�⧼u�T>	���Nþ]�پ=f��my�>b<�>���>�%û��þi�?�*�\����D����2�`�$?�/�?���?(�7?*S>��#�����\-ۼ8�^?I�?7T?�P0��������=
�j?�_��hU`�Ɏ4�;HE�
U>h"3?�B�>�-���|=E>���>#h>T#/�B�Ŀfٶ�+���3��?ɉ�?#o���>|��?js+?ji��7���[����*���,�e<A?G2>e�����!�T0=�-Ғ���
?Z~0?�z�@.��{]?Y']��i���0�;#��ʐ>C�����G���l;3� �\h��嚿
�r��ʫ?>�?fu�?�9'�	�!�!�'?馩>�ݕ�=�̾t�<A)�>��>��Q>��b��j>T����:��>���?<��?�|?눿PĢ�.��=�~?��>��?k �=���>���=c���X�=���>���=[$E���?h�M?���>V{�=�8���.�qF��R�	����C�6��>~�a?�=L?�d>�}��֨1�SZ!��3ӽ'm3��޼�>��13�>�ཏ�3>b�;>6�>_�B�XӾ��?+p�,�ؿ�i���o'��44?���>��?��V�t�2��<_?{�>�6��+���%���B���?GG�?��?��׾�@̼?>��>�H�>�ս����肇���7>y�B?� ��D��F�o��>u��?ֶ@�ծ?�i�	?�pK���W~�L�"�6� ��=��7?
5�W�z>v��>��=5mv�����H�s���>�@�?�y�?6��>��l?�|o���B���1=�I�>��k?�t?$Br���O�B>��?�������I��f?:�
@_u@��^? L>ӿJ����i��}�^��C�=�ȼ���=U =��<}B~>�L>Y�`>��p>��>��>�n=��=GfD>v�>��z��+�@ܠ���s���M��f5�?�vp�q$�q�<�bվ������L���ýٽx�e�Y���0�-S=��l?BiT?3Jp??�}�<]">����(׼��L��xS>���>�?��-?O�?�==�q̾M}�ֵr��1��!�����>^��=�#?�K ?�i�>��=�3�=�8>�t>��>A~	�i嗸K߽<
�[>j�>	�?�_�>�I<>��>�δ��1��m�h�w�w$̽'��?�|����J��2���6������{�=�b.?�r>����<пJ򭿈0H?[ ��5+���+��>��0?kcW?�>�����T�c'>����j�xs>> �'{l�,�)�� Q>�o?�Og>�t>�-3�3X8��#Q�����%>�#6?����ֶ6���u���H��uݾLN>9��> > ��4��疿�~�G�h���~=�/:?�|?n°�NC��I�u�����R>��Z>H�=/��=�M>��_�T�Ž=�G�3�+=�=ƭ^>�`?�>KdC=Г�>ME��U��$�>�R6>�?G>��7?AN?I�T�8n��^y�N=���]>���>�'�>��>�7-� j�=�S�>��U>��;���������
V>���1> ���ϋX����2b�<	L��k;>��=\�.f7�� _=F$v?�՞������ �n���'5Q?�2?�v�>N���.����j���e�?!
@Dg�?�����[��	?�`�?)���i�=9�	?F��>�ƾm5h�J��>y݁��ќ�(W���7����?��?n�.>j�b0x�y�J=EN*?0cJ�@o�>����Y�������u�=#=��>�1H?YF���O�\<>��s
?�?+G򾗠����ȿ<yv�)��>��?��?.�m�)A��K@��u�>#��?�fY?V]i>�g۾�xZ��p�>˱@?&R?�2�>�(�ك'��?�׶?j��?�tF>Q�?�t?���>K�x��^/�����o=��"j}=��:�b�>F��=������E����J����k�g�]>(=?T�>��0��('�=����楾�V� ��>0xr>7�I>���>� ?U2�>C��>P*=�瑽`��������K?���?%���2n�P�<z��= �^��&?}I4?	l[�g�Ͼ�ը>ٺ\?g?�[?d�>:��M>��?迿5~��Ǫ�<��K>(4�>�H�>�$���FK>��Ծ5D�Bp�>З>�����?ھ�,���U��1B�>�e!?���>sҮ=̞ ?͇#?�;j>��>�SE�B����E�v��>��>�5?+�~?\�?s����<3�����ۡ��~[� 1N>��x?�K?���>G���A~��	L���G������?�Mg?�彝�?5�?�x??ȭA?��f>����ؾJ���� �>K�'?��h�V�I��N1�Se��#?�B	?���>�.�;����V�8���6��"�/?=/m?�L?�N�{gJ��fǽY�*=Z�ϼ�Dj�q�u=�c>�R�>�Z>�M�;��
=X]`=��D>1g��h��C=�=!�>��=1H5���ܽ�:,?�2F�d؃���=Q�r��yD���>y2L>c���w�^??~=���{�$��dz��5U����?���?7m�?�[�� �h�9#=?1�?E?��>�;��w޾j��(bw��{x��m���>���>�Tl�	徙�������PE��n�Ž�m���?�I? �.?��!?��>��)>>���9�P��z�N�νxN������=�=<:��� ���ȩ��[���UE���@s�	P�>�%�=bD>ݠ?Θ�>bq�>/�>�Q�^�u>�s�>��g>!�W>�.�=��.>g<q> %�<�� �ЎO?��Ͼ( ����.n���w8?Q!W?�?����Ig��'���s?p!�?Ji�?�Ŵ>�p���7��L ?��0?́g�0��>��>Cr=��<)�ľ��[���D�Gӗ�4�o>�����:�[�H��D��d�>�&?O�== �g=D\���v=�h�?�%)?֣)��Q�͔o���W���R���L�f�(���?:$�=hp��������'���(�u�%=��)??�?�����҅���Dk���>��g>���>�ϖ>�#�>�G>�c	��[1�l~]��'��E��1�>h�z?k&�>�J?W�:?��Q?l�P?�!�>��>Sx�����>|4����>�{�>�44?_j*?Vp.?)�?�'?��R>.���7|���$Ծ��?I�?��?Et?���>}�����c 4�D�>:�a�ud���Z=��<k�����C�3��=.\=>R�$?Gn�0�O��2�W�A>�S:?R�>G��>�s�p֪�q��hU�>�(?���>9`��]C�����L�>���?���Vm���JM>��=�����=܉<>ǰ>B�g�C��;=mJ8;��i>_y>�U�=�tj�!u���<#	F;O��>�|?�:B>���>�0F�2 #��� 2L<��h>�\=�W��Y��b����	��	-j��i>U�?���?��þ�[�=�>6�|��ٗ��|׾Z���4��SW�>���>�H+?�$�?[7(?E?���=(���f�r�����AF?�!,?p�>����ʾ�꨿8w3�ǝ?@c?17a����<)���¾.	Խ7>�?/��3~�J���D�j�i�=���K��i��?G��?tA���6����K���m\���C?�
�>�8�>���>��)�R�g���S;>��>sR?8	�>��O?G+{?�[?v�i>e�2�}᫿(���,	�ɯ>DOB?H�?�,�?f+t?�;�>�>zn)���޾ם���&�F�齇"����T=��X>���>��>	�>���=�~ӽ�ĺ�D�8��B�=��Z>�8�>�t�>e��>I�~>�f�<r�F?���>p���p�ߣ�Ј�Y�A���p?�o�?�(?{o%<,����G�.�����>l�?��?�n)?�d����=�ϼ���.�j�S�>6�>n3�>}�=�D= w>�%�>4B�>���fW�i}7�Փ��b9?��I? �=�Ͽ�Z��))��0��*�=%yj�b�־��s>v�]=�?����*I�>
m�=������sľ)mƾAy)���=��i7?��>����QD���6=z��-�M��_,��-�=�����c��:/q�����l�a��3��?��ٱ�=HǶ=�*����|?�NV?5�-?]�a?��>29�=e��p >��4�,?&K�>Vb�2�����=����������� #���DQ������q>ޔ����K>n�~>֍>*�=w=�0=�5=�J�=��H=Tց=�����'6=��u>�x�>M(:>�Ql?Al�K���z$J������	?&�>;�`>����e>B?���>ڈ��7%���5�)I�?�b�?�Ƽ?�>6�J�Q��>/4پB��:��R�\�s����=���>H��((�>B��>ɂ+��"���������?���?��M?���dп�>�yN>�`�=H|P���/�72U��E��D���b�?Z+�$�ƾ.�i>ؗ�=�Ҿ����D�<�c>��F=���z�N��p�=\ew��w�=i��<�o>�YB>"��=�����r=��=��=5x'>LY�������:<��={׹=��K>.�:>���>�?� (?!@f?�>�F��nǾ6վ�O>{�O=�²>��x=$��=��>L@&?�@?U�S?���>p�5<�>L��>�6'�E0x�`��~�����g=��?(��?p�>d =�{����Z'��y���!?pt+?�z�>���>Ԕ�w�ݿ	�$��z.�w�it%����<�kS����W�n���약� >Yk�>�e�>CK�>~d>z�#>V?>�x�>b>�c�<P�q<���;
�=T� �Ń=g2ڼv=�BT�o:��c<8�輂���@�<��<Q��<��;�Y�=���>��=��>�U�=�N����=j���}G���m=��.1�'�e����o/?�q`V���q>Ӓ>��}Ή����>#�S>�l>t��?�؀?���>�bU���	�Ҝ���������b=��>����2�(���T�	@� ���5Ѯ>Wu�>��>ך>��(��)>�8�=��龷�(���>�a����Z�/��uh��8��i�����s�[�ֽ�%?�{��w�&><�{?�J8?�}|?�݌>�����,��W7{>�$��CO=��"�]�H���	��(?d�'?�ڒ>1��/;�~ʾ*п�K�>�6D�O�@Δ�k0�����޷����>!��~оsu2����㏿�A��?p���>`O?8�?J8]�����%CN����-����?��e?D�>fc?�?}������_���j�=��o?7\�?���?��>�~�=Ӗ����>L?-��?]�?b,o?�aW�|��>�ؑ��+>�ǁ����=���=�w=���=�M?ө?��?�֑����(��z�}b�yZ�<lJ�=��>r��>�n>^��=�zF=�?�=[Z>
�>���>u�r>�s�>��>����7���'?ܽ�=�\�>*�1?6�>wzV=f~�����<3�.�5\<��)�ך��֟��ݯ<��-�W2=�lټ݂�>�ƿX�?ӺR>M�M=?�b�sV�O�Q>��V>Upս�>5'A>��{>T�>��>�>V�>��.>��վ(�>Z;��Z"��AB���P��ZҾ��|>E���"��O�m��7[E��\���.��i�3ၿȹ<�Ӏ�<d�?p���l��+�������?� �>��5?����$�����	>+��>M��>�����!��x��V��U�?�P�?T��>).�>��Z?�&?b�#��k�1�5�*�d�P��cC�Ta��>t�a�q����2�9�Xop?�V�?$�)?�e���9>�b?�z��z��*i%>��<�Z��%����> ���
�����JA��������>�p?���?�&�>���uhm�'>P�:?ʙ1?uLt?o�1?K|;?~���$?ee3>K?�j?G5?��.?��
?�1>��=����p�(=�8���抾+cѽA1ʽ��[T4=��{=Fᘷ�<Ѹ=J��<�e��ؼ�U;����<h�:=,��=�*�=i��>��]?���>��>�4?���#}6��EվN�?傈����moy��Qþ�#��ZQ<�"R?�c�?&�]? ��=�<�
�.��� >�'�>��%>��>���>���F���%���/>d3>�=�=�
���т��e�?���vr{=�{>܋?�l�>���=�GT>�_;�Mн�|>ݖ2����ݣ�t�Ri�����.x�>hmL??V<?�Hռ�<��&=o\9���2?��-?�&a?n��?�)Q>ϥQ��^��[{�͏⾘$?��>���J���䪿�>>��N=�ϡ>��񾥓���za>u��B�ݾkn� !J�y��}+Q=T���IQ=Q����Ծ�%}�K��=�s
>�O���X �i����`�� �I?2e=�[���U��
��]8>�ș>Ү><�:��hw���?�����#�=�u�>��>>8K���G��tG�������>X�A?�Z?�߁?���xw���A����u����?��>�u?��=>F�=u���(�E�a� >�yl�>`��>_W�!tE�
��L%��"�!�rm�>'?0��=G� ?��M?�? s`?h�.?�.
?0і>X���.#���%?Uw?�&:=+����߆���H���8����>��?K_��ܺ[>�?G?d�&?k�M??�c>��W�'���>z�l>�R�Ff���a�>P?��>GE\?ppr?�I>4=�(���@�=N�R>�̜>�??�|
?�?-�>;��>gǡ�e�=i��>�b?��?q�o?�R�=w�?(2>8��>NǗ=���>w�>�?6O?U�s?��J?Y�>�ɏ<b���I��#]s��sK�Wwz;CQ<�y=���&at��k����<=m�;�����c������,D��Ԑ���;���>G�K>-�J��7=}Ϥ�'����Y�=��	��������"g��T�<;��>�U?��>a�U���;P��>�"�>S�
�~�"?��?W?���=��p����@�y�j>��=?^�W>��`�Ʊ������⽨�w?ԧj?RB��� ���a?=�[?#�:�BTǾ+qt����K�N?#�?*�R����>k&{?קo?:��>{Z��i����f_��3b�t޲=��>�m��Td�I<�>[�8?P��>Q�m>P��={l۾x�𠾬�?1V�?���?&Q�?�e!>�!l���ݿ����8Ƒ�	�\?��>�¥�b]!?/h㻖�;�_��Ꮎ��߾���rR���U�������8'�4����Vؽ~º=�Z?�s?��q?�Y^?�� �}bc���]� ����U�) �����E�ǭD��C�5n��������U=�z��;���?�*?�r��s�>ə��h����Ӿ��7>��1�=e�=Ƚ��l=�=�qg���"��ի���?õ�>�5�>�8?�E]��T=�s�/��2�`��<�C>`{�>-�>G��>��<#�6�rB��� ʾ:���w�̽2�|>��`?F�H?��k?4���e5�⌁��T���4�W�����6>�a>���>�YO������#��f:�|eo�B$����������P=XR.?��~>7�>�B�?M?u�r^��
}E0��7�<���>�l?�>c�>���OR�\��>�m?83�>�|�>�+���F���x�8ҽ3��>�ר>���>�Ht>��(��Z�ߒ���f����7�U��=g?!V���)V�E��>RN?#E,���!<<K�>o�C�|����10�5�=��?��=�#0>�OǾ��� �|������'?l��>����7�����>k�1?���>Q�?ہ�>kMZ�jel�^�>"R?\�q?sD?��u>�]b�(���������PƽX>>a<>Z�;�Ӗ"��k�X��� ����+�:ܘ�=��=���O5ļ꯽�7ݼX�=�k>��ۿ��L���۾l��w��a���*�������w�����1���'���\`�˓���P��uZ�p�m�&���ʩ^�5��?��?�r��,ˉ�Ȳ��0�������x}�>0�d�9������X��Sܖ��g۾૾�	��K���c�H_�X�'?�ȑ�o�ǿ0ơ���ܾ�5 ?W� ?>�y?w��P�"�0�8�"� >�.�<D���P��L���E�ο�b���^?nZ�>|P𾮘��R�>Q�>(aY>}q>^��鉞�4c�<�?uX-?d��>�p�jɿw���"�<���?��@�$?LE�������>ȎT?�e?w�y>nq��).���	�z�%?��?C	D?	޽6H�[
��A�-?�4�>ڤ+��.2�2)>�P>G`�=��T���g>t>�>��
<vc��X�<NN=R�'>u&�=���o^�:g/�͞�>����k;Z=��?�bW�M^��D1�����!>�X?w)�>���=o�0?*A�3=Ϳw�_��d`?NO�?J��?�m"?�Ͼ�Ǟ>��ؾwG?MT7?0�>�%�:m���	>먼�S';��о�oP����=�`�>ַ>u��9�
�c���
�J��=�����ƿڙ.�W��`/4=ճ�<]YŽ-�x����g���V֑�*"M���y���)=��=4>(m>��G>�-]>�4E?�o?Ɖ�>>7�=xw��w����Ѿ�A���Q��+�1UP�����S��ھ����\����W¾�G���ܽΪY��������(s�/�I���I?�ߗ>�m��x2���>��6��8��Hv��U��2��se.�5�0��a�?��&?󷃿S�"�_����7�E[��G?�л�W9�y�����<>Ck���J
=��>Y 
>�z�����B6�(d0??U��ѽ����&>��7=��+?�6?�K<�G�>"�$?܎*��%߽i\>�k3>���>�{�>�]
>8����}ҽg!?�S?K �H����!�>'���3{���R=F>�7�,�༺�\>�y�<�����D�����6�<�W?�p�>�)�y�󄐾�?���B=j�x?S`?(Y�>O�j?��B?�k�<�9���R�R�
�jt=�0W?\�h?�a>h΃�iо�R��x5?��e?��P>�ug���辆�.����>1?Q�n?�v?���Z,}�%*������46?��v?�r^�ts�����;�V�^=�>�[�>���>��9��k�>�>?�#��G�����Y4�$Þ?��@���?(�;<��9��=�;?c\�> �O��>ƾ�z������#�q=�"�>���wev�����Q,�c�8?ؠ�?���>������.��=1
���d�?��?Kڛ���J=sB�nIk�9�u�;���=��o�R��+��:���Ҿ���l1��;S���Ă>�@�6�����>�Q�O�߿��˿EN���Ƹ��0L���?��>!ό���� Gk��Yu��G� N��;���߾>��^>"�^ժ�b1d��C����N�>A�<'`\>�UO�����F|�w�z<��>��?c�>%훾e����.�?5���X��@�����%?2<�?���?~m$?1�=��C>SL�z9D����? Ԙ?�G?�As������ �>�j?w_��UU`�ގ4�_HE��U>�"3?�B�>W�-���|=�>}��>*g>�#/�m�Ŀ�ٶ�6���Q��?܉�?�o�(��>o��?ds+?�i�8���[����*�ȥ+��<A?�2>���L�!�D0=�bҒ���
?T~0?E{�].�dlX?�LF�� ^�S	3����֪�>��F:"<��"���LFt�iq�N���W��Fx�?�D�?�\�?�N��$���?�ь>j�ľBaž�.���[>Wt ?Ȋ�>ԋ1�iD�>d����?��OM>}�?�?f?�ꋿ5򫿞� >?�i?/��>�v�?��=\O�>��=DP���r>� �">_�=��?��!??�L?�8�>��=#w:�A�/�U�E�z�Q����f�B���>�fa?WvJ?LZ>����p�D�՘ ��ɽUG3��E�J�>�e�+�=ܽC7>/?>؆>%D�u]Ͼ��?fp�3�ؿ�i��Ap'��44?p��>G�?���;�t�n��?<_?�z�>�6��+���%�� C���?gG�?��?.�׾�U̼�>��>J�>�ԽA���o�����7>M�B?Q ��D���o���>���?�@�ծ?�i��	?s��E���U~��y���6�-��=��7?W1��z>���>��=dmv�����?�s�t��>�?�?x�?���>#�l?�so��B���1==T�>��k?�n?��z�}󾦤B>�?���!����V��f?R�
@hv@��^?��A�ӿ���������P���l�=�Ǎ=q�9>�SE=��=��>�&j>+`=օ>�2�>M3>���=�J=m��=YŐ>A�v�^�,�rD��Y���%�a�qp$�2���sC��$�_�>;�¾�t�=���,쬽��I�G�ԽP@����<��;���=٩U?�R?cp?�� ?<�x�x�>����8=,�#��҄=*0�>6g2?|�L?�*?Г=������d�Q_���?���Ň�_��>gpI>)�>|I�>5'�>=}P9H�I>�*?>D}�>�� >xc'=Y��nn=��N>(M�>c��>�z�>�D>>ǋ>c3�����0h��=t�u���Ϣ?S-����J��R��4܋��3�� ʨ=0/?��>Jӑ�<�Ͽ���"�F?����S��3���>j�1?�W?��>�n���,i��A>_�
g�SM>����Zbq�l�*��XS>�O?�k>�s>��0�Rz9���R���$g�>��5?�d��?`*�l�q���I�xݾ��Q>���>�f7�N;��2���qz�2�f�f�z=p�5?�� ?G����!��Փ�𷛾�N>KoM>��=2��=�gO>��a��Iǽ��@�iL=��=>�j>�8?�si=sy#�VS�>C�v������q�>=��>^�=&L?�a?bD�<�"��0���=�B=ik�>/��=Bж=-��>�>f�?��J=�L���M�r[S�a@��z��=�,��u��UK��3��4���>��=� ��[ ���T>�Wa?�F�v�D�H��}���R\?��N?Q��=�U�=��T��9���pp�1�?�[
@�w�?8� �"g��2?Y7�?����!<|�>�_2>��;���>�6�I�c�EwӾs\�;D�?Q��?�A;>�oj��2���m2<D-?���h�>5y��Z��z��y�u�h�#=ƨ�>9H?�U����O��>�Qw
??�^�ũ����ȿ|v�j��>0�?���?$�m�zA��N@����>��?pgY?�ni>�g۾6`Z��>��@?{R?��>{9��'���?�޶?���?��L>*��?��x?;�>��B�5�(�'ձ��f���?W=;K/�*)�>�c�=l����sB� ����ފ�/i�t��F�i>x,=(^�>	�ɽ�ϸ����=�̈́����>�O�2��>q�t>�5=>��>���>��>.��>I�=@������V�� �K?��?`���3n�3��<	��=��^��&?JJ4?�Z���Ͼ�̨>�\?���?�[?�f�>���Y>���俿�{��l��<(�K>�/�>�K�>�/���-K>��Ծ�5D��d�>7̗>�`��?=ھ�+���裻�E�>�c!?��> ��= � ?<�#?P�j>�%�>jdE�>���E���>���>�/?�~?��?<Ź�\H3������ޡ�|[�!�M>��x?R??��>D����y����J� HJ��2���?�_g?]O���?�%�?Ay??�A?��f>��@�׾.+�����>�$?�	��Z����B���پZ��>_w0?��?➤>YbV>;��=F3��"�3?��?��V??���0����	���<��_�f�u=|FW<�K��t�->�y>�%=P�>�I>-��=��n��=�=�>S��>@��p��})	>�<,?vG�=ۃ���=<�r�XwD�2�>�BL>}����^?ir=���{�Z���x��ZU�� �?��?k�?���h�2#=?��?�?g �>\K���|޾̓�=Qw��{x�v�I�>��>3Tl�
徆���ڙ��G����Ž��̼T�?�0@?Щ?ŉ?�a�>�[>]Ȏ�#�"�����¾�^B�#"����w�;�eC��޵�����?>�<��q�����>�5;��y>��	?ag>%�v>C��>U*�=�f>-�>w�->�O>��:��~�=�^">��'�E"�VWG?������3:�о�\U?�bu?z�>7�߼�چ���*��{?X�?�_�?���>�J����?��V?��'?%�6	?�>��
>�R>���r�Ծ�
��A�K�~B�>�U�<	�>�ݴ=�c�����>j?��=2$����m�A
���q=�a�?��(?�w)��uQ���o�J�W�rS��/�[�g�Z<����$��`p�/܏�Xb�����.G(��M,=rA*?��?�/�)5����j�9�>���f>tz�>���>s��>�LH>ѡ	�H�1��%^�dl'�m���g��>�{?���>�~I?��;?jhP?�`L?���>�T�>�!��	�>�s�;Q�>2��>"�9?1�-?30?�h?2Z+?)c>"A��t���ؾ~�?��?L?�4?�?���CDý�s���#h�vy����G#�=Xt�<  ؽz�v�|�T=#�S>�?�'`8� ��8�a>�6?���>�
�>"ь�Et��
}�<FU�>�?��>����(Fr����m�>�ā?�-��=u	1>7�=Y�d��/��=�Qּ��=�9�^�J�1A�:;[�=�=�=+���l����:A��;��<�#�>U�&?�>�b�>�D�w��8�kB�e|.>kq&>C��=�}˾����pϙ���m��u>��?'�?�O>���=���=(ᄾ�ɾ��
�O:Ⱦ��< �?�(?��P?���?�T-?u1 ?�z3>�'"������%q�� '?K!,?L��>Y��g�ʾ��%�3��?�Z?�;a����n;)���¾O�Խ��>(Z/��.~�4���D��H�����Rx�����?ֿ�?�A�`�6�y�ھ��[��,�C?�#�>�W�>��>_�)���g��%��.;>��>FR?�>�[M?�'w?��X?#�=>><�����蹖��u��e�>C:?��?�ϋ?4�t?�1�>�>m_#��۾�5�!�+���ᅾ��?=�zS>��>��>��>���=n	��J7׽��@�	$�={v>*��>9�>GH�>�~>u��<,�G?n��>���������α��=�"���t?i��?)�+?�<=UQ�uE�ZZ��ZI�>�'�?B5�?XF&?�@L��=��ɼ�A����o�M�>�P�>*M�>��=?<C=�>Z��> ��>8���N�2�7���2�N�?J�D?���=��Ŀv3��Ն3�X7/��𼋎��8B~���>�'���)�>��=r�`>B�>/����������;�����B�����>�e>>ͭ=v��=��+>ky`=D�~���J=��=� ���}�[I�=��;���Aչ� �=���=K�����jr�� �x?b�P?x{*?bgC?�8x>���=�|;�Of�>u���Rf?��7>U�a�>���u�N�ǈ�������(̾��žrd�7X���>�i���>\9>��=�Y<c��=�/�=���=P�s;Â=�&�=cّ=N�=%�>2�>��">Ns?O~u��w��,�K�	+�?L3?�N{>�.=�ܽ��K;?�>�N���ַ��e�H�t?�r�?�C�?�) ?����Ǡ>������h=��ý�>��=��
�MF�>${I>�R�����]���!�?t@5N:?!����ӿ&O>�G>��=��W�A�H�M���t�P�]�~o%?��(������}�>��%><�ľ�-���~
=>$>��/=x$�m�T���=ut���=�1�=V�>��S>�J >Vi���~0=̇=o��=�B�=��8�⿼�ܼ?j�<�=>D�]>�y>nc�>m#?��0?�d?	f�>x�i��qξ"¾��>���=�ϱ>j �=��@>�W�>�7?��C?�ZK?f�>��=�a�>h��>#�+�hm�0�������<��?
ʆ?��>�)<_�A�����=��;Ƚo6?�w1?��?|�>��Cs���0��8�F�
�x�輳f�=����Ϸ�$�<>�X	��෽�V/>���>^ƨ>Y�H>V�>�?>�ZY>%��>M��=�J����=oA�<վE=�'�F}�=��ټݦ8��h���4=GW�=fl���u��y�<��*=�퉼��;�L��=µ�>S�>�F�>�=ꝱ�0�.>�.����M�^ӷ==����@���c�Ա}�u~.���7��/@>�3X>&6��}�����?@E\>�F>]��?�Av?$� >:��Lؾ�]���j_��WN���=F�>2@@��1<�1�_�ڦK�Ӿ���>�֐>��>�rp>�:)���<��^y=���6��v�>�m��;��\��wp�⭤���)ih���Ը��C?����\�=�}?9aJ?���?Ҟ�>@Փ�!�۾�]'>qƄ�u=���#ss�e8��S�?d�%?E��>�f�.�D���˾>���ݼ�>eH��O�=�����0�)��%���%"�>㪾�оM3��G��w���c�B��
r���>l�O?8��?��`�|F��a'O����L���En?Ug?>��?�?���K���E��C.�=�5o?���?��?^�	>�9�=*��Z��>�F
?z�?`C�?��r?��B����>��g8�$>n�����=�>6��=���=k?%�
?Z
?����@Z�2l�C��b���<���=�I�>�A�>��v>�$�=5�W=Mh�=��\>�>�
�>��c>�>��>�=��Id���&?wA�=�ߍ>Y<2?�k�>�Y=4ઽ�x�<�kH�q�>���*� -�������<X%����P=�̼^�>Zoǿ>-�?(�S>_��P?���r�/��T>�|U>��޽ ��>��E>�[}>yC�>��>�>�:�>��'>��Ծ�>��`k!�etB���R�SҾ<�{>�T����$��'�#3�x�F�	��+p�9�i��!���8=�&��<ː??:���k���)��" ��?���>UG6?���G���>@��>(�>i���NZ���p��S�ྎ�?[��?��p>�Y�>GX?Bj�>0.>5C,=�P�桉�I�;���B�1ND��t��B����3��w���l_?���?J�-?�{Խ3�=VXX?�{`��_��'.i>cW�!W�
���ȳ�>���&�;������;�=�'�?�B�?���>Qx���i��%>�:?��1?�"t?��1?_e;?B���$?.�2>�|?B�?�!5?�.?��
?nV1>`��=Q���3F%=�~���/����ν��ʽ	���1=���=�����;N�=ט�<>���@/;Rv�����<�2;=���=�#�=�ߙ>(Ns?�^>��
?ή?��4��b�rl6�om?0pa��[)�����Fa�w�q��As?,��?���?�!!��8��MH��"]=u`>�T���s=�G>Q!?=���p�=��=x�>n�e=�s�=��<�žS�ѾX��Ak���y?���>��=5^=ص̽��W����=��:�C�ݾ�m���ݾ��Ѿ�#{�|[�>�9?��?����w����p�= �D���8?�'X?��?\ʠ?���>�ϣ��w�����]���?��>CM�\����\��i \�o�i<z��>������M<b>�����޾�n�0-J��b羴`P=���ŠU=��־5�~�?��=�	>n���,� �6���ɪ�,=J?�hl=v���JU�w����>U��>��>�^<�Z%v��@�����9�=���>Q�9>-���D�wG���a!�>*�C?�3U?�ވ?�g�M�o��/N�٭��Q��v�V��"?y�>hy�>v�>���=v�����ޔ`�'s@����>_��>����*H�l�����T3�cǋ>G?b�=v
?��W?t�?��]?05?��	?"�>,&���¾��%?W��?�sp��9�<�y�H���K�U�Ž�>Su&?I���?�>N2D?��C?�V�>=@?�6?\�>�T���b�'�b>Q�>��-��쫿0�>�1?<�>>E8?��q?/��>�S�����P>N�>��>j�?�{?�@�>1�>���> k��N�=s�>�d?��?�n?�S�=�; ?W�7>���>e�=��>.��>4?(EO?=�q?�L?�e�>�?�< /���s��	�����)����;ĠX<C��=G���g�z��|
�<��;l�μ��xk�B�L�@`&�Ds0<�_�>��s>
����0><�ľ(P��{�@>҅��wP���ي��:�:ݷ=�>{�?���>,Y#�d��=���>xI�>5���6(?��?�?�!;ˡb���ھM�K�$�>	B?\��=��l�������u���g=��m?��^?'�W�\&��;e^?��]?uF�*��������f�9��UH?&N?N茶X�>`��?J.b?%Ϻ>^P�<jK������k��~���=��>�E#���o�Gi�>��9?��?��i>��S>ؔ��L��)����+?�f�?�u�?�c�?I��>s|��ܿ����"��Y^?�9�>Ʀ�I�"?���'�ξ�ҋ�񾎾��Të��������Ħ���$�[����ֽS0�=j ?s?�?q?��_?ý ��%d���]�C���yV�j������E�ϝD�tC���n���������k��msK=E�]��3�3�?r#?郛�Ȟ�>����˾����;�r>�.۾i�����=M߽x����*=�z���;�]����?�C�>�c�>=6O?�Z�V2F���+��O%�
Z��L>h�>l�z>���>�+0�U�4�au�U|㾴����:�9v>9vc?1�K?�n?�l��(1����7�!���/�4c���B>�c>P��>�W�K��5<&��Y>���r�[���w����	�|�~=R�2?�*�>���>�N�?�?(z	��o��}ox�m�1�Զ�<�3�>3i?�A�>]�>нJ� ���>�l?���>5�>�|��mL!���{�.˽��>��>��>�o>�C-�hC\�|k��H����69��m�=X�h?����[�`�8�>��Q?���:U�V<l�>vFt�V�!�5B�:�'�I�>�Y?9��=��;>��ž6	���{�������&?*M?6iz���Z�M��>���>�^>�4�>{j?��>9�ľ�P;qg(?�kO?cNa?fU?�Y?�>l�ѾQ�����c��=��l>F�=���<N&I>r�ǾH���1�]ݎ>�R
>Ͽ����l=�
R=���=%�?>W��=��G>Ĭ��[N�Ȇ�I��4����4	���Ϻb��=�d�����Wq�����^s]�hFW=O�F�D����8����$�?)R�?�6O��N������F���d��"3#?;2�����u��= r���;��q���v4"��S��P�<�t���'?A���I�ǿY����ܾ|�?�l ?b�y?{"�v�"��v8� >}��<t������������οr��w�^?���>��������>a�>�W>�p>��'���l�<Ȱ?�^-?���>��s�]�ɿh������<2��?@PtA?��(�׹���V=3��>��	?&?>�0��9�ED���s�>�;�?���??�L==�W����%]e?*�;��F��1ܻ���=���="7=w��C�J>���>���,A��ܽ��3>*��>Cd�@�h�]�+'�<e�]>�_ս���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�~���ſ�&����������E=�����.���U_�r��;�X��e"��-�=�c�=N<>���>g;o>�g�>��_?�Fe?�ӥ>iB	>��ɽ*����8��^�q=Jڗ�_���.��̑8�@O��P վg%����X�pl�N�̾�=�/�=~?R����k� ���b�,YF��.?��$>��ʾ/�M��,<Vjʾ�r�����xƥ��̾�l1���m�Z֟?�B?�ꅿ[�V������
��긽��W?�������=3����=멜>_�=���3�r�S�v0?i�?�O���@����+>�� ��G=�+?��?%o<F�>W�$?�)��y���\>��4>�=�>X��>��>���qٽ�i?pT?x�ʜ���>m���
 z�Q�b=�r>N�4�����\>�<o����F����4�<4(W?��>]�)�h��c���C��==��x?�?�+�>]yk?��B?��<L_��P�S�: �GXw=��W?u'i?M�>�t���о���<�5?T�e?f�N>*[h������.��U��"?��n?�\?�"��g{}�,��N���o6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������#��=dǕ��^�?W�?�U��5Fe<��Y�k�(���<�<���=����"�w��.�7���ƾ��
��o��욿�u��>LO@��;t�>��8��/�WMϿM��Zо	"q���?��>=iȽ����z�j�"Ku�]�G��H�)o���/�>�~>�.��5瑾��{�rL;��G�����>������>87S���������9<��>3��>�>��������UǙ?���-ο����R��LzX?Fa�?3}�?�.?C�7<R�v���{����$G?�Xs?tZ?�%�x�\�@�9��k?�f����\��Q3�f~G�IG>��3?a7�>v�-�6�=7P>�>�L>N�/���Ŀ����% �ʎ�?p�?J�龃��>z=�?a�,?%>��y��s���-,��O�;vA?��,>���ˌ#��/@�5q���?A�/?�����з_?x�a�!�p�m�-�d�ƽ�ۡ>��0��h\��v������Ve�n��`<y�y��?�]�?8�?׵�S #��4%?�>���6Ǿj��<р�>�)�>�+N>S#_���u>#���:��h	>��?\}�?�i?򕏿k���*]>��}?c$�>��?�n�=�a�>Gd�=E�y-��k#>�"�=s�>��?��M?L�>FW�=z�8�~/�7[F��GR�d$�=�C� �>��a?ނL?tKb>���2��!��uͽc1��Q��W@��,�r�߽D(5>��=>�>P�D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?PQo���i�B>��?"������L��f?�
@u@a�^?*�ƿ�𒿾Y��V{������/��>��>P7�ɹi>�
+��	�=��Y=���¡�>O��>�3_>V�>^m>82>�Xv�M�"�FS��~&|��9g��Ҧ���쾬`ɾ�ʄ��;aj��;�����Ez$9�I��J�%��7=&�þ�� 9���=@�U?�R?�	p?� ?=Ix�ݍ>9���&�=�j#�v�=*�>�j2?��L?T�*?M!�==����d��`��;7���և�Q��>/I>��>oJ�>*�>�9��I>TN?>Rt�><� >:�'=*캃v=#�N>�(�>��>`��>D<>��>/ϴ��1��]�h�fw�/̽A�?����@�J��1���9��2���k�=�a.?w{>����>пL����2H?|��� )���+���>��0?�cW?��>V��t�T�89>���T�j��_>�- �ށl�ߎ)�%Q>�l?^�f>�%u>c�3�~b8�:�P��v���X|>�46?�嶾�<9��u���H��Tݾ�GM>i��>�8C��h�@���z��gi��{=4x:?=�?r ���簾��u�<���?R>]W\><=;�=dYM>AOc��ƽZH�.=i��=@�^>~W?��+>�=fȣ>�H��C.P����>ՊB>��+>f@?C&%?6��ͱ��,}���-�"w>uI�>1�>�J>�RJ�ɯ=�k�>��a>$�����i��C�?��VW>`�}� |_��Ru���x=;<�����=��='� �?�<��&=�~?���(䈿��!e���lD?U+?| �=F<��"�D ���H��F�?r�@m�?��	�ߢV�?�?�@�?��\��=}�>׫>�ξ"�L��?��Ž9Ǣ�ǔ	�3)#�hS�?��?��/�[ʋ�Al�p6>�^%?��Ӿth�>�x�sZ�������u�@�#=���>�8H?�V����O�w>��v
? ?�^�㩤���ȿ5|v����>P�?���?V�m�bA���@�)��>#��?ogY?�ni>�g۾�_Z�q��>��@?�R?P�>�9�	�'�J�?�޶?﯅?:3I>���?�s?Ϫ�>��w�,\/�4<�������v~=�_;��>ƃ>����sF��Փ��`����j�+����a>�$=�,�> 彆0��؉�=�����R����f�F̷>�p>��I>z��>I� ?,\�>ڙ>�]=̓������Ė��NF?�Ó?����wg��6>��=U���]�?�):?�UL<R���U �>~~x?k?�"^?Vb�>�D������簽��z���=c�>��y>�-�>L�꽔ws>=N���l0��9�>>Ԟ������@��Ū=�B>��>t�?!A�=��?�k?.�s>��;?Wf�>T��(���&�>�>�(?� �?:�	?���A�X��E��L���h���>@eS?>�?���>#e��tx���=��j<����I?��?-�Ⱦ=6C?��?� ?��?�x�>�a=�4�b@��1
�=l�!?�P���A�&��d�5b?d�?M,�>�M����ٽ0ڼIF������?�\?��&?���ma�<-ľ,R�<ǟ�R0��Z�;L(B��X>�>�܇�A��=�g>PA�=�o��F5�-т<ª�=#�>k��=@�5�%���0=,?��G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>'�l���K���ڙ���F��^�Ž�m���h�>�W?;�>���>k>�Kw>�D���6��A���F���x�dx-�nH��G��G<������[�7�A�������6��\�>��B���>h. ?ʈ�>M��>�V&>���<��>=�=�Y>g�>N9\>���>�i�<�YN�5:k��KR?�����'���辠���^3B?�qd?`1�>�i�2��������?���?Rs�?4=v>�~h��,+��n?�>�>7��Kq
?�T:=�;�;�<V��i���2����9��>(E׽� :��M�Pnf�hj
?�/?]����̾e;׽C[��j�=2I�?�zF?%�
�+-J���Z�)�%��w����=�b��-/�ø�j�z���}�|�����/���M�=9�#?<�p?�9�e�uK�`�n���c�mH>�%�>���>�~#?X!�> Q�*o8��a��m�ŬO�z�?��p?�>]OV?�Q/?p�?��[?��>n�~>�����>�}=���>v��>��9?L�@?%NG?;:?"�<?�@>�p����H
���?0?u?���>S]?lL*�3먾ܢ�t0L=�i�����<$��<w�߽�R_�̈́Y<��v>�X?)���8������k>R�7?��>���>����,�����<�>��
?�F�>1 �~r� c��V�>t��?J��Ƀ=��)>���=劅��Һ�Z�=$�����=\5���y;��a<쁿=���=�Kt�����A�:1��;�j�<�u�>1�?P�>�=�>y ���� �e�����=9�V>wT>�>L�پ�k��,���h��Gx>Y�?V��?Q�h=��=���=m��eK�� ���1����< t?�d#?�T?�̒?#>?��"?��>e0���?!��}���V�?g�:?�rU>��ᾫ�Ҿ�﮿�u�4f/?�0?K�e��	�(8�]�Ѿ ��=�:>�R�o�������:K�~iP>��˾�ܽ�^�?_��?��w�M��������x��V?X?aEJ>��>��>G���������-��UI�N��>P�?}!�>��O?�.{?1[?�$W>�8�xۭ���OQ�x">E6@?6v�?Qێ?y?}@�>:�>�n)�5�����Q�����ȁ�a�H=�DZ>$�>�Z�>��>,
�=,�Ľر�Ж>�=��=Y*a>�J�>�U�>N��>�'z>�!�<��G?A�>6������\������Q>�[�u?���?��+?G�=�m���E�����Y��>�h�?1�?m**? �T��Y�=4Լ������q��ӷ>ɼ�>�J�>� �=��G=�K>�N�>���>��*�M8���K��?\F?{��=?Ŀ�u��ف��W�����TZ��(������=d���]* ��A����6�=������	Π�_f���;��2?�|�=�ݭ=���=׃�<�[0��%9=Q��=_��;�O=��~��H�6����<p�ƽ��<ޏ<?Ȭ=�p���˾�}?�;I?��+?��C?;�y>�:>��3�ޙ�>f����@?V>ĜP�׈���;�
���� ����ؾ4x׾��c�ʟ��H>baI�*�>e83>�G�=>O�<��=�s=�=r�Q��=�#�=�O�=gg�=���=��>^U>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>N:8>9Q>�R��u1��l[��b�(![��!?��:�8�̾��>��=�2޾Wƾ2=��7>Ahe=Zp��\�p��=�?y��==��g=���>��C> `�=Z���a!�=��M=R��=i{N>	(���:4���*�|�3=�X�=�c>d�%>�|�>s�?��0?��b?�ؼ>�j�7�;!��כ�>i��=V2�>M��=�|E>ɋ�>̎8?��D?A�J?O��>��=S�>�}�>c.+���n����.饾��<��?GV�?`��>@�6<f�?�]s�G>��Ľ�?`/?��	?�>)e�,m˿<C1�v��������>�S�>N���>�Pd�t��=9��=�·�.P�>!.�> �&>���>Y�޽�	�>���>9��=������>�f�	�]�k�=%��;L7Q=�=�_J�QP����c��"����콮�ὡ�ܽ�o�=?� >07>�5�>��x>�g�>:k:=�s��w�>�ި���F�ͭ>�=Ҿ]�G�*ge�/�����9��5���ڧ=�R>�Zc<Mَ�7�>|�=���=���?�6?h��=����˾t����.|�3\X��7=R�3>ي�� @���U���P�MO����>jX<>�{?�;�>uzT�Պ^��{>l1ľ��/��?�7ξH#2�ԽP����o��xm��A�n��;
>�xv?�#�޹>lum?2�J?�U�?�6?�ʯ��j
��o>�rk� +i�I9�����z�#z#?�?5��>*�پ��O���ʾM������>��A��jO�����4�0�`�� 깾ط�>����FҾ3�h������B���v���>�qO?"��?�pb��~�� �M�^��D���@� ?��f?��>ҷ?Y?�W���jƀ�{��=�[n?�`�?���?B(>��=t�����>'��>诛?�?��j?�V�#��>�Xe=�D;>��d�1>I�!>�*>�">�?��?
1 ?�(�����ܾM	 ��@�MyG=t��=�>i>K>��>�-�=���=�ǲ=M�7>��>��|>�A>�V�>.Ɠ>�ُ��w���1?OK'=}��>��1?#�>~�J=�@:���=�_޺��/�mpǽX$��ͼx�=�����=��t���>��ƿRV�?��=���(#?a�۾��=e
�=>vt>�2���>NZ>�WH>=l�>��>���=�7�>ԔU>�J��ef>�j��X#�aOF��d�T���0�>Y����s/������$�����	��Ki�V�y�_l0�Zұ;�Z�?�r�UcL�y �C�8�3�>��>,>4?t���t�-���=)��>���>���`��������~9�?|��?<c>]�>��W?��?�1��3��uZ�3�u��(A��e�a�`��፿����G�
�F��T�_?o�x??yA?cT�<g:z>��?��%�\я�c)�>�/��';�@<=9+�>m)����`��Ӿ3�þ>8�?HF>@�o?�$�?bY?SV�m��&'>�:?�o1?4et?[�1?ـ;?\R��$?ξ3>!G?5m?FT5?��.?��
?=52>���=�����Q'=���
��_ѽ�˽���EE4=�{=1��9�m<c=�<`��[0ټ�;�P��1;�<]�9=��=�o�=7c�>��]?���>��>{�9?�n��7�㖯�/,?��U=�}�Հ��������ޝ>&�k?��?F�Y?w Y>�q@�uJ�J >�n�>�'>a�\>x��>��e�N��ψ=��>��>���=��O��[�����bx����<�	#>��>7|>Ю'>�n��b(z�`�d>��Q��Ѻ�C�S���G���1��vv��]�>��K?��?ڗ�=�]�|C���Df��()?�^<?�EM?<�?��=��۾��9�d�J�*0���>�Y�<��ſ���!��M�:���:�s>�)���ܠ��Xb>���v޾�n�R
J����RAM=�|�RV=,�#�վ�,����=�#
>���}� ����6֪�1J?��j=Gv��kcU�Xt����>�>tܮ>W�:��v��@�l����0�=h��>��:>�c��`��%~G�8�\>�>�PE?�V_?�j�?� ��Os��B�
���Cb���ȼ�?Jy�>�h?SB>��=������U�d�}G���>���>�����G��<���/����$�.��>h8?E�>��?\�R?;�
?��`?�*?�D?Z&�>��������A&?[��?C�=��ԽM�T�w 9�{F����>��)?�B�_��>X�?½?��&?��Q?f�?t�>�� �BD@�)��>�Y�>t�W�Mb��g�_>J�J?қ�>_<Y?�ԃ??�=>(�5��ꢾթ��W�=�>W�2?6#?ǯ?���>���>n���)y<X��>��q?��}?��L?��">g?	WF>p��>~E�=6��>��>�&�>�RB?eK�?i�A?���>8�<.��|�׽�	��E��>�=�p����= o�����҆���W�^��;5��vA#=H ;��z�J<�o�m�>h�r>󴗾��.>Bž^⊾�eD>�	���������Q:�qX�=4=}>R?X�>�"��ߔ=&��>nU�>�W�d�(? �?u?>r��b�̗ھ�M����>�<??���=ۺl�=ٔ�<�v���b=�m?I_?��T�Y'���^?M]{?����2�l:��I
�'C��T?H}?�*��B_�>�A�?�L2?�.�>�M�*�n�\ִ�#d�<�����d����>7�ݕ��o�>��`?��>��?���>���b	��5��I(?�{t?3?w'z?��>0���{8�y������V?���>娧�9?�P�;��ľ�����������j3����[����A���\ �I��/�̽#��=6i?��u?z�r?�?Y?T��b���Z���}��:W�/�������D���G��IF���n�Φ�T꾠ԓ�C�N=�~��pA��2�? g'?�-�]�>0���ﾼ�˾J�B>�^���Et�=�ꋽ�X@='6^=�[e���.��a��� ?^�>T��>�;?g\��=��.1��a7�*���Y�6>���>)�>j��>�Q�:v,�����ɾA�����ӽ�8v>0zc?K�K?еn?�m��(1�I���w�!�[�/��f����B><h>���>�W�П��9&�1Y>���r�����w��O�	���~=@�2?�&�>z��>�N�?�?Qy	�Ui���jx�o�1����<�/�>ii?H>�>e�>� н�� �7��>$�l?pI�>ˋ�>��"�,g� �ǽA6�>�$�>�@�>��&>��=�<�`�U𐿞.���z:�Z��=O�j?�7��֣j��y�>��K?�o���H<�s�>� &�*�����*�.�_�3>��?�g=�8>��Ӿ�&��X}���_��"?�8?fr��nd)��ϊ>oY%??\�>�k�>?��?�b�>A�����S=�?��T?ZrA?W�;?0E�>UKU<����sǽ�����;=]�>޸K>� =h`>[�+��!^������H�=Vv�=�~��ˑ�p��<s1��ߊ�L=9�I>�s����W���'����\����s�����>�ġ���=T�u��[�GS��	���^찻��9��d�pK�;����?���?�Ḿ{�3������l���F��?�̾d�ݼŵ��~Mʽp�ݾ;H ��sϾ��־����'�D.'�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾u1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@G~9?�&�FC�w�3=$c�>�f?ٙ>�{ �����ʧ�,��>%�?8��?��<=��M����=�k?6��8C��%�<��=s��=��=�T�N���D>��>���P�m�u��%[>���>�r9�����P:�+2<	9>N��~N����?�=\��@f���/�'���>�vT?
<�>���=��*? I��Ͽ�[�`b?�c�?i��?F�(?����7�>�jܾM?77?���>� %� Et��~�=�$������侬�U����=<�>� >��,����O�Q�;�����=�/ ���Ŀ��%������<ٶ@<�����������"��̔���c�
	ܽ]��=7y�=�`>>7�}>RsL>(Q>Q�]?*�a?%��>�->�6׽����dɾ�=~[�����9���o�f<���J쾀�پ	�D)����	�þF�;�:��=�S�%��q  ���b�D�D�W�/?<5!>��Ǿh�L�ǈ;<�]ʾg�a���m���˾͔0���l��B�?o�B?09��5�V�z�����`���fW?-��k���!��6w�=P�ټ��=n�>	�=�-���1�DQR��/?��?�ʾ�[Ց�n'.>�����=�,?(?�Ǩ<o��>��%?d� �N��{�Z>U\4>г�>��>%>&F���ֽ2�?��S?!z��̜�ͦ�> ޾�l�z���h=�,>�!6��F��\>��<���7���o.�����<�)W?8ߍ>��)�Q��|ِ�[x&��,>=�x?/�?���>�Kk?�C?�0�<;m���1T��j���u=P�W?p i?s�>����qо�æ���5?%e?/N>+Jh�4b�"�.���X?��n?�D?v1��=�}�;F���&���6?8w?��[����`���d����>QG�>d��>�;����>BN;?�#����V���4���?��@���?tć<�4�b��=4�?b{�><�g��y�����d���,i=��>�e����y��"���3���;?�ф?�p?<〾X����=7ԕ�kZ�?��?(����zf<���l�q��9��<���=� �?r"�W���7���ƾt�
�򦜾ɿ����>^Y@�U��)�>�?8�5⿊RϿ����WоQq���?ׂ�>�ȽG�����j��Su�ƵG�0�H�ڝ��u�>��>�"��������{��o;��������>���>�@T�:��TР��<�F�>��>ٶ�>�"��{�����?�����ͿX����)��X?��?��?�?By<l=x��d~�w�.�G�F?��s?�oZ?�����\�Xb6�&�j?<_���U`�Ď4�]HE��U>Y#3?JD�>��-�Z�|=>��>�c>�#/�1�Ŀ�ض�������?r��?3m꾢��>���?�q+?�j��7��v[����*��t.�::A?�2>����N�!�1=�OҒ��
?�~0?�x��-���o? jT�m����M��Q����6>y�ڼ������׈ƾW����f���r��%�?��@L
�?����n��Y@?]��>i����Yb���(>!r�>��><�;�����>T�&�|�;���= @�a@�?-Չ�碤���=��?��>�م?��=gQ�>��='૾U��;�>�s�=�Un�Ku?DaM?�\�>�p�=L`8��,,���D�v
S�����C��C�>
�b?c�K?J�b>w,����$����ѽI.&����/�;�Ϋ���&�7>>>�>��@���о��?�n���ؿi��u'��04?���>=�?�����t����:_?�s�>F7�*+��$���<�0��?�E�?@�?|�׾B�˼��>��>:H�>8ս���������7>��B?�%��E����o���>���?��@�Ԯ?�i��u?����kGd�{�l�@@���}�t8?>�O7?�����'>�
�>4x�<����j���ol����>���?��?_��>��h?څM���/��{��>�KW?s�?l�.�I��׀�=�?��!�=O��B��+q`?�
@��
@��f?gf��)!Կ▖�/װ�gټ����=��\>I#>\�S���=�J>E�	>2�y����={�>0+�>hgG>0� >8�V>�Q>=���$��1��Cɍ�V�7���D-�K'���U��� �K%ƾf�V��_\v��s���$���l���ڜ���=�#v?��E?�^<?�,�>|D�=w_�>�O'���<�g��Z�>Qm�>{�;?��&?'?�>'>"E���Vi��K��\�Ⱦ�W��N��>���>@{ ?!��>bR�>�]Q>t�q>��>+�=���=1��=䰢�3��=�))>,Q�>�A�>���>�C<>��>9ϴ��1��.�h�w�l̽�?���Y�J��1��f9�������i�=1b.?�{>���?пw����2H?	���e)�ʹ+���>��0?�cW?�>����T�?:>���S�j��`>�+ �$l�q�)�U%Q>Al?��f>/u>��3�Fe8���P�pz���j|>�16?d鶾&H9���u���H��`ݾ2FM>þ>FD�^k�u�����vi���{=�x:?-�?<:���ాE�u�fA���LR>R<\>Y=�l�=�XM>�ic���ƽUH�7g.=���=�^>cL?��&>�=��>����]�D�v��>(LI>:C2>�g??�#?&Xܼ3o�YR��d�+��y>��>�}>��>�RD����=r�>>�T>��.��g�����)>�{�M>yH�r^T���^�ejh=Ϡ��TL�=�]�=E����B�E�&=�~?�⦿v���
쾙�Ž�B?CU?�=6�;�6%��W��,w��T�?�-@�6�?���iU��>?0�? ���&��=\��>���>6)Ⱦ��J�^v?4�ڽ�5������ ���?Q9�?�%9�ݦ��`k���>��#?"
ҾXh�>}x��Z�������u�˶#=b��>�8H?�V��l�O�b>��v
?�?�^�ݩ����ȿ*|v����>S�?���?R�m��A���@�g��>3��?�gY?Toi>�g۾�`Z����>ƻ@?�R?��>�9�a�'���?�޶?ү�?�K>.�? �t?R�><	��}�.�����I���J=��?g�>^��=I���`H���F��-�j�1���m>`�=S�>y*��c��{�=�C���D��N�O�9�>S�f>�gB>-c�>�>�L�>�ő>�X�<B;��ha�����=[7?�'�?b

�"�u�ׁn=b>!>o}ļ�Z�Z�-?R2Ѿˎ)���>?	<?��|?��
?��D>Uj �I��tlٿ���A�c��}�>���>�K0=�M�>�*?i��^�Ͼʭ>=n??$]����<�e�j�O-Y��
�>yI?�k�>�LL=v�0?�8:?N�K>��3?<G�rѲ�9����? �>��'?��g?	}Z?;i �Y�*��8��\0��q΅�Oސ>'x?�8�>X"�>�͋���k�9�>��0�π��_?�i)?�~5�y�?�h�?��D?}?�l�>��&�T�H�vig���>�!?��g�A��P&�G��݃?�C?���>WÒ�J�ս�Dռ���	@���?[\?9:&?��D/a��þK�<Jb"�{�M����;��G�$�>��>�׈�!�=T<>n��=
5m�Q6��f<S_�=:s�>H��=�7��2���n,?/�+�Yہ��0�=h3s��E��r�>�vN>Y�����^?M<��z�H/��FZ��~�Z�p�?^I�?i��?Fᶽ�	h�eQ=?�O�?7%?�>y���� ߾OF��q�'.v�����>v}�>gN�*J徃����ܪ��n��������Kt�>�f�>��?>��>��D>�[�>8[��X -��}���k��b��R���;�=�1�}������9��(#��K������c��>`���8R�>�S	?�Y`>��}><n�>_Dw�0�>EVf>ּs>
��>:�F>��&>���="9�6��KR?������'��达����3B?�od?�1�>]i�����}��~�?���?�r�?:=v>�|h�*+�qm?�<�>���q
? k:=.����<U��t��2��+����>�8׽�:��M�mf�:j
?�.?�(��}�̾<׽��o�>`�?m ?��(�bF�e〿��H�9�r��!�������Fd�)j}�Y��KY��������5���$>��?�e?ǝ��Ҿ�u���PP���.���{>F<�>��n>W�>�0�>SJ�?�3�h�d�~"0�$I���>��o?�g>wW?�@=?�rJ?z�P?�F�>�-�>|R޾�w ?��&= )�>���>)<?�q)?�I"?e?d�?�8�=F�j�܃ ����Ӎ?��A?O*O?ޒ?�i�>��/��=[>�	>�JF��Yݾ���J�;>�}�=߬0�\#�Z>�|�>-F?��K�8�~���Tk>i�7?�,�>���>㿏�.������<G�>P�
?A1�>E��� Kr����	�>���?����=��)>k��=C���d����?�=K�üai�=Ńy���8�Ǚ<���=�@�=��k�X���\�:�P�;���<�Y?�9??��>a��L%�tp����>`[��<��>^.>���g���鰛�����h�>4��?�U�?	9v�8S�=5�>�&�F;@��v����#���[��>��g?;�k?��?Z�x?"_?[a�>m�+�mJ���C�����`��>��-?�ύ>���~3̾�먿1�3�"(?���>\&b���&���+��0ɾ�U½��*>�P(�`&y��c���A�n��<��A����?�;�?D ���4��s�Ai���=��
?B?��>5�>�>5�)�h�����l4>���>-�O??#�>R�O?�;{?�[?�iT>�8��0���ә�-3���!>	@?���?��?�y?Gs�>��>��)�)�SU������N���1W=�Z>���>�(�>��>���=q Ƚ�X����>��b�=��b>)��>���>��>��w>DJ�<��G?f��>�:�����栦���,��pu?ȶ�?��*?m�=����rF�c+�����>!��?J#�?��*?��S���=��������q����>��>�=�>��=ɵJ=�">�d�>R��>�E���e8�-F��D?PJF?^�=f�Ŀv�r�5Z}�ߺ���>f<$���gh�ئ���V��e�=�_��sk�kΤ���D�����N3��'���%l����w��Q?x�j=���=�d�=!�<������<�Q�=�Z<'�=�m���_�<�lk���y��y����9�п<�<1=}g޻��ʾ�{?�G?2�-?!E?>�2>�G�⧛>_�����?dW>M@!��Q��b"A�x���p��2پ4OԾԮb��7��$� >��S���>y�1>Tq�=5Z/<6��=�Iw=��=��D;�)(=���=�/�=F��=Tf�=Z�>&�>�~?�'m�rx���Mg�<����h?�)�>ڵ>���p�?#M�=Fc��5���	&�XQu?:B�?���?x?����>�?��n�$��@�z�P��>���=�W����>�=2}F�L���ɱ&<2�?&o@y�U?	;��TĿD�e>{�7>�n>�R�!n1��[�}�`��.[���!?��:���˾_�>�a�=�ݾ�Tƾ��.=i�6>#�i=��T/\���=ny�&?=`�d=�҈>%tC>�l�=�񯽴G�=v1R=w��=�eP>�O��qU6���)���1=��=�0a>V�%>��>h?�/?l�c?���>��j�}�ϾĿ�T��>�=綰>/F�=��E>$�>7?��D?_HL?�>��=_d�>W	�>
�+��8n����2a���Z�<�Z�?�1�?�P�>�uv<T?��b��=�y(½�?��0?6s?�I�>m.��ۢȿ.�)�}�>�Ĥ$=Q�h>#������;k����>mR�>Wǽ�f�=�߿>�>#5���=�"�>E�=�:�>8>�MV�4�:<t2��Q����<���=A�_��r'�++���7Y=�q�<��<�������'.���MA�� ���C�=/�>T�">���>�Ί=A���� >�헾�xO�tͬ=�ʯ�=�D��Lc���~�v�.�\�:�8=>��Q>Zl���� �?��`>��9>n��?gr?�>����׾����j�c@T��=�=�Q�=âR�	%?�Jo`�{N��;���>{ �>ģ>nl>�,��?�Xp=���ų5��!�>������!��r��fq�E������i�@Q���D?c���Y�=�[~?$�I?W��?1��>�ܘ�w2ؾ#�0>�_����=Nr�_�q�,�����?�&?�W�>ܬ뾐�D���9�2M�h�%?��Roa��`��*���=�j��~�=
���Ѿ�I���������+3�|�b��!�>K�K?���?;�����&#��H�O�޽!�:?Z�??�'�>��>~v-?,�Q�{;�����`�->r��?��?T��?�@���pa=�
��l�>j�?M�?M,�?/�C?(r��'[?��\<�w�=P=��@�>ߓ�=[3K<1>J@,?,�?%��>?)��e���#�۾\�
�1������=��O=�2�>��)>��G>���=���=ڗ�=�G>��>���>��W>��s>_>`(��3��`?!?���=��>t�4??�p>KӍ=�u��#�<�XV�,P,�:��#"��JT߽��=X��<�8N=9��	��>�¿|��?Z'>P.�y?H���j-5>�k>)�����>�H@>��|>娲>Jp�>`y>s>�6>K!Ӿ��>u��)Y!�g#C�}R���Ѿ�sz>uٜ��&����I���XI������j��j��'��m5=�|�<�>�?\����k�c�)�����w?GV�>�6?�ꌾ���Mg>���>���>']������Ǎ�/e���?���?�>���>,�h?�?k����dG���<�F�b�GjL���_�1^�}-��\y����x��g�o?���?�WO?n�v<ð>�с?�+/�������>Vh,�J]��=פ>/����Ͻ��о�����;���� >�v?���?��$?�A}�����u�=G/?��Y?,�?��J?
5�>��=dtk?���>���>MZ�>$�Z?�N�>ٶ�>p��=Σ>��w���5>c�������LD�Z����^;v]�����]�=/�=B�/<:;<�Ӥ�u`<g4}����Ȋ;��U>"�@>տS>9��>�S]?l��>���>>�7?����v8��4��*C/?:=����杊�aס�����>��j?��?5Z?��c>�)A��B��a>ႉ>C7%>�<\>TL�>I���[F�d�=��>��>��=��L��d����	�����;��<J�>�?Z�(>�j=	��=�EؾfՔ�}!�*�Ӿĳ�����ȃ�(Fa�bG���>\Pl?Pu6?�S�<+�Ҿr�Z>�&c��MQ?+?�?�B?�w?w�>J���w�\����=ؚ/><X�<�V,�8ξ������yP�:���ok=W����M<b>�����޾�n�0-J��b羴`P=���ŠU=��־5�~�?��=�	>n���,� �6���ɪ�,=J?�hl=v���JU�w����>U��>��>�^<�Z%v��@�����9�=���>Q�9>-���D�wG���a!�>*�C?�3U?�ވ?�g�M�o��/N�٭��Q��v�V��"?y�>hy�>v�>���=v�����ޔ`�'s@����>_��>����*H�l�����T3�cǋ>G?b�=v
?��W?t�?��]?05?��	?"�>,&���¾��%?W��?�sp��9�<�y�H���K�U�Ž�>Su&?I���?�>N2D?��C?�V�>=@?�6?\�>�T���b�'�b>Q�>��-��쫿0�>�1?<�>>E8?��q?/��>�S�����P>N�>��>j�?�{?�@�>1�>���> k��N�=s�>�d?��?�n?�S�=�; ?W�7>���>e�=��>.��>4?(EO?=�q?�L?�e�>�?�< /���s��	�����)����;ĠX<C��=G���g�z��|
�<��;l�μ��xk�B�L�@`&�Ds0<�_�>��s>
����0><�ľ(P��{�@>҅��wP���ي��:�:ݷ=�>{�?���>,Y#�d��=���>xI�>5���6(?��?�?�!;ˡb���ھM�K�$�>	B?\��=��l�������u���g=��m?��^?'�W�\&��;e^?��]?uF�*��������f�9��UH?&N?N茶X�>`��?J.b?%Ϻ>^P�<jK������k��~���=��>�E#���o�Gi�>��9?��?��i>��S>ؔ��L��)����+?�f�?�u�?�c�?I��>s|��ܿ����"��Y^?�9�>Ʀ�I�"?���'�ξ�ҋ�񾎾��Të��������Ħ���$�[����ֽS0�=j ?s?�?q?��_?ý ��%d���]�C���yV�j������E�ϝD�tC���n���������k��msK=E�]��3�3�?r#?郛�Ȟ�>����˾����;�r>�.۾i�����=M߽x����*=�z���;�]����?�C�>�c�>=6O?�Z�V2F���+��O%�
Z��L>h�>l�z>���>�+0�U�4�au�U|㾴����:�9v>9vc?1�K?�n?�l��(1����7�!���/�4c���B>�c>P��>�W�K��5<&��Y>���r�[���w����	�|�~=R�2?�*�>���>�N�?�?(z	��o��}ox�m�1�Զ�<�3�>3i?�A�>]�>нJ� ���>�l?���>5�>�|��mL!���{�.˽��>��>��>�o>�C-�hC\�|k��H����69��m�=X�h?����[�`�8�>��Q?���:U�V<l�>vFt�V�!�5B�:�'�I�>�Y?9��=��;>��ž6	���{�������&?*M?6iz���Z�M��>���>�^>�4�>{j?��>9�ľ�P;qg(?�kO?cNa?fU?�Y?�>l�ѾQ�����c��=��l>F�=���<N&I>r�ǾH���1�]ݎ>�R
>Ͽ����l=�
R=���=%�?>W��=��G>Ĭ��[N�Ȇ�I��4����4	���Ϻb��=�d�����Wq�����^s]�hFW=O�F�D����8����$�?)R�?�6O��N������F���d��"3#?;2�����u��= r���;��q���v4"��S��P�<�t���'?A���I�ǿY����ܾ|�?�l ?b�y?{"�v�"��v8� >}��<t������������οr��w�^?���>��������>a�>�W>�p>��'���l�<Ȱ?�^-?���>��s�]�ɿh������<2��?@PtA?��(�׹���V=3��>��	?&?>�0��9�ED���s�>�;�?���??�L==�W����%]e?*�;��F��1ܻ���=���="7=w��C�J>���>���,A��ܽ��3>*��>Cd�@�h�]�+'�<e�]>�_ս���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�~���ſ�&����������E=�����.���U_�r��;�X��e"��-�=�c�=N<>���>g;o>�g�>��_?�Fe?�ӥ>iB	>��ɽ*����8��^�q=Jڗ�_���.��̑8�@O��P վg%����X�pl�N�̾�=�/�=~?R����k� ���b�,YF��.?��$>��ʾ/�M��,<Vjʾ�r�����xƥ��̾�l1���m�Z֟?�B?�ꅿ[�V������
��긽��W?�������=3����=멜>_�=���3�r�S�v0?i�?�O���@����+>�� ��G=�+?��?%o<F�>W�$?�)��y���\>��4>�=�>X��>��>���qٽ�i?pT?x�ʜ���>m���
 z�Q�b=�r>N�4�����\>�<o����F����4�<4(W?��>]�)�h��c���C��==��x?�?�+�>]yk?��B?��<L_��P�S�: �GXw=��W?u'i?M�>�t���о���<�5?T�e?f�N>*[h������.��U��"?��n?�\?�"��g{}�,��N���o6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������#��=dǕ��^�?W�?�U��5Fe<��Y�k�(���<�<���=����"�w��.�7���ƾ��
��o��욿�u��>LO@��;t�>��8��/�WMϿM��Zо	"q���?��>=iȽ����z�j�"Ku�]�G��H�)o���/�>�~>�.��5瑾��{�rL;��G�����>������>87S���������9<��>3��>�>��������UǙ?���-ο����R��LzX?Fa�?3}�?�.?C�7<R�v���{����$G?�Xs?tZ?�%�x�\�@�9��k?�f����\��Q3�f~G�IG>��3?a7�>v�-�6�=7P>�>�L>N�/���Ŀ����% �ʎ�?p�?J�龃��>z=�?a�,?%>��y��s���-,��O�;vA?��,>���ˌ#��/@�5q���?A�/?�����з_?x�a�!�p�m�-�d�ƽ�ۡ>��0��h\��v������Ve�n��`<y�y��?�]�?8�?׵�S #��4%?�>���6Ǿj��<р�>�)�>�+N>S#_���u>#���:��h	>��?\}�?�i?򕏿k���*]>��}?c$�>��?�n�=�a�>Gd�=E�y-��k#>�"�=s�>��?��M?L�>FW�=z�8�~/�7[F��GR�d$�=�C� �>��a?ނL?tKb>���2��!��uͽc1��Q��W@��,�r�߽D(5>��=>�>P�D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?PQo���i�B>��?"������L��f?�
@u@a�^?*�ƿ�𒿾Y��V{������/��>��>P7�ɹi>�
+��	�=��Y=���¡�>O��>�3_>V�>^m>82>�Xv�M�"�FS��~&|��9g��Ҧ���쾬`ɾ�ʄ��;aj��;�����Ez$9�I��J�%��7=&�þ�� 9���=@�U?�R?�	p?� ?=Ix�ݍ>9���&�=�j#�v�=*�>�j2?��L?T�*?M!�==����d��`��;7���և�Q��>/I>��>oJ�>*�>�9��I>TN?>Rt�><� >:�'=*캃v=#�N>�(�>��>`��>D<>��>/ϴ��1��]�h�fw�/̽A�?����@�J��1���9��2���k�=�a.?w{>����>пL����2H?|��� )���+���>��0?�cW?��>V��t�T�89>���T�j��_>�- �ށl�ߎ)�%Q>�l?^�f>�%u>c�3�~b8�:�P��v���X|>�46?�嶾�<9��u���H��Tݾ�GM>i��>�8C��h�@���z��gi��{=4x:?=�?r ���簾��u�<���?R>]W\><=;�=dYM>AOc��ƽZH�.=i��=@�^>~W?��+>�=fȣ>�H��C.P����>ՊB>��+>f@?C&%?6��ͱ��,}���-�"w>uI�>1�>�J>�RJ�ɯ=�k�>��a>$�����i��C�?��VW>`�}� |_��Ru���x=;<�����=��='� �?�<��&=�~?���(䈿��!e���lD?U+?| �=F<��"�D ���H��F�?r�@m�?��	�ߢV�?�?�@�?��\��=}�>׫>�ξ"�L��?��Ž9Ǣ�ǔ	�3)#�hS�?��?��/�[ʋ�Al�p6>�^%?��Ӿth�>�x�sZ�������u�@�#=���>�8H?�V����O�w>��v
? ?�^�㩤���ȿ5|v����>P�?���?V�m�bA���@�)��>#��?ogY?�ni>�g۾�_Z�q��>��@?�R?P�>�9�	�'�J�?�޶?﯅?:3I>���?�s?Ϫ�>��w�,\/�4<�������v~=�_;��>ƃ>����sF��Փ��`����j�+����a>�$=�,�> 彆0��؉�=�����R����f�F̷>�p>��I>z��>I� ?,\�>ڙ>�]=̓������Ė��NF?�Ó?����wg��6>��=U���]�?�):?�UL<R���U �>~~x?k?�"^?Vb�>�D������簽��z���=c�>��y>�-�>L�꽔ws>=N���l0��9�>>Ԟ������@��Ū=�B>��>t�?!A�=��?�k?.�s>��;?Wf�>T��(���&�>�>�(?� �?:�	?���A�X��E��L���h���>@eS?>�?���>#e��tx���=��j<����I?��?-�Ⱦ=6C?��?� ?��?�x�>�a=�4�b@��1
�=l�!?�P���A�&��d�5b?d�?M,�>�M����ٽ0ڼIF������?�\?��&?���ma�<-ľ,R�<ǟ�R0��Z�;L(B��X>�>�܇�A��=�g>PA�=�o��F5�-т<ª�=#�>k��=@�5�%���0=,?��G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>'�l���K���ڙ���F��^�Ž�m���h�>�W?;�>���>k>�Kw>�D���6��A���F���x�dx-�nH��G��G<������[�7�A�������6��\�>��B���>h. ?ʈ�>M��>�V&>���<��>=�=�Y>g�>N9\>���>�i�<�YN�5:k��KR?�����'���辠���^3B?�qd?`1�>�i�2��������?���?Rs�?4=v>�~h��,+��n?�>�>7��Kq
?�T:=�;�;�<V��i���2����9��>(E׽� :��M�Pnf�hj
?�/?]����̾e;׽C[��j�=2I�?�zF?%�
�+-J���Z�)�%��w����=�b��-/�ø�j�z���}�|�����/���M�=9�#?<�p?�9�e�uK�`�n���c�mH>�%�>���>�~#?X!�> Q�*o8��a��m�ŬO�z�?��p?�>]OV?�Q/?p�?��[?��>n�~>�����>�}=���>v��>��9?L�@?%NG?;:?"�<?�@>�p����H
���?0?u?���>S]?lL*�3먾ܢ�t0L=�i�����<$��<w�߽�R_�̈́Y<��v>�X?)���8������k>R�7?��>���>����,�����<�>��
?�F�>1 �~r� c��V�>t��?J��Ƀ=��)>���=劅��Һ�Z�=$�����=\5���y;��a<쁿=���=�Kt�����A�:1��;�j�<�u�>1�?P�>�=�>y ���� �e�����=9�V>wT>�>L�پ�k��,���h��Gx>Y�?V��?Q�h=��=���=m��eK�� ���1����< t?�d#?�T?�̒?#>?��"?��>e0���?!��}���V�?g�:?�rU>��ᾫ�Ҿ�﮿�u�4f/?�0?K�e��	�(8�]�Ѿ ��=�:>�R�o�������:K�~iP>��˾�ܽ�^�?_��?��w�M��������x��V?X?aEJ>��>��>G���������-��UI�N��>P�?}!�>��O?�.{?1[?�$W>�8�xۭ���OQ�x">E6@?6v�?Qێ?y?}@�>:�>�n)�5�����Q�����ȁ�a�H=�DZ>$�>�Z�>��>,
�=,�Ľر�Ж>�=��=Y*a>�J�>�U�>N��>�'z>�!�<��G?A�>6������\������Q>�[�u?���?��+?G�=�m���E�����Y��>�h�?1�?m**? �T��Y�=4Լ������q��ӷ>ɼ�>�J�>� �=��G=�K>�N�>���>��*�M8���K��?\F?{��=?Ŀ�u��ف��W�����TZ��(������=d���]* ��A����6�=������	Π�_f���;��2?�|�=�ݭ=���=׃�<�[0��%9=Q��=_��;�O=��~��H�6����<p�ƽ��<ޏ<?Ȭ=�p���˾�}?�;I?��+?��C?;�y>�:>��3�ޙ�>f����@?V>ĜP�׈���;�
���� ����ؾ4x׾��c�ʟ��H>baI�*�>e83>�G�=>O�<��=�s=�=r�Q��=�#�=�O�=gg�=���=��>^U>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>N:8>9Q>�R��u1��l[��b�(![��!?��:�8�̾��>��=�2޾Wƾ2=��7>Ahe=Zp��\�p��=�?y��==��g=���>��C> `�=Z���a!�=��M=R��=i{N>	(���:4���*�|�3=�X�=�c>d�%>�|�>s�?��0?��b?�ؼ>�j�7�;!��כ�>i��=V2�>M��=�|E>ɋ�>̎8?��D?A�J?O��>��=S�>�}�>c.+���n����.饾��<��?GV�?`��>@�6<f�?�]s�G>��Ľ�?`/?��	?�>)e�,m˿<C1�v��������>�S�>N���>�Pd�t��=9��=�·�.P�>!.�> �&>���>Y�޽�	�>���>9��=������>�f�	�]�k�=%��;L7Q=�=�_J�QP����c��"����콮�ὡ�ܽ�o�=?� >07>�5�>��x>�g�>:k:=�s��w�>�ި���F�ͭ>�=Ҿ]�G�*ge�/�����9��5���ڧ=�R>�Zc<Mَ�7�>|�=���=���?�6?h��=����˾t����.|�3\X��7=R�3>ي�� @���U���P�MO����>jX<>�{?�;�>uzT�Պ^��{>l1ľ��/��?�7ξH#2�ԽP����o��xm��A�n��;
>�xv?�#�޹>lum?2�J?�U�?�6?�ʯ��j
��o>�rk� +i�I9�����z�#z#?�?5��>*�پ��O���ʾM������>��A��jO�����4�0�`�� 깾ط�>����FҾ3�h������B���v���>�qO?"��?�pb��~�� �M�^��D���@� ?��f?��>ҷ?Y?�W���jƀ�{��=�[n?�`�?���?B(>��=t�����>'��>诛?�?��j?�V�#��>�Xe=�D;>��d�1>I�!>�*>�">�?��?
1 ?�(�����ܾM	 ��@�MyG=t��=�>i>K>��>�-�=���=�ǲ=M�7>��>��|>�A>�V�>.Ɠ>�ُ��w���1?OK'=}��>��1?#�>~�J=�@:���=�_޺��/�mpǽX$��ͼx�=�����=��t���>��ƿRV�?��=���(#?a�۾��=e
�=>vt>�2���>NZ>�WH>=l�>��>���=�7�>ԔU>�J��ef>�j��X#�aOF��d�T���0�>Y����s/������$�����	��Ki�V�y�_l0�Zұ;�Z�?�r�UcL�y �C�8�3�>��>,>4?t���t�-���=)��>���>���`��������~9�?|��?<c>]�>��W?��?�1��3��uZ�3�u��(A��e�a�`��፿����G�
�F��T�_?o�x??yA?cT�<g:z>��?��%�\я�c)�>�/��';�@<=9+�>m)����`��Ӿ3�þ>8�?HF>@�o?�$�?bY?SV�m��&'>�:?�o1?4et?[�1?ـ;?\R��$?ξ3>!G?5m?FT5?��.?��
?=52>���=�����Q'=���
��_ѽ�˽���EE4=�{=1��9�m<c=�<`��[0ټ�;�P��1;�<]�9=��=�o�=7c�>��]?���>��>{�9?�n��7�㖯�/,?��U=�}�Հ��������ޝ>&�k?��?F�Y?w Y>�q@�uJ�J >�n�>�'>a�\>x��>��e�N��ψ=��>��>���=��O��[�����bx����<�	#>��>7|>Ю'>�n��b(z�`�d>��Q��Ѻ�C�S���G���1��vv��]�>��K?��?ڗ�=�]�|C���Df��()?�^<?�EM?<�?��=��۾��9�d�J�*0���>�Y�<��ſ���!��M�:���:�s>�)��[����b>9�z�߾��m�q�J��W�l�J=3l���P=���ԾR��HL�=G>wG��_e!�A��S����J?�t=�菉�-W�Qߺ�$�>`�>q�>$�9�4#}�0d@�����E�=z��>�9>6+����O�F�W���L�>�&D?F�^?cy�?�:~�:�p���A�_� �Mg�������?&>�>�
?+N>�ٳ=��������d�̯D�d��>W��>5���7F��7������#��r�>O�?�r>�k?C�Q?�U?8Q^?��)?��?���>[d½Iּ��A&?	��?��==�Խ��T�� 9�`F����>��)?L�B�J��>i�?ۼ?��&?��Q?��?��>�� ��C@����>�Y�>��W�[b��c�_>��J?&��>�=Y?�ԃ?g�=>a�5��袾T۩�M�=y>I�2?6#?9�?���>o��>D�����=��>�c?�0�?�o?'��=�?�:2>��>���=���>i��>�?FXO?6�s?��J?ޑ�>帍<8��;9���Cs���O�5ɂ;�rH<��y=Y��34t�%J�:��<I��;_g���G�����D�E ��E��;���>`�H>�̴�&#�>	Ѭ��f���k>��=G�þ�������rǽ��Q>�M?礥>�\ȼ/�>��5>��>&��#�?���>�?ΒG�[�v�)(���0Ž�C�>,�I?r�=?IN��(���)���gc=�nc?�bd?WI��}���W?�wy?���K�ٽ��f����F?��?v(��F�>mۂ?��f?�5�>�Ϲ�:���㢿~ab�l&G��t�%y�>dr�=`�Д>��8?3�>1>%B^=�_��Mnb��5��v?p��?��?���?�B>t�v��y࿞{���I��^?��>w>��c#?�  �4�Ͼ$S�����;�����=@��p��Ŧ$��ԃ�h׽�̼=>�?Is?3[q?x�_?�� �_�c�O/^�9��&gV��#��$���E��(E���C�սn�]`��#�������G=7h.��U;�"��?�5;?[F��F�!?�����u8ܾp#����<���]�=��4="k�>�>�p.�(��ҳt�Z�?�6=��:>�h?]��%�L�S�Q���6�]��`�����>�<3>��1?�(�>s�2�aDz�4�ܜ)�	o>�x>
Xb?��J?w�n?�U���/�끿8k"���O�j?��AB>�>E�>]�K����dX%���=���r�}E�{���?-
��^K=��1?�)�>ǜ�>�w�?��?5_��'���r�YI0���;T��>�sh?��>؍�>c�׽b"�U��>M�?�Y�>7�E>4���(���n������>.->���>��>�(�m#^�+���~��$CQ�nl�=�@l?&i��I8$�`�*>e�*?w��=k��=:�>Z���d2�LE�����§�<W�?'�=jLQ>��оD�
�Բ������FO)?|A?[풾
�*��}>�"?���>H9�>�)�?�2�>�zþ�`���?[�^?�GJ?�UA?EB�>�o= ���qȽ(�&�$m-=�}�>7[>��l=I�=�����\�ǖ��D=���=�ͼ7ٸ���<�|���H<I��<4>VS˿��N���0��C��&��%链����A2�B�ҽ�����))��U2�x�ٽ����ь��"���/�� �?X�?�w�����y�L���3���b�T>{5�s:��ھR#����ԟ���ƾ��R�W�ܗ`��!J�K�'?�����ǿ�����:ܾ! ?�A ?(�y?��@�"���8�.� >�B�<o-����뾩����οH�����^?���>��/��o��>���>T�X>�Hq>����螾�0�<��?�-?��>Ўr�#�ɿO���Ť<���?,�@S{A?�(�H���]V=���>ߍ	?��?>�g1�qL��
���L�>-7�?���?E�M=j�W��
�Vte?��<'�F�WR޻��=���=�O=���J>�V�>{x��XA�\=ܽ��4>z̅>�o"������^�E��<ц]>��ս�(���z?�L�b3\��P �Z���9��=)z?o��>a��=�*?IpB��Pο<H@���K?���?��?>�?7�Ҿ9_U>.���?UUA?��t>L� 
y��� >]ʼJ U�K?��a�T��.�=u?\w�>Iδ��������fֺ�6�="t�� ƿ,^&��P�� =�Z�;�����8̽��^����������T�(e׽�,=���=��C>ď�>R%N>0!K>��b?U�n?��>�>3ȱ������ž�ш��އ�p*)�t���`�¶���]㾢*�W�n*�����ž7%6�'�s=�=Y��������-m��.@��!#?y}
>��̾b�D�l�$=�2Ҿ�맾�LF�2N齫�88�O�l��֥?x�M?��>a���������y�ˏN?��S��ge��y�=���V�<�=�>���=�*޾�'��lD��u0?�[?-����]���"*>�� ���=�+?Ҋ?<nZ<y%�>�J%?��*��/��d[>6�3>�֣>t��>C;	>��6R۽��?ʇT?��������ِ>�c����z��a=�)>775���Х[>�}�<<�G�U�[G��yI�<�O?�?0�f��=齺n}�*��=㛋?^�A?,�H>��?՚?���<,�&�����x|'��R��S/]?��g?���<�t�=�n��)Ѿ��m?A�<?۴����ɾ�iᾧ"?� �9��Y?�d?��?�Ᵹs���5m���
 ��<8?1�v?�^�5|�����9W�C��>�+�>!{�>�m9��z�>�.>?Œ#�"=��A���T#4�~��?+x@#U�?[_:<#��.@�=0?@��>ՄQ��Oľ�Ȱ�������x=O`�>~�����v����m+��r9?��?�Y ?�=��y����=�����Y�?Q�?s��+�g<6+�(l����B��<��=����Z�u��A�7�d�ƾ��
������ �����>�G@.7�)�>��7�&�GCϿ���+�оzqq���?��>� ǽ+%��,�j��[u�ȯG���H�����T�>!�>�蔽�둾T�{��f;�\=�����>���L݈>Q�S��0��Ȃ��5l9<��>���>`��>�w���ӽ�3��?�i��Y=ο���� ���X?�`�?�s�?�r?�/6<ݻv�M�{�)���G?��s?f(Z?+E$�(]��U8�%�j?�_��xU`���4�tHE��U>�"3?�B�>S�-�_�|=�>���>g>�#/�y�Ŀ�ٶ�@���Z��?��?�o���>r��?ss+?�i�8���[����*���+��<A?�2>���I�!�C0=�TҒ�¼
?V~0?{�f.�*
^?3@a�Hi��j(��}ӽ(�>�H���g��=#�ՙ2���e�ư���g�UE�? ,�?��?h$��= ��&?�
�>�阾�8̾��<3d�>�U�> �=>�т��t_>N���4���=���?�8�??�9��`�����>1ـ?�G�>?,�?d�
=)Ċ>�̸>����E�:p0>��@>��=(��>�*[?���>־�;d%��'�Q��JV��c�$�dsE�#8�>c??�.?��)>���_	�<���z�x���h��@�1�f証��3��L�>Mo>-q>>1��\��^�?�O��ؿ�s��>j'��4?_��>y�?��A]u�t��_?�&�>8�3������\�S��?c �?�	?��׾t̼�%>ae�>h	�>�CԽTP���r�7>�pB?Q��4����o�m��>��?[�@ڮ?��h�<�?88��S��u���h@���;	��Y�=ʻ&?&�ž"�=��>A~P=��r� 4��q
f�7�>���?���?`��>C�c?Ģt��N)��;�>�|>`D�?��?�=�쌾*Cc>�P�>��8�$����<�B�?<@�@�k^?K����hֿ�����N��;������=��=r�2>��ٽ9`�=>�7=��8�e9����=5�>��d>�q>#(O>[a;>��)>���+�!�r��K����C�������Z�H��@Xv�bz��3������Q?��a4ý�x���Q�)2&�?`��1�=�[U?�MR?E�o?r] ?�zr�.`>l�����<�t"���=1߆>� 2?�zL?�*?�r�=��a�d�[��lէ�W�����>��J>e��>B��>2��>�Q:��I>Rj@>�)�>La>9s =Yk�lB=��N>���>���>��>qB<>��>^δ�_7��وh��ww��̽W��?-�����J��(���������.�=�D.?U:>���m8пd�t@H?�ٔ���	�+�<�>��0?�^W?ݴ>�찾�rU�,>b����j�Q0>` �nl�Sm)�߄Q>$q?p2o>�Wh>?J2��S6��V�WA�����>��6?�H���&�=�t�<�L��1Ծ�U>.�>^W�;Z����I:{���s��]�=64=?Z�>�{��r������u ��H�,>ֽA>��'<X��=U_>�߼�����R�G��<
>�b>-E?��+>(��=�F�>���ĒO�·�>:B>B�*>�
@?q�$?�{��̙��G��6�,���w>���>�ǀ>u�>NbK�b<�=:��>,Bb>	��܂����0)?���W>�_{���_�z@r��9t=������=/��=C�����;�F�$=�~?�w������Q��T,���TD?��?8��=�2<<k�"�n���h:��%�?v�@	i�?��	�-�V���?VM�?���.��=�)�>�ګ>��;�L�d�?K�ƽC����	��i"��'�?��?ڬ,�fˋ��l���>>I%?EӾRg�>wr��Z����|�u��0#=���>�4H?U���!P��>��v
?N??^�S���}�ȿW}v�4��>��?���?
�m�l>��~	@� t�>£�?�eY?7vi>�X۾DeZ����>��@?R?7�>�3��h'���?�?^��?I>���? �s?YT�>��v��Y/��2�������=S�Z;�d�>�}>����OhF�xړ�:m���j������a>�#$=��>�n��:��*[�=࿋��?���g����>�Kq>G�I>�F�>H� ?�^�>���>�x=�g������&ʖ���K?P��?O���3n����<3��=��^�L&?�I4?� [�u�Ͼ�ר>��\?f��?J[?�^�>����>��!迿:��V��<�K>�2�>OF�>)"���HK>m�Ծ/1D��p�>�ϗ>�����>ھ	+���Ȣ�5C�>�e!?(��>�Ů=� ?�#?^�j>�&�>�_E��9����E�i��>��>pH?��~? ?'Թ�"\3�[	��=桿d�[�0CN>��x?�T?�̕>e������ϽD��CI�������?�sg?Xd�t?�2�?��??}�A?�"f>����ؾ����_�>��!?;��A�;&�����v?#M?F��>���bZֽ��ռ���-m���?&\?�B&?ܕ��/a���¾¯�<�$���a���;�H�f�>I�>����"��=i>A�=�Rm�<}6�L�c<�n�=)��>YC�=�!7�t���=,?!�G�ۃ���=V�r�xD���>�NL>� ���^?)g=���{�r���x���U�� �?���?pk�?�����h��$=?��?(	?*"�>7K���~޾P�ྛKw��x��v���>���>�l���W���֙��hF����Žۖ�b��>��>P�?�l�>#^>s��>�m��"�'���*�~�\��I��7��+��|��:��d���6(��ƾ����y͚>^r�|��>0w?��`>�8>b��>~~�E�>s-T>x>rh�>PR>La3>X+>h�^<2*ɽ�Q?����&$�������rzA?T_?���>t���\���h��[�?��?�5�?Ԣw>��g��+��\?��?�T��M3?��(=��7�<%���,��n��-(�~E�>M�˽��:�}^K�(�`�7?{�?$qN�`�̾�ٽ����(�n=�M�?n�(?��)���Q�žo�ӸW� S�����6h��i����$�.�p��쏿�^��+%��}�(�:x*=�*?B�?Ό���� ���&k�r?�8cf>�>b#�>k�>xrI>��	���1�[^��L'�/����R�>�[{?Hq�>��H?ь<?�\P?�K?��>��>����]��>k�
<�X�>v:�>��8?��-?�?0?�?�+?
�b>��`�����ؾ`?P�?P�?(U?I?�
������"�����n���w�����V�w=]0�<6c׽2�i���X=KS>�X?b����8�����uk>T�7?��>d��>����,����<��>�
?�F�>` �C~r�c�2V�>���?% �̄=i�)>m��=���V�Һ�Z�=������=3���y;�d<y��=���=�/t�����R�:��;�h�<[h?�~-?)�>�>�;���>��=���!�>�b�>�ƽ>+��>�/���֎��R��4bp����>��?��?O�<��=� �=⶧�a-��.�w侜g�ʟ?TZT?@{4?�?�Il?�\3?o]���><��B���P���"����?t ,?Ƃ�>�����ʾZ�y�3���?gY?�9a�̷�L?)�=�¾8�Խ��>�K/�!~����D�kQ����Et����?]��?V@���6�J����~k��E�C?��>Pi�>��>�)�R�g��"��;>��>�R?�>dV?L��?LEp?��>�ཱྀ����P����ɾۮ�m��>�T?[��?x3�?���>~�'�c����۲�J>|>�%���9�=��ľ�Q=9A�>9@f>:p*?��a>�W?��3�=^�=-�ǾL��=z��>�$]>J�>$�>���=/���'<?>�?�����`���(���1���e	>sGk?w]t?G�?�sE=4��P�h�_	�2��>�Ȟ?"��?9$M?/]����4=�#�<�=5�� ��ڰ>�t?Ӷ>��>_:&>��#>^/?��> �:�-�t�L�J��N�?+�?S�X>�˿Ӂx���~������^M��~��B<���&��!��j�>!�g�B����)��}i�E��Vߓ�ꈯ��o����~����>� =��=��>s{%=�,�� /<$`=���<�X	;��}����<9W�cӢ;+F��#껴�<M�=�#����˾K�}?�7I?��+?��C?V�y>�:>s�3�J��>8R��D=?�)V>��P�������;�M����"����ؾ�׾d�ɟ��C>�YI�@�>b;3>pJ�='/�<�+�=�"s=;ʎ=�Q��=X.�=f�=x�=���=/�>�D>�n?N�k�e����/D�c�^�P�N?뽮>7;�=a���$?��=?d��	}������|?� �?>3�?���>ʑd���>�b�j�M=��I>0�x���
>��>����B^�>S��>����/��ٜr�J�?��@�C?k�v�*
ȿ�x>��7>)%>��R���1���\���b�rZ��!?�G;��M̾�3�>��=V.߾�ƾ?_.=��6>5b=�n��T\�L��=��z�g�;=l=�ω>�D>E�=?!��u�=��I=l��=H�O>������7��,�4=�
�=��b>J&>�e�>�s�>z?��n?���>'2������&ѾiZ=Ӥ��`�>��ƽ���>g>?��0?�5?P+?o�>���=�F�>��4>�sV�~�F�|��]�����=�K�? :|?�C4>�=��&�*eA���E�J,k�eh(?2?-j�>b��=�v��Eտ��[	1��(��m�=��?v*�I��>���>7�[>���=�>� �=9c�>م�=j�>x>�=�
�<J5�>\�3��4͸��U>|���<�f=���5��=R�=��<=w#��i�:��+�ߡ��Y?ż��b=m�A='��;��<c��=A��>�?>���>	��=���wD/>������L�rĿ=	J���+B�-4d��H~�/�T6�5�B>�:X>ˀ��,4����?E�Y>�n?>��?7Au?%�>U!�1�վ:Q��Ee�SS�ɸ=��>��<�^z;��Y`�S�M�C{Ҿ��>;�>��>�.l>G�+�^?�Q\v=���m85����>@Y���Z����|(q��C��M��?-i���𺱫D?-B���.�=�}?�zI?�؏?H��>$]����ؾZ�/>�ԁ�i�= �[�p�7����?��&?�{�>�I���D����n���p��>�Y���?B��n��u$�ʈX�Lb����>���]6��.#2�8����t��dA�O���C�>ge@? 8�?�K� ]r�m:����݉G=`V?�jb?y��>���>��>b�����YR���� >C�|?�?&��?��5>ؿ=�v��@�>�	?%��?K��?*�r?+B��5�>��[; >����9"�=��>���=*��=C�?��	?��
?�H����	�^��m/�	^����<\6�=���>�u�> �n>o)�=�>h=�U�=c~Z>V��>��>��e>4ڢ>�C�>|^��t� �-`S?�z>�
'>�\?�t7>%$ؼȧ9���)>Cӝ������h�ཁM�y��=�~=>z��=O�	�'@|>����wR�?�ȃ>���r9?$��}i���ʆ>��=��I����>,�7>l�D>Z�><��>i�>��q>H�L>��ʾ/M>����-�Q�8�x�\��Iʾ�/e>p��f�9���ѹ���']����7	��_j�������B���;!�?�)��ř`���.�l�c�?�r�>��2?���ƽ]��=.[�>/K�>�����鑿Qʅ�M�о��?���?
Rc>�)�>N�W? �?�1�3�3�eKZ�X�u�eA���d�M�`�qٍ�����
�o�����_?A�x?gjA?Pҍ<��y>$��?��%������>��.��;�ˏ==rA�>�����`�}hӾ��þ���[�E>+zo?-!�?��?XV��m��'>��:?Λ1?�Ot?��1?i�;?�����$?co3>�F?�q?8N5?��.?'�
?Q2>
�=�����'=�6���g�ѽ�~ʽi��X�3=�^{=~a͸� <�=���<��ʣټ#�;\%��B%�<:=o�=
�=�>˕]?�i�>���>W�7?X��#O8������	/?�;=V΂����	�����>n�j?��?�jZ?��c>>&B��C�/Z>&�>R0&>�r\>JU�>�f"E��$�=��>)�>!i�=
XO�g�߶	�DV��m�<W>8��>be)>X��=ETx>�s��?�k����>�σ� �����J���b���.��%d�d��>�Y?O2,?�Y>�>Ҿ!��ݝg��?�[�?/[G?"XQ?��X>"O�S�?�I���H�<6Լؽ�>,�)�c���{����.��X[>Vs�>����ܠ��Xb>���v޾�n�R
J����RAM=�|�RV=,�#�վ�,����=�#
>���}� ����6֪�1J?��j=Gv��kcU�Xt����>�>tܮ>W�:��v��@�l����0�=h��>��:>�c��`��%~G�8�\>�>�PE?�V_?�j�?� ��Os��B�
���Cb���ȼ�?Jy�>�h?SB>��=������U�d�}G���>���>�����G��<���/����$�.��>h8?E�>��?\�R?;�
?��`?�*?�D?Z&�>��������A&?[��?C�=��ԽM�T�w 9�{F����>��)?�B�_��>X�?½?��&?��Q?f�?t�>�� �BD@�)��>�Y�>t�W�Mb��g�_>J�J?қ�>_<Y?�ԃ??�=>(�5��ꢾթ��W�=�>W�2?6#?ǯ?���>���>n���)y<X��>��q?��}?��L?��">g?	WF>p��>~E�=6��>��>�&�>�RB?eK�?i�A?���>8�<.��|�׽�	��E��>�=�p����= o�����҆���W�^��;5��vA#=H ;��z�J<�o�m�>h�r>󴗾��.>Bž^⊾�eD>�	���������Q:�qX�=4=}>R?X�>�"��ߔ=&��>nU�>�W�d�(? �?u?>r��b�̗ھ�M����>�<??���=ۺl�=ٔ�<�v���b=�m?I_?��T�Y'���^?M]{?����2�l:��I
�'C��T?H}?�*��B_�>�A�?�L2?�.�>�M�*�n�\ִ�#d�<�����d����>7�ݕ��o�>��`?��>��?���>���b	��5��I(?�{t?3?w'z?��>0���{8�y������V?���>娧�9?�P�;��ľ�����������j3����[����A���\ �I��/�̽#��=6i?��u?z�r?�?Y?T��b���Z���}��:W�/�������D���G��IF���n�Φ�T꾠ԓ�C�N=�~��pA��2�? g'?�-�]�>0���ﾼ�˾J�B>�^���Et�=�ꋽ�X@='6^=�[e���.��a��� ?^�>T��>�;?g\��=��.1��a7�*���Y�6>���>)�>j��>�Q�:v,�����ɾA�����ӽ�8v>0zc?K�K?еn?�m��(1�I���w�!�[�/��f����B><h>���>�W�П��9&�1Y>���r�����w��O�	���~=@�2?�&�>z��>�N�?�?Qy	�Ui���jx�o�1����<�/�>ii?H>�>e�>� н�� �7��>$�l?pI�>ˋ�>��"�,g� �ǽA6�>�$�>�@�>��&>��=�<�`�U𐿞.���z:�Z��=O�j?�7��֣j��y�>��K?�o���H<�s�>� &�*�����*�.�_�3>��?�g=�8>��Ӿ�&��X}���_��"?�8?fr��nd)��ϊ>oY%??\�>�k�>?��?�b�>A�����S=�?��T?ZrA?W�;?0E�>UKU<����sǽ�����;=]�>޸K>� =h`>[�+��!^������H�=Vv�=�~��ˑ�p��<s1��ߊ�L=9�I>�s����W���'����\����s�����>�ġ���=T�u��[�GS��	���^찻��9��d�pK�;����?���?�Ḿ{�3������l���F��?�̾d�ݼŵ��~Mʽp�ݾ;H ��sϾ��־����'�D.'�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >\C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾u1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@G~9?�&�FC�w�3=$c�>�f?ٙ>�{ �����ʧ�,��>%�?8��?��<=��M����=�k?6��8C��%�<��=s��=��=�T�N���D>��>���P�m�u��%[>���>�r9�����P:�+2<	9>N��~N����?�=\��@f���/�'���>�vT?
<�>���=��*? I��Ͽ�[�`b?�c�?i��?F�(?����7�>�jܾM?77?���>� %� Et��~�=�$������侬�U����=<�>� >��,����O�Q�;�����=�/ ���Ŀ��%������<ٶ@<�����������"��̔���c�
	ܽ]��=7y�=�`>>7�}>RsL>(Q>Q�]?*�a?%��>�->�6׽����dɾ�=~[�����9���o�f<���J쾀�پ	�D)����	�þF�;�:��=�S�%��q  ���b�D�D�W�/?<5!>��Ǿh�L�ǈ;<�]ʾg�a���m���˾͔0���l��B�?o�B?09��5�V�z�����`���fW?-��k���!��6w�=P�ټ��=n�>	�=�-���1�DQR��/?��?�ʾ�[Ց�n'.>�����=�,?(?�Ǩ<o��>��%?d� �N��{�Z>U\4>г�>��>%>&F���ֽ2�?��S?!z��̜�ͦ�> ޾�l�z���h=�,>�!6��F��\>��<���7���o.�����<�)W?8ߍ>��)�Q��|ِ�[x&��,>=�x?/�?���>�Kk?�C?�0�<;m���1T��j���u=P�W?p i?s�>����qо�æ���5?%e?/N>+Jh�4b�"�.���X?��n?�D?v1��=�}�;F���&���6?8w?��[����`���d����>QG�>d��>�;����>BN;?�#����V���4���?��@���?tć<�4�b��=4�?b{�><�g��y�����d���,i=��>�e����y��"���3���;?�ф?�p?<〾X����=7ԕ�kZ�?��?(����zf<���l�q��9��<���=� �?r"�W���7���ƾt�
�򦜾ɿ����>^Y@�U��)�>�?8�5⿊RϿ����WоQq���?ׂ�>�ȽG�����j��Su�ƵG�0�H�ڝ��u�>��>�"��������{��o;��������>���>�@T�:��TР��<�F�>��>ٶ�>�"��{�����?�����ͿX����)��X?��?��?�?By<l=x��d~�w�.�G�F?��s?�oZ?�����\�Xb6�&�j?<_���U`�Ď4�]HE��U>Y#3?JD�>��-�Z�|=>��>�c>�#/�1�Ŀ�ض�������?r��?3m꾢��>���?�q+?�j��7��v[����*��t.�::A?�2>����N�!�1=�OҒ��
?�~0?�x��-���o? jT�m����M��Q����6>y�ڼ������׈ƾW����f���r��%�?��@L
�?����n��Y@?]��>i����Yb���(>!r�>��><�;�����>T�&�|�;���= @�a@�?-Չ�碤���=��?��>�م?��=gQ�>��='૾U��;�>�s�=�Un�Ku?DaM?�\�>�p�=L`8��,,���D�v
S�����C��C�>
�b?c�K?J�b>w,����$����ѽI.&����/�;�Ϋ���&�7>>>�>��@���о��?�n���ؿi��u'��04?���>=�?�����t����:_?�s�>F7�*+��$���<�0��?�E�?@�?|�׾B�˼��>��>:H�>8ս���������7>��B?�%��E����o���>���?��@�Ԯ?�i��u?����kGd�{�l�@@���}�t8?>�O7?�����'>�
�>4x�<����j���ol����>���?��?_��>��h?څM���/��{��>�KW?s�?l�.�I��׀�=�?��!�=O��B��+q`?�
@��
@��f?gf��)!Կ▖�/װ�gټ����=��\>I#>\�S���=�J>E�	>2�y����={�>0+�>hgG>0� >8�V>�Q>=���$��1��Cɍ�V�7���D-�K'���U��� �K%ƾf�V��_\v��s���$���l���ڜ���=�#v?��E?�^<?�,�>|D�=w_�>�O'���<�g��Z�>Qm�>{�;?��&?'?�>'>"E���Vi��K��\�Ⱦ�W��N��>���>@{ ?!��>bR�>�]Q>t�q>��>+�=���=1��=䰢�3��=�))>,Q�>�A�>���>�C<>��>9ϴ��1��.�h�w�l̽�?���Y�J��1��f9�������i�=1b.?�{>���?пw����2H?	���e)�ʹ+���>��0?�cW?�>����T�?:>���S�j��`>�+ �$l�q�)�U%Q>Al?��f>/u>��3�Fe8���P�pz���j|>�16?d鶾&H9���u���H��`ݾ2FM>þ>FD�^k�u�����vi���{=�x:?-�?<:���ాE�u�fA���LR>R<\>Y=�l�=�XM>�ic���ƽUH�7g.=���=�^>cL?��&>�=��>����]�D�v��>(LI>:C2>�g??�#?&Xܼ3o�YR��d�+��y>��>�}>��>�RD����=r�>>�T>��.��g�����)>�{�M>yH�r^T���^�ejh=Ϡ��TL�=�]�=E����B�E�&=�~?�⦿v���
쾙�Ž�B?CU?�=6�;�6%��W��,w��T�?�-@�6�?���iU��>?0�? ���&��=\��>���>6)Ⱦ��J�^v?4�ڽ�5������ ���?Q9�?�%9�ݦ��`k���>��#?"
ҾXh�>}x��Z�������u�˶#=b��>�8H?�V��l�O�b>��v
?�?�^�ݩ����ȿ*|v����>S�?���?R�m��A���@�g��>3��?�gY?Toi>�g۾�`Z����>ƻ@?�R?��>�9�a�'���?�޶?ү�?�K>.�? �t?R�><	��}�.�����I���J=��?g�>^��=I���`H���F��-�j�1���m>`�=S�>y*��c��{�=�C���D��N�O�9�>S�f>�gB>-c�>�>�L�>�ő>�X�<B;��ha�����=[7?�'�?b

�"�u�ׁn=b>!>o}ļ�Z�Z�-?R2Ѿˎ)���>?	<?��|?��
?��D>Uj �I��tlٿ���A�c��}�>���>�K0=�M�>�*?i��^�Ͼʭ>=n??$]����<�e�j�O-Y��
�>yI?�k�>�LL=v�0?�8:?N�K>��3?<G�rѲ�9����? �>��'?��g?	}Z?;i �Y�*��8��\0��q΅�Oސ>'x?�8�>X"�>�͋���k�9�>��0�π��_?�i)?�~5�y�?�h�?��D?}?�l�>��&�T�H�vig���>�!?��g�A��P&�G��݃?�C?���>WÒ�J�ս�Dռ���	@���?[\?9:&?��D/a��þK�<Jb"�{�M����;��G�$�>��>�׈�!�=T<>n��=
5m�Q6��f<S_�=:s�>H��=�7��2���n,?/�+�Yہ��0�=h3s��E��r�>�vN>Y�����^?M<��z�H/��FZ��~�Z�p�?^I�?i��?Fᶽ�	h�eQ=?�O�?7%?�>y���� ߾OF��q�'.v�����>v}�>gN�*J徃����ܪ��n��������Kt�>�f�>��?>��>��D>�[�>8[��X -��}���k��b��R���;�=�1�}������9��(#��K������c��>`���8R�>�S	?�Y`>��}><n�>_Dw�0�>EVf>ּs>
��>:�F>��&>���="9�6��KR?������'��达����3B?�od?�1�>]i�����}��~�?���?�r�?:=v>�|h�*+�qm?�<�>���q
? k:=.����<U��t��2��+����>�8׽�:��M�mf�:j
?�.?�(��}�̾<׽��o�>`�?m ?��(�bF�e〿��H�9�r��!�������Fd�)j}�Y��KY��������5���$>��?�e?ǝ��Ҿ�u���PP���.���{>F<�>��n>W�>�0�>SJ�?�3�h�d�~"0�$I���>��o?�g>wW?�@=?�rJ?z�P?�F�>�-�>|R޾�w ?��&= )�>���>)<?�q)?�I"?e?d�?�8�=F�j�܃ ����Ӎ?��A?O*O?ޒ?�i�>��/��=[>�	>�JF��Yݾ���J�;>�}�=߬0�\#�Z>�|�>-F?��K�8�~���Tk>i�7?�,�>���>㿏�.������<G�>P�
?A1�>E��� Kr����	�>���?����=��)>k��=C���d����?�=K�üai�=Ńy���8�Ǚ<���=�@�=��k�X���\�:�P�;���<�Y?�9??��>a��L%�tp����>`[��<��>^.>���g���鰛�����h�>4��?�U�?	9v�8S�=5�>�&�F;@��v����#���[��>��g?;�k?��?Z�x?"_?[a�>m�+�mJ���C�����`��>��-?�ύ>���~3̾�먿1�3�"(?���>\&b���&���+��0ɾ�U½��*>�P(�`&y��c���A�n��<��A����?�;�?D ���4��s�Ai���=��
?B?��>5�>�>5�)�h�����l4>���>-�O??#�>R�O?�;{?�[?�iT>�8��0���ә�-3���!>	@?���?��?�y?Gs�>��>��)�)�SU������N���1W=�Z>���>�(�>��>���=q Ƚ�X����>��b�=��b>)��>���>��>��w>DJ�<��G?f��>�:�����栦���,��pu?ȶ�?��*?m�=����rF�c+�����>!��?J#�?��*?��S���=��������q����>��>�=�>��=ɵJ=�">�d�>R��>�E���e8�-F��D?PJF?^�=f�Ŀv�r�5Z}�ߺ���>f<$���gh�ئ���V��e�=�_��sk�kΤ���D�����N3��'���%l����w��Q?x�j=���=�d�=!�<������<�Q�=�Z<'�=�m���_�<�lk���y��y����9�п<�<1=}g޻��ʾ�{?�G?2�-?!E?>�2>�G�⧛>_�����?dW>M@!��Q��b"A�x���p��2پ4OԾԮb��7��$� >��S���>y�1>Tq�=5Z/<6��=�Iw=��=��D;�)(=���=�/�=F��=Tf�=Z�>&�>�~?�'m�rx���Mg�<����h?�)�>ڵ>���p�?#M�=Fc��5���	&�XQu?:B�?���?x?����>�?��n�$��@�z�P��>���=�W����>�=2}F�L���ɱ&<2�?&o@y�U?	;��TĿD�e>{�7>�n>�R�!n1��[�}�`��.[���!?��:���˾_�>�a�=�ݾ�Tƾ��.=i�6>#�i=��T/\���=ny�&?=`�d=�҈>%tC>�l�=�񯽴G�=v1R=w��=�eP>�O��qU6���)���1=��=�0a>V�%>��>h?�/?l�c?���>��j�}�ϾĿ�T��>�=綰>/F�=��E>$�>7?��D?_HL?�>��=_d�>W	�>
�+��8n����2a���Z�<�Z�?�1�?�P�>�uv<T?��b��=�y(½�?��0?6s?�I�>m.��ۢȿ.�)�}�>�Ĥ$=Q�h>#������;k����>mR�>Wǽ�f�=�߿>�>#5���=�"�>E�=�:�>8>�MV�4�:<t2��Q����<���=A�_��r'�++���7Y=�q�<��<�������'.���MA�� ���C�=/�>T�">���>�Ί=A���� >�헾�xO�tͬ=�ʯ�=�D��Lc���~�v�.�\�:�8=>��Q>Zl���� �?��`>��9>n��?gr?�>����׾����j�c@T��=�=�Q�=âR�	%?�Jo`�{N��;���>{ �>ģ>nl>�,��?�Xp=���ų5��!�>������!��r��fq�E������i�@Q���D?c���Y�=�[~?$�I?W��?1��>�ܘ�w2ؾ#�0>�_����=Nr�_�q�,�����?�&?�W�>ܬ뾐�D���9�2M�h�%?��Roa��`��*���=�j��~�=
���Ѿ�I���������+3�|�b��!�>K�K?���?;�����&#��H�O�޽!�:?Z�??�'�>��>~v-?,�Q�{;�����`�->r��?��?T��?�@���pa=�
��l�>j�?M�?M,�?/�C?(r��'[?��\<�w�=P=��@�>ߓ�=[3K<1>J@,?,�?%��>?)��e���#�۾\�
�1������=��O=�2�>��)>��G>���=���=ڗ�=�G>��>���>��W>��s>_>`(��3��`?!?���=��>t�4??�p>KӍ=�u��#�<�XV�,P,�:��#"��JT߽��=X��<�8N=9��	��>�¿|��?Z'>P.�y?H���j-5>�k>)�����>�H@>��|>娲>Jp�>`y>s>�6>K!Ӿ��>u��)Y!�g#C�}R���Ѿ�sz>uٜ��&����I���XI������j��j��'��m5=�|�<�>�?\����k�c�)�����w?GV�>�6?�ꌾ���Mg>���>���>']������Ǎ�/e���?���?�>���>,�h?�?k����dG���<�F�b�GjL���_�1^�}-��\y����x��g�o?���?�WO?n�v<ð>�с?�+/�������>Vh,�J]��=פ>/����Ͻ��о�����;���� >�v?���?��$?�A}�����u�=G/?��Y?,�?��J?
5�>��=dtk?���>���>MZ�>$�Z?�N�>ٶ�>p��=Σ>��w���5>c�������LD�Z����^;v]�����]�=/�=B�/<:;<�Ӥ�u`<g4}����Ȋ;��U>"�@>տS>9��>�S]?l��>���>>�7?����v8��4��*C/?:=����杊�aס�����>��j?��?5Z?��c>�)A��B��a>ႉ>C7%>�<\>TL�>I���[F�d�=��>��>��=��L��d����	�����;��<J�>�?Z�(>�j=	��=�EؾfՔ�}!�*�Ӿĳ�����ȃ�(Fa�bG���>\Pl?Pu6?�S�<+�Ҿr�Z>�&c��MQ?+?�?�B?�w?w�>J���w�\����=ؚ/><X�<�V,�8ξ������yP�:���ok=W�!��'a>�
��߾t�l��L�;���Cc=Э���m=lO��3Ծ����/\�=)�>����ɺ ��7���1��`�J?Q�{=Eݪ���Y�𧽾�>�̙>@ڪ>�uH�3Y���@�e1�����=�l�>�8>9*��Ik�U�H��P���>y I?�=f?�A?xx��\�l�%;A�Hs�����yr��?��>�?��S>W�=����B���g�l�O�\�>���>b~�G�3��Y�����9��>7p?�O>l�?�V?��?��\?��2?N�?e�>����������%?�0�?�y�={��nN��17��F��N�>O�(?�lI�zЗ>�Y?%�?2�)?��R?�?��>"���R?��U�>@=�>09X��ӯ��j>%�J?`��>H�V?aN�?��=>��5�N��^������=��>E"4?�$?7�? ��>���>����x>�)?h�s?�p�?�o?��/�)k<?�T@>���>� �<x��>Ӛ2?�.
?�GL?p��?i�?~M?3S<��Ͻ����}UȽ[¹�N��=��]>:x%>�b9�§,=\�=Aۊ�%ʄ=�؎=��+�f��S �s�=Ƚ&�4�>��m>�i��x�1>��¾d����A>oc��e���Ǉ���9���=��}>�� ?$-�>�u!�d��=� �>��>f���'?D�?�?�[f;��b���ݾcN���>�A?H\�=n�l�����;	v�W�q=Hjm?��^?�`W��w����b?��]?�r�=� "ľ��a����ݬO?g�
?�G���>)�~?��q?V��>�e�n����sZb��Jj��i�=�e�>_���d�{ߞ>��7?�h�>�2d>��=�۾Sw�њ��j?��?�?*�?C+>��n�_"�
���e��o1?E�>�����$?=�����&��l@��:�Ӿ/ᾪ;���׽��|��-ޔ�o�4�I �ö�i?�5�?��\?^�1?]v���z~�c<}�>��(�I[��%F�1
S��%J�P�J�D���ɂ2�k�;F\��45�=����sE�̞�?�&?������>R&��X�ϾCȾ�$v>i����D�T=Ɗ���X=�P4=��k����$��u�!?I��>c�>z�3?Q�V�ƘA�{�8��'6�v���s0>��>�Ky>ܴ>P�ռ�V㽇rǽ<6��]I������m�v>�fl?](`?!�S?�;�!�%���|��*�$d~�,Ծq$�>!�=�~l>��#��k5�F"#��C-��(x��&#���\�z��<7[>?ܨ>���>�(�?�?�����,I�3�Y�6����>���>�Nz?��?���>��ֽ�$����>q�l?�(�>`�>���G!���{�6>νݐ�>ß�>��>�n>�-��\��{������9��(�=�<h?de��o�`�G�>!�Q?0Z9��@<�u�>�Ht�Ϣ!�����&�>	>mv?*�='=<>��ľ(��<�{�\���(?��?����c+�v�z>�#?>��>М�>�T�?��>+H��+�ػ\?�^?��I?�w@?���>R�=2���8˽�	+��+=��>�\>�w=:�=���?�Z�!\(�7�Y=}i�=�j�����j:<=�ü��<��=�,>e�ٿ�L�`׾���5��W���ӊ����������罛*��/����ڀ�M��a��WT���b�o?���h����?�h�?;ۗ�;l���ʙ�\ր�F����>�Hu��2��G,��J�_͞��tᾯ⡾�9���L���h��f�4�>?W�����οa����ྪ7?7�>�S?�r������(��E)>��Ͻ�D;���ξ�t��Ͽ�6����3?8��>����=��>oZ9>��>%E�>đʾ_"���>��?���>��?M�����ʿ����L¼�d�?��@�mA?߫(�3��O�]=��>�=	?M@@>҆1����氾ע�>+�?v�?�aN=�qW��y�_�e?ݟ<��F���ֻ���=蜧=D=����aJ>�ʒ>>|��MB�x�ܽ�4>���>V�����]�홲<��\>E�ֽ?����Ԅ?r{\��f�d�/��T���Z>��T?r+�>�3�=ͱ,?�5H�}Ͽ��\�q)a?60�?¦�?��(?�ڿ��՚>��ܾӉM?�B6?���>�b&���t��s�=�r�i?��`��&(V���=���>�~>��,�m���O�L@�����=CA��oƿ��!�Q�P�,=����w��u���������#��KX�����/Y=���=b�D>��>��V>әf>f�U?Q]i?���>}�>� Խ�q��U�Ѿ���Ӏ��d��Ս�(l!�����D��ҾV��I�R���#ʾS��j��E�M�e�z�NY��������k���M?�m=�+$;(�k�~��=�+!����{>0��<26��R�.���s�h؟?�7]?yi��A�n�d�0���Q��A,�
�>z���6�1���i���a���(Z=%ִ>'>�=�~ ��S]�W�}�ZP0?�E?�l���掾2;*>#����=�:+?+?4�T<j&�>ah%?��'�]z佭!\>��6>�פ>���>�	>�k��r�ܽ̃?r�T?"5�����?u�>lҽ�j|�ׅa=�>�4��ټDJ]>�<�M���db�,����<�(W?;��>��)����a��a��Z==��x?g�?..�>{k?w�B?nߤ<�h���S���+]w=��W?�)i?�>���EоȀ��S�5?4�e?��N>Wch������.��T��#?%�n?_?j���Ew}�O�����n6?��v?s^�xs�����L�V�e=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?n�;<��T��=�;?m\�> �O��>ƾ�z������.�q=�"�>���ev����R,�f�8?ݠ�?���>�������[ >�}����?? �?pâ�Ixh<���Ye��ﾱ�\Po<�]꽣SY�����4_E�5dվ�s��*����L�dRw>��@�"'���>��B��߿8�˿7��P����4����>
G�>�}"��ҟ�29n��Z��ޱP���L�,�x���>pk%>�Ǹ�����P�{�q++���=|��>κQ�v�>�z/�庾�/���Ǖ<c�>�.�>�Sg>� ������^�?�{��ʿ�؝���H�_?B�? ��?E5#?��I���4��φ���y:��M?�Tv?�V?=*<��G�4���]�p?J���ّ\�kbD���]�f��=��9?(��>��J��3�=�>�$�>��=�O��
���[���%�KÓ?��?�q�? ��?d�1?�R>����)�A�Q�;����O�&?�>���i��)������	?��?]`����]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?@$�>��?n�=�a�>dc�=�𰾃�,��k#>	"�=��>�9�?b�M?�K�>�W�=K�8�u/�A[F��GR�<$�:�C���>g�a?ÂL?�Kb>3��U2�I!�uͽtd1��K��W@���,��߽�(5>��=>E>��D��Ӿ��?Mp�9�ؿ j�� p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>E�Խ����\�����7>1�B?[��D��u�o�z�>���?
�@�ծ?ji��	? ��P���`~�����7�S��=;�7?t0�(�z>I��>Q�=�nv�������s�S��>wB�?n{�?��>"�l?�o�P�B�a�1=�L�>2�k?)s?�uo���&�B>I�?Z�����L�' f?��
@`u@��^?.	Ŀ +��F���᩾���	��=I�M>�x.���=j��<���=�H�=��>	��>�T>�"6>,6�>!�>��>��{�S�����|���r
8�w!#�]>7�0���uG��X1�H�"���8��i���H�7R�ZmX�&w�d{��5��=��=�U?�R?Kp?�� ?;�x��f>����E�=9�#��B�=�!�>}s2?b�L?<�*?�ד=������d�_���6���Ǉ��b�>�YI>���>�U�>�>���9�J>�4?>�g�>'*>MH(=\к�j=�-O>Uj�>U��>�~�>Ԍ�>j�>�ʿkʨ�n$W�����8RA���?��Ծ��-�����*����fl(���;?.�>�4��Uտ8S��1�H?�΅������d��ļ��P?��I?7.���þo���>y����)Q�rၽS,M�:g���K��6�>pP?S�f>	 t>��3�A8���P�&(��=�}>~&6?�����9��u�ѻH�>�ܾN�L> �>�>4�)L�oږ���~���h���w=�3:?�?����@���v�0S���)R>BJ\>��=��=L�L>��h�jCɽ{�G���3=3��=��]>��?�->��=��>�ĕ�/�_���>@!7>EF>b;?�(??��g�)��Q��������>��> ��>d��=U�>�n�=E��>%Nu>M���ߞ����q+>��=>@5s�xaa��m�M
�=~zD�5�=�=�O�Ǝ?�!s�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>bx��Z�������u�ȷ#=���>{8H?�V��/�O�P>��v
?�?}_�̩����ȿ\|v����>#�?i��?�m�(A���@����>���?�gY?Jni>�g۾�_Z����>2�@?�R?z�>�9�#�'�=�?�޶?�?x�]>�?�?��{?ڿ�=��h�?�v}��qC��7!�V��)�>��оS!����>����&�N��r����<��<��>\4>��$@ֽ�@c���U�y�*�52>2w�=�'�>7��>��>m��>�>B�=��S�l\.�\Q����K?~��?���2n�A�<���=��^�&?�H4?��[���Ͼ�Ө>y�\?>?�[?(d�>9��L>���翿�~�����<��K>�2�>�J�>����GK>��Ծ�0D�hm�>�ї>����>ھ&+��{jB�>2f!?���>Oή=ٙ ?��#?{�j>�(�>IaE��9��J�E����>Ǣ�>�H?�~?��?�Թ��Z3�����桿��[�K;N>��x?
V?uʕ>`����MhE�aAI����a��?�tg?�S�6?62�?�??h�A?�)f>Ç�ؾu�����>�??����}D��X4���.�R�(?�I,?���>:��L�g�~p!>�2'���ӾQN?�NQ?��?�-��=\�	��*,;<)F���'�<��<(���}&><��=��=�-�=��<�� >nq�w�P�	|;�e�=_Jq>Hu>T��u�8��<,?��G��ۃ�]�=��r�vD�r�>�FL>���)�^? o=�w�{�x���x��hU� �?��?j�?����h��'=?�??� �>�N��E�޾%��Kw���x�yy���>9��>~�l�����f���sF����Ž>p�Bg?>��>i��>��>í�>�U��*Q%����-�ܾ�^����I*�	!�gY�g�����Y�4j���1; �{���>}�ὟA�>��?~mu>ZL�>�,�>!׽K�>��&>.sx>��>�)>�k3>��;>��1=\j�=3R?Z����'����ð�4OB?��d?A�>��i�h������,W?z�?�h�?�cv>�^h��/+�=??�>�3���T
?X�9=f�����<���������U��/+�>W�ս�:�s�L��e�*u
?A!?T̉��H̾��׽�������=���?�<$?�'��rN�G�p�w4V��N�yaz�㧀��毾HV$���q�c鑿`������t�*�hI�<��&?R0�?(��7"�������j��i>��1K>�#�>??�>�|�>1/>f��-�e�\��L,��N���{�>Ebw?��>8�:?��7?�V�?:H<?�f�=W�>.ɾ�,?�* �]$�>r��>�l?�Y:?%�@?{�?��A?��>�_��,�ž������8?��>)`�>�Z
?U�>?"T��ؐ���l��|m�C�����:5��>vj�=�4���]��X�wvB>�H?t]�g�8�����Y�j>��7?��>y��>����[����<���>��
?�U�>����llr��c�x*�>И�?����=��)>*�=ꅼ]0Ǻ�D�=W6��㼐=�愼%�:�x]<�#�=�є=/�i�������:sЎ;\�<�t�>4�?���>D�>�@��8� �C���e�=DY>S>�>�Eپ�}���$��S�g��^y>�w�?�z�?'�f=��=n��=�|��"U�����p������<�?J#?XT?V��?|�=?dj#?�>�*�jM���^�������?A�8?Ѐ>B��g��^x��M�+�2?C_�>Z�j�����X���iI��y��+[4����꒳��+2�d�h=9��F7����?���?��A��|2�+���Ù��ľ_�4?��>Z�\>[A�>H�(�"�g�+����=�V�>��d?#��>D|J?�q�?l�m?:�Y>o)������	����
��a/=��9?�{?���?E��?9q?��=�#���/��,������O���%p�ׅ�qI�>��>Ԡ�>�;�>�q�=,��:4�[JG��a/=< �>i]�> m�>�@�>l'}>�ҽ=,�F?�@�>�ｾ62��ɢ����i�*���r?*�?ѝ)?�-=~"�`EB��/��=G�>�]�?[��?N;*?�yS�\�=����.~����a�nڷ>X��>��>֟�=5dA=b>���>��><���}��8��>�e�?��G?�>�=cմ��_��ܨ��~1�s��>��e��vq��C�>�H�c+�>6���E��>�֩��k0��hݾ�80�ڴp�kq缓�<@$?^W�=�/�=���=�=��e����<>�ߎ�Fɍ>�.ƼseW�-"����K-2<I2���%���"� G���˾�}?7I?`�+?#�C?��y>�O>H�3�&��>ץ��8D?JV>b�P�<����;�䪨�="����ؾ�u׾Y�c�2ϟ�vL>OI���>�93>�C�=��<��=��r=j̎=WeR�1=��=�Y�=�`�=f��=N�>�E>�6w?X�������4Q��Z罤�:?�8�>h{�=��ƾq@?~�>>�2������yb��-?���?�T�?>�?@ti��d�>L���㎽�q�=M����=2>o��=x�2�S��>��J>���K��D����4�?��@��??�ዿТϿ4a/>�L7>T^>��R��1�.�\��`�m�W�'�!?�);���̾/�>�>�=��޾ƾ��0=҃6>��_=j�h\����=I ���>==kn=���>�C>�M�=	����d�=��E=X��=�.O>쵥�Xp9�9*+�Y�2=
�=3?c>��$>�T�>��?�,3?�Te?P�>:h�[.ʾ�2�_]?P�e��m�>��=.��>�H�>�E?kj?+�a?���>dt�Ym�>��>�W��Y���v��!p���s>�Y?�_�?o"�>���<x�=���,Q����B??�S?�)L?+�?@B�Z׿�v������{<�=x��
��<��f=w�=�?f�
.�=�t���I�>�h�>�>�D�>;*�=��>�'�>>��=%O�=�@/>-��>*a�=$ɸ=�AO>ʚ����=I�ͽ�W>`(=�6�<�ޣ���=�}�55=}_|���=C:�>yh>���>��=l��:s0>斾��L�s)�=�צ�&BB��c���}�r�.�*h6�JWA>��U>!9��#����?�cY>р=>݂�?cHu?8 >u�
�V�Ծ�m��m>c�xT��6�=t^
>B�;�S;�u�_���M���Ҿe��>bR�>�1O>�q�=�t��| ���>o��[NU�T��>~�|�#�콜��Bv�}ʝ��U��N^����R�H�W?�c��MkX>�*J?�1?��?*�&?8�=O�)�3��>�z��o�8>���/��l�>�l3?o
1?K%?���t�>��G̾�����ٷ>�#I���O�����
�0�����Ʒ�<��>����һо�&3�`d��<�����B�wRr���>��O?�?�b�5V���RO�B��M���&Y? mg?2�>�D?-6?�������,���n*�=�n?���?�1�? �
>�$�=P{��BT�>D>	?7��?f��?sPs?yA��e�>�G\;��#>����[�=!(>J�=n��=k1?�_?�i?���{	�[�����<]��	=�=���>7I�>|�r>
��=�<^=�=�([>���>?��>xtd>ԡ�>no�>�a���� ���?d�<-L�=�b?��>/@>�9���myN>_�������>I����=�~=����3{*��K� �>�̿�Ȉ?���>�%۾���>0���c�׭�=❾>�Dp��2�>Y}4>&��<@_�>���>@�>un�>�?;1Nɾ��>����#�B���P�VԾb3t>M��t��P��7ｧzQ��v��5Y�j�����L�;�vu�<��?� �jle�ؙ)�V`��J	?s��>]�0?�����i���>�'�>ؐ>����%��v����'�F��?�4�?oBc>���>�W?)�?a�1�4�2�3iZ�U�u�#A�9�d�'�`�፿m���2�
�K����_?o�x?:kA?I��<e5z>&��?��%��ʏ�D4�>�*/��3;�i�:=�7�>�)���Ha�k�Ӿ��þ�e�f�E>�~o?#�?�O?S<V�=0j�ҧ'>��:?��1?�`t?�W2?��;?0��{K%?;�3>*G?)?��5?-f/?l�
?�z2>���=�8�`�'=%N���튾ܦѽ>;˽�J��Y�1=7�=�#:��<�R=���<n�n�ͼJ6>;�ߨ�n��<%
7=h��=��=г�>��S?���>ak�>Q�+?��e�R(�p��K�L?V�L<����@��ʽ�C�6?7>:t�?�+�?Vl?�vq>�Y�j�� >��>��=y�=��>�v��+�����=� &>�a>>%#>UM:Z��g�O���S�=3��=7~�>*"V>g}���G->|q��uWL��fr>�<�_:����O��@>��J4�R:f�0�>��I?&�"?п�=�o�:[ҽ$�]�'J'?��3?��K?7�?iT�<w�'�@���@�/3��o}>���p�=٢�gs���8��.#=_�q>���hd��a�a>�7�����Tm�~sK��\�Y=���$Q=h(��Ծ�������=RQ>�j��d�!�I����7����H?��\=ǫ���lS�&�¾��>7�>B�>S�l�ɢ��p�<��5���=��>F.>В���Y�><E����V�>�QG?��`?^��?�����ep��%D�2��@Ǟ��K�F?��>K�?�5T>�ɭ=NӸ��&��d�{�E�j��>���>z��� E�a���]��ƭ#��F�>��?ƕ!>�U?ϏW?� ?&�]?U�'?<+?��>���O����E&?x�?<7�=<�нT�T��9�I�E����>��)?F�B�aX�>a%?z�?�'?��Q?n!?� >B����h?��O�>`�>m�W�����j�a>��J?^��>9dY?���?<I;>|5��=���8�����=(�>J�2?��"?�?��>�
?{���?>�>�2?�?��?��>L�5?��T���?~��a�>���>��s>Vv`?��z?^??�'?�o㼤��iK,���{�B�5���=bh-=�0��_`�G�1<��B;+�#<�L�=?(=r-X��W��=Z��8�Y���V�>�K>F���� >⳦���-5->2Bv<�x��.R�r�_�&�=ͬ4>�$�>�c�>Z*8�/�G=ϊ�>]j�>����-?�?�?����j�Z�������p�8�>>LI?e��=�Qo����P�v��U=F�p?�:a?�LM��
���b?>�]?�h�=�w�þ�b����i�O?h�
?n�G��>3�~?��q?f��>>�e�B9n����IDb� �j� ʶ=�r�>�X���d�&A�>I�7?oN�>��b>m+�=v۾��w�vp��?��?R�?���?0*>��n��3�!�Ӿ�Џ��z=?���>K֧�B�1?���<�䢾Zc�������鮾��������H����r��K����m��+}�ᚦ=5v	?�:�?�r?�kf?�i��y�^�j�P�u{��{G��� �
�Ȳ;�{�H��AJ��i��kb*�30������+�>��%�A�n��?�'?r�+�Ҡ�>D������̾��G>ؠ��/��<�=˾��?�G=^R=��h�,��ޭ��l ?zY�>�s�>p�;?�[���=���2�a 8�a�����6>�b�>c��>b��>�̺L'-�W�{Ǿ����Lb޽L~v>dd? L?Pen?�����a0�h�����"��~$��ᨾy'C>l�>��>�MO��8��'���>��r����>ӏ���	�F5x=�2?���>�˜>�ؗ?��?�N	��{����t��(/��ڏ<
¸>��h?�>���>��Ƚ{^ �h��>(�l?G��>�>閌�*Z!���{��ʽ�%�>.ݭ>���>��o>
�,�x#\�k������9��p�=]�h?Ⴤ�B�`�J�>�R?���:b�G< {�>,�v���!�:���'���>�|?p��=A�;>f�žF%��{�98��*y(?/1?a���٠)��e>ys$?���>7�>nĄ?},�>����6��a?�1Z?��B?n>?/^�>��A=�h��]���v�+���*=ϥ�>`>ZЀ=z��=��Y�D����(r.=w��=��H� 뾽2�*<�G���h��2=�^5>�_ٿgKL���پh�Ht���	�׉��;���9���/��ܻ�ߺ��<�������O^�*Fi����C�i��{�?0M�?񳎾%n���;��R�}��+����>�dj�w{/�d������Z
���
��:�����.J��e�u�i�h�'?O쑾-�ǿ�/Oܾ*9 ?O5 ?��y?��è"�Xr8�{� >��<�����m뾋�����οO�����^?���><��󣽇H�>9��>.�X>Tq>��鞾p�<~�?z-?c6�>Tms���ɿo����$�<���?��@SA?})�%M�T=�)�>~�	?��?>��.�&x�3���9�>s��?�?�I==\W�����d?�� <��F�Dý�ٌ�=PO�=+�#=|����K>u��>u��$B��T޽zr4>@��>��/�Ǔ��Eb�.��<h%]>�oϽ�[��5Մ?,{\��f���/��T��U>��T?�*�>U:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=n6�ĉ��{���&V�~��=[��>b�>,������O��I��T��=
`���ǿ�.�Z�0����=yD�=�8:�d>50�%�J>P�־Բ ����Y=�;�(k>n����y><��=@��>8:Z?��c?q��>좛>�y�=�������z3��0���-�9.��W���\���IB�*g;�G�d�w��I'��3����Ӽ8LO���������xi���|��?J >+?>l�w��ED���H��ھ,��=��<.��+�#���n�,K�?��R?�܌�	i���������֮�fn�>S�������ܾV����>߬1��`Z>!M?>��
���v��I[�"60?�?����lY���%>���m5=T=+?��?�<<�@�> 3$?�'�Z�ཊ�W>YV4>䒤>Hr�>	�># ��M6޽~?��S?�$��[v�����>\4��m�t�3d=�/>�66���
���X>���<Iɋ�����>��fl�<2&W?���>9�)�� �5e����-�==H�x?�?�>	zk?��B?�Ƥ<�`���S����w=�W?'i?�>ň��Qо�o����5?�e?s�N>YFh��龟�.��U��!?��n?TU?����ro}��������i6?��v? s^�ts�����8�V�t=�>�[�>���>��9��k�>�>?�#��G������uY4�Þ?��@���?��;<��w��=�;?c\�>�O��>ƾ{��������q=�"�>����ev����(R,�`�8?ܠ�?���>�������S>��(�̲�?�{?�榾���=F	�+@c����)�X��G>�W!�������-�b�����������~���F>��@P�>'�>������߿4�ǿ�蕿��U�J����>�+�=��E<{<\��k��'����X��jj������0�>�=>Hwҽ`�ǀ�VI9��=���>�*����m>d��J������텣��4z>���>��j>��	��JԾ/��?�Ά=̿k晿}f�^�f?4�?=*�?�J'?q����,�oPO�$~ﻓ�J?�p?�V?iF=�/R�u (�"�j?�_��vU`��4�oHE��U>�"3?�B�>I�-�F�|=�>{��>g>�#/�v�Ŀ�ٶ�0���[��?��?�o���>m��?qs+?�i�8���[����*��+��<A?�2>���I�!�A0=�QҒ���
?T~0?{�_.�T�_?�a�c�p���-�H�ƽ�ڡ>2�0��e\��L��4���Xe����Ay����?3^�?W�?k��#�-6%?R�>$���n9Ǿ �<���>l(�>*N>�G_��u>	���:��h	>���?�~�?<j?�������&U>��}?	�>�?~�=lC�>7��=g氾F[*��^#>b��=�x?�9�??�M?dB�>�n�=��8�W/�tPF�)KR�V-�9�C��>G�a?DvL?�Qb>/⸽�2��� �^+ͽ�d1���RZ@��G,��<߽�\5>��=>O>0�D���Ҿ��?p� �ؿ�i��:o'��54?���>��?P��V�t�۳�;;_?ay�>�6��+���%���A�s��?cG�?.�?ʺ׾9V̼�>��>XI�>��Խ0���w���n�7>ʞB?2!��D��=�o���>���?�@�ծ?i�L	?� ��O��:`~���7����=E�7?�/���z>���>��=�rv�Ẫ�n�s�r��>�@�?�z�?F��>��l?9|o�:�B��1=�F�>Ùk?�l?��r�?�+�B>8�?A�������M�f? �
@�t@n�^?\ׂؿ�)��lվ5����<���=��>f\=Z�{>��>����P�=1�>���>=<>��h>o3�>�>@�&>����y4�h��R����0�_���C&���l���h?�z_5�:^i�y%}��ỽ|��;��]B�����v �;�A�=��V?g8R?�Ao?���>؏v��>�'��=�['����=��>3?�IN?&�)?;K�=솠��?d�Zs��,T��xK��o!�>DM>K��>��>���>.I�8��D>=�C>�C�>�I>T-)=�
��=�oQ>b�>��>�ĺ>�۪>�>�Rʿ;)����(�%�K�����?+3ܾ��R���G<���޾���:,Y?��<dT���GĿ�T����C?�e�S�8Rܽ��B���?�Uz?(1>2�,�J箾�V�>��S�v�彞�>cr������f�cP�>�|v>Xge>���>��6���:��VR�e4���>��2?�o��C�@�'�j��E��"ھ8�R>��>TtY��$�8_��΀���k�HO0=/=9?���>v�ٽtҭ��,z�����e�I>9R>;=LϢ=�U>�I���N�E�I�[=���=�U>nQ?1+8>$�=km�>x����jU�7ì>��F>|bA>_�7?�9'?�k+�HIϽ)Ih�W��ދ>�>&'�>!#>�WD��_�=P��>kj>��
�f�n��D� ��mx>����~o���?��8�=hL��� >t��=�j���K����<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾQh�>~x��Z�������u�p�#=N��>�8H?�V����O�g>��v
?�?�^�ީ����ȿ5|v����>U�?���?h�m��A���@����>:��?�gY?soi>�g۾@`Z����>ѻ@?�R?�>�9�~�'���?�޶?կ�?7U>���?Vă?wX�>kN��X��i��O6��� [>g�����N>�s����=�-A����8���r!��#Q6� ��=�m�<�_�>ɷ=�ש�E>G>z������օ�ɽ�>=L�>�
>��>�?D�7?��?R�N=#U1��v����`��K?翏?:"��7n����<7�=�t\���?��3?-�s���;���>UQ\?ꕀ?�Z?{�>��)A��鿿�.��ϐ�<��J>�c�>~��>�~����I>�Ӿ�(B�-�>� �>�'����پ�ـ�����>�!?C��>�D�=ٙ ?��#?r�j>�(�>OaE��9��E�E����>���>�H?�~?��?�Թ��Z3�����桿��[�;;N>��x?V?�ʕ>b���냝��fE��@I�����_��?�tg?�S�H?=2�?�??b�A?�)f>����ؾt�����>A!?�8�A�B�&��E�M<?�?hP�>C����qٽ�Ѭ�c��pQ��8?��[?�%?U����`���þ���<�[�|���X�;	�N���>�>�����j�=��>6�=nm��p4��Zp<��=���>O�=��4�oڋ�p<,?�H��ۃ�R�=��r��sD�N�>�HL>\����^?�b=���{����z��U���?���?fj�?���o�h��)=?��?�	?y#�>�P��^޾���7Nw���x��v���>;��>ڟl��徧������� F����Ž�����?5��>��>��>%YN>���>홗�wG%����څپ��S�V���/��](��.��m���Q�۽�oRӾ�Cr���>Dd��]�>�z?�G>E3�>�+�> Q���K�>�eC>,��>6ּ>&Ȋ>a�">��M>�	�< ȶ��KR?����۾'��������\3B?�qd?1�>�
i�������1�?J��?�r�?C;v>c~h��++�an?o>�>����p
?;U:=:0�e:�<^U������/���
��>E׽� :��M�`nf�Pj
?V/?���̊̾�;׽����
o=�M�?`�(?��)���Q�̽o���W��S�C��35h�,l��M�$�o�p�H폿 _��
%��J�(�Gl*=��*?�?w����k ���&k�T?��[f>��>w"�>sݾ>2mI>�	��1�^�FM'�x���1M�>�X{?V9�>d<?��??Fs�?�o?���>���>w���?l���>��>!�\?p�-?#?�v?rC?���>dG�=u˾�=�6�"?͹?=��>�;?�s!?��b�~-�@��=�|:��f�0�̼�N���Q���{:;�=��.>ֶ>�?��ʽ�t2�>���x�>zE?��?�W�>�~�L�����%>飪>)��>fc>��
�Q�^�×þ��?y?�eA;�/6=b��=�=>��?<Xյ���=2��=B�
>�U�<VQg��K��δ��Ϻ<��=�Ϻ5n|���B=�/=u�>.�?���>�C�>�@��� �B���e�=�Y>#S>�>Fپ�}���$��n�g� ^y>�w�?�z�?e�f=��=��=}���U�����C������<�?,J#?XT?[��?s�=?[j#?��>+�iM���^�������?RE?7T�>|�7��H��,����o�zv�>��>ɛ�]�V�(�V��T$V��s7���t�\��?��&�Q�8��C��2�=0��?���?�`
�������i����4g���?�=�>c\�=��?����]����0�>�>v-4?���>M�o?/,�?V�P?@ws>�����T����|�=����c�,?�jW?"l�?�B�?�>�;@��]�����C���'W�3����]>��>:�>6� ?z��> q�=�뇽zQ���!c>Ӷ�>��<�4�>A�	?�?ڨ�>�w»�:G?��>�r�	�Zv���d|�>4%���t?���?=�&?Fq2=>�b�E�c���%��>^w�?�
�?;*?��I��M�=���!g���b�m��>�O�>+�>2Q�=A_=Yj>'�>F�>#�}����8���E�D�?1D?���=?������.U�]6���?׆������ ��>H���� ?�.�-G?l���w��+�;�惾͆x�����o*��,?�|=�.W���>p(>�*��E>~l�=�@="�>mNνTc=�o���>�oN��tN��4�jPg>LKO�t{˾ʍ}?� I?�w+?͟C?��y>�x>�i3�☖>a悽�R?a�U>�VP�7g��vv;�ڛ����-�ؾ�׾Od�䟾vR>�bI�y�>� 3>W��=![�<�>�=fXs=��=��X�\@=5:�=4��=W3�=���=[>�d>�6w?F��������4Q��Y�b�:?D8�>�{�=Z�ƾ�@?��>>�2��ȗ��|b��-?x��?�T�?�?�ti��d�>����厽�p�=-���/=2>m��=��2�m��>��J>����J�����i4�?��@��??�ዿߢϿ�`/>B�>�sN>�JU��j8�[���p&�9�轃�?��/�yy���>hY=Wþy�����=�%3>P5�=�;h�l#e�(�<7 "����=�L=	�}>w�4>����ʩ;i��=�,=���=�0>`=p�u��A.=��m�g7>z�>J�S>.;�>|�?BX?���?��T>sᎾ��W��(ᾫ>Q">#��>�w�ؼc=�>�_?V�Y?��\?p�
?��>��>q��>�w8�%"U��K���������_ܒ?*-o?ܷA>�:�=��7��W�p�����"=��,?�F�>��>ߞ�>����࿟!��hE�6O׽H��<�?�����!�߼|�=8�a�:��=&>v_�>΍�>�Á>$�>�	>��r>G��>ff�=w7�=5s:=+�<fX�=����f��=�[����=�Z����\<���ń�鯥=�	�C$��i�[�I�=�p�=t��>n�>���>��=򋴾-F4>����L�$$�=.ݣ��A�Hc���}�;/�63�(�>>�*Q>�h���Q�� ?.S>�=>6��?L�v?� >��|�Ѿ�4��Y>V�72N�nq�=�L>�X2�:���\�W�L��VѾ���>�ǲ>�d�>$�=`P`�3
V�pZ>���,kL��,�>0Ih����&���i��ѭ�f쌿��w��T ��^�>�,����u>��F?�t+?�"�?�?Y�A=����>,��	��>B����:��ǒ<[<?��0?V�?\�׾�Y9̾����㪷>jZI���O�+�����0�D'��շ����>�"��2�о�=3��]���쏿�B���r����>�O?�?2�a��E���ZO����I ���I?6Qg?��>�W?V@?J�����\���T�=��n?��?0�?�;
>b�>���	�>g	?�4�?yI�?�8x?��D�s��>9����4>6�ɽp�>1>>n�=.�Z>��?.�?t�?.,������L;�}��VJ�T@�=�,�=�)l>��A>Uc�>VW�=��;��:=(�2>��>"�`>(׃>���>�O�>���������>Ld/�C���/?�yZ>��=���7����%>Z�D�dTO��"T��
=��J=|�<�%n�EFU����>I�տ�ʆ?���>}w���	6?M�JQ>���=!��=I'��9~�>A�=*/��W��>Dş>��@=q��>@��>q Ӿ7>����`!�*C�'YR���Ѿ��z>
���`&�h�������'I����}4���i�l$���5=�_ɸ<�A�?,����k���)�����L�?t�>r6?:�����A9>���>�z�>-���>��������iᾗ�?���?�6c>4�>G�W?*�?�a1�3�;qZ���u�#A���d�I�`�؍�o����
�	���^�_?��x?yA?M�<i^z>.��?z�%�������>�"/�=7;�\�;=(�>����`���Ӿ�þBV��CF>S�o?�#�?D?��V���R��O*>�99?F�/?q�o?�2?�x=?����&?�*(>ve?��	?p�5?s�-?x�?�2>��=��r9��D=B��"c��prǽ
ν��μ"�B=���=��p::�(<t�.=5ם<pM
�O5�w����N����<��)=>��=�g�=4V�>T�Y?���>���>�64?)�D�+�"�����3?8��<��h��"��Y���޾1�&>�@t?��?X�\?�8�>d}=��H�{�>A��>�;>O(�>�r�>\�ӽ��#���E=��=V�>9��=]�u��q����M!��$?<z>u��>s�Y>X��%>l��}�P��b>�7��2��#�f��@��}/�,�t�6�>�J?h�?%��=A��v稽�G^�2�#?6t9?ݜS?A�?�e�=�ӾAN8�6H�ы ����>b��<*����V��[l;���F���>�ą�	j��V�_>P����޾��l�z�H�m����S=5L��b=����Ӿ��}�aW�=,5>i뿾�� �q�������J?�qx=3奾�UW��.��F}>�>�a�>�
F�ۂp�.@����=D�=���>�F:>%��:���G��D�1��>��M?~?�Ѝ?=�������j*�Ʒ$������p"<H�>?
A�>#�!?H�>t[R>[N�n�þ��Z��k����>�K�>}I�H3]���u�SI���6�y$>ə>�>���>�li?��>�V?<)??��>f�:>,���1��?؆?)�$>ID��w�T�d��6a��z�>��M?Ԝ߼9��>W�?�=?7�!?m$l?O	H?i��>�0�2�>�!'�>�g>��R�QQ�����>��T?�@H>��s?~�?��>'�K�x�ʾNy=�����=�*?�1?�{�>��>(��>�h���e;\�>��>B	S?�J�?��R>lR5?#w	>Er(?�2>�_>?V�?gnO?M�q?rc<?�h�>ťV=��⼀��c�ý<WIU<���3�?>ad�=�/B�[)=�>"����\��O>��= , ���V=y�=yU�>+t>�ϕ��u1>B�ľ�~���A>N����?���&���:���=MV�>��?;��>�(#����=���>�+�>���K4(?��?/?�,.;ȩb���ھ�K�� �>i�A?)��=��l��x��n�u�v3h=��m?�^?�W�H��L�b? �]?3h��=�
�þ��b����_�O?;�
?Q�G���>��~?Y�q?E��>�e�.:n�(��	Db���j�Ѷ=Tr�>KX�C�d�t?�>h�7?�N�>1�b>>%�=cu۾�w��q��k?�?�?���?+*>��n�Y4�[����/V?F��>�痾��>*�9�����˾�� ��������=�Ͼ]B���}žRۀ����Ϩ==Fq>�}?�'�?�^~?B�^?����ᯍ�14Q�9�����g�N�C��DM��7k��ND��T4���t�K�վCݾ����$�=찀�G�@���?��'?cv+�%��>sw���;�_�˾��C>AើPv�6h�=�f����H=�]=�d��A0�0���K> ?�Ⱥ>\�>Ի;?��Y��Y=���1��7�4����;3>
��>�=�>�M�>�ᵺ�],����pʾR�/Խ<̇>$+q?��2?+v?�h����A�݉[���!��?=�5��n?>q��<1w$>EA��<����
�:$�q"�����|������ӹ=��e?k�B>>F^�?1��>����y����=$2	��s>��>1��?UaH?�F�>{U�='�:�C��>-0m?��>�	�>?B���J!��{�9�ֽ2��>�ߦ>M�>�c>;Q4�d�[�Rŏ��q��U�8��[�=i? ჾM�^�][�>ZFP?Ar�^�<u�>��w�c����(�%�|M	>��?��=|;>g�ž�&�7�{��v��N2(?��?u���o0%�B��>�I?��>%�>�ȇ?&��>B5��՗<��?�
]?�"K?�rE?�<�>U =G����<ν��)�_J=Ӟ�>_g>?��=�2>����3Z�@99�w�<q�=ّ@;Ő��c��������<�=##>�ֿ-(H��&׾W��T<Ͼ����!������.O��/���!�¾��Ǩo�\���ض���C�oSm��ę�����˼�?���?���2��I�����{��T�f8�>ɪ��1�T�|�����<���w �(F��ĥ��U���f�J.b�EOM?d3��A�ݿ�Z��e�վ�1?�r?�PV?��=��ɾ�,��!�<t>���<�����5���=ܿn?ν�F?mI�>.����=�D?r���ʰ>���>�������]>��>k��>�O8?����迪Lȿѩ�>��?ߚ@�{A?��(����V='��>'�	?8�?>�G1�TH�n����W�>;�?���?��M=��W���	�9~e?1�<��F�a(ݻ
�=E�=_=��݀J>�S�>́��aA��hܽ��4>Hօ>��"�t����^�d��<��]>&�ս�;��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�����/�� ��*��;~>�0>�A�}9i>�- �o� >3����=	H>�h>��~>ucA=�*�>{x�=2�=��Z?�R|?5��>I�a>��I>�������P�{�A�7�����о�1��\^�(s���-Ͼ*�(���1��*��<�X6X=�eY�ˇ���Ԫ�l-�zW�R*?�
)<����a����=B���� �۽�=���;W? �JE���{���?6�J?̓��vr��0!�;:���1��??|��7��E��Mܑ��w�Y���<�>�(�=��6�1	!���P�>F0?�,?�<�� m��u�*>�����=��+?�2?��S</R�>=�%?�r)��>޽N�^>�!:>�ͥ>�=�>
�>����Dܽ��?��S?>R��N���ɑ>����_z���N=F�>{Y.�c�ݼ�\>'��<U;���G��L�����<s#W?֘�>��)�Y��Y����t�<=��x?4�?�%�>%zk?[�B?���<�_����S���1�w=2�W?�"i?��>]Ł�^�ϾEx����5?��e?.�N>�Gh����U�.��]��$?��n?]?u���o}�Z��/���b6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������Z8�=;链��?�φ?�V����;�j�PNk��� ����;��=Ʒ.�+6=�x�w8��ǾZ
��<���Ġ����>�]@؏ս�>�%5��S�5Ͽ����IоPWu���?�N�>.�׽A����Kk��Es�2�F�7�G��1���M�>}�>��������v�{��q;�#2����>�+
�>?�S��%�������t5<��> ��>���>.��n轾+ř?�b���?ο5���ԝ�ɻX?h�?�n�?�p?�9<�v�I�{�_��{-G?w�s?Z?Iz%��<]���7�W�?c�žc�^�n(E��t�5"_> �C?~�7>��O� u>>��<nq>NC>`!V�eɿ�����y��f�?��?<Q��s?�ϯ?�D'?�GF�^㙿�����Y�]��<�n*?��>�b���u��QQ��Qf�3�?&9?�������G�_?��a�	�p�i�-���ƽCۡ>�0�8e\�c<�����JXe����h?y����?8^�?m�?���� #�46%?��>U���
9Ǿ��<I��>U)�>�*N>4H_�D�u>��'�:�i	>���?�~�?j?𕏿�����U>��}?�#�>��?Uu�=Re�>h[�=����2�,��g#>a(�=�>��?��M?yK�>�U�=�8�H/��YF��GR�9%��C�3�>4�a?��L?�Lb>���x2�%!�hsͽ�Y1���&V@���,�Ս߽�*5>>�=>;>6�D��Ӿ
�?Rp�:�ؿ�i���p'��54?B��>��?4���t�����;_?Oz�>�6�,���%��9C�j��?�G�?.�?��׾`K̼�>��>�I�>I�Խ����Q�����7>�B?}��D��{�o�,�>���?�@�ծ?4i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?Qo���h�B>��?"������L��f?�
@u@a�^?*��ٿȠ������'~ᾩq=K�K>7�F>�>�=l�l=���<�̼��.�I>��>��>_��>�Rh>]��=��n>�U��7#�e}���󙿹-6�L�����ɽ���������*�����f.�+�}�dᲽU��QwN�	�=(��=N�U?zx\?���?[��>n����T>+j����=� ����>��5>1)?��??P�'?��U>�3C�bjT��1��I7���w��'=?�"J>M��>�>8�>�Q�Io>43�>��>dh>d�>f�$>�v=��5>�w�>>��>�+G>- �>x�0>�ÿz���`e5�����
G��-�?Àھ�F/������Nc�ć���T���8?�F$>�Τ�(�ſ�K���`S?0՚��Z*�4F�2s��ֹ"?��h?a�=��˾�8�ݿ>p�Y��zþ� >TC��Ӻ��i�I��|�>�?��f>�u>Û3�oe8�a�P��|���i|>�36?Y鶾?D9���u���H��cݾ'HM>�ľ>�D��k�~�����	vi���{=Nx:?�??7���ⰾN�u��C���PR>�:\>�U=oi�=�XM>`bc�F�ƽ H�Mg.=���=��^>� ?w(>#��=g��>>难
�J��ū>w�F>�.>�=?&?��i���lƀ��,+�v>K��>���>q�>&kF�;'�=��>�`> ��������J��`=�|�O>+����$a��l���o=)j��s��=��=Z�����:�2L$=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�k�>:}�8[�������u���#=\��>f7H?BZ����O�	>��t
??;_�=���?�ȿV}v�7��>V�?���?��m�?���@��z�>���? hY?�ei>g۾n^Z����>��@?R?_�>�;�*�'���?�߶?b��?ľ�>7 �?�{?�q�>{��oO�tF�����Z�ƽ#[��>������d)�+�4��b�������_d�������>~xq<v�>:�y��ɻ�][�]�Ǻ�[�,?�<���>V��>�J|>A�>aI�>F�w>""�>����B��n���&Ծ}�K?���?���&/n����<���=)�^�	&?�N4?	�[�!�Ͼ�֨>��\?���?�[?�i�>b��"=���濿�}���}�<��K>,9�>�G�>����`K>K�Ծ�<D�qf�>Qɗ>�/��E9ھ,%���G��
>�>�d!?���>?��=� ?=�#?Ҡj>8'�>�^E��7����E�ب�>Q��>pA?��~?�?�ع�1Y3��	���桿�[�j;N>��x?*T?_ɕ>��������E��(I�
뒽
��?�sg?.?�x?\2�?~�??@�A?�#f>���	ؾq̭��>��!?��$�A��G&��
�>~?XU?y��>�㒽��ս�?ռ������� ?:'\?�E&?F��#"a���¾8�<��"��"U����;��C�Ļ>�>l��ؚ�=s�>�=�m��F6���f<�s�=֋�>��=�87��t��+=,?��G��ڃ�n�=q�r�dxD�6�>�HL>j��1�^?�l=�*�{�����x��
U�� �?Ѡ�?Wk�?�
��%�h��$=?�?U	??"�>�J��~޾���qPw�~x��w��>v��>��l���#��������F��7�Ž��ս'�?���>�J
? ��>H�>���>��Ծ5��e���B,���u�q�+�I�@��k��ž��R<�~H>��Ͼ�nW�p�G>ˎ����>N5?d�=�h�>y)�>J��<c��>)I>Dqw>���>w�~>uX�=��=Y3$���m��KR?������'����ڲ��V3B?�qd?a1�>9i������&�?7��?s�?�;v>�~h�p,+��n?|>�>���q
?LW:=C+��?�<W����$2����M��>�G׽� :�]M�nf�Aj
?Z/?7���̾-;׽�Ϟ�!r�=���?U)?1�(��S��ho���W���S�CtC�u�j����J\&�6�p�m������������&��>=.|)?YW�?9m ���
\����j���?�-]>��>�ӕ>��>?>T%
��)1�4)^��X&�Qփ�tz�>j@{?{��>`�U?�2"?SfJ?_�Q?ױ)>u݀>1���N??����>̈́�>,_p?C0?�V5?�1?EE?�� >R�z�F���Ծ��?�\-?l�?#	�>c6?vx���px��n�r���J��:/;z9^>�->��g�GT��|Q>Ć�=X?s���8�m�����j>��7?��>O��>	���,��7�<N
�>��
?�F�>
 ��|r�ab��X�>u��?��Ow=.�)>���=m����Ӻ�G�=����=�)��*e;�։<Rx�=W��=�:s��U��sU�:���;�p�<�k�>��?p�>�d�>1���� ����ڮ=�fX>��Q>�4>��پ������h���x>~X�?�n�?tj=���=���=A���O������[��dc�<m�?�A#?AT?���?��=?�r#?� >�#��N��gd��l8���?�3,?�W�>���ʾ�_3���?`L?�La��n�+8)��¾��Խ�r>�s/��L~��
����C��$f�����ƙ�2��?C��?��C�#�6��3����dS���C?-��>x0�>�d�>��)���g�i)�/�;>��>�R?X-�>hXP?�a}?`�^?}�E>��;��L��r��圏��:#>�C?�?d��?0�x?���>��$>�M���ྊ'�;��5��Xށ�W*=Y> -�>���>�̣>B��=�/��.�����*�q��=��f>|��>3ݟ>�Q�>��n>�B�<��G?F�>)���g�|Y���Ѓ�7=A��~u?���?0}+?��=�:��vE�U������> v�?n�?�)?ݪS�Fw�=�)׼7���q�w��>V�>�v�>��=s)K=>I��>��>������T8���N�Ƴ?S�E?gA�=����[3y������f6�?7���a"���>#���g�>�l��X�>2+�j�!�a�l�4��џٽ�*ʾ0����>���;+���e�=��B=&@�=��?>����P�B=KJv>�?�h]S=��a��V��1׮����=��,����=�Ϡ��˾]�}?~9I?0�+?j�C?y�y>LD>��3���>����HA?V>��P�1�����;�����!����ؾq׾��c�J̟��G>�uI���>�53>�&�=��<�"�=V*s=I֎=\�P�]=U)�=oY�=b�=���=n�>TS>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/> 7>��>�R�{t1���[�\�b�ξZ�p�!?�*;���˾��>:)�=�߾uxƾvP/=S�6>8oc=�q�=\�l��=�{���;=�tk=}>�D>�ߺ=�1����=�I= ��=��O>����^7�_�+��3=`m�=x�b>1�%>��>(s?f�/?�c?W�>���Ilξ�P¾=ȍ>�\�=<Ͷ>n�=�|D>�x�>6�8?�'E?�bL?~L�>��^=g�>7B�>6a-��m�{�ݾ	����<�c�?���?չ>:ӹ;aZJ�G��J;?��P���?<3?]?6��>M�
���1�!���:�u'#=�U>�<>���<�-��d->�n����=��P>b��>���>�g�>l3�>��>h�>R>�>���=97>�K�<��(�K�>5����Ƚ=��C�ĜS=�V*�K�j=v̿=�'�=Tz�<��'�7��= �=7ʵ�ɻ>���>�>Ŵ�> �������>f9��n�L��W�=Ḡ��=I�K�b����78���W��8�=�2{>�eϺ������?�>>P5P>\�?p�}?�H0>�|y��&���)���)���r�w��=�\^>%�ZA,�;.T� �M��t��?m�>*ɀ>��>sQ>�d�v��+�>5�*��BE����>bB����8��_l��Ą��T��g{���9k��LV>UP?�a����>{�a?ĽZ?$
�?��
?�J�<����W��>-wо��>e�������H�=�m?L�)?�A�>5h��.�CH̾L��v޷>@I���O�7��0�i���̷�㏱>����k�о~$3��g�������B�DMr����>O�O?c�?�<b�}W��CUO�n���(���p?A}g?��>�J?�@?i!��Yz�?r��x�=��n?���?=�?)>eݹ=�������>�W?���?���?b#u?c�F�}��>��@e/>zĽ](�=�w>���=�=&�?�5?��?�����H��쾀���J����<�u>=BS�>��>��w>���=ҋ�=��=
q[>�i�>ؤ�>|�p>iq�>�Z�>C&����侦Z?-�=�gD>�EI?'+u>��=XA�+	�;0>u}��������)���߽(�X�^>X>���=���>uϿx~�?f$�=R"�u��>���@	d>��r�n6�=�\�\a?LC�=&\q>���>��d>�Gn>J^2>7 �FӾ%>g��9e!�^,C�!�R���ѾN~z>1���	&�ɟ�Ew���CI�$o��g�Hj�u.��J<=�"��<H�?޽���k���)�������?K\�>O6?�ڌ�H	����>��>]Ǎ>�I�����pȍ�hᾴ�?J��?�sn>xȲ>��b?d?,�O����W���u�>�H��&{���^��p���∿K��q0�UpM?`�e?j�B?nҞ=A�]>�g�?��� Xs�	��>��,�ZD�f��� ��>�e��������sԾ(�����=*�e?��t?�
?�Z�tƳ���=�#+?�B.?!=?:+@?h�^?������(?q!>��!?�)�>-;@?�	r?���>���>.�Z>������k üw|v�P�&�'� ����i��;��=ho@>��9y>t<�0=z=����������"����|=`'*>�`�=��>�<^?&��>��>�s7?�� �p8�0����2?��==��}�H,���m���A���
>��k?���?
W?�p[>t@���B���>��>�,>
�c>ٳ>?S��QQD�X�k=+a>>��=�/�����pZ
�N������<�f>���>�0|>��ֹ'> |���3z���d>�Q��ͺ�O�S���G���1�4�v��X�>��K?��?k��=.]��)���Hf�:1)?w^<?�NM?L�?; �=e�۾��9���J��A��>u�<0�������#����:�7�:��s>s0��:����|H>����!�yU[�%�F�����2�=|=���=��G���􏾨t�=<�>@M��61��˗��;��{�K?eԖ=�t���@U���h��=}>���>(̖���8��A�l��Dn�=2��>�i)>�ߩ�����D�&��qj>1aJ?�s?���?�ԑ�����B%��|'���z�hA=��*?�G?��F?Y��>
�j>�c����쾍�N���X�.f�>W��>K�޾��@����T�2��_��ؓ>���>�ٴ<���>�B�??�?c�G?�o=?]�>�!>�p �T�n?%�?�hO>� /���I�8�b���L�(��>��A?q L�X��>�:1?6A?��L?	3f?��"?�|�>���KN�>��>ډ>��[�V���6�>%�d?d�>��?�?��D>�v$�*��;����G=i��=Z^W?��.?�(�>�?��>�C���[
>eq?�`�>��?���?"'�՛%?�*>�)0?� n= �_>��(?Mi%?kv?? �?�R+?Iz$>���<n%��������*{=	��:������QR���dfa>N����>����$���#��rؽs��=D��$_�>Q�s>�	����0>��ľ�N����@>G���\P��'ڊ��:��׷=ǆ�>�?���>�Y#�6��=u��>�H�>���!6(?Z�??/O";=�b�z�ھòK���>	B?#��=T�l�ꂔ�}�u��h=��m?�^?�W�=%��N�b?��]??h��=��þx�b����e�O?=�
?9�G���>��~?e�q?Q��>�e�+:n�)��Db���j�#Ѷ=[r�>KX�R�d��?�>o�7?�N�>.�b>)%�=fu۾�w��q��h?��?�?���?
+*>��n�Z4��S����~�
�L?6��>x!��g�@?����/��<5��c�t��ܿ�H�ܾR虾1I����ƾ�㗾�m���vb:��d>E��> |�?@&}?/vk?��;�'X���X�卙�5>L�R��f,�}�T�F���`7?�����X�sD�S�¾]:�=P���=S<��ݰ?c?MU��+�>�!���Ͼ�0о']>֭��0Ž�V�=g��U2�=�c=
�e�ow`����8�?�F�>�I�>QD?<?�/�?�$8��J7��ڇT>S�>���>���>������A�9־yn��`y�@�j>�r?�V:?6df?�W�7����I�sI�	'1>y��2 >�q<�}>��W��]���%�*F��Q�d�-��✾��P�=�-K?!sB>&ł>v�?0�>�w��t=��~>iN�r�'>pS7?�q�?ݲP?���>�y
=������>*�l?��>��>����F!�c�{�$b˽�>jG�>�p�>�3o>O-��\��s��텎�i9���=��h?�o����`��Å>��Q?=��:m�D<�g�>��v�Є!�����'��>Z~?�`�=w�;>�cž*���{�]]��є(?~�?7|����(�Њx>&�"?jJ�>4�>UR�?��>��������u.?�k_?zJ?sB?��>��=���#&ƽ��)�,�=���>��[>�Sp='�=~��2Y]���q�==�7�=(ͼ� ��a<�/����T<b=��3>��ڿ�CM��Qپ�9#�ͻ��W���u�D-��A��S�
�Mwþ����.�o��~���C�<��L�聑��k��a�?���?�G�6`�m ��)!w�����d��>�lg��K���۾��������&��>�@&E�6hw���f���M?m>ξ8Ͽ�����+"�Q
?3��>��N?G�����A<�V�1>ҍ4�`�y����H����dȿ�G5���u?(�?{��_�1��/�>q�!>՟>�>����:����S�?�~�>9��>�A������̿4��>.�@߈@�zA?$�(���v�U=���>��	?��?>�A1�FK�����BW�>48�?��?�;M=i�W��
�,{e?�c<��F��޻o��=G�=��=�����J>�W�>�Z�5ZA�Q!ܽ�4>7օ>�"����|^�鄾<7�]>��ս` ��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=ٰ�����!���U��ý�ND;lى�>H����X�ߺ��Aض����i��=�<>Z�T>��|>{O>¥,> �\?ier?�P?!k�=r�������Ҿ�RO>G��e+����������X侁���<3��7��g����>�#𾡑&���;�>:������s����i�Fm�9�7? �=�t"�i�i�Mw>o�ﾣ ����=᩼!qƾ+�J���x��j�?;>?�t���I^��������b��i;?�g=xX徜�׾>=#�	��=������=�'�=�f3�0�#��\%��r0?�T?����c���*>D� ���=��+?�?�\<m,�>�E%?o�*�I,佃V[>m�3>�ף>T��>GP	>M���w۽t�?��T?a��\5ʐ>yh����z��Ca=�>�B5�4e��[>J�<���T�W��j���f�<��U?���>�*��M�zg��GUݼ?<d=BIx?K�?��>Nk?K�@?��<p���fT�O �cHy=��X?fi?�>����̾�I��?K5?�e?�:O>�X��z��+��I���?1�o?i?(���Z{��ߐ�s��a6?�v?s^��s�����|�V�\=�>�[�>���>��9��k�>Ց>?#��G��꺿�pY4��?l�@���?g�;< ����=�;?q\�>��O��>ƾ*y��������q=^"�>����{ev����nQ,�&�8?���?K��>�������2��=�q\����?���?����,O=�����h�?�
�����Sr=���K
����A����p��Љ��=c�v>}L@B�@����>�b��4�Xɿ����Ažž�?�A�>�5,�񎮾�t�Nb�i�:��oI�Wgp��D�>�>gI���ꑾL�{�$N;�F}��� �>�w����>hS�G��6���E-<Ψ�>}�>K��>C\������-��?0���0ο����ai�H�X?ge�?�z�?un?��8<	5v�	A{�p�
��IG?�qs?~Z?Q�"�l ]�\�6��?$ ྫV{�ܠ2�BjD�\=] ?�~�>~#m�֎ =�(��Ӣ=eJ�f�b��*��v˷�|�9��W�?��?x��9=?�n�?�?,:u��j��IIɽ�"�s.q�YM�>��>y־a}����U��kܾ�4?'�>x ��׃�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?^$�>��?o�=�a�>d�=O�	-��k#>�"�=-�>��?��M?L�>:W�=��8��/�D[F��GR�\$�@�C��>��a?�L?wKb>-���2��!��uͽ�c1��P鼦W@�?�,���߽O(5>��=>�>\�D��Ӿ��*?N%��ٿ�����뽽�-?&W>��>�� �[J��#�(�S?��A>�����iΎ�_��YD�?���?�_?��оh��)�!>B=�>��w>�!����̪��{ >^}9?�;�rA����Y���v>��?}r@�p�?I]_��	?���P��Pa~���e7����=��7?�0���z>���>��=�nv�ۻ��Z�s����>�B�?�{�?"��>�l?��o�F�B�7�1=EM�>՜k?�s?�7o���u�B>��?�������K��f?�
@}u@Y�^?��ǿ%���]���PUξ��5>�ט=]�>�p�=��+>���=%�%=$��=�Y>N��>���>B��>I��>��/>�	>�0}����᯿�����F �����ĺY�L��L�U�$����&�����<h0���9.�����&%Խ1ҵ����=�NU?�8R?%iu?���>[N��(=>qJ�PS=���<��=�_r>�5?P�P?DS)?��=�s����_�	ـ��g���ڇ�6�>D�X>�Y�>p��>ִ�>�e<<��->E�X>�H�>�0>���=�n<��U=�_>���>�^�>K��>�G>�>�²��N���mU�R�����)�ݒ�?m����:�(W���0��Q(��9#U={�*?��>dٔ�l�Ͽ"���PP?V�[!���?�QX�=U�1?D�T?�V�=����Wq<���%>�`���Z�;U�=م.���w�(�3��]>� ?�P@>�`>V-��<���I�w����Ah>c�>?%"���+��)z�S�>����B>Υ�>J5Z��P�)6���,}�1�P�咂=|�:?;u?97��!�������F����.>��z>Z֝<6��=�gM>���������H�U�<H��=U�I>�?�� >iԈ=�ό>L���@�嘧>�(�>,�>v�C?^�$?��i�84h�g�~��r4�`\Q>��>o/�>�;*>�32�Y/V=
�?I�>����N�?E�<r���i>��Y� ���hŗ��=w�z�	o>�Q�<��B�~�K��r�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>o����З�����Vr����=`S�>�D?�����������+?���>+�����+����Ol�f}�>�Q�?p�?�d�uC����O�y� ?���?��Z?���>9hѾ�1=�Fۤ>�:?^?-��>����+�J�!?^ �?_��?\�X>��?��f?�>�Ż�@��r�������Y	>��:�]���z����0�5�:��������qT�Bc�l��>Zhd=���>usG�����|�<$L���~b��׈��)?��Q>��>=�!�>��?��Q>��^>Va����L�S���d���K?���?Q��1n�
e�<�=��^��&?wK4?�][�j�Ͼר>�\?{?K[?Wg�>���=���翿�|��Q��<��K>�5�>lI�>���XJK>��Ծ+1D��q�>�Η>���@ھA0���ۣ�TB�>%e!?<��>%ڮ=6Q ?��#?��f>8�>��E�w���-�D��~�>�+�>4?�<~?z�?oj���%4���������!|[�ߏQ>ܜx?��?*�>�W�������T���&�Z����?cg?��轞=?@1�?�@?E�B?,�f>)���Ӿ:��9K�>>�!?.���A��M&���?-Q?���>�:����ս�4ּ���~����?�'\?A&?O�� +a�h�¾]9�<v�"�j�U����;6pD���>/�>Æ�����=Z>�ְ=1Om��D6�kg<Rl�=I�>��=7.7��s��G=,?`�G��ۃ�F�=f�r�)xD�m�>�IL>C����^?�l=�	�{�����x��G	U�� �?��?ik�?!��/�h��$=?�?L	?"�>�J���}޾5��OQw�c~x��w��>��>�l���=���י���F����Ž<���?3h�>G)�>���>,��>�X�>���� *��!�����Y����o9�r�5�
��aB���fӽ2_<V3¾�u���Ɠ>��� ��>?<?Bx>�6�>��>�E�<3��>�eS>"N�>'I�>àS>C�?>��@>#/;ڦ���JR?�����'���(����4B?�qd?5�>M4i�����+��*~?:��?�q�?o4v>]~h��*+��o?A�>}���m
?�{:=��T�<�S�����z0���
���>rM׽ :�TM�Rff��j
?T-?c3��S�̾E8׽JǞ����=�4�?��(?��(�ȒO�;�n���W���S�)&G��i�99��R�&��1p��7��H���%��&� �E=v2)?�ԉ?d ��쾪a��5�l�k=?�k�^>WV�>c�>/�>,kC>�b
��{1�V_� %�]6����>hz?|?z>N?�R?��k?KX(?/�>��>�畾n�;?Ъ>x�>�L�>�A1?i"C?BD>?��A?C�_?����]}���;	Ǿ8?�!?h��>�?�2?�=�eܢ�a#>��=I����}X�L6_�W�=�}&�<N�Ӳ���>�?��"��C;�������p>Y�6?���>�>sT���ul��i�< ��>%�?OE�>1���A]t�)/
�.��>%�?қ �B�=��8>���='pڼ��k7-��=ܐ�b0=8Ъ��-X�K���z��=˧=q�ܭ8�����G<N�i<�t�>N�?���>�B�>�@��M� ����?h�=�Y>�S>�>�Eپ�}���$����g��\y>�w�?�z�?�f=r�=/��=x|���V��+�����&��<��?�I#?CXT?E��?,�=?�j#?��>�*� M��:^�����Ȯ?�.,?�t�>���Y�ʾ�	���3��?�7?R^a����)=)���¾��սr>&s/�'2~�l���C�w�j�����h�����?�̝?��B���6�S�d���r;����C?F�>iD�>t��>�)���g�c�G;>S<�>r�Q?�:�>�dQ?��?i^b?��0>Z(Q�x|���������(>TeA?��?u�?M?vE�>S�>��^�_��'2ɼp3����Fz���d>�T�>f�>�=�>�2.>1����۽��H�Q�l=`-�>;@�>���>��>��m>C�<��G?��>�Z������줾$���<�X�u?�?�+?�q=)��i�E�KB���K�>_o�?���?�2*?j�S����=k�ּ�㶾��q��$�>X۹>"1�>/ɓ=HrF=�b>��>��>�(��`�ip8�\GM��?�F?H��=�E��E:e��b�ʱ�����>��D�Ӿ��f>LھK��>R���>p;p%:��<��L]0�������d�Ѿ��?�m|=��=��]>R�q>�޲���g���x���4>��<��7=8'��D���ّ�h�=0g�=�=FX��˾�}?�;I?�+?��C?Y�y>�;>r�3�c��>�����@?V>��P�Ĉ��G�;����d ��Z�ؾx׾��c�ʟ��H>R`I���>�83>�G�=EK�<A�=s=�=I R�w=$�=hO�={g�=���=��>1U>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>$�3>�/ >��Q�b�0�\S�c]c��U^�$"?r�;�ŔȾ���>�K�=�ྦྷ�žN�;=�7>�Ga=�2�\�(��=�Ew��C8=:Um=6|�>�A>�´=���㪶=��R=�q�=t/M>9���P?�n�)��8=��=S�b>�#>/E�>�?�q0?d?J̹>�o��ϾV���~�>��=K��>�و=�(D>`��>�<8?�D?WL?���>Y=�=S�>a˦>��,�L�m��h侴<��[��<���?��?θ>{F<%?C����y[>��'ƽ1�?�1?�?R��>Դ���㿃�D��J<�"����&�G=˂s�?�4�L����OW��0�>(�>�,�>A��>�#N>?�[>ݓ8>�M�>��;>���=��G��ѽ��=���<g=0B�0)q8�4�?(�<Zqh����W⚽n���ڥ�S_�<鲌=��=
r�>�Q>���>��o=�Ұ�&�5>�ꖾ-GM�\Ȯ=0���t�A��c�H��,0��=�_�6>�b>Fk�:���$?<�O>~�)>�;�?��z?��0>���
ξ�e����K���C�Ԭ�=xu>%}6���6�$X�`6K�:�;{~�>��>1i1>�֎>3�i��D��8�=�c���S����>z���k�I�z���%��P|��ޗ����|�ZC->y??�ň��O�>�wJ?��3?�V�?��%?���= &��c��>c&���f�>{«����}� >$?8(? �?�7ؾ�5��̾���� ��>9I���O�����V�0����۷��|�>�쪾��о*3�sj�����֒B��lr�W!�>p�O?�ܮ?1 b�P��mXO�~�������?m�g?�	�>�6?N?��7��"���{�=��n?;��?W7�?>ov�=㇖�P�>�4	?��?�M�?�*{?�=���>�o)<�XH>½/��=A!">�=)>1�?�D?��?����f�aV������Q�~��e=ݶ�=�^�>hQ�>�o>���=o
�=!�=�h>�Ǚ>�l�>�i>���>gΈ>�͌���
��>. ���M*>��E?���> �|>��b���g=�s=�V�G%H�����]�9�N�(�f=��0>0t�=��>�˿��?�mA>=j¾FS�>ԭ��
�="�Y>���>d%�ZI�>�Ԍ>��><��>��o>T��=$\S>�p>�n��h��=��2/���&'Y�V��R�>ږ��歼b_"��}���Q\�!+Ѿ�j��]�L����CL�e6�xO�?`�3�F]����%��]#�KK?7q�>�j
?�g��h�y�w>'��>�;f>�M�
��ݮ���(���C�?>n�?�c>L��>b�W?m{?2�1���0��Z�3�u�G�A�[�e��=`�<#��������
��"ʽ�]?�Qw?�A?07�<py>��?�$��Ꮎ�u�>X
0��:;���.=�>63����a��ԾR�ľn��+A@>Do?��?�?2�S�6PR�>:n>AQ?;�J?@�X?qK?
�d?��?��1?x�u>/�/?�(�>В*?I�A?-x?���>}W�>w����c���e�Y̢����N����C�+��=j$
>���O�N=/�$=ә�=��6��<;,=�խ���a=KL9=l�>ꡬ=箦>|�]?(��>��>�7?�0�7<8�冷��g/?�;=7��`���������>�k?1��?��Y?�uc>I�A�Y�B�<�>�>Ф&>iv\>Ss�>����E��=��>��>�`�=K�R��ǁ�0�	�q{���A�<��>���>�/|>O	��v�'>[|��-z�7�d>��Q��̺��S���G��1���v�<Y�>=�K?��?Y��=^�Y(���Hf��0)?#^<?�NM?+�?��=M�۾k�9���J��C���>MK�<��������#����:�k�:��s>w1��d���#�_>�����޾%�l�aJ���)rV=�7�Ra=9�MxԾ�������=.�>�2���� ����ส��:J?�]y=�o����X�q�!�>t��>�G�>z�F��y�߫?�d���=J�=ӫ�>g;>������b�G�pr���>1B?�]s?o��?{-��9n��>�'���N̾��=�-?-n.>¨	?�#>H�%>�_������Mo���^��3�>��>��}-Z�͎��i!�@#J��L�>@��>5F>��6?"��?��_>�4S?��2?��>��>��=(S���i0?C[�?.vB>X��^���*O�wRT���?I�*?�ֽi��>��?�E?��E?�e?}6?B��>c��Gw��@:>�΋>��:�s���X�>�nd?��>ls?�P�?ɦ3>g�c�]ʠ�%!O=�!�>�M>�E?V�S?j�,?�`�>�?�>/ᇾ2>#�>��\?G �?6�?mq=+�?)�>�?�6�<OB�>��?�v#?|�_?8��?p�H?���>L�<��ɏ����c{_��bE�z4Լ�t==���ɼ�Z���<�=�a|�������	q��k�]<�U�<Jx�>�iO>/���n>�羾�^�-kV>(U��~e�������+����="�>r> ?i�>��*��g�=��>~��>B<��/$?��
?-(?1X>�xoh�Ĺھ��S��p�>��C?J��=��i�3��m{u�N�M=�j?�\?��[�����L�b?��]?h��=��þ¶b�Љ�O�O?+�
?O�G���>��~?Y�q?7��>��e�%:n���Db�6�j��ж=Rr�>GX�G�d��?�>a�7?�N�>b�b>t%�=Iu۾�w��q��l?��?�?���?+*>|�n�W4�ӊܾf,��o�`?��>�8��Ϩ.?�6�=��ƾ	���<J������ű����ڋ�<���1���5��`b�&�(>�h
?���? ds?�vh?\�O�A�g�Sy���*�D��ѕ��HE��At�vnN��p���Q��K����3=��{�6YC���?e�#?X�(�6%�>*���U뾳�Ծ��I>-0���?��"�='c�w�f={H=�\�2�&�&���@?�_�>�c�>�>?�'Y���A��D0�7�6�-�>>�>���>���>���7�.�ݾܽ�þ�����G޽Z�>v�`?n�A?8?�??Ҡ��� ���Y��R0�|@X��N̾�n�=W��_��>�ϑ���x�@4,�pH+������l����۾n�<>�I??A�;�>�=!�?�*�>W��5WF��憼Mf��eY>��>\@�?{�F?�x=�3��X]Q�7��>�)l?���>W��>�l{�� ���71$���>�ע=Uf�>�w]>9ܽGf��;���������=�Q=�W?6�d��� F>�'a?�����.��!�>��<0�4�b�Ⱦ\!:�5�=�?A�>�j�>ȸ��RӾ_����� )?P?�]����&�R}>��?y.�>���>�6�?���>�2��p|�;��?�b?�}J?plF?\%�>��f=꽾ֽ��&��]=�&�>q	c>��=gB�=�W.��C�����M=�+�=� һ3DԽ�&\:������{<J=�^>��ؿ+eK��dھ��������uV��r����d��+���D���x��I�{��������SI��a���""t��z�?�u�?�����ϔ�������~������>�{���H���d�f����6ھg̨��#!���U���m�~g���8?j����ο�?��?Ǿz�>�<�>1t^?}Y/� ��y-'���.>RA��_]��_����Y�׿2Xƽ��/?@��>W��/�����>�&��"��>(��>�����ϾX�<K�	?���>��?��޾�>׿������=3�?�@�xA?��(���rV=C��>~�	?��?>)F1�iJ���oH�>N:�?���?��M=��W���	��~e?i)<U�F�V�ܻ}%�='h�=%P=���CyJ>�M�>*���TA��%ܽ[�4>Eͅ>X�"������^����<x]>��ս$Z��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=����~�¿�4 �9�7m8>
me����`->�?���Z=4�ƾ>�,��k���>�o>�?�>aP�>hy>�A>H]?rg?��>:�}>�|O=��9��#!x���uܷ�L�ѾR�2������j����a�;��-��w���"�h�H�|郿���� �q�d+L�],?�d�=gP�eFs��=�b�8�sQE=�_E<׾޾��=���t�v�?�LX?��k���u��C1��?5������4?����������p�Op��]�½��;��>+�����B��z]���[�Yu0?�d?�]��`V��d(*>�
��y=��+?��?и]<��>�E%?��*��M�֋[>�4>��>���>��>���Q]۽�|?ֆT?V���՜���>�w��Cqz��Ca=o)>�5��輻k[>�<�쌾+	U��ŏ��x�<qdG?���>�*�$�$F��B�y=�B>�ed?��>j@�>�mx?"�)?���=��#�M��G���<�3_?�u?���=�[߽n�;�^Ⱦ;<>?��e?��J>�	�&��A'6�@E���h?c�r?��&?u4=��x�G"��r  ��u9?��v?s^�ws�������V�E=�>�[�>���>��9��k�>��>?i#��G������lY4�!Þ?��@��?��;<��Z��=�;?[\�>ثO��>ƾ{������Ǔq=�"�>����ev�����Q,�[�8?٠�?���>
���������=�)w����?��?�����=�~��)c��	���w�)י=���9� ����6)�\�˾���0����Au=�F{>Vg@�7E����>��
��r߿sPؿ5�s�}����@'�>@��>��~�(�ؾؘ}�]b�8�9��\K��5g��J�>N�>;Ɣ�������{��j;��m���	�>��	�>�S��(��&���DY5<t�>���>Ҳ�>��� ݽ�b��?y\���=ο	���l��:�X?af�?oo�?1n?��7<i�v��{��h�Y2G?R�s?�Z?nf%�<]���7�z�s?8a���c�S+6�q�n���w>��3?�l>��Q�wl4>��=�F�>n�.>HKY�#�¿�Ů����{��?���? �3w?��?H� ?݆;���p����=���=TM?_89>��۾M���Gm<��*��3?��(?ˆ����]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?_$�>��?No�=b�>�c�=G�-�ok#>�"�=r�>��?��M?L�>W�=��8��/�=[F��GR�X$�:�C�	�>��a?�L?LKb>3��&2��!�Ivͽrc1��P��W@���,�Q�߽(5>��=>�>a�D��Ӿc�?*p�5�ؿ�i���s'�[54?��>��?I���t�a��V:_?�w�>�7�,��&���H�:��?G�?��?�׾u&̼S>��>K�>��Խ���邇���7>��B?�#��B��u�o��>`��?��@iծ?~i��	?���P��Ua~����7�b��=��7?�0�"�z>���>��=�nv�޻��W�s����>�B�?�{�?��>!�l?��o�O�B���1=9M�>Μk?�s?�Qo���h�B>��?"������L��f?�
@u@a�^?*��ҿ?����y�p�˾N�=��'>(w>�G2�/:>�{�<���=u�9���,>]��>k��>�>Շ�>�hq>���=�
���� �jJ��C�4>��a�? ���2�,�v�b!	�࠶��ھ!'����<��b��M!�M�����->�V?-�\?�B�?�>T�ɽE�K>Dy����;���&ߐ=yr�=nHG?/�>?=1 ?ʖ�=#���v�?Z�����8{��M�>��/>L�>�M�>��>&��<l>��h>n܂>O�)>���:E��;��=��->�!�>��>���>ʥV>k[>C|�����KDH�j�����t��.�?�����,��왿7�v�R7ᾴ��= r.?Pߣ=HE��HпQ���QXN?�0���6(�9s�D�u;C�(?PNI?��D>�U��.uɽ�Ls>�	ӽR������<���ľ@�7�K^�>��?G�f>�u>Ǜ3�\e8��P��|���i|>�36?M鶾vC9���u�N�H��cݾ�HM>ž>�D��k�u����� ui��{=x:?��?7���ⰾ9�u��C�� PR>^:\>�S=�i�=TXM>�bc�a�ƽ�H�d.=#��=��^>�?�e(> D�=y֢>Ù���K�QU�>C\B>P�'>�@?A�$?��䓑�L��+�a�u>w��>�r�>�,>C3I����=���>�@d>�g�4t��6F�ט@�T�W>qt�7`�Ɍy�	�c=�ޚ���=?��=����=�O =�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ߼�>5��ј�����"u�Rm=XY�><mD?�A����\�(�	?�u?���X���� ȿ�u�<"�>]��?K�?'�l�K����B����>���?�	X?R�t>�Hܾ0�e��ʋ>r??��S?U�>��AZ-�s?#�?�ۅ?z�>��?�z?x�>��<`Yھ3ꭿ6I�����>}���A>��D���[Io�����,�k�E"'���%���>�X�=��m>
����9���ݪ<n}��3g�������>:ś>,x=u(�>�i?�)�>��<��.��pv���&�����K?ز�?���j%n�ۺ�<��=2_�x:?(h4?h�W�c�Ͼ�Ѩ>�\?_ɀ?�[?X��>���J-��5鿿؂��z��<��K>�%�>�3�>ޅ���MK>��Ծ(lC�U��>Ð�>JΤ�+ھ�!���쫻�7�>5g!?J��>�ܯ=u� ?
�#?(�j>�'�>4aE��8����E�
��>>��>H?�~?y�?�ӹ��Z3�����桿H�[�>=N>��x?�T?.ʕ>@���ԃ���.E��5I��񒽈��?�sg?g\�p?�1�?/�??�A?�*f>����ؾ����u�>]�!?j�/�A��L&�9��:}?qP?���>o6����սOxּ���G����?.(\?6A&?u��*a���¾u@�<��"���T��u�;UsD�F�>Њ>ˍ�����=f>cѰ=UTm�EE6�G.g<yj�=U�>F��=<27��{���<,?'�G��ۃ���=d�r�cxD���>�JL>�����^?Bo=�9�{����ix��FU�� �?Ԡ�?:k�?Y����h��$=?
�?�?�!�>K��~޾V�ཱྀQw��}x�hw���>���>�~l�p����󙪿�F����Žd��o�?��>��>f�>�~z>�-�>sƞ��!�������3�^��e�D6�F/��H�N����ZV�<k�ƾ%|��帋>�齊��>5�?9�_>m�>	�>֐~��g�>��V>��>�S�>C�T>��>7>���9󅔽�R?i���M�'�m��%����uB?��d?<��>�Lm��l���r��@?��?�U�?HBv>ph�� +�t�?-��>����
?�0>=��ۀ�<nk��/������/�緎>�ؽ��9��M��Bf��i
?�?�����̾��׽}���o=AP�?"�(?O�)���Q�i�o���W��S�g�H1h��z��t�$�p�p� 菿�Z�����P�(��*=Q�*?��?���p�����"k��*?�5Nf>Q�>���>�Ծ>�{I>q�	���1�^��D'�����-6�>R{?z��>NQ?E�;?�8?'=O?�}>��j>T�q�4�D?�=�־>�5?�tV?��=?��??��K?��a?�ފ>��#��/���&��]�?�j?�@ ?t5?�q0?����]p���]>q�3�.(���呼��7=�@�����O���Y�>:�?_;�ʹ8�cU��M�h>�]8?��>��>aI��Û��-�	=��>5?��>����Xr�L�S�>@�?~�
�[�<��)>Z��=TNJ�0(: `�=�c�����=k攼��F��<<bY�=���=�Q������6;_fD;��<�l�>��?KȊ>�3�>5(��� �'��ï=�*Y>�Q>�>SRپ|�� '����g��8y>�q�?�^�?;h=' �=�m�=�����Y��,���潾��<�?XV#?�KT?���?�=?rl#?�>&;�MD���]��f����?��-?���>���:@;jv���;0�`
?�% ?]�c��S�gs(��$þ�3��=�V2�u0���W��i!>�o��;i�������?
֛?�듽�1�=�۾�e��0q����B?C��>�њ>[R?UM+���g�Yh�w)D>eW�>v^U?�%�>-�O?�>{?��[?�&T>ћ8��&���ϙ��f2���!>s@?ޡ�?h��?�y?�l�>a�>8�)��3�ah��P��w�TȂ�R#W=��Y>m��>f&�>�>@��=0�ǽ�8����>�8b�=x�b>e��>P��>#��>A�w>0�<��G?N��>=���bJ�&���J��1�I���u?
�?��+?�H=����sD�R���L�>���?"�?n*?�yW��V�=%9ؼ,����Jo���>�r�>!��>0�=ǘV=� >[��>a'�>m�:��E8��L���?�YF?��=�+��a����;M�,�ȓ�>����y���K�>��O�ع�>T ��V�>�F�D>�;��C�Ԯ���E�>s��W����?$��<��v�@�Q>.')>��;�Y3<���W�F��;q۹=��d�Y��\6����b�=�
ɝ�5��=�mH>��;��˾�}?�;I?{�+?��C?ָy>2<>ƚ3�˙�>�����@?�V>БP�����>�;�ë��� ��s�ؾ�x׾��c�(ʟ��I>�aI�)�>�73>�F�=�O�<��=�s=Î=�Q�=$�=�Q�=�e�= ��=c�>�T>�6w?Y���	����4Q��Y罌�:?�8�>�{�=}�ƾs@?�>>�2������lb��-?��?�T�?>�?Kti��d�>+��+㎽,q�=c����=2>$��=��2�6��>��J>���	K������4�?��@��??�ዿѢϿ�`/>tj->1��=j�T��/,��*@�G�p�_0W��#?�h6�����8�p>�=5��jľ��C=g�9>��=�����Y��I�=�c��Ǜ9=��`=M��>"�E>�Ϡ=����❭=�6C=��=��A>J'9�"�]��.���2=Z��=	lp>��!>��>?�c0? <d?�*�>�.n��9Ͼ�������>Wa�=�7�>��=u�B>?Ÿ>|�7?f�D?��K?y�>w��=�>f�>[�,���m��W�S������<@��?�׆?�ܸ>��K<a�A����U>�#�Ž2k?~S1??m�>����Ὶ�/��W�w���{ �=LO1>	<�\�<�6���U<�v]�G�h=�+?�^�>U��>��>wٞ>Αu>u��>��=�1K=<��<��=��z�?�����>��x��=����>+ý5R���
���
=��O;0.��)L��y!>%i�>�}�=��>8�ǽ�X8��/�>)��\�A��E(>�*�j�K�ZSL���z�
�3�F8���=O��>:�=�ݎ	?c��=�xU=�w�?x�}?I�r>vlA=�蔾8W��f��<�SD�|�>�0�>�����!B�E�4���6�Dp���>�>�׏>z�>��G>�N���#�>����;�^�?����0�R������ ����m��q>�PU?Ǐ����Q>�ql?�I?�3�?���>�|��s׾�e�>����U4>�
������Q=Y�?q�%?��>T���e�A�vA̾2��շ>FI�s�O�����î0�2��ҷ����>*�����о6%3��g��l����B�bYr�j��>��O?�?�7b�IU��ZSO����h���s?	wg?��>�J?5??�<���m�v��(a�=��n?���?j<�?>r��=�[~����>�?��?[�?��y?��N�n'�>Cr\�/O>>�ɽ��=�	">��=!�>�`?�W?��?ق��:D����+��n�S�X=�/�=p�>�z>��h>v4�=�r=6ľ=.V[>�I�>��>7�X>4(�>�p�>[��,���� ?60ɽ;6c>�1i?���>�0:=W_Y�����=�p���=#���EK�$I׽hUҼ��B>F_>4��>�Rտ퓝?���>��м�>l����<���1��>����x=�>,>�!e>N~�>�Ƞ>R"�>���=�伉���W>I���A#�\I:�rV��o�lV�>�)���]������ٽ5u�����������i�.䅿M�=�`81��?=	��p�m�!��.!��D?�U�>��0?ه�������U;>��>t�x>m��]
���f���>辟c�?�N�?u|b>j�>;+b?�?��f.#�Y�]��jo���:��2u��X��_��m���9��+�BzJ?F�p?3~/?	�=g�p>)�?�w����w�>��!���K�l��<��>��i?^��m¾�����{X���@=Cf?�Q}?/�>�F1��`f���%>�::?�U/?NYs?0�4?�=>?�����%?��3>e�?��	?�?5?0Q0?v�?��9>���=m��9PY=dz��I����̽�ʽ���X�=��i=�ᶺrx�;�;=���<����� ���O;�ʔ��d�<35=�=�P�=K��>\^`?b�>�}>�1?-�#�`<�*���'�>?b�==y�}f�����SоR�
>�Zn?���?�iS?�`7>��E�D�?�R�>E�>��1>\t>�b�>ML �,��Tv=�>C�">�=�읽�8���v��w��j==6G^>6��>{*|>�㍽��'>�y���#z���d>��Q�Һ���S���G��1��v�S�>-�K?k�?٪�=�Y�0��6Ef��6)?�]<?SNM?%�?#Г=Z�۾��9�w�J�\�9�>*�<F	�+���>$���:�'�:��s>U.��kR�<C	>� Q�����C���J�]GϾ��n>�t��[�U��˾+bþ��$�����6<����[��(u��~���*,?&��o<B꽥�	�m�=�?��>^��m�A>�U����3	��� ?I�>o�_����X�^�I�.���>>�R?T�p?��?�Ȣ�V��ِV�{��������=/l2?�߽>��?q�">ۮ�=����7�C�b�x�V���>g�?����A���y� �� 7��լ>/6�>UpB>N�?K�C?���>�)o?�P?�y?�;�>s6a�ˉ��?&?���?	�=D�Խr�T�D9��F���>�})?�B�q��>ڈ?E�?��&?�~Q?Ϯ?c�>[� �i:@���>O�>��W��^��	`>;�J?���>�0Y?YЃ?��=>ǃ5�4梾�穽Č�=�>m�2?�5#?+�?��>� ?�v*�G3�=�ױ>[4r?>�k?W?�X�=��?�_�=�ǚ>�!v�+ �>j�?a}�>�6X?�d?�(?S-?��<(��9k�����u����8��߻u�=�ɽ���B�cC0==;=>�=���=�Z(���Z;� `= Gr�zT�>/�s> ����1>�þ����A>*��W���1`��n0:�kJ�=���>�?�|�>�T"���=~��>�m�>�����'?D�?&�?��:�db�;�ھ��K��;�> �A?���=�m��w����u� �i=�n?�v^?{W������a?��^?�G��9��	ž��i����P?��?��(�B��>O�{?�vq?�\�>	�j��cn�؀��Q�]�+�Z�A	�=F��>A��d�8�>6?6��><JU>�}�=�c侍�v�-��A�?�P�?7��?�Պ?&�->��l�uݿ3r���L���^?
��>>���#?g�����Ͼ.@���(��H
�V
���%���S���u����$�\ۃ���ֽ���=��?�s?\q?��_?�� �y�c�!^����jV��$�� ��E�gE���C���n�\X��,��b��ZG=�D��YO��K�?P�?��d�{Q0?[xZ�& �ȸ���9>�Z��S�Y ��v�X��<ʗ�<7�a����Z<ȾZp?���>_�>��N?���  *��
���W��R��1Q>��>7r�>�	?�����	ý�MR��8վ��k��]���v>�cc?3rK?>�n?�i ��x0�����#!��h�yԥ���B>Q	>���>�BT�=��6�&�bl=�/-r���� W��� 
�5w=C2?�a�>�ל>
%�?��?/Z	��毾B�{�P�1�\y�<��>��h?"r�>,6�>Hӽeb �Wj�>	On?@�>t�>2��+�!�*:o�����>���>�r?��l>��v�U��p��uȎ��q6��o�=�"h?�ہ��i�&t_>�C?Pۣ<*gK<�י>�\���	$�6����O1�y��=y�?բ�=��E>"C��\���v��\b(?~�?ꑾ�c)�^i~>�� ?��>s[�>M��?���>CľE��^?�^?�*I?D@?�D�>j�=�잽m+Ƚ�N*���3=��>�_\>O ~=`]�=���qZ\��w�`D=�6�=�տ�V�����<�r��_��<���<Xi2>x�׿�I��{�$��X4Ӿ<���򈾿w��Ȑ���2�[�Ͼ#��d������)�n�g�v�O�!ej���C�X��?���?赭�(t��[đ���t�	��g
?�?1��b�BϾb���������`������_q�m�}��Lp�B�'?���˶ǿ
���1Aܾ� ?�- ?��y?����"���8�^!>Ȭ�<�H�����u����ο��^?���>����N�����>0��>�tX>�q>D��̞�" �<��?�~-?���>��r�ŕɿc�����<���?��@??��%��>��U=H��>џ	?XF>�-����#���d�>}��?��?JC=`@[�L�=�X/f?��;�iF���>Q�=N �=�G=��'�>>�>��.�(`<�^���	:>p��>�mϼp� ��%b��N<�T>t`ǽr��5Մ?+{\��f���/��T��U>��T?�*�>X:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?&�(?8ۿ��ؚ>��ܾ��M?_D6?���>�d&��t���=j6�����{���&V�~��=\��>d�>��,������O��I��T��=� �G�ſ��#�ڳ'�Q�<=�Z/�W ��Z��������b��zγ�ր�&�>��>C�>,��>>��>V��>�T?d	v?(�>3&>�B��y���#��6�=HCY�gZ�f����pn�������
��U���O)#��k"�n�ᾥ�����=�*���n��6o��Q�ܡH�{�l?S U>�8���E���Y>r��f����oU7��9 ��d��q�<�+ڣ?N<?`F��C��9�����~���`��1P?;]��[��`*��>��+�@$����4>Z�<�H�����l�_,?P�?gϿ��@���{@>�M�JZ=Fr(?a/�>D��<=�>!{"?���*�Խ��0>!>�٭>���>�Q�=󸮾�,�08?��S?��ؽ@��u�v>�j̾��t�_W�=|v>�5�B�39Q�v>9j�;�u��������o�[�=��V?ɐ�>|�(�������E*�aH=аx?�)?��>�:k?**B?R�<13��r�S�w���Do=EW?�i?&[>����ʜѾ�Ȩ���5?�d?,qL>��i��{뾕�/��Z�k�?��m?+?I���{��3������p5?��v?s^�xs�����M�V�h=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�$Þ?��@���?>�;<��T��=�;?m\�>�O��>ƾ�z������'�q=�"�>���~ev����R,�f�8?ݠ�?���>������Jj&>><B�mE�?�?�?�"�Տ>e�
��"���v��>^�8>?��=]0�=U����w׫���%�JZyP� 7z>��@�}(=�??[�3�y0����ܿ
�^�H�&��=/?N	y>���=��ͽ�9I���V��x?��ij��|���[�>��>IP��6����{��o;����i(�>��q�>��S����V���3<�ے>���>���>}��!���Ϳ�?ZV��<2οH���M���X?�c�?�i�?:f?+�:<�w���{�3m��0G?�s?�Z? �%��M]��[8��j?w_��oU`�َ4�CHE��U>�"3?�B�>d�-�G�|=#>x��>eg>�#/��Ŀ�ٶ�����F��?ˉ�?�o����>s��?xs+?�i�8���[����*�+��<A?�2>���,�!�0=�MҒ���
?(~0?
{�O.�\�_?)�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?h�?ص�� #�f6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�i	>���?�~�?Qj?���������U>	�}?�:�>�?;��=�.�>��=����7�!�W�#>���=��7�ޥ?�YM?o��>pr�=i�9��,/��F��R�p���C��U�>{va?�!L?�5c>����,Q4��:!���Ͻ��2�����A��r+��wܽ��5>�>>�h>�E�КҾ�k ?!o�xiٿ�ؗ�g�'���-?=�o>��?�����Έ�2���_?�}>̆��ᴿz������f�?t2�?m)?P�Ҿ�bk�#f/>3u�>��>I+ӽ����~����+>m�F?X�&�L���ZBp��>೽?��@$d�?�_r��	?`��W��Ic~��� 7�_�=��7?��9vz>V��>s�=.qv�������s�8��>�0�?�v�?���>'�l?[xo���B�MW3=�4�>ޏk?�n?�8x���a�B>��?j��9���N��f?'�
@vm@��^?������ֿzZ����ž+���B�=@6@��$�=e���9��=�!�=8!�3������ݠ>8��>?��>Ec�>�=�=H��>�d��u�#�7x����ʩQ�4w"�9���X��}�	�`���i���Ӿ��о/��bD�=���=T"B���!��f����=�U?MR?��p?�� ?rp�>` >'^���=
��x^�=��>�x2?շL?��*?���=�T��^hd�
倿�Ŧ����h��>hI>f��>���>�`�>�����F>�3>>��z>���=�)=�E޺N=��Q>��>�d�>N �>�W8>��>%,��-l��]�h�7}����뽃ϥ?�M��ƜN�����P��ᴾ�N�=T1?�@�=;���mQͿr~���2F?�p��b8�i�.�SR�=�.?�oT?,�>����MZ�)�>+sؽ>f��>���H�e�d.$���C>��?��d>p�]>��?�]JP��^���оMC>��j?M�u����#�v�������>) �>�����4��|����u��KH�����[�X?���>��ܽ�Y�h����L�T��=��>Af<84k>р>L.��dU��M��8�=}�2�N�>>O�>5�J>o�p=b�>��J��>���>�O*>�k�=W�>?�R+?�.��<t�9��Z��ߠ�=���>qM>w�>v�G�/S�<AR�>.i>��<�s���(q�dF����L>2�_���R�wg�*�=��;D�>'��=��1�c�5��A�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾFj�>k9��f��]6��ܗu�$y =2п>�nH?�n��\�W�d�>�?%?
��4�����ȿ��v�~��>Ӳ�?��?7m��m����?�|`�>�;�? �X?�gi>E!۾l][��-�>��??�^Q?P�>ڞ��(��y?���?L�?�tI>��?ʄs?�d�>.Zz��[/������Y����=���;&��>To>�<��YGF��ѓ��w��ڕj���CJb>��$=�ظ>-��b���]T�=����Y��d�t�>��p>��I>���>�� ?���>���>ɓ=�i��2܀�������K?(��?��� 8n����<�g�=M�^�S6?�J4?ץ^���Ͼ�ߨ>W�\?��?R
[?j]�>
��<;���࿿�w���ȕ<��K>[7�>�C�>����`UK>�վ�/D�p�>�Η>�Ţ�@@ھ�,��˦�>�>[g!?q��>��=%u ?=�/?�[�>u��>bE�x����� ����>`9?"4>?�+y?�?>0��ө/�u�������J��R>Ow?�U?���>�������Lt����5Xѽ��?czW?d􀽚�?��e?�*3?��6?��>gUG������㶽
#|>��!?����A�R&�����U?�?�5�>�W����׽D�A��d���?�\?�5&?�t���`��¾�/�<�)(��D��;u�E�x�>��>�������=Da>�.�=Hm�{6��lf<��=ܪ�>G��=T7��6��/=,?��G�ۃ���=��r�<xD���>�IL>����^?bl=��{�����x��)	U�� �? ��?Xk�?i��?�h��$=?�?T	?n"�>�J���}޾:�ྻPw�	~x��w�Z�>���>i�l���K���ٙ���F��S�Ž>��#�>���>���>�?�E�>-��>�j.���E�����g����G��F��A��T��1"�{)��U��Bx�D]ھJ@���d>I��=�L	?/�	?p��=x�>{;�>y��=�(�>d��>� �>���>���=+u�=�ۢ>�2H>VA�=�JR?����h�'���辙����1B?]pd?�/�>oi��������N~?��?�r�?�2v>o}h�*+��l?c>�>����n
?�\:=9�5V�<�R��\��xI��k&�9��>�L׽�!:�M��gf�}i
?a0?�⍼ӊ̾�3׽����uNo=�L�?��(?y�)�E�Q�g�o� �W�)S�c��h�d_����$���p�^쏿x^��� ��(�(�Lb*=��*?��?����#���)k��?�.}f>��>0�>��>hI>��	��1�� ^�4N'�vǃ�MH�>'W{?k�>�;?ϖ>?�ka?Sh.?M��>8�>p��{Z?�`N>ky�>���>��??U�(?�	?��>W%? �1>��=<!ھ�7�t�>w'?��(? T�>ue5?�l����=[#�=�+��E)�'?�0��=���=�q��-5���"E�=g?g���8�(^���-n>�7?F��>���> ҏ��O��
$�<_M�>b?jƏ>�� ��!r��j�#c�>�^�?do�r0=	*+>q6�=y���$�H^�=B�Ҽ���=@��D�<���<h �=I�=�W���$:[;`S�;Kt�<��>"�!?$;�>�?�>������辀���sd�=�l>
��>��>����4���)���.(a�=�M>f�?���?'��=�j>�g>k���W�v���׾`�;<S�?�r%?Ue_?o�?.4?�C?vޣ= �"�>���(������?��;?�Y�>�J��8��Aƺ�&9���-?��?�6���<�k�P��Mھr¾Ը#�k�!�Ro�`پ�AP��	̾x�2���r=��?O�?��[>�A������n��5���-J?�F�>k=�>�u(?�oK��rZ�Lx��j�>u�>n�g?7�>�`�?7�?STq?��M>5E��͌ƿ.s���L��(�>�/{?�6�?.F?��E?Q��>���>�o�<A����Ͼ��b�Rt�� ��b��=�J�>�S�>?z>�su=D��>�U��,?��Hͽ��=��=sܸ>}��>'-?o �>ڄ�>v�G?��>�X�� ���⤾ۻ����<�_�u?��?ȋ+?9=W����E�>=���D�>�p�?W��?�1*?��S�8��=�ּ嶾�q�� �>չ>72�>�ד=�F=�j>w�>���>%��\��g8�#M��?IF?d��=Z���xn�ߌz�mo��&�����.�h�%^P�^�M��Q�=Oq��A�ý�$���g�
�����.�����cz��� ?jd=lY�=��=�۽<m��M��<��/=UJ�<:~=6s�e�6=n��� ��H;��g0���;�И=�浹��ʾ�T}?9I?��+?��C?�/z>{.>>�3��C�>1���R)?7@U>~L��g��J�<��C������ؾ�־��c�m����n>��J�r<>>3>'��=Č<=K�=<o=wЌ=u�=���=ڕ�=}�=���=���=|[>��>�6w?U���	����4Q�zZ罥�:?�8�>b{�=��ƾk@?v�>>�2������tb��-?���?�T�?=�?*ti��d�>I���㎽�q�=N����=2>|��=j�2�^��>��J>���K��A����4�?��@��??�ዿ̢Ͽ7a/>���=�N�=��K��@9�8v�U�F�.yl��.?zn��aھ׭�=�q{>�dľ�R̾ S�=P�	>��:EV,���H���=N
��
|<��y="(m>.�X>���=Jw.�:�z=q��=y�Q>Y1�>N
�<��ͽuJ��G	<Fܴ=.�>c5>���>��?��8?�p?o2�>�ؽ�҉��"۾^a�>�:*>�[>c+�=�:n>Q�>��0?��>?��R?�î>�7�=���>��>��1��2���[��a�����<ӽ�??8f?�"�>��+>@E����a>F���`�FF?#?�q�>��>�����X#��B���D�="�����=�i>��N�`�L���7���վ�5=�?
�D?���>[Z�>	/k>�W�>���>G	>��<��=>��=y��=
�<6�b������<��L=W&����>\x0=.�ڽ+�c��%=qӄ>]G����=b��>a>���>	m�=������/>ʆ��Z�L����=�6��&B�i-d�9^~��/���6�ސB>OHW> R��6����?�vY>��?>Ȓ�?sIu? >���K�վzC���Md�mS��=�>�s=��h;���_�i�M�Ҿ�P�>6�>��>�P>�k'�0�7����=)=Ⱦ��;�6�>s��ZJ��r+��"}�{��G�����c��P�r-?!��9��=�fi?;N?>��?�T�>Q�9�	z��"�(>������>ȸ��![��X"�˳?��?�G?_����(��(̾�徽-��>�I�?�O�f���+�0��������C[�>~򪾷�о3�\k������F�B���r���>��O?�?�b��]���8O�����%���g?lg?�>�;?�N?������,�����=��n?���? 0�?1�
>Dn >@��}��>��?�0�?>�?7h?�o���$?�%?=q�=TU��7o>��9>���q�> �?��>��?߫��]ؾ�羷��D
N��t��=�>��>>�>�b�7�?ٽ����)�*>`W�>^��>[X�>(Ϣ>g��>�Y�� a�� ?H>��>1i-?���= "�]�����=���=_=:���C�c�սM۠�B�4��B��E�y����>ߎÿSQ�?,?�=��+�<�??1ӾSf�kO�>݄�=rw�'��>����
���?�f�><1��{%�>Ųw=��þ�%�=���E0/��?�K�C�JӾ�ߚ>����ʰV��c�0�=�%��m¾K���{�]��,�|�$�H�<��?ﲭ�B}��5�����&��>�f�>E�1?&�h������,>���>P��>����{��	��Ɩ�(�?�[�?�$f>��>.�V?O�?p,��%,�f	X��t��?�m6e���_�Tݍ��Ѐ�T����Ƚ�Ha?�y?	Q@?)��<|�x>]�?9�%����酈>�j.�Oq9��|E=c�>�譾�d���پ=�ž�����N><�p?pV�?��?�bS��!�<�+>�a*?n9?O�}?8�<?��@?�eY�w�9?;��>@�?ټ�>%R6?��?~�>8�=0�
>P1��G�D>�o��f�1'ν���z�<cb<=�،=8��<Φ�<.�0��qo��� =dɺ�tL8�"Ȑ�<!�=�=jW=��S=+̨>�Tf?�z?�y�>^n%?'
���Qa����B-?�p	=|�5� �����~X��`X>5F{?a��?��q?�8�> �Q���n�a�=�$�>|��=�	�>;<�>:�������"==�=�q�=��=ZA�<&C��!�Cz������Z!>b��>9N|>�Ǝ�̸&>����_;z�¥d>�P�u�����T���G���1��v����>[�K?:�?���=���(��Q;f��(?�:<?9hM?x�?y�=\A۾��9�(�J�n�c��>��<t������X$����:�%K2;8=t>�՞�w��,�b>����޾;In���I��o羧�O=�����Q=����վT �G��=��>S����� ����s���'J?"�d=�#��,~U�gB��(�>Z�>�(�>kX:�;T{�ݡ@�����Ӕ=l��>�;>7������G�����H>Z]_?u?~6x?�o��{�h��~V�ނ��/ݾ썔=��$?ס�>{F%?8�x>g%�=(������vb�1uZ��V�>?e�>�6=�"R��K�+�,�0��>��>5!>��?��B?}��>�b?u4?5� ?�G�>H�ۼ� �� 4&?���?��=��ӽ�U�9���E����>ӕ)?��A��З>�?��?g�&?�FQ?؉?�+> ��@�N��>H�>��W��W��Ld_>��J?��>>!Y?�̓?��>>�j5��n���+��F�=l>~�2?�#?k�?��>�.?�u��k��҇?��*?[U�?��
?���o`(?� ?�_?�>r�B]�=�.?H��>��A?D�D?)*R?���>8!��[Q=~��<X"�� >�<�"<[1�<���<� ���}S���=�44<𚼣��<@��3����[��s=�j�>��s>�啾iA1>��ľo��*�@>^����雾���P:�_F�=K]�>'�?
��>�H#�X;�=�ͼ>9i�>����0(?:�?��?i�;��b��ھRUK��/�>IB?���=2�l�|����u�(�g=��m?؊^?�W�V��O�b?��]??h��=��þ{�b����g�O?=�
?0�G���>��~?f�q?U��>�e�+:n�)��Db���j�)Ѷ=[r�>LX�S�d��?�>o�7?�N�>.�b>$%�=iu۾�w��q��h?��?�?���?+*>��n�Z4�~��wJ��u^?���>Z<����"?�B����Ͼ4P��$����A��g���<��Dx��&�$��ڃ��׽�=~�?s?TYq?Y�_?״ �5�c��1^�:
��PhV��&� $���E�A"E��C���n�_��0�����S�G=�gþd�"H�? �>�厾���>�����~;�7���)j>2
[����;�z>7�^=��E>B%2=ZU��I뫾�G��f?�#?�H ?��j?��q�V�
��&j��#*����o�>���>�A>�oT?��;w���ܼ�x ��t)�X߻��v>?~c?�K?��n? E�p-1�	�����!���/��P��߫B>E>�É>��W����k/&�H>���r�����h��3�	�,�}=U�2?A�>YȜ>�K�?��?v	��q���Rx�k�1���<j5�>�i?9�>n��>]Oн�� �Sg�>F�l?���>Ů�> ����!�2Uz��6Ƚ*��>r�>��>��p>�*��K[�[b���u����7���=�gh?����`�/\�>X�P?�����!e<=��>"�w��� ��3��a'�n��=ɶ?���=3�<>r�ž����z�Vt��,l)?N�?�ْ���)�g�~>�c"?�>m�>�#�?&��>�;¾�?&�30?c�^?o�I?�_A?��>&=���zwȽ�&�3-=��>;�[>��m=�S�=�����\�����B=e��= !˼����U<[D��B�J<���<�3>�iۿhBK�[vپ����8
�!ш�����k�����ZZ��a���x��g���&�SV�04c�'���y�l����?�:�?�^��������􈀿7�����>kpq�>%��߫�4��`���z�ྜ����b!�H�O��i���e���-?����\)Ŀ���Io�R�?\�P?]�y?<�
��-��#���-e��c	�;P�M�0���ѿ�צ�q^>?D��>�-ʾ$=�=^�>��>}Q>ᷴ>�ѾIR\����=�m�>�?��
?-��+ ӿV�ȿOߘ�Y�?�@�CA?�(�f��K�c=�X�>YM	?�N=>��1�Q��⠰�,��>��?�$�?�T=��W�wf���e?}��;F������U�=/Σ=ŏ=�-�>@J>W�>����Y@�۲߽�<3>Q�>��!�ND�(\��j�<�\>
fԽ����5Մ?-{\��f���/��T��U>��T? +�>X:�=��,?P7H�^}Ͽ�\��*a?�0�?��?�(?;ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�
��=�6Ἀ���p���&V�e��=\��>j�>͂,�����O�2I�����=�6�ƿ��$�����=��޺�D[�+�罁Ӫ��T�q"��	Yo������h='��=8�Q>�g�>�W>�.Z>eW?Z�k?[�>t�>�~�:o��	ξ����8��]���������[ڣ�K�d�߾��	������$�ɾ��f�_�S��yO��C����!�����N��a�?�P�>=/�[�����>��ɾ�3��C��߭�]�:�?���΁�MӁ?���>�����9P������n�=�ر���-?B'ҽj�%�ڻ���9=�M%�?^2��"�>5؃>����@�����jl0?1F?�.������
*>ó �߶=Ƭ+?��?��e<�g�>0>%?�*�G���[>��3><	�>���>5�	>�뮾?�ڽwq?ET?������>p/���Bz�شc=��>Z+6���[>z�<�Ҍ�ږO�c��>	�<�$W?{��>R�)�&��Ew���U��==!�x?�?�R�>�pk?��B?~�<�I����S����Cx= �W?�$i?�>���-'оnr���5?�e?��N>Hmh�`��T�.��S�[�?Ŀn?�`?�`��][}�������`6?��v?s^�qs�����W�V�=�>�[�>���>��9��k�>�>?#��G����sY4�!Þ?��@}��?s�;<S����=�;?p\�>ëO��>ƾ�z��������q=�"�>	���eev�����Q,�[�8?⠃?m��>��������=
l�����?��?_������<����l��� ���<� �=�S�(	��}�ɥ6�?�ž�?��Ν���Nj�>�7@by�7��>1�7��⿳ZϿ^S��
�Ѿ5Kl�1l?Ϳ�>����㡾߭j���s�6G�J�G�̐��K��>R�>�%��h��
�z��7�(�t�>`nr��J�>�K��a¾���b��<zQ�>2��>�<�>T�n�����-�?�����ο�#�����DG\?7>�?�Ȁ?�?,�A���~�eG��S�.��D?�o?�#]?�	�+�X�[�>���e?q۱�2LW�}%:�GuT��W>=3E?�P�>�#���=r��=���>�>L�:��ܾ��]�����2*�?��?�Y��2�>H�?�q0?�������˾��9�-�r���B?���=�g����$�JP�wx����>	-?X� ���_?��a���p��-�V�ƽ١>t�0��C\��������Te����PPy�=�?�`�?i�?���I#�-%?��>6����)Ǿ��<�t�>�$�>[KN>�u_�t�u>l����:�XT	>]��?�{�?Ha?˙�������t>��}?W$�>��?�o�=�a�>qc�=j񰾼�,��k#>Q#�=�>��?��M?L�>6W�=��8��/�![F��GR�@$�(�C��>m�a?ȂL?Kb>����2��!�guͽc1��P�jX@��,��߽;(5>k�=>�>�D��Ӿ��?Np�8�ؿ�i��"p'��54?.��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>=�>�I�>@�Խ����\�����7>0�B?W��D��t�o�y�>���?	�@�ծ?ji�	?���O��a]~�<����6����=��7?{,��z>���>��=�kv�ӹ���s����>aB�? {�?
��>F�l?��o���B�b2=TN�>=�k?�r?Jp�A�F�B>��?��������J��f?��
@@t@��^?E��<���aq�����eX�����==���#a�=;����>ʖ�=<�1�`B=���=`Qo>�)R>�+:>�
j>S�q>
�6>^����Y���������+aI��?�l���3�<2�ӾC;;��~h��Gþ��X��%�\z��	$��ګ���R����=9�U?W[R?>p?�� ?�4~��f>����U =�0"��f�=^�>�{2?��L?�K*?�[�=����~�d����A�������IE�>��K>(T�>��>�,�>��9X�I>>�=>��>�F >M*)=����8=��N>N�>���>1�>ft�>�A2�]�¿ܓ���F`� %K��+�f�?�K�Ņ��ǧ��4�o����x���Z�?pf�>�̒��x˿�A��OE@?Gd~��?�V=Y j=_ .?���?o�<������=Fs�>3����Z��>_M>�G����[�mF=��B?w�f>h�t>�3��h8�#�P��l��4�|>;6?����5�9�&�u��H��sݾ�?M>_�>��C�h|�������"Yi��@{=�z:?Yx?׊��7Ӱ��'u�'N���R>�t\>Ӯ=V�=U�M>�bb�GQǽ��H�D�-=���=I5_>f�?xs>9�*>��>_a�� k�|��>�7>7��>Z�Q?<�#?�g�D���J�C��?s���=c�>٥�>@�S>B�Ƚ%�<2�>�>�Y���XJ<Xq���1��
O>�<X�h��~����&<<)k<�q>Z=����<�����<�~?���(䈿��e���lD?S+?_ �=
�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž5Ǣ�ɔ	�/)#�jS�?��?��/�Zʋ�=l�6>�^%?��ӾZh�>|x�|Z�������u�|�#=N��>�8H?�V��O�O�\>��v
?�?�^�۩����ȿ!|v����>R�?���?q�m��A���@����>9��?�gY?Hoi>�g۾F`Z����>ǻ@?�R?�>�9�:�'���?�޶?ϯ�?�I>5��?��s?qq�>�y�\/��)��M�����=ihp;�s�>]v>����YF��Փ��d��֦j�"��2�a>�$=H�>\佂<���=� ���F��7af����>�jq>9�I>(�>�� ?s�>���>��=�]��n���䭖���K?���?-���2n��N�<Z��=)�^��&?�I4? k[�}�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��H��<��K>*4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��WS��GB�>�e!?���>�Ү=b ?�$?Wo>oI�>�oE���B�C�'X�>�j�>��?�b~?I�?�L����2�?
���t���mY�vMQ>Q�x?�?4��>���M������>�F��Ǐ���?�wg?�rϽ�?���?��=?��A?8�d>�����׾�����>��!?%s���A��E&��>�T|?�X?5��>���tֽj=ּ���������?�H\?�D&?Ǧ�,a��þڰ�<�X#�.�G�r� <לF��>�>{����=�h>�R�=Ipm��6���k<<1�=�%�>`�=
�6�D#��0=,?ܿG�|ۃ���=��r�<xD���>�IL>����^?el=��{�����x��	U� �?���?Zk�?^��?�h��$=?�?R	?n"�>�J���}޾8���Pw�~x��w�S�>���>Ǣl���I���ٙ���F��b�Ž��۾:�'?�T^>��>e�?�=�:�>GR)�0S��fܾ��w�t�A$�e30��a7��A�'�վ)�۾GW��a&;�P;��d#>�M�����>�]?cd�>,�b>>2P>�-�<�֨>S��=���>���>��;oǊ>���>f�=�wl�QLR?������'����ò��N3B?�pd?�/�>�	i�K������~?-��?�r�?�:v>�}h�@++��n?�>�>q���o
?-@:=���L�<S��f��4�������>H׽�:�)M�mnf��i
?`0?Q��!�̾C=׽����.q=fU�?��(?@�)�g�Q��o�)�W�'S��P���g�rg���$�}p�V叿S��#��ˡ(�e�(=�*?i�?\��А�O묾>k�}?�u�f>p�>��>�>�tI>,�	�"�1��^��='�����`�>�S{?Bc�>x�K?��>?ۣP?��M?��>���>�7���J�>)Sv<l-�>Ę�>�9?�.?R{,?�?�-?NZ>Jؽm���P��)�?��?pP?B?V�?ģ�����23����Z�y���c��o�=�E�;��ҽ�i#�[�=�_e>\d?R��t8�������k>>�7?��>F�>�@��i���-U�<���>�
?S��>Oc��k r������>_��?Xy��:=�*>C��=�J��+�J��=s���F;�=�;��l%<�Qp%<���=^��=J4���i빡�1;k��;>�<lx�>h�?B��>ꩌ>����Y��}
��=(�a>��Y>�q >�4̾���{얿��h��r>��?c�?<8�=�}�=wz�=VL���qþ�
�h���"�
=��?N*%?MY?Gԑ?A�5?��?
�>���{���丄��H��k~?z%,?_>�����1�}[ ��3?��>%	R�T/C��T-��7�����8?w=9m*����{۵��)��6=)���
B�7��?cĖ?LI����0���Ø���펾�cD?7�>r��>|��>��I��l���&�_�,>���>�TS?�'�>�)X?M!�?[�a?U�>�93�%[��ډ���׽�F>-�7?��c?V�?3a�?�G>2N>-�g��Tݾ h��ٰ<�U�;���=�<��>�u=s#�>�*�>YP]>z����5��Hh==6�<47�=e4�>D�>��>3�>CS�=hH?� �>\���3��ꤾl:���3=�Mu?��?��+?�#=ܘ���E�����?��>�X�?=�?!L*?+
S����=�
߼R���q�(;�>:�>�4�>~�=��D=Ű>���>S��>�N��;��<8�:KG���?�E?�4�=��ſ�kc�-kg��룾��d=s䐾�3��ͫ�6Z��ܑ=�Ԍ���'��X���P�kC��b/��OG��rB��QYe��7�>Q��<s(>�=35Ļ����]��<���#%=���<Љ����`=�.���s<����<��=;�=�3���;�}?��G?�*?��C?'�x>�8>�/�� �>�V��K�?�lP>+S�������?�o~��ߪ����پ��־@c�����~A>'K���>ؘ2>(��=6e<��=R=l=�=�Ϲ>�#=k�=g�=���=���=X�>w�>�6w?p���貝��3Q�B\罸�:?u8�>Fz�=��ƾf@?��>>�2��A����a�<-?=��?�T�?]�?tsi�)e�>#��o鎽qt�=N���{@2>C��=��2����>��J>q���J������4�?c�@�??�ዿ��Ͽ�_/>S�3>[�>;�R��q1���Y��9b��,Y�1o!?4�;��˾��>1�=r߾��ƾ �"=�63>�x\=V��I�[�m.�=���f;=oKj=��>3�C>�/�= Ų���=��G=���=J�P>�^9�I5��@1�J�8=��=\�c>��&>���>�?w*4?�3n?�M�>ȋi�`z���ۡ����>��,=S?�>X �>�׳>���>���>=o)?wW?���>3|}>@ƪ>GԾ>n[徔Wn�+��}�¾AӍ>nx?��?��?��<����+�A�<�5�$���>'�>JL?v�0>�U����7Y&���.������4��+=�mr��QU�J���Km�.�㽗�=�p�>���>��>7Ty>�9>��N>��>��>�6�<}p�=�ጻ��<� ��t��=ҝ����<�vż����Vu&�%�+�ݏ��w�;���;��]<���;�l�={�>.�>���>m��=���l�.>\���YM����=���	�A�߼d�̜~�/.��p=� �;>��N> ���IL����?o�S>97?>t�?K�t?,>ө��5׾����\�,�Z�.c�=�b>��?��9�[�]�g?N��Ҿ9 �>�k>?��>��=h@��s:���>�C �X�4��O�>=]ʾ�ţ=Ŋ�%��U͈�o˴��
��l�ν��:?�I��C�>S:P?2TP?��?��k>Z����X�9�ֽ�wx��25>����/�����;S	?�_"?��?�}A�(�;��D̾Ѿ��߷>�0I�;�O����R�0�y��·�Ŕ�>��о�3��a��������B��3r�z�>˳O?��?�ib��T���OO����fi?�mg?��>P@?i1?sk���z�]�����=��n?��?�5�?L>yd�=Lo�����>n�?둕?�?��i?;�A�ɀ�>�Ƨ<p�(> m��Q��=�:>�9k=E{�=��?T�	?x�?��}�[�� ��IL�ԑW�`�=M-�=��>���>�l>��=t�=q)�=�O>6��>���>X�b>T�>�Ӂ>yľU�ʾ��?���=�5�>9��>��P>Nz��pEz�m��<M�ý��p�1�l%�=�짾IB=�_�=�l��x*#>�� ?"�ſ��O?��>�v��rw"?����� [��@�>�%�=�R�Ђ�>9=7#�>z��>ɨ�>���><�	>F��="SӾ�>���~d!�%C��R�z�Ѿ@}z>ߪ���&���E����AI��o��Kk��j�[-���==�_ڽ<E�?����Ȼk�8�)������?�]�>>6?�ی�o"��Ț>��>�ɍ>E��Ǝ���Í�Y]�D�?���?c>.�>��W?��?@\1�B73��uZ�l�u��A���d���`�⍿�����s
��<��[�_?��x?�kA?�<Doz>�}�?b�%��{��J�>��.��;���;=P�>F<��W�`�°Ӿ�þ��$�E>g�o?�"�?/=?8V��O��[>z�/?�A0?Z�|?9?Z� ?��?��w?P�;>r?u�?��<?�0?-.?B�3>A�>��=��>�@.���R��Em��²�Q�>�VrC�Aq8=��6=y5=f��=[�H=b�<}#���<[�?��?���=���=��>5��>��\?W��>�ٔ>/;?�Y'���=�+>��J�)?�Sq=t�������f����ھ�8�=Jzh?�^�?d�P?7 v>�})��qj�A��=���>�o:>ɬs>@�>x���X0��R*=
N>�<>D�=�B(�����q(�^>��<��;��0>4��>[1|>���F�'>X{��01z���d>��Q�0̺�_�S�D�G���1���v�VZ�>��K?��?G��=_龔)���Hf�,/)?]<?)OM?��?��=(�۾D�9�u�J�Z?���>`V�<K�������#��x�:��0�:ƿs>�0��kR�<C	>� Q�����C���J�]GϾ��n>�t��[�U��˾+bþ��$�����6<����[��(u��~���*,?&��o<B꽥�	�m�=�?��>^��m�A>�U����3	��� ?I�>o�_����X�^�I�.���>>�R?T�p?��?�Ȣ�V��ِV�{��������=/l2?�߽>��?q�">ۮ�=����7�C�b�x�V���>g�?����A���y� �� 7��լ>/6�>UpB>N�?K�C?���>�)o?�P?�y?�;�>s6a�ˉ��?&?���?	�=D�Խr�T�D9��F���>�})?�B�q��>ڈ?E�?��&?�~Q?Ϯ?c�>[� �i:@���>O�>��W��^��	`>;�J?���>�0Y?YЃ?��=>ǃ5�4梾�穽Č�=�>m�2?�5#?+�?��>� ?�v*�G3�=�ױ>[4r?>�k?W?�X�=��?�_�=�ǚ>�!v�+ �>j�?a}�>�6X?�d?�(?S-?��<(��9k�����u����8��߻u�=�ɽ���B�cC0==;=>�=���=�Z(���Z;� `= Gr�zT�>/�s> ����1>�þ����A>*��W���1`��n0:�kJ�=���>�?�|�>�T"���=~��>�m�>�����'?D�?&�?��:�db�;�ھ��K��;�> �A?���=�m��w����u� �i=�n?�v^?{W������a?��^?�G��9��	ž��i����P?��?��(�B��>O�{?�vq?�\�>	�j��cn�؀��Q�]�+�Z�A	�=F��>A��d�8�>6?6��><JU>�}�=�c侍�v�-��A�?�P�?7��?�Պ?&�->��l�uݿ3r���L���^?
��>>���#?g�����Ͼ.@���(��H
�V
���%���S���u����$�\ۃ���ֽ���=��?�s?\q?��_?�� �y�c�!^����jV��$�� ��E�gE���C���n�\X��,��b��ZG=�D��YO��K�?P�?��d�{Q0?[xZ�& �ȸ���9>�Z��S�Y ��v�X��<ʗ�<7�a����Z<ȾZp?���>_�>��N?���  *��
���W��R��1Q>��>7r�>�	?�����	ý�MR��8վ��k��]���v>�cc?3rK?>�n?�i ��x0�����#!��h�yԥ���B>Q	>���>�BT�=��6�&�bl=�/-r���� W��� 
�5w=C2?�a�>�ל>
%�?��?/Z	��毾B�{�P�1�\y�<��>��h?"r�>,6�>Hӽeb �Wj�>	On?@�>t�>2��+�!�*:o�����>���>�r?��l>��v�U��p��uȎ��q6��o�=�"h?�ہ��i�&t_>�C?Pۣ<*gK<�י>�\���	$�6����O1�y��=y�?բ�=��E>"C��\���v��\b(?~�?ꑾ�c)�^i~>�� ?��>s[�>M��?���>CľE��^?�^?�*I?D@?�D�>j�=�잽m+Ƚ�N*���3=��>�_\>O ~=`]�=���qZ\��w�`D=�6�=�տ�V�����<�r��_��<���<Xi2>x�׿�I��{�$��X4Ӿ<���򈾿w��Ȑ���2�[�Ͼ#��d������)�n�g�v�O�!ej���C�X��?���?赭�(t��[đ���t�	��g
?�?1��b�BϾb���������`������_q�m�}��Lp�B�'?���˶ǿ
���1Aܾ� ?�- ?��y?����"���8�^!>Ȭ�<�H�����u����ο��^?���>����N�����>0��>�tX>�q>D��̞�" �<��?�~-?���>��r�ŕɿc�����<���?��@??��%��>��U=H��>џ	?XF>�-����#���d�>}��?��?JC=`@[�L�=�X/f?��;�iF���>Q�=N �=�G=��'�>>�>��.�(`<�^���	:>p��>�mϼp� ��%b��N<�T>t`ǽr��5Մ?+{\��f���/��T��U>��T?�*�>X:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?&�(?8ۿ��ؚ>��ܾ��M?_D6?���>�d&��t���=j6�����{���&V�~��=\��>d�>��,������O��I��T��=� �G�ſ��#�ڳ'�Q�<=�Z/�W ��Z��������b��zγ�ր�&�>��>C�>,��>>��>V��>�T?d	v?(�>3&>�B��y���#��6�=HCY�gZ�f����pn�������
��U���O)#��k"�n�ᾥ�����=�*���n��6o��Q�ܡH�{�l?S U>�8���E���Y>r��f����oU7��9 ��d��q�<�+ڣ?N<?`F��C��9�����~���`��1P?;]��[��`*��>��+�@$����4>Z�<�H�����l�_,?P�?gϿ��@���{@>�M�JZ=Fr(?a/�>D��<=�>!{"?���*�Խ��0>!>�٭>���>�Q�=󸮾�,�08?��S?��ؽ@��u�v>�j̾��t�_W�=|v>�5�B�39Q�v>9j�;�u��������o�[�=��V?ɐ�>|�(�������E*�aH=аx?�)?��>�:k?**B?R�<13��r�S�w���Do=EW?�i?&[>����ʜѾ�Ȩ���5?�d?,qL>��i��{뾕�/��Z�k�?��m?+?I���{��3������p5?��v?s^�xs�����M�V�h=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�$Þ?��@���?>�;<��T��=�;?m\�>�O��>ƾ�z������'�q=�"�>���~ev����R,�f�8?ݠ�?���>������Jj&>><B�mE�?�?�?�"�Տ>e�
��"���v��>^�8>?��=]0�=U����w׫���%�JZyP� 7z>��@�}(=�??[�3�y0����ܿ
�^�H�&��=/?N	y>���=��ͽ�9I���V��x?��ij��|���[�>��>IP��6����{��o;����i(�>��q�>��S����V���3<�ے>���>���>}��!���Ϳ�?ZV��<2οH���M���X?�c�?�i�?:f?+�:<�w���{�3m��0G?�s?�Z? �%��M]��[8��j?w_��oU`�َ4�CHE��U>�"3?�B�>d�-�G�|=#>x��>eg>�#/��Ŀ�ٶ�����F��?ˉ�?�o����>s��?xs+?�i�8���[����*�+��<A?�2>���,�!�0=�MҒ���
?(~0?
{�O.�\�_?)�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?h�?ص�� #�f6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�i	>���?�~�?Qj?���������U>	�}?�:�>�?;��=�.�>��=����7�!�W�#>���=��7�ޥ?�YM?o��>pr�=i�9��,/��F��R�p���C��U�>{va?�!L?�5c>����,Q4��:!���Ͻ��2�����A��r+��wܽ��5>�>>�h>�E�КҾ�k ?!o�xiٿ�ؗ�g�'���-?=�o>��?�����Έ�2���_?�}>̆��ᴿz������f�?t2�?m)?P�Ҿ�bk�#f/>3u�>��>I+ӽ����~����+>m�F?X�&�L���ZBp��>೽?��@$d�?�_r��	?`��W��Ic~��� 7�_�=��7?��9vz>V��>s�=.qv�������s�8��>�0�?�v�?���>'�l?[xo���B�MW3=�4�>ޏk?�n?�8x���a�B>��?j��9���N��f?'�
@vm@��^?������ֿzZ����ž+���B�=@6@��$�=e���9��=�!�=8!�3������ݠ>8��>?��>Ec�>�=�=H��>�d��u�#�7x����ʩQ�4w"�9���X��}�	�`���i���Ӿ��о/��bD�=���=T"B���!��f����=�U?MR?��p?�� ?rp�>` >'^���=
��x^�=��>�x2?շL?��*?���=�T��^hd�
倿�Ŧ����h��>hI>f��>���>�`�>�����F>�3>>��z>���=�)=�E޺N=��Q>��>�d�>N �>�W8>��>%,��-l��]�h�7}����뽃ϥ?�M��ƜN�����P��ᴾ�N�=T1?�@�=;���mQͿr~���2F?�p��b8�i�.�SR�=�.?�oT?,�>����MZ�)�>+sؽ>f��>���H�e�d.$���C>��?��d>p�]>��?�]JP��^���оMC>��j?M�u����#�v�������>) �>�����4��|����u��KH�����[�X?���>��ܽ�Y�h����L�T��=��>Af<84k>р>L.��dU��M��8�=}�2�N�>>O�>5�J>o�p=b�>��J��>���>�O*>�k�=W�>?�R+?�.��<t�9��Z��ߠ�=���>qM>w�>v�G�/S�<AR�>.i>��<�s���(q�dF����L>2�_���R�wg�*�=��;D�>'��=��1�c�5��A�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾFj�>k9��f��]6��ܗu�$y =2п>�nH?�n��\�W�d�>�?%?
��4�����ȿ��v�~��>Ӳ�?��?7m��m����?�|`�>�;�? �X?�gi>E!۾l][��-�>��??�^Q?P�>ڞ��(��y?���?L�?�tI>��?ʄs?�d�>.Zz��[/������Y����=���;&��>To>�<��YGF��ѓ��w��ڕj���CJb>��$=�ظ>-��b���]T�=����Y��d�t�>��p>��I>���>�� ?���>���>ɓ=�i��2܀�������K?(��?��� 8n����<�g�=M�^�S6?�J4?ץ^���Ͼ�ߨ>W�\?��?R
[?j]�>
��<;���࿿�w���ȕ<��K>[7�>�C�>����`UK>�վ�/D�p�>�Η>�Ţ�@@ھ�,��˦�>�>[g!?q��>��=%u ?=�/?�[�>u��>bE�x����� ����>`9?"4>?�+y?�?>0��ө/�u�������J��R>Ow?�U?���>�������Lt����5Xѽ��?czW?d􀽚�?��e?�*3?��6?��>gUG������㶽
#|>��!?����A�R&�����U?�?�5�>�W����׽D�A��d���?�\?�5&?�t���`��¾�/�<�)(��D��;u�E�x�>��>�������=Da>�.�=Hm�{6��lf<��=ܪ�>G��=T7��6��/=,?��G�ۃ���=��r�<xD���>�IL>����^?bl=��{�����x��)	U�� �? ��?Xk�?i��?�h��$=?�?T	?n"�>�J���}޾:�ྻPw�	~x��w�Z�>���>i�l���K���ٙ���F��S�Ž>��#�>���>���>�?�E�>-��>�j.���E�����g����G��F��A��T��1"�{)��U��Bx�D]ھJ@���d>I��=�L	?/�	?p��=x�>{;�>y��=�(�>d��>� �>���>���=+u�=�ۢ>�2H>VA�=�JR?����h�'���辙����1B?]pd?�/�>oi��������N~?��?�r�?�2v>o}h�*+��l?c>�>����n
?�\:=9�5V�<�R��\��xI��k&�9��>�L׽�!:�M��gf�}i
?a0?�⍼ӊ̾�3׽����uNo=�L�?��(?y�)�E�Q�g�o� �W�)S�c��h�d_����$���p�^쏿x^��� ��(�(�Lb*=��*?��?����#���)k��?�.}f>��>0�>��>hI>��	��1�� ^�4N'�vǃ�MH�>'W{?k�>�;?ϖ>?�ka?Sh.?M��>8�>p��{Z?�`N>ky�>���>��??U�(?�	?��>W%? �1>��=<!ھ�7�t�>w'?��(? T�>ue5?�l����=[#�=�+��E)�'?�0��=���=�q��-5���"E�=g?g���8�(^���-n>�7?F��>���> ҏ��O��
$�<_M�>b?jƏ>�� ��!r��j�#c�>�^�?do�r0=	*+>q6�=y���$�H^�=B�Ҽ���=@��D�<���<h �=I�=�W���$:[;`S�;Kt�<��>"�!?$;�>�?�>������辀���sd�=�l>
��>��>����4���)���.(a�=�M>f�?���?'��=�j>�g>k���W�v���׾`�;<S�?�r%?Ue_?o�?.4?�C?vޣ= �"�>���(������?��;?�Y�>�J��8��Aƺ�&9���-?��?�6���<�k�P��Mھr¾Ը#�k�!�Ro�`پ�AP��	̾x�2���r=��?O�?��[>�A������n��5���-J?�F�>k=�>�u(?�oK��rZ�Lx��j�>u�>n�g?7�>�`�?7�?STq?��M>5E��͌ƿ.s���L��(�>�/{?�6�?.F?��E?Q��>���>�o�<A����Ͼ��b�Rt�� ��b��=�J�>�S�>?z>�su=D��>�U��,?��Hͽ��=��=sܸ>}��>'-?o �>ڄ�>v�G?��>�X�� ���⤾ۻ����<�_�u?��?ȋ+?9=W����E�>=���D�>�p�?W��?�1*?��S�8��=�ּ嶾�q�� �>չ>72�>�ד=�F=�j>w�>���>%��\��g8�#M��?IF?d��=Z���xn�ߌz�mo��&�����.�h�%^P�^�M��Q�=Oq��A�ý�$���g�
�����.�����cz��� ?jd=lY�=��=�۽<m��M��<��/=UJ�<:~=6s�e�6=n��� ��H;��g0���;�И=�浹��ʾ�T}?9I?��+?��C?�/z>{.>>�3��C�>1���R)?7@U>~L��g��J�<��C������ؾ�־��c�m����n>��J�r<>>3>'��=Č<=K�=<o=wЌ=u�=���=ڕ�=}�=���=���=|[>��>�6w?U���	����4Q�zZ罥�:?�8�>b{�=��ƾk@?v�>>�2������tb��-?���?�T�?=�?*ti��d�>I���㎽�q�=N����=2>|��=j�2�^��>��J>���K��A����4�?��@��??�ዿ̢Ͽ7a/>���=�N�=��K��@9�8v�U�F�.yl��.?zn��aھ׭�=�q{>�dľ�R̾ S�=P�	>��:EV,���H���=N
��
|<��y="(m>.�X>���=Jw.�:�z=q��=y�Q>Y1�>N
�<��ͽuJ��G	<Fܴ=.�>c5>���>��?��8?�p?o2�>�ؽ�҉��"۾^a�>�:*>�[>c+�=�:n>Q�>��0?��>?��R?�î>�7�=���>��>��1��2���[��a�����<ӽ�??8f?�"�>��+>@E����a>F���`�FF?#?�q�>��>�����X#��B���D�="�����=�i>��N�`�L���7���վ�5=�?
�D?���>[Z�>	/k>�W�>���>G	>��<��=>��=y��=
�<6�b������<��L=W&����>\x0=.�ڽ+�c��%=qӄ>]G����=b��>a>���>	m�=������/>ʆ��Z�L����=�6��&B�i-d�9^~��/���6�ސB>OHW> R��6����?�vY>��?>Ȓ�?sIu? >���K�վzC���Md�mS��=�>�s=��h;���_�i�M�Ҿ�P�>6�>��>�P>�k'�0�7����=)=Ⱦ��;�6�>s��ZJ��r+��"}�{��G�����c��P�r-?!��9��=�fi?;N?>��?�T�>Q�9�	z��"�(>������>ȸ��![��X"�˳?��?�G?_����(��(̾�徽-��>�I�?�O�f���+�0��������C[�>~򪾷�о3�\k������F�B���r���>��O?�?�b��]���8O�����%���g?lg?�>�;?�N?������,�����=��n?���? 0�?1�
>Dn >@��}��>��?�0�?>�?7h?�o���$?�%?=q�=TU��7o>��9>���q�> �?��>��?߫��]ؾ�羷��D
N��t��=�>��>>�>�b�7�?ٽ����)�*>`W�>^��>[X�>(Ϣ>g��>�Y�� a�� ?H>��>1i-?���= "�]�����=���=_=:���C�c�սM۠�B�4��B��E�y����>ߎÿSQ�?,?�=��+�<�??1ӾSf�kO�>݄�=rw�'��>����
���?�f�><1��{%�>Ųw=��þ�%�=���E0/��?�K�C�JӾ�ߚ>����ʰV��c�0�=�%��m¾K���{�]��,�|�$�H�<��?ﲭ�B}��5�����&��>�f�>E�1?&�h������,>���>P��>����{��	��Ɩ�(�?�[�?�$f>��>.�V?O�?p,��%,�f	X��t��?�m6e���_�Tݍ��Ѐ�T����Ƚ�Ha?�y?	Q@?)��<|�x>]�?9�%����酈>�j.�Oq9��|E=c�>�譾�d���پ=�ž�����N><�p?pV�?��?�bS��!�<�+>�a*?n9?O�}?8�<?��@?�eY�w�9?;��>@�?ټ�>%R6?��?~�>8�=0�
>P1��G�D>�o��f�1'ν���z�<cb<=�،=8��<Φ�<.�0��qo��� =dɺ�tL8�"Ȑ�<!�=�=jW=��S=+̨>�Tf?�z?�y�>^n%?'
���Qa����B-?�p	=|�5� �����~X��`X>5F{?a��?��q?�8�> �Q���n�a�=�$�>|��=�	�>;<�>:�������"==�=�q�=��=ZA�<&C��!�Cz������Z!>b��>9N|>�Ǝ�̸&>����_;z�¥d>�P�u�����T���G���1��v����>[�K?:�?���=���(��Q;f��(?�:<?9hM?x�?y�=\A۾��9�(�J�n�c��>��<t������X$����:�%K2;8=t>�՞��Ɇ�Ϭ8>ɫ�?A侎i�"(@����oZ�=�I��#��;�	���ϾNύ�L�=�>Ne��%�� ��`ޭ�ԹK?�4=�د���1��þD#>�Ȝ>qz�>j���Ѷ�{<�H���/0=��>�+>���:���k�W��u	��7�>k�N?�f?�2�?�(��h}b��V�	�$�#�	�->h�?��>�)?�h^>F�D>�^�7�o�Z�t����>�O?��Ҿ�o+��l��(�6 C����>\�>�Z0>�"?��I?L��>�/U?�w ?b�?���>?V���ھ�<&?���?Pp�=D\Խ<�T� 9��$F����>=y)?�JB��>�?'�?��&?�uQ?��?5>�� �>@�ߌ�>&S�>\�W��]��`>�J?v��>a?Y?�҃?)�=> w5�6���v��X�=4�>��2?P3#?f�?���>#�?�����P�=�!�>��y?%��?��e?;�"=B;?`�N>���>�0��Mx>�8?���>��3?1\s?�,R?� �>�]��D�Z����w$�C-����=��<�
����X�����!&�=�h�<�#�<�m��z�=,ߞ<���@�1���K��K�>ѧs>G6��BZ0>z�ľ�S��E�@>���q1���튾�q:���=Rv�>�?���>�`#��ƒ=�>�3�>.��� (?�?�"?w@);�ob��ھ�L�%e�>-�A?F��=��l�H{����u��f=X�m?uq^?�W��[��N�b?��]?Oh��=��þq�b����h�O?@�
?B�G���>��~?[�q?>��>��e�#:n�&���Cb��j�nѶ=Or�>QX�D�d��?�>o�7?�N�>�b>l%�=nu۾�w��q��\?�?�?���?�**>��n�[4��q���N���
^?Qm�>�'���#?*����Ͼ&k���+����� ������=���o��_�$��ڃ��P׽���=�?Ys?�Zq?�_?)� �B�c��2^�����_V��%��E���D�ƅC���n�U�]_����!aF=p�`���F����?��?2�?�?��f��� �y�'>����{�)��
�=���b1�=oۨ�Y��WYd��'þ�?$!?�-�>�bf?H8z�B E�)cE��R�����S�> ��>SZ�>*�?ii<�^Y=8��>�����ޝ���4v>^yc?��K?�n?Dl�w+1�������!�!�/�Dc��h�B>�g>��>L�W����J7&�tV>�j�r����w����	�К~=��2?�)�>"��>ZP�?C?�y	��m��mqx���1�縃<m3�>�i?�<�>��>�н�� �f��>��l?��>��>F~���R!�G�{�,�ʽ9/�>���>ɦ�>��o>�y,��#\��k��X����
9����=a�h?�|��I�`�uօ>R?�Ҍ:��I<���>�Mv��!�����'��>�l?�Ǫ=h�;>Hhž"���{��0���R)?n:?O����{*�M�~>�>"?ɀ�>��>01�?C�>R�þ������?r�^?J?.FA?�w�>r =/;��IȽ�'��*=���>,�Z>"�o=x��=���|\�=< � fE=Hݹ=ȂѼ^췽x<�ǳ�	�F<a�<`�3>�[ۿdFK��ھ������ނ
�'3��'j��Yȅ�k���1���|��Z^y�_ ���R�T�Pc�g�����j��?"s�?�Е�����?��`��E����>��s�����ـ��X
������Q߾����{!��%O��g�U�d�W<C?BA��g�ƿ����ε��z?�N=?��_?C���,�ۼ�@\�;�j�8�6=xS���n��9/տ�=���HU?���>F`Ծ>&F�>k�>U��=���>rS��T��Z�>���>�w(?Rf?:�t��Ŀ'u���¼��"�?��@�aA?(�HR���]=�p�>7	?}�=>�12��T�����K'�>%S�?�=�?D1C={ X�	F�,�e?�sE<�F�t'̻[v�=i�= =�c�ŚL>E�>\��ҧ?�S@ܽ9E4>�݃>H�)����~f`���<3~\>ǵԽ6��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��=H)��@���(��*�k��;�m��)��$���E��p���@Ĭ��O�	
���=�E>�US>&%p>N�b>jI_>�1V?1a`?=ͬ><�=��;֍��;�����<� �����r�w��������ྑYǾ ?	�ɔ�9��vN��o
0�$�̽5m��-����z�F���2��]?���>x��5(��<>�ؾP�žg�^>.I���栾����9�@��m�?�$?�Ȃ���L��O�=4����?-��=%��]4��;#A��m��8�>���=���NL7��!^��u0?O\?W���J[���2*>6� �]�=��+?��?��[<�!�>=L%?k�*�=�U[>��3>hܣ>M��>�D	>��\b۽F�?��T?&���������>-^��]�z���`=�,>aL5� ���[>Z��<?팾�AV�S���Y�<q%W?A��>,�)�H��>8�������<=��x?��?�b�>qck?7�B?���<Wl��/�S�8���x=7�W?�(i?b�>'ǁ��о�����5?J�e?�O>�,h�?��~�.�zQ���?��n?j?�����W}�Z�����|d6?��v? s^�vs�����H�V�]=�>�[�>���>��9��k�>�>?�#��G������qY4�Þ?��@���?�;<�-��=�;?u\�>�O��>ƾ�z������E�q=�"�>�����ev����R,�X�8?ݠ�?}��>1���ʩ�so�=���q�?rJ�?x���D��=B_�M�w�|����D=���=�2��&�<�O�|�^�����C嬾�k��1�>@���L+?m-����Hѿm񅿈��¼��r?��>�/�*ɏ���M��:S��L�ɴG����L�>�>P��������z��:��X��t�>���l�>u�R�2 ��h��4��;���>�\�>a��>�L��F ���̙?�����Ϳ�������M Y?�˞?�x�?l= ?"2<)u��5���Q�%UF?K%r?�+Z?#�+�ـa��N��r?B=˾+"T�916�)Mf���>&ZI?�ě>l�N�=+� ���>�&�=y�G��ÿj�ÿ6���k�?ع�?�� ��K�>؏�?�72?����꥔���о��8���'j3?�>�,��RO1��Z��?�����>+�6?�}��g��]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?ֵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?Y$�>��?!o�=�a�>d�=O񰾉-��k#>B"�=��>��?��M?L�>]W�=��8��/�D[F��GR�_$�>�C�"�>��a?�L?{Kb>a��9 2��!��uͽ�c1�MP鼕W@�h�,���߽5(5>��=>�>W�D��Ӿ��?Ep�/�ؿj��cp'�h54?���>E�?����t�<���;_?5z�>7��+���%���B�h��?�G�?k�?r�׾�X̼d>8�>!J�>��Խ����������7>*�B?���D��q�o��>���?�@�ծ?|i�	?��.X��^y~�e���7�t��=�7?���W z>+��>���=Ev�0���e{s�y�>��?wu�?��>��l?�Yo�
C���5=�T�>Ԥk?FB?�������B>Ϯ?���o}S���e?F�
@&T@�$^?������ؿ��E����񺾏�>
}�=��>�P-���>�?�mI۽j8Խ�@s=��s>"�k>0�>���>)ۂ>fS>E�|�����𰿙]���ZF���'����E�l�d��",þB�$���&�G����=7.����hL�Tn���=�YV?�S?C�p?�M?��s�D� >[�����=/-��v�=`�>��6?��S?E�'?힨=�B��σb���~�@��������>Ƣe>���>R��>}��>>�����h>��F>��k>J>�W�<�
�L=x~F>�y�>]��>��>[�>�q��+#������x)p�����U��B��?��)�3c�ɵ��ԯ������<��?{5>HV���Ŀ����f!<?6��!�쾿��7��?�%x?\�z=��<�<hE,>vr���?�	�|>o�}� �M��_���q���??�?h>0�s>��3��h8���P�R򯾄�|>�6?M����v:��]u���H��޾@M>Z�>�:�K��� ����~��h�E�{=b�:?7N?�Ҵ��˰���r�/E��&�P>�a]>n�=ө=�ON>/�^�7�ɽ��H��&=X�="�a>�F?�p,>���=E��><H����O���>�@>��->�@?�x$?)[�	ޓ��O����.��v>QJ�>m��>bW>�KI����==�>�w`>������9��?�҉W>x|��`��Rz��Ws=����ʐ�=F��=� �#�;�<�(=%�~?���(䈿���e���lD?j+?] �=�F<��"�A ���H��=�?k�@m�?��	��V�1�?�@�?(��/��=B}�>�֫>�ξG�L��?5�Ž'Ǣ���	��)#�jS�?��?�/�Yʋ�Tl��6>_%?հӾgf�>Oz�Z������u�ݦ#=u��>f:H?qU��5�O��>��w
?@?#_�_����ȿ�zv����>T�?���?��m�sA��@�ʁ�>ݢ�?fY?ji>�b۾#\Z���>H�@?BR?;�>/:�g�'���?�ݶ?z��?�I>	��?��s?�j�>��w�aW/�3��ǔ��	i=�b;�e�>�L>P����eF��ؓ�	h���j������a>l�$=��>&H�:���6�=�싽�E����f����>H4q>��I>{R�>�� ?�\�>��>_�=�W��oـ�����}�K?���?���2n��M�<��=h�^��&?oI4?h[�\�Ͼ�ը>�\?h?�[?d�>=��O>��K迿1~�����<��K>4�>�H�>\%��tFK>��Ծ�4D�Up�>З>����?ھ�,���U��OB�>�e!?���>�Ү=Z� ?�#?}�j>o1�>.VE�#7����E�e��>��>#U?��~?-?M����[3���桿��[��dN>��x?�S?�ɕ>ی��f����qD���H�����?\qg?-2彫?�+�?�??��A?H�e>%���ؾ�����>��!?�����A��R&����w}? C?���>z:��uؽ�Bռ���������?��[?�6&?���:a�`þ���<۟#�VV9�
#�;V�Q� �>;>�0���g�=��>�:�=�m�4�5��]t<�N�=�D�>�`�=��7��Ċ�0=,?��G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>$�l���K���ڙ���F��_�Ž�d��J?��X>���>�'?�uI>���>0�\��T-�Ỿ�ʁ�E%��]��(���]���!�����޾�n>�������ZKa>C��T��>��>*D@>{�>ɜ:>}�>ٗ�>I�P>D�>1��>�o�=�|�>֑>8ǁ=����KR?����B�'�ķ辷���A3B?�qd?�1�>_i�2��������?~��?#s�?,=v>�~h��,+��n?K>�>���+q
?�P:=!-�1;�<�U��\���4���쪎>�D׽� :��M�0nf�Fj
?�/?��/�̾�=׽!�����n=�M�?��(?	�)���Q���o�˸W�S����l6h�]j��N�$���p��쏿�^��%����(�4s*=��*?e�?Ό����!���&k��?�hdf>O�>e$�>2�>2uI>��	�p�1�c^�M'�?���mR�>x[{?�9>�)P?o�T?�5d?.F?�!>J�t>-�~���>�����ۢ>�|�>W b?Fbl?��?J�%?�D?�U>[ۊ�J���P������>��3?�?De?��"?�g����J>�M=U(������D� ���5=�0��Lf8�#8�<4)8>��$>+P?�u�Ǩ8�����4k>�7?���>f��>`���!�����<���>F�
?�F�>] ��zr��^��9�>ա�?	�\;=�)>���=%��� ݺwT�==<ü ��=����:�8!<���=���=�;u�E�E����:^��;&]�<u�>8�?,��>�D�>�?��3� �h���b�=�Y>�S>4>"DپQ}���$��N�g��[y>�w�?�z�?v�f=V�=��=}���V��)��f���\��<>�?J#?>XT?3��?�=?Mj#?�>�+�XM���^�������?��@?#">������$���n)�; 9?���>">D��-
��}<�@"����q�/h�=��<����:鴿��8�%��=�]�x������?9��?���n@��ھ�����-=?�.>f��>�+�>Q�ekc��@J�G~>��?��K?{�>��?_��?��T?2��=!�m�$W��R�j�����2��>4�?�El?Tp?^DT?�g�>���>p�= 1�@6��둽8���>�0���B�!Z�>ؾ >y"�>��>yq�>Jp��@x���.��=r8|>Z��>�أ>L�?���>�8�>��G?���>�X����-夾���=���u?���?��+?4=~�A�E��F��&D�>	m�?���?�6*?
�S����=��ּI䶾��q�I%�>j߹>~3�>'Г=��F=�V>�
�>���> 3��]�p8��4M���?�F?���=j���*�i�Hf������&�� ����Uc�afW>��	�ʽÜ���:��ɯ�ADj�6��m��QQ���߽��/�??ϖ�=��=���=8��;��)��0<��F=���ny=^��;W��=�99<|Z>����'�d�z��<��%>�'����˾�}?�H?y5+?��C?VKy>�8>"�3�Ǖ>耽%z?opR>|�Q�rE��lF>�����4��A�پ&\־@�c�9*���>�NK��>" 2>�%�=��l<�p�=W�x=�=hO�S�=���=��=�o�=j�=�>&�>�6w?6��������4Q��[�е:?�5�>���=|ƾS@?��>>�1��I���c��,?��?`S�?��?�i�"g�>^����|�=����o@2>���=��2����>��J>G��"K��򍳽�3�?��@`�??Y⋿��ϿRV/>d�)>���=]cT���6���c�>�p��[�K(?�28��RҾ\�>��=�yھ��ƾ9�w=2$>$d[=�Mܽ�U��$�=]����<��y=��>��S>U��=A�½�k�=�mm=��>��H>#�⻑�}�;Np�w�G=���=��^>΅>�|�>�	?e�;?Lf�?���>�ې�0ֻ���.�>�p�>�=��>7��>��>�?ǥ?�dj?QZ?Q�.>��>�I�> "�@v�CN������|���<g?+NY?H+?Ζ�:6� ����5�[�㱍��o>�?�=&?��>*����ӿB�'�ڄE���`�;׬=d׼�l�= �Z�J�����ed<aw>~s?���>s�9>��@>f�U>���>�.�=k�=��=��üJ����,��q�=^]Y�F	�=��#��@=ёn=�{����ý��`�5g��a)|=l�}��2�=h�>��
>���>Ȣ=є��S�=>𙗾'NL��t�=C����G�-1i�-π��o0�#�S��">��2>�L��g���
?��<>��<>�o�?��u?��>����g�Ծy��4�3��ʅ�$��=A+;>"�8�M�)��DV�)sS�'�ϾAY�>JvM>���>�A>i4�~�5���9>�	�8�-��S�>@J��´���s���l������d���gq��ڴ�x�G?l'��*$�>.J?YGQ?ѡ�?I�>��I�M�H�.죻�3���ڋ>6@L������j=��?O�H?a�?Р���;��H̾���iط>=LI�I�O�"�-�0����̷�D��>)���G�о�"3�g��������B�Kr�u��>�O?��?8b��W���RO�C����p?�yg?��>�J?A?�%��
y��t���i�=��n?J��?�;�?��
>�%/>޼]r�>Q[	?,�?�I�?x�N?u�B�![	?��`>7��<��0$>f>��\���=v $?H+?:.?����u��d�#��X>��w>YF�>:g>�#7�SR�=ZO ��M���>���>a*�>
�>:Ej>=)b>�������?���;�,�>Ѵ:?��>�	Ҽ9��5�<x��=������Q5��O���S�����;~��J�?=h��>�ƿ�9�?��>���_e8?��Ҿ?���>��=�ⒾI��>a�)>�!S>lM?~Vx>� �=��>�=��{PӾ�>���Ҋ!�)C���R�J�Ѿ@�{>*���3�&�z��Sa���YI�wB������i�"��^�<�w�<E�?������k��)������f?S�>��5?>F��������>,��>��>c���������J�?E��?�;c>��>G�W?�?��1�3��uZ�$�u�V(A�e�U�`��፿����
����%�_?�x?:yA?"T�<.:z>G��?��%�Yӏ��)�>�/�';�$@<=m+�>@*��4�`���Ӿ��þ�7�IF>��o?3%�?mY?8TV���2��)>��8?�s1?�u?|g7?�>:?l�v&?A=>��?UT?�2?^�0?�t?�8>q�>���;o�W=�)��>A���kǽ��ѽ���*�<�\Y=}��~{"<��X=a��<G6�|����;�����@�<Fp;=k+�=eP�=���>��Y?OS ?:z�>3<?�v���7����R�4?��]>��������)�����&�#=_�J?M��?٥i?�#�>�� �X�7����=��>w�:>�T�>.�>C�+�{U��6�=�|�=*D=���<X������h���Q���}2=�='>��>Y0|>���C�'>�|���0z�S�d>��Q�r̺���S���G���1���v��Y�>8�K?��?K��=>_龜,��bIf�60)?�]<?�NM?��?��=��۾��9���J�>���>MY�<���	����#����:�V?�:��s>
2��kR�<C	>� Q�����C���J�]GϾ��n>�t��[�U��˾+bþ��$�����6<����[��(u��~���*,?&��o<B꽥�	�m�=�?��>^��m�A>�U����3	��� ?I�>o�_����X�^�I�.���>>�R?T�p?��?�Ȣ�V��ِV�{��������=/l2?�߽>��?q�">ۮ�=����7�C�b�x�V���>g�?����A���y� �� 7��լ>/6�>UpB>N�?K�C?���>�)o?�P?�y?�;�>s6a�ˉ��?&?���?	�=D�Խr�T�D9��F���>�})?�B�q��>ڈ?E�?��&?�~Q?Ϯ?c�>[� �i:@���>O�>��W��^��	`>;�J?���>�0Y?YЃ?��=>ǃ5�4梾�穽Č�=�>m�2?�5#?+�?��>� ?�v*�G3�=�ױ>[4r?>�k?W?�X�=��?�_�=�ǚ>�!v�+ �>j�?a}�>�6X?�d?�(?S-?��<(��9k�����u����8��߻u�=�ɽ���B�cC0==;=>�=���=�Z(���Z;� `= Gr�zT�>/�s> ����1>�þ����A>*��W���1`��n0:�kJ�=���>�?�|�>�T"���=~��>�m�>�����'?D�?&�?��:�db�;�ھ��K��;�> �A?���=�m��w����u� �i=�n?�v^?{W������a?��^?�G��9��	ž��i����P?��?��(�B��>O�{?�vq?�\�>	�j��cn�؀��Q�]�+�Z�A	�=F��>A��d�8�>6?6��><JU>�}�=�c侍�v�-��A�?�P�?7��?�Պ?&�->��l�uݿ3r���L���^?
��>>���#?g�����Ͼ.@���(��H
�V
���%���S���u����$�\ۃ���ֽ���=��?�s?\q?��_?�� �y�c�!^����jV��$�� ��E�gE���C���n�\X��,��b��ZG=�D��YO��K�?P�?��d�{Q0?[xZ�& �ȸ���9>�Z��S�Y ��v�X��<ʗ�<7�a����Z<ȾZp?���>_�>��N?���  *��
���W��R��1Q>��>7r�>�	?�����	ý�MR��8վ��k��]���v>�cc?3rK?>�n?�i ��x0�����#!��h�yԥ���B>Q	>���>�BT�=��6�&�bl=�/-r���� W��� 
�5w=C2?�a�>�ל>
%�?��?/Z	��毾B�{�P�1�\y�<��>��h?"r�>,6�>Hӽeb �Wj�>	On?@�>t�>2��+�!�*:o�����>���>�r?��l>��v�U��p��uȎ��q6��o�=�"h?�ہ��i�&t_>�C?Pۣ<*gK<�י>�\���	$�6����O1�y��=y�?բ�=��E>"C��\���v��\b(?~�?ꑾ�c)�^i~>�� ?��>s[�>M��?���>CľE��^?�^?�*I?D@?�D�>j�=�잽m+Ƚ�N*���3=��>�_\>O ~=`]�=���qZ\��w�`D=�6�=�տ�V�����<�r��_��<���<Xi2>x�׿�I��{�$��X4Ӿ<���򈾿w��Ȑ���2�[�Ͼ#��d������)�n�g�v�O�!ej���C�X��?���?赭�(t��[đ���t�	��g
?�?1��b�BϾb���������`������_q�m�}��Lp�B�'?���˶ǿ
���1Aܾ� ?�- ?��y?����"���8�^!>Ȭ�<�H�����u����ο��^?���>����N�����>0��>�tX>�q>D��̞�" �<��?�~-?���>��r�ŕɿc�����<���?��@??��%��>��U=H��>џ	?XF>�-����#���d�>}��?��?JC=`@[�L�=�X/f?��;�iF���>Q�=N �=�G=��'�>>�>��.�(`<�^���	:>p��>�mϼp� ��%b��N<�T>t`ǽr��5Մ?+{\��f���/��T��U>��T?�*�>X:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?&�(?8ۿ��ؚ>��ܾ��M?_D6?���>�d&��t���=j6�����{���&V�~��=\��>d�>��,������O��I��T��=� �G�ſ��#�ڳ'�Q�<=�Z/�W ��Z��������b��zγ�ր�&�>��>C�>,��>>��>V��>�T?d	v?(�>3&>�B��y���#��6�=HCY�gZ�f����pn�������
��U���O)#��k"�n�ᾥ�����=�*���n��6o��Q�ܡH�{�l?S U>�8���E���Y>r��f����oU7��9 ��d��q�<�+ڣ?N<?`F��C��9�����~���`��1P?;]��[��`*��>��+�@$����4>Z�<�H�����l�_,?P�?gϿ��@���{@>�M�JZ=Fr(?a/�>D��<=�>!{"?���*�Խ��0>!>�٭>���>�Q�=󸮾�,�08?��S?��ؽ@��u�v>�j̾��t�_W�=|v>�5�B�39Q�v>9j�;�u��������o�[�=��V?ɐ�>|�(�������E*�aH=аx?�)?��>�:k?**B?R�<13��r�S�w���Do=EW?�i?&[>����ʜѾ�Ȩ���5?�d?,qL>��i��{뾕�/��Z�k�?��m?+?I���{��3������p5?��v?s^�xs�����M�V�h=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�$Þ?��@���?>�;<��T��=�;?m\�>�O��>ƾ�z������'�q=�"�>���~ev����R,�f�8?ݠ�?���>������Jj&>><B�mE�?�?�?�"�Տ>e�
��"���v��>^�8>?��=]0�=U����w׫���%�JZyP� 7z>��@�}(=�??[�3�y0����ܿ
�^�H�&��=/?N	y>���=��ͽ�9I���V��x?��ij��|���[�>��>IP��6����{��o;����i(�>��q�>��S����V���3<�ے>���>���>}��!���Ϳ�?ZV��<2οH���M���X?�c�?�i�?:f?+�:<�w���{�3m��0G?�s?�Z? �%��M]��[8��j?w_��oU`�َ4�CHE��U>�"3?�B�>d�-�G�|=#>x��>eg>�#/��Ŀ�ٶ�����F��?ˉ�?�o����>s��?xs+?�i�8���[����*�+��<A?�2>���,�!�0=�MҒ���
?(~0?
{�O.�\�_?)�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?h�?ص�� #�f6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�i	>���?�~�?Qj?���������U>	�}?�:�>�?;��=�.�>��=����7�!�W�#>���=��7�ޥ?�YM?o��>pr�=i�9��,/��F��R�p���C��U�>{va?�!L?�5c>����,Q4��:!���Ͻ��2�����A��r+��wܽ��5>�>>�h>�E�КҾ�k ?!o�xiٿ�ؗ�g�'���-?=�o>��?�����Έ�2���_?�}>̆��ᴿz������f�?t2�?m)?P�Ҿ�bk�#f/>3u�>��>I+ӽ����~����+>m�F?X�&�L���ZBp��>೽?��@$d�?�_r��	?`��W��Ic~��� 7�_�=��7?��9vz>V��>s�=.qv�������s�8��>�0�?�v�?���>'�l?[xo���B�MW3=�4�>ޏk?�n?�8x���a�B>��?j��9���N��f?'�
@vm@��^?������ֿzZ����ž+���B�=@6@��$�=e���9��=�!�=8!�3������ݠ>8��>?��>Ec�>�=�=H��>�d��u�#�7x����ʩQ�4w"�9���X��}�	�`���i���Ӿ��о/��bD�=���=T"B���!��f����=�U?MR?��p?�� ?rp�>` >'^���=
��x^�=��>�x2?շL?��*?���=�T��^hd�
倿�Ŧ����h��>hI>f��>���>�`�>�����F>�3>>��z>���=�)=�E޺N=��Q>��>�d�>N �>�W8>��>%,��-l��]�h�7}����뽃ϥ?�M��ƜN�����P��ᴾ�N�=T1?�@�=;���mQͿr~���2F?�p��b8�i�.�SR�=�.?�oT?,�>����MZ�)�>+sؽ>f��>���H�e�d.$���C>��?��d>p�]>��?�]JP��^���оMC>��j?M�u����#�v�������>) �>�����4��|����u��KH�����[�X?���>��ܽ�Y�h����L�T��=��>Af<84k>р>L.��dU��M��8�=}�2�N�>>O�>5�J>o�p=b�>��J��>���>�O*>�k�=W�>?�R+?�.��<t�9��Z��ߠ�=���>qM>w�>v�G�/S�<AR�>.i>��<�s���(q�dF����L>2�_���R�wg�*�=��;D�>'��=��1�c�5��A�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾFj�>k9��f��]6��ܗu�$y =2п>�nH?�n��\�W�d�>�?%?
��4�����ȿ��v�~��>Ӳ�?��?7m��m����?�|`�>�;�? �X?�gi>E!۾l][��-�>��??�^Q?P�>ڞ��(��y?���?L�?�tI>��?ʄs?�d�>.Zz��[/������Y����=���;&��>To>�<��YGF��ѓ��w��ڕj���CJb>��$=�ظ>-��b���]T�=����Y��d�t�>��p>��I>���>�� ?���>���>ɓ=�i��2܀�������K?(��?��� 8n����<�g�=M�^�S6?�J4?ץ^���Ͼ�ߨ>W�\?��?R
[?j]�>
��<;���࿿�w���ȕ<��K>[7�>�C�>����`UK>�վ�/D�p�>�Η>�Ţ�@@ھ�,��˦�>�>[g!?q��>��=%u ?=�/?�[�>u��>bE�x����� ����>`9?"4>?�+y?�?>0��ө/�u�������J��R>Ow?�U?���>�������Lt����5Xѽ��?czW?d􀽚�?��e?�*3?��6?��>gUG������㶽
#|>��!?����A�R&�����U?�?�5�>�W����׽D�A��d���?�\?�5&?�t���`��¾�/�<�)(��D��;u�E�x�>��>�������=Da>�.�=Hm�{6��lf<��=ܪ�>G��=T7��6��/=,?��G�ۃ���=��r�<xD���>�IL>����^?bl=��{�����x��)	U�� �? ��?Xk�?i��?�h��$=?�?T	?n"�>�J���}޾:�ྻPw�	~x��w�Z�>���>i�l���K���ٙ���F��S�Ž>��#�>���>���>�?�E�>-��>�j.���E�����g����G��F��A��T��1"�{)��U��Bx�D]ھJ@���d>I��=�L	?/�	?p��=x�>{;�>y��=�(�>d��>� �>���>���=+u�=�ۢ>�2H>VA�=�JR?����h�'���辙����1B?]pd?�/�>oi��������N~?��?�r�?�2v>o}h�*+��l?c>�>����n
?�\:=9�5V�<�R��\��xI��k&�9��>�L׽�!:�M��gf�}i
?a0?�⍼ӊ̾�3׽����uNo=�L�?��(?y�)�E�Q�g�o� �W�)S�c��h�d_����$���p�^쏿x^��� ��(�(�Lb*=��*?��?����#���)k��?�.}f>��>0�>��>hI>��	��1�� ^�4N'�vǃ�MH�>'W{?k�>�;?ϖ>?�ka?Sh.?M��>8�>p��{Z?�`N>ky�>���>��??U�(?�	?��>W%? �1>��=<!ھ�7�t�>w'?��(? T�>ue5?�l����=[#�=�+��E)�'?�0��=���=�q��-5���"E�=g?g���8�(^���-n>�7?F��>���> ҏ��O��
$�<_M�>b?jƏ>�� ��!r��j�#c�>�^�?do�r0=	*+>q6�=y���$�H^�=B�Ҽ���=@��D�<���<h �=I�=�W���$:[;`S�;Kt�<��>"�!?$;�>�?�>������辀���sd�=�l>
��>��>����4���)���.(a�=�M>f�?���?'��=�j>�g>k���W�v���׾`�;<S�?�r%?Ue_?o�?.4?�C?vޣ= �"�>���(������?��;?�Y�>�J��8��Aƺ�&9���-?��?�6���<�k�P��Mھr¾Ը#�k�!�Ro�`پ�AP��	̾x�2���r=��?O�?��[>�A������n��5���-J?�F�>k=�>�u(?�oK��rZ�Lx��j�>u�>n�g?7�>�`�?7�?STq?��M>5E��͌ƿ.s���L��(�>�/{?�6�?.F?��E?Q��>���>�o�<A����Ͼ��b�Rt�� ��b��=�J�>�S�>?z>�su=D��>�U��,?��Hͽ��=��=sܸ>}��>'-?o �>ڄ�>v�G?��>�X�� ���⤾ۻ����<�_�u?��?ȋ+?9=W����E�>=���D�>�p�?W��?�1*?��S�8��=�ּ嶾�q�� �>չ>72�>�ד=�F=�j>w�>���>%��\��g8�#M��?IF?d��=Z���xn�ߌz�mo��&�����.�h�%^P�^�M��Q�=Oq��A�ý�$���g�
�����.�����cz��� ?jd=lY�=��=�۽<m��M��<��/=UJ�<:~=6s�e�6=n��� ��H;��g0���;�И=�浹��ʾ�T}?9I?��+?��C?�/z>{.>>�3��C�>1���R)?7@U>~L��g��J�<��C������ؾ�־��c�m����n>��J�r<>>3>'��=Č<=K�=<o=wЌ=u�=���=ڕ�=}�=���=���=|[>��>�6w?U���	����4Q�zZ罥�:?�8�>b{�=��ƾk@?v�>>�2������tb��-?���?�T�?=�?*ti��d�>I���㎽�q�=N����=2>|��=j�2�^��>��J>���K��A����4�?��@��??�ዿ̢Ͽ7a/>���=�N�=��K��@9�8v�U�F�.yl��.?zn��aھ׭�=�q{>�dľ�R̾ S�=P�	>��:EV,���H���=N
��
|<��y="(m>.�X>���=Jw.�:�z=q��=y�Q>Y1�>N
�<��ͽuJ��G	<Fܴ=.�>c5>���>��?��8?�p?o2�>�ؽ�҉��"۾^a�>�:*>�[>c+�=�:n>Q�>��0?��>?��R?�î>�7�=���>��>��1��2���[��a�����<ӽ�??8f?�"�>��+>@E����a>F���`�FF?#?�q�>��>�����X#��B���D�="�����=�i>��N�`�L���7���վ�5=�?
�D?���>[Z�>	/k>�W�>���>G	>��<��=>��=y��=
�<6�b������<��L=W&����>\x0=.�ڽ+�c��%=qӄ>]G����=b��>a>���>	m�=������/>ʆ��Z�L����=�6��&B�i-d�9^~��/���6�ސB>OHW> R��6����?�vY>��?>Ȓ�?sIu? >���K�վzC���Md�mS��=�>�s=��h;���_�i�M�Ҿ�P�>6�>��>�P>�k'�0�7����=)=Ⱦ��;�6�>s��ZJ��r+��"}�{��G�����c��P�r-?!��9��=�fi?;N?>��?�T�>Q�9�	z��"�(>������>ȸ��![��X"�˳?��?�G?_����(��(̾�徽-��>�I�?�O�f���+�0��������C[�>~򪾷�о3�\k������F�B���r���>��O?�?�b��]���8O�����%���g?lg?�>�;?�N?������,�����=��n?���? 0�?1�
>Dn >@��}��>��?�0�?>�?7h?�o���$?�%?=q�=TU��7o>��9>���q�> �?��>��?߫��]ؾ�羷��D
N��t��=�>��>>�>�b�7�?ٽ����)�*>`W�>^��>[X�>(Ϣ>g��>�Y�� a�� ?H>��>1i-?���= "�]�����=���=_=:���C�c�սM۠�B�4��B��E�y����>ߎÿSQ�?,?�=��+�<�??1ӾSf�kO�>݄�=rw�'��>����
���?�f�><1��{%�>Ųw=��þ�%�=���E0/��?�K�C�JӾ�ߚ>����ʰV��c�0�=�%��m¾K���{�]��,�|�$�H�<��?ﲭ�B}��5�����&��>�f�>E�1?&�h������,>���>P��>����{��	��Ɩ�(�?�[�?�$f>��>.�V?O�?p,��%,�f	X��t��?�m6e���_�Tݍ��Ѐ�T����Ƚ�Ha?�y?	Q@?)��<|�x>]�?9�%����酈>�j.�Oq9��|E=c�>�譾�d���پ=�ž�����N><�p?pV�?��?�bS��!�<�+>�a*?n9?O�}?8�<?��@?�eY�w�9?;��>@�?ټ�>%R6?��?~�>8�=0�
>P1��G�D>�o��f�1'ν���z�<cb<=�،=8��<Φ�<.�0��qo��� =dɺ�tL8�"Ȑ�<!�=�=jW=��S=+̨>�Tf?�z?�y�>^n%?'
���Qa����B-?�p	=|�5� �����~X��`X>5F{?a��?��q?�8�> �Q���n�a�=�$�>|��=�	�>;<�>:�������"==�=�q�=��=ZA�<&C��!�Cz������Z!>b��>9N|>�Ǝ�̸&>����_;z�¥d>�P�u�����T���G���1��v����>[�K?:�?���=���(��Q;f��(?�:<?9hM?x�?y�=\A۾��9�(�J�n�c��>��<t������X$����:�%K2;8=t>�՞�N��p�a>��'g޾1[n��J���GM=�P���S=@���վ�c�|Y�=�
>����� ����uЪ��0J?��l=O���V�	x���r>h��>���>&�<�`�w��b@������,�=m�>V�:>,����)��lG�-&�]��>!SP?ڌd?Vہ?@֤��'n���X���Gn��-S=��"?���>~�>�>%>m<�=OǕ�A��u���L�QX�>OM�>D���6B������D��u&�J�>0W?^��=��>H�D?l?)�K?l�+?�	?���>i�=����:&?)��?��='Խ[U��8�V.F���>G�)?$�A�9'�>qV?^�?g�&?�|Q?t�?�S>I� ��g@�u��>��>d�W��K��=�^>QJ?$��>�IY?��?�%>>�O5�����7���E�=DU>e�2?�~#??�?M��>�?����Ã>x�L?hL}?h\�?�t?ջ>z(?^��>�)-?6�f���>�.�>,�)?� P?`��?D�?@��>)�f����R:�I@�=P��>�x,>Vd#>�O;H���jI3����j��=:eh=��->��W<�b�<�Y=sѩ�J5��_�>|�s>�	��P�0>a�ľ�O��i�@>�����O��dي�׍:��ݷ=H��>��?.��>�W#�¹�=Q��>�H�>���6(?��?�?��!;��b���ھL�K���>	B?���=��l�������u���g=��m?̌^?��W�;&��L�b?�]?*h��=��þ��b�Չ�]�O?<�
?0�G���>��~?b�q?H��>��e�":n�'��Db��j� Ѷ=Rr�>IX�R�d��?�>m�7?�N�>6�b>%�=fu۾�w��q��e?��?�?���?+*>z�n�T4࿬���u���t^?�~�>Vg����$?��;��ξ�χ��a����߾�{���띾6���$���������y��M(�=H�?+eu?sul?m�c?o��X�c�y�\�����nkV�c��Z�hD�bE���D�`Vp�����e��/���!H=�Tp��lR����?1�?�c��?�g��M�G���wZ>E����ӽ��Y>1��;�~�=��=c�<�� ��0ؙ�è?�~�>���>A]U?B�]�=�9���%�*�@�����!�=?�>T>�>�8�>�=y��v�~���hʾ��|�d캽(z�>�*k?X$O?�P?���<8������K��z>�A|��8(@>��(>9ތ>�%K�)�<�v���+��փ��9%�b�����a��<��&?��>x��>F�?o��>��%��/��9���a:�� ��ϰ�>�ZZ?=��>TI�>�n�;֓�=��>G�l?���>K�>d���4X!�u�{�i�ʽ��>��>µ�>��o>��,�%#\��j�������9�:k�=��h?������`�q��>,R?�=�:�`H<|�>��v���!�����'���>p}?W��=a�;>ž!��{�7���`#?�
�>�o��W+�U`>��'?���>��>nL�?�֩>A���L�<~�?��a?��G?Y-A?�6�>��=X᜽0����	�B�8<�K�>۲+>��=
u>�77��zC��6�w��=	8�=����i�ѽ�]�;Y��/�<�dp=��/>D|ڿ-IK�o�ܾ�������ʢ���Ҭ�d���������෕��Y|�W�����/�R�:�h�N�����t��6�?���? �����͙��E�6=���y�>�z����@O���b�@,�����7m��z�"��DQ�:�g�J�c��?Y���6Dƿ�w�������>--?�?ݲ7���_�������>0I���5��I��r���ѿ[�张|?4W?I�ƾ��{�t�>l��=�˃>��>�t�E�}���ؽ�E�>)�>?�;'?(*�>Կg���2����y�?��@vQA?�))���neS=�I�>p�	?�7@>�1��	�u��'1�>,�?��?��Q=��W��D�8fe?��<#�F�Hܻ��=���=�=���sJ>���>�O�p�@�lݽ8%5>)��>}!�� ��
_�
"�<�]>��ԽP��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6��{���&V�}��=[��>c�>,������O��I��U��=����FĿI 7�v���<">ykҽ��Խ,{��b'�=�!ڽ`�Ծ���,\���=��>�Ou>)8>�;>G�9>� \?x.S?� �>��>1r��⨾�d�>��9i��~�3۾У#��?���+!�Wv��$��D>���-���<��v$=3(S�R������uj�'6���+?T2>�u�nX��l=GQѾ`���u+�f䖽�׾c�3�Z�p�=��?�gG?�y���c���@�2�ٽ��\?��T��g��Z|��K�=*}����<�>�p������L�)�^�:�Qz0?�L?�,���%��/�)>�� ��*=��+?�?�f<�T�> %?��*��K彧�[>�4>��>���>�u	>B
��;�۽f\?z|T?�(�&����̐>s��S{��M_=0>5�D�!�[>Y�<�����b��֐��L�<�*W?ƍ>��(�A\�v�������A=[nx?��?ط�>Uk?��A?���<�l����R�L
�ֵ�=^�W?o�h?->� ����Ͼ�Ǧ�l�5?S�e?�uN>/Kj�?���.�x9��?So?�?{Z��+}�RF����d�6?��v?s^�xs�����N�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?i�;<��U��=�;?l\�>��O��>ƾ�z������3�q=�"�>���ev����R,�f�8?ݠ�?���>������M�=hX��0�?:c�?YG��U=�J
�^�~�	���R�=�[K>�=��&=t�޾�*/�+G��'[�5�I��*Q���|>��@ݤý��?��s���￹8��ڄ��Z�y ��3?N�g>͘ھ*f���^��+q�[�T������ξ�M�>��>����e���A�{��q;�g$����>��	�>�S��&��ݚ����5<��>��>g��>+���罾4ř?�c���?οS�����X�X?/h�?�n�?q?�9<z�v��{����(.G?��s?ZZ?�o%��=]���7�t�i?��<�
Lw�W�E�kZ���;�BT?ˍ?|N,��(Ⱦ���>?t�O>��G����FzͿ$�?�#�?F�?w�ɾ+��>��?��?ՁP�F��ΣǾL����=�oQ?����X��4侄K�Q�U�J}?��?yO���l �]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�$�>F�?�v�=}a�>.Z�=�󰾈�-�Dh#>$�=��>�ޠ?��M?�K�>�R�=��8�}/��ZF�8IR� %�o�C���>f�a?/�L?�Mb>!��U!2��!��tͽd1�'V��W@�D�,��߽_+5>��=>/>��D��
Ӿ"�?@i�%�ؿ�i��{o'��+4??ʃ>�?�����t�;|��D_?ps�>�4�"/���*��zm�X��?I�?��?#�׾ ̼B(>�٭>&H�>4�Խr%��t����7>	�B?k%��9����o���>���?P�@dЮ?�h��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*��ٿ�Ԣ��������b>�s=�7>���ю>�YF���S��0��@>2��>�w�>��>&x�>��h>��C>y��n=�s�7����"���� ����z���*�{��������"���t�;j�T�'@��#}�!v�R�ֽH� >��N?}U[?3#c?��?A��<��A<�x��z:�L:ҽw*�=>	>��
?��J?�2?��=x�M���h�q̊��Ņ�*����+�>�5�>�s�>��?�i�>���a$#>+�>�k�>���<Nŵ=Ċ`>�Ƚ��:>Ӑ�>7+�>%��>��3>M�>���������d�O遾�hǽ�{�?�>���K��k��I鈾����KZ�=��,?�c�=Wّ��IϿs[����H?�N��Gr���A���=~/?�WS?�y+>O�����Y�R*%>��	�3'��a4�=ON�M�����,��}S>e&?��f>�u>E�3�e8���P�?����j|>�26?F嶾?N9�h�u���H��cݾ�@M>Qľ>��C�<l����O��li�9�{=dw:?I�?�D���ⰾ�u��<���CR>6\>w{=ad�=�IM>�gc���ƽ�H�TD.=ն�=)�^>iF	?L�0>~[�=��>�ꝾT�/�%��>�DV>�[�>�G?�e)?i)�����-g��C��%	�>��>qq�>�>��E�A
Z=���>�m>/��<��} ��Z�Tk>����-W�;if�s��=����1w�=R?7=�@C�7�O����=�~?���%䈿��!e���lD?S+?^ �=d�F<��"�C ���H��H�?q�@m�?��	�ݢV�B�?�@�?��Z��=}�>׫>�ξ�L��?��Ž4Ǣ�ʔ	�')#�hS�?��?��/�Zʋ�;l�6>�^%?��Ӿ'D�>��!����7�s���	=�>�^J?�(��W����>�G?W,?�m�6j���ʿ0�w�,]�>Ä�?�^�?��l�n(��*Q;��.�>r�?�?Z?�?_>�a־�OY�W��>�>??M�T?�C�>ݍ��;'�7(?��?���?�Nc>J�?U�x?��>Mw��E�Q�'����#��y~S=��d=�h�>22_>�J����Q��vr�e�]�J V��&N�U�<�Co=E��>J�̽�پ���=� ��9ξwA=3a�>�Z�=���<� �>�h?0��>;��>�*�=�ᙽt
������K?$��?Ƒ���m��<�=� `��?}4?Zs\�@�Ͼ�Ψ>f�\?@��?Z[?dk�>����H��q῿zg�����<}fK><9�>b��>�g��%M>J�Ծ��E�{e�>���>J���jھ�ρ�wm��>�>��!?���>�ޭ=ٙ ?��#?��j>�(�>EaE��9��Z�E����>Ϣ�>�H?�~?��?�Թ��Z3�����桿��[�b;N>��x?V?zʕ>_����&lE��BI�e���\��?�tg?qS�.?:2�?�??\�A?)f>և�)ؾ������>��!?�"���A��L&���?!P?���>:4����ս#ּ���z����?o(\?JA&?���F)a���¾�5�<��"���U����;�oD���>7�>Г��u��=>h�=�Mm�QA6�A�f<�n�=��>��=&)7�*����G,?D�?��F�����=a�r�'ND��>�L>ɞ����^?9<���{����L|��/AT�)��?���?3a�?I鴽�ah���<?���?C�?�^�>嗮�);޾0��8�w�,x��y�0�>�1�>��t�~��>z�������7��k9½C(1�TY�>�rk>1q�>c*�>_e�>喚>o����fK��������=�����ɛ2��dF�������J���=�oǾ>&���&�>ֺ��߄�>d�*?&Ɂ>�ǳ>��>�ڜ�\��=�'�>v/�>u�>�.*>���=|��>(�=њ���KR?������'����#���M3B?�qd?Y1�>!i��������Հ?���?/s�?�:v>�~h��,+� o?`?�>���q
?�U:=>�{&�<�U������6�������>�C׽V :��M�aof��i
?m/?F���̾{;׽�w��gp=�L�?/ )?��)���Q�E�o���W�S�K�G�g�U����$�9�p��揿�V�������(�5�)=�*?�!�?Kx���4���>k�V5?��af>�	�>!�>�վ>�aI>+�	�Ƿ1���]�I:'�����o��>�+{?�>;*H?�<?��O?�J?ꔐ>�W�>�ԭ�)~�>��\<_Ϣ>��>s{7?}6+?�_0?�|?Lt+?I]^>>���n&���hپ�;?�i?ȹ?��?R?I����۽��ļ�h#���y�r��g��=�l�<ȷٽ�%{���R=IP>��?-��y:�^/��s�g>�4?'/�>=q�>�ْ�!����W�<�O�>r	?�>�d��\u�*O����>Yڃ?U����K�<Z4+>9v�=�˼k�0�_�=����%�=g
����U�Y�;�s�=��=��]�k�@;�6;>A;�?�<���>^�?�&�>?l�>�Ȇ�e} ��^��a�=�]>�ZU>2�>H�پ�|��}+��PBg�x�z>���?�[�?��e=���="�=�9���ܾ��L�ط��P�<
?��"?�T?=2�?�w=?��#?�r>���],���}���B���7?�$,?���>!���ʾ)꨿��3�ȩ?�f?�=a��!��8)��J¾/�Խ��>?s/�^D~�	����C�"�j��������<��?���?YB���6�7]�����?����C?���>DB�>�9�>	�)��g����+;>�u�>?R?���>��i?��|?�jD?~�=cBO�֐��ǎ��7=
��=�m2?rF~?Qw�?�Q?+.�>�<)>�AA��$��T�M?�ˀ%��uS� z�>���>���>�}�>�z�=�Wѽݾ��@�a����=֐>�?ň�>�~�>.��>��<��G?���>�q����Ծ�=���zܼ�{}?d#�?��??͒)>�`#�O�R�b" ���>��?˫�?C�5?H�����=��Լ�(���`7�ه�>j�>��>u�=��=N�!>���>a��>��a�vL8���+��Sr��_?G18?|�>r����So���Ⱦ�����
1>��о�.O����kߖ��hѽ%��E�
۪� 7��>�����q��%ھ�M���<ʾ��
?��4>p�>!l���<#9�L� >�S�=��9�F��Ѡн�>J�C�r�ջA���
\𼀑�����u��ȃ˾��}?Q<I?�+?��C?	�y>�!>\�3����>���C@?6V>ދP�����};�A��������ؾ�{׾�c�ʟ��C>�nI���>1=3>�A�=�O�<K�=X
s=>ǎ=�R�0=�<�=�[�=`�=c��=�>R>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��7>�>��R��1�9�\���b�vZ���!?D;��O̾�'�>��=�+߾˔ƾ#�.=�6>�9b=�q��W\����=��z�A�;=��k=>҉>��C>̀�==�� ֶ=3�I=���=��O>����e�7��,��3=���=s�b>g&>Sv�>2�?e0?��K?���>9�J��*Ⱦ�J���>߈>�?��M�9�>�	?-"8?G�H??uT?��>@��6��>���>�!�u�g��M,���Q�=x��?O�?Z��>��_=�U��#c/�z�[��m��S?�Pt?[H2?$ܐ>RE���ۿ�uC��;���=��M=�=��?��?л�S�7���F����W\�>�r�>�x�>Ϟ�>�G>x�>{��>}>��=�9�2� =�#��+��R׃>]�=}4�=El�֌>�R�������;p<Z���M@=��=�F�=�:�>Yx>�U�>r�=�۱�Fc->�J����M� �=�x��4E��c��}�ە/��l8��z;>sWS>+0u�����?�,R>w�C>Ł�?�=w?��>�~�R-׾�n���a�V�V��=[
>��>���9�@�[�t L��xѾ��>�ڜ>P``>�g�=�E���A����=��$���8���>��þ��0�g�R�d���i?��f��M{�j����K?%[�����="AX?
cU?{�?U�	?�k����<�<$F�=�a�>{	s�lzo���>n@?M�S?�d?7��F��H̾>���޷>�@I�0�O���S�0���8ͷ�2��>������оi$3��g��������B��Lr�X��>'�O?��?e:b��W��JUO����D(���q?�|g?,�>�J?�@?�%��z�~r���v�=�n?̳�?R=�?u>[Կ=!�ٽ|��>n5?L�?���?+oq?��6�-��>�<��!>�:��6U�=�>���=�#�=�?�Q?φ	?�`��ة	��v��G8a���=���=׊�>dR�>M�q>f�=Qd=*&�={T>��>ܕ>'*l>=٦>�\�>6���l�$�f%?�n��>�D?eƀ>��0=����P�~<��w�lN��]�]>QhO>a� ���C�>���>���=H�>��˿��?a�꼐n ����>�X��o�>w��>!��>���<~�"?�Rq>:X�>ý?�	?�P>#�>��j=�Ѿ�>�|���8�8�(���^��x��H�>�����7���p��q�0E����Ǿ������c�؀��n>����k�?��;11h�zM��fE�V�?9��>=]G?�㾈�ڽ�S�>���>t/{=��Ծ�H��V���)|����?� �?�;c>��>I�W?�?ܒ1�43�vZ�,�u�n(A�+e�S�`��፿�����
����-�_?�x?0yA?�R�<+:z>R��?��%�Zӏ��)�>�/�'';�@<=u+�>*��.�`���Ӿ��þ�7��HF>��o?;%�?uY?CTV���[�+`2>s9?p�>?�>|?JL<?}�B?d9����#?��M>��?�N�>h�3?(�0??�+W>�`/>B�<�2�<������{�?�����Z7��SX=�B�=�@�<+l�<#.=8=<����Te��n=;s˼~��<�AM=�\�=�^�=���>��Q?��?�f�>$%?����G �b�y�P�R?�D>��Tr��������~->��i?k�?|W?�Xg>��4���\�)n�=2S�>�n>`�>_ޡ>':����R�'=v��={�>�,>5�L�e�|�MH	��վ�s�SZ�>f��>�3|>����'>�z���-z�K�d>T�Q�]κ�F�S�M�G���1��v�X�>��K?�?�=�a�X?���Gf�Q-)?�[<?�OM?=�?>/�=)�۾��9�9�J�=���>1�<�������#����:��K�:��s>�1���u����d>D��э徺�k�L�N����%�=���Z�<'n�v˾	틾T��=ʎ>���*�#�I��!���t}J?��=_��4�b�6���P�>�	�>7ƨ>��������D������=z��>��@>'Jm�������J�:�I#�>�e?t�{?�r?#��u�����t��#!�S�����;)?�%>v+�>�c�>=)��&��<���D~�� [����> ��>��[�S�Ȇ)�Ln����c��>:��>\�<�]m>QC?���>]�E?��i?N��>^ſ=J.��0l�=�$?b
�?���=�C̽�1i�D;?�e�M�,��>��'?�\:�/͐>��?��?�*?)TQ?��?�H�=n[�UF�L�>���>-W�͉��B�>�kI?}��>��X?�b�?̈1>,�9��ⅾ�Kx�u��=Jb?>�8?�b?��?�7�>i	4?�R����s�w$?�{?P�m??u?C�p�[*%?��?x� ?��g��^�>�<��?S�H?u��?��M?�
�>� <�e��K�<S�}=�RL���e�C=r|=2���I��:�=��g=ei	<,(��^)��ͽ��/=R��=�_�>a�s>f
����0>�ľO��3�@>v���{O��Lي��:��ٷ=͇�>~�?C��>�V#�?��= ��>�H�>���6(?t�?�?u";b�b��ھE�K�7�>2	B?���=��l������u���g=Y�m?h�^?$�W��%����b?��]?�d��=��þ��b���龂�O?��
?V�G���>�~?��q?��>8�e�9n����FEb��j��Ѷ=Dq�>�X�O�d��A�>ܛ7??N�>��b>�+�=�t۾��w�n��y?��?T�?���?+'*>��n��3࿕���Ъ��Cg?�t�>��3?
�R�)ɾ�S��	������(8�����M��7���͇����a�/>�C?��q?\j?ݢt?~���nc�3p����97�K��9�5�L��nQ�W�Tc���ھы�Y����L9�ှ0�N�֍�?X<!??�'�"�>�U������|���)5> �����(��Q�=�}��	=�X�=9;k�*�!�x���^�?:��>���>��E?�_�>�ol:���@�-��? 3>��>$U|>+�>�#N��,��=����վ.���I���v>d?6�K?i�m?T����1����#�!�2�'�E���1B>A
>�R�>9�P�����$� �=�%t�a/�����Z�	�8-w="N1?���>�.�>p͗??:��ᮾ�z���/��q�<Ч�>"�i?�2�>��>��ν� ���>��l?���>Z�>Q���LZ!���{��ʽ�%�>�>^��>�o>��,��#\��j��[����9�au�=A�h?;���I�`�6�>JR?���:��G<�|�>�v��!�����'���>�|?���=�;>�ž�$�ݦ{�7��ec*?�o?�_����%�G�|>z�!?9��>}_�>'�?т�>㹾�q����?i�X?x�H??�A?�-�>8�(=�m����ͽ��&�7@5=��>�\>sS^=Y�=���X���&��S=b��=�������\�g���ݼ��1;�!�<�=>mFܿ=L���ܾZ���u!����� ���ր�yE$��ܺ�����8��6������]���g�4Ǌ���q����?���?�U����{��y����~�t3����>(����ݽڌ�����b��I��J��:� ���\�
ln�b^j���	?�
�E0˿JA�����{N�>�B?u��?�-Q�r�W���K���>X[ƾ���=
���]����ؿ'�I�_P?�6?�[ݾ�Y�J\�>���=�ػ>%��>.j�����1��>�%?Z,??|�?i���ɿ����c�=�o�?^�@�|A?K�(�����!V=���>y�	?�?>X1�I�����,U�>�;�?���?�sM=��W���	�	�e?�<�F�7�ݻ�=*.�=aI=���+�J>�V�>J���SA�P7ܽߴ4>�؅>p"�ת�;�^�z��<��]>6�ս�9��5Մ?({\��f���/��T��
U>��T?�*�>Y:�=��,?V7H�a}Ͽ�\��*a?�0�?���?&�(?7ۿ��ؚ>��ܾ��M?^D6?���>�d&��t�ۅ�=56ἰ���|���&V���=W��>^�>Ƃ,�ߋ���O��I��m��=+7��2ſ�8��4S����U��8���#�>�휺�=콫���?��=���N&�>E0>�H$>�j>�p>Bރ>I�N?�0g?���>��U<��%��Kо!���kJ>��?8���羙�����!޹�-q��j#�ip,��U(�z��_��F=�B���� ��ݜ�ަX���Y?f�=�%�M8p��9>E��'�~�[��E�:�� O���p�g�?T�H?��`��LE�q��뛙�%��})?����\�}�
�]��;������!c>�ͯ=C(1��a��QY�1?��?z达�o��*�*>~2｝N==��)?�� ?#�g<췭>��?w���$���\>�:>��>���>�.>�ܯ��G轺]?wS?L�皜��ъ>����˃u�.�P=f�>;�1�����5Ee>Q <JT��E0��U������<�(W?{��>`�)����`��<���k==�x?��?�.�>Z{k?��B?��<�h����S���pw=I�W?�)i?ո>s���@о������5?��e?d�N>Vbh�6�龑�.��T�h$?��n?�^?4����v}�K�����o6?��v?s^�xs�����C�V�i=�>�[�>���>��9��k�>�>?�#��G������vY4�#Þ?��@���?t�;< �Q��=�;?h\�>�O��>ƾ�z������a�q=�"�>���}ev����R,�d�8?ڠ�?���>�������ޘ=�@���p�?�?L� �$_=:�>�_ ��Mˊ�^h�=���>�X��hl�$��b�J���S�m����ʧ�I��<���>L@����?G%�����*�ÿC.��������x?U_�>룽 )���!i�`[}���z�U�*F�N�>�>���������{��q;��Z����>Y��	�>o�S��'�������5<�>ɭ�>_��>�8���꽾}ę?�a���?οꪞ�ܛ��X?�g�?�n�?5q?��9<��v���{��]��,G?��s?�Z?;z%��?]�
�7���Z?�S���]�2J5�TgQ���6>�2?Vf�>�@�g�	=5j$=0E?�.'=AL��ʿ��ÿz��ç�? ��?�q澛%�>���?N@?#d��L`��WȾ�NM����#a?��>�⾎ ���g�g�����?�8?�RA�p)�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?t$�>��?|r�=Oa�>yb�=�񰾭<-��j#>�$�=�>���?�M?eL�>�Y�=]�8��/��ZF�QHR�%���C�#�>e�a?��L?�Kb>����2�!�iuͽ<c1��D��X@�E�,�1�߽�)5>,�=>�>��D�XӾ��?Lp�9�ؿ j��&p'��54?0��>�?����t����;_?Nz�>�6� ,���%���B�`��?�G�?=�?��׾vR̼�>;�>�I�>B�Խ����Z�����7>0�B?W��D��u�o�w�>���?
�@�ծ?hi��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?aQo���i�B>��?"������L��f?�
@u@a�^?*	ۿ�����ؾ�s��K�>�s�<��>ߓ�{t^<U0�����=�`�=���=>�(�>5ە>��<>��>�eR>/	����=���^稿3�W��U$��3��)r<%����cv��*�x�,����q2=(:��-�F���E��0�ZC�=]�;>�yR?��r?.�N?�Ȭ>6�����'�<�>����=��#>l�?!A?�gO?�J>��M���r��	��r?������X�>�ƿ>�/�>f+?�y?j���M�;�>/�>˕�<f��<�m�3�b��=��?�&?F�>]^=��C>����&��S�[��U۾b	8�e��?�3޾�ҁ�j­�i�����.�=�?�e<J��iӿ�&����W?��?���1�������ŻZ�0?�=p?�G>Ԑ��̽x�G>�����-��3��=� �q�׾'�>�sq�>�")?7�f>Bu>}�3�We8�^�P��|���h|>�36?
鶾;D9���u���H�$cݾ�HM>Iž>�D��k����� �vi���{=fx:?�?�6��?ⰾ��u�jC��?PR>q:\>X=`g�=�WM>(ac���ƽ�H�bj.=��=ͮ^>�?��=>C$u=r��>e䕾�?����>a�C>84>-�??��%?�i��q�rׇ����j�>���>���>v�>'�I��n�=���>y�Q>��pЈ�����:�Z*U>�D���SV��;Y���y=�B��$��=y܆=���H�8�H.l=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿn]�>8q��X�������u���#=���>�9H?`��p`P�">�wx
?U?hV򾝩��B�ȿ�~v����>��?��?��m��:��p@��w�> ��?�dY?�ji>rV۾�JZ�Ɏ�>��@?�R?� �>k9�n�'���?ݶ?���?w>I>��?U�u?s��>���H/2������猿R5i=]�;�v�>���=Zռ�Z�>��#��P����h��e���O>L�3=l�>�����\U�=a����g��R�F��,�>��b>O�8>L��>("�>�e�>�`�>�=�[��@h��c���J?�j�?,U	���i���<�<p=�z��
 ?[�3?_���Ͼ�V�>5�[?��?��\?f�>���h��>����)�� Q�;}%U>���>�,�>��;��V>n�;�wA�DG�>E �>��8�۾��{��A<a>f#?rW�>98�=ٙ ?��#?��j>�(�>DaE��9��X�E����>֢�>�H?�~?��?�Թ��Z3�����桿��[�n;N>��x?V?tʕ>a��������kE�>BI�<���^��?�tg?�S�.?;2�?�??a�A?�)f>݇�&ؾn�����>��!?q����A��-&�����?�b?���>v����,սʣӼ���mG����?�!\?�L&?�t�'a���¾��<z� �a2W�n�;��H��>�\>�񇽥��=>�$�=�m�o[6�xd<��=�g�>%_�=k7�*>��0=,?��G�~ۃ���=��r�>xD���>�IL>����^?hl=��{�����x��	U� �? ��?Zk�?_��?�h��$=?�?R	?l"�>�J���}޾5�྾Pw�~x��w�[�>���>�l���K���ڙ���F��Y�Žo�f����>�l�>P�>�>b=>/��>~��E��j[;H���(g��
�raO�H�Q��h4��
����׽YE>��ľ8����΋>���� ə>��-?��Y>6{�>��?o���}>��D>?�>2I�>�՝>q�">���>�3>����KR?�����'���边���l3B?�qd?T1�>Si�8��������?���?Us�?=v>h��,+��n?�>�>A��Lq
?�T:=�7�R;�<V�����M3����.��>�D׽� :��M�[nf�wj
?�/?(����̾�;׽.����n=�M�?��(?�)���Q�j�o�ʸW�S�N���6h��j��9�$��p��쏿�^��%����(�Gu*=��*?Y�?�������!���&k��?��df>��>�#�>#�>^tI>U�	�3�1�.^��L'������R�>Z[{?M׫>�>?�Z&?tS?DJ?Hh�>ZO�>�˾���>��=&�>�wi>p?C?d�?�n?��?.?��o>M��+v۾J׾�k�>�?,g6?�L?,?T �������N>���=vA�p� ���E=k=�>{�/}�<4��=��=J[? ���8�D���+k>��7?���>���>����#�����<!��>Q�
?);�>����sr�=Y��W�>j��?Z&� U=�)>g��=���ֺ;�=]*¼(��=����r;�l�<��=��=w�����k��:%ʇ;��<
u�><�?���>�C�>�@��$� �Q��f�=�Y>US>�>Fپ�}���$��g�g��]y>�w�?�z�?�f=��=���= }���U�����C���|��<��?8J#?XT?\��?w�=?Uj#?��>+�eM���^�����Ʈ?�%?�j�>���3�vF���z#��?0�?�g�(D�%w0���3��`:�`l�=�H����0���C���b >L��ݹ���n�?-��?���.�(�8��^���K��&GP?Z��>!��>e?��N���l������a>�~�>�IP?�̾>�O`?�)|?�mB?��=+XJ�8���ۥ����=9>#�$?�^c?�΅?hx?5�>�D>�"J�H��L�!��D���j�T����!��1Ʊ>��>��>�-�>Z%>��ѽQ�P�)1��_�	>��>ڟ?��>�i�>"�l>�B��8%H?�G�>����i�����ꁾ�f&���t?45�?��+?ڻ=Pi��<D�����|��>)H�?�ݫ?a�)?��R� �=�����ͥu��>]U�>
q�>3�=�@M=��>IW�>���>�Q�YQ�#f8��J��?�E?e��=�ƿ��q��p�v͗�aad<7��C	e�K���=[����=ﺘ�O��Ω���[�����ʇ������ ���.�{�T��>څ�=+��=���=�e�<��ɼyý< K=��<��=�7p�0m<�8���λ���k��n\<�vI=d���x˾R�}?>I?�+?��C?I�y>4>x
4�h��>ى��eA?%
V>K
P�����{f;�K�����ۦؾ��׾;�c�'Ο��>|3I�S�>^W3>x��=A<s��=�s=wю=��J��=��="S�=偬=���=�>lU>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�7>e->K�R�q�1�r�\�֕b��qZ���!?�F;��F̾:�>��='߾��ƾ4�.=H�6>��b=%f��S\�Zߙ=O�z��;=��k=�׉>~�C>�i�=�2����=w�I=���=��O>$���´7�B,���3=���=W�b>&>�D?r}?�B?Pk?k`�>�+*��d?�M���T>�/�>���>�J��~�>�%�>/�F??FF?=Q?#��>�ӽ���>���>HUV�)yU��.���j���%p>�`�?馀?���>�M�;<�ɾ������S�9���	?`�2?�h�>��>-c�E��D�&�q�.��ՙ�C�z�?P+=w�o�j U�L �7l���޽\��=�9�>G+�>���>,Zy>��:>�.P>m��>(L>�"�<�|=�U̻�#�<�'��x��=;Ճ��l�<ͫ�/V�󮛻��"����5�6;6�;�J<��;��=���>MK>���>.�=*
���A/>nĖ���L���=RT��v/B�6+d��O~�#/�k�6�ʊB>�X>0��w2����?��Y>b?> z�?cFu?��>���KqվuW���&e��S��x�=�>��<��p;�E`�K�M�
nҾ8P�>��Q>a�>M�
>}2�K2?�<��=���at���?�ɾ�|�<V�^�0���|������m���'Y?�=����\=�+�?�[4?�-w?�G�>P�J7޾&�>������=@#d���ۻ9�;=�m?��G?��?w� &8��N̾�����>�EI�E�O�����0����Wȷ����>���Y�о�3��h������s�B��Yr���>��O?'�?uOb�3Q���MO��������sm?�~g?U<�>M0?�;?���PN�kO��Iĸ=��n?���?;�?��
>���=������>C?��?.�?�<q?��T�}2�>ܖ�<׭8>AG��7��=b��=0O�=�� >Ol?��	?��?�k�����]��}�	1K�XLC=E��=Բ�> ܁>6ς>���=�Ri=���=�zS>�ܥ>���>�mj>�=�>c��>�A��u?��A/?R幻p+>g�L??_s>�>J	��T��	���%��M=J0�= ��3�׽��V<��>k�5>-��>)̿���?�p>=�e��)?��U�<i�`>1�Q>��>R��>3(>��>���>��?��>�s&>�*)>��Ӿ��>�a�@�%���B�|�S���о�C�>���eE�M���۽�dd�/Z��O��0�j��σ��>�X+]<AZ�?.�����l�[�)�����
?�U�>`%5?/������Nd$>��>�0�>���������3������-�?�"�?�;c>��>K�W?!�?��1�3��uZ�-�u�j(A�$e�J�`��፿�����
�M��+�_?�x?/yA?�Q�<-:z>M��?��%�Vӏ��)�>�/�';��?<=h+�>*��%�`�y�Ӿs�þ�7��HF>��o?:%�?yY?1TV�\	G�h*>`;?�^2?� s?�~2?P�8?� ���!?�5>�#?�T	?M:6?�*?]#?4+:>;��=h�[;J��<����]��o���(��2o�i�_=Ξ=�<}�j�=:��f=�T�<���N�?���;���d��<�.B=\o�=���==~�>��]?���>�2�>Rs7?in�v?7��N��6�.? �>=�� �����6.�>��j?�ɫ?V�Y?��c>��A��=C��T>.��>�Z'>x
\>~˰>'��.rE�p�=��>e�>_x�=PNL�Dၾ}~	�L���׷�<�[ >���>7|>D獽y�'>;z��.z��d>��Q��Ǻ�Z�S�/�G���1��}v�y[�>U�K?��?���=Ka�^L���Ff��,)?�[<?�OM?O�?"$�=�۾��9���J��>�=�>z_�<�������#����:�ԣ:��s>,������q&a>�7���޾�n���I���}'N=����Q=`���־z����=	�>����� �aʖ�Y����J?<�o=ڥ��?S��=���N>���>�ٮ>�2�������@��������= �>:�:>K���>R��+G��M�p��>psU?��d?4��?}����{�/�U�"p�ڧ���y��8�?���>0��>"Y>*��=ج˾����'p���]�
��>/��>|���
I�^�u��6ؾ/�_̍>4�?���=	��>IT?m�?��S?.<?�?���>���w㾬�%?�N�?�u�=�i��!L���6�c�F�{�>��+?�/��>��?S?��%?cVQ?�I?)�>rA��jA��>o�>~T�i9��N\>�L?6<�>��Y?I�?|�@>Xq4��/���A����=�>ut1?Hf&?T�?��>��&?хr�E�>P�>Jq??`f�?�e?9�=�� ?B0�>�?{\<2,?0�>2�0?��A?�ky?do?G�?N�*�}���!��;x����EԽ��p� �$�cT�<��=�%rQ:����Κ<X��<�gv=9��=F�=NP7�f�=�+�=�[�>��s>Q����0>�ľ�O���@>(u���I��!ߊ��:�ط=v��>{�?���>R#�M��=԰�>H�>���$5(?.�?�?k$#;�b���ھ��K���>�B?���=F�l�����i�u�c�g=��m?��^?��W��$���Ab?��_?�\��A:���ƾ4�l���R�K?�	?A5F�ZO�>�}?�o?�A�>�Je��~n�����d���z�OA�=Z*�>����e�4�>�H7?b��>��f>���=�>ݾQNx�k���N?Dߋ?%x�?��?�u'>�zo�(�߿:�����v�b?v{�>�֦�3#?�<ۼ]������_�����m���Rӯ�����h3��H �c���Ƥ�담=M�?du?]"p?>�c?�c� hn�5�_��~��JO��E��?��X�C�ƫ?�|dL�U%|��L�K��g���h=�i��W��ظ?�?dCK�q�?�[���&ľ.�ԾM�F>' ��y;ʽ�uG=s#ؽװ�=ӱ�<m�N��iɽu���&?�"�>��>x~=?�i�) G�Q5��=/�s�ݾ7?>�B�>�s�>�>���\����*Y��q��Ô����ɤ�>&2l?>IN?��f?n���8�~W���(!���-�`⥾�:C>Lp)>�)y>I!1��ܽ�"�^>�o6���w(��l����
�a�<"�%?.ܓ>���>��?�?7& ��a�������b(�^�<ܶ�>!�j?�M�>/��>����i�3��>+�l?��>�	�>&���>[!��{�I�ʽ-�>�ۭ>z��>��o>�,�`%\�Sl��d���V9��N�=��h?J���/�`�ۅ>	R?�l�:�SI<3��>>�v�D�!�	��H�'���>x?W��=�;>gxž+��{��0���(?�
?񄒾�)���~>�A!?�4�>JȢ>���?�_�>�]��	�:pL?��^?~1J?j�@?���>h[=������ɽ^�#�0!;=p��>��]>�zD=̗�=���#a�}�"��G=��=�O��`��<`C����<�8	=�2>�\ٿ�FO��!򾁟�� ����U��A�a�Ȕ}��u#�>7��=F���"��d�>�[����
��?;�-�}��GR���?$��?����Yw�H ����s��S�J��>���"*�S���]��"�⾏����̜��*�z�W���b��\��#?�����&���ѥ��uw�>^�;?�J�?Q�<��Y�e)C�Q�>n��g_>�b޾����-ܿT�A�S?�>�˾��� ��>#?<]g>���>� ������,�>;N?ɑ"?Ж?α�a���c/�����<?8�?i�@�|A?2�(�G���V=���>f�	?W�?>P1��E�X����X�>H;�?���?�M=��W�o�	��e?-\<:�F���ݻ��=e@�=�F=�����J>�M�><���\A�&Kܽ`�4>�ۅ>�p"�o���^�'��<�]>�ս�:��5Մ?,{\��f���/��T��U>��T?�*�>W:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?7ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�څ�=|6�񉤻{���&V�~��=[��>d�>��,������O��I��V��=c������o_��sc�uw�����G��3��1͵��_��F1��5��)��,3=U���*�>��>��>?]�>��Y?��B?�晽��h>O����)�Ft1�Q�=5	H�᚛�Aݡ�ur��3��	*�S�˾�o��}���
=����Jk.�4Kʼ��Q�]ڋ��*����g���&�EPO?M<=	���}��ͅ��&/�����z}Z���������#4�1�M�V��?O+]?� S��?��M��R�!Lh��N\?b=.�����u'�w�Z>-P��;Uʧ>�
o��!Q��xN�.�:v0?O�?E���3���6**>n����5=�G+?��?�p]<0��>��$?M(����R^>��5>5�>Lz�>��>hȮ�U�ؽ5?�S?�[ ������_�>���Y9~���^=�>`3��߼�]>���<�~���z�0ڍ�S��<e W?�[�>�*�m
�,?���y��>=�x?Ɨ?�*�>�jk?h�B?���<c ����S����Hw=��W?Wi?\�>Z��w�Ͼ����6�5?P|e?�JN>�$h������.�c�AJ?��n?�a?����TV}�;
��o���Y6?��v?s^�zs�����J�V�b=�>�[�>���>��9��k�>�>?�#��G������vY4�"Þ?��@���?"�;< �Y��=�;?j\�>��O��>ƾ�z������+�q=�"�>����uev����R,�b�8?۠�?���>��������"> ��O#�?@u?����4�>��D|��d���>�*}>;���JB�!7�:a�	I̾�_��3¾sx=�P�>�@ �[�!l9?�h��HU �YϿ����(̾Zֽ��6?�`>-����h�k|���Ō��q]�$$}�&���J�>��	>����{l���m|���:�����0�>�� ��>�R��^��!⟾E�;U��>��>���>�%���5��V��?������Ϳ����R8	���W?��?���?ԡ!?�w�<��v�ju�������rD?��r?m�Z?`7��]��7��Hj?2Z��f�_�b5��F���I>��2?��>i/�&�s=ک>��>�>�6/�)4ſ�ٷ���a�?\g�?<#�d�>�;�?��+?8@�JW��="��2	.���.��'B?"3>f¾e~��_?��p����
?�P0?�����X�_?)�a�O�p���-���ƽ�ۡ>��0��e\��M�����Xe����@y����?K^�?f�?ҵ�� #�f6%?�>g����8Ǿ=�<���>�(�> *N>RH_���u>����:�i	>���?�~�?Nj?���������U>�}?�.�>a�?��=�}�>q�=������.��L#>���=q5?���?��M?��>���=�8�2/�PDF��TR�sF�~�C���>f�a?��L?-^b>�����1�!��lͽ(�0����vX@��-�h߽@5>b�=>�>�D�!�Ҿ��?Op�8�ؿ j��p'��54?,��>�?����t�����;_?Tz�>�6��+���%���B�_��?�G�?>�?��׾�R̼�>:�>�I�>?�Խ����X�����7>/�B?Z��D��v�o�v�>���?	�@�ծ?ji��	?���P��\a~�%���7�;��=��7?�0���z>���>��=�nv�ܻ��N�s�ڹ�>�B�?�{�?��>-�l?��o�S�B�b�1=�L�>��k?�s?�/o�/󾺲B>��?I�����L��f?	�
@ru@P�^? ֗�wP��0F���$޾�(>���=N��=��1�&2���S��=�=ܻv�R>�A�>�(s>�=�>z�p>Y��>Pc�>,���A= ��M���ݦ�R�L��;�ۚ<�I����^'�>h�^���+7�*-�����=�������9n�MnJ��U>��>pXf?.S?��?��>�F�+ƽ{>�<�>�'�=6�R=�"[>nq�>g.T?h�O?�=�@H���|�����y�b����Z>�F�>d�>\��>�Ve>E�MJ�>M�>�tf>��=m݀>�Q@=�#���y>�ĩ>��?2�>��@>�mb>>��������O�����/����?K¾x�k��m��(��8���jW�=jk?�*	�*P��k�ο,��{}E?+)"�`����[��|%�k>)?�f?�n>f���H��0�Y>��м�_<�BK>��*��Y���a%���>�v%?�%W>�g>��7�i~5��?N�nf���H�>�l3?�Ψ��EE���u��cJ�0���>>��>U��j)�����x�ng� ^=�<?Ƿ�>��������/$c��C��2�O>��u>� 0=���=��Z>ч��;�����Y�@�=��=^�a>� ?��)>5�=I8�>���:L��p�>G�A>��->??��%? e
������T��7r(� Hy>�>�>��>k7	>��I�eP�=F��>�`>���d*������n>�5R>�ل��C\���h�2 �=������=Fߒ=�� �
�<���=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�h�>�p�"Z������u���#=��>p;H?�Y����O�>��x
?0?MY�,����ȿ�}v����>��?��?X�m��@���@�b~�>,��?kgY?~ji>qg۾�VZ����>L�@?L	R?�>�9���'���?�޶?S��?`x{>LИ?��?v?T��h�W�9Wǿ�I��(�ٽ��>�?�Mv=ƙþ)��xО�w4��!�l�K[9��<�CI=M��>i<�NfƾF`>r<�m`��M� =р�>��=�- >-w�>�>.?-�?�ـ�|Z�< /��
9���J?�ۏ?^����i�ҕ�<�ty=�jj�#�?��1?�ʙ��I̾���>2Y?N�?PN\?��>֗�g���&����l����;`'C>���>(.�>�:��i>̃̾��C��׆>�q�>��ھ`g���aY���>J�&?�I�>���=�� ?��#?N�j>3)�>�aE��9����E�	��>��>�H?��~?��?�Թ�bZ3�	���桿��[�^7N>�x?�U?A̕>%��������lE�SNI�����#��?�sg?�R�F?2�?7�??��A?�*f>���jؾ㨭���>��!?F@���A�-8&��	��Y?�G?(��>�*����ֽ��ؼY������s�?e\?�2&?�����`�n�¾�s�<��$���*����;��@�X>{�>������=~Z>��=��l���5���o<�L�=hB�>?��=�7��덽g9,?I-H��胾�՘=��r��uD���>'CL>������^?Wx=��{�4���x���	U�r��?3��?j�?����h��#=?�?�?(�>�N���~޾���x<w���x��v�)�>��>nik������ŗ���C��Wƽ^�>�|&�>��<>�>�C�>)p>L��>�=���������-��g��5���5������������׽�#���ض��Cx����>���%��>�{�>S_�>>��>js�>^�=��>�l>�x�>
��>�0I>�\�=���=j�<۵"��JR?s���>�'�������z1B?\qd?3�>�i����?��}�?���?Gs�?;v>S~h�X,+�on?�?�>v��Kp
?T_:=�.�AK�<�U����6��5���>�>׽ :��M�Tnf�xh
?�.?s��)�̾z9׽Q����Xo=�N�?9�(?��)���Q���o��W�lS�-?�7h��i����$�1�p�����`���%���(��p*=E�*?��?�����9,k�x?��^f>2��>�"�>�>lsI>+�	�g�1���]�CU'�����0H�>�G{?���>��I? =?�V?�2N?o��>�,�>�����>�.�=�l�>~��>C,?��?}X/?.`?��2? ��>�)̽����Ͼ�l?�?:+?h�?D�?����nV���t���=�F�A4A�3	>�a�=��۽�+�y+��>t�?��!���:��Z����r>{o1?9b�>R��>W��N�����/=`��>��
?���>9����n�c�	��]�>�k�?�S�ȟ�<�C4>A�=�0;/Z��T��=��e�kƆ=k�[�
�L�$�<x�=~X�=�����2�;>�T;���N"<�c�>�?�t�>~<�>1B��1� �9���s�=X*Y>��R>:�>5Qپ�����!��d�g�^y>Xs�?�u�?x�f=Q�=�|�=b��0b��)��:�����<s�?E#?2_T?ᑒ?��=?�j#?��>%�aM���Z������?}d-?�q�>i^���Pw���H�Y� ?(!?���a�G��S/����Q&�e�=M�S�w��K\���0�� `>�����@�{�?!��?*���wY'��:)�a�'l��^[?��>�1>z�?~m]����n����[>$K�>�<5?u�>��m?�uz?i�R?/l�=��J������k=�>��'?�Yp?��k?"�k?~C�>G��=Q����1�IaS�cO�B�z���k����>/��>�1?���>$�
>Ȑ�(��2��n�=�>D�?%��>x��>�o>vnp='�G?pX�>S��6�
��*����~��u<���s?�Đ?�.??F=t��jjB�g����p�>섧?�ҫ?��)?U�S��<�=o�˼/R��r�w��>堿>M:�>�E�=yu=��>���>��>�k �{���7���]��=?�sF?�=�k����o�ڋ��)̾����<)��[w�H��=ai>Ro���P��������As��B4��6_� k��Bӽ�^8����>W"=�!o>.�>-�<>E<���<��=X`=�X���c��Md�=��=A��=!oQ�J����=���=F���˾��}?�DI?��+?̱C?k�y>�>n�4�/9�>�ǁ�N6?�U>�R��@��R:�k��͔�A�ؾ}�׾��c�t����>6�H��l>8j3>y��=�v�<d��=6�v=)'�=̥T��I=8��=���=9�=R�=�v>4k>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>���=��8=�jq��$��K��w��H8���?U��K��e�7>�7n��)���;e��;�;K>��y=f� �@�v3=�o��L47>�=���>���=I>�<4��X�=x�<�>��>�ʢ<��x�,���Z=���=�H
>�;>]��>'??�4?Hq?��>�
&�D�پ�������>�W�>���>��k=a��>m�>�t4?9�>?/�J?=��>S��i��>X�>8��,|�lھ5���o>�C�?ej[?�̮>��G�����3� i��D'�ʞ�>ШT?8/?���>�����ݿ��-��Z9�.M��{�üѥs:Z�,v���ن�r�=�t���>,T�>�3�>��>f_�>��V>��\>���>�>[.�<�f==�LJi=�.黆�f=HV��<E ż"��;���<�����ƼxS�;P_n<[�8;3z����=Ӿ�>��>4=�>	9�=����.>+���L�B�=�>��1QB�Y0d��P~��/�@�6���A>�W>�ჽ���?Y>��@>a��?@"u?{�>�=��tվ1L���d�`T�4�=��>p�<�XR;�`��M��UҾ ��>���>3F�>v/=~���VP����;�N�N�z�1��>��h�>�ѽ��%�ￇ��K���ޯ����yd���E?w��l�o�xx?�<^?���?�;?	)�����"4�=L2�VG9>�ce�/l�
ͽ�?V�<?_a?�/۾��&���;?�½֨�>K�X8P�t���P~0�U�Ra�� �>����jоr�2��f���Տ��A���p�mɺ>1�O?���?�|a�rV��	O��q��ʅ�~h?��g?���>��?�?�K����见���=�o?k/�?.��?��
>�] >�T��[��>6?��?���?yy�?�V�1��>N_�=U�->s�D��I%>,�D>���=ٳ�=��?0�?] ?�Ľ�����پ���MD���=5�f=���>V�q>��T>&�n>�ނ=|��X�>�H�>M��>E;T>�x�>Q�>�����I��?�,�<��>{] ?��J>��l��Խ��1>�.���~���L�Ѣ/=(oѼ�����mF=Fw�=�I>=h�>?gǿp�?���<:�^\.?��
�z-o>1��>@�}=��7��d6?l�>��>�w?s��>o6Q>���>J���Ͼ��>����#�B�?��3T�S�;�#�>�s��:}C��y�;�̽e_�����΃��zl��-����?����<���?�׽Z�i�v*��	�U�?԰�>�d7?���������>���>�a�>��1��<�������?��?�c>���>̓W?j�?��1�&
3��jZ�&�u�uA�"�d��`��荿ϡ���
�Z$��[�_?m�x?�vA?��<Xz>蟀? �%�(���}U�>�!/�U*;��,<=eP�>j��K�`�ǆӾ��þE���F>�to?��?�V?�V�/C>���>��"?��B?��?P�\?L~[?�d�r]�>۝�>�X?��>}�;?m=?�?�g>�d>����o9<�<>�H�� ̖��I:��2�S��;T$��S�� $8>�ֺ�=�N.����=���=�M�� ��i�<8Vȼ9��=yu�>{;_?�?�m�>=S.?8���@����]1?o�>3ft�W i�N����1�N�>F�_?j��?�\?ޘ\>8�<��A<�Wy>J�|>!�U>}�>��>#H��;�������*9%>$�>&/�;���y�`��G�������=+�P>���>�)|>r/��e�'>�|��T1z��d>��Q��ƺ�]�S�l�G�Z�1�W�v��V�>��K?3�?4��= Z�p1��mFf��.)?�[<?OM?,�? �=��۾=�9�E�J�:I���>Ҕ�</��+����"���:���:@�s>�2���n����a>���ٰ޾�4n�P2J����P=;�@�Q=h���վU��B�="$
>�n��"!��#��cĪ�&/J?��m=;��LRV�Lk���z>uI�>�ˮ>��:��Cz��u@��K�����=_��>X;>�w��
g�/�G�">��\�>eP?��^?���?ۚ��v�b9S�=
��ё��X���?K��>�
?�0>ѫ�=`�����[y[���7����>_�>"����Q��`��Q�a<�V��>V7�>	��=���>tB?46?��`?�C?��	?.^>�'�~��R&?��?@�=*�ѽ�(O���6��+D�Q�>��(?�>�" �>��?0�?�'?ʺQ?��?	�>Gh���2@����>���>�nY�į��e>I?�,�>~MT?r�? D>$�2�����w��j��=�W">�1?�F#?�F?�I�>� 2?���#��=h�?��h?�<�?Y�s?¾-:��?rZ�>T��>��K<��>��?�/?{H?�b�?�~7?�R^>X��=�8�\3w�Pv�;*n3=4V�=eb�>;g*�F;��2��Ci�`��=-T�>���<��L�MO�3f>��X��_�(��]�>��s>W����0>��ľ�J����@>���O��vЊ�ň:���=f��>��?���>�P#�i��=쫼>;E�>����2(?��?�?��";��b���ھ�K�H�>�B?���=��l�r���e�u�L�g=��m?�^?ՄW�����b?b�^?����3;�U�ľ�h���W�M?��	?��G�wβ>N�~?KYq?�U�>K�b��m����әb�A$l����=c��>4 �h�e��]�>�e7?C��>me>��=�ܾ�Ww�8L��h?���?��?1�?#�&>��n�_��������o?ns�>�氾�11?>E����Ͼ���nG}��l�d��Pvʾ�N۾n�������S��KU����=Pj?�R�?]V?M!_? '��OY���b��҉�~�N�(A�ڮ�ߞX���*�fH���i�3���.�Xۥ��鼞A|���J�Z��?��#?D?4��P�>�랾��龇�ž�J>0��p����=M=yNϽ�@R=��`=npW����
X��t{?~G�>��>�:?X(]��8�fk4���7�B��B�>4�>Ĵ�>���>���iz �1ֽ��̾�A��M���q}>��m?��K?�e?y8%�`8�o����l�rpr��˩�j�?>�-,>%y�>BM��9ý���ViC��(z�����$��]���=�?��y>ٛ>f��?U�?j 
�#����[Q��t'�%��<}u�>�?o?=�>�ٓ>���;3���>��l?���>��>����Z!�J�{�ůʽ<%�>U�>���>G�o>��,��#\��j��"����9�<r�=��h?����{�`���>�R?) �:gG<u{�>Z�v�8�!������'��>�|?��=�;>ž�$��{�v7���X2?8!?�Ș�����۱>*Q$?;��>�rZ>��z?���>��v���w=�%?hn?��F?<�<?Ը�>�ޏ=+w��
�����佭
���ɠ>ᒓ>�W�=*Q0>��W����pɽ��;��Mk7<�Jڼ���M�{��0<S���),>bܿ=M���ܾ^��O�����V����|�T|�f	þy<��+1t�/�HO!��K���n��9���s��F�?��?�{��'A������� ��9r�t:�>2�l�[ ��,7��RI��Un����پ�����+ ��"W�9cl��]c�ak?ato�">Ͽh�� ����+�>�A�>eV�?
��)�h�q}!��[�>�L��νa/��Į��Aο��ϝb?S�?����c��9?&��=��>(�>Y=�����Z׾���:?W�?��?�	���̿\/Ͽ�'�=�?�?�F@��A?��&�1b�m[=���>}�	?�A>�7�]^��~�����><K�?���?��h=DU��K�:�e?�1<`F��A�����=���=�$=n��>J>Rْ>v����D�Amѽ�:4>[Ѓ>Ϥ�`x	���]��'�<��]>QMݽi��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=s6��{���&V�}��=[��>c�>,������O��I��U��=���j�ɿԾ5�""9���>m���R����<���=<
Ľ�����Ҿr�o��a���1�=婃>�oG>���=j��=�G?0Sf?j�>r�#>Y�>��p���=՚h�G�վy��}�N;�g���/	�����j���0<�mD+��=վ�n��]^���@��ʘ��L����~��TW�s`B?RP�>�K��6��v�G���Ӿ1���/��:�K�j��ƞj�6�f�(%�?�xN?�!P���r�$��L����{�!�8?��������I�g>�l���=`�x>(�:�>��d77�މ>��|0?�e?�o���(���*>Ml � �=��+?��?�;`<�Q�>E>%?,_*���&�[>��3>?�>4��>�	>g񮾩۽�c?IxT?�R�uӜ����>�<����z�:Ta=�>qg5�Ɔ輣�[>�А<W���\W��Đ�aм<�(W?�>��)�6���M�������==��x?f�?3.�>`}k?�B?���<6Q����S���>�w=��W?ii?��>Q��?#о�����5?M�e?3�N>��h�s�龥�.��K��?�n?�i?:F��p}������eg6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?r�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������<��=�ď��?p�?b�����k=e�8�_j��:D ��=Ca�;ϲ%�����=��6���ʾ-+�I��x��<�M_>#�@*)�v#?���k��ޣ���]|�)٤���&CP?��>AE=+��V�w��n�M�Y��K�59���N�>m�>鰔����Z�{�=p;���p�>^���	�>ӸS��!��>���Т5<-�>ǯ�>l��>�"���罾�ę?�`��>@οq���ޜ��X?�f�?�l�?Ap?��9<��v� �{��5��/G?�s?.Z?�g%�@]�\�7��NO?�kǾA���5s��t���ۼ	�I?(V?�v2���s�"�>�>�>o�=J;��!ٿ	�ȿOS����?/��?�wʾ���>0�?y�I?58�|샿$ʻ�w^F���i>�2�?��v>3�X����d���p�|�<?��@?���7��]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�$�>��?3��=u_�>�;�=�����/��[#> �=O?��?��M?�M�>SR�=��8�D/�]F��KR�;)���C���>��a?�xL?cEb>~����1�� !���ͽc1����R@�$,��߽�>5>�=>->5�D�zӾ�?T���yٿ�;����-��-?�F�>Y�	?�p�e7���X�:^?m>�F��\��닑�k��ͫ?�)�?�7?J"ؾ�-��>�8>��>�0r>�K�����1���:>WbC?��#����^�h���d>�o�?�@2�?�^c��	?���P��Va~����7�c��=��7?�0� �z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�O�B���1=7M�>Μk?�s?�Po���h�B>��?!������L��f?�
@u@a�^?*Z�׿��C�Ⱦ�ܾ�=K>�z�>�"̼��N>Μ�=�<Χ���1���f�>Bb�>e��>�@(>�{#>S��=#���)�k��7����;;��3��t�sϬ�]H��qn�C�"�s��dK��_�E������Ҕz�@8b���ν�->�!N?�[<?
@?۸�>�
<�·�=[���v��G<c��=�j�>ߖ9?_+�?6W?��[>j����v�`揿rC��:���Ƣ�>;eo>%��>�
?ک�>�����>6��>���=H���n#�J�˽oG�;�sn>��>�?���>.%�=��>ů�g庿N�Q�������p�?�%����`��6���c�>�پ�=�=��!?R�=qҖ�Adѿ_����N?^�p���#�X4H��ϴ=�+?�A[? Os>F�¾�趽��P>�r��?�����=��%��г�������>P�?�f>�u>��3�^e8�L�P�f|���i|>�36?�鶾�C9���u���H�Acݾ�HM> ž>�D��k�����vi���{=ex:?ل?7��rⰾ��u��C���PR>�:\>T=�g�=XM>=dc�P�ƽH�ig.=���=H�^>|L?{�0>���=k;�> 5��ӛH�X*�>brB>�l7>[@?��$?�F ���v(��G&�2z}>���>�	�>N >v8H����=���>0_[>h����tP
��:���\>vW��pZ�-zv��Eb=�q���~�=��=q��ˊ9�w�9=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ	g�>����i�����Z�u�x#=���>�WH?>p��b�T�W�=���
?��?V��M����ɿ�v�" �>,
�?��?��m��"��Ժ?�8��>q}�?	iY?��h>�]۾�:Z����>��@? R?���>�\�w�'���?cֶ?���?]�B>ڒ�?\�x?�}?{�@�_.J��!���3����<��=1̻>��f>K�����/��J��;���~:f�����N>xD=f�>}r��۾̭->l���Ǳ��Z=/S�>��>�/>��>�F?�?�i�>�Q�=�k���ɰ��K?���?�o�Ʊm���<�Y�=%B_�ӥ?�I3?�,S�,�ξNv�>�\?D�?"B[?���>&�J��O���6�����<�rK>���>|��>����B�L>վIYC�mˊ>�+�>dܩ��"ھ0Q���"���;�>z{!?���>8ʯ=/� ?^�#?��j>5R�>`oE�x8����E��r�>��>�E?o�~?��?XϹ��f3�9��L᡿�[��	N>��x?�J?��>����Mr���KD�L�� ��"��?�kg?�#彜?H6�?��??�A?Vf>s���ؾ�խ���>��!?���A��G&�����}?�P?���>]���ս�ּ���k���?�*\?CA&?���}+a�þz.�<�*#�e�R��;��D��>��>r���Ι�=>��=�fm�lT6�gKf<	X�=Z}�>���=�#7��Y��/=,?.�G�yۃ���=��r�;xD���>�IL>����^?el=��{�����x��	U� �? ��?Zk�?c��>�h��$=?�?P	?j"�>�J���}޾/�ྰPw�~x��w�U�>���>��l���J���ٙ���F��J�Ž5	C��]�>�@�>a�?���>�+^>5��>������9��Xо ����l������,�3�QT�����Z:�+O=�%Ѿ�����> ��d��>��?\�>5r>L��>).7�e�>��>�oU>�b�>��`>&">q�=F׫<�{ٽ7LR?�����'�Ƶ辙���g3B?�qd?�.�>�i�{��������?���?ds�?Y>v>�}h�_++�Cn?b=�>p��"q
?�I:=��8I�<�T��̺�@2�������>�G׽� :��M�kf��i
?�.?i���̾�;׽=�����u=�]�?͌)?�*�c�Q�)p��/X���R�����e�������$�R+q��돿�8�������(���,=�*?�V�?�7�=T�)���8�l���>��Jg>
�>�A�>�:�>ץM>���׎/���]�'�1o�>��z?ǆ�>�K?c�0?>0N?��R?/�>wt�>�������>��=���><�>�B?�6?��/??��.?��^>� �����˾��
?LT?e|?Q�?�'?f�m������%���P���6O���=��;�I�*�m�O=�M>*[?��O�8�Q����k>ŀ7?~��>x��>��+��S�<e
�>º
?}J�>�  �;|r�A^��V�>���?9��v`=��)>�=-O��W�Һ��=����ѐ=�4����;��l<^z�=��=$�x�-�v����:���;S,�<�s�>�?[��>�K�>�D��� ����r�=�<Y>�6S>�> Lپ}��v ��1�g��yy>4z�?�y�?��f=	�=ϥ�=�x��6Z��{����[E�<�?�O#?sNT?4��?��=?�\#?��>�&�UK��y\��P��ɱ?�,?��>���F�ʾiچ3���?*c?w<a�����2)�¾սЏ>g/��<~�����D��|�A��3���R��?[��?��A�5�6�F`辡����Y����C?�(�>�F�>��>�)���g����L;>Y��>�R?%�>�dj?�i?�08?ۄ=��K�ʻ��%��z�T��S�=`�6?�y?gR�?�Va?�K?E�I>�z��(�+�3�� [���F�������v��><��>x0?�s�>E[¼{K��1:�9bJܽT>�j�>(�?�_�>��?r>+>K2��F?>��>�#��2�T���$(|�ߔ5���s?Ed�?��,?r�=$�F�������>�4�?��?�O+?��T�#��=3����-��b�u�u��>�:�>���>�]�=k�z=>I��>�t�>������6��rb�&�?�GE?z��=��ſD�q���o�2ӗ��Of<����vMe��� �Z���=J���N������\�Ɣ��c���µ�ti����z�x��>�ͅ=���=R�=r��<�ȼ��<)�J=Vj�<��=��q�s�o<l�:�«��?��v�	�}GV<:]H= ���˾��}?�;I?ە+?~�C?�y>;>��3�^��>�����@?XV><�P�툼�J�;�3���� ��J�ؾ'x׾��c�ʟ��H>�`I�*�>�83>�G�=�L�<��=Ns=�=�Q��=0$�=�O�=rg�=��=��>+U>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�7>�&>Y�R�M�1�ԝ\�ڝb��}Z�1�!?�I;�I̾�8�>��=R)߾ʐƾc�.=��6>hb=?l�7W\��=�z���;=Fl=Yى>.�C>M|�=�3��M�=�I=���=��O>�����7�i&,�2�3="��=��b>�&>���>^?ܒ9?b^?�ˠ>yJ��˱��nʾHi�>���>b�>�Ӣ>a'�>5�B?«Y?��f?I@�>Vo��H��>� �>|�
���4�?i���if�EҊ=$=�?Y��?a��>�ۇ=���,+��&G�/����g?N}W?��4?ū�>SY�I���d&�|�.�pc��~���,=Rr�:S�7���y���e�@}�=�c�>h��>'��>�@y>��9>��N>���>׭>�>�<'�= h�Pį<�E���#�=�b����<!#˼�G����[.�8���c͍;0[;s�W<���;'��=���>&�>���>�r<#嫾�s>�꨾�R��
>���F�LyK�*/v���3�VU>���1>ʀ\>���<J쒿�t�>�k>^M>��?M��?TH>?)�ؤ�m�������⣾�s�=�D>�W�o�#�[CX�J�A���Ͼ���>1c>�Av>gb�>��N��`D�`A>d���6?�?2����=xф���o�0W��������P��i�=Ĝa?s��̻>��?�)9?!�?	� ?�����E��<LP"��~>��8�d�����<Ҹ-?0-D?��>�T��,8��H̾����޷>�@I���O�q��0�5��lͷ���>�����оJ$3��g�������B�Mr���>P�O?z�?x;b�tW��UO�����'��Lq?�|g?��>�J?�@?�#���z��r���w�=��n?���?=�?�>��=��>+�>�}
?�O�?W�?;)q?��E�H��>԰�;ʂ4>GO���>��>��=d>�?�\?�9?�چ�׃��g�����i_��E�<J'R=�`>Np�>m�v>n��=oI�==�=�Ks>-��>?L�>�[>���>��v>An˾�+=�pv+?��u=��>5�:?��0>WPr�����.>�)�p�#��f��}=����?��Z��G&=���=pLl>���>E�Ŀ�1�?Ep�={���]z?��3�Y�=���>��>+�q���?f=:�!$��\p?`^�>r]�> �C>���ʋݾ[O>#�p:�o�2�+[�1TѾ1��>�ǘ�B���@�L�������Ϊ��7���e�?����A����Qސ?D�׽��u���͈	�D?�H�>!N@?�m����Rn>_��>�u|>�� V��.���i+־��?���?�@c>��>��W?u�?��1�e 3��rZ�̮u�1"A��d��`�t⍿̘���
��ÿ���_?��x?�sA?��<�/z>�?*�%�wȏ�] �>\/�g";�c�<=/=�>�����`��Ӿ��þ�X��9F>��o?(�?�b?�6V�׽6��/>�7?��2?��u?`�2?=�<?ϩ��"?��8>(?��	?)r8?x/?��
?(H6>���=CD��=�D��S���@�ӽ�ͽ���$�0=&�{=2S���;��=��B<��?FǼ �Y;��ΰ<��-=$�=��=i�>��]?,X ?�Ӗ>W�?#�}��"�Q2���M?�X>��C�������<�Ӿ��D>!n?]}�?\�`?*�?>k+*�SD%�!>��D>��#>�"Z>� �>���İ�b�:<o�5>C�="����<��x�*���s���f2=�i_>-��>T6|>�� �'>�w��'z�d�d>3 R�к���S�V�G�h�1��zv�`a�>��K?��?$��=Oc龖M��&Ff�3,)?�^<?�MM?1�?` �=��۾p�9���J�[2���>��<x��@����"����:�,�:��s>�&��Io���j>b�;S:;b<��2=�0)Ӿ�}�=̂���������������h�L<�p4>o�}�)��yJ���ȧ�hF?�>����y��پ��\=�5x>���>�=9��?-_��P��z�>ї�>L5�=B�Uu�zK��N���>B\?�,a?M�?M��|��0W��x	�_O����w�_!?J�>�H�>Vef>��M=�:���4�T�p�H�U����>3�>�&��\��@�U�ݾv����>���>u�S��>�r>?�x�>W�Z?��7?�?�"�>{�B���Ґ&?��?��=Bzʽ�2X��;�*�G�_w�>�S'?�E���>ߕ?"?\&?��P?jv?�N>�f�iqB���>)#�>�~V�M���A�b>ƽJ?tگ>,Y?%#�?��:>x�4�#��z墽`��=��#>�+3?�[$?(�?��>�?p�Z��J��x?η�?���?��?y���X>�b�>���>1��G�L?��?<?��a?��y?��=?Hb�>�p���t�J�H�=�zX=��C�-sA=��缸�ӽ7¸��V�}��=G M=�X>�p>�J�=}�=�E�<�uO=m��>Q*d>�G����=>`�������o,>�U��\O���]��Â��2>Ê�>�i�>:�>����p=-�>���>1
��t'?��	?�h?��:0)b�Ѿ��Vm�>�?8?�ٴ=-Wo�x����1p�77=�h?��P?m��������ha?k�s?�O��Y���㾳9Ӿ���y-?�
�>�f)����>��n?Y?G�?�/c�ǲk�;כ���l�T�����=���>��!�H8w�m2�>J	!?)�>34�>)��=1���t�q哾SL?�'�?}ڲ?吏?�HR>�,~��=��p��7��i�]?e�>�㦾�"?[S�j�Ͼ���	��A��ª�oE���M��\��$��Ճ�׽�?�=��?�
s?nSq?]�_?l� ���c��^�y��2	V�%)��,���E��*E�b�C���n�qN�3s��2t��9D=G>�Ga����?<*?�@_�{�?V⸾����}N߾t�>ъR�z�\�=���?�=�i�<��� ����~��l?F�>o:�>DdD?�e��)-�3�X���Z��,��`}�>�|�>)!�>)��>a�|���4���B<@����_���#�4��>Sg_?Q�W? �o?z�.��>�����]��$�d�9����%>&ϝ=G�:>�a�	��}���[(���x�0�8��-��[��b1>�J?q�A>!��>-��?q�>CE��X���^���4�	��F8>"�J?���>���>6����>��>7�l?1��>��>z���T!���{�v�ɽ)k�>?߭>Ϯ�>�o>ζ,�4\�kd���u��t�8��;�=�h?���2�`����>�Q?^d�:Z�K<��>��w���!�ּ���'� �>"o?�H�={�;>už(��{�]3��`�&?�q?�y�����)�>QS*?�	?��>��?<v�>�é�Etk�3r%?�^???iE?q��>�(a<ש�`��R��~��=�ת>1�6>
�=��>�9��85�Ta#�S��=�Խ=�˼WS��p�*2���<M��F3>�[ؿ�H��;Ծ�����7��h;���s���烾v���v��wٓ�kȁ�8I����UOH��mf����Zv��d�?43�?B<��J��c��������/D�>e�S��l��&⯾N��셖�Y�ݾ!'����!��M���i���d���>?9>�ȿ�m���_����;>(�?zѯ?%L#��(���Y����>��(��ݾ��n����S��hC'��/?W��>��ؾ�n��u�>t~>��>Oj�>�y����Tq�3&?�!�>j8�>�%D�!Bֿ��߿j���[�?g�@Ք@?�x(����;`=T�>Yr?Y"=>��0��\�l�����>���?���?y�N=ӈV�j��{5d?V��;xeF�,����E�=r��=9	=O���QF>�'�>Ѥ�ue;���߽)@2>]�>�8����O_�-e�<��X>[�当���5Մ?+{\��f���/��T��	U>��T?�*�>U:�=��,?X7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=c6�w���{���&V����=\��>a�>,�ߋ���O��I��P��=z~�\訿Rl���0�]��<�X=SӚ��sf�!��K6�=�I�Hj��=���ma��, �>�i�>|V�>|�C>�::>�M?��j?��>r>6O����r��ˋ�]���+��>C��㘾�����Ǿ��þ_
��-����t����I>���Wm��R��RC[��2,�R�N?�ݻ>'�	�8#e�YK>*��Rӿ�U2��[d�.�澠=Z�������?i�K?5}���g���1��fI�bX��pQ?,B�<;����u�>)ӏ=�d=.�>TP��w��d"���B�~�-?9?6��`7��{2>Y���<�''??� ?#i�<.	�>�?/�����D>�-0>s��>�u�>��>�?���L�be?;K?��ƽ9G��ǹ�>�'Ǿ̐����=K�	>��G��O�.�U>��=���	��0��
]�<ѺV?	��>�L(��<�w}��@���K6=��v?[6?" �>Vyj?�??��<����.Q������=
�Y?��h?�?>۟��sXѾ����4?�h?�sU>0�p�����w*������?��m?Ȉ?�Z���z����7,��3?H�v?dp^��r������V��?�>�Z�>���>X�9�nn�>�>?�#�vF��E����W4����?˔@��?�'<<�,�ʔ�=o:?Z�>�O�]5ƾdk��x����q=-$�>�����ev���LJ,���8?ꟃ?���>ᓂ���X�D>�ʴ����?�Y�?E��LX=��T����HA�,�>ꄃ>T>��~;�?Q���F������2�
��<�=�>E@����g?���
p��|�̿}����/��h:V��
?�4�>m��0�[��N���Ɂ�I7�V6F�����"2�>R�>.E��[ȑ��{��s;�u��2(�>l����>k�S������՟��w3<f̒>���>:n�>qư����B��?"����ο��������eX?kU�?�y�?-�?��2<��w��|�p�%��G?_Gs?k�Y?:'�� ^�$#;��:k?N���ԣ`��f5�,�F���J>�|3?�r�>!_,��0M=�
>r��>\�>��-��ƿ���XO��9�?C��?o5�R��>Ň�?�,?vc�����!��}l.����;�&D?U+>}��f��<.<��B��u<?�@1?�9����]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>dH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�,�>��?U��={O�>��=x����5�GQ#>��=�n?�Q�?M�M?�:�>���=G�8��/�9OF��WR��<��C�Y�>��a?NkL?ub>&�����1�� �dͽ�)1�nO� �@�eX-��߽k[5>}�=>8E>��D�g�Ҿ��?Jp�9�ؿ j�� p'��54?/��>�?����t�����;_?Lz�>�6� ,���%���B�`��?�G�?=�?��׾�R̼�>7�>�I�>>�Խ����Y�����7>/�B?W��D��s�o�u�>���?	�@�ծ?fi��	?���P��Ua~����7�U��=��7?�0�%�z>���>��=�nv�ݻ��Q�s����>�B�?�{�?��>�l?��o�K�B�|�1=9M�>˜k?�s?�Uo����B>��? ������L��f?	�
@|u@`�^?'C�ؿ�B�����k��C��<�y=��=�Y���D>Q��=𙺽�P����5<�A�>��>��k>�4C>�{>�g>����Q��y梿����3�K`�g8���,�İ�p���v�n n�}±���v<J�ܼ�g��������$�n���wK>zaU?�k?#6y?���>�L��&�	v���_�����>+>�?��>?�(?�~�<H�v�=�|�uD���m��E������>i.c>C<�>#&?�%�>�yڽgS-=�h:>�u�>=>���=�+ٻ.�W�J>�n�>�@�>6��>�&�>98�>�ĥ�uT����L�^���hU����?�m��y�g����!#B=�վʇ�<:�2?�b)>>ښ�b'߿�͹���N?���ֆ3�kF���[�=�6?9?�^>�s߾���B�>�o�����x�>��X���ھ)�=�@ѹ>�?j�d>��t>�23��F8��IP������z>͆5?VƵ�c9�%uu���H�ۺ޾(K>dP�>a�@��v�����~���g��y=��9?f?�B�������fv�g����sR>�PZ>[�=���=NfN>�b�ʽ��H�s;&=;`�=S^>�P?X�K>��=ޗ>�g�_��.�>ͫ7>ͬ(>L�@?�N ?����������Ҿ~�z,l>H��>s �>w4>>�w^��6=���>s�#>��5<��>P�*��3����=:��<2.��K}'�ɹ�=P*���@�=�d~=��;�=�Ë���~?���(䈿��e���lD?S+?^ �='�F<��"�D ���H��G�?r�@m�?��	�ߢV�@�?�@�?��K��=}�>׫>�ξ�L��?��Ž3Ǣ�ɔ	�/)#�jS�?��?��/�Zʋ�<l��6>�^%?��Ӿel�>W��$���c;���:u�g=���>�I?���gig��>�� ?�k?:���줿�zɿ�pw��S�>M��?���?��m������?��Q�>nb�?{WY?'�c>��پהU����>��@?U[R?޶>�.���'�^V?y�?��?�KI>��?��s?y�>�Cy�Ux/�y9�����e�~=,�R;q�>u>+����OF��ɓ��_����j�����+a>�t$=i�>@j佫p��Ƶ�=�\��BW��˂e�T��>��p>�I>�T�>� ?C^�>r>�=˓������ٖ���K?�X�?��
�r�h�7�<��<=����O?�0?��y��ȾcA�>9Z?*�?�bZ?�Ώ>#��߹�� ���(��������S>TH�>��>�4Q�[>�|ξ`)6��ʎ>��>9��sݾ��q���<���>T7"?� �>;)�=L"?��3?DB�>���>�g[�#З�9ha���@>J��>�,?�4�?�?�����%(�J٘��N��q`���0>�kf?�?��>,h��#��  X=�=��G�=a��?�V?�{�����>@\h?L�"?�Zm?%h�>�?��2߾��s�Hm=�K!?up�d�A��;&�$��2?�?���>U���Aoֽ�Sͼ�!�O���'�?T[?,�%?�7���`�/�¾It�<��;�!�B�
%<����p>��>�����R�=�'>��=��l��^9�g_<���=�"�>���=S;6��3��#=,?��G�ۃ�U�=��r�awD�4�>tJL>� ����^?�i=���{�E���x��QU�� �?���?dk�?�����h��#=?c�?}?t"�>tH��|޾є�;Qw�=|x��w�>�>��>��l���ԏ��u���F����Že�W�>/:�>��?���>�r>��>����!��*Ҿ�����b�*��0�;��d(�XN�Vݎ����L/���^��Tm��q��>����B�>�?Ƒj>2^>S9�>��<��z>�j->�w>�@�>PFD>@>�>rњ��h�CR?D���d�'�o��C����(B?'fd?�'�>��i�ቅ����"�?H��?�n�?Q<v>�nh��)+��g?�2�>5���p
?��:=���;�<�]��������p{����>P׽�$:�fM�smf�]c
?1-?q���@�̾ob׽�����n=�D�?X�(?��)��Q�c�o�|�W��R��H��_h�Cl��7�$�m�p��܏��N������(�q�(=ڑ*?��?g����P?��)k��?��g>.�>��>��>0�I>��	�)�1��^�'V'�r�����>W3{?�Ï>�sF?>9?�N?�K?���>UX�>����5O�>J�M<|��>Z��>A�;?k�*?��,?��?_d-?wc>L������׾~?�
?4�?2?��?q����ͽ�+�������+{�����2 V=�p<:�ν�̉���D=�rR>.�?$��#g8��_���+n>��6?x��> ��>T2��hށ�"4�<�;�>�
?���>���{�p����q;�>�?M��c=��,>�C�=��W�O����=�Һ���=���S(7��N
<�.�=�=�n���;��M���9:�@�<M�?�!?�l�>%�>[4��4%��	�GN�=!�>L�g>��(>ܾF�������zEd���~>|Ñ?(�?��=
��=A"�=>9��J>��**���ɾ��%=m?�f%?HG?l3�??�4?�i"?���=T9�	����������;R ?��@?�!�>���4��4���q7��2?p�?+{<�����M��S�<le�<���=�Ǎ�)���o����H�>�	��!�,��?T�?KZо�Q�xx���������P�?�T4>(}�>%�.?C,��>R��諭���>Gr'>�aL?;B�>�d?t?�KN?�7>�zN��ȴ��狿�7�����=m(>?�wv?w[�?��r?�>|>g$<�G���%�����=�f�M���;�>*�>,��>�=�>R`�>�4>j�G�$ɽ��I�!+x=�v�>��>Ъ�>���>��z>�.<��H?��>R㫾��ԟ��߅���j��ynu?c��?%I.?���=&J�TF�����>X��?��?cS1?��1���=.w��$	���$s���>&��>��>uf>��=·�=#�>&R�>Ќ�*<���7��G���?��C?q(>w6���f�^ㆾT<��,�ؼ�JG��68��"U�^���Կ;����g�Q��gž�䍾}�A셾-^��wD����u�T#�>A��=�z=�1��� �}�AnϽ-��=�c=sc!>��W=�D2�䛦�
<ň��r�<|�=��E=�ύ=��˾}?-I?̋+?4�C?��y>�#>:�3�Q��>�����:?".V>N�P��~��i�;�ꢨ�1��Ӭؾmx׾��c��Ɵ��H>�#I���>�)3>�e�=��<���=�s=]�=��V�n�=w>�=�L�=�z�=���=��>�m>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��B����4�?��@��??�ዿТϿ6a/>:w=)L�=�R�:����"��8����h:�>�/'� ��Y>��5>�(�kw`��䯽"vB>�$�=��(��Y:���=S�Б�=�b>��>aa�;4��=�׽b�3�E�:�vG>B��>RX�=�<=B�=��Q>jc��}>�B>�;�>N
?<�0?��[?C�z>o]�h-Ҿ1�־�?>>�^/>]�#?�>�~�=�1�>?��3?��O?b)�>�Y��"Լ>��>��%��?u��"��ԾB�;6W�?�V�?��>�О����/�9�ZF���E���?��=?��'?vd�>�L��IѿE�B���}�Ǩ��Ծ�=�@z�]�R�O�>�QE��M����־�a=���>�J?'d�>�%>��=�Ƒ>h�>�\(>��
>!}�=��=��O=�N�=�<㕁�i�=��<)��U�v�k��h<��%=�1>��$=�����m�=Z��>�>���>��=�ұ�d�/>[����:L�s��=�া�wB���c�P�~�Hh.���5�Q�C>�,[>H���8ꑿ?��Y>6Y?>�S�?��u?�	">����wվ�����f�.TU��ϼ=r:>��=��:�=�_���M���Ҿ�p�>���>n"�>��>gP�XA4��>*�쾴H#�y��>����=U�>�;w��絿
���WJr��?�b1m?�.�����r?p�b?��?� ?�ػ�]��U~7�Z���[�>`�X��h�j+�6Q)?-M-?[!0?�����Q�nS̾����Ǖ�>ҺI�)�O������0�:��hB��^�>z����о3�a��g돿�qB���q����>DrO?D�?q�a�Y���\O����%}���=?�Ig? �>80?88?ξ���>�(��v�=��n? ��?�&�?�>l{�=�Ȝ���>�=?�N�?�i�?��t?�SE��J�>�e'=a�1>�����J>��0>�M�=6>C�?�?�q?/�:��~�� ����U����<x|�=��>�k�>ZDF> ��=��=X�=��>�>�^�>ݑ[>���>7}y>Zt���׏M?�{> �Z>�0?��=a:=,܍��]�=�́<>�H��=U�/����&U�o�����<�,I�͕=���>F�ӿ?@�?�F>�� ��#?u)��q*���J>댥>���3t+?���>B�q>)�?���>\�Z=�j�>��=<oӾZ'>[g�A!��B�E�Q�7�Ѿ&�z>�њ��h&����L~����J��7��y	��ni�(��	%=�8˧<iC�?:���Q�k�D�)�uE���?:ҧ>8�6?����\���)>�m�>/T�>����J���H���K-���?XS�?�(c>��>�W?�?�}1�k3��rZ�~�u��&A� e��`�፿����
�����_?��x?tA?�<�9z>���?J�%������-�>T/�A&;��F<=-!�>�,��z�`�ׅӾ��þ�<�IWF>l�o?�!�?�U?BjV�n��\ >�P2?��0?�q?O7?x�F?@4��rd&?L�)>��?���>�h<?�%?nw?]�V>�I>qF��QF=����vo���ݽ������H%=�E�=��:�g����S=�g�<��G�	��5��դ̼��<��;��==&
>J�>}RR?��>j��>�y#?�LA��3��죽��l?@�>�%��ϕ�a松U0�W#+<��F?�ģ?�Zo?�ݾ>0�Q��V��
<'[/>F�>�ۋ>�C�>w|8���þ��= _�=8r>ȸ�=��ܽ�!����8j��@�<8>���>�t}>U���{�,>�\�� {��)a>6�S��;��x>R�=G�r�1�ix�T��>�L?�?[��=��꾟���ܝe��z(?
d<?fzM?#"?c�=Rxؾ�:��L�K��'�>=�<x��)Ģ�B�����9�z�!;Wq>���R1��l�b>ݵ�6�߾#9n�\�I��辳�\=�����_=55��վq�~����=�
>���`� ��J��(���
�J?�Yo=�A����V��~����>>a�>��B���w���?�𚬾8*�=�b�>`49>���H���fG�f���݇>�3@?rRj?0X�? '��iπ���@�B&���㾝01=�h ?-��>��?�P>�@>���������t�j'\��@�>%~�>�h/�1^�p���edǾd�	� ��>%r?���>|c�>�P?���>�%d?�Y(?hQ ?�#�>�������p&?~��?���=mtf��n��}�öA�H��>5R?�0��=6>��?�_?��"?_tU?<�#?��3>�U<��`�]y�>�d�>�a�J(Ͽ�$%>S(m?��>��?�?�>rv.��ݾ��n����>�k=��t?>?M�?��>[��>������>�4?�h�?6�\?�x|?ɽ==�?��p�S��>�l��w~>>?�?�H?�_?�k�?>�8?�t�>䵁<�X�����h뼎�/�ѵ����nL>�/n=Meӻ9R�i�<���<��|#�]���<��)������_�>9�s>�
����0>��ľ�O��\�@>�~���O��ڊ�/�:��ܷ=M��>��?���>�W#����=��>�H�>;���6(?��?�?n�!;ɡb���ھ�K���>b	B?���=�l�����j�u�R�g=��m?i�^?3�W�R&���b?/^?�m�4=�^�þ��e�ef�OSO?f8?��G�T��>�=?SHr?�G�>hmg��!n�7���>Tb�=�j� ¶=c�>J'���d�}מ>7?f�>t�b>gE�=>�ھ�zw�$���??��?��?���?��+>^�n�@�8E�����U_?*��>�/��#?�+��Vɾ�������x�������T��������&��ԅ�ћ����=q?8dp?�t?7]?�N�ߠd���`�ɡ����U�ư �7��ܘC���A���@��m������ ������Q=aa�y6D��&�?u�%?p�@�W�>�����uξv���j>�r�������=`���=6+=�e|���Խuw��H�?�Ҭ>��>I1?Vli�I�B���A��tA�����7V>�>m�>f��>�3�<��1�+��T�����p��U�|>�\?ַe?�n?9	׽�(M��u���?�2��4���6�>��>�/�>���<Z�6���,��3|��<�tޟ��̵�=�X?�N0>M��>-�?�h�>$L�m۾pʽ��c�|%ͽ	jO=�o|?U�Z>2�Y>hZ罯����>8|o?�\�>Җ>J���j#�)�z���ܽTh�>���>�?tw>9�)�͑^������k��@����=�Bj?����PUZ� �>"�M?�Ƭ:�ꣻ淝>Y�����8�}0��!$>��	?��=��4>Dh��=��_�{�~E��eD)?�$?��}���N��z>>�|:?o�>;�W>�?�� ?��y�r�#�<�>�U?yJ?��e?r ?���<%K�զܽ�%���i<8̩>,�>�F�=/�7>�4w��[t�:3K�s�=� >{Ʋ<�gG���<�T���M=��=]
o>��ѿ�G���׾(��Ѿ�=�����%�y���Z��=����Xh�[.)�����y�ǶS�{XT�|ϕ�T��D'�?�g�?3�w��T���,��'2��z���c�>�S��Epi��)���劽[���cR�6������^�N�j�n���l�\G?#㞾��п���X�Q�N?Y��>��?M$پ��J�(�g��>/�}>��V�<��ʤ��\¿�����A�?t�?r�"����??��S>e��>���>�����4��ae��6H?��!?,<�>��Խmο��ƿ�<Q�?`�@}A?�(�����V=;��>!�	?�?>�S1��I������T�>s<�?���?�{M=��W���	�)�e?v<��F��ݻ��=�;�=F=���єJ>}U�>����SA�@?ܽL�4>Fڅ>o~"�@��ς^�=��<��]>�ս?;���Ԅ?x\�ff���/��S��^>X�T?�'�>�K�=�,?�4H�K|Ͽ��\�w*a?0�?ڦ�?�(?�ڿ��ך>��ܾ;�M?�B6?��>�a&���t�ٌ�=�H�ю��%�㾋%V����={��>��>��,����O��a��L��=�-���_¿Q�"����V�<�F�<����y#ý��/��H=�0ݾ�g�&p��l�=R��=�<>-Ά>7�6>�5?>9�]?<�t?N�>��=u�ټ�aQ	���<�^������V��3,3�݇����Q�����	�^����#�վ�n'���=�2B����I�X��Y�)W>?�њ=j�[�Yu����=)מ�>����#��ƽ?;aK��*~��D�?�~S?�l���H_��Q��/=T�&���r?A���d�ᘍ��\�=����&K���)m>�x�<V��A��T�ex/?��!?i7������B>��g��=��?�-?�+	=�.�>�n?�MY�<%��}}s>fW[>�;�>SF�>��>�k��d�ڽ��?�rZ?*T���<��E˗>蟽��ጾi�@����=q��[_�=�Kr>��<����á������\,�<w'W?e��>��)���{Z��<���==�x?q�?#9�>{k?��B?�c�<�\����S�t���w=+�W?�%i?�>ʃ���о�p����5?ڝe?x�N>�dh�%��,�.�dS��%?�n?�_?�����x}�������n6?�v?�o^�s��C���W��E�>nr�>��>Y�9��f�>Қ>?�"��F��׶���`4�<��?��@��?�=<���?��=o@?Y�>��O�6gƾb����{����p=�2�>2���yiv�N��I�,�}8?~��?_��>ﮂ�_��|J>p��PB�?f}�?�5Ⱦ���;���AV����e��=͠<�Nu�|IT����sl3�z}Ծ�w#���s�ʮ�;X�>��@0:��.]�>�����L��1Ϳ*���T���m�P���?�<�>ª�U.��)�{����Խ_���K��zA�.[�>0,>R���đ��{�w;����E��>O���.�>��S�2ݵ�f����6<�>���>Q��>�ⰽU-�����?c	���CοQ˞�~����X?�P�?č�?��?c�8<�sw���z�����?G?�{s?FPZ?�9$��f]��7��[�?��Ǿjw�����v��	�>8dZ?���>O>9�K;����>I?76F=K��HĿ�ū�FiP���?`��?.C �EO?+֟?��?\=�੿@����
�D��0V?PUV>!uξu�?��RX������'?Z^?���=�U�_?��a�;�p���-���ƽ�ۡ>��0�/f\��J�����eXe�����Ay����??^�?g�??��� #�X6%?��>U����8Ǿ��<���>�(�>0*N>�H_��u>����:�2i	>���?�~�?Aj?���������U>��}?~"�>�?���=jj�>�c�=4����-�<T#>��=X?�ͤ?�M??P�>�C�=C�8��/��YF�XIR��'���C�Q�>�a?��L?8Db>�#���1�+!�	�ͽ�Z1��z�fl@���,�ժ߽g$5>M�=>�>4�D��	Ӿ�C;?��*�߿�����Gf��T?��>�?v`�d���j�=�_?���>!z�������y
J�u[�?1 @]9�>|�ľw]6=�9'>�69>�@`>Ng�=�B/�ѷ�Ĵ >��M?��E�yԍ��V���$>���?�@�G�?�zl��	?���P��+a~����7�;��=�7?�0��z>��>��=�nv�ݻ��[�s����>�B�?�{�?'��>�l?��o��B�<�1=�L�>ɜk?�s?�do���3�B>o�?�������K��f?��
@zu@a�^?�gӿdd���<Ӿ+ɔ���=���;�&>>:H��_'=�Y
��ڽ�g8�P�=���>|�J>5�T>|�Q>_�7>���=x#��X�2?���͒�Ǽ5���������a�Ɣ	�˳��hh ��ʢ�D↾�L��顽ᆹ�-W,�Q���1P�2E�=��T?��S?!ar?^��>x��is>a@��A<8�'�zt�=[y�>��2?��H?I5*?�%�=zU���:f��6��(t���,����>�J>���>E3�>��>�䀻m
A>��H>�:v>�W�=�=�m���&=x�R>&�>��>(�>�J>�q">'�������O9d���a��U�<�?�*��@�5�jћ��ˀ�e���$[=&?f�=����"�ѿ<.��uV?k��%(��&�q�=G4B?�X?[
L>���v ��l�F>͋དྷ<�ۏ>~,�	퍾�+�X�K>�"!?��f>�Cu>&�3��o8���P��j��B]|>36?A˶��9���u���H�0jݾ�bM> Ⱦ>@��a�a���U��ni��{=�r:?�{?z?���а�Ɖu��^���mR>�W\>f=ժ=�	M>s�c���ƽ��G�hX.=L�=³^>Y?~L,>�L�=C��>5"���rO����>�0B>��,>\@?1.%?6��֙�IN��/k-���w>4��>��>�O>�ZJ�笯=�_�>�db>d4������\���?�ھV>�^��j�_�=t�p}=�:��_��=H�=c ���<��&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾL�>ʔ�B�����u���;=���>i�H?)����[��<��\?ߪ?�`����7ɿ��v�-�>�o�?&��?�n�H�����>�h��>I�?5JY?�e>��ھ�`]�U�>��??��P?P�>�a<*�_�?搷?��?O�>,��?��q?��=O��6�d�۵���t��,�>�5q=a��>�Kw>��佦g�_��ԉ�@e���������>�[`<���>�\��_藾�d>����J���S-�r�?I�>��z=�v?jO(?�E"?��Y>�$j>��">���*8۾U^K?S3�?N#��s�H=<��=H�^��W?i�6?��4;(gϾ���>9�T?)��?{oY?�H�>��������������8�<�&H>���>��>A�M�jZ>!b߾�i(��ǐ>�=�>OT���Z�=�����!�>`p?�B�>o3�=�3 ?��$?�p>�>pF�J���Z�F�բ�>���>R�?M~?�?s�����5�,N���3��Y ^�kP>|y?��?���>^����P��M��P�#l�����?/�i?��N�?*�?�>?>?�]>�|�O�վ�ǩ����>	"?�D��w�>�-M*�nc��S	?x?�>�>
iQ�������`���!���?�L[?zY)?�(�k�^�fzǾ�<G�9�DX�����;*B8�@,">��>P/�����=vt$>�غ=J&v�i/J�Z<+��=_�>�u�=x�!������3?�,:������=������A�u<�>��>Ki��]?y0s���l�5���.E��@6����k?g�?א?���e`���4P?�u�?�>O� ?� �����q��E����>c���)��5���>7Fq��׾�d���ٵ�]Z���fB�S�����>��g>�	?��%?�o>_��>y����0�)B@��_Ⱦ�E�u%�0 t�+�E�vI�1�Ǿ�������<�@���)��3�>Q�i�Ƚ�>W(�>�H�>_��>�q�>u��=k��>k��>��h>.|�>���>�1�>T�K>���<%���KR?����*�'����Ĳ��k3B?�qd?[1�>ai�<��������?���?Rs�?=v>h��,+��n?�>�>D��Qq
?lT:=g8��:�<V��l��;3��=�)��>�D׽� :��M�@nf�pj
?�/?�����̾�;׽N�d��:�=@�?��?�=?��*R�g�t�[?F��Z���=DMI��5��8� �t����ߏ�z⇿�d������>�-?�I�?�Y����}㠾rn�C8��t>�x?�1>?t�=��,:�]�w�� 9��ˎ����>�St?>n�>oN@?�*-?�E?��p?g��>|�?_���>�5�W��>s��>I*?FFH?�Q?V�=?dZ@?�|>jx�s~��\����<?�U?��?�aq>��>A{�F�+���8�[�̽�8^���
>�У=4�J>�����;���l>��><?�:�?�8�]y��s�k>�U7?|��>�P�>y<��ҿ���|�<���>z
? ��>� �-jr��h�G�>���?����=�*>��=pꆼ;뺙��=���&�=`2u�� 9��0%<�i�=%�=i�Q���9��$;w4�;���<�t�>2�?���>�C�>e@��-� �I��g�=eY>�S>�>�Eپ�}���$��z�g��]y>�w�?�z�?U�f=��=���=�|��zU�����B�����<�?6J#?6XT?\��?r�=?Tj#?�>�*�[M���^�������?v!,?��>�����ʾ��Չ3�۝?j[?�<a����;)�ސ¾ �Խȱ>�[/�h/~����<D��텻���Z��6��?쿝?iA�W�6��x�ۿ���[��|�C?"�>Y�>��>S�)�|�g�r%��1;>���>kR?C)�>�*]?M?%??\�Z>u�f�W6��n���e��=�|a>�5?���?ä�?�g?�!�>1y�=�{:�Ap��|�za��O:�kW�Y�>+(G>7�>���>�H�>8ѷ��K�<;�h=����f=�K�>��*?�"�>I �><AT>C���#D?�#?w���Y�E��I��
����t��>D?�ҝ?�^?ط�=�7���~��#��Ƥ�>���?*	�?s�?�؝�~�=V��	+��2>!����>W��>C��>$7���e=��F>���>�߻>�t��Κ���\�%� �	?91?.�@>��ſM�q�H�q������Y<�����Rc�/��8Z�C�=U���j���-����Z�ß�򒾵@���`���{���>�=m��=}�=�,�<Ƚļ0n�<�}L=9�<��=��x�BHy<$P5�=˻�����X�Q�^<TXG=\D �i�ɾϕ|?ًJ?˰-?�xB?�p>c">b�[�#X�>F���h?��P>/-8�P
����5�T����uܾ�(ܾ��`��R����>��B�P>�w,>�?�=�d<sN�=R�=\=�=w��� =G��=&��=3Ǵ=���=�B>-�>�6w?V�������4Q��Z罦�:?�8�>_{�=��ƾt@?��>>�2������wb��-?���?�T�?>�?Cti��d�>M���㎽�q�=<����=2>{��=x�2�Q��>��J>���K��J����4�?��@��??�ዿϢϿ;a/>�7>��>ĪR�_�0��Y�0�b��W�xW"?�F;��ξ_��>�Һ=�߾�uȾ�#=�05>��[=Ί�Ɯ[� �=�;��@=��l=	&�>Y�B>Y4�=K ����=�`W={E�=fVP>Ɨ��,.��4$��8=���=Dc>Y<&>C��>h�?�a0?�Wd?�4�>�n�Ͼ�@���H�>�=\E�>,݅=2qB>Ɛ�>��7?#�D?��K?߀�>q��=r	�>��>Û,��m��l�Qȧ����<̗�?�Ά?Ҹ>}|Q<��A�+���d>�U)Ž�w?OR1?�j?Q�> )���J˿��"���پO<�<dٸ�FK.=*n���7���f�|�ξy�����=R��>���>���>�|\>�s!>_�:>]�>`�>yI=�m��ċ���==d<q�=2,=SF*>4���J�<$��<��-��(̼��6��t;��O�h�O��R�=���>X=��>��u=�︾�zX>�.m�n�h�g�^<�`��{�f�@dl��W���CK�h ���G>8{>��M��噿�.?1�a>�(>,t�?ˡq?�=/�ֽ4͑������V����A��>4繼�|��%����j�=�V�¾���>M�>��>·l>�,��?�x=��j5����>t������L��Bq��A��=���)i���ɺ �D?TH��@��=V~?y�I?1�?���>�6��OxؾP0>�k��(=��.q�������?|'?�l�>���D�vG̾{��8ݷ>�=I�+�O�8���0��<��ͷ���>������о�$3�h������ҍB�~Nr����>�O?��?�;b��V���TO�����#���p?j{g?��>8L??@?6'��Yx�o���}�=	�n?~��?�<�?.>�̾=�����>�P?~i�?��?��t?��?����>z�Y���">�3��Zs�=��>��=L��=��?w	?��	?X-��b�
�����ﾣ�]��G�<�ǘ=�o�>��>�vp>i{�=.Nc=ؐ=�t]>x��>�_�>�a>3�>�+�>���M���j�?ڜ->t�>`�!?㨣>�S�>vqz�;;�<*��7�[��H��L����K�S:��`L=g�S>E�=�_�>�ȿ��?�>��1�.+&?lJ�duJ�d��<��>
��;"�>؊>���>|�>+7�>��=�Щ>���=������>���&�,��A��1?����/��>b�u:�0����]�&�����f���d��{7J���+���?"���?}�H��F�o@?Tq�>J�5?N]�{�̽�QZ>� ?�W�>�ؾŬ��͍����
A�?��?�;c>��>H�W?�?ے1�03�vZ�+�u�l(A�+e�U�`��፿�����
���.�_?�x?1yA?�R�<,:z>Q��?��%�[ӏ��)�>�/�&';��?<=v+�>*��-�`���Ӿ��þ�7��HF>��o?;%�?xY?=TV��u����h=N/L?��f?Q�?��.?�Z?"t<�l�1?EKW<=��>ٞ�>ק?&X<?j�0?�j�>m�>^�����=e)B�֌���� ��o���|��7Y=׊=]�
>iӓ=��G=��{=M���Ѱk�;�<�p��C�B��Ż��H���5=��>�"^?3��>�-b>�w4?�Wέ�/��g��R!4?%��=-mg�Q���翾Њ㾔'>��o?n�?�]S?�[>��B�>�>\s�>s�A>KT>h)�>[����X^�5#�<��>yd*>i�=��Û���������"<F�,>Z��>>|>�	��N�'>o}���#z��d>m�Q�º���S���G���1�p�v�*]�>��K?{�?X��=�_�[D���Ff�h.)?�[<?�KM?y�?t�=��۾O�9�,�J�^5�#�>_��<������m"��l�:��ݜ:��s>�-��˰����b>rt��Fྜྷ0n��9I�I��ޥY=��f�X=hH��)ӾQ�~���=qm>�)��K;!��4��%調n}J?��i=Lp���
X�����5�>苙>�N�>�F���q��:@�Dt��{��=�)�>�<>y��8�PG��o�$�u>4�N?]]F?��z?sc��-�� S����r􇾾����?��>��?�=+^>����]�t�\�J��-�>��>DK��gJ�M?Ͼ����r�ھX\\>��?`�=>�)�>W�a?*�?"6�?%�J?�'?%`�>����������/?)��?�4�=�,�5�t����:�-�PM�>R>?yW���6>��+?�@?quE?4�X?� ,?��2:����M����>�I3>/�>��������<
�d?R?�Oh?��q?�e>N�I��%���k὎��>G�>�W?I�?ٝ
?�y>��>���GN�>B3	?G>y?q�q?(�?�����>p��n��>c�<�d�>�?WW:?��[?pR�?�H?DT�>E艼I
J� f�w,��h!$=�D�=m�-:)��=�s�=�䰻��W=���=i80�}׼m$3=	=>��N�Y7w�]Ew=�9�>H�u>k��b�2>}?žŊ�ǿ=>� ��қ��kf8��&�=�h�>�s?E��>2E%��M�=�H�>���>�(�SA(?JE?�=?��<�b��ܾ�O�Y�>l�A?��=N�m�W��u"v�=�o=�m?Ѽ]?��Y��(��BQb?�w\?�_��	2�bB־�a��\�΂T?��?�G�)��>�҃?��q?��>�Nk�m���s�_��>W�J,�=�H�>����zb��å>�5?�}�> �O>d�=�:辅#w�G3���	?��?�u�?*i�?�G8>*zp��y޿�������q?u��>��˾��(?����;x���k�Z>�NȘ���˾�%���
��R�O�Ky�ʚ��#�=��?\f?Z�~?�K?c��Ab�Xp�.���HL��n��$�B��FG��>�Gek�v�����꾸�N� �<u�~��B�ɑ�?��'?{1�7�>ir��H���;!C>���Dq�4�=����<=a�V=h��-�����< ?N��>���>�<?L\�A>���1��8�\���D�3>L<�>�>�[�>2�:�.�W���ɾ�5���1Խ<aZ>|Qh?8?&$f?�q�ԧH��V������퀽#�����Y>�Q�=b��>	ؓ��)��^%�j�C��Rz�Rc�&����?ﾎN2;�l?;��>�*w>�Y�?�ȵ>b	���������w?�VO���Fb>]�|?�2�>9a(>-�&�PW'�P^�>W�j?ﮠ>�X�>��Η*�]�_��-X�>L"?N�C?�?���<�R}�y�'�y����Y�b*�>���?	�#����
ш>�7z?��[�P���>|�>VP���wӾ���;�A�>��6?�<=��>�$þ�u�ુ�X�q��K?=�D?�<���T����=�jV?��>�-�>��?\?��ھ�To�4��>#f?�BP?]�_?+a!?109��ی�D�T�+?�<x���>|>U®>�D�<A�S�ʣg�����NF>p7 =��H>P���0����>�0�>S	>u9M>�8ۿ4�K�9�׾�T�����#�2������?ā����������y4z�u�Yl5��UQ��a������i�.��?\
�?�@��~��uq����~��c�R��>�z�m�o�E���s������]�dZ��%��6O��>k��g�3Y-?�v̾�ѿ�T��f�྾�J?���>'�Y?���2�ߢD�jެ>p�=��d�8��:Q����ҿS$ž��u?B�?W�i�����?�^[>�˛>��>�]D��;�-nP�[�<?,�)?\�?q揾Ϳ�%ƿ�x�����?��@}A?��(���쾘V=���>��	?��?>�R1�xI������T�>�<�?���?�|M=v�W��	��e?�z<��F���ݻ��=q;�=�D=���ٔJ>/U�>W��nTA��@ܽ��4>څ>�~"�r��r�^�.��<͇]>[�ս�<��=Մ?�z\�qf���/��T���U>��T?�*�>M;�=��,?M7H�E}Ͽ�\�+a?�0�?��?%�(?\ۿ�nؚ>��ܾ��M?%D6?���>�d&���t���=�5��}��'�㾟&V���=$��>��>*�,�؋���O�G�����=���+Ŀv�������=G�
� ��G��]����j&Ͼj|���4���=GN�=*�N>��w>tN>`�l>B�]?:�f?��>(5�=Y)Ƚז��y߾�3�=�"d����������ν��{��U��}���� ��sd׾�cM��p�i A������0���H[��=]�b [?�d>�V���g��._>�۾y����?���6���Ͼo�=���h�.�?tN?"K��*ll�~��)��=�i�\T,?V��B$�������*<��ѽS)���>*}�<��	�G�X���m��l0?��?䦿�%��k�*>����h�=Q+?��?��<Rp�>��$?o�'����}\>>6>���>*��>�>jr���
ܽ]?%�T?�] �����k�>�-���p|� �Y=+�>��4��MǼ�z\>�h�<r����h�׌��ٴ<�'W?��>S�)�0�d���)�E==u�x?��?�1�>�zk?��B?���<2d���S�s!��:w=��W?�*i?�>x���о�z����5?�e?��N>�ih���#�.��R�#?��n?�^?����v}�,����+m6?��v?s^�~s�������V�+=�>\�>���>��9��k�>8�>?�#��G����Y4��?z�@u��?s�;<z#���=�;?,\�>��O��?ƾ
{������c�q=�"�>⌧��ev����S,��8?٠�?s��>��������=�A���/�?@��?�V��PEV<h����k�x�����<U�=��I�yl�i��\8�koȾ�u	�Lx��u{ռֶ�>E�@2��U��>o9�⿼%Ͽ\N����Ѿ��w��_?�T�>����A����l�u�m���A��J?��쉾�=�>}0<>o4���W����r�,�4��M��#�>ߜ�<d�>t�U�}��U�����h=] �>���>��V>����˾�v�?�����ÿT���0�8f?d�?��?b$?D��<�N���P�{�"��Ad?c�t?�?m?N�	�LuI��S��[Jr?6	پ���$��L`��_�>��4?��>:.�Ǡi�L��>��>Ѵ<|��m�Ŀ�9��0����?>�?p�����?$�?<�?�
&��9��kRH���.���?���V?�ъ>����@�m�D�"��j�(?��X?y�>�UG�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?ֵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>bH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?�r�>�B�?�>�=�?1t�<c�ܾGQ����g>��>r_��"�?o_?}��>5�=��Q��5��?�&eO�ԙ��(G�s��>�{N?��1?�õ>����Ƨ��Pb/��A�7�L��/нf���Gk�Id!��Ra>d�f>b�>���������.?/~6���1���vXb���M?Ù_>��?�%��ÿ��J�<�2l?^�}>p��D��w�������?<@�= ?S"����Z;u�e>�AM>.�=p��=:ͽX���Bm>�7]?v��>��	N���g=��?)@�ӵ?β`��	?���P��Ta~����7�h��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>!�l?��o�N�B�}�1=5M�>Μk?�s?TRo���m�B>��? ������L��f?
�
@u@a�^?)�࿞�������j����>��}=���=���Si�=�$��D�c=_�Y�Ҩ�=��1>�B>n<}>�}D>�>���=K�{��B�>���A���(�2��/��&�\�]�O����������9'���Ⱦ�W%���A�����h�v�p��L�;]��=N�U?�'R?�&p?� ?�mx�Jk >j���.�=g�#�e]�=�(�>�h2?��L?g�*? �=/����d��_��s9��P뇾@��>īI>�\�>��>e�>-� :;I>l�>>�o�>;>̡%=��� \=O>Pf�>C��>�|�>�6>���=�D���ʸ�9�_�t"*��8k�*�?�Ѳ�b7,������<� �ȾSe�=�f?Ҵ�=�����տb���+y]?���*1��K��?^=>O?T�[?-L�<䕾w\���u>���P��~P>1�堬�710�B%>��(?E�h>�u>�t3��z8���P�7���E}>�6?/.��׎7���u��H���ܾ�P>d]�>m$&����@>��Di�eV}=�9?�3?������S|v�|*���Q>��\>u�=9�=�fL>�Eh�.�Ƚ�#I�K7=.�=��_>�Z?	�+>
��= ܣ>�s���UP��u�>v�B>�I,>]@?b*%?j��B����|����-��w>&N�>��>�d>mkJ���=(f�>�a>��e���r��6�?�XRW>6�~���_��Du��y=�C�����=�?�=Nx ��=�;`%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿxn�>4��]������u�sH$=��>�6H?�N����O�j>��{
?�?-^򾢨����ȿڀv�:��>��?���?��m��@���@��{�>՟�?#hY?Mqi>Ya۾cyZ���>G�@?�R?��>>@�K�'���?��?_��?"j1>}�?d1`?���>��=�F��ݶ�[���cR=%���Ӗ>.-�=L���Y�R�������p�F'�V>�y=B�>kF���v���n�=d+{��:��Ws��>�>�d>��/>4¥>��>�º>��>T��=�M��Z������]V?�8�?`��'p�v�L��>L�z�?��5?��=���r�>X\Q?r&�?{�`?���>���e晿M���Hj��z[�<�c>1��>9��>�C����:>�(þ�R��}�>+f�>����ھQB��r�ؼ �|>8,?�i�>T]�=�Q%?j!?Wj^>���>)�S��ڕ�?����>?��>��)?���?��?�Q���q+�jz��k*����b��fn>�L�?��?��{>�*���Ȋ���K��+�&㜽��?��U?��o?�ؗ?�3<?��7?C�8>���T����E��JD>X�0?�>��ߝ7�6;,��fd���?��?u;�>5���z#�qRֽl���ᾃZ,?��b?�3?Ǹ���d�+�� =�ݻ�X����߽�/E>=Z>�C��Ri9=�4>/�=R��ցL��s��W=��N>SVH>���+���*?$�p��ԭ���E=�����J���>��>�p����P?�D�-ƅ��)������͌��U�s?��?�?	V'��"{���I?&��?�S?'<�>���h���=��4���c��$�N/�<?�>J�"�xpؾ)@��L�������XL2�m����C�>�S>
� ?��	?)����>��;� M�7"$�R����x��x�J�Y��G�+�+�1���%26��ك;�j��SBo�6�>�Ի�;�>�%�>aAS>�?�>��?���=P��>8è>�r>J/�>��>6��>�N>�k�<�`콯KR?����Ͻ'�O��C���0B?�od?�3�>�i�ȉ�������?���?r�?�8v>1h�u,+��l?�>�>���q
?�P:=0q���<)T��%���@��j0����>�O׽^!:��M�dpf��j
?�/?!���̾J׽؛��Ё�<R��?=((?��/��L�9�l�	mW�UlX�Z�Ik��AϦ���'�7r��莿`؂�;����� �=:�(?��?����W�-߫�"p�&9D�ѥZ>���>@�>vR�>�k1>9���5��\a�b��jRp�(�>�Au?h�L>b�C?�E?}!Q?��P?J�>W�?L8�ͨ�>Ж̽n^�>�:�>»d?&B;?�H?
HF?Y�f?�6s>6���ﾷ�� �K?= B?e>�>��l>�E(?;�������J��"=�P#�R�� r=�>~�
��}=�"/>��4>�X?���ɬ8�����Pk>n�7?
��>y��>���#-��5�<w�>�
?
G�>E �!~r�c��V�>���?���E�=��)>���=?�����ҺZ�=������=�5��!z;�ee<���=@��=�Mt��&���7�:���;�n�<��>��5?�xA>R��;$/$��m�J�,�����6>���>	�>������9f����t���>�"�?�I�?r�(>��>3��>�{Ǿ�Ⱦ��׾��Z��x�=0�R>|�h?��l?ꃈ?�.�>��Q?f��>��Ͼt��n���p[[��&?w!,?��>�����ʾ��҉3�ӝ?X[?�<a�и��;)��¾�Խα>�[/�l/~����,D��煻���u��1��?￝?�A�W�6��x�ҿ���[���C?"�>Y�>��>Q�)�p�g�x%��1;>��>iR?K�>��O?�-{?֡[?âT>��8��3��|Й��Q4�J�!>g@?��?c�?3�x?�n�>w�>�)�u5�F^��K��s��2߂���V=<Z>���>� �>�ȩ>R�=��ǽ�f����>�0H�=��b>G��>Ǳ�>���>�gw>���<H?O5�>wk��|��_뤾{�����<��su?���?�+?c=�o���E��y����>�d�?U�?t�)?d)T����=м�ᶾ��q��q�>6��>D��>%h�=��H=Z�>��>Gp�>����x��m8���M�z?�E?&¼=Kpƿs�q��p�v��Yϔ<Z���c'f��)����W����=
������먾�RY��ڠ��D��Z��w"��{�v��W ?��=��=���=i4�<�Z׼Ex�<��h=���<�1=�Ӎ�8��<��B��,�*􌽍�Ӻ�{<��<=\��;�˾��}?�9I?��+?��C?��y>�=>}h3����>�����@?�V>A�P�䋼��;�٬�������ؾ�v׾-�c��ʟ��J>�[I�3�>u93>UJ�=>a�<>$�=�.s=jȎ=�P��=$�=�Z�=t�=%��=�>T>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>_)3>�v>,�R��0�4	Y��(f�B�X�4�"?��;��y;\҆>��=/p߾��ȾX0=�V3>�x]=��؉[��#�=�O��qA=�^l=04�>|E>ּ�=�f����=��Y=�B�=9�S>�I��d�4����B=�i�=e�b>&&%>���>6�?�d0?<Yd?�8�>�n��Ͼ�?���@�>��=E�>���=�rB>T��>��7?��D?c�K?Ո�>讉=��>��>��,�K�m��e��ǧ�{�<~��?�͆?�ϸ>ZXQ</�A�,���d>��Ž�u?P1?�k?��>��S�׿�P�X{%�終�� �i�]�q�9��z\���#c���<x)�=S?�>y��>���>+�&>�X6>��k>Ɯ�>�r">sI�<6����<�����:RA>��l=,� >�O���>5�Y<�� >�qĽ�}���g8���<�3I===k��>�y=�ث>�/����?�F>7jp��&}�S�ȼ�Y��5c�J�i���*L��i��i�=7a$>�u���ܚ�c?%R|>�dY>�h�?k�U?���=j��<A�׾3٣��m���]P�-HY>b��=#��9�/p��SO���þN)�>F�>ɱ�>��>��*���G�*�;�I̾��,���>ބm�y�o:���v�k�W���&X��,�c�'��H�;?B�����	>�+m?�m7?'�?���>��lQ���=^y��#k��2*�>���1���?[�(?ȩ�>����"�J�+N̾p
���շ>�I���O�S����0�Z��w����g�>�㪾S�о�-3�m��������B�h/r����>��O?��?�b�O��SO�[���̅��_?�dg?a�>(J?;?ж��	���a��ᠸ=��n?���?�6�?�>�F�=�^νe��>�$?��?���?)�}?��U����>kyJ���>HY���.>�(> ~>��%>��?A?{T?����������S辒?A� �G=֟�=�+�>]��>t>j��==]{�=8~N>��>gc>�'>���>�!�>�+̾�Z���	?<Z>�|�>�O?� �>ci>�K���7�\g=�,7���r��G}��R��tz�9��<.{=R��;�G?hTѿgx�?�"1>9"�1�F?�o�z.~�'>Z�>���aU�>�;�=�6�>u�>ǡ�>�#>�×>>�
>��ξF�
>j>�c0'�u�B�W�J���׾��x>i�������4޽�tN�w����j�wg�� ����B���;[N�?�X��]o��#�� �.?x��>�/?M ��lC���#(>�b�>(˗>y��������U����
d�?ǩ�?Ef>�>�X?80�>�C���x��/d�i#a��)c���N�'[��"���(��z�3�&�|��=?<�i?0R\?j>�<�u>[��??�X�'���e�>�(�~�E��%�=FS�>�}���ٟ��c��hP������<�h?���?h�-?���ǆ!���t�[�\?n?��|?�2?��h?1��|�?�t<�5?���>@�A?��?�E?p8�>��I>��ż.K������Gw����������8Ͻs�����m4 �У�<�`c=�Ov�)���iSD=`t���W�퟽��-ۼ�b�~F�<���>]�]?�a�>됆>տ7?��{�7�Gخ��/?!9=儂�����n�9�>�k?k
�?�+Z?1xc>YB��FC��&>kt�>z�&>�[>�Z�>��FcE���=�1>��>���=LL��a��ۘ	�ģ��^��<a?>���>d:|>C��S�'>�����z��d>��Q�Bĺ�f�S�i�G�)�1��}v�e�>��K?��?8��=c�W���Ff�f/)?AW<?�HM?�?|�=O�۾��9�-�J��4��>�ɩ<���<���D"�� �:�؄�:��s>�(��3١��Y`>����h߾{m�=VI�b�辅Ve=��o=G=��#�ԾDq~����=��>[羾+� ��<��!O��i6K?��o=�x��J�V�^R���e>m��>�o�>�BA�Öy��@�ͬ�[��=�k�>�\6>q,��f��2G����>�A?M�??�%�?�2N�����5���
�����n�����<?�3�>���>�&�=܂�=K
���#��f���7����>�P�>���AY�G��:2ʾ��$����>3\.?��h>[?�Wg?�	?�@l?��d?&�&?]]>0׽�ƾ�(?���?���=��(���a�+�1��A�!��>Ӥ*?����]>� ?�!?E�6?��S?�(?/��=*U���O��~�>T��>�.I�.貿7cz>�S?�{�>�Z?�u?X>I.A�����6L����O>��9>1?�b?�A?�Y�>��>�C��Ӡ&>z�>��X?,�w?zmv?5�=W?�9>���>�<�< J�>0��>[�(?W9Q?Bs?�??���>�S8������ν_�g�&�C<��=��<ܞ�=� �QB��q,]��=Hb
<�G�K���a��M��y�����<D�>��s>� ����0>�ľXT����@>v����V��/�����:����=ar�>2�?W��>Hv#��z�=v��>,[�>\��]9(?��?�?��+;��b��۾[tK�-�>�B?3��=)�l��~����u�ٯh=;�m?��^?��W�l(���1\?��\?��Ǿ1�/����l���"��� ?�` ?�Ӕ�1��>��?��n?w6?�B��>B�����Gz��״���I>d��>�c޾5��Y�>��Q?R�>K��>0>�D~�����V��c7?�D�?�d�?/I�?��7>�f�J�ڿ;׾�~���^?L&�>BQо��??������J{�������� W���g���A��ۖȾ��-������gݽ��>A�?��c?�?�F?"�	�^�N8���GE��f�=Pʾ��$��~T�,�S��� �f�Y�Š�-%�i�p��]�=�!|��YB��>�?�'?p04�)&�>WX��)2��;��A>�V��3�� �==z��9�+=|VV=�(j���-�꫾�M ?u�>��>��;?��[�t
>���3�%�5��;��A�6>Y�>�G�>Lx�>U��;P-��
�!�ɾ�w���̽n>�Y?a�:?]�p?=�d�Y�;�e�o�[O?�����H�����F>zX�=��>����J���K��C�Ou� 徵졾����*<�7H?�Ϝ>��B>���?���>J�"��`w�i��r�)�L�0;R%�>6??b��>6\�>���J��}�>�?��>��8�Q��;x`A�=
��;/¾�?�=>�=1>Xl>�2���s9�݅���ݔ��r���> ��?�c���lr�90f>��\?�w��xT��'��>oC����y���f���4><K?���Z?t=��ݾ�������WE�590?��G?�B{���P��L>�6?�Ŝ>2��>�<�?�#?D���]�b�f�?��}?tNS?��W?W��>��o<���z���*,���>�}i>������=>vE��]F�ƽP�脐=O�>���=�|˾��/:�=,�y>eɐ�#��>6~ۿ��K�5.־Q���R򾲍	�����5d������-��y�������\z����f(�n
W�g�Z���.k����?&��?����^"���v��~~������\�>��n�����'h��+���>���R�񒮾���уM�Qlh��vc�d�>?B�˾2׿����s�ľ#C?���>?�?Y^��뾪KH����>���=�@N�K%��X��5�ȿ�(���f?�?U,�Ws�t��>�(J>���>�^�>�������N�<�#��>��C?��>�F��'ÿC�¿��<}�?.@}A?��(���쾈V=m��>�	?�?>�S1�\I������T�>[<�?��?d}M=?�W���	�@�e?�t<��F�q�ݻV�=j<�=�J=��S�J>�U�>���UA��?ܽ��4>Xڅ>�v"�5��w�^���<��]>�սy;��5Մ?*{\��f���/��T��
U>��T?�*�>a:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?$�(?8ۿ��ؚ>��ܾ��M?^D6?���>�d&��t�ޅ�=w6����{���&V����=Z��>\�>,�ߋ���O��I��[��=t��zÿ�A	���q�;v���ZEȼ��ܽ:����8����p��g�ň/=�y�=I=5>�_3>��>˂ > OV?Hw`?q��>ֶ�=X��Z�e������3d=�q���Dy�=��D��^K;~����5����6�NӶ�Y�+��dO=r�W��V��`E����\��[�#�\?��V>�p��wR�t�.>9ӏ������5%�
\<l�˾ez<�&.��(�?ie3?�Ð���]���Ҿ�&�=�y��B�N?�L1�\��s���>{�> y�=&��=;Uw>��>?���N�N�Xe�OU0?�#?T�������$7>�C彚�=�'&?��?��Z=8	�>��#?�m�����c>�-U>ȉ�>��>D�=�v������;S?�+Y?�ܽ'˟�ۿ�>GȾ؝���X=�A>�?�l�=ߠK>&d<%���E<�{���Ѓ<�bV?�4�>p(�F�&���˖&�,N=b u?
;?С>��i?B;@?*?/<����oT���
��?q=�{Z?��i?��>��i�D�;������4?{�d??Q>�Iu��徉--�=���?p�p?8P?�׼_\~�+��j��P6?T?*.f������k �����>k�?�D�>~cR�o�j>S;]?c� �D���Cſ&�F��̒?�@#��?��<�?�"�>�4?�B�>�Ɯ�.�(�R������s��I�-?���
����w��P��l
?�ۓ?~�?����"����=�,��\B�?D͆?�¬�C`�<wk�F~l�ѓ ��<���=b ��q1����DW8��0Ǿ��6��wx��Ӫ�>p"@f�ݽn��>o�8��"�X�Ͽ򁄿�Ӿ��l���?���>h�ֽ�J��Hqi���t�%|F���F�ń���>A�>"7���	���{��};�u���;�>���dM�>I.T�񵾂���X0<���>NK�>$f�>�C��Ar���?����2ο4���i��yX?�?�b�?F�?�<Q< �v�+�z�96�>G?��s?DZ?Z#�x�]���:�5q?7ʾ��l�"4��TT���>��-?Ƙ�>�5�Gmw��0>�]?��e=N9����s%����վ.�?�s�?���-g?���?ID(?�1�y%��O[��+�ެ.���6?
Y�>'����.�,F��覾�f#?��O?ND��2�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}? $�>��?�o�=�b�>�]�=���-�qe#>I�=�>�Р?z�M?L�>�P�=F�8�u /�:[F��GR��#�
�C���>g�a?i�L?Mb>^���	2��!��~ͽ�a1�0�<X@���,� �߽�-5>n�=>3>��D�?ӾDb@?2�F�e��S4��LEL��K_?W�>�?���ɐ�����wߏ?To5>d:"�;������A��׭?4w�?�`�>�ξJ3�=�>�.�=9{K>�d�=	<��s���k��:f?
c��@���́���B>��?��	@�[�?n�]�I?>��{����S}��y	�8���d�=�5?a����c>��>.��=��x�3
��Qt��G�>$ �?���?���>A�f?vFi�}d=�n�D=9��>�#c?��?��F�%����0?>�x?��i����x���_?�P@lY@ɤ[?�פ�b~ῠ�����������>)�=q�2>��H�]�;=1�<������ј>���>*6c>�+�>��U>�z2>z�*>}�����|X���J���6��
��U����4g���y�����#��O��S+���jӽ���v�d���	��l�=0�T?�R?i�p?�, ?ކt��=%>m��,�=���p�=���>��2?*�L?�G+?)�=Lw����c��B��/����-��/��>�J>)D�>��>O)�>/�:|�I>�=>/�~>�T >K=9��O�=��M>�y�>F��>��>�~R>�)>8������vM�/�@��h����?W����3?�s���Cw��F��K0�=�?�3>Ӭ���ӿ�娿{k?HԲ�\*1�a�+ޢ=��E?-)N?v�>�Ұ���q<*J�=�� ��pc���>ځO�������)��M>I�?�f>�u>w�3��e8��P��{��ki|>�36?�趾C9���u�ŲH��bݾJM>ž>{D��k�>������ui�e�{=�w:?��?�4��Jⰾy�u�5C���QR>;\>JX=
i�=XM>ec�d�ƽsH��j.=׾�=n�^>T?v�+>4��=�ң>�E��(BP����>�nB>� ,>�@?"%%?0��S㗽�����-�w>7V�>��>�\>jJ��=�j�>��a>P��c�������?��mW>J]~�	�_��3u���y=����=��=d� ��=��&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ#��>!G�vp��/���u�Z�'=�K�>[KH?�b��;�N���>�L�
?g?Sg�Ҥ��~ɿ��v����>Z�?��?!�m�j#����?�)F�>>��?�^Y?��h>K�۾ [�회>��@?Y�Q?@��>2��'�)�?�?}��?�+H>���?~l?ȫ�>��-��~6��&��a��.�=s?�:)�>ٚ�=�h��x`C�q��9���j�{q���Z>Eo=䅵>�,��
˻����=peƽ3j��Q���t�>�p>�]m>5��>�i�>$�>nװ>-�=R��f�x��ܙ���N?�?̾Jǈ�w�ޤn>z�f�
&?��9?�_�>IP�fU�=��T?�}�?Sc?���>���{\���˿�ҩ��1�=4>�%�>b��>��>��Q>~t��S�'��v�>�U�>Ŀ��][�h�A����8�[>n�?a?r�> � ?l�#?-�j>#/�>�XE��=����E���>Z��>sC?��~?*?^ʹ�:U3����3硿�[�ON>y�x?<X?�ȕ>ĉ��C����#H��H�)�����?�}g?K���?T2�?E�??��A?{f>T3�8 ؾ]ǭ��ـ>��!?6��{�A���&������?#*?���>觑���ҽ�5ؼ��9 ��1S?�1\?�G&?�����`��þ#�<����r��u<��@���>��>�Q��T�=">>��=�`m�S�6�m�Y<���=5j�>ʵ�=�E6��͌�00?ӛ޼f�=X=ƴ��r0`�R��>��b>}����Z?ځ�=��o�)%��Q���wK�����?�c�?��?"�Ƚy܆���b?e	�?��?��2?be���G�������J�r��Jt�<DV�>!'
��׭�X���lh�����������'�� ?q:�>�?(�?�3)>�t�>X>U�(R2��-��Pپ\I�����cF�)!3��_���|���)����x�Ǿ���I��>űP�7��>\�?d6Y>���=��>�=�O�|>��>�ܬ>��>u�v>�>�p�=��<�ِ��KR?�����'�~��Ͳ��l3B?�qd??1�>�i�9��������?���?Qs�? =v>	h��,+�~n?�>�>B��]q
?�T:=+9��:�<&V������2����7��>E׽� :��M�:nf�uj
?�/?�����̾�;׽DN��`�M=s��?�'?�7*���M��En�%gU��T��}N��q��£���$�UEn�^W���a���̓��&��gZ=�e*?|�?D�������*pl��IA���o>�)�>��>���>��F>)�
��0��jZ�S�$�53}�G��>�(z?�2�>i~=?��!?�:L?b�6?�s>EE ?�|��e��>�:�>�ʜ>C�>��v?i}+?�$G?�/0?>�I?欌=7�����J 
��\?[hR?@��>�g�>��5?֜����(�C���F�D�����Q�=�f>��)���ֽ�>^>7X?,�Ϩ8����k>}7?�q�>���>���Q%��|��<"�>j�
?�B�>� ��}r��d��e�>L��?��u�=z�)>��=�����r׺YQ�=\V¼m��=x�����;�B<[��=���=��x��+��l��:I2�;�ï<���>�~*?�(w>�y>��
�-���	/�&��=��6>��w>1+>�J�4��#���X7d��"y>Z��?O:�?�g6>�_�=G�f>�$������b����c�>�m>O?9?�IA?1�u?#�-?ZUK?y2>���/+��zV��
#����?w!,?��>�����ʾ��։3�۝?i[?�<a����;)�ߐ¾��Խѱ>�[/�i/~����>D��텻���W��6��?�?MA�W�6��x�ۿ���[��{�C?"�>Y�>��>U�)�~�g�s%��1;>���>lR?!!�>��O?�<{?l�[?1cT>>�8��-���ә�'^3�Z�!>.@?.��?��?�y?�v�>��>��)�ྵU�����+�+Ⴞ�W=�Z>P��>z#�>�>{��=�Ƚ�O��`�>��L�=��b>���>l��>u�>2�w>�,�<�JG?S��>�r��"���ӟ�-y���Nq���t?kʏ?�M+?1=]o���G�O����-�>f�?�9�?�G,?��N�_��=�p��ڝ���1w�#޼>Hl�>u=�>���=�W`=�<>���>��>�L�9��8��#G�c?�wD?~��=oLɿ�i�M��S��F.��"	�7��J�F=�8��� ���e�����֌���Hh�%ʙ�a�ɾ6 �j篾T�
�/d?�*>ԃ������Y=yT��6q��p>f0�=.ʠ�P������5w��{�ĝ� (��-�<Q)d=V��=܉˾��}?�;I?R�+?:�C?��y>3?>X�3����>ʃ���@?�V>%�P�_���)�;�K���|����ؾYx׾��c�.ʟ�K>_I��>N83>�F�=�G�<V�=s=[��=��Q�U=m%�=�S�=g�=$��=��>�T>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�)7>h�>��R�:K1���Z���b��2Y�e�!?6o;�w�̾�>1�=t߾�=Ǿ��)=8@6>?Ke=Ձ��\�kS�=%k|��>=�Nl=X�>�E>���=Fų���=��E=�G�=�P>�{A�·0��0)���2=ʖ�=�sb>�=&>���>��?�`0?�Ld?.�>�%n��@Ͼ���C%�>�G�=�6�>$�=n�A>Sw�>��7?Z�D?��K?�Ų>���=���>I3�>O�,���m�r徢⧾X(�<���?nц?'��>�T<lA�f��Nc>�� Žr|?#S1?;y?�О>���ڿLk��O����;��O:��=NF��cM��
 ��!V�h���:>�ß>&|�>z��>��P>�T>]R>�>�>��>�ǧ=�8;aR�����%�x�tT�=!��jҼ�`���3=�
	��4-�WǊ��f������>e��삽��=���>е�����>
a�=����X�>IT<g�x��*=zt��G�A��+��+���[�C�ώ��~ �>�=>��������?RL>��H>���?� v?��s>T�M�=�f��j��C:��Y��'A>BU>Jd����;��KV�#�D��������>J�>��>%�l>F,��%?��0u=#I⾐B5�;��>ZZ��Ӆ����1q�6:�����Ui�g�Y�D?�<���Z�=��}?��I?ď?]g�>1(��=�ؾ��.>^��%�=P�Eap�]��r,?��&?���>+��E��l־��̽�4�>��P�Y�F�������,�C��<����,�>�Q��;έ.��s���q����C������Z�>lAR?���?�O�{���e�L�\��[�½_��>8d?�w�>��?�(?tL:���ᾄl����=P's?���?"�?���=ϥ�=���r�>~�
?��?H��?��s?5�B��Y�>�#�;((">���`�=5/>��=VD�=A�?�
?q	?`>���	������Z�c=L�=AD�>�P�>%&m>���=�Wm={C�=�tW>\{�>���>0�c>k�>� �>H������6��>!>�Ѻ>�@<?�ϟ>f��q3���Ľ?�=\Y˽�W��hA�.�o����<Ih=7A�=��<=��?��ֿ=z�?C
f>�3�PA?CO+����ㅏ>䖮>�����s�>�1>n��>�t>1ȅ>Ci?�ʇ>.;>?(��Nm=ya�$� �BD<�J��-��CZ�>�o����¾�7/��b�xoE�L����lg��s��?��k�<���?=����p���������>�a�>�*?�ɓ�����>$�?x+�>+ �
���e���L���?T�?&	|>�9�>|�X?~�?��e����~�y��hK��SY��1�(�J�������O���OS��5?F\?edX?T�(>u�A>�[�?%@��������>O�[�g�E�?�>�-�>���A����z;45�5i|��v>n�k?
�?�L?�*G��E��Tp�*�o?
ׄ?�;1?&�>�)�?�%��v ?�=>�1)?��}>�RD?�,?��j?L��>�N�> Fj= _O�1��#Ԟ�Ӄ�7�ཇP�;���J����:�������;I�>c��<#����z� z��w��]ݼ���<��=Z��>�e^?ݤ�>>�9?���s�9�MD��*;.?�Y=�i��ӌ��ħ������=��g?X�?\�]?
nl>D�A�d9��>�r�>7�+>�4Z>�H�>o�/�<��P�=�
>�>�6�=uD>�$��K�%㗾q��<��">���>�j|>,2��3�'>j��	z���d>��Q�����o�S� �G���1�Jv�+b�>��K?I�?��=�d�4e���Df�5 )?�Q<?WM?]�?'ѓ=e�۾��9���J�0�T�>a�<��'����"����:��:�s>X+���H��S�j>����^�+Og�4UI���쾜�a=�6��;5=����CѾ�>u�A�=\�>��=z!�������(�K?�"y=�ۧ�W��<���>eq�>ل�>��O�A�u��@��C���&�=s�>�D>?��(G���G��:��s>-H?��:?��x?���7.��l�A�:$Ҿ�о�j�x�?�ٖ>W?�� =�<F>O���Q>��o��A��!�>���>�/�	VT�7#ɾ�a�����e*>�"?'�>\�>��C?(<?[?�T9?6�#?�(S>��4����B(?m@�?c�ѻ�p,��Ԛ�Ͷ0�{kF����>G)1?{��us?>�~�>�3 ?M,<?Z`?�'?u���j2�ZN�t�>�m>������C {=�o?n��>?H?$�?��=�E������=�b�?yjh=O-p?��?p�>ZwM>h��>~������=Z��>��b?j�?w%p?���=g?(}1>m��>W��=Nz�>���>~9?��N?ɉs?pJ? ��>CA�<ͭ��������s�e�V���{;|j6<k�z=�����t�(\�h2�<�P�;�~������_d��{�F��N�����;O��>��l>)?��~t#>�2ɾ���� PH>}�}<���]�q�Wi��P�=��S>��>$rm>e.�4�=��>Pp�>m$*���+?G?�<?uL-=�d���Ͼ<)?��2�>� A?��=6o��|��D�t���w=H�k?��Y?sw����@�b?]?W��-�6�5"þi;��xL���E?@?W�G��y�>���?7s?�>�a��$Fo�v��=�_��{E��qL=�5�>@����V��A�>�42?�y�>�wt>��F=<�߾�Nq����F?��?5h�?�s�?ˏ:>��p���޿+žͧ�G�n?���>�y��=A?D3�<����)ﲾ�X��|7�0�x�<J�������Z���xn���������烼=��?	QK?ʑp?�'?���&�.��|�xk��,�\��%۾��5�AO��Ie��nK�p�W���پ�績��ҽ\��=8o}��A��_�? �)?*�-����>9菾�0��VMо_.>��������h�=���&�W=e�3= j��5-�@���?M��>7�>Ĥ9?��Z�2�:���.���5�����c�#>+��>.d�>3-�>,�8���8��=��ž�|�t��αh>|Z?eV6?��j?�e��g�:�����_���������̄>$�>�r�>�zo�F�
���'���;���o����>��'	�Q+�=�1?
ԉ>Nc�>� �?���>��&���1@?�~O<�4�W���>w?>��>���>���g�#��`?X�Z?"�>�ׂ>���R<�!�O�o�}�dk?���>-?�r{>��}(�Y���e��&rT�O~�>�Gr?�9���GݽO�>H�"?-X>O�����=��->�����(��%5�%��>y�?�6���}�=�����n!��!�}�.�,?K�%?��-�	F��6�=�Q#?�>��>�O�?af�>`!���I=�D�>Iy?�,A?r�p?n��>ns6=D�$�Ͳ.�4�z�|=(��>��T>9{=Z�=;���N��(��J�?>��?>�Q��ߜ�Ф=���>,u=�)�=�f�>�jۿh'K��_پi�U>��.
�����pҴ�x���k�QY��Ӂ���x�F���)��T���a� .���Sn�Sn�?� �?ޕ��-��
��f���z���>��o����ǘ���
��B����߾�ᬾ� !��$P��6i�@Je�kJ?���*|οj�U��M�{?�=�>�΄?U8ž�{	��_��)�>��>���?r�˹����Ŀ%o��!�?��>�0���� �?h��=F��=���>3�q��G����Ľ�7$?qA?�F�>%k�@�ǿ��¿���r#�?��@�|A?�(����YV=���>F�	?��?>�T1��I�S���mT�>U<�?���?�{M=+�W��	��e?<��F���ݻ��==;�=lE=���|�J>�U�>ɂ�}TA�#Bܽ��4>�م>@�"�b��"�^��|�<��]>��ս�9��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=s6�􉤻{���&V�}��=[��>c�>,������O��I��U��=�}�����
����#���=��@��ս��⦈:��=ڳ���_g���P�(=ma�=X�_>2��>��\>��>l%^?�Fj?NV�>�p�<�$�<l6�vvϾ�h���A���&�������Y���Ѿ@��NB��������/����J�g�=�	O�Z���=�c��~:�/3S�D+�>�}�>ˮ��N�r�+�=�㏾m�=�4)��}b��%8����*��?n��"�?%OO?%���(�l����=�	.�FX?��?��o��&�Jk>���=��R>��>G�v=��
���Q���&��/(?o�2?�‾�߼��>�|���	(<��O?��?��=vS�>�A?��M����Y�>�u�>5�>���>��>`�پQ-��gP ?��r? 9�<Dɾ؄�>g��"پ%<u��/�=S��n�s>�#�<���=M�����v��[k=G�W?>g�)�0������ELJ�$�;=ar?ø?pަ>��k?N�>?�<�<q#��U�(���I=i�Y?t�i?�>Im��8ʾ�����q4?#�`?�K>�}Y�.��k1������?��n?�]?��7S{�?��.��5?��v?�]^�}g�����:�V�@�>5��>A��>H�9�=_�>ĉ>?�B#��Z�����Nd4����?z�@ڑ�?tQ><����E�=�?w�>��N�r2ƾⲽ�����Ft=�[�>�6��ydv���-�+��f8?;��?���>�_�����2�=2A���L�?���?�԰�O+�<׺��:l�R� �Xx�<���=.J���;�/���:8��ƾ��i���{��&?�>�m@yL�����>�u2���Ώ�Ͽ���+)Ѿٿp��G?V�>��ཧh��~�i��]r��*D��E�í����>Ú>mט��&���{�><�������>&a��_z�>��R�이��]��͸.<B�>\��>|�>D¾��뾾���?:����cͿ�4���J	��Z?��?En�?�!?��<��{�${����� J?Ȯr?�R\?��/�dF`�i�H�.�y?��׾惿!h#�<Q�;%M>�r"?�_ ?[���C��`(�>E�"?z�=�"*�`��O���9Ծ-��?W��?8�]7 ?�ѐ??,��q^��͹3�Ŷ�Y�&�I?��> �e�`�_[��:�b�?w�Z?ĽZ�K�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?߮>�V|?W�J=b�>s9>>�ᾷ����">���=�꯽_R?|�F?c�	?�\�<v�+��3�i�B�ÂO��B�c�U�XF8>F�H?]|N?G��>�佰�ϼ���0E�(��'G=�ƫ�"�߽]�����>��Z>�*>�T^����*�?wp���ؿ7���4+��B5?�'�>��?G�6 w��N<���`?���>����ճ�yY��� ��B�?� �?��? �վ��ϼ7�>�>� }>�ͽ}ء��:����5>�OD?ۨ��㋿{�n��y�>=��?fz@�?wh�P	?b�*4��XA~��g���6��t�=D�7?.A���z>���>��=j�v�㻪�e�s�y��>HV�?U��?��>^�l?o�W=C� j-=b%�>	_k?h?��w��ֲC>�	?���㎿����e?�
@�t@Ŷ^?�Ӣ��hֿ����^N��Q�����=���=φ2>
�ٽ:_�= �7=��8�T=�����=r�>��d>"q>@(O>�a;>�)>���P�!�r��]���P�C�������Z�@��Xv�Yz��3�������?���3ý�x���Q�2&�*?`���=bR?�R?{�p?\ ?�rc��I(>� �$��<�k)�1�=�*�>Q-2?
 L?7D+?�3�=ꘜ�;c��À�\뤾Jƅ�-r�><E>Ȏ�>��>��>!��:�AB>31>59y>��>LS=�#���<�E>�t�>$1�>C�>NIH>E�T>���I���J�=���]��d��O��?�?��Y4�������-��TV���>��?��4>}+���̿�����rt?�����,��B�<.����\?S�S?��>�z��T�=�]>ea����m����=G@�.,e����6 >Z�,?��f>�*u>
�3��b8�e�P�3����Q|>o26?�ᶾTJ9��u�N�H��_ݾ�]M>�Ⱦ>I�B�Bl�����Z��qi���{=ww:?�}?h#���ް�ңu��6���OR>�C\>8!=�i�=eEM>_{c�X�ƽi�G�E�.=���=��^>�w?��*>T�k==t�>[��-S����>��'>�7>��E?�%?�Os�x���|��x4��c`>r��>���>pF>CWK�+��=�u�>i>3�.��ͮ�B?�01�mR>�����W���Y� ��=k����^�=��`=�s�t�H�IA@=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿl�>r~�][�������u�0$=���>[:H?�Q��ǼO�E>��w
?�?�Z򾀨����ȿ
|v�b��>�?���?��m��@���	@��|�>���?&hY?pi>�f۾�^Z�y��>�@?{	R?��><��'�S�?�޶?F��?�G>��?d�q?z`�>Ĭ^��#1���������/�]=�jN:sX�>_Y >gF���JF������(����j���$]>{,(=�J�>7��C����=�=/��4���Fae�Y��>T�o>�8B>[#�>z3 ?�r�>S��>��=6��Y큾�핾�O?:�?��ھ�����R�y>§��m�?�AX?�Z~����#�>��'?�Ҟ?�RS?�v?w�	�n���������c�< ��>��>�I�>o�o</[=>0/���8�te�>IH�>�`ƻa��v�u���$����>k=?^?;�>V�%?j0#?�G>�L�>O�ǽ��l�:��!�>���>J?u�?6
?�����8%��"��{ڣ�jb��>sY{?$?_��>|6��"4���o=�'��0���*�?��\?�:�1�?r.�?xwA?�.?��'>���X<�6[G�87~>��!?�P�4�A��`&��'�wu?'?���>�c��k�սm�ټ?��|���7?�\?wj&? ���#a��.þ���<�i"��@�
��;^C�)�>�x>Ꮗ�H�=��>8�=�m���6��Fa<Ǻ�=_}�>�#�=Qa6��̍�m�3?H.�ɯ��-"�=�My�B�=�g�k>��=U���#�y?NWཱུV��(���/����j����w?Mۻ? ��?INؼ�+b�V	8?[<�?2�?���>!BѾVľ7�¾�W~���O���(�=	��>��պ�M�涣��f������ۭ���S��|�>�l�>l?��>��)>l=�>CLD��uT�E-*� ��[���J=��C,���(��Ҁ������;�ξ][���a�>� �#�y> ��>��8>�ڇ>���>��-<P(_>�=g>!7�>�S�>��>�@A>��=��'<���LR?����&�'�.��񲰾93B?zqd?1�>|i�(�������?���?�r�?�;v>%h��,+�Yn?_?�>���7q
?�S:=
-�?�<�V�����*2������>�B׽� :��M�anf�Rj
?m/?T��O�̾T=׽H���r���A�?&?��9�N�A��Oq��Y��?V�x�3�r��������0)���t�N��vÁ�5X���b�[h=��(?�-�?���C���K��b
k���M�]%m>�
�>o��>�:�>l�(>����3��dY�lg��PE�M�>N�v?e&>�~`?lH?шJ?�@?w�/>�?�9m���f>#��<ʑ>���>1>Q?�r?3d\?��??�"[?[&-> �$�����Oƾ!!?�B?|��>��>1O4?'���L,�y���������޾쇼�9@>?�F>A�����=�v�=�s={W?x��r�8�b����k>�|7?u{�>M��>?���-��v\�<Q
�>ߴ
?$C�>2����}r�?c�QQ�>ՠ�?�����=��)>���=����<Cֺ�]�=�����ސ=�;���;��V<�z�=��=��q���|����:r�;s�< o?nv?��t=#��=�A��١�_I�YT���>��.?�	t>��&�ts��1�w�6q��n^>"�?Y��?�V>�AR>�Ӈ=HM��n8�N�#�I���0�>��>(�/?O�z?%�r?�v�>�=?�v�>�إ�渫�gӎ��~���� ?�&,?Y��>�����ʾ����#�3�Ė?!F?:(a�0b��+)�"�¾�ս��>�^/�5~������C�����q���K����?���?�>A���6��g�u���]Q���vC?B!�>i�>I�>��)�g�g��&���:>�d�>2	R?�	�>��O?� {?֦[?��T>��8��$��!Ù��;�0�!>�'@?ʟ�?��?C�x? �>&p>��)��3�	[��.���s�9Ȃ��5V=��Y>Jl�>g#�>�ة>:P�=:#Ƚ���o�>��=0b>Ӧ�>r��>p��>Cw>�u�<�C?���>�۵����O(����S��)�'�f?u�?
�"?�~=m,��j��V�If�>;L�?ܭ�?��E?GP%��>��=��w���!��>�=�>Ol�>y�
;�6?>܄�>rv�>�"�>�������]7�x����r?s�F?PJ�=����1x��b����@�/�!>��������E�TH?�H	'=eD���-��Њž�Ǽ��cW�1�s�ޢ��B;��F�վH�?�"�=�3X<Ȑ��d7�&	�53��
@=,��> >�>np�=]�>2<d�.|�=������=��a>�k>��ȼ���T�E?QP?��D?'@?��S>�M>�oM�����n�b���?�ˀ=�}��Tk˾3���^0¾Tp��Uʨ�}4��yg��j��:��=n���|>^��=�\�=QM�����<���=�ئ=�P��@:Z�"=1;>�I�=��=&h�=w�>�6w?K�������4Q�Z罠�:?�8�>�z�=N�ƾ�@?��>>�2������rb��-?x��?�T�?d�?	ti��d�>H��n䎽�q�=ظ���=2>���=�2����>v�J>��� K��C����4�?��@f�??�ዿ��Ͽ*a/>��2>�>P\P�p*�SF����)e���?�=��f̾_��>ܸ�=�پ�3ɾ/�V=a�$>z�!=J�)�j"[��n�=�~F�VOL=��D=5��>.�3>1��=����2$�=dJF=&��=8�L>�m��^������TH=���=6S>W�">d��>2�?d0?�Wd? 0�>��m��Ͼ�E��>�>���=�B�>kم=�fB>���>\�7?�D?9�K?%��> ��={�>[�>/�,���m��k徎Ƨ�Ļ�<@��?ʆ??ȸ>x6Q<F�A�����h>�FUŽ�q?�Q1?	m?��>�U��߿��$���-����;�"���=lr��A�POӼ�c����N�=d��>.��>ĩ�>�~>�-:>WfF>���>|2>w-�< �Z=�$����<�Ͼ�4j�=�黠�=A����J; | :2k�͈ļ�U <�6�;�˒<@c�;>�=���>�bѻô>�G6>�꾋��>�y�G7o�s|�=�$/��0�"�]�����~�M�yH����w>:�J>z�Y=ת��}�>o�>į�>��?�1f?v>Y���?]�4�����������VL>�ug=�ӽ�3���^�C�G�����>�r�>Z�>�c>8$�ƐF�x�F;lXξml*���>�Y�<k=�E��Z�m�����Dŝ��e�����.B?O���.�=�Eo?�qL?2�?�"�>�u��Ǹ��ڞ=]x��oD=�����E�R��LL3?��$?N�>���e�S�9vʾwʽ&Ը>6H��oQ�����x�1�[R=����\%�>M.��A�о(�4�F����ޏ�+�A��q�Ї�>��O?�K�?YpT���
�O���N���� ?��g?��>)�?]�?�����'��{���b�=��o?(c�?ɚ�?�>w�=r������>�7
?��?���?%�s?�!E����>`�麯3!>	����|�=<�>���=h]�=1�?<�	?�k	?���]��t�p%��`����<�j�=��>狇>��m>���=��_=	��=%3W>��>>�>�Vd>|D�>�Љ>V���a6�>٫%>qRg>X�?攫>,�>�׽� �����U�=Ƚ��Q�Ԣx�:���N���t-$=�\j=�G?���yî?D�6>;xE�;7?$�l鍾�)�>��>++���N�>t>�Rx>or�>;��>���;��^>�T>�Ͼ&>����"��oB��xN���Ҿ�S�>���"\$�޻
�e��#A��Ұ�
���$h�'��@">��h�<�Ր?�]
�7�k��P&�_����
?��>*6?ca���y����>g��>�6�>���Ǜ��4���	�ྺ��?���?�~>�=>�L?8S?2=��Ǫ����v�U\�e1I��]S�εh����/����+���M���O?G�q?iMY?*��=��u>��?m\�<�;�,?Z0�6�B�@$>w��>_,����x<2������ɽ���=�ք?o9�?�EB?�u?�i�o��g�� |?�dn?
�W?bR?�:�?CYƾ�:h>uS�=��#?W�=�%?��@?6�M?�#>��y>��ܽ��~����箌��˽g7�l{��.�=�S��=J�����҅=�l�=�>�����6G?��"?��ԽM��<�=� �>��]?Xh�>��>��6?G��Q+8����?�/?4�A=�����磾.���>Ük?�˫?�Y?Zc>qAC�a�B��>O��>9F'>��Y>��>�콥H�B�=z>K0>���=34\����̇	�s�����<5�!>���>>|>E썽/�'> t��9)z���d>o�Q�Wɺ�t�S���G���1�erv��V�>��K?��?֪�=�\��)��EHf�-)?�Z<?ZRM?/�?���=��۾v�9���J�DG���>�<$��׾��� ���:��h�:|�s>�0��5�����q>l{�����eE]��sQ�����=�H��( �����ݴ�rox�V~=��>�󪾹2#��ɕ��I���~N?̪=�f���.}�J����- >Ax�>���>Ǫ�f����L��̱�i��=#/�>/�>!�Ƽ���H�l��{>��9?��h?�Ջ?������cN��,⾹��*Q̽=K)?偼>��?�J7<u�=B몾����o�]W��!�>\��>3,�w�[�h���*Q��L���f�>(�?.��>'u]>λ\?0O�>��}?0�A?/:>?c�>����ľۼ+?�w?�>k�6�Z����"��Z��)?�?��وٽT-?+?��-?�,Q?��+?*k�=I�;���V��p�>��>��H�ſ;E>�c?e~�>Pe?��?/��>�a��6��'�����>y�0>��X?@�>"?��>,��>tK����=��>�(d?^�?�mp?x��=�f?c{->�"�>ĝ=R��>��>^r?eO?w�s?�J?m��>��<
c��#ܺ��@f�sV$��ĉ;��3<*(�=��bDs��6��#=%��;��ԼcY��!��-G�5ґ���<$b�>�s>�����0>��ľ�n��3�@>(���_^���Ȋ��J:�F�=I{�>7�?ڍ�>�#����=H��>�S�>���a6(?��?I?�2.;�b�r�ھ��K���>�
B?Q�=
�l�������u�ZBh=]�m?��^?��W��:���b?��]?1f�=���þ¸b�����O?:�
?b�G�>�>��~?�q?k��>��e��8n����Eb���j�Uض=r�>{X��d�V=�> �7?�L�>�b>)0�=
s۾��w�jp���?��?��?6��?F**>K�n��3࿚D׾�/���#~?���>����
�0?3ѭ<9ɾ~舾�S]�$�ؾ�/��י��d��'���l6��X��Wɠ��Q�=
a?�n?�s?<�B?���@NU��i���q��iBM�3��!�+v4��O�rkM�{f�!C�B�����z��]>��x��iD��Ŷ?��(?zK��6�>2Y��m�J�ʾ�<E>�ќ���
�U��=Nۏ��#=�?=Ghn�TH(�W!��4r!?�δ>���>�9?��\�9�9�b�8�E�:���=>>$B�>5��>���>h�_�ٽ+���Ͻ�Jξ	����!���Df>!�V?� F?�v?��>���:���x�����
��G�!˅>?w�=c�t>�.ʾ�-���6�|�5�� _����a���	��V>0D?ё�>��h>�[t?U?4:��{ľ꩸�7�'���>���>�vh?L0�>|�>����U����>�Fo?���>��>f�ھ6��u��7׾��7?hz�>���>�����5��4?'�]�r���	,R��^�>7i�?/k��}���^{�>v�h?��e�b���V�>�ߟ>�<6�&�;�1ڽs��>y��>��q�XŇ>-����U��y���t�]<-?$�1?�a�s<;��I>�GS?Ab?aL�/"?�]S?��@�"n��+?�ׇ?�*S?�pM?r!
?�Lb�tYξ�b����&��� �2]�>���>����>����냾!�	��h>��>z�>F���b(=�,f�<�>*�<,T><Uؿ�AI�3�ھi �g�۾,J�BZ��[����Ib���'�z��� ܃��ye�>�(�샴�r�3�5[b�c^��|�m�0��?���?�։�iO�����/>z�����u��>R�d�ʛ������꽳���&龷����jM�B�e��|b��<?2��/Gؿ�`����¾f�M?s5�>��?6ʾy� �S�4�>c��>����,nվ�B���οپ��j�G?�>����ʽ���>�=��B��=���>:�ܾ�����襽5R�>�O'?�1�>��̾.9�s~׿k.�62�?��@�|A?3�(����8 V=���>ԑ	?�?>|Y1�vI�����EU�>�;�?o��?�M=n�W��	���e?"O<�F��ݻ��=S3�=�c=w��e�J>lX�>���MRA�RFܽʶ4>�څ>�`"�_�� �^����<��]>��ս�7��Մ?�x\��f�y�/�U��o\>q�T?r*�>�<�=ͳ,?�7H�^}Ͽ�\�},a?80�?���?W�(?�ڿ�eԚ>�ܾ4�M?C6?���>�c&���t�ؖ�=*�ἄ6��@�㾑#V�W��=w��>{�>��,�ƌ���O��!��H��=}B���o��-&��� ���>���
8	��읽y��=ʫ:�jʾʙ��3��:L5Q>�$�>��i>:g>�+Q>�~c?j�?0�>�#=�*�wc���p޾�=]߽x�O�L�����!=D�}���6>�ɝξ�R%��'�����$2�BY�=TaD��Ȍ��Y��m� V?��G1?�[�>L������>>q>���߾��u=ߟ=��׾�&8�Z�b�?�	M?>�l��`�`������_���<pK?�u@���Ͼﭸ�mD8=������=�%>*Pٻ����N,�KC�ds0?�f?Ք���F����*>�� �7�=��+?�d?�"m<3�>�7%? y)�����[>>%4>�;�>tq�>_[>�����۽~?x�T?)���)��D�>�k���Pz�	:\=I>�c5����M[>>i�<��eS��b���X�<(W?��>��)����Z��ӷ��==p�x?0�?44�>yk?-�B?���<�d���S����kw=E�W?�)i?u�>����о5~���5?�e?D�N>�dh���龰�.��S��"?��n?_?Ψ��Ww}����x���n6?��v?�r^�_s�������V�j=�>x[�>���>��9��k�>�>?�#��G�������Y4�Þ?z�@���?��;<��휎=o;?\�>��O�w>ƾ�z�������q=�"�>ǌ���ev����iQ,�N�8?Ġ�?Ŕ�>˓��������=����g��?[7�?�ż�z�< ����h�����<~`�=sż0G����n�7�! ƾ�M�v����	y��܈>��@A��h��>�}����8�ҿ�����;��}�9\?*8�>y��AV����l�H�l�H	A��J?�4x� -�>��>���>T���{���;���ҼT��>e5��z�>�"Y�r��������;<! �>UU�>H�>vǽQ������?0n��O�Ϳoߟ�,��wY?v�?pą?!?́�<B���T�w��ʇ�d�I?�ys?\?۫#�,�_���8���m?�#��P��'�� �r����<x�4?z}�>�h#� �Z��9@>�?cc>�<��ɿ�ſ�i"� ՛?��?e� ��
?�U�?��,?���A��͟������5�t�^?7!�>�4ľ_�F���8�	�̾�?bG]?{�ֽ���]�_?�a�=�p���-���ƽ�ۡ>�0��e\�uM������Xe���Ay����?F^�?g�?е�� #�J6%?�>O����8Ǿ��<���>�(�>Z*N>J_�a�u>����:��h	>���?�~�?Lj?��������V> �}?��>�?��=��>���=�F��ϟ8�!#>���=M�C�[�?YbM?#%�>S��=f9��</��AF�}&R�Y$���C���>(�a?4�L?��c>j��F5�P� �Pн�`1���dh@��@(�x�޽��5>�C>>s�>`E���Ӿ��?Hp�9�ؿ�i��dp'��54?9��>�?����t�����;_?Nz�>�6�,���%���B�]��?�G�?2�?��׾%Q̼ >5�>�I�>��Խ����l����7>8�B?e��D��r�o�f�>���?
�@�ծ?ji��	?���P��<a~���y7����=��7?j0���z>���>��=Hov�ֻ��e�s����>�B�?�{�?K��>��l?5�o�v�B���1=�M�>ʜk?�s?ϱo����B>��?d�������K��f?��
@wu@|�^?
ܿԎ�����+�q�e!8=�	�=�c>*��%��4E=,��IQ��m�=�<�>\��>�q�>'�>�>�>FN>Ѯ���Q ��㡿�>��s��CW���J逾_���[�a������־^0뾒꛼� H=�N����c8����<Z}�=ةU?x�Q?`�o?� ?`�w�� >H����(=FY"�?�=��>Ù2?r�L?��*?y	�=s��7�d��_���I��������>�UJ>�E�>���>�E�>�#	���I>>>�f�>�� >N�'=�*��=}�N>^�>��>���>6 e>$�Q>���e��f�)���K��>K�/��?z_^�}�F��Ǚ�����,0v=/9#?�F>���� ͿW���!X?�3��v3�}���=|�=86\?9=?��>v��n9�<Dc>��̽���b>�ݲ�����5�%��ׁ>��?<Pj>U2y>2��u9�clQ�� ��m�x>��5?ʖ��,!/�Џv�m�I��q޾\�X>~��>z��ҳ��c�����K;i�-D�=��8?��?j粽b쬾7ei�H����0K>-�`>�iD=�֜=jnO>3kb��~Ľ��N��u?=C{�=�l^> Z?�=,>�l�=(��>���w�O�F��>��A>?;,>$*@?$ %?�9ؖ�F����-�%w>w�>I%�>�>QfJ���=,t�>�Fb>� �Z��JQ���?��W>~���e_�5gu��y=��h��=u��=� ���<�F�&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾRh�>|x��Z�������u���#=Q��>�8H?�V����O�f>��v
?�?�^�੤���ȿ6|v����>X�?���?g�m��A���@����>9��?�gY?koi>�g۾=`Z����>һ@?�R?�>�9���'���?�޶?ׯ�?CiF>�k�?e�s?fQ�>�\�e\0�唳��7���8@=�zB��\�> �=�ļ��IH�af���_��t�h������T>w
=��>�Ͻ�綾��=CA��V����-]���>h�u>�N>�{�>,z?���>��>_�C=�������֜�&7N?��?QܾQ1���Ƚ��^>.���WW	?�d2?�"1>�M��zT>�&?\֓?�V?o��>����������댣�M��=�>9Y�>�ܶ>́�=j��>�/�[pi���>� �>�}�u��٩��,���>o�?wC?�ɀ=� ?3�#?��j>&�>jaE��8����E����>5��>I?��~?��?Aֹ��X3�����桿F�[�UBN>�x?�T?-ɕ>?���.�����E�O`I���㜂?�rg?�e�C?3�?`�??K�A?�(f>���ؾ������>>�"?�k�k�=�<�(����s�
?��?Y��>Z,��Aˬ�YH�?������>?��[?q(?Rv��`��ʾ���<��f�ƙ��`�;wb���'>9/>����B�=�t&>�l�=X�}�9�0�fX�<1�=��>��=(�"����0=,?��G�{ۃ���={�r�1xD�s�>�IL>����^?Zl=��{�����x��=	U�� �?���?^k�?(��9�h��$=?�?L	?e"�>�J���}޾>�ྡPw��}x��w�?�>���>:�l���I���י���F��S�Ž��F� <�>�%�> ?B�?���=�~ ?p�����h�}��dX�� W�p�:��7��=G���@�����7�k�g6ֽ(8���쇾J��>��C�BΒ>!�?\�>��w>k��>D֒��.,>} h>�A�>�{�>=��>��/>X��=�)=}d��KR?����$�'����²��g3B?�qd?Q1�>ii�;��������?���?Ts�?=v>h��,+��n?�>�>H��Wq
?}T:=�8�
;�<V��u��3���1��>E׽� :��M�Dnf�vj
?�/?
����̾�;׽)����۷<�?H�'?42:�6y?�'�i���K�MeL��gּ�V��2���t�&���q�9�����z�}���v����=F�%?0��?�������W���o���_�?um>fZ�>�W>+ե>�>�G$��3�$
f�V��6�2?��z?09�>��.?u~@?}�p?�v?=c>�8? ��uK�>�E>��>T%�>5�k?тF?/�]?!�7?��?�,>�`��s������P?�7:?���>��>�\�>G�Q��Vq�~�x�#Ʃ��`�'@X��#=�y�>M:ʻ+=���=��>�X?�����8�����k>5�7?|�>c��>_��O)��F�<V�>}�
?�F�>� ��}r�/b��Z�>q��?����=��)>i��=�����}Ժ�^�=B���O�=8���x;�!p<�=���=h�t��݊����:r�;���<��?Ȃ$?u1�>p�3>�.=�)sǾ�����"�x�>��>��>?��<~��
Q����j��sX>"k�?�w�?Q��=K��=hx>�+��/���s9��f��_&=���>q�'?�MS?���?Gf'?��+?�
8>G_�B������R���D?�#,?���>���ٲʾP��3�ڜ?�\?�8a����9)��¾�Խ>�_/��5~�	���D� ���\���m����?��?3~A���6��d�����q`����C?d"�>�T�>w�>t�)���g��%�;;>���>7R?��>k�O?|:{?��[?�|T>��8� ,���Ι�+�6���!>�"@?ի�?%�?sy?�n�>!�>��)�K�4a��F�����ւ�k?W=�"Z>�~�><�>��>գ�=�ǽ�C����>��ʥ=��b>�>���>��>&Ew>�&�<��G?���>Ѣ�����S���Pa{�fHn���p?���?��+?s��<�Z�uI�+����p�>GB�?���?��,?�P���=ܨ���w��ex��'�>�#�>'>�?=k�]=�)>@i�>g@�>��	���x6���l�k�?GzF?���=uÿ��j���s��B����<�5���Gr�O�D��1�M(=)�����ڽ|f��-w� ɓ��o���|��������|��-?�]�=�)�=��y=L��9w�̷<	8i=��<�g�<�,�\�J<PRz����i>���r��N���(�$=6���s˾X6}?��H?��+?��C?S�x>�:>=70�c��>�"���t?�fT>�NX�켾��<�Μ��g����ؾ��׾��c�ڨ��"A	>��H�5><%3>�\�=~3�<~��=% s=ң�=5p��� =�Z�=L�=�<�=�)�=џ>s>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��4>�s>�_R���1��5\��$e���[���!?(�9���;�U�>�'�=��޾-�Ǿ�O4=�7>�,\=J9���[����=dk�95=j�Y=e��>�]B>T�=Ȋ�����=�lJ=��=C|M>��ƻ��0��<4�J�'=���=.�`>,�#>��>��?4a0?�Ud?'5�>�n�_Ͼ@��G�>�%�=�D�>��=�oB>/��>��7?I�D?��K?���>���=��>��>;�,�3�m�Oh�̧����<N��?�͆?iѸ>�Q<J�A����f>�[.Ž�v?UT1?;k?��>�u��c�Qe�Z3վ���=����E�d=}L��Y�&P5�()E�m����=$ִ>G?�1�>��>�:>��>��>��>>�Xc�݄һ98�=(���?�P�=,E>��;})5��"��/�����`��w�;�X4�1{;\c=���=�m�>��=�m�>'��=���vq�>��*���t��$�=̰ӽ�02��f�r����C�mՕ���/>Q>&�R�b���CP�>��|>�m>���?/&�?��4>��&���辽?��ׁ��^1����)�
\H>Tu��_,�BI�\L�X����H�>ʦ�>�P\>z�}>��1��?b�M�>AϘ��H��?�> �ԯ=Ʋ@�Ȣ������ߠ��JT��;8�D?-���l� >�~}?(}I?vQ�?���>��K������B�ӫp�,8�=w*�;ّ��㲽H�?@Q)?�?�Y��Da���Ǿ����QR�> MD�#cP�󚔿�W1���[����O�>�J����;el4�y��i쏿��@�*�u��ü>6�P?��?�pI�������P��)�^�����>#�e?R��>�?��?�Ƿ��1��^]���+�=�n?v��?tf�?G>���=-q���E�>�=	?�Ö?s��?Ĉs?�a?�5X�>p�;�� >�p�����=+�>�М=�9�=�t?i�
?��
?�"��c�	�'�����]�,�<���=<��>Ԗ�>��r>��=�i=J7�=@�[>���>�ۏ>X�d>���>VQ�>�㝾\�!�)?�ł>S�->�?=��>��E>ԯ�Ů~����=F\ҽ羥�!����Z���	���;�)=&����>��οĦ?�+>�C�<�)?	+�̆<��|�>�2�>�R�[0�>�Ŕ>��f>��>���>�<l��>��>
?Ӿ�>����f!�0)C�G}R�=�ѾQ�z>����%&�M��c���8I�%k���c�,j��.���<=�4b�<�G�?�����k�s�)�<����?e^�>Q6?�،������>���>]ˍ>�I��$����ʍ��c���?��?[Ñ>ｫ>P�Q?���>�z����o���X�E��;LF���T�sz��qY����l���jF?��S?{c?f�K>�;o>A)�?�T�y:�{��>>_�O%D�}����>&�i��z��k�����w�b8�=yW?���?9>?�
x�m�P���6<��>?T�R?K�?��0?�LM?��ͽh^?��=��>
�?Ͽ6?��&?\�?��Y>=.>d�<��V<��� Q����
�
ڮ<��j=�$";wJy=�c�=o�n=�h�<� �=�<;��������Ws<�D<��=�I�=�>,�b?�F�>VM�$�B?/�=��U��4��yR?�t>��;�Z�'�˃����ξ>R��f�1?���?'͍?�ˢ>z�Jνtƶ=5�/>:��=��x>��>3冾�/3��c:>��>��#=���>�\�=~f�sk$��*־�Q =%7>�2�>�}>�T��f�$>@^��нv���c>�Q�b��ҊP��'H��K2�r�w��	�>!�K??@�=�8龀ߛ���e�' )?��;?|M?nf?Vg�=z�پi�:���J�=����>��<8h��}��9ϡ�_;��+2;�hu>ۯ�������72>���q%�dX��8��8�i6������=��
�������I�=��=���#�(�_����Ȧ���F?���=W-��:{G�ق��t>��>��>��8�|½�D�q譾�8�=��>9�<>�����|�8��Ǿwl�>W�E?O�^?v��?�R��w�r��mC��a���R���|��K?Z��>��?�fC>7�=K@���j�ӧd���F��}�>�j�>9���9I�����E
龾#��,�>��?y�>?GtQ?�e?��`?�**?r4?��>�ý�Z���$?Pd�?��&=�=�z����Q�B�m��>F6 ?!��>�>]N?��(?Y�.?�[O?ޅ?N�=iQ�=Q��i�>^̉>��\�oݰ��eb>$[Z?���>��D?]h? �o>s��k�%W�=L�>��3>ޗ2?�?@<?@�>��>�q��?�=�`�>|�b?� �?l�o?p%�=D?Z�1>/��>ބ�=�ܟ>`��>�6?NO?�s??�J?��>0��<�r�������s�m%U�BO{;��I<!{=�����r�������<��;Mֵ�N���8Z���C��������;z�>x�r>ˀ���:4>Qrž�h����A>�G���F��L���!�9�p��=�~�>�� ?���>������=�W�>�%�>����(?��?�?�?=;²b�u|ܾX9J����>�JA?�C�=�ul�􂔿�5u�/�l=�l?_�]?�V�5s����U?�%e?OOȾ�%���Ծ�P�7���`B?-�?��о���>z�O?�8^?D� ?�_4�4�V�MT���<c������>o��>L�<�.Q|�Z��>�u?N4�>/f>���L^�;W�"�R��l"?'Ό?J�?:��?j�V>X6q��⿧0��������]?�X�>���6�!?P]���ξ�ދ�IZ�����#�|�����͠�!'���t�t8н�؞=�?*�r?��o?5�\?J�����`�cSZ�=瀿��V����R"��@H�F6D�0�@��0n�������㕾��+=�A��U;A���?�q&?��/�x�>}����e��;�A>')������ь=X��>fC=�S=f�y-0�&`����?��>�M�>��;?�Z��=�b�1�u38��[��˜3>W��>+ɑ>j��>��o;-0��=佦�Ǿ�'���ӽr�k>]Uj?\�R?�ju?F�9���S�xކ���y>8ª��>��=Au>� �͙�ܗ%��C��)c�:�Ծ��^���(췼�?��>R�?=�?q
?�V����p�	%J�=�=>̾>�!J?�� ?v�>�o��jX�3��>I�t?��>��P>\��E�O���_���3>���>��?WR?ՎK>��)���/���pH��3�C��&6>�m�?�n�26f�f��>�Vx?�RC=�(%;�Ɩ>mR������k������1�>���>3ҭ<;��>e�>�
���)ϥ�!�"?*�!?�2r� =8�{l>�(%?��?K�>�5?�G>'T[���,>�S5?�g?��H?|<?��>�ڼ�����~��2��U�=R�>i�>c;�
y>�׽�������\���D>d��ʼ��#=,T��q�
���=��>ilۿ��L��ɾΛ��p�a����Vj�J!�#E��!$�*Ҿ����m����D���4� �V��@���o��#|����?��?o��=ܞ�k���x�y�����e�>�����:��pN���8�]��������
�������M��c���p���?kڠ�t�ÿ��ċ��),?�S?e�{?ߤ2�&o��X�Ӄ6< ����>~pо�Z����ƿ�#ž)�k?1	?� �zѾ躐>�W�=�^�=}
E=�%e��<��o>|�?%Rk?0�2?��ǽ��ÿ�v���d�=��?S@ȜM?�7���
�š>[��>� ?�ޝ>�	��G:*�s�W�V��>8�?Z�?Ƴ�H�S�G�	>L	p?�'�=/C����eb>Q�>�8�=��p��k>VL�>Oh��ݏ<���">�>.&=�����!�Qa�<o�x>�u߽����5Մ?*{\��f���/��T��$U>��T?�*�>W:�=��,?U7H�[}Ͽ�\��*a?�0�?���?-�(?$ۿ��ؚ>��ܾ��M?\D6?���>�d&��t����=�5�"���x���&V�m��=E��>_�>��,������O��I��T��=�4���¿ɦ����=,�v= g���7�D�ܽC��+̾8���q��4W�=X��=@�6> �F>�>��D>�W?�5q?�ܹ>C L=<�� /��G����3����� �jH���-��ɾ�Xg��.����|E��K辿>=�<��=8�Q��k��B��yb�]F��.?��!>��ʾr�M�#��;^�˾���0���e���B�;cu2�A�m�脟?H`A?���o'V�Ap�'�F]��#�X?����K��@����=�P��DO=E��>$�=;��I,2�ԴQ�{a?մ?DNɾ�
R��'�>6Խ�[�`M"?Gi�>Ia�����>��/?!N,�����N(>�J>��>���>�˼�����!�N�9?�1?|��m޾Psy>�WO�Ԝ<�2�`�ľ�=3�9�t>Ͻ�e�>�h>���͆,��(��&�=�Q?��>P���^0�Уݾ��-���7�<�?�~?�{�>"�r?�/?�y��dӾ	`c� ����<�gZ?��b?��>��T�_%Ҿ9�i��{?(1V?^�>VMO� �����z)����
?76i?��?���<�����n��[��'�@?�
�?��������;2<�\�˼�c�>�B ?�7�<��o�hя>��2?�
�=�6��$���|2�d��?���?p�?���Gۓ��P%>}�>�\?���� �!=�1���"'>��?�׾y n�}R��{�оɺ?�#�?���>iU������=dٕ��Z�?)�?����Y;g<����l�Sn��Nv�<�̫=���Y"����|�7�/�ƾ[�
��������c��>2Z@�T��*�>{D8� 6⿼SϿ�� \оMTq��?�}�>�ȽD����j�;Ou���G�h�H�ݤ�����>w>Jt���M��}�z��:��Ѽ�\�>�G� ��>�nO��Ӹ��m����b</$�>��>��>&
��PB��Z=�?OX����ο�Ҟ�ݓ��X\?��?�6�?�k?�H����v�\nz�ET���pG?�+s?2Z?�0�C�a�9�g���j?/b��rV`���4��DE�'U>�!3?C�>�-���|={">��>e>�"/��Ŀ�ض�S���?��?���?Fm����>���?�u+?i�i7�� [����*���-�8;A?�2>6����!�2=�fВ�J�
?O~0?�x�</�]�_?*�a�M�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>hH_���u>����:�	i	>���?�~�?Pj?���� ����U>
�}?�>ō�?O�6>t4?7z�����+n�	�>�]�>�>�?��I?��>�=N趽{*D��K��pD�8�W��1@��Qu>�j?�M?���>�����-���<�A��/��� g�=^��xa��D���>���>r��=o�y���ݾb�6?B�6�Hyݿ[��.)#>��-?�h>0�-?��&��c��>1��?���>9"��O����:���>a��?�~�?@�?�^	�Wǽ=q��>\��>�eH>�󽹉��*��d�e1U?q&�<L���E���I>���?�@���?ǜ^�iK	?y]�Vd��{~����M6���=�7?��U�y>�&�>X�=T7v������s��r�>�T�?l�?��>��l?Ďo�P�B�J�:=�ѣ>�>k?�@?�ٷ���dB>��?���p玿ø���e?�
@�Y@j�^?X�A=տ���[�P�~,����=A�>>�>��c�,k=ț���ro�wR���=pO�>(;>�*0>4��=��=��=V����b#��虿gy��R�2��y��A�����7�E�� �e���5�پ���cv�	�)�a��f���������=�=W?8�R?A�d?u?��e�<l">|����=����)�=�i�>��2?�FK?��@? ��=�:��؇]�1�}��T�������>Ǿ0>KB�>>	�>]�>�LǼ�i>�.K>[�e>���=Б�~q/��͍=�R>���>���>���>Y�=kL�=�x��p����1�'�O=r=ym�?�;۾�S�}������>�Ak>F�?~�B=���uϿ�͘��K?�ؑ��`3��D��B>{�H?u�?}w�>c����V��\�;��B�)wV�*�\>�`��Jn��2���~>�w,?��d>t7t>7H3��e8�[�P�Iﯾ��|>�5?n����j9���u�I�H�L޾��L>恾>��J��r�]���>�ZNh���}=:;:?i,?ؘ��e�kw��T����R>H�\>ׯ=���=��M>�X^��ǽ��G��.=���=��^>��?$n>�(�=%!�>����44��Q�>UB/>��">�=?��?�kd�p�ܽ%7���`�	�~>��>2S�>GX�=	�H��,�=6;�>��d>��T���|�)�Y��U>�n���1~������V<�e��D��=��=㴸�1�0�*=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿl��>�:�����Ƌ��@c� @�=���>��M?w ����<d�c�Η?��?�B��M���gпZPs�bA�>?��?��?�i������I3�� �>o2�?��,?�ԃ>�j��c3�I��>�T?7�c?�P�>ާ(���V��V+?-u�?z?�hH>��?V�s? ��>����93�W��~ߋ���=�M><��>�;>a��j�C��3���6��:=k����t_o>�~=p�>�DԽg��n��=�Jy��A��"1Z����>�[>��J>Iߔ>M� ?*��>���>j02=ˊ����}�����'dE?[đ?O	�~s��3��S?>���^��>�+?1��Gj�1��>Cw?pU�?��U?�9�>Z�
������������2a�<�PK>b�>P��>돽��>�-����Ѐ�>.�y>V{�=n��H�P��h&<o��>:Q?��>��O>�= ?�J%?Gj>�8�>�I�6���E�d��>�:�> �?2�?�!?K���20�nؓ��Ƞ��X��Y>~�v?D.?뺔>~������,����:�~]���?�c? ɽ��?gI�?�*@?|�C?Mtb>��)��-����Ț�>i�!?����A��c&�h4��?�I?z��>?�����׽c�μ��������?L!\?�;&?����&a�@þ+a�<�� ���U���;u=���>�>ɵ���ƴ=�>�w�=�/l�_a5��,k<��=Rv�>X��=�R6��i��vB1?4�Ƽ��l��>�Gs��q��ls>{�g=H����-m?Og�\�U�����%I����e���?���?�h�?�
��:p�9�f?��p?���>-?� ̾I+��Z��e� �8y���ež��>q�?>ʎܽ�V��֠��룿G�h�2 ���	��>���>S�?�� ?u�O>?��>�Ř���&�I�����\�]�|d�~�8�;�.�
^�u|���!�u��>¾��{�fL�>�[���n�>�	?�ig>1}>��>W���mE�>��Q>c�}>�M�>�Y>n3>�f >���;8�ν5R?���~�'���辐��B?�d?D=�>%�e��z���g�1�?3��?My�?��v>�h�-+�� ?n�>�9���$
?i�?=���ۘ<s����]��������>Tٽ	:��$M��hf���
?�?�}���*̾��׽	����hn=�F�?h�(?��)���Q��o���W��S���/h�����$��p�p㏿�V���"����(�R�(=@�*?W�?2����} ���k��!?��kf>��>�"�>�Ͼ>�I>��	���1���]��?'�𻃾�(�>;V{?�>KiS?I|:?�@!?�-f?D1~>ɸ�>��r��?<ù���>�	?`H?�H>?yun? "?��>ɱ�=(���P��{ݾ�5?Z?k?ps�>�g�>ɒ�`�;dFh=��=N��_T�4���R%�>�9���7�=��	>ZW?U���8�I%���j>��7?���>���>˻��i�����<���>�?}��>����<,r��c����>L��?�~�v�=j*>��=�lw��l ����=|���=��y��<=��](<y%�=�z�=.a��e����:*�;�}�<���>�	6?˲�>���<޾�=���M����>=�>��>���=J��; ��b䍿�}|�*R�>��?�(�?7��=�c&>& >�kξ�H��$�i0����O>ɖ6?a�??�>|?
�?�O?>�?�h�>�?	����� ���\��?Q,?��>����ʾ�����3�Պ?�r?�a�P���#)�zp¾Rս��>bB/�{M~� ����C��%M��������.��?xɝ?�>� �6����;ɘ�䫾!pC?���>�o�>���>�)��g�k��5;>��>��Q?�w�>X�P?(_{?�\?�G>�\=�W������u8<�t)>�8A?S؀?�B�?T�v?���>F>�O6��Y�K��&�N���z�=O=��`>�(�>��>ܩ>(��=d_��������O�$ܯ=Q.f>S��>���>���>��u>��D:F�G?E��>z�����Rɤ�Z���U?���u?��?�x+?�=�]�gF�;P���R�>�T�?���?�,*?�T���=/ּR}���q���>;Ϲ>��>i	�=��D=�2>&��>	3�>��@F�2t8��lL��	?#F?o�=;�Կ ��Ojλ��<�~�:�G�� ��)羒����;���'��U��!��=S��ʓ��-��|%��\-#��1�%��>5�H>�7�����EK�=d&z;C7�!��=�l�<�����-�	�&={�l�t�<2lȽ�3	<���;�#p�5�<[�˾��}?\=I?��+?9�C?y�y>�>>\�3���>~���??�V>�xP�����};���������ؾft׾v�c��˟��E>�MI���>t23>�6�==�<X�=(s=�ю=�}Q�4=�%�=>L�=�f�=/��=e�>�Q>�6w?_�������4Q�/Z罨�:?�8�>1z�=ہƾ`@?��>>�2�������b��-?���?�T�?T�?[ti��d�>!��j㎽�q�=东�G>2>n��=��2�[��>�J>����J�����m4�?��@��??�ዿǢϿ�`/>a�7>{�>aHQ��%1��XZ��\a�}�]��<!?��:�@�˾=��>�=S��}6ǾK�4=��4>&1s=4,�z\���=��y�`�N=+En=)�>+C>���=�Z��n$�=�D=C��=�J>^�#@.�I4��[6=���=n�a>P%>Y��>��? d0?Bd?F�><�m�IϾ�1��x^�>��=(1�>x؅=DB>s�>R
8?Y�D?5�K?z|�>�R�=��>�>�|,�Y�m�i�徂ʧ�N�<��?<Ɇ?���>r�N<�A�����]>���Ž�n?�Q1?�Y?���>�U��࿁U&�h�.�����}��d+=lwr��YU��������㽀�=�q�>���>J�>qHy> �9>��N>��>ݲ>��<@U�=E7����<󼔼稄=�ϑ� �<E\żR��	A(�^�+�Dt��
��;օ;��]<?i�;/=>���>WϠ;#�>K>�g�s��=�1���=1���>$.�WM��4E������0��5���j�>�>�H�D ���$?C��>FW*=o!�?�gM?�J�=X{]<�=о-���߽R�뽻)<��A�=Â��_V��~�̚C�����Y�>���>���>Y�|>TG?�0�N��M=�ܳ�Xx��?�n��� ��>{�tc�(w������oh�ę%�'KW?����؇�=7{?9�W?E�?��>�Z�?V�}�>-���(�<� ��9�|@ý��,?Ό#?}a�>�K�5�6�zH̾+���޷>�@I��O���^�0����#ͷ���>������оv$3��g��������B��Lr�Q��>�O?��?k:b��W��CUO����6(���q?�|g?�>�J?�@?|&��*z�kr���v�=�n?ĳ�?E=�?�>0��=�}��Ew�>P	?���?��?Us?GN?����>j�;�� >�ޗ����=b�>��=7��=�A?\d
?�
?�坽��	�,S�T%���^�]��<^s�=�>�>��>Axr>���=�hg=�@�=�\>쉞>�>�We>Ȣ�>%��>)҇�ޱ��?"ԍ=��>0�?-��=w5E>�L�b��=;Z������c%0���l�s�(��)�=�2�=T���m�>ڿÿfc�?Ṳ=>�B?�M ����>�=��~>}�t���>?���U�>S�>Y0�>��>�X>Ɍ(>Zcھ�>u�	�d]#��K5�ÝI��_˾v>�r����3��F��` �'l�B��}� �G�f��Ղ�h*E�B�?<�~�? ���d�o�ǻ#����<�?��>��B?����;Ľ�.�=Q��>j�>�澟���IL��}�ݾ؉?Bw�?��j>��>/�Y?���>�v
��%���bt��IY�-1.�=;T�~�S�qB��7.��k�
�\�C�P]H?�a�?F:?��b�J>V��?O��PY�ol�=sFK�1�=��ғ=Bў>����]�þb&���#��h������y?�b?~)?��]�:������>V�|?�I�>�11?���>4?��?!C?D�>-u�>{0�>]=H?m4?D�l?%�>�����ﶽ�^>LB�U���R�*<�RX�������ϼ>��<����L>��=ĵ��Jl�<k��=DR���̆�,�=s���L�=pK�>�$]?�+�>��>��7?��48�mB��R\/?�8=|��.'���b���U���>x�j?�t�?�VY?�b>>�A�U�A��>�f�>��#>/y[>�X�>����l_E���=[g>�r>Ƥ=��A�n����c	�p��]Ƚ<$# >���>��{>�+���(>����Dy�A�c>��R�g��(R���G�k�1���v��"�>�K?�?���=�d��֗�:>f���)?$0<?��L?��?�c�={ܾ��9��J����>� �<E!	����������:�$��9̊s>�I��똢�38M>�W�ðѾ��b�aL��߾��y=-���#/=(���־�� >�>,˾ʽ"�J���$��tTI?�̔="n������ƾ�E0>��>���>Z�x�������>�_(���.�=FJ�>��?>��~���D�t����$�>R�E?�r^?���?���R�p�wE@������(���%�)?7>�>�?V;C>r��=�H��B��D�f���F�`p�>���>�]�ȯG�%᜾a���%��8�>G�?Z>
�?]dU?΃?-�]?�(?�?���>ˋ�����>&?��?��=1ս��T���8��F�O��>9v)?�B�-ė>�?��?N�&?noQ?A�?�z>� �dC@�|��>'K�>ɼW�qK���`>�J?���>�Y?j˃?��=>'w5�GŢ�|T��7~�=	
>{�2?�1#?X�?y��>
��>���
�=@��>��b?U�?��o?/*�=�5?�3>U��>jX�=��>J��>�,?-?O?��s?��J?f��>�5�<i`���V��Ijr��5E����; �D<�yz=�}�(&s��1����<���;�N��zU��y]��\D��g���@�;�i�>�t>7畾��/>V(ž�v���@>A�����+:��j�=�X�>��?�<�>�#�O�=ٸ�>�.�>
��53(?N�?�5?�;�b�s	۾�K���>{B??��=��l��}����u��nh=��m?u^?M�W�x����[?$�^?�Ǿ��3�qH���_��:��jXN?���>~�J�u��>�L?��]?l��>��c��8u�����
�x�:t����=���>j"��@d�<�>hKJ?ԝ�>�N^>���<����w���ձ��$�
?#��?~N�?��?\A�=��n��ٿC��ג���U?MD�>�*��cX?ᢖ��e׾����x���5�ӭ����Os���I�����⪂���u��=�?�>{?��p?Ib?���$a���\�
\�ȵZ�Na �?��C�P�J�\zC��=n�����������U�;oEl�x�E����?�;?c��*�>k�������ž5e>�߬���
����=D:����&=f~=Ij>�]������?˄�>�-�>�K>?��[���?��:#��s9�����}>���>L��>�)�>K�=~�D���Y����u�n������>��d?iG?W�^?Sa6���+�}�x�!��,��z����rm>w��=Lm�>Y\��5��!(�:B>��!{�MY
�ǆ�2��V�:=O!?^q�>`��>�a�?{?{|��(¾X����6��=��>o�k?���>�Y>�D��< �$�>�I|?���>kl�0�\�1���UH���>���>կ9?�6�? �8>譣��)�l���܉�,��b�>�%?�	Q�ɗ:�؋�>�c^?vX�={�=�>��K�Z���ls��1ҽ���[�>�J�=H >!���[�2�����T��)?ܟ?Ý��4*�Dv~>ͮ"?���>DP�>�Ճ?3�>X�¾�x�;�u?�%^?�tI?zj@?{��>��=����q~Ƚ�&��A;=�ч>�w\>p=J��=�@� bX�'��5�6=�{�=�7ּ�����0<8᰼)7<��=[�3>x�ܿ�aN�U<־
B�j�ƀ����/�׽�N����3ȶ��F���w�H���V�L^T���k��3��Cv����?���?�����w����A�|�uz����>@/��do�񰠾=��n��>z����aZ$��S�i�k�`�h���&?Q�����ǿA�����ھxb?�G ?)zy?���j� �2�7��>FZ�<���ր꾲4��.�ο�V����`?
�>?2�Ѽ�v��>Y7�>�\>_�l>p0�������[�<�?��-?�T ?kq��-ɿ�k���t�<YP�?�1@n�@?��)�5�W_1=��>+�	?.�6>ew/�8&�J ����>�p�?��?��F=R�V�/6����e?��U<H�A�^�4�=���=-=8�#KC>6ʕ>�}"�0�9���ཊ�2>v��>V�?�r���b��`�<�
a>=Ͻ�U���Є?�;\���f�2�.�C���v>?T?ϗ�>�5�=}F,?�G�fϿ��\��x_?"�?0��?i�)?������>�1ݾ�M?+�6?T�>z�&�.�t�b�=,5���:���w[W�t�=5�>L(>z-����p,P�	&�����=���_�οg����A�4��� �y/	>t���6=��Vw��tþ5�R�P̪�3N)>�U>4n{>�Xm>\�=��L>F�[?1D�?��>��R>D�Z�9�\���n��:�����q�C��=���ܾ��"�#c������+�ê9�*��].=��j�=�kQ��ԏ���5Mc�ZF���.?�q>��ʾr�M��F&<ұ˾8���q�j�1ά�:�̾tj2�T�m����?/!B?�օ�~$X�|Y�R��r!��E�V?��-X�n ����=������
=oS�>�7�=a��u�2�z1R�Rg0?Q�?)���u���bw#>6��C=�l,?{� ?=�^<��>ʾ%?�Q+��余dT>B#0>�Y�>���>Q�	>�4��<�ٽHz?��T?F�u1���)�>ծ����x�8x=�@>� 6��rp[>���<F{���U^�y�����<��P?�>	w��Q��˾?���[��=��?��>��O>c1n?�J?��x���u��)��n�=�iO?�Va?��	>ǋ���?ž�夾s\?��Q?ȁ> ����ྥ��Y�����?�s?��)?E$��`O��2��H�e�-?6�?�GU�~����s��1�F���8?6�>׳�<Ջ��'�>�N?�1�c��l�ǿk?��8x�?�@���?q�=�R��%�5>�?��> �$�l��ZN(���	��v�=6��>��ؾ�h�~��4��'�r?=b�?���>�[�.]+����=�ݕ��Y�?*�?P~��tg<���zl�Yh��l��<���=��l"���e�7���ƾ��
����À�����>KZ@�E�S4�>�@8��6��PϿ���Tо�jq�i�?s�>��Ƚu���h�j�DLu�%�G�u�H������X�>^K>9���瑾��{��j;�-��x&�>��Z��>ERS��q��ڇ����6<;��>~�>O5�>��Pӽ�Y��?	/��]#οE����j���X?�r�? a�?�?o�&<��x��|�����;G?�s?��Y?#�(���]���:� �i?{|���.]�Ϥ:���I��#B>��1?��>�,�Gn�=�1&>�A�><Q>��,��HſP5�����+��?�z�?��{�>��?1�.?j���p��������%�܈v;B�E?�95>I�¾@� ��a:��n���?�-?vI���]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�k�> �?���=��>Æ�=�<���&^��Z>��=�jJ���?��N?d�>$M�=��8��c.��8F�+R��f�7C�쯇>�a?f�L?G�c>(���Z2�:� �|`ɽuc1�k`�ke?�؋*��X�4>Ծ<> ?>qB��Ҿ�S+?�%���G4����ƽߵ9?�s�=� ?g��ϻf��ߴ=�?A?���>�5���˰�ퟛ�F󞽙+�?b! @�v?�Aپ������>��>K��>Ěl�9�9�z8ﾷ����4?O`��P��㳁���:>���?��@W�?l��O�?�^��U���q��������=�N6?�[�� o>���>��=A�l�BO��#Fu�~߫>u԰?�V�?w,�>>h?��h�P�7�"�=�ӑ>?"q?Q�?uA��ݨ��L)>TD	?g
�x��('��l?��@��@�\]?�⥿E�� ��z���y���$�=�;>N��>4|��j��=&\�;f�:�<IB>�~�>�U�>\g�>{3>��>�݊>rԄ�Rj&��㭿�S��6�A��	!�Ⱦ�������C��e���c�[I���Ƣ<���vs=�� �����s=��>��Y?@KG?-XU?�w�>���<S�6>���Hڧ=$�E�<
�=�\�>�B=?�:?p(?Mŝ=����[�4v�ߏ�����7��>�H>�h�>�T�>)�>��;��K>�S>��>��=;:}=m�=槇=R3>+��>(��>@߾>mW<>��>J´�,��4�h�=�v��y˽���?+�����J��0���Y������欟=�`.?{H>����Bп �B'H?D픾�)�j�+��>��0?�[W?Jg>i���^U��>�z� ]j�ii>%���el��)��Q>�\?��m>¤�>��-�$�7�5�P����[Ǉ>Qb4?�"����G���t�WTI��ZҾ`�T>I��>�����#�Ꮩ�y}��e����=(U4?�H�>�����B��,݀��)����[>fiP>{W=��>��`>��vE��
7��F2=lv�=lP>�x?��->�`�=���>t֝�[�W� ��> jH>0�.>4@A?:.&?���� ��僾�M4�$�p>��>��>.C>_�H��=���>P�i>� �3I~�����(H�t6\>�{t���Z��~�x�j=����(�=�Ø=����l>��F"=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��>��:��頿�v��b�=��+d=﩯>�oO?�{�X�P>ҽdd�>�b?�;������D&ݿ	c���+�>� �?�?<�[�!䶿%S��?�>�`�?j�?���>��j���<ݬ�>�W<?-�v?�ڥ>2�0�9�i��X	?S�?#+�?(rK>e��?`pr?��>7�~�o�.��*���s���Ղ=�)�j�>�>�X���>F�C���F���gj��3�mZ>h�"=�%�>�s罦&��7��=Y���}���0��uE�>��m>�L>
'�>�y ?���>Bǖ>�=Iv�4�y� s����@?���?)�ؾ�Xr�.���R�=LbT�m�>x?����K��E��>�r\?�MT?*�C?GB�>s�*����� ���J��B�A=8�=���>d��>Z��uU����v ����L>�k�>�>�甾�پ�����h�>C2?8~?{۱<� ?��$?P�i>��>��G������uC� H�> �>4W?��?�d?͚���2����p���"Y��{O>�w?y0?=�>c���+��r-���[�w~�����?,f?6�ѽ��?F�?��>?D�@?�Wg>�����پ߽����~>�� ?)�����0��j%�� 6��?�,?s��>~�ƽ����_���%��L��?�X?8�?x=��t�!�ɾ��<֓o;|���!�Av�< �N>U�>�&�~L�=���="]�={����ؽ�H�<�A>��>{�=�K"�Sv���,?���;�Ӿ.)T>ēp����]��zx��Y�Ⱦ^5?`ľ�F��(���R�����7��?L7�?,x�?� W���q���Q?4/�?}{�>�s�>�q�Q�뾇����T�>�����':��=�Q�>���Ԑ=��g��}���r��r�R�q�I ?�{_>�L�>�
?�$�>1��>�)��������^�+W��͈�;]���/�&e��2���+6�
� ���t���gVX>��p���>� ?#SB>Up#>֎w>&�=�>��>���>=��>e��>ӽt>ZR>z���U�2�QKR?������'����Ⲱ�u2B?@rd?�/�>�i������}�?��?]r�?�9v>�}h�-+��l?�;�>���-p
?�a:=o���L�<�V����S(����Ӫ�>�E׽�:�rM�@if�8k
?�.?I-���̾==׽�����Nn=DJ�?��(?�)���Q��o�]�W��S����+Ch�ug���$�h�p�]叿u_���#��k�(�"*=��*?��? ������B��k�`?�xXf>���>��>ݾ>^WI>��	���1���]��O'�ﺃ��K�>!Z{?�>0�O?gL9?z�<?D?X �>�P�>��ؾ�v?��½a-�>@
?zJE?��"?�'?�x
?�?-�:>=� ��b�_�ξ0�?�?�?_��>i�?����Y��*׼Ќ���䚾d0�> ��=�%��Ӛ��:�q=�@>J?��7�3����X>q�3?H��>�n�>;<���9��74!=�t�>+�?#��>���q���
�1��>Z�?�P����=W�+>�F�=�(ļ��Ȼ�7�=�D��Ȯ�=�jQ�w�"�s�L<�M�=e��=�M�:�V��i���=;���<�^�>��>?��>����z�����#�T�(��ϟ= �0>b�7>9��<����G��Ug���E���{�>`ל?��?_%Ի��>$ >�a߾8/�@�>������>�K?�=�>%H?v��?��p?�KM?�:�=ç.�p��@���&�ԾZ�'?� ,?�đ>
��=˾����3�Q�?��?�%a��x���(�F5¾�Vսx�>$�/�o0~�Oﯿ0�C���~�i��K��W��?ŝ?BLB���6��辆����+��R�C?(�>�>���>��)��g��8�;>lC�>c�Q?���><�V?cQj?X�??^�@>�t'��i��Rp����<��o=�$E?�Ӌ?���?��T?'Z�>ٳ >�,>��0�����+�A����Q�=Sr>�"�>�� ?Z7�>	��=F���kF޽/eK��o�=��h>h�>��>���>�؎>@*^=�G?��>諭����[g���.���qC��Tu?�p�?��+?b'=eM�C�E������>�I�?��?�G*?cU�(��=�iҼϵ��qp��P�>m�>���>���=c�J=s�>ȿ�>A��>�v�����8��N�m?)�E?Nۻ=�潿By��8��9|�=�W�>'R��ց�Yտ=o�*&���IȾT��Z�����<y�k�����B��uy�7~羟�?�A�<�b
>�P�=Ɠ�>�d{��]�:2$@>�'����="j�|)A=0xb�kM@>�J�=ٴ���ʤ<v�=���_= mƾF�}?'�G?�M(?��A?�Yz>wS>�`l���>Mh��Ф?��h>� �_4���4;�f̥�u��d�پ�پ�vb�A%���D>��8�>H8>h&�=��:<^u�=��l=ӆ=s:��ؔ$=C�=ø�=ץ=�\�=�>"h>~;w?���Nɝ�7�P�����:?��>��=�nǾ��??,;?>s0��u}�����
e?D��?�l�?q#?��i���>WV������yE�=p!���1>j��=(�2���>)�I>���!T���W���	�?c@&�??�^Ͽ�7.>9�9>��
>)Q��a2���Y�5>_���^��?59���ξI�>�=Y�۾�|ȾS�=�{7>oGP=E}��M\�>��=�uz�c�2=�en=�ϋ>.�A>ٮ�=�s���f�=�M=�s�=�V>|܎98r2�T�'�3=�=#�e>�[%>A��>��?�b0?Nd?�7�>�n�j/Ͼ�D��QN�>z�=�,�>Θ�=�KB>3��>v�7?]�D?v�K?���>���=k�>c�>��,�1�m��x徃ѧ����<=��?ˆ?-ٸ>D�R<%�A�d���i>��;Ž�u?�O1?�f?|�>���k-�]l,��7�����a=Y��S�>wk���U���1:B�;���2>���>A�>
6�>Kex>C�>��>);>0f�=]<	;�|!=[����v��p&�s��=�<�<%����|н�k��'�<[�M�Cfɽ��S$�=����<�y��3�=���>��R=0S�>Zi�=����^Q=����P�(�K&�����{=_�d�g��{����4�Q�	��L:>�j�>��E�>���Г�>
0>��>=�i�?�oo?�p�>�r�M���I��	��r�r�!/�=A�="Ɠ�`
=��8u�tK��u��Ln�>���>�C�>Ĩj>�V-�6�@��p=�@޾�4�S��>�����!������p��R��W4h�v$���C?݇�
��=F}?rbJ?���?U��>�㚽V�۾�34>�F��!r=W��#�q�8�����?��'? ��>��뾕�D�oH̾J���޷>AI�.�O���V�0�<��+ͷ�G��>������оh$3��g�������B��Lr�c��>�O?��?]:b��W��/UO�����(���q?�|g?;�>�J?�@?=&��z�mr���v�=��n?���?G=�?k>ɬ�=�Ѳ�-��>�?���?ⓑ?��r?j+@�8��>Z�2;UC>�[���k�=�->� �='��=�?dj
?V
?����	�#M�6��]����<<�=E-�>��>/�s>j��=g�o=oV�=��]>��>�$�>SNe>���>�ɉ>� ��3H���6�>b�� �?��/?�
սh���`���Y���ov��w@�����Vb��w�HH->{T�=��6>�e�A'�>l̿��?<X�<x*�n�>%��Vt=�B�=�>F �Z!?�� >���>|�>�7L>_x�>��|>u�C=QDݾ�[�;[E���h���
���S�_�>B�>7��W爾Q����E��`���W�%�¾�����C|�[mV��b�=�A�?��=I���*N\�C��x+5?�ȸ>��"?�AZ�pkV=2�j>߶�>�?��������̍�-�@k�?��?穀>묓>xR?�
�>�p�{�~�+$}��4����0G���~�ſ����=$�GZ��#S?��?'S?�Y�w
<>�)�?ٍ���1�+��=��Z���0�5j�O�>�nþg\S��M���(���v��^=��U?yy?�d?z�K����=�4>�yj?k�-?w�?4?w�!?c���9|?�.�>(`I>"�?��[?�U?P~:?�ʈ>$;��eq��->�;�����F��<$G�=9�p��P����<2��=�7=���=Ud�;�(���!���=�=���<�w=� >�>͝�>��]?B��>�R�>��7?T�m8�&殾/?��4=w��������բ�-��c>�j?�ޫ?MZZ?Wc>_�A�3CC�;�>���>�#'>3\>@�>$�)F��͈=�c>B>J�=M~H�I���	�\+��y��<4L>`��>�B|>}׍��}'>����nz��d><�Q��ú�� T���G���1�V\v�2R�>��K?�?cA�=kq龃����=f��0)?�R<?KCM?��?Ԭ�=F ܾ>�9���J��L��2�>Q�<�������� ����:����:`�s>-��xؾ
�=q�澋A ���V�dh�G�J�#o>B�7���<���r�־���!�\>�?>�!��/��䡿�6��0�N?�I�={�̾�� �Ӿj.=>���>�$
?I����컽�7����ܡ�<��>}�>���޾#�Q��g���_�>L?��H?�݈?x�Ծ����VWJ������У�Ŷ��B�'?=7�>�?'5h>g�	�ѥɾ
���1q��wO�X�>e��>�m+�FdK�� %�qⒾ�%���>�m�>�&���+?L�L?�	?��E?d7?�9?�~>�!�u���;R)?�8�?U�k�����W��Ʉ%��Q��{?��>�|���!?9=??9F?|�"?ƨ?���>t��=���FV���>b7�>��_����d�>1sy?��>*�,?�Ub?-2>D*��A�P}>K�>�4>>*4-?��>t0?�1�>��>ӏ��ݥ�=���>y�b?�,�?W�o?�*�=/?k�1>���>��=U��>d��>�?�GO?ǥs?�J?w��>�<}��lL����r�5�M����;�hE<D6y=��6�t�>]���<��;gZ����{����8�D��-��}��;fX�>`x�>�	���M>�&;>D����2>�f��`��?.����@��=<�>�?n~�>���%pA=?m�>}��>���^�!?�?�T?>����_��pܾ�[�LȺ>�hF?	 �=T�q�����W�v�BU=�!h?^Y?�0W�!.��b?$A^?���0[<���ľ�Qc�@>���O?}�	?�J��ҵ>��~?�Rr?��>�g�ӻm����zb���m��Ͷ=r�>ge��e�;v�>_8?7m�>,�a>���=5�۾7�v�����R?���?п�?[��?G�&>e(m�SB߿9=m��,���.O??�1?�(3���	?�Ƙ�@a���a�d�̾�+��Xپ�� ��c������)^��n��ޗ���ZB�}��>%�L?uVV?��S?����		�һ��<�d�C�f����f!8��a�6���Z� �d���-����kڼ��y��:퀾��A�o�?�/'?�=+�p��>������pR;H@>,f�����g�=zˏ�A8=��[=f�^]/����1 ?�I�>w��>�;?@�Z�Ч>��0���6��M���.5>"��>V?�>T��>�,�;l^*��$�V4Ǿ�V��dֽ�P�>� f?�LC?P-t?e^n��D�����գ�E`��+y��2l>���=[-�>��+�4�f���-��24��Ey��������� �9E`=Q2?�K�>���>^��?��	?���=ؾ��W��1���Ϻ���>��h?ـ�>�>���n�6�i��>h�l?���>G�>5�ʾ@5+���l���;�*�>��> T?�ƌ>Pƽ�&<��ʒ�e%��+C@�u>�=CQ_?2|���d���v>!Fd?9Ļ�k:h��>%R���@ �-�Ӿ΋��-�=��>Ճ�=Q8c>�K�����O���T���="?�q?-)��LP+�Pbh>s ?���>���>]��?o>Ҵ���C=�3
?��Y?�G?_�8?�n�>1�=l�I�b�ٽ~$�'�=(ȅ>��_>�B2=J��=�N�*�>!�t�J<k� =j���;��;�e^���<�1C=:>>q"ۿ�K��2׾����2�Q�у�������("��ص�0/��.�z��y�z���wY��a�����ao����?�z�?)͕�K)�����W��VO��F!�>Uu�SLa�I�������N��s�پ	G��HK!���M���i�U d�[p?H!��,ȿ5�������B��>K�?q�{?�.����L��!�=f�N��	��ξ����[�ÿr��!��?�?��徲Q����>]]>%�>�2��Ma��W����>��?�OJ?_�&?�`z�d�Ϳr�����;���?��@*yA?�'�s|���F=��>٣	?�O=>�8.��)�"���*��>� �?!W�?�W=#QW��;�)d?;��;yG�$���z�=-�=׸	=�l�ϠN>6��>����a=�
oݽ��/>0�>�"�&��l6Z��|�<`X>�ν�6��a��?��b���j�7����p�Ǆ>��/?��n>��= �>?��A��sȿ0I�@�/?è�?�h�?dO?��Z���7>H��\s?�D?���>vZ�������iY6=�J_>�����v�~�Q<q�>,�>#H�����?��9(�8'>�� �ƿ{�$�np�:r=��ܺ?�[�������}&U��'��jo�Ҫ�Yrh=���=W~Q>�b�>�
W>_Z>rbW?�k?�Q�>�>x'佡v��H�;�$�_Q�����������[��߾��	���������ɾB+@��]9=�L��
��-��dmf��M<�C/?1�=J�ǾI0L�2�g<W�̾E��� #�忽TȾ�t5��^l�x�?�u=?���N�\�`��97�����N�^?8Q�bn��슞�:��=�=���Ȇ=�k�>l��=�ھ�5��:N��g-?��"?+���)w���@�=��	��'�<�t.?d ?x��:݆�>F�)?<���r��,>��>I�`>��>
->4��-Xݽ��?<W?������p�>܀Ѿ/�8�Z�>i�=�>��ւ�іI>L�R=o-m�4b�;����=R�O?fQ�>#5�p�H�j���M�꼵P�?{� ?o�U>?w?׆@?��=L���� ��P���Sܽ�rj?QF?-�+>p���"/���6?8w?G>0�U��V�X�,�œ���o?��o?a7?��a=)Q��F"���
�y�/?69�?�7��DЦ��r0�]N%>���>�&?f�]>.m�&?�MN?C�^��ML�|ɿ��_��Q�?�9@�'�?�e����
�=��>3��>8o9�(� ��cA�s�"��s�>K;?���D�i� 澻y��sHc?�ؗ?���>6���uI�O��=�ٕ��Z�?�?@����\g<���l��m�����<"ɫ=��2R"����s�7�t�ƾ;�
�g����������>QZ@�P�/,�>�C8��6��SϿF��D]о�Uq���?�>��Ƚ8�����j�(Pu���G���H�����$4>�H=���@�{�t{U��rD��P\=���>�z��R>3��YT���ű�+ф<"W|>���>��d>5V-���� �?.[�*�ƿ奔]��t�5?��?65�?�f�>�=>��Ƚ����^ץ=�`?�Ȅ?�E?sW=#��������j?�Ң��z_��y1��/I��'D>�U1?T�>{Z*����=>(>]�>�V>6�)��ÿ�ﵿ���V�?�>�?��9~�>�ޛ?tg.?�������2����-��J<��D?�*/>x��Z���`9�$����
?�1?�(�8��]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�4�>���?
F�<�*�>z��!��s�=a[v>iS>�ؼ�,$?�O?k?Am�>�u���+�H�L��T7����u-���_>�k?�+??�>��g����"�.�f��<K��N����s�何)�T�>8
>�J�>����M�,?��=�rٿ֬���D(�3�?�#">I4?Hc)���=e��=�&??�ǎ>Z�ɾ�h��˕�1,�=�D�?Ǣ�?/6%?�N��lgD>�>��>ŀ�>�Y	>����u���V�B=N�p?�+���o�(�m��~�>%b�?��@AB�?�rt��?OX��䈿:�w�$���T< �?�	>�:?�0 ����>�a?7j�=��n�%u��h�q�ʱ>0G�?��?�N�>Qk?�%p�7G:�� �=���>F~d??@/��t��6�A>�1?�q	�����\��	lm?R@":
@��_?����?ԿE����+���`�\�=Z:Q=В	;�뽿�>7�7�y��I����>eq�>�1e>4�j>i�$>��L>��=|i��P�"�5����y}�3���\|�{��v�_3�����������۾�����2R����k������4�+{�=�L]?�J?CO?E�>%I���w8>���%��=���݂n=e��>�,6?��P?��3?�W�=h����Z�nox����"���1�>?�g>���>���>���>g�R�={>��>�V<>�^>�u=�';4��d>5��>aY�>���>�q>���=�Q��p���n�c�50�����D��?~��y6I��U�������Ǿ�B�=��.?���=ҭ����ҿ��)�I?���������:�f>Z!8?�$R?�.>v��CC���l�=@)���s����=Pl�g�z��R*�6�>>\X!?�nf>��u>�3���7��P�t쯾�x>��5?���=/6���u�V
I�Yݾ jI>�>ҡ$��,�'����~�x�i��}=�:?	�?���d����u�GH��M�O>��Z>Z=a��=�I>yg��XĽ�fI��3=��=j>]>�?v�5>�=�f�>oW��,�G�cx�>ѧ8>��=>D?�?�;��d���y����2��>���>j�{>k>�`W����=�}�>�N>�A��G�Z���6�D� �?>�ӗ��T]��G����<���u�=�=��5E����<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>q�f��F�����?9O�E���Ԃ�>f�N?�
�mʈ=,f��?]e?��Ծ�Ԡ�7lп��p�s��>M��?5�?!a��D��r�&��_�>���?Ԃ*?d>�>O������+��>��6?A�\?�_�>��3��l;�=�(?���?`�w?X>I>)��?)rs?f��>�����/�����q��	}�=l�e;��>�V>tf���
F�kߓ�Mg���j����+�a>�%=��>���\����ٶ=�>��ɡ���Pd�^��>�yo>*�I>���>D� ?��>ؙ>s�=.:����&����RH?60�?����o�+Q9=��=s�J��d?8�'?#�^��xI�>��d?�ۀ?�T?~i�>�E�|�����!l��yR�<&|>T��>�I�>�0��Ie>�پ΄��^�q>gd>o�@��7ھjk_�3�;=�>�?���>���= ?<�&?8�g>$��>�zL�jn���MB���>���>|�?|b}?x?����1�ӯ���!��i�W�֍d>m�t?�?�{�>���	d��#U����(���b��>�?�p`?#|�C?��?��D?�F?�[>{�8��o�T���;.�>�!?��	��JA�Tw&����8�?߿?�\�>YL����ڽ5ļ ��÷���1?�[?�%?��Fk`�XH¾���<���y�6"��;'�X>?�>�&��g��=Ž>f-�=��n��a9�̝`<!��=��>b��=�#5�y����g/?�O.�)Ṿp� >�as��(�<�5=^l�=,�s���q?�jž4����Y��{��y{L�ց�?0��?h��?$���Sw��li?�CP?���>�C?����~��D3^����;:�׽����=��>f���,�3��哿
f������:F�=��I���>G�>�.?(�?ω2>��m>aâ�I��Fƾ����n�9�%��&M��-�&���ќ���<��kz�����1����B�>bKa����>�P
?�@�>��{>�0�>J�b=�|�>���>��P>��>~M�>��>.�M>sK���ѽ��Q?������'�i���N����A?��a?~!�>��p��4�����n�? �?^C�?��q>6�f��)-�Q�?e��>�����	?��\=k2���<󙳾�A	�[����ļ�؎>�U�*<8�XeL�b\��?��?齼�0ʾ�%��Ȇ���Ѽ6��?�#E?$��G� �Z�f�U��L[�[�r��������P���{�mѓ�$���r�~�81�||4�]�)?fUw?������Wa��X_t�S�ە�>5��>��>���>���>�Ͼ���fG��V��b�J��>A�?���>�!J?�;?��B?��C?{q�>���>����9?K!�����>�h�>�2?��*?'�/?�y?�\?q�[>�?�������־�?�?z�?{��>ɞ�>$߇��	��O��+Ӽ���I��<=8=��<t ��bT��Sw=uU>J�?՘Q=í0�0=
����>PB?'�>�8�>������j�=-��>��(? &�>�xɾR�_�
�&��> Bc?�#��\#�=�W�>h��=���;�S�<�5>�,���/>O� �0������f'8�,�=`%�=s��:�E6��"
=[
z=E��>�?>?)�>�!�=����<���/� �=���>�M>�3P=��	��[��Rܕ��Á��L�>�Ѝ?6ν?��'���=��c>�Ͼ<a�quJ�ù� t�>�QJ? %?[0?e�?�>k?!UN?Xx^>��*��_��S���H����%$?1 ,?�$�>
��
�ɾ�+��U�3�g?��?~x`�� ��(�d����#ѽ��>�/�E~�,��
�C��麢���5��U>�?�?�BI��F7�i����������D?8��>�+�>���>g()��(g�1���f=>v�>j�Q?��>�O?{?k[?�hS>e~8�L������0#�l_!>@?)��?p֎?��x?07�>�z>��)��	�����o��"����-aW=a�Y>�z�>n��>���>T��=C�ƽn����?�dM�={.b>�t�>���>���>@Rw>R��<�G?ۻ�>������أ��Ё��eK�+�t?�_�?��+?��=��3�E�<����>�a�?f֫?p�)?�FU�`��=��׼���Hnp��ڷ>-׸>�>�}�=@�>=��>�>���>}��/t��8���M��%?@ F?϶=8�ҿ�Tl�u1��l��<��1>��U��3l�2�u�A��`SE�Oq�Ԑоt"�)'Ǿ�
߾��þ' о�þ�Sվ�� ?��=���=�:=��=���`�����=�iG�@�a��U~��J��#i���u�k_A�1<V�=ܯ�<0ޢ=����`z?.FJ?�0?R�7?�y>;�>𨜽��>M뽌?#�L>-ڭ�_E��O��Q���诙����o����c����s�?>K�=<�:R>�� >���=#��<>��=xR�o�:'�8<��Q=�g�=1S�=��=W��=ޠ>l��=�x?RX��T ��0�M���ѽt<?��>�E�=U�ȾVeB?�@>=����Ƿ�e"��:�?��?M��?�a	?.�r��ǜ>��)�x�yԊ=>����2>�f�=-�3��Y�>�oF>����J��I������?
}@�J??����Aοqw.> �:>�>�S�|�0���T���X��jd�µ?g�8��>Ⱦ���>
��=־mLƾ�F=��8>K�C=���#[��p�=��Y���l=Y8=���>�P>B��=ۻ�i��=�"3=��=Q�K>���wV"�M��.=槺=��c>9�)>�J�>�?0L0?�c?$��>Om��ϾDE����>��=Md�>�+�=�lB>5��>��7?�~D?pK?8<�>�=���>߶�>�?,��bm��8�˧��<�S�?�Ȇ?�g�>qR<2�C���9�>�h�Ž	Q?�1?�Y?1D�>�U����9Y&���.�$����{4��+=�mr��QU�M���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=$�����<�vż�����u&�:�+�1�����;r��;B�]<^��;��>O��>U����>�x�=ở�B��=9����*�1͇>��Ͼ
�M��"F��+��*�(��<s�-9>/�Q>��D�?Ҏ�{Z?��;>�G>�b�?�Lg?0��=^۽7:Ծ]����%?��d�8XD=p�J=�i��cG��Op��K�6^Ⱦt��>���>���>O�m>��,��?�l�v=Q-�j�4���>������3f��[p�hD���響��h�	�P�όD?�����=D~?H�I?Θ�?��>:u��՜ؾܫ.>����5�=<�csq�#����?ʮ&?��>���D���۾#��=��>J.���C��5���)�ϔ���þ�L�>o���{�վX�6�A��� ���!TB��)z�G�>��I?�׭?�%q����I+W���*l���%?��h?��>Σ?��	?⼁�Ѿ�H�Rj>��i?��?���?W>���=�%���s�>�	?��?���?lhs?��?�x��>bmu;[� >x�����=},>胝=Kt�=�@?kh
?_�
?y����	���:���K^�{�<|H�=�F�>�w�>E�r>�T�=S�g=�M�=�D\>F̞>�><�d>��>b�>#E���hY�>!���"�>]�F?�=��"=�C��wn>e�ؽ������~k����v�o�@>��>A$=o%��/��>�9Ϳw�?��<�C�?ŇϾ�j�<�r>H�=��>��"�>/I>���>�>ʹ>	��>I��>�%C<��侞?=�v��P8�.#�I�F�|�����>{��$T���(�}ہ��¥�d놾V��I[u�z�u��Se�	>��?�q��^z��v&��~=f�?/>1
?;�U���<�A�<A��>���>�A���������2�����?�
�?�F�>6,�>H?*�>��w����%���2ts�C��i9(��Za�}=��/���$�E��o?{�?+�P?$U���e>�ӡ?�!վi߼��= v��0<�>+���[>^+������3��q��B������4?W}]?*�A?�M0�y�W��Ow>Fm?h`�>�Z?�Z+?�h:?�9���a?pӗ�`W�>�j;?�%?��A?L�1?A+[><e�����YR9>��J�����ߐ<x~=�ɉ�D|n=@.�=?�Y��+=�+�=P)=�3���;0��=���<�N<�L=��k<�ߝ=z��>��Z?��>�-�>�5?*���<=�ٮ��-?3n�=�n���\��rn��{���)�=��j?Q
�?��R?XmV>ƹH�vT6���<>��i>*~>�n>oZ�>Ե��ޠX�Fi^=d�>��>��=Xr~��n�����R��Au<B)>w��>Q�{>_W��&(>Dd���*w�m'Y>P�Q�֧��W7D�;�H���2��?t����>8rI?�?u�=��澨����e�0T)?q';?��J?H�?`��=�m۾�R8�0)J�mn�T�>��<h��8���a��GV;����'m>����ᵠ�R2g>S��ǰѾ�k��I�_k��A=�H�{/�<����E׾�����=��>�徾��!�Z���������H?NP�=���wXm��\þ� >�4�>w�>1TC�5v��N@�����؍=)��>�Z>��x�v��PfI��%��{�>�H?D.X?A]�?�����m��@6�
q��s�X�/�Y�?�W`>Hp�>l�->*k>l͢�+O��x�tYO����>Jn�>�R��]d�wQо;������G}>��>��=�O�>Ζ;?��
?��m?�`N?Ac
?g2�>%U;�Xlݾ)*?���?�d�=Ȗ/�}泾�d"��%<��o�>#�+?����˗�>��?��?�0?��f?��?![=�+�5�[��׋>^��>��M�Z%����>׵m?�K>$-E?:�}?1�=>}�����"}�=7S>k�N>��/?:*?_?��>�j�> ���J-�=�!�>�)c?��?ɗo?A�=��?I:2>�
�>�v�=~-�>ـ�>�?�6O?��s?3�J?�S�>[�<�
���˵�b�r���N�N�;��K<1t=���Vu�������<���;�庼� �j|��LB��"�����;.8�>33s>����EU0>�yľ�E���+@>/<���0������s;�A��=��>��?鬕>`A#��_�=�̼>��>��%U(?��?b4?V��:�b�ϙھ�PL����>Q�A?"��=%�l��t����u���e=��m?�v^?.W��X���b?l�]?Q��>�<��PľjFc��d龋�O?��
?XlI�߳>hj~?*�q?���>��d�5�m�����b�Jl����=Z�>BA�xAe�Sc�>ٯ7?�M�>l�b>\��=�S۾��w�o��!-?��?��?Q��?G*>�n����򾤟��)0]?���> x���8?"�ؼ���&��u�3���X��u���?���}��g�Vb��닽?3�=��?�z?�l?��]?����c�&X�CZ~�JW�������C��E��lI�sUo�`x��&�ZU��C��<J�{�lzB�oG�?"?�!�RU�>�F�����Y&˾s�>>e���i�&�v=Yu���d=-bk=�^V�������I�?�E�>X:�>T'<?��[���=�p/��i8�� ��&>���>^e�>���>�n����8�Uh̽���Ō|��&�Pw>`?Y�A?參?q�z:�P��C���_<NŸ�O��>���=�kE>��t�����<O=���u��D��Z�m���>��?!$>&�>�p�?T_�>� ��$����� _A���)��_�>`�p?)��>�X>j#H�[�-�-l�>_�i?K��>`�i>Φݾ�+(��gz�%�=O��>r��>�?�>��>�IY�o*�厃�#ɋ���H��U=׽q?6�e����=)�>֭w?�>�XV"����>�½Cl(��	;tH=�Nu>��><K0=00�>��L���u��G\��?3?�ͽ3),��Z>� /?h�>���>[~�?i�=4�Ծ�>�8&?��S?U�d?"�>?�t�>۝��Of��q⽡/�$o>?��>,�Z>"��;Σ!>^@�p�>�����6���B=\Ѷ��ڽl��<ݬ��ln<�P=N�N>��ܿ�K�7&׾�{�Yu�@H
�	����,�����������n���u_��Q\��"���T��2i�-x��-!r����?~1�?����֋�d����S|��B�����>� u�)���/����B1��g"ݾ�ݨ�<�"�L�O��\g���_�u�?X���Mǿ����V�;��?�t?!�x?EK�~}���8��>�=�?���^�ݛ�>OϿ
����sd?���>
��\����>!'�>l�f>��m>7�������l�|=g�?|:.?��?�vZ�� ʿQ��VC�<���?>�@!�K?�MN�����=��
? ?|I�>]#���H��|��5�,?ɦ|?���?��=|ge��λ/u�?t�> ��߸?=Vax=�2">�/+>�# ���8>���>���������S�<�t=���>H�K��;���I�o
�>q�>c��ku��5Մ?,{\��f���/��T��U>��T?�*�>R:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�݅�=x6�ԉ��{���&V�}��=[��>b�>��,������O��I��U��=�����ƿ�,$�g��]*=���G_�,�� ����U�j���#�m�ܻ�'�i=���=�fQ>�7�>I@V>�X>|W?S�k?\�>�>T��5����D;��#�z����ꇋ�<Y�����F��޾�:	�Er���yɾ��=�ф�=��Q�~����< ���b�aVF��c.?A�">�ʾ�xM���&<˾�y��R��pʥ�G~̾��1��n�6��?�B?�1����V�+��#+ ����~�W?������묾��=�����+=pO�>W`�=��2�2�R�R�/?� ?͊��6�����=�8�>y�;��5? ?�0=+�>	�*?�w>�����8B>�� >mĆ>É�>Y;6>v}��8x ��?��_?���(����>�T���U��ܲ�=��R>�e�NE���B=>3�Q=����c;��Ľ�d�;�tF?w#�>u����@��|߾�b���q ��2�?:T?���>�,U?Km1?yL��!5ҾHK[�h������)C?ǂT?�6>+x���S������)?a?~�=��4��3��F�Q��>�j?�]7?>?��.x��.����[��P?�H~?�~��˗��	���=Z��3�>��S??�G>j�d�>U�D?��2�?0}�G>��8�@�O�?s]@��?���=�HS��*F>�?���>���i��<����o	�C�>>��?�I�*XB��|;���& 4?YB�?�y�>>��r�e��=Tە��Y�?��?�{��+1g<l��Ll�n��lc�<���=#���~"�|��T�7���ƾ�
��������*��>^Z@uS载+�>�S8��5�4RϿr��7]о]Tq���?x�>&�Ƚ0�����j��Ju���G���H������V�>>�H��`ʑ���{��q;�Y�����>m|�rÈ>��S�A;������d5<���>���>���>������l��?TJ���1ο���î�u�X?�b�?�d�?�i?si7<��v�Ӏ{�m���;G?šs?�Z? B%���]�l9���j?����`�84���C�_�W>��3?�e�>�&.�Qrt=�%>�!�>^�>c�-��Ŀ쩶�op����?x��?��[��>�X�?[�+?F��.ۙ�l�����)���˻�h@?R6>�Y��j!��=��:�?	X1?�	���]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?���>3�s?��=%o??4]��	�eT����>�N=>�h�=yC5?�j?�\�>�GL=��6���)�D�&eL�뿾�5(�>�T>��L?�]X?�%�>�}��,��{�~��.���}iF<<����u=��$�։>ZM�>Z->��o��#�e`?VY���ܿ����֏�=�uM?�>#��>���.�轥�>�б>*f�>��9����3����t���?�/�?R�?>=ʾ��>Y�E>v��>�94>��!>�P=�ľI���j?�f�-�t�yiY��۳=j5�?�@�v?�[~��	?.(��Q��Y~��x���6�&.�=\�7?B���z>���>�٪=ncv�����Y�s����>�C�?gx�?���>2�l?�{o�^�B��p2=AJ�>t�k?�z?�Us�s�_�B>��?������Q�'f?��
@�r@)�^?$颿��ѿ����%���[�$�>���=�<>�$н���ΰ�<�q�I >v�e<�P�>JS5>�W�>�g�=���<B�;-=z�����h���`������S(��g�����DE�!�����̾���"���
�������q���
���;��J�=�&R?��p?�1?���>�k�=�M>�8��қ�>�룾�|�y�>��B?��6?&�[?�U>����O�\�Pq}�S����ċ�,.�>�v>~L�>8hs>�~�>Cc&�S:�=��i>�>L�=�F�<s���6[<v5;>���>p�>m��>XC<>��>Aϴ��1��c�h��
w�m̽,�?����S�J��1���9��ݦ���h�=Gb.?|>���?пd����2H?����)��+���>��0?�cW?:�>��s�T�":>?����j�E`>�+ ��l���)��%Q>l?�f>�Nu>�p3�b8���P��Q��EW|>:/6?ɛ���9���u�"�H��<ݾg]M>"��>TC@��a�~���]�Kxi��D{=�w:?��?�z�� ���u��?��9WR>�\>�=oR�=\mM>
�c���ƽ,�G�'�.=���=��^>E ?�B->���=�_�>�����T�"��>^B>S->Y�??�
&?�C������|h��#.��@t>	�>-�}>�u>q�I�7�=T��>��b>x�����o��q�?��V>������_�k�����{=�ߚ�9#�=Z��=Ae��_e>�ƚ=�~?���)䈿��e���lD?S+?Z �=�F<��"�C ���H��G�?r�@m�?��	��V�B�?�@�?��B��=}�>׫>�ξ�L��?��Ž5Ǣ�˔	�%)#�gS�?��?��/�Zʋ�;l��6>�^%?�Ӿ��b>�����%���+~�g-�@��=�0�>�]=?�����=�BH��l�> � ?��x������ϿA���j��>���?��?A�r������9���>���?��B?���=%SR�o�8=�"�>��*?�b?�t�>��*�Т��1?���?2J�?��H>TX�?Hs?�I�>8�w��/�~����"����=
�;��>�>�^���F��t�������j����`>
�%=p�>y߽���|N�=�;���V��u�a�K��>6k>wF>\��>K} ?�]�>���>]�=4��t����ї�@�E?/��?{,ҾJ�v�"q����o>v)��b�>	�F?�ow��u����>j�p?��z?�Um?D�>���������὿�	�����<!b�>�w�>[M?�w=zT>�����=ƽ��R>E�8>�O=󃐾�Or�4���:0t>�?D�>�>�r ?��#?kj>훰>��E��i����E��>22�>ۮ?��~?w�?F���03� �������H[��bN>ؑx?D?���>����\���mA�}�A�r����T�?	g?�V���?U�?֑??��A?4�d>���.-پ����轁>��!?�C�A��L&�����?�M?_��>���#ֽ�VּA��gn����?�)\?m?&?#���'a�7þK-�<#���O��q�;�D���>z�>}������=�>��=kBm�nC6��e<�z�=���>��=*7��s����)?q��������Oh>�����b�����>�ͅ��G߾�t?��O�tOD�������� Nx��Ҋ?��?�G�?bh���e�#7v?�;a?^?]L�>�}þ�S>�<���k��=�IQ�.c��m����>Z˾��cR��F��+�[�"��R�I��j�>XE�>�"?/� ?Z'=>@�y>�j��s �]�Ⱦ���j��Ԛ�]�F��1�����+���{���P =uû�헾q)�>��P�N��>(Z�>� �=��>��>kO�F=?>��>� �>GG ?L'�>�T>�=b	�N��7�KR?,�����'�%�辵���!4B?�ud?9�>�i�����8���r?$��?�q�?`v>	h��+��r?5?�>a���k
?�:=M<��Q�<EU������%��4��/��>�׽H:�-M�ҋf�h
?9?����U�̾N׽������n=�M�?��(?��)���Q�g�o�̸W�"S�9��D6h�Vj��n�$�֛p��쏿�^��%����(�p*=��*?e�?��,�!���&k��?�ef>	�>$�>�߾>�sI>��	�B�1�%^�M'�p���R�>�[{?��>��I?Z�B?��A?|�D?n�>�A�>���R?mJ�]f�>�=�>N�>?7c,?2;?�?��"?�#3>�M"������־i?�M?Oc?..�>7q?7����սѢ�y���j[}��&���5=��<��Wr�+�q=�jQ>�i?k����8����c$k>�p7?]��>�b�>����-��2�<#P�>�
?�w�>U? ��kr�0����>���?t��J�=�I*>��=���HiӺup�=3�¼~h�=��}��8�� 5<D#�=͈�=B|B�Z	�:Ѥ1;0�N;�O�<���>?�2?�g�>���=cþ�TA���-���~>Wu�>���>�>:���o��ݪ���/T�.Y�>?)�?3r�?	�\�_�>Liw>��վ3��W&��'��A=+D?o�P?ke?.ƛ?+%F?�?`>�:2�����恿�Oɾ�
?�,?ʳ�>���,�ʾ����̖3�ns?i�?�a�!"�	)������ս�>M/�n3~�� ���D���Y�������_��?�Н?�@B��6���羮����w��F�C?ǽ�>���>3��>Ծ)�\�g�}
��e;>S4�>�Q?Zл>�O?q�z??�\?��S>H�8������p��\��z">|@?��?ו�?�=x?Ӻ�>%>��*���������F�𽈗��kT=3$\>�֒>��>c	�>9"�=h�ϽH��Y^B��å=�a>��>߾�>7��>du>칛<$�G?3��>�]������餾�ă��=�W�u?�?!�+?K\=����E�+F���H�>�n�?���?E4*?3�S�|��=��ּ�඾<�q�s$�>�ٹ>�2�>=oqF=�c>�>J��>�)�.a��p8�+@M�~�?�F?I��=%Nɿ��v�Vv)�Yά�V�>A���8�r�f!�ڂ~���=[����tս�Wξ�p1��݂��9��7z��v��j����f�>���=|v�<F=Zߍ;>a=K==0y�G]l�`V39��ŅD�����ዼjǤ�Jj���)�<m�=�⼺�˾�Z}?�I?�D,?�lC?{%w>Hl>��3����>�n���o?W>
O�_~���;��R��vf���"پ�9׾�Uc����OY	>��J��?>��3>0��=3�<xK�=/f=�Ҋ=`���%=�+�=��=�z�=�$�=��>�\>�6w?X�������4Q��Z罥�:?�8�>Z{�=��ƾq@?~�>>�2������zb��-?���?�T�?>�?>ti��d�>J���㎽�q�=S����=2>`��=z�2�V��>��J>���K��H����4�?��@��??�ዿϢϿ5a/>J�7>��>��R�j�1��5\��Mb�� Z�ś!?�M;��B̾jb�>蒺=
߾&gƾ��-=�T6>�7d=���<\��)�=� {�E�<=_m=։>;�C>��=i���6�=��I=���=�	P>7���9�¡+�{�5=�~�= �b>i�%>�}�>6�?pb0?C>d?�%�>�0n��6Ͼ;��_E�>���=��>�2�= �A>Z�>��7?z�D?u�K?!��>�`�=���>�>�>x�,�ԟm��往	����<P��?M҆?��>��V<ðA�ܘ��a>�[�Žvm?�B1?�Y?M؞>�Q����8N&�W�.�/��v�ҷԴ*=��r��AU��u��A�������=�r�>���>��>�ey>� :>��N>: �>ܧ>^�<di�=pЌ��<?����<�=Y�� ��<�Ƽ�\/�
,�D�����;a�;b�_<��;@K�=)+�>�W=v;?x[t��Ō��>�˾d-=�Ȏ�>�?��l�`�,.V��!���`3���N��'C>䅆>:�f�E�����>ҪP>��L>���?C?�+�=�;�#���h���>��KE���t|>b$e>2f��M�A���x� uO�1�����>� �>�͢>��m>`d,�Y?��Uv=8ᾓ5��g�>1o���������p����^럿Mi�J���D?u&����=3�}?�(J?�Ϗ?B��>E~���>پi0>|��=۸�O�p�"����?m '?ʑ�>����D��H̾b���޷>k@I���O���]�0�1��ͷ����>	����о0$3��g������ƍB��Lr�f��>#�O?~�?2;b��W��tUO�~���(���q?�|g?"�>�J?�@?�#��az��q��ly�=�n?���?5=�?<>9�=�����>��?���?#��?Cs?ŧ?�g(�>k��;H�>G����V�=a�>�̜=Q��=Sb?ט
?�
?𝜽#�	���ﾨ�r]����<!ҡ=	
�>3�>e�q>���=�k=���=Y\>�'�>�+�>ye>��>��>'絾��	�6g?��v=S��>�(?�@�=a��=�猽��<V:�0���S�罏q��|9��=@=���<��>�1�=���>��ÿ#�?b;f�*ा�F�>��Ǿj���\(>VDr>�v(�;?����"��>?g�>V��>K �>T-=Np9��%�<����/��;���{8��1��pj�>�l�~\r�<����p�:ͪ���u�*ܾ��c�?����N��ִ=T��?v^��)��
L��Tͽ��?���>��M?d��>�O=�̋<���>��>�����������-��<�?T*@4=>פ�>�S?r�>v��/�\��W��쀿�	8��N���m�����!������;́��T^?�y?�M?t1S���e>�?����9��y�<�P���;��j3> �>�Ez�s����
�6%Ծ۝�i�U�/_h?$Wj?B ?d\J��IǼG݆>�`?�'?��Q?�26?�_?����>8?��x�l(>(?"1A?.c?��=?[�>��=�6���~����酾e��"fǻ�=�m =�W]= �����2�\A=��e��L��� �ؽz�{;`Gb=Z�>�Վ�=dҮ=؟�>.�]?���>�y�>:�7?	8�[K8�����>>/?e�6=qA��7ъ��Q�����->X�j?i۫?�Z?%oc>7�A�IC�� >Ah�>�y&>$�[>�&�>�c�_�E���=a2>�{>�ݥ=��N�����u�	�k���n;�<�>l��>|>�Ս�
�'>�e���#z��d>R��ƺ���S�k�G���1�'�v��T�>��K?�?ʙ=�K��@��%Af��6)?�Z<?6MM?&�?�ܓ=�۾��9�6�J�zJ�0�>��<y��V����"����:�~p�:L�s>�9�������72>���q%�dX��8��8�i6������=��
�������I�=��=���#�(�_����Ȧ���F?���=W-��:{G�ق��t>��>��>��8�|½�D�q譾�8�=��>9�<>�����|�8��Ǿwl�>W�E?O�^?v��?�R��w�r��mC��a���R���|��K?Z��>��?�fC>7�=K@���j�ӧd���F��}�>�j�>9���9I�����E
龾#��,�>��?y�>?GtQ?�e?��`?�**?r4?��>�ý�Z���$?Pd�?��&=�=�z����Q�B�m��>F6 ?!��>�>]N?��(?Y�.?�[O?ޅ?N�=iQ�=Q��i�>^̉>��\�oݰ��eb>$[Z?���>��D?]h? �o>s��k�%W�=L�>��3>ޗ2?�?@<?@�>��>�q��?�=�`�>|�b?� �?l�o?p%�=D?Z�1>/��>ބ�=�ܟ>`��>�6?NO?�s??�J?��>0��<�r�������s�m%U�BO{;��I<!{=�����r�������<��;Mֵ�N���8Z���C��������;z�>x�r>ˀ���:4>Qrž�h����A>�G���F��L���!�9�p��=�~�>�� ?���>������=�W�>�%�>����(?��?�?�?=;²b�u|ܾX9J����>�JA?�C�=�ul�􂔿�5u�/�l=�l?_�]?�V�5s����U?�%e?OOȾ�%���Ծ�P�7���`B?-�?��о���>z�O?�8^?D� ?�_4�4�V�MT���<c������>o��>L�<�.Q|�Z��>�u?N4�>/f>���L^�;W�"�R��l"?'Ό?J�?:��?j�V>X6q��⿧0��������]?�X�>���6�!?P]���ξ�ދ�IZ�����#�|�����͠�!'���t�t8н�؞=�?*�r?��o?5�\?J�����`�cSZ�=瀿��V����R"��@H�F6D�0�@��0n�������㕾��+=�A��U;A���?�q&?��/�x�>}����e��;�A>')������ь=X��>fC=�S=f�y-0�&`����?��>�M�>��;?�Z��=�b�1�u38��[��˜3>W��>+ɑ>j��>��o;-0��=佦�Ǿ�'���ӽr�k>]Uj?\�R?�ju?F�9���S�xކ���y>8ª��>��=Au>� �͙�ܗ%��C��)c�:�Ծ��^���(췼�?��>R�?=�?q
?�V����p�	%J�=�=>̾>�!J?�� ?v�>�o��jX�3��>I�t?��>��P>\��E�O���_���3>���>��?WR?ՎK>��)���/���pH��3�C��&6>�m�?�n�26f�f��>�Vx?�RC=�(%;�Ɩ>mR������k������1�>���>3ҭ<;��>e�>�
���)ϥ�!�"?*�!?�2r� =8�{l>�(%?��?K�>�5?�G>'T[���,>�S5?�g?��H?|<?��>�ڼ�����~��2��U�=R�>i�>c;�
y>�׽�������\���D>d��ʼ��#=,T��q�
���=��>ilۿ��L��ɾΛ��p�a����Vj�J!�#E��!$�*Ҿ����m����D���4� �V��@���o��#|����?��?o��=ܞ�k���x�y�����e�>�����:��pN���8�]��������
�������M��c���p���?kڠ�t�ÿ��ċ��),?�S?e�{?ߤ2�&o��X�Ӄ6< ����>~pо�Z����ƿ�#ž)�k?1	?� �zѾ躐>�W�=�^�=}
E=�%e��<��o>|�?%Rk?0�2?��ǽ��ÿ�v���d�=��?S@ȜM?�7���
�š>[��>� ?�ޝ>�	��G:*�s�W�V��>8�?Z�?Ƴ�H�S�G�	>L	p?�'�=/C����eb>Q�>�8�=��p��k>VL�>Oh��ݏ<���">�>.&=�����!�Qa�<o�x>�u߽����5Մ?*{\��f���/��T��$U>��T?�*�>W:�=��,?U7H�[}Ͽ�\��*a?�0�?���?-�(?$ۿ��ؚ>��ܾ��M?\D6?���>�d&��t����=�5�"���x���&V�m��=E��>_�>��,������O��I��T��=�4���¿ɦ����=,�v= g���7�D�ܽC��+̾8���q��4W�=X��=@�6> �F>�>��D>�W?�5q?�ܹ>C L=<�� /��G����3����� �jH���-��ɾ�Xg��.����|E��K辿>=�<��=8�Q��k��B��yb�]F��.?��!>��ʾr�M�#��;^�˾���0���e���B�;cu2�A�m�脟?H`A?���o'V�Ap�'�F]��#�X?����K��@����=�P��DO=E��>$�=;��I,2�ԴQ�{a?մ?DNɾ�
R��'�>6Խ�[�`M"?Gi�>Ia�����>��/?!N,�����N(>�J>��>���>�˼�����!�N�9?�1?|��m޾Psy>�WO�Ԝ<�2�`�ľ�=3�9�t>Ͻ�e�>�h>���͆,��(��&�=�Q?��>P���^0�Уݾ��-���7�<�?�~?�{�>"�r?�/?�y��dӾ	`c� ����<�gZ?��b?��>��T�_%Ҿ9�i��{?(1V?^�>VMO� �����z)����
?76i?��?���<�����n��[��'�@?�
�?��������;2<�\�˼�c�>�B ?�7�<��o�hя>��2?�
�=�6��$���|2�d��?���?p�?���Gۓ��P%>}�>�\?���� �!=�1���"'>��?�׾y n�}R��{�оɺ?�#�?���>iU������=dٕ��Z�?)�?����Y;g<����l�Sn��Nv�<�̫=���Y"����|�7�/�ƾ[�
��������c��>2Z@�T��*�>{D8� 6⿼SϿ�� \оMTq��?�}�>�ȽD����j�;Ou���G�h�H�ݤ�����>w>Jt���M��}�z��:��Ѽ�\�>�G� ��>�nO��Ӹ��m����b</$�>��>��>&
��PB��Z=�?OX����ο�Ҟ�ݓ��X\?��?�6�?�k?�H����v�\nz�ET���pG?�+s?2Z?�0�C�a�9�g���j?/b��rV`���4��DE�'U>�!3?C�>�-���|={">��>e>�"/��Ŀ�ض�S���?��?���?Fm����>���?�u+?i�i7�� [����*���-�8;A?�2>6����!�2=�fВ�J�
?O~0?�x�</�]�_?*�a�M�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>hH_���u>����:�	i	>���?�~�?Pj?���� ����U>
�}?�>ō�?O�6>t4?7z�����+n�	�>�]�>�>�?��I?��>�=N趽{*D��K��pD�8�W��1@��Qu>�j?�M?���>�����-���<�A��/��� g�=^��xa��D���>���>r��=o�y���ݾb�6?B�6�Hyݿ[��.)#>��-?�h>0�-?��&��c��>1��?���>9"��O����:���>a��?�~�?@�?�^	�Wǽ=q��>\��>�eH>�󽹉��*��d�e1U?q&�<L���E���I>���?�@���?ǜ^�iK	?y]�Vd��{~����M6���=�7?��U�y>�&�>X�=T7v������s��r�>�T�?l�?��>��l?Ďo�P�B�J�:=�ѣ>�>k?�@?�ٷ���dB>��?���p玿ø���e?�
@�Y@j�^?X�A=տ���[�P�~,����=A�>>�>��c�,k=ț���ro�wR���=pO�>(;>�*0>4��=��=��=V����b#��虿gy��R�2��y��A�����7�E�� �e���5�پ���cv�	�)�a��f���������=�=W?8�R?A�d?u?��e�<l">|����=����)�=�i�>��2?�FK?��@? ��=�:��؇]�1�}��T�������>Ǿ0>KB�>>	�>]�>�LǼ�i>�.K>[�e>���=Б�~q/��͍=�R>���>���>���>Y�=kL�=�x��p����1�'�O=r=ym�?�;۾�S�}������>�Ak>F�?~�B=���uϿ�͘��K?�ؑ��`3��D��B>{�H?u�?}w�>c����V��\�;��B�)wV�*�\>�`��Jn��2���~>�w,?��d>t7t>7H3��e8�[�P�Iﯾ��|>�5?n����j9���u�I�H�L޾��L>恾>��J��r�]���>�ZNh���}=:;:?i,?ؘ��e�kw��T����R>H�\>ׯ=���=��M>�X^��ǽ��G��.=���=��^>��?$n>�(�=%!�>����44��Q�>UB/>��">�=?��?�kd�p�ܽ%7���`�	�~>��>2S�>GX�=	�H��,�=6;�>��d>��T���|�)�Y��U>�n���1~������V<�e��D��=��=㴸�1�0�*=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿl��>�:�����Ƌ��@c� @�=���>��M?w ����<d�c�Η?��?�B��M���gпZPs�bA�>?��?��?�i������I3�� �>o2�?��,?�ԃ>�j��c3�I��>�T?7�c?�P�>ާ(���V��V+?-u�?z?�hH>��?V�s? ��>����93�W��~ߋ���=�M><��>�;>a��j�C��3���6��:=k����t_o>�~=p�>�DԽg��n��=�Jy��A��"1Z����>�[>��J>Iߔ>M� ?*��>���>j02=ˊ����}�����'dE?[đ?O	�~s��3��S?>���^��>�+?1��Gj�1��>Cw?pU�?��U?�9�>Z�
������������2a�<�PK>b�>P��>돽��>�-����Ѐ�>.�y>V{�=n��H�P��h&<o��>:Q?��>��O>�= ?�J%?Gj>�8�>�I�6���E�d��>�:�> �?2�?�!?K���20�nؓ��Ƞ��X��Y>~�v?D.?뺔>~������,����:�~]���?�c? ɽ��?gI�?�*@?|�C?Mtb>��)��-����Ț�>i�!?����A��c&�h4��?�I?z��>?�����׽c�μ��������?L!\?�;&?����&a�@þ+a�<�� ���U���;u=���>�>ɵ���ƴ=�>�w�=�/l�_a5��,k<��=Rv�>X��=�R6��i��vB1?4�Ƽ��l��>�Gs��q��ls>{�g=H����-m?Og�\�U�����%I����e���?���?�h�?�
��:p�9�f?��p?���>-?� ̾I+��Z��e� �8y���ež��>q�?>ʎܽ�V��֠��룿G�h�2 ���	��>���>S�?�� ?u�O>?��>�Ř���&�I�����\�]�|d�~�8�;�.�
^�u|���!�u��>¾��{�fL�>�[���n�>�	?�ig>1}>��>W���mE�>��Q>c�}>�M�>�Y>n3>�f >���;8�ν5R?���~�'���辐��B?�d?D=�>%�e��z���g�1�?3��?My�?��v>�h�-+�� ?n�>�9���$
?i�?=���ۘ<s����]��������>Tٽ	:��$M��hf���
?�?�}���*̾��׽	����hn=�F�?h�(?��)���Q��o���W��S���/h�����$��p�p㏿�V���"����(�R�(=@�*?W�?2����} ���k��!?��kf>��>�"�>�Ͼ>�I>��	���1���]��?'�𻃾�(�>;V{?�>KiS?I|:?�@!?�-f?D1~>ɸ�>��r��?<ù���>�	?`H?�H>?yun? "?��>ɱ�=(���P��{ݾ�5?Z?k?ps�>�g�>ɒ�`�;dFh=��=N��_T�4���R%�>�9���7�=��	>ZW?U���8�I%���j>��7?���>���>˻��i�����<���>�?}��>����<,r��c����>L��?�~�v�=j*>��=�lw��l ����=|���=��y��<=��](<y%�=�z�=.a��e����:*�;�}�<���>�	6?˲�>���<޾�=���M����>=�>��>���=J��; ��b䍿�}|�*R�>��?�(�?7��=�c&>& >�kξ�H��$�i0����O>ɖ6?a�??�>|?
�?�O?>�?�h�>�?	����� ���\��?Q,?��>����ʾ�����3�Պ?�r?�a�P���#)�zp¾Rս��>bB/�{M~� ����C��%M��������.��?xɝ?�>� �6����;ɘ�䫾!pC?���>�o�>���>�)��g�k��5;>��>��Q?�w�>X�P?(_{?�\?�G>�\=�W������u8<�t)>�8A?S؀?�B�?T�v?���>F>�O6��Y�K��&�N���z�=O=��`>�(�>��>ܩ>(��=d_��������O�$ܯ=Q.f>S��>���>���>��u>��D:F�G?E��>z�����Rɤ�Z���U?���u?��?�x+?�=�]�gF�;P���R�>�T�?���?�,*?�T���=/ּR}���q���>;Ϲ>��>i	�=��D=�2>&��>	3�>��@F�2t8��lL��	?#F?o�=;�Կ ��Ojλ��<�~�:�G�� ��)羒����;���'��U��!��=S��ʓ��-��|%��\-#��1�%��>5�H>�7�����EK�=d&z;C7�!��=�l�<�����-�	�&={�l�t�<2lȽ�3	<���;�#p�5�<[�˾��}?\=I?��+?9�C?y�y>�>>\�3���>~���??�V>�xP�����};���������ؾft׾v�c��˟��E>�MI���>t23>�6�==�<X�=(s=�ю=�}Q�4=�%�=>L�=�f�=/��=e�>�Q>�6w?_�������4Q�/Z罨�:?�8�>1z�=ہƾ`@?��>>�2�������b��-?���?�T�?T�?[ti��d�>!��j㎽�q�=东�G>2>n��=��2�[��>�J>����J�����m4�?��@��??�ዿǢϿ�`/>a�7>{�>aHQ��%1��XZ��\a�}�]��<!?��:�@�˾=��>�=S��}6ǾK�4=��4>&1s=4,�z\���=��y�`�N=+En=)�>+C>���=�Z��n$�=�D=C��=�J>^�#@.�I4��[6=���=n�a>P%>Y��>��? d0?Bd?F�><�m�IϾ�1��x^�>��=(1�>x؅=DB>s�>R
8?Y�D?5�K?z|�>�R�=��>�>�|,�Y�m�i�徂ʧ�N�<��?<Ɇ?���>r�N<�A�����]>���Ž�n?�Q1?�Y?���>�U��࿁U&�h�.�����}��d+=lwr��YU��������㽀�=�q�>���>J�>qHy> �9>��N>��>ݲ>��<@U�=E7����<󼔼稄=�ϑ� �<E\żR��	A(�^�+�Dt��
��;օ;��]<?i�;/=>���>WϠ;#�>K>�g�s��=�1���=1���>$.�WM��4E������0��5���j�>�>�H�D ���$?C��>FW*=o!�?�gM?�J�=X{]<�=о-���߽R�뽻)<��A�=Â��_V��~�̚C�����Y�>���>���>Y�|>TG?�0�N��M=�ܳ�Xx��?�n��� ��>{�tc�(w������oh�ę%�'KW?����؇�=7{?9�W?E�?��>�Z�?V�}�>-���(�<� ��9�|@ý��,?Ό#?}a�>�K�5�6�zH̾+���޷>�@I��O���^�0����#ͷ���>������оv$3��g��������B��Lr�Q��>�O?��?k:b��W��CUO����6(���q?�|g?�>�J?�@?|&��*z�kr���v�=�n?ĳ�?E=�?�>0��=�}��Ew�>P	?���?��?Us?GN?����>j�;�� >�ޗ����=b�>��=7��=�A?\d
?�
?�坽��	�,S�T%���^�]��<^s�=�>�>��>Axr>���=�hg=�@�=�\>쉞>�>�We>Ȣ�>%��>)҇�ޱ��?"ԍ=��>0�?-��=w5E>�L�b��=;Z������c%0���l�s�(��)�=�2�=T���m�>ڿÿfc�?Ṳ=>�B?�M ����>�=��~>}�t���>?���U�>S�>Y0�>��>�X>Ɍ(>Zcھ�>u�	�d]#��K5�ÝI��_˾v>�r����3��F��` �'l�B��}� �G�f��Ղ�h*E�B�?<�~�? ���d�o�ǻ#����<�?��>��B?����;Ľ�.�=Q��>j�>�澟���IL��}�ݾ؉?Bw�?��j>��>/�Y?���>�v
��%���bt��IY�-1.�=;T�~�S�qB��7.��k�
�\�C�P]H?�a�?F:?��b�J>V��?O��PY�ol�=sFK�1�=��ғ=Bў>����]�þb&���#��h������y?�b?~)?��]�:������>V�|?�I�>�11?���>4?��?!C?D�>-u�>{0�>]=H?m4?D�l?%�>�����ﶽ�^>LB�U���R�*<�RX�������ϼ>��<����L>��=ĵ��Jl�<k��=DR���̆�,�=s���L�=pK�>�$]?�+�>��>��7?��48�mB��R\/?�8=|��.'���b���U���>x�j?�t�?�VY?�b>>�A�U�A��>�f�>��#>/y[>�X�>����l_E���=[g>�r>Ƥ=��A�n����c	�p��]Ƚ<$# >���>��{>�+���(>����Dy�A�c>��R�g��(R���G�k�1���v��"�>�K?�?���=�d��֗�:>f���)?$0<?��L?��?�c�={ܾ��9��J����>� �<E!	����������:�$��9̊s>�I���꾸�9>jsپ�Y'�~Gr�&�p�Ȣ�����>Q��Ǥ
>v	��3��{���u��>�>V菾�����GY���L?�Q=�^����`���&�y�z= w[>�]�>9��
og�FEK�����x�<���>��A>�ʹ�*I��N�H=�n)�>�'E?f�_?���?�v����r��B�֔���^��m¼��?>T&?��@>�=�=m���%�e�0rF����>�t�>2���G���������#��e�>e\?��>̛?��R?`�
?ra?�*?�?Nސ>����S��ǀ!?�z�?(�R=�뽍�*�r7��Q����>�<$?�Fc�[ː>��?߶?#?W�V?V� ?�q8>?%�dZ=�芑>��>]�Y��۱�P�>4nK?g��>VBV?�?��]>�|1�搏�.�;.�=w�C>b]1?�� ?Z�?���>Q��>n��0$�=gy�>�
c?5�?]�o?%�=�?yB2>6��>��=�L�>m�>��?5O? �s?�J?2��>Tm�<�d�������r�NwO��@i;�G<��w=�+�YCt�D����<�ح;k���������LAE��Ս���;m�>�Y>�ٓ���+>,վ�K|���D>����␾�*�����Is�=Q9�>��?��>��/��V=> �>6��>�|"��#<?e�?y?���=��k��%������>g�B?���=3�k�����V~��I�<Ld?j]U?j!T�t���i?˼L?��W���}
���̽P��(F`?���>T�.��?s�}?��h?� 
?!�	�g�l���o��u���>�Qy>i�C�Lew��?�>�J=?�ۮ>q�>�#�>�#�!�c����m��>ص�?�A�?��?��P>#K�u�࿚��(7��+c?`D�>򬙾?�?< Fླ'������.�޾x���7�������2��#gP��<��Lg��喟=C)?2m?�|?��P?�@
��X_��l���l�1�N�M���)�PH���B�mE� ~f�uM��GǱ�����	�=omy��K8�'��?��0?��3�om�>롙�$���^پT�U>=���,��;��=�[ٽ&�H<i=��c��Z<�zޱ�&c?�T�>[#�>v�9?)]U���7�h
1��3�����1'>I�>S�>��>OZ���1+�����(ɾ�������O�u>PUc?��K?��n?w����0��x����!��5�������A>��
>�|�>� Y�ë��&��!>���r����������	���=n�2?o@�>D��>��?�?��	��K��2�y��71�v}�<{��>V�h?�I�>��>'GѽȬ �?�>�)j?$��>GA�>�x�����T�x�.������>k,�>v�>��X>qH-��^�����ڈ�h`0�#��=B�^?ީ��d~�@F�>��T?��g;�;=��>�xƽ,�*��ؾ�Qd��4>j+?%}=Ә3>��Ծ���%c���ԅ��e*?��?TG���V)�8N�>�z!?9Y�>�>y�?���>�帾�Ď<Fj?
�\?(�H?�>?,A�>��<g��EϽ��"���7=��>��e>�G=�=X�%��X���_)=���=�����Ž�T�:������<b` =î@>�߿ν@�_4����%y�(�������U@<�e����eA���฾LU���3ֽ;L���p8�9A��T|���I��|�?ګ�?^�q�,U����o􃿚㱾iU?��Ӿc���hM������ޝ~��݃�������uF�綈�/ry�0�'?�����ǿ鰡��:ܾ! ?�A ?�y?���"���8��� >�B�<+,��۝뾨����οY�����^?���>��%0��g��>֥�>?�X>�Hq>����螾4�<��?&�-?��>͎r�(�ɿZ����ä<���?0�@X�C?b5��`���=�S ?�?�9G>�Q���_������>�#�?AI�?ٺ=TtO�S��5�X?�V�=�E�LX����=�ٳ=�S�<C[H���$>���>%��CO�n{� �=���>�s�����b� q�<�ZX>Gλ����5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�}��=[��>c�>,������O��I��U��=���bs��"]�� �1Y�&�
� ޸�5aʽU3c�0��;�
��wޔ��U���*=֏�=��4>(M�>�Ӄ>�@p>��S?��j?��>��=m��T����!����x=<����B��~����K(��[���wnʾ����!���v"�4�ξkOD� �=D3H��y����'���f�_�>��'5?�x>^��_G��x`��,ɾg��)�����Q~ƾ�2��m���?��B?n���X�X�O�	������]�]?�t �&�����T�>Vf��,j�=E.�>��=|��*@��n]�m>?3�?,����W���>�	�%B>��0?;�?��7>�Q?')r?Dϡ�5�����=�i�=�P�>C\,>��>���Z���n?��5?�lu�i�־e�{>U�Ѿ_A_�*+>� >�^���${��9>>�ѽH�S�{T�<�f�=�t>�(W?���>��)���`��p��b_==Ȳx?�?e.�>�{k?��B?�Ƥ<g����S�j��cw=��W?�)i?�>����о����2�5?��e?��N>�dh�h��p�.�U�d$?��n?�^?���^v}��������n6?��v?�r^�`s������V�T=�>�[�>���>��9�El�>�>?)#��G��غ��mY4�"Þ?}�@n��?��;<����=�;?U\�>e�O�H=ƾ4{������v�q=�!�>����ev�����Q,� �8?��?���>(���ש�Ƌ�=Jѕ��[�?!�?����Lg<.��l�0n���O�<İ�=:�j:"�����7���ƾ��
�񟜾/ҿ��>�V@�����>n_8��1��TϿ�
��l\оXdq�z�?�g�>M�Ƚ�����j�>u���G�G�H�!��� خ>e>Lm@��[r��怿��0�Z=q_�>$܋��>=p��~D���1����=쵈>0��>��h>�Z��K��y�?;����տϘ���g�j�]?Z�?��?�'?�+�sxR���k�hy�<M�O?:z?2�S?�RüO5X����%�j?�_��xU`��4�tHE��U>�"3?�B�>S�-�o�|=�>���>g>�#/�y�Ŀ�ٶ�>���Y��?��?�o���>r��?ts+?�i�8���[����*�u�+��<A?�2>���H�!�B0=�UҒ���
?V~0?{�e.�Qe?~��w{��1��l]=

?�@��6p��g<��	�C[G��;����m�八?o@_��?�N�p#���)?,��>}T���<���Y�=���>��>B=Őͼ��>[��H���B>l��?��?���> ���#y��d� >Ղ�?3��>��?���=���>�1�= :���{�
�%>��=':�!	?��M?�g�>r'�=��7�.�.��E�4MR�2���C���>'�a?�!L?)d>
~��i�6�Z)!�3F̽�/�	��@)?�Q2�lRὄ�3>��=>��>n^C�x8Ѿ-�?ao���ؿ�h���p'�;04?F��>��?|��I�t�����8_?s�>j4�-���$���B����?7F�?�?4�׾�}̼�>`�>OS�>HսR⟽�y����7>=�B?��4D����o�J�>��?��@S׮?�i��z?&)
�5f���Jw�/�쾃�)���>�&?�7�����>�*�>	I5=��w����|�w����>	n�?���?�q�>� �?���1����<k׬>W
�?��>!FN:����S�=��?�� �ƻ�����w�?:�@bk	@��O?����ڿ|&����t���G1��;�\>���!i;>��<�b�;z�����=+k>�@G>�=a>��F>@��>���>i��%���Z�����B�N��'����NN�Z?��Y������� �@��2FI��%�7���5l���d�<KΘ��{�=2pU?��Q?�4p?	� ?�gw��� >���4� =��#� ��=9	�>�C2?�bL? f*?t��=s-��t�d��B�������ȇ�#f�>��I>���>���>1�>��,:]J>?>�\�>� >Hj'=�����=-O>*�>?��>+(�>�*7>�p>���dt���h���}�YV̽6T�?�w���'I����RF��t���n�=0�-?Y>����aпT���C�G?�@���~���(��=
>yG0?��V?|>	���m�S� �>�8��}j����=%.��k��)��R>c�?��;��(>��l�U���3���6
{>��J?�D̾�)�hg������{�>��>eC =V1�q��c����^�`$_���?�"?j�Tk��ؽR��/ג=R>>O�>/O����M>�yH�6�g�zx\�;��<��P>hX�>�U?4>�mo=:��>s
����X��4�>�L>�y3>WB?*?�L�#��|rw��%2�wn>e�>�@u>.�>��K��Ǯ=g7�>�&j>�����x��BM��><�n�S>E�K��S�)�r���y=Oڎ��=|l�=п�6x8�$�,=�Yz?�g���^��>������>��?b�>��=n�=������h�H��^�?V�@%�?T,�9Y��\7?�s�?�^��=�A�>�t�>�Ю��Ѽ�8f
?8�<v�־������C�?��?N�0���x n�~�C>�/B?	��R'�>;��P��W����u��d!=m��>H?����I�L�=�=�"`
?q�?H*�촤���ȿQzv����>Y��?�?��m��:����?���>���?�AY?(�i>?4۾*�Y��e�>��@?'�Q?t޶>�(��7'�?K�?���?�F>U��?i�w?�>@�~���-�ب��7|��S�1=�2�;��>�>D���H�ۓ�!��Tj�/����_>��'=Y�>�۽�a��V�=d��������E�|z�>'g>�S>��>���>�>�ŗ>� =����n�zw�� V?��?D��MY���S��">т��s-?�N4?�1��U?M��4�>1�G?��t?X\?
|>��!5������I���E�=�$>���>��?�Խ�p<Xþ����ݡ>��`>w"=J��?G������O�>)�$?���>�ރ>��?�P?�>�>4�?tYN�- ����"���>x�e>��?u��?}�?Ȯ���S&�ތ������Z�[�wC=&?��4?���>�����ܠ�lL�bN =,S>�S�?��n?����oG?��?UH?"�q?�O�> ���׶�G��(�>@#?��
�F
B���$����A^	?��?@M�>)���X�ڽ_�U�PL����_L?�Q\?�$?�
��a��Ⱦ��<�R컒��c4[:{�:-�>sR>�z����=q�>s�=��h�K�<��\<��=��>�\�=� 3��Z��|"?f�=g��(!>��l�-4<�%�7>#u;>q⦾�{N?Wb��aqx�iD���%���	�?��?���?;[��\��)?@�?/B3?�}�>k�O�3aľY(
����l�F��^0��
>���>5������g|��N̬��T��\���#�[(�>��>`�&?��?(�U>s��>Z�$�<�#��� � ��g8���վ]�&��l#���4��\�;WŽȶ#>W̾�ʃ�_��>:؆=�ԡ>���>�O�>��>!I�=SS�<��>o�K>�o0>�s9>@)>��1=�ͼ]\�f,�O5Y?�*%��(��r��F1ܾiY?�w? :�>'B�Lg���\�q�1?)��?톢?���>9�g�%%�KG3?,�?�͑���??��>�rϽ�����˾��������=z�;��S�Qoo�Ż}�6=��M
?��?n1��[e߾`v=�)�����=��?eN?w�!�N�<�s�i�1V��Yt�G�:@=��*�����/8~��̑��
���À�p2����=�,&?��v?.����DѾ�q��J-c�����>	��>`en>5�?�O�>�^꾵��LF�"��{���ɍ�><̈́?���>��I?5�;?�vP?�iL?��>�f�>�/���k�>���;��>�>ޜ9?-�-?x20?�v?�r+??0c>j��H��e�ؾ�?��? G?�?K�?�݅���ý����f�y�y��y����=���<-�׽�Au��T=�T>�S?P��Iy9��}�kՉ> �(?���>G��>��n��Z���=:�?�n�>�M�>�]��%�f�$(����>X|?+lA��"�<S,&>��=��>���9��>T�6�g8=­7<�!��m�<��=��=�޼���9�D�ʅ<�w�<�J�>�� ?��>�>օ�+��#�Iz�=y�^>�}J>v1(>,۾=���W,���g�l��>R�?�Q�?�G=`)�=9��=�d��r��L	�_�����	=�?d�?�yU?>��?�:?��"?|>�o�Ye���ȅ�������?�,?;��>J��q�ʾh憎�3���?b\?+<a���:)���¾nս��>+[/��*~�$��D��S��h��L���>��?c��?�'A�U�6��p�R����^����C?o&�>�O�>��>��)��g�)%��0;>��>�R?f#�>w�O?�<{?�[?�gT>��8�p1���ә��k3�#�!>z@?���?��?y?t�>��>�)�V�T����������EW=�	Z>��>(�>.�>:��=�Ƚq[��`�>�8`�=��b>>��>���>��>��w>S�<�4?y}?o�ξ��*�%)�ځ`�����Y?/�?/�
?R��=G/�Y�A� �'�>OZ�?fݲ?�
?1ރ�q�=N�P�RH��~�[�C׏>��>��>�2�=A>г�=u��>��>ԑ�4���>�U垽��?�/C?,TI=�]ͿyQd�9w2�ܩ�����~mƾ[�Y��v���{���f`><�������*��6�O�ݽɾI���Ĵ���VR�~������>���=Q��=��=	�O��l<$%�;
P)���e��v=Sd0��M�����;]=��AL�Mhǽ�rT��`B=9OJ=�XǾ��j?t�.?a4?2QH?��x>�ʇ>�h%���P>�q��TQ�>p*(>O� ������b���о�tվPw�����$k�7ղ��+*>?�<�h�=[:
>K �=ʇ=�l�=��	>%��=ű�<��K=�P�=��=��=�(>/� >��<iy?y���Af��kH����8!K?��>��@=�̱�^v@?��X>����Զ���|����?zS�?'��?�F?DRl��y�>ׇ�����w�>��=6��>dIt<<p`�}�>.ϻ�A�?^����<$��?ّ	@X8?nj����˿A�O>$�/>�Z>ɬP�eq3��UY��Yl�� Z�HC#?a9�n~ǾE#�>���=O�߾�n���w:=��9>�wM=�%�p^��֖=�&���8=��~=i�>��D>��=hŽYn�=�gH=~S�=��N>���ʗM�n[F�n�-=�/�=��f>)>ES�>�l?Z�.?�Jb?c�>Q�p�r�Ծ�)��s��>%��=䓯>��h=��>>�-�>��8?�F?-�L?-߯>匄=�&�>Ա�>� -��n�@J�X������<��?��?��>G4<�q<���D{>��B����?��0?��?<*�>;��D�ڿ���dS,�� �db���$M;��m�;�1=G~=�C��4�/��=��>Q��>�Ҕ>�7�>,x|>�	i>�]�>��>��=��<�_��%��<o� �M��=��J�`=�Ҫ�}�f�$�;3��g� �i���4�f��%<��B�U��=p��>7Z�>Yf?a\�;�c���=ǯ��Y�N�ب@>0ޤ�N:��>T�+􂿳v;�@8�h�O>�x�=t#������@�>�-�>n�v>�$�?�s?�K�=�g�v4�ѭ��ćɾ����^�=�@C=�&���K�1�j��\X��#��2��>��>3�>�
m>1�+�~?�وw=fU�gS5�?��>䛌���,��.q�X9���럿Si�r&κ��D?B�����=>~?��I?�ݏ?���>����ؾs�/>�����=h��q������?��&?�C�>�(�g�D�&�ʾ�{��q{>�Z_�R�C��Q��mt��A�"������>����輾K[1�{i�������C����ZJ�>O\P?�|�?������w���B����؎�=l�>c?���>��?|�>=���� �yk�����=uq?Q��?���?T\>3��=������>�S	?���?���?��s?��@�.��>��R;��>`����z�=�u>��=F��=�?z
?��
?������	���F��]^�'9�<H��=���>/�>@�r>��=�g="4�=��[>ب�>ԏ>j�e>�֣>˨�>�ަ����p"&?�V>��>�y.?v��>e\�<������<8Oq���6��b�#���@������~Ѽ�hc=�����>�q¿�F�?�9W>�P
���?Y� �l�wS>�U>�W۽{��>D=>2g>r��>�a�>s�D>I��>�*>�`�`9�=g6���!�?�i�\�3n��9L0>�U;�-��ˌ���L
���L�n����z� �c����҇B�Y�,�c �?����Nl������*?�5�>�I?�����<��>���>�n>#y��~A���R���＾tE�?a]�?=<7>�Y�>��`?r�?�?�򽆾Jke���]��:���k���1����`.d�	Z�k�V���X?5�v?@\/?�-�=I	�>��?�b<�:�����>(L%�ߘk��/,>1�>#�о6�)D�^�¾����G��>砒?���?q�>5W��LZ���)>KL8?�O1?H�s?F�/?<?g��a$?�Q8>�?�&?$3?ua.?aY	?�->�:�=H�ٻ��8=_̔��b��64˽ek��	q����"=R~=z˴��
<��'=���<.f鼡�м@y;�[�����<�
B=�	�=v��=@R�>+H�?�bs>XG����3?G�0�Fw�^���d?q)�oy�<B���vIʾ��H�{�k>�}�?x�?m�"?]�2�c��6�Y��
�>���>4�y�4V$>f��>�;������L�=�΅>U��=)�9=g�v�����1/���m��a >�f�=��>��p>��Ƚ��0>�@��Y߁�W3>	!�H}����ؾ4�h��'.��R1�I&�>�=?��>���˜���<2q�RX?��4?=4M?-^�?Њ���׾m??��0����=�g�>ې���D�S������3������/>F`I�n�߾�
2>���ݛ���}�]�V�|ﹾ/�]>.���>��񾳾�x�ٝ6>�Q�=0T������k���q��g�H?��;U���y�@�����<�U>���>t�x��@l�A}P���E� <G��>W�2>����R���U��V���>��D?
�`?���?C���_is�B�s������e�K��?i��>�p?786>[n�=/������Zd��0E�H8�>���>b��*}I��ţ�|�!��m�>�y?��>��?��R?a�?A@b?!�(?�y?���>S�Ľ�Ŷ�-H?-M�?�	=t�_��<#H���U�:��>��"?cԟ�!��>'�>��?��?4e?h-+?�� >����*��И>��o>a^��?���Y>��G??��>jB_?���??'>q[(��닾����Hr={!:>�7?�V?F� ?vm�>���>����N�="��>w
c?�/�?`�o?d��=��?�<2>Q��>��=���>ϋ�>�?WWO?P�s?q�J?���>_��<8��
0���6s�[P�~��;��H<��y=u��z!t��M�V��<��;l���V��G��M�D�@쐼���;��>�7>���Y��>c����I����=[���~��;U�������+D>uÞ>��?�3�>A�3�ۅJ=%�?E�>�\A��W{?�l�>��1?ԶS>��g��a ��D,���l>c(Q?�*=po��������ǡ=Q[S?��E?��;�y����jh?ϝP?��1����q����*G��nY?��?��+��ܶ>�-y?��|?Y�?�=��Dw��~��{p^��)��Q�>��|>��+��a]�}Qj>-T?n1?�͍>���>)� ��R�˘��qx?k��?�Z�?�5�?��A>;�[�B�޿u��x=���^?Q��>��� �"?�����Ͼk��t��8�|��r���b�����r�$��؃�}ֽ� �=�?�s?`q?h�_?,� ���c��*^�����oV��
����E��E��C���n�,T��,��^��p�G=�,�o�>���?�*?UC$�^�>ۏ��!��^QҾ�U>J���͓�=#����=�Y=�i���(�h��PY?��>�R�>��<?S:W��g=��R.��6�=��b:>>6�>���>��>��9D80�@r��r�̾��b濽i1v>�wc?��K?��n?ik��*1����ޘ!�4�/��Z����B>�k>���>'�W����8&��X>�m�r�����y��|�	���~=��2?-�>s��>�M�?�?,~	�i���hx�/�1�ڃ<-�>bi?$;�>�>�нE� ����>ǧk?KG�>^#�>������!��|���ʽ`B�>�i�>��>{�n>g/��]�.�������\8�1�=�f?Oc��1�^���>�R?Z��;�<�:�>ISx�nw#��4�2�'��]
>��?y��=_W7>�$Ǿ�3��z��w���+?�?S̖� w,�?��>�?���>���>���?��>𵾯�G<(
?��^?2�F?�9?.��>��|<1����Ͻa"���'=V��>(�`>~C=o�=�$��Z��h���9=�<�=�r�[˹���:rx���~<�
=�7>�2��5��߷�~.#��	�,[�R��T�k<$T��MK��;4r��ZA�p���d��2��W�K\�T4���?��?Q���ՙ �OP��}���bվ&�?"a����0=��
�Z��?馾���*Q���� ��Q7�!v��	]���'?����{�ǿ�����;ܾq ?�B ?b�y?��c�"�F�8��� >B�<���Ǟ�X���d�οܧ����^?���>��z7�� ��>l��>�X>�Iq>����瞾>�<��?Ȇ-?��>Y�r��ɿʊ��6ͤ<���?��@j�A?G")����U=a��>h�	?�,@>��1�+N�=g����>�G�?�,�?rwR=R�W�:(��3e?�<��F� �h��=���=��=Ԅ�a�J>Oq�>4\�dA�`�ݽ�5><X�>�g$�����v^�OS�<q�]>��ս���8Մ?Y{\��f���/��T���U>��T?�*�>�9�=��,?47H�f}Ͽ�\��*a?�0�?��?�(?`ۿ��ؚ>��ܾm�M?KD6?���>�d&���t�Ä�=�9�V���`��'V����=���>Æ>�,���~�O�	K��d��=����:ſZ�"��J��l�<'�;�^G���SX����K�-ؙ���j��޽̒e=���=��N>'߄>*�[>��Z>��W?�j?�L�>�\> ���G���eɾ�U�;�ă�:�x_��p��b��>�#�ܾ�t��|�:��cȾ͌E�If�=�LK��듿h(��b��R:�v�5?�>�7��I�J���<Gľ�ٙ�D�h�Bz�� DǾ�1��Uh����?��7?fQ����W�^������B׽�g^?�������Ⱦ�I�=&���h="�>i�=G�ݾ
;�5
W��_6?�%?ꁳ�﷾��v>n�D�<�_>R�?�?���=��>a�)?l��d��=O��=!5�=��>�b/>VU��㯾k�
���&?�qI?=��I�m��^�>�4߾������m>!=�=J����b�ê�=К��oI�3��<�N=ޕ�=�(W?���>��)��0a������Z==��x?ϒ?	.�>r{k?��B?�Ӥ<�g��\�S����aw=��W?�)i?Z�>Ǉ���	оn���b�5?��e?��N>�bh���1�.�YU��$?��n?!_?����w}�o��W���n6?�|w?��a�����0�8bI���>>��>i��>j�9�	�>b??�"��y��"���4��7�?}�@�I�?��<>�y�A=��>���>gDB��`���p���꺾��=���>Z���՝z��I���"���>?,?�?���>����������=Lו�N[�?��?�~��0�f<���-l��r�����<���=���N"����l�7���ƾQ�
�����;⿼���>\Y@�W��'�>�B8��4⿔QϿ����\о�Pq���?߁�>;�Ƚ������j��Pu��G�9�H�z������>=�+>���b	��*-��� /���r=M��> �ϼ�>�9*����i�HkL<�2Z>��>e�I>���M��<�?�����MԿ�ş�3��*lq?���?�:�?��A?���c���mb��l�=>�a?��?1MH?��L�P�����j?�_��nU`��4�`HE�U>�"3?�B�>Y�-�İ|=K>���>�g>�#/�o�Ŀ�ٶ�H���[��?ۉ�?�o�,��>r��?Xs+?�i�	8���[����*���+��<A?�2>����L�!�00=�4Ғ�ϼ
?d~0?{�g.�1�i?.��X���"��Q�=��?��n��X����Ž{�a�O�������c���?�y@@f�?v��6
 �c�?x>ٳ���١��e��T�>��>��;=����>d>&���2t�	7$=U��?�I�?�?DY��.����A|>���?�F�>0|?^�w>��?�`��T�Ⱦ*�.>6�!>�$A>���=)'?�@?睛>j��=b*u�4P��?3�%(<�${��O����>��e?-+q?��T>��k<W{\��S�4�A�Wo��3��=�"�l�>�MJ�ԛ@>�z�=fV��Y�B�G�ɾ<?UG���ֿ����+�mK0?G:�>Y:?�%�)1g�Ri���_?�ۄ>�W��Ӵ�n���/� ��H�?+	�?�}?w�ݾJh$�$�
>��>�&�>KU⽦���!���9>&5D?�L�����q�p���>�.�?�%@3v�?��h���?S?�`k��o[���L޾��(�4]/>�-?f�	��}�>�Q�>K�C>w�s�߭��c����k�>{p�?�#�?o�?I'�?�>��:\�TL�=
B�>�Ń?M�>�I��NȾ��+>��?v�!�("��Ž�^*l?�@�C@MQ[?�̪�׿%*��YU���9��x�w=�V�=-��=�����=Ł[=� ="IA=�}>~��>�oJ>��Q>�$7>�;>]|%>�F���o�DM��l▿��U��
"� ����`�n�
�?��c�|-���U��@'����ѽxי��U��Q@��A%����=��U?:�Q?��o?�n ?dcy�W  >�@����=�r#�.և=ik�><+2?�}L?X*?8��=z͝�B�d�`[��1i���������>�
J>�/�>�Q�>�ͭ>���0I>u�>>���>3� >��(=Q���d
=��N>�
�>���>�T�>�!;>sN>i����2���h��w�he˽��?������J�d*�����I������=1M.?nf>���??п��4H?�Ԕ����>+�%>��0?�eW?��>����V���>���Vj�=>Mj �9m�,�)�h�Q>y�?��=_�F>�]��ZH�ZZT�`0߾�{�>��J?�ѿ��Wνnu��-��:ᾓ,�>(�>5����z�E)��������q��!�=2�-?J�?[��c��PG(�T���L�>��>:f�=�+�=\�@>��~��]�k���Í�9u�>�Ў>�L?E�D>�ĭ=�>�����e�r��>�=>|S>�TC?�	(?"sW<D��.�L�@�U��h^>���>�eY>�I�=��f�Kp�=�Q�>��>g���G������d�&�؀0>�1м��P�撽�yx=@Q���=o�r=s������B<� �?�pĿ 핿qھ����>��b?���>�������m�\�������o��?�@Ą?_�-���N��P?dږ?�퉽l�>S��>�p�>�J�2���F"??�J�Ҫ���]C�
��j��?�?\E��͓�=�R�t��=x�4?�侦P�>��#�l���҆���s�K��;;_�>��G?�+��3�H�?��?L��>!��"����8ƿ��s��\�>'v�?oɚ?��q��?����=� ��>�$�?��N?@YJ>r�۾i>��r�>��>?��C?��>����
��G?��?��?��8>Ȥ�?��z?���>84���3�Ҵ������m�-<,x�=ԡt>��>Ze���{O��ӓ��j��?-g���� �\>Ҋ4=8�>���\��q��=\m��I���0�N��>T�d>�]d>�!�>�k?e��>'�>��:�����[������%�Z?��?	>��ak�M�<��>%�=Ȱ(?*�R?������	��|�>G/3?.�{?�PJ?��>o��������J��F۬=��=�~>� <?@޲��"���gž��@��*>>C�>p�����SN�����V��>u�?ǳ>��&>�?2�"?��>���>�4��莿i�.��ú>%�>��/?�[?N?Tw��d?����������:T�s��=�kg?R�3?��>��Sb��f�v��=7x1>�R�?�!�?wF����0?1�?.�K?F=m?VG�>Q|x���ɾct�N�:>��!?nyٽ�@�Ϭ#��Y��>?u�>׎�>�a��a��b��������t?y�c?�U,?B�����d���þC(=`�������h2<�����*.>�f>�#Z����=�1>5z�==Uk�wO�1�I��j�=�3�>&t�=��#��ڸ�H�?[��=E���!�=�:o��<�Y��=��>`��wY?��9��Xo��M�����k�냁?;Y�?��?.J�n�[���>ұ�?�UB?/�>#����E߾��#���)��p�=�3O���>�{�>�ֽsCھ-G���F����m�E�Ľ�锾\�>KQ�>&C(?/�?s�c>fY>�O�f
e�AlξJ�(�;C�?��q E��'�rU!�g9�l��=Bt#>�Ϭ��B��
8�>Mq~�2c�>#	?��>�A�>'�">�����b>0`>Z��>���> :o<S|�<<�Ѓt�Qo:=��Z?���E�,���Ծ���}UW?�(g?LN�>�vS�ި�����H?�l�?��?::S> ga�0�"���?5�>�����D?l�>0��<�9ü?շ�/�l�J���B�;RW�>���U�!�k�u�j~��XA	?S� ?҅�=��;UD��n!��)�=�h�?�%2?\��!�U�'Ol���N�=�\�t*H=~���ٕ����z����/��&��8�"���@=gM(?���?n_�����޸�̰`��')�q�r>���>��>���>�[>w{���Y��:[��,��������>�x?k��>�I?��;?|kP?�`L?���>Ot�>(��t�>ً�;��>e�>��9?�-?)0?�q?�l+?c>Q�����y~ؾ�?�?�7?�?ح?�ⅾ�ý~]��7g��y��v��k��=ƚ�<թ׽�:u��U=T>s�?�h�:~8�����o>��5?���>F��>ʔ���Ā��=��>�#	?�> ���q�������>1i�?֟
�ʞ =�*>���=
������D��=@|�^��=��_�\'=���*<&��=�#�=�b��`â:�!;���;2��<��>�1?��>��> *��� �5����=��e>d�U>�>x�ܾK��7s���&f�>�}>Q��?���?�=S=4��==��=���%`����h����=��?Ѭ?9U?2J�?��<?Jp"?+��=�!�D쒿jヿ����?`!,?	��>`��[�ʾ��׉3���?\[?�<a�V���;)�¾��Խ*�>�[/�B/~����"D�����������.��?�?�A�M�6��x�ӿ��V\����C?�!�>'Y�>��>R�)�d�g�q%��0;>؊�>aR?R�>C�O?�%{?$�[?ӜT>��8��5��~ϙ��2��R!>@?���?��?iy?C��>�S>4�)��8�+���i��5������V=�Z>���>y�>��>JX�=8Ƚ�0���>���=)Qb>���>���>/��>1w>P�<cv2?E� ?�}���پT������� ���L?ݵ�?��=zU�<�$Z���g�V�#��\'?� �?� �??�>4�U��@�=�K9��#�;�d�9�>y^�>�o�>[��>��>�"�>K��>U�>\��`����H�yn���,?ڻY?L�8�l̿<�_�Y�;�^ ���������,N+��II=�>[��>!����侽v|��� �ў���y�]b��R����^�����>ni=hw�={d=�ug<��V�|�T=�C�=:����;�[ѽ��<o��}��<[�U�����SB���3�<B���@��q?��? �?Hv?Ǫ�>�}�=�d�xt�>b$1��+m?8w�>��=r����酾�^ξ��	���쾳� �h膾ec��@*;>����H�,>b,�>�Ѕ=����c�	>�B=,�)<��Q�ƌ@=��=Z�==É =��,=��=�!>V�?�)���a��G�@��3@=��Z?}�w>��<:Ѿ�LB?��>1���aȴ��<���i?�(�?.��?(?]L��g�>�EᾺ��ѠE>*�<�k�>�I\��ԗ��=�>IE>J:�\+���^�I��?&`@Ӑ3?�;���ۿc��<�/?>�*>R���2��H�Qkk�BPX���!?�4��;-�>Z�=ԏ⾥I���hR=t76>��]=��)�:�[����=`���>�:=�~�=�'�>ˆA>�޷=�K��I��=vZ_=�D�=q�L>d��aH�S�I���0=�|�=�e>'?&>�Q�>M?��$?��X?�<�>�?��D�Zƾ^�>ֲ�;�W�>H|k<��(>gm�>�F?�AS?�I?Ï>��=ݻ>%Y�>+�2�� h��N۾����8਻��?�B�?�%�>��<80'��� ��(>�Mw��_x?��*?�r�>w�>ig��U���%�[.�N������:��-=�;r�gHT�����eo�gs�#?�=�(�>��>��>u�x>x�:>!�N>���>-�>"�<��~=
�»��<�i���щ=Ȝ�����<H^ռ�H���%7��H'�e��j=�;W��;faZ<B�;���=w�>�bY>SG�>M�>JϿ�
8=T믾�P�J�4>�;ؾ��7�9�Y�7���2<%���"�z�*>�Y�>��n�hᎿ�t�>���>	-�>V�?T�V?��>�� ��^��O���<_�2<N�o��=���<?+P���7���m��Q@�֫�U��>hߎ>��>�l>g�+�,!?�1w=���d5��%�>����c��@�@q��:���쟿zi�^�ºۓD?�D�����=�!~?q�I?��?v�>^!���ؾ�/>�#��_j=j��q�������?!'?�g�>Z���D�m;�$��2�>N�t���K�4ԑ�g�+��<nž6�>�慨L���Tj*�3u��"��}�C��N�%A�>:f?F��?�e���̀��J����6��8��>k�R?�_�>�?z?���
��&���C�=��p?��?���?\�>	�=H����<�>+�?���?d��?�@s?��?�Y�>ԭh;��>ݘ��n�=2>���=���=�?˴
?�.?�����	�ʎﾓ:��]�\��<�N�=�p�>�(�>��r>�s�=A�c=S<�=?�\>��>���>�wg>/�>a��>�0����v?ɼ�=��>�8?�:�>�=$:R�D�$������8��[��^���=��Nc��z��09�=���=��>�������?)�=3a��[3?�A��<�;�>��a>>�ϽY�>��">�\�>�{�>��>�?�>Ob�> ,>R��[��=��۾��1��]A��L]��PE����>�b���@r����Z/p�Y*3��$V�n�f�b�y}��i7��0>-ɍ?M�N�� `��9�۞����?1�>~��>��w������c>iE�>���>�O��ؙ�F	��ӥ��0��?�@+>�ȸ>��D?�R�> �d�5����Eb��v��d7��ax��kW��2��T��{辂�t=|Z?�!f?V`3?i<J>9r�>qD�?gx9��`t���>�h�m�]�Hoλ�A�>�;���%�������ֶ���?;A�?�y?�.3>z�����f�%1(>EM:?��0?ōs?q^1? �;?�S���$? �4>��?��?�c4?�.?�	
?C�0>���=Ujػ*$=����;Ί�c:̽mcƽ���2=��=9~��xt�;�9$=QD�<�wܼ��;�}���:�<��9=#	�=A*�=�>�	Z?¶�>�iy>�@0?�{L��WB��>����/?��<�2w��b������:t��C#>��o?d��?��I?J>��=���C�,y?>�$�>�>��R>q��>g�˽]�a�,�>��>-�#>�V�= ���;���5�	����'g�<��>W��>2�|>=����h+>�2��߉z���a>xW�sb����S�U�H��v1��u���>S^K?F5?�U�=�w��C����f�2*?@<?�IM?M�?#�=�ܾ��8�L�J��.�
�>�Xk<��	�U��в��:b:�ou���r>i<����߾�b,>'���ֈ�t�y��y��&���y�=g8��l#>�n������뛾2>�=����p����pr����"?��<�m/�+�������5�>���>
�X>�Խ����fA�tσ��w=�N�>��6>�􅽌�ػ`�����>�D?��a?���?h���[�n��YC�J���*���Q�i�s�?�ά>q�?Jj4>��=i����`�p�d���C��Z�>��>'��h�H��G�������P�>��?p>��?bLS?0?A$b?
{(?W�?�D�>�����]����"?D��?e&=�[Խb��Y�?�d�L��f�>>+?NᒾCc�>���>��?�?C
e?�(?�f.>����*�t˟>+~�>��\�3����o>�M?p�>��b?�h�?��>�
,�G����xͽ�C�=��H>��2?D�?s��>8\�>L��>������=>��>(c?.�?_�o?½�=��?�C2>���>^�=/��>��>�?BRO?��s?(�J?���>�v�<�#���A��Xs���N�b\�;��G<�y=t���Dt���\��<̆�;�n��F������"�D�����v��;��>�9>�֎�Ѹ\>L��0HE�γ>'��T�������$~����>��>�+?d��>ad�1�|=��>��>^r"�ٗF?Q?2�?�7>bq�x �i}}����>u4>?q"!=R������r��M\�=x�c?̷M?ҭ!�L#;O�j?�N?DEӾ��*�t��_�Q��`�_?��?��½{4�>��s?�u?7�?�7��s� ֓�{zl��Ѿ{�
>Z�d>PR:���\�*I>	4?��?wօ>e��>�m⾨}�M3���?��?ǲ�?~��?�<#>�nM�{�ܿ����s����C^?�2�>񪤾j�"?��_�7	Ͼw� k��ə�����E���h������^�"����&�̽���=�*?��r?9fq?{_?� �9f�f�^��E���S���NL���F�N<E�-�C�2Jl�l��B��������8=d~�
3?��I�?�'?��&����>�ڝ�D�쾆8Ͼ�2F>�3������=�m����-=��E=N.i�M%(��8��� ?��>(��>B�9?[�%@�P�1�r�5��h�?�0>�I�>���>)��>0��<�'��Wֽ�������kٽ�6v>�xc?�K?��n?So�S*1�|����!���/��b��h�B>�k>%��>�W����$:&�nY>��r�!���v����	�ɧ~=�2?�'�>���>�O�?\?Q{	�l��jx�f�1�r��<�0�> i?M@�>S�>Nн � �0B�>��h?}�?k?�>gm���c�:���$f�%g�>�{�>��>�@>�E@�9qg��,����+75�e�=�re?R~�H'd�䬙>�F?�K�<���=�b�>4������n��A���bQ>�p
?"�=o�>��վ��d�z�#Mo��*?��?y8����)��Uj>kx!?���>�2�>�Є?W_�>�����;�?V#]?��I?Z�=?�$�>Z��<lӽ��ʽ �%j=�<�>�e>'�p=�/�=�b�
>^����W=P�=w��nͽ��<K�{���<�f= >>`H�#M���Ǿ�/��%!�5��ӁU��r̼u�Q��ﺾ�H��)y�����_���X)��So�(g�u����?*u�?���!Y�Ɵ���胿a݇��!?�zֽ��=J�Ӿ��O���a�)�o������
�� ���P�#�K��P'?ё���ǿG���]ܾ׾?�R ?N]y?c$���"�;�8��� >ה�<�❼M�뾺�����ο�����_?a�>C�ऽ?��>�>͡X>�p>yC���瞾i�<�?|a-?�h�>��r�*�ɿ���g�<���?x�@E?#�5�` ��'�=w��>�R?�SR>3M#�;V�r�ƾ|,�>U��?��?�
>HgW�������Y?�%�=x�L��F��
>vm�=,U�</w��$!L>g��>��=�:�#	��e>i��>��x�
�*��rc�z-2=H�R>�����ս5Մ?+{\��f���/��T��U>��T? +�>b:�=��,?X7H�a}Ͽ�\��*a?�0�?���?&�(?:ۿ��ؚ>��ܾ��M?_D6?���>�d&��t�ޅ�=Z6Ἔ���x���&V�z��=Z��>c�>Ă,������O��I��P��=��{�ƿ>�$����&�<6�Q]��I�����V�����;o��齷�g=�E�=�sQ>��>;W>m�Y>agW?��k?Ӿ>�)>/��Ӊ�aH;d�廀恾�$��6������أ�t��U�߾�R	�9��@��o�ɾ�/J��g=ыN��|��e�0��{j���5���5?]'$>����,I�Hv	�e�¾{c��QS&��B������,�9�n�!G�?��D?�X��*VV����.���.��;U?�Խ�Yپ�����=�~ۼ�z�=�+�>W�=��ʾ��,�U�J� x8?�L/?��׾y穾��>���Ǜ�><�c?��><�6>>�"?*s?hp�<�2����=�x�<���>q)�>��7>�#�����L�>.R\?��������T;>����L����=f�廠���uڽ�?�>}���t�U4����>7&v>3-W?���>>�)���:P����9L?=@�x?y�?BD�>ϋk?�B?=��<�i��d�S�$�9ax=f�W?i?�~>���� оN}���5?�xe?AHN>�7h��꾐�.��)�;?A�n?7?�֟�b}�/�����x6?��v?�r^��p�����ֱV��,�>�Q�>��>��9�Ƅ�>��>?�2#�
I��ѷ���T4��Þ?i�@���?��;<>�6�=f-?Z�>i�O�l�ž�r��.�q= ��>G����gv�x��8,���8?���?���>j���߰����=zؕ�aZ�?��?c|����g<v��(l��f��N{�<�ë=��6J"����z�7�`�ƾ��
�|���7H��ʪ�>�X@8�!*�>�J8�'8⿕RϿ1��Qоx]q���?o�>I�Ƚ������j�!Eu��G�m�H�y���Ş�>�>:H����� ~��n8�>�»v�>�C����>G�,�����~�&��;��>�=�>�C{>h��l���X�?����gXѿ�ߝ�&��p N?�ܣ?~�?ZB*?�%"��ah�īy�ƪ�<��P?Nv?AW?�	�� a�3����j?W_��mU`�Ў4�dHE�}U>�"3?C�>E�-�-�|=>���>�f>�#/�l�Ŀ�ٶ�����C��?މ�?�o����>q��?�s+?�i��7���[����*�!i+��<A??2>���=�!�#0=�PҒ���
?0~0?e{�P.�%(f?�����:���d5���:2|�>�ـ�竜�#ƽ��ν�Hh�׋��W���e7�?A@+��?��Q��g	�S�?h)�>�=��a;վ� �<�y�>3��>k<>DE����=�a���Y����=(��?�v�?<N?���������B>?�|?�)�>_6�?��X>9�?�P=
�E�<>oQ�=��t>��8=��!?a@E?E9�>��>эx�i����$��nO�L�ݾ��H����>���?xSS?c�3>�:9=	��7L�rF�=�̾>�>s�"�H�y=I��Z\L>��Y>��/���<�T�?Kq�}�ؿpe��T0'��3?T��>��?���ԥs�ա��_?�+�>L4��5���"����D��?�J�?~%	?/�׾kvѼί>�#�>���>�yս�Ӟ�lI���|8>�vB?�_��<����o��C�>Y�?�@��?�i��?[��nx��k�����Ҿ�����r
>��?����]�>� �>i�=q�x�WE���?|���>L�? �?U?-�?7�|���L��*�;���>]��?���>[�=e����:>Q-�>"`��u�� �����?Z�@�@�VN?�����޿�����ޏ����a=M�=%S=b5'�,��$9m��:=F�=��=��j>��3>�G0>c��=B��=N��=_���g�.є�m���I�T�̵�y��X���R���v�F@��ɞ��ƾ|��_�C�N��~R�}�ƽ���q��=m�U?gR?"Sp?,  ?z1u�V!>�����=
{$���=���>822?
ML?�*?P�=:���e�S_��������U�>�eJ>�T�>P^�>=#�>���I>�l<>��>�1 >7�)=�,�6<="�N>�v�>X�>s�>��2>��><�������h��f��x��l:�?o<��9�I������ċ�j���&k�=��,?=Y><!��мп� ���2G?d������~%��r>�0?βW?>�;���n�*Q>DQ��oi��L�=�&���q���)�WnM>�?,'>�bZ>�Z(��D�3�V�q��+�>��1?��� ��q�Q^:�]�z&`>lo�>�G0<#��W����1th��=(P8?�a?�7��������$�ee���5>n��=T��;���=��>>�x��<ǽ�g�J��ޥ=�Ă>j�?oPQ>}=��>�˔��?]��0�>�z>��>@*C?�+?;�x;ol��di��E���H>R�>_�c>�9>�jg�k�=y��>j�>Qe���V[��S��s��Cc>�@�z�9HW�#2=��R�]��=Ӓ�=���|=Q��4N=��|?A%ÿ��������7�>�lW?�_[>��YS��3�����g-����?:m@�`�?�!(�c9L�^�<?� �?�9d�J�/>�x�>ye?����Q�%�'?U�'>f6�b�$��7�	��?E��?׮�<�񣿢sw�
�`>մ?�
����>0�DȘ������u���=���>��F?�N��	�K��z>���	?��?������ȿ��v���>Z,�?��?;^m�,��rB?�;1�>���?��W?%Xf>p�ھ��Q�sp�>�??�P?>6�>\���(��?�з?��?�~F>��?��|?e,�>�?I�� �������/��.�0=B�>2J >����N��]��}����i�����ds>�_Z=-`�>M?ƽ�3ƾp��=�1�l,��M�෹>vY>��>+��>1�?�:�>��>�7�;k$��X���NU��2�W?��?�:	��^��4���>I�=�?��V?=��=�r���y�>�HS?��l?�&Y?K�j>8z��ϓ�/l�������G�=�<�=�6�>��?����5��=��7ׄ��>I2�>7���z���˾WIr���>5*?�O�>�M�>�8?: !?Qw�>w5�>l	G���g�88�n>�>`3>�p)?F�{?��?痾�<�䰐�ϵ����R�g�9=r�d?�,/?t(`>(ʜ�k���a�c�-�e�=Y�>\�v?��?:��J??��|?`�S?��n?�>�-&�7���c�Ui=�V#?��	��o@�K�$�γ#��V?cC?L��>j1I�##ʽ���������<?ę\?��#?��lVa���̾ߧ�<�M�L\5� ]��/����!>��>J#��>�=*:>tS�="i���=��B�;��=-�>��=l/���w��O?���=%�۽C �=Mk���$�)T�=ڗ�>����P�[?��'��?��Ì��B��ռZ���?�$�?6�?�E��\^�-�?0��?�T?Ω�>�u���a�4����%��W=8�2��F�=��>�g��
����m\��P�=��<���?�e�>�v,?X�,?>*�c>���wiT�8��"�P3@�k�K93��y�i�4����|j=|ri>�}��_����'�>��1��>��4?�~�>M��>�:c>.-����>���>�>�g�>_a�=!.=ʳ-;Ln+���</xY?,��3�����Xxվ�5R?��X?�>�ٌ�����߶�z�a?Vש?!��?�>��a�����)/?�K�>�s��$�=?S�:>4�<��V�����E�T��|��<�q>/Ͻ�4H�f3������lo?�z?
�h򾾐�<�Ϟ�3}=�q�?�p(?j�'���L��dp�H�S��nV��¼�Hf�Ɨ���%$��r��ԏ�р������>(��Y_=�+?��?�a��r񾶬����f�Zw9��C^>\��>j��>Ď�>��X>/��'-�b]��'�t����L�>!y?I��>f�I?��;?�wP?�bL?���>`p�>�*��xl�>��;��>?�>��9?;�-?D-0?�r?�o+?�c>�f������yؾ�?��?�E?B?S�?��bCýb-����f��y��k����=�-�<h�׽�u��pT=|�S>��?��	��D8����c�j>I�5?���>���>PA���V{��T*=-��>�
?#��>>���(Vq�-h	����>�ȁ?v��l =a�%>��=m��}��a�=�.��~�=D�%?7��%<��=t�=��}�뺴�s;�<�N�<C�>�?u�>=��>�񅾯 ��F�"��=äT> �U>�)>9�پ5e���U���g��	x>D+�?��?�xi=]4�=v��=iȞ�Φ��������x��<�'?�u"?��S?6h�?� >?u#?��><#��<��;k��������?!,?芑>n��ݳʾ���3��?c[?r<a�����;)���¾��Խ��>�[/�./~����vD��
����������?࿝?oA��6��x�׿��\��#�C?�!�>Y�>Z�>X�)�d�g��%��0;>���>�R?"�>*�O?={?;�[?KnT>��8�w0��"ә��2�Y�!>W@?^��??�?�y?�s�>��>��)���aQ������₾� W=BZ>��>�&�>��>���==Ƚ`����>�&`�=��b>א�>�>� �>W�w>M�<k�J?��?=_;����0��W� �&+ؾ�z?!Q�?�5>�m=��C�݈g���)��l5?�ִ?[��?�Ζ>9S1����=�ǭ��[�yÙ��:�<�
�>֑>r9�>��=>m��>;�v>PZn����*�E��`o�z�?D�V?z_��^�����L��T����RxY����;8:�V:�=���V>������������6��ڴ�=�D��^�'*������vi?�M7=���=:
>!]�=��7�t����,����<�R<>ǽ����r="x�ݬ6<��ҽ�͗=�;=�Ҽ�ƽ�����jp?<�?�l?�:6?
3�>��4>?����?5	��a?R,�>d�> �������p�w��x��5������Q��p�=���̶,>��&>f�k��-=1��=%8�=
���� 5����=U$e=�]|=�_H=���=(KG>�a�=�{w?S�������X�S�׼��1?��>�''=�P����A?G��=����&��xB���~?9�?QZ�?
�?3�0���>����>�{c�=X5�%O�>�}�8l�9��>�B��)��g��8=�I��?]8@pG?zy���LϿ���=e78>|�>�#R�ֻ2��]��og�%�S���"?ƨ9�wCƾ�Q�>�f�=��ݾ�ž��'=ο4>�	y=����[�^b�=eu��<:=�}=v��>�j=>���=闰����==t?=���=a�N>ѭ�$�:���;�@�0=t*�=Wa>;$>��>D�?g"?�zW?���>L��	�辖���:T�>��t����>ó<i2>�1�>�K?\�V?��J?�͍>J0�=w��>dܒ>��-���c���վ�����U3����?��?iܭ>k�X<C�-��&��<�#���J4?�'?-��>� �>�p��,߿���,)��V罏 ̻��;9����=������	�����6R�=&G�>R۾>���>I�S>neA>�m3>$�>"E$>�=<hi��A_�Q���꣗<��=/m+��g7=���!�{��M���v#�֪�l�<*�=<H��<�<��=so�>̪>k��>">}У��	�=�˱�u&R��_�=��Ѿ��A���X��Uy�	�#���G���
>f�>��f���S�?~�s>��Y>�G�?�"q?��>F�������َ���+0�{�T����=��e<�?���D���m�"�E��L�����>�>2�>r�l>R,�f ?��w=���b5���>���E��,�/8q�0>��/����i�֪̺ �D?F��|��=�!~?�I?x�?Z��>| ��.�ؾ�-0>�E��5�=]��'q������?Y
'?ĉ�>�쾔�D�D.Ӿ�!�{��>������:��������X��Aھ��>�Ƣ��N���G5���t��~��u�V��N���|�>�?��?�7��y����=�#�����<-�>��S?Y��>��3?��>>���t��sA��}ߖ=�Mq?�&�?���?�@>]�=�o��>I�	?IŖ?��?.�r?�E����>�t|�s1>���� �=�>y{�=}��=�i	?O�
?|3?����1'�x���]��r
a��s=�y�=$Ė>�@�>�v>���=IDz=�١=ý_>ϝ>w>�>��h>���>Oш>�屾eO��[4?�>���>~�I?��w>LH��uM��~���O=��@�LQ��mf�;�h�S]��K�=��>���>9&���E�?3c�=�8
����>�J���=�ܙ>V��>*<s=���>��=�]>�Ӯ>���>�>��u>s�>����=����-�Z�N�R�t�LX@� >pѸ�I�2����� ��݅�ph��9��[�_�)���f��e =�?��D��V����+���!?�ђ>`��>J����E��5e>���>?i>���4��M����ʾ���?�� @��B>���><hR?��?�q/��ƙ��#i���f����sd�\�<�)��*wf�χ �d�=tUk?�s?	0?��>�>4�?�9�j{��ܸ�>�/`�L'�����s]l>���.Q
���	�!X־�cv�;��>#��?��r?K�>�_�Ge��IO>�T?�bK?n�w?q�5? (?�X���'?�w�=�?�?E8?�v?��>%�>������:�<R���]�����r��s�Si�<vM=Aϫ��3�����<���Dfa�v��w�)=�@�;+��<i_+=�C=�~�=�>{]?G��>a��>۰4?lJ�%:�����$�1?sZ=Ϧ}�����ު�_���!>'�l?�ڬ? \W?r3[>K@��E��j#>i��>? >H	\>v��>rWݽ��J��j�=�7	>��>�ϝ=ުq�2����D	�L��'�=*_>q�>O�~>��\LT>4��K�k�O�F>K���C���w�u��;T�b�'��d����>�	@?Q�?A(}=�%����|�M�l�^/=?[5?ǦJ?R�?�w@=�/پȡ3�� N��Oн�w�>vl��)������E9���%��@|>zo�|࠾]Ob>߽�s޾n�#J�]�羍dM=]|��_V=l���վE7�	��=�#
>����� �e��[ժ��0J?�j=�y��0[U��n����>���>^ٮ>X�:���v���@�.���F3�=���>Q�:>?;������~G�	6�n=�>�UE?v@_?�a�?�傾!s��C�8���.ɢ�C5Ҽ�?r��>�]?��B>^@�=r���$����d���F�)�>H8�> #���G��N��mw��d%��y�>&?I�>ة?��R?8�
?(�`?�C*?�??��>����<D��vr?oل?
�<0���ս5;��b��|�>4?rH���Ԋ>P �>�\?��4?��e?o?�:�=�\���{�kY�>>^|>E�Z��谿ìh>�K?DZ�>��I?:3�?�[r>��2�Q���D��vJ>�T)>��?�$?��
?=v�>0��>����|�=J��>nc?�0�?��o?Ԁ�=��?D92>���>$��={��>���>?XO?��s?��J?&��>N��<�7���9��B@s���O����;rzH<o�y=L��16t��H����<�;�n���L����@�D�	��L��;tW�>�Y>G[�gȲ;�龒�;�-��=�X��-7ƾp�þ�F��6u>g1�>�y�>��>I�㽯��>��
?�$�>��B�lj?�x�>�f?�hd=��e�b�˾�=���>��<?-/�hZ��_ȣ��Ҋ�`p�="�L?ڰQ?�4�=c����<n?��6?4��g�8��=���q����s?ZR/?�(Ӿ�}�>8xs?��h?Y:�>۳��b
�������F�X<���N�=��>��\5;��	7>�JU?u&�>�4V>n89>5������ԩ�J�>u�?.U�?Ր?��=�P���s�~I��`.��W8^?U��>�e���"?�T�5�Ͼ����ZҎ���;��mM��	8���b����#�t���b�ս�=��?i�r?5Xq?l�_?�� ���c�<^��	��aV�� �M�4�E���D��PC��^n��
��������� H=�q���9��o�?�&?�S����>F~���n�Bᾄ6A>�+��V�=�<�ʒ�Y
= °=�t;� \ٽ-���]�#?!��>V��>�4?0#U�n�4�cJ/�B:��O��g�>v�>.Ps>�i�> Q�<]�˽N��	r�����D���5v>Zyc?��K?N�n?�t�(*1�D�����!�r�/�+`����B>�j>q��>��W����<9&��Y>���r�>���x��i�	���~=m�2?z(�>���>"N�??c{	��j��Nhx�φ1�c��<-�>i?�?�>2�>zн�� �ٴ�>��l?��>��>����7W!���{�R�ʽ��>V�>��>\�o>��,�3 \��h��Ձ���9�s]�=�h?ώ���`�a�>�R?�M�:i7H<qs�>��v���!�����'��>O|?��=g�;>�|žE)�y�{�v6���(?�?�y����)���>)q"?&@�>t��>w�?ӌ�>�P���ﾼ��?�b?� N?�!A?J��>�=š��2���h(�Hw=/C�>2�Q> g`=�N�=�'�B�P���$��FG=j�=$� �?˽�<d� ��ц<(֞<Oj'>.mۿCK���پO	����A
�!戾���a����'`�����M]x�����'��V��9c�Ǣ��6�l�K��?=:�?N����+����������[���Ư�>��q��������:'����R���ib!���O�|$i���e�Q�'?�����ǿ򰡿�:ܾ4! ?�A ?:�y?��4�"���8�� >EC�<1-����뾪����οJ�����^?���>��/��k��>᥂>��X>�Hq>����螾�1�<��?4�-?��>��r�0�ɿb����¤<���?/�@��J?!l��/پA��)�6?�6?E��>VSY��M0��qؾ�k=o�?bL�?}��>#�q��K���Hy?I+e>�؉�e�<��I>�g>wMr<I�,��N�>�5�>�:��>�
	��}�>
�?�д����9����>x9C>�����Ч��?�S[��@f�l�.�a��bf> nS?F;�>�=B�*?XVG��HϿz�\�	q`?GK�?9��?��(?O¾Y&�>�(ܾMUL?7�6?H��>y�%�+�u��j�=v1�� l���c(U�j�=���>C�>�..��i��dL�������=��<+ƿ)�$����{�<CT�zm���⽤ġ��E��S����o�����!e=�f�=.^P>�M�>�eW>�zZ>ZW?Mj?��>g>� �t�����̾������������"�������S��ݾ}���S��5�}#ʾ	(=����=�5R�3����� �w�b�t�F���.?w�$>��ʾH�M�$D-<1sʾ��������祽�(̾��1��n��Ɵ?��A?������V���si�F���ĬW?�B���D䬾2w�=�ձ�F�=��>���=����3�hyS�[8?�6?pݳ��lȾ,>��L�s>K/@?C�?�v>3Q�>��?J������$�=��>�|�>z`�=v�=��ξ$�޻.�)?(^?LNf�n鵾>y�>.�ʾ	ľQ=>G>������Zg>�QJ��3��W�=���=��=K�^?4F�>9%�?}"�k×�D%\��3>��?Ԍ?���>�!�?�A?Lx�=V��P1]���;���`�X$M?�i?�/>@=��9㾪�Ӿ�/?�π?�v�>3�[���l�����^?�s?S�,?�>.=Lu�H�����#?��v?�r^�Ys�������V�T=�>�[�>4��>��9�Yk�>��>?�#��G��庿�DY4��?��@���?��;<�#����==;?�\�>'�O��>ƾ�z�����+�q=b"�>̌���ev����DS,��8?���?1��>����������=87����?d��?�I����?<�����k�z�:�!<%��=m6�_ ��l�+�4�����A	����#�l��ɇ>hb@�4����>s�)�E��UϿ�t��о�@x���?��>�)��G'��ثe�[Ss�j�G�` J��S��9��>^>�d��ԓ��{��Q;������W�>���ԉ>"jU�uQ��p���<�~�>���>��>5����Ǽ���?����
EοZp��t�sLY?�?R�?�?�b+<�w�*@}�e�'�~'G?y-t?��Z?
���r\��!@�%�j?�_��xU`���4�uHE��U>�"3?�B�>S�-�j�|=�>���>g>�#/�y�Ŀ�ٶ�?���Y��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�B0=�UҒ���
?V~0?{�e.���O?�|C��[a�����_�=.{�>a�۾	ƅ�j�.�\Ŗ��pI��R���E��S�?j��?�ְ?��r� 2��7?I��>[څ�1��
	���?�˯>������r���>d���;�+�p�=#��?���?��&?����,��HȆ=o|?f��>Hh�?�M>'�?a���m������=
�x>*�v=Q��=�H?}6?�>�.�<��q����[�<�l�X�H����R�>�QZ?��v?>�&>l�	�[����1!�T����x��ů�=��-�N�=��C��B>jL,><����f���Ѿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji����>M�����������l�3d>�A#?S��v��>ⰸ>S
=^�t�����P^r��i�>�5�?�1�?Be�>+��?�j���^���?�S�>�y?/��>���=���$�>�J�>���U�����˾�Gz?,@9	@��N?@Z����ٿ����ݰ�*� �ha=o���s��<;T2�eH�>��=�ن���H�?�<�K5>��->�.>	�$>u��>�
>�����_��E��u���l�C��s)��w#��� ��`���1����O;�]޾�R���L�EܽE[F�Ҭ������=��U?� R?�+p?�� ?2x�,�>F�����=Q#��ޅ="3�>�V2?��L?Պ*?A��=＝���d��\���B��I�����>�~I>&��>�Q�>��>}F�8[�I>�?>l��>�� >��'=�l캫�=R�N>�H�>���>Zm�>N�<>N�>̴�8'��(�h�Qv�g1˽�
�?����J������v���I�=�X.?N�>����?п0���sH?ǔ��!�N�+��C>*�0?!W?Rz>t��
R��>�����j�C4>*  �8�k��n)��vP>mn?�ӌ>�@y>u7���=��F�˚��}>�D?����h �
=d���8�&�־��">ɋ�>a��<e#�������x��Ny����=�9?v��>;�%�ڐܾTx��X����=�R�>�+o�E
�=��>ʾ���e	�tU�Y��= �=;J�>hB?p�8>)��=&Ӣ>|㟾z1X����>��H>��(>4oE?z�?ä��x�̽�S���-8���n>"��>��i>���=?v]����=���>q0�>�5���G`�xv��O�2'J>-ۓ�EO�a4d��؅=���lK�=j=@���� I=�ls?JQ���㍿!��9�>��i?�K�>Rt�=L��H�,����^��b�?�@fH�?�4/��]\��&?El?[x�!
�1��>���>���z=��%�?8�XJ_����t�#��?^Z�?
a� ���DY��
7�>��?
�o��>yV�fQ�������u��$=���>UVH?�����#Q��N=��
?�?6�򾓦��Mɿ�v����>���?d�?X�m��6��@��/�>*��?�tY?�^i>�3۾��[���>Ͳ@?2R?W�>�Pu'���?���?���?I>���?��s?l�>�&x��Z/��6��Ė��cc=�[;bd�>�U>����}fF�ד��g��ںj�@����a>��$=��>�H�)5���;�=��G����f����>H-q>m�I>wV�>� ?�a�>W��>hn=zm������^����U?�Ճ?!����m�nQ\��%>���_�&?��M?Tȼa^�����>�$G?n�W?f�G?%��>�8$��~���#���c����==Y>�@�>s�>l*v�W�=�߾f������>n�6>0�����R��
��1�>�)/?[=�>�8>�N&?�D ?��\>���>>"F�������#���>ۣ�>=�?���?��
?�d����A�Υ��΅����B��:�>3qq?�k#?��z>Qݔ��g�� 5B=ύ�<�/��Jg�?�hf?�z_�]%?��?��N?ς??�e0>�	��{��/��D��>�?��>�IP�T��]�=�*?q��=� >�'�%u���Pt��S��t��[�N?��?Υ/?\5�$T��9;>�=+I��M�����<��"�=>Bs>Ȝ~=�Mi>hZ>L��=\=!���$i�I�\=��>o�L>������[�B#,?��B��h����=��r��oD�ڢ>3�K>A��2�^?�>���{�*���r����T���?'��?t]�?/v��O�h���<?0�?�?���>?���L6޾���)�v���w�ד��>4��>Ky�o>�W����r�����@�ƽ�A��n? �>�u?�v�>�U>0��>����'�������ZQ���u�9�K�-�����sG�Km�:̡��a�����Ol�>�b,��d�>���>��?>_6s>!c�>��y���>9nQ>�?>7��>��>1� >{��<�tp��ۼ��[?ֈ�� ��:������t?&�m?Rl�>%���n��ѕԾ�o?��?i��? >�S��<��@�>[O�=�s����,?��<a}���)���Q۾	�����0x=�M�>���&8���h�ǻE�C�?*.?o�<���/�C>���sk=5�?x�(?��)��R�zPo��W�T�R����[Ah��u����$��lp�z�P��@��|r(���-=&�*?l�?�=�'�����(�j�n?��~f>@v�>��>���>9jI>_�	���1�d�]���&�=��h��>�{?���>;�I?= <?�tP?�hL?��>�_�>�6��~h�>7��;]��>_ �>0�9?~�-?�60?�x?�v+?~Ec>Mw�������ؾ?�?AJ?�?�?�څ��ný�r��N�f��y�������=d��<[�׽�Qu�N�T=�T>�E?�?�d�8�H�����k>_�7?���>[��>X現�s����<؋�>�
?6k�>�[��M�q��m����>.��?y}�r}=�:)>˻�=��uܐ�L3�=
����?�=k���DZ:��, <Q�=���=(�����!:�s�:�Za;�?�<���>�E?b0�>�C
?j�پ���8w��>��tN]>c�>24=�����膿ߤ��JW��4>�%�?��?�㽼��o>cQ�=c��+�>"�k��`��=�]?�J\?��?�n�?x?sd<?jq�=�����R�l��ݰ���%?� ,?P��>H��t�ʾ�樿��3���?m]?W5a��a��6)�~�¾kս�y>�P/�U~�s����D�����7��Ix�����?���?5�A���6��]��Ø��m��ǦC?���>Xb�>c��>��)�5�g�Y/��[;>��>y�Q?eP�>�-R?8`q?`�U?�nr> �9�˱�𬗿�A �^C�=!;?��w?���?�p|?C�>� >g5�l�޾1o־�������Ȍ����<�;`>�g�>��>��>�B�=$񕽯Uƽl"J�b�=
�i>v��>=u�>Q��>��k>b)=W�G?���>i(���n����]��W�N�(�t?xȏ?�E(?ir=�L�)�E������x�>��?�g�?��&?l�L�Dl�=q"�V����k�1�>l��>�K�>��=].=�!>X�>HI�>���/x���8��>��?>�C?�^�=M`пV�_�پy�{!w�ShC��0*��G�����L=�=���>�Y���\�K�������wԾRo��%�Ǿ��I��Nƽ��?)1���=��3>s��� NF��r?>�)�i�r��`<� ���%�f���|vл��<����oG��c =�#�=��¾�?!�?*ǂ?�?�q�>�H+>^6�=��q>:�<9F�?)}�>��<
��t�y�%�e���þ���SO��Ma�܌>��G�>x;��r#�>�Ύ>ډ�=?/�;��>���<�o:>�X=d,�=�=���=�Ǒ=��=>NF>m�)> mm?݄�����4Ca���O�J�0?�3�>�7�=j���b�6?G�=h���������H`q?�h�? 0�?1?]mS����>ӊ��뽔�=Ron<
W�>�f5��16����>��=������QB��w��?�@�f7?߭��h���wR>� 1>̲
>�R�320�|�]��L\��Z���?+�:�u�;K}>7"�=�ݾmȾ'� =}�/>/ϋ=H�n"Z�-��=cx��0=Q�=|Ɗ>w�B>�l�=����=�r9=>�=� F>`4��C�W�L��=3��=JrX>�8$>�?�>��?�\0?�kd?�o�>j�o���ξ[Qľ^��>��=�ά>QE}=�<>r�>��7?�QD?	L?>�F�=���>��>��,��"l��2�J����Q�<���?���?y�>�Q�<��?��m��T>���ý��?F1?��?N�>J�+�Ͽ5H%�$�5��N潼���ڟ�X|*����=0�p=M��U����x=寐><t�>�q�>��s>^�O>��Y>��>A6�=�!�=���=���<�&M���M;��=�.��E=A�׽���<e�R�V*�q��<��<�.!;d���E �K��="��>C�>���>��[=������ >7U���H�w+�=^ᶾ��<��\��|�y)��{7��r>*X�>�<���-���W?#�8>0V>z��?V�o?xY>x��O�ϾQ���|W���w�}�=
��=��L�d�:��:\��!I�XWҾ��>���>�	�>��l>',��"?��w="�b5�}�>�}�����_1�A9q�?��N���1i�(�Ӻ�D?+F��^��=�!~?R�I?�ߏ?*��>�����ؾ�90>9I��M�=�
��%q��x����?�'?��>�쾍�D��d޾��u�>A�w��L�	���a-��Ÿ�M�˾x7�>]ª�H�ƾ+.5�T|�������*�4yb���>�M?��?,)���C�r��㾸��Z��>�f?ۺ�>�W�>�n�><l���[쾪P���^�=�U~?��?���?�o�=���=�ڴ�S(�>�$	?7��?㵑?vs?��?��n�>��;�� >�	���>�=d�>Μ=�2�=n?��
?7�
?�[����	������Q^�B��<��=c��>q�>�r>n��=��g=�R�=\> Ӟ>��>��d>u�>�G�>E��I���)?%>��:>&Y%?
>��*�L�F�d�ʦν�0�ݓN�����i"��0���s<�c>��=iQ�>�N˿���?�8>�/��:?T��Z4S=�z�=��`>�z;��>9�>���>d�>�2�>P�=�%>���>�HӾ�z>����c!��,C�R�ʼѾ�zz>=����&�r��2x��(DI��n���g��
j�".���;=�MϽ<H�?3�����k�6�)�o���Γ?�\�>6?ی����{�>���>�Ǎ>J������Ǎ��f�2�?���?�Z>��>%�k?�?��l�A�&��`�nvn���S��[�LG������m��h�]��~�m?v�i?*~8?��=�?�>��?�2��iV��/�>�@>�� G���x��0r>dNܾ7�1�vV�B�l�ZC���;�>\
c?�7a?�7�>4���dR�� tN>zC?�7?L&x?n�8?��7?�`
�1�(?B>>Ɉ?aU?�1?SM'?W9?��">Ȅ�=��`����<�,y�֬���SڽX�轷z#���?=%.=��	�yF��\�<n��<]��u���z���������<"qL=�'�=�=ID�>�HT?�$�>$��>M?.<�v�&���޾g?^�=JȾ���կ�X���5�=O�J?�©?L�e?�1=>y[�4�(���=�q�>v<>2�k>���>�t*�A�̽O��<?_�=��=|*�<�w
�+����!�|� ��<<��=|��>a�>�Ã<��> ]@��龚�>	�^����_�6�� B�uc߾sV@>@qX?�Rd?��C><K&���H����>�~?��X?aE)?�0�X}3�a�;�5pe����>.���w�>��:m���Ű���@��oa=�s�>��D꠾QBb>���~t޾��n�J���羬EM=���ɓV=\�9�վ7/�	��=I
>����*� �+��	Ӫ��1J?1�j=x��lU��q��g�>��>Qۮ>x�:���v���@����Y%�=a��>��:>�u��� �9~G��1�x
�>�3E?��_?�|�?X��� s���B�
����٢��ض�4�?�^�>�?�@>lH�=�ӱ����z�d���F��b�>�s�>���H�屟����$w$��Ί>�W?Nu>� ?��R?'�
?�`?��)?�?"��>3:���Q��f�%?�l�?#�~=� ٽ3�M�=69�x�G���>��(?(�H���>�9?�?��$?��R?Ŭ?Ӽ>
� ��$?�$P�>{�>8�W��Z���f>�lJ?1U�>uuY?X��?�>>�j5�����,r�����=�>�P2?�"?�?�C�>x��>:���u�=���>�c?�0�?�o?��=C�?�:2>k��>}��=���>Z��>�?GXO?.�s?��J?��>9��<Z7���8��sDs�M�O�Ă;�tH<'�y=W���2t�K�[��<� �;�g��bI�����z�D�������;s޸>z�K>�ڒ�|�N>���.�e��3>I���3tǾܕ��$��#��=x��>.i?�4�>�f&�n�s=C��>N��>�7���n?sM�>+�?���=5_h�!9̾A�)��>cFL?~5>ӈ��ޮ��ʒ�E�=}vY?�@?�z��'�o?�C?����:�,���ݽO����aV?��?�]��2�>�Ѐ?o�t?D�?ߣ^���q�{w���-b�������=��]>5$"��XX�쾐>y�T?�k?�k>=�C>�p��r�������?��?��?���?VS->T_�?��A������/�^?�	�>á��8T"?C��hоZ�������������h����,�������$��P��p�Խز�=:7?ZMr?.�q?�`?4 �1�c���]��!����V�����u���D�w-D��C���m�p�|_������E�E=A�v��+�0d�?h"@?����o�>0�����є�7��>�iþZ!�B�<yW��9z:�<DzS�6 ��Ц�Y�	?�>XZ�>(KC?�>��G�Ч(��?F�������>'�i>��>}��>�܀<{,��#L�yQھ�韾���,v>�xc?J�K?\�n?{��)1����T�!���/�{g����B>Es>ʻ�>"�W����8&�X>���r���,z��=�	���~=��2?*�>R��>�K�?�?�y	��t��mdx�͇1���<.�>�i?w7�>a߆>н� �|��>+@l?��>�͢>8��w:!���{��̽B}�>��>ڥ�>%�o>j�-�#�\�-0���C����8����=��g?K�����_�c[�>�WR?0�;X�<���>�݂���!��𾄢)���>c?{��=V�:>rƾ�^���{��䉾�:-?tP?�n��B-��ex>.#!?�.�> �>�9�?V��>W����<��?j8^?S�K?�4:?fq�>�<Mcʽ-�ҽ�	���E=E'x>�5_>�@=0��=Y���V|�dx��Q=�!�=��� S׽�9�<߼�3�<��O=�D>��ۿ�XK���پ>9����~�5�������^���"���N���Ә�R�w�&��4��WV�>d�V�����k�'(�?���?�;��~����՚������8��K��>N�q�n�p��ޫ����eH��E �i��J!�	P��i���d�n�'??�����ǿ���#>ܾ� ?A ?��y?3���"�ƒ8��� >� �<�✼��������οc���U�^?6��>O
��-��a��>�>�X>�Cq>h	���瞾���<�?Q�-?m��>)�r�X�ɿ�����<���?��@8~A?W�(����� V=_��>)�	?=�?>ZG1��G���
K�>E<�?' �?v�M=��W�X
��ze?�<�F�K�޻z<�=S�=I0=4��N�J>�M�>���XA��=ܽ�4>�߅>Q�"���w�^�K��<X�]>i�սE��5Մ?-{\��f���/��T��U>��T?�*�>U:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?$�(?8ۿ��ؚ>��ܾ��M?_D6?���>�d&��t���=q6�ʉ��{���&V�}��=^��>i�>��,�����O��I��Z��=���ƿ��$�������<~g��oX��'��@����S����� wn��X�-�i=M�=T�P>z��>{�V>�Z>�UW?(�k?��>�>��W����;�L��Z���=�����Y�����O!�}߾xj	������qDɾ�=��.�=E3R�����û ���b���F���.?yT$>
�ʾ��M���*<�oʾu̪��J���_��N̾�1�^n��ʟ?j�A?J�����V�F��"h�����9�W?&�����מּ���=����N�=)�>���=6��m"3��uS�G�J?C?'"�������=R�;���*>��K?uV�>��l>��>��?u9���p�8�u>�:9��>��7>��B=�ɾ܆��!?0�F?�VQ�q�оb9�>h��
{��0u;> L=P�S�6����Z=�@5�F^�/x=*�����>�(W?���>��)�o�%a�����c^==4�x?��?C.�>�{k?��B?�Τ<�f��U�S���*gw=�W?9)i?H�>�����о
����5?��e?��N>�bh���龊�.��T�J$?5�n?E^?e����v}���k��o6?k�v?�M^�PZ��M	�PHV����>���>O�>F�9��;�>�>?��#��Q��󴿿-;4����?�@���?�E6<������=�^?��>�vP���ž�l���ѵ���o=�2�>����&v���3A,��O8?���?�>抂�ў����=�������?}5�?���A�Y<� ���k�n% ���<xU�=s�y�%�W���7���ƾ̊
��V�������3�>l(@�C���>_7��[Ͽ����о�xo��X?4��>�sǽA��pyj�wZu�ۮG��H�:t��ib�>>:���U:���V���1���z=��>��V<��>:���B��߱v��n�<��>k�>�<*>��L�OM���B�?���ۿ�.��?�]�?�a�?�$�??�??�kZ�v�;�����!>��j?Q�p?=?�(��b�:�i�|��j?G`��nU`���4��HE��U>#3?�B�>Q�-��|=<>���>j>#/�D�Ŀ|ٶ�7���R��?�?�o꾆��>k��??s+?�i��7���[���*�c�+��<A?�2>)���6�!�0=�ZҒ���
?W~0?�{�j.��~`?ч��D���#��mc=(�?F�L�C�[���=Ѧ�pUT�����V���?S�@��?y�V���K�?���>^Ƙ�󫾿�>o�>6|�>�~c>^'���>�����X����=���?�@��	?�����R����>�!�?�2�>�{? B�>�_?yN����ɾ��>$�(>�5>�J��%?n�P?��>��,>e}��<"�Ӡ`�v���PO�e.�>W?T�c?�Z>[�;�P�����_���V ���<�@C���=�	�;4�>ˋ�=�R������=��{G?6 "��!пc꘿�m�J
?���>AB?��bX�n����e?��K>E��~���m8������խ?���?=,?���9¨����=v��>8&�>
�#���1�y�QzK>�{F?[>�8���w�6�>�޿?Ĝ@�,�?��l��i�>���-F�����i�߾=;����=�*?���.u�>��>>-[���Ğ�������>���?P��?g�?#@�?뀿n�N���=�	�>gЀ?o��>���{	����=Y?��7��N���-�ɯw?�1@<7@іT?����U޿�ꌿ�絾>�����>2��]&]>������6֩�p�Ƚ�(�=$>���>�.=Z~6>	y>��(>Sӷ=�Nz�A��aj��ډ���Mb�_mC��ɾ�{N��'����W�=�LG��Z����#� ye�!����t�.\N�y_����=D�V?��S?�8s?��>�$���.$>u���=ڎ4�Ѫ=�҈>B.1?>_K?C&?�#=:��X_f��灿jx�������>B4F>��>y��>.x�>q�#� B>,�/>LT�>���=��E=~P�
�=��C>�,�>&�>@�>,f<>,�>ʹ�2/��١h���v�ܚ˽� �?�f����J��-��y*�����t��=Ib.?=g>��� >п����w.H?H���U)�c�+�� >*�0?�]W?9�>���/�T��E>�����j�{c>�	 ��jl��)��Q>Cc?kk>Ziu>��3�+�8���P�����<n>U�6?|h����5�u�s��GG��tܾ��N>�v�>�i�L?�6�����~���i��L�=�:?X�?#
���V��L�w��㝾b�M>2*^>'h=�C�=��J>��k���ɽ-G�/*7=�_�=�+b>z�?3fV>{n�=�s�>f���'�����>h1z>rg>M�S?�v)?E�f<�$��h�o���<��CH>?��>0*4>R�>�뉾���=�?��>A�G��O��a�Ƚ�x��J�>�˿�˟X��e8<_T0=�Y/��U=5��=�4#�H�x�:L]y?9콿4���D��X9b�y8l?��?�\�=�����%������g����?��@;�?p����X��G?��?S?��Ѣ_>�$�>�>���ۜ�P�?�9����Ӿ6������{�?O��?��e�sv��D]n�0�9>6�?ㆬ���>ڍ#�py���)q�	MC�T��>�QE?U�G-y�8�L�-�?�d�>��+v��^Tǿ��w�e�>h�?��?el��A����;����>���?��Q?�n>��Ծ�6�̍�>3c;?klE?J��>;��S�#�yd?�A�?�@�?U�A>\p�?�z?�B�>ɽ[��<0��񲿨݋�/=�3E=���>^>�Wþ��I�P���w���f�����X>�N"=ط>{�ν㭷��J�=����8��=��2�>Rhp>��J>�>Ѷ�>T��>���>��<�̔�I/��y���,Te?��?u����k�ў���G>P.� C+?��H?��=�gb�U��>�$D?�`~?X�c?Q�:>��޾����;��m���#>�(A>�N�>h	?R:{������뗾斻�0V�>n��>GU�;|Z��齝�~齼F�c>�y&?���>9k�>[? �?��>�k�>�+J�V)���v9����>�ɶ>E%?�l?7<?�����B1����.����T����=�?s?s"4?r�d>�?���@�������-=#��=�ԍ?5>x?�c����(?���?�*M?MZ?<�I>�'����y>��fr>�&?Nd���A�IS%��1�y?a�?��>=���*۽E����q�뾍u?��\?� ?����d���ؾ�G�<��<�<2�=t;U�:<^}>���=:d�lG�= �'>�(�=8�p�
<@�M�9<�d�=���>!�=��C�8���̟?�lg;�0��ͻ=��R�`\#�u��=���>^����[?��<��{g�Y쫿�Ԡ���{�0��?���?J��?������Y��,?'��?s�[?+��>�ƌ�*ړ�TO2�쾛>
J[�l�>�X�>�b�W�Ts��2��Ć��7����u��j�?��>�?�8?�r>�l�>���V�������ɴZ�l7��11��/���"���ϾY�=�!>>��þ�[����>�@����>��?���=��>���>�K����>78#>��>�p>�=w@�=0ջI<�%�A�b?�� � '��%ʾ���y�k?�q�?�/�>���=~z�%��ZQ@?yϣ?�>�?���>�HZ���KL�>;�G>b~��mf9?)�=�V���@�=Z���1Z���ى�V�A�p��>�Ƽ���_���l��F?Z\?�G)>g����e��h��?��=��?C3B?�Y�]�E�j���X��Ea��P> 闾�K��E�)���y�h����*��Yo�>�"�2��<,E1?�+y?��S�pG۾�`�]�����>y��>4�,>�T?��4>,��� ��0X����/���!�> hz?��>͉I?@<??vP?�aL?Y��>Ck�>�*��\k�>}��;��>	�>J�9?x�-?�00?w?Is+?fc>����M��|ؾ'?C�?xG?;?e�?䅾�Uýᤙ�B�f�ӣy�q��+�=	��<=�׽8�u���T=3�S>�^?���L�8�������j>wx7?7��>��>������B�<�>�
?gE�>G����{r�QW��@�>��?�F�u�=�)>R�=g)�����<^�=��¼Π�=�I����;��<��=��=��|��g��&�:��;UG�<F�>��?Ŋ�>���>���U� ��g����=?�Z>'$P>�>�۾�݊��<���sf���{>wN�?���?�oV=5��=��=˃��5��6�	��G���a	=��?� ?΍T?Y�?o1>?g5"?v�>ZD�0̒�aY���r���?f!,?��>���8�ʾw񨿅�3���?q[?�<a���2;)�&�¾�Խ��>x[/��.~�(���D�3������~����?���?�A�e�6�7x�还��\���C? �>Y�>��>#�)�7�g�X%�w/;>ȉ�>-R?"#�>k�O?�<{?�[?�gT>I�8�:1���ә��J3��!> @?䱁?��?�y?t�>��>��)�ྻT��0���������W=q	Z>���>"(�>��>���==ȽfY����>�Xa�=��b>��>��>�>��w>L�<��.?#?Y۾�!�8�>����N���?�y�?%�^>�|���E�0SQ�H�+�d\/?i<�?B��?�u�>�L�gM�=	�b�y)X�����ӧ�>�ӛ>yH�>�v�>���=���>pz�>W֞>քf�Q�׾��3���i��?80J?W��%�ӿO�k�r���;B}]��=�@�˽_hv�U>���@>/�оұ㼫ӕ��P��MO�����-�ݾ�Я�M%��/?�_�=o>�=�ͳ�6{߽���f������<+�}�2>ZD5�@B=�Ž5�b���"�Q�#��Ȼ:�K�#>����)@y?�<I?�k?�7?m�>���<Bն�+D�>n�����j?2h�>=�,>���j����u��ud�YEﾃ�!�����᝾m��;y�ؼ͆�>�x>񝕼n�=��6>��=�Q@=<����X�<.��v��=�	>LJ�=z�=�{E>�wn?�T���"��2M]�j�k�{u=?�5n>��b=��;�:?X�3>����D���l���l?,��?E��?|Q#?�E8�{t�>ZѾ;y��dF>q�-<`��>:�:�EX�]L�>I�N=ƫ�YѬ�(�G=���?��@��P?���O�׿4
�=�A>��>j)R���2��=Z�.�a��)V��#?
�9��YȾCv�>A��=�޾��þ�CO=
�0>P9z=����O[�~�=t�i�`�G=v9d=�A�>��9>rĲ=޷��Ϡ=��_=Rq�=~�J>�]���5Q��cF��93=Qr�=pZd>\�*>�6�>�?"�/?Sc?�5�>��o�q_Ѿ�t��z��>*��=+�>��y=4�@>Z�> �8?`�E?9L?�7�>?��=�f�>l��>��,���l�P�⾭צ�g��<P��?��?)��>:6<F>��S�ݳ=�N5ý�X?*1?I�?G-�>
V���X&��.�,���k��i8+=#ir�p�U�i���|�d��C
�=q�>���>��>jGy>
�9>��N>��>ʥ>�'�<xX�=������<n����=�Б����<��ż^b��}(��+����ה�;h�;��\<�#�;��=���>� >nI�>��=)޶��F1>"h���K�r��=ǳ��QC��Ub���z�"+��<��1>^Ƅ>����ǐ�tB?	�X>wAA>��?��l?��>�(���¾�~����>�c��H�=�l�=>�d���<�y^`�[xD��Ⱦ���>ݎ>z?�>*m>9 ,��?��Lw=/�o5�gL�>���6��"P��Aq�W7��6쟿��h�g"Ⱥ��D?�A�����=5*~?)�I?�܏?�Y�>�<��)�ؾ��/>���=�=���j�p�vy��M�?_�&?�]�>��$�D�P־+���>�h�5�K����Β)�l�=���Ǿ﫻>nί������2���o����D��H��Pi�>!^Z?�q�?Ȯr���|��K���l�U����>�Mc?W��>�?��?,����O�|;���ɡ=��h?���?��?��>�}�=v���X8�>-.	?���?���?�~s?W�?�Fx�>VB�;� >˘�jP�=)�>p�=��=�j?��
?l�
?-W����	������^���<��=��>hj�>��r>9��=.vg=/{�=3+\>�ܞ>a�>��d>���>'K�>�Oʾ�W�?!?�G>�ݝ>Å+?c�R>Aڽb��#��<�Ͻh�����ì���ZoV��J��F9=,�=��>��ĿKT�?^��=��6�?�o	���p<$V2>@S,>�wE�"Օ>��>D 8>�M�>ik�>K��>�rz>/R�=y�
��g=Z
�2�4���L��k����;Bs>��׾��?���s!�t_�J����p��}d�A����:��R)>�j�?���*Q�/"��¿<m�?��>�r0?����}x�:�7>}�?B+;>�fھA�[������l��?���?o|
>Q2�>��M?dg�>z�A���a�H�|��ld�m�1��n��;��)���c�\�(��4)>)�?�>z?�?\1�=� �>V6k?{�=����6�>w[<�}T�r�>�Q_><U��	=�E����Ĳ��3_�n5�>%��?y?W��>�\��¨��c5>��1?�7?��v?\,?�.?*��,2?[W>(r?z?q�1?��?�? F:>{z2=`�;�3y=9 T��E}����hԽ����j�=��=;A�=�6=���<�Y����ۻ!g�Y�&=��:y�#=5�f=�1�=��
>���>PTW?Z~�>��>�D?�I:��I�fd$�[�5?��I�T�A�b�p Ӿ�E�"�:>��p?u�?l�]?�^#>G�6�����dlq>��>�C=�^>c��>���Ck��U�=2�>Q�;>,#=S�u�˥��8v�?�����=��=���>g��>䊚��8>Ώ���N�B{d>��{�DlǾ�{O���L���/�����v�>�#H?��?f�=$�̾C^�3i��06?s6?WJ?�?�?�K=�-Ӿ��-�ߊA�r��Y��>#�=k�҈���0��ٿ7�"^u�ē�>e�����갴=n���Ⱦ�v��Ao��Ǿ���=_0$�N�{='�C!Ѿ�Ǎ�6q�=/w
��+���m0��@��%٢���v?}�6�	v�:���|
� �'>���>қ�>oB����<��<��`Ͼ�aJ=��?+
j>i������b;��.��%��>��@?f?Sr?���Oq��(G��K��A���Iv=�/?_m�>?�|�=�k�<�ɾ7�	�0�l��9�Gr�>���>�����?���޾��ҾZ�����>�i?��u>Y�?�P?��?a�b?��"?��?.ѐ>�:A�r�־8A&?��?�Є=&,ս�HU���8���E�5@�>*~)?�A�E̗>6s?Y�?��&?�hQ?5�?>�>V� ��[@��>�T�>�W�rI���_>g�J?p�>YYY?���?��=>Y5����-����=�>��2?O##?��?E¸>���>���ꂀ=�_�>_ c?4*�?��o?�[�=u�?2>�>_/�=m��>��>�	?�EO?��s?��J?R��>1��<Q欽Ͷ�*�r���O�^�;��F<F�z=;U��ct�{E�r��<� �;j���D���t���D�Z�����;�V�>�YA>�K����:>l���Gԡ�d�=��Z�t�Ҿ�*���v��Tc��>�?���>��<� >E�>؉�>y��z_%?\��>l��>_�=s�G���{�p����>٘c?���>�v��f�����^�=�=�V?��c?%M)�^���b?U�]?d�=���þ��b���	�O?��
?t�G�L�>��~?Z�q?���>7�e��9n�M��zEb���j�۶=�p�>KZ�;�d��8�>�7?AS�>��b>�%�=$q۾v�w��q���?��?j�?O��?,*>��n�;4࿺�'�Lы�x�^?���>�᣾�[?Ӵ�����g���	ti��q׾[ۭ�ہ���ˢ�x�׾Oi��y��9�O��*�=ͭ�>�8V?�Si?hN?����h��d�7����Z��l���q��YB��=���:�!d�����*��Χ=��j�"*?�E�?�-$?sF)�;��>V[��,1��[/ɾ7�>�������K�=��a��ӂ=�X="JB��s2����?lc�>�>�>��B?6Q[�`=�>�4�wD/�3���%�'>�ʓ>���>���>?��<��!��o��(Pξ$���iĽb-v>�rc?�K?L�n?	\�L-1�����!�&w/��F��z�B>�`>Ƹ�>��W�Ϯ�?&��R>���r�(��M`����	��H~=آ2?�>���>xL�?&?�o	�J:���x��v1�?ƃ<
=�>qi?�L�>��>��н3� �I+�>,h?G��>���>�8h�\%�o�~�е��`5�>m�>���>��K>�j%��b��_���[��A�1�~��=wu_?lWx��uf���|>q<?x*�¾K�oҏ>�_c�V���ι#����� >�?܇�=-X2>����
��B��/���|'?n�?�⓾��+�^�>XD?���>D�'>�w?UrO>Wr���<z�?J�X?�G?N�/?���>v�=qģ��g���,�ǈ=�Ȥ>�*>�=M�y<ⓕ��d�rJ;�g�X��=<
<�G`��	<ǥ�<9�#<^<�u$>��ۿXK��,پy��� 󾁙
�� ��lD��-���!�������䙾%�x��#�4 ,��9W��c�������m�܉�?��?;��&�������hh���\���>��q��~��7��}���֕�~߾tL��,/!�ǙO���h���e��>'?d��q�ǿJj����ܾ]�?�d ?ɂy?c�T]"�]�8���> E�<���ש�
�����οOB����^?�)�>�O�~������>/��>�^Y>r>�'�������Қ<��?�h-?��>6�r��|ɿ�Y�����<O��?��@�C?�+��>�ьú��>2�?�w�=6x�0���Nܾ,ݚ>�8�?��?lZ�=y�@�mx���yl?���=tB��$<���=D'�=t�=7�5���&>/�Z>-ٽ�Tk���+�m�>)�x>
P�����JE0�Εu=��p>�s��$ڽ�ф?
f\�Zf�U�/��L���,>4�T?�"�>G�=*�,?�H��ϿI�\��a?�+�?���?�)?2���k��>��ܾ$�M?K6?� �>m&�"�t����=��㼏u��ľ�g0V�֜�=���>��>��,�-r��O��*���+�=X�7�ƿ�$�}�@_=.�ݺg�[��~�}�����T�y#���eo����Ջh=��=шQ>xl�>�%W>�3Z>gW?h�k?�N�>��>7�d���ξ�w��G����i���,��F�mR��߾d�	���������ɾFD���{=̵M�93���� � ,f��D�{+?�5>G�Ǿ8�H�F�<ʓʾ!媾��X˽Z;̻5�zo���?��8?�ֆ���V����3|�#�x�F�]?KK�0 �Q���5x�=VO���%�=볞>�[�=���61�7P��D/?�/?�6¾�H)>��ӿ,=��(?0��>K<K�>ܻ#?ؚ�r;׽U>C�/>�B�>���>�� >§����?IS?cj����l��> ^���Vw��p==s�>&<.�M���#O>9��<����c�;ڣ�N�<KT?	R�>��-��|��y���5&;�W >y�?!��>Ѵ>�ro?P�5?��W<�9徱�P����Ci=�P?� f?�X�=O���$��m��Q�;?� c?�!b>ĆY���>4�7��A�?�^`?P�?���I�w�ό�`�x�8?v�v?]q^��r��J��0�V�O;�>�\�>���>��9��l�>�>??#��G�� ���V4�Ğ?��@U��?7�;<B(����=�<?�\�>n�O�b;ƾv������y�q=� �>C���(bv����c,�%�8?���?���>ѐ��������= ו��Z�?*�?ׂ���Hg<���-l�el���<�ѫ=��F"�Q��2�7���ƾü
������޿�s��>�Y@K��(�>G>8��5� TϿ~��5WоQUq��?���>ݜȽ�����j�8Qu�޳G���H�E���I7�>�C<��м+�޾~���}>�|�@>�v�>
���:�	?�$�����05��pé<e��>(��>��>%)&��0��%�?��ؾ� п�y��81ľ gt?8{�?c'�?F;�>I�)�#����'׾��;^0r?�?�mo?���<+D�=+j<��j?_���U`���4�[HE��U>5#3?�C�>}�-��|=*>>��>�f>�#/�\�ĿWٶ����!��?���?�o�>��>D��?�s+?1i��7���[����*�4V,��<A?�2>w���)�!�*0=�hҒ���
?B~0?�{�q.��l?�z�������g����.=�>�kӼԹ �ݾܽ����`�XR����f����?Tu	@wZ�?a�Z������>���>l)׾'���/0=��?�B$?�F�ٟ�=��>S��q�H�z	>#p�?�
�?�,�>٢���o��)>>�G?�Μ>Ȉ�?��=1�>�c>�؆��Q=�r>f�>��$��?d�F?#+�>z�8=J�����NI�Q�fx����B�1q�>��e?�[E?#�>�Ľ/7����Ԫ�<jD_�]����� �#,8���I><>�=M?�=��@�$����?\p�4�ؿ�i��
p'��54?/��>��? ����t�����;_?�z�>�6��+���%��~B�]��?�G�?7�?��׾�P̼�>%�>�I�>�Խ����^���i�7>0�B?��D��j�o�q�>���?�@�ծ?oi��	?���P��<a~�g��7�U��=��7?�0��z>T��>��=�nv������s�㹶>�B�?y{�?���>6�l?m�o��B���1=CM�>��k?�s?�2o���D�B>O�?;�������K�+ f?��
@mu@w�^?vܿW �����ޫ�� ֡=T`�;o8�=a�+�}�;=}ۍ=�o߻����Y�=��z>��>cq4>� �=���=��!>��������ؗ�+^���D���+�ت��r�����?a�24�����Ǟľ=b���A��\����8z��Sk:�G��=ƬU?;R?p?� ?�Mx�j�>8����'=�o#���=U0�>8d2?�L?d�*?�=ڤ����d�`��DE���Ƈ���>�uI>�~�>�B�>y�>�N 9l�I>�.?>z�> >�W'=yE�7a=��N>8J�>\��>�v�>ו+>��> ʳ�ڮ��+k��Ղ������?6z���G�oה�,������Y�=��+?R&�=���ѿ����f�I?,������=�P��=��1?B�X?��>Dj��V;���>���{�m�@�>����&�h�۽)���O>80?��f>�5u>|�3��S8�-�P��\��/�|>aC6?� ���
9�`�u��H�\ݾ�AM>㤾>ƇB�ud��������i���{=�q:?U�?zӲ�{ް�λu�}Y��5MR>w/\>��=Z��=�HM>��c�6�ƽI�G�z.=�j�=�y^>z��>fԥ>(��9�>�m��_$=Ö?8;�>,���~T?��o?h�=�Ɣ�����o��-�>m��>L�=���fݾ��~�=˝$?Zb>��	>&�꽬����������>�I6���,�2�=��|=L���=�y�=�L�E�y��<�'�?5\��ޛ��I8�#���|�?#U�>˲=�Zm>��h跿w�Q��F�?��@���?Ƨ�b3J�&%5?�|?^��p+����>j�>�U���oc��$�>m'��6��|nN�*Ƃ���? ��?r:��BE����>��>����b�>S��MZ��H��B�u�O�#=���>�7H?>]����O��>�zs
?`?�Z�!�����ȿz}v�;��>�?���?%�m�7@��^	@���>ɡ�?gY?gi>pc۾:TZ�⌌>��@?}R?��>:��'���?�߶?���?�)>��?q<z?lO�>�<�6�����G�r��Ƣ=E�R=�u@>�1}=�ѯ��S�n��T�����Y��!�M c>�2�<�̐>¾�ah˾��<=ֿ��.��`x�����>�{�>�H�>ԑ�>���>��>Oύ>��x<;j޽��9��T�K?Բ�?v���.n���<���=X�^��+?D4?�`Z�_�Ͼ�Ҩ>��\?���?��Z?Hf�>���=��濿�~��˖<b�K>�6�>�J�>����GK>��ԾC:D�4n�>�ӗ>6ڣ��=ھ�+������dB�>d!?��>2Ǯ=�;?��"?�.}>���>�jB������MG�=��>��>�G?�={?Q�?zt���5��D���¡�`�X��5>��u?�?��>ۚ��υ���DN�)�"�n�[��_�?_�e?ϫ����?$��?W�=?qlB?�+e>|��VEҾ��
�i>Ǵ!?^X�[�A�sp%���w�?��?;G�>���uѽKN��<��|h��z�?c[?�&?����i`�����V��<!Y ��G��E0.<[��F�>/>�����c�=,�>��=Gxk��97���Q<�=`�>`�=u�8�M�����$?��C=L��h,>Z�]�/Z0�<ݤ>�>����l�H?�l<�01~�2W��-���$L��?���?jT�?�0Z;]�a�&�??5h�?���>:�>I(��� ��m��,t��u���?�3�>q��>�\p�Q�%��i���������c}�9 �*�[F?��>�?7	?�6G>\6�>�я�^C��r𾍞���cS�2I���>��(*�qX�ޤ���e�t�>9������}�BS�>d��"��>?1 1>�LT>P��>�����y>ڰ/>�h�>��>�M>l��=o�=%�A�a����m?PH��kG���2�E޾�F?�
&?7
�<ѻ;���� !�Mރ?��?���?�Ml>(oW�%�(?B��yܱ��j�?��=��b=|o��w'�qaJ�������n�3��>�ͬ=��!�Y>R���i��D?c?g3���䙾���ޱ��v]=Q�?�e(?��(��T���p��)Z���R������]��-��+`$��p��l�������v���'-��k=x�+?���?;Z�0������.h���7�k�w>9�>M��>�A�>�G>7��M�.�$(\���%�?�t�l'�>:�w?g��>=I?X�;?��O?�LL?�}�>�a�>�尾�/�>3�;qX�>��>�9?a�-?V0?.?3�+?g_d>����l��{�ؾ��?p�?�?U�?�?܃��hTýp���8�v���y��Z�	��=ӗ�<j�ս��n��uP=*�R>UZ?Rn��:6�O��؎l>i�%?9��>T)�=Q�!j��=[ѽ�>��?[Ϭ>N�Ͼ�aZ�rC�\D?�Lu?Xe�]�#���j>���=�ֹ�� ս ��<fv*=0Iu=��ͽ�=z
;i�=��T��_������c=/(<�������>�?z��>9��>�����E����=GT>��P>'�>�پk7��匘�,�g���j>e3�?Q|�?�e=f�=G��=|���9L¾�q�D���<�?+�#?��S?���?��;?��$?o8>6<��������&��̗?!,?���>����ʾ��S�3�f�?�[?�<a�����:)���¾��Խޱ>�[/��.~����0D�Rօ�a���~��ڛ�?ſ�?IA��6��x�Ϳ���Z��P�C?#"�>_Y�>��>7�)�,�g��$�2;>̊�>�R?���>�	8?v�`?/Y?��A>fu3�ǰ��G���cu�&�*�:U?�Jo?�?��{?��>QsH>�<Ͻ����S���x�v��������>A>�?>���>R��>I᫼b`	�Z@3����=���>Wu�>zx�>��>.�1>iU�=E;D?�}�>��оG Ӿ7ט�����_>��u?m�??�8?"g>��W���H����q?K��?�9�?�U/?)h�>��<�_�=5��A��!O>��>��>�<֚�=�H�=/�>:�>m���Z�Q��*���>�b
?(xb?v��>�*����q��_���ע=4����v־�cY�b�&��"վ�r>�*Y�}\O�9eپ.y/� �پ�ֳ�X+����OýVr?��.<��==Ύ=
ᒽ_hͽ���=@�;/�>�>ݺ����=�F�gg�������=�@>�m�>W,�="�QO�?Eh�?��!?��?=��>XP���=�KK?�ľ��$?Z��>U���}�.��[�lգ���c���n��@ >��/#����=qE	�ST�=�q=�~ۼ�L��.�sV����A��BJ=�ܤ���<�	>Q =Y">C��=��=mLv?<���&~����Z�}��(/0?�ɨ>���={־r�??&}+>�����<���r��[�?{��?���?�	?4J��*�>�5����9�<b+�
|>�y�=s�K�>�S>�P�,����H�"��?��@�=?A�4tɿ���=��9>��>ǘR� j0�}~Z���]�5�S�S7!?8�:�Pʾ<�>e�=u-ܾ^!ľ� (=5>g�j=� ���Z�XƔ=�ԁ�<wG=��}=xʊ>X�@>�*�=�7���x�=6:=�(�=)KP>��n���E�'��7=�%�=\>p>K�>�P?vb"?��`? C�>�C���hݾ�髾-�E>�o�=�>�>Jx��c>�_�>/�A?_�K?��K?_��>Eh>=���>ҷ�>�'��]e��L־���L��=_a�?��x?y��>Z��=N���
4��j9�<����?�a4?o�?�u>�U����9Y&���.�$����z4��+=�mr��QU�M���Hm�2�㽱�=�p�>���>��>9Ty>�9>��N>��>��>�6�<zp�=ጻ���<� �����=$�����<�vż͗���u&�:�+�2�����;s��;C�]<]��;U��=�H�>vd>;��>���=dɱ�-�>Apg���A���=���Z�7��X������R1�y�9��[R>�g>'�_�fÏ�0�?�A�>%E�=,��?�>T? #��Ǿ��ũ���w��k7���3�o{3>���=��a�o+a��sr��sI��Ⱦ���>��>��>�l>�,�9?���w=��1Y5��>Jp�����m!�77q�=>��2�;i�5պ;�D?`D�����=�#~?�I?�?u��>�R���ؾ�a0>/R���=���q��s����?;'?��>��R�D���о�TW�	�>$O��8�h���+x�V6���xо;H�>�e��Fþ'7�*�h�U���}�)�(Պ�j�>�xW?r�?J�F�N�L��!��|�_����>W$Q?�Ց>q�>��>VἽ���v�?��;U>�k?���?jݾ?�}>��=����+�>r#?Xʖ?y�?Hp?��C����>;f�Q
 >�����V�=>�ҝ=���=�y?�?�g
?!O���
�w������YX�S�=Ɗ�=3:�>w/�>�Po>��= f]=�l�=~�a>���>���>˽d>O�>��>s �����0?}��=��>^(?d>���[���qh��;����#��Q��Ǟ�����������=�ŵ=/����>��Ŀƣ�?�_`>��?U? ��0��F>T�#>.����>C�Q>��u>���>r��>�]>�s>��>Ƴ��<���Ԙ�۹X�S�������~>��
�νM�(HH��|{�)n��� �4�g��5��&�_��)=�O�?�-p�bfb� ���+��3�?@'�>�6?v���/<<��>��>y<>7��K��b�z�'c��X�?LA�?k�c>���>�W?Q?3o1�O53�+yZ���u�e�@�R
e�0�`�#���nS���J
�1���y_?vy?oA?���<P�z>,i�?K�%�vA�����>`�.�xH;���>=/��>�|���vb��Ӿ�þͶ�G>��o?�	�??�V�[j���m0>�Z<?H�0?�1x?��3?�P2?\�(�(?:� >��? ?-.?�%&?��?t>.>	��=�?���k=Є������̽�в��M"���6=G��=��;��;5D=��<"6��|gڼ�[r;�,���:�<�@$=9��=�0�=�>�>�fY?.��>��>M8?���@0B��궾GX*?�Լ4/����|�s��_��>�Z\?]ר?�eY?�!k>�0���J���>4\�>�(>z7g>�L�>�,7I�s<=��=�[�=ǈ�=e��<H�_�I���ӫ���w�<�,>���>�]|>�L���&>4��K�x��e>��R���R/S��G�EJ1��St����>6�K?��?Ր�= 辉䓽�9f��)?��;?5�L?O�?`ŕ=��ھ�h9�V2J�HU��ҟ>�ؒ<h+	������ء�NJ:�z�K:�dt>�읾̙�1Zk>���_վ��s���F�ӣؾ���=w"
�iҩ=�i���վF���S�=l��=����I#��+�����J<G?tƐ=Dh����J�TB��v0#>I6�>8Ю>�G����z��t;�$ȵ�o`�=���>P�0>��@<���~�B��@	�SF�>�QE?�W_?�b�?
k����r���B�lX��3���fü;�?�^�>�B?ƭA>^�=�����
�{�d�G���>T��>E�� �G�&Z��,���$�$��>�?�>b�?��R?��
?�`?��)?Xe?��>(帽XK���9&?ɂ�?	t�=�fӽm�V��8��E�Ϝ�>�j)?%A��*�>g5?�`?��&?<Q?��?��>#��@��a�>���>U#X��!��74`>�J?*�>1Y?���?�=>�55��q���E��F%�=Ϋ>��2?�4#?d�?&�>�Y�>��|2�=��>̙c?��?pmo?�"�=�l?Ev1>	��>�ٗ=���>���>W)?{fO?is?ǿJ?�X�>�,�<��������˵s�ÀS���;��X<��x=g��Dq_��9	�s?�<⧳;������������_uJ�y㗼�^�;P=�>��l>����3>�ɾSɇ��z;>����z��\Ύ�[�?���=���>o�?��>�o�J �=�>^��>a�-�*?J��>Qd?G+�<�1_��ؾ�J��q�>�??C�=|qk��8���o�2ĉ=3�i?t\?�O�������`?:j]?�~��m7�Ӿ�xc��� oR?�|?׼&����>Q5z?	-j?���>(q�Mg�����]�f�M�s��b�=+>%��`��ݓ>�@9?\��>Ϡt>G��=Y�ؾ�;s�e|���	?ع�?g�?�͍?ew&>��o�N8�y���#�����[?���>Xc��D(?��t�>ξs�������?⾩����j���������O/!��2����۽f�=	�?�;q?��q?�H\?���c��8Z���}��W�������+E�$�E�]A�wMo�G��E�������1zL=O��8�¸�?��?�?!��>u��i�"�ԾA��=�����f��B�>�)���=	�Ӻ���۩8��mƾ:�?@e�>�:�>�Y?O�]���<�?+2�J�1�-���m;>�p�>�ט>2��>Iμ=����ܴ�ew�;��?��Ycu>�nc?ʹK?e n?� ��0�p\��� �.(�ަ��XD>�u>"�>r$Y���H0%�3>��5s�����Ï���	���x=�=2?��>_ڜ>�X�?�?U-	�GQ����y�W\1�\�y<q,�>a�h?�4�>.�>�nνU� �Uy�>q�l?c1�>��>�g��iz"��R|�*ǽKN�>���>��>�cl>�V1��7]�lݍ�J�����6��1�=;,j?C���}�b�8�>1�O?���uOm<�o�>��8���G5侉X��>h�?y�=�',>{��\���{�*����(?j�?�����h1����>�(?�S�>E0�>��?�^�>��ѾZ�2=��?� Y?0&C?��7?�\�>�p=��
�R�ý"X�L��=M�u>)Q>DU[=���=Nh-��9���,�|�[=|J�=����n�o�/�����~�<6P�:O:>0�ٿ�L��nԾ���\�������|��7��f����н׉�������jt�z��P0��ֳK��fn�"�����X�x�?U�?�;���̌��Ś�C�}�b���J�>�����Ҽ��9]�R󢾺ؾ\���k ��CP�"�e�M\`�O�'?�����ǿ񰡿�:ܾ5! ?�A ?8�y?��5�"���8�� >cC�<�,����뾬����ο>�����^?���>��/��t��>ߥ�>�X>�Hq>����螾n1�<��?7�-?��>Ŏr�0�ɿc���]¤<���?/�@�.??��#�6���Ҿ���>Lx8?Gr�5U�
���;�t��Ps�?5�?F�X>j��1��믅?�ϫ>G쀿�슽͵>黴>���<%nS���>�4Y>�C����]��ţ��b>_m>�k1��h�-��q]=z��>߿��J���Ԅ?�w\��f�N�/�RT��Q>��T?�)�>f>�=�,?6H�\}Ͽ2�\�'-a?&0�?ͥ�?&�(?0῾dۚ>��ܾA�M?�B6?��>�c&���t���=x�dt��h���"V���=��>jy>#�,�5���dO��9��R��= �e�ÿ>��Z����<� `�?��۽B7�W�ǻ��[�c�[|ݽ��U=�v=��Q>Od>Q�;>�xi>�9]?��c?m�>��=��'�ũ��Ú��e�I�u���֡�����tv-��9���۾�8����}��D�̾�	=��e�=:)R������� �ºb���F�F�.?�v$>J�ʾX�M�k�-<�kʾ.���xf��Yo���3̾�1�R)n���?�A?� ����V�T���S�ղ����W?׏�����鬾n��=���n=��>7S�=����3��S�K/?�V?(Ͼ�1�����'>92��~.=�k,?�A?�j<�U�>�$?�&+�B��JY>� 8>�`�>G�>}�>�=��A۽��?� S?���l㜾9`�>	���VCu��)H=$�>x[3����a�V>|m�<�׍���W����rF�<�W?�>��)�l��`��������>=|�x?�}?la�>�k?��B?s*�<�n����S�F�
�H(w=ܴW?�i?ߎ>�Q��4оk����5?�e?7�N>�Ah������.��F�3?#�n?�P?�Z���h}����U��6�6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?o�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������XG�=�;���o�?�?�]��c�c<�q�ܓl����c7�<��=G'�#6+�;z��6��Ǿmj	�����K���D�>]@�%�x��>�r5����5Ͽ����7о1�q��?k��>*�ĽUK���uj��Xu�tH��eH�"���c�>ѩH=�������s��y�U�_.>��>�)�
�>��9��l���辨�]=L$@>�?`�i>����w}��T�?y߾H��-զ�Sо��r?��?t�?<p�>�h1��P���̾kg=Pj?�ڈ?�t?�չ=��8���w�W�j?�a���U`���4�mHE�U>�#3?jA�>}�-� �|=�>���>gk>V"/�E�Ŀ�ٶ�����,��?ƈ�?Bo����>%��?�q+?�j��7���Z����*�ٖ+�<A?�2>���y�!�r/=�lђ���
?�}0?p�;.��"c?��u��ko�ɺh���۽�F�>����[����*����'�p��|���ǂ�<��?B�@�8�?MS����˾l/?�H�>\������ �=?qD?Ji��
>l��>��6�P�'��<�<�#�?���?��)?^ԗ�����:>>v\?R�>��?bc�=���>��=�Y���L�G�\>�t>z�V���?�@A?g��>�=Y�&�q���E��1E�A5���D�ѯw>��d?�Z<?�>.�н�]!��.�^C
��c\�����5���������;>�>�>�,�X����?Qp�8�ؿ�i��&p'��54?6��>�?����t�����;_?Uz�>�6��+���%���B�_��?�G�?=�?��׾fR̼�>+�>�I�>)�Խ����_�����7>4�B?R��D��q�o�x�>���?	�@�ծ?hi�R	?O"��N��>_~���2+7�`��=��7?�;��z>߿�>��=�pv�������s�/¶>@�?�y�?D��>L�l?�~o���B�C�0=?M�>�k?�q?�j�x��הB>l�?>�����}B��'f?1�
@*u@͟^?�뢿	�ؿ����R��Z���+><�=]bn=��R��Ω�ʄ�=�z�<�\׻��<���=�q�=��=���=K߼y]�=����>Q"�_���z􄿸�2����7���L��L2��x�� �\F۾�n���7��� �潎Lt������L�7�=�3V?(S?l?с?WDw���>������=#R#����=9��>�--?U�G?B+?d;�=M���Re�����X���ŉ�r��>@�K>d��>�4�>Q��>'�x<J�M>ţ'>�o>� >o�=ʲ<�=�`L>�)�>E�>7��>C�<>>R>ݩ��������h��v��ɽQ�?_+���9J�o长;f��gٷ���=�.?k�>O	���Hп}��:�G?�m�����-+��D>��0?F{W?R>'���aU�K>��	��9j�]?>sH ��/k�07)���Q>�?K�f>Osu>$�3��<8�y�P��X��o�|>H6?Aö�D�8���u�֯H�?pݾ8M>�>e�8�	h������bni�@�|=�6:?��?m�������3u�GE���Q>�
\>�8=��=8SM>ڑc���ƽ6�G��/=���=�^>d��>��>i�Ľ�)�>w����
���?���>���=l�L?0'n?5*���ɽ����:�0�>
�j>	�=��k>ٷ�����=ԁ�>w8>W�b>��ҽ�E\����B��>/p��j���]�=�"�=���ëy>�:��w��z�n�"�F>���?g���,���0���vN>_��?"��>���>�9>�-"��6��cR��+��?q�@�6�?�p;��YT�F'y?���?����`�,��-�>��?������F�>n ���ɛ�B�	��*̽��?��?枙�v'��К�T�>��?e���<h�>�x�|Z�������u�6�#=n��>�8H?�V��s�O�i>��v
?�?�^�㩤���ȿA|v����>T�?���?c�m��A���@�z��>-��?�gY?Qoi>�g۾+`Z����>ɻ@?�R?�>�9�M�'���?�޶?կ�?ׅC>f��?���?H��>�7|��.4�>��ބ��=+>�}�rm9>",�<Nоq�S��x����B�. ����>M��<{C�>�7ؽ �����=|"��������=�ԭ>��u>n�>���>��>)�>�0[>��]��悾�uJ���K?h��?J���4m����<�y�=Z�VR?��3?j20��g;4�>�[?x�?v�X?�ϕ>�S�{6��
��*���%�<@�F>]r�>0��>Ԗ���M>@�Ծg�G���>i@�>�FƼپ�	��������>��!?���>Fq�=)�?�Q(?���>�d�>B�N�$s��O�P��:�>��?-+?of�? �?Kľ��=�r��h����&O��1>�J~?��?��N>򶑿����	�Z���@=�7A<9��?��A?mQ�=�-?
>y?4	#?��H?��=H(=L9��Eꔾ�<�l,?�꽅�S����[�m��>5?B��>!�ֽ.C�D�|�J�ƀ��T+4?Q`n?v�*?d&���^��թ�-�<�F�=��#8=�(��Y�>H��>=",B>��>z�>�O��M����=�o>m��>2��>5��O�<d+?n���Zy�2R�=r�q�x�B���v>$?>7���#]?�f?���{�	v���՛���N�mp�?q�?`(�?�W��\#h���=?_�?�?��>|��T��
ྈx��(w����_>���>���޾徕Q���a��� ���3�����3��>H�>�?#� ?v�I>�#�>����#�����a�d�]�6���$9���+�A�������}$������'z����>�����>Z?�-g>��>�%�>|L��W�>��S>[6}>E��>�.V>�+0>��=�%q<��ɽ�1^?�.߾��/��z�����Y�H?�/G?�iM>@BZ����z��DL?��?��?���=�<e�����??�ł>�+����h?�M�;��¼�PѻE��/���t��(�p����>-�j��H��%���ƽ��?ǧ+?�ږ������I��}4=c��?e�&?�>*��T��f��LT�0!X�nP]�w�n�ٛ����%�Ql�7���9g���T��K`*��H=�-?4,�?C��������3i�uZ9���V>G��>yZ�>!��>E	B>�d�.���Y���%��Ņ���>�Yz?W��>w�I?#<?�O?�L?W�>���>dv���u�>�^�;�:�>U�>�8?M�,?(&0?��?��*?��a>�;��F����zؾ�,?�_?�H?��?I?�V��l���������x���x�n������=�B�<jٽ$;t��Ua=GcR>�D?�n�d�9�����.?l>�58?�6�>>��>����т��&�<���>��?��>-����q�����>�m�?I��	�=�,>_�=7؇���Q��=��׼W�=������7���#<yѻ=D�=�`������(;�S:��<���>��%?�п>�<�>�脾q�
�Û�rc�=b��>�PI>�">O>ԾK���x��S}Q�M�>G�?p8�?�� >�s�=���=����:������Pf�����<,,?�?M�f?��?'
F?�?0� >8�R-��7���rl��S?g!,?@��>���Z�ʾ�񨿹�3��?�[?r<a����e;)�ߐ¾(�Խs�>�[/�#/~����0D�����������?ٿ�?�A�B�6��x�տ���[��I�C?�!�>	Y�>k�>P�)�T�g�l%��1;>��>RR?�Z�>��+?H n?i>i?�>��)����}D������D����>�g�?�?L�?��>�:�=�c�<�A�Ͼ�❻�
�zx��6�w>b!�=eNa>L�?��>驋=�	�= ��<t����h%��k�>��>�<�>DG=G�g>o5�>�%A?���>�9ľ�B�ܽ��AR��ϖ=+�?k�?)�=?]�,>����%D�����	��>�\�?���?��>U����=��;=Y�%�-�I�>j[�>��>�k<����t>���>�>������� �+��8���"?�W?��>�п�/l��>n�ձ'����=s��,���@�ֽ2�Ǿ��d>#���]%��膾(����"���X��-��׾ �Խ��?�V�;myD>��>E�F��<���>��=A�Y��b>�8�����1�1�:�>#a0�M٘<�H���j>K6>�DѾ�r�?��d?*�>��?*>i�D���P>1�-?=X�=l->?��>E?վ-�'�xm�=�	>�b���־=���V�����*�A>@���W>�f>+m�=���xq�=�C>�ܹ�E k=�t��(�=��=��Y<^��=��;x�=Sv?������G�V�k"���5?	p�>�9�=$̾�??20+>����Ӹ�Կ��]�?r\�?y�?�=
?x�Z����>&���k���]=N�`�y3]>�ܴ=W#%�>��>��->���ҳ��:Px�0��?*@&�;?���J0Ϳ�,>�w:>j8>��S�]�0�|�^���W�&US�; ?�9�&>ɾ+ �>�B�=�rھa�žs=�:>��l=�����]����=�,e���,=��h=4��>#�C>Н�=_Y����=<:=���=1�L>7��J�N�}I0��4.=(M�=�
d>71->0{�>�?��.?�f?-]�>\�k�x�;��ľ�t�>�=9#�>��q=ذG>��>]!8?R�@?%b@?���>@4�=��>ύ�>��*�ezh�P�pp��uq|=�?���?��>���<�f���O9�}䪽��?o�&?w�?���>xu�n�Ͽ-&���!���~�� 	<K�Y�m%��?�;���0�
��I�=�5>>��{>if�>�sh>=�q>��W> �>�q>f Q<|Cg=%��<�ֺ���<	��=$=���iuQ<�$=��;�o�AaV=���<�<�<��<Jp�:M�=��>>�>$m�>��=�F��qc.>����1K�B�=$�����A���c�-~���-�3�|�@>XX>r���� ��0�?��]>�<>b}�?#�s?��> &��IӾ��%f�a�Q��=�(>|;�};���_�X�L��Ӿ���>=�>���>��l>,�~ ?���w=��2b5���>w���u�g�I2q�z<����ri�6�κU�D?F�����=~?��I?)�?���>MK��i�ؾ80>�H���p=;�q�Tp��,�?�'?���>c쾯�D����:�x����>���i!`�X��m����q��3���W?�椾x�Ӿ��E�9�\�;D��y!��>Ͼ8�>��]?7�?�w�W�}���S�G2
����t}�>�?K?n(�>���>�*�>u�����gj��'��>~��?���?a�?��8>贪=OK����>�n??yۏ?��p?�F)��'�>J�
<��+>�J����=�o�=�~�=���=��?(�	?aP?�V����	����A����\��<�Ѥ=���>�	�>e�> �>F==G�=�L>�&�>��>�oT>/�>	��>u	�����$?v�=��> J/?�zk>{Y�<i��ɻ��h�(��{�����e�˽��W<c"=*4J=��e�y��>��ƿ�)�?�o>ˠ�0�?�E��=G�=�@>p�A>�3��C��>(9> 1�>*�>i)�>�3>��><*>z�Ӿ�u>�1��� ��+C���R���Ͼ��y>dr���"�������ߪJ�Y ��8/���i��{���n=��{�<�[�?5�����k�N/)��Y ��?F��>T5?���������>�'�>ᔌ>}���=7��/���p�,��?e��?Z�b>�%�>wF\?-?�2��1�`�\���x�_�6�;_�^�^���������}�6֢��W?�ey?�A?��=��f>ѳ�?�A�����A��>s2�>�{�I=T��>�(����j���Ͼ� ��3�B��P5>Jd?L�z?�6?P�@�dQ��q�2>��=?��.?�aw?v80?��9? ����'?,�.>pM?�
?Gq-?�))?$�?ר>><��=˯�;�/=U����ӌ���ڽM ʽu���JI<="��=��ݸS��<�ˆ=Nk3=2�����ռ�Ӯ�,�ͼ|�D<(X=]�=��=I�>��\?�w
?Sd�>�Y0?��!���=��u��d�0?1="A��G���\�����o9><+X?���?
�R?��v>C5H������/>%T`>�0>vm>�Ù>:���(�:���=��=%>�C�=�ݽ�߁����b���W�<��9>��?%�>a�=�M�>��ʾF� ����>�F���軽Ң`��@,��D�"+��X��>�`?�i?+��>�}߾�&=��]�yM*?2&O?5�?�S?t�=����V�,���r�C��p>�>�d�%���o���vH�iR>��>�%��O'����V>���)پ΃n���J�z�/L5=k���x�=��	��1Ӿ�~����=A&�=Q����!�c����&L?��<=᣾��N��Ӽ�%�>8C�>�"�>��V�O�v@������,�=���>k�5>��z�Q�, E���WV�>�'E?s_?1O�?����s���B�"��l���ng̼ٝ?�ͫ>V�?��B>���=����(����d��F��>O��>���.iG�eC��,o��^�$��l�>�	?+>�?��R?�
?x�`?��)?e@?ی�>n����O���B&?D��?���=;�Խ��T��9�F����>�r)?��B���>O�?*�?;�&?ڀQ?«?�>�� ��0@�H��>�T�>�W�[��`>��J?���>,KY?�҃?#�=>]w5�V����ک��f�=�%>��2?%#?Z�?�Ӹ>b��>������=���>c?S0�?��o?at�=Y�?^62>���>���=���>j��>�?�UO?��s?��J?��>���<�>���?��Js��cO�@7�;�)H<̹y=���p3t��H�|��<�ɳ;Sy��HC�����D�1萼Z�;�>��t>�����W >}ž�M�y2R>���xOs��
��4҅����=uݑ>�"?��>�$��!>� �>���>���y�,?9~�>��?iĬ=��g�����j��1n>��F?v�=�o������h�/`q=֝U?"tX?Z/��EԾ hk?�X8?q�߾l�,�ܤ�ni,=�i��h0v?�?3����>��?�nD?A��>G܃�_��������~��E��?�=r��>a����8�@��>s�=?�>�<�>���=f�"��'�ğ�����>�z�?���?�Ɇ?�.�=�w���@��߃��J���	^?��>wE��K�"?|S ���Ͼ�L�����0⾭��s���B���}��ͮ$�o���U׽F�=	�?�s?L[q?��_?�� ��d��0^�����hV�_%�!��E�A!E���C��n�&b��2�������G=�\m�e�>�pʯ?�� ?4P$�pL�>���U����7ؾL->�⩾ �����=�%�mU=�)=ҞI��t"�������?Q��>���> �>?�\���A�4Q0���5�<���;/>�>p��>��>ě�<�j$�9䶽F7ʾ�1��󠻽6v>ryc?.�K?߹n?�n��*1�����+�!�'�/��c��O�B>�j>V��>��W�d���9&��X>���r����w����	���~=V�2?�(�>���>(O�??�{	��k��#lx�5�1����<?1�>/ i?-@�>��>�нv� ���>Fm?��>�>V���%;!�`>{���ý0;�>�Z�>P��>Gyn>v0,�<=\�wd��7H��a�8���=�og?�ф���^�g[�>�&Q?0pz;�<���>�|�|"��X��(���	>f�?K��=U�;>��ž���_{��l����%?�)?�����S(���>��"?�T�>g�v>4B�?���>�*�s��9�A?4^?��:?ץ)?��>e ,>#�Ž��齘B�u��:yfu>�u�>�u;��J=Υ5�b��o�1���D=�_�=hU����G�<�
���`���M=�AQ>S�ۿHL�־����+��PJ�����2���?���<���=��ٞ����~�����3C���L���g�}����{k�]U�?|G�?)��Wۅ��n��wu��P �, �>�dm�i�f��O������E�ܾ�u���!���Q�2(h�[&c�R�'?�����ǿذ���:ܾ! ?�A ?�y?��D�"���8�c� >	H�<�(����뾢�����ο�����^?���>��E0��r��>>ԡX>�Hq>-��螾//�<��?��-?��>��r��ɿQ������<���?1�@lJ<?	A ����=�F�k��>�1�>C��<kh��F�����=�=~��?7��? �l>�	0�Pj���`?�|>�+����;�h�=&w�>-L=s���=�>[/��]�H���g�M�>(��>��:��� ;]����=>`������vӄ?�j\���e�<�/�dF��h1>��T?G�>�ՠ=��,?�3H��Ͽ��\�d<a?�(�?Ƨ�?��(?^���(�>>�ܾ>�M? D6?���>\I&�e�t����=8㼈7��f�㾠V�,�=k5�>�(>L�,��w�߾N�����s��=Oe�]ſ3�k'�3憼�;�F�t�V�u�ƽj����ߜ�d�y�$�����<#��=om>B6s>V�=>�OJ>� W?Ҹd?�>67>�;�T㤾ğվU��<z�d�������@I	��Փ�PW޾�v�2�	���!�\I�Ӿ�K=�iN�=+%R�=���G� �"�b�yF���.?�3$>g�ʾ��M���-<�mʾx���V�����%;̾ł1��n���?��A?�����W�������������W?i��%��Ǭ�U�=�?���I=�Z�>}�=�{�a
3�,gS�X{0?��?�ľ����Z>C���=�-?k��>V�L<j�>�"?f/�,���*U>�6>8��>Y��>�
�=ᚱ��1ƽ�0?�+V?2��Y������>�����{u��zq=S6>�6�{����O>��;�X���,,���U���=\�[?���>�^�F���7; )r<Lxf>�4y?��?�f�>b?S�H?� ּ`]�5�f������e=�>?��y?�bN>2�A*�&���0�(?M�?��>�k	��'��xY�>�����+?.�n?Q�R?j����Ջ��L���U!�#?��v?s^�xs�����T�V�h=�>�[�>���>��9��k�>�>?�#��G������zY4�%Þ?��@���?D�;< �^��=�;?o\�>��O��>ƾ�z������A�q=�"�>���~ev����	R,�d�8?ܠ�?���>������e��=nؕ��Z�?��?$����5g<3��Nl��m���|�<�Ы=��*C"������7���ƾX�
�̪���鿼J��>Z@�R�*�>B8�G6�TϿ��E\о%Tq�K�?���>�Ƚ5�����j�^Pu�5�G���H�����VC�>��u=��½�[վ��y��7��e�=v@�>�,o�m��>?�[��N��ϻѾ"t߻�Lq>P?v'�>oW���y�|��?j)���uǿ�^����ђS?L��?u2u?y[ ?+�<�ᚾVN��_Z���@?.�?��u?��زg��j?(^���V`���4�oEE�^U>j 3?|;�>r�-��|=>!��>k>� /��Ŀ�ٶ�������?��?fm�Y��>݁�?�q+?=h��8��W_��(�*�9�o:A?�2>���϶!�.=��Β�ʻ
?�|0? ��-�z�a?!}|������s��A�=�g�>#�|�J�˽V�=>M=�b��z������?��@㓾?<"����?Gx�>pp¾0������>��7?���>f�ؼ��>Y|�>�4 �˾D��_ͼu5@���?�S)?z���#=��'у>}LX?S�>�Ԇ?�L�=W�?Gz�=����F>���;>&p>a�6��?�\F?�V�>�_�=2-M�Q,��B���M�$�	��BC��o�>�b?;�E?�n{>�C �����u�����"z=�9�1�ѷ+��r<�@�ݽ�y3>/�%>��
>N�B�;?Ӿ��?ip�ږؿ�i���q'� 54?Ĺ�>��?b���t���?;_?y�>�6��+��v%���B�2��?oG�?��?�׾�X̼�>�>�H�>��Խ��������k�7>K�B?x��D��	�o���>���?Ѷ@|ծ?�i��l?���ا��@�~�:c�Ҭ9�n�=;�6?���],�>���>���=�v�����u�s����>�ݮ?c�?���>�Ym?��m���B��=�<���>Qzi?�
?X�D������B>)z?�X�]f��H�C�g?@��@�]?�ˡ��>ؿ"b��]�&����=wG��_T�=b�����N6�=Ӆ��vX
�o2�|�&>��_>6ڿ>;>���=��>�}��X�"�C��좏��!C�Q�����uP���92���ս�t�ʌž�bپ���<2��+`�<��*�����9N����=c�U?HR?�p?ڏ ?)�x��|>}����3=�#�k��=3�>�c2?I�L?��*?)Г=h�����d�y_��D>��4ȇ����>�tI>b|�>~A�>�#�>�"K9��I>�/?>�~�>�� >�p'=�M��f=�N>�I�>0��>�>�<>.�>\´����U�h�S�u���ɽ��?�H��1�J���#���䷾]%�=rv.?~�>����UTп�����G?�R���W�68+�y>��0?�W?�+>�[����Q��H>��	���j��� >!I �T�k�I)�$bQ>;7?Zq>��|>#�5�X�4���R��>��7΂>f);?�u��c�9���i�'�G�]��)�C>?2�>�I���+����U���0q����=�f4?�s?c�½Y������do���"H>�f>��Q=e�=)9P>�#��xW��6<�
�f=�>�Hp>u��>)�>n3�j�?��޾v�q�@{�>J�>�Ԅ>�n$?��T?K�-[ٽ&���+K��+M�>�{�>�hS>rה;�Q���r{>*?�m�>��>4k����$�q�_���>�5����V�ּse>�G���-<TE��<GE��i��*�=���?����ڛ����澌��>�yX?���>���>6�>����K���˾ޚ�?u�@ƞ�?ڍJ���e��4M?/(�?r��}�=�ؾ>r?�>�n��ֽa�?nJU��`����W���C����?k�?U���Ѥ�5s�� w�>J?g�ݾ���>c1�h)�������v�� &=��>	KH?r���qG�t�<��
?K�?��γ����ȿ�v����>5��?��?��m�bK��(�?��D�>6��?�Y?qj>(�پ*8]�C6�>�A?�R? ��><H�mK*���?hU�?|��?��H>K��??�s?�	�>�v�1X/�����U��%��=��D;�ܐ>	(>0����}F��͓��T��d�j�å���`>�s#=k��>ű��R��U2�=歌�3ݨ���i��ζ>+#p>�XI>A�>`� ?�A�>���>��=����߀�����]�N?8�?�G���]�.<���j,>
�!$?ٸ'?fW#�i�y���>��8?�oj?��Z?"�>#�w���7ſ@н�0�>��=8�?�,�>��ǽm��=���m�~�\2�>:�>�Q��ξ@ ���E��)�>s(?���>���=�A!?Ӎ"?�8g>Q��>��F��𐿩�A�is�>[*�>��?=�}?�?O鹾��4��	�������X�=tO>�y?�?���>�@��ˏ��O�G��L�r�f�!S�?oi?9}��c$?���?�,@?͇D?�Y>4�#� ��`r����>D�1?��	��0��c���'j�>��2?�|?�A���8��[0���A�����cR,?�1t?V4?\����x���%��֙=�"�;��Y=[T8���&>+�=߲��������>�d�=5��i��H
,���`=^�>�H�>\햾��)�@�(?w*=&���u�>��u���4���>�v>�J��`�V?;hӽ�y����R����p�\�?e��?z��?ؽ�l�MA?��?m?#��>�\̾m�Ӿ6:ھ5�7��i��(�{>>��>œм�4�4٠��ŧ��Az�~Q�����*x�>Ӹ�>9P?�a ?�dO>�'�>�И��&��H��g���^��<��l8���.�g��;h��V"�m���O¾�Z{�٣�>:���h�>�
?��f>b{>���>�ٻz�>�tR> =>�/�>��W>!4>
%>o)<�н|eU?w���.���׾ڇ��i ?hS?��7>�K�>��������-?Ez�?_o�?�`N>�G�=��v�-?���>��F��?��<iq׼`�^飾��=\2>f�����>4�W-\�ڸ2�14�?V?��Ὓ�վ�rǻ@���i=�6�?��(?$�)�$!R�w�o�{�W��R�I��L�g�E����$�6np����#D��k9��ו(��8)=�*?�	�?�~�R<�/�����j�;�>���e>?q�>7�>p
�>�oI>��	��z1��]�I'�`���HH�>��z?���>�I?�<?�wP?�kL?���>W�>^6��*f�>���;���>���>��9?H�-?I50?Ex?�w+?R:c>8���������ؾ�?ݡ?H?/?x�?$�����ý���[Qg�ҩy�R������=��<��׽�*u�3�T=T>3;?����Z9�������k>X7?p��>Q��>rS��{}�����<l��>P�
?�ُ>F�����r�D��[��>oQ�?�|�n��<1�)>&.�=Gk������7�=g~ʼ�&�=�c��[G8�*�<TԾ=R�=L ;��ݺP�?:��M;k!�<��?g�?:r�>�i>����͕��g��"�*>U�=��>��=�Ǿ;��`����
T��A�>�R�?��?�>/Ap>A<)�I� ���޾S����7�?>��*?uO?F�R?l��?}(B?C�?���<�i,��K��a��撾�?c&,?Sʑ>F ��Fʾf���� 3�Ϙ?.�?�a���Ϩ(�Ѷ¾a-ֽ�>�D/���}�ͯ�SD�R�������t���u�?#ɝ?1+B��6��s�
�������C?��>�	�>�6�>P�)�� h����Iv;>�7�>7R?�/�>2�8?� R?ǥL?�`2>�F�Ͳ��II��C�#��l=��?�~�?��?��?���>�N�=n�������z���f�<�d�⁌�7h >�R>ْ=>^y�>2��>�d�=}0�܍�=��U�c��=ߓ> ��>ˌ�>8�&>9�>Lt�>�+H?\�>Ӿ�9�'v����K���#}?��?2�#?�U�=���-G�ɉ��`#�>ᘤ?!��?��? ��*��=Y�<����݈0���>�c�>=��>z�<l�5=j�2>��>Dt�>*�����i@��q���?'pS?��>�پ�1�t��˽�aM���־GF�c����=��7����t1?ȣ�V�Խ�h��]&F��6'��Ӄ������޾[s��3�)?ቨ<EP�
>���T��=��>"U�=Z�>M��=�e��,�<?�<���=*�ϽCý&d�bѹ=-��=�j����?�̈?�'-?�>H?�>l�οA��>��׾��,? ܛ>D�G���1��� �Om8���=�>r��	��.�f9��N�N>Nz��#>��$>�D�0� ��h�v��;���e��=f ��lm=k>�=�&>~��=cI�=�!q?�	��氙�"It�9B�`r-? �>�=Y�˾a�J?��>����޽�"��~�?y�?-�?y�?,9-�)ǽ>7�¾��"�_C{�݀M=E<�>���:�����>wn@>���&[���L�����?�@�iI?��Y�ſ���=��;>G�>�S�t�/�t�c�v�X��V�N�"?�r:��W˾�W�>pv�=���ƾT�(=E8>�tv=��W]�sl�=.�[�`�:=VF�=Ɠ�>��>>Ș�=�2��B��=�TX=���=�OK>�Ȥ8�~R���P��==��=�n>U�/>>��>'�?c??�fW?.��>��s��þL־�<�v$>�L>ċ=�(�=�́>Q�,?��A?ϋj?B��>]�>#N�>ul�>	#"��}l����'��T��=	��?�Xu?T=�>�
;>n���+��Ol�T��?u�?���>,�>f�Z�ٿ���WO:����� ���N=w���#�&�=[��F(��P��|m>��>��>�l>�>�E&>���>{`�=�o	=_���뽪��G�A�11>�н=�ܟ=:X����<p��;��C����urʼ�E��|,<	ĺ���=u�>�>w�>�P�=@���P2>����ЬJ��2�=w��4B�7Qc��_~��N/���3���B>0�W>7戽�=���f?�4a>�@>��?:5r?�>$��IJӾ���i���P���=r�>sU=��;��?`�*#M�
RҾ��>�ݎ>Y�>V�l>),��?�`�w=��za5���>��������0q�R<��D���%i��ڿ�-�D?C���j�=�(~?��I?�ޏ?�n�>�S��d�ؾz0>�H��� =���q�tI��|�?�'?u��>,(��D�:���8�&��ژ>�`���P�;ߋ����RT�;KM����>i×��#ƾH{4���v���0���z�Yb�>�)X?5�?��-��Wv�S�z��6 �pc�����>T_?��O>S��> o�>�㳽z����K�+>.�}?��?��?Հ@>\��=�Գ�u�>1�?|��?U��?;s?�U@�k��>'{;�>�;�����=�>��=U��=H�?��
?i�
?Vٝ�M�	����s����\�J��<��=��>ƈ>8r> ��=df=;�=�[>+Ğ>�g�>bd>R	�>Ȁ�>�b�����ʰ"?���=��>:�/?t}>5�)=�b���ٵ<d2p��<���$�s�����K<�:~.x=��ڼ��>�%ǿǢ�?&�R>z%���?؃���|;�S�H>K(S>�Bн��>�tH>�.�>���>�c�>��>v4�>Ŷ&>�oҾg#>8a��u��hC�5�Q���ξ�wv>A������`��N����+J����$�:Di��避�<����<`F�?:=��^�j�}�*�F�����?��>��6?HÊ���'�>���>���>jL��1l������ʏ߾|�?j��?Q�c>��>�JY?sH?��*�A53��yX��v��DF�c^�~�c��B�� Ā���Q��|H^?6~?|�>?�i=��q>��?0��H9���]~>�,���4��>=���>������O��ɾ�ľ�@��B3>�	i?�2�?�?�K� do��F(>�';?�1?�]t?��1?��:?@��$?�X2>� ?�r?Z�4?H/.?�
?�22>���=���x�$=���������ѽl�ʽ���v�5=y=�H���<��=��<�m� �ۼ��@;�����H�<o/9=���=�W�=� �>'<Y?^( ?���>TX0?<��r5�>6ƾ��?�/^=�����m��������羢�>j#d?ů?L�T?�5>�|C���Θ5>%{Z>���=n�@>>��>�h���(��O1�=m�>�+>�e=����}�����bm�l~=��+>}�?�@a>8�Ϻ�9�>6�9���N��NM>����.��wV5��F���U�N ����>��W?��E?Y�Z>Օ����=�Sc�N8?��L?�*?��D?��\=޻��i��<��?�L�=Q�V>,���C���p��G�)�N�>^��>vYվ����b>���֥޾n�S�I�7�羹�I=���T=>$�b�վ��~�^��=
>]���� �s���
۪�� J?�j=MाptT��L��6>�y�>na�>��;��&u��O@�������=@}�>Z;>	������@zG�P"�hL�>�EE?LT_?n�?5���	s���B�Ф��a��]Ƽ��?M�>)s?�:B>>�=�n������d� �F�2�>R��>�����G�6��&����$���>�.?͘>1�?3�R?]�
?^�`?}*?�D?:��>���۸��A&?j��?��=��ԽɻT�i�8�@F����>��)?ӱB�췗>j�?|�?��&?�Q?T�?��>t� ��@@����>�Z�>=�W�b���`>�J?8��>�=Y?=Ӄ?f�=>��5��뢾fݩ�K\�=�>3�2?�2#?ʮ?߯�>���>
����=��>�c?�0�?:�o?Z��=��?(;2>���>��=̛�>���>(?sXO?��s?t�J?w��>���<�7���9��LCs���O��΂;�fH<��y=%���7t��H���<hֳ;�d��H�����ؽD�����E��;���>�}>e�Ⱦ��>����J���p�=�����r�,���qܡ��=>yD�>(H
?o9�> �o����=��>��>V����&?G��>�?@�=?�o���Ҿ����� �>8IA?�<=��[� ����m�q/�=��W?V?���ʛ��p�c?�jY?�
��)C����,Y��ܼ�V�i?2��>(q~��H�>\�o?oC?�u�>9!s��d��Z���q�-�$=i��>�w6�WXA�u��>lK0?[1�>[� >��>6-׾o�Y���s�0��>�z?+X�?�R}?� >t2���~��7��S@��ݺY?��>7�����?��=eB۾��x��WھԆ���)��'���6N��]���ㅾEν8�=d�?y=o?2�o?��_?���'e�!�[�󀿪�O�e����r���D�-�G�-�?�.�h��Z���Q�����<�#���8�7��?�k?`�Z�P��>�l��8r��*�>��=I�ƾ+zj��,>�DһF]�=�ӓ=b��/�6��� ?�Ԓ>a��>��i?]�G�L8�|o���;�Q�R��>�h�>��?>[�>=@=������=�E侼���m%�=�v>��c?N�K?��n?�I��1�݂��8d!�%�-��{���LC>�>-��>��W��y�v%&��G>���r����T�����	���=�m2?���>��>\<�?��?�	�,����w��k1��S�<�G�>�i?���>7��>�н� ��5�>{m?��>>ԡ>���!
!�t�{�'Ľ���>�G�>�q�>�dp>E-�F\�E9��&��`f8��7�=��g?����`�e>�P?(i�;~1n<�o�>�w� �!�����ؼ%�C�>��?�k�=D�<>�nž�n��3{��c���&*?�"
?|A��O �>D?XU�>�)�>�r}?x�>��ʾ�N��?�2a?fUM?�cC?�Ͽ>&��<|�q���˽w��(�=�8~>݃D>�qf=���=b���i��(�x�X=���=u!X�B'��,�8<�猼�m�<�=�|3>lۿo\K�$Eپ����#�m
�����p���I�����5V��l��G%x�̨��K)��RU�Vtc������Jl��i�?��?2����������_����Y�����>&�q��C~������"��%��S�ϧ��l5!�ʴO�mi���e�P�'?�����ǿ񰡿�:ܾ4! ?�A ?4�y?��4�"���8�	� >�C�<,����뾬����ο>�����^?���>��/��v��>ߥ�>�X>�Hq>����螾�0�<��?=�-?!��>Ȏr�1�ɿe���D¤<���?/�@�D?��6�s����㄰>!�?��쌾�c �n��ӂ�ƹ�?�{�?3M�>�X�]�ݾ?��?��i=M��fl=o�>/��>z����o��>���>ڽ�����f�T���>�>����Z�qs����o>G��>F&��}�b��҄?j\���e�/}/��C���3>��T?j!�>�;�=�,?Q-H��Ͽ��\�C<a?�*�? ��??�(?b濾u�>2�ܾAwM?e)6?��>�w&�*�t�?�="�el��h��	V�U�=U�>�>�`,�Y��yO�/+�����=��Ihƿ"�#��v�OX�<��ۻ�S�8���4��8�J��T��I p���潠�\=�~�=�NT>+#�>�T>�qZ>�"W?��j?�X�>�,>U���׉��ɾB�������
�����'O��ɡ�n�꾪I߾: 	�����k��Sɾn�<����=�@R�����7� ���b�~F���.?w�$>��ʾ8�M���0<<}ʾ�����h��2$����˾�1��n�ҷ�?@�A?�ꅿ!�V����������vW?
Y�ڙ�������=���`�=>?�>�+�=�z��3��S�SF+?�
;?������۳�<N���d��=1J4?m?Vv�=���>J*+?A��������>x(K= �>]֯>9�Q��n���ҽ��6?(�N?��{�S5Ǿ�>����|�½�m->mz�=������}=�>�'��g�T���=V��<F�%=�5Z?�>�9�W0�>�ᾅ��<2�W=��?�F�>��>�j?�[/?��&��A�_>j�����r=�.a?��u?�Z >]�]����|�ؾ��0?�p?�j=>���������J�w/޾&)-?¨_? �#?�=���jɜ�� H�.� ?��v?s^�xs�����M�V�e=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?U�;<��R��=�;?k\�> �O��>ƾ�z������.�q=�"�>���ev����R,�f�8?ݠ�?���>������?��=�ٕ��Z�?~�?����=g<7���l��n��c��<�Ϋ=f�F"������7���ƾ��
����-࿼ݥ�>?Z@�U�[*�>�C8�U6�TϿ!���[оXSq�s�?'��>�Ƚ����/�j�|Pu�H�G�!�H�ʥ��(�>�%I=r5��u�/�V�b�u�&_>d>�4=>��>.^�������v��;z�N>��?͹�>*�p�|v���u�?��ھ�Dƿ�Π��^����q?T��?��?R-?Y��i6z���'�<��}?�A�?��K?s�ýe��U<�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�^�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*�N�+��<A?�2>���I�!�C0=�TҒ�¼
?V~0?{�f.��Y?( a�~j�0G��nĻGNw>��F=�����>=~L��V�>X������l�?��?��?U�2�%+(���?���>[�����[�R>�S�>:`?~=���=>D�>��"���S��!>3a�?�1�?�R?�_���ک�vc3>���?f��>�ن?`K�=�\�>Ϙ�=�ߘ�Ȕļ�Q>�a>���tK
?i:K?�v�>&�o=��(*�Y�@��X�ʘ	�*A�uS�>�}V?r�C?�>T����9��"�A<ƽ��0�m_}��(���_��(��N>h%>�o>03��Ҿ��?Tp�1�ؿ�i��p'��54?K��>�?��`�t�����;_?^z�>�6� ,���%���B�^��?�G�?A�?��׾�Q̼>$�>�I�>�Խ!���`�����7>.�B?F��D��h�o�e�>���?�@�ծ?ii�c	?���L���b~�m���<7����=��7?�#��z>���>�=�qv�t���"�s����>2A�?�x�?��>
�l?�xo���B�-�0=�Y�>��k?�s?z�j�a �4�B>ְ?���N���\E�.#f?+�
@�r@~�^?&뢿?�׿D>����l��T4���>�L�=�E>3���N�=;D�=�ݽ&����G=�>��%>N[�>�+>��Q>7�j>r:��c�#��j���gy�x�G�y.�H��FOξ��	�hK#�K,�{~����f�������=�w����-��E��]��=ӕU?uR?,p?�� ?Ĕx�A�>�D��t�=��"��ׄ=(��>�n2?��L?:�*?Uk�=�*��~�d��.��2���q��l�>��H>͢�>�O�>�8�>�?:�7I>Ɋ>>iu�>�r >�%=�:��jw=��N>�ܪ>��>���>U�<>�>,Ӵ��%��l�h�mev�*�˽��?�]��/�J�^��j���ͷ��ў=a_.?�R>���Hп�rH?ᡔ�fC��'+��(>�0?�FW?t>hհ�V&S��D>	����j�\� >1���Jl��`)�hQ>3,?abj>S&}>��5�37�2oP��<��z�z>07?*ҳ��9��0r�fF���߾*�E>�<�>��j����������~��$k��=�I7?l�?֫�B��{s�񮠾�U>�Cb>�=7�=�J>-�BǸ��JG�U;N=ڜ�=�xU>���>P�>���I�?_� �t"l���>/\�>��>V�A?�G-?U�-��i�ZSھ\�@�N�B>���>�r >�����R��?�C=jW*?��U>jJ�<����t.��5�޽��>�-��q$�Rå�$�=[�5��A���;>�b��x<X�cƫ=��?rd�������ؾuՕ=�46?@��>vBx=�C>���G���"��ݗ�?H�@�ǋ?�E#�t-e�2|#?ޡ�?�_F����V>�>Ǧ�>vB��ue���L>��G=�����:����G�?nR�?�\���x��Ҭ��&I�>��1?3`�Mh�>wx��Z�������u���#=U��>�8H?�V����O�S>��v
?�?�^�ᩤ���ȿ2|v����>W�?���?b�m��A���@����>7��?�gY?noi>�g۾O`Z����>Ի@?�R?�>�9���'�x�?�޶?ѯ�?
I>���?�s?Yc�>s�w�S/�&5�������=\U;Ir�>�c>�����gF��ӓ�7f��B�j�I����a>Cl$=��>a(�>��]��=ǿ��E����f�㗷>
q>��I>oV�>�� ?e�>0��>@=����߀�>�����H?|�?�/��<\�+<�ŕ>hi��1?�/?Zb,��E���>�7?v�^?v�X?{gc>?��UB��iS���蹾�6�=��=��?u��>�Y���>>���V�� �>w��>�^�<r�Ծ�Ң��~=���>�^,?p��><�Ҽÿ ?"�#?��i>�n�>��E��ޑ�ֆE����><H�>�:?'�~?��?����p3��+��t����[��P>�!y?eG?dƕ>|�������A�:�L�?�������?�Sg?r!���?_�?�l??��A?�e>����nپ�,����>�1+?P|�����"Ծ� \=Jb�>X ?�Z�>�^/�R��=m`ʽ>cB��mx�&?@�k?�F?��:�l�d����S�;�_= �8�hE��د�0�>�4>(&A=DE<@B<=#��=s������h�=��>g2�>��>{k���V���:,?+F��ڃ��"�=��r��vD�ֿ>\L>v���A�^?HX=��{�$���x���U����?���?'g�?�#���h�7!=?3�?F?F(�>zE�� �޾t��+Kw�בx�8s�g�>���>�l�2�#���ŗ�� E����Ž{����>�t�>�A
?���>4S>t\�>�ב��;#�������
[�uM�L�8��,�~q�ԥ��3*�d��J�¾�{w����>F���r�>&?�Ue>b�q>���>�D�����>��R>�w>�\�>O(^>~G)>R��=��<�gŽ�eP?|����6��������R?ݗ?��>8�-<����'���}A?���?���?#I>��m�Dd;���>��S>C���ǘC?B����
>��=�� �\������P�@>�s�>�	�d�B��'5���'�uZ6?�B�>�!�G��6o漁����n=vK�?��(?Z�)�"�Q��o���W�oS�'��1,h��o��A�$��p��폿tY��� ����(�6�*=��*?��?���K����&k��?�PZf>�>% �>�;>2ZI>�	�F�1�'�]��A'������P�>�O{?�"�>�I?��;?��O?4L?��>[��>a|��ؔ�>�Ǜ;v&�>��>�8?x�,?��/?t?[�*?��_>���/���	�׾{�?&_?~R?&a?-n?C��9xǽX����I�;Ey����C�=�}�<1�۽:���=LR=�U>�X?�o��8�����q�j>}7?�x�>���>���'���3�<��>֭
?7�>����9|r�b[��M�>���?!�t�=d�)>q�=I	����ຈz�=�K¼��=xY��n�;�6-<���=�Ӕ=5u�b���#�:g֋;*h�<��?@�?���>Y��>�O޾tϾ���?X>dT�<���>��)>"�����ٖ��d_��D�>�L�?�!�?#>#�h>6K�=\���`n���������5>��?U�[?��$?�?�XE?j��>��>J<A��Qv`������?e!,?ꋑ>�����ʾ\�2�3�s�?[?�;a�e��;)���¾��Խ��>BZ/��.~�����D����|�����ϛ�?���?
%A��6��x�x����Z���C?n!�>�W�>��>��)��g��$�3;>���>�R?�j�>la$?x{w?wZy?io>�`�ES��D	�+]�>z?ɂU?(��?�Et?k�>��>��_��D��7������@�r���>���>��6>��?��>��>��>)1N���ݾ,F>���>}��>���>?�>G�)>��>��G?1�>ۅ��]�](���F���A��nu?�?z�+?�=���x�E��������>Y`�?�ǫ?Z�*?�R�+�=�ּ����ɔq��N�>I|�>��>�S�=�H=?�>oI�>";�>>������8�M>N��?0F?i�=#�˿_lv�χ��1R�m�6����:r>I)��_7��/�>�EH�^i��Ĕ'�>)��H���F����>>�K�Z=�?���=�5�=��==������w� �D>`2��k�1=ҽE>�ھ<4 ���'����W=�'�J䡼]�h=HAy=��<�cݾ��?Cg?rYh>��?@o�>#�c�wɱ>�y?��^}?>g�>z���}��ݒ<.�a/��e�߾����u)M�ò��>6i��s�A>p}�=@/�=���a=9=��<=��=������.L�=���=5�=t�=([0>~n>��u?^��̥���T�"�ݽ��5?X�>$R�=�\þNA?��;>>Ʉ�p���+�	���~?I��?R=�?��?��g�;��>�����|��/��=Gŉ�W|F>�B�=x*�w��>�H>s���7�������U�?#�@"<?{ϋ�jϿ�0>��T>��U>+~j�e]��p�E�C��&l�j�?�%!�U�¾�'y>�|&>C�_�̾²�=
�=���=�+��pc�aSI=)�a��Z�=茕=�pw>Up�=
>�e���=+��=���=�Ab>,���P�ؽ�&����<��.>���>fY�=�p�>y�?j>?fYu?���>z2�üϾ�/���<�)o>�2e>@챽��{>��>�H:?M�W?��?���>��L>	��>+Ϝ>�l�	�P�������\>�,�?[�r?q��>��=�_����a,5�>���
?��?H�?��>�Μڿ��{������gn�CO=Z��َ�������z1��X�\l�=�A�>��>6�>�k=>�>w,A>���>�$'>�<�=�J�*r�:�Y�=�>Xᆽà�<v.=w-�b�"=4�Y�gkJ��s	��L��� ƻ�����=p?��->�p�>w�<�����U�=������@jk=��C�F%�x=X�_���P)��?�{�Q>�� >i�۽]��d��>�Ջ>��<��?�z?-�=j�����0���Y���Y��=Am>>�ɽ�C6�;�f�k�@��0�����>\ގ>�>F�l>5,��!?�Q�w=��	a5���>|}��������6q��>��U���ni��LԺ%�D?�E�����=�~?��I?��?ň�>U��Ёؾ�;0>,E��I�=
��(q�ob���?�'?���>��w�D��MվV�؈�>��6�sqO�Ġ��Q&	�a���?���P�>�7��V�ᾅA:��	��y���&��B.�9�>�hC?t��?�t�dTn�h�j���澉�̽���>��`?☦>���>z��>q7���	�>����
>��x?���?J��?���=1)�=�Է�V��>#>?+ǖ?9Í?_�t?�z>�vJ�>4�<��>-�ڽ�D>��#>��=�9>�i ?�F?�?j���|���N��[Y_�KP�<���=O�>nO�>ӽa>Ru�=�M'=#<n=�*d>㡠>C:�>�-a>�L�>X��>`���t��E#?��=�r�>U,+?�Ax>��<�Ͻ��	<\���l�*����r������<��<���=���N�>�ſ{@�?b>|"�k?$�����X�;>��U>�|ƽ�>��S>؛|>c�>8�>kW>l�x>n[(>�PӾ�u>����e!�+C�g�R�m�Ѿlxz>\���&�ԝ�L����@I��n���h��j�,���8=�u)�<�G�?u���k�k���)������?�_�>�6?ь�2���>-��>iȍ>cC��􎕿ȍ��d�3�?]��?�4f>:��>��Y?�}?�6�Ë'���^��o�E�F��\��_��_���
���
������a?��r?MxG?G�=�r>��~?2���+��̍�>�>*���3��f=+�>�ڢ�� _���ѾC���2�A��.>-�l?��?6I?�V��bn��]'>��:?�~1?�Zt?u�1?ci;?5+���$?/3>�a?�y?�%5?q�.?7�
?�1>���=ʦ��(=�<������ѽ�-ʽ'`��3=�1{=�A
�9�<��=^w�<o-�ۼs;�ܠ����<1�:=��=�8�=A��>��Y?��?+E�>�'?�����F�����?�̣=jo��竗�u6��n���oC>n�m?���?�^j?@`>4w>���$��K5>?�}>j�>7�c>�h�>I8��4m����=[|	>4��=�I�=A������3���7fs���=��>]v?�R>�k~=�ڵ>L�� A���=D�k����.�o�S��9A�s�?J"v?��>?�y������@b>�ZU��K!?��(?C�?�B?OW >��@�����9��-�w)P>��3>��p��*�}���'�B >���>����������5>E���-Ǿ�u� �?��h��y=D,����=�+
��׾:�[��v�=���=�KϾ�h$�_B��X����P?$�P==���i^�k��	/O>\ٸ>���>�O����c�v`:������u=���>�CI>o-�cPþ�WD��#����>��D?S*_?u�?A|���r���C��0 �.���dҼU�?'�>��?��E>MX�=�e��r�Nd�G�hQ�>5�>�����E���������K�$�Q��> 1?��>~�?1S?FN?�`?��)?�?mM�>y�����B&?���?U߄=��Խ�T��8��F����>�~)?��B�	��>�?ӽ?��&?��Q?"�?��>D� �xE@�듕>&X�>��W�>`��V�_>D�J?֞�>?Y?2Ӄ?o�=>y�5�/񢾗ީ��J�=�>�2?<7#?��?\��>r��>�������=ʢ�>c?�-�?��o?~��=?F2>*��>:ɗ=��>\h�>�	?8UO?��s?��J?u�>��<mS��t��X�r��lP�K�;�9G<��x=���4t�]����<���;���Գ��X�4�D����g2�;��>P[i>(�����~�s�阾��_5Ht�Jb�>�5�K����K�D��>�	)?�.�>�>���.ڽ�B�>yR? �!�?�?}?|�>�|a�#���㰽��>�cb?�p�>��J�����2M����ٽ�$I?�%J?c�|�����>�`?�	O?��޾4�=�[��x�Λ�-�\?�F�>��(��>}Us?ӄN?�M�>L�����a�T����m��k���>�Y�>cB9�3�I�?�>_?9��>-��>��C����e�W�4���w.�>�y�?S�?���?�-�>:�w�������*��Ϡ]?&��>����7�"?�޻��Ͼt:����]E⾫C����%���RN��w$��̃���ٽ�ؽ=L�?A�r?ːp?��^?ne ��d�3^������U������ZmE���D�iEC�0�n�P��3����%����G=�1�=�2��?[�>�+D��L�>��s0!�}�쾬��=�q���̬<bKS>�.�=2g:>���<��v}	��*��=�"?m,�>�>�jh?+bi��DS��	8���=�ș�əԼ���>$��>
?��,>�q2��c����~����{7v>�xc?S�K?{�n?Kp�+1�����?�!���/��c����B>�j>*��>%�W�ٝ�F:&�dY>�=�r�t��$w��/�	���~=q�2?�(�>��>�O�?�?�{	�rk���kx��1�,��<01�>� i?A�>�>�н)� ���>��l?���>��>\����{!�O�{�^�ʽ��>W­>2i�>��o>�,��$\��a��_����9����=ȱh?Wm����`�~��>��Q?��	:��C<[��>�Us��m!�/��Ҫ'�>�w?4�=��:>}�ž�B��~{�f���x)?q<?���*�ܕ>g�!?Y�>kI�>��?Υ�>qVľ�P���?!�^?�J?��@?���>�4"=(���Ƚ��'���7=>�jZ>U�h=��=���o[����sL=࠸=7@ۼ_a���[<Q⵼lQ<!��<�X3>y�ݿ�T���ȾԆ��� �m���ꉾ������~�/���v¾n�����v��)x��=�^ӡ��ú�O���G�?�"�?QN��EY������:�f��N�����>Y��ұ�=��h���L��������5�(�r�M��?a�O�-�P�'?�����ǿ𰡿�:ܾ1! ?�A ?2�y?��9�"���8�� >�C�<�,����뾬����ο6�����^?���>��/��j��>ܥ�>�X>�Hq>����螾l1�<��?1�-?��>Ǝr�0�ɿa���u¤<���?0�@�B?�J�nO�p�=L�>LG? =�>�<�%��`���9?�)�?�'f?��<X�Y�CC��(��?�Z��[�������e>��<��>�.���:>P�[>�i[�L?��&���>�>R>��
�ji��?��2�U�骋>�0�;yh�=5Մ?{\�vf���/��T���T>��T?�*�>�9�=��,?H7H�]}Ͽ�\��*a?�0�?��?�(?+ۿ�ٚ>��ܾ�M?mD6?���>�d&��t�>��=n5�#~��7�㾶&V���=��>��>�,�ǋ��O�eK�����=���5>ƿ5	$����2o�<�#ʻz�b�A������ju>�y��`q�S߽cjJ=���=s�O>��>��M>O�[>��X?�Pi?u�>
�>���=O���BɾL&������֊�������
��s޾� 
��0�K��Tž�=����=YR�)���� ��b��KF�3�.?
�#>�ʾ6�M��P-<6Bʾ������������-̾v�1�8*n�3��?��A?���j�V������E�����W?���������շ�=�᰼��=�P�>�m�=�T�"3�.uS��<0?y�?m���8+���!$>[��\%=V�,?���>9�;6ɮ>?v#?��+���ƵP>Vr->�E�>�m�>tK>�Ѱ��Խ�?XzS?8����n��>����@�s�iUS=Y�><7�}jۼ�W>�4p<�ȋ���Ȋ����<��V?�:�>|*�<��Cg����A�M=J y?��?���>��l?Y&B?-~�<����T�������=�6V?��g?B�>�,u��	Ͼ~ܥ���4?d?XM>�Gj��D�75/����r�?knn?F�?"����}��&���p�:�6?��v?s^�ys�����T�V�Z=�>\�>���>��9��k�>�>?�#��G������}Y4�*Þ?��@���?��;<�����=�;??\�>˫O��>ƾ�z������֓q=�"�>쌧��ev�����Q,�n�8?䠃?���>$���������=�/��`^�?��?��:�B<�v��&l������}�<��=�����)��&�7�z{ƾ�
�Ww���̹�x��>-G@��+�>G�6����%Ͽ5����Ͼ��q��?���>��Ž����j���u���G��VH������[�>.>������+���u=8���?&�>��e�u��>�C5�����p����;��n>���>��~>?0ٽ)`��2�?����S/Ͽ����jk	��Pe?���?���?�l?�$��x`�/zw����:\�N?7/w?H�Y?ʒ��=ҁ����j?�V��$V`��4��HE��"U>�#3?�H�>l�-��r|=5.>
��>�b>U"/���Ŀ�ض�5���r��?φ�?�r꾩��>���?�q+?�h�D7���[��E�*����99A?�1>0���ѵ!��/=��В���
?�v0?By�-�Q�m?*���ow���7�]e/=~4�>�XQ�鲾� �}K�;�@U������>��²�?A�@��?�G������?|m�>w)��벦�cOK>���>{O>�׶���O��Њ>g���d��R>�D�?���?.�?�������|�t>�t�?̍>颊?���=�j�>f�����S��=q)�>�%�=0 ���@?��?��>#�#��,������z/�r�T�k���a����>'j?��?���>�څ�iWw���9˽�0>�s%5��B��G�`��,�;>�mA>Z��=�����Ⱦ��?Sp�1�ؿ�i��Pp'��54?H��>�?���t�:���;_?>z�>�6��+���%���B�_��?�G�?N�?��׾�T̼U>A�>�I�>�Խ-���a�����7>,�B?5��D��h�o�J�>���?	�@�ծ?ei���?�p ��$t�����Ya��j�>�w*?�9��5�>#��>^�{=�dy�t˞�l�{�WF�>�&�?�[�?ԫ�>?c�?�t�c�J��a�1�>E
d?�?���<����@>��?��٘���辙_?�+@�@�"K?`�����׿�����������=��=&�#>1�ؽ�м=C�H=�����¼�x>�Q�>�\>w�r>H	>>�Y.>��$>3m�0+ ���������K�j���Q�=�b��#�G�X�-<�f��>W���н&��1��3NS�M�0�(h*��p�=j�U?]R?��o?ѐ ?�by��>���L=�2$���=GL�>V02?�NL?�U*?ʓ=$H���d��`��Yc��?������>�*I>��>pE�>a�>n�:YJ>?�?>��>R�>σ'=t���=��N>��>r��>DJ�>��E>��>l���
����j��e������?�:��ĝI�Ӣ��%���`0��z��=)\,?%P�=���Іпi���� F?MX��'��%��^�>?�2?1W?�/>�	������>^�E!l��x�=�(߽Hfd��o!��D>'�?��k>8`y>�3��E6�D�Q� 婾��>I�8?P���[�>�u\q��]G��ݾ5�G>�ú>��I��u�}��dɀ�p�n�Nы=߃7?M�?,7���|����u�c���^�S>��T>�g0=�q�=2_H>�}�)�̽�C�AmX=��=�c]>xU?��>bؽV��> �ѾX? ���>e��>�7=K��>��I?�c���ֽ�G����Ͼ��=ɣ?� �=7d<�b���?>�C?��M>2Z����C��:�Dj�k��>g��ڝ��V1�����=;3���=ܬ>�������&=�ы?�͸�*È�U�Ͼޑ�=�N?���>嘼��=~?徘խ��U�P��?L@�ʩ?���Ŭd�ҡ8?1�?>ƽf�m>H��>��^>�����f*?���>�zd���2�Ǹ�����?�1�?���x��F�y���=�i?����g�>�w�Y�����z�u��#=��>08H?SV��V�O��>�]v
?�?�_����2�ȿ�{v����>��?���?S�m�mA���@�r|�>���?�hY?gti>�j۾�]Z���>�@?�R?[�>�8��'���?ܶ?/��?��H>d~�?�s?��>�iv���/��C�������{=E�a;���>7K>�$���pF������Y���Yj��n��c>l�#=r+�>�T�������=2������2^�S��>3�p>}�H>�*�>p� ?���>��>H`=w菽�=��=ϕ�[L?�i�?����m�s�<���=U]Y�0Q?}
3?��s�F9ξ�V�>H�[?mQ�?�jZ?�ғ>ؠ�ق��PG���e��gV�<�F>I$�>�H�>6�����J>i|Ӿ�C����>5�>v���'Lھ����ƻsɜ>��"?3��>���=Ɇ?>f?~�>�Ҏ>�oF�ר���X5�~��>��>��)?ڀO?R�
?��Ծ9]@�N<���柿��Q���]>4�?�&?�5>�T��͂��L�2>ш,>yɊ?:
(?��=q@9?�C�?L�/?7IK?�4�<��˽���j����=I$?���|�A��"$�:��?'v?x	�>�ҽ��ʿ��@L����m�	?E�U?��?;K���i�澈T�<<�<+3K�,�0=�}�<�+>J�>�J#���=8��=�T�=m�z�/D@�����'�=v#�>�,>O�7�a'��g*?����m����=bo��DE��we>uT8>z�ƾ?!]?�~<��w�є��%E�� �P�.Q�??+�?�Փ?�~��OCk�vA?�?i'?S7�>�����f�sjݾV{�mA|��t���=�n�>N�	�p>�K��Wd���ʁ�qT��]��=?N�>S=
?���>��A>\��>y�g��� ����1[�1�U�)�°5���6�׹�������<��\��yZӾ̵[�Bc�>/k��WH�>���>rD>q?n>V��>9,�芈>�-I>��e>��>�X>G_/>�A�=&t�<� �\?iؾ��4��G��[ɾ�2?>��>�_n=W�/�ꭅ�~�9��[�>��?9�?�i�>�wC�Y
R��7N?=;?/�;�LZ?T���������O����˽M <[���9Ҹ>KnX�
dV�R0<��M��8�>�\?�/�=�/߾	{�=�ݝ����=���?�(?��&���U�C	r���V�@�Q�o����q�����ܩ%�?hp�2V��L����؁�L$���l=��'?���?�u��k����I�j�9���y>N��>j�>P�>�G>%���=1���]�q�)�S׍����>ZM{?Ɣ�>��I?8<?iEP?>�L?�>iP�>�h��[��>�a�;��>���>]19?q[-?��/?'R?��+?$Ib>�|�����imؾ��?ɣ?�?G?�?6υ�����Gތ��Q\��x�Z>����=�h�<@ֽ��x���S=�T>6J?�&�m�8�����TRk>�T7?`'�>B��>m��k��Y�<���>�
?oL�>�����kr�,E�n]�>j��?���[=��*>2�=�y�����G �=��¼�ݑ=��>9��F<�w�=P�=���̆�_��:�6�;q��<���>��"?@N�>�H�>�VX���'��s(�`�<��>|�C>\�=w�߾�~������Z�X��#>��?4Y�?G8>���=�_�=�i���Iྖ�
��Ͼ$'	>��#?��A?&�G?�}?�1?�B ?��h=�2�ڔ�	����(j�83"?�",?���>���z�ʾ�憎��3�-�?�U?&9a���2)�3�¾��Խ��>�P/�Z~�����D�����4���w�����?l��?�	A�o�6�Mi�ʸ��7=��C�C?�*�>?a�>��> �)�>�g����H;>w�>c�Q?Q(�>)/?�[?Y�L?G>	0V�V۹��/��w�i���Ҽ�1?�V�?��?aZ�?��>p4�=AH���s{���	���^<D�D�Ⱦ��C>�1B>b�>��>Kr�>�B5>ؘs���o;��x��=_`r>���>�q�>�uv>w�>k�>�
H?��>����N1�4����|�;���bw?���?ʳ)?:�7=����E�${����>���?���?��%?��a���=]匼�g����g�@ù>i׸>�G�>�>�=rfA=�>)��>�=�>T�s�':���\�=�?$-F?�u�=liǿt[]�4l��̏#>�����߽<K�;
���ԃ>k̨������zP�kθ��k��r'��0|���jᗽ�C7?9���0����O>%�ս�B���=9`��1�$=�b�=#����ʠ<�=�����=��E=R��=���F��"=}?ٞz?S?��d?Cϓ>���=���>�?B?+/���L;?ȵ?�y��e��\V�;�T��<f>�l��gx��郾͜��|�H>���<]e>wd�>�_T<'�E� ފ>�K,>��$<l|�=�W�<)>�=�Z>BI�<�)�=`E�=b>J$|?5K������1~�=�n��rG?�Q�>��1=�۾�+_?�e>)�\�ɿ���d|n?@2�?q;?�/C����>�侳� � ��<*�$>x�>4gJ�ǽϾU��>�8�=���\Z���ɽ��?�`@�d'?e��Yrֿ�\
>ڋP>ĉ>\�S��)�{x}�0*����E.?}�<��о_�>Я=���3þSX�<�v$>M�=d�S��[g�P�L=u���C�9<np�=�K�>��D>t\�=`	��+ǹ=��<��>��2>lr����Oڛ�R��<�
>��k>�
;>��>��?�c0?LXd?C�>��n��XϾ�f����>���=��>p��=/3B>�p�>X�7?��D?��K?J��>�E�=�>�"�>8�,���m��E�F槾.�<_��?�Ɔ?���> �J<��A�A��d>��Ž�D?�"1?�x?<�>�U����1Y&���.�%���w�4�|+=�mr�OQU�����Vm�F�㽵�=�p�>���>��>Ty>��9>��N>��>��>K5�<?p�=�猻;��<T ��k��=����l�<wż����@q&�n�+�􏦼��;���;ϧ]<K��;"��=uB�>��K>E0�>��=�iľ���=�ޣ�B6O�.�=쉤�ַ;��fi�_	{�>�(��+�3o>�II>8�N�*+����?a>��>V��?֥^?e��=������;+?��Ĭ���n�<�=]f�=_|N��vE�3�]�CyA��฾���>[�>�Ƣ>/�l>�,�:�>���x=�ᾭH5�F��>V3���M���;,q��@���㟿��h�b�RkD?yK��c��=-~?��I?ҏ?��>S���i�ؾ��0>z:���=���Z�p�b
��=�?9'?�)�>]
쾈�D�#>����H��=�>i���9KT�~o��V��s��vO��j��>p����Ͼb$��8z��5��k%����> �<?�z�?�v���̀�l�i�t龣�G����>n%c?Pk�>Y�	?�?߻u�����n��!���1x?��?t�?".T=�+�=͆��h��>	?���?^��?Zs?�a>��V�>��;�]!>����&�=�
>�2�=؂�=8�?zP
?�^
?<����	� t�_�E�\��;=N��=l��>�i�>5st>2��=x�l=烤=&�[>7 �>��>�^c>��>OP�>�z��Z��>1�X�U��>�i
?��<8��߽#�>Xm+�[�������tED=p2�:&��*˼v:>�p>�2�>_����ů?���<i"$���?���;L��̓=J%�;��=��?q�[>��>)�>�v�>��=SU3>�$�;��ؾ�8>���7��΄D�|R���ξ
�v>�ˡ��|������ �@�4^��o���i�����e>�2=�J�?P�e-i���&�m����?ė�>64?����	#c���>���>�Ռ>%���@s�����q�ྍ�?@{�? �^>�r�>+\?�g?��%��iX��a�+&v��-D���[�ў]�{���	c��V�� ŽDZ?�Cz?�N;?R�<R�U>�ǂ?�H!�{W��)ޒ>�u3��;�S��=�]�>�v���耾N�ھ>#���,���+>�Y?Kw?|�?�B/�� !���k>�-L?�p+?E��?�3?u'*?�Y��6]V?FHH>�2?e):?�Q?���>�, ?�X>�g>�'^�Z1����&���U�������v8=���;�௽���`u=�����3X�,$���<=Cp:4G=�Q=D��<�{�=k9�>��]?-�>u�>v�7?���4
8�5ԭ��x/?|5=C܁��ډ����#4�@ >�j?�ګ?F�Y?}\b>��A�1!C�B>(�>��&>�.]>���>��Z�?����=xp>޵>��=(#O��ɀ�QG	�l���x�<� >�?��7>�F�=_H�>��վ��Ǿ��=E%���ɾFa���`���n����3�>�(3?x�>?��3>xA���]8<c)�M�!?)_?��Q?]C|?=N�=���]4�~k(�%~{�UF>|>Z�4�sv��0瑿��&��!N>�J>�^������TU>O~�Υ�g'��%����%��=� �m�>Ԭ%��O���R^���=��>,g��
��O��h����K?��>���XA��Mg���h>[6r>�l�>�p;<�޼V�B�}Ca��v=�R�>��->d�;r����8�����5�>�D?��n?J�?����ƀ����(�qj���@��Z����?T�>��>(�G>8�>�ڔ���;�M���U����>��>%7�\�@��뎾
� �����>'=�>�[>=k?�/?���>_k?$!.?���>�d�>)�ؽ�\���#?ǆ�?��+>6��Ӛ9�e<C����8�>��>���(0�>Y�?�?��#?��S?C|
?�Ü>*վ_F�I2�>	��>�X�k���v(1>#]?g��>�T?%Nx?�u	>&#�������!��=��y<s!?9�?S�?��>.O�>������>�:0?�(U?�r?{t�?O��>%?>�>��?��;Fti>U�?�@??di?�}{?�1?vf�>wvI=���"<	�v=���\X.���w�l�C<�_���$��� �����"1����V�<�0�:�b��nĝ=g�#=X�>��s>����0>�ž�J��4�@>ߟ��	������W]:���=I��>��?R_�>ø#�Y�=J��>RQ�>����)(?��?�$?��;��b��ھ�EL���>HB?���=Q�l�4~����u�^�g=n�m?��^?�xW�0��V�b?��]?���==��dþ��a���B�O?E�
?�WF�pP�>��~?��q?�u�>�e�3n��	��o;b��j��X�=列>�8�We���>^�7?�9�>Qc>���=��۾��w�Q/���?�ӌ?o�?'�?�;)>O�n�t#��վo���9[?���>�j�\h?�=�۾���T���⾴���DU��ɜ�.޾�[|�����f�p�3>G�?T�R?���?<_{?���5�Y�8�a�����Y�M�+3־&d�.B���9��3B��e������۾�˾��9�es�]9A��N�?:S(?��I����>�ؒ����/t��>�1>�o��˛�u�=�:��d�<#�=T4j�&@6���e ?{�>�R�><ZB?O/Z���>���5���A����p�;>8��>k-�>x��>��d�q?0�̔սXǾJ]��8���>��i?�m?��n?�nȾ�D>�Ę��\�V�^>������]>�i�=R8?Ae�Ɖ]�SN�n�(�5'b�W5��2���6����>��'?��>��>�Ϩ?��)?\�%��&�n!$��+㾊U�=ᇼG�?�"?N�?m��;���EF�>��d?�ʹ>3�q>�h� �)��-9�b�X�%�>�k>��?�O�>Wrk��`�@e�������B��%>vi?l�L��۶���>�m+?L<޽v��;IR_>�i9��K�� ��h����J<?�ޓ>9x>^���CY��� Y�,�|?)?L�?^����)��|> }!?$!�>�֤>,ȃ?�Q�>0��������?7�^?��I?�@?��>�g)=-+��� ɽZ�'�r[%=@ކ>v[>o�z=���=��-\Y��� �̠A=3�=3ͼ|���T��;ֱ���y<���<z�4>�Rۿ)^K�fھ�(�����	�����h���	���������<����x��D�@�%�g�V�*�a�3���Rfl�>�?��?����"���Z���8��������>9ip�vo�:���Dq�b��uP�G��I!�n!P���i��We���J?*f������[��P甾*�W?lL?B�?�.�T��(:n��`�>����0������B噿*ҿ���ܔf?���>�O�,c>{�.?Vy>�E�Ŝ�>:�K�����k𺽯_*?X�a?w�W?e�ȾL��qG¿q���b�?F.@KzA?��(�����U=���>��	?��?> ;1�)K�gް��A�>B9�?���?~aM=1�W��	��xe?��<��F���ۻx7�=��=�=�����J>P�>�p��+A��6ܽy�4>�څ>Ќ"����x^����<Ek]>��ս�&��4Մ?,{\�wf�y�/��T�� U>��T?
+�>U:�=��,?L7H�`}Ͽ�\��*a?�0�?���?.�(? ۿ��ؚ>��ܾ��M?YD6?���>�d&� �t�a��=�5�c�������&V�w��=1��>5�>��,�Ջ�h�O�hI��R��=\?0��H�+�S����<�Hμh4#����&}�=8S�V]Ǿc�t�`�8�;>~�H>=�H>�>Z�>�:>��>?-Q?wT�>�<W���K�r�վ�=�N*�U�>!��$V�=Dih�gҾE��H������'$�|�̾�z�sp�=xb�|b��م۽%��@$g�x�&?�²�Y>@����">9V��zA��x;J<W�� Ҿ�I���j��Ó?lbN?Z�e��tp�����$�8>��$��&K?��Ƚi��w�ƾ�^>u���U�\Fg>�"�=�}
�9��S:�:?(?��#?��ž�#����=������=:b#?*�?��<��>��*?�n#�ǗP�'D
>�A�=#�>K�>)>�踾�4���:?�SN?}�൙�p��>+Ǿ,�V��.$>\�B>/J�᎟�B7�>�ٵ�IN���o�<��C;�q;=gW?���>��)�A��ϙ��m����==C�x?��?Dߟ>�hk?��B?P�<�d���S��5��u=��W?�i?7�>�����Ͼ�Y����5?�e?��N>1Vh�	p���.�3����?��n?)c?�T���<}��������[6?��v?�r^��o��$��&�V��8�>d\�>��>��9��c�>�>?m!#�QH��G����P4�zĞ?�@��?��<<����=�9?�X�>ޫO�Fƾ����z��O�q=�>#���{`v����o],���8?o��?���>D���3����5>�^���ū?��?	��]���W��@��#E��̊����e=����MC���
�z�W���.T
���ؾ�Q�<r��>�@`��<7�>R:+�#���y����?���XDC���0?��>/܋��ܓ�?)F�^AH��lZ�BWH�!վwL�>�>�r��}��v8{�� ;�/���@9�>QJ���>��T��յ�����5<���>'E�>(k�>�~��S��i��?����/ο�������X?5�?�c�?jv?7�C<�)w�|O{������F?qbs?��Y?�W(�o\�~>5��n?���V�P��4�~>���>��0?���>��4��
=��>�r?��>UJ��ȿǯ�������?c��?�� ����>[�?y[4?�,�𘡿�m���Q<���s;��)?/��>.�aD��B�]8���u?\�"?A��D'�[�_?)�a�J�p���-�_�ƽ�ۡ>��0��e\��N�����Xe����@y����?K^�?i�?���� #�d6%?�>e����8Ǿ �<���>�(�>
*N>"H_���u>����:�i	>���?�~�?Tj?���� ����U>�}?�f�> i�?p��=��>��=ڂ���L�;��&>ؿ>�����E?cRN?���>\��<B5Y���4��I��M�$�p^E����>UZ?*�J?`(U>�)���5Ӽ��"��b��K�����<uz!��N����n�K$>U/ >n>>#�xr˾��?\p�7�ؿ�i���o'��54?��>�?#��ϴt�.���;_?Az�>�6��+���%���B�[��?�G�?6�?��׾�S̼�>&�>�I�>9�Խo���G�����7>�B?���D��k�o���>���?	�@�ծ?ai��	?���P��Na~����7���=��7?�0��z>���>��=�nv�ֻ��F�s����>�B�?�{�?��>�l?��o�U�B���1=M�>k?�s?�Jo�n�w�B>v�?+�������K��f?�
@}u@]�^?!9&ֿ���d5��Q?��:g%>�G��d��=�{\�{��2;�d�y=&҈=.��=�>[�=>B`>ʲ=}>S�W>����(�!Ҹ��'��� �2��\E��)���B���P����7��*�Ⱦ�g���]�<�ʽǴ��#w2���@=�/�=}U?>B]?�q?Z��>�νH�>�L�\a[=�[�׺�=��>Q�0?�??�^*?���=���,hY�(^���l�� )����>��->x��>�"�>���>m/=�$(>�>���>V�">ƈ�����V�=K�m>d��>���>���>���>փ�>���)¿�I;�;٦=��M��ڥ?a(���[��¥����B��s�����(?3g�=�����Bڿ�Ȱ�R<D?��:�pm���C[��I
�/�"?�8l?Nv<>��ž4<+�c��=��ལ����t�:z򽏲���^C�I�)�?�We>�,t>��3�ba8�Y�P��1��;�{>�"6?56����7�ڲu��H��ݾ`�M>��>7�E��K��Җ�o�~���h�G�|=y�:?�q?�ױ� Ѱ�lv�Ǟ�C�Q>��\>7P=}�=Q�M>I�_�|�Ž~BH���+=�?�=!^>��?�!D>�=r�>&)���LW��>U6J>?W+>��:?�(?*��Q����}��,��o>�+�>u��>��>ЉH�v՝=��><rL>AS)��P4�[+���5�Q`>ȳ���U��w��d�j=�5m����=���=�*�u6&�y=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ	f�>ur��W����v�u�ۍ#=��> 6H?.I��]P��>�Lv
??Y^�;���	�ȿgzv����>��?{��?�m�<��}@��x�>���?vdY?Pi>�`۾�`Z�	u�>ȯ@?�
R?{�>w8�ŋ'�c�?�ٶ?䭅?���>�U�?o�s?y��>�T����U��D��������>�q̽\ʽ>m�Z>�Rᾘ� �௙�Dd}�;w��,#�Ŭ=�@ =���>��R�����0>v��c?�#���{��>�.v>�΋>z>M�?��G?���>���=�3�}���h��{�K?���?���2n�YM�<ٟ�=l�^��&?�I4?i[�[�Ͼ�ը>�\?f?�[?d�>6��H>��@迿3~�����<��K>4�>�H�>�$���FK>��Ծ�4D�]p�>�ϗ>K����?ھ-��ZH��QB�>�e!?���>�Ү=�Z ?l�#?;�j>j*�>-�E��9��h�E��G�>A�>|�?+�~?NP?c��߇3�,���꡿��[�%}M>�x?��?<�>x'��V���LM�L������Q�?�;g?����?-�?�??�GB?n�e>!C�V�׾����]�>��!?���h�A�
X&�'��9�?Y=?���>ټ����Խ(>ؼZ��-u����?�\?I6&?����'a���¾r+�<�� ��e\��~�;�E���>*u>�a��� �=M>i�=�#m�{A6�=�e<���=���>%��=� 7�V��2=,?U�G�tۃ�'�=}�r�:xD���>�IL>����^?Zl=��{�����x���U��? ��?^k�?7��7�h��$=?�?O	?b"�>K���}޾%�ྫྷPw�!~x��w�Z�>���>��l���D���љ���F��W�Žc,�!��>:J�>Y�?C�>ZN>�r�>r����%����O���]����q99��/���mˡ��]#����#�¾�(y����>���\P�>�T
?Ǫh>-kx>]��>q��>�>�=S>=�{>HҨ>(�V>T+3>r�>�`P<�ϽJKR?�����'���辵���2B?]qd?�/�>��h�S�������?���?Yr�?k4v>�h��,+��m?C@�>����n
?�r:=j��h�<�S��e���I����`��>QS׽�!:��M��mf�+i
?1/?����Ǎ̾~;׽�e����o=�N�?�)?@�)���Q���o���W���R��r��h��6����$�M�p�F�M]��F#��k�(��+*=c|*?(�?Ѕ� ��	���+k�j=?��f>K	�>��>"�>ǿI>��	�V�1���]�s5'��탾�G�>.{?��>@{G?D�;?%A?E@+?��a>�!�>�'2�H��>7��y��>�]�>d�(?��#?	?L8?37?�L�>]R���~G��)�>Կ
?��@?�U%?LP�>X����7=���$x���I8�v�!�%�=�
�=�a��S|��I��=K!>�?�^�8�����Ve>��5?���>g��>����f	}�q�=9��>�t	?�u�>�O��Ws�����t�>I��?��	����<�P.>{��=
����֔���=ʫ��Ϡ�=�{�ʺ.�"�5<ۣ�=ľ�=��ڻ�-�AA+;VN�;��<�s�>��?䔊>�D�>�A��7� ���a�=�Y>5S>><?پ�|��M$����g��Uy>�v�?�y�?+�f=q�=��=�y���T������������<e�?H#?MXT?���?��=?�g#?��>�*��L��]�����3�?�l6?W[�>�|	��ݾP����%��j?�i?��^�����W*���#��5�<�"��pcF�<���}��8�3�O`>r����ê�?A��?L��_����暿8U��q�&?
(?�0�>c�?#�2�zen��D���.>��	?��K?�3�>}mV?Ł?�Y?�=�?K�����z����.>���=�>?��e?5�}?y�m?��>eP$>Z���־1����*�R����X��X�<_�S>7	e>S<�>ϳ�>��=7*`���dH5�m>Ѣ�>�:�>��[>�?7�^>�~y��G?YM�>쨽����JB��(�����2��}u?
�?<�*?��=���'F�q���L��>(�?�?[O+?(SQ�,z�=C�˼r\��7�q���>c�>c
�>uh�=Q�M=��>�D�>��>K7�ga�R�7�
�F���?~�E?a�=�X����n�IK���K��2�=죃�}��m:h�e�3�� &>㥺��<#�S쐾z��K�{�T�|������{��²���8?3��=�&�=z\�=���=�\L�n���:�<&ـ�Td�=���˓�=<"���7��������<�ť8N;����J�{ɾ�}?�WJ?h�+?M�B?��p>1�>2B����>���G7?][>U�N�7��8��ݥ��#����־  ھ�a�J���9�>"wO��>o�+>^��=��<�e�=�ns=�;�=	�7��=Fn�=�=�=�=�y�=>��>�6w?U��� ����4Q�7Z置�:?�8�>1{�=��ƾc@?��>>�2������kb��-?���?�T�?E�?-ti��d�>^���㎽Kr�=ⷜ��=2>���=>�2�(��>��J>����J��d����4�?��@��??�ዿŢϿ/a/>!�7>�N>��R�,�1��Y�!�`�p \�B�!?sj;��ʾ`�>��=��޾Cƾ%�-=��5>b�_=�p�%,\���=��t�}�6=4Cb=��>� E>F��=�����ù=$kN=pT�='Q>VB����8��K+�75=gt�=Ukb>'�%>{��>q�?�@7?�{b?���>�.��8Q��ɰ���l>z��=�a�>��=�<><	�>��9?�??sT?i��>'Í� ��>R��>	m-��`k�bپ����SO=�h�?�`|?�#�>MR�<<I�&e�q0�Hܽ�?R[-?�$?�Ǧ>G���|ؿwY�Y�,�����ؽ�à���J����<������(�Ծh/l��I�>�z?��>k��>�~�>�>��>m�S>�^=Q�j=������;Ք�<E��<��J><pU>1J���[�lo�=�f>�ò=�D�=�q�=���<�����=��>4<>���>Î�=����C/>������L����=�G��;,B�{4d��I~�N/��V6��B>�:X>c}��74����?��Y>-m?>���?PAu?$�>� �6�վ�Q���Ce��US�jʸ=��><�<��z;��Z`�a�M��|Ҿ�E�>���>9{>(_>��4�kB�fd�=�撾	M+��h7>�����=�f�=ѝ���������������j�X?����"y$>'c#?��Q?�X?���>澔�N�����>��~���_>! 3��c��6�^=ؑ.?z�)?=�?������6S̾�A���ҷ>KEI���O�����f�0�*���շ� ��>!�����о@#3�Tf������ŋB��Lr�J�>_�O?D�?J<b�iW���UO�����#���o?�zg?��>�K?F;?�A���~�@n�����=��n?&��?�;�?�>���=���@��>Oc?���?Rp�?4�x??nU��H�>�(��^l>�����{=��>���=�s`>~&-?�l?���>�K<��-�[	����	<�1�=2J>w�e>��=-61>�k����=�xD>��V>�%�>��>�	J>���>��>����I��}?��=�)>Qt?+��>�[=9�$�H7z�oN�9!,�ټٽ�ڽ�I���y������8=t<=�X�>E]ɿ^��?<@�>S1�	?�ྷ"$���M>��G>�m�[~�>��>��r>�3�>�T�>�<<>�$<>�y$>x���@> ��I(�4�h2��	꾮׉>�c�U�<��<ٙ��s9�x��-���x�Y�єs�	YE�L���W^�?��h��{�t�E�m
<�0?���>Ct;?b����<��">Ui�>= X>���l���� �����S�?�1�?��c>՝�>��W?s�?��0���2��Z��Ju���@���d�+q`�nꍿD�����
��ͽ�
�_?y?��A?���<�3z>ь�?��%�������>I//�u:;��==�$�>TY��¼`�F�ӾPľ%��,F>�~o?&#�?=E?hV�b����D>>�C?�<5?5�k?�%?��A?��۽�s?42B>�?�4�>�7)?U2?H�?u�A>+=>w =2&�߶��#`���湽����x�b�Y<d��<��D�~p=��n;7��������MYY�zĽ�A&�8��=q�~=)�=rڧ>X]?�W�>���>0R3?�z.��b1�r����+?��!=��l��v~�*���F��>��h?Mv�?[�W?�J>^�:���@���>��>�9>�Q>�J�>ݸŽSC�Q�o=�
>[�>B9�=K�!����v�
��2��v��<pv">3��></|>9
���'>_{���/z���d>��Q��˺���S��G���1���v��Y�>��K?@�?ݟ�=�^��.���Hf��/)?$]<?%NM?��?7�=?�۾��9���J��=�N�>�Y�<��������#����:���:R�s>02��N���\b>?L���྄�m�M�H��hH]=���d=����Ӿ����t�=�V
>~��� �+�Nߪ��)J?_Dn=����aW�������>:Y�>f��>,K�b���L@��;��3��=�$�>�!;>4����QsH�Vk��n�>��A?�`?~P�?������,R�3���f��DRͽ	�?m.�>8��>�I7>���;+���-,���c��G�6�>[5�>
���9H�X����㾊�&�b��>�U ?!m">E�?�J?k?��e?�(?��?��>4뽧Ҿ�"?��?=��==_����W�l28�W'>�4��>�D'?��.����>�	?Oe?�;(?C�N?�?�+>�P���w;�p֒>�>��W��0��aU>��K?}�>�
[?V�?p,>�[2�����C��/4=v@><1+?Gt0?L?i�>��	?s$��DT�@�?��e?!�Z?�w?6�>� 4?]zX> V?�P2>b��>�?G�'?��(?#o?Nyb?|`>�a���U��9�;m�d�<����;}�=pη��)��B���ʙ��Iٽ�-z�]/Z=[&�=�K����=�<�_�>z�s>.	���0>��ľ�M��(�@>>���,M���׊�-�:�b�=ˇ�>X�??��>�T#����=��>�H�>l���5(?a�?�?� ;��b�o�ھ��K�h�>�B?3��=��l������u�	�g=��m?	�^?	�W�t"����b?h�]?�c��=���þW�b�,����O?F�
?<�G�W�>��~?��q?2��>jf��7n����Db�{�j��ζ=�q�>V���d��<�>w�7?�L�>��b>�#�=)r۾]�w��q���?��?��?e��?�/*>��n��3���������� _?�\�>D��i� ?7��;�׾!U���m��c�f��&���m��������a�ba����ڽ-��=�'?�2p?�br?�bb?������b�@�]�������Q���?�[�A��A��:=�*(m��N�`�����{:=j�`�J�:�?�*?v
��+��>=�w�v��"�;�2>�������@�=��ν���; �=xcm�NS1�װ���N ?�w�>���>�zG?�<S�b�;��<2��?�{��t��=�a�>߆�>/��>IkW=�@;�$ܠ��p۾�Eo�P\ܽ.9�>��W?��\?=d? ���`BF��N���9*��MI�?]̾��q>�b>���>�ը��]�Zp��i>��p�� �ᙾa����> >�?�e>�$�> *�?�?��i��������2�&�o>���>�`�?$�>"϶>.ə�Om��-�>��l?���>��>�I���t"�hWz�Tbս5�>>x�>JD ?��i>�47�j�\�V����u���#9�v��=�i?_���l�g��9�>/�Q?�|�:Z^<�ϟ>}O��" �꾐�&�jm>D�?tj�=G�9>�"þDg
��z�mǇ��P)?�e?E[����'�Q��>m�!?���>�>ީ�?>�F��ɏ;?d<^?h`I?S�??�A�>�=7=�鶽��ǽTa'�<�(=b�>�_>�=}=��=dJ��[�� �Q�G=X�=%��G���
<:�ȼ�#<L�=Z
4>�ܿ��Y�!��E�N�þ�������)�K����ؼ��%��1���]J��_���57��i�b��
U�y���x��_�?5�?\��p��԰���w�¨����>)%��;�<�;��B�i��q��w�.R���%�x�V��@t�s�l��5?[��_
˿eV��A� �8�4?1g)?��?���2���E�'��=Y	M�bS��0Lݾ����<п�S�>�G?�B�>�:ľ�*��7�?R�'>��Q=>h�>I��lq� �\�O�?�[�>�+?u����bڿ��Ϳ�\�<���?�6@c|A?��(����%�V=���>�	?��?>?>1�`;�A�^�>":�?���?c�M=��W�C�	��e?Z�<9�F�d=޻�=4�=H#=���{J>\T�>���RrA��Bܽڲ4>Cׅ>ȃ"�S��u^��(�<|m]>i�ս�(��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=`��yUٿ�n7��G�&>�k�=f�#��p����\�A� <2�	��諭/�H�� 5>S�`>�9>�w�>+�>��}>5&f?��d?)�o>'��=��=x�m��󾮬$>��&�;���;���S:�(��|�þ�]־'����.�Ya@�9��Z<'�s��;Uqt�쩥���Q��aʾ�Ё�j�S?`�u=&Ʉ>�ǈ�I��>iݾ��ɾ2ư=d�=\5��¸$���{��5�?ƗX?��J�//���1�u~<ԁ���I?�e���k޾��_�%d>lS����ѝ)>�L�>B����%��91�Ot0?�4?�s��4 ��S�*>�w ���=��+?��?�)\<a\�>�G%?0�*��P�]�[>��3>X�>���>F�>C���S۽Ry?�ZT?���Y7��M��>�h���:{��`=-(>�F5������[>`d�<�����r]��0��,U�<`(W?���>A�)�A�5[��^��Cw==l�x?<�?�.�>O{k?��B?"��<ue��c�S� ���w=\�W?�'i?��>@����о􀧾6�5?4�e?��N>s^h���龌�.��S��#?"�n?.]?c���u}�L��n���n6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?p�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������m>H񥾑(�?�<�?4" �J�����Q��C/�r���ٵ=�w<�]���c��O��L�����@Q��-f�=���>8�@0t� b�>`C��
�s�ݿx�s�(󝾠QžX� ?��>�>�d�M���j���a�F�_�G:��ͬ��.�>��>����e5���{�uF;�����.�>� ��l�>�&T�x絾1���Թ2<t�>��>���>}3���������?[$��(2ο;������ݯX?�]�?h�?�U?9<<(�v�!{������F??js?A0Z?��%���\�:�7���j?����E`�>�4�6UE�ͥT>,3?�2�>�-� �z=>�>\�> I/���Ŀ�㶿���ަ?���?���+��>ϐ�?�+?
a�{;������w�*��˃��A?z3>���l�!�4=�ߒ��
?Qj0?Dv�=%�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?$�>��?�r�=b�>mc�=�񰾰�,��j#>1$�= �>��?��M?gL�>�Y�=%�8�%/�[F��GR�u$��C�2�>g�a?��L?�Kb>���G2��!�%vͽ�b1�P鼧V@���,�&�߽�'5>b�=>/>��D�Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�P��=��7?�0�.�z>���>��=�nv�޻��V�s����>�B�?�{�?��>"�l?��o�M�B�q�1=0M�>͜k?�s?aQo���j�B>��?������L��f?�
@}u@_�^?)�Կ�螿{[��밦�K��=:'=��>��&��a�=�<��[��½�9*>�W�>��n>�*�>eW`>B��>U�=<��'��ŭ�O�����D�W������<������r��Y��
־�,��o�7��ʽR�#��'�d����=��J?�i?(`?��>reO�`'>ف߾�r�=�G߽"�=��>� N?�lT?�f4?�h>�����)P��D������81��ĭ>�.>�?�>H3�>���> e/��Ox>�h>�T$>��;>M�۽�rG;<��=�;4>��>1?�>%�>ң�>��k>�l��.�ƿK�R��;Ѽ�)��W�?���<%-�Yw��+MJ��G�o@���-?���>]%����~���m�@?�vདྷc�ܗc��jڽ7.?1�{?r,%>�=¾����N�> 4��7`о˻�>,۽n\ʾ��K�m��M�"?��f>u>̛3�ve8�Q�P��|��j|>�36?�鶾�D9���u���H��cݾ~GM>�ľ>�D�l�i�����#vi��{=Px:?̈́?�6���ⰾg�u��C���PR>�:\>cU=�j�=bXM>@bc�	�ƽMH�/h.=���=�^>�H?��(>�p�=Q�>�U����K�7<�>��@>Y�1>��>?^�%?�s�H����{�dF%�*z>Es�>�C�>o>�JI����=��>_�\>B�Uě�A&���G�eU>)����j`���~�9��=��	+�=��='G��U8�bN<=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿh�>Ix�oZ��~����u�D�#=0��>�8H?�V��5�O��>��v
?�?_�ߩ����ȿ&|v����>R�?���?��m�lA���@���>2��?�gY?oi>�g۾]_Z�J��>λ@?�R?��>�9�r�'���?�޶?¯�?]>���?�p?ձ�>T���/P�P���A����=���ԥ�>�Yr>�%پ��<�a����8|���p�d���{2>l%=�θ>�꘽�Ͼu�]=�읽�nҾ_�!<L��>�4i>-�q>>'�>�X	?���>��>�)�=r,0�霾�vϾV�K?���?����2n�.G�<���=N�^��&?mI4?�i[�(�Ͼ�ը>6�\?m?�[?'d�>��?>��>迿W~��
��<��K>�3�>!I�>�#��hHK>m�Ծq3D��p�>gϗ>����?ھ -��="��DB�>�e!?���>�Ү=Oj ?�"?[o>�g�>EF���� G�≯>l�>��?�}?-�?ް����2�C���/<��~�\���J>qx?8�?[)�>���.=��满*y��>���Y�?�Uf?��ｨ1?$��?`=?A?��`>C���1ؾ�κ�D�s>��!?U�)�A��M&����~?�P?:��>�5����սiBּh��.����?�(\?[A&?����+a���¾�9�<�"���U�h��;�D���>]�>G�����=">2ְ=`Om�AF6���f<Bj�=���>a�=E.7�)u��0=,?��G�}ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?`��@�h��$=?�?S	?n"�>�J���}޾6�྾Pw�~x��w�Y�>���>'�l���K���ڙ���F��]�Žs�i�K?�\�>���>Ca�>8?�����>Cn��0�:�9�8��g�T�w��VE�u�`��(I��<b��پ�]��٠ >c/Ҿ�����>|=!�> ��>w>f[�=���>vf2>_Pl>E��>�$>+�> �b>���='�>���=�>8�9KR?"�����'�F��(���A6B?�td?2�>5�h��������<�?؄�?(r�?KEv>|h��'+�?n?5:�>���vn
?Oj:=���ܕ�<�`������^�����\��>�A׽f:��M�wYf�Qi
?o3?zz��W�̾�$׽����=�3�?�U(?|@*���U��o�om[���Q��k��4W�������'�-Dp�됿���.O����%���i=$(?3 �?�+ �����T���j�T�B��_>̽�>;��>.��>g�`>�2�C�-�	�[���!�⏁����>j�s?���>�Q?G?�A?ͥ??3~>Yԭ>�J��e�?��_=3��>�f�>_7??>?�Z$?�<?�h>?`��>���;��۾l�о��>��?";?�#?A?�>�Ѯ�0FG=Aؓ<t֌=Vb��v�Z�^-=�n/��z(��[���Sg<v��>;Y?��v�8�v����k>G�7?���>���><���&�����<��>n�
?hI�>����Jzr��\��Y�>���?	�:u=w�)>D��=ϔ�� �Ӻ�Z�=v������=D^���w;��g<�x�={�=��s�κa�f��:��;���<�t�>D�?ߓ�>�C�>v@��#� �>��%f�=&Y>@S>�>Fپ�}���$��O�g��]y>�w�?�z�?�f=��=p��=(}��MU��^��������<��?MJ#?XT?W��?G�=?Mj#?��>+�`M���^�����ɮ?T�8?h4�>����
�� ����!���?X� ?������&��-�����I���e�~Ɠ�����GHJ�c�>�:�oˏ�]��?x�? ����
q�x�ѡ��`�>�?	*?��<)?�;Y��!����.����=�q�>��Z?a~�>�iG?�)�?lN?R�<��N�N���0ˌ��������=qs5?��?���?"�?�L�>>NG>OTH����1�����ܟ�yG)�mCA��uT>{�>��?|��>y �=��=�B��-��?O>BVZ>ؿ?���>e?ӄ>��<��G?��>�达_��ä�����9T<���u?���?�+?�q=�_���E�!���[�>�U�?c��?OA*?�}S�y��=6�ռ8����q��V�>&�>�$�>��=r�I=�H>���>X��>'����_8�=AM�a�?�F?��=��ſ��q���p��ɗ��=c<1��e��蔽2[�n̤="�P��ʩ���[�6������ �[�����{���>ؖ�=���=���=�)�<�wɼ�|�<�J=��<	�=kAp�x�n<��8�`�ϻc�S���[<��I=>��A�˾��}?�<I?o�+?�C?d�y>D2>��3����>�v��b@?9�U>�4P���f};���������ؾM`׾�c�Ο�|.>��H���>@O3>��=���<5�==s=8�=y�J��=�p�=�<�=D�=���=��>L>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>k@7>�5>A�R��1�/�[���a�Ď[��!?�(;��˾Ǉ�>2��=?߾o�ƾ%!/=��6>��b=l��F\���=��x�M�:=Of=i��>�C>1ƺ=Uo����=d3I=4�=(rP>Y����b<��$.�Ri:=�p�=5�b>U�%>��>;�?�)F?��X?�X�>Le���|���]�>�>�۬>]��=��x>���>�
3?	6=?��S?�۴>��[=M/�>���>��3�Dnc���Ҿۛ]�O�p=mq�?�Ä?jљ>�aw�,���I��cS���ɽ���>�N?��?� �>���쿱�+�V�'�����r0=������q��P�y<�U��X��z==��>�7�>nh�>�N�>�6�>�|�>!��>�G�=�퀽�I:t�=>"��;�D>*�E���<�i\��b�<@�>���=��<C���e`=&�ӼW�>��=}��>27>���>�t�=���F/>������L�#{�=4;���1B�l6d��L~��/��q6��B>+1X>&`���3����?��Y>lw?>��?�;u?R�>E�߱վP�� ;e�]BS�;��=)�>��<��x;��N`���M�	Ҿi9�>�ξ>5�>�>�>�m�F��~b=]�꾮�Z�`L>{
��h����n������p��B����������gY?�������=�Lf?�7]?/��?'L�>����MҾV�>ƭ��}�x>;���rϾ��J��h3?��?Ӥ?������T��Ͼ+�l,�>��>��2P��q���$,���E�ھ��>����ʾ$o9�C7��˂��'�K�<{�Dw�>�T?G��?���ITs�t@�_�.���?_�Z?�)�>!�?[��>޳f�(Ѿ.�t���=�w?^"�?�u�?7 >��> <�	��>g?҄�?]�?TS?^!%�҅?q#�=@�>����uC>c>�[�=U)�=u�?zf?��?R������*�m'��d����<�\>ɕ>��Z>D�>�!>�H->/��=�ڢ> �>�x>�/,>��>A>&��o��=�?i[>zF4=�{?̼�>���3:-�BvQ=�w�<��;�1���΅�4�p�;�ݽk}d��q5<8>wy�>g#пf��?G�><y.��+)?���D���Px>|P>�w����>�4�>���>���>��?=�.>>>�'�=�_Ӿ�<>���\v!��B��ZR��Ҿ��z>N���9%����(����wI��Q���I�jj�� ��w@=���<�K�?����k��*���y�?�?�>6?Aь����>~�>�Ӎ>����؃��d���:��?���?�;c>��>Z�W?�?��1�93��uZ��u�1(A�e�0�`�y፿��
�����_?"�x?:yA?~T�<:z>>��?�%�Aӏ�*�>�/�';�y><=�+�>*���`���Ӿy�þ�8��HF>W�o?,%�?xY?kSV�L�e���A>s�2?��1?3+c?�^?��0?��/��s6?1p2>\�?G�?9�>?=.?r�?z|h>��->�At=O}*= �a�o�9&�����SN=���=��>=(�ۼ�s�HA�=�*c=o�<�R�B�=�F������=��=cz�=ZΣ>YS_?0�>�>!�5?	��n�,��)��f�5?��z=�Sr�&���G��Nh�d�
>��a?�k�?��Z?�Ã>#;�.PK��v�=�*�>ٵk>��>(�>����.�?�=f�(>���=˔�=3�4��߈���	��*����6;� 7>���>�2|>���&�'>.|��~0z�n�d>��Q��ʺ���S�	�G���1�؂v� Y�>�K?k�?|��=\]龬(���Hf��/)?�\<?�NM?2�?��=��۾��9���J��=���>�6�<o�������#����:�C$�:D�s>>0�� S�b�>R�)�^y6���QV��*/#��i>��޾*Ȍ>� G�n�ƾ��e���<ըK>m�վ�W'�^v��ͷ���H?U]w>���(������9>�EQ>C|�>iNX�����K��˿���׽� �>WAE>������ھ�)4�Q��K�a>�;?v�z?�]�?���V	��R��G�������k�=1�?�>��:?B�N>9�h>�<I�ؾ�Y��,a�``�>}�>u�'���9��ԃ��ﾒB��(�5>݆�>���=�"?��_?]�?�ua?q�O?�v�>�E�>��b=�8�(�?���?x�>�b���Ӿ�&�O��|�>�?�Ρ;�A�>�o�>��2?u�?�Ym?Ё2?R�>i\���9W�a^�>D��>f~k����h?�=y$�?���>A�+?�?�W�=��"�sB��@��%�>�oǼ�X�>��C?��@?�]�>T�>�������H?D�B?H�?6A�?Zx�>C\�>`s���A?�1!>�/�>B8?��#?�A6?��?�%?�B�>a��Ow����y��l��T��=I��<��F�l�
�<���=�Ʊ���d=�}G�oh��6o�;�y�<�<=ؑI<��=�_�>��s>Y��w�0>.�ľ9H����@>1G��2E��QҊ�4y:��շ=���>� ?���>'Y#�#ɒ=D��>�G�>R��M/(?��?L?$&;u�b��ھv�K���>t	B?���=��l�A���!�u�*h=h�m?ֈ^?h�W��"����b?F�]?xj�=�b�þۦb�Í���O?�
?t�G�]�>��~?��q?Y��>j�e��9n����*Db��j�ض=s�>xW��d�:�>��7?�L�>��b>w�=u۾x�w��o���?��?^ �?I��?�(*>z�n��3࿣뾜P��ϲ_?5�>!/ƾ��?�i�<�P�F,a�캡�p�׾�{���ԭ�h���d����i3��>���߽�*�=��?��h?K n?.]^?�g�c���i���}��cM�������<�?�D�$�4��ja�cV	�k�%�����;o�l�I|B�|��?�y,?�0p�Z�>6��0������>�d��my�M�u=0�ĽoX<zd�<r��.�n~��E#?OI�>��>�=?=Z��&>�
=�i�8���|�=��>�z�>�>�<�<,��wAͽ�sžN��,\��=�>N�=?��?�`?���b�Y����;�)>,>t`^�Ya�>rĥ>ɸ�>�m���j(���Ⱦ�� ��v���پSeѾ����-�d>�\3?T3�=���>Q��?�d?�K?�7M>T|�@�]����>�̹>r>`?K):?�Z�>�kս�7ξ\�>��k?�#�>SI�>
)��^r$�p+~�AU뽧��>���>���>@8�>�@.�VM[��%��|ʍ��H8����=�xa?�х��h���>ȟQ?tTX�8�J<� �>b���$��hݾ��"�[�>_?�3�=SH>a���j�	�h�z���~�9�'?��?QS���q(�_)->�[*?\��>��>���?��>+e����k��2?E�c?��G?��6?7��>���=a��'�����F	n=j<{>�>[^�=n�>��4��76"���=��==��p\����Y���ؽb��q��;g>�^ۿ�:K�u�پ�v��W
�8��u��~���>������왾��w�����&���U��c�縌��m��p�?Y,�?6������������۲��	l�>0r�Y���������ޕ�B�ྶ���U!�X�O��!i�v�e�/l6?z(ʽ�쾿O���R�׾�)?��?!�?��,�A���Y���>�'Y��-��n��'���տH��M?n!�>8-Ҿ�Nu<��?��?>�LD<im�>���~�������B?T]"??�?�꺾�߿�t˿Qo�߫�?Qq@1zA?j�(����ehV=E��>��	?��?><11�C��
���Y�><�?���?��M=��W�c4	���e?�<1�F�I!޻��=�k�=�H=g����J>�P�>�Z�f`A��sܽ}�4>�υ>�l"�܇���^�a?�<�]>hֽ8r��5Մ?,{\��f���/��T��U>��T?�*�>U:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=r6�щ��{���&V�|��=[��>d�>Â,������O��I��V��=	���G���n\�C-.��g�>>@0���+�=>�l�M�>������*��<Y�>D	|>8�t>r��>i9> ��>	�V?�\k?{��>�����>H�<Y������>�ʓ��>!�����w��=XX����=�� ��ݗ.��8�z�*� ��=��T�������;6�%��*T��.%?��>����V�a���<F"������t�<������߾:>�R�c��K�?�VM?���ԜW��}	�g��<�����D?N֥�� վ)ž�!�;׮���=��>�|�<��&}%�|NF��0?4�?>������#>��T�!=f�*?W�?a�<��>�"?�$���ͽM]>�/>f�>S�>/	>�����཈L?�T?�V�Wd���"�>����/w���i=��>��2�i��H&b>w4S<$��F�Ƽ������<�W?�B�>��)��yߐ����y�>=jbx?p�?>6�>�jk?�B?���<Đ��C{S���
�,�}=S�W?1�h?�9>�ွ��Ͼ�}����5?��e?'rO>��g������.�pE�$�?��n?��?����@�}��
�������6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������0>j%���i�?=�?X^ ��(��
�*���i^���E%��Ԝ=ڬ�<߮����ͷ>���׾����O��}�c�QL�>è@��½�'�>"�u��NῸa���a�<��n��a2?�2�>�ǝ������Q���k���G��?��$��i�>�e>R����d���){�f;��x��"��>��	�T�>S�Q�C����ޝ���Q<,�>��>ȭ�>��������Lm�?�"���FοVj��:x��UX?�5�?�q�?W�?]�<�Zw�1�~���G?n[s?��Y?Q@$��[�(:��)j?�_���hZ�~3���B�OO+>Y�/?���>�7��c-=f6>���>�J�=�q9���ɿN���	�
���?z�?�g��"�>ȃ�?,5?���왿p;��it3��om��i;?F�p>�־&?�`	:�h����
?N/?5�	�ZK!�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>cH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?u4�>�?���=b]�>�	�=��	3�:#>��=��@�U�?-�M??5�>���=p9�4 /��VF�3FR�Y+�+�C�'��>n�a?΁L?�b>l��5�1��!��νY�0���"@�\�*���߽�]5>�>>U>E���Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*�z׿?���"�ƾwٜ�;�=?�><+�=Q����1��+�	ے�Y=̼3�=�>@��>��|>��>nk>7�>l���G�(����ꋿ��<��\(���$��Ȩ����!T���D��n�;��"�F<hv3�j<�ȣL���%�D_Z�N �=�vU?(�R?�*p?t�>����MZ >�����=��!����=j��>�#3?�ZL?��*?�f�=؜���d�����}⦾�ˆ�$��>GH>u�>��>�	�>8;F��F>z>>>��>"�>G�+=� �9V�=� O>�5�>W=�>RƸ>j�> ��>[ʰ�]Uƿ�z'���-=��m��?��������ʵ�(�a���g�ѽ?ѕ�=-(��	ݿ~׾�)B2?P�l�3־LP��R�`��^�>>�v?[��>������>��=�������w��
��*H�g=W�?,�f>tau>W�3���8�bsP������R{>�76?�׶�q8�W�u���H�>ݾ=�L>u��>�H��g�e�������h�aD}=�c:?�N?�>��Ѱ�[�u���d�Q>��[><=�2�=�M>�f�w�ǽ4�G��-=gD�=8�]>�8?Xj0>��=���>����-J��|�>j�A>Y�2>�y??�B%?y��� ���R��W*��;u>�@�>]r�>�>�EK�1�=E��>_c>�ռ�c��G�	�=���X>��x�Uh^�� r��u=����7��=���=����y?�U�,=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾNh�>yx��Z�������u�z�#=T��>�8H?�V����O�c>��v
?�?�^�੤���ȿ5|v����>X�?���?i�m��A���@����>:��?�gY?moi>�g۾>`Z����>һ@?�R?�>�9�}�'���?�޶?֯�?�K�>懆?��y?b��>��;iS����^������>2�Ͼ���>�>\����C�7��������N`��J�}U���=�x�>82���mѾx�;>3籽cѨ��˼*��>��>�\:>��>��;?�v�>ޟ�>g�=�F=���W����K?���?7��8n���<�ߜ=}�^��(?qF4?^jZ���Ͼ"Ψ>Q�\?���?�[?�^�>&���>���翿�w��y��<��K>�*�>�=�>�D��#JK>;�Ծ�LD�fh�> ��>����Dھd4������F�>a!?��>ȣ�=� ?0#?%�n>f(�>��E�9]���F��n�>��>��?�~?�U?���\�3������ܡ���[�)�J>j6w?�?gk�>�县xŝ��I��b�B��Ă?Fg?�I?�$�?�<?qF@?Bc>���׾Z����|{>��!?�<�R�A���&��X��'	?ь?(�>� ��l�ѽ������V����?D\?��%?2��x1a��Hþ���<�c��ld�g��;I�c��>>q>Pׄ���=r�>f��=��l��6�PfX<�0�= Œ>�2�=^T8��N��0=,?��G�~ۃ���=��r�>xD���>�IL>����^?jl=��{�����x��	U� �? ��?Zk�?a��@�h��$=?�?S	?n"�>�J���}޾5�྽Pw�~x��w�Y�>���>��l���K���ڙ���F��[�Ž��3�U�?��>��?���>�A�=|@�>Br���4��J�%���J�/D8�J@Q���J� �'��������=x־����ֈ>7�I=� �>�?(%�>X�=���>]�=�N>	�d>��>.�>-o�>m_>�v�>b�n>�KV<?KR?8����'�������:3B?Wrd?L2�>4i�����w��D~?酒?s�??v>�}h��*+��o?6>�>C��>o
?�!:=�Z�;�<�T��@��K5��2�����>D>׽�:�UM��pf��i
?�.?������̾�9׽�v�(�v=�a�?)�+?��5�m%Y��v��?b���1�f�<�3�E�\�K��\@��Bn�G��5*���\����%��o<�a'?%/�?�N����	��]O��t�i`�Tړ>e��>q�N>+�>(�>3R��,��T���)�谇����>��Y?��>,&[?��=?oL+?�M"?�>�m�>'_�!t)?#>�T�>eτ>�,9?X?R?a�$?���>�+?�ƚ>D������
��;7?DI?n�??t߅>1�?8�i=(�F��=��Ż���lK�,4�����J=tr���W�t(>JV?����8�0#���Zk>��7?���>���>�ڏ�������<���>��
?��>|��{_r������>ߏ�?4���=|�(>X��=#ҁ�W�
��k�=!cȼj�=7o�~�8�WA/<��=�)�="3Z����99t;>�;�<%[�>]�?���>�H�>T.���� �����=�Y>�!S>(>�Oپ�z���!��W�g��y>�o�?�u�?Bg=��=���=�r��&C�����彾G#�<!�?�J#?�TT?���?&�=?`m#?��>�)��F��$_��� ��v�?��4?Yη>����~㾮Z���+���?3`?�p�T5��/,�l.���#��)��~W�����fķ�Xy5��FE>$��ݣ�o��?톧?�2���hX����fۥ�ģ����#?Sx?�&'>�r?�);�=����-��/>�?��O?�-�>q_O?*2|?��[?4�M>6�9��䬿嶘���4���#>��??-B�?xH�?�w?���>7�#>:''���o���]!����임���N=��X>XU�>�L�>t�>�'�=L�ƽ�Q���9����=6vg>*�>U��>���>o=z>�Ł<��G?��>c-���i�����`6���M7�+6t?���?d+?0y =e��pD��6�����>��?Q!�?D�*?�)U�^�=y̷�����zv�{��>���>���>^-�=J	r=T�>>
�>µ�>Z�����[9�^�l��?��E?�X�=����V�]�`3����Ⱦ�(8>u��O��'^�;���h�=��ƾ<�=Z.�����n⮾8w��b��SK��8���	�?x�>�>qx�;�>�=��<��q�D�i[&=lI~=��GK�=�T��1�����E�D@%�r���>?�$SR=cs˾�s|?��G?��*?�C?�St>(>�vd���>�S���?_dB>M��֚ž�Q����ΐ��Ͼ5�˾��c�Mͥ���>M�-�'o>� A>:�>� 0�8�=]�=�7�=�����8k=s��=K�=�3�=�7�=v�%>$�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>F)>��=�eQ�3�K�B��5P�8�f�7�!?��;�EZƾ/�w>���=��Ҿ�ɾS�=��5>��^=��#��/\����=b�C�{v^=B6==)��>j:F>J�=��ǽ�k�=��L=A��=\Y>�~����r�ڗ8��|!=_"�=��Q>7�+>d(�>-�?�/4?��b?|�>NB����þi��(u>d� >���>h��=�f>,��>�??v�L?#\H?7��>�Gn<���>��>�$2�_�s���꾃X��u�<��?ӧ�?��>�\�<z�,�!J!��7��<���.?Q�3?�?�W�>����A���5�����ŽCF��z�*�j���p�<�-�@%�|�8>�l	?���>�j�>��j>>݆>/�>8��>B>�$����=f�s��=�����c�>��=�U�=�Ǻ�O�=p��=4-�<aG&=nL�5R�=k|���U�<���=7��>�@>S��>7��=����C/>R���Y�L�L��=�D���+B�]5d�AJ~��/��Y6�)�B>�3X>�|��4��a�?��Y>�q?>��?�@u??�>����վMP���De��PS��ɸ=λ>��<�Qx;�ST`�N�M�\zҾ�>���>�i�>eC;>�?��E���X=a��t�M����>�Q���C� 퍾hz��Ep������%(��Gլ�ݣ@?u����V=t}?��\?/6h?T��>��н�<Ѿ/ٶ>2�g�,�`>�	�j-�� �==R�9?�G?�$? m��Cr_�9H̾ ��A߷>�>I�5�O�R�c�0�F��̷�e��>����f�о�$3��g�������B��Mr���>.�O?/�?<=b�CW��*TO���� '���q?�{g?��>;J?b@?J#��-y��q���x�=��n?n��?�<�?�>�+�=<��%>?�?3{�?/�}?�(�?��ʽ�˜>Z���y>y_G��Qs>�Օ>��=�L�=�%?��?2n?��%<���� 8�����/r����x=���=f�>�o#>��;��Wڻ	Q�%_���>�B�>��Y>�\�=h�>GN�>}���.���&?w�V>JP=Y6?�.�>KG��-a=:���{=ȧ���p�qx��s�� 
�DO��WX�=jmA>�<�>s�ѿ��?�P�>�M�z`�>�)־��Z��h�>�/:"��l��>Q,\> P>T��>[��>5$=<�=�c >EBӾ��>��Aj!��C�atR���Ѿ�{z>������%�ѥ��g���<I��o��3b�;	j�l-��~>=��t�<CG�?tr��Z�k��)������?U�>p6?
Ό��鈽��>��>̹�>�<�������ƍ��fᾶ�?���?�;c>��>R�W?,�?W�1�33��uZ�+�u�G(A�&e�7�`��፿�����
�����_?��x?yA?�S�<H:z>F��?��%�Aӏ��)�>�/�.';�@<=]+�>K*��d�`�y�Ӿ��þp7�!IF>�o?.%�?`Y?�TV��oi�%}%>��:?m�1?Bt?jz1?�;?���:3$?fk3>��?٬?q5?�/?'�
?:2>��=����m-=����������ؽNν����4�2=աy=T�K;��<r�=�p�< ��9��;�g��<�i4=��=,�=Hg�>�T`?4p�>L�>Ft0?�W�f�3��}��v3?~O=G�v��퐾`x����侩�
>�Jg?�>�?�\?f>#E���>�*<>��>�L;>(ra>�P�>�ݽ.�.�k\�=J�>uM>֠=�	ڼ�3��y�8Y��"Ċ<�	->���>2|>�����'>�{���.z��d>e�Q��ʺ���S���G���1���v��Z�>��K?M�?N��=^��,��If�8/)?&^<?POM?��?q
�=��۾
�9���J��<���>Qe�<�������#����:��z�:.�s>�1������P:>��
�����X�m�>�����Kf�=���_o�=����龘������=�>�Tž���x\������ɡM?���=�����Hk��ν��>��>���>T���̻�<A�eT��{ y=��>�F>��$�,���יH�o=����>�vD?,G^?"�?�Č�rcv�G��B	�"̅� 9R�>D?�η>���>wi?>���=Tq���t��2_���F���>��>����$J��(��������*��-s>�O?��@>�P?P4H?�M?�)i?#�"?J�>�&�>*W���￾s?��?�7	>\�\��I�]�B� �1���>WD&?�;V�}d�>�u?��?�?�ZV??�,?�:>����Z@����>�f�>vRQ�l���ܚ(>$�W?CG�>�'P?�~?�>~�/�������ͽʔ&>��T=z6?B62?�)?��>0�>����r�>�V?�#R?��t?xyx?�F�=�@??�߆>��?����˻t>~g?q1?��N?(�?2�a?.��>_��"ս�m==9�i"�<�*�=�ʼ;)�=Ue��!��E�=s��= /ڼ�W���XK=�`<�^��Lz�����6�>�*t>L���͌1>f2ž��-�@>D����E�������9�'y�=h �>2?�>z#�K��=0��>���>����(?��??�RV;(~b��ھ�kJ�߰>g�A?��=M�l�s��0v��m=��m?j^?��W�|��N�b?��]?<h��=��þ��b����b�O??�
?2�G���>��~?c�q?X��>�e�):n�)��Db��j� Ѷ=\r�>KX�S�d��?�>n�7?�N�>)�b>%�=au۾�w��q��i?��?�?���?+*>��n�Y4�H����N���v]?���>�����l"?t��ۈо�)�������Xᾟ��+T��������������C�ֽ\c�=FI?L:r?F�r?`?��J�c�z_�_߀���S��F���(D���E���B���m��������b��6=��[�#BG�\^�?f�3?������>��U�^���jЮ�L<�=e���Z���C>�;��_	W<�f>cjn�Ø&� n���#?�m�>���>7�B?��[�!�=���>�v;P�<nľy�?>��>���>#
�>�%��17�Hf���,߾�͚�o�v݀>*�_?�mU?x7f?�t�(	/��C���<�T��:g��0�>&ek=I~�>��0;W�� �:��~BU�(��)��J��g�<��&?X9�>�+�>5�?3?�7 ��\��K@����-��;�=�PB>�J�?�4�>���>���Z��0#�>:/l?�j�>Ai�>�|��\�$�� g�����Į�>D��>�T?\\>	C+�.H[�UV��'Տ�\(2�3�.>��g?����Έ}��oo>P�M?Kq�;�a@=�ʟ>k�[��V%�t�5�H��>Q?_M�=||c>`Ħ����S�t��{���(?6?�R����)�_�|>��!?���>ˋ�>�"�?C�>�X��x{���U?r�^?Z9J?lA?�P�>��)=谴�ĵɽ�((�0�(=%�>Z>dEz=���=�����Y����#?=�n�=.�ּ�۶��c<TY̼'(< � =5M4>zRܿ�gR�߶Ͼ[f���ɾ���fb�������1���q���Jľr]ӾR5��m8�~;��x���d��6����r��l�?D��?J���z��م���zo�3j�Qд>�D�!�;��վ�G<���\�Ծ疾�!'�.b���m��c\��]?j�7���Կ���v"���W?�1?��?!/�׬��X�`�>��
>�%f����>֏�M�ſ#*˾�*z?{��>V� ��#���.?���>S=(<iei>�����>[���<����>n?'?>����ٿ������$��P�?��@�|A?@�(���쾨"V=D��>��	?��?> U1��H�M ���S�>�;�?V��?�sM=C�W�J�	�-e?E�<��F�pݻ2�=�F�=�T=T���J>�R�>~��QOA�?ܽ��4>�څ>	�"�;��3�^����<��]>/�ս?��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=[���oͿ�������	> �S���Խz.ٽ}��s��<�X��)���'?�sϮ=���=��(>���> > >\[>C�e?��v?���>T)�=̈=��:����<�j�82<W�߾%���ϻ��ޔܾ�z��Z�3�)�	��������&ە;�>W�j���zC���S�}�H�܏6?z�=��b��i������ܾ.����ݝ=i+�	Ǿ��O��g��E�?�`?��l�rAf��J���׼j�����a?Ќ���7��֧��v��<�;�'�P�>w�>�m����:��W��k0?+a?�����S��g *>^���=��+?��?<[<�8�>�@%?m�*�~R�/[>qa3>ף>���>rM	>�!��P}۽P{?�~T?���'朾�ߐ>ZY��^�z���_=>�5���輓�[>��<�݌�'�T����Q�<Y[U?���>�j*�>��Q����7��`=|mw?Ҵ?���>Ԍk?0*A?�c�<wK��WT�����w=�Y?Ti?j>?�����о�`����4?��e?�N>4f���뾩Q2�C>�?ho? 6?�-�˦y��ԑ��=���5?��v?s^�xs�����N�V�e=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?��;<��N��=�;?m\�>�O��>ƾ�z������1�q=�"�>���~ev����R,�f�8?ݠ�?���>�������(>�����f�?.��?U=��Yb���~���g�V��:>��=�@��; �s7��V����V����?8|u>��@�VS��K�>�戼H�޿w��8R��cM� (�,D-?���>þO�N���_���v���D�3t8�Y�ھ�0�>u�>eܔ������{�4f;��D����>hq�#�>��S��)��1����5< ؒ>*��>g��>� ��-ٽ���?�c���6ο���ؕ��X?�c�?�i�?�a?j�4</�v��^{��X�s%G?rs?AZ?��$�P']���7���?�4���$k�l/�"��,s�=i*/?��>�P/��zw��,�;��@?l��>&nU��ʿX����8�ظ�?n��?�!�N �>���?R�.?9$�2ʸ�	�u��a��:��9?y�>��E/��8M��ɺ��%�>��!?����"�\�_?+�a�N�p���-���ƽ�ۡ>�0��e\�'N�����Xe����@y����?N^�?i�?Ե�� #�f6%?�>d����8Ǿ��<���>�(�>*N>dH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�"�>��?Ks�=1c�>�[�=��ܢ,�h#>��=��>���?��M?�K�>U�=��8�2/��XF��ER�$���C�*�>�a?"�L?�Pb>p!��
2�H!�tͽ�h1��;�P@�Ǟ,�߽ͨx,5>��=>x>�D�	
Ӿ��?+p�0�ؿ�i��Kp'�u54?e��>�?����t�����;_?Jz�>�6��+���%���B�b��?�G�?#�?��׾iS̼
>#�>�I�>��Խ����s�����7>�B?&��D��]�o���>���?��@�ծ?Ji��	?���P��+a~���7����=��7?�0�Z�z>��>t�=�nv�Ի��Z�s�=��>�B�?�{�?7��>�l?��o�>�B���1=M�>֜k?�s?�Oo��󾴰B>K�?��������K��f?�
@mu@.�^?Ahֿ�����N��������=F��=ą2>6�ٽ`\�=��7=��8��8��x��=N�>��d>$q>�'O>d`;>{�)>����!�r��N���.�C�������Z�8��#Xv�z��3��2���3A���/ýQ|���Q��2&��<`����=��U?)�T?��t?WS�>,q���&>�^��>�|<S5
��>4��>.�3?�=?�T9?��'>F�]�9aW�
!~������J��>��K>>�>}�>N�>(|=�,h>ޯ>aJ�>e�+>��8<�ޠ��\=�*�>���>ge�>&r�>���>�)�>�ϭ���¿{CR�,:�:����?��Ͼ�1��T���û�)���b܏���.?��d>������ӿx
����U?X��s�.��f�E��f�)?uR?��>筡��=��U>8��Jq���=��S���;3���G>O>%?9�f>ju>n�3�zf8���P��v��}]|>936?�궾�99�]�u�M�H�qfݾFM>�ž>c(D�Zk��������ki���{=ru:?�?'H���߰���u��>���MR>q8\>x[=�j�=$UM>9dc���ƽH�tl.=��=�^>��?vU8>�~=��>oa����_����>�2?>?�,>+�>?��&?��'�y뙽�7�6�~a>�p�>E��>�h	>�T���=���>Zr]>?rüdMn��
��a;��J>K��X�[���Q�v��=r����	>���=V�B�2��i1=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�K�>&��W��	��q�u��V"=V��>1-H?LE����P��=��d
??n������ȿ>dv���>���?G�?��m��7��j�?��f�>͜�?WY?]i><u۾H6[��J�>�@?�R?;
�>����&���?�ʶ?$��?�f>AB�?�m?���>r��gp?��湿�Y����g>�h��R.�>�b>F���o.�*J��5Gv�t�d��W�5�>��<q~�>�b��;ﾨ�!>�(ӽ�޾�o�b��>��>܆>|�O>��>��#?i��>NU��r����Jh��۶�{�K?���?���2n��M�<��="�^��&?I4?3j[�`�Ͼ�ը>�\?i?�[?d�>.��I>��C迿>~��]��<j�K>)4�>�H�>%���FK>��Ծ�4D�Rp�>�ϗ>
����?ھ-��FM��WB�>�e!?���>�Ү=� ?�#?izj>�=�>�oE��=��;�E��H�>*��>�?��~?F�?e��9V3�$���ۡ��[�hN>��x?�?y��>a���-�����=��	J�wܓ�\x�?]g?\O佳?��?W??��A?�=f>���I�׾K������>�!?3�ӺA��R&�����?�H?u��>pp��,�սj׼��������?�%\?�7&?����+a���¾���<>�"��]�Oz�;��F�̭>1>x����=J>�ְ=d[m�^6��e<���=Bz�>L��=�E7�����/=,?��G�ۃ���=��r�?xD���>�IL>����^?hl=��{�����x��	U�� �?���?Zk�?^��@�h��$=?�?S	?m"�>�J���}޾5���Pw�~x��w�[�>���>�l���J���ٙ���F��]�ŽD&���?ˑ�>�l?��>�a�=��>X����	��|Ծ��˾�@W��|��7���9�A�.�Ə��ж� ��<ʡҾ#ㄾIQ>2���	�>�U?h�>|�k>�G�>�&�N)g>g�e>M�>i��>�Ж>$hs>��.>�58=�����KR?5����'���辿���e3B?~qd?1�>�i�0������J�?j��?�r�?�<v>�~h��,+�n?b>�>v���p
?�R:=`8�!*�<V��7���3����᪎>ME׽� :��M��nf��j
?�/?���W�̾�<׽b���)$n=(F�?�(?G�)���Q�C�o��W�%S�z���dh�D���l�$���p��㏿n^���!��m�(��)=�*? �?̂�������Fk��*?��Af>��>{?�>̱�>�dI>��	��1���]��O'�ꃾZ$�>�E{?:!h>��V?�_E?��>?��>�.3>���>ᝧ���?�E�=���>��>�?ә)?�
C?�?�)Z?��>�t���΄�^�>��>2�?��>c2?�f	���1=�(�=�T�)]������,r����=[4��½i<>iF>�O?���_�8�/���OHk>#�7?Gn�>���>) ���,���U�<��>W�
?�B�>����#zr�`�[D�>@��?ѥ��V=$�)>���=�K����׺9�=�����Ð=I~��OC;���<<4�=xɔ=��g�V�˹W"�:�;P��<�t�>:�?���>�C�>�@��W� �T���d�=vY>�S>>�Eپ�}���$����g�]y>�w�?�z�?��f=j�=��=B}���U��g��I�����<��?.J#?XT?\��?T�=?(j#?��>�*�[M���^��s��}�?>t,?/=�>�Z�B�ʾ睨��.3���?��?0a�[�Uc)�3N��fѽ��>�/�6_~�)���[C�Xo�����\����?Д�?�yD�A�7����0���=ڬ��tC?}��>�Ҥ>p�>�)���g���Sr:>+S�>,�Q?m��>12P?�Ax?\�Q?��<��G�cɲ��C���L>i�O>�4X?��Y?�z?1D�?���>���=����žu��]�ｙ���������J*"><�>�#�>�!�>�,���
=�U��'�����>���>��?�{p>��?�'t>��D=��G?p�>�-��N~��夾�σ�Iy<���u?Ȗ�?0{+?ҧ=ws���E�"��m[�>p�?f��?/3*?��S���=��ּ��5r�m�>K�>�B�>/�=�G=O>k��>�|�>�D�:D�yp8�InN���?$F?�ۻ=|���U.q���k�����?]m�=���U=�ھ䭁>���Sj���09$���s��8_���X��;⎾�f?���<�t��M���=���=+l�=��=�az<n�Ž����	>�(g;�W���.=�2:K�d����9E*<;˾*�}?�;I?K�+?޹C?��y>vR>�3�y��>�s���C?#V>܉P�Uy���[;�����;��ҝؾLx׾!	d�6ן��O>',I�>�>�33>�J�=��<'�=��s=���=�zO�=7�=�E�=�^�=|��=��>,]>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��5>�>�uR��1��W���^�|r[��p!?�_;��q˾�D�>}�=4�޾X�ž�s/=��5>}Da=����[�/�=j|��2=pb=Ma�>��C>Ǿ�={���X�= �B=�8�=��O>�Z����:���&�.�/=~��=�oa>t�%>�$�>�?��2? f?`L�>�/��CľvR���>Vļ=la�>W�=X%Y>���>'k=?�qM?KN?�צ>���<k�>�9�>�)�+l�G�۾�c��yG�<�D�?&��?�>}�<�q>�q���Z4���U�?�4? i
?IЛ>V?����Ϟ �����D�����<ꜳ=Yuw���z��1ڽƌ��
�=k��> ��>�τ>Ym>�j>�!>��>���=�_=~%=�>O���,���<}=_"��\>.���?y����=���� ڽ�K0�X��=H�R��;�M�=��>=�>v��>c�=����5>���*�K���=�����A��lc���}���/�p�=� �A>'�_>v^x�<����?FOT>.�>>��?�u?gX!>���Jp׾���;&g�v�O��)�=�h>H5��H9��}^��iL�,mо���>�j�>�xo>i�^>�%$�S\m���,>|w��7 ���>�;/��ח��'m�����z���o���"k�̊>[J\?�"��@�Q>;)?�4?{2?�5�>tOd<K����+�>=z��Ь>��/���v�r-9>>?���>�2?n����N]���ɾh ����>�cD��P��啿1,��ƻ����q�>󸣾��Ҿ�v2�A���1�E�� s��ٽ>�:O?LF�?�CV�e��v8N����q��Q?��d?�?�>7�?K	?t��9��
j���=��k?O~�?I�?�>��=�|����>6�?�ɖ?7��?I#s?��>��&�>�ܒ;�q>����v�=�.>��=j��=nh?vj
?�|
?�5��ͼ	���!5�	�]��n�<l��="9�>e�>f�q>�}�=Plg=>�=�~[>��>��>�d>���>EZ�>����	�x��>Ԭ%>P��=	�?4�>	H�=ȃ�8}�#���Y3�5�<�z(��[��{7=w=�f�=ߴ�=�\�>~̿!(�?���>!�-��;%?G���|�6��#|>Z���)�����>�K�>3��> .�>�,?Hd>���:"�=9�Ѿ�q>�G�B�!���B�ddQ�kLѾ'V}>�ʜ��Y%�5�������_J�z���p��Ӗi�1��v�=�1�<�[�?C� ��l���(����à?�@�>±5?ᆋ�I��k >th�>�>[������(܍���ྍ��?�	�?�;c>��>G�W?�?ʒ1�>3��uZ�&�u�j(A�%e�L�`��፿
�����
�D��.�_?�x?(yA?*R�<*:z>P��?��%�[ӏ��)�>�/�"';�@<=y+�>*��#�`�v�Ӿ��þ8��HF>��o?8%�?qY?>TV��2�r5>�?V?��=?
e?Lw2?��D?h*ܽ��'?��]>E�?I�	?�%?��0?�?-�>�_>_�=4����|��[\���_ν�o�.),��j�<�ߊ=�S�=@��̥��"v=(=�_;�A������c�$;4�(=�']=I�=Z�>I`?�^�>P��>��3?�b���2�l���#�/?�$=�Dr�D���ޝ�%i龟�>^�k?���?7_Z?�W>�B��qD�ޕ>E�>9�>1�o>�j�>�|뽆.9�%ċ=l>ȁ>���=�w$����9J�Ч���/=w�!>K��>40|>����'>�}��2z���d>��Q��˺�N�S�:�G�h�1��~v��Y�>*�K?��?���=�^龕/���Hf��/)?Q]<?�NM?�?&�=��۾�9���J��>���>�r�<&�������"����:�n��:��s>72���k��LQ>������o;���_".�I���'����>B�,�D��ۋ���b�=7��=d;!S0�W�|����.S>?֑�=�߭��sO�9Ws�9h%=�w>A�>�� =�[�<�7e��<ʾ�Z<>q��>�=��X�z2վ;0!������>��F?�^?^��?�P��R����M�vd�N�u��rk?VA�>��>.U>E�P���������h��=����>�
?����I�mp�m���o5;��"X>?j��=E�?+Xn?��?��]?vM'?]��>���>+�r��f����?Î�?��D>5&p��P>�S�2���-����>O*#?TJ��ܞ>��&?�+?�?t�X?�U?�>�)�b�C��/�>&<�>)�]�!T����>ҍS?n�>��U?r?w?�F1>f&-�����;�tm<C��=e�1?O?p�?Q��>J*�>�e��.g!>��>?1?`4i?/^2>1�/?)�]��?�Ȭ=�Ш=MÞ>�;?��D?�و?�A�?�Wl>���<o(��v��I���<����i�� �<8��������S�=��;�[��{�@<��:����1��={��=%\�>k�s>��G�0>"�ľ�J�� �@>�7��eG��[����z:����=Fz�>��?ؔ�>BP#�_��==��>�K�>@��1(?l�??z�;O�b���ھ��K�b�>�B?n��=��l��|��;�u��2h=��m?d�^?l�W�/)����b?��]?-k�M=���þV�b�h�龺�O?��
?ԲG�%׳>0�~?6�q?0��>r�e��7n�����Cb�k���=�}�>�T���d�9-�>ђ7??P�>�b>[>�=]}۾2�w��e��r?4�? �?���?�+*>.�n�h2�2��6S���T?�W�>	˾a�?`�=I5۾�W�����'þƅ��ǌ��O憾w����ݽg���d�
��&>��?�?d?TG}?�<r?b��}�e�,,i�����e�Q��������R�:�f*<�e7�u�i�r:�H��������Px�%�B�)ʳ?Y|(?G�=�V$�>�u��n���̾��<>jG��֡�8Л=_��c�=0Yz=�Ul�5�3��g���W ?��>fg�>p�@?��Z��>��)4�L�9�;��K*5>���>O�>���>�X;r81�N�ͽ�aǾ�,��El�8�>�e?��Q?Ğm?-�D��:����4��-M��\���@�>TC>o{�>3֩�TH��2��=�(�j����(˕�i.����=�&?�`>�(�>m��?L@?c4�����\�	<:�"�b=m"�>��s?Ʊ�>��>�b��M���z�>ypj?���>���>`����$��P��}��W=�>O��>��??�C>�S��eT��Ɛ��U����9�^	>ĕp?|hb�{��D�_>]K?��6I=���>*�H�1��}kݾI���N� >��?��>�6�=�S��N�޺d�͞2��'?6�
?����ë,��>P�'?�$�>�[�>Zҁ?�#�>��ʾ�P�W2?:�[?=F?��<?��>fP9=j꽽��9�!��=��>J�Y>�k=�U�=(���{V��j!��X=�X�=w��v���K
�;	�	���}<��=�s0>a�ӿ�G�Vᾡ���2ݾ`��{���p����P���F���s߾`����i��Tg��$��w��&���쇾6%�?�e�?����i���LH��%�Z� V�]U�>��^Fc=�̾ Fh��Ծ���Iھ*y)�%�A��ჿ��e�;�D?a�`Ϳ~ӟ�K]�s7?)?��o?�S2�5
�#�Q��I7>&ٖ��\u����_�����տn����I?��><U���ѽ�E ?���=���:���>.qھ�־�m	=ze�>f?�$?Z������5�Կ(;޼��?Ʌ@�|A?6�(���쾝V=���>֑	?G�?>�R1�@I�7���AR�>b;�?r��?!}M=��W�-�	��~e?8�<��F�'�ݻ=�=e<�=�D=r����J>�U�>C���RA�?ܽڳ4>lڅ>{"�Ѫ�Y�^�ꋾ<އ]>��ս7A��/Մ?{\�qf�~�/��T���T>��T? +�>�:�=��,?A7H�X}Ͽ �\��*a?�0�?���?2�(?ۿ��ؚ>x�ܾ��M?UD6?���>�d&��t�p��=c7��~��3���&V�`��=M��>4�>��,�Ջ���O��J�����=���Sп0�)��p�/51=����>UŽҚd�\tp�)1��=>���#=��0;�� >Ǒ�>�>�(�>Q�>]Q?�/R?�B�>�?>�=�j��ӏ���>�\꽲�m�+3��W�;��?���_��h��*���A�674�໿�����d>8%Q�7
������(�*|Y��b1?��C>�}ؽ1��7����֫���X��݇��p>�>rɾ4�<�9���?��n?�vN��_q�u&��k������JR?F�{�Y� �Mz��ݍ>i^X� ���r�>kB�>��ľ�Si�BSF��9*? ?���k����2">*��+�=œ-?�$?�[�:V��>�$?��D��}�S'8>�<>h��>�2�>^�>�?���ٽ�?kL?��֙�@O�>K<־�[l�玿=LQ>I%��,��x�f>��#<�����a�1���Z=�cV?�t�>��)������� (&�L�K=�x?�{?���>8k?�B?9�<�`��*,T�����m= TW?vmi?�
	>'m���ϾE;��]�3?�Oe?�N>O�m�L���+.��C��?��n?�a?7��_�|�

��{A���6?��v?�r^�hs�����b�V�W=�>\�>���>��9�ok�>�>?�#��G��𺿿KY4�#Þ?��@{��?e�;<d����=�;?8\�>_�O��>ƾ{������q�q=�"�>���sev����;R,�h�8?ࠃ?y��>W��������3>�����}�?�݌?���+���	�΃������>�p��˝���ú�j�U�������ܾ�?2=ֆ�>�k@���<���>�^��|��Y�����N�l�A/��?�?E���
�{�dZ\��q�3�4���D���Ӿ�J�>g >�ڜ�J͕��Mz��49��^ڼL�>�U��$��>7�W�!ݸ�Q���z<#ِ>�S�>>��>��Y_��6��?S����̿g���n1��[?zZ�?Q��?G?��<~j�$�q����"*E?�Xt?�ZZ?��F��aY�*�(���j?�@���J`���4�NEE���T>/3?bM�>��-���}=�>X��>1D>|U/�/�ĿL������?Ŗ�?��꾄��>ꗝ?x�+?�X�g8��2�����*�Ew]�X.A?y3>3����!�H=�w�����
?]�0?,6�f$�N�_?�a�N�p���-�*�ƽ�ۡ>��0�!f\�GO��L���Xe����@y����?7^�?X�?��� #�O6%?'�>^����8ǾL�<���>�(�>�)N>G_���u>����:��h	>���?�~�?<j?��������V>��}?�>�?�R�=ZS�>�,�=���&�ˤ#>(~�=�?���?��M?��>~��=�$9�%/�&QF�@4R�����C��>T�a?�lL?�b>�	����0�v!�ͽ��0�b��|@�ۗ,��0߽D5>��=>!�>K]D��Ҿ��?Ep�4�ؿ�i��Fp'��54??��>	�?����t�����;_?Fz�>�6� ,���%���B�[��?�G�??�?��׾ R̼#>�>�I�>G�Խ����c�����7>,�B?Z��D��f�o�r�>���?�@�ծ?^i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?�Qo���i�B>��?"������L��f?�
@u@a�^?*�XܿFj����(]�����<���� T>Ң�==��=���m̽���=�,;>��0>��Z>��>���>�T>�i�>�%�� �B��q���вD�ܡ� ��.6��-���rɌ����� ������w���,���"=�R��p,��K
=���=�>O?`�r?�s?�Y�>�f�0�J>�M��U<����w_>�N�>SQ;?�T?3?�+�=�¼�s�Q���p�Ŗ������Hc�>�v>rl�>;��>�3�>|O^==�i>�˟=���=��%>�z5��?���=�">�3�>�$�>�>�]�>vw�>W����¿�%+��G�M�S�&�?Y(������О�9)��=� �vI='2?�>Zt����ݿa��<
I?b:��W!�ٌ��Ť*��z?5Fb?|e�=���=�ͽ���>%��=�+�T%Q� �-�Kw���i���U=�:?�e>59u>��3��9�2�N�%����u>kI5?v�����2�?�u���H��޾G�K>߽>��^����������~�S�f��y=��9?�?Xo���ί��Qu�H`��~QP>x�]>0t=�o�=��L>�a�O2Žr�G���=��=#�[>OZ?�,>/[�=S[�>�����$T�g\�>�yL>�:>�77?�#? �J��g��ň������>�X�>�U�>B�>�aB�5�=c-�>��T>�1���~��W��V�H�`>�ּ.�R�8n�>�=�9�����=�Ֆ=�����8�%�}=�~?���(䈿���c���lD?4+?v �=�F<o�"�H ���H��;�?k�@m�?��	��V�<�?�@�?�
����=}�> ׫>�ξ9�L��?c�Ž.Ǣ�͔	�Y)#�dS�?��?i�/�Pʋ�9l�s6>�^%?�Ӿ͓�>i��EL���`���:v����<!%�>�OE?��3V��$1�N�?�� ?�a�Ƥ��ɿ6]v�>��>,��?~ޓ?f�p����:�׷�>�M�?f�V?�R>Z�ܾ�^�$��>�>?�R?�ݹ>q������?[*�?.O�?Fa>ɚ�?G.p?���>��RuD��踿[���:	>������>��>�<���,�xj��yE����f��q��rS>*�<���>������Ѿ���=�a�$ľ`Z��}˷>UT>l�>�*�>��?U%�>��>X���Gv�Np7�̜�_�K?೏?x���4n�cu�<	��=(�^��'?pI4?��Z���ϾJҨ>�\?���?�[?�c�>J���>���迿�z��=�<��K>/�>�B�>�+��XIK>��Ծ�2D��i�>]ї>ɣ�~Aھ�+����pE�>jd!?���>�Ϯ=U{ ?�#?�>j>��>;dE��4��H�E�}��>��>�?j�~?��?�ﹾJL3����硿m�[���M>p�x?�1?ȁ�>#{��,\��`JL�y}H�ܹ��q[�?�Yg?�L��?�'�?�|??�A?Rf>�;���׾Fج�t��>e ?�<�;�B��&)�P�ٽ;�?��>#��>�蜽����U�H��d!�G�����?͜W?dM!?���?\���ľ%:=����5��=��;�'t�֓>�!>BNN���=1�>m8�=pg�3�-��ן<X�=|��>C��=�`5�Ε��,=,?B�G�tۃ���=��r�2xD���>�IL>�����^?Cl=�	�{�����x���U��?���?Uk�?���-�h��$=?�?E	?l"�>�J���}޾7��dPw��}x��w�V�>���>��l���A���͙���F����Ž\����?q@�>���>4�>ǽ>#��>Z���2���� ���ݾV�U���#��n9���5��+����SqA�ĩ�<��̾�w8��I>8����>
�>A��>��=*�?j�	>*f7>�{>�K>d.�>A"�>'C/>|�!>}�2>�?~��BR?����2�'�~��@��6OB??d?�+�>��i�=g��[��VI?%y�?i�?�v>��h�<0+�9e?���>���E~
?w�:=�@�|E�<L����j�y̆��O�_u�>�ؽ��9�M�,\f�hj
?�$?���n�̾�Kؽ����07o=BL�?\�(?��)�(�Q�	�o���W�S�����%h�Y��\�$���p��폿{\��+$��٣(��w*=Յ*?o�?��ۗ���'k��#?��Af>��>��>�>'�I>��	�ʷ1�*�]��M'�'���>P�>�Q{?�z�>�Z;?�=L?]EQ?��H?�~�>ػ�>S����� ?�.�="�>���>��W?Q�?�61?v�$?��G?��>Ʒ0���ɾ(��`��>o�?SL?g?)�>�� �9����W>c<;eZ�����<]�>���S�R����#>��C>�??%	�m�:�c����>��@?�E�>�@�>u��w�8�������>�?d8�>J����wr�26���>��y?����]*=�T">��=�]��ו��l�=j�a�\�=������O�<�G�="G�=r���Ed��*-��iSI�=dE;��>?�1�>��>#3���� �'�T�=X�Y>��R>Jm>Y'پ!v��d
��_�g��w>&7�?�F�?Qk={S�=n��=M����!��� �����u��<��?c#?>jT?9��?H�=?�[#?�9>Z��(���\��MA����?��G?᩟>��#�M^�4����G4�29?�@?<���;{�v�G�&'���_2�����|]�\���5��?I����>)��v�|`�?��?|�r=jxe����4���
��YfC?R�?�zi>#?�*�F���?�"����>��?�	m?��>��Y?��?,:b?'=�:�a�T���ҭ��O�<=��<�ye?�R�?���?��?�Z�>���=<����Ӿi�<'̽�6�����q9��L>Ҹ>�?=z�>���ѐڻf�ݽ�����}
>cT>T�(?�>�.�>Nq�>7b��-{G?�M�>4��-Z�K{��t₾F+���t?��?@|*?O]=����E�����w�>;��?|�?e9*?�BS���=�`ͼ����Fq�m�>��>WĖ>H�=&�\=�� >g�>o�>�#�0d�_�7�+�X�1;?�:E?>��=	Ӱ���Y� ���Ҿ1�^>9�6��O¾嫻�l|�ؕ>�-̾>@���_����B��t��݄��#�;=����ҋ�> ?ֻo=\Ñ=���=-�u=﮼�td=p3>=(=I�)�����<Z�S=ݦ��Vb��&�J<�/�=�+��Rɾ�}?ϑE?})?�A?Νj>�&>���?|�>N���}?ܭP>㏁�-7��i�D��!���Q��`>վu�ξie�����6��=� P�k�>��.>��=2�	���=ޜ�=�O�=M�Q:�(=��=]Ȱ=�Y�=���=.�>4>�6w?V���	����4Q��Z罡�:?�8�>r{�=��ƾi@?��>>�2������xb��-?���?�T�?@�?Fti��d�>F���㎽�q�=g����=2>c��=x�2�U��>��J>���K��/����4�?��@��??�ዿϢϿ2a/>Q�/>�8>}�P��5��y5���)�œx� �?I;��޴��z>�q�=��MǾ��2=��,>��=��v�Y����=�����.=�Ă=��>¸P>=�=h�νd��=���=L��=3B>ov���%�%�+�3�=�-z=i�j>H>eX�>v�?�<8?�e?���>�Iu�
c�������+�>�9�=g\�>��=�:>-,�>1�;?IF?�G?�Q�>~%=9�>��>_l/��l��ʾC1��:=Q�?�a�?�L�>�8��>;�0\��?�ˊ۽5?faA?@?��>%����HQ3���<c"��U���,��\F�50��' m�]�_�w(��|�=�_>n��>q�>6��>��>�1�>�R�>�52>��>�5g;�O����=LP=;�ջsV��}F���G��½H�K<�1">��)�����6����+=%�4�{��=���>`!>��>5��=�ܳ�A/>b�����L�o��=k7���*B�15d�nF~��/��u6��B>��W>3i��,����?W�Y>�k?>Z��?jFu?��> I���վaB���*e�&S�Pl�=��>��<�h;�V`� �M��zҾ�G�>Rd�>���>��2>?l:�o�O�H��<���-���uώ>����@��0W�}(��>f���-��81w�ұ,�|j?w��KL >$�h?��U?��l?Ʒ�>������?�"�o��>���W n�Vk>�03?_?M?�(?�iԾ��m�L:̾C���_ʷ>P;I���O�����n�0�l��0���`�>=⪾9�о�$3�|e��9���G�B�*Zr��պ>�O?��?�!b��U���HO�����慽�|?�]g?�>�>}L??4?y����t�J����=�n?n��?b8�?	>��=�l���8�>Tz	?Y�?;�?g;s?U\>����>�D�;�$>�x����=��>���=��=`�?��
?�	?N�@z	������X��=D��=@�>��>~w>���=�6S=޳�=�6]>MÛ>���>n�j>�Ӥ>⤉>�r��F�۾,��>����=>��/?2�h>: ������)=p�=χ`��\����۽1�`�]�g�˦���;V^>���>�ſ-��?ob�>�Dɾ�4?�~��qY��E��.9n>������>u'>�i�>t�>�?ع*��!>���=DҾ�:>�q�!���@��)P�,Ӿp�w>�X��U�����w� ��VJ�����v���i����>Y<��ָ<E�?j?��%pk��?)�0����d?��>kO5?G����m��� >K7�>�s�>����)��(R��9���΋?��?�:c>�>��W?&�?	�1��3�vvZ���u�0(A�Ae��`�\፿ٜ����
�b���_?�x?xA?�2�<�;z>���?�%�aӏ�K+�>�/��&;�dB<=�+�>�&����`�{�Ӿ��þ�5��EF>q�o?�$�?Y?lSV��<���=&Ia?�oL?�n?t�+?t/<?"�����<?u�>�?���>b,?�+?Q�?��>�B�>��e>8z����B��ț��,��X���T�e�p=�h�=�=��=?� ;\E�<���"޽/<�Xa�f��w�M=n�2=b�=�Ҧ>t]?���>ē�>K7?����7�)��hv/?�D:=�����슾j����?>��j?��?_HZ?/Ed>i3A��C�|�>�܉>^�)>�s[>q�>��;�C���=�R>?[>�Ʀ=��D��)����	��(��y'�<�$!>���>A2|>���<�'>x��z�Ϙd>��Q�|̺��S��G�G�1��v��U�>��K?d�?Η�=O_�0��Ff��-)?+]<?�MM?��?,�=�۾4�9��J�c1��>���<���ݿ���!����:����:�s>�0��+%�o>�a��ھ��p�էC��!��(=/�==w=�1�ܾ��p��t�=��>þU!�e0������\�H?f�\=6Ϩ�ǽZ� ���H$>���>�>�A�_�j���<��Z��P��=�2�>~yD>�?��辟/B����È>anR?��L?��_?'X�5:���^�>�+��''�R��>�Y�=
#?Ӫ�=nZ>]����#�y�u�ktP��D�>=n�>���uwF����Jp���#8�r�>���>oZ> 5�>�.?�qA?w?y�(?�?w�r>&�<1홾�~%?���?�W�=V,ؽ``���4�*�H�~��>~�&?��I�`�>(�?mj?�%?�NR?{�?q�>[��@�Mϖ>o�>l�W�u����i>��J?�K�>KZ?�/�?�?>�2�����l֌�i+�=��#>�@1?f="?2�?��>��>���a$�=���>�'f?��z?p�m?�t�=?T�`>���>�=�#�>���>e�?F�N?�/t? �A?@��>R"<ٌ��Zý�퓽l��Z��:(��;{k=0����&Q�w�!��pq;��<��w�����k�-�N���u���3���H�>%r>�󔾝�.>�	ƾ�@���L@>�����Û�zԊ�G�:��q�=�Y�>z?&=�>A�#��ҏ=J��>"�>�k�"(?UH?�S?��1;�}b��ھ�~N��ޯ>�0B?%Z�=اl�׬��5Ov��~`=�5m?G�^?��Y�����2�b?I�]?�s�;=��þ��b��龈�O?�
?��G�z�>��~?��q?a��>F	f�z7n�y���Bb���j�N��=�r�>wV���d�^�>��7?B�>��b>o��=Z�۾��w�Oy���?r�?^�?F��?�*>��n��/࿺�Ӿ乏���[?�ߓ>�3ﾒqG?YV��ZɾHg�����6mپ7렾�i��'ݽ�~־�g@������	�|�P>n�?�tc?�?Fc?�l꾝+Z�3/N�ړ����V��"���g�#@��j`�)W��r����<n��B�;>�=9�w�$@�ѩ�?x�%?�W8��n�>x�����@ʾ��D>����!)��=cia=i�=W�d��[4������?-�>r��>�%>?_nW�5E9��,��95�?���~�@>ܱ�>Ͱ�>�{�>��+�^�2�� ��ƾ�ǉ�^���u>2�d?�UJ? "k?�.�W,��炿_�#���4�����4+><O�=��>1hn���x'�d�=�Dw�Z��_m���@�Y?�=��'?岂>a��>2�?so?f>	�8�����p'0�է=�u�>eg?N��>b>_-���<����>�l?C��>F��>�܌��)!���{���˽��>�)�>"��>vp>��,�q�[�$_���P���8�0$�=��h?~���`����>�R?���:�E<��>-�q���!����(��>I[?��=�g<>-ož?��{�������!?�P#?�4b�����X�>�]?���>5�Y>��??B�>�����;T��>Q�J?��&?�Q?a�?C��=r�.<gؽ������=4�>?�>�Q����\>�B4=�-�1gG�m�;����.�=�)�	0>A��=��>��K��g�<kۿ�cK�lپ����S�JW
�j��a��O���N%	�9��X'��"�x����^*��LW��bc�����1Im�Z�?,��?R�����ć���I���S��[S�>��p�}�"3�����!�����b���e	!�ـO�}�h�0|e��Q?7���߆ؿ�{����ý|�&?6?��?k���D� ��0!=;�^=e�!>9V���V���kݿ����9F?Z��>���j���>�Ρ=��B��v�>��㼋{q��]Q�.p%?���?),?}Ľ����qw⿣���*�?��@�xA?��(����q	V=д�>��	?m�?>�b1�5:�%谾D�>�5�?5��?"{M=�W��x	�A{e?Ռ<��F�+s޻��=@R�=��=���L}J>Ix�>�d�9A��`ܽJ�4>�م>��"�|�� �^�.�<~m]>��սr&��5Մ?+{\��f���/��T��U>��T?�*�>Y:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�܅�=x6�����z���&V�|��=[��>c�>��,������O��I��V��=�5Sſ���S����J=�~X��� ��_��߽.���%Y���I�;3��i_ =x'V=L_�=�}W>�r2>#n2>�W?��{?���>�2_>����c�Aȯ��00���c��0ֽwi潂Ud�A����W�����r�%g�i���r����(��:��I�@��\r�k����`W��k)�Xk8?�+c<X�,|*�sݍ�,e������a��/ֻ:q�����싿aT�?˯?pۜ��Y��/&�Y�>_�ý�8=?����t2��I˾�=6�P=� �w�\>���>�ex��O�.�[�0k.?��&?_���x��C�>�޽xϷ<Qq?�_?�B0=�C�>o�"?����ۤ��J>=GR>i��>���>}F%>$����c���4?8�R?�D�����J�>�̝�^�[�o^<���=�d#�r�üAFP>�v=/	��2�C���}t%�Y�V?׻�>@#(�N�[��#��z
=�/t?��?�s�>�j?b�B?Ǧ�<��XqT���Oߓ=��X?wj?C>�|��kѾ�O���4?�>c?g=a>�]��E���/�P�S�?��k?��?m����|�d?���$��4?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?t�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������h#>�Å��9�?��?��v��=���?q�4��n�W��a>����մ��0��nQ���(��W+��
�<=�@>c@-𗾪�*?5����jIڌ�����oy��	?!�y>��ľ����������K��oQ��v��բ>Gz�=��
�C᛾Fu��-������>J+�����=^�Q�<X�����V���bD>�M�>*��><��7��	�?���ο����G��K�h?���?�x?�H?�j���Vx����4�a��??�5z?�1a?UZ���/������h?�nھ�6���R0�O�W�vv=W�5? �*?^'h��o��5?�]?jݺ=0�	��i��oh̿�'��7�?�:�?�x	�m�5?uÆ?TA?&*������Ǟ� )7�h฾.dl?���>�OԾ�8�]�j�Uo�;��>�^F?g�����`?ib���q��i/��C��p��>>�,���V��6�E�$���d�?����z�ny�?$��?7�?�!��&$��B"?>9�>�.����Ⱦ�Q�<"6�>�˴>��H>ּ@�˫v>yU��9���>3�?���?�C?vÏ�Τ��>G�?�#�>��?w�=Ic�>[b�=갾D-�5^#>�(�=�?��?M�M?$S�>�W�=9�8��/�dYF��ER�#�s�C���>Z�a?��L?Pb>"��V�1�!�Sfͽ>^1��Z��D@�}�,�G�߽�+5>T�=>�>>�D��Ӿ��?Sp�:�ؿj��#p'��54?A��>"�?��Ѵt�v���;_?[z�>�6��+���%���B�g��?�G�?3�?}�׾�P̼>��>�I�>�Խu���}�����7>J�B?P��D��s�o�X�>���?	�@�ծ?Si�	?+ �jP��_`~�G���7�d��=�7?/1���z>]��>P�=nv�㻪���s�b��>&B�?3{�?��>˯l?рo���B���1=�J�>��k?�r?�$o���!�B>_�?���"���{L��f?��
@=u@��^?v�ۿ�A��h��-nѾ�l=���= U>����>_&�=��Z���y�]�!��>?T>f>>�y`>p�=���=b����k!��5��/����4�f��,��m�	��������y����Ѿ�}ھ�����Q�T�۽�r���4T�:���B�=>��B?�??�x?�/�>w-�=v瓼'���'���VSԼ�ch> J?�$?k�B?AV�=��9�� a��@|�^\���Y�1�>��n>���>FZ�>N<E>l+���>��^>��`>���=/>�<�眽y�A>���>�<?���>��>�b��Z$��=��XA�U)=���<8��?M0Ӿ=�e��?�����N˾-;=�,?�m�>�����Ϳ�i��s�P?������ ��nj�?[�>��#?�6-?so>^&��=��=�c��n-��B�>��W=B���3)_��q/>k�;?�qg>Yw>N3��8���P�G���/Hv>ϣ5?����_�:��Wu���H��(۾mP>��>b��y�p��~�Big�ts=0�9?��?�����ï�38w�_Н�2S>�l]>�0=c��=o�M>�pW�Q�ýC[G�_�8=˯�=Z`^>��?n]<>i��=�>ڹ���PR�(!�>��> TB>��??O�?�C�L���ʁ���"�>9��>�,s>|�>˱A��m=hr�>�hr>�ü��z�����&���R7>S����Zl���S��@k=C}��w�	>�'�=ڕ	��^D�=V&<ǖ~?����㈿�뾏k��amD?+?��=�F<��"� ��^G����?i�@�l�?��	�C�V�J�?�@�?=�����=��>A֫>ξ��L�s�?2ƽjǢ��	��'#�	S�?A�??�/�Zʋ��l�,8>�^%?f�Ӿ�f�>y�IZ��<����u���#=���>z8H?�S����O��>��v
?�?�X�!�����ȿ�|v�p��>��?��?!�m�>��@��w�>��?�eY?afi>ge۾�aZ����>W�@?nR?N�>�9�b�'���?p޶?���?�+L>�u�?h�U?Jm�>�Ȥ���$��-��ʟ��K�<�zĽ[�e>:�n���F���n�U���(e\���H����=Z�-:�>�aͼ�徬ץ<�V$��վ_<���>�b�=%L�<_�@>�D5?�;�>��>k-
>X�Խ��[�Z�ɾ��F?WC�?f����M��ۼ82Y>����>�
?㒽L�˾G�O>��n?�E�?q?W&H>�m�,ݙ�4��?1���3c�4�#>c�?&��>�2����=B��5�h�>Jb�>Np=;ݗ�͉��'<^��>A7?D��>c�#=ؙ ?Ϝ#?��j>@(�>XaE��9��x�E���>��>I?�~?��?�Թ�iZ3�����桿2�[��;N>��x?�U?�ʕ>]���ƃ��LpE�CI�����P��?{tg?�T��? 2�?��??Q�A?*f>��@ؾl�����>�!?~�FA�{&���a�?.�?:��>�ؓ�0Uؽ�༌��G��8|?Z|\?�w%?�w��)a�Xþ�E�<��B����:�<����Z>��>IT�����=�]>��=�5k�<�4���}<���=)o�>!|�=,�6��l��C=,?t�G�݃�(�=��r�yD�I�>�JL>:��;�^?�_=�(�{�L���x��/U�e��?���?k�?� ��n�h��%=?j�?�	? "�>J��p|޾і�?Tw�uxx��w�d�>���>��l�"徂���7����F��� ƽ~����??2>R=�>�?mQ�>�q�>�9��.����P��WJ_�����;��3'�|��7߾�⟾H�e�ITƾ�����=�>��/����>T�?f�>�_.>�U'?�bйŲ7>��.>��\>Ʉ�>k�>�)>���=�@�j��e�Q?)����&���龹���QC?��c?]`�>e��u��b��?�=�?�Ü?�Nr>�!h�N�+�=�?�}�>ד}�m�	?fY=\���M�}<�b�����v����N!�>��ҽV:�MxM�B%h��	?K�?��[���;mFԽ�y��U;o=�E�?�)?�)�
�Q�	�o�/�W��S����^h��e��d�$�+�p��菿Wb��`��/�(�� *=qy*?�$�?���m�� ���1k�9?�f>���>u�>sǾ>�NI><�	�ɸ1���]�FQ'�=���)-�>�-{?�'�>d�J?�	G?��Q?��(?��w=?G�>w	�vL?�k�=��L�>�)?َ3?���>UR?��"?Y ?��>;*�=7ؾ�n����?��>�|?��s>�X?iY���/��
�=/�=�N�=�@Z���>>�i�=Vv9�R�����&=端>gW?����8�J���mk>�7?�~�>��>���h/����<��>��
?�B�>�  �7}r��d�QM�>���?�	��V=u�)>���=�����ҺvR�=���� �=���;���<I~�=��=o�q�6[��]�:�!�;�U�<�� ?z�"?�@�>�Eg>�������ӳ�8�t=��o>�1v>|q0>H�Ӿ�E���}���m�Vu�>��?g��?yA�=q��=ҩ >2��I��^��uҺ����<d&?��#?}L?*ʐ?�9;?��?��> ����i�������?�,?j�>���p˾��ZL2�^?'$?��`�(��+)�%¾kJӽ_�>��/� �}�����B�C�����]�������?x��?��C�jk6�b<��ۘ�}�����C?��>擤>��>6�)��h���TE=>d�>L�Q?'Q�>z{P?tp?|]?�X_>z��s���0k�������:$>+3'?��u?3Ж?�k?x��>�1>�,
���ɾ�V����I�l?Ͻ��4�}P=S|f>��|>b�>�]�>�T�=��p�s��ߠM��X�=��>>���>A�>��>�'�>D�F=vOG?Ū�>���/���h��s�w�b�Ž� h?��?��2?�Jv=�����?��]��5�>%��?<�?�>-?�$.��R�=v�T���ľ�Rt���>�-�>Ք>���=�҄=��>V�>_��>}2���� Q5��Ct�W_?0D?���=%ʾ��Ro���F��i�=@�� �c�P������>Qw��!�T>?�>ɦr��H�#����Dپ**��Qi>��|�?��=t��=���=�=�=5�	�*�=ɮ�=W��ؠ�$�����<v�d�:�o�l,��1�=&-�<^�>�V���ʾE"}?I?�+?�D?xdy>h$>�u5���>��|�h�?�:U>�7U�1p���:�����k���6پ�0׾дc�֪��^>�I���>2>s�=�~�<7<�==p= �=r���=���=շ=�e�=���=d�>>93s?:���㠿Ƣ_�Fg��G?�*�>@-
>�\��J	?�>�������e��1�j?���?�ؽ?``�>kϾ\.�>"���o'��G� �Џ3�|F�>�>�=R��$�>�K�>K�����N�0��?�Q@��,?�D��$Rǿ1B.>�*8>(�>��R�=1�M\�u_��^�**!?;��̾�u�>^�=Wݾ��ľA59=��3>/X=7D� \��i�=�Ɂ��i5=1�p=΀�>�oD>���=l)��
�=V�O=�h�=��P>�����*���#��]3=*��=�gb>*�%>��>�g+?H�D?�Z,?�{�>a��{���R�>ñ>i>-`>��?���>�G?l;?�oV?'�>���=yf�>!��>vS��!���M��^U��+���}?��{?��>1��>;��2��m�@�O5�}�?��f?��>D��>��n���$�8mR�9�s���x�i�=��ĽZݽ䗉�W�T��W�Q�;1r�>�V�>�>�(2>�T�=��A>$O�>J��=�,:=¬=i=�m�� I+�a�>6ߍ�]}��1Ƣ�閝=�5>>f���	�=�	sV���c=�N�=j�m=���=�"�>6&.=9��>�2�=4����K>a�\���a�h�v=�r�5�:��Z�Hu��v�=��i��z�=e2>��:�����N?�v=>�'>�8�?�?\>������`{���'��z���T>�>��ν9���]�a�q��~O�>�U�>U�=u�B>�1,���>����=�㒾�uc�8&�>��1�L�a�AO���y���t࠿�o��i�<��O?6���d�>��Y?J%?�e�?ՙ?e�����Ѿ�l{>.�ƾ?�[��9#����+���?i79?��>+#�
�?��̾L���÷>��H�źO��ƕ��t0�S(�W���!"�>�k��y�о=3��h��I���vtB�`Lr�x7�>�<O?��?Ab��a��nO�����܄��5?(Xg?�˟>3�?��?�ԡ����ό��Oն=��n?&��?�
�?�	>���=��t�r.�>��?E �?0�?�"z?��h����>؏�=���=fL=����=`>/��=�*>D<?f��>�H�>pٗ�����0������[;�@�<��q<�ˆ>gD�>u�=>��=��=���=`ӈ>�fo>#4�>k>�~�>j�>8o�����_˥>�*��>��D?�tu>,�>tP�;���?���b�=�����=�"&�K$�00��v.�<w} >�5�> �տ��?	E8=֜^�ā*?��޾`yT�sؗ>S�>��D�c��>z~>��>��@>�s�>�)>P�>s�>>FӾ�> ��d!�A*C�]�R��Ѿ�z>�����
&�������XAI�n���f�Kj�\.��&<=��н<GG�?����N�k���)������?JY�>�6?�Ռ�#	����>��>ɍ>�C��8���>Ǎ�f���?���?&c>n/�>6�W?�T?[(1�1o3��(Z�L�u�}�@���d���`��͍������i
�����_?��x?CFA?�'�<�y>�i�?Q�%�̏���>�/�}�:��<=c2�>����?�a�"Ӿz�þ��z7G>��o?)�?�&?+4V�@�%��)M>�J?�@?D��?x��>��+?����Q?��>�
�>U�?P<?1`>?kn�>�>Ɉ>�f��-�=*���zYl�����٤���ƽ�v�=��v���X=���>f�^��*�<�l伖��9�b�<ت���e���v�7��<�rI;���>-�U?�?���=�>���G�����$@?��>6b��R������X����=g?��?Ċ/?��>��/��1Z����=�{�>���=�=͋?�!�;�����:0�:��;uu>cO��o1����<�l׾!5ɾ�OH�LIH=�w�>�\{>u���*>�̢���y�8�g>{0S�X���,�P���G���0��`v�Yn�>YAL?n?�ƚ=��龾����e�o�(?��;?wMM?Ԩ?%�=�>ھ<�8���J��C��m�>�4�<�	��H��u���	;���9'�r>�Ο�h}��/� >v����ξrq�:�/�lOɾҡ�=�P�K���n�5�_�5F�=f�>¾���?��^��S�����L?���<E���C��7��W�d>��>ޖ�>ѷ������.(A�}����=K��>i�H>q���,���G=�a�	�m�>cXV?ϙ??Bq�?ß� �n�}�?���e!��۴��s�	?�u�=V�?�|Y=��=�Q����"^����`��ݸ>�q�>�x׾�U�a���Ծ�
�3�=l?�O�>�*�>&�/?�t?^�I?��
?�y?�o>e�;�r���v%?�p�?$ˏ=&�ӽNV��[7��|G�#6�>�(?��G����>*?6�?%�#?�1Q?�?��	>���g@�je�>;j�>)�V�q���]Oe>~J?���>�X?4�?��D>9�4��`������p?�=:�>�I1?u�$?MI?���>�k�>mL��H�=�+�>��h?78t?�Aj?dK�=5�
?�>>�l�>Հ�=��>m��>Y?�K?��m?��F?�<�>�k<J��a*��D�C��lz�X�<z��<&��=�붼ɆJ�����o<�o'���6�/6s�v; �˱���߼��Y:*H�>��s>�畾�B1>Qgľ����'�@>q������⊾�N:��F�=�~�>�?-��>�#�e�=�x�>-=�>����+(?ʶ?�?�nA;��b���ھ��K�<\�>�
B?�6�=A�l�=�����u�r^g=��m?��^?ʹW���u�b?��]?�j�,=�{�þ��b�9����O?I�
?[�G���>��~?P�q?9��>% f��:n����Bb���j�Oȶ=�t�>�X���d��B�>D�7?�M�>0�b>�1�=et۾O�w��q���?��?/�?���?�+*>��n�u3���Ⱦ����N=]?��>�M�QiF?&1�=9��n� ��&��K������;����ʾp�T����	���u�>�	?R~d?7E?�d�?q����u����t;��8LZ��h�����&�W���b�'�#��c�<���:]������~��U����?H?J"~�s		?��Ѿ��$e־j�>�1���LI���=`k����=7�<�͏�A7S�t)�d1?ki�>�f�>��C?��W�2q@�8�0��8�#� �	�u>4��>9�c>�9?�{ļ�r�/�<3�Ӿ�|�p�����>0c?�B?C2]?�J�$p(�Ÿ��	��$�#�ւ��.��>"6 �J�
?v�����,���㾘K��!z���/���p��ξ�&@��AO?s�!?�l»YΚ?ך?�ܾ�`��K��f�y�%=��>n
?z��><ѳ>��T�g�侟��>��l?U��>��>���CX!���{�J�ʽ4%�>�߭>���>��o>*�,�$\��i��҃���9��t�=��h?������`�"�>AR?�K�:��G<G}�>��v�~�!�?��b�'��>a|?���=Ӡ;>�}ž�$�!�{��7��2'?��??���O�'�v�>k?g�>`�>,�?b�>A�ľQ�M<��? �^?�K?/�@?c~�>E8=���YBȽf&�O)=<+�>�qW>�qm=�f�={���V�m!���M=���=v6���X��ܤC<�G�����<,i�<��2>a�ۿ��L�p#ʾ�p���:�&��x��>��c�����Yl��˰��Ƭ~�j��ҡ��\�5~T�q��xs��#�?T�?~�}���_��y��	���v��OS�>�百��b�ȗ��v�k���>־����"�B�RX���]�^"E?�a��$迤����wվ�(?�?g@�?
	3��G@��K�?�'(>�I�<i �?֛���ڿ�y��=�<?1��>Ϝ��Kl	�v��>�.>4�˽L�6>=b<`�G���/���:?ՠ�?!tM?�W˾���0�׿�DZ���?}3@K|A?�(�����V=d��>Js	?O?>�K1�B(�^װ��;�>�/�?y��?DL=h�W�%��C�e?e� <��F�)��E6�=b��=��=����dJ>A��>h���A���ܽt�4>Sׅ>Q�#�����^��I�<Hz]>F�սa��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=9�8�ſ���M��Σ�=_=��w�T�	�b}��0�ӽf����������FA�<�>=�w8>�*e>��=2�&> \?��v?<��>3��>��ҽ�������Q�=`ಾ�Ī�? �U���7����������h����G����+�8�|�<��L�����\+��'`��81��m9?�:�=���g�8���#<�Ӿ5S���ߐ���ɽ��þ"��o��F�?�y1?����Y�����=P����?J?F,A�O�
��������=N�V�26�>��=��޾%�3���Z��+=?��(?K�þ�9 �5�[=18=,�׼a5?kd/?�n޽�>��H?Ƿ�=������>��>?�?Ȱh>�ξ�ؽz�?"�d?DV�=�����?�lh�	KA�4�d�6Η=
Ԏ����>�B]>��+=�/��̙<
����W?�^�>�`)�,������1�
�Q��<'�u?m�?[��>m�g?�SD?���<����ŠS��I	�{��=�X?�%i?i>��/%Ͼ�$��V�2?��d?�db>��i�h���m1��� ���?x�j?��?!�4��}�����wu��V5?��v?�r^�_s�������V��=�>a[�>���>U�9��k�>Ǒ>?�	#�nG�����Y4�	Þ?��@g��?��;<!����=u;?�\�>X�O��>ƾ�v��������q=N!�>����Sev����S,�È8?젃?���>����Ʃ��1>�#��O��?�5�?D�����<;޾�w�w�𾉦��5���]�%�Wm��l ����:�����6E⾋�t�T�v�T>b�@������>r~���׿,qȿ'y{������ۋ����>��>�9z�n1�9"-��T�ְ(�f�k�a����j>Oeٽ�]E�� ��h�������t6>3� ?c���ٽ��<c4������v�-�=�>'/9>ؼ{��
�]S�?��	�y�ʿ�X�����I+�?ޫ�?��H?m_�>:3��\&��P'��9	���?�2i?��A?/	�lۦ��蟾[z?a\�䆿��h��i���e>��5?�JQ?�g�t�/�%�,?�t�>;F�>����Ϳ2ؿ$3���?0��?+p��6?���?�M
?��y~�Yђ�uY��W�D�L?���>2�ؾ>X'���L�Y�Ǿ��>�sA?����~��_?{�a��3q���-�2KȽ'��>&d/�_�Z��2�� �vPe��<��jPz�q �?�:�?�߲?�I�] #�A$?O-�>O�����Ǿ��<���>)J�>��M>��[�qv>x��=;��4>6��?zo�?A?������`�>�}?~�>�$�?���=��>S��=zͲ�N\8���!>���=�@��?eL?}'�>*��=��:�@,.�u�E���R�k���C��s�>�^a?�	L?�b>O���+���!�f��S�)����4�>�g�0�%�ڽ��3>�u>>�Y>��B� �Ӿ��?Xw���ؿ�l���'��04?dă>Z?����t�����8_?���>�.�v+���,�����W��?5G�?�?�׾�+ʼ�>wɭ>�M�>+�Խ����Y����7>�B?���B���o�F �>���?��@�خ?��h��|?�������|��r���7�œ�=��8?5����q>b��>�0�=�v�wv��%!t��z�>p��?���?���>Wpm?�~o�a�C���=&��>��l?��
?G�����@>(�?O��E�t�.�e?��
@4�@�q\?���Ó俧�Uw��������=d�=�w�>l���H��=�m>���[����;��>8��>���>�f>�V>�0*>����K&��ח��`���~:�����A��f���{�d���
�����R�¾���|����F�������<��RP>mB^?t�I?�k?0��>�A ���=��
�(M2=����\ӿ=�)H>=�2?��9?gB?�X�=���	kg�6���Y���Bv�bL�>^W9>Y7�>S��>Cn�>�$����^>�R�>���>$>�A>�p�<�g=�}}> ��>ۓ??ĥ>��>+��Ǣ���T��L�b��`�=M=���?�]��hC��^������A�b��>:�3?�^�=	v���bʿ�ÿ��J?HF��K�;�Ŗ��5B>G�?�A+?0u>�$i��'��C��+�£{��,W>��$�1L��f:���[=_3'?ڶe>�4~>0�.�H 9�c@Q��L��Z�k>�2?����B�NAr�_�G���ݾ�?>\y�>�ܨ�.���Ŗ��u���d�?�t=r�8?ƭ ?�q��9>���4y�?d��a)H>8R_>��"=ĕ�=K^>1@��x�˽'
?�\�)=���=��S>��?]�->�ު=#s�>i����h��j�>��.>�3>�B?�|%?f�5�7Q��8�����!�坂>c�>kZp>��>q�E�P��=y7�>�[>B4�bIG����S���L>'��sR�r�}��=�Z�����=S�}=���*$>��Q=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ3T�>����T��q
���u�#=���> FH?�s���Q��=�ko
?t?�B򾝩����ȿ�qv����>h��?���?X�m�5A���@�8q�>���?RcY?�_i>T�۾֜Z�$|�>"�@?=�Q?��>46��s'���?+Ӷ?x��?��<>U��?/k?��>�ӓ�@�ZZ��u����D=�����0
>�TP<$��KT6�BI9��~���\�C�\���h=*z�;���>��<ʘ��g=�� <��m�O=���>xkb>ڋ�>��>k�'?�>A��>w�#>$�J���r���Z�K?+��?���in�/)�<�7�=��^��?,54?az_�E�Ͼޭ�>�\?沀?@�Z?>X�>*���?���俿Cl��85�<U�K>�&�>FY�>����VK>�Ծ&�C����>���>墣�I"ھ&�� 䪻�A�>�g!?9��>�]�=ҙ ?��#?��j>�(�>EaE��9��M�E�z��>Ţ�>�H?��~?��?�Թ�lZ3�����桿��[��:N>��x?V?�ʕ>Q���􃝿�kE�BI�3���T��?�tg?�S�/?82�?�??<�A?	*f>���Gؾ������>K!?o?
�{�?���&�ӭ�p:	?�b?Oo�>�Ɣ��ݽ�Tϼ��z�����?X\?E�$?j����`���ľ�h�<U�5�)�S����;J2���>��>l�����=��>�1�=�	m�.�i�<�X�=���>T>�=q�2���<,?�G�ك�U�=��r�ZvD��>�HL>f�����^?�u=���{�:���w���T� �?��?l�?	��^�h��"=?��?.	?�+�>;O��|޾o���Pw��sx��x���>��>�k�h�Q��������D��)�Ž���D?�#>>Y�>��> �>Ձ�>��O��(�Z�¾ �ݾ�[Y�f��X%�f'�?
,��Wʾ�-��8]=I������>{飽�0�>A?�0M>D>�> �?��=�oG>&�g>	�F>j1�>Dh�>y�v>J�=>Ԗû��ϽhKR?=���;'����&���g3B?Oqd?u0�>ci�򉅿����?���?�r�?�;v>�~h��,+�7n?�>�> �� q
?�T:=���@�<'U����4�������>�F׽k :��M��lf��j
?y/?g
�� �̾�9׽9���/o=hI�?��(?��)���Q�a�o�˷W��	S�����Wh��y����$���p��䏿�^�������(��*=��*?��?S|�1�%���"k�?�jf>x��>��>�>v�I>��	�Ϻ1���]�jA'���f7�>�F{?�~k>�C?��:?p=?T�e?�6�>�>�,վ3�*?�2=����t�?K��>��?|t&?n5?�B1?���>�*=��޾w����D?�2�>��?0��>��?�P��]e���$�=={Ҽ<F��ei���-E> �ֽ�k���U��ƽ�9�=Χ?���x>�?�� u>h};?�U�>�-�>+���6�k����<��><�?��>7 ���s�rQ�]a�>��?$�&���=a7S>�
�=ϔ	��:c<�g�= f�ե�=#H2���A�?= w�==��=�̔<�.+<䰿<r�U;�ɜ<u�><�?���>�C�>�@��� �����e�=?Y>S>>�Eپ�}���$��~�g��]y>�w�?�z�?�f=��=��=}���U��������K��<Σ?J#?XT?W��?v�=?:j#?ҵ>�*�pM���^�������?\!,?��>���L�ʾ���3�s�?v[?~<a����3;)�Ȑ¾H�Խ)�>�[/�t/~�����D�G텻����~����?���?�A� �6��x辩����[��`�C?R"�>Y�>��>�)��g�%��1;>
��>�R?k�>EhZ?��o?.\i?���>��A�f���sƚ��;@y�>�_C?�ob?�ݓ?��l?'��>g>΀I���辠��)(������,���=�5>ر�>�9�>D�>�>i���\�9���q$>��l>��>�s�>�M�>i?�>5��=�V?e?�>�鱾ew	�Qwg�������i?B͞?�\?7���+ƾ����I>�%�?���?�~?�齽��>j�v=L��~��T��>�=�>�3�>�$`����=�
�>!�Y>Q��>��p����ڱS�`�O��B?�8;?�>�ÿ�gk�飯��1=a<���̓x��$�=ď���Od>Ԅ�=;���w����|�/�־�Њ��/���u�mL����?B��=�<��=>·��]0�hz}=��Z>HqD���{=��.>,�w=%�g�>�[J������H�;��=>�y
���Ǿ�tz?�7I?�+?��E?A`j>�!>�e����>��+���?.�c>�^O��軾75�����e���پ5Ӿ�_��蛾�(>��Q��>LgA>y��=���;�.�=�T=:�=�A�;l�9=���=4͹=��=ܾ=��>�>'t?c�����:�N�w
�@�@?���>ͣ�=
ھU�2?�3D>�����)�����m,{?�[�?��?} ?����)��>e������F�<�,g��Ui>�	�=�S/�￼>��h>����v���M���[�?��@�@9?�׊��8ο3e
>4s7>$&7>b�6��-9���}���	��5��w]?�:4���޾�>�_=�ZԾU�j��=|�>��~<�<6���c����=�l��A�,=�c=Bg�>$�h>�r=+C���N=Un�=�T�=�9>�(�='R���3���a�=\U�=Y{�>i�=. ?<�?��,?}�y?��>du���w �{�����>k>��>�M�=^9?k�>Ah+?�]?/�-?�E�>,
X=i0�>���=�3�@�~����o��`Ѿ�N�?���?.ׇ>!Kz��/��C��^�;����S�>�D�?��?��>w��X]��	�Du.�j����=�X>&�L���`��R�����{������4��>�v�>z�>� >���=�q@>���>C >?�=�<���;���=Sm�Q�(=)��<p�;��n���Ҽ_���刽�	�!>��/��z�<�jP�-�=���>��>O��>ۈ�=�Ⲿ�r/>����o�L��q�=�
���B�H�c��}��l/��9:��?>
eV>f&����o�?GW>��?>��?#Eu?'>&��&Ӿ� Hg���R�P�=�,>��7�-:���_��7N�6ҾQ��>�"�>��=0P�q�!�P� ��=�'����S�d�>�0��������K����䫿0t��n�=�yK?.Ћ��%�>.[8?�E?�?�?i�?rT��������> �t��U��[��ӻ��VK�=_�/?R�S?P��>�s$�-5���̾H���Q�>��G���O�/����S0������F�>z���!Ѿ�3�9H��2����vB���q����>�_O?[�?ֵa�/����N�o��G��+h?�ng?6�>�i?5t?"7��9:�=��iU�=o�n?>��?�?��
>G;�=}h��JW�>i�?�"�?y�?��p?�>�Z.�>@��;k	>��T��R�=>���=,��=�
?�T
?S�?5؛��z�Qu�p�뾿?Z�ˎ�<p�=��>�'�>M�y>%n�=�[=3#�=�T>Q�> Ύ>��g>�P�>��>��������$?�&L����=�c?eyk>��>ۧ����A=x��&�Ž��4�]=��pr�;�
��#�=^�=�f�>��ֿ�7�?;�
>�3@���?N;ھ�>��&�>��=B*�g��>>>�]>���>oY�>�x=��>p�;-�Ծ��>���x\�!�C�m&S��ξ�Ҁ>ܞ��@(�l��Խ����J�Rڰ����<^i��j��;�y��<���?�����nk��w)�����1	?Y�>2�6?����Mޤ�Mg>+�>���>r���-������E⾌��?j��?�?c>3�>ҽW?^�?�2���2�"QZ���u�WA��e���`�{ލ�����q
��f��Ņ_?�x?�/A?U�<rz>i��?|�%�q����(�>b /��8;���;=w.�>�5��[�`�o�ӾH�þ��E�F>�^o?}�?}?�V��2����=��5?��?�9�?��8>Em@?�'����?̳>�>�FI?!k>n?s�>>l�>�VU>+�T<3WE>��V�F���T�.��ue������WR�a"Q�I�B=�{�=Ӊ���<���=�>��6�k<uJ�=���GH�<a�=�@>To�>�^?l��>`g:>>�8?P����?;�U2 ��f[?���>]��,I�=��V�ѻ�+�r>�gh?i��?��R?5?,�M��1��i�=��=�� <�=>���>��8B��k�p9f>P�>S2e��.�z� ��t��e�g���gL	>Z��>y�|>�����(>�I���Bz�sid>��Q�y���
NT�t�G�D�1��
v�7�>N�K?�?���=��-���:f�R!)?�U<?�=M?��?�#�=߸۾Y�9��J����ϟ>�T�<	������ ����:�%̟: �s>��w�#S>+��q׾to�T?��&׾�م=Hq�����=���޾'M��/o=s6�==���Z �V$�����3�S?k��<s�Ծ)\���ר��O>̷�>::�>�{��A��ݿA��Ѿ�]=��>��z>�ч����}S�S��r�>�O<?ya?Īu?8e���};���T�s��������{�o� ?]�J>� #?&��=|i>Ϡ�����c�%XN�Ʈq>�e?Q���J0�/:�=wj�tb��{>��?t؁=��X>�sa?�'
?�mY?���>�g�>��>���<jľ�&?\x�?���=�ҽ��Q��F9�O|F����>�)?�vC�:��>��?}�?KO&?Q?��?�>� ��@�h�>�5�>�hX��篿��a>�I?���>ǋW?��?�$?>�>6��a秽=<�=i�>0�1?^^#?z�?��>IY�>�ޠ�9�=�]�>c�b?V��?��o?�O�=;?b5>nv�>ҡ�=�>�!�>��?�?O?hds?.J?hf�>x�<�������o�)c�0/C;�sT<��{=v��?�q�
���<hV�;r�����~�-�PD�RG���l�;W�>nt>�ԕ�|\1>�cľp��X@>��������);����=�À>��?���>L�"�S��=���>z��>���M+(?�?M(?�i;b�b�)Aھ�K�lN�>��A?b�=�l��e����u���f=�m?r^?�>W��%����b?��]?^g�X=���þ��b���)�O?�
?J�G���>f�~?��q?���>�e��9n�"���Cb�K�j�/ζ=�r�>�X���d��@�>ƛ7?�O�>��b>�)�=u۾j�w��p��5?��?��?j��?�+*>��n�
4��ľ����L?�q�>���a?͗�=}L��	���	������9����Ǿ�Ko��žO?W��W��1U����=R�?�hP?��;?Э�?���d�h�+�K������Z�� ��oO��>��b�:+�G7Q��q1�먾ˑ�w,�������F?��|�?jp(?3	1�w�>Z���f��Z�Ⱦ�\I>�ȝ�<��@�{=�����dy=6�h=Y�f��3�����?_��>ae�>�0<?>[��<��m/�yM7�]P��]2>�d�>��>���> A�:؂4�<����Ǿ1��;tӽg��>�R?�_g?q�[?B�̾�q��8}����'����̃��f�>V%?��	?���|D=Z��5�H�D8d��+#��h��O��h �=��?���>ȝ>�	i?�E?����p��C"��t�+�v�4>Q>�L?��$?B*t=r��ҋ	�C��>׹l?�N�>0t�>�~���8!��{��vʽ���>�ڭ>č�>$�o>�-�H�[�Fe��R����"9����=��h?cӄ�Z�`���>��Q?�w�:�U<���>�v��!������'�=*>�?��=tT<>�žB%�S{��9����%?P�?�ۉ���(����>��?���>b��>=��?���>r�ľX�f;�?R�Z?�+J?�A?�5�>��=k┽�Խ�(��?/=��>97R>!�r=@|�=![��"e���%�>�T=/ܸ=�Tּ�	Ľ�\<������;���<�++>|�ڿOY�S�ž��þ�cپ �	��V]���_���˾����܅��Ӿ;T��C�_
���]�o���z��ܩ�\��?'��?/?���������h�FrھL��>0��GT^�i����� ����3־ob��hi�x3��
E���h�{I?����ڿ���3[u��8?:�?���?\L�^�I�C���W'>�k�>��>Z߶��u��^�ҿ9G�cP?%.?����ͷ�=��>V�R=k�@>�i�>�@��g$���Z��2?t&�?�?����{���	@¿Ċ=l��?��@}A?�(����x�U=���>H�	?P~?>Pk1��0� 谾�=�>�<�?���?�TM=��W��\	�{}e?f`<��F��E�U(�=9ۤ=�=>���J>�y�>ٖ�^A� ~ܽ�|4>�م>&�"�o��%R^�lY�<]�]>�vս�R��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=w6�����{���&V�}��=[��>c�>,������O��I��U��=�P�nNſ�g�d����.=�5��V�^�ҽ{���z}�xZ���,���,�ݠ�=@ϟ=&E>f�[>F�Q>��>;c?�y?t��>}?1>P������.�U��"����C�H�\�������{\о��I��$��}��˾�4��5��%�H�D�n��(���\��H5��'?uj�������8&���,���þ������-�����/������^��#=�?�3 ?�ߊ���m�y��b+�=^F��*�E?��R�.�4駾�g�=���Lý���>f�&>'8ľ��S�oQi�6?��&?�V̾U�U�J�;>���8C��s{�>b?�@5�K� >��T?P(��sU�d#�>U?�>e+?�?�O�>�i��!�5�h�?t'r?t}0=+���B?,�9�z���f�25�P���sV��B>��t>+d��Kp��<Y�ѽ��W?-ߐ>7^)����aH�������<�zt?�8	?:�>�i?֒D?V�<�����T�"���_�=R�U?"�i?L�>S�y�2Ӿ������3?	f?�zS>V�s����r�,�h��2*?�o?��?���=���������q�4?S�v?��^��v��4$�$T_�w�>Gr�>���>�;���>z�A?�&�wD��� ���7�|2�? g@��?<�i<(9��=}*?��>EO��yɾ�Ľ���k o=@��>訾Kw�xI ���,��:7?<�?f��>mw������5>y����?��?�;=G���x������VC�7w�����K��!ܾ�94�����V�þ�(��!o>HL@}��7�>�ۄ�7w�mÿ#�{����!�T�,�?_�>�9�vG���![�����$�%=H�������>m��=�+�h䑾i8{�i�0����.y�>�ý�M7>�A���ž�î�8��?��>x��>�g>e������?����G^ҿm���K��^C^?�ٝ?��?��?A:���4���衾��ＯO?�zy?�[P?����I��z%C���~?A+��7��boa�F�g�~�G>0�X?�C?�?\�
�:���?HR?)X�>}0���ƿ�����Q���?��?���n�?ʒ�?�0?\�%�/u���+��;&��n��RF�?g��>����-��sd��R��?��v?�Sc�7t��_?��a���p��-���ƽ�ݡ>��0��`\��g����0Xe����By���?j]�?��?��=#��3%?��>ѝ���;Ǿ���<̓�>�(�>�'N>�(_���u>r���:��j	>ɯ�?�~�?�i?��������;X>!�}?�ʴ><��?_	�=���>�A�=0W������A�">�5�=��F��� ?�L?o�>���=��<�KB0��:G�c-O�����C�ل>�\`?o�K?Ŕi>J}����&�p,�c\½�<6��	���<������ҽq�;>4�E>�>>��7��oӾd�?�y���ؿ�k����'�=4?�ʃ>�?�����t�Ţ��G_?ߎ�>�+�X'���(���Y����?F�?��?
�׾�˼�>�ŭ>�=�>��Խ0��������7>s�B?���B����o���>��?��@<Ϯ?�h��	?���P��Ua~����7�a��=��7?�0��z>���>��=�nv�޻��W�s����>�B�?�{�?��>!�l?��o�P�B���1=8M�>͜k?�s?Po���c�B>��?"������L��f?�
@u@`�^?*mֿ@����q��?*�� L�=��=��2>�cٽ�]�=�6:=�
E�Ͳ��d�=��>W[e>��p>R%O>Q�;>��(>p�����!����KR��S�C�?�v�>�Z����Ou�x�j%�������a��u#��UΣ�N0P��&�B�b����=�4f?�<?��y?>X<?/X���>�$	�S>�m�
Do�ݱq>��L?�W?�8?��>]����H�,��z�����J��>�9>6��>pF�>�.�>���V+Z=X�}>Qb�>W��z����>��νaP�>��>@��>���>�]>s8�ڔ�������W�K���T@;Y�?|�;_]b�׉�զ���ؾ-��>��?O�=cԿ�����Gn?p��ۦH�z����>+�/?u�;?�!�>�0�L��<�,a= 0�����/r�>r�缱�y�u�1��K/>��N?:�f>�u>�x3�wK8���P������|>,6?cȶ���8��u���H��tݾ�SM>H�>��@��\�#�����~���i�e�{=q:?��?V����󰾷�u�zC��vR>�-\>��=oa�=�DM>U c�x�ƽ�H�.=���=��^>X�?->��=Ҟ�>f���guY��>�3>�3>R�@?�"?9���q���_������}>���>f�x>s
>�,M�ս�=it�>"�a>yc�p3����
���C�A�L>�Ek��M���Y��?n=���A�= ��=e���&3�O�,=%�~?�����舿)�
f��SqD?�,?���=_*E<I�"�a���s��S�?��@g�?�	�d�V���?�A�?;��}��=��>�̫>@ξ�L���?��ŽyԢ�~�	�;�"�U�?��?��0��ɋ��"l�
�>\j%?֎Ӿ�g�>$w�iZ�������u���#=	��>�8H?+V��ƿO��>��v
?V?m^�Ω����ȿT|v����>$�?��?�m�
A��?@���>��?�gY?Goi>+g۾�aZ���>��@?	R?��>9��'��?�޶?���?�i>��?�Jb?�?����<g�+���K���/=�Z��B��>-a=��ϾJ	��胿	W��į:���8��
�=��0<l�>�g5=�q�b&�=T��r;����;w�>> >��>L��>��4?�j^>,ٟ>�>a���I:�T���QuK?��?�+��l� ��<��=�Z`���?�4?�s��VSѾ���>�]]?.q�?]�Z?��>�3��Қ�&׿��˴�M��<E�F>���>��>F�����N>{7׾�>��q�>Z��>�T��	�پ'B��t��a�>�!?��>��=o� ?c�#?��j>�*�>�aE�{9���E����>L��><H?��~?v�?Bع�JY3����6硿ܑ[��5N>��x?�T?�̕>t��������gE�>I�o���ɛ�?�tg?�T�Y?�1�?k�??h�A?�(f>����ؾ�����>(�!?��o�A�vJ&�A��S{?Q?���>�	��X�ս?�ּ1��|���
�?5*\?+B&?ҙ��,a�?�¾�<�a#���T�̶�;�E� �>�>����Ff�=C>��=�Jm�G6��f<�l�=�|�>+��=m07�[���<�0?
i������i�=��e�Օ�>қ>s�l?��=�|����e��u�ؾ&�]?'�?O��?�H:�ax�߼`?�?�6
?r ?������л��㎝��v��6�� �=!?>�}X�bǧ��$���`��}����<b�,��VL ?�%�>�V�>u��>N>>��>�,V�C���������f�7����M��
3�$2��ݾ.����F�=��炇����>�ֹ<�.�>�?�A�>��>Y�>�!��mC>��V>K��>�^�>!�>���>V8�=��=T;��JR?"�����'�2��A���d3B?�qd?2�>)i�ɉ�������?���?er�?
9v>�~h�[-+�&o?�>�>���vo
?ic:=����3�<qS����H7���E��>�F׽p:��M��lf�_i
?M/?�卼r�̾.@׽e��,\=_Q�?��8?��3�:�L�Ԍ^�X�]���P�>�P�Pq{�A���b�9��c����X���,�~��P0�f��<\�!?mC�?v����0޾�g��"�n�{�=�ld>?��>���>
��>8Q2>���7� �6�W�9�.��W����>��k?�rj>�L?��?��I?Wi?�0�=,��>\�����?�?f=�ǽ�#�>"��>ŷ?q�S?Hi:?�WC?#6�>o,>�
)�m���k�0? �>ؐ	?�ɡ>J=�>"���!�A#w>Ȭ��di��j�IGB>�F��mwK����q���"|>��?���RZ8������"m>�`7?9�>���>�������W��<4h�>�+
?u��>d��� �r����&�>ӂ�?�G�$��<w3.>�2�=6������:Xp�=x��T2�=�r���j<�}<��=X��=[TP9%1�;R�';��<�]�<�y�>��?֐�>�8�>�>��Ϊ �ǽ��b�=�-Y>�(S>�>8پY|��$��M�g��yy>�x�?�v�?��f=p&�=��=����F]��G����j��<l�?�J#?�YT?.��?�=?�m#?׮>7.��M��_[�����?>!,?#��>�����ʾ�񨿈�3��?N[?N<a�����;)�y�¾��Խֱ>�[/��/~�����D��ͅ����&����?Ϳ�?�A���6�Mx辜����[���C?�!�>�X�>�>��)���g�%��1;> ��>R?>��>�M?��|?��Z?��'>Ħ)����Jr���܏��t>��B?_�t?�ɐ?��c?��>��>��G��K�q� �(�2�K�0����i=�Cf>���>w��>�X�>���=y�轚Wؽ�P����=p�V>��>���>5"�>�j>��o<�O?�f�>����X��ޔ�yꚾ����r�Y?��?w4?�d�=�¾mt8����Jx>���?rH�?��?`�n�+#>�,=�1����)z�>���>��C>^��	>���>�H>D��>K�=!��/�J�D�J��\?_�O?<%>e�ο�M��(\��G𕽒Yc=T�3ԍ���Ҿ� >�P���Ĉ�����z��F&���Z�xҮ��8ɽ3����?9vʽܭ���^�>)=a����W�r(S=�v��� >�)��<C���Y<���=�x= �(�ę!;���=����A�ʾ*�o?��W?�;?�`B?�k�>Ԅ@>�#>��3�>4�=���>�}�>Q��h�?����h��}���Ц�]"K� �ʾ��>ңb���=/u>R�0>��۳5=k��<��P='P=c�-;VE~=���=Y��<OG>�	,>��/<�6w?Z�������4Q��Z罣�:?�8�>{{�=��ƾQ@?w�>>�2������wb��-?|��?�T�?&�?�ti��d�>O��~䎽q�=����!>2>���=T�2�^��>��J>���K��H����4�?��@��??�ዿϢϿAa/>�7>Z0>��R��1�U�\�*�b�:TZ���!?TC;��>̾E/�>"�=,߾[�ƾ�B.=�f6>0�a=�Y�JJ\�y��=�{�0J<=�Kl=$ۉ>D>���=���!�=U(I=]��=��O>Jˑ��7��+��4=���=��b>>�%>�u�>!�?�8?�I?Nl�>��9��g��ٚx�M�>ў�=!V?��=���=��>,�?I<o?�L?k�>�k=t�?⭱=C4�FŅ��#�$�ƾw�;简?�՝?�:�>9�>��<i�4��V�T�轚�4?p!E?�O�>��?�"�zd����|+�����d�Ľ?��=��A�?;����C=H������/=�r�>���>���>N��>��=G�=��>���='�Ľ��<?l!�i��=�����=m�^=��=��;r��E̹-�$�i�;�l<rs�� �<��=��>���>������&>�@ۺ���%�/>l�6��E�b8a>3�o�n�B�<Lw�m[���dP��H��a�=i]>n��={���T�?bqm>]�=���?9�{?чr>�_V�i���������ƾ���`�<<�>��*��C'���z�8'C�����x�>>�L�>PVK>�a)���?�A�=4�ؾsm3�Ia�>i����=���*��q���������Kxh���:9VE?"��`��=�B{?tqD?R��?��>2�[��n׾�I>�ʆ��~U<�;�lFe�0
B�(@?�#?�H�>�3较A�9J̾� ���ܷ>�9I���O�v�X�0���=з�u��>p��� �оM#3��f������	�B�=Mr�b��>D�O?�?T:b��W��kUO����"���p?�{g?��>/G?�??g��Jz�v��1l�=��n?��?;�?��
>�Ic=ۿ����>bC�>Mё?^�?etn?�m����>8�=�=��A��j$=��=r%>9�>	?���>�� ?'�̽.>�PCھ�c���!|�������=��>ֵV>=�V>c8>zX���}�<D�>��>K��>�y`>X9�>p.m>:���J�ɾmE?��%<S�>�NE?8N�>��>�ޤ��m%�f
�X�ͽ�=��������������:>1�=P��>p˿ᄎ?�k�>&9�ǜ#?
�ξU���e��=Vy,=v?½���>��=5�b>�ܖ>���>x�*>s^2>,��=s/Ӿ�K>����i!�� C��qR�8�Ѿ��z>{���W*&����& ��/.I�	;���a��j��/��AC=�_ݼ<�K�?	����k�o�)��f����?�K�>-"6?<Ō�&��p�>��>��><�������ƍ�r���?���?<c>��>t�W?�?��1�G3�	rZ�V�u��'A��e���`�����������
�2��>�_?�x?�sA?f8�<�5z>��?��%�?Џ��#�>K /��&;�,C<=-�>7(���`��Ӿb�þ�-�UDF>��o?�$�?,W?*WV��ʽ��!>�KJ?�{*?ד`?.�?�.??� E�ck&?��>�`�>��>[�?R�?�R'?
Pq>Ɉ�=�)��a[w=������q��9���WD��p����<�=6��bwf��(-=�'�=�����t��� =�����A<�(=6n�=��=�ƃ>��^?��>恝�'�5?�;���)�����n?rm?�c������U����6�.>I�Y?.&�?/*?ù ?������&�>̨=�4>W��=S��>x�>[�>���n�$�f����=Ǳ�=P\->K+5� �/��?��k�����̕�<?��>-�}>����~*>W'��f�|�v�c>�]P�����T�,�G���0��Es�h�>4L?�?�ؘ=�v�v����.f�WO)?�l;?��L?Z�?:�=`ھl:�ǟI�T}�7�>��<�	�U���L�����:��ր���s>�P��w�#S>+��q׾to�T?��&׾�م=Hq�����=���޾'M��/o=s6�==���Z �V$�����3�S?k��<s�Ծ)\���ר��O>̷�>::�>�{��A��ݿA��Ѿ�]=��>��z>�ч����}S�S��r�>�O<?ya?Īu?8e���};���T�s��������{�o� ?]�J>� #?&��=|i>Ϡ�����c�%XN�Ʈq>�e?Q���J0�/:�=wj�tb��{>��?t؁=��X>�sa?�'
?�mY?���>�g�>��>���<jľ�&?\x�?���=�ҽ��Q��F9�O|F����>�)?�vC�:��>��?}�?KO&?Q?��?�>� ��@�h�>�5�>�hX��篿��a>�I?���>ǋW?��?�$?>�>6��a秽=<�=i�>0�1?^^#?z�?��>IY�>�ޠ�9�=�]�>c�b?V��?��o?�O�=;?b5>nv�>ҡ�=�>�!�>��?�?O?hds?.J?hf�>x�<�������o�)c�0/C;�sT<��{=v��?�q�
���<hV�;r�����~�-�PD�RG���l�;W�>nt>�ԕ�|\1>�cľp��X@>��������);����=�À>��?���>L�"�S��=���>z��>���M+(?�?M(?�i;b�b�)Aھ�K�lN�>��A?b�=�l��e����u���f=�m?r^?�>W��%����b?��]?^g�X=���þ��b���)�O?�
?J�G���>f�~?��q?���>�e��9n�"���Cb�K�j�/ζ=�r�>�X���d��@�>ƛ7?�O�>��b>�)�=u۾j�w��p��5?��?��?j��?�+*>��n�
4��ľ����L?�q�>���a?͗�=}L��	���	������9����Ǿ�Ko��žO?W��W��1U����=R�?�hP?��;?Э�?���d�h�+�K������Z�� ��oO��>��b�:+�G7Q��q1�먾ˑ�w,�������F?��|�?jp(?3	1�w�>Z���f��Z�Ⱦ�\I>�ȝ�<��@�{=�����dy=6�h=Y�f��3�����?_��>ae�>�0<?>[��<��m/�yM7�]P��]2>�d�>��>���> A�:؂4�<����Ǿ1��;tӽg��>�R?�_g?q�[?B�̾�q��8}����'����̃��f�>V%?��	?���|D=Z��5�H�D8d��+#��h��O��h �=��?���>ȝ>�	i?�E?����p��C"��t�+�v�4>Q>�L?��$?B*t=r��ҋ	�C��>׹l?�N�>0t�>�~���8!��{��vʽ���>�ڭ>č�>$�o>�-�H�[�Fe��R����"9����=��h?cӄ�Z�`���>��Q?�w�:�U<���>�v��!������'�=*>�?��=tT<>�žB%�S{��9����%?P�?�ۉ���(����>��?���>b��>=��?���>r�ľX�f;�?R�Z?�+J?�A?�5�>��=k┽�Խ�(��?/=��>97R>!�r=@|�=![��"e���%�>�T=/ܸ=�Tּ�	Ľ�\<������;���<�++>|�ڿOY�S�ž��þ�cپ �	��V]���_���˾����܅��Ӿ;T��C�_
���]�o���z��ܩ�\��?'��?/?���������h�FrھL��>0��GT^�i����� ����3־ob��hi�x3��
E���h�{I?����ڿ���3[u��8?:�?���?\L�^�I�C���W'>�k�>��>Z߶��u��^�ҿ9G�cP?%.?����ͷ�=��>V�R=k�@>�i�>�@��g$���Z��2?t&�?�?����{���	@¿Ċ=l��?��@}A?�(����x�U=���>H�	?P~?>Pk1��0� 谾�=�>�<�?���?�TM=��W��\	�{}e?f`<��F��E�U(�=9ۤ=�=>���J>�y�>ٖ�^A� ~ܽ�|4>�م>&�"�o��%R^�lY�<]�]>�vս�R��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=w6�����{���&V�}��=[��>c�>,������O��I��U��=�P�nNſ�g�d����.=�5��V�^�ҽ{���z}�xZ���,���,�ݠ�=@ϟ=&E>f�[>F�Q>��>;c?�y?t��>}?1>P������.�U��"����C�H�\�������{\о��I��$��}��˾�4��5��%�H�D�n��(���\��H5��'?uj�������8&���,���þ������-�����/������^��#=�?�3 ?�ߊ���m�y��b+�=^F��*�E?��R�.�4駾�g�=���Lý���>f�&>'8ľ��S�oQi�6?��&?�V̾U�U�J�;>���8C��s{�>b?�@5�K� >��T?P(��sU�d#�>U?�>e+?�?�O�>�i��!�5�h�?t'r?t}0=+���B?,�9�z���f�25�P���sV��B>��t>+d��Kp��<Y�ѽ��W?-ߐ>7^)����aH�������<�zt?�8	?:�>�i?֒D?V�<�����T�"���_�=R�U?"�i?L�>S�y�2Ӿ������3?	f?�zS>V�s����r�,�h��2*?�o?��?���=���������q�4?S�v?��^��v��4$�$T_�w�>Gr�>���>�;���>z�A?�&�wD��� ���7�|2�? g@��?<�i<(9��=}*?��>EO��yɾ�Ľ���k o=@��>訾Kw�xI ���,��:7?<�?f��>mw������5>y����?��?�;=G���x������VC�7w�����K��!ܾ�94�����V�þ�(��!o>HL@}��7�>�ۄ�7w�mÿ#�{����!�T�,�?_�>�9�vG���![�����$�%=H�������>m��=�+�h䑾i8{�i�0����.y�>�ý�M7>�A���ž�î�8��?��>x��>�g>e������?����G^ҿm���K��^C^?�ٝ?��?��?A:���4���衾��ＯO?�zy?�[P?����I��z%C���~?A+��7��boa�F�g�~�G>0�X?�C?�?\�
�:���?HR?)X�>}0���ƿ�����Q���?��?���n�?ʒ�?�0?\�%�/u���+��;&��n��RF�?g��>����-��sd��R��?��v?�Sc�7t��_?��a���p��-���ƽ�ݡ>��0��`\��g����0Xe����By���?j]�?��?��=#��3%?��>ѝ���;Ǿ���<̓�>�(�>�'N>�(_���u>r���:��j	>ɯ�?�~�?�i?��������;X>!�}?�ʴ><��?_	�=���>�A�=0W������A�">�5�=��F��� ?�L?o�>���=��<�KB0��:G�c-O�����C�ل>�\`?o�K?Ŕi>J}����&�p,�c\½�<6��	���<������ҽq�;>4�E>�>>��7��oӾd�?�y���ؿ�k����'�=4?�ʃ>�?�����t�Ţ��G_?ߎ�>�+�X'���(���Y����?F�?��?
�׾�˼�>�ŭ>�=�>��Խ0��������7>s�B?���B����o���>��?��@<Ϯ?�h��	?���P��Ua~����7�a��=��7?�0��z>���>��=�nv�޻��W�s����>�B�?�{�?��>!�l?��o�P�B���1=8M�>͜k?�s?Po���c�B>��?"������L��f?�
@u@`�^?*mֿ@����q��?*�� L�=��=��2>�cٽ�]�=�6:=�
E�Ͳ��d�=��>W[e>��p>R%O>Q�;>��(>p�����!����KR��S�C�?�v�>�Z����Ou�x�j%�������a��u#��UΣ�N0P��&�B�b����=�4f?�<?��y?>X<?/X���>�$	�S>�m�
Do�ݱq>��L?�W?�8?��>]����H�,��z�����J��>�9>6��>pF�>�.�>���V+Z=X�}>Qb�>W��z����>��νaP�>��>@��>���>�]>s8�ڔ�������W�K���T@;Y�?|�;_]b�׉�զ���ؾ-��>��?O�=cԿ�����Gn?p��ۦH�z����>+�/?u�;?�!�>�0�L��<�,a= 0�����/r�>r�缱�y�u�1��K/>��N?:�f>�u>�x3�wK8���P������|>,6?cȶ���8��u���H��tݾ�SM>H�>��@��\�#�����~���i�e�{=q:?��?V����󰾷�u�zC��vR>�-\>��=oa�=�DM>U c�x�ƽ�H�.=���=��^>X�?->��=Ҟ�>f���guY��>�3>�3>R�@?�"?9���q���_������}>���>f�x>s
>�,M�ս�=it�>"�a>yc�p3����
���C�A�L>�Ek��M���Y��?n=���A�= ��=e���&3�O�,=%�~?�����舿)�
f��SqD?�,?���=_*E<I�"�a���s��S�?��@g�?�	�d�V���?�A�?;��}��=��>�̫>@ξ�L���?��ŽyԢ�~�	�;�"�U�?��?��0��ɋ��"l�
�>\j%?֎Ӿ�g�>$w�iZ�������u���#=	��>�8H?+V��ƿO��>��v
?V?m^�Ω����ȿT|v����>$�?��?�m�
A��?@���>��?�gY?Goi>+g۾�aZ���>��@?	R?��>9��'��?�޶?���?�i>��?�Jb?�?����<g�+���K���/=�Z��B��>-a=��ϾJ	��胿	W��į:���8��
�=��0<l�>�g5=�q�b&�=T��r;����;w�>> >��>L��>��4?�j^>,ٟ>�>a���I:�T���QuK?��?�+��l� ��<��=�Z`���?�4?�s��VSѾ���>�]]?.q�?]�Z?��>�3��Қ�&׿��˴�M��<E�F>���>��>F�����N>{7׾�>��q�>Z��>�T��	�پ'B��t��a�>�!?��>��=o� ?c�#?��j>�*�>�aE�{9���E����>L��><H?��~?v�?Bع�JY3����6硿ܑ[��5N>��x?�T?�̕>t��������gE�>I�o���ɛ�?�tg?�T�Y?�1�?k�??h�A?�(f>����ؾ�����>(�!?��o�A�vJ&�A��S{?Q?���>�	��X�ս?�ּ1��|���
�?5*\?+B&?ҙ��,a�?�¾�<�a#���T�̶�;�E� �>�>����Ff�=C>��=�Jm�G6��f<�l�=�|�>+��=m07�[���<�0?
i������i�=��e�Օ�>қ>s�l?��=�|����e��u�ؾ&�]?'�?O��?�H:�ax�߼`?�?�6
?r ?������л��㎝��v��6�� �=!?>�}X�bǧ��$���`��}����<b�,��VL ?�%�>�V�>u��>N>>��>�,V�C���������f�7����M��
3�$2��ݾ.����F�=��炇����>�ֹ<�.�>�?�A�>��>Y�>�!��mC>��V>K��>�^�>!�>���>V8�=��=T;��JR?"�����'�2��A���d3B?�qd?2�>)i�ɉ�������?���?er�?
9v>�~h�[-+�&o?�>�>���vo
?ic:=����3�<qS����H7���E��>�F׽p:��M��lf�_i
?M/?�卼r�̾.@׽e��,\=_Q�?��8?��3�:�L�Ԍ^�X�]���P�>�P�Pq{�A���b�9��c����X���,�~��P0�f��<\�!?mC�?v����0޾�g��"�n�{�=�ld>?��>���>
��>8Q2>���7� �6�W�9�.��W����>��k?�rj>�L?��?��I?Wi?�0�=,��>\�����?�?f=�ǽ�#�>"��>ŷ?q�S?Hi:?�WC?#6�>o,>�
)�m���k�0? �>ؐ	?�ɡ>J=�>"���!�A#w>Ȭ��di��j�IGB>�F��mwK����q���"|>��?���RZ8������"m>�`7?9�>���>�������W��<4h�>�+
?u��>d��� �r����&�>ӂ�?�G�$��<w3.>�2�=6������:Xp�=x��T2�=�r���j<�}<��=X��=[TP9%1�;R�';��<�]�<�y�>��?֐�>�8�>�>��Ϊ �ǽ��b�=�-Y>�(S>�>8پY|��$��M�g��yy>�x�?�v�?��f=p&�=��=����F]��G����j��<l�?�J#?�YT?.��?�=?�m#?׮>7.��M��_[�����?>!,?#��>�����ʾ�񨿈�3��?N[?N<a�����;)�y�¾��Խֱ>�[/��/~�����D��ͅ����&����?Ϳ�?�A���6�Mx辜����[���C?�!�>�X�>�>��)���g�%��1;> ��>R?>��>�M?��|?��Z?��'>Ħ)����Jr���܏��t>��B?_�t?�ɐ?��c?��>��>��G��K�q� �(�2�K�0����i=�Cf>���>w��>�X�>���=y�轚Wؽ�P����=p�V>��>���>5"�>�j>��o<�O?�f�>����X��ޔ�yꚾ����r�Y?��?w4?�d�=�¾mt8����Jx>���?rH�?��?`�n�+#>�,=�1����)z�>���>��C>^��	>���>�H>D��>K�=!��/�J�D�J��\?_�O?<%>e�ο�M��(\��G𕽒Yc=T�3ԍ���Ҿ� >�P���Ĉ�����z��F&���Z�xҮ��8ɽ3����?9vʽܭ���^�>)=a����W�r(S=�v��� >�)��<C���Y<���=�x= �(�ę!;���=����A�ʾ*�o?��W?�;?�`B?�k�>Ԅ@>�#>��3�>4�=���>�}�>Q��h�?����h��}���Ц�]"K� �ʾ��>ңb���=/u>R�0>��۳5=k��<��P='P=c�-;VE~=���=Y��<OG>�	,>��/<�6w?Z�������4Q��Z罣�:?�8�>{{�=��ƾQ@?w�>>�2������wb��-?|��?�T�?&�?�ti��d�>O��~䎽q�=����!>2>���=T�2�^��>��J>���K��H����4�?��@��??�ዿϢϿAa/>�7>Z0>��R��1�U�\�*�b�:TZ���!?TC;��>̾E/�>"�=,߾[�ƾ�B.=�f6>0�a=�Y�JJ\�y��=�{�0J<=�Kl=$ۉ>D>���=���!�=U(I=]��=��O>Jˑ��7��+��4=���=��b>>�%>�u�>!�?�8?�I?Nl�>��9��g��ٚx�M�>ў�=!V?��=���=��>,�?I<o?�L?k�>�k=t�?⭱=C4�FŅ��#�$�ƾw�;简?�՝?�:�>9�>��<i�4��V�T�轚�4?p!E?�O�>��?�"�zd����|+�����d�Ľ?��=��A�?;����C=H������/=�r�>���>���>N��>��=G�=��>���='�Ľ��<?l!�i��=�����=m�^=��=��;r��E̹-�$�i�;�l<rs�� �<��=��>���>������&>�@ۺ���%�/>l�6��E�b8a>3�o�n�B�<Lw�m[���dP��H��a�=i]>n��={���T�?bqm>]�=���?9�{?чr>�_V�i���������ƾ���`�<<�>��*��C'���z�8'C�����x�>>�L�>PVK>�a)���?�A�=4�ؾsm3�Ia�>i����=���*��q���������Kxh���:9VE?"��`��=�B{?tqD?R��?��>2�[��n׾�I>�ʆ��~U<�;�lFe�0
B�(@?�#?�H�>�3较A�9J̾� ���ܷ>�9I���O�v�X�0���=з�u��>p��� �оM#3��f������	�B�=Mr�b��>D�O?�?T:b��W��kUO����"���p?�{g?��>/G?�??g��Jz�v��1l�=��n?��?;�?��
>�Ic=ۿ����>bC�>Mё?^�?etn?�m����>8�=�=��A��j$=��=r%>9�>	?���>�� ?'�̽.>�PCھ�c���!|�������=��>ֵV>=�V>c8>zX���}�<D�>��>K��>�y`>X9�>p.m>:���J�ɾmE?��%<S�>�NE?8N�>��>�ޤ��m%�f
�X�ͽ�=��������������:>1�=P��>p˿ᄎ?�k�>&9�ǜ#?
�ξU���e��=Vy,=v?½���>��=5�b>�ܖ>���>x�*>s^2>,��=s/Ӿ�K>����i!�� C��qR�8�Ѿ��z>{���W*&����& ��/.I�	;���a��j��/��AC=�_ݼ<�K�?	����k�o�)��f����?�K�>-"6?<Ō�&��p�>��>��><�������ƍ�r���?���?<c>��>t�W?�?��1�G3�	rZ�V�u��'A��e���`�����������
�2��>�_?�x?�sA?f8�<�5z>��?��%�?Џ��#�>K /��&;�,C<=-�>7(���`��Ӿb�þ�-�UDF>��o?�$�?,W?*WV��ʽ��!>�KJ?�{*?ד`?.�?�.??� E�ck&?��>�`�>��>[�?R�?�R'?
Pq>Ɉ�=�)��a[w=������q��9���WD��p����<�=6��bwf��(-=�'�=�����t��� =�����A<�(=6n�=��=�ƃ>��^?��>恝�'�5?�;���)�����n?rm?�c������U����6�.>I�Y?.&�?/*?ù ?������&�>̨=�4>W��=S��>x�>[�>���n�$�f����=Ǳ�=P\->K+5� �/��?��k�����̕�<?��>-�}>����~*>W'��f�|�v�c>�]P�����T�,�G���0��Es�h�>4L?�?�ؘ=�v�v����.f�WO)?�l;?��L?Z�?:�=`ھl:�ǟI�T}�7�>��<�	�U���L�����:��ր���s>�P��R����8`>�����ݾ�-n��J��N羀�P=���k�N=,���վ��~��,�=�I>���^� ��ݖ�uિ��J?Egf=�Z��'SV�@빾T>W�>DP�>z�=��Iw��`@�𓬾 ;�=L4�>�:>A풼S��ޓG����rts>��@?M�]?�z?PK�QL���G�D�Ⱦ.����-%��"?%��=+�(?��7>*�n=-���N���7^�/J��k�>��>����L4��ڝ���s��	��>��>�Dz>Y	?�P?���>�;W?c<?`�?�e�>7r�<U����&?x"�?��={6ս��T�g+9�z�H�M,�>��)?O|8�˻�>��?(�?܋#?|Q?�@?��>?I �D�?��U�>Wc�>sY�x���=\>��F?ǝ�>I
W?ze�?cRE>�5�ț�Ť��Z��=�>��2?��%?�#?���>��> ��C>�=m��>�i`?U��?T\m?�ٺ=Y�?��<>��>�â=ZI�>�D�>��?��M?׽q?TzJ?���>�͙<װ�ଧ��B��PҼQŻr�D<��m=<�?�³u�G�����<��2;Gż4��� �G�`�17��;r�;���>�2�>���K�E>����������,>��<B���7���k"�LƔ=�$�>�y�>"|�>Ga��>=x׹>�>���`I'?cH�>;?��l=�k�{ƹ��.X����>�H?#Z�<�;X��X���ck�n�Z=�h?�r]?�V�!��I�b?��]?3h��=���þ��b����a�O?;�
?3�G���>��~?`�q?L��>
�e�':n�(�� Db��j�"Ѷ=\r�>HX�H�d��?�>d�7?�N�>�b>7%�=Yu۾�w��q��a?��?�?���?+*>��n�W4��ݾSV���:O?�u�>⠾��W?͛�=b�⾾^���
���+뾐����_Ӿǯ"������#������S�	
�=v?�~?�bP?�|?�>WX��~H�0⏿��Z��NǾ�о8^9���H��"P�/�v�OC%��Ⱦv���88�<�v�n6�#ճ?��?4��
�>�V��]�����A^S>�>�����iV=A�L����=Δ�=w�K�\�5��y�?�&�>��>3�B?m_�v�<��Z.��A;����AY->"�>Å�>���>F�';�"�$0齑J���	P��Lѽ�M>�7V?d'@?�?j?��˾���΍��*�]�u���q�	��=qK>=U��>��ľ�O��R�@:O�ryy���(�ℾ1��Is�=g�?%��>{��>�,?�n%?�Eݾ�����@��	~�6��=��>	=?:#?e7:>�Cp����H�>ֻl?���>j��>WP��r5!��{��pʽS��>,��>���>2o>g�-�/;\��X�������<9����=%yh?����[�_��9�>{�Q?덟:+�F<h�>(�v�O� �� �oi)�9
>��?6��=��;>I�ž���Ym{�=_��$Z?=_?�0W�7��T>�>��?'��>�/�>�Å?�q�>�E�E',:��?:Ok?(�K?�C?��>��@=L�������(��-�=z�f>/�<>�aF=�LF=��/�P�V��V���9�=��=[1{�wy�Z*T��Q�NdB���?<��$>��ٿ�KR��c־ž边r���$�VD���h������&�V���+W����V�QG�vm��Bl�cW�,�7�U��'�?��?�Ӽ���z������X��&��^�>�}}�YrF�G����r���5�}�վ��ݾ���SH��AZ���t��{K?kP���Կ����eN��+?�(!?D�?\9����%����=;��=d7=>�4��<��q_ѿ'�@��@?R(�>�3��ɹ=�}�>�:��<S��>�w��5(��Ӳ��>;�>��G?a�?�N�@�ȿ{�ɿ�L>|��?��@�B?�E'��쾉�F=7��>��?@4>��5�I��jC��^?�>�n�?Ox�?��Q=%�W�� 
���g?���<��D�1����=���=��4=���GK>�>G��H�G��B�5>�@�>��)�!V��ET�iA�<��X>�E̽@Ӌ�5Մ?+{\��f���/��T��U>��T?�*�>V:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=~6Ἳ���y���&V�{��=[��>e�>Â,������O��I��X��=>��+,��b��~����'&��(���/^��ڽ]���l+���������t�=��	>�eD>�B�>̙Q>-�.>eH_?j�T?+1�>4��>1m��ç�M�����U=c���_�Ͻ0򻽟&H�w����ԾA��I(�9"�+�������,�x�6��lV��Rp�q�$��P��/�/�*?6:����D���<��{������~���H?�0þ�U�sL��?<��>F��Zdu��۾M�A>p�<�a0?m�}��R�%
����:>���,m�S6>+��>o˾��T�ֈ{�t�<?k�?����[1�`��<�׽S��f7�>"X?k=���>�>?��'=�H7���~>�<!>��?��?�t>����n"����?��}?@��gX��K! ? �+�%���u>�ѿ0>�1&����Q�D>QZ�>��*�z�o�Ƥ����<��^?�a�>W��w)�q������?��W?�m,?�0�>:�X?�\\?<�C>o+��%�e���۾��>W�O?@<V?��>���q��ӏ�jI&?cGf?��`>Ӭ�� ���,��|��֜�>q,o?�v/?�r�膿XC��S���!�:?:pv?k][�`����y�4�����>��?���>�nG���>�pC?�L�=���m��Z�A�޻�?�@�N�?�%k=����>#"?��>Fi:��־֎��c��i��=/-�>V���Goy�|�%�6M�~7?���?���>�^�]V�<.�=�À�;u�?ө�?7u̾8]#>��?�}�[���;j���7>q �Y���M��^�I�����
�63оf�6�h>��@�ᮽ���>�<f��<�yrοI�v�~�Ծ�C��Q`!?qל>|Hs=K0��O�Z�b傿?s>��a,��NK����>�V�=fL�������y��7����� �>��T�{�n>.�J�5�������eA��Ƅ>b��>��>��Ƚ�-ξf��?�G���3Ͽ]&�����z\?�]�?BK�?$1?���<�^s��a��i��y�A?��s?[?�1��@m�=�{�1x?�1�`z���Y]��Kf�bL�>A|h?C?��k���=�s�>�D�>�]�=���O+ɿ�ֳ�N^�pt�?1M�?�}��}:?xw�?��(?�&�A����x�Z}2���N��#l?_�L>�)�[C6�\�f�,���b>?��]?�P��A���c?��u������B�^�"��>a��r��qw��A3"�_�R��ɝ��X��'ԧ?�l�?� �?��i�,�>a�>*A�>�!��J�ؾ�O=�c�>	7�>�\>��=��>n�����/�&>���?#��?��?s'���U���+>@ˌ?�H�>���?�D>[�?��H>ǎо���"�2>�>�u�6��>��E?�<�>���=��>�u�"�~&B��K����$:�+�>�Y?m�M?:vw>��#\E;*�P����ؽ$սEO%��ma�:s����K>
8=>V�><�v��jܾ�?�t���ؿDk��	�'��64?�Ń>#?�����t��O��:_?�{�>'0��+��:(���9�g��?AG�?��?/�׾��˼D>��>9G�>m�Խ��?�����7>%�B?�(�&D����o�H��>���?�@�Ү?��h��	?���P��Ta~����7����=��7?�0���z>���>��=�nv�ݻ��c�s����>�B�?�{�?���>�l?��o�S�B��1=6M�>Ɯk?�s?�Wo���~�B>��?&������L��f?	�
@xu@R�^?)�?ӿ`o���ذ�LZ����=�!8=�y;>��UXX=��5=���x��:;�=F
�>��>�s>`hK>+�7>��4>�p��Z� ���������zyI���#���1y�����0������-����Ѿh�ҽ����r�s�x�6������S��==a?"Q?���?](8?�/���g>�6׾h��<%R=~9�b�=�6?D)F?;3?d��=uy����f�(T��ꨂ�9��!��>h�D>�^>�	?�jo>tk=��=+�>�Ѩ>�e�<��j>:{�G��=�-9>���>���>���>��j>�G[����������T�]�̽��[��?$ҾFzY��h��rD����ɾ��/�ȟ?��_>)
��L�ʿ�̽�]VR?�����*��5��3jV>>F?&3S?��!>�K��<p�=��=V�]������L>��=�bJ���*���+>d	?��f>)u>��3�d8���P��_���~|>�,6?9ֶ��E9��u�.�H�kݾKM>���>ĲC��i�����A�r_i��O{=�x:?b�?WK���˰�S�u��W���6R>B\>*�=�m�=�JM>�-c��ƽH���.='��=��^>�?\^2>��=e&�>�@�T����>�u:>jI1>(j>?�?�������?`��#�@My>Br�>"�>�=>�H���=9��>	m>����PX���f��V�=�HP>�Zu�3�a�^�f�ݣ\=Ic�� �=-�=mv���B���=��~?@����ꈿD8�2����iD?�4?�ّ=��B<��"����|&�����?3�@e�?��	��V��?oB�?@(����=8��>«>�cξ��L���?�ƽ�碾ݑ	���"�!N�?��?,�/�I׋��!l�0�>�k%?_`Ӿ�d�>=o�.Z�������u��#=m��>�9H?>T��t�O�&
>��u
??0_�0����ȿm|v�:��>%�?b��?Z�m��>�� @�Y��>G��?�fY?�si>d۾JfZ����>!�@?\R?��>	8�K�'�w�?`ݶ?ڭ�?�:>���?,q`?ׯ�>�s����+�������N�Mֽ([u>`��>��2��d�Y��e����7i��q>�e�:>Em/<،�>[��������b�>��;߾,3(����>��M=�kk��M�>���>��> �>��.���'��Ij��e��D�K?Z��?F��%0n����<^��=��^�8'?WH4?g�[���ϾҨ>��\?���?�[?�c�>���|=���翿>}���Ŗ<��K>�4�>�K�>�8���LK>D�Ծ�/D�t�>˗>�����AھC+��F��zB�>�e!?���>>Ю=� ?��#?d�j>�)�>�`E�9����E�z��>��>�G?��~?��?�ӹ�|[3����硿�[��4N>I�x?�T?�͕>ȍ�����4XE��jI�2�����?�tg?S�>?�2�?ފ??�A?l*f>���ؾ�����>��!?�]��A�gQ&�<��o�?�T?��>z-��vֽ��ؼ���~���?�\?;&?͝�6a�*�¾��<�U&���A�n<�F��>>~쉽�=?�>��=@m�Q�6�E%h<vH�=
r�>I�=QQ7������f*?D;��}V��Ī<LGv��?���>�^j>V��d?7g�馅��E��U��g��k��?���?��?Q�={�u��@]?F�?��?%�?Bm�����HʾJ㒽�I��G�bcr=i�A>�7L�厜�����3��#)��er���M5��?�HK>2�>
8�>VT>d�>Ԁ�n��sOھ�3ξ[�V�!>�=�<��0�Cy(�b�ݾ�1���=Z<�������>\��>S}?���>�ޜ>%�>Yo!����=��><��>�_�>)TO> P�=�϶=a����^-��FR?r���@�'��辂���t;B?nd?�/�>3i�牅�T���{?ځ�?Fs�?Av>uh��)+�l?_8�>c���g
?��:=0��(�<B����s���:G�?��>�*׽O:��M�b[f��g
?�,?�����̾-P׽Xۖ��D�=�?X+?ڟ,���I���g�� ]��T���*�ܪ%�4Ǩ�� ���t�r����� ����\*���.=Fs!?��?ݰ�zI꾎w��էv�
YP�Tl[>�><��>ɲ>B�|>����^6�[�P���)�����$�>��u?�I�>.u=?ų?�h?��9?J>���>�a��)+?��,�m�=�x�>dp(?)�U?S�r?��.?n�?���>��(>d[�x�9��n1?�:�>�.?+��>�?P_G�.�l<�}=��H�ҍ���%�6�+>�=׼�+S��+T��)�z>IM?Ae�y�8�����Hk>�|7?���>��>`��[-��� �<���>0�
?�-�>� ��r�%k��H�>���?9+�Q
=
�)>���=�>��>��L{�=7���5�=�n�<��#<�N�=8�=]Yr�	���ٖ�:Iʇ;̉�<�u�>^�?���>B�>�@���� �����f�=_Y>�!S>b>�Bپ<}���$���g�kby>-x�?qz�?�f=��=���=�~��-V��������{��<��?�J#?�WT?���?&�=?�j#?ڷ>,��M�� ^�������?v!,?���>�����ʾ��͉3�ڝ?g[?�<a�!���;)�ڐ¾��Խͱ>�[/�m/~����6D�U녻�����3��?翝?�A�U�6��x�׿���[��s�C?�!�>$Y�>��>R�)�}�g�u%��1;>���>kR?��>*�O?&{?J�[?)�T>�8�e
��x����2�� >��??�p�?�ߎ?��x?���>>^�*�2�"x��,����`݂�_9Y=��Z>���>�l�>[�>*A�=��Žް��J<>��ã=��b>�~�>൥>&��>�#w>E�<�;P?o�>�c������ѯ�"�������T�h?)��?
Y?X\'>%���C���#�Ǩ�>j��?q;�?{�?J�R���>�N�<V�T~���ء>�{�>�,]>�Ͻ���>�\d>�_c>�d�>��ף�5^�%�8���+?+??�	
>(�ܿycx��"�����8ƽ>�����B=Ե���D0>�_�+X�3�۾�h�%)s�rH���	J��=�<Ŀz��?��-=���^>_�<��（ϭ<�N�=�pW�u�=AK=sLX=�c"=��o;p^��g�U�e;i$>������ɾ�m?BJR?���>a�W?o�>ȥy>Q����>{��<	�>h"�>��l�:ہ��Y�q.b�x�Q���.���vS�m����}�<ʱ)�;�=E��=��$>ZL>a�L�ˍ^��2��ɷo��jC=+�$=��>?��=4��=̞6<N6O=�t?�a������x�i�6̽�bX?��>���=g���?��@>�i��������Pl?"��?k��?�(�> 侷��>�.��J�$���6��܏=j�>���=�|	�K��>��>P$�
3���ӝ����?
b@��%?:��n����`>c7>��>l�R��1�k$\��\b��Z�7�!?!);�$1̾c3�>pJ�=�v߾��ƾ�--=��5>��_=�y�;\����=�Y{���==��j=׉>�D>��=ޟ��o·=��G=]�=#OP>�=w�;66��+��;3=G��=6�b>b�%>|��>�'?�[8?��X?G�>�]\����b��Y4>}�|> �?�<�v�>��V>d�+?t�V?)#0?�{�>�T��4R�>�A>��K��텿��LVӾ����^z?&�?g��>��>�n>Pq%��BP����=A8?�Dm?X4�>G�>1$�1�ۿ���÷,��S����}���<|��r�����v#b�Y��R�=l��>bB�>^�>�Oq>��6>��K>O�>-_�=�L?=�c$=��7=�{�=;������=�M�:���9�b=	;�ְ;�Z��@���5e<��K�A��ǎռN��=���>�����>@�u=F��@�D>��*���P���0>�@�C�`�3	��o����5��
(����=�p>�B�=&���Hz?"z_>���=4��?qnf?34�=����8�����?'�?�$�<�">�޽��F��rw�;r�:oɾ��>��>���>
�l>,�� ?���w=l��_5���>5p���-�9��8q�W=����.i�Ϻ�D?�C�����=L~?��I?�?�w�>���Yؾ�[0>$@��M=��-4q��`�� �?Y
'?���>��I�D�cR̾R%��2޷>W;I���O�OÕ���0��^�η���>��k�о0%3��f��������B� Ir�A��>.�O?��?g7b�LV��QO����/6���o?�{g?�>.L?�C?����y��v���n�=T�n?v��?�=�?p >�[�=@���Ps�>��?,�?Ў?��q?�VG����>�צ<�h�=�`����=$>x��=.<�=S 
?��?6R
?�ϓ�9�<3߾I{�LEh��0 =c��=3,�>-�>Ⳅ>
��=��h=
)~=�jJ>f��>���>*h>�P�>�p�>�3��>־gy?KQ,�I�>��Q?}L�>�GK>[�$<���po��~��g:�ޢ�<�"��;��<��۽��)�ߖA=���>�^˿{ڠ?)N�>���.?�޺����L��<�
�=i�=�S/�>�'>r�>!�>�'�>'q>x��>���%GӾC~>����d!��,C�K�R�W�Ѿ^~z>휜�V
&�����y��BI��m���g�nj�6.���;=�[Ž<DH�?�����k���)�����Y�?z[�>�6?Vڌ������>
��>�ȍ>�J��`���ȍ��g�b�?���?c>�#�>%�W?-�?�Z1���2�mMZ�P�u���@�2�d�3�`��̍�i���&
�Fɾ�ض_?��x?�|A?�l�<8Xz>ђ�?��%��y���Ί>B"/�;���:=
ߦ>+��=a�l�Ӿ{�þ�
�OF>k|o?y�?�l?h>V�R����j>wd?��)?>Da?+��>�3?�/���q?)m�>O�>�� ?���>�	1?{1?�Z>�ɐ=Q���6�R>+�ܽ�R�`v��w�=�d=��%�4�����
滷��=@��<`�Ӽ㛃<頼,���f�p���<U�>g.�>reN?�]�>�H/>��?ѵ򽭫8���� C?�^o>�I��ɝb�����.D��n��=v�M?�?X*`?�r�>G8�G-r��9�=y�>Z�<V>V}�>R+�;���;5`�29D>�~�=p=fq�<3������jK���@E=HM>kb�>YU�>:�y�^}&>R��/eu�Dg>�U�8ֱ�/�M���I��0�S�n��,�>ӰK?��?��=\��Rky��>e�1/'?06<?> J?n}?��=z`޾j�9���H�d�]/�>���<�
�� ������S:�IM��9_n>�柾�࠾QQb>/�� q޾��n�?J� ���M=܀��tV=����վ�2�L��=�)
>������ ����`Ԫ�2J?�aj=Cp��soU��k����>���>@�>��:��w��@������+�=��>P;>������}G��6��<�>�QE?�U_?Ek�?�!���s�u�B�����_d���*ȼ7�?nw�>dg?B>��=H�������d��G�/�>۞�>����G��6���/���$����>�9?��>C�?l�R?m�
?�`?h*?kE?/&�>���5����A&?���?F�=u�Խ��T�� 9�aF���>˃)?��B�鷗>}�?	�?�&?ǆQ?`�?0�>�� ��C@�Z��>�[�>��W�}b����_>��J?��>�>Y??Ճ?'�=>��5��ꢾ/٩�!P�==>n�2?L6#?q�?���>u��>T����=���>�c?�0�?�o?u��=$�?|:2>#��>���=���>^��>?\XO?4�s?��J?ܑ�>���<�7��e8��XDs��O�-˂;�pH<��y=����2t�L����<���;&h���G��g���D�������;�@�>��s>�*���<1>�ľq��ePA>a��RJ������E<�;�=bt�>6�?Eҕ>?�#�ٟ�=�>r��>B!�wk(?�?�?Gz;��b�)b۾�WL��ٰ>��A?y��=,Ll�/p��_�u�~g=��m?�L^?�W������l]?7�^?�.ݾw�;�7�̾�Mr>Dxؾ�?$��>��˾'Ǻ>���?�]�?4��>��˾L���g��3[�>�=9��=�ݫ�S�+�Z0>�]�>1�?�=+�Ž{6\��g�������>�Ԋ?���?�Ճ?�� >W�X�s��}~��}K���^?v��>�?�� #?������ϾYP��)����V������B���w��>�$��݃��׽��=H�?�s?U\q?d�_?� �8d�62^�A
��MkV��(�&���E��'E���C��n�4b��/�������G=g,~��A�E��?�m'?0z.�Bl�>Ɨ��g��;�AB>]K��*��6ǝ=�}���XM=%Kf=pg���-��\���2 ?�;�>��>Q<?��[���=���1���7����A4>�S�>Q�>>��>��X:�+��G��,ɾ�փ��ӽ�.v>~wc?�K?��n?�g�)1� �����!�0��a����B>�j>$��>5�W����6&�{T>���r�����y���	���~=)�2?�-�>��>pL�?V? p	�-l��&Vx�ʁ1��d�<$5�>�i?0K�>��>�нl� ����>4�l?ۡ�>���>���jE ��|���� 	�>��>d��>��q>~k-�	\�����e8��P[7��F�=��h?�����n`��G�>�R?���:��3<��>Y���!��2��:3+�<�	>��?%$�=F=>��ƾ��4�z�4��P)?wK?�蒾��*��4~>�$"?��>�-�>Q1�?�*�>tqþ@CE���?G�^?OBJ?lTA?6J�>E�=���=Ƚ��&���,=��>��Z>um=Ȁ�=Z��s\��w���D=�s�=O�μrO�� �<ȃ����J<��<��3>~-ֿ�/E��s��������!�.u��v�������"��h�����h�VHp��N�l���w�kt������J�E�?�i�?����i��M�����Y��Ծ�H ?����z�]�ƾ[���ط���FӾ/���!\��NT��jy�0&V��'?�ȑ�һǿ�����ܾ ?N> ?l�y?z��"�ڊ8�@� >��<x��մ�$���p�οn�����^?K��>;'� �����>A��>u�X>W�q>�����)�<��?��-?l��>u�r�8�ɿȁ��j��<g��?��@�|A?;�(�Z��(V=���>]�	?��?>Q1��H�����T�>Q<�?���?�xM=��W���	��e?N{<��F���ݻ��=q<�=0M=�����J>SV�>����TA�"@ܽ�4>�م>=�"������^���<�]>��սg?���3�?U�_�]P^��w(��{�T>x�{?��>�h�<��3?��l��Wп��/�ź�??H�?�-�?Hw?Ɵʾ�>\)��ulS?�-3?�X�>8?�2���t��=���<�p�$�øK��q=��r>Zc�<�ݽ������L�wծ=�����ſ%#�9��_f�<��'��[l���<����;�j��lj�F@��2n=dc�=v�K>���>$;Z>,?Z>�Y?�l?��>
>�<��z���ʾ�>;h���FN��~����Cӣ�r��`ݾ�	����~�e�Ⱦ��<�W�&=�/H�r�H���s]��&?��-?�6�=W7���;A���H=J�;>q��ۘۼ��潎4۾|B5��c�G�?�5?4����Z�.���l�����e?��.�K�>���o�$>��7���=�s�> =+8��h�6��C�'0?��?؀���V���">�:���<g�+?��?�?<�>P�$?��/�{齔T>j2>�>���>"E>�谾�%ٽ��?V|V?�4��R���!�>����g w���>=�>�0�����=^>���<L���&RH��F���M�<��L?M �>��)����?}��#�>�y�oT�?M�A?�I�=2v?9lh?���=��	�Q�j���$�4���gD?KT�?#�V>+�<�����h���b?+��?$>�=,_�<�-0�,�&�1����?�d�?:�?�ι�|�y�2d��x�4�n�G?W5w?}b�� �����V�'�I(�>m��>��>&/>�-��>�R>?��U���྿��0��͞?�@j��?�d�����=�R ?���>z-U�m����q�!4��@=&�?ɻ��N�������C?�x�?��>UI���
����=�ٕ��Z�?��?~���lDg<R���l��n��U�<�Ϋ=���E"������7���ƾ��
�����࿼˥�>EZ@�U�w*�>�C8�]6�TϿ)���[о�Sq���?M��>V�Ƚ����@�j��Pu�a�G�3�H�ť��qL�>��>����G���3�{�s;�I����>���	�>��S�r.��ޤ��05<���>���>���>/��X꽾�Ù?�T���>ο�����V�X?[d�?�p�?Au?��9<i�v���{��f�y'G?��s?�Z?�G%��5]�8�7��j?�]��U`���4�=HE��U>"3?3E�>��-�l�|=�>2��>�k>�#/�j�Ŀ�ٶ�������?"��?�n�J��>7��?s+?�i��7���X����*��/��<A?�2>t����!��.=�bВ���
?�}0?^|��/���f?#��iH���$�5��<4��>E��������!�O�n=67\�̦����c�H_�?j�?|��?���*?�!�>�np������ �<��Z>��>(8>�r���'�>\~�כi��hi=H��?��@�
?Q8��X���-�=��r?�0�>ux?�R�>m	?�9��U����->?fK>�!#>����4
?�R?���> <5>Q���u�J���x�En&�
�d�v>��Q?0_?��j=�h��.ǻ:�8A�o"���>��=���M�3+,�a>-	>%��>�;f���n�� ?tg&�1^ٿ,͙�O���`?�>?�?���MB��}_����g?Șv>��O{��
E������?<�?�?��������I>L�>n<�>;W��'"�ڥ���$g>��F?�3�47��.�r�彋>��?��@�?��e�d�?W��Z��}p~��"��(�*�n5l>81??��]<a>#r�>�A.>�1p�����x�倭>�b�?�G�?�F�>�e?j*��9���>�E�>jփ?�E�>�B����A�>�:?��9�N���ݸ��i�?��@n@�R?�뫿�pֿ�����5��/���޶=���=�h2>�bڽ4Z�=��7=�Q7�_������=��>�d>
q>O>�F;>��)>Q����!��l������8�C�A��w� �Z����=@v��~��=������d��D\ý����Q�8-&��s`�I�=$(V?�S?��p?b��>`����#>0���>
=��&���=D��>�
2?�K?De)?�ۊ=e����pe�k���'����8���1�>*vG>�(�>�,�>W�>���sJ>H�>>s
>��>�)=��$��=�jN>O�>���>��>�C<>��>Eϴ��1��h�h��
w�x̽1�?����Q�J��1���9��զ���h�=Eb.?|>���?пd����2H?)���)���+���>x�0?�cW?+�>$����T�-:>-����j�3`>�+ ��l���)��%Q>xl?a�f>2*u>ے3�9^8���P�!f��r|>�76?�޶�/09���u�آH��^ݾcRM>���>�D��q�L���d�9�i��F{=�x:?b�?by���밾b�u��P��5TR>�D\>'u=�*�=�CM>�<c�Ұƽk�G�2�.=���=l�^>�'?7*->-��=�^�>uY��bKR�9��>=B>�6->�r>?��$?����Z��!$���60�Qv>�2�>9�>� >ȎL��,�=wi�>��f>s� ��Ǆ�}���C�bX>�ވ��`��j�	�q=�M��ѵ�=���=E ��*<��&=w��?��������|޾u=��O?��?�颽仚P⾇U��5Oݾ�e�?t�@�J�?�$��PI���?4�p?J��(�>��?���>	A �@:���F?�m���
��<�V�ľWђ?�L�?aO>S,��ڢT�7=h;?�Vi�j@�>�A��K��^���I_P���R�3��>sS?�����ҽO�?��"?���>]��i����rȿ�x����>��?> �? �v��ݡ��-�O>?�&�?�og?$�?>P۾Z�Z��ǈ>�n<?Y�H?�?�>c!��"�4 #?:x�?���?I>���?��s?*l�>b1x��Z/��6�������n=�j[;�d�>�W>-���ggF��ד�~h��I�j����p�a>`�$=�>E�i4��;�=D��H����f�j��>l,q>N�I>(W�>^� ?�a�>|��>,z=�n��0ှ�����L?�D�?���O�l��L�<�z�='yX���?�T2?vTd�@ ˾�Ȯ>HXZ?Y�?;�X?���>8��gΚ�`\��u����	=<��T>��>.V�>Vy���L>��Ծ�_>��<�>m-�>Ě�5.��G{��Z�;B�>�� ?G��>e;�=�?�/?i�=>�I�>�DA�H���k�F��-�>i�?�E ?\K~?Ѣ?��̾�*:��
����c�M��c�>X.�?lW"?�,�>��蒦��n�t��=.	��΋?�\i?�߽� ?+��?�YR?�=?TH<>��,�2���(�}��>p�!?e��A�L&�����?�N?1��>Y8����սּ����w����?x$\?%:&?@���+a��þ��<7�#�P�8 <�dE�.�>H�>8���)��=}+>}԰=�Xm�'f6���g<���=���>#�=�37��Ύ��$&?)ʁ=~DQ��F�=�cr�NR>�n%�=�>�,z�|Y=?=᩽>;h�'������ #���M�?���?��?P	���g�;g.?��o?u�O?vh�>&(ԾvTɾ���x=;�[������B��>ᯒ>S�=�-þ;c��~E����I&�;�b��T�>��n>g1?�	?��s=�+�>;�ľ$>�fW��v��[V�Ec	��,�1y��,
��^y�������mP˾|�����><��(��>���>,o>~FB>	f�>$����>�qR>f>��>��>��>�b >�7�Q)��ZW?T���R-��x߾�7���YT?>'�?���>�����<Z�2Z0��.�>���?	��?;��>�#R���)�C��>(/?nѕ�;�?E�>�R��*f�S����=�0;=J��ԫ�>xw��vN�r�X�5�<�kA?ZH?^2�<���",\�!���M�n=�M�?��(?�)���Q���o�͸W�S����6h�Pj��M�$���p��쏿�^��%����(��r*=��*?k�?Ҍ��!���&k��?�wdf>a�>a$�>7�>.uI>��	�q�1�b^�M'�G���`R�>t[{?��>�I?�<?GyP?KiL?���>"e�>r7���d�>CR�;+
�>���>F�9?��-?+40?*s?�p+?�#c>���l����ؾ�	?�?-H?�?خ?�ⅾ�Uý�2���Xg��y��x���!�=>1�<��׽oPu��T=ZT>�Y?]��K�8�d���	�j>׋7?�m�>O��>
��%9��mh�<6�>��
?=�>! �M�r�j��K�>���?k���#=L�)>���= ��p�Ժ^��=������=�3���<�mz<I��=r�=Br�V̌��:���;u�<���>o6.?��M>9 �>G�P�����L����=Ll�>{ٍ=�s`>X9��(���_��PTi�\�Q>M�?�g�?3]�,46=$v>��Ҿ�P���K����Z���=X�>��5?5(?V�?�L?�?z��=F��F��u����t�\�:?h!,?��>4���ʾ,򨿘�3���?�[?;a���;)�k�¾�Խ�>	Z/��-~�V���D�\��� ��p|��P��?5��?.1A�2�6��w�󿘿�[����C?k"�>-V�>��>��)�6�g�|$��6;>Ј�>�R?v#�>n�O?9<{?Φ[?;hT>~�8�N1���ә�_V3�~�!>�@?ϱ�?��?y?�t�>b�>g�)��ྙT�����C������W=�	Z>6��>�(�>��>r��=HȽ$Y����>��`�=}�b>���>���>}�>��w>�H�<�99?���>,]���=��i�E�S��Ì�Yo�?�p�?�Z?��+�M��s�A!�2��>���?�2�?y�I?�>�u^�=v��=������@�>~j�>��J>�>��C=�%�>�V ?��>`4�~��w�X�+���6?�g?b����ɿ�Hr�3�L��`��ye
�(:��s���0���/G�92�=Ūv�4�������?�7��b��H,��fାu#y�RZ��	?��=�^�=���=��<ߋ]���2=C�=m�8��=U���l\=�cl�������{6��㹻��=V(л������?W��?��b?"
?��5<?�>	u���>Ŧc��iK?���>p>9>$t��m�վ���d2����C�������:c>a[��>��=A��=�J�<5�7=�
3>)j�=(��Ǣ;=|��=���<Nx�=K��=�RQ>+��=7�y?a���#����]G�w��={D?�<c>8v=#��~S?��^>00y��Ƶ������u?�w�?O_�?_�?꽏����>3gؾl�'�� �=Y��*�>�۽α��2a�>׆�>59-�=u���<����?�S@�"9?i�eտ�$�=j�7>�M>�R� g1��<\��b���Z��t!?�X;�6̾��>���=;߾��ƾa�.=x6>�b=�]��M\�}�=�|�m�;=��j=��>��C>���=�A��ҷ=�H=[�=��O>6Q��,[6�_�*�i5=���=8~b>��%>��>��?W1?(�K?�'�>RQ����׾�oϾ�w�>���=kPt>�v��Y��=j5�>]nP?�=\?�4D?��>[7�<��>E-�>��6�U�o��n�f���hb�	�?�3�?��>x�<��P+���=���ʽ��?>�.?	=�>f��>B���ƿr������r��5�ݽ�8�����߼��D�},<�|l�˱�=x�>�C�>+,o>�Ut=ю�<Q
>>�>nx=�1���ԁr�2��-���
�<�U ��3\=?8���4�=}��U����#�� ��D̼�$�=��<��=@`�>��=d{�>j�=��Ͼ�A�=ኜ�6N��u�=jk����>�E^���y��|,�_[@���n>�nT>�w�m͑�(?�f>��n>�N�?��d?B��=�V��Ǯ�BI����������u=���=@r#���/���M�D�=��Mվt��>��>���>�m>�+��5?���v=�(�͊5��0�>C���1���$�Z2q�a+���柿z�h�OѺ��D?�G���=L�}?o�I?!�?R{�>������ؾz�0>��=����.q�����}�?S
'?���>d��p�D�[H̾���޷>ZAI���O���2�0����Zͷ��>������о[$3��g�������B�FMr�>��>2�O?��?�:b��W��*UO����"(���q?�|g?�>�J?�@?Z%���y�r���u�=��n?ų�?\=�?�> ��=1��-;�>+	?Կ�?���?Ăs?��?��s�>�~�;�� >ɘ�G�=��>���=�7�=�r?/�
?(�
?�a����	��������^�v��<š=��>�n�>��r>���="�g=�m�=S/\>�ܞ>��>��d>G�>�N�>��Z}����?i$�=�?�>)��>��>w����e����}6.����!��	`��a!>i�Q>�+=,-λ6�߽w��>ܖ˿(��?�b=e���4?�
���-.��D=>?a�=p���|I�>�=��z>E�>��?�s�=�2�>�>M����=)#��0@����ǟZ�rǾ�պ>�b����;�چ����U�I�m�3���S��zam�����A���L=FS�?�?n���8$��C =�a�>$��>-�9?�G����B�hH�=�;?ր�>M�x�fӊ�wl˾^݋?�e�?rKw>�zo>��V?���>�g&���t���R���t�*�4��9L��j�F����ڀ��m����>3@~?��f?Op2?�� ��/�>��?�6����l%>�;!�dsI�9�>��?LC����8�).��}���S���?>zGs?ԍx?Í?	�a�1/��ߢh>p�P?A6?�o?Uw&?��A?�6�(�?��Q>��?��?ac3?��(?�?�w�=7&�=��a���|;�ԕ������7a������̼��j=*�=X��;t=�Z=L�����ϼ_z����;i"o���=���<��=���=]��>�Z?r�>ꧪ>7y!?��9��l=�����e�4?L�b���[��r��#;����I=d�Z?���?��^?{#>�s����]-�=E��>�RI>#_J>��>��K�n�'�����d!>�1P>�S=���kyT�I��H߈�;��=,�">��>v�>�"��=>W6������o�>#B�_���}�����?J�"�j��>�[Q?���>���=K�پ�X�<a���om?�_?�U?0��?B*j��;�O9�S�A����?Q�8>����̾�����}u!�x�=ӯ�>݈��4ϟ�̸`>I�
���ܾQ	n�d�I��n�<�==�����U=����־�T~��$�=��>�G���� �-���������I?.4h=X
��t�U�S���^Z>���>���>*b9�SL���I@�`����ؓ=$��>��;>�=|���F�`��A�>�=E?�a_?hh�?x'���s���B�:����w���mȼſ?�d�>d? hB>=��=�b������d��G���>���>�����G�et���%����$����>�/?#d>	�?ǯR?��
?ݐ`?�*?�M?N�>r���k:&?2�?���=,ڽ|OX��19���D�O@�>|)?�zC����>/E?�?Y%'?�Q?i�?ʴ>� ���?�"��>A�>�W��Z��~�^>��J?��>HY?W��?)�>>y�4��Z��B�KB�=��>�s2?�"?��?�ڹ>o��>?�����=מ�>�c?�0�?�o?��=7�?�:2>K��>��=���>U��>�?GXO?7�s?��J?��>��<�7���8��Ds�	�O�Vǂ;GuH<��y=ݘ��2t��J���<r�;�g��EI��[���D�j������;��>��t>�`��$3>�1ľ*���a@>�)���{��������;�T�=�>�?Bߕ>�t#��w�=�=�>���>]#�V(?�	?�?u{�;�Mb�K�ھ9K���>�cB?�S�=lTl��~��%Gv�x�b=�?m?^?XrX����e?�g`?U���b8�.�'�w�)=5Y��@L?�G
? ��J�>���?�n?'��>P���Tlt�����+tl�L!ͽ��2=�̧>���vA�|Y>s׺>�Μ>��|>��ܽ��e��f�Ͽ�OW>�<q?6F�?5�?FP>퀿��w����H���^?'c�>�)��a�"?P���̏Ͼ�<���A���ᾢ���c�����Ꙧ�5�$������ֽ]��=�?as??\q?!u_?�� ��d�^�X��XV��j+���E�iE�9�C���n�fY��F���G���[H=�:`��x>�d�?i&?']���>,���l.	�fe׾�*5>�|���F#�ԃ�=.ٺ{��=�W�=�u�Jz�A#����?0��>�U�>5?$�k��4��0�U ��F����=�6�>�_�>���> X�<y���=�(ʾ��f�=O��z9v>�c?sK?8�n?�����0��j��vq!�41� M��r�B>lz>#�>�@W��n��D&��N>��r�O��5���<�	��]=+�2?���>o?�>i7�?�?lb	�u����Qx��}1�{y�<��>��h?!3�>�ӆ>��ν�� ���>L�n?K��>�U�>�
��é%���|�����>�>�0�>ƿi>%8��O]�Pm�����T�.�[>W�b?�	���HR�11�>�aT?��;~�<��>>���������>�B�/�>��?���=T�@>7�˾�@	�[\y�-?���O)?{K?M蒾[�*��3~>M$"?��>�-�>:1�?�*�>�qþA9F�w�?�^?xBJ?�TA?�I�>q�=��W<Ƚ��&���,=���>l�Z> m='��=���Mq\��w���D=vt�=ܥμP����<�}��M�J<���<n�3>��ٿ�M�d䵾�4�*d辸V�y�f�r�r��`���)��v䎾`u�hQ����̽��U��9m��X���`����?���?��i�㭴�24����M��J��>�ㆾ���糾�
��S����ھ����B"��R�(�e�qaJ��'?ƺ����ǿ���(;ܾ�  ?�A ?�y?���"���8�X� >�D�<�+����뾰����ο���6�^?H��>���/�����>h��>�X>�Iq>u���螾�,�<��?p�-?Ϡ�>��r�	�ɿA���yĤ<���?�@^}A?��(����OV=h��>��	?��?>�L1�fH�����HS�>�<�?���?B�M=��W��	�C|e?�V<}�F�k�ݻf�=�>�=3Y=�����J>�U�>Ȃ��UA�0;ܽ��4>}ׅ>��"�4���|^�M��<҄]>��ս7K���τ?#S\��f���/�T��7\>g�T?��>��=�},?�I���Ͽ��[�Bb?���?qL�?4 (?�"��:�>Aeܾ�(N?�@6?�B�>��&�>�t��S�=,�༤�������V��c�=���>C>�-�rz���M��M��D7�=�L��+Ŀ��˲�,��<�,¼�	��ǽ�ڣ�U8��d�����[�?Fݽ���=��=��@>-Wv>tT>��O>7Z?�hg?p��>˜�=�	���똾z����K<�d{����a���!�*��t����ﾎw����������K�ƾ=���=�5R����� ���b��F�]�.?ru$>��ʾ�M���-<jpʾ:���-����ڥ��/̾M�1��!n��̟?��A?c���B�V� �*c�nz��z�W?�I����鬾V��=�ޱ���=7%�>֏�=���s 3��}S��b0?C�?͝��	א�<�(>�����	=�+?�f?@|A<Q��>9+%?ٞ+�E��%4Z>L2>`��>���>��>�Y��l�ٽה?\�T?�V��[����>�ľ��a{��\Y=dn>ͤ5���㼒�[>���<�ތ��K����H�<׏W?�n�>Ȅ/��J$��ʊ���f>$ҽ�ё?��?�zN���|?Z�c?� �>�3���c�l�/�v�����?'��?�v>J쑾�`<�
ܹ��?4S�?���>SXW��վ:.�|�ݾ,_Q?���?�3?2���.s�)��fn�T�F?�/v?x�_������C���I�Q�>���>Or�>2T:�n\�>F�@?_W �Ig��P���R83��6�?6�@7f�?�#;���p�8=��>���>;�6�q����l�7�����M=?�>c[���Vz�1' ��	'�h�=?���?� ?�����	����=�ٕ��Z�?��?}����Dg<R���l��n��i�<�Ϋ=���E"������7���ƾ��
�����࿼ͥ�>EZ@�U�v*�>�C8�]6�TϿ)���[оSq���?M��>T�Ƚ����A�j��Pu�b�G�3�H�ť���j�>�~>6-�����1<��)A�O�<���>_y��_�d>������˾���ܗ=ֱ>z?��o>U:��f���>��?�`���jʿH����!R?f[�?h��?�]C?0�<=m�釃��,��m�/?Ug?�KQ?iد���u��o�<x�j?fZ��6S`�ʍ4�EE�U/U>G!3?9D�>Տ-�	s|=�>0��>�{>!/���Ŀ�ٶ�����J��?���?Dm�"��>Y�?�q+?�d�7���^��j�*���'��?A? 2>c����!�,=��͒�O�
?�z0?Z���-��\?�Q���R4��*>l�?�M
�:}��}��0`j>Y�S��p��������?� @��?��T���O�ZZ�>#��>A,��ؾ����Tk9=�'>h�>�>��>�h$�3D{���/����?��?�d�>PЎ��<��H�c>��?��>�͂?��=2�&?�����@��Ay�:p-j>�ӂ�b����>;�P?Z	?k�>o
'����F�A�&ex��2F��hK�&�q>u�p??K[?j�1��p���4;�I6�
Z�Կ���>L�*��)>`���t�=�>ƅ�>��ǽ�**��?�p�}oؿ���(��4?2�>?���5 u����gK_?\�>�G��3�����w�.��?�C�?	?��׾3wӼ��>c�>��>��ӽk��aZ����7>:�B?���J����o�F]�>��?��@]Ԯ?�i��4?����Aq��=������#9�7N�>i#?J�����=-?��>/�w�T������A��>��?���?�� ?�z?�dx�"����#n>�8?q�?��>�<�������G�>`O?�/�ֲ��^	�ܓ�?�"@9@t�A?�����ؿ����\�����V->��=e�\=7c6� l�=Ao=wp�1������=!��>�^(>��L>K��=��=5J1>�)���"�PQ���邿 �.�Ml���"�^?��6���&��}�U���>Ⱦ���a��qㇽb�E��=�6u�����=��\?��Z?29z?���> d��[+>�D	�Ⱦ�����l�=�O�>��=?Վ??{�?�S<�����h��t�Yղ�B倾<��>�r'>	a�>aA�>Nd�>���9]>>>}�a>Qe>���<wd-;J[=gg0>��>u��>���>�F<>U�>�δ�t1��4�h��w�*̽�?����j�J�~1���6��Y����k�=�a.?Vx>&��?пs����1H?�����(�`�+�J�>O�0?�cW?��>a����T��9>���"�j��^>j' �zl�{�)��#Q>�i?Wj>��y>k83�˪6��dP�9���ez>/7?�Ʒ�`�7��t�g/F�VܾyXM>�=�>��p�v���1���l��5?k���o=z�:?cJ?&ɽ�Ų��Wo��8����O>�eW>�h!=�=�Q>��b���Ž�u?�~0F=���=��Y>�^?�30>P�m=	�>���>Q��>gM>>B�!>cyA?^<#?޶7��С�����}�*�r}r>(g�>�;~>�>W�M�6]�=���>�m^>�μ}Ћ�P��nA���W>n�x�<�\�c�z���t=�@����=r��=�4��<A�Y=��? W���ϋ��(���\�p4F?t�?�ۧ=�K�=���=췿�����?1@G8�?tվyP�9*�>kU�?崲�S��>>
? ��>�,��º��C?��ν)l��@1�c$z��?��?|��=�懿��]��S>Q�5?�����I�>�r"�Z����㋿"�w��~�h)�>�`F?P���b�g9:�R�
?u� ?k��-w��?dǿK�z�b�>qQ�?�'�?(@e�B䖿ܤE�OG�>�K�?��\?�ah>P�޾ȉk�G(�>L�I?5	G?1 �>��������?>s�?���?I>J��?��s?�t�>�Ex��`/�T4��l���b�=HN;�X�>�S>.����hF��Փ� g��>�j������a>{z$=��>�4�>'���E�=K䋽=���f���>�q>!�I>�R�>�� ?�]�>��>�,==h��W׀�U���5�L?=4�?�z�[bi�Kc�<�R�=�Oe�eo	??5+?�F���Ͼ��>�T?�|?F�T?˂>����Ĝ���������*<��R>�?�>B ڽ=]>��Ǿ`R_�*&>U��>�i��ܾ7��<�<��>eL ?L�>�:�<� ?�%?WAa>�I�>��D��r����F��4�>���>�j?��~?�?B���4�b���l���0rX���Z>��x?�+?UF�>%E��/8��g^4��s޼攽2i�?U�d?�ٽ?�L�?��A?�@?�]a>��g޾y���p�>�!?�����A�qC&�z��<z?�A?���>|x��8�ս�n׼����x����?�\?�+&?���#3a��þK��<��#�ltN��<��I�Ag>��>iS��,B�=z�>sİ=��m�a6���f<�ż=.��>��=�67��S���d&?�4>)\��!��<��\��9Z�Mk=�y>��#�?k ۼ�a��
������d<��&�x?���?���?����^f��VI?��w?5<?��>�귾$��]�%��*����ھ�� ��R>3�>��@=#1���d��ET��G�*����?a?��)>�`?��?4>~j�>d2��w;�r�P�����(o��;���%���	�@I{�UMJ��,��fƾ v����>�o����>���>:��>a�%>]��>��<�V�h>}�>e�{>���>�f>��>q^=t����B۽;{V?܇������v�����`?�qN?�`�>l\�<q������6??�?���? U>	w�6@A�&H�>�B?�yt���?�$Q������=q;Äl�R�������S�>w�/��5���U��H.�*�?�8?T,.����ط%������n=�L�?9�(?T�)���Q��o��W�AS�����4h�:a����$�p�p���\���$��)�(�@�*=�*?��?��[��9*��"k��?��df>R��>_&�>׾>�I>��	���1��^�R'��ǃ�L�>6a{?!�>ڧI?7<?��P?m�K?2\�>b1�>�[����>�t�;��>��>��9?[�-?��/?��?c1+?3rb>vN��������ؾX�?�[?2�?_�?v�?���V½�y���3h���y�������=S�<�qؽ�w�N�Y=e�T>z" ?��ڽ|�.����G�Z>;O?��>#��>�i�,&���BQ=�6 ?�� ?P��>�p�[�|���F��>�]�?�uȼT�o<�.>+��=���<��<t�=e�~v�=�J=γѽ�ƻn5�=�>>碞<ֻ���N#�dҽ���<���>'O5?U�>�"�>N�v������Z'>�ֽ>ܲY��^2>>Ⱦ}���8�����h��1>��?���?�A��rm1>�>d�ؾh۾>?�����+֕�j�.?�?�0?�<�?��H?ɐ%?�~=:������4ƃ�Rd�xD-?�%,?�ґ>���/ʾ=����V3��~?i�?�#a����h)��¾Z
Խ��>�//�2�}�����h>D��ƻ6���������?�ҝ?��F���6�辖���S:���QC?AK�>f�>���>\�)���g�����D<>�v�>7�Q?��>��O?.n{?�[?��R>�|8�j4ܙ�| F��!>q???�َ?��x?���>'>j�)���߾�M�������O���U=	�X>�N�>���>��>�4�=�u˽�{����>�w��=Ĩb>#n�>�ǥ>�v�>�Ex>���<� I?���>�폾�CB����|���1>B��?� �?�<?�(��^`�2�z�s���3��>.W�?��?R~!?����v�=���=AY��0YM�Ǯ�>�r>n=��=&�7>��>�[&?*c�>��%��9G�+�w�O�:�u�H?�/d?j�D�5�˿K[v��/1�]�~����<�U��P����v���iM�Bl�=���D����&�����C���ΰ�Y���3�f�Cp�>v��=��=bێ=�}�:��k�D!?=81�=.�!���=<�)��0,=�j����/��t¼>�;z�k=�к�;�r?��u?�M[?ӟ?��P=��>�q���'>��@��m?$�>���>Op���<��_�Za������R-���H��A��<�=�&ս��}>�:>">��=��=�ϫ=J#�<��-�A4����<��	<��=�8�=t4>�=_}q?���6��S���>�r?�2���W龄���j?�$�>��^�ٺ�=�<���?(n�?�-�?m�> ��*dp>�\����=Io%>y\=��>Vʬ�%��H��>��>������<oӯ?M7�?�?�B��گѿO��=�7>4�>�R�1��[��b�`Z�p!?\l;��_˾���>��=�N߾�ƾ�D/=$6>ֈc=���u6\���=ܧz�<= �j=��>BC>�:�=�q��k:�=��J=��=F7O>lh��X!8���+��R5=���=8�a>B�%>��>Y��>�C?b�F?��*>�c��EP���d����>���<�q=�4H�w�>=r�>�P?JEg?3 ?4��>aM|�p��>h#�>�'��Lz��T�H/���~�=��?��?�Ƅ>�O����.�+�>�.�A���?�n?�:�>�i�>���N���9���LȾ7<6����-��*�`�o32�$~ܽ��=��;�˙=���>��l>��=U8�=�|^>ɬ�>X۶>E��=nO�.�3=@t�~���}>��=p��
A�(�=��=�<�u�_������ߥ��=c0=�=�F�>���=�h�>8��=7���l) >�C����O�`s>C饾�}E��Lc�Lz���'�yE=�'EP>�R>M���2;���F?� B>�bE>�<�?�Aj?�K>7����Ӿ�H��	�E�bJT�vU�=c�=�?�3�6�y [���M��Ѿ���>z��>��>��l>V,��"?���w=U��b5���>�|�����+�9q�6?��r����i�f�Һ��D?fF�����= !~?*�I?N�?���>�����ؾ:0> G��s�=���*q�m���?~'?;��>��
�D�K�ƾ ���5�>RE���V��r��ӿ�D{�<�f˾���>1 ��F���(�����㞖�inH�I������>�a?��?�f���L0Q��G
��3���U?�W^?O��>���>�D?��;L��.t��at�=(�t?c��?8#�?:��=ڥ�=n��w8�>�,	?ƿ�?���?^�s?�|?�rt�>�(�;Ƿ >�ǘ��J�=a�>鈜=��=�q?�
?(�
?�j����	����O��^�=o�<�ۡ=���>>m�>��r>��=^ug="v�=�.\>�ٞ>d�>��d>��>PN�>R����
(
?���=t6�>�>�&�>�{a�.,0��b >�>p��@��J�p�Q=ܘ�=Gf!>>ż%� ��ý��>F)ƿ�ڰ?,�=�Y��:��>W���CVD�\\>��̽�^����?F�>���>��>4?U=D¶>C2�=��ﾙI=ը����5��>�/Z��B��H�>�$����#�����`���)�+�l���1�A�d�ʪ��H6.��)>>���?Mc3�B>K�D�M��Y��c�>>
�%?S�����f�>� ?��>0���}V��󷎿�����B�?�n�?�c>wT�>�X?��?�82��4��Z���u��A���d�@=a�𩍿?J����	�Jt���`?�$x?9A?/z<�z>�[�?VO%�>���z�>)�.�x�:��zO=�
�>ջ��}Aa�5�Ӿ��þ�O�i�F>9�o?ȃ?� ?��U�����4�W>�%]?��G?�b?�x?O;?�����2?��_>��
?H�?��@?q�?^��>�L=G�=�Hy���W=6�|�����<�M�ý�<B�n=��R=���{�:<*f�=��+=�)���G�g���s�I�<L�K=1��=^cZ=o�>'Th?�e�>��>H_ ?�����>��sܾ{�0?1h
�&���Xn������ޠ�WX_=L�F?!�?�:S?�J> �A�����>�D�>_->�W>�2�>W��4�)�T�����=2;>���=:����Yc���Q���$f=c>}��>޾s>�L��6]> ؾ��G�!��>��O���޾ڬ�k�d��N�Ќ#��+?UvI?y��>��=� ��S߼��u�QL?,� ?Ʌ^?.��?��������v+"���h��J�=S�?V/�=NuA�п���|�5��C >�$p>3��<ҥ�B5Z>�Z�ݾ;�q���K�ý�`�=�<�U~`=q���dվ�{��=��>��%!�OĖ�1����EK?�Gh=�����Z�B����l>���>��>���)O{��=�*���{��=u��>�0>zᐼd9�
H�0���X=�>;+E?�[_?�h�?pA����r��B�	��������ʼw�?�2�>�Z?S�B>�Ϯ=V����}�d�4 G�c�>�_�>O���G��&���%����$�"ϊ>(?�%>��? mR?��
?
�`?�
*?�J?��>pҸ��޸�^K&?���?�jz=e罛O��9�m�A����>Ԟ'?&Q�$��>�y?��?
+?��U?��?��>R���9���>mV�>�;V�����g�k>��K?[��>��\?߆?��L>��4�)���io���=�Z&>�3?�?(o?�!�>ߨ�>ԭ��O�=l��>tc?{0�?#�o?���=��?�:2>���>���=қ�>Ԋ�>�?�WO?�s?r�J?P��>g��<C7���9���Cs���O�2��;@yH<L�y= ��p/t�"N�<��<Q�;�g���I��o����D�����J��;��>٥_>��¾s�g>ԩ�d񧾯R[>�_<�]����Y��e���=>���>�	�>NDO�3�=���>T��>�-�w�^?v5�>I�)? �>DOR�S��7M½�C�>&h[?�[>5c��U���!���hW�<܎I?�(B?)[������l�f?2:U?���5,;�������'>�F��`?Vd?P�����>H��?&�N?��>~Щ���Z��o}`�w���c=��>?����9����>��>MP�>��>S��=�8L��Ea�Ǚ��u��>�o?a��?���?.�G>Y�����꿟���`J��^?փ�>vH��N�"?�m ���ϾNR��)�����������>���s���$�.݃��׽��=?�?ns?�[q?��_?� �ld�E2^�U	���iV�E&��#��E�N&E�όC���n�>_�Q0���!��i�G=�a���?���?Y�&?�8j���>Y料����35>�����
���=���6�=]��=�A�[�ݽ�W��9T ?��>$`�>�;?��_�@�/���:��*�����i>Q�>n�V>� �>�P�=��ܽ|�	��Ļ�������o�m>�9b?�AM?app?%��?�,�q*}�ND!��?�#(��XR`>�1>�ˎ>��Z������$�D�8���r�	:���������R�=D-?Dm>Ϭ�>Ar�?��?����5����X���2���=���>m�a?N��>[�>�}��?� ��H�>y�l?�i�>3E�>Ę��k:!�V�{�gʽ���>�>�|�>Fm>�d,��\�(<��.���19�v��=I�h?[j��:Pa�ձ�>-`Q?�a�:��L<�ߢ>myz��� �E�'�+>�g?���=hP;>GLž��6N{�5X��6P)?XJ?I璾1�*��5~>!"?�|�>*8�>"1�?`&�>.vþ_NO�B�?��^?]EJ?/YA?XG�>>�=����^7Ƚ@�&���,=�|�>W�Z>�Dm=�|�=J���P\�1i�5�D=���=�8ϼ�����7<+6��5K<���<��3>E]ܿٶH�UEѾ"D�	u�-l�'G��7��������v��t�����{�Gw�J�
�t�O���f�S�i�r����?Sa�? o���b��Hl��E�~�5���a��>�h���2��ޤ����^Ɠ�H@۾�X��T��6KQ�}h��i`�֒'?#��� �ǿ
���R<ܾ[ ?7A ?�y?����"���8�Ҷ >k9�<p(��*�뾏�����οܦ��\�^?���>��<�����>���>O�X>�Rq>S���ힾ8?�<��?.�-?��>̐r�ǕɿY����$�<|��?��@cA?��(�S��i�U=j��>Ƞ	?�?>�1�i=������K�>,=�?���?� M=��W�+�
�9ge?�C <��F��o޻m5�=]�=F�= ��0MJ>�X�>�w��VA�r�۽��4>U΅>E#�ř�AO^�ᐿ<��]>�)ֽ�㕽g��?d\�O�e�ά/�@��t>�uT?�Y�>0-�=�,?7iH��WϿR�\�`Ja?�?���?��(?MQ�����>GEܾ��M?��5?�A�>h�%���s����=�.ϼ�<��e� �U��b�=���>3�>A+�����O�f���H�=#�m�ſD#��L �)�<��%�4�a��3�t뫽ӝ_�A��
^p�p��p/m=J�=�kP>�|�>+GR>bmS>�{W?9$l?D
�>LJ>����芾�8ξ�YI��q�p���,��f'�7��� k�ޡ�'��U���j��Ⱦ0=����=RR�C���2� �|�b�n�F���.?<c$>T�ʾ��M�]"-<fuʾ����N���[᥽JT̾��1�0n�f͟?{�A?�녿�V������46��Z�W?��R���ݬ����=,����w=+ߜ>��=����3�fLS�81?�!? ݿ�����v>��ؽ��1=��0?#9?�Z=���>�n)?n6�3^��whZ>� 1>R��>[��>/D�=�=���R㽛�!?��T?ڊ*������Q�>�s����|��B=�>_�1�҇7���[>�^.<.���!K<L:X�+�*<�Y?���>��,��>�N<�v�>Ɍg��6�?�?k�=��g?�e�?��=G7��.~���!���R��Wh?�͛?h�d>��09��#���'?Ks�?uK�>������U�)�������>��o??ª<�ڄ�֢���~��?�v?�x^�7p�������V�x9�>p�>a��>�9�>m�>?�##�BF��洿�hZ4��Ş?�@���?�<<���.c�=0?Fd�>YO�1�žN��>���ahs=@1�>6����~v����,/,���8?௃?���>DĂ�u�����=�ٕ��Z�?�?�����Cg<U���l��n���~�<�Ϋ=���E"������7���ƾ��
�����࿼Х�>BZ@V�r*�>�C8�Y6�TϿ$���[о�Sq���?6��>Z�Ƚ���9�j��Pu�`�G�8�H�������>&��=8��~���{�˿<�e�`��J�>B왽��U>s��Ѿ3��w��=d��>�>�*�>Eɽ�J��Q�?��6�οz���"��I?� �?ev�?҄&?�!g��n�ş������F?�m?�y[?��E�����9���j?����g`�Y�4�j)E�2�W>�2?]��>�D-�e~u=�&>L��>�>�/��zĿ�嶿�G���Ȧ?�z�?�A����>�C�?�M+?�/��3������3�*��yعXjA?�1>����-�!�

=�
9����
?�e0?Q\�V���g?O�t��+}���A�=���>B�u�*4��:<� �<l`^���ƣc�q��?@�@�լ?��5��a�=�?�s�>��)ž�->��>h]�>��=��-���)>h���d��5>�&�?�� @�]?ѣ�L����Zk>�j?���>�e�?}h=a�>\�۽�Lڽ�)=���>�*>RJ�=�?w?�5t>VC�ӿ������i��y�~;\��\D�uY�>��?��I?u��=�^��*�j��32��f���D���4>�b�*��=�7�֭>"r!>�$�>��׽�|a��v?��ؿ1���̀(��#3?�Ԅ>�@?%9���r��K� G_?���>}���o��� ����n�?�4�?F�	?�OؾR��� >�c�>Tʆ>P0ϽL�������9>�B?X��$����o��C�>��?��@��?P�h����>�:}�)<���>��oD�Wɀ>��8?��Fâ>D�>[ >QPj�(䟿�;���?�>�s�?�0�?�a?@{?�Ee�az\���=�?�>���?gM�>qbr�����M��>n� ?l^4�F덿j��R�}?N:@w>@a�R?A������n���[���G���j^==��l>�f>�}��<���>u����Ӽ~�>�Ҏ>f�\>o8>w��=&�,>��
>J^�� \ ��T����S*����]c��9��w�	]� ������⋒�K���2K���Xѽ�l����A�o-U����=|�R?j0V?m�s?r�>��S�z�8>>����,4<�G%� >O;�>O�2?��<?��"?.�B=�׌�4pd�e+��]�������e��>qf7>���>`2�>��>��
=2�=��=���><6�=T�=BL�<�l�<KOC>�>��>�\�>�C<>��>(ϴ��1��@�h�w�s̽/�??���:�J��1���9�����j�=Zb.?�|>���?пF����2H?����a)���+���>m�0?�cW?�>l���T��9>s��Z�j�*_>c+ ��~l���)�8%Q>Ml?��i>d�x>�)3��I7��LP�.A��i�|>�+7?�״���4�>1t�W1F��ݾ�J>�i�>�X2��m�d;��e��̩k�'r=O�:?T�?��Ľ�@��r�s�����O>(-V>�{)= a�=�RP>�D_�ʽ%`E�j�A=R@�=N�[>^H?�G,>�C�=Z��>HV���DP��E�>�sB>ջ+>X @?%?@��k#��������-���v>�%�>-�>?>-�J���=��>_�a>�}��Ѓ�T��X�?��W>��~��A_��uv���x=Q̗���=Z�=� ���<���%=��?�*��I����;~��>� *?�??;�[�R�����O��&���)�?�E@���?<��~F��`>?�9?����>�,�>��=3� �p����1G?p��Pt��*�w똾ߚ?
+�?!���jl����.����=��>���=_�>��O�¸���p����n��.߽
��>+L?�����ؼ�3>�jH?aM�>�ھ�F��Q�ÿ8�{��c�>j�?m̚?Jr����c�2�2^�>�r�?�0f?��n>��:8�D)�>L&?��6?�x�>���:��5;?���?r	�?I>��?Ӕs?�n�>��w��Y/�*5��"���3=wh`;�W�>�3>����ogF�bՓ�i����j�Ľ���a>̈́$=�> �n:���Q�=t���A?����f����>�q>��I>�U�>�� ?i`�>ʡ�>�\=���N߀�F���m~L?e͏?���k��4=+#�=>X�3 ?n.3?��<m(ʾi��>��T?�oz?�!X?���>|������Y2���ڳ�·�<E�a>Ѝ�>���>��ýY�O>#�;1�D�_��>�6�>���aSپW�z�IŢ;���>�� ?)��>��J=��?�4?��#>�Ϝ>�I-��a���e���>�L?C�>_V~?�> ?9̾�:=��������F����>~?j�)?]�>ɋ���H��[=T�P>yν�?�I?gɪ<��*?K��?�Z?@p'?�L>f�/�\����o�i%�>�!?���Z@��l&�	���?�?W
�>�|���߽�F�ܖ�\J���I?��]?�r)?aY�@a�ϊ�����<!��9�������̻��">o	>
�b�9�=��!>�	�=�b��yB��C.����=/z�>���=��8�[���ep?ě�=����B5�=k�m�x#E�s�:�>�L��"?� ���4i��Q��H�������V��?���?���?��E���f�,%8?�s?��P?���>����%�׾� ��Y���7�2�-�~�>>L��>���=�_߾U��ޘ�����М�\c�=C?Ze>�w?�?���=}�c>4⋾ c5��������r���A7�! �E/�x�ӾMA�=��>v���:`��P]�>�'�s�>�7�>I��>��>�>.�ҽ�.�>ӕb>��>R��>�.:>� >�-�=9�C��nR?^Z�by?�8�-���<3?�?ZD�>�č�� ��n�&�8F'?��?֔?�r3>��b��..���?�d�>����5?�h�=n3>��N��o���0;�=�}(�/��>h�^��a0�Kwu�i�¾0�>y�>Đ�<)7��,})�2���Y�n=�E�?��(?��)�6�Q��o��W��S�����Uh�-Y���$���p��叿CV��s&����(���)=�*?�?����������k��?�ƴf>��>'
�>�ʾ>c�I>��	�R�1�y^�FI'��΃��8�>qZ{?-Ռ>�gI?3V<?/�P?kL?�g�>¾�>ူ�z�>�#�;��>$�>D�9?�-?��/?��?�+?�Y_>�o�������5ھ?3�?�R?N�?�t?~8���˽p��>�3���{�^x����=���<׽^�w��V`=8�Q>ܞ?�8��5�;�*��*�\>�]T?�,�>��>/�~��"��{O===1�>u�?7�r>{i	�U���Q ���>J�?P	޼�0��5�=$>�����.<�c�=o����=�11�L��-7�w�=ꎨ=��=o��6Lj:KQ���PK�p�>�Z0?�b>̻�>�S�6#���|$���ϼ���>�l"���>�Ⱦ�ᎿZ���:f�Zaj>�h�?Ҵ�?�7=z26>��>�Sž)� ���������l!1?g#?J�Y?qB�?8�[?��.?���=]i�Ew��>��>;�V�6?!,?���>C��G�ʾv憎�p3�ݚ?�j?�a����0")��I¾�!ս~>GL/�3~�}���#D�aϠ�����0��?���?�.C�G�6�wg辀����a��zjC?�L�>�N�>2�>̭)���g�L�K�;>���>�	R?M(�>-?K?O�{?Rw[?�#A>�8�u���4͙�d�l�>�;?u-~?��?i�z?h�>"x#>I�$�s;ܾ�(�����j���B����R=�U>���>��>�]�>�=��νk��HFU��3�=��v>l�>$�>x��>'1`>�V�<��@?���>�K����O�|����,����Ľ
G�?��?�6?
�H�,�EN���E��ߕ#?��?�ޠ?Q�>I�޽�,>=��>;Ѫ�Xl#��KD>Xă>Z�=�1½�b>��$>*�;?�;�>�0���,b��L\����KJ?
dV?�M�Q̿��M�>	��;7ժ��S�r锾;��� M��=%��O�&�����4�ZB��#�x��վ�O׾�ʗ�܃?�1)>�>��=yW��c���=���<j�9=�j�=�������=��L�E�i��qS�D`a��l!�������<��ľY�3?�я?)?K?�w�=���>0菾���<��=�
v?k�=�j>�Ծ�q�5�f����P�=�&�q��}����b�H��=�i�m�>_(�;�ٔ=kV=�=��=Pz½�1Ͻ��6?�<K
=t�=�Ӄ=Q�>��	>�>p?Q��h���.a�/W�<��9?���>���=�t���g?c�!>�ꆿ�ݰ�?�
�`Ek?x��?w��?J��> P�b_�>L�������zr>v�D=8t�>	��	�U�M�>J�`>�y#�Щ�~���v��?��@�#F?�]���<Ͽ�[\=�7>4>��R�:�1��\���b��wZ�
�!?9E;�?>̾I3�>��=�-߾v�ƾŚ.=��6>�#b=�t��X\�WΙ=��z��0<=�l=nʉ>��C>3{�=s9����=+fI=���=пO>	�����7��=,���3=���=X�b>X&>��>A�>��?��B?�"u>�x��<�þ�}�%"3>i�����>G7���=S�?��Q?4�h?h�0?�N>nG>2e�>���>9J�Pw��3�}�ج|�z<�= ��?��?"#�>@�}�x�	��22�t;��gW��G?��?�>�_�>��4�׿L��*3�~]��T��E�a���K�Ž/Y�=�>���!�B�=
�>m��>ߙe>���=_�=���=g=�>L�|>L^�=��#�|���+_��%�=,��="w���6=��]���ӹ8�G�;7E�<:U<F��;�)���=5�>���=d�>�=�񾾹��=�>��g�J�v��=1���f[G�h�`�*�|�s,���N�\�F>=�>*��\;��b�?�i>�?@>��?�^n?B!>?��0��)����?q��Cp����=���=z�5�l�;��a���C��Zľ�d�>�+�>��>3�s>��*�~|?��4o= �I8�kH�>�؏��C��a��-p��̣��J��-�g���Z<O{F?}4���W>��|?	EI?o�?y��> ���tԾ~-:>ăv���.=T�[H~�������?~0$?,��>���^A���˾;nǽ��>-P���O�˕�F�.�!X������O�>�'���̾tm2����d���=C�@�u��N�>Y3Q?A�?}{f�g��0�N�53�r�^��?�Ef?lМ>�?��?jƨ��x��ځ�0��=��n?��?ɳ�?�!
>��=��D�>b0	?۽�?ݴ�?d�s?�?��o�>�?�;9� >����j�=�>F��=��=�q?��
?��
?yY��"�	�s��V��}^�Z��<c�=H��>EZ�>�tr>B�=UCg=��=^6\>1ў>8�>��d>2�>6F�>�2�������?�>rً>�Y�>��>����dW�f����v7�s�Z�JNӽ�w���)��X<�A&�̭�>�Q�=Qq�>$�ǿ�]�?�tE>~E,��>�~��"�Y��=�i<�����	?��=�&�>tP�>�?�H�>���=}��:�������=��޾�9��W��in�A־?�~>������̽�	�΄��g�_�:,��a����Z�����/�O��?=�ȗ?R�`�d|[��(�>�z��{�>�6�>�oI?��������&>�?�>(�ؾ���\���*Ѿ���?-U�?�l>`݁>��Z?X�?9u�'FK��U_��xx�N�I��d� �a��g��ٝv�x۾o����Ma?��n?:):?���<�G�>��q?�{(��ȉ�d��>ʬ)�?�4�Cn�=�4�>�n���YI�V������q����]>�q?��u?&e�>R�?��ѽ�dF>8�L?RB?��c?�R?HfB?�>:�0R?MW>��?c�>z�.?�A?M��>���=J�>{�p�煀�%o��ES��ѽ?�强�1;�,�=� =i�`=�L�=@���z�;s���J�������;��==�@�=�Ϫ=�}�>0Ke?��>c"�> 5%?��X�9;>��,뾲@?1J��܊�T���[���5���h=D�U?&O�?�+J?��>G�@�ɵ��m>���>��l>�>��>M���祽\����=�'>��=,-�;��F��l�n���	آ=o�Z>�n�>�t~>�����2>�����΁��a>n�Q��ƾT�F���H��2�+�p�N��>9qI?��?���=k/۾��S�a�f�]m/?��:?WM?۬�?��=�澸#5��C�a��u�>9�C*��֣�Qc���P:������}>/Z��࠾�Tb>O��s޾#�n�"J����9M=��Q_V=����վ*4����={$
>����D� ����֪�D2J?Z�j=�x���gU�Kp��q�>"��>=�>��:�1�v�~�@�Ϭ���1�=!��>X�:>0a�� �<~G�*7�G7�>mGE?BG_?Zj�?����<s� �B������r���(ȼ��?FO�>�^?�A>%�=f��������d�*G�7�>I}�>$���G�
1��/Q����$��X�>�@?�u>�?ֽR?��
?u�`?�*?�M?�9�>�����Ը��B&?<��?�=��Խ��T���8��F�a�>4�)?��B����>;�?v�?E�&?�Q?��?�>į ��E@����>�Y�>�W��a���_>A�J?���>}=Y?�ԃ?�>>"�5��碾�٩�EU�=�>7�2?�5#?��?"��>���>����qO�=n��>Nc?Q/�?n�o?�q�=2�?#2>U��>��=Ҥ�>��>h?�OO?��s?��J?���>M��<���C$���Ns���O�9�;�I<�y=f��(t��o����<�4�;�����s��F��<sD��ѐ�p��; P�>�Et>�̕�
�1>E�ľ+�����@>�s��ࣜ�Ώ��|d9��S�=��>e?+��>t�#��ڑ=�=�>�(�>q��P!(?�r?��?�W
;�b�T�پ��K�}E�>j�A?���=��l��I���cu��j=�m?�]^?�<X�����e�b?!�l?� �)O��9 ���
���߾;g?�w??�U�.њ>�v?�8r?��?g,���i��M��ɇw�.؃���g>�mD>T5��w�3/>� z?��-?Q4?� >ۣ�i��R���)?�O�?���??ř>=�`�����h���B��/^?�~�>�����"?6��m�Ͼ�j��k#���*�O.������I���\��8�$������ֽ�м=��?��r?�lq?�_?� ��d�&^��
��LeV���8�d�E��)E�}C�8�n�M5�4��[혾'8H=�j~��\A�Sn�?ߗ'?��.����>D���񾶜;��B>�*������B�=�4����B=tb]=>�f�,�-����{ ?�5�>�=�>AO<?L�[�e>�ku1���7�����4>�l�>��>�B�>� ;�-��6���Ⱦ:փ��6ҽ:Lv>�tc?6}K?��n?^�'1�?�����!��0��Z��X�B>5�>�̉>��W����"8&�X>�0�r�����|����	��~=I�2?��>���>�L�?��?�~	�
���vx�d�1�A�<�3�>�i?�(�>��>3�Ͻ�� �E,�>�Wr?}�>���>�ԾzC��⍿��Ի,�>�Z>�?Ø�>_X��[��@ ��|���/��g�w>��[?�����Ρ>�L?���=�.=��=-φ��6�a�9밾�Ή>�E?�'�=�1>��\9��8���ޯ�mZ)?�a?3��m�*��y~>�K"?���>�c�>
!�?b�>�kþG�:�?a�^?�J?�-A?��>��=Ђ��k{Ƚ۰'�.i,=R�>�Z>��i=���=
��+l]�	��xJ=[,�=V�̼�ٸ�u<�e���+M<o��<��4>�
ѿ��<��������-��$���@5���ս�둾/�ǽY������k�L��_q��W3���q�:�y�k���M�V�C�?���?{�徢1ľ뭎�0w������S�>����S�����ξ���;�#���
ݾ\轾-g ��_��ue�p�F���'?�œ�Z�ǿ�b���DԾ�?`U"?&�z?���x�!��N7�R(>jQ=�0�3x�����(�οǥ��w�c?q��>�����ýK8�> Ǝ>Ec>f>@���M镾��<�?4�-?���>Mr�{Nȿu��z��<���?��@q�A?�'����\=D��>�D
?��6>H�-�ݿ��Ů�K��>0��? ي?��W=��V����>c?�P�;��F�������=�'�=�(=����F>�#�>ɦ!��8G���#(@>(��>���:�,�\��Қ<��\>mȽ;/��$��?��i��Hy��A0��ߌ�Ӑ>�k?c �>?p0>"�)?Qx�1uӿ�>V��jo?r�	@���?h??�~��އ>\>����t?P-0?0�>��P�_K}��q�>�>ڻ��R-����V�ީe����>��g>�
��b-��#W��*=�% >��ɑſ�"�q��V)�<�����HJ�H���ܴ��N�J���ӯt�x_�T��=e��=��L>Lm�>$QS>(�Y>?�W?�zl?+�>D�>�0������Cɾ�v���⁾�j�/��������_�뾇{޾"	�s4��=�PYȾ,=��ۍ=`R������ �r�b�_UF���.?��#>��ʾy�M�:�+<�Gʾ�s�������H̾˓1���m�2�?�B?��W�`��eP��*���W?�������&����=M䱼��=���>ۛ�=m-��3��BS�.�1?�F?۾��T���&>�l�;��ؽ�"?�U�>��K<dM�>l4B?:�$�a=�s^@>4��=�W>ﱸ>?��=�R��HU&�{s?��S?uis��׏���>i о ���X9�~��>��|���<�,{>ޯY=L[��ЂQ�2<�>W?�-�>��)����65��/�'��3=9�x?'Q?�D�>x�k?7�B?�
�<���PT���ϼz=&X?\�h?V�>����cϾ�0��<5?̤e?V:M>� j���龟�.�'%��B?�Ro?&5?�ɖ�,�}��Z��%y�͇6?	?��m����;���|=eE�>���>LN�>y��b��>�-7?������9G��)�@��Q�?�@��?W��|� �y�<�Q>?��>���nܸ���$�K����?�<�X?�٫�����V1�Dg��F_?7��?�?�R��>A����=�ٕ��Z�?��?}���,Dg<S���l��n��E�<�Ϋ=���E"������7���ƾ��
�����࿼̥�>DZ@�U�u*�>�C8�\6�TϿ)���[о�Sq���?N��>U�Ƚ����@�j��Pu�b�G�4�H�å���L�>��>����}���A�{��p;�(I��1�>��� �>��S��#��W���5�5<�ߒ>ʩ�>b��>�8��⽾�ř?]��d@ο����Ɲ���X?�g�?�p�?"n?'�8< �v�܂{����.G?��s?Z?��%�|=]���7�$�j?�_��xU`��4�sHE��U>�"3?�B�>T�-�9�|=�>���> g>�#/�w�Ŀ�ٶ�>���Y��?��?�o���>r��?us+?�i�8���[����*�'�+��<A?�2>���G�!�A0=�PҒ���
?W~0? {�e.��m`?P�b�hr��.�lQ̽Ȕ�>� -��a���޲�f���E5����?J @噳?*D���!�Q�#?B3�>�����ľK�<x�>���>�`>c&R���z>���&=����=��?��?��?�`���Ҧ�hz>�}?(�>�}?j!�=�g?b;_<�娽�':<��(>:�<�)��~??�?e?��?P��>K���İ.���9���D�e�ƾ.�F���>�Ɔ?ZvH?��]>���4�x>� ��њ=�{��|Խ�x��
=%��5ta>t�>ߟ7>�`��^���t�.?��.��]ۿ?B��ƹ5>l�4?�>�C�> &վ`h�i3C<��b?7N�>��𾅗������� ��B�?�k@��?��
,;�Q��>\`�>fT$>��g�0�B��<� �>djB?8�D�h푿N�����>�
�?#@<O�?�o���?�b�O��hd|�FW��,�Eu�=un5?����Q�>� �>��=�dr� ��g�v��е>&N�?W��?S�>sj?qo���=����= �>%�a?��?�7����㾤T>��?Yk�=���+��I�d?؉@��@�EX?A���Y�ؿ
њ������ܺ�ء����>��=��վK��aq�=&�=�#/�M@1=`��>�9J>�F�=�(�=m�4>�@[>�����)�����O2����+�h��3J"�X���=��žQ� ��a��ξ}��ҷ����}�2}���ӽ������=��\? V?��?=�?�u�&~>b�ξy��=�y�ǫ$>l��>�{E?-P?U�"?���p�����o���m�����/�h�	��>�|)>��>5�>��>�䢽\X>4m�>�5�>��=�U��I ҽ�=Ż6�H>��>H��>���>=F<>p�>ϴ��1����h�w�2̽��?�}���J��1���7��Ԥ��t�=\b.?B{>��?п����2H?^���n)�ֺ+���>h�0?cW?B�>���ֲT�R6>Ӿ���j�`>�& ��{l���)��%Q>yk?Ϲf>5u>@�3�-H8���P��s���c|>�6?c����/9�~�u��H�"Uݾ�M>�Ǿ>(E��]�B���/��di�B�z=�:?e?��������u��k��NxR>��[>�Q=���=LM>�5b�`�ƽ��G�F/=��=)�^>�%?��+>9��=�H�>�E���;P��2�>wJ@>Q�)>��??x�$?�!��%��������,�U'v>��>���>�>�I�g��=��>�_>��o�������B�R�W>���� �_���s���v=����B�=Zh�=�m���:�f�,=�~?���(䈿��(e���lD?U+?_ �=/�F<��"�E ���H��F�?r�@m�?��	�ߢV�@�?�@�?$��`��=}�>׫>�ξ�L��?��Ž:Ǣ�ɔ	�.)#�iS�?��?��/�[ʋ�>l��6>�^%?��Ӿ�[�>�t3�2������e�L��,�=\d�>z�\?!����	�D�ٵ?C?|������¿����U�>�?��?-�����j.��W)?���?C9?��=:#���.��>i>+�E?c8O?4��>u�$��8�ĭ?��?���?��F>j��?��l?�=�>�r~�چD�{���H���2�=�m��4Nv>H�Q>�۾�Ad��i��j����Ng�}�G��>3+=dй>I&�.�о@!>f�@��װ�b*彲��>��>@��=ͽ�>��?��>��_>!��-�1y��Y�8�2�V?3d�?-/+���~���Q�2�	?'����i?Įt?k[<Š���?�[?��r?��I?��x>6�!��~U��Μ������1�=0�?g
?�cr�"�����3%پ�0?�ʗ>�d:>���J⯾��t��Bl>Q�?���>�>�a?�z6?NHg>P��>�t2�Dk��U�o��	�>��?X֤>�^?��?�K���F��䜿ꅨ�s2l�5�=]��?A�%?w��>Ǽ���Z��� ǽ[�~>��=���?wn?I�o��z?,6c?�8s?=9f?ɛN>߂<��O ���V��p#>P�!?M���A�{P&�p���?�P?���>�󒽻ֽ"�ּ���Tt��?�(\?`>&?����.a��
þ4,�<��"��W�"�;]D�J�>-�>�q��K��=$+>5��=�Gm��G6�I�f<���=���>��=�'7�����,?j��]Ƃ��g�=�.s���E���w>��P>�`��G^?n/6�c^z��謿����Z���?�+�?Kܖ?�����	h��<?��?��?8a�>FB��\�߾z��*�w��Wx����:�>��>�1f�I��IŤ��F��ʄ�V���������>4��>��'?-.?�@>U��>���imL�S���'W	���g���EP�ۉ�b��S����W�l)-��Y���"���\�>�P.�<��>��>��O>��=<D?�y��@��>?I>��>c)�>��!>ҡU>�MJ>�O<\���w0R?����'��������xB?M�c?���>��m�W��������?��?�d�? Bv>�oh�K-+�W0?z$�>ΐ����
?��E=���@r�<�r��4�$[�����+R�>�oؽ�/:���L��Qe�t
?��?#��b�̾~&ֽǊ���o=�M�?<�(?��)���Q�%�o�ȷW��S�����5h�<g����$���p��쏿,_���$����(�4�*=q�*?��?	��ߖ�C��&k��?��]f>�>U!�> ۾>�yI>&�	�:�1��^�WM'�����3M�>�[{?<��>O�I?��<?%-Q?,FL?D�>B��>�J���u�>�|b;B��>���>E:?��-?/�/?��?�B*?�\>X-���d���y׾?�?��?\?�?��?����ƽ}����B���y��+����s=iP�<�vսlFm���V=�uR>�Y?z��8�����j>�7?�X�>f��>'"���3��2Q�<�+�>%�
?�R�>�����yr��d��M�>�?����{=J�)>p<�=+�����ͺ��=��¼S��=<2��Ԕ:���<q��=�#�=R�l�o�����:UI�;�ʰ<��?�W+?}*S>z<>����
,H�_�!��@�>9�i>�W>ɣj>f���g������R���B�>T��?��?X�X�1��=��8>����=��s��fq�,С��1�>��>�p@?��?b+_?Z�`?~�t��q	�5%������h��M ?e!,?��>���ղʾ�񨿄�3���?J[?�<a�}���;)���¾s�Խ��>�[/�L/~����D���������~����?保?�A�-�6��x�̿��	\��)�C?}"�>�X�>��>L�)�N�g��%��1;>���>R?���>�PO?��{?w@\?�"W>ɺ7��ѭ����Gd���!>ڍ@?���?��?n`x?�k�>M�>2*�E�߾�E��a(���&Z���N`=��Z>~%�>���><_�>	��=�н�٭�C�>�p}�=`ha>��>� �>�O�>t*z>� �<=?��>��0����}o�`�r�m�n?�͇?�w�>F�v��
.��ꐿ�h��T>��?�V�?��Q?zƾҨ�=�$>T^ʾ�-�����>��O>�Cz>�>�q=�jy=�S?(��>nć�r>&�;,:��4w���?��V?��=�?ƿ��s��7Q�쇞�� �&��C'S��Rｷ�e����=
�~��<3�����&��7[��V���嬾V���CP���>�N�= ��=f5�=D_=�7¼��<��u=zn=(�=(���� =�r��c:�5��FP����<C�=Ŧ���&����u?�1g?�-8?��J?��>&��>�����a>�m����'?�Ɯ>�Ω=�ʭ����,��	f��7�~ʾ�6L�N��Hp>�r���&>g�:>���=��;=~"�=E�=�!=�׽�P<��=�0=1~�=Ef�=�&>S.>�9�?'��ҡ�	�6��Bd=�	=?��>>%E�;�o����k?��=
���᯿�'���?~�?��?��>����`y>}�����W���ʾ
�>p�=����{Uj>��==L@�����CQ����?s�@ 10?�5��M�˿抋>��7>v4>�R�9m1�Sg\�pb��Z���!?�O;��,̾�+�>��=�߾3�ƾ��.=�_6>�b=�~�IV\�i��=`�{���<=��k=vω>e�C>ǃ�=����\�=VhH=�r�=U�O>$c��2�6��3,���3=I�=�b>�,&> ��>#5?P�/?�wc?v�>�@t��ϾО��@ċ>-C�=�>x(u=��9>�ط>K57?�F?�L?�z�>�z=u{�>���>�B-�ghm�=�㹨����<F��?���?�@�>bi<��A��� ��0=�E*ʽ�?t�1?�g?u-�>c���ɿ����Bi=�zN��asB����Yi��v�+DN>%#<O,����=䗸>�'n>��=4.�=�p0=bk�>{��>��>	Z=Pd,=�'�lK���>��C>���=��=M�=?D�=�z=^I�<9<(<�<)��<�?4�r�.����=���>���=#��>
K�=���D0>Q���a��� >���%F��_^�S������i�M��,>�@>U��9�����?�n>�wd>�o�?�Zj?;�=e�+�`ھ9Y��w��H/7�
��=�=�K��|?���U��GO�@�����>"�>���>��l>
,�A?���w=��j5�J�>��g���$��;q�Z:��R���i���պڙD?NF��b��=�"~?��I?q�?P��>w����ؾ�30>.H��=Q	��q�������?"'?���>�쾲�D��G̾���߷>p?I��O�����0����>η����>�����о$3�pg��K����B��Ir���>f�O?O�?U<b��V��cUO���l-��q?[{g?�>K???�#���z�wq��gv�=��n?^��?=�?�>d�=�y��b3�>W�
?Ж?�E�?��q?/�@�:��>�<�;��&>������=iU
>��=��=�;?k�	?V?ܾ���
�]Z�4�TZ���=7ћ=�̒>~G�>��i>'j�=Dd=6��=�Z>L�>�B�>u'g><1�>��>���"���Hl?�3>�I�>�?2{�>���Z$���;���)H����*��^��ob�4��<��b=��&=`\x��o�>4�����?�V=���Z�>�޾��+��J>j�E>�[\��0�>���=��>�S�>�_�>4�L>�(�>.c>�T���{>���9*6���?�8,D����<ʬ>��;�e��7�"����*�
Q���)�}d�� ��Of>���=�=�?��#Ӌ�l6:��;�)�?�C�>��P?fe���o�/�3=N�?4a�>�~ԾjF��#��F���Q�?D(�?e��>�6>��H?|�?��@��Nܾ��2������0@�Y/��+��0���~���@D�<��?hǀ?�g5?ul5���>��U?�i�����I5�<��)��X?�!��>e��>(��-<��%s����4�쩧�{W=��?,�u?�X?��������{>�>��?�o?��}?�Y?�@?[�b��]�>��=��B?}�?�qO?;�>W��>�ҽ�O=G�o�>��F�"~���%�;q�R�K��o��9I_�����	�(��<�=�̕<}f=��q}�b�0:4i���|<��c=|�7>� >#Φ>�]??�>�g�>J�7?�����8��c���-/?v9=s肾�D��l��*򾾉>k?��?܁Z?��c>{�A�+�B���>Z,�>�s&>��[>�Z�>xR���E����=>b�>7��=&�O�x�����	�rV���<�;>v]�>]�\>'�%���y> �]fU�7Θ>r����T��8�c���E����"�>BrT?�_?��s=�ľ��i�2�u���J?��<?�Eu?Ow�?��q<q��E�/���|�ww�����>8}*>��ݾ��������\��ꮼ��=�ž�T��j�`><=���ݾۄn���I�/[�ÖC="�}\=���־z/���=t>����~� �'���8����J?��l=MG��oQV�3���ݘ>MT�>n�>�4��r�N
@�)���,��=E�>��;>>���B7G���5�>�NE?�X_?vl�?a ��s�-�B�;���Z����Ǽ�?�x�>Hk?�B>G߭=e�����{�d��G�A�>���>��X�G��;���/����$���>e6?Ȥ>f�?s�R?��
?�`?�*?�A?�$�>����񸾆@&?Ć�?��=4ս��T���8�zF��
�>&�)?��B���>Nz?c�?�&?��Q?f�?��>�� �V=@�I��>�l�>$�W��`���`>��J?ߏ�>?Y?*׃?��=>Vz5��~ ����=�>b�2?�3#?ݦ?Y��>y��>P�����=Þ�>�c?�0�?�o?���=5�?�:2>3��>��=���>m��>�?TXO?6�s?��J?��>���<h7���8��dDs�K�O�vɂ;�vH<h�y=����2t��J�&��<���;�f���H�����D�v������;}��>
�k>|퐾��+>�jʾG���K�E>�P¼Y���σ�M�J�6Ӟ=�Fu>��?`T�>ή�<m�=��>���>C����)?~?��?���_���Ҿ�}2���>��@?��=�|m�����r��q=��m?�]?�m^�P���Z�b?A7]?������;�7U���!E���߾�O?<M?Ծ9��ڴ>V	�?'�k?�8�>R�r�?Lq��Ȟ��Q`��f�F_�=���>y��_\���>!�-?L��>ʞ^>�Y�=�ɾ1r�ʄ��ʺ?ʊ?_�?-a�?j�>S�m����^}���I��9^?��>�>���"?�� ��ϾCN���,��5⾸��p��SD���w����$��؃�׽�޼=A�?�s?bZq?�_?ϰ �d�;1^�9���kV�/.�;&���E��$E�ҏC��n��c��*�������G=M~���A�3K�?&z'?��0�@��>E�����_;�C>�M�����ɝ=x0����J=C�b=4�h��,�.^��� ?8��>Z>�>L)<?xA\�@=���0��6�x����5>�}�>�ޑ>0��>�;��+�R-佇�Ⱦ6��Sս��u>�fc?pVK?Χn?"'��#1��}��@�!��#0�����B>�4>}��>��W�*t�V7&��;>���r�����f��!�	�Gw�=}2?"�>�?�>�J�?I�?ER	�3���k�x�e1�k�<�M�>ki?�b�>o��>H=Ͻ�� �/��>��l?:r�>G�>!n��uI!�
�{���ʽ
�>��>f��>z�o>!�,��\�:d������09��!�=̤h?煄���`�'�>�R?���:B<8��>Դv���!�x��L�'�~�>f?$��=�;>+bž."���{�tg����(?Xv?����F#-�m> �?�>��>=ֆ?&��>�þyᴼ�?��Z?|�L?�E?�O�>O%�<*(���ĽQr��+=���>9hZ>E��=E~�=	�;	V��n���c=�F�=�p��g�ν���;N�����Z<�2�<g>3><�ۿ@�J�Y׾�;�a����W�����"g���P	�ͳ��e����w���D4�!V�)f�z����7i�">�?���?,�拾�̙����0��6'�>��p�D$���X���A	�\i���s߾͸��0�"���O���f�g�b�M�'?�����ǿ򰡿�:ܾ2! ?�A ?6�y?��7�"���8�� >JC�<�,����뾭����ο>�����^?���>��/��i��>ޥ�>�X>�Hq>����螾i1�<��?9�-?��>Îr�1�ɿb����¤<���?0�@�A?��(�G���WU=���>۝	?��?>�1��E� �WU�>�<�?���?�7M=��W��x�Oe?� <��F���߻dd�=���=��={ ��BJ>�X�>,����A�P~۽H�4>7��>��#�_~��B^�X�<U]>yAֽ�����G�?,�Z��/c�C#0��ꀿ��>�V?���>���=�z,?�H��BϿ��]�dVa?��?O��?� (?�ؿ��>sھ�IO?�4?���>��$�'ps���=�Ԏ��w<��⾠,S�EK�=���>�G>�)��`
�>�J�YXƼB��=����ƿG�$��~���=#�
�F]\�/�罼'��+U�|��8oo���?vh=78�=UoQ>�K�>tW>�7Z>LmW?��k?*�>�@>�佲~����;����=����-���d��urD�p�߾�	������c�ɾ<=���=�3R������ ��b�q�F��.?�y$>��ʾ��M���,<sʾ̹��o���̥��*̾��1�Gn��˟?��A?����e�V���� ��Je��A�W?+<�#��zꬾ��=nױ�=�='�> ��=7�⾰3�#{S��o0?�u?e"��������+>�k��j%=�+?�?l�x<d�>�<%?�n+�Í�[�Y>�0>���>��>�		>����?�ؽ_�?I}T?���ԝ����>69���l}�AZd=MD>hr5�����(�[>���<g���|?Z������<sb?���>�9�.q��Z ���> �=��?Ś�>�߄��Ps?m7}?�߼==�;c�_����=�B�?k?d^U>��'��}������|�O?�@�?�ň>�eU�(�þ,Z�W� �A�+?�Ɗ?�/?��l=i�y�����>��d?��v?��^��|��s�1�S��!�>n��>FA�>1�9���>��>?Wq"�]��I���XH4����?��@H��?H�-<w��\�='�?�?�>�+N�oPž�U������s=%	�>q����ov�	����+���8?���?�%�>aw��������=�ٕ��Z�?��?}���}Dg<R���l��n��[�<�Ϋ=���E"������7���ƾ��
����ῼ̥�>EZ@�U�v*�>�C8�]6�TϿ)���[о�Sq���?M��>R�Ƚ����B�j��Pu�a�G�2�H�ƥ���ˣ>>Q�S�kǒ��s�ݟ8�*eZ;w7�>(ϼXH�>�$v������`��1�Z=��>�y�>:�>#����_�����?�߾N�ǿ:���0�	�[|Q?:��?~�?
�'?1�P<pYV������OV�B@?��n?5�[?��ż�q����j�j?9����`��t4��B���[>pT2?i��>�u,�`{=e�>���>��>Y�.��Ŀ��Ğ ��ĥ?��?�����>퇜?ל*?���j_��㨾Xm*��Lϻ�B?A0>����i#���;�C����4
?�.?�^�e���j?oU������<��K�>J��>(��l`��z����=��|�{B��Z�q�ʏ�?w%�?٥�?�bK���/� �7?���>��R��o��e��<:�>m��>nN�>?�=�G�>�Z۾]�R�]����{�?�7�? e?:���2䥿@�[=�{?w;�><^?�1>=2e	?N-��-h��"!>�o�>�޽.)=��?��T?��>���=�y�.�2�g�f��f��4L�n5�2\�>�f?1m?&"�����s�w�g���鑽֝H���<��V�g��=q+���95>�j>��>�I�dy�O�?�k��qؿ~����h'���3?/P�>?!����t�����C_?R>�>>!�C.��-��(�j��?Y@�?�/	?P�׾�μ�w>��>cv�> ^ӽi$���l����8>��B?Z��C����o���>F�?߽@lٮ?vi� ��>���i��%����u��|�~c?y.?]��}ɐ>�O?p�}>���_%�����¯>|��?��?�`�>��?T���uz�	J>��?R�m?y��>���|��,�>N?B�	�Y������Z�t?fQ@0�@]�@? ��-�#>���p��7�%�2=�K���+>oˈ��D<�5=2��ca��y,>��>'�>�GY>�,Q>7�^>���=ڡ~��u ��������%=��U.����~|�����ㅾ%�������Ⱦ_�X��^����i��X�F�?�p���=�V?f�Q?��q?m0�>������>J��rd�<��"�bה=@�>��3?��J?�(?�ˀ=�h��D�d��D������B���(��>��D>y��>5��>���>ߔɻ;�I>�U>>6�>v� >}Y)=��a7o�=7`K>�o�>n��>�\�>�C<>��>Eϴ��1��j�h��
w�e̽1�?���Q�J��1���9��զ���h�=Gb.?|>���?пe����2H?#���x)��+���>{�0?�cW?"�>��q�T�5:><����j�3`>�+ �ul���)��%Q>tl?�f>rUu>�{3�\8���P��d��z�|>m<6?Q���P�8�E�u���H�͕ݾ/:M>iݾ><�=��`���~�nXi�7�|=�u:?r?P���zذ�B�u������R>)�[>�=	ܪ=�?M>�6d�ƽO8G��.=��=�Q^>�K?Bn->�Lo=���>(떾O�R���>�d;>H�'>�NA?ؤ"?��)�����$���.(�Oxp>���>G�z>>�I�fҤ=���>�Z>zg輸����Ҳ<�.�\>R|���fa���e�Ss�=�ƌ�ϫ�=aȣ=�����7���=u�?�墿�0���غ���N���z?�J?�_>���>����U����Yh�?�_@��?��JW�at�>y�?|�����>�%�>R��>$.�����8/?���D$K��&��G�����?�6�?�Û��D����M��P\>:?�K��=�>S��j��ge���?s����<���>�F?*���]�{�N�;�4�
?�� ?�.�~���9ȿ2�u����>��?�p�?j<m��Ș�JbC�'��>�!�?�]?��z>f�پ=Q��]�>F&D?9*M?��>o�X ���?iT�?ԭ�?�H>���?�s?<��>�*x��[/��3������w�=�`];�y�>	o>Ġ��gbF��ғ��e�� �j�q����a>~�$=;�>t3�51����=���UA��e�f�<��>�q>(�I>-N�>[� ?�]�>}��>Un=�c��Iـ�����`�K?K��?;��u0n��$�<-��=.�^��'?�F4?*[���Ͼ�ר>f�\?���?�[?�`�>.��7>��x迿�~�����<��K>�8�>�A�>+���DK>��ԾY0D�Kn�>Oϗ>e��:ھ�+���ע�GE�>�e!?ҏ�>Ʈ=
� ?ĝ#?rj>��>	`E��6����E����>���>�6?��~?;�?�۹��b3�~	���㡿Y�[���N>��x?�Z?(��>�������.BD�XIH�習�,��?Z]g?��?<�?T�???�A?*'f>o��.ؾ����>�� ?ǥ꽶;6�|j+��M3�l�>[q?}��>+��f:��G��*#�wZ���?�8a?�0?*���3c^�c��a�<���<n��.��� :�">��=W�n��=��>֏�=jPr��h9��3��t��=���>J>�=r!A�+p��<,?l�G�Lڃ���=b�r��wD���>&LL>� ��b�^?�l=��{�����x��	U�!�?���?�j�?����h��#=?��?p
?1#�>�K��T~޾_�ྶUw��x��w�d�>
��>�l���G�������E���ƽ)�h��>]%�>�[
?Ř ?�>��s>���� ��P�������W������=��������M�@� =d%���(���Q�>��ɽl��>5��>,�>�^>�?�> h��i>K�i>�=�>Bͤ>�ht>�]>���=(%=F�
�W?�؍�ʄ2���ﾒ	�n�e?6�P?h�?!
��E!}��ݾƧ2?`�?{��?���=�Ex��2D���>�g&?�ƌ�Z#?�f�c�o��/S�h� �i�I��.���P�>���xmA��c��#1��V�>y��>d3��9����,S��w~k=%"�?>>(?k�)��AR���o���W�p.S��v�n;g������$�%"p��̏�T%�����>(���-=��*?H�?�������j�g>�Tg>Eq�>��> ��>;:J>��	��a1�ф^���'��0��d��>�{?免>2�I?�<?�xP?EjL?���>g_�>�4��k�>���;W�>b�>��9?��-?u60?�y?nt+? 1c>h������ؾ�
?��?�J?9?�?�����zý�����6g��y��x����=���<��׽K8u�E�T=�T>�W?To
�!9�V���d�>��@?�J�>{9�>�ώ�;g���''=L��>�?@��>���`t����Y�>J�?}6�}\&=�o%>��=����	b����=ʨ1��\�=`<=�����3�=��=-�;�Qc��yټ������<���>��#?�)4>�RV>������|����,>ڂ�>�a�X�F>~�Ѿ�U��#Y����w���`>ڑ�?@�?gIٽ\��>���=4����@u��q��2'*>b	N?���>�NP?�'�?��?i?������n*�������y-?�!,?�>��5�ʾ����3�K�?s\?�<a�"���9)�(�¾c�Խձ>5[/��.~����D��h��m��{��>��?+��?�FA�z�6��v�վ���Y���C?	!�>�U�>��>��)���g��!��4;>��>�R?��>��O?(<{?��[?�WT>��8��.��"ә�؏3��!>N@?���?��?�y?q�>r�>(�)���"T�������Cւ�0�V=-�Y>���>�&�>;�>e��=��ǽ.O��t?��A�=�b>���>���>���>؁w>-\�<��4?+�	?��ݽ��;����Հ���7=rb�?x_�?�7?�E��CCV�+K��ba˾{=(?[Y�?S�?�n�>d*ѽ]P�=�4>a���2_��tB�>m�><�=��>��=��>tS�>�G�>ؑ���$�L� �WBo��	�>��?kp�=�kǿA�q��zp��)��v�<l_����n�7���i\��x�=IF��:��$姾H�\�[���T����؜��T{���>�ɏ=�2�=~`�=�z�<��ڼR��<Χ\=ڍ�<	�=��E�趺<�2��j3��Z��=5����<��N=�l�J���Le?�?��n?�W�>1t���� ޾� 8�0`l���S?�L�>��?�R���X��2��5����sӾ�,�\�,��|�Xj>cpý���=O��<�W�<ň��?�;C�=LF�=�Z��~^�9=��-=%��='�'=�>��>/�z?���������h8����>�H5?
�>�����ξF�U?�7>IS��h�����|�d?�'�?���?~?. ��46�>wnݾ�!]�et�>�Y����>���X<`��=~>&�=�<C�k���#Be=���?H�@]�%?�K���Tؿ��y>�"7>-z>U�R��'1�f�[�W�b��[�u@!?�3;�{˾��>�F�=ii߾�Ǿ��.=T�5><�c=�����[�㙘=��{��>=[[j=^0�>��A>V;�=�5��a�=�UE=�>�=b!P>����@&8�h~*��Q5=,��=��b>�%>)z�>>I�>�y/?49?s��=O5}�3 �?.��۹�>�A>��=����UA=�?�"J?YS?.�+?���>HB����>�3�>L���v��t��.����>�@�?7h�?g�>Q�>'��-0>���'�W!/��M ?�*?镭>��>��� ܿ���$?4��x!�snl�����	ƽ�P�����U����8ѽi/�=�ߖ>]��>���>��o>>6�=���==��>�3!>��A=�4�=��b<�飼�+k�A��=ڧQ=u�3=�r�='թ=*���q�ӽv⟼A�	��9��N�����#��=���>��>%��>��=H���N�.>.Ė���L�'�=�@��)B��0d��H~���.���6���B>�W>?���J-���?&�Y>TV?>���?��t?��>�;�K�վ�=����d���R��?�=g>�=��i;��@`�o�M�v�Ҿ���>V�>���>��l>,�?�Z�w=�	�)a5���>�x��i��r-�T7q�n=��S����i��qغ�D?�D�����=�~?ƭI?�ޏ?�|�>���_�ؾ�,0>hA�� �=�
��6q�zj��Q�?c'?R��>��v�D�dnھ�ҽ{�>;��s�G��B�� ���s1<�ɾ��>M���c?����.��wz������G��4����>�0`?v��?������q��#[�u������J?��n?�Ò>�g?��?K��<s9��0���$�=�;m?c��?�j�?�~�=���=4��t3�>	+	?�?G��?�s?��?��u�>��;�� >�ʘ�;�=��>�=i �=r?�
?��
?�f��@�	����a���^���<<�=�>yo�>��r>%��=��g=$��=%8\>'ݞ>@�>��d>��>OK�>=��'�s��>�<�=끛>P^�>��Y>E��
]ϽS�o��}����R�����b��&��=�{�=�>Z��#�=s�Y�LM�>0ܻ�Ӽ�?��=��J?U:��:�����=K%>���K�>1�G>^��>i(�>т?=���>�X�;/F�f(�=*��W�.�K;.��_i�bȮ����=�;�k��龜�?O�kO������2`��Ҁ�G�t�?>���?�~��7]�`�C�����M:�>�:?��D?�{�u��N��=֣?*�5>��;wG��d ���Ⱦ�e�?�I�?�nC>,�>��S?�g!?������m��Ln�Lk��� ��넿w\���o�n����^��~�_?⚄?�@?�
�J�W>F�^?��&����c%�>��0��#���C���>��<�%�c��7�������n6���4?a�|?ަ6?=>��)u��(>Հ;?�22?�Qs?�0?�:?`;�x$?V�5>��?�y?�5?C�.?78
?�@/>��=l�ջHk#=�䒽U���Rͽ��ʽ����i7=�<�=�K�;��!=��<!𼥗ּ�W;����<��:=a<�=���=쁢>��[?���>�t�>�4?�?&���<������-?�c:
��՜��񛤾92󾂿�=�k?^9�?#�W?U'A>�0@�UB��>��>+�)>eG>y�>����>�r�s<�J>�a>���=�@V��s���;�^g��1�n=,_
>�i�>���>���Y>4`߾�wͽ6R�=�۷�� =��[��E�S��:>�� ��_ؘ>�>?O>?�)>����=�gm�Ur ?o�>��`?�\�?��h�M] ���Y���Y� ��p�>:�>>����^��U簿MC�93>.j�>iE׾����/a>S����޾�n�(�J��v徿�b=����N=�����־-1{�'��=��>d|��z7!�p����ᪿ��J?�1�=[2����b��˾���>t�>��>�	u�b�-`A�Ր���=���>�.=>nԁ�'��^I����$��>ߵK?�KW?�`}?����(/v��K���	�������;G8?J{�>I?�.>��-=�G���(�=md�Y�I�b��>&;�>��r�=�_����,!����>�?�[6>�g?H&R?��?��b?��.?'�?΁�>B��ƌľ�&?2��?���=~�н�W�29�S^E�>{�>��)?)T>�n��>?�"?3!&?ãP?�!? @>`����>��X�>B�>xOV����G]>/�I?��>6�Y? %�?�8>B}6��꡾D@�����=;�">��2?��"?�>?��>��?!+����>/l?ޥ?G�?�
Z?mս`�?>�?�R?O��=���>e8 ?��?8�J?�	z?`�L?�&?�0C<MX�'.�=�w��,)y=��;<� ��o]��!��m)>���>~g><>$�P�0�=ĺ�=Mi���x'=V�<�Q�>�tr>Ɖ��Y�1>�2žZ툾�A>U�e����L��+�:�+��=$n�>�j?��>�"��g�=���>���>���((?�?'#?&;�nb��.۾8L���>D�A?���=�l�����G�u���e=��m?T^?LpX�������b?�^?PX��=���þ��b����t�O?,�
?��G�4�>]�~?��q?̠�>�f�8n�����Hb�#�j��ֶ=,o�>�[�g�d��D�>O�7??D�>��b>�C�=�d۾˼w�Gj���"?\��?��?���?�8*>f�n�c4࿓�������õ]?��>Bɪ��C"?�"���Ͼ�V�����բ⾂����ǫ�����W��u��2�����ս1�=xZ?��r?�sr?��^?� ���c�_�� ��T����Ս��D��bF�F�\0o��������K��]S=[Jf�{K���?O�+?��i�e��>f�s����9���h&^>ik����x�*�=C>D=���=1}�=zL����l找�$?t��>�i�>�;?�eU��q=��98�0�6�����>f�>�9�>�a�>�ћ�r�H���x��������t�lz>�lc?��K?��m?t\��1� ���~9#����h����H>6�>�#�>�zH��4���%�b�<�z�r�~%����x	��=�2?G��>���>�ߗ?�V?p>������:k�AM1�0�}<V�>�b?�q�>���>R����C��u�>��l?7�>��>�Ό�u!�;�z��3Ƚ���>�C�>���>h(o>�*�_[��2���.���`8�+��=:i?�o��wYa��ׄ>��Q?��T;-�m<�T�>~�~���!����W�&��l>�R?%0�=�:>�ƾ���D|����)?CM?�݋�7�&�Z#|>K�"?]��>_N�>G`�?��>�S��I�y���?�;_?iNH?L�@?���>��B=����Fɽ�<&�09=X��>&b><�=���=�f"�4Z`�k���o=�ݾ=	�Ƽ���<�ʼ$�6<]��<�)>H�п�@H�:�侅���ʾG��TO��0&���&�7�)�2Ծ,w׾�M�?�,�C�\��f�����̠��C����?�Y�?�e�u觿,
n�'��`�>^�پM�k��K�z�����"�Ǿ����7@(���D�iȉ���u�JS'?Ñr�Ibȿ���r��Ӕ"?H�+?�X�?g}���%�b�?�p'>�� <���ޅ��j}��F
ҿ�թ��Q?��>�G�}�����>�5^>>92>:z{>�cp��̢�&XU���>Ck?Q�>���~�ʿ����Mr��	�?��@�yA?�(����R�V=���>��	?�?> Y1�U.��Ӱ��C�>6�?���?ZO=<�W�g:	�5xe?Oj<h�F�G�ۻ��=�b�=�=|��J>�>�>؂��MA��Gܽ��4>�ͅ> @#�l���^��_�<�]>�ֽV:��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��=���y�ÿ��9�`�$����=6H�}5Z��\ü�;��f�Z��s���Dw�l�����=*;_>GV�>��>��>0�A?;N?���>{�>w��jV�:|׾ngv��ћ�����r;�!7��Q������M���5�H�-���cط��L1���=f+I�Px���/��
m�.�&��":?5��<�d��#�h�R�E��u��S���_5=�E��9��i]���~��ٟ?ȨU?쎁��Ӆ��&/��-<��kPi?�dƾ����ۉ޾({�>�H��>d��>x�>��ƾ��L���j�	O3?Ln!?n���)����>��(.L=X*?8\?�=��>U?։��Ө���D>@1>��>�D�>GG>$�������?�[O?=	��<���qR�>h�ƾ]큾�	b=]d�=�4=�GGӼN>��;�ĕ���s
���+�d�W?��>�
&����ב��'�+�J=��w?�&	?�u�>��h?>�@?���<���[R����iA�=��Y?��k?	>Q�����ξ���g5?�ve?dO>*�p�wr�)�,�!-��?4}l?��?Dzɼ=\}�󶒿~�
���4?��v?s^�xs�����N�V�e=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?��;<��V��=�;?k\�> �O��>ƾ�z������=�q=�"�>���ev����R,�f�8?ݠ�?���>��������>�d��L1�?�<�?��������,���b��桾E_'���r=��=��1��E	��^�c���kI��K���z
>/~>p�@�.=�<x>��c�g�;|ؿVgw�����H�ѾbI#?��>=����&������4����t�LK�۞��<:�>1�>�W��1A��K�{��x;�/���[�>#�
���>�wT�V��z��Rp:<M�>���>R��>30��A���Ù?���s?ο�Þ�7��g�X?�L�?�q�?97?��@<��v��z����Q-G?'�s?�&Z?s�$�Z]�A�9�"�j?�_��vU`���4�xHE��U>�"3?�B�>U�-��|=�>���>g>�#/�w�Ŀ�ٶ�N���V��?��?�o���>s��?zs+?�i�8���[����*���+��<A?�2>���K�!�B0=�eҒ�¼
?[~0?#{�e.�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?ֵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>dH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?F)�>��?P��=m`�>�N�=[��,�1c#>�G�=º>�d�?;�M?�P�>:��=��8�$/�YVF�yAR���i�C��>*�a? �L?�\b>�긽B�1��!�x�ͽ2a1��輠_@���,�f�߽�$5>j�=>A>��D�7Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*U����*���[����{>��f=��o=cͮ��f\�M'��=M��=$=?>R�M>M�>��>p��>�5b>ZD>$���Eu"��d�����6'���&�A���U:<!.	�9&;ݶ�g�����;S���3�p�-�Cv;q��+��'>	N?J�Z?z�n?���>��ݽ6��<�#�а=��%�v1>��K>�H1?��P?�	?Qӟ�R�w��c��������Վ�$�>��>*�?s�?��?g��=xY�= &@>���>�W�����qS���T���>�	�>�@�>_s�>�:v>�&�>E�ĿyRؿ/$v�X���rR=%t�?�*��p�������z+>����̚>U�{?&�>�c��m�Ϳ¸����6?>��SO�y�?�
�=3FK?z�R?CJ!>�Ƚ,�q��d>3t�_���}��H 9=�҇���N�X��>��?u�f>�,u>�3��j8���P�Vn����|>�96?�鶾�U9��u�>�H�rdݾQ<M>ؾ>+�D�yt�������si�X�{=�|:?s�?]���氾V�u��6���BR>�\>:4=.�=�PM>U�c�`ǽ19H�)�-=��=��^>�?��W>5x>���>#ٝ��IK���>�e>��>?�??s�?
0��@o����^���/��J�>���>���><�c>�5��<�=bB�>/�=>�6ؼ{���и��[,��|>ԝ�����b3b��<ڸ^�&��=��H=���$C����=�~?���%䈿��7e���lD?T+?Q �=�F<��"�D ���H��D�?r�@m�?��	�ܢV�?�?�@�?��2��=}�>׫>�ξ�L�ޱ?��Ž-Ǣ�Ĕ	�()#�iS�?��?��/�Xʋ�6l��6>�^%?�ӾPh�>{x��Z�������u�y�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?toi>�g۾;`Z����>һ@?�R?�>�9�~�'���?�޶?֯�?�6�> G�?�p?�g�>����s�a�)e��h���U���ؽ�8v>��
>s����u�tR��O|��yׅ�$D��'�=D��=���>�ϩ��9Ѿ�X*>fT���������.�\>�Ŋ>�=���>0?H��>��?���>T7��ѝ��YI�'�K?���?���S	n�⇼<x�=�_���?524?U<X�9tϾ��>��\?H��?�[?!=�>����7��a뿿,e����<��K>L:�>�$�>�J��wqK>�Ծ��C�4j�>i�>����~�پ�؁�О����>^u!?2��>ȸ�=�� ?o4#?<Nk>�߳>�&D������E�y<�>�>�>^u?ϟ~?G�?�����-2�"}���}��E�Y��O>��w?ѝ?��>�P��FE��/G��]+[��-����?�jf?V���$?k��?�??�@?�h>I��+Xվ�\��'�>��!?��)�A��L&�@��~?Q?J��>H/����ս|Xּj���~��� ?;(\?XA&?ۛ��*a��¾�=�<�"�S�U��c�;`D��>^�>����ώ�==>fڰ=EQm�I6��f<@k�=l~�>���=�/7�u���=,?MG��׃�@�=�r��wD���>sPL>=����^?�j=�e�{�{��(x��TU�� �?���?Jl�?������h��#=?��??�!�>�G���z޾���Iw��x��y�M�>���>�sl�w徶�������gF��t�Ž�,�[��>;A�>�?Z�>Z�c>��>_ ѾC?"��� ����j��>k:�<�I�`(A�b�"�.�ʾ ����@۽z)��m����_>�5�;�n�>�#!?���>��(>��>�!�=W�>z�>��>:1�>%~>� �>_��>�m>iŪ��KR?L����'���ȱ���-B?�nd?�)�>�>h�������z?���?u�?N"v>Suh�F!+�Lp?*L�>��~e
?B:=�5����<�7�����[��9x����>׽�:��M�^f�De
?S)?����ʡ̾��׽4�����y=�v�?��(?�*�=LR�f�p���W�C�R�����f������$� cq�}������+��˔(���1=/]*?~l�?����X�d��h�k�.�>��c>UW�>�]�>uɾ>&OH>�7	�p�1��?]�Eh'����LK�>�z?��>�S=?�1?�K?@D?��>�*�>�Î���?�='�>Ar�>�d?��=?*&?��>��-?�Ax>v��;X��� ���>��'?=�O?-@,?,� ?���m�_���ǽ9A�=�駾�$|����a0y=#M�͞�<�ٽ\ʼ9[?�p�e�8����K�j>Iz7?��>���>쏾N���$�<���>z�
?A�>����yr�\L��j�>���?3+�sT=��)>��=įֺ��=$������=f%��s6;�#<�4�=�}�=�s���޹��:I�~;�3�<�}�>��?ź�>g�>���Ł �����=8Y>K�S>�n>Ƅپ$s�������g�q!y>�o�?0t�?�,h=���=bq�=SU��it��������I�<Ů?�4#?�BT?���?W�=?��#?��>�!�3L���Q������n�?�x ?�d�>�$���X����0/?D5?;�`��3¾�J��о�=��q���u<����ſ�<�k�W����=����?�2�?�{=.�R���!��"�����?�O�>��D>#�>��;�9���P&��t�>��>��B?��>��_?rA`?��8?����)
]����Z꧿ h�<��B>D�B?DEj?���?��y?N�>{=%l���J�|x@�fB9��늾�Pͽ�C>f>��>[[�>�y�>h�:>�����P=�4�;�=�a�>䚺>��[>[	?P��>P�B=E�I?*��>����N2	�\��A��<�/�@{x?=��?�!,?|`=Mm�Ԋ<�D%����>O��?��?��3?:8��p�=��c��L���U{���>���>��>A>�=�=��=DE�>�:�>��<�
2�&�.�%���
?��E?(s>���������ol��&Al>d
����ȈC>�ļ�+dt�>�����&>��	���N���[ؽG���˽��Q��>#.�=}u�I�Y>�v�=�I����>$>�L�>�W<��X������]�=!y=[�= ˼2r����CZü�-˾Do}?�BI?��+?v�C?��y>�u> 6�7q�>�7_?N�T>1(P��M���]<��ը�TŔ�n�ؾ�W׾��c�d矾��>��G���>g<3>G�=m�<E��=�x=�܎=�r���{=�=�=�Ը=�=C�=��>m�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>Sq7>��>]�R��1�|w\�d�b�
�Z���!??;�'V̾ �>(�=�H߾�ƾ�[.=�6>N�a=PT�?L\�k�=�z���;=(al=�ԉ>.�C>gɺ=����U�=��I=���=��O>�k��x�7���+�"�3=���=��b>�&>O�?U�?��$?ò]?y��>Jg ��D���ޟ��t�>ʢ�>�q?�>���>6�>
��>ch8?��I?���>�eb>]�>3��>���)y���᳔��v2=���?�Ӆ?{#>=I�rm�0��Y�!�}|#=�G?�?�#?�ݡ>��ɼݿ/sU�#8C�ό�}M<}�ݽ�e%��t�8D���%f����Ʈ����G>��>�>%��>�"�>�O9>���>��e>Aff>P<�=�3����;���p�e�"���E=��0>��\<���0����� ����J�����t�=�>=���=���>A>I��>tɖ=_󳾁Y/>ⴖ���L�(��=�D���/B��2d�V?~�j/��V6�ϿB>1X>m��1����?��Y>�?>a��?�Eu??�>�8���վ?O��4)e�CuS��]�=��>�<�q;�jN`���M���Ҿ!��>�}�>���>fW>��*��9�<^=��ξYb8�ٟ�>���Ľ�!c�zo�����p����u���s�O2?`�����0=�[~?"�V?=�?�2�>��ͽ�����3>"�g����=�'��[����q��?�3?��?����@��B̾����޷>�1I���O����� �0�Fa�V˷�!��>�� �о�3��e�������B�{Br����>��O?��?f0b�cW��<TO�����?��yn?Z~g?��>OI?�=?� ���o��p��V��=��n?���?�=�?�>��K>rK'���?�(?���?2݂?�[?m���N�>��a>|v�>˰ľ��=ъ�=f���*j��)?��>��?��ȼ�)꾻��!�2��j���=��>�c>��>;��=��=��>]9>t�L>mD6>y^>���>�R�>�_���h��	?<I(>�5>?0?���>Y.=��]�{�+�`���#%�'�Ƚ��>3P߽*%T=�����=�~�����>H�ÿ�ʌ?Л�>��!��}�>�����o����>��>@D���+?��>�?�>��>��>U��>H��>��>�FӾ�~>����d!�e,C�;�R�ӾѾN}z>���Y
&�Ο��w���CI��n���g�^j�2.��<=��ʽ<H�?������k���)������?\�>�6?)ڌ���G�>b��>pǍ>�J��S���;ȍ�:hᾓ�?��?�;c>��>A�W?2�?_�1��3��uZ�.�u�R(A��e��`��፿𜁿�
�	����_?	�x?yA?rS�<\:z>C��?��%�\ӏ��)�>�/�';�/A<=`+�>�)��F�`�:�Ӿ/�þ�7��HF>��o?1%�?�Y?�SV�7޿�<?#>�a<?O1?��j?p1?��=?���҇(?�ZF>��?(V�><6?�[-?^�?�N >��!>���<�|�=�L	��b뽽i����E;�Z=��=��N�L=��~��TD=��=�=�?=c�<�bW=� �=劳=��=���>à`?q?�3�>��?0v&��A���w�MIJ?й=�Wu�:��7��(ݾu�=��b?F��?p?���>f/B���E�E%>��>�lE>Ա�>���>4�>��*���Q=���<k��=2H_=w %=�g��}������׽��B>���>� y>�̊���)>[6����x�5f>�;R��<��ER�ԻG���0�s v���>�K?t5?���=!�辧�����e�N�(?ȟ<?�:M?\?�c�=Փܾ��9�/fJ�D�rs�>0N�<ڃ	�fݢ�����ޓ:�Kǖ:�p>�����!����a>��g�޾�wn��(J����eMN=�d�T+T=P�w�վ������=:>
>�~��e� ��!��"ͪ��4J?�m=|m��N�U��˺�&�>a��>>��>�w9�D[v�x�@�����az�=���>6w;>�Y��ﾴ�G�h|��2�>�ZD?��e?1;�?M��Ef���B����{w��!�Ҽ�Q?���>C?ƾ$>zv�=�.����Ƞ^�[E����>�+�>_���1J��1��)4��PP���>��?�M>л?�E?���>6]?�(?-�?�s�>|��������&?f��?]��=�Zν��W�g8�?+D��.�>�)?�?��R�>Q?�I?�o%?ANP?�s?W>>$���2>��(�>���>}�V�O߯��1V>�>I?�t�>s.Y?�Ń?t�;>e�3��9�����0b�=b+&>�u2?�!?>q?d��>{��>��վzr�98�>s�?I�?�l?�^+��>��>�?�W�==`
?x6?.l�>�2?�uc?ZU?�1?��=��<��x="輻��:\=�	�"-�����]� =�� ����<����<n�U�<�=�h$<i-=��L=���>��m>룂�%{<>�����"~���<>�͞<������}���1�ƛ�=�)�>�h ?>ߙ>Ë-�oѱ=�]�>"�>4��k$?'X?�V?0�[<�L\�]|�L�q��b�>��C?�[�=F�e�xۑ���q���r=F�n?��[?�B�
2����b?��]?sf��=�[�þ�b����?�O?��
?��G�-�>��~?��q?`��>g�e�:n�����Cb���j�g˶=Sq�>�W���d��?�>��7?�M�>��b>�#�=�v۾��w�r���?��?G�?#��?,*>Z�n��4�������ĭl?�i�>-�Ͼ�m6?��+<qpӾD�i�������)�0�̾T ���.��l�:�����V�-��<>�?�*v?܀?;CS?�H���?�V�\��Yc�3�,��!��'���W� ��j�<�e�n��;J�u������4	>��-��6���?^�)?_^���?�a����pϾ[lw>�N���Ľ��=	����ڮ=�t�=U��s�3���-?V�>xM�>d6?��9��%<�M�&��i*�c��}�`>���>v]�>�@�>ךz=T��?��;����t���&�7e>��f?��E?��X?+�G��:c�bj��^�N���'����xv>��T>���>ڟ`�n����z]��$e�㯀�Q\�n�����"��o.>>? o�>��?3�?��>�) �����	�#�.��=[��>ʽn?��?��>�p.��&'�G�>�gm?K��>��>����zR#��|�y@ս�y�>5A�>���>�r>��*�<F\�CS���	���):�QW�=RYg?�׃�
�a���>C�R?9{�;"P<%3�>�%u��"�z�����*�Gk>6?�;�=W�<>O��I���{�K���)?�		?Fф�!��hc~>�?:��>��>�ۆ?���>P��Y���"�?O�X?O�S?��<?��>���=�{��ە���X��
!=�ʐ>��v>\H=�6�=
g��E���6��i�=rQd=L3�<�����4t��D��;�W=�Z>Өۿ'PL�~پo�����Uʊ�<�����B �Rn���p��u�	r�PT>��QT�QCg�׋���h��5�?+��?����c���n��鑀��x�����>�"n�^M��Y8������ �����{��i���N�i�])e�۔'?�����ǿ�����;ܾ�  ?�B ?e�y?v���"�q�8�� >r0�<'.�����w���(�ο������^?~��>~�'��.��>ҥ�>��X>�Hq>��Ꞿ�!�<X�?*�-?j��>��r� �ɿ�������<���? �@��S?Z��,��>�s?ʨ?Yр>��=��2C��>1��{�>�Ʃ?�R~?�:>�;�5�=Nj?ʳ�;�83��
�=}>�=���]}@=u1�*4�=�>���@����ϼ4
>L�>����5ډ�K���h(��Ȓ#>�~���%�2Մ?{\�if�v�/��T��	U>��T?/+�>+;�=��,?.7H�b}Ͽٯ\��*a?�0�?��?�(?�ڿ��ؚ>\�ܾ`�M?_D6?���>�d&��t�/��=�0Ἦ���h���&V�k��=f��>S�>O�,���W�O��H�����=;�
�K�׿��=z5�c¼Xo���d���f���7��Dk:��ݾ�>ؾ����=t��<\�>j�=<S��=:��>�L?�}C?���>>��=$\�;��Ǿpp��O_�9�4S���D��K����+>�8V�6o��&���"��i� �Z@����o�����bX�����\��y��u�%�#?uIo>Ф	��Ζ���I>ca�������~)=D���X���1�����?M:z?!�z�D%�|~�=z�(�}OA?��+;J�������==�O>�m=ڝ?t� >J"ľKu+��=��@=4?�}?�t��(���]4>�_��xJ=W�*?m��>mS/=���>e�$?���IL��"�e>�C7>��>��>��>}��.kսV�?P?��Y��c<�>����Z����=p�=��0�����V>2�!<f��l"t��'��;P?5s>/�ي
�V���;��>��k?���>�Ǘ>">r?9�6?��<0�߾&�H����i��=ii?ɰa?���=|��Bg��h���P?�Dr?ͰU>��0�v辮�6���7�?�b?\� ?9��<�jo�ۀ�����פ&?/�v?/r^�`s�����&�V��<�>�]�>���>g�9�Pj�>��>?�#�G��+���Y4�?.�@���?�<<'�ښ�=�9?u\�>��O��=ƾXt��O���`�q=v"�>J����cv����jP,���8?���?6��>�������=P��,��?�z?֗�&#�=m����h�����9�	�	�����+�������Z��Z���;����>"Iw>��@��,��0>��U������jȿ;=y�L;��y�;H?�^e=�<�������@ꋿ�Mo�w_^�5�,��A�>|$!>��S� ����|�4�5�L�T� <�>Ƃ�;���>�E)�⊹�h`���sκ�ɓ>r��>�n�>�&^�7���|b�?����y]˿~A��dP�K?*l�?�3�?~z?���<L�e�:)v��hr<��E?-}p?�R]?C���x���XW�%�j?�_��xU`��4�tHE��U>�"3?�B�>T�-�e�|=�>���>g>�#/�x�Ŀ�ٶ�=���Z��?��?�o���>q��?ts+?�i�8���[����*���+��<A?�2>���H�!�B0=�TҒ���
?U~0?{�f.��^?cQ���e�I4'��s��$}�>SV9�C�O���%=��۽~Z�)�w�U����?I�?M�?,�id�p�#?�w�>䵰��|޾���=�T�>�>�Q>K)��#k>�?�E/.�6�U=}��?w��?-?P�����P	>��q?;_�>�`�?���=�9�>u�=q���6�8�?�!>�=ˢ �g�?��O?���>���=�2�S-���C��Q�rK	���C���>�<`?��J?Дc>+�����?�:z"��ﹽ��*�� ���F�i=�$�� 2>/7=>Z>c�B�Dv׾��?3p��ؿ�i���p'�}54?���>��?���t�j��u;_?�y�>�6��+���%��uA�i��?�G�?O�?Q�׾�e̼�>��>aI�>��Խ����c�����7>�B?:�RD��3�o�t�>���?�@�ծ?Zi���?��T���}���Ǎ5����=)7?n�𾒊y>���>�ܨ=�jv��_��K{s�/Ҷ>b�?�?�?
��>�l?@o���C��4=pݢ>
�j?��? �U�@>iJ?���x�������e?H�
@'G@�_?�����ֿy���~��y���`35=S�=,�D>6R.��=���<@�Ӽ#�ǽy���D�>�R>�[|>��W>ճI>�!>]Q��j�'�0ߴ�ge��c�V��z%��A��3���%���a��r�O���8[�i��<T������}Y��-O�Od���0�>�N?��7?'sk?��>꽫9B>���\E���,=cҷ=iX�>��J?�)U?�X?��=�x���P��u�����ŋ��!��>�.>&ڱ>�$�>T�>����hV�>��=�ul>V��may=����Q�̆>���>ȅ�>
��>G�[<)n�>X�ڿF��޻j�,�w� >����?Dy�=>\K�̳���*>�s�P����^?�>+���Y|ǿk�ֿ[�+?����F���1>�I���?1F�?r�>̉���,���=��9�ǆ��	7U>w��1���Ų�za>�'?��]>i�q>��3�ą7���O�ci�� z>��4?�ƹ���H��]u�_�I��I�|�?>#��>FC���w�DҖ���}�{ck�{�V=QW8??��������7��U̠��yX>Md>#V=r�=3zN>'l@�T�ν��A�RNi=�y�=�Ma>.u4?�1�=��>>�I�>k��������>!��>����L6?�
?��`=��L>�VV=�; U,>���>�ɿ>P��=�V��=��>�=>�ý ��<EH���Ƚ4<=�y��s�\��]M=f/ >����0�=iM^�E�.�C�������~?Y���㈿���]���lD?�*?B�=[�F<�"�����wJ���?;�@+m�?X�	�>�V�~�?�@�?�����=�}�>�׫>�ξk�L���?0�Ž�ɢ�Q�	��'#�
S�?��?"�/��ʋ�3l��8>�^%?��Ӿh�>�x�jZ��W����u��#=ĩ�>}8H?�V����O�7>��v
?s?�^򾯩��F�ȿ~{v����>4�?���?�m��A��n@����>Т�?�gY?pi>�g۾�_Z�d��>��@?�R?��>p9�]�'���?߶?���?���=�`�?"Qj?�T�>�{�����}����ґ��=�Ž���>�">��ھ/���/Ӽ�����A4��A��h��>��_=���>�a�aX���6 >�ޙ�=a��*�����>G.)>��s>[@�>\�=?��?^�?�=����1����M? �?t��U�i�n��<3�={�R�I#?�/?	+y�[�;�>//]?�#�?~(Z?��>�w�a��b��ǘ��ٕ�<HL>��>��>s#��&�A>%پ��9�)��>���>Cv�^�׾
���Y�Ố(�>C�!?���>�T�=� ?Μ#?7�j>�'�>=aE��9����E�ϯ�>���>RH?��~?��?1չ�[3�����桿
�[�o;N>��x?�U?�ɕ>m���e���i�E��KI�� ��?�sg?�S彼?�1�?��??(�A?�-f>���ؾģ��6�>;�!?/��ˢA�&�����n?�Y?���>)����2ս��Լ����#��?6!\?2&?����a�D�¾Z�<�"���U����;bsC�*�>��>u~���մ=��>�K�=��m���5���d<�U�=�D�>��=�F7������v"?��"=��O�!��<�O���IH�],f>Cwh>1b��G�\?�)�x��۔����X����?j��?f��?1{��?Y��^7?�{?��?�H?��ğ������X��#ͷ��-��.�=���>�N�/�德������.)���ĽZo���>�/�>��>��>h�3>1�O>�'����"�O��Y���!p��<���=���-����f��tK�qS������s���3PV>��=,ǟ>�-�>�Ƽ���=(�?�H>���>�->���>F��>6>n�[>��>��a>�V<eiR?����w'��C����nB?�se?`��>Ý��x������ql ?���?G�?~zu>�|f���(��v??��>����"�?�FB=����6�<�ڱ�4�|���L4���>����}9�n�I���b��M
? �?i�|�m�Ͼ�轜ǣ�x�>t�?i"?�q5��[��Xs��U^��KD��ý��C�V���f5�/�����*���@∿��*���>)�?��?��	r��묾�߉�Ja9�:NJ>���>+ï>���>�:>>~վ��C�/Ro��:%�~��v%�>²z?�r�>�vK?e�7?��M?�F&?c�P>'�>�=N�N��>q�y<�*�>�>ЎI?e%5?b�?�=	?QV*?\g>�)�9���+��?��>��>���>�| ?�x�>���>f;9�}�;p���b�.fZ=�"�=�D>�,sA���>�U>��?F����:�6����;V>�K3?�~�>T��>$F��$mu�{@_=�&�>�?�>mL���Ym������>��? ��{r�<��%>��=�w�;駓<]��=�d�n�=�93��@6�0�<}��==��=��d���<���
�j�D�[<���>�w?�ޅ>��>w���/��1�
�bH�=e.T> �M>bu">
�پ�ۉ��'��U�f��y>TQ�?��?2�}=i!�=��=���5����DH����=��?��!?��S?䇑?i=?��$?/�>C�ɶ��7������#?���>���>ޡ���l��"�#���C?��?f�U�����j���̾Բ����>�/����v�5:¿ �m��d*��Q)��@*�h��?	ͮ??U>f��j�9������>�N ?F�j=�ټ>��c���J�0��P�>0��>mij?R�>�O?I�z?:�[?0�U>��7�]i��3Z���b��#>�??-Q�?�ǎ?�x?��>�>]�%�� ߾(b��x�#����?9��:&T=k�W>w�>��>qn�>n�=Jf˽x髽�_@���=�2b>�e�>E�>���>f]x>���<d�=?�P�>�Ò�����Cg���t��ٯ��j?�?z;?�#	>��/�%t���ƾ�+�>D2�?�W�?�7?����>�9��Q��f<�ֶ�>Ą>Eɟ>��v>kl��}>�a�>{n�>��-�U��i�1�pʽG�?@�A?v��<
�ɿ�]|�<-|�樨��<�<Op������-}�0O��x�<�:��Y���y̾��l��o������&Ⱦʵ���H�}"?��=�z�=2�=�3�=�1�����;���=##W= Ȁ��m���;�=��ռ�I<��U��<!�<�H�<���<V�;*���6v?�VW?߳,?�U=?/8�>a��=����6�i>�'ٽ�?�\V>����<ɾz�G�4kž��N
ϾϷ۾�MQ�����>����d��=X�I>A�=L�<��=�� >b��=�n�3ɼ���=n`�=O�=B�>'+5>�# >�6w?���ֲ���4Q�RZ�v�:?8�>{�=��ƾw@?p�>>�2������nb�.?d��?�T�?H�?�si��d�>���v掽
r�=����>2>���=&�2�g��>��J>���K��g���m4�?��@C�??�ዿ��Ͽ#a/>��'>� �=��V�7�%���w��kZ�Y,=��?�0��
̾�>��=�ھy�����;m�%>���=ԁ���J���=ZX��%�C<�z�=��>�9>[f�=c?����=b��=��>��r>3<�=j�3�m,K���<n`�=t��>��>U�>EU3?��@?y:4?�#=>!��]���7�����>��$>w��>+(��
> n1>@�?2p4?�UM?.��>�H>É�>D�S>��$���}��n��eؾ0C=G��?w��?���>'w�=�HֽsZ�D��^Q>��[?_cS??�/?l��>WQ���7D*��3�B擽�Jr<��"<L�H��?o���!�e%-��M����;)��>�#�>Y�>78V>9?,>D�a>�־>�>��=��m=�P�<�=���^�=�Y����=�$W��1*�7r'�����&a������e���U =2/�=���=�}�>'$>U�>��;����7�>�Ds�f<6�/@�=I�����G�^ ]��w�3���C��56>x�h>����ي�a& ?z2W>(a>��?��k?�A�=��ڽ�kھ������p���M�G�=#��=YqS�ٰG��rs���X���۾��>c"�>�͒>VM>y*�rg8�`�=��վ�N@�	Z�>5p�����;�'%~��硿W"��em�M]��:�7?lǈ���O=�t?YOQ?��?K��>e:�����>��n��g>V���o�oإ�<�
?qK(?��?%L˾��7��̾����}�>�vC��J� ���X~*���Ѽ�ѹ�:��>�5��M�ؾ�J5�gZ�����t<�]�a�P��>s�J?�{�?�/l�J���:�D�U��-7�����>*�`?�>�>@�?s�?�a̽[E�+Y�H��=�*n?�W�?�_�?TR>C��=a
�)��>��?z"z?@�?�*d?�]��.�>���=�>��/�=9�=��;m>۱?�y?��?L�%��B ��Q�;F]��8��=�b>2W�>���=��F>�� >1P�<��)=�(f>��>d�>�J�>Ì�>R?�>E:žݖ'�Z/�>��>�^>�t?��=�e����F��D�<CRO=�� ��y���F�T�x1�=a	=N��=K��=0�>ccĿ��?±�>D�����'?&�<f��\��=,�>�s��u�,?��>���>.8�>�M�>�>�[�>�\}>5LӾ�l>���`!��)C�%R��ѾRnz>Ꮬ��&�������RLI��l��'j��j��+��G7=���<�D�?�����k���)������?$Q�>�6?�Ō��Ո���>"��>�ٍ>`0��ύ��č�q\��?M��?�a>z�>n�W?��?1
4��73��_Y��u�޹?��c�F�^�砍��Y����
��9����^?��x?T�@?^d�<B�z>��?�&�����I�>��/�Q%9�k�S=�>�Y��Y3`���Ӿ�(þGI���I>k�p?VE�?��?��S�ЀQ>�>�G?�9-?�`?G�'?�@?1��B�>��Y> � ?���>��J?��,?�"?��=�/8>#�<��!㽈��S.���0��JW<��=���=)�P��4>H�W>/�'�����!_��}�e㼗P1�������3��=:_�>[�^?�?s_>� ?��4���+�s����@?x��=?�vƍ��逾�뾮�R>.�q?�W�?��Z?y�l>��-�8�p��)G=��S>�0>�N>zE�>������*�=/�=��+=���=��޼�����l���B�=�>���>2�>ӗ{�2>ɩ��&��K�Z>�MB�_+���`R��E��)4�\[u�� �>��K??f?�ϗ=�>��3����b�#(?�:?�M?�?��=\�߾�5��K���=�{ۛ>J�<�a
�����8����w>�gM꼧�]>�k��Ҽ��cdQ>`��=>ྕ�g�cL�bS㾷\=`�-u=Q��y�ƾ,���Hh�=��>�ۺ��\�F��Wި��I?��=?���@\��Ķ�T�>Z��>�/�>���fV��arA�R���+�=�I�>�o@>*���C"��s�H�ٮ	�-~�>�"E?W)_?Jq�?�Â�M�r��B������l��`[ļ��?��>g�?�|A><)�=�L��i����d��G�S�>z��>ƪ�E�G��󟾥�����$�Oъ>/]?��>1�?�OR?��
?�`?�A*?Ar?h�>4+��Ps���&?hS�?w�=��ͽ��Y�`�9�PF�cg�>�'+?�;�}��>��?�?��&?�(R?�z?Ӑ>0���@���>8w�>ғV�����[^>�>I?�&�>��X?Jۃ?�=>�u4�uܠ�\ ��Q+�=!| >�2?a#?>�?���>���>������~=n7�>JӇ?���?r�c?��m;�4�>[m>7�?� j=��?d\�>�
?�f?�?�}f?3.?�L�<3���X��
mM��N��=u�>gc>�d%>���=hǽ�L��Z:O=X�мQ��;��,=j��<�=��>m�>}�z>�핾��%>��ƾ���ЯE>�Zl������1���x5�Ј�=��t>���>���>��1�=��=E��>���>�
�%?�?(�?,�vrb��,Ӿ��T����>#=?m��=��p��򓿳Su�K��=sn?�b?��Z�(���I�b?�]?h��=���þ��b�ŉ�E�O?5�
?(�G���>��~?Y�q?'��>a�e�&:n�#��Db���j�%Ѷ=Sr�>EX�=�d��?�>]�7?�N�>8�b>Y%�=�u۾%�w��q��e?{�?�?���?�**>q�n�U4��׾�I��w�q?�o�>d�۾R�.?2�=:cƾI����:��[ؾ�ʹ������k��a����ǽs5l�n�w�)�9>�O?-�?T�z?�M?���(\���R���X��;k��,&�8�2/V��Q���;��Ĉ�zL:���j=���6>���'�L�g��?�&?/K����>�+��JK����˾p�a>P�����4P�=���H�=0v�=bV����v��'s?�	�>n��>a0:?@X��W7�ę&���,����>���>�ˈ>���>D�<=�lZ�W*��۾ρ��d�v��F�>�Ak?��L?��j?)ٯ��
:�mO��&P4�ɞ<����>$>��e=��X>�v9�KB3����~>�lb��(�Ժ�������=�7?��F>0�>g��?tw�>?-������U�1�>�(��A0<��>�u?���>�֟>]���Y�����>��l?99�>n(�>�e���!!��y���Ƚm�>��>m9�>3:m>�f/�M ]�`*���h���g8���=��g?�܄�-�`����>�R?"�:��<�#�>�B}���� ���V-�a�=X�?���=.H?>��¾�4	��,z�����s�)?��?Q���&�=�h>/?r��>T:�>�ʆ?���>}ȹ���Z;��?�E^?��L?��D?��>Mr[=�-����̽�N"���H=���>� a>=}=1��=�f"��`�����;N=���=T`¼�½���;j���_=<���<b5->ۿ4fK�%oԾ�z�X9ﾁ��ke��տ���쇾v
�jش�����q\��<��a2�LV���f������e���?��?P��{���f���l~������h�>Po�#u�������ʑ���۾�����!�t)N�(2j���g��.?��ٽ�Կ#Ͳ�D�m�{&I?�tR?la�?W*+��B;�U�Z���>'� �^�=��&���"�ӿ�z7�f%?g�>F�Ͼ��>���>2� >θ= ^�<�4�㤞��]��r7?P�*?�?�Ce������E¿�r=���?l%@G2E?BE/�K־�s�>֙?o\?�>�#���!��dP��6�>,�?3��?�}
��Q��3�f�Z?j%�5/�{�R=�?(>�8Y�i����H��=�0>�������tN��*�=Z�7>�	>.��1��A�3>�W�>���xw�4Մ?{\�nf�y�/��T���T>��T?+�>?;�=��,?A7H�\}Ͽ��\��*a?�0�?���?2�(?ۿ��ؚ>��ܾ��M?`D6?���>�d&�!�t���=4�^|��n���&V����=1��>|�>��,�Ջ�k�O��G�����=�:������R�����'��=W��l�q��fX��?�M����7��p4��n���+yi>�>5�=>) N>G��>I)�>J?� K?�>��/>�X�D���p��~}C��Db�zЦ�j�p���n=����&�����r�r�@�ԁ@������.�7�=��U�w'�����՟l�����7?Y�L>$p���:W�tÂ>�*��zu����=6���j־3G����Ε�?��>?�C|�F	V�%���gޞ=�7�$p?���?�}
�̐>� >E:
���>� <� %�K�L�@]_�])?9�?p���?����>�g	����=�)?���>�Ơ>=l?�{E��d,�IEC>��>�>��>�>�c��A��U?˯X?�a��/렾�n�>є��͟D����Sq�=Ht�6�T���E>��*=4���:i=S�{�i���x(W?��>h�)�o��`����JZ==:�x?��?!.�>c{k?��B?�֤<�h��U�S���<cw=��W?*i?ں>T����	о����\�5?֣e?f�N>�bh�6����.�-U��$?=�n?�^?(����v}�D�����n6?��v?s^�xs�����I�V�g=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?a�;<��[��=�;?i\�>�O��>ƾ�z������E�q=�"�>���ev����R,�f�8?ݠ�?���>��������>��p�͆�?$<~?����"Yb=�7߾lX�J "�S�Ǽ-�>�SJ�LbU�C(��=�g�S���g�����`>��>@��1����>����ۿ�ӿ�Z���R��8���g�(?��>*"��0y���턿����:\P��=o��d^��E�>�>��������A�{�q;�\����>w���><�S����o����6<��>F��>���>'3���꽾�??U���<ο^���ĝ���X?�e�?hn�?(r?]:<��v�az{�a��&G?��s?TZ?�M%��7]���7�}�[?�R���W��C���3�an>G�)?���>��>�>ż�|>�?���= ,+�-������a�	�?��?K� �ߓ�>�?��S?�v(��c���񣾒GV����=�,3??��>
�o/+���C�D���?��G?/H�#��\�_?,�a�L�p���-���ƽ�ۡ>��0�f\�N�����Xe����@y����?M^�?i�?ӵ�� #�g6%?�>e����8Ǿ��<���>�(�>*N>\H_���u>����:�i	>���?�~�?Oj?���� ����U>
�}?;"�>T�?
x�=�N�>�;�=����K-�iO#>��=_?�ݚ?E�M?3�>��=�)9�#/�0XF��@R�����C��>��a?��L?�Fb>4B��P�1�M!�\�̽�1��,�ߑ@���,��߽�U5>
>>RG>Y�D�FӾ��?Gp�6�ؿ�i��)p'��54?1��>�?����t�����;_?Hz�>�6��+���%���B�^��?�G�?8�?��׾HR̼>2�>�I�>'�Խ����M�����7>+�B?z��D��u�o�|�>���?
�@�ծ?ji��	?���P��Sa~����7����=��7?�0�	�z>���>��=�nv�߻��V�s����>�B�?�{�?��>�l?��o�K�B���1=2M�>Ɯk?�s?�So�~�J�B>��?)������L��f?	�
@u@\�^?*���l�������G�� ��>6�=%�Y=���+>s�t=S�u=�Ci��j>��>l΅>y��>�j>��g>�<!>? ��YU�Ҫ��"i��	���L���,��%��,!�G_�!-߾^о����hI�~'���Żiw)�I�5���ǽ�<!>+�K?�CS?�u?>��>Բ5�q�%=��F�.=��*�LI>I>��?�1U?Y<"?^�O=S/�� �l�t<r�^��\�Ѿ]<�>w��>�;�>�{?�I�>��=i�j=Ԇ>'ѷ>��z>yV�<Hb�w֊<��>���>	>�>��>�vx>h��>��ÿQ���� � X�%��=�?���0�^����i��;�ܾ�.�=�<?�$e=�o��qϿޓ��$^G?X9�g�5��(־���>�a?��|?2�k>����t��fgB=V@�����<>P��u���=�{��>�J?��f>4"u>�3�Ea8���P��|����|>�/6?�ڶ�3e9���u���H�bݾ�
M>V��>�,F��b�3���zui��T{= r:?t�?�(���ݰ�o�u��>���dR>w\>�=�=;zM>�Xc�E�ƽ��G�S�.=���=��^>��?a4>㇛=��>oc���^����>�lE>�K>#Z@?CQ%?�'��:q�[҂����u�>�X�>ѩ�>�$�=�L��!�=;t�>n^a>/ל��b��&�W�I�c8N>�Oq�<�Y�������=~��a��="�=Tl�m:���=�~?���$䈿��8e���lD?V+?P �=t�F<��"�D ���H��E�?q�@m�?��	�ݢV�B�?�@�?��_��=}�>׫>�ξ�L��?��ŽBǢ�͔	�#)#�eS�?��?��/�\ʋ�Al�p6>�^%?�ӾPh�>}x��Z�������u���#=Q��>�8H?�V����O�_>��v
?�?�^�ߩ����ȿ3|v����>W�?���?i�m��A���@����>;��?�gY?qoi>�g۾6`Z����>ӻ@?�R?�>�9�~�'���?�޶?֯�?U;�>ő�?��n?�3�>���G��Ǧ��쒿ثC=5�c�8��>q�s<sYQ��M���|��'Z�!D�rˑ>�_=z��>��@��bm�6�>�M*��c���R��|�>��
=�
���7}>���>W|�>�M�>�^>ZP��5tx����q�K?���?���~2n�@N�<���=�^�Z&?vI4?Wo[�%�Ͼը>��\?u?�[?�c�>&��Q>��/迿~�����<G�K>W4�>bH�>P"��gGK>]�Ծb5D��p�>fЗ>�����?ھ�,��O>��.B�>�e!?���>Ӯ=�� ?4�#?˭j>Q*�>VdE��7����E����>g��>�E?�~?��?WԹ��]3����硿�[��#N>��x?T?�Օ>����������D���I��7�����?:vg?�;�?�1�?��??n�A?� f>��� ؾS⭽��>��!?���A��L&�2�(|?Q?���>4.���ս;Nּ���;z����?�%\?L>&?{��J)a�>�¾�,�<'#��RU����;1iD���>Ԋ>+������=�>�ݰ=�Lm�};6���f<�v�=��>��=
07�
y���I,?l��y�{'�=�~r���D���>��H>�h���?b?`�1�G{����J��%�D�,��?��?��?��Ƚ�`g��]:?鶇?��?�L�>�ʧ��ݾ�㾊ǂ�O���Z��A��=oӿ>m�&V�Z�����%��@�ʽ����V�>2˘>�8�>m��>���=�� ?��G�Lx���(��n@l����T�V� �~-���B������1�xC���ߚ��&�>r<�=�k�>�k�>�"�=��5>��>��c��ʔ>�ә=��
?�>Yj`>o!�>��Y>͞ۼ7;��KR?�����'�M�辊���c3B?�qd?31�>�i�*��������?���?5s�?�<v>�~h��,+�wn?~>�>=��Zq
?�U:=;��3�<NV��н�3���M��>�D׽� :�}M��mf�xj
?�/?�����̾h<׽������=M9�?R;(?Z�-�feO���n�/�X�FER�����T�\,��sE#���r��ғ��$���s����)��̌=�h(?2�?�������Ўm�'SD�?>�L�>��>�q�>u-W>�
�m�0�CC[��u&��φ��>��s?{�>?I?��<?�N?�zB?`~�>"F�>����o?p�T=��>��>��9?�)?��3?�s?�0?aCq>y��B����d־��?5�?�0!?��?&��>U���v��F��ls��-y���~�f=7�;��b�����=H`H>/-?S���8�`����;j>w?7?���>P��>���gف���<*L�>�
?Hn�>�����r��'��q�>��?U���=}*>�J�=>Ӄ�[W��ʡ�=f�¼*�=檆���:��<���=��=��h�bF9^;���;�w�<�t�>3�?���>�C�>�@��,� �R��f�=�Y> S>k>�Eپ�}���$��q�g��]y>�w�?�z�?»f=��=���=�|��rU�����:������<�?8J#?XT?\��?r�=?nj#?Ե>	+�bM���^�������?��,?
��>�2�5���c��1`���?P[?�~g�+C���(�!ڂ�ׯ���Z�=v^,�FP��/���1'�V�>=��u���S�?�e�?=�ٽ+�>����d��� ܢ���>?n��>H4�>�{�>kO,���x�x���[>u`�>%�^?�u�>��O?�{?x�[?W}S>[#8�(���ҙ����:$>P�??�w�?�?�?�,y?��>�>W*�o=�O�����;���i��Z�h=s�X>�9�>�"�>�]�>M6�=ܬ��Y����x<�V�=��c>�\�>
�>j-�>�sx>g�<ޓK?���>�ԅ�l�;s�ﾼԾ�I��Ιj?{ �?��L?�9>3���h�;í�z�?u�?o��?�7?hn��B�=Z��;Pa��,i��'��>�'�>�o�>�/	=YӦ=��>��>���>�������������?]�<?���=G[��*�]�)Q��&��c�<"ؾ\9˾�6��������=W}���������>���t���̹��r����X�܇?;��=!
��&����<=��7�F�G>;�`>� =�R�=�lֽ#L>/��i3��P%��$%=a4�=H���G�{�˾I�}?D;I?C�+?�C?>�y>�.>��3�[��>O����>?IV>f�P�y���S�;�����z"�� �ؾ�w׾v�c�_˟�;J>�4I�[�>b=3>�4�=5�<y�=)s=ν�=g�R�a=B;�=�k�=Yv�=���=��>pO>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>ĵ.>���=u8R��<1�Z�Y�WDi��W�sY ?0�9�axȾP1�>�I�=���<(þ�('=�3>�Co=��pWZ�¤�=!�u�=��h=�؉>}>>�9�=������=�E=�5�=\�Y>�b���PO��1��(I=�ۼ=�Z>J�>&;
?�g?�~?ڗj?M�9>Ip�����M㤾�ٿ>���> �>���r��>�Ρ>�b8?�WW?̸]?4!�>��3u�>���>?��t�n�>:�L(������?���?B��> ���Z��Á(�=\����>��?��7?x#? w�>���W翐�(�<Q*���,=`�]=�?����AH��h�~�B�ٽg�/���g=�b�>g�>�'�> ��>��:>�f?>|Z�>���=�3S�i��=){��x�5=5�<n�=����Br0�;˛�h��<e��Q���9���C=cKQ=XD*<�cX=r��=���>�->���>�;�=���Ot/>�����L��X�=bG��k-B��/d�tP~�� /��w6���B>�KX>�s��/��b�?`�Y>��?>�}�?�2u?��>n(���վ�R��]e���S�K+�=��>.�<��o;�6@`�(�M���Ҿ���>Y��>Y�>^E>`?,��8���=sIϾ�2�̀�>V��l�� |,��w����&���We�Id<S�D?�$����=�Wy?[OT?^х?��>���U�K�l>y卾%�4;�$����^hսd�?,S*?�?H��b�G�|H̾����ݷ>AI�c�O�<�ί0�r���̷�K��>������о�$3�'g��������B�QKr�w�>��O?�?W:b��W��TO����Y)��=r?|g?X�>pJ?�??�!��^y�t���x�=��n?���?�<�?�>Z�>/�����>L?���?U��?+�c?Եm��!�>$
�<#�b>S��.R>%Ғ=�M=o��=V�?܃?ͦ?N�$�+d�v}�����6�?��=W��=��>��v> U�>��=&�=�$>��>:�>"�>`ƃ>*��>�K�>*���#�U3?3(Y>�[�=��0?bؚ>�8+��p�:<�=/�L=�T<���.>�y[��n���	>���=�b�='�6=�G�>�Z��>�?���>ۢݾ�'#?r'���G��ov���?�v �q�?�҄=z��>C��>�0�>�=^0�>�Y�>y-Ӿ>g>����G!��C��oR�!�Ѿ�Cz>������%�n���<��hFI�Js���_��j��%���>=���<KC�?�^���k���)��!��a�?te�>�6?�댾T�����>��>,ɍ>9y��B������S�t�?���?u;c>��>��W?Ӛ?��1�c3�wuZ�îu�(A�'e� �`�o፿���F�
�%����_?��x?yA?�T�<o9z>"��?��%�{ҏ��)�>�/��&;��><=�+�>�*���`�K�Ӿ�þ8�~IF>`�o?W%�?\Y?<UV��k�8�&>�z:?��1?o�t?�2?�D;?���D^$?A2>��?'x?�5?7G/?�
?b�2>�y�=o�s���+=>�4���q�ӽ�νs��@7=�(|=U��:��<�C!=�/�<l]���bؼ�5�:�J�����<�H>=���=���=��>�qZ?�t ?�_�>��?`���#�����VU?�6q>t��!Ć���V��SϾB�>��?i��?w�_?v^>+aR�ZP1���T>�"�>1�>��>s�>�.O�TÎ��*�<���=�ȫ=mU�=���	�����	�������=q��>�={>�ǀ���/>�����v�Xb>�WU��o��]^N��}D�E�0���u����>�vK?�8?��=��.���Bd�.%?;�9?'�N?|��?~t�=��׾7x8��IK����{X�>���<*�U���u����x:�|��:$�t>6������/a>S����޾�n�(�J��v徿�b=����N=�����־-1{�'��=��>d|��z7!�p����ᪿ��J?�1�=[2����b��˾���>t�>��>�	u�b�-`A�Ր���=���>�.=>nԁ�'��^I����$��>ߵK?�KW?�`}?����(/v��K���	�������;G8?J{�>I?�.>��-=�G���(�=md�Y�I�b��>&;�>��r�=�_����,!����>�?�[6>�g?H&R?��?��b?��.?'�?΁�>B��ƌľ�&?2��?���=~�н�W�29�S^E�>{�>��)?)T>�n��>?�"?3!&?ãP?�!? @>`����>��X�>B�>xOV����G]>/�I?��>6�Y? %�?�8>B}6��꡾D@�����=;�">��2?��"?�>?��>��?!+����>/l?ޥ?G�?�
Z?mս`�?>�?�R?O��=���>e8 ?��?8�J?�	z?`�L?�&?�0C<MX�'.�=�w��,)y=��;<� ��o]��!��m)>���>~g><>$�P�0�=ĺ�=Mi���x'=V�<�Q�>�tr>Ɖ��Y�1>�2žZ툾�A>U�e����L��+�:�+��=$n�>�j?��>�"��g�=���>���>���((?�?'#?&;�nb��.۾8L���>D�A?���=�l�����G�u���e=��m?T^?LpX�������b?�^?PX��=���þ��b����t�O?,�
?��G�4�>]�~?��q?̠�>�f�8n�����Hb�#�j��ֶ=,o�>�[�g�d��D�>O�7??D�>��b>�C�=�d۾˼w�Gj���"?\��?��?���?�8*>f�n�c4࿓�������õ]?��>Bɪ��C"?�"���Ͼ�V�����բ⾂����ǫ�����W��u��2�����ս1�=xZ?��r?�sr?��^?� ���c�_�� ��T����Ս��D��bF�F�\0o��������K��]S=[Jf�{K���?O�+?��i�e��>f�s����9���h&^>ik����x�*�=C>D=���=1}�=zL����l找�$?t��>�i�>�;?�eU��q=��98�0�6�����>f�>�9�>�a�>�ћ�r�H���x��������t�lz>�lc?��K?��m?t\��1� ���~9#����h����H>6�>�#�>�zH��4���%�b�<�z�r�~%����x	��=�2?G��>���>�ߗ?�V?p>������:k�AM1�0�}<V�>�b?�q�>���>R����C��u�>��l?7�>��>�Ό�u!�;�z��3Ƚ���>�C�>���>h(o>�*�_[��2���.���`8�+��=:i?�o��wYa��ׄ>��Q?��T;-�m<�T�>~�~���!����W�&��l>�R?%0�=�:>�ƾ���D|����)?CM?�݋�7�&�Z#|>K�"?]��>_N�>G`�?��>�S��I�y���?�;_?iNH?L�@?���>��B=����Fɽ�<&�09=X��>&b><�=���=�f"�4Z`�k���o=�ݾ=	�Ƽ���<�ʼ$�6<]��<�)>H�п�@H�:�侅���ʾG��TO��0&���&�7�)�2Ծ,w׾�M�?�,�C�\��f�����̠��C����?�Y�?�e�u觿,
n�'��`�>^�پM�k��K�z�����"�Ǿ����7@(���D�iȉ���u�JS'?Ñr�Ibȿ���r��Ӕ"?H�+?�X�?g}���%�b�?�p'>�� <���ޅ��j}��F
ҿ�թ��Q?��>�G�}�����>�5^>>92>:z{>�cp��̢�&XU���>Ck?Q�>���~�ʿ����Mr��	�?��@�yA?�(����R�V=���>��	?�?> Y1�U.��Ӱ��C�>6�?���?ZO=<�W�g:	�5xe?Oj<h�F�G�ۻ��=�b�=�=|��J>�>�>؂��MA��Gܽ��4>�ͅ> @#�l���^��_�<�]>�ֽV:��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�򉤻{���&V�}��=[��>c�>,������O��I��U��=���y�ÿ��9�`�$����=6H�}5Z��\ü�;��f�Z��s���Dw�l�����=*;_>GV�>��>��>0�A?;N?���>{�>w��jV�:|׾ngv��ћ�����r;�!7��Q������M���5�H�-���cط��L1���=f+I�Px���/��
m�.�&��":?5��<�d��#�h�R�E��u��S���_5=�E��9��i]���~��ٟ?ȨU?쎁��Ӆ��&/��-<��kPi?�dƾ����ۉ޾({�>�H��>d��>x�>��ƾ��L���j�	O3?Ln!?n���)����>��(.L=X*?8\?�=��>U?։��Ө���D>@1>��>�D�>GG>$�������?�[O?=	��<���qR�>h�ƾ]큾�	b=]d�=�4=�GGӼN>��;�ĕ���s
���+�d�W?��>�
&����ב��'�+�J=��w?�&	?�u�>��h?>�@?���<���[R����iA�=��Y?��k?	>Q�����ξ���g5?�ve?dO>*�p�wr�)�,�!-��?4}l?��?Dzɼ=\}�󶒿~�
���4?��v?s^�xs�����N�V�e=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?��;<��V��=�;?k\�> �O��>ƾ�z������=�q=�"�>���ev����R,�f�8?ݠ�?���>��������>�d��L1�?�<�?��������,���b��桾E_'���r=��=��1��E	��^�c���kI��K���z
>/~>p�@�.=�<x>��c�g�;|ؿVgw�����H�ѾbI#?��>=����&������4����t�LK�۞��<:�>1�>�W��1A��K�{��x;�/���[�>#�
���>�wT�V��z��Rp:<M�>���>R��>30��A���Ù?���s?ο�Þ�7��g�X?�L�?�q�?97?��@<��v��z����Q-G?'�s?�&Z?s�$�Z]�A�9�"�j?�_��vU`���4�xHE��U>�"3?�B�>U�-��|=�>���>g>�#/�w�Ŀ�ٶ�N���V��?��?�o���>s��?zs+?�i�8���[����*���+��<A?�2>���K�!�B0=�eҒ�¼
?[~0?#{�e.�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?ֵ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>dH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?F)�>��?P��=m`�>�N�=[��,�1c#>�G�=º>�d�?;�M?�P�>:��=��8�$/�YVF�yAR���i�C��>*�a? �L?�\b>�긽B�1��!�x�ͽ2a1��輠_@���,�f�߽�$5>j�=>A>��D�7Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*U����*���[����{>��f=��o=cͮ��f\�M'��=M��=$=?>R�M>M�>��>p��>�5b>ZD>$���Eu"��d�����6'���&�A���U:<!.	�9&;ݶ�g�����;S���3�p�-�Cv;q��+��'>	N?J�Z?z�n?���>��ݽ6��<�#�а=��%�v1>��K>�H1?��P?�	?Qӟ�R�w��c��������Վ�$�>��>*�?s�?��?g��=xY�= &@>���>�W�����qS���T���>�	�>�@�>_s�>�:v>�&�>E�ĿyRؿ/$v�X���rR=%t�?�*��p�������z+>����̚>U�{?&�>�c��m�Ϳ¸����6?>��SO�y�?�
�=3FK?z�R?CJ!>�Ƚ,�q��d>3t�_���}��H 9=�҇���N�X��>��?u�f>�,u>�3��j8���P�Vn����|>�96?�鶾�U9��u�>�H�rdݾQ<M>ؾ>+�D�yt�������si�X�{=�|:?s�?]���氾V�u��6���BR>�\>:4=.�=�PM>U�c�`ǽ19H�)�-=��=��^>�?��W>5x>���>#ٝ��IK���>�e>��>?�??s�?
0��@o����^���/��J�>���>���><�c>�5��<�=bB�>/�=>�6ؼ{���и��[,��|>ԝ�����b3b��<ڸ^�&��=��H=���$C����=�~?���%䈿��7e���lD?T+?Q �=�F<��"�D ���H��D�?r�@m�?��	�ܢV�?�?�@�?��2��=}�>׫>�ξ�L�ޱ?��Ž-Ǣ�Ĕ	�()#�iS�?��?��/�Xʋ�6l��6>�^%?�ӾPh�>{x��Z�������u�y�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?toi>�g۾;`Z����>һ@?�R?�>�9�~�'���?�޶?֯�?�6�> G�?�p?�g�>����s�a�)e��h���U���ؽ�8v>��
>s����u�tR��O|��yׅ�$D��'�=D��=���>�ϩ��9Ѿ�X*>fT���������.�\>�Ŋ>�=���>0?H��>��?���>T7��ѝ��YI�'�K?���?���S	n�⇼<x�=�_���?524?U<X�9tϾ��>��\?H��?�[?!=�>����7��a뿿,e����<��K>L:�>�$�>�J��wqK>�Ծ��C�4j�>i�>����~�پ�؁�О����>^u!?2��>ȸ�=�� ?o4#?<Nk>�߳>�&D������E�y<�>�>�>^u?ϟ~?G�?�����-2�"}���}��E�Y��O>��w?ѝ?��>�P��FE��/G��]+[��-����?�jf?V���$?k��?�??�@?�h>I��+Xվ�\��'�>��!?��)�A��L&�@��~?Q?J��>H/����ս|Xּj���~��� ?;(\?XA&?ۛ��*a��¾�=�<�"�S�U��c�;`D��>^�>����ώ�==>fڰ=EQm�I6��f<@k�=l~�>���=�/7�u���=,?MG��׃�@�=�r��wD���>sPL>=����^?�j=�e�{�{��(x��TU�� �?���?Jl�?������h��#=?��??�!�>�G���z޾���Iw��x��y�M�>���>�sl�w徶�������gF��t�Ž�,�[��>;A�>�?Z�>Z�c>��>_ ѾC?"��� ����j��>k:�<�I�`(A�b�"�.�ʾ ����@۽z)��m����_>�5�;�n�>�#!?���>��(>��>�!�=W�>z�>��>:1�>%~>� �>_��>�m>iŪ��KR?L����'���ȱ���-B?�nd?�)�>�>h�������z?���?u�?N"v>Suh�F!+�Lp?*L�>��~e
?B:=�5����<�7�����[��9x����>׽�:��M�^f�De
?S)?����ʡ̾��׽4�����y=�v�?��(?�*�=LR�f�p���W�C�R�����f������$� cq�}������+��˔(���1=/]*?~l�?����X�d��h�k�.�>��c>UW�>�]�>uɾ>&OH>�7	�p�1��?]�Eh'����LK�>�z?��>�S=?�1?�K?@D?��>�*�>�Î���?�='�>Ar�>�d?��=?*&?��>��-?�Ax>v��;X��� ���>��'?=�O?-@,?,� ?���m�_���ǽ9A�=�駾�$|����a0y=#M�͞�<�ٽ\ʼ9[?�p�e�8����K�j>Iz7?��>���>쏾N���$�<���>z�
?A�>����yr�\L��j�>���?3+�sT=��)>��=įֺ��=$������=f%��s6;�#<�4�=�}�=�s���޹��:I�~;�3�<�}�>��?ź�>g�>���Ł �����=8Y>K�S>�n>Ƅپ$s�������g�q!y>�o�?0t�?�,h=���=bq�=SU��it��������I�<Ů?�4#?�BT?���?W�=?��#?��>�!�3L���Q������n�?�x ?�d�>�$���X����0/?D5?;�`��3¾�J��о�=��q���u<����ſ�<�k�W����=����?�2�?�{=.�R���!��"�����?�O�>��D>#�>��;�9���P&��t�>��>��B?��>��_?rA`?��8?����)
]����Z꧿ h�<��B>D�B?DEj?���?��y?N�>{=%l���J�|x@�fB9��늾�Pͽ�C>f>��>[[�>�y�>h�:>�����P=�4�;�=�a�>䚺>��[>[	?P��>P�B=E�I?*��>����N2	�\��A��<�/�@{x?=��?�!,?|`=Mm�Ԋ<�D%����>O��?��?��3?:8��p�=��c��L���U{���>���>��>A>�=�=��=DE�>�:�>��<�
2�&�.�%���
?��E?(s>���������ol��&Al>d
����ȈC>�ļ�+dt�>�����&>��	���N���[ؽG���˽��Q��>#.�=}u�I�Y>�v�=�I����>$>�L�>�W<��X������]�=!y=[�= ˼2r����CZü�-˾Do}?�BI?��+?v�C?��y>�u> 6�7q�>�7_?N�T>1(P��M���]<��ը�TŔ�n�ؾ�W׾��c�d矾��>��G���>g<3>G�=m�<E��=�x=�܎=�r���{=�=�=�Ը=�=C�=��>m�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>Sq7>��>]�R��1�|w\�d�b�
�Z���!??;�'V̾ �>(�=�H߾�ƾ�[.=�6>N�a=PT�?L\�k�=�z���;=(al=�ԉ>.�C>gɺ=����U�=��I=���=��O>�k��x�7���+�"�3=���=��b>�&>O�?U�?��$?ò]?y��>Jg ��D���ޟ��t�>ʢ�>�q?�>���>6�>
��>ch8?��I?���>�eb>]�>3��>���)y���᳔��v2=���?�Ӆ?{#>=I�rm�0��Y�!�}|#=�G?�?�#?�ݡ>��ɼݿ/sU�#8C�ό�}M<}�ݽ�e%��t�8D���%f����Ʈ����G>��>�>%��>�"�>�O9>���>��e>Aff>P<�=�3����;���p�e�"���E=��0>��\<���0����� ����J�����t�=�>=���=���>A>I��>tɖ=_󳾁Y/>ⴖ���L�(��=�D���/B��2d�V?~�j/��V6�ϿB>1X>m��1����?��Y>�?>a��?�Eu??�>�8���վ?O��4)e�CuS��]�=��>�<�q;�jN`���M���Ҿ!��>�}�>���>fW>��*��9�<^=��ξYb8�ٟ�>���Ľ�!c�zo�����p����u���s�O2?`�����0=�[~?"�V?=�?�2�>��ͽ�����3>"�g����=�'��[����q��?�3?��?����@��B̾����޷>�1I���O����� �0�Fa�V˷�!��>�� �о�3��e�������B�{Br����>��O?��?f0b�cW��<TO�����?��yn?Z~g?��>OI?�=?� ���o��p��V��=��n?���?�=�?�>��K>rK'���?�(?���?2݂?�[?m���N�>��a>|v�>˰ľ��=ъ�=f���*j��)?��>��?��ȼ�)꾻��!�2��j���=��>�c>��>;��=��=��>]9>t�L>mD6>y^>���>�R�>�_���h��	?<I(>�5>?0?���>Y.=��]�{�+�`���#%�'�Ƚ��>3P߽*%T=�����=�~�����>H�ÿ�ʌ?Л�>��!��}�>�����o����>��>@D���+?��>�?�>��>��>U��>H��>��>�FӾ�~>����d!�e,C�;�R�ӾѾN}z>���Y
&�Ο��w���CI��n���g�^j�2.��<=��ʽ<H�?������k���)������?\�>�6?)ڌ���G�>b��>pǍ>�J��S���;ȍ�:hᾓ�?��?�;c>��>A�W?2�?_�1��3��uZ�.�u�R(A��e��`��፿𜁿�
�	����_?	�x?yA?rS�<\:z>C��?��%�\ӏ��)�>�/�';�/A<=`+�>�)��F�`�:�Ӿ/�þ�7��HF>��o?1%�?�Y?�SV�7޿�<?#>�a<?O1?��j?p1?��=?���҇(?�ZF>��?(V�><6?�[-?^�?�N >��!>���<�|�=�L	��b뽽i����E;�Z=��=��N�L=��~��TD=��=�=�?=c�<�bW=� �=劳=��=���>à`?q?�3�>��?0v&��A���w�MIJ?й=�Wu�:��7��(ݾu�=��b?F��?p?���>f/B���E�E%>��>�lE>Ա�>���>4�>��*���Q=���<k��=2H_=w %=�g��}������׽��B>���>� y>�̊���)>[6����x�5f>�;R��<��ER�ԻG���0�s v���>�K?t5?���=!�辧�����e�N�(?ȟ<?�:M?\?�c�=Փܾ��9�/fJ�D�rs�>0N�<ڃ	�fݢ�����ޓ:�Kǖ:�p>�����!����a>��g�޾�wn��(J����eMN=�d�T+T=P�w�վ������=:>
>�~��e� ��!��"ͪ��4J?�m=|m��N�U��˺�&�>a��>>��>�w9�D[v�x�@�����az�=���>6w;>�Y��ﾴ�G�h|��2�>�ZD?��e?1;�?M��Ef���B����{w��!�Ҽ�Q?���>C?ƾ$>zv�=�.����Ƞ^�[E����>�+�>_���1J��1��)4��PP���>��?�M>л?�E?���>6]?�(?-�?�s�>|��������&?f��?]��=�Zν��W�g8�?+D��.�>�)?�?��R�>Q?�I?�o%?ANP?�s?W>>$���2>��(�>���>}�V�O߯��1V>�>I?�t�>s.Y?�Ń?t�;>e�3��9�����0b�=b+&>�u2?�!?>q?d��>{��>��վzr�98�>s�?I�?�l?�^+��>��>�?�W�==`
?x6?.l�>�2?�uc?ZU?�1?��=��<��x="輻��:\=�	�"-�����]� =�� ����<����<n�U�<�=�h$<i-=��L=���>��m>룂�%{<>�����"~���<>�͞<������}���1�ƛ�=�)�>�h ?>ߙ>Ë-�oѱ=�]�>"�>4��k$?'X?�V?0�[<�L\�]|�L�q��b�>��C?�[�=F�e�xۑ���q���r=F�n?��[?�B�
2����b?��]?sf��=�[�þ�b����?�O?��
?��G�-�>��~?��q?`��>g�e�:n�����Cb���j�g˶=Sq�>�W���d��?�>��7?�M�>��b>�#�=�v۾��w�r���?��?G�?#��?,*>Z�n��4�������ĭl?�i�>-�Ͼ�m6?��+<qpӾD�i�������)�0�̾T ���.��l�:�����V�-��<>�?�*v?܀?;CS?�H���?�V�\��Yc�3�,��!��'���W� ��j�<�e�n��;J�u������4	>��-��6���?^�)?_^���?�a����pϾ[lw>�N���Ľ��=	����ڮ=�t�=U��s�3���-?V�>xM�>d6?��9��%<�M�&��i*�c��}�`>���>v]�>�@�>ךz=T��?��;����t���&�7e>��f?��E?��X?+�G��:c�bj��^�N���'����xv>��T>���>ڟ`�n����z]��$e�㯀�Q\�n�����"��o.>>? o�>��?3�?��>�) �����	�#�.��=[��>ʽn?��?��>�p.��&'�G�>�gm?K��>��>����zR#��|�y@ս�y�>5A�>���>�r>��*�<F\�CS���	���):�QW�=RYg?�׃�
�a���>C�R?9{�;"P<%3�>�%u��"�z�����*�Gk>6?�;�=W�<>O��I���{�K���)?�		?Fф�!��hc~>�?:��>��>�ۆ?���>P��Y���"�?O�X?O�S?��<?��>���=�{��ە���X��
!=�ʐ>��v>\H=�6�=
g��E���6��i�=rQd=L3�<�����4t��D��;�W=�Z>Өۿ'PL�~پo�����Uʊ�<�����B �Rn���p��u�	r�PT>��QT�QCg�׋���h��5�?+��?����c���n��鑀��x�����>�"n�^M��Y8������ �����{��i���N�i�])e�۔'?�����ǿ�����;ܾ�  ?�B ?e�y?v���"�q�8�� >r0�<'.�����w���(�ο������^?~��>~�'��.��>ҥ�>��X>�Hq>��Ꞿ�!�<X�?*�-?j��>��r� �ɿ�������<���? �@��S?Z��,��>�s?ʨ?Yр>��=��2C��>1��{�>�Ʃ?�R~?�:>�;�5�=Nj?ʳ�;�83��
�=}>�=���]}@=u1�*4�=�>���@����ϼ4
>L�>����5ډ�K���h(��Ȓ#>�~���%�2Մ?{\�if�v�/��T��	U>��T?/+�>+;�=��,?.7H�b}Ͽٯ\��*a?�0�?��?�(?�ڿ��ؚ>\�ܾ`�M?_D6?���>�d&��t�/��=�0Ἦ���h���&V�k��=f��>S�>O�,���W�O��H�����=;�
�K�׿��=z5�c¼Xo���d���f���7��Dk:��ݾ�>ؾ����=t��<\�>j�=<S��=:��>�L?�}C?���>>��=$\�;��Ǿpp��O_�9�4S���D��K����+>�8V�6o��&���"��i� �Z@����o�����bX�����\��y��u�%�#?uIo>Ф	��Ζ���I>ca�������~)=D���X���1�����?M:z?!�z�D%�|~�=z�(�}OA?��+;J�������==�O>�m=ڝ?t� >J"ľKu+��=��@=4?�}?�t��(���]4>�_��xJ=W�*?m��>mS/=���>e�$?���IL��"�e>�C7>��>��>��>}��.kսV�?P?��Y��c<�>����Z����=p�=��0�����V>2�!<f��l"t��'��;P?5s>/�ي
�V���;��>��k?���>�Ǘ>">r?9�6?��<0�߾&�H����i��=ii?ɰa?���=|��Bg��h���P?�Dr?ͰU>��0�v辮�6���7�?�b?\� ?9��<�jo�ۀ�����פ&?/�v?/r^�`s�����&�V��<�>�]�>���>g�9�Pj�>��>?�#�G��+���Y4�?.�@���?�<<'�ښ�=�9?u\�>��O��=ƾXt��O���`�q=v"�>J����cv����jP,���8?���?6��>�������=P��,��?�z?֗�&#�=m����h�����9�	�	�����+�������Z��Z���;����>"Iw>��@��,��0>��U������jȿ;=y�L;��y�;H?�^e=�<�������@ꋿ�Mo�w_^�5�,��A�>|$!>��S� ����|�4�5�L�T� <�>Ƃ�;���>�E)�⊹�h`���sκ�ɓ>r��>�n�>�&^�7���|b�?����y]˿~A��dP�K?*l�?�3�?~z?���<L�e�:)v��hr<��E?-}p?�R]?C���x���XW�%�j?�_��xU`��4�tHE��U>�"3?�B�>T�-�e�|=�>���>g>�#/�x�Ŀ�ٶ�=���Z��?��?�o���>q��?ts+?�i�8���[����*���+��<A?�2>���H�!�B0=�TҒ���
?U~0?{�f.��^?cQ���e�I4'��s��$}�>SV9�C�O���%=��۽~Z�)�w�U����?I�?M�?,�id�p�#?�w�>䵰��|޾���=�T�>�>�Q>K)��#k>�?�E/.�6�U=}��?w��?-?P�����P	>��q?;_�>�`�?���=�9�>u�=q���6�8�?�!>�=ˢ �g�?��O?���>���=�2�S-���C��Q�rK	���C���>�<`?��J?Дc>+�����?�:z"��ﹽ��*�� ���F�i=�$�� 2>/7=>Z>c�B�Dv׾��?3p��ؿ�i���p'�}54?���>��?���t�j��u;_?�y�>�6��+���%��uA�i��?�G�?O�?Q�׾�e̼�>��>aI�>��Խ����c�����7>�B?:�RD��3�o�t�>���?�@�ծ?Zi���?��T���}���Ǎ5����=)7?n�𾒊y>���>�ܨ=�jv��_��K{s�/Ҷ>b�?�?�?
��>�l?@o���C��4=pݢ>
�j?��? �U�@>iJ?���x�������e?H�
@'G@�_?�����ֿy���~��y���`35=S�=,�D>6R.��=���<@�Ӽ#�ǽy���D�>�R>�[|>��W>ճI>�!>]Q��j�'�0ߴ�ge��c�V��z%��A��3���%���a��r�O���8[�i��<T������}Y��-O�Od���0�>�N?��7?'sk?��>꽫9B>���\E���,=cҷ=iX�>��J?�)U?�X?��=�x���P��u�����ŋ��!��>�.>&ڱ>�$�>T�>����hV�>��=�ul>V��may=����Q�̆>���>ȅ�>
��>G�[<)n�>X�ڿF��޻j�,�w� >����?Dy�=>\K�̳���*>�s�P����^?�>+���Y|ǿk�ֿ[�+?����F���1>�I���?1F�?r�>̉���,���=��9�ǆ��	7U>w��1���Ų�za>�'?��]>i�q>��3�ą7���O�ci�� z>��4?�ƹ���H��]u�_�I��I�|�?>#��>FC���w�DҖ���}�{ck�{�V=QW8??��������7��U̠��yX>Md>#V=r�=3zN>'l@�T�ν��A�RNi=�y�=�Ma>.u4?�1�=��>>�I�>k��������>!��>����L6?�
?��`=��L>�VV=�; U,>���>�ɿ>P��=�V��=��>�=>�ý ��<EH���Ƚ4<=�y��s�\��]M=f/ >����0�=iM^�E�.�C�������~?Y���㈿���]���lD?�*?B�=[�F<�"�����wJ���?;�@+m�?X�	�>�V�~�?�@�?�����=�}�>�׫>�ξk�L���?0�Ž�ɢ�Q�	��'#�
S�?��?"�/��ʋ�3l��8>�^%?��Ӿh�>�x�jZ��W����u��#=ĩ�>}8H?�V����O�7>��v
?s?�^򾯩��F�ȿ~{v����>4�?���?�m��A��n@����>Т�?�gY?pi>�g۾�_Z�d��>��@?�R?��>p9�]�'���?߶?���?���=�`�?"Qj?�T�>�{�����}����ґ��=�Ž���>�">��ھ/���/Ӽ�����A4��A��h��>��_=���>�a�aX���6 >�ޙ�=a��*�����>G.)>��s>[@�>\�=?��?^�?�=����1����M? �?t��U�i�n��<3�={�R�I#?�/?	+y�[�;�>//]?�#�?~(Z?��>�w�a��b��ǘ��ٕ�<HL>��>��>s#��&�A>%پ��9�)��>���>Cv�^�׾
���Y�Ố(�>C�!?���>�T�=� ?Μ#?7�j>�'�>=aE��9����E�ϯ�>���>RH?��~?��?1չ�[3�����桿
�[�o;N>��x?�U?�ɕ>m���e���i�E��KI�� ��?�sg?�S彼?�1�?��??(�A?�-f>���ؾģ��6�>;�!?/��ˢA�&�����n?�Y?���>)����2ս��Լ����#��?6!\?2&?����a�D�¾Z�<�"���U����;bsC�*�>��>u~���մ=��>�K�=��m���5���d<�U�=�D�>��=�F7������v"?��"=��O�!��<�O���IH�],f>Cwh>1b��G�\?�)�x��۔����X����?j��?f��?1{��?Y��^7?�{?��?�H?��ğ������X��#ͷ��-��.�=���>�N�/�德������.)���ĽZo���>�/�>��>��>h�3>1�O>�'����"�O��Y���!p��<���=���-����f��tK�qS������s���3PV>��=,ǟ>�-�>�Ƽ���=(�?�H>���>�->���>F��>6>n�[>��>��a>�V<eiR?����w'��C����nB?�se?`��>Ý��x������ql ?���?G�?~zu>�|f���(��v??��>����"�?�FB=����6�<�ڱ�4�|���L4���>����}9�n�I���b��M
? �?i�|�m�Ͼ�轜ǣ�x�>t�?i"?�q5��[��Xs��U^��KD��ý��C�V���f5�/�����*���@∿��*���>)�?��?��	r��묾�߉�Ja9�:NJ>���>+ï>���>�:>>~վ��C�/Ro��:%�~��v%�>²z?�r�>�vK?e�7?��M?�F&?c�P>'�>�=N�N��>q�y<�*�>�>ЎI?e%5?b�?�=	?QV*?\g>�)�9���+��?��>��>���>�| ?�x�>���>f;9�}�;p���b�.fZ=�"�=�D>�,sA���>�U>��?F����:�6����;V>�K3?�~�>T��>$F��$mu�{@_=�&�>�?�>mL���Ym������>��? ��{r�<��%>��=�w�;駓<]��=�d�n�=�93��@6�0�<}��==��=��d���<���
�j�D�[<���>�w?�ޅ>��>w���/��1�
�bH�=e.T> �M>bu">
�پ�ۉ��'��U�f��y>TQ�?��?2�}=i!�=��=���5����DH����=��?��!?��S?䇑?i=?��$?/�>C�ɶ��7������#?���>���>ޡ���l��"�#���C?��?f�U�����j���̾Բ����>�/����v�5:¿ �m��d*��Q)��@*�h��?	ͮ??U>f��j�9������>�N ?F�j=�ټ>��c���J�0��P�>0��>mij?R�>�O?I�z?:�[?0�U>��7�]i��3Z���b��#>�??-Q�?�ǎ?�x?��>�>]�%�� ߾(b��x�#����?9��:&T=k�W>w�>��>qn�>n�=Jf˽x髽�_@���=�2b>�e�>E�>���>f]x>���<d�=?�P�>�Ò�����Cg���t��ٯ��j?�?z;?�#	>��/�%t���ƾ�+�>D2�?�W�?�7?����>�9��Q��f<�ֶ�>Ą>Eɟ>��v>kl��}>�a�>{n�>��-�U��i�1�pʽG�?@�A?v��<
�ɿ�]|�<-|�樨��<�<Op������-}�0O��x�<�:��Y���y̾��l��o������&Ⱦʵ���H�}"?��=�z�=2�=�3�=�1�����;���=##W= Ȁ��m���;�=��ռ�I<��U��<!�<�H�<���<V�;*���6v?�VW?߳,?�U=?/8�>a��=����6�i>�'ٽ�?�\V>����<ɾz�G�4kž��N
ϾϷ۾�MQ�����>����d��=X�I>A�=L�<��=�� >b��=�n�3ɼ���=n`�=O�=B�>'+5>�# >�6w?���ֲ���4Q�RZ�v�:?8�>{�=��ƾw@?p�>>�2������nb�.?d��?�T�?H�?�si��d�>���v掽
r�=����>2>���=&�2�g��>��J>���K��g���m4�?��@C�??�ዿ��Ͽ#a/>��'>� �=��V�7�%���w��kZ�Y,=��?�0��
̾�>��=�ھy�����;m�%>���=ԁ���J���=ZX��%�C<�z�=��>�9>[f�=c?����=b��=��>��r>3<�=j�3�m,K���<n`�=t��>��>U�>EU3?��@?y:4?�#=>!��]���7�����>��$>w��>+(��
> n1>@�?2p4?�UM?.��>�H>É�>D�S>��$���}��n��eؾ0C=G��?w��?���>'w�=�HֽsZ�D��^Q>��[?_cS??�/?l��>WQ���7D*��3�B擽�Jr<��"<L�H��?o���!�e%-��M����;)��>�#�>Y�>78V>9?,>D�a>�־>�>��=��m=�P�<�=���^�=�Y����=�$W��1*�7r'�����&a������e���U =2/�=���=�}�>'$>U�>��;����7�>�Ds�f<6�/@�=I�����G�^ ]��w�3���C��56>x�h>����ي�a& ?z2W>(a>��?��k?�A�=��ڽ�kھ������p���M�G�=#��=YqS�ٰG��rs���X���۾��>c"�>�͒>VM>y*�rg8�`�=��վ�N@�	Z�>5p�����;�'%~��硿W"��em�M]��:�7?lǈ���O=�t?YOQ?��?K��>e:�����>��n��g>V���o�oإ�<�
?qK(?��?%L˾��7��̾����}�>�vC��J� ���X~*���Ѽ�ѹ�:��>�5��M�ؾ�J5�gZ�����t<�]�a�P��>s�J?�{�?�/l�J���:�D�U��-7�����>*�`?�>�>@�?s�?�a̽[E�+Y�H��=�*n?�W�?�_�?TR>C��=a
�)��>��?z"z?@�?�*d?�]��.�>���=�>��/�=9�=��;m>۱?�y?��?L�%��B ��Q�;F]��8��=�b>2W�>���=��F>�� >1P�<��)=�(f>��>d�>�J�>Ì�>R?�>E:žݖ'�Z/�>��>�^>�t?��=�e����F��D�<CRO=�� ��y���F�T�x1�=a	=N��=K��=0�>ccĿ��?±�>D�����'?&�<f��\��=,�>�s��u�,?��>���>.8�>�M�>�>�[�>�\}>5LӾ�l>���`!��)C�%R��ѾRnz>Ꮬ��&�������RLI��l��'j��j��+��G7=���<�D�?�����k���)������?$Q�>�6?�Ō��Ո���>"��>�ٍ>`0��ύ��č�q\��?M��?�a>z�>n�W?��?1
4��73��_Y��u�޹?��c�F�^�砍��Y����
��9����^?��x?T�@?^d�<B�z>��?�&�����I�>��/�Q%9�k�S=�>�Y��Y3`���Ӿ�(þGI���I>k�p?VE�?��?��S�ЀQ>�>�G?�9-?�`?G�'?�@?1��B�>��Y> � ?���>��J?��,?�"?��=�/8>#�<��!㽈��S.���0��JW<��=���=)�P��4>H�W>/�'�����!_��}�e㼗P1�������3��=:_�>[�^?�?s_>� ?��4���+�s����@?x��=?�vƍ��逾�뾮�R>.�q?�W�?��Z?y�l>��-�8�p��)G=��S>�0>�N>zE�>������*�=/�=��+=���=��޼�����l���B�=�>���>2�>ӗ{�2>ɩ��&��K�Z>�MB�_+���`R��E��)4�\[u�� �>��K??f?�ϗ=�>��3����b�#(?�:?�M?�?��=\�߾�5��K���=�{ۛ>J�<�a
�����8����w>�gM꼧�]>�k���6���3A>g��R����o���I������=�e�ج�=%f��#���y�,>s, >B�Ͼ�x �NC���Q���K?'>�/��(�H��ɾF�=�k�>�N�>j��AA:�U�:�z��!�<z��>��?>��5����A�S�H
����>�E?�:w?ǭ�?_�����m��}7�{Ͼx�������?��>}A?�ܒ>��>$ƾ)16�����,����>���>�|;�G��žƟE��n㾰|?H�w>Q�>6)?�Q�>��8?r��?JGH?{� ?�j�>Iv"�J� ��-?℄?�-=�y=�G־��S����EGB?}?�lQ��O�>妳>a4?uF?V�d?m{�>w�A=� ��X��T�>qQ�>�h��ҫ�<�=|�C?T ?�:U?��?�$�=9�%�c7��è���"�=�mZ>��!?�!?(�5?m߯>)s�>G���7�=��>�xe? �?Y'm?��=�
?��+>&o�>/&�=���>Ȋ�>ڲ?�O?�Gq?]J?��>n��<�箽C ��M)q�q�����;�8�<\=�3��+w�F�(����<�̥;��� �����;�3�󂼵�p<'j�>�t>���1>+�ľf����@>K塼�7��%����:���=���>�?ӕ>W#�ޞ�=>��>43�>���� (?�??#_7;͍b�K۾�K���> �A?*O�=�l��u��}�u��0i=,�m?�x^?�W�q����b? �]?V�=���þ��b�}��K�O?��
?A�G�M�>��~?�q?{��>��e�?7n����}Fb��j��ض=�o�>5W���d�;3�>C�7?qW�>��b>��=�v۾?�w�
w��g?��?�?^��?.*>��n�"1�4`���@���^?��>�1��M�"?���ֽϾu3��>뎾e�\���,���Z���~��|�$�V���ֽ�W�=�?�$s?�@q?��_?�� �/�c��=^�*���qV�t�����E��E�H�C��n�im�D6���'��LUG=DZB�8�1� p�?�?�rν1j�>$*���eվ�n���4{>I¾/�������m��B=1ˠ=+,,�Y�ν���� ?�/�>�>4�Z?��a�-�8�՟H���-��L���>�ø>>���>Џ�u:��K9(���ݾ���7#�z+�>8pV?ǡR?��?�#����Fw�����5��=p]ؾ�Xg>�G>-Ӕ=449�iBH��QH��O�e��y��凈��U��%/>3�?	A@>{?�/�?mߕ>�b�h�����J
��>�*?t�v?q��>��;>��������>�s?D	?�z�>^��u8��|�����<�o�>�|�<�� ?P�e>dR��h�]�5���>���6��=�R?�pX������,>?�O?O����+���>������+O��ylN�->�>C�a>3�Y>`�׾�v�$�g���"���)?6�?a����#�Fh>2?{�>lS�>���?2�>N/��[i�<�P?ʰb?�oN?P�8?J��>�i.=�.ǽ��Խ	4�1�'=@��>�p>��=��=�0��^X���&Ih=b��=[���,�����мd��<O[p=L�A>�
ʿ4�W�*���ހ-�>&۾%�����*�=�-��򘃽Ӷ��큾b��NC?�tm뼥�_�׻m��ӕ���佋J�?@��?+O���૾����>S��qY�3��>�z�+#>!��f����N������຾�/��R�HҌ��
?���"?����ÿ����*Ҿ1�?�)?G�^?0<�>v	��p<��\�=F<���ӫ��>��%�˿9Ϣ��=z?z�>k�ԾĜ�
�>7#d>b�g>�<>CN��mB���̨<~j?�;?�?��|���˿�渿TJ%<z�?�4
@[|A?A�(�0��	V=?��>ё	?��?>�U1�\H�k����Q�>q;�?���?�TM=X�W��	��e?r�<��F�޻��=cB�=�5=��ȖJ>]V�>1��MA�'>ܽ�4>�Յ>o"����&�^�|�<�]>�սiA��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6��{���&V�}��=[��>c�>,������O��I��U��=�A�8�ƿa�#��Z!�L@=X��;\L�_&ǽ����'�j��k���_f��Fн��{=���=b�P>5!�>GW>V�Y>ίZ?9�k?�A�>5>�����А����R1�;�ɑ��������+k"�n���y�MB徠�	�&��g��ݾ��<����=��S�y;���N"�5b�$C��s0?8�>��ž3�M�2�;�ɾ�t��D�x��y��x,;��3��l����?lD?`3����T�f,�W�����V?�Y��{�T���_K�=Ł鼍�=��>mÚ=�S��{5�ɴT���1?�-#?[L������>$��ޅ= *?)8�>w�='w�>�"&?���f�$�G�>��>�~�>W��>I��=5Բ�����!?sQ?����?����m>���a�� 5=�Z�=\�0��xp���H>�E7=�|�
��Ow���9=(W?o��>��)�d�,b��Y�?==u�x?.�?J+�>d{k?��B?���<Vg����S� ��bw=��W?^(i?�>����	оc�����5?w�e?t�N>�ah���龲�.��U�%?I�n?5^?�}��v}�!������n6?�҇?�G�%ư�]���0��3�>#�(?���=h�h��*?�?�M�势 ���ZV���?��@���?��L>�3ộ�ռ��>$#?Ħ۾vUu�}^����u>�-�>��	����@�"�O���p?�}�?J��>c���|*x�u�>��q���?�?߳��� s;�1�}�Y�>~ɾZ;>���<}��S��=�2E:��w��b�ܾ��j����&	�>�.@��4�>�?�|��gMп!ʿ�C����ɵ��s�<?��>1X��;��:���~���?�֥?��م�8�>��>m}���0���|�(@�ý��q��>�M!��)�>�<�B
��6����=���>N��><�{>Ȟ�uKȾ#ܘ?��b�Ͽ��L��|�S?�נ?���?�?��;�Zp�4|���KܼU�J?�qw?�W?䇽�ΒJ�=�|�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�M�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>lH_���u>����:�
i	>���?�~�?Qj?���� ����U>	�}?)�>	C�?���=��>���=P�����:}(>}>�aB���?<K?�e�>�X>���"-�M^C���L������@�t�>�Ie?WOI?M�m>.벽ŵ�����pý�<�y8���C���,���你<K>�BL>�\>�O���ɾ �%?����g�տQ������'?�ݼ>�.�>�j#�'D9���V�b<?��S>U��弿�3��b�ڽ5�?-$@"�?־��ݽL=r>�R�>�G�>�Y���A�<>7���6W>�1K?ɢm��,����f�O�<>���?}�@���?�銿?���$^���p���.�R"q>�[?%��k�>��>j��bt�����m�����>�E�?���?��>�m?FRs���?��g|>�\�>4g?�j?x,>�x��p;>j�?|���{���#���T?��@|�@4�Z?aS���;׿�᡿�����*о�X�=v��=Ԟ=�Ѳ��>_���S!>�1H>9y>f�>Q�H>��2>�o�=�KK>��J>�Q��r�'��蝿���J����Di�>k���e꾇��dH��d�v���U��������ӽ��_���[��0�8>uW?�LU?�]?lG?C�G=�X=;��&1	>�:����>��>�a?(j?�9U?T��=`Q����X�G���!���є�J��>~��=���>���>�܁>齢Ί>GB6>�Sk>��>�F�=]g��8����H>&Å>ߙ�>���>��;> �>Ӵ�GJ��v�h�}�w���ƽ�?�螾��I�h��/���*b��:h�=�!.?�1>x�Jп����7H?�Œ����*���>00?3PW?>�>�Ĳ�
RT�Kl>��
��k�ۍ>���dyl��S)�(VM>�[?/��=M)>�E1�n�3��N��� �*��>R"?a�>�G�&��i���v�����1�>&�y>�$��������a���#���<!�;?@{'?1˼=��ݾ��)�f/��lW>���=_ =K
�C��=�r��W���.�=�vI>66�=i?��?>���=�%�>�Ҟ�9�`�鯨>2K>��*>YE=?�O*?t������+a����ysg>h��>Í�>L��=4]Q�p��=�u�>R�g>�$Żvń���#��8���\>�S��Me�C���V�=����4f>`ǣ=_S��:���Q=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>�[�S����J���Og�d����>H�(?M��6��<0q`�O?���>�������4˿�~y��/�> t�?�A�?�:\��L����6�M��>N��?&�F?�q0>Íپ��)�Z�>WBD?��M?L�><�%��/�H�?փ�?o��?��t>�U�?'>|?z[�>���5/�􅿿,/����=`���L�>hW��k�z�@�ak�����Ϥ6�L����>�*<kI�>I
��0���>�d3��9���;��>��V>��>j|�>��y>ͭ?>���@������sI�[,P?���?���<���I������zq�J;)?�"(?���Eb���V>%MO?�܅?�j?*f>���Z�������s��#_�<��>{�>E��>�7=֢<>y���
�6�>�ޯ>�I>0��p��5��])�>P�?��?r�>�� ?=�#?�k>抲>\E�*��DAF����>�R�> �?�~?�|?;7���L3�n���{ء�f;[�)O>zx??Fܕ>�g��-S���<4�_K�b������?�Zg?+�轳�?7�?�A??�A?H�f>���@'ؾ45��4�>N�!?o��ɃA���%�IS���?1�?���>씽��ӽ%lμ,��:����7?4�[?´%?�y�	a�MUþ�y�<C*�1Q��E<�-���>Y\>������=j�>x�=@k�e6�x�o<]�=_&�>��=�45��L����@?X�;I�Ǿk�>�l���L��ns>oL���Ͼ�d?a1#���E�k﾿����N�#��?a�?D+�?��5>/�y��e?�y�?'�>ڨ�>\���_E�8���j�=(8�A&�C5>r�+>Hb���h�� ���������w����_뽈�?j��>��>�K?���>a*�>8���9�	�����j���U�����V���2�ə ��!P������?�~��'E��A��>�^1���>�_?,��>yf�>S�?\�i�=_]>8R���>~~�>�>Q$/>�I>Ѣ��yv��KR?�����'�d�����E2B?�qd?�2�>�i�܉������?w��?_s�?�?v>�~h��,+��m?=�>$��q
?�W:=�A�mF�<U��J���7����Ҫ�>�D׽ :��M��nf�5j
?c/?:��\�̾�8׽�T��/�u=�R�?r?)?/;*��sQ��*p��W�T�R�w
��De�M��#�$���p�m������Ȇ����'���=�)?� �?�q��\������j�Mb>�HOg>UV�>��><H�>��D>��	���0���]���'��Ճ����>h�z?�ͣ>�N?7
8?L�O?��:?�>>[�{>]/����?�M�:��>�@�>(�A?u�J?|�[?6�
?�}?�>Q�1�/��ξ=VD?D? �=?��'?+% >�Ӿ��'�d���#:��v���:>9�`=�>��<�S��ȷ&���+=T[?Y����8����T�j>�j7?���>.��>8ŏ����ԯ�<0�>��
?��>�f��
Sr��M�1?�>���?�����=e�)>�<�=Cn���Aк��=	�¼���=� �� ;;�1 <n��=��=�5r��m�S� ;U͒;/�<�@�>��?N�>Ш�>\Ώ������
�a��=��Y>� �>k!$>��ؾNX��I����Jc��P]>�?(��? 7��ø�=,U,>����D,��3����Ⱦ�_�N�?�??�L4?`�?�?)?G�?�l,>�������~� ��{�
?�,?��>���[�ʾ�Շ3���?(\?COa����<)���¾��ԽG�>0O/�%~�M ��d(D� ���Z���������?��?Y�?�H�6�no�Ø��N��6}C?��>�5�>i�>��)���g�p��0;>͋�>�R?��>)�M?���?��U?�-�>�������י���I=�П=��9?�K�?Z>�?�@~?e�>�C:>{�C��7�W���)�N���h����<R�G>ٽ�>���>�J�>ڧ6>����W���Rv=�3<|L�=dg�>D��>T��>?_�>�� =n�G?{��>-�����x֤�_˃���<��u?��?k�+?x�=�r��E��2���[�>�b�?��?w1*?��S����=��ּ۸���Oq�r��>�ù>�>q�=�HE=�>��>��>n5�NN��i8���M��?j	F?�P�=si��"Sa�-Or�QT��p=/�ܾ�6�]�ν�b����4>�H�������A��f9	�����u���}M��\V������f�>q5�=0��=o��=��=Wyy�n$�=E=�2<�>>�����=l?����):W-�˫�:=��?��=�U<Ag˾�k}?�(I?�+?=�C?�x>U>f3��[�>8A���4?�'U>��Q�:\����;�������a�ؾ��׾x�c����77>�H�[>63>Ճ�=�<	/�=��s=	s�=�rI�K�=<�=��=�_�=���=>�^>#9w?���������%Q�v��Ѽ:?�B�>��=1�ƾ�"@?�>>�/������j�&?J��?;X�?��?�Ci��W�>E���?���r�=����'2>/x�=�2���>ٶJ>����F���೽�/�?~�@y�???���l�Ͽ�a/>�
1>�2�=��O�i,�J�[��~��:�&%?k=��d¾&t~>�IB=�/޾�ۼ�m�=��'>N�F=�.+���Z�I��=����\�R=��="č>�O9>���=�(���=�Ɠ=/��=O�G>��B�\d�x�M��>=>D�=�(o>uU>a�>?��8?	�\?K��>"�=�Y�վ �Ͼ�f�>e�U=]ı>�k�=X�y>���>|??E?��<?�W�>/1�<P۰>z�>C�%���i�yO�	������=m��?䍉?-�>��=8�d�Y�2���O�Й*��$?^ .?{?*��>Hl�|��k�QS�#�;�/?>�û^G����+>�W����=�ϐ>�>�V�>�f�>��~>�=6w >A#>�T�>�]>G�<
7=b%=�U1=z�<sx�=M�ͽ"O��`��
ǽd�<-奼�.<��(<���=��c�V`ټ��>x�>&�X=L\�>��>8Dy�(f4=�pؾ��6�� �<��쾘��(�x��̐�W�-�� ν�h�>���>2�ٽ ���ͭ?�k=>�q�-��?
Ry?�-7>��<rŌ��l��bS=^��c�>��=�ʏ�ƖN�}�p��BF�c ���>���>*	�>`�l>�,��!?�A�w=}⾮_5���>z�����Q.��7q�?������=i��KԺ��D?�E�����=�!~?b�I?�?}��>���d�ؾY70>�I��߻=��� q�}U����?t'?Д�>�쾝�D��F̾��-߷>W>I�9�O�/�u�0����gͷ�4��>���[�о8$3�hg�����"�B��Kr����>��O?��?�5b�oW��9TO�s��+��q?D|g?��>�H?�A?�)��<y�p���r�=2�n?���?U=�?�>1V�=����K�>;6?N�?w�? r?�@�d4�>B.;�">�p���,�=�i>l�=u��=�j?$�
?N�	?�ϝ�^�	�����j��P]��-�<V��=�f�>�ъ>�r>�|�=�mU=�-�=��^>Vj�>�Ϗ>��e>ޑ�>�[�>n�j��DԾ*�,?+E�y��>�'3?gr0>������>�>����c�ľ읮�����a�,��1 >��J>��K>�+
� �>1Iɿ*�?j�g=V� ���y>�qվ�=�i>��>�Uν�?�q=Uy�>�?��>�'>�V�>Nh�>N����b>���%�����/Q]�u�콃J\>���EX�=r���*���쏾&���u��<�e���v��'J��5�=�a�?���<0�p�ZR��!<���?b�>c�?�i��s̽2��=��?��>�����H���6��R����{?l� @�	c>X؟>rW?W@?�,���-���Y��Gu��X?�T�d���`�A��㍁�-��=�ǽ-_?��x?`A?NAL<�8y>i�~?��"��U��i�>��/�dW:�?�A=Ө>����dza���Ծ��þ����CI>p�n?�ԃ?�
?�Q�J�=��*>:�>?�Q�>\�?���?��
?]�p=��d?C���?�>>?��6?�:?��:?p��>yE�s4|�}ж=������o���2l=vH>��=#;b>�y�ar=�"���,	=��/�S���-;�<9�h�#�=�v>�Qz>��>��Z?u��>��{>�a9?hh���6�K���/?��D=?Z��"󉾉��������=�i?u�?�Z?�4S>�)@�"cC�Ӎ&>~��> �>nW>��>���CL@����=v">�U>5t�=�C$��y��a��)z��Ν<��>s��>�S|>~	���'>ɋ��ASz�t�d>�Q�Ǻ�
�S�e�G�D�1�idv�dj�>��K?��?�l�=ae龻���=f��$)?Z<?BM?��?�J�=��۾2:���J��0���>��< ����������:�o�:��s>d$���Ȼ�L20>c��3ﾅ�p�/�C�������=�:�+��=����g����>��{�=�9�=�վn+�vۗ�vۘ��`C?�/�=����w�q�N�NtE>� �>צ>q�6��ԭ�E�6��[о�Ù<�>Bk>�EF:���0�B����ٖ>�.?Mn?�?���h�E���-B��N�i�1��	?��>l��> g�>���>c�ᾚ�%��z��%E����>�w?#�.�l��;ľ����ھ���>��]> D�<0��>��[?�s�>��?�8?z�>�Xr>��>��N���p&?��}?j"�=����ԉ���<��r���?\�? �Ҿ�mX>Aq&?��?;?�qe?:��>3D8���"��vG���>,�>��r�����>j3C?���>�J?>{v?��e=y1�+-q�S>D'�=�l�=ׂ(?��%?2$6?��>��>~㡾�	�=xC�>N�c?�P�?C�o?��=?,>׎�>|r�==N�>m�>�u?g3N?s�r?}tJ?���>$��<ȫ��@���>w���T�8S�;YP<��l=� ��p��n���<a�;�Kڼ�]��T�ʛE�㻜���;���>ʙ�>9����vH=�
��m�k�>�Ϝ�8j���tw�0{���=�x�>߱?3̟>��o?|=+��>P��>�
�.�(?��>�?R��ck����!W�A��>F-P?�6>��`��W���|b��< `?��M?�k����Өm?�,m?�V߾J)N�
�����Q�@( �^,?{H?W໽��>�#{?�?��?��7�ӼZ�����SZ��s���=���>�~��"�@��0�>>�+?U@�>��>�~>-���5=^�Vt����>�Ê?G�?0}?��>�q���S���W��o�[?��>� ����"?�,W::mо�1��Hݍ�J
��㮾�r��"������~�%����m�(2�=d?Kzq?^o?a�_?V� �Ɖb���]��>���U�����0�x�D�B{D���C���n�����񾪼���}q=�V��5�a5�?$�	?MyK���>��Ҿ ˾�L��F�=�*��&ǹ���=�v���xѻM�A��G���e4��gվ(?���>X�>�B?g䋿��D����D7�����>}:
?I�>�{�>����7��V�S� ���`4u��{�=��h>�*N?ʯP?�Ӄ?�ԁ�D^+���u�wH�Б�=��̾�`H>���=N4>��m�?A���#��FR�Vhi�!C��AW��#=$��o�=kUT?&�H>z:?]��?�#j>��Î�B�Ѿ���c^m>���>ES{?H��>�+x>tG|�=+����>Ҭe??Uԫ>8�¾��_�g����q�=���>���>k 6?�2U>5,վ VA��2�����jI8��><�T?p���1w��d�">�$L?p��=C4>�>�ԃ�����������>E/?g->�,[>桾����_��5!�8�6?k�?��V�.� ���>��,?aw�>L�>+Ą?~J�>~�����=[�?�9^?�K?�x-?�H�>,�μ��(�GɽL
;��\�=�Н>�C>��I=v�
>���K�*��týB�v=v��=z"3�#�"�爩�����<#��}eF>ʟֿ�M�X��~�?x�	 ���O����������G��;͝��	���a!������׽z������1���ս�o�?���?kG����}��*�w��̼�9��>*&ž�Z =�f����s��&r�$��H�Ѿ��,���`�̧s�j�Q�'?Ǒ�O�ǿY����=ܾ	 ?�K ?��y?^!��"��8��R >^"�<W���S��I�����ο㯚���^?���>��~�����>���>��X>�q>:'��l➾���<1�?��-?��>��r��ɿ^����z�<���?��@<B?�G&�ѿ��s0=�~�>3e	?
�9>47��R������0�>�ƞ?�V�?�\^=SV�?���d?�< �D��������=�գ=b]=<���D>�ԏ>����j4���˽18>TL�>{�yF��a�vߺ<4�Y>Ӫ��ҡ�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=t6�艤�{���&V�}��=[��>c�>,������O��I��U��=̓����ÿC�$�����D���l�kT���0�����]d����� ⃾l�k�c�<̜=��3>>�n>11>_?�>��[?�3|?Қ�>�y�=�O��⟾rz���Ƨ�����j��G�c��D���L_�֧۾YS�w����'��&��q���.=��@�=/R������� ���b��>F�C�.?��#>�vʾ֒M���<Zʾ,���^����G��fx̾B�1� �m����?��A?腿� W������r��?�W?f��Ū��۬�e�=H����=�3�>�P�=���"3��S��*?h�!?����F�j�d�=�Ѝ��E8= H?��?Un��ҏ�>��=?�+�;Q�#=��>�
>�>ޕ�>���=�����Y㽬�?�S?��=���U��>��v����]�>h�>V��j:��*�x>�;�=X�"��	�=�r���Y9�`2W?�͍>T�)�� ��b����0�;=E�x?��?[>�>�{k?I�B?\ҧ<�8��*�S���w=�W?-i?��>�.��� о�k����5?�}e?eN>8Sh��o龘�.��<�(?,�n?�\?�8��,g}�A�����\K6?�p`?B4����e��򉾤�?;.?���=W�}��)?H�><ľ�����̿��h�ͭ�?7�@���?x�=�,�<�K�<��>ǳ?��}�v:c�,�7> ����K�>|��"�_���ʾ�h?�>�?̢�>��~�y��#��=�╾�Z�?��?�E���m<)*��k�#m��*כ<�Y�= ��$�Z����7��$Ǿ̼
�Q����0ü�߆>@@����>�h;��@�	Ͽ򅿈jо�)p��f?�٩>��˽ ���<�j�pXu�|�G���H��{��a]�>0>�������8�{��h;��_��1��>oN����>�S�����k����:<��>���>���>_����Խ�ܻ�?�2���9ο⥞�ȏ��X?DV�?�m�?%v?��8<��v��m{�����(G?ws?�Z?��%��[]�'�8���j?�\���T`�
�4�HE�U>�!3?'@�>��-�,�|=�>\��>Uk>�"/�̍Ŀ ٶ��������?���?�n�-��>���?@s+?�i�8���\���*�ԙ#��=A?�2>?���/�!�X/=�Ӓ�E�
?c}0?�~�/�`�_?�a�H�p���-�z�ƽ�ۡ>��0�f\�uN�����Xe�	���@y����?J^�?e�?ҵ�� #�j6%?!�>T����8Ǿ��<���>�(�>�)N>�H_���u>����:��h	>���?�~�?Ij?���������U>�}?P��>�?}!�=�"�>�X�=�����Y(���#>���=|�=�L�?$�M?��>��=΀7���.�]"F�+R��.�-�C�g��>��a?�}L?b>������1��� ���̽1M0�z��G�@�TC.�M�߽�c5>w�=>J(>MFE���ҾJv?���ؿk��Z�{�̃)?�j�>�)�>̞����lҽr/?AE>���������U���Ӳ?�c�?�C? �˾�f��c�>v��>�s�>P��WC
=	t�I�!>*6K?�2��٪����U���6>�&�?�@�2�?)ǅ�u? ?����i���U"	�[Ƚ�U
>�?.�a��>?2�>@Ԅ���|�%{��Z�}�>��?��?�8�>��k?��]�6�1�ثl>M�>w_?}�?��>G=�ĳ2>��?�־L���Q��g�8?��@S&@ouR?i꫿�ZԿ������Ͼ����v#>:�'>�\>�>��]?�=idϽE��=->��[>p�>��I>�Έ>Z�k>s�j>�H�>�
����+�Ы��w��>[+�1E��I��@���S�����Q����򽾨��k����aD=��p��{E=�dU>�S?s�B?+�W?���>;s¼C=>
i����>��w����=�j�>C=?��Q?��C?�a�=V_���W��ms�����I،��>@>1��>���><W>�A�56_>C�M>$�q>ܮX>f>-���y3���1>���>˅�>���>�Z:>j�>����&��9�h���v�%Iƽ���?w���?J�X� I������ŵ�=��-?*>���`3п𫭿��G?A:������4+���>K�0?�|W?��>Yﱾ�yX�8w>[
�T�k�u2>:H��Yk��')�i�P>��??qS>h�f>��3�%�8���O�P:��Ċ>�U2?���;�2��r���L��ؾ8�J>]�>_��G �u����{��kb���?=�%7?��?�ʢ�F���-n�\F����A>�R>���<�O�=x<>H؁��@���N<��+`=_�=H�]>'�?�$:>�G�=a�>�-��z�o����>nO>�2>pk<?��'?���
ܸ��]|��C(���f>h��>[�{>��>��E�::�=���>5c>�����ĉ��(�q�5�E8u>��*�#�K� ���EqW=����y8>���=�<���6���=S�~?�|��ވ����7����pD?+?V��=�G<>�"������+��G	�?z�@�l�?�	�3�V�h�?�@�?������=�q�>)ͫ>�ξ {L�T�?_-ƽ.���~�	��#�pR�?��?{}0�xɋ�Jl��/>,W%?Y�Ӿ�Z�>�e��������M�v���&=�2�>��>?)������DkN���?�K?dY��,,����ȿ˴u����>�%�?�k�?*d�0����D�ͷ�>9P�?��R?�+c>U�־>�N��!�>�j@?�.M?���>���.7��+?eT�?�f�?`�r>���?*&{?mT�>��K/x���Ŀ���5%b>�?�=�� ?-=�e/�"�:��R��P�����;���G��>�F�<-`�>��[�����=.�y��B��f͑�)�>/.�>�~>tu{>�)�>_��>}h>�=<$Yܽ�3������g?h�?��Ǿ@g�6��=�WR>X��V�>$ON?9�=I*����>vmi?�O�?{!Z?ߪm>c�	�j�����ÿ�o���.>�[�>�?^#?�>>�Q�>�����x�$h>2 :>�-<O���c��S�=�Al>ܫ?fX�>�����?�K"?(��>@ï>�F�w����)M��\�>�
�>�\?C��?��?Љվ�R0�����)��V�P�?fI>+�r?�9?5�>����y���b�~<Ƹ���}�(��?@n?^Ɲ��?,�~?�C3?p79?d�q>Z�����ƾm�s�6�{>��!?���A�LT&�	4��Y?)I?h��>��Hս��Ҽ��{���p?>\?�&?��Ra���¾}t�<��%��;P�	<]!C�-�>D>}��0�=�m>DV�=ԡm���6���g<ȼ=ـ�>;�=PU7�N���"?ta;`��^�y>R�s�\(��U�>�������a}?7� �����ͦ������|8���?��?��?��=��d��:?̺�?��>��>����-�pRL��R)>!����5���>�n>��2>O裾����(��L$��(�0��|/�w��>���>�e�>�`'?y��>g��>F����������d�L{��!D�1]4�Z���v���T6���佣&������6�>��ν�)�>��	?�L>��>��>F9Q���>-��>�M�>�?F�n>��=����9�)~���Y?Σ�����+�	�홾�I?�|[?so�>�!��g��[?�m�?T�?"��>��W��� �I�?�
	?`J�S�?Y�K@⽛Q�"�����6<���.��>�>��Ľn?�7��R�aC�>��	?]�\�xĮ�%ڮ���h���1=�e�?�B?�6�-�W��
s�&{.���@�չ����̽�H�5:��_�?ƈ� Ʌ�\bv����`J�=U<$?�?*� ����|� ��Ɏ�D[�٬�>��>ǂ�>�@?�剼��0���%�0�N������s�>�'x?�m�>�C?�t2?kS?30?�.>�v>\�]�5?,$T<�U�>�i�>8#%?(7?�DM?�?#�?��>��W�5���kӾ�'?�6?�'"?B�?���>�_Ⱦ�5��'���Ê<q�8�˂�`Ƽ��>=�#�����ɘ�;k�2>C?ȧ�J�7�c����k>��6?�O�>r��>W���ă� �<��>/4?��>R7����q�`:�@q�>4�?���w�<H�(>���=���fL��]��=�඼t��=��U���6���?<��=��=� ���O�:ڣ';�%�;���<E��>�`?�>1�>8M��7��Ȱ����=�b>=�[>"�->g�׾>苿�;����f�Dj>�L�?(��?��f=�,�=���=o}��0p��E��m3���w=�?�<?<�S?B_�?��=?Y#?�V>��6Z�����_t����?w!,?<��>���׳ʾ�񨿯�3���?G[?q<a�;���;)���¾I�ԽC�>�[/�B/~����-D�=煻���+����?ֿ�?oA�6�6��x�̿��I[���C?"�>1Y�>��>7�)�z�g�\%��1;>���>FR?�P�>�O?�-{?�Z[?q�U>�.8��	��g���\���~!>�@?m��?V�?��x?���>We>k�)��8�Z�������u��v���Q=M,Y>�b�>���>���>_��=��Ľc���C�>�3w�=`>�Y�>� �>G��>��v>F�<(�G?��>�S���� 뤾����_�=�h�u?W��?��+?{=kv��E��%���H�>�f�?d�?�.*?�xS�}��="�ռ�ܶ�O�q���>��>��>N��=�vH=��>0�>��>X���S��q8�b[M���?UF?��=�h���j�Q����ԫ���j�@�l�ĉ�;Qj̽����8"�=���-��D����<����Aգ��fݾ�p޾Q�P�r/�>Q���=g>��n=�@�=$~=s1G�ceϽ �I��W�'������m`�m�缇�$=��=�y�=�FO<Yk˾��}?�?I?��+?�C?N^y>��>�E2���>.E���I?�V>T�Q�ӄ��kz;�{��������ؾe׾_�c�����.>[�I���>� 3>���=�<�^�=��s=���=	WR���=���=�)�=�_�=���=M�>'P>@%w?_���uƝ�:�P���轆�:? �>6`�=�.ǾV@?�v=>F���������f�~?���?f�?n?u�h�� �>���������Ə=$����0>���=��2�ٹ>~BJ>���8:��ѳ�h�?��@�Z??q勿ǌϿ�(/>�/>�a�=Q}R���1���_��_�lhK��( ?��<���ɾgE�>3��=�۾�kľ�%=�c0>C�>=�"�n�Z�Qy�=����6=_�z=��>�YJ>л�=�^����=1�9=��=7�G>s�,��@������D=$t�=ˍd>��#>9��>Ռ?�D,?(Q?��>�\R�m�ʾ�qɾy�>D�=ݜ�>c�=/W>�!�>�7?;�??�F?	��>;��=��>���>�0���n�����P���T=�5g�?n�?7�>��<�
N�2���_8����?�+?޹?s��>ex	�J0������� �>��
>��G=�T��N��,���{���q=#DE>jο>���>�ɣ>*>B�>��r>>Ű>��s>�G)=]R�=k���ʵ<V�=m!�ߘ���Vk=���?�J��Y��{�U��I�V'���(�+����$<j�=lk�>5M�=a��>=�C>*��D��=Ŀ���9��}=�
�$�T���_����ť;�s4�w*�>cI>E���2��|��>��>���=�4�?�h�?Z�>��e=�؄��Ψ�ND^=��ƽ��>�G>�>����Z�XCd���Q������>��>\:�>m>�,�#F?�51u=3��65�b��>� ��Y�����$q��1��(��i��ߺ��D?7��0�=��}?b�I?�ޏ?
��>����{Xؾ�0>������=�F�p������?�'?c�>�쾣�D�!���\�����>�Д��PY��􍿥S!�}ʽ.zپ�\�>BȾ�X쾊g,������^����R�N��ik�>�`l?2ī?6G���R����P<��1��>��_?���>	�?���>ha������^��'L<w�V?g��?i-�?�6�=�`�=�����F�>>�?R#�?.(�?P�q?j>��I�>T���T/>�6�f�>��%>TB�=��=Nx?�	?�?�X����%�%񾌣\�h�+=�0�=���>���>Ehr>k��=���=+�=ޙ@>$�>� �>,_>���>{�~>$	������Q2?�*)?��2?�G�=M��=�.C��뉾�-��fP�D�7��~J��#w��r�a���5?�4���)�>��:�?�W�;}p��N�?�T"�R�,<���=�0[>�i���<?E)�=�?�>��>�TY>�s�=F˒>��=+����=.�
���E��j)�EM� >K<ʫ���+Y�Z���n������x���v���e��Du�+M!��w�>���?�6�='9}�stC��*K�f��>CC�=۩�>))k��dA=SF���?]r�>as����qÑ�2��]��?�'�?9Dc>��>x�W?͙?��1�+|3�zZ�9�u��A�C�d�ޡ`�ۍ�ϡ����
��J���_?��x?�oA?gݒ<<.z>O��?�%��ŏ��6�>�/��);��==II�>�����`���Ӿ޿þ<2�GcF>ѐo?�#�?�[?O;V�^c$>�kv>�;?��?�Ym?��1?��?#=�|G?Ԃ�=�_?M�,?$�H?�*1?��;?9>�a���$��Tcʽ����>5��0��' �p����/K=�Y�.�>�=|���s�!���(��a*��k_=�`=p��=�8>I�>��]?�D�>�}�>k]7?V�[�8�o���)#/?�>=�s��q̊�����az��>
wj?O��?xZ?e>�\A��B���>��>Gr%>��Z>J��>T��B���=�@>�I>�z�=:K����	�,ő��8�<�F>���>�B|>t����'>kz���-z���d>��Q�Eú��T���G�3�1��gv�t`�>E�K?��?��=�\�2.��qDf��+)?�X<?iGM?.�?�&�=�۾��9�'�J�2/�Q�>Թ�<���
����!��v�:�h:�s>�*��������P>�u�o�۾��t���E��̾^�1=���Ų=�n�Y>�
�R����=Q��=�����{%�7����Ч�w�B?V3�=-���5y)�����ms�=lњ>���>)��^�V��C<�O�Ҿ(�<��>"f>k<�EK���an�>Ї:?�u?M�?�^��uv`��-��ұ�� ��a!<�#?5��>%��>�g�>��>���f���q��H�:�Y��> ��>���7�9�����8��������>s��>�5�>;O�>�?�Q?�p?�I?%f?�b>���������?7?��?���=�I��w�Z�tl
��a=?)�0?`&���g>CC?�?~4?L&d??]�<Ά���F�։�>rr�>�'�b>��'�>�mE?_8�>pjd?�Z�?<�;_%��� ��P�������6a>+�7?�?�0!?�W�>��>���1��=a-�>l�f?U�?�l?!��=�?�->`�>�l�=SH�>rY�>T?9�J? �o?�dI?f��>�0�<����ѷ���b��1;��
<���<��x=�':��s��E���.=l�<���e�����Oh���ƕ�<nN�>�	q>񪘾�,><�ɾb�����F>(ͦ����|����6�/�=��>D?���>��%�E�=W�>^��>��N(?-K?��?�Ѫ;K�a��ؾ�O���>.�@?b��=~�o��ϔ��u�,�X=s�m?ؼ[?��_�/u����b?h�]?�N�2=�J�þP�b��龬�O?�
?��G��>��~?��q?���>T�e�74n����REb���j�f�=���>�f���d�*"�>~�7?�j�>�3c>.�=�q۾��w�����U?,�?+�?��?}'*>��n�b0࿄a���͑���\?Ws�>�v����!?�џ��Tξh;���׋��Tᾁ����+��+#��uF��x&�� ���e۽�ۮ=]v?�s?��p?I�_?���nd�H�\�q �8�U����m��F��E�jC�1n� 	�I���ݜ�%�>=��S�e�B��"�?X��>p[Լl��>��~�%Ѿ��ྈ6u>*��;I�z�,<^��5����=���3���)
�w�?
�>X|�>shG?�u�H�N�H�.�Τ'�l�
�v>�>Y�>"�>C�:�B��@�����
T׾�h�;�7�>ȇ\?��j?�o�?��{�����z����$e=q�ʾ_p<>|9�>�G>�L�˼˽k�=���Q�y4\�����Pz��BC���:��$?��&>5��>�?�)?^z���ݾ�F����B�f�=Y?��?K��>��>��_��9A�ؿ�>��k?pA?}��>ה��G�#�`��j�\��Z�>�1�>�i/?k�>������Y������Ό�F�L�`��=Es? �e��N�H�>WQ?��S=�=�=���>���C��Y�<��5Vx>�?
�j>H��>Js˾d�g_��W���4?�?�_����/��)>��?q��>T��>���?p�R>���\Zi=���>q�[?�nK?gn@?��>�x=H���Ͻ��2�񀐼�f�>*��>7z�=q��=�/6�܄���[Y�=A�=1��=P�#�����M��=���=��b>�9ʿE*J���	�T�������:T�tb���ٍ�����K�����������D���u�����(2���F�~�?�@�?�37�S��� B���Ri�y����>�����<�ux��Y��y�����龔���D�V��h��rg��'?U���	�ǿ����*ܾ ?w@ ?M�y?�� "�,�8�$Y >'��<v ���뾻�����οѓ����^?6��>���,������>���>�Y>�'q>+����ږ<-�?[�-?���>}�r�E�ɿ����&ǥ<��?�@<A?��(��?��N=x��>։	?
�?>j�0�>L��B���x�>A%�?���?'
M=��W��	��re?�<��G�ǂɻ���=an�=�L=����ZH>i�>DD�3B��ؽ,�4>\߅>�_�6&��^���<ޥ[>\�ڽ�R��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=.*��_Ŀ�U8�����z&��ּ�7��]
���aȽQ���Ŝ����:��=�>�4>��c>`�@>��j>>Y?�"�?e��>�v'=��Q��n��f.���떽Ss�Z .���^��1��/u��5侯��c�����]�ឹ�c=�'ލ=�:R�����i� ���b�s�F�p�.?�M$>��ʾ�M��
+<Iʾ�����ʄ���7̾Ŕ1�Sn�|ǟ?[ B?�셿��V����h�����n�W?���U���߬�A��=�����Q=�>���=O�⾱$3���S���E?zK9?}Vپ�h����>U�G�UW�=+O`?�?�,����>�D%?~�,=��=*o�>��n>���>B]�>!{}>������7��t+?��O?�y�=v�G�W�Q>�3�������0>șo>����E�>B�>�k�=�1��j�i�;C��v]���W?�ߐ>)*�����A���*���G=�Yz?��?9��>8�j?�B?�ߋ<L�WqQ��K	���t=�W?��h?�#>����6�Ѿ\���7?Ede?�L>��i��b�x.�O(�w1?&=p?}~?��Ҽ�d|�z\��u��I�6?�fj?�*�8���䑾7'~��N�>*�1?�P2>�O�����>vV.?����� ��A¿U�W��δ?��@�@3�w=��W<���<�M ?d�>��������r7>C���ֶ��=?���/����U��l�]?J��?��>ܺ¾�����=�u��?��? z?�������O9��"]�%�����=��=4��;zJ��df꾠�?�.Pվ����2����ӽ.ۀ>�E@c��>i���y6޿Ɔҿ�큿W]���L����+?6�>��پ?�e���z��3N�@�J�";/�딼>��X>@e�yCE�ޙ��Y�Q�p��<�?��ü.�>�%�����Ar����=�O�>q��>H�,>��	`۾���?Z����wտb���L�"O7?^W�?~)�?��?�6�&I��R㜾�䘽��<?=ن?Ȟe?������Ž"C���j?�J��^[`�-�4��@E�R4U>q3?�#�>��-���}=�>�W�>�V>G /��Ŀ�׶�����=�?2��?G[꾌��>)x�?u+?�a�t5���N��m�*�RRI�u+A?2W2>����A�!��1=��^�
?�0?�<��B�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?]>�>��?.��=l��>d@�=U����+�MV#>H8�=��A���?>�M?@�>�`�=�7�T/�OSF�qAR����C����>!�a?-gL?�a>⎸�V21�4� ��ͽ�1�����?�\�.�*�޽u5>��=>>��E�67Ӿ&�?�o�]eѿ[����z ��9?ڙ�>�>�>n��N.Z;� ��<?��o>�y
�i���0��&�Ae�?���?�P	?�t��W����!�=���>��y>�9�G2�s���=3�Y?�b�����y-k�4ZX=�a�?��
@b0�?�Cv�?%�־	���R�o�7u쾸 �d>�?F���Ś>p��>�I��y�v�����S����̡>�b�?�?���>��\?��^�f5�}�f>�3�>&_@?z�?G/T��v�Q�>b?,��O����3��)??��@Q@ZXI?�ҥ�*|׿I���⫾2��r�;Up=���=B���o�:����<�qk��`=Z��>��>	��>�^%>��=D�>\����%�a����j���J�pd5��]��R���;�Ծ�Z�1*ɾE̞��1=�RW=D�.�ħh��p�۠����=�U?}�R?Oq?��?�u?��>������=��.����=���>Y�1?R;L?�,??F�=BF��ǅd��D������������>��G>L1�>Z��>���>PK;��K>�>>#
~>�r�==^=����_=�\M>�	�>9��>:��>�H<>ǘ>Cδ��1���h�hw�̽��?{��z�J��0��u7������]s�=�b.?�>=���=пT���p1H?�����*���+���>�0?�`W?��>t�� �T�=>@��f�j�"Z>3 �b}l��)�x&Q>�l?o>�,>�6�A{��#T��þvv�>,W?�6�o�m��\���t�F���,'>^d�>D0<��,��.��������\��<�/?
?h�>z���Spb��Ӱ��a�>1�<>�%�uJ���x�=�.轆�u��pý`>d�<c�=�W?��+>�T�=�̣>�^���YP���>�B>�#,>�
@?�#%?~��%+��9`����-��w>|>�>��>+H>@eJ����=K��>�a>M�i������@�T@W>��}�nW_��au���x=�헽��=��=�� �:9=�M%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ&��>�q��񙿌r���e���Z=[:�>)�,?(����=�(��y��>�Q�>�H徝Q��HvƿN�m�c{�>���?(4�?��Q��~��l�I���>���?�	I?��@>J�ھ��!�Ŗ�>X�:?�\D?�k�>�,�Y�J��?O{�?D��?۩�>�V�?#i~?_��>��h�8�S� kٿo����+�>��r>�N+?�C>�V/�5�k�K⏿�ʄ�i�h�1?���>Љ�=7C�>�ф���&�x�=�ï�bqm��'��!�>�>#�>��>���>���>��>.[�=\]�׽;���'��L?ջ�?����Fn��7�<�˚=!�]���?y}4?/~e���Ͼ�>�h\?t��?�[?7��>������k¿�KO��!��<akJ>��>���>����J>�վ�C�=�>���>����aھ$I����û��>�q!? ��>ꬰ=�� ?��#?�8k>s#�>7KE��6���6F�B�>=��>uS?*?z�?y0��v3����g᡿��[��	N>e�x?sF?]ڕ>z���a����C��H��A��6{�?�]g?�佺?�!�?d^??ΊA?Dgf>xU��ؾ(��)�>X�!?,���A��4&�B���M?(Z?a��>�ᓽ��Խ�3׼��0��?�?�[?�&&?����.a�$9þr��<U�!���I���<�7�З>t>��Y�=��>?��= �m�c~6�b�b<0ֺ=�}�>�v�=_\7�qɎ�_P(?��=�����;>�y�C`-���>1�v��J�L΄?#pؾ�~�[���k_��iŞ�p3�?���?��?P{�>�Gf���/?��?%$�>x�?�� ��&?��%�Ņ>�����>�PpI=ae_>���< 烾�ͧ�����Q��Q�-�3��>��>��>p?�P�>���>Y⏾��[����Kl��A+���T���.� n��Q���O���Q�ۑ��a_�����>t���d�>��$?О>�RU>�y�>���,|>���>��>i��>�*>!�>�B	>���<죁�qIR?����a�'�ʶ辪���/B?�pd?�1�>i$i�d���0��}?���?Ir�?�?v>|h�R,+��k?X:�>����p
?��:=�{��s�<�N��Y��GO���U�P��>k2׽� :��M��mf��i
?!.?͗����̾
b׽��u���=z��?�?^�%��Q���_�G��j1����m.���QM�]7�ڐu�a�����6s�)�'�Vrf�k`?�?�q�:�¾9+��5n��yt���=�?E�s>�Z?|��=U�(���X��E�!� �dᢾ^��>06y?�S�>��O?I�+?]P:?	�[?�/�>�M�>��b�>C2�q��>:�?�pR?6gG?C�Q?�?��?X�>�%g����v�龗PI?��"?(�3?�D6?�/�>K���W2�@x�+3==U��S�����89>�}���;�Q� �̴�=^Y?����8������k>�7?~��>���>y���-���!�<�>�
?II�>*���"|r�b�4V�>��?���=��)>���=/i��T�Ѻ%]�=����N�=�3��Xq;�zY<\��=���=\�u�X������:Ç;��<�t�>��?۔�>�B�>5?��� �c���d�=�Y>2S>>�Dپ�}��u$����g��\y>�w�?�z�?6�f=��=̖�=d|��NT���������'��<��?�I#?BXT?)��?'�=?5j#?��>�*�.M���^�����̮?k,?By�>���R�ʾt�9�3�G�?�M?�Ca��d��+)���¾u�Խ�>S/�4~����D�E������^��8��?���?X�?���6��f�ʻ���T��~�C?���>���>3��>X�)���g��#;>Q�>W�Q?Y(�>��O?�C{?1�[?�qT>�{8�a!��ə�̞1���!>�@?8��?�ߎ?;y?Sv�>@K>q*�i0�RH��|���m�ꂾF�V=�|Y>Jj�>:�>���>��=×ǽ߲����>����=��b>���>��>��>�v>D��<��T?��	?|þ+� ��X�Kj��N�<�~�?���?P�?��N==���C�Xb���b�>���?�Ӗ?��?�HA����=v��I_�J,F����>���>dh\>Y�_�/_T=B�Y=�K�>���>
���`E���m���?02A?lJ>�>���e�~Ε��Z��=�����aͽ=�f�B�>O�о�X��	�y��'F�����������)˾_t��ˑ�>���=<�=4�=@�#=�����<�J|=�
U<�������P�=���)Q�<�0�������{=��=��>E�ʾA}?v}I?�C,?5�C?0�z>>~�7��?�>In����?�6V>0�R��û��9�
����Օ��Yپu�׾g�c�B3��s�>:|J�h.>>1>Pl�=�<�<���=)cx=��=�fn��1=[I�=瑻=��=�H�=�G>{->�5w?c���߲���*Q�]��V�:?nO�>`�=k�ƾy!@?�>>2������Vl�6"?���?GW�?/�?�Bi�E^�>B�����:]�=�㜽�2>��=��2����>:�J>����G��>p���.�?�@e�??!ዿ��Ͽ|/>*�1>;��=ѳR���.�ѢZ���e�P R�&�?��:��xž��>��=�ھ�Dž�!=�6>�L=	r#���]�S��=��~���/=��y=�]�>�A>Aθ=���)2�=��5=���=�EN>�F��@/7���b�' =��=�[a>�}.>��>��?�d0?J]d?��>	^n�?Ͼl��uC�>+X�=YJ�>x̅=s�B>���>g�7?�D? �K?�_�>#N�=��>4+�>�,�|�m���
⧾��<���?�Ɔ?���>,�M<��A����BS>��#Ľn�?�J1?)u? Ğ>�O��v㿠7���e����9�=2���.0�<��������W�����>�W�>E��>�]q>*&�=K�)���=k��>���<�R]�/O�>d�޼*�T=���<䛡=�9��j�j>v�;����+�=�ɼ�0����1���v<���=e�=d��=���>��>.��>ɖ->]U��S�=;��S�<�~�m=��ؾ��J�T�o�&݌��1��'��R}>f`>b��<8Q���r�>��>���=�p�?*�~?-�'>��=6i��ű��)���B����=�5>��#�j���lN�Ğ���o�>��>�X�>:$l>�Q,�?��{=��Ὰ�5��K�>.*��tH"�=���p�5���۟�>%i�{�(��3D?~"�����=�4~?�I?�̏?��>�T��%�ؾ�/>u��m.=����r��a��#�?�!'?V�>���E�M�˾ى����>��I�N�O�a���1T0�*�/�DH���5�>����XEѾw�2��A��������B�_r�F�>�P?fݮ?7�`�@H��_wO�m��`ށ��3?Hg?׼�>�J?�G?£���N�����u�=\n?r��?y�?��>�!�=�񴽲`�>/@	?��?M��?7gs?ь?�x�>w};�� >�Ɨ���=��>U2�=�[�=�P?vq
?�
?O��%�	���]���:^����<�L�=���>IG�>��r>|�=��g=�T�=�u\>
��>�Ϗ>t�d>���>�!�>-F��S�����<?Wj��|�>��<?\:�>��#=^����_�
�:4�yd��zS��s}�Ǵ����=�m">�ҥ����>=�οu��?�$�<ax¾^�>�I�b۬<�\>��>�=2�@I7?v��>��?��F>���>��r>̼�>����?�ľ��=�����*�*�O�."����>�翾u�,�Z$�����������E����c�8Vm�w$B��5�=܃�?��Y���g�@r=�E����?�Ă>�3?V���. =ގ>2?�:>�Tؾ_��������*ľ;��?#��?�;c>��>D�W?��?B�1��3��uZ��u�^(A�<e�T�`�፿����
�a���_?��x?yA?,O�<3:z>'��?��%��ӏ��)�>�/� ';�e@<=u+�>�)����`���Ӿt�þ&7�oHF>��o?A%�?�Y?UV�5�`>�z$>$4?�7?Z��?��?}?:�= �V?�/�?iaP?��m?pL?.N?V8>x#T=�`ļ�޴�[�����X����:���)Q=�,[;���<�@����s~@=�J)�]���g��<;^�+�g���M�o�<��=���=���>��]?�I�>��>t�7?����u8�뽮��+/?J�9=o���g���Ǣ���i�>��j?f��?�cZ?�ad>��A�C�Q>�Z�>`x&>�\>�b�>U���E�k�=�N>�W>��=vKM�ρ���	��������<`(>j��>|>y��r�'>�����Ez��d>T�Q�*຾^�S�k�G���1�lQv��N�>s�K?f�?	�={t龄ϖ�;f�%)?�[<?�QM?��?u�=[�۾��9���J��1�/�>�Ѧ<� 	����� ��r�:�Tw�:�|s>E��:���8�l>�s	�s/ϾI�r���D����ӟ�<����7=S��؆ɾ�Wu�/3�=�h>þ�"�*����v����J??�J=ѩ�FB������>���>���>6	�W���"!>�
:��Mv=g��>s�Q>�Hy�U9�y�A�Mn��C�>I4E?�@?�2�?a���x�B�5�_�9��������</�?�d�>)+?v��>��M>�Q���#��L���jY��|�>|Q�>�$����a־<t ����A��>�b�>�X�=�+�>5�?��>D�]?-4;?��>��<>�ν����p!-?�_�?�u�=A����}[J�f�1��?��,?���7M�>�5�>�?�EL?g�b?�K�>ی�����sz�܀�> }�>VwF�����NB>��!?M�?=�?d�B?0y�= >��s(��U7� ����=#$?�/?��g?�F�>��>�����>���>��f?���?`2\?�C�=��?>��=���>��>{=�> ��>G�?d#H?ݟ_?;)B?e��>���<qה�(.��f��3�<���<��E�,Z�=p���Hx�X����L<O�S=TT�<����J����d��?=Y,�<��>�Gp>5��q_2>B�¾>A��x�G>�5���U���y��Lm;��L�=��>�?:G�>V�&�ퟎ=!��>3��>i���'?"?�U?��<��a��۾[^S�@�>Zz@?*�=w%l�\2����u�%UV=�nm?��^?�#Q��(��/\d?+0^?���r
-���辀�O��O���D9?	b?&�5�{��>�B{??xm??�>V��2k��F��g(b�Ffp�"�>W֑>/���S���>Q�8?�ܧ>�7>��>������r���r���>�9�?Q��?��?E�>��b���ݿ!����M��	K?mc�>�`����?��=K�ƾ�ԡ�q�v�Y�����r���c9y�nP���H�0���*Է��3*>�?p?��m?��U?
�߾�bZ��LY��Ã�6oQ�`2����qF���J��nG��mn�3L��*;��a�>��=�,m���7�	�?�+*?� +��F�>�l��F���5���`i>�p��zG9����=A����M���t�����G���X?���>���>��D?1Kf��J����7B���Ij>Ld�>�أ>4��>X<�<?J�����|	ܾ+g������Mݐ>!Mb?�cA?)�p?�#���#�ui���2�V��<@嶾J;L>FL>S�>��1���ӽ�y"�ŽA���v�N�ۅ��n� ~�=}d*?��>6q�>��?���>����o���3�q��S%�����]�>_2^?��>j)p>���d���7�>3l?��>f��>�M��e���{���ݽ��>��>�X ?��v>��0�w[����v����9�0�=��e?�����V��N�>9�O?n�n�;N�>/Z�f��]��K���	>g?1�=V^3>��þ.��'�{�n��,q*?�?P4��s{'�K2e>t�? �>�@�>�?��>�����j<�?�
]?�oI?��;?���>R�5=�u��[�ʽ��.�K^�<Zi�>f>� �=?�=�����|�� �÷x=�;�=2.ټR_��>�����1�e��<�

=}�M>�	ؿK�O�;�辷���ܾm1������w�D�����������7mq��P���3�#_�^�W�����Ɂ�Y��?�l�?�m¾S�z����'���۾0W�>:��z�3��ҋ��n�*���A���u��v5'��V�Wf[���8��K ?�엾f�ǿ����־A�?7�!?@�}?������6��>p��<;!>�Ě�l�̿����rE`?�;�>��;��"�>>x�>q�9>��>n���s�=�) ?�'?�a�>�g�Nǿ����;��?�o@>wA?��(��;�Z=5��>��	?�7?>z�1�����K���"�>59�?J�?��M=]�W�9�
��-e?��<�F�:ݻSj�=#�=�s=���3JJ>eI�>�`��UA�l۽=�4>-�><�#�����^��<�+]>#ֽr��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�z ��Pſ\G#���'��d=��<�jU��T�����k�m����ӱz�ۛܽ^�=~��=�E>���>k�A>0{>.X?�6l?�L�>�>fx�����?��uؚ<~h��?��Df�k��<u���8Ⱦ	��X������A�����a=�1�='R�_���� ���b�W�F���.?�$>s�ʾ��M�0l(<Ӂʾۭ���Ɇ�w��m�˾v1�Fn�(ğ?��A?������V���������|�W?�������̬�&F�=���@=&�>��=�����2�>1S��$6?��5?���/`w�*��<dZ�$2|>��D? ü>��;>��?�?�#��1-3=1��>�cN=Ҽh>�Y�>���=~���#���?}�V?�K������~�>bP���V���!�=���=����gL�=�>��̽����m�=P�&a�=2aW?��>#(��P������A��v�=9z??6�>�wo?��A?ӂ=��꾧2L������S=e1U?�,b?��>����E\վ����5?�$g?�	_>�@a������/&�w����W?�i?xd?����.}�M����J�JF:?��V?r��b˿p&�64�~��7�c?h�?�k����?��7?݀��ꡱ�㸼��n���M�?��@���?�@>�<L�=gL?��.?�k���ξ���=�Q��V�=�C�>F,��4�r�uپ� ��8IB?��?ߏ�>k[��Fh����=+᏾�R�?7��?�Ѳ����<����%m�o@�M�=��=���b3�r��i>��پZ�
������� �rH�>� @�ݽn��>����C��DM���?��!L־h�7�7#?ߙ�>�����k��{zd�ӡm��I�/ U��q�0��>>���%���)}��:��V¼��>Ñ𼐿�>�UQ�o�������6<i+�>�h�>�m�>��������p��?;���ο�Ý���O�X?$P�?�?x�?J�2;qx��s�^m��VG?��t?��Y? C+�V[���N��j?�_��{U`�Î4�:HE��U>#3?�B�>q�-�Ӵ|=8>��>�f>x#/�d�Ŀ�ٶ�)���?��?��?�o���>e��?\s+?Ui��7���[����*���+��<A?(2>6���W�!�N0=��Ғ���
?n~0? z�#.�]�_?*�a�L�p���-�{�ƽ�ۡ>�0��e\�N�����Xe����@y����?M^�?h�?յ�� #�f6%?�>c����8Ǿ��<���>�(�>*N>\H_���u>����:�i	>���?�~�?Pj?���� ����U>	�}?Ü?��?�1�=
?�{m���+��}���[��}�>=�N���#?c�d?|��>H�5>���/�9���X�%yh�����1��[2>�/?�?�ٟ>��������2^����ػ^���!�Zp'�nv�>"�=���>F~>Pw�=�������??��!��lտMˑ�6yݽu� ?�Y�>u8�>�i�8�P��*x��*H?��g>[��μ��S7��u���(�?�)�?% 
?,j���:���=sQ�>�Ҁ>�b�b���7d��fb>-�2?����e����x�(;D>?��?'�@�F�?0$\��,�>�о�헿`ו�h^���㬾3�.>�/?�$�Y�>m*X>���b����ᨿ+���|�>Y��?{�?;?�j?��*�Q�b����<�g>� ?�?Jzf>�a��wF>��,?$�Ծ���n��_?�V@e:
@�S?#1��ǚڿ>Ǥ�� ��9*ؾ�x�=��к>�+���4�=���=��K������=���>��D>O�>�a>��+>>�u>ks��/�0����敞��5�BD ��߾�qa��_4��:������T��Y���d=����hS]��@}�-2������[@>a�V?��_?G�c?�z ?�r<�뻊k�3 >��{f�=i��>%.0?~s-?�?�@y�3N��h�a�<C��(���[?���4�>Z��=�m�>���>6��>T��<DH>u3$=��>(���s���"�y����=ed�>L��>Ng�>�6<>߅>6ϴ��1���h��w�p̽��?ʆ��`�J�0��:��ߣ��<��=6_.?�l>���3<п󭿈3H?Q���++�˭+���>d�0?�dW?��>����T��5>U��8�j��d>=4 ��l���)��$Q>Sq?W�f>�u>N�3�~�7�H�P����F/>5k6?X\��V�6��Ou�7�H�ğܾ$�N>��>X\��8������M~�_i�b*y=�:?5�?I8��tt��&�u�����4R>�\>x=/G�=��L>��f�&�ɽc�F���/=r�=�O_>�?yC�>U#=�h�>i���B���Z?7d�>R:�=1OU?!(3?*K�W�{=WQ�����b>�g�>ˏ>��=�Hu��8=�o?��>��>e��`M���j��|
�>~���ZM��k�;�>�,0����<T�[>�p�Ն�� �;�~?���䈿��pd���lD?E+? �=B�F<��"�@ ��tH��D�?m�@m�?��	�ۢV�=�?�@�? ��}��=}�>׫>�ξ�L�ֱ?�Ž.Ǣ�Ô	�P)#�dS�?��?��/�^ʋ�;l�N6>�^%?�Ӿ�E�>��[�����u��"=-��>}3H?Qw��a�N�R0>��_
?�?71򾩤����ȿsv����>�?�?:�m�r7��+@���>��?�XY?�i>xj۾�VZ�Lj�>��@?$�Q? ��>�?��'���?�ݶ?���?�4�>�7�?�	d?D��>I����� ��1�����.��=D�>�9j�>G>}�ž��A����"9���Zl����?>�1�<��>�<ӽ����T��=X��hi���c �f��>'r>;��>Ɵ>d��>���>K�>�x�<_S�� p����e���L?�|�?f9��WW��Ԅ��t�<O�4��{?{/?k����q�>l]W?�{?��[?NN�>������!Ի��I���:<��>t��>=1�>�<��5U>��ľ?�����>�F�>i�0=!��������8�Z��>��?P��>�U:>.q?�C!?!��>���>n�j�e����D��%3>���>M�??|Zs?�U�>�ad���>��摿!���U��N�=:#j?��=?���>ڧ���4��\*W�f���$�m[?�@I?�4j���?��?��:?��p?�>�>w�|�C?ݾ� F�>�3"?C���2A��?%���M�?��?R$�>����˽����:�UO��?%?��[?�s$?څ�*�_�(\¾rm�<rUA������9<F)��n>��>V���Z��=*z>�^�=̟n���7��8�<%��=��>�=��8�f����?�8�=�x�� w���S}�ygc�`�>�eN=+���si?��BȈ��������*��9�?&3�?U��?�Q>\�p�$?<<�?��w>'?Ǻ�=��4��Ҿf1�=1l ����Uħ>T�>YD�=L�U�ʢ��?����臿~E-��.���>��>� �>��?O��=S$�=��9��� ��0�*>��fx��@�{�P�4�n����8�sE��1廋��4�|����>��<Ԍ>�s*?���=�.�>�?r�>�>Uw�=���>�
�> �b>�9ݻ�p-<a�;=E���sLR?���x�'�B��+����,B?�Zd?�>�Wh�{���+���?���?sl�?Gv>�{h��.+��\?�&�>s���g
?�):=����[�<O��d���^��t����>�D׽:�_M��_f�[e
?�*?7)��݋̾�F׽�枾y�q="�?(�)?�*���P��ap���X��2P��4��<�e����L(#�r�������踃�V(��6=-�*?�.�?���a��Am�o�:�o�]>���>Z��>H�>WR>^���s-�5�[���%�Nr��Ҝ�>vz?/�>��>?�=?�cY?�M?;��>!��>t�����>g(>=k��>�>�`>?n�)?�*?�?�i?|2>�̽/�쾾�����#?߹?�j(?�2?ն�>�����uG�L^Խ-	��V/��*==�[=.����'�4�n�;��=��?����7������a>˙5?���>O��>�i���u���.=}T�>
?uY�>����v4r��
���>9y�?*P����<W(>Ȟ�=ҥo��5v��+�=ϳ��
�=#ZM��D��m�:Ԙ�=[%�=��7��u���r�;��?��<K��>�?��>�v7>W��Hީ���C�2�m>��w>�'>��\��n]��Or���Lm�2��=�R{?E7�?�u={�=aS�=v���g�҆%�U~��0˼qWt>��K?��o?!��?��%?_�Y?c=	���Ǉ������=��u?��+?{��>�9��_ʾC�����3���?�?�ea�5]�-D)�U�¾ԽxX>�H/�w/~��ӯ�G�C��ݺ*}�q?��cp�?�Ý?�p9�h�6�k�~ۘ��>���:C?�B�>�Z�>|��>]�)���g�Y��]�;>���>eR?e�>ERR?/p?_?��D>��$�6"��r���.�k=^,�=�/<?"Ѓ?`Ë?�vn?GU�>g�>��l�H����9�A�����0���=��D>�U�>�i�>�G�>P�=YJ�h�����M�Y=>�q>��>a�>�6�>�(2>�|����H?{��>�c��5��<��	���<ؼ�x??�?	�(?�e�=��&�<���X�>(�?gf�?�#'?�[g���=�z��C��˜�z�>Lv�>
�>�7�=[*7��(>���>Q��>� �T��19�w�p�a ?2�I?��>����l�~�a
Ǿ�.˾)	�<����ۼ�>���~^A> �����r������G�������ľ]о�N������$�?HM=K�=�݈>�d)>�� �v=}�˽�]����=�����w�\"���<jsB�)g���
U=>��=Qc����p?,�[?��2?[V?��>���=�ѽ�v�>_�1��?.�D>��󍶾6��M���4���V徴����K�Iз���R=�a�i2>�2>M>��:���=��>	V>Ʌ�l�<U��=r�1>A?=kd�=I��=��N>�6w?W�������4Q��Z罟�:?�8�>^{�=��ƾr@?z�>>�2������}b��-?���?�T�?A�?5ti��d�>H��[㎽�q�=W����=2>Y��=~�2�]��>��J>���K��J����4�?��@��??�ዿ΢ϿEa/>g>>��>��P��p/��N`��ae�9*[���!?
9���˾;��>���=�n޾"�žN.3=�2>`�T=A��.�Z��)�=H"���{ =�s=���>��I>b��=������=�=j=��=ŖM>VY����+���4�F��<uK�=��b>�/>pg�>�O?�A1?'Zd?k̾>�t\��|Ͼ3'ľ���>���=�D�>���="aH>���>�6?��B?)�H?ږ�>��= �>ߑ�>ͥ,�X\n�R��l����'�<r[�?��?뗾>aX�<�<>��<��R=��軽qZ?4�0?&<?��>�h��X�it��B ��.U`��7<���;S70�17��*=�c�~�q\��M�u��ko>���>�>�j=�]��ˏ=u��>K��>)�p[���i����8=k���c�=U2=of�<2���v=�?=��
��r�<S>}�3v�=⒒����?ģ=���>��>{�a>�<�=�ͯ��P�=�����I�"⽮"Ͼ��>���~�dr���9�x��o#�>�n�>������>#�N>��I>�?ͬ_?9�����=9+���E��	�$���l�d�=��8>�ވ���t��3p�ͥW�-����9�>P��>mբ>�p>
+��V?�E�=���Q�4�X�>\Ԉ������nTo��S����h�_h���C?.���Ĥ�=y?�]I?\�?���>#�ܾ�6>([��\4 =e;��m��W��H�?\�'?�*�> ����D�p�Ǿ+�a<>Ĝ���t	��U��-��o+�����/��>n�����*:��9j��t���EB�V⽴}?Ė~?��?�۠=�肿}���<#뾶𐽙Q�>�
J?���>1:�>���>�H��'�� �nD�X�v?�|�?��?\<pH'>����[p?�d?B��?�]�?i90?�m����>�X�L�>�9>h�>[��=��> S}=|��>2�>d�>SZ��3'���H�(�`%�������T�=X��>*b>M��>�A>2�'>�p=	�/>�>a��>V��>�{�>�)>�B�����IW&?G,�=q��>��1?�N�>�HX=v��nL�<��G���;�Z)�+�����۽��<Q�����L=�ɼU��>}ǿ�'�?��O>��B�?�Y���2�=	V>�rV>���@L�>�E>H8|>�J�>p$�>k�>�}�>�H)>y~�:��=�j�C
.��1�`�L�q`���t�>y����s������H��H<�"��bb ���k��oz���-����=�G�?�A����u�����j�7�>���>�g3?�#��A�q<��>ۿ�>}Y�>g;ξ������b��?�[�?��`>��>lpV?M�?��+��<6�{�Z�Fs��A��f�9a���\=������*˽��^? �x?�XA?�y�<�ly>n?�l%����%��>U�.���;���[=(.�>P����\e�V�վ�@þ��2�E>e:l?~~�?��?\WV�q�(>���"2\?j_?�Y?}|?�P�>.��G
4?(��XL�>O:?�CJ?-'?��&?��=	잼�;:�X>Y߾��.����W��:�!<ͪ�=Y��=(}=���A�\=���:�?��� 0=���=f���N��=F��=�6�=mhH>团>J�Y?��>D>*�8?-N%��/;��¡�a�)?��<X�� ��~᰾����E��=I�g?Q��?>Y?:�c>d�=���N��D>j�>_Q/>QhU>;��>^r��C�:�,!�=@��=�L�=Ru�=��/�z��r��>��
��<�>2��>��|>rˍ�8(>:h����z�o>e>ƀQ�H�����R�ΌG�L�1���u�x�>˵K?2�?9�=�F�@���-*f��	)?~t<?:M?�?��=�lܾ�:�p|J���`*�>�l�<���h������A:�gHP:�Ms>5��7Ⱦ�>��	�9��͙H�F�,�믏�|g޽����Z=lz�9���$;��=�Ҟ=�����[=��0��%t���]K?�P�=W������yM�����='?���>��u�5 �=l�B���:��~��>�
>S2��A�f�B��d�2�>.�@?�6s?��?T���ؐv���H�
��j��F2��?!�>5&?Ѭ�>��=�޾gT8��?��B�E�tA�>��>��A�u�,�r���ڍ#�����s�>y ?��X>��?ՉA?���>�Yd?�cT?6�?͏?>T/:iѾ&�0?�?؉=_�W�0����BM���g�8?!@?�����>�**?r�?�dG?��p?H#�>�c��H�E�:��>^w�>Ҥ������M�>�X?m<�>��G?��l?6N�=q��i�罰���v��<G��=5n,?�??��;?���>���>m���*��=Ǟ�>c?{0�?�o?*u�=��?/*2>���>��=M��>b��>�?WO?O�s?��J?&��>���<�J��|,���is��N��:�;CH<�y=d��-'t��U�GP�<*B�;�����`���񼑮D��������;Md�>�t>�Օ�,1>��ľQ{����@>)���!������n�9�%��=�{�>2?��>ff#�,Z�=���>�>���v.(?n�?;(?��;��b���ھ�K���>�A?�T�=��l�lw����u���g=��m?z^?�SW�}����b?�]?�e�=���þϼb��龲�O?p�
?>�G���>L�~?��q?(��>��e��9n�G���Db��j�#ٶ=<s�>VZ���d��>�>m�7?Q�>#�b>�)�=v۾�w�~o��>?~�?!�?j��?�+*>9�n�K3࿘
��Mޑ�6_?��>����$'?�μ�˾uЉ�)j�#3��"��󂘾�⨾��#�G\�� Rֽss�=��?�1u?�n?Ri\?ZF�<�c�,_��~��sR�?�����
��pH�o�D�E��{k�-	��?ﾭ���&�6=c:e��yN����?�?<5���?����O�ʾ7�Ͼ�J>v��h�ǽ�Q;�}ֽ���+Rp=�|X����G���?�2�>�R�>Ҍ-?�vo�1�3�!%@�.>6�nؾY�o>�,�>x>r�>\���� �|�R��r��A`��USܽL�i>�<^?�JO?��m?��ӽ��$�Ȩ����(��}�ʾ]�E>�>�a�>�J�M�&�`�*�R�>���v�~��Љ��s����=�'/? $l>�߲>xL�?W��>O�����������/��=à�>��\?��>�z>QC���Ӧ�>�(q?�5
?	�>jΑ�!�>�[����y=/�	?f��>�l.?h�>桃�*^�?%��;ǘ�+=��,�="�?�s�y{�2eY>�m]?[=@A<��>�`9���~��xQ/�4;>F�"?y-�>p:>��оw�
�Y�����6��!+?G ?���oY(���w>�?���>u�>Ϧ�?R!�>�z���C=}?"�^?H�K?�=?��>B�5=B+��pM̽�*�n�=���>r`>���=�z�=��*��Ki�5��q2= �=�{<�?ɽN��˧��{5=�h<=Rx=>��ڿ3 J�kaپ˝���c\	����� ʽ8������P ���%��x�q��7���-�o�T��!k�3q��j���?g��?D���������W|����4*�>Zŀ�(�V������%�ݙ�@�#����[�#	Q��Ij�U�e�GR?,Ї�ˣÿ+�������?x�?�b?g|����J.8��S�=OT�;(<�;!��F����ȿ�σ��Df? ��>���|�AT�>�Y�>�6c>�^>��7�ն��	{�=o?��)?�^?0b�( ��tx��X=���?�	@XzA?@�(�����V=w��>H�	?�?>�H1�I�����I�>>;�?���?OmM=��W�@�	��|e?H�<;�F�a�ݻ��=�P�=>B=���J>]I�>n��|NA��ܽi�4>1υ>#�"�O��>^���<�}]>��ս:;��.�? Q�6�r�[��p��';>�f?��F>5t�:��E?�T���Ͽ��[��:A?R�?�K�?�8?�����>Y辭}S?R�A?���>��$�mZn�.U�=Y�m��G>�����q�߶l=�S�>%Yk>As����Ё����x�=���i�� }�P	0��	�<g�D�jϽ�>�{8D��뽉����hL�(�D����=�(�=ӈ0>�>>~�>|�R>�PU?��k?���>���=��QX��G����޽[F��e	������ƾ��ɾ����V�������(���#��ľ(=����=�(R������� �)�b��{F��.?�$>d�ʾ�M�%�%<:ʾ-���Ӆ��ƥ��f̾H�1��n�%Ɵ?��A?�酿?�V�p���v�ื�4�W?�-�<�������=`a����=��>ԍ�=����.3�k�S�e�8?�)1?����D�Qf"=J���ͼs>�yZ?U�?p>t����>��>?�ī=F]4>�N�>I��=@-�>�z�>~��=�����?J�3?nn?�9��о+��>�R��Ʀ���l>J�=�T���6>Ϲ�>�K�v2e��2�=�r:=B���s(W?���>�)���``����IZ==��x?��?m'�>�{k?U�B?gˤ<�b����S����]w=c�W?�'i?L�>j����о?����5?ɢe?I�N>hh���#�.�~S��#?��n?�\?樝��t}�������o6?�{?G�Z��s��S>־3Hc�^�y>k?���> bs��>�[#?����� ����¿�qW�й�?
@ Y�?�$�<O��<��<5-�>�F?~���mH��i�=�����*�rE?Ů��r^���Kj��wOZ?�{�?
)�>���Tָ��J�=�����I�?��l?oy�Ԣ >��/�w�]��l�H��=I��= ���� �����3�T�˾����r��f3�H�{>��@҇ὂ��>�՝����~5ſ7����H��!_@���B?��+>�f�:z���Y��|n�Ʊ�Ɇ.��'���m�>��>����T����{�Q�;� ��ԅ�>ǘ�a��>��R�w�������N<z��>��>��>�f��0j�����?S����jο]�������bX?�z�?���?Wr?Z-<�v��z��4��NG?!�s?.Z?�.#��l[�T�6�%�j?�_��zU`��4�qHE��U>�"3?�B�>V�-���|=�>���>g>�#/�z�Ŀ�ٶ�6���[��?��?�o���>o��?ws+?�i�8���[����*���+��<A?�2>���J�!�G0=�XҒ�Ƽ
?]~0?{�j.�`�_?#�a�X�p�t�-���ƽ�ۡ>��0�{f\�QP������Xe���Ay����?J^�?s�?t��� #�6%?�>=����8Ǿ��<���>�(�>�)N>NH_�B�u>���:��h	>���?�~�?cj?���������U>��}?�r�>�j�??.�=`��>(�=#d��anQ�_(>��=��i��+?XBL?���>{��=9�y/���E��7R�WR�<B���>\�a?.9L?�^>������H�C!�50ͽA0������?����ν��4>�=>>�H�+Ҿ��?� ��)տ�����6���?�+g>+�>�%�"c�<��N��?�u1>(��	���VH��ǙĽy��?h_�?��?�~۾Y�.����>�>4>�A���Ұ���i[&>tA4?*�*�f����0�=r�?��@���?�j��?ҹ��$��v�v��'�өS�eW>��0?���Bȝ>�6�>��;Tav�����!z���i�>*��?��?��>
~i?u�m�=�>���1>�pv>3`\?;�?�������*�8>_1 ?V8	�EՊ���)�χR?�y@�m@��J?)�՚ѿ&۬�����\��A>>X�>h42>!�/��?>c=�O5=[Lp�a�?>+m�>���>v�>�6>��5>%>�?��#}#��7��6׍��m-�H&
���'�>����~[��Yﾘͷ�����:��{�q��7��\	�aȩ��>!R?~�T?��q?w�?��.�0�=���z�="IW�f��=�:�>��??�}R?"4?.n�=�垾Q�d�&�~��%��A���u��>�>5I�>8��>
�>!��:~�P>�X,>��.>�]�=�I=6k�;�r<լ6>d��>���>���>6;>�+>\������MLh�=Lw�PCǽ���?�)���BJ�7'��D󍾷���rϟ=t.?�>b���Dп+��U(H?Ǐ������+���>O0?K�W?6)>�����vP�ګ>�e	�I�l�Q�>u� ��m��;)�7Q>�4?Ov9>�_>}#1�L@��F�J���g9�>?�ξ�~ ��lt���R������U>,��>���Y�)�<ߛ�������)�[�=�!?�5�>��Ȫ��\����z-�>��o>H=�TD=A��=N���tL�/Ow�{w{=|�*>�8�>G�?��H>�=y�>&ԭ��ʕ��^�>��> %G>�26?)2)?~lk�T���8%�����`>�0�>�W�>�8�=�uO�嚒=��>Ȳ�>�<ݻ^-a���=�,r�;�I>׍Y��'�X�j�/��=��m�>�>�=*���vR�lN/=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿt_�>��nI��C��#=m�b�=x�>�B?1���>]��	)I��_?�r ?�O辚 ����ǿ�u��H�>�{�?�/�?��i�����79��-�>�V�?�[P?�oz>{�辈7@����>�S>?q�P?'T�>�a���0�[�?�q�?븈?�[@>���?$�|?��>3����&��籿��t��!�=���2؞>"��=�Ư�?.8��ҍ�Ԉ���lf����b>q)G=�7�>�W��S���?�<=��#�<�����L��>"$�>�h>���>��?/��>b"�>�;���ڌ��Xk��L?��?����n����<���=�&^�Hn?%k4?�m��>ϾhY�>5�\?B?r[?K�>.������Ŀ��Y��-:�<�K>���>3d�>�P��|K>1վ�hD����>C��>򼠼Ҵپ�e���ⶻ�3�>��!?J��>I�=��?�C$?y�n>-0�>��D��3���*G��
�>���>T�?��?%>?ü���4��Ò�Iġ�s�Z���O>	{x?;�?&M�>�펿 ���1���P�����z�?R:h?���4m?�
�?�@?�RB?�kf>/L���ھw���>ԓ!?�����A��c&���<?F�?OU�>֔���Խ�ܼ�T�����?N�[?�&?����Ya���þ���<���Ns�.��;RE��]>��>G��,��=�v>린=h~m�|E7�A�l<�޺= �>Ry�=Aa6��<��a�.?^�2<[6����]>�{���!)�:X�>��;�������j?�h׾�,��f���{i�������?���?2�?&��=��p���B?\�?�H�>`�?�8þ�K	X�5Ԋ� � �����/>G�>�x�;����6�����o��>b�(�=��>TK�>w�?�R?A�>�Y�>����[�ڪ���pQL���z�@��E��������{�Q9n����gԐ��e�>������>��?�[*>��.>8՛>(p���c�>|�>�ץ>Jp�>�#>T"$>��>������?��KR?>�����'����`����1B?�qd?�2�>Ui�牅������?���?js�?�=v>m~h��++��n?�=�>U���p
?_:=;��;�<V��p��Q6�����>GB׽� :��M��lf�%j
?Z/?��X�̾9<׽�ݜ���x=�6�?�%%?�4&�ɞJ�[�s�68W�iP�c���rT��}����(��q��!��낃��5`&�P��<�(?J��?h���6Z����@q�@<�o�Z>��>y��>�1�>gs1>���0��L\�h&%���j�`�>�=v?M�>��A?�@7?c h?J"*?q"�=Q�>e�a�Ȝ?5�|�>_�?xV? �K?�9B?<�?~�?��1>[��ﾼ��B1#?���>�8?k�2?��>��e�Q���?�գ9=~ꅺ��<0]����>�e���6���$�V >B[?t���8�-���q�j>iy7?ր�>��>� ��.7�����<}�>��
?EO�>a���Hwr�N^��S�>���?���W=�)>i��=�M���?κPx�=�¼;��=ks�;���<Z�=��=A�y�@��5�:�;hۯ<���>�/?��>�v/>����"��kx-��}�=X�'>ⅈ>�A�>��侨P��v+��A�g��C�=\t�?���?����j�=0�>�6�������־�K޾n}ݻ*?��;?r{?'�?29?�?;�I�Ѷ�9.���퇿n����*?v!,?��>�����ʾ��ۉ3�ޝ?m[?�<a����;)�Ր¾��Խ��>�[/�c/~����6D�s���b��3��?쿝?2A�R�6��x�ٿ���[��v�C?"�>Y�>��>M�)�u�g�n%��1;>��>fR?M�>@�G?�|?�f?��>����]��kA��̘
>i���4�F?��?���?��?�?�g.>)cK���f��ȇ=�aT ��)��5��@�a>ɽ�>�'�>+�>�E>4�	�Y����F�k��=��e>�յ>�`{>H�>wW0>84����G?k��> X��ȓ��뤾̃�V�<�x�u?<��?�z+?=-k���E�)��<W�>�f�?W�?�-*?j�S�a��=3�ּ!趾
�q��)�>��>j6�>ˆ�=�"F=?�>� �>!��>����c��p8�M�c?�F?��=�eĿ��n�znt�pA���}@<�*��ZV�`_��~�b��p�=:���ƈ"��z���U��������/���BK������V ?�1�=�?�=B�=��<^�мъ =\�;=�2<�d8=&ń�������܆�����q�����<l�/=W�\��@?u?��O?_.?,�;?BJ�>�=b����Ɛ>^e%��]?�UH>���:����!I����e����'��Rо��P�!Ꜿo)+>+:�����=�2>o~�=[L���x�=��Z=���<���z�=��'>N͔=tp�=�h�=QS�=�j>�}?t�x��Ħ������y��6?EK�>X}������k?�Y�=N���oꭿ��-�p c?��@��?m�?9�o�$ۉ>W�U�����&3>7[���_�>�)>�H��E�?!�e>�4;����2�����?J�
@�I?����Jɿ�â>DW3>�>�+R��H2�S�\���d�^�J���?d�;��Ⱦbc�>��=8��\�þ�c'=��2>�*9=�%�A�]�$f�=E�p�m�)=<�R=���>{a@>	�=���4��=\~Y=��=۾J>+�e��(���C�B�=]\�=�f>!�)>��>G=?<1?�Cc?w�> �m�V�Ѿ�A�����>�
�=�̲>�x|=�,8>�&�>�6?h:C?.CL?���>?f~=P�>�8�>C+�Z�l���wn��R2�<�C�?x�?�t�>6N<U)E������=�4�ǽ�.?n�1?�	?���>?�����ɬ���\�����{e>�-�=V��^�=���K�:��<;���>�D�>��>4��>W�G>��>�$]>Q�>�:]>	�u�`�Ͻ�r�&rG�w<.=b5�=�G	���H#:��5=��S>&��ּ l=+-���-����;���=��>�	�=��>�·=�����W>�I����9���< ��4!A��]��������� ��C�?>�9k>��c�������>�ȓ>���=ү�?�It?j=��켃�ھȪ�\�M�u�����=Y�=zQ���ML��~V���L�D���[��>cߎ>C�>һl>�,�A#?�n�w=��>b5�H�>~|��w��)��9q�@������Ui�rҺѠD?�F�����=i"~?�I?S�?��>����ؾ�:0>�H����=Y�C*q��h����?'?��>�쾕�D��̾x�����>\4I�p�O�?���F�0�:�!��ҷ�ަ�>������о�U3�d��b���p�B�~q���>$jO?Ӯ?j�`��7���$O�����戽�r?Ycg?[��>I;?�6?C������x��=��n?m��?{6�?�>���=������>		?��?��??�r?^�B���>�e�g�>յ�����=9�>��=��=q6?�	
?d	?Iݜ��
�/��3�(�V��=��=�=�>�(�>�ds>i��=I"�=4�=`[a>j��>��>��d>Ŋ�>d�>�(�������?���=>�6?0�V?�)D>��S��1���꽾i����Q=��:����e<��(>r0�=Z�=��5���>��ǿ1~�?*��;Y#���9?�,�y�+>Gy�=���>~�뽚��>+���8m�>�< >�:d>�=5�l>���=��þ{�	>CS�s@��C-���D�A�����=Pg��r�HG��[��F��ǐ���1�?Bf�h避�)?�|�+����?�ܽ90k�5\+�C^��
?m<�=�//?0R��_�;�B>@��>	�>�fؾ����R���K����?�D�?��\> g�>�x^?��?Re9�Y�*�K�f���k�-�9���J��<�_ǉ��&���\��D���E?�,z?-�8?|�}���m>é�?e+�������E>G��� �yљ=�M�>������C�n�꾂"۾�s&�Y�>�c?(��?!?
9�q���#>�9?}&?��s?
a<?��%?3a�zw0?�>\�?yA?f�.?*y*?k?25>��=��Q<�:�<?t���'���,�����f5
����<w΍=K�h<2��<� =�m|N=Z�=�,"��9�:M�;�J=c��=l˩=�">٥>�]?�R�>��>�4?���s�9�N���A,?��O=�'{�V���<J��g��E/�=D
h?v�?@Z?KZ>��?��;�<>[c�>�N!>CM>�;�>�v��nB���=��
>�.>y��=�i��b��/��P����<!�!>l��>x$�>�L����A>���Ɋu��x>}�i��h����J�Q�P��A5�Pa}��Q�>�L?��"?SH�=u�پAN���h�VR'?X�B?ߊC?bo�?,�=o�\�(�)�E�v�c�/G�><4d=��Ȧ��ޣ�&nC�u����#]>������<d�<�
�8<�K��n-_��|� �j=��#9�>:�%��K�d���i>�J=�A���*��˓�f��RH?�C>�b�p����V�=[E�>��N>�|��V��=\j��柾�^>�H�>K��=���}���T���#� H�>xOT?O�]?�?�/��G�`O�I�"���P��-A����>� �>J�?|��=:lb=�{�
R�nzM�U�>���
?㱼>p#E��j�*ѾBま�NG��5�>��?r^�<y��>��V?+�"?,X?S'?F� ?"�>V�I��}Ծ�H&?�?hj�=�#ս�T��8��5F����>��)?01C����>"�?��?��&?Q?P�?{|>̺ �vC@����>dG�>��W�Hj���_>�J?�f�>�[Y?�σ?��=>s5�墾�悔B��=z1>N�2?�"#?��?���>\��>�3-�=��>r'c?�%�?f�o?g��=a�?w�1>%y�>�4�=K�>���>�;?O?-as??�J?��>�X�<����c����p�:M���;�F<��u=^T��:s�,�=��<�;�;�z���낼�A��F����G��;���>Ԟw>����A>K��Ϡu�N>E��~��	D����3��3�==�>�H�>��>�0*�ߖ�=�o�>Gj�>���D�+?��	?	�?e���1e���̾��T����>?�B?��=z�l��K����o��U�=�;i?P�Y?��Q�O!�2i?_~j?�
�;<�uɬ��$�<68���@?R�%?^�-2}>��h?�[n?Q8�>օ�=^�8񛿳�p�*��U>�f>�B�����}�u>�E?G�.>q�?�>{� ��XF�uٙ�L�3?��?U��?�a�?P�=l�������+����(��24_?���>[��$7#?�P��JϾ���!ק⾃ޭ�~}��꒾�P��do"�i��۽u�=��?^�r?op?D�`?�D���d�ʨ^�$����U��g�8��?'E�1�C�S�B��uo�y�����8h����Q=�^A��D�\��?�(�>���:���>Ny,�a���3��E>����u�����ŽV6�<
z�=���=�W���q�x���?�N�>���>��^?�j��Y�m?K��5����D>_��>ل�>��>'���˒��oS�{���
_���9�P�v>.�q?:EH?��k?�C�)��끿�=�P =dlȾ�7�>��E>\Kf>j>���V�V�3���?�y�b���!p���}����=��??��>(��>�o�?rV�>�L!�����G2��Q3e�:��))�>�;d?io�><�N>R_d��L-��4�>X��?�_�>�&h>t��T���ӆ��! ���K?$e=
�;?r�5?F����"��ւ��zJ���7�IP�=�͖?Nsn�N	T��E�>r�=?m��=� >��2>���o��k�������#����>[ܲ=Z�[>������ �/k��ɻ��o?��>5P�q{B��ߧ>KP(?�?�r�>�~y?��>X�ܾ�D�����>�Y?�jQ?7!>?�>�ь;��ȽT������=�׉>RV>�C�=��=�o�k�M��Q �,k�=��-=�%<�3p�h�ż
/��xU�7Y"=v�>)ݿ��N�A;޾���(����mu���Q�́�����y���Q���^�[���U��,���}��n���7�c��?,1�?����1����� ~�0Q�|��>9������Ⱦ����i���׾���D����L�5�m��u���'?񹑾��ǿ����u9ܾ�! ?A ?A�y?����"�%�8�'� >�W�<O:��y��V�����ο᧚�*�^?��>K�/����>R��>3�X>:Lq>���螾�?�<z�?�-?1��>r��ɿF����Ԥ<���?��@�R?��H.��\>��?�MN?��c=��;��=�PZ�>���?���?�,ڽB��f���zJ?.���A���� <��>�_>������J>�/?C$��b���4S>A�=��=?�$�d!��es��}4�Uܲ>��J>��=�`�?ߺJ�,y���3�߶S���<�T?��1?
�>�e?27y�,ѿ냃���?@�H�?�/d?G⻾e��>@��Zlf?��I?X|�=�f�Z�I��>g$Z>\*�=����b�%a�=�u�>9E9>�kx��<$�s�R�S}�@�d>$�=�ſBA%��u#���x�:ȳ��!8��Ž���i����-��S�q��׽��V=�'�=w�\>�zx>�dP>��K>L	V?��h?y��>'>���[���7Ǿ~{B�(��A"�Ψ���"�6���XS�	�߾e��ӷ�/��\�ܾ�G��|
=��Q��ԑ���*�o�c���>���/?��&>���<�L�v9��/������im���Ҿ@�,�}�i�i��?��;?Q���T�����q����VR?,�-�ێ��;�¾��=�7�
=Y�>L��=Df徆8�q�^�hg2?a�?��̾~����nE>����/=]�*?���>���A�>l&?P�	�t�.4J>��">C�>��>׳ >�q���@��c� ?�7U?���­��/o�>"�ľK!U�w�=nN�=U�J��6$��/l>\A�<�������hOK��K=a�V?���>�J)�����J��N	%��3=D�v?"y?���>OSl?��C?�R�<fI��|CT�l��h@u=� X?�j?��>�~�Aо�j��h�5?��d?)�K>.Vg��Z�m�-�����?7�n?v�?�檼��|�#"��u�EF7?��t?�&[�K������{r�YE�>�c�>��>r�A�v�>��A?R6�k�/߿��4���?��@Cx�?��=���fQ8=���>��>�5?��������ʾ7�y=��?�c��a���Q�)������J?jԎ?�?������>U��(�?�eu?�����z��{���d�������<���=����s��g�Ⱦ� ,��������׭��@��Ǉ>U=@5�4���?�5˾����̿���ӹ־�����4?���>��:�¾�Qn�y�w���#�z��
7��̣>7>�*��_��/S{��w:��Ͻ����>����A�>�ET�g/��?����R'<�ϒ>��>��>���GF���љ?���wο�'��T��v&Y?7��?�م?��?(�<��v��{��K廂LG?��s?�lZ?��)�A`��>:�.�j?�[���V`��4�}CE��&U>p#3?�A�>v�-���|=4>h��>Fr>l"/���Ŀ~ض������?��?Tp����>���?�s+?�h�y8��8Q��>�*�^� � >A?�2>����!�q,=��͒�4�
?�{0?�v�+���_?Ԡa���p���-���ƽ��>*�0��6\�i���o��Ye�2��B�y����?�a�?�?"O���"�./%?��>v���Y%Ǿi��<?��>J�>l&N>�{]��u>�*�:��3	> ��?���?7o?a���������>��}?3�>8��?ʫ�=�?tPt>�J<�T��=�/>\?2>�X�=��>�'A?�?�s�=�#��*���&�� 5�9����b:����>7N�?C�E?���>�C�5�a�\�p�(�
92��9o��M�;*$�4������>Y?>�=UE�d!쾸�?�a�Ńؿ&Y��Q6(��4?v�>�!?���t��z
�-_?;<�>QM��2�����w� �ϥ�?�2�?�3	?�F׾��ټ�>�Q�>���>�@ֽ8/��]� �8>�B?��?Y��W�o�;C�>p�?��@%Ү?B�h�S� ?1��i���}g�vN��k��|�W>>?�Q$�["z>du?���=�h� ��r��W��>���?i �?yS?ہ?CO��U�B��=~�]>���?���>0aԽ��A��>��?w�@�y�������w�?��@��@ŮY?�.��>yǿw���;���Ƹ�9���7�<Ev>{��K>RQ
>(AI="qs��c>��>��<>-qX>�@�=1h�>LuX> 7��>7�Ὕ������H��'@��l��vK������<�0�����e¾M8	�� 5��¨=O���v`��v�R��=mKW?�yQ?47r?"�?�AL�m&>���k� =�P)�ĳ�=��>1�3?w�J?��)?\�=�M���ab�z�G��撄���>��I>t�>���>^��>�\:PJ>��D>:�>B�>��=q�C =ɪL>��>B�>���>�ML>�)>!Ĵ��$��-e�oV�]y��6�?2��K$P�Q9�����)���ե=I�-?�w>��V�пШ���XF?����ř��e2�>>2"/?5kR?u�6>A���Ry�a">i��bG� 0�=����(M�ԥ&�U�<>¢?L䶼���=�R"�
_'���c�����}�>,
-?�J�N��=W�^�p�9��{��F�>��h>/��=�k�R���6��x7a��E�=n@-?��?�K=5��O��&�D���[>�!�=���= ѻ="g�;�|a�ʍl��Wm����='�>���>\<?E7>A~=���>V%��(A�֫>�Q6>�o3>OH;?�N%?��弩*��僾m�/���d>ή�>���>��>^�K��=ͣ�>��d>9�2���`�����F��f>���(8_�C�\�#t=���5u�=ӌ=�@����.��<*=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�'�>H��>G��#	����u���"=��>0H?����v�O�E>�~s
?��?�s򾚱��:�ȿ!;v�U1�>���?���?ρm�rQ���
@���>��?hBY?��j>z�۾�^Z��@�>��@?"�Q?���>�0�2'��D?�߶?��?.\P>+#�?�m?z��>����}�%�aD��D����">��C�os�>��L>v����eQ��%���w��%b�ߠ�At�>ؑ=&r�>~��1���s�=���(>ľ�孽Oi�>&�D>��>��>��?䤿>���>Q��;����!��}G~��]?9-�?�:��!a���=-�>{��3}/?6c,?a��������>Ά}?�sG?��??�<�>b���X��Є���Ҙ�q�ｘ��=�?��?����f�>0ݼ�������>Ej�>,>���$&���R�}�>�5?���>�>=,�?��+?Y�r>Gϧ>�F�^s��}dC���>�f�>Y?�B�?v�?￾U�9�i����;���[Q��}>)lz?�?#q�>E��Gi����e��M%�	���9*z?K�k?�n̽Ղ?h�?Lg=?(�5?��E>�<�[8׾թ��3��>A	?��9��e&��k5��y����
?2G?���>:o��$�����g"�'��q�?1}_?{�%?����}]�8C����<= ��j��<}T<<��;�K>aK>�2����=�)>{��=�G{�V�$���=R{�=�5�>`h=�l&��%���<,?��G�Qك���={�r�xD���>�LL>}��*�^?�q=� �{����Gx��CU�� �?���?�j�?����h�#=?J�?�?�#�>bI���|޾���|Kw�M~x��v�c�>#��>�l��)���#���RF���ƽB�O�>��>��>�H?�mD>�L�>� ��A"��%�s
�@_�����5��E&�+G�hힾ�T.�F&�R���9���R�>ó��5��>j�?D�_>�p>���>��4<n��>'�I>g�_>�V�>2?M>J�'>���=�6�;4S��R?�Ķ�lS+��jӾ	͝� H?�e?�^�>��3��ȃ�����y?'ؒ?.�?Ftg>�f�0�"��;?}��>"����?�ı= 8M<"9<bsƾ#QٽIo��_D#�]��>�����R;�qrH���N��w?TJ?J�ԼѬľ%`��ݜw���=��?�?�d+�~�P�)�b�)?V�]�A��d�;?�Ľ������'�Va�w����~��ps����y��=�??���?���Ǿz$���d�	q(�$F>[�>�~>{g�>�P�>����@��Z��Z(�<ѿ�1�#?n?f��>'P?��<?�&]?�?Z?ۡ>u��>� ���+�>i�P����>���>�@?��'?S.-?�n	?\�%?	�c>���������Ӿ�?P�?,Z?�J�>���>�h��H��� �<=^j:^��Op����=;V?=◲�ë��g�;=�N>�Z?Y����8�:O��/xk>t7?�@�>Ա�>�ԏ�6��zo�<<�>�
?
d�>�����}r��S�8��>���?%���=	q)>C��=���6T޺9�=�i��"�=v^���:��[ <ܶ�=Z)�=��y����,;N��;���<;��>3�A?���>��j>
̾y���7���5�z��>�!�=&��>����Ɇ�[d��_h�uՕ=Z��?��?��7>��=�]>n����Gྌh׾�y�������>7J?Fy#?�ׂ?�r?E�?1�@��ǌ����l��"z��8?f!,?���>�����ʾ��ԉ3�ޝ?i[?�<a����;)�ܐ¾��Խ�>�[/�X/~����ED��������F��/��?꿝?�A�N�6��x�ӿ���[��o�C?"�>Y�>n�>M�)�t�g�r%��1;>���>jR?�L�>�rL?�x?S}\?ԭ`>��4��/���җ���R;�!>��@?`�?B�?2]w?ֆ�>�>��1�\�Ӿp��A�缤9�H��|P}=6'U>�Ȏ>��>��>�h�=��½����#+���=��a>��>��>���>-��>M�9;C�G?���>�C��^�� ��˃���<��u?��?7�+?4�=
~���E�@M��=�>�e�?~��?i4*?ţS�u��=�,ּ�ڶ���q�e"�>�ݹ>�.�>	��=\G=�>>��>l��>?F��a�\o8�UyM���?XF?���=���k4e��<>G�z�.�� �,vn>*���g{ݾ\��>@Կ��l��e��MC=�`ž�N�z񤾄O���ԾZr�>����_
>xK�= `>�˹<=�_����<��$��ܢ�� o=G�
Jj��A��2�����B>Zj�>���}#�?�H?��3?tK?T*�>h�%>���Ü>,��q?~_>l~������Z,�p���j?��f�Ͼ_E۾I3g�Ԗ��gc">�&�P%>݁/>2��=� <&��=;�=k��=��	<���<j �=�J�=Ks�=�z�=:�>J>;�y?}��^��{/�#Q�>\?�>��<v���R?}>}����H����ޔ�?�Y@��?�/?�Y����>+5ҾvD�������=��\�dн��;��W�>�
�=�b��㖿{���p�?͜@�OK?gĕ��ҿ~�==�Y$>� �=��P�'�/��<f���n���O�qf!?ɴ=�����M�>)Q�=�yپ����C�=��8>�_=��(�6P_��p�=�?y���S=��|=6�>_I>�0�=�̳��-�=�7=���=�ZL>/����A�����	=h|�=��l>$�/>���>��?6t0?�"c?��>��r��mξ�.ľ��>U�=��>�=�7;>��>�Y5?>A?�cJ?�>>��=�>0R�>��,���k�L�羘@����<ق�?�?_�>��<X�1����!'?�p�̽�r?�j2?H�?/ܝ>�1�n{���%���-�$ח��'�IM/=J]r�/&Y��+��r���㽯�=�D�>���>[�>��x>��9>�M>!'�>��
>�<�<�=?ď���<�b��5@�=�G���<�lʼa�7���$�0	.�B�����};B��;�k<��;���=���>�>|�>2%�=���y�/>31����L�N��=Z§�>3B��Dd��*~�r�.�B�5���B>��W>8 ���&����?c�Z>H�>>ȁ�?i>u?5�>z��Mվ�0��ήd�� S����=�0>Rp=��{;�+�`�7�M�ӴҾ��>=�>
�>��l>	,�E?��hw=$�lV5����>3f���W�w)�<q�>�������i�Hպ��D?�D����=�~?��I?���?���>䘽+�ؾ0>)@��ǁ=K��Lq��h����?G
'?���>�	�F�D�! ȾX���-�>*"V�J�I��������Q<Mtݾ��>/Щ�����tB!�T���x�I��21�I��>�U?��?' ��4�O�j�1��h�=�p�>|�z?��>�?�>o�*?o."�b��j��M�;jlS?��?��?wL�>���=����q��>=�?���?p�?w�V?N�C��I�>/�@<�W>]�Ӽ7�;>��2>E\9>¬<���>��?B�>�:d���*`�R̿��V��#<?�d=��>�j=>M�f>qs>��>S5A>��[>|0�>�\>��C>���>x>�ʋ�:���b<?d�Ƚ.��>�?Qé>�_E>iA)�`m� �I��֋�x����|��d<�7�=�����aZ���g�>>:��ʎ?l�=��o�2?�oܾܯ�y�T>��>2���?�>bb�=b
�>���>4�>�<c~{>���=�پ�=�`��J��5:��UR��4���J>6茶�4�*r��_߽�BJ���������g�# z�)�-���=�A�?���9�h���0���J��
?�;�>��;?����\���n>,��>�:�>�� �"/���4��Iɾ���?+�?�d>�3�>S�W??_?�k4��/5��Z�g�u��@��d���^����������
��ý�|^?�Tx?��A? #�<�y>�?4&�.����ǈ>
�.��a:��b/=Z��>XM��X^���о�þd��ҢC>�n?�K�?�?a�T���>J�I>&4?�v?��?��*?o?�>�T+(?B�=,$?�-)?]�d?`?z?�ҽ�Ę=��x>����LC�ț��|���}Ѽ�]b=��<��ż�<\��x>=Ek>e7�=��g=�Q�<Uy�='�%;���=/��=a�X=n8�=�¦>,�]?pR�>��>-�7?-��m8�Eݮ��*/?�e9=� 	��6ޢ�0%��>��j?���?�lZ?�qd>��A�.�B�� >�<�>Vn&>x\>.U�>����%E�|x�=�\>�>���=B!N�Iف���	��}���=�<M@>�7�>N�9>��=5�S�S�{�	P����>;=
w��u���O�v��C��ﺾ<Z�>�j?�H3?hg>�u⾢f]=B�m����>m? $
?�z}?�Y>i����7����h	����>Df�=�)��6���v��"J�祕�]9!>X+龨��$�>�㷾Z��Vǁ�3�o����En�={� ��19>܃���Ѿ�{�q>"�S=�͛��%%������򳿟w7?���=��%����;|���G>��>��
>�j��oB�/�C��j���u����>ƈ>� ��H4���^������>�"K?��\?3%�?W!_�Db�~w;�A��(T���F���?ѹ�>��?�">ճ�=�������a�тH�A��>W|�>h���d?�|#m���ݾn)�4x>V�?�G>��?�qT?��?��i?�:,?�`??��>��e��}Ⱦ�?$?���?�u,=럴��F2�s,9�"�L���>�n#?&Wz��l�>j�?��?6V+?��Z?h?Ҡ>�'��&1��Տ>�Q�>�T�������^>F?{�>�W?J?�?�.>it/������4⽜7=O�&>_6?
�?��?S2�>R��>~�����=n��>vc?0�?T�o?t��=��?':2>���>��=қ�>��>g?OWO?�s?��J?o��>^��<�5���:��BBs�A�O��W�;�H<��y=>��~1t�H����<�(�;�f���H��l��V�D��琼���;���>�1_>�吾6�>�P��b����I>IrD�4���Z���`�LU�=�݅>�J?%j�>8^@���=�[�>�.�>�j��R"?��?;{?�R=l\��Ծ�);���>b�F?K��=�so�����kUw��^�<g�d?��S?y�b�����N�b?��]?@h��=��þj�b����f�O?9�
?=�G���>��~?b�q?B��>!�e�,:n�&�� Db���j��ж=fr�>GX�H�d��?�>f�7?�N�>�b>%�=\u۾�w��q��g?��?�?���?�**>��n�W4�������C]?9R�>3Z����#?o'�=�پ�Ύ�\i���?꾿G�������ۍ�������(�A燾��ǽ�?�=�?U�t?S;m?jc?x����c� =[�
m���V�z����%�E��#B��#<���f�Q��m�پ����j{=v�v�Ao>�4�?/�?���R�>#����5 ���Ӿ�/I>O��n1�ԟ�=�8��I=��(=�2r���"�{`��X�?�t�>�(�>��>?��_���=�^�0�,�4������#>��>E��>Xk�>oF�<2���h��o��77h�v�}�LHt>�d?YK?�Wn?����Q/�;���� ��1&��r����E>LF
>���>��`��#�K'�?>���r���������4	��g�=�D1?�F�>rk�>@ǖ?�$?,��Zڭ��wr��0�P
�<�_�>S�h?b��>¡�>%�ɽ�E!��P�>Y,m?J��>k��>%)��N~���g�r��Z��>�3�>2E?��>-���"c�ڪ��b}���(���=*�f?H镾������>��X?�լ��+7��/�>YƼ�}�?�Ծ��F����=�*	?�.�=��,>�bɾi���Ly��O��G�'?k~?�t����)�U��>+�?���>�Ɣ>�U�?|j�>|�ľΈ��$
?��]?��O?�J?�R�>=�<���yʼ�.t&���=�=�>5M>HM�=���=A����X��]��7=�~�=q����սl�
�S�༢��<_��<�->�濎�W�>��������N�6���c�7�C=6�Ͼf�[=�O���e�����Q�t��F�:\G�&��Je��vx�?`��?ڱi��ѯ�M��!����bܾ�f�>�$h�ZF�=F����0����sc���gR�!
�� %8��\��a�g�t�'?CÑ�B�ǿ5���3ܾ�  ?�E ?��y?c�	�"��8��� >��<۳��ƒ�����οʦ����^?��>�� ��0�>-��>��X>)Vq>���ើ�<��?��-?���>��r�ĕɿX����$�<G��?�@`�A?�W(�����MT=Gy�>m�	?�i?>l /����;���S�>i\�?���?�)D=`X�AO��le?a�<_EF�N������=�=��=P^�� I>Hߓ>O���B���۽84>���>�����uZ^��W�<U.\>kڽ ���5Մ?+{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?_D6?���>�d&��t����=Y6��z���&V����=[��>a�>Â,������O��I��W��=��L�ǿH��W��b��<n$��Y�Q�7���7��(J�t���B^�f፽M��=c��=�a@>u�z>�AJ>�6>��\?s�o?�p�>�G>W
�D���v��7� =Ć����$o��p����?�i� ��"�� ���j0ľ��=���=�-Q�z���!�7�c��rE���.?�� >=%Ⱦ�tM�H�<��ɾ��������z����˾�22��qn�
��?�B?X{��ȞV�Ͷ��������6�V?����d�
X��4��=������=�N�>ҡ=Cu�l�4�l"T�1�3?{X?�!Ǿ�w��S��=U
��A��<�%3?�O�>V�B����>4�9?��#���0��\>��=�>�n�>�bJ>�ø�>��=?��`?�f�ة����>R���O��7j�=�>�=��'�c=hPu>�L�;QB���(������	=R#f?*bn>�b@�9�5�>Ǿmm>�G���l?\#?֌>e��?��r?�Z��9� ~�]�Dc�>knt?�fC?ϓ=��>J�9�#{��1��>��?��>r׽�u�5L��vѾN?�S?^��>�q�=D����֖�6$N��hR?;9{?�B��P��ώ��v{�t�?�v�>]�?t\���>��_?�B�=���v���[��ƞ?�@\b�?�c轈�#��m�;�t�>��>+�I���Ӿ���r{׾O���P�>!��ƱO���P�V��?�@?���>���Y������=�ו�CY�?~�?;����Rg<����l��r���a�<o��=
K��<"����G�7�i�ƾ��
�q���MY�����>zY@Cm轓6�>�P8�:6⿍RϿ��
^о�dq�w�?|�>��Ƚp���d�j�LGu��G���H�j���z��>%�_=�,��J\�5�o��KB����:'�?�"a�kC�>��p�����:_���<9Ý>F�>���>V��;��i�9�?�!��)ӿ�������w�?�3�?ۜ�?�M'?4�6>��=@�����"��- ?�Ia?�5�?̪�`Ƚ�$�ʔj?���}Q_��q0�w�G�o)[>£1?b��>�E+�j�J=�$->��>t>(�0�m,Ŀ���� ����?:��?b�� ?꼛?�$.?����͙�R*��?"+��ķ�A?h(>�ʿ��e�29����F�?++?�v���Re?-l��Ћ��^ �c޿=�F�>�8�=�=%=Wr#>�P�>��8Kv���?���?Ow�?ђ��� �A�?�0�>�i;n6뾀�5>r��>���>Q:�>6Hn����>�A�-H4�㧎=��@�K�?=\�>K���ec��:*T>��?dG�>܅�?���<�u?��{<�{���>BQD>��E=C,̽<�?�]?��>��F��ؾ�NL�"l/���D�cо��I�>c�>4gV?�,?+��>�� �н�t�{Z����������վTF'��	u��p�=~�=�1�{�a�k����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�$�?7�2��@W~�����V8���=8?����|>u@�>rU�=�~v������s�eͶ>3�?�J�?_��>��l?o�o��MC�Qc/=�y�>S�k?�?������=�C>1�?������hQ�aBf?�
@�R@�f^?sآ���ɸ����??��=E�<,�G��=q���G&>��+>��μ�?���/d>�Ş>�N�>J�>5�=a��=Ώ�=dǄ��(�䩛�����5��!���� g7�� �0�i����fG��TA��b(���{ ��Ǜ����gX��2�����=�&X?�;R?�Wn?UM?�=�H�>v� ���=P&�Oө=��>�2?�G?}M%?��p=s���]kb�	��ҭ��e��-��>��I>`��>a>�>zɝ>�<�zL>�.>>]��>#�>��:=Q��<�K%=RN>��>���>��>C<>��>4ϴ��1��p�h�Cw�q̽&�?����>�J��1���9��Ԧ���h�=5b.?|>���?пi����2H?%���`)���+���>x�0?�cW?�>��f�T��9>T��Ҧj�>`>�+ ��l���)��%Q>vl?�_>�s>��1��v8��-Q��㲾"]{>�%5?'g����6�ƻu���H��ݾQ�M>��>� L��K����������g��Wq=��:?P�?�}�����-ns��H���AQ>�NW>�?=dǥ=7�H>�a\��1ŽOI�2w=�(�=�a>�/?�(2>�
�=ޛ�>L��#�Q����>=�F>@k%>� >?��#?؋�0���
��g>1��Vp>��>�{>��>�L�ֵ=�^�>��e>����̓����]�G�O>w2M���i��τ���t=�+���B�=�g�=�l��t7�'D=uԂ?����#��s�t���?���i?�j?�a�j�,>]Dܾ�m����о�s�?T�@D�?���`��I^?x��?��i���1>�?	�G>�M(�C!=�&�>�f���Ⱦ4�T���N�?�A�?o =�!��i΄��-�>��%?��оPh�>|x��Z�������u�o�#=Q��>�8H?�V����O�f>��v
?�?�^�੤���ȿ4|v����>X�?���?h�m��A���@����>;��?�gY?voi>�g۾:`Z����>һ@?�R?�>�9�}�'���?�޶?֯�?t/>���?�>s?1~�>f3���0�o⣿�m���'�=����>��>ᡠ�"�O�bޑ�����wkd�jA�!Y�=��<d�>	xؽ����r>>ڲ�;����V�����>~�>�ϗ>|��>а
?<��>�_�>c��=��,:F$� ?��v�K?���?2���2n��Q�<���=�^��&?uI4?�y[�|�Ͼ~ը>��\?e?�[?�d�>��E>��!迿~��ϩ�<@�K>4�>qH�>$��;FK>j�Ծ�4D�`p�>�ϗ>9����?ھ-��X��!B�>�e!?���>dҮ=� ?��#?S�j>�(�>EaE��9����E���>'��>sH?�~?9�?�Թ��Z3�����桿ݑ[�2;N>��x?�U?�ʕ>�������E~E�iAI�4�#��?Ctg?VR�S?2�?��??n�A?�(f>��3ؾ������>��?�:����A�O"��o�����>�>��>�vy��}����^������?��r?��M?���wdY�����q� =!㼦q��SV���I�b>��=�Q=���=�k">h��='�K�j�]��f\��E>=!�~>���=�� ����@I,?	H�C�����=A�r��7D�}�>��L>C�����^?�<�a�{���|����U����?8��?v�?8���~h�=?a�?��?N��>zh���t޾��?�w��y�{m���>���>�Oo�y�侠���I����B����ĽyQ�E,?���>��?���>l�5>_~�>7\a�H����c�ž-�I�o	�S�b��0E�I*D�5f۾t�������tƾLji�*��>|������>�Q?��.>�q�=�z�>.җ<C�>�$>�M�>nվ>���>-^~>�B�=����.���J?�~��4D8��8�K��.�)?Յd?��ڼ��Ͼզx����T>?QϠ?T�?�'�>�`��3,��?�&?��ľĀ/?�|_>��#�3��>�	�1��'��X!�t_�>�?��pL��mr���۾c]�>��>^V½����(7���¡�#�_=�b�?�~(?/�*��R��#n��BW��S������j�ⵢ���$���n�aN��񖃿�n���>(�^a-=�/+?�7�?w���K�1���<j��#@��i>��>���>wB�>7zN>���N0�C}\��@&����Q��>��{?/\�>J�I?<?��P?�L?Î>��>������>fR�;o$�>���>s9?n�-?�0?�B?�S+?�Gc>%�������Zuؾ#?��?�T?i?a�?85��ռýꖘ���s��gy��׀�q��=75�<��׽�w�
�T=hqT>�k?��i��R��b+�U��>+$?�Ĥ>.��=M΍�{���g%a�*�A>��>(��>-Ͼݦq���9����>)Yu?C���I9����~>�ֳ=�ȼ
��=W>ݽ�$�B�}<}�;�Gp��=*�=|�=�K��S�=/�=̹ؼw�ȼD��>b�?�T�>��>^J���� ����1��=u,Y>TS>mp>��ؾXz���&���g��]y>u|�?�z�?��f=#�=���=�`���<���������͈�<�?'#?!#T?��?)�=?nV#?˷>�fP��`���-��W�?3 ,?���>X����ʾ�쨿��3���?�S?T=a����.=)�_�¾&�Խ;�>zU/��/~�����D�����M���|��g��?'��?It@�j�6�Ur����@E����C?��>�A�>t
�>Q�)��g��%�m;>�{�>R?엻>��K?}(j?��^?E�f>d�4����^F��.�M���=0y1?*zl?H��?0ʀ?N2�>��L>�� ����U|־���Ӫ�� ����==���>w�>�ܼ>�|�>��>>����T��� ���=�se>t�>{�>�~�>^�>>���<mUX?M�>lc��t#���־>��=���?km�?f�3?->�>�U����_��|�&�3>��?�X�?;i{?����"�#>J#9�D��S��+��>�d?%(�=x�=bL�>+�>�y?���>�7=��+�)����=��?=ta?�p��ձ�lQ����>*r�����;�,����<��0��YݾwO�=6���Sо�U�/݀<1��[|���� �%�_��U?!嵽�� >�=@>>&D9/U����<���ܝO�ܪ=ַ��V-�zx��ɐ=� �#	:=U�>���>�>��
g�?cYp?L\?Ɔ?xW�> ����-�;8H?uF���^J?+�x>6�=�*Ѿ�w��d ��z*�ɟ_���B�N�<�����	-�=����ec�����~>!��=�T!>�=46�����"�~��4>WM>�>��=�w>�^�>��o?և���r���T�!���P\!?xd�>��>,���Jrs?��>�ً�5���w7ܾ���?�<�?��?��>%u��o�>clᾲ��"	�=$�C>Y�>��a>3�A�'3?t�P>������ጤ;PZ�?@�@yw@?�����ʿ�;��7>]>��R�E�1�E{[�8�b���\�r!?�	;��̾v��>]��=g ߾�žD�5=r�8>ʲb=Ȼ�?�[��=`j{��Y:=A�l=5u�>,�D>Y��=�����m�=E�J=�5�=;�O>����Q:�>�-��2=5i�=YMb>X�%>�^�>8?+��>Lo?���>���Z���ϙ�E;�=I?��� >��=,P�=���>��f?Ԑ]?G1N?*R>�TT>��>FG�>�X1�l	���e��O���9�<���?��?��Y>���>�U�f'��U1��ϻf%?2�?C/�>�L>>7�X��x���4#�����4�+|$=t�r�e𚽱��;�����>3y�>���>�R�>�`>�X'>�|'>89�>��>ըa=�C�=!�9�>�<���=F��=��
�s�����<����eO�l���#�	M=(R�<~��j��=���>l >K�>�^�=9~��X�9>>�����J����=�ᚾ��9���`��8���4���P���4>��D>f㐽#��:J?�,h>�68>:��?��n?6�=L�G�о�\�������yu�?��=���=��:�5':�m_�E�J�ע޾]��>���>(?�>��u>ڵ)�6`:�fΛ=4.۾��3�ϊ�>&b���;�����]rs��t������f�dZ2�g�A?pÇ����=�x|?۠E?q�?,��>s����iؾ��+>s}����;���%~��V��Q?r�!?��>�뾭�H�ޑ˾�u(����>qY���\��h���'���<@ྼ��>�亾�hľ�2�6[\�I��8+�g�$�q��>B�I?�ɯ?���������4W�����W�)��>�n�?:�J>K!?	|�>��M�7��Q���}@�=bg?W��?'�?@>=�=.���3�>XQ?�Ֆ?���?~r?5yA���>��[;�t>�C��ٰ�=ܡ
>�ۚ=}z�=8�?�.
?�	?�杽܍	���#�Z/`����<��=$R�>�-�>ܲu>���= b=�8�=;�\>�ў>$a�>�h>��>="�>�c��Zk��'?w��=Ι�>��/?�c�>�eD=����;�<Q�^�B�F�+�d�����y�<���$>K=@��f��>�lƿ���?ЬN>!�0�?�����$�e9P>��Y>�ٽ���>�hD>�}>]��>�ݣ>�+>e��>4M+>&rӾh�> {�s?!��BC�9�R�Q�Ѿ,�y>�ۜ��0%�����X���I�=���W�l�i�����5=�H�<�F�?;@����k�x�)�����|g?�Ĩ>0*6?�ތ������>��>���>�����i������U����?���?#�z>�Ê>Y&A?X ? 	��:���X��e��z�S��CN�Vi�!g��X�R�Ϥ���Н<ÉE?��d?�6'?V�Q>�H�>�$�?5�7�Ify=�� >�GM�,6��ŧ�KKZ>���l1��xᴾ�#��bt>-��>ˆ?**�?�}�>@����ս�e{>� N?�!?�gn?�u?1+?��V�/SC?�0%>̒	?/7�>9T*?�K?��>1H>��>Dme=H�G<	�a�sm���彣G���ze���`����=?2e=�u�<�OQ=08=�R�<����aOa<��X�=��_=�	>���=K1�>�:M?���>���>��'?`~���W�ҕ�al�>�q��Ѿ.Ԅ�䲽�+��5�>ѭ|?�k�?.?X>�>�h ���5���1>�^�>�a�=�=>y>�>�߽?}~��	N>�<��3>{��5�ѽd�E�6$�%R6�y
>a�i=���>f@�>{])��2�>�F�8򆾴����p0��D���o���*;���o~��$��>�Y?��'?� �>�[���p=��Q��?z�U?�U�?B�O?�+2�,��ۃ �N�P�a)b>�B> ����о=6������X`�>->� g>Π�S�����I>x� �&)о _o�'�P�P���/=.�J�=!i��Cվd���c�=c�=�'��� �����Y��YJ?���=}̘�B6�5��j >���>.*�>x�F��D�'@����)��=�P�> >Ň��"�4J����>�E?�h_?�N�? !���-s�]�B��s��Z���2�ļǫ?��>�6?�B>]�=�b������d���F���>z��>)����G�ͽ�����%�ߒ�>�/?��>�{?,lR?,�
?I`?*?BX?I�>��������u>&?���?�Ԅ=�ԽA�T���8��F����>w)?R�B�%��>�?�?��&?�Q?ܻ?7>v� ��<@����>�Q�>u�W�_���`>/�J?8��>�>Y?փ?�>>^�5��⢾D����=
>��2?`/#?��?���>f|�>�@���}=Ou�>޿b?��?��o?�&�=��?�0>��>�2�=���>s_�>�g?�O?�t?�K?��>�U�<� ��T��U�p��@��"�;O	+<�*{=����<Gk�*���E�<���;�K��}!�����P�G�\���;��;��>�@6> K��A��=�w�� ���^V�=�=�1M���䇾�؀���S>�5�>l�?ҷ�>���	=�E�>B��>z|,�|p-?���>�`?�G>sg`�7h����|�>$C?�㽪〿�ᓿTq���p=�Q?�@?4M����ݾG�b?��]?Sh��=���þR�b���r�O?%�
?��G���>��~?O�q?��>��e�>:n�4��	Db���j��϶=�r�>"X���d�P?�>G�7?�N�>��b>�%�=iu۾�w�r��N?h�?�?���?l+*>��n�I4���֒�%�]?O��>����!?��=�վ�.��}`��~�ླ$�����V����E��k�?��<���=S�?�r?�[m?n�W?���Y#c�3[[�(�x��U��,�:�)�?�ʝ>��y;���d��V��_㾇���^F�=7����U^�Ϥ?�3?T�R�T!�=_»=��
��~ݾ���>K禾��m���Z=�6�=Y� �/��==,c���/�J���,?�v�>s��>w�?�dR�9>;���(��I� ����y=��>
�J>I��>o��=���/��<����}�<�><Ac>" h?�4N?��h?�3U��;*�{������¶;M'���8>��>m܇>'x�>M���)���C��t����ѕ����X�=/�2?4�x>�u�>���?��?kG��6����?<�-0$��e(=k��>dg?���>u?�>i���z$�r��>�8k?4��>+[�>�7�������|�>Ó���>SS�>9^�>,�> 7'�Q_\�����^��ް>���=�Ll?� ��Q|T��<�>�tR?'c׻�f����>F鋽,�����>n8��h�=�?��=C/>WľŔ�t}����و(?��?���/�(���}>�i ?���>o��>��?Z��>��þ�ျ��?��]?�kK?JtC?(�>6�9=2����ʽ$c%���=o"�>y\>��z=tf�=2��ѝX����zO=�=�6⼑ý��ф;!����R�;L��<w1>݉ؿ�VI��쩾�/ �x��/��Єw�r�ӽc���߿�{i��1~��L�u�eѽƵ��e#�2�Q�Jd���~j�8��?ު�?f/�����["��/%w�n�	����>J~X�Qđ�m>¾?t �Z��LԾ�۠�O���A��=b��D]�r�'?�����ǿ����9ܾl! ?_A ?��y?s��"�
�8��� >~F�<�8��7�뾭����ο����M�^?���>\�2�����>���>c�X>�Dq>Z���螾�C�<�?��-?���>J�r��ɿ(���`��<L��?�@��S?��N�)$��#���>��?7��>*&�t�B�8���?���?���?"��>��R��y��\h?�[н�삿Է_���c>n:N>J�⽶uo��K�>��>�DоsL���'�=4%�>S�?����b۾a?��u?�<y��>��Ǿ|ɼՄ?�z\�sf��/��T��sT>��T?�*�>�8�=N�,?7H�F}Ͽ'�\��*a?�0�?ۦ�?2�(?�ڿ��ؚ>��ܾ��M?KD6?���>�d&�,�t�9��=!)�����"���&V�_��=e��>�>��,������O�|D����=��̙ƿ�$��J����<��b�?]]����Hͫ�B�Q�/��\o����h=�j�=�+R>o�>��U>1!Y>�EW?��k?d�>z>g�彈뉾��;��
�3�����@ꋾ����<�쾵�߾�G	�l���<�bYʾ=�ˋ�=#�Q��d���!��c�wF���.?��">�>ʾl�M��(<	Mʾ*/��$��� Z��J�˾d1���m�ֹ�?��A?��_W�^d����;漽 X?��[�髭���=ᛸ�N�=>��>Ǒ�=ye���2�2FS�7�/?Nq??���������(>>�$P=B�*?�f ?#�2<���>Ԛ#?��/����G�^>L�6>�ӥ>M9�>c	>�î���ֽj�?sS?��JR�����>L"����z�DW\=>ga3����-W>]
q<k����0h�i�����<|Qe?�9�>)I'��-w��]��?��!=ḋ?���>^X(?h�?O*l?�r��*��Ndd����N}>>*�c?-X�?��=1������w��"?]|?S��<Ӟ[�c�
������w�>��I?T}?Q�����l��T��[�1�H�$?��v?�r^�ss�����y�V�j=�>�[�>��>��9��k�>"�>?�#��G�����xY4�%Þ?��@���?��;<Z���=�;?(\�>��O��>ƾX{������6�q=�"�>܌��fev�����Q,�C�8?ʠ�?d��>���������=ga����?z�?�w��*��;u��t\l��� ���<��=%x!�n!�8�8���ľb
�*o�������݆>:L@U��B�>
�8���῝NϿ�ׄ��uо�r�}�?~�>��Ƚ�䡾�i�W�s�՚E��|G�>��fw>M���E"�<�*��������S��`�ҭ?�Fo�举>�T���3
���Ǿ ��=hܞ>ܧ ?B��>da�\{�����?�J�]�ο�(������r?�r?oЋ?bF?������^��e4�-�:?���?�X�?>8��>Tv���彨�f?�Uo�]�`�(&P���� �T>��>��?�"��r+>��>%�?]�>�O4��ſ�6����0� �?��?���F,�>�M�?�:?����5��qfҾf+����m�G? �=8�s���.��������>�?3���%����]?e�x�C����%�:����a>�����7ʻ(F��P^�&�c�]	��S懾�׵?H@3��?�n�����?�L�>w�˾�+���=1D�>�>{��>	�ؽH/�>�fH��& ���d>��?�@v
?u᛿a����Qx>���?�ɫ>鳅?*��=���>D�/>��fC<��R>��$>���ϯ�>�d9?
}�>��E;��I�B���U�&�l�d��EvQ�>��>�u?O�R?��>�2�ݖp���.�^G�<!Ǟ�����p���� �&4�1�>�>p�%>��:��l���?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��&a~�A���7����=��7?#0��z>���>��=ov�ջ���s���>�B�?�{�?G��>4�l?��o�|�B���1=�L�>ڜk?�s?2�n��󾏳B>��?������L�xf?��
@cu@��^?��m����r������]�=G�H�6�=5������D2=e����U+���=���>HG>�;�> >���=�'>�X��qf����V1��W�S�p�=�
��1O.�u���r>�:���hо5ɽ�6I��q6�2�t�����dD��m�=A�U?*BR? �o?j�?�Rv���>�����R=�r"�)b�=�Æ>�
2?JWK?c*?_��=k螾�d�#�vy������6��>�%K>-��>��>�a�>d�;��J>ta>>���>�v>ӕ+=y���q
=��Q>�>U~�>��>�C<>��>Fϴ��1��i�h��
w�o̽0�?���S�J��1���9��Ҧ���h�=Gb.?|>���?пf����2H?'���y)���+���>}�0?�cW?!�> ��q�T�4:>:����j�4`>�+ �|l���)��%Q>vl?�Xf>31s>�s3�h]8�c�O�����|>�e5?]��R�9��,v��DH��ܾ8�L>�ҽ>��R�V�����up��i�aov=h?;?��?FX��yA��5u�O���]Q>6]>p0=AΨ=��K>��Y���ƽUUE���3=���='�_>��>:�b>mA=:�>�ٜ���{��Ü>��N>1.�=�*?�?����
�( ���½	}>]Y�>��>�>aDO�~��=	�?�� >��	��Žжν`T��	b>�U�Y���>g���=w�b$�=A!=��Խ����Uq=�a�?�s��ߚ�wٽ�Q+��O:?�?��L>��=�U�A����Ǿ*z�?�@R�?�q��ZT���&?��o?�$����=eN�>�o�>L�J��)˼o��>�3������k�=<M�?��?�-O�kը��[��Y�>y�?qlJ�Th�>px��Z�������u��#=P��>�8H?�V����O�M>��v
?�?�^�ߩ����ȿ3|v����>W�?���?f�m��A���@����>5��?�gY?soi>�g۾;`Z����>ѻ@?�R?�>�9���'�}�?�޶?կ�?�[>0H�?Ms?}��>��(>��������|��*>Y�� �">Ubx=v����V�8Q��6Z����}���,��o>C��	�>j L�r����">�ϽW�������2�>:�>�Pq>��>{?�!�>0��>��=1(C���?�|}����K?e��?5���0n�W{�<|��=[�^��#?�H4?��[��Ͼ�ը>�\?��?6[?�`�>���=��迿9������<\�K>K1�>8I�>����LK>��Ծ�/D��n�>�͗>&���Aھ1��?O��?�>2d!?͐�>߾�=� ?��#?rvj>��>�RE�H/��E�E����>ݝ�>�C?`�~?�?"ɹ��[3�\���桿m�[��4N>2y?nK?Fĕ>F���N~���tE�J�J�����旂?:gg?Y����?)�?�??G�A?�e>%��+ؾ�᭽��>�!?5	�Z�A��5&�����k?r@?��>�����ֽs�ڼ;��)r��N�?�#\?�D&?nu�(�`��%þ>�<��%���Y���;ou@�.�>�W>GӇ�'�=�z>;�=�<m��}6���a<[̻=���>��=�7�v����,?n�9�����D�=��r��yD�wr>qL>�$��_^?hN=���{�c���^����S�r�?Ռ�?�c�?N��}h�*=?��?p�?�>����޾7�߾��v��x�Ӛ�R�>Q	�>)���� ��|��bt������OŽ����z�>(ֆ>�/�>�?]>VG>�签�ݾ������0��&6�a!�4�9�g=���)�Eɾ^r(��0��jԾ�ۏ����>�S>����>u ?兆>1�>� �> �N=��m>�X�=�2�=M]>��>͋/>��">ռ����"�T�Y?Ce�_>�A�B�վ~�@?�d?�d >�h��uQ��0ǾSqi?s�?�\�?�Y>�yR����0�>��>JƮ��%?J�<��<-8�=0���I	��m�е�=ٯ�>sQ���:��<��}��/M?�?7�n�Q`	��=.=�S��7�^=fZ�?��(?*�NS�9�m�wW��S���V�f�u���]M$�_�n�����қ��^p���(�!�+=RQ*?�r�?�	�3������qj�L�@���m>2��>%ؕ>W�>3�F>ۏ	�p1�Ly\��?&�U���0��>�^z?�>�>"J?��<??N?/#N?��>�Ʃ>���,�>�};\��>��>г7?�*?�/? l?|H)?��e>���'���<nؾ��?h?��?��?7?����dν�����9�2({�������=C �<a4ؽ都�U=NM>��$?������7�'���>M�b?.l�>q?����~����Ӏ>Mt?�Q�>�h>���Z�y���޾˺�>)�?�]������;>6=�*o=�W��V]�=���=��= ���W�Vb>��/>��2=�4<�	r��c�.�"�!?��?{�>l�m>����������� >��u>��~>F38>8ξ ��� ����hf�ކ�>���?�#�?R{=�>h��=����ξ�q � >��q�
<$?8�?�V?)�?@�<?j|)?�A>�g�zޓ�C"��l����:?�!,?`��>���y�ʾ��3���?I^?�:a�����9)���¾��Խ\�>�^/�C1~�����D�ڂ�"��Yk�����?!��?�?A���6�8{�5���zZ���C?[�>�L�>[�>�)���g��#��/;>�|�>}	R?��>�oO?��z?�[?��O>(48�o���~���r����>U�>?��?��?��y?�$�>~>,� �mU޾�����G!����fŅ���Z=�X>��>D�>�F�>�#�=vHн������=��Ř=X�c>�v�>�s�>υ�>=�r>�4�<=�C?��>L�˾[E�@;߾)�O�tR�;�i|?ڦ�?��;?�!>O2��h�iz��/�>p�?c>�?�^?������b>�Խz��Q����ҥ>�F�>��>�7�>��>���>��? 3�>����]�"��U����xƴ>�/]?�Ψ��տ��{� �>�{->?yf���!�H!�=I-�h氾_,�>����7Β���!P���	O����ؾS*����L�?�&�b4>{��=`�)=�#��E>�QQ=塛�K���g�H��"�9/8��
>�(�G�z�=��p=MV�ؑھ��?o�h?���>}i�?g.>���3Z�<āW?U��<?���=tU<���O&@=.O���#;5��p�c{^��@����m=���~J���V>qc�>�R#�	��=���;E>�+��K!=�Bf><�=��,>��x>2��>�v�<�5v?[��������\P�o� �g�8?��>��=~
ɾ�@?�7>F����j���
�R�?�(�?Tz�?�?bk��}�>Nݧ�&櫽�L�=����Q:>$l�=�F0�/b�>�A>���z���a��֗�?T�@=�@?X^��[WϿ��->щ7>hE>:�R���/��Y��b�=Y�X�?�:��@;�I�>X��= Q߾��ž)�@=}9>�q=�q�f�[��ݓ=��}��C=�;a=W��>�D>�7�=.������=D�W=�l�=�tN>ѥŻ�J��;��2=���=��a>�">pv�>��?�W ?y�c?VB�=�՜��x�@�޾��0=S�V�XDl>��������> Y]? �J?2*�?�=�>xd.>O��>�LJ>�T<�� X���վ��j���>��?�N�?+m�>?��=���./�4�O�k��"�?�?ӆ?��r>�U����3Y&���.�D���~:6�y+=�mr��QU�����Mm�6�㽡�=�p�>���>��>,Ty>��9>��N>��>��>�6�<�p�=�⌻N��<E �����=@����<wżƘ���v&�+�+�����P�;ȭ�;)�]<���;��=�f�>��>=��>lÛ=�m����+>1엾��K��q�=�䩾 .A�Y�b�_}�K'.���7���>>�W>Mh��-��Ζ?�Z>�I?>G5�?"�t?�">��	���Ҿ
�Th�KW����=`�>�?��d;���_��M�1�Ӿ`A�>�f�> ;�>u�9>��q�-�Nt��x����$�w��>���8] <"���,�s���������v�W��0V?���4L>�*�?a�`?��?�ڻ>H���3[��<�v>ft���S�<ȋ%���������? ?��?���R��Uξ��ν��>�B��Q������.��cݻ�﻾7�>7[��&�Ҿ��1�@����ꎿ?]>�4�k�S��>}�L?�`�?�]�s!��z�N����6�l�͵�>8�j?p��>t�?�8 ?����¿������=�o?�P�?�a�?/�>��=�ԭ��w�>��	?�S�?uq�?�r?N�E�G��>>��;�= >���[��=��>
�=�(�=�r?w�
?�+	?�M���Q
�#c�)�͆a��=���=
n�>���>��u>x&�=�me=^��=�Y>���>�׏>��d>@3�>���>���-=Ҿ�q6?W�>���>��0?�b�>�T�Ej*>�+�=+��(�{��j�{�ίe�9z?�]���u=.v����>�N����?p��>�Q�G��>�骾l��dc>T�>O�)�(Fe>�}˻��>>_�>a�>;?>H��>��>�K����=���R��U>�b�T�⯾�}r>yϝ�'����y��tX���z�ٱ^��F~��dG�oV����?���
�j����jG�\?��>��$?������B2>���>}��>�=��8��Ն�¢Ӿ@�?d�?��m> ��>^�P?He?%_���a�CKH��3{��I��l�u�Y�K ��@�W��\��ҿ�=QV?Iw?��E?�=yV>9��?O�+�ن��K�<=�V&������:���=^�����'�ž���7=�k�>0 Y?��?���>�kW��4����>>�~<?��*?u�y?@�2?l�8?-"��g-?��">L�?�?�2?��&?2�
?�+>��=��h;9�&=����
���l��9���w����=�)�=IM�j���\=�r�<���������<)���#Y�<��<D��=���=hB�>@�D?c�b>	~�>��?��P���2�كȾ!��>kJӽb��]���4(�r渾��>~�{?��?�Y?3|�=k;������qD>.v�>��=��@>��8>Rʽ�Hg�b��=��I>+>�c�;�����������z��j���0�n>�q�>�\>��&�m�B>Vn�`jp��>VY��;G���́�Ɖ]��2���;Ƚ>�3C?Sb?%��<5������O6g�I�!?'?2�A?�Mv?��=�T��M#���@��00>]��]7����Bo��б;�#1���L>$ڹ����	>���/�������VOT�r澔�
=Xx�Ui'>��� )���w�/� >_��=1�۾�>����ã��q]?��A=��־��$>��_S>&�>s��>�Uҽ�a���<��z����<�װ>�2=>�&ŽD���L�T���=�>_OE?>V_?Bj�?i���s�T�B����mg��^ȼl�?#y�>Xf?P B>��=����	�k�d��G��>��>���o�G��>���)���$���>�8?��>k�?8�R?�
?�`?(*?F?�$�><2�����C?&?3��?��=V�ԽA�T���8�$F���>Xl)? �B�N��>Շ?'�?��&?��Q?k�?n�>� �g!@�ߐ�>�J�>Y�W�}[����_>\�J?Ό�>2FY?�Ѓ?'�=>ju5�W袾[d��5��=�'>E�2?�,#?��?=��>*��>w�����}=���>�b?�X�?\�o?.^�=�!?1�2>�(�><��=K�>��>��?cYO?��s? �J?�T�>�A�<k��7ڶ�A x���Z��6o;��L<l�y=�T	�U�u�[4���<�ջ;�Ƽ��c��
P��l)C��?��NI�;޿�>:�(>k���&2������{�K\=�"��o���Gڽ��9��>%p�>,�>�g>�ũ��$=�L�>�)|>�Q2�V?�e�>l?t��=M�h�A\�JD;�Es>���>\X���!��|Ҁ�o�7�>t&]?�`?��l=&���W�b?��]?j�5=���þ��b�j����O?��
?��G��>?�~?��q?9��>}�e�I9n����Db���j�kǶ=ou�>�W���d��>�>͙7?�J�>��b>�%�=�t۾�w��s���?��?��?���?o,*>�n��3�Tu�6l��\?!
�>�iZ��?��U=����=�_��_���)��1⼾����������'m�썾?.��x�<��?��W?5]w?�9_?]���&J���Y�9����'b������&�"�A�ũB��?���p��l������ό��@=�%O�xG6��/�?�?�&P����=�Ұ��;=��Q���=�֯���<M�>��7=���;t�L>������N=�EG��?��[>���>Z$O?�y�h�R���/�xeC�w!�--�>OS>#Z�>@
!?{�|>��>!O�=�v���L�'">�v>Дc?dK?n�n?�� ��1��~��#a!��-��^����B>>m{�>8nX����6Y&�AI>�~�r���������	��=l�2?�1�>���>�>�?��?�a	�󶯾�x���1��<s�>i?��>���>��Ͻ�� ����>C�m?L��>V�>F��* ���{�E��e3�>iʭ>���>v�m>+P.�M�\����	��T8�r��=�g?If���_���>�Q?O�;u�k<�>eBs�` �.���c�,�,w>t<?ӥ=��<>;ž���
'{�ړ��'�)?	?�A���*�7P�>��#?ɥ�>d2�>(̄?�c�>l1�������?��\?�;J?�:B?�i�>֣=�赽ǽq�&�7]4=�%�>�[>�^�=��=���3c]�`�!�1Y=y�=Iͼ�������:EҼ�"�<��<�7>����N��{����{���������޽r���1=p:ľ�;���i�H���B8ʽJnz�{�������ҁ�l �?�Z�?7g���ٽ�(��׿���龯�>�F��`�?���ؾ��?��ʜ��BվM���Ԃ.���c��o��UW�P�'?�����ǿ򰡿�:ܾ4! ?�A ?6�y?��7�"���8�� >�C�<�,����뾬����ο<�����^?���>��/��m��>᥂>�X>�Hq>����螾C1�<��?7�-?��>��r�0�ɿa���t¤<���?/�@��[?z)S��S'�l�Q=��?�?� !?o��z������p?��?�Ͷ?0q�>�Nl���Z��ǐ?:/��<��@�켹g�>�MI>B���h�^�i�>�y�>U����!����>p��>l�?'m��O�N�����>G�8>��ƾ���;BՄ?�z\�cf�5�/��T��(Y>��T?J+�>PD�=�,?q6H�2}Ͽ<�\�?*a?�0�?���?��(?#ܿ��ך>	�ܾ��M?�C6?���>[d&���t�t��=H�Ґ��@���%V����=��>C�>�,���6�O�zP��+��=���ƿ��$��v��K =�	�f#\���&����R�|*���o�Lz���h='�=�ZQ>$D�>I�V>�Z>�tW?��k?�?�>��>��佬���ξ����t��
���ҋ���5�IB��߾��	�������9�ɾ�g=�=��=��Q�v��| !�v�b� �F�f�.?�b#>`ʾR�M��#<�Jʾ�w������O����̾H�1�Wn�pٟ?i�A?����FxV����G��򤸽ɘW?���������a��=%�����=f�>3��=�1�03��TS��%?|	?/q���9Q>	�}�<+�?r�>e?�ȱq>�&?q�>�S��M�1>�>�~�>C[?z�l=.���NĽ߆?_W?�&������o�>����p��b��6(�<0��0���*�>^G��/���lU:� ��=t1W?Y��>F*��!��M��y��y�==�x?n�?�7�>��k?J�B?�̠<����_�S�b�
�C�y=��W?�i?�Y>�����Ͼ����\�5?�`e?�O>��g�+���.��3��?�n?�%?eޡ�^l}�������Rg6?pz?hD�aZ���|�MoY���>�U�>��>�g%�f�>�V?�e
�t���
%2�T�?� @���?y�O=丳���G>��?o� ?��{���&��}!(�:ӝ�eK�>e剾��Y�d�𾵜�s?@3W?���>�#'��Ͼ���=Oٕ��Z�?g�?����Eg<)���l�_n��E}�<)ϫ=��-G"������7���ƾ��
�����%⿼ۥ�>.Z@eT轁*�>�C8�/6�TϿ(��"\о�Sq�=�?��>��Ƚ����(�j��Pu�C�G��H�����V�>���CT�=
Ņ�����ϸ3��	r�4�?��D���>����6����ƹ��7X>�? #?g��>t�m��x��B��?zN ���ſ�v��Es�Q�R?���?�&�?%�@?O��;fu�z�>�0���A]F?���?�;=?W?V�'E�"j����j?Ȧ��^=`���4��E��PX>	(3?���>=-��=��>PG�>6�>�/�@WĿ�O��\���0�?x9�?���*�>�E�?q�+?�}�J����Ω��m)�ׄF�HA?��1>������ �E3=�#���R�	?>20??>�n�߹[?�v�h_\��:�������`>�跼�;��k$f�a7y�Z
��k=���?���?�m�?Tu��� �0D&?t��>��ؾ.>���F=���>V?c9�>����o�>GjQ��`B���>U��?��?�k�>������ٯ>�w?&Z�>.��?P�=l ?e?>�瑾�~���Yg>��>>l@�Z?�u5?ɖ�>��4�9dW��eA��5��&K��$��U�I�s�>��^?P�:?���>�� ����X���+Q����X���x�%s��8S��F>*6>Ϊ�=�k�w����?"p���ؿj���m'�U54?��>��?���ߴt�^���;_?`z�>�6��+���%���B�9��?UG�?(�?�׾DC̼p>�>�H�>�ս���������7> �B?"�_D����o���>���?�@�ծ?�i��	?���P��ja~�ւ��7����=��7?z0��z>���>�=�nv�ɻ��B�s����>�B�?�{�?���>�l?e�o��B���1= M�>��k?ts?y�o�����B>}�?��������K��f?�
@wu@j�^?	�@�ޘ�������5ȼ��=��	>V�	��,n=��>�/�|�(�B)�=3o�>`�!>��@>">m� >c_�=�[��œ!�˒��D����d�?�7�K}���R��.$���ɽ��L�޾H�о����k�#����x���"�L��I{�^�=,�U?qR?M�o?J� ?�w���>�i��//=<r#�6��=W�>[D2?L?9�*?�U�=���I�d��V��E9��FǇ����>��I>Qt�>F�>?)�>�g�>+I>�>>JG�>�� >�&=���\�	=6rN>�=�>���>\g�>lk<>ϊ>˴��/��~�h���v���˽��?HV��ڮJ�,��Y��ټ��$W�=q.?,�>w��8п|i5H?C���-�|�+�3>��0?�mW?۹>ΰ�$�S��V>Q����j��>E �uLl�U�)��RQ>;K?~�f>jBt>��3�f�8���O�|��^~>5�5?A#����9��yu��CH���ܾ�DL>[��>�"Z��H�F�����~���h���t=��:?�?Z��4���sKv�{��S>C$\>z�=Mө=��K>#s]��>ǽ-^E�-=z��=�_>��?�E,>�v=���>����N�K�璨>��=>�p,>
=?��"?���7x��R���K�/��0q>N��>1�>��>�K��b�=;^�>�oa>�μ}�R���C�3S>.f���'^���|���k=W��g�=U9�=�#����6��j2=���?8#���i��(���a'���1?/�)?�&l>�TW=�r�邫��a��U�?h@�ɑ?�t��d�&^j?`�x?a�<�2�=i3>$��>]���5#���>A�P�N���I�b�(>���?�5�?��Gc���l��59�>��?�fE�Ph�>{x��Z�������u�y�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?roi>�g۾;`Z����>һ@?�R?�>�9�~�'���?�޶?֯�?n]G>���?cs?���>A�m���.�ӳ��n��o�=�@;'A�>��>\0��`sF�����O\����j��s��a>�s$=d0�>���Z޼�~�=Cl���m���df��ܷ>}/r>emI>�N�>�� ?���>ә>�=�&�����閾	�K?��?A��C5n��.�<활=�^��#?G4?��Z���Ͼ�ܨ>�\?T��?�[?Ud�>���O<��@翿�����2�<��K>�7�>K�>--���EK>��Ծ�5D��g�>�ȗ>ƌ���?ھ2��Fᢻ�@�>ff!?&��>8Ǯ=ٙ ?Ӝ#?��j>�(�>9aE��9��8�E�9��>���>"I?;�~?��?�Թ��Z3�����桿b�[�	<N>��x?�U?J˕>T�����^VE�DI�k���%��?�tg?(S��?#2�?��??Q�A?�)f>����ؾȫ����>t�%?����E<�g������4�?ǉ�>A;�>�;<��������
�I��f�?��a?|�3?W����a�����'�<V!��}F9=�<�Y;A�Q>]�>b�����=Zl>���=&�X�2G��`�<�.�=%xt>�O�=
I��j���4?L~�=����c��=�Wh��R��7�>�j�>����W�d?� �=��O�<r���"���簾P�\?�?��?��8=�tq�$�{?j�^?ny6?ܯ�>q�-�L���n9��,:�[2���K���=I�>q�=�1ɾ�L��1|����Vֈ��*�U�?��>���>@�?�RO>,۩>e�t���޾[ �BVվ��J��_	��k;����=-�'��Z�
��^ԽTƾDX¾U�>'77��ݽ>|��>��P>GZA>�B�>�T=/;`>���=J�	>䠻>�R]>U�u>��=���c w�l5\?.޾P@���#�C����N?��k?R��>��+C��:����y?}�?-]�??�=��U��<#����>\�>rÝ�s�*?�8����N�������a��*�[)�=qa�>M`��9���N��W<�!{?I,?��)�0Л�!'�=���N^]=�"�?�*?*���Q�8on��jW�Y`S�)
��j�~t��ʓ$���o�n���E���Y���!)��z#=.�*?�P�?4��[��C��Оj��j>�\�b>�`�>�-�>�4�>��K>1	�F1��^�g&��ʁ��e�>8�z?Ĉ>�!J?[�:?iL?�^L?���>���>�!���z�>���;���>}��>��6?�-+?p�.?��?��(?E�\>�#������3׾\D?Ȥ?I�?%�?�C?�9���M߽x �bs��t�~��ݎ�!�=cI<�$콍zl�>[S=3rQ>/�?!C�ol8���tŊ>O@.?y�>?%�>1?���P���ƨ����>��?|��>�k �P�k�j�
��>�>�&q?zR�s�;��u>�2=b�=�0��7!=����=JWͻ��t&<�-�=���=���S	�=>�<��B<y�=�?L?��>�!�>H����s��?�
���=z�U>�tV>��)>}�־g��ku����g��>{>�?Af�?t�z=��=`�>��.����q�\<ɾ&�<(�?�>?��S?C�?"R<?D�$?jC�=�����������럾�?N!,?Ɗ�>}��t�ʾH񨿚�3���?�Z?#<a�����;)�s�¾��Խs�>�[/��.~�����D��텻o��6~�� ��?ѿ�?wA�b�6��y�򿘿4\����C?�!�>>Y�>|�>��)���g��$��2;>F��>TR?��>F?z�Q?�YS?s�<B�Q��"��O���`^��~0����>aTV?k�?;[�?�?�?��1��>ƾ�?>͘�����'7��0�	j>�V�>K,�>F�"?m�=��2�����e����>��>�ϳ>�D>=�+<TŃ> s?H�f>������.!��?�榽�$a?Z��?)�S?6�>h�&���o����h?w�?%�?���><p���!�=1ȧ�y+��ʓ��]Ė>aE�>!"�>Y}�����ُ>��?W�>}�D�!�� zR���E����>k�2?*�E=h`���I����>@��>��澅�3���=X�����	��4\>S��}/���q��V,ֽd$9�G����+�bo��G��XJ?���S p>��ǹ�B-=o���=�����n�=�H$��p��I�=(���&�;�(�Ab�>Q�}>�}>�_�<�f���o�?��?�>��~?�+�>�f<;M6���%?2L9�or?�Q�2�վ5<*�����;��L�8�*�tF��l�~�:˹�wY�>'��]�A��}=ح5>G�E�u��=�]�=.#$=	�<�O�=��N>���=��F>ϊ�<��=5q�=/7w?k�������_3Q��P�4�:?@3�>���=uwƾu@?��>>�2������vb�//?���?�S�?��? {i��d�>������oy�=P���K2>���=��2�㤹>y�J>)���I����� 3�?h�@��??P���v�Ͽ�^/>�8>��=_ U��6���,�U�W�/��u?�_1�x�;Ti>��=�ɾ7�žBK�<˪>��6=M$�[ X�%�t=�h�����=��<u��>e�8>>��=�ئ��^�=O�?=O��=l(>�����ʼ�S�$JU=«�=��E>�:0>���>�$?��)?�Z?C��>|Nv�#�$�{֥� ��=��B��'>�Q�=�	>�-�>*qU?]�R?ȇJ?�ad>��>雹>L�>�0/�j�Q�1*��|�>�fd;r8�?�{�?���>�8\<��[��6���#�}��<�h?�?pٺ>��R>�U����,Y&���.�d���!�6��+=�mr��QU�Y���Fm���㽷�=�p�>���>��>CTy>�9>��N>��>��>Y6�<Gp�=ጻ���<m��ȴ�=����a�<�vż����nq&��+�5�����;���;N�]<S��;�j>�?D�};h�>��=!���͗=�սN�$�pQ{>�׽���W)N����?�0�޵�X8>-{z>�g<����8(?�$>�RM>]��?()a?���<��q��^����D��M#`�f��<��=���<��[���`�&2⾸��>�ȏ>�>�Zm>��+�C�>��t=+��E�4�e��>]2��0��eU�MLq�k"��T�����h�4�`��~D?B_��+��=�}?�I?���?�f�>N��ؾ4�1>����y =���SWq�*n��Q�?Yu&?��>2��f�D��h̾�����C�>�bH�SP��Ǖ��|0�[d&�"��\ͱ>�����о��2��B��}􏿡LB��q�9ú>�O?u�?�9b��=��AXO���n(���8?x�g?џ>�J?�&?�ϡ��+�+��k�=2�n?��?\�?_>[ض=lq��v�>�?���?���?or?�A����>�6%;y >m�����=�>�	�=�3�=<	?�r	?G	?;O���
�jq�p��.U���<�=���>=�>��s>!��=ɮu=�=�)a>zŠ>&�>J�g>�ţ>!��>c&������M%?���=��z>��?�F�>;L�f�ƽU�A<׮��x�2�&���o����=�݅=��0��T=NC=��G�>p&�����?�-G>&����	�>�t��ٹ��d5>L�^>yG���1�>ܬh>r�>M5�>� �>�Ce>e��>�5>L�Ծ��>�c��� �
�C��R���Ѿ(�y> �����#�k������oFI�ⴾ�o��+j�g~����=�E�<�W�?R����l���(�L����?�>��5?����E���1>yu�>_�>)l���E��'�����ᾖ��?\��?`�e>F�>�R?�e?��,�7��|\�v�t���=���d��w^�5?����z�X��台�e^?��w?$�D?9
�<@�{>��{?����u��Ru>;:2��A����r��>0����Sc�F�ľ5Ʒ������H`>U�q?g�? )?b�A�h�n�cr'>�:?��1?dTt?%�1?��;?��q�$?iS3>�H?�\?G05?~�.?��
?[�1>޵�=R���@�'=�A���芾"�нtʽ���4= |=�&4�V�<��=^s�<!����ټ�,";/y���A�<�&:=��= �=Ò�>�TP?�s�>���>̪/?�B�=p��t����>3������c0V��Ӕ��Zʾ��>�a?S�?u�d?�6�>�K���Q�ġ2>�Y�>;�*>�%>�v5=�����k�����>��t>s�:��7��ä�����X�����eX>:��>�v>������)>����Ho�IE�<;G����ݾFe�%�^�>��ΨB�p��>e?�#.?H�s=�ޥ��W+>�[��U?CM?f#?Jyg?��=;־&�g&�����˖>xۿ�,7 �Wn��ဏ�kVJ�>>*p�>�ʾu��ܱ�=��ܾ��Z�G����W�c�#��<m�.���>!� =����T��O�=ଟ=#�ľl;��������?p��ξ�v�C�����=���>�>�>Ņ�4eԽ�T���վ�ʽu��>[��=�댽Wz�q�H�q��WL�>�?E?�=_?VZ�?����s�_�B����L���:sż�?g��>��?fB>p �=ˋ��B��d�>G���>=��>����G�W+��c����$�z+�>,?!�>(�?ާR?��
?#�`?w"*?AH??�>Pѷ��ø��A&?͈�?��=�Խ��T�� 9��F�{��>��)?�B�ܹ�>Ɋ?�?��&?�Q?t�?v�>� �+C@�В�>�Y�>E�W��b��Z�_>H�J?���>�;Y?tԃ?S�=>̅5��뢾�٩�gW�=>*�2?�5#?@�?}��>ϩ�>����C4�=��>M�b?�,�?L�o?�J�=n�?=Y2>���>ݨ�=B��>�{�>4?�`O?��s?��J?2��>z��<��(%��m�s�D�P����;[�I<��y=P���s�f��A�<Z@�;�����3�����DD�5+�����;r��>f�&>�����\'��Ӕ��M�p��p��>��8(�[��\�>"��>��+?r��>[ࢽ0�=u��>�?�c$�T�!?+s�>H��>��=�5��f�~�/��i�>x�?���m���ܓ�L{v�Ј6=�X?�j<?"P:='�Y�ձe?hnU?�K�/�6�hT����G��1��6i?��?��o��N�>VO�?��k?k�>H둾;x�,���W���νP@Y<Ȁ�>���r�U���>e�?H��>�B>�"R��R*�a�`����>�>��?;�?s�?v�1>��m��ܿWi�Tȑ�*�]?q�>�ʬ�jN?V쨼��Ͼ'����������k1��Aqꦾ]�%��·�������=nx?��l?��l?�N`?���@�d���[�>}�s�V�R�����EG���E���A���m���d���ʝ��a-=eHD��%"��?�?'��>n�򽋝�>�Ǿ S1��	�+o�=�f׾�dk�$�#>M>�S>�qP>��1L����ҽ��?a�s>�L�>0�x?��s���'�)-���8�rB1� ";`�>���>��>�b}>�P=�6`=�Wt�����#�k7v>�wc?s�K?��n?*p��*1�چ����!��/��e����B>i>Ѽ�>��W�x��q8&�6X>��r���Lu��}�	�1�~=��2?$%�>���>RO�?�?+{	��k���lx�ن1�bz�<l0�> i?A�>y�>jнg� �j��>x�l?��>���>)Y��=U!���{�Ηʽ��>���>��>��o>�,�*\��f��p}��9����=��h?cz��Ώ`�u�>��Q?^U�:M�C<:>�>�v�e�!����c�'��?>f?���=��;>�|ž\)�B�{�����:'?]{?ʈ��r,�uр>$k?@R�>6��>B<�?m�>EǾ u����?��]?��I?�r@?�@�>f==V͙�D8Ľ�$���k=pj�>+�^>�ޅ=%��= ��_T�1���p7=���=�����\�o;�����G&<�N�<IF.>�lۿ�BK�y�پ�	����@
�ꈾ����[g������c��v���Xx�?��5
'�qV�k4c�:���Զl����?C<�?���J4��ͱ����X���+��>ŏq��u�����%)��������b!�G�O��#i��e�V�'?�����ǿ񰡿�:ܾ>! ?�A ?:�y?��@�"���8�_� >�C�<�-����뾮����ο?�����^?���>���/����>ߥ�>�X>�Hq>����螾�1�<��?0�-?��>��r�(�ɿ^������<���?-�@M�A?��(���6HM='x�>��?�C>�4�5��N�����>�g�?xh�?�a=u�V��m
��Od?莕;��F�Q�����=.�=@=;����B>3��>�#���D�^Uֽ��5>͠�>���=C�pJZ����<I*[>h�׽�Z��Մ?d|\�ff�>�/��S���S>|�T?�*�>=�=��,?;6H�'}Ͽ`�\��+a?r1�?���?v�(?*ܿ��ך>p�ܾK�M?-E6?���>�d&���t����=�{�����='V�1��=µ�>E�>��,����:�O��#��� �=i���=ƿ��$�N��m=��T��|b��%�:����KS�4���zp����%�k=RO�=�R>�>K�X>�\>�V?�k?:��>�S>?�߽����u�̾tj�m����|��틾~��k`��љ�7�߾g^	�������Eʾ<�=��F�=��Q��J���!���b���F��.?�_">"/ʾ��M�_�<�ʾ(�������*����̾��1�~bn��o�?�SA?}���5�V���j	������W?������s[��D��=�P��{*=��>]�=U��43�%iS��\0?�~?�ֿ������+>hQ����=��+?lm?V�a<�5�>�%?L%*�5�㽥3Z>�}2>�1�>\u�>�<>u`��@ٽ��?U�T?�`� ��Z��>Q~����z�m�]=�7>�?6����FY>�ё<,ƌ��sM��
��l*�<�G|?[�N>��)���R�2oe��Z?V�Z>��V?��0?&����W�?�a�?�i�=*�꾗,r�&?�m�$>�E?[;g?�">�O:�ɹ����F�u ?��P?g��b����T���	:�`����-&?��X?�D?�ʼ��h�"�����0�.D?�v?mr^��r�������V��;�>�]�>��>��9�o�>5�>?K#��G������`X4�HÞ?��@���?R�;<T�c��=9?�Y�>�O�=ƾ�q������ɕq=:"�>����4ev�c��R,�ǉ8?���?��>�����͞�=�֕��Z�?��?p�����f<z��l��m��Pn�<}ʫ=���Q"�^���7���ƾͻ
������������>�Y@?I�}%�>48��5��SϿ����Zо�Zq�]�?t��>âȽ����j�\Pu���G���H�����=��>�j><�)��b��U�e��M,���<#�?����Y�>�*�����־��ݽ�$->��>X��>!�>�w��.�?O��BҿC嚿��$�N:�?�å?�#q?Xe%?ܦ�=ī�<׃齢��=qB?� X?<2?��Q={�0��\ν�j?�?��f`��4��)E��U>53?�x�>�l-��2{=�b>6��>ԧ>�/�Z�Ŀ�ڶ�[���a�?ۄ�?�r�#�>ys�?�_+?S�-5���?��ü*��k��TA?�1>���B�!��=�`���f�
?�i0?���%B�-4]?�������kG%�]�(��{>}3�;����R�W{�=��=��!���Fq�.!�?�6@k�?|X,���(�=U�>�+�>�O���w^�Q��=M��>��>�z�>i6@�>�^$��<��M4>�1@	�?� �>B{��Q!��9�%>���?���>�?�?O��"(�>�*�>(����ㅽIR�>�g*>��4���?��?���>�V5��Ѡ��4���A�"+u�w7���E���>b5]?�\K?��1>��K��M������X��ᘾ��a�릊�2K���ھ+;>��>�*!>	�6�i�����?Lp�9�ؿ�i��p'��54?+��>�?����t�H���;_?Rz�>�6��+���%���B�_��?�G�?<�?��׾�R̼�><�>�I�>B�Խ����\�����7>/�B?b��D��r�o�{�>���?	�@�ծ?ji�?g�e���Gw�y��UhS�h�=6�??t��#�>���>kh=�)y��o��k��k�>��?[4�?���>��q?=uc��K�q��<(ڤ>6j?"�?��<@vо��W>��?��6��� ��?q?��	@�	@�]?9��ɲſ�胿�ݽk((�o��(��<E�ødm�����>�4[=�(�f�P>Qt>�+>�G>��>�'=(�4�������9��E�b�&�u�Z�6��8��G��.B�u�	����4񾄮��@�����9�9a�E˾�L��	�r���=U�U?�R?Kp?�� ?Ԛx���>������=�#�@��=�.�>�f2?��L?��*?j�=����d�A_���;���ʇ�E��>��I>Mr�>�E�>"�>��g9��I>l4?>y�>� > 	'=7�,V=��N>�L�>��>�q�>�C<>��>Fϴ��1��k�h��
w�q̽1�?����S�J��1���9��Ԧ���h�=Hb.?|>���?пf����2H?&���z)��+���>}�0?�cW?�>!��v�T�4:>9����j�5`>�+ �~l���)��%Q>wl?�f>ʬu>��3��J8�ԇP��=��k|>:6?�¶��D9�\�u�E�H��2ݾM�L>pu�>ξK��l�������W�i�)~=�t:?��?���:���Tv�`k���R>oS[>Ȕ=,�=d�L>xg�xƽ�H���-=���=�h^>�)?�
'>w��=m�>�=��2�=�L��>��*>��:>�]D?�Y?*B��C�Ľ錾I�<�PK�>Ҽ�>���>T� >&O�q8�=��>�y*>��輅崽���>��F2>��y��G0�.ʧ�(pt=�n����=k�<@�꽔+9��+�8��}?XZ�������)���R�g�F?5�Z?�M����>���x����>�����?@�ޙ?@L�C�K��o?[��?Kh弽�T>Pz?X>q��*�<8�>+�A�����;$,��ʂ��v�?抒?a��=�������wX>�9?Q������>?��8��5���u��a%=���>�9H?[����wO�O�;�ky
?�?!��I�����ȿ��u�3��>���?���?�m�OL���3@��\�>E��?:�Y?0�h>6�ھs�Y�Ʋ�>b�@?�YR?q��>C�0�(�4�?���?\��?g5>���?�v? �>�$]�q0�ׅ���m��w�=MF,��A�>!��=tO˾��K�o��������,e������O>�L.=W�>"6��/~þ�%>,���2���*9���>+rD>�@>�³>�~�>��>�<�>��=�×�&s�cm���K?�u�?S��n����<�*�=X@\��?�.3?��P�̾�O�>4�\?�t�?�@Y?�0�>T��F���6��@����J�<{\O>��>�U�>������I>7=־KG�I�>zK�>
%ռ�Xھ-��3�U����>�q!?�B�>_Ħ=8p!?�m#?��h>�ʭ>g�C�@퐿_�C�x@�>��>	?��?��?�;��T�3������
���W�[>�w?��?�v�>���O����Q޼}ɼ�:n�ڏ�?XLg?g�ڽ�?M��?2�A?77B?)Z^>���Ծ�?����|>&�!?��W�A��P&����%y?�I?���>�*����ս��ּ���u���?H&\?�>&?���;$a���¾��<�"���L�.�;uC�T�>��>�t�����=<>X��=Zdm�<R6���e<�P�=�{�>���=�27�𚎽+!?��<��߽�{/>�Do���,�6��>n��=Lڡ�;^?����� ��Λ��ъ�#̊?��??��?Sx޽@�d�4D?���?"/�>�c)??�辇#��vYȾڤ��7Ⱦ�l�hj�=7�> ��E�þ����ج���G�n��; ��� ?���>�>�>	+?���=<�>O���zU�����@����V��B�KW;�TC)��}��Ӣ�(����9Vv��;�L�nޠ>��ҽ�r�>�d�>�6/>i�>���>�h��`x>X�{>h9>�[�>�I>d� >���=U�W<���M�T?X�̾"�1�ۤ �ߐ��T&?S�i?H
s>�)L�q#2�-^��<�X?Z8�?�+�?�ye>@�V�:"�Z=�>���>\���?�L?ܓ">�((� �=t5&�d�Ⱦ4���EӲ���>���=�{�g�"�mYJ���>3�1?�;���󾌂,�V=���#R=�:�?�)?q�*�K�R��dn���V�u;S�f:�7\m��򢾫�$���o�/֏�����惿}�(�QA=��*?�Έ?�9 ��<�P���y�j�^?�b�_>�
�>DV�>ި�>��J>�9	�N1�8
]��%�L�bV�>�{?���>f<I?_�;?/cO?�OL?�ύ>�N�>�E����>3�;�q�>���>2_9?��-?H40?4_?u�*?k�d>����e��K�׾S�?W?y\?�W?�?-��W����ޗ���s��{�������=���</Tؽ�w���R=�hR>p�)?l|���H�0�����{>�O?)�>� ?����뿾��	>��?=7?l|o>�������R�>��?��j��L�=�%�=� =>�P<�d�#9�=��$=^�I=N�=��ɽՐ�0>��>�u�=�M�?\��3��\z��d?�*?6 �>���>������!E�&x�=��j>]e>��>�X۾��ҕ�,f��ď>Ӓ?���?K,�=oQ>��>���ɐվ���o��Yq=�?��?��P?k+�?!�7?i� ?dq�=$*�?��z�%��=V?�!,?0��>�����ʾ�憎N�3���?-U?�>a����5)�݁¾=�Խi�>uW/�4+~���|D� ���8��iW�����?p��?�A���6�I�辥����_���C?�>-Q�>}�>��)���g�� ��(;>V��>!R?��>EG?�{?:zX?��?>:7����+���m���v��=�C/? 'w?��?O�?ku�>>$@>}����Ծ��������H���A��~o>&!>��>�5�>��>b��=��ܽ�8Ƚ��%�o�D=�BU>_��>+ԧ>���>2P\>4r>��gF?���>G��m��y8��,aa��P^;`�d?%V�?�2?��9+���JG��p���>�Ы?j�?��*?ĩ��7�=�b=��!���Р>@��>(�>�X�=:�=\�#>6y�>�%�>������&7�00��w?)X6?6��=cSſN�p���>#(4>;Z'�b ��v[M�����f>����ݾQ�־T�\�=��"h)�(zо9�ؾ�����"?�"�<U>�>X�J����<�5�;1ބ�ԊL=X��<J��=5�<��=�=������m���#>`�>�9�>٬5>Y����0�?���>�-�>^��?� �>fj�<?�>��4?W�
�6g#?���>�ɮ��"�u���h���������b��)������">�\;�#>/�=�e!>\g<��$>:B<���<�)�=�o`=�!>."6>j�
>�7>�>u(D>ss`?�Ȃ�W����:�b�`�a�
?��>�i�>΂��>�t?��2>�����������?�2�?*$�?|	?�����=�>����	���b=$�|>7�>�-�<f���@�>O�Q> � ��8��᳽ƫ�?��@�u7?M_���Hҿ�!!<�@7>u>v�R�0�1�:�[���b��
[�aN!?�;�N,̾}΅>���=��޾�jƾ�/=�6>�a=���Y\����=sy��n@=i�k=!��>aD>��=�T��	��=�GI=qN�=]!O>-W����9��p-��3=u+�==ob>�z%>���>9I�>��B?ʐ?{�=�(��ħ��.�[Ҵ=I��=K��8�˽,��*��>��.?B�?q�Y?���>��l<�=�>�@Z>,2���������[���F}>��?���?0;#?R�=s�t��)��z�����H?T5?R��>21�>U�[��3X&��.�����Q�{���*=�rr�ESU������r�y���=|p�>���>(�>�Qy>C�9>��N>�>�>uw�<�k�=?g����<�씼���=.|��F"�<�}żȓ��e='�w�+������ȍ;ڟ�;~�]<<�;5�=aA�>�ow>���>h��=9H¾�A'>E1����=�
�=�䡾urH���b�"1���a/�ή!�8S>.T�>?��S���q�	?�D�>��=(�?VaN?E�<�M�diž����ی�$�὾G�=��>�23���J��y�Q�5�C���6��>K܎>m��>��l>�,��!?���w=U⾭d5�(�>�r���I�}���,q�H:���񟿆i�oܺ٘D?�E�����=�~?�I?;ߏ?�w�>�y��H�ؾV/0>1J����=(�!+q�/m����?�'?��>��ȷD�nǾ!����>��I��F8�(W��o�=�^�=��۾R)�>����Važm�K�"y��v�Y��b�D=��>c�!?<�?��,��y�h�B�����}>;L?V(�?v�>��?�3@?�};���M�~�ǡ�=vfK?~��?�4�?݊w=�S�=�˴��{�>v�?�?���?yEs?->@��a�>͝�;��>	�����=��>�˜=���=�T?"�
?!�
?B����	��-����MX^�3z�<؛�=�F�>��>Hfr>�O�=2�g=f��=t�\>��>��>}Le>��>V�>��%����/?�!��%�>�?�]P>K��ș���š<:��X��Y,�ҭ������eeM=�Ν�p
>q��=H=�>�0�����?��b>d���6
?���pq���=�7>����W�>L�R>��>��>Vq�>�C>���>y�)>�^Ӿ�f> ���W!�c0C�#�R���Ѿavz>����7�%���e����EI�Ak��ig�3	j��/��C=��z�<�E�?����8�k�0�)�����ې?�e�>F6?H֌�� ���>W��>r��>aD���dō��d���?#��?�~`>�_�>^�Z?2�?,����>�BX��Ks�N=��4c�x�`����Y�����Nkʽ�7]?��t?�C?���<^��>��|?ƃ$�1菾��>�?+�ϝ7��/�=)Y�>�ͬ��1R��%ɾH�ƾ����]=>E4l?sF�?"?fA���w�2�+>��:?D.1?��t?l�1?Ǌ;?*����$?Y�/>/�?�-?��4?��-?��
?o�.>���=�;ۻ#= ��U���ƐϽ=<ɽA��v4=(�{=������;�a=���<��ݼ�����9򩮼���<�;=�5�=�(�=Mo�>��X?e��>�o> X4?�a'�S7��຾W�+?}S=�u���������ݴ��E>��h?{ݧ?��Z?��>%C=�H�.�Y=>�	�>��4>ؘk>쑴>�:ʽ��'�6��=*>�%�=1=�D��26��|������_�<NJ>
��>B�{>xn����>����~��2[>>.\�r����XQ�|TH�6�1��Iq�D�>��K?J�?%w�=��㾬���d�:�(?��=?;cL?o?A�=4�׾��6��\F�g���e�>f�@<6�	�Vs���T��d9�m�����p>�㠾����F>I�����x�xLJ���Ծ�&�=?�
���C;�����8���� >�f>�㹾 $�Mg���򨿖$I?�@�=Xܟ��J��H��&��=�5�>��>=�d���C�;��~���Jt=i��>�)>����s���}H�T���r�>��C? W\?��?���Wrn�F�K�ޛ�P���=�<�?|�>�?��(>]M{=3���+*�t�`��SD�Y��>#6�>M���Z@��Ύ���k���m�> E?xM�=¨?wL??��?��^?/?̶?���>"*ǽ���.m&?0�?H2�= �Ž� X�!�8��;F��>Bp)?��B�<!�>��?7�?9�%?�Q?>�?߼>3� ���?���>�5�>�V�S8���]>n�H?���>Q�V?���?��4>�C6��䢾㨱���=E,>�3?� ?�?��>_��>�2����= v�>�q?ZM�?`�Z?vN>=$#?�/O>���>���=s6j>��?�#?ܡ[?�s?>E?W�>D?�<���;����~����ֻK��;��=����������=�#=Vɷ;1��<I�L=��L=�� ���=1�8=�m�>j�s>=땾�.1>��ľEX��Ʃ@>MO��;,��񓊾W&:�U�=lm�>�?�ҕ>��"��D�=1��>��>=��UJ(?��?|?T3;u�b���ھ�vK���>��A?�u�=P�l�nr����u�Y�h=.�m?��^?ctW�����>sb?	�]?(�𾐸;��ľ�~c�'e�V#O?ui
?�G�-�>��}?� q?j��>J�c��m���*>b��n��׶=��>�z�c��ޝ>�7?���>H�b>R�=t�۾�=x�d���0�?�w�?��?��?�(>B�n�CM߿��Ŧ��b]e?���>�U��t�?e^����ξz����Kk��I��ħ���0���料�d$��򀾺��hč=$�?Fu?��k?ad^?#)
�v�T�A]������X�w!�C�B�9��:�ҿ?�tUk��h��c��p���U��-�f���Y����??��>[�1��>ꣾ�1�~�ʾi̛>����+�y-���S�i�:�@Q<G�d�S~�Yž�x?oY�>�9�>X�B?,�v�R�B�:���C�<6��S<��4>�^�>���>6��oU������#ƾ�Ѓ�-�>A�Y?��@?VRW?l兾Z'�J3��p\	��*��g�X��Ҡ>�>��>�z-���ݽ�B�wHY��En��>�DRW�����b�
?�>���>Ћ?��?��R���оk���İ/�iO����>�z?8j?l�e>'�L�O��(��>�l? �>��>����^l!��O|�o�нO��>f�>�>�p>�,��\��P��#_��p{9����=I�g?������_��Ǆ>��Q?��M:n@<��>��l�b"���~%�BM>+�?�D�=��<>՜ľ���2{�!���;y1?R�?t]��;	�"�>ɑ?+��>p�>��?�5^>TG\���U>z?��T?I�H?��=?)��>z��=�ܽ�ϼ�L�2�q�=��>��[>o��=��=av�+�P��G&�6í<L�>p��<��=^ӿ<�Y��y�=w�=��=<�ؿ�V��V��?+�%	�/,����&������4E�1��=Ծb���i�ݽӄ;nh:�_���d���#<����?���?�ø�q� ���W�Iy���x�>���� �.����ZQI���������Ͼ�J?���(ƈ���X�,?��#��ȿ�ؔ�W,о�f?�m?��H?1?����U���ڼo/>w+�ǉ(�B�����Ϳ3�۾%|h?�}?��ξa�e�F�?I�>��>b�K>Q��(5̾]�5>-��>�K]?Y�Y?��4��SԿ�����u�=���?.�@�A?�(����"�V=���>ڎ	?/�?>\�0��-�M��4q�>O@�?&��?ʵM=W�W�!��;ve?H�<��F��޻���=TQ�=��=����J>79�>[v�=;A��ܽ��4>�߅>x�!��:���^�4[�<ۈ]>�qսZ���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=����;�ɿ���(��ߦ�<�؎��0<��I��_ӽE$��g��|��^��U&�=���=��h>V݁>�a>�J^>U?��q?��>|��=����.P��z��#"ϻ�n�����~���'��������
�B �l���)�>v��߹�
^\�0�5�S
_�Zt����8�L�Y�U$'�n�1?vv>[ �^�\�+�r�ɺ����a�I�;=m�r��P;g=�}c��g�?��G?V���]�$9&�Pս���<�3X?����~�
���̾�T5=��a���~1�>&V�<[y�\L���Z��c3?%�#?O8��̠���ZF>�Ľ��U=�4?Qg?>r¼	�>�2?�署�˽�8k>v�@>cA�>[��>� >6)������Z?��Q?����鉾�c|>�lľ��o�@�3=�	�=Ѕ0�'�ʼ���>y3a<ߊ���;W����r��R3^?���>N��&�Z�G��,��'�=$��?�?_c>�z?F�V?E�>a�����������>'�L?��e?;r >C�0��g��!���<�0?�w�?埿>��&���V*�����2?���?ܵ�>�!��Յ�U���R� 7?��v?�r^�zs�����`�V�p=�>�[�>���>��9��k�>�>?�#��G�����~Y4�Þ?��@���?��;<1 �_��=�;?i\�>�O��>ƾ{������d�q=�"�>􌧾}ev����R,�d�8?ܠ�?���>	���é�Yb�=
J����?f�s?� ����㼗t-�6�t�Y�侪�y=P�<�m<��㽄����u2�s��������P��Y�>��@]�G�1?Yj��.�Ϳ�cӿrS���!��Kj2��*?��> hռ�'��>�f�.m�+B��3N���l�dO�>h�>����%��{��o;�U��7�>�����>6�S�j%��8�����6<��>��>���>s)��lｾ���?�c���9ο����.����X?�c�?o�?'v?t:<L�v��u{�f���2G?Z�s?[Z?�x%�3$]�&�7�9�[?vcj����1@���R��W�>��'?��!>��,�m�>���:H?��
>�Wc��ÿ����F���(�?���?7��q]�>���?�!?������/��?<"��b�=Hu#?n)�>uB��aL���9�~b`��"?� ?O8���@�]�_?+�a�M�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�f6%?�>d����8Ǿ��<���>�(�>*N>^H_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?%D�>�
�?oI�=�V�>��=1���C�:�\#>;T�=E�>��?fqM?H&�>�q�=	m8���.�i{F�2XR��=���C��·>��a?OL?�wb>o����d/��� �sʽA�1�9��0�@��/�E�޽�;6>��>>�>�wE���Ҿ�?�r���lݿ�������@o?��>���>��2命� ���l?ߍ?-�/��Ƚ��Ś�*`���?��@+?�����>��=�+t>�2�����k�6��wV>\�>?$�U�	^���$��I�>�?�<@�$�?F�H��	?���P��2a~�ɂ�7����=��7?�/��z>���>�= ov�����-�s����>�B�?�{�?��>�l?��o���B��1=�M�>b�k?ns?�o��󾾲B>*�?�������K��f?��
@\u@)�^?�׿/U����ǾrZ�	@<���<&!�<�*���`I�o.�Vf����۽�~>yp�>K8z>M<�>z�>�m>��3>El������ʵ�������W���'�c�3�1�R|��p̾[�J����Ǿ�A�=�iN=�����4������7k�{N>�B7?��<?f	o?Y��>��߽ڿ='��b��=ԫ���=��>�r�>88?ly$?=��=^3���s�����Ғ��٧���>R�3>���>��>��>4����t
>��P>ʑu>���=,�����=�)]���=���>ӯ?�1�>���=q,�=�㴿�}��s�x�N����9�����?����@V��՗��]��1(��0�=�-?��>�ڐ���ѿ���� D?0������������=�O"?F?��=W@���*u��$&>��#��Jr�ь�=�
��0^��&�}�>>�Y?�Lһr��=��>��W��m�p�߾t�[>��/?P���v�����y��Y�<5ھD��>K�>��<"��ܛ�މ{���J���1F?��,?��=��{�
V��v���	&>�]>��>ͯ�=.E>\M7��4����F�=�4b>��>�?�#>&��=Ѩ>�ꌾ� T�=��> �>>p�4>��@?�g$?�弴4����a�i���>���>^�}>I��=0C��,�=��>A�_>��6��M�&x4�ٵH>������L�D�x��V�=�;��N��=���=V`ݽ�+�{:>=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾI��>�����+Y��_�b���=��>�/?N����?��+f?�!?�k���^���Wп��}����>� �?�?;g��y���V4�UW�>��?�K0?�+>#ﹾ�����i>x�X?�$U?�W�>�����g�?�$�?>5�?�e>g@�?�is?	�>]�m��,�����o��D��?j>��>W�y>K����}D��狿����@�u����^�=qa�=�T�>��v�-���&��;yѽ��H�`=��>{�r>��>�O]>��?d��>r%�>��=�X	� pj��b!�B[K?0 �?E��4g�kq<f�=,�c��4?Q�7?+~���̾��>�V?_�}?wH[?�)�>�K��霿����'D��*�;<A>)�>�7�>_����ZS>��۾ScD��Վ>��>k�$S���~�o��9���>�"?���>gx�=� ?��#?i�j>�0�>�fE��7���E����>Ј�>�R?4�~?c�?�ʹ�Z3�t��?㡿ۘ[�uN>��x?�R?�ɕ>ƍ���~����E�K[I�T�����?�^g?�m��	?)�?P�??N�A?w?f> o��ؾժ����>�"?��/�4�O��ߖ�,��>��>�q�>w�<�qLս����6�x���s?��[? �$?�����i�о���<���㈼�<��<�*>Ͳ*>��ͽ���=0e+>�4=�R~��Y�[=�<ȋ�=��>��=�D�aLf��+,?A!A�6M�����=��r�._D��>��J>�����^?I�=�N�{������1�U��֍?���?�x�?�����h��	=?�=�?5�?�/�>k��-�޾�b྽�v���x�L=��>}?�>Di����y���S����5���SȽ��`�VK�>�|�>+?�X?�6>��> ���O�.�����&�r��%���F�/H�d-�ug��������Wƾ�㳾�>�!4��-�>��>T�>���>���>�U>	C�>��(>�$�>�\�>O�w>��L>��>�V�=2Q7�LR?������'���簰��3B?zqd?�2�>!i�P��������?���?s�?,>v>~h� ,+��n?�=�>A���p
?hY:=���7�<�T������8��X��>5F׽� :�7M�pif�-j
?f/?	��ً̾l?׽x
��e�r=i�?�'?O*�?�O�9^w�@]�A�K�g����Gf�Dc��q%�vo��6������o���W�'��n<��(?��?"����Ӿ�޻��f�HlD��@A>jZ�>���>�3�>�Y>�d�i_0��)^��"����c��>�Iy?3�>��S?�f7?2�U?�V?(�?C^>l�q��?�hF����>_(?�Z?�1?�6?n�?8P:?zMj>��G���ݾ��پ]�?���>��>���>���>����' ����=d�����a����5>�W�<�O��T��=¿��;+�=�b?�
�Z�8�����3k>�~7?���>��>7���!G��	�<^V�>t�
?\.�>b���X^r��Q��d�>ܚ�?F
���=�)>��=n��7A�� #�=/���M��=�r��^<�~+$<WԿ=��=�����f�1�:�W�;@a�<.t�>��?���>5D�>@��� � ���f�=�Y>eS>w>1Fپ�}���$����g�\y>�w�?�z�?�f=x�=���=�|���U���������3��<��?QJ#?�XT?r��?��=?>j#?�>m*��L��t^�������?U!,?���>�����ʾ�񨿷�3�ޝ?'[?�<a����;)���¾s�Խ�>�[/�d/~����D�KՅ�������.��?߿�?(A�T�6�y�ο���[��e�C?	"�>�X�>:�>2�)�_�g�c%�u1;>���>HR?���>$�L?@�u?��W?e�#>��6�Ԧ���9����B���<>=C?�Xy?���?�}k?�>��>�1Y����,��ۊ�pD꽠 ���=��b>q�>�e�>�`�>#;�=W�	�$���@J�V.�=�~>]��>�#�>S"�>�-g>�)d;:[M?��	?ë���辒k��������%c�?�?$4?�1>�- �Z 5��ݾ�!�>���?�z�?q.?��� �=r~g=$<��V섾5��>���>x�>"�= �<w��=/��>��>� ����-���/�U��a��>N,?��<>W�ƿ��x�	�{�� ��jͼ�$��v�`�k����=U���*<�����F��ڲ��%�b���Z��:;��p袾:��>��<��0>J0&>�}�=�^�<"�<���I�"<�^�=��)�|�<��v��  ������R(97�=���=j��<�dɾ
�|?��H?��+?d�C?�v>ښ>�>�a��>�t}��Y?��S>��Z�z6���:�+T��B����;پ��ؾءc�O0���>=�Q��>&�2>S��=SG�<��=_[j=�
�=Ⱥ�b�=��=���=�4�=f8�=Ou>O>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>5�9>%�>��Q���/�S�X��Xc��Z��� ?n�9�խʾ�}�>��=P�W�ľb�2=�;6>��h=HT�I�\��/�=W����7=��c=�j�>��B>Wz�=�������=��J=T[�=AGQ>^���1#�4x*��&4=�p�=qOf>�M%>T+?�?�?H\`?���>����\U۾�Y#���>W��=�B�>/>�=���=Y��>3�K?a�\?�X?9��>���9ķ>�u?����G�F����꽐����?=gq?��=���=��t�������e�Ct0<!(?V�5?z�>ȱ�>�$�o��" �]������]żɚ�=vŪ��6���׽��I�:�i�}��<K��>���>cl�>g�}>�#>A�=>�s�>���=���=$�>��a=]��=P>� ����X���j>j4�;h��;�8˻�����4d���{�<4�=�K�=��=��>��>���>��=�/��7�>v/���VG���=����nSA�b|e�O�����5��]�� >X�r>��yz�� ��>��>��J>c~�?��r?�>�����־R�J8Z�|׌�C�=��0>��1�H:8��F[�.nP�xi�+�>�ԝ>�'K>�k>9+.�Z�>�)�S=��	�»(����>� ��a��[��������圿Y��{>/�L?:,����g=.g�?\4@?�S�?�r�>�"��>���**>I�����a=��8�	[��а�<�?3s?{u�>D��
Z���̾�s��Eз>,�G�M|O�G���o(0�{�
����)f�>2��$Ѿ-3��M������f�B��q��Ȼ>ekO?]��?��c�1񀿍gO�L��B�����?�Vg?�u�>��?Sf?hu���U��A]�=�o?Jf�?��?��>t>�����1�>j
?7�?#�?�-[?�����> a=�2>Ƿ���-�<��T>A�=<�=ѹ?� ?�/�>y���iv�V2־Ի���g?���<�=x��>��>��>sx�=[B$>���=�,�>�S�>$­>C�K>�Q�>�"�>Y�ɾK�.���*?�[ =�>�>xK�>��:>�>`fF=.�>S��=�=���&�����8�%�L��<�L�=���>&�=�3�>z����o�?��q�b�!��>�	�	Y�1W�>/�>�^S����>ba�<���>� ?Z��>�P�=C�>�2>,�>�z�<�٦P���4�
J�^>;�þ-�v��M%�bh�����`uӾ���lj�oύ��[���<�Z�?���<A5����K��>��> 8?�#���ٱ�h�=_��>��>p��S���G���M9ؾc�p?x��?sCc>�>��W?Q�?S�1��3��rZ���u��$A�e�ʶ`�a��������
�;����_?��x?"rA?�<�3z>���?��%�Dӏ�Z.�>�/�B$;��c<=�(�>�'����`�%�Ӿ��þ�*� 7F>ҏo?
&�?P\?�UV���>�v�> uG?�P:?J=q?��F?�\?ܨ�=��G?���=�?ӌ?�i@?R93?�f#?�~�>6�>�<��v�������љ�����Z��Ê<���<�_=��9;+(�=��W=�� <���;�Q`�%�ϒ�;��!=L�=��=�>�_?�n�>̉>fZ6?�8&�7�W&��~�/?�'=��n����k2���'���>��l?Sƫ?�lX?�|e>�<=�31:�>L��>y�&>�Mp>=#�>�罧xI��߀=��>�j*>t��=�⃽�ʅ�<�
��ǒ���<��$>y��>X�v>Yk\��bO>�z��K�r�U>}�u��C��$-�SY>��2��d��d��>�'J?S,?��O=�����_ֽ��\��}?��/?��I?΀?�sv=�̾L�:���P�����c�>���<�H	�ﳛ��M���<�M�= ��>񩝾�g��2LO>"V�$�߾�k��sB�ưվ��[=����B=ޡ��<��Ԁ���=�}>��t �sF��c4��SwJ?�[�=F��<�o��F���!>���>V�>�Ǎ��Ø�	�>�������=÷�>_�4>������[J�c@�1��>;<?�kX?�%�?0�\�c�d�:4>��kﾑ��O_*�F�?lH�>9 ?C�}>kz�=����?�	�-�\���F�v��>���>"���uM�����3����}�?��>�?�C�=��>�A?��?̩e?�1?�
?��f>o/��0L����2?Bc�?Ѿ";2b;�+ D���E�h�=���;?֊C?H!���G�>���>���>ʺG?d�s?ن'?-�;>߫��DR����>�r�>��e����P��=wf
?e�i>�y?�M�?%�h>�=*�&��,Y��r��=>�Y.?�]5?��?=z�>�`A?�����0>��7?�a{?���?G�%?���>T�?tU�>��?�b+>0Ў>��?�+ ?��G?���?Y?�{>�f=;�<����>�=x =��<@���/^>�u>�q:�T���a4=�� >ၽ��8�FOԽ��=�=s��_�>n�s>�	����0>_�ľhO����@>�y���O��U܊���:�[޷={��>,�?���>�W#�ܳ�=���>fH�>���6(?k�??{;!;<�b�2�ھ��K���>,B?���=��l�,����u��h=��m?a�^?8�W��'��-�b?<�]?iX��=�+�þ��b����f�O?��
?��G�!�>��~?��q?I��>N�e�<-n����>b�C�j�w��=�v�>�Z���d�r+�>)�7?K�>c>};�=�۾O�w�*p���?��?
�?7��?.*>6�n�%-��(�����V `?���>s՝�iQ?�ɻ�Ҿ_����3��Z}޾�����G��U݌�6��|{���4��<�=/O?dr?Z�q?��b?����0e��r`����'�U��d�����C�`�F��.D�7�p�����=������ֆ=`����X�FĶ?q��>�F.<��>��{��󨘾d��=|�������<�=3��=N�X=�v>G�>��,L�㭳�.�?V �>�w�>��P?V�c���O��D�?��c�b>�h�>s�>�T�>us3����=�nV�rKV�`w�一>&%Z?��L?�~k?*�D��8D��쇿�n+�/G*�2HT�d�R>�H2>�]�=
)^�����a`��,D��Mm�g���y��Y7����-�?�f�>ӛ�>���?���>e�ʾSH��[���*��]=R1�>%�f?@	?�ِ>:�:��B��>y�k?R:�>D��>ď��"��}���׽��>G�>�� ?��y>i�3��]�Nߎ����O�8�D�=ݗf?p̂��k^��ǅ>:�Q?R�q�?�<v/�>
�]��!�8~�!��+>��?�y�=(�@>��þ�3���z��L��J#;?�84?L���>q.��=�>��?��>ɝ�>���?�s=����'0�=Ӳ?4 Y?��Q?�V?+?��=�:�o̽:�@��>fr�>4'�>��!>�{5>��f��s��%☾�Dk>�Bz>鯈=�t~��Ĉ=��$�֨���F=&}`>�ۿHTU��>�N���������T�N2��gf���V���վ��Ѿ��[���u��J����b� z��#�a��O�?��?����������,\�L�Ծ��>����|*���þ��I�����"̾ʃ��e!��Oh�-4��`�_��P�>@
���Pο�������gxA?�57?V)?+HB����{i���=:�>��S��9�F&��-�Ŀh+𾂕�?u:�>��׾1�<��V�>�(\>����fW>��������VP=�R�>qeA?"�1?�f?��!��嫿sW���?ہ@�A?��(�G�쾉�X=H��>Ҙ	?�?>U�0���6İ��P�>�1�?|��?HN=)�W�����e?!K<��F�#߻h�=g�=ܭ=<��P~J>jh�>���AA�+�۽Cu4>*��>��"��5��M^��L�<��]>j�Խz䔽5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=u6�����{���&V�}��=[��>c�>,������O��I��U��=�i��[Կ�I.�K�	�������o�߾>'EY�,�x��=QU��B�Ͼ�5�i��<X8	>�>�v�>#+>eCU>�AW?)s?4,�>�N̻�Z2<����$������
۾IԾ!��bz��D6¾e
þ��۾�	����=��O������?�&�X=¹R��ҏ�.� ��u^��t>�Yl-?��>l�̾�P��y���!̾���(?�����ݽ̾��5�Ԙk��@�?��D?�_���\Y�}���҇�6���q�S?��se�``��_��=Z���oW=���>�=�����7�E�Q��O5?�y'?4������#WU>���;�<�^4?Z��>�lý��>�@+?� 꽵>t�,��>X�c>��>�{�>	.�=F)�����4!?�#c?v�ʽ����y��>���?$���jv=�HB>���dN��JC>�K={��D[�I����<-)W?Y��>y�)����]����AN==Ӳx?�?k'�>vyk?��B?��<�b��l�S��F�w=J�W?�%i?��>j���Aо1~��J�5?�e?��N>�nh�w����.�eQ�&?��n?�]?({���t}������xn6?��v?s^�vs�����;�V�i=�>�[�>���>��9��k�>�>?�#��G������wY4�$Þ?��@���?��;< �T��=�;?h\�>�O��>ƾ�z������+�q=�"�>���ev�����Q,�e�8?ܠ�?���>���������=�թ��3�?��t?�ߜ��V.�����zy��hϾA!�;_ 2>z�
>��p���x5;��x��A����1��S��>�@ϗ�~%?(��$�ǿ..߿�	����b�D<̔ ?���>��x��Cz����M�K�� \�7aP�hc�>j>/I��gN����z���:�mT�� ��>����G�>��R�-������ڜc<�T�>���>���>؋���<��}��?Dc��*
ο����9��6X?�1�?���?�6?��<F�w�a�{���� �G?��s?� Z?J{-��^�NL7���T?K4���s��y6�K��u9>�*;?z�>�@�%�;5Й��?���> 9=��ɿ�7��g��zۗ?��?�����>���?l�4?U!��������C��";'D(?���=m��!H���I�vԂ�P?$� ?/Y�����_?��a���p���-�2�ƽ�ۡ>�0��d\�H��+���We�����?y����?�]�?�?^��� #��5%?l�>]���B9Ǿ���<M�>�'�>j*N>�7_���u>#	���:�
h	>Q��?�~�?�j?b��������S>q�}?a$�>��?p�=	b�>c�=��X-��j#>}"�=��>��?��M?tK�>�V�=F�8�d/�E[F��GR�n$� �C���>?�a?��L?�Kb> ��O2��!��tͽQc1��T鼰W@���,�S�߽�(5>J�=>W>��D��Ӿq�?�o�?�ؿ�i��Ur'�+54?��>�?�����t�k;��;_?�}�>l7�<,��&��*G�֙�?H�?��?��׾a*̼�>��>yF�>� սf���၇���7>��B?z�6D����o���>A��?��@�ծ?�i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?�Qo���j�B>��?"������L��f?�
@u@a�^?*��տ��3ξ�D���?��>Xh�H�F>Z�\�� >n|r>{�j<j2��c3>Խ�>��>�^�>��>"@t>��=ku��ӎ!�vH��ӆ���;f��:A�
��=�t�*���20<}%�z�����޾A �ߕ��1��*0(�<�.�o�=���=�
E?{�K?��o?QZ�>�:��h�=�4�ǵ�=3���T'�=�t�>�?��E?�+(?��=}��	�c������{��O͎�9�>�_]>���>���>���>:�~�G>��#>m�n>��=�H=9fݼ`�#< >=�>-�>�.�>��=�2�=1��	v����e���"��q=�y�?��ʾ-G�� ���־�����=u�%?�k>��5+ֿ�� NK?-0,�Yn�򣁾�R�=Y�8?6�L?&,�=cr̾��2��f>��ҽ1f+�PZ=2}7��z���9���>1 ?�|f>�t>�3�Bj8���P��Z����|>�-6?���#Y9���u���H��`ݾG5M>߿�>�-C�q�J����>i���|=Qm:?�o?UY������=�u��O��q+R>�>\>P=e��=mM>�-d�L,ǽ�@H��}-=���==�^>I7?�)>���=�>�>i����L��ۧ>��?>µ->�@?:�$?�	��қ��M���=+���v>�"�>�.�>o�> PI�O[�=M�>Ża>Ό��~}�]���>=���V>���"8_���|��7=�W�����=�ݐ=��I!9��#=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾUd�>fp�g\�����F�u��#=w��>�1H?(a����O�">�t
?�?ob�D����ȿ�~v� ��>U	�?	�?��m��=���@�)s�>Л�?�cY?I`i>�d۾>RZ���>0�@?�	R?��>�9��'���?�޶?Y��?R�E>�x?���??�-۾.�`�m��AR��lB9��:�>�R?A6 ?u�*��k�\p��/l�2U�6���	i=���=d�>�tM���m�We;r���3F����<�7>��>0Q�=X��<��>N�>� �>;��=j�q�Ja�$0L?�я?����m�g��<P��=_��(?��4?3W�ξ�(�>�[\?H��?�d[?ð�>ڽ�Kۚ�v������sT�<5L>S��>&N�>���.L>�վE�E�ύ�>�6�>l ���Rپ�����ǻ[ܜ>�!?���>Y��=�� ?#?�j>�,�>�bE�#:����E�6��>���>�J?��~?��?$ڹ�I[3�����塿�[�d7N>	�x?�T?�ɕ>ߎ�������OE�CI�,������?Arg?HO�K?�/�?L�??��A?+-f>e��
ؾ������>N�!?e���A�5(&��}�z{?&5?���>�����pֽO?ռ��tJ���#?y&\?b8&?ۄ��a��þ��<����Wo���;�J��T>�>t���K��=�A>���=�Um�K�5�w�p<�h�=c��>���=3[7�r��0=,?��G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>$�l���K���ڙ���F��_�ŽwM��W��>�>X`�>ya�>$�[>��>֗7��!���C�ɾ47]�X
�	33�`6?�H�R�����L�=��>漯����c�>���5N�>_��>��">�W�>�{�>��>v�
?�\�>''�>n��>� �>Ż�>��>�E=�J�aHR?����ϲ'���U����-B?jdd?%3�>��h�ˉ�����]s?���?Ux�?�`v>cjh��#+�ea?��>����t
?]�9=���mo�<�o������Y��ū�Z}�>�e׽�:��M�^9f��u
?�4?�:���̾7a׽�\��M|=S�?Pd)?��*�G�R��qq���Y�mP��K�+Z�2��Pw&�p�n�(̏�R����S���g%�UE=h�)?rn�?1����I����g�Z?C��g^>A?�>��>�b�>2�P>�
���4�;�[�w.(��Ѕ����>j�z?�
�>V�@?0;8?�(Q?��K?겒>р�>4����>�H=#��>m��>��,?q6*?�/?�i?�r,?�^K>���"8����׾�4?�`?[�?��?��?���/ý��B� ���oe�FB(=���;�F��`���@=�=X#O>&?���$9��=��}'j>�u7?f��>A��>���R/��ŀ�<=��>�c?�L�>� �Q�r�a����>���?����5=��*>u`�=����� ��~��="Ƽ.{�=�}��B���=<���=��=;���b��D��:}��;��<�t�>!�?ߔ�>aD�>dA���� ���s_�=6Y>�S>�>�Cپ�}���$��k�g�	\y>Nw�?�z�?o�f=��=���=�|���T������������<ݣ?�I#?_XT?F��?(�=?�i#?t�>v*�:M���^��\��ɮ?!)?|3�>����Ͼ6�����.�%�?Wp�>SId�NU�ϯ/�������m�M��=��5�����6��r�?��0T=P���z�����?B�?����;�&o�!I������%�??���>���>��>[,��d�����7>j��>ȭN?|��>��5?-n?�W?6�.><�3�"lL����5=%D�>rM0?�Jt?^?��g?Q��>�[6>�������*�<ွ(H�[����U�=��>	��>��?U��>�V>�;M��>½-�]��ʻ=�y>���>9�>g=?}hq>� =~�O?y?�Ѿ�I�:������E��K��?_P�?K{?�#�<�r�_'8�ؠ�����>
E�?�;�?Ś?@�����=�<�����Ql�J'�>��>蠰>�Z�p���7>ݰ�>V�>I�Z�����M���ۼ��?�B?�c!>�ſ��q��p�آ����h<qВ���d��g����Z�H�=���@���۩���[�3���fY��I�������`�{����>�q�=��=���=9�<>Ǽq��<�#J=)�<��=K1p��g<t�8���׻zf��dJ(���Z<�J=�����/ž��u?�F?��.?D�F?:ă>�l>�~��˚>�VT�B?ScM>u��l�����3�<ݦ�(���iCվnpݾq_�[��	�>>78��>}�5>�n>2�<��=}�=m�=�#1��GF=ͨ�=R�=��=���=�%">Ɲ>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=J����=2>s��=v�2�T��>��J>���K��C����4�?��@��??�ዿТϿ7a/>�Y7>�>p�R�wm1�]i\��Zb��|Z��!?	1;�u8̾�@�>���=�߾��ƾW�-=|�5>Ǆb=���3\���=B�{�Z<=1^k=c�>�D>�^�=u���ζ=z�J=S��=�$P>���C7��P*�4�5=U��=��b>4&>W��>�A
?Q?"?\\P? X�>�Q��������`�>�����>6�5=/V>�8?r,??�[B?�$7?�H�>)�¼�\�>5�>�P3�z�y�'� �\�⾋kZ�*��?J��?�nv>`��&�Ȫ��%�ݹk=��?�?ܙ�>0b>{�2��i�&�>�,������s�J=.�m�?�>�#�w�F�����B�=�>R��>�ɡ>p�>e;>�N>bk�>�>���<Ŕx=[�;��<W
���τ=�"ļ��}<�����+���^�
�4�hvѼ��; A����HRP<���=:��>#<>���>Ԓ�=���~B/>繖�|�L�Y��=H���+B�
4d�:I~�$/��Y6�^�B>?;X>�z���3����?(�Y>m?>G��?wAu?!�>#���վlQ���=e�>[S���=�>	�<��z;��X`�n�M��}Ҿ݀�>���>�=*>��(>98(���4����=�;���N��	�>Z��ߜ�t��=r���ˬ�᳥�:y�>r�=�m?(`��ԩ�=菙?C�@?��?�,�>Z:@�}�����[>����ִ�>�LK���6��<֧$?�
?~��>�َ���u��I̾����޷>�AI�3�O�����?�0����ͷ�N��>������о�#3�Lg�������B��Mr�#��>��O?W�?�;b��V���TO����()��q?�zg?��>L?PB?����s�o��$��=��n?��?$<�?q>�@Z>Y���\�>�f?y6�?2?��_?����?/_�=8YA>�.��� =��T>�1d>JKe>n�?JY?�~�>��r��T
� ��V>Ծ�oٽJ�	>s>t��>>��>���>u��=��=�x�<��>YK�>��>_v>���>/ �>.Kž�O�-O'?������> ?H�>��"<]�x��7��y;`=�`�����<���<X����W(=&�=�Tf>8��=t�>�X¿�?vi=��P���>K���p����>naH>X�B��O�>v<>=��>�p�>�]*?)�R>b��>��h1����>�="�<D��TJ�`)��J^��7U5>w�����O�sc)�9:��f.:�"�Ӿ����q�Q�c׆�|ps�8��=��?��=�	d�0.6�T½|�?#�>�?3
t�Q璼8��=��?�{�>eJ
�[���ć���Z�'��?c��?�;c>?�>�W?7�??�1�3��uZ��u��'A��e��`�R፿������
������_?��x?�xA?�G�<�9z>"��?��%�2ӏ��)�>r/�d&;�BC<=++�>�*���`���Ӿ�þ�7�sHF>$�o?%�?~Y? TV���O�2D>�8?��5?:w?�I3?t�4?�)�%?`�<>̴?��?�)?L�'?�%?C+(>�U>D���><g��5k������������û��N=)�=��;��)��;�u#=�~�'z�D�f:���<<�[:=���=к�=�B�>��Y?�.�>fl�>�8?�"�p�7���H�/?N�X=*��-ᇾ>��)��3>o�h?�׫?��W?}U>s�@�T�B�S�>K�>�/>��c>l�>�:�� <I���m=p�>>{
�=Ғ[��Ă�i^	��H��y=��>���>4�{>F���2(>N.����y��"d>`eR������FS��G���1�:�v��C�>t�K?\�?b�=c�W%���,f�q)?�C<?dFM?��?�P�=�B۾(�9�B�J���k�>��<����������:��b�:�\t>����׾�'	>Pa�}�۾k;S��4?�̾��e:(�)�96=�b����ʾz��=D�2>æ��/E1��V������1�I?+�:>S�����</�lg0>]�>�ĕ>D9����:���o��e�C�;���>�Q=�Z���� ���J�˩쾗؍>y�A?N�V?΁?A&s�_V_�K�;������by��#��P?�y�>��?�Ή>���=	���#��[�T��H�6��>�p�>���$�N�jƾ��!�
�f��>���>]�>�?r�]?� ?��p?��$?w"?�F�>�(<s�����2?��w?�Q�=�� �پ�]=���K�I?��2?�����>)�??g	=?BqP? \M?��!?�Y�>�P����D���>���>�^��a����A>}?5Q�>�ׂ?9o?E>�2��Y���ý )W�hK|>�k6?�'+? v
?��>�]?2E��e*
�r�?މX?(u�?93r?J��=��)?���>�hp>�H<c�>�3.?	vB?��_?
�`?(#+?P�>���<QE.��糽W��:��=@�M>����̃�қl�r߬<�Ș�� �;n�u�<N�e���#�m�=�%�=d9X='P�>jDt>z*��1�0>�žHY���~@>���Y���⊾�;���=�h�>��?�]�>�~#�3��=���>o��>���n(?�?:?��,;Ūb�<�ھW�K�=�>d�A?��='�l�Y�����u��Bi=��m?Jl^?��W��`���b?��]?{f�%=���þ �b�Պ龎�O?��
?��G���>��~?��q?ʶ�>��e�*:n����Cb���j�ж=r�>/X��d�o?�>��7?�N�>��b>�'�=�u۾��w��q�� ?i�?��?���?�**>w�n��3�\��������^?K��>�t��	"?�NĻ0�о�ˉ����x�߾M;�������U��m���C#�ׁ��ҽ#��=��?�3s?�5q?n$`?�� �#d���^�/��P*V�������`�D�,^D�ED��m�M��Ҙ��l����==
z��V�dh�?�
?I��<^��>�>^��N�6����s�=z�?���,���=�p���*4<�q�=I�W����Q��7�?�$�>���>z�B?�hP��!F��	E���;��(�9c�>z*i>��>�v�>Z���2���8�s����("�@�>�i?EK?�LT?�^���2�����=��=�=�!=���»���=n$)>�Ӊ�{v����A��Y�A���B��N���9A���"?�
u>�c?wɏ?���>u�����=8���a��=Z��>��Q?" ?t�>�罏��v�>�Ad?��?�=�>>���U`1���������J��>`f�>�?p_>?�3�zj��Џ��K��0k4�a��=��V?��k��1��G1>�2?�+���,=�
�>�ħ��*,��'�i]ӽ��D=IQ?7�6>���=�뾾�;���t�kr��(E?��)?!]ž8��S��>?���>�B?�~}?��+���ʾ���>'AE?��O?�C?��S?�-?|�m>��a�rڽ��I�9hR�֝�>EP�>�&�>I�4>��[��׬������=|F�=��{=�	�濽��Y���u�kP=]�[>�aۿ�K�@�ܾ'���"�ɝ��↾�b���o����
�F����l��M܂���,���M�bh�Ob���%r�W��?a�?H���Ɖ�+噿����N��n��>o�g��Ր�H���a	����CH߾�����#�v�P���i��Ie�L��>��ҽBͷ�
K��{f뾨"?�>E?��5?M�/����Ea�U�����<�2�P%������ӿˡ�����?��?����/;��W�>��>��=f��>57[����:��>�`?��W?:���Կ:�¿�|C>��?ap@>}A?3�(����GV=N��>��	?��?>�F1�F�(��T�>�<�?x��?8�M=U�W��	��~e?��<��F��ݻ��=C�=�9=�����J>�X�>�u�XA�G3ܽ]�4>�م>Br"����S|^���<ʊ]>U�ս':��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=u6�����{���&V�}��=[��>c�>,������O��I��U��=�E���ɿ)pM�t(���=ʇ=�9��`��г���;���;�hs�GY��o�=-��>푿>$yf>��E�& >�ZU?�Op?	��>�0�=Zac�~�+�"U�� ��=�Sڽ)�i�v��$}��}���˾V�ҾR�891��/�w�߾�t=���=�:R��b��$[ �̀b��%F�G.?�� >jnʾ�M��k<�˾Se���w��o���;�-2�5Tn���?�7B?����W�&N�'���G���)W?�����M/�����=���d=���>�D�=�}�q=3��S�y+;?׮%?�aʾF(��cw�>�����=�G?�/�>��Q+�>%U<?�E�<�����s>g>���>���>��=����G�UI)?��T?���@�e�~|�>����	{��L�=p}o>,�|�����>F{'=�����ns��?����/*W?Ҧ�>��)���T_��r��Pf==�x?��?&�>�rk?�B?��<0Y����S����w=��W?�#i?7�>���о�z����5?�e?��N>)hh����.�$R�� ?�n?�V?i۝�7p}�������3o6?��v?�r^�ss�����<�V�A=�>�[�>s��>��9�[k�>��>?{#��G������Y4��?z�@���?��;<�"���=�;?�\�>�O�\?ƾ�{�������q=y"�>x���zev����Q,�x�8?堃?���>��� ���!�=�Y���J�?�<�?�KM�`�9�|�'��Lt���Jc~>t��=Y��<�P����0���ؾ�ھ�_z�g-���Ɍ>�@H���w2?!����ѿ����W�/&޾��g>���>+ �>��A�w��(�X�,I���U�b�I������`�>��>�0���ӑ���{�ya;��ß��>���r��>�;S�P���3���C<��>H��>;��>j���� ��Ѻ�?�O��c-ο��������pX?'a�?�?'X?��:<��v�{�i�5G?�zs?�Z?Q�"�#�\��Z7���_?�`~���f��<�1�O��%N>�-?�>��/�׫�<M��<ju�>�\>�G��,¿/��axǾ�˪?H.�?�&��h'�>�+�?{8?(�7ܜ��H��R�(�b[1=|�3?RZa>�Ͼ��4�!�5�1F���?�0?�����1�]�_?+�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?_,�>��?���=�\�>��=x����2�xH#>2/�=-�>��?�M?3�>��=�8�//��^F�MER�,(���C�Q�>��a?D�L?�ab>0����1� !��)ͽX�1����pA@�[,�QD߽>D5>H>>�>��D��
Ӿ��?�ƾ��Կ�*����Z��d?�~n>3��>��	��h���c���iN?*4�>�,��n���ŕ����wR�?z�@���>3*��-a%��&>��>Ɠv>&�žz���Ph�x�>�$?D��w⌿������>=2�?@@r*�?�$i��	?B��O��b^~�Ҁ�1�6�4��=��7?D2��z>���>�
�=fov�E���.�s�!��>�B�?${�?8��>��l?�o��B�=�1=�J�>�k?�s?��l�+󾟹B>�?��������I�4f?��
@-u@�^?��Q#ѿ6����;-W����><|�=2i>wy�����=^ix=l�C=�A�=��>��>�V>�ۇ>d�d>�D@>*M>^����l%�����L��`q8��+�1��WtI���������S��aˎ���6�Y˽������r�?u���2�>S�R?�mM?Q�r?w�>,g�t6�=@H�/�=�_�2.i=���>��0?A:J?��$?a�=*����`��,��r���'|�����>��%>B��>�>���>n7.="��=�>�3�>�S>a�=���=,?R=�A>²�>�D�>�I�>D�2>��>�,��Oİ�	Xh�>�w�(�½|p�?^����J�%���������H�=8 -?s� >w����п����3sH?���4���q6�p=�=��1?KQX?��>������c��>nx�s�d��8�=�b���s���*��oO>�L?��b>��r>Ԛ3��s8��P�?����5{>�5?a���9�Hu���H�Fo޾��L>޾>s<��}�C&����~��h��y=>�:?��?L.��}4���uu��읾��Q>��\>^a=�ȫ=W�K>�e���ʽ��H��.=YO�=K�]>CM?��,>z��=d�>�����O�辨>�@>�.>{@?�$?���N��i�����-��;w>"��>�S�>kl>��J�䌭=���>Ѡb>{^�˯|��;�֨?�m;X>�����]�z�x��E{=ݮ�����=Η=9���I>��"=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ>p ���f�����|i����<��>2:?S���K������f�?"$?�l�5D����̿��x�J��>x��?0�?��g��'���<2�ͭ�>�S�?�f9?��y>����Ĥg�:��>��N?�P?�a�>J��v�P] ?���?	i�?\�>8̈?'�?���>;�����X�E7��.wf�^�����>�L�>�߼���ʓQ�~&���ŕ�JYw�L��Y��=鉤<9�>�Y�'����!>����UG^���|�[>Y�<�k����<>=��>7��>G��>R�=
9�����f��B�K?}��?����+n�=��<?O�=�^�F?�R4?�^���Ͼ��>>�\?D��?;[?	~�>��S-���޿�ot��@�<ogK>��>en�>f=���JK>��Ծ�8D�j�>Կ�>9��<1ھ�M��:?�� A�>�Y!?؆�>(o�=��?(�!?ɲ�>ɑ�>��M�� ��T�R���>v �>�!?I1~? ?:��Z�;�����v��%�X�v�E>�m?i?�d�>�B���V���ٸ�-��7��ߢ}?݋N?�J�dW?y?��=?:�L?y8>1/��+뾡B��{{>\�!?��,�A��J&��
�,?O?8��>P����սPpּ���R|��{�?�'\?OA&?���*a�� þ	'�<A0#��V���;m	D�7�>�>`������=\�>g�=�Rm�MA6�Vug<�s�=���>��=�27�3{���4,?�D�"郾Ϩ�=��r��wD�>�>�"L>����^?�=���{�G
���}���8U����?U��?�o�?Dk��ˤh��=?�'�?�?p*�>�a��nv޾`��w��x�a���>���>�Ah� ��܂��*���E��e�ƽ��,����>C��>�R?�>?��]>4�>�ꗾ��(�A���!���V^������7�'�/�=���q���J���x��^���`��5ڊ>�Q����>˒?|�>ii�>���>�>=yޮ>�QF>~u>��>z!c>_mX>��8>>��<%���NR?����'�"��t����4B?@qd?�I�>$�h��������Z�?���?r�?~Fv>loh�5 +�_q?�2�>�!���i
?;=���P�<F����������ָ�>��ֽ�#:��M�?f��h
?Q&?Z��]�̾vW׽jn��f|=�ˆ?�4.?m:,��U��t���W���L�9؃<o/`�NY����#�ۯu�d���]���Lˁ��G%�uw=8�'?䖉?�#�,y�aK��d�h���@�`kp>8��>D�>�Q�>��>>;U	���0�vN^�SQ*�gP���8�>k�w?E��>��D?.�4?�`?P�H?�w�>��>�hb�O?�"��h�>���>�G?�A?,s6?��?��?
�?>^;�$��q���־.?N~9?�`�>Y ?���>�7Ӿ���=�2+>d�|�j_�����)��=�+>�	��K@$��Mǽ��=[?����8�e����k>׀7?{�>3��>k���7����<9�>a�
?{I�>�����vr�P^�[�>Ϡ�?N�o=��)>�=����̺�k�=�¼�ΐ=|���R;�W]<r��=��=4u�곐����:a�;\G�<�5�>�?Q�>��>B����I�����%�=�Y>19Y>�N>�RؾXQ��f����g���u>�(�?8$�?�kd=��=���=������D\��ͽ�$��<��?�k"?�S?&��?��<??#?K>�q�EA��AI��%ޢ���?t!,?��>�����ʾ��։3�ם?e[?�<a����;)�ې¾�Խ��>�[/�h/~����4D��ꅻ���b��7��??A�X�6��x�ڿ���[��v�C?"�>Y�>�>O�)�y�g�n%��1;>��>eR?�W�>��O?��z?8�[?B�S>�Q7������p��֍��A>�??�I�?���?��x?��>��>%�*���߾���16�N������)�I=u!V>�L�>z��>�#�>x)�=��̽D����16��²=z�k>�S�>��>���>D�{>�<LH?���>�u��à��A�����<�Cv?v��?��*?�v=Y~�1E������>�_�?o�?6*?�T�H0�=GҼ褷���q��<�>2�>��>��=��C=�]>�~�>_B�>���_���)8�saK�p�?��E?���=(ɿ:~w��E�������0d������Z���)�~�־�>�"�ږ�]c�F�S�a���*�c������1{���%�>q��<2.�=#A>�.>3g���=LjP=�{�M��=���=���=L�㞀���ӽTj��cŻ��<�;�ַʾ�m}?�'I?7�+?sC?*#z>��>�9�㽗>$M��\�?GU>e�Q�Ж��;�������s�ؾ�
ؾ�?d�?����>}�B���>5�4>��=x�<|��=�Tf=��=;$�=��=g^�=?��=��=�>~>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�47>(�>��R���1�y�\���b��tZ�j�!?�H;��4̾�F�>~��=/I߾v�ƾ~/=��6>�a=^���Q\�Cƙ=9Z{�8�;=зl=	��><�C>q�=�#��2Z�=J=N�=��O>�ј���7��c,�D�3=���=��b>��%>���>\U?�[.?1�_?���>��k���˾Һ��zA�>���=�'�>y�=9e>^�>�{5?�A?c�G?ԫ�>�j,=<~�>�>��*��(q������}	==$p�?Ƀ�?戵>]m�<R�!��.�]�/�{Ѡ�S?��5?|�?��>�0�h��I/��1���O�� f��z�<��v��Ƚ+��!�������=g��>l�>s�>B��>�O,>��J>n��>��>��=R��=T=�<���<���&=���+ Y=��1<G|�����.l��3ɻ�������5\)�ɜh����=���>A>���>��=���^/>Z���x�L����=xZ���"B��/d�AR~�K	/�)a6�t�B>IsX>����4����?6Z>��?>n��?�-u?��>�8��վ0N���e�ʀS��N�=.�>r�<��l;��V`���M�$�Ҿ��>v��>E��>�tA>��6�*�>��}<b��3�0��>�ȫ�U޺��>$�O+���w���G��-[L����=F�L?Y����>�=`׊?��Z?"�?䔣>����ޡ�Fh>B������=8���y���gL;kG?��&?���>í����M�6Q̾�*��nַ>��H���O�����	�0�Y��䷾�W�>bݪ���о+03�c�������B��q�b�>x�O?��?�b�Q���XO����р���w?�g?i'�>�Y?�^?00���a��K����=i�n?s��?�4�?��
>�L=A;�.�>)�?I��?Q�?�Ai?i/��c�>�%���B>���A6��5�=�!�; �=S?�7?'�?�م�oj����	�ڛj�Gu���>�(�>�Y�>�N�>!a�>R�=��=��>���>_�>���>*J�>�0G>�ֱ��X.��0?Z��<�S�>:,?Nմ>���<`�i������G>z��E�����潤�R��|n=#
�>$ʒ>3�G=F��>lƿ�Ӧ?�-μ�St��G�>�=���Y��9v�>��6>/��<y6�>t_�>�l>e��>+��>�	�=�>J��=���j>[���i3��I��z<�9���j3>x5޾�dX��!�c��ʹ�v���� ��_[������_�ӊ��_�?fc=5�L�y>��4�h�?�}�>�?DY��ݗ��C����>4�>J���d��|�����Un�?�� @<7c>Y�>k�W?��?��1��3�itZ��u��(A��e�ݺ`�l፿E����
���n�_?	�x?�yA?dc�<�8z>桀?��%��ԏ�/(�>�/�%;�e<=�+�> &����`�ˮӾw�þb3��JF>͖o?�%�?�Y?gWV�_7N=�C>�,:?�N\?twn?�4P?	�C?M����@?���>�>�>��?2�/?�'>?�e?��>���=�����p/�0�ٽ�x���u�S�!�(p-;��=��=��=�8ƽ��%=Y�N=�[A��J��;Ԇ;T�;x>��ҥ=���=��>iɦ>�]?B�>��>��7?2���p8�S���R3/?ǎ9=����L������e�]�>��j?���??XZ?�4d>��A��C�)>�c�>ɕ&>�@\>/l�>]��J�E�tb�=�i>�=>��=��L�����غ	�������<�>���>]-|>}��:�'>�z��/+z��d>��Q��ʺ���S�Q�G���1��v��Z�>=�K?��?5��=�]� +��If��/)?(^<?�NM?��?��=X�۾��9���J�z<���>�d�<�������#��Z�:��+�:��s>�1������`>�u��ݾV�n��XI����� \=gP��#H=�=�Z�־oE����=�	>���(j ��떿ڊ��O�I?��e=\���O�T��e���X>#Ƙ>���>h�,���u�I@�\����Ö=��>g>>E���3���G��9����>�$7?�6?r�f?�t���R�m�6�0Ҿ�����=_?Nw}>U�>E	�>{V">���#]��k�@]H��A�>���>���U�!D;�
��:	��>Aq�>j~>�N ?�'m?3��>�AG?�N?��8??�>q��zx�#�!?�(�?�w:;�����U�(:��|<��S?=s?�]��OW�>}P?MX
?3�1?��e?��?�� >Uz�a�H����>�p�>"�G�I���z>�*.?!$�>q^b?T��?�� >R��1��mj����0�>�A?{�,?T$?���>m�A?�����)�>pX)?ʥ@?�}�?�X?�ǭ���>mv�>�1?5��>���>:k�>! .?\�s?e�T?��>{�>[~�=b�%�Wt�<X˼_j˼,D�=gV�=,��=���?	�!%B��0��d�g���a���;.$��*潪���x_=+T�><�s>I/��x1>9fľ�܈�g@@>�v����� T����9��ߵ=[��>?-??��>u�#��Ȑ=�+�>N��>:���(?��?��?߅k:��b�_ھIK��%�>��A?Yh�=�Al��^��Y�u��_m=�Kn?6i^?��X�I���bfb?�]]?��^<�?�¾�`��z��RO?�|
?g�D�%5�>��}?�Uq?���>�ld���m�\����b��j��ܶ=k�>���,e��R�>��6?7��>g�c>�>�=��ھ�u�G0����?��?��?�y�?{.+>{�n��࿚)������&�\?��>�5���$?E�~�Rʾ ��k���ol徣���ᐨ�瑗������*�vU���r��6��=�?�z?��a?��c?�/��5Y��V`�s����X����I�
��F���>�ΐN���r�|��W���a����k=����Jhl�[�?��>���׌�>f�g��T^�(�%�O8>:�ھė��_o~={��<j�Z=�Ǌ=/-H�������� s?��>Egn>&�D?�c\�1���T�фg��(�F?�>���>���>t_�>�]V�Ѐ���C��ל⾡�]�B�����>��z?tO*?mW?�c�z!D�v����Z ����s�J�(�>�ѻ��&>��ؽ��wG�i�Q��5X�	�	��l�����A��=�?sM�>�I�>��?��?x�ᾧ�ξ�>��ط$���<>Dk?[u{?�V�>{�>a�M<���2{�>�m?���>���>��r�!���|�^?ν��>�ݮ>O�>�Hn>��.�#�[�}H��F�����9����=�"h?�ꃾ]�_��>`�Q?^;; �@<؍�>��r�Ƌ!�"��B'���>i/?��==>W�ľ2���{��g��&?Sq?�x�����՚>�?�2�>&�>��y?���>������w=��?�T?��X?�/<?'�><.��_���#3����<��>��>I� >�=9c:�e53�^�E�p�c=�=>:f=K8�3&{���3���0<;�c=��T>޾��b��ھ׉��{���QKT���=ލ�>+_�{Ͼ>F��چ��#�$�S_�L]�<S��dǝ��ł�)��?��?����,������d�i�Ӿ֭>;�|�e���,;�#l�":p���پg>��t.��P�|�i��=��?95��xǿ{4��ξM?��*?>�X?׆��/��+C�.��;��=#猽���;��qϿqQ��I1~?���>˾�2���>!�>�S>d%>�k��:\��)��=�p�>��)?F�?�{�Gſ�⩿�FQ=1v�?�2	@��A?B�(��9�p�W=q��>��	?�h@>Aj1�-V� j�����>d4�?�ߊ?o�M=�VW��-�Le?��;8�F�)�ϻ��=�s�=W�=���DJ>��><�_
B�i۽�5>Pʅ>:M"�Ak��^����<]>��ֽ�m��6Մ?){\�~f���/��T��U>��T?�*�>2:�=��,?O7H�]}Ͽ�\��*a?�0�?���?$�(?<ۿ��ؚ>��ܾ��M?[D6?���>�d&��t�؅�=6�܈������&V�f��=[��>Z�>Ƃ,������O��I��`��="���ƿl�$�\�����<���ՉR�$g��Ϭ��f�?o��%hr�-x��b=���=�P>~{�>+T>��W>�AW?3�l?,h�>��>���Iԇ�?;̾{��������43�� �~n������{�4/
�>�##�6�ƾ��=��f�=��Q��M���!�;�b�U�E���.?�'#>�̾ɻM�pe�; �˾�W��ꆼW��jJ̾�1��m�?�?��A?tⅿW�����������G?W?"��H	�����G�=@���j=�U�>(E�=C��A�2�ŨR� .?='?��Ѿ&�����>�Z��۲=�0?
�>�/��7�>�>?F�2��䧽���>AK�>[h�>[ƹ>�a�=����~I��?�*\?�MA<m�E�_?�>���󲊾e7�0�=H�����=��c>6�����w
�;F���h���W?��>r�)�I��>ݏ����f<=��x?�~?�>w�k?�-C?е�<�(��m&S�M�
�{�w=��W?z�h?��>�Ё�}�ϾaƦ�l�5?��e?�TO>ji����F�.��0��X?a�n?f?�妼jX}�N���A���G6?>^?�P�����ќ�bVi���\>G��>A�>�I�^�>�;,?��E�턙���ſ�A��?W@ @h/�=�Z���=
J?���>x�������։�Sh����
�?Bx���q��x'�,1ڽ��?Czw?:?s������џ=�ᠾ�>�?�i?��Ͼ>�3�7w���b��߾�Վ=�_H=	��<~��:vN�R;�
�پ����l�Y*J�f��>��@g(���?�����ƿ
Uѿ�����Ծ�&�`�(?G&�>i�	������Gs�������T�9�6�[�d��w�>N�>��������{�� ;� Û�'�>�U��>�uT�P���eڟ�4$E<���>H1�>���>�������ъ�?�<���Ϳ�E��A�W?4�?�D�?K�?��C<��u���x�"l��G?��s?�bZ?�f"���\�Zh>��j?�^���W`���4� GE��U>D"3?�@�>A�-���|=�>���>^>"&/�P�ĿEض�{������?���?�n����>u��?et+?|l�F8���Y����*��S2��<A?�2>����ܺ!��.=��Ӓ���
?��0?�|��0�Q�_?6�a��p���-�1�ƽhۡ>��0��e\�DJ��&���Xe����Ay����?A^�?d�?���� #�L6%?%�>f����8ǾU�<À�>�(�>�)N>DH_�z�u>����:�Si	>���?�~�?3j?󕏿����	V>�}?�*�>��?�H�=g_�>a��=����+�S�#>��=��>��?&�M?�[�>���=ѧ8�/��CF��ER�4,���C�,�>��a?pmL?f5b>X긽��2��!�i�̽�$1�o#�ϩ@�7�-���߽h/5>v>>�>�E��Ӿ6Ƥ>����(�I���<i>"?M�>���>m���ாO����?�>��I������r�xyg�t��?
@s?�ٸ��4�-A�>���>�<����_��;dqN��C<>'�<?Lo!>Q���wl��+��>/��?x@���?(Mb��*�>^*��J�����z����e�T���=��(?����V*1>�x�>�u^=��x�c@���Uv�ֲ>ǰ?�`�?#/?��`?�a�e-�'8	>�J9>�!E?�k
?�!�;d��jC>��?*��H��l`����O?Y�@?@�T?�����ÿ�d��5c@������<0B1=/�R>���8m0=�>=��h<��0������C;>I,>XY>4��=�,>W<�;��� ��ۨ�����;Q��4@�%F˾�+��:c
�������@��)�����H�qM�K|#�&mξ�����!�j>�	T?�=?E�c?X7?\��e>�	���=�ֽvV=s=>��0? �M?)�'?g"[=�u��bc�3���������F�>�/>>���>@��>8��>��K<9n�>`wR>Rn>T�6=(��=ʧ�<i�
�Yx#>�ȥ>h3�>5L�>C<>^�>.ϴ��1��b�h��
w�̽)�?����E�J��1���9��⦷��i�=9b.?|>���?пX����2H?����m)�L�+�7�>B�0?�cW?��>���|�T�J:>���~�j�1`>�* �q~l�o�)�w%Q>Sl?��V>�,i>��1���5��sR�vt��sT>�6;?â��&�M� cv��:I�q�ྞ?K>q��>["��N��ݕ�a}��Wb�?\=��9?�?�ﲽ�𵾄p�zΙ�7Hq>��^>4�
=�g�=M�L>��7������E9��Y?=T`�=�sT>=E?�)	> �
>A�>N��U	��S��>@�=~��=d�D?v�>?��&=������a�g�u��E�>�>��>���=����x�=C��>j�C>��Y��@�5�H�P�=v5>Sq��,�Y�쿵��bM=y�Y�� >=��=�]�0�1�;le=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�-)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾC��>����q��!M��^Tu�z�'=�_�>�sG?N�����X�/6@�1I	?�)?���Ȥ�y�ȿ��v��P�>nL�?�ؔ?�Em��,���?�j`�>�<�?O~X?�i>tھV�W��,�>�@?�;R?�A�>@K�O�%�W�?%�?�?��3>��?jsO?�h�>t����
d���׿�Ǉ�wP�>@)�>��>F͋<����IJ����1���� ��ΰ	�NoO>���=���>b#Q��B����>�n���,�@�w<�4�>{�%>	�w>e�;Z�>���>ž�>�a=L��Oȣ�׃G�ޑJ?�5�?Z��vl�^��<��=G}_�2�?�]0?�eS���¾���>2Y?w�?��]?T�>�$��x����� ��(%�<�,H>���>��>�唽�F>�\ʾ�+3��|�>�̙>w��9�'׾[c���g< ҥ>�"??��>��=G� ?�#?��j>9'�>/bE�L9����E�S��>���>�J?��~?��?w׹��Z3�.��}硿=�[�Y9N>�x?U?�˕>F��������EE�!hI�1	��J��?�rg?�I�K?�/�?c�??��A?W+f>���ؾᶭ���>?�"?����y5��C��q׽ݻ
?��>B]�>�	�����~>=���!�g�?\SY?��?~���_��ܿ�
h*=��:�呺�;;��$����=B>��:�j=�>�s>��%� 3���<N�>�|�>�1�=��K�X�ѽur?g��;�L��n#�<d܉�<z\�X��>���=��
�� @?{�F�N	w�t:��*����ľ��?�?��?��B��a��B0?��?%��>��v>:�����˾�t̾`�A���Y���Т�=q�>��>Q_ݾ����Po���H��z2]�5���1��>{��>�c�>N��>�o}>p�>����P4�"�/���{�d��&(�2��7�Fx�&z��Ig������3���Z���ۂ>�n=^�>�7?6s>�?���>?Ӿ�=�<>>��:>c4�>�L�>䁂>���=�d��.
��R?�u���'�p������oB?5�c?���>@�e�[���\�-�?fK�?Mq�?r�u>Noh��O+���?���>Ē��6
?�g<=U�0�_`<�e����������XX�>kUѽ��8�;�L��e���
?��?"��sf;ZKܽJP���=� �?��?G�:�bFF���r�Gu_�'>�괔<��d�"灾�b��v{��P��`�k���.`��y�<-%?��?�2����þxb����a�0�S�J�>��>�s�>(��>V_>YH��+���S�s;��q�����>$q?�Ɯ>wFG?�c%?OBH?ǟW?�_�>�T�>1"��(|�>v��;ǽ>�a?�TA?�S,?oL6?#�?� )?H� >��<����EϾO�?�;?)�?!��>F��>�H���
��V�n<Lf�;y��������=��ͼ�޽"���{<�>Me?(j��$:�����+Ⱥ>%�-?.��>)�>�G�����.<'W>a$�>4��>�Qܾ��~�]U����>0�n?s����9�@� >�;s=����Ul�<5�>\���<�E�<La>�	�<Rx=�EF=B�T�|�=�)��=����<�t�>1�?���>�C�>�@��<� �[���e�=TY>*S>e>�Eپ�}���$����g��]y>�w�?�z�?�f=��=��=�|��}U�����J���4��<�?7J#?(XT?Z��?l�=?Vj#?�>+�hM���^�������?w!,?��>�����ʾ��։3�۝?i[?�<a����;)���¾��Խӱ>�[/�i/~����>D��텻���V��6��?�?PA�W�6��x�ۿ���[��{�C?"�>Y�>��>U�)�}�g�r%��1;>���>lR?�&�>*$P?~7z?�H[?qUV>�68�쭿<o��<�"��`">j+??C��?n��?�$y?h�>Q�>F+��߾�S�����������mW=�\>�%�>7B�>���>>w�=Xǽ^����?���=̚e>�,�>̉�>\��>��w>��<"�F?ɼ�>����Kf����ba����L��7y?�ʎ?��*?pFi=aN���A����qy�>a,�?[��?Ӕ&?�FX���=�˼�3���c��̿>�F�>��>ĉ=\P_=��>���>Y��>-���&�R5��d1��?RF?���=��ſ�hq��o��+��>�;�Y��`�`�Jt�� Z�	8�=>8���Q�/뫾�7[��ߠ�(���@>��;X��[|��4�>��{==��=U��=��<��輽�<�`=��<�!=�s�)��<�g5�qm��3k��~;e��<�T=8m�l�ʾ�u}?�H?�|+?,�C?'�y>K�>�1��>H���r�?D+T>>uN�^G����:��]���L��`ؾ�N׾��c��-��{4>��H�_P>�4>Q6�=�<�<y��=��v=o?�=�Ί�&�=���=�=���=s�=��>R>�6w?W�������4Q��Z罧�:?�8�>M{�=��ƾr@?��>>�2������wb��-?���?�T�?9�??ti��d�>K���㎽�q�=L����=2>Y��=}�2�Q��>��J>���K��F����4�?��@��??�ዿ΢Ͽ8a/>�;>�>+[Q�:�/�8X��Zi���Y���'?Lh5���þn�>52�=��پ.Ӽ����=�I>Њ{=���"6Z��p�=�t���(=�=�=�+�>��I>7�=2Q���b�=>�<
F�=�Ap>�PZ<�r�����i�^=���=P�p>��3>�:�>�s?@0?d�c?Ϲ>",j���;Y��D8�>���=�|�>�,�=7#A>]�>
�8?�BE?w]K?�O�>c��=�!�>�>WG,��nl�O�i������<q\�?�{�?���><��A�����=���½�?�<1?C\?�Ş>�U����4Y&���.�y���4��+=Smr��QU�I���jm�n��e�=�p�>���>��>ITy>��9>��N>��>��>�6�<�p�=�ጻǿ�<c �����=7����<�vż����t&���+�Q���U�;~��;�]<���;g^$�s&�>���=���>Ԑ�RkȾ�9>G9��{Y�{��ο���B���a�N~���F�{)X��-�>��>]첽Y<���f�>g=�>��!>�.�?me�?n�)>ք=���W;������8�Y��>]�g>�ݠ��UF�=#��w��:ܾ<��>ߎ>!�>�l><,��!?���w=C�$b5���>}������+�b8q��?��k���mi�Һ۞D?�E��!��=�"~?��I?]�?&��>���?ؾ�80>�M����=���'q�\����?'?���>�쾘�D��W̾�.���˷>�SI���O�����2�0����Ϸ�}j�>�	��M�о:!3�~d��.����B��Hr���>��O?	�?VBb�U�� HO���uG���h??|g?v8�>QL?3;?�衽�l� i��bǸ=��n?7��?�;�?	>��=�R����>8)	?�@�?���?7�n?^}<�<��>�t<��!>����
�=`C>���=+��=�?&n?=R?fg���{	��*�R^��l=%1�=l.�>�r�>W:u>s�=��c=���=�\>�Z�>�K�>��_>緞>�$�>k��<�x{(?��'�P�%=���>�~�>��?��>��þ�^���{�����.�l<uC���=f�	>��:=�X��>7����&�?�+6�ĳY���(>h����]��j
?��>|���&? &�>x��>A��>д�>�1O=��>b��=&?��*=1�!���K��*I�o^,��M=��F�=�@˾y���	�#����#j�O�ξ5�ړj������N��<>�?L7>��{�x\?��n<�:&?���>p?ɷ�������i�=ӥ>kr�>`��Y���*���@%澉�?ag@2;c>��>1�W?�?R�1�3��uZ�ծu�R(A�Fe�]�`��፿����
�����_?�x?yA?sQ�<9:z>=��?��%�Jӏ��)�>�/�';��@<=�+�>�)��3�`�R�Ӿn�þ�7��IF>��o?4%�?|Y?lTV��o>{�+>KM?�c?�]?E�&?�]?԰"�;�>�_>D�?�s6?��?_�>?BP?՟>ʇ�>J`���Z�Z��n��T�=��6����.E=*h�=��~�cV#��7�=��O=<���oj��=�pʼƞ$=G�U=,N�=b�=~�>b�]?5��>G��>��7?�\��I8��S��&/?��:=K ��4r���E�����)R>��j?8׫?UZ?�c>s�A�	C��>���>�G'>�\>�p�>K��cfE��Z�=��>�>_ק=`1N�p@����	�]��>$�<�L>���>�)|>�����'>z���.z���d>4�Q��Ⱥ�~�S��G��1�uv�QX�>��K?��?���=�\�O1��lFf�,1)?PZ<?�PM?��?I�=#�۾D�9���J�%<�b�>^Y�<���g����#���:��|�:��s>�.����׾�'	>Pa�}�۾k;S��4?�̾��e:(�)�96=�b����ʾz��=D�2>æ��/E1��V������1�I?+�:>S�����</�lg0>]�>�ĕ>D9����:���o��e�C�;���>�Q=�Z���� ���J�˩쾗؍>y�A?N�V?΁?A&s�_V_�K�;������by��#��P?�y�>��?�Ή>���=	���#��[�T��H�6��>�p�>���$�N�jƾ��!�
�f��>���>]�>�?r�]?� ?��p?��$?w"?�F�>�(<s�����2?��w?�Q�=�� �پ�]=���K�I?��2?�����>)�??g	=?BqP? \M?��!?�Y�>�P����D���>���>�^��a����A>}?5Q�>�ׂ?9o?E>�2��Y���ý )W�hK|>�k6?�'+? v
?��>�]?2E��e*
�r�?މX?(u�?93r?J��=��)?���>�hp>�H<c�>�3.?	vB?��_?
�`?(#+?P�>���<QE.��糽W��:��=@�M>����̃�қl�r߬<�Ș�� �;n�u�<N�e���#�m�=�%�=d9X='P�>jDt>z*��1�0>�žHY���~@>���Y���⊾�;���=�h�>��?�]�>�~#�3��=���>o��>���n(?�?:?��,;Ūb�<�ھW�K�=�>d�A?��='�l�Y�����u��Bi=��m?Jl^?��W��`���b?��]?{f�%=���þ �b�Պ龎�O?��
?��G���>��~?��q?ʶ�>��e�*:n����Cb���j�ж=r�>/X��d�o?�>��7?�N�>��b>�'�=�u۾��w��q�� ?i�?��?���?�**>w�n��3�\��������^?K��>�t��	"?�NĻ0�о�ˉ����x�߾M;�������U��m���C#�ׁ��ҽ#��=��?�3s?�5q?n$`?�� �#d���^�/��P*V�������`�D�,^D�ED��m�M��Ҙ��l����==
z��V�dh�?�
?I��<^��>�>^��N�6����s�=z�?���,���=�p���*4<�q�=I�W����Q��7�?�$�>���>z�B?�hP��!F��	E���;��(�9c�>z*i>��>�v�>Z���2���8�s����("�@�>�i?EK?�LT?�^���2�����=��=�=�!=���»���=n$)>�Ӊ�{v����A��Y�A���B��N���9A���"?�
u>�c?wɏ?���>u�����=8���a��=Z��>��Q?" ?t�>�罏��v�>�Ad?��?�=�>>���U`1���������J��>`f�>�?p_>?�3�zj��Џ��K��0k4�a��=��V?��k��1��G1>�2?�+���,=�
�>�ħ��*,��'�i]ӽ��D=IQ?7�6>���=�뾾�;���t�kr��(E?��)?!]ž8��S��>?���>�B?�~}?��+���ʾ���>'AE?��O?�C?��S?�-?|�m>��a�rڽ��I�9hR�֝�>EP�>�&�>I�4>��[��׬������=|F�=��{=�	�濽��Y���u�kP=]�[>�aۿ�K�@�ܾ'���"�ɝ��↾�b���o����
�F����l��M܂���,���M�bh�Ob���%r�W��?a�?H���Ɖ�+噿����N��n��>o�g��Ր�H���a	����CH߾�����#�v�P���i��Ie�L��>��ҽBͷ�
K��{f뾨"?�>E?��5?M�/����Ea�U�����<�2�P%������ӿˡ�����?��?����/;��W�>��>��=f��>57[����:��>�`?��W?:���Կ:�¿�|C>��?ap@>}A?3�(����GV=N��>��	?��?>�F1�F�(��T�>�<�?x��?8�M=U�W��	��~e?��<��F��ݻ��=C�=�9=�����J>�X�>�u�XA�G3ܽ]�4>�م>Br"����S|^���<ʊ]>U�ս':��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=u6�����{���&V�}��=[��>c�>,������O��I��U��=�E���ɿ)pM�t(���=ʇ=�9��`��г���;���;�hs�GY��o�=-��>푿>$yf>��E�& >�ZU?�Op?	��>�0�=Zac�~�+�"U�� ��=�Sڽ)�i�v��$}��}���˾V�ҾR�891��/�w�߾�t=���=�:R��b��$[ �̀b��%F�G.?�� >jnʾ�M��k<�˾Se���w��o���;�-2�5Tn���?�7B?����W�&N�'���G���)W?�����M/�����=���d=���>�D�=�}�q=3��S�y+;?׮%?�aʾF(��cw�>�����=�G?�/�>��Q+�>%U<?�E�<�����s>g>���>���>��=����G�UI)?��T?���@�e�~|�>����	{��L�=p}o>,�|�����>F{'=�����ns��?����/*W?Ҧ�>��)���T_��r��Pf==�x?��?&�>�rk?�B?��<0Y����S����w=��W?�#i?7�>���о�z����5?�e?��N>)hh����.�$R�� ?�n?�V?i۝�7p}�������3o6?��v?�r^�ss�����<�V�A=�>�[�>s��>��9�[k�>��>?{#��G������Y4��?z�@���?��;<�"���=�;?�\�>�O�\?ƾ�{�������q=y"�>x���zev����Q,�x�8?堃?���>��� ���!�=�Y���J�?�<�?�KM�`�9�|�'��Lt���Jc~>t��=Y��<�P����0���ؾ�ھ�_z�g-���Ɍ>�@H���w2?!����ѿ����W�/&޾��g>���>+ �>��A�w��(�X�,I���U�b�I������`�>��>�0���ӑ���{�ya;��ß��>���r��>�;S�P���3���C<��>H��>;��>j���� ��Ѻ�?�O��c-ο��������pX?'a�?�?'X?��:<��v�{�i�5G?�zs?�Z?Q�"�#�\��Z7���_?�`~���f��<�1�O��%N>�-?�>��/�׫�<M��<ju�>�\>�G��,¿/��axǾ�˪?H.�?�&��h'�>�+�?{8?(�7ܜ��H��R�(�b[1=|�3?RZa>�Ͼ��4�!�5�1F���?�0?�����1�]�_?+�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?_,�>��?���=�\�>��=x����2�xH#>2/�=-�>��?�M?3�>��=�8�//��^F�MER�,(���C�Q�>��a?D�L?�ab>0����1� !��)ͽX�1����pA@�[,�QD߽>D5>H>>�>��D��
Ӿ��?�ƾ��Կ�*����Z��d?�~n>3��>��	��h���c���iN?*4�>�,��n���ŕ����wR�?z�@���>3*��-a%��&>��>Ɠv>&�žz���Ph�x�>�$?D��w⌿������>=2�?@@r*�?�$i��	?B��O��b^~�Ҁ�1�6�4��=��7?D2��z>���>�
�=fov�E���.�s�!��>�B�?${�?8��>��l?�o��B�=�1=�J�>�k?�s?��l�+󾟹B>�?��������I�4f?��
@-u@�^?��Q#ѿ6����;-W����><|�=2i>wy�����=^ix=l�C=�A�=��>��>�V>�ۇ>d�d>�D@>*M>^����l%�����L��`q8��+�1��WtI���������S��aˎ���6�Y˽������r�?u���2�>S�R?�mM?Q�r?w�>,g�t6�=@H�/�=�_�2.i=���>��0?A:J?��$?a�=*����`��,��r���'|�����>��%>B��>�>���>n7.="��=�>�3�>�S>a�=���=,?R=�A>²�>�D�>�I�>D�2>��>�,��Oİ�	Xh�>�w�(�½|p�?^����J�%���������H�=8 -?s� >w����п����3sH?���4���q6�p=�=��1?KQX?��>������c��>nx�s�d��8�=�b���s���*��oO>�L?��b>��r>Ԛ3��s8��P�?����5{>�5?a���9�Hu���H�Fo޾��L>޾>s<��}�C&����~��h��y=>�:?��?L.��}4���uu��읾��Q>��\>^a=�ȫ=W�K>�e���ʽ��H��.=YO�=K�]>CM?��,>z��=d�>�����O�辨>�@>�.>{@?�$?���N��i�����-��;w>"��>�S�>kl>��J�䌭=���>Ѡb>{^�˯|��;�֨?�m;X>�����]�z�x��E{=ݮ�����=Η=9���I>��"=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ>p ���f�����|i����<��>2:?S���K������f�?"$?�l�5D����̿��x�J��>x��?0�?��g��'���<2�ͭ�>�S�?�f9?��y>����Ĥg�:��>��N?�P?�a�>J��v�P] ?���?	i�?\�>8̈?'�?���>;�����X�E7��.wf�^�����>�L�>�߼���ʓQ�~&���ŕ�JYw�L��Y��=鉤<9�>�Y�'����!>����UG^���|�[>Y�<�k����<>=��>7��>G��>R�=
9�����f��B�K?}��?����+n�=��<?O�=�^�F?�R4?�^���Ͼ��>>�\?D��?;[?	~�>��S-���޿�ot��@�<ogK>��>en�>f=���JK>��Ծ�8D�j�>Կ�>9��<1ھ�M��:?�� A�>�Y!?؆�>(o�=��?(�!?ɲ�>ɑ�>��M�� ��T�R���>v �>�!?I1~? ?:��Z�;�����v��%�X�v�E>�m?i?�d�>�B���V���ٸ�-��7��ߢ}?݋N?�J�dW?y?��=?:�L?y8>1/��+뾡B��{{>\�!?��,�A��J&��
�,?O?8��>P����սPpּ���R|��{�?�'\?OA&?���*a�� þ	'�<A0#��V���;m	D�7�>�>`������=\�>g�=�Rm�MA6�Vug<�s�=���>��=�27�3{���4,?�D�"郾Ϩ�=��r��wD�>�>�"L>����^?�=���{�G
���}���8U����?U��?�o�?Dk��ˤh��=?�'�?�?p*�>�a��nv޾`��w��x�a���>���>�Ah� ��܂��*���E��e�ƽ��,����>C��>�R?�>?��]>4�>�ꗾ��(�A���!���V^������7�'�/�=���q���J���x��^���`��5ڊ>�Q����>˒?|�>ii�>���>�>=yޮ>�QF>~u>��>z!c>_mX>��8>>��<%���NR?����'�"��t����4B?@qd?�I�>$�h��������Z�?���?r�?~Fv>loh�5 +�_q?�2�>�!���i
?;=���P�<F����������ָ�>��ֽ�#:��M�?f��h
?Q&?Z��]�̾vW׽jn��f|=�ˆ?�4.?m:,��U��t���W���L�9؃<o/`�NY����#�ۯu�d���]���Lˁ��G%�uw=8�'?䖉?�#�,y�aK��d�h���@�`kp>8��>D�>�Q�>��>>;U	���0�vN^�SQ*�gP���8�>k�w?E��>��D?.�4?�`?P�H?�w�>��>�hb�O?�"��h�>���>�G?�A?,s6?��?��?
�?>^;�$��q���־.?N~9?�`�>Y ?���>�7Ӿ���=�2+>d�|�j_�����)��=�+>�	��K@$��Mǽ��=[?����8�e����k>׀7?{�>3��>k���7����<9�>a�
?{I�>�����vr�P^�[�>Ϡ�?N�o=��)>�=����̺�k�=�¼�ΐ=|���R;�W]<r��=��=4u�곐����:a�;\G�<�5�>�?Q�>��>B����I�����%�=�Y>19Y>�N>�RؾXQ��f����g���u>�(�?8$�?�kd=��=���=������D\��ͽ�$��<��?�k"?�S?&��?��<??#?K>�q�EA��AI��%ޢ���?t!,?��>�����ʾ��։3�ם?e[?�<a����;)�ې¾�Խ��>�[/�h/~����4D��ꅻ���b��7��??A�X�6��x�ڿ���[��v�C?"�>Y�>�>O�)�y�g�n%��1;>��>eR?�W�>��O?��z?8�[?B�S>�Q7������p��֍��A>�??�I�?���?��x?��>��>%�*���߾���16�N������)�I=u!V>�L�>z��>�#�>x)�=��̽D����16��²=z�k>�S�>��>���>D�{>�<LH?���>�u��à��A�����<�Cv?v��?��*?�v=Y~�1E������>�_�?o�?6*?�T�H0�=GҼ褷���q��<�>2�>��>��=��C=�]>�~�>_B�>���_���)8�saK�p�?��E?���=(ɿ:~w��E�������0d������Z���)�~�־�>�"�ږ�]c�F�S�a���*�c������1{���%�>q��<2.�=#A>�.>3g���=LjP=�{�M��=���=���=L�㞀���ӽTj��cŻ��<�;�ַʾ�m}?�'I?7�+?sC?*#z>��>�9�㽗>$M��\�?GU>e�Q�Ж��;�������s�ؾ�
ؾ�?d�?����>}�B���>5�4>��=x�<|��=�Tf=��=;$�=��=g^�=?��=��=�>~>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�47>(�>��R���1�y�\���b��tZ�j�!?�H;��4̾�F�>~��=/I߾v�ƾ~/=��6>�a=^���Q\�Cƙ=9Z{�8�;=зl=	��><�C>q�=�#��2Z�=J=N�=��O>�ј���7��c,�D�3=���=��b>��%>���>\U?�[.?1�_?���>��k���˾Һ��zA�>���=�'�>y�=9e>^�>�{5?�A?c�G?ԫ�>�j,=<~�>�>��*��(q������}	==$p�?Ƀ�?戵>]m�<R�!��.�]�/�{Ѡ�S?��5?|�?��>�0�h��I/��1���O�� f��z�<��v��Ƚ+��!�������=g��>l�>s�>B��>�O,>��J>n��>��>��=R��=T=�<���<���&=���+ Y=��1<G|�����.l��3ɻ�������5\)�ɜh����=���>A>���>��=���^/>Z���x�L����=xZ���"B��/d�AR~�K	/�)a6�t�B>IsX>����4����?6Z>��?>n��?�-u?��>�8��վ0N���e�ʀS��N�=.�>r�<��l;��V`���M�$�Ҿ��>v��>E��>�tA>��6�*�>��}<b��3�0��>�ȫ�U޺��>$�O+���w���G��-[L����=F�L?Y����>�=`׊?��Z?"�?䔣>����ޡ�Fh>B������=8���y���gL;kG?��&?���>í����M�6Q̾�*��nַ>��H���O�����	�0�Y��䷾�W�>bݪ���о+03�c�������B��q�b�>x�O?��?�b�Q���XO����р���w?�g?i'�>�Y?�^?00���a��K����=i�n?s��?�4�?��
>�L=A;�.�>)�?I��?Q�?�Ai?i/��c�>�%���B>���A6��5�=�!�; �=S?�7?'�?�م�oj����	�ڛj�Gu���>�(�>�Y�>�N�>!a�>R�=��=��>���>_�>���>*J�>�0G>�ֱ��X.��0?Z��<�S�>:,?Nմ>���<`�i������G>z��E�����潤�R��|n=#
�>$ʒ>3�G=F��>lƿ�Ӧ?�-μ�St��G�>�=���Y��9v�>��6>/��<y6�>t_�>�l>e��>+��>�	�=�>J��=���j>[���i3��I��z<�9���j3>x5޾�dX��!�c��ʹ�v���� ��_[������_�ӊ��_�?fc=5�L�y>��4�h�?�}�>�?DY��ݗ��C����>4�>J���d��|�����Un�?�� @<7c>Y�>k�W?��?��1��3�itZ��u��(A��e�ݺ`�l፿E����
���n�_?	�x?�yA?dc�<�8z>桀?��%��ԏ�/(�>�/�%;�e<=�+�> &����`�ˮӾw�þb3��JF>͖o?�%�?�Y?gWV�_7N=�C>�,:?�N\?twn?�4P?	�C?M����@?���>�>�>��?2�/?�'>?�e?��>���=�����p/�0�ٽ�x���u�S�!�(p-;��=��=��=�8ƽ��%=Y�N=�[A��J��;Ԇ;T�;x>��ҥ=���=��>iɦ>�]?B�>��>��7?2���p8�S���R3/?ǎ9=����L������e�]�>��j?���??XZ?�4d>��A��C�)>�c�>ɕ&>�@\>/l�>]��J�E�tb�=�i>�=>��=��L�����غ	�������<�>���>]-|>}��:�'>�z��/+z��d>��Q��ʺ���S�Q�G���1��v��Z�>=�K?��?5��=�]� +��If��/)?(^<?�NM?��?��=X�۾��9���J�z<���>�d�<�������#��Z�:��+�:��s>�1�������:m>x��P$��m�+;D��Q�A�=y��]=n���׾�o���`�=w�>A���f���`��熬�oEK?ZS�=���{R�W�¾a,>�>�>G!�>9����;5C�'/��^Ks=���>�oC>�g��������N�<�����>~"J?��k?���?;�w����5�1��K�O����κ���%?�>>�?f�>��>_���
�	���U��-D��T�>�
?���u�F���ž>���.-A�!`>2�??J>�B?�\? �?� Q?b�*?�O�>S��>j������2?K��?Xk>�&���gR���"�Wq��U�>JYC?i�4����>��8?h4?��7?�V?�� ?�P|>����đR���>��>�d�������>@+u?V#p>;�6?z܇?�ȕ>AO-���N�'�����=c�>
T?��o?�j<?�n�>�)�>�3��ra>���>�?�n�?�]?�#�<��>{F�<0'?��j=�`>~�8?��,?�a?�]~?�i?5��>G��<�p$�����ٴ�������;Reֻ �y>�z��=�h��ұ<�@��(&�0�w���(����������<M�;�^�>��s>)����0>V�ľ�N����@>����xQ���׊��:�9׷=䋀>D�? ��>KX#�䵒=���>�K�>����4(?P�??��#;��b��ھ��K���>PB?���=H�l����]�u���g=G�m?Љ^?��W�%����b?��]?Ž�ę<�ľBDd��F�}bO?��
?�7H����>��~?�~q?&�>g�Yn�*����a�Ϙj��Q�=�>�h�d��t�>�7?�C�>� c>G1�=&�۾��w�pg���?l�?}��?���?��)>}�n�-2�2��֫��`�]?f��>�%���"?"��<��Ѿ�����F��k��Ń���:��9����^���m$�s݂������=��?Q�q?�p?�`?o��7�a��"^���}�[ZU���p���]F��F�OA���o�V�����\b����=�j�^�H�͛�?��*?��>���>e�C��S���*־�o>���ņ6�(</>{6��~�=�{3=	�[��n4�\u�
?�O�>0��>�9>?�A��T5���*��0�����g+>�:�>��i>7V�>�ͼ�'>�5	�6پ������<�>��O?`sF?ƾf?���'�8�W8�����(�< -۾F$>*�>�@>�!9��Z�Rl�e�D�#�O�z�y�~�	�� >�p?[S�>���>ȑ�?u?{k���Ծ�n���	���z=���>���?Rv?2.�>����C�<���>F?f?�[�>���>k��L)�O_~����>���>�C	?n\�>eaX�EZ�� ���Ì�N�;�� >�h?Zv�z�S�Ɏ}>4�G?&�;-���c�>y'�@��{�ލ_�@4�=� 
?r��=�m>�𫾀#�<<r��6��t�)?v�?4ȏ�/+*��*�>\J#?<I�>�Y�>T܄?W�>ʿ��*<�?]t_?�&J?h�B?�^�>O�H=b̸�Y�̽\�(���%=�Q�>��`>?�=G��=it �%|Z���[A?=
e�=-ϼ<����5<R*��I��<�=g�>>W�ؿ*�G�X�۾�x�ra޾,��� e���N�b:��򹵽n{þ����(�e������ �E�J�H�x����k��?Vr�?����R���ӝ��T~�T���m�>�Y��A�f���N�9��z��A�#�Q� �&<R�,n�y1g��%?�4f���¿�B���3���.?1�7?�9�?J�)���/�NA5���%�H5ѽFμW�����ӿ̛Ҿ�P?���>���a7=���>�r�="Y=<ԭ>��G�3|ؾ�|�� ?��?��>���:Tǿ����k�;[��?	@�yA?��(����=XV=���>P�	?E�?>i1�!D�S簾K�>�6�?I�?�L=��W�s�	�V}e?�9<P�F�T�ܻ���=ob�=�=���&�J>]�>h���YA��ܽ��4>,Ʌ>Xj"����{^��*�<Xs]>��ս#��5Մ?,{\��f���/��T��U>��T?�*�>Q:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�z��=[��>b�>,������O��I��S��=Y5�ʿ��L���<����>�̆<֪;��r>&�_>[?�|�Ey�:�>��軍�&>y��>��>�s�>�c�=�:=?R0G?|`�>�� ='�#=�N�f���׭�=;���VÙ<3��(�Oqe�n�����A�m��cu���	��F@�ق�=FuP����/'�~8�\m/���:?DQ>��{��^e��ؐ��Ǹ��Ə��Y=�N������7����9k�?��\?,#���}_�^4���ǽ��P���3? qu:G*���ubX=`i޽A�:jI�>`�={��@;U��NK�D�0?#?{@��%c��G�)>c�k�=@�+?�6?O)2<��>�o%?��*�h7⽣�[>Ű3>��>T�>��>vH���uڽt?�JT?�� ��Ꜿ���>ý��W{���b=ޥ>�5���ۼ�x\>��<~n���EA�}�Z��<�(W?Q��>C�)����a�� ��Y==�x?m�?.�>p{k?��B?�Ѥ<�h����S����^w=��W?_*i?��>򈁽	о ����5?h�e?�N>�ah�w�� �.�?U�$?�n?�^?Pw���v}�I��i���n6?��v?s^�xs������V�^=�>�[�>���>��9��k�>�>?�#��G������uY4�$Þ?��@���?��;<��V��=�;?i\�>�O��>ƾ�z��������q=�"�>����pev�����Q,�a�8?ؠ�?���>������v�>-=��t��?jM�?a� �o�=l$�B�q��7�~�=��=@E��m�=`��v��a?ӾY������v-=�p>�@gk����>#�<�ɿs+ܿ))����ľn���`�)?tF�>^8ľD :�fX��Ʌ�E�)���ؾL�>�>��������Y�{�	q;������>J
�
�>�S�&��星�eo5<��>���>���>K(���潾�ę?�c��?ο��������X?�g�?2n�?�o?A�9<�v�"�{��J��,G?��s?�Z?�l%��=]�G�7��j?4_��0U`���4��HE�U>�"3?�B�>��-�.�|=�>��>&f>�#/�}�Ŀ�ٶ�n���
��?։�?�o꾧��>d��?�s+?ki�8�� \����*��+��<A?�2>n����!�@0=�LҒ���
?o~0?�{�F.�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?���>�N�?��>�H�>�n�=_��I�߻hF$>���=,օ���?�KM?��>:��=��.�m�*�x:D�SO���nB��T�>�-_?��K?<�f>$gҽv� �ZV ��ս=#�>��I��qڼee½�o5>V�:>TI>=iN�r{˾��?Pp�9�ؿ j��p'��54?(��>�?��o�t�����;_?Vz�>�6��+���%���B�_��?�G�?>�?��׾�R̼�>?�>�I�>=�Խ����a�����7>0�B?A��D��p�o�v�>���?	�@�ծ?ji��	?���P��Va~����7�[��=��7?�0�%�z>���>��=�nv�޻��W�s����>�B�?�{�?��>"�l?��o�O�B���1=9M�>Μk?�s?1Qo���m�B>��?������L��f?
�
@u@a�^?*�|п�~�����=�۾V��=�M�>4wS>h���9�=��μF=�e�=	�>G��>�*�>�v�>an�>�S>B�=>h��q�'�¿e��~W��D+�����=<��۾2D��n#��i��v���8  �O��=U=�����0��e�L�]>�;>?\�Y?i�l?"��>4S1�a;(>@����������0O>�A�>�H?ԦD?uj?�-�=
!���F�����\��W6���>L��>���>H�w>n�>�[{�k��=��p>��>��=_�A>�>��=�3>���>�ה>i�>�$>�V�>*���븿�pd�a#��":[��١?�c���7�	﫿@�ʾ�e�6l�=y�4?�x�=�x��5n�>���V?�吾��2�i=�N<��0?`�U?p��>Sb!��cU�x�>�L������Q=��|���V0W�4)>~.7?��f>�u>�3��g8�;�P��j��8�|>�=6?o���w\9�]�u�$�H��mݾPBM>XǾ>6�D��s�5���i	�-gi�<z{=={:?�?�g��G𰾦�u�(;��)R>�-\>D�=+]�=�[M>rc��ǽX'H�[.=P��=��^>�K?��>,�=�d�>.����X@�&��>E�(>�a>SjB?xK?��k�����Y��0i��vk>���>�'t>f#6>�5;���=u�>�Qr>���;K2|����P�;���E>�t�X�[�L��LU=�Ѳ��	�=�Si=���oN��3�<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾;`Z����>һ@?�R?�>�9�~�'���?�޶?֯�?v��>��?�_?^]�>o�(�M�5�i���_����L=�m���>`f>�s��I��X��|���il���о�>ףx=`;�>)�ҽ4���7��<��*�첾��Q=�5�>+t�=��=��y>��?��>���>���=�O�A��)z��f�K?ʲ�?c���/n�Z�<���= �^�<&?�G4?%�[���ϾMר>��\?���?�[?�c�>���P=��迿�~��X��<��K>14�>�H�>�*���JK>��Ծs6D��p�>Eҗ>9��";ھ�)���㢻�A�>he!?1��>0Ԯ=�&*?;�?{�>�k�>��7��b���h;��e>>
�>�y�>u�?���>	��_q;��A�����YWe���w>@8y?�}?1�s>i�������j�ʽ�3ǽ{Ի#tx?#B[?������?Kd�?��5?H�6?�WJ>t�4=mO��Q���ɗ>A�!?�X���A�O:&�X��|?4e?6��>\|��qqս*�ּ]���>����?`,\?�6&?s��%a���¾���<�#�]�J�n�<��?���>5�>����U�=>LҰ=I~m�[T6��e<�-�=�k�>b��=�K7��Ȏ�0=,?ؿG�}ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?^��@�h��$=?�?S	?n"�>�J���}޾6�྿Pw�~x��w�Y�>���>+�l���K���ڙ���F��a�ŽP�0����>r-�>D?�^�>��=�1�>fI��'?�9��gժ���T�9�%��,�&�0��6�?梾�! �[�<Luƾ�C��$o>9R �!�>׋&?���>��>v��>�6
�/��>R.>Lѱ>���>��>��>�*>�+x>�"½�KR?�����'�%��ʲ��S3B?�qd?1�>�i�������`�?���?#s�?�=v>�~h��,+�gn?�>�>(��2q
?bV:=w2��@�<�U��(���2��S� ��>�D׽� :��M�^nf�bj
?�/?���Ӌ̾F<׽%�:���>��?l|0?!ھ��0���z�'�y�Z�T���*���뜾tq:�J���9�����������Ծſ�=�'?̧p?������
��ھ��D�x��\>�>��>��>k>�8�<��n�e4�� ��C�>fe?2:�>Y�_?N0>?y�8?�_Q?:	�>nLx>��Ҿ�!?�*�=I�>�W?��@?�-H?ŝ4?�-?��O?��>����6��̹�
�?D(?[�?�"?)o?����Y��_k�<�)�;4��˩�q�>��I=���������=�r�>,[?n��q�8��}��Ԛj>�b7?���>p��>����
����<�>E�
?3�>� �uor�2c� <�>���?i���H=�)>�,�=�ჼ1A�p��=�)��d"�=�m��=;�[<տ=) �=� m�h�j�{��:��;dޭ<�u�>+�?���>I�>$7���� ����=)�X>S>>�Dپ
��%����g�*y>�q�??y�?�f=q3�=|��=����Z�����5����2�<��?/H#?FPT?F��?��=?�^#?�>.-�QK���]�����خ?�h&?���>_a	�^a޾�1J?��/;?�3?�����c\�j�'�$��
g0�i6>|h8�7���Ȫ���_���8>	{
�l���*�?y$�?�`��8�v����!گ� ���oK?蓣>�M�>`?��(�WO��ޘ5���>�R�>�<?���>�P?�{?�L[?iT>�'8�����������@!>��??W��?VЎ?q�x?x�>S>��'���޾�����T!���{����V=�[>r�>��>54�>�M�=�kŽm��4'>��S�=zc>j��>���>���>�=x>�÷<��G?��>ɤ������Q��g����QE���t?��?��+?�=+��C4E���.��>y�?! �?�*?gsT��K�=��ڼ�궾)zq�&��>��>��>Pʏ=�CG=K�>ޖ�>gi�>�������68���K� 4?�LF?�c�=C�ſ�z����cU����=���wK��-0��+J���>�㳾�p��ky��Mxy�A����t��Д������`�����>�3f=|�>� �=��h=�hQ;�l�<�JX=(����=��@�kо=��Q�67=§��j�ɼ$;�<DY�=~��� ɾ�|?�I?��+?C?"�v>I>��.�x7�>ݠ���?��X>'=L�=ֺ���8�!k��@��T�׾#پde������>I>�P�>X9/>%i�=��s<���=��}=�I�=)ͻ �)=hW�=���=�U�=���=��>�u>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��6>��>��R�wz1���[�߾b���Z���!?��:��˾��>���=-�޾i�ƾ7'.=��6>U4e=����;\�p��=o{�_*==�^l=1�>׉D>A�=}"����=�bM=t�=q�P>_��3�`*+��M3=�Z�=�b>�%>`��>
5?�0?wDd?�Թ>1bn�1�ϾUi��3��>�b�=���>�S�="uC>��>8?6�D?��K?�p�>Շ=���>6o�>��,�_n�>�d榾���<iz�?yن?���>õK<�@��v�f<>��EĽެ?�1?�?l��>6��@ܿlR�5wA��R��\Q��B�=�
�n=B�Ǽ�*����>�=�p�>9�>tB�>�F�>�c�>3[�>ڜ�>d��=��.>�we=�~�=���:���eZ>t��=^<:>:A;�l���=I��l�;�`��=�]�/J���=���=���>t<>��>2}�=A��2?/>i�����L�k��=�<���)B��5d�&J~��/�0f6���B> (X>�m��33����?��Y>Bw?>��?*Cu?��>�+�`�վTQ��� e�{QS�'��=R�>��<��m;��U`���M��|Ҿ�e�>i=t>N�>��u>�lB���e�Ŧ<�D��� J�Z&�>�҄�������S�Y�p��h����fDX�ɉZ�W�>?B����(}=q�k?��`?Z�?!��>�����,��>�l���s>RPؾ������=�k�?��>?���>2kb���E��.̾㾽z�>�I�0�O�+�����0� ��շ�!{�>�ߪ�s�о�33��g��)����B�#zr����>��O?V�?�8b��U���JO�����
��?u?�sg?�(�>�@?H?����u�<Z���X�=��n?���?r4�?F>�ڿ=� �����>3:
?+��?��?0ws?S�E��V�>[>�;8(>Ĕ��C��=�>]��=/5�=ع?�?td
?
�jC�X���L�j�\�8�=��=J�>@�>O�j>x3�=Z=�ğ=^Q>в�>�ݒ>ppd>�6�>��>� �����h?��^>S�=ߏ?t7�>�ڍ�?(��To=�
_�<�=��=�tB��L�<fV.=�Xh=��=��9>�U�>�¿�H�?��u>�o���L?e^�ތ��:7����>b|���>�u?����?�>�<>9>8�>�CӾ�>���ve!�%-C��R�C�Ѿ��z>7���t&�9������II��n���e�'j��.��X==��Ľ<�G�?c���\�k���)�����X�?�_�>�6?�ތ�����>6��>�ō>pG��-���^ȍ�%i���?y��?�;c>��>D�W? �?Ē1�G3��uZ�+�u�i(A�(e�@�`��፿�����
� ���_?��x?+yA?IS�< :z>L��?��%�Wӏ��)�>�/�';��?<=+�>*���`�s�Ӿ��þ�7��HF>��o?3%�?|Y?(TV���S�4�)>:i;?4�1?��s?�u/?z�:?�7�{�"?f�*>'�?�
?kp4?Gv/? �
?ש4>���=I˱�;}=������� Ͻ�̹��9ܼ�-=��=bӆ�'ι;t�#=��<�i�)���"��;yʙ����<}�?=���=w�=��>�c?wt�>,~>w�6?X���;�����c5?M1i=u�q�UOl�	C����߾�I>�%n?t=�?�O^?/S>��F�`�G�]�>�ĉ>NM:>�N�>��>r��J�?���=÷>�[>Y̠=*� ���~����9��h�B=OIA>�:�>�	X>��I���<>����g�4�>�]��}��x�9��eE�I4��`F�Ef�>��L?��?���=�%���"��b`�	�*?�;?�GN?P[�?[�=����?7��I�?�'��L�>�4e;?�+k���袿�:�跾�H�l>�	��O!ξ�x�>�=��٥��Z�b�K�n���6��Ծrt �v�<�� �*� *=����cgR�<����.�A���#���tM?��v���޾�r�������>\��>�O�> [}����HN�j=��'��=W�?��+>h5d=�~��"#�?�+�N`!>�?�Ai?ucj?ˇ���y��6�L���ޚ�[�=p&
?���>���>a�>��=a�ҽ��ky��a����>1�>���:a�����t�0�ØJ���=��?�8�=`?���?<�?y[o?��$?�K?���>6x!�Alξ� ?Dcs?O�y=w0����O�qfT��V��x�>�?�qT�s��>�Q4?�*?lo3?�$O?'??0=>���g<T�:*�>�Z�>�c�D}��]ڡ>A�G?��>�O?J�?��=H4�$����A���:ok5>D=/?��7?��G?Ȇ�>���>�v��W����m>��?�X?��:?��=�J?�Wϼ���>�(�>2d�=.F�>�b�>%�4?�k?V-_?���>��=x� ��j�^��;����O=�V�=N)����9����=n|c���t=g��^�D;����(ܧ=��=7��<�E�={�>$xs>AI���0>�e¾�@����@>��������U㊾�%8�%�=��>�?P��>;� �S��=���><��>�S�܏'?Z`?�?9;�Gb���ھ�aJ��ް>�A?43�=<�k�1��K�u���h=Qm?��]?��V�St����b?�^?�P�#=���þ�b��w龖�O?��
?�G��>��~?��q?ӻ�>��e��4n�0���3b�|�j����=�g�>QD�E�d�6?�>�7?=�>p�b>T7�=�e۾βw��^��*?1�?)��?R��?�*>U�n��3��� ��㕿�`?���>Ҝ��gc!?�}�<��׾�ۚ�8m���jž-���fO��q-���gF����e���=�?Z�s?$'v?q^?����Ier���^�'�|�x�X�oy�����:^D��E�=A���l���	�rE�����
=0D��lEd�w,�?��*?�s���b�>E��<�y[���ɔ>dz������Gq�>�����=����	���=�(���a��d(?�&�>L��>�9?��L�=S�/�#���<�S��a�>)YY>z�3>j�>	Z��.g�e��n#���h���ɒ���>�M?l::?�[?2�4�N�?��T��8�+�W��������=� ���>-?6��=n�d6�'�=���p���J�G1x�_����o=�R:?�&>��>{Δ?�>9?r=���������-����L>�K?/�?�
? �K>����7?����>M�l?;��>��>@����Q!���{�Rʽ0�>�>���>�p>f�,��\�2d��,���9�i��=I�h?�����`���>GR?���:5�I<�k�>w���!����$�'��>��?��=}�;>��žN(���{�Y����8?��?�p���"��ܘn>���>���> ��>�R`?��>����l�=�)?��I?I0?A5?��>6�> "��8���S����=$>Aw>;�=�h>2A���
`�uA5���(<�IR=���'�'����<�0���E�<��=Y>�@��x�������$�D:��
����ؾ*�;@���V�<�c��Te��^��x� �;��V�ІX���˾�h���?j`�?3tx���ؾ3���Gz��6 �uX?�����r=��0Ͼ^�v�n�о���ݙ����1�+��('����m�_��>����Ҕտ�?п@��a�>L�>�C�?��`�A��2�m�`�h<�c���}��>������ݿ�¾a�e?5K�>�hӾ2@����?��K>�_R>���>�y��/1��`�;�N?1�?B'?�0��s��ο��P����?/�@�A?�0$�T����,2=�*�>�?�}Q>	��v��B��3��>���?ގ�?N{a=�Q��M���c?M�9��<�ͳ����=j�=!g=�I,>��>� �d�C�dSս9�,>Q��>��#��3�E�Z�c=J�f>���&Մ?z\��f�C�/�aT��gV>)�T?3*�>G;�=U�,?�7H��{Ͽ��\��(a?o/�?���?R�(?�ۿ�-ٚ>v�ܾ�M?�B6?���>�e&�*�t�J�=�W�u0�����@'V�r��=��>�>�},�(��j�O�d;��0��=�����ӿ�H9��(���>s.��pn�����ߣ׽�S=gT�F�0���w�)��:��>UH>=K�>HR$>`>�pK?"�e?v$�>�%>t��𰉾�Rо齌=Q�s��Wb�is��C�)�����D��,�־���p�0�W�"���Ӿ"�V��ꄽΝF��駿r�,��r[��ld�7�T?Lb��0���։�9߼��� ��zd=�)	�=A	��m��]l�F�?)�t?F�|��Q��ǯJ��m=�ɳ';? �?�Q˾|�����σ�'D�Ѭ���>;TR��	8� �*�}A�v�C?q�*?Z���]yн�>��|�qƾ=��?F�	?���=��>j9?]�Ҽ� ��|>�zR>���>�w�>�yb>0��ܼ$�I!�>�&T?�����ѣ��>�쑾C7�?�=Pc�>��.�O�*>�`>%$�c��(���,�D�q�S�Y?�ߢ>Z�$��,��g��=�'�x�n=��w?�u?���>�8j?�lA?�<iU�
�L���ǝ�=��W?{*h?_�>�<���!Ǿg㜾Vk1?9Tb? H>t]��?�wk+������?T�p?��?��̼ ���㩒���k�.?s�v?�o^��o������V��M�>�h�>е�>n�9��n�>7�>?�#�JA��o����T4����?��@&��?a=<fP�䑎=rC?�j�>XzO�Eƾg���s��J�p=�	�>C���pv�6���,���8?o��?��>�v��T������{ʾeI�?�߆?F����L	�c�O�q��_ �Y��=����㕾@�=��*��	$��}���"�/K׾/�)<QP>ѝ@#�<0�>��:=T���*��h���fk��׾5?�m�>��澮�A�O�n���;��-��fp���˾{P�>1�4>���ſ��b�x�n�<��������>첵����>�$:�ô��l���#��<l�>��>��>�������Lś?K�޾"ͿZ_�������S?�]�?2Y�?�Y#?79?=��l�o�s���;dVA?��i?JT?��K��;P�)AD���j?l_��^U`�Ύ4�HE�U>�"3?.C�>6�-�o�|=_>y��>Mh>�#/�T�ĿZٶ�����
��?щ�?�o꾍��>c��?�s+?�i�8���[����*�+�|<A?/2>�����!�e0=�
Ғ���
?R~0?L|��.�]�_?'�a�K�p���-���ƽ�ۡ>��0��e\�N�����Xe�	���@y����?J^�?g�?ʵ�� #�d6%?�>Z����8ǾL�<���>�(�>�)N>�H_���u>����:�i	>���?�~�?Oj?���������U> �}?Y*�> �?��%>2.�>*A�=���:�<�C>�1>�3-=�y?`�V?E�?X�>=���k(�95<��_7��o	�]f;�ng>hk?~CD?+�c>o��5a��}t�Y����)�~�v<���O��z�^;F>Kts>��>s�Z�G�����?;p�3�ؿ�i��_o'��54?c��>�?����t�����;_?xz�>�6��+���%��{B�L��?�G�?2�?��׾�Q̼>*�>�I�>��Խ����G�����7>�B?~��D��}�o�i�>���?�@�ծ?xi��	?���P��Na~����7����=��7?�0��z>���>��=�nv�ڻ��P�s����>�B�?�{�?��>�l?��o�G�B���1=/M�>ʜk?�s?�Po���Q�B>��?�������K��f?�
@u@c�^?%��̿�Ԫ�N�y��W�k>1=�^��W������j��>�h��Ƭ=;H�>�ɼ=3N�>�/z>�ɖ>��=YG>���
q%�����;��.�ǾC>�2�(����Ao�}�����j��D(��i��
O��nļ|ý�҅��z��|�6;isB={C1?�Q?T�t?P�>R&����=�*ؾ��<��s�k>B=)��=�`?�">?�	?G�6='~��OP��j���,���g~�o(�>yz>�>���>���>C�j=��=�L>{z�>�T�>J���͓�ae�=?�>Bw�>|��>Z8�>�g6>�F>�ô��b���Qi��Xx��սJң?�����	J�2G������������=�-?s��=�����пC�����H?+�������51��(>��0?��W?��!>�ִ�}b��>��L�j�c>*�66z�W,*�-1X>��?�i>g�p>?o2���6�`�P�G%����y>�g4?@W��b�8��Ju���G�_۾�M>�W�>��vN�����}�/f�]=*�9?�5?-׿�/簾�-n�w7��A�J>�IV>=��=,�O>�xV������G�[y=�S�=KUY>�?���>�CS=Q�>gׇ� ���g�>v�X>ㄆ>f`D?D;#?�+�=��K�I��ƽ%Ԉ>��>���>ؠ>ϭ&�Ccz=���>㱅>?�`���n�F�=���,>5C��Z�6��r��D��=8�[����=��3%6�91�P ��~?���(䈿��e���lD?T+?` �=�F<��"�D ���H��F�?q�@m�?��	�ߢV�?�?�@�?��I��=}�>	׫>�ξ�L��?��Ž5Ǣ�Ȕ	�,)#�jS�?��?��/�Yʋ�;l��6>�^%? �Ӿh�>�x��Z�������u��#=J��>�8H?�V����O��>��v
?�?�^�ᩤ���ȿJ|v����>K�?���?a�m�{A���@�d��>*��?�gY?�ni>h۾�_Z�勌>��@?�R?��>�9���'�h�?�޶?ᯅ?��0>\��?�q?���>����4�dn��H���|�>=C��;Uق>��=3�־-�F������Ĉ��i��=�w�>#4K=�>��������N�=�DT�.������)��>3j>��:>��>eg?���>MZ�>r͘=^�����j��̓��L?���?���m�é�<�,�=�g^�p*?�U4?�M�xϾ�*�>��\?z��?��Z?5P�>������ۿ�O������<�ML>��>�?�>%����J>��Ծ��C��>ת�>@�����ھ�5��i^�����>aj!?�[�>���=�� ?@$?��i>�n�>�>E��4����E�ց�>��>z?!�~?Y�?�w����2�G���V����[�ӦN>-y?L�?zA�>`����m��&�D��XI�&���w�?��g?#�߽��?��?z�??k;A?ed>$��Rؾ�@��I��>�t*?����5=��x���(�� ?)D?���>ki�bU��>ס��
�^$پ%� ?��P?�l'?x�澠�O��ॾ�7=<��<k�;Ƀ!=�6��캡=�>��Ž���=(�=o=�7��N$��V�:߶='`x>#�=���\��s=,?k�G�;ۃ���=��r��vD��>�JL> ��F�^?�h=�e�{�����w��U�� �?���?+k�?���؝h�$=?��?�	?o"�>L���}޾���:Ow�;zx�cu�h�>���>��l���\��������F���ƽD���W;�>Ɓ�>|S�>=�_>��=�U�>�	��[�)��f&�tz���X�����Q���,�9�����aSK���[�����yY����>��j�?v?75{>��=�n�>�ǔ<>�>��>=�>���>6]>���>��=�=�����<R?,�����'���2���~`B?�nd?J!�>0�h��m��E���R?���?
U�?�v>,h���*��5?���>0��#*
?�X<=_s����<�k�����:��k��]��>M_׽�~9�5�L�r�g��6
?='?Q���C�̾�ڽY���V5>ܝ?X;	?���3��䧿�J��>e9��,�W߽c5���[�m∿Ԛ�7{�� ����_���"��!?]��?#�߾sP��D���+�P_�렂�֖�>n�>_�>`��>A�*�N㾬T��Pྞ�W��c�>B	?6��>�b1?�0?dI4?��2? ?3>�נ>�Z��m?�G3���>���>z�>�H?H?{W'?� ?���>i�1�T��
��P ?%*?c?��?1��>�R��� �V͞��,�, ˾'���
>Go�=�����G�,:�Ao>�!?��齿D�����$�>�GR?��?ח�>o]}�I̐��{=3֒>�4?l�>�Ҿ�2=�~`�
A�>٨�?_ٻ+�<&��=3[�=��<R�>�.�O=3�?��=�L�<���<k�=�>�=7�%=�^ܼ�=���=CQ��[d��z�>f�?G��>E@�>?��a� �F��cz�=Y>�#S>Y$>�;پ�{��� ���g�by>+v�?*y�?�g=!�=��=�~���J��������O��<2�?+H#?]RT?���?��=?_j#?Ʒ>�'��N���]�������?�a�>2u>?��N�!�r���bq-�Q��>7�:?�b��m��Un9���۾˜�������AH���"¿W>#��`�> �<�Ͻ���?=�?6ۑ�pIK�l������n�|�޸?-�>�J>�H?�,��<P��'���>���>`�I?>@�>�C?.2[?�^T?��k>�=�J!��F��\�;��=��D?LB~?���?>�x?P��>�o@>��Ľ�����J���7?�$I�Gq���<5=��R>��>�A�>1�>�A�=�+��󛺽�S�����=��^>�(�>�×>
i�>:Hy>��v=VR?o�?0ü������dD���_�b?�M�?�`<?��=CL�#�?�4Ѿ�>g�?��? I.?���H,J>� '=Nv��yQ:��-�>WL�>nz�>{$�=F��=ea?>���>�9�>a�����4���?��5?x7B?D��<�¿��m� Z����~p��o��.e_�p�����c�W�=Y斾��!��~��
&P���腓�����r����J�� ��>˄�=2>,g�=yc=d;��$(=^�Y=B}C<�0,=�HG�UV=��G�8�ռ�q��	T�<�e�<��d=�9/��ʾ@7}?}@I?=�+?=�C?�g{>��>�C.�T�>L�����?<U>JM�����<��Ч����Īؾ�׾8 d�<��u�>�oJ���>H3>b��=/m�<5h�=<�q=G��=p���'2=��=�/�=�=%��=�=>!)>�6w?V���
����4Q��Z罡�:?�8�>l{�=|�ƾm@?��>>�2������pb��-?���?�T�?>�? ti��d�>?���㎽�q�=�����=2>3��=l�2�W��>��J>���K��a���~4�?��@��??�ዿˢϿ'a/>^�L>_b�=�S��%���N���p���[�vi?i|1�	�ɾR�>:�=n��Ö�����=��M>Cޢ=z���Q�aǇ=��t�om8=��Q=�1}>�C>*H�=�\��
$�=��8=�m�=>N&>��/<�'6�ؔ1����<,�=�yc>E >��>�\?!_?�"?��>`6���ƪ�cP���-�>�5'<���>Z�K>�ɧ��^�>�-?k�G?��L?��>��\>}�?���>k�Z�@MW�q����3��1� ��kx?6$k?|�>���=�=^�_I�l�v9��*a�>�(
?E��>�P�>R����w[&���.��}��̎G��5+=Efr���T��[��9S�;�����=r�>��>��>SYy>�:>��N>t�>�>'�<�G�=l닻�ö<ʷ��?��=����v�<��ż��+�#���+�G��Wz�;�b�;�^<d��;{��=P��>BJ>,��>5k�=V��AD/>����A�L�
¿=XF���*B�k3d��D~��/��R6���B>�0X>s����1���?L�Y>�c?>i��?�?u?r�>�-��վ_N���8e��LS�-��=V�>��<�*l;�CW`�8�M��pҾ���=H>���>��d=����T�E#4=�&�F�t��=�پv���N*��AҶ��a������,s�R�k?�댿IE>b�e?IKR?��?���>�~=�D/�^�?Of��"�=)����Ӹ�0�>9_?�_V?!�?cS�~x�٘̾�ݾ����>�9I�pP�
����0��!!�\ٷ�w�>$�fѾ6"3�Af��������B���r��Ӻ>��O?M߮?R�b�H@��2O����S����w?�Ag?�>u?�8?Aj����M����ù=�n?(��?�"�?�>׬">?�4��]�>G��>��?�Ŋ?[�f?4W��7��>��6Gt>��_�Ӗ=yk>d->t�&>
�?q�?�d?о<gK�)�3=��͌���=�)>���>΄�>��&>��U;�E=]B3>���=�,�=&�E>w�{>�ư>�K�>���%�T�#?�	>�9=�P?�+�>Bd�<�1���Y� ��������q(��ل��Q��G�+u3�a�=H����>�]пZ̉?Xj�>^� ���A?rm��vꐾ�t�=��&?�����P>���>�W���?���> >��l>bȜ>�T�!t�=���+�P�Y�O�SN���T8�>9AѾQw%��m2���-�tT}�i��l���o�*[����T��̼^��?�3�D���5�J��h?�Z�>��:?#xƾ�M�T�\>\��>:�>}>ᾀ���p蠿J\���?^��?Y'c>	j�>�vW?�Q?|00�=F3��RZ���u���@�U�d�iG`������m��vR
������_?��x?(wA?�ݜ<y�z>��?�3&��1��*d�>�/�qs;��?=K�>ư�I�_�!�Ӿfoþ�����G>�*o?D�?�E?��V����>��&>c�?Iy??�~�?,i?��4?wn=�F0?�� >oȼ>`�>7�#?-�5?���>�B>�(@>'�N���0���cͽ�R=�;B�:�)=�_�=S�l;�I��J���Ӻ%V��O�D��u����<�f-;��;=1�=�ߥ>�Y?���>��>wN6?�A5�v-��ң��*?��;l�G���u�K͠�_�¾��7>��i?H�?��]?��_>QE��DU���=\˗>	�->��Y>hI�>1ཽ��U�=��=_`>��=�=�)����`�~6
��͍�{�m;v1>���>�|>[��5�'>�c��<�y���d>��Q�G�����S���G��1�mv��U�>��K?��?`=�='�c���9f�$)?�K<?�RM?w�?�v�=��۾��9�U�J����]�>C­<
��г������:�/�d:�@s>Z��l䘾�|�>h��V����h�3[:���߾!�=�D�\2�=u��g�ܾPX^���=�j%>B0���y��r���'��ޏM?D�=iSʾ�V��ƾw�B>:P�>n��><䨽\���4�E��W��,��=���>��.>t�ż֬���S��h�^1�>��?�/S?-��?�`Ⱦ�X~�=�l�&��ڎ�k�";�GH?w�?��?]Ԝ>�q�=��ݽ���O�]�u�I��E�>ـ>�W����H��⸾����(#T��M >���>g&���=?Q�?�L?ʞQ?��/?�K�>�С={�I�$+Ͼ��0?��o?�@ >=�U��9��$7��X����>�N-?/	��R��>v�?|?n*9?7N?��?p�=��	�"�R�겉>�7�>�O�h����U>џP?~�>�U?�]�?�Q>��>�<�۾�=���7�=e��=�,?�3?�,?Y�>O�?&���t?	�U\�>�0C?�b@?B��?�sG>��#?�Fݽ�~�>A�?1��<?�?D��>��z?��?�߂?�?��W<�Vƽy��/�(��R =�lx��O?=o��=���=im�<eM��q�<��Y�����۱�����l�<�j�;�E�=���>��s>����9�1>C�ľ4I��~�A>H������1݊��;8�|W�=�4�>>?Sq�>ҹ!��ؓ=V�>��>���m�'?�f?l�?*U;�b�g�پ��K�3��>ǽA?���=Al��p���av��Fi=�m?T^?&[U�5U����b?q�]?�V�
=��þ��b�S����O?z�
?#�G�L��>l�~?!�q?x��>��e�x2n���Fb�P�j�l�=Nm�>�T���d�5�>՚7?�:�>��b>�f�=4z۾*�w�z��5?��?���?��?�5*>��n��1�i��%����h`?wM�>�{��3�?��%;{qҾ�i������������(�ͤ��k���I�)������ҽW��=!?V�o?��p?S�c?����mjh��W`�����>X�=�;��A��wB�xGF�(m�,G�����������6=E�~�K����?�t?�����>�*��f¾"�Ѿ+��>��ƾ�,�Y�=MN�
�;>�p�<ư���
��H��Y)?�O�>�O�>n$F?QeF�9 P��;,�!� ����cwt>�Or>���>we�>'��RϽ9��[Ҿ��\��7�>��q?�je?�l?MǇ��JK�ꉿ�$)�5�2�h�ֽ��(>5�S�M{�>����-�)q-�k@0�>�|�j�=�}� �#���,���d?��#>��>��?K�?���[�Z������$�:Mt��'�>�R?�E?d�>μ��̾y��>��l?%��>��>����J^!��{���ʽ"�>��>��>r�o>ѣ,�I\�Si��􂎿69��C�=��h?�����`���>�R?hن:%�G<Xt�>��v���!�H�򾜻'��>�}?���=¡;>�už��Π{�\0���+?j+?ߒ��w�"��&d>8�?@�>��>
?�5�>�V��L��<)Y?�a?ݜG?U�A?���>�xe=�Lѽ�ڽ��w-A=�Q�>-)e>ԟ�=t��=���b�p�,���E{=�;�=����=ʽ�rx<������<}1=OG>I�ٿ*�I�2վa��D���P������Ȑ�-ゾa�߽R����䚾r;�����ȝ���M�rj\�x���Vk��3�?�Y�?�����"���g��Փ~������R�>kJl�o����O�����ct����߾襾J_��xK��3h�q*g�b<,?�(�$,ӿ�L��,��@:?VB?zB�?~*��N�\a��rʽH5>��T����g6�ۿ��Ǿ�(?���>7���t%�=���>��=Lր<(�3>e_ �6jƾ~b:��?��9?g�?��;��ҿ��տ7d�;���?�l
@��A?ݰ(�#=�+�Y=�K�>�	?T�?>WP1��������ϊ�>%3�?�ӊ?�VR=7mW��5��te?��<��F����0��=�0�=�|=���;LK>�>��hA�D~ڽ�/5>Sh�>�3"����~^�'��</�^>aҽ�R��5Մ?,{\��f���/��T��U>��T?�*�>R:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=u6�����{���&V�~��=[��>b�>��,������O��I��V��=*����(gA��>���=����T_�L��=�bS>��V>��+ݾΰ��z<�mY>(��<_S�>,V)>|�g>T�:?Q�?$x�>�J�=���<r8��?�o���������0=H-��݆�!�k�Y�~���:�����:�J>�GH.��x)�ȏ>W3���ž�M$�Iz ��N?�&>����0b���9�{}��$m׾`z&>��Ǽ�<��e�&��j�2�?Ӫq?+$��ke|�_B��|�=1�`�??՝d�6+������S<��&>sKj����>0�<�7�v�P�ů|�i1?�,?�㻾a뎾��">�g�� 	�<Tu*?�?{6<R�>z%?�$�Ýн&�]>�7>I�>��>5�>W��~׽-�?QqS?l���R?��b�>3"��:g�]Mi=�>�Y2�|���NY>���<�ڍ����S3��T��<Q(W?r��>1�)����X�������==��x?՗?80�>xk?y�B?!�<}]����S�A�.�w=��W?�)i?��>є���о.�����5?��e?O�N>#Fh�S����.��Z�' ?W�n?�^?�ȝ�dt}�������g6?��v?s^�vs�����>�V�h=�>�[�>���>��9��k�>�>?�#��G������xY4�%Þ?��@���?2�;<	 �P��=�;?m\�>�O��>ƾ{������U�q=�"�>�����ev����R,�c�8?۠�?���>������[	>s����?��?}F���H~�,���i~��+�o@x=�a�;�E�<��d��A+��#����g�$�����.@l=r<S>�@�Ͻ>��> �=�3�m�/�����
p����#?���>������9����h����A�6o7�)Ҿ��>9�>n���6����{��W;�S���',�>����>�T��%���z��?�3<���>���>_��>�3��1۽�f��?�<��@;ο�������&�X?\Z�?�n�?�l?�Z:<(Bw�'�{�����G?�|s?OZ?�%�
J]�R�9�D�j?/���8`�K�4�ukE���T>�3?�K�>��-�\T}=��>�z�>�>^E/�X�ĿQ涿������?[��?���j��>ы�?u�+?�^��?��
���+�s&��$A?.[2>	@��_�!�c=��풾�
?�0?B��?�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�'�>��?��=�m�>�J�=����GQ.��Y#>�,�=V?�M�?Y�M?.D�>^��=��8��/��TF��=R��"���C��
�>��a?�zL?�bb>N긽)K2��!��Fͽ�i1�ȗ�X,@��,�߽߮�,5>6�=>R>��D���Ҿ��?�q���ؿVk��p'��34?��>]�?���Űt��L��4_?/{�>4��'���#��+���?%E�?l�?
�׾oW̼�>1��>�`�>]�Խ����sm����7>��B?��o=��-�o���>���?��@�Ӯ?r	i�&	?A �OQ��/b~������6�L��=.�7?a-�v�z>���>�=Emv������s�߷�>fB�?�z�?���>q�l?�o�d�B���1=�N�>��k?Ps??�l�O �'�B>@�?���P���IL��f?��
@"u@�^?b��ڿ�K��]1׾��㾘�r=��=�j >���Å=��+=
��<�2��i^���F>֩2>�T�>�� >��w>h9q>������I��0R��8�3�ݟ
����޾���t}�rm羥������E��I��J��`F�����t	9<��.>abM?��G?�?���>s*��@�=Ҷ���P�;�3��?��=�>��"?��P?��?�݌=����RV�8iu�������iU�>�A�>ܖ�>2�>0��>��;F&�>�� >���>[:>2���dR�P)�;;�>���>��?��>��w>���>9�ſ*Y��v�V�M��=MZ���?���<R�5��oo���G��q��4?�>u��O4��پ�ɹK?#����K9�u��<h�=E�&?�H:?��T>�ɾKkM�706=.��&%�j�ռ{}�����6B��?z�=�E?ޤf>2u>��3�_f8���P��q��3b|>66?"ض��-9�A�u��H�VUݾ�HM>�Ⱦ>�ZD�td������`ii��y{=]z:?�?O��\㰾Ʈu��L���@R>�Q\>%g=jS�=_M>.c��ƽ/H��).=-��=ݤ^>��?�!0>O�=�y�>����>�Y����>ɜ9>��1>��>?�)$?�	�����	 t�S,���y>�`�>b�~>���=�F�kz�=��>^b>.���U�q���*C���\>�T}��;G���"���=�Y�����=���=�p ��#6�U�.=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�c�>f{��Z������u�q�#=���>{8H?�T��$�O��	>��u
?Y?C]������ȿ#zv�g��>��?6��?��m�3A��@����>���?�fY?�ui>�c۾�\Z�ׇ�>��@?�	R?]�>e8���'�$�?�޶?���?וw>���?���?N&�>�2��w�?����m��}"߼�H�����>j����g_�>%��%���Y���M�Z��0��	ws=���>��:<���<��#�=�훾��+=�5�>嶠>^>�#�=���>	N?��>�K>��=j���2���L?4w�?�m���m��H�<[A�=�`��?*h4?�i�v�ξ��>Ŗ\?�׀?��Z?�ٔ>#�������󿿶����<ZK>���>F\�>L��j�K>?AԾ9�D��؊>,��>�ᨼ�پ,2��ε�����>�!?N��>�Q�=ə ?��#?�j>;*�>aE��9��*�E����>���>I?��~?f�?oԹ�Z3�����桿d�[�Z:N>�x?�U?ʕ>��������gE��@I�R����?�tg?RU彤?M2�?��??ŤA?�(f>W��Mؾ���;�>Q�!?��ʵA��E&��
��}?DQ?���>$*����ս#�ռ<��Ku��1?�'\?D&?����$a���¾��<�"���U��t�;�fD���>h�>a���yo�=>%߰=>m� G6�D�d<�g�= �>E�=�!7��W��0=,?ƿG�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?a��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�[�>���>+�l���K���ڙ���F��_�Žv!=���?���>���>�M'?�pQ>ع>,Y��|�#���@�:��hX0���6���"�T�4�BE1��+����+���=\Hվ�e��@`> X�uc�>qc?d�=��;=Dw ?��-�1�>��2> �q�h_>���>4�>�H>��<���AKR?m����'�Z��|����8B?md?�-�>gFi�e�������z?��?�t�?Qv>�th��&+��l?v3�>`���l
?��9=nh��<�<�X�����6E�������>{/׽=:��M�?�f��m
?1?�5���{̾S׽�������=���?g*?6K&�
�V�CSr�XwZ�K�S���=�N�d�T����T%���r�ќ��Y���{����'�{C&=�'?7��?tm����b���0j�� A�y_>��>sF�>$/�>��:>��(�-���b���%������(�>��s?�M�>Z0!?4E?��P?��#?���>$��q�m����>&�Խ��?#�>��d?J2b?*3&?b}?h1&?�Q{>A����G���.��x�>&?݇3?��?�6 ?����(�uy+��M.=Gf����<��_=��<Û޽%h����;Hp>�X?�����8�����k>�7?c��>���>d��,.����<��>��
?K�>b����wr�_^�Z�>��?�����=��)>���=w��^.Һ X�=�����=
��iu;�9�<q}�=�ڔ=SCu���}��L�:��;n|�< u�>6�?���>�C�>�@��0� �b���e�=�Y>@S>~>�Eپ�}���$��u�g��]y>�w�?�z�?ʻf=��=��=}���U�����G������<�?@J#?'XT?`��?|�=?^j#?˵>+�hM���^�������?��+?��>���3�R+��F��8 ?H�8?ML���<��MA�pվ~�G>Q�C��@i�; ��կ���I��>��� (]���?β�?Ž?��t�����ϥ�����d�#?<9?"�?��>����k��Y�>�Ã�>`��>]w�?@��>D�'?�^x?JS?��A�l-����P���p�=�`<KM?8^�?�ۈ?�&�?���>Bu>
R)�k2�T�%�@	R�6��� t�0���_>Y��>��>��>�t.>~�0��'1��L��bv=�7`>�H�>,�>�r?��>���<C�G?ɫ�>k��xf�������l?��bu?���?^+?�e=U>��E�/���@3�>�f�?�?�)*?�kT�1�=aռ?�����q��9�>��>� �>��=U�D=��> �>�e�>����[��G8� �N�|?FBF?���=n}ƿ������.�����=|�k�B�
�1,�=�|�)B>����Ϡ���ҾzV�lf������!ｾ�9���=ݯ?�w)>Ff>���=�K>>?>�;�=wa�>͘�=6>=b��%u)>�o�=�H���<���=��=�sY=Q("� g˾��}?�-I?��+?�C?IJy>�%>��4�ɓ�>����e5?��U> �Q�ac��T�;�e���� ����ؾ�`׾��c��ڟ�!>I�"�>kL3>���=,�<� �=�s=/܏=\P6�Bu=�H�=�P�=^�=���=��>�(>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�G8>��>�zR��R1��k]�tQb�Nk[�Rm!?��:��D̾Z`�>��=ջ޾D�ž��/=J7>�c=���
h\�T�=&�y���;=&�k=��>�yD>�ź=7����=�L=�Z�=E�O>`2��T�8���*��V1=�;�=��c>C�&>��>Ci?��,?��b?~�>�/���¾�!���-r>��=|�>"-z=�g>#e�>�=?@�E?]QG?��>�<P="U�>ҥ�>@N.��~k��z&��Z�=W��?��{?Ӎ�>ZX}<�9�D���1G��I{��e?d�,?�4?o��>*�k�ٿ+s/�s�5����u�C�<�<����Z�<>%<�u���m�0����S>�^�>D�>*�b>O�@>��>�1�>>��^=��=	3b=�Z*�$����P=�(��}�<ei����ý�u��q%���v�������<;`#���u�<L��=�P�>�<>���>���=d,��<4>쓾��M�,m�=u�����?��=c��{���/��0@��x:>}�S>�Ws��C��e?�aT>r�8>ӓ�?Z3v?"*>RL�S�;�s���X� P��m�=��>1�� 9�F?^��J�DӾ\�>-�>1��>|cB>οA�CE��aM>�'ʾm�u�5G�>D�����<=-��q������E��_�h�����B�f?c���w�J>�ZU?�>? e�?m��>�K<����>�>�#�t�L>[�ƾ�����>ޱA?PC?��?������@���̾�W�����>�wJ�n�O�����0����s���L�>�"��(�оt3��G��Wݏ��zB�o~q��>��O?c׮?-Kb��K��z,O�l���e���[?*�g?���>K?��?����Ӯ�򢀾<b�='�n?W��?�&�?H*
>�r�=�Ц����>��?�.�?�Փ?�$k?',��2�>�n���P>K�����>hP>Y��=PZ>x�?��?�!?���
b�����]���o���L��;n>���>z-Y>|�w>}�=L�=��=23>�ά>f�>��Q>�6�>+�>ᴾ��ܾV�?!�=j�>rF,?�o�>�9w��������+a�I%��`��Tn$�=(��Px��+@8��; ��=w��>Sֿߤ�?uZ�>1C�J��>������<��>s"?�dD��1�>��?�G�<�?+z�>!X�=��>�M>��Ӿ �><���!�=8C�X�R���Ѿz0z>a_���&����L����I������B��i�����'=����<3�?������k���)�Σ��c�?	�>T�5?D���kӈ�v�>���>b�>�����m���Ѝ�����?���?�;c>��>>�W?(�?A�1�^3��uZ��u�M(A��e�@�`�{፿����֗
�0���_?��x?�xA?8Q�<o:z>O��?��%�Jӏ��)�>�/�';��?<=�+�>�)��E�`��Ӿp�þT8��HF>��o?$%�?cY?�TV�/Q`��+(>=w9?�7?%�w?�d>??�*?Ö꽗?CI>_�?� ?��;?�:?�O?��D>ޟ>Z�V<��W�����?���8��|ٽI/��{�=`*>Կ�1��1=�<G�-��<c��	�;���<*X.=�� <�ު=%�>���>"]?��>dӆ>>�6?`6���8�4����9/?�u5=G��y������4��
�>��j?���?8Z?;�`>�B���A���>w�>*�'>�]> S�>����2G�g��=ӑ>�5>�Ȩ=�M�������	��G��Y��<^�!>���>�%|>�썽	�'>����O,z���d>��Q�:ƺ���S���G���1��sv�_]�>��K?v�?ꠙ=*W�@���Ef��-)?{Z<?zLM?J�?��=~�۾D�9���J�G4��>�r�<&��ڿ��� ����:�*1�:��s><(���x����Y>��
�	�w|o��G�^��A�k=�{�mTD=v��?־y�~��'�=Bc
>DZ��$p�w���]���nJ?��=>����Z�{���l>�>��>.X�<��V�>����I�{=]^�>J>Θ�����H�r<�Oԝ>�B?��k?@��?*����0�����i}�����>E?��>��?�5x>��^>�mH��0ھl�Z�lX���>Ok�>$)���4��J���ɾM8��->�e?gKJ>���>�e?F?�#^?��C?�"?��Y>i��u�}�o2?�-�?ҝ_>��<G�R��b.���<��S�>4�?�c��M̼>�C?��)?�?v��?�)?��y>�Mž=@)�NX�>P�>�d<�Y,���Ԯ>��?�c�=��k?��?.2��n��q���'��H <cƫ=��?ݾ-?bC?v�?��%?c�������>�Wi?oڋ?>�?Y�=��?��J��5?S��>8� �C�??�>��l?0�d?6K�?���>��-=u&�&N�#������/ ���p�=��=\�0�7�֎���C�=K`"���7��<D�=X�T��b��.��>��s>^땾��0>��ľ!���A>���L*����:��η=&�>� ?�.�>f�#�q�=���>A�> ���(?	�?�?�U�:'�b��ھ��K�D�>�8B?���=�l�Eh��:�u��jj=f�m?=k^?�OW�s���J�b?�]?h��=��þ��b�҉�R�O?>�
?�G���>��~?n�q?U��>��e�(:n�%���Cb�/�j� Ѷ=Lr�>OX�@�d��?�>n�7?�N�>Z�b>�%�=gu۾�w��q��f?|�?�?���?+*>~�n�S4࿓r���T����]?���>6��#�"?���g�Ͼ�#���x��0�n`����� Ε��*���]$�Wr��c:׽���=��?S!s?:�q?�_?ܴ �@
d��H^����QV�e;�f���E�� E�كC��n�<���;��H����jA=�z��TJ���?�1.?'�K��S�>E�n�~���yξՎ�>����`�?��k>�0�p��=k=P�?��z������@?^�>z}�>��??`�J�KD<���2�Z&5������.>�M�>zw�>���>�&�bI�����@������0e��>�>��m?�U?��r?e���?��a�u����ͽ�!�Xk>���:�>���V$�\{�E^���]���5�D�h�w���1�='/_?xQ>η>�_�?�k?4O?�&�ɽ�۽7�0�U���f>�J?���>S�>
7��;%�Ϸ�>��l?-��>��>����\!���{�V�ʽ �>��>���>_�o>�,�	\��h�������9�AX�="�h?�����`���>�R?◁:� F<=��>��v�d�!����c�'�C�>�z?E��=��;>^wž	 �l�{�[3����)?��?
l����&����>I�#?+��>��> Ƅ?�v�>|���P�<�?�b?��I?}�A?��>�w�=�'���)Ͻʮ)��C!=�L�>�YU>Ӎt=T��=�(�i�]���$��8=C�=:�ؼ6��[�;����g<�n7=@55>aEѿOU����c� �@AоH⾡��H<�������F龜��k�۸H�я��!��i/�A[��:*�����?hj�?Y��\q�ˆ���҂��k���Ƴ>�u�3f��-f�8w��¾$�d���o�9�P�M�u�~�`��4,?�m�-(ǿ���k���i?"�&?Z�?�-�O�/��A�]~=r큽V�Ͻp�ھ�X����ؿsd��L\A?K�>`�ݾ ء<2?�O >���;�$w>����u��E!���?ʊ$?��>�pb��=տ̿�=�,�?P�	@\B?�(�*���c^=���>�
?V3G>-��������%�>�,�?=��?�F=��V�P�ܼ�f?mm<L~F�򗻆N�=���=}�
=M���G>L��>���c�D�?�۽}?;>�Ç>t?�A�^�{�<��]>�!ͽ�j��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=v6�����{���&V�}��=[��>c�>,������O��I��U��=]���:ȿ��h���R�Ҷ?�B>%F&���c<���>a?P>��@�W�ɾ��c>VY�<E�>���>k!�>���>:$�>?d_?�t8?�A�>;Aq�����9�樾��=7P	�����h����������
�e��w���( ���$��X	��S3��B�K;�����S_5�� >���@���2?Աx>��ɾF�a�y���8��N���u�r�ν`���*M�����?�S?�~f�r�P� +�ŭ�<65(�X�O?�5^��}�?���2�Q>y�B��'u�Q�>Y�=S��#L�$�3��K3?��?�ž�߆��y<>ߓʽ-ɋ=DU)?:|�>a~;��>])?ةS��	�j�[>�L>b��>:A�>�>fA��>�ؽ�"?dO?��1���4�>7���m�t��=��=@�g��j���1�>�=m͊�b?��΁�|�H=�)W?Θ�>s�)����X�����k�==y�x?[�?�(�>;~k?��B?�<f����S���K�w=P�W?�'i?>�>�����о�~����5?қe?�N>Qch�:�龯�.��T��?S�n?c?�1��\s}�S��4���o6?I&{?�@Q��s������׽��>�?���>W�,�^�>ٸQ?]`�<���Y���z�)�U��?���?���?��;aB��m=���>���>J��� ߾M��B�����==,q?%q��������JF�4�2?.�n?@��>4�S��{׾a�=韾�R�?��?�������z���m����?[�=��<����(��=R='�&��&�׾|+����>w=�Ut>zD@���=eN�>k�v��ܿ����Q��vҾ,�ۋ?�]�>�I���OK����������q��k����gL�>��>P��������{�op;� 0����>����>��S�&�� ����5<��>ϭ�>��>m;���꽾�ę?i_���?ο⪞�g����X?�g�?�n�?Go?Hg9<��v���{�޼��,G?N�s?�Z?ŏ%�+B]���7�<j?�0��<�_�<�3��?G�f�J>$�2?S��>��/��|Y=�>��>kP>�70�`�Ŀȓ����:��?��?�3���><�?O,?����b���¬��	/������A??>>���g�!�`=��ё�Ɓ	?ө0?��x��]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>+�?�~�=�W�>�M�=}̰��y*�Nk#>�0�=�@���?]�M?s�>R��=eo9��/�OSF�e<R���ʶC���>��a?/pL?}�a>DU��S�1��!��mͽH�0�J�=d@���,���߽KX5>�>>�>�D�4�Ҿ��?Mp�9�ؿ j��p'��54?0��>�?����t�����;_?Oz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>;�>�I�>A�Խ����]�����7>1�B?X��D��u�o�x�>���?
�@�ծ?ii��	?���P��Da~����V7����=��7?�0���z>���>��=�nv�ػ��N�s�й�>�B�?�{�? ��>�l?��o�V�B�(�1="M�>��k?�s?�Ho���_�B>��?������L��f?�
@yu@a�^?"�|ٿ�����8���渾��'>��>�ů=^�?�e��=������\��-&�q��>$ϛ>a(G>-�>p�Q>�d<>���v� �U��6���S�!���	����#C�#��0`�F�-�M�����o&��ӕ�ti��������o=u��=:V?a�R?q?�
�>����O�>d�����<k3��q�=���>�3?��J?W	)?K��=l���ںc��������R���M��>W>��> ��>R��>E�;��:>�/I>��>��=	9=B��V�=$�U>��>���>\W�>	-d>��>�=���N��M�v��	�o�t�)�?���DN�p ��";Y��`ξ��(�ׅB?`�J>Q���(տ!䫿M�L?����<��tF��C>��?�_?���>������}>�F^��\h�,�K>�}��-���<p��r�>��?c�f>�u>��3��b8���P��s���j|>�16?bⶾ�O9��u�/�H�vhݾ�IM>b��>��D��k����;��oi��{=�t:?	�?�^���㰾�u�ED���ER>R\>��=wR�=�SM>�c���ƽ�H��R.=���=�^>�~?��>�@�=AU�>��N�0y�><9>$>!QD?T�!?T�j�iY'��#������Jt>�>�x�>�>^�?�5y�=ٓ�>={r>@���T������H�TNE>�_V�%�p�ײ_��J�=��J>���=��=F��=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾;`Z����>һ@?�R?�>�9��'���?�޶?֯�?%e;>��?|G�?�O�>�����_�n�ȿ�n���Pr���N=�a>R�6=B�h��X��)��<���g,Z���)�]��<z�=VG�>꽫ؾD��=O��;󨽾K�<��>m+�>'��=Z��=�}?t ?Z�n>�Yk��'���E��z����K?&��?]����m�6'�<!��=^�^�p?�U4?u�V���Ͼ���>$�\?��?��Z?�_�>����1��m翿�d���ۓ<[�K>x��>�W�>9)��WeL>4wԾ�D�Y{�>�ї>�ꧼTfھ�E���e���K�>&�!?�B�>���=ٙ ?��#?��j>�(�>BaE��9��Z�E����>Ԣ�>�H?�~?��?�Թ��Z3�����桿��[�h;N>��x?V?vʕ>a���񃝿�kE�$BI�G���\��?�tg?mS�0?;2�?�??b�A?w)f>և�&ؾj�����>۽!?|�ЭA�'A&�g��~?�Q?���>i���6ֽ�~Լ������ ?}\?�-&?h��.a���¾���<�j$�ZrU����;��H��>��>�݈�Ci�=ʆ>�D�=�qm��%6���c<�=���>���=�7�RB��M=,?-�G��ۃ���=	�r��wD���>�IL>���V�^?]j=�p�{�����x���U�� �?ܠ�?ik�?G���h��$=?�?3	?�!�>�K���}޾��4Pw��|x��w���>���>N�l��!���ؙ��jF����Ž8B�o��>?��>�{�>DQ�>�X>uϵ>�g���pu)��`����G�E�C����S�o/-��Q�{�k�;�=6�Ǿ�1�òr>""����>��?}�n>��u>k��>D�c���j>�E>o
�>�R�>M��=�g>6݈>+�<|R��KR?�����'�`�辤���e3B?�qd?@1�>�i�9��������?���?Js�?O<v>�~h��,+�nn?�>�>;��<q
?�S:=�9��7�< V��=���3��N����>�C׽� :��M��nf�j
?�/?�����̾�;׽�s��qY�=ù�?\F)?�)�L�S�4�p���Y���S�f�&�=�d������$���p��ޏ�Hv�����-�)��=/X)?���?� �]��媬��i��A�l[>;Q�>1�>}V�>�hK>�>
�L	-��t^���'�?���5Y�>� x?���>�~V?��=?a}??,�D?`��>��>�x��ő?C��Ǵ�>[6�>46(?��@?n�2?�?'|5?���>����^��Ǿڣ�>��?+�?):?L?����8½�琽�r�;�;��&n�4R>�we����8�J��;1>I�y>��?�E���1��z��4f>	|6?a�>���>��������p
=I��>�>���>��
��Mr��Z�B.�>��?�I��=ʪ!>S�=*���]l�:��=�b��}�=�-�<N�н�<B�=�Jl=��h;7܄<)-E<>d�<K�q<hu�>��?ꒊ>�C�>�?���� �ʵ��f�=hY>GS>m>�Dپ~���$��.�g��^y>�w�?�z�?�f=��=q��=�|��?U���������+��<��?J#?@XT?7��?��=?!j#?ܶ>�*�EM���^��s��خ?�(+?��>t���վ�ۮ��6:� ?�e?�x�򪆾I] ��ʡ�qa�5�<��N��荿�ȶ�E ,�m)>.G��?�����?k��?{p��I�<�u����2������8?E�?'��>�>*G)�R�i�-)%�	�>v��>ϿX?�a�><Za?�,~?7cI?R�>��@��篿Z"��4JW=�w]>��/?�=a?�3�?�?k?�b�>�oF=��I�`@Ѿ�%9��$� ������>�J�>��>��?��>p;>��ؽ��<����"��=40)>���>ι�>���>�2>�=J�?FH?:r�>�*�����aP��XO��^�;���u?�h�?d*?t"=q����D�5������>0b�?/ޫ?Dz*?�}R��^�=��Ҽ�ַ���s��Ÿ>؝�>�>,��=R�M=�%>��>C��>�u����i�8���M�!�?ՇF?�6�=*ſ��p��r��!���\�<�g���ra���ixS�Y��=�V��GS��M���V��������_Ҵ��U����s�:w�><у=cn�=���=a��<A������<��>=��<��<=X�^<@1'��Q������.e;#�:<ܰG=����˾�%y?42F?�n)?ʛ@?�.�>�>N�!�b��>���~�?ҍW>�������V�Ϭ��얾��׾�Ѿlc�,����>�~W���>0�,>���=�<�=/,�=�=Q7��m3=s�=���=�/�=u��=�c>mj>9w?����$���"#Q�,�潬�:?�U�>���=�wƾ+@?�%?>�#�����4a��#?��?�M�?g�?XWi��T�>;���h����r�=5+��=�1>���=+�2�P��>�K>��YQ��:Q��55�?\�@�??�㋿Z�ϿΏ/>�6>��>�#R���0�\�?`�fHX�E!?��:��;ц>X3�=�	�ž=.4>"�[=�~�4|[�˷�=�h|���:=vpj=Z�>Y3B>�C�=�����=^�^=�5�=N>�Ɗ���?���"� b;=�T�=R	c>?�%>r�>8?'�2?rHh?x��>����
�Ǿd������>p�>���>�ȶ=_&]>q��>Ƶ??#�F?�H?�z�>I�-=�ݻ>,�>A�)��w�� ܾ镈�!���6�?��?aZ�>y(9<q
�_����>�!ߗ�p@?�Z1?��?���>$����࿭�&�((�2��f�=�{�<��O���������T���u��+�=��>1)�>\��>v��>Rce>�/�>�>6��=�������<���=%ı����Ɓ�=��>%6�=��A���½��=yt� a���d=�k�=��<���=>��=^Q�>YX>jd�>�7�=�峾GZ/>���\�L�҈�=|Ȧ�3B�ۭd��~�>/��7��,@>�V>�9��!��ۜ?FZ>��?>��?=xu?KR >Le�aaԾF��ff�.oT��n�=d�>��<���:���_�|�M��ҾP8�>�6d>�k�>�	D>ʾE�2B�(<�=�3Ծ(S�	�>�H��̮�IΓ��Y~��[��j����{�ۺ���J?vU��As8=�I�?�H?+�?]��>NνK����>=A]�}�=�� ��,��k�$=�K!?��8?���>�A�xN��H̾_!��Oܷ>4I�.�O�U���`�0�]5�"˷�3��>�몾��о�#3�Ze��j���_�B��Vr�m�>T�O?F�?2gb��S���IO�����D���s?�ug?��>CT?�7?Q���]������ȸ=��n?��?[:�?�>y)�=�]����>�u?�ٔ?@w�? @s?�61�t�>�<輗p7>���N��=��>^sN=U��=��	?	Q
?�L?h��f�Ӏ��k��I^l��LI<ީ�=,C�>e�}>[�>��>	��=%Os=��8>�j�>W�>��b>���>G�>�\�����pE? .:>��=��?M{�>?ͷ�/S���=�ʓ=�����8�]�������������x+=�]>��>*ο�M�?3A�>���ey�>ũ��Ҳ����z=ak�>ӎ��M]>� ?❽��?�5�>Q�>˱�>�/�>FFӾa>#��e!��,C��R�$�Ѿz>!���9
&����x���BI��n��5g�jj�n.��l<=��Ľ<H�?J�����k���)�W����?�[�>�6?�ڌ����Y�>D��>�Ǎ>�J��t���ȍ�7hᾼ�?9��?�;c>��>I�W?�?ْ1�53�vZ�+�u�n(A�,e�U�`��፿�����
����-�_?�x?1yA?�R�<,:z>Q��?��%�Yӏ��)�>�/�&';��?<=s+�>*��-�`���Ӿ��þ�7��HF>��o?<%�?wY??TV���e�n�)>~:?�1?�[s?�2?z;?Ie��@%?.>�o?�K?V!4?=F/?�s
?�3>�+�=���9��7=���(��wϽɽj����6=;Uz=	�]:�|<��=煗<�t��n�:@�����<�;=ts�=���=�Ϫ>l_?̺�>Bq�> 47?��
��6��;��z�1?,=��s����ԟ���㾶�>J�j?zr�?�\?_�m>�D�
�A��H>���>�0&>Oza>K�>����pB��xj=g�>d>yƑ=�i�����I��(N��?�'=r%%>��>�.|>����f�'>�{���3z�=�d>��Q��̺���S���G�@�1��zv�8V�>�K?w�?W��=�^�_1���Gf�d.)?0^<?aPM?P�?1�=0�۾��9�>�J�!8���>�:�<��������"��^�:����:ټs>�1��cf���VK>1\�/Z�B� %V�ߧо��>Z����jj>��������8p�&�&>��a>A;�����鍿m[���j;?�_�=�þKJ�ǣ� �R>6��>Eh�>F׺�Ę;� F�X���'��=z?�>Rw>l�=L��H�F��J��}�>#�D?�~a?a��?]�X�q�t�JjG�����G��w�7��_?{�>u�?3�0>�|h=K5��O�
�'�e�@�I�}��>�>��r=K��1�����;� ���i>cX?�>�e?=�S?�?U�`?�*?A?o��>p��-)����$?�Ƀ?0�^>���DU�(H.��#8����>�#?���\q�>�&?�'6?&n#?_$Q?#?�y$>�%���8�~��>*��>�r?��O��R�>"�`?*��>Rb??O?O�$>$(��֯���e��R�=2>u5?yh?fp$?Pc�>���>���S��=�^�>�
?��s?�ߌ?��>M?>�����Q?>3?>�&����%?��#?�V?�T?�d?jX�>P��������O� �Ǩ\=3W�<��;�T<�<eFv<'���r<`�}=p��[���!\�즄<�?Q=v���!4�>��s>$��}�0>��ľ�1����@>�8����� A��Э:��2�=)*�>+�?�x�>�#�֒=��>=�>(���'?[�?o�?'�;X�b���ھlQK��9�>7B?���=<�l�#Q����u���f=!�m?�^?UOW����L�b?��]?5h��=�	�þ��b����Z�O??�
?G�G���>��~?c�q?M��>�e�):n�(��Db��j�Ѷ=Xr�>KX�M�d��?�>l�7?�N�>*�b>:%�=gu۾�w��q��j?��?�?���?+*>~�n�V4�g�Ѿ�s��}(X?���>P�ʾ2}?Ώ�� �ʾ�Ub��@�d	�5�Ծ�2�{�̾��ľ�s8�{N���˽3�*>s�?u�Z?Y�x?qk?6о��]��l�|7����n��þ�1���N���"��=J���c�U&���" ƾ�u=�wx�e�C�`س?ca(?~d=���>[��D���ľk�H>\���|����=C몽��=�TR=E�[��)�[K��� ?F�>HB�>R??�6Y��=��2�7�7�9����oK>N��>7�>e��>�G���/�4��E�̾�%��2 ½�j�>��p?ǒN?Ufa?T��$7>�zޅ�gBJ�XZ�=�ݭ���>�f)>i�>�t"��>g�:N�C�4�N�|�s.��
��������<��3?m��>�Tq>蟗?�?y�������2�~��"����=�q?4Cw?L� ?Y�J>^���3|�s��>R�l?N��>��>c����Z!���{��ʽ�'�>�ޭ>���>a�o>�,��#\�k��F����9�gl�=Y�h?������`���>�R?젇:��G<�|�>��v�<�!�S����'�x�>f|?r��=՝;>~ž?$�æ{��7��%)?af?�N��8�)��z>�|!?1��>�C�>�L�?��>^K��>��:�?{�^?u�J?��A?�x�>#]7=���ZȽ��&�l�%=+�>��Z>�Sw=�]�=�����Z�uy ���A=\ʴ=,��&c��b <z综a[Z<i�	=�G4>M׿b�D��Nܾt�����������)c�5|��	ܚ��1��M�����z��R�5��uo;��U��^��=�q�ch�?N��?C���Lb���9����q�M�'ˤ>Q�n��6��U������jљ���)����4 �z�B�"�c��^f�	�0?T�׽:ڿn������Y?�� ?���?9�0�����S��^1=��u>������������o�,3b?�1�>�z
���>�=0?C?>m�#�N�>��¼2�վ����w�?|y?�&?-����VݿpϿy���W�?0@�wA?f�(�!��2cW=��>�	?g@>�,1��T��	��Z��>09�?V�?�O=ưW� 5	��ye?�<��F��W㻨��=*x�=�=d���{J>|1�>����mA�$*ܽh�4>>�J"����3^����<ل]>Iֽ�锽5Մ?+{\��f���/��T��
U>��T?�*�>P:�=��,?T7H�^}Ͽ�\��*a?�0�?���?(�(?,ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=6Ἠ���w���&V�q��=Z��>]�>��,�ߋ���O��I��`��=m���������!���<���=z_����!��H�in����>:�����Խ !3�e��=u�M>�Y�>�\�>��>�H>�{?qyw?]u�>�T�=��޽�U�̈��j(��!ý�A>��C��f]={9m����1�4����T�����X.���=>��S�h�����h�C�*��
�5?F�=M�]�@��,s��yǾ�����r<�J��B���i)���`�qא?.xU?i���� v���=�X��>��;�?ٮR�#4,�-�׾PAн��� �~�3 %>W/"=�n޾�G�`WR�Pv0?�@?Ƚ���y
)>9���=��+?]� ?��J<���>ܴ$?�J-�%	ܽ'�]>v�5>bL�>�[�>�v
>\��8�߽`?�jT?2� ��蛾F%�>ɇ���w{�FW=��
>�4�M��(\>���<�K��z�[�^0��2��<�W?T��>��)�7�lH��e��==�x?��?|g�>�qk?C?V:�<-P��+�S�:���w=g�W?� i?`�>Z@���о\x��>�5?ՙe?�O>�h�u��q�.��R�_?�n?�g?����p}�������Hl6?��v?�r^�Ys������V�w=�>O\�>���>��9��k�>$�>?#��G��Ѻ���X4�0Þ?~�@���?��;<; �Y��=�;?H\�>G�O�<>ƾz������G�q=�"�>|���cev����DR,�@�8?���?���>����~���10>`ѹ���?~��?�����>Z ���v�ru��4?>N�b��捾j�4>��&�kQ�����W�,�۾I.6=�>�@ކ`�!��>�6�=�Ŀ)�ۿp����d���1��j? ��>[�/�S�"��1Z��z��H��a����`>�>Z�> ����/���{���;��Ԟ�a�>Ɔ�_b�>U.T���1�����:<�6�>�$�>?N�>χ���ؽ�f��?c���pο-v������X?�<�?;<�?W�?��<y}w�ͥ}�o���kF?ƾr?"�Y?~E)��y^�ؾ9��k?����a5e��4���k���.>!m?�.?	nX�/I�=?�Q=�/%?��@>4Ja�.ȿ`�ƿ��0�W��?�d�?\1辁��>���?W�M?��'���������8H��Yټ�)?�#�>�橾FxP�ٙ.���b����>1X?.��F��]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>`H_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?�#�>��?|��=�e�>���=R���K�-�ig#>�?�=m?��?��M?KP�>�b�=(�8��/��XF�~FR��&���C���>��a?ĂL?�Mb>����"2�	!�uvͽ\1���輰J@���,��߽�.5>t�=>(!>4�D��Ӿ��?;p�5�ؿ�i���p'��54?!��>-�?3��m�t�F���;_?gz�>7�,���%��IC�X��?�G�?/�?��׾�L̼^> �>fI�>p�Խ;���b�����7>7�B?$��D��p�o�j�>���?	�@�ծ?Zi��	?���P��Va~����7�e��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?\Qo���i�B>��?"������L��f?�
@u@a�^?*��п����Z@������Fٳ=ɬ=m9>)G�Tٕ=���<GPe=s���:�=^.�>��>	Mq>��>�5q>��3>�"����$��T��^���5�d �?��99�F�ee��&4��s����Ӿ�μ,s��KC���Bt��᡽|>����>ּa?x�[? 6v?{-?�^�������v���Ӑ>��b�O=��7>\�S?v^G?���>���=}����R�@��������B�����>��>��?b;�>]�[>��>��'>�H>Q"�>�HD>�C��*<�{�=�	>f.�>�?R¡>��O>w3�>öĿ\¿��v��۹��2�����?h1����1�/p���U�%���YV��J'?���=�0����ؿ�*���[?�����}8�����:>'�N?��'?W�u>7Ⱦ��x=��V������7=��U��H���ao�ZCd=��2?
f>��t>Q�3�q8��qP�Aϰ�G|>3Q6?�����7��u���H�?ݾ�M>���>��C��m�떿��~�e&i�{b}=n%:?>v?C����c��w/u����v�Q>P�Z>R=.�=t%M>u�g��.ɽEG�o.=D8�=A*^>5�?�Y>��=���>�v��2�=���>�=>Ź>�=9?�M*?>�����½�l��J��X�>[��>��>�s>�N�ݙ�=���>o�O>V�4���Y��,�(;�L�X>�\z�f�`��|���p=u���"
>���=o���+�J=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾQh�>yx��Z�������u���#=Q��>�8H?�V����O�h>��v
?�?�^�੤���ȿ6|v����>X�?���?h�m��A���@����>9��?�gY?qoi>�g۾<`Z����>ӻ@?�R?�>�9���'���?�޶?֯�?��R>j$�?|�k?�,�>�%>Jq,��(ʿLQ�����>�)��"A�UJ�9�1�ҙF�Nd��{�����>��g�=ގ��s_<���>N�Y��ž�	��.ĽXh����xF�>�@.=��>i��>rx�>��>)�o>��@>m�A�V��p��~�K?���?���#n�b�<�5�=z�^��?�O4?��\���ϾoŨ>,�\?���?��Z?Eb�>���o<��N迿�}��\�<�K>�B�>�e�>�D��*K>d�Ծ3%D��h�>�֗>Z���DھS"��cE���8�>f!?X��>�ɮ=Й ?��#?ؖj>�(�>aE��9��l�E�<��>Ǣ�>�H?��~?��?LԹ��Z3�����桿��[��:N>��x?�U?�ʕ>P��������`E�gAI�:���A��?�tg?tT�A?@2�?��??{�A?V)f>����ؾ���f�>h�!?zt��P@�'�$�$��!?]�?��>r����ѽU,�����^���?��[?��&?[��t%_�|����}�<n��k��D�:;�����>��>�܉���=�D>n��=h3d��Q5�9�K<� �=7l�>���=��3�oƑ�%=,?��G�5ۃ��=��r�xD���>�IL>�����^?m=���{�a���x��$	U�� �?��?Jk�?R
����h�u$=? �?{	?r"�>�J��(~޾&�ྯQw�m|x��w��>;��>�l���H���ș���F���Ž[��u�>�l�>�
?��>���>��>R�����F�6�����O�m�*��&�rL2�2r��������j�l=7�־��Y��vt>�؞�Θ�>���>^�S>)�>�(?(����x>W;>j�>�(�>�uT>W��>�>"�C�z�'��KR?����Ѿ'����d���\3B?�qd?�0�>�i�B���@��t�?2��?:s�?�<v>�~h�s,+�`n?_>�>���q
?�N:=KE�=8�<�U�� ���4�������>�E׽� :�EM��mf��j
?�/?3��o�̾E:׽�J���[s=n0�?�h)?��(���Q��,p�>�X��+R�$��tom�����4#�h�p�� ��ߎ������D`)��� =�(?`ۉ?������ ���$�i��@��b>�Z�>�V�>�R�>N>"

��u/�^A]�'('��[�����>Ynx?���>!I?6xM?��E?��(?��>r��>
1����>G4�x8�>R�>?B$C?��:?�2%?I�)?�f�>�ü9?��z���Ó>3l?�?�J�>��#?���D�L9$���>�՗�#g��3�I>�<@8�2���Xd8>�ki>LW?�����8�m�����j>�~7?Ԝ�>���>���#(��z��<��>�
?zT�>����a_r��X��\�>��?
�/u=V�)>���=X�����ʺ/Z�=;���
�=+ȁ�Y6;�n7#<qk�=Uؔ=T�i�BѸ!f�:�;Mɮ<�t�>/�?���>�C�>�@��'� �\���e�=�Y>�S>R>�Eپ�}���$��t�g��]y>�w�?�z�?�f=��=(��=�|��yU�����^���O��<�?EJ#?=XT?Y��?r�=?pj#?��>+�]M���^�������?�C/?*|�>-N���־���W!�
�	?5?Fl�����A+�mv��ɲ9�R U=��:�����@��Y%9�ܴ�=]S��ܽ�<�?r��? �н]�K�<����첾��:?�]�>]�>�D�>p�+�v+g�j�$�wp>�y?�(X?餻>�kY?��?�g?��>:T��5��c���I�i>p>3�,??Ü?�e?��>,�->�r�w��l�&�ׇ�� �<*����iȆ�牦>�k$? �g>��'�hΝ<����Ƈ�|>�1�>��?��>�\�>�� >�3>*�G?�_�>���yu�r��o��4�s�s?v��?�)?�xC=B���'F�����g��>���?I��?ܚ-?��L���=<�ؼY4����n��V�>B��>C��>C��=*g=4>��>K��>;������5�Q��;?�pF?��=���c�b�وѾ�ӥ=nY־�~���G�;���/�>䕌��@�<O���&�W�N�|=��������~Ss��?r]%>�!�=��=��=��I�Su >�>�HS=�����Ҽ~����y��=�~�<ŽPf��4}]�4=�^˾8�}?�:I?��+?��C?V4y>>ޗ6��Ԗ>z����?�V>c�N��t����;�ר�+����ؾ[�׾��c�ժ���E>ZJ�I�>�63>~��=��<P��=
�s=�"�=�
J�rk=*��=l|�=���=���=>�S>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?��>>�2������yb��-?���?�T�??�??ti��d�>M���㎽�q�=H����=2>s��=u�2�U��>��J>���K��B����4�?��@��??�ዿТϿ7a/>yI7>�>jR��[1�r�\��3c���V�);!?��:��ɾ��>{L�=S߾��ľ��@=+�8>vh=s� T[����=�\w�.)5=w�g=W�>��D>�L�=٨���=T|?=y[�=�K>�x��d=��%�q�7=��=�Gd>�%>'��>�?o7:?�^?8C�>tp\��ž4s���ۆ>s]�=}E�>�)�=�Ud>��>��8?�I?'�H?б�>�M�=� �>G��> x*��l�W޾>���f��=E#�?}�w?4�>i�=yjd��.��j/����
?G\,?�?�Ѵ>���ص�nYU���:���<��ݻ"��=��=
Ǌ��HX����L�z��5g���>8A!?���>Ą�>ͣ�>���>h��>�c�=���=�YǽI�A=���;��"�>�J�;�N>ֽ��)�C=|$T= >�y���=�>�=o���T�KH�=3��>��> �>���=B5����->ly��тL�M�=�ꧾ�B�Y�c��J~�A/�d8��eA>t�V>Ą��*���d?t�Y>��=>�~�?�,u?��>p���2Ծ�U���d���Q�$�=
�
>��<�);��_���M�C6Ӿ'��>��>�Rc>K�>�,o�_|<�����¼���Q�&Q>����O+=#ܢ��N��U����H���k�.�J�X?Ԉ��>�,c?��U?��?f�?�j=	&-��-�>S���	���,�|���a��>�&*?CAA?]�?��Ҿ4T��G̾e��Dٷ>@I�@�O�������0�jg��Ʒ����>9����о�#3�Gf�������B�MGr���>��O?��?>@b��V���SO����D+��]o?}yg?q�>�K?�>?h/���o�}���S�=�n?\��?�:�??�
>���=��Fc�>X�?t��?mG�?p?�9��{�>R�y����>�/��O�;��X>	��=�B>�l?M�?�:�>�w�dI	�;w�<����ؐ��cK=�&
>w�j>�e�>,-L>�ʻ=�kR<�ެ=�8>��>%�>��Q>�Ӭ>���>�����8��?T<>{��=e�?��g> r�<�>9��!��Z�|��^:���m�ú�=E+�=��/=~7=�H�>��Կ�x�?@�>$��`��>��b}���W2>�o?�cl�J�>
�?�7.�,oo>7#�>�Ne>�~�> B>d=Ӿ͗>5���p!��*C��rR���Ѿ��z>�����%�a��C���j/I��t���`�kj��0���E=���<�G�?=���"�k�j�)�L���'�?M�> 6?䌾� ��=�>���>�Ս>�U�������ō�/~ᾙ�?8��?�c>�>�W?p�?7�1���2�9\Z��u�0�@�l0e�@�`��ٍ������
�o���/�_?��x?�\A?/��<�z>���?��%�F���
�>�)/�a;�J'==�a�>c���h�`��Ӿ�EþN���F>��o?�,�?1L?7jV��0���'>�9?�[-?s�l?�8?p@?j_��kL!?�O;>�?�u?��,?�M0?�?��9>���=�)�<bk=`m���]������ؽ�fS��8=��#=��R�ǁ�<�*=(�E=p���n��y�<.�ּ�;�~
=v!l=-;�=Ĵ�>�]?�o�>�N�>��6?^�� _6��ݫ��Z-?� -=��z�4���K�;?�f>a�j?:I�?�-Z?ωe>C��lG���>혋>q�'>!`^>HT�>���<;H���{=8)>`�>Pl�=OJ�p��	��^�����<:�>u�>�?|>h㌽G�'>���Az��Ce>@�O��㺾3S�W!G��1���w����>��K?��?Z!�=!���̔�O�e�:�(?��;?}M?AC?��=9�ھ��9���J��~�΄�>sN�<�	�򱢿Y=��Xp:�D��:��s>��������F>I�����x�xLJ���Ծ�&�=?�
���C;�����8���� >�f>�㹾 $�Mg���򨿖$I?�@�=Xܟ��J��H��&��=�5�>��>=�d���C�;��~���Jt=i��>�)>����s���}H�T���r�>��C? W\?��?���Wrn�F�K�ޛ�P���=�<�?|�>�?��(>]M{=3���+*�t�`��SD�Y��>#6�>M���Z@��Ύ���k���m�> E?xM�=¨?wL??��?��^?/?̶?���>"*ǽ���.m&?0�?H2�= �Ž� X�!�8��;F��>Bp)?��B�<!�>��?7�?9�%?�Q?>�?߼>3� ���?���>�5�>�V�S8���]>n�H?���>Q�V?���?��4>�C6��䢾㨱���=E,>�3?� ?�?��>_��>�2����= v�>�q?ZM�?`�Z?vN>=$#?�/O>���>���=s6j>��?�#?ܡ[?�s?>E?W�>D?�<���;����~����ֻK��;��=����������=�#=Vɷ;1��<I�L=��L=�� ���=1�8=�m�>j�s>=땾�.1>��ľEX��Ʃ@>MO��;,��񓊾W&:�U�=lm�>�?�ҕ>��"��D�=1��>��>=��UJ(?��?|?T3;u�b���ھ�vK���>��A?�u�=P�l�nr����u�Y�h=.�m?��^?ctW�����>sb?	�]?(�𾐸;��ľ�~c�'e�V#O?ui
?�G�-�>��}?� q?j��>J�c��m���*>b��n��׶=��>�z�c��ޝ>�7?���>H�b>R�=t�۾�=x�d���0�?�w�?��?��?�(>B�n�CM߿��Ŧ��b]e?���>�U��t�?e^����ξz����Kk��I��ħ���0���料�d$��򀾺��hč=$�?Fu?��k?ad^?#)
�v�T�A]������X�w!�C�B�9��:�ҿ?�tUk��h��c��p���U��-�f���Y����??��>[�1��>ꣾ�1�~�ʾi̛>����+�y-���S�i�:�@Q<G�d�S~�Yž�x?oY�>�9�>X�B?,�v�R�B�:���C�<6��S<��4>�^�>���>6��oU������#ƾ�Ѓ�-�>A�Y?��@?VRW?l兾Z'�J3��p\	��*��g�X��Ҡ>�>��>�z-���ݽ�B�wHY��En��>�DRW�����b�
?�>���>Ћ?��?��R���оk���İ/�iO����>�z?8j?l�e>'�L�O��(��>�l? �>��>����^l!��O|�o�нO��>f�>�>�p>�,��\��P��#_��p{9����=I�g?������_��Ǆ>��Q?��M:n@<��>��l�b"���~%�BM>+�?�D�=��<>՜ľ���2{�!���;y1?R�?t]��;	�"�>ɑ?+��>p�>��?�5^>TG\���U>z?��T?I�H?��=?)��>z��=�ܽ�ϼ�L�2�q�=��>��[>o��=��=av�+�P��G&�6í<L�>p��<��=^ӿ<�Y��y�=w�=��=<�ؿ�V��V��?+�%	�/,����&������4E�1��=Ծb���i�ݽӄ;nh:�_���d���#<����?���?�ø�q� ���W�Iy���x�>���� �.����ZQI���������Ͼ�J?���(ƈ���X�,?��#��ȿ�ؔ�W,о�f?�m?��H?1?����U���ڼo/>w+�ǉ(�B�����Ϳ3�۾%|h?�}?��ξa�e�F�?I�>��>b�K>Q��(5̾]�5>-��>�K]?Y�Y?��4��SԿ�����u�=���?.�@�A?�(����"�V=���>ڎ	?/�?>\�0��-�M��4q�>O@�?&��?ʵM=W�W�!��;ve?H�<��F��޻���=TQ�=��=����J>79�>[v�=;A��ܽ��4>�߅>x�!��:���^�4[�<ۈ]>�qսZ���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=����;�ɿ���(��ߦ�<�؎��0<��I��_ӽE$��g��|��^��U&�=���=��h>V݁>�a>�J^>U?��q?��>|��=����.P��z��#"ϻ�n�����~���'��������
�B �l���)�>v��߹�
^\�0�5�S
_�Zt����8�L�Y�U$'�n�1?vv>[ �^�\�+�r�ɺ����a�I�;=m�r��P;g=�}c��g�?��G?V���]�$9&�Pս���<�3X?����~�
���̾�T5=��a���~1�>&V�<[y�\L���Z��c3?%�#?O8��̠���ZF>�Ľ��U=�4?Qg?>r¼	�>�2?�署�˽�8k>v�@>cA�>[��>� >6)������Z?��Q?����鉾�c|>�lľ��o�@�3=�	�=Ѕ0�'�ʼ���>y3a<ߊ���;W����r��R3^?���>N��&�Z�G��,��'�=$��?�?_c>�z?F�V?E�>a�����������>'�L?��e?;r >C�0��g��!���<�0?�w�?埿>��&���V*�����2?���?ܵ�>�!��Յ�U���R� 7?��v?�r^�zs�����`�V�p=�>�[�>���>��9��k�>�>?�#��G�����~Y4�Þ?��@���?��;<1 �_��=�;?i\�>�O��>ƾ{������d�q=�"�>􌧾}ev����R,�d�8?ܠ�?���>	���é�Yb�=
J����?f�s?� ����㼗t-�6�t�Y�侪�y=P�<�m<��㽄����u2�s��������P��Y�>��@]�G�1?Yj��.�Ϳ�cӿrS���!��Kj2��*?��> hռ�'��>�f�.m�+B��3N���l�dO�>h�>����%��{��o;�U��7�>�����>6�S�j%��8�����6<��>��>���>s)��lｾ���?�c���9ο����.����X?�c�?o�?'v?t:<L�v��u{�f���2G?Z�s?[Z?�x%�3$]�&�7�9�[?vcj����1@���R��W�>��'?��!>��,�m�>���:H?��
>�Wc��ÿ����F���(�?���?7��q]�>���?�!?������/��?<"��b�=Hu#?n)�>uB��aL���9�~b`��"?� ?O8���@�]�_?+�a�M�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�f6%?�>d����8Ǿ��<���>�(�>*N>^H_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?%D�>�
�?oI�=�V�>��=1���C�:�\#>;T�=E�>��?fqM?H&�>�q�=	m8���.�i{F�2XR��=���C��·>��a?OL?�wb>o����d/��� �sʽA�1�9��0�@��/�E�޽�;6>��>>�>�wE���Ҿ�?�r���lݿ�������@o?��>���>��2命� ���l?ߍ?-�/��Ƚ��Ś�*`���?��@+?�����>��=�+t>�2�����k�6��wV>\�>?$�U�	^���$��I�>�?�<@�$�?F�H��	?���P��2a~�ɂ�7����=��7?�/��z>���>�= ov�����-�s����>�B�?�{�?��>�l?��o���B��1=�M�>b�k?ns?�o��󾾲B>*�?�������K��f?��
@\u@)�^?�׿/U����ǾrZ�	@<���<&!�<�*���`I�o.�Vf����۽�~>yp�>K8z>M<�>z�>�m>��3>El������ʵ�������W���'�c�3�1�R|��p̾[�J����Ǿ�A�=�iN=�����4������7k�{N>�B7?��<?f	o?Y��>��߽ڿ='��b��=ԫ���=��>�r�>88?ly$?=��=^3���s�����Ғ��٧���>R�3>���>��>��>4����t
>��P>ʑu>���=,�����=�)]���=���>ӯ?�1�>���=q,�=�㴿�}��s�x�N����9�����?����@V��՗��]��1(��0�=�-?��>�ڐ���ѿ���� D?0������������=�O"?F?��=W@���*u��$&>��#��Jr�ь�=�
��0^��&�}�>>�Y?�Lһr��=��>��W��m�p�߾t�[>��/?P���v�����y��Y�<5ھD��>K�>��<"��ܛ�މ{���J���1F?��,?��=��{�
V��v���	&>�]>��>ͯ�=.E>\M7��4����F�=�4b>��>�?�#>&��=Ѩ>�ꌾ� T�=��> �>>p�4>��@?�g$?�弴4����a�i���>���>^�}>I��=0C��,�=��>A�_>��6��M�&x4�ٵH>������L�D�x��V�=�;��N��=���=V`ݽ�+�{:>=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾI��>�����+Y��_�b���=��>�/?N����?��+f?�!?�k���^���Wп��}����>� �?�?;g��y���V4�UW�>��?�K0?�+>#ﹾ�����i>x�X?�$U?�W�>�����g�?�$�?>5�?�e>g@�?�is?	�>]�m��,�����o��D��?j>��>W�y>K����}D��狿����@�u����^�=qa�=�T�>��v�-���&��;yѽ��H�`=��>{�r>��>�O]>��?d��>r%�>��=�X	� pj��b!�B[K?0 �?E��4g�kq<f�=,�c��4?Q�7?+~���̾��>�V?_�}?wH[?�)�>�K��霿����'D��*�;<A>)�>�7�>_����ZS>��۾ScD��Վ>��>k�$S���~�o��9���>�"?���>gx�=� ?��#?i�j>�0�>�fE��7���E����>Ј�>�R?4�~?c�?�ʹ�Z3�t��?㡿ۘ[�uN>��x?�R?�ɕ>ƍ���~����E�K[I�T�����?�^g?�m��	?)�?P�??N�A?w?f> o��ؾժ����>�"?��/�4�O��ߖ�,��>��>�q�>w�<�qLս����6�x���s?��[? �$?�����i�о���<���㈼�<��<�*>Ͳ*>��ͽ���=0e+>�4=�R~��Y�[=�<ȋ�=��>��=�D�aLf��+,?A!A�6M�����=��r�._D��>��J>�����^?I�=�N�{������1�U��֍?���?�x�?�����h��	=?�=�?5�?�/�>k��-�޾�b྽�v���x�L=��>}?�>Di����y���S����5���SȽ��`�VK�>�|�>+?�X?�6>��> ���O�.�����&�r��%���F�/H�d-�ug��������Wƾ�㳾�>�!4��-�>��>T�>���>���>�U>	C�>��(>�$�>�\�>O�w>��L>��>�V�=2Q7�LR?������'���簰��3B?zqd?�2�>!i�P��������?���?s�?,>v>~h� ,+��n?�=�>A���p
?hY:=���7�<�T������8��X��>5F׽� :�7M�pif�-j
?f/?	��ً̾l?׽x
��e�r=i�?�'?O*�?�O�9^w�@]�A�K�g����Gf�Dc��q%�vo��6������o���W�'��n<��(?��?"����Ӿ�޻��f�HlD��@A>jZ�>���>�3�>�Y>�d�i_0��)^��"����c��>�Iy?3�>��S?�f7?2�U?�V?(�?C^>l�q��?�hF����>_(?�Z?�1?�6?n�?8P:?zMj>��G���ݾ��پ]�?���>��>���>���>����' ����=d�����a����5>�W�<�O��T��=¿��;+�=�b?�
�Z�8�����3k>�~7?���>��>7���!G��	�<^V�>t�
?\.�>b���X^r��Q��d�>ܚ�?F
���=�)>��=n��7A�� #�=/���M��=�r��^<�~+$<WԿ=��=�����f�1�:�W�;@a�<.t�>��?���>5D�>@��� � ���f�=�Y>eS>w>1Fپ�}���$����g�\y>�w�?�z�?�f=x�=���=�|���U���������3��<��?QJ#?�XT?r��?��=?>j#?�>m*��L��t^�������?U!,?���>�����ʾ�񨿷�3�ޝ?'[?�<a����;)���¾s�Խ�>�[/�d/~����D�KՅ�������.��?߿�?(A�T�6�y�ο���[��e�C?	"�>�X�>:�>2�)�_�g�c%�u1;>���>HR?���>$�L?@�u?��W?e�#>��6�Ԧ���9����B���<>=C?�Xy?���?�}k?�>��>�1Y����,��ۊ�pD꽠 ���=��b>q�>�e�>�`�>#;�=W�	�$���@J�V.�=�~>]��>�#�>S"�>�-g>�)d;:[M?��	?ë���辒k��������%c�?�?$4?�1>�- �Z 5��ݾ�!�>���?�z�?q.?��� �=r~g=$<��V섾5��>���>x�>"�= �<w��=/��>��>� ����-���/�U��a��>N,?��<>W�ƿ��x�	�{�� ��jͼ�$��v�`�k����=U���*<�����F��ڲ��%�b���Z��:;��p袾:��>��<��0>J0&>�}�=�^�<"�<���I�"<�^�=��)�|�<��v��  ������R(97�=���=j��<�dɾ
�|?��H?��+?d�C?�v>ښ>�>�a��>�t}��Y?��S>��Z�z6���:�+T��B����;پ��ؾءc�O0���>=�Q��>&�2>S��=SG�<��=_[j=�
�=Ⱥ�b�=��=���=�4�=f8�=Ou>O>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>5�9>%�>��Q���/�S�X��Xc��Z��� ?n�9�խʾ�}�>��=P�W�ľb�2=�;6>��h=HT�I�\��/�=W����7=��c=�j�>��B>Wz�=�������=��J=T[�=AGQ>^���1#�4x*��&4=�p�=qOf>�M%>T+?�?�?H\`?���>����\U۾�Y#���>W��=�B�>/>�=���=Y��>3�K?a�\?�X?9��>���9ķ>�u?����G�F����꽐����?=gq?��=���=��t�������e�Ct0<!(?V�5?z�>ȱ�>�$�o��" �]������]żɚ�=vŪ��6���׽��I�:�i�}��<K��>���>cl�>g�}>�#>A�=>�s�>���=���=$�>��a=]��=P>� ����X���j>j4�;h��;�8˻�����4d���{�<4�=�K�=��=��>��>���>��=�/��7�>v/���VG���=����nSA�b|e�O�����5��]�� >X�r>��yz�� ��>��>��J>c~�?��r?�>�����־R�J8Z�|׌�C�=��0>��1�H:8��F[�.nP�xi�+�>�ԝ>�'K>�k>9+.�Z�>�)�S=��	�»(����>� ��a��[��������圿Y��{>/�L?:,����g=.g�?\4@?�S�?�r�>�"��>���**>I�����a=��8�	[��а�<�?3s?{u�>D��
Z���̾�s��Eз>,�G�M|O�G���o(0�{�
����)f�>2��$Ѿ-3��M������f�B��q��Ȼ>ekO?]��?��c�1񀿍gO�L��B�����?�Vg?�u�>��?Sf?hu���U��A]�=�o?Jf�?��?��>t>�����1�>j
?7�?#�?�-[?�����> a=�2>Ƿ���-�<��T>A�=<�=ѹ?� ?�/�>y���iv�V2־Ի���g?���<�=x��>��>��>sx�=[B$>���=�,�>�S�>$­>C�K>�Q�>�"�>Y�ɾK�.���*?�[ =�>�>xK�>��:>�>`fF=.�>S��=�=���&�����8�%�L��<�L�=���>&�=�3�>z����o�?��q�b�!��>�	�	Y�1W�>/�>�^S����>ba�<���>� ?Z��>�P�=C�>�2>,�>�z�<�٦P���4�
J�^>;�þ-�v��M%�bh�����`uӾ���lj�oύ��[���<�Z�?���<A5����K��>��> 8?�#���ٱ�h�=_��>��>p��S���G���M9ؾc�p?x��?sCc>�>��W?Q�?S�1��3��rZ���u��$A�e�ʶ`�a��������
�;����_?��x?"rA?�<�3z>���?��%�Dӏ�Z.�>�/�B$;��c<=�(�>�'����`�%�Ӿ��þ�*� 7F>ҏo?
&�?P\?�UV���>�v�> uG?�P:?J=q?��F?�\?ܨ�=��G?���=�?ӌ?�i@?R93?�f#?�~�>6�>�<��v�������љ�����Z��Ê<���<�_=��9;+(�=��W=�� <���;�Q`�%�ϒ�;��!=L�=��=�>�_?�n�>̉>fZ6?�8&�7�W&��~�/?�'=��n����k2���'���>��l?Sƫ?�lX?�|e>�<=�31:�>L��>y�&>�Mp>=#�>�罧xI��߀=��>�j*>t��=�⃽�ʅ�<�
��ǒ���<��$>y��>X�v>Yk\��bO>�z��K�r�U>}�u��C��$-�SY>��2��d��d��>�'J?S,?��O=�����_ֽ��\��}?��/?��I?΀?�sv=�̾L�:���P�����c�>���<�H	�ﳛ��M���<�M�= ��>񩝾����F>I�����x�xLJ���Ծ�&�=?�
���C;�����8���� >�f>�㹾 $�Mg���򨿖$I?�@�=Xܟ��J��H��&��=�5�>��>=�d���C�;��~���Jt=i��>�)>����s���}H�T���r�>��C? W\?��?���Wrn�F�K�ޛ�P���=�<�?|�>�?��(>]M{=3���+*�t�`��SD�Y��>#6�>M���Z@��Ύ���k���m�> E?xM�=¨?wL??��?��^?/?̶?���>"*ǽ���.m&?0�?H2�= �Ž� X�!�8��;F��>Bp)?��B�<!�>��?7�?9�%?�Q?>�?߼>3� ���?���>�5�>�V�S8���]>n�H?���>Q�V?���?��4>�C6��䢾㨱���=E,>�3?� ?�?��>_��>�2����= v�>�q?ZM�?`�Z?vN>=$#?�/O>���>���=s6j>��?�#?ܡ[?�s?>E?W�>D?�<���;����~����ֻK��;��=����������=�#=Vɷ;1��<I�L=��L=�� ���=1�8=�m�>j�s>=땾�.1>��ľEX��Ʃ@>MO��;,��񓊾W&:�U�=lm�>�?�ҕ>��"��D�=1��>��>=��UJ(?��?|?T3;u�b���ھ�vK���>��A?�u�=P�l�nr����u�Y�h=.�m?��^?ctW�����>sb?	�]?(�𾐸;��ľ�~c�'e�V#O?ui
?�G�-�>��}?� q?j��>J�c��m���*>b��n��׶=��>�z�c��ޝ>�7?���>H�b>R�=t�۾�=x�d���0�?�w�?��?��?�(>B�n�CM߿��Ŧ��b]e?���>�U��t�?e^����ξz����Kk��I��ħ���0���料�d$��򀾺��hč=$�?Fu?��k?ad^?#)
�v�T�A]������X�w!�C�B�9��:�ҿ?�tUk��h��c��p���U��-�f���Y����??��>[�1��>ꣾ�1�~�ʾi̛>����+�y-���S�i�:�@Q<G�d�S~�Yž�x?oY�>�9�>X�B?,�v�R�B�:���C�<6��S<��4>�^�>���>6��oU������#ƾ�Ѓ�-�>A�Y?��@?VRW?l兾Z'�J3��p\	��*��g�X��Ҡ>�>��>�z-���ݽ�B�wHY��En��>�DRW�����b�
?�>���>Ћ?��?��R���оk���İ/�iO����>�z?8j?l�e>'�L�O��(��>�l? �>��>����^l!��O|�o�нO��>f�>�>�p>�,��\��P��#_��p{9����=I�g?������_��Ǆ>��Q?��M:n@<��>��l�b"���~%�BM>+�?�D�=��<>՜ľ���2{�!���;y1?R�?t]��;	�"�>ɑ?+��>p�>��?�5^>TG\���U>z?��T?I�H?��=?)��>z��=�ܽ�ϼ�L�2�q�=��>��[>o��=��=av�+�P��G&�6í<L�>p��<��=^ӿ<�Y��y�=w�=��=<�ؿ�V��V��?+�%	�/,����&������4E�1��=Ծb���i�ݽӄ;nh:�_���d���#<����?���?�ø�q� ���W�Iy���x�>���� �.����ZQI���������Ͼ�J?���(ƈ���X�,?��#��ȿ�ؔ�W,о�f?�m?��H?1?����U���ڼo/>w+�ǉ(�B�����Ϳ3�۾%|h?�}?��ξa�e�F�?I�>��>b�K>Q��(5̾]�5>-��>�K]?Y�Y?��4��SԿ�����u�=���?.�@�A?�(����"�V=���>ڎ	?/�?>\�0��-�M��4q�>O@�?&��?ʵM=W�W�!��;ve?H�<��F��޻���=TQ�=��=����J>79�>[v�=;A��ܽ��4>�߅>x�!��:���^�4[�<ۈ]>�qսZ���5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=����;�ɿ���(��ߦ�<�؎��0<��I��_ӽE$��g��|��^��U&�=���=��h>V݁>�a>�J^>U?��q?��>|��=����.P��z��#"ϻ�n�����~���'��������
�B �l���)�>v��߹�
^\�0�5�S
_�Zt����8�L�Y�U$'�n�1?vv>[ �^�\�+�r�ɺ����a�I�;=m�r��P;g=�}c��g�?��G?V���]�$9&�Pս���<�3X?����~�
���̾�T5=��a���~1�>&V�<[y�\L���Z��c3?%�#?O8��̠���ZF>�Ľ��U=�4?Qg?>r¼	�>�2?�署�˽�8k>v�@>cA�>[��>� >6)������Z?��Q?����鉾�c|>�lľ��o�@�3=�	�=Ѕ0�'�ʼ���>y3a<ߊ���;W����r��R3^?���>N��&�Z�G��,��'�=$��?�?_c>�z?F�V?E�>a�����������>'�L?��e?;r >C�0��g��!���<�0?�w�?埿>��&���V*�����2?���?ܵ�>�!��Յ�U���R� 7?��v?�r^�zs�����`�V�p=�>�[�>���>��9��k�>�>?�#��G�����~Y4�Þ?��@���?��;<1 �_��=�;?i\�>�O��>ƾ{������d�q=�"�>􌧾}ev����R,�d�8?ܠ�?���>	���é�Yb�=
J����?f�s?� ����㼗t-�6�t�Y�侪�y=P�<�m<��㽄����u2�s��������P��Y�>��@]�G�1?Yj��.�Ϳ�cӿrS���!��Kj2��*?��> hռ�'��>�f�.m�+B��3N���l�dO�>h�>����%��{��o;�U��7�>�����>6�S�j%��8�����6<��>��>���>s)��lｾ���?�c���9ο����.����X?�c�?o�?'v?t:<L�v��u{�f���2G?Z�s?[Z?�x%�3$]�&�7�9�[?vcj����1@���R��W�>��'?��!>��,�m�>���:H?��
>�Wc��ÿ����F���(�?���?7��q]�>���?�!?������/��?<"��b�=Hu#?n)�>uB��aL���9�~b`��"?� ?O8���@�]�_?+�a�M�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�f6%?�>d����8Ǿ��<���>�(�>*N>^H_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?%D�>�
�?oI�=�V�>��=1���C�:�\#>;T�=E�>��?fqM?H&�>�q�=	m8���.�i{F�2XR��=���C��·>��a?OL?�wb>o����d/��� �sʽA�1�9��0�@��/�E�޽�;6>��>>�>�wE���Ҿ�?�r���lݿ�������@o?��>���>��2命� ���l?ߍ?-�/��Ƚ��Ś�*`���?��@+?�����>��=�+t>�2�����k�6��wV>\�>?$�U�	^���$��I�>�?�<@�$�?F�H��	?���P��2a~�ɂ�7����=��7?�/��z>���>�= ov�����-�s����>�B�?�{�?��>�l?��o���B��1=�M�>b�k?ns?�o��󾾲B>*�?�������K��f?��
@\u@)�^?�׿/U����ǾrZ�	@<���<&!�<�*���`I�o.�Vf����۽�~>yp�>K8z>M<�>z�>�m>��3>El������ʵ�������W���'�c�3�1�R|��p̾[�J����Ǿ�A�=�iN=�����4������7k�{N>�B7?��<?f	o?Y��>��߽ڿ='��b��=ԫ���=��>�r�>88?ly$?=��=^3���s�����Ғ��٧���>R�3>���>��>��>4����t
>��P>ʑu>���=,�����=�)]���=���>ӯ?�1�>���=q,�=�㴿�}��s�x�N����9�����?����@V��՗��]��1(��0�=�-?��>�ڐ���ѿ���� D?0������������=�O"?F?��=W@���*u��$&>��#��Jr�ь�=�
��0^��&�}�>>�Y?�Lһr��=��>��W��m�p�߾t�[>��/?P���v�����y��Y�<5ھD��>K�>��<"��ܛ�މ{���J���1F?��,?��=��{�
V��v���	&>�]>��>ͯ�=.E>\M7��4����F�=�4b>��>�?�#>&��=Ѩ>�ꌾ� T�=��> �>>p�4>��@?�g$?�弴4����a�i���>���>^�}>I��=0C��,�=��>A�_>��6��M�&x4�ٵH>������L�D�x��V�=�;��N��=���=V`ݽ�+�{:>=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾI��>�����+Y��_�b���=��>�/?N����?��+f?�!?�k���^���Wп��}����>� �?�?;g��y���V4�UW�>��?�K0?�+>#ﹾ�����i>x�X?�$U?�W�>�����g�?�$�?>5�?�e>g@�?�is?	�>]�m��,�����o��D��?j>��>W�y>K����}D��狿����@�u����^�=qa�=�T�>��v�-���&��;yѽ��H�`=��>{�r>��>�O]>��?d��>r%�>��=�X	� pj��b!�B[K?0 �?E��4g�kq<f�=,�c��4?Q�7?+~���̾��>�V?_�}?wH[?�)�>�K��霿����'D��*�;<A>)�>�7�>_����ZS>��۾ScD��Վ>��>k�$S���~�o��9���>�"?���>gx�=� ?��#?i�j>�0�>�fE��7���E����>Ј�>�R?4�~?c�?�ʹ�Z3�t��?㡿ۘ[�uN>��x?�R?�ɕ>ƍ���~����E�K[I�T�����?�^g?�m��	?)�?P�??N�A?w?f> o��ؾժ����>�"?��/�4�O��ߖ�,��>��>�q�>w�<�qLս����6�x���s?��[? �$?�����i�о���<���㈼�<��<�*>Ͳ*>��ͽ���=0e+>�4=�R~��Y�[=�<ȋ�=��>��=�D�aLf��+,?A!A�6M�����=��r�._D��>��J>�����^?I�=�N�{������1�U��֍?���?�x�?�����h��	=?�=�?5�?�/�>k��-�޾�b྽�v���x�L=��>}?�>Di����y���S����5���SȽ��`�VK�>�|�>+?�X?�6>��> ���O�.�����&�r��%���F�/H�d-�ug��������Wƾ�㳾�>�!4��-�>��>T�>���>���>�U>	C�>��(>�$�>�\�>O�w>��L>��>�V�=2Q7�LR?������'���簰��3B?zqd?�2�>!i�P��������?���?s�?,>v>~h� ,+��n?�=�>A���p
?hY:=���7�<�T������8��X��>5F׽� :�7M�pif�-j
?f/?	��ً̾l?׽x
��e�r=i�?�'?O*�?�O�9^w�@]�A�K�g����Gf�Dc��q%�vo��6������o���W�'��n<��(?��?"����Ӿ�޻��f�HlD��@A>jZ�>���>�3�>�Y>�d�i_0��)^��"����c��>�Iy?3�>��S?�f7?2�U?�V?(�?C^>l�q��?�hF����>_(?�Z?�1?�6?n�?8P:?zMj>��G���ݾ��پ]�?���>��>���>���>����' ����=d�����a����5>�W�<�O��T��=¿��;+�=�b?�
�Z�8�����3k>�~7?���>��>7���!G��	�<^V�>t�
?\.�>b���X^r��Q��d�>ܚ�?F
���=�)>��=n��7A�� #�=/���M��=�r��^<�~+$<WԿ=��=�����f�1�:�W�;@a�<.t�>��?���>5D�>@��� � ���f�=�Y>eS>w>1Fپ�}���$����g�\y>�w�?�z�?�f=x�=���=�|���U���������3��<��?QJ#?�XT?r��?��=?>j#?�>m*��L��t^�������?U!,?���>�����ʾ�񨿷�3�ޝ?'[?�<a����;)���¾s�Խ�>�[/�d/~����D�KՅ�������.��?߿�?(A�T�6�y�ο���[��e�C?	"�>�X�>:�>2�)�_�g�c%�u1;>���>HR?���>$�L?@�u?��W?e�#>��6�Ԧ���9����B���<>=C?�Xy?���?�}k?�>��>�1Y����,��ۊ�pD꽠 ���=��b>q�>�e�>�`�>#;�=W�	�$���@J�V.�=�~>]��>�#�>S"�>�-g>�)d;:[M?��	?ë���辒k��������%c�?�?$4?�1>�- �Z 5��ݾ�!�>���?�z�?q.?��� �=r~g=$<��V섾5��>���>x�>"�= �<w��=/��>��>� ����-���/�U��a��>N,?��<>W�ƿ��x�	�{�� ��jͼ�$��v�`�k����=U���*<�����F��ڲ��%�b���Z��:;��p袾:��>��<��0>J0&>�}�=�^�<"�<���I�"<�^�=��)�|�<��v��  ������R(97�=���=j��<�dɾ
�|?��H?��+?d�C?�v>ښ>�>�a��>�t}��Y?��S>��Z�z6���:�+T��B����;پ��ؾءc�O0���>=�Q��>&�2>S��=SG�<��=_[j=�
�=Ⱥ�b�=��=���=�4�=f8�=Ou>O>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>5�9>%�>��Q���/�S�X��Xc��Z��� ?n�9�խʾ�}�>��=P�W�ľb�2=�;6>��h=HT�I�\��/�=W����7=��c=�j�>��B>Wz�=�������=��J=T[�=AGQ>^���1#�4x*��&4=�p�=qOf>�M%>T+?�?�?H\`?���>����\U۾�Y#���>W��=�B�>/>�=���=Y��>3�K?a�\?�X?9��>���9ķ>�u?����G�F����꽐����?=gq?��=���=��t�������e�Ct0<!(?V�5?z�>ȱ�>�$�o��" �]������]żɚ�=vŪ��6���׽��I�:�i�}��<K��>���>cl�>g�}>�#>A�=>�s�>���=���=$�>��a=]��=P>� ����X���j>j4�;h��;�8˻�����4d���{�<4�=�K�=��=��>��>���>��=�/��7�>v/���VG���=����nSA�b|e�O�����5��]�� >X�r>��yz�� ��>��>��J>c~�?��r?�>�����־R�J8Z�|׌�C�=��0>��1�H:8��F[�.nP�xi�+�>�ԝ>�'K>�k>9+.�Z�>�)�S=��	�»(����>� ��a��[��������圿Y��{>/�L?:,����g=.g�?\4@?�S�?�r�>�"��>���**>I�����a=��8�	[��а�<�?3s?{u�>D��
Z���̾�s��Eз>,�G�M|O�G���o(0�{�
����)f�>2��$Ѿ-3��M������f�B��q��Ȼ>ekO?]��?��c�1񀿍gO�L��B�����?�Vg?�u�>��?Sf?hu���U��A]�=�o?Jf�?��?��>t>�����1�>j
?7�?#�?�-[?�����> a=�2>Ƿ���-�<��T>A�=<�=ѹ?� ?�/�>y���iv�V2־Ի���g?���<�=x��>��>��>sx�=[B$>���=�,�>�S�>$­>C�K>�Q�>�"�>Y�ɾK�.���*?�[ =�>�>xK�>��:>�>`fF=.�>S��=�=���&�����8�%�L��<�L�=���>&�=�3�>z����o�?��q�b�!��>�	�	Y�1W�>/�>�^S����>ba�<���>� ?Z��>�P�=C�>�2>,�>�z�<�٦P���4�
J�^>;�þ-�v��M%�bh�����`uӾ���lj�oύ��[���<�Z�?���<A5����K��>��> 8?�#���ٱ�h�=_��>��>p��S���G���M9ؾc�p?x��?sCc>�>��W?Q�?S�1��3��rZ���u��$A�e�ʶ`�a��������
�;����_?��x?"rA?�<�3z>���?��%�Dӏ�Z.�>�/�B$;��c<=�(�>�'����`�%�Ӿ��þ�*� 7F>ҏo?
&�?P\?�UV���>�v�> uG?�P:?J=q?��F?�\?ܨ�=��G?���=�?ӌ?�i@?R93?�f#?�~�>6�>�<��v�������љ�����Z��Ê<���<�_=��9;+(�=��W=�� <���;�Q`�%�ϒ�;��!=L�=��=�>�_?�n�>̉>fZ6?�8&�7�W&��~�/?�'=��n����k2���'���>��l?Sƫ?�lX?�|e>�<=�31:�>L��>y�&>�Mp>=#�>�罧xI��߀=��>�j*>t��=�⃽�ʅ�<�
��ǒ���<��$>y��>X�v>Yk\��bO>�z��K�r�U>}�u��C��$-�SY>��2��d��d��>�'J?S,?��O=�����_ֽ��\��}?��/?��I?΀?�sv=�̾L�:���P�����c�>���<�H	�ﳛ��M���<�M�= ��>񩝾�g��2LO>"V�$�߾�k��sB�ưվ��[=����B=ޡ��<��Ԁ���=�}>��t �sF��c4��SwJ?�[�=F��<�o��F���!>���>V�>�Ǎ��Ø�	�>�������=÷�>_�4>������[J�c@�1��>;<?�kX?�%�?0�\�c�d�:4>��kﾑ��O_*�F�?lH�>9 ?C�}>kz�=����?�	�-�\���F�v��>���>"���uM�����3����}�?��>�?�C�=��>�A?��?̩e?�1?�
?��f>o/��0L����2?Bc�?Ѿ";2b;�+ D���E�h�=���;?֊C?H!���G�>���>���>ʺG?d�s?ن'?-�;>߫��DR����>�r�>��e����P��=wf
?e�i>�y?�M�?%�h>�=*�&��,Y��r��=>�Y.?�]5?��?=z�>�`A?�����0>��7?�a{?���?G�%?���>T�?tU�>��?�b+>0Ў>��?�+ ?��G?���?Y?�{>�f=;�<����>�=x =��<@���/^>�u>�q:�T���a4=�� >ၽ��8�FOԽ��=�=s��_�>n�s>�	����0>_�ľhO����@>�y���O��U܊���:�[޷={��>,�?���>�W#�ܳ�=���>fH�>���6(?k�??{;!;<�b�2�ھ��K���>,B?���=��l�,����u��h=��m?a�^?8�W��'��-�b?<�]?iX��=�+�þ��b����f�O?��
?��G�!�>��~?��q?I��>N�e�<-n����>b�C�j�w��=�v�>�Z���d�r+�>)�7?K�>c>};�=�۾O�w�*p���?��?
�?7��?.*>6�n�%-��(�����V `?���>s՝�iQ?�ɻ�Ҿ_����3��Z}޾�����G��U݌�6��|{���4��<�=/O?dr?Z�q?��b?����0e��r`����'�U��d�����C�`�F��.D�7�p�����=������ֆ=`����X�FĶ?q��>�F.<��>��{��󨘾d��=|�������<�=3��=N�X=�v>G�>��,L�㭳�.�?V �>�w�>��P?V�c���O��D�?��c�b>�h�>s�>�T�>us3����=�nV�rKV�`w�一>&%Z?��L?�~k?*�D��8D��쇿�n+�/G*�2HT�d�R>�H2>�]�=
)^�����a`��,D��Mm�g���y��Y7����-�?�f�>ӛ�>���?���>e�ʾSH��[���*��]=R1�>%�f?@	?�ِ>:�:��B��>y�k?R:�>D��>ď��"��}���׽��>G�>�� ?��y>i�3��]�Nߎ����O�8�D�=ݗf?p̂��k^��ǅ>:�Q?R�q�?�<v/�>
�]��!�8~�!��+>��?�y�=(�@>��þ�3���z��L��J#;?�84?L���>q.��=�>��?��>ɝ�>���?�s=����'0�=Ӳ?4 Y?��Q?�V?+?��=�:�o̽:�@��>fr�>4'�>��!>�{5>��f��s��%☾�Dk>�Bz>鯈=�t~��Ĉ=��$�֨���F=&}`>�ۿHTU��>�N���������T�N2��gf���V���վ��Ѿ��[���u��J����b� z��#�a��O�?��?����������,\�L�Ծ��>����|*���þ��I�����"̾ʃ��e!��Oh�-4��`�_��P�>@
���Pο�������gxA?�57?V)?+HB����{i���=:�>��S��9�F&��-�Ŀh+𾂕�?u:�>��׾1�<��V�>�(\>����fW>��������VP=�R�>qeA?"�1?�f?��!��嫿sW���?ہ@�A?��(�G�쾉�X=H��>Ҙ	?�?>U�0���6İ��P�>�1�?|��?HN=)�W�����e?!K<��F�#߻h�=g�=ܭ=<��P~J>jh�>���AA�+�۽Cu4>*��>��"��5��M^��L�<��]>j�Խz䔽5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=u6�����{���&V�}��=[��>c�>,������O��I��U��=�i��[Կ�I.�K�	�������o�߾>'EY�,�x��=QU��B�Ͼ�5�i��<X8	>�>�v�>#+>eCU>�AW?)s?4,�>�N̻�Z2<����$������
۾IԾ!��bz��D6¾e
þ��۾�	����=��O������?�&�X=¹R��ҏ�.� ��u^��t>�Yl-?��>l�̾�P��y���!̾���(?�����ݽ̾��5�Ԙk��@�?��D?�_���\Y�}���҇�6���q�S?��se�``��_��=Z���oW=���>�=�����7�E�Q��O5?�y'?4������#WU>���;�<�^4?Z��>�lý��>�@+?� 꽵>t�,��>X�c>��>�{�>	.�=F)�����4!?�#c?v�ʽ����y��>���?$���jv=�HB>���dN��JC>�K={��D[�I����<-)W?Y��>y�)����]����AN==Ӳx?�?k'�>vyk?��B?��<�b��l�S��F�w=J�W?�%i?��>j���Aо1~��J�5?�e?��N>�nh�w����.�eQ�&?��n?�]?({���t}������xn6?��v?s^�vs�����;�V�i=�>�[�>���>��9��k�>�>?�#��G������wY4�$Þ?��@���?��;< �T��=�;?h\�>�O��>ƾ�z������+�q=�"�>���ev�����Q,�e�8?ܠ�?���>���������=�թ��3�?��t?�ߜ��V.�����zy��hϾA!�;_ 2>z�
>��p���x5;��x��A����1��S��>�@ϗ�~%?(��$�ǿ..߿�	����b�D<̔ ?���>��x��Cz����M�K�� \�7aP�hc�>j>/I��gN����z���:�mT�� ��>����G�>��R�-������ڜc<�T�>���>���>؋���<��}��?Dc��*
ο����9��6X?�1�?���?�6?��<F�w�a�{���� �G?��s?� Z?J{-��^�NL7���T?K4���s��y6�K��u9>�*;?z�>�@�%�;5Й��?���> 9=��ɿ�7��g��zۗ?��?�����>���?l�4?U!��������C��";'D(?���=m��!H���I�vԂ�P?$� ?/Y�����_?��a���p���-�2�ƽ�ۡ>�0��d\�H��+���We�����?y����?�]�?�?^��� #��5%?l�>]���B9Ǿ���<M�>�'�>j*N>�7_���u>#	���:�
h	>Q��?�~�?�j?b��������S>q�}?a$�>��?p�=	b�>c�=��X-��j#>}"�=��>��?��M?tK�>�V�=F�8�d/�E[F��GR�n$� �C���>?�a?��L?�Kb> ��O2��!��tͽQc1��T鼰W@���,�S�߽�(5>J�=>W>��D��Ӿq�?�o�?�ؿ�i��Ur'�+54?��>�?�����t�k;��;_?�}�>l7�<,��&��*G�֙�?H�?��?��׾a*̼�>��>yF�>� սf���၇���7>��B?z�6D����o���>A��?��@�ծ?�i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?�Qo���j�B>��?"������L��f?�
@u@a�^?*��տ��3ξ�D���?��>Xh�H�F>Z�\�� >n|r>{�j<j2��c3>Խ�>��>�^�>��>"@t>��=ku��ӎ!�vH��ӆ���;f��:A�
��=�t�*���20<}%�z�����޾A �ߕ��1��*0(�<�.�o�=���=�
E?{�K?��o?QZ�>�:��h�=�4�ǵ�=3���T'�=�t�>�?��E?�+(?��=}��	�c������{��O͎�9�>�_]>���>���>���>:�~�G>��#>m�n>��=�H=9fݼ`�#< >=�>-�>�.�>��=�2�=1��	v����e���"��q=�y�?��ʾ-G�� ���־�����=u�%?�k>��5+ֿ�� NK?-0,�Yn�򣁾�R�=Y�8?6�L?&,�=cr̾��2��f>��ҽ1f+�PZ=2}7��z���9���>1 ?�|f>�t>�3�Bj8���P��Z����|>�-6?���#Y9���u���H��`ݾG5M>߿�>�-C�q�J����>i���|=Qm:?�o?UY������=�u��O��q+R>�>\>P=e��=mM>�-d�L,ǽ�@H��}-=���==�^>I7?�)>���=�>�>i����L��ۧ>��?>µ->�@?:�$?�	��қ��M���=+���v>�"�>�.�>o�> PI�O[�=M�>Ża>Ό��~}�]���>=���V>���"8_���|��7=�W�����=�ݐ=��I!9��#=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾUd�>fp�g\�����F�u��#=w��>�1H?(a����O�">�t
?�?ob�D����ȿ�~v� ��>U	�?	�?��m��=���@�)s�>Л�?�cY?I`i>�d۾>RZ���>0�@?�	R?��>�9��'���?�޶?Y��?R�E>�x?���??�-۾.�`�m��AR��lB9��:�>�R?A6 ?u�*��k�\p��/l�2U�6���	i=���=d�>�tM���m�We;r���3F����<�7>��>0Q�=X��<��>N�>� �>;��=j�q�Ja�$0L?�я?����m�g��<P��=_��(?��4?3W�ξ�(�>�[\?H��?�d[?ð�>ڽ�Kۚ�v������sT�<5L>S��>&N�>���.L>�վE�E�ύ�>�6�>l ���Rپ�����ǻ[ܜ>�!?���>Y��=�� ?#?�j>�,�>�bE�#:����E�6��>���>�J?��~?��?$ڹ�I[3�����塿�[�d7N>	�x?�T?�ɕ>ߎ�������OE�CI�,������?Arg?HO�K?�/�?L�??��A?+-f>e��
ؾ������>N�!?e���A�5(&��}�z{?&5?���>�����pֽO?ռ��tJ���#?y&\?b8&?ۄ��a��þ��<����Wo���;�J��T>�>t���K��=�A>���=�Um�K�5�w�p<�h�=c��>���=3[7�r��0=,?��G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>$�l���K���ڙ���F��_�ŽwM��W��>�>X`�>ya�>$�[>��>֗7��!���C�ɾ47]�X
�	33�`6?�H�R�����L�=��>漯����c�>���5N�>_��>��">�W�>�{�>��>v�
?�\�>''�>n��>� �>Ż�>��>�E=�J�aHR?����ϲ'���U����-B?jdd?%3�>��h�ˉ�����]s?���?Ux�?�`v>cjh��#+�ea?��>����t
?]�9=���mo�<�o������Y��ū�Z}�>�e׽�:��M�^9f��u
?�4?�:���̾7a׽�\��M|=S�?Pd)?��*�G�R��qq���Y�mP��K�+Z�2��Pw&�p�n�(̏�R����S���g%�UE=h�)?rn�?1����I����g�Z?C��g^>A?�>��>�b�>2�P>�
���4�;�[�w.(��Ѕ����>j�z?�
�>V�@?0;8?�(Q?��K?겒>р�>4����>�H=#��>m��>��,?q6*?�/?�i?�r,?�^K>���"8����׾�4?�`?[�?��?��?���/ý��B� ���oe�FB(=���;�F��`���@=�=X#O>&?���$9��=��}'j>�u7?f��>A��>���R/��ŀ�<=��>�c?�L�>� �Q�r�a����>���?����5=��*>u`�=����� ��~��="Ƽ.{�=�}��B���=<���=��=;���b��D��:}��;��<�t�>!�?ߔ�>aD�>dA���� ���s_�=6Y>�S>�>�Cپ�}���$��k�g�	\y>Nw�?�z�?o�f=��=���=�|���T������������<ݣ?�I#?_XT?F��?(�=?�i#?t�>v*�:M���^��\��ɮ?!)?|3�>����Ͼ6�����.�%�?Wp�>SId�NU�ϯ/�������m�M��=��5�����6��r�?��0T=P���z�����?B�?����;�&o�!I������%�??���>���>��>[,��d�����7>j��>ȭN?|��>��5?-n?�W?6�.><�3�"lL����5=%D�>rM0?�Jt?^?��g?Q��>�[6>�������*�<ွ(H�[����U�=��>	��>��?U��>�V>�;M��>½-�]��ʻ=�y>���>9�>g=?}hq>� =~�O?y?�Ѿ�I�:������E��K��?_P�?K{?�#�<�r�_'8�ؠ�����>
E�?�;�?Ś?@�����=�<�����Ql�J'�>��>蠰>�Z�p���7>ݰ�>V�>I�Z�����M���ۼ��?�B?�c!>�ſ��q��p�آ����h<qВ���d��g����Z�H�=���@���۩���[�3���fY��I�������`�{����>�q�=��=���=9�<>Ǽq��<�#J=)�<��=K1p��g<t�8���׻zf��dJ(���Z<�J=�����/ž��u?�F?��.?D�F?:ă>�l>�~��˚>�VT�B?ScM>u��l�����3�<ݦ�(���iCվnpݾq_�[��	�>>78��>}�5>�n>2�<��=}�=m�=�#1��GF=ͨ�=R�=��=���=�%">Ɲ>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=J����=2>s��=v�2�T��>��J>���K��C����4�?��@��??�ዿТϿ7a/>�Y7>�>p�R�wm1�]i\��Zb��|Z��!?	1;�u8̾�@�>���=�߾��ƾW�-=|�5>Ǆb=���3\���=B�{�Z<=1^k=c�>�D>�^�=u���ζ=z�J=S��=�$P>���C7��P*�4�5=U��=��b>4&>W��>�A
?Q?"?\\P? X�>�Q��������`�>�����>6�5=/V>�8?r,??�[B?�$7?�H�>)�¼�\�>5�>�P3�z�y�'� �\�⾋kZ�*��?J��?�nv>`��&�Ȫ��%�ݹk=��?�?ܙ�>0b>{�2��i�&�>�,������s�J=.�m�?�>�#�w�F�����B�=�>R��>�ɡ>p�>e;>�N>bk�>�>���<Ŕx=[�;��<W
���τ=�"ļ��}<�����+���^�
�4�hvѼ��; A����HRP<���=:��>#<>���>Ԓ�=���~B/>繖�|�L�Y��=H���+B�
4d�:I~�$/��Y6�^�B>?;X>�z���3����?(�Y>m?>G��?wAu?!�>#���վlQ���=e�>[S���=�>	�<��z;��X`�n�M��}Ҿ݀�>���>�=*>��(>98(���4����=�;���N��	�>Z��ߜ�t��=r���ˬ�᳥�:y�>r�=�m?(`��ԩ�=菙?C�@?��?�,�>Z:@�}�����[>����ִ�>�LK���6��<֧$?�
?~��>�َ���u��I̾����޷>�AI�3�O�����?�0����ͷ�N��>������о�#3�Lg�������B��Mr�#��>��O?W�?�;b��V���TO����()��q?�zg?��>L?PB?����s�o��$��=��n?��?$<�?q>�@Z>Y���\�>�f?y6�?2?��_?����?/_�=8YA>�.��� =��T>�1d>JKe>n�?JY?�~�>��r��T
� ��V>Ծ�oٽJ�	>s>t��>>��>���>u��=��=�x�<��>YK�>��>_v>���>/ �>.Kž�O�-O'?������> ?H�>��"<]�x��7��y;`=�`�����<���<X����W(=&�=�Tf>8��=t�>�X¿�?vi=��P���>K���p����>naH>X�B��O�>v<>=��>�p�>�]*?)�R>b��>��h1����>�="�<D��TJ�`)��J^��7U5>w�����O�sc)�9:��f.:�"�Ӿ����q�Q�c׆�|ps�8��=��?��=�	d�0.6�T½|�?#�>�?3
t�Q璼8��=��?�{�>eJ
�[���ć���Z�'��?c��?�;c>?�>�W?7�??�1�3��uZ��u��'A��e��`�R፿������
������_?��x?�xA?�G�<�9z>"��?��%�2ӏ��)�>r/�d&;�BC<=++�>�*���`���Ӿ�þ�7�sHF>$�o?%�?~Y? TV���O�2D>�8?��5?:w?�I3?t�4?�)�%?`�<>̴?��?�)?L�'?�%?C+(>�U>D���><g��5k������������û��N=)�=��;��)��;�u#=�~�'z�D�f:���<<�[:=���=к�=�B�>��Y?�.�>fl�>�8?�"�p�7���H�/?N�X=*��-ᇾ>��)��3>o�h?�׫?��W?}U>s�@�T�B�S�>K�>�/>��c>l�>�:�� <I���m=p�>>{
�=Ғ[��Ă�i^	��H��y=��>���>4�{>F���2(>N.����y��"d>`eR������FS��G���1�:�v��C�>t�K?\�?b�=c�W%���,f�q)?�C<?dFM?��?�P�=�B۾(�9�B�J���k�>��<����������:��b�:�\t>����׾�'	>Pa�}�۾k;S��4?�̾��e:(�)�96=�b����ʾz��=D�2>æ��/E1��V������1�I?+�:>S�����</�lg0>]�>�ĕ>D9����:���o��e�C�;���>�Q=�Z���� ���J�˩쾗؍>y�A?N�V?΁?A&s�_V_�K�;������by��#��P?�y�>��?�Ή>���=	���#��[�T��H�6��>�p�>���$�N�jƾ��!�
�f��>���>]�>�?r�]?� ?��p?��$?w"?�F�>�(<s�����2?��w?�Q�=�� �پ�]=���K�I?��2?�����>)�??g	=?BqP? \M?��!?�Y�>�P����D���>���>�^��a����A>}?5Q�>�ׂ?9o?E>�2��Y���ý )W�hK|>�k6?�'+? v
?��>�]?2E��e*
�r�?މX?(u�?93r?J��=��)?���>�hp>�H<c�>�3.?	vB?��_?
�`?(#+?P�>���<QE.��糽W��:��=@�M>����̃�қl�r߬<�Ș�� �;n�u�<N�e���#�m�=�%�=d9X='P�>jDt>z*��1�0>�žHY���~@>���Y���⊾�;���=�h�>��?�]�>�~#�3��=���>o��>���n(?�?:?��,;Ūb�<�ھW�K�=�>d�A?��='�l�Y�����u��Bi=��m?Jl^?��W��`���b?��]?{f�%=���þ �b�Պ龎�O?��
?��G���>��~?��q?ʶ�>��e�*:n����Cb���j�ж=r�>/X��d�o?�>��7?�N�>��b>�'�=�u۾��w��q�� ?i�?��?���?�**>w�n��3�\��������^?K��>�t��	"?�NĻ0�о�ˉ����x�߾M;�������U��m���C#�ׁ��ҽ#��=��?�3s?�5q?n$`?�� �#d���^�/��P*V�������`�D�,^D�ED��m�M��Ҙ��l����==
z��V�dh�?�
?I��<^��>�>^��N�6����s�=z�?���,���=�p���*4<�q�=I�W����Q��7�?�$�>���>z�B?�hP��!F��	E���;��(�9c�>z*i>��>�v�>Z���2���8�s����("�@�>�i?EK?�LT?�^���2�����=��=�=�!=���»���=n$)>�Ӊ�{v����A��Y�A���B��N���9A���"?�
u>�c?wɏ?���>u�����=8���a��=Z��>��Q?" ?t�>�罏��v�>�Ad?��?�=�>>���U`1���������J��>`f�>�?p_>?�3�zj��Џ��K��0k4�a��=��V?��k��1��G1>�2?�+���,=�
�>�ħ��*,��'�i]ӽ��D=IQ?7�6>���=�뾾�;���t�kr��(E?��)?!]ž8��S��>?���>�B?�~}?��+���ʾ���>'AE?��O?�C?��S?�-?|�m>��a�rڽ��I�9hR�֝�>EP�>�&�>I�4>��[��׬������=|F�=��{=�	�濽��Y���u�kP=]�[>�aۿ�K�@�ܾ'���"�ɝ��↾�b���o����
�F����l��M܂���,���M�bh�Ob���%r�W��?a�?H���Ɖ�+噿����N��n��>o�g��Ր�H���a	����CH߾�����#�v�P���i��Ie�L��>��ҽBͷ�
K��{f뾨"?�>E?��5?M�/����Ea�U�����<�2�P%������ӿˡ�����?��?����/;��W�>��>��=f��>57[����:��>�`?��W?:���Կ:�¿�|C>��?ap@>}A?3�(����GV=N��>��	?��?>�F1�F�(��T�>�<�?x��?8�M=U�W��	��~e?��<��F��ݻ��=C�=�9=�����J>�X�>�u�XA�G3ܽ]�4>�م>Br"����S|^���<ʊ]>U�ս':��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=u6�����{���&V�}��=[��>c�>,������O��I��U��=�E���ɿ)pM�t(���=ʇ=�9��`��г���;���;�hs�GY��o�=-��>푿>$yf>��E�& >�ZU?�Op?	��>�0�=Zac�~�+�"U�� ��=�Sڽ)�i�v��$}��}���˾V�ҾR�891��/�w�߾�t=���=�:R��b��$[ �̀b��%F�G.?�� >jnʾ�M��k<�˾Se���w��o���;�-2�5Tn���?�7B?����W�&N�'���G���)W?�����M/�����=���d=���>�D�=�}�q=3��S�y+;?׮%?�aʾF(��cw�>�����=�G?�/�>��Q+�>%U<?�E�<�����s>g>���>���>��=����G�UI)?��T?���@�e�~|�>����	{��L�=p}o>,�|�����>F{'=�����ns��?����/*W?Ҧ�>��)���T_��r��Pf==�x?��?&�>�rk?�B?��<0Y����S����w=��W?�#i?7�>���о�z����5?�e?��N>)hh����.�$R�� ?�n?�V?i۝�7p}�������3o6?��v?�r^�ss�����<�V�A=�>�[�>s��>��9�[k�>��>?{#��G������Y4��?z�@���?��;<�"���=�;?�\�>�O�\?ƾ�{�������q=y"�>x���zev����Q,�x�8?堃?���>��� ���!�=�Y���J�?�<�?�KM�`�9�|�'��Lt���Jc~>t��=Y��<�P����0���ؾ�ھ�_z�g-���Ɍ>�@H���w2?!����ѿ����W�/&޾��g>���>+ �>��A�w��(�X�,I���U�b�I������`�>��>�0���ӑ���{�ya;��ß��>���r��>�;S�P���3���C<��>H��>;��>j���� ��Ѻ�?�O��c-ο��������pX?'a�?�?'X?��:<��v�{�i�5G?�zs?�Z?Q�"�#�\��Z7���_?�`~���f��<�1�O��%N>�-?�>��/�׫�<M��<ju�>�\>�G��,¿/��axǾ�˪?H.�?�&��h'�>�+�?{8?(�7ܜ��H��R�(�b[1=|�3?RZa>�Ͼ��4�!�5�1F���?�0?�����1�]�_?+�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?Ե�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�i	>���?�~�?Qj?���� ����U>
�}?_,�>��?���=�\�>��=x����2�xH#>2/�=-�>��?�M?3�>��=�8�//��^F�MER�,(���C�Q�>��a?D�L?�ab>0����1� !��)ͽX�1����pA@�[,�QD߽>D5>H>>�>��D��
Ӿ��?�ƾ��Կ�*����Z��d?�~n>3��>��	��h���c���iN?*4�>�,��n���ŕ����wR�?z�@���>3*��-a%��&>��>Ɠv>&�žz���Ph�x�>�$?D��w⌿������>=2�?@@r*�?�$i��	?B��O��b^~�Ҁ�1�6�4��=��7?D2��z>���>�
�=fov�E���.�s�!��>�B�?${�?8��>��l?�o��B�=�1=�J�>�k?�s?��l�+󾟹B>�?��������I�4f?��
@-u@�^?��Q#ѿ6����;-W����><|�=2i>wy�����=^ix=l�C=�A�=��>��>�V>�ۇ>d�d>�D@>*M>^����l%�����L��`q8��+�1��WtI���������S��aˎ���6�Y˽������r�?u���2�>S�R?�mM?Q�r?w�>,g�t6�=@H�/�=�_�2.i=���>��0?A:J?��$?a�=*����`��,��r���'|�����>��%>B��>�>���>n7.="��=�>�3�>�S>a�=���=,?R=�A>²�>�D�>�I�>D�2>��>�,��Oİ�	Xh�>�w�(�½|p�?^����J�%���������H�=8 -?s� >w����п����3sH?���4���q6�p=�=��1?KQX?��>������c��>nx�s�d��8�=�b���s���*��oO>�L?��b>��r>Ԛ3��s8��P�?����5{>�5?a���9�Hu���H�Fo޾��L>޾>s<��}�C&����~��h��y=>�:?��?L.��}4���uu��읾��Q>��\>^a=�ȫ=W�K>�e���ʽ��H��.=YO�=K�]>CM?��,>z��=d�>�����O�辨>�@>�.>{@?�$?���N��i�����-��;w>"��>�S�>kl>��J�䌭=���>Ѡb>{^�˯|��;�֨?�m;X>�����]�z�x��E{=ݮ�����=Η=9���I>��"=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ>p ���f�����|i����<��>2:?S���K������f�?"$?�l�5D����̿��x�J��>x��?0�?��g��'���<2�ͭ�>�S�?�f9?��y>����Ĥg�:��>��N?�P?�a�>J��v�P] ?���?	i�?\�>8̈?'�?���>;�����X�E7��.wf�^�����>�L�>�߼���ʓQ�~&���ŕ�JYw�L��Y��=鉤<9�>�Y�'����!>����UG^���|�[>Y�<�k����<>=��>7��>G��>R�=
9�����f��B�K?}��?����+n�=��<?O�=�^�F?�R4?�^���Ͼ��>>�\?D��?;[?	~�>��S-���޿�ot��@�<ogK>��>en�>f=���JK>��Ծ�8D�j�>Կ�>9��<1ھ�M��:?�� A�>�Y!?؆�>(o�=��?(�!?ɲ�>ɑ�>��M�� ��T�R���>v �>�!?I1~? ?:��Z�;�����v��%�X�v�E>�m?i?�d�>�B���V���ٸ�-��7��ߢ}?݋N?�J�dW?y?��=?:�L?y8>1/��+뾡B��{{>\�!?��,�A��J&��
�,?O?8��>P����սPpּ���R|��{�?�'\?OA&?���*a�� þ	'�<A0#��V���;m	D�7�>�>`������=\�>g�=�Rm�MA6�Vug<�s�=���>��=�27�3{���4,?�D�"郾Ϩ�=��r��wD�>�>�"L>����^?�=���{�G
���}���8U����?U��?�o�?Dk��ˤh��=?�'�?�?p*�>�a��nv޾`��w��x�a���>���>�Ah� ��܂��*���E��e�ƽ��,����>C��>�R?�>?��]>4�>�ꗾ��(�A���!���V^������7�'�/�=���q���J���x��^���`��5ڊ>�Q����>˒?|�>ii�>���>�>=yޮ>�QF>~u>��>z!c>_mX>��8>>��<%���NR?����'�"��t����4B?@qd?�I�>$�h��������Z�?���?r�?~Fv>loh�5 +�_q?�2�>�!���i
?;=���P�<F����������ָ�>��ֽ�#:��M�?f��h
?Q&?Z��]�̾vW׽jn��f|=�ˆ?�4.?m:,��U��t���W���L�9؃<o/`�NY����#�ۯu�d���]���Lˁ��G%�uw=8�'?䖉?�#�,y�aK��d�h���@�`kp>8��>D�>�Q�>��>>;U	���0�vN^�SQ*�gP���8�>k�w?E��>��D?.�4?�`?P�H?�w�>��>�hb�O?�"��h�>���>�G?�A?,s6?��?��?
�?>^;�$��q���־.?N~9?�`�>Y ?���>�7Ӿ���=�2+>d�|�j_�����)��=�+>�	��K@$��Mǽ��=[?����8�e����k>׀7?{�>3��>k���7����<9�>a�
?{I�>�����vr�P^�[�>Ϡ�?N�o=��)>�=����̺�k�=�¼�ΐ=|���R;�W]<r��=��=4u�곐����:a�;\G�<�5�>�?Q�>��>B����I�����%�=�Y>19Y>�N>�RؾXQ��f����g���u>�(�?8$�?�kd=��=���=������D\��ͽ�$��<��?�k"?�S?&��?��<??#?K>�q�EA��AI��%ޢ���?t!,?��>�����ʾ��։3�ם?e[?�<a����;)�ې¾�Խ��>�[/�h/~����4D��ꅻ���b��7��??A�X�6��x�ڿ���[��v�C?"�>Y�>�>O�)�y�g�n%��1;>��>eR?�W�>��O?��z?8�[?B�S>�Q7������p��֍��A>�??�I�?���?��x?��>��>%�*���߾���16�N������)�I=u!V>�L�>z��>�#�>x)�=��̽D����16��²=z�k>�S�>��>���>D�{>�<LH?���>�u��à��A�����<�Cv?v��?��*?�v=Y~�1E������>�_�?o�?6*?�T�H0�=GҼ褷���q��<�>2�>��>��=��C=�]>�~�>_B�>���_���)8�saK�p�?��E?���=(ɿ:~w��E�������0d������Z���)�~�־�>�"�ږ�]c�F�S�a���*�c������1{���%�>q��<2.�=#A>�.>3g���=LjP=�{�M��=���=���=L�㞀���ӽTj��cŻ��<�;�ַʾ�m}?�'I?7�+?sC?*#z>��>�9�㽗>$M��\�?GU>e�Q�Ж��;�������s�ؾ�
ؾ�?d�?����>}�B���>5�4>��=x�<|��=�Tf=��=;$�=��=g^�=?��=��=�>~>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�47>(�>��R���1�y�\���b��tZ�j�!?�H;��4̾�F�>~��=/I߾v�ƾ~/=��6>�a=^���Q\�Cƙ=9Z{�8�;=зl=	��><�C>q�=�#��2Z�=J=N�=��O>�ј���7��c,�D�3=���=��b>��%>���>\U?�[.?1�_?���>��k���˾Һ��zA�>���=�'�>y�=9e>^�>�{5?�A?c�G?ԫ�>�j,=<~�>�>��*��(q������}	==$p�?Ƀ�?戵>]m�<R�!��.�]�/�{Ѡ�S?��5?|�?��>�0�h��I/��1���O�� f��z�<��v��Ƚ+��!�������=g��>l�>s�>B��>�O,>��J>n��>��>��=R��=T=�<���<���&=���+ Y=��1<G|�����.l��3ɻ�������5\)�ɜh����=���>A>���>��=���^/>Z���x�L����=xZ���"B��/d�AR~�K	/�)a6�t�B>IsX>����4����?6Z>��?>n��?�-u?��>�8��վ0N���e�ʀS��N�=.�>r�<��l;��V`���M�$�Ҿ��>v��>E��>�tA>��6�*�>��}<b��3�0��>�ȫ�U޺��>$�O+���w���G��-[L����=F�L?Y����>�=`׊?��Z?"�?䔣>����ޡ�Fh>B������=8���y���gL;kG?��&?���>í����M�6Q̾�*��nַ>��H���O�����	�0�Y��䷾�W�>bݪ���о+03�c�������B��q�b�>x�O?��?�b�Q���XO����р���w?�g?i'�>�Y?�^?00���a��K����=i�n?s��?�4�?��
>�L=A;�.�>)�?I��?Q�?�Ai?i/��c�>�%���B>���A6��5�=�!�; �=S?�7?'�?�م�oj����	�ڛj�Gu���>�(�>�Y�>�N�>!a�>R�=��=��>���>_�>���>*J�>�0G>�ֱ��X.��0?Z��<�S�>:,?Nմ>���<`�i������G>z��E�����潤�R��|n=#
�>$ʒ>3�G=F��>lƿ�Ӧ?�-μ�St��G�>�=���Y��9v�>��6>/��<y6�>t_�>�l>e��>+��>�	�=�>J��=���j>[���i3��I��z<�9���j3>x5޾�dX��!�c��ʹ�v���� ��_[������_�ӊ��_�?fc=5�L�y>��4�h�?�}�>�?DY��ݗ��C����>4�>J���d��|�����Un�?�� @<7c>Y�>k�W?��?��1��3�itZ��u��(A��e�ݺ`�l፿E����
���n�_?	�x?�yA?dc�<�8z>桀?��%��ԏ�/(�>�/�%;�e<=�+�> &����`�ˮӾw�þb3��JF>͖o?�%�?�Y?gWV�_7N=�C>�,:?�N\?twn?�4P?	�C?M����@?���>�>�>��?2�/?�'>?�e?��>���=�����p/�0�ٽ�x���u�S�!�(p-;��=��=��=�8ƽ��%=Y�N=�[A��J��;Ԇ;T�;x>��ҥ=���=��>iɦ>�]?B�>��>��7?2���p8�S���R3/?ǎ9=����L������e�]�>��j?���??XZ?�4d>��A��C�)>�c�>ɕ&>�@\>/l�>]��J�E�tb�=�i>�=>��=��L�����غ	�������<�>���>]-|>}��:�'>�z��/+z��d>��Q��ʺ���S�Q�G���1��v��Z�>=�K?��?5��=�]� +��If��/)?(^<?�NM?��?��=X�۾��9���J�z<���>�d�<�������#��Z�:��+�:��s>�1���g��2LO>"V�$�߾�k��sB�ưվ��[=����B=ޡ��<��Ԁ���=�}>��t �sF��c4��SwJ?�[�=F��<�o��F���!>���>V�>�Ǎ��Ø�	�>�������=÷�>_�4>������[J�c@�1��>;<?�kX?�%�?0�\�c�d�:4>��kﾑ��O_*�F�?lH�>9 ?C�}>kz�=����?�	�-�\���F�v��>���>"���uM�����3����}�?��>�?�C�=��>�A?��?̩e?�1?�
?��f>o/��0L����2?Bc�?Ѿ";2b;�+ D���E�h�=���;?֊C?H!���G�>���>���>ʺG?d�s?ن'?-�;>߫��DR����>�r�>��e����P��=wf
?e�i>�y?�M�?%�h>�=*�&��,Y��r��=>�Y.?�]5?��?=z�>�`A?�����0>��7?�a{?���?G�%?���>T�?tU�>��?�b+>0Ў>��?�+ ?��G?���?Y?�{>�f=;�<����>�=x =��<@���/^>�u>�q:�T���a4=�� >ၽ��8�FOԽ��=�=s��_�>n�s>�	����0>_�ľhO����@>�y���O��U܊���:�[޷={��>,�?���>�W#�ܳ�=���>fH�>���6(?k�??{;!;<�b�2�ھ��K���>,B?���=��l�,����u��h=��m?a�^?8�W��'��-�b?<�]?iX��=�+�þ��b����f�O?��
?��G�!�>��~?��q?I��>N�e�<-n����>b�C�j�w��=�v�>�Z���d�r+�>)�7?K�>c>};�=�۾O�w�*p���?��?
�?7��?.*>6�n�%-��(�����V `?���>s՝�iQ?�ɻ�Ҿ_����3��Z}޾�����G��U݌�6��|{���4��<�=/O?dr?Z�q?��b?����0e��r`����'�U��d�����C�`�F��.D�7�p�����=������ֆ=`����X�FĶ?q��>�F.<��>��{��󨘾d��=|�������<�=3��=N�X=�v>G�>��,L�㭳�.�?V �>�w�>��P?V�c���O��D�?��c�b>�h�>s�>�T�>us3����=�nV�rKV�`w�一>&%Z?��L?�~k?*�D��8D��쇿�n+�/G*�2HT�d�R>�H2>�]�=
)^�����a`��,D��Mm�g���y��Y7����-�?�f�>ӛ�>���?���>e�ʾSH��[���*��]=R1�>%�f?@	?�ِ>:�:��B��>y�k?R:�>D��>ď��"��}���׽��>G�>�� ?��y>i�3��]�Nߎ����O�8�D�=ݗf?p̂��k^��ǅ>:�Q?R�q�?�<v/�>
�]��!�8~�!��+>��?�y�=(�@>��þ�3���z��L��J#;?�84?L���>q.��=�>��?��>ɝ�>���?�s=����'0�=Ӳ?4 Y?��Q?�V?+?��=�:�o̽:�@��>fr�>4'�>��!>�{5>��f��s��%☾�Dk>�Bz>鯈=�t~��Ĉ=��$�֨���F=&}`>�ۿHTU��>�N���������T�N2��gf���V���վ��Ѿ��[���u��J����b� z��#�a��O�?��?����������,\�L�Ծ��>����|*���þ��I�����"̾ʃ��e!��Oh�-4��`�_��P�>@
���Pο�������gxA?�57?V)?+HB����{i���=:�>��S��9�F&��-�Ŀh+𾂕�?u:�>��׾1�<��V�>�(\>����fW>��������VP=�R�>qeA?"�1?�f?��!��嫿sW���?ہ@�A?��(�G�쾉�X=H��>Ҙ	?�?>U�0���6İ��P�>�1�?|��?HN=)�W�����e?!K<��F�#߻h�=g�=ܭ=<��P~J>jh�>���AA�+�۽Cu4>*��>��"��5��M^��L�<��]>j�Խz䔽5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=u6�����{���&V�}��=[��>c�>,������O��I��U��=�i��[Կ�I.�K�	�������o�߾>'EY�,�x��=QU��B�Ͼ�5�i��<X8	>�>�v�>#+>eCU>�AW?)s?4,�>�N̻�Z2<����$������
۾IԾ!��bz��D6¾e
þ��۾�	����=��O������?�&�X=¹R��ҏ�.� ��u^��t>�Yl-?��>l�̾�P��y���!̾���(?�����ݽ̾��5�Ԙk��@�?��D?�_���\Y�}���҇�6���q�S?��se�``��_��=Z���oW=���>�=�����7�E�Q��O5?�y'?4������#WU>���;�<�^4?Z��>�lý��>�@+?� 꽵>t�,��>X�c>��>�{�>	.�=F)�����4!?�#c?v�ʽ����y��>���?$���jv=�HB>���dN��JC>�K={��D[�I����<-)W?Y��>y�)����]����AN==Ӳx?�?k'�>vyk?��B?��<�b��l�S��F�w=J�W?�%i?��>j���Aо1~��J�5?�e?��N>�nh�w����.�eQ�&?��n?�]?({���t}������xn6?��v?s^�vs�����;�V�i=�>�[�>���>��9��k�>�>?�#��G������wY4�$Þ?��@���?��;< �T��=�;?h\�>�O��>ƾ�z������+�q=�"�>���ev�����Q,�e�8?ܠ�?���>���������=�թ��3�?��t?�ߜ��V.�����zy��hϾA!�;_ 2>z�
>��p���x5;��x��A����1��S��>�@ϗ�~%?(��$�ǿ..߿�	����b�D<̔ ?���>��x��Cz����M�K�� \�7aP�hc�>j>/I��gN����z���:�mT�� ��>����G�>��R�-������ڜc<�T�>���>���>؋���<��}��?Dc��*
ο����9��6X?�1�?���?�6?��<F�w�a�{���� �G?��s?� Z?J{-��^�NL7���T?K4���s��y6�K��u9>�*;?z�>�@�%�;5Й��?���> 9=��ɿ�7��g��zۗ?��?�����>���?l�4?U!��������C��";'D(?���=m��!H���I�vԂ�P?$� ?/Y�����_?��a���p���-�2�ƽ�ۡ>�0��d\�H��+���We�����?y����?�]�?�?^��� #��5%?l�>]���B9Ǿ���<M�>�'�>j*N>�7_���u>#	���:�
h	>Q��?�~�?�j?b��������S>q�}?a$�>��?p�=	b�>c�=��X-��j#>}"�=��>��?��M?tK�>�V�=F�8�d/�E[F��GR�n$� �C���>?�a?��L?�Kb> ��O2��!��tͽQc1��T鼰W@���,�S�߽�(5>J�=>W>��D��Ӿq�?�o�?�ؿ�i��Ur'�+54?��>�?�����t�k;��;_?�}�>l7�<,��&��*G�֙�?H�?��?��׾a*̼�>��>yF�>� սf���၇���7>��B?z�6D����o���>A��?��@�ծ?�i��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?�Qo���j�B>��?"������L��f?�
@u@a�^?*��տ��3ξ�D���?��>Xh�H�F>Z�\�� >n|r>{�j<j2��c3>Խ�>��>�^�>��>"@t>��=ku��ӎ!�vH��ӆ���;f��:A�
��=�t�*���20<}%�z�����޾A �ߕ��1��*0(�<�.�o�=���=�
E?{�K?��o?QZ�>�:��h�=�4�ǵ�=3���T'�=�t�>�?��E?�+(?��=}��	�c������{��O͎�9�>�_]>���>���>���>:�~�G>��#>m�n>��=�H=9fݼ`�#< >=�>-�>�.�>��=�2�=1��	v����e���"��q=�y�?��ʾ-G�� ���־�����=u�%?�k>��5+ֿ�� NK?-0,�Yn�򣁾�R�=Y�8?6�L?&,�=cr̾��2��f>��ҽ1f+�PZ=2}7��z���9���>1 ?�|f>�t>�3�Bj8���P��Z����|>�-6?���#Y9���u���H��`ݾG5M>߿�>�-C�q�J����>i���|=Qm:?�o?UY������=�u��O��q+R>�>\>P=e��=mM>�-d�L,ǽ�@H��}-=���==�^>I7?�)>���=�>�>i����L��ۧ>��?>µ->�@?:�$?�	��қ��M���=+���v>�"�>�.�>o�> PI�O[�=M�>Ża>Ό��~}�]���>=���V>���"8_���|��7=�W�����=�ݐ=��I!9��#=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾUd�>fp�g\�����F�u��#=w��>�1H?(a����O�">�t
?�?ob�D����ȿ�~v� ��>U	�?	�?��m��=���@�)s�>Л�?�cY?I`i>�d۾>RZ���>0�@?�	R?��>�9��'���?�޶?Y��?R�E>�x?���??�-۾.�`�m��AR��lB9��:�>�R?A6 ?u�*��k�\p��/l�2U�6���	i=���=d�>�tM���m�We;r���3F����<�7>��>0Q�=X��<��>N�>� �>;��=j�q�Ja�$0L?�я?����m�g��<P��=_��(?��4?3W�ξ�(�>�[\?H��?�d[?ð�>ڽ�Kۚ�v������sT�<5L>S��>&N�>���.L>�վE�E�ύ�>�6�>l ���Rپ�����ǻ[ܜ>�!?���>Y��=�� ?#?�j>�,�>�bE�#:����E�6��>���>�J?��~?��?$ڹ�I[3�����塿�[�d7N>	�x?�T?�ɕ>ߎ�������OE�CI�,������?Arg?HO�K?�/�?L�??��A?+-f>e��
ؾ������>N�!?e���A�5(&��}�z{?&5?���>�����pֽO?ռ��tJ���#?y&\?b8&?ۄ��a��þ��<����Wo���;�J��T>�>t���K��=�A>���=�Um�K�5�w�p<�h�=c��>���=3[7�r��0=,?��G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>$�l���K���ڙ���F��_�ŽwM��W��>�>X`�>ya�>$�[>��>֗7��!���C�ɾ47]�X
�	33�`6?�H�R�����L�=��>漯����c�>���5N�>_��>��">�W�>�{�>��>v�
?�\�>''�>n��>� �>Ż�>��>�E=�J�aHR?����ϲ'���U����-B?jdd?%3�>��h�ˉ�����]s?���?Ux�?�`v>cjh��#+�ea?��>����t
?]�9=���mo�<�o������Y��ū�Z}�>�e׽�:��M�^9f��u
?�4?�:���̾7a׽�\��M|=S�?Pd)?��*�G�R��qq���Y�mP��K�+Z�2��Pw&�p�n�(̏�R����S���g%�UE=h�)?rn�?1����I����g�Z?C��g^>A?�>��>�b�>2�P>�
���4�;�[�w.(��Ѕ����>j�z?�
�>V�@?0;8?�(Q?��K?겒>р�>4����>�H=#��>m��>��,?q6*?�/?�i?�r,?�^K>���"8����׾�4?�`?[�?��?��?���/ý��B� ���oe�FB(=���;�F��`���@=�=X#O>&?���$9��=��}'j>�u7?f��>A��>���R/��ŀ�<=��>�c?�L�>� �Q�r�a����>���?����5=��*>u`�=����� ��~��="Ƽ.{�=�}��B���=<���=��=;���b��D��:}��;��<�t�>!�?ߔ�>aD�>dA���� ���s_�=6Y>�S>�>�Cپ�}���$��k�g�	\y>Nw�?�z�?o�f=��=���=�|���T������������<ݣ?�I#?_XT?F��?(�=?�i#?t�>v*�:M���^��\��ɮ?!)?|3�>����Ͼ6�����.�%�?Wp�>SId�NU�ϯ/�������m�M��=��5�����6��r�?��0T=P���z�����?B�?����;�&o�!I������%�??���>���>��>[,��d�����7>j��>ȭN?|��>��5?-n?�W?6�.><�3�"lL����5=%D�>rM0?�Jt?^?��g?Q��>�[6>�������*�<ွ(H�[����U�=��>	��>��?U��>�V>�;M��>½-�]��ʻ=�y>���>9�>g=?}hq>� =~�O?y?�Ѿ�I�:������E��K��?_P�?K{?�#�<�r�_'8�ؠ�����>
E�?�;�?Ś?@�����=�<�����Ql�J'�>��>蠰>�Z�p���7>ݰ�>V�>I�Z�����M���ۼ��?�B?�c!>�ſ��q��p�آ����h<qВ���d��g����Z�H�=���@���۩���[�3���fY��I�������`�{����>�q�=��=���=9�<>Ǽq��<�#J=)�<��=K1p��g<t�8���׻zf��dJ(���Z<�J=�����/ž��u?�F?��.?D�F?:ă>�l>�~��˚>�VT�B?ScM>u��l�����3�<ݦ�(���iCվnpݾq_�[��	�>>78��>}�5>�n>2�<��=}�=m�=�#1��GF=ͨ�=R�=��=���=�%">Ɲ>�6w?X�������4Q��Z罥�:?�8�>f{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=J����=2>s��=v�2�T��>��J>���K��C����4�?��@��??�ዿТϿ7a/>�Y7>�>p�R�wm1�]i\��Zb��|Z��!?	1;�u8̾�@�>���=�߾��ƾW�-=|�5>Ǆb=���3\���=B�{�Z<=1^k=c�>�D>�^�=u���ζ=z�J=S��=�$P>���C7��P*�4�5=U��=��b>4&>W��>�A
?Q?"?\\P? X�>�Q��������`�>�����>6�5=/V>�8?r,??�[B?�$7?�H�>)�¼�\�>5�>�P3�z�y�'� �\�⾋kZ�*��?J��?�nv>`��&�Ȫ��%�ݹk=��?�?ܙ�>0b>{�2��i�&�>�,������s�J=.�m�?�>�#�w�F�����B�=�>R��>�ɡ>p�>e;>�N>bk�>�>���<Ŕx=[�;��<W
���τ=�"ļ��}<�����+���^�
�4�hvѼ��; A����HRP<���=:��>#<>���>Ԓ�=���~B/>繖�|�L�Y��=H���+B�
4d�:I~�$/��Y6�^�B>?;X>�z���3����?(�Y>m?>G��?wAu?!�>#���վlQ���=e�>[S���=�>	�<��z;��X`�n�M��}Ҿ݀�>���>�=*>��(>98(���4����=�;���N��	�>Z��ߜ�t��=r���ˬ�᳥�:y�>r�=�m?(`��ԩ�=菙?C�@?��?�,�>Z:@�}�����[>����ִ�>�LK���6��<֧$?�
?~��>�َ���u��I̾����޷>�AI�3�O�����?�0����ͷ�N��>������о�#3�Lg�������B��Mr�#��>��O?W�?�;b��V���TO����()��q?�zg?��>L?PB?����s�o��$��=��n?��?$<�?q>�@Z>Y���\�>�f?y6�?2?��_?����?/_�=8YA>�.��� =��T>�1d>JKe>n�?JY?�~�>��r��T
� ��V>Ծ�oٽJ�	>s>t��>>��>���>u��=��=�x�<��>YK�>��>_v>���>/ �>.Kž�O�-O'?������> ?H�>��"<]�x��7��y;`=�`�����<���<X����W(=&�=�Tf>8��=t�>�X¿�?vi=��P���>K���p����>naH>X�B��O�>v<>=��>�p�>�]*?)�R>b��>��h1����>�="�<D��TJ�`)��J^��7U5>w�����O�sc)�9:��f.:�"�Ӿ����q�Q�c׆�|ps�8��=��?��=�	d�0.6�T½|�?#�>�?3
t�Q璼8��=��?�{�>eJ
�[���ć���Z�'��?c��?�;c>?�>�W?7�??�1�3��uZ��u��'A��e��`�R፿������
������_?��x?�xA?�G�<�9z>"��?��%�2ӏ��)�>r/�d&;�BC<=++�>�*���`���Ӿ�þ�7�sHF>$�o?%�?~Y? TV���O�2D>�8?��5?:w?�I3?t�4?�)�%?`�<>̴?��?�)?L�'?�%?C+(>�U>D���><g��5k������������û��N=)�=��;��)��;�u#=�~�'z�D�f:���<<�[:=���=к�=�B�>��Y?�.�>fl�>�8?�"�p�7���H�/?N�X=*��-ᇾ>��)��3>o�h?�׫?��W?}U>s�@�T�B�S�>K�>�/>��c>l�>�:�� <I���m=p�>>{
�=Ғ[��Ă�i^	��H��y=��>���>4�{>F���2(>N.����y��"d>`eR������FS��G���1�:�v��C�>t�K?\�?b�=c�W%���,f�q)?�C<?dFM?��?�P�=�B۾(�9�B�J���k�>��<����������:��b�:�\t>��S���h^>O��vc�.�l�ӨI�2龄vG=���M%T=�$��Ӿ:'��V��=V
>3����C!�����T���׀J?/+p=˓��ӀT�-����>�8�>q5�>�9����i�@������{�=���>��4>�#���P�{_F��<�]�>�8Y? V?5Rt?c��sf��EM9�xJ���Wg��f��S?4D�>њ?k�d>��.>�R���z)�u�i��B;��	?�j�>O�S�(qa�A"�Rz"�b�K� r�>�?ٳ�=,�?�<�?�
G?�pQ?K�J?] ?j�$>w�Y翾,�5?FT�?�ｼ�~��"����xe�ĨD�:�2?��G?����߄�>�a?&o?Xn=?h�?�U?¶��Z"���D��ɉ>'��>�)l�p���%�N>r3?NT�>��?ڞ�?48|>��F�ޢL��J�=�G.>��>��O?�s:?�?1.�>�)�>�0��	6�=eJ�>�;Z?�q�?_Tx?�-�=!��>��a>	/�>�)a=�M�>���>q�?�.C?�`?�b8?7\?S�i<B����̶�L>ý���S�XHߺ�p=M�l<Z\���x��h��5<W憼��L��2���偽C�A����A�>��r>����V�0>��ľb>���mB>몖��B���Ɋ���8�ב�=9��>�?��>�m"�/O�=��>V��>����I(?�?G�?�K���b��ھ��I��-�>�B?>�=��l��C��au�ŏh=G�m?�Y^?X�W�����F�b?��^?����<�_Ⱦ��l�/\�$�O?n�
?�JI����>��?,s?���>z^���k����2�b��o�a��=t�>@
�~=g�c��>��5?���>��m>��=�ܾrkv�����'[?�K�?���?�D�?k+>__n��8߿*�پ����ɮU?ɰ>-���",?G��=�4����Ͼ�M�f�6��������&�$���rA���;�JT���,>gG�>4�?,�m?g�O?�x���{_�"�t��m|�<*S���Y<���}2��wB���8���l�s$��V�s����3e��q~���@�mi�?8�'?ź0����>�ؗ����̾!@>j���^����=e��u�@=��X=�\i���/�� ��g�?�~�>EW�>{<?P�[�@>�o2�Ѳ7�Q���3>T��>s�>Ë�>�j���+�B�뽣ʾ�=��QDҽ�ib>>/^?�`?_pn?�5��;�;�SW�_+����^�j���b>=��=��S>������)�5��N7��x���c����~�6;�b?���>���>[d�?�?? @t�/�ݾ�^��k�m��..>\�?��|?.�?/�p>�Q�6�,��E�>1�l?d��>K��>Aጾ��!��{���ֽ��>|�>J ?ogs>�/�܇[��i�������<9��U�=�-h?
���z\b����>$�R?{�w;B�0<���>Ss��� �`���'��>}H?���=��:>R�ľ�?��z�B����)?��?�����*�"Lu>pO ?�>�1�>|�?���>g�����j���?��^?�!J?A?�h�>9� =?ާ��Ž�!���)=cY�>@dR>_�Y=��=KM�\�W��"��D=t��=��Լ8~����<����o<\��<�4>��<
S��M�x6�*¾���Α���Ū���-��oP�¬�!���݁�+5ؽ2h?<r!���U�TĖ��3��_��?E��?�������5���W�� c�O��>9,���罝|�C`�1<ξ�����龅B�~�`���s�x�z�;�'?������ǿ���b:ܾ\! ?�@ ?�y?+�z�"�T�8�ܯ >�E�<R<��}��ᚚ���οǦ��x�^?
��> ��<��	��>��>��X>�Cq>���4鞾%0�<�?І-?2��>Òr��ɿM����̤<:��?o�@]{A?�(����~V=p��>��	?��?>�I1��I����V�>;�?<��?�yM=��W��	��~e?j�<q�F�A�ݻj�=�N�=5=|��3�J>vR�>_��>SA�YDܽ8�4>Iׅ>��"����w^�0��<�}]>��ս�8��5Մ?&{\��f���/��T���T>��T?+�>k:�=��,?W7H�_}Ͽ�\��*a?�0�?���?#�(?8ۿ��ؚ>��ܾ��M?aD6?���>�d&��t���=�6�񊤻y���&V�`��=Q��>`�>ʂ,�����O��I��P��= �~�ȿy�'�D@"�	6�=K�=���LS�U�/��둽�`����|�]R�J��=�)>l�k>|&�>��J>��H>lb?P(q?��>�H&=����i��!�㾛��<K�C���N���	����া>9��K�����yG��������V�,4=?�N�*��Q�
�|Eg�PS��@#?ϵ>U�ؾ�D���We=N� �yA��Җ�:��U�G�����-�DD���-�?hPE?&7r�U�4�=� ��v�_轳CE?�i�=�Sh�#">��������� >��h�����/�'�G�Mq0?�]?�?��i���;�(>���=Y�+?o�?��a<��>g%?Q�)���^\>�W4> ȣ>�n�>QE	>���y�ڽ�?�1T?�g�����[�>M'��I�z���a=�G>��5��=�.�[>@�<_e1Q�ᏽ`�<�(W?a��>��)���a�����PZ==��x?��?.�>i{k?��B?l֤<�g��e�S���Vbw=��W?1*i?��>�����	о����"�5?ȣe?��N>�bh����%�.�SU��$?�n?1_?#~��w}�t��j���n6?��?�:O�M������J派�?�H�=O?�7��4����?����"�޿j%���|?�r @�l@F&�=V�~�2��>��?VӮ>����bӾ�ג>�$��A�����>ZD����\�������-.�>���?�dD?Q}��Q�5���s=��B����?)�m?PI�����=�Y���b�!!�u��A>�ݼm1	�~���_E�k�M�S����x���1>Ph@�����>�tD��mӿ{rտ�-���a��m��
�>�u>1�u=	Zo��5u�j��I�a�6P�-j��$�>{ >�œ�����u|�q4<����
3�>�� ��-�>apQ�|����	���{X<�ݓ>���>z�>���������?�_����ο��������W?(��?2Ņ?�H ?0�<�:v�L�u�0����G?*_t?�^[?%0"��b^��V;���j?c��y[`�*�4��KE��0U>A3?sG�>�-�r|=g>�y�>hH>"//�k�Ŀ�ն�E���f��?���?�u���>��?o+?�q��5��IE����*�k�@��8A?�2>R�����!�h9=�cҒ��
?��0?W��3�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?! �>��?�h�=\d�>X��=��^_'�J�#>s,�=jU?�U�?��M?U2�>Y�=�p8�M/�?AF��<R��*���C��ɇ>��a?��L?/�b>N*��D
1�GB!�U@ν�P1�w6�e*@�C�-�j�߽��4>C�=>�*>uE�0�Ҿ!�3?X ���޿'������c�6?�4=��?Y�߾�����+���L?=u>��)�R��曑�<��cP�?G�?��"?ȷ��(�q��E�>~K�>y�w>�z��S�����i�0>��f?ʮ��}򗿨�e�Kf�>B�?5�
@w��?�)i��E&?F��`��x�h�@���䏷��酽��;?o'׾��1>�>�3��ă�٪��)g����>�~�?�T�?(,?�ff?wlj�"�+���(>ĉ�>}c?'�?G>;�J����=K
?+�!�C󏿼��[1a?!�@��@~�j?���!gֿ"����L��薺�$��=���=��2>��ٽ�[�=%�7=�8��4�����=��>��d>$q>�(O>�a;>;�)> ��$�!�7q��ȣ��S�C�K��~�g�Z�&���Rv�>y�&4��n����6���1ý�r���Q�w3&��=`�v��=�7L?��d?�U_?�g�>�W�?R|>ϾC�k=�w����=@��=� ?��H?Y�?���=ߙ��g��rl�õ��m��%�x>�	(>-�>��>B}�>M1����>�Kj>T�]>#�&>j\�=e�r�de�=apE>4e>̽>+M�>o>�u>�岿$㴿^�c�5]���[�r��?��e��vH�㚿�#}��{ɾ�X�=�))?��>Ґ�\�ɿ����2cG?f���n
������!>�1?�[P?�� >_��fr&���=�~�0�Z�̇�=M� �pri��\ ���>i@?v�C>�ln>��4�u�=���K��
���Y>��4?;s��\/@�~�ՒA���ן@>�>�H�T�L����6��Z�`�zm�<�9?�'?�p������e������d>L�X>)��<ܤ�=��^>򉏽�ýj�F��eD=Q�>��P>�'?_Z>;D�=䲒>���$�W��m�>�b>7�>`7?O$?���
�J��kS�n,	�Y�>y��>'�>y9#>X�;�o�=It�>�>����Oν�����f>x�����P��	����P=��?����=t�=��ɽ��?���?=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�E�>�n�ģ��]��DOU�b*>HY.>)*K?������_:���?Wn�>�5	�04����οK)��L��>�/�?''�?��Z�����x?z@�?��?jI�>8T�(�x�?^# ?1J#?1��=z��zR��'%?k��?OΠ?z��=�p�?��?���>Mި��K7�����⣥�(է�!b>F&�>��>jb��t�����<���-��C�aY4>�,b=��@>]�d����렮=�]Z�����,�>���>�׎>���>�i�>N��>`�>��=ӂ�<��{�g0�y�T?�;�?���@���0br�s��՞m��S?��d?:n�=y8þ���>�~�?؊�?�f�?��	?�����f���f��;�Ⱦ��'���>^�?�_�>8���Si>�bξ
���빚>�V>� ��4;'��t���2!�r�=��
?�� ?��W=�� ?��#?z�j>5(�>8bE�:��R�E�ư�>���>^H?��~?k�?(ҹ�Y3����T桿��[��4N>��x?_V?�ɕ>����񃝿�E�{SI�/���H��?ug?�U�s?�2�?N�??ߥA?�/f>�}��ؾ㬭�G�>�s!?A��%?���%����/�?��?	b�>M̐�gн׬��P�t��>�?�[?Z�%?���^��E����<%9T��)��)��B�ּ?M>�>Vy��z�=�">��=��o�65�c�<�;�=���>"��=?�7�㈽�p7?��2=Є��~k�=1t��//���e>�"�=" ۾�g?��� w��BM��W��� �?���?�>�?x
�aǂ�M�:?p��?���>�L"?�Ҿ��@��������n�<rh���^>���>Xz�>���e���ݦ�Wə��R��M�<�#U�>^�?>kZ?�C0?դ�>�i�>�o�`R<�g8���|�O.g�*h���(��"L�͵�����l,��*'�;���㆒�yR�>�1����>���>\z�>(k�>�*�>�<2���>�8>'��=���>�t�>��h>Yr>��;\N.<=R?N���Ţ'���辗����B?cqd?�B�>�wi�\���ۨ��q?�{�?*k�?0~v>#Yh��+��d?kD�>����~
?�:=o�����<z��^j�9���Hf��̎>��ֽ#:���L��e�p\
?�,?�ˋ�+�̾x׽�3��kD�=v��?$�%?�&�{	K��co�РY�ZmU�&i�U�U�6��e�!��m�-퐿X���pe��(K'����<��#?�H�?	� �6U�e���b�p��KD�
�D>��>̷�>!�>U%>l�ϼ(�g�^���,��&��[x�>��t?���>&�M?�MB?=�M?D�7?�vN>�g�>����.��>��f��,�>f�>_u.?�/?�_3?{�?��?Ƀ>$94��	���依?l??P$?��?J�>�w߾.^���<��"��Y��}�R;<�Cȼe`̽��>�Z÷:��a>s>?G����7�Ϛ��\g>F�6?Z�>��>-������9��<�X�>,�
?'&�>8��#Tq������>+��?]����=��(>�B�=q�������1%�=����5i�=�6Z�v9��"<��=ܩ�=v� ¥:��M;��W;OS�<�t�>5�?���>�C�>�@��-� �_��f�=�Y>BS>�>�Eپ�}���$��w�g��]y>�w�?�z�?߻f=��=��=}���U�����L�����<�?AJ#?'XT?^��?x�=?[j#?ӵ>+�hM���^�������?�!,?T��>j��ֵʾ��]�3�ʛ?�_?|6a�ر�:)�o�¾��ԽP�>�U/�0*~�V��<D�	���������j��?���?�A�I�6��p�n��� d����C?�#�>�R�>0�>D�)�t�g�'��0;>Ċ�>u	R?��>��O?�K{?��[?G
T>�8��)���ޙ�i>�$k">.,@?��?�Ȏ?G�x?���>�v>�*��Oྼ3���]����Ă�M&X=:Z>qs�>���>[�>�M�="oɽ㲽;�?���=^c>���>��>��>�Tw>`��<��G?��>�V��������C҃�˦<�ʠu?`��?	�+?�y=�z���E�n,��X�>Xm�?���?9-*?��S����=�0ּ$Զ�"�q�X�>�ɹ>b3�>1Γ=`�F=Ht>.�>��>�<�	Z�on8�hWM���?[F?s��=����Tuv�N��=Wؾ�BF>����Ⱦ������>X��<v�G�e�=�����虾w,���7����+�H�[��>��@�^�&>��,>�?G>��U>��8=�A��	9�Ea$>��S=1�=M�'���ǻ��κ����N�P�*��=R�ʾ��{?;�G?.#+?��C?�r>�>�D#��N�>Jtw���?��D>Z���6�=�nE���ő���ؾ_�վ�ye�⟾M�> fE�r�>�g0>Ԣ�=�r�< F�=�e=�$�=?J:O�=���=8�=���=*~�=O�>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�K5>�(>�R��h1�~(Z��{c�H�Y��x!?	D:���˾$�>���=&u߾�Bƾ�j*=)H6>ϼc=[L�$/\����=�;��ר?=~�n=<u�>�C>�C�=D����=s�K=�)�=9nO>6��>f9��(���6= e�=1�b>�h&>�,�>��?;/?[_b?cJ�>��m��yȾ.y�����>6V�=��>� �=�oE>Q��>8?�\C?A�J?��>G��=��>�;�><+��o�Z��<������<| �?�Յ?��>�zw<D�Ƃ��:�����XA?��0?��?M_�>����a�5�"�W*@���<���=���<��Y��2�u�N��~��0�o=w�>/��>ڮ>v9�>��+>e8w>���>kG>�q�=N2�=��<5�=NZ�;�5�<W=_��."=�������d+�E�`�?G����<ޛ[��Q<���=�>�(�>$���>�e7>��l�R9>G���T`��^>�6T�t�V�=�G��Ɓ���X�~Y����>���>_�½4������>5�Q>��I>/��?�O�?�n>�.����쾥3������ ˽(��=���>�R�JR�	��J�\�������>��>��>��l>�,�]"?���w=� �*e5���>�j���[��7�t4q�E?�������i�Iߺ��D?�B���q�=�~?f�I?M�?��>ZA����ؾ�?0>�C���Z=���0q�R��R�?�'?���>���D�"̾�"��{��>E�I���O�����߿0��#�����s�>���s�оs3�&i�������B��~r�'�>��O?��?#Xb�M_���/O�v�����R?7xg?��>*L?�j?���������y��=��n?��?NL�?0h>���=%���l��>Ɔ?���?�?t}s?�~*�C��>i�<�LF>߿ݽ�}�=�>��=��=u�?��?1�
?2�ǽ=	�q�ܾ���Z�k�ۛ��T��=O�>��>8�c>Kӷ=$�9=��k=�\> ��>\	�>�i>�=�>4`�>����YB�)�>���=�y>��7?�0�>�JC>�88�?>I���>�W��~�Ƕ%�MT{�A�=��`>��">Ԥ=e��>̈́п�z�?:�=e�3���<?�ȴ����pA�=���������?f�L>���=�?�ƶ>������l>->�̾rQ=d��C�m'�׻*�v����B>�1�Գ_��8A���/���T��6��
t���g����U�5�%1���?q6%=�:����.��_��U?��I>W?A����c���I>b��>k��>����ԟ�蟚�F"�@��?P�@�;c>��>H�W?�?ڒ1�83��uZ�#�u�k(A�+e�O�`��፿�����
�s��)�_?�x?+yA?�R�<+:z>Q��?��%�]ӏ��)�>�/�&';��?<=s+�>*��&�`�x�Ӿ��þ�7��HF>��o?8%�?tY?6TV�����
�j���?8\Q?u�=?�:?G�t?M딾��J>�	?8��>$��>Ɗ1?5�B?�|?:A�>��>i��<���>�|ӽ�l��;P�%�ٽ�~c�Hn�9긼ӝ�=�����w��=e'�.�<���̒%��6�;�S=�>��=a��>Q�]?�.�>	��>��7?���e8�ܲ��/?5G:=ِ���*���٢�w
�
�>��j?H �?�^Z?smd>��A��%C��5>RM�>�E&>��[>2e�>�)��bE����=a3>R>Y��=zM��Á��	�c{��� �<~6>�G?�^�>��T<iu�=b�徊s很kc>�߱=�A<�b0�l[(�����1��h�>�m`?�?x10=O�ݾK��Mq�V�><�]?��s?dg|?��>�3B�B�W��q����{��>V���/.�V萿0��3~E���T=�@W>l���ߠ�$`b>����n޾�n��J�>���}M=z��V=e�� ־��d��=,0
>̦���� ����֪��0J?z�j=Ou���aU��s���>R��>�>C�:�g
w���@�=����K�=��>"�:>w����wG�!1���>_�E?��e?��?�ƾ�z���*���;�T�������?� v>r4?��=�wK>k<����'�n��Ki��?�Z�>2�2��0+���þ�q�z*��d�>iS?A=�`?��?�S?2@&?L�L?�[�>�2>����%?�z?<?c��?~V^�� ���T��w�7�͗��^5?g4?�Z� �S>�?�#B?�?M��?&:&?�v�<��	�[\V��+�> �]>fv����dK�> [h?Mk�>��b?t�x?%ס=G�L�AξĆ<}�>���={�?�s�>�{#?��>���>=�ʾŞ�>�?��?m��?#9�?�r�mBW>A�>Pe�>)j>�d%�l1?�?�_?�1�?:�?�2 ?B���������Ɣ���8��P۶=z}=�q3=�ؽyΙ���$�)�<M�Q��f��
OI=q����a=��=������>TBu>#����l/>��ľ����U(<>����ꚾj���<��=j��>o�?� �>�#��:�=u4�>Ԁ�>n7���'?�D?�?�}�;�b�",ھ��P�P��>�A?���=%�k������t���n=��m?i�]?�[�}���`�b?2�]?�j�8=���þa�b���龙�O?@�
?��G��>f�~?��q? ��>��e��.n�5���Ab��j�(ζ=�n�>9Y��d��C�>ɕ7?N�>��b>�)�=�}۾	�w�n��I?��?���?M��?*>��n��-�)_뾈*���X?5f�>��!��F:?�E ���Ӿ�by�闾⬾U��Ib�����;K��e���J����0=1�+>��?��?Y��?�'D?�+���n�[�B����Ysw�IXʾ�n�RsF��("�oE��d����:����ĳ�v%ʽhw~�dB�r�?0T'?��)�L0�>�ј�����ʾ[@=>}u��\:��F�=���tx>=�i=��h�F(�9뫾Lw?�o�>�W�>a�;?��Z�T>��~0�I(8�jI���'5>�F�>�P�>c��>��s�%1� ���
;Q����۽9u>*�o?�K?��T?Kii�;\D��u���7���>��[�^9>��E>}v>$�����#����v�z�I�7��ϗ�[��%NN=�G?�'�>�VO>8U�?_?��о�&���	��_��j�=���>��6?���>���>�R��?��m�>̈m?!��>�<�>rv���_!� }�8�սO*�>D�>֌?�t>�S+��B[��ێ���hL9�&��=�g?e΃�r}c��N�> $S?L\i;r`<&��>�r�G�������2�5�><0?色=K6>��þ�y	�� {�\{��'Q?En?��Ͼ�Q��d�=7�'?���>��?|&�?\��=�:�M�5>�X?�Y?��I?7�?&ȁ>A�=��6�T����E��2�U�Q>���>���= i8�*���ܙU�nU:=��)=��5>�4�v�[���B�/^0���h=��e=H*�>�����O�U*��E�-��7߾zI��Ǔ�{6����~],��d��O����{��a��ņ+<P���X�㽔͂���Y���?���?����P�߾$����v��j��f��>̧�p��;~e;�޽�M������ò�����=��L�ZX��N*?!���Rп^푿������C?X�>+�?�*������(�mB~>Á�=����(6�ڭ����Ͽ
;/��ـ?У?=F�?�?�|�?oS>�eA>��C>�{�^��jJ=#�1?�b?�h?����@�οI�ƿ=Ir�0�?�@�mA?�^(�(���[=��>��?��@>�p2�1��y��Q�>�E�?k�?�S=W�W����Ze?7��;h�F�٪�?#�=]�=��=֓��H>���>|2��iA��rڽ
�5>`j�>�. ��J���_���<�`>�ս�Ж�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=��������4*��;8��?&>=ݺ��ڽ�����[I>��*�^TܾIa��s�ҽ�&>?I\>A�>���>.�*>w>�	g?	�n?��L>��:S~:��x������h>$�><E��U��~DH��]ƾy������0������X��k୾��E�57�;�S���Xv	�~#Z�fI�W�/?T��>eʾ�c�豼<*5о�q��.B=6�������7/��]����?s�W?������J�g�����=I�7��Kk?�XE�N�Ӿ�R���X>
��Wμ>b>ݬ�.�"�a�+���7�{!@?MO?�۾F���B�=	����Փ�y4?E�?�0ϼ��W>��5?5(V�ǋ���#h>���=t�s>�X�>k;�=��ľ�Ͱ�Z�?�h?�!��P"ľq|@>w��M��K>=��=yc��|-��[>�H=W�P�1�`���<�G�0�T)W?_��>2�)��b��3���_==��x?.�?G*�>�xk?��B?H2�<�d���S���Qw=��W?�'i?�>X����о�����5?A�e?4�N>�eh�v��>�.�ST�Y$?��n?�]?����w}�Y�����o6?�v?s^�ns�������V�k;�>�Y�>���>:�9�k�>�>?Z#�QG��һ��Z4����?��@��?3C<<.8�n��=�<?�X�>1�O��Bƾ�m��k�����q=��>����ev����QX,�E�8?���?��>;���ת�'��=5N���i�?��v?��_�]I=�(�(�w�t ���J��n�=��;�'�_����L�X��r����c�U�����a>��@ӎx�=�>�鮾g��0�ĿL}�>����S���>��y>�Ep��Ծ�j���b��ρB��>g������ �>�K>�i�i�@�>R��:L�燿���?��z</�>�����]���:�� �3�>�]�>�Y>Ae �F��,�?���3�׿�����X��:V?B3�? �? _(?b0�������3�+�=/cT?x�{?�tS?k.����,�����v?��	���U��oa��d>�1�>O��>QG��%�="E�>�!>=M,>��k�,���ue������?Q��?*/�?f?��?.Q�>��7����Ze���U�y0Ѽ|?�B�=3��_�[��Lj���.�n�4?5�G?Zׄ�X8B��_?��a�*�p���-���ƽڡ>��0�#I\�����_���Xe�2���+y���?d^�?��?���n #��0%?��>О���;Ǿ�G�<!��>�/�>�+N>�K_���u>q�&�:��]	>ϭ�?�}�?�e?镏������`>�}?�5�>�	�?b�.=V/�>���=o
����㽻B&>�>���>;�]?O��>��
>����H�;?���R�N|	�0wM�f��>W�t?knZ?W�>S1G��=�g>����Z�j���ѽ�8)�$����3�>E>`>�c>�����q����+?a�;�9�ݿS�p�*����:?6�=M� ?z��i9g���=7�A?>m�>���� ���6��|݌��;�?Q/ @f�?l3��lf_=EƇ>=�=��=W�H��C)��]��nb`>�7J?������v�$�l���>��?���?���?̓c��	?���P��Ga~����7�A��=��7?�0��z>���>\�=�nv�Ừ�Z�s����>�B�?�{�?%��>�l?��o�B�B�I�1=%M�>��k?�s?u\o���Z�B>��?'������L��f?	�
@}u@Z�^?*�ѿ�6���Z��Z~��rh�=eS�=�4>���b`�=���<��:�;q���>�'�>�G>�ޅ>�%�>R�J>,�*>�ԅ�κ"�����_T���<�ؒ�I��03k��<��!��~��_��S�վSbؽ4����_�}\�>@��$)�ًK>�dL?29Z?��t?Q�>�v�CQ�> ��F��=fvv��?��i�>�e.?=^?�� ?�3;>���b|�^������I�j�3��>��p>(>��>��>�=%� >(r>hi�>�|�W!>CÔ� j�=��>���>�f�>D�~>.Jq>S�5>�;��c����Cg��Mf��W����?�{���Z��������b���'�=�:?�t>���4�ɿ�I��?ZE?~�����}���+>��:?@>O?�G>�i���0����=����O� �&>r�.�Ɗ�&G%��{>J{?~}h>��u>t�3��q8�V�P�!��Z|>��6?㵾��:�H�u�"H���۾:N>=Q�>B�=��m��Ȗ�J�n�i�@gy=FF:?�?~����n��/�u�Qힾ*�Q>Yu]>��=<M�=IM>
6a�sɽ4I��11='_�=ec_>�T?��+>)�=q��>cF�� �P����>q B>n,>E�??�%?�e������K���-�'�v>�`�>�ր>S>�cJ�t��=�h�>��a>p��������C�?�dkW>�
}�X3_�;�u��x=����i��=�y�=�( ��=��k%=��~?�~��䈿}�Fj���lD?a+?��=8�F<R�"� ��G��i�?+�@m�?Ё	�ȢV���?�?�?���E��=�{�>�ӫ>Qξ?�L�b�?�ƽ�Ƣ���	�D'#�!S�?\�?�/�vʋ�{l�58>_%?�Ӿ�p�>��fa�����O�u��s%=Xl�>TKH?�G��� P��>�|}
?V?K^�?���m�ȿ��v����>��?���?=�m��A��C�?�Kn�>ƙ�?�UY?~li>��۾�AZ��Ì>Ч@?�R?��>\L�n(���?�?V��?���=�Ӣ?'�v?Rf�����i�$��䥿�����Ծc��>)�D?f�D�Yq���a�՗��� ���񘿃����>���=us�>T������s5��@(W��3��Ƴ��L��>�&�>{0�>���>�H?�J ?5	?�4�>gW������~m�� \?�?+��y�e���Ǽ'��=#DS�S?1f6?���~��9�>	m?o`y?)`?�/�>�-��s�����޾�au�;"!{>���>�K�>��_�,>w8�ECJ��K�>,�|>���<�]оh�?��۞���]>��?z��>��>H� ?�#?՚j>�%�>�aE�n9����E�3��>���>HK?Z�~?[�?Թ��Y3����a桿�[�g6N>	�x?oU?6ȕ>܎��8���]>E�lPI��������?[ug?�_�g?�1�?��??��A?A$f>����ؾ%�����>� "?`�/�A��d&�:��w?[?��>�X���ؽx1ܼ�������?SG\?�5&?��a�sTþ�#�<��(��d�6Z�;�:>��f>1�>����5�=KE>	�=n�l�	�5��6k<Z&�= �>>��=6C6�@����F,?�WN��9���=.s�C�D�φ>9rK>�Y��#r^?�<��K|� �������U��Ǎ?�f�?%��?+&��Q�h��M=?��?�?ܓ�>������ݾS���Vw��y�!���[>Et�>&ca�X���Y��UL���b����Ƚ��R�8��>}�F>���>�?܈�>���>�ꉾ��7�`���p�;��V��M#��V<�;G�?t&�����L�\�>C�=`�˾/����>��ý��>U,?S>$^>�?�Z�=Aɬ>}�.>	)�>z��>aP.>��{=k[�=O��=���=��T?]���u_)�������=B?��]?���>4.�W���X�|�!?���?�?atu>��f�m�*�"�?fP�>hf����?ns8=��i<�9�<"��R#.�̗��31��.�>��ֽ�6��1O�*h�M1?�7?. ����оժڽ�!��ˉ�=�;�?$D ?�!�uAJ�-o�tK\�P^�y�n��
O���)���z�,y��?B���E���9 ����<�{?���?������N�ܾ��p���@�ӄ�>@A�>t[�>km�>ɖ[>�o���4��R�y�&��-��Y&�>��m?\�>GK?�+C?�U?�4?�>>��>��ƾ�?��I<N;,>
��>�M"?�8?��#?��#?�_/?j�= U����%پ�?�4?�?��? ?�.�u*��ٻ�J>ƨ��@��$���Z����c�=i>]��>�#?�����8��z����k>��7?%�>�f�>Y@�� �����<P��>�
?:�>�$ �jnr��	�t��>"Q�?�z
�w��<�F)>6B�=ȶd�����|�=P�̼	��=~f��6���<��=&�=g���)���L0�:?B�;��<�t�>"�?{��>�C�>a@��� �C���e�= Y>+S>�>�Eپ�}���$���g��]y>�w�?�z�?��f=*�=���=�|���U��}���������<�?JJ#?5XT?\��?u�=?rj#?�>+�iM���^�����Ϯ?�,?���>N���~ʾ@ۨ���3���?:>?� a�T�}W)��;¾�Խ,�>#B/�R~�h���� D�ױ��1��c���t��?仝?[$A�<�6�*�9����^���{C?}�>?�>T�>�)���g�0�l�;>Rn�>x�Q?k�>�!V?c{?#�P?��>;�@�p|��`��� �e�Z>�YD?0��?`��?EZr?��>hs�=j,$�)g򾳆 ���-�������L�=��Z>`!n>I��>�0�>eH+>���>#�R�*�1��=��>?��>:��>Xq�>��J>n%�]�G?=��>�b��C���菉������<��u?ԛ�?5�+?�
=�~���E��9��U�>�m�?���?�0*?
�S�J��=�׼>ⶾ{�q�'�>�>�(�>P��=2nF=M~>~�>��>��<\�t8�F�M��?�F?Y˻=��ʿ��D��$��U�!��½Gξƃ����ռ��ռdf>B�޾q��M˘�G������"�j?�(�O��^6�k6�>�?=��f>7BS>c�H=��=:�<�%���=���=Z1��=^�=X��;\g׽NG��	���f�<a��=jV=U�˾/�}?_;I?��+?��C?-�y>[@>؜3�n��>�{��
@?FV>u�P�e����;�{�����i�ؾlu׾��c�r˟��G>%UI���>f83>�>�=%J�<��=�s=Yǎ=7R�=� �=�O�=�c�=���=�>�S>�6w?X�������4Q��Z罦�:?�8�>a{�=��ƾq@?�>>�2������xb��-?���?�T�?>�?>ti��d�>L���㎽�q�=B����=2>q��=z�2�R��>��J>���K��A����4�?��@��??�ዿϢϿ3a/>�R7>:>P�R���1���\��yb�^Z��!?�;�?̾}�>���=��޾�dƾ��-=�k6>%�b=��<0\��b�=�{���<=��l=��>KD>ݐ�=�6��齶=�K= �=��O>�����8��
.���1=���=��b>l]&>���>t�?'k0?Z\d?��>T=n�Q�ξ3T���N�>�+�=�"�>�'�=ۊB>F��>T�7??�D?��K?c<�>��=�>���>��,��m��f徿����=�<8��?�ņ?ڸ>Z�V<_SA�!��	c>��Ľ�x?�?1?/p?��>���4z׿J}���6��Cu=6�<h��=��c�*��߭��T{��8D�<�V>���>S�>���>���>>N�>���>�Y=_�ͽ��=]�'>9�(�������=��,>'������,:�q���f����:>V�ݹ�꼋���h�D���=pF�>t�ӊ�>ƛb�pž��u>>����j�А<f����d�X������$M5��XY�s�M>'v�>WD��3�����>�y2>��=֏�?��?���>J�z�'+۾g��.�W����<�	>�x�>�E���"���3��\�=Ǿx�>!Bu>��|>=�~>=�>���C�W|g=R�侑9�ӫ�>�z�33��]�d����ס��/����\�d�>��D?5	����8>�{?��2?�ُ?���>Ϯ����q�>�̐�C��g�
派��"�j%?X� ?G��>%	�W�L��H̾`���޷>�@I�&�O���N�0�ԭ�)ͷ�D��>������оh$3��g��������B��Lr�j��>*�O?��?�:b��W��5UO����8(���q?�|g?0�>�J?�@?5&���y�zr���v�=�n?ĳ�?O=�?�>���=h�
��G�>�\?���?�Q�?	�?Ww[��2�>��=�[?>����ˠ��2�>>N��=/*C>�%?�q?�?�󅽼j��P澅⾣[����<��=u��>�_�>xy�>��=�ޟ=��>fk>��>�t�>��>�{�>�>8Ų��&����>�
>��>��S?ߖH>�=}?��.�X�=>����&~�?��_+���;Z�=u>��!>M��>��ƿ���?<�\>m ־8�?{��� ?�>N	h�H�Hb�>*��>�,[>��>4�?ѿ�<B�>0�=_ۿ����=c"���+���)��!'�)� ���>Ġ4���L�}�!�k��!TP� Ġ�ߝоj%Z��8����:���[<�̞?��ｺ�����X佨�5?i>I?
��
�Ջ>-?YE�>��.Ӓ������(�r��?{�?�;c>��>J�W?!�?�1�63��uZ�(�u�n(A�,e�Q�`��፿�����
�v��-�_?�x?+yA?�Q�</:z>P��?��%�Sӏ��)�>�/�'';�(@<=r+�> *��"�`�v�Ӿ��þ8��HF>��o?:%�?sY?3TV�t���00�=��@?�1?�o�?1<?u�R?��K�I�?#0�>g��>;��>l�?s�3?D��>up�>dY>*gֽ �1>��Ľ
��������7���=[�=��X<o2E�'�[��H�=�^�<�����V�Q���Gn�i���ia=���=te*=���>;�]?�V�>���>}�7?���`8��Ϯ��%/?��9=ϸ�����㾢�z����>��j?���?bLZ?�Qd>{�A�[#C��4>�_�>�c&>��[>
f�>�z���E���==w>�H>)��=�GM��ց�i�	��f���Z�<�>���>�k�>�|���*>;���]~�[�`>�U�M��S>[�C�I���,�uq���>I	L?�?.:�='�쾸��vNf�I�'?B�??��M?�6?yHu=�IϾAn;�ۜI�E�!����>���<��薠�;ơ���:�\�<�l>�	��Ȱ��`�j>-��tؾ��l�%G�jR侳x=�l���=b�
��پ�逾-��=��>�C��)##��+��g����lF?gZ={���V�M�NZ	>=��>ʣ�>I],����?�<��֪�R��=���>hC>�Vo�C$供MD�Y��͋c>!AG?�jb?�ax?���n���Ƨ������z���?�ۧ>�>�l�>��=�{���C��k�h�ȴX���>k��>��
��1��)���>���p��>"?���>u�?��T?��?�Od?�:?�?��>ͷ\���F&?�~�?7�=M1ѽw}U�p�8��E����>�*)?\GA�gj�>5�?�?G�&?��Q?w�?��>� ��C@�ZE�>M'�>��W��'���_>שJ?�-�>�<Y?���?�r@>��4��g��*�����=?�!>�Y3?�.#?ݑ?�=�>T�>������=���>�+d?ڐ�?�p?H�=�?O�@>fU�>�7�=�o�>��>��?v6Q?Att?��H?�5�>a6�<̽��W��F�m��as�0"<�P<ݍ=���\ہ������<X�:�yϼ����I���qj��ۑ�#��;Œ�>�r>�t��Qd1>@mľT0���w@>$��������`��n/;�O�=��>�&?qa�>n+#��Q�=�^�>m��>	��5(?�5?r�?��:|b��Qپ��N�Y�>�A?�T�=��l�����]�u��	k=��m?l�^?W/W�E���b?�]?�g�9=���þr�b�9��)�O?l�
?3�G���>��~?��q?���>��e��8n�T���Ab�{�j�zŶ=�q�>uU���d��A�>a�7?�Q�>�b>��=�u۾�w��o���?��?R�?f��?�-*>/�n��3�����F����Z?�>��y�أ??���<�q� �~��,
ʾc�;E�c�t=�� ���R�k���41��ٔ =��?d;�?+al?�<L?{�?/e���]�ԥu�IB��,�E9���&�p[N�+�O��τ�M"��y��$ɾu�)��d��$�1�y�?y�/?��w�G��>!�{`ɾ���1�_=�O��KM��p��<���=I�6><d�=�R����o��+��/?���>:��>�eC?O�p�[���'�Az��*��kHR>�?&*�>Ő�>�����r��;�������su�<7� >56Z?��_?^R�?�o!�T�3���t��E&�ƴ��J��7�=^k�=�d�>]Oy<ߟ4����8:���u��Q"��_n�rQ����=us&?�?�=K��>ݍ�?L6?CK���ݸ��s�=O~�`��WW�>TlW?u�?hv>B��$��'��>݊l?�>�>V�>��x�7�*��^l�/(�q|�><�f>�W�>�\�>�
4���^������|���-��R�=΀j?;\���I�d5�>��W?�� =\0ݼ��>�s���2�q����D��ja>���>��=Y�$>�}��"
�JE~�c��X�(?�8?����)�:�|>�0"?���>Zm�>tك?\s�>��þ���G??�	_?~�J?|�A?17�>�N=S����UǽWN'�M*=�	�>�q[>s5n=[��=٬�ȲZ�z����K=���=�̼���8Y<ۮ�I�P<1� =V4>�jۿ @K�2�پ�	���08
��鈾qɲ��c������`������^x�q��Oe'��V�&@c�����
�l�m��?u=�?�����3����������������>=�q�,������/���ྭȬ��g!���O��&i���e���?���O�ο�^��r�����2?W��>���?y�W�𾡛6�5bL>���=K��=~?ξ����Dʿ��j���S?h?���5��u�?Ǆ>7��> r�=w���ڬ��|��=-�?C?�\�>`�Ǿ<Ƚ�+ż�����4#�?�@cVA?��&��d��n=��>%\?�IG>S�2�B�������>�?��?�zE=wuW�����e?�/-; �E�s.���=��=��=�]���K>pP�>D�$��C���Ͻ[:1>��>��!�ū�\[�9��<�)`>�ٽ����τ?ky\�f���/��V���A>��T?��>(Z�=X�,?X0H��zϿ�\�V�`?�/�?ޟ�?��(?�{��	�>9�ܾ�M?wG6?rߘ>I[&��t�#��=���S��|���V�L��=��>�`>T�,�`|��*O�����=N�����ȿ��Vv���4=�+�=ҳü��x���*Pν�?��Ǌ���r��%�=�>Y`>ꅅ>sZm>	fC>�*P?��g?sZ�>X�>�w��㉾<�˾p�?��`Q���I��O��Ǥ��<��'��ͯؾ�� ��\%�8`�ˁʾ#+a��է�ĕW�i]���S��g�d|I���4?-cE>����Ud�M{L=����1�+�ղ�<��>�ޣ���2���i����?�G?@��̣Z��="�9V<��=�m�R?T�<����־L5>={=�>���>�b$�x����4�4�E��KZ?�t,?������G>U_��=����O?w�:?-EU�=��>�eN?�u��󡾾eh��&>�׊>	[�>��><	¾�4��^(?1�c?f���$ɾ2��>���p𾦭��fO����!�B���>�Ƽ����t+<:̗�u
���z?��>�����#��bؾ[&=c'�%$�?��=?G�\>�.�?�G?۷�>�����O�x!,��cɽjGP?�bz??->J��� �龒� �~�V?NWy?N�U=!e�6J��Eq]������?��\?U �>&t����u�޹��v���HE?�Si?�k��i��+5ܾ{,z��Y�>ְ�>�C�>��%�J^�>�n ?4V���|���q¿®����?���?j��?��
>d�7^k>��?�I�>�ʑ�=V�q Q=ހ�w[�=)��>�q���j�TI6�A;���A?Q��?��"?�fQ�3��F�=O���F��?�ł? ��YJd={���m�����1��1�=:<���N8�V�T�=���ξ�t�p��G�A��)�>��@3ݽ4*�>�L^��C޿�^˿����!�ྋ�C�}f?��>V��q���r�(�z��M��J�)勾 8�>T�>p燽� ��T�{�5�:�ziI����>���Q�>T�R�D�(���f��<^H�>�&�>�̆>�(���~���B�?�G��!uͿ˝�Y���W?W��?}��?�) ?�}�<h�n��zw�Z����F?x s?yTZ?�:�!fX���+�6Th?����d��.��A���a>�+?:-�>�.*��Q�=�K>��>y�>��1��1��Iд�^��;��?m��?�\����>�s�?��(?D�������m��|1���'<�Y;?�->��ʾ�O%�IGB�IA����?=-7?\ؽ���X�_?,�a�O�p���-���ƽ�ۡ>�0��e\�*N�����Xe����@y����?L^�?g�?ݵ�� #�c6%?&�>h����8Ǿ
�<���>�(�>�)N>DH_���u>����:�i	>���?�~�?Nj?���� ����U>�}?塸>��?���=�B�>��=������7�&>�=�e���?��O?kV�>�M�=��<�J!,�~�D�ܣQ����]�C�x܅>B�c?��K?|�a>�w���:�i�#��E��V�3���O��G��6�ʕν,52>�D9>�T>�T���վ+$#?�e5�տЁ����j�B?Yڼa6?׷�ۉ��L<w';?�q�>�����������߳n��]�?z��?���>*6���)=P�V>ENk>5�=E��<�X~�g*��g{>�Y'?m\��]t���)���C�>x�?��?�h�?�`+���?S�	��y���Lx����zZ(����=��4?q���݈>��>�H�=�r��󪿥-n���>g��?��?(��>8i?,Jf��i9��"*=�ޘ>��c?m�?-���t��7>ES?B��䏿g���g?�?
@8@�^?�7���i���l��ϟ���8��,�>�5�=,xU>��];��
>@�>���ek'=��>qy�>�j�>{?�>f2&>�=��~�������V���h�4�B�4��l=�r6���lؾ?�n��'�X���������	 <�� 輨ڃ��Vh������E�FR?�Hc?�!3?w7�>�8����;����	�3���	�=��a>�<?Oa^?��<?���=���W(r�ď�D�=����>ٸb>���>fܯ>��}>�e�=:�m>;RX>$TB>�g.= v�=�d�=a>=��=R&�>�+�>�B�>�g�=��;�+�������nT�:]a��7)��/�?������-������ S�+��>>?(1?�1>G��{ǿ?¥�u�c?�̵�OA0���Ľ��=�kI?�_9?�8G>�mӾΆ�x�Q>p�d^���ǳ=g��0EѾ�E?��<�>Qb)?j�`>��s>:�/���5�ˊO�������>u�5?a[��nD>��Xv��xK���޾�*U>S��>�|��R��ᖿ�����c���m=�8?P�?u%��bﱾ�m�W���7�M>܋V>�:5=#�=Q2J>^\��+˽-�I���7=!~�="�]>�?�.>&|�=��>9����P�p��>{G<>�A*>)�??�#?-����8��w:���7*���z>���>��~>��>�GJ��°=]��>}`>ZX�{�IY�s�=��Z>|[�b<Z��Gp����=�ǋ�I�>�= ���'P;���=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>�T��U�����u��V$=��>CH?K��kP���=��z
?�-?�e�ꥤ���ȿ�}v�b��>U�?��?;�m�A=���@���>��?=RY?/xi>|X۾x�Z�3r�>d�@?��Q?�>c4�D�'�O�?Kڶ?ȯ�?�=ѥ�?;7q?xB�>-΅�*�7����\��S=g���r�(��>.?>�׾`2��ʉ�$�|��B��D�.��yG<�<�<�O�>�q$��<���=�,r��B��G�z��ފ>��$>��>���>���>���>�<�>u�#>އ�w����ܾ}�K?���?����2n�K�<*��=e�^�s&?_I4?W_[�`�Ͼ�ը>ʺ\?g?�[?�d�>���B>��3迿'~�����<v�K>�3�>�H�>�#��6FK>s�Ծ�3D��p�>З>����6?ھs,��v)���B�>�e!?���>�Ү=�21?��&?{�j>�k�>4�t�+M��ϊ.�<f�>�)?��?^�?�r	?;T���]₿���;�D�jI>$h?��7?(�>w��~���B<��<N�R�O�?��?e��Ɗ!?z��?�i?ҏ�>�}�=2�u�����V=S��>\ ?��C�>���$����p	?��?���>mv���ݽNo	��U�����X�?4]?g�&?�@��va��(ƾ��<P�L��y����;�v�S}>�>����u�=
h>q׸=Wn�S7�&zy<��=�ː>�h�=K4��Ս�jN?]���	��۱�=b�x���7���|>��=#p��3,h?�LQ��-��z���ެ���8׼b7�?E��?���?5�����o���U?���?���>V�>���C���*I���ʟ�����y����
>_�>�󛼛M�_���������9t��-��1�>c<�>f��>��?!+�<��?�zϾ>�>�xh���~3�d�2�I�+��#�|l�����	��Zm�h�8=zA��2���2�>��8�`�z>}�?\|>�7�=�Y�>�p}>a��>f�=��G>��?�݊>�@&>7�l>�u=H��lRR?������'� ��h����3B?Vdd?�C�>�:h�������l�?���?3j�?"v>$�h��-+�mq?GQ�>���(l
?�:=
#���<�V��h�������O��>�D׽3:��M��~f��g
?�/?�茼��̾�)׽���Ĕ�=wȁ?�?��+���-���`�� ]�MES�c �]�3�����\%�(�b������w�����%��ռ�Z?֔?������W[ھ�&i��$8��Z>�:�>J8�>j��>/��>�����(�P�O��1$��淾�\�>6�f?��>i�G??1C?Y�^?�5?&��>��?�~޾�3�>�L�>�~�>��?��3?�<?p�Y?7GU?�T?O3�=Yv�~����پ��?�|�>9�A?�?`��>�:ӽ�rd=�e>%A�=��j��	�JF�=1��=5�#�猤��� >��>�8?հY���2�e��B�A>��2?���>��
?�J2��i���A9>���>I\)?{��=U��}y��'�1��>���?�H�2J�<\@�=>��=H�<W��0qz=�52����=a�	=�r���������zw<��;�r�=
�>�<8�;(u�>V�?g��>}D�>j@���� �;��ha�=�Y>�S>�>�Dپ�}��{$����g�0[y>�w�?$z�?��f=�=���=+|���T�� ������<O�?�I#?jXT?��?��=?�i#?��>"+�aM��0^�����1�?�,?�(�> 9��FɾIw����3�#�?p�?a���T�)��\���K׽9F>c�/���}�랯��fD�^1Q����ǚ�l�?Sl�?|�K�-N6�����#��������C?H��>H�>\��>x>)�J�g�i��0<>��>x�Q?B�>�P?zE{?�DZ?gQ>�>9��ʬ�����r���n%>9�>?��?
�?Ly?�s�>�v>
e+�PN�{G�����rW��-��-��=�	U>ٷ�>���>,T�>j��=:����,���D��¯=D�e>���>:D�>g��>gx>���<��G?���>�Y��V���菉2�����<�+�u?���?�+?�=Ix���E��I���K�>l�?��?�3*?I�S�%��=�lּ�۶�l�q�� �>�ѹ>o-�> Ó=��F=|u>��>@��>/�1Y�~f8�!�L���?4F?b��=A�ÿW�l�����wY���>�}y��Z>�R^O�Uh��>�������m����6�Fd���Ɋ���,�y�n��l���>q���Y*>@Y�=��<+�J=�m@��ʼ4H�=�#;G���[Y�=��*����=��R=F>��]�=⢓=��Ѽ�˾�}?RSI?3+?�C?;x>\�>�;��&�>ע��7>?dV>�eR�K��|�;�i���?-���hپ�;ؾ��c�OL��cb>Y�G��2>M�1>���=�r�<O��=��q=��=�,��N=���=@��=��=�$�='1>k�>�6w?X�������4Q��Z罤�:?�8�>[{�=��ƾr@?|�>>�2������{b��-?���?�T�?@�?;ti��d�>G��㎽�q�=K����=2>z��=x�2�S��>��J>���K��J����4�?��@��??�ዿТϿ-a/>o�6>(>��R�<�1��[�mmb��&Z�Tw!?fS;��5̾���>$��=�F߾ppƾ�U+=Wd6>/_c=�[��%\�cI�=��|���;=��k=f�>��C>�w�=����嘷=D�J=>��=_�O>���ǈ3���*�63=ݸ�=@yb>H[&>�p�>@?M1?9�n?�p�>�����e��A����>.�=�}�>�L=�;>���>=E7?�@A?kF?�>7=7��>��>u`2�*la��4���8�� lɼ_��?0��?�}�>q��=�S˽�9?��sͽ6\
?��0?��?�j�>S2��q�L&�H�.��쑽+�:�W,=(�q��W�Z���,b�M�罓�=��>��>���>��z>�\:>�O>��>v	>���<�օ=�ד�_��<�$���C�=�s����<*��V�����,o)��8��gY�;t͖;]]<���;G�<��>���<ɟ>�@�=�ŭ���k>�Ҕ��oM��E�=�K��xE���j�舿��.��
��e��>�4�>��}��H��G1�>��>Zy�=Ҷ�?)f?�1V>J���=���X��{����_�>P�=�>����6�c�R�Qn�~+����>Z��>�Y�>`cr>��(��@���=��ݾ!�3����>������ļ�4��3q�6����C���Eg�𬻧CD?���(��=�?I?!�?�V�>g�z�g�ݾs�>����(9�<�Q���q�}{��¨?�j%?fo�>8�VE�*5̾s&��ӷ>aI���O������0�����̷����>V���о
!3��e�������B�N:r���>��O?��?�#b��P��KO�����5��(w?�eg?J�>�L?iB?G��qx�2y��J��=�n?��?T:�?E�
>Qؽ=JЯ��>X	?���?Y�?
yt?��B���>H��;�Z>��j �=O�>�=K��=�P?�D	?�	?�ӝ��u	��2����?�\���=-r�=�O�>ݭ�>m�x>{�=�o=擨=�Zb>-!�>L�>��f>���>觇>ܭ��3��W�>���<$��>?�R?Au�>� C���A��������ޞ���e�<=>���0�D<�W>533>�p�<d��>/Ҽ����?�f>FM ���-?�����
�5oD>��Z:��՝�>W��>�=�>.�>jz�>A�^�lz�>*�ؼ�5оR�>����mD�tQ�_0Ͼ5��>T���3�!�������i8D��3����]f��'���<���|<ȇ�?u����Un��%�ʎ���?~�>�+7?/N��'%O��0)>��>\�>�6 ����������A��?@D�?�Ac>��>�W?�?��1��3�>pZ�g�u�"A�C�d�K�`�+⍿5���ɠ
�����e�_?��x??�A?	C�<�$z>ץ�?��%�Nԏ�I�>& /��;���;=�)�>p,��L�`�$�Ӿr�þ�K��YF>�o?z'�?rS?vrV�+N�R0->�};?U3?��v?[23?�=?�h��M%?L�N>�%?�g?�~4?��/?�o?�H>�$>d���Ϣ.=���B��>Ž��Ž�~�C�Y=/=�Ed<٫�;��=���<]���t0�O5�9׼���<+�=�q�=@)�=�K�>	�]?4��>��>z7?� ��u6��ͮ�b�-?k� =�ᅾ�Ȉ�/=���E�=p�i?	m�?)6X?��d>"A�$�C�R>�׉>j!>�[>�۲>�E��ZG�3V�=~
>o>��=H�F�˷��[f
�꽏�Nܻ<Q�>3�>}�>����X,>�Z��mY��Gh>Z)P�%1���w[���H�m�/�+�v���>�0J?v�?_�=���q��8�e��(?2@=?�ML?Y}}?��=�׾H*<�pK�P<�fU�>T�\<s/	� ���!Ρ��P;�߽Y;�vm>)���נ��c>M��ݾ�.n�iYJ�����DJ=���L|P=�t���־`���k�=0�>�c��0� ��(�����\�I?��g=p�����S������>�6�>� �>��8�ٜy��X@������=,��>�:>����V�p(G�T����>RI?�P^?U��?]�E�,Cw���"�(�j���n���*?֘�>}U?�/2>�T=�q��B���`��F�#w�>H�>��Dh@��7��Zg���/���>:}�>��}>.�>K�3?2�?*`?"�E?���>�Г>{���n�˾�/&?�d�?�9�=lսT�V�8�9�E����>��)?ڗ@��>�8?��?~?'?��Q?�?L,>�� �x;@����>ta�>T�W�S��M=_>�eJ?mO�>�
Y?��?#�>>6�5�`����榽���=��>��2?,c#?t�?���>���>�6���'�>Ե�>�P5?"�?��d?�A�=���>I��>Xݒ>�[����@>�I?��\?&��?�v\?]�?<�w>Ì�=�
��н6*�=好����.��k�=ѱ<�!=`F�=/T�<fH��6O�;U�=t�=�h=��%=3`L���?� �>r��o!�=_���=(���=X�>���'o�+y���Xi>gP�>�K�>�̉>�#�p�=F��>m��>���i /?���>[�?p��;�T���sR��A�>�|M?��L<A6z�;���Tt�9A�=��e?;\?��$��Z��S�b?��]?�S�3=��þ��a��Y龎BP?��
?�I��<�>Z?,Fr?'S�>ӳf�`^n������a�o�h�%�=�C�>bQ�$�d���>_�7?���>Lc>y�=��ھ�w�R>����?���?��?<(�?3+>��n���i��]1���&a?b�>N����7?;Pӻ�žk�a�g�;�������U�m5���A��=qڽ��P�'��-3�="�?s��?��?�U?{�ܾ-zb��.T�w���b��'	�u���};��s;�a�L��b���|�r	�1�ݾ�LG���x��W:���?$�)?Y�D��-�>Ah��� �n����>K����8�3L�=�*&����=�pl=�0m��
B��x��� ?���>���>h7?}^��.<��&-�]<-�����S$>ĸ�>�ό>���>˗v��m�s��mS˾����ҝ��n�S>�7r?��X?@�i?;�@���I�b2[��1��|�<M�����>l�<[��=ay!�59�;�0�X�d������I��&��ӂ�Ң�<�,@?q�n>�D<��?Yt?��;��ؾFt"��44��*��7E ?s��?���>��>����u<�l�>4�g?�x�>B�>�鍾.�>��0�%�b����>��:>$]�>�5�>һh��@�����9$��߇)�?��=H�q?$��+�R���>�:T?L�={���?4�������kG��m>j�>��>k= �ܤ��"���lb�$�|�c�$?.�>(���>53�W2>C�#?�:?�9�>)�?r�?�ľ�޽���?9��?�܃?xo?�?V=�����X���,�L3���Y><�=>*=�AG=#gν�<��7Y����=p�4>\��=�sn�lb�<&֣;G2:=`�=���>j�ۿ��M��7޾>��T���N�}��������y����ۼ�����fs��) �����U��Y���hTp�;��?*-�?�c������ڳ��?��������>��S��e��AD��;�R���tBܾX���R�ٔJ���b��b���&?�G��ױǿ�m���wؾ��?6�?D�y?�"��k"�~�9�iY#>}�<�%��$��n��G�ο)ܚ��0_?���>'�C{��{�>N��>M�^>��k>�)������ƽ<kM?QK-?���>�x�ɿs@�����<J��?�C@�A?�P(�U�6O]=ɢ�>	?�C>V�2�W
������>C�?��?
�K=q)X����-�d?
z�;HF��&껪��=��==����K>��>���C-B�[�޽'4>0C�>�- �:[��^�ʩ�<��\>�mս_5��Մ?�z\�`f���/��T��<V>��T?�*�>`@�=2�,?;7H�}ϿF�\��+a?1�?���?��(?�ڿ��ך>��ܾ9�M?ZC6?��>�d&���t�΄�=�0������'V�2��=L��>&�>��,�f����O��E�����=(4�7w���$�;"���=�m�AS�c��%�>KM�=�]¾�i�I:��#��=d@>�3>��>�'>� R;��J? �k?�j�>)��=�y;�����ھ�׸=�U�����C�׾�qm�4�����ɾ�U��'�����3�,ݩ�+A���ͼ��N��萿p���NZ�d#O�r&?��>B�޾��j�k$!<b1�p�����u<�r-�[�о9���g�EP�?$,T?4"}���l�kL�?=�Pܽ�,c? ������?q �K<�=�&c��ei=>[V>�f���h�=������N?J</?'���Ę�	>��;�����N?j�>�=�F�>��.?x|��96��c�9>-�>��>���>ܳ>Y�⾛�}��2?(Ua?&�{��
��?v�O��R�R����X%=�Ⱦ�o��:0�>�'���;"~��i�:��s���X?aW�>��(���2G��;a�_H;=��{?��?�͕>>l?��G?�]7=G���nT������:=��V?��l?@�>�)����о�Q��9?�Hi?g6I>"�T�y�/���?�o?�Z?�ࣼ?�w��Đ�4��`\7?�~?��O��6���@���9��ȼs>%N�>��>�9q���i>ǹ?���t����տYI%�}?���?f[�?;wK>�cѽ��G>q�?�&�><
�k8��>h�־ur�<�ˑ>��H���C�2ʾt�G���>�4M?O�?���fP�9&�=�HS�޻�?	v?�=��}�o=7�	�&�]���n�S���>�򠽾��<�3�D�K��=��g`�a���^�E0q>}�@������> g9���E�˿��u����� ��Uc?&�>��F���¾����g�t���d�4u�(M�>S�>���E�����{�r;�y�����>�����>��S��)������}�5<0�>Ů�>=��>~8��'뽾�ę?�b�� ?οk������ �X??g�?�n�?�p?m�9<r�v���{����*G?��s?Z?fn%�"7]�'�7���k?�=��w?b�1�A�D�_R>�/?S��>ڮ/�ߺi=��>�>�|>�3��!ÿ�X�����=�?���?��C�>p>�?�+?�i�-���ޡ�C+���;,;??�->>����!��;�\}��I#
?C.?`����.�_?��a�i�p���-���ƽ�ۡ>��0�1e\�@:�����jXe�����?y����?]^�?z�?Ӳ�� #��5%? �>ɝ��J9ǾN��<��>M(�>o)N>F_�I�u>��:��h	>z��?T~�?-j?����p����U>��}?@�>{��?��1>;?q�>�˾vt>�e���=≾���>�)c?m��>�P:=s���)��B��A�7�߾�G<�>��>ޅU?��=?=*�>m֔��9=���)��@���ֽ��.�u>�i�R=�½~��>�h>��=�\Z���yC?J� ��Ŀ�U����I;��;?�]=o
T?�nľ�Ȼ���=Z��?��>?���������oPa��Ț?��?��?��žir����>�Z�>���>D-�#hu<�(����>C�:?x#T��j������ݰ>�>�?R4@Ys�?�D�D�?�U�i7��{Cf���i���
Ի��:?J��i��>���>N�}=K샿h�����`�/��>9�?��?*U?+Xm?�n�0�7���G>���>W�_?8�?�J/�u"����E>��?��*�,�~��	�0Y?�3	@��@�Et?����f�ſ�/���<Ǿ��7��i6;�>f�@>у��w��=R�	�z��\9=�k\>�׵>ȥW>i(�>݉>�	>���={�~���#�A ���Ҁ��>R�Wq&�jP��X�"�ᾓ*.�#ܾ�{@�_���=�<b�I�Լ�OG��T9�<�����={p`?=�V?;�?���><��x��>=V)�^�=�H�\�:��@>��?dF?�tJ?�S=RȰ���x�󩎿�4��(g���>e�>��>Й�>R�>�X�=fEO>�F|>m0>��.=	>r�=���=G,�> )�>�)�>PW�>��;>\>���7��f"h�5?w�qͽO�?�+����J��K�������tz�= K.?��>����6п�孿�SH?�V��F��-�n�>m�0?�&W?uz>�ܱ�ATV��>�8���k��,>ɪ �,0m���)���P>��?1�e>|t>>k3�U8�V�P�e���[�{>�6?�w��y19��u�ԱH���ܾ��M>z��>�)>��K� 閿��+i�9!y=�:?�?A��㐰���t����ÏQ>m�[>M�=��=�\M>��d��Iǽ��G��/=�h�=��^>�e?r�+>P��=%	�>OO��Q>P�n�>��A>��+>=�??�$?C��X!��h���Hf.���v>�,�>��>>�JJ� ��=��>@�a>���H��G����@��PW>�U���{_���t�e�x=�S���^�=c��=<� ��=���"=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�I?[i������:���F�c�%b�<R;�>Xr?؍��\Z�2H8��??�!?�eվ휿�2޿,�����>#��?��?�Sc�G����G?��'?�@�?X%?5\�>?��nk����>W�n?xlX?{͢>���ִ��*?Ȫ�?Tϐ?[��=�>�?�^�?�;�<k_�����\쬿���g¸��b�>�P?����5����(�)��կ��]᜿,uj�'�5<G��=���>/	�)���]
>΋��0I�aM�,��>��>Hr�=�j>��>��>��>�K��%��v�A�O���g�K?���?����2n�S�<���=R�^�I&?bI4? f[���Ͼ�ը>ܺ\?\?�[?d�>��G>��7迿1~���<�K>�3�>�H�>v"���FK>X�Ծ�4D��p�>�ϗ>�����?ھ�,��WB���B�>�e!?���>RҮ=ذ)?�3"?��g>3�>��e�����53��$�>.�?s��>��|?$V?�`����2�?֐�T߫�M�b�oV:>��w?QA.?�lc>Q���I��$�j=:�=�����i�?�W?I!��u!?\�?�GO?�9?�
>Y9��mN־l1T=��>��!?���A��D&�&��Ĉ?�[?z��>[��=RԽ�׼>���]��i&?�L\?b&?Lh�Ia�#þ(n�<�� �:Zc��[�;.
H�P�>�r>�G���8�=�/>1��=E$m���5�pih<ԭ�=By�>Y��=*�6��/���)?'=)*��:��=����]G��Р>�#>�۾�)\?�y�#�v�����r���śX��(�?��?U֜?�$���r��wP?�i�?�-�>X?�x�kWʾœ��D���gf �t��gC>�K�>%ZF>���>Q���D��� ���B���!�U@�>�<�>z?T�#?�M>���>ʠ���Q0��\ ��&ᾘ@I�=M
��z�p�D�K�f�*៽�*k<�ξNG����>�W�����>��?�*[>>B��>I��?>_&�>԰�>��>@�n>!)5><9�=��-=��ս"m]?����^'��Z��
:���VH?p�M?�1?���X��0'ྚ;?�H�?n�?��V>�=Z�%��?2??V�~�7w??��<��<��=m�	�M����pɛ���>n��@��Z�*g�?�?<$=+������0����=Eu�?��(?9�(�>O��p�K�R�4[�����x��U����;�j��O��Q������%/��,�<�T%?���?Y�A��T���6i�dRL�a�O>]��>�*�>��>y?M>�����-���T�Ua.�����K��>�j|?�s�>��I?��;?P?�aL?Eۍ>�W�>����
V�>�<� �>���>K�9?}�-?�~0?�e?h*+?��_>a��������׾y�?ӏ?�d?�?�a?u��C��ٍ��W�Y�1�x�>́���=8U�<�ʽ��\�b�U=��R>�J?KW�;�8�������k>��7?�y�>� �>�)���d��(�<�5�>R�
?T�>� ��[r�pA��c�>T��?Bk��	=�)>0��=}����@��~_�=S�¼��=�k��0,<�� &<Ľ=8��=�#Q���:Y�;7��;��<���>d�?Q�>�N�>PN��]� �n��JO�=��X>}S>�>voپ	}���+����g��Ny>�w�?[}�?;]g=��=���=n]���@�����E%���r�<�?jB#?�@T?���?�=?�b#?ו>n&��H���^���#���?��,?���>��	�E���Si��Ɨ4���?�9 ?�6]�y�/%������꽆O>��0��~��f���@�z�<���������?���?�D�Α=�1࿾����D���<
<?Js�>��>9��>~A�;n�:�!��?)>'��>اO?Q��>��P?e�z?�\?j�X>��8����9����_��/>�Z<?R(�?�D�?�w?���>�>h�,����X��*)�U�͊���z:=7Z>���>���>ᯪ>���=ݘ��������>�h��=ZUh>ĳ�>��>��>2�r>���<�G?K��>>쾾���򿤾Qr��S:�xu?��?ʻ+?ot='}�V�E�wm�����>�w�?F��?*?�
T�N+�=��Լ"��hkr��ҷ>��>��>W��=��J=F�>��>�{�>�:��/�B8�"�L�s?x�E?�?�=D������U�v�<�޾�Iܽ1g������A<���=Y"9>cu��� �4���T[U�e��ja��q.��Q��ڴ��5�>�%<g�g>T�>->p'==�=/��=�&����D��{�=���ȅʽ����{G�<2�9<�x<w�ɼ n̾\z?9�A?9*?�HK?�l�>:�>t�:�ZK�>(
���?+�:>\�3��y���O�&���̋���ϾP�Ѿ�m�͔��U�>��\�->j�?>�2�=�S7<�h�=�U#=c�O=�^<(�=�=�z�=nƜ=���=K>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>s��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�3>>	�R�A�0��}Q�I�\�F<U��| ?��;�U�̾:0�>��=fK߾��žM�=��5>�?o=e��!�Z�R��=�}���b>=�ad=T��>Y�E>���=ra��꯻=	�7=&��=2�T>
M5���A�����z3=���=>Re>Z�%>�Z�>y>?��1?�4^?���>�a\��_¾.㻾��>�D >1ԫ>}d=C�>>���>])??�"I?�>M?t�>��X=�h�>~B�>ZM-�Ln��S��_���Ǭ<^��?8?�?oJ�>C#k��+@�.=�[�7�H5��4�?B+3?cY?u�>���X�b�2��������5�s�g,���$�	�=]�u>goT��%=�4>��>�˽>�w�>j�>�O�=ZR:��>��>��<#鐽��E>��=�,��t�
<�(�=0�>]�f;�����U9��% �\Mz<�a�8m���<��%�P��=�i�>��f=45�>t!>y���h�d>SW����Z���>�'X�� C��f��m��?�O�߽g��>��>6���
/��᡿>_>aO>\$�?�w�?xr�=8��� r޾����[=�Xtv��E�>���>1鐾�L9��yz��Q��椾\^�>���>v�>���>�&��>A��
>�?�Y>/���>O����7;�P���j�f榿���?5d��m��jE?�W��ȃ�=y{?C*I?�f�?��>PX"�-�� >�C����<*�	�+�]��d���?�>!?�2�>�	��_D��̾�(��N�>J���O������0�\F��跾�{�>P-��v�оdL3��`����|�B���r��
�>��O?a��?vb��^����N�����Ʉ��O?nbg?�>�c?K|?Fɢ��^��ڀ����='�n?��?�g�?�>N�=�(���ˮ>+J�>�^�?+3�?g�m?�:�k�>Up�=�
>��ܽ*��=x�>���;�l�=�?d�?�D?�ů�����վ/꾠�Ќ�=�>��t>k��>H� >��=>�>֐���$>J��>T�>��F>�0�>�L�>�@����	��9�>c��=F�U>��B?2B�>���<B� (�?��<ب�k����Д�����=���=K�m>kRm<}��>z俿 ��?>Ų"���?�� ���P<�a�>���=X�=��>!�>�à>��>�՛>Ow�=͸>��=�a��U�C>�jϾ�a��?<6�f�����P�>�N�����0-�`�T����{���(�Ѿ4X�;酿�K�:�f�*�?�ҽ뇿��%�Ö���j ?vR�=�c?�����@�="e�>$
"?�7�>xI��Ǧ����L�ž��?@=c>�>_�W?J�?�1��3�6uZ�֮u�(A��e�׻`��፿�����
�����_?Y�x?�yA?;V�<E8z>~��?��%��ӏ�Y)�>�/�e&;�,A<=,�>�(����`�P�Ӿߺþ(6��IF>��o?`%�?/Y?�UV�7A��%>wP?	?�ji?A�c?yN?�\����?[>���>�7�>FDA?��U?�%'?Z��>B^K>�j�a,�<��(�����~��X��r���)��=$�ż�B{=VY�=,�
>�;)�Z��m���!4�D���{=	*x=->��
>\��>ƕ]?U&�>蓆>�7?l���Y8�鹮�/?ߺ9=Ҥ��� ������c��C�>��j?���?�\Z?^d>��A�=C��>3=�>E&>5&\>bj�>C��QfE�i�=>��>s�=��M�������	�h����+�<.>���>ʍ|>^m��T(>�����yz�9�d>Y�Q�>���,2T�#�G� �1�D�v�%�>��K?��?�_�=R�&���6f��)?�i<?dM?#�?
��=U�ھ�0:�R�J�/��N�>��<���͒���4���:��a:N9s>aힾ:渾S�>>m�
�]U ��eX���L����'�=o��%=�-�G�ھ�����>��6>�����h��Ɣ�,:���G?��=l򡾫�N��{���7>��>B��>�$������eLA�e���}�=f�>�2>F�K�����.A�5����΁>�[B?�_?m��?�&��j�q���,���u���P��	?Y��>|�?4�g>��= ���b���c��G�Ik�>T��>�����=������A��,��p�>F`?o:">h0?laM??�M?�j?�3�>�|�>��5��	���H&?���?[Ƅ=��Խd�T���8�*F��>��)?c�B��ɗ>�?	�?��&?)yQ?�?m�>G� ��1@�듕>�]�>7�W��`��h`>��J?䖳>�/Y?r̓?�>>��5�����ꩽ��=99>��2?A8#?,�?��>���>vٴ��#
>�)�>�`?�8�?^_{?R�=��>m�>�Y�>�"=_~�>��?�S$?	9T?�#l?/�7?T5�>c��<�����_{�u�m�$2�Rt�;_�3=�7=SØ�엽�O��� �U�<jd=�m���h����8%H�U��;���>�\u>�����*>�8ƾ�І�}d<>�D7��.����� I2���=�7�>�. ?T=�>������=#�>k�>պ�Zx(?�e?ß?�;�_�ùؾj�P�F?�>�DC?a��=��m�蓿�v���=�5n?��^?bN�p�����f?vY?=��t:�A�;l�^�Q����X?y�?o�S���>��?pxt?�e�>�����j�N���w�Y���,����=��>8t�R�j��y�>�a=?��>L�H>���=*��Sw�8���j�?�x�?)��?�'�?Լ6>z�`��ܿ���jߑ�T�k?Z�>�%����-?&\f=цӾ(O�Y6x�(���x3׾�(z�s}�������?��k��z���HC�=g]
?X��?l�n?�U?���:�Z��hV��w�R��	���w�I���=�w�B����7b��rʾ5�˺<]|���E��m�?�)?��#��W�>gqw���󾆀���5H>�rq�'�6����=�0��Q[='�=�]f�MN�_���?k��>҉�>��9?�[�(Z?��E+�/�)�.a߾dY6>d@�>PY>�@�>��ϧe���Ž�qپ������1�,>�m?��d?7�T?�,6�yt�5�Y���C�� ��(��qhk<?��=�O�>�O\�e?u��Y2���X��J������#�޿
�<O�</�U?, >4C�>B�?�~�>�㷾�2ƾ1}�h)�%?}=��?ȉ?T��>�ӡ>������Z��>�2o?e��>�=�>�f�ь�lS[��m��i�>���>4�>��>!s�RU�0ы�fË��1��g�=��g?����V�]�ҍ�>xK?�����@=���>������ �%��|cK��-)>��?Q�.=��(>�M���
��{s�����Jf.?�I?#����{*��e>P�%?���>E�>�	�?\��>����h�i<��?�S?~�H?F+B?f�><�=Cy���ȽD:�uxH=}��>\�K>�pW=�R�=P���U�� �"JG=C�=tؼ��齩��<]��Ae�<�=�'>W�ݿ�ZM��߾F��S��m�R������m�MO'�yR˾���(b������m/�L�D��,N�����{�i����?9��?����;���j���y�5h��D�>�X���ٽD��η��*�r��4ھN쥾gK ��LD��Q`���a�u�?����ȿ�L���莾
�2?*��>f��?�������c=�rU5>b�=�����}ǾH����ƿFy��i??:?n}�N#H�A�?!ƙ>)��>ۊ�=���@?��
�=��#?�/?�>er־�ſ?z��n��=�r�?��@��A?��(�]��(�U=���>��	?�?>�1��7��簾Y�>B<�?W��?�M=��W��	��pe?f�<�F�(:ݻ�>�=�w�=��=���&�J>�R�>Q��FuA���۽��4>C��>�q"����h2^�#�<��]>biս����5Մ?,{\��f���/��T��U>��T?�*�>J:�=��,?X7H�a}Ͽ�\��*a?�0�?���?'�(?3ۿ��ؚ>��ܾ��M?aD6?���>�d&��t�څ�=�6Ἀ���w���&V�t��=Y��>e�>��,������O�J��V��=�n���ſ�! ����1<e:c�w�xc��%Y��!h�Q���BR� g �v��=J >s�`>v��>]�+>�wK>��Z?�t?�ˍ>eW�=�X�fQ��n�Ӿ���=�;i��^g�����s���_��F�D�پ���$�������оB5\�(��<��\�z ��=Ѿ2�U��!F�ȲD?'Í>y�ﾘ�p�if>�����5�sq>u�W�􅅾U�)�|@_�cX�?��V?�_w��z��$�d���.�D�8�s?JL������h楾�^;=��˽|�">ߟ`>{?��ƹ����z�A�x�Z?x*D?ಾ��z�,��
�׽8�<�
D?��#?��>=P�>��K?2���Ǿ�7>�I>v3�>,�?,��>U�Ѿ��<���>D�5?_T�=�X��aG�>��御�\���g�2�b���-����6>�U�G���z�<�{o���N���`?���>�S*�9n���9��ug�;�O�?��?X�u>�Lx?�~W?���=�~龪Z��]����<[K?�|?�T>�r�����hy���D?=�n?UZ!>�^u�������E[���?�)S?�?�&�f�a�Z4��y򾺓%?E\�?M|�N���M��?�����>��>k�>7"}�?��* ?��޾Dm���οЉ��c�?Y�@{� @`l0�@���k~>�M?�Y>&����Bо��=������>n>Q}���p�^:�����Xg?�Jo?x�?�y��.� y=���D5�?/Yz?-����>���>o�5��X8Z��q�>�
u���=iuо�U��ƴ��A�Il��U���e>R�@��+�j�>Kݽf�ֿZǿ3\]�:�Zپ��>7��>�i�U�T��j`��ؑ�VY��9\������N�>��>H����z�{�9t;����/�>T����>��S��!��'�����5<��>2��>겆>�0��m㽾Yř?%]��\>οk���.����X?�c�?!q�?�t?!:<��v��{� C�:'G?��s?�Z?�S%�l&]��_7��k?󎩾N%`��4�<YE���U>�d2?<��>Ɖ,�Ł=r�>�o�>�>G/�tTĿ^_��Q����Ѧ?�~�?��龫,�>`d�?&�*?�������q����+������A?�0>[����!��h=�k����?S�0?F��D�\�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�f6%?�>d����8Ǿ��<���>�(�>*N>`H_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?Ę�>ZN�?PY�=B��> >(ϱ�j�<�\>��=%遽X��>6�P?��>���=�-F��/�KB�M,N�Vv��]�?���>�*e?9_H?H�N>�����G����#�����.���J�db*�����Y�!�0>��F>��>B[L�u�ξ$�9?'%��Eп	N��E�[��f4?�¨���!?X޾eȽuw�<&�P?�S�>I��_̞��&z�*#�UB�?:��?�^?�o߾h��<	�D>m
�>r�v>bW�������[�����>d4?�ƾa~��aG{�~�>�6�?w;�?@�?ѪT��)?aW$����>�X�sD��=��-f���-?���E\�>��>��$������+_�!�>
1�?���?�?!�[?��_��)��T�=��C>�#T?=f!?�ߓ�����
�=a�?�L��d�����cM?+�@�@� c?W,����̿f����E��C���d�n�Œ�=/�O>�Z�Ä�<L�]>��ϼɇg�iн<3_�>�q�>��>��m>:��=�BV>�J{�)M�Z���C���ؿc��x�(��F��й
��엾-~ �9���	� ��6���Ҵ=��=�:[��ݽAƯ<��=�E?��[?�K�?Tʸ>7�ӽI��>=��Ю�<�7B��w/��=>�:?BGe?'R<?|�>eоs�q��܀���`��j�� �s>b��>��>�Q>��> �~=�=<>�2V>��>5X,>�(=�/�=�&ɼX��>,?�>�i�>�u>T�> ��=�X��:��1rZ�����g��Sן?A����-H�V.������Ǿ��={�3?M��=巏�8�̿����a{O?[e���M��V%����='=?�mM?�(X>ܾٝ�Qh��>P5Ͻ���_>��������p2�4�k>?lyk=�6>I�7��fi�]�-��S�{�=�D?�5�1ҽ��}���0�Ԏ�ؤ�>�v�>m�s;{�a�����T�Z��O�B?�?��6gɾ�^��Ծj��>���>�=����H�=>����ۧ�O���x=�� >�?}�G>�	�=%��>�%��w/�r�>PZ>c>I>�A?��%?��f;pYe�Gא�7)�2��>��>�|�>�->tH����=#`�>�ck>>�`��?꽿�N���D>h�6��_��c���m=��ͽ�>nl�=j�̽ -���<�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿj��>� ���������@o�2Ic=��>�L?/���c�S�=��W?�?�6��]��;ȿ��u�'��>�H�?꽕?�m��̚�S@8�0��>İ�?[Q?,]>�ܾ�H�b��>�>??�@N?,��>�3����;�?x�?��? q=5��?�܉?�K>�iM�U+�N���|� �.�0��<��>}��=��=l��p٘�Ll���b��L�D�{t>�I=X�>d�H�ja��D�o;Z�N���ʾ�?�.�>n��>\
�=�6�>w1�>u�>#�>I9�=>ט�am���t�W�K?���?����2n�rY�<���=��^�-&?�H4?�w[���Ͼ֨>Ӻ\?]?�[?�c�>+��8>��#迿$~����<��K>�3�>�H�>�#���EK>��Ծ�5D�p�>"З>k����>ھ�+������B�>�e!?J��>Ϯ=l�2?N�?2Po>�`	?$����=�����s?��4?���>dÎ?:�?���$����L������|qI�f>
t�?0�;?�>>�d��fY��/��Q�n=���Y%�?���?d-1�UoE?%�?��9?�t�>$����=�����k��=��?�!?�����A��N&���>�?H?���>�璽�[սռ����c����?z\?�?&?,��Ea���¾�H�<� ���M���;�@D�O�>��>ƈ��`�=�*>9��=vkm�d=6�v�d<��=΋�><O�==�6�>����-?A1��󙟾�uI=������J�mY>���=8���?�� ����i��������� �� �?��?`�?�Xq���k��4T?�;�?��>��?����;վ}���k����=�:ʾ��>�$�>���=�����>�1{��ˊU<3��I?#�>���>��+?iŅ>QD�>>q���L+����*�˾�}>�G��Z.�M>B�E���#��b佗�����ʾa�j���>5�/��>݃$?�T�>�SC>�b�>m��S�#>&��>7�>5��>��k>�:>��O>}�=o��R?�����'����f���,�A?�Wc? X�>*�V��R���q��g ?���?D�?�<r>h��!+�|Q?� ?��~�K9
?g;=oIT��@�<�ϴ�{��s$��`;�p��>�D۽=!:�^�L��Mi���
?��?A�{�W~ʾ��ڽ!��a	�=�2�?�>.?� ��KM�� e��T���O��r���2�����a�H	`��%����Ҍ���[)����<��%?�?&�w��&,��gDs���F�_�>c��>3�>>y�k>�t���(�?�W���4�����>:�~?�v�>?J?��;?�O?L?���>�E�>g����>���;��>s��>��8?Ǆ,?>�.?�&?��)?_I^>������6׾1�?�3?��? ?$P?F���wԽ����ծy�Chz�Pc�p�=���<��ֽ��q��L=�J>��?H|�l�7��*��d�h>H87?���>��>)u���~�H��<A�>[b
?�ڌ>U-��Kq�����H�>Ɵ�?8���*
=�6+>e��=�{�����c��=IѼTp�=�ad��>�
�<���=g��=Y�":�A�:;��;��<�t�>.�?���>�C�>�@��>� �?��.e�=�Y>*S>\>�Eپ�}���$��i�g��]y>�w�?�z�?r�f=��=���=�|��QU��`�����<��<Σ?J#?;XT?Q��?r�=?lj#?�>%+�aM���^��(����?� ,?���>i��>�ʾ�7�3�+�?�W?�8a�(���;)���¾�սj�>�[/��.~�-���D�d������������?Ծ�?�@A���6�}p�뿘��\���C?��>�[�>��>F�)���g�F!��';>_��>c
R?�t�>O�P?֖{?�mY?nT>�8�����뙿n����$>�>?��?�n�?=�w?u��>7�>@3����Γ�����\���́��e=N�U>ൔ>���>3��>��=��ֽ�c���"@����= �_>���>��>���>�2v>� l<}�I?��>�.��f,��ݦ��-���J�`Pv?~�?b-?�6=(��K�B�~�����>�ǧ?���?��*?��H��Z�=n����{��lno�b�>x�>�n�>��=��:=X�#>0��>?�>���jO��4��-.���?��F?�ϰ=�q��3Ig�46�����ɠ>�rܾ
��\;��$<�+�=W,˾$�'���m|����N[�2憾5B����ʾPc�>�<�8>۟>2ea=rƆ<��=�K�^G�<EM��0��3ܽl�н�tB�ϕ��y�����~'�EY��z��~?�I?�&?�R6?��U>I�>&�`_�>������>��>:I���-ǾF�V������'ھg���(�X��^����>��3�_:>�� >`d�=�`ؼSb�<u�=�=Ә+��k>�>k�>	��=Nx�=��=�u�=�6w?�������,Q�ݫ��:?�8�>Ҍ�=��ƾ�@?��>>�6�������n��(?1��?xW�?a�?��i�Y�>3�쐎�b=�="✽�2>E��=��2�N¹>��J>5��AK������0�?
�@і??ዿ�Ͽ�Z/>�<,>I�>��R���4�L{U���i�;b�r"?��6�5�Ⱦ_s>��=��I���\�J=p�5>Wwt=���]�	Ԙ=���:�Y=U�=�k�>��>>欹=r����=�pU=/:�=FC>GE�~<����M�6=� �=��]>cH >���>��?cs3?�bq?'v�>?���7���=Gƾ�w�>0^�=��>1�=o�P>E��>�6?M<?m"<?���>�6�<>��>�M�>��*��Be��� �����!��>��?z��?Lk�>6u�=D2(��.�}�D����}��>�.?�:?�ֻ>�H��4�n���)��o��$=�D=s_��ы��U��4�4�8�ֽ����>4q	?eH�>{[Q>��>��>���>/�>d���O=g_=��<[�&�8�^;&��<1�+��%ν�m=���=�0[;��9B��CIx�l�(=I�<3�>?��>��"=
��>>�4׾ R$>��w�F���a> �I�4K�9�a�_����;�f?�t��>�f>���VQ��Y?~��=�<U>)�?�o�?_�j>�������&�|�������$��=���>{���Ե@��R���]�l9��~��>��>��>1�l>��+�u?�z=;�J;5����>��K�E��kq�V1���🿙�h��F�Z�D?d9���3�=�4~?q�I?�Ǐ?â�>���=�ؾ��/>la����=��l�p�����1�?d'?hC�>y� �D��B̾K
���ݷ>6;I��O��,�0�M$��Ƿ����>��S�о�!3��f�����ӌB�Nr���>?�O?�?i4b��V��0UO����%���o?�|g?��>!L?B?�,��9x�Ov��Uu�=T�n?���?5=�?�	>ۨ�=/C��9��>�?�ǚ?^ő?@fs?I�X��>���</T*>G����=���=�5�<���=}�?p\
?5��>�������X۾�h���r^�֊=�=��>%o�>��*>+��=��=o�=��[>S��>ص�>Wvv>~�>)�{>|������?[�=-��>��s?f�>���O��%�xQ�=H6
����� l��f<���n=wV>�3I>��/�{,�>;ϿȰ�?�h>�~)����>5`ܾ�*��w�>��M>��	>H�B>�õ>�]�>
�?���>���r2p>F"u>0LԾ�/�=���120�ҿ'�{�;�\aԾ#��>q����@�6E#��V%���G�u�|�{�Ⱦ(yi��ρ�V;�S�>��?����ހ��~�멯�7�#?��h>ªJ?��޾&��rk>@?���>fE������ۍ�~����?���?�;c>��>H�W? �?ܒ1�43� vZ�+�u�m(A�-e�U�`��፿�����
�|��-�_?�x?0yA?�R�<.:z>Q��?��%�Zӏ��)�>�/�'';�@<=w+�>*��%�`���Ӿ��þ�7��HF>��o?;%�?wY?:TV����"�<kq7?�D?�os?�8?v�?��j�J��>���>a��>�?o:?N5a?'=?�a�>co>Ξ彲'������v��� -��AF����@�T=��=kB<��Fr�<?�׽��W��<&<U`�=��R<[Z=�d+>?L>��=zͦ>0�]?p��>4m�>Y�7?(��8�7����/?��:==���g���Ƣ��4�()>��j?�֫?q9Z?f�d>L�A���B�-�>�K�>%�%>�?\>���>�G�wE�}��=ɓ>m;>��=аN��b����	�h4���R�<��>���>�=|>W����
(>zw��AOz���d>zR�ӽ����S���G�
�1��qv��i�>��K?��?EP�=Eh�=|���6f�b*)?:U<?dHM?
�?���=t�۾��9���J��7��*�>	�<$��A���w!���:�� �:��s>����H���t>9`
��$���L�X���T�Ο=�eþ]�q�<���ƾ�~��o�>�!>Gv��đ-�:������ �=?�^>zsʾ�ɸ�/�Ծ�5>޾]>b/�>���}^=F��ͪw��t�>�?a>�$4������1��1��>@�E?!�Q?��y?�>��w�Y���H�d����h�<j� ?G��>g8	?�gE>�}�=J���!�о�R�;-1����>�?��3bg��J��YV�n�%��	c>;��>r� >)�8?�V?�,�>E�L?�K*?!��>=�)>ax�{Ȋ��L/?���?K��q�<�yr|���)���=�<�>�?�R�=�?�?�� ?K?�2X?Ab�>���=����C�>�}l>GPr����>��8?	��>+h?Q^?#��=�=0��ɾm�h��C >m�>Z�5?���>�ȳ>ʇ�>_��>�g��~0�=�4�>�c?�q�?po?r��=��?��.>���>Gԓ=B��>�w�>M�?Z�N?��s?�'J?B��>�ٔ<I!���º���z��Kz��m$;��0<��o=
p�Xe��c!��Q�<&<����v�22׼��4�a���t;*��>s>╾>[/>\Nƾ�튾�eA>&0��@��}�����<� ��=$��>H?[ߕ>�"��x�=>6�>?��>%��G�'?i�?2�?��;Ga��۾_N��ӱ>�`A?�t�=��l�����j�u��j=ݻm?K�^?d�Z�����b?� ^?\f�C=���þ�b��z�-�O?|�
?l�G�p �>��~??�q?���>Lke�on����Bb��j��Ѷ=�R�>�[�e�d��.�>��7?e�>�(c>�'�=�c۾��w�������?9�?���?}��?��)>��n�F�%o��E���^?v�>���Q�"?)>����Ͼ�)��o9����j��`C��^<���]���Z$��у��׽6�=u�?`s?XGq?��_?@� �X�c��^�����XV������E�� E� �C�Ȣn�D�*;���O��K�F=HQ[��C�}_�?N�!?�?�#�>½��v���v얾���=��Ⱦ7���`�>�BL�g4>���<��p��Z��8پ`?Pb�>:ƶ>�,?ܛ��>�*��N�o�:�@'�Y��>3�>���>���>&�� �����>��r����[���ǽ�׆>"�]?�)J?�m?�a�=W/���������Ś��1���>�O�>���>��ži��(R"��8��P��(�OԒ�k~��o����?���>��?K��?q�?J��+��.��ܭS�x��;��>�?e?@�?y�>����U8�����>0k?G�>Ǯ>=��\b#�݄���1	�rb�>���>�"?@�>Ԥ!���X��e��n=���70�l�>�H]?��~��KN��KM>�6I?�����.�����>{X`:|�#�?�(\2��r�=�>?RXq=�&`>����ܶ��Z��[W��{�)?��?�v��/N*�#)|>��!?�U�>�	�>>��?@��>n9¾�?����?��^?[J?�YA?��>�f=�{���ɽv'��+=�,�>�4Z>��k=0��=d!�D�]���:-:=��=�ȼ1����c;T袼�B><G��<0>NaؿR�F����"�\�վ�!	�>�{�l�������Q�m�����ꆾ�g�A'<��B��@�8Zd�l�:��W�?��?�����S������g>���i�f�>̱��[���;���㣽��������5L!��}T���d���j��'?���L�ǿK����Wܾ?�?�H ?��y?��#�"���8��� >��<�1��ω�ԕ����οP�����^?��>������>�o�>AaX>"cq>���P���a��<Z�?��-?���>N�r���ɿ3x��Q�<���?��@iA?M�(�Eu쾘�X=h��>W�	?1V?>y1��#�Ȱ���>$�?}��?�N=�W�(
���e?���;��F��{ϻ	H�=3��=�=B��L_I>Mے>m����@�.�ڽ��5>�%�>�#�l��)`^�iܻ<�S]>�|ս����TՄ?�v\�@f�.�/��S��5X>��T?�/�>3/�=	�,?�4H��|Ͽ~�\�+a?=/�?ԥ�?��(?�ݿ�fٚ>C�ܾO�M?sC6?`��>c&�,�t����=���������^&V�u��=«�>T{>��,����D�O��F�����=�,���zǿ��;�h�=�A�+>{��=4��<�&<�c�>m�>C�ڽ��孾�-Լ�0=RD�>^1?��?d*�>�Ml?ǅ�?}�>s��=9����v���"]=�����`�!�a��=�>��;r�0ބ�w��nI7���7��
��~�*�c$=�nD��Ն���־�.m�/��ĉ?4�I>_Ᾱ�M�=�/��j�?���� =F�W=`��ŀ/�#�t��t�?mH?7M}��B]�vE���e�<��jy-?" ��>�A瘾�\>A�=e��=��>���<���>�1�,�X�"�0?�y?�r��% ���(>�����%=�,?�^ ?y _<m��> #?�e-���ٽ6k]>��6>7A�>C��>c
>��� #۽�<?�|T?8�����+��>�-¾,}�;�]=*X>-B9��Q޼#�V>��<Dp����q�2����<�(W?�>��)���Sc�����^M==Ȱx?��?�*�>.|k?=�B?B��<}d��5�S�9�QLw=�W?�)i?��>m����о\���g�5?أe?.�N>�Oh���龟�.��V�# ?��n?�^?�3��Nq}�o������o6?��v?s^�vs�����;�V�]=�>�[�>���>��9��k�>�>?�#��G������xY4�$Þ?��@���?��;<��:��=�;?q\�>�O��>ƾ�z������x�q=�"�>����ev����R,�f�8?ޠ�?���>$������yQ>���VǴ?�;x?4%�����=�5�h쀿͡�ͦ>�>��f>I /�F��H�5�a���׾�pi��Eཡ~�>{�	@��	��`�>�j!�Szп˚ۿ�ށ���׾(vw�T?��>T�;�sW��卿����|F��ھ��Ľ7�>�U>�P��_Z��-{�X;�7��2�>�u�>׭P�&���`��_aC<`��>��>�y�>��������>c�?�q��ο�,��H��X?	e�?4y�?R�?N�5<?�y�xX~�}�5�z�F?�`s?OXZ?b5��_���,��j?~_��pU`��4��HE��U>�"3?�B�>S�-�m�|=>���>�g>�#/�\�Ŀzٶ�����F��?ۉ�?�o���>v��?us+?�i��7���[����*��+��<A?�2>Ռ���!�F0=�"Ғ�ʼ
?L~0?!{�\.�H�_?�a�=�p���-���ƽ:ۡ>j�0��e\�:K��z��qXe����JAy����?:^�?b�?r��� #�E6%?+�>*���
9Ǿ?�<���>�(�>j*N>4G_�,�u>����:��h	>~��?�~�?Qj?ە�������U>��}?"�>p�?��=3�>.S�=�j��6�)��#>"%�=��4�8I?��M?�(�>���=�8�c�.���F��BR�}��5�C���>b?iTL?b>@綽.5��1!��;̽��1����2A�J+����p�4>��=>gW>��E�;�Ӿ��?Fp�1�ؿ�i��p'��54?5��>�?����t�����;_?"z�>�6��+���%��lB�b��?�G�?;�?��׾+Q̼#>8�>�I�>�Խ[���9�����7>�B?T��D��b�o�x�>���?�@�ծ?mi��	?���P��Sa~����7����=��7?�0���z>���>��=ov�λ��Q�s����>�B�?�{�?��>�l?��o�<�B���1=CM�>Ĝk?�s?�Po�a�m�B>��?&������L��f?	�
@wu@K�^?(��Կ�ơ�1�ؾ������=k(>��a>4~=Y�>����6�t��3��f� >ǋ�>=��>�ۺ>�>���>Ͻ�>Ӆ���"�Xࣿ�i��B@�"��BE��W�)�j 很pb�" �o�׾�ƭ���v����Zc`���߽� ����=�U?�R?�p?ݏ ?odx���>�����z=ћ#�9��=�#�>�b2?��L?�*?Ϯ�=ꨝ�n�d�N_��A��Aև����>�wI>ԇ�>}Y�>z$�>��9��I>L?>�|�>�>�&=��亶�=��N>�L�>D��>�r�>�:Y>-m->>>��|�����b�⓾��o�Al�?���tq<�����f��	�����K>z�%?�`�=����h̿�ڬ�
,??V��nU�p:�d8=<g?�NU?D9W>����_�� ��=����n$�f�=dbͽi�W���)�f�S>�z+?�>�>[/�>ۿ;�jE��-K���Ӿi�>��B?̩����uw��D<�����xֻ>nM�>�,�����Xڔ�$�~�<�N��?<՛?�	?n�H������N+��d�b�>h��>��^&�=P�>6TֽfꐽC"��[�@>��>��?�(>S�=��>Ǘ�*NT��>�E>�)->�??�X#?��'��������,�y>��>!�>$�>!�F�VZ�=���>Sd>�$��-��le��iB�
�[>c�|�C�^��>���=D���׏�=���=fx���F�Q=�~?}��-䈿��f��nlD?i+?��=�F<V�"�C ���H��;�?n�@�l�?��	��V���?�@�?P�����=�|�>c׫>'ξ��L��?�Ž\Ǣ�m�	�o)#�RS�?��?��/�5ʋ��l�.5>_%?دӾPh�>{x��Z�������u�u�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?V>��?���?S��>;�ս�Z$���ǿ�旿�T�;��>�`�>nC�>�f��38:�,R�+G��þ%HN>A�=3��>yS������>^?��.��B=�J�>&&>y"z>Q�Y>,��>Y��>4�j>�2�=Q����0g�+�����K?5�?���<p�"��<℈=m�W�Ǌ?�M3?�/<�FpҾ�}�>��[?Y��?��X?�j�>�o�A���C(������]<?Y?>��>�V�>�ҏ�LHM>��Ⱦ�C��I�>a�>�M���Ӿb}��G#�Õ�>Q8 ?^�>��=�f ?$? �o>>8�>��D�^����_H�郻>��>2a?zA�?H!?�;��BI2�ƒ�@�<�X�؏P>�w?=�?�З>&����<��)8d��	l�Ґ�4T�?�Me?��� ?w�?�X=?ۑ??��j>����Jپ0ȴ���>�<?#�=}Q��:��}K���?
?cX'?*l��������=j��5��i�?4�y?��0?TI��k�`j���y�<X��3��l?�=34�<��J>���>�<CK޼��>Z'ýD�޾���\�=����s�>�)�=���
�,=,?]�G�}ۃ���=��r�?xD���>�IL>����^?ol=��{�����x��	U� �?���?Yk�?r��;�h��$=?�?T	?o"�>�J���}޾7�ྯPw�~x��w�J�>���>��l���F���ڙ���F��s�Ž����(��>�E�>˱D?H�?��>m]�>�n¾AZ>�Aj�� ھ��b�>��1�u��s`�ϊ�7�L��"��{2r=ղ��h��G��>o#�=H{ ?50? &d>��\>F0 ?�0;��)>eN>9�>�!>�!H>2����-�>۲2>@>�HR?������'���0Ұ�6�A?�jd?���>Yi�zm��y��
_?ׁ�?���?= v>S|h��*+��/?��>Q���@
?�8=�"�q߁<Pr���2�����?��Eێ>x�׽�:���L���f��b
?�&?�r��IL̾_FԽ걙���r=ю�?��'?1/��lK�M�t�g�\��U��\1�,�O�0��W?!���o����Y���.���"�^��<�'?Qa�?�j�������xj�'H��qP>U��>��> �>��e>!_�>!*���f���,�u�r����>�r|?��>�I?�<?�P?�fL?w׎>@�>���<4�>���;n�>���>x�9?T�-?�0?G`?cm+?!Hc>����s����ؾ��?��?e?=?��?����.�½�꙼��h�[�y������݁=��<l�׽f=t�K#V=�MT>�V?���u�8�K���Yk>i|7?1��>���>��g/����<L�>Q�
?�M�>(���xyr��^�V�>���?5���Q=��)>��=���C\Ӻfh�=�������=~���;���<�s�=���=vGv��i�L��:S��;uܮ<Zs�>��?�>�H�>�J���� �H���
�=��X>�7S>�0>�%پ�y��n"���g��%y>Nv�?�x�?��f=~�=|��=~��=L��
��+��qe�<�?�I#?�VT?ۙ�?�=?8g#?��>�1�)M��+[������ű?�](?�j�>����ξPܳ��/[�$"?�?rW���d>��L��x�0v>r�>�6��HN�����)2����=��.�ֽ�1�?hP�?�&����W�0���v����\?��>�'�>�V?��I���"��B��A�=�:�>�P?Rz�>�+O?�}~?G�\?(�6>�y8�ݶ���$���M�=�9>��L?];�?��?�k?��>���=�s��ľ\c���m��ɽ]���v6=QP>V�r>]��>���>b�=�x��и�1lb��$�=^I>�v�>^c�>"{�>/e9>���7h�G?K��>�^�����b뤾�ă�l�<��u?%��?Đ+?{W=���E��D��$K�>�n�?���?�2*?S�S����=��ּ�ᶾI�q��$�>�ٹ>T2�>տ�=�uF=�a>|�>���>�(��`�gq8��>M���?	F?ģ�=%���5?e�'����	3=�ꧾTA�1+뼘�a�J.=������,$¾^��뤾�s���y���i�X o���?�l=FL>��>ݶ�<9S���2=G��=�V=xN�;����N=@����=5��\ �;ᴟ<�=����-z˾ti}?0HI?1�+?��C?Bz>dB>�)3�ë�>�}��:,?y�U>3UQ�䢼��5;�|�������ؾ�y׾��c�bԟ��^>}YI�ȟ>~3>:#�=���<#%�=�\s=���=�A���=:P�=u�=���=��=��>�Z>5w?4���g����3Q��L罳�:?�9�>���=�~ƾ@?E�>>y2�������a��,?	��?'T�?��?wi��e�>6��_掽�t�=۱��V;2>���=��2���>��J>q���J��w��33�?L�@Y�??I⋿=�ϿS]/>Z�=��=��A�q�7�R뺽�!���b��a)?( ��Ҿ��6>
��=2e��iH��+��FK>�>��G=M&H���>Ù����=�l7>�>f
>�|>�#e�(,R>�$,=��6���=��L��[���<�P&>���=˫�=�t����>�?�'?B4g?�j�>D
�sVھ�Oƾ�#�>�y�=#��>��=�a�>�y�>#�&?�/?�"]?Z�>�$ =���>���>�$��R����7i�
���9�f?��x?���>�K>UpB�ϯ#��P��`�����>Ւ?�8�>�ۥ>������XdB�M�3�#xM=^�">�	>_s����=A]���E�v�A����=���>�r�>
�?d�>�e�>���>���>ګ�=ϿQ�1�u�^�!J��D���偼�o�=� >>�50=���ڟ� ���98=�b<��=N_V=���=���>ѯ>���>N��=�ͳ�0/>�Ȗ�"�L�|�=�o���1B���c��P~���.��j6���B>��W>8��]&��H�?�UZ>@>���?�[u?�r >���-վ�Y��.e�5�S��X�=�->��<��s;��`�W�M��>Ҿe��>�	�>�`�>�r8>"8M�*�C��U�=����$��|*?�u̾Y�$�@�?>�O�zU��z����i�
_)���?d3~����<��?��<?�M�??#��2S�ev�>��H�R=LL3����"?��?��?H.?R���_W��H̾���޷>�@I�!�O���P�0�9��Eͷ���>������оg$3��g�������B��Lr�m��>�O?��?J:b��W��+UO����E(���q?�|g?4�>�J?�@?�%��z�_r��}v�=��n?���?P=�?R>�֫={����>>�A?�Ӟ?��?*ZL?Fq���׼>�	��Dl=<���[>q����	>��t=�� ?�i�>�\�>����Y���:�&ꁾi�n����<��>�Ұ>��>ʲ=X�=,�x>!u�>��>ѿ�>c��>8$>�	>���3��Fq:?��3>˓�>H'?�=�>';�<č�=>��@���*l��p�E��g�;؆���5�R�j=�k����>����ʑ?�i�>I[���?�Ծ�R3=�>�G*=���#�>���^>+��>5,�>U��=1v�>uߧ=f5Ӿu�>���k!��*C���R�ƭѾ��z>t���u�%�֣��{��a$I��F��	c��
j��,��f>=���<<D�?����;�k�K�)������?Z_�>�6?�ތ�q҈�}�>��>�Ӎ>�I��񊕿�Í��jᾗ�?f��?�7c>��>[�W?Ś?�1��3�qZ�ȫu��%A��e�X�`����������
������_?s�x?wvA? �<*;z>8��?��%�(Ώ��*�>�/�q$;��<=�-�>i&��l�`��Ӿ��þ@��GF>1�o?�"�?gS?�RV�"t���>�7@?j�1?u�u?#�1?Ǥ9?�w�U�(?��>Ba?�N?^W,?g�(?^�?��'>� �=6�G��<�9���͊��B���i�mg�ڽ^=��$= 2�����p<=�_e<���:>T!�.b�;=ƾ����<9�?=h�=E�=�Ŧ>1�]?�X�>�>��7?| �7Y8�񮾃�.?;�7=۳���>��<����p�u�>��j?^�?�IZ?�d>4�A��$C��L>hY�>{�&>�@\>8�>~����D�;.�=b�>�t>��=|�N�`���\�	� ��5��<i>��?J��>��㽳F@>{s��� ���>����h�J�ko8���U��K�'ps>�?\�5?N���i��8$���;Y��b�>��p?U�h?�|?�oa>�Ҿ
�\��M4�����>7IԽSR��ݮ�����X(���;ꖦ>M��?̍�k�z>�������=�d�9NO��vܾ>?�=@����=��p[Ӿ�:q����=�>}þ�"�́��"	��׹E?�b=����G�������=�U�>'s�>}A޽/�<�{4������=�R�>|�6>����'=־g�A���a�>"�D??mM?1	t?�@����O��='�����Ϊ�XEw=۳�>�h�>�<�>СG>��6<Z�;i�ɾ�V��<�V��>\�?�)��y�x`�����/��*>}g�>P�+>�'?�yj?R�>�}?$h?�<�>�/�>���3��C'?�΃?�f=D�ཤ�Z��\8���B����>$(?Y�H�� �>�?8�?V�)?kAN?,�?�x>�G�Q�@���>���>�Y�������^>1	G?��>�[?p�? >��1��⢾�,����=��>U8?>/?��?D�>|��>�����=0?��?�^�?h�~?h6e=��?��=~�>Yzq<�	�>nT�>	�>�oa??g�?�nS?],?`�*�^�����>�>�|ڼ���֋<5п���t�1��<#�D>�Z>D�<Rٽ��w=��_�+;�/�;4��>�mm>�j��֥+>M߾�[���'*;>K���B晾�ω�6�=����=R�>� ?_@�>b���@�=��>�H�>g��ݹ&?��?�1?N�;2__�A�׾��G����>,�=?�e�=��m�-��Wpt����=
tn?��]?H4_�����-Gb?�b?��;�9���̾{�p���۾ܸF?8?�yE�L�>�r?Ķ\?��?u!h��f�4��ۇb�'�w�m��=	�>�o �ql�[�>�E%?�W�>,��>�!>���j��㜾��>�S�?�?�?c�?`�=�6l�I�㿠w��rF��
^?j�>�����"?D��Ͼ�����x-�'��*���X��R���$��냾�ֽ7��=��?�s?KKq?��_?'� ���c��=^�� ���TV���� ���E��"E�C� �n�)k��:���7���G=��[�� >�}�?wM?���}H�>5$������u����J>� ޾�W�J%�D�i��{>yNQ�ǰ��Gc�����~�?'�>�D�>7n�>tl���8�;!X�E�+�e��T�>���>�i�>�>��=P��������j�ʜW�f���vde>�8U?��J?B�h?�[��)��r�w�1`)�����\@�wV�>�H>�S�>iن�6[��,}3�����M��2Ӿv㐾����L����B?�}�>�y�>�{�?w:?B��K��h� ��`b��� ��H#>���?�0?'�Q>lҚ�b8¾���>�l?�z�>u��>$!��x(!���|��ѽ���>���>�=?�:v>"(���Z���ⷎ�38�"��=�{g?Vt��WN`���>��Q?���;�t<��>U�q���!�2��n(��>Q�?���=�+=>-�þ�N�>�{�����ִ-?��?6���M'���h>��?Z��>��>��?�@y>�-��cb!��c?��^?�G?(&D?�.�>bZ�<Li���ž�U�1�Q�=^x�>0�F>( �=�A�=a����X�/���w�<(γ=�X���:�?o�<٫$���<xk�<'�;>Q�ؿDSK���ݾz����辋b�ᬎ�Q[���X�E8�oȺ�.ۓ���~��O�U��x)G��u^��҇�R�a�oJ�?�2�?Q����
������W���j��º>9R�S�������c�]R���iԾ������$���W���m�6z`�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >`C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾�1�<��?7�-?��>Ďr�1�ɿc����¤<���?0�@pZA?'�(�$2�+�\=!�>�	?�o@>�)1�q� ���A�>��?M�?�7G=9�W����C�e?�~<wF�L�껗l�=�q�=c�=C��6�K>p�>����A�q!ݽ��4>ie�>��$����eL_����<�^>��ҽ�t��5Մ?({\��f���/��T��U>��T?+�>]:�=��,?X7H�`}Ͽ�\��*a?�0�?���?#�(?;ۿ��ؚ>��ܾ��M?bD6?���>�d&��t�ޅ�=u6�牤�x���&V�~��=\��>Q�>,�ދ���O� J��i��=���O��2
A��F��=u�7<�n����,�Z�->	����C��
����j��
>�� >0�>7r>ᆓ>��>�%g?*�}?3*�>'�/;�k �4���-���W�=�)_�bc��}Xվ�t���2����F�0���ھ�*��F���
��= C�R���e����]Y�:�M�3�?��>�"ܾ�Y��T��e��m=�HM�<kܼ�����H��]��,�?�D?�z�q�g��<��� n�L|<�u;? ﱾ#V��N��9N=wmB��Ӧ=mI�>fV;f)���T��d�%4?�\?���F@���>�2��	�=��6?q�?�*���M�>�F?D)!�p���`>Gg>	ʛ>	K�>ź�=?Ӳ�|�⽗;)?��Z?��ཞ������>Ïž�o��X�=Z�=�./��y;;Zk>$�L��׈�3x+=��P�.�=l(W?��>n�)����`������Y==Ͳx?��?�-�>B{k?��B?�ڤ<�h����S����fw= �W?S*i?i�>_����	о]��� �5?��e?��N>Uah����3�.�yU�G$?��n?�^?	x��w}�U��l���n6?��v?s^�Ws��N����V�1>�>\�>���>��9�k�>ؑ>?�#��G��
����Y4�
Þ?��@|��?��;<�����=�;?�[�>'�O�O>ƾ�z��ۂ���q=["�>0���sev����LR,�[�8?���?p��>
���p��&��=圾KI�?��{?�����:������g������Ya=,E�:�C�<�:ӽ����^-��߾��������th�0B�>��@�&�SF�>�F��(տQ�Կ̀��.cᾂp۽;�?T��>2X��qR���u�߂z�S����4�!<���G�>"e3>������� 4y��/9��LX����>�|��-}> �`��J��9#���.a=ؔ�>�"�>9'�>~P齪¾dj�?���'�ͿG���9�ͨL?H��?�]�?KY!?�'{�jh��L����J�K?�m?'-f?����_5n�Z��%�j?�_��xU`��4�uHE��U>�"3?�B�>T�-�^�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*��+��<A?�2>���I�!�C0=�VҒ���
?W~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�>��?-��=���>ܕ�=f̴��a!�7>���=�|�$�?�L?F��>_��=�u4��z/�yCF���R���wC�_Q�>�2d?��L?��e>Yr��6��"�Ҵ½�V5��ּb�?��YV�����}:>Jc?>�>�J@�|zо�?�<�>7׿�閿-���0?8K}>�� ?�Y���u�n����~`?��>��(���jo��DI�q��?���?H
?fξ��R�}�>�}�>%��>H⽋����φ�=�.>VeC?���±��Ul�l9�>���?�H@
��?��m��	?���P��Va~����7�`��=��7?�0��z>���>��=�nv�ݻ��X�s����>�B�?�{�?��>"�l?��o�N�B���1=8M�>͜k?�s?Ro���h�B>��?"������L��f?�
@u@_�^?*�忄P��Co��%�ɾ�]>�IN>F�,>��H��؂>d�=N'>�|P�x��=�}�>���>���>m��>{��>ٳ�>*^��n�$��<��	H����8��	�I���Wɾ���?�	��������8)¾ґ�T� =�0�!v��۽T�Ǽ��=�U?)�Q?c�o?&0 ?�}���>����*��<V>"�y{�=��>jX2?u�L?�*?4]�=�ӝ���d��S���X���߇��N�>�J>���>���>F��>Qہ�PNJ>�O>>���>�� >]t!=iJ%��=�O>��>8
�>It�>�5]>�W\>� ���O��҈R����۽�T�?�����0A��5����{�1'���d�=��#?��=֭��k�̿�D���B?�n���f�H����=o�	?ǻg?kUZ>�{�٩P=�t>\-�leڽd�>oR���}=��h��4>�"�>Φ�>��>j�:��;�xeU�#%���>��1?���	gn<`cE�	.>�`v���>*N�>�G�{������@���zg�HFt��V^?�&/?qS���ו��D�1ľ�(P>p*�>�ӌ���=�}k>�];�b������Ǎ=��Z=���> �?~�,>Q�=���>-���e+L�Y��>(D>{->��>?�X#?i.�W�7*��v�+���w>"��>H�~>�	>��I����=l5�>��`>�H�O���n��B�rV>Үu�2\�Ӑu�6gt=�?���`�=�̑=�G���:��G&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�g�>�x��Z�����}�u�s�#=��>�8H?<V����O�">�w
??�^�詤���ȿ9|v����>L�?���?
�m�kA���@����>��?[gY?�ni>�g۾q`Z����>�@?�R?*�>�9�Î'���?�޶?���?�e>�q�?�0�?�Ө>�$���"�ݨǿu���2i�5ڒ>��>���>�9�"s5��G��!��� 9N�s�}�/]=�U{=d��>�����J|�;���-T����Ľ]�>!Q>��>졝>�0?�>٢�>	{��q揽������F��L?�|�?[���n�6Q�<�0�=Y�Z��&?�{2?�֌��ξ��>�[?�<�?��Z?Д>������I����"�����<�zL>
y�>��>����N>��Ӿ�G�V��>b��>*���>־����अ� r�>��!?B�>�د=~ ?t'$? �i>�r�>orE��_��q�D�Gþ>���>-\?�|?N(?H���s?1�H���ࡡ���X�0&I>�w?Ɋ?���>�ď�mp��K�j��q�ju���΁?9f?ul뽓�?�'�?U�=?�NC?��c>�[�׾@���as>��:?�)>=qX���fQ��>D?f8?���=���8r<���k$���J?��-?*�V?�`��b��-�&�S=�J+��£�xTP=w\<��%>`�>�aw����=�\=��=w'�������7>uي>�=닂��E��0=,?��G�~ۃ���=��r�>xD���>�IL>����^?ll=��{�����x��	U� �? ��?Zk�?`��?�h��$=?�?S	?l"�>�J���}޾6�྿Pw�~x��w�Z�>���>�l���K���ڙ���F��`�Ž�*�6x�>�>�>�?x��>��>}��>���������'G�%o������<�;��j�u���?(�L�=o���8m�f�>��`���>���>L�>X4�>�I�>�����ep>�:>�_P>�ۢ>�(8>XA\>� �=-_�<��ý�KR?���z�'�������3B?%qd?m0�>�i���������?���?�r�?P>v>�~h�,+�zm?F>�>����p
?�H:=:$��;�<�T��-��n)�������>WL׽�!:��M��lf��j
?�0?+���̾<׽� ����=A�?�??:*��L�i~{��Z��O����<yс��RN���#�SKl�XY������z���b_��n&?D��?ܽ �^�����{z]� �S�dj3>ul�>b��>W3�>�$>�+۾]&��a�D&�7V1�N��>��f?�Ѝ>�`I?+�;?��P?%�K?�ߏ>��>�\�����>|�;��>.6�>�O9?�,?�.?�?"S,?�>b>���g���16ؾ��?�	?��?��?�?����g���@y��zB=�e|�黄��;�=��<�7ܽ�]��Vh=T�U>�X?����8�����P k>ŀ7?8��>���>`��
0��}��<��>��
?XE�>s���fzr��b��R�>e��?���k|=�)>���=(����Ӻ�X�=���n�={9��3�;��0<���=�=xkt���|����:G�;Ax�<_i�>c�?߭�>�K�>�R��� ����='�X>�@S>��>O3پkv�����u�g��y>�o�?4o�?2�f=�H�=�/�=����i�����O���r�<ϊ?<3#?bT?G��?*�=?�s#?|�> -��I��M���󢾽�?�N*?E
�>`���;j�����:���?���>	�d�)(Ƚи&��A��A4���Z'>��(��?}�������G�xӳ��_�Ѳ��NF�?��?}�0���*��P�:虿�e����<?U�>ip�>i6�>e(�I\��>�Q�*>[��>
�Q?��>fN?7I�?C�??x��$+���������1~��ȸ>((�?n~�?���?Y�c?�k�=��(�C�Ž�eҽH��3Β�l�׽�=��7>�a�>���>��?M��>dω��a����a���s=��H>(��>�
�>$��>A��T�O>�G?'%�>Ǿ�H��.Ѥ�l킾��5�yu?tu�?��*?t8=,c�]E�X��^Y�>HQ�?�?�)?\�R��(�=��ּ�����n�eٸ>���>�>~ҍ=�B=�>z�>��>�����}�8��UV���?yF?�5�=�2��7o��������ĺ-=����4�`��Bl�_E$�7��=;ǳ�
L���*|��@��^��l���˾ɉ��=�k�?��=gS>g>3�y=h��������:��9jғ;8q�����=4�%��h�;n��o�E=��=~:/=�*��q�˾(�}?l;I?��+?�C?��y>�=>5�3�w��>\����>?�V>ܬP�9���V�;�㪨�� ���ؾ�t׾��c��ȟ�uG>�bI�b�>A53>ML�=,R�<	�=Js=���=�R�E=�&�=L�=n�=l��=��>�S>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��H>��>ǔT���0�h�]���e�#�I��$?�C6��Ծ���>wx�=�$�����O=��D>9=V�$���]�쑛=�����W=.�=���>rT@>ۮ�=˵��0��=��e=K7�=1�G>���;�H����	��Q=a��=��]>VD%>��>i?�/?�uf?@�>�>B��ƾ����^!w>qF�=��>�'0=�9>�k�>��:?{�9?PWH?�7�>O��=��>I�>�>,�C�]�@�޾�Y�����=j��?$��?A!�>��I�-����$��;�k��?	�%?CX�>���>��ɸ忲�/��g,��b��R�=��,=�獾�|a��
�:���{w �!��=b��>;s�>�(�>��>��>�}�>��>��>�"�<>�b=�ߝ<�5=�.���o�=Q���B~=�J<*$��JS��\�<Yʊ<
q#��փ<�:;,^�=(|�>Ӡ>a��>R��=����.>FҖ��L��N�=执��A��c�K2~���-�7/8��-C>�V>J�{��ԑ��?�=W>`�B>���?Z2u?	�%>���оw]���k�"�[���==�>�59�y�9��:`��N��7оۇ�>!l|>}�>�Q1>��4�3>N����=���#C��~
?tS������?���?���{�w��{f����J�?��~����zn�?��Q?�"�?9�?y�Ǽ���;-�>.�þ��<�����ʖh�uX(?J(?��>W�v��73��3̾B��<
�>�:I�	P�����S�0��9!�u׷����>8�����о3��b��Q�����B�53r����>��O?��?�a�R���JO����l#���I?.bg?	�>a?[V?����11�R����=[�n?!��?2:�?j�
>�>��콡f�>�b?"s�?�̣?�~m?d��=�&�>�W��A�=�ʏ�v�R>�Ꞿ�x�Rk>�R?�J)?��H?^��ԉ��y��Aҧ�k�c>�<�=Eg?��>��9=�1Ӽgؽ�轣d�=�ry>��J>j��=���>P��>�0�� D�p�B?�=>]�>� ?�S�>�����Tő=F(۽S����ɷ������=���H���36=)*���>�k¿�i�?�K>�S��y�?����l�=��>�2�=�FC�j	�>��A>��F=��>�:�>=��=��>F>�FӾO~>���We!�U,C�G�R���Ѿv}z>���>	&���Uu���AI� n��Hg�=j�c.��+<=��ǽ<H�?p�����k���)�"���c�?v[�>P6?>܌����ذ>��>ɍ>�I��B���ȍ�g�;�?a��?�b>~1�>��W?;�?Y�1�e�0�Y���t���@��sd�'�`�����r���
��:���Q_?xex?��@?�X�<��z>��?m�%��2����>Gn/�@�:�)!4=��>⯾9k_�M�ѾF�¾R����C>��n?�%�?C�?JW��m�l'>h�:?��1?�Pt?H�1?�;?_��R�$?n3>�E?�p?�N5?^�.?��
?1
2>|�=k���z�'=47����ѽ�}ʽ���j�3=�P{=�i˸I�
<
�=q�<�c��sټ�l;�Y��'�<�:=��=��=(�>��Y?���>���>�{/?杽u��y���:�&?�����*�#����O��u
��~=a�^?TJ�?��K?��r>WLQ��pG��/8>i$�>+Qt>�>b�>�'6���G��`�=}LZ>?��=W�A=zr?;� �����&��8;>ВB>t�?Oɐ>^�Qi[>�����WC��>^?���ቾE��L���%��p@���N>)L9?�t+?��=N:���>�<�`�S�?&�M?&]?}?��,>�޵�,�L���=�K����̢>r�ƻ�����������<�<�9>_��>]�B��H���t>9`
��$���L�X���T�Ο=�eþ]�q�<���ƾ�~��o�>�!>Gv��đ-�:������ �=?�^>zsʾ�ɸ�/�Ծ�5>޾]>b/�>���}^=F��ͪw��t�>�?a>�$4������1��1��>@�E?!�Q?��y?�>��w�Y���H�d����h�<j� ?G��>g8	?�gE>�}�=J���!�о�R�;-1����>�?��3bg��J��YV�n�%��	c>;��>r� >)�8?�V?�,�>E�L?�K*?!��>=�)>ax�{Ȋ��L/?���?K��q�<�yr|���)���=�<�>�?�R�=�?�?�� ?K?�2X?Ab�>���=����C�>�}l>GPr����>��8?	��>+h?Q^?#��=�=0��ɾm�h��C >m�>Z�5?���>�ȳ>ʇ�>_��>�g��~0�=�4�>�c?�q�?po?r��=��?��.>���>Gԓ=B��>�w�>M�?Z�N?��s?�'J?B��>�ٔ<I!���º���z��Kz��m$;��0<��o=
p�Xe��c!��Q�<&<����v�22׼��4�a���t;*��>s>╾>[/>\Nƾ�튾�eA>&0��@��}�����<� ��=$��>H?[ߕ>�"��x�=>6�>?��>%��G�'?i�?2�?��;Ga��۾_N��ӱ>�`A?�t�=��l�����j�u��j=ݻm?K�^?d�Z�����b?� ^?\f�C=���þ�b��z�-�O?|�
?l�G�p �>��~??�q?���>Lke�on����Bb��j��Ѷ=�R�>�[�e�d��.�>��7?e�>�(c>�'�=�c۾��w�������?9�?���?}��?��)>��n�F�%o��E���^?v�>���Q�"?)>����Ͼ�)��o9����j��`C��^<���]���Z$��у��׽6�=u�?`s?XGq?��_?@� �X�c��^�����XV������E�� E� �C�Ȣn�D�*;���O��K�F=HQ[��C�}_�?N�!?�?�#�>½��v���v얾���=��Ⱦ7���`�>�BL�g4>���<��p��Z��8پ`?Pb�>:ƶ>�,?ܛ��>�*��N�o�:�@'�Y��>3�>���>���>&�� �����>��r����[���ǽ�׆>"�]?�)J?�m?�a�=W/���������Ś��1���>�O�>���>��ži��(R"��8��P��(�OԒ�k~��o����?���>��?K��?q�?J��+��.��ܭS�x��;��>�?e?@�?y�>����U8�����>0k?G�>Ǯ>=��\b#�݄���1	�rb�>���>�"?@�>Ԥ!���X��e��n=���70�l�>�H]?��~��KN��KM>�6I?�����.�����>{X`:|�#�?�(\2��r�=�>?RXq=�&`>����ܶ��Z��[W��{�)?��?�v��/N*�#)|>��!?�U�>�	�>>��?@��>n9¾�?����?��^?[J?�YA?��>�f=�{���ɽv'��+=�,�>�4Z>��k=0��=d!�D�]���:-:=��=�ȼ1����c;T袼�B><G��<0>NaؿR�F����"�\�վ�!	�>�{�l�������Q�m�����ꆾ�g�A'<��B��@�8Zd�l�:��W�?��?�����S������g>���i�f�>̱��[���;���㣽��������5L!��}T���d���j��'?���L�ǿK����Wܾ?�?�H ?��y?��#�"���8��� >��<�1��ω�ԕ����οP�����^?��>������>�o�>AaX>"cq>���P���a��<Z�?��-?���>N�r���ɿ3x��Q�<���?��@iA?M�(�Eu쾘�X=h��>W�	?1V?>y1��#�Ȱ���>$�?}��?�N=�W�(
���e?���;��F��{ϻ	H�=3��=�=B��L_I>Mے>m����@�.�ڽ��5>�%�>�#�l��)`^�iܻ<�S]>�|ս����TՄ?�v\�@f�.�/��S��5X>��T?�/�>3/�=	�,?�4H��|Ͽ~�\�+a?=/�?ԥ�?��(?�ݿ�fٚ>C�ܾO�M?sC6?`��>c&�,�t����=���������^&V�u��=«�>T{>��,����D�O��F�����=�,���zǿ��;�h�=�A�+>{��=4��<�&<�c�>m�>C�ڽ��孾�-Լ�0=RD�>^1?��?d*�>�Ml?ǅ�?}�>s��=9����v���"]=�����`�!�a��=�>��;r�0ބ�w��nI7���7��
��~�*�c$=�nD��Ն���־�.m�/��ĉ?4�I>_Ᾱ�M�=�/��j�?���� =F�W=`��ŀ/�#�t��t�?mH?7M}��B]�vE���e�<��jy-?" ��>�A瘾�\>A�=e��=��>���<���>�1�,�X�"�0?�y?�r��% ���(>�����%=�,?�^ ?y _<m��> #?�e-���ٽ6k]>��6>7A�>C��>c
>��� #۽�<?�|T?8�����+��>�-¾,}�;�]=*X>-B9��Q޼#�V>��<Dp����q�2����<�(W?�>��)���Sc�����^M==Ȱx?��?�*�>.|k?=�B?B��<}d��5�S�9�QLw=�W?�)i?��>m����о\���g�5?أe?.�N>�Oh���龟�.��V�# ?��n?�^?�3��Nq}�o������o6?��v?s^�vs�����;�V�]=�>�[�>���>��9��k�>�>?�#��G������xY4�$Þ?��@���?��;<��:��=�;?q\�>�O��>ƾ�z������x�q=�"�>����ev����R,�f�8?ޠ�?���>$������yQ>���VǴ?�;x?4%�����=�5�h쀿͡�ͦ>�>��f>I /�F��H�5�a���׾�pi��Eཡ~�>{�	@��	��`�>�j!�Szп˚ۿ�ށ���׾(vw�T?��>T�;�sW��卿����|F��ھ��Ľ7�>�U>�P��_Z��-{�X;�7��2�>�u�>׭P�&���`��_aC<`��>��>�y�>��������>c�?�q��ο�,��H��X?	e�?4y�?R�?N�5<?�y�xX~�}�5�z�F?�`s?OXZ?b5��_���,��j?~_��pU`��4��HE��U>�"3?�B�>S�-�m�|=>���>�g>�#/�\�Ŀzٶ�����F��?ۉ�?�o���>v��?us+?�i��7���[����*��+��<A?�2>Ռ���!�F0=�"Ғ�ʼ
?L~0?!{�\.�H�_?�a�=�p���-���ƽ:ۡ>j�0��e\�:K��z��qXe����JAy����?:^�?b�?r��� #�E6%?+�>*���
9Ǿ?�<���>�(�>j*N>4G_�,�u>����:��h	>~��?�~�?Qj?ە�������U>��}?"�>p�?��=3�>.S�=�j��6�)��#>"%�=��4�8I?��M?�(�>���=�8�c�.���F��BR�}��5�C���>b?iTL?b>@綽.5��1!��;̽��1����2A�J+����p�4>��=>gW>��E�;�Ӿ��?Fp�1�ؿ�i��p'��54?5��>�?����t�����;_?"z�>�6��+���%��lB�b��?�G�?;�?��׾+Q̼#>8�>�I�>�Խ[���9�����7>�B?T��D��b�o�x�>���?�@�ծ?mi��	?���P��Sa~����7����=��7?�0���z>���>��=ov�λ��Q�s����>�B�?�{�?��>�l?��o�<�B���1=CM�>Ĝk?�s?�Po�a�m�B>��?&������L��f?	�
@wu@K�^?(��Կ�ơ�1�ؾ������=k(>��a>4~=Y�>����6�t��3��f� >ǋ�>=��>�ۺ>�>���>Ͻ�>Ӆ���"�Xࣿ�i��B@�"��BE��W�)�j 很pb�" �o�׾�ƭ���v����Zc`���߽� ����=�U?�R?�p?ݏ ?odx���>�����z=ћ#�9��=�#�>�b2?��L?�*?Ϯ�=ꨝ�n�d�N_��A��Aև����>�wI>ԇ�>}Y�>z$�>��9��I>L?>�|�>�>�&=��亶�=��N>�L�>D��>�r�>�:Y>-m->>>��|�����b�⓾��o�Al�?���tq<�����f��	�����K>z�%?�`�=����h̿�ڬ�
,??V��nU�p:�d8=<g?�NU?D9W>����_�� ��=����n$�f�=dbͽi�W���)�f�S>�z+?�>�>[/�>ۿ;�jE��-K���Ӿi�>��B?̩����uw��D<�����xֻ>nM�>�,�����Xڔ�$�~�<�N��?<՛?�	?n�H������N+��d�b�>h��>��^&�=P�>6TֽfꐽC"��[�@>��>��?�(>S�=��>Ǘ�*NT��>�E>�)->�??�X#?��'��������,�y>��>!�>$�>!�F�VZ�=���>Sd>�$��-��le��iB�
�[>c�|�C�^��>���=D���׏�=���=fx���F�Q=�~?}��-䈿��f��nlD?i+?��=�F<V�"�C ���H��;�?n�@�l�?��	��V���?�@�?P�����=�|�>c׫>'ξ��L��?�Ž\Ǣ�m�	�o)#�RS�?��?��/�5ʋ��l�.5>_%?دӾPh�>{x��Z�������u�u�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?V>��?���?S��>;�ս�Z$���ǿ�旿�T�;��>�`�>nC�>�f��38:�,R�+G��þ%HN>A�=3��>yS������>^?��.��B=�J�>&&>y"z>Q�Y>,��>Y��>4�j>�2�=Q����0g�+�����K?5�?���<p�"��<℈=m�W�Ǌ?�M3?�/<�FpҾ�}�>��[?Y��?��X?�j�>�o�A���C(������]<?Y?>��>�V�>�ҏ�LHM>��Ⱦ�C��I�>a�>�M���Ӿb}��G#�Õ�>Q8 ?^�>��=�f ?$? �o>>8�>��D�^����_H�郻>��>2a?zA�?H!?�;��BI2�ƒ�@�<�X�؏P>�w?=�?�З>&����<��)8d��	l�Ґ�4T�?�Me?��� ?w�?�X=?ۑ??��j>����Jپ0ȴ���>�<?#�=}Q��:��}K���?
?cX'?*l��������=j��5��i�?4�y?��0?TI��k�`j���y�<X��3��l?�=34�<��J>���>�<CK޼��>Z'ýD�޾���\�=����s�>�)�=���
�,=,?]�G�}ۃ���=��r�?xD���>�IL>����^?ol=��{�����x��	U� �?���?Yk�?r��;�h��$=?�?T	?o"�>�J���}޾7�ྯPw�~x��w�J�>���>��l���F���ڙ���F��s�Ž����(��>�E�>˱D?H�?��>m]�>�n¾AZ>�Aj�� ھ��b�>��1�u��s`�ϊ�7�L��"��{2r=ղ��h��G��>o#�=H{ ?50? &d>��\>F0 ?�0;��)>eN>9�>�!>�!H>2����-�>۲2>@>�HR?������'���0Ұ�6�A?�jd?���>Yi�zm��y��
_?ׁ�?���?= v>S|h��*+��/?��>Q���@
?�8=�"�q߁<Pr���2�����?��Eێ>x�׽�:���L���f��b
?�&?�r��IL̾_FԽ걙���r=ю�?��'?1/��lK�M�t�g�\��U��\1�,�O�0��W?!���o����Y���.���"�^��<�'?Qa�?�j�������xj�'H��qP>U��>��> �>��e>!_�>!*���f���,�u�r����>�r|?��>�I?�<?�P?�fL?w׎>@�>���<4�>���;n�>���>x�9?T�-?�0?G`?cm+?!Hc>����s����ؾ��?��?e?=?��?����.�½�꙼��h�[�y������݁=��<l�׽f=t�K#V=�MT>�V?���u�8�K���Yk>i|7?1��>���>��g/����<L�>Q�
?�M�>(���xyr��^�V�>���?5���Q=��)>��=���C\Ӻfh�=�������=~���;���<�s�=���=vGv��i�L��:S��;uܮ<Zs�>��?�>�H�>�J���� �H���
�=��X>�7S>�0>�%پ�y��n"���g��%y>Nv�?�x�?��f=~�=|��=~��=L��
��+��qe�<�?�I#?�VT?ۙ�?�=?8g#?��>�1�)M��+[������ű?�](?�j�>����ξPܳ��/[�$"?�?rW���d>��L��x�0v>r�>�6��HN�����)2����=��.�ֽ�1�?hP�?�&����W�0���v����\?��>�'�>�V?��I���"��B��A�=�:�>�P?Rz�>�+O?�}~?G�\?(�6>�y8�ݶ���$���M�=�9>��L?];�?��?�k?��>���=�s��ľ\c���m��ɽ]���v6=QP>V�r>]��>���>b�=�x��и�1lb��$�=^I>�v�>^c�>"{�>/e9>���7h�G?K��>�^�����b뤾�ă�l�<��u?%��?Đ+?{W=���E��D��$K�>�n�?���?�2*?S�S����=��ּ�ᶾI�q��$�>�ٹ>T2�>տ�=�uF=�a>|�>���>�(��`�gq8��>M���?	F?ģ�=%���5?e�'����	3=�ꧾTA�1+뼘�a�J.=������,$¾^��뤾�s���y���i�X o���?�l=FL>��>ݶ�<9S���2=G��=�V=xN�;����N=@����=5��\ �;ᴟ<�=����-z˾ti}?0HI?1�+?��C?Bz>dB>�)3�ë�>�}��:,?y�U>3UQ�䢼��5;�|�������ؾ�y׾��c�bԟ��^>}YI�ȟ>~3>:#�=���<#%�=�\s=���=�A���=:P�=u�=���=��=��>�Z>5w?4���g����3Q��L罳�:?�9�>���=�~ƾ@?E�>>y2�������a��,?	��?'T�?��?wi��e�>6��_掽�t�=۱��V;2>���=��2���>��J>q���J��w��33�?L�@Y�??I⋿=�ϿS]/>Z�=��=��A�q�7�R뺽�!���b��a)?( ��Ҿ��6>
��=2e��iH��+��FK>�>��G=M&H���>Ù����=�l7>�>f
>�|>�#e�(,R>�$,=��6���=��L��[���<�P&>���=˫�=�t����>�?�'?B4g?�j�>D
�sVھ�Oƾ�#�>�y�=#��>��=�a�>�y�>#�&?�/?�"]?Z�>�$ =���>���>�$��R����7i�
���9�f?��x?���>�K>UpB�ϯ#��P��`�����>Ւ?�8�>�ۥ>������XdB�M�3�#xM=^�">�	>_s����=A]���E�v�A����=���>�r�>
�?d�>�e�>���>���>ګ�=ϿQ�1�u�^�!J��D���偼�o�=� >>�50=���ڟ� ���98=�b<��=N_V=���=���>ѯ>���>N��=�ͳ�0/>�Ȗ�"�L�|�=�o���1B���c��P~���.��j6���B>��W>8��]&��H�?�UZ>@>���?�[u?�r >���-վ�Y��.e�5�S��X�=�->��<��s;��`�W�M��>Ҿe��>�	�>�`�>�r8>"8M�*�C��U�=����$��|*?�u̾Y�$�@�?>�O�zU��z����i�
_)���?d3~����<��?��<?�M�??#��2S�ev�>��H�R=LL3����"?��?��?H.?R���_W��H̾���޷>�@I�!�O���P�0�9��Eͷ���>������оg$3��g�������B��Lr�m��>�O?��?J:b��W��+UO����E(���q?�|g?4�>�J?�@?�%��z�_r��}v�=��n?���?P=�?R>�֫={����>>�A?�Ӟ?��?*ZL?Fq���׼>�	��Dl=<���[>q����	>��t=�� ?�i�>�\�>����Y���:�&ꁾi�n����<��>�Ұ>��>ʲ=X�=,�x>!u�>��>ѿ�>c��>8$>�	>���3��Fq:?��3>˓�>H'?�=�>';�<č�=>��@���*l��p�E��g�;؆���5�R�j=�k����>����ʑ?�i�>I[���?�Ծ�R3=�>�G*=���#�>���^>+��>5,�>U��=1v�>uߧ=f5Ӿu�>���k!��*C���R�ƭѾ��z>t���u�%�֣��{��a$I��F��	c��
j��,��f>=���<<D�?����;�k�K�)������?Z_�>�6?�ތ�q҈�}�>��>�Ӎ>�I��񊕿�Í��jᾗ�?f��?�7c>��>[�W?Ś?�1��3�qZ�ȫu��%A��e�X�`����������
������_?s�x?wvA? �<*;z>8��?��%�(Ώ��*�>�/�q$;��<=�-�>i&��l�`��Ӿ��þ@��GF>1�o?�"�?gS?�RV�"t���>�7@?j�1?u�u?#�1?Ǥ9?�w�U�(?��>Ba?�N?^W,?g�(?^�?��'>� �=6�G��<�9���͊��B���i�mg�ڽ^=��$= 2�����p<=�_e<���:>T!�.b�;=ƾ����<9�?=h�=E�=�Ŧ>1�]?�X�>�>��7?| �7Y8�񮾃�.?;�7=۳���>��<����p�u�>��j?^�?�IZ?�d>4�A��$C��L>hY�>{�&>�@\>8�>~����D�;.�=b�>�t>��=|�N�`���\�	� ��5��<i>��?J��>��㽳F@>{s��� ���>����h�J�ko8���U��K�'ps>�?\�5?N���i��8$���;Y��b�>��p?U�h?�|?�oa>�Ҿ
�\��M4�����>7IԽSR��ݮ�����X(���;ꖦ>M���H���t>9`
��$���L�X���T�Ο=�eþ]�q�<���ƾ�~��o�>�!>Gv��đ-�:������ �=?�^>zsʾ�ɸ�/�Ծ�5>޾]>b/�>���}^=F��ͪw��t�>�?a>�$4������1��1��>@�E?!�Q?��y?�>��w�Y���H�d����h�<j� ?G��>g8	?�gE>�}�=J���!�о�R�;-1����>�?��3bg��J��YV�n�%��	c>;��>r� >)�8?�V?�,�>E�L?�K*?!��>=�)>ax�{Ȋ��L/?���?K��q�<�yr|���)���=�<�>�?�R�=�?�?�� ?K?�2X?Ab�>���=����C�>�}l>GPr����>��8?	��>+h?Q^?#��=�=0��ɾm�h��C >m�>Z�5?���>�ȳ>ʇ�>_��>�g��~0�=�4�>�c?�q�?po?r��=��?��.>���>Gԓ=B��>�w�>M�?Z�N?��s?�'J?B��>�ٔ<I!���º���z��Kz��m$;��0<��o=
p�Xe��c!��Q�<&<����v�22׼��4�a���t;*��>s>╾>[/>\Nƾ�튾�eA>&0��@��}�����<� ��=$��>H?[ߕ>�"��x�=>6�>?��>%��G�'?i�?2�?��;Ga��۾_N��ӱ>�`A?�t�=��l�����j�u��j=ݻm?K�^?d�Z�����b?� ^?\f�C=���þ�b��z�-�O?|�
?l�G�p �>��~??�q?���>Lke�on����Bb��j��Ѷ=�R�>�[�e�d��.�>��7?e�>�(c>�'�=�c۾��w�������?9�?���?}��?��)>��n�F�%o��E���^?v�>���Q�"?)>����Ͼ�)��o9����j��`C��^<���]���Z$��у��׽6�=u�?`s?XGq?��_?@� �X�c��^�����XV������E�� E� �C�Ȣn�D�*;���O��K�F=HQ[��C�}_�?N�!?�?�#�>½��v���v얾���=��Ⱦ7���`�>�BL�g4>���<��p��Z��8پ`?Pb�>:ƶ>�,?ܛ��>�*��N�o�:�@'�Y��>3�>���>���>&�� �����>��r����[���ǽ�׆>"�]?�)J?�m?�a�=W/���������Ś��1���>�O�>���>��ži��(R"��8��P��(�OԒ�k~��o����?���>��?K��?q�?J��+��.��ܭS�x��;��>�?e?@�?y�>����U8�����>0k?G�>Ǯ>=��\b#�݄���1	�rb�>���>�"?@�>Ԥ!���X��e��n=���70�l�>�H]?��~��KN��KM>�6I?�����.�����>{X`:|�#�?�(\2��r�=�>?RXq=�&`>����ܶ��Z��[W��{�)?��?�v��/N*�#)|>��!?�U�>�	�>>��?@��>n9¾�?����?��^?[J?�YA?��>�f=�{���ɽv'��+=�,�>�4Z>��k=0��=d!�D�]���:-:=��=�ȼ1����c;T袼�B><G��<0>NaؿR�F����"�\�վ�!	�>�{�l�������Q�m�����ꆾ�g�A'<��B��@�8Zd�l�:��W�?��?�����S������g>���i�f�>̱��[���;���㣽��������5L!��}T���d���j��'?���L�ǿK����Wܾ?�?�H ?��y?��#�"���8��� >��<�1��ω�ԕ����οP�����^?��>������>�o�>AaX>"cq>���P���a��<Z�?��-?���>N�r���ɿ3x��Q�<���?��@iA?M�(�Eu쾘�X=h��>W�	?1V?>y1��#�Ȱ���>$�?}��?�N=�W�(
���e?���;��F��{ϻ	H�=3��=�=B��L_I>Mے>m����@�.�ڽ��5>�%�>�#�l��)`^�iܻ<�S]>�|ս����TՄ?�v\�@f�.�/��S��5X>��T?�/�>3/�=	�,?�4H��|Ͽ~�\�+a?=/�?ԥ�?��(?�ݿ�fٚ>C�ܾO�M?sC6?`��>c&�,�t����=���������^&V�u��=«�>T{>��,����D�O��F�����=�,���zǿ��;�h�=�A�+>{��=4��<�&<�c�>m�>C�ڽ��孾�-Լ�0=RD�>^1?��?d*�>�Ml?ǅ�?}�>s��=9����v���"]=�����`�!�a��=�>��;r�0ބ�w��nI7���7��
��~�*�c$=�nD��Ն���־�.m�/��ĉ?4�I>_Ᾱ�M�=�/��j�?���� =F�W=`��ŀ/�#�t��t�?mH?7M}��B]�vE���e�<��jy-?" ��>�A瘾�\>A�=e��=��>���<���>�1�,�X�"�0?�y?�r��% ���(>�����%=�,?�^ ?y _<m��> #?�e-���ٽ6k]>��6>7A�>C��>c
>��� #۽�<?�|T?8�����+��>�-¾,}�;�]=*X>-B9��Q޼#�V>��<Dp����q�2����<�(W?�>��)���Sc�����^M==Ȱx?��?�*�>.|k?=�B?B��<}d��5�S�9�QLw=�W?�)i?��>m����о\���g�5?أe?.�N>�Oh���龟�.��V�# ?��n?�^?�3��Nq}�o������o6?��v?s^�vs�����;�V�]=�>�[�>���>��9��k�>�>?�#��G������xY4�$Þ?��@���?��;<��:��=�;?q\�>�O��>ƾ�z������x�q=�"�>����ev����R,�f�8?ޠ�?���>$������yQ>���VǴ?�;x?4%�����=�5�h쀿͡�ͦ>�>��f>I /�F��H�5�a���׾�pi��Eཡ~�>{�	@��	��`�>�j!�Szп˚ۿ�ށ���׾(vw�T?��>T�;�sW��卿����|F��ھ��Ľ7�>�U>�P��_Z��-{�X;�7��2�>�u�>׭P�&���`��_aC<`��>��>�y�>��������>c�?�q��ο�,��H��X?	e�?4y�?R�?N�5<?�y�xX~�}�5�z�F?�`s?OXZ?b5��_���,��j?~_��pU`��4��HE��U>�"3?�B�>S�-�m�|=>���>�g>�#/�\�Ŀzٶ�����F��?ۉ�?�o���>v��?us+?�i��7���[����*��+��<A?�2>Ռ���!�F0=�"Ғ�ʼ
?L~0?!{�\.�H�_?�a�=�p���-���ƽ:ۡ>j�0��e\�:K��z��qXe����JAy����?:^�?b�?r��� #�E6%?+�>*���
9Ǿ?�<���>�(�>j*N>4G_�,�u>����:��h	>~��?�~�?Qj?ە�������U>��}?"�>p�?��=3�>.S�=�j��6�)��#>"%�=��4�8I?��M?�(�>���=�8�c�.���F��BR�}��5�C���>b?iTL?b>@綽.5��1!��;̽��1����2A�J+����p�4>��=>gW>��E�;�Ӿ��?Fp�1�ؿ�i��p'��54?5��>�?����t�����;_?"z�>�6��+���%��lB�b��?�G�?;�?��׾+Q̼#>8�>�I�>�Խ[���9�����7>�B?T��D��b�o�x�>���?�@�ծ?mi��	?���P��Sa~����7����=��7?�0���z>���>��=ov�λ��Q�s����>�B�?�{�?��>�l?��o�<�B���1=CM�>Ĝk?�s?�Po�a�m�B>��?&������L��f?	�
@wu@K�^?(��Կ�ơ�1�ؾ������=k(>��a>4~=Y�>����6�t��3��f� >ǋ�>=��>�ۺ>�>���>Ͻ�>Ӆ���"�Xࣿ�i��B@�"��BE��W�)�j 很pb�" �o�׾�ƭ���v����Zc`���߽� ����=�U?�R?�p?ݏ ?odx���>�����z=ћ#�9��=�#�>�b2?��L?�*?Ϯ�=ꨝ�n�d�N_��A��Aև����>�wI>ԇ�>}Y�>z$�>��9��I>L?>�|�>�>�&=��亶�=��N>�L�>D��>�r�>�:Y>-m->>>��|�����b�⓾��o�Al�?���tq<�����f��	�����K>z�%?�`�=����h̿�ڬ�
,??V��nU�p:�d8=<g?�NU?D9W>����_�� ��=����n$�f�=dbͽi�W���)�f�S>�z+?�>�>[/�>ۿ;�jE��-K���Ӿi�>��B?̩����uw��D<�����xֻ>nM�>�,�����Xڔ�$�~�<�N��?<՛?�	?n�H������N+��d�b�>h��>��^&�=P�>6TֽfꐽC"��[�@>��>��?�(>S�=��>Ǘ�*NT��>�E>�)->�??�X#?��'��������,�y>��>!�>$�>!�F�VZ�=���>Sd>�$��-��le��iB�
�[>c�|�C�^��>���=D���׏�=���=fx���F�Q=�~?}��-䈿��f��nlD?i+?��=�F<V�"�C ���H��;�?n�@�l�?��	��V���?�@�?P�����=�|�>c׫>'ξ��L��?�Ž\Ǣ�m�	�o)#�RS�?��?��/�5ʋ��l�.5>_%?دӾPh�>{x��Z�������u�u�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?V>��?���?S��>;�ս�Z$���ǿ�旿�T�;��>�`�>nC�>�f��38:�,R�+G��þ%HN>A�=3��>yS������>^?��.��B=�J�>&&>y"z>Q�Y>,��>Y��>4�j>�2�=Q����0g�+�����K?5�?���<p�"��<℈=m�W�Ǌ?�M3?�/<�FpҾ�}�>��[?Y��?��X?�j�>�o�A���C(������]<?Y?>��>�V�>�ҏ�LHM>��Ⱦ�C��I�>a�>�M���Ӿb}��G#�Õ�>Q8 ?^�>��=�f ?$? �o>>8�>��D�^����_H�郻>��>2a?zA�?H!?�;��BI2�ƒ�@�<�X�؏P>�w?=�?�З>&����<��)8d��	l�Ґ�4T�?�Me?��� ?w�?�X=?ۑ??��j>����Jپ0ȴ���>�<?#�=}Q��:��}K���?
?cX'?*l��������=j��5��i�?4�y?��0?TI��k�`j���y�<X��3��l?�=34�<��J>���>�<CK޼��>Z'ýD�޾���\�=����s�>�)�=���
�,=,?]�G�}ۃ���=��r�?xD���>�IL>����^?ol=��{�����x��	U� �?���?Yk�?r��;�h��$=?�?T	?o"�>�J���}޾7�ྯPw�~x��w�J�>���>��l���F���ڙ���F��s�Ž����(��>�E�>˱D?H�?��>m]�>�n¾AZ>�Aj�� ھ��b�>��1�u��s`�ϊ�7�L��"��{2r=ղ��h��G��>o#�=H{ ?50? &d>��\>F0 ?�0;��)>eN>9�>�!>�!H>2����-�>۲2>@>�HR?������'���0Ұ�6�A?�jd?���>Yi�zm��y��
_?ׁ�?���?= v>S|h��*+��/?��>Q���@
?�8=�"�q߁<Pr���2�����?��Eێ>x�׽�:���L���f��b
?�&?�r��IL̾_FԽ걙���r=ю�?��'?1/��lK�M�t�g�\��U��\1�,�O�0��W?!���o����Y���.���"�^��<�'?Qa�?�j�������xj�'H��qP>U��>��> �>��e>!_�>!*���f���,�u�r����>�r|?��>�I?�<?�P?�fL?w׎>@�>���<4�>���;n�>���>x�9?T�-?�0?G`?cm+?!Hc>����s����ؾ��?��?e?=?��?����.�½�꙼��h�[�y������݁=��<l�׽f=t�K#V=�MT>�V?���u�8�K���Yk>i|7?1��>���>��g/����<L�>Q�
?�M�>(���xyr��^�V�>���?5���Q=��)>��=���C\Ӻfh�=�������=~���;���<�s�=���=vGv��i�L��:S��;uܮ<Zs�>��?�>�H�>�J���� �H���
�=��X>�7S>�0>�%پ�y��n"���g��%y>Nv�?�x�?��f=~�=|��=~��=L��
��+��qe�<�?�I#?�VT?ۙ�?�=?8g#?��>�1�)M��+[������ű?�](?�j�>����ξPܳ��/[�$"?�?rW���d>��L��x�0v>r�>�6��HN�����)2����=��.�ֽ�1�?hP�?�&����W�0���v����\?��>�'�>�V?��I���"��B��A�=�:�>�P?Rz�>�+O?�}~?G�\?(�6>�y8�ݶ���$���M�=�9>��L?];�?��?�k?��>���=�s��ľ\c���m��ɽ]���v6=QP>V�r>]��>���>b�=�x��и�1lb��$�=^I>�v�>^c�>"{�>/e9>���7h�G?K��>�^�����b뤾�ă�l�<��u?%��?Đ+?{W=���E��D��$K�>�n�?���?�2*?S�S����=��ּ�ᶾI�q��$�>�ٹ>T2�>տ�=�uF=�a>|�>���>�(��`�gq8��>M���?	F?ģ�=%���5?e�'����	3=�ꧾTA�1+뼘�a�J.=������,$¾^��뤾�s���y���i�X o���?�l=FL>��>ݶ�<9S���2=G��=�V=xN�;����N=@����=5��\ �;ᴟ<�=����-z˾ti}?0HI?1�+?��C?Bz>dB>�)3�ë�>�}��:,?y�U>3UQ�䢼��5;�|�������ؾ�y׾��c�bԟ��^>}YI�ȟ>~3>:#�=���<#%�=�\s=���=�A���=:P�=u�=���=��=��>�Z>5w?4���g����3Q��L罳�:?�9�>���=�~ƾ@?E�>>y2�������a��,?	��?'T�?��?wi��e�>6��_掽�t�=۱��V;2>���=��2���>��J>q���J��w��33�?L�@Y�??I⋿=�ϿS]/>Z�=��=��A�q�7�R뺽�!���b��a)?( ��Ҿ��6>
��=2e��iH��+��FK>�>��G=M&H���>Ù����=�l7>�>f
>�|>�#e�(,R>�$,=��6���=��L��[���<�P&>���=˫�=�t����>�?�'?B4g?�j�>D
�sVھ�Oƾ�#�>�y�=#��>��=�a�>�y�>#�&?�/?�"]?Z�>�$ =���>���>�$��R����7i�
���9�f?��x?���>�K>UpB�ϯ#��P��`�����>Ւ?�8�>�ۥ>������XdB�M�3�#xM=^�">�	>_s����=A]���E�v�A����=���>�r�>
�?d�>�e�>���>���>ګ�=ϿQ�1�u�^�!J��D���偼�o�=� >>�50=���ڟ� ���98=�b<��=N_V=���=���>ѯ>���>N��=�ͳ�0/>�Ȗ�"�L�|�=�o���1B���c��P~���.��j6���B>��W>8��]&��H�?�UZ>@>���?�[u?�r >���-վ�Y��.e�5�S��X�=�->��<��s;��`�W�M��>Ҿe��>�	�>�`�>�r8>"8M�*�C��U�=����$��|*?�u̾Y�$�@�?>�O�zU��z����i�
_)���?d3~����<��?��<?�M�??#��2S�ev�>��H�R=LL3����"?��?��?H.?R���_W��H̾���޷>�@I�!�O���P�0�9��Eͷ���>������оg$3��g�������B��Lr�m��>�O?��?J:b��W��+UO����E(���q?�|g?4�>�J?�@?�%��z�_r��}v�=��n?���?P=�?R>�֫={����>>�A?�Ӟ?��?*ZL?Fq���׼>�	��Dl=<���[>q����	>��t=�� ?�i�>�\�>����Y���:�&ꁾi�n����<��>�Ұ>��>ʲ=X�=,�x>!u�>��>ѿ�>c��>8$>�	>���3��Fq:?��3>˓�>H'?�=�>';�<č�=>��@���*l��p�E��g�;؆���5�R�j=�k����>����ʑ?�i�>I[���?�Ծ�R3=�>�G*=���#�>���^>+��>5,�>U��=1v�>uߧ=f5Ӿu�>���k!��*C���R�ƭѾ��z>t���u�%�֣��{��a$I��F��	c��
j��,��f>=���<<D�?����;�k�K�)������?Z_�>�6?�ތ�q҈�}�>��>�Ӎ>�I��񊕿�Í��jᾗ�?f��?�7c>��>[�W?Ś?�1��3�qZ�ȫu��%A��e�X�`����������
������_?s�x?wvA? �<*;z>8��?��%�(Ώ��*�>�/�q$;��<=�-�>i&��l�`��Ӿ��þ@��GF>1�o?�"�?gS?�RV�"t���>�7@?j�1?u�u?#�1?Ǥ9?�w�U�(?��>Ba?�N?^W,?g�(?^�?��'>� �=6�G��<�9���͊��B���i�mg�ڽ^=��$= 2�����p<=�_e<���:>T!�.b�;=ƾ����<9�?=h�=E�=�Ŧ>1�]?�X�>�>��7?| �7Y8�񮾃�.?;�7=۳���>��<����p�u�>��j?^�?�IZ?�d>4�A��$C��L>hY�>{�&>�@\>8�>~����D�;.�=b�>�t>��=|�N�`���\�	� ��5��<i>��?J��>��㽳F@>{s��� ���>����h�J�ko8���U��K�'ps>�?\�5?N���i��8$���;Y��b�>��p?U�h?�|?�oa>�Ҿ
�\��M4�����>7IԽSR��ݮ�����X(���;ꖦ>M��?̍�k�z>�������=�d�9NO��vܾ>?�=@����=��p[Ӿ�:q����=�>}þ�"�́��"	��׹E?�b=����G�������=�U�>'s�>}A޽/�<�{4������=�R�>|�6>����'=־g�A���a�>"�D??mM?1	t?�@����O��='�����Ϊ�XEw=۳�>�h�>�<�>СG>��6<Z�;i�ɾ�V��<�V��>\�?�)��y�x`�����/��*>}g�>P�+>�'?�yj?R�>�}?$h?�<�>�/�>���3��C'?�΃?�f=D�ཤ�Z��\8���B����>$(?Y�H�� �>�?8�?V�)?kAN?,�?�x>�G�Q�@���>���>�Y�������^>1	G?��>�[?p�? >��1��⢾�,����=��>U8?>/?��?D�>|��>�����=0?��?�^�?h�~?h6e=��?��=~�>Yzq<�	�>nT�>	�>�oa??g�?�nS?],?`�*�^�����>�>�|ڼ���֋<5п���t�1��<#�D>�Z>D�<Rٽ��w=��_�+;�/�;4��>�mm>�j��֥+>M߾�[���'*;>K���B晾�ω�6�=����=R�>� ?_@�>b���@�=��>�H�>g��ݹ&?��?�1?N�;2__�A�׾��G����>,�=?�e�=��m�-��Wpt����=
tn?��]?H4_�����-Gb?�b?��;�9���̾{�p���۾ܸF?8?�yE�L�>�r?Ķ\?��?u!h��f�4��ۇb�'�w�m��=	�>�o �ql�[�>�E%?�W�>,��>�!>���j��㜾��>�S�?�?�?c�?`�=�6l�I�㿠w��rF��
^?j�>�����"?D��Ͼ�����x-�'��*���X��R���$��냾�ֽ7��=��?�s?KKq?��_?'� ���c��=^�� ���TV���� ���E��"E�C� �n�)k��:���7���G=��[�� >�}�?wM?���}H�>5$������u����J>� ޾�W�J%�D�i��{>yNQ�ǰ��Gc�����~�?'�>�D�>7n�>tl���8�;!X�E�+�e��T�>���>�i�>�>��=P��������j�ʜW�f���vde>�8U?��J?B�h?�[��)��r�w�1`)�����\@�wV�>�H>�S�>iن�6[��,}3�����M��2Ӿv㐾����L����B?�}�>�y�>�{�?w:?B��K��h� ��`b��� ��H#>���?�0?'�Q>lҚ�b8¾���>�l?�z�>u��>$!��x(!���|��ѽ���>���>�=?�:v>"(���Z���ⷎ�38�"��=�{g?Vt��WN`���>��Q?���;�t<��>U�q���!�2��n(��>Q�?���=�+=>-�þ�N�>�{�����ִ-?��?6���M'���h>��?Z��>��>��?�@y>�-��cb!��c?��^?�G?(&D?�.�>bZ�<Li���ž�U�1�Q�=^x�>0�F>( �=�A�=a����X�/���w�<(γ=�X���:�?o�<٫$���<xk�<'�;>Q�ؿDSK���ݾz����辋b�ᬎ�Q[���X�E8�oȺ�.ۓ���~��O�U��x)G��u^��҇�R�a�oJ�?�2�?Q����
������W���j��º>9R�S�������c�]R���iԾ������$���W���m�6z`�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >`C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾�1�<��?7�-?��>Ďr�1�ɿc����¤<���?0�@pZA?'�(�$2�+�\=!�>�	?�o@>�)1�q� ���A�>��?M�?�7G=9�W����C�e?�~<wF�L�껗l�=�q�=c�=C��6�K>p�>����A�q!ݽ��4>ie�>��$����eL_����<�^>��ҽ�t��5Մ?({\��f���/��T��U>��T?+�>]:�=��,?X7H�`}Ͽ�\��*a?�0�?���?#�(?;ۿ��ؚ>��ܾ��M?bD6?���>�d&��t�ޅ�=u6�牤�x���&V�~��=\��>Q�>,�ދ���O� J��i��=���O��2
A��F��=u�7<�n����,�Z�->	����C��
����j��
>�� >0�>7r>ᆓ>��>�%g?*�}?3*�>'�/;�k �4���-���W�=�)_�bc��}Xվ�t���2����F�0���ھ�*��F���
��= C�R���e����]Y�:�M�3�?��>�"ܾ�Y��T��e��m=�HM�<kܼ�����H��]��,�?�D?�z�q�g��<��� n�L|<�u;? ﱾ#V��N��9N=wmB��Ӧ=mI�>fV;f)���T��d�%4?�\?���F@���>�2��	�=��6?q�?�*���M�>�F?D)!�p���`>Gg>	ʛ>	K�>ź�=?Ӳ�|�⽗;)?��Z?��ཞ������>Ïž�o��X�=Z�=�./��y;;Zk>$�L��׈�3x+=��P�.�=l(W?��>n�)����`������Y==Ͳx?��?�-�>B{k?��B?�ڤ<�h����S����fw= �W?S*i?i�>_����	о]��� �5?��e?��N>Uah����3�.�yU�G$?��n?�^?	x��w}�U��l���n6?��v?s^�Ws��N����V�1>�>\�>���>��9�k�>ؑ>?�#��G��
����Y4�
Þ?��@|��?��;<�����=�;?�[�>'�O�O>ƾ�z��ۂ���q=["�>0���sev����LR,�[�8?���?p��>
���p��&��=圾KI�?��{?�����:������g������Ya=,E�:�C�<�:ӽ����^-��߾��������th�0B�>��@�&�SF�>�F��(տQ�Կ̀��.cᾂp۽;�?T��>2X��qR���u�߂z�S����4�!<���G�>"e3>������� 4y��/9��LX����>�|��-}> �`��J��9#���.a=ؔ�>�"�>9'�>~P齪¾dj�?���'�ͿG���9�ͨL?H��?�]�?KY!?�'{�jh��L����J�K?�m?'-f?����_5n�Z��%�j?�_��xU`��4�uHE��U>�"3?�B�>T�-�^�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*��+��<A?�2>���I�!�C0=�VҒ���
?W~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>gH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�>��?-��=���>ܕ�=f̴��a!�7>���=�|�$�?�L?F��>_��=�u4��z/�yCF���R���wC�_Q�>�2d?��L?��e>Yr��6��"�Ҵ½�V5��ּb�?��YV�����}:>Jc?>�>�J@�|zо�?�<�>7׿�閿-���0?8K}>�� ?�Y���u�n����~`?��>��(���jo��DI�q��?���?H
?fξ��R�}�>�}�>%��>H⽋����φ�=�.>VeC?���±��Ul�l9�>���?�H@
��?��m��	?���P��Va~����7�`��=��7?�0��z>���>��=�nv�ݻ��X�s����>�B�?�{�?��>"�l?��o�N�B���1=8M�>͜k?�s?Ro���h�B>��?"������L��f?�
@u@_�^?*�忄P��Co��%�ɾ�]>�IN>F�,>��H��؂>d�=N'>�|P�x��=�}�>���>���>m��>{��>ٳ�>*^��n�$��<��	H����8��	�I���Wɾ���?�	��������8)¾ґ�T� =�0�!v��۽T�Ǽ��=�U?)�Q?c�o?&0 ?�}���>����*��<V>"�y{�=��>jX2?u�L?�*?4]�=�ӝ���d��S���X���߇��N�>�J>���>���>F��>Qہ�PNJ>�O>>���>�� >]t!=iJ%��=�O>��>8
�>It�>�5]>�W\>� ���O��҈R����۽�T�?�����0A��5����{�1'���d�=��#?��=֭��k�̿�D���B?�n���f�H����=o�	?ǻg?kUZ>�{�٩P=�t>\-�leڽd�>oR���}=��h��4>�"�>Φ�>��>j�:��;�xeU�#%���>��1?���	gn<`cE�	.>�`v���>*N�>�G�{������@���zg�HFt��V^?�&/?qS���ו��D�1ľ�(P>p*�>�ӌ���=�}k>�];�b������Ǎ=��Z=���> �?~�,>Q�=���>-���e+L�Y��>(D>{->��>?�X#?i.�W�7*��v�+���w>"��>H�~>�	>��I����=l5�>��`>�H�O���n��B�rV>Үu�2\�Ӑu�6gt=�?���`�=�̑=�G���:��G&=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�g�>�x��Z�����}�u�s�#=��>�8H?<V����O�">�w
??�^�詤���ȿ9|v����>L�?���?
�m�kA���@����>��?[gY?�ni>�g۾q`Z����>�@?�R?*�>�9�Î'���?�޶?���?�e>�q�?�0�?�Ө>�$���"�ݨǿu���2i�5ڒ>��>���>�9�"s5��G��!��� 9N�s�}�/]=�U{=d��>�����J|�;���-T����Ľ]�>!Q>��>졝>�0?�>٢�>	{��q揽������F��L?�|�?[���n�6Q�<�0�=Y�Z��&?�{2?�֌��ξ��>�[?�<�?��Z?Д>������I����"�����<�zL>
y�>��>����N>��Ӿ�G�V��>b��>*���>־����अ� r�>��!?B�>�د=~ ?t'$? �i>�r�>orE��_��q�D�Gþ>���>-\?�|?N(?H���s?1�H���ࡡ���X�0&I>�w?Ɋ?���>�ď�mp��K�j��q�ju���΁?9f?ul뽓�?�'�?U�=?�NC?��c>�[�׾@���as>��:?�)>=qX���fQ��>D?f8?���=���8r<���k$���J?��-?*�V?�`��b��-�&�S=�J+��£�xTP=w\<��%>`�>�aw����=�\=��=w'�������7>uي>�=닂��E��0=,?��G�~ۃ���=��r�>xD���>�IL>����^?ll=��{�����x��	U� �? ��?Zk�?`��?�h��$=?�?S	?l"�>�J���}޾6�྿Pw�~x��w�Z�>���>�l���K���ڙ���F��`�Ž�*�6x�>�>�>�?x��>��>}��>���������'G�%o������<�;��j�u���?(�L�=o���8m�f�>��`���>���>L�>X4�>�I�>�����ep>�:>�_P>�ۢ>�(8>XA\>� �=-_�<��ý�KR?���z�'�������3B?%qd?m0�>�i���������?���?�r�?P>v>�~h�,+�zm?F>�>����p
?�H:=:$��;�<�T��-��n)�������>WL׽�!:��M��lf��j
?�0?+���̾<׽� ����=A�?�??:*��L�i~{��Z��O����<yс��RN���#�SKl�XY������z���b_��n&?D��?ܽ �^�����{z]� �S�dj3>ul�>b��>W3�>�$>�+۾]&��a�D&�7V1�N��>��f?�Ѝ>�`I?+�;?��P?%�K?�ߏ>��>�\�����>|�;��>.6�>�O9?�,?�.?�?"S,?�>b>���g���16ؾ��?�	?��?��?�?����g���@y��zB=�e|�黄��;�=��<�7ܽ�]��Vh=T�U>�X?����8�����P k>ŀ7?8��>���>`��
0��}��<��>��
?XE�>s���fzr��b��R�>e��?���k|=�)>���=(����Ӻ�X�=���n�={9��3�;��0<���=�=xkt���|����:G�;Ax�<_i�>c�?߭�>�K�>�R��� ����='�X>�@S>��>O3پkv�����u�g��y>�o�?4o�?2�f=�H�=�/�=����i�����O���r�<ϊ?<3#?bT?G��?*�=?�s#?|�> -��I��M���󢾽�?�N*?E
�>`���;j�����:���?���>	�d�)(Ƚи&��A��A4���Z'>��(��?}�������G�xӳ��_�Ѳ��NF�?��?}�0���*��P�:虿�e����<?U�>ip�>i6�>e(�I\��>�Q�*>[��>
�Q?��>fN?7I�?C�??x��$+���������1~��ȸ>((�?n~�?���?Y�c?�k�=��(�C�Ž�eҽH��3Β�l�׽�=��7>�a�>���>��?M��>dω��a����a���s=��H>(��>�
�>$��>A��T�O>�G?'%�>Ǿ�H��.Ѥ�l킾��5�yu?tu�?��*?t8=,c�]E�X��^Y�>HQ�?�?�)?\�R��(�=��ּ�����n�eٸ>���>�>~ҍ=�B=�>z�>��>�����}�8��UV���?yF?�5�=�2��7o��������ĺ-=����4�`��Bl�_E$�7��=;ǳ�
L���*|��@��^��l���˾ɉ��=�k�?��=gS>g>3�y=h��������:��9jғ;8q�����=4�%��h�;n��o�E=��=~:/=�*��q�˾(�}?l;I?��+?�C?��y>�=>5�3�w��>\����>?�V>ܬP�9���V�;�㪨�� ���ؾ�t׾��c��ȟ�uG>�bI�b�>A53>ML�=,R�<	�=Js=���=�R�E=�&�=L�=n�=l��=��>�S>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��H>��>ǔT���0�h�]���e�#�I��$?�C6��Ծ���>wx�=�$�����O=��D>9=V�$���]�쑛=�����W=.�=���>rT@>ۮ�=˵��0��=��e=K7�=1�G>���;�H����	��Q=a��=��]>VD%>��>i?�/?�uf?@�>�>B��ƾ����^!w>qF�=��>�'0=�9>�k�>��:?{�9?PWH?�7�>O��=��>I�>�>,�C�]�@�޾�Y�����=j��?$��?A!�>��I�-����$��;�k��?	�%?CX�>���>��ɸ忲�/��g,��b��R�=��,=�獾�|a��
�:���{w �!��=b��>;s�>�(�>��>��>�}�>��>��>�"�<>�b=�ߝ<�5=�.���o�=Q���B~=�J<*$��JS��\�<Yʊ<
q#��փ<�:;,^�=(|�>Ӡ>a��>R��=����.>FҖ��L��N�=执��A��c�K2~���-�7/8��-C>�V>J�{��ԑ��?�=W>`�B>���?Z2u?	�%>���оw]���k�"�[���==�>�59�y�9��:`��N��7оۇ�>!l|>}�>�Q1>��4�3>N����=���#C��~
?tS������?���?���{�w��{f����J�?��~����zn�?��Q?�"�?9�?y�Ǽ���;-�>.�þ��<�����ʖh�uX(?J(?��>W�v��73��3̾B��<
�>�:I�	P�����S�0��9!�u׷����>8�����о3��b��Q�����B�53r����>��O?��?�a�R���JO����l#���I?.bg?	�>a?[V?����11�R����=[�n?!��?2:�?j�
>�>��콡f�>�b?"s�?�̣?�~m?d��=�&�>�W��A�=�ʏ�v�R>�Ꞿ�x�Rk>�R?�J)?��H?^��ԉ��y��Aҧ�k�c>�<�=Eg?��>��9=�1Ӽgؽ�轣d�=�ry>��J>j��=���>P��>�0�� D�p�B?�=>]�>� ?�S�>�����Tő=F(۽S����ɷ������=���H���36=)*���>�k¿�i�?�K>�S��y�?����l�=��>�2�=�FC�j	�>��A>��F=��>�:�>=��=��>F>�FӾO~>���We!�U,C�G�R���Ѿv}z>���>	&���Uu���AI� n��Hg�=j�c.��+<=��ǽ<H�?p�����k���)�"���c�?v[�>P6?>܌����ذ>��>ɍ>�I��B���ȍ�g�;�?a��?�b>~1�>��W?;�?Y�1�e�0�Y���t���@��sd�'�`�����r���
��:���Q_?xex?��@?�X�<��z>��?m�%��2����>Gn/�@�:�)!4=��>⯾9k_�M�ѾF�¾R����C>��n?�%�?C�?JW��m�l'>h�:?��1?�Pt?H�1?�;?_��R�$?n3>�E?�p?�N5?^�.?��
?1
2>|�=k���z�'=47����ѽ�}ʽ���j�3=�P{=�i˸I�
<
�=q�<�c��sټ�l;�Y��'�<�:=��=��=(�>��Y?���>���>�{/?杽u��y���:�&?�����*�#����O��u
��~=a�^?TJ�?��K?��r>WLQ��pG��/8>i$�>+Qt>�>b�>�'6���G��`�=}LZ>?��=W�A=zr?;� �����&��8;>ВB>t�?Oɐ>^�Qi[>�����WC��>^?���ቾE��L���%��p@���N>)L9?�t+?��=N:���>�<�`�S�?&�M?&]?}?��,>�޵�,�L���=�K����̢>r�ƻ�����������<�<�9>_��>]�B����BP>a�	�G��j�g��J���'Ɗ=�W��5w=����zƾ�����=?>�u�����$���@��wUI?Wd�=�$����[�浾d >p{�>���>����}桽Z�<�ܹ����`=�r�>��:>Ƥռ�����gH�����h�>�e>?�cs?��?\Mg��0D��`0�&��7؁��f>��%?��>M�*?�`>��	>f���mS���R�)]�s��>/��>Ď���1��蛾��߾��%��Y�>�?�Č���>N�M?���>�yt?�!I?��	?_ܢ>��:������'?M�{?:eN>H��cL�,y#�k7G��A�>�s2?HEP��͊>�-?��0?��4?��X?9�?�>g>U*�/Zl���>+��>�&K�FѬ�xL�>��J?�?�>��t?d*�?l�=�FY�K����>�S�
>��<>�D?�$ ?��>P��>���>�˾�˙=>��>Q'~?��?J�f?�o����*?�Z�=
��>��پ��>��*?��F?��M?�	C?��,?��.=�ck=߈��Z
���!̼�ym���7�w-�1�b=�����׻@}Q=�QW=���=�4�<�sսFU�mF>=��_=13=i_�>��s>(����0>��ľ�N��L�@>҈���O��ۊ�Ռ:���=���>��?Q��>�Y#�~��=Ʈ�>�I�>���*6(?m�?�?*!;-�b���ھ��K�P�>XB?���=��l�/����u���g=!�m?��^?��W��$��B�b?��]?�g��=���þo�b����>�O?2�
?��G��>��~?h�q?G��>��e�:n����Cb�T�j�FѶ=>r�>CX�O�d�s?�>f�7?�N�>x�b>�%�=su۾�w��q��g?}�?�?���?0+*>h�n�Q4���ؾ噉�ͩF?���>y\оt4%?��<P�Ӿ�ue�<���m̾m�*����P���湾�bF�#���H�?>1�?<k?}�?�yb?�����g�mV�~��In�]������Q0�5n5��z>�x,m���� ��$	�����=�~��}A�mk�?��'?��0���>������M�̾�B>�]��A���ڝ=<B���o>=LxY=�Oh���.�8쭾 ?��>,��>��<?[�[�	(>���1�	8�8`���e3>�i�>��>�>!�:7�-���ҨɾJ���2�ҽ2t�>��~?��o?T{?g���Z2��Yz���6�:Ck��w�����>~gD��7->��L��o���H�mz:���M�/ﶾ�>�������~��>�ٲ>}?�?��>M(��Hh��w�s�6�4��Z�>��>�Ղ?��+?��>aCӽ�8��z�>n�q?���>��>2&���L��a�u���>�>�<�>��?L>�:�s(]��܌�d�����(�!`>i�u?˻r��߾��*�>ژV?+�����>R��>S�=�N�ž+��?s�Z�>�8?(`�=�>��ľΕ��҇��V��'?�
?R�x��|���>$%?���>gϞ>��?�> �ƾ��"?$z`?_�K?��B?î�>��R<��: ̽k���5=�h�>��q>�ޮ=Ki�=X���i��T/��=2�=z�}��媽g�,<6�_��; #]<Z�?>��ؿ�Q���ھ�x�&оa���;���8H�>�l�+=$��Eվb���#ă����^ü��2��=R������9L�`�?;��?�{������͔�t���
�A��>�&���U�7OϾ�/��t��f��gܽ�l�!��B��a�>-f���'?����s�ǿb���_ܾ� ?%& ?�y?�s�"�|�8�&� >�Q�<\��R�뾍���� Ͽ3�����^?���>F��_^��c��>�_�>a�X>��q>\܇�������<S�?�-?���>#As��ɿ�������<��?]�@ kA?��(�6�쾟uV=�[�>��	?Q@>iA1�Y�=4��XK�>�C�?T݊?B�J=;�W��
�%Xe?���;��F��8ػ��=v��=�y=,��Z�J>�1�>���KB���ܽ��3>+�>�E#���\�^�@m�<� ]>1�սP���5Մ?,{\��f���/��T��U>��T?�*�>U:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�ޅ�=t6����{���&V�|��=[��>c�>,������O��I��U��=C��	wſ����i�=�0��J;�7Cֽ�D��*齽������{����4��=Ϡ>��u>#�>.y�=�Lx>sW?��c?���>�M�=�����ȧ�/���f�(>9&�dv�˳��T����A��B��Ր���#��y�dҾ�C����4���d'��u�e���x��cL?̩!>�����?��.�T>ܾje�/۹�13��9�ʾH�j���k���?pe;?�T���}���d���׽��Z?h@�����:��nE>D�D�V��=vz�=E�׽��c(��L���/?�]?��������|'>�^���E=�9+?U5?D<<]�>e%?�-�;v��kV>�1>��>��>�>*q����4�?y�T?>
��қ�f��>�g���Bv��\=I�> 0���ٖY>h�<�O��kk���z��x��<�\U?���>9w+����h��f+)��y>='�v?��?VǞ>T�l?�
@?��y<J����T�p�
�x�=��W?�j?�>#���ʾ�����i2?7(e?d�E>d��۾�-��#���?c�m?�?C]��F{�2���`�
��6?	��?p>�����C35�X�ǾEt�=��?$�"?J1y��B�>�}0?�=h��_}ͿdQE�W��?��@�?&[�=�f����=5D1?��?�ľ���Ĝ��$k�/�=)?yx��ӻ���?�M9�	?��X?�?�H}��,/��!>�j;�_�?�c�?�t�����������V���f]���=� �=<2�����*)H�r�
�H�#�"���4J>V=�>�A@5>��
?�Jo��@�ƿx����^����&'?��>�5���J�m�q�S���9Z�f/�$P��M�>��>��������{��q;�i+��~�>��
�>,�S�q&��������5<��>���>F��>c,��"轾ř?Lc���?οC���Ý�4�X?h�?�n�?�p?ҁ9<0�v�(�{����(.G?��s?QZ?�q%�>]���7�%;k?4A��� b��D6��?F��N>�3?��>V0��}=�9>O�>H�>�\1��SĿ_ٵ����<d�?��?`��3��>�ϝ?d�+?�������娾h5,���o���B?L/>y�¾j#�=<�
��c�	?;1?:G���]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�#�>Q�?"w�=�b�>�[�=����,�d#>M&�=S�>��?.�M?�L�>�K�=�8��/��YF�GR�1#���C��>(�a?W�L?lBb>��8%2�!��zͽ�k1�m��I@���,���߽�+5>��=>�>��D�?Ӿ&�1?��	�<4⿚Т������?T��>ִ??{�,� ��ő��r�?猝> �@��3���І�ӽ��?F�?,�?�DѾ}Z�K>Tf�>�RU>Jx�=&ŽVѾ��>��d?Wvz�|�������.�>�y�?�@�Ϣ?qV6��? ������ׯ����
�]�K�}�>xrK?rc�wn>>ݠ�>�1N>��u��Ա���u���>~��?���?'?�>a?]d�<-2���"=�߈>yQ?z�?�떽� ��C�>X�?�����������g?�2@]@��W?���׿���2���J*ھ���wC�=IC>�f���Z=�|ҽ�"�;t�����K=���>�`�>{��>��)>۱w>�,>�`���#�=菿鞿� 2�����_��S��$�������|�L�־�J��w����ͽ.�=��q�z���*==��>t�N?e�S?�e?��?��=�>�%�	�=L���e��=P�b>��K?�P?M�1?��>�R��:�d���{���wŪ�HF�>s�z>�I�>A��>���>`�ؽ�I>\x>>΢>�l>�{<^H���B�<�<>�Y_>f�>O6�>�<%><>�'��%0����^�y5�������?Ӈ��ʠI�[���.�i�ƾ��=j�&?Ks�=��ԿJ\����L?�kt����u�J�&=Q�(?Z�S?�>>h���*���Y�>+���E�.�=�%��T���{2�Aq>��?8�e>Vt>�}3�Rw8�`�P������z>�O6?'u����8�� v�^H�d7ݾ��L>���>-B�P4�f���~���h�w}=I�:?�-?Cȴ�����i�u��R���Q>�]>[�=E��=eJM>��c��Ƚ�H�2-0=�`�=5]>*C?�8>��p=�>��{�N�@N�>��>>�%>�D>?vH'?p�&�g⠽�����:�4�l>-%�>+ȃ>T1>-J����=l�>��g>����f����NA���l>5���qZ��y?���=����X>y��=x�
��ME��aG=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿг�>���JW���z��b���
��Ε�>��t?�b�܂�Q[���o?Y."?Qi�"����ӿ�Z��?	#�?�O�?�\P��"����-�03�>�|�?�Un?Z��>�	��P����>�|l?rSN?�î��C��j�NN;?���?0��?f��>�ը?F��?В?�����]�9A�������:�K�=�&?�N>����G/��u��bŢ��ݎ� ���>��;�D�>ѓ�=5_\��>���U����"<��>��`>?"[>�$>%-�>���>���>@m�=v�U<[�%� <����K?˭�?ͨ�H�m����<���=F�^�%?kR4?�f�K�Ͼ���>^�\?�ŀ?q[?v��>#���8��C߿�>}��F�<swK>^�>�i�>�r��9�K>C
վ��D�Es�>�З>;4��ھ����,����>�!?L2�>C��=� ?��#?�k>Wi�>ېE�0>��j�E�p�>�8�>�;?��~?��?����\3���N�����[���M>^y?�5?�K�>,K���a����>�sqL�Y������?��g?T\��O?{�?H??�A?��e>O]��ؾ�̬�E��>\�!?��9�@�"{%���b�?��?>P�>ѹ��5׽�*ټ�y��=��oR?gF\?o&?a"��`�L�þ���<��S�H�.�<��(�M>�U>�Ԋ�=��>�/�=r�o�ov7��t<��=�M�>���={�6�����;?wI�=�3ľ.�нp��r��/�>+�>V���y?i�>�� �����������ھ�!f?��?Ԣ?�9潕�g���T?ł?�E?��?��a�$��l�0���g�������>�$�="��������q����b�������^�	?^c�>��>��>�[2>���>됌�:0�?���ؾ�a��~�+�:���;�����Og��P��������ɾ�Vi����>2`����>�?P>W�Z>Q��>KW2�Q�>2 4>���>Rȴ>���>œP>��=���S^Q��KR?�����'�3��ز��p3B?�qd?1�>i�8��������?~��?%s�?�<v>�~h��,+�Sn?�>�>��!q
?�X:=$4�C1�< V������5����˪�>�F׽z :��M��nf�Oj
?�/?m����̾�:׽������>T�?2�/?�:�~�V�u`h��b���T�z���A(�sP��>e(�#�o�������6r���&�j�	>�_"?,H�?�����Ӿ-��V�w�eL���z>E��>��>�Z�>��>{����;gW��U(��ؐ����>	�f?��>o�F?�)D?j@?AI?�F�>��i>eDi���?��ٽ~�7>�u�>Ab?ΜA? �:?߃!?�q?�j�;����ﾀ{���>�'?�?�A!?�?봾���Ѥ�=�e�=ǃB��>-��=>n��s�Ž��K��&���>X?���+�8�������j>́7?���>��>���b1���<��>ٲ
?@�>� � }r��a��Q�>���?����d=[�)>���=����oҺ%S�=�¼1̐=�P���;�D# <�x�=��=�\u�
���&��:�]�;؎�<ö�>�
.?)0>PX^>"�y��K������F�=��#> @?>�>�f⾖e������vp��C>�ޏ?)�?��=�=�E�=4��Jى��z�����>����>�uN?�??"͋?ȉA?��&?i�>z�˾����A�� 6%?T,?�S�>���urʾw�D3�q�?�/?��`�
x��)������ս�>�`/�|~�ﯿ*D��$Q� �����?���?�&E��6�Ku�'�����mwC?���>g�>��>��)�k�g�.�[q:>eW�>�R?
��>O9P?K�?��]?�]D>v+�Ya���7��Г�j)�>[�F?��h?��?Y@f?�S�>2� >�%��C�Ƥ �fǼ�P��=q�|��<�B>$:�>T��>��>���=�0��3⽛�έ�>V��>�q�>sJ�>��>�U>���~�G?���>�]����줾zŃ��=��u?���?��+?�W=I���E��G���I�>Co�?���?4*?d�S�[��=V�ּⶾL�q��%�>.۹>R1�>�Ǔ=A�F=�a>��>���>t(��`�Jq8�lOM�8�?_F?���=����SQr��q?������r�<	���T�ؾ��;=����(.>�{ �����76��R�Y�騕��]�k�Z���޾_��K�>�J�=<�&>�%�=cF6<_Dм�@=�G��4Z� �=�Yh�]2�=U)�� "=e	Ὡ*��c��u�<�8@�A@ʾ\j}?�I?�+? C?�+y>op>�B�3�>��a�}�?��R>5x;��M���X:��I������1�ؾ�6ؾ�tb�㎠��H>��O���>��5>�7�=*Ҁ<���=V�c=�,�=!��:��(=��=��=�a�=�2�=�>�i
>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�7>Q1>ǴR�č1��D\���b�2�Z�}�!?�-;���˾Cۅ>��=�1߾��ƾa�*=�6>[�f=�i�@\�]��="ly�ǥ<=��m=܉>�D>-w�=�ٰ�y��=E�H=hq�=O�O>������4��)���4=�R�=0�a>)�%>���>�?��0?�]d?8Q�>O�m�8�Ͼc����t�>�@�=���>��=�6E>�q�>�8??D?i�K?�j�>V�{=��>�A�>8�,�X�m�s��𺧾$Ҡ<x
�?E�?��>�<�@��U�0-=��I��Q?�U1?j?��>�l��Yӿs�侘>�/�JO<o�<�ӻ����1ހ�|�2����ٽg��>>��>�v�>wb>��=�J�> ��>��>��U=�)}>��/>ȫ���=���ͤ=�5=]ʕ=�$4��V�=��X���ҽ ���޼;E���2q���`=(p&>�D?��-�/ч>�|�<��Ӿ�>�O��r���C>\���͖4��q�ȿ����Q�A!��k�>��>�����i���/?E��=�Zn>^�?���?�8>ng�S���������=0��9?> �>����2�p�G���N��������>8\�>|ݢ>��l>q&,��4?�(x=� �?y5�~�>��] �����>q��F�������h������D?M6�����=�~?-�I?�?m�>�n���Iؾ��0>#`��9�=	.�R�p��<��z�?��&?�B�>��뾽�D��H̾R���޷>�@I�0�O���Z�0�U��(ͷ�2��>������оk$3��g�������B��Lr�M��>$�O?��?N:b��W��MUO����a(���q?�|g?.�>�J?�@?�%��z�r���v�=�n?ɳ�?P=�?Z>-Y�=�VŽd�>�W
?5ߖ?� �?r�t?bB�!(�>b�|<��!>@����~�=�>t��=��>�
?�O
?��?;K����	������%��kV�_�<�j�=ƌ�>�Y�>;<z>q��=��J=U�=6�Z>��>1g�>�`g>ִ�>�o�>�������\�>Kj>R26>Q-?�Ս>b�=]��<LSn��>=#9T��J�2::�ll=���������$=�=',�>��ȿ��?Q�>z()�� $?��˾�5=�e��=��=^B���N?ͤ�=^�$>�/�>cR�>ױ�=�@>��>Y����v>[��>�G� 	J��X�M��th�>AS��׿W��S3��x���G��,�����}u��Ɣ�ݡH�(��(��?���<�"���M�X�ɾ.R?N��>XB?�z��8!���8>��>��	?O�.�R1��+��Xz�a��?�Q�?�;c>��>H�W?�?ϒ1�*3� vZ�+�u�l(A�-e�U�`��፿�����
�u��-�_?�x?1yA?�R�<+:z>Q��?��%�\ӏ��)�>�/�(';��?<=s+�>"*��-�`���Ӿ��þ�7��HF>��o?;%�?vY?8TV�/'�=�c׼�%?�8?���?B{x?�c?����k;?�4>M��>$�>�&<?�7?�D-?��> ��=n�:�s���
��n���+�8���"��� ���2�\�6>�����@=�9M���*���M�����&=�p<��=�4>���*��>W�]?p�><��>��7?����W8�;��vQ/?�4=�ς�~芾����#�G�>��j?\�?��Y?��b>��A�ޯB��>v��>�'>�]>DN�>�f�^E��)�= >�y>�c�=��K������	�eۑ�$��<�� >���>Q.|>�	���'>�z���+z��d>��Q�`ʺ���S�'�G���1���v��Y�>�K?��?Ξ�=�^��.���Hf��/)?�]<?\NM?F�?h
�=~�۾��9�7�J�B�%�>�W�<X������I#��I�:����:��s>*0�������a>\���޾$~n��J�M6�Z�P=�o���U=KC��rվ��~�7�=;:
>u���� �����窿$>J?<�k=���3�U���X>Р�>�I�>�<���w���@��c����=,��>�3;>�ݛ��ﾃ{G�04��m�>��<?Yn?]b�?M�7�x4Q���*���y_��5�=�?�>p>�?Bi�=<�C>��P�iu��l�ɍ+��P�>4^�>��=�'�M�����w/��%�th�>ǒ>Ǖ����?��o?�4�>���?�~?���>V��>��i=Ƀ����.?�e�?hx=��+�24��?;��!�ٜ�>D�?�̤��ɪ>�H?Q�?3K?Xn\?]�?���>����yl)���>�>!Rh�#����Z>j�M?]B�>�"[?��k?Q�c��3N�IF{���=��>�?>�?. 
?0�$?,Ű>&!?�o��=�>�$�>iǂ?�K�?gN?�+����?��q>�?Њ�����>�T?=2#?��j?�.s?�G?��>���=d`���u�O�=���=Kj�=7��<'�=�!�&��K�����<!{>"R�����1�:&V�L翼�(�<i^�>��s>\
����0>��ľ4L����@>�����K���ۊ���:��̷=ۃ�>K�?Ʀ�>�[#����=���>�I�>P��w3(?_�?�?�$;L�b�R�ھX�K��> B?���= �l�������u��h=��m?��^?ٞW��#��N�b?��]?;h��=���þv�b����e�O?<�
?D�G���>��~?f�q?V��>��e�':n�(���Cb���j�Ѷ=Xr�>KX�R�d��?�>s�7?�N�>'�b>E%�=lu۾�w��q��i?��?�?���?+*>��n�X4࿵ؾ�(����P?�?�>��վh�?l =��%�����J��Ǿ_G���#����ƾ��v��ߺ��B����>R?��f?�)s?�e?�Y�>nV�$�L��4����m��Z�_8!��_7��E�j'/���O����H������=��{���?��V�?h3(?�/�5��>{���	��oʾ��G>�Z�����/�=sy���5G=Д]=C�i��4�z4��T?#Ϲ>��>>�;?�+[�r�>�~1�Bi7�Ic����0>�>8�>N��>��%;P�,�t��*~Ǿ����>Ͻ�dj>��i?�q_?:1p?<�)��S,�ކ~���%�n�ͽ,��E��>��R=��>�KP���1�u��WM7��[��o˾J����c�}\=2L�>�̭>2?qV�?K� ?�������A��j/B���=b֟>��n?�?_��>�-{�4�/��0�>��f?~��>h�>���-���{c�mн�>�P�>�?�f[>��Q��^��͒�eZ����:���>�g?�!j�䨓�1��>-mI?9����0'��ɛ>0����Z$���˾�N���%>qt�>��	>�>&Kվ�
�$c�����E.?�?AJ�����>�%?���>���>��?5��=q~Ӿ�����"?M�f?��L?>M@?��>��Q=&⭽��ڙF�ho	="��>��>��>\��=�\�`�⽘M
�_ ����%���r��v��<��+��Y�<��&��V >��ڿT�L��׾����Y��������ة��~�����o��ͅ��T{��0��R7�XD�Yᒾ�ؑ��Z�?�l�?&.��q	��㈘�T��-�9��>jVg�$�㼠���%��`x��>�w���y�#��6���h��m�G�3?MR`��,Ͽ�챿f���>.�?��?&�/�E�D�1�S�W��>���<��\<8�̾���,ѿB��QqC?�=�>j	޾�X8�0�>��>�+1>��?�Ǿ����O=2N'?�"?։�>d�F���ῒ�ٿ"7==\�?.&@1}A?6�(�>�쾌V=E��>��	?�?>�R1�I���� T�><�?
��?��M=t�W���	��e?��<a�F���ݻ��=�7�=eF=���C�J>[U�>��bQA��Bܽ]�4>م>5n"����T�^�k��<م]>��ս�9��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=���{�ƿw����,�~y=�F=��ٽ��M�,��jM�9Yžw`�r�����<�F> L�>9�>��o>���=��Q?&�z?Am�>34/�zH�t���B�˾�x=�И�L��5�`�2a>�<����Y�Op�}��F�(��*�m�D�z�`��M����A�$�b��Ȉ��^M?Oz�=Z|���x�OV�>M&T�����O���7=	�<k:W��9���˚?\*0??w��wH�C���6��q/����?獂�'ܾ���j�i>��;7�<8<�> FF=�f�_�?��1F��{/?v�?�w���Ɛ�&>N�����=�*?A�?C4d<kH�>� $?�7-���$T>�R/>9^�>�[�>�>�֭�k����?A�S?�S�����H��>�����{���p=�	>Ow0�5,���^>[<mю�^�i��ن�P�<=W?z��>L�)�1���_��5��S>=��x?{�?��>�vk?��B?�¥<GA��l�S�N�pGw=��W?/i?��>9߁��Ͼ^q����5?f�e?��N>�h�&��B�.�(h�z?5�n?Q?=����h}�Z�����,\6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?r�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������9�=P����ħ?Є?r���9���.
�<�q�d���,<o��=$XH��f�m��m�=��.ҾV�j���zC�;s��>�F@U/L��+�>I�#�G	��"ɿ���2�Ծ1�m���?`�>��нD���f�]�g��?�@�=�E��oN�>�>X���v�����{��r;�Uz����>���>D�S�'������N6<n�>*��>���>7?��A꽾qę?h\��f@ο몞����ѴX?Af�?�o�?"k?u$8<f�v��z{�C7�3G?h�s?~Z?�P%�/(]���7�G�p?@��A�|�ɈI�0sh�Ȗ�#�?�j	?�}���>i��=�D?�c��Q2���ο��ȿ	���̶�?���?r�ݾ��>��?�*c?��K�St��#�T��Bl��PK���z?���>�'��1X���6�(TľI��>O�-?Z��P� �]�_?'�a�J�p���-�w�ƽ�ۡ>��0��e\��M�� ���Xe����@y����?M^�?h�?ɵ�� #�f6%?�>c����8Ǿ��<���>�(�>*N>]H_���u>����:�i	>���?�~�?Nj?���� ����U>�}?%#�>��?Ά�=Bd�>U�=����|s-��`#>(�=0�>�&�?�M?q@�>U�=m9��/�=\F��ER�����C���>��a?��L?�Ob>����/2�r!��uͽ'd1��S�X@�a�,�ڠ߽�/5>��=>�>�D�K
Ӿ��?�n�ؿ�j���y'��/4?�Ń>�?G��p�t�_W��?_?�x�>�6�9,���'���Q����?�F�?%�?i�׾��˼''>d�>@�>�Խ/��∇�X�7>"�B?D�*E��6�o����>/��?Ѷ@Aծ?@�h��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*e׿�C��q@ƾA;˾4d=s��=cPS=���&>�#>=�<{��y>��>�$n>K��>K�z>T�t>	Ge>7��}�%�7���}���r��/"��#�Ef�t�ۄW��:%����3ξ	�'=�������b����jbG=���=d�U?p�X?rin?ZF?��輝�->����P=�*(�
�=[>�p)?�G?Է(?IY�=�����a�m�{�ܠ��S��\<�>��J>G��>��>I�>I�;K8`>��T>�Z>��=f^�= ��}�=+Xm>,��>?m�>L�>Y�?>���=�۰������6[��Ȼ�K"��� �?�ξ��U���ɬ �ҧ�1��!�<?�>�u��:�ٿЕ��*�W?�;>��"������<�2?1�z?�K>G��~�#���>Xw�K����>�������p����>U�E?��f>�u>Û3��d8�	�P�d{��{i|>A26?�綾uD9�Կu�m�H��dݾ�@M>N¾>�,D�l����8�ui� �{=�w:?Ȅ?^8��
ⰾe�u��B���PR>/:\>�i=�l�=EVM>^[c�p�ƽOH�[q.=���=Q�^>,8 ?6+>��q=`�>����OI�3߫>�5>�	3>�=@?��)?V���#׽Av����W� �I>'_�>�U�>uS>�:��o#=��>� p>��q��I��av	���C��#>��O��π��bL���<	�R��$�=�i=F����:��r=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�g�>cu�iZ��6��g�u���#=
��> 8H?NU����O�� >��v
?�?"`�賓�b�ȿ|v�E��>��?��?P�m�X@���@��~�>��?XgY?Vpi>5h۾�ZZ���>�@?lR?��>�:���'���?�޶?c��?|{i>��?��?y?@|�b\��ۣ�����.���N>���><�)>�����U���CJ}���{���
� ��>��h<���>���;��k����>�E	���վ���<?�>lv>!�>-C�>��?_X�>�B�>7��=��=�r�`�R�.�K?���?X��?&n��-�<��=N�^�T ?�L4?a�`���Ͼaè>G�\?�Ā?B[?l�>����8���῿�~�����<��K>(;�>=M�>O߈��0K>��Ծ�D�k{�>HǗ>襼&@ھ�!���L��LB�>\d!?`��>>��=|� ?�#?T\j>b�>aE��,��a�E��y�>x��>�??B�~?��?�����\3�3��:ߡ�`�[�x8N>��x?H?V��>hm��Pn����J�(tJ��������?�Qg?'I�?�/�?�m??6�A?��e>���1�׾�ʬ�+�>��!?��T�A�>&�@���|?�K?c��>)���6tֽ��Լ����l��+�?z\?�3&?}��ea���¾L��<��$���S��<��D�$�>|z>������=�.>�N�=�Fm�BP6�6i<��=�n�>4�=� 7�wU��2=,?c�G��ۃ�s�=��r�ExD� �>�IL>O��ì^?el=���{�����x���	U�� �?��?`k�?���@�h��$=?�?V	?k"�>�J��~޾T��@Pw�~x��w���>���>D�l�{�7���ܙ���F����Ž>K�t
?Q�>#��>�b�>�OD>��>�T���_����l����R\������L�zZ.��g�-U���F�K�o=�s���zv���>Q�&G�>V2	?�V>��w>;��>�����>3
C>�F4>'�>�M >�)O>5�8>`�X=�W���LR?������'����)����4B?0md?q)�>h�<���n���x?ψ�?�s�?kSv>Lqh�� +�`k?W5�>C���f
?FD:=g<�7�<C:��������p[����>�l׽,*:�>M��Wf�Sh
?C,?L���b�̾k>׽P����=c��?��+?͟0���M�U�Z���`��W���D�SJ����6��nf���u���oʆ�x�"����=�)!?�ʑ?5���}��,��{z�e�A��s>_��>b�>���>0�g>K��&��$�U�����{�z�>N'p?T��>K_6?cM?��R?;`Y?Լ�>�ެ>^]���A"?����'�=@w">�Sg?̡O?�xH?�]%?�7?�2>ˋ���:��K�?�(?ȩ+?�?G��>Y>���n�=w&r>+��=Ó�T��<D�=O�B=����UY��HY�l˘=�?}S���9�����>Y>,J4?�J�>��>Ρ��]�z�N,=�U�>��?�>|>�5�%�p���/��>�U�?(����X�<h�2>��=�.�ֽ��=��=��ڻ�,�=� 4;�Vʼ�|�<O�=IY�=:
�y��k�%;�(�<�/�<���>�&?+g�>�!�>�q��ޤ���J��Ъ=��[>�bS>�p$>��ؾ�B���0��#�h���s>�?���?��|=0��=���=�眾[�����Ͻ��N�<PZ?g�!?�T?T�?2>?�?"?<u	>��`���Є�p���;�?�?,?XB�>�W�@]˾2ਿ3�3�f�?�?q�a�����4)��G����Խ�>X�/�܊~�����aUC���%�i���%�����?)؝?	�F���6���}Ԙ��Ҭ���C?���>df�>��>�)�Hh��	=>���>[R?��>\�P?�%|?�_\?�T>�
:����Cs��� ��oC'>�A?3�?F�?��w?�M�>�>��.�x�྄3����&�2���9����/E=WT_>��>��>ψ�>���=��ֽ�����TD�qҶ=u_Z>�j�>��>ٍ�>f�v>�/�<F�G?���>8[��A��#夾X���s�<�K�u?���?p�+?�c=��j�E��<���M�>�n�?���?�4*?�S���=��ּ:綾��q��'�>��>�1�>�̓=��F=aU>��>��>�
�qc�q8�LM�(�?�F?2��=H�ſ�3q��%q�F"����M<.C��Fh�.	����Y��ˢ==,��n����O_�ɠ�R���kH���J�����w�>���=���=���=o}�<���o�<�W=	)�<Z�=��y���<}�)�#j��6������ ϟ<h@=��B�{ݿ��0|?��O?��*?~�C?7�>�s.>�C���z�>�W���@?��>zɕ�S�����#��v��������ھ�Aо (Y�Kp����>����>��V>1�#>��=B� >L��=�#=�ؚ�s= v�=`>�`>W.>�]�=���=�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��2>��>�ES�߬/��`���]�<�T�B�?%�6��rʾ6ԍ>��=�]��̾D�=�".>�=@={|�<W����=�3��N�D=�v=�҃>��@>)��=����Kl�=P[i=��>>bX>��|K��#]���=���=~l>�?'>=��>�?K>0?�d?��>�Hp���ξ����ҋ>N��=�y�>��=�B>`V�>}<8?ΔD?��K? B�>�M�=��>�1�>k�-��m����%���UH�<��?��?�]�>��?<l�<��3���;��`���!?Us1?^I	?�N�>U�����X��*2���R��<�=��.n���AX=�S��liq�es���f�=?��>+��>Q3�>v�>�_�>��>�a�>�gh>��=l0k=P�>�u�<"F= �=����c/���޽Z�T=TA���8����<F�=�D�<��=:苽���=�z�>�>��>kړ=����/>����L����=�Φ�BB���c�7�~��/�n�7�WN?>�%V>[��������?{qW>�5@>���?�Gu?��>>]�OZҾ�Y��!�_�|9V�>��=4�>^:�h :��L_��N�w�Ѿ���>bf�>�%>�\�=)�T��=���i>�ξ�	C�J?��[+=hЕ��낿�a���(��� x����=H�E?�Έ��؋>�N?��=?�]�?L�?NG������?��ǚ=��c��ȃ������v:?+PU?���>��4�B,��F̾����շ>G?I���O�;��� �0��]ŷ�P��>5骾=�о�$3�h��7�����B�_Tr��>��O?<�?�Ab�T���QO����2/���p?�|g?F�>sL?q@?���Dx�i���R�=B�n?L��?P<�?�>KZ�=D)��Y�>pB
?}y�?���?]�q?NyD� �>iVP<�\">3_��[R�=��
>H{�=���= ?�s?��?��<	����<���`��<|$�=eŏ>���>�`t>�j�=MHm=��=�H>J��>�ԏ>��^>~F�>�{�>PD���5���?���=��5>�r$?b�>��D=��Z�r2�=��=�2�V�f��� �v�N�K�p�c��\"�=���<#��>{lƿ�`�?�|>�
���?�澬����:�=IP>�aZ�#�>j�=s��>r:�>K�>c��=d�c>�2
>�$Ӿ�>^���F!�>'C�VLR��XѾ��y>�&��d�%���H�����I�U۵�����i��%����<�U8�<�*�?!���fRk���)�����a?�Y�>�)6?�䌾3
��@�>�$�>G��>�������a͍��T�A�?r��?�;c>��>3�W?'�? �1�63��uZ�P�u��(A��e���`�_፿"����
�X
����_?:�x?�xA?GY�<):z>z��?R�%��ҏ��)�>/�';�D=<=�*�>*��a�`���Ӿ^�þC6��GF>A�o?%�?AY?�SV�ҤT=��9>`S?b N?�r�?��l?�*?F�}��M?w��>%��>�>��P?�?]|?�>�u�>��;�-�KÏ�ʣ��g�w���M�D2����U+m�������=�N:>���<ą<�Ů=��=��Y>���=�^�=>�'<��=�ͦ>�]?�B�>���>l�7?�j�EQ8�9����//?�>8=8����-���m�����KR>0�j?^�?�?Z?�Dd>��A�'C��>uU�>B\&>i3\>�=�>v��B?E�B9�=�$>C>~o�=�M����ٳ	�q�����<$>���>t/|>�
����'>�|��R.z�٥d>��Q�̺���S�9�G���1���v�Y�>h�K?��?晙=-_�*���Hf�H0)?�]<?OM?F�?��=K�۾��9���J�>�;�>4O�<N��i���e#����:�� �:��s>�1��!����,a>���s߾�n�lJ�I�辒�R=B�e,R=�I���վ'7����=TF
>�T���� ��-���֪�WGJ?wl=������T�&Ǻ���>�z�>V��>��<�|{���@�S���O�=���>�;>1������m�G��+�D{>��F?�^]?.�?y^���m�p�E��I�9���yc��n�?%M�>�c?�w>5q�=/���.����X��D�P��>u��>oI�JH�R���޾
d��Ė>D�?��>	D�>i�M?J�(?�u\?8�,?_�?���>7g��z:��!&?���?Ɨ�=�ӽy T�l�8�:
F��8�>�k)?�7B����>֢?��?��&?A�Q?�?R7>�w �u�?�ho�>咋>cW�%=��C`>ۍJ?�ó>�JY?�σ?�>>^5����㐫�i�=e
>�	3?��"?(�?��>]4?3�� �`��>W,@?Y�o?A9p?�$���B�>��>GV?o�=b"W>b��=rB�>3�h?A{?t`b?�	(?s{�<�����@5�O�>��lּ�v׽E�n=�A��Z^�������=�#?�>K�緡=�S��������<�D���^�>�s>�㕾�1>��ľ3��>�@>����`�������Z:�D�=���>��??��>a+#�B�=2��>�Q�>o���6(?4�????";Жb�)�ھ�K����>��A?���=	�l�����u���h=<�m?q�^?7FW����G�b? �]?0h��=� �þ��b����Y�O?7�
?G�G���>��~?a�q?X��>��e�,:n�)���Cb��j�Ѷ=Zr�>>X�U�d��?�>v�7?�N�>J�b>�%�=Uu۾�w��q��y?��?�?���?�**>}�n�P4���苿��K?��>'��?�d�<�Ѿ�"U�A`��0�§ܾ�O�\��f~�� �a�蟾�vL�B5�=�8?)U?�p?O `?R1��v���m�4�}��%_��<�{q�۾9�iKJ�U!�B�m�������:���g=<�}�_�>�x�?>�&?�:����>_����+ľ��B>�^��2��
h�=E@1��G/=��4=Y%k�;�;������%?�U�>���>QG;?N9_��A�VV4��7��>����0>��>$�>SF�>*g<��,�����"���SS��*IֽLV>��k?��I?�q?wT����=�'�~��r&�/�o��3�����>NG3>X|�>>q�����,�~1>��b�`<�S����J����)>��	?��>C�>�G�?@�
?kq��?{ ��#�i|*�Q�Z>�`�>��a?��?G��>�3ڽmt�"��>��l?���>�k�>ء��ي!� �{�k ̽�A�>�N�>,��>�o>f�-���[�.���D����	9���=�Ah?�r��v�`����>	>R?�B;~C<�֡>i�x���!�y��.%�>�>Y?�8�='�;>azž��6F{��ъ��T)?�1?�Ò�lv*��q~>e "?Qv�>��>)/�?S�>/)þ������?��^?CEJ?~RA?�e�>�=�����2Ƚ�&��8-=�y�>4�Z>�m= 3�=�x�2*\�x�1 E=�D�=��ϼ�=��&d<+���+M<3��<��3>}翀4Y���� 4!�~i��4���ю�cX��6�c��P1��=پ˹ξ���I,	���}�F�D]T�j������d��?<��?S:e�6A�������_y������>�� 
=�ܧ��Z��^���ﾡ汾W�A�E��X��K���+?��gϿ� ���g��?��>F7?�}�?�����H���E�p��>�����>����\�����ʿ�|��,?%�>P��� ��=�c�>`�W>Q=�Ӛ>�����o��N�2�?�D?ࡰ>v���¿����$����?�@wA?��(�0v�~W=B��>�	?&bA>�1�Nz�%(���~�>Y��?3��?��G=��W�1����e?�<$IF�+�ջ���=0X�=��=K���0J>qڒ>�g�o�A��?ܽ0:4>C7�>z^&��s��^�wo�<�%]>�9ҽxJ��5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=l6ἧ���{���&V�|��=Z��>d�>��,������O��I��T��=���t�ɿ�%���-�/��{�4����Yӽ������Խ/`�����I����W=�3�=�G>k�}>*�>��>�SY?ux�?��>�1V=Z�E՗��׾b��<�*������D���=���F��A���߾l��X�������*ly����tlP����2d��}d�Jω�, K?�K�=�<��?c��=1���٨�m#�=��<~#��^�s��j��d��?uZ9?�o�:�%� ��9�9�z�A�H_�?��6��/(��+�(V�=0�l=��=}��>0�f=&!:���n�΃;��w0?cU?����fU���?*>E� ���=��+?׌?�aZ<�3�>P%?q�*��+�Fo[>t�3>��>���>�I	>���A۽�?��T?��������ː>e����z�FIa=�5>�/5���輚�[>�>�<�􌾈MV�f[��\P�<.(W?Y��>��)�Q��[��в�q�==�x?Ӎ?�1�>�xk?��B?�9�<�s���S��E�w=E�W?W+i?��>󐁽$о���� �5?�e?G�N>�Zh����f�.��T�l$?��n?�]?Hĝ�"v}����^��8q6?�av?J�^�l��%/��cM���>���>�(�>p�;�j�>�??pd*�i���	o��&�2��ڞ?�#@ ��?�Π<�	�;ґ=MC?�L�>CYO�����ћ�������q=���>����ǵv�8# �R1���7?-�?�M�>!���q�#�=;t���?<�~?��辏������@�g�9���:����<��?�b|i� ����I����:)��Fƾq]�aK�>��@�Y�����>4��߿�W˿�q�C�
�د���s#?�b�>bg��<�Ǿ��n��M��Eh)��#&�P~�� �>��>��������{�o;��~�����>����>1T������a���t/<S-�>o �>r?�>�ﰽ�z�����?�:���/ο���}H�+�X?�u�?h�?��?�#<hw�X�|�l�fG?��s?{6Z?�["�N^]���8�"�j?�2���;`�Ȃ4��fE��T>�3?R)�>��-�p~=.�>(��>b>�B/�ܕĿeڶ������?��?:��C��>T��?��+?�^��1���}����*���G�LA? 2>������!��G=������
?�r0?���v(�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�#�>��?�s�=�b�>�c�=��C3-��g#>��=��>��?@�M?�K�>>Z�=��8��/�zZF�]GR�f$�x�C���>��a?��L?�Mb>����*2�W!��wͽ`b1�5&�T@���,�.�߽I*5>;�=>v>��D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	? �{P��q`~�c����6����=D�7?2���z>���>o�=Knv�ƻ����s����>�B�?i{�?���>��l?�o���B���1=M�>��k?rs?�o���-�B>!�?�������cL��f?��
@8u@Y�^?Um׿�Ƥ��M���u���M!>���=��\=Խښ�=L�<Aّ�'����>ᮂ>2�G>&ch>\>�Vw>��>�n���.�:>��D�����=��������L��:�\ˎ��/�`�۾�,�&�ҽ�^Ži���]�ܽ�"�Kt.�f�=�VY?i�^?>k?��?�L�	�>�q���N=�.�h:>;��>=UL?�T?t\(?�G�=�흾"Y�F�w��7�����\�>tտ=�I�>�<?ޗ�>-=>;>y��>�9r>j�\<�W9=��8�p�X=��>+��>�S�>���>�>+zR>�e¿f���f	�����Nt����?է���w��
����<���H�1�<��R?�A<s/����Ͽ����
f?0��y4���ü�=�G-?�y?��|>�S����(�|�!>����Od��i�>�[��V��/P(���?k?k�`>u>:�2���6���P�W���ņ�>��4?#ʲ�~�:���t���I��n߾��O>8�>�z�����}����}�6�d��gL=�v:?͔?C,ǽM˱�Xiz�<���r�L>�|b>��=S��=}$A>�K�P)ƽ�*J��f.=��=��W>4�?�$>�k�=&!�>�d��zG��>u<>�[ >��@?�h%?.�&��s���,����,�R�~>���>��>��>�|H���=���>�a>�}	�:z��0�n�?�r�U>��v�b�Z�����g=~`��K}�=�أ=���]t8���=�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾMh�>rx��Z�������u�j�#=S��>�8H?�V����O�i>��v
?�?�^�੤���ȿ5|v����>W�?���?g�m��A���@����>;��?�gY?voi>�g۾D`Z����>ϻ@?�R?�>�9�w�'���?�޶?կ�?�7>3%�?�ZL?�Q!?^;=0T�BT��[Ց�����@}��)�?��=X�*���%��䍿������A�GQ�P���x3<�ʟ>J`�ZW��G>>�I���Z���C��$$�>�V4>��6>z�>΋�>�u�>H	
?B��=&��=�����Y�K?���?���Q5n���<���=7�^�k*?_G4?�\�l�Ͼ2ب>m�\?q?�[?_�>U��|=���翿{���Җ<��K>�1�>EH�>�.��ALK>��ԾG1D�m�>�ӗ>����:Bھ(���£�<�>bd!?���>}�=�� ?Ȝ#?��j>)�>,aE��9��h�E�!��>��>�H?��~?��?չ�dZ3�����桿��[��:N>Z�x?�U?�ʕ>:�������XE�|CI�����A��?^tg?�S�V?52�?�??#�A?_)f>և��ؾ"���i�>��!?w��5�A��E&��pz?.Y?���>�䒽d7ֽ�.׼h��wv����?�\?81&?^���$a�b�¾Kr�<�(��P�[�<B�F���>�z>؞���w�=~?>���=%m�	�6���g<y��=�~�>]�=�$7��쎽1=,?��G��ۃ���=|�r�3xD���>�IL>����^?_l=��{�����x��	U��?���?[k�?��8�h��$=?�?L	?T"�>K���}޾&�྇Pw�~x��w�I�>���>f�l���H���ܙ���F��g�Ž�3q�� ?D�>Ɍ�>c_�>#�>x��>�$���������}0������m�2�D�� ��վp�Z3�=Pw��/E��W>Z���f�>�4?k�>껉>\�>����}Z>]�=f��=��>���>���>y�.>ڍ=��L��KR?�����'�w�辡���]3B?�qd??1�>�i�-��������?���?Js�?#=v>�~h��,+�rn?�>�>(��Rq
?�T:=*5��:�<V��}��D3��'�'��>�D׽� :��M�onf�pj
?�/?���i�̾;׽ϑ��θ�=��?�7)?',��zT�&�m�ڢW���T���b�Z�f�䄬��v*�E�h����V兿Rw��,�)���
=�'?�?�8���s׾W���!l��FB�=U>��>�;�>��>�tW>����4��]���*�C�f�e��>`Ll?���>.fY?00b?S�D?p4N?��>�Ո>c㧾��?�8�=`��>��>��.?�?.(@?�G?�:!?\Wy>�v�*$�"��<�
?B1?-�'?�(?K�?;�C8 =A+�={�8�#ߟ�.d2�i��=wޯ;��3�2�Y�SN�<+��=�X?i����8�t��� k>��7?���>���>���'���&�<�>Ѵ
?-:�>b���qpr�rY�o]�>���?��{i=|�)>���=E>��ʡԺ�;�=+����="y��}m;�!�<�b�=��=I�q�Tɔ����:���;^l�<u�>&�?���>�C�>�@��� �M���e�=Y>lS>�>Fپ�}���$��m�g�^y>�w�?�z�?�f=��=ߖ�=}���U�����?������<�?CJ#?XT?T��?w�=?\j#?ĵ>+�cM���^�������?�-?Yt�>�����
��i���
U�c\�>��8?�GX��5���8����=���U >��(�9���P���q۾s*>��D�ԽŢ�?Z��?7����s5�K���ƿ*����?���>��w>8�>fhx�x���� ����
�>r�{?V_�>vV?Z@�?4U?[>�>+��v��펖���<�� >��6?�O�?A�?�v?n)�>aN"> ���Ծ4\�#�ȼ�C�a�P��7<w�Q>�>K��>���>	>�_��6���v�a��)=��>��>(@�>��>�T�>�^H=��G?E��>�6���I��t��3t��J�2�5u?b,�?D�+?ٞ=ғ��\E��L�����>焨?���?�(*?�gR�K0�=jۼ�|��s���>v��>��>�=�dK=n�>��>���>�-��[�[�8���N���?�F?�F�=]ο�q�LꃾV�̾1F��:��vU���J���7�=z��Ƣ#��������ړ��݄�����J?��v{��?��=���=_�6=�==J��f�� ��=<�9��m=)$H����=)�=G���dׇ��0=bCX=^��;��.�~�˾�}?N�H?�+?�KC?��y>{�>J5��
�>�Ղ���?�(Q>z�J�00��B�;�k����ʕ���ؾo־�(c��5��R[>xWG��~>�k6>�	�=��<C��=u�w=�d�=�W$��I=��=���=���=~��=1�>�q>�6w?P�������<3Q�R罡�:?6:�>5x�=7ƾ@?E�>>�2��ܖ��1b��,?��?�T�?p�?�mi� d�>h���ݎ�n�=yÜ��82>���=��2�D��>v�J>J���J�������4�?k�@�??j⋿-�Ͽ_/>��7>�=>D�R�8�1�¤\��b�8]Z�<�!?]?;��R̾3*�>঺=^)߾��ƾa7.=Ox6>hb=&u�wM\�e�=�i{�<�;=�0l=�ω>��C>"o�=�.����=d�I=���=�O>G��y�7�N�+�N�3=���=��b>O�%>S��>�A?^�??o�Z?��>G�J�F8Ӿ�NѾ�@�>�)�=V�>�>+c�>U�>��??�>?�G?���>j��=;9�>o`�>gL� e��Ծ�ۧ�"��<��?�h�?K=�>`��;reo���#� �A��^���3?�[)?t�?�d�>�V�͚࿐V&�>�.��㙽��J��$)=�Ir�8�T��������㽥��=/:�>i��>�ݟ>eZy>1�9>�9N>�(�>��>��<��=���'�<:����=U���]�</+żu�!��A��.-�u������;+u�;qQ\<�&�;\��=��>e8>��>�=�(��/>�ǖ��L��1�=b:��3B��2d�q;~��/��6��pB>y�W>䓄�B+����?C�Y>g�?>ǉ�?N5u?��>|�V�վ�M��]�d��CS��ø=/�>��<��m;��/`���M�ƞҾ�
�>�M�>w�>��e>��^�ap�|
�`����U�D�?ࡾ[g:�*ҽ]��51ÿ�f��^݅��,�ki@?uA��Z.(>��-?�f5?�۝?��>��=*@���>�_����@>*9`�Q��Ш@<���>K�?*S.?В#��G�LH̾����޷>�=I���O�����0�����η�4��>������о�$3�Og��+�����B��Mr���>˴O?�?�8b�iW���SO����)��\p?�{g?:�>zJ?LB?x��y�1s��Aw�=�n?���?�<�?��
>\�=?L�c5�>�J?7��?�?��u?��T���>@}�=�Q>M���[#>.8�=�=��:>;�?�R?�?�E��X

�S���Q�
�e�R�;�=�t�>˺c>^�/>��f=4�=3u�=��=>��t>��g>xg>m�>��>�ܰ�[��M?O�=R#F>�'?�)�>�v9=x�A���ͼ�5��Ẑ��c���_��1�����·��T�ռ}������>FPɿJc�?���>Da�
H?Z�������!>�>�l�����>��Y=�u�>���>A�>��>!iS>�M�=�;Ӿ�>:���l!�~.C�M�R�˻ѾD�z>~����$&����>W���?I�Xa���^��j��.��9;=����<�F�?����k���)������?�a�>�6?8׌�^ ���>��>*��>(9��z����ɍ�.c��?���?C;c>��>��W?U�?ڔ1��3��uZ��u��(A� e�N�`��፿0���e�
������_?��x?�wA?�H�<M9z>6��?N�%��Ϗ�:-�>�/��';�b7<=(�>_*����`�A�Ӿ!�þ$<�%FF>Ӕo?S%�?�Y?�YV��)��:�=4+v?5�/?$�?7�S?��?�o�:a3?���>R�?:v�>�67?�P7?�w�>:��>�A[>[���V=�a��z²��20�r%W�ξt�z��=w�=EJI�x���5��-^Y�ˢr=M��;��6�|�(�dK��j>+�<�܆>;��>Į]?{�>8��>��7?���%h8��î��./?5,:=m���&�����H��G>��j?���?x]Z?דd>�A�@C�">^�>?�&>/u\>�w�>i���9E��ʇ=n>�>��=�FM�:ā�ɰ	�������<�>���>��|>�F���%(>'񣾸{���c>��R�P��dT���G��2�L�w��v�>�PK?Jg?e��=�龨7��$f��Z)?b5<?KiM?��?�[�=�Oܾ�9��K���eˠ>x�<���������� �:���;�Mt>�����ᠾ�Kb>\��9�޾�n�2J����"O=|n��vT=����վ��~�"�=j
>���?� ���� ܪ�:@J?̥j=���U������>��>��>#�;�#w���@�Ŝ���Ֆ=H��>�z;>�#��h)��G�P��>�>"XE? W_?�k�?���`s���B�"���`��X�Ǽ&�?���>�Z?�@B>=s�=H���R ���d��G����>�n�>�����G��&��v ���$��~�>8?��>i�?��R?��
?ߟ`?�*?ZQ?�7�>H�����v@&?m��?��=8�ԽǻT�i�8��F���>;�)?D�B�M��>�?*�?9�&?��Q?0�?�>� �A@�V��>�Y�>C�W��`���_>:�J?d��>�<Y?	҃?��=>Ȇ5�?颾�֩�8f�=K>:�2?z7#?��?ͫ�>�I�>|α�xY�>�?�>��}?O�?h)o?0=u����>s؈>���>i�L�>#0 ?�'?�_?[�?^�a?%�>v�%;i��Z�����88f=D/�=�_
=������ѽ��0�	r��!ży�0�u礽$�A=���=>�Z�=+_�>�s>�	��J�0>�ľ�P����@>Ҙ��)Q��xي�ʊ:���=���>��?���>g[#����=��>�H�>���^6(?0�?.?��!;��b�A�ھ�K���>	B?��=��l������u�U�g=��m?�^?�W�&��F�b?�]?
h��=���þ۶b���W�O?:�
?�G��>��~?P�q?M��>;�e�0:n�#���Cb���j��ж='r�>QX�B�d��?�>i�7?�N�>+�b>J$�=iu۾��w��q��w?��?�?���?:+*>{�n�R4�������4P?6��>vη�ˋ?�`s�
�۾��r��Gt�ݾ�P��)Y����������*c��!���V�9�=�?qek?���?w�V?���=�`��?d�����~W�v׾���w�'�b�[��z2�CDe�q�!�g���_���ᒇ=�Z}�R�A�5ȳ?�)(?_�5����>託��h�x�ȾKD>��7��z�=b���i7=�8=�l�O�/�=����D?��>n��>��;?f�[��=�К2�.9��Q��]�:>+�>�
�>�&�>.��;l+�`���]ʾ���!�̽�w>�Nh?�K?0uv?6%�R�J��䊿�K��������Ϸ�>a��>��g>lst��z�'e+�i�&���X��G������ߘ}���	?�U>���>��?��>v�*�H"���Y���09�b�=�D�>�u]?c@?r�>�%彄�/��0�>@Ps?4I�>���>.���j(�	���d�Խ���> /�>�T?�}�>�#B��5W�'������*�7�I%�=E�h?}5��1�t�G�w>Y�N?7�(=��,;o��>�F#���$��)��F����!>��?�.>�.E>��������u�������(?Z�	?T፾�R(�6�>R�$?G#�>�>��?���>����BF]�E?D�_?�,K?($C?[O�>$	C=R��B�ý!+)�L-=uK�>�
a>uz=�^�=+����T��)!�6&=:Ա=kS
�9�ν�3�9��<�!'=��8>�߿��S�q�Ӿ���-������ ��#�i�|OQ��Z��.ܾ{q��_�'���ô�[�=��f'�c u�^��A�?VM�?�A��6ľ�S���Ԃ�my
����>��*���6񶾉���zb?� ����#�����'F�*�z������'?�[����ǿK���2vݾ�b?
b ?z?����"���8��^ >���<�[��\��Ja�� �ο� ���#^?�8�>�g����f=�>���>�V>��m>�҉�Y���o!�<LF?�c-?�'�>�r��ɿq���Zؕ<>��?~�@�|A?S�(�j�쾽V=���>H�	?8�?>�T1�J�z����V�>C<�?���?R�M=3�W��	��e?#�<��F�8�ݻ��=�:�=o;=2��ҘJ>XV�>7���TA�f;ܽ1�4>�ׅ>��"�5��*�^�a��<Ň]>��ս�>��5Մ?,{\��f���/��T��U>��T?�*�>Z:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?7ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=l6Ἕ���z���&V�x��=X��>]�>Ƃ,�ߋ���O��I��Y��=�a��dͿ���#)�U=�S�=~%��U�����b��m�]�ƾ>X��K髽-��=B�/>��>�I�>pH�>Y�u>Y?��q?_׳>H�û��A�D֎��پ�,>�܎��\������˽H�Ͻ���X�������� ����M�Y�x�<_^T�B���$�2�B�єG�d�9?��>mC��+[��]�;@߽�*о��컔C�<~s��<1�����jӣ?��M?m&��R�N������M�� �X�h?��	�df����7�,�>� ּ��彧l�>��^>[+����z��;� o0?�S?���"J���*>�� ��=L�+?��?xZ< �>>B%?��*�U<佂T[>y�3>?ϣ>ڱ�>�G	>��Kh۽��?T?�������"ΐ>�h��J�z��Ka=B">|�4��q��[>PJ�<+����W��+��ͫ�<v(W?ӛ�>,�)���a��L���^==��x?��?^-�>6{k?l�B?�Ӥ<�f����S�y��gw=5�W?�)i?Q�>Έ��Z	о����D�5?ݣe?Y�N>�bh�����.�dU��$?��n?"_?�w��w}�������n6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������:��=��!�?W�?α���;�N�=o�����f�*=���=)O��i������	l7�ؾ��xW����t�a؆>��@�~�I\�>Մ9�cN߿��ο���ǄξŦL�S?寨>Q������Cl�B�s�̅G��C�#�pI�>7�>�ϔ������{��p;�E\���>\��� �>w�S�!�� ���55<�>ͱ�>Ӹ�>+F��T��ř?�`��w@οq���Y��b�X?Th�?jo�?m?�X9<��v�f�{����?-G?��s?NZ?�%�AN]���7���j?�]��U`�1�4��HE��U>4 3?�@�>�-���|={>E��>|`>�$/�z�Ŀٶ�����z��?��?�q�i��>0��?�v+?pe�~6���Z��.�*��(��;A?Z2>u���>�!��2=��Ӓ�2�
?~0?)r��,�]�_?+�a�O�p���-���ƽ�ۡ>��0��e\�)N�����Xe����@y����?N^�?i�?׵�� #�f6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�i	>���?�~�?Pj?���� ����U>
�}?�$�>�?�i�=a�>�X�=����׋-� f#>f��=�>���?%�M?�F�>�T�=*�8� /�6[F��FR��"��C���>J�a?قL??Qb>v����2��!�4tͽ[]1��@鼓e@�x�,�b�߽%5>��=>d>T�D��
Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*��Ͽ%x���h���췾��=���=��G>i��e=#��=���<������W>�!�>�_>\��>.qq>4�X>\|>>2.����#���������F���D���`��A��ZN���
�K*���?Ǿ�꡽������ɼ'��� ��'�L��=2lU?T�Q?>*p?+) ?�=��~>���y��<��#�)Ę=$�>��1?�gM?�[)?N�=�*���d�����y�����פ�> C>��>�C�>2ܯ>
��\�F>� A>�~>��=A�=��4�g=�cN>�1�>�#�>���>:�>ѳ�=P¿�Y��"��RΑ�"��;@4�?�����́�걙�����Q�4]</�_?N@�>=��3׿Iʪ�+�X?��v�\��(���a���>�Yv?ۃJ>1�=��� �V��׾��>l݈��V���eb���=i�/?=�g>�t>K�3�%�8��Q�յ��f$}>��6?�z��,s:��u��}H��Rݾ��M>+�>?G����	����~�03i���{=�:?XD?�?��L��q�v������P>DI^>/8=B)�=j�K>��b�9�˽�5J�@�)=Ҙ�=�R_>��?�o)>R��=;�>�����N�m�>K�@>H�/>{G??5o$?���,�������-���t>���>3F�>~�>|H���=�>��`>����?�����B��FU>�<t��_��{W���\=�挽:��=�ȃ=�� ��:���(=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?�A�>��?"0x?F�?=rV��E��u��y���qA�>�in>���>�W>�1�"DM�o��;�����m�f��Dp�>���;^U�>�ֻ�����Xr>T|��Z���9>(�>�5=���>r��>fh?���>�L�>��4<�ON=����T|���K?���?-���2n��N�<Y��=)�^��&?�I4?$k[�}�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��H��<��K>*4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��dS��GB�>�e!?���>�Ү=�� ?��#?"�k>#��>{.E�F���AF��?�>���>>?3�~?E3?�H��ZE3����g�����[��	N>5�x?�?6S�>#m��CN���S+�]�K�;��I��? g?7��
?^3�?��??��A?�|f>�g�Th׾�a��	��>:�!?��\�A��L&�r�]?�Q?B��>�.����ս(Xּ���f}����?�(\?B&?ݛ��*a���¾S:�<��"�~1U�ݞ�;��D��>��>�������=F>=Ұ=�Mm�YK6�2�f<�c�=�~�>9�=�)7��n��0=,?ֿG�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �?���?Zk�?_��?�h��$=?�?S	?k"�>�J���}޾7���Pw�~x��w�]�>���>�l���K���ڙ���F��^�Žv�����>?uB>?�)�>9�>��>�Y��ݫ�'��� �7����8��g!e�;�b����|��:QU�e��$�ž���Q��>�%<�k>,�?�Xj>�Lh>%�!?Rę�݆>�+>m��>I��>�ٙ>r3s>}>^[	=sF��KR?�����'���辶���g3B?�qd?N1�>Ii�:��������?���?Ss�?&=v>h��,+��n?�>�>G��Oq
?�T:=�8��;�<V��z��I3���6��>E׽� :��M�Bnf�uj
?�/?%����̾�;׽˄���g=��?��2?ߟ-�לG�F�n��h��C���=Q�W��9�iI�z�e��������������� >�?>�?�u��:�Ҿ�����k���O���>~�>���>�C�>2�>�f���0�f�"��Vz����>{p?��>�`B?*�A?z�7?.\T?�
�> �>rz����>X<D����>4^�>�.5?�C?u8?Q�?N.?M��>����yd龈���1�>_:�>Ȑ7?Y!3?c��>4V������ه='ޚ�n��t�=7z�<��G=�zv�B����W=�i>�V?Û�ʬ8����b�j>�7?S�>l��>���,��i��<_�>1�
?�?�>� ��{r�	c�jR�>ꡂ?m��sh=��)>e��=����Ѻ	L�=x������=�����j;��y <�m�=��=b�q��C��ʍ�:�҇;7��<�t�>(�?���>�C�>�@��'� �W���e�=�Y>+S>i>Fپ�}���$��r�g��]y>�w�?�z�?7�f=��=���=�|��{U�����8������<�?BJ#?'XT?Z��?��=?Hj#?�>�*�kM���^�������?@j9?|T�>�1�
R	��A���'@�Yt�>�?�懿	��5�o�q�n�+���>W=#�e{q�Z��lZ�J��W��)�.�?��?��=�-��T!�_񨿒u���@z?3�?�X�>�<�>�(K�*����0��-�=L�?S�U?Jֶ>&�O?mUv?Ʋ^?jY>L
?���������邽B(>8U?l�?�.�?�A|?'*�>���=����׾v��pcy����4�����;�A>ѳ>J=�>nN�>��*=VE��a茽+ ����=[�m>/w�>�>��>�Cw>'�����G?��>�E�����ߤ�t����<�}�u?ʚ�?A�+?��=d��y�E��.���O�>m�?���?�7*?��S�P��=�nּ�ⶾ�q�;�>�ʹ>];�>���=LGF=4>{��>��>Z+�bX�
k8�5FM���?�F?ѱ�=5�ſ7�q���p������c<�����d�;֔���Z����=������$ĩ�\�����!�����������{����>�I�='�=�	�=�I�<�Zɼ�ռ<�tJ=f��<�G=r�o��q<|�9�l1Ȼ$^��I�*��[<�I=8��؈˾Ύ}?�:I?#�+?��C?��y>V9>�3�"��>�����A?�V>�P�)�����;�񫨾1��_�ؾUw׾��c�Eʟ��H>�kI�μ>'?3>[M�=xE�<b �=�"s=���=ȁS�=w'�=MU�=�h�=���=4�>�R>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>Β7>$>!�R�ho1�x\�a�b�MZ�@�!?8;�F̾��>M�=�߾��ƾ�q-=ƈ6>9�a=k}�,@\�=��==�{��j<=�=l=��> D>!K�=v.��շ=�J=C��=��O>w���*Y6�<%+�>u3=���=�b>�#&>��>8O?�'7?��^?��>�F��H������d�>qC>ʅ�>�Л<�e:>���>
�8?��B?��T?��>�a=�j�>��>8�&�_"g� ��������*=��?���?2�>�p��$;�d��u+��Ný?��@?��?WD�>�����ܙ"��j1���\��� =��s=�Ɗ�����Ԋ<���I���=Ϩ>uc�>Y�>t��>��h>���>�9�>�>�L=D�L=;t�*$=w�R�>>�3�=�=�9P�ǋ�<�xN=��k���Y�A�����<�ָ<�11�6��=ȴ�>��>��>`��=(@���/>{���	M�=�d��%B��d�d�~�:;/��6�e A>	BW>����$��z�?��X>Ӹ@>�{�?�u?��!>�����Ծa���f�^�V�;�=��>S�;��:��l_�3�M��zҾ���>���>��.>�CU>����E���z��оPZ`�"��>7r��<��<ՅT�������kJ����y��M��q�3?�����ǜ=��_?��n?�+�?͈?�u=!fҾFߋ>F��e��,B��3������?�**? �?3Y���.�{H̾8���޷>�@I�'�O���L�0����Kͷ�0��>������оi$3��g�������B�Mr�D��>�O?��?_:b��W��1UO�����'���q?�|g?E�>�J?�@?�&���y�r��w�=�n?ʳ�?K=�?`>�4�=t߮��r�>?�D�?>�?8�s?ցD�7U�>mD�<��%>�}���o>
�5>��=��>>�?�2?��?�ܡ�������(�%�:�\>�=��=��i>l��>:�}>��=�tJ=�5�=��G>�~�>�;�>G�y>�՘>f->�{��|K�=�	?q�4>��T>|k#?M�>r�=~�=<+Ơ<~
i���V�i��:�g��O���x�f^O<���<ڑ�>�S����?�^M>8*��M?�j�m��3�J>A�>,h��D�?t�5=(�>�3�>j��=�2�=M��>9=/>&FӾ�}>���-d!��,C��R��Ѿ�|z>��8	&�ǟ�zv���BI�mn��;g�kj�?.��6<=��ҽ<�G�?c�����k���)�X�����?�Y�>�6?ی������>(��>7ō>WI������ȍ�4h�e�?���?�;c>V�>��W?�? �1��3��tZ�/�u��&A�xe�ƺ`�g፿������
�� ����_?��x?HyA?BM�<�:z>��?��%��ӏ�L'�>/��%;�FN<=�*�>E+����`�ͮӾ͹þ�4��GF>�o?�%�?+Z?�SV���a��q>��:?q�0?~u?y�3?إ;?S�x#?g9>$?��
?P6?[/?oK?�F9>���=k��:1=񬓽����ҽ��н}&鼜�4=�y=�`����;8�=U��<32���sؼ��;���ĳ<�C=�ߣ=l��=Mا>;�]? �>���>I�6?��À5��ʪ� �.?j�'=�-������s;�����B2>�4j?#=�?W�[?b>l�?�+�A�UZ>c�>�E(>�[\>	7�>�罫�G��o=��>y�>�o�=!;��F~���	�ha��|�<� >:��>�(|>|����'>���/z���d>��Q�tɺ�3�S���G���1��v��V�>�K?k�?���=R_�o$��Gf�/)?.`<?�MM?��?'�=��۾�9���J��3���>���<�������"��l�:��˚:��s>R/������Sb>���X"߾�qn�+�I��P��P=T����R=�'��|վ&�~�X��=Xj
>�#��͕ ����;��3J?�m=�����U�cO��VO>	|�>���>!�9��-z�tt@�����P8�=b�>�$<>�昼����G�Z0��ň>(H?a6a?!�?�{���w�9�F������������?q�>[Q?�\7>��=�µ�a���ub���>��1�>���>Y����G��V�����D6'��)�>T�?>�$?RqL?g}?Nyg?h[(?�?��>iM�N���3>&?6��?�,�=/�Խ/�T�B�8�FF����>�x)?��B��͗>b�?�?}�&?zzQ?_�?��>h� �X?@�Z��>�K�>��W�a����_>�J?���>�7Y?zԃ?�>>߂5�7��橽��=�:>��2?�-#?_�?Ɨ�>N.?���]�=K�>ې|?��?��h?��<��m?�z�>�nT>m�	�X��>��%?qS?��~?*�?��F?���>
g�=���_ꂾ"����<�J�<�/�<��=BH��W���|�ྲྀی�c{�=Q��=gY�=)%�<�x:=r��=�zL=�7�>KNt>P䕾�81>��ľ*,��)LA>�У�0���⊾!�:�>��=�F�>�?k�>��#��=��>6�>�����'?��?�)?KY�;�Rb���ھc�K���>��A?ݲ�=:�l�G�����u�L�k=�n?y^?�zW�*%��C�b? �]?h��=��þնb�ˉ�C�O? �
?�G��>��~?d�q?B��>X�e�*:n�#���Cb���j��ж=Ar�>FX�@�d��?�>{�7?�N�>W�b>�%�=�u۾�w��q��X?y�?�?���??+*>~�n�P4��Q�����9]?��>I����+?]o��sѾ ��2��'�"��5��Qǚ�3���b<��[��X��R��=#�?��n?�Qt?�pc?%��u�d�%1_��΀�c^X��7���
���<��6E���@���e�R���������St@=�[p��9��i�?�R%?]�V���>���w��b�¾"�H>�����3�aKX=oǳ�/x`<���<ky�6�5��k��-?���>�[�>D">?+�a��.@�p�3��]:�o �}H>�W�>C�>�U�>�������ʍ
�K�оj1y���ͽ4�>=U\?)VE?�r?�Ӽ��5�\����$�I�ͽ�t����>��>>�Ɔ>�)��S���Re)�L�v�;����O���� �@=��?�w>Ι?���?�?u�ܾ�������uM=��#�9�5�>��W?�p�>=�>A�4��/����>,�f?h��>Ls�>]���	^ �~�s�X���>iͭ>-��>
�t>�=��Z�k(��z<��V�9�m��=�f?
Mx�:W��>�jS?&D�������>輽��$�g޾S�%��>T��>B�=B�B>�u̾�����q�7���K)?�"?|���9*� �~>�5"?�;�>�֣>�4�?ɤ�>þѼ ��?s�^?�3J?�jA?��>��=�y��țǽb�&�p�*=ls�>S�Z>ĵm=Rg�=����F\�X�u�D=�@�=`�˼n����9<�K����N<>5�<N�4>�uؿ�K�)ݾ�U����0���>ʀ� ��������%�p���Ǫ���y��-�O�Qe����5���Y�l���=e��lP�?b��?���*���*����s�6
����>�7�鹁����g�_�f��+h�ё��O��܏=��b���q��M7?�U��Ͽ	\��sf �"��>��?b7�?��Ӿ)�p��fR���>�}y>{`0=�N������zCͿ9r�*,>??����?<?*��=�o;=Ͳ?v煾H_�Xc<��?؎#?	��>����B࿦$ֿ׌��	b�?�@�|A?��(��쾈V=7��>�	?w�?>ET1��I������T�>R<�?���?�~M=d�W���	��e?�w<��F��ݻ#�=@<�=�C=^���J>�U�>ۂ�`SA�[>ܽ�4>*څ>"����^�u��<�]>��ս�;��5Մ?-{\��f���/��T��,U>��T?�*�>b:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?)�(?'ۿ��ؚ>��ܾ��M?UD6?���>�d&��t�م�=�6�&���o���&V�<��=b��>��>��,�ڋ���O��I��E��=wZ ���ǿ/a%������=ld����;̽�XG���ԽV����q��NO�+��</
+>��g>�)�>~JE>HR>�wO?�t?q��>��$-���K�I课�<=&�$�k�:�(t�������۾0 �ޔݾ�2�Ӷ$�M(�@�־D�@��L�=��C�������n�@��aj�8�'?�x�>��޾Y.F��j=>uᴾ���>�<5�>\��v�>�<g�����?&+H?|�P�I�\	о��!�Q$k�'"k?E��=���H��e��=��2>����F�>�x�=�辕�2�B1F�YT0?�H?�D��N���R)>,���=;�+?��?�]<�Ъ>�"%?��+����6;Z>]�2>�d�>J�>#�	>�Ϯ�z�۽��?�VT?���5���Z�>2���<�z��8d=�>��3�/��][>A��<<��_��q�����<�(W?s��>��)��}a�����4Y==��x?��?$.�>m{k?��B?Xդ<'h���S����aw=�W?4*i?��>����	о^���@�5?�e?z�N>�bh���:�.�^U��$?�n?4_?P~��)w}����m���n6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������^>-Ut��w�?�>�?`�Ҿ��Q�4�	�r��f �r��=�#5=V�λ��<��`��O�5���.,����I��<YU�>:@�Y|�
�?Lp���ٿ}�ȿ�9��7/� �'�Y2?�!�>=aC�@��?�N�u�e��]I�n�2���v��L�>�>����������{��q;��>��1�>����>d�S��%��b����b5<��>a��>���>�0���齾ř?9b���?ο#������ӻX?�g�?�n�?�p?hl9<U�v���{�q��-G?҉s?�Z?�z%��>]�!�7�yVk?�r�2�Y���1��f���=ʐO?���>��N�6I�=s��=8S?�>Ն#�i�˿1缿�[�si�?��?Zi�w��>��?�H?{V'�Š��g�־��]���i�OKt?)/7>~2����KE�磱���?��%?�cQ�s��D�_?�a�l�p�#�-�k�ƽ+�>³0��f\�������We����Z6y�
��?V]�?��?�����"��5%?�>󠕾=Ǿ���<�|�>q)�>C'N>7X_���u>����:��R	>���?��?�k?������T>�}?� �>u�?@��=`�>`��=����7-�!A#>��=:�>��?��M?�(�>Y��=#9��$/��[F��AR����C���>��a?�L?��a>�|����2��!�r�ͽ5'1�]%�b&@��P-�k�߽�;5>�=>��>~�D�} Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*5¿����̞�"��I� >���=ި�>5jۼp+���D�֩��99J���Q�>��>�L>D�d>c��>i<>�Q�w�'��˲��酿�p3�ґ.�IV����|��3E�U���2#�4�d˾vP��&��iͽ�����ϑ��ּ�U>�H?I�[?�i?��
?�=���=���� M=4��*|T>�wX>G�!?�C?�K"?��=�c����\�L�u�PO���Dd����>���=�-�>��>!��>�@P=쉙>�|>��C>,�y=s�;���&�>TB�>VJ�>���>H&�>֠<>�c>J��X���eB]�9Ս�ޱ`�{ʶ?C����q�C���>
.�]����d�X�T?-i&>�␿T�ؿp��`?�i�RG(�}���^�<_1?�v?�	�>�;�67��"�<��0�ݐ	�-�s>��׽���dxU����>	�J?|f>�u>�z3�F8���P�"t��vG|>26?ێ��R9��u�T�H���ݾ�iL>_V�>��H�]^��ꖿ��~��i�
Z{=��:?%^?�y��0���-v��N���@R>��\>�0=0Ԭ=�OM>ƭc�~ƽ{XH�O .=�C�=�`^>��?��0>T��=�֥>�5��HaM�歨>;�2>o�8>5=?�j?ɯ�Ѡʽ������>�,]>�a�><�k>	�>�F<���=� ?U�X>����������$���I�F+L>���?^�ϴԼP�d=����i�=�]K=P$�z*��*=�~?���(䈿��e���lD?S+?] �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��J��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>yx��Z�������u�t�#=S��>�8H?�V����O�g>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>:��?�gY?qoi>�g۾:`Z����>һ@?�R?�>�9���'���?�޶?֯�?�3i>E�?`ez?pU?��ֽQ�W�G���%[��]�ҽ��>C�
?���>����~X������+��<�t� (��9��>��@=�O�>l���<nܾЯ>H;u��*۾���=N��>H�[=U�
?O��>P�!?�B�>;��>��>VƇ=�*��&Pz�`�K?x��?O��?2n��W�<��=��^��&?zI4?�S[���Ͼը>��\?`?�[?Ld�>���%>��-迿�}�����<��K>�3�>�G�>X)���DK>H�Ծ�2D��p�>Tϗ>0����?ھ�,��8\���B�>�e!?ʓ�>�Ү=�_ ?/$?L�m>Wͳ>@�D�e��SF��D�>XH�>�P?l�?ٲ?ﺾ��3��Ւ�Vԡ���[�S�M>��x?.�?�y�>����<���o���X�>[�����?�Eg?L��)V?l%�?�>@?$�A?�Qf>����վפ��h�>d�!?�	�A�EJ&�Y��V~?P?���>a+���սA ּ�������A�?�%\?�?&?���+a�z�¾�;�<�,#��(T�`��;��D�z�>|�>����ѝ�=s>��=TNm�]K6�aqf<�{�= ��>B�=,7�{��/=,?��G�|ۃ���=��r�>xD���>�IL>����^?ml=��{�����x��!	U�� �?���?Yk�?Y��>�h��$=?�?S	?f"�>�J���}޾7���Pw�~x��w�`�>���>/�l���K���ڙ���F��^�ŽBF�u��>��>c�?HE�>�>>@��>%钾��U��E���1[��G$�}:���5�#���{���T���<����>-�����>
����>��?rC>&U>3��>I:p=���>|E=>���=�Ζ>C�>�;>��=�2�<d�۽�KR?����*�'�y��Ѳ��C3B?�qd?d1�>�i�>������w�?���?<s�?i<v>h��,+�qn?�>�>I��0q
?<U:=�-�:>�<�U�����3����Q��>�C׽� :��M�anf�jj
?�/?\����̾Y;׽J�����=3o�?s�.?�0�­Q��Kj�5']��O��z<ƚg�Wg��N�5�n�q��2��HƄ���� �#��m�=+`$?L�?"���ʺ�����Ͳk��yA�@>���>$�>�5�>�e>�#��3��P�7#����+I�>�br?F��>Q�:?��^?^S?��L?�m�>�->H�¾�?�i>.��>
��>�.?=G?#� ??]5?&�S>���?پP��}�>?9e,?��'?�A ?�?��R�1���G�U�=�"���
:��>��O������(��=��>~U?�����8�������j>�|7?���>t��>m
���+����<��>=�
?9�>h �\{r��b�FH�>2��?o���.=��)>f��=���/�Ӻ�>�=�¼e�=�_���';�J <�K�=��=Mjp����#�:܈;�b�<�m�>v�?���>nG�>�D��/� �����E�=�Y>8S>%>�Aپ8��o#����g��;y>�o�?6r�?�	g=|%�=�f�=�X��4S������ ����<u�?�B#?�XT?,��?��=?d#?ح>�#�XL���\�����N�?T�8?�I�>��"��B��z�C�1A?�`'?"�s�%�'��*���p�
E>��P��?��d+���|����>�1��Gǽa��?L��?q����<�e����L�����6:�?o��>i��>ͱ�>�1�u��A����
>�×>N\?+��>�+U?J/y?�_?���>��S�T��iە���Ƽ�>��h?Tn�?CJ�?��q?D�>*��=VE�'��~@¾b*���4� }���7T=��v>�k�>y*�>�E�>�N�=�e�)�N��(�=;Ġ>�{�>���>��>T�>l,}�`�G?��>�\������뤾 Ń�q=�՜u??ב+?U=2����E�,G��yJ�>[o�?���?�3*?[�S�~��=�ּⶾ��q�u%�>�ڹ>31�>�Ǔ=I|F=\b>a�>Y��>l(��`��q8�QM���?�F?���=I�ſ�Up���r�<'���'0<�*����h�Fƒ���S���=�晾��1�+�b�s���O됾����<w���K��7m�>��=RG�=:��=���<>7ݼX��<�VQ=0}�<��	=n�m��<��"�})��p���o�%����<Z
K=qm6������r?��J?]P+?�[E?�U�>%�>E]���o�>��]�*�#?-?>T�`���ǾDP�h���29����� ޾
�M�X5���&	>J�F�>}�i>��>�S==L��=��=Gv=R˕�u"�<�}=�@>?B�=ڜ>t_�='�=>6w?����Ʊ��J2Q��E���:?�;�>�x�=�}ƾ�@?�>>�2������5a�8.?	��?TT�?&�?oi��d�>F��U�j�=�����?2>���=��2���>��J>��PK��p���5�?-�@��??������Ͽ�^/>��>x�>��P�=�6���c��g���o��(?~�/���ȾQx>�=��ھ��Ѿ:�=� A>�`�=5��r�`���=,�)��_:=��=���>�7>껂=S���E�=��=���=u`H>�g<	o*�%�'�!=z<�=��_>�>A��>b?�1E?.�a?��>��6�\g¾�W��t�>�->��>�"�<�lH>���>�G>?��B?�>J?E�>}�K����>�o�>�h���^�C�꾝^ӾA����?��?$��>j�׼�=<���a1��
���H?��;?��?�>,����k/7�c����<���̀i=����c��J[��z�Q������;���>��>%��>���>���>պ>��>+xU>>�>�ٕ�����;{��C��=��L=�*�l{�;��<>�6�=�Ƽ5�»�ǁ=��z�`���=̽���=���>3>N��>�p�="��Dc/>������L��h�=[X���*B��-d��F~�q/�In6���B>��W>�9���.��<�?��Y>�?>���?:Au?!�>����վwG����d�*�S�ً�=ڟ>b�<�_;��H`���M�ՂҾ۪�>��>ؚ|>x?>n�h�.�F��>W�׾��F���>�a��D>
	O>�ul�ﹿ������p���μo=[?Ã|�Ԝ�=';:?��R?�Ȥ?�?��������$?������q�3qU�����v^��%?��A?�n?G�)Y��M̾���uշ>�WI�~�O�4�����0�c���·����>������о�%3�uh�������B�?r���>l�O?b�?(b�^T���WO����B���h?oxg?�)�>�I?�>?����j�"t���\�=��n?{��?c;�?]�
>8��=��̽<�>��?��?H��?xns?Ӵ?����>�<u<U)>�`ʽ^��=
>=��=N�>�?�7?�
?�I���
��m���&�f]��f=���=m�>�^�>kw>fɧ=	��<Al�=��>�ؤ>ڇ�>U�f>�(�>��>/휾j��I�?R�>i�|>��(?u#�>\�==wU�/�	=/�n��(A�L�a�� ��5�.��6��Hn�<"R�:.=�>�¿���?��>>���?�w��|��'�C>t>��ҽ���>�p9>*n>�Y�>D�>#)�=z��>�w%>]/ӾG�>��jn!��-C�&{R��Ѿ��z>���@K&�b���*��I��m���V�vj�S/��;=��<�<�G�?����Իk���)�W0����?�p�>6?�⌾r��ʦ>���>Ծ�>�"��K���Nҍ��r�3�?���?K<c>5�>��W?,�?S�1�`3�uuZ�[�u�'A��e�%�`�>፿�����
�� ���_?��x?cxA?8�<�9z>&��?W�%�	ӏ��(�>o/��';��@<=?-�>�(����`���ӾW�þ�7��FF>]�o?R%�?iY?�RV�=w=��h>7�Z?�9?��r?��??$�?u8�-�#?�u�>��"?��>$?��?��?�i>yR)>��\G���U���Y�&� 9�a&=�z�=��=��,=8~�=�м��@m�����D�=1�,<��=�n>�>>���=�§>��\?�.�>8�>>W7?.�\�8������1?�0x=��{��W�����͸�?�>��j?ZΫ?��W?��X>=?�)H�U�>�e�>��(>�d>�~�>R��(J��(�=ޮ>�i>���=ce�U���S�	�����:F�<�/>O��>�0|>�����'>���l3z�!�d>��Q��˺��S�4�G�I�1�݋v�JV�>��K?�?䐙=_�"&���Gf�f0)?�]<?,QM?��?A �=��۾��9�2�J��7���>�h�<-������^"����:�Ì�:��s>�0����#b>6���޾��n�{�I�o�羍�M=I~�u�V=L���վ3�X�=t�	>����� �����Ϫ��5J?��k=�p���JU�Rg��"�>̴�>%ۮ>�|:��{w� c@�+������=ĕ�>-�:>be��*��*YG�n9�퇇>8C?��`?�݄?����gr��VC��n��tX���눼k*?�ȡ>k? �L>�x�=k�����i�`���E��0�>�4�>���XD�k����iV$�;J�>X�?�>Ǝ?08M?��?
_?�v*?O�?��>�Ԧ��Ϯ�N�)?O��?�|�;h�Ѽ��	���@���F�x�>E�A?���Uv�>a�$?��>Z�?�bC?�>?�d>�������΁�>E]�>D�W�9���㉨>��D?Şg>5>?2cz?�r�=Om1����%��9�¼k�i>��??�;?!��>sť>t��>����Uk~=�`�>�c?�,�?�p?o��=Y
?�72>���>炖=Mן>�~�>�
?�)O?��s?��J?h.�>�%�<M䭽{���|?s�K=S�^��;��H<_�y=�N���t�}��"�<���;Wr��������(�D�����2�;&\�>b0t>�����0>�ľ���1�@>��g��ѩ����9��ʶ=��>��?I��>P7#��=jӼ>��>�����'?a�?�$?�kM;��b���ھ��K�|7�>��A?��=Q�l�v����u��<h=��m?g.^?�X������b?��]?�h�=���þF�b���龊�O?l�
?��G��>��~?3�q?��>�e��:n�����Cb���j��ж=�r�>xX�:�d�3?�>u�7?�M�>
�b>+�=�s۾
�w��q���?@�?��?���?�**>��n�"4��&��L��i�]?w��>'���"?����ϾK��1�����|������:������)f#�l+��ў޽���= ?�[s?7�p?{�_?�c �Z�c�*^���[V��W����E�N�D��MC�-	o����ȸ��`p��g�?=�.��'>��U�?��)?�k��;�>q�׾�Ӿ&)�S��>\�f��#���9=I%��>�P>~7 �c������[�?��?Z�y>,�\?2�g�ǣ.�D����8����sy�h1�>��A>O��>{��=3ע�y� ��_ӽ1�A�GxP��8v>ixc?�K?�n?�o�:)1������!�l�/��f��]�B>L`>d��>ġW�p���8&�tV>���r����&w����	��~~=;�2?S+�>Ұ�>�O�??�x	��k���]x�	�1�	��<�.�>{i?�>�>>�>zнc� ����>z�l?��>J�>v����Q!�b�{��˽���>G�>�j�>�lo>:7,���[�]�������8�J��=l�h?9�����`��ޅ>�R?GZ;c.M<(C�>�w���!�/� (��)>�?zI�=�;>Už.%���{�@���2\(?��?�����|(����>��"?�H?��>~��?ȝ>�/��ڲ�`?.�Y?��G? t9?�@�>�$�9-1ͽ1m����+�54=�z�>ÂL>R��=��=<���qs��E$��dL=cH�=J�<q�콄����aM��<��	==�>|Bٿ�M���پ��"Aݾ}�	���<�Ĉ�?�Ͻ�Ⱦ,Ο�=R��|!�����R<>����B��է��a��?ɩ�?����_���C���倿�
�t߾>�JQ���нƙ��旽�O���뾉E���a
�S]Q���S�f�b��'?ຑ���ǿȰ���9ܾ�! ?0B ?�y?���"��8�K� >�J�<�(��}�뾸�����ο���]�^?���>��1��6��>b��>8�X>�Hq>���瞾�<�<��?�-?&��>��r�:�ɿ5������<���?��@LjA?+/(��=�HuM=��>��	?�A>/Y.������a��>�&�?���?;dG=�W��6�,e?��<I�F���	��=���=Z#= ��q
J>�?�>�,�s�@�NٽoZ5>�˅>/S(��S�NA_��<�]>��ӽ���5Մ?+{\��f���/��T��U>��T?�*�>Q:�=��,?X7H�a}Ͽ�\��*a?�0�?���?$�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�م�=|6Ἆ���y���&V�{��=]��>c�>��,������O��I��b��=~ �xɿ�|$�� �⬜<�>�=1��H߽��ܽ��=�{���K���	5�l�==��=��=��>|N߽}�=>X�K?��p?��>I6>���;�ȾcѾ��/�m�����潰_Ǿz-��WϾ�ξ�'ھ�������R3���J!����={�;�i_��|&��0B���5��CC?s��<�ő�"�p��%t>�g��,	�A�q�sv�=t��!��5`�@��?\hu?(;f�]捿�VF���=68P=���?n�m�Ԙ��yr�X�>u�<�y����>�!<�w3��e�<$<�rk>?Q�=?S[��Ir��0>�$ �s`�=
P?��$?���Q,�>TmW?�˿�2z��l��>�I>�>���>�S�<o㳾z(���S?W�)?!��Ҩ�b?;9���XžD�A>��=�S���jS=�)�>�0�i��5� <#�>zjܽ�$W?B�>��)�
��"
��� �Q�;=�x?��?Rk�>=k?	C?U�<5{���S�x�
�ºz=|�W?xi?��>2䀽) о������5?N�e?��M>"nh�J�龇�.��Q�>P?N�n?�?~��}�4�����9J6?`�v?��U�	%��IE
�r�j��ʟ>���>�(?�_;��>ά4?�1�����@���8�/:�?��@Y��?�ꦼǠ)�"Yz=:Q?�A�>�PC���Ҿ���	b���7=3�>#���]t����L4��_=?��{?�n�>��~�Z�����=�7ˬ?�0�?�ͩ�:P)<W�p?j�����V	=��=7�F�? �\��Y5��p���.��-��q����>�@#���{��>��K��P῔=Ϳ24��KNξ�ۂ��?[Π>�`��a2��u�g�t+r�v�C��GC��F��qV�>�>�Ŗ�\����|��+;��x�����>W��"�>g�T��������H<��>��>��>Aè�?c�����?9p��&�Ϳ���TS���X?�8�?���?_�?T�F<�Us���z��S�
�F?�Sr?��Y?C� ��Y�3I?��j?�Z��oV`�א4�hIE��U>�"3?�I�>J�-��|=�>��>�X>&/�ލĿ�ض�@������?���?�o꾨��>́�?=u+?h��8���[��y�*���1�^=A?�2>/���͸!�/=��ɒ�2�
?}0?�z��,���^?�Xa�a�n��_-�;4Ľ#��>=12�]�Y�}����L9d�������}�
��?E&�?B�?�t��d"�i�#?@p�>����q�ľ���<U��>���>&pI>b�bVu>����A;�'>G��?�\�?�?���������>DE~?*�>��?���=Ef�>�4�=������*�{c#>�M�=�?�p�?�M?�4�>@�=��8��/�'QF�8R��"���C�N
�>��a?��L?�*b>D8��.y1�P	!��ͽ�!1�(�鼻w@�aG,��c߽�5>��=>L,>L�D�;Ӿ	�?����wؿ=���N2*��4?�߃>5�?���ett�a,#��m_?� �>�b��"��勿-P�/��?O��?L-	?[�־]ܼ�>D�>�z�>5OϽ�q��#r��;�7>.�B?Lk��p���so����>���?��@־�?�i�R	?}���V���~�B���5�*�=��8?��a�y>���>��=��u�B���Bt�fP�>��?�G�?���>��l?�=n�GQC�C<3=*�>-:k?kS?��\����rB>R,	?����R������%d?x�
@�1@K�^?~Т��,пyӓ�륻�zA־%�B<����=E	I����=N�>ś�=��>��j>(�s>Y��=��=�6<q�=���=,;���!� 6��%���� Q��f0�q�F���������e��bJ	�cs����x�H���]-���b�K��ʺ|�0)���=��T?�Q?��o?�?E�Y��C$>Ǵ��K��< '�s�=��>2?�M?S�*?���=�����d��Հ�8Ȧ����{X�>��D>EE�>�h�>z�>:3�9"�O>�@>	�>�>�=��ݻ��=hR>!ҩ>���>�ܹ>CM<>y�>bʴ�j9���h���v��̽l�?g����J�m2��N ������ƞ=�I.?�p>����)п����:H?�ϔ��2�R�+��>��0?�sW?z�>�����T�!�>נ�>k��k>-\ �l��v)��~Q>cN?~�f>]u>?�3�id8��P�%���p|>v36?m涾�-9�Y�u�y�H��gݾONM>cǾ>H�C��j�������wi�dO{=ow:?��?�#��4۰��u��C���QR>�=\>�@=�W�=�dM>C]c�]�ƽ6�G�F.=E��=ٲ^>�7?v>%�">��>n���^�u�#�>B*�=��:>�7?n�?%D��9%@���;��=�@��=[��>�G�>>B�=H=I� ԙ=��>��p>�k�=w��� ���z�챩=T,�<�x���2��$>z'�=�n�=�Ԯ<�O��VU����=�~?�~��P㈿��9C��LpD? .?���=�vF<v�"�����H��)�?�@�l�?��	�L�V���?~?�?���Z��=�w�>�ϫ>ξ�L�3�?��Ž�¢� �	�+#�,R�?W
�?��/��ʋ��l�9>V]%?ɭӾp`�>N�SX��7����u���#=,��>�EH?w\��R�O�3>�c�
?a?�p�m���2�ȿ�tv�x��>>��?A��?V�m�m?���
@��\�>-��?�rY?�yi>Eg۾�TZ�Ħ�>#�@?a�Q?]�>o<�|�'���?�ݶ?���?DI>���?��s?gl�>9x��Z/��6��ᖌ�mw=��Z;4d�>�V>�����fF�Vד��g��K�j����A�a>o�$=�>iC�#4��;�=��MI��E�f���>C,q>��I>#W�>J� ?b�>��>ep=i��Dှ����K?���?8���2n��Q�<���=Ͳ^��&?�I4?�j[�]�Ͼ�ը>ں\?d?�[?�c�>5��P>��;迿&~�����<\�K>4�>�H�>�$���FK>��Ծ�4D�Xp�>�ϗ>7����?ھ�,��KP��eB�>�e!?���>�Ү=2{ ?��#?��g>]��>-D�B0���LE�|��>�>�?h�~?�>?|I��b�2��Ē�b����Y���M>idx?-}?�=�>׏���r��g-�:�X�&���qj�?��g?yy�$?�T�?��<?~�=?
?h>�����Ծ�����>�n?�O��R�ـ!�.=Y/?Œ)?U~�>�� >��;�^%=�@����?�X?hz�>��
�r��˾e��<Y�=����J�<A����=��]>� ˽�C�=���=f_�=M�=�򽦨��y>���>+��=��i�h8S�f�,?h�;3g���8=��t�_�F��r�>2�o>�ʾE�\?#+H��]p��}���蝿�X�蟈?��?�<�?�`����g�.�6?c��?ْ?���>�.��_p޾����S�I�Y����8�= ��>%T<��о���ا��ւ���������x�>�}�>�Q?! ?keN>t^�>yҙ��&�`�𾹩��^�M����7��.�+��!����������!¾J�{��9�>'���[o�>�
?�g>�Wz>�H�>�l��[��>��Q>��>`|�>R�W>W�4>�y >��;r�˽
P?�Yþ��%�K6㾐D���HG?!�f?߉�>�j�����!g���?�X�?��?�!r>H�k�,	+��c?+U�>x|���?���<����*�<B�����N�������E�>\ӽ�9�Z7M��J`�$�
?A?��㼞TӾ����ȡ�)�f=�Ԅ?4I(?#/)���Q�ho�ʑW� �R�x�Rii��o����$��Up��я�+ۃ��B��|�)��j"=+?�_�?f�����)���Ak�ވ?��vh>�4�>M��>�վ>8�L>|	���1�k�]��&�h����>Juz?g�>ѿL?�0G?ZY[?�q1?�o>�~�>Q��M��>�D���> >�>��<?E0H?w+?�ȭ>�"0?z�>'�:��ﾋ�޾4x�>�?Y�=?A(
?���>�r��^������g�~����=LX[>Xd�=�g��:�n��CM>�?�i��}A��V�����>G[?݂?i��>/D�6c%���+>�j�>�1?#��>SG���������>�bX?�a��UI=�L_=�+Z���㼠ɓ�P�]<;� <�_&>�O�=����'���=�r=���}&=�\��Z'���hz�>�?��>�O�>�S��� ����E�=J"Y>�S>�>*پ�v��{����g�8y>,v�?R|�?Zf=s��=��=[���9�����vｾO��<5�?*2#?FjT?���?�=?�r#?��>�'��K���O��ݢ�Q�?�/?nħ>1+�]f��y���y:��y?6C"?��h�ý�/�if�QYc��7���O,���z��>�����������8�ν��?� �?��"vK��B�#������PsK?�k�>�>�7�>���F3�wN�G >�F�>�9F?u��>��P?��{?�;\?��C>-i4�\\���`��&+���
>�w5?��y?���?Drz?YH�>�>l��Ծ`J㾌.1��X �0��F=��`>�0�>��>���>�|�=���S�u���M�Z��=�Ci>��>q��>jP�>�Sr>|u��.H?���>��žz�`����у�i�l��Xs?EÐ?ν ?׭=���E�e\����>핧?���?�$?��N��N�=�9���ֺ�8�p���>���>�>�=�'A=8">u��>1V�>��������4��M�v?5�@?���=5῅~����۾{��Ȋ����D�l쐾M��ֱG��>�t�h��Cb=�����4�}��~R7�X�����ͽ���>����g�'>��9>��<("h>��@>�{�>�엽�ۯ[:��~�:S�Z�۽��=	�>>��>2y�=1>��˾Y�}?l9I?+?��C?w�y>28>�3����>����@?OV>ިP�ˊ��>�;�§������ؾlv׾8�c��ɟ�F>{dI�/�>�:3>�F�=�D�<��=-s=�=��Q��=2 �=DN�=�h�=e��=B�>zR>D�v?=����a�P��R罇�8?O��>s��=E�Ǿ��@?�A>N��>����|���~?���?���?��?�hl���>�Q���	�=w��.�3>���="E4����>�M>va��;��7寽#�?�j@}v@?r܋��iϿ\%1>�v�>�R�>}m�q%l������뇈���[?��>��r���7�=�+�>S�����{��EP>i��=�#�=�gz�n9>��m���K��7>Ǩ�>��T= u>[�4�XTr<G�=(�=t6�>�$c�����3f��M���E>h�}>��=L}�>U�?�~&?|�{?�s=���]| ��ݾ!u>�\��?H��o�=j�>`�?<?	35?_�>9ߒ>zZ�>ܗ�>~�9���H��˜�a&��"��+�Y?Cy�?١�������Ja>z7�MN��H�H5�>>H�>��h>�'
?Vn��
㿾�&��.��o��j�=ײ�=�D�����6[�,C�������>��>��>[[�>�;>�Y�=\0Q>��>I3>�OB<'�=��<�	Ӽ�����������h�=� ���󼶝��P��;s�u=��<]Z=X���x&���=�u�>��>o�>m!�=ݨ��<�1>@;���L����=�����A���c���|���.�`�7���C>��[>����q���+?/�Z>��@>1��?��t?3�>���(�־w?��q�e�5R�zm�=kV>ү:�r}:�m7`��|N��jоJ3�>���>��>4[�=��3�'q���=8X�4�Q�j?6���0M��zھ��Z��ǉ�ܜ��q>��v>���><������	�??�e?�Ŕ?�/e>�Nc��$�`A>T¼,08>��C�f{���p�>�k-?�Y?d�>������Ҿ�ν=��>QT�kjO����]�/�Q��@�n��>����nl;]�0�'<���㐿�cB���z�q��>E.M?a�?�xa�=��R�L�/b��b�l+?T�h?���>��?f�?m��Ɵ��҄�s�=f�k?K��?��?Wf>X�>�NN��ݥ>�$?��?�7�?�_�?�ꁾ��H>�����9>�W(�rv�>�6�>��>��5�q7�>�|�>�w�>]kj�w!�P
�Q�E%���>?=C1�>禨>m��>��>B�B=,U��?<��=xN�<���<~9s>�.K>գ��S ��??"f�=�u�>u�>�}�=>>��g����>۞�<�s���%��j�=��#>�T�>,[�~j�=����e�>Ğȿ:Ғ?�ȸ>�1s���`?��� ڽ�>Z�t>�Ba�R~�>��>�*>�P�>���>�O�<��:>A�>��վl�>�9��!���B��-R���ѾJx>�R���]#�8Q�62��MH��������i��V����<����<	�?<����j�
M)����i�?m�>x�6?\ތ�9G����>w��>��>����'��������ݾ�*�?�~�?�]i>EC�>��Y?�5?Y�Q��g7�)�^���u��(:�K�d�ǉZ�����l�����㉽�0a?�Uw?c#??QR�=�8s>�T~?]���K��>�E.���9�-O=r��>����%&����˾I=�������>>܌a?�ń?��?(��)��o�>�.?�1?�?j�@?iD?G~{�� ?��=�?��>g.?a5?��?�k>�_
=�M����<O��������=�/,��]�Ҍ<ۄ�< �=�2>ٚu=t6V�
�=���ONZ�=)��K��<�=sw�=���=AU�>��d?0�?c�>76�>G�W���`�OL�V5=?YG��7A �H�'����2b�+~�>�oJ?��?Y?��@?���i1���D<Yj0>�>'К>ҟ�>x(��s��>;��<Vx�=�WL>��=���+վ=P�ØU=V4Ƚ�'�>��{>o���\,>Pע���w�sla>{�T�H̹���T��#G���2�m�q��x�>�L?'�?���=E��V��Ze��B'?�j:? 3M?7o?֎�=�Jؾ��7��H��:� ��>Eά<	W�cq��RE��1z:����\�o>���������3d>���p߾Z�n��.I��I�;`R=
��b[=�D���վ3Py�ֻ�=N>4L���[ �m���ɪ�r�I?�k=J���lV�.���O>U�>��>r;���{��@�Lժ���=1E�>�\9>�q����
G�yW����>�AE? 2_?A_�?����	s��A����E��ֈ����?�;�>.�?�yA>5�=8#�����vd�O�F�nH�>c��>�%��^G�Mݞ����l$��C�>c�?�� >�? �Q?T
?`?Sq)?L�?�b�>�峽%���u&&?���?�b�=.k̽Y�T�${9�wF�=��>7�)?52D�S��>�h?0�?�c&?@�Q?�:?PD>\�����>��̕>�Ԋ>��W�#�����[>z�I?�>>%Z?8%�?,�B>i�4�Bң������P�=#�>�2?�#?�l?m9�>���>����Tǁ=��>,�b?]'�?��o?@�=��?�)2>&��>��="U�>}�>��?�PO?��s?��J?5c�>���<X­������s���E���;�L<]�y=����w�W�����<�u�;�ֺ��0��o� F��А����;4o�>���>j왾YV�=�Ծ����.>9z:<�ߒ�,7��<�P��K	>߂>���>���>��
�Y��=X��> ڴ>��� $?7J?!�?��̺kvh������J�\@�>�D?���=�_�u�����r�{��=�i?*�W?�eP����b?��]?�j�o=�k�þA�b���4�O?��
?��G���>��~?��q?���>1f�m9n����f>b���j��ݶ=�r�>!Y��d� ;�>��7?FM�>M�b>�-�=�w۾�w�;j��0?J�? �?���?�)*>��n�o3�c���$N��#�]?�L�>릾<�"?q0 �£Ͼ�>��ꎾc�᾽>���/��ݞ��=�����$�i����`ؽ�S�=�?�Fs?~Bq?۞_?�� �k�c�/Q^�i��)V�M���@�X�E�xE�pdC�(nn����*�������]H=��6�(l+�J�?3,?F�i�1� ?It����辡�0���V>�n"�:U��so>�O�<mX ��5Z>;�u�'5��}��b?xM�>��>�C?�SW��+����j-s����U�w��}�>y��>���>x	ͼ�<9��@��=ܑ�I*T�=9�� �>_<b?��G?+�m?#��r4�(]}��!���ȼῙ��B>]�=�h�>�"Q�n��zT ��7���p��o�s����n
��gR=�{,?�t�>�z�>���?�?H�
��~���Z�5�-�e�<��>�L^?���>O�>@E	��" ���>��l?5��>=�>�����[!���{���ʽt'�>��>���>N�o>J�,��"\��h��Q����9��c�=b�h?�����`��ޅ>�R?�ŉ:P�G<���>!�v�5�!�Y���'�f�>�{?���=��;>6}žL$��{�;��h�(?�?k���xI$�@&�>U�?g��>���>��?B-�>˾�����?�]?1J?��;?,)�>Y��<�i���ͽ�<'�~�R=F�>	S>w�o=�6�=��h�G��M���=pɨ=�bǼ��� w;˼cC0;6=�g6>1�׿-|H��Q���4������r蝾���AL*��Gn�ʝо){�������u�]T �M.�Ld��Q��i�|���?���?���Bಾ}?��7L��\-���>"� ��#\<f�䴙�b@[�*����y�i��6?�i<�5�N���'?{���h�ǿͯ���5ܾG" ?�B ?��y?w�o�"��8�� >~\�<�����뾉�����ο������^?G��>�
���/��>b��>ǝX>�Cq>���6鞾�\�<�?2�-?=��>�r�ڔɿ����Ա�<���?��@��8?��˾A�
��}��C1>u� ?��=e�=�� ��N�����=Zl�?�ʠ?�*��E�������1L?��g>1�f�R��=��->Ѽ�"�<(�8�a{�=��>�n:����=���Ǒ2>բ�>�qg��n�Ng�n�4>�K]>�a���=5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?:ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=u6�扤�{���&V�}��=[��>c�>,������O��I��V��=�x�,�ƿ���P�$;�=n�<�|'�� нqw��9���t;������L�b��� �=*,>&�z>H�>��6>�Y?piy?�]�>f!�=B�������g�j���(�8���ڽ�S���� �L��/��ٹ��Y�۾����MﶾX�N&s>\3���6%����8y�!?50`>_�@��x��Y��	�<�m��E�f���������������b��j�?�^?��x�����XP�d�.>�o?���<��3���JG>`*�>E��=�ȼ�|�mv�2G�{*]�k�6?�5?�`о��*����Q� �=C�M?xX�>O�>��=ۭb?��t�^�d�"d�=�Pm>���>c>	?��G�������,?Fy�?皽������>�7ƾ�|ƾ˖�><D>���܊V�:�>���>�������=�~z����mI?�A>��A��$��T:�� �=�>��a?Z%�>��L>�Z?~�:?*,]=�'�x�zf(�T�>�)V?�VU?�q3>IC�����r���xO?o�\?<n^>�0{�	�Ӿ�Z'�6��w?l�n?7K?->�M��o*��%�Ծ۔"?��v?3C^��j��l��7lW��>�O�>���>��9����>)d>?�"�jF�����G4���?ˊ@��?/4<�k�*�=�P?���>VVO���ƾo���F���%�n=�r�>Ch���`v�1��D,���8?̇�?O��>���������=O/�����?=��?t��s��<F0�ׁl�4�{w�<��=�$�����G}龁O7��������Ș�ތ��zʆ>��@�a��t�>��>����ޗͿ�����о�~�� ?{�>��Ͻ�ߦ�ͭh��0q��A�{CG���� Z�>�`>S�������D�z���:��7ڼ9��>x��3�>�(Y�����6���Bi<�|�>���>9�>6#��'���y6�?!=���nͿ X������X?i)�?ա�?��?�kj<�o�H�y������D?�-p?��X?�v!�76`�~+_�v�j?D��;T`���4��QE��U>43?�X�>��-�Q�|=��>��>�Y> #/�ߋĿ�϶�F������?$��?�d꾒��>o�?�+?Tf��=��m<���*�C��DA?�"2>�x��a�!�.=�ߧ���
?�{0?(n�'(�"�_?�a�r�p�l�-��ƽ�ڡ>��0��f\��I��1��Xe����G>y�)��?�]�?��?Y���#�6%?M�>f���M8Ǿ��<��>�)�>Q+N>{F_���u>e�7�:�Yg	>a��?,~�?-j?���-����U>��}?�O�>/�?�j�=X�?\��=⹾�!�=���=b29>/#�{�>�:?=�>�h_=�Խ+(�r(E�{Z������<�,��>`�e?�>?.�A>����˛��@%�o�W�c}��,ü��%��ؽ��#�6>��>׃>$Ч���3�?dg���ؿOk���~'��74?�ƃ>R�?=��X�t�K��)8_?w�>I�q/������#�z��?d:�?��?��׾��ͼ�>T�>�4�>R�Խ�͟�����_�7>[�B?m��1A����o�-��>���?��@	Ѯ?S�h�	?��\P��Aa~�4���6����=	�7?#.���z>~��>p�=�mv�+���H�s����>)A�?�y�?o��>��l?~o���B��1=!I�>r�k?u?_,n�]�¬B>m�?���*����O�f?��
@ou@V�^?�좿���X_�����#˾k��=y����/>����+ї<ы[=��b<+%
�8=���e>��=03�W�Ļ`ߧ=��1>��� 5'�'���������Y��P2�TQ"��XD�����KuJ���Ѿ���h�����k[�	R2������
��y>>��E?��G?��b?v�>�L�:?>�����=�m�=��C<h'�=�M?R{:?j�;?f�Z;u����S�-Lh����������g�>X�>Y׭>o�>Υ>�ʽ��*>j��=f�i>�˹��ad���=;�H�Zc>>}��>|�?U�>�C<>L�><ϴ�	2����h�Q
w�3̽6�?P���0�J��1��#9��W���th�=�a.?Z|>����>пd����2H?����_)�T�+�7�>7�0?�cW?E�>��� �T�r:>k��ݧj��_>1+ ��~l���)�Y%Q>�l?�*h>/Cv>u�2�o�6��aP�c߰�=�|>75?�K��K�5�6u�0ZH��`۾�tL>��>�M��d�[&���X~�X�i�&ez=��:?R ?be��uf����r�랾�&T>��Z>L�=�ݩ=+K>lNb��;ŽG�H�  )=���=M]>ޤ?O5n>�I>z��>����������>��=��=I?�_?��N��2��R�7��~P=wm�>��>V񞽺�{<��9��3��i��>D#J>T���T>�6�=�T�Je=0f���F����V~>��s���g<I޶<�+w�*����>�~?���#䈿��Rd���lD?]+?�=ɣF<��"�= ��hH��B�?j�@�l�?��	��V��?�@�?��G��=}�>�֫>�ξ/�L��?p�Ž+Ǣ�Ȕ	�I)#�^S�?��?��/�Qʋ�0l�t6>�^%?�Ӿ�=�>�?!��I��U���%Oh����=�p�>+A?���Y�z�X9���?s��>�d�X���vlſ;&g���>���?���?��a��$����C��(�>��?�4X?��}>�:�ur���>_*H?�\Q?*�>��"�x{$���?�2�?��?)I>V��?��s?5��>��x��d/������#7�=`�n;7Y�>#�>�����;F������d��$�j����{�a>�?$=��>���(���U�=���nJ����f���>\)q>5�I>�>� ?Pp�>�w�>�W=^������S���J�K?nV�?��BWl��<$��=�]��\?Co3?���"�Ͼ쟧>�M\?�G�?�%[?�P�>����2���v��Rߴ�?��<m�O>��>�8�>�	���K>��վ��@�8��>��>Pd��;�ھV9���}��H�>2� ?v5�>8r�=љ ?��#?�j>Q(�>1aE��9��9�E����>���>�H?��~?��?CԹ�~Z3�����桿w�[��;N>��x?V?^ʕ>a��������mE��@I�����a��?ltg?�S�0?12�?�??D�A?l)f>��ؾ]�����>j� ?����P�Jd�l����2?/�	?d�>з���Խ<U�<��#�義�?�PU?Ko?G��ug]�9U���(p<�ӣ�$�l=3�=l����>,k�=dg���>�F>)�*=�x�T�:�����>�=��>�%�=ia�g�/�d�-?���<���	�_=�lz��P�rt>�x>�fȾhl?%[�+~a��|��0���
+2�P��?��?���?3�3��^e�.�+?�u�?$?f� ?����J��}���ji����B���HYS=�w�>7��<鿾�栿ZB������)����ƽך�>���>�r?��>�*d>�	�>i=�� n޾����/
�?q������e����J�׾aX���0f�3��"b��j�>Ԟ����>v-?��>H�>j�>�dM��T>1*�=e�+>A\r>nD4>��>��=��+�0k[�o�F?��оVl��c�����<��g?uy?��?𻏼�,{�닦����>��?�׏?�zB>��r�Y�:�`??���>�J��O�>"S����=b��>>o��ڧ��^�=���>�ș>����GO��nG������I3?��D?� W�/����������n=M�?��(?�)���Q���o���W��S�M���=h�fj��i�$���p��돿{]��^$����(��f*=��*?5�?Q��������&k�?�0`f>0�><&�>�׾>&yI>��	�8�1�1^��I'�����_V�>�Y{?�S�>�;?��<?F:M?�k#?��>wG�>X�ѾFr�>}W1��D�>w;�>�
?��6?!;6?~�?r%?e�[>T������5�2��>3�?�+?�O?���>xڎ�l����_�S\�e���U붽�H=ս	= ��D��#�=DO>dD?x��gfK��~z�Sy ?�hb?ʑ#?��?&d?>C�'� �<9"S>֮ ?���>�A�����@L�V�&���[?���k��:!7?x3>�M����%�x�~=0��C����<�75�ش�>�o\>���=�!�!�o�) ;�L�l`�<�t�>k�?旊>�G�>�@��� �s���&�=��X>��R>�<>�*پ�y���&����g��y>{�?v�?�6g=��="��=X���N��d��F���i�<͞?�P#?IOT?މ�?@�=?,`#?@�>� �	F��[�������?�D-?�H�> ���Fоه��$�9�p?�?M]�f���,����������=��(�IPv�x�_5��H�/��<��`m�?�U�?DG���I<�I �W˘�߄þ2�I?���>���>��>+4"�.�U����t�M>���>-�@?ƫ�>LiN?�	v?�_?Z]�=�a;��L�������
PZ�b??G�n?�`?��v?&��>9�d>4��GR����n���W�1�!��������=_"r>Ƕ_>�<�>Ug�>v��=���;`�ͼ�텾��`=�=�>��>�J>|3�>^'|>~�߽l�F?�c�>�~���0�9Ŭ�&}z�OGN�0�t?~�?�A)?D?�<
O��@�ӌ����>P�?�g�?�(?�3_����=���d��i�Z�*��>9K�>���>f��=R`=r)>=�>vU�>Fy+�^���2���y�?Px??�,�=Hڿˠ�������벾b��<�1��Ӈ���=����=��\�2@��@�}����ȿ�l0��칗��e��'2��'s�>���=��%>�W�=xO=�T�=�c�;E_��8=���=�Ԅ��܃=�]]=��a��p)�c�=-`�=���;	����-˾�~}?�/I?R�+?�C?��x>�>�b6�K��>�4��F?�sU>��P�$r��/�:�����JR��h�ؾ�v׾d�妟�U�>��I��>;3>~��=iӄ<���=?�r=�l�=��]���=���=��=�۫=h�=o�>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?Ati��d�>M���㎽�q�=J����=2>s��=w�2�S��>��J>���K��A����4�?��@��??�ዿТϿ6a/>Sq9>E�>�7R��1��2^�f�_�Y��E!?�x:�O4ʾ̈́>
�=^�ܾ�;ȾH=H7>'5o=6;�\�&3�=jz���0=�wh=4��>��D>(��=z�����=<�G=�)�=DbS>��c�)�?�,�2�"6=�8�=��`>�'>�)�>&�(?�ZB?F=p?�0 >�%ܾy�!��#5���;�����?��.>;4<�d9>ԫ=?��B?=�u?���>���>��>���>@9�Y_A���Z�:�¾�߽�b?�?ހe>�H��-�[���,�E���!�/_?`�2?��=a�>]����	����{->��\%�ڲ>5�j<������:O�R�x��W��	~�>�i�>1�i>5�=&�=�U= ��>%E�=ʍ�˝�=�; =Ĝ,=r.K�o�>����{�=j>�:�2�f��o#��G�d��<���[���@=U��=���>��(>H��>��=ó���>?>Ϙ��6B��ڷ=����9>�{b��:s��B#��(��7>RhR>���o��
Z�>KM>��0>�_�?;�|?x�>����پHB��.�{�x?m��S�="�>M� ���5�Ryb��L�zžl!�>'۞>[�>�U>�12�סO����<�����?���?�I��� =�\�~d�Q���N��$�N��F�<��?�܅�{+�<���?�Q?�?�,�>*-9�Wy����@=r���H˹=��*��4���g=@A?9�?j�>����0��Fþx�"�>[KZ�#�D�?)��2�����E	��i)�>nh���վ,�1�8��A���bB��^�g�>a�G?\ʪ?��G�����~�X���P.���*?�Rd?#�i>�,�>!N
?��;	ؾ�����]����k?�1�?~>�?$��=�7�=�Z�����>B3?F��?�s�?�u?�7I����>cR�^(�=�.�b��=�	>���=IC�=���>�L??�O��q��G�����SY,���=�=~֠>�X�>eNH>Lي=��<Ь�=٦Y>�'�>�Gn>ӕ>-5�>kI�>\����	�)�'?���=ҏ�>��.?/"p> ��=Se�GmL=�L5��G�x�2�|%��D˽��%=�<7}E=�� ����>?ſ��?8EZ><���?�6���W�[�A>y�<>�½�'�>��I>{l>^)�>8^�>�� >�Ǌ>0F>TEӾ��>x��6o!��C�/zR�g�Ѿrz>臜���%�K��ov��aI��W���j���i�"(���*=�|.�<
J�?�,����k���)��W��-�??S�>*6?������>3��>{�>d,������-Í��S��?��?��c>�˞>�Y?�?^r6�[�/��.Z�=v��WC��3d�]��>��6W���w	��½�T`?�y?.A?��<wbz>(�?�g&�B�����>//��f:��+$=W��>���-KU�9�ξ�5ľ��D>��o?��?�?-�S�_3i��[(>��:?+�1?NUs?�1?�;?�`���$?�{5>�?�a
?��4?3/?!"?l/>��=zf\�q�$=g'��]P���ѽ��ʽѿ�]�7=I�y=�	:���;y=�Ҧ<j� �Uּ�;X���
�<619=7��=��=(��>;e?�  ?�L�>t�>s�����K������>�پ�����UE>�<��UҾ&o�>�A�?+I�?�C1?�/?F�5�_�@�d�=%m>���=�o>���>%�����F�<�~=��O=�0=$�>��%�n� �m�þ-�Ƽ�E>E�>"(z>zt���$>)���� ��̟;>�I9�Ͼ�����A�߅+��1y����>��K?IQ?���=���,��N�c��\?�A?x�H?�C~?HI	>�(־x	8���I�q�7��;�> 6м�=��R��k���07)�Af�<1`>uv��1���?d>X���k8k�p�G����)1=ݩ�M�}=���nپy)����=l�
>T���օ �`T���w����I?�{z=���� �Y�����>,�>iO�>��A��a��
>��J���ؔ=�X�>Ʀ@>㩽�� �k�E� ����>-KF?�\?�G�?��F��It�Oe?����v��r����$?���>J<�>�C�=�G>�������U�a*@����>���>�-���@��}�����٠�>K�>�v?T�'>q`�>5PB?
	�>'&W?�,-?:R�>���>K�V�L�Ⱦ�2!?π?��=@O�;��O.E�j4���>�@? Eֽa��>Y��>4�>��?��Z?�X ?쉝>����M� ��>9}Z>�6G�����>�>?\�>�z\?��y?yq>�7���پ}��ת�>l�Z�u�?S�?[�?��>0�>�	�=)��>��b?�͂?Xo?���=T�?�1>���>�ϔ=Z֞>d��>��?4O?zDs?Q�I?J,�>Rh�<�F���7���m���0�В;�=A<U�{=����wv�\=��0�<��
<�)��d�n�r�����L�͈�c�;� �>Q�>0�*��V)>��	����=ZoJ>+���zZ�1R���<;.�>�`?N@8>b���"e=�?}�/>��,��q?��"?���>�ZI>��I�ClT���v� (�>��Q?:1�=5f��!���~��In>��?gP?B�n��ě���b?}�]?Ie�=���þ}�b�����O?��
?��G���>^�~?`�q?���>'�e�9n����Cb���j��ʶ=�p�>�V���d�^C�>��7?�O�>T�b>y�=�s۾#�w��m���?a�?��?���?R(*>��n��3��(��6���^?���>ø��0�"?	����ξ����1��oQ⾭W�������֕�1t���l!�͖��C�ӽؿ=�?t�r?��q?��_?���:c� �^��U���(V��^��k��lE��D���B��n��S�s����똾�E=��_�B�6�vT�?2A3?������>�ڬ�@>Ⱦ#$վ��=_L��4�뽴,"=W��e�=�?o>r,��e*m��{@��6?��>K��>��F?��`�!���4U���j�ʋ��5f�<���>�R}>��>�l.=�	n���q=~nϾ>"���$����>�\?�0G?ߠo?�f@�^t-�Osa����Ǝx�����&#h>3#\>�K>��]�QY~�n��D�<�i�6i&�����A'�d8�=��?"��>�>78�?D8�>�l�=����[x�P�	�!�J=Q��>�j?:;�>GP>����P,�Q��>B�l?w��># �>����V!���{�� ʽ�1�>Pƭ>B��>y�o>sg,�$�[��d���x��.9��\�=��h?�r��� a��ԅ>R?�
:�ZG<�r�>�3v���!�I����'��=>�~?G5�=o;>}JžS.��{�_#���?�?r����
4���o>*=?���>Bw�>
Ņ?s%�>��ξ�'��Q?�f?'{C?E4?���>��=�%��T|�OJ���<��e>��;>��=rk=+���zz�_�$��݀=�_�=�������[&<���9�Y�<�"=	g>I�ѿY�6��¾LC$�ɗ������[�������A��=˭��Gf�8l��aJ���y!���@��^���m�\ ��I�?��@��̽J�ԾRy���p��);��'2>X��#�{=,���۾�b��V��d@N�_��RD��3��x�Y%?���x�Ŀzj��o.;�-i5?�3?��1?�0(��T׾Z�(���c��� > �	>��Ծ�s���Կ���"o?�\�>jQ������>`F>o��>(��>WM��J΍���Ž��n>�[=?HB0?a�n�HMÿ�ƺ�4ǔ=g;�?�@�>A?��n��C��f��>�$?\l�>�$n���%���;?)W�?��W?s��ȶ��͊0�O�Q?�~Իmy8���s����=R�= H�=����I=+�>��;ʫ��Q�0��N�<�x>#e^�:�(��5b�!#q>z��>�{��^F�5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=r6�����{���&V�}��=[��>d�>��,������O��I��U��=�"���Ϳe�+�����p�=e}=�@C<ޮ�^H�=ҋW=�Iž���<9P�&)ҽQ��=g"d>z�H>Π�=�bv=��Z?H�i?�>v�.>��ǽ͐A��Z׾*=&��&��LB{=*v�/х���u�y7پ����^оn��<ﾝ.����4�_�>P�A�*��g���L�̷R�~�
?�Ԇ>�PJ�8YU�'1�t���?�kg�ߋ��Rթ���bG��Ɯ?��G?	=���eY�r���%	=�	/��fF?	���������Yd�<}�<���=�)�>�4o=��ʾF���t6�X�1?Z�?����Y�"�uh��6E��=\�(?�?~���v�>��?�)����/D#>E~w> �y>س�>>��=�ĝ����ͳ?p1J?��<�y����>rO���j��w��N�>��J%9��{>���=W.�aw��z���s��{N?9�>�B*�Dg8����6\='aݼ&{?<f?zň>��F?NZ4?��>/qʾ��]�������={�T?�dO?�'&>��ѽ��þu�b�Z&?�N?H�t>ի��B�о&�S������&?��z?�|-?̨�8������5;߾�&?��v?�q^��s�������V��A�>�^�>���>��9�lm�>��>?�#��G��M����\4����?��@΋�?֘;<�%����=4;?|Y�>��O�~?ƾ�y���~��Euq=��>�����cv�X���W,�[�8?N��?��>L���y����=�ӄ��e�?�Í?�־:�]<G�#���v�0�������H�="�̼d���a��2���;%�+��\)��5�-�q>}�@��1�t��>���
]ٿS"̿�_����	�����"?j��>p����ĕ�:B�t�[� 4���L�Ws���L�>C�d>�ͽ�P�	o� � |�q��>�!=xq�>�߅���ܾ�[��[=i�p>� �>CØ>�������]�?�Aܾ�kſ{ꖿ��fvV?���?�<�?�?Z�޽0�Q2(��ٱ=8c@?	�H?��@?ip>���<�L�|��9d?���$a���,���4���><�A?�j�>���Efb<��9>C"	?�R>5I=���ſ�]���H�C�?��?'�ξr��>�W�?h!?k�y6����־��)��ʑ==]^?��>D���?,��52����`��>�)?����0&���_?�a���p���-�Ktƽ��>��0��|\�*^��|��Le�n��Fy� ��?LZ�?\�?����	#�04%?��>g����CǾ�*�<"{�>�(�>,N>�_�Ѭu>5�C�:�^	>I��??z�?�c?��������^>��}?��>���?���=D��>/�=�Z��9V˻� >�*�=Z�C�}?5N?��>�=��2���-�]�F�?R��l	��&C�~]�>.�`?IK?g>�ǯ�+)�f!��f۽f0���߼"�9�/�&���۽D�8>�8>cn>�F��%Ծ��!?����.ѿ�Ӎ�8����A?���>�~�>�D¾�/��Q>��^?c7.>�($��w��U����VS���?�M�?oo?Ey�����Bk�=h$�>�t>׋9�	�齒��&��>u�i?��i� i����Y��N><��?��@m��?k��	?��_T���U~��h�=l6�/x�=5�7?��f{>:;�>�)�={zv�y�����s��[�>�2�?�h�?$��>ߙl?�bo���B��T1=�s�>Ѕk?\g?�0h��!�C�B>t�?���O���0R���e?��
@ku@1N^?�碿ъѿʔ�����\����u�=��=@BK>o×����=�ѐ=�l<ߏƽ��B=�s�>U�>5�{>��N>n�>3�=�m��J9'�V
��ǚ�)�>������4W�fu�oLZ�
�G���F� ����򸽺락��O��ᐾ�j˽�]>�N?��N?��l?a�> q���m>�P�*HN����Y��=���>U|?�WA?Η<?��<��ƾ��`����设�>��S�>�s�=?�?���>�}�>{+���L�=m;>��U>I�>͎�=؉�= B?=�8�=t��>P��>�g�>�o<>��>㰴�����V�g�U�t�9�ǽ֬�?�\��>J��ϕ�g�������1q�=�0.?�4>4��SпX���s�G?��������+�W�>e0?%�V?�>e=��>�K���>�}
���j���>_z����m�x*���O>��?g>��t>�3��58�P�P��>��^�|>�6?�ڶ���8�bu�i�H��MݾJYM>ڕ�>�V@��e�k���B�~��+i�'�y=�.:?w?^����c�u��K����Q>�2\>��=&��=4M>��`��Ž�H���)=��=�_>�?7J>���<��>I��]Zb�Y��>(a�>d��>�V?6#?x-��"K0�����{��^=�>�r�>R��<fB=brK�D��� �?��}>8��� �Ͻ��H��.F�=�y�����>g=���=�tx�I�>3b>g���&��nP���|?q~��N�����\ˈ��H?S�?�P=+�i��E�����X0�?��@"��?/��iBZ��K?-�?�E��^��=a��>��>Zо.P;�G�?zh�����������/���?_J�?O�N�^����m�f� >��+?�?ʾMp�>�5��S��&��N�u���&=(��>�1H?���P�*=>�vj
? 0?�*�٪����ȿ7_v����>���?�?h�m��.��=�?���>��?4NY?�	j>J%۾2[�(r�>��@?�R?�;�>TH��(�a�?�Ͷ?w��?'I>≑?��s?Ej�>�v��_/�E,�������=�h\;,}�>r>"���_F�ؽ��lY��_�j�����a>w'%=�>��佾H��$��=�ڋ�}4��#ie��z�>�"q>��I>�F�>�� ?�0�>�Ù>�=�o���	���Җ���K?A��?���+n����<(��=٣^��#?�F4?t�[���Ͼ�ܨ>��\?9��?[?�b�>���J=���翿�}���w�<_�K>u0�>EK�>x���NK>��ԾjCD��m�><З>H���];ھ�*��]롻�<�>0b!?q��>W��=�� ?�#?�Xj>y��>�_E�*��k�E�X��>f��>.D?<�~?��?����T3��	���㡿��[��cN>=�x?KT?�>K����y��g�G�i)I�����k��?�lg?�彷?�.�?�??�A?R�e>�����׾���;ր>�R?��4��MG�Y.���=eq?�k?ua�>m~����=H�>g�9�p��]�?�K?�� ?x�-�:���ٹ;��s=o͋�4�_����<�<���r=��<=5�,:#=:f�>0��=b��������9>^>�Ɂ=A ���Rgv>�b*?�j'�6B}����=c2q���D�:�{>�AU>C�����^?%sE��z�����������L�n��?9��?���?����T�h��l9?��?E(?���>�^��pݾ���w,f�(�x�y*��`>�}�>	����޾{���⨿�݄��}��n�����>�$�>+?���>j�K>���>{h��f�%��~��9��^�^��Uk8�_-��#��������@�Ʊ¾��~��R�>U�aD�>��?O~f>�Yy>��>�3�I��>�1R>W&~>��>TuZ>"6>���=_�6:�ɽQIJ?處�7'��,������J:?��???�j������e ���#?炥?j�?A�=3;s������?�O�>��t�&p�>LId>-�>�:������ɽ��=� �<�c>�n%�1�+�-G���B���?9y�>�oX���+�	�N�􎠾�o=�L�?��(?�)�<�Q�h�o���W��S��T�]?h��k����$�"�p�쏿�]��j#���(��|*=Ћ*?��?���:��B$���$k��?��Wf>��>n&�>�ܾ>�[I>��	�m�1���]�iL'�纃��T�>7]{?"Ŋ>��H?��>?�P?6�I?���>�>���_��>�}y��D�>���>�
3?-U*?�M1?1!?�Y-?�g>�ܽ.�����پ�?|J?m�?��?��?i����j��}̼��$��o��i����t=���<�LོX��|E=2S>�?�n���L��¾c&�>/f�?,�H?�!�>۵�5ʾ������>$;?E	B>v���D���'��M�>fϖ?��ؽ�g���a>{zC�@�/��d�B��=�#m>�^#>S�d�X'w=�ac>�w�;B���[���Ｚ�1=״p>R��N�>��?H��>�0�>�ㅾm� ������=�Y>S>8�>�Eپ�q��J����g�Cuy>�n�?[g�?�f=�N�=7}�=�⠾�~���������O��<�?�#?g"T?���?@�=?�Z#?J>���<��<V��90���l?&)?Jt�>�8�ZL¾2L���.9��_�>I?
5_��S�8�1���*_=�bu>�8�R��{����q�ͽ9���׽j}�?`Y�?m�» ^�>M������q���kL?`c�>�5N>4��>,�$���H���Ͻ>Hs�>�a5?�I�>�Z?ZI�?t h?1�>�sF��a������3�;Ī
�"?m�\?q��?��h?�6 ?���>i�����;@AGY����~���K����v�>��}>p��>Z�>O�	>����Q>1��a��_�=���>mƹ>�*i>���>�0W>BG�=��.?cQ?�V����8�vV��͗7�8AZ��E?��?)I?�¼��:�~..��O߾}E�>��?���?b*?gW&��5C>R`)�w�վ�]���J[>GA�>��>J�>������<�[�>���>�wJ��� ���D�d23<"�?+/*?���А߿O���el¾(��x�<������ ����;�
7�E�>�G�����<���������8��#f��羾����g��LQ�>�T=`+>(>��f�T}��T�R=ƨ�=Q��=4=��\'>���=�*�K�z��N�<9
���">M��=q�˾�}?[8I?d�+?i�C?o�y>�7><k3�r��>Ռ��lC?cV>��P����Mw;������ �ؾzw׾�c��Ɵ��;>�^I���>f73>3K�=*��<+	�=�s=;��=�O��L=�%�=�c�=NM�=<��=G�>�D>e6w?蚁�X����3Q��U罧�:?29�>���=�ƾ�@?��>>
2��+����b�!,?���?6T�?$�?fvi�d�>���Վ��w�=����62>���=��2����>��J>q���J���{���4�?��@m�??�ዿR�Ͽ�_/>�
`>�e�=��I��J(���7��X���D��x*?��0�(�¾p��>�=�'Ծ�ؽ��ka=�+=>��Z=K0��gX�4�=�-��"|=���=���>yN>���=�攽�=n@2=,�=��l>�^=�����o��G<6x=�1`>V0�=� �>Ӛ!?�3?Z�_?*��>�D��v�������Y>�;���>D$=ab=a�l>��L?�n:?,�F?,��>fwd=���>��>}�/�a���6џ���;��z?�t?F�>����W�j�	�!���X���>�t/?)��>�\>2/�Q�C�/��J(��T6�*y=��=��۽0�#=VEq���C�mL
>s>��0>�8�>�2�>\>, {=J��=h��>F�=�[=�'> m����=�I����_�D��= @K>y�*��b,=�L=]��* ��`�=X�d;�&�=�w�. �=���>��Z>�6�>l��<M�Ծ�>��/���C�� >x὾�8��Wc�δr����	�ؽ�b>�R�>�G��(����>,�>��f>���?�w�?q�!>n.�PJz�Bm���k���OD���<�P�=8���*��RD�w X�Xy�����>���>)�>b>?�7�\iL�=V=ѭ�}eI�`�>I㏾ڰY��`۽��_�����^��(�\�n}�=�.?�Ȉ�M٣=�^�?�,=?���?���>�(��)QھOJB>=�l�<�=�~F����P�&?�2?,(�>Ԋ�G-�E̾.����η>&�I�c�O�����D�0�T������~��>;����о3��\�����ƅB�,r����>��O?K�?�b�JT���VO�����څ�c?zwg?,�>D?NB? 9���d�����h�=��n?Ԭ�?P3�?��
>���=h&��9#�>{d?���?f��?I�s?h?��1�>��u;22>ݣ��*��=/�>���=�U�=�#?
?�-?�\���n	�z{���3`���<y��=���>�3�>�^n>+��=��f=�!�=7xZ>���>�r�>;2d>XV�>���>�ݡ����9?��,>+�u>�M?0�R>�>*ȸ��yP=���/jJ���>�T������1�=�%<^��=��=��>~�¿�T�?z>7v�O�,?)��mC��{>��[=&�k����>`�^>u�S>���>Xշ>�|z�[P>w�Z>Ӿ�>����!��B��%R�u�ѾmMy>KQ��FS$��;w��S�H�aq���=���i�l#���+=� o�<�6�?2{��ϳk�Q�)�����^�?bը>��5?����Ҽ��+o>�t�>�.�>����[k�������Kᾮ�?���?4_>��>�Nd?��"?�v=���E��9a�FG{�x�I�Ueh��K�ql����r���	�d{ ��'j?a9n?�}6?&��<�c>\�?��(��쎾J�>�8��=���/=�(�>����X�c���ɾ9ζ��jｇ�i>�X?�/�?1�?�+��X�5#>�n9?�0?��s?M�0?��:?ץ�	�#?�P1>��?L�
?��4?{
.?��
?X2>,��=����-�=.����鉾Y,ս��Ž���,A=�(�=$��8v�	<ɭ=	�<F¼	\���^;O�����<�\/=_j�=���=���>�f?X$?��>9�;?��ϾI,L�����Z?7��=,���q����	�"�T�q>ә]?�v�?�(-?Zg�>+������/��
>�>e�.>#8�>5O�hM�����=��k>$��=5i������݊����#x��m�=t�<���>��|>�3��� )>?��s�z��4e>@�Q�/�����S�SBG��o1��w�.��>��K?*�?P�=�/�\1��!f���(?�R<?��L?>�?���=��ھ	:���J����Rȟ>�W�<���=l��M����";��69�&s>"+����#b>6���޾��n�{�I�o�羍�M=I~�u�V=L���վ3�X�=t�	>����� �����Ϫ��5J?��k=�p���JU�Rg��"�>̴�>%ۮ>�|:��{w� c@�+������=ĕ�>-�:>be��*��*YG�n9�퇇>8C?��`?�݄?����gr��VC��n��tX���눼k*?�ȡ>k? �L>�x�=k�����i�`���E��0�>�4�>���XD�k����iV$�;J�>X�?�>Ǝ?08M?��?
_?�v*?O�?��>�Ԧ��Ϯ�N�)?O��?�|�;h�Ѽ��	���@���F�x�>E�A?���Uv�>a�$?��>Z�?�bC?�>?�d>�������΁�>E]�>D�W�9���㉨>��D?Şg>5>?2cz?�r�=Om1����%��9�¼k�i>��??�;?!��>sť>t��>����Uk~=�`�>�c?�,�?�p?o��=Y
?�72>���>炖=Mן>�~�>�
?�)O?��s?��J?h.�>�%�<M䭽{���|?s�K=S�^��;��H<_�y=�N���t�}��"�<���;Wr��������(�D�����2�;&\�>b0t>�����0>�ľ���1�@>��g��ѩ����9��ʶ=��>��?I��>P7#��=jӼ>��>�����'?a�?�$?�kM;��b���ھ��K�|7�>��A?��=Q�l�v����u��<h=��m?g.^?�X������b?��]?�h�=���þF�b���龊�O?l�
?��G��>��~?3�q?��>�e��:n�����Cb���j��ж=�r�>xX�:�d�3?�>u�7?�M�>
�b>+�=�s۾
�w��q���?@�?��?���?�**>��n�"4��&��L��i�]?w��>'���"?����ϾK��1�����|������:������)f#�l+��ў޽���= ?�[s?7�p?{�_?�c �Z�c�*^���[V��W����E�N�D��MC�-	o����ȸ��`p��g�?=�.��'>��U�?��)?�k��;�>q�׾�Ӿ&)�S��>\�f��#���9=I%��>�P>~7 �c������[�?��?Z�y>,�\?2�g�ǣ.�D����8����sy�h1�>��A>O��>{��=3ע�y� ��_ӽ1�A�GxP��8v>ixc?�K?�n?�o�:)1������!�l�/��f��]�B>L`>d��>ġW�p���8&�tV>���r����&w����	��~~=;�2?S+�>Ұ�>�O�??�x	��k���]x�	�1�	��<�.�>{i?�>�>>�>zнc� ����>z�l?��>J�>v����Q!�b�{��˽���>G�>�j�>�lo>:7,���[�]�������8�J��=l�h?9�����`��ޅ>�R?GZ;c.M<(C�>�w���!�/� (��)>�?zI�=�;>Už.%���{�@���2\(?��?�����|(����>��"?�H?��>~��?ȝ>�/��ڲ�`?.�Y?��G? t9?�@�>�$�9-1ͽ1m����+�54=�z�>ÂL>R��=��=<���qs��E$��dL=cH�=J�<q�콄����aM��<��	==�>|Bٿ�M���پ��"Aݾ}�	���<�Ĉ�?�Ͻ�Ⱦ,Ο�=R��|!�����R<>����B��է��a��?ɩ�?����_���C���倿�
�t߾>�JQ���нƙ��旽�O���뾉E���a
�S]Q���S�f�b��'?ຑ���ǿȰ���9ܾ�! ?0B ?�y?���"��8�K� >�J�<�(��}�뾸�����ο���]�^?���>��1��6��>b��>8�X>�Hq>���瞾�<�<��?�-?&��>��r�:�ɿ5������<���?��@LjA?+/(��=�HuM=��>��	?�A>/Y.������a��>�&�?���?;dG=�W��6�,e?��<I�F���	��=���=Z#= ��q
J>�?�>�,�s�@�NٽoZ5>�˅>/S(��S�NA_��<�]>��ӽ���5Մ?+{\��f���/��T��U>��T?�*�>Q:�=��,?X7H�a}Ͽ�\��*a?�0�?���?$�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�م�=|6Ἆ���y���&V�{��=]��>c�>��,������O��I��b��=~ �xɿ�|$�� �⬜<�>�=1��H߽��ܽ��=�{���K���	5�l�==��=��=��>|N߽}�=>X�K?��p?��>I6>���;�ȾcѾ��/�m�����潰_Ǿz-��WϾ�ξ�'ھ�������R3���J!����={�;�i_��|&��0B���5��CC?s��<�ő�"�p��%t>�g��,	�A�q�sv�=t��!��5`�@��?\hu?(;f�]捿�VF���=68P=���?n�m�Ԙ��yr�X�>u�<�y����>�!<�w3��e�<$<�rk>?Q�=?S[��Ir��0>�$ �s`�=
P?��$?���Q,�>TmW?�˿�2z��l��>�I>�>���>�S�<o㳾z(���S?W�)?!��Ҩ�b?;9���XžD�A>��=�S���jS=�)�>�0�i��5� <#�>zjܽ�$W?B�>��)�
��"
��� �Q�;=�x?��?Rk�>=k?	C?U�<5{���S�x�
�ºz=|�W?xi?��>2䀽) о������5?N�e?��M>"nh�J�龇�.��Q�>P?N�n?�?~��}�4�����9J6?`�v?��U�	%��IE
�r�j��ʟ>���>�(?�_;��>ά4?�1�����@���8�/:�?��@Y��?�ꦼǠ)�"Yz=:Q?�A�>�PC���Ҿ���	b���7=3�>#���]t����L4��_=?��{?�n�>��~�Z�����=�7ˬ?�0�?�ͩ�:P)<W�p?j�����V	=��=7�F�? �\��Y5��p���.��-��q����>�@#���{��>��K��P῔=Ϳ24��KNξ�ۂ��?[Π>�`��a2��u�g�t+r�v�C��GC��F��qV�>�>�Ŗ�\����|��+;��x�����>W��"�>g�T��������H<��>��>��>Aè�?c�����?9p��&�Ϳ���TS���X?�8�?���?_�?T�F<�Us���z��S�
�F?�Sr?��Y?C� ��Y�3I?��j?�Z��oV`�א4�hIE��U>�"3?�I�>J�-��|=�>��>�X>&/�ލĿ�ض�@������?���?�o꾨��>́�?=u+?h��8���[��y�*���1�^=A?�2>/���͸!�/=��ɒ�2�
?}0?�z��,���^?�Xa�a�n��_-�;4Ľ#��>=12�]�Y�}����L9d�������}�
��?E&�?B�?�t��d"�i�#?@p�>����q�ľ���<U��>���>&pI>b�bVu>����A;�'>G��?�\�?�?���������>DE~?*�>��?���=Ef�>�4�=������*�{c#>�M�=�?�p�?�M?�4�>@�=��8��/�'QF�8R��"���C�N
�>��a?��L?�*b>D8��.y1�P	!��ͽ�!1�(�鼻w@�aG,��c߽�5>��=>L,>L�D�;Ӿ	�?����wؿ=���N2*��4?�߃>5�?���ett�a,#��m_?� �>�b��"��勿-P�/��?O��?L-	?[�־]ܼ�>D�>�z�>5OϽ�q��#r��;�7>.�B?Lk��p���so����>���?��@־�?�i�R	?}���V���~�B���5�*�=��8?��a�y>���>��=��u�B���Bt�fP�>��?�G�?���>��l?�=n�GQC�C<3=*�>-:k?kS?��\����rB>R,	?����R������%d?x�
@�1@K�^?~Т��,пyӓ�륻�zA־%�B<����=E	I����=N�>ś�=��>��j>(�s>Y��=��=�6<q�=���=,;���!� 6��%���� Q��f0�q�F���������e��bJ	�cs����x�H���]-���b�K��ʺ|�0)���=��T?�Q?��o?�?E�Y��C$>Ǵ��K��< '�s�=��>2?�M?S�*?���=�����d��Հ�8Ȧ����{X�>��D>EE�>�h�>z�>:3�9"�O>�@>	�>�>�=��ݻ��=hR>!ҩ>���>�ܹ>CM<>y�>bʴ�j9���h���v��̽l�?g����J�m2��N ������ƞ=�I.?�p>����)п����:H?�ϔ��2�R�+��>��0?�sW?z�>�����T�!�>נ�>k��k>-\ �l��v)��~Q>cN?~�f>]u>?�3�id8��P�%���p|>v36?m涾�-9�Y�u�y�H��gݾONM>cǾ>H�C��j�������wi�dO{=ow:?��?�#��4۰��u��C���QR>�=\>�@=�W�=�dM>C]c�]�ƽ6�G�F.=E��=ٲ^>�7?v>%�">��>n���^�u�#�>B*�=��:>�7?n�?%D��9%@���;��=�@��=[��>�G�>>B�=H=I� ԙ=��>��p>�k�=w��� ���z�챩=T,�<�x���2��$>z'�=�n�=�Ԯ<�O��VU����=�~?�~��P㈿��9C��LpD? .?���=�vF<v�"�����H��)�?�@�l�?��	�L�V���?~?�?���Z��=�w�>�ϫ>ξ�L�3�?��Ž�¢� �	�+#�,R�?W
�?��/��ʋ��l�9>V]%?ɭӾp`�>N�SX��7����u���#=,��>�EH?w\��R�O�3>�c�
?a?�p�m���2�ȿ�tv�x��>>��?A��?V�m�m?���
@��\�>-��?�rY?�yi>Eg۾�TZ�Ħ�>#�@?a�Q?]�>o<�|�'���?�ݶ?���?DI>���?��s?gl�>9x��Z/��6��ᖌ�mw=��Z;4d�>�V>�����fF�Vד��g��K�j����A�a>o�$=�>iC�#4��;�=��MI��E�f���>C,q>��I>#W�>J� ?b�>��>ep=i��Dှ����K?���?8���2n��Q�<���=Ͳ^��&?�I4?�j[�]�Ͼ�ը>ں\?d?�[?�c�>5��P>��;迿&~�����<\�K>4�>�H�>�$���FK>��Ծ�4D�Xp�>�ϗ>7����?ھ�,��KP��eB�>�e!?���>�Ү=2{ ?��#?��g>]��>-D�B0���LE�|��>�>�?h�~?�>?|I��b�2��Ē�b����Y���M>idx?-}?�=�>׏���r��g-�:�X�&���qj�?��g?yy�$?�T�?��<?~�=?
?h>�����Ծ�����>�n?�O��R�ـ!�.=Y/?Œ)?U~�>�� >��;�^%=�@����?�X?hz�>��
�r��˾e��<Y�=����J�<A����=��]>� ˽�C�=���=f_�=M�=�򽦨��y>���>+��=��i�h8S�f�,?h�;3g���8=��t�_�F��r�>2�o>�ʾE�\?#+H��]p��}���蝿�X�蟈?��?�<�?�`����g�.�6?c��?ْ?���>�.��_p޾����S�I�Y����8�= ��>%T<��о���ا��ւ���������x�>�}�>�Q?! ?keN>t^�>yҙ��&�`�𾹩��^�M����7��.�+��!����������!¾J�{��9�>'���[o�>�
?�g>�Wz>�H�>�l��[��>��Q>��>`|�>R�W>W�4>�y >��;r�˽
P?�Yþ��%�K6㾐D���HG?!�f?߉�>�j�����!g���?�X�?��?�!r>H�k�,	+��c?+U�>x|���?���<����*�<B�����N�������E�>\ӽ�9�Z7M��J`�$�
?A?��㼞TӾ����ȡ�)�f=�Ԅ?4I(?#/)���Q�ho�ʑW� �R�x�Rii��o����$��Up��я�+ۃ��B��|�)��j"=+?�_�?f�����)���Ak�ވ?��vh>�4�>M��>�վ>8�L>|	���1�k�]��&�h����>Juz?g�>ѿL?�0G?ZY[?�q1?�o>�~�>Q��M��>�D���> >�>��<?E0H?w+?�ȭ>�"0?z�>'�:��ﾋ�޾4x�>�?Y�=?A(
?���>�r��^������g�~����=LX[>Xd�=�g��:�n��CM>�?�i��}A��V�����>G[?݂?i��>/D�6c%���+>�j�>�1?#��>SG���������>�bX?�a��UI=�L_=�+Z���㼠ɓ�P�]<;� <�_&>�O�=����'���=�r=���}&=�\��Z'���hz�>�?��>�O�>�S��� ����E�=J"Y>�S>�>*پ�v��{����g�8y>,v�?R|�?Zf=s��=��=[���9�����vｾO��<5�?*2#?FjT?���?�=?�r#?��>�'��K���O��ݢ�Q�?�/?nħ>1+�]f��y���y:��y?6C"?��h�ý�/�if�QYc��7���O,���z��>�����������8�ν��?� �?��"vK��B�#������PsK?�k�>�>�7�>���F3�wN�G >�F�>�9F?u��>��P?��{?�;\?��C>-i4�\\���`��&+���
>�w5?��y?���?Drz?YH�>�>l��Ծ`J㾌.1��X �0��F=��`>�0�>��>���>�|�=���S�u���M�Z��=�Ci>��>q��>jP�>�Sr>|u��.H?���>��žz�`����у�i�l��Xs?EÐ?ν ?׭=���E�e\����>핧?���?�$?��N��N�=�9���ֺ�8�p���>���>�>�=�'A=8">u��>1V�>��������4��M�v?5�@?���=5῅~����۾{��Ȋ����D�l쐾M��ֱG��>�t�h��Cb=�����4�}��~R7�X�����ͽ���>����g�'>��9>��<("h>��@>�{�>�엽�ۯ[:��~�:S�Z�۽��=	�>>��>2y�=1>��˾Y�}?l9I?+?��C?w�y>28>�3����>����@?OV>ިP�ˊ��>�;�§������ؾlv׾8�c��ɟ�F>{dI�/�>�:3>�F�=�D�<��=-s=�=��Q��=2 �=DN�=�h�=e��=B�>zR>D�v?=����a�P��R罇�8?O��>s��=E�Ǿ��@?�A>N��>����|���~?���?���?��?�hl���>�Q���	�=w��.�3>���="E4����>�M>va��;��7寽#�?�j@}v@?r܋��iϿ\%1>�v�>�R�>}m�q%l������뇈���[?��>��r���7�=�+�>S�����{��EP>i��=�#�=�gz�n9>��m���K��7>Ǩ�>��T= u>[�4�XTr<G�=(�=t6�>�$c�����3f��M���E>h�}>��=L}�>U�?�~&?|�{?�s=���]| ��ݾ!u>�\��?H��o�=j�>`�?<?	35?_�>9ߒ>zZ�>ܗ�>~�9���H��˜�a&��"��+�Y?Cy�?١�������Ja>z7�MN��H�H5�>>H�>��h>�'
?Vn��
㿾�&��.��o��j�=ײ�=�D�����6[�,C�������>��>��>[[�>�;>�Y�=\0Q>��>I3>�OB<'�=��<�	Ӽ�����������h�=� ���󼶝��P��;s�u=��<]Z=X���x&���=�u�>��>o�>m!�=ݨ��<�1>@;���L����=�����A���c���|���.�`�7���C>��[>����q���+?/�Z>��@>1��?��t?3�>���(�־w?��q�e�5R�zm�=kV>ү:�r}:�m7`��|N��jоJ3�>���>��>4[�=��3�'q���=8X�4�Q�j?6���0M��zھ��Z��ǉ�ܜ��q>��v>���><������	�??�e?�Ŕ?�/e>�Nc��$�`A>T¼,08>��C�f{���p�>�k-?�Y?d�>������Ҿ�ν=��>QT�kjO����]�/�Q��@�n��>����nl;]�0�'<���㐿�cB���z�q��>E.M?a�?�xa�=��R�L�/b��b�l+?T�h?���>��?f�?m��Ɵ��҄�s�=f�k?K��?��?Wf>X�>�NN��ݥ>�$?��?�7�?�_�?�ꁾ��H>�����9>�W(�rv�>�6�>��>��5�q7�>�|�>�w�>]kj�w!�P
�Q�E%���>?=C1�>禨>m��>��>B�B=,U��?<��=xN�<���<~9s>�.K>գ��S ��??"f�=�u�>u�>�}�=>>��g����>۞�<�s���%��j�=��#>�T�>,[�~j�=����e�>Ğȿ:Ғ?�ȸ>�1s���`?��� ڽ�>Z�t>�Ba�R~�>��>�*>�P�>���>�O�<��:>A�>��վl�>�9��!���B��-R���ѾJx>�R���]#�8Q�62��MH��������i��V����<����<	�?<����j�
M)����i�?m�>x�6?\ތ�9G����>w��>��>����'��������ݾ�*�?�~�?�]i>EC�>��Y?�5?Y�Q��g7�)�^���u��(:�K�d�ǉZ�����l�����㉽�0a?�Uw?c#??QR�=�8s>�T~?]���K��>�E.���9�-O=r��>����%&����˾I=�������>>܌a?�ń?��?(��)��o�>�.?�1?�?j�@?iD?G~{�� ?��=�?��>g.?a5?��?�k>�_
=�M����<O��������=�/,��]�Ҍ<ۄ�< �=�2>ٚu=t6V�
�=���ONZ�=)��K��<�=sw�=���=AU�>��d?0�?c�>76�>G�W���`�OL�V5=?YG��7A �H�'����2b�+~�>�oJ?��?Y?��@?���i1���D<Yj0>�>'К>ҟ�>x(��s��>;��<Vx�=�WL>��=���+վ=P�ØU=V4Ƚ�'�>��{>o���\,>Pע���w�sla>{�T�H̹���T��#G���2�m�q��x�>�L?'�?���=E��V��Ze��B'?�j:? 3M?7o?֎�=�Jؾ��7��H��:� ��>Eά<	W�cq��RE��1z:����\�o>���������3d>���p߾Z�n��.I��I�;`R=
��b[=�D���վ3Py�ֻ�=N>4L���[ �m���ɪ�r�I?�k=J���lV�.���O>U�>��>r;���{��@�Lժ���=1E�>�\9>�q����
G�yW����>�AE? 2_?A_�?����	s��A����E��ֈ����?�;�>.�?�yA>5�=8#�����vd�O�F�nH�>c��>�%��^G�Mݞ����l$��C�>c�?�� >�? �Q?T
?`?Sq)?L�?�b�>�峽%���u&&?���?�b�=.k̽Y�T�${9�wF�=��>7�)?52D�S��>�h?0�?�c&?@�Q?�:?PD>\�����>��̕>�Ԋ>��W�#�����[>z�I?�>>%Z?8%�?,�B>i�4�Bң������P�=#�>�2?�#?�l?m9�>���>����Tǁ=��>,�b?]'�?��o?@�=��?�)2>&��>��="U�>}�>��?�PO?��s?��J?5c�>���<X­������s���E���;�L<]�y=����w�W�����<�u�;�ֺ��0��o� F��А����;4o�>���>j왾YV�=�Ծ����.>9z:<�ߒ�,7��<�P��K	>߂>���>���>��
�Y��=X��> ڴ>��� $?7J?!�?��̺kvh������J�\@�>�D?���=�_�u�����r�{��=�i?*�W?�eP����b?��]?�j�o=�k�þA�b���4�O?��
?��G���>��~?��q?���>1f�m9n����f>b���j��ݶ=�r�>!Y��d� ;�>��7?FM�>M�b>�-�=�w۾�w�;j��0?J�? �?���?�)*>��n�o3�c���$N��#�]?�L�>릾<�"?q0 �£Ͼ�>��ꎾc�᾽>���/��ݞ��=�����$�i����`ؽ�S�=�?�Fs?~Bq?۞_?�� �k�c�/Q^�i��)V�M���@�X�E�xE�pdC�(nn����*�������]H=��6�(l+�J�?3,?F�i�1� ?It����辡�0���V>�n"�:U��so>�O�<mX ��5Z>;�u�'5��}��b?xM�>��>�C?�SW��+����j-s����U�w��}�>y��>���>x	ͼ�<9��@��=ܑ�I*T�=9�� �>_<b?��G?+�m?#��r4�(]}��!���ȼῙ��B>]�=�h�>�"Q�n��zT ��7���p��o�s����n
��gR=�{,?�t�>�z�>���?�?H�
��~���Z�5�-�e�<��>�L^?���>O�>@E	��" ���>��l?5��>=�>�����[!���{���ʽt'�>��>���>N�o>J�,��"\��h��Q����9��c�=b�h?�����`��ޅ>�R?�ŉ:P�G<���>!�v�5�!�Y���'�f�>�{?���=��;>6}žL$��{�;��h�(?�?k���xI$�@&�>U�?g��>���>��?B-�>˾�����?�]?1J?��;?,)�>Y��<�i���ͽ�<'�~�R=F�>	S>w�o=�6�=��h�G��M���=pɨ=�bǼ��� w;˼cC0;6=�g6>1�׿-|H��Q���4������r蝾���AL*��Gn�ʝо){�������u�]T �M.�Ld��Q��i�|���?���?���Bಾ}?��7L��\-���>"� ��#\<f�䴙�b@[�*����y�i��6?�i<�5�N���'?{���h�ǿͯ���5ܾG" ?�B ?��y?w�o�"��8�� >~\�<�����뾉�����ο������^?G��>�
���/��>b��>ǝX>�Cq>���6鞾�\�<�?2�-?=��>�r�ڔɿ����Ա�<���?��@��8?��˾A�
��}��C1>u� ?��=e�=�� ��N�����=Zl�?�ʠ?�*��E�������1L?��g>1�f�R��=��->Ѽ�"�<(�8�a{�=��>�n:����=���Ǒ2>բ�>�qg��n�Ng�n�4>�K]>�a���=5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?:ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=u6�扤�{���&V�}��=[��>c�>,������O��I��V��=�x�,�ƿ���P�$;�=n�<�|'�� нqw��9���t;������L�b��� �=*,>&�z>H�>��6>�Y?piy?�]�>f!�=B�������g�j���(�8���ڽ�S���� �L��/��ٹ��Y�۾����MﶾX�N&s>\3���6%����8y�!?50`>_�@��x��Y��	�<�m��E�f���������������b��j�?�^?��x�����XP�d�.>�o?���<��3���JG>`*�>E��=�ȼ�|�mv�2G�{*]�k�6?�5?�`о��*����Q� �=C�M?xX�>O�>��=ۭb?��t�^�d�"d�=�Pm>���>c>	?��G�������,?Fy�?皽������>�7ƾ�|ƾ˖�><D>���܊V�:�>���>�������=�~z����mI?�A>��A��$��T:�� �=�>��a?Z%�>��L>�Z?~�:?*,]=�'�x�zf(�T�>�)V?�VU?�q3>IC�����r���xO?o�\?<n^>�0{�	�Ӿ�Z'�6��w?l�n?7K?->�M��o*��%�Ծ۔"?��v?3C^��j��l��7lW��>�O�>���>��9����>)d>?�"�jF�����G4���?ˊ@��?/4<�k�*�=�P?���>VVO���ƾo���F���%�n=�r�>Ch���`v�1��D,���8?̇�?O��>���������=O/�����?=��?t��s��<F0�ׁl�4�{w�<��=�$�����G}龁O7��������Ș�ތ��zʆ>��@�a��t�>��>����ޗͿ�����о�~�� ?{�>��Ͻ�ߦ�ͭh��0q��A�{CG���� Z�>�`>S�������D�z���:��7ڼ9��>x��3�>�(Y�����6���Bi<�|�>���>9�>6#��'���y6�?!=���nͿ X������X?i)�?ա�?��?�kj<�o�H�y������D?�-p?��X?�v!�76`�~+_�v�j?D��;T`���4��QE��U>43?�X�>��-�Q�|=��>��>�Y> #/�ߋĿ�϶�F������?$��?�d꾒��>o�?�+?Tf��=��m<���*�C��DA?�"2>�x��a�!�.=�ߧ���
?�{0?(n�'(�"�_?�a�r�p�l�-��ƽ�ڡ>��0��f\��I��1��Xe����G>y�)��?�]�?��?Y���#�6%?M�>f���M8Ǿ��<��>�)�>Q+N>{F_���u>e�7�:�Yg	>a��?,~�?-j?���-����U>��}?�O�>/�?�j�=X�?\��=⹾�!�=���=b29>/#�{�>�:?=�>�h_=�Խ+(�r(E�{Z������<�,��>`�e?�>?.�A>����˛��@%�o�W�c}��,ü��%��ؽ��#�6>��>׃>$Ч���3�?dg���ؿOk���~'��74?�ƃ>R�?=��X�t�K��)8_?w�>I�q/������#�z��?d:�?��?��׾��ͼ�>T�>�4�>R�Խ�͟�����_�7>[�B?m��1A����o�-��>���?��@	Ѯ?S�h�	?��\P��Aa~�4���6����=	�7?#.���z>~��>p�=�mv�+���H�s����>)A�?�y�?o��>��l?~o���B��1=!I�>r�k?u?_,n�]�¬B>m�?���*����O�f?��
@ou@V�^?�좿���X_�����#˾k��=y����/>����+ї<ы[=��b<+%
�8=���e>��=03�W�Ļ`ߧ=��1>��� 5'�'���������Y��P2�TQ"��XD�����KuJ���Ѿ���h�����k[�	R2������
��y>>��E?��G?��b?v�>�L�:?>�����=�m�=��C<h'�=�M?R{:?j�;?f�Z;u����S�-Lh����������g�>X�>Y׭>o�>Υ>�ʽ��*>j��=f�i>�˹��ad���=;�H�Zc>>}��>|�?U�>�C<>L�><ϴ�	2����h�Q
w�3̽6�?P���0�J��1��#9��W���th�=�a.?Z|>����>пd����2H?����_)�T�+�7�>7�0?�cW?E�>��� �T�r:>k��ݧj��_>1+ ��~l���)�Y%Q>�l?�*h>/Cv>u�2�o�6��aP�c߰�=�|>75?�K��K�5�6u�0ZH��`۾�tL>��>�M��d�[&���X~�X�i�&ez=��:?R ?be��uf����r�랾�&T>��Z>L�=�ݩ=+K>lNb��;ŽG�H�  )=���=M]>ޤ?O5n>�I>z��>����������>��=��=I?�_?��N��2��R�7��~P=wm�>��>V񞽺�{<��9��3��i��>D#J>T���T>�6�=�T�Je=0f���F����V~>��s���g<I޶<�+w�*����>�~?���#䈿��Rd���lD?]+?�=ɣF<��"�= ��hH��B�?j�@�l�?��	��V��?�@�?��G��=}�>�֫>�ξ/�L��?p�Ž+Ǣ�Ȕ	�I)#�^S�?��?��/�Qʋ�0l�t6>�^%?�Ӿ�=�>�?!��I��U���%Oh����=�p�>+A?���Y�z�X9���?s��>�d�X���vlſ;&g���>���?���?��a��$����C��(�>��?�4X?��}>�:�ur���>_*H?�\Q?*�>��"�x{$���?�2�?��?)I>V��?��s?5��>��x��d/������#7�=`�n;7Y�>#�>�����;F������d��$�j����{�a>�?$=��>���(���U�=���nJ����f���>\)q>5�I>�>� ?Pp�>�w�>�W=^������S���J�K?nV�?��BWl��<$��=�]��\?Co3?���"�Ͼ쟧>�M\?�G�?�%[?�P�>����2���v��Rߴ�?��<m�O>��>�8�>�	���K>��վ��@�8��>��>Pd��;�ھV9���}��H�>2� ?v5�>8r�=љ ?��#?�j>Q(�>1aE��9��9�E����>���>�H?��~?��?CԹ�~Z3�����桿w�[��;N>��x?V?^ʕ>a��������mE��@I�����a��?ltg?�S�0?12�?�??D�A?l)f>��ؾ]�����>j� ?����P�Jd�l����2?/�	?d�>з���Խ<U�<��#�義�?�PU?Ko?G��ug]�9U���(p<�ӣ�$�l=3�=l����>,k�=dg���>�F>)�*=�x�T�:�����>�=��>�%�=ia�g�/�d�-?���<���	�_=�lz��P�rt>�x>�fȾhl?%[�+~a��|��0���
+2�P��?��?���?3�3��^e�.�+?�u�?$?f� ?����J��}���ji����B���HYS=�w�>7��<鿾�栿ZB������)����ƽך�>���>�r?��>�*d>�	�>i=�� n޾����/
�?q������e����J�׾aX���0f�3��"b��j�>Ԟ����>v-?��>H�>j�>�dM��T>1*�=e�+>A\r>nD4>��>��=��+�0k[�o�F?��оVl��c�����<��g?uy?��?𻏼�,{�닦����>��?�׏?�zB>��r�Y�:�`??���>�J��O�>"S����=b��>>o��ڧ��^�=���>�ș>����GO��nG������I3?��D?� W�/����������n=M�?��(?�)���Q���o���W��S�M���=h�fj��i�$���p��돿{]��^$����(��f*=��*?5�?Q��������&k�?�0`f>0�><&�>�׾>&yI>��	�8�1�1^��I'�����_V�>�Y{?�S�>�;?��<?F:M?�k#?��>wG�>X�ѾFr�>}W1��D�>w;�>�
?��6?!;6?~�?r%?e�[>T������5�2��>3�?�+?�O?���>xڎ�l����_�S\�e���U붽�H=ս	= ��D��#�=DO>dD?x��gfK��~z�Sy ?�hb?ʑ#?��?&d?>C�'� �<9"S>֮ ?���>�A�����@L�V�&���[?���k��:!7?x3>�M����%�x�~=0��C����<�75�ش�>�o\>���=�!�!�o�) ;�L�l`�<�t�>k�?旊>�G�>�@��� �s���&�=��X>��R>�<>�*پ�y���&����g��y>{�?v�?�6g=��="��=X���N��d��F���i�<͞?�P#?IOT?މ�?@�=?,`#?@�>� �	F��[�������?�D-?�H�> ���Fоه��$�9�p?�?M]�f���,����������=��(�IPv�x�_5��H�/��<��`m�?�U�?DG���I<�I �W˘�߄þ2�I?���>���>��>+4"�.�U����t�M>���>-�@?ƫ�>LiN?�	v?�_?Z]�=�a;��L�������
PZ�b??G�n?�`?��v?&��>9�d>4��GR����n���W�1�!��������=_"r>Ƕ_>�<�>Ug�>v��=���;`�ͼ�텾��`=�=�>��>�J>|3�>^'|>~�߽l�F?�c�>�~���0�9Ŭ�&}z�OGN�0�t?~�?�A)?D?�<
O��@�ӌ����>P�?�g�?�(?�3_����=���d��i�Z�*��>9K�>���>f��=R`=r)>=�>vU�>Fy+�^���2���y�?Px??�,�=Hڿˠ�������벾b��<�1��Ӈ���=����=��\�2@��@�}����ȿ�l0��칗��e��'2��'s�>���=��%>�W�=xO=�T�=�c�;E_��8=���=�Ԅ��܃=�]]=��a��p)�c�=-`�=���;	����-˾�~}?�/I?R�+?�C?��x>�>�b6�K��>�4��F?�sU>��P�$r��/�:�����JR��h�ؾ�v׾d�妟�U�>��I��>;3>~��=iӄ<���=?�r=�l�=��]���=���=��=�۫=h�=o�>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?Ati��d�>M���㎽�q�=J����=2>s��=w�2�S��>��J>���K��A����4�?��@��??�ዿТϿ6a/>Sq9>E�>�7R��1��2^�f�_�Y��E!?�x:�O4ʾ̈́>
�=^�ܾ�;ȾH=H7>'5o=6;�\�&3�=jz���0=�wh=4��>��D>(��=z�����=<�G=�)�=DbS>��c�)�?�,�2�"6=�8�=��`>�'>�)�>&�(?�ZB?F=p?�0 >�%ܾy�!��#5���;�����?��.>;4<�d9>ԫ=?��B?=�u?���>���>��>���>@9�Y_A���Z�:�¾�߽�b?�?ހe>�H��-�[���,�E���!�/_?`�2?��=a�>]����	����{->��\%�ڲ>5�j<������:O�R�x��W��	~�>�i�>1�i>5�=&�=�U= ��>%E�=ʍ�˝�=�; =Ĝ,=r.K�o�>����{�=j>�:�2�f��o#��G�d��<���[���@=U��=���>��(>H��>��=ó���>?>Ϙ��6B��ڷ=����9>�{b��:s��B#��(��7>RhR>���o��
Z�>KM>��0>�_�?;�|?x�>����پHB��.�{�x?m��S�="�>M� ���5�Ryb��L�zžl!�>'۞>[�>�U>�12�סO����<�����?���?�I��� =�\�~d�Q���N��$�N��F�<��?�܅�{+�<���?�Q?�?�,�>*-9�Wy����@=r���H˹=��*��4���g=@A?9�?j�>����0��Fþx�"�>[KZ�#�D�?)��2�����E	��i)�>nh���վ,�1�8��A���bB��^�g�>a�G?\ʪ?��G�����~�X���P.���*?�Rd?#�i>�,�>!N
?��;	ؾ�����]����k?�1�?~>�?$��=�7�=�Z�����>B3?F��?�s�?�u?�7I����>cR�^(�=�.�b��=�	>���=IC�=���>�L??�O��q��G�����SY,���=�=~֠>�X�>eNH>Lي=��<Ь�=٦Y>�'�>�Gn>ӕ>-5�>kI�>\����	�)�'?���=ҏ�>��.?/"p> ��=Se�GmL=�L5��G�x�2�|%��D˽��%=�<7}E=�� ����>?ſ��?8EZ><���?�6���W�[�A>y�<>�½�'�>��I>{l>^)�>8^�>�� >�Ǌ>0F>TEӾ��>x��6o!��C�/zR�g�Ѿrz>臜���%�K��ov��aI��W���j���i�"(���*=�|.�<
J�?�,����k���)��W��-�??S�>*6?������>3��>{�>d,������-Í��S��?��?��c>�˞>�Y?�?^r6�[�/��.Z�=v��WC��3d�]��>��6W���w	��½�T`?�y?.A?��<wbz>(�?�g&�B�����>//��f:��+$=W��>���-KU�9�ξ�5ľ��D>��o?��?�?-�S�_3i��[(>��:?+�1?NUs?�1?�;?�`���$?�{5>�?�a
?��4?3/?!"?l/>��=zf\�q�$=g'��]P���ѽ��ʽѿ�]�7=I�y=�	:���;y=�Ҧ<j� �Uּ�;X���
�<619=7��=��=(��>;e?�  ?�L�>t�>s�����K������>�پ�����UE>�<��UҾ&o�>�A�?+I�?�C1?�/?F�5�_�@�d�=%m>���=�o>���>%�����F�<�~=��O=�0=$�>��%�n� �m�þ-�Ƽ�E>E�>"(z>zt���$>)���� ��̟;>�I9�Ͼ�����A�߅+��1y����>��K?IQ?���=���,��N�c��\?�A?x�H?�C~?HI	>�(־x	8���I�q�7��;�> 6м�=��R��k���07)�Af�<1`>uv�N��g>5��2㾐�k��BJ�r���v=���&F=A��Ӿ���OU�=���=O˼��"����׳���5J?�wh=�<���P��.���h>��>8��>�,Y�@f��>� 歾?4�=��>��:>Ԇü����F� |���>j�9?�k?[��?�ʆ���t��7��'
�Nc�yԘ>��W?s�2>�?t*>��>�1�W�����H�.{K���>5�?�Y
��x?��P��9b��X�#U�>�?���=f��>H�>?oL?Ԅ;?�?��>2M>9r�t��x�/?��?���=gM/���Լ2Zb�ީ|��V4?pm?d>}��>�V?ɲ�>�$?
c�?�H?6�8>�վ*<����>���>��B��u����7>AV?2�o>@%U?w��?��=�r�]�������ٽEL���!2?�&?��%?'�?���>�ݾ"1��V�=�b)?Q��?�j�?������=�c���@�>�c)>v�>p��>br�>,�4?筋?Uu?-[?ެs=���S#���\�����$��[�:W��="h��żM=y�<�^�=�+�=�!߼�l��ꢼ� ���[	�G��;&�>U�>��}��"�>���̯���ʆ>��;���Ⱦ�OT�:gZ���=��>�?Kʍ>����ծ=�C�>�4�>k@��>?�
?̝%?׌]��@i�����4t�衔>Q�a?.>�����+���(i��>�� �m?�Fc?^R�b�ݾM�b?��]?9h��=��þ~�b����b�O?;�
?9�G���>��~?j�q?N��>	�e�':n�*��Db�
�j�,Ѷ=`r�>LX�S�d��?�>l�7?�N�>-�b> %�=fu۾�w��q��j?��?�?���?+*>��n�W4�$w���G���^?ى�>�6���#?�� ���Ͼ�P��<+����%������R���}����$�H⃾=*׽/�=2�?�s?�Xq?��_?�� �r�c�C.^�����eV��+��"�W�E��$E��C���n��]�|.��y���G=�k>�qu3�?<�?��1?d�}��>?.YѾ�Ҿ�擾,F���- �j��=QR��Ӿ|׆<�TR>1)���F�PcԾQ>?I��>�o�>�s*?2�H��^�����/�_���V�>�Е>6�r>l�>k	>$�<߉�l츾����_��փ>��k?�`=??�k?�4���3��nd�:�+�,�*����c��>���>���>	Vǽ"���a"���,���c�����t�����S.�<>�L?�_�>�X
>�x�?�X?�7)�\�rk��Qc�O���l��>��A?�;�>i$�>J���|ݾ���>�+l?��>YF�>����Q���u�Ci����>�1�>
  ?�X>��+��xZ�ٍ�ϋ���5�k��=,f?]���&�d�l��>��S?&��<� =fe�>�!��(�������DO>��	?R��=��:>v\ɾ]��Q0{�`I��R@)?"�?x���yz*�'>�u"?`:�>=1�>��? �>	�¾�wf�W?E�^?��J?�_A?[��>,!=vF��^(ǽ��&�$�.=y!�>h�Z>Evl=E��=?!�ϔ\�3���?=�o�=	�ݼ����w<FG����;<���<�3>��ؿ�TO�P��H� �(߾aw�5N��"��q�o��,�ϩԾY����$o�b��s����t���/���x�&�G����?���?�_;mCϾ�⃿J�b�����޾>}9��l��~KT�/�׽���)�V˾��JB��^��HZ�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >UC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ďr�1�ɿc���}¤<���?0�@��@?��'����F�<=���>�C?��U>J�4�����O���I�>�J�?���?б+=�!U�݈��tl?pXW=G/9��*q�KJ�=���=PA=T����F>Lߎ>͒+�w�B���\9>C�>�XT�Б���n���;�n>�ޕ��@��3Մ?({\�f���/��T��:U>��T?�*�>-:�=��,?P7H�[}Ͽ�\��*a?�0�?��?$�(?,ۿ��ؚ>��ܾ��M?_D6?���>�d&��t�ȅ�=B6�Ɍ��s���&V�Q��=H��>5�>߂,�ߋ���O��I��u��=������n�W�*�P�9V�=�"ʼG���\v<iS�<M����龮F��4�؉<��A�=�v�>��S>m�Z>L�V?�t?�$B>&�|;F�K=�#b���Ҿ4�6>v�~�eÑ��{0�:�=�s��nR
�����������I���@ϾD�-��EE>�ꁿ;˧�䄾=�E�Iqp�,�C?��>K���Ƨk�b�>H��1���G3����=N!�r�L�>�R�?c�?��r?�+c�~4-�ѐ��;S[���)���J?j�\;�:���)��tI�<e�����=�.�>�>�H��yG�.t�Z�0?yq?6��*����(>���J�%=`E/?,?Q =M�>��?SE/�!�罧XU>��8>M��>���>I�>���������?H�V?�D��7y���S�>3fþ]����p_=�b>��.���?��_>��|<P��������7����m<!�V?䑉>T�'��~��d����ü�|=vss?��?>�>mi?[�C?
��<�	��\QR��'�v,�='g\?�k?�5>1�z�i*о㏡��5?O�_?	I>�\���⾟v,��� ��?�6p?UX?�����jy�����Z	�fm6?��v?yS^�F��L��MW�3��>��>	D�>�9�7#�>�m>?/"�$�������Q4����?<�@���?�O<B>�_��=?�?���>jO�� ƾ}!��ձ���"r=�d�>����v���;�,��)8?�r�?+/�>S���x����=#ݒ�礫?��?���-V�<c�ire���޾V��,=�=�t$<�0��a��b�&��{�� ��H���ō��a�>��@�f���Y�>�A��c�2`Ŀ;��&���D4�d�?�O�>��<E-q��bT�Ev�lJ?���;�A"��@C�>c�>IŔ�-���*�{�]m;����d�>����>��S��'��c����5<�>��>ݵ�>R)��3彾Cę?�[���?ο������t�X?0d�?�n�?.r?�:<��v��{{��^��%G?˂s?XZ?�I%� 9]���7��j?>`��T`���4�QGE��U>9#3?�@�>�-�B�|=>���>�l>&"/���Ŀ#ٶ��������?���?�m꾯��>���?s+?�i��6���[��-�*�J�0�};A?~2>2���Ը!�/=��Ғ�j�
?�~0?2x��-�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?'�>}�?{��=�m�>K��=c㰾I�,��J#>���=t�>�i�?+�M?%I�>W�=\9��/��YF�]DR�� �A�C���>�a? |L?KVb>6Ÿ��"2�+!���ͽ�1���cH@�D,���߽�4>3�=>�>o�D��Ӿ��?Pp�9�ؿj��p'��54?'��>�?��s�t�����;_?Lz�>�6��+���%���B�^��?�G�?A�?��׾�S̼�>B�>�I�>M�Խa���M�����7>.�B?B��D��u�o�k�>���?�@�ծ?gi��	?���P��Na~���^7����=��7?�0��z>���>�=�nv�ֻ��L�s����>�B�?�{�?0��>�l?t�o�M�B���1=,M�>��k?�s?eo�x�3�B>��?������L��f?��
@zu@p�^? ��ۿ���̾bܾ��K��M=�}>�ʴ�Yn�=D���߽�ӽ�>G��>۰�>�t!>NA(>u�.>d��>���|�%�릿��a�_�:D �C�׾�Z����xˊ�-$C���Ͼ����� &<_��=dX<�|�S��xýbN=���=��U?%'R?�r?���>Yy��Th+>u����<Z���%�=��>̖1?�L?��(??�=�@��	8d�H���Bx��l������>,PL>RW�>���>���><R��XN>�`O>Q�~>��=�Y$=�*��~l=��Q>���>g�>�[�>Ìl>e�>�ȿ�`���G
�^Ⱦd����ӯ?�SZ�ɖE�~��E�۽Y��_�=�j�>E�>=����Hֿ�<��L?b������i���N6�a��>J�k?.<�=fW9�ϔ�=�Zx>��V��0�� �>0�w�c���t��;�'<��X>�f>�ju>-�3��8�ɺP�����q?|>�K6?P*��%<9�F�u���H���ݾW�M>�8�>�VD�(��s	���'�Ji�VHz=s�:?>�?�������t��N��ȣQ>��\>�+=w�=-eM>`�.vƽ!1I���/=�w�=�]>bI�>�_>g�'>{5�>@f��,����>���=�o�L6S?]�D?��|qZ�BPP���9��χ>���>	"9>��=4�@�F�=q��>3�x>�hѽ
R㽐�!���D��ވ>	�>KO=�wM5��
�=��K�)�>���=�{߽8�_�ܘ=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿsg�>�y��Z�����q�u�d�#=ި�>�8H?�V��"�O��>��v
?�?�^�ĩ����ȿ�{v����>/�?���?�m��A��@���>��?2gY?�pi> g۾<_Z����>һ@?�R?u�>�9�ڎ'���?�޶?���?QP>���?j�r?���>-��q{*��ϲ��ً���|=ɂ�4�>.o>Pu��QF�{ǋ�A�|�� m�'s����=R�X=?��>�U��lǾd�=@X���h��Ԉ����>�bW>ga>�ף>�g?���>[	�>��E=�bc��)r��×�i�K?���?���A2n��U�<���=��^��&?�I4?&c[� �ϾL֨>�\?:?�[?�c�>���>���翿~��Ţ�<`�K>X4�>�H�>�%��JK>��Ծ!5D�6q�>�ϗ>���@ھF,��If��rB�>�e!?���>�ծ=ә ?��#?ޖj>�(�>9aE��9��[�E����>Ģ�>�H?�~?��?�Թ��Z3�����桿��[�4;N>��x?V?�ʕ>Y���烝�hE�CBI�w���V��?�tg?�S�+?>2�?��??A�A?f)f>���ؾ(�����>�!?���A�
7&����`�?��?��>�+����ս�м���H���?)T\?BS&?�<���`�:B¾���<kl'��9��<K�B���>})>�]����=��>GU�=J�m��8���W<��=Di�>���=�!8�1v���4/?�=*�e����=Z9d���D�"ǅ>^�>�剾�r?��!��R��SE���4����W�L�?^C�?��?"8�-T`���&?��?!'?�u�>�E����ľ���Z;=�t�P;��,>RC�>�;<.�Ҿ8X���m���C���m"��Q<{��>�)?��1?�?��>��>�{��B�2�A��������
�mUw�r]��,���x�<������/���� �[>�hὝ��>�;?�ʠ>���>,�>�99��NF=yΨ>-G��*	_;��}= G.>�X >c&@> W�>�8R?k�����'����N���QB?
�d?�~�>bj��n����8w? ��?_t�?�v>�:h���*�ρ?Hv�>���6N
?(9=���[��<kٶ�����p���i�5�>Ebս�:�"M��Kf���
?�?#����;��ٽ$T��@_�<o{�?M�*?a�,��1<�-p��;O�H}N�՛��Ь[�R��^�%�5ms�<�%���w膿�n*��*���� ?}?����m־ۤj��WP�r7��r�>��>_�f>G��>�b�>�>�w�?���L�������\�׷�>G��?F��>��I?�7<?��Q?RSL?xߌ>��>YT�����>A�u<��>?@�>�O8?��+?�#.?�?�c)?��\>_��z5��#�־O�?��?|�?x�?�?�È�s�̽ޘ�q�Q���{�,ف���n=�qP<>�ؽ��q��H=��Q>	� ?��?�T�"��ɾ��>A�9?,�?p�>����h������<B	?*�*?E��>��	��Xs����9?�ۇ? ��ٚ��W>]�K>��˽x19=�Sd<��)��Rýv�0��Y��$Ä��Q�=Z�>���gA����=�8ż��'�	 ?Fe?��>��>�����K��m��1�=�\>oBU>>>��ؾ�-�����jg�R�z>ѐ?���?"�z=/��=�'�=X�����ӧ�%����,�<�/?�/!?1�R?i��?l=?w�#?��>���В�=���1Ǣ���?�$?��>G^6�Vq�������b����>��?⠂����<�0��t
��_��j	�>��K����+��m��a��=j�Aj?�Q��?�W�?���<��m�Ͼ����3����9?z��>:b> �?�/�����!�b���>�,?b�>3��>=�i?�k?1�F?�v�=-�e���&������;�t<=8Q?��?1��?��:?��>p�>p���5[þ���/�ԼD�(�+ʏ����<j�>�M'>��>|P�>�ʟ<�;��+��RM�T�1<h/�>4R?%X(>���>���=�6N>.�J?��?����
��E;x�
������7g�?է�?p�[?؎�9>1��xY���lz�>V`�?�ˢ?��.?N�<�c�=;��@*��AT�f$/>G�>	�	?@�	>�V���`>(��>/��=��Y����K�yLŽA�>*�X?-hM>��Ŀ/�r��ƍ����)�<߽����s��Z���L���=���~��U���{j]�����˗�:�\����`p��Q?�l�=�Ƶ=���=��F=1<̼� �<M.�=�O=11�<�.v�.%5=N�X� ������UK =A:<~�=�����˾�}?�<I?Ԙ+?žC?��y>�=>�3�掖>ri���D?BV>cP�%�����;����[��#�ؾ+y׾��c�)Ɵ�GL>�dI��>o13>�6�=�9�<�/�=,Ls=$��=y�S��%=�)�=_�=*d�=���=M�>�X>�6w?X�������4Q��Z罦�:?�8�>[{�=��ƾp@?��>>�2������wb��-?���?�T�?>�?<ti��d�>M���㎽�q�=K����=2>y��=t�2�S��>��J>���K��N����4�?��@��??�ዿТϿ1a/>m�6>x�=��I���+�Ja�N�L�3�f��V?ϵ8�^ Ծ�	�>�^�=C�꾻�ؾ6a=pWC>B�'=�� ���[���=>�R��6=��f=><>h�=�[�� �=CDV=?��=�Oc>�k��V��u�:�=w)�=E�n>�Q$>�s�>8�?G�/?�@f?+��>�Ǚ���ھ�q��ű�>��5>�+�>S=�k&>���>˘B?=?�~D?U�>N_
=c��>n0�>"	/��w��QվD���lJ�?ݐ�?�X�>'�_�K�ʽ.Z��@����D�
?{(?��?�Ȯ>Z1�XC��X	�v� �9��ɱ7��E�=3�n�"�\�Q����1��p��T�>�u?�?x!Y>+ov>>��>.j�>o`�>ʢ>�I>M�1>��,=6^T�ȓ�p_=��<�[���x�N<`��;�5��7��2|<�zļG�L��v?�4h>�/?S|�>_?*JH>ws���^>g(M�8�>��$�>����{�9��A�%Oe����og�M��=Iq>�u���~�p/�>�J�>A�>N�?_�?ek�=+��u1!��]���0�{�B=�m5>`_���'�s}h�X�_�����>;_>�A�>��z>c�x����R�Ž�O��6�@��Y�>�$��ܮ_����W��3��.F���K����3�x�>8-{��H=���?�M?�Ԛ?G?<�*��x��7��>S����=������׊�9��>�%+?o��>�y~��׾u&Ѿa�Խ�>	�S��N��M��$c0���G��h��J��>¬��UҾ�1�-����S|C�\l����>�/N?�®?Q�[�����eR�ӑ���n�( ?�h?5��>^_?�N?!���P��R���E�=a�m?��?R��?^*>p
> �H��>Kg?ń�?:.�?��?�3���l�>��k��4]=&U�4>^=�}=E���p��K�>JS?��(?�{�&�(�x�#�p
�x㻾J�����:`�g>kZ�>^x�=���=�6���;>R�?b?n��>�X?�?�a�>D���h����'?�=�D�>�s2?<��>R�V=�F��E��<*�D�SM>��S.���ý�v佷ӳ<߭���E=����W�>��ƿ��?��S>�e��?���@*��U>9�R>�>ֽ2��>V'A>�x>+�>C��>��>ٴ�>��+>͗־3`>|���!�;�B��Q��1Ѿ��v>0����.%��v	�v���9�G����#��:j��J��{�;�r�<pI�?���|�m��!,�����?���>��5?�݋�Fs�jH>���>�D�>����F�������E޾5Ћ?���?�2c>��>	�W?%�?A�1�z�2��wZ�f�u�.A��e��`��΍�
���ν
��5����_?��x?=WA?�u�<v)z>��?��%��̏�J+�>�	/�i;�K�<=5�>#��*h`�tCӾ~�þ}�� @F>Z�o?�#�?BX?f V���l�X�&> �:?�1?�Nt?x2?��;?���$?�\3>�9? W?�.5?��.?��
?y$2>:��=|.����)=�R��f芾̢ѽ�ʽ2h� 3=xz=F^E9��<��=��<7L�b_ټ��	; ����-�<�d:=�¢=���=L=�>g�]?d�>�͆>��5?���h�4�I{���~1?֒�=	Q��q��oা4�򾎢�=��j?���?��Y?nbj>g|B���G�"�$>�Ə>�$'>��a>Ė�>����X���=�+>�`>*�=��B��R��m�
��i�����<[�>5�>��>��"�?BJ>`���6;n�Hbk>8�P��q���w'��
:�//��w�8�>.5G?Ʀ?�3j=i/�4Q���b�UZ(?0�;?��H?��~?8>8ھ5�G�]M�B�C�즢>��i=6b�x��������Q6��F��qqN>5Ԡ���u�t��>�������+g��a�Q�پ���>p��]⣽��tA���]뾶�<>�Y=˛��~�1���^�����L?L�q=7 �����<����=o��>��>@@��,>7 6�����f=�7?e/>��𽔜Ѿ�:H�>�	�*'�>�_J?�Hq?!��?K޵���a�=(M��1��(��-���2?�b�>L�2?F彬���?�J�6-꾋�V�,X����><�?�5���U�?���7�n���5n>�U?)�k=!�>G�^?w��>:(*?}�?��?�&�>�y;�]E��)00?���?̄=]U��N=V+�tY��T�>�V0?��W�`�c>�rI?��>�$?�fV?�w�>�+�=������ݷ�>���>�Fc�e��r\�>��w?��C>��2?"k�?X�>��\�dm�p�!�/�K>�|�=��?ИE?���>mB�>��)?����՛<8��>��*?�ل?��i?=�?�M�>4'�>T�1? Y=D�v>WN?�tr?��T?�jS?:�?$�)?e��<��8��=���=����vv�����]�=N�<����:*=�[��=���<���<>��=i������=�װ�@�.����>3nu>.���	/>�LþCx��_�@>Ĭ���Q�����u�:����=�z~>�?���>3"�V��=P��>��>n���'?i�?C�?BA:=�b�HپZ�G��ܰ>�jA?���=��l��Δ�wv�f�p=A n?'e^?X�T����M�b?�]?h��=���þζb���T�O?.�
?6�G���>��~?P�q?#��>d�e�:n�%���Cb�g�j��Ѷ=or�>pX���d��?�>��7?_N�>l�b>%'�=�u۾$�w�bq��0?s�?�?���?U+*>x�n�!4࿿������޹Z?�|�>����� ?����˾ڭ���������K����M����OĤ�޳������H۽6��=�?&�t?MWr?n�^?�m��d�)p^�L4��W�֮������E�QE�*TD���o�������o���%�@=�5j�}?�~�?�!#?��=�	L?6y�O�������.�=�����v=L���P� ��uý}�����{��ƾ��?K�>e��>@N/?-R`���F�6U��M��$
���=C?�B�>F�?v��=���=}��9�����`���n�M1u>�&`?��K?�}?Jp�mv/�I?p�X�)��I���Ő��qz>�,�=���>�1�����y$���3��k�m���V��C����=�:?�>]ԉ>� �?�-�>p��a����_�J-���=<��>��a?��>��s>��u@�b��>*�k?�~�>�ի>���!���v���޽`��>;L�>>�?�^h>17)���X�@������2q6����=��f?}�d�eg�>BT?r6H<m�;��>���T'�pU�!��A>=C?���=�V<> bž���+*}��ዾ=�6?�!?�M���m0����>.@?���>�k>�)�?�X�>k �"��=��>�W?5W)?�]?�g�>-#=Ʃ>'$}���[��K�t�{>!�`>Ό�>�Y>������hq�y�Q>s�q=2�R�V���!���_=!	��J�_>l0>��ӿaA��$۾�3��Uƾ������v���"Z���t�7�þ��i��gy�ŷA�8:��)g�T��W��BkZ���?�)�?�`��'��.���炿��	�j��>?栾(����Ӈ�Fڿ�#˾<Ѿ
Ⱦ�*��iB���d������'?����c�ǿW����:ܾ� ?iV ?�y? ��}"�f�8�<. >���<�ɚ��<�����ο'y��/�^?��>W
�*[����>�Ƃ>��X>5$q>Z��m)�����<?�-?���>�3r���ɿۊ�����<���?�@�A?�(�����IT=h��>í	?y+?>N]1����?����>�3�?/�?�M=P�W��	�-ge?5 <��F���ݻ{��=���=K�=��e�J>���>����&A�@Kݽ��4>���>~3%��sR^�i��<�G]>��Խ�Ĕ��ӄ?�s\�f���/��R��;_>`�T?��>+g�=\�,?�3H��{Ͽ\�\��*a?�/�?��?��(?ȿ�E�>��ܾ2M?�:6?��>V&���t��o�=e��r���Ⱥ�JV��F�=w��>��>��,�ɔ�̑O��9����=m�|ٻ�y�:�2l&�zXL>��t�þ��fZ���L=@�z����O��$꨼���<6\�=
\�>s��=�E7>ao�>.R?��q?�Ʒ>nE>�xý����X�߾�|K="�w��Q|�Wv�8Ϫ�&�������p��p$���5�w��������6�
��;Y�]�ܚ��ný�Гf���S�:5K?�R>)�־eW0�3��>+�۾%ϑ���_���=<y���4�~\���?�?F?+Vx�b�D�c1��f���N=��t?�, �����q�?"1>m�����_>�͒>��<t}Ǿ�N������C?g�,?{Y��Yh��{L�>�=�Y�=�tV?N68?�1e�dV�>-�?��þ��u��_>�M�>`�>1�>Ev�>�k��Ś��8-?�0U?�ꀾ��־6��>�L���0��kN�>S�V>2��Q�=��>�~8���ýZ�>NT>��d�*W?ܱ�> �)��
��0������<=��x?��?�9�>eNk?��B?<�<�0����S�����w=��W?�1i?��>"Ɂ�hоo��W�5?��e? �N>�h����.�*B�?��n?b?�Ρ�zh}�������[6?�v?�o^��r�������V�?�>�\�>���>+�9�th�>k�>?�#�4H������)W4�$Þ?�@���?�m<< ���=�<?R^�>ٲO�WBƾ~{�������q=9(�>T���fv����O,�؅8?���?���>�������G��=�P���,�?��z?09�i�=�5�b����L.��YU>&���� >�$�|
&���㾴�D�-;��;n�~y}>��@j��t�>�����ڿ��ȿ$u~���-��J:&?�a�>,�=�	��N�4�/=���"��@T��þD>�>6>Hʕ��8��F�{�ǐ;�Y�����>-	����>�VS�Xõ�>$��{�:<���>ר�>{��>=����D��0Ù?h���.ο���o��M�X?[n�?	k�?T6?�G<{�v��T|���JG? fs?5�Y?��$�v�]��2:�%�j?�_��xU`���4�uHE��U>�"3?�B�>S�-�_�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�TҒ�¼
?V~0?{�f.��_?q�\�0�n�>�-��ڽ���>#\��gi��jR�?/��zb�Q����N�?���? �?�$2�H�E�+?_�>=V���)Ǿ8HM=�b�>@��>��D>1�ϽmGD>����+�GZ#>a��?�J�?�6?�䐿Ġ��Cm6>�j{?㕶>/��?_:�=�E�>w�= ű��%���Q>!��=��#���?�L?�_�>1�=�M7��/�mE�QsR���C�B�d^�>�da?�\L?�Mf>1ݿ�c�!�	� ���e�)����_�?����Wѽ�L7>W�<>�>�K�12վ��?8p�1�ؿ�i���o'��54?(��>�?�����t�7���;_?4z�>�6��+���%���B�Y��?�G�?7�?��׾�R̼�>�>�I�>��Խ����Q�����7>3�B?[��D����o���>���?�@�ծ?Ui��	?o��P��Ia~����( 7� ��=�7?�/��z>���>Y�=ov�̻�� �s�깶>�B�?{{�?g��>�l?u�o��B�%�1=�L�>K�k?�s?��n�_󾧲B>��?!�����JL��f?��
@lu@f�^?��ߏӿE����l��+Ѿ�g�=U��=6��>K(�Ѭ���<��;<���Zr=��^>r��=�	8=�h�>�*w>�'G>�x����#��λ�����:�4���qk��\D��E���y���?�h׾���k�d�313��|��҃�&౼-�V=�#�=N�O?˝Z?��?~�?P�,��>�i���?�&�<�I>TE><4?�V?��?o�0�;N��Bi��q�������V�4	�>0v+>�E�>%��>Mٱ>4�=)?)>7�R>7�9>�$�=<+�;�����<ւH>L˶>���>Zww>_.>J>�]���#����`��n��Sɽ�ͤ?� ��;�G��d����x�OG��g"�=,+?�!>%�����οC�����E?H������! ����= �+?Z?>�ΰ�s�]�B>i�'���k���	>���qn�4�%��@>!?�x>�n�>8�3��>2�"h�A����>CC<?kپ�(���p�KM�q���7�>Oۖ>#�����#������Nf�6��<��??-�?�^�l���M�F�d9۾=�R>Y�>i�Ž�5L��o>�&��g/��*��Z[��5�s=~/e>A?��1>N��=$�>_���'I�L��>��>>��3>5�@?dz$?�)�}���$��#�,�F~>D��>l)�>@>�zL���=	�>~e>V�ټ˹x����pVM���P>;�Q���Z� *~�my�=!T�����=۹w=�����>���
=��~?�{��f∿�뾍s��kD?�1?Vː=��G<Ay"�����T�����?3�@sn�?Ry	���V���?�B�?+������=os�>�߫>GξU{L�m�?�Vƽ�آ�ڍ	��"�S�?��?ܖ/��ȋ��l��.>�f%?��ӾMh�>}x��Z�������u���#=Q��>�8H?�V����O�{>��v
?�?�^�੤���ȿ1|v����>T�?���?j�m��A���@����>=��?�gY?oi>�g۾7`Z����>̻@?�R?��>�9���'���? ߶?֯�?x)H>���?��v?c�>�Sӽ�-��a��6��c	=l�D���>#�>�����#O��f�����O�`�C6���>F3=���>K���������=�6���L��:Xo�\�>Cn>Ӹ3>���>��>A4�>�/�>��~=a(��U��눁���K?���?E��h2n�C��<%��=V�^�%?EK4?E�[�8�Ͼب>��\?���?z[?�b�>���$=���忿�|����<S�K>W3�>�D�>\���QK>4�Ծ;2D��j�>�ї>N��+Eھ}/�������C�>7c!?0��>�ۮ=\+ ?}(?;9>�Y�>*`1�\����-@��R�>@�>\?��{?�F?�c����+� -������BZ�p�E>>Nm?�� ?eˣ>�����0�����<""B��b0��~�?�
o?>=�`��>e$�?�1?ne-?r1�>z���H�fp�����>O�!?�\�e�A�9&������?��?��>�9��
Rѽ�fڼ����}��<?�y\?
B&?��)�_�����[
�<�F;�H_{��y+<a�!��E> �>P������=��>Ev�=�8i��#6��kl<:m�=C
�>��=4�0�H����=,?{�G�ڃ��=D�r��vD���>�LL>����q�^?�j=�{�{�#��?x��1	U��?���?�j�?�����h��#=?B�?�	?�!�>�J���}޾J�ྒQw�mvx�~v���>e��>0dl��ԏ��-���eF��� ƽ	W0�~��>��	?q@�>��>�/�>���>��B�����v����<�n���ɾ.��(r���v��\\��)߽�ͽ?�⽶��������]�>�c��(��>�W?��>(�>�2�>�����>M�j=P�>-��=ɇ�=�`�>���<T�>}!�;�R?�����'�2��򃧾��D?�
a?$��>�"��h��#�D�?�Ԑ?&a�?P�q>��e���)��3?V  ?�~�xh?O')=�����(<��������>�L��e{�>�����d8��Q���w��A?��?�ƪ�&Fľ�pǽ�䟾�r=)��?��(?�*��BQ��cp���W�:S��&���c�2���w#���p�鷏����D�� ;(�a�=Z*?�W�?r��mK��\Yk��>�`�d> =�>�)�>{Ͼ>i�L>�	���1��/^�1�%�6���?�>6\z?�g�>9K?�6?ŧ_?Y3?>>��>Ҿ0i?JiP=���>�*�>o�?p�?�	?��>��&?��X>h��u��נ����?	KN?Q�?���>1?����Ũ�= �>���=�l���ڙ�w^P>ؼU<�:���'��Hs4��E]>}�?Q���r8�����)m>G�7?�R�>.U�>�M���R��!�<��>��
?	�>]b��t�q�����>B��?����A�<��(>��={���J:��=ht��Ī�=8~��xL1��d!<�O�=�={����E�:ȉ[:�U�;jƬ<u�>;�?ȓ�>�C�>m@��� �=���f�=�Y>uS>�>�Eپ�}���$��V�g�^y>�w�?�z�?�f=v�=���=�|��BU�����:������<��?J#?,XT?M��?K�=?tj#?�>+�VM���^�������?�?�|�>\��}����ÿdbX���?�>�#b��h;o�N�{ ��׶�	��>��-�����C����|�������hW��t�?O=�?����� ����޾Jᓿ�eH�: ,?QP�=��>�*�>v\6���T���9��;�=|'�>p U?�P�>u"e?�Ar?�[:?��>��8��[���|���� =d,R�ɩ>?\Ax?���?��2?o��>>+K>[_��1�`	�Z�
��OɽG{��Ն^=��|>�ac>��>�ۧ>��u>��E�⽥V�X����Ш>�E?�~�=���>���>�U>�H?���>��>T��m���8k�e���Cv?���?G�#?�r=i����H������>��?�Z�?��)?k�9��/�=&h�h���;�c����>���>Bɞ>��=��1=/!>��>p��>�G&�g�� 3���IX?�"G?���=]Nƿ�g��g��f�۾<>�j��H���P=�Z�����=`S޾1�s]��_��i�b�5�o��Dؾ������4��;�>G�=�!>�l]=)"h=����.=o��F,=`d�v=#���e�s˼��b���=��\����=E��=~b˾��}?�EI?,�+?�C?�y>̫><�6��
�>����S?�U>��N��#��04;�漨�D	�� �ؾ�{׾@�c�����ZK>�I�G�>��2>Ĵ�=Ʀ�<G��=�s=�F�=��\���=x9�=�c�=��=~a�=��>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>?)4>ê >TS���1��FX�Db�4�Y�>�!?5�9�[z˾ǡ�>T�=�O޾Y{ž �7=��8>V�O=�����[�t3�=��x��uA=y�l='ԉ>��C>Y��=t����=�\2=�=��L>Dn��`�;�Nj,��7=C
�=S'b>��&>(��>��?��4?x9}?��>:����{��\����c.>��8>��>��<��A>S
�>��&?�*?�_H?Z��>�C�<��>�=�>I6,�i�r�jپ����'#����?��?2�>��;�ֽ���G�M���#?p?V�?�y�>F�	���޿�H��<L��g��!��S�=�T�!>U��t��Xj��gd��y�>_�><��>A��> 9t>Q��>��>�v�>e>�K�=f?>oTc�FP˻*gI�� 8=;E�=�	�=-��=jF�=M��=�������<mc\>��̨ѽ��P�.��=��>�e>���>�o�=�����_/>k�����L���=�;��.B�!-d��@~��/�t�6���B>;!X>����h/����?��Y>�?>t��?�;u?� >M�W�վ�C��0(e�QkS��=��>z�<�Hs;��M`�M�M��sҾ�Y�>Y3u>l��>�l>�D�v�,�_mJ=�:Ѿ �6�=��>B�ܾcf	��
��l4b����n��M�\�����9%?Q���(Us��&?U�>? ��?5%!?Շ9;!���J>Z=w�D]=Ց��	5�7���t��>��?�c&?c�e�E��O�˾*ý>͹>KF���O��t��N/��������:̱>�ͮ�{Ӿj�3�����^��ʽD�
)l�Y��>ΧM?:��?��g�yi���FN�3Y� Z�,q?�h?��>8�?�?>a���뾲���P��=n�m?���?���?ɻ>���=�Gv��{�>��>.ޕ?�9�?0�l?Fv5��s�>6����W>t�d��=�4>�=���=�,?��?�?-*��~$�U��>�d�d�Ф�<�x�=7�>�)�>9�Q>B[>M	�=_+c<��>�ĥ>�g�>��l>徵>�%�>G$�������&?G �=9��>P�2?R0�>mf]=΀��3E�<��N�X�A��9,������彺}�<Ќ���T=��ɼ[�>�>ǿ$�?SuT>�Q��?jq���6�+FR>��R>0�׽���>��F>�U}>6Ů>�d�>_O>�>�?'>�<Ҿ��>Ҟ��� ��D��WR�LѾJkx>3b��� $�E
�m���� N��V��]���j��L���E>��!�<�K�?[��Ti�H�(�*Y�Nc
?N�>d�5?��������
�>ym�>�ލ>|)��t��������8ݾL@�?[��?�;c>��>p�W?"�?�1�"3�'vZ�!�u�x(A�>e��`�i፿Ӝ��:�
������_?��x?�xA?H�<�9z>]��?��%�Pӏ��)�>�/��&;�F?<=d+�>*����`�ٮӾ0�þ�8��GF>��o?Q%�?Y?TV���l�7Q'>�:? �1?�At?��1?�;?fY�&�$?�24>+_?�N?&M5?l�.?w�
??�1>4�=�ĵ��#'=����̊�?eѽrʽ�J��1=BV{=�؞9i<��=P£<֎��ۼ��;뺡��m�<[>;=�+�=�Z�=�ͷ>��^?i��>`9~>#:9?��нe�3�
"���r9?��=/����Ń�����Q���=�
d?���?X�M?9Ё>X�I�#f@�<3>+�>$&8>�ق>���>��3��>��J�=���=���=��=5�����a�����٩�<V��=?�>�w><��9D>b夾;o�6@z>ʤ[��o��nGB�!AF�R4�u�z����>/oO?*??
�k=��9:��a�Ț$?��7?].N? �?�m�=��پ4�>���N�]����>z>#=���M���#栿~�=����r��>&��N��g>5��2㾐�k��BJ�r���v=���&F=A��Ӿ���OU�=���=O˼��"����׳���5J?�wh=�<���P��.���h>��>8��>�,Y�@f��>� 歾?4�=��>��:>Ԇü����F� |���>j�9?�k?[��?�ʆ���t��7��'
�Nc�yԘ>��W?s�2>�?t*>��>�1�W�����H�.{K���>5�?�Y
��x?��P��9b��X�#U�>�?���=f��>H�>?oL?Ԅ;?�?��>2M>9r�t��x�/?��?���=gM/���Լ2Zb�ީ|��V4?pm?d>}��>�V?ɲ�>�$?
c�?�H?6�8>�վ*<����>���>��B��u����7>AV?2�o>@%U?w��?��=�r�]�������ٽEL���!2?�&?��%?'�?���>�ݾ"1��V�=�b)?Q��?�j�?������=�c���@�>�c)>v�>p��>br�>,�4?筋?Uu?-[?ެs=���S#���\�����$��[�:W��="h��żM=y�<�^�=�+�=�!߼�l��ꢼ� ���[	�G��;&�>U�>��}��"�>���̯���ʆ>��;���Ⱦ�OT�:gZ���=��>�?Kʍ>����ծ=�C�>�4�>k@��>?�
?̝%?׌]��@i�����4t�衔>Q�a?.>�����+���(i��>�� �m?�Fc?^R�b�ݾM�b?��]?9h��=��þ~�b����b�O?;�
?9�G���>��~?j�q?N��>	�e�':n�*��Db�
�j�,Ѷ=`r�>LX�S�d��?�>l�7?�N�>-�b> %�=fu۾�w��q��j?��?�?���?+*>��n�W4�$w���G���^?ى�>�6���#?�� ���Ͼ�P��<+����%������R���}����$�H⃾=*׽/�=2�?�s?�Xq?��_?�� �r�c�C.^�����eV��+��"�W�E��$E��C���n��]�|.��y���G=�k>�qu3�?<�?��1?d�}��>?.YѾ�Ҿ�擾,F���- �j��=QR��Ӿ|׆<�TR>1)���F�PcԾQ>?I��>�o�>�s*?2�H��^�����/�_���V�>�Е>6�r>l�>k	>$�<߉�l츾����_��փ>��k?�`=??�k?�4���3��nd�:�+�,�*����c��>���>���>	Vǽ"���a"���,���c�����t�����S.�<>�L?�_�>�X
>�x�?�X?�7)�\�rk��Qc�O���l��>��A?�;�>i$�>J���|ݾ���>�+l?��>YF�>����Q���u�Ci����>�1�>
  ?�X>��+��xZ�ٍ�ϋ���5�k��=,f?]���&�d�l��>��S?&��<� =fe�>�!��(�������DO>��	?R��=��:>v\ɾ]��Q0{�`I��R@)?"�?x���yz*�'>�u"?`:�>=1�>��? �>	�¾�wf�W?E�^?��J?�_A?[��>,!=vF��^(ǽ��&�$�.=y!�>h�Z>Evl=E��=?!�ϔ\�3���?=�o�=	�ݼ����w<FG����;<���<�3>��ؿ�TO�P��H� �(߾aw�5N��"��q�o��,�ϩԾY����$o�b��s����t���/���x�&�G����?���?�_;mCϾ�⃿J�b�����޾>}9��l��~KT�/�׽���)�V˾��JB��^��HZ�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >UC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ďr�1�ɿc���}¤<���?0�@��@?��'����F�<=���>�C?��U>J�4�����O���I�>�J�?���?б+=�!U�݈��tl?pXW=G/9��*q�KJ�=���=PA=T����F>Lߎ>͒+�w�B���\9>C�>�XT�Б���n���;�n>�ޕ��@��3Մ?({\�f���/��T��:U>��T?�*�>-:�=��,?P7H�[}Ͽ�\��*a?�0�?��?$�(?,ۿ��ؚ>��ܾ��M?_D6?���>�d&��t�ȅ�=B6�Ɍ��s���&V�Q��=H��>5�>߂,�ߋ���O��I��u��=������n�W�*�P�9V�=�"ʼG���\v<iS�<M����龮F��4�؉<��A�=�v�>��S>m�Z>L�V?�t?�$B>&�|;F�K=�#b���Ҿ4�6>v�~�eÑ��{0�:�=�s��nR
�����������I���@ϾD�-��EE>�ꁿ;˧�䄾=�E�Iqp�,�C?��>K���Ƨk�b�>H��1���G3����=N!�r�L�>�R�?c�?��r?�+c�~4-�ѐ��;S[���)���J?j�\;�:���)��tI�<e�����=�.�>�>�H��yG�.t�Z�0?yq?6��*����(>���J�%=`E/?,?Q =M�>��?SE/�!�罧XU>��8>M��>���>I�>���������?H�V?�D��7y���S�>3fþ]����p_=�b>��.���?��_>��|<P��������7����m<!�V?䑉>T�'��~��d����ü�|=vss?��?>�>mi?[�C?
��<�	��\QR��'�v,�='g\?�k?�5>1�z�i*о㏡��5?O�_?	I>�\���⾟v,��� ��?�6p?UX?�����jy�����Z	�fm6?��v?yS^�F��L��MW�3��>��>	D�>�9�7#�>�m>?/"�$�������Q4����?<�@���?�O<B>�_��=?�?���>jO�� ƾ}!��ձ���"r=�d�>����v���;�,��)8?�r�?+/�>S���x����=#ݒ�礫?��?���-V�<c�ire���޾V��,=�=�t$<�0��a��b�&��{�� ��H���ō��a�>��@�f���Y�>�A��c�2`Ŀ;��&���D4�d�?�O�>��<E-q��bT�Ev�lJ?���;�A"��@C�>c�>IŔ�-���*�{�]m;����d�>����>��S��'��c����5<�>��>ݵ�>R)��3彾Cę?�[���?ο������t�X?0d�?�n�?.r?�:<��v��{{��^��%G?˂s?XZ?�I%� 9]���7��j?>`��T`���4�QGE��U>9#3?�@�>�-�B�|=>���>�l>&"/���Ŀ#ٶ��������?���?�m꾯��>���?s+?�i��6���[��-�*�J�0�};A?~2>2���Ը!�/=��Ғ�j�
?�~0?2x��-�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?'�>}�?{��=�m�>K��=c㰾I�,��J#>���=t�>�i�?+�M?%I�>W�=\9��/��YF�]DR�� �A�C���>�a? |L?KVb>6Ÿ��"2�+!���ͽ�1���cH@�D,���߽�4>3�=>�>o�D��Ӿ��?Pp�9�ؿj��p'��54?'��>�?��s�t�����;_?Lz�>�6��+���%���B�^��?�G�?A�?��׾�S̼�>B�>�I�>M�Խa���M�����7>.�B?B��D��u�o�k�>���?�@�ծ?gi��	?���P��Na~���^7����=��7?�0��z>���>�=�nv�ֻ��L�s����>�B�?�{�?0��>�l?t�o�M�B���1=,M�>��k?�s?eo�x�3�B>��?������L��f?��
@zu@p�^? ��ۿ���̾bܾ��K��M=�}>�ʴ�Yn�=D���߽�ӽ�>G��>۰�>�t!>NA(>u�.>d��>���|�%�릿��a�_�:D �C�׾�Z����xˊ�-$C���Ͼ����� &<_��=dX<�|�S��xýbN=���=��U?%'R?�r?���>Yy��Th+>u����<Z���%�=��>̖1?�L?��(??�=�@��	8d�H���Bx��l������>,PL>RW�>���>���><R��XN>�`O>Q�~>��=�Y$=�*��~l=��Q>���>g�>�[�>Ìl>e�>�ȿ�`���G
�^Ⱦd����ӯ?�SZ�ɖE�~��E�۽Y��_�=�j�>E�>=����Hֿ�<��L?b������i���N6�a��>J�k?.<�=fW9�ϔ�=�Zx>��V��0�� �>0�w�c���t��;�'<��X>�f>�ju>-�3��8�ɺP�����q?|>�K6?P*��%<9�F�u���H���ݾW�M>�8�>�VD�(��s	���'�Ji�VHz=s�:?>�?�������t��N��ȣQ>��\>�+=w�=-eM>`�.vƽ!1I���/=�w�=�]>bI�>�_>g�'>{5�>@f��,����>���=�o�L6S?]�D?��|qZ�BPP���9��χ>���>	"9>��=4�@�F�=q��>3�x>�hѽ
R㽐�!���D��ވ>	�>KO=�wM5��
�=��K�)�>���=�{߽8�_�ܘ=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿsg�>�y��Z�����q�u�d�#=ި�>�8H?�V��"�O��>��v
?�?�^�ĩ����ȿ�{v����>/�?���?�m��A��@���>��?2gY?�pi> g۾<_Z����>һ@?�R?u�>�9�ڎ'���?�޶?���?QP>���?j�r?���>-��q{*��ϲ��ً���|=ɂ�4�>.o>Pu��QF�{ǋ�A�|�� m�'s����=R�X=?��>�U��lǾd�=@X���h��Ԉ����>�bW>ga>�ף>�g?���>[	�>��E=�bc��)r��×�i�K?���?���A2n��U�<���=��^��&?�I4?&c[� �ϾL֨>�\?:?�[?�c�>���>���翿~��Ţ�<`�K>X4�>�H�>�%��JK>��Ծ!5D�6q�>�ϗ>���@ھF,��If��rB�>�e!?���>�ծ=ә ?��#?ޖj>�(�>9aE��9��[�E����>Ģ�>�H?�~?��?�Թ��Z3�����桿��[�4;N>��x?V?�ʕ>Y���烝�hE�CBI�w���V��?�tg?�S�+?>2�?��??A�A?f)f>���ؾ(�����>�!?���A�
7&����`�?��?��>�+����ս�м���H���?)T\?BS&?�<���`�:B¾���<kl'��9��<K�B���>})>�]����=��>GU�=J�m��8���W<��=Di�>���=�!8�1v���4/?�=*�e����=Z9d���D�"ǅ>^�>�剾�r?��!��R��SE���4����W�L�?^C�?��?"8�-T`���&?��?!'?�u�>�E����ľ���Z;=�t�P;��,>RC�>�;<.�Ҿ8X���m���C���m"��Q<{��>�)?��1?�?��>��>�{��B�2�A��������
�mUw�r]��,���x�<������/���� �[>�hὝ��>�;?�ʠ>���>,�>�99��NF=yΨ>-G��*	_;��}= G.>�X >c&@> W�>�8R?k�����'����N���QB?
�d?�~�>bj��n����8w? ��?_t�?�v>�:h���*�ρ?Hv�>���6N
?(9=���[��<kٶ�����p���i�5�>Ebս�:�"M��Kf���
?�?#����;��ٽ$T��@_�<o{�?M�*?a�,��1<�-p��;O�H}N�՛��Ь[�R��^�%�5ms�<�%���w膿�n*��*���� ?}?����m־ۤj��WP�r7��r�>��>_�f>G��>�b�>�>�w�?���L�������\�׷�>G��?F��>��I?�7<?��Q?RSL?xߌ>��>YT�����>A�u<��>?@�>�O8?��+?�#.?�?�c)?��\>_��z5��#�־O�?��?|�?x�?�?�È�s�̽ޘ�q�Q���{�,ف���n=�qP<>�ؽ��q��H=��Q>	� ?��?�T�"��ɾ��>A�9?,�?p�>����h������<B	?*�*?E��>��	��Xs����9?�ۇ? ��ٚ��W>]�K>��˽x19=�Sd<��)��Rýv�0��Y��$Ä��Q�=Z�>���gA����=�8ż��'�	 ?Fe?��>��>�����K��m��1�=�\>oBU>>>��ؾ�-�����jg�R�z>ѐ?���?"�z=/��=�'�=X�����ӧ�%����,�<�/?�/!?1�R?i��?l=?w�#?��>���В�=���1Ǣ���?�$?��>G^6�Vq�������b����>��?⠂����<�0��t
��_��j	�>��K����+��m��a��=j�Aj?�Q��?�W�?���<��m�Ͼ����3����9?z��>:b> �?�/�����!�b���>�,?b�>3��>=�i?�k?1�F?�v�=-�e���&������;�t<=8Q?��?1��?��:?��>p�>p���5[þ���/�ԼD�(�+ʏ����<j�>�M'>��>|P�>�ʟ<�;��+��RM�T�1<h/�>4R?%X(>���>���=�6N>.�J?��?����
��E;x�
������7g�?է�?p�[?؎�9>1��xY���lz�>V`�?�ˢ?��.?N�<�c�=;��@*��AT�f$/>G�>	�	?@�	>�V���`>(��>/��=��Y����K�yLŽA�>*�X?-hM>��Ŀ/�r��ƍ����)�<߽����s��Z���L���=���~��U���{j]�����˗�:�\����`p��Q?�l�=�Ƶ=���=��F=1<̼� �<M.�=�O=11�<�.v�.%5=N�X� ������UK =A:<~�=�����˾�}?�<I?Ԙ+?žC?��y>�=>�3�掖>ri���D?BV>cP�%�����;����[��#�ؾ+y׾��c�)Ɵ�GL>�dI��>o13>�6�=�9�<�/�=,Ls=$��=y�S��%=�)�=_�=*d�=���=M�>�X>�6w?X�������4Q��Z罦�:?�8�>[{�=��ƾp@?��>>�2������wb��-?���?�T�?>�?<ti��d�>M���㎽�q�=K����=2>y��=t�2�S��>��J>���K��N����4�?��@��??�ዿТϿ1a/>m�6>x�=��I���+�Ja�N�L�3�f��V?ϵ8�^ Ծ�	�>�^�=C�꾻�ؾ6a=pWC>B�'=�� ���[���=>�R��6=��f=><>h�=�[�� �=CDV=?��=�Oc>�k��V��u�:�=w)�=E�n>�Q$>�s�>8�?G�/?�@f?+��>�Ǚ���ھ�q��ű�>��5>�+�>S=�k&>���>˘B?=?�~D?U�>N_
=c��>n0�>"	/��w��QվD���lJ�?ݐ�?�X�>'�_�K�ʽ.Z��@����D�
?{(?��?�Ȯ>Z1�XC��X	�v� �9��ɱ7��E�=3�n�"�\�Q����1��p��T�>�u?�?x!Y>+ov>>��>.j�>o`�>ʢ>�I>M�1>��,=6^T�ȓ�p_=��<�[���x�N<`��;�5��7��2|<�zļG�L��v?�4h>�/?S|�>_?*JH>ws���^>g(M�8�>��$�>����{�9��A�%Oe����og�M��=Iq>�u���~�p/�>�J�>A�>N�?_�?ek�=+��u1!��]���0�{�B=�m5>`_���'�s}h�X�_�����>;_>�A�>��z>c�x����R�Ž�O��6�@��Y�>�$��ܮ_����W��3��.F���K����3�x�>8-{��H=���?�M?�Ԛ?G?<�*��x��7��>S����=������׊�9��>�%+?o��>�y~��׾u&Ѿa�Խ�>	�S��N��M��$c0���G��h��J��>¬��UҾ�1�-����S|C�\l����>�/N?�®?Q�[�����eR�ӑ���n�( ?�h?5��>^_?�N?!���P��R���E�=a�m?��?R��?^*>p
> �H��>Kg?ń�?:.�?��?�3���l�>��k��4]=&U�4>^=�}=E���p��K�>JS?��(?�{�&�(�x�#�p
�x㻾J�����:`�g>kZ�>^x�=���=�6���;>R�?b?n��>�X?�?�a�>D���h����'?�=�D�>�s2?<��>R�V=�F��E��<*�D�SM>��S.���ý�v佷ӳ<߭���E=����W�>��ƿ��?��S>�e��?���@*��U>9�R>�>ֽ2��>V'A>�x>+�>C��>��>ٴ�>��+>͗־3`>|���!�;�B��Q��1Ѿ��v>0����.%��v	�v���9�G����#��:j��J��{�;�r�<pI�?���|�m��!,�����?���>��5?�݋�Fs�jH>���>�D�>����F�������E޾5Ћ?���?�2c>��>	�W?%�?A�1�z�2��wZ�f�u�.A��e��`��΍�
���ν
��5����_?��x?=WA?�u�<v)z>��?��%��̏�J+�>�	/�i;�K�<=5�>#��*h`�tCӾ~�þ}�� @F>Z�o?�#�?BX?f V���l�X�&> �:?�1?�Nt?x2?��;?���$?�\3>�9? W?�.5?��.?��
?y$2>:��=|.����)=�R��f芾̢ѽ�ʽ2h� 3=xz=F^E9��<��=��<7L�b_ټ��	; ����-�<�d:=�¢=���=L=�>g�]?d�>�͆>��5?���h�4�I{���~1?֒�=	Q��q��oা4�򾎢�=��j?���?��Y?nbj>g|B���G�"�$>�Ə>�$'>��a>Ė�>����X���=�+>�`>*�=��B��R��m�
��i�����<[�>5�>��>��"�?BJ>`���6;n�Hbk>8�P��q���w'��
:�//��w�8�>.5G?Ʀ?�3j=i/�4Q���b�UZ(?0�;?��H?��~?8>8ھ5�G�]M�B�C�즢>��i=6b�x��������Q6��F��qqN>5Ԡ�N��g>5��2㾐�k��BJ�r���v=���&F=A��Ӿ���OU�=���=O˼��"����׳���5J?�wh=�<���P��.���h>��>8��>�,Y�@f��>� 歾?4�=��>��:>Ԇü����F� |���>j�9?�k?[��?�ʆ���t��7��'
�Nc�yԘ>��W?s�2>�?t*>��>�1�W�����H�.{K���>5�?�Y
��x?��P��9b��X�#U�>�?���=f��>H�>?oL?Ԅ;?�?��>2M>9r�t��x�/?��?���=gM/���Լ2Zb�ީ|��V4?pm?d>}��>�V?ɲ�>�$?
c�?�H?6�8>�վ*<����>���>��B��u����7>AV?2�o>@%U?w��?��=�r�]�������ٽEL���!2?�&?��%?'�?���>�ݾ"1��V�=�b)?Q��?�j�?������=�c���@�>�c)>v�>p��>br�>,�4?筋?Uu?-[?ެs=���S#���\�����$��[�:W��="h��żM=y�<�^�=�+�=�!߼�l��ꢼ� ���[	�G��;&�>U�>��}��"�>���̯���ʆ>��;���Ⱦ�OT�:gZ���=��>�?Kʍ>����ծ=�C�>�4�>k@��>?�
?̝%?׌]��@i�����4t�衔>Q�a?.>�����+���(i��>�� �m?�Fc?^R�b�ݾM�b?��]?9h��=��þ~�b����b�O?;�
?9�G���>��~?j�q?N��>	�e�':n�*��Db�
�j�,Ѷ=`r�>LX�S�d��?�>l�7?�N�>-�b> %�=fu۾�w��q��j?��?�?���?+*>��n�W4�$w���G���^?ى�>�6���#?�� ���Ͼ�P��<+����%������R���}����$�H⃾=*׽/�=2�?�s?�Xq?��_?�� �r�c�C.^�����eV��+��"�W�E��$E��C���n��]�|.��y���G=�k>�qu3�?<�?��1?d�}��>?.YѾ�Ҿ�擾,F���- �j��=QR��Ӿ|׆<�TR>1)���F�PcԾQ>?I��>�o�>�s*?2�H��^�����/�_���V�>�Е>6�r>l�>k	>$�<߉�l츾����_��փ>��k?�`=??�k?�4���3��nd�:�+�,�*����c��>���>���>	Vǽ"���a"���,���c�����t�����S.�<>�L?�_�>�X
>�x�?�X?�7)�\�rk��Qc�O���l��>��A?�;�>i$�>J���|ݾ���>�+l?��>YF�>����Q���u�Ci����>�1�>
  ?�X>��+��xZ�ٍ�ϋ���5�k��=,f?]���&�d�l��>��S?&��<� =fe�>�!��(�������DO>��	?R��=��:>v\ɾ]��Q0{�`I��R@)?"�?x���yz*�'>�u"?`:�>=1�>��? �>	�¾�wf�W?E�^?��J?�_A?[��>,!=vF��^(ǽ��&�$�.=y!�>h�Z>Evl=E��=?!�ϔ\�3���?=�o�=	�ݼ����w<FG����;<���<�3>��ؿ�TO�P��H� �(߾aw�5N��"��q�o��,�ϩԾY����$o�b��s����t���/���x�&�G����?���?�_;mCϾ�⃿J�b�����޾>}9��l��~KT�/�׽���)�V˾��JB��^��HZ�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >UC�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ďr�1�ɿc���}¤<���?0�@��@?��'����F�<=���>�C?��U>J�4�����O���I�>�J�?���?б+=�!U�݈��tl?pXW=G/9��*q�KJ�=���=PA=T����F>Lߎ>͒+�w�B���\9>C�>�XT�Б���n���;�n>�ޕ��@��3Մ?({\�f���/��T��:U>��T?�*�>-:�=��,?P7H�[}Ͽ�\��*a?�0�?��?$�(?,ۿ��ؚ>��ܾ��M?_D6?���>�d&��t�ȅ�=B6�Ɍ��s���&V�Q��=H��>5�>߂,�ߋ���O��I��u��=������n�W�*�P�9V�=�"ʼG���\v<iS�<M����龮F��4�؉<��A�=�v�>��S>m�Z>L�V?�t?�$B>&�|;F�K=�#b���Ҿ4�6>v�~�eÑ��{0�:�=�s��nR
�����������I���@ϾD�-��EE>�ꁿ;˧�䄾=�E�Iqp�,�C?��>K���Ƨk�b�>H��1���G3����=N!�r�L�>�R�?c�?��r?�+c�~4-�ѐ��;S[���)���J?j�\;�:���)��tI�<e�����=�.�>�>�H��yG�.t�Z�0?yq?6��*����(>���J�%=`E/?,?Q =M�>��?SE/�!�罧XU>��8>M��>���>I�>���������?H�V?�D��7y���S�>3fþ]����p_=�b>��.���?��_>��|<P��������7����m<!�V?䑉>T�'��~��d����ü�|=vss?��?>�>mi?[�C?
��<�	��\QR��'�v,�='g\?�k?�5>1�z�i*о㏡��5?O�_?	I>�\���⾟v,��� ��?�6p?UX?�����jy�����Z	�fm6?��v?yS^�F��L��MW�3��>��>	D�>�9�7#�>�m>?/"�$�������Q4����?<�@���?�O<B>�_��=?�?���>jO�� ƾ}!��ձ���"r=�d�>����v���;�,��)8?�r�?+/�>S���x����=#ݒ�礫?��?���-V�<c�ire���޾V��,=�=�t$<�0��a��b�&��{�� ��H���ō��a�>��@�f���Y�>�A��c�2`Ŀ;��&���D4�d�?�O�>��<E-q��bT�Ev�lJ?���;�A"��@C�>c�>IŔ�-���*�{�]m;����d�>����>��S��'��c����5<�>��>ݵ�>R)��3彾Cę?�[���?ο������t�X?0d�?�n�?.r?�:<��v��{{��^��%G?˂s?XZ?�I%� 9]���7��j?>`��T`���4�QGE��U>9#3?�@�>�-�B�|=>���>�l>&"/���Ŀ#ٶ��������?���?�m꾯��>���?s+?�i��6���[��-�*�J�0�};A?~2>2���Ը!�/=��Ғ�j�
?�~0?2x��-�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?'�>}�?{��=�m�>K��=c㰾I�,��J#>���=t�>�i�?+�M?%I�>W�=\9��/��YF�]DR�� �A�C���>�a? |L?KVb>6Ÿ��"2�+!���ͽ�1���cH@�D,���߽�4>3�=>�>o�D��Ӿ��?Pp�9�ؿj��p'��54?'��>�?��s�t�����;_?Lz�>�6��+���%���B�^��?�G�?A�?��׾�S̼�>B�>�I�>M�Խa���M�����7>.�B?B��D��u�o�k�>���?�@�ծ?gi��	?���P��Na~���^7����=��7?�0��z>���>�=�nv�ֻ��L�s����>�B�?�{�?0��>�l?t�o�M�B���1=,M�>��k?�s?eo�x�3�B>��?������L��f?��
@zu@p�^? ��ۿ���̾bܾ��K��M=�}>�ʴ�Yn�=D���߽�ӽ�>G��>۰�>�t!>NA(>u�.>d��>���|�%�릿��a�_�:D �C�׾�Z����xˊ�-$C���Ͼ����� &<_��=dX<�|�S��xýbN=���=��U?%'R?�r?���>Yy��Th+>u����<Z���%�=��>̖1?�L?��(??�=�@��	8d�H���Bx��l������>,PL>RW�>���>���><R��XN>�`O>Q�~>��=�Y$=�*��~l=��Q>���>g�>�[�>Ìl>e�>�ȿ�`���G
�^Ⱦd����ӯ?�SZ�ɖE�~��E�۽Y��_�=�j�>E�>=����Hֿ�<��L?b������i���N6�a��>J�k?.<�=fW9�ϔ�=�Zx>��V��0�� �>0�w�c���t��;�'<��X>�f>�ju>-�3��8�ɺP�����q?|>�K6?P*��%<9�F�u���H���ݾW�M>�8�>�VD�(��s	���'�Ji�VHz=s�:?>�?�������t��N��ȣQ>��\>�+=w�=-eM>`�.vƽ!1I���/=�w�=�]>bI�>�_>g�'>{5�>@f��,����>���=�o�L6S?]�D?��|qZ�BPP���9��χ>���>	"9>��=4�@�F�=q��>3�x>�hѽ
R㽐�!���D��ވ>	�>KO=�wM5��
�=��K�)�>���=�{߽8�_�ܘ=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿsg�>�y��Z�����q�u�d�#=ި�>�8H?�V��"�O��>��v
?�?�^�ĩ����ȿ�{v����>/�?���?�m��A��@���>��?2gY?�pi> g۾<_Z����>һ@?�R?u�>�9�ڎ'���?�޶?���?QP>���?j�r?���>-��q{*��ϲ��ً���|=ɂ�4�>.o>Pu��QF�{ǋ�A�|�� m�'s����=R�X=?��>�U��lǾd�=@X���h��Ԉ����>�bW>ga>�ף>�g?���>[	�>��E=�bc��)r��×�i�K?���?���A2n��U�<���=��^��&?�I4?&c[� �ϾL֨>�\?:?�[?�c�>���>���翿~��Ţ�<`�K>X4�>�H�>�%��JK>��Ծ!5D�6q�>�ϗ>���@ھF,��If��rB�>�e!?���>�ծ=ә ?��#?ޖj>�(�>9aE��9��[�E����>Ģ�>�H?�~?��?�Թ��Z3�����桿��[�4;N>��x?V?�ʕ>Y���烝�hE�CBI�w���V��?�tg?�S�+?>2�?��??A�A?f)f>���ؾ(�����>�!?���A�
7&����`�?��?��>�+����ս�м���H���?)T\?BS&?�<���`�:B¾���<kl'��9��<K�B���>})>�]����=��>GU�=J�m��8���W<��=Di�>���=�!8�1v���4/?�=*�e����=Z9d���D�"ǅ>^�>�剾�r?��!��R��SE���4����W�L�?^C�?��?"8�-T`���&?��?!'?�u�>�E����ľ���Z;=�t�P;��,>RC�>�;<.�Ҿ8X���m���C���m"��Q<{��>�)?��1?�?��>��>�{��B�2�A��������
�mUw�r]��,���x�<������/���� �[>�hὝ��>�;?�ʠ>���>,�>�99��NF=yΨ>-G��*	_;��}= G.>�X >c&@> W�>�8R?k�����'����N���QB?
�d?�~�>bj��n����8w? ��?_t�?�v>�:h���*�ρ?Hv�>���6N
?(9=���[��<kٶ�����p���i�5�>Ebս�:�"M��Kf���
?�?#����;��ٽ$T��@_�<o{�?M�*?a�,��1<�-p��;O�H}N�՛��Ь[�R��^�%�5ms�<�%���w膿�n*��*���� ?}?����m־ۤj��WP�r7��r�>��>_�f>G��>�b�>�>�w�?���L�������\�׷�>G��?F��>��I?�7<?��Q?RSL?xߌ>��>YT�����>A�u<��>?@�>�O8?��+?�#.?�?�c)?��\>_��z5��#�־O�?��?|�?x�?�?�È�s�̽ޘ�q�Q���{�,ف���n=�qP<>�ؽ��q��H=��Q>	� ?��?�T�"��ɾ��>A�9?,�?p�>����h������<B	?*�*?E��>��	��Xs����9?�ۇ? ��ٚ��W>]�K>��˽x19=�Sd<��)��Rýv�0��Y��$Ä��Q�=Z�>���gA����=�8ż��'�	 ?Fe?��>��>�����K��m��1�=�\>oBU>>>��ؾ�-�����jg�R�z>ѐ?���?"�z=/��=�'�=X�����ӧ�%����,�<�/?�/!?1�R?i��?l=?w�#?��>���В�=���1Ǣ���?�$?��>G^6�Vq�������b����>��?⠂����<�0��t
��_��j	�>��K����+��m��a��=j�Aj?�Q��?�W�?���<��m�Ͼ����3����9?z��>:b> �?�/�����!�b���>�,?b�>3��>=�i?�k?1�F?�v�=-�e���&������;�t<=8Q?��?1��?��:?��>p�>p���5[þ���/�ԼD�(�+ʏ����<j�>�M'>��>|P�>�ʟ<�;��+��RM�T�1<h/�>4R?%X(>���>���=�6N>.�J?��?����
��E;x�
������7g�?է�?p�[?؎�9>1��xY���lz�>V`�?�ˢ?��.?N�<�c�=;��@*��AT�f$/>G�>	�	?@�	>�V���`>(��>/��=��Y����K�yLŽA�>*�X?-hM>��Ŀ/�r��ƍ����)�<߽����s��Z���L���=���~��U���{j]�����˗�:�\����`p��Q?�l�=�Ƶ=���=��F=1<̼� �<M.�=�O=11�<�.v�.%5=N�X� ������UK =A:<~�=�����˾�}?�<I?Ԙ+?žC?��y>�=>�3�掖>ri���D?BV>cP�%�����;����[��#�ؾ+y׾��c�)Ɵ�GL>�dI��>o13>�6�=�9�<�/�=,Ls=$��=y�S��%=�)�=_�=*d�=���=M�>�X>�6w?X�������4Q��Z罦�:?�8�>[{�=��ƾp@?��>>�2������wb��-?���?�T�?>�?<ti��d�>M���㎽�q�=K����=2>y��=t�2�S��>��J>���K��N����4�?��@��??�ዿТϿ1a/>m�6>x�=��I���+�Ja�N�L�3�f��V?ϵ8�^ Ծ�	�>�^�=C�꾻�ؾ6a=pWC>B�'=�� ���[���=>�R��6=��f=><>h�=�[�� �=CDV=?��=�Oc>�k��V��u�:�=w)�=E�n>�Q$>�s�>8�?G�/?�@f?+��>�Ǚ���ھ�q��ű�>��5>�+�>S=�k&>���>˘B?=?�~D?U�>N_
=c��>n0�>"	/��w��QվD���lJ�?ݐ�?�X�>'�_�K�ʽ.Z��@����D�
?{(?��?�Ȯ>Z1�XC��X	�v� �9��ɱ7��E�=3�n�"�\�Q����1��p��T�>�u?�?x!Y>+ov>>��>.j�>o`�>ʢ>�I>M�1>��,=6^T�ȓ�p_=��<�[���x�N<`��;�5��7��2|<�zļG�L��v?�4h>�/?S|�>_?*JH>ws���^>g(M�8�>��$�>����{�9��A�%Oe����og�M��=Iq>�u���~�p/�>�J�>A�>N�?_�?ek�=+��u1!��]���0�{�B=�m5>`_���'�s}h�X�_�����>;_>�A�>��z>c�x����R�Ž�O��6�@��Y�>�$��ܮ_����W��3��.F���K����3�x�>8-{��H=���?�M?�Ԛ?G?<�*��x��7��>S����=������׊�9��>�%+?o��>�y~��׾u&Ѿa�Խ�>	�S��N��M��$c0���G��h��J��>¬��UҾ�1�-����S|C�\l����>�/N?�®?Q�[�����eR�ӑ���n�( ?�h?5��>^_?�N?!���P��R���E�=a�m?��?R��?^*>p
> �H��>Kg?ń�?:.�?��?�3���l�>��k��4]=&U�4>^=�}=E���p��K�>JS?��(?�{�&�(�x�#�p
�x㻾J�����:`�g>kZ�>^x�=���=�6���;>R�?b?n��>�X?�?�a�>D���h����'?�=�D�>�s2?<��>R�V=�F��E��<*�D�SM>��S.���ý�v佷ӳ<߭���E=����W�>��ƿ��?��S>�e��?���@*��U>9�R>�>ֽ2��>V'A>�x>+�>C��>��>ٴ�>��+>͗־3`>|���!�;�B��Q��1Ѿ��v>0����.%��v	�v���9�G����#��:j��J��{�;�r�<pI�?���|�m��!,�����?���>��5?�݋�Fs�jH>���>�D�>����F�������E޾5Ћ?���?�2c>��>	�W?%�?A�1�z�2��wZ�f�u�.A��e��`��΍�
���ν
��5����_?��x?=WA?�u�<v)z>��?��%��̏�J+�>�	/�i;�K�<=5�>#��*h`�tCӾ~�þ}�� @F>Z�o?�#�?BX?f V���l�X�&> �:?�1?�Nt?x2?��;?���$?�\3>�9? W?�.5?��.?��
?y$2>:��=|.����)=�R��f芾̢ѽ�ʽ2h� 3=xz=F^E9��<��=��<7L�b_ټ��	; ����-�<�d:=�¢=���=L=�>g�]?d�>�͆>��5?���h�4�I{���~1?֒�=	Q��q��oা4�򾎢�=��j?���?��Y?nbj>g|B���G�"�$>�Ə>�$'>��a>Ė�>����X���=�+>�`>*�=��B��R��m�
��i�����<[�>5�>��>��"�?BJ>`���6;n�Hbk>8�P��q���w'��
:�//��w�8�>.5G?Ʀ?�3j=i/�4Q���b�UZ(?0�;?��H?��~?8>8ھ5�G�]M�B�C�즢>��i=6b�x��������Q6��F��qqN>5Ԡ���u�t��>�������+g��a�Q�پ���>p��]⣽��tA���]뾶�<>�Y=˛��~�1���^�����L?L�q=7 �����<����=o��>��>@@��,>7 6�����f=�7?e/>��𽔜Ѿ�:H�>�	�*'�>�_J?�Hq?!��?K޵���a�=(M��1��(��-���2?�b�>L�2?F彬���?�J�6-꾋�V�,X����><�?�5���U�?���7�n���5n>�U?)�k=!�>G�^?w��>:(*?}�?��?�&�>�y;�]E��)00?���?̄=]U��N=V+�tY��T�>�V0?��W�`�c>�rI?��>�$?�fV?�w�>�+�=������ݷ�>���>�Fc�e��r\�>��w?��C>��2?"k�?X�>��\�dm�p�!�/�K>�|�=��?ИE?���>mB�>��)?����՛<8��>��*?�ل?��i?=�?�M�>4'�>T�1? Y=D�v>WN?�tr?��T?�jS?:�?$�)?e��<��8��=���=����vv�����]�=N�<����:*=�[��=���<���<>��=i������=�װ�@�.����>3nu>.���	/>�LþCx��_�@>Ĭ���Q�����u�:����=�z~>�?���>3"�V��=P��>��>n���'?i�?C�?BA:=�b�HپZ�G��ܰ>�jA?���=��l��Δ�wv�f�p=A n?'e^?X�T����M�b?�]?h��=���þζb���T�O?.�
?6�G���>��~?P�q?#��>d�e�:n�%���Cb�g�j��Ѷ=or�>pX���d��?�>��7?_N�>l�b>%'�=�u۾$�w�bq��0?s�?�?���?U+*>x�n�!4࿿������޹Z?�|�>����� ?����˾ڭ���������K����M����OĤ�޳������H۽6��=�?&�t?MWr?n�^?�m��d�)p^�L4��W�֮������E�QE�*TD���o�������o���%�@=�5j�}?�~�?�!#?��=�	L?6y�O�������.�=�����v=L���P� ��uý}�����{��ƾ��?K�>e��>@N/?-R`���F�6U��M��$
���=C?�B�>F�?v��=���=}��9�����`���n�M1u>�&`?��K?�}?Jp�mv/�I?p�X�)��I���Ő��qz>�,�=���>�1�����y$���3��k�m���V��C����=�:?�>]ԉ>� �?�-�>p��a����_�J-���=<��>��a?��>��s>��u@�b��>*�k?�~�>�ի>���!���v���޽`��>;L�>>�?�^h>17)���X�@������2q6����=��f?}�d�eg�>BT?r6H<m�;��>���T'�pU�!��A>=C?���=�V<> bž���+*}��ዾ=�6?�!?�M���m0����>.@?���>�k>�)�?�X�>k �"��=��>�W?5W)?�]?�g�>-#=Ʃ>'$}���[��K�t�{>!�`>Ό�>�Y>������hq�y�Q>s�q=2�R�V���!���_=!	��J�_>l0>��ӿaA��$۾�3��Uƾ������v���"Z���t�7�þ��i��gy�ŷA�8:��)g�T��W��BkZ���?�)�?�`��'��.���炿��	�j��>?栾(����Ӈ�Fڿ�#˾<Ѿ
Ⱦ�*��iB���d������'?����c�ǿW����:ܾ� ?iV ?�y? ��}"�f�8�<. >���<�ɚ��<�����ο'y��/�^?��>W
�*[����>�Ƃ>��X>5$q>Z��m)�����<?�-?���>�3r���ɿۊ�����<���?�@�A?�(�����IT=h��>í	?y+?>N]1����?����>�3�?/�?�M=P�W��	�-ge?5 <��F���ݻ{��=���=K�=��e�J>���>����&A�@Kݽ��4>���>~3%��sR^�i��<�G]>��Խ�Ĕ��ӄ?�s\�f���/��R��;_>`�T?��>+g�=\�,?�3H��{Ͽ\�\��*a?�/�?��?��(?ȿ�E�>��ܾ2M?�:6?��>V&���t��o�=e��r���Ⱥ�JV��F�=w��>��>��,�ɔ�̑O��9����=m�|ٻ�y�:�2l&�zXL>��t�þ��fZ���L=@�z����O��$꨼���<6\�=
\�>s��=�E7>ao�>.R?��q?�Ʒ>nE>�xý����X�߾�|K="�w��Q|�Wv�8Ϫ�&�������p��p$���5�w��������6�
��;Y�]�ܚ��ný�Гf���S�:5K?�R>)�־eW0�3��>+�۾%ϑ���_���=<y���4�~\���?�?F?+Vx�b�D�c1��f���N=��t?�, �����q�?"1>m�����_>�͒>��<t}Ǿ�N������C?g�,?{Y��Yh��{L�>�=�Y�=�tV?N68?�1e�dV�>-�?��þ��u��_>�M�>`�>1�>Ev�>�k��Ś��8-?�0U?�ꀾ��־6��>�L���0��kN�>S�V>2��Q�=��>�~8���ýZ�>NT>��d�*W?ܱ�> �)��
��0������<=��x?��?�9�>eNk?��B?<�<�0����S�����w=��W?�1i?��>"Ɂ�hоo��W�5?��e? �N>�h����.�*B�?��n?b?�Ρ�zh}�������[6?�v?�o^��r�������V�?�>�\�>���>+�9�th�>k�>?�#�4H������)W4�$Þ?�@���?�m<< ���=�<?R^�>ٲO�WBƾ~{�������q=9(�>T���fv����O,�؅8?���?���>�������G��=�P���,�?��z?09�i�=�5�b����L.��YU>&���� >�$�|
&���㾴�D�-;��;n�~y}>��@j��t�>�����ڿ��ȿ$u~���-��J:&?�a�>,�=�	��N�4�/=���"��@T��þD>�>6>Hʕ��8��F�{�ǐ;�Y�����>-	����>�VS�Xõ�>$��{�:<���>ר�>{��>=����D��0Ù?h���.ο���o��M�X?[n�?	k�?T6?�G<{�v��T|���JG? fs?5�Y?��$�v�]��2:�%�j?�_��xU`���4�uHE��U>�"3?�B�>S�-�_�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�TҒ�¼
?V~0?{�f.��_?q�\�0�n�>�-��ڽ���>#\��gi��jR�?/��zb�Q����N�?���? �?�$2�H�E�+?_�>=V���)Ǿ8HM=�b�>@��>��D>1�ϽmGD>����+�GZ#>a��?�J�?�6?�䐿Ġ��Cm6>�j{?㕶>/��?_:�=�E�>w�= ű��%���Q>!��=��#���?�L?�_�>1�=�M7��/�mE�QsR���C�B�d^�>�da?�\L?�Mf>1ݿ�c�!�	� ���e�)����_�?����Wѽ�L7>W�<>�>�K�12վ��?8p�1�ؿ�i���o'��54?(��>�?�����t�7���;_?4z�>�6��+���%���B�Y��?�G�?7�?��׾�R̼�>�>�I�>��Խ����Q�����7>3�B?[��D����o���>���?�@�ծ?Ui��	?o��P��Ia~����( 7� ��=�7?�/��z>���>Y�=ov�̻�� �s�깶>�B�?{{�?g��>�l?u�o��B�%�1=�L�>K�k?�s?��n�_󾧲B>��?!�����JL��f?��
@lu@f�^?��ߏӿE����l��+Ѿ�g�=U��=6��>K(�Ѭ���<��;<���Zr=��^>r��=�	8=�h�>�*w>�'G>�x����#��λ�����:�4���qk��\D��E���y���?�h׾���k�d�313��|��҃�&౼-�V=�#�=N�O?˝Z?��?~�?P�,��>�i���?�&�<�I>TE><4?�V?��?o�0�;N��Bi��q�������V�4	�>0v+>�E�>%��>Mٱ>4�=)?)>7�R>7�9>�$�=<+�;�����<ւH>L˶>���>Zww>_.>J>�]���#����`��n��Sɽ�ͤ?� ��;�G��d����x�OG��g"�=,+?�!>%�����οC�����E?H������! ����= �+?Z?>�ΰ�s�]�B>i�'���k���	>���qn�4�%��@>!?�x>�n�>8�3��>2�"h�A����>CC<?kپ�(���p�KM�q���7�>Oۖ>#�����#������Nf�6��<��??-�?�^�l���M�F�d9۾=�R>Y�>i�Ž�5L��o>�&��g/��*��Z[��5�s=~/e>A?��1>N��=$�>_���'I�L��>��>>��3>5�@?dz$?�)�}���$��#�,�F~>D��>l)�>@>�zL���=	�>~e>V�ټ˹x����pVM���P>;�Q���Z� *~�my�=!T�����=۹w=�����>���
=��~?�{��f∿�뾍s��kD?�1?Vː=��G<Ay"�����T�����?3�@sn�?Ry	���V���?�B�?+������=os�>�߫>GξU{L�m�?�Vƽ�آ�ڍ	��"�S�?��?ܖ/��ȋ��l��.>�f%?��ӾMh�>}x��Z�������u���#=Q��>�8H?�V����O�{>��v
?�?�^�੤���ȿ1|v����>T�?���?j�m��A���@����>=��?�gY?oi>�g۾7`Z����>̻@?�R?��>�9���'���? ߶?֯�?x)H>���?��v?c�>�Sӽ�-��a��6��c	=l�D���>#�>�����#O��f�����O�`�C6���>F3=���>K���������=�6���L��:Xo�\�>Cn>Ӹ3>���>��>A4�>�/�>��~=a(��U��눁���K?���?E��h2n�C��<%��=V�^�%?EK4?E�[�8�Ͼب>��\?���?z[?�b�>���$=���忿�|����<S�K>W3�>�D�>\���QK>4�Ծ;2D��j�>�ї>N��+Eھ}/�������C�>7c!?0��>�ۮ=\+ ?}(?;9>�Y�>*`1�\����-@��R�>@�>\?��{?�F?�c����+� -������BZ�p�E>>Nm?�� ?eˣ>�����0�����<""B��b0��~�?�
o?>=�`��>e$�?�1?ne-?r1�>z���H�fp�����>O�!?�\�e�A�9&������?��?��>�9��
Rѽ�fڼ����}��<?�y\?
B&?��)�_�����[
�<�F;�H_{��y+<a�!��E> �>P������=��>Ev�=�8i��#6��kl<:m�=C
�>��=4�0�H����=,?{�G�ڃ��=D�r��vD���>�LL>����q�^?�j=�{�{�#��?x��1	U��?���?�j�?�����h��#=?B�?�	?�!�>�J���}޾J�ྒQw�mvx�~v���>e��>0dl��ԏ��-���eF��� ƽ	W0�~��>��	?q@�>��>�/�>���>��B�����v����<�n���ɾ.��(r���v��\\��)߽�ͽ?�⽶��������]�>�c��(��>�W?��>(�>�2�>�����>M�j=P�>-��=ɇ�=�`�>���<T�>}!�;�R?�����'�2��򃧾��D?�
a?$��>�"��h��#�D�?�Ԑ?&a�?P�q>��e���)��3?V  ?�~�xh?O')=�����(<��������>�L��e{�>�����d8��Q���w��A?��?�ƪ�&Fľ�pǽ�䟾�r=)��?��(?�*��BQ��cp���W�:S��&���c�2���w#���p�鷏����D�� ;(�a�=Z*?�W�?r��mK��\Yk��>�`�d> =�>�)�>{Ͼ>i�L>�	���1��/^�1�%�6���?�>6\z?�g�>9K?�6?ŧ_?Y3?>>��>Ҿ0i?JiP=���>�*�>o�?p�?�	?��>��&?��X>h��u��נ����?	KN?Q�?���>1?����Ũ�= �>���=�l���ڙ�w^P>ؼU<�:���'��Hs4��E]>}�?Q���r8�����)m>G�7?�R�>.U�>�M���R��!�<��>��
?	�>]b��t�q�����>B��?����A�<��(>��={���J:��=ht��Ī�=8~��xL1��d!<�O�=�={����E�:ȉ[:�U�;jƬ<u�>;�?ȓ�>�C�>m@��� �=���f�=�Y>uS>�>�Eپ�}���$��V�g�^y>�w�?�z�?�f=v�=���=�|��BU�����:������<��?J#?,XT?M��?K�=?tj#?�>+�VM���^�������?�?�|�>\��}����ÿdbX���?�>�#b��h;o�N�{ ��׶�	��>��-�����C����|�������hW��t�?O=�?����� ����޾Jᓿ�eH�: ,?QP�=��>�*�>v\6���T���9��;�=|'�>p U?�P�>u"e?�Ar?�[:?��>��8��[���|���� =d,R�ɩ>?\Ax?���?��2?o��>>+K>[_��1�`	�Z�
��OɽG{��Ն^=��|>�ac>��>�ۧ>��u>��E�⽥V�X����Ш>�E?�~�=���>���>�U>�H?���>��>T��m���8k�e���Cv?���?G�#?�r=i����H������>��?�Z�?��)?k�9��/�=&h�h���;�c����>���>Bɞ>��=��1=/!>��>p��>�G&�g�� 3���IX?�"G?���=]Nƿ�g��g��f�۾<>�j��H���P=�Z�����=`S޾1�s]��_��i�b�5�o��Dؾ������4��;�>G�=�!>�l]=)"h=����.=o��F,=`d�v=#���e�s˼��b���=��\����=E��=~b˾��}?�EI?,�+?�C?�y>̫><�6��
�>����S?�U>��N��#��04;�漨�D	�� �ؾ�{׾@�c�����ZK>�I�G�>��2>Ĵ�=Ʀ�<G��=�s=�F�=��\���=x9�=�c�=��=~a�=��>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>?)4>ê >TS���1��FX�Db�4�Y�>�!?5�9�[z˾ǡ�>T�=�O޾Y{ž �7=��8>V�O=�����[�t3�=��x��uA=y�l='ԉ>��C>Y��=t����=�\2=�=��L>Dn��`�;�Nj,��7=C
�=S'b>��&>(��>��?��4?x9}?��>:����{��\����c.>��8>��>��<��A>S
�>��&?�*?�_H?Z��>�C�<��>�=�>I6,�i�r�jپ����'#����?��?2�>��;�ֽ���G�M���#?p?V�?�y�>F�	���޿�H��<L��g��!��S�=�T�!>U��t��Xj��gd��y�>_�><��>A��> 9t>Q��>��>�v�>e>�K�=f?>oTc�FP˻*gI�� 8=;E�=�	�=-��=jF�=M��=�������<mc\>��̨ѽ��P�.��=��>�e>���>�o�=�����_/>k�����L���=�;��.B�!-d��@~��/�t�6���B>;!X>����h/����?��Y>�?>t��?�;u?� >M�W�վ�C��0(e�QkS��=��>z�<�Hs;��M`�M�M��sҾ�Y�>Y3u>l��>�l>�D�v�,�_mJ=�:Ѿ �6�=��>B�ܾcf	��
��l4b����n��M�\�����9%?Q���(Us��&?U�>? ��?5%!?Շ9;!���J>Z=w�D]=Ց��	5�7���t��>��?�c&?c�e�E��O�˾*ý>͹>KF���O��t��N/��������:̱>�ͮ�{Ӿj�3�����^��ʽD�
)l�Y��>ΧM?:��?��g�yi���FN�3Y� Z�,q?�h?��>8�?�?>a���뾲���P��=n�m?���?���?ɻ>���=�Gv��{�>��>.ޕ?�9�?0�l?Fv5��s�>6����W>t�d��=�4>�=���=�,?��?�?-*��~$�U��>�d�d�Ф�<�x�=7�>�)�>9�Q>B[>M	�=_+c<��>�ĥ>�g�>��l>徵>�%�>G$�������&?G �=9��>P�2?R0�>mf]=΀��3E�<��N�X�A��9,������彺}�<Ќ���T=��ɼ[�>�>ǿ$�?SuT>�Q��?jq���6�+FR>��R>0�׽���>��F>�U}>6Ů>�d�>_O>�>�?'>�<Ҿ��>Ҟ��� ��D��WR�LѾJkx>3b��� $�E
�m���� N��V��]���j��L���E>��!�<�K�?[��Ti�H�(�*Y�Nc
?N�>d�5?��������
�>ym�>�ލ>|)��t��������8ݾL@�?[��?�;c>��>p�W?"�?�1�"3�'vZ�!�u�x(A�>e��`�i፿Ӝ��:�
������_?��x?�xA?H�<�9z>]��?��%�Pӏ��)�>�/��&;�F?<=d+�>*����`�ٮӾ0�þ�8��GF>��o?Q%�?Y?TV���l�7Q'>�:? �1?�At?��1?�;?fY�&�$?�24>+_?�N?&M5?l�.?w�
??�1>4�=�ĵ��#'=����̊�?eѽrʽ�J��1=BV{=�؞9i<��=P£<֎��ۼ��;뺡��m�<[>;=�+�=�Z�=�ͷ>��^?i��>`9~>#:9?��нe�3�
"���r9?��=/����Ń�����Q���=�
d?���?X�M?9Ё>X�I�#f@�<3>+�>$&8>�ق>���>��3��>��J�=���=���=��=5�����a�����٩�<V��=?�>�w><��9D>b夾;o�6@z>ʤ[��o��nGB�!AF�R4�u�z����>/oO?*??
�k=��9:��a�Ț$?��7?].N? �?�m�=��پ4�>���N�]����>z>#=���M���#栿~�=����r��>&���w~�Ɖ>~U�"���9�h�$�A�JC�T�>lN�ja�=?,��s���F��F�*>��>D�������@���ՕH?U.#=�&����@�Z�Ծs�>�)�>���>a᯽wU}��d<����B�=\��>Wgx>�ĺ?���Fa��q��5m>MD?��l?:z?]+���p���"�+gӾ�(:���d���?,�}>v�?��y>��=��ݾ��t�X�B�U��>lj�>z�$_P�&����@��qb(����>��?��I>��>E�n?�?�@n?�|2?-�?j��>)�8�Ⱦnq)?�Ȃ?��I=ʨw��]�����N�@��>��0?'3g��>B�?l�,?�L$?, N?�k�>F�->W誾��'���>���>P\a�����"�>0�@?�[�>�2A?̔a?�n�>-A�
վ�+��d=��M>?'e1?�&?���>���>�O����,��z�>!W0?�Q?j�?(j;>��?KD�='n6?�/�WE�<�����h>��q?�/l?�Y@?�R?�;=��s�=���"���4����w�>����?�*$���::�$����<��*>��>e98�[�$�3��W��>M�{>���>o6>쑺�@
���f>>��U���8Ɔ�m,=��p�=각>�:?H�>��"����=([�>���>��HK%?\`	?�?�t�:��_�_�վ�N���>>>C?��=B�m�t!��_�t�1^k=�o?��Y?��T�j���Q�b?�[^?���Br<��&¾�c��z�lO??WZI��Ʋ>y�~?f"r?4��>�4j��m�������a��Gm���=&˜>UN�Yd�S��>V�7?P��>P�a>Ɗ�=�ܾ��w�ʝ��~�?=�?�گ?K�?Va*>�/o�n.���������:]?���>+H����"?L+�cϾ�)���
�����&���W���>���"~��v�!�\?���-׽�F�=��?}�r?�Zq?�[_?k/ �zc���^���~�%,V�<��,��F��D���C��Fn��u��t�1;���A=�n��dJ���?Hs?ǹ;�G}�>�X����4��hj�=�Q���ls�4YX>`6ν
c�>���==z����c�(���݈	?@��>�>��E?��;��C��A��DL� �xĺ�U?0��>�[?Z��=V�?�t�⽖3����>�<V�y>��c?g�M?�o?�=׽�.��G��=� ��r���Ⱥ��B>S�>�j�>q�O�����'�;�;�ɕj��.��!���e����=Է0?��f>(��>��?��?6W�m�����t�\�*�gZ<���>;`j?w��>��>������v��>�l?���>�R�>G[��zD!���{�.C˽(A�>&�>��>ޘp>ؑ+�
\�Z��4�����8���=w�h?����Ja���>�R?}.:S�L< ��>av���!�Q��^�'��>�\?�ܪ=	<>"�ž����r{�m���.)?*�?X����c!�a�>��.?���>��s>'Á?W��>��;��ֽ,?UR?�3C?�~?\�?���=�
��ʽ��&��J=�h�>S0@>щݻrh&>l��oa8���j�bK��P+>�d��눏��cN���?�R=�Z��� g>1Nѿ�jA�y�K�����@/��|�@)��X[��x���'ǾF��3����.����'�H_Q�j7o���c�$��?G�?��g�����Z�Mv��1��%�>�0W��������8,��"���`ݾ']���a'���7���Y���l���'?)���R�ǿ����>EܾB ?B> ?\�y?��1�"��8��� >��<�n�����o����ο������^?��>A	������>Ҙ�>��X>�\q>����ٞ���<��?��-?u��>�r��ɿҊ���:�<���?��@A?�&�;��s�h=G��>]�?�S5>3C5����������>$"�?O�?ٶ@=�>X��A��|d?��2<��E�@���P��=M��=�#=�g��_K>�Β>5��?���佽�/>G�>����f�[�e�<V�`>&ZϽUl��4Մ?*{\��f���/��T��U>��T?+�>e:�=��,?S7H�^}Ͽ�\��*a?�0�?���?%�(?/ۿ��ؚ>��ܾ��M?]D6?���>�d&��t�օ�=Z6Ἂ�������&V�{��=V��>r�>��,�ۋ���O�J��&��=*��>y��n�A�d5����"
�=�)޽J�<�sl�X&�=m����h��#l������q��=���>J�2>��N>a�R>�Z?��p?�1�>��r�%߽�l�����b�ؼH]���&,���f㹽��������jľ���f��Y��e ��W!��PW>[�J��S��q �C���^��b??YP$�6���h��?x�=P��X��	*�ۍŽ�����e,�1�z��?��Z?)�G��M��(��bս�fQ��5�?Wk�<.���l
��N:>�M�=Q�=O/�>�M
�w��>y�����-0?� '?�X��y}|����>Hfz��X=̟?�d	?�{�:��\>��?'ͽ,T���N>m�q=џ�>�h�>��s>�������~�.?ܓg?�L��̳�1Î>]ܿ��,p���
�(��=�5��~嗽�"�>U�$���T��<��[���j=h�V?5v�>�*�{�������/��?==b�w?�4?2-�>p�j?!�C?���<)����S���	�zu=X,W?��h?O�	>Qp|���ξ���F6?~0e?U�M>.zg��2龞.�#��8?�m?u�?QX��S�|��.��7�ļ5?�vv?PU^��J��_��ppU�R'�>��>���>��8��>�>��>?$�J&��]����J4���?�l@I=�?�ڋ<��[�=:�? ~�>ASM�"�ž�ߴ�1*��7�r=g
�>i⦾s v����a�,��8?�r�?x��>��B����=,H=���?x�{?�N���,�<,�V�N�'�޾6*�
��>h��=q�>�¾W������B�����	=�-�>�-@�+��(�>uG�=�����������5����{��� ?9y�>�,���������Z�u+�����9��2�>F�>x唽k��I�{��a;�Na�� ��>�1�'�>o�S�����(���m�8<��>N��>
��>Aخ��Խ�t��?�b��`)ο�������|�X?8L�?	_�?�\?hD<w���z����$"G?3os?�Z?%[&��]]��a7�
�j?_��EU`���4�HE�U>�"3?SB�>�-�Ͱ|=>D��>/g>l#/�N�Ŀhٶ����C��?��?�o꾧��>y��?�s+?�i��7��v[����*�T�+��<A?{2>����<�!�0=�1Ғ��
?�}0?�z�..�v�_?��a�C�p���-�e�ƽۡ>+�0�0c\�"Y������Xe����PAy����?V^�?=�?2��##��5%?��>L���L8Ǿ��<��>(�>7+N>�G_��u>	���:��h	>{��?v~�?#j?��������gW>�}?�$�>��?��=�d�>{s�=b밾�c.�[#>�,�='u?��?��M?�T�>s]�=��8�[/�WF��?R��!�`�C��	�>��a?ɁL?�Fb>���n�1�*!���ͽ@e1�E��T@���,�d�߽<55>O�=>c>��D��
Ӿ#�?Ip�ږؿ�i��q'�/54?<��>��?�����t���;_?mx�>r7��+���$���?���?{G�?>�?l�׾#_̼�>=�>VG�>.ս
���H�����7>�B?��D��u�o���>���?Ķ@�ծ?3i��	?���P��?a~�*����6����=8�7?�0��z>o��>��=�nv�������s�C��>2B�?{�?;��>�l?�o���B���1=AK�>[�k?�r?�`n���Y�B>��?���$���L�{f?��
@?u@;�^?��8Tܿԕ��W龾�������=O
}<t�Y>��N��=7��=��7=n̼@��=�FF>cEY>��>J�U>"�>�.�=뷅��D%�����V뎿&�9�����H�^���㾭b[��M���Ѿ);־c&��>�W���b����r����I��=�Q?@�U?�5p??�/:��>!���t=�K� =�t�>_5?U�P?u�.?��@=3W���a�������:����Ʊ>n�2>	��>��>�+�>��C<vl[>S�R>lu�>���=U�;�Y;<��<�d>��>�>V�>*s�>���>�U��?,��q��o�x��8���P�?��1�:�r�b��UM�<J㾉�>�e^?V��=���c��=Jÿ0�%?��������7= �뽻ǻ>�Zc?�'[>b����d�;�q�>@�m��^�����=���=��e�}�E���>�?�р>
�}>d�7�#�=�شP�1ڮ��t^>l�=?�Ҿ���l�s�V�2�J#龺U�>G^�>� <�O#��v���~��:[��ن=��<?��	?��ǽ������Z��R��<�l>a>1��<gp=p�F>o^J�Wcý�*c��4�<�f'>K�i>K�?��>7=���>nu��d5�ps�>x�:>!t7>XM9?�{(?*�'���̽�B���J�YT�>�t�>L�>_V>s�=�Y��=T��>��U>9���!���!/%��w��?^>ڪ6��+U�󛥽�=�3ս׫>�*�=Ҳ�5�&�L"=�~?���(䈿��e���lD?S+?` �=	�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�y�#=Q��>�8H?�V����O�d>��v
?�?�^�੤���ȿ4|v����>X�?���?g�m��A���@����>;��?�gY?roi>�g۾9`Z����>һ@?�R?�>�9�~�'���?�޶?֯�?1�Z>��??�m?%��>V�}<�v-�#��.���;>��p��ގ>��4>m��q7S��t��䱀�h�Y���
�X'>�Α=͙�>u��I��� �9>CR_<�ر�>rν҇�>�D.>l��=�ܠ>��?���>
��>���=��3:킙�ܵʾHL?���?����@n�x=�<�%�=_�d?m�3?�vM�e	о��>z�\?�ƀ?f#[?KK�>���
R��w�:X��݀�<=�K>�E�>9�>N����K>��Ծ�C��C�>�
�>���{ھ����4���!�>�%!?���>��=�) ?L%?Nln>�>��A�ᑿ��H�P��>_��>??�~?t?# ����5�&����Π�g�Y���P>G7v?�?���>]h��'
��#-;�'#��ӧ���?eoi?z���	?��?�DC?93??;�Z>��ٹξ�~��x�k>��?���qE��)������?"�?�,�>�IȽi��Gcμ-���
� !?��S?�)?o��7^�%徾��<�ך�%A�<�<
^<C�>CE�=������=Ћ>|3o=����7�:����<���=Ë>���= ,�Z��=,?N�G�܃���=U�r��wD���>�IL>1����^?Ak=���{�����x��q	U�
�?͠�?<k�?�	��֝h��$=?��?	?�"�>�J���}޾Ô྽Pw�o}x�uw���>j��>|�l������ҙ���F����Ž��
��U?y9?&?��>�҅=7�>¶x�[�
�ۼ��վl�w��� +��0*��s=��ؾw/�$T���-߾��o�u��>����k�>d]+?Ɗ�>^ �>Eq?��<-�k>�{C>���>P��>a9�>7><>�)}>��=�½^HR?�H���h'���C��:�B?)�b?���>1]����o��k?���?��?�y>+�h���)��u?�{�>˗�љ
?�,="{��黮<�ܵ����Ű��	��L?�>ʞݽ�:��-L��-h�ӌ
?v�?-'���˾��ѽRX���Sq=>M�?l�(?)�)�&�Q�/�o�Q�W�L�R�0���f����$�$�ԛp��菿tA����2Q(�,=��*?�A�?o���9��@����j�Ɛ?�?7e>޷�>\�>�4�>SI>y	�202��^�C'�����I�>?�z?��>��A?��Q?�Jx?:_E?��>��g>�)��z?L Y�Emk>�@�>'�:?. "?�	?���>F3G?���>2V>B �<��&�A?��9?���>V��>7�?Gl���S��I3=�N>��x�����x�O����=�08>��h�����R�O?�[�#4�$��ldi>��8?x�>m��>ퟄ�� y�4ڃ=���>%?H��>� ��l�4��،�>=�?�nӼ6�=�n>x��=UD伏˗����=���e�5=�\���;��GW<yҥ=�g�=�0	�~�4<���<e��^�=h�>��?���>\�>� ��#� ����J<�=�<Y>S>$f>Eپax�����\�g�oFy>�q�?�t�?�kg=�=�z�=9����v�����=�5��<��?�E#?�IT?ӓ�?j�=?&x#?å>-.��@���W���
��J�??K?t�>��ʾ�,¾W�пI�����>6�4?:�z�Ѓj���$��ި���)�B��>֛��6��������[�s���,�uռ����?�0�?�0�<�Hv��2ֽ�b���S��vt�>8^?+���7�>���O0��i�3�+�=���>e*)? �>�g?��m?�j?`?i�ܾߏ���<��r��>�Dݾ�1 ?n�?���?��,?�(>V��=�½����l�	�n�1�De����*V+>C�=w�>� ?T��>���<+<e�W�P�Iq�79=��>a�?���=-:�>�C->+��=m�F?=�>�P�����l��f��Ǣ	�6�s?�P�?6�)?@/F=mH��\E�S��2ֽ>�è?���?c�*?r�5��`�=I	�Wr���"r��K�>p��>�+�>o3�=I�d=EE$>���>0t�>p�+�<5�u�"�&?*CE?�	�=~ŵ�X�a�B*���Y����0���I��p���ɾ�
>w�T�]�'���^����k��A��
��v�!�a�)��?�~�=�b=~��d~Ͻ�Jk���=9�=F���� >����>_7n�P�=�災xL�=��=� �=��:��˾��}?�:I?��+?U�C?E�y>�@>��3�ۛ�> ���B?� V>L�P�Έ����;�n���,��)�ؾ�s׾��c��ɟ��F>�sI�e�>�93>P�=�T�<�	�=s=M��=�.Q��= '�=mN�=i�=T��=��>�U>_6w?7���ݲ��=4Q��V�k�:?�9�>9�=M�ƾ@?��>>�2������*c�{-?h��?�T�?j�?�oi��d�>���S⎽p�=����<2>���=�2�9��>��J>ރ��J��⁳�m4�?s�@E�??�ዿg�Ͽn\/>�z�=-���!i���bf������;���>�)��>�g�S�=쐄>�g�>�{!����Z\۽��>=�:`R��id�	�2>��;�&�=+��=���>��m>�YD����)��<�9>F����9@>Y9����)>������=�� �������=6C�>��?;� ?�=g?���>U\(=��D����>d�9���>H/�=w�>��>.4?C��>��@?�x�>��=3��>�:�>H�V����ž"]`��ϻ�_?!�`?k;&?G��<�� �6-�uڽ���>�3?��+?���>,���꿟�"�~F���^g����=	ýc��=��m���Ὤ�����`fݽ��*>��>��&>�P��â�=���>ɣE>x���J���kt0=�51���RQc�! �=��Խ}ab���=;���-�=2��<"�ǽ���=�'=7�=U��>Q�>c)�>(v�=���� .0>�$��b�L����=l���,B�w$d��~���.���5�rC>�Y>Z�����(z?=�X>e$>>=l�?�Su??�!>S��cpվ���W�e���S�+�=��>X�=�&�;��Q`��M��vҾ���>\��>h��>*��>	�)�X�~���>;&ྫྷ&:�Fd�>g�B�<��e�Vd�������������kR?3mp�=m�?��T?^��?�}.?�������1�> r��<q�=Z��Y�Q�`h~�S?��?Q�>�u�,�n�ؾ;<�	�>M�r�NBO���*'����f�¾�o�>q����˾X�6��s�����:}4���k����>�L?�q�?��=��Uz��J�c�� �n� ?Ĺi?A��>ٲ?�?}�i� �վ Hy��mk=�k?��?��?�=*>���T��>�y?]�z?�O�?�s�?���z�><�M=�N�>+���YV��^�4���6)=o�-?�1#?�&?�������������S��/=�^>bJ�>�c�>�	o>�0>WV�=��g=р�<�A�<Q��=u��=��>�,�>���P	���V?���=�\>@I ?�R�>hT>�>�5�=�鄽�V�И5����=M��=�U�;sJv��X(�[��k�>PvпB ~?��2>Gξ�e#.? �����<�9�<܋8>7;��ފ>-�2>�>�H��>@?`m�=p�b>�>�FӾC>����d!��,C��R���Ѿ6}z>�����	&�ϟ�Bw��cBI�Hn��Rg�mj�>.��,<=��˽<%H�?`����k�.�)����7�?�[�>�6?�ڌ��
����>���>�Ǎ>�J��V���Iȍ��gᾦ�?,��?�,c>	�>�W?,?#]1���2�ZrZ�q�u�a4A���d�(�`�jՍ�Ҡ���~
��m��l�_?��x?�lA?'B�<Tz>ԥ�?!�%�͏��&�>�/��<;���==!�>��Mwa�K�ӾQ�þ�O��F>kqo?p$�?�W?��V���F���,>T=?��6?�cq?ex.?��:?�R#�V�$?�,(>�A?�H?��2?��(?�	?��S>�>~��;Qus=S���� ��e���r��3�#��*=�ɀ="��;�~����<9G�<É���_#��`�����=	�K=�g�=���=D@�>*}\?��>b�>��C?�¼����1ؾi�+?<n�=�?f�{Ǵ�[�2�a�׾�0?>�J?��?W�[?g�>�A��l����=� �>\�>/8>���>��$�_�a,^<<7�=�$>�y1��1޻�_�����;�#�e� ;|%>^/�>��z>�u��^&>�آ���y�Uc>։R�ƻ��R��?G��1�*�v��I�>F�K?Z?L�=����!���e�N�)??a<?M?}�? #�=��ݾ(�9�zUJ��M�)\�>���<���b��������:��?7;[u>�����L��-�>����½e���B�[T��{�=y���1>�*�����������+>A3>�u��z*�,6��:���B�F?O�=�6��8>��ĸ��h�= ST>���>��������L�Wݨ�m�)>l;�>�E>����Npھ��R����+�>��H?��r?��?V$s�ˮ���d�[��X������Y�N?�[�>@�	?�F���ϭ�o�E��r�Pl��+g�O5�>�;?�d9�\!;�ʟ�d��Al9��>�?g���?�?I?�b�>��b?��?Rk�>g�>Ȃ���ᾢ9 ?���?�y*>�?=Q:̽�u;���l��Ǳ>�{?�c;M��>j�?��?���>X#?��?��'>����k�ZM>��>�P��,���l�>�xw?q/�>G�7?#��?��>	M`��ܾ����>S�>@��=�j?�t?~A ?4�>���>�o߽2�2<I��>T�@?��z?q�^?�������>�e�=�\>	R#�p~�>3߫>�, ?�c?��|?t�E?)��>��=Vڽ�Z�%1�2�%����=�w�<���3�=ƌ�<�I��K�t��=I�_=f��=��ս��	�ͱ>�e�>f�s>%���1�0>� žK���<A>���*��ӊ���9����=���>��?bu�>+�#��ב=/��>W,�>���}(?v�?�4?��P;ˈb���ھ�ZL�`+�>-�A?b��=B�l��x����u���f=��m?�^?�W��L����b?� ^?���)=��þ��b���{�O?A�
?�G�Le�>i�~?��q?���>�e�An�����db��Uk�T<�=�x�>�4�~�d���>Wy7?��>;�c>���=}C۾L�w��z��x4?A��?Q�?v֊?2	*>y�n�5�p��E���|�^?��>!<����!?֔�Eо�v�����_��������#���֦�:�#�ׄ�iؽ�Ʒ=��?�xr?�$q?e`?o ���c�e�^��L����V��Q����/@E�� E���C��m�۽�5����ۙ��;=n�H��,5�b�?=n&?FS$���>��b�p��S��@�>v2�4�w�<4>� ��Lj�=��=-9���]�����?��>�>��U?!�L��1<�9wY��`�����g�>�&�>�A�>�]�>A.��Q콈�>�T��s��N�%�}M�>W�`?�J?c/h?Qb,���=��\������8�R���mK>�-�=BC^>u�c�����,5�J�H�u]u�XH��ť�5��Ix�=�A?��>���>��?��
?��0����۠�d3N�Aܼn��>�P?�]�>G�\>��	H�ø�>��l?x��>Q�>����A^!���{��ʽ�"�>f֭>���>s�o>�,�� \�i��[����9�Q�=,�h?7�����`���>�R?�!�:H�I<��>�v�\�!������'�B�>�x?y�=a�;>�wž�"�J�{�
9��	)?*?�u��F(���>r"?�G�>�l�>��?1ޙ>^�¾��6��?��^?��I?\�A?n�>��=۝���ɽ~'�U^3=�1�>e]>��p=���=v���"Z�cT �0C=+�=)���⿽@�;�A��/�"<��<�.>O�ȿ��:��	����D�������^͚�7��=E�r�A��'v��꫾kI����u<�t
��\v��K���"?��d�?8�?�K�6ʟ�����0������>�� �ꐜ���龍%�����y^ؾu�����7�X�T#}�K�o��^3?2k��)ǿD?������?Q�?�ߊ?�`����vA6����>�$=�"�=�q���Ǖ�p�ѿޱ����Y?��>���a���]��>mx>���=�u�>.�)��i��i��zH?�
?w@?��7�Q��껿��}</�?�@�lA?��(��n���W=���> �	? �?>�H1�`1��F��g,�>�5�?��?-yM=�W�<	��e?�I<H�F�t|ػ�G�=�ߣ=[�=ʥ���J>ڀ�>N����A�۳۽=�4>�>"������^��y�<�]>�dս�锽5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=\<���ǿS�$�a.���6�y�<cL�;;	���Y>���>��)=�����۾F೽x����p���>��?,m?;�>?��e?��>�'8�����#�����UG߽'C�Av�=�ý��ݽ+������<@���쾊��@H�z2��|,�ڂ>�Of�'蕿�A��M���S���?~�=�cW��:X�L�>� ����}��>?=��S<�B�'>���Z��L�?ΦV??�C�X�P��6���H*��f��^;{?4��������K�>�m�=�� >� �>�^����,k�w�x��r0?�[?�q��2��?*>߄ ��=3�+?E�?~[<?�>;%?pK*�;�㽆[>��3>��>ʲ�>�e	>���}v۽�?�}T?���7󜾅ؐ>"\����z�d`=+K>�C5�����[>ԓ<
錾+�Z�v��=�<)W?��>s�)���tc���.Z==E�x?��?./�>zk?��B?.פ<_d����S����Cw=�W?�)i?B�>҇���о����5?��e?��N>�\h�H��<�.��S��#?7�n?j_?D���w}�������o6?��v?s^�ws�����J�V�g=�>�[�>���>��9��k�>�>?�#��G������wY4�%Þ?��@���?��;<��N��=�;?j\�>�O��>ƾ�z������(�q=�"�>���~ev����R,�f�8?ݠ�?���>��������>�o���ʶ?���?�����J�����u��M�h�#>��/>�V���2�;���l6�b�\�Jo��ȾÕ��4�>��@QL8�3G?�j*��ؿ�*ܿl�q��(�㸾�O4?���>`���1�׾�.o�V�V�����/mD�g����>��>�Ͻ$��[z��5�A���j�>i_y�M�>�QI����� �����[<�H�>���>}�z>X��Ԧ��L��?�����ο�ޚ�@T�y)Q?.�?�s�?�??�z�<`Ii���]����,J?/t?��Y?u��[KA�<m�!�j?�^���T`�Ɏ4��HE��U>�"3?�B�>0�-���|=4>���>
h>#/�1�Ŀ�ٶ�������?���?bp����>���?Dt+?kh��7��A[��X�*���)�<A?�2>���'�!�.0=�;Ӓ�i�
?�~0?�|��.���_?ca�\q���-��DȽ✡>.�0���Z������RMe�[ʛ�Gy����?c�?��?����"��0%?v�>V���6Ǿm��<��>!��>�kO>E�[���u>	6�)�:�5!	>��?�j�?��?ڜ���妿z>}�}?���>DA�?��="d�>F�=�ʾ�i��_�">0��=�_�Q�?i\R?_��>%��=��=�¬6�d�F��9O��g�E��+�>�?f?]U?,ʃ>� ������%��1B�9e	��:M�94b�����Z >,�:>�_'>��[��ھ��?q���ؿ�i���p'��44?N��>��?���c�t����q;_?�y�>�6�L,���%��WA�X��?�G�?�?A�׾�L̼�	>��>II�>ս!���ր��A�7>�B?G!��D����o��>X��?�@Zծ?�i��	?���P��^a~�#��7�U��=��7?
1��z>���>��=�nv�ͻ��'�s����>�B�?u{�?��>,�l?c�o���B��1=tM�>��k?�s?�_o�L��B>��?��������K��f?�
@nu@i�^?���׿�*���'���ﭾ�|�=�>Q,V>����h8>=l:�~�z��N��x�I=]��>��">�:i>Kq�>���>Yx>
���*�F#��k_��#���:������I����t���j�������.H����\ʯ��V�v�Լn�'�4G�=WCW?�R?G�o?��?59m�$�><+ �5�0=��,��=�N�>�03?��I?J$?�ȴ=�'���nb�&#��楧��>��S3�>�#8>�b�>X�>Lү>N��O>��S>��q>��=��;=/�D<ve�<+�L>Qx�>���>�H�>6�>���>8���?˶��nh�R���`��O��?��I5�������=�K����>:�?�[c�k���#�ڿ�����2?j����s�����k��)r?`p?p�>�̾�v���U�>�	=����p�=B=�qk�s�3�f�>\�=?�f>�Ku>ס3�Kv8���P������{>�G6?��¯8���u��H��VݾR�M>bӾ>�	G��w�Y�����2i�:�z=�d:?�z?Ŧ��'а���u�X���R>�\>�=��=�M><�b���ƽ�XH�:�.=X�=�^>0�?�+>��=�(�>�k���Q���>$kC>\�/>8g??#%?`������EK���A0�(t>��>�~>p5>��I�F"�=�b�>�S_>f	��M����m�D�+EX>��q���[��Ot�²~=�������=��=pr �L�9�E�=��~?uz��M刿��r����cD?�*?���=�D<~"�����&2��8�?��@�p�?��	��V�k�?�?�?��.��=�}�>ګ>b(ξP�L�{�?�ŽHŢ�̙	��#��M�?�
�?��/�ċ�Il�7>#`%?*�Ӿ�a�>�{�UZ�����)�u���#=|��>�3H?�\��!�O�� >�-u
?3?v_򾶧���ȿ�zv����>��?���?��m��C���@����>���?�bY?�hi>xc۾�OZ�E��>Z�@?RR?��>5�tz'���?l޶?į�?Z#I>_��?�s?��>Q�t�kJ/�";��Ֆ��.�=�b;���>0U>o��QF��ٓ��A��.�j�i���a>��#=D�>Y��oC��`S�=x슽���#Lg��s�>�pq>��I>*z�>�� ?��>Y�>M�=�z��J���⅖�Q�K? ��?%��!8n�t`�<�^�=� _�+4?�=4?��W��Ͼ$٨>3�\?�ŀ?�[?2P�>���D���迿>l��>��<g�K>�,�>�-�>�����7K>��Ծ�MD��e�>�ŗ>b����-ھ9%���ަ��!�>gc!?ۂ�>�ۮ=� ?��#?K�j>�(�>EaE��9��T�E���>���> I?�~?��?�Թ�zZ3�����桿��[�A;N>��x?V?oʕ>[���郝�'nE��BI�m���`��?�tg?�S�<?82�?�??d�A?�)f>��*ؾ�����>��!?����A�C&�e��q�?R?���>Q���ս��ּM���n����?�#\?zE&?r��p'a�,�¾`�<M�#�ԐS�ߙ�;�tC��>�>\���^��=� >:ɰ=T\m�cn6�#�d<�5�=���>q��=�+7�C���0=,?��G�}ۃ���=��r�=xD���>�IL>����^?ll=��{�����x��	U� �? ��?Yk�?`��?�h��$=?�?R	?m"�>�J���}޾5�྿Pw�~x��w�V�>���>z�l���K���ٙ���F��V�Ž�뽝��>�J�>3�?z��>�@>�H?2�A�^���f���羘bg����va0�M�/���.��2ʾ���X���2Ͼ賾�u�>��M�>�0?6$>ᨍ>ѓ�>��=�{�>�s>K�>	Ϟ>�4�=��p>{|B>j��=��G��'S?A����(�Ѻ�yQ���??��c?U�>g���}����� ?~�?Ĝ?�W�>pph���,���?m��>�~���	?�C=y���P��;������%�u���D��>R�Ƚ��9��J��7c�-�?#?���˻Ⱦ�Fƽo���.�n=�M�?��(?��)��Q���o� �W�wS�,���-h�^i����$�ќp�r쏿g]��g$��̡(�<_*=��*?o�?����b���%k� ?�	df>A �>& �>��>�I>�	��1��^�YJ'�)���#Q�>2Y{?��>6�,?tv*?Y�d?�P?�
�>}�>�%��xD%?P��!c�=���>��U?��<?_!?WR?˒B?`�g>g�D��	��y@̾��>�?cX�>�'�>rt�>!��j,3<xI���
&��S~��X����'�����V�.���� �<��=�X?���i�8������k>j�7?���>���>���%�����<	�>��
?�L�>9����sr�<Y��V�>���?��m=��)>� �=�3��$wպ�_�=�¼ѐ=����C;�`/<w��=��=;�o��Յ����:ﾃ;��<�t�>��?���>wD�>�>��� �~��^c�=�Y>�S>>�Gپ5~���$��[�g�`^y>�w�?�z�?��f=��=v��=�|���U�����X���H��<ɣ?�I#?�WT?	��?"�=?�i#?�>U*�PM���^������?kP?_ķ>\��������s�i���?�l?�΂�ztٽ��վ���<�<��>�������-�����?
u> �����P;�?ㄣ?�2���g��ݭ��!��k��dd�>�?��v>H��>`�������-�K��>��>�� ?�?�>E'g?o�?��M?�&�>u���8o��6���u��<_�/>�:3?k?�<�?g�o?/5�>���>Ox��f̾r�(�\����:O��Z��e<��=�޿>8��>
D�>rJ�=�C�D>4������>~p�>�z?*�>��?�ŝ>��;t�G?���>j ���?��C���!��9�HJu?��?�L+?�o=��F�E�Xm�����>�q�?<�?q
*?�S�^D�=ټ������q�j_�>��>N8�>2ɓ=�E=��>���>Z�> �\���l8��P���?o�E?�ؼ=E���@�v�AaǾ�a�K��\+�ڿ󽩽;��Tƾ�J>?�ѽ�LS�C��Hj��Ⱦ�⾾���J"��?���?�>M��K�c=YzS=����^B�G��=�(���<A��`2> X�<9��=����i>v�D<��:l-&�׀˾��}?�<I?�+?�C?�y>�H>/v3����>����:?�V>LhP�u����;�U���b���ؾ�v׾��c��Ɵ��F>�I�3�>�X3>_�=n��<���=as=PΎ=�+S�U=K
�=�'�=:y�=��=\�>iH>�6w?X�������4Q��Z罥�:?�8�>a{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?>ti��d�>L���㎽�q�=K����=2>o��=v�2�T��>��J>���K��D����4�?��@��??�ዿТϿ6a/>�A,>���=�LR���2�I7e��Z�l�V�2�?��=��7ʾ��>\G�=G��Q~ǾM�/=,62>4�E=s���*Z���=]j�O�<tYp=��>��D>��=�ٰ� �=X�W=���=ҭ^>�G�:"�+�C����=��=`�c>yl)>~�>g�?��4?�]_?��>A��[j۾^�¾�Z�>�5=�>��=ފ�>���> �;?�H@?��X?�ɴ>.���r�>�El>?"1��]L���������=���?I�?��>K�)��Z7�uN�cK.����5�?��B?	g?��>������J(�^�'����2�赏=ь^���ļ�
ļ�Sͽ�ء��?�=}��>Z��>{�t>m�p>�_�>��>"��>��>�b;Z�b= ,<�-�:��h�;Up=s'������p��L<3�=?�Ȼ�*���΃2<j��<��
=V�=���>e>���>��=�س��/>Ļ��5�L�l��=�<��T5B�:d�K~�/�d$6�֧B>+�W>�e���*����?%�Y>��?>G}�?�Ou?� >��שվE���le���S�N�=�>=�Aw;�<G`�a�M�hDҾ�>��>��>��Y>�:�'�w�>� >]����$���>+㿽�p�=����ZkB�C���g���%Sj�g����4?7���*��=x׀?حx?,�?n�?�=���w<v>�����쬽�/7�=��_U�B��> "?�.�>��|�B���Ӿ���h�>1�y��O����>'�M�͵Ӿa�>8)��Oɾ+V7�,���F���7�Љ~���>�K?z�?�8K�,�����B�<|���-��Ic�>^nX?/��>>?";?�^�<�پ;�>��9>�v?R�?�%�?�J4>�o*>.~ս�G�>�?1�?Ld�?�3s?�B�����>����C��f۾.$��<�;D�<�>��?j�?�4�>�䇽�p�X|�����t즾\���#W=�A>�>P�b>gE�=��
>)��=V��=Ԯ�>5�:>�w">Y�>]��>8#��w��ȗ7?�>��~>�1?k�>���=�#�D�0=s�<��j������ǽ=)��,�����ʻ�g����>�w¿M�?��>��߾O%�>�1������m>���>g��U�>�<x>�AO>�2�>�~�>� ><�>��<E:Ӿ<{>��Nl!��-C�:yR���Ѿ��z>����P�%���8=��vVI�>c��3^��j�E.���<=�<ý<�F�?����N�k���)����]�?6^�>k6?�Ԍ�눽��>���>�Ǎ>�2������u����a���?���?;c>y�>j�W?g�?Tw1�;�2��jZ���u��!A�
e���`��፿8���}�
�����_?��x?8tA?�N�<)3z>��?@�%�]ӏ�g.�>/�";�	6<=q&�>�(��v�`�k�Ӿ4�þ*P�CF>׍o?�"�?�X?<;V�Z;��bA>��:?�A?5�p?E5?o�*?ۗ�Ą1?�ՙ<��>�?�;?�_+?�?�0>�\k>�T=Lh��w�d��Qb���нQ�"��=br>+��=��;C�a���a=�5=����Ngj��娽�Ύ�H:=w�=g-=k�W=#ä>�ia?wk?M��>��E?��|o?��𽾇�5?�����^p��M����n�4�ھ>�5=ޔi?�&�?H;E?���=\J�m/�Z�.>�2>�\�>]d�>�u�>.�c�Q���'>��>�~>���=�����hl��  �ȥ�**=�Q\>n��>Y|> i���?*>zZ��,v��;g>��R��f����T�,tG��'2���v���>j�J?X�?Ŝ=Q������Z�e��w(?|<?��L?;�?�ʘ=9�ھG9��?J�����W�>,|�<)�
�������v�:��';��s>�ܝ�}Й��>˦�i�~j���'��>�>��+�+<�>K��w�Ê��HII=���=���1
�������I�F?�<>�f������d�־:mR=w(>'��>�齽g�=�J(��'�`>)�>��>d�žmmJ����%@�>��C?��e?�"�?{��/���+\A�4B���f� ���m�%?.�t>�C�>��>7�P�V���(�ˤ{���O�94�>�?�� ���]�$��~'
�"��)Mi>7�	?�=�|?�*Z?���>eq?bB4?t��>V��>©�� ���"?Eqw?L��=0&<��罪�&��XN�(�>�d?��)�=�>+�>@?��5?��T?Ż%?1E�>�om��6@��C�>5-�>�9a������>��4?T>�?��G?Wq�>׀3�\Ҿ6��=��>Ld@>��?/3?(E?��>H��>����*>;U?/|?Kކ?�2�?��=�?�6X=��&?\�x=�i>6e?:4?fN_?u�g?[�@?���>4����O��]���ٽC�=3?=x	Z=`/Y>�	>F+
������>�#ꧽ!���w��~6�������,=�G�=�N�>��s>J����0>-�ľ%8����@>���B_���Ȋ���:���=$t�>��?t��>�S#�M��=둼>?�>���2=(?;�?�?��;��b�1۾O�K�5�>=B?m��=G�l��y��>�u�ah=��m?��^?��W��6��I�b?��]?)h��=�
�þ��b����W�O?=�
?@�G���>��~?Y�q?T��>	�e�:n�)��Db�)�j�Ѷ=^r�>JX�R�d��?�>n�7?�N�>+�b>F%�=^u۾�w��q��i?��?�?���?+*>t�n�V4�[s������]?}t�>�C��W"#?���=Ͼ�ϋ��������|̪��X��@g��
���˪$������ٽ��=i�?3s?�eq?8�_?�� �Nd�4^�����JV�x������E��D��WC��En�G!�:����%����A=`�R��F���?Z�:?sG�	?Ԁg�n�پق�V�X>�Cľ�������f \��������<���T���fۦ���?k�>OTg>&�N?�k���.����%h��P��՚=z��>+ >���>��k>杉=�w����������'�5�s>�d?�7L?z"m?�*���9�i���P�$�G���#j���=P>Gv><��>_=�\��Η� �?��>s�$��S��N���Pp=�,?Xy�>���>��?T�?�n�P�����t��$5��"=�f�>]�l?��>���>|8��Z�ŵ�>b�l?]��>��>ፌ�M\!���{�sxʽ�'�>�>آ�>��o>��,��,\��n��N����9��v�=X�h?������`�V��>RR?��|:S�I<sz�>�Xv�^�!����'�p�>�~?4��=��;>Qyž����{�Y4�� �(?5[?p񄾫]�g�>��?�=e> ��=��z?�d�>�]r�WR��'?��q?[�N?uvF?�-?��>V�������*���=�}i>�TG>|wi=kC�=���A�7��^A��'�;��Q>���,<� ��=aIb<z͆<*gY��H=>�ٿ�B�WR�9S ����n������(K�签ū�������~��p�����GD6� ��l��Ո�R<<�x�?���?�'(�Ŭݾ�ϙ��i[�*��f�u>�B��a�=�Z���)_��Y�����A14����`�6��[���\�;?�Z��e<���(��^��e3-?�_9?��?�Ծ��,���M�i�>B��=���=T�Ͼ(p��s;���Z��5��?k��>�T��拮��u�>ˌ�>���=dea>c�@��n־?	�<O?B?�@�>���mſX����"D�yB�?o�@I}A?��(�����V=���>��	?g�?>WQ1�JG�����vR�>�;�?e��?y�M=E�W�4�	�\�e?E�<~�F�{ݻ[�=�5�=#A=�����J>`V�>|���PA��Gܽ��4>J؅><x"�$���^��]�<q�]>��ս1��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=���w�ʿ�<9�-f$�`M5<��<k]������I*J���}@��i���l���=tv�=YU>5kx>��;>b$W>�{^?&�t?��>Ӹ�<��|�n��51Ͼ,½Fz*��\�*�`��n�z��1^�NO���������73�͐��pY=�D�=I�Q������7"��X���C��(?�:>L!����L�kCL�&ʾU4��5����q��ndž]�2���j��2�?d�??n�IFT���|y���墽esW?�S��v�X@���R>�<l<��[=Fz�>͘�=��Ѿ^�3�B�N��F0?�'?8����h���8>�u �cR�<2$)?�A?,<�>>`%?5%�x�ܽ��m>bC>Gگ>܉�>-m>�����佔/ ?,V?3���D����`�>���.�y�[�T=�V>�=,�˕�-�H>��<����;�Ļ�������<)W?���>��)���*m��d��vm==ѵx?��?5.�>+qk?��B?�y�<c_���S��"�tJw=��W?+i?��>ʵ���
оTs��ߺ5?h�e?V�N>�Uh������.��V��"?��n?�^?���v}�������t6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������0>�"��V�?^��?l2ؾ�1)�����Pr�>D�ܸ�<�1�=k<}��l��4����<:�����������P��e�}>�@�_c�'b�>W�����c�ÿ�ׄ�fjھ�����T<?���>v:y���E��R��<�6C�H�r�	ŕ�@>�>�Q>���Y����{��>;�����<0�>�k	�'{�>�T��ص��W���3<x�>,P�>[��>r�Tý�\��?vu���%ο����ͦ�6�X?�]�?�d�?o?i/<'w���z�+���)G?�Ss?��Y?��#�h�\�\�5�%�~?].��b�Z�4��*5���+=XDA?��.?]o@���9��Z�=�)?d�%�/��"���rS׿IE�f^�?��?t ��ؒ?�Ӟ?]1'?�$��v,�����V��#+�1{?��>-�澻�J���q���p< ?��>�͘���F�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?��>��?�[�=AQ�>�T�==尾z�,�:l#>q��=/�>��?�M?�>�>�@�=9�8��/��YF�xIR��"�V�C���>{�a?r�L?�Hb>�D��dd2�!�ЃͽvG1��r�@i@�MP,�Y�߽g25>�=>E>��D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?�Qo���i�B>��?"������L��f?�
@u@a�^?*x�ܿJ媿���P�����G>=��C>ҏ�����;����z;�30�<w�u>�V�>#�>+��>͝�>=%�>5v^>Ԍ��̓�P��x���!���c��q��;-��멾��@��r����H��մ;�3)���Ͻ�M��cY/���\��>0'i?d�W?��c??�k����C�����>��&�`��>t�ZW?�U? �?D>/cվ�S�:�����x�!ց�;��>_}W>�p?*L?j�>�=:�N>��F>��7>(��=t�=���9!�=�
>f�>��?��>"C>8z>����Bʲ��wk���c�cT/��]�?�DҾ����ύ��1C�V����=��3?H�v=	ǌ�x�ѿֲ����E?����($��5q�!�	>�/?V]=?N�+>����)*�V�j>��:��B��|�=UJ�C�|��01�y27>��=?�6@>w,v>�&1��?���K����r�v>W�1?��ɾ[�	m�%:=���ྨ�(>'��>����A�����s�~�G����=]t=?X�?Iv���A��򏆾@D���&.>��{>��<�R=�i>�|T�u��.�;���M=��=j�>2?A(>1}�=aD�>���ߖU����>�c@>��)>8@?T�#?>�6���Uh��߷6�	�s>�h�>ȼ�>��>�lL�U�=�!�>� a>����v��A��	9���W>yd|���b���q�Cy=D��d7�=�7�=���!>���=H�?����7������m�}?F?�@?��='� =�7(�v����u��U��?q@ �?>K��S��u?@��?����?�=b��>G�>-Hɾ��E��z	?5k���ˢ�ª�r��޸�?O˜?�r�������n����=��(?��þ֌?�z��&��+�������>���>c�n?,#���0e=��̾9�4?��9?����y𐿜���9(K�O�u>M��?7.�?�D���x���<��}C>���?���?�0�>m-=�&"�>̽^&?٭_?�?��-��}���q%?E9�?@�z?aI>�K�?v�s?���>ϸ����4��k��Ĭ���+�=V����5�>�H>{¾�dC��Ԓ����|Jk�+�'�N>��=�U�>��19��ѳ�=LU���訾�`�:ҹ>u\n>�|D>fG�>�� ?��>G�>E=�}���Lv��k��X�K?���?����2n��Q�<���=)�^�s&?�I4?5h[���Ͼ�Ԩ>��\?_?�[?d�>F��<>��7迿�}��]��<��K>�3�>�H�>�"���FK>Q�ԾU4D�jp�>�ϗ>����m?ھ3-���E���A�>�e!?ؓ�>�Ӯ=Q� ?D�#?�nj>|	�>QbE��3����E�1��>��>�U?��~?�?mȹ�'W3����(塿p�[�[N>v�x?�X?���>Ŏ���{��&G�SI�I���К�?@yg?r�{�?V/�?��??ڢA?<�e>[��y�׾�k�����>͹!?a#�x�A�]&�*���?�O?���>���3�ս6$׼���َ���?�\?7,&?���q1a��¾��<2 �;�F�B} <��@��>(S>*���-Z�=�R>�ް=�^m��L6��e<Z!�=�s�>�}�=�Q7��w���<,?�G��ك�c�=A�r��xD�K�>�IL>���ˬ^?�m=�0�{���y��U�R �?��?�j�?���h�8$=?��?�?� �>4I��&}޾����Mw�@}x��w���>���>�l�H�
���S���@F����Ž+�ڽxҚ>��?��?��>Y�==��>Ħ6�$�����B�����?��1M��7s���h�4���E���]�c��d~Ǿ�}�O?�>�<5"/>FO*?�er>)�>%�>�p�� �=���=���>���>��I> >�>S�μX���^?�N��1��:�Q��K?�?%�?<��=�a���1&���.?�ɖ?��?ϑK>��w����;j?�9?Tz]��K�>b,�=YS�=Z7=u����>�_�Wu|�0>ԏ���0�W�dkE�-?�>z��>>o��Pg}�q� =����rPd=�h�?o�(?]�(�FeR���n��V��@R�\��j��Ҡ��c&���q��z��o���#����'���$=��(?u��?����T�"j��N>��m>�9�>�1�>֓�>��J>�v�[U1���]�='�y����v�>a�y?���> �=?�P-?��I?�b?e݄>�J>T��� ?�{X��?�>��>ZI-?��0?�bK?Y'?cfF?���>���b�澭�ʾ�\?��"?h?���>me?S�R�������N�\=�c���@�9�-��*�=��ռ�O��m|���>4�?���8�9y���i>߿7?қ�>�>�����)���w�<�/�>�&
?q�>O ��Qr�R��5�>a|�?�M��a=�'+>�S�=|sw�l\ܺO_�=vȼ���=E�i��:�k~<7Ǿ=W7�=$s�� Q9�\i:Ԟ[;ZЫ<�t�>��?z��>�C�>�?��s� �5��Hg�=Y>�S>�>aEپ,~���$���g�"\y>Sw�?�z�?h�f=U�=ٖ�=�z��3U�����W���M��<��?qJ#?�WT?镒?/�=?dj#?��>*+�UM��~^�������?1C,?,'�>���|�ʾ"꨿�V3��?��?�a�m��wT)�:���jսX�>�l/���~����
�C�����s��cؖ�'��?���?�H;�7���辙����(��v�C?;��>KG�>
G�>��)��g��P�N9>���>V�Q?9�>�S?�Ex?uX?�I=>PH��ث�L̘���= ��=�~@?�n? 3�?�ix?��>��->!I�4��Ĺ�ǐ.��~ýVo��]u�<JƏ>N5�>��>[`�>���=�}��쏶��Ry�� >�ʐ>s��>�ʖ>�g�>YD�>��"<'�G?)��>�Q��<���Ť����z">���u?-��?�+?�=<}���E�"���`�>�l�?e��?B*?��S����=�qּ޶��q��,�>fҹ>$#�>}��=JF=�h>r��>2��>m�U�Vb8�rRM�"�?�F?Ļ=����1�G�ꔺ��g�Y���}�'9��X��<対Q6�=�m���4�?x��L�������>���<���?Ӿ��Q����>3C>y�a>�9�=\ݐ=)���X-��|=2!����=�����z:{�c�/&�0O��޸�I-Ѽ��@�f,{������-v?�JK?2?y�J?��a>2D�=�y��Hv�>�|U�x?b�8>'�����Xw�.��KÏ���ľ�:���l��	���/>}9'<
">5@#>�6+>ςU<��=��<��>��=:=�%�=w.�=�w�==
1>PE%>V�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�%|�l50=w#X��0X��dҾ#��<��^=%w#?�UQ���ǔ>@��>�Q����ľ��<o>��>��|��K6�B�>��ѽVQ<ד<�l>��>!�=�N=]=�'���=��:>�o�� ��<�i5��Nm�|;�����=1>CB�>e4? �*?N�k?���>�����e��@ ̾�r�>w�<���>���=�p>�ŵ>e�6?�P?��K?D�>}S:�h�>���>MH:��mq�����O����8���_i?��c?g�>y���Xvw��z߾���\9@��.?�(C?�?-��>����뿙�@��)�+.+<��R=S=�!p��HL��T�rm�/X��3>s��>�N�>o�>�i>�wG>�]R>��>u�>��<�*E���ٽ��;t�2<��=��%3>F.�=υ�����F/ǽ<�!�{`\��p���s������={u�>�>[!�>���=���j�,>���}L��K�=����D"A��Uf�Ǣ�+1�78��<>��W>�m�� ⑿��?�ne>D >>��?Zu?�4>�4���Ӿl���ji�F�O�d:�=��>W�?�݋:�_��HM���Ӿ���>�&>t��>�*�>߲̾��i����<ܚ�a�	�?R8��(��H��ړ��ỿ�U���<e���=�3?�-~��cf�Q��?LL?�qb?��>��ҽt����>Un!�?����"�T�h��^<�T��>E/Y?>.?����
c��D̾�$����><3I���O������0�������>��>W ��t�о�'3�jj��?�����B�MSr�-�>ƲO?��?�:b�S��oMO�c���녽�p?�xg? !�>=G?D=?UO���k�m��w��=��n?���?�9�?m>���=ŬȽؚ�>+a?Ͽ�?���?=�v?��9��-�>�����D>�r��3�=j>i��=>�>��?s3?�a
?]Ҩ�9����_����X���=L��=���>�~�>44o>�s�=�,=!E�=mD>J��>^ڏ>d>*)�>`��>2���� �[2?� =ҔQ>3L8?m�}>�==�6����k=S����iC����8p$��� �{�r<�<&< }��e�>�:����?vPs>�	�v�?ͣ��=@�<E_�=���=����*� ?U��>>d�>vƨ>�GM>.�c>���=Gݦ����>A��S�:�&�E�J�7�&$��r�>�ؾ�(=J�����<E:��P����Ǿ.`f����j9T��Χ=}�?}0��s��y�,;��Q?�^�>y0?QA���>���=�� ?���>rv뾶���B��AǾ�C�?e�?c;c>��>��W?��?/�1��3��tZ���u�>&A��e���`�t፿������
����I�_?��x?�xA?aG�<W:z>���?;�%��я��&�>/�}&;�&<=R(�>�)��Y�`��ӾƶþB.��QF>�o?�$�?LY?VV�ɪ�*G>p�F?t�N?�?�"?�S9?����i�?�)���;?X�??:?72)?�#?��>8�'>f�=;�*���N�7^���	��X���߽��P=#�>:�<��(�%���L�=j�	=%V%�1���+X���=���=#�=aJD>��>�]?�e�>`p>�!H? �����G�G:ݾ�I+?��=�Z������/����\���> 6l?22�?�6y?A�>Z)5��7��)>�P_>��9>�kK>�X�>�):����B�	=��=z�0>�f�n����K��+߾�Y;�����"1>���>:0|>�����'>}|���0z�:�d>.�Q��̺���S���G���1�C�v��Y�>�K?��?z��=U_��,��eIf�20)?�]<?�NM?��?��=��۾��9���J�K>���>�X�<��� ����#����:��I�:z�s>-2��{p����o>#-�&���h�������W��=��enx>$3,��Ǿ+����>N='>�/���Z#����l����N?e�>;�i���L�ȼ�b�=0,E>���>I��;� ��Q�E�������9>Vj�>�*H>�������0�;��ɛ�>KR?��g?�Ď?[畾2��q�J����۾�鐽)�C?N��>4��>�Q�>W��;�Ŵ�d���x�]f�]��>-z?�)��%E�O�������1����>>�>( �AB?��?��?�� ?`?R��>Fu�>�G;a���X$?�?�W>��=>����i`��k�p��>��9?�U���?�$?�?�?A�?[�?��>�⿾�a���oO>T^&>��B�����l>�P-?�">��V?Jڪ?�ϝ>
ue�H~Ͼx����=xρ>_]?,;?��W?]Ϋ>��>�_���.�À�>ځj?ǆ?/2�?辦=�;
?�g����?��Ǽr,�=�?�1?��!?P�;?t�+?/P?얡���P������b�.D!��8�_K#����=<{��<e>�a9>���=����8��	���l�������C_�>g�s>�	����0>5�ľiL����@>A���gO���݊� �:��ط=���>m�?3��>�U#�l��=k��>?H�>��+5(?;�?�?5Z!;[�b���ھ�K�U�>�	B?��=b�l�т��I�u�h=��m?��^?�W��#����b?>�]? a�=�H�þȾb���Q�O?��
?��G�Nҳ>�~?9�q?��>c�e�t9n�����Hb��k�%�=�z�>�S���d�",�>,�7?:G�>�c>I�=[y۾/�w� s���&?��?��?��?*>��n��1�s���G��$^?-��>�1���#?<���K�Ͼ�T��I4��#�K(��3 ���8���s��p�$�d؃�p#׽���=v�?s?Lq?#�_?�� �P�c��(^�Z ��+kV��,�T$���E��"E�i�C��n�f��J�����AzG=�9i�6�4�	m�?K|6?�,н ��>VM����㾣Q�����>q���F�aRm=X�.��TV����=$?��w1_�:M��'L#?�&�>rla>IU6?��T�p�9�M,��Q����dL=�h�>Ѫ\>ë�>�R�>q= �{��j�󹊾�M�`-v>�sc?�K?z�n?�_�)&1�����i�!��/��J����B>aZ>`��>�W�f��m6&�UV>���r�����u���	��n~=�2?�%�>���>1K�?X�?>z	�d��cOx�|�1�]*�<�E�>�$i?OP�>=�>��Ͻ�� ���>��l?��>��>Ζ��bZ!���{���ʽ?&�>U�>��>`�o>X�,��#\��j��G����9�u�=�h?�����`�C�>�R?>!�:F�G<�|�>�v���!�l��a�'�*�>h|?���=ݝ;>�ž�$�a�{��7��M6)?�?C咾�w*��~>c'"?��>�!�>0�?��>�þ���"�?}�^?�J?�6A?{�>>�=G���&�Ƚ��&��-=\��>[>�l=\��=���a�[�b_�;RE=�=��Ѽ�����Q<����6J<!r�<U14>1�߿v�`������?�Q�"���K���%$�c,���땽p�oϥ��/w�7��'�s=Py��X�����Ծ-��ȵ�?U� @Ί���/e���9�� �ʌ�=�����	.>6\��� �XK���C��As��"���3�r��6�t�A?��7�����բ��4���?�U?!Y�?�����P��5n���>��>h�*>�����塿�1���8���3?`g?�A�+@v�h?�L>�[r>J�?X�z����������?�VS?Q��>{.v�7��ª��>Ӧ�J�?qd@�|A?A�(�p��� V=���>��	?��?>�S1�EI�2 ���U�>�;�?i��?\�M=��W�i�	�Pe?8s<y�F�B�ݻv�=�2�=}E=d����J>�T�>j~��QA��AܽA�4>Bڅ>a|"�g��Ă^�w��<c�]>�սM;��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�+�%�Ͽ��5�t���i �j�[��61��ֽ@�����ӽ(�z�}�U��c�3�.�EL�=��4>�܀>��7>��A>��`?T�X?曥>"�/>6�c��ʮ�W�Ӿ�[=��T�����V��1Z�I���w���l̾e�$,���qϾ���Q>��:�����]8�F�A�)�G�Q-?~{=��!�L�|� 'C� ��R|a�M7�=/7=��~��A~[�>����?<>i?(�B��Q��&�fY�53��3{?��|<��>���b$=��z>3*>5��>Ƿ��]���'�][�v\0?�#?v޽�H?���\,>�I�!=�7*?Pj?l{q<�]�>��$?�S(�X8��[>�U8>ե>ؚ�>dh>(����ܽ��?��T?n+�L᛾b'�>὾i {���@=�V>%5����l�]>�<O���>�	��pH�<^&W?���>��)�����[��i���v== �x?�?��>7vk?\�B?��<�`����S�P�f�w=��W?<&i?�>����8о�v���5?��e?
�N>=Lh������.��T�^ ?V�n?�Y?�u���w}����V���n6?��v?s^�ws�����F�V�d=�>�[�>���>��9��k�>�>?�#��G�� ���xY4�%Þ?��@���?��;< �]��=�;?i\�>��O��>ƾ�z������)�q=�"�>���}ev����	R,�c�8?ݠ�?���>�������u>��}��H�?��?�ے�_#]�ŷ�9�n��N���=�!�=���7b�3T����6��蝾t���վ��ｚ �>�@wun��e�>R��ۤ�v�ƿ�ǉ�
��T4¾_�9?�*�>�+۽��t�U�F��7���)�WN�!�;?��>�N>d���#��+�|�:�:�K���>��
�>�r[��^���Ŝ���~<���>g��>���>IT��!_����?������Ϳw6������X?�'�?�C�?kW?��:<s�u���z���Ӻ{�F?��q?��X?-K�p�X�zf*���j?�]���U`�`�4�LIE��U>�"3?H�>��-�ڦ|=�>��>ki>X!/���Ŀ�ٶ�t���D��?\��?�q�\��>���?rr+?*f�U8��a����*���4�f<A?�2>v���u�!�0=��ؒ�ܺ
?Y}0?My��,�]�_?*�a�M�p���-���ƽ�ۡ> �0��e\�N�����Xe����@y����?N^�?h�?ֵ�� #�f6%?�>e����8Ǿ��<���>�(�>*N>TH_���u>����:�i	>���?�~�?Qj?���� ����U>	�}?]$�>��?o�=�a�>d�=N񰾊-��k#>�"�=��>��?��M?L�>SW�=��8��/�D[F��GR�\$�C�C��>��a?�L?�Kb>&���2��!��uͽ�c1�Q鼪W@�`�,���߽=(5>��=>�>c�D��Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?nQo���i�B>��?"������L��f?�
@u@a�^?*p㿣d���ɾ�����={��=^~E>x	���4=�O==w=�=���=�[r>(Vs>�T�>�G>c�3>��Q>�i��zO��Ǥ���nUM�Ȇ'�<6��0R�Ǒ�������n���_�ž�6��_��@^�����3{���ɽ���=r�U?�R?Zp?^� ?��w��X>����M=_�#���=r�>^n2?o�L?�*?�B�=�|��q�d��Z��]5���̇��w�>�\I>^�>�N�>���>����I>tl?>���>�@>&&=���R�=!O>�S�>ζ�>�d�>>T�>iҠ�~f��冿��5�J����?[Q[���%�d\�����(䃽Ǒ�>�=?R`�C��R̿�ܷ���c?h`��n�'��	�=��<�*?q�g?���>�X��dͽ�Z,>cüm4�=M#>?�{�Q��O�ƾ�ś>u�+?�T>�d>K�6�B���I��3���&Z>R�+?�6˾���Oy���C��L��n�J>�(�>9���d�:Ĕ��;w��?��C�=@�>?��?e6⽳�þ睂���v�x�H>A2>z1�@��=�wd>vC�qfѽ��[��	<�i�=u�=�9?�o,>���=p��>�蘾H`O�O��>��@>M�->r�??8�$?Ee�A���ᝃ��J-��ux>]��>�
�>ơ> uK�=�t�>(�b>,��S�������e?��W>�E��b�^�0�w�N�s=���^�=Q��=�9 �pV=���(=\�~?�|��l䈿��򹶽bjD?6/?3K�=>UG<~�"�� ��M2��m�?}�@k�?��	�&�V��?�?�?���&��=�p�>�۫>�ξ��L��?��Ž�ʢ���	��#��R�?��?t�/��ǋ�l�
>kc%?a�ӾQu�>�p��G���#��6�v��#=���>fI?;��A�N�$B�' ?�b?���XQ��+ɿ�v����>,��?��?tn��=�� ?�=y�>
S�?�kZ?0gh>^ ۾W[����>�@A?g.Q?Ft�>h!���'�?��?��?�I>��?�s?gq�>Ox�'X/��4������v=5�`;�c�>�P>����;lF�lؓ��f��@�j�F���a>֓$=��>WS�y/���6�=bҋ�hI����f�2��>�)q>��I>-U�>X� ?�l�>ޮ�>D�=�w��+܀�D�����K?���?$���2n��N�<蟜=^�^��&?�I4?k[�n�Ͼ�ը>�\?j?�[?!d�>.��F>��I迿7~��	��<��K>4�>�H�>%���FK>��Ծ�4D�bp�>�ϗ>�����?ھ�,���O��]B�>�e!?���>Ӯ=ۙ ?��#?��j>�(�>CaE��9��X�E����>آ�>�H?�~?��?�Թ��Z3�����桿��[�q;N>��x?V?sʕ>b���񃝿�kE�9BI�=���^��?�tg?vS�0?<2�?�??`�A?|)f>և�(ؾl�����>��!?rV���A��V&����;�?�;?s��>hĔ���ӽ�ܼ��I�����?s�[?�&?Q���a���¾�F�<K�$�b�8�%�<ebF�L�>@�>{������=�>��=��l�:�5��Gf<�O�=�'�>�-�=~W7�vn��=,?K�G��ڃ�#�=��r�NxD��>�HL>;���^?l=�q�{�&���x���U�+�?��?ck�?*
��J�h�$=?��?e	?�"�>�I���{޾���PRw�[�x�jw���>L��>Тl���;��������F��K�ŽbF=��
�>�� ?��?q'?X��>���>����@���k���T�d��T�;8Z��_7��������o��ֹA�ً��L*���Nr>�4�=��>� ?6c>�^>�;�>iM<���>Ϋw>�6�>���>Rk�>�d�>��=�6�=.�`jl?����^KE��y��$���%?h�{?�=?/t��s�_���a?���?���?��>�C{��JN�?�� ?����k5�>1v ��z�� vF>݁޾�u�ˡ��L\d��s(> i>�9��7v�vd2�Jv�>���>hzq��[0�lȼf�����n=Q;�?��(?��)���Q��o��W��S�B���0h�4�����$��p�M���^��� ����(�x�*=�*?Q'�?���ݻ��Ǭ���j�L?��!f>���>M�>Ͽ�>�H>��	���1�N�]�9'�r����M�>{F{?��>'�J?�J?�XK?��??�U�=�O>��־Lu
?Bʾ��W>>�H?-P�>@�?��3?s�_?g,�>�p<B�y�(���>��?��>��8?�A)?ks��w����A��щ=�
��B��˥�>Tg�=I;w�H�������=9p? ��y�7��"��Ծu>�_7? ?�>���>xɎ���� =�C�>џ?�r�>k����<p����B�>��?{)���<\o#>��=z�z��-��D�=�8��t��=�c��hE���<���=nĎ=��X:��-;p�.9m�;K��<u�><�?���>�C�>y@��(� �_��e�=�Y>JS>o>�Eپ�}���$��g�g�^y>�w�?�z�?V�f=�=���=�|��yU�����1���?��<�?.J#?XT?W��?r�=?Oj#?۵>
+�dM���^�������?�B?>�>�|�6H�RZ��j	N����>A	M?5@z����a��b	�= �@�K�>��T��|���ϸ���[#'>�q@�6�&�#w�?�4�?4ϗ>bmX��c*�����M���m>?�S�>rZQ>H�'>� >�����/U3�uM$>��>:�f?n3�>J?U?px?�z]?&h4>l�D�3���I�����E=�L�=-�G?J��?�v�?H|s?x}�>�L=>���1˾�s�kG�{��п���F�<	�V>[��>��>x��>V�>�%���н� ���="e1>"E�>�T�>�R�>�^�>n&Y=�yG?�T�>|β���fǏ�t���a�&Y`?�q�?x,)?�#=�����0�߄�!��>�^�?��?R�6?R����=���<�߹��{�����>]��>kј>s�F<�eS=!'u>G��>҃�>7C�!��HD�j$���?�`[?�A�=�W�����aV龷60�v��s0e>J!G�f�����%�?������J��#��j�/)�����Da�����؃�Qy?4g�����=q"�<��<���<N��9C�O>!�M=��=F�T���'>������<9w����>^ :=���=���C˾^�|?B�H?vv+?d�C?�{>3|>��4��ҕ>�ȅ���?9�T>�$R�l/���};����Wg���dؾ�׾j d�L����>H2G��6>DA2>�L�={�<�Z�=O�t=3��=$�ۺ�=g��=�O�=��=C��=��>��>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�'>��>XuS��P4�?b[�iL���Y�
�?͕<�2⾾!�>T6�=��>�ž:6=�u->�uB=gZ!�C�Y���=�|�F�H=/�t=v��>��F>zܺ=�I��̷=�(;=4�=�?W>�h���-��C5��D=��=�Bf>]�>Q��>�_?��0? ?U?���>��$�ln#��ѾT��>1�:g��>E��=9�>��>B�]?K�[?�Td?�Ú>p��=��>ߩ�>7PJ��	��&ʾ�ľ����eT?0�u?��>�@���A�}����P�耹�i�?��'?О?�l�>�I��뿻�;�5����ĽIK��W=U|��oZ��Ž�ѽ� ����=>�Q>h;�>��>&y[>��>	�>�m�>|b�=6��=�'>Bf��ie��%a�ɂ�=��ͼ�C=��+�+�{?�=�<�������B��~�_,�9@�� �=j��>!V>��>r%�=آ��+0>Nޖ��L��ѽ=1��d@B�1d�b~���.�6�V�B>lX>qჽB���y?
Y>Ԣ?>r�?)Eu?�I >�b���վ�O���e�`gS�Ʒ=_�>]=���;�j�`�O�M��bҾ!g�>T�>�"?�<F>�a�C�p���=WUm��+O��F�>�Ӿ�&�<zƾk�����ۿ릿�����ʽ�cF?D핿5�2�?�}?�Y~?i?JO�<l�f�>��5=ڢ���C�1�w�j��C�?��b?�h?��'�!�L���;���	"�>�5N�7QP�����i0���a��ù���>>�����ҾU�3�1��O���B�vs��>�HO?��?��X�zQ��,�O��,�%:f�R?��e?r��>Q2?4?�D���?��x���[�=H_n?���?��?��	>mP>n+���xX>�k&?z�?�"�?��?��'�E��>J�۾�E3>|㖾(��;��8>��=H��=���>·�>7�>�$��D!�sx�;��	��0ٚ=f��=u��>�=�>�GO>y�=1��=��;MV>z7�>{Ԅ>޸�=�m�>�f�>��ߓ
�=�(?�y >���>��2?��>�A@=U���!�=��@���I��F/�s	׽s��[�<С��O+=:���<�>�-ƿP)�?�oW>�/��C?����=��_G>@�H>�Խ>�>�4G>>�>��>��>�N>��>��>\�Ѿ"H>~����&�rH���L�^�Ѿ�[|>>֞���-���}�Q�=�ȫ�����<k�q����<A���p<�ɑ?6ս�m��(��Ľ>?�9�>[e0?���!�L���	>!��>��>f������9��!�Ծ��?��?Qc>Z&�>v�W?��?�t1��3��~Z�M�u��A���d�G�`�/ߍ�m����
�P���6�_?��x?�A?��<�3z>l��?��%��菾�2�>�/�;�nt;=p&�>�����a���Ӿ��þ�r��F>��o?C"�?�j?�CV�t���~��?�3?��?��6?�I?˲��&u?��=��?���>�C?&�#?�t?�]>(��=Z`5���=�L�F���XO���佮>�<� [=MW�=ZE���|9�h>!I��4��oJ������щ9<c+��ٺ�<!��=�~�=�W�>P$�?s��>;�G>�p-?�X��J�[����dR?�Y>A�we�R�,����[�,>�E�?�}�?gB�?�F~>Yꦾ�b�+�i>-�t>��d>�[>V�?$*�����6�@O�<��	>o�=�ĳ���J�v�����h��G�t�_>���>V(|>����D�'>fp��z���d>��Q��ƺ��T�x�G���1�C�v�AW�>�K?!�?���=�X�{���Bf��)?(Q<?&LM?��?�H�=��۾��9�;�J��X���>���<Y��ͻ��� ���:�f"~:V�s>.��Y�M�
f�>m�
�@b0���W��r۾�@�uC�=�Y7��y�>2	$��r4� �̾1�=�*>���v6-�.ş��$��ϵ:?˘
>㍾AR^�@��i���$=g�>��j=هH���P��턾
C>���>!�a>�@���*��T.���+�Fb�>P+K?Lh?�i�?�o���M���`R�*���|��\6N�h�:?z�>z��>�P7=[<<�᫾��F�P�$�T�|�>�c?�)��UQ�I���j׾����>0>� �>�x8=A?^�Q?ϵ�>��Y?
�&?e!?��>M����[��� ?��?X�(>��μV[G��fH��N��)�>�R-?c=ɾ��>��>��
?bE?��;?��)?��<��E�A�V�>�\V>`zM�fך���>+I?��>�	_?G�?��>Z�8�� ������>�|b>'"C?�?O)?���>��>\uþ�%�=��?.�s?XRu?���?KH��5�?6{����>��<Gm�>Ž?��>p�6?'�h?�??�J?-�-��?�׻&�u!1<�56��%�;�
(>�q��w�m1~=Q��=��{�������$�Н�� ��<A u=[a�>�s>}	�� �0>(�ľ)O��Y�@>�F���H��V؊�^�:��ٷ=���>��?㬕>�L#�ݽ�=఼>�F�>���5(?�?G?�V#;)�b�+�ھ�K�Y
�>�B?J��=#�l�s����u���g=1�m?U�^?u�W�� ���b?%B^?j��ʅ=�G�þ�Zb����<�O?�
?΢E��C�>	�~?)�q?�$�>�d��3n�?��T�b��Wm��ȷ=by�>O���d�3a�>�7?��>�Xd>�h�={=۾Q�w�h����U?XȌ?ѯ?��?n�)>P�n�r࿚���+��p�a?r��>p���8�?�������N����۾�z��{ښ�����ꩾ�w �t���s���*�=�`?Ԥn?ro?�e`?	3���c�q�_������Z������PB�$�@�6H�(�j����n���������<��^��VE��Q�?<0?�\\�A��>?�対�ԫ���T>"����W>�	\>4����Z;4r=�ʂ��H���E���\ ?���>x�>�EB?oQ�X�7�
6���5��K��F>�p�>U�|>-�>{���l6��i"�w�žw�㽏!N���y>ce?ţL?��l?��5��e��TK!���亾])b>e>�M�>$�^����ْ��P?�Ąr�z7�믍��c�^sZ=/�-?݁>���>���?ot?̚��/�����6|8��a�<��>ǭh?g��>O�>P�ӽ�~����>2�l?���>��>���8Z!�R�{�Ԙʽ�%�>0ܭ>ߴ�>��o>I�,��"\��j��;���n9��i�=ɧh?d�����`�v�>R?	6�:�G<;y�>�v�k�!����%�'�y�>�~? ��=(�;>@}ž5#��{�B8��MH)?�?]V����)��b~>��!?���>���>z��?���>�����*���?G�]?�qJ?*�@?t{�>?&=�����#ɽ2['�k[6=V�>�K]>�<r==h�=:��+_��@#���2=U��=���m��m�;11׼���;�a�<�q7>��ֿbN�%�߾S=��Gؾ��ƾΊ�1�ս(�پR����/̾��þ?ƾ� c�/��<a��󜇾�/̾�A��.�?��?��e����+똿=�c������>8�g�y=~d��|굽0*���
Ծo+��s�/��e>�Ҧq���p�Z�'?�^����ǿ����=tݾc�?.~ ?6�y?=�� �"�C�8��g">���<Z+��:꾟���n�ο����%k^?L�>�ﾩ���;��>��>F�W>�"p>@�������7]�<��?s-?��>4s�Wɿ]l��@N�<��?��@eA?��(�[@�V�X=�>�	?�C?>�1���� ɰ�.�>��?F�?�K=Y�W�A<�E�e?0�<j�F��&Ի��=덣=-=$����J>`!�>�|�#�@�Lݽ� 5>��>i7%�����^�B��<��]>�Zս�J��'Մ?�z\�sf�r�/��T��UU>��T?�*�>;�=̲,?�6H�[}Ͽ��\�}*a?�0�?��?^�(?�ڿ�ٚ>s�ܾl�M?*D6?��>od&���t�ч�=9�B������&V���=���>ƅ>��,�����O��M�����=�Q��ʿ�?�w�-��x=&�=.4����^�t�8� D��Ŧ�$Ь�vb���厽]f�>x�><b>��>��>�T?!jd?�A�>���=f�S���w¾��Ͻ���2*⽈Ҟ��G�j�����辑�����#�8�$�U ;�n�˾�d"���G>CQD�bv��X��tA���O�U?�,�����X��Z�;b�	�k$�����=ܥ����羝A_��c��?=�i?OBs���Q���K�s�C���Z?��-ZԾ�D��M�t>|�>M�J;���>��|=Jd���~�+h���.?��?��������\@>�н���=?�#�>z9g=��>E�?�JC���۽-�i>�>>4}�>���>M3>�A�����t?|X?�9�ŏ�
Җ>��ʾ�N��ʫ<̵�=S^�� <*��>�>h�e��D9���ƽ�"=K�V?���>��)��5��J�������R=�2v?R�?�g�>J�j?��A?�Jl<=��O�Q���	�xώ=2$W?(�h?�?>H#��u�̾3��I5?� e?�nQ>Q�m���꾃`/�I�ػ?�*o?�'? �ɼ�}�%�����K6?��v?,o^�Jr�������V�>�>!X�>Z��>��9��p�>�>?(#�^E��x���PT4��Þ?
�@e��?,9<<�%����=�8?yQ�>C�O�|<ƾ�]��E����fq=;&�>#���%ev���VZ,���8?C��?ِ�>咂���.;%>�|�����?���?w���ƽ0�v���Y:���G�?1>��â�=����6�'��$���m�B�>ڙ@���I|>��R��濺E׿`?���9۾���9�C?]?Uj���贾$VG��t`��OC��bD��O��JC�>4�>w����̑�Y�{�U-;�y���X��>����>��S������D��>�.<E��>Y��>R��>���߽����?s����6ο&���A����X?�P�?�X�?aU?�d;<�u�"{��x"��G?b|s?%�Y?ތ!���\��,6��j?>_��9U`�Ў4�~HE��U>�"3?�B�>[�-���|=>��><g>�#/���Ŀ�ٶ�O���W��?̉�?�o����>o��?�s+?Ei��7��j[����*���+��<A?�2>ь��[�!��0=��Ғ���
?-~0?{�.�H�_?ۚa�8�p�_�-���ƽ�ۡ>��0��f\��N�����SXe����xAy����?"^�?H�?��� #�n6%?��>{���58Ǿ�<���>�(�>U*N>�L_���u>����:�|j	>���?�~�?�i?땏�����T>��}?�#�>��?�t�=%b�>Wc�=a��,�nm#>�&�=�>���?�M?�K�>�U�=��8��/�Y[F��GR�$���C���>J�a?L?�Gb>���y#2��!��sͽ�`1��E鼺V@�ǉ,���߽L)5>��=>>��D�@Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Ua~����7�b��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B�y�1=7M�>Μk?�s?`Qo���j�B>��?"������L��f?�
@u@a�^?*�ؿ�͡�k�Ѿ������=�W�=,bG>��Խ��M=�$���^ƹ2醽N�J=,>�>�w>[ >�U%>�T>f>�h���b'�S�������fG�-�[����F�y^��_��+���þ��D�A�B�Ͻ���!�1�q�i�)]����=��U?�R?��o?,H ?�J���>����*o=�O'���=��>��1?\�K?$R*?��=�w��{Nd�N9��:̦�Hg����>/J>�`�>tc�>0��>.7;oM>��B>Ҵ>�S�=͗%=��"�h*=�O>�4�>�y�>�3�>��>��>i�����z���^�z�:ob�a+�?q%��R$<������~>Ø<1��>�|T?<HH�>����_ӿWd��I.4?}	¾z�
���>�����\�>��?9��>{��<��[����=�R$=�Q4�ŧ>���<@}��V����N�>ɋ?���>O�x>��9��v8�]	Z�a�����>��9?�����-�pz�%�6��{Ѿ��f>@��>�����;���]h|�F�c�E5�=��9?�A�>����+��@���R����I>27>��=&�=�<>�Jy��ý�eS��A��6>��t>�??�n0>�a�=Q��>�땾��C��>�a7>}�0>i�A?��%?'�K�Dޔ������]��>���>l�>�>>�fI�İ�=r��>�aW>h��Vt�S��	�A�b�G>�[�2Yc���v��h=-���=�h�=a��5=�*d8=�~?�]�������뾍Q��w4D?�K?;!�=�	M<�z"����S���H��?�@�x�?ʄ	�ԠV�Γ?�?^r����=���>���>M�;�L��u?�$ýc㢾>�	���"�R=�?�?�91�����}l�=4>�%?q#ӾLh�>tx��Z�������u���#=O��>�8H?�V����O�h>��v
?�?�^�ީ����ȿ2|v����>V�?���?b�m��A���@����>:��?�gY?zoi>�g۾6`Z����>Ի@?�R?�>�9�s�'���?�޶?ԯ�?�M>	n�?5>t?���>���/D5�$�����ܴ]=�����K�>�Z>9���a�H�z��������j��<�~�D>�� =j�>�3���¾Q��=YIy��ף�� ����>��[>DP>-8�>/��>��> �>�p�=�	j��)��Cr���-L?:��?����Gn�0��<�d�=��]���?db3?ݿB�f�Ѿ8��>k�\?��?qh[?y5�> �)?��*ӿ�MԳ�d�<��K>���>RF�>fN��
vK>��Ѿ�C��͈>�q�>#ԗ��uپ:������
�>�] ?XC�>�P�=�� ?Ĝ#?��j>�(�>�`E��9����E����>	��>H?;�~?�?�Թ��Z3�����桿��[��:N>��x?�U?�˕>e���ꃝ�)fE��HI�����Λ�?/tg?�W�Z?;2�?W�??-�A?'*f>'���ؾ,����>��!?dF�W�A�gy&�����?�?��>-�����ӽ��ڼ>��>���P�?6\?�&?ӑ�3>a��2þ���<�*$��JB��e�;F�G���>:>2P��!�=�9>^�=#�l�36���p<�=��>u��=��6��䎽a0,?iA>� ��%��=Dr�VD�-N�>�K>���<�^?.�<���{����Q����S���?D��?;S�?T/��ch��<?��?�-?�/�>�Ԯ���ݾ���x��*y�����>��>��H��h��{������>J��<Ľ����y�>�v�>I�?�>�7>�~�>��.��& �u:��^�AU���'�w�>�K�4�����xҾM�X�.����ɾ�`w���>�ڼ���>QU ?M�Q>�>�M?D�ͼ��>~mH>m��>UY�>��>[/[>k5>�Ᵹ7:ɽ��V?RF���W/�ZZ输7Ѿѓ6?�ng?�?_��~��z��8�(?��?��?�s�>�
f��\-�t[�>Q��>>���
?�ڻ=4I��_ =Qڻ�=�:��; _���+q>	J����2�f%I���k�� ?�?? #~��թ���u���jo=JR�?'�(?�)�f�Q���o�R�W��S������g��V��s�$�k�p�=菿�[��u'��Ő(�1)=]�*?�$�?l��a��	���/k��(?���e>%��>��>��>��I>}�	���1�H�]�C'�Y�����>={?Y��>��)?�$$?�4M?�W?�:�>���>�;���e�>��Zv�>t�>Qb#?�8?��?k)$?-q3?֡>;.5=MO���S����?�=?<�?��
??`���Af̽�b�c�e�P�d��>Y>JAa�����GP�`>q��EK>�Q?+��Ӭ8�Y���^=k>6�7?՛�>E��>���c#���<H��>"�
?/N�>� ��kr��O��g�>5��?&��s=,�)>��=w�����ݺ2�=����ܐ=�r��Er;�fl <��=@ؔ=��t�w�j���:g	�; ��<u�>%�?���>tC�>%?���� �����a�=�Y>�S>">�Fپ�}��_$��)�g�a_y>�w�?�z�?��f=a�= ��=g|��)T�����/���m��<�?-I#?^WT?���?��=?�i#?�>+�*M��m^��:��Ѯ?�Z??}0�>@��A�ľ�d���Bq�t��>�Hf?iJ��_��;S#�0��=r�P=���>�W$��C���좿`
޾�$�<�$z��F�?\l�?*��>	�f�l$������񾤿@?�6?k��>^�|>��#������J���>@�?,�_?#X�>o�U?YOz?��W?/@>�7C�ok���씿Ӹ"<': =�N?�#|?���?�Y`?櫼>�rH>jP��$���#����޽���=�$=� h>��>7��>43�>y�.>����R��j:���N�=7�>Q��>��>S��>0l>��=�B?���>jx�������P��(�K��+o�y�T?[U�?i8?�j>�-�%B0��?���>qJ�?��?�6?���t�=xO*<k7������I��>�ī>�.�>�Vt=�c�F�d>��>��>!����������ӽl*?�%2?B�=)ƿ�q�UHs����S�Y<hÑ���d�����\��K�=Ȋ��������h?\�F}��C{��(�������y�/8�>eވ=>U�=)��=ŗ�<{¼4��<I=�<�g=��l�y�v<�9���л�E��b�ߺk=_<rfL=���%�˾Վ}?$<I?��+?L�C?ְy>n4>��3�Z��>����pA?pV>��P�-���9�;�.���-"��e�ؾ�v׾��c�g͟�SG>/GI���>�73>Y<�=ma�<o�=�@s=�Ǝ=t�P�H:=�&�=&U�=i�=���=��>�S>�6w?R���	����4Q��Z罣�:?�8�>E{�=|�ƾv@?��>>�2������}b��-?���?�T�?C�?&ti��d�>@���㎽sq�=����=2>���=t�2�?��>��J>���K��v���~4�?��@��??�ዿʢϿAa/>��	>�LM>�M��G�?!z�t�ټ��T��"?�oY�����;�e>�>67�L��$>�=��=���=Fґ�hkJ�xv >9�m�9��=�
��g>��>�K8=�; ��u
>�=��>l�>�2Q�(=N�����#>�5*=Fgj>!��=F��>���>��?a\?�4�>�}�p����þ��?~=���>N������>i�L>���>�Q?ܶc?��>__�<�;�>���>]�j�;����Њ1�,��=�YW?AC?$��>u�c>���g=����_^b>��?�+/?�� ?���>1����u�Y�?gE�V�c���p7�&��;��vM�|���F�&M��ST>RE�>��|>̓�>�>>��>��>0�T>L R>�㊼^%ڽgd�=����m�=ɛh=B>�>s����3���G����	�};Θ*��=��}<1�=�/�=���>\s>���>�@�=`ó��0>_���|L��
�="����B���d�E0~�o/��S7���@>��W>�4��d���?�fZ>��@>�k�?1�u?8O!>Eq���Ӿm��|+f�`�T����=]&>܏9�	z:�2`�g=N��#Ҿ���>��>X��>]�>E��$�j��(u=�q���;�^��>C�%���>�b��-�V���ƿ��ĭr���=��%?��&S���(g?� S?��?�L?/_�=�������>��������:�T��񾆟��I�%?��O?LK�>�L%�¯9�
_̾F���ў�>g�K���O����h0����\���{g�>���bо��3�Jt���s��M�B�h(q�k��> O?��?|�]����pO�����/���??��g?m*�>�B?2o?uD������%���6�=q�n?���?b��?6m	>lU�=��T�/��>GR?�t�?-��?�v?(t��LI�>f��9��_>��%�Uo^>��0>�\Ӽ�h>D�?��?ul ?|uu�֏����j�
��JM�Ӱ=�.=R��>��}>j,B>�%>���=��Y���@>�ƅ>��#>�T>��>+Ł>}R�����B?]�I>~�>>x2?���>�_N>�o�=�*�;��[:��G��C��؊�����+M���{ѽg���@nW�p��>w�ÿ�5�?P�>�N%��b?KO��l/<:��=�W�>d�m����>���>y2�>��>۽>6�E>���>���	7Ӿ��>N���d!��3C�R�>�Ѿӕz>���e&�:��A?��7I��`��V[��
j��,��/>=�`V�<ZE�?X���M�k���)�������?kR�>�6?�ڌ�r.����>(��>�>/K������ƍ��h��? ��?�>c>��>��W?��?p�1��3��vZ�'�u�*!A��e�o�`�Q፿������
�H��%�_?��x?wxA?�*�<6z>۠�?��%�gЏ��,�>/�#%;�&F<=y,�>�����`��Ӿ��þ>�JF>��o?Y%�?�[?)GV��<���=��&?��??/Co?�5?�^?�=�?)�5Z�>�\�>�p-?�uO?C��>��q>o�>�;�=�)�>�z̽��v�/�u�S�����<�˪���x=D�=���;A��מ<�6��>��_L���ߤ<�A�=O������=�->Р�>d3?֔�>��>$�I?�>佳���_��A�B?%@�>`4@������E8�U(� й=yΈ?>��?S]Z?W7@>�%K��d��5�<>�E�>.�>`Z�>�x�>�GR�x�s�\�">dM�.�>�@>O�=����
��S�ϼ���'/>C��>^5|>�獽��'>[g��
Dz�fzd>��Q�]����T���G���1��/v��@�>}�K?S�?���=D+龒<��oAf�)?�m<?�IM?��?�C�=��۾h�9���J����-Ο>�q�<c��J����'��k�:��~�:�s>
���aþ)�W>p�
�z��Eg�d�<�O�wbb=-;���=J��ԝ�@���)iA= )>�jھ�{������ি$�F?ؐ�=䁙�U�>��פ�͙>���>ܚ�>i.o;҂6��eN�񴾾Bt=,��>��4>1/��v��"�D�ވ����>��@?2#]?>|~?s-���Gm��@I�����L߶�S�-��F?.\�>���>�>�	�<֝��U��Z$`�]�A�K��>q�?�~��@��흾���/#�,��>B�
?K�=	?H�P?<?�HV?4�?�^?=�>+�������u%?܁�?�,~;��J�<����r ����>'�)?����_(q>ß?���>��>vv'?�6?�mf>I_������>�x�>ac��²��,�>17Q?���>�*d?�J�?��Y>�nJ�-�澅C
�|Q$=�6>��T?b�2?�\�>��>R�>�s���L�<E_�>��<?vۉ?4,�?h�ļ��?"��=�,?@\�<;o�<�J�>�C?|�R?���?N	Z?��0?��<I"��Y@��E*Ͻi_=����?�H�=#@;�%=0I�=n�=o����(��Q�9<�[�@���dP>߭=_�>t�s>����1>��ľ�E����@>���WF���ߊ���:�v�=���> �?g��>X#���={��>�G�>Y���3(?��?b?2E!;y�b�]�ھ]�K���>�B?���=��l�������u�e�g=�m?I�^?c�W��"���b?��^?48��A�>������b���,�Q?S�
?^%K�7�>�]?Tr?�_�>��Z���k�]���ۏa��ps�X�=�ћ>%��?b����>�W7?���>��k>���=h:ι�s�\F����?���?��?Ɋ?bA>0zl���߿��������^�^?WT�>�ӡ�4"?>��ݡξu���
*����̩��^���*������r�&�E����ͽ͘�=��?Js?��o?��^?AH��a��^�:W����V���Ob�qD�dD���E��l�=�����Y<���$=]Ex��+`�M~�?|�?�G=��>����2�߾�����>������慱�h壽�,���l�����"ҽ��T�s�?�[�>{�>y0?�_����'�5���J�-��!��<�5�>s�>��>"�{��_���T���b;��l��U��0�~>e?��D?\g?���\�%��Ă���"����ܗ��UD>��5>Z�{>��n����W-�C{8��^u����� �����7d=ս3?Ā}>�(�>Ζ?��>~t㾞������h
0�0�4=;h�>4rk?��>Gz>S���E����>s�l?��>%�>�����N!�)�{�l�ʽ|(�>�ƭ>���>��o>ŭ,�� \��b��t|���9�<�=F�h?�~��h�`�څ>R?���:��I<f��>��v���!�����'���>�z?���=��;>]�ž?�H�{��.��Me)?�}?����e)�ʍ�>z�#?���>���>Xx�?�t�>!�þ��\X?�![? �H?laA?��>��/=?����ǽx�&�V6=Tl�>
g\>�]=���=$g�� ^��N��$_=�R�=&���a��Yq^<�i���;vi2=S�4>�޿ʟG�U%վ�!�������p���輽?*�������¾s���t����g�)�s�������S�����l�A�jo�?�.�?�Y��
��l�����e����ހ�>�9��U޽\���V�w�Q[þD׆�3�%���a����������'?\�����ǿ!����`ܾ� ?; ?��y?���ɧ"�Q�8�ê >�?�<d���X�6���)�ο����N�^?¿�>+��#��"�><p�>]X>��q>E��������<A�?�c-?���>�q���ɿ~���:~�<���?J�@cvA?�(�٨쾩mV=G��>Ό	?Z�?> q1��8�8$���I�>�:�?���?y�L=a�W�Ce	�ale?C��;��F��2ܻ�E�=C̤=q�=�����J>8h�>����@�UNܽ*f4>Ʌ>�"����^@^��a�<d�]>��ս�唽6Մ?&{\��f���/��T���T>��T?+�>i:�=��,?T7H�]}Ͽ��\��*a?�0�?��?�(?0ۿ��ؚ>��ܾ��M?]D6?���>�d&��t�+��=96�鏤�X���&V�?��=\��>��>�,�ދ�w�O��I��`��=���ƿY�
���b=�E<Z6��p���֞�Ln��z����g��qD�H2ۻ!�=e>S��>��>f��>��[?fst?Mߢ>.�x=�u��Y�{�͎⾩.�<#6��L�5�KC��[佣~��$=ܾ��ľn��_&�4�&��о'���qM>��S�Q8������$�U���j�>w6?|>�oz���l�L��=��l�����m ��QF]���޾��4��/L�yo�?��<?1�o�.;�e�Qd�=1⛽I��?kMǼ�8�:/��;LM>w�N>���<l�?]�>M���& �>�Y�+�-?za*?�Ժ�,�`����>W�=�Ԅ=�~ ?±?�����>g	?V���ѽ�͆>KMU>���>���>��y>�m��g
�42?�Uc?����3���M>s�Ⱦk���,�=UX�>$�żJ�>s��>Z?�=Z���п�Y63����;J(W?.��>�)���[��r��&u==��x?��?:+�>Wxk?p�B?���<`h��%�S����w=S�W?!*i?��>Ǌ���о�}��1�5?ןe?I�N>1ch�����.��P��%?��n?@a?2H��2w}����6��Fm6?��v?s^�ws�����K�V�h=�>�[�>���>��9��k�>�>?�#��G������xY4�%Þ?��@���?�;<��T��=�;?k\�>��O��>ƾ {������+�q=�"�>���}ev����R,�e�8?ܠ�?���>���������=R��=j�?��o?kc�\&N�k�FZ��(�ת�=x(�=2��<���:	�� D�`ľ���r�o��qw�  �>%R@P�R��ݵ>����Կ�ȿ3o�Zʾ�wľ�?�ƪ>�h���˾RQ��>�T�:��M���Ǿ}�>�x>����Y���{� I;��Ĥ�z��>���P��>XT������䞾��7<=�>|t�>J%�>�����/�����?���� ο���������X?LW�?�z�?46?*�4<=�u�:L{�����G?Pes? Z?H�%�]�Y�:�"�j?�_��qU`��4�mHE��U>�"3?�B�>T�-�ײ|=�>���>g>�#/�y�Ŀ�ٶ�@���X��?��?�o���>q��?ts+?�i�8���[����*���+��<A?�2>���L�!�F0=�SҒ�ü
?V~0?{�d.�k�_?�a�h�p���-���ƽyۡ>��0�Ee\�K�����Xe����H@y����?L^�?\�?j��� #�,6%?�>�����8Ǿ�	�<[��>�(�>�*N>CH_�(�u>w���:�bh	>���?�~�?j?�����V>��}?�5�>M�?\��=(0�>�&�=�߯��K�"6!>� �=��I�/^?!�M?���>���=�7��y.��F��qR�2��1rC�n��>��a?�L?�%a>?&���@*��c!�ǽ</�Z��m	B���(���޽��6>]�;>9>M%B���Ѿ��?Mp�9�ؿ j�� p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>D�Խ����\�����7>1�B?Y��D��u�o�y�>���?
�@�ծ?ji�X	? ��P��Oa~�?���7����=��7?�0� �z>���>��=ov�⻪�-�s�%��>�B�?�{�?E��>��l?��o�@�B���1=�L�>��k?�s?�Po�i�R�B>r�?/�����L��f?��
@qu@=�^?�翱�������ʾ�9����=\�}>�X;�o�=��==-W9�a����.)��#�=��r>�J�>@?W�?!�>������͇��D����O��@�����6����od��r�����M0������I��LZ�=#��;9�Ƚ��M5 >�X?��K?Fi?���>c��iA�=�C=,bU��)y=gM�>J$,?�>?��'?ᘸ=:��>=i��|�륢�AV���_�>�-_>MD�>!��>��>�kF��{>�>I>a,\>E�=��~=!_л��=�/>�j�>�G�>*&�>�3�>���>d��]ĩ���Y���p���U�iC�?4B��4�c��\�k���Y^�8��=7�v?�*1>A����毿_ȵ�kI?�VǾ���� �=��9�?�=�?`�>��������̙]>�d��^IϽ���>�d���'�4�#��x�>���>��c>^Ft>r�3��t8��aP�Fد�0{>��5?U���E�9��v��I� fݾ�SL>�Ѿ>�u�@��Ȗ��/��ug��2y=W�9?��?���4���I�t��n���P>�]>/�=f�=��N>��W���Ͻ �H��/=��=�C_>v�?�w.>�Z�=�F�>+�� �I�禧>��8>H�2>Ѓ>?�3$?����z��_���lS'��Ku>��>�>8�>��J��=���>�Ui>XI�V/��~S��@��W>��v���^�����ʀ=���IT�=t�=���W6�0�%=��~?�h����e��^��&FD?�*?f�=]�J<J�"�t馿�B��>�?��@�d�?�_	�Q�V�j�?��?�����=�l�>D�>^Cξ�+M�*�?טŽ�4��1	�z�"��'�?���?�r*��틿l��>�E%??~Ӿ?h�>�x�eZ�����h�u�&�#=,��>�8H?�V��E�O��>��v
?�?{^�⩤���ȿ3|v����>G�?���?c�m�nA���@�ׂ�>9��?pgY?Foi>og۾�_Z����>׻@?�R?��>�9�l�'�s�?�޶?߯�?�8c>+q�?/�f?^�>3��u�2�'̷�������_�b��"w�>L�|>� Ծ;�J�B���, l�;_��$�7*>w=�v�>WK�[S�����=Z�'<�}��F�w��X�>3(X=��=ɳ�>���>���>1�>��=��<K������5L?W��?�l���m��<Jڛ=g6^���?J4?�L��uϾԨ>��\?���?	;[?݈�>�+�����⿿l��Qa�<~gK>#��>1��>�Ί��IN>�Ծ�XE����>깗>�i��,پ� ��ɽ�Ʊ�>ph!?��>�=�� ?V�#?³j>UB�>�XE��,����E���>׌�>E,?��~?�?5ƹ��Z3�����]ޡ�%�[�9%N>y�x?UT?*�>�������iE�GI��㒽���?Ddg?Q
��?�0�?�s??��A?�e>+J��׾�^��݀>[�!?����A���%��y��	?�d?AB�>u㊽ƽ۽sy�ʱ����u�?�w[?��&?��a�K�����<���Y���ȡ�;� �\>��>����W�=5�>�W�=�0r�z6�w5}<�Ǻ=ٯ�>���=�1��ꉽ0=,?��G��ۃ���=��r�4xD���>�IL>����^?gl=��{�����x��	U�� �?���?Zk�?-��;�h��$=?�?S	?j"�>K���}޾5���Pw�~x�~w�r�>���>+�l���J���ؙ���F��X�Ž_w���>3��>�?g��>�X>+Y�>Ö���M �������]x]�.P���6���(�����Ԥ�qT�C���8����x�HĖ>�儽e��>S?:�q>�>0��>�=��2��>
�Y>J�>���>ǝM>U$>y�>�G<�ҽ�cR?r�����'����$��	B?jad?��>��g�@���k��a?ː�?�t�?]�v>,Kh�^F+�e?p��>���nA
?�:=x�l��<����G��8ۆ�g&�;�>f�ֽ)2:�.�L���d�J�	?M?�����k̾��ֽG��q9b=��?�Q?I���5N�T\q���P�E�S�e�I!m��5��&�&��eo��͎�i����M����(����ǟ+?��?ˢ
�#W辧���o�p��K��rh>M��>_�w>;%�>ns�>���-�$���[����3Nc���>wr?�c�>�)??�E9?��o?X�?i,�>O��>�
�a6�>!M&��D�>�y�>��$?2b?U�6?�%?rk?�Nu>ȩ��쾇�ؾ�4(?�Q?ZΛ>.L�>>Y?ϭ̾X��V5�={��=ُ���=��$>�6]=��ͽ�����=ܡ<�Y?�f�h�8�O���_k>��7?��>���> 񏾡0��+3�<P��>�
?G/�>���Qjr�<S�kW�>5��?����m=�)>���=}ք�3ٺ:I�= ���~ِ=W��~;�Wu<"�=�=�=;p� r�����:睑;z��<0�>H�?�e�>G.�>���s� �ؙ��=�=�mY>��R>(�>:dپVx��=����g��y>�u�?x�?��g=���=_�=�W���5��0��������<m�?�'#?�ST?���?��=?om#?�$>���M��f\��Т��?VF?kl�= �1�3��c�m{��?;�M?�{�k3>C�Ͼo���Ҵ>��?��9��G���!$��ƾ���Iw�o�?��v?�[>e
Y�Xi����t�2>��#}?�<>�:.<�-�>��0���PAQ���R>;2�>F�H?Sۼ>�Q?�t?c�V?3�K>�U/�?���w*��8񫻍)�=�:?�E�?�?j*j?[��>e&>��*�4��
���T��o�ٽ�����`�="^>���>~�>���>B<> �ڽ1��Һ=��|�=�[>M��>�ٚ>`�><s>�'=�G?8�>��¾KN��坾@�l��K���q?���?r&?Q�<�-��HD��������>�?dh�?��%?�C�Dv�=��ļd����Fz��g�>��>Aw�>��=�/g=��(>bG�>IL�>�l�%���}5��t4���?�~I? ��={}��J�Om���jӾ��
> ��2���j��I���o-�=!m�qc]�L)��)�^�['��! �w���X�Ҿr���s�?26�=��=�J�=���=��87m���=�1�<���=.bF�9�=�c�=�Z=ş�qw�:���:!��=sF�=}ɾڇ|?1I?��-?�A?��~>a�>K^����>�����?_�P>@+Q�������2��<�����g־&�Ծ��c��៾>�	>�'�?W>�2>{�=F�<}+�=�d=;Ɋ=��n�]�.=<�=b��=^N�=|�=�\>�\>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�8>X
>�_Q��0�%Z�*�`�ia��?'$:�fZϾKr�>H`�=��޾�JǾ�W#=4�8>�:^=#!���[����=0�p��j3=v�p=�>�>:RL>3�=Sⷽ۶�=�a@=�/�='M>�:o�3�O>
���2=���=�]a>rQ(>AU�>��?(�'?�Bw?37�>^.�Х��+���>J#v��.�>�\>��U>��z>�K*?A?<�1?z��>Y��=���>��>/'@����ꩲ�-��;�=î�?��a?y�s>�r�;"�z�'��=�L���?��_?{J�>��>�U����9Y&���.�#���p4��+=�mr��QU�E���Hm�:�㽨�=�p�>���>��>9Ty>�9>��N>��>��>�6�<sp�=(ጻ���<� �����=.�����<�vż疉�u&�8�+�+���`�;���;��]<1��;��=k��>
=>���>ݍ�=]���A/>&�����L����=JG���+B�Y4d�KI~�/��U6�:�B>�8X>�~���3����?n�Y>!m?>f��?rAu?��>� �
�վ�Q��JEe�|US��͸=_�>��<��z;�9Z`�(�M��{Ҿ|3�>�\�=V*�>i�(>�>�NM_���=����J=�Y�!?8�����H��B��R*�$o��aH��*7l�C��<H�A? 悿�?��T�?�&*?�R�?df?�r�t*���Q�>2�1�̈́d���þ�#��Fֽ�� ?3�	?���>�.��4K۾�J̾5���ҷ>�TI�(�O������0�����ķ�Y��>�����о�!3�.e�������B��Pr��>.�O?U�?,&b�V��$TO�+���>��ij?og?��>J?�=?�����h��k���g�=��n?L��?99�?�
>@7�=O�H�/�>�Y?�ې?̄�?ԙu?��K�D��>�����> ҽ�]�=;��=%A�=Ͼ>�&?[?�.?oE���C�ۋ�������0�i�=�)�=y��>���>�ހ>���= R�<�tr=q�Z>�>��>�#S>p9�>��>�0��	-�xa7?�ڶ=�T�>d�?�fp>o�=���Q>5O���uC�J�O��O�;�`�ʱ��@�`�E�=s��=���>������?�Ks>QԾ��6?S �5=��M7>��8>�6���?�@ =r�=�h�>	��>e�D>���>�6>��e�=����'�1��t�P�����;N>�↾5	�C� ��N!���d��ױ� q�ۚw��8y�A�C��Þ�Qt�?8���o'b���%����
�>N�0>�K2?xp������7�=�^?v9�>HdѾ�\���₿|žS�?�A�?�;c>}�>q�W?1�?j�1�_3�MsZ���u��$A��e��`�2ߍ�9���{�
�y���_?��x?dwA?U\�<.=z>��?=�%��؏��(�>x/�$;��m<=$(�>�-����`�ŧӾ��þ:;��<F>��o?�%�?EU?�RV��쀽� >�qN?F�c?W+=? �6?�V?�s���U�>��=(M0?�??�6?l@?�?ap�>�X�>aˑ=�r�:J���ű�������Y���b�+>�e7>;c����j�泣�+���2=>�4���<�L�����O��=� �=�7>n�>�w^?:�>�i�>�4?��i3� �����2?���<CW��t߈�����������
>Eh?w��?�$S?��l>�@@�͇F�q�!>ゔ>��>"X>+�>d���2�'�=�B>�>s[�=�V�9�i�r�����݉=�J(>F��>�6|>�ߍ�U�'>8����z�d>�R�_�����S� �G��1��ov��L�>��K?u�?CZ�=�T���`Cf��")?�^<?4SM?l�?��=��۾F�9���J�3��>�9�<���j������	�:�-�:��s>�!��H����X>w7
� ����i�P=D�Lzܾ���=�=�F�0=�*�I�Ӿ��Y��t�=�>�������{�������J?�2�=�ן�z�g��g��ԫ0>�ې>��>v��Myx� a9������_=��>�QA><M��W�羦C��1�'_�>�:E?0�Y?�s�?[4��}WV���G�
t��2��	ǽ�FU!?�{�>�?����5]>�8������U���M��S ?��>��?��ze��kr����h���Q�>���>��>�>�G?�8�>��^?�')?���>On�>�!�w7�|-?�u?Z�<.$���Q�/4 ��^7�q��>�!?
8�tӛ>P�'?�.?�V?�Jb? '?��=�z�� 
)�8G�>��F>"e��Ľ�S'�>��I?q��>!\?O��?�6><b]�+ޠ�g���?�>[�=:7H?E)�>v�?}OZ>f/�>���F��=$^�>�bc?�>�?�Ip?���=��?��5>���>��=�B�>���>u?PO?�t?3 J?W��>ͩ�<j����T���q���Z�_�$;S_<w�v=`���~o�"��S�<�5�;�8��g�������D�#��.� <
L�>�l>�U���J.>����~����H>�F���࠾z��>�6��ü=mU�>$?tݓ>��$����=���>	&�>�,�!�&???�b?T�<��a�[�ھ;�Q����>$�>?g��=�Al�p��yu��l=B,n?��]?BsZ������b?�&^?���uq<��þ��b�`)��
O?��
?G��M�>?~iq?Ч�>͇c���l�V���JSa�j��`�=�j�>w���Hd���>��7?��>��`>���=��ܾ�,x��T��j?Ռ?5��?��?��+>��m�n�A[��e���&�b?��>����'�?���<��̾s����Q���׾j����'c������'��ց�ا��O*�=7�?FNm?9�o?��V?�y���c�I_��H}��DP����7��C�.E��{D���k�GW�%��4������<P�s�o�D�vº?O�?�	��S�>��k�6�ݾ����~�=!y���A0!=)��#N����9<�S�����|��E�?�_�>�>�a!?H�j���F��rH����ݾ��]>%��>#j}>ɱ�>��*���>���!�������ɲ��]l>�"s?�T?��?�u�!�
[��@e%���=M	����>H'�>4��>ˀ��0��Cپ�b#�L3����8���r�B@C>�?�<>�W�>�k�?�A�>��g�߾����1�2��_�=Q6=�r?���>'��>��-�euR����>`�n?���>���>������"�����˽5�>A?�>�?�Vw>�z7�$Z��
��M���M9�K8�=m�h?/ꄾzY_�]�>�8P?>-�:��<w�>dg���>��Q��+1(�ui>O�?Bܺ=��H>Ŷ�����TFz��m��ԁ.?C/?aġ�d�2��M�>��#?�z�>ZU�>�*�?��d>AӾ��=�?:�k?��R?R�>?q��>�%:<�go�E{��������<��>{
e>q0�==J>��N9�|��ꔾ�����=?z��7Y��8>�C����=�s��&R"=m4ۿ��J�ωھU��tz�p�
�MZ������Jم�D�
�����sB��1q�ؘ���%��0O���c�����v\i����?a��?����X%��zD��Q�~��:���	�>hIp�,V��F�����������O�����n"��P���i��d�2?���̷��v���\)��1?��'?��u?%���)�-�"�{b�>T�=`�h�J��s���֦Ϳ��3�ԑk?�t�>(��	�`�DF�><�S>�y>*p�>g-[���ھ�H�;�?�] ?⋚>X�0�}N��V���C��	��?{� @0&A?�(��`�:)4=�M�>F�?�R>>�_-��P�$���̯�>�7�?�Ȋ?|�L=�W�F��",d?v�*<�E��䵻���=�ϡ=��=�]�j�M>iȓ>$~�	�?�����c7>��>��V��a�U�<�[>�jӽ���5Մ?({\��f���/��T��	U>��T?+�>S:�=��,?Y7H�_}Ͽ�\��*a?�0�?���?%�(?;ۿ��ؚ>��ܾ��M?aD6?���>�d&��t�߅�=�6�F���|���&V�_��=X��>V�>��,�����O�J��S��=�9 �6ο�Un�~ݑ���>.wþ7��=��@�n��>w^�>~e,�_�[_2���#�и(�0�F?E&?!��=�]�>,�0?H�U?��>��8�����PA�����͘>A����i��ɚ����JF��4��s��㠾��+����z�s��;�klf=�{K��b��w��]T��7��0?��->�/žRYU��A�;6���.̵�#��r/r�e�˾��A�b]��5�?f�<?�{�āV���
��a�<��ؽD�L?u������	��!�>��R�>=�ז> �K�-�ھg�$�V�K��*5?v�?#�¾>����I>Y]��W��=�:?�j�>�2����s>y�&?��:��M��W�>�>>2�>�9�>�3���g��]0���f$?K�f?h�z�lI��U��>@[¾%���iE�C: >������h��=J�=IL��܍�<7}����Z�T?&q�>Ɲ(���:�@��k��Y��Lt?�}
?��>�MP?��X?B1>��Q�Y����W�#=ͲM?�^?i 6>a��۾�艾}s�>4t?~��>���,s��7�0���B?�#r? � ?{��r��5��ྟ�=?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>���������=��vQ�?5��?*����85<% ��+k�bF ���<�=���Yw)�*���
8��MǾڗ
��1��?س�6�>"T@����>#�8��
��QϿ>����QϾ#�n��7?j�>�&νt����i��t���G�EH��Ҋ�=��>��>Ӓ��2��H�{��1;�$&���P�>K*	�2��>e�Q������ƞ�,�<Q��>F��>"��>�>����,��?q���Eο�ޞ�U"�NX?y8�?T�?$�?�L`<�<w��8x�)��ԋG?�9s?��Y?�(��G]��F*��x?�W���5G�ĉ�	Za��O�>��?��?0W��A���>w�>�*!�(	���:��p�Ŀ�%G���?؞�?�aᾇT�>;o�?��,?�����9���`ھ��,;��B_N?���>(��Jc��e��ʄ�2��>�2?������9�_?|�a���p���-���ƽ�ܡ>��0��g\�OK����2Xe�!��/Ay����?G^�?(�?
��� #��5%?��>�����8Ǿ�	�<d��>�)�>*N>�T_�ٳu>����:�Mf	>C��?�~�?j?ԕ������9W>�}?��>��?0��=<��>f�=���JT��">4A�=�"C��?ڭM?>k�>w��=�Z8��.�uF���Q�A��b�C�]b�>\�a?5VL?�a>�綽#�0��!���ʽ(�3�}��1@�-I'��D�y�6>�>>��>�E���Ծ��?l��ؿ�g����'�A?4?m΃>�?4��J�t�i��>_?V{�>�3��)���(��h�����?[F�?��?��׾��˼�8>��>IB�>;սiǟ�����7>{�B?�h�oJ��U�o���>+��?��@�ܮ?�h��	?���P��Sa~����7����=��7?�0��z>���>��=�nv�ܻ��V�s����>�B�?�{�?��>�l?��o�J�B�k�1=DM�>̜k?�s?�Uo���Q�B>��?!������L��f?�
@}u@[�^?,Wgտ�-��Ҁ�(�6� �>>�s�=U'�>󘾗��=�&�>��l���ڽ��]>�Ĥ>/+�>WB�>���>cv%>X�G>ܱ����&�^T��F<[��� ��>�����C��쾴�G��I�2����.����mĽFԀ����=�J�����; S'>U\?�O?P�t?�	�>��L>�!�>�'�e>�=bM��>�=DaH�͊?��[?9(N?Xtd=)܊�\KV��ay�{F��%�E��г>�(b>�?��>�:�>�y��,��>���>��t>9���������>h4�8�>�>+�?Q�>��=4�>1���崮�ģ[�R�2�fX��5~�?s���N\E�>I���Ą��_��	��<Ʋ%?���=����ҿ࿢��GM?e<U��:�\�`�x�'>Mr)?�!,?�=G~��b���ʸE>B+P�z��,�>��������N,��v�>�?�`i>{>�;1��}6�74L��?���L�>�7?E۱��P��4u�26B���پ�L>x
�>��5��P�喿?��[�^�d�=�k:?��?�ԽHZ����x�����Fv;>��P>H�x=�+�=6�>>�%��M�ŵ\�P�#=x@�=*�^>��?��'>�n�=a��>�����}O�-�>�B>'/%>��>?m�$?�*�bᖽ{!���.���s>���>=�>ȶ>%�K����=Q��>�]>?����|��>��kB��X>B~��K�]��x�0en=������=�X�=n���2>�L=�~?���(䈿��e���lD?S+?_ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��L��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>�=ٽ&������݃��s>2]�>��H?6�þ�)�����R0?��%?�������Z¿u|s�`��>��?G�?"�e�Lً���OCq>��?)2s?��a>�d� �����>�X ?�3,?t��>�
�5���j�>���?[s�?wl>X��?�Id?���>��׽�>A�gG���ru�Z7�<j_';��>
�4>� ���?�
6��}��>k��P���	�>d��<�e�>�A��$����C�<�V=b^Ⱦ^�P�
2�>��>�dm>���>�$? X�>a�>�7>�Z���鈾�䡾��L?�ڌ?�c���k���k=d��=��<�X�
?Or3?��@�׾*N�>��T?��?��a?/��>A��W���������Lں<�Q>�M ?��>%bo��_>BB¾ �a��R>;��>�iY��g��C��><=�Y�>� ?A��>�OQ=T?�'0?/$z>ۤ>R�/�O����i`����>�J�>��?�.�?�6?o��k<��څ��T��˂U�ه�>��v?I?���>O���z��-��(�<q���'W?0Zk?��L�aX*?���?1?�:G?ua>[Y���оxfd���>,Y"?D��W8A��&�CV�'�?+O?��>ZB����?��?�E5��!�?`R]?�&?LA���_��.ȾJ��<���/��@�<Fw��>Ѽ>Gim��ޢ=��>` �=U�p���=�@�D<OO�=m.�>M��=
;;��P��0=,?ҿG�|ۃ���=��r�?xD���>�IL>����^?jl=��{�����x��	U� �? ��?Zk�?e��@�h��$=?�?S	?k"�>�J���}޾6�྾Pw�~x��w�Y�>���>6�l���K���ڙ���F��]�Ž�����>�]�>�&�>��?q�@>�!�>Ӑ���9�˕��@��FbI���P1��*��[��O����׽�����	ɾ�u�@p�>����N�>�x�>�>��<>O�>�R���>�(>UV4>0&|>G5>�NC>��>���8�9�zR?�����-'��3� ���ɫB?Z�d?��>9�r��r�������?1�?���?�-r>��h���+��c?A��>o/��^	?�@=&������<�|��P��jh����'�M�>�̽��:��N���b���
?8�?�4��?Ⱦ� ׽D)j����3�?�e�>ʁ���i�BAa��K��pt�dR��λ� x�A)���v���� x���_������H�=P1%?���?�^-�T����Ҿ�u��5m��ܣ>�@�>K`�>ܔ?L�>	���^8��2���c�¾�`�>)p�?�?�>��C?p�F?G�k?w�e?aU�>���>\*���?i��=>�Z>�rT>|�?��d?��?
�?��G?���=����u���v�?P�?�?J��>=�?�Ϛ��@p�=��<N�6�, �=��>�3����=1��<lQ�:}�s>IR?���ׂ8�����^�k>n�6?`��>g��>�N���̀�%2�<���>7v
?�>����Spr�f3�V6�>v�?�� �#,="W)>�O�=�����н��8�=�w��0l�=�܉��8���6<��=���=Dڳ��f �;�;y�;U��<�T�>ѥ?Q��>j�>A���w� ������=Q�X>��R>��>&�ؾ�m�������g�7Qx>UK�?DS�?��e=���=ԯ�=�;������	*�z,��ah�<c�?�A#?S T?�w�?�=?r�#?i>�@�0���)���Ǣ���?�&,?s��>����ʾv騿~Z3���?c[?E+a��_�M.)�׀¾l*սi�>�/��~�t�vD�|]��2��d!����?)ŝ?�6B�@�6��b��Θ��p��f�C?�^�>�ɤ>[��>��)��g�6$���:>{z�>�R?P�>ؼT?��v?��\?7#>�7�����0����7<V=
>ybJ?�K�?�܊?C�l?l��>�w!>*S0���Ծ���SJ��O��n� �=�h;>"��>���>�t�>�>�����P ��11�>"�W>�?�>�(�>8��>��`>�c����G?��>�\�����rݤ�Yʃ�Mc=�C�u?��?��+?V=t���E��=��<�>Tf�?���?v0*?8�S����=7ּ�߶���q���>Jٹ>!3�>h�=��F=E>z�>+��>r��#W�\u8��_M���?�F?⽻=(���-C�(S���Kྐྵ��=���3N��=1e��1"�=m��ٝ��U�����E�s�|�Q��U�����K�Ee?]�D=��0>�!ǽF邽b(�;��V�=�8�;ב=�U��X"�=Į���\d=�H��kL��=@�=!�R�˾r|?�J?\�*?LWD?>�x>h�>4^6��=�>�O5?JV>JY��Ѽ�f�<�ʑ����S(׾fBؾ�d��Z��� 
>3�S�x�>~/>���=�<t��=B�n=�a�=� ����= �=���=?��=��=�y><�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�c$>�6>SxN�j�D��$�79:��%����?�J�^/��6�>�r/>%��:%־5�v=21�=]媼�xF�@�� =>�@��:�e=�!�>ܳ�=QtE<�8⽙&>�V�=�C>���>�����k��������>�N�>��:>d�>�?b41?�e?�B�>��Q���ʾ�̾E��>���=r�>��"=n�5>"?�>ִ8?�d@?m�J?'�>-v(=�>�P�>�o*�u�i�� ھ�Ԩ��Y�<$��?�0�?w:�>lR;;�X-����O:��-�?��5?�?2/�>�T����)'��-�]䕽|�Z�Z(2=G�t���C��HǼ�ƭ뽑b�=��>w��>�z�>.0>l�:><�O>���>�>���<�=�����۳<3�����=�}��y�<:Xؼ�8"������1:��ȼ�q�;�9�;^��<:5�;���=q��>��>_��>���=�ﳾ<�/>������L��'�=� ���	B�Id�h0~�m�.�m6���B>�{X>p����/��b�?�Z>c&?>Ҁ�?@$u?��>�����վBQ���$e�3wS��ٷ=/g>��<�G;��6`���M���ҾO��>*:
>���>�k*>�j�)�%���w>q�C��+u��~�>��Խඛ=V)�X�M�O����h�W�)\c>��T?�ĉ�>cֽ��?Dr?�ߗ?o��>�@P>�v���-7>I����u�'�����s�Ьؽ�??�=Z?�H?� ��h���˾�,��o��>~J��O�9���ż0�M�u��
��>���Hо�&3�!W��f揿�B�"Jr��ܺ>5�O?�ۮ?4�a��/���bO����bm��Y?�zg?iG�>�'?3?���h����-Y�=Z�n?ܒ�?��?�.>�q>��&=$~?��+?���?<��?u�q?������>�k/>9��=�w����<͆�>�>4� >�?.��>u��>��ݽ86�h����Ѭ�����w��ȟ=/�>�
s>7�>_��<��$>�M�='�{>Wr�<
�>��>��>]|#>����>����*?Nm�=���>rp.?0�>G�R=��ܽ�A<ݍ,�b�4�y.��pý�<�jl�<�\ͻ�Ps=.H�a��>�rĿ~Е?�:C>?;���?���[�E�r�U>7�J>�Uҽ�x�>Џ8>�|m>{v�>z�>ʌ>���>�}>��¾t>�_��1���4���?�̝Ծmʅ>�����&5����o����)�2h���X�� �d���|��W;��j�<^�?�Υ��!e��#��'߽�A�>��>m>%??
m�=?����K>:�?k��>���h��� ��-�۾?2��?G=c> �>��W?��?yz1���2��oZ�Y�u�:#A�\e�)�`�*⍿�����
�����_?��x?SuA?q��<2z>ڟ�?��%�HϏ�/-�>�/��%;��o<=�+�>%����`�p�Ӿ��þc4�6%F>��o?�&�?�U?�^V�Ȍ\��p#>a�>?�U<?��w?��5?�yD?��W�R�!?D�h>D�>���>r:?�>? �?%�O>�$>������ <⮜��䏾�fͽ������F��<W�=�e@�e˕���X=�Q�<��߼z<0l;�������<L|�<�b�=���=p��>*]?��>#�>+#<?�<�7�1�I|��w0?�y=\?���u��I��J־-�>]Vg?��?�hT?��B>dsD��N��!>���>`�.>n0M>u��>Uh۽�k@�UB�=]�>C<+>i��=I�=��	���� �J���M�<��>w�?�ə>�;�ʚQ>=�����7L�>,���y���D����=�>�(��Wz�6S�>xji?o?���=�R��R|�S_�׈"?��P?Qe?K�O?�kE>�!˾�Rp���>�(X齟.�>s�Q�kL�!6��I��o�4�dk��6e>�'�`Ҟ�ډe>�������h�D6K��>�pG[=�
�y�i=]����Ӿ7���(�=�W>K���3!����#f��f�I?K3~=߱��W�����%>>M(�>�u�>�P2�̣���+?��@��Т=$��>sIC>�1�����F�Vv��
�>NF?�hb?`A�?+O��<^J�B&Q��T�`�&�ɽ,??{�>�8?�Hӽ�`�=�%��2���B+�V�A� ?a�>G�0�ʇA���u&���X��>g%?h0>d��>!�?� ?��D?86?�t(?V��>h�����h���>?�ދ?z� =�5��m%��
�2/H���
?B,k?T�!�k'=>L�X??�F?3\?�?��>(��6�0��>�7[>F�d����C�W>#D?&�?� �?��b?��=zP��u���^5� �> Tz>h?\@?pU�>u#�=¦�>����%��=���>�cb??�?Fp?jW�=5�?{m1>um�>��=S��>���>g?�0O?��s?�qJ?���>�6�<�&���I���ts��oQ��̚;��D<Fdp=�,���g�;���f�<j��;�X����k�K�ܼ��<��B���<e�>�It>����K�1>1ž������A>r���'���͊��S:���=Ց�>��?��>K#��ݒ=�u�>�c�>g���(?\�?P�?!;smb�{�ھ�qL��7�>*(B?��=�l�Wh����u��i=�m?�^?��W�����Y�b?�^?Ƀ�3=�}:þFb��B��+P?7@?�&H�?߲>=�~?��q?uS�>��c���m��㜿)b��l����=^��>�����d�>�7?�V�>�_d>���==ܾ��w������?6Ɍ?0ٯ?;܊?��(>=Dn�a࿨q��:F��4^?-p�>����"?����Ͼ�d�����G�B#���"���<��ꎦ���$��ރ��9׽��=��?�r?�`q?9�_?�� �2�c��^�� ��PV�n"���E��(E��C��n�T�.7��T蘾FCG=�YO�K�B�9�?��>��qvk>�^��l��iK��F�>�;)��N�z2+>J��<n��n,m&�s�*�Ƥ���4?ͫ	?,)�=_~0?|e��
J�T�[����	��ꇯ>��?`Q�>$?3�u>�ûM@��y~�C%�:�G�e�u>�Fb?ԃM?��o?�W�'E-��s��uy#��h8�;���X�M>��>��>�h�^D���%��>��lm�=7�N;�����c�=�/1?h�~>�>��?�l ?�����-���[5�.�<qV�>��d?r��>�}>u�սo�%�N	�>��^?'�?��>��� ݾ�,��(���N�>�F�>�^I?^��>ԁ&�P�l�?P��[���_2�@�> ��?,~�a�r�i:�>G:?>� =W5>Փ>7�����ʾ�ﾹ��b��!t�>�z�<�ќ>�����ؾ�$[�����<�6?4�?���"�-�޼�>�%'?���>��>F=�?LZh>�hྩM@=��?p�h?�aS?�C?�C�>R_��A�H�\l���Y�w�����>_�`>�]>��F>TJ���y��^�^���[����<�.��ˌ!���=���<�#��~Wc<���=�ѿSpI�����n��Ĥ�U����r��h�����������AžT�l�c9���ò��p���ڄ�l\B�줪�����?2�?б���ξ�쀿�ɏ����%2�>Q�D��#�n����R��e���|���p��=�~k�`�G��`��u,?�~���ǿX������|?� ?��?�S� �U!��z>�=a1�<����1���RͿkҦ�z�P?GH�>���Uu��T��>�"b>��>V�>�w���Ҿ1>�Y?�?!?�4��οᲿ�Y�=Q��?7@O{A?��(�A���V=��>�	?n�?>�K1�lL��밾6^�>:�?��?��M=��W�:
�#|e?^<q�F��ݻ_B�=�'�=�{=�����J>hO�>���JA�Lܽ��4>�܅>-�"���}^�e'�<\{]>t�ս��8Մ?{\��f�u�/��T���U>��T?R+�>�:�=Q�,?o7H�I}Ͽ�\��*a?�0�?��?�(?{ۿ�fؚ>��ܾa�M?kD6?g��>�d&��t�+��=<�-�����㾭&V�X��=���>�>[�,�͋���O�ZL�����=8�@꼿��*���ܾ�Ù���->8�.�����F��|�;��>���;����j��U>/�=��>ux?�Ճ>)ģ>n*B?��T?3I�>2y�={6�=R���⻾N�>.L<�P	��[���d��ˌ��z�M�����]�PdD�ص��|���0�V>3�<��蝿h�x�=����tT�h�,?�{�>.4;��wQ�])�<¥ʾ��i�B��M}����q��}o�'�?�A?��_�1�?�e��M��ͪ�[]?^C�U�P�c��">�z�=Ɋ���X? >C.'�s�"�j(�j�0?W?���z%��F�,>�<��F$=*,?PI?<��;ᄨ>x'#?w2��(���]>1�6>d��>��>� >����xڽ��?|WU?E���e�����>�����q{���Z=L	>�:�1��:�[>X�U<�R��U�J�^�����<w�V?�>k)���}D��D&�q8=B\x?��?R�>��k?*�B?T�<�@��TT�Q��h�t=\�W?t=i?��>�5{���ϾS���OX5?h�e?��L>�fh�C��Z1/�'��\?x�m?��?C��0\}����Y��6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>�������i�=�����?R�?򸫾dߋ:���:fh�(���0=�ǿ=3X'��j޼�4�W�9��"ɾ���BT�������>�@�k����>��H�w{��οYǃ�[Ͼ=pg��? +�>%X���ܛ�M�e��>t��F��D�5����r�>0<>������ź{�ob;�؏��8�>U����>��S�bᵾmt����7<��>���>ȇ�>롯���[��?=Z���9ο��������X?Cg�?�n�?UU?sC5<��v�b{�����)G?��s?NZ?�%�tL]�Ԕ8���j?%����X`��_4�՜E��R>"
3?�q�>�.�G}�=N3>�r�>հ>�".�SĿ߁��x��'�?r9�?�����>ӝ?9�*?���S���C���,�ӕ_��u@?�}*>���W"���=�%����	?�V0?�����]�_?)�a�L�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?M^�?h�?Ե�� #�e6%?�>b����8Ǿ��<���>�(�>*N>uH_���u>����:�i	>���?�~�?Pj?���������U>
�}?@϶>ǻ�?˴�=��>��=�F��N�����>��=M+:���?o�M?=0�>��=8	9�S�.���E�jP����C��І>�5a?m�K?4c>0�����/�\�!�8�ҽ�2���ąH�-�!����ح4>�@?>2x>��I��Qؾ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�h��=��7?�0� �z>���>��=�nv�޻��Y�s����>�B�?�{�?��>"�l?��o�P�B�}�1=7M�>Μk?�s?KQo���l�B>��?"������L��f?�
@u@a�^?*˜ѿ�򞿇���ݙ��t=�*>���>�V����1��,=���z-�=���>��>J�H>��>���>�S�>vư>����W}%��B��&i��p�>��1���&���ξ��0�꽾ӈ.���y������Q=�񠽖8Q<v��&���_.��bB>g(Q?��W?�~�?���>���='U�>��ɾ��)=A<þ飇=��ֽAQ ?�1H?�
)?[��=�r{�C1^���f��-��82��>�>��6>m�V>�]�>�F�>�}Ͻ��0>��>�3`>�u">�Zj>J��<��>ߌ>��>g?��?�Υ>؟�>�񳿌���`�R���վ���E�?%٭���V���y�Z��z���?,=z�Z?�~�=Ш���ҿ�Q��B?K�ƾ&�L�<Qmp��B?��?�=�=�"��Mu;H�>������>mҽ�Q�������^>O�?�W�>T�|>�{3��E.���C�����\]�>�[=?�D��q�m�6�x�=D���s�3>��>�n	=R3��헿u�����{�5�%=W)>?�u?s˺��ܴ�3d�CǱ�?N/>P<>7�=�V-=L%>L���\��G��=�(�=n>I?H�/>��=%r�>�z����y�-q�>ҤF>���==�K?j�/?�6$���Ҵn� C�)J>W'�>l�>�D>��6�Y)>���>{�|>b>g���v����"GI�1(e>�n��nJ.�D!��)B=O5��Ao�=��6=�&����Z�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾQh�>Xx�{Z�������u���#=>��>�8H?�V����O�>��v
?�?�^�ީ����ȿ/|v����>T�?���?T�m��A���@����>:��?�gY?`oi>�g۾d`Z����>ӻ@?�R?��>�9���'�y�?�޶?د�?+L>k�?��?oG?g�M���[�������=�9���@�>�H
=e�����Y����P9��яl�����7>��r=(>�>��潱Ҋ�8��=ި?�P�~��P.��׶>-� >P� >��C>��>X��>'�>p=+��8�/�kָ��\??8�?	�|�f�]��=m�@>�"ؽV�.?��;?p�2�����>Y;?�x?��r?���>�=��ݕ�a�ÿ���������>�g?�y�>�M��ͦ>���͋��CT>�d>�\Ͻ&#���k;�<��>��?�u�>#�4=�8?C!?Iה>&�>7Z��咿]R@�bM�>'�->�i>?�*�?u�?�r/�S�!��咿�ޤ�j[D����>+|?��?gS�>v�s�gpl��TM�C�(>٧m�ZeP?�	k?�أ��p	?(��?z�>�S�>?Z>��u�\<�Ϙ(=I�>4�#?h���A�ô&�Bc
�[�	?W?���>�w��佚�g�*���ߝ?^r]?��&?����v`�ɾ���<j/�����V/Q<���z#>o�%>��s�L��=E>��=b�r�5<�+f;�,�=�ē>���=�_9�gך�3=,?�G�kۃ���=p�r�&xD���>�IL>��s�^?al=��{�����x���U�� �?���?Bk�?���?�h��$=?�?[	?T"�> K���}޾W�ྰPw��}x�hw���>���>��l���L���љ���F����Ž��� �g>��?���>�"?�T=Mm�>�%����0����~�����b�М6�8F�ʊM�|!�(\��~֨�+r�l�ɾ>疾;S�>;"���B�>�?��;>v.>i��>���=�-�>)�">�OE>X>��<�Jr>��~>�T>4n,�NR?�����'��辬���h3B?�od?A;�>Ҹh�M������À?[��?�s�?qLv>�wh��*+�!j?q.�>,���k
?:=�@�BK�<XI��ɡ�E���V����>�[׽,!:�sM��sf��j
?K/?W��=�̾RW׽kI��\/p=1̄?zH'?��*�gxS���m��PT�(�T�x�Q���Q�<��&���Lm�Vȏ�DT���ւ�4�#��F==��)?|��?���a����Z�h�>?���b>��>�ۑ>(s�>U�O>:����0�.�Z��r'��(����>P�{?1��>��L?��I?�r?��"?���>�?���Ms�>`=�:Cw�>8w�>ג#?<�"?�)I?�@?�(??U�=�D��B�������?2?���>?$�?��>�	ʾс���>��<�Ay���3�R)=�+0=d�=�Ø=�5�uVJ>9W?��2�8�E����k>9{7?�v�>���>n��9%��&��<��>��
?MF�>� ��|r�b��S�>��?����=��)>���=����r�Ժ�R�=m��|��=iM���;�w#<��=�ܔ=��r��1��!R�:p��;if�<�n�>:�?��>/5�>u0��:� ����YV�=_�X>�5S>@>�Dپc|���#��:�g��Ly>t�?�w�?o�f=$�=��=�}���U���������Q��<��?)F#?�WT?j��?��=?p#?�>�%��K��`Z��8
��֩?{�2? ǎ>%g*�!�ھ�v��T�'�!4?Q�?�`p�zb�=�9�ؾ��(>���>ˑ�k[��2��2�6���=����9!���?��?�U=.1�7aؾ�R���%�3�U?�t�>�G>Ug�>0k$��@���S,�F�>KE�>3�S?�̻>��O?L�{?�\?t�N>+l7��>������X:��q!>�Z@?�-�?��?��v?���>��> �+�V�ݾ�-��� ����ԁ�X�[=3�Y>"5�>Ġ�>$��>y2�=�˽bl����D�v�=�_>(t�>!�>���>W�t>OZZ<��G?��>�a����s䤾-�����<��u?���?��+?��=�}�3�E�A>���R�>�n�?��?�+*?c�S����=�.׼�ܶ���q�q �>�ٹ>8�>ܺ�=�'F=GS>��>Q��>F4��`�/q8�::M�F�?�F?Ϣ�=�<��FL�c��A��	u�>�\d��_{��UнX$�=��a>��վgk��T���"�e�̾��ľ\�����@��� ?Y=�=�|	>�2��>̜F�H=�;k >�n�<��>#����%>�ci<~$���ܽX +������6e5�˾|i}?��I?�+?��B?�4z>�>��;�KF�>2����J?@�S>WcL�Tq����;�A#���Օ�n�׾��׾c��`��!�>A�E���>T�2>F��=.]�<�M�=��m=�h�=&}��M0=���=�[�=u4�=�%�=��>N�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>}�5>5�>�R�|R3� mG�&l���a�P�?k7���ž��>�̻=	8㾟=þ�=X;1>"\=���l0\�nP�=8b���S=M�R=�+�>IK>>��=�埽듿=�vI=�A�=��J>�2;`�R�t�%��=
 �=m�e>H$>D��>�k?ez0?%e?j��>��k���Ͼ�E���>R�=@ڱ>�h�=_F>Nǳ>�q7?�
D?HJ?�I�>.u�=��>c�>�-�p�m�FE�>\���>�<Ӟ�?D+�?' �>Qm?<�[4��y�<�<�ڶ�7�?#�2?�T?A�>.3
��CY1�i5�1�E���s>/`V<��ǵY�!�c��ǒ�J9=W>ʱ)?Zq�>I??u� ?�b	?L��>޿�>	�K>[�2=�i�=ze��p=<	g�,�3>�`=#ѿ:���=s��*(l�3E��1w���1=���<��K����=6��=���>V>&��>衖=���W/>Y�����L�0o�=�A��0B��3d��=~�>/�[6��B>"X>6���u2��G�?50Z>.y?>���?�2u?$�>/C�@�վ�L��n;e��uS����=Ҽ>�=�8z;��T`���M�}lҾ��>6�<>�h�>y��=.��� T�>�>'nɾ�[���?6��`�ϽR8��ߜK��������{b�԰ڽ�(?�����A&��6�?�+?Sy�?.�g>P=s�U>�ɾ]Ԓ�����Ҿ*�F�0��>� ?]|�>p�n���D��ʾ
!۽!�>E�O�6�J�����m�+�e>o�v���d�>����|#Ҿ��2�y��Z��UGA�Vp�:
�>�lM?�*�?mV��G���N��K��~���m�>r�f?�ћ>�	?�$?�=��	Rݾf	r��'�=x�j?>��?� �?pG>0F�=��T���>>�?��?�Ҝ?5F�?G�c�$H�>���V>Bt���
>��>��=��>ޝ?�P�>1f?�y���	�%�羻��6����=���=7(�>~�s>��>��=�F^=m��=�G<>C�>B=�>��l>�>tǑ>mq��N��4)?�S�=g��>��-?�@�>�N=�����<�oj�X�E�R2�5�½&~���NO<+]�<�O=�μ&��>x�ƿG�?�U>�v�}�?:}�]0���R>�R>°ؽ#�>q<>Ͷr>��>a	�>Ɔ>Ѕ�>�(>ӾO�>j��WZ!�{C���R�_�Ѿ�z>j����%��h�5X��V�H��A���q��	j��!��=��K�<�;�?+Y��ڪk�,�)�e����?N(�>6?/���i����>F��>X��>�T���{���}���?��?�:c>*�>��W? �?Θ1��3�ttZ���u��&A��e��`�፿a�����
�����_?��x?GyA?��<>?z>,��?!�%��я�y*�>�/��%;�s<=\-�>�$����`�ףӾ�þ6�hLF>�o?%�?HW?�QV�6Qm��'>��:?_2?Gt?x3?��<?��eU$?�z2>P�?tS
?~R5?B�.?�
?bS3>�O�=[h��g.=N��}����ҽ��ʽo��C�C=��=`}�8e�;��=�5�<+���U.Ҽ;��:�5��rV�<��9=�%�=�y�=2Ҧ>�]?W,�>�Ն>�7?A���.8�����W$/?x�6=����r���o;�����,�>-�j?�ث?<�Y?�bc>B��VB�$>-=�>�%>��[>)�>� �*0E�Z�=�>a�>���=L�稁�|�	�ڲ�����<��>~s?oa�>&νE�>�LC�[��7O�>
�P�-������vF�$6�Ɠ��>^L?�J/?0^�=�:��&��J�d��?�[^?�~?QO?�-]��"پ@�[��'8��">���>��M�����~��ޢ��B�N�=rW>�$�N����us>ly�_7�T;>���V�����=��tҞ=~S� ׾��)��=�C�=��'��ώ�4줿TJ?]�>Y{�jo��V��l��=6�b>�L�>8��=�h�T�7�����}�=��>㾁>�������G�Z@뾣��>�D?�J[?Å?x��Iui�n�7�-���2���_ݫ���?���>w�?��=>b��<�nϾ��
��Y���A��W�>�J�>���kM�8������$���>�?
�(>��?lY?��?��W?��&?O�?���>�"ƽ�媾+J-?��?j��;O6����E���H�f??��:?ڄ\���a>��0?�?M$?��??�f?1��=��ж-����>�W�>�GP�����[�>�7L?S�>��m?/S�?�>>��F�¾�����->���>~�7?�r?���>��>4N�>�����\B>��>+�!?��|?(q?ΤT��f�>�,�=��>G_�>P�!?";?�4?�gv?\�?��x?��?U���g�<���������>�G>��<���>�J>�M���Z)��Ka=r�>VR�=JT��D2Y��]�<��,>E��=r��>�r>�X����.>>Lƾ�����
A>j���zM��� ��H�4��ص=��>��?u��>�*"�I�=���>�6�>��	l'?(:?	�?ȗ�;��a��ھ�P���>	�A?'��=�+l�&x��۱u�vb="nm?�^?��Z������%f?�}s?o ��0��Kk� n¾^
��rX?y+?��m�@�c>I6�?��k?���>	�]�H�8����]�
Y"���>�Ĉ>@�#i�l�>Y�9?Ᾰ>Xq�>���>'������� ;���>�	�?��?֊?�$�=�u�PпJ������o^?s��>6���y�$?�G
�mξ�3���ꉾH`޾�_���ݬ����G����N#��郾dg߽���=N�?��s?�q?>`?6S��e���`�{~�fV��|�Xk�e�E��B��qC���n�9���Y��5+��*�u=�i��RU�s��?�?B ��J ?;�y�F�ؾ�����>Yj��}���x���#�,Z�<C�=<9g�F'u���Z� d?!2�>ۖ�>�HA?k�l���C��R_�
�t����">���>a>�y?ӟN���f���D�y˾(�,���=�r�>b�h?�@F?�g�?/�p�����݁����t��"Қ��K�>gX>l}�>�O3����/>4�i�!��}O�u۾��������O�=��Z?�X8>ط>��?�2�>@n0�2�1�=v��<UD�����R�>�?mN">�y�>xn�;]|G���>�Ln?>^�>���>�?����`�|��ؽ�c�>D[�>4G?H@�>㣘�5gM�F�������q�,�~��=��a?4��m�؄�>qA`?)�l���]=2k�>��K��j-�4��i�:��]|=�y�>a3�=2�=���F����b������`)?�n?��l�)�7D�>��!?�E�>�x�>�Q�?1Ӛ>=ľqK�:�'?z8_?�J?�sA?|�>E=�ޱ��?Ƚq�&�3z*=�ن>�[>��x=�Z�=+)�UA\��� �.0;=�@�=�{μAL���#<�о�4�[<4k�<��/>#Nٿϱ?�k���9��۾��Eo����9��b���( �Uj��<u��KZ���cd�����f@j�P/�6V�@��p��?#��?�r���Dd�*����t��ྍ��>>��%߽O���29���k�qT��|��~��BJ�f�����H�v�(?"A���Jȿ�|��N��$*?�?8�z?'����!�V6�t>*��<i�H���{����ο����1�\?�E�>	��Oğ����><#�> U>�Hu>�������<�Z	?l�*?�W�>"af��0ɿʹ��<���?�@��9?�_�9ƾ*�3>���>G?Tp> |+��%0�in��>r�>���?�n�?�p=��p�?9N��GX?H�O=ٖ;���(<�q�=���<В���� #>#̫>8��i1��P*����=Ϲ�><���\�i�Y�Ƽq3M>��u�)�b�Մ?�z\�/f�`�/��T���S>��T?�(�>�8�=2�,?�6H�}Ͽޯ\�-*a?�0�?��?��(?�ٿ�Oٚ>a�ܾy�M?D6?���>$e&���t�4��=�Sἒ���Y���%V���=d��>;�>��,�����O��d�����=aV��¿���]�(��"����;��ͽl�����½]�z=Ȥ��<Ў��+��$W�r��=��=n)�>�s�>0^�:�db?�ņ?�T>�3�</P=]Ҿ�O��J��ΰ߾�|���ǽ-/���˾x{ξUgھAJ�P��C��4Y۾�^�P�D>�b��l���U)���o`��E@?Q��>�8>�y�d��Qt�Gҕ��������OY'�S9���n����?F�<?�@N�_U��o�U�,�\��\T?���;` ��U��"�>q�=���=)�>���<l�4��),�U�)���0?�a?�=��M͎��")>g���t =�>+?�H ?��&<���>�t$?W�+�k��y\>��4>+͢>�6�>ř >�D��q�߽�2?��T?I�W��7Б>;¾44����_=zL
>Q�:�NF����X>~�"<�Ɍ�cJ%�Ϲ����<�W?�ˍ>��)�WM�W��Z�@=�bx? �?w��>�k?��B?��<" ���MT�����,x=!�W?�h?ֽ>����,о����=e5?�ce?�>P>9Kh����/�md��G?��n?,?����l}��꒿S���76?�v?��]����G(W��>�>"��>P��>>97�s��>O0>?�{!���� ����3���?�@���?�r<4���o�=�`?L��>�^R�=�ľ�9��a����Ts=_��>�����v�u��#|1���7?s��?���>Ώ���'���=r���ژ�?��t?6H��,�=���FY��{���>YF5>�Z⼾*��D��"�8��ɾ�B
�2~�����=��>Φ@��i ?�0������tտχo���ɾ˂��K�&?f9�>z;6��Q���yp����HR�q�(�0E
��Y�>��>B0��@��כ{��P;�����_�>V��ٿ�>HsS�s[������[�-<��>A�>�W�>�鬽s���d��?����z"ο����#��SX?�_�?W&�?�?9�O<L�u��%z����I+G?1zs?�3Z?��)��1^�DY5�-�j?``���V`���4��ME�� U>� 3?7H�>ڙ-�q*}=�>>3��>�j>l/�8�ĿLֶ�a�����?���?�q�p��>\��?it+?�a��6���\��9�*���<��=A?�2>����4�!�k,=��ג��
?4�0?��� .�u�_?n�a���p���-�A�ƽ�ڡ>�0� n\�Zf����hVe���?y���?�]�?��?���o�"�6%?�>垕�d6Ǿ���<�}�>�'�>�,N><W_���u>��!�:��p	>ί�?F~�?Jj?ܔ������cP>��}?�Q�>�?���=%��>���=�а�T_���6!>���=�&�O�?��N?{��>�3�=�-7�n�.���E���Q�8.��C���>sta?�0N?�=a>�~���6"�t� ���ӽ@8���t�C�$+*��ڽj�/>�;>��>�+D���վ��?Mp�8�ؿ j�� p'��54?0��>�?����t�����;_?Qz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�>9�>�I�>C�Խ����Z�����7>1�B?_��D��v�o�y�>���?
�@�ծ?ii�8	?��O���_~�����6�4��=�7?�'���z>W��>~�=Mlv�h�����s�[��>mC�?<|�?���>��l?�o���B�[�1=/G�>3�k?xr?��l�����B>�?`�����QN�f?��
@yt@y�^?0좿sm޿s��*:d��ܿ���x�
s�=��:>3UF�X�>�s�=i,-�p�(��к=A��=Y��>He�>0Ō>8�'>��1>2����U#��[��
u��u�Y��v�Ȯ�����ķ��P3/�Q�R�ʾ^��Й��A�<��F�S�m�;����=F-U?��R?Z q?}V?�a���'>���Ug�</(��G�=�}>}�/?<�K?�h)?
ڑ=�Q��G�b�B@��ǧ�˧�����>I>��>��>/e�>r)ϻ;�I>|j=>��~>���=�"&=����j=lKJ>�(�>)A�>�̼>�N�>9�b>�fĿrٮ�h�j�f�ܾiŚ���?k��Q�/�Z^u��Q����#�>ed?B�%��̣�݆���J���YA?2��]�Q�~=�4�H?��b?=!Ҿ���� �>������J�/4>�мr�f��!���>�c?�Z�>�|>tc3�Ƴ*��B��Z��;x�>|�3?C(��ƝY��"o���@����Ƕ8>���>E*�;�I�����ㄿe\p�e� =26B?���>�۽�~����R��͹��U>8A�>n��=�}��$F>��ּ�}"�@2P�	{=d�@>���>� ?���=��=N��>�;��L&�D��>q���v�=�z.?�#?�(��J ���g�Q���J�>'(?靓>�>��_�N#�]�?�v<>�}F�$�ܼY�བ3m�n��=M��y����a�=��u>�X�<�>�=IO�O�g���d=�~?���'䈿��;e���lD?R+?k �=O�F<��"�A ���H��E�?q�@m�?��	�ޢV�>�?�@�?(��K��=}�>׫>�ξ�L��?��Ž8Ǣ�Ô	�$)#�fS�?��?_�/�[ʋ�:l��6>�^%?�ӾLh�>�w�QZ��@����u�G�#=v��>�8H?.W����O�F>��v
??�^�������ȿ�{v����>!�?���?C�m�|A���@�*��>��?�gY?"oi>�g۾@aZ�:��>ݻ@?�R?��>�9�3�'�l�?�޶?���?g�`>�y�?Sp?F��>�@�چ8��Gÿ��P�~<̟>�Q
?�y>�ڧ��it�v���.���ti�����?�K�=MK�>Tbl��˙�h��=�X���4��kG,�3��>��>�z!>E��>��?��?f��>�$X>s3=���9ͳ���W?Iԏ?KY#�V?��{p>�=	M����N?�Q?��5�rI�j��>W�K?dy?��{?c��>�Y��ڕ������ȭ�8���8>�E�>�r�>�o8=��>����׾\��=n-k>�x���������;�@>od?F��>�薾8z?ti6?IL\>�I�>��P�O����g3����>]d>
7�>	E}?��@?,v但�,��%���\��n�8�&�e>w�l?��?X��>�ۍ��^���*>�S������٠\?��?�*>礡>�ӏ?4>?�u ?�۲>�a>Z2پ�ߒ�E�>/�"?t��E�D���&�7� �j�?#?y!�>������۽�ü� �'��wm?M]?��#?���=Ba�c
þ���<�����-��:�;�)m�K�>��>��x�� �=�#>x)�=�t��4�td�<��=E��>���=3�1�s�j�Jc*?���B���Sa�=5�m��A��G�>��!>�S���6Y?�}2�e�y��`��X����q;��+�?D��?�ʕ?����(�d�� 2?��?��?�]�>�?��E ;W��{����dR�����e0>�r�>#�<�h۾mV������Z��nU��½�����>���>t�?]Y
?���>WS�>�￾6�1�M�����޾#?h�}e"����J(���!$���W5��ܹ�M8ξ'+f�q�>H�'=@
�> �?g�^>��=d��>�ܝ�C�_>��.>�l>��Y>���=� �=�>�F>��>�eR??���v[(��� g����A?�d?�*�>�vk�TU��e.�i?Z]�?Kj�?�Ow>�dh�!�+���?���>�d��-�	?��<=�R�C��<
���h@����x[���>��Ͻ �9�b�L�6�c��	?�+?c���c�˾�gѽ�%����!=s�?�?�-.�RA�]h}��0�g�W����=�q�:п��JR�B߂�XE��s����[��.c���>��&?f-�?������~<Ѿ�ل���U���>z��>>t�>Ny>A�꾘�@�KIV��P��'�� �?�r?ID�>��@?��Q?��p?�MS?D�>��>뎸�g��>�m�Z��>支=P_?N#?K�?(8�>U{?wv>y)�<��������'?&X8?`r?��>r�>5��z�tw����"=��=�j]����	>t�J>�Xڽ��ֽRX�<�g�>?����Z7��=��3�d>Ԥ7?�8�>��>a�����=��>W?	�>����s����Ϟ�>���?r� �Y�=W'&>U��=�a����3�a��=rǼpd�=L���]�E���l<���=Q�=P����<����:���;�س<���>��?��}>$��>	�u�2���A�0.=�iU>ʀ6>>�����&��+aX��>�֓?5'�?���=��=}��=�����G��2���о6B�=�b�>�?��\?O�?��A?�2? �>�D����+憿ّ��

?�r4?�o
>�XA�����r��0��` ?��,?z�c��=�Q�.zƾ�璻�V�>M���bR��骿J�I��=�t�H�����?g��?CB�=�9���/%�����C�k? ��>;�|>��>4�Ծ�Sq�U�Ⱦ�^�>"�]>�:?�>�>ߙV?:*i?��M?�7�=��2�>ݴ����ύZ=��>׾W?�ي?�G�?��Y?�)�>a��=7��cϾ����G���<�S!t�+Jj>O%=>��>ܡ�>-�X>?�=J��(������7>��>���>8m�>���>�m2>P����C?�f�>&Ƚ�����ѣ���U�$Z8�NCq?z�?��(?S�;=?�r�=��K�����>�E�?K��?�8?��3�T�={�=�,'����b��o�>8�>��>�{�=�Y=q�Q>6��>�ä>��&��4�zy1�CC�;;?b�A?&O�=5���xC@�]签��Ӿ.T=ʨ���1�����ѱ��{><٬��ॾ<׾X﴾I���U�ń�z���r�ž�a?��=\Z$<�|�=y;>މ�%��;;1>XΎ=W�	>�֋���=���=
s�="X����<�ѽ��R�vg��N)����z?��P?�q6?39H?��{>��7>��9�_!�>�ճ���?U#>�2��P��� i)�a����ґ�q�˾����j�k��@����,>Z�H�d�>9>�%�=�������=��2=��r=�l�<"�<�m�=:�=�ޞ=�&�=�o">�>|�u?�#���Z��d�J�A~ݽx8?��>T�=*�þg<?%�=>�I��Mҹ����3~?�d�?���?�6
?��b�	R�>3A��"����Մ=uB��ڥ >ne�=�.D�x&�>;�\>(��iř�}�{����?��@2QA?�H��UϿ�6>�>)>�Q�u�2�_`R�Ǐc���a��[?E5�&l¾n�|>�=[W��P̾�/=��7>�zb=�#�9R]���=,h���=wS�=[�>3F>}��=�睽�M�= ��=�T�=Y>��/<���#Za��/=ݦ�=��e>��!>dZ�>��
?�,?8�[?]G�>=��d��vW��!ߞ>]V�=P��>���=Q�`>Fa�>�T3?`�F?�T?>Q�>|��=Iv�>l̞> {*��#h�R#�=���ey<�	�??X�?���>/��<�nb�ű�C�A�����?��2?m?��>'��i��i ��1�Ў����>T >������_=ּ֑��Ǿ*���i@�:�j�=��>��>�I�>-�a>{ӽ=���>��>yeս�=֐�=�Ը=�������`>����|=��=/c�=��,�n��L���m@������x>����B��="��>��>[$�>���='賾��.>�|��jN�hI�=u���q�A� ]d�C�|��V.��6��N>>�N>\7��#ۑ��� ?�j`>��=>��?)�u?+%>�-�p�Ӿ�����k�6dP���=���=p�9��:;�c`�:0M�ڮѾf��>gd>�Ț>12>I�(��@���U=.!־�kJ���?�u<���h�BH�KH�`C���Ĕ�%�b��"��4?#����C=���?V�:?fқ?p.�>	�s�x��+>:Ձ���Ž���˩�D�9�.~?W+?>�>������I�VH̾Q��'߷>[@I�5�O���y�0����Iͷ�1��>?�����о_$3��g������.�B�SMr�V��>Z�O?��?9b��W��UO����K)��nq?�|g?N�>�J?�@?%���y�r��&w�=��n?���?D=�?A>���=�ی�%u?wM	?�D�?��?�=w?�웾��>;�7����<�n���=X^>��=�:>t�-?of1?�{?Un��ی�[N߾�۾񔤾�1>@�T�Ks�>�Ǘ>\FU>��=���=l�L�aL�Z�>��>=A�>Š�>:�9>_����!�..?�=ZW�>V�:?�Y�>�H%���:��X*>q�l���孨���̽#�<�/~�7���)ļ�1�>���m�?�B>3l쾆�,?��ξ�ػj��>
@>u�ϽH~�>�,E>z>_�>���>��<>�ޤ>�z>+?Ӿ w>����e!�F(C��R���Ѿ��z> �����%�=������yDI��g�� d��j�.���<=��R�<;E�?������k�!�)�b�����?O\�>6?�ڌ�������>h��>�ō>�?�������ō��j��?���?�nh>���>��`?[�??��;�o=��*��ie�����k�Z�P݋��.��� ��tҽ�
X?rC�?_�X?��=i �>}�8?r��)��ʾ>T�/�PK.�T�<c�w>N.!��+Ͻ9�־ӧ򾷧_���J>?�?Ґ�?Ը
?�O��7t^���->�x=?[D5?�Ju?�0?wL<?�����#?�'>��?��?�x1?�}/?r�
?��->���=B׺�L=�ښ��놾e糽|�̽��ܼ�F=��n=��ɻ%�6<S�=��<��������;��<�[��<0J=���=˕�=>F�>��W?�w�>R1�>?3?F���_.��o��I)?H�&=�z��q��d��s���a>0p?*9�?[?/k>��C��*R��> 9�>Dv>nM>��>:@�O	[�
��=�>�A;>�	>R���t�&�������&��j(>:�?A3N>q1���	>��^�E�I��;�>�c���g���<�,��^ �GF���3�>Q%?F�?��\<�0�kƫ��6P�X�>��h?PJ1?��p?�l�>8{���p�G)>�����<>5�����$�
��h����)����;�D�>t^T�.l���}�>m_	�,���O�� H�^ ��)?A=�`�,�=љ��Ϋ����s�=��>�Ҵ�����4��㣦�[DN?sE�=)���� 	ǾM��=T��>��>��辽O�(��ǐ�[��=0��>�oS>��K=:ھ�K�~��<��>��B?Lx@?��?�_l�-(Y���Q�r�]B���~����/?�̔>���>㫜=���=��N�~s���Z���#�7V�>h.�>^"'���i�=�ʾ���`R"�,�>\�?��3�F�>u�H?�?��|?�!+?���>J�k>+�C�S�Ⱦ�^6?�?eH�g��̽[\4�q�8�f��>X7?����޽E>.y�>W	�>��/?�(J?�"1?A�콅p��b/�N_�>aDQ>_^H�=��;��>��-?��?��u?D�{?���=��j�⌾�1[>�8�>�X�=��?f(1?fk'?U���K�>m����6�=bK�>@�b?�ބ?�o?A>�=�?j�,>5��>��u=/2�>XH�>i�??�L?�t?�)L?PJ�>�`�;�������G~��=����:��@<=�=����{�'����4>=*�<Hi��ַ�(���-�Ü��v@6<o��>ws>�����.9>�lþ������B>Iӷ�i����X���Q3���=w�s>�?bU�>1�5��a�=�i�>II�>%f�>X'?
C?��?o���Hk_�D�۾��b��@�>MGB?k>��o�;�����r���?=7k?�dX?��J�M�o�b?�^?���Un<���þz�c�^�7O?��
?~#J��6�>[C~?yp?3�>0�c���l�����b�5Oj�ݞ�=MU�>ȭ���e�eD�>3�6?:��>��f>���=ܾґx�X퟾ͅ?��?���?H��?S)>gan���߿G"��M���o^?���>1����`#?D>���ϾB猾����߾-9���D��m���J����!-��^����ӽ�l�=�z?eHr?�rq?1`?�� �ڗb��]�{À��SU�Y'��	�JUG�	�D�j�B��vn����t����㕾�1^=\U}��=J��Ͼ?��?�I�����>w"6��%ӾL���AIf>O�u�y�V����=�uV�Ս)�{���#��h���c��?}%�>uE�>��&?��[�:L��Q�8�=�[7��Q}>~�t>z��>��?#�/=E������㢾3U��V-�a�>�]n?�s6?�u?g����3��{��,>���=C���ϽX>�?>���>@q����)���� ��y��q�~����J��i=��3?��>-j�>�L�??�s-�I��x/3�bK�A�2�=L�@?�$�>꾹=��}�������>��l?��>K$�>Ὄ�^!���{��Y˽o9�>��>���>�p>y,��\��d��z���9�c��=i�h?������`��Ӆ>�R?���:�I<���>�9v��!�����'���>fd?��=�;>:mž�(���{��E���S;?�?}�����(�_�>��?̯?�L?�s�?>ͻG���˽�� ? ?�?>??hZ?3�>w�=������%z�����=�C�>�BN>�+�=��E>���=���8��_������=���;#?�s��=�Z񼭁�=�̽��6>cK޿�w\��,߾��� ;�j��v`�ٴ3=�! �no�VOƾ�x���Y��7Ͻ��޽q�d*�Nd��5���"�?9� @��оP�Ӿ$Ά�e�bT'�H��>T��<D��w�b��⃾v;���2�*z�oFH���_���Q�<N7?�[ھ��ǿ�Ĕ��;�!!?��!?}̀?��=��;Ȣ���n>�˚�}�>�+��(��j�տ��ֽ��S?���>UϾ3�Y�]��>���=��J>�h�>GQN��lо�O�=�U(?ë�>�H�><�3�'ؿ�+��@�K�{H�?��@|A?I�(��쾭V=���>l�	?��?>�V1��E�����hS�>�;�?A��?��M=*�W�W�	�~e?'j<@�F���ݻ��=^2�=G=��̘J>U�>m��/PA��@ܽ�4>�ׅ>�v"�����^�G��<M�]>��սDG��>Մ?sy\�Lf�%�/�.S���U>;�T?#/�>�<�=ܮ,?c8H�N|Ͽ�\�l+a?z0�?f��?��(?�ܿ�՚> �ܾ��M?�D6?7��>/e&�d�t�$��=�]�Υ����)&V����=s��>T{>�},�?���O�����g��=/��DҿΚ�X���=�M�l?Y:�ͼ��=�����ʾ�c�������+>d0���5�>���>y�]>�7�=�g?j�_?��>½=�A��ؾN}��Eo�=��F�J�l4h���/g��笾8���~:��}'/����*;��9��0>&@J�+����Ż���J��#L��?OJ7>�#��eNh�x|�=�^������q2(<�\�;泛���@�w�n��d�?��5?>0j��\G�_7���<�/2��B?kx�vǾYӗ���L>qm��O��#��>�m�=^ʾ��7E�o3?�=?�ľ�ܒ�9�N>�9�E�=�L4?P ?յ1�s��>_3?��>�\}��8�{>��I>�!�>�G�>8C�=ު�����S?�T?�'�������>�:ž�����ME=)�=�pE��Hd�s�%>0�=`Ũ���v;����x	=�(W?q��>��)����a������V==��x?Œ?8.�>{{k?��B?�ؤ<�g��e�S����`w=�W?<*i?��>����	о%���"�5?ףe?v�N><ch������.�_U��$?�n?8_?a����v}�m��x���n6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?n�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>������yC�=�`����?0m?����/=������Z�4��S �=��=��=Г�=p��|s7��.� ���Q��;#=(�>fK@�œ����>�����M��R��=�����V��?,��>��2:0|J��TC�4d�|;���$��+��{��>�E>�蚽&8��J�z��:������>�7���>�CJ�/c��;ܤ���<�q�>gy�>�ǀ>�cý�N��_Y�?L����Ϳ|ߟ����pT?�L�?u�?(%?����5��7Gw��к��H?�sr?��X?��,��a���O�""i?p=����a��i$�j�g��(Q>~�8?6��> �5�0Ֆ=C s>���>j��=)8��¿���t1���?G��?! ��
?�`�?�C?�2����R��G�*��sܽ8wd?��ۺ���)eӾV>��R�*��>j�=?��<��˾]�_?$�a�M�p���-�s�ƽ�ۡ>��0��e\��M��.���Xe�
���@y����?L^�?h�?ݵ�� #�a6%?�>g����8Ǿh�<���>�(�>*N>HH_���u>����:� i	>���?�~�?Pj?���������U>�}?%�>��?�s�=4c�>�V�=��,%-��d#>�$�=��>�Ӡ??�M?"K�>�V�=��8�(/�NYF��GR��#��C�T�>��a?ЂL?�Gb>@���2�q!��ͽg1�I'鼯_@��,�ѧ߽�$5>�=>.>��D��
Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�d��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?Qo���i�B>��?"������L��f?�
@u@a�^?*��ֿ���"P�������>�=�=�=�y2>�cٽE;�=��5=��@�ӗ�̘�=�ɗ>tgd>�p>�P>+�;>Zl)>�	����!��W��������C�����T�5HZ�ё��v��k�M��X����R����Ľ�X����P��%��[_�a3�=mU?��Q?�mp?^� ?D�^�m">�������<l�$�Y�=�> �0?6^L?\�*?o=�=✾W�c�/��c5��Lˆ�N]�>;�H>�@�>�>DT�>��s�I>#�A>��>��>p&3=q,	���=0gQ>/I�>/�>���>�~>=�>)�������d�2M����6�?Cą�8�?��݋���Ƚ:<G�(��=��P?r;�=%���M�ſ�4���k?tg��D0��B1�/�~�1?�]?{�8>�w;�����mɻ>X�ӽ>8���E> �=��֩,�=s�>_E?eg>��u>��3���8��K��ĭ��{>�>8?����(D�x/w���F�& ޾�<O>�3�>��:������~��Ii�� W=�b:?��?N�ý����}�x�nl����A>Ka>,�=7�=�E>}B��ƻ���[��`=2��=C�\>U?�/>?��=�f�>~m�� 6A�V|�>��+>w� >d=?�D&?�nJ����3����-��w>��>w>��>g�O����=>$�>.�c>V����i�����}F��sR>^�f�*=J�$��C;=�������=�ǘ=1�
���3�X .=�~?���&䈿��=d���lD?S+?� �=0�F<��"�A ���H��<�?s�@	m�?z�	�ϢV�9�?�@�?�����=}�>�֫>�ξ��L���?��ŽǢ�ϔ	�\)#�_S�?��?��/�Uʋ�$l��6>_%?"�ӾPh�>|x��Z�������u�z�#=R��>�8H?�V����O�e>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾;`Z����>һ@?�R?�>�9���'���?�޶?֯�?��S>�y�?O�f?�S�>�+o����۰�P.���.=��= ��>�!�=��龡IT��֋��v��Mn����'r>��Z=Z=�>����)Ӿ�>�=�H�������:S���>��,>
eN> ��>��>���>���> !�<sW���5}�q��'0N?�?&w�oRl���~=ޅ�=��D���?�6?P1��׾�>nZ?���?l+X?�4�><
�Q蕿x5��76��%�y;[�N>}O�><H�>�U�w&k>6��IK)�z�t>��>
�T�a1Ͼk�Y���|�8�>��'?�j�><eL=�?+N?Hm�>���>�u=�,S��_���>�>�>2�?q�?��=?c�8�c>0�+����휿%B��Й>S6y?T�?@�>1Җ���~�E���Fk�)o�t4M?Y�?WxP<��?���?wQ4?VKN?Y�y>Ձ��?�����ՠ>D�"?
�;�A���%�=��^�?�C?� �>�~��4���K��6����?Yr\?z'?�?�\i`���ž���<�{��ȱ�:�o8<�jp�+>,�>�ч����=�>(2�=�dn�4:�+]�;���=id�>��=�0=� ��"=,?~�G�oڃ���=2�r��wD���>9IL>[��ѫ^?�k=�O�{����sx��_U�w �?Ϡ�?#k�?���O�h��$=?�?�	?�!�>�J���}޾u�ྞPw�N|x�qv�Z�>4��>W�l���
�����6F����ŽM�/��O�>�l'?�V*?¡�>�\�>��>;E���95�쿾�U��}��7A���1�)
��K�I���ۻ��ʞ=W���9�O�e>Sƽ��>+4?�0E>W����>1�>f�>�H7>E�=5`>�ٖ>7��>�	�=]�=�ܽNR?j�����'���辒���&/B?�sd?�G�>��h�Ս�����x?�}�?�s�?_v>�nh��#+��c?�!�>L��Sb
?�:=7b�WS�<�K������_�����Ƣ�>�H׽D :��M�u�f��j
?�?H�����̾�׽�x��f�m=sW�?��(?��)��Q�ɫo���W�� S�4���g�3ؠ��$�i�p�`᏿�]������`(���+=t�*?�&�?��A�gO��$Pk���?�M�e>���>��>���>4dJ>�	��v1���]�P5'������a�>/8{?N��>�	J?H@?��Y?;�L?R�>|�>M�Ѿ�4�>żI�>���>�?t�"?�\:?��?�A4?J�>m���8�� ľ�	?+��>�<?O�>L�>$:O��������G�=0g@���߼B�W=R��=����vh�;�>��_>�X?���Ȭ8�����dk>k�7?	��>v��>���*-���<r�>�
?G�>C �~r�c��V�>���?����=��)>���=卅���Һ8Z�=������=66��7z;�ee<k��=h��=�Lt�c#��48�:t��;)n�<�t�>'�?Ǔ�> D�>a@���� �\��zd�=:Y>S>>Fپ�}���$��O�g��]y>�w�?�z�?%�f=M�=3��=�|���U�����@���4��<У?1J#?�WT?\��?F�=?4j#?>�>�*�UM���^�������?�-?P��>�I�4����(��	01��L?Kj?�Cg��z��.��X��t���9>��>�����=���)�c��=G���O��?Jg�?���K��bվDH��ž%�T?�(�>�P�>�	?4�+�it����b�>��>gxO?�2�>�Ba?�1I?^`]?�ƽ<�?�8��������s�>��?�9?:�?(�?c�V??��>i��>̞�<`b�����V=�Ly<K��� �=�'���> ?���=�&�<>z�Gq�>���V���(>�>��>���>�������G?���>�n��L��Ԥ������z=��u?��?>�+?�l=M}���E��5��0I�>No�?���?>-*?J�S�h��=��ּ�Ҷ���q�n �>W�>$�>���=��F=!�>���>���>&��W��i8�9�M�	?�F?P\�=ү���OJ��씾�-˾Yu">>5��7γ�L���^ǽ�&5>�������bp�wI��D�����d��v��zq��	�?��=J^�=Nͼ!ރ<����G*=�x[=�������yw��Ĝ*=g(F�'��=��м��?� ��lv�y/?�˾J�}?�;I?��+?5�C?f�y>�J>�4�g��>킂�C?�U>��P�È��Bq;�������^�ؾ0r׾�d�sğ��K>�I���>s;3>�,�=�q�<I�=Ss=	�=A�H�8)=]�=�l�=�P�=0��=��>V>�6w?X�������4Q��Z罥�:?�8�>c{�=��ƾq@?��>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=L����=2>q��=v�2�T��>��J>���K��B����4�?��@��??�ዿТϿ5a/>l2�=Ҫ>��U���<��G��ue�s{���"?s������99>�>�=i˾^f۾n�C=A6w>��=i)�ɬ[�ڄ�=��P�u)c=^ �=�c|>+K>� =D��+��=��>���=Q�j>)�<�(q��|.�^<�fy9>_/n>�>��>��?�+0?5yd?�>֖m�Q�ϾW����T�>L@�=Q�>$x�=Q'A>{׷>��7?�D?LnK?��>D�=��>4�>{�,���m�ʃ��է��B�<?��?ۻ�?�(�>{�G<�!A�~^���=��Uý�j?\1?R�?�U�>�R�Y뿎��x�)��m=��=���=� )��`��Ƚ��^���6�ѕ�=ר�>+��>{��>���>=q�>3j)>]�>Z	�<�=�@	==d[�{^�<�c=�A>�d�=��w��r�e�g�����_<F4�uD�=��<�rJ=��&;=�>�_�>3�>l*�>�9�<�	��7?>��ž��C����=�Hv��t7�V�b������-��y���h>���=�����,���7�>hJF>-s>���?.�|?6�>�(�����/��H1��Ƒ�W6�P=��.�Ac"�4=i��N6��v�����>�3�=���>���>G50�{��i�>=?�Sр�c^$?�\��/���U�=Y]�ƻ�f��I�UL>6�|?l����B���?�?0�?=��>�F�j���?�=7J��������0�������?Gk4?��?{����M��J̾Z��vݷ>1II�Y�O�e���n�0�FE��ɷ����>h���Q�о{"3��g�����H�B��Gr���>'�O?��?{/b��V���TO��������l?)yg?M�>�L?>?��Wv�gt��~�=&�n?v��?<�?��
>���=��=3*?�T(?D�?+��?FNx?�إ�ia>��g�MP�>!�S����ϝ
>7�>7`Z<!�?�!B?���>�U��ﾣ=���ľ;L�� �_%�=�@s>��\>�>>�I>t�>Q�=��=>��>�z�=ND>1��>�%�>�\���V��2?�}�=�Γ>��0?�-�>ڶ�=x��O)=��輏�6��D0�����R
��N<Ћ��"`v=Ni
<k��>1������?'y/>N��F??Yh���uy�mP>L�Q>�"�<��> Z>�r>�Ȭ>X/�>��/>Pg�>�>�*Ӿ�b>B���h!��5C�|wR���Ѿ֙z>^���L&�l��o'���'I�[��+O��j��.��J<=���<�F�?�E����k�I�)��<��#�?�p�>f6?�ٌ�6���>���>
��><1��S����Ǎ��o�W�?3��?�?c>��>��W?��?�1��3�sZ���u�'A�Ke�g�`�⍿\���&�
������_?��x?�uA?�M�<2z>ڡ�?;�%��ӏ��)�>M/��$;��:<=�,�>�'����`��Ӿ7�þ)�CQF>��o?�"�?�W?�WV�#lm��P'>��:?V�1?XMt?2?��;?�����$?AM3>�L?�X?/?5?�.?��
?w�1>���=�l���'=���銾�mѽ��ʽ,�3�3=�4{=�Cҷ�'<��=a=�<0�꼄�ټ+�;�{��׌�<�V:=�W�=A>�=ϔ�=��;?�ߘ>9��=��"?�f�-R�1و��D?7�P>V ;�_L�`�����=U�\?s�?ÆC?#<�=�n�B̊�Hb>�9�>�rm>UaK>k�>�����ȉ��:>|3�=�>u�_>�+-=����2r%���,����F>�O?��e>(�޼m`G>V_;��T���>k>�A��:���I�T43�*�����>Q�N?du�>�CB>���O�j��jo�2�>��e?�a?�� ?��!>}&�U�o��Y���
�?�$��$`��TP��Ҵ����h�E����r�>^������(�b>�j�g9޾�n�M�I�<�� �L=<��O>V=��"C־W�~�#'�=�b	>��{� ���z���hJ?s�j=�����T�f���Ƴ>�}�>�ˮ>vG:�T�v�0i@�ݬ�'��=���>�:>o!��jw�/�G���K�>>E?��c?Hm�?B)���g�G�D�������c�A��J?�)�>6�	?�b9>��='������c���?����>�x�>�P�?�;�����������c�>�
?�Z@>7D?X�S?e�?\^?"8*?�6?��>v��z���A;&?n��?}��=eս �T���8���E����>փ)?ҺB��ؗ>R�?W�?��&?��Q?�?r�>� �&=@�ɓ�>%N�>��W�b����_>�J?���>�<Y?�Ѓ?�>>3q5�"���dS��?��=�]>�2?)#?��?̸>���>+�jW��Q��>��w?&�?t��?��t>�n*?=�X>�?�ҹ=p֢>��?��L?'�>?)B@?�O(?e�>�"=ɂ����#�6<o�=�Z���}��4�=+�:Q��<N����%�۲��*�=�=[Vн�3��pl�=���<�T�>��s>0̕��d1>��ľc0��� @>����[/������:��˶=z��>��?���>�M#�8�=ݾ�>��>����P(?=�??���:d�b��ھ�K���>|�A?L��=n�l�ؐ��v��.g=��m?d�^?��V��5����m?�d?�.�0�V���I�u/C����\lj?��?���3�_>H��?[x�??EzP�5\��ߍ��?�[��$���=�Q�>�O9�4q��f�?3�U?�bp>,+ � ܍>zH����z�ah�4��>�Ǆ?y[�?I�?޾S>����������ͩ���^?rJ�>���K#?��;��ɾB,���!�� ��ɲ�XC����������`b$��gv�x��.��=�w?lu?�m?mK_?��	�`ng�0,]�����Q��g�-]�xF�F��:D���m��3�6��݋�E�="g���@����?�+?2��?�������=�����=Z<ھ
�{�1>����jb=�l�;�������LX&?�?�>]��>��@?�8��lZN�-�A���-��.���	=GK�>�1>[~�>�߹�_�6�������L��v���Qv>�tc?��K?~�n?�	�0�����%�!�ә3�-<��&DC>�
>�ۉ>�W�1���S&��N>���r�����K��F�	�^�=D�2?��>��>}:�?7�?>`	�R<��z3x���1���<�6�><i?�5�>We�>�н� ����>Y�a?@��>*>�߾��پԊ~��u>�a>�/
?F!*?ue�>K֩�V�S���j�,���0�2Q�=â$?~�E���n��#�>�a?��+�㥖>|G�>�4d����o�������u?4n�>��<4'���2�����N���n�?CO�>��ƾ[A�Z��>|2)?z�?���>�4�?}	�>��G�;A�<(_?�sh?�tr?�2?�z�>��0=S ؽ.B��q�TL�=��>�~�>��R�*P�<y�����D�ҬĽ�;t=>�=an{�H&G���+=y�����:)��=�E�=,�ۿX�K��>ھ���S�
����m��T��_����s�ihx�j��>�,�U��c�뭌��$k�[>�?C�?7������i���uu��I ��=�>�@q���s��f���}����>�����$A!��$P���h��Rd�N�'?1���]�ǿ*����;ܾ2 ?0? ?\�y?���"���8��� >k�<���ӣ�����ο7���j�^?9��>v�|-����>7��>��X>�Iq>�
��垾i��<��?��-?��>�r���ɿˊ����<1��?��@�yA?��(���V=#��>��	?��?>�G1��L�j���J_�>(8�?)��?��M=i�W��\
��xe?š<3�F��m޻��=�[�=�R=����J>7Z�>'����A���ܽ��4>﹅>�'"����Z�^��{�<�\]>��ս�8���K�?��[�=XD�����7��d�R=35_?p��>�,�sL8?�:p�.Կ��b��4Q?��?-?�?~�0?Ĝ���@�>`�'�I?�yO?q��>d�1���\�?ʥ=����N[=S����f�Ms�=c+�>�0>�y�HZ�Ð��=�ս�V�=��C�ɿ�#4��b�l&�=��`��b�<��ɽ	�����=�L����������S@ ;�d=�bV>
�_>Qd>��p>\#R?d�~?�\�> 5>"?r�ᐈ�������Ž��{�g�<ns�c�@���N��y������$��2��Jk�3#=���=B4R������ �P�b�?�F� �.?�j$>��ʾ��M���.<�pʾ����ɥ������5̾��1�	n�͟?`�A?g���%�V�������dm��`�W?�W�L���ꬾ���=%���	= #�>Y��=��⾟3��xS���/?�#?�o���ӑ��(>e��n;�<GX-?�V?���<*ʯ>8W%?�*(���?�`>!�*>jϣ>7��>-�>���8;�#�?�
V?;��+��dd�>�8�������L=�	>"4�:;ü��d>*#�<�ב��Ւ�$e��x�<�;X?R�>�#�K���Ǘ�����4t%=z��?Fu ?�>�m?ЍF?��_=����O�0��x�<��P?�]o?��>�pO����\�d�<?P�e?U�?>��c�GWᾂ3��`��?!�s?=�?����{�����6}	���-?�Yn?�T����K�پZ͓�7�b>>�?U�>��L�wS>A�0?�<���{�����<�<�xҨ?*2@���?H�#=�ce<���:�?�H	?�y��3�v��-��C�h�齚K�>�l�	<��0V�Tm����G?�s~?�?h葾g%
�Ӳ�=	��U�?�?K���l�l<�>���k�^)��h��<���=����� ����k�7��ƾD�
�1Z��K�¼&ֆ>hS@Gy�e:�>��9��7⿽,Ͽ3��<Pо��q���? �>Y&˽����j���t���G��}H��͌��J�>	�> ��������{��g;�����<�>����>͞S�~��)����b6<Y�>X��>��>=G��\佾�?�b��@ο����N����X?g�?zn�?}n?�:<��v�{��<��,G?��s?�Z?v%�]�X7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�y�+��<A?�2>���I�!�C0=�VҒ�¼
?V~0?{�f.�O�_?(�a���p�~�-���ƽ١>4�0�Ki\��~����Ze�p���Dy���?I^�?��?x��	 #�w6%?��>���w4Ǿ��<,}�>(�>�)N>�H_�E�u>&�u�:��g	>���?C~�?:k?[�������O>Q�}?��>�]�?��=�>��<>������=��={�=Pt5���>F�@?A�>+m>>['�ܿ%���;���]��t*��@��:f>+�u?yeY?�?�=��,>��E�[���a�#i�<����}.;ԧW�Ɇ�=G�H>n�>��&�Z:����?W��3�տ-f���:�܊)?�Ƃ>K�?h`� <j��7��T�]?B]z>�d��յ�����:��ƪ?��?I�?��վ	���>�>9��>WA�>Nl��{;���j����;>�A?=���'��r�F�>u�?1{@⊮?��k��/?ei
�"�z����)��c`ؾ�C�> ?�Ѿ�_�>���>��>Hx��[������3B�>��?��?�q?�W`?��C�N�)�E8)>䅡>��w?�(C?�ܧ����'��5#?�rȾeΌ��''�ҡl?+�@:�@&r?2˒��]ݿ]d��r� ����gJ>}��=��=o�OJ>���=�F��tԫ�.
>3D�>�w`>"x>�;>C�>�h>?'��B+�I��䛏�_*�[71��k'��[O��"žk ����qu������C�� Žʹ̻#�#���gg��c1K><:R?KP?�?�+,?Y}�>{:i>{]�ᎀ>���=�G>>Rs?Z��?A� ?�=�a�����"�������vT�)��>��=>�ĳ>x(�>�b�=Yp����$>��w>TJ">��=
P>�������N>��=�ؒ>$'�>�C<>��>Eϴ��1��f�h��
w�Q̽/�?z���Q�J��1���9��ͦ���h�=Ib.?|>���?пe����2H?%���})���+���>{�0?�cW?%�>��S�T�9:>@����j�9`>�+ �vl���)��%Q>xl?�f>c]u>J�3�D8�֞P��N����|>�6?aܶ� �9���u�[�H��6ݾq�M>�þ>��F�td�����I*�Q�i��*{=��:?[�?����̰���u�T&���pR>��[>�9=Tg�=�hM>�{b�ǽN�G�Q�.=j��=ͩ^>�?��/>Pϛ=5R�>�����jI�0>�>��@>� >u�>?&�%?6�*�~���^���x1��Nm>�E�>$C~>�>��H���=1k�>Md>���7������?��CU>~���J�^��A��GB�=%�����=�U�=k�
�߇B���@=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>B���藿������t��T9
u�>"mI?s���Pu�{�<�|?7: ?Z��i���ȿ�y�5��>��?��?Q�g������g>�+�>M��?&�W?Y&h>'�Ծ.;p�z��>r9?AL?�l�>:F�j}1��?���?b�?��O>y.�?y?��>�ֽ-[�����4䇿a���Nx;��>��=�Ȫ��TA��ɑ��r���h�%)��X>O�Y=\�> _���6����Y=[���(����Qz�>�>�F>lŐ>���>�&�>���>�p=H�� ؈��d_�C�S?��?�T9�2�i�p��>��>�` ���>�'?<zý����>��>�Q?��?�/S?�= V ��d��t<��?���&=��7�>'�0?�P�>�D����>��������L�����>B���J�����ؙ���>� :?H �>�J�B�-?t�%?�)�>���>�\��͇���!��?�EQ>�C$?�?h��>X�3��6��G���>���h���=���?�&?�Џ>C��P!��ՀD>3��u_L>�0�?�|f?�2���>���?Jk??;�B?��>�6���v�a�9=l��>"B!?C��vB��~%�0��E`	?.2?���>rhn�KMҽPؕ���+��}/?�^?��%?���s2_��f��@�<�~�"7��{B<ں���D>�>�/|�lK�=y>Gާ=��n���8��,k<�f�=��>^��=�P4��L��$o*?�Hs��'����=L(~���D��^�>�=����<c?'ž�b������E��6ŧ�m=�?.��?���?P^I�gj�Ɋ=?�j�?�l?a�>�]r����6Mݾ4�8�Թw�0���)W>c��>�!Y��5��?���X���8|�3��^%�R��>���>�I	?g��>�k>&��>�z���*� ۾W�Ń^� ����6��/%�te��ɕ�PB$��.��E��~	�����>�9/�(7�>��?�c>�m�>�!�>�ʀ���>�.>�>ܴ>4�]>�}>�=k6L�.���]JR?	���(�'����骰�,4B?Gsd?�0�>��h���������?���?�r�?2Kv>Dzh�f++��k?�9�>��qo
? :=�p��f�<U��������_�����>�A׽i :�	M��ff��k
?).?���T�̾,׽�s˾A��<t?5)?< )�n�P���k�^3T�]J�Q_�=g�����^����n��搿�J���0��-#�r@C>l�,?K�{?Q�۾��Ѿ!訾?�x�w[-���>.��>�}>���>'"�>c���t]O�
o+�_���)�>|p?ԍ>#vI?ì;?�Q?:�L?���>˘�>���_e�>��-;�/�>���>б9?�y.?Z�/?h�?b*?�]>a�����w,ؾ�?f�?��?:?3�?*^��f����U���:M���x�x~y����=B/�<?�ֽ,�y���O={-U>�Q?E���8�Ϭ����k>ą7?���>5 �>΋������;�<g�>
�
?���>!S���Kr��V��;�>匂?}�ma=�)>���=W<��0c�����=\꿼�=�܁���;���<�%�=G�=<�i�4�� ��: D�;�m�<��>fEh?o0�>S𹾓lܾM���BM8�i��<���>熑=�>p>7] �!y���y��)UP��Wz>�n�?�ǩ?t��!�=��D=������}j��ʇ���qj=J)�>� F?�~~?�Ho?�BI?Һ?�D>cRϾ��w���B�$��k!?H!,?���>����ʾ��ш3��?[?6=a����:)���¾��Խ0�>�[/��/~�m��D����c���}����?���?�A���6��x辔����[����C?d!�>�V�>��>��)�	�g��$��,;>��>�R?Oܻ>S�O?+;{?�|\?PW>�;6�=D��%9��� $�"F>}�??I�?�E�?.�y?���>��>a�-�o4����U�!�����Ɓ�w�E=��V>儒>W��>�l�>�]�=wʽ�����<��ǫ=a|b>Y?�>%`�>��>v>��<��G?�?�>�������k�����?�`nu?%|�?�D+?w=����F�l�����>�\�?���?Y*?:T�ur�=��м5ƶ���r�>߷>n�>0k�>ܜ�=}XH=w�>��>���>���Q��f8�;iN�'�?1�E?�H�=�ſ�i�ib� ���򹕼�x� ⍾�D)���p�+�W>�d���ǽ�����鈾V���0����O����Ҽ��?��< ��=ڟ�;���;7�
��9w=�5>����?��<�\����>�[�8�a>ĩ���Y���}�6�r='�6�J�˾�}?<I?��+?+�C?��y>�9>��3�噖>*���<@?�V>$kP������;�����J#��5�ؾ|׾J�c��ʟ��K>�DI���>�63>p?�=� �<L�=�Hs=ώ=x1R��=i�=�N�=-e�=���=n�>}X>�Cr?/|~�`2��F_��=��"?�_�>:����N�&?rq��13��C4¿����i?���?$g�?-�?a[� �>�����>��=8|[�?=�{�=o�\��j�>V�>	�s�,����f >�0�?d@�w<?�����࿇�{>�7>m�>*�R���1���\��Bb�ڎZ�N~!?82;��]̾�@�>�:�=�J߾�ƾY3.=��6>Yld=T��yK\�Ž�=�z�-�;=A2j=���>��C>r��=iU���ȷ=@�J=J?�=f�O>F_��%p7���,�@3=���=Vib>##&>:�>�s?�0?�$d?��>#k���ξ����뵌>���=��>��=��C>a��>��7?�hD?��K?ұ>s��=r!�>��>� -��m��u�x���s_�<\Y�?!n�?*q�>��<�A����->��L����?h1?	?޲�>	#�|��baw�'���'
>�����7A=	!	��b��1�$�Î���I��tY>
�D>!i�>*�>Ic>j�1=�Eo>���>^��=�m�=�*�=J?<�퉽$A�=��=�B�%��=̟���v�<����lѽ��<G=�M���=kg�=��>���>߷�>�`���q�o�=�G�(J[���(>� �#�-�q�Z���q�3�������Ċ>'X>¯v��(���n�>�(�=6�>���?��?�Y�킙�4g���s��/�̽s�{�P"C>%��=툆�^`���n��J��ľ+��>j�>��>$�l>�,��?�vw=F��Xx5�p�>AE���$���� ,q��:������`�h�&/غ��D?	>����=D*~?�I?�ӏ?ܩ�>�����ؾ��/>z���=C*���p��Ⓗj�?M '?�?�>;��D�먾�҂!��w�>�����_�l3���N�棵=��ƾ��>�ǳ�a\�?7�&i����bx^�h0���>�y?3ɮ?���ߧW��)D����%�=�a?J�#?v��>���>��>�h\������ƾ�"4��3s?;��?��?۽C��=�䩽�[�>�o�>�?z�?Mz?^R����>P�����>�@�=��i>'x>&�C>�K,>]�>%`�>���>�伃�	�u�9��J(���������=>���>�p>/�>p�>mߟ=|~<��o>�=�>S�>�u>O�?+A�>�i��R��=�6?�( >��>��E?m��=�=d����=R�o�Xχ��|��Խ��3��-1<�N�<ñJ=S��@�>�����#{?�x>�˾v`?�%-���!>�K�>EJ�=�����̱>V�>���>�E�>{�\>X>h]�>|A>B\��y��;����"�_�4��4��р˾��>Ǿ�=�޾Q�:>^jl����|
'�{mp�D���#�tV�>3B�?(����U���'���q�̾�>4��>��K?�W���"���=ѯ�>`yS>�ö��������w�̾o��?�G�?�[w>�&�>��V?�V0?�B�����"���A@!�'/(�����N�%���9m��!��:����L?�At?��j?��H�z�r>�ߨ?�d�=�ܾ��>\c(�%mƾz��=��=��¾F�E=.I���A?�u��&�C=�*^?�j?f�7?�q�;�<\��=�j�>�-?���?#+?�H? �9=��>?�Ad>��?�B�>!*'?5D?�BF?�B:>W��=�K�;*i:�`D����r��L�;BM�b�4�c�� �<?=��-�����=�-=��f��郼if�<�e���`g�:�<=�p>���=7g�>�xb?�W�>_f>��,?�4���8�	.���S*?k+�<��x�����J���S�!6�=��g?>O�?�r]?��R>:�@�;O6�3�>c�q>��>a�Z>�&�>|���'���=\�>�&>�i�=��D��p��k��:+�� }�;u$>��>��3>5��=!L>H׾{�~����>���f߾����$r��}2�r/���X�>�M?�R8?�0>�ž���co���,?��=?��,?��y?��\>?��`3���2��?S�{��>�r.>�%�8��������[�V��og>b���ޠ��Xb>4���t޾�n��J�G�羾CM=���ZV=^�3�վ	5���=�%
>��� � �4���֪�\1J?Ϥj=)x���aU�ip����>�>�߮>d�:���v���@�����5�=��>O�:>�\�����~G��8��s�>'�E?�\_?G\�?)���ַq���B��������T�ռ��?Rԧ>d�	?tH?>��=�=��A���7d��C���>t�>�� G�1���+x����$�9b�>0�?{�>�?�{S?��	?q�`?�+?�#?�}�>���(���A&?>��?��=m�Խ��T�v 9�SF����>Z�)?��B�E��>N�?�?��&?��Q?{�?%�>� ��C@����>�Y�>��W��b����_>��J?���>-=Y?�ԃ?>�=>P�5��颾ש��W�=�>m�2?�5#?�?m��>���>ۮ���=���>Xc?�/�?B�o?I��=��?C2>���>��=���>��>�?cXO?3�s?�J?��>$ɍ<�2��S���]s��xO�?�;M�H<8�y=���/t�9����<�ڴ;?p��/���e�	�D�h���"k�;YH�>�8s>����o�0>ž㈾$�?>����F!��A���W�:��Ŷ=�G�>#�?�ŕ>�;#�)�=,��>\i�>$��R7(?��?-?1V?:>�b�L�ھ;MK��z�>g3B?��=��l�������u���i=�
n?E�^?�V������S?��?!0�*B��#��]6��l�%T7?�{�>�ᓾ�>?Z��?GKp?Nk"?IV^=�X��}`���c��=����<(�>T�¤��z��>�D?��>����U�=�k��*�s�B�|�s��>��?�"�?�?ʑq>�t���=�t	��a4��x�]?h��>�����"?_���Ͼ�؊����:o�>誾Y������xP����#�����z�ֽ�~�=�?'`s?j<q?']_?�� ���d�u%^����JV�n��h��̱E�c�E��D��Go��@������k���
S=M�r�<�F����?S5?�5)��	?�6ʾ�Z����ǾK�=I毾�%X�t�==vx���=r�=��R��) ������&?|"�>���>r7?�����$D�Q���$��I��Oב>�L�>�ݥ>Gt�>$�|���p¼�9��D�;������7v>�xc?��K?۸n?to��(1�ƅ��k�!���/�(b��m�B>K`>�>F�W�R���:&��Y>�Y�r����av����	�	�~=��2?H%�>屜>>N�?H?*z	��n���ax�6�1�,��<�.�>i?�<�>��>m�Ͻ�� ��>x_?��?���>����$��2U����Ҟ�>=�?gb�>%H�=z���4@��E��8Y��8;=�L,-=�E|?�A��
ؼgk�>"<?���=���=�>���=@I��k%���]�B·�֪!?�Y�<jB�=R¾��!�(�w�Q��J)?5X?�����*�,�~>&"?2z�>�>n#�?4�>�ZþD�6��?��^?�CJ?�CA?4!�>�C=�W���ZȽb<'���-=���>t�Z>�m=Av�=0L�-V\��� jE=rG�=��ϼ�}��cL<������K<��<�4>�ٿ7�F�`A�w��?Ⱦ��
�7����s��">X�pJ�5оW���Q�w��˃Q�(T��FV�=�z���C���?:��?�m�����i��6t��.����>��>��/�<�����p�y���������Y@�"�H�n)�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >YC�<	-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾w1�<��?7�-?��>Ŏr�1�ɿc���{¤<���?0�@BA?�(�
���U=K��>y�	?+�?>�>1��C��𰾇Z�>�<�??��?�M=I�W�9�	���e?��<��F�G޻�!�=��=-="����J>�P�>i�AA��Eܽ��4>��>*8"�|��R�^�丽<�u]>8�ս�(��5Մ?,{\��f���/��T��U>��T?�*�>@:�=��,?Z7H�a}Ͽ�\��*a?�0�?���?&�(?8ۿ��ؚ>��ܾ��M?aD6?���>�d&��t�؅�=�6�։��y���&V�{��=]��>e�>��,������O��I��T��=Q��¿�68�%���=�6�=�w��2#�L�~�3�	���о%�� h|�T�D>���>�q>�NS>��9>���=[�a?FA�?�_�>A��=󶃽���e�侞��<ڽh���������#�
c�HU&�K�	�ξP���w?澸ge��=�؍=�AR������� �`�b���F���.?^(%>��ʾ+�M��9<n�ʾ� ���f�������̾@Q1�\�m�}ʟ?�A?"�����V���P_�s��n�W?'� ���t���?�=B��F�=��>o�=z~�I�2��[S�
=?�?�Xƾ���+<ˎѽ��>+0??Kh8?�$:>fc?`�V?�����2�ٺ=�(0=��>��>�>�>þ�(��r�,?�K?2qw��;ub>�f���tȽ���>E|�=)2����=䯮>�P�oپ�D�n���3$=PJc?��R>O0��x��s��F:=C->^�?�
?���> tv?�P`?3��e�TRP��"D>>�	\?��I?�=����8L۾�P��>?1?WK?�>�'U�uR��0�"�񭏾��-?�xi?�/0?kb@�����ț��ih�&�/?��i?eJ�,��� ܾɋL���>$(�>��?e7E��1�>�:?%"�����`��,�-�(�?o�@S��?SG�<+";u��q�?y?��3�z����=�&�C��~��>�L׾<�����
��G���DA?�?�q	?l����辬��=p��\�?.�?~Ѫ���d<m���l������ţ<��=���+$� ����7�xƾ��
�pv���Y_�>L@�
�r��>��7���&gϿ�녿.�Ͼp�q��?�~�>gWǽ����/�j��{u�?�G�k�H�4w���[�>�p>�O���ɑ���{��@;��n�����>?�8�>��S�"!��k����u1<� �>��>��>���\���+ř?�'��s-ο���l��ҔX?�o�?2g�?�x?(D<��v��{��7�}�F?�ps?�+Z?��!��C\�g�8��j?xW��*K`���4�JPE�B�T>_$3?7C�>Ym-�~f~=h>G��>h>N/��Ŀض�/���p��?s�?Ex꾛��>e��?�t+?�m�8��tU����*���@�2LA?��1>���c�!��=��ג��
?�c0?��C#�]�_?+�a�M�p���-���ƽ�ۡ>��0�f\�:N�����Xe����@y����?N^�?i�?ӵ�� #�g6%?�>e����8Ǿ��<���>�(�>*N>lH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�K�>|��?&9�=���>Qq�=�E��Z���">�W�=(�=���?MM?�Q�>H��=��7���.��#F�ZR��q���C�Y^�>�/b?��L?Uga>�Ӹ��1��� ���Ͻ�1��x��$B�65,��v߽�
5>�Z>>�->�<D���Ѿo�?˳�Y�׿�)���(��?��R>&.
?���E[�o_H��e?h�\>���ó������z_�?���?�J?�SԾ59���>�N�>�[y>������8�EN���#>�C?�^������j�B�>���?tT@'�?��g��o�>O����*�����ʾ	u�������`?�	�� &q>�f�>��>J�����)�w���>n�?���?V��>/�c?R5I�����Z�>�{\>�Q?R|-?g1�<h#���8=��?�N�uv�����\?e��? �
@��`?�ě��8ҿ(���6���l&����>��<��Q>E����TP=L��Ǻ�<�*B���>|��>쏃>_{p>@IC>��B>�{>������)����u���C�D���#�7��QT����8��c�����B=��� �r���v���?!D�0t�@0Y����=�M?�7?¯g?��B?�cR><��>����ܼ����ن�=�^���7?@LU?F6A?H,>f{վ���01��{�����eN�>%I�>���>G˨>D�>γI���>ѱ�>N�>�:�e��=���P�0���6>��n>�"�>7�>�C<>��>Eϴ��1��c�h��
w�f̽.�?���T�J��1���9��ͦ��i�=Hb.?|>���?пg����2H?.���v)�߹+���>|�0?�cW?-�>����T�::>6����j�.`>�+ �pl���)��%Q>wl?\�f>�Fu>��3�+W8�A�P�N��Rv|>�+6?b߶�I�9���u���H�=ݾ�~M>y�>94B�@i������ ���i�xz=݄:?��?iv��Dְ�Qtu����=MR>C>\>�G=Cɪ=�2M>/�c�Joƽ��G�C�-=��=��^>R�
?�s>�ߛ=ò�>z�þ�np�H�>��+>�_�>�*`?�#2?��<}h_�k���]���>��>�ʃ>�� >:�w�h��=|�?z��>�m9�2�ｫ��a����`�=�L<�	��`���d�=�ԼAˎ=�G?=�KR���]��ײ=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿe�>Ax��Z��.��M�u��x#=���>9H?&P��?�O��>�Vx
?L?�`�/���K�ȿ�zv����>��?���?.�m�`A��
@�	��>k��?�eY?�wi>�f۾g_Z�6��>��@?QR?'�>�7��'���?�޶?{��?��D>�b�?�N{?��>�Fý�} ��F���u�]����	=��>���<S�����@�����Gq��d:o�w���>9*2=s��>=���o����v=�9���a��Zi�=
��>r�=:*�>�Q�>�?�S�>;P�>Ó��Y��wTP�V魾�.5?^u�?���j脿�(�>m�<>D텽��">�9�>9�H��ѣ��s>�4Y?���?8�j?�k>�0�~���t�Ͽ>���-�~�Hc>E�?�O�>��/�!aQ>��O�<d��bl=Һ�=��_������d��L_����>)�5?j��>�����?w7?�$�>���>��5��S��a6J���?�b�> �>ON�?��>E��������꫿��y���
>.�v?@�?!ݝ>�����Փ�S�=u�b��a4q?�Tg?)�����?C��?�?�/Q?2��>	������t��<ii�=��!?>|�ݳA�1x&�^����?B?�@�>5l��M$׽�/ռt������ *?B\?=&?����^a�J�þ(�<�/��uN��<�JD���>��>>����a�=��>J��=\�m�O6��ua<{��=���>3e�=�	7��Ϗ�?'��'p��C�>��v�̾7�^��>h��;��?K?�辣�������܉�B �ل�?n�?X��?O�ۻ�PX�c�>x��?�i�>㭄>��ýU�����ڽ����GI��j�=�?J�=����\%��"ء�U�~�_r�%<,��`�>�c�>Dj?�?[�>Y�>�N��b3-�"��W��g��H
�nn-���2�����N��il)�M��IA��¿���x>���f�>6�(?{*N>�#v>k'�>���-�>��">G+�>��>o;G>�A�="B�<ݪ=�F��KR?�����'����_3B?�qd?�0�>�i�-������v�?���?Ws�?�>v>�~h��,+��m?�=�>L��q
?mU:=�:�M:�<�U��\��M3����
��>�F׽� :�yM�nf�lj
?�/?`��ȋ̾$?׽ B����E=��x?�4?���/�X��l�tIP�4�B�����]���1���'�x;p��^��/�x�h�}�����=դ0?�X�?O���ٍ��dB��֎x���B�A�x> 0�>)��>��>�TZ>u�JF=��l�H�)�f:���>�>�?8�>�zI?[�;?KP?yL?��>U��>�����>@�?;Ԥ�>O3�>�i9?�.?U�0?�L?T*?�y]>K��e��~ؾǊ?e?E�?k{?��?ʅ�6½-��T2t�|�|��%���=���<ӌֽ�t|�G�[=�6T>W_?t����8����(�j>F|7?���>��>h쏾���݉�<#=�>&�
?Q+�>v ��ur�fR�r[�>w��?�P�Y�=�)>T�=1��c�ۺ+7�=������=)�����:��F <ӵ�=*k�=��r�+�E6�:ǂ;Q
�<�Y?&�?ur>��`>b���fwᾳ�Ⱦ�٭=��e>T�>nX+>ݯ�/���Ę����X���>�ݑ?oP�?��= ��=�4>�󾫺۾N�ξ���y̹<�?��?)8?��?LL?�0-?8>� ����k���ұ��?�",?Ʌ�>M��\�ʾ󨿪�3�O�?�S?�"a��K�))�{¾b�Խ��>�]/�r2~�f���D�ޅ����aZ�����?@��?�&A���6��t�����eq���C?��>�7�>3�>�)���g�S!�,�:>Ev�>R?�#�>��O?�<{?��[?�gT>�8�J1���ә�WY3���!>@?���?�?$y?�s�>��>G�)�A྾S��P��p�6Ⴞ�W=�Z>N��>V(�>��>���=�Ƚ�X���>��b�=`�b>��>��>�>�w>�F�<�#Q?���>q�.���վsz�-�ڽ'�z=�(Q?�U�?QW;?(C���"�yO�Q�!�=�>lt�?�ϰ?.~E?���I>%I�����i��Cg�>�:>�v�>ʕ�=�v#�W�J>��>���>����\+��l=�������>��U?稼Ŧſt�q�Y@o�����Ӆ<�A��%�h��ѕ�9C[�ޝ=<����-�����݊[��r���̓�,���! ��L�y� ��>A�=,M�=?4�=Y2�<���HҸ<هN=Hu�<9=s.g� k}<=��<{�h��T���uV<^NQ=����˾4�}?(8I?2�+?��C?/�y>מ>�6����>�����3?Y�U>XcO��^���R;����p%����ؾ�׾��c��ɟ��>/FI�j�>�E3>���=��<jO�=G�r=���==aE�3)=���=�-�=b�=�1�=�>�[>83r?&�z�#��xM;��h
�Ѻ#?�J�>� �=WR��6?�m4>�|���H������s?\X�?ӧ�?s?d�N�r��>WJ���9C<tp>�`�T�^>�K>���^<�>%\>C-�|P��o�¼��?fA @�vB?w"��2�ҿ��:>.�7>z>��R��1�B�\�f�b�T`Z�Т!?7;�/3̾�G�>=K,߾m�ƾA�-=w�6>p�b=�?��K\��ٙ=�z�r�;=l=xՉ>��C>h�=lï�K%�=�eI=�*�=��O>���#7��,��J3=Ͼ�=��b>]&>���>�X�>>�F?ǡY?U>OEֽ�Bh��sʹ>��=��m>�"�<}��=R�>��7?m�>?�P?vM�>C6>R��>4�>D���NH���h	���V>�~�?N(�?�
�>��,=����(��[`�	�p��,?�	X?�c.? ac>G��I��GR�e,�� ��M�=��.>�?��Y=6�u�O�@��K���·>8�?TB�>�{p>OR;>.�1>->H��>�W.>��\=���=�S���׋=�5�x����Z=�@�=���5�=�X��R���� >�@�=�+=��������E�=���>��>�@�>��"���������𲾹�L���=�>���"B���O�ѻj��] ����Wu�>E2>I�<A����_�>
�=B����?S��?}O��9P�N����,��M�ɽ+M\��Qn>�2�=qۃ��|\�ed��HK��ڵ�H:�>T�>;��>�;�>B82��?���=�_�?"���?��X�+n���C�ٝd��R�����b��'�:~vC?�z���%>몀?�I?oU�?�h�>����Ԩξ�d�<8�����''�d78��ʎ��?^w"?�^�>�������p۾Tν?�'>V�Ⱦ��&��𡿲WL�s�=���UC�>�ʪ�ӥY�n#J�w����k��n}"���Q�d��>�[a?�U�?�2���x�HCF���((��ڱ>��o?}R�>��>P�?\�>e������p=y�B?׬�?���?�q>���=�W��|�>p 	?ʾ�?�֑?	�r?u�?���>�P;+>nl���=]�>"�=|��=�K?xh
?�
?p霽@�	��_���񾕢^����<h��=�k�>T��>%�r>�F�=�g=$p�=kU]>�]�>
ԏ>*cd>�%�>�Ɖ>hL��X����.?��=��>-�L?�#�=%RO;�X	��ս��
�+<����"�R�g��� �+f��T���b9:=M0�<Y�>ѱ��f
�?+7>l���?y�ܾ
�Ҽ��>�\�>��!��W�>��=��><��>s+�>�>�c�>�Ln>V�־S�>,�@8"��f@���T��Ӿ�aw>�3���T �t	�x"��P�����[���!g����f:���=�i�?�?�vj���*��2�?�E�>&66?X����o���>tz�>��>�T��}?��텍�J�߾U0�?�]�?��^>S�>��\?B?��V���1���X�8�t�~�C�&CX��|j��������RH	�˸���_?�Kx?��=?��=��a>�?�)�Z���1�>�F%�BH��T�=�ȸ>&����nE��Iƾ-��%��B6>yX?C|?H?��F��Qq��E,>�c:?Rg3?^w?��2?|�=?h}&���"?�1>z�?�I?06?�.?V�
?�5>^
�=�ڢ�;7�<����銾�ڽ�wȽ�@���^A=��=vo��P�]<�=�G�<ת���>��<��<!����<9T=���=���=>��>�]?	R�>���>t�7?���Uy8�4Ȯ��&/?"�9=궂���~ˢ��x�>��j?���?�bZ?@ed>q�A��C��>(N�>�&>2\>�X�>Tk�7�E��=�T>sW>�ݥ=fM��с�=�	�Ō����<�#>U��>��z>�
*>�C���z�l�c>|[S�M���"vR�T{H�,�1��w����>"�K?� ?ᱜ=��[��� *f�R1)?e-<?YL?��?��=�ݾ3P9�-�I�����>�X�<O��z����^;�%�8YXr>����ޠ��Wb>A���t޾+�n��J���羥DM=���ZV=_���վ�4�ڤ�=%
>����� �)���֪�p1J?H�j=�w���aU�Mp���>>�߮>4�:�u�v�y�@����45�=��>[ ;>\��*���~G��8��~�>`I?:�S?x�|?�,u�+�i�%	7��辞��_8彊W?:c�>�,?�wL>Va<�N�F�%�ݗX�mL+�Q��>,6�>Y,��B�?@���_���Q2�Y�>��?C7I>�,?Qq`?��?�`?�;?	?��>�L�ۛ۾2B&?q��?w�=H�Խ��T� 9��F�|�>,�)?9�B����>e�?3�?'�&?K�Q?��?��>"� ��A@����>�Y�>{�W��a��[�_>��J?}��>^<Y?�ԃ?@�=>]�5��梾�����e�=g>��2?l3#?��?���>��>����ܮ�=��>��s?�ی?��|?]s�=J�>2v>��>��)=h_�>V��>0�?�J?�bn?E�;?L��>���<�Z��du���Žr���և(�񛸼��=i���^��施eE=	^=z����J��dG��gG���ȼW�U��^�>E�s>6ҕ��Y1>i ž�&����@>h禼8��Ŋ���:����=�|�>G�?=��>{l#�ۚ�=7��>uG�>����,(?a�?u?�	�:��b�"�ھ��K��@�>B?޳�=*�l�-}��g�u��h=�n?^?�AW�+��T`o?-�m?��]>�0���֒�4�;�wl?'5�>�Ɨ��&?Ï?���?)�,?��5�Ŭv����PuX��ۥ��>�I�>�1'�}u|�Q|�>:K?��>VBU=.3>��U�E X�:����>�>�?9�?�-�?��d>튿�M�ɪ��o]��7zZ?�f�>�3��q`!?&�C���Ͼ+����P����+~������㓾�����["� %����ٽ�$�=�?.�u?b�q?Š^?):��Nf���_�ĭ}���S��H���Y��vG�ΠG�8E���p�mJ�?��A͔�~�a=(�J�XZ3��t�?��5?"&K��,?��ƾ�7�{�[0	>���;>����<�4�{�&���ǽ���%D���O��M$?�d�>-Ύ>�{G?�掿>�1��2�Ƚ%�AY�!�P>Ʀ>0s�>��>�U��s�ᔥ��Ս��'Ͻ�Њ�f�v>ˆc?}tK?��n?v)���0�^0���v!�5��]��!qB>O>�
�>��W�5���k&�Y�>���r��`�ȇ����	�-�{=Ō2?��>�A�>=Q�?�?��	��°��x�Ls1�gE�<|��>�h?��>�9�>�ҽ�] ����>��v?z��>艈>�/��a�:�R�~m�:7�>b�>> ?���>|�����G�왁�����6��z�=�C[?F/��);z���>'_?U��=��=5�?�w��~�0*��7��y����g?=Ѐ>u�=���+��z��`�P)?eF?iؒ�g�*��~>�;"?Q��>�>�(�?c�>oþkiG���?��^?x>J?�OA?�L�>�%=�S��7Ƚ��&��Y-=e~�>��Z>�l=�Z�=���!�\�h|��D=Td�=��μ�c����	<�L�� N<��<��3>��ҿ�O��3������׾���y����ƽ�S���3�^�ھ���ؠ��� �Q<O�7�:�K��*���|_�,i�?��?�V��ln��7�����#Z�>�`�� >�v��DJ�ޥ羐{������!�� N�s>�+�.�A�'?�����ǿ氡��:ܾ.! ?�A ?*�y?��;�"���8�)� >E�<�,����뾯����οL�����^?���>��/��j��>祂>
�X>�Hq>����螾�.�<��?#�-?��>��r�*�ɿ`�����<���?+�@u|A?�(���}+V=���>��	?��?>�T1��J�J ���R�>=;�?���?�|M=,�W�	
�|{e?�*<��F��ݻ��=E6�=�<=����J>�S�>���WA��]ܽ��4>BՅ>@m"���?�^��<��]>��ս�,��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=�y��>2Ŀ}H��&"�z�=��=���U������;� �NEȾ�|��Z�d��=�$i>:%H>�*U>���=��8>�&P?�1d?�I�>谍>��D�����~����@��M1�BXB�+�I��Dھa�H���<�����վ|N��;!=���=47R�[���	� �A�b�)�F���.?,w$>��ʾ��M�|�-<pʾ-���L؄�qॽ�-̾�1��!n�U͟?z�A?������V�B��Y�����W?Q����ꬾ$��=(���G�=%�>튢=&�⾡ 3�p~S�`1?/(?�i��q(����>����w�8?$�#?��=���>Gc=?<��h"��f2>.�>�C�>+��>z^ >���y���$9#?#�Q?J�!��U��4o~>�о�=�����=�=?Dv��)��j>߈�80���ӆ�t�ٽa�=�aR?P5�>�P�8^$���t�?�޽�Yɽl~�?�G?d��>I2�?�^w?`e<�-�)�>���ʾ,R�=v�T?�rX?^�=Ȉ�v���O;���m?�XS?e6�=)G�7%��?d��m�մ�>�l?�3?��S�(��bC���y �0F*?�b?N�X�큿�yǾ�վbX�=8?y=�>��0�D�?6>(? �H�ț��9��)^E���?�j@?~�?r{�[ ��۩�=��*?;q�>�'Z�꽬��<�g&����X��>"Q����״.��s��Y?�}x?�y?�'�IN�E��=�ݕ��[�?g�?���S�e<����l�zk���ס<���=I���"�����7���ƾ��
�1����'��ڙ�>�V@&g��>�-8��+�=QϿ)
��aо�\q���?�{�>;BȽ�����j��Uu���G�r�H�����(O�>��>�����䑾��{��n;�S��
�>r����>��S�M(��7����3<$��>��>���>�殽�ݽ�n?�U��>οX������z�X?�e�?o�?wp?7�9<��v��{����&G?�s?�Z?�%��$]���7��j?L_��PU`�Ԏ4�ZHE��U>�"3?�B�>c�-���|=>D��>Wg>�#/�v�Ŀ�ٶ�|���A��?��?�o���>\��?Ws+?�i�8���[����*�Ԝ+��<A?�2>���A�!�0=�BҒ���
?4~0?�z�a.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?*�>��? ��=+c�>5��=kⰾ��)�U#>���=�?��?9�M?NY�>�S�=�9��+/�`F�PER�����C����>��a?EwL?^Ub>�ʸ�e�1��� �d�ͽ��1�	&�7|@�,��+߽2�4>l�=>��>��D�N�Ҿ��?Lp�.�ؿ�i��Tp'�w54?)��> �?����t�+���;_?,z�>�6� ,���%��gB�b��?�G�?@�?��׾S̼�>&�>�I�>h�Խl���Z�����7>.�B?;��D��t�o���>���?�@�ծ?bi�a ?4���p�nY�����Ѿ�#)>0R?�[Ⱦ'H?U�?���=�z�q���.�}���>q��?	x�?S��>Z_?}�c��#��0�=�H>�vd?�c1?����7��I�>���>����'��EZ�1m\?�@@j@�}Z?hX����Կ����I߾v:�F	>L��=˘G>�C�<8�>��r��g3��6=w$�=���>�(�>KO�>��=��=�)i>ڄ��6(�Aw��������I���!�x����.�Ѿ�ya�Z	��湾n��hƽIR�=S��:������$��<�be>9�O?�pQ?�2t?�vC? �>��>ԕ>�L�e�������l;�(>oM?`}�?3�(?�v�<�2�4<s�����p��5���'?��>S��>u�?��>;a���$=9(>c�>�$����#�_c<0ӽ��W=��2>�>��>�B<>�>Hϴ��1��M�h��
w�k̽,�?&���E�J��1���9������Ei�=Hb.?|>���?пQ����2H?���p)�K�+���>b�0?�cW?�>���R�T�Z:>�����j�s_>-, ��l���)��%Q>�l?��f>�/u>��3�Fb8��P��p��\w|>e06?W嶾�X9�s�u���H�tSݾ�\M>�;>4IC�be�
���,��i�w{=i~:?��?0��5䰾=�u��L��~<R>�>\>�=�n�==XM>�c���ƽ�H�ӄ.=���=��^>�B??�*>gB�=���>�E���yS�~��>�;E>�,>��@?v�%?��ً���w��W�/���w>B�>�`�>N�>�)I����=6t�>�b>�7��&����
��CA��U>�����`��w�Ju=������=n��=-~����;���"=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾUh�>9x�xZ�������u�[�#=^��>�8H?�V��v�O�M>��v
?�?�^�ީ����ȿ;|v����>T�?���?^�m��A���@����>2��?�gY?soi>�g۾�`Z����>»@?�R?�>�9���'�w�?�޶?ѯ�?Z]>Á�?/'n?�x�>��>�L&��H������,3��g�� �>��=�񤾦9�����q���"u��s��7�>,{=�#�>���}ߺ�mt=�tｲ���Җ�k̺>�e>�{a>N��>H�>Ś�>���>{�&=���l�I�V����]?R�?̦�(1j��?�>+�>�>�Q��>���>\@v��Cؾi��>/�k?��?Jb�?E�>S���>������+Q��t�н�
�>j�?.��>� �� ��>��P�'������=;�=�y�B ƾ�����wޭ>��<?��>�/]=�"??6(?c�h>���>%�;��؍�P=��>�>fc�>�~�>�}?ߜ	?vl]&��둿"���n�g��&<>�Sw?U�?�H�>ڮ����n�M�����x?/�e?�$���H?��? B?�C?�B�>��ǽ�ξ��f��/>��!?���A�fN&�����?�N?���>�;��0�սOּo��Cx���?*\?'@&?0���-a�þX)�<ֻ"��!U�=�;6$D�O�>!�>���(��=	>ð=FSm��H6�W�f<-p�=���>��=m.7�$����??1{ҽ*=���B>�}��WD��J�>-熽�.Ⱦ�t?���
n���D���!���÷�Yӎ?4��?���?�,�:1O�, ?�?D}	?�?�p��G9ܾk��5��t[�I�$���+>\U�>�c>�k���ő�A⠿B���(�=��9��>�5?^?::?~H�>M�l>v.���MR�����X��c�N�w3���8��a6��徊���x�=cϞ�K����k�>b�<�G�>�;?�]=9TD>�˦>��-��V�>/5>�&>�n>`�>��=�>yض=�f��KR?A���׽'��������2B?qd?�/�>�+i�f���`��;?n��?�r�?�6v>��h��-+�m?�?�>����p
?�L:=jV��5�<9V��|���.����_��>�>׽� :��M��jf��i
?�.?"��ԉ̾)?׽�Ҩ�ɹ<i�q?�"?��&��[�Zfz�?E�$9I��&Ի��z�־�)��i�Fݍ�*�|��x�4��E^�=�5?i�?�\��s{ݾ�A��Q��<�$��>���>���>�O�>��>���9E��|��w�"�:�u��?+�?��>7�I?`�;?�'R?��U?��>��>wd̾���>*���>���>�sB?�"A?��/?]�	?�'?y�>�R\��F����ڮ?�' ?2?�G?V��>�J���N��c���m�;���;���A0�=�w���x���xW=u1�>?�?w�¼o �j�ž�o>�}(?(��>u��>�Ⱦ;������=w��>8�?XU�>>��	G��p�$�)s�>厇?HF��Ɓ.<��>ES%=�I��:����;�O!=J��=��
��Lx=��轐c�=ޛ>t�R����c)g�0�8=�x7=]?�?č>p�i>Ovq�H��H"��`\><�>UT>�ő>[��ue��W��� �J�J@�>��?��?1�=*B�=�,�>�;t���A�R�y�����?��2?G?�m�?��W?s�c?��=�/Ᾰȍ�s��;hݾ� ?v!,?��>�����ʾ��Ɖ3�ޝ?_[?�<a�T���;)�Ӑ¾{�Խ�>�[/�n/~����?D�k녻������-��?忝?9A�M�6��x�Կ���[��f�C?"�>�X�>��>=�)�x�g�x%��1;>���>hR?>$�>J�O?]<{?x�[?�qT>��8�t.���ә���3�=�!>;@?N��?��?Vy?�q�>��>�)�}��R������߂�OW=OZ>���>y&�>��>��=ZȽ�U��8�>��T�=�b>���>��>���>#�w>�x�<�C?|��>���f��'~��׮��짽��x?
Ë?�r?|{!>6�#�Z�ms�ڐ�>�x�?�/�?'16?6d:�!#�=�I>HT��ž���>D��>�uZ>W�'>�γ=W��=}��>�?k潵� �F7�\r��|i?��7?&�!=lkſ�{��}���#��+��=X�|��wO��q<������<�����k��u��qC��`�����-	˾]ׯ��s �m��>+��<d��=E>��'=C+���&J=�m�;�;�O�|��K����>=���<4� �r��˯�<�=�S=ހ-=�˾8�}?8=I?p�+?i�C?�y>�6>��3���>ɂ���<?�V>ʫP����0�;���%��:�ؾEr׾��c�3˟�K>�]I�_�>�H3>5�=�N�<��=��r=WƎ==�Q��=$�=;a�=�c�=��=��>/I>�6w?X���
����4Q��Z罢�:?�8�>O{�=��ƾr@?r�>>�2������zb��-?���?�T�?A�?Cti��d�>K��w㎽�q�=;����=2>n��=��2�T��>��J>���K��B����4�?��@��??�ዿϢϿ6a/>�7>!>��R�ˉ1���\�>�b�|Z���!?RH;��I̾�7�>�
�=�+߾$�ƾ��.=�6>�bb=�g�JU\�'�=0�z���;=M	l=�։>��C>|w�=�2��,�=b�I=,��=$�O>C���7��',���3=Y��=�b>�&>�Q�>`�?�0?4�i?��>u�uȾ�ݪ���>ms�=ד�> �=B��=�(�>��/?)�Q?gnK?���>��=/f�>D�>k3�t z�ν��o���-�Ս�?"�?惒>y��=��Ͻ��"�@�<���[?�{4?�?t�>����!ӿ%�v�x�t�d��:���=g�Y>c��=7�]=`yq�E4����яx>`��>5�!?���>g�=L�1.r>p��>(��;{o��E��=�.��n��G	�J
�<>���Yμ�����ݽh��<bm�=�t=<5{��>���=��!�)N�=��>R��>��>��<�x̾��B>�?��O)N��I�>q�˾�Q6�ʁW��f�o?��0k�ة�=S�]>I��=꬇���?M�>sf�=�W�?'��?Z
���1�����񛿵Ǐ�Ə����I>��D>��S�7(^�����+j���m����>ˎ>�N�>(�l>��+�� ?�ԟw=�M�Z�5��
�>������?�iq�>��:���ui�Z>ۺ��D?�8��o��=��}?��I?4�?��>�ᙽ�ؾ(�/>���nW=
�fq�����R�?�&?�A�>��뾱�D��?����U��>
���ce�����3G���=�s���?�A�^*Ͼ�M�Z���}�����1�ԧ�Ӕ�>�F?'��?�km�
#D�����*��]I�$�!?/te?q�>5�C?@�?l@ >�=žwś���-=��b?�[�?�\�?$�=���=�"����>��?i�?_Ô?y�w?��=��x�>��Y�$� >��=�N>ē�=y	�=�v?B�?�
?��.���,���{Gh�����[=LE�>�P�>y_{>ε�=᎙=\W�=��^>�C�>�$�>!�e>�&�>e3�>f�;�
�~/?�	>�+�>>�6?�\>��m<le��ɂ<Yꃽ�zQ�7�<�W̽�����o��M��Y�m=<Ө�])�>(�¿a`�?wg>�f�k�?L���z�/$s>��<>�蝽q��>M�E>�3>T��>�I�>/�*>k�>��>�NӾ]S>P��R!�}#C��R���Ѿ�}z>u�����%�x��i���LxI�Ks���p���i��&���*=�` �<?H�?����a�k���)�����B\?�*�>�6?����>f��(>_�>�x�>Wy�������Í�]]���?��?�>Q`]>]X?&�T?%�	�=�ܽ!R7� io�(�ܾ:|���<��׈�E�x�0:)�9c��q?h�\?��V?�l�=�eq>J'r?f7��̟��g�>x�X�(O	��C�>>R�>ib���X<�Ƞ��%��_ҽ�o�>��?�}?Z}?�������r�>��1?��-?���?��W?�MU?��I�_�?�C>/��>�� ?
�8?6�7?1?eC>�q>]c]�lLP=�d�%�e��4T�ͼ�; ��1=�=�j�����!⻄���Zⅼ�x��l�7��4ɽ�F=�'�=��==gڦ>��]?��>,S�>ݰ7?�1���8��8��ee/?��:=i���`���Ţ�Q��>��j?��?�hZ?�td>��A�`�B�
�>��>S,&>�\>q+�>�/�6E���=�C>Ho>��=��J��ā��	��������<�T>���>*D|>-����'>�i���z�s�d>��Q��Ⱥ�[	T�T�G�S�1�ijv�c�>��K?��?d��=�f��y���Ff�+%)?�c<?�OM?r�?���=`�۾T�9�_�J�[.��#�>{Ȫ<��������!����:��h�:z�s>#��:���na>M��v�޾�Xn�/�I���tN=l���U=���վ�'�ُ�=�	>����;� �����v���-J?��g=�s���xT��[���1>��>�Q�>��9�.]y�2�@��ାE�=���>�;>k4��=�HG��$�nN�>LWE?0V_?f�?�#����r��B�f���k��V�ɼ��?�{�>�p?�.B>��=wͱ���%�d��G���>��>~����G�d9���/���$��x�>E9?��> �?z�R?��
?.�`?>*?)C?�/�>�䷽�긾�A&?8��?�=J�Խ�T�} 9�@F�i��>o�)?A�B�ܹ�>M�?�?�&?�Q?ݵ?[�>� ��C@����>�Y�>��W��b�� �_>��J?ݚ�>d=Y?�ԃ?o�=>^�5��颾i֩��U�=�>��2?6#?B�?�>b�>�ȡ��5Z����>\	�?W�?�c�?M؈="�?�a>s�?��>vS�>Jp!?G=?��2?�%H?'�?�0�>�=To;����c�i��ί�!�!<��>j�$��y�ׯw��޿=�SN=����U�=��=v
=I��ź[��+�>�s>x7����0>��ľ����9@>�j���^�������,;�%�=$6�>��?��>��"����=ϸ�>�9�>;��!n(?~�?f�?0�:L�b�۾-~K�˶�>��A?Ω�=�l�����20v��sf=N�m?��^?��V�(0���1o?e�l?!�^6� sܾa�����о��]?'��>*X�� ��>��?�d|?�?�1���v������U�����=K�>M�-��2?�U��>��'?�]�>�*�=��=C=���YQ�В+�!�>�3�?H��?q��?ž=����ݿ5����4��j[?�~�>OA���� ??i��.�˾磉�w^������֫�􌫾]���o������G��Иͽ��=��?�s?�#q?yo`?�����e���]��w�F�T�'O�g=�DG�(�E���B�
j�/�K�������L=�Wr��c6�ȶ?�$?(�T�+�>�о���$����u>��;�\�t��=�㟽R.�=Dɞ=��R�����I����&?Ȣ�>u��>�#k?T����>�2 �w8;��޾5H�=AN�>iQ>5��>*�X�I�P<�Z��S&�������v>m�b?UM?q?����x.����n�$��>�n���`�<>�e>�H�>�$Q��!���&��'>�Tt�V���Q���%�JbX=�1?��>�+�>�`�?н?.2��h��M�r��1�ZO<�Ƹ>(h?1��>�>�:���_���>L�l?�2?�(�>�{�_�����P�U>7�:?ͮ	?� A?��Z>ѽ���L��ک�L����D��0>ڨ<?��b�8U ��u�>���>�$=�R�>��>i9i��숿�E;��W��v ���u�>gL�>�����6�iA/��L������=)?�?�钾��*��R>�\"?���>w�>v*�?qF�>��¾ͱȸ!�?3�^?<QJ?�7A? <�>�=�?��C�ǽ�&�Z�,=�s�>��Z>�ul=.��=�}��I\�y���+E=���=��ϼ6׹�9=<\x��:�P<�h�<�4>�ͿY�Y�p���,�?ƾ?� ������_=����6�I�A��5��;
���w���=�����U� uH���9.�?��@��*�)���7��S��O�>q��AP;���˾\>��=���$����b�x��j���V�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >]C�<-����뾭����οA�����^?���>��/��p��>ޥ�>�X>�Hq>����螾v1�<��?7�-?��>Ŏr�1�ɿc���z¤<���?0�@�|A?�(�����V=���>�	?��?>3V1��I�-���nT�>7<�?���?9�M=��W���	�e?vH<��F���ݻ�=;�=<?=���"�J>mU�>���uSA�>ܽ��4>uم>q�"�?����^�m~�<��]>��ս�<���Ԅ?�y\��f�h�/��T��J>��T?�*�>�.�=��,?�9H��}Ͽ<�\��&a?�.�?���?��(?�տ�6ٚ>Q�ܾ̈M?uE6?���>c&���t��y�=(�%{�����0'V�V��=6��>{�>�,�G��O�c��a��=������̿�7I�P��d�=ʟ��k��h��]���u�~����ׁƽ���=l4>�:>x�>>|u(>4K]>	�V?]�i?Pˠ>�n>��L�]ھl
��﫻r����C��L�Ľb�����Ⱦ����tt�FY�)i�UK;�.>�-i=iaS�S�������yb���E��@/?�@>o�ʾuL�<�W<�Zʾ�����+}�᪽½˾�/�sk�
��?�1??���lS������?���2�Z?ݻ�~0�H��%��=ڧ��2	=A�>L��=xU޾�00�1�Q�4v0?�]?х���[���*>� ��x=!�+?r�?�[<�.�>�M%?L�*�sK佨`[>ܞ3>�ѣ>k��>r@	>���cZ۽ɋ?`�T?:�������ߐ>}f����z��Ha=�.>95����B�[>F�<!���>\V��i���<�zV?X�>k�'��S��k��EJ`��ɹ<�|?1�?��>�yo?ڝB?���<����uR���
�4�K=�X?�@h?�#>�<��:Ǿ�6�� 5/?p\e?�0Z>��s�徏�(��2���?�m?(<?^�����v��#�
�YO1?��Z?��?��퐿�m⳾l�{=S/�>G?ݺx���>���>���ỿ��ſ��ᮣ?��@���?)�>&��=���=���>ɵ>
�6��1_���>i���@>w�?D�Ѿ��c������.ͽ��?,��?|i�>�6|�E촾���=�ٕ��Z�?��?�����Cg<U���l��n��K~�<�Ϋ=���F"�����7���ƾ��
�檜�ῼͥ�>AZ@V�b*�>�C8�X6�TϿ ���[о�Sq���?U��>��Ƚ����9�j��Pu�^�G��H�ʥ���1�>v�>���>���-�{��p;��^����>se����>K�S�o��ɝ��ߤ5<��>��>��>a��kܽ�Rę?�l��b<οT���'����X?�d�?bs�?�k?L�7<{w�<�{�	�z)G?�s?> Z?!$%�V(]��7�%�j?�_��vU`���4�uHE��U>�"3?�B�>T�-�T�|=�>���>g>�#/�z�Ŀ�ٶ�A���Y��?��?�o���>q��?ts+?�i�8���[����*�$�+��<A?�2>���G�!�B0=�SҒ�¼
?U~0?{�e.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?۝�>^J�?��=���>�f>o���Jf=���,�]<p�uz�>�D?���>��x>�����)�w�R�P|�qy���<�=:>��x?�M?��D>�j���9��(1�M����FA�{VU=�I�������@��E�=h�=#�8>�� �Q폾��?Gp�1�ؿj��cp'�h54?�>*�?2����t�����;_?�y�>7��+���%��(B�c��?�G�?M�?��׾�Q̼�>�> J�>��Խ~���|�����7>=�B?J��D����o�9�>���?�@�ծ?Zi�޳�>�3�Z��3����������[.��S?/�$��eF>��>���j���7Z�W�>:w�?B��?Y�>�q?C`]��$�l�v=�>�ˁ?/$?Jς�>L �QV>q?�S��������L�0?��?��@YCF?6����~ܿ~��i�����>��0>`Fe>���E�=r��`���<�	>�o�>Z�U>5L>�N&>���=Q�,>I݆���-�'W������Y;����]�1Q���_	�I��}����i�f�?ȽQ��P�ɽ^q!�z>a����t2Z>��b?�&�?�?��>��f=Zmu>��}�)<�D�ྺ�<�4]�>C�6?cD?�x�>`�y�7�O$�������ƌ�>s��<)�>��>.��>d?�q�>'x�5�>00M>D�9>^p�;K����Z"�����X�=`�>�*�>E�?�><>2�>Yϴ�r1��:�h��w�8̽#�?����"�J�L1��8��P���k�=�a.?gz>���j>п�����2H?����*�ʳ+�b�>��0?scW?�>����T�p3>+��x�j�eb>^' ��xl���)��%Q>+l?��f>R;u>�3��^8� �P��{��0r|>5&6?궾�Y9�}�u��H��Qݾ�ZM>���> �D�An� ���V"���i��O{=#}:?��?h)��1۰�"�u��V���DR>(\>�/=��=�MM>�*c�!�ƽ�)H���.=���=R�^>S?��+>��=L��>sp��ՈP��z�>ˋB>,>� @?f�$?���$N��������-��w>���>�'�>��>JhJ��˯=���>��a> i�C_�������?���W>�}�"�_�b�u�R.z=������=���=� �%1=���%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ)h�>�x��Z�������u��#=A��>�8H?�V����O�9>��v
?�?�^�۩����ȿ3|v����>P�?���?i�m��A���@����>-��?�gY?�oi>�g۾_`Z����>ǻ@?�R?�>�9�2�'�{�?�޶?ί�?J�]>"t�?_�u?��>S�ֽw."� _��(Nz�l�<�;���>,K�=T��@�?�������� u�&@��?�>��?=�m�>�!�'&��D�=�	�dy���7}���>�lg>,�>��>¥?3��>D�>s�T=wl�ý���oj�P�U?�?���oL@�e3=ƺ� ؽ���>B�?B��A����?�dT?�3t?Jth?@�d>�s7�LN����ǿ�P��F�o:�>
?C�>������>��*���e�c�>}��< 9���3оi��6^�
�>J7?�TL>���Q'?l�6?��>�3�>�Q��]����>��?���>u=�>�k?��?WK�]��j��ǭ��&�}���=Y��?)�?o��>���\~��4\��|��|Z�=J�O?�?a?��>�L?u}�?D�D?k�P?(	�>��d�����gL�=�>s�!?����A��L&�y��?�Q?���>�1��&�ս ּ���@{��� ?�)\?�@&?Ӝ��+a�E�¾�3�<�"�jzU�J�;�nD�p�>L�>#���U��=�>�̰=2Sm��E6�$�f<8i�==��>��=�27�8���EJ?mڮ��Yټ��߼@m�?�_����>^U>�־]Y�?I�6�
<���c��_q����`���?���?Zу?G_>5K�6?is�?-��>4�>1��c�ľ�Ͼ6'Ǻc�:-o��>�?��A>���^������������?�<C�#��{�>�W�>C��>�h ?�\B>[�>����fx!���� <	�y�Z�^!���3�\�3�����K������G�cT���*�>�����r�>l�?��>���>5�>	�A��׆>^k2>7E~>M�>j e>$>'R�=�}�<(-�~QR?���>�'����F���|B?dd?a?�>%�h����_��,�?���?r�?��v>�vh�@+�P?J�>.��vs
?�f:=g�
��V�<�S��jq��뇽=���>|�׽�.:�oM��f�g
?�??X����̾Cbؽ����$"o=)N�?t�(?��)���Q���o��W�0S�����-h��i��(�$�:�p�3`���%��W�(���*=J�*?�?���������&k��?�cif>��>`"�>"۾>�zI>�	�7�1�� ^��J'�����qL�>�[{?ʃ�>�|I?�<?��P?�wL?��>Jx�>���\4�>�u�;@ߠ>/��>��9?��-?A0?%K?vF+?�}b>�u������;�ؾ��?<~?�c?�)?-�?ꕅ��'ýC���<`�$�y�]�����=�w�<T�׽�t�kEW=�"T>T?����8�'����Ck>,�7?���>���>����-�����<��>b�
?�\�>���epr�8Z�uE�>?���px=5�)> ��=�N��_���r�=� ��Q��=My��>z;��V!<���=�Ք=ep��?"�Y��:�y�;�ݯ<QM?�8?�kp>PP�>��޾j����^� ��>6R�>�^-=m��>�ݾB������t2��Ǎ>�k_?���?_q<�@�=c2K>?đ�m��Ӿ�{�.�L�3?vv?:m�?�V�?�Qr?+"l?�>kJ��z���葿��;i}?�!,?���>'��İʾ�憎�3��?X?�;a�b��K;)�i�¾��ԽI�>�Y/��-~�O��|D�����.��F���ě�?���?�A���6��y�9���4[���C?T�>�R�>|�>�)�B�g�w&�@6;>@��>	R?��>��O?��{?��\?�+U>�n7�k5��uE����\��z>]�>?_L�?��?��x?��>�p>�),���⾨�����!�����;���4Z=�h^>㫔>_��>��>=��=3Ž]����?��J�=�'a>
��>j��>�g�>E+z>��<�G?�i�>�r��c8����6z��ȧB��u?���?�*?��=l���F�a�����>�O�?��?�*?��R���=�@ɼ������r��,�>�\�>@I�>XU�=דB=�R>4f�>FJ�>������I8�U�L�4
?/F?�=��Ŀ�K��f�۾�<��SS�=���(�k��8v<��n��|X=��@�g6)�����E� ��i�����v������k��?�`u�+,̼H��>tq�=���x��=)�>6=���Խ�u���Oq�7��=��A=�0#>�V.��+�=��^<w�Ǿ��{?�8J?Z�.?�:E?��>K >XR���>W���`�?�T>-D1��]���-<������V��ibܾ͏վ$9c�K���G	�=��l�Y�>�<>,��=�Q�<p=�=2�k=���=�L�,J=��=�n�=�f�=��=��>N�>*�v?�E���D��"iQ��:�$9?$��> \�=3Ⱦ��@?�9>ct�������a�d%~?���?}��?�a?g����>g�����2�=1𜽟�.>,w�=�!2��ͺ>ZbN>������*�����?�
@ē??T����mϿ�n->��7>� >��R���1�f�\��b�l�Z���!?`U;��=̾��>!z�=Gd߾H�ƾ�.=4�6>i�c=��G\��0�=�{�p<=)=l=�ɉ>�QD>׺=/�����=�I=t��=��O>�5��Ӿ7���+��n4=�R�=I�b>�&>6��>��?v0?3e?��>S�m�S�Ͼ:9���k�>��=>i�>�Q|=ܾ>>��>��7?��D?��K?B��>_a�=�+�>���>�F-�v*m��2�����ô<m��?�a�?~�>�3�<<'A�ZZ���>�1�Ž��?�X1?P�?y��>_��T��H]V���j��ţ:L5�=tѠ�l$ž�#F��F���ʽU�<eAY>�E�>��^>T��=�">u�=W��>���>��>I=��=.�H=A�S���6���X=�𢽖�7>�
*>�a<>-��7v����<�;Ľ��Ž���==�m=o��=���>{��>��1>��<
�پ��>
&��L�/�i�>�I���@��J��p�Uv=���r��> x\>�JY�-�����>[T�=&J =��?t}?��tR���0n��L�A�U��;$8=9�]>1yZ�w�^���k�� �ô"����>�>	�>õl>?,�!?�L�w=�⾬[5�2�>�r��	���!��7q�B��}���}i��Ѻ��D?�D��B��=@"~?Y�I?=�?p��>>��͇ؾ	0>_Z��u�=9�$q�0C��2�?]'?k��>�쾃�D���ɾ����`>t▾w�N�hI����=�N>�5��Z�>�(۾/w��f�P���z�o�L� �Gf��#�>�,B?_[�?K�Z���O�V�[��'1�{h�����>�f?��>E�??1���0�D{�N���;�R?S�?I��?�h�=���=|֑��\�>u]�>\w�?��?��}?�S��Ӵ>�� �`Z�>m5<�B	>!2�>i��=Ck�T�>�s�>g��>%,��������A��y&�|>�M	>T�>"��>���>�q>�F�=��'=	*;>�[�>��>8�>���>i��>��������?���5t�>�?*��=+��=F����;D��Sd�o,�����q�0�v�f;�	<$,�= ���@�>˻��=3�?X�>����8?�O�)�7=��p><��=��o�c(u>%�L>Vӌ>���>re�>�)=2�>�>GӾ~>����d!�y,C��R���Ѿ�}z>��	&�{���u���AI�n���g��j�B.��'<=��н<H�? ����k���)�%����?E\�>k6?�ڌ����1�>+��>�Ǎ> J��&��� ȍ�#h�i�?���?N��>l��>ʭb?k�k?܏���)�@�g�<S�� �Mw��>U��ݚ�
����� ���=��m?*(a?W}\?��d�&��>KI�?)	Q��#��>?>u^3�b�߾{W>�D>�ȾюS>D��3��k�lf>I�??*ot?�=?�Y��=M�0;A��>:��>ؔ?�*�?v�n?5��Q�?�<�>-	?[�
?h�4?�xX?C�=?�,D>e�>��y�1>��<�L�Ȭ��k�"��l��5e�=cJU=r��=�n=�f�<Q�;�o�=��t�(�<�����c=���=
�>"2�=ܕ�>�]?e^�>1C�>Q�7?�~~8�ò�� /?�:=�킾�7��xӢ�k�&=>��j?�?�TZ?�#d>c�A��<C�D>�"�>�v&>]>{��>>�@E��Ȇ=�7>�	>��=4�K�����w�	�jđ��:�<��>���>�*|>�;��g'>����iz�(�d>��Q�����mS�\�G���1���v��$�>�K?,�?�)�=�F�]���jGf��0)?�H<?�(M?��?X�=l(ܾ��9�(�J�k���4�>3��<"������7��|�:�ܾJ:d�s>t��"ܠ��Wb>����n޾��n��	J����7M=��O.V=Q�B�վ�$�װ�=�
>����� �g��-Ӫ�x1J?<}j=B}���XU�^m��O�>j��>#ܮ>��:�Q�v��@������:�=���>�;>.d�����1}G��4��V�>/�F?�^?�H�?_w����n���=�0��������Op?+�>��?2B>�|~=A��h.�o�d���>�{a�>���>�.�a@E�����6h�/��ۆ>��?>9%>��
?@�U?~e?A�a?p�-?��?�*�>e�ǽۮ��rB&?���?�݄=U�Խ��T��9��F���>9�)?�B��җ>*�?��?��&?�Q?K�?��>�� �9<@�>��>yZ�>~�W��b��>�_>֡J?5��>	6Y?�у?>>�|5��٢�󙩽]o�=�>��2?�-#?5�?���>�(�>-m����=:@�>�Ad?GX�?�q?f��=��?Tp0>�C�><�z=H;�>���>-I?��L?r?�4F?���>M��<�ԭ��Ӹ�\��ţp��T�;� E<"G|=_��oo������M!=�<kc����9/�P��i��}+�T�;�G�>S�s>}����0>Z�ľB��D�@>jɣ�V��6֊��y:�kY�=���>�?���>�H#�Ң�=n��>�@�>\��D(?>�?`?�";M�b��ھGtK�H �>\
B?���=��l�'�����u��rg=��m?��^?LW�M���e?dyk?"����?��k����H۽��?b��>�_��'�>��x?��|?1C?���=E���J���k��<W��'=��t>�4�#vl�3g�>9�!?'��>�>���<�־uG&�r辽�F�>[��?a�?�_�?=�#w�A�࿠���_K���]?Iy�>�*��;�"?W�j�Ͼ|G���$����wӪ����J���H���{$�ֵ���ֽ璼=u
?�)s?�Gq?v�_?�� �rd��,^���+V�H������E�qCE��C��n�6T�{�������>�G=�_�(h5�Q�?W�(?ےp���>T����p辝ㆾ�~
>�/¾yt3��m=r��j��=�1�=�,��q�`ӾhF?\��>�m�>�FT?�Ë�WbS�L:U��U)�{K<���>���>J�=�T�>o�ػ�k?����U�ݾd�O�a1�k�w>�~c?�K?Go?�����0��5���!��A4�"Ĩ���B>E�
>Ԇ�>	�Y�$!���&�G�>�ݍr���������n	��}=�1?`��>��>R�?j�?n�
�����|�y���0�)��<�p�>�{g?�$�>��>�Dҽ" ���>�Jm?Ȟ?��>�����A��xf����i��>N �>��?c��=
ǽ��X��ꆿ�}r��H��Z=1pJ?�R���z0�T�>�,;?=-����>���>E�]�w���9�]���ξ�hx=���>֪�;I�����������7���>��	F)?�6?ů��ډ*�q�~>�Y"?ظ�>0ۣ>�#�?�"�>_3þ�#����?L_?�9J?q6A?dE�>�p=�ձ��5Ƚ��&�TQ,=@�>��Z>�$m=u�=��Fg\����bE=�j�=l"ʼ�a���<ԩ���wT< ��<�3>�ǿvJ��)ؾw������W㴾kB�=�9���#r��쑾#����ݾ����P���I�R�o���@���ӽ]J�?6�@_ �����`���씿V-Ͼ!?��h�>�=�����y�Lپ�:�(��)�P�֍��e+�%	�$�'?y�����ǿͰ��x;ܾ�  ?KA ?��y?��ٞ"�y�8�w� >�;�<�2��|��ٚ����ο馚�-�^?-��>���1�����><��>ҢX>�Fq>����螾�1�<��?Ɔ-?��>;�r�$�ɿ=���~��<���?�@}A?��(�f�쾫V=T��>��	?�?>SX1��I�����:P�>�9�?���?rM=1�W�T�	�,{e?e�<�F���޻���=�D�=)=���C�J>L\�>��LA��;ܽu�4>5؅>Ep"����}^��ھ<�]>��ս�G��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6��{���&V�|��=[��>c�>,������O��I��U��=�S��˿�H3�/��<>��G=�G�o���(|�������WE>��>�u�>�|r>"x�>�`>��=��>�_?:2>?��>s(B>�*�%���=��ټ=�k6�>r�0i��~5���������;L[ ��u�n���ś��!=��э=�4R�+����� ��b�9�F���.?If$>	�ʾ=�M���/<pʾٳ��X�����!̾�1��n�͟?�A?����V���X������Z�W?�A�����ᬾr��=�i����=��>�7�=��⾬3�{pS�=3?�!?ٱ�C}����>�M����/<�w;?Ae1?��=>p?&�?����B��C>d.>%*}>���>i��=tУ�p���̓ ?d�=?g��BX�� ,�>g��Ϟ�����=冕=��]�m�6=��J>K�P���]��qͽ�X<�@U?א�>��#��=�wL���M�Oﻶ�?�O'?4��>^�?��>?��7��i����C��'��#�3=��V?�__?2:>$~;���˾<žp�*?j<I?J��>����7lܾ��Do��r?��p?�?|6��4z�R���p�y�#?�l?��M��v���Z�*5Ⱦ�;�>�V�>���>�'�*�?-I+?W7�]S��p�ſ�#�r�?B\@U�?g�=�����ۨ=�%?Q�?�uY������U��s�F�9�0�/>���q}���T�ZQs�G#?~�?�#?����&����=hٕ�[�?��?܆���Ug<��xl�k��O��<Tɫ=���H"������7�C�ƾ��
�W������d��>�Y@o]�u,�>�J8�p6�TϿ����VоIq���?{}�>��ȽO�����j��Nu�c�G���H�m����X�>(�>蛔��ۑ�.�{�g;�"�����>��^�>p�S��,��و���$4<]Ē>��>���>L஽>Ľ�|��?6S��K=ο�������X?Fd�?�g�?�q?��<<�v�o?{��%��"G?u�s?Z?}q%�K�\�w�7���j?/`���U`�9�4��IE��U>"3?iE�>��-���|=�!> ��>�a>�%/�1�Ŀ�׶�h������?��?Qo�h��>���?:r+?�h��6���Y��8�*��,�):A?z2>����Y�!��0=�OΒ�0�
?L�0?Wv�Q.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�b�>�?�G�=�7�>&,�=����G�#���">9`�=��@�b�?ikM?�N�>��=E�8��/�ieF�dUR�0�@�C��χ>�a?�ML?(�a>�㷽W,0��� �D�νC�1�7=�A��+�M�޽��3>:�=>��>s�D�&�Ҿȣ?���iѿ�'�������l*?�2�>`�?���	��=��N?��>�K!���������$Ͻ�B�?.�?/??�ܾj�N�*�;b$�>,��>�g��)���d0�{�o>Ys<?>�y�Q[��bia�Z��>��?�@zo�?�b�\�?�G�R ���y���6�E��?x>Ơ??�ؾ7��>?�?�x�=�c��&��I�k��6�>��?ߓ�?
��>n�U?~c��G4�j|��{�>Mh?���>y��ǾG[>�g�>�3���i�����1n?�@t�@a,b?�%��|�ؿl�����ľEž$n�=���=�>���� h=��Y<�ͼ-���P!>M2�>�Iw>��q>�UI>e�->u�
>9̀��G�� ������*;���f��iMm�֎��v�u���e��������ӽ��˽2׊���C����?6`�a��>kc_?:�7?�u?��,?���>�?������A���'?����/?��u?�"?��=����B؍�����$������J�?>+�>�ձ>i��>�O�>�U7=^�x>�>�=K �x�=fÉ>��=���=��i>�9�>M�>�C<>��>Fϴ��1��i�h��
w�|̽0�?����S�J��1���9��Φ���h�=Hb.?|>���?пe����2H?&���y)��+���>|�0?�cW?�>��d�T�5:>:����j�5`>�+ �l���)��%Q>vl?�g>ړu>�t3��18���P����V<}>X6?������9�l�u���H�^ݾ)N>}޾> @��d���YI��j��z=f�:?��?���㽰�H`u�����B�R>?,\>r=%�=DM>��_���Ž�/H��-=7
�=m^>d�?�[G>ǣ�=��>OȖ��j��O��>�o>s��>��L?O7?�p������V��K�*�UHq>Nn�>���>^[�=#9H��K�=��>�"_>��W��������=�y�?:>XS�Jw��׶��8�=?����$�=p�a=f��ڞO�s�<=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�:�>3Z������Fs��ρ��J��Ti>]v^?Z���T=�-����>sK�> �H欿�Q˿/:d����>`��?,|�?
�h��'����'���>���?�\E?��*>�1Ѿ�G�UB�>cC$?�J?sW�>$��t˽f��>e��?�Bh?9�s>� �?7�u?|
�>:\��h���ꚿ�Z|���׼ra��gԊ>���oT��H�4��k��^��c�u����>l_=-d�>��X�V�¾̺=����Ђ�O�9�"�>�X>�>2Hu>/��>1��><x�>1G<дɽY���.�1���P?���?X����G���>�#>����8v>���>�ER��븾x��>cHJ?�p?t?�;d>�Q9��ޫ������,վ�n���HE>�H?��>g�K=��=ba��:T��A&>ɵ<(
�Gh��VV���l���9�>��^?��{>5����A!?nk)?�g>W��>�);��-��ʦ-�F��>�}�>��>zj^?���>3u�����&��b����a��*�=�<�?�W!?"�T>�/��w}��B�F<c��D����c?��N?60@���	?��?R�>?&�A?7�>GO�@2�������>��!?K��m�A��y&��b��l?��?�)�>R��8`ؽn�ʼ<F�R|���H?˿\?��%?Q7��wa��þ,.�<-�!��#}�x�<�!.�J�>Җ>�c��SQ�=�4>�f�=�<n�^@7��eU<���=���>���=}O9�
U����?1)Q�U��-.�>�r~�PP?� �>�"��<���;6;?�M�����e+Ŀ`M��#�!����?���?���?������;7?�Ғ?�?GH?C��� Ǿc1��86�ݩ�t0���>�ƾ>�>�������-ݝ���t�A[��N��Fh?���>�?A}?�PT>�b�>����?�Yt�����Ga��z�G6.�6�,���Q��(/�m%=F�)���� ^>&p��(p�>ְ?�A�>�)�>DL�>Vuӽ���>�#>��>���>��W>��>w[�=�����C��aR?������'���龞��^�A?��d?��>i�o�;v����-�?�e�?��?
�|>
>h�8,���?5E�>{H��Q'
?W�3=p� ��̞<J|���i�w'���,�E��>��ܽw:��'M��3g��I
?�?}���sξ�T�ok��l�o=�=�?�(?�)���Q�ŵo�sW���R����h��R����$���p����l�����8�(�f@-=̚*?2�?U��.^�QC��Sk�/?��\f>���>��>�ƾ>�=I>�	�<�1�� ^�|X'�6���\;�>�T{?�>T�I?~�;?ѣP?��L?;�>�ث>װ�m��>���:Ǐ�>�3�>@�9?,�.?�0?Y=?�x*?��\>ږ�������ؾ�?^�?�?;�?$J?�焾]���S+��j}��^�|�4߀����=$��<�ڽg�{�f�^=�T>RX?
]��8�������j>�x7?S}�>4��>���d2���~�<���>��
?�7�>� �%�r�@i��A�>���?���t=��)>5��=]����Ѻp�=3���z�=h[�;��<��=�8�=�el��0n���:4-�;�[�<�>?��?ﱋ>{w�>����p�%��c4�S��>��?���>���>�lܾ`f���t��-�0���>��o?5Ѳ?���=���=m>E��#	�I�:��_����>[X1?�W ?��D?e{�?p�g?��?��F=x쾖����r�&۾& ?t!,?S��>a��5�ʾ�񨿌�3���?G[?c<a�����;)�N�¾�Խٲ>�[/�%/~����QD�� �����R��5��?保?~A�*�6��x边����[��S�C?M!�>SX�>K�>
�)�4�g�i%�31;>���>ER?y$�>��O?�<{?e�[?_eT>ܛ8�0�� ә��3���!>@?���?��?�y?sn�>0�>-�)��ྶP��g��6�r₾��V='	Z>֑�>�)�>��> ��=�Ƚ�Z��\�>�cg�=̏b>��>���>W �>N�w>�k�<6�G?I��>5 ���u�˦�����#1i��5v?^�?�,?��H=b���RF�ځ��if�>'�?ԧ�?��+?֒Q�Z6�=����.����y�~:�>2j�>�>��=�k\=�>���>T�>�;�����6���Y��?�]C?��=;=ƿZ�}�)����y���o6=�鉾h��Ty��G���/"=쨙��k�+u�����I?��h0������[E�����n	?�&=���=���=�˭<�>z��Ɣ�ts={Fy<�Y�=��Ǽ1"�<���|�������%��=��<z1�=�W�;ǂ˾��}?9@I?��+?��C?��y>�D>��3�㊖>͂��0?u�U>��P�܇����;�������x�ؾK^׾^d��៾�+>�I�/�>�N3>�l�=n�<��=��r=���=I�O�J�=�^�=oi�=�P�=���=��>�W>�6w?U�������4Q� [罛�:?�8�>={�=��ƾo@?R�>>�2�������b��-?���?�T�?E�?Fti��d�>D���⎽Ur�=)����=2>���=��2�F��>^�J>���K�������4�?��@��??�ዿ̢Ͽa/>O�7>7>��R���1�X�\���b��~Z���!?�F;��:̾8�>�3�=�߾��ƾ�S.=
}6>�\b=�Y��M\�8��=��z�L�;=K�k=�Ӊ>q D>遺=-����=D	J=���=w�O> ���% 8���+���3=_>�=��b>%
&>���>�(?;lE?N$?�B�=`�w���������> �J>ꅦ>� ��O�=>8�'? sM?z@?��>�跼���>�\�>��K���L��о�H�o}}�b��?ܒ?�i?HΑ>[V�9�$�o�F�%.�;�?n<	?� ?���>
�0ۿ_g�M|�T\�>J:�>� =lվڍ���r��Kj���>�G�>x��>���><��>m��>:A<�=���>�&=�փ<��R=ǌr�2`���9=m�U>F�:��>��2;ɕ->��2�����13 ��)�=�L�=��;��b>��=�{�>���>���> ��=%���&>�\�c�-��հ=�����4�Kh��5z�!#�Ț"�
N�>��>�볼D椿��?��:>z�=�F�?c9p?&g�ڽӼ�Ϩ�ܔ���ֽ�hI���e><��>�'Q��47�y:V���a�ޞb����>��>��>u�l>�,�?��w=]��%\5����>�i�������5q��C������i�r�ٺءD?0@���q�=	
~?��I?�ُ?���>Xv����ؾ9�/>sT��[�=-��p�!����?u�&?�|�>��ʱD�G��)� ���>�X���)m�������I�>�{>p���XN�>!8X�Oo۾�V(��Q��S8��g]��Q����>�Jh?��?j?���zr���9�Uu���f�=B�/?��"?�(g>�?� ?��½�Mt�n����O�=�?xZ�?�ҹ?��<�Ȯ=��,��>��?/a�?;c�?��r?H�\�$�>/50�*s>�N��R>7K/>���=�K>G2?�) ?:�?�Ư������羸����V���m=�8�=o��>��}>�B>8X>��=��=��o>*ί>�ߚ>%=~>���>��w>^-���[ ��E?�=���>�:? �>��;wz���׽��*��S�O�F�S]νHZ���_�=c�>(�=8�Ļ�2 ?�bɿ?ۈ?w�=�10�s`?�J�F�<
��>'D>.V2���>��G>�>PR�>Mf>c�=!k�>fD��:'Ǿ�A>��	+%��K�G"f����>Tt�������𾺨X�4���{��Z��8���U�^�R�&�2p)>#�?�B��N`�T
��o����>~�N>,�/?2샾� ]��o >cY�>r�>����Ĝ��-����-�?�F�?��c>2��>RX?�|?�T6���2�D[��]u�N~?���c��D`����of��.1
��W���_?��x?6�A?Z�y<2�|>��? �&�pc��5��>$0�~j;��"F=*��>����)�Y��Ծ�Bľ���8:D>�io?5��?%?�S���R���$>e�9?M2/?c[u?�7?Ӂ=?��U'#?61>��?�F?�7?>�2?�R?��0>�N�=+Z�`�(=�J��������ҽ�x�R� ��9=`�w=�;�:eI�;%s�<�5�<�z���t�Q7<�50��&=�#v=Q�=Q�=h٦>r�]?!�>X{�>��7?z��u8�n.��Wm/?j?== ��n����Ϣ�@��>u�j?}�?�aZ?id>��A���B�Q�>��>�\&>�[>���>11𽋓E�ց�=�i>{>zݦ=��K�.ׁ�@�	�y���>��<��>1��>*Q|>
����'>�a���z���d>R�к�dT�*�G��1�[kv�Bb�>K�K?8�?O�=cu�f����If�%)?�]<?�NM?��?,�=��۾�9�Y�J�X<�O��>�w�<B��̻��Z"����:����:�s>�>���࠾�Tb>.��|q޾R�n�[J����A6M=N��>V=f��վ�8�C��=$
> ���Y� �m��Zժ�f0J?��j=yx���dU�|n����>���>�ݮ>�:�B�v�p�@������.�=ڲ�>��:>UU����|G��7����>��V?#=?��u?�b�@Ju�y�V��s
���f�.���B?��>��>rej>&O�= ��������e��50�H��>�H?� �AWR�GFؾ�� �x�`��
x>�?;��>.4-?~�_?cUF?�P?57\?��?;"�>�#��@�ľق)?i��?���=v��Y^���8���X����>F�(?�HC�	�>��?�*/?#�*?i<Y?y?��=�d��E�6�>5��>.�M����P�>��W?ᦣ>n�D?�y?o4>�@��۾���~�c_>�1">ZU'?30?H?Q5�>�/?�Ҿ��d�I>�oU?�M�?��?*D�>J�9?�Ւ���x>>��>U��=J8 ?2�K?�{Y?ީz?[??��>���=bM<=
U��6(�3~�	�~Z�;mԱ=#$a��Z
<�Z��$��S��=h�<��"=�G��Y�N"�]�μ_�>&�s>�	��r�0>1�ľ{O��o�@>�����O���ي��:�ݷ=���>q�?���>�X#�M��=���>�H�>���6(?��?�?o�!;��b���ھ�K�E�>G	B?���=��l�r���F�u��h=��m?��^?N�W��&���b?�ih?�޾�7��hȾEp���B�	�E?�)?�@�?��>bǂ?�,�?8�?}���`�������g�V���J��={ߦ>/}�3$l�<+�>!A?f��>��a>���=�v径�z��ծ�$p?�H�?q�?QM�?z�1>FVh�|�ۿ��������k?��>�4���?��e=!y�}xs�P�J�����ش����i���L��������|�]W���=�m?A�g?��L?7e?8�־H'a�?|N��w����]���#e��6�*���9�b�0�KWm�W�ڏ�����(�>삈�=N��[�?�?^T����>�R�ES�Wǫ��o>0ɾ� A�2.�=%�Z���4"�=�F�(R��Ի��N?ޣ�>|�>,eC?%�@�D;�`(��3I�y���=�Z�>�>���>���\�e�#x#�������of��5]>��f?�5?@o?�H��3�|�b��0��|��Ȱ���>@�	><Z�=3g���K�0��,G�c�z�p�������,�R��=�G?�>q7z>��?�9�>:#�5�����ly6�~Z�B	�>Z�_?�f�>�t>ra��7L����>�@�?!��>=B=>�Wa����'����n`���?��?��G?îk>1RX��Q@�o҄����9��%'<��~?��v�N;����E>�n?�>>�ڋ�� �>FD �U~\��c1��a���݃>�9�>3w�=�4�>�5������삿����"�5?�?/����e'�ณ>\+?��?ci�>K�?n>�l��=L�?�/`?�uP?�}I?w�>�@=7���3�����=V�>�3a>��/=(Fl=��2�?���齼�=v�+>>�
=�+:��c�<j�����^=�>&�ݿ�L��ؾ=���{��������R0���{��:��kp��X��=H��Bl���"���c��8l�?_����c�[��?��?�x���Ã�㴗��H��iU�L̵>�yx��>������.�vϛ�	�辉б��y!�OP��|h��b�U�'??���d�ǿ象�Z8ܾ� ?�? ?�y?��4�"�E�8��� >U�<�x��F�������ο������^?���>���a�����>��>[�X>Eq>��f잾u��<��?��-?��>F�r���ɿ�����ͤ<��?/�@}A?��(���!V=���>E�	?��?>S1�^I�>���iT�>t<�?���?̀M=��W���	��e?x<��F���ݻH�=�:�=�C=����J>�U�>��{SA��>ܽb�4>څ>�}"���&�^�Ņ�<��]>��ս;��5Մ?){\��f���/��T��+U>��T?+�>�:�=��,?U7H�X}Ͽ	�\��*a?�0�?��?+�(?+ۿ��ؚ>��ܾ��M?bD6?���>�d&��t�ƅ�=7�A���n���&V����=b��>v�>��,�؋���O��J��K��=e��J�ÿ���  ��G#����[+����S��?'�Xѐ�i0���<E�6�J=w��=�� >N>�A>�`>0�U?�[]?ڰ>��0>��ؽ/w��V:���l����3a��{>�:�<�)v��g�	�k�򾜖�����f�¾$=����=�5R�ߗ��I� ��b��F���.?"p$>��ʾ��M��-<sʾ�����߄������1̾Ė1��n�͟?��A?6���|�V�$����1~����W?�W����I笾\��=sֱ���=�"�>\��=���3��zS�,�0?�>?�z������&�*><m��)=�+?A�?~�P<�ު>�J%?��*�W��+\>��4>�$�>9��>�	>�ா��ڽ��??�T?׌����Bm�>�%��� z���a=�R>��4��c�g�[>�b�<(���c��\����<�(W?y��>��)�	�sa��F��Y==��x?��?).�>m{k?��B?Mդ<h��w�S����aw=��W?3*i?��>����	оO���F�5?ڣe?q�N>�bh���9�.�TU��$?�n?1_?|}�� w}�~��p���n6?�*\?�
_�R7��	 �{�Ut>]>	?��:?><W��d?c�,?	R����t��Nſ�;�\q�? @��?o[��ܑ�o�=�q?>�?�t¾���Xoj>�9�pH\>��?c��� �.��7U�-1q����>H��?(�-?�Ӯ������=w$�����?ro�?�ܥ�q�<���(F��������<J�"=�)��}?�~{���>���Ⱦ"~�&�eo��x>T�@\�<����>�w'���׿Yƿ�x�@���P���?!s�>�(�JU��?>o���{���K��'L�:�L��M�>��>����]���S�{��q;��#����>��	�>A�S��&��䚟���5<��>���>l��>�*���罾7ř?�c��@οS�����g�X?5h�?�n�?q?-�9<��v��{�j��;.G?��s?gZ?�o%��=]���7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�e�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�9�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?+�a�N�p���-���ƽ�ۡ>��0��e\�N�����Xe����@y����?N^�?i�?ѵ�� #�g6%?�>b����8Ǿ��<���>�(�>*N>iH_���u>����:�i	>���?�~�?Qj?���� ����U>	�}?�>��?���=�~�>k��=������.��#>��=�=@�R�?�M?�	�>��=��8�P/�[F��PR�!�e�C���>�a? sL?�!b>�`m2�B� ��1ͽd1�l�꼭8@�qx,��y߽�5>��=>�,>n�D�N!Ӿ�?0��>߿vԣ�cl���6?X�S>қ$?�s,�"�w�E�j�?�}�>Dr$��������"��?�}�?
�?ˌξ:�K��\=>��W>��>�1�%�>����BV>��/?JΣ��ou�W~}�s�>k��?7�	@�0�?����>G
�ǿ��5����-� ý�=�uh?�y"����>��>��C�8I=�M���ji�YӤ>���?�8�?�O�>cb?h��G:�%�P>*>#�=?9�?E5�=�Ⱦ�9>�-?}����D��W#���_?sl@7�@��C?`��0���s���+����ܾ��^=g����|>�ҷ<��=lxi=�e�]7���ٹ=-��>^�|>�M>g`>/>�8>Dz���8�¤���?��zMX�`�f�Ѧ�!�^��(��[�m쾹N�'���/L���%�ຂ�����eF�t����>ߑE?]b?���?�GP?׊�=9&���~�=�z �=/.=&�$?s�9?Qwt?�yU?1N>�K����i��뇿��|���˾�Y�>�|>&��>d= ?�d�>�q�<S��<�I>dh>7o>x�=�>"��-��t>.�>���>��>�C<>��>Eϴ��1��i�h��
w�s̽0�?����S�J��1���9��֦���h�=Gb.?|>���?пe����2H?"���|)���+���>�0?�cW?�>$��J�T�4:>B����j�/`>�+ ��l���)��%Q>xl?=�f>�"u>3��[8��P��}��=\|>r.6?�涾�Q9���u���H��iݾ�LM>��>��D��l�r���y��hi�@�{=�r:?�?�L���᰾p�u�_C���UR>1F\>_�=%��=�[M>1�c�F�ƽ�H�.=t��=/�^>`�?)>��=���>������N��u�>\|A>Q{,>@?`�$?���RL���ރ�7m.��w>�t�>A�>�>l�I�?H�=&w�>R�a>1��%��&� S@���W>�z���`��Gw���t=�X�����=풕=���L�<�@�#=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ��}>��D��D��w���&�b�%Ic=�i�>WK?4
&���k=����v�>��
?sX�r���cdп~�k�><��?�o�?#KQ�	ը�|:�9�u>���?�;?���>}���l�;N�">�)0?I��?�*5>7�8�ٽ��?���?A��?�<>h�?y�K?�!>񑯾���ʫ��*��{��>��|>B|�>�Ƚ���W��N��������n_�!i�h;1?@w�=Y/�>�]�o%�Ã�>�OV���̾;7���?�k�>r��>���>
M�>h�>D��>&�=yJ�һj�pv���kO?�+�?-���G�֔�=W��=��	Z�>��9?������þw�>�	v?x�?	{?�(�>������Ŀ��O�D�'>+.?�?n�k�>����ؽ�';AP=��@�+i�Rz�;�X�=s��>�G�><��>�^�=��?h$?]�j>�O�>W�E�m푿�F�T@�>���>�j?E�}?Jy?�칾�2��8����a[�lM>��y?�?SJ�>�L������E�[�$PM�9욽f\�?�h?L\��?F�?q�>?}B?LRg>��ɵ׾�ᦽ5��>��!?�8���A�VF&����ڍ?pm?���>�G����ֽ�Q׼{���m���?�1\?J&?~i��a���¾��<���?����;TG�y�>�x>������=p>�=@�l��5��mj<�v�=Lx�>7��=sH7��d����?��ٽW��pÿ�M���a8U�f��>z/r=qڽ����?��<�IU�(خ�XP��l&徠��?b}�?}��?ei��V���?��?!��>%k?�%�2SӾ�}����bM����
����=���>� (��Ņ��0������Ƀ�Z[�=�=$����>IE�>��?�8�>��S>�6�>�B���W'�OU�����Z�8@�"/;���1��1�E�����l�0�e}¾�0��2Y�>`�.���>�P?�y>>U�t>�>y����>R�W>u��>���>�V>kk>� >�{�:�����KR?����(�'�~�辅���s3B?�qd?\1�>�i�?��������?���?Ks�?�=v>�~h��,+�~n?�>�>+��\q
?|U:=�>��7�<V��R��)3����1��>�D׽� :�wM��mf�uj
?�/?&����̾�;׽�����=}v?;�0?��5��E-��OB��|��c���;��������'�D�_��ќ����z�y���S1>��?0��?�y�X��F�U�M��\���>��?�֫>Y>�Eo���ܱj��$W��*��$��1�>o��?B�>�PI?�<?�)R?�!N?O �>R��>�ޭ�(*�>S{ �e[�>K�>9�9?��.?��0?�1?Ǻ)?�e[>O��E�����׾KZ?��?ĝ?��? ?N"���;½�.��	�h��aw�Hp��g�l=���<��ֽ_#j��x]=��U>�Z?���ԫ8�4���'k>��7?���>���>	��q3�����<�>��
?�K�>�����ur��[�2T�>�?���z�=��)>e��=:����PպjK�=� ¼��=�$��^w;��H <o��=3��=&�t�b������:�A�;,U�<�t�>3�?���>�C�>�@��.� �`���e�=�Y>FS>j>�Eپ�}���$��v�g��]y>�w�?�z�?ۻf=��=��=�|���U�����B������<�?=J#?$XT?`��?y�=?_j#?۵>+�jM���^�������?v!,?��>�����ʾ��Չ3�ڝ?h[?�<a����;)�ߐ¾��Խ̱>�[/�g/~����=D�/���_��6��?�?(A�U�6��x�ڿ���[��x�C?"�>Y�>��>R�)�~�g�t%��1;>���>kR?���>�GT?�~w?�UT?�Q>-*5�˯�qԗ�P��:��>T??:5�?yӐ?o'y?���>�>
�.�@���"����D�0c���1=�k>��>|_�>��>��=���M��<dR���=nh>S��>K��>���>��o>�ՠ;��G?���>^��E��
뤾
Ã���<��u?ɛ�?P�+?JV=���W�E��D��L�>So�?���?�3*? �S�c��=3�ּ}ᶾ��q��%�>�ڹ>�1�>�̓=�zF=�d>+�>(��>�(��`��q8��KM���?OF?窻=�Cп��}�rdｐR��B^4�3�(�2%���h<����9���i���þy�������r&��ԥ��+����6V�$�?���=��A=L ���=��=�C=��>:�7=��������K=�Ty��0A�����rv�Qu^�f�=y7��gŮ��p?W�:?h�9?��5?}I>���=�ӽ*
L>4��9X�>u�;>��-������� ��c���մ����ѷѾq�H�����78�=����u�<g1>y���o�=��B>�=��#=.Ǭ=Ѹ.=`�d=��e=Ť�=c�>��>]2�=�6w?X�������4Q��Z罤�:?�8�>b{�=��ƾr@?v�>>�2������zb��-?���?�T�??�?@ti��d�>N��w㎽�q�=C����=2>p��=v�2�S��>��J>���K��=����4�?��@��??�ዿТϿ:a/>"�7>�H>�R��d1�ւ\���b���Z�l�!?�;;�SY̾N �>�;�=3D߾Rqƾ�|.=�Q6>|Ma=f���G\��=��y��~;=�pk=>��C>V��=�Y���,�=��J=&_�=GP>; ��Ǥ8�
,�}�3=��=��b>�&>|��>q�?vc0?�[d?rD�>�m��Ͼ16���C�>���=�A�>M�=�zB>t��>��7?�D?��K?�u�>腉=c�>��>��,�ñm�Bi徱Ƨ���<��?BΆ?Lи>�Q<�A�����e>��KŽp?�Q1?/l?��>�U�3��kW&���.������8���+=ukr��WU������l��㽓�=4n�>���>��>�Py>q�9>��N>��>ީ>�=�<�o�=�X��<�����=������<��ż�a��='���+�䐦�>�;���;��]<&j�;�ɗ=��>>�9>���>b����}�o>K�����H���4>vȾ�C�W��;��k7�țý:C9>�>}�P��j]�>��>�q>���?�~?���<H�������;�]=\��En>B�>��f�dJ���f���f�,ʾh��>�؎>��>ŭl>,��?���w=��;`5�>�>bx������$��:q��?��N��i��aк0�D?�D����=V"~?@�I?F�?��>�@����ؾ�<0>L���S=^��q�J/��a�?�	'?���>:�P�D��P̾����ط>�HI���O�����4�0��b��η����>�󪾟�о�#3�(e�����g�B�^r���>��O?�? b�*X��$ZO�������.i?�wg?Z"�>�N?�=?�J���p�d���i�=��n?=��?5<�?e3>��=���r��>�?�Z�?�)�?x?ݝ�e��>�ꎽ���=í�;gu�=��1>V��=jw >5b?:�>�|?h����+���
��-��)���~t<��$>Vѧ>��>fNs>(y�=��r=��=ZHy>��>k�{>��`>w��>�C�>%͵�V+���:?2�=KG0>��,?��a>�z2��/½O�=�c�<,h��l-;הi��j���S�<���< e�=j�䪡>�1��֥�?X��>�O�p�?<�۾k�u����>�>ԫ��,�>�2<>���>ު�>؍�>�%q>s��>��<=� MH=&A��:�p�'���W�W5���r>�Ҿ�w+���ƾ4��y[������,���&��₿�c*���=�`�?l/̼?���l�A��D+��9?��>�l-?e�;ʆ1>5j�=��>X�>[�&F���Ǌ��Ͼ��?;)�?�:c>5�>[�W?�?��1��3��uZ��u�2(A��e�F�`�|፿省���
�p	����_?��x?yA?:O�<:z>F��?��%�wӏ�)�>�/��&;��><=�+�>�)����`��Ӿ}�þ�7��HF>N�o?%�?YY?"SV�F#�=�X>[�D?>�K?C�?�[?��,?ە���?u�q�@��>3H,?�B8?�/7?�(?�{o>ي�=V��������Ž��w����$Ͻ��
��4a=�>�dϽv�E=���=��O�����	���������qI<s=�=���=|')>˾�>)�]?�M�>>��7?���|w8��Ů��+/?��9=�X���Ȣ�r��>@�j?���?�cZ?H^d>"�A�0
C��> Z�>Ps&>\>�d�>��o�E��=�J>y[>Sĥ=.lM��ρ���	�E�����<(>x��>d5|>I��T�'>x��`0z�5�d>:�Q��ɺ��S���G�h�1�k�v�]�>4�K?�?ꓙ=�`龨9��fHf�<.)?^<?�PM?��?	�=�۾��9���J��;�8�>���<���:���$��^�:�KŞ:��s>�-������<�T>���T!߾r�l�O�M�i��==����H=`�	��gپ)ր��W�=� >Z�¾P#��׮��
8I?�=O����.[�Jv���l>�Ó>�V�>��F��Z�#>��ܮ��j�=��>�B>�������H��6����>�a?��O?]?���c�8KU����S���z��T1?�م>5�?��><+�=p��iܾ��n�e�K����>1��>�J�F�C�;/�)����m�5y4>�?�>�\^>�f,?>�}?��)?ws?GH?���>�Z>s��ޕ��^x*?���?Ig{=�*ν�P`���5��,k�@�>0$?�^}�cu�>}�?�3&?�=?R�\?�?A��=����]�D��>��_>��T�!h��mQ�>w[?�n�>�T?e�?�`�=	�V�4j�����G�=m'r>j�K?=r ?��?�݅>W�?UH��<DM��ܲ=��?��?�?�n?�PR?K_R<x��>��>��>��?��4?Ec?Ѩ�?(?���>�v�<0硽�`�����ν��;�X=��=�	8���?<���9,��j[<�g�����=��?r�"�=�Ӕ��^�>A�s>����0>��ľ�O����@>ą��YP���܊�)�:�Dз=o��>��?;��>tY#���=���>F�>����5(?l�?�?,!;(�b���ھݵK���>�	B?��=�l�큔���u�;�g=��m?ً^?��W�\'��&Eb?Eb?���`�7�0�ɾV9|����E?zu?��S���>��{?��r?�E?��C��Sj�SE��� d��䈾�=�?�>]����e��2�>P:?��>�d>��>>����}�ި��?�)�?�ǯ?�&�?�z>4j�� ߿!ﾬu���	l?���>�C����#?���<JzǾ����b��������Ԫ��׹����������Kvk�tՐ���x=;o?~�m?yi?�]_?�C���\�� S����T�B��j� (	��j@�KB���5��[i�?��	���5V����.=��p�!'Z��^�??J��c�>:ba�F��@¾|%;>�\¾��%�?}��\�����r�=eC��ת��㺾�	?{��>�Z�><?�>s��_8��+��-?�� 龿9~>��>p"v>��>Ot�<)U���n���b;v(z�So��k>"�a?�.?���?��D�Q60�s~S�_��ؼ�Ͼ�1�>w��=�����&�J��6��i/��%b�"�Ǿh�`��O��+�(���%?<b�>ϱ>:T�?w�>��F�\�@��}��#7���<�V�>1+E?¬�>RO�>F��,=��@�>��p?ˁ�>��>�+���<0�!錿G�i<�#?/��>��I?��>ܷ�Y1B��|�ш��\;�f��=�>k?�EW�-���	>�>l?1�>R��Dw�>����x4�f��6f��f�=wߪ>���=�H�>��ѾK��dl�O�����3?���>:v��ļ2�@�>��5?hp?Y��>5��?k�>�C�����=���>�H[?��M?��B?-��>�{=~{���󽱊)��r�=#>�>��>]#�=ǹ�=�ٽSbV�ѽ���'<���<��X��׽U�-_�;��=�Y�<�6>f@㿅�Y���ݾ���e<�-�H�G��̽����p�i������˞��9��^ ��|�'���A)���tl����?~��?yl��57������B~�5��Þ>�)��;��<�~m���S�l�b��j��r�i�D��U��=b�x{_�c�!?~���E�ǿ���W	վ�I?;�?n�x?�����,�/��\�=���<\v�~�zU��rZп�D��b#b?�u�>��j��R�>1�v>[j�>�jr>�Γ�����M!=Џ�>��&?�?��s��ɿ�����h<��?��@�sA?��(�-�쾥�S=��>��	?�,@>�1��E�k谾y%�>�6�?��?��K=��W�S�	�"|e?�e<S�F�������= �=p�=�;�}�J>�,�>����eA��ݽ̹4>.Ņ>H!�����*^��_�<�P]>P/ֽZ��5Մ?,{\��f���/��T��U>��T?�*�>R:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=�6Ἲ���{���&V����=Z��>b�>,������O��I��T��=\��ƿ�����;�r������S½��N�wrL�V�۾�`�l�n�[�=�oM=YX�=�r >�*>��A>9h?q
V?��>�O>���<B�1˨�F�������-����wu�=L��>d��%D(�"9뾓N���!��$� B��t�=�u�=�'R�j���� �M;c��6F�œ.?�h#>6�ʾ�nM�m7<�{ʾ���rׁ�tj���̾t1�� n�.��?B?х���V�_�ܠ��ẽJW?$���n������a�=����dd=��>�N�=�j㾁K3�MxS��|0?�G?�{��O|���|*>D �?�=��+?�?NfY<�>�>TU%?+��Z㽅�[>N�3>}�>���>�t	>h����۽��?�zT?O�\Ꜿ?А>�/��g�z�c&`=e�>zv5�,-�SU[>�I�<�Ȍ�_R��f��R��<�%W?���>��)�|	��f��q����==�x?�?2�>sk?	�B?���<�p����S�C�V�w=n�W?�%i?��>g�����Ͼሧ�;�5?2�e?T�N>�Nh����Y�.�>Q� ?��n?\?�����s}�:����nk6?��m?��Z��꨿���'����>��?�?�M����>��?�lj�lw�/���<"���?��@� @Y6k<z��$��=��?���>$@����
�R�>�u�ff�>D��>&���� �!6Q��匾p� ?�`�?N0?�X��Tq!�ϭ�=�����?�M�?��,.=���y�QS��p�=����HĽ�6�����l�S��u��F����s�����+K>T�@K=����?���5�ҿE�ÿ8&���%߾��R��Q�>��>�嚽�����nz�l2x�4�D��jd�m��<�M�>.�>���� ���0�{��q;��%��Q�>	��	�>�S��&�������5<��>���>@��>�+���罾 ř?�c���?οE������j�X?0h�?�n�?�p?w9<y�v�/�{�i��=.G?��s?\Z?	q%�;>]�7�7�T�j?�l���h`���4�KE��JU>3?ed�>ƣ-��~=��>�Z�>��>\./�+�Ŀ�̶�����J�?r��?o����>~��?�z+?Us��8������*�לܹ7A?;2>U_���!�-7=�������
?��0?�Y� D�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?�"�>W�?!y�=�j�>h�=N򰾡�+��k#>��=�w?��?<�M?(:�>q�=��8�1/��XF��IR�$��C���>�a?e{L?�>b>���-2�j!�`ͽ�O1��m��s@�w:,��x߽T5>��=>�>0�D��Ӿ�?�@�D�Ԙ���h�($U?^=,>�.
?a0��E��� ��?'�?	�����z��Vν
��?o��?o-?ѕ�<c'��=�>gr>\*+>�D����=B�m�\�_>-?�"�Ť���/���w�>+ �?p?@9�?�x��>"?�+��͍���w�P5���9�=��@?q�~��>�>�>�S=)Eb������Cm���>`�?<��?���>��`?" m���/��u�=�>��V?r�?0���ܾ�9K>C?_��"���	��%f?�@�+@�\?�L����ҿ1Θ�eㆺ��V�=%V�=X?>���%�=��R=��?=�/�����=�֠>~^z>Z8w>ŻL>��Q>�>
0����'�Q���p��}�H�C� ����`�����6u��O��緾�[Ⱦ�Q���˽J�����u�Qg����w�>V?h?g H?�P�?(@.?��s<���<񬳾�/>��|�g=��?��.?��o?
eO?��>T-&�+7q�����pY�����<��>7�Q>9~�>Y��>�T_>�
�����=F+g>��y>8+j>ԇ>����Q<���rO>� �>���>�Ɣ>�B<>R�>8ϴ��1��a�h��w�p̽$�?����6�J��1���9�������h�=Eb.?�{>���?пS����2H?����)��+��>��0?�cW?��>@��R�T��:>d����j�5_>, ��l���)��%Q>�l?�f>^�u>r 3���7��kP��o����|>��5?$ɶ���:�k�u���H�-�ݾ��M>kY�>PH��?�|����~��i�-�{=�a:?>#?�A��n��Z�v��|��9IR>y]>�y=�G�=C�N>�c��ɽ2�F���0=L��=}�]>�M?j	,>.�=�ܣ>Q��.P����>\B>o,>��??��$?t�������n��(.���v>�8�>jˀ>�>�BJ���=���>�}a>A���/���.�,�?�8OW>�n}��_���u���z=;T��7<�={y�=�o ��=�J%=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ\�>�����4�Z��D>�i�>/?+9)��(�=w��l?>�&?T���6���ٿ2��Xu?���?j��?��L��[���0�*q�>us�?:�E?���=��I�]���c<��1?�҄?n�>`o(���v�I�3?x��?>S�?��	>H�?^Rb?B̥>�\��b�1�A���퀿��Y>�6�> ��>�=7�ξ:�/��ꕿ�ez�;6]����+�>Zc<C��>M_)�= ����#>g���ؾ�R>s;.?��>PI�>+�>⿑>�<�>b��>Jf�X������Wm�+�M?���?����>	K�'0�=��=ʩ����>	�6?.�3�Q
ྀk�>�Z?�ц?�Xo?S��>�[�#˙���ÿ+ߧ�X�1���W>�>?4,?��x;k�>��w�Nr-��F7>�a>���=�ϻ��d��]m0<T,�>��?>'�>�LE>�?G�'?Xz>���>��L��7�K����>�b�>��?�#|?��?ܕ��/�����˞��X��<=>G+?��?���>��������<��^���߽MƄ?+�t?����?���?�[.?��??�s�>��F�Ҿ�OG���l>��!?�_��~A���%�ۚ�[?mj?���>r����׽��ټ,������O
?\?�&?�w�t(a���¾")�<��"���4����;:&J�(�>K�>o���.,�=�>x��=<n��m5��k<`�=x��>��=\|7�/z����?J+����¾?��Ћ�W3����>i��'����[~?�ù�V&����w���A����5r?���?2g�?����S��S,?:��?hk>,��>r����﷾.�
��!٧����NɄ>1e>E����t3�ř���Q��K����
�/d�L�?�o�>q�?\��>%y>m�> z��!�i��3���Y��'�����B�&���*���t��������*Tw��>L��9[�>�T??AD>�[>���>'�=�\d>�m�=��>�Ƚ>&�>��|>�> 霽�r2� LR?�����'��辵����3B?&rd?2�>�
i���������?x��?8s�?>v>7~h�,+�`n?�>�>���Dq
?>N:=gZ��'�<
V��=���0�������>�A׽A :�kM��nf�j
?/?v��g�̾@=׽[2�����=uԂ?�:?��9�c�E��2j��Fp��Q�e��=WF����;�����i�����Ŋu���|���$���>V�?wO�?1�������Yܾ��p���=�0�i><�?k��>�>�	>�� �����GE��/�\ٖ��װ>i�?bQ�>��P?�@?��d?��Y?�ڎ>��>����>}���L�>g�?;i@?�)>?�@?,�/?�
%?��=��n�����`�˾��?+P?K�?C��>H3�>-���6��\L���^��D�����z�<z3�<�=�����Г;=j=>�`?��;�8�M���3	k>a�7?-��>}��>]ݏ��%��g=�<�%�> �
?3T�>����lfr�OQ�\Q�>���?���O�=B�)>3��=U΅�Q!Ǻ7��=p����=�����:��;<�-�=���=�t�������:�l�;�d�<�n�>��?΀�>,�>a��� �P��꾯=1Y>pTS>��>K(پ)���&��$�g��Qy>#y�?�z�?&�f=&��=�~�=AD���m��'��h罾6��<۝?}@#?=BT?Ð�?��=?�h#?k�>�8�M��ua���0��Ѭ?v!,?
��>�����ʾ��Չ3�۝?g[?�<a����;)��¾�Խֱ>�[/�g/~����?D�����T��5��?뿝?WA�U�6��x�ڿ���[��{�C?"�>Y�>��>T�)�~�g�p%��1;>���>iR?�>�>^;T?��v?��W?��:>;�C*�� ���-����|>��D? ��?�Ŏ?�|{?��>�>f`'���辉��S�O��
ۋ�z~�<�i>�Ö>U��>���>,��=���ò�e�E��.�=�~>ͼ�>i0�>���>��m>S4���G?h��>:b�����Ӥ�⩃��<��u?(��?�+?�U= r�>�E�j-���W�>|m�?���?n0*?d�S�B��=�+ּyﶾ�q� �>�ɹ>�.�>��=�F=.w>��>V��>�0��`�?o8��M���?GF?�s�=R�ϿQ�r�b/��u�-�׽!o����|-��j��҅�=L4u��W��xb��ā�d�&�ݲ�����Q-���n��w�?��>���=7�&=R��a��HżT��=�\���>��<(C��H�o=ύ�<j�5=yl����ս˽�+=�ʾ�i}?FI?��+?yLC?�Px>		>q�8�C�>;7��#c?nlQ>j�X���<��0��┾�ھuؾ�	c��랾z�>�L�;=>Md3>��=Zo<�p�=f�|=�q�=TW���$=�3�=נ�=~��=�=r>�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>�7>�4>��R��~1���\���b�qhZ���!?qE;�GT̾,�>rº=H1߾�ƾ�n.=U�6>Mb=���U\�K�=�z��<=��k=&Ή>��C>�3�=�E����=��I=���=�O>������7�Mo,��3=n��=�b>��%>���>��?<`0?�Vd?[7�>�n��Ͼ�<��oJ�>�=tB�>Gׅ=AoB>���>��7?��D?��K?���>���=�	�>��>��,���m�`p徚̧��P�<L��?M͆?SӸ>G�R<ۅA���� g>�s7Žat?�P1?�j?���>fU���࿅V&���.�������p+=�xr���U�5���?h�����=�e�>���>Cȟ>��x>/�9>o�N>?0�>�>Ǿ�<fC�=�i���ƴ<�!����=U�����<�^ļd^����C|+������;�5�;ҧZ<���;*� >��>��>SC�>�2c;�����m�>lXȾkpD��_>�����(��3\�ʵ��gzE�A�;�_�r>B�>�s~�P�����><0�>4�=x>�?8�?�\�=f��K��i֣���9��7c��O>���=�
K���2��+d�kT��4¾���>�Z�>�>�Bj>��+�w�>�#�~=��⾧K5���>�،�Cx����jq�cW��|̟�M�h���
��ZD?�&��@�=�W~?/I?��?�:�>N����H׾QJ/>W9��"@=���,�n��ޓ��?��&??��>mR�0�D�.F̾E���[�>�6I�AP�����Z�0�B���Ƿ�͜�>s���R�о�"3�Jf������ߌB��Tr���>��O?1�?�'b��V���ZO����G4��Ql?<~g?�-�>�I?�E?w󡽟w��i�����=�n? ��?=;�?�
>�=����S<�>�i?(��?w��?��s?�+<��r�>&�7;�}>M����=�7>�z�=-��=@�?�d
?O�
?�_��U-	����3�a���<yZ�=���>���>�ls>y�=<k=-l�=D#Z>3��>�]�>@�a>*��>��>"�p�)�9��7?�=�0�>c�;?B��>��,=_�G�q�s��p���e��h���Ͼ�n���Wr=m�>{�+>ɂ����P>v�Ϳ�.�?�*�>����?;l��OT>�?>��=�K���>�ڳ=��~>"d?ug�>��<n��=��=����P��4��U�.�׍(�8Y��cľ>��>|B���
Խ��m��ʱ��??�����WS����v��퐿`�0���=�l�?-���Y����R0���=CQ?�o.>�K@?�վ��D�][>��Y>.t>��A�M=��cȏ�����?_��?�<c>��>�W?n�?�1�j3��nZ�4�u��$A�@e�ι`�j⍿�����
�0!����_?K�x?�lA?g��<�:z>��?��%�GЏ�T�>`/�^-;��<=|#�>"����`���Ӿ�þ�?�59F>a�o?�"�?�X?,PV�_��J2>w�<?�q7?!�?}�5?��1?^��'?� >Z�?��?Z�6?�06?=X?�v>`�)>T�߼��;W䤽~���Tѽ��ӽ�p'��L<=��=�H�Y��:@��<�p�:��n�x<	��<e���1�<�`�=s��=Ci�=��>O�]?+N�>��>��7?i���v8��Ů�+/?�9=�����iȢ����>
�j?���?�_Z?Xd>�A�VC��>�W�>�s&>�\>+a�>���E���=�O>�Y>ɥ=enM�΁���	��������<#>m��>�H|>�Ս�@�'>ur���.z���d>��Q�Ⱥ�+T�O�G���1���v��]�>��K?��?���=zq�k��k>f�t,)?�Y<?CM?$�?@�=M�۾��9���J�;��$�>&v�<������� ����:�X٦:޾s>\1���⠾Eb>X���o޾�n��
J�7��#M=�~��+V=~���վ�?�S��=�
>a����� ����$ժ��.J?<�j=�q��h\U��n��	�>��>"�>'�:�m�v���@�����V�=���>�;>�0��}�{G��6��\9>cJ?Tb?�sj?�6�w� ��X��	ھ�M_�v+	��?��>d*?���>�`�>�߽���Md��>�Py�>k�?�D�.�=�X#� ���X��>�U�>�Л<a�0?O�s?��?Yϖ?�J�?��>n�X>M����t���41?���??FҼEI/=�X*<~��/�A��7�>�,?�灾���>�� ?�
?�&)?�Q^?�+?�2B>���'[��#�>3�>rsV�#�����R>u�I?}"�>8-?YHb?0o�>�K.��'ľ0F�Ie=��>�dI?��$?&v�>��S>�YA?�!'��=x>x/�7�A?Z0u?�O?���>�E6?�f�<U��>/0�>�ӈ>1�?@�9?ݓA?��g?I�5?~W�>�E>r���]V�TJս8ؽ�k�=�O=��<FIռ�>=0�9?}��_�Ž�E,�Fg��v���������=�v2=/f�>��s>�����0>i�ľ C����@>؜���F��h׊� �:�޷="��>��?D��>�K#����=>�L�>Q���7(?m�?|?a�!;V�b���ھ��K�B�>�B?���=��l�"���b�u��	h=R�m?�^?�W�� ��!�b?�]?hg�\=���þ��b��龩�O?��
?�G���>��~?��q?޸�>��e��7n����Cb���j�|ն=�r�>�X���d��>�>a�7?jP�>��b>�#�=r۾��w��r��=?k�?��?��?<.*>��n��3�����WK��d^?��>o���= ?l�2���;r勾�`���n꾇���	o��ZΘ�\d��A�(��q���wֽ��=�?V�p?��l?�!`?����b�n�[��>|�cDX�ν �G��jnH�#�A�XTE��l�������ޚ��;�=\���Gh����?|9?���(z�>~��]���vȾ@�	>�����{� ��;�IL���2�7�=@�Ҿ�O�:@����?�v?|�X>3]?�]r2�s�� ,�o���>���>���=a�>�{�|=����UW���yC���P>�>]zd?F�-?��r?�Zz�7--�2c�)-��
]�l���{�V>��=���;�M�Q�|�{�B��#D��~�]4��t��8����=ȭO?'��>}�>77�?�\�>���>��n�my�E7>�ޱ>q,v?GA?�j�>V���J[M�W'�>��q?�J�>�Y�>|����c%��y�ا ��#�>!1�>�q
?��;>�%���P�j��n㐿�A��,=��l?����]�i����>yQG?C=�=:!=�`�>�i=��e1��@��2�I#>���>��=�gk>�Ǿ9���]~��/���~A?��?Fթ�A���¹>:W>?�!�>/F�>��?�b�>V?n���=Ǝ�>�T?lyJ?0�V?E�>�e|���K��vƽ�i ����=c�8>�`1>���=���=���b�0���Ž���=Y��=��轴hѽ���h���m�v;uF�=�kS>�lۿiCK��پ�
����>
�`爾����=d�� ��d�����Xx�^���'�sV�;c�|���X�l�8��?�=�?���X,��\������R���1��>�q��w���E���'��>�ྐྵ����c!�$�O��%i�V�e�n�'?������ǿ䰡�f>ܾ� ?�? ?��y?����"�8�8�U� >�B�<����!�������οΥ����^?���>	� D����>A��>}�X>�Cq>5��m垾q��<M�?/�-?���>P�r�s�ɿF���?�<���?��@>A?��(�����U=���>�	?a�?>�N1��B�����"U�>d;�?!��?�M=��W���	��~e?GG<��F��wܻb�=�!�=<=����J>-T�>Ո�jNA�{4ܽ'�4>�օ>L�"����^����<��]>��ս�4��5Մ?,{\��f���/��T��U>��T?�*�>Y:�=��,?X7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=y6�􉤻z���&V���=[��>d�>��,�ߋ���O��I��S��=5����ƿ�6$�o��v6=�{�H"Z��<�}y���Z�GF���Bo����y6d=\��=�Q>��>�W> �X>fW?/Fk?�=�>�>�C⽰`���rξ�{��������쌾q������6�쾠g޾�l	���%����ɾ�(=��Ս=|6R�@���`� ��b�F�F�h�.?W$>��ʾ��M�F,<�vʾ=ɪ��U��)9��o;̾��1��n��Ɵ?0�A?�����V�� �e���~���W?:_�����묾�y�=bٱ�1�=��>�S�=L��E3��vS���4?_�$?㗼��;{�%s�>'�+<�y =��!?�6
?|���$�>�?Ф��&�jC�>"�t>�s�>�8�>�S�<;¾��/�W�?"OI?з��O<��_��>~4���n� �b� >{�i������F>n�]�I_�������;�=�W?qό>l)��V��f�������J=K�w?H|?ii�>j�j?~tB?84�<���N�R���	��+=��W?��h?��>$|�t�о覾�'5?	�f?�N>�k��I较�-�`��\�?�:m?��?�3���	|�E���fc���5?yGU?�Kg�j�����ª��m�z>ĝ�>d�?�EZ�K�?�<?.k������%R����;�D3�?O�@A��?�P~��L����&=�*?{�?�Ί��
���=����x>��?%ұ�=_�Hr��*潾�?�%~?���>�+������=�����?⸈?�籾/�?<����cn�w��zG�<�3R=�&��@\P�!��T�8��¾D��n���&e�;���>x�@��2�O�?�q�,&��ÿ0,����վ�#D��?q�>�Ӎ�����?q�JOl�]t8���C�V�5��ģ>/�>�����6����{�	�:��	�� ��>f����>�S��������g�9<��>���>�҆> ���������?Y��n-ο����P��|�X?�P�?H?�?:i?��<<�u��i{��� ��G?^zs?Z?�&�G�]���7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�h�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�c�_?'�a�J�p���-�v�ƽ�ۡ>��0��e\�M�����Xe�	���@y����?J^�?h�?ĵ�� #�g6%?#�>X����8Ǿ��<���>�(�> *N>�H_���u>����:�i	>���?�~�?Sj?���������U>�}?w%�>��?�g�=~e�>��=��$O.�Ef#>.�=�?���?�M?nG�>k�='�8��/��XF�iGR�E#���C�
�>.�a?�L?�Ib>�����1�p!��kͽ@e1�ڇ��T@��,���߽;(5>
�=>�>^�D�*ӾOЛ>�#��b�1������y?�%:N)?f�.���;c� �f|�>V��>�,.��&���\�����w%�?Y<�?�?���I�νڠS>���>2��>hꢾ�Z�=V
ξү�>�%?�����O����I����>���?!�
@#�?sc� [�>�0��l��<<���>%����30��Gd?'�=�')?r��>��@���G�_譿��n��]j>ZͿ?H^�?�d�>�\]?��h����$��=�>��/?�p,?��>5���F�>�v?9���m����U�G?6X@��
@bY?�t��F���W
���☾᪾�P&=p?�0>�e<.H�;w��{�[=ŮǼ1Z >o�Z>8>;K�=��Z=K��=�K>� ��5z#�h£�"���_�"�R��r����!?�R�����M �xP쾰0�����\V���!�Wyu���=��/>��R?g�;?&n?�?�^M��GA��޾��=R����L;>��>x�*?\�Q?��0?{��=�ޖ�Emi��	}���x�]���>N�2>"�>!�>;�>M�=׭�>߃,>�>��=�!�=�폽������X> ��>��?��>mC<>��>Eϴ��1��k�h�w�v̽0�?����T�J��1���9��ۦ���h�=Bb.?�{>���?пb����2H?$���|)���+���>z�0?�cW?�>��5�T�1:>6����j�`>�+ �~l���)��%Q>wl?.�f>�u>��3�1e8���P��{��j|>�36?�趾�D9�r�u�q�H��cݾIHM>�ľ>�D��k�h�����<vi��{=-x:?��?47���ⰾ��u�C���PR>E:\>�U=i�=,XM>bc�Z�ƽeH��f.=��=��^>��?��+>hF�=:K�>����!�L�=!�>�iB>�F.>��??M�$?Z�x��������,�k�w>MI�>�?�>v�>��H�4g�=f�>�a>V1�gY�2�7@���W>$�}�͚]��x��qq=����y�=�1�=�� ���=�dj)=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾP6W>�aJ�]���ˏ����{���]���>�D?�<�v���c�+���>�k?�1��ؤ��ͿZ-z�K��>�h�?�W�?��N�]���7�>��#�>���?�5?ZS\>�Ⱦ��Z���w>�*,?:�o?�]�>{t��	�	?f%�?ݐ�?��>�?�m:??�Q���H��=��!���*i�<|�=�N�>2��#��,.��ڗ�_���+�e�T:
���?�@</��>�5�����,q>X������IM�>��u>
Y�>���>)B>D��>^��>-p߽���-e־�꥾FYM?8p�?@���4\�P�=VH�=eW��#w�>�/?�C��e��&�>��W?1��?��]?%��>Ip�R:���f���_��˝�<�:>[K�><x�>�[f�j�?>� ɾ{)�뉖>���>��d9뾳ڍ��I3�~w�>%�?(��>}��=�r ?�#?D4j>ɼ�>�|E�l>��x�E��1�> B�>oB?v�~?��?䦹�8K3����eڡ�L�[�8N>y%y?�>?j2�>t���~��hD�J�G#�����?�mg?�
潮?;�?AC??|�A?@�e>�����׾[�����>��%?�5�|�@�%�$������?�?3i�>"�R���Ͻ4�:���������?�\?�M)?�5��m_���¾x3�<���:����8��;��(���>��>�a�����=�j%>u��=��g��14�PL�<���=?7�>�8�=D�>��������>��M�7vǾA}�=�k��r�p���>Y��=�K���X�?���[���$���ў�����|�y?�	�?=�?u�n�&�O���??O��?�-�>�-�>T{Ⱦ��~�|�z�M>o4����R�R��>R|�=��#�n��ߋ����3:��6��=ߍB����> �>3?���>�:>�x�>�bþs[&�.����0�()P��7���̸�U�����y@��
� ��+���×���>�ǽRWR>�V?7͒>\��>���>}�f��g>��|>��>f�>dϧ>��>�S�=�ߤ=���cR?����/�'�^��֏���TB?Ftd?�&�>�tf�}~�����u?*q�?�j�?6Vv>�Ph��	+��t?LF�><���n
?x�8=q��c�<Lⶾ �����xM�ī�>6Hֽ1:�-M��kf�ee
?*1?�A����̾�׽8,��U�=�!W?��i?��A��sW�K�$�H�k��Q��T�=u���Wl������
&_�0����fa���y��f�|E�>fO?�3�?�Z�ƥ����վr�|���I%_>���>�\{>�\�>5`n>��Ǿ+;�Z_�}�+�����>�%�?_�>�tK?�<0?юG?>�P?Pء>�>�y�����>����R��>R�>f�&?aP,?��0?��?�h*?OU?>��$��Q�f߾�?�?¡?�X�>d�?�"b��н��0�7>;߃�xD��a�z==\<�X�8���[��=�!p>E\?��,�8������	k>�~7?H��>���>� ��-�����<��>��
?'R�>����=tr��Y�+[�>]��?���t=k�)>���=�Ӆ��DҺ<�=L¼p�=C&��F�;�1�<�z�=��=0�{�[�^��d�:�)�;��<Vt�> �?D��>wE�>�A���� �յ�pa�=Y>?S>Y>"Fپ�}���$����g��\y>Ww�?�z�?��f=�=���=}���U������������<��?:J#?�WT?6��?;�=?j#?Ƕ>+�oM��w^�������?w!,?��>�����ʾ��։3�۝?i[?�<a����;)�ߐ¾��Խѱ>�[/�i/~����>D��텻���U��6��?�?LA�W�6��x�ۿ���[��{�C?"�>Y�>��>U�)�~�g�s%��1;>���>lR?B��>�ba?�+Q?a�C?A!�>Z���N�z�V4�=��\��U?��?��?A.�?��!?��:>(K=�A�0�'�����=C"��梾��>Dd�>�>�x>�5�>�s5<m�Y5�!07�s<���;��!>Б�>fZ�>>9�=8�<L�K?�>q���/�65��Ya�G}��dr?]��?X�(?��=���^E�
��a��>���?M��?�]*?1�F�r >�蚼XA����m�61�>��>՗>?^= �_=UB >���>7��>.��;����3�
"�n�?p)??�I�=3躿-I����e��]Ҿ݃�=���b.�3�8�a%����V�����X!�;J��Y����Z;�H����پ�-v�P7��;��>��J<�>��K>���=�f�=}Xս��>)Zݽ���<e����s��}�> �)=�a�=0B��˽���J��Y�ɾu?}??H?;L+?�^D?U}>�>nf,��\�>OL����?KV>��f�����88���L��WپؾWe�KT���c>��C��1>�\1>D@�=���<��='�j=$=�=UK���j=���=rε=̉�=��=h^>��>[�?=?x�9���tS�C���W?#ʦ>q�=��g�5?UnI>-wx�Z��^�����w?:��?�}�?�K?�|6�2��>����8�ѽ�f�=�w���>to�=h����>�oj>���I���̟񽅓�?q6 @S�B? 0��o�Ϳr#>{8>N�>��R� Q1��	[�V2a��lZ���!?��:�6A̾��>=Ż=cV߾hƾ��1=�d7>W�d=E�3`\��
�=�|�<z<=�Yk=�ʉ>1�C>��=�k��	�=B�H=$ �=�O>����'�8���.�X�1=�G�=8�b>��&>��>۷?+B0?��c?m��>�2l�X�ξ����D�>�n�=w�>���=,�C>M�>�O8?�pD?aL?O��>��=�Q�>'P�>�C-���l������:s�<@F�?�t�?�M�>D�Y<�HB��u�>�ŖŽ�?��0?P?hΞ>�U����)Y&���.�ш��.5��+=�mr�:QU�_����m�4�� �=�p�>|��>��>Ty>�9>��N>z�>��>7�<�p�=ތ�\µ<������=����I�<.yż����g&���+�ێ����;આ;)�]<W��;����>X�+>9px>�[ʽ8�پ���>�z�'@0�_��>p��`y3���o�󨅿�P8�����d(>}�>�>���ȃ���>sn�>����Q��?��?&X�>ƁB�?t޾�+��#߽�n��mN<��>�h��#�#g��z�������>7��>y��>�l>,	,�%(?��Jx=kR��X5�+�>�g�����5��:+q��9��.�
i�7�t�D?�6����=�~?:�I?Q�?���>M����uؾ�/> �����=���1q�
	���?��&?�e�>gI��D�ر��=��$R>"i����W�T���!�Cd=�����>��7��(�'��ʌ�O㏿��d�4ڮ��B�>�X?�\�?2�
��ā���I���q�~<��>"lK?�e�>�%?���>��N�p�*�I�c��͡�o�f?���?w��?�]i>"D�=&��F�>6�?�D�?�?փs?�b8���>A6�:e4>:v���V�=��>�6�=X[�=CR?�
?�	?���M����"����]���G=,��=��>���>�s>�c�=��W=i�=:�W>H��>?��>8@_>��>s��>̺۾��9��XC?�!/�ULh>\��><x�>VU����;�B��-@��G6�jOϾ�k��yݏ�_ȇ=֠����=.��<�>�Rÿ[�?�BQ>����s�>�c'�S!>�Z�>ݳ��e���Ǽ>N>���>���>.�]> 3=�>���=P�!�4D��2T�7-.�	J�?m�ېѾmq�>n
�>H��| ��x��=$���
����鋿3[��ص7���=Q�b?a�8�~q���)��V�`��>gڠ>h�?������G<ݻ=U��>݃>@�%��P��
[���sξ�́?�E�?�9c>��>r�W?��?��1�3��tZ��u�w(A��e��`�O፿{�����
�l��B�_?��x?xA?؁�<O:z>���?�%�.ҏ��'�>}/��&;��C<=x+�>})����`���Ӿ4�þ�4�EF>�o?�$�?�X?�OV�,�=�G_>��-?�N?�;y?��:?�?�8:��;2?8�%<Y��>Q� ?A�6?N;?$� ?}�>~�>��(�/����,��b���?л]��q
�z����=�G�=��6�M=��_���=��뼺�ܻ�#=fw>��>;�<ŧ>��]?_��> )�>p8?-P�eB8�YE��K]/?��7=�<���܉��"����
�>'*k?�ʫ?l8Y?�j`>��B���C�*�>�ډ>�*&>�l[>d��>Ma�S,E�ڽ�=LH>�R>N�=?N�@�� 
������r�<�� >���>k2|>�����'>;z���,z�U�d>��Q��ʺ���S�E�G���1��v�
Z�>�K?��?��=\_��1��!If�?/)?q]<?dNM?2�?k�=��۾��9�Y�J��?���>"I�<H��x���#���:�U^�:.�s>/0��y���{jc>e�
�n4޾��m�J��N辦^C=v��)L=j[�K־=M�˾�=�b>���!��������I?��o=�S��H=U�I���jR>)�>1��>F�:�
yz�O)@�b���=||�>%:>t�����G���<��>i�c?V?q?���?���� �$k��.�s��^�o����>�L�>~�>+�>3��=i��j_/��怿΢M���>�>�a���U�F`��-�K�+��b@>��>���>��$?[�I?t�"?��?�5?��>���=�r.�����&?�ل?&��=4���EW��(9�dG�(�>Q�%?��M���>y�?�& ?�,?�-U?q?��=�=���G��>�߅>o�X�"�����y>p�M?¹>�\?HU�?��">"9����k��$��=&�5>Ya2?�� ?RU?,�>�b(?f4���#ľ��7>h^Z?K=�?�?�?��6>hR?b�kPٽ*��>�}�=m7�>��;?�v?CBK?k?
�>�
���Ƽ&������s���LK��C�=3KI=�� =�����Ļ��G<�T;��=+A<䓚<C�N=	��=Fm�> �s>�����0>�ľ7��cA>�����2���ߊ�4^:�數=k��>�?�ȕ>z#�|!�=S��>)F�>���l+(?��?#?`:';��b�O�ھۗK�a/�>��A?��=f�l��x����u�o�f=��m?�v^?�W�~���3b?�a?����`7��Ǿ\Ss��@�Z/I?Hk?��I�?ְ>v�}?V�s?K+?iP�`�l�C˜���c�\�����=GΘ>\��Q�d�^D�>�;?��>mu>���=b���|�	r��G�?ˊ?�{�?d%�?t�)>�j�L�߿ <���D��_Kd?�A�>e�����?DK��O�u�'֜�2U���Ծ�a������V��c���7&T�N�u�U��=�?�k�?�W?@��?@�0�|;m�^�\�-,���YL���ľ�X!�:)}�a14��9��f��`1�&M-��Z�����=�$��.�O��b�?�?� ����> e��a����FǾ�"H> �������=[����L=�z=�4�W�>֜�9x?3�>�k�>�.M?n�a���5��&��93��9��\�>��w>��O>W��>��<=B������⾂���^���c>��o?O�^?[�k?5Ƚ�I*���n�YI9���G�`����z>��>�:ż��oy?�Y�(�&�i�2{�+|���XU
�5u>:�;?�?�\�>�?8H�>3Y��}"��O��4�$�:$=�M�>+�g?��>%�]>N�qWa���>q ~?���>�Р>�f���*��A��
t�V��>��>�?'��>�f^��uR�����o��M�d��;/�t?Kl����g��z�>�zF?�c=>]R�<���>b� ��}>��q%��-M��\>	)�>��!>[>֜��;���z�ę��?�+?�]�>�.����#���>�e'?b_ ?*��>y<{?�È>������=7?>�_?��O?JC?�
�> �=����ʽ��)G�=0��> \H>�	���ޒ=x%�I�>��"�6��=�d�=Qk�	��)�=l�CIS�n=��5>J�俺_E�j����8'����(� �����<�ɽ����$��_�����S��v���f��3gd�~gq����Q����?V��?O�Q�o�پW���o����I
���>g������ppվЗ%�ü��3u����g�"��J��L�O�M�'�'?���x�ǿ���D:ܾ�  ?Z@ ?�y?m�u�"���8�>� >"B�<sR�����&�����ο	�����^?���>�=�����>z��> �X>�Hq>b���鞾�p�<��?T�-?���>��r���ɿ�������<f��?8�@��@?�/'���Ϧ�=���>�?%WO>)\A��<��_��g?�>�(�?��?��}=��R��𐼍td?4�*;�H��߻mx�=	�=O�<*���T>�͘>����7��mｬ2>�f�>��J���/��id���y<v�P>�����g�&Մ?�z\�xf�~�/��T���W>��T?+�><�=\�,?=7H��|Ͽ��\�+a?�0�?��?y�(?�ڿ��ؚ>0�ܾt�M?JD6?���>�d&�d�t�=��=�;ἱ㤻���&V�e��=���>��>܀,���z�O��M�����=�	��?ȿ���� 2��=��]n形�Ͻ��U��f=�+ҽ��޾%Ԏ��iu�tTm<��'=�<>t<c>1�$>z�;>8AR?��y?�_�>�Y>��݈��u��1`R�|�νC۽��w�m��T̾E� ����e��pR+�'����Ǿ+�=�8'�=��Q�V����� �c���F�ze.?Ņ&>��ʾ��M���<_ʾ����b���ܧ���̾Y�1�T�m�\��?B�A?����@�V�:��u����mHW?4�����ʢ����=����=lv�>-v�=d'㾫3��<S�c
1?�2?����Ւ�ޑ(>f���-J=�'?� ?"��;�O�>\')?�'%�X@����r>��?>��>7-�>C�	>����;wϽ�?^UU?R���Gߨ��p�>$���e���6=�|
>Y~0���켘�6>�m;hۄ��sü�h���N=��V?�j�>��)������������>=}�x?�]?+�>��k?�B?`�<W����	T���@y=��W?.i?BI>���Jо{0��h�5?ߜe?d8N>��g��$��.��x�$?�n?=�?�X��D}�u
�����o6?�h?�_S�$����������{>���>��1?�Hb��x�>�U^?��������ȿ��2�f[�?4�@%2�?��d=W�9�+9�=�?+?�hQ��
�n��=F������=�{?'8���.7��Z�i���.(.?�W]?+�?�7���{Ѿ�e�=+��t�?�7�?vPƾ�_�����|g�����u=�}c=���Z#Z�����N0��zؾI��n��z�<�6�>��@멣����>l��.�޿�Ϳ�$��&���q��O?֖�>8z��ү�9bq�����NQ�4]F�{v���>��>�l��z����{��K;��'���6�>1�
�R�>ƌQ��A���F���j<�7�>Ar�>�.�>���O���i�?6����οC9��?-�@�X?���?Ci�?� ?��'<�/y�; {�_���G?�t?��Y?��%��\�n�2��j?�_���U`�ю4��HE�U>�"3?�C�>��-�g�|=�>-��>�f>�#/�i�Ŀmٶ�j���i��?ԉ�?�o���>{��?�s+?�i�8�� [����*�41+��<A??2>y���.�!�0=�ZҒ�s�
?Q~0?|�1.�^�_?+�a�N�p���-�<�ƽ�ۡ>��0��e\��M�����Xe� ���@y����?K^�?f�?���� #�c6%?�>W����8Ǿy�<���>�(�>*N>�H_���u>����:�i	>���?�~�?Dj?���������U>	�}?�	�>��?#�=J��>��=}簾�R3�%�">q�=�A�ͣ?S�M?���>�[�=�8�/�KyF��FR���4�C���>��a?�rL?��b>P����2�� �8�̽Ȁ1�����@��I)���޽�n5>��=>��>i�D��^Ӿ��?#v����ݿ��� @q��/?���=Y&�>��ؾ�g<�'��&?�	�>�{$�����w�����)��m�?��?�?��ξ�4N��>a�>��z>��:�(=^����x�=�D[?��#�����IDq����>���?�#@�S�?�r�.��>������Du��@/�}��#����@X?�3(��g�>��?����6e�����z�v���>9��?�n�?ه�>12P?�p��V,�a�>%�K>KW?7�0?���>oa@��.�=�2?�9��<3��<X�'�_?��@�@�B<?�~����߿�����q����ƾ��=Ѝ�<��>%���i�=  =4�d�-Q��ӽ=���>gRF>�>�4>*,>�".>����a+��������ުP��
 � ��22�V� �52P����C��5���%�ѽ������\����p�Kw��Ǥ>16X?��$?���?��2?��=�o>n��S�ڽ4�˾�Y>���>�*b?��?�W?�R�>4Ǝ��o��L��lك�*���jF@>�-u>z?��>vS?b�����<�0>>L>E<>K8
>pA��m#����>�x�>�s�>���>sC<>��>Cϴ��1��f�h��
w��̽-�?q���R�J��1���9��Ӧ���h�=Ab.?�{>���?пc����2H?&���z)��+���>��0?�cW?�>'��t�T� :>6����j�`>�+ ��l���)��%Q>vl?�f>9u>M�3�Fe8�*�P��{��j|>36?綾�E9���u�3�H�cݾ@HM>�ľ>J�C��k����c��ti�$�{=`w:?!�?L4��{ⰾ��u��C���NR>�9\>6_=Ti�=�UM>/bc�J�ƽ?H��i.=���=x�^>�?�i%>�N�=���>�,���P�~�>� E>4>��>?k'?�~ּ�2��Ǉ�p8�Ġv>�z�>[9�>�|>[�M��=�-�>Gd>9��6�z�"���v:��Jc>�����d��Nc�Q$f=Q��0
�=l=�=�H��C=�{m2=�~?���(䈿��e���lD?U+?] �=O�F<��"�E ���H��E�?q�@m�?��	�ݢV�@�?�@�?"��N��=}�>׫>�ξ�L��?��Ž/Ǣ�Ȕ	�.)#�hS�?��?��/�Zʋ�<l�}6>�^%?��Ӿw�>��̽Ad��پ��[�h���=L`>T�1?D��e&�=c��@Gq>�??q`�β����ϿD}�/?�~�?��?�E�%U���*�]ҙ>p8�?�4R?\$�>�"��P"!=���>am?5<c?��>���1�H� �?N�?|�?,K>:��?�`�?t�>�&w�m%����q��/H�==*<>��>M8C=������+�tI��F#��I�h����8�>DY�=Y�>s�`��a��<�=�[&������=(�>��2>�E>$��>	ʦ>b�>��y>q��<.A���Ҷ������uK?d��?�b�dB�I=���<�i��܌�>m&?����aھW��>�T?Z1�?�Rp?l�>�1�៛��FǿY��� s��R[>���>k1�>/J˼�a�>��ƾ�v�l�s>���>?���LԾ���S����(�>+?���>C��=*�?W�%?�{t>��>��G�*����F�sԻ>M��>�^?9~?
�?�ָ���2��Β�3<��`[���I>H\{?k�?h�> ������#7�C�^����Wg�?�ch?��Խ>�?)��?�x<?�Z??��a>��v־Pu�����>�c"?G��j�B�K ��cɽE�?��?���>���Li����K�u�����N?_�X?Ԩ*?e+��y[�����o�<�n��۷��I��F/�c�	>̼�=�������=�b'>��=.�����S�1��<���=^�{>�C�=�B)�)���֫?T���@���>�3��D�g��%�>�}?l��[��?ag�=�/e�eU���l���U���8Y?�2�?s6�?!�=��Q��?��?U۽>��>CYþ��]�};7��x��F�w�O}��	�>�>�l�i��p���Tݢ��c��+սH9$�<��>���>��>���>�W:>WT�>�ב���-���_���P�e>&�=>��`8�����ϔ�M�����g�ƾ���H�>=}D��%�>mZ?Z�F>�h�>�}�>��鼈j>�vY>�Xu>���>�"t>�?>�(>�G+<�����KR?=���<�'�������6B?�sd?,�> i�C������-�?7��?�q�?�Cv>zwh��'+��l?�9�>���Uo
?K:=�f�{"�<R�����������Ӥ�>�?׽�:��M�tf�Qg
?�,?q_����̾�׽現j|>�+�?��)?�f<�K/J�i�l���\��F��r�=SR�پ7=�ti�Q���剿�ւ�A���v>Hu,?��?-��х���þx�j���F�w�>>� ?ak�>H��>?�t>r��e(�;�h���2�
呾#ȹ>���?ib�>ŀF?t9?�[S?�P?'0�>�˭>�����>�L�N��>ۉ�>4 >?!�0?O0?Í?�z)?ޒP>���B�����ھ�$?��?��?g?Z�?����"��%���G�Pq��!��WB3=Q�<�}ս��D�M�v=�JV>n?�-��8�����]k>p�7?�>l�>Xt��n&����<}��>�q
?�Џ>+n����q���[H�>p�?R�]'=�U*>�i�=�5����<�>��=�~��-ؓ=�����8�#7<nu�=7��=�{��p=h�2U�:�Ȑ;ҧ�<�k�>f�?71�>9�>_p��#� ����1e�=7X>r�S>��><Uپ�{���&����g�Gxy>���?炴?j�g=���=���=d/���	��w���?���a�<��?�Q#?�hT?J��?�=?*_#?R�>#�>Q��K��iM��t�?w!,?��>�����ʾ��։3�۝?i[?�<a����;)�ސ¾��Խұ>�[/�i/~����>D��텻���V��6��?�?JA�W�6��x�ۿ���[��{�C?"�>Y�>��>U�)�~�g�s%��1;>���>lR?���>��i?�:|?�/Z?���=�JI�o笿�-��y������=v*/?x?|��?���?)��>�c=[�����d�$�n���6J�l ��ϧN�+'�>�b�>��?_X�>��=D,�ׅ��O�i���6>�f>�K?��>���>`||>�@"���G?���>�b�����⤾Y���ə<�;�u?���?ƌ+?�(=�z���E��7��bQ�>vo�?���?'2*?��S����='�ּ�ٶ���q�z�>�ɹ>�$�>ḓ=]+F=d>U�>���>,�|[��i8�N�M���?�F?�{�=��ǿ�:������h��b���襶�������>��<��¾�ʬ�ߢe��4��p�Ӿ*������Ʈ�lhL�y��>~�>�9�=\)�=���=Fp�=�E���g�=I~��oR��#���>�;W����zW��r}��}�����\r�����m�y?��Z?��:?O�C?�[Z>i�=����x>�'���?[�Z>����p���4*.����/󹾗%�M`��R�.��z��=��~�|Q>}4>|>g=-J\<dy�=�5=���x�(��=�]�=/}�=�<�,U>��> =�6w?X�������4Q��Z罥�:?�8�>h{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?>ti��d�>M���㎽�q�=I����=2>m��=v�2�T��>��J>���K��A����4�?��@��??�ዿТϿ5a/>mJ">7`�=��F�rB9���p�"m���(� ?ҀH�g������>���=�c��J���.�y�/>_�=����Q�(�-=�v���v<�̈́=3��>X�U>��{=m҃�&#>�%�<0u�=# d>8t�S�;:O���	�=���=��Q>��0>
��>H�?X,0?tld?H�>��l��DξU���u��>��=�ʰ>�ʈ=� D>}��>��7?U�D?��K?��>�=bǺ>v�>��,�>�m��h��J��A�<Ol�?`��?ĉ�>�9O<F8A�����>�Vǽ,?X=1?�l?⿞>>����~�%�g�.��q��ژ8M�(=Gzo��3S�����,���_��=�=���>c��>&��>`�z>�;>��O>��>ќ>5��<��=2F���ο<HZ���1�=
鐼�"�<�K����!�B9 ��+������;�H;�.O<jS�;�'�=�f�>�dB> >�h콱�۾��>�4'��|�(�j>�;�<y���܃�����\5c��8I�b��>:�>x���������>[ĳ>.)��V�?_s�?oe><k;�	eǾ�����S����e<����nmr=���a�U�Y�t$X���ؾ '�>^��>��>|\>�L,��G>��f�=7ݾ�'6��7�>`傾ސ�H4+���r��k��;9��-Fd�q�y:KgC?�͇����=E�y?MEJ?e�?��>������Ѿ��G>4���<���JJn��?C�6j?b�&?�J�>��辆�@��1ξ���{<�>�da�@�M�XM��y�2�i�T��7��μ�>� ���h޾�.�=���A퐿�`H�������>LvP?�خ?�?Z�� ����M�_r���:�
;?��f?���>I�?�	?��Ƚڙݾ6�q�Bw�=��l?��?K"�?[�+>� >���!��>1N?��?K?�?,?�<����>���*��=���;��>6>y9�=��>>$�?���>��>}B�������#����CM��Qi=��=v�>E�>��R>�=g��:���:$u>�U�>R�>S�5>ߣ>T�>�}ξ8�8F ?�%����>>�?xx>��>�S�y�;�z�=ɘ4=:�����a� C�˶�=j>f>XZA>��%>+O�>}���{�?I>?�'���?�}�q��=�"�>�a>u���V�>��?!�>�F?l�k>8�&>��>�A>�+���(>7��F�L����K�������=vü��J��RE��ᠾ}jL��p�s4����e����8�b�.=Ȏ?�(�Dew�o������>?U�_>�?�Y����,>zb�<�@&><��>)���C��o*��B������?V\�?:;c>��>��W?��?�1��3��uZ�`�u�)(A�we�*�`�፿꜁�t�
����s�_?��x?�wA?=�<�:z>��?�%��ӏ��'�>�/�u';�,A<=�*�>Y*����`�˯Ӿ׺þ�5��GF>��o?�$�?XX?TV���|=g�>;-?a�F?*%�?��8?��C?����f&�>9�*=�R�>֭?��O?Y??��?�>��>?砽�W
�I��� ���Kp�95�X���̶=(>�g>=��V=q�D<�sY��!���y��]K��������<���=�B
>���=���>N�]?�G�>*��>��7?����o8�ˮ��%/?�9=����������r	���>n�j? ��?�_Z?�Nd>��A�]C�r>�Q�>yi&>1\>9e�>�j�r�E�]ׇ=�G>�V>ک�=D�M��ҁ���	�2���r�<�+>��>�,|>9��4�'>�x��W'z�(�d>;�Q�˺�\�S�j�G�J�1�v��\�>��K?��?w��=�]龷4���Gf��.)?�\<?�LM?P�?���=��۾/�9�/�J�Q=�6�>��<I��/����"����:�W��:��s>�2��_Ҡ�Ab>{���d޾��n��J�޽�� M=���DV=x�t�վ%�~�p�=!
>Ů���� ����Ѫ�#&J?��j=r��FU��[��Z�>���>�ܮ>��:�s;w�ɂ@����� y�=���>��:>�m��r��uG�r0��*�>�'e?Ӏz?[��?u���p�g������~��~��C?��>@**?���>��s<D����"�0�d��P��;�>I��>��?�#��_ؾ�-	�j�8�<:���K>df=>P1?K?��?��]?��'?i�>}�o>ޣ߼�v��a&?4��?�v�=O�ҽr�T���8�?JF���>��(?T�C��\�>�?BD?�y'?��Q?21?�>,%���@�0�>�~�>wW�5����a>UK?h`�>inY?���?��<>l6�����]��2�=;�!>��2?#?q{?{a�>�	?C���yº]��>�w?��?�#w?�`>?')?Fˋ<�h�>���>O��>�%?G�8?$�<?��j?D�C?,��>[� =����k��"��iiƽ��n��=\��<�U&<}Y�=�=?M=sP\=��==��<�!<�������C_�>��s>�����0>H�ľIP��7�@>�����O��`ڊ�ލ:��ݷ=��> �?P��>�Z#����=l��>�H�>���W7(?I�?�?r+";R�b���ھp�K���>�B?���=w�l�:���=�u�i�g=��m?Q�^?ƗW�C%��q�b?H�^?�*�ܹ;�u�þ�d�w뾃�M?gY	?H,J�v�>A�~?��r?,? ?�_�4�m�㪜���b�5�p�~��=\��>N��e��֟>z99?�0�>�Yg>f��=�R۾�Oy��蠾�?�5�?��?���?a�+>�o�s�߿�,��
O��s�]?X|�>~)B ?���1Ͼ�����	��Ly޾�ۧ�AA���F�����;8%�p���W�㽐/�=;?��t?y)n?��`?����b�� ]���~�1�T���e����E���C���A�Kmq�yC�������Q=�r��>��9�?��&?M8�A��>Þ���;�'�ξb@>�i��>���k�=F���d�-=0�d=�s���=��)����?f��>���>v<?��U�>A;��1��|3�����K)$>�H�>��>K��>Z}�;-B����O̾=���Oǽ��>`�k?GKS?^�m?�i����#�՜r��Q ��g��>�Ⱦ�r�>H*H>��>
X��8(��4��tK���e�|
Ծ~����<��^�=�6?2t�>��>�?0��>����ھ�w̾imP�ڤ��NĎ>[cc?J�?Q�I>
v콅�%��j�>I�?�?���>A����g�U�q�tPƽB�?��>�J?�?U����#�x3��Fœ�;�=��;��?O2�����!�x>��`?^�>d�=�s�>������a�Te��ۚ�Iǌ����>��->��=��׾�:�F�6�&y���N)?_�?:���*�\�>�#?ȍ�>ȣ>�>�?+Ț>l�¾���:�W?��^?^GJ?^A?���>��=�O���	Ƚ�(�ޝ/=��>(GY>1wp=� �=W��"]��z���B=���=��ļ�����#<�鬼�M<�	�<��4>�`ۿ�`S���ݾ���C������#��L֢�lȋ���-����c`��J�m��bý@ ��%b���\��_������_��?���?]Y<�����ί��CԂ����N��>U�4�kO <���9�K�<��a��2j��5��H,S��Ff�}<�;�'?����߽ǿ�����:ܾ"! ?�A ? �y?��-�"���8�� >0B�<�-����뾧�����ο�����^?���>���/��P��>���>��X>�Hq>����螾�2�<��?%�-?��>��r�,�ɿ]����ä<���?+�@tA?��(�H���V=���>B{	?�?>rV1��K����U�>�4�? �?�eL=��W�V�	��\e?���;��F��x���=f �=�K=ê��vJ>(2�>f�wlA�"�ܽ��4>�ƅ>6b!�����^��@�<�>]>Ԥս���k̅?��Q��k����*�|
����=..~?P�?�Չ�!5?%�F��M׿��g�n8?��?L��?x�B?:�彮��>������6?�*9?0��>_J;��Ѝ�!��>�OC�v� ��W�)W:�s�_>�"t>We>�=��6�;�U�)����l�=r �%�ĿȐ$�e���0=q�<+ĵ���׽�Խ,�� ҏ���[��#뽁�=#��=*�$>Ep>��->��=P?�v?5i�>E��<��>�[>����־q�9���E��C�����X���������-�˾*��������솾�!=�7׍=�*R�����P� ���b��F���.?��$>��ʾ:�M�d~+<�uʾй�� "�����0̾2�1�7n��ǟ?d�A?��u�V�m�<���^��*�W?~>�;��䬾X`�=�U���G=��>?W�=�� 3��hS��p0?tQ?_��xJ����)>���=��+?=�?��[<.�>�J%?8�*�\y佹H[>s�3>츣>p��>�'	>���s2۽��?�T?����������>�R��N�z�"i`=w:>�5��v�ѯ[>��<����1�W�6_��Aa�<�'W?<��>;�)�F� b����B==�x?"�?J2�>}k?�B?s�<g���S�C ��Pw=��W?�*i?^�>�����о~����5?��e?I�N>bh�m�龮�.��T��#?[�n?6_?�����v}����w��7m6?��u?RI\�>�����S��>�)�>���>N�:���>�j;?9�.�\?������x�1��ʟ?~!@���?Ǝ�;f �(�t=���>N�>��X��,���.��'����mH=#)�>8����3x��0��1%��<?��?���>&��������y>����k�?��?Eث��H��
�ib�Fu�C�<���=v�X�T�=ǋ��|�<�R�žm-�g��>c�zKi>��@��å�>�C����пw�¿����������h�	� ?�~q>3����˂�%n}�	�;���3���[��N�>G�>�Ҕ�������{��n;�eo���>�1�d�>�S�+��᚟�=S4<F�>��>PĆ>����轾�ę?fe�� ?ο�������0�X?h�?7o�?Wm?-w9<��v�F�{�z��{-G?��s?Z?�_%�&C]��7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*���+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�^�_?'�a�T�p���-���ƽ�ۡ>��0��e\��N�����Xe��� Ay����?M^�?n�?���� #�k6%?"�>n����8Ǿ��<���>�(�>o*N>I_���u>����:� i	>���?�~�?Kj?���������U>�}?S�>��?��>�F?:��=Q�����;�&>"o>Mt����?DdE?xg�>�>�yR��I-�(?F��nR��>�v�7�Ҭ�>zRY?y�H?�8>���7���!�����a�(�X�d*��ˆ��Ї�4/>��H>_n/>W�g� ݾ7�?�g���ؿso��Wo'�)4?���>��?���J�t����&_?�g�>�6��*���#��*5��?�B�?��?ϝ׾ϼ��>s�>eQ�>�ս3z������0�7>>�B?F�C����o���>���?W�@�خ?ki��*�>��˾ ���󑒿���� :E� ǽ�GJ?;Q;/P�>��>�7��j�������k�S��>��?���?���>��q?�tY��ex�ý)>o�>��|?*a�>=��>Ճ(�c93>�W?n���k��|M���w? _@�@�O?M���)Կ����Fվ[�����k>i�9>�q>?��Q]��������!��Z>��>�rq>6�">�&K>kM�=��4�J��U�%�/ ���H(��a��BM�V�½���������Ծ0ۨ�%u�d͛� ?��Tt��1���ل�t�A>}�_?_?*�`?Cu�>F4,��=!6쾗���Y���Ȼ�R�>F�A?�V?��L?��=d����y�ʢ���B���O�����>v��>1�?*4�>.�>�[k�s�>��>�}�=���=,�=�Ҡ�tr�<Svy>�p�>��>�a�>rC<>��>Fϴ��1��f�h��
w�a̽0�?����U�J��1���9��Ϧ���h�=Hb.?|>���?пf����2H?'���z)��+���>}�0?�cW?,�>��t�T�>:>/����j�%`>�+ �zl���)��%Q>vl?�f>��t>Qq3�G8�E�P�h���.l|>�6?���9�ߡu���H��0ݾ��L>ꪾ>iB��i�g���
��ri���{=�l:?3?�Ҳ�°� �u��0��:R>W�[>��=0��=5N>��b��Mǽ�#H��*-=h�=	�^>���>Ｆ=s�B>*��>�ô��f��£�>i�=E�=�2?��?ڀP<��=�����7�>W]�>~��=�B�<bJ��L=7�>T�I>�{<��{���o��� ���>=*�̑н�s>=���>�!��3,����[<[�V��5U����=�~?���$䈿���d���lD?V+?x �=��F<��"�C ���H��D�?q�@m�?��	�٢V�?�?�@�?��$��=�|�>׫>�ξ$�L��?��Ž,Ǣ�Ĕ	�%)#�fS�?��?c�/�Wʋ�8l��6>�^%?��Ӿ$h�>�x�vZ�������u�K�#=��>�8H?\V��)�O��>��v
?�?�^�ީ����ȿ"|v���>J�?���?:�m��A���@�j��>$��?�gY?poi>�g۾�_Z����>��@?�R?��>�9�{�'���?߶?ӯ�?��\>r�?(g?8(�>Pc�<�V������|�n�>
�;>���>g�_>V{��.�q㟿܃�5�\���T��>�%�<o�>8t��G��ES�kq7�����=P�?���>$6�>pf?]��>��>ڤ�>��<h'�<
,$��Y;EML?�A�?�	�di����<9�=��`���?@3.?ҍҼ��о�Ū>·^?3��?�J`?&v�>�������������w�;DrK>S��>���>mV���O>��Ӿ�3�H��>�#�>vV��B�׾󣇾f/��)E�>��?���>���=;H?r�.?��>$�>�_6�|���ԁJ���>-�?zy?�N�?��?0ŭ��M.�'q�������W��{'>�=�?�\?�d�>�҄�	}���?ӽ�ۼ,Px�Y�?��k?G �<{'?Aʑ?e�=?��;?���>������;��Ζ�>@�!?3"�M�A�@D&���v?cO?G��>F��.�ս��ռ=���j��<�?("\?�?&?y���+a�`þ���<�]#��zR�3��;+D�,�>gm>;p��	z�=��> ��=�.m�l�5�gg<�:�=w�>���=�47��Q���}5?����7�ݾ�� >{���'l�*�.?�f�>������?�«�����I¿/��C����G�?0��?��?�^>r�Y��8(?���?�^�>���>�Ⱦ\��f��Cw3�A �@���0й>/�>#���x �Y���������}����U7�>#�>v�?;O�>3(>��>hx��y�%���˾3& ��:R�hW��
=���#�������;�s��ʚ���������> �N�aú>5?s�2>�->���>wEY�5~�>�m�>Ib�>#��>-�u>y]]>��=�z_�Z��LR?���ؾ'�ĵ�鯰��4B?�qd?�1�>+i�+���V��9�?���?us�?�@v>~h��++�|n?I>�>����p
?rG:=�8��,�<�V������1����A��>T@׽�:��M�lf�gj
?y/?����̾R=׽w����=��?�w9?���I�!�[�(�V�!J�pH��M��˒�E���Zj�!���V���m����)�]Ӷ<#?|��?7#��?K��9@��H�5�:�w��=%�?���><�>AQ�=��'�[���py�QM/�c�N�|��>��?쎍>6yI?B<?6qP?�TL?���>Eg�>�<��cR�>1��;���>��>�9?��-?�00?�t?<\+?��b>.���������ؾ�?�?�B??֙?!҅�"Cý���\�d��gy��(���1�=���<d~׽�u�vT=0T>>W?<��u�8������	k>Z7?7z�>���>l���,���a�<0�>��
?�=�>�����rr�8b�B�>{��?�O�=_�)>f�=e���Ӻ�%�=������=���k;�u�<���=��=�{��k��W��:ٽ�;>ï<jt�>�?���>�B�>`@��)� ����Kd�=�Y>XS>v>�Eپ�}���$��z�g��\y>ww�?�z�?�f=��=3��=�|���U�����n���;��<�?J#?XT?K��?R�=?hj#?��>�*�OM��^�����Ѯ?Y!,?���>*���ʾ���3�ܝ?+[?�<a���f;)���¾\�Խï>�[/�/~����!D������������?Ͽ�?�A���6��x边���I[����C?�!�>LY�>��>��)�=�g�S%��/;>?��>�R?���>̆q?���?��M?9|�=��8�@���������Uo<�d]?{x?��?�n�?�`?9�=!|��`	�� %�7�Fk�����E�&ë>��?���>���>x]�=����^о_�v��L'=�<>�?q��>~N�>�w%�kU+�V�G?+��>Be�������"ă���<�Ϟu? ��?*�+?�5=L��"�E��G���O�>Iq�? ��?�6*?��S�w��=D�ּ=ݶ�M�q�y�>SϹ>?�>���=�oF=�m>��>��>	0��\�+r8�2eM���?�F?���=�+���0`�̓�M��vc>\o7�:��Fe��}��=�B��#����F� ľ )���b�(S���¾�K�[��3��>�!>��>X�!Y=��̽�,��bu<:�0>��>����n2z���;�����U�������<"�>4�>��Ⱦq�}?V�I?�?,?��B?&�t>�I>�N)�5@�>A^��5?#3U>`r;�h渾�\?�^���\��0�پyվ�a�%&��K>�>G��\	>U�*>�w�=��<��=�h=�ӕ=���-=���=��=���=+,�=��>>�>�l?��Z�����2�c�~�7��i4?��6>N�?,^���:?��,�OT��Hh���UA���?�x@�'�?�L?>���$��>Y.��Ƚ��c>͜���
,>�g	?N�6�ũw>��>-�������b��t�?!��?�T?k鋿퀶�^�>��7>�,>�R��*1�k0]��c��Z�$!? ;���˾p'�>ɮ�=4޾��ƾ�i-=��6>I�]=
Y��$\�{�=�(y���;=PIm=��>�mC>���=Y����@�=�]E=��="�O>�5��_6�o^3��N.=�~�=4fb>�b&>��>��?b0?mXd?z6�>n�aϾ|?���J�>p�=
F�>��=�sB>3��>+�7?ȳD?��K?���>Zŉ=T�>�>^�,��m�Dn�;̧�F��<|��?�Ά?aӸ>�R<E�A�����e>�N,Živ?3S1?�j?2�>F7���ۿt7�����=��>��=��ŽJ��`���΢��'Q���=K��>-R�>�V>�OF>��=����|x�>��=�t�=�a(=��i�-�p��A�n�zX��v+=�)	=��;�ѽ�:C�`B��Vr};�	g<fD�=�כ=E>���> 	>�ܾ>���o߾�y�>s�s���[� @`>����>����'��MU*��,�/�.>�u(>�/��Z䆿�u�>���>:\>ы�?��v?w�=�gc�`��?���AM���Խ�ӊ>G�,>ZO�G1+��zq���F������>�0�>�.�>^m>",�>N?���=�y���5�c��>�{��^!����Bsq��䤿ꃟ�i�h�X�'�H�C?�퇿�.�=os~?�I?L�?ӈ�>8����پ�L3>�#����=���Зh��卽)�?��&?"%�>^��'E��˾�D��l"�>����=>@�uq��-.7�&IʽZ�0����>�k��%����(�\o�,͐�RCA�~9V��3	?�L?�?q���c����I���ھk@ܼ���>)f_?�qJ>��?�^�>F�b���A�޾BG.=�Ua?;��?c��?�>+0>[�N�?��>ڊ?��?tt�?�v?�Ͻ��?%� ��ǹ=b��=��>�ғ>�/u>s>r?&?��?s!��M��7�Lþ�ǆ�?%�F�#>8�>3]�>�H{>���=�b=K�b> �>x��><�>��>��>�>*��<���'?���=�0�>wM.?IF�>�C1=87��z�=y�O��<�S*��<ͽQRڽM��<bB�n�+=Y�����>��ſ���?�O>�����?���*�D��F[>7�K>>�ʽl��>��f>F�>�#�>)O�>�->���>��&>��Ծ,m>p
��%�:�@�XqQ���վ�Ep>����(�#���
�%��Q�M�uδ����+�h��)��I�7��F�<
Ď?E� j��)����F?Dz�>D6?���
i�F�>���>8�>�����:���!��b�پ$�?2�?�9c>+�>=�W?Ƙ?�1��3�vZ��u�'A��e���`�u፿՜��ї
������_?$�x?�yA?�f�<�;z>I��?��%��ӏ�*�>/��&;��L<=�)�>Y(��*�`�t�Ӿ|�þb=��GF>b�o?�%�?�Z?�SV�P��<5U�=�0?��(?0!�?�a?$F5?����5?�V=�
�>i�?��?+6?Z?�6>��=���-�C=r����Χ��zT��C��e(��Eo�=�'Q=ު
�ki;���<敘���;۟=5�=�=Б=�Mj=�?�=��>޽�>0�]?N�>���>+�7?���v8��Ǯ�*/?��9=2�������Ţ����>��j?#��?;aZ?S^d>��A�		C��>;W�>Pn&>�\>)`�>�m�Y�E��܇=eP>m[>��=0_M�ҁ�C�	�U������<�(> ��>!�z>���t�(>gӣ��&{�ȯc>}�Q��m���HS��G�1�}�q�k��>b�J?fk?U�=���'Q���e���)?�;?u{M?И?I �=0�۾�x9�zkJ�T��N�>�w�<<S�=��`���A;����s>LV�������ya>'��I)�Cbr�mJ����ޛ�={}�!�<���o�ѾyD��K�=�>�M��Y��tA���Ƭ���M?	��=���]�C�����9'>N�>9ܱ>����%?���x>�R���A�=�g�>6QG>y9<�T �/�R����5>'�Y?�Zv?�w�?��1���c��U�V�s�����Uw,?kM�>��?bh>�;��Yc_�����a���3�U��>MV�>j��bD��uz���`H��i�>�5�>I)=�,�>�|?��*?/V?�b?�G?�x�>̰ȽȌ��'�%?�r�?$��=t*;�!32��b+����>��%?t��cv>(?9
?x�3?��\?P�?V�>R���*��i�>�v�>V������m>�N?���>��[?C5�?-��=n�G���K��Rd�=}�A>q6?[�?�.?���>]�>�_��y�=Vޯ>�9_?��~?3�f?L��=L[?In�>y��>E��<���>��>J�?�q/?��}?��Z?���>o��<ɹ��z��Z�^�&��[�a�&�k��7=�	��f?I������>�RØ���<�|����O�o0�$a��{��>�r>���IW0>��þ�j����A>����{K�������H:���=J�>��?�ٔ>�$���=���>���>/����'?v}?��?�[;5�b���ھ�\K���>��A?��=s�l�0����u���j=�m?�^?�W�{���[ob?c_?��m;�&���krb�8P侕yO?ʑ
?lyM�ϋ�>��}?B�p?�� ?��Z��l�����{�_��c��1�=�/�>܅���d� ��>[8?q�>~�g>v��=8e޾�y��#���H?�y�?w��?��?&>�Ho��X�� ���aS?4?�@ɾ��?���9k����Q0�@�����_���#6�ۢ���|��'�����
~�=�v?-�5?b?��~?���'K���H�8����J�#�t���wgJ��U@���B�Ԗu���	�˾*�G��w*=��w�̭C�Б�?�0?�N�#��>a�����O����M>9���0�*��<�=�g	=�D�<Yo�!;��覾|�?ϓ�>F��>�/A?��Y���9��L*���8�S��\>䲢>>�t>�Y�>ċ��(G��u��������o�cͽH.v>1wc?�K?��n?�8�N1�f�����!��'0�KU����B>�>2ɉ>.~W�d��Q3&��O>���r�����z�� �	��)~=զ2?�*�> ��>�P�?�?�	�_h��VBx�8�1���<?�>ei?f�>�>��ϽR� ����>��l?Q��>6�>m���|X!���{�
�ʽ�&�>@߭>���>_�o>��,��"\��j�������9��x�=��h?]����`���>iR?���:��G<�v�>��v���!�G��m�'���>�|?���=��;>�}žs$�E�{��6��I?��&?��y�� �И>5�?�B#?���>��t?�J>k����r���?�fn?�h?�nF?��>�?<W@U�A(ֽT������<�|G>S�y>^zT>T>9��r��k�o��<k�	>��ҽ��M��DO�=�S/,�����K=Q�޿�6O��I޾8�G�龄t
��3��.ɘ�����E�0�U�Ⱦn���%4���D�Ř!��KM�f^��䋾�Me����?�g�?�e��6ꕾ���[�{������>�5P����gr�����46����ؾ��j��fM�~f�H f���'?!���s�ǿҰ���?ܾe ?�? ?թy?�H�"���8��� >�K�<_�����W�����ο������^?���>M�)��8��>���>_�X>�Nq>���螾�E�<?�?I�-?���>�{r��ɿa�����<���??�@m�@?*.�z����=�4�>E>?'T>��4��n!�ԇ�����>X�?HΎ?�Tg=�fQ��r����j?�r4=ߪ5��*�I�==�F=�Y={�	��):>0ƍ>/��
�K����.6>���>����p}��1M��hĻ;eR>u�ɽ)��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�����{���&V�}��=[��>c�>,������O��I��U��=����ÿ32'�_s��=��� ���U ��]��uQz��O�3������H�f�=!dF>��t>��;>]�N>a?�K�?�>H�@=p�����֯�faU>q���v�tCо" ��2?�P�� ��\��$�f#�*`���B�k{ �מf����ԟ=�q6}���o��a?P}�>���:g�%�~=;��}.0��ny������HK�#V���������?gx!?�`K��Y=�	��C">�����B?���4�󾓣I�#�Y�g���+>ʧ�>�T<Q����j���o�y?0?�?͇��;o���,H>�%����=��%?&?��]<�g�>��&?r7:�]�-E@>q�!>S�>��>��	>�*���m��/"?c�W?�Iὀ萾��r>�j۾��w�(K�=�$D>%]�l'���L>B�̼8׊�������u���=�W?�5�>��)�!����*n�&C=�7x?��?��>�'k?e�B?	~�<u����PS����À=�W?6gi?�t><�����оk���]5?Ee?��N>l�h����9�.��	�(?v�n?)s?������}�ݒ�I��NJ6?��v?�u^�dm�����!�V�H�>[�>���>��9�|�>0�>?r#� ?������Y4�U��?N�@���?L�><sD�6��=�4?�X�>�O��Nƾ�����|��<cq=J�>7���Fiv����a,�D�8?e��?�~�>���4��g�=6>�N�?NÑ?W����3����w,����QN�=���>@�7�'�潐s��
�B�fBϾ ��ֆ���k,���=>�@���="3�>�Ҽ=��ſ�QϿ��J��������
?Щ�>�6>fփ���P�!�'��4M� ?<��7��}£>:4>����`��nz���:�ʝ��B$�>[��9҉>�6V��;��i����g<OX�>���>��>_h��Uƻ�?b�?6-��ο~H������W?���?m�?3�?�><�Iv���z�kh2�?pF?	ks?1�Y?6**�e^��?�NId?O;;�%Q���,��s$��p�>�91?	�>���Y�>^T)>�(�>���>�.��t��D��^���t"�?���?8U����>�w�?�)?�t쾯o��"��������=�D'?�c>1Oݾ�GE�t|:������?��?fc���~.�b�_?��a�g�p���-�g�ƽzۡ>!�0��d\�N��Ƥ��Xe����@y����?K^�?a�?Ͷ� #�*6%?O�>m��� 9Ǿ��<���>�(�>O*N>�H_�Ĳu>����:�vh	>���?�~�?<j?򕏿����V>�}?/�>��?���=*R�>��=^ΰ�U5(��I#>��=�V>�j�?��M?_@�> l�=��8��/��QF��;R���W�C�*��>`�a?�hL?B�b>�r��C�1��!�|ͽ>41�����@�|�,��q߽]95>�>>�>H�D�T�Ҿ9�?�}��ؿ�\���&��C4?�ʃ>��?���t�׊�^/_?���>�&�)���,��{�m��?&C�?��?��׾S ˼�A>��>���>ąս����lM��&�7>��B?l���V����o�M�>9��?��@�Ů?�i��	?���P��?a~���M7����=��7?Z0��z>���>I�=�nv�ʻ��M�s�{��>�B�?�{�?4��>�l?�o�I�B���1=3M�>��k?�s?Ro�m�5�B>��?,������L��f? �
@mu@I�^?/]hֿ����;N��6������=Y��= �2>
�ٽl_�=��7=v�8��<��5��=F�>��d>�q>�(O>�a;>��)>���B�!�r��W���]�C�������Z�P���Wv�Nz��3������:?��H3ý3y��nQ��1&��>`��0=�z]?�=?!1<?HX�>F���|�>�#�}��=��2��%=R�#>�c$?�K?p1<?���=o�ɾn�o��jp�+ؾN>���Ų>�^�<���>r��>��>
<;�> �F>�I�>z�.>菽��P=d>���>���>�ݺ>d��>��>%�G>���v�R��=΂��vz��]�?����B�x�n偿`�ɾ�^Ͼa�=�1Y?�В>�q����տ�I��q�e?n����&�
�P�+q =��?W�H?ޣ=��=��$x�.м������=7o�>�F��,H��d�K� >8u$?��a>�>�2�F|;�=�L�����(�>H�3?���O�*���i���H��`׾SHk>���>�2p<�o&������z��On���<�8?�?�,ݽ	J��^�p�=N��+aD>؃m>ށ=S��=�1>�0����⽉7O��?�=-��=�lh>�
?�K�="h =�#�>s�{���%��ѭ>�)%>"f>�E?��?-ē�Y8�/p�2�:���B>E�>�>�0>c�,��=t�>�de>h�ؼ$�?�}\<��T>�h��nK��@�����;�[��_[>r��=_���_6�n��~?���'䈿��e���lD?T+?c �=�F<��"�E ���H��F�?r�@m�?��	�ߢV�@�?�@�?��D��=}�>׫>�ξ�L��?��Ž4Ǣ�Ȕ	�0)#�iS�?��?��/�Zʋ�=l�6>�^%?��ӾPh�>~x��Z�������u���#=S��>�8H?�V����O�f>��v
?�?�^�੤���ȿ3|v����>X�?���?g�m��A���@����>:��?�gY?roi>�g۾=`Z����>һ@?�R?�>�9���'���?�޶?֯�?v�H>6��?![t?��> o�f�.��'��?����Wb=�_;�˒>m>����E�
�|z���j�A���`>��=��>>�۽T����S�=�k�����z�`��Ͷ>��k>�F>�]�>N7?��>��>�(=D����{���2�K?���?����n�=[�<P�=ɣ]��(?HB4?]la��
о
è>��\?`À?/[?�y�>���i*���ѿ�<s��ƫ�<��K>��>�T�>Y���T;K>R�Ծ�C����>mȗ>R���Yھ7���ٴ���>�Q!?���>��=ș ?�#?�j>:)�>�`E��9����E�)��>��>�H?�~?��? Թ��Y3�j���桿�[��<N>��x? V?/˕>m���҃���E�	LI�/򒽋��?�tg?OZ��?�1�?��??{�A? ,f>���ؾШ����>�9?G�޽�<�0�%��^����?��?�'�>��p���ѽ=Y��4�uZ�,?��`?�((?g��=�_�>h��e�<l���֗���;x�Ļf)>��>����*��=;�">�W�=�yZ�[�B��ۘ;�>�=��>}�=�88��U��+=,?��G�cۃ�X�=p�r�"xD���>�IL>�����^?Cl=���{�����x��T	U�� �?��?Sk�?8��;�h��$=?�?T	?~"�>�J���}޾P��Qw��}x�^w�j�>���>�l���<���͙���F��6�Ž��#��� ?��>��?�~�>��K>�A�>�����!���aF�z]������0��-&�`��}E��s[8�ܫ:���ϾW5o�~8�>�8�렾>��?��>ǐx>���>R�]��^�>]<U>�Rj>���>��q>,�W>H�=b�׺q�0)R?{ֿ�|J'�r��eG��h�A?R�d?D��>4La����ռ�D ?]�?%U�?&�v>A/h���)��?�d�>�m��
?��3=/�����<暶�����6��2v���>Զ۽�9�� M�06f�(X
?�n?<��C�̾e�߽䟾X�c=O�?Z�)?�A*�_Q���n���X���R����  c����6n%�«o�q叿�B���݃��N(�N�+=+�)?ۚ�?5���X��a��k�j�6X>���g>���>xB�>2_�>�	D>S��l1��|]�vm&�=��7��>x�z?��>�U>?��U?��\?�]?�^�>8#�>K:����>��~=�&�>�l6?P.?aR?}=�>��?|J?���>����A �<f ���?Y�?�.?��(?�?��i���N�g;����$���d6��Ws^>ذ�<�浾�)�;#�u=��!>?Y��&�?>���M�>:4I?� �>o�>I���Ş���U=�V�>֦8?M��>����%-���E�?��?]{y���=��\=��=G��<�Yi��X<=��TD\>�^̽2=
����;c~a=]R�=����>�O�E�<d;@w�>��?��>�D�>Q-���� �"��Y�=8=Y>�S>�>�4پ�|���!��N�g��Ky>Wu�?Yy�?P�f=��=�O�=�g���>��������<ʐ?�D#?�XT?ԙ�?��=?�g#?��>�0��I���Z��S
��ެ?
�G?
X>%2��ľ����6F��3�>��?I�]�op�H|C�,�1���Z�a��>� ���g������*]�jk��_�A�-GI�|�?/v�? Ь<�'0����}P���F־��?��\>=c>���>�Z��3Bc��E�N��>_��>O.6?a�>��t?j�?W`?Uu>�EH��2��l/��/�QI>�l?K=�?�o�?.:?��>4r?��aȾc��(e��T}�0.��JW<}�9>^�z>���>�O�>G��>x�=��
���<n��������>H5�>R?�Ǥ>B7>;�J?���>�CƾO��V㙾�.y��ڼ� n?�s�?��/?J<C����:�0���>�h�?���?�J1?��9��L>׸��=ľ`~c���>�(�>dڌ>��=%Г=�,>�T�>U�>�M���[�1��/@��
?�@?�b�=t�пi�io���־��P�_�վ�����<ѓt��4��ؾ�4�iYξ@b�(ܾ��ֽ��h��6�D�)��'�>�Y�=;�	=��=�TJ��/[��d�Jd>R��<:1<�#�=�&Z>
�Q=r=���=���=�g>L#޼�˾�}?�:I?�+?M�C?�y>C>?�3�C��>Dw��K@?UV>,�P�ǂ���};�K����"����ؾ�v׾#�c��̟��F>�`I���>83>�J�=�J�<�=�%s=Tގ=�TQ�d�=�+�=SS�=Xk�=-��=��>�Z>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?~�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>q��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ5a/>��6>�_>4�R��1��[\�ߕb���Y���!?;�e�˾�9�>;_�=*߾�eƾ<0=�7>�m`=R��#8\�B��=��|�7�;=�+l=n��>.�C>���=P��^�=��J=�P�=j3P>�椻Xk6�WL+���3=X2�=k�b>�J&>W~�>_�?J�,?�'d?~��>�7�+F���¾N�>6�=r��>�Ti=�-Y>���>�'?iG(?��D?j.�>�>Em�>^�>�A��wb�M����qm>�+�?��?�Q>�T�JV�<��h�{#�=�M
?L?B.�>2��>����%ܿ}'���2� Ԯ���/����<�\�N��Jǚ��K6�ޫѽ���=\b�>݈�>(��>���>]�K>�Y>:(�>st>4�/<v�=�~J�y�弤��g��=����Bu<���;�[=�9�<�!Ƽ+����b�/t�:��/=��4��a�=���>D�&>�p�>N}>=$	���l7>�M���4M���=�퐾��C�6�`���q�1�.�JxP���'>� =>��p)��<�?FGx>'>���?p?R>$����Sʘ�CG?��xZ��!>�Q�=�-*��-��\���G��ľ���>st�>��>�>+-�U�:�dx=-�׾u�@�S�>p*��W�A����J�|ƙ��R��e�h��ͽ�?u5����l>[�?�� ?1d�?��	?_Q=I����>w9��@>�0¾�95���3��+?�!?WU�>�.־1}�_�;Q���y�>��J��O������0�"8�*϶�=�>����4Ѿ�/3���������L�A�bq�dκ>
LO?�Ů?G�`��*��UO����숽�?+g?�>�?�R?&_��u��}��䜶=��n?R��?C)�?/]>�#�>�]̾��?'b�>���?���?�A_?w�3�;�J>��>B��<fk=�8x>Kh�T�p>�!�+�<?|o?�_G?s����P���9��鰾i�y�l�=�Ǚ>!�Ż[�>֖���T��^>MX�=&N�>�D=��>�z�>e��>�t���*徬�?���=�^�>P?�С>g�6���;=So>̬�=�#��5�i�A��<9<>�<�;��E���@�ݻq	�>�Pʿ�$�?�'�>���z��>���Ev���pg>@U>�x'�9�>�M=';9>��%>R�=n��>��>K9>�FӾ.>����d!��,C�T�R��Ѿn}z>�����	&���)x���BI��n��wg�vj�F.��Q<=�"˽<H�?�����k��)�����>�?�[�>�6?kڌ����$�>���>�Ǎ>�J��a���Iȍ��gᾢ�?7��?c;c>��>��W?H�? �1�3�}tZ��u�(A��e��`�[፿����
�8��Y�_?��x?=xA?hZ�<t8z>��?��%�wӏ�,�>s/�^&;��K<=n&�>�)����`�\�Ӿ�þo8��GF>��o?^$�?�X?�SV��a�hT&>��;?Ł2?�=u?�3?�N;?׿�~�"?.D5>e?d?��4?Jq.?�b	?�->SF�=�k��|/=u�������5˽NȽ��ټ��J="=�v�;��t:�.=om�<O-�����:*93�U�<�L=^��=���=�~�>�x^?n$�>
g�>��7?&��}�9���� �/?�G=�Zv����������2>;_o?���?�`X?'2f>��E�
rG���>R��>u�+>{i><��>����eP>��}=�>�2>�4�=�=��?���I
�r?�����<�!$>�?s��>����5z">ydv��p���>m��������S��Z���"���o��>)�:?)�?�p=zƾQͺ�y2m���?\�A?��B?�U�?(�=>�e��R�	��� =�-�>�>è������]�<�h:<=���>h�|����M�a>N����q���I����d~�=ɂ�5@�<����Ծ+���b�=�3>������]��������J?.�e=8D��=�P��׾���>���>S=�>��b����*�?�dy��v��=��>�B>%�F�#)����M�)��y�>hma?x�j?Jq�?8�z�~��&c�T������Ȗ���8?�D�>�?���>Sk>��?H9��f�J�P�c�>A� ?�D�8[M�]����O�q�=��a�>�?���=s"?&�a?�'?�OP?j�,?��#?��{>�#:�������&?S�?���=�n�.�[���f���>II
?�hy���u>�U�>�?��@?�i?l��>�>�̾�$��G�>�r>01r�}���`>]?�-�>�\?}�?��U=Uz@�������ۼqc�<�/j�dZ?D�?�Q?��>d�?'La���*��!�=��k?mf?ӴM?E8��ٗ>��>fW�>�=]%:>I>.�W>��L?���?��h?a�-?�P=�A�  �(����
 >n�>�4=�;�=�V�<j�x�U��u��o���S��
'L������ý@ӽnj�����>aVt>�|��%�/>�rľ���v�C>^{������b��"W<���=��>Zv?kX�>��#�m��=�y�>���>��ܤ'?�@?y#?k�;;��a�Y1۾�
L�<�>�oB?7`�=�l�5}��K�u�X�^=��m?��^?�fW����O�b?��]??h��=��þz�b����g�O?=�
?3�G���>��~?f�q?U��>�e�+:n�*��Db���j�&Ѷ=\r�>LX�S�d��?�>o�7?�N�>/�b>(%�=iu۾�w��q��h?��?�?���?+*>��n�Z4�7����~���$\?)��>{2��gO"?,�#�t�оԀ��U��?W��F���h��C?��G����*�W����ͽ�R�=��?�p?;�p?�Lb?�'��0d�^����*�Z��5������@��.>���B��m�7��i������t�G=_gy��K���?�
4?=�l�%�>0&������݌�.�9>Xn��\o���2=� �U&�:�OV;J=P�?�I]��mq?��>�?�>>�N?��d�,B��_4���9�3��m�>�Y�>� �>m?���;���ѽ&��\� Ͽ��v>�6c?�ZL?�4o?Y����0��􁿗U"���;�����g�E>ch>Ef�>�M�m���/&��&>��r��"��f���/
���w=�R3?�Z�>���>��?��?��	�����z�|��s1�5�<�߸>�ri?E��>��>�kϽjR ����>_�l?	��>��>B����Q!���{�ٞʽx"�>��>V��>�o>��,�U"\�<j�������9�ň�=��h?e���g�`� �>�R?��:�QG<gu�>��v�E�!����,�'���>�y?���=j�;>�yž�#���{�4���v*?��?'r���.&��q>s"(?��
?��>p��?ܗr>Oվv*8���?�Y?<C?0�,?��>i�=G�������7�[4$=�cW>RNY>�>�=/�=�����.�y���<3<�=]�E��
0���Ƚa��SsZ=M�=+ba> �ٿ�]U���ݾ���{B����&��8���ԍ��>�r�̾+<��x��K��螽2S��_�҅���du��n�?���?�夾���0�����k���1��>Ҋ������U��������|������zվ�k�U�3�-RW�\q���'?a���Ȼǿr���o8ܾ�" ?F ?X�y?W�֠"��8�`� >.��<�휼���\�����ο������^?��>��.�����>O��>u�X>�Hq>����ើ=%�<�?]�-?��>�r�O�ɿۈ��"�<Y��?d�@�hA?��(�2^�	+S=��>j
?�A>4�2��dɯ�*��>�ޞ?+��?r�H=��W������e?<�.<��E�%ۻ��=b��=��=Vj���I>5ɒ>S��1?��޽�1>nq�>�C&��7�"_��V�<=\>Kսvߗ�5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=cI��Wؿ�*�-�+�����\��k���⼢?�@ �����񤆾| ֐����=�R��P��=Z��=#9>>�T?��o?��>R�<>#�������j�,>����Տz��g�����������i�����ԛ+��1޾��0�T��<�U}��V����(�{�k��?r���o?�4>���MWI�`c*=�u����#�f�;��xw���4�������	�?��C?X3���,Y��`7����=a�@�^�w?�s�^�$�b&���.�=� ��
����>�%>Xֿ�3O��􏿝�2?�
?_����z���'>ϰ���4>a*&?��?n#��%�>"?Wr�{���>�<>���>`m�>�'<>Ȥ�d.���)?�.X?�ռ�}����b>G���օ�Ä+>��,>���۵��m�7>��"��.���0=�yԽ�=�'W?���>��)���~Տ�^+�h�>=:ux?;�?�>,4k?��B?œ�<z����S�8�
���y=0�W?�2i?��>�̀���Ͼ����!�5?!�e?m�N>��g�%�龒�.�ɝ��?��n?>&?Hu���X}����c��16?��v?�r^�1s�����U�V��=�>3\�>Q��>3�9��k�>��>?�#�jG��Ѻ��zY4��?g�@V��?{�;<��W��=�;?\�> �O�^>ƾ|��$���ݒq=Y"�>*����dv����@R,��8?���?R��>��������=?Kn�pѥ?oە?[�Ѿ�0{����G�v���*�?��<*�>��<>�'<��ʾM4�,a߾�("�z`��5N>���>�@�Q�=���>����I1�r�ֿO����,�����+4?}n�>r5$=��Iw�� k�c0n�3�Z��Z�i�>�X>�B��9�����{��D;��Y���"�>�^���>��S�8��gO��S�D<	[�>�f�>˨�>C�������ʯ�?�4��<Cο{���E�`�X?p�?�n�?Jo?��-<�lw�^�{��v�^�F?Fs?9�Y?�&��\�.�7���j?cQ���`_�O14�ΙD�&�X>V�3?�'�>
�,�.-u=�>9��>�>��.�
jĿFn��?��1�?;�?9��W��>���?��+?)��O����	��̓*�A���A?��3>�����"�2�<��/��^a
?�0?ah��%�[�_?�a�?�p���-���ƽ�ۡ>��0��e\��N��1���Xe�
���@y����?K^�?]�?ε�� #�a6%?�>_����8Ǿ��<���>�(�>L*N>�G_�Ʋu>����:��h	>���?�~�?5j?���������U>��}?��>�=�?��= ��>���=	���^x��(�>�D�=�Ռ��
?;cK?�r�>	=nSC���&��E��zV�����E�j��>tb?RyC?�6�>8Cw�E��Or��'�K�.��f�;������}ܽ1�:>�4>�>E%�J�����?Ap�.�ؿ�i��p'��54?R��>�?����t� ���;_?Uz�>�6��+���%��zB�^��?�G�?7�?��׾Q̼�>5�>�I�>�Խ����X�����7>+�B?8��D��w�o�O�>���?�@�ծ?Pi�0	?�_P���`~���s7����=d�7?�.��z>���>c�=Tnv�������s�j��>DB�?<{�?���>u�l?�o�a�B���1=�K�>�k?Is?�o���*�B>v�?��&����K��f?	�
@uu@��^?��k�ٿ^���!O���wݾB�=�-�=m	>�ܫ��Ƥ<�7�=ʃ>'��=2�=1��>���>�X�>�r�>sK�>@�V>OG��*5%��䛿h��Mj?���$�)� �0�]�?����Ҿ̊*�w\������۽��ݽ��\��qc�n����R����=�JP?`�K?q7d?���>:�s%>�����[=qW+��=��>�N<?��A?,R.?&�=A߸��b�/t�h���v�����>aP>��>t��>Uڷ>���=��>E�>[�@>�֍=���:��o:@l�=>�H>���>p(�>|��>fHk>��>fXƿ�չ�J����茾����"��?��ž�ތ��t��8º�hJ�a�?�4?
�y>�b���`޿kÿK�E?/����ᾴ��:"�d<+e?�x?��=Qh����ɻ���=���Vj���1�>�kd�������Q��	<���>+f> 
u>+�3��h8���P�e���,|>N 6?[Ŷ�A�8�:�u�A�H�sDݾC�L>韾>�t@�[l�[�'���i�=�z=;w:?Gk?$��7ð�Ĝu�X��K�R>�C\>��=��=�M>��b��Ž��G��8.=7��=_>�2?�H6>�=>�J�>K�k�]���P�>t�B>�";>̓<?�?�,�"�2���q��f>�X?��><�Y>�@�V�=7�?(��>��_=<t��0�5�_U��[<>��=ѩ�	�=2-�<
��%�F>���=x�Dꑾ-S=��~?q}��.㈿���d��[mD?#.?��=xG<z�"�����K����?��@�l�?]�	���V�$�?�?�?���ۮ�=�x�>�ϫ>%ξ!�L�@�?��Ž7�����	��/#��Q�?X
�?� 0�ˋ�ml��8>N_%?��Ӿhh�>x�sZ�������u�ڹ#=���>�8H?/V���O��>��v
?�?�^�ǩ����ȿ|v����>A�?���?Z�m�vA���@���>0��?{gY?+oi>�g۾`Z����>��@?�R?y�> :�W�'���?�޶?ٯ�?�I>4��?.�s?�h�>W�w�X/��3��蕌��\=\�[;�Z�>:Q>����rfF��֓��h��Ȼj����^�a>��$=��>:F�b2��$)�=��kK����f�۪�>g/q>d�I>�V�>�� ?�c�>4��>S�=�u���߀�i���o�K?�?����0n�cB�<׸�=1�^�9&?9I4?�\���ϾΨ>��\?:��?s[?�[�>+���;���忿�|����<��K>�'�>�K�>h���TIK>�ԾD�Ul�>�˗>�ƣ��<ھ�7������h@�>1e!?R��>I��=� ?��#?w�j>m(�>�`E��9���E����>���>�H?��~?��?�Թ��Z3�����桿��[��;N>��x?�U?Hʕ>L���Ѓ��tE��GI�����N��?�tg?gR�l?%2�?�??Z�A?�)f>>��ؾ𨭽��>j�!?5��/A�z&����W�?�P?��>mM���pڽ�`�
��8��ش?��[?h%?o$�N�_�2���cC�<�<�7U�����;�[A��C>!�>�ӈ����=/�>m¯=u�k��6���<���=��>Č�=�G4��܇�?=,?x�G��ڃ���=��r�wD�o�>vIL>T��Q�^?Jm=���{�d���x���
U�� �?ݠ�?<k�?`����h��$=?	�?{	?�"�>0J���}޾ǔ� Qw��{x��w�Z�>���>#�l� ����������F����Ž�����?ݻ>�s�>�?� h>���>4���:� �O ˾���=,T�j��#�9���.�4��/����m �.#��f����i����>!�y�Q��>�ܲ>%�3>?Zq>��>6�)=���>T�W>Eυ>�u�>�tY>s��>�ԩ=0=hn�C&R?�����'�L<�7ί���B?�e?���>��N�ꔅ�W��??s�?b
�?k<w>�h�'c*�Ф?ԅ�>�`~���?מ5=��m�i��<������Qw��
����_�>G�ݽ�9�7lL���o��`?�x?�Y���Ⱦ��ɽ�����m=�C�?"�(?��)���Q�8�o�8�W��S�(���dh��w���$��p�p돿�^��9&����(��~*=��*?�?n��`��:��Hk��?�ۦf>�>�+�>
�>4I>��	��1� �]��?'�����"^�>"N{?�p�>*�N?[�U?b�R?�5?Ys>;�>�pɾX��>r��=���>�3
?��:?E�=?4�0?��>*�"?	;>�A����X о�)?(�?�p/?jH)?�?T��V㽜=Cg�;��S��Q���>�>��A�e9���=���C>Gq?g,
����I���>j�D?~?8>�>�(:�I�E�vE?��¥>���>U~7>����r�'T��+.?�?"-����<�P> ]�=��)�)A������=�T0>8?��^���ļ'k=�wJ�{�E����:R(��M%=� <D~�>g�?��>7�>`+���� �ě�m�=GY>�S>��>LFپy��� ����g�%#y>�t�?�v�?�mg=��=��=�X���1�����t�����<י?h?#?x`T?���?�=?�\#?��>� ��C���V��Q����?{'?�b�>�:��ξb1ƿE6A���>W:?�+k�}k"�m�7�&Fj�����t�>F��hp��⮿%�z�
��2��G�=��?kɛ?L�=����t�w������eۍ?��>���>e�/?���kX�Q����3v>��>��q?e�>>�i?�3�?'�r?_�W=p�@���.���({��p> �g?�ߖ?���?m�?X�?*��>򓶾5	�}̼�6��`h_�V����^|=��='�>��0?uK�>5��=�=����G_�i*=�+>�0�>���>�\�>���>�wf>��K?��>*[��������xo���;�Th?]<�?x(?�	=����58����7�>b�?¸�?Ǖ+?�c����=L,�/�ž�M�Q�>R�>{c�>�@�=���<�!>��>ju�>E��l5��!�P<��!?7?-�=�ʿ��y�Vﱾ������X<:��1�]�tȎ>ٰr�� P��̾�-d��W&�N�ξM-��Qۃ��<򾿡c��.���>��]=� >��=�n��`��9޽�e=��_>��'>��m=e~�=�Ԯ=���=܀
>{78>��=�>�z:�wӾ�q?�`2?	`?�H?�7c>c�>ru��g*�>xKf=�8?1�<>ڥ�=ԣ�L<d�S���*��	s�����}���U'ȾX�2>3��=��^>��!>�=0��=���=�_6=�g'�(���G:|�O*>�%=�"r=��>�D>F5�>�6w?X�������4Q��Z罤�:?�8�>l{�=��ƾp@?}�>>�2������zb��-?���?�T�?=�?Cti��d�>M���㎽�q�=N����=2>t��=v�2�S��>��J>���K��E����4�?��@��??�ዿТϿ3a/>q�0> 2>�RQ�o�0��V�b��"Y�U� ?�X:�pmȾ�ʅ>@�=a߾�}ž�=��6>�fa=!>��[���=q��,C=�;k=<k�>t�C>Ҹ=�����0�=C�G=���=7wN>�T�5q0�/m!��T;=���=��e>s�)>Q�>��?�0B?�Pu?m�>srD��l��2_��ȴo>���=R��>Ż{=<��>���>yw?�-? K3?᎟>��=�Ҳ>���>��B�Ӄz��jݾs���Q>\z�?�^?��>Z�=sY��Ѵ���:F2����>�m4?�?��>�������$�U�)��T���=��yk�;T�?��7 <y<��+.�tȽT��=�m�>���>5�>�GB>xg->9J>�T�>E�=�#8=87�=�=h�d�`<=���mӝ<����{ܼ�A<�eB-;��&=zrG������b���<yך��۪�s8�=��>m>�m�>O�=����wJ*>9����1L��z�=EA��Xy=���]�V6~�r/���+�d�;>�ED>��O����?ܔd>�.>��?W`u?��">���sž�替c�U�P�4��B�=�p�=�7�2�7�bM]�8�H��8Ǿ2�>UՖ>9q�>�]>v�/�q<��RJ=���=����>���,�@�'B�-�l�>�����\Wf�pZ��T3?�房�Q>鍀?�;?ב�?\��>�ܘ�6B�qO>�u���=�#�x7�����h�?�(?��>B�۾�h3�m�ܾD��ϳ�>��U��"L�
H���n-�{��<󭳾��>Y�����оM�;�����D���B��f}�j��>=4K?욬?�M���|��P�����$��M��>��e?Q�>�9?�	?��~��2۾�u�T��=��m?>u�?X�?��>j�u>��K�w��>���>�|�?.�?�>k?�ޒ�D%�>�a*>��G>�6a��i>1�>B�����=f?0?Dz(?fΟ�E
�����f��I��X�'��s���>*+O=x�r>`~�=����:��=�">���=���>���>a��>>��>㡲�6_�˳?>>�>�"?�_>ԢH�,>+	�=[����Ɂ��ߟ�)0?�#F��*��}�=��<����_��>H%����?�۹>�p9�Xy?N!従�ͽ���>,�=fw	��2�>�-�=���=[��>$�U>���=Ò�>�SO>�NӾNs>D���b!��&C��}R���Ѿϋz>�����&�������XI��t��g��j�k-���:=����<&D�?�}��t�k��)������?gW�>�6?t�����=�> ��>�Ǎ>#O������Z��[�Y�?���?�Ec>6�>`�W?ї?�1��3��pZ�E�u�W#A�Ee��`����������
����u�_?�x?yyA?
ʒ<�8z>���?��%��ӏ��)�>�/��#;��W<=(�>�'��l�`�%�Ӿ[�þ�<�#FF>��o?D$�?�U?�TV��Ɔ<�`U>��H?��??�n~?�|M?-�C?67!�Yr0?�Gk>�@?Ew?�?:\?�|?��>��	>Y�+�
>ݥ���/��ҼԽ옽���=]�=�p��?��L��J����>v\�;�Q�<R�<�}���=W>�<���=V�>��>@�[?��>0-�>��7?D|��G3�	����.?c�6=o�������AX�� ���-b�=�pi?_j�?�uZ?��m>�r>��+?��H>�+�>�->^H`>��>�콄�H���=8!>��>p��=�u\�������|������<�>�t�>N�>�
��%� >��l�}��[>�#Z��Eɾ�:�)QC�?�0�d�"��>��C?�4?��=Qb��^�˽S�g�|"*?��??0�C?���?��=��ؾ�9>��A�
����>���=M���p���������2��%<Q�y>j���:M���YX>�j*���վ3v���H����/�G>� %�K�ѽ�վ>��D�Ѿ�a<B<>�����"�+���S��1�D?�C4<`]���*���*�-L>�6�>�J�>�Ø�����C�tw��'�=��?_�l>GD��PR�g�j�&u��s>��W?wH?4w?E���1Z��n��4*�MX�A;)�A?�e�>��?O��>��=X���U<�es�g�N��2�>��?F�徾���cG'�z��Xo���t>
�>���=��$?Q�=?�4�>5Mp?��G?Ǟ?zU�>E���ٺ�ۑ ?�Æ?b>�ዽ�B#�'_(�CX$����>4�2?�����H>>"?��??;?8Il?�N?5�>���)6���>��>�+P��د�n{L>�C`?L�>GkX?/ӄ?oj�=��F��䏾�q�X�9<�u>%�7?��?�� ?I��>20
?��L�	��=X�=PYf?�р?8a?Iɡ<�*�>{rf>���>_��>��?��>3�==�s?���?P6?�s?-=#������X�(g���h��0ӽ��A�>0����Ce�����<� ���ɼ
7�����>	$=К�<ε[�+��>\m>������1>����|���A>�N��	���$���D��k�=��m>(Y ?L�>�m)����=�ϸ>s��>Gb�"o$?'??�?&(��8�a�e'۾g�9�<��>k�=?%�=yk��£o���=��n?�]?^�������b?7�]?d�K=��þ��b�#��5�O?R�
?��G��>�~?-�q?F��>9�e��9n�e���Bb�8�j�2Ҷ=ts�>�W���d��>�>��7?P�>9�b>��=�t۾��w��n��/?��?��?Q��?(*>��n�P3����l(��m�]?���>�@����"?�<���ϾW��;��4�ᾇ���mī�B%�������%�瘃��Aֽj�=T�?�)s?tkq?�_?BF ��d�D?^�����>V�q��h����E��D��C�u�n�������:u����E=mz��r@��G�?\�%?#�.����>�-����ﾏ˾�F>FW��N��:x�=�W����>=�T=�We�aQ-� T��H�?C"�>c��>�v;?~Z�f=��=1���6��E����6>?;�>���>�b�>ֽ:��)�u��6'ʾ+B��?b۽p$v>V�c?��K?��n?\��/1�����&�!��3/�W��{C>a>���>��W��G�,&�`%>���r�����y����	�\:=A�2?Mk�>
�>�e�?�?U	�u���Tx�Q1� d�<���>( i?���>d�>�5ν�� ���>l?��>$=�>���v- � �z�<Vν%j�>$߮>{R�>Rl>+b1�yb\��d��Ԅ��#8�NF�=�h?>+��d�`��3�>�&Q?@�:�a|<��>��|�h�!���+(�d�	>��?
��=e�;>�ž	���z�`���O�'?��4?ЄK��|!�;ظ>�3?�!2?�ֵ>�-�?��=Ǜ�X��~�?Z�f?_��?��5?6�>�|輠Kǽ58��A���|G>4�M>.;|>}��=H;.��5���r;��=���=�T�;T��QxQ��u=a��=�vP����=+ܿ1&P�n�Ҿ�3�����	��p����e����]�Ӻ�����pr�����E7��&r�!kt�����^mn���?f��?��������vR��N|��b�����>�Yn�����_���ʄ
�lƈ�Ȭܾ(}����!�7\M���f��%g��R'?_�����ǿfQ��D0۾��?�?�\x?("��'!�Dx7���">[�<�9�����񩚿��ο֙���]?KY�>�J�K>��~��>�>?�X>��p>�����A��<B�?�9,?`�>G�n��(ɿ�H��t�<���?��@�e@?�C&��j��q�=���>�	?�q<>a�8��x�i\��]��>�?{��?R�s=�iT�:�g�|t`?���<0?A�~�P�~��=L�=�Ƅ=���7rG> Ԑ>R^��;�f׽`�'>-!q>���[0���h��b<"�N>�jؽ�o�k҄?Rz\��f�e�/��R���Z>��T?� �>�p�=ů,?!3H��zϿ"�\��*a?�+�?ϡ�?��(?3㿾�֚>s�ܾj�M?]F6?R �>:k&���t�-B�=z=ἱR�����1"V�Q/�=e��>�k>�,�'��5iO�������=��/M̿N������ ��+��0���U�'���8������ԝ��3��9��a�¼�$�=cco=���=��l>ttK>7�T?�a?�L�>�W�<���u)�1����<�7��oa�~:����f���7���ƾa��t�-��L*�������q��X�l=� k�1�����C�S����M�(��?AA=��9���/�H>������V���<��=��^���������?�(7?:���V�&�:�K�=�_���[?����&�8�)"�~P�=���������3�>{e>lf�7��rĚ�R�4?s�?8��Iߧ���K>mŽ��z=p?��>W��<,��>��?�i�#�ΰ>`�>>�]�>�Z�>s0>N�����ϽR�?�J?z���+����>q����A���=@	�=��P���̽Y��={㿼����烛��P��á@=�wX?Hu�>�;$�Ӏ ��-��Qڼ%�7=� q?���>(�>	�f?��9?�Jt<e����|M��w���z=��S?�d?"�>��l�q�پ!����n3?�f?�9c>�r�����(�Bw ��?�rq?\?�ҁ��Qx�u���S��50?��v?�r^�Vs�����[�V��=�>6\�>���>��9��k�>�>?�#��G��躿��Y4�Þ?|�@l��?T�;<�����=�;?\�>«O�5?ƾ|��X�����q=d"�>⌧�Oev����R,�v�8?젃?1��>N��������>e?Y���?�h�?V����Z�"+��Nw�&��}N6=;�]>�o=n�=$Ƶ���>������K�k�8�ZNI�ٱE>��@ɜ�=C̬>�7==�ؿMwԿ6󉿻�(�A�6���<?�n�>u���pa�� S�"*`��.h���A��벾c�>n7#>AM׽�ꟾ��t��3�S��(��>�z��'��>jP6������ɵ�Uʨ����>h�>vtl>�ƽ��Ծ0�?}���c�ѿ�����辦)W?�D�?~��?F?�+&=#�,�?�x���@��N?5p?!�H?����,�{�ڼ'�j?����x�_���4���D���U>#3?y=�>di-���{=d�>�x�>O�>%9/��iĿǩ��y����Ԧ?o��?�*�Ѯ�>>|�?WH+?_�� ��aE��T*�TG�:�A?N�0>ާ��m^!�m�<������
?bQ0?_��&3�&�_?Ța���p�0�-���ƽ�ۡ>0�0��f\�^P������We����By����?^�?��?��� #��5%?m�>*���:Ǿm'�<��>�(�>n)N>�D_��u>C���:�:g	>j��?s~�?�i?ݕ�������V>
�}?�-�>���?�A�=��>
�=�����1��">\��= �;�ۜ?�zM?g�>�F�=��8�'M/��aF�bR�B�Q�C��Ň>��a?l�L?<b>�۸�ql1��� ��bͽ��1��켈 A�K�+�j߽��4>5>>�>�9E�]�Ҿj�?p�ٕؿ	i��x'��/4?��>��?���u�t����:_?�u�>�7��*���%���@�~��?�E�?5�?��׾Lx̼�>n�>�=�>hս�������7>�B?T�C��@�o�r�>P��?ض@{ծ? i��?���L��_^~�C��aJ8�L��=��7?�	���y>ƻ�>���=�Sv�6���s�s�|��>�9�?�r�?bm�>��l?g9o�?�B�թ0=k
�>_dk?z%?g�C����A>A�?�������+k�U�e?K�
@yc@{�^?S����ۿc����阾G9���I,;��G=Ə=>�a̼U>�E=:,�����=��f>rwh>HO>!"�>�Z3>&�o>��s>�5��ג*������]���/;����
ﾃ�����p�g����������>GX�r�ڽ�1�K����ŻA��= V?�R?U�o?�� ?jy�I>�����=i"$���=KO�>�`2?�L?�*?ou�=�뜾��d��<������z߇�0��>�%K>���>���><B�>ސ9��J>�?>��>��>�!=A���r=ߧM>��>y)�>p��>a�=>é>�)��|�����i��!{�b�Ͻqɣ?�T���[M�)���H񋾏ʽ���=ȣ.?>>�ԑ��XϿ����G?�A���V��%����=��0?�X?Ԭ>�G���=���>����`h�z�>V���g�j��*+�+?>H�?�g>(�m>�36�َ4���O�lӭ���w>>4?����=5��Ot�d�H�3�޾vyR>̠�>��$��b������|��"h�w+s=��:?��?�ǽ������z�>@����a>�yP><=��=ۑR>K�t��ν6A���D=���=�\>g?�W>'��<v�p>�T��{Ͻܲ�>)��=܄5>h�<? �>yi�9YJ���b��:��">�o�>�J>��L>�6�,��=/2�>�Z>)�ѽ�����.�~�н&��>�P��&��{��<��=�\���F�=�
�=[����6���ü�~?���-䈿��ee���lD?B+?1 �=0�F<��"�> ���H��:�?l�@m�?��	�ϢV�0�?�@�?�����=*}�>׫>�ξ0�L�˱?�ŽǢ�˔	�)#�jS�?��?F�/�\ʋ�5l�m6> _%?��Ӿ�d�>�h��[�������u��#=���>8-H?�]���5O�1�=�C{
?�?�M򾃢��S�ȿ}wv����>���?���?y�m��G��.�?����>���?qcY?|i>T۾AZ�,��>��@?R?�)�>6�y�'���?]߶?4��?OlI>~a�?�:r?�;�>Wwc�H/����������f=Ȭ;��>}>���+�C�Z���L���k�J��`\>�%='0�>o�ͽ����\��=ֈ��Λ��~�l�lF�>;�l>?�Q>@�>�r�>�J�>N�>�'*=y񝽲b������|�K?w��?����n�F�<��=�]��,?4w4?�h��/оF��>�\?�Ȁ?8[?�o�>��j3��jֿ��[��b��<��K>-R�>�A�>�ㇽ�K>�
վ5�C�Ӟ�>U�>>���@ھ� ��9c»��>�]!?y�>���=9� ?��#?��j>��>�ME�N,����E�z��>w��>.U?��~?�?r繾�V3�����ࡿ%}[�N>��x?�Q?ȕ>
���	~���uC��6H�����x��?Gg?�佚?,�?�??�A?3Ef>����ؾ���1ƀ>�� ?��ÔH��E�����;t?Y?�W�>�&��s��"���%��b��V�?��W?�?;n ��6Z�F����3�<Jټ�-<��;�wZ�s�>�D>��a��F>E6�=��=�[h���,���<3�=*�>v�>��?�Mi��?,?��F��҃����=۾r�JnD�T�> 4L>9��{�^?�{=���{�����w��$U����?$��?ce�?̴��h��=?�?�?7$�>QK���z޾O��{*w�_Lx��t���>��>�Wq��徦���;����B����Ž4�=���>��>���>B?`��>�ݬ>eػ��M��i�h�����A�Y{6�?�5��o9���4�9�P�9���g>�J���y���>‷�7c>�>��z>�F>V��>��ҽ�2�=�>掙>�<�>�>��4>RB,>��k��b��7R?�����	(����g��N&B?N>d?W��>R�i��W�����UF?�b�?�m�?�Tv>��h��,+�RV?��>����4
?�:=!��ք<�3��p~�2S��~=��7�>i+ؽ�%:���L��f�xU
?->?X����̾eֽ�����>|=8��?G�'?'	*��5P��o��KX��T�I�� Sl����[$�q�o�Չ������HB��)�*���=ˮ(?��?#>�]0��?g���)h��|=�O f>�#�>L��>�~�>��V>��
�v#0�.\��c'�pJx�a*�>��z?���>`�`?�/P?��a?��O?ګ�>�"{>Ǽ��5 ?HϽ(-~>�?�'?��%?(�5?��?;*>?!�J>�o����	���?�]9?�?"?��,?Wo3?tk�1A���#=�z�<Ω�"� �f�޽���Ě���{��GR>"�f>�!?���ܢ�����m�>��M?~��>�ف>ꧾ��E�Sm��T�>�' ?e�4>�I�
cw�����M��>�z?O�����=��>N/�=T�<���<^P>oT�{=B=�"+:ǅ��������=���=�����̘=�`Ӽ�ü9 =�O?Dg?�>wUh>{ux� m��3��_N�=�Ln>%jm>��>q��o ��vk��l)b�+ o>�M�?$h�?]_�=�i >�~�=����m�ƾ0�����_;�:��?��?W�V?�v�?�j1?� ?c��=���w���2M��!���9	?Y( ?�i>���d��
Ϳ#�5����>4y	?nYi�@���L�7��[W����o>�:ʾr�,��l��a���о�qr����?-�?-��<����%���u�ҿ�N��F�?�/|�'�O>�E?xt|�aC���=���>��u?�,�>_8�?�jf?/C?��U>U5Y��Ŀ	T����ZO>�݃?��z?�ۑ?�5�?.&�>�`�>��o�0}�"�
�U�k�bV����a���>��e>��>=�>��>�+z>�K˽��}�&�{��`��=b���>d!�>pf%?�X�>�C>��H?��>�Բ�OB�����I}���8��q?R[�?��-?Ǿ
=h���F��s����>o��?m�?P�&?�lG�B#�=�����y����z��>8Ļ>_��>ꍍ=�3�<M~(>�Q�>�@�>~���O���2�p��+
?�%B?TY�=���/��٪!�����~����M��W��g>��W�>�ʽ�T����̽��m���оK�ξ^��~l���+�>�P��B?�n�=��a�ԉd>5�`�/]�eO= N{>�F>�Gn����=� �=���!�!�]<!;�=]�6=���=B
>E˾l�}?:.I?�l+?��C?N�y>%[>�D4�2b�>�f��;1?��U>�MP�Z����`;�������٘ؾ�c׾�c�Ƹ����>��H���>0@3>:�=�%�<@v�=��s=Ŏ=�R��=���=�/�=���=9��=��>�s>=/w?V���߸���.Q��D车�:?"�>:��=��ƾT�??7?>*�������q�Y,?���?B�?��?Z$j�j�>���z[�����=����Hh2>��=�!3�܋�>6K> ���U���K���:�?x�@��??�苿�Ͽ�`/>�G>=�>�L�	)4���N��T���O��L?-<�� ���c�>n��=r�޾{�ƾ0�='S1>W�=����"U�/��=��k��=�g=M��>�E>n��=w������=�v=!D�=FM>9h��]y�+,2�XI=O�=�6]>ki$>C��>�E?�<?ac?"��> �{�lb��7�����>�:=��>��z�*~P>�A?~�C?�k+?��B?���>9<�=ּ�>h�>��)�_g�i�󾋒��ރ�=���?���?"�>.K�J��.&��7)�,{^=�4?0F ?ى�>I��>w?�Y�-&������Go��V�	<�R%�a����<���
�I�hw=T�q>A��>���>M>�mn>�R[>�>h��=L�:<H=xE;=)���}l׼*�=.�����7=Qb��������];p}��fܭ�@4��g�Q�g�F�w_B�]��=���>;>AM�>��=i����/>������L���=����FB�Dd�?~�D�.���6�(�B>��W>�͂�=񑿔�?qtX>R�>> J�?�'u?�7 >��@־���wd��R���=��>�<�!�;��J`��M�2pҾ���>֎>���>8m>��+���>��Nu=�m�E5���>Xk���a��	�&�p������i�Ty���\D?�+�����=;~?XI?��?�P�>p@����ؾ�/>�����=���p�Ԏ��W�?\�&?�a�>P�뾭�D���߾���Ҙ�>�Q�|tQ��×��T ��>�)��s�o>!㐾eר�+�2������І�	T�tq��|�>�yH?�Ϣ?��r��&t���G��G
��ǐ��%�>�"[?�Am>=�>�m�>�����Ӿ�K���=qn?Fq�?0��?��<;1-y>*�ۼxQ?  	???G �?gр?K�B�p ?2>�>���=C�c�@>Q�.>�1��=}?s��>��'?*&6�h�� ���
�r,��G�/=�^�<ع>�VZ>"E#>$��=x=8�;>3}>���>P��>�.y>}pG>Կ�>^���d�R	?��>�(�>�_.?z�o>e� =x����[=l/I��(S�דH��G�Q���1�:�_����=糂�MJ�>�K���X�? �t>!n�\?f��� ���-�>8f#>�����r�>AU>�k>�p�>�Ӭ>�k)>fe�>��(>����N�>�^#�����)���.�QžX��=�q��+ç�{ʾ$=ς����r��ܷ��n��u���)��b���?�S�e������h!�=<�?w�>��4?�5��� =���>&��>`�N>����X��֫�����
�?"v�?��h>�"�>��Y?�?��-�L�.�oW���t��=� b��xa�=������k�
��ǽ4^?��x?�V@?�3�<D>y>1�?cu#��I��B��>�d/��;���i=sZ�>�����eW���׾�8þ����^L>w4n?���?��?��_���T��#*>�m:?��/?�:t?L2?��;?����$?`8<>��?V�	?��4? �-?s1
?B�1>	��=���c�0=�4��4�����׽��Ͻ����75=F^�=^:(�w<�k.=<3�<���j�ļ>9�;px���u�<A/4=�u�=���=�x�>�R?I��>QQ>aN7?V�罳� ��	���� ?���=6��Ĭ����־�_�j,J=(zR?u��?�
E?�D�>>�*�&06���>Ixz>)v=>��R>�R�>Ї۽�2�KJ>��>d1�=��E=(����b�����$ ��/P=�S>o��>Uk->'�?�"��>��پ��=��T�= b������;+���C��B����`��>��0?���>)
ʺ�w�#,�X�S�X�7?��H?��4?r�?o��<h�E��-�/l轠��>Cݞ>�1��2��t��b�?��,!<���>mo���U���WZ>����v��>Zt� �J�g���=�L�׎+�J!�#�ԾӜ��UCc=���=Y������1��=w��"mJ?*k=锠���)��þ��>�2�>��>�9�7Fm�>�������=��>��J>�4�yF���O�����!Y>��R?�#n?��{?�䐾�wp�Uth����O���C:��43?u�>�O?��>�=��+q���?�s�h��N;����>��?����.�8�|������v%F�-��>��?��?=q5?D(??��>Y�p?�96?�)?��1>w��/��>&?ۉ�?C.�=�Խ�T�]�8�!F�i��>�)?&�B��×>��?��?r�&?�Q?�?|�>� ��<@�$��>U�>��W��a��V�_>f�J?���>;DY?у?@�=>'�5�����=��>��2?:#?и?��>�.?�R.�����d�=R[?��p?�s?��L��>hľ>:�>Q��=5�>�>��>'Q*?���?��_?�7?��>^�v�����=�W�=M�=�瀽!E><�t�=R�żB�0=��=ޝ̽Ò�G��<�Pu��ͧ�K
��X�>f�s>�����0>��ľbK����@>tӣ��P��ъ���:�&�=̌�>��?试>&[#�p��=ߥ�>5?�>����5(?.�?%?�~';
�b���ھʭK���>=B?��=�l�(���Q�u���g=��m?ي^?%�W�����b?��]?g�=��þǳb���l�O?��
?��G��>>�~??�q?ȷ�>��e��9n����kCb���j�lѶ=Or�>LX���d�;?�>=�7?�N�>��b>(�=:t۾%�w�Nr��@?|�?k�?c��?L)*>��n�	4�\�����*�V?#�>�����#?4L�Wx̾���� x��&������;&��>���qŤ��?�d���_������=��	?�)m?��l?��S?R�����f���Y�T>v�bMS�a��E��vR?��@�3�A��-i����&Q���H��n3!=Ӌ��� d����? gL?l����?1u����2�����=��:QB�Rm2=��ݽ� ���y�|�����нJ�~�0]?s�>��>*�3?)�:�I�<�b"��V7�e����>�I�>�`�>G�>���QY%�
���gپ�姾Է��v>nwc?��K?��n?	�q1��v����!���1�����KC>WH>\,�>��V����6&��U>���r����\����	��~=��2?�1�>�>�Q�?��?-d	�k*��ǉx��r1�r��<�
�>Yi?N�>���>�н�� ����>B�l?,��>���>�{���I!���{�=ʽ]2�>h�>h��>��o>¨,�\��k���x���8�L<�=�h?�u��8�`��ׅ>KR?D��:�kM<֚�>�ku��!����z+(��>�?�T�=e�;>mkž�$��{�z-���$?S1?�X�����Џ>@�!?�{?�6�>���?�r�>��Ǿ�4!;��?59U?��w?�c?�D�>��]=9g�n���D���lK��l>#uB>y�����<����X�y�����K�0>4�3>%���Oo%<Ļ7\�����=�f�=[$�>Ή�[�!׾[��	�־Α������d,���Vyl�"L������籾���}���5�@�9li�]~t�B'e�c�?�v�?>T��F���eV��Q�g�뾹v�>�L�8����b�<��˾p	���Ӿ����|<��h]�ڌk�R�'?�����ǿ��:ܾ2! ?�A ?/�y?��.�"���8�� >�C�<-����뾬����ο9�����^?���>��/��Z��>᥂>*�X>�Hq>����螾�1�<��?>�-?��>֎r�-�ɿ[���ä<���?-�@��A?��(�K��KT=>��>��	?/�?>�E1�2��̰��J�>�=�?���?M=ǷW�[��e?��<c�F�\(׻���=rģ=��=,��J>�K�>����=A�ϝܽr�4>}�>g������^��g�<��]>�ս����5Մ?,{\��f���/��T��U>��T?�*�>R:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=~6�$���{���&V�|��=[��>d�>Â,������O��I��U��=��.Aȿ�>#��a�ݸ&=G��W��� w�����}��yt����i�����c�<þ�=o1N>�}>�jW>�U>[�R?�yn?)<�>��=O��垾�̾f�=�Y��l/�������,��U����#���"�����>ξ��Y���w�H!d��=���%������1D�R�r?�E���5�T�\�7��FE�;�F�nR>��C�=��h�:?�\���i�?��H?����)f�5�G��Ɔ=G�ν��Z?ه�,��ș��5=B��=ב<�#x>h��>�E��&�I��_����/?_�?ݸ����?4>�����h=�
'?�?���<�P�>uG'?}���i?t>�7>�z�>"�>�r>3�� ��j?��P?!�뽐���,ʇ>�Fƾe��`(5=�I>ͧ �@$��;^>�5�ۿ�� WF��*P���=NGl?T5�>G>;�d���:$�U!�=���=$h[?M� ?Y�>v�\?�D?���<F]׾�4;�2_���	>�:d?|Ss?��0>�1!�����͸��%?�c?�t/>������� %�e'�=�!?��?�?A�����p�ѧ���v ���.?.�v?�r^��s�������V��=�>�[�>���>��9��k�>��>?
#�NG��޺��wY4�Þ?��@r��?O�;<H����=c;?\�>��O��>ƾ5z��<����q=:"�>茧�4ev�r��9R,�%�8?۠�?�>�������u=������?��?g7��v�=8����q�F�u�=6�K=~�v��R�T.ھ�#X���ݾl��� ���xo�Oċ>��@��=��>|&���	ٿ5~��<���;?��>0��<j�ɽ�hQ��P3��P���e����H�>p�>e��(	��M�{��d;��`��w�>Ç���>��S�$������'3<��>`��>���>�0����!��?oC���5ο�����~�X?�d�?�f�?�n?!�9<L�v��"{�����G?2ts?K Z?'>%��]�j7�/�j?�_���U`��4�kHE��U>�"3?�B�>P�-�a�|=�>���>[g>�#/�u�Ŀ�ٶ����Z��?��?�o���>j��?js+?�i�8���[����*���+��<A?�2>���9�!�@0=�XҒ�ż
?X~0?{�`.�[�_?$�a�H�p���-�q�ƽ�ۡ>��0��e\�5M�����Xe����@y����?O^�?e�?ӵ�� #�d6%?�>_����8Ǿ��<���>�(�>�)N>�H_���u>����:��h	>���?�~�?Uj?���������U>�}?�#�>_�?t�=�a�>�h�=�<�,��e#>�"�=��>�?�??�M?N�>I_�=��8��/�@ZF�3FR�#��C�$�>��a?_�L?�Mb>����2��!��pͽra1��K��X@�x�,���߽�%5>0�=> >��D��ӾN�I?![�yt����܄����I?��>��>��澧�@��o�<��{?���>���PШ�ޛ��]_>=���?��?�D?Oɾck�d�G=�XP>/�>��x�.4�<(����=,�,?5w<�+�K��b���*>O�?mi�?��?۬J��	?���P��Va~����7�f��=��7?�0��z>���>��=�nv�ݻ��X�s����>�B�?�{�?��>!�l?��o�P�B�x�1=6M�>͜k?�s?�Po���f�B>��?!������L��f?�
@u@`�^?)'p����������rP�"��>6r�=�G
>����nV��/��ͽ�B|=.��=���>8��>
��={2P>��p>�j>mT�ߍ��B��Q���~)��08�P�&�}m����0�����A��~���(
�ԗa����:g�����R�ʳ����= \S?�Q?�=q?��>�~6��>���#^�<��	��]�=���>(�9?U�K?O�/?p�W=p)���9b�F�}�&S��b��cg�>�5>��>9��>�Z�>�@�;Yec>�/O>��l>���=��<L	��`E=��Y>۫>���>�P�>�>���=�g���²��y��A���&K�ES�?�YӾ��}�Y���І��p�վ���,?�6�>�����տ1����/@?B��˾���=�<t;sA�>��>?���=^�R����=�&=z�Ⱦ5��|G�>H�=^���W"L�⦺� ��>?g->�->rN2��}'�l���ܾ�� >��3?����6F���q��]�B�;��>2�>��n�.�>���"���p��{D�=b�K?�f�>ͩJ=��Z�[ ���پ�U>���>6-�=��>�S>@��^�½:K6��:�=}FQ>v2�>S(?;A>
�=��>̶~�+�1�勇>[�J>ߣY>��<?�>?R���[��������`�'!Q>���>	Ù>�a>�&9�C�u=�/�>��K>S����3��z�W��ty>'8��Q����޼$!
>����-�>���=O;���6�]�K=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�@�>!�����o����t�a0=��> �G?�x����J� �<�U?bi?���a����ȿweu����>���?Ɣ?|km��h��$@�Q�>�S�?�Y?؁k>D۾./[��%�>��@?�R?��>^�RH&�7'?�i�?~�?�'G>�?(t?���>���1�/����^���O�m=D;ɫ�>?�>����&D�d֓��M���Vl�R]��~^>��(=��>4�߽�����ѱ=ˣ��p��&~[��X�>d�k>.�R>R�>� ?��>���>��7=t�����}�������K?��?��� 0n�Q{�<���=��^�,&?�L4?��Z�`�Ͼ�Ө>��\?���?Y	[?S^�>���;<��k忿{��͝�<��K>�0�>@F�>UA��'=K>��Ծ�9D�~n�>�՗>����8=ھf'�������=�>�e!?��>�=֙ ?��#?��j>�(�>aE��9��"�E����>��>�H?�~?��?�Թ�wZ3�����桿^�[��;N>��x?V?Fʕ>P�������TjE�W@I����c��?�tg?PT��?32�?�??,�A?	)f>���ؾ������>L�!?8�2A�� &�0����?��?��>1���ѽ|�伊���d����?��\?a�%?�\���`�˫¾d��<���7N��: <�1I�N(>��>Ǩ��?<�=~>�ΰ=�m�[�5��+�<h1�=�Ǒ>�G�=%8�#8��0=,?��G�{ۃ���=��r�>xD���>�IL>����^?hl=��{�����x��!	U�� �? ��?Zk�?^��?�h��$=?�?R	?l"�>�J���}޾3�྽Pw�~x��w�\�>���>9�l���J���ڙ���F��_�Žƻ?��O�>ȶ>��>���>F�H>���>%�����yԾs� �R�V���E�1�E�-�t�&���<�=�zD}�;Bľ6�u�˞>/�N�Gp�>b?��{>��Z>���>�]Ժ1�|>x�.>�]>��>�$4>R�&>�>'�g=�	ǼLR?5�����'����p����3B?rd?�0�>Ui�S���|��I�?V��?�r�?I@v>�~h��++��n?�>�>���p
?9C:=J=��8�<�T��ȼ��2��@�f��>bG׽ :�\M�%lf�k
?�.?���p�̾�:׽&����o=2K�?��(?�)���Q�ýo�l�W�S��t��6h�cp����$��p��ꏿ�]���%����(���)=�*?.�?~�t�����Vk��?��>f>���>#�>:�>U�I>��	�t�1���]��='�˾��gT�>2T{?�=>eQ?cqC?ƲK?�c??��j>��>ྫ��>6`�=��>��?8X;?�5?P1?W��>%'?��W>@�|���q.�e�?� ?3�?O?�l#?)b��ͨD�aw�=a҂���)�x +=3�(=N�;h�/��@����=��>>�?�(���5�����p>�6?e��>��>�;����w�:�<ԧ�>�?=Ս>�w���r��&	�H��>�(�?���9=�f,>0��=4�t�W�����=6����Ư=L�>��]��B0<V��=N�=�����C<�h:���!�<�]�>�?�Պ>��><���� �Q���.�=3WY>s�S>i�>@پ^s����_�g�1Wy>�s�?�u�?~fg=�!�=i��=�e��Z[��Y�����>��<��?,#?@�S?�g�?��=?f#?b>�6��0���F���v��ۢ?��?9�.>���.���;/��xsY�?�> C?C�K�v�M��8�%�&�o��>�����r�P㫿p�������a*����?�v�?N==#�����4������
m?�}�>ER�>��>�����M���!��b>9"?��\?@�~>��m?�Q�?��d?:>�7+�T5��%����נ�|�>��?�υ?�֌?��?��>�L�>f�¾+C����ľX���@�ս���g��=^��>�f�>]u?��t><q�=�O�=,h`�̞�����=|S�=%�?9� >:�?d
^>:�=`AD?�	�>�����{�Xd��_탾�^����q?R��?~-?��x=ښ��F�u��o��>���?zת?R&,?R�G���=���,6�����ϲ>hl�>�͢>'	�=��5=^�=�V�>q[�>�k�r�e&>��'9�y�?�M?mp�=�Ŀo^o��p�X����*�<�����SX��>��ІK�� �=����$�쩾��U�Ď�����䕳�Ki����x����><�Q=�$>_��==� =����=b�<~�3=W��<���<'L����n���j�#<�m��X
����<���=VU�;�\˾�t}?",I?�~+?�C?�y>�x>� 4�?Ȗ>
΁��&?$V>��Q��}��:�;�����x蔾�}ؾ�7׾��c�����c>��I��>�F3>9�=�݉<jE�=v�r=���=8�O�Զ=���=��=o�=���=h�>ٙ>�6w?V�������4Q��Z罞�:?�8�>�{�=��ƾd@?q�>>�2������b��-?���?�T�?5�?_ti��d�>K��㎽�q�=i����=2>s��=v�2�S��>��J>���K��*����4�?��@��??�ዿѢϿ+a/>���=�>VA�{6�]�}���4�n�g�
?'�$��5����X>d�=Efþx�޾A�㼩�>�Ƽоk���W��5�Γ;��4F=5��=2Y�>���> �S>����ȸT>Q�b=4��=y�)>����~\<!��>>��N>P�v>��> ��>�=%?ˀ=?�<Q?���>�#g�,��`ƾ���>mQ�>��>&�<RB>�>~3?�3?��D?���>���=ӭ>�#�>j���䀿gξ��Ⱦ�}�=s�?gmw?�"�>���<�R��=(F�E�X����?�Q?1�,?J	�>�U����5Y&���.�݈��S�3�+=�mr�4QU�����Tm�z�㽇�=�p�>n��>��>-Ty>��9>��N>p�>x�>�7�<�p�=�ی����<]��a��=���� �<�wż7ʉ�4&�:�+�M����ލ;]��;��]<%��;��=}��>�1>���>�h�=����K/>R����L��ؿ==D��'B��*d��D~�{/��:6�F�B>�X>4����0����?��Y>�g?>څ�?'@u?� >�$���վ8J���@e��IS�˷�=�>i=�Jp;�@M`���M�fZҾ�>�/�>�f�>Ml>V�,�K-?��^r=ƣ�[�5�m��>���h�'�`����p�bि/ٟ�2'i��@��xC?v.�����=O~?C�H?�
�?i�>/�����پ�N/>�逾h�=���v�o����/�? S'?PB�>����C�T̾)1���ط>�JI�k�O�+Õ���0�����з�A��>�����о�'3�Pi�������B�)Or�D�>]�O?��?Eb��U��;YO����+/���q?p~g?J!�>;F?�@?���U~�G����Q�=��n?/��?�9�?��
>#>���φ�>���>Ql�?z?�?H5u?��ؽV��>(�=�Y�=`Z���=���=���=�^�=��	?�?|?ty3�g������Ծ�7�1�=�y
>X3�>t�>��e>����'+[=Ղ.>D�b>c��>L�l>��>�fB>`i>(J㾥$+���?��>W�9>��1?rW�>Y�p��fV>���nA��W�R���IK���I��fh�Fm����=?һ�~�>n8�����?2Z�>en<�
�&?8Ͼ������>��½�L潥^�>���=�� >�N�>��=YH�=kc�>���>�Ӿ�e>˧��!�u�C�ԀR���Ѿ��y>Zd���%�J�������H�9f���� j��0���p=��V�<ҿ�?CW���|j��5*��y��4B	?I�>��4?Sˌ��H��[>>���>��>M����9��J$�����B,�?���?�;c>U�>Y�W?ך?�1�c3��uZ�ήu��'A�}e���`�s፿���ȗ
������_?�x?+yA?ET�<:z>��?��%��ӏ��)�>�/��&;�J<=9+�>�*��2�`�S�Ӿ��þ�8�<FF>\�o?1%�?�Y?DSV����<,1`>bY-?ɔ?�k?`N!?�DC?��1?Iن>r?��?��+?�T2?�)?T��;�@4>/U�=��=�C��������(� n���<E\�;Υf�oO�PŽ�F�<���=��]�{%�듳<�f���"��a=f�>	0>|�>!._?�}�>F%p>?�4?&����)��Ú���-?M�==W�����R���/��z�=��c?��?��]?�5i>�k3�ţQ�	J>��w>0t >n�t>��>aw8�c@�Fe�;T�=��(>���=-%���u��z��d��aj�=ě%>G[�>
�{>^l��Oe'>8H����z���c>X�Q�-��.JS�t�G� 2���u����>��K?�z?8��=|�龫F��%;f��,)?x~<?��L?�
�?0�=��ھ:�t�J����k�>ȿ<T��������&-:���:�6u>f1��5����$b>=����޾ݩn�J�����oP=�o�M$R=S$�p�վuv�S�=�"
>�v��i� �d��|ܪ�0J?29j=�n��n�T�*���s�>�ۘ>a®>��;��x��[@��۬�	ו=��>��;>�q���Oﾍ�G��2�<X�>�P?=�j?�?���j��+?�w��I�Ծ��<��"?�/�>��?�7g>��[<}B��y.'�j�[���4����>�&?����L�EV���ھ9'�b�>�7?o�>r�?]�\?�?J^E?~�!?E�?�>���譶�1�%?��?ے�=%xսIT�Կ8���E���>j)?�oA��f�>:�?ǣ?��&?}}Q?�{?��>
	��2@��Ô>ֲ�>��W��Y���tc>6J?���>SQY?�փ?�>>4���/����=��>�53?.R#?o?%~�>͜?��K�^{�=���>�v?~�?���?5�6=T��>D��>�^>��,>�(�>pp�>bt?��*?cɃ?]c?��$?�X=:�����΍K��t�<d�@=�(==`f�=-K7<�����t�bM"=�Y�l����	=n�D=M����v�8=2��>�Ht>u}��Í0>�ž ����?>���te��Y���~z<�6��=��>��?��>!&�=��=���>,5�>	���(?�?�Y?y8<%�a��پ�I�/�>�B?��=U�i�C���:v���n=�o?zu^?3�W�+m��O�b?��]?>h��=��þz�b����f�O?<�
?2�G���>��~?f�q?U��>�e�*:n�*��Db���j�$Ѷ=]r�>LX�S�d��?�>o�7?�N�>0�b>-%�=hu۾�w��q��h?��?�?���?+*>��n�Y4�6J�)����MT?�F�>������9?qq=E�Ҿ��)�Ч����Ǿp�Ⱦ�.��fx��ڦ��$��Z��_J�J>��?�i?x�x?ռk?����j�x�S��q�ak�t�����r2��]4�M2F��}��Z�i6�����J��=�5|�sGF�v��?�.)?Yp4�-z�>�p��]Y��̺�r�<>����%+��=i���%=v�E=8�Z���aA��\�?�O�>�s�>dA?OW��@��8/���4������(>��>��>ʕ�>�m��kyN���ý��Ͼ���o����.v>	yc?J�K?4�n?�j��'1�`���I�!�Y�/�M[����B>7>���>o�W�8���6&�Y>��r�:���z��i�	�Ȉ~=��2?�?�>/��>aP�?�?�q	�#a���Cx��x1�}'�<�%�>i?�P�>8�>н�� ����>��l?���>��>󖌾qZ!���{��ʽ;&�>�>��>��o>5�,��#\��j��R����9��u�=)�h?���J�`�U�>�R?��: �G<�|�>�v��!������'�E�>c|?���=e�;>#�ž�$���{��7����)?�?|ˑ���)�[�>��"?,�>�`�>�̓?�%�>4�ľR�N;��?T	^?�4J?��@?^��>��2=z���`ƽ�I'�o1=���>��Z>��s=�6�=���Y�����VD=G�=PA�ڀ��)~#<*p����S<T�
=�Y5>�]ۿ��K���ھHT���ZE��ꉾnC���e��^k�������������&V�f0�'W�խ[�E����(g�=��?���?�)�������f�����f|���n�>oc�xW��6������0��>a�R%��<� �6FK�b�e�o�f�P�'?�����ǿ򰡿�:ܾ4! ?�A ?8�y?��7�"���8�� >FC�<�,����뾭����οC�����^?���>��/��q��>ޥ�>�X>�Hq>����螾�1�<��?6�-?��>��r�1�ɿc���v¤<���?0�@�|A?"�(����V=���>��	?v�?>�U1��I�[����R�>�;�?���?�{M=O�W���	��~e?kF<��F�޻
"�=	=�=2=,���J>NV�>��'PA��9ܽ3�4>ޅ>"�ܮ��^�^��<�]>_�ս�2��5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=u6�򉤻{���&V�}��=[��>c�>,������O��I��U��=4� ��
��a
"�Ae*��ұ=�`�������� Q�P)Ƚ���k#��p�³N����=�T8>�S�>��>�{>VV?��g?���>~�=�bJ�~��l�Ⱦ>��=>R�,�.���Ǿ���=Ey�g�
c��z5��CӾ�ྫ��Q�*�-��p��ܞ��q�$lJ�e�[�O�f?��>3��� l��K<�s��8U1�ʘ��o�S= �o<ó⾏�n�;ۜ?ӧ$?�:��1�6��p:�hd�=�����X?�Y�Mq5�nൾ��<��ͼ��B�/��>�UN>�C�k�9����\0?_?�X���t����*>�N ��q=��+?w?vg<��>ja%?�+�\%���[>�I3>�ޣ>΅�>��	>���ܽ�j?XiT?|.�Nx��I�>e:��pz�d=b= >h�5����t\>��<D2����V�0�����<�4W?Gȍ>y�)����������iB=.vx?�W?"r�>I[k?C�B?'�<�`��Z�S�`�oy=�W?ECi?��><����Ͼ`R����5?z�e?u�N>-h� ��:�.��!���?/�n?V??彙��m}�+��2���_6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?q�;<��U��=�;?l\�> �O��>ƾ�z������2�q=�"�>���ev����R,�f�8?ݠ�?���>��������=-s��'ۭ?���?v��<]%;>|�B�p���&�l{S=$�>������N�����[�R�n�������犾�5�=�Ë>�@Ͽ >�e�>E�޽C��\�Կ�+��A~��G�6?''�>�^�<��|�)\Z�ەA�;Y���L��貾�G�>�>s�������{��i;��J����>�%���>��S����L�����1<!ג>u��>���>p���; ��q��?�H��^7οP���u����X?�c�?@l�?ph?h7<�v��N{����U"G?-�s?�Z?��%��}]���7�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�?���Z��?��?�o���>r��?ts+?�i�8���[����*�l�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.�]�_?&�a�V�p���-��ƽyۡ> �0��e\��M��w���Xe��� Ay����?J^�?a�?��� #�N6%?�>c����8Ǿ�	�<���>�(�>:*N>yI_���u>����:��h	>���?�~�?Tj?���������U>�}?��>��?�l�=Y�>Fg�=�ﰾ��,��`#>��=G�>���?�M?UJ�>�H�=R�8��/�0ZF��JR��$�E�C���>��a?yL?qb>��/�1�� !��Fͽ�U1�~p輗2@���,�:�߽-5>�>>~(>��D�y�Ҿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��[a~����7����=��7?�0���z>���>��=�nv�߻��_�s����>�B�?�{�?��>&�l?��o�[�B���1=M�>ʜk?�s?CFo�p�G�B>q�?!������L��f?�
@zu@K�^?1J�ȿڧ���μ�����u>�=%#>���yY�r�e=�y�=��.=�޻;p#>���>�N�>�G�=�<>�^>��{�����E���?��U �x��g!*�0x��|�¾��վ�:��ab	��'.�A���Rr�����S�k�l���y=	DZ?8?�@?:��>(�����O>$��\�T=����t�=�	�>� ?��,?,�1?���=`$��N�s�L�r�|����Kb�3\�>F��=��
?�9�>���>�3�=շ�>:H\>�
�>��F>��"���<�?h=�,�>���>Z��>~�>�ˁ>l��=�㸿 ����{�����
S�"@�?p�����<z�����h���Y����5?+C)>�����hҿ�����@?N$�������1�=3T�<���>׈a?�T�<����?���JE>�4��~m�����>�^�=�;�vF�V�1=ܦ?��i>�q>|4��N7�� R��O����x>�B6?;��� h?�Ҝu��TJ���޾#�O>5t�>�����g��S��p���/i�f}=zD;?bF?���������m�����FN>vd>�o=�ۥ=��O> K�B�ǽ�%M�F
)=���=��`>TS?P�+>и�=ΰ>Y&��T]O��ȩ>,6B>�Q,>L@?z%?:F��I��j����-�v�v>5X�>�)�>F�>�'J�!^�=(\�>`b>���Q삽�{��?��7W>�}�c=_�`v��fy=d@����=�ԓ=�� ���<�={'=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��ӾPh�>{x��Z�������u�x�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?soi>�g۾<`Z����>һ@?�R?�>�9��'���?�޶?֯�?�dM>v��?.8z?86�>>�{�|�0���Xʍ��r<�e�;��>��>
7����;��Փ��(��ko��l�
�b>��J=��>�f����O�=`���<뺾�L�q��>�Y>�~@>�N�>�?<�>$�>eS=b��G�v��ӡ���K?Z��?b��'n��x�<�z�=\�^��?J24?��Y�1�Ͼ��>��\?T��?l[?V�>���@���࿿����?��<��K>g��>}��>�.����K>��Ծ�C��z�>8�>3���~Eھ�;������M�>�k!?h��>1��=ՙ ?��#?��j>�(�><aE��9��T�E����>���>�H?�~?��?�Թ�{Z3�����桿��[�4;N>��x?V?�ʕ>Y�������fE�BI�X���X��?�tg?LS�2?A2�?�??L�A?�)f>l��ؾj�����>��!?����A�xL&�?��N~?�R?$��>+!���ս�5ּ����}��U�?7(\?I>&?����)a���¾�/�<Da#� bU����;D�
�>;�>J���ߐ�=�>ܰ=�Um��E6�Dg<`b�=�z�>"�=�7�W��0=,?¿G�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?b��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>%�l���K���ڙ���F��_�Žٲ�ܞ�>?��>s`?E�>��M>�ܰ>\���'�:�V�ŝ]����<7�`-�2=������)��g�
mþ�As��f�>\����>�K
?Ck>q)|>��>�@����>q`>�t}>���>H�Y>'A>59>LK<�5��IR?'�����'�7��}��� /B?�ld?H&�>wei�C�������z?2��? q�?�?v>p�h� /+�$f?�0�>d���t
?��:=����Ԋ<�M��E���5�����!��>�׽�:��M��f��i
?�6?C���f�̾�	׽f���Eo=�L�?�(?��)���Q�t�o���W�8S�D��&9h��i����$���p�돿�^��N%���(�$O*=��*?��?��������#k��?��bf>��>q&�>��>s�I>��	���1�l�]�VE'����bN�>[{?�\�>IG?�<7? �H?�K?E��>�>I����o�>5=�<@��>��>�84?��,?uY0?s�?k�(?�aL>B����}��(��l?��?��?�a?�?�`��[���xC���ۼKM��ޖ��>��= �<_��EI�f��=u6a>�q*?��o������ �>�{X?��?�C�>���&n��osһ���>���>�R<>>����Yt�>o�/q?H��?t�?�8-6<"#>�|>uS�=��.=b�=�f_���=j�<���?��;@�O>M��=ˌ�<���#��<?,�u�6=u�>6�?���>�C�>�@��)� �]���e�=�Y>FS>~>�Eپ�}���$��r�g��]y>�w�?�z�?�f=��=��=}���U�����?�����<�?<J#?'XT?_��?x�=?`j#?ϵ>+�jM���^�������?B1?�Y>)��SǇ��۷��@����>��>�W��c���A:���=��L��>|��i_���!���uf�켏�q���p�?�?U�?j�=$��Ke��e����Ծn�r?�>���>L�?���s�S����	F>�>+{O?%��>�fx?P�?�Qo??]W=r�4�'L��k6���5�=t�t>�Z?K�w?8q�?��?9��=-��>R�y��l̾�8��sl������(��v$>%��>8��>��>�:^>]�+>�F��ky�������6>h�?��>�I�>kѺ>Z�,=��G?���>�]��$��$줾=Ń�!=��u?囐?ȑ+?T=6���E�mG���J�>]o�?���?4*?*�S�3��=��ּ?ⶾ��q��%�>�ڹ>�1�>�Ǔ=�xF=3b>��>���>Z)�!a��q8�PM�r�?�F?Ҫ�=,(ǿ9�s��u�����x�<�-��3i��z�g�f��ؗ=>���4��̱�.c��ќ��Ȍ�����
���l����>�t�=�@�=z2�=E*B<�����<7��=��<�C�<EE��Z��<�F=����`��&���J~�<X=�#7�)�˾o�|?A�E?�[&?b\C?��n>��&>Y�.�%a�>}T���?=�j>ٻO�J���%�*��M��0�޾�վ@<d�T���*�>�5���>6�7>r�>4.�<ɏ�=o{�=�j�=7߇�&l�<j��=*R�=�͓=s�=`#>R>w5w?`��������6Q��r罊�:?�1�>��=Oƾ�@?o�>>@1������f�b*?���?WS�?x�?i�i��g�>���뎽���=;ɜ��62>���=]�2�\��>�J>$�lJ�������4�?��@�??I㋿��Ͽ�Y/>��6>	7>��R�7�1�R�[��b�b0Y��a!?X�:�O�˾�(�>྾=��޾`ƾ 3=��6>�b=����+\�.Ϙ=X0|�N�:=��j=�V�>��C>��=އ��m��=Y�K=���=�eO>�\���M4�!�+�^�3=���=��c>~8'>AX�>�?,S0?�d?e��>K n��ξr��l�>zz�=d�>][�=e�B>�y�>��7?-uD?*�K?��>V�=���>�+�>;v,���m�@�Е��]�<���?oƆ?�>�\<ќ?�ۤ�d>�"ý؝?�H1?#U?�n�>}?���߿� $���+�:J=�y߼,ND�dQ1��	��<F�Ͷ��-ý�����7�>�>���>7�1>f;@>�#|>�߰>�w>6�><�����p�J�c��c���>��;��1�5ս�u<�H�ݰ���3��eWĽ0O�=�D�=���<���=���>�:>{��>y�=���0>/>/�����L�fǿ=�K��_*B��.d�E~��/��e6��B>�"X>�����3����?��Y>�Q?>+��?�>u?�>����վ�M��o)e��&S��Ǹ=!�>�<��n;��T`�+�M�ToҾ^��>e�>��>[.n>U�.��:�]Y=!�澷�9���>`��� ��v����e�pԝ�T����vk��8�&74?�����>'B|?7?��?v�>��d��R׾��9>��W��}�=��TZ�Ք��z�?��2?���>����2���̾�\��a�>�#J�Z�O�y����0���	�s�� $�>���=�оn33��p��쏿\tB��Dq�^K�>C�O?]�?e]a��a��VO�����"��6?��g?,��>6#?g�?Q��2̀���==�n?��?T�?R	>F%�=NϽ+H�>�� ?�&�?�֒?��v?giV��s�>�Bs=d��=���7��=�,0>o>=!=A%?Me?e�?H�g����.�޾��ľ3cy����=�g�=�^�>'X�>�P5>��=��#���x=�tI>���>0�>Ii>�J�>3��>5��*a�n?kC>���>��E?�H�>�O����=i}�=�C��dP��:n1� �q<26��{����=��=�M�:)��>��ÿ^�?��>�����*?��;D;�w	K>�,�=�6A����>"->(:>��f>ܖ�>�2>�Ƨ>�]�>�FӾC>����d!��,C�J�R���Ѿ}z>��	&�����x��BI�Tn��]g��j�R.��g<=��ǽ<H�?R�����k�,�)�g���\�?�[�>�6?bڌ��
��b�>Q��>�Ǎ>K��U���0ȍ��gᾔ�?<��?�;c>��>H�W?�?ڒ1�13�vZ�,�u�n(A�,e�V�`��፿�����
����,�_?�x?0yA?�R�<):z>R��?��%�]ӏ��)�>�/�&';�@<=v+�>*��(�`�}�Ӿ��þ�7��HF>��o?<%�?vY?:TV�+rŽ�3>�w,?^?�@n?�V$?D?P���L'?`Ru>A&�>wj?M�$?�6.?[�?���=0>�m3���=����⮾�}������i9�6�$>�[�=hhR�`�3=$(=�~�������H���=�L��i��=z!H>S>M˦>��]?CE�>���>��7?.���[8�hŮ�"/?��:=墂�P�zâ���G>�j?(��?ObZ?s�d>��A��C��>�O�>̊&>�3\>�l�>�kｷ�E�y�=9D>�<>�ӥ=�DM�P���C�	�~���,J�<�?>��>U�{>卽��'>���Qz�jd>!�R�)���nS���G��2��Hu�VQ�>J�K?�?�|�=]��)q��>f�g)?�l<?n|L?yD�?K=�=�4۾�9��YJ��Q�Ơ>,�<َ��ˢ��ѡ���9�ݸ;�8s>L�����8_>
 ��D޾M�m�Q�J���� �R=ζ���^=j����վD2��T�=�		>����:A ��Ӗ�Jw���
J?�ay=������X�iŻ� �>m��>���>��5��u�б@�:^��Z�=��>�;>�?|�Jz�
�E�Ӎ��5d>�7>?MO?��{?v��bW�}��������MS���!?3�>c6?��>@U=�$��_����[�gk6���>x��>�,��Z���C4پe�	���>�Ʒ>S�=��?.j?�v?�UE?�%?��?Jۓ>�1��2���<&?���?�߄=p�Խ��T��9��F���>�r)?��B�:��>{y?j�?/�&?t�Q? �?��>� �&6@����>V�>d�W�\����_>F�J?ᦳ>wBY?̓?��=>Vs5�ü������U�=�>��2?�6#?W�?֣�>��>VKs��fT�J�>�6a?Ĉ?�|�?�&�=s(�>�43>#�?as>K,�>�C�>�_	?��M?awz?�R?w�>�X�<Ҧ�E
c����m�=W��<ǒ����=��F=9ͨ=�bI�`��u��pG��옽��h�vt=.��<L�����>�,>^E���>:@�GC��'�>�Y�:^0־!����~]�gE`�9~>>��>X�}>�Y���r����>��>��
?�$?�a*?�o�<��W�@v޾]5s�4K�>�%?ЬM>o�n�ȧ����c��5=�p??�R?�����}����e?�@e?�lþ�hE������N���ľ�d?d�>ۧ��ܯ�>K�?��;?�>����0���U>������*#��i�=�v�>k��z�^�e>p�W?0�x>���>��9L�C��������>�ڀ?ZI�?cAu?�O�=\�z�#����y��qᑿU�]?M6�>�|��!?<�dξ�G��f;���t��q���������U٥���$�3�����ν�L�=�;?; s?�q?ɂ^?&� �mPc��9^����T��������nE��+F��C��hm�;����oI��E)M=��~���A�ǂ�?��'?V0�S��>����V��;��B>�[������=�
��;�?=Z=Ìh��..�Z=��  ?�"�>�S�>h�<?%�[�(>�g�1���7�����33>���>�|�>��>��:�0-�E��QIɾ�ń��9ӽ�-v>�}c?��K?ٯn?�b�l1�/���d�!�(�.��=��6�B>�o>�ɉ>\�W����|3&��R>���r�������v�	���~=�2?�4�>��>�L�?#�?*i	�?h��_Yx��v1��5�<�(�>�i?W=�>���>��Ͻm� �<h�>ȏr?؇�>cU�>�i��@h�-�s��
w���>�t�>?��>�-_>c;A�_�a����8�����=�|b>y�m?샾�p�픑>�V=?29���M����>L��{�(;˾�(��n>�r?Ν�=�	�='=Ӿ��� Ʉ�ĎO�wE)?R?�Ғ���*�!0~>�$"?��>�:�>b,�?|@�>�Jþ�E���?&�^?�.J?�IA?=�>�=�G���OȽ��&�-i,=���>	[>�-m=ߌ�=����\�1W���D=�κ=o^ͼP��,�<�ܴ�O<}�<b�3>��˿��M�D$�1A�v̾�t$�����"5���R����款���7�r�8^�n	C��g��AA��ڛ�/|w��:�?nt�?_"S��Z��v����z�����6�>�W�(KT�豵�R]�����L������h��J=���G�9Q�O�'?�����ǿ񰡿�:ܾ5! ?�A ?6�y?��7�"���8�'� >|C�<%-����뾬����ο?�����^?���>��/��q��>ߥ�>�X>�Hq>����螾�1�<��?7�-?��>Ǝr�/�ɿa����¤<���?/�@&�4?|���` �i$�=�Q�>��?���>�m4�!�!�����A?�ѧ?0�?̟��$!J��'�;}�b?�	�=u@3�cސ<�� >��=#Nb=�䷽�Z>{h�>
j�m�e���R>�f>�ۨ��>�L3\��=���>�m�>|�gӄ?Hn\�8f�o�/��P����>5�T?��>Y�=��,?�5H��|Ͽ��\�<a?�0�?���?4�(?�忾�Ϛ>��ܾ)�M?�>6?��>�\&���t���=��޼z���+���V�	��=��>�>،,�����XO�+���#��=�}���ÿ�1�5�.��A>}�=��l��zn�Г��ӱ=�n���3z�[$ӽ@r=c�@=�1>9,y>lҭ<�Y�=3sf?�6\?{Z�>_h>��-=�3y��0ľ�1ƹv���5W4���þ��5Z��y5�P���!�����5
��\þo�6�k�F=,R�����7��gk��OH��,?W]
>>亾�vI�����ݴȾT���	��������i���p.��Vi��@�?�C?�����[�����y��ݱ��.Q?82�L��ܼ�,�=J|�fҝ<T�>��=��վ�t&���H���)?�@?͕þ�|����I>�٠�(��=��#?�W�>KP=�.�>2�,?�@����WS>C8>��>x�>N2�=����Y�n!?�M?�������F>-ľ��Y�I�u=��=]7^�M�O�DP`>��;�ޖ�T����H��1�o�V?	��>E�)����w+���i��fA=vx?n?��>��k?-C?+�<�l��a�S�G�
���x=§W?��h?�>�`��IBо�����5?cue?J�N> h�&
�=�.��;��5?��n?O2?M���+D}����R���76?��q?DUT�Z)��+� ���7���>+�?V>�>#�6�w�>�2G?��轈��Fн��4����?�*@{8�??Sa<I*���=x?hG�> I���̾S��~J��๜=��>z߸�9�v��x�$:3���,?_Y}?���> ]���d�~��=�ԕ��X�?�?|�����f<��l�@l��Q�<�ʫ=A?�>o"�_���7���ƾ+�
����䠿���>�Y@q8��&�>�H8�x3�;QϿ����Yо3Pq���?2��>:�Ƚ����j�qMu�ųG�<�H�՚��Pݱ>_�|=��'��|Ǿ�����1J�7����>3����>����,ܾ�����k�W�>���>��>g��IH���}�?T��!ÿ�����6�M&�?=�?:dr?;�0?���7�&��������wK?�p�?�6u?�T\�9U;��_>��h?�����YT�؂2��\U�,�O>1D,?�x�>k�9�u�C��E;=b��>-,>Gx!�Oz���ﱿ_� �u��?<��?1}���I�>�؟?��8?W���Z���!���H%���4=��T?��>:�߾�%�`~H��C�����>�?��潝�%��qi?{pl����(2W�@2¾ �>- K��ާ�~�=1JR��X���S���<Y�5��?�@�+�?��������Q?=��>3x��f��%S�����>�(?���>2��{�u>�:����v��=�?e�@U?]ߕ�����>��?u5�>7�?N}>.$�>�,A=�Y�0��6��>S�z>~*>���>�o)?���>}!���9��0 �3lA�@R�m�9��G�6��>��Y?�`?���>th�օ:��1�>������������Gm='��%�=��z>G�>U����x�?�l�O�ؿ�g��
i'��64?Ń>�?J��!�t�c5�B@_?�z�>�6��)���#���<�7��?E�?"�?��׾�[̼�>k�>WN�>�Խ5;����7>��B?d��D��.�o���>Y��?8�@&֮?: i��	?z��P���`~����7�R��=��7?61�Y�z>���>��=znv�������s����>�B�?V{�?���>��l?�o���B��1=�L�>�k?�s?^o����B>p�?
�������K��f?��
@Yu@��^?���a߿�����F��o �֗r;�ȴ=7_>vy=��.>{{3�O�?� ����m�=�m�>U�_>X�:>q\�=�<�N%>�F��� �<���k˛� .�����d*�
ɵ���ƾi�����GӾ�ѫ�>��;_Y����:��?�L�s�����=j[[?�W?��h?q��>�}!��T>ܥ޾֩=�
ν9�n=yЄ>�j3?[>?� ?�ߍ=L���Ha����{�������>_}>EP�>�n�>J��>dռ j> �5>��>->F�]=��V���<�~R>�K�>_
�>��>�D<>�>�δ��1����h��w��̽-�?с��ֻJ��1��[9��l���2g�=�a.?Wy>���?п�����1H?�����(���+�!�>��0?cW?V�>����T�)9>����j��_>) ��|l�@�)��&Q>1k?�!}>�$�>�g�<�>�!�R�� ��4T>_�G?�����(wh��B��˾�>`=�>�Bz��j-�ډ��*뉿`��#�=	xB?��?g��9U���b��W���>���>h=�:=7vy>O��]�����@�=�A>�6i>�s�>�s>GV���K�>&��Z�E��&�>Y#>Σ
>FhA?�|??�v>�m�� ����ynn>�1?Ru�>|1]<Q@H��=���?>
Z>C���F��͞���P����>ֶ��s�޾�-Q���=O�<H��=6���p��g
��#N59mɇ?�ȸ�����:�D���ۼ�?P?$�>���>f��=��P�玦�W���!�?ys@Ć�?�"���k��,[?2b�?6"��8 >�+�>�A�>ᴱ��$0?������j/�Ak��s�?eך?�z��%����Q��R�=3�0?�:���a�>Cl�IX�������u�>�#=��>�1H?�U����O���=��|
?_?�]�q����ȿ�vv����>��?Q��?��m�eC��E@�R��>ß�?�gY?�pi>�x۾�xZ�?��>��@?{R?��>�2�~�'�1�?�ܶ?���?��I>t��?�Ds?y��>�y�WD/��	��ߌ��&~=́};%J�>�%>����t�F����[���j�S~�Ac>Ko#=�u�>=7⽭}����=󮌽�:��{�a�e��>�0r>�IJ>���>
E?���>�Ƙ>�=�ۏ�X ��A땾�)D?���?�{��p�	�b���>j�h�ؚ ?t
#?hM�=1Ⱦj؁>�&J?��]?�J?9�Q>�c"�v9���Iƿ��;o]�=~e�>8��>e�?<���tc>��|z�l?�>R�>�}��9��莾�mɼt�>P�%?���>�>�X$?�=?�K>
��>�4N����������=���> |?��f?��3?GH��@�4���������l�3>��?k�?S,>�e�*���L�7�q��~�x<�H�?A�\?a�3�G@?>L�?�.?<B?�Oi>���j(Ѿ�k��-'�=��!?���̣A�%?&�]��@?�$?�~�>0���O�ֽ^�ּ+��;���_�?H<\?gt&?�v�m%a�h�¾���<��!���N��4�;�1C��>��>5��0��=�">��=@m��[6�Ըj<E�=:y�>1��=��6��/����1?�t =D���t� >��V��<�ɞ2>9=����_WH?f3��mn������}��r;{�_��?_��?�Y�? �߽pd�"�V?Dso?�?l�>�ޘ�4�̾N��70��a[,�u����>B�>������Ϋ����~È����=@�����>4.�>6�
?~��>��P>1p�>3S���/%�������]�6Z��8���-����	��FF#�� �'þ��{����>��x����>7�?QUf>6�w>�k�>�MN�.��>�,T>T�>�F�>�JT>�8>��>x�9<\Ƚ�\^?�Z�:�6�����'��N?SYM?Q
�>����f���2�8�?�?��?���>jQ��~"���>?�Q4?�����LI?n9<>��m=��˽���HL����H�M�1k�>+��5�/�3�~�QC	���>��>���=�ľR����p���n=10�?��(?��)���Q��o�%�W��S�t�Hh�h����$� �p��䏿}U�����~�(��\*=v�*?�?�g�����d���k�?�KBf>��>��>:��>WvI>��	���1���]�*'�ި���K�>�N{?l�=>Ǚe?��_?�`?�T?�5�>��>�Nd�
D:?9S@>aD�>���>�68?Zn�>U�>�?�s?>��=փ���������;?��=?^9?��?�c2?��¾ڿ;�V(�R�t>�	G���+��x#>���=�쀽ى⽇(=	ǡ>�,?ь�l�8�T����k>s�7?��>�L�>Ϡ��U0���g =�s�>r�
?���>������q�k�����>ς�?���k=R�)>:�=��z��p�����=�&����=i`���4�o�<@�=Q�=9����V�9d�h;��;4��<
t?�?&?�eT>Ń�>H�d��U���g������^>n�K>@�>�پ���V��f�p�1}I>�V�?��?f��=�><=�ŋ>� ��Yf��1�
�ڬ�J�=~K�>���>�T?�܉?�Y??a�A?�(>L�0��Ә����H���8?�w,?�ԍ>I�
���̾,Y����-��K?7�?�.c���(�Z�+�p�¾�V���
>m5,�X�}�E	��#&6�^B�<���������?!��?Rj���_2�~u�<E��ß���I?��>W��>N��>�i,�k�e��Z���$>+9�>��F?�!�>��O?)7{?��[?�_T>$�8��-��&ҙ��L3���!>;@?u��?,�?yy?�t�>��>��)���Q��D�����₾]�V=�Z>j��>�(�>2�>���=Ƚ�V��T�>��h�=Čb>v��>���>���>�w>ِ�<�!P?���>�/���ʾ�O`�>��6�����&?:�z?k�>`�ƽ��B�^���J��`	"?��?+�?�Y?��CM>��}:�����?)��_�>@c?���>-��=��M>
��>]��>6N�>�&^�hi$�c
9�����w�?k��?�/�����$��̪�<�U��?����P����<�����>m����	J�,eξ�n��⾱�ݾ��j�=��O�Ծg�-?؊=�ӂ�9�>>K�s;H�����=�����X���=��a=�����@{�;�������0��=��=�0�<J����?�Ή?tR]?�xK?��>D±>�νY��>˙�=��9?�f�>��B=𜘾��'�e���I�Fξ�j���o��Ӿ�a�<5�a� +�=���=��=�t߼j�?���׽{B>2H
>��1=�|>Z��=��V�(��<�>F�B>�w?�h�������DQ�*���9?^��>Ћ�=�4ƾ�??�t;>�F��Li��h8�Q?Q��?��?�_?�g�� �>_��������=)O����5>>�=�1��`�>��G>���$���/��� �?��@@?����JTϿ��1>�m >1'>kV�́"��%1���ڽ�X^;]3?.�J�`B��2�>L�>K!��pcվ5�"=��F>���=1��D�C�u�>���݀��`]�=��>��>b�j>�rJ��+��k5=���>&u�>F����	{�DI�<���=��>���>:>;�>>�?.?E�`?��>�����Ӿ��ž��>�O�=}�>�Q=��1>�j�>R:?J^J?R�K?!u�>b�=���>�ʥ>�Y*�~�k�6��9��0�<k�?m��?޽�>jR<R�9�����:��hȽ��?�1?`�?�۝>;���޿��'��&5�ņ�U�/;5��6�MY�Y��c_k��	�E���= ��>'M�>(�>��p>�>�q6>��>	�=���y%�=�'+=�D=C�s���0=	�'�(�=sU��
<u];14i����y��;m��<��B��<~����=���>L1>��>��==���*/>iٖ���L��̿=A���(B� 4d�!L~�3/��_6�S�B>�QX>VY���2��s�?�Y>}o?>�|�?�8u?��>CC���վRI���+e��9S�y1�=6�>r%=��~;�\j`���M��YҾo��>a�{>Cu�>�?s>z1�\�4��Rb=�ȾM�=�$b�>f����J.��Od�����ݞ���k��˰=7�B?�Ά���=���?6\?��?{�>{�޽�5��.:>}B�ߐ>1*�{6�������)?�6$?��>T�(�K�M��+9���U�>�Gg���E����!]8��?�;�iþޘ�>�`����Ծ�f.��+�������8��G�@v�>ųB?�J�?�#��m��	X�x�&��o����>Q*[?�1�>�%�>�8�>d� �LE�S1����=��v?��?c�?X%;>㈲=�(��F�>״?�m�?���?�o�?��>��L�>i��<�M�> �=I1>Qט=r�=xF>`�?�_?y?��7�%��������f�1��@�=p��=���>�L�>z�>�T�=K;d=�3�=[JV>���>ތ�>�@m>��>�>�>1*���>���#?F��=�> 1?7��>�rF=�V����)=()��Y.����;L��������<�-�ǝQ=,��x��>��ƿ��?�P>M%�Bu?���v�4<^>�!V>��޽���>��O>쁇>O0�>*o�>5�=��>��7>pAӾ�r>���_!��#C�ہR���Ѿ�mz>P�����%�b���?��P,I�pn���e�Pj��(��o9=�Й�<OF�?q�����k�!�)�����G�?YO�>6?�挾�F��7�>���>~��>�N������l���wX��?���?ߊ�>�ʄ>L�H?��?d��R�޾o�y��Є�?>����]E����������v
�mmg>���?T�e?A\?qV��$g�>��d?����+� ��>�`@��`=�=���ށ>a��΅�ή���I����}��>H-�?��w?���=�~v��ֈ�3��>�sL?�^\?/6?n�3?�=,?>�ɾ��B?�Ʒ>�D?
�
?@#?��>��|>����K��=+Z>K*={���RM��n��'��vt���)=��H�W���T�l3�<_ ���T=t�<��ݼ�FZ=ٚ!=�x�<%+�=�!�>��X?���>g~>�/?O�P��t<��ʰ���+?��<�r��$����v��`3��0>?px?�׬?ouP?�TE>"8���5�Jq>$�>I�)>kc>a%�>�L��:��K��=�k>�T>0�v=o�.�<Ҋ���>w�S�b=�>F��>�6x>o���) >D&��~�w�pf>��G�ey���a��kI���0�o��k�>x`J?/y?���=�w���x���e�V�)?��=?$&M?Vh?��=zH۾�8�`vG�l�t��>{<S�
�����2��o9;�A�l�e�r>�Ġ�q��� Z>:���ݾ�g�t�I����d>=����Z=���r{Ӿ��{�@�=���=��uM����T��N'K?޲a=����(}X����3>K�>�>�|����|}C�4款AQ�=�I�>��9>eYR�]�龛$F���;Y>��_?��f?ks�?������p�A�=�H��Jhu���<�9� ?r|�>z�?kS�=`��=��ɾ�0�����L�t�>g�>�+ݾ��g��*��AM��A�!�Fk�>�	?��[>�S	?��?��>v?vn-?,+�>���>��ʽ�c��
&?⤃?�ȇ=TkԽV�U���8�AF�8�>��)?�BB�t|�>�6?��?)�&?�\Q?�^?��
>*��Z@��q�>��>_vW�^��|�_>��J?Y��>�Y?ƃ?�>>�(5��Q��d��D��=��>��2?S?#?$�?'��>��>$���ۀ=��>3c?�3�?�o?0��=��?�G2>�7�>@�=���>���>?�2O?�s?��J?���>�l�</��aC���{s��-M����;�G<��z=���Ut�?U�3+�<�N�;�$��
��#�񼉫D�I�����;dB�>�G>@�f��G >�5�+c�9�T>����mǾzv��E�N�i	�=�^�>�;?�)�>.G��=h��>~��>X2��72?�R?�$?�b#<�S��"�!�@���>(P2??#�=a�z�����W;y�-H_=��s?=�\?I�7��HɾG�b?�]?)h��=��þ��b����`�O?<�
?3�G���>��~?b�q?B��>�e�*:n�,��Db��j�'Ѷ=\r�>BX�Z�d�|?�>r�7?�N�>`�b>H%�=Xu۾�w��q��b?��?�?���?+*>}�n�U4�k�澣���ʲd?�>{̾�)?
�������z	��O����[߾�*���E��d���h���wJ�r9|�C��x^
>�M?��t?Z}t?�~^?m����_���h�ߥy�\�O���L���Q���K��[B�ܫa�O� �˾����A��=~��bA�r�?LK'?!�1����>�䗾�C�4�;��?>�����Z� ��=������:=��O=bh��-�c���'�?�)�>���>7�<?�!\�Sm=�P�1��u7����ZG2>�F�>�4�>�C�> ��:��-�|�<�ɾ�2���"Խ��k>x�i? �N?��i?9K�)�/�v�����r˼�-��(�9>d��=y��>�\���E�&��D�uf{���5���A��+�=r�$?><x>KI�>{s�?:#?~������E�c���4����;
��>��d?�J�>Q�>�ӳ�ٰ�V�>�+�?�>��>b���Z�Q��/1�i9����>�E�>/x�>Df\>����w����a����p�̻5��2ż$�?�}��ֽո=>8]r?W2׼�9���V�>=z�<���� ��E�0q�>�#?:o�<�ZT>LȜ�@�[��Ɠ���l��@)?�G?(ϒ�]�*��"~>�*"?���>s)�>�.�?�7�>�þI63�V�?C�^?BJ?�CA?��>�$=����NȽ��&�^,=�l�>�Z>?l=��=N�]s\��f�2F=;�=��μU]����<%��R�L<gN�<��3>ƅӿ&GG�a������¾c��M9�����Iz�<
��~;�+��k���7����)S�zP�$y��U7�5T�?�L�?1C����������}��&�[��>�w��瑼�ه��Kƽ���&��V��$
���L�&gR�h!N�O�'?�����ǿ򰡿�:ܾ4! ?�A ?8�y?��7�"���8�� >oC�<�,����뾭����ο@�����^?���>��/��n��>إ�>�X>�Hq>����螾�1�<��?6�-?��>ǎr�0�ɿb���h¤<���?/�@��Q?}�U����f�<8b�>�?�>��^>��>=�Y$�����}�>�=�?���?(��>��=�f	���W?v�E>N�l�{�]��Z�>�lK>B�(>V����A=��>w����Ӿ��=IbG>|ѻ>ӈ��kx彿,��t�=Qj�>��]�\�,�5Մ?'{\�{f���/��T���T>��T?�*�>/:�=��,?[7H�_}Ͽ�\��*a?�0�?���?*�(?5ۿ��ؚ>��ܾ��M?UD6?���>�d&��t�!��=@6�Ԅ��g���&V�{��=T��>a�>͂,�݋���O�I����=����+ƿ�5%�(��/Q=!໻H�h�
e�7���z<J�^0����m�t�/�e=`��=��O>	+�>.fT>.�Y>�qW?�>k?$��>0�>���⬉��Ͼ6+��D�������_���1����f޾�	�ޏ��'��8Ⱦ<'?����<�OV��!������Ni�)�F���,?��>	ʬ��)S�$�<�0������T�����5�����1�H�`���?�K=?�u{�k�T����#���N���c?-�ƽ���0٭�/��=�����<2��>��=�G۾s�$��	;�*c0?�3?���ꪑ�g�)>-v �Re=��+?�?�_E<��>�*%?+z*�ۅ��Z>�M2>�ƣ>���>x	>�N���Fܽ �?O�T?������F6�>�6��k8y�Bh]=>
>Y�4����:?[>ݺ�<�����a�O̒��;�<(W?���>$�)�0�b��F���h==Ʊx?%�?�)�>^yk? �B?j�<�f��c�S�� ��cw=�W?X)i?ö>p���EоL}���5?��e?J�N>dah���x�.��S�X$?��n?u^?٘���w}�Y��T���l6??�v?�K^��g�����.eV���>\2�>D=�>t�9�^P�>GY>?=#��R��>����I4��̞?��@e��?Ĉ.<q? �2
�=75?���>�O�+Rƾ��U;���r='�>F?��S@v�5����,��?8?��?8c�>I�������=�ٕ��Z�?�?a����kg<��l��o��]�<�̫=��D"�F���7��ƾL�
�����ȿ����>Z@�O��*�>sC8��5�9TϿ���[о]Tq��?�~�>I�Ƚ監�i�j��Nu��G���H�_����e�>���=��罣����9~�9�,�׽jF ?
υ<H7�>��r�g˾O�����s��>�X�>�>��g��d����?5��*ֿ�Z���"�4q?�f�?�v?Z=!?7���������r�.� #T?V�?�b?l.��k��A�/��)j?(֪�&^��y4��VF��X>�3?��>7�.�c`=�Z>Bb�>�C>��-�N,Ŀcƶ�j���ͬ�?	�?A���I�>1��?O+?C'�:��M���E*�K����??��2>-Hþ�"�!=������v?О0?Μ��y��rl?��u��y����K�T!�	`�>Ta6��j��,�=�4��j��`��y圾6c�?]@=�?����� ��DE?��>%�����྆�ֽ���>\��>\��>6��s��=G;:�&[��6>5��?�N@�4?fq��E���|>p�_?Z�>3�?���=�j?L�=�ҽ�a;;�Z>q��=-T�T/ ?�M?��>�(�=J���*���I��ZU��� �8�B�`�>��b?��I?��[>_��(>��Ȇ�Ƚ��]0��yX�x,�yo���U˽��8>N�6>c��=�QX�(�޾��?Lp�8�ؿ j��p'��54?'��>�?��x�t�Y���;_?Nz�>�6��+���%���B�^��?�G�?@�?��׾;R̼�>/�>�I�>[�Խ����Y�����7>1�B?^��D��u�o�x�>���?	�@�ծ?gi���?r6�Gʂ��䂿��
��t�a���_H?�?̾���>Cr�>�u=6u������n���>�W�?�i�?-��>)�?w�y�[RQ�ز�=��^>�?�?-�)ź���=u��>�*�pC���'۾��s?��	@(�@��R?GZ��7�׿�덿wx��[C���$�<%��=mk7>j�ܽ*+l=j��<S��c��=��P>�<>�4>H-">$�?>.��=_���uꝿ�ʔ���9�H��А�&�q��V��?���5�D߾�g�������c�8)��<;���,��[��	.�=y!a?�Y?��d?���>��M��8>fH߾L��=��񽈧�=�U>��)?��>?&�$?�&@=0,���p��~�|���^J�����>��(>L�>�]�>�~�>�c=]b>�V>x]�>��=��<�~�<�=-�V>�6�>�q�>j0�>�B<>5�>;ϴ��1����h�Dw� ̽�?{���/�J��1���9�������h�=
b.?�{>���?п[����2H?����)�'�+�n�>O�0?�cW?�>�����T�	9>U����j��`>�+ �l��)�_%Q>|l?�f>�#u>!�3�fb8���P�Qu��af|>D26?鶾�S9�t�u��H��XݾFM>ܻ�>��E��l�������kri�@L{=)w:?�?�f��Ͱ��u�s2��ZR>;\>њ=,J�=eTM>�(c�D�ƽ	H��`.=���=��^>�?dB,>@Q�=�΢>�y���1N��ت>!�B>�%(>}�>?�L$?Z0�/��$���.�N�r>L�>�h�>�F>T�K��ͪ=�q�>�d>���( v������>�~=Z>�˃�t�[�~+o�G�~=Y���0��=c��=8�B�?�Wv=tw�?cp��7�����*�޸�=�B(?y�>��>W$=��O�U\��0ް����? �@��?+�#�D�:��wH?�*M?��Ͻ#p�zq?��?�/�s�Ͼ�w�>�};"��������=��?RM�?ߍ��ﻛ�����
y>��W?GK>�Mh�>�x�Z�������u�m�#=N��>�8H?�V���O�y>��v
?�?�^�ީ����ȿ.|v����>S�?���?d�m��A���@�p��>8��?�gY?|oi>�g۾8`Z����>̻@?�R?�>�9���'�~�?�޶?ү�?|>��??f?��?�@��p�C�N���������=Oh#�4H>ށ�>�Ɛ�QIa�}׌�!Jy�P���O%E��>>0����>���=>����<�f=U0�-g=4��>aE[>��>��T>f�?���>�>�|���齒顾g�ݾ�K?���?R��y2n�H>�<
��=��^��&?�I4?2b[�3�Ͼ�Ԩ>��\?&?�[?Kc�>����>��)迿�}��o��<��K>�2�>_H�>����FK>	�Ծ�3D��p�>LЗ>����?ھ�+���Q��~B�>�e!?���>-Ԯ=Й ?Ҝ#?}�j>�(�>:aE��9��8�E���>���>�H?��~?��?�Թ��Z3�����桿~�[�A;N>��x?�U?�ʕ>N�������hqE�5DI�4���H��?Atg?�T�1?42�?��??$�A?w)f>,��ؾ����&�>��!?���A�aL&�z�f?Q?���>�=����ս�5ּ��{z����?o&\?==&?М��)a���¾q,�<�*#�(�T� ��;cE���>�>������=3>	�=%Pm��E6��f<�f�=J�>�=F-7��m��w"3?Jj=������=Q�Y@��?>�#R=�u��K�L?��x�e_p��߳����"��==�?>�?K��?,�K��$f��nR?aq�?�}�>��>��ʾ3[�dz����ݫ��ܸ�g��=ⳮ>�K���b
��\��nH���rr����<4��l�>m��>��> ��>�E>$��>��Oz2�?��d��	JM�����/��/��="��%��/~���8һTC˾{�����>�H<<<�n>m�?��">�t>�E�>�bT��7�>>^>V��>�ў>�l'>���=�d�=�ǉ��(�8�^?Å����HQ�,�߾w`�>��V?Dj�>�����������{D?01�?���?�,>}�\�,о.�+?ds�>
 ��I�X?HT�>zt�R��x����ټg���^�����G>h���L�H��߆��pȾT ?�P)?Tּe]��ݢ>q���o%o=SK�?��(?�)�A�Q���o�=�W��S�b~��@h��_��5�$��p��돿5]���$��.�(��w*=�*?��?���6�,��<!k�^?��zf>u�>Z'�>2�>�iI>�	�I�1�a�]�K'������O�>�V{?{�>��I?[ <?4tP?gYL?��>��>+����>u4�;Z?�>���>�9?{�-?920?�i?�T+?��b>�J������ӑؾZ�?��?�F? ?�?����'ý�S��Wd��ay�lz����=NR�<��׽�Bu�N�T=N
T>�?�"7���������p=�>?*�>8k�>�B���k�����;J�>��?�6�>�O�iH���6���>.q?�<��rӼ�$e>0��=�Խ[>J=ߘ6=s��;ݯz=\"_�2��;����9*�=&ݎ=�l��N��<�
o��9�]�=K	?)?z}>��p>�k��K�]����͵p>�Ʉ>Kܼ=������+���F�v��s�>�~�?���?ϕ�<ެ_�`�>l�L�����d�c�΍<�.�><c�>�DN?,˛?8'?��!?}6�==N�9���j2��թ�u�C?�,?Hv�>�����ʾI먿yo3�|�?X?�Ma�-�A>)��¾��Խ�>?]/�7~� ���}�C�,Ё�=��7���!��?Ͼ�?�C�r�6���U����%���tC?�4�>�B�>�>Z�)���g�j(��:>N�>��Q?��>7P?�N{?&�[?GVS>(�8��������*�f�!>��??���?#܎?\�x?d�>�.>g�*����?������F�噂�q�R=��Y>��>	�>��><��=�<ƽ�S��t�?�{��=lJc>�v�>��>�%�>I�w>���<�.T?1��>�o�������5��Я����-�ŋ?\a{?��?��!��\���d�PK��?�>�Z�?@(�?�
<?F%��I�=�3�<a���������>*��>�P�>,u=�v>���=��>���>��K�n�8�bP^�J��ŀ?W4V?9�=�Fп%�J��������T��>_魾]��|����Z���>/�ʾ�̽��++w�R���ʎ���&!پĝپ��?J�8�e#ܽkeg�G�K>~��a͎�@#>�=��>mْ�6��=������a=�����:
l�=O�M��=�Ν���?]�q?l�?���>ړ�>Ui�>MU8>'?�y>�6?~�����q����e�L�����H6��g�ս)���>+�:��>��]>Y��>�5�>E<�3g>���<�%�>/� � �2���=�	=���=c�->���>~R>�y?��������8 X�NE��.?6{!>�]<>S
���M;?���=D~��]������c�?W_�?:��?���>�b��>x���v��^`=��`����>F�z>�ka��k�>��<���*ǟ��㗽�z�?��@KN;?N+����Ϳ�RN>�7>�>J�R�(�1�ݿ\��b�YfZ�7�!?�K;�BZ̾�+�>��= ߾��ƾ]:.=�]6>�Tb=�W��Q\�	ݙ=�>{��<=Bl=�É>��C>9Z�=[��|��=v�I=w��=��O>������7��F,���3=���=n�b>R&>��>�?N2?��a?s�>�3w��SѾ辱�c>��=p��>�F�<�*�=�K�>��L?@^?| Z?���>=t�	��>�L�>��8�9�S��gξ�P��X��=8�?)B�?�(�>�x3���5�I��r4�+d%��%?S]9?��?O�x>h��Z=տ=�s�5��c���G�;����`��?7�������]�-�㽽۸=$��>���>��>��f>��>�$>���>il�=�$�<���<�!1=�Jg=�Ž*��<�D��j�=��j�I��=k��<k6���GҼ���"r< "׼N�ͼ^,>_N�>�Q>��>�Ŋ=�ᶾ$�j>�\���X�x�<=ӽ��G�9���Z�zpt��-�.�J��?>�>B\���|���� ?�o>��p>�c�?py?�3>{ؽjE��y���WYK�D���=ĭ=+F`�c@���`�%TU��P㾲z�>�n�>mj�>�V�>�+�j9C��Ƥ=���$�5��~�>�R��$T�[�o�u��뤿�J���g�
�]�kEJ?������=k]v?��O?p��?j�>0$Y��0ɾ?�)>X���Y�<ٝ�P�S��o���)?9�$?6/�>k���*2C����r�ܽ6�>:{��L6� ��
S��Y>�q��t�> �Ⱦ頌��y*��U������5C.��cP�lۧ>��`?��?p>L�iG�>^?�:`F���>=%�>�1^?1�>�\?M?lRW���Se�����=C�m?���?�0�?q�>��=cի����>�
?u�?��?;�t?��9���>���;'+>����c#�=I�
>��=eU�=�P
?jR	?yi
?�0��ߴ
�����mﾭjX�E��<W�=L��>U?�>�Bk>q��=8�=a�=��[>ޜ>���>ռc>���>��>�B��ҽ� )?&(�=�K1>+�3?���>δ�=��W��� ��$ $�j� �������s���B�[��=���\2�>W2Ŀa��?��>���+"?<X���;��A}>��>h�%�8�>�z\>ֹ}>�@�>Mv>�ܵ=]&O>p�>��Ӿ�E>5����$���7�%,X�>پŚ�>uW����
�L����ν��D�q���5A��e�U2~��;��'=~s�?ͽ��\��w+��	3�Z�?�;�>}:?V!��u@���%>���>�b�>H��C��k܊��}�<u�?I'�?-V�>k�w>��~?��?����'B�v�d���n���g�R-��o�\�ǩ��$t{���о�71>o?*�?\&?E�(>���>��_?m �r�����>��B�&��+����>��R=S�����}��6��xB�$� ?5W�?욃?��>)Ծ�r�<[PH>Jt�>'GR?��V?dAq?b\`?v�=Z�1?�X<>7�?��<?,7?�?��?v��=Rw��M��d�>r����q�-i9�ڕ��q�=f��]����~�hZK��<�!9��+
>�[�=�F���Y=�tW=W��=�� =�����>�sZ?���>�`�>�u6?��`�5�O���5�.?/�,=�?���������73��X��=j�o?6��?'~]?�aD>�fE���)�s2>Y}>R,>�\O>�>&ٽ�86��ŏ=�>ő>a��=qW������
��덾u�/=*�>3� ?a>�4-��1�<�đ�r����t�>�C1���!j��sxP���&��e���>�??f)?T_�=_K��W�F=��m��y5?h�E?�;?<vn?֭M>�þ�B��d)�z�,��y>�2J� {�,
�����(]D�[��C.>�詾�2¾�S@>����=Ծ"I^���M����>�������<\���ٯ���f����=���=ﹾ9!�mb�������A?Ve@=������X��0���]*>��>ٷ>Y�
�O��ʅK����;(L=�>��6>k���6�龇�C�=|���=�>oOE?�X_?�k�?Q#��,s�@�B�õ��Hb��5ȼ�?�p�>�f?�B>-�=�������d�HG���>��>����G�{9��\0��t�$���>@<?�>(�?P�R?j�
?��`?f*?�E?.�>�������A&?7��?/�=Z�Խ�T�| 9�?F����>}�)?�B�ṗ>L�?�?��&?�Q?�?��>� ��C@����>|Y�>��W��b��D�_>��J?ܚ�>o=Y?�ԃ?��=>U�5��颾�֩��U�=�>��2?6#?R�?>��>i����5�=��>�c?@�?�+p?Q��=��?L3>x��>$�=>ݚ�>�?�2O?X�s?̼J?�o�>�|�<'�������Eu�kH���;iUO</�s=a���{s�s��.��<c��;�.��hr����1E��ꏼ�o�;�>޹i>�ҏ���4>Yʾ�����>>���=o��J����:����=�@~>2�?�>�>�&*���f=��>'��>�2�t9&?�?n�?x��<	Vb�Y�I�Z�&ܱ>ZZ??��=��i��瓿F|x�?=�rk?��\?�(U�m��G�_? rb?����[+���ľ��o�Z�ﾻ.B?�_??�+�D�>�z�?p�j?1��>�o��oy�;d����a�ߵ`�I�;=���>#!�4�W���>U(8?�n�>>>�dc==K��I�������0�?� �?u'�?���?�>9�q�h�;��ԧ����Y?���>e����?up�;������+��-�Ӿ ,��ӏ����������?#��2���{�p>�=�P?Bg?��g?dh[?�7�Ybc�=a��~�?�R�:��
���=�҃D�PA��k�wi�:^��M��wk=:�n�t�=���?d�)?l�:����>X���n���׾��3>1���t�C��U�=�ɘ�6�E=�M�<�ƅ����@�����?�o�>��>�zD?�LN�BJ<�vE8���=�]BҾB60>���>q��>��>��^�$�2��zĽ����g5��Oզ��u>�;d?p�K?�*o?TH���0�+���:!��(1�HR��UC>��>�!�>FY��=�ra&�	�>�LFs�N%����^�	�o�=7�2?5=�>���>��?��?=	��g���u��N1����<�=�>�h?��>�/�>Z�̽�� ��
 ?ȡb?��>'w>ҮѾ�K��j�0V=$��>�M�>�MD?��?�Ǫ�ʔZ�ו�������>�v?8D��xz�C��=��?;���Ǩ�=��?>�1�����Fp��bP9�cQ�>V�?!>�T>����d��BC���;SO)?UK?6璾�*�?6~>H%"?̂�>�,�>-1�?,�>�nþֹC���?��^?BJ?'TA?�I�>,�=o ��9;Ƚ�&�h�,=2��>.�Z>I%m=���=����u\�8w�d�D=�u�=q�μ�L���
<4����J<O��<�3>�gۿ�;K�\�پ�����d:
�{����OU��ݗ�ub��J����Jx������'�hV��?c�O�����l� ~�?C/�?����A���'���9���Ě�>F�q��w~��竾�������ྣ���hX!�H�O� i�ߪe�8�'?�����ǿ鰡��:ܾ5! ?�A ?$�y?���"���8�� >�C�<<-����뾤�����οQ�����^?���>���/��%��>ե�>��X>Hq>����螾Q7�<��?&�-?��>�r�!�ɿR����¤<���?,�@}A?��(���쾃V=��>��	?��?>�S1��I������T�>j<�?���?�zM=��W�!�	�!�e?ʃ<��F���ݻ}�=n;�=�E=���ɔJ>gU�>���SA��?ܽ �4>Fڅ>/}"�D����^�4��<$�]>(�ս�;��yՄ?��\�mf�g�/�ZQ��e>>�T?�5�>�
�=W�,?�6H�t|Ͽh�\�D1a?�1�?��?i�(?Pٿ��>�ܾB�M?�D6?��>Sj&���t�S��=�B��]���㾷%V����=���>��>��,���s�O�f������='���ƿ2�$�m��=Ẏ�[�X(��K��;�T�02��<+o�Գ��Uh=���=#tQ>�E�>��V>��Y>�jW?�k?��>6P>2�㽆����3ξd���>��\k��������ϣ�TO�B�߾�w	����N����ɾ!�E���T=-sM�����x�e�yI�x�?!�
>�"̾��D���P=�������:���Ι�?�̾0K5��p�Ԅ�?X7?!s��;)S�b
��6������O?�T�{>�Lݾ��={���Q
=���>w�=µ�3!4��O��z0?k?�	��K⑾�<!>ԭ���=��,?���>|�<'��>H�"?vz,�$Z㽱�Y>kK->,��>�e�>!>�ﯾ$^ؽn�?=\S?*Z�ۛ���>֣���gv�x�k=�>vf2�(@ܼ&X>��V<M^��������<^>W?d�>�8)���������-��>7=*x?H?r�>/�k?��B?۵�<�I��g�S���@~�=�?X?T�i?O�>��{��Ͼ픨���4?��d?�HL>XFh����TF.�^���_?�~n?�?K����}��'���R�m�5?6�v?Om^�Ko�����w�V��9�>�R�>ڲ�>s�9��\�>Ê>?�&#��G������f[4�Ş?Ė@ˍ�?;<G��H�=47?�T�>j�O�R<ƾ�Z���r��C�q=�%�>L���av�P��BI,���8?�?���>D���.��En�=�敾�T�?<"�?�ɪ���^<a9�K�l�p=���U�<羭=�(&��S%���"�7�UǾ������;���ˆ>�@����>�7����c8Ͽ������;rr�PU?��>z�ʽ�F����j��~t�|F�"\H�'���:U�>��>.-��~���{�A^;�����m�>���%�>'�S����#�����3<Z��> ��>g׆>�Į��ڽ��Ǚ?փ���<ο�������	�X?d�?Sh�?�q?�U6<��v�z�{����/G?8�s?�'Z?��$��Q]�\8�m�j?����|`�{x4��E��vT>l�2?b�>��-��w=6`>h*�>¾>j�.�pKĿqȶ�|�����?Jr�?e�꾁��>\m�?�)+?�v�� �����ܳ*���z95A?f(3>�2��s!��1=�N`��84
?��/?C��DV��h?�����h��RIK�0/s;��>7�>�8�s��a{��G��/nX��x���u��}ۯ?� @w�?@�&�T,��%6?���>:4о'!���y�<<�>�~�=iʰ>�}�<����7�#P*�p�<�?g�@�2�>֙�#�����>6p?�̚>A��?݅�=�?ƀ=+ͻ�w䋽�d=�k�=�:,� ��>��C?z�?�5=�I|B��F��|R���o��b�GP�Ҿ�>�z�?Ŝ7?Rz>�0漫ъ=H��V��0�]��\!��>���,�=yn���q>9�>�b�=�qa�2����?@o���ؿj���i'��44?��>��?!��r�t�.��:_?y�>
7��+���$���B�X��?�F�?�?m�׾]f̼;�>��>PJ�>�ս�������b�7>ܝB?���D��p�o���>���?�@v֮?�i��E
?cx��ɷ���y���J���V��I,���2?�ݹ�Â�>���>4��=vr�����%�c�ٮ�>��?9r�?rA�>���?�����aE���1���V>��?V�?�9��񯾍[c=l�>�
��떿�Tξ9U�?2Q
@?U
@��H?��!п-(���/��tg��4\�=y�T��0�=�͈����;ćK=Sb>�6�=�2]>U~>��!>kfo>��+>l��=�hH=_o�����R���x��8I.��.@��m4�����W���Ͱ�(%���)�@٬��{	�׺4��I��G$���_���m8�[	g=Gx?2�k?�چ?���>?n����6>ž!^�<��k�u�>�k�>��O?.�?G�?�l�<�֪� �h�TƂ��a��2���G?T�T>G�>N��>�,�>uk�=F�>���>�S�> x{=�0]=�T�=d�1���>?"�>S	?��g>�;>�i>�ȴ�")��7h��w��0̽R��?�k���J��*��O������U�=<F.??�>����9п�ﭿ�3H?�����/�P�+���>p�0?�aW?�>?���RU�>����j��_>�/ �4�l�k�)��Q>i�?�;g>�'u>I3��F8��#Q��o��\|>	�6?�巾fe:�3�u��I�jGݾ�AM>㋾>�H^����{����^~��1j�?�z=&{:?�]?���gx���Ru�M���{�R>#�\>�=���=�fM>�'f��ɽ��H�D''=���=E�\>�?�,>�W�=տ�>�ՠ��Q����>�[L>VP>��;?��"?;U��������`+�+ei>�1�>�7�>�>g�N��ٲ=@�>�8`>�q�������<D��$^>�d�!�R�q�d���}=,6����=c�}='F
��A����<s�?�Y���3��)�<�����0W^?��*?O�{=T�:�F�*����P�޾��?�?@�G�?�����WI�|�?���?A���_�>[y.? L�>��M�P�ν�9?��'�B�
�����M��Y�?���?��=:�p��Cf��>�?8Sʾe�>�w��Z��Z��e�u�r�#=��>K7H?+T����O�h
>�1v
?:?[^򾏩��9�ȿX{v����>^�?:��?
�m��@���@�}�>j��?�bY?fqi>5e۾sPZ����>��@?R?�>�7��'�_�?l߶?��?X+I>���?�s?]`�>~x��\/��2�����]=9�\;Cw�>>F>[����gF�pԓ��g��۳j���Q b>�$=��>������=����Q��x�f��>kq>�I>i�>v� ?K�>ǒ�>^=�x���𴖾��K?���?-���2n��N�<Z��=)�^��&?�I4?!k[�}�Ͼ�ը>�\?k?�[?d�>=��P>��G迿7~��H��<��K>*4�>�H�>�$���FK>��Ծ�4D�cp�>�ϗ>�����?ھ�,��VS��GB�>�e!?���>�Ү=f� ?��#?�8k>v°>�xE��\����E�G�>�t�>�<?A~?ʕ?}亾��3�����T󡿲�Z��O>H*y?�l?Ȩ�>!��".��D5t��H��M���*�?��g?�K߽��?No�?�#??�AA?r f>����}ؾ�|��_%>��!?	�"�A�2M&����{?�N?I��>jh��=ֽ6wּ���#����?�&\?�;&?\���%a�7�¾��<]z"��_S����;�E�$�>�>w�����=�>u�=%Jm��@6�<<f<�H�=v�>���=�27��2E,?P�A�ꙃ��ݗ=g�r��aD��F>��M>�����^?�=��|���E����T�θ�?p[�?�m�?�Ա���h��)=?��?��?$Z�>�
��@P޾A��Qv��cw�!����>��>���ϓ徃���ᘪ�7,��Voǽ��I��>f��>��	?��><tI>���>�g���*��0��V��I�a���>�5�N�+����������3��ɽþ8~v��y�>�y��\~�>f�?��`>C�m>��>oi�:�>!�R>�y}>���>�H>�3(>2��=?�@;E3㽶�Y?�v��o!�ѡ�p�J�@?Y}�?�?MO��k��-�5����> ��?��?s��>�xM�d��,�?��?ϧf��
,?�X�=o~>�/�=r�������<#����qR>���<�I�h�e��y¾���>�?��X=q����Y��ƍ�{�=1�?�'2?P�(��OI�wr�lJh���I���D��:������!�ek��z��M��@��Ӝ��Qt=|H'?�b�?���dƾS�5i�1�E�i�<>!?$p>H��>� m>P�
�|?C���Y������x��>�1v?/�>��I?]<?A�P?Q^L?<�>,�>�k��zJ�>��<y4�>��>�9?�-?��/?�%?�H+?`�b>����A���v�ؾ��?{M?�T?l@?^�? υ�5�½����n�:x��k��=��<>�׽MDu�R�U=<uU>\?#J�?�8�������i>�U7?.W�>�>�>���Ji��n�<�e�>̎
?�8�>1���r��d���>R��?g���S=9$*>��=>F���=źtS�=ǂü���=7�}�U�8���!<���=���=-����{�Чt:��x;۫�<C�!?�~?�`�>�>>$z�F!�)��e
�=��'>���=�=�>�	Ծ%9��A�����e�;b�>JӦ?h��?.e�>���=' 1>ʦ���,�x��*1������?'�>{�P?�I�?�^?���>��>�˾�r���&��+����f=?�*?e�>k����Ⱦ�譿ܯ*�j?�+?JDq�2�K�/� �0�������>E ��Ɂ�������!�=�p=m���ӽč�?Nۖ?L�̼~�#�sMݾj"���-����A?���>?��>���>:�$���a�l^���=$�>�B(?^�>�O?�>{?�[?�cT>��8�Q.��nљ��@3���!>x@?گ�?/�?y?kp�>W�>|�)���/X�������mڂ�qW=#Z>���>�'�>!�>���=�ǽ�R���>��U�= �b>��>y��>��>s�w>��<�G?���>����"��򣣾�K��R5F��Zr?iϏ?��(?�i =���kF�֡��'�>@�?�3�?N�+?�9V��5�=t����Bir�R��>�q�>k�>i¢=P8F=� >�>�>���-�D8��[5���?�bF?�~�=T�����6��W��;S���?~ξ��������א�*ݽ~�ھ<�>�灾Ҙ�����vI,���þ��#�k�(�?Υ=%������`=P�>o�<?�">�˝=5�0>����<�*��ݧ�%3㼌���������<L��=�%>��¾.�?�|?@\?��0?y$�>�>X:>3�	?,Ը>? ?�[>�>�����_��Q��F������`��oQ��ݟ���=��Eց>y�>ثl>��;'��>'��=�-�<;<�=޷��� >�� >��<?��=m�h>�<�>c�x?�N��I���3�j�z���9J^?;�>�Q�=�|o�7�=?��=�q��S��a��O>�?Y�?R,�?�B�><<��>"���J&�h��=]�r<ݒ^>�!>��"�>��>l�=�����ٮ��ޞ�?q�@vC?
��K�ۿ��_>�6>�>bmR�^P1���]���b��!Z�F�!?�_;��̾��>:��=��޾X�ž;*=@�4>H�[=U����[�q��=�cw�:;=i=���>��E>�}�=�i�����=�8O=���=ܚN>����e<�fK4��;)=fJ�=�a>۱%>ϗ�>��?j�0?afd?F��>�Jn��Ͼ����\�>b�=H"�>�S�=x�A>/׷>��7?umD?̸K?���>D��=�3�>�`�>�,�*�m��8�x槾��<�|�?=Ȇ?q#�>�SF<=�@�0��(�>� �ƽ��?{�1?�~?F��>�T���࿿W&�5�.��i��A�H��+=�\r��5U����v�ߥ㽖��=�m�>.��>��>�Fy>��9>"�N>T �>�>���<�u�=N���O�<@甼b��=�����|�<�`ż����'�R�+��Ϧ�@N�;4��;�8^<��;�?�=a�>�	>21�>�6�=����c.>������L�lw�=�;���OB���c���}��.���8���@>TY>�ڀ������?�xZ>i�>>2��?��t?��>���վX����
d���S�lC�=��>�j>��d;��`���M���Ӿ���>hǎ>���>�T�>�:���.�)@�<�F־A�;�� �>o"V��/�t��h�R��ё�K*��g�r���=X�.?��y=#�y?P�^?��?�$�>����-#�V>>i3k��Qb=�'	�F�&�)z�E?A ?���>5��I�T�ƥ���3��Yq7>�I���d!�����1B���;�c���9�>�h��F%��t���t}����w0���~�ƣ>�T?�5�?��P�_�o��Mr��p!���3�1��>~�Y?�*�>�=?2>�>��0�SU��«��#>tq?��?���?�[>�u�=7O��%��>`�?}`�?�/�?�lu?/�D�o��>2�S<�E,>+t��n��=�U>��=c��=� ?��	?p�	?�9����	�+������5X��'=|R�=�K�>>8�>�Cq>�L�=�$r=��=�q_>2|�>72�>��`>�F�>�3�>:w��/9�9�&?*��=�d�>ő1?�΀>nFC=윲�_��<HD�>D���+��!�����K�<;�*�S=m�μ�K�>F�ƿ�0�?�X>��?T��P�J�^X>T�V>Əٽf��>��C>�cv>�D�>�T�>�>�y�>U�(>��Ӿ!�>���� ���=��jN�bӾ�!w>������b��J����D�Z2��l����g��T��u=���<�y�?/�')j�iZ,�@���?+S�>��4?Ŋ���,�c�>pu�>+�>����ȓ�j���_�ܾ�C�?	!�?�C�>���>�T?��?��c�r�e�.�b��E������w|��D��Ì�\����06���]�ǦK?���?��S?5��;ȑ�>	De?�/�T���>�6��9�`��=�y>�9��H8���J��5�о��y��4l�5Ō?G��?�K0?�N���3��X1>%h/?bY1?k?�3f?�_�?��<��<,?���>�DC?h�?�. ?��?Z�?ƺ%>�u	=80�<��=�jμĉ�����ͽ�-W=��M=ӓ=p��m��x�x��]���~=�?R=��=��=p�b=#�<	Y"=u>/>(˨>\�\?�R�>y��>6?�]�8�7��o��\�-?��=;��ॏ�����{��mq�=Y�l?��?��[?|_>�<�F��>���>Cs#>�EY>�r�>5ٽt.D����=��>�>>;۠=K�B�����K��W���o�<�>#\?��->�ṽ��>i>��b��NeJ>O�����5��վ��N��A]��j]����>U?�i?V��=�iK�E�>��X�+�N?�[D?~�"?8�X?������	�\�7���ý˪�>H��dv/�'L���#���@�z��G'�>����s���Gb>��	}޾cin�;J�~���OL=�v�HW=�3�վ�9�d_�=��	>p���� �����̪�u&J?��k=�J��!�U������x>H��>3��>�:�vv��}@�㋬��Ɩ=V��>;>�˙�����iG��.��S�>��Y?�NR?�~?ukc��au��N/���)����齙,??ۮ>�
?>�>m.=ז�w�s�i�+JZ�ܩ�>ɠ?Xj����f��5̾龌�	�Ä�=S��>{�C>�'?%�`?J/?9�R?O?0?�P?�j>�6=�t۾A&? ��?\�=��Խu�T�s 9�6F����>9�)?d�B����>J�?��?��&?@�Q?M�?��>�� �kF@�撕>Y�>��W�fb����_>ҭJ?���>�;Y?�ԃ?x�=>`�5�u袾�ҩ�cS�=�>��2?c6#?�?z��>̈�>������=���>��b?�2�?~�o?3�=��?�12>���>}ۗ=8��>���>��?wCO?߭s?K�J?��>��<��������z�s�z�T���;��J<&Hy=�-���s��f�̀�<4�;����ɀ�:��|D��������;���>��k>�X��p�,>#�ʾ(����E>�?I�,�����t�=����=���>�1?�Ԙ>J �a�=��>"��>�R��)?��?^�?w{-;�sb��ݾ��R�,a�>��B?.}�=��k��[��Ovv�� :=|�m?�*_?J�[��M��\�b?�^?�D�1�<�D�þ_c��g��O?M�
?�4H���>]�~?{�q?-o�>`9f��Kn�}���Fb�O�k��a�=<��>2�6�d�C0�>��7?:T�>�b>���=x[۾��w�@H���?��?���?���?�*>��n��+�?�2��I_?�%�>����M"?&�0��޾�㓾e�����Ѿ7D��R쨾V���S��bDU�w5���lٽ��>5^?�f?�l?�>h?:s쾟MX�w^�!w�+�Q�8 �$��Q<���L�~�@�\�l�	��־����-=c�{���@�B6�?O(?�3�J��>����.'�Hξ��=>������_�=Im��7�+=�k0=��l�\�-�����?Gc�>��>_z>?�eY��<�,�1���6������q0>/q�>�F�>	V�>�d�s�1�q�Rbľ6���1Խ�Hw>fd?��H?�7o?�W��0��ǁ�FH�nB��諾5�B>�>y`�>xQ_�d7'���'�ͨ=��q�
������N�
b�=�p1?��>��>c�?��?/��ޞ���X}���3�λ�<�0�>�9i?���>.z�>�F⽟�"����>��u?�>O��>�3����)��R��%���?A�{>{?�h�>w���Ub��-���5��A�� >B�K?-˾Թ�Ћ�>�h)?m�>�x4=.�T>")>o� �'B�vT߾uT=�� ?� �=�F>.���]*�۸��A��O)?1K?p蒾�*��3~>�$"?��>U-�>1�??*�>=pþHeD�t�?��^?�AJ?2TA?J�>��=����`<Ƚ��&��,=݇�>	�Z>@ m=,��=���~r\�8w�<�D=�v�=��μ�P����<d���G�J<���<A�3>zտ~I���Ӿ���Tؾ�����S����Ð�T�w�2ľ7/��y��������,�7��pm�$ښ�2�C����?&b�?�U��鮓��+��孄�S�`�>��N�J����B<J�Vy��{�(������2D�ISZ���U�P�'?�����ǿ򰡿�:ܾ5! ?�A ?8�y?��7�"���8�� >sC�<�,����뾭����ο?�����^?���>��/��p��>ޥ�>�X>�Hq>����螾o1�<��?6�-?��>r�1�ɿc���k¤<���?0�@�}A?Q�(�9�쾋$V=���>ʏ	?!�?>�]1��G������Q�>�:�?���?�eM=��W���	���e?��<W�F���ݻN�=v'�="=O��4�J>�V�>~��PA��;ܽ~�4>�݅>��"�z��&~^�cW�<"�]>v�ս�6���҄?q�\�@�e���/�����Y�>]IU?���>�٩=Y)+?!tH�cZϿ��[�"-a?��?�`�?�(?fν���>݋ܾe�N?O6?z�>��%�o�t�g��=bU��LXྠ�U��q�=���>8�>�A3�M�� �J�����(�=�� ��ĿA#�}����.=Pּ����	뽎
½�˼�����X� R��k=�o�=�-W>�p�>�C>�_>�Y?��j?"(�>�]>�۽����OԾ*�<�|�����ݒ��X8�6O��yx�W޾���C��������t<����=�rP��������me�}H��0.?��>	B¾��N��3p<�m̾�R��7����+����̾t�1���i�1�?CB?\���:�W�7u�dRD��ݽY?m���<�������=TF�>�<��>�=�Hݾ��.���P�pP0?��?/���Ғ�i >G����=L,?���>Cj<�ب>�!?.z'�����]Z>��.>ԣ�>`�>D>�T����ݽ��?N�S?d ���A���)�>,Ӿ�r�v��wV=�>h�0�����."X>�m<����ϥ��c�����<��W?��>��)��o���k=�B1=^�r?$?�t�>��m?��B?4[{<�j��^U�p �Mp�=�iX?�Ai?94 >�,=�o,˾Ks��F5?qb?HL>6t�k�8v0�N~�x�?zn?m�?��żu�~�i锿��
��M5? w?�`]�g�����EV��0�>���>�S�>�{8���>56=?/Z!�����*����3�Ъ�?��@&h�?=��;á����=�?���>s�M�{�Ⱦ����ۮ���v=���>I`���t������1� G6?;��?�O�>Ϊ��1����=ە�Y�?��?������i<����l��x����<��=T���"���� �7��Ǿ9�
�ۤ��"̽�2��>�S@���;�>_58��-⿻MϿ�	��Vbо�]q���?ʀ�>+ɽH�����j��<u���G�<�H��������>I�M=�5(���ɾ��y��U�
�U5?��O=��p>���"q˾Vؾ�?6�}+�>s�?��>�߁9�����?ޟ!���ٿ�������?�h�?��`??� �6�Y���� N�NQ?ሓ?(w?
�=��8c��j?�Z��0P`��4��JE��U> 3?0G�>��-�э|=�>/{�>i>r!/�t�Ŀ�׶��������?4��?�q����>ၝ? q+?�e��4��3`��}�*���(��8A?� 2>M���Ƴ!�:/=��Ԓ�-�
?gw0?M���,���l?^)��,ڐ���S���c�İ�>9&��M�l�_�0���Rj����ޠK�U�?(�@�-�?���&D�UO9?�µ>`$��GZ��A_e���>���>>��s�Vj���5�y�۾�j
>^��?37@�?�˛��A��MŅ>�g?a�>P��?:��=�?�G>)Q;�6��R�,>
�>�nU�[�>hp<?cI�>:�;p.��,EO��MH��S�pS)�'�8�J��>ˠa?��?I(>���|y=�h&�*�5��#�Y/����N��ɝ�w�ź��>�0>1��=���0�����?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji�}�?M5�@���gV���r�O�UI�=��;?+���y>G�>��=çw��é���q�Yӹ>'�?���?�<�>�p?q�q�,�G��[�<n��>�o?�?��λS쾽�,>��?X|� ō�U��zj?��
@��@��_?�.�������g���c������!�g>T�s>��=��#DZ��>����b�~�r�=}>q@>M��=�A>�c�=(��=Z�}��3������������x#�j?Q�DP8�nB$����NK?�� �U/��E$�%nb����5�6��0���]@�=�<?�O?�??�>x�x�(a>R���>���A%�=.��>%�-?�M?��?.o��{ز�ʗl�za��1ذ��i���	�>3�>>� �>6?�>?�=��>��>��>�=<f@=wB�<��</��>��>�d?X$?�C<>��>Fϴ��1��k�h��
w�u̽1�?����R�J��1���9��Ԧ���h�=Gb.?|>���?пf����2H?&���z)��+���>|�0?�cW?�> ��w�T�5:>6����j�5`>�+ �}l���)��%Q>wl?k�f>H�t>�3�\f8�*�P��{���<|>�,6?b�;?9�#�u�f�H�Uݾ%GM>j��>IE��i�������oi��${=�r:?
�?���۰�C�u��G���UR>�\>;'=ӫ=koM>�Oc��ƽ~H�@#.=9��=J�^>�?W->剣=,��>n?��f�R�"[�>SKK>��>P:?$$!?86x�;���<����+�~ f>f��>��>�\">�)S���=���>��g>ʼ��V�,b��cH��\>t���KD���G��T�=�=����=0Y=}���K��
=LQ�?]���闇�*�0���G��,(?�?��>��ľVRa�E���A��#&�?i�@-y�?�8�#|^���O?N��?�o��4>��?C$�>��پ�C �px?F�<�����O ��H��9ӂ?#^�?�V�=p�f�^瀿,o=@�K?	m��Ph�>{x��Z�������u�v�#=R��>�8H?�V����O�f>��v
?�?�^�੤���ȿ5|v����>X�?���?h�m��A���@����>;��?�gY?roi>�g۾<`Z����>һ@?�R?�>�9���'���?�޶?֯�?��E>Pԕ?=�m?'�>NWq���2�	����Ȍ�	��=R�����>_�!>����B�����t?��jym�Ћ�Ʋ>MA=���>^=��~�ݾO�l=�%�3X���Ľ\׹>�O�>��7>���>	L�>W��>C��>&�={�k�F�������R�K?���?��+n�Q�<sJ�=Ӏ^��?fH4?4^�T�Ͼu�>�\?W��?0�Z?�;�>���A��~���Z�<>�K>(	�>�G�>�%���_K>��Ծf�C����>[ė>}ߤ�6)ھg$���꡻YW�>!m!?���>�a�=[� ?µ#?��i>7{�>=tE�j1����E����>���>b?_	?b?mӹ��i3�B��Y⡿�O[�x�N>o�x?`?Q�>e_��s���T7�G�J�ᒽ�j�?�\g?��ơ?�+�?/�??E�A?ݐe>���G�ؾ�ʰ����>|�!?��A��M&���s~?�P?���>s8����ս�Dּ���U����?�(\?;A&?���,a�<�¾U8�<��"���U��;(�D�T�>��>�������=�>�װ=Om�{F6���f<�i�=��>��=1.7�u��<�3?tn�<�	���/>�v���B���X>8O'>?R��!f?�Xy�sa��Ȧ�G̝��8�����?!��?�˗?j�2�r�`�t4L?�?^$?f��>�ũ��mԾ�����Z���H����	&>c�>J,E=h���r��|�ϗ�����%��>���>l�?SQ�>��Y>窚>�g����'�^�������c�F��p2���+��!�諾����e=�g����~�g|�>I��;n&�>?X	?�c3>��Y>�Q�>�X{��ۗ>p�S>�pE>s��>��)>��>��
>>�t;6�ڽ�_?���.+��h�s
$��Y!?��}?:�I?��	��e�����Ս>���?H��?�?
H���7��3?�
?@y��6	?̸�<v�>�3���\�T	?��U�� ��>謺>P:��r�"����'�?/�> �3?t�>0���򊽢v���z=w�?J�%?ki!�AN��ir���R���Q��F��ZKm�뚣���$�7�g��"��S���B����%���=�-?�̅?����޾z᩾@�l��&F���>9E�>1Ł>qv�>�*>�I�	�2���V�t6�|�J�ng�>$2p?CO�>�I?��<?�wP?N�L?���>��>�!��Y��>,�<�q�>v��>�9?�G-?ӧ/?��?��*?�a>����:����uپ��?��?�?0�?ؠ?�����[ǽ�U����\�ksv�����H�=)�<�zԽa�u�t�S=%�T>K?����8������j>��7?���>��>���\+��:G�<(�>�
?�V�>�����lr�!d��8�>���?a��7�=+ *>)E�=����P�����=b�¼ɐ=�����B;�%� <�q�=:��=_�}�[����k�:H�;�˯<G"?�T?d�
=o�>ᯠ�|{�aP��>�`�>?��>2C�>���8�0U���]�Қ�>�}�?��?�`�<��=J��>%B<������4����,�m����>r"?�_?*Ѧ?��.?+�4?�>��9�7E���\��b���A�-?4�+?���>8	�;�;W��ni2�v�?U?c��_�,7(�l�̾�ƽ7L>
�+�:6|�༭���<�q�<���e4����?X\�?E��1�U�7��N�����>?�	�>�!�>���>X�(���f� ���#>�	�>ǑM?���>	9P?�{?M[?O�S>@�8�񭿩ؙ�	�*��� >��??,��?�؎?��x?��>f>h�*���@2��O��hi�E��+aR=�Z>�8�>�&�>[��>��=�FĽDc��ަ>��^�=�"b>[g�>���>�G�>��w>L��<
�_?_��>��6���'@������ܒ�w?��o?��>�s~��s�L���z�_u�>�:�?���?lTY?)پa��=��;>l�Qz��>�'�=H��>tF�>œ�=^��>Y��>�j�>��L��~(�A��+�J�V�
?(�>?+�>�KĿX%Q��悾��▐>��j���#�A�h�>˾��>��<A�-t�6Ջ�d�;q�s�䘧���2�@���� �>��e=a2=d>�{��y����Zw@=�y�=k�=�VA�V"w>��_<aM�<Tڼ@��=�ɋ�T�;�ܱ(>v�Ӿ�˕?�ˆ?6%?�pM?#��>���>���l�?䎩>��C?�e�>714>V6���1R���^����D���B���Ͼخ�>�Ѕ>���>���>y8a>��=p��̣�<��>`�=�=R��=-z>ǘ�=�Ԍ=�>�
�>�Lx?l��^���*�\���=��O&?�Mw>��>���!c,?�>�=����D��[��!��?���?,(�?��?*FG�y�> Ҿm�G���-=����(`�>�d>�^��J�>i�=���R���ޅ���?��	@�	F?�G����˿b�h>�:7>-�>6�R���1��\�D�b��Z��v!?X;;�1̾ �>#F�=O߾vpƾ`�-=`�6><�b=���lV\�x�=�L{�v�:=�*m=3�>M|C>�P�=j���%�=V�I=��=��P>Վ����7��+�%�3=���=��b>��&>���>>�? �.?d?�׸>�:l��оe�ž���>^��=[��>��z=3:>[,�>0I7?I�F?��M?���>|xi=ǃ�>�!�>��.��n�h=��%��`��<~�?E�?�N�>J]I<�U9���q�=�����F?631?S�?jb�>���2�&��S.�9H�������=�et���V�\�����׽��=�`�>e��>��>&�v>a�5>N>,��>O�>a8�<a3�=�i�U��<���J��=Mۖ��9=�7ļ-��:�V.��l/�5!��j��;���;�hm<�g><a��=_��>�l>)w�>_@=Qq��5&(>�ǉ�8�L�P-�=S��qD��F]�i�y�,���B�n"6>V�c>�]��+��G��>,�q>N�?>+��?яr?�	>u��|о�1����I���H�� �=N��=�oB�P�=�ӣa���N�9CҾ @�>���>鴲>�Q>�5���3��Q�<u{վ4�1�F�>M}�O#�����*)`�d�����h�r�~<��N?w �����<Ӭu?zc?f\�?\}�>w���)��kI>"z��j�=,t����̡�F?�?��>8D���@�R��������ĝ>�D��1�/��!��:cV��p>?���/�>��澧R���2A���|�����#���[�9��>vS?'�?�?���|���^�%�0��}�0E�>��n?8�>�̋>^��>{�~�#���m����>�$f?��?��?�S)=<9E=�ȁ���>v)?�S�?��?<\s?��w����>��9Ʋ�>iG��$�=�=,>�>�=��=�K�>��>`��>�劼,��o���m���x�[�M<�1C=�9�>��y>��`>�Ϡ=nu>�}�=��c>���>=�>�5> ,�>���>L����
�0�&?o��=Ť�>4�1?i<�>��9=c����Z�<�1"��?���&��U�����:�<$B.��48=y��!"�>W�ƿU۔?L�[>���@�?�����Z.�{mP>/ S>v
׽�>�/@>�tz>��>�Ѣ>��>�W�>�i(>�GӾ�d>'��]b!�C�i�R�7�Ѿ�z>������%�@��L���XI�Ik��h���i��+��9==��Ҿ<�I�?;k����k�b�)������}?},�>A6?.Ì��<���>���>ۦ�> V������Í�Sᾃ�?���?l�>��_>,-I?��7?�9z�T�*�ڐ^�ϩ��93��sg�>U0�⇿Ҁ�m�����Bk?��?!�F?ޅ�d��>�aO?8�\����� ~�>?:����%�Ƚ���>��\�.}Ҿ4�g�
�Ⱦ���Ƞ�>l�?���?��&?f)�M�e�]81>?�J?e�V?@q??w-�?�pk����>��g>�X?NR?K�*?�#?��>��)>�j��Iz��6>}��<U���ѽ~Lս�^�Q�<�$�=Ҵ�̊���UU�1��O�<� &<f!�:/:��#=]u\<(A>�`�=�*�>%e]?���>���>k�7?����n8�A���/?U7=[΂�����p��:&�$>'*k?"�?-�Z?a�b>{|A���B���>�ɉ>�I&>i[>���>�,�%E�E8�=�w>�P>T��=��O�<����	�U4��f��<��>=o?��(>�����b=G`�緘�My>R�z �������
H�s\�N^���>o�>?wp?�9=� U�:ms>/�R��	a?@�X?�<?8c�?u�=�->���>���n��^=�:�>eD4�ܧ �{���I'����B�Q
=E��=����g��;)a>�^��ݾ[m�b�J�v��V=��0�[=���@վZ�}�я�=�8	>�y���!�����,c����J?ncj=���W��q��2�>�J�>�0�>��;��X|��@�[������=��>��9>����qk�p�F�yP���T>�a?~8V?�J�?ʫ7�SCu�%m�����e�9��ϵ?v�4?h�#?M��+n�<�׾H�!�� ����N��>- �>����+2J�̾4����f�O�q>�U
?|k�>��U?��"?p9&?�a}?3H�>��?��>_c�h����%?��?ڈ=xѽ�HT�%�8�Q�F����>�)?'A�[��>Ѧ?s\?;�&?-Q?�]?	x>#�F�@��,�>�'�>�xW�'/���=a>>�J?��>�Y?tك?�\A>�e5�Fe������zz�=��>@�2?�d#?�%?��>B��>59��~�x=`q�>��b?��?�o?9�=y�?��/>�T�>G��=�c�>u��>��?~�O?�t?�]K?���>r�<j����D��Ўx�i�6����;��\<MM�=I��o�s�cC
����<�lm;�ȼ�
����L/A�;�?��  <%q�>f�p>ە�&�/>5�ƾ�⇾�eE>]�������ꋾ��<�α= $�>��?h�>Ϧ�J��=�>&'�>�j�q�)??ã?�3�;7�b��3޾(�O�%��>�^B?� �=;�l�H��W1v���U=7�m?e�^?��W�R2��@�b?�]?$h��=��þ��b�ˉ�O�O?-�
?6�G��>��~?^�q?��>$�e�5:n�&��
Db���j��ж=Yr�>FX�.�d��?�>Y�7?�N�>v�b>�%�=zu۾"�w��q��r?u�?�?���?�**>}�n�U4�E.�V󍿨e?�G�>�*����"?ػ4�;ܿ��ٛ��Ҡ�<�׾T���*���ˑ�H ��c;�ku��{�ӽ���=π?�/u?��^?��]?�]��-Q[�� \��ڄ���X�0���~�
�g�=��ZG�ޞ?�J�s�a�_Ͼ
ى�=�i�9�3��]�?F`?w9���p�>����kW��(���<L���Kg_��Q�=�^��%��=m��޲��-�*�r�����?�V�>���>��B?�X� <+�,.%���@�����*>\w�>��>	�>`I �ܓ������r�{� �|��y��c>Cj?�bB?Mt?�uٽ�4�gG~����K6����qH>�S^>�}�>�����"���*���>�5dv��!������'�t=E�7?!�>|��>膒?m�?��I���z���X#�y�=��>�i?��>�>�>��ѽ^�&���>��t?�>��y>�zپE|�&,i�p��DIo>8(�>s*?��,>-�k��pH��j�����d
*���>e}?����y��_Z�>��0?���8��<߲�>�!�=%�n���� �G��>Q�?i
�W)q>�c�Đ)��叿�����O)?'J?�Ⓘp�*�73~>7%"?�|�>�(�>1-�?� �>omþQ���?�^?�AJ?�RA?�K�>�=����5ȽT�&���,=8��>8�Z>$m=ې�=x���`\�f}��E=쎺=��μ�X����<r��*K<Q��<� 4>eۿ�J���پ�����r:�X���@������2,�w����/���v��l�a�*�N�U���d��ڌ���l��r�?I��?�2��nf���ٚ��t��e%���ͽ>�q�li��������
�Y����<�~���X!� kO�YRh�w�d�O�'?�����ǿ񰡿�:ܾ1! ?�A ?8�y?��6�"���8�� >�C�<�,����뾭����οA�����^?���>��/��l��>ץ�>�X>�Hq>����螾d1�<��?5�-?��>ˎr�0�ɿb����¤<���?0�@�A?��(����N�V=���>}�	?[�?>��1��S������>�(�?�ʊ?$�K=��W����+�e?˿<�F���ܻUy�=T�=J�=����CJ>lN�>����@�<�۽� 5>���>�"��0�.�^��ֽ<|e]>9�ӽ�E��nՄ?�z\�If�̡/��U���[>��T?�*�>�,�=�,?�7H�%|Ͽ�\�.a?�0�?��?��(?pٿ���>��ܾ��M?E6?;��>Y]&�o�t��;�=r����!��V����=Ӗ�>Yp>�,���utO�.]��O��=�����ſ1{%�� �N;=2i;��\���𞔽?2�Kz��:xr��G�]T=���=b�P>d��>{�S>��V>7�V?�j?1��>�S>U)ڽ�ŋ���̾#�E�%<���������颾}~��uݾ�-�4��&�(u˾�<����=��P�%d��BM���f�x�E��/?Ÿ$>��¾�O��e�<��ľ�J��]3�����A+Ͼ!�0�L�k����?��>?����F	X��\�3,���̽��U?����મ�+C�=҇O��4�<xʘ>ތ�=��޾�b/�a�M��}0?�_?����,H��8T*>4� ���=�+?Xn?63W<�Q�>%H%?[}+�Y��::[>f 4>�/�>�#�>��>	��x۽_�?�xT?���_��fА>eF���sz��Zb=32>:�4�����7[>1?�<����gXW�����{��<.)W? ��>��)����e���Y��==�x?��?�=�>�|k?t�B?*��<yh����S�%$�ߺw=,�W?�.i?&�>tB����Ͼ����s�5?��e?��N>�ih�����.��L��?	�n?�c?����}�O �����lu6?$w?0�X�Py�� l���J����>���>���>�7:��׬>�h@?�z��b�����}�2���?��@��?8:2�����~�=�� ?���>�P���Ⱦֻ�����Ά=ފ�>�У�ϙp�г�}q9��]2?0<�?ѯ�>^�t�5����=ĕ��`�?��?�ª�gvm<D��}�k�}���E
�<!�=����"�m���7��
Ǿ	�
����!j����>�Q@�U�m3�>��7���ABϿh.��.�о&�p�`�?Er�>�ʽ옣���j��u��CG�p�H��ƌ��k�>m>�y��k��5�{��s;�'`��>��>�%���>�S�C��趟���0<��>��>���>�����Ƚ��Ù?����>6οӟ�������X?�_�?7l�?hr?I4<&�v�N�{��#��,G?5�s?�@Z?�^%��]��6��j?�^��;U`���4�HE�U>�"3?�A�>L�-�ٶ|=�>��>
f>�#/�w�Ŀ�ٶ�����I��?���?�o�P��>f��?s+?�i��7���[��f�*���,��<A?2>����!��/=�7Ғ���
?�}0?I}�.�3 q?^���y�id$������^�>ݫ��@��<�,�=�k�,u`�iNn���[�{!�?�k@���?$ĉ�i�1�p:E?�(�>�����y��?>8�>?^�>xޱ>���=�ȃ>T!$��)E�i��>��?��?�),?|��d����_;>6eV?D=�>�T�?�N�=r2?�}>Sʾ�d9!>���=?�Ľ��>�~]?���>�(
966��2�j�H��`U��e� �>�d�|>�z]?m�P?�b�>n�νj/��7��19�iB7�~Ⱦ�������<s�꽂�S>��a>|/	>�Z��l���?Np��ؿ�i��Ir'�)44?/��>��?����t����k;_?�y�>67��+���%��]A�*��?gG�?��?3�׾)`̼�>��>�J�>��Խ����
���E�7>w�B?"��D����o�L�>���?�@�ծ?�i��.?F���Ň���x�1��+���4�l=��+?X�ؾ���>*M�>W0=�o�����vh�&m�>��?q��?��>đw?�h��K!G�=��V�|>�(�?�?[���W�վT�	>��?Γ�t������}?�O@f�
@Z�J?~����Mÿ�j��^K߾����$�=�>�m?>�'�r�->��4>>U=����|��=�~A>�uU=e�9><y9>�=�=,t�>�qx����橱� ,��<-7�A1¾(����<��K�ฤ�$�=�Q��"�ݩ���v�0�w�W�9��D �Ͷ<=I��=��g?�]?G�n?�?��<�8�=��뾄f->_=�V>Q>d�S?�A?��
?��`<K�m��F[��ʊ������l�j��>_>n��>Q��>��
?����VK>�P{>�Ec>i=��w��������!>s�>��	?��>gC<>��>>ϴ��1��S�h�zw��̽-�?n���9�J��1���9������
i�=2b.?�{>���?пZ����2H?1���~)�;�+���>a�0?�cW?�>����T�3:>-����j��_>�+ ��l���)��%Q>~l?w,f>�{t>�2��O8�,�P��̯�E!|>�N6?�S����:�x�u���H��
ݾ:M>��>�S������G�~�i���x=8;:?��?�϶������t�q睾u�R>`�Z>�I=�ޭ=r+M>iVf�ôȽi�G���/=���=�:_>>j?(,,>O,�=�ǣ>0)���O��P�>eA>�"+>��??�'%?����虽����v�-�Zqw>7��>���>Y�>[J��*�=�:�>��a>[v��都�q�?�H�W>�}�H�^�8�s���x=�s����=x��=� �j�<���'=<��?N����^��zž���/'4?<�H?L?�K=�me�>���)����?|B@���?����Vcq��C?n:�?�)�|
�=�S�>���=|$��L��9?Q��N��^'!��J�3�L?M�?�[>ʒm���m��:>��-?㆙�?g�>5y�Z��#����u��x#=:��>�8H?�T����O�>��v
??�]�^���A�ȿd{v����>G�?P��?�m�"A���@�Zz�>���?�eY?ji>�f۾�_Z�T��>r�@?�R?��>09�ҏ'� �?�޶?���?�.2>��?}�h?��>v|�	`5�t���������x=�z&�,�>}p>�����R��Ɍ�l�����k��i!�^g<>�7=֫>L�G�y�����=߮P�pž����>S>�>
ST>zY�>�t? �>�U�>1Ff=�{����k�����K?���?���V1n�yZ�<��=��^�U&?J4?�[��Ͼ�ը>�\?6?�[?�b�>���A>���迿�}����<|�K>3�>�I�>���vNK>��Ծ32D�s�>ϗ>�#���?ھ�,���m��jA�>�e!?��>�Ӯ=�� ?3�#?��j>� �>eE�6��v�E���>���>JK?��~?Y�?`ع�X3��	��-롿q�[�|>N>��x?�G?[ӕ>܈��~��[F�l<I��璽⛂?�hg?��彵�?�1�?��??��A?P6f>���dؾ�+����>��!?�"���A�5L&�@�2�?�O?���>�i���?ֽ]�ּ9���v��L�?+\?�:&?����"a�@�¾3O�<^i#�;�U�<�{F���>۝>7s�����=��>�ٰ=�,m�k<6�a9f<�B�=}�>��=97�E����,?����tރ����=�q�`D���y>X�:>\3��E�^?��2� �y������؛�QC_���?���?;ǖ?x�����g���<?A�?��?���>4®���߾ɛ�)�x���o�ɢ��y�=ͫ�>�E��Aa��饿i���1���ԥ������,�>�I?>��>�
�>�4m>Ra>�0G��K��Q��d�ﾰo��i�	�����.�z9'�T�̾��G�8�Ľ�Ծ�Cn��>�8�=P�>��!?�I�>���>�?��Y�b!>>��>���>��>\<�>���=a/�;�̽��k��<\?����� �f���)��=?�?��!?+���
���2�j��>^@�?G��?ͽ	?mK.��2���?\�-?O�B���:?Q�=�]#=Ͱ�<��~����aŽ���>5lӽfh>�`�G�4���G�>%,?(7 >}߾��ڼ�s���n=�W�?��(?�)�q�Q�âo��W�X!S�h3��h�����q�$��~p�׏�P[��@��3�(��*=B�*?��?¥�vQ���k�_?��/e>p��>@2�>���>	wI>�	�±1�^�D('�a3���\�>&0{?ڠB>#�`?j]?l?2�O?2$�>���>v}Ǿ{?�>��>&��>��Q?l+*?��?-��>��?�>>	���2� ��:���3?�c#?	�?*�>� ?�Ɍ�cF8�|���i+=n�+�~�%����=:�=
���ى���=	_?�X?�����8������k>h�7?��>���>���f-����<F�>�
?�F�># �~r�c��V�>���?b����=��)>���=I�����Һ;Z�=����&�=�6���y;��i<���=���=abt�;���G�:���;�o�<}7?NJ(?���=ee�>u�7��Zݾ(羰�2�z�=��>�=�>�	u��1���S��Ipl�hb�>4C�?~&�?��e=��`=�[!>{x"�@N� �z+ ��;��^X>Q�?�eo?��]?���>-?�|S>[3��:��.3���	���Q?� ,?W��>%����ʾ����3���?�[?�<a�R��k;)���¾�Խ>�>�Z/�=/~�����D��I��������?῝?�#A���6�Dx辍���V[��ϓC?l"�>�Y�>��>8�)���g�%�~2;>���>>R?p�>��f?�+�?` _?�,>�#��E�� ���9>D)g>K�Y?\�?��?,�a?gb�>�V�=��8��u"��01��_�*Ľ��D��u���Ȓ>3��>^2?n�>�#�>T�S>�}Խ3辧`
>�I�>[��>m��>�i�>���>�M���Q?�8�>�]Ҿ�O뾾�W�:h	��$��3?�kb?0�?JD>���a�9n�F�>3��?��?�J?8������=U�
=�c���Pz��)�>ԛ>vߘ>�'V>�(�=�>���>�_�>:�2��W�N�3�l01�`? 9f?�l�=ъ���3���˾���:B�>����z(��t�=z��>$�>v�
�c��m�;/�O�~g��!�Z��gt������7ƾ0��>}A�=�8�=�pq>�u�=�s˾�A��_;�<Bѽ�X��%?�lx�=1n=t"�=�~�< ؋��P�m�E9 � �<6Ծ�Hz?DI?98.?�G?�h>��>�r��,�>���1$?�]>Svڼf豾ӞG��@�������^پ+�۾%h������">뤼�:>�k.>�I>�}<��=��e=F��=ou����=�|�=���='�=��=�>��2>|?�؅�T����U�r+��'.?Wg>p�>py����+?D�>]r��|���1��;y?�l�?	��?d_�>������>������Lg=O5= �?�G">{�Ҽ��>�%=*��F��/5���?��@�Im?=���Iӿ3w>f A>�	>^HR���.��RT�F�W��Y�|�?	<���;���>/˵=-��G�ƾ�"1=�B>S�=#��H\�^ѝ=��i���.=n\=���>??>J'�=HU��}��=(<Q=S��=�eU>R��uO�R�<��5=�g�=ܱn>L'>`0�>��?ZQ?�]?)ݸ>�q9� U˾Gg�F><�=�;�>>�=��="ج>��1?�YK?k?_?���>ӣ�<��>3��>4�*���g��#ʾ�
���uI=�?��?O\�>ez=}M����`�2�"���A?ȷ-?hV?�٪>�
���߿�&�.�a���w��;B�&=m�p�+�D9�����ź�%��=�b�>b��>�1�>��w>A�5>��I>���>*�>a�<Uu�=�	m;�5�<(�����s=Ȇ¼��<�����:������.���Ѕ�;��9;W<��W;09	>���>�'�>Ua>��T=�)��m��=TU����h���=n����\W���a���p�7��OhW�_�">�>�_Ľ/n��oN?��>�=
>%o�?�x?d�=���1���8���)��j�AR>�>'��N�H��h��u4�(�ھ�8�>r.�>L�>���>��*�~!>���.=4Z��43�p6�>�G"�{��=KC�,0}�/���ʶ��K�f��汽U@?�ڈ�Xo>��J?�j?�ܙ?��c>���j��o>��⾰{b�{���(�ǽ�a��'8?g�8?,�>���BuX�������>P�o�>�R�%礿��4���"=𪣾��><G���UF�����-��ےJ��S���>d�L?ǻ�?�K����}��I��@*��\-; ��>S�=?�Ñ>���>�1?@?A��r�;U��:�>�p?��?��?<05>���=����g�>#C?�w�?e��?��s?�C�(��>P�9<�*>�ܒ�x�=Z>�U�=]�=�?tw	?��?I�����
����?�ﾋ\����<H�=4��>M�>z�j>� �=4}{=�S�=q�\>c�>�/�>y�`>?��>cߋ>���������2?W�=�Z�>3?B�w>���=�W��J+�NT���v�?��V�����[�������e��sy=�����>RN¿b,�?���>��Ɩ?d-پ�5���n>�F>��ν���>� J>l�T>�>�{�>��>��K>��A>��˾BU�=g4����~�)�f�s�
u⾞ �>fჾ[|�� � �� f���н�|����[�c�V�|���2��H�<���?:v:���g��l5�lU��\�>��{>�� ?c�������R >�>2p>m����������pɟ��R�?�1�?�S�>�&�>�6?�6?+�L��-=9G��u�����Ćc��k!��k���`~�����w�ͽR�??߬�?�1:?;�,����>�r?�Q��c�,�	�>!���������>���f �*���5��:�_�5>L�?cI�?�R?���U؋>��o?Լ`?%�s? -??��[?�X�k~?��>|-E?'�?��L?�y8?:^�>9s�=��;=�;���]>��ٽٻ�H�Ľ�g	��Լ�����
>+��/�������&6>E�>(X:=Ss�=}�:=���[59���<��2=^��>��Z??�>j7�>m�6?�絽��)��2þ�>?��s�N����p���ؾ������=Jgq?�?*\w?;�>��1��{�>|>X�>_�$>��>Jxr��z
�v�=Z�'>b�E>Ş=�g�����t�����o.�=��>��?Z�>H��û9��r\��̓>1L;�`������C�2�N�ᮅ���>�j\?��.?���=Q\��^ֳ=��[�x(\?:r?���>�5�?Xo0�@�D�k�:�G���M_�=���>U�"�u�P��v��᯿��;�o�_=��>�����q>�L��X�#�t��u`�4����B�5�9��=��� J��1�m��=4>^T�=�z��K��Ӓ��b��A�3?�v6�;����c+�|��숃=D�">$%�>���=z� ��M/�x���3H=���>��>|��]M���|C���~M�>	JE?yU_?e�?�����r�3�B��e��8��ZʼD�?6��>�?,�A>�=;񱾵�6�d�%G�v�>2p�>/��/�G��'��)��N�$���>�,?�>C�?;�R?m�
?E�`?A-*?pD?��>�%	��hF&?Ã�?=aս�T�X�8��E�~%�>��)?��B�ρ�>v�?��?��&?D�Q?�?��>�� ��L@�+��>@Y�>�W��Z��G�_>��J?,��>�,Y?E܃??>>J�5�l٢��
��V��=Q>��2?�/#?�?���>`��>���`��=}^�>�fc?��?��o?���=��?�42>D�>�i�=\�>(��>m?�
O?9�s?��J?I��>�ӓ<���������q��YO�&pz;ccP<��}=���>t����:,�<��;r:���Vu��f}D�6.����;Ap�>�s>o��d�0>��ľ�.��A>H��ۛ����$�:���=D��>�?�ѕ>
#�k��=I��>��>����=(?P�?G?4k;z�b�f5۾��K���>��A?���=Y�l�����]�u�?_f=�m?
~^?]X����
�]?�q>?��̾q!��Ԭ���)�J*��Du?��?PȾV�>��q?.�?�g�>L��4ws�靿������L1>
r3>�<A���e���v>s�?6"T?���>Aē>����ޔ�8萾b��>��?W�?�Ô?�{8>ane��п2��a"���^?���>Ey����"?�{	�tоv닾;ߎ���ᾓ˪�k���<�������$����:x׽|�=�{?k�r?�8q?	~_?�� �Ad��@^�
���V�$�Z����E���D�q2C���n�V�T����^��>C=&&e�7�A����?�6?��7�t?p������W;�l<>
����?�q�=⺽D�5=`��=��e���罩	���~%?F�>*s�>��O?]�i�q&6��J�� 1��D���x=���>'�>B��>���H.)���a�xc���4��A����v>�Yc?ĆK?��n?�M���0����&!�T-�⧨��C>9W>��>�0X�C���&��~>�Sr���X��Ŷ	�QW�=�R2?-6�>]�>�'�?J?`	�}��@y�PM1�z��<nu�>�(i?,�>`��>�ϽH� �g�>�2\?���>2#�>}]��V���%���
�e��><9p>[a?У>�λz�_�g��餖�%J�	�!>�W_?)������-��>��O?�/=*�=�ω>�ˣ�$�-�TVվ��,���;?�> xO>P������&�S��i˾zg+?4�?�8��:�)�`�v>�!?�?b3�>딈?�҉>M1׾W�<�u?t�`?gP?�"??<Q�>!L=W>꽻�˽<����L=Y��>?�K>�z=3�=	��p5.��S�ck_=n�=Y���*51<�%!<��<�W�;B>��ۿ�I�%�־�7�z����
�4'����Ž8M��������l���b�x�`��^_3��W���e�#����q�u�?l��?aے��U�������뀿�� �5�>�fl�u�y�#ǫ��������>�ܾ5�����!�NHO�q�i��f�6�'?𺑾߽ǿ찡��:ܾ�  ?�A ?=�y?���"���8�o� >EC�<t/����뾲�����ο$�����^?���>��0��	��>>��X>xHq>v���螾0�<��?:�-?���>ǎr��ɿY����ä<���?!�@�|A?��(����V=ΰ�>�	?�q?>!)1��4�����e�>�;�?4�?��L=q�W�+R��`e?R<��F����a}�=i��=G�=����J>=I�>���!�A��(ܽ�4>R��>S!��|��f^��:�<:�]>Raս���7X�?�Z�����a-��=N� �(>&�G?��@>�!��.X?�]��ÿK�c���?�|�?c��?�?�잾�t�>�ƾˀw?�5?� >d�n��j��5��<I�7>pcc�FW྿�P��iv>�
>�(��$dB�� ̾B�Q�:�#>��g>g���ƿ��$�b|��'=��D�[�Qp������T����Xo�����h=��=-vQ>j�>iW>�+Z>�fW?<�k?gN�>�>\:��~���ξ�F�����۪�����ꣾ�Q�|�߾��	��������ɾ'�L��5�=D��(��X�"��pb�M`F�M�?�ӹ=@y��Rd?�ٳ=�ɾ������Ԩƽ=�Ҿ��0��q�b�?�7?%��UY��������"�l�L?=�Ľ�<��)�����=Ѽ,9�=w��>��N=|�߾��9��Y�fj0?�e?�a��U�F)>6^ ��={�+?b�?�D<)�>�?%?�)�� ��[>Q�3>b�>-�>!C>WS����ٽ	�?�T?�p��ɜ�$ �>����d'|��za=zF>�p5����ou[>���<茾p�P��J��/�<��a?ۖE>������˾�$Ӿu����&�?܉1?"7=Ej�?0�w?/���X\�?���E��γ�k>?��?"�=D��V��!P��� ?/*Y?Xj��f�U��Nj���&�\-�M�$?O��?�?@=�f���f���*�'�?��t?N�a�u���{Z��
O��4�>��>[^�>!�;��w�>��>?ǌ(��}��BE��XP4��?	�@� �?��;�Q���=�R�>�{�>�e+�修�yrͽ��žo�D=RO�>h.����z� d$��)�h�A?�I�?�Z�>�z��������=�ٕ��Z�?��?}����Dg<R���l��n��d�<�Ϋ=���E"������7���ƾ��
�����࿼ͥ�>EZ@�U�w*�>�C8�]6�TϿ)���[о�Sq���?L��>S�Ƚ����A�j��Pu�a�G�2�H�ť��tT�>��>�ǔ�.�����{��j;��e��?/�>���U�>l�S�����g����5<��>���>f��>����9񽾳?b���?ο����Γ��X?1p�?n�?�v?Q�7<�6w�~�{�(���-G?��s?= Z?�%�XR]�'T8�`�j?ϩ�^�_��>4��RE��"T>P<1?���>�&,��q=>n��>LY>>u/�p�Ŀu��fz��a��?�=�?|��)
�>�]�?��+?a��h^��Lp���*�6.����@?��1>޶¾����<����
?��/?�,�*h���d?'a��y����w,��8>d�?�N�T�վe�?��K�=b��̧�A���}j�?��?!ر?��� 2���?�K�>�3����x����=3�[>�!�>�>5�����>-�C6�°5=�^�?�U�?XI ?��L������<w?_�>�1�?%�=M?�k=&Ձ�V]��V>j�>mP�m?+�@?c?��D=�It�Z�*�Q`F�lF��i��H�_��>%6j?�vD?��>�!���sI=��"�Ir����3�'���Ƀv�[W��C�6;>P��=�L>�4��9�Ѿ��?9�5�˿`���Y��7M�>�rv>g�? ���T��F��=��]? aw>\���0������~C�8��?�5�?��?�Ѿ�`�<��=�lt>�~�>>f�B7��f����>�G?>_��Ʉ���[��.>�6�?��@���?��u���?hQ)��N~�,?����������)>PD<?_��oG�>o�?9
�=��f�P*���Xt�Օ�>���?��??~�>�Ei?�{N�O�y�<TO�>�d}?$1�>�M=������Q>J��>�=�����1��ob?��@5@��T?����ѿ�3��:x���̾�g=��1=�>����:-Ͻ�=���=�%:=�N�=ƾj>i�>�:>0>�,>g��=�D��2������v����X�/�,�Q&��;��G����F��w�������ܾ,i��G-����@���<����o���!=�o?�AN?�cu?E0?d�׻�>�WҾO��S'��F*=pg>ݣ?`�C?�"?�«=�I���r��邿Aؾ�����D?Ä�=ݴ?0�>�W�>̔�!�D>�ڱ>�Q�>��>�~̼�!<�x�;�r�=ߐ>H?G��>�E<>�>ϴ��1����h��w��̽f�?2~��ʼJ� 2���7��'����n�=�b.?�{>���k>пh��� 2H?2���C)�.�+��>a�0?dW?H�><����T��5>���j�Lb>�' ��yl� �)�:"Q>Yl?��f>�ju>��3��A8�n�P��N��:�|>b<6?d���Z�9�s�u��H��2ݾLgM>�̾>��>��i�T���:�y�i���|=�x:?p�?�����ذ��wu��e��ҧQ>�9\>�/=a�=��L>Wqc�A>ǽ�H�/�.=�X�=t�^>�W?��+>���=�>�^��88P�[W�>��B>W*,>%@?	*%?���9�������.�~�v>10�>��>�[>�\J�h�=�w�>V�a>���湃����'�?�VPW>��}�4�_�a�u��x=񗽏�=�'�=
y �p�<��O%=u�~?����.���U�����z�D?��?��=��/<��!�U릿�����?��@���?����UV�fQ?<#�?�q����=���>� �>��ξ��M��?�D��"d��ib	�W*#� �?NĠ?��0�����άk�h�>��$?�^Ӿ3Ⱦ>��'��I������� p�]?<�(�>��I?%�������*5�Lg?��?�!����*�ȿ�Oq�b��>���?���?S�k�tЙ���A����>��?�T?�4o>Eq־C�Y��ɐ>O�@?��N?���>�]�"f4��)?o�?9�?�<c>잋?J�o?}�>�_���*ȸ�Վu�oF�=�K�/ٟ>��:>t�F�ɔA�P���w7��i�o����r�F>#�=�c�>!ۨ�^�¾5P�=���c؍�'pa<޾�>pgd>Zw>���>zR�>YC�>��>\=���`�_�8⟾v�E?0��?����F�����Ĝ+>�銽b�J?X�?�����ᾈ��>�1_?�q?�T^?¸�>�B�i��:Ӳ���㾕I^>q�>��"?X!@>^P*�,U;�޾'Oؾ�P<��?�����b����=����>K$?2�=C ��� ?*#?K�i>��>e>E����p�F��r�>��>S?��~?g�?�ܷ�x�3����d���c�[��N>ky?��?N��>�7��f&��
�K��=�ѓ��1�?�f?bN�J?⦈?�@?��A?�rg>�=�Esؾ{@��	�}>Θ"?���*B�>&���4�?`�?���>fg�o���&��[�"[��?��]?�%?�0��v_�@nž�S�<aڻϻ�\��;�}�"�>W>C�����=H>`�=(�m�#f;�W��<���=�>�*�=�=�烽MH,?�/R�^ ���7�=�r��HD�l�~>��J>9���^�^?O$A���{�����r(��WR����?^d�?(;�?Ӿ���h���=?e�?�E?A��>{+��!�޾���;$x�~�x�n��S�>+�>=��k|�t����d��'��oŽ6���Z?$ߪ>A|?<?2U>V��>�H��$�-
����� �m�j%��9�C�����(��45�B�<�ɾ ��+��>M�,�,��>Vy?��H>�]>G��>��t��>��Q>�zu>�q�>�+>Ul>ҏ=>��<K-���7U?l��/�+����Ѣ�%=?��t?��?�6�=�w��V �T�$?ř?ԁ�?2�>Q�N��0��
�>��>��r���?�lL=�9���Sͻ�p��������(�=�}�>O!�c2��	P�NW,��q?�� ?eb������Y��^��9#o=/A�?�(?��)�)�Q�3�o�2�W�?S���k�g������$�op�ݏ�IP�����	�(���&=e#*?��?Le�^���M���9k�>6?��/f>7�>O�>���>ASI>��	��r1�i�]�BN'�	�����>��z?�l�>p�I?�;?�P?�>L?�ӎ>���>��zH�>�Ȼ;y�>2��>�9?��-?/!0?W{?.P+?�b>t5��Q7���"ؾ�?��?�o?]�?�?]9��ZŽ�ˑ��mi�u�y��]��:`�=���<��ؽ4#u��4V=/T>=O?@��0�7�m���@j>�-7?(;�>��>�*��t遾iG�<��>!�?q�>�� �Ks�9����>�7�?��7�=�+>���=M�o�36��W�=���S�= �p��AC�Y�<���=ٰ�=�A��rU�9P�;{�;h��<<�?G.?(fA>5��>�Kؾ��
�y���=>���>���=���>04վ�B���Z��抆����>�֝?�H�?#�W>�P>�%>������@�姾Y�,��ҽ��+?6^?%5F?�!�?S��?d_�>�ƣ���&�I!��Һ���˾�O�> !,?��>1���ʾ��Ĉ3���?�[?L;a�2���:)�[�¾��Խ��>�[/�j.~�h���D��d��0���w��͛�?���?A���6�4v�翘��^����C?� �> W�>^�>Q�)���g��%�31;>$��>0R?฼>m]O?��z? N[?} S>��6�S���_����$���>�??��?Ə?�8v?͏�>l�
>-�1���ھ@���y6�����/����@= bY>E�>R�>D�>�\�=6�ƽQ��b=�,�=��f>�h�>y��>s��>M�v>�[�<��G?���>�N���p�S
��㲃�=���u?���?�|+?(l=�����E��P��a"�>�n�?��?�J*?��S�%��=�?ռ$�1r�� �>I��>���>�R�=�H=O�>��>��>Ǜ��a��}8�"M�L�?�F?إ�= �ƿ��B�����׾Z���jT��t��a��Hؾ�ߦ=�.��T�<'��׭��f#N�=��d����J����?�Q���ռ�#P>r��<4�޼��A>i�>,�N�\��=�w�����te�����&����<�J=��=���>���̐?�X�?�3?�$m?���>�L�>Zc	�;�>+10�!��>��>*�~�Y"�D,н�ޗ��#��^��ܝ�BR�_m��@h>�|�a�>�)M>��9=��C����=��+>�I�9�X9=e��=�a�=�1�=��X<��=�!*>��U>w:t?�󌿮"��`�X�#��=\,0?��]>��]<����U?O�>���r��Od��ly?Ј�?���?�?IӃ����>埰�a�Y�^D>;�*>���>u�Y����5Ǌ>�>=�8��ݥ�(��S�?0�	@xbO?�)����ҿ�[;>�/7>�>:�R���1���\�:�b�G�Z���!?�L;��5̾CC�>�.�=k ߾m�ƾ�o.=�36>C�b=;��Q\�^�=��{�x;=�Wl=oƉ>��C>��=v߯�!�=*J=��=��O>8��S�7���,���3=<�=��b>~(&>��>f?�c/?��h?`��>>c���˾÷�� �> E�=�K�>q�G=��;>��>]�3?O�E?��O?^4�>�=8R�>��>�-�R�n����I������;K�?^ʇ?SY�>�$�<��9��3"���=�nh�Z�?�41?� 	?���>
�4M߿��%��#.�W�r�<+=�=q���d���	���ڽ���=��>+S�>(�>'�y>�y2>I�E>v�>��>3��<���=Dz8�	h�<іZ����=��V����<����p0�6�`���*�V湼��<_��M9<WS<p<�=~�>M�=d��>T��=̀��}x>WS��u�G� xV>y6󾙼Z��l��{�Wx�["�Ge>�1>�5�<T���c�?b�E>�49>+��?�re?I>�l*��N��IC��:��])a���p=��=�����=�Un��XH��	����>���>[��>Ac>��,���8��)*���Ͼ��$��r�>ced��s�;p��=r�Q_���΢��1o�'؎<F�B?Y6��x�>^�~?	OL?g!�?���>:����پ�~�=tw���=C���,��	,��?�9?��>UӾ��P��gξC��mg�>2"L�I3L�q@���,��>�;aۻ�J��>K�uȾh�/�傄��<����C�#�h�9�>1|Q?oh�?9�n�u.����P�)l��4��� ?� h?ZȞ>qF?�?�;��U!�Ս����=��d?���?nE�?�`'>_��=E���x��>�?S^�?q3�?jFs?NE����>�¥;��$>������=� >���=-��=��?)e
?pj
?��C�	�����a�p[�!0�<���=]3�>-�>]�p>S.�=�x=O��=�Y>���>N�>�d>���>��>:����g�2�?��Z>�q�>�,R?z>J(�(�	���=����վ�y��"d�x�ͽ�I'=��!�6�=�G�=�D�>�"ڿ� �?[�>�E&�)�8?;�����½&?7>ϰ�0�=w��>��>]Od>m�j>3G�>��>�_�>�?>4�C���l ����)+0��\c�Vߤ��	�>����"~-=���P�u��h8��7��2���	f���W���1�"*#>��?|�x���o��J6�#�=ӝ�>�V�>A+G?h�U��d>��Q>yl?N"w>rF������.��������?��?�a�>��=>!�P?�?ԡ��)'�=�7 ��^q�@�%��Fb�BA�&�[X�E7�S��Q�k?�?H�t?�i&>��>�O�?v93�s��e=JU�"�#���x>���>�rݾk�<�S��z%�^�)�r�n�^�W?�v�?��.?��a�▊��d�>9�n?�C?�v�?��:?aOT?� ����?�r�=�R�>:?]�8?$�?�z�>>��<��=�� ����=#=汛��죾w袽/F�;��l�>d�[�<�6��e43>��=���=&�>)A=�!��9�P���ϟ=@��>�U5>���>�]?|L�>t��>��7?7��"x8��Ʈ�b+/?f�9=ݮ��9��Qʢ����>��j?M �?�dZ?:cd>&�A�
C��>�X�>s&>r\>�d�>|��E���=M>Y>ť=�aM�tρ�2�	�����5��<'&>)r�>�*�>P@�ֱ%><^Ͼ��Lu0>��I���վ����jt���=��;���a�>�N?�2'?R�=y>��(	=��q��f?d,?mJU?8Å?*->�s��i�F��
?�˟�ŧ1>�VE�D��p��A����P�"��[c�=�`��GE���a>5���n޾W�n�qJ�,��/J=-��F�U=A�o�վ��o��=$�	>������ ����Jê�
'J?��h=�y��QkT�`/����>b��>r��>��=���w��W@�L������=���>>�:>�=��Q ��xG��:��[�>�D?XN`?	ބ?�H�s�irC�����~��5���T?�e�>��	?�=>>�@�=5Ͷ�%���c��D���>2P�>��܌I�9ܟ����[$����>x�?D<>0D?�R?3*?�"a?4�)?|�?檎>�Ž�G���E&?���?�=^0ս̳T���8���E�Y=�>�)?�C�~�>#�?��?_�&?��Q?ץ?F`>D� ��S@�4��>Ri�>��W��Z��N$`>�J?t��>$!Y?�ۃ?�=>��5��Ң��G���q�=x�>��2?� #?�?��>~��>P�����=Ş�>�c?�0�?"�o?��=;�?�:2>Q��>��=���>g��>�?UXO?=�s?��J?��>Y��<t7���8��'Ds���O��ǂ;�uH<��y=���2t�K����<A�;zg���H�������D�;������;�_�>:�s>4	����0>��ľIO��9�@>,����O��bڊ�v�:��۷=���>��?M��>�V#���=Ѯ�>nI�>����6(?��?�?ͮ!;��b��ھ>�K���>�B?j��=��l� ���)�u�8�g=J�m?a�^?��W�X%����`?� T?����
�#�]���Ļn�5���z��?Jx�>9�}��_>b�?�"�?D8?�Q:���y�}Ě��K\�륞�]��=賠>|fD�D�v�s�>h�R?�?�Ӡ>���>W<�*��������> |�?�0�?	ٚ?s�3;,CK�T_ֿȂ���A����]?z�>�8��� #?�
��Z�Ͼ2e��k-�������,��#4��a��+�$��郾�|׽�t�=�
??�r?�Oq?I�_?�� �i�c��2^�,��VV�t��}��E�}E�%�C���n��U�I�����4�I=Kn�P�<�?"�0?L�.��� ?�ځ�
���	Ҿ+s,>�歾�52��1=��5��=�n�=(�_��'�裾�Z$?�$�>���>8�G?5oa���9���3���6���־�@C>o��>��>���>�?$9�yQ�sc��X��-0W�r���3v>(yc?��K?��n?j�](1�ń����!���/�d����B>�c>˺�>G�W�ږ�P9&�?Y>�,�r�����x��*�	���~=��2?A.�>{��>[O�?�?E|	��h��Ghx�L�1�O��<�/�>0i?�:�>D�>^н� �-�?&Z%?wy
?�y�>�����߁��Or�v�6>���>��>Q'T?���> =vD?�{m���咿�3#�Ն>)	l?7.���h���ș>��j?I)�<���>r���=������K�v#��2@>?<�>>ϳ]>�������w�8j���+)?C?M-���*��i~>("?��>nj�>x6�?���>_Sþ����?��^?z$J?�@A?��>N=�P���bɽ�&�#0=���>��Z>�Qm=��=���8\���3�F=��=-}ʼ
5����<�Z���M<��<��3>Pwۿy�J�_�ھ3 �����
����������}	�bm���R��6v�nz�O�%�'�U��Pc�Q����f�m��?��?c��W���6���=���8 ��p�>,�k���U�t̨�v� ������-����� �:�M���g��e�Ï'?G���ǿ���8ܾ: ?�; ?�y?G��"�*�8��� >�
�<�S��ȡ뾣�����ο����<�^?=��>��w�����>§�>q�X>�?q>���잾?|�<u�?��-?���>K�r���ɿ񉻿N��<���?��@�A?�(�x��ûW=a��>�
	?٨>>�*1�P���į�u��>B�?(؊?<�C=l�W�����]e?��,<sF���ػ��=@��=6�=F��vJ>���>���[�B��5߽�W4>{	�>֓���۾\���<�Z[>��ֽ�ꑽO4�? �f�	$Q������W��%V>�Fv?x#�>oщ=B�5?Y8��7˿��^�,qw?a��?ɾ�?L?nݾ�u>\׾؜o?/=D?D�i>W����)}���=R��<V�=W���}��hT>�%?��s=��ͽ�7��ܩ-��ߍ>�[�>R4��"���+�p,��;��Kڰ��������N�W�̽z}��F�y��Ӧ���>���=��.>b�N>�"2>�A�>��Y?H*_?��>�\�=!�vh���n쾙�E�����<��-�
�=�������1���p�����:��3�ξ4#=�2�=�6R�ɗ��� ���b�?�F���.?co$>^�ʾ�M���-<anʾ����턼⥽�-̾ϗ1��n�Y̟?��A?z�����V�=��Q�܍��ȪW?�V�$��:款���=wz��|�=� �>ʊ�=���A 3� ~S���*?�%?�mɾ!���4>��ԽZ�m<N�-?��?ו=�UK�>r�"?�K�N1㽜�U>_�7>~��>-��>�=���t��T"?�6P?����ĩ��lD�>������q�&��=O�>'8����_ �>@�=������ػ����<�[Y?�{]>cξ˙��;��w��U����-?��F?j1?h�e?n�g?����I�~�j������>���?&O?�/>�@*�����[�r�M>?>�*?�ϥ=��C��"�s}H�����~�?�_?f?��n=��J��@�������J?��u?��`�+
��u��9�.��˪>�p�>Lw�>��;�ſ>N;?Q���?��+���{2��~�?@��?`�v<��ph=&�>~>�>�$%�U`���!ٽ�8��R�=�A�>jӣ�vzt�������r??<]�??F�>Ő�������=wٕ��Z�?��?G�����f<L���l�<n����<�ԫ=���9"�����7���ƾ��
�!���iܿ�
��>Z@JQ轍+�>�A8��5⿻SϿ����\о�Rq�x�?��>�Ƚ�����j��Pu�߲G���H�>����O�>�>2���o�����{�Sr;�J��<�>����>�S�D$�������4<H��>X��>G��>����罾Cę?�a���>οW��� ��h�X?h�?�k�?Oq?��9<��v�S�{�k��#-G?��s?KZ?Z`%��:]�)�7��j?Y����_�Q4�]E��5R>h�2?&��>�>-��~=�z>Þ�>V�>j	/�G�Ŀ����X���b�?R��?(P� A�>3X�?�+?�m��R��pЩ���*�[Cĺ�DA?�%2>���(%!�!�<�����,
?>30?�� Y�,�_?��a���p�I�-��½Id�>-/��]����r��d����i�z�l��?�O�??!�?C��5K#��$?��>TȔ�a�ƾ��<+ߥ>��>�XO>�S\�sUv>���A ;��>��?�@�?��?�Y������i>{�}?1�>�w�?�(a=o��>B�>�߇��j�igT>��T>�ս�	�>�TA?��?�T�=Τ��A�^�9��/P����	�E�X~>�Wu?�D?��j>�����X/<M�!�Èڽ��*׺�:E���G�D��:��g>��=��=n޽��þC?��!�:�ͿTԝ���F.$?`��>��?�1��q��q�<� a?h�V>��5 ������ę��G�?C��?м?OlԾ<@ɼ�>�=�Ƽ>l׃>��߼�=c�D���J�P>�+9?��Nv���wm�xb�>hT�?.�@%�?��c�@	?����w��h��8��4o>K�&?Q<��J�>m]�>+�>>T'{������n�3۞>��?��?�� ?a�w?X�t�L�J�Q�,>V��>��o?���>qf��A�־��>#H�>n������h��+1t?Wz@%i	@6�E?۵��D�ǿk����﴾�?����L>��=�ۥ>e�I��J����T���vK���=���>�]>_�>���=� *>Do�>Ӄ{�����Ѵ�8���N=�(���|�J�/�lK+���Ǿ�-����$˾�m=ĝ��CP���k���͂@=�e�<��v?�|[?B]?��?Zt=�"J>��Ҿ���=�-t���<��j>zT1?!L?�y*?4�J<����$0`�dQ��u���42��L?�yz>߱�>�`�>+��>�O��ͤ=3G)>Ƈ>Hn�=�¦�w��<��<�+=��>�X�>�E�>�C<>5�>ϴ��0����h��w��%̽�?Py��7�J�U1���5�������W�=�`.?>�>W��7?п����M.H?�����(�G�+���>��0?�_W?@�>���v�T��?>���p�j��_>�2 ��l�)�)�*.Q>Ik?�c>��>�6��7�{pJ�io��ڨg>o�7?#���s�M�Hys�߸C���Ѿ��<>h"�>T�}���1����~�*�u�3)_=��8?JH?Ӗ��wU���\t�m-��rjN>u�h>�1^=Y��=W$Y>u�4w˽��K�N�=
�>��Z>�'?��&>�Q�=+�>qڢ�
?V�F|�>5�.>RN>P�E?�3&?9 ��������B�L�4Fa>x��>��>��>M$C� ��=�"�>�`> @&��!4�����<�	R>�g���}e�nV���=p骽�">_x|=���Z�4�Cg=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>�������MM��Q�t�d�=�`�>�G?D���K�4���;�I?	�?^c�Rl��D�ȿ#du����>���?�/�?ːl����#A���>t*�?@�X?�Tl>��۾k>P��*�>�}@?$hO?k$�>�j���(�Y�?O�?���?�S\>׍�?V�z?-Q�>�N#�4�8�]��勁�&�=��=X��>��>j"����F�3̐����"Xe����oB}>�%=]��>��̽�ѾSa�=�8�����}-���>(�t>"!>d�>?��>C6�>#�(=Lն��Ǘ�v��6?���?BE+�MTa�#��=� �>��*��!C?B)f?0�ھ|(��b?W�m?\�/?�LV?N��>c�@�^���׸�Ԋ��sR>�,V��	�>��>��f�Ћ㽪���o��w�>w۱>��f��<�R
澜�-�5ѳ>,�*?8W>��%>��%?ω?Y#�>��>a�,�6��|5T�O%�>6��>9�?:�?Ē?�qG�g5�����3����Q��Z>��?.?~��>�J��
���Ak��I���D?�?�7C?����O�>�)n?�G>?�X?!�K>�餽����t�B�]>##?��t�A��#�j�Z;
?
�?���>����@3���M��#�� ���?`^?�e)?U��4Dc�E�ɾ��<>��:�|;屴;V���>�%>0[z�\��=X}>���=6�v�8+��a�<xz�=j͒>��=�C5�NPe�oQ,?>�P�Y?�����=�Ms��*D�2�~>�I>YS����_?��:���z�bȬ�ʝ�� Y����?`��?\��?�ӷ���g�==?�χ?�?vR�>@����AݾZ'�Ets���w����N�>KX�>��z���q9��39���΃���ýC4�x?��>��	?��>�v>䀾>�B���//�C�����rb������7����A�_v��=&�� �L�Ǿ0�~���>8�2���>
�?�Ɗ>E��>�ը>s�< ��>�Dk>"��>\�>��->�>���=Չ3�2��HgR?�R��_b&��F�Ĉ��u�A?��f?L�>Y�	��q�
���#?�Ŕ?�؜?�7�>jMe��/�ƽ ?�>�1~��{?���<
w����<�9��6B	�b%��V���S�>�zｩ�5��'N�(��1Q?��?ڗӼ�;���ò��H�e=�?�7(?Z�)��rQ��mo��_W��S��o���g�+��{�$�iAp�ҏ��_������S|(�xG/="+?տ�?~��i�ﾧU��Pk�K�>�EDg>��>g�>v�>L>
��h1�^���'�W_��x#�>�{?�PT>�^?&�1?��<?��J?��>|��>ꎾ8�?H�P�V��>C/�>5D?��4?�1?ϫ	?�?z>�KK�� �_5���)B?�?�<?sC�>G ?`˘�\��q磼��h��D|�QI�@��=,U�=�<E��D���;=2lA>�X?���ɬ8�����Sk>k�7?��>{��>���*-��\�<z�>�
?G�>G �"~r�c��V�>���?���'�=��)>���=f�����Һ(Z�=������=�5��z;�%e<���=`��=Mt�c2���7�:V��;Yn�<K�
?��>�B�>.��>OF��E���5�@6M> ��>���>(�>��� ��(����y��"��>j��?#:�?��>Q>�%��	���!���}ľ�ڷ=��>��?2�`?���?��^?ɫ?�ώ�����Ԕ��*-��W����>>",?��>���ʾ��J�3�˙?�\?q8a�}��2)���¾��ԽD�>o_/��0~�4���D�K!��8��t�����?W��?�A���6��s�N���\a���C?��>�W�>:"�>ҿ)���g��)��0;>���>�R?TG�>��O?WT{?p\?rbT>��8��"�����uV9�gU">6+@?l��?7��?��x?���>�>c�)���߾M���v�A��2|���GW=PWZ>��>g��>j�>�%�=ǁǽd�����>��-�=9�a>���>V:�>ƽ�>��v>̹�<�G?���>tN�����K�о�(��v���i?-�?�#>?�>���PH����U�|>OR�?���?��>?hZ�x�>��G��V��
�����>s��>_d�>H/���=٨^>�-�>���>�Y�����/����S?H�@?�%(=ꢾ��AQ���ھ y��Š �lD����߾���~�о�<��f�&��������_��]��Hژ�ޜ׾6ں�81���?vw��=��->cr$=6��=�=��9pѻ ��<W�= S=��:;������f蜽o�.��o�<҉��[���v�?M+�?��5?5_?
b�>��>F|���4x>�H ��'�>��=붷�׉���0ؽ�þ�ƾ��羪5;_:%��ص���=�<4#?>�^(>�"=L�T=���<��M=c��=�:=�����=IKZ=�I=M��=#�>�8W>�w?�Y�������$���>i>?&%�>gh��|���?xC?�͜>�5c��)��eݧ�5t?O��?�H�?�k�>��ؾ��>�˕�׉`��Vp>����x�8>	��=��k�.T�>���=�������������?y*�?R>D?_[���ӿt���]4>w>��T�Z0���O���T���e�@�"?{�3�.IӾ���>��=��Ծ�ɾ�n'=]:>4�M=�d,��f\�=�t=���`�U=�w=5��>� B>) �=���=A��=��>��F>K.<� ռTn0�XU=�d�=�	z>��">��>n#?YL7?q��?3�>�!@���޾�˾aq�>e��=��>���j�=Ey�>�|?�Z?K?{A�>��K>���>�>��3�8�l�{�%���f"����?=�?�u�>�l>	�5��8 ��@���	�?l�7?*�!?���>�@��s����B��3�=�̽��;���=咾ʣT�Zd��$�{�3�����>���>��>=>ߢ=��=o�>�x�>G�>
� =n�}�YT��@��y��I>���<��=�JG�n��=�׫�>Դ�>�j�q�.=�ib=�1�4QƼ��=�S�>D�#>n}�>NJ= |��a�8>o���4jN�ܮg='i��/FI��i���x��lN�#a!>�MW>����C����?r�P>�8I>	U�?a�m?p�K>43�����6��k$�;�1�=Ns�=U6S�Λ;�
1f��"L���X��>2�>&��>g�>�)�׭I��[B=�Nվ��1�Ͳ�>k�#�����7l�y1��z=��c�e�B%<��@?5`���>��}?~pO?��?��>�՟���־�i>�O~�CI;�A�u�C�Mi���e!?r�?��>��龫f@��¾�; ��ɞ>�ћ��&@�����L)��b���ϾF-�>#��s$����.�95y�Xa���ZP���a��г>lb?���?cZO�,5g���[�^;���ﹽQ�?��c?b=t>I)??1dJ����J�r��
=�]?v�?]?�?�YU>K��=�㴽H�>�,	?���?���?��s?y?�,t�>Uԉ;� >�՘�Y;�=�>���=s�=�m?p�
?k�
?�X��-�	�q������^���<���=怒>lj�>��r>��=��g=yk�=�0\>�՞>�>��d>d�>�V�>"����f�c�9?  J>Ӓ�>�VB?Z��>��ý�#V�hUf�p�	��������5&��Gb<�p�=�_I����������>gCʿF�?�J�>���}�?�۾������>Ӊ_>�D<��T�>b�->/er>Yk>��>	֊>՟�>糶>H�վ�tE=�>���!��b7�>�A�B.Ͼ9Q>�s���/ǽ�����A���J����
�:Ll���x�9�6���=ø�?v7	�O�K��6��{��z�>˅�>��3?�Ǜ��I�=��(>c�?,�:>��꾭���@�������s~�?>9�?>�v>�J�>�-b?]�??3�Z������@�mʁ��$5���V�|@f��i���z�: ��:����m?��l?J�8?��=� �>}hs? �%�ܽD�E�0>��@��P��H>B�>&�x��X�z�߾�ߑ��[�!0�<�kr?<p�?]�'?X����q��(>'<;?��1?�t?LN2?W�;?���L�$?&�2>8?2?,E5?&�.?o�
?��0>���=੿���(=�y��k����fҽ�Qɽ=^���3=��w=�2�86 <�E=;�<�-��ڼVh;�����</x9=*U�=?C�=�ݧ>,�\?dp�>#��>n�5?�����7�����D�0?��Z=0>��熾� �������=��i?�$�?��[?�7c>�?��@�+N>-y�>�^+>)�\>�3�>ܮ�}\E���q=�>|�>p�=-V���}����A���W�<[6%>���>�s�>N"�=W!>�C�?��B>I#о�%ɾlZ��>g��A�9������>@�k?&�.?�>˄��5�I�e���V?�-?0x'?��y?�g><j�S�C�'�U�Y����?�>��a���#�<=��y���\eD�a�1��\>
꾔ޣ�ka>}w�X߾] n�I~J����c�C=����P=�$��*־���T6�=��>W ���!��M������o�I?ݎf=Dx��۟U�򎹾%\>e�>cu�>t6��ǀ���@�Q�����=I��>��:>~���s-�JG������w>F�F?��_?ik?t�W��d��*;��9���Ϛ�1�[��?2�>#?я?>��=�*��d�1�c�ht>����>X
�>��$���I�W���u��-�/��X{>.�?8�>��?��V?��??T?��!?8�?�w�>f˽k��R@&?Շ�?*�==�Խ�T���8��F����>1�)?��B����>��?�?��&?h�Q?(�?%�>/� �G=@����>�S�>|�W�Ha����_>ȨJ?��>�?Y?-؃?��=>q�5�]ꢾ�驽��=A>�2?�5#?!�?���>��>ٙ��]-�=��>��b?X.�?��o?@��=��?�c1>���>�ٕ=��>j��>� ?�;O?ʶs?]K?-��>��<�3���7����r�vsN�9-i;�bC<��y=����s������<4�;'��%Q��z��` E��'����;��>M�h>�5��G�X>K�ľ*<]��SY>󺐽�b��� ���*J���N=���>3�?��>�!�W��=!u�>��>���T�&?j�?=&?ED;�]��o־�
2�(Χ>{�3?0�l=Q�j��|��@�q��T=�d?HT?��3�� ݾ�nb?._?�Ͼj%f�?�Y��&<ko�JXW?��>�������>F��?ƅ?��?�#Ѿ.�]����I��	y�P9�;8_�>���?)����=`�J?D�>I3�>�=���l�`��Ǿ��?(�?j��?*m?�>�|O��aٿ��������0\?���>�}����#?�,��EѾ�����_���7�>.������8��TQ���%�B߃�9+��a��=�<?��p?�s?�^?Q���-Od��y^�ټ|��
T�������>�E�ՒD�(�D� n��?�f���h�� �{=����8���?�W#?P����>;n��Dn�tUɾӔ=>�瘾�g	�2�=x�z� �^=C))=��l�ڽ0�;5���Y ?0��>�f�>�4?]]P��r;�C�8�,�6�qF�A?6>E�>�x�>XP�>�����1�G���%¾�Ć�Mײ�6v>Ryc?4�K?f�n?�q�5)1�q�����!���/�]d��(�B>�g>E��>l�W�V��<:&�UY>�R�r���+x��
�	�*�~=��2?(*�>ϲ�>�O�?�?f{	�5i��Glx��1�ҍ�<�0�>�i?m?�>1�>�н� ����>��l?��>V�>�ǌ���!���{��ͽT��>�[�>t�>��o>�/��F\�C���=����8�y+�=�?h?2����`���>�R?P�
;V�M<�ݢ>�[t��!�9y��'�.�>��?V3�=� <>��ž�4���{��	���=)?NR?�͒�U�*���~>�1"?Ue�>(�>W'�?��>�Iþ�h�P�?b�^?�6J?�?A?�&�>�2=����ǽ[�&��`+=�w�>�[>��l=ę�=���[\�o���E=_��=qм���:6
<����\�I<&t�<��3>mۿ�AK�A�پ����?
�M눾P���e��*���f��h���cx���TN'��0V��=c�����ϯl����?�:�?.����5����������������>ҍq��W����m"����ྀŬ��b!�[�O��!i�e�e�I�'?�����ǿ𰡿�:ܾ2! ?�A ?0�y?��8�"���8�� > C�<!-����뾭����ο>�����^?���>��/��f��>ۥ�>�X>�Hq>����螾�1�<��?6�-?��>Ύr�/�ɿ`���X¤<���?0�@�G?��6����u�	>{0�>
 �>6z>�c�)�3������>��?ʀ�?X�3>�
C��X��>BU?8�Z=3�9��-
��H�>�nw=�=��sbV>��O>�Pm�Q�a�K�C-~>\=�>Y��S���q�����=��x>�/L�*,�5Մ?-{\��f���/��T��U>��T?�*�>M:�=��,?Y7H�`}Ͽ�\��*a?�0�?���?$�(?6ۿ��ؚ>��ܾ��M?`D6?���>�d&��t�߅�=y6����{���&V�o��=]��>j�>,�����O��I��^��=��.�ƿx�$��|��=g//\�{��GЪ��NU�A��]uo��齣�g=���=�
Q>:N�>��V>nCZ>4hW?T�k?H:�>]8>0�`���lξ��>����酋� ��Cͣ�2M��߾o�	�������"�ɾ�VX���Y=G� ����Pnj�[K�N?�F�=�)���+D�C�%���Ⱦ���ǔ6�����0ϾN�@�b{�iW�?�$)?����X�u���۽י ��I?������oɾ_I�=(�I���P����>^L=����8��=Y�X0?�@?�5���ѐ��t)>o���u�=�r+?`?>y.<�Ϫ>C�$?e�*�W�!N[>3>Y�>�W�>ï	>�5�� �ڽ��?�`T?�y�;k��hH�>�н�|Fz�D_=M�>I�5�v!���Y>-8�<B;����b��.����<cY?T:�>� ��!���s�i���M�?+|?�(�>�̪>�Sn?>�Q?hR=2���]�X����T���N?��k?W�>ᠼ�ؾӨ;7�F?��s?l�>h�q����@��}�Ou?|~?��.?@�f;o��3��4d��(?�v?Au^�1I���)�Y��.�>?H�>�$�>g�8�ٴ>�!>??"��f��������4�bΞ?Q�@�d�?�61<~\���= k?�x�>	�R��>Ⱦ��������F�a=��>H/��U�u�5� �4o*��8?(#�?�~�>�-��D����=*֕�dZ�?v�?-����g<��:l��l�����<�ҫ=���*:"�K��2�7���ƾo�
�֫��^���j��>}Y@�m轢&�>Q;8�"5�nTϿ����Yо!Qq���?-��>=�Ƚ������j�Nu��G���H�d������>�u>����^��o�{�Ȏ;�c쬼���>.y�yF�>�V��5��o|���?2<˥�>���>���>BϬ�5��Į�?%���Mο ���<{��X?��?���?ُ ?,m]<�^v�Qj}��&#�HQF?��r?,Z?�9!���\�"�;���j?_���T`�ڍ4�HE��U>�"3?9A�>��-���|=�>��>�f>�"/���Ŀ-ٶ�����|��?ω�?Mo꾑��>=��?Ys+?]i�)8���[��A�*�C-��<A?a2>J���ȸ!��/=��ђ���
?~0?tz��-�E�d?����X��@���>��>�T������:f�W�
�P�~*�����k��?,� @��?��;�]H��w-?��>Q��D̾bs�=�K�=�*�>͚o>\�ѽ��#>a8�#1#�Cu��$�?3{@�*?�E���調��>�b�?��>@�?��=�|?�ª���S�H_>5E�>��=�h�i?�	0?���>���=������M�<�^��*�E�S���{>��p?$�R?fǡ>57��#�=�V��7��\���������(��I�@�삶=�I:=�=k>:�a�R���<�?p��gؿ.���s|'�If3?p �>G?j���?s��&k_?5 �>�Z��#���
���� ����?[�?�Z	?ؾ��Ƽ>T��>@�>�ԽT�������9>dTB?�)� 8��ʞo���>D%�?��@0߮?�Ni�K��>����{u�
Z��'�F�ؾ��:��nJ?z�׾2��>t*�>��2>�m�>᥿�{�0��>5��?���?XV?�τ?R�t�'�-��$�����>��g?�+�>�տ� ��3�>��>;'���y�q0ɾ9�X?�@[�@��R?
ո���ҿ:����]ֲ�==�������=�I/�v��I�O=�=��i�ϼ=n*}>9�,>,74>Hw">��X=5�=� �� f�#���"畿��9�RE�WE*�sb�I-�{����e ��Vݾ��ƾn�	��q�:��K;���~���ȇ���X��	i?�pm?��`?O�>Y�>^��>V����~<�pN��]�>��g=b?[)?�*?�Τ�P}��e|b��<��"N���?ƾ�$4?Mz<`�?77F>U�>��e�(e�=� �>�T>?�;>DQ<�>9����Oل>�k>��>.��>�C<>��>'ϴ��1��h�h��	w��̽@�?T���T�J��1��89�����aj�=2b.?�{>����>пk���m2H?����_)���+���><�0?�cW?H�>�����T�:>P��Ŧj��_>
* ��~l���)��%Q>,l?d�f>�Mu>��3�oZ8���P�;b��Zu|>\=6?g߶��r9�ڱu�§H�}Jݾ�OM>�̾>h�D��p�����1�J�i��{=2x:?�?,9��?ܰ�Itu�nL��=>R>�%\>�]=��=>3M>��c�Иƽ�H��.=��=�^>�
?�5>c��=5G�>&?��9�a����>�'>0#>:?7?�~(?�
���߽+]����.�؟w>���>6/�>�(>�jK��E�=g��>S�j>䊼�P��������2�"B>&b����a�.o���=�ꪽ�)�=?�f=��M�X��1=�ԁ?l9��fÖ�앾D<g��?�t�>]ӎ:�@��l#۾Q�������(�?m�@�-�?>��V�?�̍Q?�4�?D����@>�+?I��>m���y���>?�����`%��b�=�?s�?_H*=������DD<>�?j����h�>w��Y�������u�s�#=���>9H?�U��ŵO��>�Yx
?�?�^����n�ȿQ|v����>*�?D��?l�m�A���@����>��?�eY?oi>�f۾�[Z�O��>�@?�	R?��>C9�Ȍ'���?4޶?;��?2�H>挑?ߘs?jT�>w�v�C/�B0��������=k0_;sp�>N�>����`F��ϓ��c��>�j����K�a>�%=
�>����2��J�=s勽�d��g�6��>�!q>S�I>�\�>Q� ?^?�><��>��=�q������K���+�E?Jޓ?��R�@�4�H�?>�'��I?�B%?͆V�մ��?��>�f?J�u?� ]?xGh>KL)�.!��J���iѾ/�>M�9>J�*?�{g>��x��>�����8h�=��>����:���H�����>�T�>��?���>�=;)?F�?s�u>��>JJ�r����H�/��>��>�
?l��?}9,?�'���;��ᕿ�圿�[U��,;>�Aw?nA?�ʀ>�l��5����T�=>\�i�<��?�K?6L�=$C�>B!�?�+n?}8[??�=@=m���ݬ�V��>|�!?a��A��M&�i
�?�O?���>;��{�ս�Mּ����{��w ?(\?�?&?{��t*a�G�¾U(�<)�"���U���;��D���>��>?���{��=�>n԰=�Nm��F6���f< x�=Ӏ�>���=�,7��w����8?k:>�y�`����=�I���Do��Z>(��=ٻ����g?��=q1��M��9ٕ��^��� �?���?]�?3�I�B�A�� �?���?` R?��>���Zپ���3��d.��Ι��H�=��>����4�}9��g#���f!�f������>���>�x?��>�[>A�>���Vu*��� ������a�h�h�.��**�^��J������F�0ӿ��w�wK�>^�g�g�>#r�>�xU>��o>��>�<�>~>�O>�=}>#S�>1�T>��6>�3>5�;<*L��!�S?bѾ~A�W�۽y�ʾML/?��V?g�=�e��Ȅy�鈢��41?g��?j'�?b9�>`]:�bA����>�2�>xa����W?[�>����f��۽�"ؽ��޽2!ƽj8;����ΈC�d�N��7k�g�>��?#T�<ZJ��f�ﳾ*�=�{?b�?�� ��P���m��^U�{,N�����l�����Y&���o�cS��^}��0\��[;*�H�=�20?�P�?�{����������.Kn�5�@��n>���>��>>��>�t>C����/��l\�wb!��{��o�>Y��?C�>BI?h�<?�P?{K?˨�>B\�>ֳ��~��>�;?ݡ>��>W�8?��-?H�/?�`?P�)?�c>����Е����׾��?O�?��?�� ?�P?B셾�Ľ�Z��KG����y�����j=m�<��ֽW2�� d=}rV>&'?<O�`\(�K�׾h�X>�X6?!5�>k��>������y)�;���>:�?	�>L���Ml��=�ݷ�>/��?��'�\�<)	O>�%�=�����ŕ���j=\��{�=)l�<����zwR<�#�=��=ٿ�{ά;�>�;:��<�6�=��?�?(�>���>v6��,�����%�l=�&9>@G�=�6�>�ï��ΐ� �����Z�h0W>
>�?�X�?�`=[�>dS!=GV��W�����~٧�"L��B�.??��G?��?"B?��4?�>ւ��f�����C���X!?��+?#�>���_ɾ�Ȩ�u�2�ǽ?�"?#a��+�Q�(��	þ�BԽ9�>�.���}�vЯ�Y�C��"��4�gP��ڙ�?���?�	:�?�6��>農����K��7_C?ۛ�>�٣>?��>��)�G�g�z]�E�:>Nw�>�*R?�!�>m�O?�;{?�[?�pT>�8�I0���ә�YT3���!>�@?���?�?�y?�s�>��>m�)����N�����x�_䂾�W=�Z>�>~"�>Z�>D��=�ǽ�S����>��Z�=��b>���>���>v�>��w>O�<WS?V��;)���!�޾����Y���AH�
��?��?�/k?*4ɾ<�}���޾�R$��w�<�1�?�Z�?.r�>Ї�aI>x��ِ��D����.>�V�>IE�>�f����>�f
?�L�>���>�b���9�a�)0ٽj2 ?כ�>�m��o$ڿ��?� ���������<�澍F���S��f��ԣs�͵�9����������ʾ�T
�S#�9]0�����؄?1Ɔ��{)��t�=�̞='0�=Z)�=H�=p�=[��<4��c>=�Ժ�93����o��8�i<]>�6�>jm��v?ֽ�?��?ِ�?Q�3?���>�ɪ���>�_�=v(?l�a>�i�F2W=*Ⱦ�䲾��þ"#��Tg�2���<f�=� �=Y�躴�5>����m�=^p=�^=~FH;z����:��=�Ҩ=�$���t>rY,>��>�Oi?v���P����Aj�m >
g?w`P=�=ڪ����V?kn���:K��Ѣ�}��h�X?���?�E�?{��>�Dj���>a��{}��2��>/�Q>)`�>�`)>nY��>(��<���Fu��R5�5��?��@�pP?�W���ɿ3� >�7><>�R�i�1�a\�ib�e{Z�^�!?�B;�2F̾V<�>�1�=q!߾��ƾ?�.=�z6>#b=�q�@H\��=o�z��Y;= �k=���>��C>�
�=ZD��Y�=0�I=A��=�O>�՘��Z8���,���3=���=7�b>�&>L��>J1?��?�o?�(>"1��3�۾B���T>���w9~��;��D>��>(�V?�Ke?6P?��>�&C>8��>)�P>&�6�u�c��e;0�[��7�?��?^��>E�нZ@��T�p�`����6?�6E?���><�%>rU�I�࿓X&��.�􄙽�:j�� +=�nr�G^U�����w�ʹ���=Hk�>���>+ߟ>KKy>�9>9�N>��>��>U	�<�t�=�x��Ӷ�<*��F��=����J�<�sż."��)�%���+����HN�;�5�;��]<��;��>���>��>E7�>ݛ]=̾�u�%>"՚��vG��+�='����[=��i��[��6.�X *��DM>�G}>󚇽�,��o:?��b>��[>y*�?\s?�1>_:�]�ܾ�����f�>�R��K�=z5�=$�#���9�y�`�%UO�i�ҾK��>�ގ>��>��l>`,��?� �w=��Vd5���>�}�����&��3q��=��`���Xi���Ǻ��D?�D��ʝ�=� ~?D�I?+��?ׁ�>� ���ؾ&00>�B��{�=�
��#q�Bl����?�'?��>x�l�D�\=�Ӫ��iS>a�ɾ?o0�n~��M�@���=Cm��e̻>|ƞ��D�I!��ׅ�z����BW��z��w�>Ņ?�V�?��V��mU��Q�2�����E��>� �?�ĝ>��??ǀ�=^_�������=�fz?JE�?��?yC�>��=�<V��>:��>���?cp�?�g?}�[���>��<��7>$d���8	>,�	>��=�\=W|�>���>�Y	?72�,���L�����H�ƽ���<�L��f\>q��>7l>�A>Ji>+E�=�" >��p>+-�>%sU>6
�>
.�>�ݨ��:��)?���=��>z�4?���>�Z6=�¢���<t.,�[=3��C�M����ɽ`MQ<��H�\�=�j����>��ÿ
?�?3<>|���7�?@��sW�z�W>5U>rh½��>S�B>��h>��>�!�>.>c�>//4>e*�}��=�4��O$�+8�AP��ؾ��V>#���o!�(��w���\d�yR�����Fp�O8��!B>�`ք=�Ɛ?�8��+�c��,��-�2U�>}��>�:2?Dʃ���ؼnW5>�X? ��>���`��"F���n׾��?�o�?�h>�S�>��K?�<(?�I���$�3/=���u�C�X�+�t���f��ŋ�ą_�R0þL:E��O?�a?7�S?��>���>�dn?@_(���T���>{O�(�:�H��=��>��z��R���&��_���o�=�>�S�?Eވ?]�>M|��2彟�e>��G?)?.y?��A?*,9?�7���?̒<>��	?�"?p%?2(?��?|#�=�Մ=��IQ=^xj�m8���n#�����:�ټ}�_=�Oy�m� �̉�<z�=>��<����4׻0p+<���!=%��<�I�=k>��>��[?��>���>�//?�v9�K2�EZ��*?�=�T�3|�����������=g?hJ�?`N`?��W>��B��7��&>E3�>pD4> �[>|��>�qϽ�^S�9��<i5>��>���=�pt��qr���
�3Q������1>���>)�t>E-н�Yv>���u���6�>�$���[��4�ԾM�<�C�3�{P$��? r??�E?F�=�������b�0u?Xg`?A)?|Zq?� A=L⾿��8j ��l�l·>��6��f!�ҏ���Ԙ�O�>�gQg�fg�>st!�B�ǾYO>�'�WѾ�'l���Y�Ւоָ�<���8p=������־Wj�U��=_�=�þ�� �J���Ǐ���H?'��=*ڞ���[��UǾM��=w5�>Z�>7AZ��[X��6�����}�=	�>�PT>�'����_�J��8�<�>PE?�W_?�j�?h���	s�v�B�����sb���+ȼi�?�w�>�h?�B>���=~�������d�$G�� �>��>(��0�G�g:��R1����$����>D8?Ҭ>��?�R?��
?*�`?�*?zD?�'�>�����PB&?V��?u��=
�Խ�T�9��F���>��)?��B����>X�?¦?F�&?4�Q?I�?��>�� ��D@�ӏ�>�M�>�W��g��&�_>ԠJ?j��>\=Y?ރ?�>>p�5�C�񩽵7�=��>��2?%/#?��?���>���>�(����<�G�>_?�݄?�.f?C� >>�?/�]>���>�и=���>���>�@?�N?�~?!M?R��>>�;#�r��(����f�Ǩ�$�t<G��<�H=H_�&�#�����$6=�9������i�̼|��x�n��و<(3p<]�>�t> ���1>��ľ�?���@>:��-F�������:���=d��>��?ᶕ>�:#�d��=A��>:�>,���5(?��?�?�;��b���ھ��K�8�>=�A?>��=��l�ˁ���u�Bkg=��m?��^?"�W�'���j_?�Ie?0��&ܾx��+@齆��}g?��>Bt����>���?�;�?G� ?əS�r���Y��b�Q��:����/���>G澿$?���>U�?�4?l�>���>atD�������n�>}�?�L�?�;�?7�1>�c[�j�ӿ����:G��_^?��>f=���"?<�����ϾyO��&*��z�:�����=?���q����$��܃��׽��=��?�s?[Uq?��_?�� �Qd��)^����YlV��!�$���E�.E�r�C� �n�C_�`$��@��щG=�ǂ��C6�L��?B�#?)���>v����w��I�ľN6&>����J`��'�=炽�@=f#L=�n�ԧ(�����O�"?Sܜ>)�>sVA?��T���;���2�P&0������R>�ڱ>��>��>�
><��<�ڽ���S�V���ǽd1v>�wc?u�K?��n?�z��'1�ۄ��J�!���/�tf��U�B>�W>��>��W�Q���6&��W>���r�K��v����	���~=��2?`%�>W��>GN�?�?�z	��c��BYx�o�1�i �<�1�>�i?k?�>��>�Ͻ�� �P��>I7]?n�?��g>�ؿ��yI�Eʒ�C=��>��>��<?��>M�P���p��T��h@���2����>iyU?����V��G>�7.?�oܽu�)�K��>f^�=g,�rt��J��d�T>�\'?,=C�%>��� �6�����4��:*?<�	?q����<+�x��>��#?�r�>���>�<�?�/�>��þ�p�:s<?��Y?�)F?{MA?�'�>�>=�ý��ɽ!�N�$=*��>4�W>_�|=)�=�H��_�A���[=��=༊滽���;�j����<�-=$�3>r�y�E�R
Ⱦ���\l̾kz��I�J����B����ٽՖ��������k���zս2u�5�{����ؽ�����?�~�?�j���6K��������ǁ��l$�>�9��W���B��b�>�sc���W��[ ��K<�6�`�$�j�1�'?����ݽǿ񰡿�:ܾ'! ?�A ?=�y?��#�"���8�/� >%B�<,����뾴��� �οE����^?���>��0����>ĥ�>!�X>�Hq>x���螾 3�<��?E�-?��>��r�(�ɿ^���p¤<���?.�@�
B?l�(�����7=}��>�
?��=>��-��j�@I��"�>���?^g�?�f=�OX���~g?��<�lG�c ��,�=�Ԩ=�
=��xH>��>�����D���ֽ�+9>K��>g�5�`����_�Ͽ</�Y>�ǽ�����w?lcx�_+j���ϾI�J�13�<��t?���=7�W=�eF?�	?���ѿ�iE�\;�?�1�?�I�?�?���}e�>���5��?CZ??*�?>����J���,���Ly�<�t��W۾5O���<�>��>/�M��=YM��#��#�=]�=�&�#iƿty$�����=�E��P]�:~轮���T�c����-p�~��o�h=C��=��O>i�>�U>��W>�W?k?oֽ>�>�]�o��
˾��YR���a�$���E���9����R���R	�Lq��n��Cʾ~2=�y�=�/R�\����� ��b���F�i�.?�#$>_�ʾƵM� �+<�cʾ'���Eم���k1̾ޚ1��*n��ʟ?O�A?��j�V���3��p����W?�v�]���֬�}��==밼+�=�(�>���=����&3�y�S���0?��?����-����)*>�A��fU=�
+??~8�<봩>gW%?�c*�����!S>(�7>�ҧ>2$�>��>�I��vҽ�=?9�T?�x�(ɟ��?�>�ӽ�%�}�0�X=
>!2�����DZ>F5S<Bp��O�f�	��"��<��V?檐>�9$�g3�����,�~��ۼ,r{?$?|O�>RNs?#H?��Z=I�����W�:}�Դi<4�N?�eo?̹>�?�t��m��Y�6?�Cq?"�2>(0f�2��3��G���?�yt?��!?�k�<&H~��Ƒ�>'�	?7?8�v?�X�I:��m��fE-���>��>Z$�>&���>�%?�q���s��G�����A��z�?�@���?�����{��D��=��?v��>;_��+�G��PW��´0�*��>�o�o�W�3�\�(�x�?%t?ɷ�>������羨��=oٕ��Z�?d�?a����5g<\��~l��m��ʄ�<}ѫ=:��K"�Z��%�7�X�ƾ$�
������ῼq��>5Z@�S�L*�>D8�P6� TϿ����\о�Tq��?怪>��Ƚ�����j��Pu�ɳG�&�H�����i�>:�>ڏ���ޑ���{�\�;�����`�>��U�>gT�0�����89<�Ւ>7��>���>�������쮙?u���53ο>Ğ�7��ЯX?�Y�?Y�?��?8<D<��v���{�nX�>�F?gs?�Z?��$��Y]�,Y7�1�j?�_��U`��4��GE��U>k"3?B�>�-���|=$>ӊ�>f>R$/�x�Ŀ�ض��������?0��?�o꾂��>{��?�s+?�i�68���[��J�*���-�<A?�2>&�����!��/=�$Ӓ�G�
?�}0?Wx��-��GY?(q��L?����-�3�>s�>�w�?�羠�����>Z�B��{��C���ɹ?��?
V�?w�7l��f?��m>T����T�\.�>&�:>ە>��?��U����>eG��<	��:e�m��?��?��>�q���ڗ�sO;��?��>�̘?;�ӻLK$?Y��;戕��ė>���=�~ >�fk�>�5?0b�>�q<B�}��9��&q��8�O}���n�>X�a?��?^h�>j佌7�<�CS�{�y�0�j=�ħ��LԾ�n��������=���,��=ڳN����G?Uv%�>1п�?��,is���.?�*�>�?'��A�`ߐ<sTe?�~U>��汿*��BȽ�ު?��?�%?�оN齳!l=:�>��>nDƽwȯ��jx����>��)?)����Ǉ�Iu��\>���?K�@橱?�Q��Ҥ?ǣ�*��][�������t��5>k<A?���b��>���>��+>��y�4���u�yr�>�E�?���?���>��v?�rc�'�H�^��=��?L�_?�@�>W>ʽנǾE9�>��> ��叿F��gTy?�~@~�@��B?�ک��hֿ����^N��P�����=���=Ն2>�ٽ,_�=��7=��8�>=�����=s�>��d> q>:(O>}a;>��)>���Q�!�r��\���S�C�������Z�C��Xv�Wz��3�������?���3ýy���Q�2&�)?`�ݕ<�\y?z_?�g?��?o��,�>��	�Y]_��G}���t=�_>/!-?�=?ǰ$?D_p�����:�f�6`y���оF��-��>�z8>`�?��>햖>�,��eUH>��~>B_>>>��<5�����<W�D>+�>� �>d�>uC<>��>Dϴ��1��j�h��
w�k̽/�?����P�J��1���9��Ϧ���h�=Eb.?|>���?пd����2H?+���w)���+���>�0?�cW?,�>��n�T�%:>;����j�5`>�+ ��l���)��%Q>{l?�f>�1u>��3��\8�/�P��n���`|>6?綾x^9���u�P�H�hݾ�5M>�̾>M C�h�O���L��i�2u{=�~:?�~?�,��.ް�5�u��/��jAR>�J\>I=Ku�=>\M>��c��1ǽpH�x-.=���=��^>Ĉ?��$>�Q�=��>� ���ZF��e�>+BB>�;>��@?�#?��F���?��]u9��}>�<�>'Ǉ>���=��K��-�=v��>4Of>E���������h>��M>���7\S�ϡb�h�J="������=��=���Q%2��1=�}?�$��NW��Z"�vg�c^D?9�?�%=)�R<���v��WcϾ+��?�@YI�?�����S��9?�?"v�����=�F�>���>�rھ�EX���	?'��^`��sJ
�\�)����?��?��0��H���i�T�>�f?��̾� �>E?W�����⏿�y��$=8�>2QT?����:���:3?��>��˾����Ͽz�p�#��>��?��?��^��p��T�Q�:=�>s�?'�K?��w>�O߾����>�"I?��9?L��>���k=ؽ��,?��?]Tl?�I>���?T�s?Pk�>7x��Z/��6������Ep=�[;�e�>KX>@����gF��ד�oh��Y�j���%�a>��$=b�>PF佢3���7�=%񋽘H��Դf�٥�>�,q>j�I>wW�>�� ?�a�>��>�r=�p��‾ⷖ��@F?��?{���I��<-ݺ=:6ѽtB+?��1?ב}��z��p��>`�p?IIu?�U?>�|������I�����.�=��>z�? �>�{=��h>پ� T���></�>ۏ��w����˾�ݼ���>�5'?6{>m��K}#?e7?'�>�ª>��L�
"����`����>��>C�?���?�z(?���/>��f��Kϥ��ib�HM>�?n�?^�>}���O����=�� >ѽ��q?<pA?�J5��m�>��w?(�T?F?}ϋ>���_�[���ү>h�!?�S���A��%�\�6�?�B?���>&��)Hн�Լ� �����3?�\?�r&?�q��`�+���E�<��Yh7��%<b���%>�Z>�x�ʍ�=�@>N�=��k�~�6��GV<D�=�ԑ>
@�=I�8�2����2?�<�C�S�Ld�=5�a���8��K>��I>1u�=_?�`���R�ܺ���i�����⽈?m��?R�?*���[���I?$Ή?~[?�>�W�cb��+f�����z��������	�=Me{> ��<Zf߾�j������rAo��L����+��h?6?��>���>aBh>w{�>��Ⱦ����������l�c_�-�,��V�D���p��
C����:Yʾ	!��
 �>m��ʢ>�k�>�n_>zF�>�@�>EÄ=a�>�s>��>��>>֌=ƍ>���=-u⻃���FR?�����'�^v��p��B?�pd?h�>Ӹf�#���ܨ��r?y��?�y�?�v>�Wh�zA+�2 ?p��>�C���f
?��:=��#�<�,��P���[�������>�ٽ�9�6M�2�f��u
?�J?ɭ��l�̾�aؽ1�����n=�L�?��(?��)���Q���o�/�W�NS�v��|2h�i����$���p��돿�^���$��Т(��k*=��*?I�?O�����!���"k��?�$lf>��>�#�>۾>qI>��	�j�1�T^�&N'�����gR�>]{?��>��I?�<?�vP?jL?x��>�c�>'7��Bj�>�b�;d��>���>��9?
�-?�70?�y?�r+?.c>xz��B��l�ؾ�?�?J?�?�?*܅��uýU5��ٗf��y�x����=���<k�׽4Cu���T=b	T>�k?���8������2k>�7?�Z�>;��>+Z��ȸ���p�<\�>�
?���>� ��8r�������>lw�?q�g�=�)>M��=�8��I���<��=�¼��=I� �9���#<���=���=F�{�������:��;�/�<�]?߉?���>�3�>���v��8&���>2��>���>ﱯ>H�e��N��o���aۃ���M>���?�N�?�%E=�1�;ƒ>KZ�#b��+��(0��(g�*.?߳�>��?���?�e?f�?k>>;��X���Ђ��ո��^!?`!,?<��>t��s�ʾ�񨿬�3�՝?E[?w<a�����;)��¾�Խ��>�[/�?/~����DD�P����<��(��?ݿ�?RA�?�6��x�̿���[��t�C?("�>�X�>e�>M�)���g�l%��1;>֊�>ER?�#�>h�O?�<{?��[?�gT>8�8�]1���ә�mF3�`�!>6@?���?��?Wy?�t�>^�>W�)���>T��=���	ႾW=�Z>,��>�(�>0�>���=� ȽTY��g�>�Xa�=�b>$��>��>��>S�w>KL�<ĿO?�]�=Ծ��+��6>�ڊ(���/���e?��?�$?K?���|⾗�%��e��8,�ﴚ?���?i�??Sؾ:s	>�S��9
��b���*�h>
N?���>�ܽ&B>��>V��>�.�>~I>%�6���D�.x��!�? �?N�<p?ڿI=�y�A�@M<�'�����$��A7�Q��ѿ�+��=-1˽�i�+i���ŀh�Q���L�߾����I�*?G��i=��-> ^L�.;-=��[=�G�=�H����Q=ږ�Y=B�<
���Mn��˽���<�z4��
#>�����?�;e?7/?<yU?�>>ċ>���pz>U"�� 	?�?W>�D<t碾�����Ǿ���/��	�˾��� e���܂>�̼`��>$�d>I��=/��� >��>���=�N�=��H;�Ɉ;a()=W�>U�=�/>�e>[j?�*���׬�B�h�i�A>�Y>?�">a�= ���Si?��=1�a������.�i�w?�:�?[6�?�?F�[�!ƣ>T�޾y8	��NE>� h>��=_�=X޾h6�>z8>;
�)7�� ���-��?_�@�nH?8I��,̿>��=��9>��>��R�Ƴ1���Z�
N_��%Z��p!?��9��iʾ�7�>�z�=,�ݾ>�ǾE$=��7>"u=����|\��==v���9=u�k=���>7�D>H��=����
��=u�N=���=o�P>VT��]k:���,�E�3=pB�=�ec>�&>��>d��>��&?/�?���>��������"�G�>p9�<��=7��<����}�>��F?�J?�9^?�d�>�c���>I�>�:�א��)@t� ��X�<.<�?i��?�z�>*ge��x ���F�����jA�H?��?4�?u�>5V��࿞U&���.�vl���E��<�*=
lr��AU�����um�H�����=:m�>���>���>Hy>z�9>��N>�#�>̙>���<瞅=����YQ�<���ݤ�=<���oQ�<��ļ�֍��"�[�+��%��5�;f؆;�'^<��;�4�=_$�>_>��>��=���w!/>^_����L��~�=:��2`B��/d��~���.��5�m]B>�~W>��	5����?r�[>��>>V�?�t?%�>z���վA��Cd�W^S��¸=�	>�>>�Ss;�dI`���M���Ҿ���>��>��>�l>3,�"?���w=�⾳a5���>]{��m���&��8q�c?������i���Ժ��D?G��ӥ�=�#~?-�I?;�?���>a����ؾ70>�E��B�=��(q�=a����?W'?J��>쾃�D��=̾<��z��>m1J��
P����0�W��D$�����>�˪�]yо�3��I��������B��er���>��O?���?Rb��Z���\O�����9���]?�cg?�>�k?�(?s��g�%���|�=i�n?���?LL�?�G
>�������<J?k��>"v�?�u�?��r?Vu����>�����K>{�e=/2�>EUV<�G`=7�<	��>2d�>��?�sA=Y�0��V%�H��Q�i���j�*��L>�̈́>N�e>(<�>��A>�FP>M�>�י>%ӥ>1EG>��>&t>����X��uP?�>(�>4�;?���>p��kY���F���&l�<U3�3_����EY�
�<�M����=��u=�@�>�g��f?���>������>o5��v��;��>a�>"��=u��>/�>;~>nކ>Q�>
�m>p1�>XW>����Ǽ�4꾉���7G�E	<����|�>�徬����Ծ/𩽾�<�LI��5T ��〿7.p�b?G��iD>�}�?ێ{�g�B���O�<G<���?��>/V?�b��0S�<AyC=���>sD�=���
��Hd��	�ǾhÕ?��? �Z>��>#�d?�H?h8���
�Q���d�8�M�S��d��҈��`�Z���28ż_?Z�x?��5?�]>=iµ>jW?��:������>�>�;6�`8J�V�l>�>Z��Rud��	��\^�O��#K�>/_?���?�)?f��a<���g$>99@?��'?IOx?r�5?�Y2?�h���?�>qb?�S?7~A?�#%?�>?��>�QL=�-�;g�=O}¼nY��N}��8��_�J�h�
<��<d�B���A�ݚ�=��=a���̴�'Fa<Z:~��P�;8��<���=���=p`�>F�\?�R�>	��>��7?p���,8��$���/?��@=E��̃���6������ >��j?��?��Z?��a>�A��A��J>[%�>��%>�[> ;�>����E��a�=e�>g�>��=��N�r��%�	��w�����<�>���>��>�a�<L�<>p���B��!�=>��d�Ͼ����C\��R�N�LI��e�?��?l�7?<��=󪾾�|>O��ްH?�M?�/?R?�O�>���>.��Y��	�#�>/B��n�,s��\���&0�2g��M�{=�]�������x[>?9
��]ܾ_�m��iK����+3=j$���L=g�	��<ԾP�|����=�?>n���r^ �O��.p��,\K?:tS=���frS� �����>[ڗ>w�>9~:�o|h���=�BM��.h�=�f�>ڄ;>6]��g�gF���EB�>�DE?OO_?�j�?%6���s���B�����}|���Dȼ��?zU�>Nk?
fB>�w�=W���`��*�d�kG�� �>o��>,��C�G�%$���?��6�$��u�>f8?�>z�?��R?u�
?Ǧ`?�*?�@?��>	|�������O&?q�?:x=�0ؽ�4V�N^8���D����>hd)?R:D�(��>?6?V�?�2(?#nR?$�?q%>I��A>����>�ڋ>Q�X�aI����a>�K?��>E�Z?��?��<>��4�X�������7r�=�>>Ac4?�^"?d?���>���>2���$�=���>oc?�0�?��o?��=��?�72>]��>o��=U��>��>�?WO?$�s?��J?���>���<�<��^;��	Ds���O��ʂ;1`H<;�y=3��*2t�0@����<�;ea���D����񼷾D�������;�K�>�[>�m����7>��о�搾�CY>�㥼$˞��
��E�M�[?E=�w�>B:?:ʣ>L`
��͊=���>��>�h �:�.?��?4�?<ʼ��^�4�� N���>��9?+�=��c���Wq�3w�=��k?�4_?�P@�ٚ�GUR?��h?`��5IH�6�۾@h���(��=?mg�>���>�>���?�w?��?����Y���m��4u������_(���?v��E�c�qrI>�g;?Q6?ąB>��>��:�Aǝ�Mgܾ�C!?u�?�B�?��`?�)>��L�X@����VJ��X^?�~�>A��$�"?� ���ϾHS��9+��5⾱��c��[@���v��>�$��܃�׽��=M�?Xs?i[q?��_?_� ��d�q.^����8jV��%�W#���E��&E���C��n� b��.�����xRG=P�=��1��U�?�x?gX��y�>�᧾���!1�<�>c@̾���v��=�H<�P>���=K+�6�2���=���?� >�5�>7-Q?2�>���l�i����I�YZ���>D��>4�>���>�>Q������\��˾J%I��4v>�yc?F�K?��n?!q�a)1�S���`�!���/�"i����B>�f>뻉>(�W�Ɯ��9&��Y>���r�	��{��o�	�q�~=3�2?�+�>���>�O�?L?�z	��j��Mix�9�1����<�1�>�i?�<�>��>��Ͻb� �B��>��l?��>?��>$��;r!���{�+̽@(�>�s�>���>o>�-�VA\��f��~o����8�)8�=�sh?����s`���>�R?���:�lK<��>J�s�y�!�	}���&��{>�^?i��=dD;>Z�žw�no{��!����'?�?Ď���*�mh>#?��>g�>��?��>u�̾6����?I[?0K?�:@?g��>��v=,���|I˽�/��uL=���>�R>ݧ`=(#�=H
���^�}���Kz=d��=�f弽����;'O弰��<	�<��.>���:2G�m*��ߕ��A�f(�����f�'�����BB�+a��~�$
�����u��3�X�r�Z���k*b��v�?-��?5:��n7�>�����f�5�>l{��5"�A���@`��;��ַ�Aھ����jE�ͬi��v��K�'?�����ǿ𰡿�:ܾ,! ?�A ??�y?��0�"���8�� >fC�<L-����뾮����ο=�����^?���>���/��T��>٥�>�X>�Hq>����螾�1�<��?;�-?��>ώr�/�ɿ_���ä<���?.�@��A?*�(�{��O�N=s��>љ	?�y:>�.�C���:�����>D�?W9�?�3=ayX���m�f?�S9<��G��u	�+[�=�)�=��=s��`�K>���>t(�iVE���߽sd8>��>&J&�h��a��C�<��a>z�Ž#���[�?8�^��?^�@���~��T*Լ�Jf?�~�>.�
=��+?%�?�/1ҿ)�%���e?��?�{�?�?�@��#��>���80}?��K?��">y$G�><q��������'�#�f	ľy�r�}��>D��>oΪ=EƖ�!�ʾ�j#����=���=���w�ÿ�H� U(��C=.۔�Ž̋$�^�ǽ�Dս���l�E��o��֯=. �=u^@>�>��C> �>^k?7�?���>c�'>�Ƚ�\��rľu{ �� ����"�s�l��p��о<�龝����7�a��f?���z-=�s<�=�R������ ���b��F���.?f$>��ʾ�M�u,<Xjʾ���^]���b��S-̾��1�n�E֟?�A?煿v�V��	�����B�W?86����ʬ�(�=A~���"=�>��=Q��J 3��[S��20??�;��=�&>�����
=�+?$� ?�8<��>}�#?�_+�W0�e]>�H4>r��>C�>A�>'򮾿Y޽��?oT?��R��I�>ȇ��h!{��h=�D	>��3�L \>�<?/��2�I����ڸ<�&W? ��>��)�t���~��~b!��5=y�x?��?�>�k?~;C?;�<.y����S��V�j�r=�nW?�i?Y>��H�о�0����5?��e?A�M>|	i��I���.�'��o;?��n?ą?�Ǣ�D}��7��u'��D6?��y?.MO�n֗�iM�H/�O��>ʓ�>�x?u��3��>��4?����ď�:�ÿ�Z;���?#M@���?厙�b�Z�s�=���>�&�>�M��c����%=�=s��`�v�><�����K�HD�N����A?�HP?���>I#�0�ɾ���=�ٕ��Z�?��?~���gDg<R���l��n��a�<�Ϋ=���E"������7���ƾ��
�����࿼̥�>EZ@�U�w*�>�C8�\6�TϿ)���[о~Sq���?L��>S�Ƚ����A�j��Pu�b�G�3�H�ť���>��=���� ���nq�w%2����<��>� ���3C>�Ϛ�
aо8���qw>��>�?) �>���L�]�a�?d�����пز��`sϾ�/n?��?m�?=�c?%����Yo�Eѽ��+����>S�Q?S|?"Ռ��}����l�%�j?�_��xU`���4�uHE��U>�"3?�B�>T�-�c�|=�>���>g>�#/�y�Ŀ�ٶ�>���Z��?��?�o���>r��?ts+?�i�8���[����*�=�+��<A?�2>���I�!�C0=�UҒ�¼
?V~0?{�f.��]?��t��x��?ᾒ+／X>�򽘸;b��$8>lR��@��k[��ٶ?s��?&�?ꔝ�4��^!#?�M�>�ī��f���Ob>�d�>��>�"�>��1�=ެ>���1N2��O�=�P�?<��?���>�#��o��T8����?,��>���?JD.=B��>�'�;wV^��2�=O�g>܆>�m���]�>Z�'?r^�>���<9
ֽ!���]��i�i�E��rf����=q?�1V?mƅ>�����e�;���#t(���y��*>⍛���ý�M��L�>��o>��>lZ,����Z�?@& ��
׿����O/�Y�/?��{>��	?�)�ٗg���;�_?&G�>�@����������S��ZG�?���?�@?-�վ�)���=���>F��>"�ƽz����C��E>
�A?U��@����(o��ɂ>g��?��@�$�?�	h���?����Ո���������z��m�=�6�?�4�S��><<?[]>�k�T����Ft�J�>B��?,��?sj�>oz?3ZU�SVc���?t7L?���>�����H� ٨>��>z��d
��/�:�r?I@t�@��C?����hֿ����]N��M�����=���=φ2>�ٽ_�=��7=^�8�R=�����=t�>��d>q>7(O>va;>�)>���P�!�
r��[���T�C�������Z�B��Xv�Wz��3�������?���3ýy���Q�2&�?`�#��=Pb?!M?`?_c�>b�<�Ms>e㾇�0=�����u�=ޙR>�O*?	J6?$�?:H	<�#��.�b�"�~�,zԾ*��Γ�>|�4>�<�>���>�A�>&%��^�`>ޅP>y�c>�>�j=>dJ=$��+
>�+�>���>�ڷ>�C<>�><ϴ��1��U�h�o
w�̽�?����[�J��1��}9�������j�=Fb.?f|>��� ?пO����2H?����X)��+���>w�0?xcW?i�>?��c�T�,:>ÿ�0�j�Y^>^+ ��}l���)��%Q>*l?Bhf>wx>�Z3��18�n�P�������|>�6?l@����<��^u�l2H�Heܾ��L>�y�>c?R��������t��>2l�*dw=��:?�?ң��Yu���t��ӝ��Q>�Z>A� =�q�={L>�i�'�Ž��F��.=���=��`>�D?T�,>�ُ=_,�>󯛾�Q�7f�>�q@>�(>�*??>�$?tV�����A^���0.�$v>���>{Ӂ>,>SRK�~��=ܤ�>��c>_� ��W������>�)�T>$�x�M�\��u��x=̔��A�= ͏=����l!=��#= C~?$I�� ꉿ�!������4?	4?�p
=YZs='a��kN��4�;T�?��@�?�㺾�d�BZ�>��?���b>Ĉ�>vڲ>8�.���ž@�>?�ϊ=�N���3�q�Ѽ9��?+p�?`�1�����M�Ո�=n�?�L¾5Y�>��T�/�������u�7��aș>�ma?����o���ܽ� ??�5�����ȿ)zm����>�k�?���?�`��l���sR����>�	�?��I?m��>�̾�(�7�>�J?W�I?�%�>= �����{�!?"[�?��?�I>팑?�s?E|�>�mx��[/�M5��W���f�~=Y�Z;4l�>L>�����hF��ד��g��#�j�x��s�a>Ó$=��>�3佦3���T�=�����O���bf�J��>2=q>��I>�\�>�� ?�b�>���>�/=�~��Dှ������??��?CH�g�y���g�=�%�ņ�>˲/?օ%�N#��;�>��b?�ہ?':?0h>�� ��:jο�8޾բ�=�>7��>�#�>�Խ�Ė�>�?��S<��y^>�O�>6���?����4{;>�[�>�h�>��>���<2�%?��?b�V>u��>v@����Vn�0E�>�U�>�z?���?��/?���d9��G�����{�G�L�>��\?�3?��d>�l������<=Hu==4�}���P?}�~?+�w��>�7�?oJJ?@�D?˃�=�hT�V�?��᛾ +�>h�!?$y��'A�fM&����L�?��?���>�O��K�ٽ�����U���?�D\?&#&?�O���_�^#��~x�<��>��� ��7<YQ���>V�>暊��p�=��>x�=Al�VZ6��Ot<�	�=���>�B�=��7�t���;?BQռQ�Y��K>��j��lf��d�=Zʣ>�n1�J?q&>���׶��ߜ�
x��w?s��?�9�?5�ƽ��r�9T?�x?�;?֍V=�/Ծ[wþ��ӣ�m����/�F��h�>��޻����ݧ��=��(:��p��<;i �ő?[�>�
?���>c�[>�ӻ>���g!�C������j\����}p2��7(��襩���4���g�G�վq�}�}��>phv�j/�>��
?�v{>�L>7��>�w�<��>�2I>=|>}�>g3>��>�2>�&>=����:9T?�۾�5*�|¾3�Q1?!r?i��>�"�sYw��������>1/�?��?���>��U��*�|��>?�@~���?�N�=г�X�ӽ�z�>.��wC�����B�r>ءͽg�2��U�̀m�4~ ?�?܍=�p����d����Rn=�H�?��(?��)���Q�ݺo��W�S�`���h�g��.�$��p��揿]���!���(��)=ʘ*?�?�������0���k�c
?��f> ��>�)�>ھ>eVI>9�	��1�o�]��O'�����W�>ZW{?ek�>��I?�;?imP?�^L?�̎>s��>���8[�>��;t��>g��>֘9?��-?�#0?�_?�O+?�b>����i&��Ҁؾ�?͗?�Y?�?^�?9����ý<,���g���y��I��%|�=?��<�ؽ��t�� V=<T>? ��7�7�����(f>>�7?`��>�y�>ِ��`��d�<��>
?\n�>s���8xq� ��~7�>Ă?���n�<6+>J��=?v��E��$��=�iμ��=�iQ�9o.�GD1<ӡ�=
�=��H�ͺ��?;�24;��<�X?�k?|��>���>VF��DL��=�v��=�b<�@>�2�>dfǾM���ߗ�<Gk�S�>WP�?�֪?y=���="K=x�s���̾>�Ѿ�|Ǿ��뽩?H�(?� _?�q�?	U?�	?X�:>�9�k��������H��q�	?,?��>���I�ʾ���3�G�?Z?�9a���/>)��¾2�Խ�>�S/��(~����D��m��������ۙ�?S��?�A�n�6��u�K���+\��\�C?O(�>�S�>��>>�)�,�g�#��4;>��>�	R?y8�>�zO?�z?l�[?��R>��8�z쭿뙿,kQ���!>��??�P�?��?��y?�M�>�6>3�(��߾n���N���)���J�R=B&[>�!�>h��>х�>�#�=Y>Ƚ����n>�	e�=�@d>�g�>8��>��>Ԑu>鲲<��^?^�)>V���
�(��rO�Tᴾ��?T�?��@?��þ�1c���׾V�0�X�>��?�}�?�y?�
����==D �C��cn���>�>������=T�F=���>C��>�T�>$U�<��L��z���G8��U[?aM�?��t�Msɿ&cH�[�j�������%� ��P���~������|��:�!��g��lӽ����LԱ���ξe� �^
���5??��N��Q(+>��
���u�n�޼�x�=��{���>���=v$S�l�;IU�=�>=.f���^��`��6�@=�]�x��?
T�?�u8?���?�8X?g:>?f�˾��>�ಾ'�>���>��D�F���[�ޞ���}�����w�� �����f�=(��.>aW>��<t��tY�=z h>��L=�k�=��%��Ѓ<���=1�)=̴>�lN>�Xk>��s?Sȉ��
��{�t�~��=��?A�'>D	l>=����r?3@k>Y�i�"��P�
���t?s��?Lc�?�f?�~�G��>��˾=�tb�>D��=���>\>��쾉��>��l>�8�Uϭ�)�x��D�?g�@؏N?\���mͿe�8>�7>9>.R��1�Ir_��_��[��R!?PS;��;ƃ>ۯ=�
߾�qƾT~8=�*7>X9b=o ���Z�;l�=����{hA=>�p=��>�'C>���=�P��+��=��R=M6�=�P>w����3��0�?�.=D'�=Z#a>O0%>�b�>E�?�f?Q X?)|�>�}��aw���Tݾ]�_>���=*�>�A�J:X>��?S�G?_�D?ߴD?/�>���=ֈ�>��>��@�'�x�����XX�w���b~�?���?���>��b�)��H�*��9@�`ν�#?7�?�)�>���>i���� ��6����I':!�<�!���eO�]�j�� �WBɽt�%>gK�>�*�>���>�iw>k�=>pς>���>C?A>�4<R �=��&=�=P���ܝT=��������g��[F<��%��7-�[^���L)�I�"<L���f��]�(>k��>xd>�?G����R۾��=�����aY��6=+xZ��{9�r�n�y�����5���A�\+�>�g|>B�\� )��_?�ȁ>[�>��?�og?���=}j��~�ԃ��Ym�zC��y3�=T�> �3�ȲA���K�ȹD�s�����>���>��>C�l>w,�>$?���w=���c5�)�>�w�����S4�\:q�z>����5i��VκP�D?G�����=!!~?Y�I?5��?Ԏ�>�$����ؾ]0>L��0�=�&#q��`����?
'?���>���D�N����CS�>�p��9�P�����1����=P-��M�>��a����#�g���4���	L��i���>.�O?N�?�bZ������/\����*y�0?u�d?�C�>-?#�?�u�WP�\݉��P=��t?Y�?]��?�f�=w޲=o�����>	�	?P�?[ޑ?��s?�]B�	��>�b;�F!>!����=�>�=uL�=�
?V:
?2?hJ��K�
�����񾑻]���<�r�=���>_�>��q>���=2q=Bw�=�Y>���>>W�>v�d>q'�>��>����V�
��%?+�={�>s�/?�p>m�N=�\ɽ�2q<�(��;qW��*.�����2�����<�
��tx�=r3#�Xd�> ǿ��?#=_>��.k?���.�
�F>�(e>�����N�>�9D>S��>���>zt�>��>�f�>��>�~��zɽV(޾[�8�D�j�\�W�׾
k�>C�˾y����F�w���^j�č�~���w�yj���6�`��;��?
����[�>e@�p�z����>a>p,k?�sJ����<�$>�=�>�@�>.f�<L���6���J����?N�?U"c>8�>�V?ю?zC��'��ZZ���r�� B��*d���b��'���n������X��e�^?tRv?uC?`�=\�y>��x?�#�9o�����>�\2���7���=1��>�K��|vL�`"˾V����`��7H>�l?�ȃ?@?%�\�����|i>Y
J?�N4?6��?$sD?��C?��g��?�.�=nG?��?6�?8?�2�>�8�<� =t�<"0 >�7������6����e�.��M�<;��<cy��t;��g};��j=��`=�e;J:�;�;���r=z=w�=+��=wɤ>�lX?	��>��s>��(?����+8�?���Ծ$?�݀<�6���I��4���P��>3�g?cy�?�0`?��>4KC���S���)>-�>�!>0�Q>X&�>x���IL��S�=��'>1>蝓=�r������A	�����IO<��>�]�>��6>j��)�=iH���}�֘\>��B��O �6(n�������\�~�4��@�>D��?U�7?U4�=�ɽˊm>�h��!==?Q�(?2~�>�fL?�C�>�.�%����"�}�r�>�~	�<5�K��灿��!�9o#;��>��8�B����u>���¾q��L�E%�2cg=XX�DA ��/���3ھ���r>� >�ٽ�gp!�����1�W�E?]��=�?��U���l)��Vh>3��>A��>[u�U�ܽ$�>��@��J��=��>��!>M�<��Ѿ��U��B���>{P6?��[?_x�?�R��V�o�V�P�ɡ��K����C��N2?t�>���>.�y>|6>�Aξ��$���\���M�#d�>���>P�*�o8N��+����ɾ�$Ծ�P�>�[!>>%�<���>`,?��>.�R?�l4?��?&�>/���+��'"?4|?�?"=6�R�7Ѵ��4�"9�xr�>���>� ���>���>
r?/?ֱG?5:
?}~>Y�S�W쀿$ �>e��>}9����G�>�[?��>t�*?�HE?ף�>���QW����p=Q���-f(�QM?)�?�p?[�j>�M�>hM��Tx>�p�>�iC?�%u?�j?,�=�i;? ?3ԅ=	<����>E��>{�,?�	X?��@?m�D?3��>���<gqսY^���@�!�[jF<q$d��
���������WҼ�,�=.�߼���-r=|#`<u =2�K;M'8+��>�W>�+��R�>�����@J��q>������B�f��E.��W�=Xz�>3�
?��>����i=#��>��>�^$?�4?u�?�g��c���þ��К�>��E?��>�e��ޗ�ӆs�I_3=�1k?��d?h�j���=b?�P^?���:�|ƾ'@j��?�NM?�	?��J��Y�>'�~?�p?�o�>oi��m�@���a���n����=
��>���e�8�>b�6?M��>�s]>�`�=H�ھ��v� 6���z?���?ݯ?�?
�%>Yp���߿���(T��`-Y?���>�û��?
$������t���i��ܾZ���J���:�����0�Lc��d@�vt�=��?�=c?��x?�d?L���p��h�������b���㾫7�oJ>��:�/�B���p�H��|b��4��K�pZ��G����?-$?1]�S��>�����ɾ�;��^>L�����"�.@==dű��>�:�h=TP?�)˽����M;!?ʿ�>q��>��@?�a�&L�i#>��lJ��N�c�q>��>e%�>���>9�X���V�n��")׾�7�����z��>�r?��\?<�h?�8��w��*����_��ʽ�=
�P��>GS$>���>��=�I���x�r�x���p�9��h�������;�5?r�3>���>.r�?� ?�����쾛�:�O
&�;U�=�̛>�Ŗ?���>�I[>�������C��>��l?�L�>Q��>����%!��{���Ƚ���>�2�>&��>��p>X{,��C\�'f�������9��!�=��h?-����8a�ER�>�/R?X�:�_D<�`�>i7u��i!����P;'�_�>�|?b�=y<>��ľ���W�{��B���Z&?�&�>�����I��>ϴ#?���>m˃>�˂?O�>�ٯ�8@R=%'?�Qa?��L?]LA?�E�>�� >Uk��%7彲#�,�|=@�d>�jS>aj=���=�a�2�^�#Z$�D��<F��=xۄ�G!|�f�<qQ=x��<S�<WD!>6rӿbvO���(���־�-�v���m�Z����x� ��sھ9������LZ%�x𮽄BM���+��g��C7v�i;�?��?tKC�Af������~�����B�>��Xx��?UӾ xB�S¾g�������&�#�[��s��Ol���%?6���iƿI㤿��־��?e�?�*z?�z�i> �e�F�>�b�;��z���������ҿj+��,f?D��>���5�@0�>�s>fu>�(s>��z�n;��v��H%�>�|3?i5	?��v�>BǿzԺ���x<5��? �	@�oA?�(�Ӳ�IW=.��>[�	?v�?>2�L �*İ�X�>XR�?��?G�P=�oW��	�}e?x�<;�F���t��=�o�=ҍ=o��qYJ>�?�>�U��EA�dHܽF4>م>q*���jq^��м<]]>+ս� ��5Մ?){\��f���/��T��U>��T?�*�>W:�=��,?W7H�`}Ͽ�\��*a?�0�?���?%�(?7ۿ��ؚ>��ܾ��M?aD6?���>�d&��t���=�6����{���&V�~��=V��>i�>��,�ދ���O��I��Q��=���L�ȿG�H�W\)���!>jZ%�4I�oC���&����8���)��S���=ݹ<�cn>���>�{>F�?>bdu?;+Y?ku>�l#>��1<���j����K->k&e�{�t�l��|��wu ����=$�����})�O����4�V^=xJN�����_��?�t���P��0?�g�=}gľ�k�����%�	˾�Iֽ�Iʽ��̾n�E�S�l�:��?�f?w%C��LX�Z���a�f:��rG?�U��u��#R����=�U�����9.o>V����u�B�?gH��*?=90?�q��:�b�L2�>&DӽI��='�!?R��>�T<�3�>P�><�A��Sg�6<}>��n>�c�>��>�|���؝�<-z�w/:?�>m?B[����.5�>�C����<A��;�1=��ý��2���>¤h>D'Z����Hd�<d��;�W?�s�>�)��#�Z���=���;=��v?��?A��>��k?s�C?��<�����R�.�
�@�o=��W?<i?+>.����Iо�٨��e5?P�d?YK>1
j�a�X�.��5�Z�?k�o?��?$u���}����1���06?"�v?��]��Π��O�!�[�n��>���>���>Q�:����>b�>?m#��Q���i���75����?��@�s�?�Z<nw&�Qc�=�W?���>NL���Ⱦ�I���|���O{= ��>^+��ߜv�����:-���7?���?��>����6��'J><$���v�?�?e��Ou� ;&��UK�'�����=��O> ~d=�災^T"���a�B��A[�ת�N����[>��@lc<��>��=��2ڿ8�ݿ����H��D���p?�%?�7N<,�ƾ�o�ۇ���<��<�&Y���Q�>��>8���ڑ��{��s;��N����>R���Ԉ>Y�S�G#������F8<O��>��>ß�>[ѯ�q������?AJ��s?οk������.�X?%a�?�m�?�U?�y5<*�v��{��]��G?�{s?jZ?$�$�Ę]�V�8��}p?����}6����M��b��R.>��2?�o?�LR��K�=�C,>�p�>���;l�,�PȿD��2(W��?��?HI��?�>63�?��i?!������Y��ss��~�w=y5?h��>��@}�rM����|?�??�)0�n�>�M�_?�a��p��-��ƽܡ>�0��f\��H��0��6Xe�����@y����?)^�?D�?���� #�N6%?4�>}����9Ǿ��<h��>�(�>W(N>�P_�T�u>n�j�:�;j	>���?�~�?	j?敏������V>��}?��>��?�=L�>o��="��&!��%>��=C`I���?�M?�>���=�9�P@/�LVF��R�ʬ��C��H�>(3b?��L?v�a>b����2�Ә �;�ȽD�0�]�E�?�z�)�$:ܽ*$6>f\?>�9>��D��Ҿ�z.?A��hܿ?o���ժ���(?�/W>�?v�<�����Lƾ6r�?��=`�L�CP���᝿~�&����?�8�?��?s޾�Z��;�T>���=:�m>H��=W����ൾ��>�Ċ?�tF������y���y>���?{@�x�?�N���$	?���[��%v~�B��w�6��X�=l�7?	���z>��>Y��=lpv�谪���s��+�>{J�?|�?���>6�l?fo���B��6=��>G@k?�m?'KW�^��\C>e�?���f󎿔���e?Y�
@,r@߂^?^����}ܿd֢���Ͼ�𹾍4�=1j�=.�=k.��\;u<�=5�ٽ�غ���g=�!�>�}>��>!%s>)�>r�>� ��(�"�+䣿�ݞ�DF9����ݕ����y��N����龺eھ\�þQ|����=���{P�Ǘ~���=$+1>��O?e�W?G�~?�`�>9*½�ړ=�澫�=�u�j�>GQ>��?\.<?L�#?�=�����Y�kn{��Ü�������>��[>v�>}?9�|>�bA�4
�>�(�>j>��r=wqU��t�e�<N�:<�>��?��>�<>f�>辴��*��?�h�=�w�mͽ���?����y�J��9���{���F��O=�=4.?�C>����Aп���+H?�x��F���F,��y>��0?�NW?�>�z���1S�8r>t��[oj�k� >�h �m�#�)���P>n?o�f>��u>bs3�OF8�$~P��p��`|>�6?����9���u�>�H�ZkݾvL>-��>�F;��H�����g'�2i���}=h�:?x?�c��򍰾u��?���R>��\>��=�=[�L> c��=ƽVGH���+=���=��^>g�?ۛ5>u�=8V�>�M���+E��B�>>>>m)>S�@?Z�#?70a����U[���+����>���>UY|>���=�}H����=�P�>D�s>�]Ǽ�4�������9���d>h�{�c�X�_7p�_�=����Ģ>���=���3��0=L�~?�~��]㈿P�V���mD?�)?;�=� G<��"�����G<����?	�@�l�?K�	��V���?W@�?�����=i|�>uЫ>[ξ=�L�ű?��ŽqǢ���	��1#�/R�?��?��/�Tɋ�kl��1>�]%?x�Ӿ�M�>�-���kΛ��4b�,�E�k.�>R?�=�Q�	�L��?-Q�>7\*�͏����ӿL��!�>�j�?d��?X3^�X���l5���>���?YFM?X�|>��ԾMa���^>_�d?ߓZ?��{>��� H�E[?,��?|)�?��j>CQ�?�Pu?�s?K��r�T�k��}����f|=��Ƚ��>�>�U��~�A�u���!��|bb��G�5�=.��s(�>;]½�nھyBo=����2=���$P��'�>[qR>��6>��>��>�?� �>�	O>	�<��;��򂲾C�I?�=�?�m	���g�qd�<?s�=ޯd���>�?�4���V���Y�>]?]�o?7�R?-V�>�S�|����¿���~t=��:>�S�>��	?�wc���!>��Ӿ�.��'�>D(�>,O���	پ�掾7�p��Y�>��?e6�>�q>̗ ?�#?��j>O�>�qE��A���F�wn�>7t�>�6?��~?�?Ͽ���p3��������[�]`N>�x?�A?',�>ׁ��z��mF��IJ�mJ���|�?\�g?����?<4�?�??�A?;f>#v�Jؾ�����Ҁ>��!?K4���@�K�%��
�2]?��?B��>�����yν����P������2?��Z?�O&?}���a�jhž�4�<��뻺׀�!�/<P�ả_>��>J����=�>�M�=��o�։;��<,ͺ=�<�>n��=��2���L�2?�<=�&��:�<�x�)�P�kA�>x�>i���9JL?��.�m��ʬ���︾þ_?�c�?��?����ko�ʝE?�(v?��?�@?�Y����Ͼ�5ƾQC�Mq��)Y���=3D�>"2�C�ʾ%�.h�������D��>���Z?�g�>E?Ľ?7r>E�>�g��"����r���oH��9�4�D�F/���(o����"�,\�;��ľj��U��>��<1�>N'?�of>[*�>.��>���V�>Y	e>v��> 
�>�6�>�(e>�>��;��ֽ��J?�þ!���Ҿ'�{�i�M?E�Z?���>�y:��l�A�����=?+�?I��?��>ƑT��1�31?� �>U���>??�=�!ؽ�U��1��cջ��;�k�t��>E|���Y���M�U�y��{�>�?,�W=G]���нx�����w=a��?9�"?�b'��U��sq�
QQ���S�����~����}/��tr��Ï��J��"���Q�,�Di�<d)?��?��C����籾|d�U�<���Z>2��>WΘ>R��>&�Q>��|2�"�\��*�#唾���>� y?~�>��P?�I?WL?�RJ?�ߡ>Г�>���V?�L�=v��>�p�>��?��$?e�9?�?(�?�Y�=xly�]W㾢�����'?O?!?D?��?�c��E=��<����Pk�I�ս@ȑ=\U�;�4�����5
>�>xO?^y#���3��~�!��>��<?���>�>-o�+Nj�Q.=6�?��?/e�>����?f����'5�>�;�?߾H��=��1>�%(=���WP#�EZ�=%~�QeQ=�^�D8Ͻ'��<�e>���=���
ʼ���^[�:+�;u�>-�?���>�C�>�@��0� �W���f�=vY>OS>�>�Eپ�}���$��x�g��]y>�w�?�z�?ӻf=��=	��=�|��\U�����]������<�?8J#?XT?\��?o�=?Vj#?��>
+�bM���^�������?,!,?H��>���t�ʾ��3�ޝ?�[?X<a����W;)���¾��Խ߭>�[/�o/~�����D�����������A��?��?�A���6��x辑���aZ���C?"�>~Y�>��>��)���g��$�c1;>���>�R?��>��P?�Zz?�o[?'�>��>��t��@���:��C
>�C@?(5~?>1�?��x?I��>��>>[�)+߾�d ��.�c��J y����<=5=>�Ԓ>��>&ɘ>���=\�Ľ����@sT���=[��>�/�>이>���><�@>�d��V�G?�/�>^$���~�S���K��+�?��;u?�G�?҆+?}�=S���xE�GB��G7�>JW�?zث?/�)?�T��H�=ZbҼr���łp��>F{�>��>T��=[\J=��>��>��>^�N��8���K�h�?��E?o��=E�ſ+�r��tv�����t<�,��P�h��̘���[�Л=���9f��]���rU�.�+��2x��泛� �{�F(?nn�=1��=r�=��=���M��<��]=\��<=+=��x�B�<��;�y��~򛽈b޻��<:E=����Iɾ�q}?.�I?�(,?��B?G�y>}">U >��w�>C����?i[Q>ЌX��T����7�����>���� ؾ�ؾ�c�󙟾f	>�BO��P>k�7>k��='އ<�2�=��=�H�=Ra¸�x=�X�=�]�=nA�=��=�>�>�6w?V���
����4Q��Z罣�:?�8�>i{�=��ƾr@?}�>>�2������wb��-?���?�T�?>�?=ti��d�>K��u㎽�q�=J����=2>v��=z�2�T��>��J>���K��X����4�?��@��??�ዿ΢Ͽ3a/>�W>�QF>rHE��,��3
��-3�d}~��?̮?�a;��<K�>�ڻ [�Ծ2=�<Z>���=��W�)�c���=r]ؼ���<N�=�'�>r+>E��=>O���>ez�=$2�=n,>י�a��rQ�i��<|>�.u>1@`>��>�?�0?��c?���>�l�PϾ������>L��=���>`��=��B>Oҷ>��7?�D?��K?���>ɀ�=论>�"�>�G,���l��>�g�����<�t�?ʆ?�ȸ>�Q<�A�����O>��%ý+<?�21?�[?��>���n6� e,�k9�����s���n� �������;�G$<�S<��Wa=%�><�>���>Z��>Z�>["M>g�>#�>	��R=�i=A��w�� @@>����޽V��=��=2i3=�B����9�i|��S^d�D�����6>��>+�p���>�Y�=�g����R>�i޽l�Y��$i<��|�e8�(l�: ���mH��У�T>���>t��<:^���]?r��>�s>cW�? ��?rK?>�[D��gv�5Ԥ�!5�����V?>�<C�\��N.�5��-�U�&���3�>�L�>6>Ζ>���o���{
>���=�7�Fb>����<� A�ؘ���Τ�����n5f�u��<HEM?���<J�=�?�OM?�֜?M�?�D�9�ʾC&�>y^���P3��;
�ѽ�Ԉ�y<?�/?��>e���,��̾n�p��>�I���O�9���Xu0��}	������$�>9�����оF3��`�������B���q���>�O?��?��c�m��b+O��C����??�?g?���>i�?v?}ǣ�T��U���i�=4�n?=��?=�?H
>&�0>x���v��>)S?�o�?_�?�h?ҕ��%�?	\>�UB>K��;c�>�>Q>��P>��'>
L�>^E?p�?~��������e �E�2�Mw�<����=��->��t>�o>��>	)�>�A�>�O>�xF>���=�>���>���L2־-_�>��>�O�><�(?P�>�=�>����8�[��c�<)4r�EX+�{�h�X�r��ǽ}��=��>�u�=�'�>~�ٿ���?��>��h��q{>�B �[�����=�� ?�ո���+>���=�-�>]wD>'&�>w?�>���>K|O�U���W>�����Q�0�)��`��W�4�>C�E�ּu�8���}���+���+��w�"Й��k���h=�=�?��T=V|q�1�T�3��*J?L��>u.#?Ƕ��1���;;��&?��?���� �+^���N�TYv?�q@$<c>��>�W?�?ё1��3��uZ�߮u�@(A��e���`��፿✁��
���$�_?�x?�xA?dN�<�9z>5��?��%��ҏ�*�>�/��&;��?<=�+�>�)����`�S�Ӿ�þ�7��IF>��o?&%�?PY?�SV���>�G�>=�d?�5?T�b?N6a?��m?iv>\j~?]a�>���>�,�>�74?��3?�
,?���>�(�=�)�G �������������Ἐ���8;=����>S>MYf���ͼp
��j�=�D=g�3�j��=�9�=n��<M�6>�}�>��^?f�>� �>��:?�����6�����(?��_=w�m��d�����������>џi?�Ϊ?�Q?6bK>�?�_�6��5 >�ړ>'�/>�`I>���>܎ݽ'
'��~=��>);>�{f=��Z���i���)_��v��<��!>�>+�~>�?��Ya%>�e����w�bWb>B�Q��﻾�R��F�3*2�Ϻr���>�SK?\(?���='��3n��(qe�^�(?��;?�TL?���?H�=�wܾٖ9�7�I����5a�>i�<��� �������Z:�O�3;{�v>/&��ǟ����{>v����@�k�?>��߾��˼������=���꾮�����E=��=�(��K;�����g���B?�W�=�8��0d��W<��~xE>��>G߳>qT5��	���fP��g���P�='�>�D>�}='�ݾ�GL�{���C�>�D?a4\?��?93���q��L�����򲾒�<^�?���>���>>*dW=�e���X�Aa��&I��t�>�T�>����lJ�B-��>�پx��he>�(�>�>ȃ�>.$9?��?(�S?�R&?Sf?!�>8�Ǽ;Y�&?�!�?A��=�柽��a���1��-B�a��>�a?��D[�>�8
?~?�N?xK?Q7?P	>��F����>�>t�U������^>��N?<�>��W?�ǃ?T�#>HA��]�������X�=��)>!j7?m!?�?đ�>��>툾�L>2ּ>?h?��]?v�/?%�<=�@?6��>m�>����]��>���>g$??2M?W�g?%:F?��>+=c㭽����{��@`�2&���螽���:H��y�޽|ڻ��T>݇@>���<{�<K�^��{.�hk�<w�=|k�>&rt>pk���X3>�)ž�r��Ҟ>>۰������B�-�6����=1�~>�>?@�>�$�i�=G��>�~�>���]
(?�v?�?o)E;tb��ھ��M�)�>>3B?ۍ�=�$m�|d���u�W�b=��m?^?WRV�Bx��E�b?N
^?-��#�<��/ľ-�c�!X�1O?��
?�G����>�?��q?���>��f��"n�;��'b��k�9�=>b�>1f�G�d����>[7?7��>��b>�B�=��ھOyw�������?��?�+�?�?�8*>$o�������f�=?Z7�>>�l����>��;�����Ź��v�������b�`?Ⱦt���qԾ?C������-Ҽ�~>i�?/�s?k?�a}?^� �v�m�# \�tt���k�卷�a�پ�H���B��O�[ތ�V�4�L� �&�վ���z���c1�j�?+?2?������?�&���7���h��yi>��]�e�{=���=�R�ɝ�=�.�<�9������b����?��>5@�>�V?�n_�_���H�,�H����W�>��>��=�	B>$�ؽziN�n�I��߾`ke�w�����>~f?]MG?�`n?m^:�1�>�;���Ju9�oƷ�ǆ�l�r>��3>�Y�>�1��<��:���<��>w�~�*�������s켙�?q��>'�> F�?87	?���nr�8�M�CG����<MM�>�.�?{m?Xܫ>1���$����>��l?"��>�#�>����W!�~�{�G�ʽ	�>�٭>C��>V�o>W�,��$\�i��ƀ��m9���=l�h?t���`�߅>�R? �:qF<}h�>#�w�T�!���ض'���>iq?�Ū=��;>SUž����{�)T����$?�P?�f�	�^�>�{?��>+Aj>$x�?���>k㠾��I=�L?�p`?( T?�A?��>j �=	��������	����;ht>j|8>L1�<�P�:��y������+���>�'�=�R�=R-��W�=�V<�0��=|<�>��ڿ��K�,�پ���p��a���釾����Ԉ��4������{��?��F����9�/�Y�Y�g��F��U�l��-�?w��?����G���
��*����H���X�>CHw�:�r��Y����������h��^���|"�T�O�m�i���e�9�'?T����ǿ�����Pܾ�?�; ?�y?K!���"��8�� >Z��<᧞�o����=Ͽ
���Y_?c��>���纥�(��>d+�>`;Y>�>q>d݇��Ǟ���<��?Y�-?��>�Pr���ɿ`����<���?�@<TA?o�(��H���X=�7�>i�	?�8?>pj/��O�ݼ��� �>�D�?ފ?c�U=�pW����z�e?F��;�nF�9_ǻ�\�=8��=h�=�\��?L>*�>`��BB�߽J82>^n�>׵ ���$`�:c�<i�]>��ս����̄?�"\�U�e�;�/�E����>U?o�>���=�S,?�H�2�Ͽ�\���`?!�?���?�(?�r��,��>b�ܾ,bM?G6?���>u&��t��&�=HNҼr���pV�#��=Ԫ�>rT>�m+�l���N��`��_��=�����Mǿ�K/�2�(�F=�=zm=�dԼ����y�Ž�܈�h+��D���{�r��#�=�=g�>%	->���>�rb>�W?��K?%�>���>���=��Ⱦa���_�%=�Ǿh=��_���X����(��b��->���*�Է�޸���=���=G3R�Փ��� ���b�N�F�k�.?9`$>D�ʾ��M�V�*<b�ʾ~Ϊ�$���㥽
,̾}�1�$n�a˟?��A?9���M�V�?��Џ�3|���W?�D����D���=�5��V�=,&�>�m�=���� 3�yxS���*?D�%?��ƾ�ԝ�G@A>����N�=��1?9��>����R�>O''?^G���'��I3>�
>�>���>��>���e��T.&?QZ?u��=O��p/l>55���)���>W�>	1�Pn�B�>l�=gQv���`<4^a�GQ;<)W?R��>c�)���l���"��==ϱx?�?�,�>t|k?O�B?(��<�^����S�-$�}w=N�W?/+i?J�>�b��^о�{����5?��e?��N>�Xh������.�`V�2%?��n?#V?�����o}�[�����m6?��v?s^�xs�����Q�V�f=�>�[�>���>��9��k�>�>?�#��G������{Y4�#Þ?��@���?��;<��O��=�;?m\�>�O��>ƾ�z������6�q=�"�> ���ev�����Q,�f�8?ܠ�?���>��������L>>o��/ˢ?���?�<�{$L�Y�0���O��P��&r=lK.>4f�=d��5$ݾ�p?�4��~���A��)o�<��n>n�@�+"�m�?�+h��p�:�ǿ�����Ѿܣ��U?���=�h{�)L���z�m�uX@��6�k�F�>�O|>z����y;�5&r������=�=�G>�������>�X��_� ˾^�M�0��>]{�>s�>�ݥ����׃?��Ѿ?���UK��dھ�_?���?�͑?��1?�=�7q���鶾28ֽ��$?PEt?�P[?ْS�
���衽��i?P_#��J���"P���a�Q1B>�!y?SE ?UL��
�<C��>'��>�&>�z��%ǿ\Y��{ɐ�ף�?۹�?kN��L��>�Ι?��<?�-ƾG��h�z����}0>�w?~Ē>������!< �LR��K?o?zd-�����_?��a���p�G�-���ƽQҡ>۷0��<\�p�����v^e����Dy���?�\�?R�?����#�?,%?��>����# ǾF��<1��>"�>�N>�m_�$�u>-���:��l	>��?�z�?k?G��������g>�}?h$�>C�?��=b�>�F�=&찾C.�ic#>�=�?�)�?��M?J�>{1�=�	9��/��WF��?R�� �E�C���>F�a?��L?�Hb>�?��r�2�!�E1ͽ�D1����G@�?�,��r߽_:5>_�=>�>�D�$Ӿp�1?�������]\�������� ?F��>=�?���Rs����5V?�-`>���zϷ�]���Nؗ�u�?�R�?��?��Ծ+�-�"�<�.>��>_�@>�:���'����}>}�d?��i��d��'���y>1�?�x@{ٱ?�x��	?���P���a~�r��7����=��7?T1���z>���>��=�nv�������s�a��>�B�?�{�?���>��l?m�o���B�@�1=UL�>t�k?St?	No���ͲB>�?`������WK��f?��
@|u@��^?I�Uڿ����7����Z�W��=C�>��=�aH���=���<�D�;~0�#�S>o��>�i>m��>H��>�F>�(#>+���\���٤�j����E�������_q�7G����F�G׾/�;-�V�����l=�=:�G����x��6>�X?s�_?�{?�p'?+q�=�=>ry�H��>��?���c�b>�w?��?�2??�;�>�ϗ�D�i�la|��鮾�A���X�>�K�=.��>��?"��>��˽�g�>���>���>ub�>$ͩ=_x�:�lK�>� i>)} ?��>RG<>Q�>�ʹ��0����h���v�I�˽B �?;���'�J��2���A��i����R�=�a.?C�>4��F?п�����0H?����)���+�Q�>̿0?�bW?T�>W����T��3>�����j��e>" ��}l���)�g$Q>�j?�Ǟ>�<�>F]�E��]� �����,�>~{h?)Y�	۾\ɛ�\Uh�lb���=y��>��(>퇒����?���UPy�_Wm=�!D?}"?A}0>RK�q�߾g�A�- ?�#>̬<#�|>5�>��>%>Z�ڽ𺓽�}>>�e�>�U?�5.>(\�=��>�����J��:�>8>�z%>P�??�b%?Z�������+\(�*�u>Z��>�sy>��=E�G�p��=�a�>��Y>�#��#	j��e��E���P>(�x���_��Jz���w=�"��U��=E��=n2��~>��Q=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ���>�P��R���{�b ��%��G��>NRK?��L��<x���t�>�}>������,�п�Z�����>�P�?�?�:�驩�y_�=�0>_l�?=?TW>�غ�T�{�=zY?0��?�>�(�}�h��R3?���?籓??��>�@�?��n?��?$�n�~�<��ҹ��D��������<æ�>ŉ�>礬���7��딿�8���~^��"��(�=���<���>�u"��K��^�5>�Ƚ�����5h��0�>��L>�
>̑>���>U*�>�^�>��H>�1���&��c�߾B�K?���?����n�?�<c��=g�^�2?�Q4?;7]�I�Ͼ���>�\?���?�	[?0w�>����>���忿�����<�L>=6�>�V�>�ڈ��3K>�Ծ��C���>ݗ>�Ǣ��ھ�+��W%��xJ�>WQ!?��>a!�=t� ?ؚ#?�j>�'�>\`E�|;����E����>���>*D?Y�~?��?乾�Y3�	��b硿
�[��0N>J�x?�X?ϕ>����Ճ���dG���H�钽z��?�qg?�G���?]2�?.�?? �A?�f>���
	ؾ�m��]�>�x"?�8Խ:�9�W�!��1�q�?�.?���>T��������UŽ�,�N%���>d�X?)�'?[`��¼i���۾���<����	ټi'��C<��>4K(>�H�<���=�d�=t3_=��X���V�&=��>~��>�o >��/�9��/?,?��F�탾Θ={�r��xD���>�TL>W����^?�L=�	�{�����r���-U����?���?Nm�?bӴ���h��(=?��?	?�8�>�@����޾��o?w���x��y�E�>R��>)�o�j�e���	���=J��?�Ž���i?q��>�?
�>��q>L^�>�����&�����?���Aa�ab��A��,�����m����7���Y��`¾]�s�{��>ߟ��w�>�)?V�j>+��>3E�>[��)p�>\,O>	Uj>a�>HCv>B@>g�>��%<o�)MR?������'�i�農˰��(B?�{d?�6�>�i�������3z?F��?@r�?��u>Ɇh�6"+�xx?GJ�>((���v
?��:=�	��_�<�G����t�����.w�>�t׽F:��M�c�f��b
?]4?U�����̾�׽�Ν�������[?Ѫ<?�6 �����^�q�T��4a�6V����t�A�Ҿ�8V�}~��Q��ԃ�Gބ�E�"��fE��W<?��?1��^ʾ�����Y� A&�/{$>*��>��>o�>��=�����'��e\���(�I�����e>i�Y?���>��;?j�@?�N?�?�V�>��>��s�|��>ӭ༧�m>��> �2?*	=?�?��>�@I?AP�=�ti�P����޾�["?&��>��?~h$?} ?L:��t!<ٜU�i�����"�<w�����=��J�c�D���e='83>�X? ��x�8�\����k>=�7?{�>���>C���,���
�<k�>9�
?@G�>�  ��}r��b��V�>}��?!����=��)>���=�����ӺGX�=���]�=�0��w;��c<���=!��=�"t��΀����:=��;�m�<u�>3�?���>�C�>�@��2� �j���e�=�Y>eS>�>�Eپ�}���$��l�g��]y>�w�?�z�?`�f=��=��=}���U�����E���\��<ߣ?-J#?&XT?\��?c�=?Rj#?��>+�_M���^�������?�,?�ݑ>+��ϔʾMè��c3�r�?/�?�
a�f���T)�-�¾`�Խ�>?6/�� ~��쯿RD�T3��p��'����?Ƹ�?pe=�%�6�!����'z��d�C?��>Q[�>i�>|�)��g���&d:>���>\R?LN�>��8?=�R?�qA?x��=f�)�����w �e������>+�n?SoI?�h�?R�?=�>"�>S�}�ڛ־���8^̼-�Ƚ�k潰�=�>�&�>@�?Q�>DD�<�����-�����t>�n>�N�>m�=&f�>�Z�=���ǅG?:�>7��5p�����b�i�d��r?��?l$?1"� H!�Q�K����~�>)�?Gf�?��?�Fv�g��=CҼ����*t�#d�>�@�>���>T�>5J�=� �=��>5��>Vn ��m�J0.��*H��"?�B?��=��ſ�q�aq�ۡ����i<JR����d�_7���V[���=,���&�����[6\��ڠ�����+��ڗ����{�H��>�B�=�;�=�e�=��<�˼	�<�J=:͊<}�=�o�v�j<�c:�ֻb@��PD4�D�Y<�G=n�����ƾ='|?J?.*?*�E?�@{>e�>;o#�I��>�u�L?W_\>5�2��I��5,������N�ؾ�p׾`�����I�>F�.�
>��4>$i�=�8W;~��=獃=��=��7�}t =�=P��=Gɵ=���=��>rD>�6w?��������%4Q�#]��:?�:�>�y�={�ƾ�@?��>>3������c��-?#��?�T�?��?�xi�d�>����掽�m�=ᴜ��<2>���=�2�b��>��J>���J��a���'4�?w�@R�??JዿR�Ͽ `/>��7>8.>��R�(�1�b�\�U}b��bZ�K�!?F;��L̾�&�>gܺ=�1߾1�ƾp�.=,�6>��b=��dY\��ۙ=�z�v�;=.l=�؉>��C>Fa�=0�����=�rI=��=�O>���>�7�R�+���3=���=��b>�&>`s�>�?�P0?dYd?�E�>�b�TѾ�Tʾ�]�>��	>0��>�(o=��0>H��>V5?�jD?�H?k�>��X=�X�>�£>�|,�?�l�G�c��ՠZ=�7�?��?f�>�����b�Y�vx:�ֶٽ�?�	2?RH	?�=�>�����x�6��9���G�]t���r=�^�&�,��{�����i���_>���>/�>,�>F�>O��>E4�>F!�>�T�=z'�$m�=���<����P����=�g=�0��A�K���"=]�����D�`󽷼 ��[@�!��=�ʶ=��=��>�(>�_�>�n=����.>�ܝ���N���=����B�Yd�����/���9�F�A>oL>�ۜ�:V���?��T>x�>z��?�w?i1>����;�<��)�����O��=�S�=Z�9�z�.���[��Q�^�׾u�>�y�>�6���<������Wn�>�`�e�L�]t	��>���<ʈ�������������TS��(>�nW?Y��~�>���?��?�#�?��?~�D�8p�v��>���mu��������ݽ�Y���?�YP?p[>�|�k9-�%B̾����۷>�0I�)�O��=�0�'%�$ѷ����>��j�оr%3�Wg��������B�Or���>�O?F�?-0b��W��UO����6���r?wg?��>UJ?�??l;���w�zu��m\�=�n?Ĳ�?�;�?>�
>���=8.����>1�?>��?�?�k?�v%�?��m="8>�4L����=� >>3�7>�P?+y�>
1�>�a��}��#^�������ߦ<��o=��{>@�s>��>��>�ek=���=֮u>�P�>~�L>_�q>\X�>NC�>1�j�y�ξ9��>�!s<��>�8?+Х>8x�>a�L���Q<&m=�>�E���0�Wa3��O����<=wZ>��>W��>���ͮ?��>�K+�x>	?F3����@s���ނ>N�/��r?��Z>�i�>���>̱�>�l>���={�A>1��z�=�w�b����#��쁿�B���^r>ūϾ�<X�MU�}w����āؾ7��}�(씿0�>�ic�=Fx�?���;�����@��
��n�?7Ȳ>��P?�@��]�����N?d2�>�K��q����~���
�U�?�9@�d>�h�>��W?�?��2�3�XaZ�&�u�}OA��d�G�_��荿)�����
��H���y_?�x?v�@?f�{<3�y>v��?��%�۽��PJ�>�^.�+):�8=�Ϧ>0�� Sc�Ծ�-þ��E>>�o?'�?ٵ?aX�Wݧ=��>�:V?�?'y�?S?��>����{?���>6F ?��?�3*?x��>2�3?#:�>L�����	��&����Q���R�1����Q=ӽ~�������%����z4
>�F�=�<Y���IX���E����WpW=O9�=V�a>���>Q5]?��>��>��7?2��x 8��]����/?ʣC=A��Ј��6顾"��.>�k?C��?��Y?n'c>�A�~C�l�>��>\�%>�V[>o�>VF�ΈE��͈=}�>��>���=��I�lʁ��	��������<%�>w��>�\�>s[��k@>�i��炾Р`>�!)�鷫���]���L�ߊ4��y��&�>�jN?��?Z��=������Ͻ�c�:�&?�C?�'P?rM�?�B�=|�߾S;�<��Q �7�>#��<����0̟������W3�H1�xȃ>m��� >2�oJ�>���+���`9��y*�"��@�8�#&	�g�z� �$�&�����վ�2=�S�=������ �䤞�u����P-?��	=�ل��d�þl�=i?�P�>L=��<6=V�l���>�?E��>�~�����
IB�:A����>S0?�Q?���?<���^�i�"\�u����Ⱦt&d��?:?k�v>�Ʋ>L\>���Tu����\Y\�Fm���>SX?~�,��b�����'޾,�I���)�0�>6X>yF?��=?��>��>,��>��?�;>��
�ݨ�H&?�փ?��=� ̽(�N�x�6��J�.��>t�%?p�N��t�>��?�?��!?�~M?`?�{>!��P{B���>7V�>W�<v���4f>s�J?꾶>{W?o��?O�7>|�8�x���.[��!<�=�� >�*2?�A ?$|?��>���>,���>�d=wT?7'w?�0H?z3>D&?Q�!?@��>����?�-?g�C?��?��T?��>?5#�>e؃=��O���ǽ���ѧ�<��˽����s᫽����a�:��;�Ե=qL>~�;�{<J�����a�¼^q�;5�>�ft>㳕���1>u�ľ�6����@>]\���;���(���{9��d�=�
�>w}?f
�>9�#�8͒=΃�>qy�>���9�'?�?�9?�S�:�b���ھoxK��}�>�B?���=V_l��q���Tu�1�i=Gn?@$^?��W�w-��Jvb?+�]?Xo�[*:��gľtd�؄�iL?!S	?��H��{�>�?̅o?w#�>�vj�:�n������`��:k�p��=���>�����d��ۜ>��6?qI�>�k`>�s�=�fپd�v�ę����??�?�,�?0�?�.>
So�7�࿈��������Ed?�q�>5�jfN?�ڼؾZ@��o�F���e���㵾x����ʾ^�<��'������R>P�?rO?��?�.�?@���W�s��֊�>b�$s�����K��6���(�r=���	�G����gʽ|t:�V84����?�uN?1ǆ���>�����꾄���-��=��|�A����8�</=���;����,��UX��	��x�?f�>>X�P?�[��'Q�\"�z�+��2����
>�%�>u>Q��>���<�Xg��k�=�U�����=�N�>B�`?�;5?�{b?4P�B��������W�������� >x�)>���=	垽drf���$��kI���c��/��Ѓ�O����0��� ?���=h��>H��?T+?
P������g��Y/�@>�>��?�1�>���>��e�M1���>?�l?w��> /�>1���KS!��{���ʽ���>���>l��>3p>/�,��\��f��߃���$9�*��=I�h?�x����`�Vͅ>��Q?�g:DG<�z�>��v� �!�!���'���>�a?���=�<>�ž��0�{��k����?��>���{���>�4?�(?ظ>ڈ?�`�>UG �`V��[iE?;�p?��f?�{Y?7��>�؍�L2��_��@q8�U���[>܌�=�W�= #>{ӽ�`�u�3�Ve<�"�[p�=҇��b&�Z�=��=�c�<Z��=pQڿ?J��}־.��ּ�!�Ί��P��@���v6
�HǮ�7���z�+��S�(���U�%T^�қ���h����?Z0�?�Ւ������H����}�����>o�b�n]���������:
���M߾���N�#���N�Ȼi��d�Ŕ'?/���6�ǿ����:;ܾ ?Q= ?ߤy?�K�"�ؓ8�� >@�<�۝� �뾔�����ο����j�^?���>�3x�����>ԏ�>�X>�Jq>������<�?�-?Ѯ�>y�r���ɿ������<*��?��@�xA?��(���9�V=��>�	?��?>hM1�fS����n�>�3�?��?K�M=��W�^K��e?�<S�F�z޻Ѿ�=�f�=/=r��}�J>#V�>0��A���۽@�4> ʅ>."�:���S^��`�<��]>5�ս�3Մ?{\�wf���/��T���T>��T?�*�>K:�=��,?k7H�\}Ͽ�\��*a?�0�?��?�(?eۿ��ؚ>��ܾ��M?[D6?���>�d&��t���=i2�z|������&V�B��=u��>��>6�,�ً���O�TJ�����=�� ��3��.��D�:�+5ƽ�
����'�R:$�_S2�Wу=n%��b����-ᅽ���=Eb�>B�>}�>�R�>�9R?�ą?b��>^j�=������4�{Y <���w����v�p�ڼR���т���v��3��Ǿ��6ѾqF��=��h�=��Q��v���Q ��Kc��^F���.?{`#>��ʾB/M�Ǟ<ɜʾ�;��de���t���	̾5_1�xn�A��?��A?�ᅿݜV����(������pW?���U��¯����=�v���=h��>d��=�b⾓I3��1S�U/?{?�K��>x����.>�d�<8+=@�-?em ?<���>1�#?N�+�4V��U>�/>��>�M�>�>ŭ����>=?	T?		��"���ˍ>�S��wHj�	�=�$>_'������`>$��<.���������<Q%W?��>��)����V��.���==ȱx?]�?F$�>�vk?H�B?9L�<�v���S�#�Diw=��W?�-i?#�>�u����Ͼ����I�5?�e?�N>�Wh����n�.�UX��?��n?�W?�p��t}�M�����Wo6?�v?6^��Ƞ��]�<�X�(I�>߄�>c��>�:���>_�>?Y� �h0��,s����4�N1�?�@3��?�
\<����Ս=&?��>0�O�Դž����Ҙ�� r=i��>�a����u�(��'3*�Q8?���?g��>H���Bd��F>�������?���?���d\�=W�3�C�v��������y�=� >�0b�,����Z���־��8����w���N> @��$�Z�?'p�����#)׿<˅��"ƾȨ����$?�>�E���|���e�9长p�K���-��[�T`�>�?>���������{��^;��������>�|����>kT��;������6<��>���>r��>!����6��%��?�Z��(οo���0��T�X?(f�?z�?8�?H9<�w�	�{��X�#:G?��s?�Y?�#%��]]� �7��Ow?�Lq�M#��`�(��2i��kr>��\?�3)?s�\�o��=��>�0?r�>>[�!�Ҕ��祬��RX��=�?���?YR�P6	?R��?�T?����q��J���L���>8N?LIT>Og��˲ԾElA��"��E/?���>?���&
�U�_?ٚa�!�p���-���ƽdۡ>��0�;f\�4N������Xe����@y����?8^�?M�?�� #��5%?��>a����8Ǿ#�<���>y(�>*N>�A_�ڳu>����:��h	>���?�~�?�j?䕏������U>��}?��>���?���=�w�>�=�=Y���,g��#!>��=rC���?�M?�>W�=��8�5S/�B�D�[�Q��E�y*C�3��>M�a?,EM?K`>`����|6�Y ��ǽ��1��F���iB�pl=��۽��4>t?>��>vG���Ѿ\�5?�c򾝍��횿.P;�"/?��}>Z.?��@�+�����=5W?�0	>�V*���������S>QY�?'�?�t?,@վ�H"�vՃ=D�]>�;�>r��=�=�VᾈA�>��X?�g�=	��x�����>��?�	@��?�W��q?PL �n������ȸ�)���C�=n�=?���ia>���>
��=*>v�1��,pw���>_�?�:�?�(�>j?W�l���B���=�]�>m�o?��?␜<|����Db>��?z���̍��W�V�c?R8	@��@�4b?ؑ��	�ۿ�S���ܿ�M������=라� �=����k=}����'���4�=��>KB�>�v>���=8��=��{>!���H�!�$E���{���_A��$%���P)�����䂾�`���1���B�����<�l�f�v�G���"���g���<>��b?�U?2=�?��?^+=�H�>�����>/��l���\���8?	�-?��D?� E>��+��s�C;b�ܰ��\�K�Kn?�]U>gi?^C?I�>/>�=�>��>��>^��>F=�=o�������Z|>�t�>�/?�?�C<>�>/ϴ��1��M�h�w�R̽�?q���C�J��1���9��⦷�^i�=Hb.?|>���?пk����2H?���])�\�+���>V�0?�cW?�>���H�T��9>]���j�|`>�* �jl���)�{%Q>ul?[͆>�>!�"�:�0�S�B��{��j~>9?�+��w]:����	%M�#�۾X�>�W�>��л����������٫t���=�@5?;q?�nS���þ�,H��C����>��>���<��'=�ƙ>�j�<���=��.�[!=��=���>��?�0>~�=�+�>+���KN/�im�>�;3>k�>9?��#?�f���9����n���-��M[>[��>�s>�9�=�H����=�>�>�>a_��ܒ�\���R/�Y�h>qR��*)f�����0*�<[r�����=�­=VM	�cRO�5m+=�~?���$䈿��	e���lD?V+?s �=
�F<��"�E ���H��G�?q�@m�?��	�ܢV�;�?�@�?��1��=}�>׫>�ξ�L��?��Ž6Ǣ�Ɣ	�))#�eS�?��?��/�Xʋ�0l��6>�^%?��Ӿ-��>���M��x:���4s�m����Ř>�A?� �av��I׆�о>�#?��[p���	п����j��>���?�X�?�9H�����z?��`3>pq�?��L?U0�>���&@�l�>#�V?�V?�'X>�� �U���C!?��?�?�1�>q�?y�R?��?������Vtҿy���1Z�A�s�}�>���>�U��u;�ox����~�ǹ���9y�:_�=���>+t��O���ߝ>��<��S����z�>�>��u�7n@>�c�>���>���>*�C=Y0{��������M�G?[(�?��{�U�a�=���<��?�!�?i6?��f�U_�1�O>�XM?b�?\f?���>}b�1��E�������<�C�>�}?F� ?ٱ����J>.\o�*�=��C>$�>3Fn��
��|�q�}�=mկ>�j? ��>��$>�� ?�#?*!k>��>�lE��,���8F����>I@�>>�?��~?�#?� ��zR3�$��`�����[�<�N>��x?6?t�>����=k��F'3�}�J��쓽j�?_Sg?}����?��?�u??�A?/�f> n�!�׾i/��nπ>f�!?��k<��R&�l��;�	?p?2�>�S���Ľ�B.�9���c7?��]?|'?�1���]��)��d�<V<໢f����;ш�nL>�p/>�]�3��=�>�Ã=,�w���3�10�<�>�=���>��=�C��+����0?J�0=�ܵ���=�_}�I�J��>���>i�辠&M?���яR�el��$i��@Ֆ���}?��?�&�?v���U�s��F?7��?�5�>�?2���ؗ��G���H���h�ݨ�=S�>jX8�O\ԾM:���W���;�����������X?M�>�V�>��?�>��>y���V�!�z���V��^S���g�c��`1��"��������"�>�,��$?���о>��A�.��>r�>��>���>��?L��=f�>�9n>0@>oٻ>�g�>�)�>��>\u�;BV��{KR?y�����'�׷����=3B?�pd?�0�>��h�Ј��u��D?c��?Rs�?Dv>4|h�>,+��m?�>�>��q
?�W:=�3�\�<#S�����;+��������>�Q׽� :��M�$nf�dj
? .?�0���̾�F׽j�1�e=ʌ�?f (?'�U���o���V���R�	�*��Z�M��)�%���m��M���׃������'�ث�<;�*?���?������թ�M�g��?��-^>�H�>m��>w �>I>�����3���`�u[*��H��Ì�>�gz?w��>�m=?5%J?5�K?�8<?���><n�>-�_�e�?� �=�]>Ke�>aQ?�#?Z�2?�?��?���<���{�վ�=Ծ�u??�y?7]�>/��>K챼�����P4�f�*�����ɽ7�:f�&�(=�����������;�>=V?�{���8� ���E'k>+~7?���>M��>
V��|�<���>f�
?6K�>R���ucr��_��P�>z��?���ҕ=&�)>���=����:Ⱥj��={���Pn�=�̃�@)<��<�+�=;��=��j���e\�:X�;w�<�t�>B�?}��>�C�>c@��7� �;��ig�=�Y>�S>�>�Eپ�}���$��o�g��]y>�w�?�z�?�f=��=ە�=�|��[U�����&������<ܣ?^J#?BXT?^��?��=?/j#?�>�*�>M���^�������? ,?+��>���>�ʾ�-�3���?�]?R<a�����:)�!�¾i�Խ�>f\/�0~�����D�-t��8��_���}��?@��?1�@���6�ez�߼���L����C?w�>(R�>l�>��)�<�g�6 ��,;>��>IR?᭼>f�H?�q?H�[?��>e������I������WJ>hC?���?x�?2[~?,-�>�{�=����ھ8D�Kb�/���n��Rs=�/>���>���>�_�>�L�=6�<�!�����W�>��>���>��>���>��1>��o<��G?��>F9�����/���ɐ���<���u?p��?��+?<�=���m�E�`+���_�>Uo�?���?�-*?W�S�B��=�4׼�඾��q���>�͹>�>?Ɠ=� F=t�>/1�>���>��� ]��g8���L���?!F?�ݻ=wV��)aM�hn��Iƾ�Zz>����S��3��cѷ�3�C�
��
����j�E;'�_�6���޷�1⑾s_�J�?3A=�=��=���=�!��8:=�@ջL�����ɼ��=Zt�d�^���=��.�ǒ?�1�u=>��<A��B�ƾ�{?��H?�,?�>??�>��>��K�>@�>t=��Z�?o]>�c;��p���d=�
ǫ�>��g�־"�ؾ�e�-��� �>W|2�=>$7>tW�=�h�<l��=^�=5W=Z���=.�<s��=n��=�A�=l��=��>۵>�6w?W�������4Q��Z罥�:?�8�>[{�=��ƾp@?y�>>�2������yb��-?���?�T�?<�?Eti��d�>M���㎽�q�=O����=2>}��=s�2�T��>��J>���K��=����4�?��@��??�ዿТϿ4a/>VQ4>C� >��Q�N1���V��Ll�g�Y�� ?�k;��5̾=t�>���=t���ľ�z'=4�1>��U=]��'"\���=�tv��`2=�Bn=hw�>�?>�'�=����t)�='�C=��=�N>�|�?F��K�?�=
��=�^>o>$>�?�>b�?��0?�.d?�t�>Om��@ξh���K��>`��=��>��=N�E>)�>�8?8�D?�tK?S��>�9�=��>�I�>�7,�g�l��_����O�<���?[Q�?���>��<$�E�L��v�>�V,Ľ�u?.�0?��?���>y	���Կ����F��6N��p���ܼ��c�p�;S�m=�B�чX���>��>�P�>0�>>�c>KC >a.>�~�>rwP�����^=�݋<�]�<�.�=�)�=�t�$�>���=_��<�M���*���$���<Vr�=w��N흽�>�X�>�A3=�W�>�#"=I@���L�>�NW���X���<]Å��%#�*X������;���y���A>�r�>�N;<�>����?:��>	�=�,�?-gr?�&�=y�齨�\Ԣ�����C����J=-C������A��u�KJU�xמ����>�=�>��&>��=*Z�w�/�Ҟ=>h���U�A���g>yH�������
��,��(O���/���_��ί=��[?Q���K�=���?D�#?�
�?f�>�$��R��M��>�瀾'D?�@�)�(߃� ���/?Ϧ??P�>��⾍�� ̾%S����>cI�s�O�X�����0�y���ӷ�O�>[ת��о�3�Kv��N�����B��Sr�w�>O�O?P�?�zb��H��0@O����㊅��_?ng?��>�c?JQ?K���՜�A���'�=��n?���?e5�?��
>��= �<X�?G�?���?mg�?�o?�-轢?
?���=Y	>bΎ;��;>���=� ">�"8>��
?���>'��>c���J�� ��^4�Gyn�yJd=]P�;�p>>��U>0t�>X�u>ϩh>��>R�>�>�g�>��\>0��>�&B>�Uh�{�{��>�ȥ�<C>�@*?�m�>��h>&<�D��=غ�=mo>ͅ������;�VK���-�<%�@>fYW>�y�>�\�$��?�>&6I��%Y?�������O&>6�>�H�c�?u��=ZC�>�Ob>c��>�l�=:]>��}�,�����=�:�Z>�����g��x	Ѿ�}K>�Q����K5��X��˛������g�(��텿Sl��|?�7t;O��?/��<����l+�.����?HMs>�'?�$D��}l������>R߹>�A%�R��%✿N���Iy?l��?_Cc>��>��W?��?�1�H3�.xZ�c�u�s%A�Te���`��ݍ�����>�
����]�_?�x?�jA?��<9;z>���?��%��ɏ�� �>�"/�G$;���;=S�>�%��M�`�2�Ӿ��þkC��)F>��o?n�?&O?skV�,��<a�j>DO?iL!?6�?H�9?�-:?;d�<H?&�?��>�S�>��T?�v'?)?NZ�>)��=�W��o���zޅ�"Վ��-���V�"X��T����~��R�v�ws���@>�K�=����W�8��
8>8x,����=�Q=ʞc>)�<+��>!�]?g"�>�l�>_ 8?�$� �7�F�����/?�H@=R����������b����>��j?��?>cY?K�c>�A��-C��*>+܈>݇%>ֻ\>8m�>�2�6�E���=�+>�<>���=��J��ρ��r	�l'����<��>���>�S|>�����'>Xb��Q-z��d>R�Q�����E
T�Y�G���1��_v�b_�>��K?t�?�f�=G|�"���@f� ))?�[<?�QM?��?g%�=C�۾��9�شJ��K��>Y��<�����������:�^��:6�s>C��u���o�5>���"ھ��\��q]���
�6��<y���b�<T��׾�C�����=�&�=GҾ�,��`�� ���v�K?�P>��|��4x���Ǿ�&><ژ>Y͆>�r��5J���;�@���;�\=*��>�%�=z��2�޾�wD�4��Ӕ�>{�2?��@?�@�?c�v��s��ĵ\�$� ��w��|X=�/n?NK�>�g�>g��>3��<�]�����/v��\�<�>�:�>��F��]-��#���ƾ	sҾ�1>nݍ>ХJ��)(?Bwr?�s�>��?�"?*�>� �>���;�k���'?&�z?H�j�&��=D�4��+8�2/%��ь>;��>�����>T�S??��>��?��H?|�>P�;=�i��om��>�k>z&C�$A���E>37?u�?��A?Qb�? R�<�o����)h�������>+�?X�?���>-�>Q�?ե������<��=3_?l_�?�Pg?{�>�c??���>^�S=���<Km�>+��>��7?x�j?��S?R�2?cf? �ż_>����9����.����"�
�=x���L<�i�=��'<�ć=(e���ѽ]1�qvܽW�;W/M��|�>u�s>E���0>��ľe"���uA>;���	��nÊ�;���=��>3�?�ו>��"�8��=ߙ�>�>���*(?�?��?v,;��b��۾IUK�H�>xB?*V�=�l��g����u�Xi=��m?�h^?�W�?�����b?�]?�Z�U�<� �þ�c�ߒ�c�O?΢
?��H�\�>2#?�q?
��>�e��#n�+��kLb�u�k���=Eg�>�T��e��#�>ۓ7?���>�b>f|�=��۾��w�s'����?nҌ?��?�?�!*>�n��#��$�!8��{h?���>9о/�!?k���ڭ����������۾���S$��H�������T��i����É�U>��?�Hh?��h?�xk?Z��U�S��Z����;sY�����.#�B�P�2*1��+���z�a���O	��O������l2�
/���?S�=?ț{��?|�q)���>��(p>�\�f�����-=:�5=��=i��=��������BBL�KQ?��y>^�>�X\?(�1�~�r�jw0���\�W^"�I�>�p>���=t?�6>�Ci����!� �ؿ�-����z>f�P?u�:??l�?�q����4�9�o�w<�� R�d¾(h�>�<q> p�>�k齱%�x��~-��|�S!+��cp����[sc>�p&?���=.�>�Ę?�9>?3^}�|zj��ž�R5��?����u>�wg?
J�>���>*�8������>�l?���>��>�c��m:!�m�{��н(�>���>��>�so>�,���[�􃏿Sa���W9����=�Th?������^�p��>��Q?S�&;&�<<�1�>2�{�c"����#%��U	>��?�f�=��;>`
žo����{���5-?� ?��۾zpE�=�>6,?���>?�!>��r?"��>����S�o=aCT?�N?iot?{j?���>k@�>�Î>��9������=s>�*^>g=!��=z����ǘ��->���=��$=Ϙ�=�|�=��o=��>0�>�v�=��@>�ԿG�V���߾`���;�3��:���5�����I?e�Ҳ��尾g��JO�G5"��ms�X��9ن���_���?�?�?�ƽ�S��撿-�w�_�)�|��>0�s�HK¼�����*�?���l��w¾~L"���W�K{�(��Cj'?ΐ�:�ǿF����ܾ�m?7�?�y?>���"���8��� >���<�٧���eԚ���ο�>��:_?�X�>��߷����>�|�>?_Y>�}q>�����~���n�<�?ؤ-?��>��q��pɿ�����ɬ<�?7�@|A?�f(������X=!b�>2	?�@>�1�H#�d8��8��>�S�?­�?�
L=LW�b�
�1"e?Ŭ�;17G���ۻ���=~Ӥ==�U��dJ>�>eK���?�1e۽��1>s�>�M!�h��-�]����<ch]>��ֽ���Ԅ?x\�f�/�/�2Q��$k>��T?S'�>�E�=2�,?�7H��zϿ�\��&a?�.�?5��?w�(?�ֿ��Ԛ>��ܾ3�M?A6?�>Xh&��t��p�=�>�ڤ�W��$V����=ݴ�>ly>��,�'��/�O��ߘ����=9���M/ҿ�-������]>�7�\�4˽ �⽯Ie�s�(���½�X��^>y=@�>=�l>D�>�S>��S?��D?��Z>#�>US���fԾ��ξh2`<#����Us��s��z'.��|���iľ�յ���N��R`�Z�t�4=�Y��=5�Q�q`��nV ��Uc�kG�]f.?��">�˾��M�dc<�[˾�����扼x6��<�̾��1��Dn�9��?(1B?�z��k�V���|���ӹ��V?{4�E#��F�����=����Q�=S��>��=���3��bS��[0?kM?p���`ј��A&>np�)>=��&?�?���<��>��#?5�7&ӽ+5m>k�A>9U�>��>q�>"P��S)Խ�]?VN?�"�Q5��F)�>���&j����=�>/90�G��#1i>�� =�����m�~���,=(W?���>��)����i��e��-h==��x?��?�K�>@_k?a�B?_��<�`����S����nx=��W?e&i?��>_����о>t���5?,�e?R}N>�jh������.��:��?�n?�f?\��J^}�^������v6?]9y?raW��ҧ�����+h���>1^�>��?�V�)�>H�*?�巽������ҺG���?,�@	��?8Ɏ=�����ww<�C�>YM?�O��¾�yp�`���g�=��>�hG���|������0�2?a�h?|^�>�b������>`ǜ����?�|�?�i��/=��Ir�����wkO=1�<���e���ľ7KQ��ϸ��&�������<i�9>�4@�����+?�i4���п�̥��ޮ�4�(�y�v�A;?�>0X>A�����x�o�ӐB��Xm��v��U�>j >x���K���(�{�ST;��h��^�>X9���>ΩS����Oz����/<J�>���>Xφ>}���3Ͻ�ᴙ?#d��\&ο�������X?�E�?le�?)q?><��v�9E{�.w�)G?��s?�Z?�$���\��,5�	1p?�s��~���>�'D�~H>mC$?���>>�P���=E�D>hP�>�!������ȿ�^���tP�iQ�?s?�?qj���?��?j[?��\�� �g����W�=��W?>ͧ>�j�B�ھ�N:�e�b�*-�>s�?Qm��U����_?ώa���p�Z�-�T�ƽ�ܡ>r�0��\\��x���L��Te�k����y���?�Z�?��?����"�$:%?Pۯ>%���8Ǿ�7�<�j�>C �>�N>8g_���u>�����:�v	>��?�z�?�q?����1����I>v�}?���>e�?���=���>�}�=�B���t��H)">ko�=rTU�:�?W!N?�^�>	/�=W�6�f�.���E�N�R�����fC���>%�a?�	L?q�d>�>���!�+���ȽG)-�h+�E-E��3*�o|��L7>8�=>_f>5�E�Ifо]D ?����dؿ����P����?\@_>:�?<��&dC�r���pd?��=xR��}��|O���	�4x�?5��?dQ?�U��2ڽuV=�r�>�X�>�Wý�'� �Ҿ@��> m=?�l��&-���dT���r>���?V�
@>�?�k�7?��Ѿ�=���v��6,��*����=(/X?�����>�l�>c�F>�Ì��������k�O>�~�?��?dd
?zk?����;�Ѷ)=��>�v?���>ޟ=Z����5>�L?�H�̰�������hQ?=�@�*@�{a?����ݿ�Ț�{���3��iH�=�س=,����x���v=x
�=��H�`p罭�=���=�^>�Շ>C��=z�	=w�>~ԅ�.������]������G������)��w�������⾏���������	?�~�&�xE��8���t����b>�ia?��Z?�]?j�?P��=Gf?�����Ŷ>
���Q�%��ͻ4!"?@�?�&0?D�>����_q��ŀ��}�.�?�Q��>�6>��?�A?j��>"�7>Z��>���>�V=Zoλi >��'�V�����=9��>d��>1��>�C<>�>"ϴ��1��!�h�|w�>̽� �?[�����J��1���8��̦��	h�=Ab.?�{>���?пf���m2H?����+)���+���>w�0?�cW?�>���K�T��8>��C�j��_>�* �&l��)��$Q>�l?ah>�w>��2��6��LO���p=�>�5?�V��>�=���u��sH��ݾ4K>Ľ�>�1N�B����#�~���i�Ȁ�=��:?պ?"���C���I�p�G���U>�^]>q�=�c�=�M>�b��dƽ�1F��-=E��=��^>r=?�6>�Mq=n�>���)�C���>]L>U05>B@?~�?@f2�-��<n����!���x>э�>���>c�>�=C����=�+�>\lG>�w�5���`*�k65���_>�2���L���E����=s�G�i.	>��=d*���.���=�~?���'䈿��"e���lD?T+?G �=��F<��"�@ ���H��F�?n�@m�?��	�٢V�@�?�@�?&��S��=}�>׫>�ξ�L��?��Ž0Ǣ�є	�*)#�fS�?��?��/�Uʋ�-l��6>�^%? �Ӿ̾>9Y���C��Պ�2?��\�ͽ�q�>�L?�� �(v6��:��A�	? �>fL������ֿ�Mm��`�>���?���?�(\��ל���J�U�>iJ�?�M?��>*����sX�>��F?��?��>u��r$]�7E,?��?���?�P>���?4�h?���>�d��j"�#ަ�~����g+��N���Y�>h@>����.*������9u���x�v��k�=��:~�>������9I>Aj���ƾ�{ʽ/�f>��>��>���>��?T�>�~�>��=�S˼�(����⾧�K?{a�?Ϧ���k�7�<�ߕ=m�W��B?�w3?�J���<оω�>�m[?��?p�Z?f5�>�}�v��G̿��C��-s�<�M>[�>"�>O߁���Q>"Ѿ/?��!�>^s�>8����ؾ������}��>�| ?Ɍ�>Dۼ=�� ?ѝ#?p�j>�#�>�`E��9����E����>���>nG?��~?��?׹�=]3�����桿��[��AN>��x?oU?�Ǖ>����������E��1I�v�ٛ�?asg?)E�q?42�?n�??n�A?�'f>��"ؾ������>f�"?t��A���%�����?E�?�:�>�k�E���+B#��%�=N�?��]?��&?W��'{Z��'��As�<����ջ溺��lѼf<>��>T��Ҫ�=�� >�I�=-�j���]6�<���=�G�>�=x�6��z)�� 0?�#=��۾}<k�o��P�~Ѓ>��>������?;�ی�uҭ��V���/˾� ?�?R�?%%t<��}��_?z��?
6)?"�>��ھ��+���\�< 16��+�1*�W�>Ҿ\Ao�p����~��nq��0a��o*Ľ��%?Bf�>��>��>��>��?��ֺ��q�����hx�j;��n�=������ij��r���"J��˾�B'���>�z �!�>�b?�ł>��O>mk?���<C�>�a>
3�>e_�>='>�_�>EZ>�*>��QHR?ߊ��k�'�Hn����� B?K}d?2��>�+h�2��������?mn�?�J�?��v>lKh��+��)?E��>��gf
?�:=~����<n*���E��ׅ��2���>�mؽ�D:�F�L��Kf�~
?k?��p\̾��Խ8?��-�c=�"�?�t?�3(��[��q��U���S��6�s������\�)��Ji�9h����L����(�|_<&�-?��?����z���-����ib�_Z-���h>���>"�>�>��B>m6�ZN4���g���!�u�\�V�>�,{?�l�>��F?U\??�N?�~I?���>���>�\����>F��;�+�>���>HQ;?�[/?^�0?�?�_!?��A>����N3��PIپ�	?I?�?���>ny�>G}���餼+���^g}�DѠ��e�=l�$=T̽����0='N>�\?���F#8������j>�7?@��>n��>`���t}��*�<,��>�n?�3�>e�����p��H����>�̂?	����=�>(>	�=�ۉ���W����=ϼ���=uV���2��G8<�X�=�=�A�:�h9z;��;���<�$�>�?J�>���>W)��� �W�ճ='EY>7�S>�>�`پdv���D��F�g�g�x>�y�?���?.7j="?�=~7�=�,�����J��������<k�?�a#?�RT?|��?�=?D:#?{P>����钿���������?r!,?튑>d��&�ʾ�񨿺�3��?b[?V<a�'���;)��¾��Խð>�[/�%/~����DD���������~����?ؿ�?�A���6�#x辷����[����C?!�>�W�>��>�)�*�g�Z%��0;>���>eR?u\�>.�K?<Ad?Hc?I�>�v8�,5�������A�tgd=�q^?l�?}ވ?��v?�/�>d>�ǆ��h���N��t��J
�:1o��=?�> ng>~��>�>.>�����^0�R��=��S>�N?܏>���>���=�J@�})H?"�>��������{��U5y���I�q?腏?l�+?l�<*��?�������>��?v�?�R*?�V�߲�=����sC�������[�>~��>PԈ>Ŕ=FiP=L�#>B4�>0A�>�r�x���n3��zG�vG?i�F?%��=ʷƿ��z�*����t���7�=���߃ҾK!�����!���젾9�6��[˾lF���4c��;���[�����?Xܾ=:r�=��@<�^��zm����=��%<�~��z<��I�p��.1Ľ���=󖝽+ܔ;��<<�<X��<�p˾ޔ}?SBI?g�+?��C?��y>��>��3�麖>!8���4?/V>��O�M����A;�f����'��k�ؾ��׾�d�9՟� 1>uqI���>�'3>c!�=G�<�/�=��s=��=O;�Q�=�=�=Ƅ�=J��=���=�>��>�6w?F���	����4Q��Z罘�:?�8�>X{�=U�ƾ�@?�>>�2������kb��-?v��?�T�?G�?�si��d�>,��䎽�p�=?����=2>���=k�2�;��>��J>t���J�������4�?��@��??�ዿ��Ͽb/>��8>,7
>��Q��g0��$[���d�DR���!?�9���;{х>��=��߾�ʾs�'= �1>ql=�L��a[���=)倽�<=��f=���>��D>���=z��>��=�a=���=�M>�|��j#��3���P=5r�=��_>�+>3	�>��?CW(?��X?q��>�L�ut���񻾸ʐ>��=�{�>��a=4lU>!K�>��7?\�B?�H?)��>��N=�S�>r�>��,�
r�a��������ⰼ`�?��?�A�>���;?b:�dY��J9�,����
?�,?u^?�F�>���W�:��;j7�ϴ-��4�<��X��۱�&��/�A?��*����&>�֔>��>��>�B�=P��=�<;�>cD=�^�=RE>2)�aL.��O�=��0>;��������<��*=��
��[ =VQR=�'��А�R^<>>�;?��=���>YU>���>�Y�=�����/>6����L�B��=M���:D�Ϝd��j����/���B��D>�]\>U�y�F����?Éa>r�;>_�?;�t?� >��
���Ͼ����a�i��hO�a��=���=�4��8��ba��M��xѾy�>0D�>�an>=�">[S$�mzC����=N:e��"1�F	�>��v�lb���x�M<���z��Ƹ��BM����=$B?�h��_�?>���?��"?�y�?N��>!�ɼZƵ���>��¾�3��8ݾg��8���w-?T,E?�΢>71Ⱦ�30��ʾ)�����>9�N�u�P��ʕ�	+0�櫚�������>`���k�ξS4��Q��d��:_D�ttr����>��P?Ү?�c��^��@�O����F{�WH?`�g?	Û>��?w�?2���B���|��e�=��m?��?S��?9>�Z6>��*�`��>?�E�?P�?��?�f#�|x�>(�=	����Î��#�={�=��=>��N>o\?";�>S7�>�Qy�0+�{����*X��Ȯ˻��#<t�d>CC�>)��>�=e�=���>l�>��>1k�>S.�>m�>�N'���ž��6?�t,>w3�=�F)?xcq>:d�>���=>�`>��8:0�]�Bք���ɽ�I�=�!I>2I�=�� >}��>�P׿x(�?s��>L�����7?5�� �k���<>��`>Hi��a ?�:���݆>��>W�?Na7<�&�=���>��ľuI\>wQ�im4�X�E�M}���`�>>�ټ�	T��h?���/�ϭ����?�-���o��pg�#�0��㈼��?2ˤ= �o�?�1�r����$?��>7SG?�*�A�p�4v;;���>�<q>��`ԯ����[����u�?L��?�<c>��>��W?��?�1��3��tZ�R�u��'A�6e��`�1፿k�����
������_?��x?uxA?�H�<�9z>��?_�%��ԏ�Z(�>?/�m';��H<=f,�>2)����`�ѮӾ-�þE7�TIF>Εo?�$�?�Y?,PV�q( ;YH�>W�@?J$"?4΁?��2?�"?����SJ?��>�5�>�$?�I\?��"?� ?"~�>]�<�ʶ�#?��N��H3���*�e��Ǒ�g޽ɹZ��Ї��m��������=�	'=�x=� �>�y�=��<��W�z=�0�=�Ҧ>�]?��>Ѯ�>��7?����7����H/?�#>=�U���b�����ش�ƴ>�j?�?�yZ?��e>�A���B��>�J�>�'&>�[>s�>'G�h�D�+��=�>wp>���=´J�6O����	�n.��cf�<�T>���>�3>���X*> ��jx���k>`�O�B�����U���H���2�u�v�)�>D*L?Y.?)��=����旽��e�F])?` =?/L?�c?yj�=%wپ�8��I�yq��>Fe<v������ԡ���9��g�:b�v>�S��x���2v;>* 
�!��l4j��sG�k�վ�D	=��Q|<8�1龹<�����=�!�=�_ɾ��#�����PZ��D�G?8QZ=¾���)D�h��>~��>��>�Q��T&��;i7������:��>��,>��������R��~���>rK??'�f?��?t햾�k��gF����至���ټT!?�>�?��j>cG0=�����S���b�MjN�lR�>��>�.���>�+叾�U�V�"��h�>�z ?3J�=&?�+M?�2?��W?�x5?�/�>�v>����Ⱦҭ%?��?M�=�p�D�I���3��B�!��>��,?'�+�8"�>~�?]!?�v'?�SQ?Y.?@>z��K>���>V��>�Y��̯��:a>k�F?�r�>�U?���?�A>�3������wQ�=$8(>�E5?�|?V?t8�>X��>�UH��@>p~>��b?̋r?�m?�&�>��?@�)=�5�>�S�=��? ��>��=?��k?���?VYg?m��>�X=�		��B����"z/��Ӯ���B=xS9>MP:��ǹ�~ڏ=�S=���=�R>VӚ�'���y�9$��>��=�V�>5t>=����2>5�þ񇈾m�A>V����_��/���	�9�{��=[��>��?0;�>�� �h�=t8�>z�>��� �'?U�?d�?�]�: b�:�ھWwN�Fï>/�A?p��=3tl�����W�u��h=��m?�^?�V����(�b?R�]?5&�W=�ߗþwb�HF龌�O?��
?�F���>�?�r?��>�me��n�Q�Mb�'�j��i�=!&�>
d�;e��!�><o7?���>g(c>M�=N(۾�w�(R���	?��?p��?��?��)>}�n�!�a�{��6^?���>bA��_w"?���#Ҿ*M��Ŕ��r�߾`��ד���w���X����a��S��rt�=��?-�q?v_j?��b?n���i�t�_�<��~Y��| �z �PD�u
A�D�E��t�88����I(���r^=�x5���^�n	�?Pl?^�_��^?�8��U�徧���gU�>��r��G(��� >C�=�/�=�AS��چ�C"߾�]"?3u>�k|>�6U?O�e��J]���<��"F���)���<'E?Hǐ>d��>�7B��
���ս�Ӿ��un����>Vd?��1?ۖ{?��g��1�Ez��'`��)��>���1>�i�=O/	=[���_Z� 2�r&&��B����)�N��yr�D^㽶�?t��>��>�?� ?;��μ����	S;���?���]>�.d?�Y�>>E�>%\ �K�žwf�>��m?a�>�>U]��NP"�>�~��ݽ���>���> ?�=u>��.���[�y���w��i�8����=4Wf?p����`�nC�>�!Q?�L;Q�g<ԥ>����D!�O��J,��#>�]?I�=�N:>��ľn�	�W�z�����l!??r�!���8���?v�?�5>�ss>��?�:�>
J�7O>�a?�/k?D�c?E�v?��.?�G�>��<Q��v�k��̽��!>	��>�a=i[�C�=�b������6������=%��E���3=� �=��?�|i�<x�>��b������9�����3��Ɔ=�ܰ�R�e�aq��}�Ǿזr�tqŽC�ؽ�D���`��y<�Dl��L��?.�?�O���WY��ā�p�hξ)ʂ>&��N����L��vþH���*�s&�N^��Hr� �g��'?����A�ǿ�����<ܾr ?>> ?��y?1���"�ݍ8�d� >&��<J,�����n�����οe�����^?l��>���|������>���> �X>�5q>���Gڞ�N�<��?ډ-?��>�hr��ɿ%����s�<���?��@6{A?�(�W��C�U=���>��	?
�?>�L1�@;��갾�Q�>�<�?��?�M=6�W�$�	�!�e?Q�<��F��$ݻk��=��=s�=4��x�J>B�>����1A�N�۽�4>j�>�"�����v^�8Ѿ<�w]>��սX@��5Մ?*{\��f���/��T��U>��T?�*�>[:�=��,?Z7H�a}Ͽ�\��*a?�0�?���?%�(?7ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=a6�Ӊ��{���&V�u��=Z��>a�>��,������O��I��M��=���dѿ�m.�@I5�_�/����k��$w������hM��z P�Ho���>��="�>�f>v�v>*>�f?kv?"��>;�O=�a=��|��TM���f=b!����3���n�H�L��z��s����x�|��ξ��p&˾�j>�U��= �R��ؐ�
� ��c�� E�ic.?��>�T̾�=L�ИW;��ʾ�u��6]��,�����ξ� 1�Z�n����?�`A?� ��e�T��Z��y�!ż�zIT?y��U�b���ր�=3���=t�>SY�=�i��'5�źS�50?�q?�˯���w���N>����@JK=��-?�8�>���;���>W?|
,� p�"ԅ>�^>���>E�>��=���ر���#?��Z?d�콂�����>�g����A���=t2>�V����<K�W>P8=EO����<J���x.�"W?���>��)�%�.Q��
��(�==��x?��?u6�>#pk?��B? ��<>X����S�g��yx=#�W?�#i?մ> {���оЇ���5?j�e?��N> �h������.�X�#?��n?�X?^���o}�,��	���k6?�v?�@^�ه��B���C`���>��>���>��:�U�>n$??μ#�gՔ�����&q5�R�?�@Az�?�AP<�(�լ�=�U?%��>e�N�o�Ⱦ����&����n=Z��>�=���u�ٔ���+���7?$�?� ?�҃������>�Oʾ��?��?�?�������.���|���	>fK�=s<�=��ʼ������G�5埾�Y�@�Ӿ<�%�G�>�@c,��?𹛾L���vÿ5���T	��j��w@9?~�>���JZ��Cv��+��2�C��U���[���>��>A����y��@{���9������t�>
��/�>C�Y��ʶ�q��n�<��>��>���>�S�������
�?A[��9_Ϳkʞ�Ah��QY?�X�?�6�?q ?(2+<����^y������G?)�s?.�Y?ܘ#��U_��H-�ϭ]?黵�
�k��t1���e��~*>NQ9?i��>E=�2�J=�YZ>4��>���=�#�tǿ��������H�?��?�Y�B}�>%�?cU-?���V����E�k���#Ƽ�t^?�"�>ڼ�N��9�+������N?��D?��+��K"�\�_?*�a�L�p���-���ƽ�ۡ> �0�f\�N�����Xe����@y����?M^�?h�?ҵ�� #�f6%?�>d����8Ǿ��<���>�(�>*N>eH_���u>����:�
i	>���?�~�?Qj?���������U>
�}?KO�>��?���=���>�]�=�z����,�+�#>j�=#�?���?�M?���>��=�7���.��dF�:R�p�R�C���>��a?ÞL?ODb>!���h�/�o� ��;˽��0�Sp�6H?���'�-߽�b5>?�>>��>��C��%ӾV"	?�<�Z 远���fmݾA?"�<>��>���� ������6?�A>��Rl���d����!�߱?,�?i��>qP���=�j�=6y"=mw�>M01��0��ɚ�e׌>63?S�@�'ZY�@�A��/>���?t�@�p�?�Ё�d_?u �Ɍ��L}����|82��� >��8?J����A>��>ٌ�=�l������c~�� �>���?A��?��>�_?�|l��c&���=���>~�X?(�?j�=����[��>e?a��뉿T����^?x�@!�@b�U?l����߿쩩��I��u�Ѿ�ɣ=/��=��> ����E�=�{¼�����>�8>P�}>��o>H&�>��_>� !>V�>>!͆�`�!��J���ߐ�}>6�j0����zS�������q�|���⵾L���ͷ�������뾽�Rj���#�\���� >P�8?> ]?��?^��>�E�=%�>R�oT|=�7*�O�˽еE>�?��T?��1?�L�=�u����i��F�����A���YM�>;��=�,�>!0�>a;�>ۘ=�k�>�u > �=�B>�oE����=PN�=&zr>�c�>�>�Q�>��;>�d>�ʹ��2���h��Hw��˽���?�����J��'��qY��I����M�=P.?�D>F���6п����E3H?)�l�_{+��3>!�0?�SW?g:>,��&�T��M>���j��U>�3 �1�l�4�)���P>�X?��e>�it>~~3�3-8�i3P�Z����|>6?RW��0#:��Nu��H�.�ݾwL>�>��F�\��H▿S�~��i�9�z=��:?�?6����1���$u�������R>z]\>��!=���=3sM>�Ua��Ľ��E�u/=}c�=�]>؂?m/>���=n?�>������G��>�yG>��/>!�>?�w$?�A �5L�������$���{>�x�>�(>(e>��L��K�=O�>�b>���i~�b��B2@�y�]>��c��|W�{�R��{�=������=�=�O��7�>�=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿh׏>�W�Ҙ��'�w�%�p�&��T�>��E?��T@����A����>���>Ҽ�zR����Կ&�
?���?p��?�:2����`P�-�U>��?��%?��,>���}�U�dp>u�7?��v?L@�>��)� ����?�P�?.ׅ?���>z�?�f?/��>��a�u�T���п!�����<��+>���>�d>7��e�6�.牿�ׇ�.�o�~�/��F=4=�
�>����;˾���=o»&���Z�ڼ�;�>xٻ<a��=�Q�>H(�>��>�>��I�`�<	�U���	�K?F��?t��7.n� �<�ʜ=~�^��(?O4?eGY��Ͼ�>e�\?��?�[?n�>)��9��2俿�~���`�<8�K>�*�>G�>�*��61K>��Ծ�"D�m�>�Η>IP���>ھf#��N⟻ET�>�_!?���>&Ʈ=� ?#?��j>�,�>�\E��7���E���>Ȣ�>N?��~?��?�ѹ�RV3�k���䡿�[�)-N>��x?T?�ҕ>����8���tF��I�0,����?msg?_��?O3�?�??�A?�'f>����	ؾڷ���>��!?�	���A�5&���|�?OG?���>+���~�ս�ټ����m��?�*\?�9&?���+a�	þ���<��$��Y�M��;s�C�W�>�w>�^��Ҵ=m�>�=Zm��g6�ȋg<{��=���>��=S7��E��ˊ?v��hn���Е�D$��c�[����>U��>� �tb]?�!1=+�`������r��nҾ\�e?Ŷ�?�?���:0�i�~EL?ׅ?'S�>�0)?J�ھ1ľ�"뾁)��ܲ9��9�x0>@��>@ێ���� l��U꧿�ᒿH]�<k�2;���>�>���>@(?�Y>�1�>��ȽoZ�����B���g�<�]}d��A��R��-žQmž��=�qϾ����"{�>S&��D�
?�=?{lK>y��>Pz?���=���>}�>�(�>w?�y0?�~?,);�($>��KR?����X�'�'�输���k3B?qqd?N1�>Ni�h���F���?���??s�?�>v>~h�,+�"n?X=�>A��xp
?$K:=|�0<�<�U��m���/��u
���>�E׽Y :�QM��kf��j
?f0?-����̾*>׽�Zg��f=�[e?%1?�u$��Bp��v�y�q��>O���r=�B����ݾ`�@��fd�$̍�m��Vā���<�TźL�.?�C�?2e߾�뾪{����z��S�"IK>���>�>���>`�U>˶�X>���N��[C�����ݘ�>��a?�'�>��2?��,?mJ?�DS?��>M�>%��$�?�:B=���>:t�>	&?��?��A?��6?5N
?EWY>w!ѽA[�����:�?#�?���>���>��?8
��pT��ռ�����O��Ƚ��/��.ļIὮ>��=D��=�Y?����8�����Jk>i7?R��>@��>���R.�����<��>�
?<X�>+����rr��[��i�>���?j �c=V�)>���=�Յ�Q>Ժ�_�=����Ґ=����X;��<��=��=�At��(��v^�:��;�w�<��>�?�Ԍ>��>6Zx�����(	����=��b>�O>�b>eoپ͈���ٖ���c�%sw>��?�a�?� r=-o�=���=�i����þ�e�lھ��6�<
?`�$?
�W?��?d�@?z�(?��>���c=���ׄ��D����?x!,?��>f���ʾo�`�3�̝?�[?N<a�i��l;)�ʐ¾$�Խ��>F[/��.~����0D�b������D~��'��?뿝?WA���6�Wx農����Z��t�C?�"�>�Y�>6�>�)���g��$�X2;>T��>�R?%�>�@8?��?P~?�j<��(��ڰ��i��];>��ub=a?�+l?��w?cl?��>��S=(>��3b���,�����+�0�n��\>���>�?�>)��>�>��p>� ���J�����>>eF>��?�n�>�i�>�-A>^_=�G?R��>�߼��5��n���o����;�԰t?���?�X+?"
	=���LB�]���2�>>��?;0�?��*?/R����=�_��hc��wiq����>t-�>���>�a�=��_=�>ͅ�>�a�>����e�{8��PD��J?3?D?<�=:�ſ��x��þ�'վ��B;���(���]PG�n�X����v��:���B�W�D�;NX޾���fݾ����~�>:�	:�i*>���>#C�=��|�� ���Q��<�X��&
=�Ғ�}��%��o������X=�g��!�=�~˾֎}?w:I?Ř+?�C?�y>�D>�3����>����a>?V>gP�놼��r;�����E��ݱؾ�m׾C d�Kʟ�mD>yI�Y�>�.3>�?�=�D�<u�=��r=�=�ES�<=(�=OG�=%\�=���=��>`>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>��6>�>��R��1�'O\��c��Z��w!?#e;� w̾zI�>CV�=�i߾�ƾ��-=K�5>�U^=2���h\���=k{�9�==/�o=d��>P�C>;@�=]w��0�=\�I=.��=\rO>6��@8��+��%4=���=c%b>e�%>	��>�-?B2?�a?��>+�W�/�Ⱦ� ���(�>�Z�=C3�>�r�=�M>���>��8?�^C?gL?�V�>J�`=ȴ�>�i�>~�,���n��޾i���0�C<wY�?*�?�_�>����]1��S�i�7��ٷ��f?fj.?�$?���>�"��y��-�J�8�7ȴ�;���3�;$E�1�8�n�S�p[��S�;CY>w�>r �>J��>m&R>��2>1�>�3�>�>	�|��[H�NL̽v&�:yv�<N!�=F�����=�c�|�0�M;���=�Vc��˽��_�=Q���H@�=���>8O=���>�y��U�Q~>��d��gL��=�*���](��wU�z���:I�Cꏾ�%m>��K>���=���?\�Y>��>BH�?�V}?��<��[�}�g�������ݾ�-��֑%=�ӽaӱ��H9���� �j������>|a�>��~>�>��#��7>�0�=�;{w0�OE�>[,��R7����*�#w��-{��<G��c]�e0���N?�!��K{�=��l?S�B?���?�{?���/侫^�>Y��������$�C;���w����0?�(?Z�>����;�70̾�;���>r�I��P�������0��������!��>����h�о�3�]���	��k�B��<s��V�>i P?	�?H�a�PZ��PmO�y������\J?l<g?y5�>/1?�?�������5Z��!��=,�n?��?B6�?��
>�>�h
=\-�>μ�>�Ǐ?9�?�Gh?�]���?���=c�D>��=@ui>Ɲ>�v>~v�=B�?$�
?�8�>��)�'ھk꾳W�e����Y���缞`>��>7��>o�#>:l�>���>ٚ�>�؉>ّI>@��=��D>�">�Y��^�	�
�?�����>� 7?*O>2v.>���<I��>����O��`�Q�����l�^=PZ�/�P=�Q�=� �>V�׿�^�?ʈO>۲��	?����۫=z��=�>��L�z�?j�I>�h�>���>���>��=��>�<2����5�= �GE��a3�/��,}����T>�꾞�����̾�3���H꾖j����s"���a����D����=�a�?#lL;0Av�����@��?��>4�R?��M�,��)b�;'�?s��>S�پ�j����f��1��?�@�:c>u�>�W?��?z�1��3��tZ���u�2'A�+e�>�`�;፿g���Y�
�������_?}�x?�vA?��<�8z>q��?#�%��֏��)�>i/��$;��C<=�.�>%)����`�k�Ӿ�þ:1��KF>��o?�$�?�W?�PV��V�=;mq>߼1?�W*?d?F�A?�EU?]�N>�C?�:><<�>?�>R�7?#<?_�,?#��>LI>�Z-=p��=���\4���<�:o����$�=B�4>��=������ܽu�R�N6ѽ���<����)����b��x�=�]c=�KA>8��>O]?�S�>�B�>�D8?Z�o�6��ܬ���/?�b6=t����f��iZ�������>1�k?x�?`QZ?L�d>�qA�;�B�^e>��>ށ&>(}[>��>-V���A��֊=�|>��>��=��J�ׁ�y�	�[i��m��<)H>���>'/|>v����](>8���sy���d>�Q��l���gT��G��1��Bv��>��K?�?��=�I� ˕��8f���(?�9<?qM?��?K[�=��۾�:���J�����>1y�<�	����+��e�:� X ;��s>��������jt>�q�����K�f��E�+���N�<���sU<=�3�zн�叾ZG>���=������#�T�������uL?�_�=U^��;�c��(Ⱦ*g.>�#�>���>c��?}���;��踾�P�=�G�>��<>
�-�Q3�1O�Z���϶|>H>?�fp?��|?Փ��b�ȑc���2���c},�s�?P�>�M?�Z�>
\=�z׾d��HHf���L����>���>�Y��)2������G�=�-���<>�`?�^U>gr?��K?�)?�Q?i�?/�	?.p�>Lf�������&?,��?�q=5�½mS�|�7��9C�n	�>�r*?�?����>�Y?R?@3$?-Q?�i?��>�`���A�Th�>��>�X����b�U>W{G?�$�>��Y?
��?�C>F�4�hM��>W���d�='�>�2?"?�l?Ŕ�>�Y
?�_�j�>�\?�=?��p?bZ?(D0>(�?���>�c%?�d1���N>3U�=�?��K?HZ?��g?���>��Y���<ԁ�� M����;~7=��&>�
/>)h�zw�����{n��<�<�k>	'=<���b��=�p��a�
4�>{��>�a���->����ÿ�� .6>�
�<[L��������s�=K��>� �>&Go>��A��h�=�u�>���>?&�e�?��?FR?��鼈_X�+�4�W��+�>d�M?�>�Ug������h�r?>W�s?�Ud?K�e�����A�b?�]?Kh��=���þ��b����p�O?4�
?��G���>��~?r�q??��>`�e�2:n�$���Cb���j��ж=Ar�>JX�N�d�i?�>r�7?�N�>�b>�%�=>u۾��w��q��X?��?�?���?X+*>��n�O4�}Ҿj8����a?�/�>?)6���.?��a�?4��D��GRX�._پڅt��6þ�$=�g`�F~d�$JX�%/��Wk=*4�>柄?l�^?.`p?����I6I��a^������R��� �W[�e�S���F��u>��.�R&�������;�`�����@���?�$?� &���>e���q����	о��:>�ܟ��y���=}ug�|�>=��=�lc��H7��Ю�7?!��>eg�>c�7?�V���>�^}4�n;�\)���w0>q�>�7�>�}�>���<��6�¡�]�˾�����?�pcq>��_?�K?�k?,s��.���~��/��W��pD����^>J�">A�>=�G�U��We�/�6��v���rᇾ{~	���.<v�/?v�m>$F�>���?�9
?���F,���W���F+�&a�; �>�b?� ?��s>�w`�6��7��>�l?=��>��>^����Z!���{�Mʽ��>���>\��>�o>�r,�!\��m��6���S9����=ԩh?o�����`��܅>MR?�yx:4I<i�>��v�Ǫ!�߷�Q�'���>�p?���=;�;>rdžg�c�{��6����8?�u�>wľ�E��,���I��>�o?���>民?��h>7Lh�%x���%?��X?��n?�?l?(\�>[�D>+�i��l��׍>V�=r�0>n��=?��=��,���Q��G'�iߪ>5��Ei��D�=�;)>U�/��<��
>�ۿS5K�d,پϪ�'j�|r
��a��W����[��������:u��0gz����]�,��)U�y�c�D��%0l�b �?*��?0K������M�����~�����>wq�)Y�������5��S߾�d��Ǥ!��jP�ui��Ff�/n7?M�^�@�Կ%Ũ���"� �)?#�??qA{?�$$��U���E�] >�� �d��=��	�S䗿�ؿVY�`y�?!��>Z2���Ƚ�=?�~=�d
>���>u��<�2�����&G$?�d?��>���@*¿.i��;��ń�?�.
@�sA?��(�����PV=���>�	?I�?>�81�>��mT�>C6�?���?ZqM=ݭW�(�	�dve?[�<��F�/�ܻf/�=Ia�=#=���J�J>�U�>���aRA���ܽ[�4><ׅ>/#�L��
x^�q��<�x]>O�ս~��%Մ?#z\�Gf�u�/��T���S>��T?_+�>�C�=*�,?{6H�}Ͽ��\��*a?�0�?զ�?'�(?{ٿ��֚>�ܾP�M?D6?C��>7d&��t����=.6�#������[&V����=��>�>��,���q�O�gE��,��=\��k���.T��:+�Z
>YK�=�k��4J<���;�д��N۾��.�%���s�;>W�>y�>q]d<N=,>�>M?oT*?!��>��=?J�=�Oپ���[f�+G徸�=���Y^/> :4�v������:��%��T)�?ɳ��$��&�=0�?������̾&�T���?� ��>>�= i��y�
�>���q����A"�8=��uj��&C���p�)E�?J�r?�~���iV����	�%>_ؤ<��3?���	-�9q~���2�A��VH�=&rY>�o��� �pU�6!a�s�0?�?:����܋�Ь,>Vp��i%=PB+?	?�<~�>ˮ"?xu+�����)`>f�>>oL�>�^�>�A>o�� vѽgO?��S?'�𠙾.c�>캾�bz���y=}�>[C/��8��V>��;y����7�	����=^(W?9��>n�)���a��!�Xs==c�x?�?-�>�zk?��B?s�<�d��2�S���Grw=Y�W?Z'i?K�>򑁽о����W�5?~�e?��N>1\h�G����.�S�k%?l�n?�_?^`��t}����f���n6?��v?s^�ws�����K�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���yY4�%Þ?��@���?i�;<��V��=�;?l\�>��O��>ƾ�z������2�q=�"�>���~ev����R,�e�8?ܠ�?���>���������=Y���c�? ��?���}��=Y+��jz����a��o�U=�{_�X6��A��:)����i��X������tZ>�(@�W��8��>���9ؿ��ѿ ���6ƾ���gG?"A�>��P=�GQ��7l�'�q�n2:�gP�F���g�>2�>�Ֆ��l����{��_;��
��6;�>Ig��و>��R�ײ��p잾MD+<���>nx�>�F�>i���5����?�c���
οZz����u`X?�.�?�Q�?�x?W<av�e|����?G?��s?$%Z?��"��x\�G�8���j?aҥ�,6a�gb3�-�G�I>�y4?��>l70�9+o=;>�D�>&�	>�-�]ſ&@��X��\�?~g�? ����>59�?�p-?�������}���+��eƻ��??B5>
�N�p�=�(c���[	?��0?�� �4�]�_?�a�I�p�n�-��ƽ}ۡ>��0��e\�J����sXe���w@y����?E^�?f�?���� #�J6%?�>�����8Ǿ��<���>�(�>�)N>�G_���u>����:�ki	>���?�~�?Yj?問�����U> �}?7$�>��?8p�=.b�>�b�=��*-�j#>a"�=�>��?R�M?RL�>�T�=m�8�Q/��ZF��GR�5$��C���>E�a?˂L?�Kb>F��3 2�R!��sͽc1� O��W@�4�,��߽[(5>�=>�>��D��Ӿ�2?����?ؿ�斿�%�_3?O��>��?�W��z�عݻ�^?'�>��#`��`F��m��"3�?r��?�F?��ؾ��̼T>Ht�>0��>"j۽���wV��N�=>�HC?x��TH��+gn�m��>���?��@��?�jh�9	?���P���`~���s7����=Q�7?�/��z>��>�=Dmv�������s����>[B�?{�?o��>q�l? �o�8�B�z�1=�K�>��k?kr?[�o���'�B>"�?���(����J�M!f?��
@]u@9�^?����ڿ�+����߾K��ȣ�=��>>XP)>Iⷽ��>��>5�V�Ѳe����жN>�>>�}>2g>�y>��Q>����<�䄦�"֚�c�2�+����z,�X�$�ţƾ��4���ؾ�����n�X��DUۼᗀ�Ï�J%��<.�=W�L?`_K?^,p?�o�>IC��U2>���V�<�f�Wؚ=Ie�>j;?�;?U�'?�R�=�֘�@]�\x�Zf���_��S��>�]�>��>�&�>��>��{=�x>�G6>�D->~�R=��¼lΛ����;{�u>-~�>�
?}!�>q~T>�8�>��)�����d�6�K�G�ѽ�q�?r�����<�SQ���[�w%ھ��3>��?��=�����ܿ���x�Q?H,J��Z(��	������54?PXg?%\�>��Ǿ���t8>�^T���=����=i�⪄�
�-�Q >@)C?��f>"u>e�3��d8��P�|���k|>=36?涾�B9�2�u���H��aݾ�GM>�ƾ>o�C� k�������iui�|�{=gx:?A�?�3��bాԯu��D��dOR>n<\>�S=�l�=�TM>�{c���ƽ�H��c.=��=Q�^>?�>v8>v0>R��>����qؽ�L�>�˜=)�K>�s?��*?9ԛ�Xӓ�����Ŝ��ڕ>T��>��>��>�h#�/R�=:��>EQ&>��6<����=�-��=;->�⽡�M�^<(<��6<������>_-)=}��'n5����<�~?���'䈿��e���lD?S+?c �=�F<��"�E ���H��F�?r�@m�?��	�ߢV�@�?�@�?��J��=}�>
׫>�ξ�L��?��Ž6Ǣ�ɔ	�0)#�jS�?��?��/�Zʋ�<l�~6>�^%?��Ӿ�d�>_f��Y�������u��#=t��>,;H?�V��)8P��>�6t
?j?`�+�����ȿQzv����>$�?��?<�m��@��r@��~�>��?�bY?�ni> U۾^WZ�P��>k�@?PR?��>�4�p�'���?K۶?<��?TH>Q�?G�t?V��>���tz.�����E���p=3*�:��>��>{����A�. ��)���qi�C`���W>�!=�U�>�/߽)ȹ�/��=�᝽⎪�=�{�L%�>�t>�NR>D�>'t?�>d�>J�+=�}���f��/�����K?갏?s���-n�b�<���=��^�_'?;L4?��[��Ͼ�Ѩ>��\?L?t[?No�>����;���翿|��IT�<��K>�.�>�F�>���$DK>��Ծ3D�s�>�ʗ>�i���Cھ08���(���E�>�b!?I��>��=�� ?�#?h�j>�%�>�[E��8��J�E�׼�>;��>�=?��~?B�?8����Y3��
��硿&�[�V@N>�x?�Q?v��>��������C^F�k I�;�����?�wg?�
彡
?�.�?�??j�A?�Lf>�f�5�׾�ƭ��>��"?����>A���!������?��?�,�>�LC�o��=�޼-:��� �?0�^?2�*?S���e\���Ⱦ���<3z��n <�:0;/���9!>��>�ʨ�[�=��>턡=�U���@�!W��{�=>��=�:�-i��C=,?^�G�ۃ��=��r��wD���>7JL>�����^?k=���{�i���x��U��?���?_k�?����h��$=?��?u	?A#�>WJ���}޾.��#Qw�<|x�?v���>���>1�l���_���w���'F��O�Ž����7
?rR�>�?���>��>݃�>���	���*�buʾ�BL�"�.=���G��&�����w.-���= %��`Շ���Z>���-%�>�I?���=&Nn>0�?
�s=���>z��=�N >gP�>���>��}>3$�>z蔽�ǽ�!R?�a��y�'���辣f��~�A?�[d?]��>�i�/������7T?蕒?�S�?��t>�h��+��l?�f�>�!��28
?d9=������<&����2��_���
�I�>=Fս:��M���e�_�
?oO?���)�̾X<׽��L�n=�M�?a�(?r�)�U�Q���o�j�W�S�(��:h�Ag��}�$��p��돿w^��W$����(��g*=��*?b�?�������$���&k�1?�8\f>b�>#�>O�>�sI>M�	�g�1��^�|L'�n����O�>_Y{?���>l�D?@n:?|kR?3�D?ŏ�>���>�乾�{�>rj��~i�>��>�:?i�"?�7.?Q�?�V'?��`>�#�������sھ��?L�?�?��?���>ޅn��.��L���'�� ��S���Ą)=_1<0����S�\q�=��S>JN?����8������6k>7?�a�>^��>��������<�>��
?�^�>�����{r��N�gS�>��?� ��2=/�)>S��=�+�������S�=��ļ��=�݂���;�D�<�׾=���=�x�.��H��:V��;�Z�<� ?�\?�>�>i"�>�x��;V����Vֳ=�[>3	V>��>��ؾ�<��c���f�D`|>��?Ws�?Lf=�3�=J�=�	��t𼾊n�#���K��<ۚ?(m"?2CT?�?�=?
V"?ѕ>������LƄ��桾{?�<?g2�>A�8�ݵ��)���_�B�4�;?�&?�����E�.H������`�;!W>4Kd�~y���ʿڔ����>�� Ƕ�H��?cް?i�D�A��S���q��EMܾ�?��>ճ>��?��.��cl������v>�?4?���>��E?oI�?��R?���=9�2��ε�ܓ��.�[��ܥ=(FJ?�c?Uӗ?"i?��>�b=�D����n��JR���+ؽt����ɯ=>d2>��>��0?E*�>���=u-%�_��T4��&�">�� ��>�>�?���>�0U>]T�=mL?��>�������N����4�Qa=P]?�u�?��.?N҄=�O��&��#�2L�>XD�?���?��/?����ڵ�=��< C��(#�2�>��>�Iz>�u$>S��<H6u>կ�>�H�>��'��=��h�=�ɇ%����>SmJ?SP>�t��$r��t禽tJ
�P�>���.��Q*��7���H ?�S�
K�>�޾;� ��'c�iq��i�������j��Dw?�S(>꫏<��'�|(�%w��Wg�;8Z��,�=��?=�a#��>т��^<���S*=�_*���=�)=� þ�lr?��J?�\0?��7?�"�>��>;𙽹�>�}��]F?��6>�M�J�ʾ��5��Ǜ��:���K����ξa�_�����>Жr��=J�0>��=�<�7�=���=��=k���л�<$ԯ=ԣ�=i��=I�>��$>*!>�6w?W�������4Q��Z罤�:?�8�>h{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?Dti��d�>L���㎽�q�=T����=2>w��=r�2�U��>��J>���K��=����4�?��@��??�ዿϢϿ5a/>�8>J>��R��P1�>�\�Lmb���Y�^�!?��:�� ̾ &�>hI�=7�޾��ƾ"�0=�C7>"�c=���Q\��ʙ=:�z� w<=��k=IƉ>�D>�^�=��"��=(�J=X�=�O>k��S�8��F,���3=���=��b>��%>���>
?$�?<g?�`�>D:½�O����ž���>����>|�0��[>vPQ>y�2?�<?�X?{d�>�	�����>匱>K:U���I�g'ݾ�(ݾ��=�އ?֊?���>�"����I����-�����?(?��+?���>�#^>p9�A��o%���,��΄��10=���;��t��޼�k���<��1=� kۻ-�/>=η>�a�>ʶ^>�l>�a>Á�>�^>��=�ڲ=bI��[�S�񁛼�:�<ȹܻ��K=}��<[�=W�L<C1�Lk=f#=E@�<�Ĭ<0a�=
�=���>�>���>R��=�����/>.���O�L��z�=����<B���c�}m~���.���5�d�B>o�X>j��������?˴Y>0d?>d��?a-u?| >��N�վV@����d��R���=�2	><��y;�r�_���M�ϺҾ.ھ>]��>�pr>3́>��)�7׉��;>ڕI���w���/>��V�f0�;G��=)�q�N���3���{~��,>v�J?[����=_b]?�%"?´�?��?��M�䛾C!�>.�˾��=���4��=�x?�i?�o"?%�C?`7��}@N�HC̾H������>'3I��O����Ѩ0�@������]�>Vɪ���о��2��b�������B�F'r�@�>�O?2�?[�b�6K���JO����酽�R?Wag?;/�>�j?�R?�)������L���ҹ=��n?��?�)�?��
>�P�=-����p�>��?I�?Q�?}�m?�zK�hk�>z>5���!>銸�� �=�k�=���=���=�	?$�?��?iq�����S�:�龟nb�Z�)=.��=��>X��>�(v>ـ�=CE�<'#�=�S>�U�>8��>5�j>S�>�w�>�Å�!�>t?of�=auc>��?p�1=�1l>��/��>N9>����uD�CL={�0;����>%s�=��=���>(|п�ѝ?�9�=���.?�f߾���z@>���>Z�n���?@ջ��3�>j�5?i�>�>:N>֨\=�ѾGA>���"��FC��Q���оDz>�뛾�,%���	�Z��S=L�����fp���i�a8��E�>��ֺ<PN�?�l�� l�o�(��)���?��>�7?>���������>��>�ˍ>L!��&>��m�����⾔݋?�V�?�2c>���>��W?A�?��1��2��QZ��u�>�@��e�Op`�s΍��{����
�k���ն_?��x?�xA?�o�<�!z>q��?��%������>�>V�.��;���<=��>�'��dE`�czӾl�þ��	tF>!co?��?;?�uV���ۼ��=B�C?��-?��g?_<?kV&?��	�S?A�>:s?K�?x)?գ$?0�?b�>�(>��=/�_<��L��'a�O�ý)G9����<� =�=���9ئ<���<�Ө����!�c��-<�Lf�N�<��H=4e1={�~=�ި>-!Z?̪�>�Ō>*J3?�F��P3�e��_/?�g$=7%p�o*�����4�����>ewj?��?�CZ?PkY>Q�<��7��>.�>�93>�_>�m�>�Dܽ�hD����=}�>A!>�i�=��.��~��
�Ǌ�XA�<�b>W��>|dx>�`����)>r���^nu�
Qh>q�P�/H����O��F��0�~s��r�>��L?�?��=�澤t����d�E+(?�X<?��L?HV?c��=��۾<$9�J�I�5��׎�>#��<V�	���H���:�:�:9�x>|�!e��H�>����@���F���R�G���%�(����>��]�`��㡾��W>�
�<�K��/���+���ק��C?��5>"O�����������j>>�t>{��>	)����<�gRD�#վ9_-<��>Cy�=B?۽�L��{O�q���Y�>��H?�@`?R��?X?l��7j��0I��\�R ��L���+o?	c�>�]?�O>Mn�=���I����`��K���>6�>9��A�>�z[����ʾ��v��>�!�>�c>Hu?IZ?��?�zi?�*1?I< ?,ߝ>$M������5�%?Ww~?�P�=��ȼkD��"�[1����>J�?l�Ƚ'��>}�?��(?R(?q�N?<?/�>���2����>(/�>��L��?����=ŪU?���>�CZ?�iY?,�.>L0������%�J8>���=Y�?7K+?�3	?�a�>�7?y`%�?�S>��?[:?ޱu?��\?J}�>'�G?��>L~?�p���>u�c�گ&?��W?p	x?"}?���>3Z�<���迬�����(�����<N� ��6=���CL=��=�l����F�F�F&���2��y��=x;�&j�>p.t>ٕ��Q1>C�ľ�Ո�[lA>9��������i(:�⬶=F̀><?���>��"�QO�=�Լ>9�>U����'?��?��?$�D;��b���ھ�kK��6�>XB?���=�m�{����u�iMl=�
n?�{^?iW�S�����b?F�]?�g�7=�k�þ �b���x�O?K�
?"�G���>��~?��q?'��>	f��:n����pCb�3�j�Ͷ=<q�>mX�`�d�Y@�>��7?�O�>��b>,�=t۾�w��r��,?7�?�?���?+*>��n�4�a�ᾍ���&a?���>W+��ݍ#?㡃�/�;F���=K��оS��e����腾�~����]�����r�qG�=��?��w??�r?��W?��?Z�eZ�jۄ�}�X������2��v;�Ox,�!W@��xi����7��J�����,=�a�4WI��S�?��?�a�<��>�$�����ž*>"�����ٽ�:%<m�м3�A=Pf�;0p�+O�2<��9�?�Y�>�\�>4�5?8R��8���,�UC�ܖ�V%>� �>���>�f�>+����YD����}�Ծ�K���	��x>*�`?�P?��m?>���(-��[���e � ��{ɬ��]M>=->��>�@E�������~:���m�ȳ�m����S	��gX<S�-?w��>=�>6t�?�}?y����񨾆,u�n�=�ReC�Y4�>#�f?���>��>�����B�[�>�m?W�>3�>�+��W�!�{�y�ʚ��eB�>T|�>~�>)th>�)���\��ꐿ�z����8���=�g?����d�&�>gqQ?Q�<�|�<���>�r����w��xh,��j�=vO?Na�=��F>�㿾^
���x�쌾$O)?��?���h�(�B�{>Į"?���>m��>E�?Uu�>$����?::�?�_?�tI?T�@?�Q�>��#=�e��%�ǽ�j%���*=�I�>��[>0t=Z��=���V�W��`!�<=�!�=6Լ(챽��<Xoü�h~<��=B{3>l�ݿP�Q�Cؾ����t��
���!�ڽ�́�|4��e橾2�d���~���P|O�aVN�H����}�7o�?р�?��ƾܐ��ߑ��ly��N��+�>(G������Um�F�|���}p���0�G�I���h�ij�?9?�(��?�տ�����b@���?*:?�s�?������F���=��G��Y=�1��K���mٿ0e�0^?���>����l���P|:?���=ĉ|����>���*�)��,�L?h�?/��>p�b��N��Y�ҿ�,&����?�I@b�@?l(�Q��f�E=N�>�q?0�>>�{1��������V�>1m�?�h�?m�]=Y(W�V���{md?��;�hF�qs��J��=���=�Y�<�0�15O>�h�>�D���@��7ڽ�"1>1�>��$��3��a�\Q�<w�]>��н�蒽5Մ?,{\��f���/��T��U>��T?�*�>S:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6�񉤻{���&V�}��=[��>c�>,������O��I��U��=p�DH����-�;F�"�=/�=Y������u�ٽ��G>}.5�>sS�ǟ�����>�`e>ܩ>�#�>o��=F��>тa?Bq??�z�>�I��S��=����T�ʾ��T=Me��_�>1���ω�=�ʱ�1PT���ھ�G��U��
�7u׾C�"��Q=+9T��ߥ��Q־�K�y�O����>D����S�{ք��I#>?���<$V�CtŽ�����V�Ɔ�N�?�y`?薿s�K�0�I�Y�w=Ǳ�=a^\?a�v����WѾ�ԕ�����`��B�Y>��;A	%���k�\j:�'c0?�??�z���ڏ��z*>[b��l6=]r+?�T?vd<ݡ�>��$?Q�'���彔$[>
c5>O"�>��>�J>������ؽ�+?��S?�E�t��㬐>f��Z4z���`=�>��4��(�Ll]>X��<�쌾8�A�����:��<-&W?���>��)�f���L���*���==ɭx?`�?;�>�uk?�B?�ڥ<K��]�S�v�W�w=k�W?Gi?��>�H��e�Ͼb���Ա5?��e?��N>*jh�e��U�.�xP��&?��n?5c?�J���p}�������Nn6?��v?�r^�Ls��T��6�V��=�>�[�>���>3�9�/l�>$�>?-#�aG�����4Y4�Þ?r�@���?@�;<�����=s;?�[�>;�O��>ƾ4{��܃��C�q=�"�>k���,ev�����P,�Y�8?ʠ�?���>����[��q�(>?�����?�	t?�F���C�=`���$t��v���1�To_=P}��G�X���ɾ�N+� ~�����Qо�Qy��
>>�u@Qs��/��># Y�yѿ�̿�Α��߾��:��>��>*5>+ؾ�9�v�o7\��mN��
6����S5�>sL>�O��!z��T�{�I;�J��]��>k]�9�>�T�Iӵ��<�;<㐒>&d�>�R�>@a��L����?����)ο͞����9�X?�V�?�p�?]I?��3<��v��y{�j� �r"G?8xs?��Y?_�'���]��5�6�j?�^��U`�܎4��HE��U>�"3?�C�>�-���|=�>5��>�d>�#/���Ŀ�ٶ�S���*��?��?3p���>���?�s+?�h�8���\����*���*�x<A?\2>������!��0=��Ғ�̼
?�~0?V{��.�T�_?+�a�M�p���-�Z�ƽ�ۡ>�0��e\�EN�����Xe���Ay����?J^�?d�?Ƶ�� #�g6%?%�>`����8Ǿ��<ʀ�>�(�>�)N>�H_���u>����:�$i	>���?�~�?Fj?��������U> �}?�$�>C�?N��=]e�>�k�=����,��f#>.�=:?��?5�M?�J�>M�=��8�y/� YF��CR��%�h�C���>��a?��L?�Jb>�$��:?2�!�xͽ[X1��R�AX@�F�,��߽3+5>��=>i>��D��	Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Va~����7�f��=��7?�0��z>���>��=�nv�޻��X�s����>�B�?�{�?��>"�l?��o�P�B���1=8M�>Μk?�s?�Qo���i�B>��?"������L��f?�
@u@a�^?*�ؿ8���!Z�/:��Y0��yb<ɉ	>y^	��<�=k!F=���<�$�tU<8�>|��>��8>(*>_m#>dP=>	�����]f��}Y���z,���!����
����]e������4�پe1�oP��7����㓾Qm�����;���=D�T?ܙP?�o?A��>t^_��� >-���@�<�N�'��=}i�>+A4?��I?\X*?���=����1b�����񢾠���v��>;8>���>�p�>� �>�?w< �8>��?>�sw>T��=U@=0�<H��<��E> {�>���>
�>��i>W��>/��������0���%c�1zĽo��?�˙�*�;�������h��5���=��?���=п����ٿ�(���Q?"pv�!�%�q��j���?ss?��>U=��֑)���x>˚P�C|�����=�ݚ��ū�o<��lp>v�<?� d>w�n>�~3�$�9���M������
x>Gu4?θ� 11�Lv�٥E���޾��T>�_�>�6�S�������~��0e�nz=uq:?$
?�G��o����ns��q��ظL>��T>��)=�ҿ=�LO>��m���ҽ�sB��0=*S�=*OU>��?B'6>���=��>�:���B<��`�>G�>>f�*>��<?��%?o���y;���������̄>�P�>�5�>x��=��>��[�=���>�UN>6C��9M�� ���6��_@>�N�A�\�
�H�S��=kz7�w��=(�_=̠ܽ-K9�"^b=�~?���(䈿��e���lD?S+?] �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�-)#�jS�?��?��/�Zʋ�=l�6>�^%?��ӾMh�>ix��Z�������u�K�#=R��>�8H?�V��"�O�^>��v
?�?�^�ᩤ���ȿ4|v����>U�?���?j�m��A���@����>:��?�gY?noi>�g۾3`Z����>λ@?�R?�>�9�o�'���?�޶?ӯ�?�Wh>1�?��{?���>MĽ`�+�Uÿ*m����H��k��'��>�u.>h�*p5����_���{j�)�/�/�=f�=ϋ�>�ߒ�����~�=Z�]���ܾ���>漘>��>��>�y?9�>N&�>;qR>����e�����v�K?���?���j2n��M�<���=$�^��&?/I4?�c[���Ͼ�ը>�\?X?�[?Ed�>���*>��迿�}��⫖<�K>v3�>"H�>�"���GK>+�Ծ5D�p�>�ϗ>r���Y?ھ[,���^���A�>�e!?���>uӮ=� ?��#?ڔj>�(�>�`E��9��/�E�
��>l��>�E?M�~?@�?+ӹ�?[3�{	��H硿8�[��:N>�x?�T?�Ǖ>'���߂��N*E��)I��钽ě�?�tg?$I��?�0�?Ĉ??ФA?k0f>9��sؾU���5�>��!?�����A��8&�����s?�J?���>����ԽxAּ̺��6��P
?\?R>&?L��Ga�~�¾�(�<�l �>�N��,�;�MI�<�>F>:��[г="�>r��=��l���5���m<�a�=^�>�={�6�����2=,?Q�G�ۃ�S�=U�r�xD���>"JL>�����^?l=��{�����x���U�� �?���?^k�?g��(�h��$=?�?G	?m"�>�J���}޾�ྑPw��}x��w���>���>�l���G���ԙ���F��!�Ž�����?���>��?wR�>>��=��>�"�i����\�}�ؾ�a�30�-LI���S�D�7�h̲�,����J�]㹾�ᶾ�U>}�ɼy��>��?�~�>�.d>,��>���=Q�K>T�=�i>�6�>
�>��>p��=�*�^�<��KR?$���$�'�B�������2B?;qd?[0�>�i��������ހ?E��?Zs�?�:v>�}h��++�Zn?�<�>����p
?eR:=t?��V�<qT��T���4������> G׽�!:��M�tof�j
? /?���T�̾~9׽�K���3p=�M�?��(?/�)�d�Q���o���W��
S�����nh������$�rdp��揿�g��:����(��(=o_*?�2�?�y��c���Qk��N?��e>���>cl�>뢾>�%I>q�	���1�k^�W!'��僾��>�{?��>DZD?t1+?�M?��:?嚾>��>�^��f�>AZH��{�>�Ҭ>O�I?�0?�	(?'�?��1?�>�V��|�\,ھӷ ?qI�>{�?���>�>�*����J @=S����Ͼ���G�0��\>_��<��=�%>�_>�]?]���l8��[���bj>�7?S��>���>rE�����(��<��>��
?-��>����6.r�L�%G�>e��?��݊=��)>%5�=�s����L5�=������=� ����<��<��=�Ȗ={؃�H�����;��;H�<Eu�>��?���>�D�>w>���� �����i�=�Y>�S>�>8EپR}��%����g�o_y>�w�?�z�?�f=.�=p��=|���T��f���������<�?�I#?�WT?䕒?��=?�j#?*�>�*�M��S^�� ����?ܜE?$��>>=���5�ǿbsk�gm:?��I?fE��(������ʹ�/hվT�>Q�Q��蛿��˿U�(�A��>�u�����p�?�ȸ?�F>L�k�Z�&�V[��c�ܾ�B2?�#4?��>W�
?a@���{�?��<�>(?gI?��>A�K?���?�O?�Ώ���)�l����*��s�d�T�>��C?(�?���?�{?���>�d	>6HS��@�������g��|�]�3�,�b>Qc>|x�>�?ܭ?��g>2,��-�:���d>d}�=��?��?��>��>\��=��G?���>�E���V������K��c�:���u?*��?ˑ+?{=�n��E�?����[�>�e�?��?/F*?۲S�0��=�Kռ7�����q��>?��>�!�>~ד=O,F=9�>���>,��>F��`��l8�a�M��?�F?Qٻ=r�ÿ?����6����ξ���=p�#.���c�:N��#R �`yվ����k��`Ya���t��W��v¯�{&ƾ��̾nX�>[G�=�)�=�#0��4=���-0������j������ð����=�R�0ɫ�F�4�Ɣ<�V�=ȟ>9��3ľ�d{?ϸI?`�-?q�B?`�m>��>�H�cx�>=꘽a�?dMM>��;�@��/>8�!��Z����Ͼ��޾0[[��A��I>���p>sU$>�<�=]�<�N�=��==�%��r	�<ݵ�=-�=�>�=��=Q�=�>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>v�(>Q��=)4I�
?���/��皾\�m��[?@�A�9���J�E>�&_>�&[���䒺z'K>���<?�#��yb�e��=��#�Cܳ=�,;�Mo>u�0>��o=z�ٽ�ͣ=�=���=�yw>���&ca�%Z��tj�; ��=dn>%�>��>'?�e2?��d?S��>D6M�}�������+�>��=.�>`�=]�>o�>�7?�+F?��??���>�2=�T�>��>d�5�<kf�F�þ����#;�=�p�?6&~?��>ǅ�<�ۉ�O�"��>�V޽��?ц.?ό?_�>�T��^ӿÃH�	��j�=���<pħ��z��I�˽�i��'X��������=I�`>���>.͢>{ܫ>m�h>H�Y>��>��>&y�=��y�&���\f�>b`m=�1缲�(�=���̰=}f,��N&��̏<H����q`<YW=p$>���=���>�;>��>�y�=����?/>P����L��|�=^C���*B�1d��I~�W/�m6���B>r7X>To���3����?�Y> r?>Є�?ZCu?��> �&�վ�O���Ne��bS��ָ=@�>��<�Vw;�lV`�}�M�\�Ҿ:��>	C?�ܚ>�[>^�E��c}��o��ȗ�cB��1�=Т*���Q*��j}�uG¿�%����o��~Y�l�\?Λ���=�m?�DW?���?�w?���o����0?Js��O��&�?o >,����>�'?8�G?q����s��H̾~���޷>j@I� �O���1�0�'���̷����>�����оU$3��g��������B�
Mr�G��>�O?��?�:b��W��+UO����^'���q?�|g?/�>�J?�@?&��"z�/r���x�=�n?���?8=�?*>��>Oِ�7L�>�4?:ϒ?�ё?h`n?�n�.(�>H9=e=>�܊���"><�=�ȵ=�c>(�?��?\�
?����І�÷ܾ���8�X��Ʌ<�;w=�mj>��>�B�>Wi>Ғ=�$�=8d>`�>�a�>{~> ��>Y(�>��{��
�;�?S>��>>�`?f��>��)>�=�^������P��b��c	O�����5l �j_��7�B��̓���>:޿9�?��=�ξy�2?�<���F��F�=ۏ>�p½0?����|�>�
?q��>��b>8�7="�><Ӿ�Z>����!�yC�=�R�j�Ѿ�	z>̜�4}%�V��h���I��﴾���r�i�>*��q8=��Ը<|=�?R1����k���)�U_����?�D�>��5?-ǌ�k]��~�>�S�>�h�>�/��@����֍�Ƅ����?��?�;c>��>I�W?*�?��1�E3��uZ��u�N(A�&e�,�`�~፿ ����
�e��0�_?��x?-yA?>O�<.:z>K��?��%�1ӏ��)�>�/�)';�F?<=O+�>�)���`�r�Ӿ��þ�7��HF>p�o?.%�?TY?'TV�ڜ$=�_^>�5?��8?(X?« ?f�:?B���(?gY�={U?�]�>��6?�?T��>��>>�)�=�b�� ���K�d����i�F�=��zy�� �:�h=��9=�e�:�}ŽE5�A<�i2Z�����؈=$�n=;ǃ=;/�>�,]?Z��>�2�>|�7?y��u7�?����.?�==�h���ˊ�Y⠾��|�>n�j?�f�?�Z?��`>�A@���@�;�>��>�$>xl[>j�>.)��NG���=P�>�i>.U�=�4A�Xw��K�	�(�����<f� >_��>"|>���٣'>r��/6z�ٛd>�Q��κ�o�S�n�G��1��v�a�>��K?�?���=k_龏4��tDf��.)?�\<?�LM?��?��=��۾)�9��J�IF�z�>�ת<�������#����:�#��:պs>T9�������V>9G	���OUh��>M�?I�z�'=�e���=$���ɾy���"�=��>ER��p ��1��O�����I?�D�=� ��xFd�CU��8�>`@�>�<�>���ѝE��C�����=֗�>�p5>*������лB���Ʈ�>BIN?Xa?t�l?����f;^��_����$�m���(��?4�A>��?	�]>���=�������{��|�]��W�>[��>r�޾�r8�(�d�q� �u�(�� %=ʈ�>&F^>�U$?#Y6?�,?& r?U�?j�>e�>�X�4��#?�Z�?��=�����x��/;���H�E��>�+?H1Z����>Ͳ?��$?��)?��S?B�?>g>�t��@DD��U�>2W�>%V�Z���TQ>�xE?q'�>��]?[�?)	>�<6�����I�w���m=OX>�|3?�k?�#!?
��>ؽ?Hо}�>�4?���>Oc?�8?Om���<?8�>V!?P#ؼ��O>6񀾆+?K�K?pu?a�O?���>�a=?1A��=�E�(��9R��u{=��i=�)�=���'�I�q<���27=ӗx�Lv���A˼u��Y��<�<j�>�b�>��e>�����x*>�������zt8>�?s<U���h����7�"g>��>G?�:�>i6���l=�A�> ��>m���,?�?��?��d<�"[��J쾆Am����>N5?��=�p�έ���v���x=^�o?O�O?�l���� ���b?U�]?�f�=���þE�b�0����O?t�
?K�G�!�>1�~?F�q?���>�e�X:n����yCb���j�8ж=�r�>�W��d��?�>
�7?�L�>h�b>�#�=�u۾n�w�Or���?��?��?���?�(*>v�n�4��辫`��x{^?��>�%��C�?�,��<����p��-޾]O��Nn��L���)^��j4>������6�4c�=�?�}?��b?7�g?e����X��i����P��g
���gVT��D��G���`��:��J(�����k+<� w���>����?RO$?EL/�fH�><������^;�1?>៾�P��T�=��i���I=KK7=��n��%7�{�h?!�>���>B�=?�`X���;�'25��;�`���G�,>�آ>��>�5�>�Zӻ��'���Ľ��ʾ;����o�E�u>Ђc?_:K?��n?F �� 1�fZ��G� �c.��O���=C>�	>���>GhX�`���%��>�+`r����U2����	�E~=	R2?�c�>�.�>,�?u%?q	������ w���0�-x<�:�>CFi?B��>��>� Ͻp� �̑�>�l?-n�>��>�W��7i!���{��|Ƚ���>�A�>��>��o>*�+�)	\�]f��-���A9�S��=�h?����ica��ʅ>��Q?|1f:#O<��>�x�x!��F�g'�1>N?#�=.=>L ž�+�{{����)?I�?(l��H�(��xx>�!?F�>���>��?yv�>w�����:.?+�]?
J?.A?�X�>�-=80��L�Ƚ�%�>�(=2��>�^>fzp=C�=XS�D�]�3����M=��= ��Q��[�<M���!�C<�o�<>u3>�wۿ��K�X�۾m�~����	����!_���ሾ���s%��q���N|�����T"�VS��ld�:&���Km�y-�?=��?�[��gd���ݙ�n��Ze���Z�>QSl��Ln�(���@K��Z��}�޾gs���`!�w!N��"h�Of���4?dQ	�.Cǿ���4�S??�*4?Yjq?����O���B�'u޽r�s��F���L,�ܫ���ڿ"���]��?� ?b���|8��?:"�=^̀=��?R�9=O\$�u�@��E?��?��>�頽x ��2�����P��<�?��@�lA?��(��-�KW=�0�>�p	?�U@>؆/��������(�>�i�?׊?�-Q=oW����cGe?�<�/F��8軻�=�j�=�=a���H>깑>V����B��'ܽ5e6>�k�>m �b)� �]�u��<�J]>��׽	���5Մ?,{\��f���/��T��U>��T?�*�>W:�=��,?X7H�a}Ͽ�\��*a?�0�?���?%�(?8ۿ��ؚ>��ܾ��M?`D6?���>�d&��t���=j6�=���|���&V�{��=Z��>c�>,������O��I��V��=�f���S��i�B���?�h��>�,̽�@���m�j�o�=J�ܾ*Lx�MC����>���=��m> �!>VU>ф!>�K?��2?���>	���ɥ=���X���E~μ>�&���ͽ�Rƾ΋�=�2{�dEӽM�ؾ�w��Y.�\�����2&����=�j>�����yþ�U�l�E��U�>�3>����L������=�Z����=�]2�^x��֧쾵%(�߶x�zѓ?��?�����jz�<=�A#�>��+���/?GJ=�1��˾������"���S�Q_��'Z��&��nG�J�`��/?�,?�뻾>b���)'>b���U=A+?��?�*#<:"�>��#?�%�0��^�]>��3>�M�>t��>^Z>
`��P�ؽ,?��S?���X ��R�>�K���~��=y=�>�L5����4+T>怘<�����u�9g���-�<(W?���>��)����a��v�=]==�x?�?d-�>zzk?��B?��<ff����S�K �]w=��W?�)i?Ⱥ>�����о�����5?&�e?4�N>#bh����#�.�U��$?�n?�^?�j���u}�������m6?�v?�r^��k�����t�V��K�>r]�>%��>��9��y�>��>?h�"��A��1����P4�?T�@���?v�=<�b�s��=d6?Pi�>��O�Bƾ����Q���%?q=V#�>�e��6]v�_��u!,��8?ڠ�?4��>������}*>V�w�4�?'�~?�ƭ�GXE��S!�t�V�������L=��J<:L���Kپ��"�!rϾ�v�hqž���>�h>�@�=	�֯�>�Z��Ϳ�|ӿ����B�Ҿ���T�?�>S��0����Q��>K��xI��K^������>��>�֔���u�{�Љ;������>G����>�:T�9õ�����w�<<j��>N�>lO�>b߮�N���[��?;=���οO���8����X?nP�?4J�?��?+K<�w�F{��o �oG?��s?K�Y?6%���\�CZ9��k?����aa�DI5�ǍF�{,S>��4?ß�>��/��dR=�>��>�>�-���Ŀ�����쳥?�5�?��8!�>�/�?��-?���ѿ���=��$�(��V�B@?�7>!＾8�!�;3;��I���
?F0?���,��]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?|	�>�ք?$��=��>�c�=ɏ��Gu��O">W��=jwE�g�?H0M?���>�+�=67���.���F��R����<C�C:�>�(a?�VL?KX`>�Ÿ��K�~$"��ѽ�/��-̼�6E�	�+�kὈ�4>*@>ļ>� I�c�Ӿ��?Lp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>A�Խ����[�����7>1�B?Y��D��u�o�z�>���?
�@�ծ?ji��	?���P��La~����7�z��=��7?�0�2�z>���>��=�nv�ܻ��Q�s����>�B�?�{�?��>�l?��o�M�B���1=-M�>ǜk?�s?j[o���o�B>��?�������K��f?
�
@~u@_�^?)i߿���r¾@款�'>�>�8�=�������y[:������tѼj[};,4�=�k>w�>N�>�\�>�]>���0!�^A���J�����O۾���z��(=-�6�.�� �'�����9K=��ֻ�����Ծ�]d�� �>VXV?ƕO?�zn?<�>���v�>�N����<�2�t��=�b�>��4?G>7?v�-?�Y�=y���bZ�ˁ|�j����X���	�>�Q&>��>�x�>���>_ݦ�,�$>Pr>��{>&r4>���=���=��?;[�?>�p�>��>_��>&�<>w*>��������wh��2q���ԽIڡ?�ƛ��;K����������z�=IT+?ʸ�=	@����п֭��H?EP�����S�+�IA�=�k1?��W?��!>yD��3x���>3���1k�f��=�����v�0e*��I>�/?��f>1&u>ُ3��[8��P�ux��5+|>>)6?���S9�F�u���H��[ݾ�9M>ž>��D�Xp��������ri�pt|=�q:?��?�Q���ܰ��u��b��P.R>�D\>��=���=�TM>N�c�нƽ��G�[I.=�Q�=��^>9.?�7=�L[>0
�>¦�=X��x�>)��=I�>\@<?��/?���=���<3���)%��>f!?�}�>��3>-�O��=�U�>�>$|�<~i��1F��1��s��K�<�yp=nT�����<���<-l>��U>|���9\X���ͽ�~?���'䈿��e���lD?S+?d �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��F��=}�>׫>�ξ�L��?��Ž7Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�<l��6>�^%?��Ӿh�>�r� Z��"����u�K�#=��>�9H?�V����O�
>��u
?�?�]򾵩����ȿV|v� ��>��?���?��m�q@��@�Ҁ�>���?�gY?pi>�f۾�YZ����>Ի@?�R?@�>7�-�'�_�?�޶?���?mJ>���?w�r?y��>ba����+�R����/���s�<o�:fɓ>)��=����[r?�Z���Y����j��b$�<�5>:$ =��>�S���;��4��=_���<����ѽf�>*��>_�>��>D�?�L�>O�>��==B��{ψ�l����K?s��?����1n��-�<˛�=��^��%?�H4?u�[�m�Ͼ]ը>�\?���?�[?�c�>��+>���翿�}��콖<��K>�3�>�G�>M$��-EK>	�Ծ,5D��o�>ZЗ>���>ھ�-��~���B�>e!?��>�Ӯ=�� ?��#?,�j>�(�>]E�H9��`�E�ļ�>���>^@?��~?�?ɹ�rX3�����桿Ò[��?N>!�x?�S? ��>5���򂝿L5F��H�	ْ����?�tg?�彵??2�?=�??a�A?�Nf>�w��ؾ]���8�>��!?����A�S#&����h?D?��>�U���ֽ��Լ���OK����?K%\?�=&?����a�&�¾���<N� �I�N��</ =��>�U>�M����=��>e	�=*Jm�U�6���^<�s�=㍒>���=�d7����=,?3oH�փ���=�r�BsD�L�>�6L>����e�^?�U=���{�|���v��C�T�<�?��?;k�?:	��ڜh��#=?K�?�	?<'�>K���v޾b���\w�T�x��t�V�>[��>=_l�j
�D���r���F��1�Ž8��@?	-�>�?:�?�=�w�>$=��#�Y!�3�*T��}��}�$�� <�.P2��5������&W�<h�ľ���b}>��C�7N�>'T?���>?�>�k�>g��=���>�2Z>��4>��b>�f�>�>�>�K<�	�=ߥ��M�N?]Fþ$����l{���@9?i�^?���>������Z��e/?��?U �?�Sr>��i���'���?��>9'u��x
?�=���<ZO=����D�?������V��z>�fѽV9��DI��dm� ??Z�?���zپ=K��~���\o=DK�?-�(?��)���Q���o��W��S�u���Ch��c����$�2�p��㏿�Z���%��X�(���)=+�*?G �?��-�(���k�6(?�	�e>���>b'�>��>uI>��	���1���]��='����
'�>�E{?Q��>\8L?fG/?�sC?�t?^�Z>���>�˾�?ä��1f�>+��>f�W?`��>��)?��?�-?�R�>�} �ļ��X��޺�>���>�76?��?��?x����m���j=�c�����gV��(�ӸȽ�h���!<�G	>'\>=�?m���5��=����c>�5?\,�>J+�>�����{�[�<Ø�>?��>T����[s���2��>5b�?�X��t�<��6>���=+Z�B���E�=����^X�=�:[�J�=��o�<��=�7�=MT�;�:;-0;���8g�l<u�>��?���>�D�>@��� �>��f�=)Y>�S>�>-Fپ�}���$��d�g��`y>�w�?�z�?�f= �=��=�{���T��I��+���)��<�?;I#?�WT?K��?��=?"j#?�>�*��L���^�����Ȯ?�p=?}i�>��0�����Y���C�P�>�8?��H?#ޙ�Z⾙)	����%��@4^>ʀ�2���ƿ?K����>su�Sx߻74�?^�?�ɽ�����Ǽ$�|q�<Ƴ�� ?�\�>�N�>W?7z���h��OѾ�>�g�>���>{��>S�Z?�`y?
G4?_�����G��Q������ם=*�&�Te7?0�t?^C�?YI�?�a?�S*>F�s����v=���@���Ð�<1t=��
=�O>�
%?�D�>S��>�䟾�k�z"0��T`>hf�=�4�>*�>��>�?�AE>=H?���>�7��.��[�� 怾d-���t?kא?[�+?Б=����<E�����PA�>�&�?�߫?�*?�O�Փ�=@;ͼr��Z�n�jr�>���>N�>��=�}A=�J>�a�>`S�>SD�����#8��A��T? �E?"d�=�ǿ�>��"�$�����>�z��~����<�x���{�>��0��D)ܾqE���j��oĝ�s2����A��r���h?�P>U�!>�f<�m�N[���=��=��>��K>Ѣ��+>�{Ǽ%�`�oM�p杽�y�=ȁ�=�m���ʾ��}?"I? �+?$�C?/�y>X>�<6���>�D���%?&(T>	L����&�9�����a����Aؾ:{׾A5c��m���I>'%H��f>QU4>\D�=Kha<���=�?{=���=�A����=5��=^b�=��=�s�=��>�>�6w?X�������4Q��Z罥�:?�8�>`{�=��ƾq@?��>>�2������yb��-?���?�T�?>�??ti��d�>M���㎽�q�=H����=2>s��=w�2�S��>��J>���K��D����4�?��@��??�ዿТϿ5a/>%�7>��>��R��B1�ca\���b�pIZ��!?:;��s̾�6�>+��=x�޾@�ƾ��/=Ws6>��a=4<�I$\����=A{�:�<=8ml=B�>�jD>��=�ı��ߵ=��M=W�=Q�O>mw����9�� *�H.6=���=�b>w%>Qy�>�?�/?x�b?`��><[^�T�þa�¾w%�>*]�=c�>,�x=&�O>7i�>W�6?F�C?N�L?���>��.=ĺ�>��>0(�
f�Q�������V�<���?݃?p�>]8�<N}L�u��C<�{*���5?N�0?�3?�e�>|2�L�׿} C��*�T�<�`���W�=c�)�w�ý ��=y[C�|�u��=iي>Xµ>L�>~�~>�t>�Z>6U�>�>*(>>p~A<h<=��ؼ�V��ѣ���j�����;Κ��j�!<�8R��v��C�~=�䊽<�M=�叽��4=K��=���>�C>��>n��=#��/A/>5�����L�1��=<A��s-B��.d��K~� /�SI6�]�B> 4X>����=1��j�?��Y>o?>���?FAu?2�>�6�;�վ�K��@:e��MS�굸=�>�<��t;��X`�,�M�=Ҿ��>��>��h>�>\>3�u��&��TŽ	(Y�jŇ=)���u(V�ɉ���7�Q��� ���-9U��#׽c=?�㈿��.=��e?�J?©�?�t?+{H�ʖ�o�>���������s��c�>6�x�@?��&?��?.��YI�eH̾{��t޷>@I���O����0�ڔ�	ͷ�T��>������о�#3��g�������B��Mr�b��>�O?n�?�;b��W��gUO�����%���q?]|g?��>dK?g@?�"��Pz�+r���{�=��n?���?=�?z>��>�W����>�?]
�?�E�?��k?`RK��-�>�<��G>\��ǔ>��p=��=��>�?�?Rb�>���*��O�ؾ|$;r쒾�����!;AΕ>��>��R>E>#�a;mu輽�>�ë>kj�>O��>K`\>IŃ>�3}�	�־�!	?~~�=/>�?�W�>�Y�>��O�,���T�H�;��$���k����,1��ܽ�p�=m��=(z�>��˿�0�?J���D����?�b���Ƀ�}�2>4I�>��m��A*?ۻ�=2�>V�>1�>݊c>��/>ݺ>�=���߉>� �'�L�C^F���!�Θ�i�1>��q������5�(z}�$���:�ɾf�&��<s��h����m��wo���?��=Sj��j�aB����? $�>.qB?CԶ��A���>�R�>veY>���p̓������c�̰b?�@9<c>��>��W?��?��1�,3�ZtZ�4�u�E%A��e���`�@፿����Q�
�~���8�_?:�x?wA?z7�<�8z>���?1�%��Џ�|*�>f/�';�A<=�&�>$���`�%�Ӿ �þ�=�`IF>e�o?�#�?�V?0WV��$���mZ>�b8?_3?Wo?��4?�(1?�抾�`?�kL>�f?R�?k]9?� ?��?�kU>�>]�E=]���m]�oZ���u̽���׾�<;�z=Ad�=,B��!=)ր=��i;�w�;������D=�����_���=���='�i=�ܥ>|I]?'"�>yѓ>��0?����/�M����/?:�=r�a�_`���l����>"mi?�v�?�2Q?bJO>�4���9��>^�>�^B>�zt>�E�>:�#�&�f���=N9>Y�">A�=�p��clu��@��N���]!<�l	>d?�>�~>�z��ŏ*>ƃ����z���c>��P�����OW�~F�,
2���r��8�>��K?ܴ?�M�=ǂ�
���oe�#�(?I�;? �L?��?뎛=m�۾�9�øJ�N��<"�>��<B�	��Ң��d���}9��z)�Zo>�㟾`��XC6>�c��kG��S���X�������+�6�G�=��&����o�����a>B�E�A{/��9��p���1I?��>|G���מּ,����Cx>�d>�ST>�F��V�<�E�����z��=�t�>�B$>��'��ʾL�O�_z�b�->j�2?0�m?l}?�ˀ�4Ov��x�iF�������;��?=��>֌?���>��w=�ͽ�����^�x�K���>h��>\���>�b���V(��d��Ly>!��>26>@�?��J?M�4?�&�?��9?�ݷ>}4�>C�D�Lc���%?Ն�?G�=\Sҽ��R�oj8���E��d�>�(?ZCA��S�>�b?�y?�C&?G�Q?�?m>#� �n@�r��>x[�>��W��=��y a>N2K?���>�3Y?���?�a=>H5�_K��ZA��_��=�>��2?3u#?�?2��>6^4?�z��S=�,0?%�?qPh??)A?|�>�%?W>� �>=D���S�>�]�<;j?��Q?4�b?�o8?G�-?{g�<��7=�Wɽ5���v��L�i��K�;�,�=1=@>nD���9�=@�=�!�L�һ���-gF���:g�@��>��p>_"���4>���4��*d@>�ڪ�pל��׍�"(2�/��=ޑ�>P� ?M�>� ����=�B�>ij�>�0�4�&?�?��?�M%;�a�i վb(=��ܯ>�@?@��=�l��o��۪v��\n=��n?֋^?��P��W��L�b?��]?4h��=���þl�b����_�O?D�
?+�G���>��~?[�q?B��>��e� :n�"���Cb���j�Ѷ=[r�>GX�S�d��?�>j�7?�N�>��b>�$�=nu۾�w��q��a?��?�?���?�**>{�n�R4࿃�	������l?ߤ�>O����E?�N���"���n��@]`�����7������8z�����V����Ǿ���8e<dw�>l��?�S?8?M0c�y�L�2Nl�%�����0�s����mP:�ރH�aY����������gP�w���ۥ�{2:� ��?�;?]*��
�>0��j
���Ծ�]>�Ig�q�<�1�=��F��=�ڭ=H���W�$��B很?_��>��>�:?w�'�["�3B@�m�L��ě�8t>�`�>�;�>+m�>a�ϻ�`����?����&T��8�B��3F>��X?�fH?'1k?w�Ľ
/���}��#��ݷ�3L��x>EEU>���>�W� H�����6� �f�C���
��&��*�<);-?[>}>L��>Ḟ?�??�ո��䬔���6���]��{~>�hd?�?���>Z������>��l?H��>��>=����N!�x�{�#dʽo)�>(ڭ>��>�p>B�,�'\��i���}��� 9����=��h?����W�`�Bم>�R?�Ҝ:]�G<l�>��v��!�L��N|'��E>�g?Dw�=�{;>�mžO��{��%��2�-?�?����|p��qo>�c#?��>1��>��?&Ԟ>{���_���?FV?9�I?-�C?���>"�=Q����ν1U��=�ц>$i>gQ=�ҹ=�����_�������<�ԏ=;�L�����>C�<Y������:N1�<��>��ۿn�K�� پ�7�&L�P���񉾿ݵ��3��s���r��B噾�y~�n��l;�R.Z�͢g��B��h�o��q�?���?�����E����������>)av�@p��㬾�������2޾B��/�"��P�j�Gtf��+?��^�)>ƿ�)��� ��A?�/?�xr?ʇ�hU3��?�i�+>��_��	=����'4��Dпڹ��h]P?���>]~�f$����>�b>��>=Qr>��U�u젾ϼx���?�3?t��>#R���ÿ-��\���%�?c@I�Q?tH��$�_o�=�(�>���>�� >s>潑��Ɔ�NX�>B��?��?l^(=�]�c�o�-�e?1L�=6���p.;K��<��#>6���*�K2�>X`>�9��_���� ��|>C7P>�,񽫂�;KI����=�{>�!�E=g�?�cZ��d�h<+�v���>r�T?z��>}��=}Q/?b�E�Z~ο�Y��9]?�G�?g	�?S4)?vR���[�>�ܾ_M?Gr6?���>x\"��*r�]��=����b���߾��T�;	�=z��>��'>�9!�k���MP������=����ƿ�$��i��1=1��_[�ȣ�Rg���JU�m���'o��罞�h=t<�=e�Q>�X�>�W>��Y>VXW?��k?�V�>�m>9������"ξ\���
��������-��o棾�6�y߾~�	���������ɾ��`�1F�=�aI�LV��Mz ��Sm�և5�-޺>v�ӽG!�d�������,��������1ۨ�
��n�}�|��\�? �c?G���zn��YE�XW�=&-;��?��� �¯��j��=27-���=Lh>��C��$��B^��7�o�4??t?3��5C���>q�����q=��(?K�?޷�=���>�?�.��F*K�WbK>E#>(;�>���>Y@>q��51����?I�(?~{�W���J�&>�}ھ����n�;p�>;�!��h�0�g>+�H�y�o����<�8�g�9=��[?eł>4�4����/��v�&��ʘ=��s?��?m$�>p�b?��8?Ɠu=>Z��<�M�*��!�=p�]?\�n?�v>8V/�O�¾v^���4-?ٵ]?�+L>�^���Uj(����r?�`d?(-?�me��*|��׌�8��X�2?w?�Q^����)#�E+S�#?�>~c�>��>��8�~��>��=?��%�nv��p}��E3��j�?�^@l�?�{g<aj��=�-?��>=.R��mƾE��,���Q^z=;��>�P���,v�S��T2-���7?懃?T�>�3��t�2鑻^ҹ�`!�?��}?�-~�4(:��C�0xp��V�}�μ��=���<�.�� ��C����6"����2�;�~>��@Yt���z�>4]��޿� ڿ}��_!ƾnMG�Ӵ;?v��>��^=�`H���Y�Z�s��d�N�A�NĐ�^Ѳ>�'�=��-��Dp���I���w�=s��>�e�;9��=�*>������M��r�z�>�l�>&n�>ΏV<��z�j��?:�����ο菿�� ��"9?M9�?V�?WP$?(]��E��Ha���w��$55?YRh?jfJ?��n�l!\�}ߙ< �t?�ܕ�e!v������6�0�8>Ч>?$��>dR�\)�=U'>c��>ˊX>�?+�w��޼���ɾ��?DT�?�Ӿ�# ?j�?��?.�������N˾,���I���/?�X�>�i��!��]+�����>=�:?]�U�bX.�ݶ_?��a���p�Y�-�dƽ��>��0��L\��������DQe�1���|y���?�[�?��?�����"�p;%?���>Š��SǾ��<�z�>�>r8N>��^��u>Z���:�|P	>˧�?Lv�?�i?����}���t�>>�}?��>C�?���=�d�>��=����vd/���">���=">>��?9�M?�7�>���=��8��/��RF�H7R�=(�q�C�o)�>��a?ׂL?�`b>�a����2�!�-Wͽ�31���缜K@��N-�\�߽�m5>��=>'�>�D��Ҿ�_?J��V�ؿb'�:�3?���>$?Ћ�Ns�����Z_?�B�>�)�������Y �V��?�
�?�?ڲ־�Gɼ?&>�N�>j��>�۽�y��	����Y7>�oC?ն�*���Uo���>3[�?��@Y�?)Yi�o	?��|R��UO~��m���6��,�=N�7?>��mz>���>Xת=Wv�X���h�s�׸�>�=�?
y�?���>ųl?s}o���B��72=L5�>�k?Qq?��e����a�B>)�?���}����J��f?��
@�o@g�^?碿����aǉ��t��徾"ZG>.Eݽ��>*�=<�Z�=�V�=������=@{�<ah�>��=D�q>��>��>=>B����c��ˣ�����W�0��W��8��o� o��M%�J�B�y��j���z�� 8e���<�?�	���;�MH�ya�=�%U?��S?ӯj?j(?��f�ǋ�=�u�E
M�-����>>��>Q!?K.%?mXF?r��=����jR��-x�[Ӆ��:B����>�1A>���>��
?ڤ�>m� <�: >�<>Ip>��=s�<��Q��<W�)>���>]:�>�1�>�l>��e>f ��׸�<&y��W��4e���y�?�d���V�Fr��戾羧@�=6?#�U=�v����տ����H?�-��������p�=�?�cU?"e>�)�����6�3>׌q�Ӄ��")>���gj���/��.�>�_?`2R>	Jw>��0�Ӥ8�&O��8���v>vX4?�L��S:N��{s�H�H���ݾ�}L>�۶>/���旖�.��-e��I=Bx9?�X?a�Ž�#���|�����d>eCb>	d�<�6�=!#Q>��#�N�ʽ��X�7�@=5�=�U>�?N_>z����D�>�Р�'����>q϶>Ǉ�>9C?��)?V��;Q�O�����9�����>E?�%�>�'�>�AZ��9�=RZ�>f_9>��;4	�c1L��ڏ��>���;�E��~ν��>�S%=�rQ>�z�=~�������'>*�~?���/䈿��`e���lD?j+?F�=t�F<x�"�7 ���H��8�?]�@�l�?x�	���V�Z�?�@�?�
����=}�>�֫>�ξ�L��?k�ŽpǢ���	��(#�^S�?��?��/�Vʋ�Dl�q6>�^%?�Ӿ�j�>:x��Z��}��^�u��#=��>�8H?|S��ĿO�M>��u
?�?�^�(�����ȿzv���>:�?��?W�m��@���@����>١�?-fY?Wqi>3j۾�`Z�玌>�@?�R?��>�:���'�%�?�ݶ?���?��H>��?��s?y�>�fw�^[/��/��ݠ����~=`�p;���>Y�>y���_SF�}����U����j�7���0a>�%=�;�>��(㻾�y�=����V��V�h����>Kq>C
J>�C�>� ?
=�>)�>^\=E��c����N����K?���?#���2n��O�<���=�^��&?�I4?#i[�p�Ͼ�ը>�\?`?�[?d�>/��G>��=迿7~��I��<��K>4�>{H�>I%���FK>��Ծ�4D�Kp�>�ϗ>�����?ھ�,���]��"B�>�e!?���>�Ү=�� ?��#?�j>�(�>�`E�e9��n�E�Ʋ�>��>�H?�~?��?\ӹ��Z3�����桿j�[�p=N>��x?�U?�ɕ>
��������ME��@I��������?�sg?zR�r?m2�?Ј??��A?(f>��|ؾ����1�>y "?����A���%�rT��~?D�?��>�L��e�սW�ؼ��������?��[?�&?���Z_`�[m�����<V��T����<��@�E;>d�>� ��~ʹ=�>���=�gm��5��CY<��=O�>n��=��6����B,? �G��ۃ�`7�=��r�`D�K�>�}L>�����^?zR=��{�L��pt����T�j�?m��?Bj�?�c���h��#=?��?p?,�>B���{޾נ�1w�ex�t�;�>��>^�h����ψ��`����?��+�Že��YW?p�>2w�>���>�~�=m�>r9��w8�����Ѿ�h�����73�i�)�������Rf����D���ȾW3����>�҈�Ò�>#�?Y|D>Cq>�.?c�˽"-=>�>E�>O�>4��=���=�3�>T)�=L�x�ƧT?�^ƾ1�)���ᾥʯ�B?�c?�w�>�5�O������?^��?�ӛ??vn>�a���#��?w?�p���?���=o�,���M<QU��ht��W'��뼛ۊ>���T�;��K�R�]��u
?y�?����|ʾ�_ӽ�9���o=�:�?��(?޺)���Q��o�C�W���R����Th�>a��
�$��<p�K揿0R����ӟ(�!� =\j*?�و?z3��:� i����j�;?�C}e>�/�>m��>�5�>t�J>߄	��!1�k�]���'��@���D�> {?1��>��N?L�<?u`B?pO?q��>Sf�>֣��h��>JEB���>���>B�1?U?`�)?�?�,?�r>�!���C�Rؼ�^3?�L?:?���>J#?Ɏm��M���<�-=�\O�FYZ��\���%=w����ҩ�i��<��R>uk?� ��"@�_Y��h>�	1?5��>|�>Kk��@�i��>=��>#�?$�>%� �|Jn������>fڂ?}s��	=��.>U��=T��z�;�U�=J�
�Ңw=��t�
��/V�<���=ͬ�=8��2*��:<�;Z�����<��>��?�1�>�R�>�x��n �� ���=�[>�R>�v>��ؾ�≿�����g���x>?h�?�F�?��n=q��=���=L՟��@���=��Ľ�NE�<�?E"?&�S?���?ؿ>?f"?u�>����蒿�񄿂�����?�~�>u?.���21���ſ�zs�l*?C�?G^y���_rN����j���R�>��I�����
���{j��T����������?f�?+��=cS���{�p�
 �""U?���>�5n>�k?ϴ*��])���̾�>E*?�/?b9�=Ω-?5��?=U@?:
>HH3�	W��T>��n�,�p�=��O?�!�?L�?��?/d�>�e*��@��q �C�����;�)����ؾ��=߲�>$�>0�3?X�>�7�3b���"<������	�+;�g>B��>ȸ�>�|�>g�>��I?��>������ ��9��+!^�'`�N7u?i�?�;(?z!=o��5�j� �y;�>���?�٧?�;,?��#���=j:��Ԣ���z����>w£>³�>�BJ=�E�<�>c��>]��>���/��,>��'��[N?ڸG?sB�='�¿�Np�B�N� ڔ�:��9:���Y�#���o�3�=�b������oN�7u�����M��)��r���2v�>�n=Z#>�H�=.�<�6мŨS<�=��=�b=bU���E*<��$�>v��F�+��
 ;�h��$J=Έ�OB��w�?�p;?�X"?�;P?��>"�w>9����<S>�O,�q�?k<I>�@4��Ӿ5�E�Io����h�>��F�ݾFD�޴���-�=���i�>�,>y�>?�=�>��:|�F==��<AԖ=�e>̜����/=ReB>�}>���=Kw?����#���dyP�ޣ�s�:?��>�W�=E�ľ�>??qm?>w򃿦���-�~?���?g'�?��?��b�/ޠ>7$�������=���X3>��=�,�c��>1�H>�U�u^���h�����?xO@��??�w���*Ͽ�0>:'>+��=�[D��%���N��ao�M�3���?O�>�5�ӾW��>]�=˾�!Ǿq��=W.k>��v=�j���^��4�=d�s�Ↄ=ʡ<��z>��.>�`�=�NϽL��=V7�=�{�=�L.>H�;�)���}]<��9=��=γS>_D�=>��>?ct!?��\?4�>�:E�����'¾_GZ>l�B=w�>���=K�`>�>hB-? �;?��??�	�>�v=���>�Ǒ>Ȉ7���^�&�ȾQ̖�\�>���?OX|?��>�����`�`�ص=�l�Ik?z�+?�n?�_�>FN���࿈A&�>�.�Ns��o�Q�a�+=skr�#�V�h ��]��}�tb�=}f�>�	�>$�>�My>8�9>�ZN>��>O�>g��<��=(���ꤴ<V��v�=�������<OżJ[��+C$�/.+�����m�;�T�;;�[<�X�;BE�=���>�@>w��>Hm�=�&���:/>]���N�L����=�9��0B�(5d�\<~���.��W6��]B>��W>؄�_4����?(�Y>h�?>���?CTu?��>���|վtP����d�s�S�g�=�>��<�l^;��.`���M�<�Ҿ8�w>hC�>o��>S�=�H2���a���=���ynm�K'�>���R�ĽA{��T�C�M�����=����??-�����i��n?�2i?�Ơ?�o?/{d�V�ξ��l>=����@B>�;��ཤ�(��=?��C?�!?����{=�W�;�޽��\�>m�A�]�L������/�����к�:�>L[���Ǿ)�0�ޡ��u���?�Y:q�׹>�L?]��?̒b��A��^�L��h��샽4�?s�k?1��>��?u�?�ζ��h�(���8�=_�p?0�?(!�?��>��=H�:v��>V�?6��?�R�?�Z?!mu�yj�>2��9��>X����<>IYս*�>`S#>�0?G?=�>�4=�	�C���.��n����w%���!>���>M��>X� >�l�<i䴽v����H>(�~>~��>�=�>��>8:�>I�����9�>P?N��\n(���?K}�=Ui�=tyҽ�ފ=R'��kӽ��=��Q>����;��2���<�<��>cϿ�f�?�4>U����"?������=(��=�L�>0\��݉�>>���>�?�L�>�C�=YG�>U�>e���2>����.���J���Q��=оlj>�5���h������ט}�Ұ���(�Yis��P���HF�,��#��?��2���Q�v��
�F��;�>mΘ>sA3?mO��t�����=��?
6w>��˾}���TX���Vܾ*ъ?hZ�?�*c>~�>��W?�?J�1��3��oZ�6�u�j(A�	e�q�`�]܍�������
������_?�x?�vA?#��<8z>��?�%��֏��#�>H/�p;�_�<=$�>I$��	a�/�Ӿڸþ�;�eF>�o?�#�?	Z?TcV��戽0>ˈ8?R�+?(�n?]�+?��9? ����?� >�?��?7�1?�!?��
?*+R>*A�=L!<� Z<cKw�["���ߥ�{����Ӽ�C=!�s=����a�<�n=V�p<v_�N�\���p<�ga���<)^'=ܑ=��=���>a(W?�>���>%�(?^븽#��i��a:?g�I=S
E��<����n�9 ��>�-Z?.�?GT?5�w>��>�� ��E>�hU>��>��#>�p�>h���}� =��@>R�e>C�G=;T��[������%k��[�=�@F>�
�>jU|>�ό��Y(>�2��"�x�}d>�P��฾��R�
~G���1�S�t��p�>;�K?�?��=#}������e���(?�c<?�L?��~?jҐ=@H۾~�9���J�* �'.�>�1�<���񄢿�Q����:��s+;wDu>Y���rH����a>�����޾X�n���I���羙=L=�i��U=�/�}]־��$]�=�x
>�n��"� �����Ѫ�NJ?j�h=ͼ����U�>����>�t�>Ǯ>c9���t�W�@����R��=2��>��:>����}ﾋoG����>ӕD?H1_?���?R ����p�JL@�
m��F}��T� �G�?���>M$	?��?>�	�=���k@�WYb��6G���>���>�E�Z�F��'��RV��!�Ƥ�>��?�!>�P?��Q?+�?_N^?��*?Ճ?��>�>���ܻ��I&?Q|�?<��=qӽ�T�q�8���E����>l)?�OB���>�t?I�?!�&?�Q?7�?�L>�� ��f@���>5]�>��W�<T��5`>I�J?�>��X?�ă?\�>>co5��좾W����l�=P
>�2?F=#?�?˂�>f�?C�M=���=��?�wS?`4S?+c?���==Y ?~c>��$?��Z��>��:>�:?t�f?ӭg?��>?O4>"i8=�IǼ9WѼG���F�=�N�<���M�O<��=É� `/�c����[`��9�=.y�=a/W�EВ=�������=;`�>C�s>\���1>��ľ�I��;�@>�����P���܊��p:�S�=o��>�?���>-F#�t��=��>L:�>��|3(?�?�?� ;��b��ھ<�K�c�>�B?���=��l�K�����u��;h=��m?��^?�W�s&��I�b?��]?�g��=�*�þc�b�1��'�O?R�
?	�G���>��~?`�q?l��>�e�>:n����Cb��j��ж=Mr�>HX�7�d��?�>O�7?�N�>��b>
%�=&u۾��w��q���?��?�?���?#+*>_�n�C4��Ծ�����g?���>FK����?��D౾�}���o4��y쾔��������9����^I�9�u���X���=Q�?�
|?��c?�E`?��� f���b���@�V�'��s����;��~9���F�T�t����ʌҾл���=f�a�[L����?��?�-��}�>dZ���(۾��ƾbvk>�񨾸6彰��=y���T�<���<a���嫾�?7�>&��>��7?�^��4B��@2�/,9��+��[$:>�Ş>)�>��>���l@I�2?�՛��.w��������>'&W?j\?��p?=x��O0�����F�9��p*;����\>�B>Y��>.@���L��	�
,�'�[�6O�����x����s;?�m�>�m>N��?��?r0���Ӿ��@��:4����=�4p>�<D?��8?IV>���$�����>��l?��>��>�����Z!�?�{���ʽ6%�>�ޭ>���>�o>Ϭ,�$\��j��e����9�;q�=��h?惄���`�D�>�R?��:�G<�{�>��v�Y�!�x��`�'���>0|?*��=��;>�ž�$�	�{�g7��
(*?0�?�L��GN%�zj�>{e#?���>�x�>ʎ�?g��>ދ���L��Ա?ʠZ?�K?/&A?�f�>��4=�ܾ��Ľ�< ��1=���>ջa>~L�=U�=�H�e]�Jz�)AI=���=-؀�*͠��46�O�ż%eC<,=3�8>�׿F�H�L[﾿���aؾ���z)��RcP�����!�'�+⾗/��e|���*��D-��Z��Ӈb��;¾�ɽ�N�?���?GȾ�������m�V�%Pվ���>�2���1��z����/�]���R��E����@��]f��䌿��n�2�'?�?��ںǿ5ס�Y�ݾ��?10 ?�z?ɖ�N#���8���#>�<���V>�׆���Ͽxӛ�B�^?���>���D��>^��>T>��p>����cO�����<��?f�-?ڰ�>�.s�6�ȿ&*��3��<̰�?��@�XA?�g(���N^=��>|�	?uA>0�0��K�M%��K=�>��?��?��J=?W����K'e?��<�9G���ǻ/��=~��=e�=�/�m1K>���>�f���A��sڽ3�6>�҅>�'�*W���\�^<�<�^>A;ӽ"���5Մ?,{\��f���/��T��U>��T?�*�>T:�=��,?Y7H�a}Ͽ�\��*a?�0�?���?%�(?9ۿ��ؚ>��ܾ��M?`D6?���>�d&��t����=t6��{���&V�}��=[��>c�>,������O��I��U��=x��-ѿ;�Y�ˈQ�\�>}��(���|�[Gʻ�&�>��ǌ�J/��-��>g��=�=�>�,�>��>V��>ɕ5?�R0?���>/��=?�l=_�q���̾�Ֆ�r(h�W�<CKM�C>])�Q��>�)��R!����x��!��H3��>]q�������6�t�B��Z4�f�?��>�}Yg��j=hz�J�e��:�![���dNo�{�V�֥?
/b?伆�O?c��`7��S�<��2<���?��<;�>2��Ƨ��h�>����T�=t��>{�<F�c#.���M��z0?�J?\%��ѐ��+>,e ��=�+?��?�\<�b�>(%?,*�˒佰�\>pq5>�X�>���>n
>�����Aڽr?�UT?Ec��؜����>J��z�&3_=~>��5���켂�[>ě�<wԌ���R��/��#�<�(W?���>��)���a�����A\==K�x?��?�.�>e{k?��B?�٤<h��9�S���4dw=��W?�)i?y�>����N	о����D�5?ߣe?��N>zbh�.���.�3U�i$?)�n?Y_?z���w}�`��8���n6?��v?s^�xs�����M�V�f=�>�[�>���>��9��k�>�>?�#��G�� ���zY4�%Þ?��@���?n�;<��U��=�;?l\�> �O��>ƾ�z������4�q=�"�>���ev����R,�f�8?ݠ�?���>������o $>-\��VU�?_�z?x!Ҿ��l��P'�X"]��a��x<��B9��o�G㊼���
�Y��_�h��P��4��
�i>܍@Z��	?�Ð�q&Ͽ#�Ͽ�Q���λ��Hɾ�?��>��L�m ӾMn�p��n?4���e��ʛ�#H�>��>�Д�<�����{�ul;���j�>�����>��S�� ��������4<��>X��>���>ZF��轾�Ù?S_���=ο���+����X?�f�?�m�?n?
9<�v��{���D,G?�s?8Z?�:%��,]�J8�$�j?�_��tU`���4�tHE��U>�"3?�B�>S�-���|=�>���>g>�#/�x�Ŀ�ٶ�>���Y��?��?�o���>r��?ts+?�i�8���[����*�+�+��<A?�2>���H�!�C0=�WҒ���
?U~0?{�d.�]�_?+�a�N�p���-���ƽ�ۡ>�0��e\�N�����Xe����@y����?N^�?i�?յ�� #�g6%?�>d����8Ǿ��<���>�(�>*N>fH_���u>����:�	i	>���?�~�?Qj?���� ����U>
�}?^$�>��?*p�=�b�>Gd�=���,�ek#>!�=��>�M�?}�M?QL�>�V�=��8�/�[F�tGR��$���C���>��a?��L?�Jb>����2�G!�1wͽ	c1�)C�@W@��,�ҟ߽�(5>��=>�>E�D�Ӿ��?Mp�9�ؿ j��!p'��54?/��>�?����t�����;_?Pz�>�6� ,���%���B�`��?�G�?>�?��׾�R̼�><�>�I�>C�Խ����\�����7>1�B?Z��D��u�o�y�>���?
�@�ծ?ji��	?���P��Sa~����7�e��=��7?�0��z>���>��=�nv�߻��U�s����>�B�?�{�?��> �l?��o�Q�B���1=8M�>ќk?�s?[So���o�B>��?#������L��f?
�
@u@a�^?+�Bҿ{6��׃�� �о�q��5�=Ȉ�>DkӽjZ�=[�=h�������"��i�>2��>'��>�G�>� �>��>8&��M������=<��;�M���� �N���Q
��WX��9�����c��C�O=��۞=ӊ�ڡ���썾��=?wQ?��R?��t?�y�>�	��"�2>�?�����<9,?�ګ=��>��6?�F?LD$?���=KJ����[�
�|�/��_������>OTI>Q��>��>6�>�p=~�+>W\,>w1�>� >8<�#ܼ��h=V�Q>J�>d��>J�>�qC>7�e>4��i��S�|��N�1ʡ�拢?��D��^\�X]����-��ؾz�	>�t?��m=~{��q�Կ�¢� �K?��t�����06:�d��=M�?v�T?���>c0޾-���~�L>-lU�(���7e>L�O�<��>��n�>n�?��f>#u>(�3��e8���P�l|��nj|>?46?�趾�F9���u���H��dݾJM>�ľ>gD�el�����J�ui��{=�x:?��?Y5��5䰾b�u�NB���KR>;\>/`=m�=�UM>�dc���ƽ�H��X.=���=Ѱ^>��?	3>��=K�>�����A4��x�>�/>�E>�F9?�g(?���*�t��,�������>��>�t�>i�=��:��c�=l�>zM>������O�J��X��Sn>�`Ӽ�|��t��W�E=����y�>a�X=���tA���(=�~?���(䈿��e���lD?S+?^ �=�F<��"�E ���H��G�?r�@m�?��	��V�@�?�@�?��K��=}�>	׫>�ξ�L��?��Ž6Ǣ�ɔ	�.)#�jS�?��?��/�Zʋ�=l��6>�^%?��Ӿ�e�>�w��Y��m��/�u���#=y��>#9H?�X��n�O��>��u
?�?�b�Ψ����ȿo|v�E��>=�?���?��m�NA��f@����>���?�fY?�hi>ge۾�YZ���>�@?�	R?
�>O:�y�'��?}޶?���?x�>dy�?Q��?���>�R���S��ɿH���)�='�O>�5n>���:�S�Ǡ��?y���<O���+��Þ='�w="��>R>�3f��1��= <=�Ͼg���J?֌>�R�>E]�>�j?tr"?^�>iS=��Ǻ���!���K?���?��z2n��P�<��=C�^�^&?zI4?�[[��Ͼyը>ͺ\?>?�[?d�>���'>��F迿~����<�K>y3�>�H�>\#���FK>��Ծ�4D��p�>�ϗ>@���??ھ�,��1k��#B�>�e!?u��>�Ӯ=� ?��#?��j>-)�>�aE�u9��s�E����>��>2H?`�~?	�?�Թ��Z3����硿b�[��8N>��x?�U?�ʕ>ێ������b[E��;I�7���ԛ�?�tg?�M�(?2�?l�??��A?-f>���ؾ����>�!?�j��A���%�����?�n?�Z�>�f���
ս(�̼߬�����^�?�1\?(?&?�L���`���þz"�<����+p�0�;�A�GI>ޣ>�(���T�=��>���=��m��6��yh<Pջ=�V�>R�=0�6��捽0=,?ƿG�~ۃ���=��r�?xD���>�IL>����^?kl=��{�����x��	U� �? ��?Zk�?c��@�h��$=?�?S	?m"�>�J���}޾6�྿Pw�~x��w�Z�>���>)�l���K���ڙ���F��_�Ž`bF��y�>�q�>�?�1	?�cX>�g�>:m3���5���7<ǾצN��B���U��"��V�4�̾�����ǻme��Ϛ���!;>#���G��>n�3?�ud>3�>S��>�J�=��>�I�=�#�>���>���=�s�=���>k��=�ʁ��KR?�����'����@���,2B?iqd?V4�>�
i���������?���?Us�?�;v>�~h�.+�)l?%?�>����p
?�z:=e�PF�<�Z��E��J'��F�r��>3׽�:��M��of��k
?G/?�_����̾7.׽;���p=�P�?�*)?zY+��Q�@>q��W�_(S�0v,��Vj�MQ��F�#�55r�C	��5���ׂ���)�D� =�)?⒉?�� ��������Si��-A�	L[>
��>��>Mֿ>aH>&<���1���\��'�D������>��x?�Z�>�F?��9?�)S?F�H?���>%a�>]㶾-��>�~�;���>o �>�@>?��'?F<(?�? �%?T�c>U[�I��#�Ͼ��	?PK?�z?Mr?��?�/Y�ǩ�}A�S@�<UGr��耽p:k=��5<�����FZ���=}A>[?7z��8�#����k>�7?��>���>��������<���>�
?�R�>� �mur��W�Q]�>���?�<U=��)>���=����V�ӺMK�=����{�=쥂�v2;��� <A��=��=3`|���y����:���;�ڮ<u�>6�?���>�C�>�@��,� �`���e�=�Y><S>�>�Eپ�}���$��s�g��]y>�w�?�z�?��f=��=��=}���U�����E������<�??J#?)XT?^��?y�=?]j#?е>+�jM���^�������?%�?F��>�u
�� �>�����v��-�>�WI?�\w�����O?�q��=?p��r!>� �SPx�VJǿ�)a�:�u> ���-Ƚ�r�?1	�?J�D>�9c��/��3h�+�p	%?'|9?�`7>߶>�]�/#�N���OZ���?�0^?�9�>rN?Wf�?�Y?h�>��,�$��^替~�=��>�7?���?�s�?Ӻu?�\�>c�O=�{0���־a*���h�Z@�%�����=_��>1\j>**?��>��?=]�����˼��L�`�G>��~>;��>���>n��>)�>.�;��G?E��>�R��2q��Ǥ�ۆ���;�ru?���?ޔ+?dx=r���E��E��m�>�e�?<��?�**?FT�H��==fռO׶�
r��*�>D�>g0�>a��=TF=Q�>5��>1o�>Q���C��k8�SM�B�?�F?��=�;ƿ7�v��|�㠾
�<���$f�����Q�<��=�Ѥ�c�5�}ͭ���:�1��}����׫�-���Wr��/�>�[=���=e�=�	=����	�;9=�'~<l=Ut���0�<jm"���:, ��n���v�;��R=�%<�ʾgC}?��H?a�+?BgC?+�y>+j>��1�!F�>���e�?��V>�I�������9��n���˔�o�׾Qyؾt�b�9���>��K�'�>4>1 �=�߉<� �=��u=�=)+k��]=	��=E0�=�{�=�.�=��>Fd>�6w?X�������4Q��Z罥�:?�8�>e{�=��ƾq@?�>>�2������yb��-?���?�T�?>�?@ti��d�>M���㎽�q�=K����=2>r��=w�2�T��>��J>���K��C����4�?��@��??�ዿТϿ6a/>?:>a#>1�P�R�-�{Z��N]��O�I� ?�<��+;"�>�c�=�۾=�ƾ6A=�I;>NQa=�a��]�*�=�p|��9-=Y�]=os�>#=G>��=.Y��&[�=]�X=���=L>	�nVB�ë'�6�4=�t�=C�e>��">��>�?��,?�Jk? �>��S�ꀡ��7���i>��J=�.�>��=��q>V��> e3?�C?&�>?��>+����t�>�j�>�0/�^cd�]u�-���Փ=~:�?�r?���>�e�=�(�{"��J;�����B
?,4?M�
?�o>U���c�(�I�0��z���ٕ�8�=��x��HE��*��5�*���Q�=���>�+�>Yȣ>3��>��?>�NK>	��>��=��<va=�<ʉ�<����|=z삼o�2=B编,<lQ;�^�
�E���Y/��&U<:�<���=��>Q<>ܬ�>h��=����C/>���2�L����=GG��4,B��4d��I~�/��V6���B>�:X>�{��(4��\�?F�Y>Qn?>���?�Au?i�>]!��վ�Q��De�8WS��θ=�>��<��z;�-Z`��M��|Ҿ��>+z�>�6�>�$A>��c�a���<&1C���W�`H>��轣��<���������⍿Fϔ�"������"|`?1I��z�KcO?��y?q�?[�%?�J������>U�ro�=�:��<M�<�B?��!?o?i~���_M��K̾	���Է>)I���O�!����0�6W��۷�x�>媾f�о'#3�mk�������B��rr�2�>[�O?�?]b��W��SHO�������?p?�mg?a �>N?(5?�W��|X��h���L�=��n?a��?l;�?��
>'>�|%��A�>^#?�b�?ɷ�?�s?O�8����>ã�=�=�>&c��v>$h)>��J=U$>��?�K?��>�Eý[��������`���c���=2��>(.�>G�R>���=$y>OQ�<�*�=��>*E�>2�@>8��>X��>̕��+�)�A�>]a�=ڠ>(�J?�6>��>>.�;�O9��Np���4�Yc��)`\���Y���P#����=���1�>P������?,�ļB
�g��>w�ܾ]x��姛>@�>h����M�>��`>�g�>��>��>�>�>�^�>�O�=IӾ�{>���xh!�{-C�;�R�%�Ѿ�~z>6����&�ܢ�pv�� KI��d���f��	j�z-���==��<�G�?l�����k��)�Y����?�Z�>j6?܌�?��q�>��>c��>�D��f���wǍ�Bm�t�?H��?�;c>��>A�W?%�?֒1�3��uZ�'�u�g(A�%e�C�`��፿�����
�>��&�_?�x?0yA?eQ�<-:z>M��?��%�\ӏ��)�>�/�$';�"?<=�+�>�)��\�`���Ӿ��þ�7��HF>�o?<%�?jY?ETV��ѻ��B>vO2?ov8?��j?�K0?�A?'$��5?�>?�?��? z9?	_!?Ur?T�W>^�>�$=٨4���Z� ��� � �=�􋮼_ؖ=v�=���<�2����\=�t=h��mMM��d���r����<�0�=��=4�=K�>4]?���>���>=�7?I�.5�V<L/?3�W=F�}�������^%�
�>G~j?m��?�OY?��]>��?���>��<>.K�>��*>u�^>���>Pm���F��'�=�>w�>���=�)1�X1���#	��d��IO�<C!>��>�0|>���t�'>_|��a0z���d>r�Q�x̺���S�W�G���1�k�v�wY�>/�K?��?읙= _龬-��JIf�!0)?�]<?�NM?��?9�=Z�۾��9���J�>���>uU�<��������#����:�'|�:��s>2��
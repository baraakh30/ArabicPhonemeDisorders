�   �   �=�>�� ����;��U�]�(���'5<z��>ؽҼ2���vj=��G>���=ф$=�d�=�eн��>^q�=��<|�>�r�<� N�$�=� U>b�e�b�h����<s�þM�V�6�h>6�5>p��<6Z���༐~C>wE+>q���v��#2�=s"?Q�?�!?��">�ؾ6�����2�ʁ:�n*>�-q��Ǫ�m*������~�h�����5�W�>1����>��[>T���q��=N�=w��Zp�IP=�NI>��:8{�JN4>	>w=�u�=�ǿ=iv?��ϙ���ۿ����}���Ӿ\�$�
�Ǿi���Egl=�^=&72��o=.���]ʽ/�=�$>�3ӽ����h->��¾+���ܾ!��6��[�ھ"�վ�\a>�LL�������2�@��/��h?B��Z��9�����(������x>,��>9u�>�9�=V�>d?�F�>7n�Ei�>�"?�(ӽ42-�ϳ�=�7=d`=Um">22`=b�R=�5=S�y��IF�Epv>�3�=����m�)><z>��4�QM�>5U=�=ɽ��a���O#c< N�=�Y/�Rƽ/v(>*�3>~��>ֈо���ֻ���
�N��=Z>g>�/�>�dw=z~�h|��6�>��<&;=�>>�j>O�%�t =�3�;�{>S�="�&>��ս6��!!��CE[>�p!��Y����꼣�ؽ�@<��=M��=�����S��Խ��>p\
�B%�O�J?H��>�l?���>�U������e���V־A	=��>�˾I$
����}�������y�®���n���پ6+=���=�Ut>0�=����m߭�p�>QZ=Z���uL;>�Ϟ<uUƼ8��<�]�=�`=��#��W�5m�������������ھ��2��x=�7��%*H=�j>J ;=X�>3ϟ=�!�����:ư���=wy>�����Ƚ�#�>�%ݼr�}�5�x��~a��p��f�>>���F�s�սx�<	m���V�������;`�E�����[�A���>��>v�>;�>T*�>�Ȯ>���=GA��=���>�Ⱦ>�D���=�IN>�&�=�H����<w�<��G>w��<hn��t��_=w�>d�>���׌����t=�r&>)�=�/�D3<�Li罿.t=���="4�="�齢�E>|W�>y6��4LM�v򁾰���>�=S>��=v'T>�ǽ"��~R	=v�I=V��>�P>��>��=��=g�:=�Q�>�j�=�E��r(=%�\���
>@�=�=>��p�AH=+���*=K$�=����Ω>���H`����=j=�mE=X/7?<z�>�6G?.�<���.�QD��8���\M=ar>�AT���< ��� @���c����v������`������=X�=%1�=�����5J<C�ŽӮk���>�cP�E�>q�,=�$=�V�=��r=�!O>-�,�Zo{���Ͻ��տ�����V�=M[���0> ��u/ξq�"�8��=9U��=���9��jӾ�7�e�ؾe�:�M��k	r�t�>��ξ6�T$��.���S��!���{�o�?����Ǻ�N� ��k��wUe�n$�<�4��������v=O����A�>Ԡ+>�T�>hK�>5�M>��?���>c�>���<V>>�]0>�">G+>s��=~��=��ƽ��,>%�>Ⱦ��W��fYu���J=���=y%�=뮲<$�F=ןG�2ν��=+�0=c�� ҕ<d�=9н|�ɽ�V�=a��/#=�=�>�� ����;��U�]�(���'5<z��>ؽҼ2���vj=��G>���=ф$=�d�=�eн��>^q�=��<|�>�r�<� N�$�=� U>b�e�b�h����<s�þM�V�6�h>6�5>p��<6Z���༐~C>wE+>q���v��#2�=s"?Q�?�!?��">�ؾ6�����2�ʁ:�n*>�-q��Ǫ�m*������~�h�����5�W�>1����>��[>T���q��=N�=w��Zp�IP=�NI>��:8{�JN4>	>w=�u�=�ǿ=iv?��ϙ���ۿ����}���Ӿ\�$�
�Ǿi���Egl=�^=&72��o=.���]ʽ/�=�$>�3ӽ����h->��¾+���ܾ!��6��[�ھ"�վ�\a>�LL�������2�@��/��h?B��Z��9�����(������x>,��>9u�>�9�=V�>d?�F�>7n�Ei�>�"?�(ӽ42-�ϳ�=�7=d`=Um">22`=b�R=�5=S�y��IF�Epv>�3�=����m�)><z>��4�QM�>5U=�=ɽ��a���O#c< N�=�Y/�Rƽ/v(>*�3>�=�>�� ����;��U�]�(���'5<z��>ؽҼ2���vj=��G>���=ф$=�d�=�eн��>^q�=��<|�>�r�<� N�$�=� U>b�e�b�h����<s�þM�V�6�h>6�5>p��<6Z���༐~C>wE+>q���v��#2�=s"?Q�?�!?��">�ؾ6�����2�ʁ:�n*>�-q��Ǫ�m*������~�h�����5�W�>1����>��[>T���q��=N�=w��Zp�IP=�NI>��:8{�JN4>	>w=�u�=�ǿ=iv?��ϙ���ۿ����}���Ӿ\�$�
�Ǿi���Egl=�^=&72��o=.���]ʽ/�=�$>�3ӽ����h->��¾+���ܾ!��6��[�ھ"�վ�\a>�LL�������2�@��/��h?B��Z��9�����(������x>,��>9u�>�9�=V�>d?�F�>7n�Ei�>�"?�(ӽ42-�ϳ�=�7=d`=Um">22`=b�R=�5=S�y��IF�Epv>�3�=����m�)><z>��4�QM�>5U=�=ɽ��a���O#c< N�=�Y/�Rƽ/v(>*�3>��?�>���/�%Q�3���ؽ��>�])?�'��=Qq���Q�>����Ⱦ_���̾Z� �DH�>c�G>y�w>�>�7����<a�q=:~><E�=n�.���<�> >��=���A�y>S��S���������_���!>���>hj>¹-?1.?G��>@�u���þvXM�eY=�:�XH>�,6�}�6<Ht�#�`����eW���Ծ]� ���q�
@7=k�U>*z=��=�๽�������=&K&=V�M<-#�=�:�=K�=<�>�Q�>�,u>��I>�8u��ڌ��Kۿ���+�U�M����=�a���44�dq�=��ԎP���g�I�����ɓo>���>
e�>�(�>ϭ	>�E����f�ʑӽ(_�=�Kp����D����ϳ�t�=햧�@2ļyP����= ���(2��B����� �`�ξ��L���d��>M�>�NB>u?���>,�>P��>�j���zA?}���7?��ƾ���>j<�>!O�>��#?�-?�O�����=nu�m��tjW>0C�=jyV>�z>m�O>C�H=3>�'��`=�[�wT���mȽ�T��c�;!!>Q�>���=pJ?`���{�k�W�$>¾���� �>� <?�xپ4�q�࢔����>�	ž����оOl��/*g��)?R4>tN�>LM�>@����B��W�� {>�j=Iu���#�?���T4>
lнF�R=�C�1.��z-���S@=�>[jC>	�n>��?��.?{F�>*|L����F��	(�Y�ƾ$�=M����c��AH+�+(��7p��
>3�~���	� Wh���=��4>@7�=_�"��/���=���%���_>��c>��4��t�W>��V>ց�>x��>5�e>�.<=�+&��>F��0ȿÞ���"�!�y��Pa�ڕ�<6	<找� �=E| =�~B��ż�#�=d��>u��>5ѭ>��$>�ý�~�=�Ѥ��W��X���[�A����q��<��z,��%a��Pӽ��P��1�<�0�}$��y�R˽E�C�Z�k��Y_�l��>R��>���>(Z?��??ռ>��>�=��+?a �=�.�>YK����>O��>^&�>/��>`�?	$�����%�ݽ�v�]�>꣄>-�s>�c>$F�>*Y�:�=�;q>�z=���y8�� �<��e�2^���'0=F�<�>��>��o=�@o[��^�����r��=>I?I�"�K�|<,h���<�>�//�0�H��p���)>���>�i>?"�!��>�Yy>0�*��L�=w�A���_>N�&��H<�2r��U�=c�">.nj�I`i=;󆾚�����=;�5>���=`�`=�g�=o�T?��6?���>�+[��#�duI��]��Z��kP����H������%>���x���'���%�=6"��2>�}�<�Jm>�=Ձt�&�<)#��K*.�	%Z=�ӥ�%��ϖ!>�gm>I��>j�O>*��>]�>2�<�p˽)\=��u��%����;A����=F���U#�={LF>���eSm���\�z��=蓈�#v>)��=�żC.��a�=��[�?6ھȧ��T�#�L�k�v1��V �������=ǖ3�)f��q������Ǿ?$/���e椾�����&��F���j>�>�{~>dN�>u�?��6?�J�>�R��I,?>�J�>p=�I;?.?�??�%�>��>>,
��G>�:J���T�_	>;��=�H>>{��=��[>��<�ZS>g{��k=�#��5���R>҈=E��<-�
=�L�=%T>F��>)�̾ɱ�Ț0�\�վ����P�>���>�]#���>}G�=8�A?��`ľ!g�����>���>k�?W��H��>H�>Yد�\t��g���3>�8>�M��AT�M�p>,k�=��n�Q?ν��:�OU���~=F7S>	��=�!=�*>Q�>,1C?�I*?�Y
�A0�����&K��E���~�=�M������d�;Cm��U�N��B�U����ѾRi(>�)�<�z>e:�<s��=�i��j�ʼ��W���r=׷)>83��|�=O�>vŌ>���>�`�>+��=�y�Tw�)��H���F݉�n���2���q>&��Wℾ\>�a�=E��B�C��>J�+�4�?>�J�=c�R>ܯ;��Hb���Ǿ�½�����|�<�׏�Z�[�����L��m�<��7A�� շ��y�=�q"�����׌%�Q���Y��B@�Z`;�u�>)-?�=���>}f�>��?q?ƕ�34?�e��7d�>#�=�?g�%?�&�>�>��>�<6�h�2>.�9���\�aM�>$�#>��>��=���>���:��*>���;��=�ޠ�����ƍ�=�7���훽 3-=֏G=Z�=>�?�ʖ��wI��@����>�����)�bZM?���5�:?�� ��e���T�N�$���I >Qn�>�E?����c>4�T>��<���=x�όl=`�N=Oz9<�y;����׽⸽�়�i,��\׽�jN=<�L=K�r=� �Lم>�K?"?'K�>�������2��=������ ��CG��)>��>܍������0�]�4�[?��B���=9��;>���<���Cy�>[���I6<��M˧>���ͩ}>��M>�.t>�!�>�K>�C�=�>��(n��&J�����*���毾�KϾD�B��;�NS��{,j�u���9�#}�����<�>��>&�>�t>H�B>���>-�|��ν�&Q��xw���u��������Ub�=g����0Խ�*�����<�cV�����j�9�F��k=���\.�"em>D>ǒ�><?׻�=�]E?O�@?/���rH?�2���)?O��=Z�?��P?4-?2�H>Պ<�k�QG>9��OA�������=������=Gb@>u��;n���i
>ef�<LlϽ�n���
=��=�3��ʵ.=�@ >N�(>���>2uC>���8������/V��"�����>H�p=Fr��0�Ⱦ�/��P������߾|�q���ؾJdg��'���>Y�,>��
���4x�r�<��~�>�)�=B��*h�7��=F줽/}ӽ�}==Ã=�>A<��h<�ǎ=ЈW>�`�>+?��,?�
�>��4>o�þE�ϾkL�f:�=���>��>�9?�O1?�.=ɓ������p���M-�C�
�5�<�2�>x��<<�$�x>���=�3����=�t~>Ɓg=P]��b���^>��P>���;��9>���=i^3�%���*J��Ä��q!4�5��T��p�\;!����H���0�;g+�[
��im�>K=?n�?oN@>]C�>�3?L�����5ɽ��;5����n��4Lu���ϼ��4N��g'��/<f蔽�!;��C��hT�Z/������(�J��>j��>�
?�k�>�[�>KM?D�&?7Q=�]>yr�>Da>����S���t��|�>B>"��>�1�>5e\>�g��S�rq�={R>��$>,钼��4�|�.����M�=��n<���=ˑ=X5-�I��;��=�F�=}��=mf�>�~�=����$A*���؛�꥾�P�>jn�=� ��U/�7��@'�/{��,4�����Ƶ�ȫ��6�%��>��,>v�<*0�<�ȍ���S=}2>��s����E9�2V�=�0-������A=g!���������=�����m�>�w?5XM?a,?������t�j�L�����޼8��>�\>��?h\>>��@��� �����;�������(D�=Y*>�{�<Tc4>�|�>>�S��f=�2S��a��9>��>��>_�>��="�J>�x>�)+�y�Z=Ѝп�����O��Y*�$��-ж=�.���޿>Q�
�m�L=�b���Ľ2S�P>�~�>�Q�>B�>>��>�R�>�ј��z�0��7�,�=a�AN��؇�̆=�C#�ḗ�ԝ�]`���D�%.� �j�lw�:��I����H�l�?1�>f��>ѥ�>h`M?O�??�0���a>��C>H�>;y[>��A>000=��>�\>_�?�|?�
�>J훽� o�MP���O�=K">��8�_h�=�F��b�=�6�>@��m�b���м��>ޖ�&>��>��>�'O>)�?<f0�)d,�vd7�����Xܻ
�#?w( >�;���z�,C��i!�1M���M>�1��A�6�:�پ��྆�7>��<A$=�� >�F]�&7�=Rb+=� �旅��&<(��=�|�<csL��=�d�=�Mi;�޽��'�q��=��>'�>��Z?x,?�睼~N�+L�#�"��m#�"��=��J>��>�o?�[>Wj�������~���;%�k���>�����<��=���� �=��o=4~2>'�!����p���.�=�n~>��}>�->(��=F�����Dο��P4��6?����=�W����4�k��=��x�톮�U��&�f��%��f�O˧��)ѻ��=��o>9�:>���=�1���=��	����a;��|`�@9�<�⺼����c��7pɽ@ҽ~I��?j�df���"���G�Jy�pD ? ?���>��?���>�G?L�?�	�$9�>b�>�R�>8���_�>�!i=K�>�?l ?JX�>���>�99���*�"��@D��[D=w�=��<i�;?{=v��=��E>^}�=���<�ˤ��cN���=�sy=�J!>�_>�t�=�M_=_[5��wC���Q�f���~�;17?f��>�'�(��1za��&���F�=o���(�WJ/�EN�J䖾r�`>��$�
>'؇>~^ݽ
O�0�>L�$p8�L�u�׀S>�;��+����=��=���|�xp>t�~>z�F>�?��D?*$?�M�=k�վ��*���@�~�o��=�p�>8�p>��=�� ��_u��4�2Xƾ��'��ڬ�݊)= 'L>��\<>+{=�^ >�b�*T��`�,>kp�=s�=`N��>�����>�Ha>a��>��M>6�z=��Z�,A���~��|����Ǔ�F��g�l����j�����c�ap��S9<��R>h����,׾�%�<I�5>���>Pg���dn�m ��x� ���C�����½�aR���n���Ͻ�{��Ƚ,-q=gѽ�n�����0���g���7L���o��?��>ޥ�>:��>BJ?�0&?�W?bp��]օ>�?W��>�KԼs�	>9͂�o�?�_2?��?��>ߗ?��M�,s��
ϼ%��;Va�=O�>��;1��<,=\�݈Ž,��<:��=k製m �}&r=S��=�r>P�>��=�Z��M�6�>�W���پ���t����W7?u�>�Y��J���޾���O���������<���(d!�`C���>�66>��=v��=��½yi��dx�>N�U��-���ཽ%="��=`jW>0ż=�yt������U��8N�A��D�>>*�7?��m?3�2?b��=�w����9<Y��8(����=Z��>�
?�?+7Y>GB���/� �;P-�ƿ��k@�����>�N;>�&=�,S>r��=��"�o���5Q^���=�a<<�d,=��]>Rc>�W>��>���=��۽�w��� ÿ4���KϾ��������/���d�m���'�����=����B|���p��'Ҿ����`�
�7=�^R����=<�оaW��t�C�b��#���;�Jw���S��� w�R�I���n�f�D�(S��Jk$��X�#D)�튧��;8��eu�N~?e��>h�}>�:�>5��>~�?~�?���=�6<>�3N>�[�>Ih!>r�5>�>���>��>n_?T{�> �>�6�=�u>� ��6��<�B~<�F�<ږ�=c9�=KA6>H�b=+��=���<���w�ֽ�t�=e��=��*>bo7>? `>�6�>)郾�/�5� ��Y�n>3�r>F>��>��9�<�?��Xf���{��*m3��5�D ���>��>�ݎ>�С>ц>huL=��>u됽
k=D׼�>ƽa�	>p�w>��!>���e۽�닽�����2�p�=ߛ'>g3�=O��>�kl?�W+?�a?YY#���]{�x�l����>��>CB>`�>�O�=���X ��S����	8���ü��R=��)�Sē>K=�>Fp<=+P��f��y���w�� ����=d.>!�>��>�T8>.��y6����Ǿ
��B��+�����~�
=S:μ��"����bD½Z q������*>�ҁ<���>��I>�D�<��=�b<��>R����9v�q���vd�� �=��\/�>s`�q��켛�XR�� }���N���:�M\�elA�R���)޽.L�=��+>�z�>��>�gn?8��>�`�>w���0?�t�+��>���=h�`>U�>y?�?�M>]4<A��2��K��oD>L�N�b�=ޱ�=��9>>S��=
>QS�=2�ѻH���V��=r���H�`�M�<VL�=�">��U>�o?w�r���;o�F�<��	�����>����=x���_J�x��=�I(��&�e$��� �F���3e>he�=��>t :>0����h=R����:�=sZF>�L=S=�=�=��ER=�kݼ�
���>v�=��]<@���5=�2y=3<��>� ?f"w>�-?�������V�;�6�p�v�����>1B�>��ҽMa�cd�����#]����[�����=��B��z�<m�M>g���׏>@��=�֘�*>>��)�(v�<\B�=���=q�>�_>JA�>��> L�a޽��Q�R'ͿeT���͚����O�;��$�̍�%K�=���[yp>�Z��{&P�?(\���2><^�= ��=���=��n�ɜ����>�N>�>�vU�;	Ǿ������&�;>�@Z��1G>Ќ��~W���@v�T�q�M�t�Mg:����;A��=����5x�>��$?��>ke?�� ?`V?��qs4?r���CX�<s��=l�?c�@?w?��?�?��=�O�t�_�� ��WM�=1�=�Sr=1�=�l�<�6��jS�<ܤ�K��<
x�=jה�9}=�Wν��=i��="v:=C�=K�3?2q�H^�������B�#�=��=��>P����Ǿ���62��j� ��D�#%3�H�*>���>��+?�SQ>mi�>�$>�ظ�>L~ �!/Z���>=�aA=2#=Ċ�=�]> �<f��<6j= S���pC�����������R=�.�>&"g?N��> �?\���0b���"��1�����>�y�=�Uw>8��>���m%�<��w�,+R�\�O���̾���h-^>:Np�%��<)��>��>�u	��o���5ؽ�1�ws����x>̟�>�h�>��>�CE=^}��˾Ϳ਩�[�Ͼ_Z.��܋��h�1h�֢�>�t>���=;־��)�/t�.Y�<U-9>��n>��=ٛ��yһ��v<����i���K����`}�jQ����=�C���V���b����<{O�ѺX�Hx��#�н5M�[Eq���.�µ����>�5?�?�_]?�'?ȯ,?��t�h�*?�〦>�e=h��>��??��>cџ>^q=��\�4x�=��L�D�j��H�>]����<�=�.{>���%>hS�=Gy;�kM��`�<!�ν�6=�zn=�#>
M�=�qh>��?�4�=͹����[�縝���)�$?z�ӯ=v<����ܫ@����[b����g��}�ѽ70L=��>zhd>&��� �9��:<��=�ϥ��b��<>�v�=Hq�=�f�<x���q(��C�:��B�Rd=���<���>)�a?�?`�>���xG0�He����M}�V�>�{�>�θ=� �=M�Xn�+fD�v�7�J��Udc<���ɷ<>���=z�>�\>X��=<�ڽ3�����9�%���z���ڽ
�(>��>��>bZ>�{��Y�
�M~ܾw�� ���X���K�o�%�F�Q�3��X{^��*>�2��jL��I�>#��>��F>`��>hő=_�L>n�>�;�>v�m�;���C?u�-���1�鮾iI>��\�,���e/��#~�ۗ���c��'�1�d	*��3��D<�#d����
>
�5>�!�>�Q,?ΥD?�v.?�N?k6��Tg>�+���b�>��>�E�c?~p?�e?�-?�>Z5p�r��^�G��5>�=c=�"�����=�"�<�5>ޛ�:���=JZ=ق=/]�<'u�=O�ɼ�u>��=��7>?���O	��*̾�.�^�m��=<�?Q�ﾽ\>�q�y�/�<��j#�e�xh>y��>(��>-�=��>f*�=�
��֟=G3��BEg=���,�o���=��<��=��F���P`����l�ȋ
�����(�<�1>ʔ>v[N?��>û?�������:�2�G���tm�B�x>��9=1�>Aͣ=�^;N�a�2C��U1�f��,Zo���Y���*>J�=����L�/>y2�<�{6=.d�=pɠ�HM��*
d��}6�U�>W��>K'�>��>���=��^K��D*��9���w��HbN�d��f��K����e�a���v=��½���=���=�!#>�bv>jz�=$>7�ƽ�2=G��>BD�=v���������R����ؾ��I>�!龻����h*��H�%���扽L4@�
q0��Q�;1���W[�F��>3��>\��>��_?�}?c�?T�����C?�08��2a=<�6��?b*.?�?I��>0�=Uᴻp��B9��������]>Ʀ*���=���=�>?ý<[�=sj{=��[=��=e>?<뫴�v�a�'q4=�+)>5�>*�,>�[�>H����W�y�G��^v>�S�>Xn?�,=�t[���B�m-����L��N8>�>�*>{�����<	t�>��=�$�;D���D��o�=N
>�?���f߽k�X>��}>2�1=���=u��{�=����N��<��=k���jl���k>��>x>_?��O?�h5�}���*K�p G�13<��&�;�*�>O7?/�>���;��*��!�����}n �?,����=�]�=K =���=ƪ�=��#=~�>D>��K��[/>L'3=>�C>1�>O�8>�(��"	u�����BԻvPԿ�%=�{��;�,�����B�Ⱦ(�;��)�T}��7�Ѽ���=f������)(��$+�E<N�3A>P��<W�<�~?�-ýr2�}�=xZ̾�����=�%�K����[�*�5��dR��v_����ҽ�`J�M�����B��^=��k>*d�>�Ty�,s�=J*?��>��>��>�<�>��m>�w4�9��:L�}��ӽ*ؼ��x'=���>��c<b�s=���n�o�Z��;& =.->̀��(kJ=J[�<�p)=��&�R���� ƽv����d�<|=��=
�ϼ��_=�)�>�߾��!�EN��� ��}>3�=i��>���T�S�̾.� �|7�>`��>����������9o>x�ɽ�@
>����A���a<�>5��>�pQ>u˽�=�=�P;>ሪ=T�Ͻa��B�8�I'��'�<N�=�f�=��<?]}>�N!>�a?�S=?�3��h�+�Bn��M��K<�Y�> H?��,?��H>�W���ɾ��L>Z�r'V�w�B�v�[���=f<>��i�J�o�*Hs�c꘾���=U�&>*@v�$8>a=Y>�q<�@l>�>����ݚ��8-��_ֽa5�}���া��L���ܾ&x��P�^6��c/�2���[�T�?~�>k�]w>�E�=�̙>`v�=y'��(�O?���=�/���R�;���ֻ��8}�i���Ѿ��t��#w����<����c���n=�я=j�ؽ;_�� {� �L>�"?it�=#�|>�;?O�>W?�nb>d�> �>�&���Fd���������ψ>��׻G��=�F�>�y>g�Ҿ��a���<�J-<�*�=_1=���=�ͦ=iV���=�%u��e�eP=ù ���o�T�<I��bǭ<�?�㯾�0�R��N��g>�>k��>?@��N>�!Ӽ�|��=�
�(ѧ�h8<�ʭ>��>�"�><ߎ�V��=1�=ܥw��Em��[���Hӻd:&=Al�;Sw�>�5�=~"��nm>9y"���7��	�.,Z���߽dOL=���<贤>��>�)R?[<?��ǽO��ٷ)�Ny5�Eی���n�Ի=����=Ac�>�L�>�n�%����,��ȗ���>�L�� �Z>6�=�'�>�Å>F���J��;�<��,�襫�4�=.�7+�>䎵>9a�>��>���;�_��j3���пI2g���?��Ac��;G^�����հj���Q�����Q�9a�g����f=Ԩ�lㇾ%L� �=Cͽ��?{���7@��O=�ʣ��c�� �oga������c>��ܽQ�@�G���,6Ƚ-~��g8=��'=Wq����?>��?�=���=Ct?���>�߸>CK>>�>dd>_��>ny�>m�j>cS==���<x'�=i>��*G�=�I��şR�C}><H?�(X�;��=p��=�t<�T
�jn7��>�c������켼oǼr�-�ql2=� >���=D��>����E~����-�>*�A>��/>���>a��=��t>�'1�Ȑ����"��W�<�d�=e�ʼ�����>�k>�!>~��<�X)<���9�+��<��m=�Sn=��e>��>�.P<bO$>1Τ>�/ٽm���[�a=w�=�6<�\�=�co=u;?��A?��C?��<���þ100��k�ڭ���fA=�}>f��>�~�D�ξ��վ�����*��%l��垾V����>zl�=��1=|�3>�Z�<S�=��;��r="fU�v7=�z;���N�5>��R>��1>����`�@L��]�̿yM��L��2"�f$��@&�3K��a��c��{��W�-��9�=����=������>�د>R7Q�cvT�r�=gm��������g��4���H�bo��
=��u��V�[s߾g	 ���#��5�=�8C>�?�=�_X���>'@�b �>@��=j��=��`>z�[>��?1>�>��
>�>�>*Y����<����O�+>t��>Qk�>�p�=!#�=O��=�|�=�ǽ7�u�_x�=��X>���=�T/=5����ǽv�!�s�q�)�t>��ν��^�4��΂��Ơ|>C�>�!�>G'V>�#?T2Ѿ��������x��a۔��8�>�{���ľ39��%�ܽ����>ZY~=B���>EV庹�>���>r��<5�v����" ���>U��;�@)>�<ʧ�	B��o��=j�0>;�
�A�ӽ������ս��S>k��^9�>ꝷ>�<C?y�"?�����$�0�v�4��þ��+��nU?K�)?�' ?`ľ�@j/�n���r���A��a����>�>0W">AM��k��F=�ą�1�h�|m޽M-�>�6�=Ѧ|=ضe>���=���<�o���]н�W �|/�Zz��/Qľ>��W����6����Ҹ��ײ����=���i5=q1F��:��,��N>�jh>�@��h�;c�>�i�����>��+ɾg闾�e��'����O��jm}����z�v����<�T��d�Y���_��8K�<r�?��<�~�>�u�>�?w��>ᾴ>$��>z>�>��뽪?��%�6���ڽsˍ>b�>sq�r-�>�x�>�sB��=!�,>�j�>
�4>�Q�<P��<1U^��8M>b�>��;�t��u��B�<�֦<��=0O�=��ý�b�=!{�>/e>v94�iM�F�ƇܽS��>
z�>��A��	*����$�)���#A�� ��1>L&�>��>Z�=�͠>l+>�]��SH��X��L'>�	<>B�j����>y
����� *=T=�7A�n�3��=�b�=�x=T`�>= '?q�A?��)?���7��m����	��3���sܾ�`�]�>�������37ݾOg@��)��$�N�=�7!�.�=��<>ba<�
>i���/K�[�>zѱ>�@ϼ�S>H�L=��=��D=���>4^>����Q���Y��<Ǿ�l}��㾴����$s�Kܯ�X->Ә_=�)�=X�ټ�����t�=v�>��?�5z>/-�=�b(=H.��FC��LN=�M����YF���"��U�B����=�냾ϛȻT4��Ҫ�-�Y���̾/Zs�T�X���a��� ��,: S�>�F3=���>�E>�W?�?6?Q�:>g�
<˓B?t�>� >7?�.?��?�>?൲>��U>��>|�S���|������_��=��=(ה=�=lL�2�j��`�w��<�|>^c��XAE>�$�=�7P=��(>�S=��=��>�=�B1��� �9*�� D�oA�=�h,?��2��.�=��=d���I������ ��= u>��>N"?��>`�>c��=��B�� >�rt�=���>[��:�k�=�L�=C_W�40�=��m>�&ռ�=I���u��t*>��>5_^>���=��$>�G?�|F? �n?�3ʽ62�L��c|/�*�0�����ɖ>��>}H0�뿶�%w0��^?��[��%���6���X�'�?>��f=1F?>=��7T�M/>.!A>sG�=\��=�>��b�>��F>���=�/�=�0��_p;ۯ����/���\���쾊��=C.=���<�ȏ�)�:�����NG>��%�=ؒ�=�	�>��>O�z=�KO���徃re� �/�-��-fO����`Y��%�����D�Z���@;1�~�߁����&���%��E9ƾ�6־<�ɾ4�*��~�>$/�>���=��L���??�+3?*��>͋4���?|�^�����.>h��>A� ?�C/>�e�=��]>>M>l��>ߝT�&ј�D�s>��9>��>�C>�u=K])�J�7=��>^l����<Չ�=���>02U>
;ئe�m�=<Ů=!{�>/e>v94�iM�F�ƇܽS��>
z�>��A��	*����$�)���#A�� ��1>L&�>��>Z�=�͠>l+>�]��SH��X��L'>�	<>B�j����>y
����� *=T=�7A�n�3��=�b�=�x=T`�>= '?q�A?��)?���7��m����	��3���sܾ�`�]�>�������37ݾOg@��)��$�N�=�7!�.�=��<>ba<�
>i���/K�[�>zѱ>�@ϼ�S>H�L=��=��D=���>4^>����Q���Y��<Ǿ�l}��㾴����$s�Kܯ�X->Ә_=�)�=X�ټ�����t�=v�>��?�5z>/-�=�b(=H.��FC��LN=�M����YF���"��U�B����=�냾ϛȻT4��Ҫ�-�Y���̾/Zs�T�X���a��� ��,: S�>�F3=���>�E>�W?�?6?Q�:>g�
<˓B?t�>� >7?�.?��?�>?൲>��U>��>|�S���|������_��=��=(ה=�=lL�2�j��`�w��<�|>^c��XAE>�$�=�7P=��(>�S=��=��>T�>O�4����MF��n�In�>��>������G�p���&�e=�罽���`���ĆV����<��>���>�v|>�R.>���p"�x��=`L>��x#���=𼊽��=&>0���ǽ-~;ַ��n=��>��I>?u>� ?>H?�;?T� ���)IL�MUо�x��M�0���:1�žUt��D)��&���3�îH���-��Hռ$,��-�=�3>B��=ۓ>�y���=)�D>6m$>�fJ=V�D>��N=pk���G��Pj�>�v�>k�R��*�';�=P�֡���x�����'L���I���ؽ����O�*�;���4AL�ٔн��=|�Z>�Я>���>�V>�\;US_������=cB�=��ν	���.Ǿ��[�h�a�`�¾?�U=Ѳa�ǿ�m[缨���|h�R��X�ľ���k6����h>�'p��ߛ>�u�>�v?��?��G>��M=J)?�>!�;>�A�>�>A?�q?��?���>��\>jT����mm�����=��=�=->8�W>_�=�#���B= ���n
��h�=N">�x4>� �>�h�=�(.>��>FK�=[�?��>N�R�B��WZ��yG��S=>@�>)�;��\����9�n�@�ӄ:��(� '¾Q0ۼ%�	?���>��>�>a`���`�<I�B��>�5�>a)-��}½up��G6�:K�x�F��h��L��d���z��=@�n<�s6<W�>k�9?d%7?���>?�,�ވ��3?����G|��>WV��m����rw�3e�o�'�@��d$7�N%Y��2 �v��0'>�1�>���<VT�=���w����x�=L{�>�$)<�)�>e��=�T=ڹb>�f4>�#>�<��2�h���%���@�����*�<~�{���`��I�;���=-
>��N�f�����=*Zy>���>9�>�-!>�Χ:N:�X�,�^�y�@��*? ��;Ǿ15���J���/ɽ��f�ͽ!�c�s��n,0� �)�m聽�,��Ѯ��SlF��T����>6?W��f�>o ?�gc?$?n��>�}��Q�A?�x?g��>�+F?L�	?��/?�7$?,?�`�>�r�=Hw(�IP���sQ��﻽L�(=9m>�a->��=ؗ�<�������=��=͝=c�=�-�=��9>��>}�B=�t�=f=��>��.�%F&�p����=�\>��-���l>�
��u�>ȇ���1C�c��qξl���BD���Z=��=
eb>�W�>������*�=���=�I�=��>�>ɼ�N�r����v��X�=S�=;J\������z+=�=���7�=?r_>�Ϩ>�? �I?�J7?�h��bt?�\�оD����=>��\�U�e>ю�>b�<i�$��⿾g�&�ŧ�G�6��*�=W����>8#�=�:�3"<Ǘ��	�:�>�W>'�;����>K�B=��=Kj�>��>C������_=,w�J�տ�������=�
�>���=9�L�g���$�)ӊ>-��x畼�A>Hv=�E*>e�>UE ?���=����������V��������+�m��#�往a>).� ݬ=q7F�8ѽC�r�}�P��"���Nɽ#V��H��E	*���>���>/Ϟ>�ޗ>.MV=VB�>T1?c��>�pf>� �oǚ>&���J��>��,?��-?1�>�-�֘ν�L���}���+=ԩr>C�m>>'���>4�o=6΍�ne��ʌ=v$�?����s@<[�=5cɻ|��=�	>y�����;���>��.�%F&�p����=�\>��-���l>�
��u�>ȇ���1C�c��qξl���BD���Z=��=
eb>�W�>������*�=���=�I�=��>�>ɼ�N�r����v��X�=S�=;J\������z+=�=���7�=?r_>�Ϩ>�? �I?�J7?�h��bt?�\�оD����=>��\�U�e>ю�>b�<i�$��⿾g�&�ŧ�G�6��*�=W����>8#�=�:�3"<Ǘ��	�:�>�W>'�;����>K�B=��=Kj�>��>C������_=,w�J�տ�������=�
�>���=9�L�g���$�)ӊ>-��x畼�A>Hv=�E*>e�>UE ?���=����������V��������+�m��#�往a>).� ݬ=q7F�8ѽC�r�}�P��"���Nɽ#V��H��E	*���>���>/Ϟ>�ޗ>.MV=VB�>T1?c��>�pf>� �oǚ>&���J��>��,?��-?1�>�-�֘ν�L���}���+=ԩr>C�m>>'���>4�o=6΍�ne��ʌ=v$�?����s@<[�=5cɻ|��=�	>y�����;�d�>kҾP#J��=�(|S>���>Tkl�ca8>���;��h�ؾ� >MC(��O;X�𾻗����C�>t�>�S�>_����
>��[>��o����<>4w�=G(R��D������V>�;ɽmZ.��_��	�����,>ͥT>Ն�>��>u3?��5?8��A (��뾑M���A>7���v�p>8͠>^7���Ǿ�ԾLn��F۾��,���7�������=��#=A��U�&>:�=P��{�Q<�(e>���춒=q	8��x�<�L�>3��=T�=Ǔ���^h��������	l	���!�'>=�V�<s����+޾"��<_�?�Nc�M����#�%�=�
�>�a�><��>U8���r����=[�=q^��QRྃ�+�2^>����̋=�Ot��[�=�]���нӹ6��Ye��zg�����Dg��_���S���=���>�?�>|Qu>�u�>��B>��?30�>�z{>���-��>�C��,?__;?�(??�?�C�>ڟX=�����ƌ�t���=9;>]B<K>�=�J>� ��0�=r�>J;�=�R��2>�+=P��>�%>�Fc>Re���������>��@������O��н��?>v�>�ݏ>���i�l���#6��D;�0Ͻ�?�,H1�\݊�fm�=רb>8�>����={�=b��i�+g�>�½sim�k�_��M��4e;�Ǳ=��H�f�ս͂����	;�x">3�=@�>s�>"#&?�H ?ֿ����&�X�Z"ؾ2�^>�=��>�8�>h�����m�W[����w����1μ{ΐ=s�E���=A�B=8�=�y>�Y@=�̴��6�=I[>H|̽ɼI>�D(>h�=Aq�>N�!>0�<�#��p���؎��M�Ϫ|�0;)���&�qI<Io�=�G9�c�s����== >)���|Ӯ�J��<��;��F=l�\>�[)>�Z��׽��>���>�����Yؾ�����*�=��\D7>�}F���=D���2:����>�0oO��E��Z����k�B��0P�*K����>W$�>7ְ>���>��>�ӹ>��!>K��=�O �"+:<��ͼJ3n>8]�>e?+?&2�>t#��_���.���\*�Ҟ���I<��>��7=>5=��ҽ�[6>-��=S�6��5��Z3����I�9=4�#>]�>>޽�q=��?Ua"�mf0������m�J�>/���$t�>�ھ�X;$��j������̾0�<�(� �l����mǼd̈>�_�>L��]��=F(d>�����f����=sSW=8�\�ȁ?�`J =f��3}�<Ҋ���y��i�I��8�<-��=��=�+�>�>��%?�3'?{|��g�ߘ��#���Q�9��o��ަ�|/>�����վ���þ>���J���%�;i�W��(>S��=�b<�TM�#�F=L��<Ԟ�=%>���6�2��6=�,=�0>}I=쇝<_��<*!��ֱ�� ܿ;>���*0�&�U�	=�=دY<�ġ�L����9�>f?�H�0HǾK��|�=:��>~غ>>�?(��>ڵ޽,{(>f>>�[�����i�����<���V�-��
��,V9=~�� D����f��k�&���g�.����N���(��rL�}e�>���>c��>� ?2��>��!?޻��??>)X9��|>�#�>�U�>{	�>T?�
)?E�
??u&>�Jb��ke���������g��#�G>�4�=��(>�ؽ��^=&>0>>-,�=�ۮ��e����=�U�=S׼=�I=�m>k� ?�ƽ-Ý�`�>��!T��Sq�.��>?��>�W->�8�M�^��$۾�V¾�{;�i>�f�>���>��>�5?��>��h<>Ԇ�F=����5�=p=+>�ȇ>���jb=#B�>vi�=�4?="��=���ӽ�$K�4=�q{>��4>��8?2[?Ƕ?���=X�ڰ�����;Wm���<���>���>���<����X9��������ٟT��7��M�����>5�>l�^>��D>F�����Z	��rJ>���������*=�#�=g� <�%4>���>:w1>JO�������տ�'�������Vs�>�?t�=���s=��>�zm��7c;��>���=#M/>9[��$�=6�Ľ����«{��
~�_�$�7��[����=J)��>�*�����2=I�=���ܛ�����_���+ȑ�����~��V��Z�n>b��>��u>�?�=q�/?���>�-v>���=8
�������v��սa�>���>���=z�v>��p�p��#p��떽��`��ɲ>�C>ό=�?8��>�R��qO�>�\w���~<M>�!�=o�!����%2�<Yp&>'��>�9>W�?k��k�
�.��E(�� ��ˈ=���>���=���8;`�о���
=1����=^��>w��>�d�>ow�>儚>��0=C���=�W<�$�2���X>��=i�!�(�>�3N>���MX8=��'>�죻���=�hR=��=P2��*>�; ?�n?�Z?�����*�(�
�C'<Z�D�d=�¹>�?�>���=-�8�;�վ��@/�����DU���^��j> 9�=�ҥ�/<�>��=�i���*�s�>�^/�e���z�(>��u>��=	�i>A3>0�=~AD���~�Z�˿Bp��*=�A�2�ގ>���>��:�����<�!�?�7=>Ѿ5|��M��l�8=4�=9tؽ�߮��U��k�㻉>;���=69�����>d��7������!���S_�K+=�C��'S�����kK�����A�����r�@I���v:�}����s>F��>��>�S??���>1��>�Չ�Z��>J{:H��>��>g�>��>��i>�Nd>?x>��=�P���_�N�r9��D��={��=�̕=�u>��>��4=)7C>��C��=���=3��?ֽ�Y �H
 �&�����(>*�s>z?�z�=Kѱ�r����R���<L�D>jT?����Eo�=���D	��=������Q�>�t�>�6�>��>H`?R��>�q�=-W��Q��*���-��X=�3&> J
�n7�=�A�=Ԃ���P=�	�=����]���cT{;o"�=}5=z�4>��4?�9!?�I?	�W>�T&�+��hᦾ��t���ɼI�>��>f����������� �L仾�7������ׅ��&Ds=��/>Y�=E^)>���=`P#<����1�<�٘����=�+�=�>��=q=%>eK>�W�=�e;�� k��AԿf0��O��n���w�Jt�>�=�o���XV>C���R����=��S>��>M�S>6t��P��=���<u���ָ��S���pV�@.���x�I�;��n�������/�=ء�C[���(�2��1�� �8�7]�j|���h=�Z�>I8�>+m�>�S#>v95?��]>͒1>�L��'��$^<��M�4%�=�9>�>���:-�~=�%�֚�F
����V���?��>�_�>�\�=K�<��B>3d=lI>�ʽ���=��=[벽2����E�9�<�(<^�=�=�?mQ=2������&�P]��)Y=af�>��2������Ǿ��Ҿ%_��7��ڹ>��>��>��>%"�=$��>;,>�=���>>_�Ƚ��A���
>Q�>6Q�7�B�=
�½}I�������&>�Rx>α8>mO��:�v�a>6�8?�9?��/?�&��+e���,�����]�=ȏ>Ԟ�>Y��>I�>77��\�������J�'�ü���{>�2V=C�����>R�=�7���U���X=a]X>:�>}֒>���>!n>��=;���������|��0߿�軿�=�����# ?>��>"�p<���i���c��=����sef�J�>��>k�>U����$�/$�d����_��r���b���n��S�����t�о��6J�B�R�����H}�/��W·�%b��n9n�xO�,<�:�o=�w>Y�[>���>co�>MD�>�?> ?�f9�˿B>$�#���>s�<>_
�>��>x��={'��^ĩ=���;(O���	�`(��!�=b�n��R�=d�[><`>�_����=�L�;wD�=3��<�6�$��������	�۰/<�m>T�=>�@?�R�+D�VF���+�6�p�T�w>	 ?�x��,����r��O���D���0��[�>�?�Ǐ>ϲ�>��>�>O��<�n��6��=�����;�%B>�t]<)�?=ʂ�=��>=ES�+�]=�>�q�<�7>>	�=���=6܈�/�=0+?� ?*��>Ict>�'���1���Ⱦs�>��h>�>�=D��>>?�I���:����b�վ �оr���T��lZ="i�>[��<�0�=�Z޼��^��(���=��G<���=e��>�w�=�,�=A��=g�F<��=�d��s^b���ݿ����D����J�v�>��|>�IٽP���T��z��=�I���!�,�:}��=���;�8��Չٽ�E��8�>�`�>2@�<�M��ԑ��ѽp�ɾ��C�Q����;=
���b�ۿx��������כ�+�m�ۅQ����4����-(>Y�>НY>�_�>�t ?�%�>�]���O�>�.=�J�>妹>Ƿq>��p>�Ԧ=�L��]J�=Q���E�)��Z>�ǲ���p�;N(1<��>Z�=h.F>[�x=}޶�#�P�KC���V=�bU���Խ �=�W���e����=��>~k�>f�:>z�o�t�o�췠>)���㹽��;?���h���������,e�W�.����PZ�>��?lE8?�L���>�*�>:��=0��=�즽�i����@�)눽c�h�&F�=��=�0?�C��	F���%��gP<,f�;�US�*X��&�>��A?��?��(?������#_�\��y>J�a����_ԝ>���=�ś�CY �
pN��{<�.<�/>�u�½��=�0�=v�2=ƅ�=�n#>�l5�Q�-�l�=�2޽l��=4P�=8�3>�I\>C�>��=��EԽY')��,�!ȿ"q۾�I��� Q�=��>��n�ui����=$0���	/��V>���>��>���>\�>�
>�2?>�q/�>Lw����$�������#��춽���=�V~�c�h��AS�}��u?����)���>�Ek^�x<	���2=��Լ��>I�&���>⩾>�^>T<?�?�'Ӿ&��=8�>{T>wS8>4��>���>��>��>�c�=��b;e�>�H��.�}�u�<� =����1��=F}/>IN�ak�=�'>�p��֜9��	>��=����I�5=�S>x=(�=�h>W{�>ͬA���P�qp�=��1�:���U9?���X�\�n�7L)���@��'����)9|�U�=�/?��;���>H!>F�����=����W`��I�4/�=8�w�R>>-u~>�K�=����,�Ze��KW�+��w^�=o��>2�O>-�Z?io?Ѫ'?���&!�.�g�"������!�;��y>e��=��>���<���9�[/J���N��L��߸ŽI6��X�Q>��=���=�v�>3t�=�If������L=��<��u<��#>�K_>rC�>�z�>��V=m�&�C�3o�EmĿ	7.����R�=�v= k>K>�h ?���1ᾭ.��,=�(=�K}>�/>��2>0�=ݺ�=�Y��z����2�t�� ���a��l��F>�g�<�K����¾H��'C�I �pdT�]f���Q������	���>�7��sL�>'�>?4!>FFD?��?��G�?����X�>��E>��M>��>yR�>�?��>HӒ>�̢=&� >�����O:�^]޼o�A�dHW=C�<��=Y�G�"�>ZP �lj&�:��՞�=ӓ?=%��<#=4	>�s=�~k�>f�:>z�o�t�o�췠>)���㹽��;?���h���������,e�W�.����PZ�>��?lE8?�L���>�*�>:��=0��=�즽�i����@�)눽c�h�&F�=��=�0?�C��	F���%��gP<,f�;�US�*X��&�>��A?��?��(?������#_�\��y>J�a����_ԝ>���=�ś�CY �
pN��{<�.<�/>�u�½��=�0�=v�2=ƅ�=�n#>�l5�Q�-�l�=�2޽l��=4P�=8�3>�I\>C�>��=��EԽY')��,�!ȿ"q۾�I��� Q�=��>��n�ui����=$0���	/��V>���>��>���>\�>�
>�2?>�q/�>Lw����$�������#��춽���=�V~�c�h��AS�}��u?����)���>�Ek^�x<	���2=��Լ��>I�&���>⩾>�^>T<?�?�'Ӿ&��=8�>{T>wS8>4��>���>��>��>�c�=��b;e�>�H��.�}�u�<� =����1��=F}/>IN�ak�=�'>�p��֜9��	>��=����I�5=�S>x=(�=�h>W{�>ͬA���P�qp�=��1�:���U9?���X�\�n�7L)���@��'����)9|�U�=�/?��;���>H!>F�����=����W`��I�4/�=8�w�R>>-u~>�K�=����,�Ze��KW�+��w^�=o��>2�O>-�Z?io?Ѫ'?���&!�.�g�"������!�;��y>e��=��>���<���9�[/J���N��L��߸ŽI6��X�Q>��=���=�v�>3t�=�If������L=��<��u<��#>�K_>rC�>�z�>��V=m�&�C�3o�EmĿ	7.����R�=�v= k>K>�h ?���1ᾭ.��,=�(=�K}>�/>��2>0�=ݺ�=�Y��z����2�t�� ���a��l��F>�g�<�K����¾H��'C�I �pdT�]f���Q������	���>�7��sL�>'�>?4!>FFD?��?��G�?����X�>��E>��M>��>yR�>�?��>HӒ>�̢=&� >�����O:�^]޼o�A�dHW=C�<��=Y�G�"�>ZP �lj&�:��՞�=ӓ?=%��<#=4	>�s=���F=�=۾X� [�oO��@:����#?�1���A��+����%�L�Rے����=�K�>���>փ�>�s)<��>�?	>�L�=H'>{�z�%E��w�=���Z獓>Q��=�����ߜ�<�%>O>�->��]<>=>e�>i�O?/R�>a�(?�4��H��?�<����1ް�~��E��>�W�>�,�>rę�>���3�A���5������z�<�^:��=|{�=Q��=j(�=yp*>I�<p�I;��c�����<�;GFm=�=(>ew>>۵�=pC�=&烻��`�ݥ�տ�����N��r����=6�>�^�>%��=�Dv>R&:�~�ƾYE� �Z=6�>��<>g3}>��=�=�x��X���k�5=<��Ծīa�����6�����=�m�=�t������r�0�N���[~��r]��ޕ��-\ҾP���^��̏>q��?���>��M>�A=?Q�2?ٚھ�9�����>D��>G~�=�m�>z>�>���>}�>���>���=��Լ����+2y�,�\=�R/=��=�w1=>/>��u=Bo>C�K=�:�=FF>x'�=��μڌ�н���=��>>�.>d�?�ك��^	�@�o�`Y�<�?�>BT�>����¡���񽈊��zި���;<��(<���>�g�=P����4Ⱦ��A>>��=����0A=8�V����=�.]>�ͦ��%>k���w1=��>���=_���$�<Y����ѻ��=�A���@>��!?�?��??��=R� �<�=���!�u����=�!�>���=���>���h��VL�����8k�d_�=P��� !>`�=�>�<>�f�kü��">g>�:�xV��N%>�/B�6�<c��=~>���=gK3=Im���p=l*¿����}���&�v	�=ն���K��4�>:�y����>4Q;��8�5�>��w>׏�>���=���>J�n>���=�=C�_�Fӽ�ɼ����� ��e��>aAh�$J~<�JH������׽(��3E���m�?�����K�����>bn?p�Z>4 >��>��a?�/�>2��MI?�����=��>�ѭ=[g
?7�y>�k�>ٿ�>�h�>,x>|wN�2ݽE
%>n�!�Ӌ>o�J>���<6O=��=���=�s��8�<QU��=�/>�W���o�="��=���=�>d�?�ك��^	�@�o�`Y�<�?�>BT�>����¡���񽈊��zި���;<��(<���>�g�=P����4Ⱦ��A>>��=����0A=8�V����=�.]>�ͦ��%>k���w1=��>���=_���$�<Y����ѻ��=�A���@>��!?�?��??��=R� �<�=���!�u����=�!�>���=���>���h��VL�����8k�d_�=P��� !>`�=�>�<>�f�kü��">g>�:�xV��N%>�/B�6�<c��=~>���=gK3=Im���p=l*¿����}���&�v	�=ն���K��4�>:�y����>4Q;��8�5�>��w>׏�>���=���>J�n>���=�=C�_�Fӽ�ɼ����� ��e��>aAh�$J~<�JH������׽(��3E���m�?�����K�����>bn?p�Z>4 >��>��a?�/�>2��MI?�����=��>�ѭ=[g
?7�y>�k�>ٿ�>�h�>,x>|wN�2ݽE
%>n�!�Ӌ>o�J>���<6O=��=���=�s��8�<QU��=�/>�W���o�="��=���=�>��>TQ��v"��վJ�1�#<G�>�n?�F�Q�\�P�Ծֈ�T���ҏ����=�=7���T��9/��왁>E�>�=���=��B�>
3>�	�< B�ПO>��<[o�=E,>�4=XB�8����g{�ũ	>9D�>;�1�6�}>k�,?	�?W>?�k�"�J�=�#�)�x4�=�=j��#�>���>���>4����	���Ͼa`�����U5M>��D�T!>|X��y�b��\!>��ɽ�Z�<e�I<(^�9�%���>«�&P�>���>��%>�*�=ߡ:=����-/ǿ|������/���@(>�������I�=%z��1#��,2[�&�>�v�����=�%Ƚ��w�9˫=Z�>��	>.B�=a`�U٠�tF=H�K�|�3mD���V>z*���r�<YP��`��.ç�,�<��=J���췾P��ޕ)�MlK>���>��>%O<�(?p?���>�C�#\d>�p�>�0�>b@�;���>�{�>��?.J�>�U�>�_p>��>���� 8��[��=-�Ž/�F>K��=�q%=&�=�Y�S�<pC����=�ʍ���s�����'>,}=�Xh=�je>(�>���([�@��aC"�o��q�B:#f?O�����~��</�1�lȾ@H��ѭ�=������䯾إ~�Q>�>{+>{��<�4>�,��;>8:�=@�9�����f��=��>�g˽XS�<86�i�������=)`�<n�W���p>��>j�??#���WF9����4ټZe=��~<��v>E�*=E�߾M	-��X�i���8��o�I������>����&Ἳ90>�ڽ>(��+>N�f=G�;��� >��Z�h�=���>kT>��$=Px=��u�TT�z-�!���(��6꾖�=ul�h�A����ǆ*�ӎ�>�����n��������>�>�����8>M;>�B�>�[�������N�x@��Ї��e���u>J���3�F��C��5���S����ڽ�s���8�= a����=z�>+�}>5�5>�7?-}�>��!?iL��� ?���EM>MCn>���>T��>߹�>Y��><��>�r�>�B|>�9#�VdF���;��9��H>�mH=ܹR;��K>W)7=���ecD>�@ż[Bl��'�����=4�����A=e��>�?�,���	�bWǾ�O���Լv;�=���>�|����|M�v����k�cێ��[H<DCս�j
�Е���n���z�>�%>�ޕ�h'C>�	�.!>ŉ�>��7��J�=�R����0����:��<&^D=�C��`4<>�އ�As{��<:(>VJ?ơ?EuC?u(����⾌���l/��W�Q3</�>S��=�>L����f*��*о�f'��.�![>A�>�:��>(�>��=�@M>�S��8�Z5��{�)=zD7��=��w��y?�>�I">	{�����=�Q��-��;�j׿�I���\������[��=f��̿��>�>uf� �o=��
�FD�="����=���5h>5�G>��>ppW����pg���s?���h����(꒾I�ԾK�>2��Td"��7�B5>�g��<'20���������ʽ(m�=ԡ�uQ=���>�(<{�ս"�q?,�=?��-?󼜽�>�`}=8��>D��=#/$<*:?�%4?�k�>l!?/��> �>�*��{��ir�<J��p->��<n�U���=�f����C>j:�=���<	~��A׽��r�giϽ+BS>��'>�d�=�)�>Y7��H޾��/���O��5>��>.�,?��+����=�����v ������ܽ�bھ>�J�_�6��;�>�/�>�eR>BJ�> �<C��=��ƽrț�H�_>��ӭ���>�~B>��z=���<�Ҭ�����*�a>�=��Y>���>4(>
�B?�MR?�>0?��7�f3����$�C���0��%�?@��O�;~0�	��ƾ�۾��8�l$�=N��<��=Lys=O~���<����1:���=���=��^Q�^�>���=R�[>���>2v>D�>�y	���Ծ�ۿ�a��j�`��U��P6�J�Q�Ы>��R>�O��b�P��+��Z��;(����#=w>w��>�s>��-8��ʵ��P���M���C��ڭ��tf�c���%�:>.�!�}���s��-6�-1��Q�w̢���B�h���=Pe� 2��Υ	?��>Y
�=���>n�[?�>�r�>#��zV?ځ�>˔{��?�O?�#M?:{2?Y�.?5{L?a>�>ɯǾ�� _���%�;c�=��>�>�ON>��p�-��;����=]�����耼�&1�R��;��==�=��>�(�=��־/$վ ~9�>�:�[H/>
q�>��>�%�|&꽝"���b�����<��s��y�+5�L(��Ye�>'v}>���>'ʶ:Y?>�AG��|d=#�
>*f	��YW��8;#q_�l��<���^�2CN����v׽�U�=@Y�=��|>�Z<?U�;?ZD?�G���?��y�p� �i��	?�wa�>s=?��>h,m�%�c�M�H������y��������=�u�=��">,���5M<X=GM@��go��+>���=��L>�>�c9�:��>I��>��>�}->,�U>���:�����ܿV巿����!!���,=������o=6�D>~Ƚ:����Ͼ=�B�4���>�`e>�)��1�^��`�=��>w�����Ͼ��h�����ܾ��H�1�о��=	Ƚ�;��d�'��;6�H��6�<�(�ܽ������-����?�?>�n�>YMR?Hj�>c֞>�DT>��6?���=�*�=���>߾�>��>2�'?��:?�[?�+#?7�8m�����|��=u =�<U>��7>��>y�����2<.w1=��=�M�=y�N������>���C��Y>>��=��>�)�>Y7��H޾��/���O��5>��>.�,?��+����=�����v ������ܽ�bھ>�J�_�6��;�>�/�>�eR>BJ�> �<C��=��ƽrț�H�_>��ӭ���>�~B>��z=���<�Ҭ�����*�a>�=��Y>���>4(>
�B?�MR?�>0?��7�f3����$�C���0��%�?@��O�;~0�	��ƾ�۾��8�l$�=N��<��=Lys=O~���<����1:���=���=��^Q�^�>���=R�[>���>2v>D�>�y	���Ծ�ۿ�a��j�`��U��P6�J�Q�Ы>��R>�O��b�P��+��Z��;(����#=w>w��>�s>��-8��ʵ��P���M���C��ڭ��tf�c���%�:>.�!�}���s��-6�-1��Q�w̢���B�h���=Pe� 2��Υ	?��>Y
�=���>n�[?�>�r�>#��zV?ځ�>˔{��?�O?�#M?:{2?Y�.?5{L?a>�>ɯǾ�� _���%�;c�=��>�>�ON>��p�-��;����=]�����耼�&1�R��;��==�=��>2~�>�1��z�O�}��La+�-�>�ٔ>�t�>׈Ͻű���ľ��c��b�/��=^���?�]��#�>���>M��>xB�=�}J>W�C>��D��4M=\��>x)����~=z�:���=��!=����?�콴���~e�=��\>F��=;�>t8>K�??orX?0~S?����Tꑾ�����=�8D��!p>���>q���}��n�)��@̾��㾌�������<̲?�<׃>��B�&ۯ�^~>���EE�����>�T�� w>?	f>�����>C�e>���>4bD>d��=p���oǾ����k��m�d�H10��>+=�[��3��I���-z�>�q>���8�T��(;aB>��>�JX>=*�=/+N��Y���3�?s<�U�v�ľvǚ����������>�
��U�2�Ѿ�B�=�߾��鼺�{��B��޾�z�u����?ܢ�>�e�<�p>��`?p��>��>���>��>������>!�
?��0?R��>��B?|G?�cT?`�=�q���5ܽ}�U���>�y)>�q>���=�>��*�}�=;�	<�0��̓漯5�;�ʽ;�<��$!����
�>�C>�=>#*�ǻѾ>��|9��rG��� �{�?6x�����a��������ҾYG�2��M����+����=�x��%�P>�	�>*�=�}=i��=��%�B>�{1�N�.�Z#�/�9bR;�0���)��3����	ཇ==�PE<>�'�>D����;I?rb?+x*?[a��{;0�Q��v�:����f���j�>,r̾������yF�'�4�*ݴ�R���m;N>�j�=�=A ޽w_����u;�v��_���g>��=|�=<X>�,>iQ�>UZ�>A��>l�5>͎Y>2����о9���ٖ�o�*��'��~6=�Ԁ=-��:s�4>�ɐ��:�=n���ߍ�17>ݶ=�}�=oU>�v:�r���!?��H���^�/�d����׾�
��\�� ݬ=�r�=bl?��5Ҿ'�#��.��21�P�1<*�N�ƾ��L�i��R&?E��>٩ӻ�[�>�.\?P߷=�� ?�
��V��>C[�>T�>6c%?��.?�k!?�(?L+7?��C?��?��I���[D��j/�=��>��">R��>T�:>�|���w2=V�Z����=��v�H��=�;�o����}<���=� R�mĝ>�5?�'�o�����c�b��'��i�Y�N�)?	���7�=>�����g�����K󵾓��'�۾ʔ ��?n7�>`�d>��,>'�p���7�=���<C>{O�=/��m����B}�M��=�L>�Y���A�<���E*M=	O�=H�Sh>�W?��>��?�&��OV߾(.
��A������C��<In==�u����n=�����B�-�Ͼ����. ��哽-��ӗ�=���<�^L>�� ���ｵ���>���<% �=%�7> �J>�3>�>�~R>j]U>���<haɾ3髾[�ؿ�v���kA�l��՚�9F�D���%e��+=��h���$v�별�m�e=v�2=��=��0>h��<��	=�V�l턽#�]�BA�����L}�٪�%�=�a��%���^��z�+���Ǖ���*���5�]a��$��=��O>��?Bh�>l�C>[�3?���>�j/?gM��T�?;��3s=�kj>�0?!7?��!?�]2?���>�������]�%�'&u��'>���=���=��[>p�=�x��߅>�U=���=Ap�6r�0qD>�s�<"Hk=k��<��>�XG>�5?�'�o�����c�b��'��i�Y�N�)?	���7�=>�����g�����K󵾓��'�۾ʔ ��?n7�>`�d>��,>'�p���7�=���<C>{O�=/��m����B}�M��=�L>�Y���A�<���E*M=	O�=H�Sh>�W?��>��?�&��OV߾(.
��A������C��<In==�u����n=�����B�-�Ͼ����. ��哽-��ӗ�=���<�^L>�� ���ｵ���>���<% �=%�7> �J>�3>�>�~R>j]U>���<haɾ3髾[�ؿ�v���kA�l��՚�9F�D���%e��+=��h���$v�별�m�e=v�2=��=��0>h��<��	=�V�l턽#�]�BA�����L}�٪�%�=�a��%���^��z�+���Ǖ���*���5�]a��$��=��O>��?Bh�>l�C>[�3?���>�j/?gM��T�?;��3s=�kj>�0?!7?��!?�]2?���>�������]�%�'&u��'>���=���=��[>p�=�x��߅>�U=���=Ap�6r�0qD>�s�<"Hk=k��<��>�XG>_t�>��9��ㆾ/��]پwJ�$L���>Y���C<�\�=�@�=�~��,Ͼ.�m�Ӽ� ���K�>g}{>9lx>$��<�P"���= [+���n�~��</��|?=��=��>�.>:<�����E�=�>|�@������B>x?�Y=?d�?���=����x��6־	�ѽo�>��K=e	����	�҃�lM&��h�~�þ�Lξ����ؓ���=N >rv><`XC>��=�`q:\���s��96b�;�;ET�=�6N>�-�=�1b=A��ZE>(�=s�D�c�߿���/�=��3Y��|
��ܠ����=��e>�^�������C���Y��d�>b
->�a$?uy�>ˮ��Ñ"�{d��U=�0���Ӄ��U��R������e2>���ɽW���9Z �1�־�͡��Ց�D�$���'��L9���ޚ>���>�\>��=a�?
�?�U�>� P���=�)��A�>�V>%��>�Z	?�+�>̏�I�>Zׯ=�w;�́��:#W�
�>O��=��>�>�)>�O��+
>e���mo>���;�#��=�n!>΅�=a�F��~Ǽ�N�t3�>�5?�'�o�����c�b��'��i�Y�N�)?	���7�=>�����g�����K󵾓��'�۾ʔ ��?n7�>`�d>��,>'�p���7�=���<C>{O�=/��m����B}�M��=�L>�Y���A�<���E*M=	O�=H�Sh>�W?��>��?�&��OV߾(.
��A������C��<In==�u����n=�����B�-�Ͼ����. ��哽-��ӗ�=���<�^L>�� ���ｵ���>���<% �=%�7> �J>�3>�>�~R>j]U>���<haɾ3髾[�ؿ�v���kA�l��՚�9F�D���%e��+=��h���$v�별�m�e=v�2=��=��0>h��<��	=�V�l턽#�]�BA�����L}�٪�%�=�a��%���^��z�+���Ǖ���*���5�]a��$��=��O>��?Bh�>l�C>[�3?���>�j/?gM��T�?;��3s=�kj>�0?!7?��!?�]2?���>�������]�%�'&u��'>���=���=��[>p�=�x��߅>�U=���=Ap�6r�0qD>�s�<"Hk=k��<��>�XG>iw�>q�ƾ+/龊�̾��\d>?V=]��>#k�=4��C�f��<�����N�= __>��h>�o>hc=o��>���>22н����C/R��
��ç̽!��>�X9�G�L=�k>��i��R���_̾�����=��=v�!>�{>w>B��<�d~?�c(?w�s?V4�>f=�����_D��iݽi�r�>6��>
��>b2e��*���c��D�M�ݾO�����c�F9&>SQ�>x۠=�N�=�qνW�F1�Y�/>0�<�a��> �>��>�Tn>�4I<�	��O��&���Ͼ�n���n���Hs��{ɾ!�d��K����½����V��'P�=aR�z����h������
�C�K4<��>�N�>&�/��d�����,>tT�=�1�y��;}�U�3F����m�2�a�7~���#�#q�8se��.��6�Y�q�R�^�]��N(��u�>��d>��<(��˕�>��>׭�,i�>3e>�C�>���<m;��&>~��>]�?̷?V}S>���6��A�;p'b=���Ö�=b��>�UB>b���%��>��ĽjX�<�_��T�>l2P>�E��Y�>�����=zm�(��>0��>��z=�FK��\¾�T�պR�{=n�=.藽}��o�;��� ��������=�͐>��<>Ƌ��S༣�>�c2>�P2�h���=LM>�`=J�W=����_�#=�� >�A���<�-��]d<�\>��>���g]N����=j�'>��9?MyA?�?�B<~��=�C뽧���e��p���E�>���>��O�����h��E;��������̼��Ƅ>��:>%@�<��i��H��=֓j�>��={ʂ>3�=Ӏ'�C㶼s�h=��>:��=^��;Q�B����i˿W���<��إ���>o׾������>`�>��>��=�"(>��>�2>ǩ��n���
�b�'>2>8�=p��c�۽��=UB��M������Bo=�6��ه��)��=�<]N6�%��+����<u=Ƚ}��|	-<���>�o>n��=�+�=�]6>@@�>^��>6��ݭz>��[�U%f=,� ��e(�*�c>a�>K�e>��n>)oH> ���A̽�	��0��=��Q����;�>��=��y=�Q8��'��g�=�r�=GE$>�jK=�i���i�9-�=1�G>��u>���>�&@=����oѾ�������>]�Y=40>�� =Cvʾ,	�����"̺�G�>7��>o��=�+��(X�=��L>��>w��<�2�=�| >}���]%<wh��ޒ��:����/>�=����}�)�dKm�|����<e�9>sa<�O>54R?o@V?M9?�s�>릤�W�ؾ�, �^"�w�ɾ�T>>b�=�Ʉ�ڸҾ�������S����S��n�>ҍ�>�$�=�g�=��ʽ���:�<r��=�k&>��P=4^��4=3�=,y>,�>�.�<�{��o㘾H˿�����Σ�#�H���[�颔=W��U�>�i;�� ?��>�8�>Z֊>Lc>|=��"Uh���6s>����<y00��k���hK�zw�ر��1P���T�=�Y���Vv�S�m�0�=�'$���޽Ƨ潮*b�˅�:콽�z$��F�>�A>�痼Wic�> r#>K�l>��E�>��A�C1�,YE=�$>�қ=W|�=��9>
��>�>�ԋ��&���i�d��=����|x�2
>�͔>�;� ��8k&{��^Q�����m��=q�t>n�>Y����	4����=յ_>q6�>�Qb>PA�\���(i�=r��^4=@���� �������hzr�G>���;L�>��O>.=˜v�q	�={��=�l=��a��?=��J>�8,�d�;���>w�������>���=�,��|s�U����Is=�=���<�!�;-��>;?�&H?��?;�:>��!�vS߾b$���E�����=PC>�o���yC��ľ�	����͔�"�:�B����>��7>�Σ�X�ټ{t�=�@����V=/�>��;��	��ݼ���=�p=
_�=�U> A6>YT�3����Lп�����6��;)��`Ƽ�$������P�>���<�?ע�>�,�>�z�>'�=	(ֽ(Fu�F���s�sm>?�A����s����н�	��V����̐�BTI==�����g���C��sj<:�U�͕۽g�-���ܻm�ֽs���;��"^�>���>�=�=�z�=�qh=��?>�͏>��'���>/><a��Ϋ)�����c=��>>�V�>���>I�6>TŁ��2�;����,> /=I�;`>xc>sl�<�r�<���=o'������>��=��= `��,���=���=і�>�ɔ���e�Vk�����[>D0g>�s<Uܼ��Ͼ����@�>��\�J>�A�>�)�>�b$>e�L=�G�=�>����,ƽ|Ѽ��Xk���F������հ=�X!>� ��9�ĵ����2� �=ީH>�P�=�nU�if���>��Y?�(?Y==?9`>I�����A��de��TB���p�>�^�=}m(=d�̾���2o�J¾2i;�9ž]>Z�hUF>�G>Ш�=E�)>x�>�j=>[�$Z��� ���oV>�>��=A�=��>7"�<ª���q��.���N˿�e��.��@:�:[=�N����)�>nB\>�S?bM�=�&?��>�j2>s�����a�v#D�ot=���=PA�=��u�}ޠ�b�8�����B5���0������.ּ�W<~�x���Z�w�ѽS���^ֽ�ӳ�B�ὠ�,=�ض����>�/=�" =�=<�i>8��>p��>�+�<�Q�<��2�@���wu����=��>���>�$\>�/�=�C�=�uS>r<ż_�Ƚ��U>^�	>D��="t�>)�6>e�>s��c޽eX�=�:�=���>�B>&L���S��.�<�+#>�:>q6�>�Qb>PA�\���(i�=r��^4=@���� �������hzr�G>���;L�>��O>.=˜v�q	�={��=�l=��a��?=��J>�8,�d�;���>w�������>���=�,��|s�U����Is=�=���<�!�;-��>;?�&H?��?;�:>��!�vS߾b$���E�����=PC>�o���yC��ľ�	����͔�"�:�B����>��7>�Σ�X�ټ{t�=�@����V=/�>��;��	��ݼ���=�p=
_�=�U> A6>YT�3����Lп�����6��;)��`Ƽ�$������P�>���<�?ע�>�,�>�z�>'�=	(ֽ(Fu�F���s�sm>?�A����s����н�	��V����̐�BTI==�����g���C��sj<:�U�͕۽g�-���ܻm�ֽs���;��"^�>���>�=�=�z�=�qh=��?>�͏>��'���>/><a��Ϋ)�����c=��>>�V�>���>I�6>TŁ��2�;����,> /=I�;`>xc>sl�<�r�<���=o'������>��=��= `��,���=���=�j�>����� �x��,��)���>�?VQ��n<u>ԅ��'QԾ��f��=��e�̽����]r�>{��>i�>��>L�j>�H>�Uc�������k��ߟ=��0�.9>�T��V��je=;s����j���,��l�>C�}>hH�>l.�>��(?�O?A�=��˾.�6�R�T����OU=�!l<wft��k����'�[��E���+8�5�o���R��w��)�>_ˀ�g�1�w�>Vyf>A�e�>�O>W*Ⱦl�=� �>zgW>�j>���>��>�J>>������9�ǿ�����:�����Il��0?��>r��IR�>�֠��o>�>#Eؾs��>�^�>Y=��>�/�����>�{�#۰�u�a�F�������-+��~���ź73����c����|�Kߣ9D0:�4�o��i���V��<���>g+9?D���)��~�C?E�>�(ʽ���=��>��=Y��<
�x>�1?MZ�>O�-?�8?��?p�ٽR+��巽�	 �Є>T��n�=��=�n�>��ս�{��]E�>刄<S'D������S5>��>�?0=�m�=��>w�>�??�/&��R�=]4j��s�u���?=U�>��/���������"�A��~ؾ�� �d%�>��B>���>���>�*>�>O�9=��<�z,���罭���N�����=EE�<�=��|<��f���<P^_��ŉ�`w��L�<�u��Cy�>��v?M��>�>5J2�(��-��ݳ��)�F�A�(�~=
M�>Tn#�y>�%�ᾀQ0��Z�\�7�S����Y�?�<��.>@��?L�>Op�>:V���߷��m>k�󽌢9�/ ���%y>b�+>��r>��k=���ȕ���[�c�ÿ=����� !����=�Za>Q@�g��-���	�>���>D���G
�>q`�>�d���'��H�>q�p=�q=9�Dր�����o���¾��a��>����
<RA,� j�2H\�z,��i���=�ǽ�$��"/��r��=c�y>;*�=���>eR?Z9?��>�����F?�w=�(`>�W>��A?�y�>Yy�=�bp>f��>w�D��$蝽�h�7�-=Յ;=�5��"�=F�=�.�=�%��G=	Z�=����K1=%���z�N�D=؇/>�fN>k�I>�j�>����� �x��,��)���>�?VQ��n<u>ԅ��'QԾ��f��=��e�̽����]r�>{��>i�>��>L�j>�H>�Uc�������k��ߟ=��0�.9>�T��V��je=;s����j���,��l�>C�}>hH�>l.�>��(?�O?A�=��˾.�6�R�T����OU=�!l<wft��k����'�[��E���+8�5�o���R��w��)�>_ˀ�g�1�w�>Vyf>A�e�>�O>W*Ⱦl�=� �>zgW>�j>���>��>�J>>������9�ǿ�����:�����Il��0?��>r��IR�>�֠��o>�>#Eؾs��>�^�>Y=��>�/�����>�{�#۰�u�a�F�������-+��~���ź73����c����|�Kߣ9D0:�4�o��i���V��<���>g+9?D���)��~�C?E�>�(ʽ���=��>��=Y��<
�x>�1?MZ�>O�-?�8?��?p�ٽR+��巽�	 �Є>T��n�=��=�n�>��ս�{��]E�>刄<S'D������S5>��>�?0=�m�=��>w�>���>4�%>����KZi�ޱ�����ݡ�>�&�>��"=�Z���1<�'�����ѷ�i_:���{>���>��> W��D�=_�}=^��='J���阽 �=��9=��=jW>uw���<b��=�+�=�~��G9�;;5����[��>��y>�Q�>�?0�?U��>�{�>��o����L��^���CP����~=5?
߅>�j4�֜�����*ؾ�1�>.����=�fB���<�؈>��<�v=�Mƽ���@�=��=�&�7D�=
'k>�K>'�=�ו=�����֔�u�տG����.�9�	�6혽��<��C��e���]j>e�>m�$>�J>���;Ǐ�N�2=�O������pqν�'����>�K�=�{��}ҽ5�	��v���v�uŽ��w��w��Z��P2�-}��+�~*E�ǐ��8�3�#N+���н�\�>D>cħ>ĝ�>�kx>��?���>v�~=6�='VH>��#��!��4=�w>��>�.�>\��>
~�=]�<��b��!S��q)>�7�=��4����<=��<��=ct�=�*=Z��=���=�rD;�i3��'�;���<��W=�N�=M�=�??�/&��R�=]4j��s�u���?=U�>��/���������"�A��~ؾ�� �d%�>��B>���>���>�*>�>O�9=��<�z,���罭���N�����=EE�<�=��|<��f���<P^_��ŉ�`w��L�<�u��Cy�>��v?M��>�>5J2�(��-��ݳ��)�F�A�(�~=
M�>Tn#�y>�%�ᾀQ0��Z�\�7�S����Y�?�<��.>@��?L�>Op�>:V���߷��m>k�󽌢9�/ ���%y>b�+>��r>��k=���ȕ���[�c�ÿ=����� !����=�Za>Q@�g��-���	�>���>D���G
�>q`�>�d���'��H�>q�p=�q=9�Dր�����o���¾��a��>����
<RA,� j�2H\�z,��i���=�ǽ�$��"/��r��=c�y>;*�=���>eR?Z9?��>�����F?�w=�(`>�W>��A?�y�>Yy�=�bp>f��>w�D��$蝽�h�7�-=Յ;=�5��"�=F�=�.�=�%��G=	Z�=����K1=%���z�N�D=؇/>�fN>k�I>.
?�;^��e1�p� ����݄��D��KH;>�Y���M>�ߎ���Y�2�߾����0=";	��
�Ę�]�e��<f>\��>|�@��f��>P!����<��$<o/��� ><2y�-A�䛁�|`�=%�B��iB��tY>��al� v�=��z>]Be?�sR?���>)��͇������B���j
��Q4>�$Ҿ�/<��,�����4���Ǿ���ʝ˾$F��u(>ؚ>L3=�p�=.ç=j���h"���=����x>X�}>���>#��>��>�O>X>�}�XU4���¿�Z��U�D�髀��\^>���<mB��E�>I�uI�>;������>��;�s0>�
���n��NF>�a>���>4�z�3���_�Ф~�s��E���m���d>I�8��J>y���Rp>�Ԗ�2�X�����cν��쐾eE�o����V�>�*�>���>��	?n�?x;�>��>�(���L-?��н}��>?�B>�/?�j(?2��>�u?�n!?�?U�=>4B";�B�'߾;L��=+�=`(>�ɂ>D�Y> 
,=s�>	�=����[^����|��D��Y{���>�=�O�>_��<i��>��ؽ�E;�'����ݾ���`U��Ə�>��&����=��þ�Nd�%#�����"���,����׾;�v��
�� �>N|�>5;͸�<����ôټ��]=��v�r��Q���)Z>���D)�<�N�D��Z�<ƚ��!���ս�w>!o?�!S?��
?"��g;��H"���w���F�h��I�]>����>��>覘>݆�{U� �,�C�#��0ݽ�fO>�s�=2:�=U�,>�)g�[\��T���%�>+>��>���>x'�>TS�>���>�$�>D A>>����ӽ:mѿR|��C��Ҍ�J��>w���Bl�=	?a��6Z?�P�9�?�g���˙�>�Խ6�>��"�2rZ>�)�������輫�>{=��m��現��>{�(>^˾K$=F,i��S�M=�BJ������v���=��J�>�z�>���>���>F3>�?ON7?��F�U�?v�B�N�?id���>�'�>Fp>�&?f�?c�*?���>:i�,ou�?�������<�m9>'�>���=�8=L�=M����ӽĿƽ������:<���=,E:>T`>�E)?��vJ?���6�+i����<�)�=H;�=p04���>����8���@����I��Q̾z�Ӿ62)���>�L'>��n>/�@>(��=^�>د���㢽�r>7ݘ�9���5����=�:��GD����սP����o���^��lU>��>_�{>��]?4G?��$?�d��.�������?��S����B1U>��Ⱦzm����E�.]��wƾ�Ա�d���YG��nr���:}=OZ=� ��TI>��3�}�9�}��=.��>� M>�u>^�>>c�G>s0�>,��>U^s>�
X>�tb�q�a��ɿ+m��Bb��ou��Ҷ>��>yg��{�?
� ��>a꾮E�>�C�>�Ɩ><3�>-�=�r�>�0���=��轣����VF��(�\ o<��C��T��f���G��:�=�����w<p���`�2k��իٽ�H��wc���ix��*K>�>HQ�=9�>��>���>@��>�>(IO?x�G>�5�>8��>I�>��?���>�=&?�?;�=�	������G�5ے���=���='7_>�L�>�->Iݡ=''�����=O�ɼ �ŻzV����O��u=�!t>{��=&Z?��}�0_-����KM��.�������>n}���x>aV����Z����ֽ5��Ҿ��0%��^�>��>��i>�b>�c@��=F%��\w�=��
>�4��aܵ�pr3�q�>�^�l'�<sb½	P��G,�@����I>9��>$z	>��Y?�{=?�?lV���_�'���6�s�<(�۹��Q���k�=T�����
�*��fP�F��`�:�	*>�¿;c=?��=I�`���	�Ŭ)�հ�>�h�<��%>@ƍ>�g>�]�>%�>��>Dq8>3� ��R���ѿ�Ҥ������D�F�ǽ��<m�=��>���8R=�1���>�F`>抍>�4�>zw�>�>v��<�=p����00��7h<�&��tZ�d8v�����O�o>h���Mn�������Ƽ�nJ�=�(�kކ�c�F�s^��ݩ�b�K�p0!>S�w>��>�?�ޝ>�?��?�����?�D�>B ?���=�"�>�E)?�4?Ց??��D?bp���O���q�A���/��<u��=�Α=�%a>[9>u���9����`>�Nd=�eͼ������1`��po�T�<u�=�<�=�y�>�0���l����t9޾SP��a=��=�&��>��l���p���������܂����RQ�Y}�>YUE>uv>��X>.6�;��4�0ė�>>�ѽ�m��v����<>�}{��T�=��������Ɔ���	>���>�d�>lJ?}5O?BJ?�\��(��x��.1����������>҃��ߘ�= �����Ub��2ɐ��2�jh��M-�a[>7`�vY<D�v=$A�߭�!� >�B>h�3�>>,��=��,>�N�>c�>!>�Y�<cd����̾��ʿ�b�����X��+)`>��=�C�>׿�>v��<e�=Qp��sw> Gܽ��>yA�>��>W�2>m{�=��=Ԉ��xE��k����=�L��O��� �>E���	>L,羳YR>�儾�6�����y�A�@�*d��1wf� �>[�[>�s6>�
>Cv"?8��>';�>��>��+?n4A>��A>�[�>s��>O�?�*?#?�,:?/ʝ>���qt���S���<>k6�=ha>B��>�o(>�:D����;�<��Ǽ��½��-� ����f��y�	= �H>�]T>�@�>9��>��{�8��*x���)��t���u=�l?�p�i��\����6�<��2�E�<�:��M?���!�=,0��O���>���>Z��=;�=mG+�Ħ�=d>b�<�<�ҷ�=Ϊ�=�w
>��Q=;��9�q�=���bܻ�2�I�Q��}>�W?�t\?'J?�ۼa���@��3"�gξD��>�2?���>-̖>��Z�uþ;[��[Ya�c���v� _>����=d�">�nj=f\�>��L�V夾葂=%�>�t�=o��<��=�2V����}>�I.>�-�1IK<��$�h~3>x2ݿe����i ���3��	�j����O=F���o25��8��`���J̾gŽ ��>�!?��>n͋>��6>�x�>�H������sb���i�1�-�gg@�BkJ��V=b�%�$�:��d���<�ZΞ�^y��i
������Z��	=�,�=ճ>�0�>S��>���>T�'?�p?��>�Q��?�;>A�<����>Ng�>���=>ϔ>�L�>��(>Г�>-�&� �V����<��9"�8=�n>X8>�0νʌ�q�'��)A���m;,C�;��<憲<�=!E�=��=�9�=�Tp=��o��� �y
E�Τ,��jȾ{6v>��?�-,� |�ک��n<��B�1����=�2��-���	��ዾh�N>���=[��	) >�
�=��d>�S�=�YP�xX|�z�T=���=X����������@K<��_�[���P���=��!���k?�Hh?mV�>����rҾҵ&����K`Ծ��^>MЍ>4u�=`�>���=p͓�<9���.����|��y�P=�<M>�:�x>79�=��{�v���1>ɯ@=�}>�>�>����O�>C��>O�m>d�I>�q�=����ܟ�ăQ���\�vL��|�=V�*�&��=~X?�D�Z�o���~���슽�'��,�=��ؽ�6;�9�=�s?��E>2˾����f�v�:���޼�*��>���<r].�l�q������.>y�h��?'�P��:�&%=3���j$�_�[�"�>@��,=��?]�?�*?@�=��1�n�?DC�>S�>��Z��>2?�S�=�+�>��?���>�?�>5N��J=Y�=�ӽ	�=����]8>r�`=�W->��ۼ{Sϼh >��μ�ڽ<��<�rս��x=���=�`�=9��>��{�8��*x���)��t���u=�l?�p�i��\����6�<��2�E�<�:��M?���!�=,0��O���>���>Z��=;�=mG+�Ħ�=d>b�<�<�ҷ�=Ϊ�=�w
>��Q=;��9�q�=���bܻ�2�I�Q��}>�W?�t\?'J?�ۼa���@��3"�gξD��>�2?���>-̖>��Z�uþ;[��[Ya�c���v� _>����=d�">�nj=f\�>��L�V夾葂=%�>�t�=o��<��=�2V����}>�I.>�-�1IK<��$�h~3>x2ݿe����i ���3��	�j����O=F���o25��8��`���J̾gŽ ��>�!?��>n͋>��6>�x�>�H������sb���i�1�-�gg@�BkJ��V=b�%�$�:��d���<�ZΞ�^y��i
������Z��	=�,�=ճ>�0�>S��>���>T�'?�p?��>�Q��?�;>A�<����>Ng�>���=>ϔ>�L�>��(>Г�>-�&� �V����<��9"�8=�n>X8>�0νʌ�q�'��)A���m;,C�;��<憲<�=!E�=��=�9�=�G ?�6޾��0�B[
��QA��+��HI�>�u?>ncټj�j�Oo����G�M�꾝��L����;	���S�G<p�a=x�H>L�x>#*�=$�x>W9�<��=n��=S�d�Q��=u��;�#v���M�ϽGY�[���^i�R���p�<Ʊ�=�gO?�(?b
?�R�Ϻ�p%�^��X���"{>�P�>��F<�w>���4�2��]ʾ�i&�;)�:}��豔>\)5>�}�<�=>�~��}�#V>q��=��;��>�>�
2>��z>�r�=�D�>e��>�ڧ<����h(¿I��t�侄�8�mԼ����p�;t_�>�y�<�о̩��J�������i�#����>pc>j�=�q<>t�->���@��n\����Z
ž�6+��D���*6>#N��qN�=
��h*>G5���0���:>~�u�"�����V='�Q�N-�>���>3��>?�8?z0�>7�>���t��>-J�>�>�^>�m�>!6?�4=Uĭ>I0?���>(�;>8���u�u �.��<dW�=��_>.5�>l�P>ݞ=)d��
e.��G��(�;�������=��!>��D>9��>��{�8��*x���)��t���u=�l?�p�i��\����6�<��2�E�<�:��M?���!�=,0��O���>���>Z��=;�=mG+�Ħ�=d>b�<�<�ҷ�=Ϊ�=�w
>��Q=;��9�q�=���bܻ�2�I�Q��}>�W?�t\?'J?�ۼa���@��3"�gξD��>�2?���>-̖>��Z�uþ;[��[Ya�c���v� _>����=d�">�nj=f\�>��L�V夾葂=%�>�t�=o��<��=�2V����}>�I.>�-�1IK<��$�h~3>x2ݿe����i ���3��	�j����O=F���o25��8��`���J̾gŽ ��>�!?��>n͋>��6>�x�>�H������sb���i�1�-�gg@�BkJ��V=b�%�$�:��d���<�ZΞ�^y��i
������Z��	=�,�=ճ>�0�>S��>���>T�'?�p?��>�Q��?�;>A�<����>Ng�>���=>ϔ>�L�>��(>Г�>-�&� �V����<��9"�8=�n>X8>�0νʌ�q�'��)A���m;,C�;��<憲<�=!E�=��=�9�=�H�>�-�����`0�~��������>U��>��X�wAʾQV�>�g��Ѝ�b,�\7'�a`��i��>��?Eg�>��>),>�����'���?��mU��� ��5E����>ޕ5>��˽_O)��v7��!����F��:˯�=!I>@�H>,}[?F�?��>�跾���O�p�w�C�����O��==��>��Ǽ�g�=�R����F����F�ݾ��b���ʾ[\ǽbX�=�=�ᗽ�8r>�K�=��ƽ��]>�	=�Q�/���<x�3>��>��>�J9>˨�>w������5�տ����_�:�g��)I�>,-"��� 5����<>+���,y���7�"�#�UYq>�}\>z��>`��<�C=O�$��bK�J���s�3�?���L��3��A�q~=S�ܽ#^0��Fʾ��=C*� )U�O��;�U�7M۾FsJ��_}�qM?��>�?�?|�?��>?JJ�>�<*>N��>i��>�?�����>�ј>��?��?}�5? �l>����,�,�
��&��w8P>��x>Ҡ>��>a�彘�)=|$B� �>�&=�l >D�=Q�i�p9�=�|L=��=gG>��g�VI�G�۾Z�>����撾����n?�H���+["���>n�?��D�����hY2�ˌ@��>e}�>֔n>���="�>鐤��SP�I���m>����z�/��>ͤ<>R�d��v�=st������&��/�ͽ6��6;�=���=c�4?�~V?*�>p����+�R�S��,2���@����=z�%>��7���8>�Z<�C��g侐��Y�>��C��VM���w/>�a;,"۽M�d>q4�<��ƻ\�_>�U�>�����hG�=tN�>PԶ>@�?��3>V(6>�V�⃿��ڿ�����۾�+����:'�Ľ=3}��S�>�#��AJ�D�&�qYp>J< ��i�>��>Jr�=��=�sV>�|>0ܾ�7���g�Eо��m��M��/B�3D�>r��م$����<\=���/�� ���"ܽ����������4��#?O�>�ï<��?��7?"S??�;`��9�>�
�>�p�>�͉����>�p0��?��?G�0?�ߧ>�,
��[�Y���(Q��s=�:>.�->�~F>�d�=�9(=K8�=��ؼ�ʺ}�(���t�����.>x�P>��N>"8]���%�R#��3����վF��<Q#?�IѾ�Yž���E=L�1�"���Z2���{����{姽��>5��>�*�>�=��>I#��d�[�>����e���J=$J+>@�=)����N��L�=쉾DO��kѾ]H��!X=~f�>*Kl?�T?�?rU���DK��bn�5C�&վQ�>o�>9�A=:ҽ=��H?����8��6��}�6�)�MI�>�=�+��-�K>��	?d�>���=��=:�0>Ԫ!�̳%�]I޽�>k��>��??6�>� �>1N�S�>�ʿ΅���!���A��:w��_�:eK�s��t	\�p/���������<���=��R>�aO=T��>X>c�>�P�>dK������罙������+�7�c���Q�/�xZ���R��9W��_�=Ƅ�p�'��9K����G赽��ƽŞ:����>&�4>��">3�?^"?��+?=�?�@��q�>�>�C�>V���4�>�<>�?��>)M?��>^7�<�V�����yW�=%F��\��=�M>y�>��=O3�<Ɩ�;mˆ=Eu<?�;�:b=�H��i�t=��>�7>�s�>- �={��)*5�
4��;����Hu0=�%?=䞾���5>���ҍ=�J��W����/�� +��- ��k>�w�>\ġ>�'>�d<��t>?��f�)=.E>~YT�
�J<��>
��>S�s=$��;�D1���e���J�!�>_��>��>y&>K�C?��1?Ƒ'?7����.�X{K�' %��-���u6=�<�>J9}>6�~>��T��w��մ�������x�����,{>�Iػ;;����>,��D����==�ֽ��Z�(l>t
�=1V�>3�?��?<��>Z��=�0�����iNʿ�h���������=`�=@��WC�=@�>�4�;�"�N�̾����������=J�>3'G���r��r�=���c��>�F��m4-�8�־]n5���=�E[=<WϾ�����Q�<�g��?Ѷ��!:�����۾bϾ锦�:�?���>Tuj>��>i�?m�+?�t�>7�F���>�	�>I٬>�З<��>��?y?*,?O�@?��u>]V����=]���jƽ���=q��=!.s>X��>��:��:�;�=���	�&�s��H7��0?��x�=qd8>��S>�?�\`>m�M�$��X��NtҾ)kٽt?t�X`c�RȾt.?��(Yھ�Z	����h���=_�=)�>���>�J���=!�־A�{���޽���m�>��>��K�Q�<:>i��M�쾪����c�Fٌ>@h�>2-�>�?0?��D?��1??����*�Dk%�k�־�ܾ��.�%B�>^�b>}�S�'�P�4T��Q;�i�)f>�BB�^t���\E�ww�=4��5*i>��+>j�ۼ���>u��=v�Q�?<����7����>��>��o>d�>p9l��E���Q̿k���\��b�𿂾,��=ߞ���H�oeL>��<�L��gh���H��'8J>��>�iZ>M��=i/Y��>������;Nゼ{I��A�"`轳�D�� $<v�d�
ܚ�������b��a)���ս4�ڽ�������]����2�`��>��=!����>��P?��1?v�&?*=�<nx>��(>Oǁ>�X����>g�>/[>#k?�>,?��?^�_>��ѽ�=���`�>��>��=�X>C���>q����^-�<��K=m�G=��=�>��>ݧ��h�y<G��=��?>��p.�����,��8l>��< �M?.�����=4��R�=��+�:�����f��I6�^��>{5�>�|i>!^^>
�;73��*0�,=�VD<"�J�>s�Hh�>��i��o������k�����|O�r�4>z�E>�$�>w�Z?8�K?c��>�mI���f���Y�p��T���\g�<b��>�C�>���>ՠ�}���E!���@��2�0D���Z��/	>�����W<��>N��<��}�<Ͽ�=����5�<�WL>TJ?>�ħ>�W�>�z�>�2o>)�b�����QͿQr������D��E��=D|߽���;V�f���2�{�����W.���ߒ=��>(�`>@�>
�>��V=��K=�<����;����~Gv�&Z;�[f�'У�~�"=�����ͱ=Gћ�Bq=�����t����ݽ���H*.��+�菴>�p�>���>��M>) <?">?��*?�\��9Y(?X��;�fq>��i�����,{?�:?�Z?�F&?�A>{��g��`>���v>�}�>11>ѻ	=�f>���T=�P�2�=\#�b���e�=���=����(�=�>�4> ��>�8S��|	��$��������< s�ML>�u�(!N�O����NP�3�پw��o��>��>���>��>`������<ݳ!�5�+�?��>��=���<S�==��>HIὉެ=r4t=�SL����P牽�L�=�
>JV�=q@1?+U�>Ap?�D��i�%/'����<���E��6�>�9�=�1>h���0 ɾ�!�u#�M���0�Gl�4l/>`+�=ƾ���d�>	@	>�X�������=��"���ν��6>�t�=AG>��$?�#�>M��=������1[Ͽ�L��(��Y�����T=��A<F��{2>0,�
�?���7>��/��%��O�M=���<�&=�F�=_\��.ly��%>����X˾qb!�3,�QJ�������=��5��I�=�8��9�F���v�nĽ��a�����=��e�>�_>�[�>Fb�>�O?�g?��;?����>�:#=@{>>�A=d�	?�E'?�Q?u�9?Ǩ*?ƨ��<`��D�+�&d�ʃ�=�AJ>&>;_�;(�_=5���U��͸���>[�����3<0�"��ȉ�/��\{�=�U�=���=ħ?Pd&��?����*��0�ü�Ǹ���?ؑ���f��g�E�>!�#�{i�������k]=4��>��>��>i�>U������;>�s��~��=c�=�R{�䥱=ƨ8=�nʽ:v���Ͻ� 0����<͉�=�c> �=`�Z>� 8?:��>�?�>��,<φA��4����y��-O���@>ŧ'>��=�Ӄ���wE�7<��uʾb�!>4���nЏ����=M��=�����==!/�<@K>,z�<R=4�.>�g�>q��>,?�$,>�.�:}������Ͽ�����.�x���+��==�º|�˽��� -����_�,���b���޼Tv��Ƃ��7#�Z2#�%�=��>�}<������щ�5]���&���꾶��=�l$�\���N���v���n9���ʋ�����2���<=�n��ń^>�u>���>��>��>H�>|$?�$����?k�>L�>�A�TJ?�#.?1�N?�e?=�>5�3=0�����'��V�Q=��Y>�~�=Ġ0=���=�E��I;`�{��{>�W�<�o=:u��
G���N���T=���=R�?>lo?xeT��,��9�T�"�1>>�����F>�@�;���>��]�wgh��*���w��)���-��-$��}�>�|?Rm2>�7Z>U�'��C�=""Z<����`>g��=_��<b�U=�(>`�,@��=�F=��ƾpȽ�/��k!>Od>4J>�v)?�8>�E�>oX)>^�Q��~�B�4� ej��T�*��>*T�>��>�c�������!��j�_2ƽ؋��6z= [�=$]V=
B>�##=v�
�Ҡ�=$[μxO�5��%3=uj>��=��$?�֫>�8=<����Ⱦ5�ӿޝ�������*S>��h�Z�B�O���"o�=�܊;�M����ӽ9�����4����<��?��n��		�> ��Q�����g"���3=�`�Q ��
'>�Ʊ=ǚ�"��=�̜��m�=�j5�aEx=]�0�1��2F⽲;�=ް�>�1?�>�T�>�y�>F�/?�%����p<^���w+>�z���;>�?F�2?=��>}�>Z���������W�,�`>7'>��b=�q[=f�>@�Z���ｧ��;�=�(�<}hǼ\4��!�6e(��I�=M2'>��>J�?�#�=x����S���N��C�=�(����>�ka=�f}=Μ����R;�ᕾ18���Ⱦ��G��Y����=�R>x�z>�E>6@�������pf�="
1=�K�j�[�mu>r��=pQC�$���;��<�˾|�5	�=*v�>X�>�� >F	?�*?�-?S����K$��=���OE����I����l�>���=������|��є.�3L�����:��-��-���0M>e�=ɛ>��=��j�|>�S��I�� �8>�F�>�s>*� ?���>Z�>�Ӿ�%����п���c����i�0�T>��q��D~�ʭC=U��=]����.|�3/@=L���G�=��>���>B	f>-)�:��>����]k�=Q�$0�� ��M;k�����d��=k&�<����'%��%����L��eV�g����}�_�����`��$�`"�>��>3sx>1*6>�?zJ?7�?��NvK>� �>X�g>���3|�>��?9�>t��>}<?�Lr>~b��52*���s���;>��>B��=�V�~��>2S ��&>�$���=�>�n�>zcl�� $>�F��>�=���=��d>K��>*6%��#&�꘳�� ���bN�D=A<�%�>0�ʾ]�s>YD���9�W1h�Ī���o����$<�>� ?z^�>�+�>�g->aS�����=������m#`=!�>Ӛ�={=�=q�J>v�.>2�=��@�.v��z_�`���S��>�� >��>7�.?-i�>�6�>�}��J)�^2�u�7�b>��潲��>^��=	�	�l	+�B��³�������/ݾ���~�����=IQ>���y>��!>�4�ꭞ<��ǻGc׾Q�x<c��#>L��>Ϛ�>��>#��=�\������nܿc���a���q�=D�q<�4H>�\�<n��abw�<�5�t�>�Ձ��ō�WrC>��+��0��c�~�;6�^��k��-��.��ً����_��	(����������v�����彵Ц�}H�� ���
�]P�o���WpL�fH�>�5�>�c�>3𙽍��>@��>a��>ZY�(�>���م�>���>w�?n`�>��P?xn
?os�=�;�h��տ���e;��a�>�Z>)��=����}�=���sm�=��>�H��B�� ��;V�C=�2�Bn(<Pn�=q�E={F.>�!�>4�B<����M�W���q��'�̾O�>xF
�'��=մ���¾�}���`�=�о���sT�>5?�[l>Udn>E�> �lY˽�@��gt�oL�:�.>e�>-�+=��&>�����=S��]��7�W�;��>M;=H�>vaB?�d�>*R>)�ҾHc�����x,����;��S=�H�>X��|��9���4оR�o�ə2������v½�R�=�v;�i��e�>�Ĩ>eP���H��=���^�R�a���+>��>�=�{�>��@>qR�"w�D �s@�O@��}_���p�ϹP>�����> �=~~��K��G󿾯|»:f��_k�>&�i>�U�=�޽�1����n�;1���H���<�@�����Ⱦ��{��9=����|���y3��F��-��� 9�\&�vVU���	�W�����G�D��>�W�>D�
?��>�r�>B�?2�>TgA�k�:?�=G]�<z��>��?a�>��?��>�+�� u+=�Ad�� Ƚ�Tu�)> �>+�=Q�9=��>=bP�=(��=�FK�{���F��T�1>�o
>�_=��=�!5>�E>��d>�Tо�^�3<��ѵ�A,j��{����>F
���>������վ�;������i�ۨ�>�o�>�e�=�j�>q\>�6���kѽ\{��4
�	����L>���=��>��1>"B >yr>Z6�=1����;��R�B>(9>4�q>�p8?�r�>��?�� �q'D����Q���c潧s�>��Y>'�>�*�=^!�<T����`M���N���K�o
>�ٺ<upZ���>�={0޽�o����O���!�V`�=��=�vn>�l>Ld�>5D>̕)>P���f��̷��t���������={�=Kg�<y�1��ѣ�����g���ľ2(��(���50��=\�h�dս��������+_���܀��3=�����Ū�M�9�����-����Ǿ�a��Nj��>��������is�E��������3>(�>@��>�N�;�v�>-0?8��>$���$?�<���x>�I�>���>���>�?`��>ؖO��;��=K��YE�U{�>=Y�='\=JG�=���=�ཛ6>��.=�Rƽ��X��~&��Z�����=*��<<M>=f�=�D�=�nc>�����-/�料?m��ên��ԅ>ˬ�=gg���>:t�=�����5���2_�q���$3�Tb>�r?=�>ڟ�>�ݘ>$���E�b=�|��OL�p��u�9>���>�n�>�aD>�2��
�=I��`��& e��(���{Q>�>�D=> $?�9�>�:E?1չ������!c����=AB�<O�>I����Ͻ���_�x��[�*!�I���|���@�ǄǼ֡d>��)��>��=��4�]J�=do�=&��E(=/�=�t>J5�>�>fL>P�,<����y�dpſ򗈿��<�k���]�>�8��uf�҃�;Ut�o��gң�>T=C��5�	>�J>��>���P���k꽥��$�V�:�s��:��;���	3����L�y<�����&���x"�mM����Y�'��B+� d�^��Po�[�'�++�>���><�>l��9ϻ>�d&?��U>8>��?�������>?�?߰�>�C?�p�>�+}>�+A��̾�d����9�g��>��f>�9>�=�Ç>��U��۩�hq�=��G��/�=�༣�Z�}j=�b*>���=yC?>�>K��>*6%��#&�꘳�� ���bN�D=A<�%�>0�ʾ]�s>YD���9�W1h�Ī���o����$<�>� ?z^�>�+�>�g->aS�����=������m#`=!�>Ӛ�={=�=q�J>v�.>2�=��@�.v��z_�`���S��>�� >��>7�.?-i�>�6�>�}��J)�^2�u�7�b>��潲��>^��=	�	�l	+�B��³�������/ݾ���~�����=IQ>���y>��!>�4�ꭞ<��ǻGc׾Q�x<c��#>L��>Ϛ�>��>#��=�\������nܿc���a���q�=D�q<�4H>�\�<n��abw�<�5�t�>�Ձ��ō�WrC>��+��0��c�~�;6�^��k��-��.��ً����_��	(����������v�����彵Ц�}H�� ���
�]P�o���WpL�fH�>�5�>�c�>3𙽍��>@��>a��>ZY�(�>���م�>���>w�?n`�>��P?xn
?os�=�;�h��տ���e;��a�>�Z>)��=����}�=���sm�=��>�H��B�� ��;V�C=�2�Bn(<Pn�=q�E={F.>/��>��˾*Ϳ�����f���V��=O�>��H>�<�����!b���8�oN=,��>2��=���<kѽ��=��<=���>�=��Z�<�Ƽ�8>W˅>C���IT�y>�iP�{}4�6�@�Ț�=�>� o>w��<Uĭ����~ؽ��=�?h9�?y�_?�m�����&;�I3�`Z ���o�3�ƽ�۽W���e۾d��C�־ �ʾ@ľ�$$���1�A>���=��=��=>ھ<Y��� �f=�j6�,�=�g>&?�;�=�W�(��=o��<d�+�j+s��]�=v<�JB��-%�b�޾�e��\�p�AŽ#�]�u>��A>��0�ھ��(����<㲃��!=��=�F�>T>;m���Y�%�x���Ⱦr~��>��f a���=��W�1*�=|�m�
|7��/@�o|����&���ʽ�t��t�a��j<���>@u�>w������`(?�Q>��>�W�>���>��)�7�>:%�>�!d=���<=��> h>i��>��+����{�K��>"�4>��,�����O>���I�=��=:�=��>�A��e���Lk�đj�wg>�l�>Eҗ=0��>6������%���O(���>[F;�0=b�Z�����)������Mj�=f��=�iϻ֯�4]>8��>��>�%�>�U�={���t��=�z"=^u�=�	G�%3k���=x�"�y�M����<�%=Ba6=�4>���=oNO=��=�N|��9ҽ��?`3C?��\?�w�=�Gľ^¾�	���:�g��=�E�x4~=��C��5�_�վ��оB$��,�p�⽋_�J*B>&`>n��=��5>��=ŕs���=���e�rӃ>h5�<�kq>��O=lb�=�V��+1��~�[6d��Kڿ�D_�� V�*g1������3���=�1P>���>�=>��W�)Vx=��ߺ	X�>1�=(��=g+`�o�̽�:E��ƽ!�3�	����������#QQ��_�>Hi�`�=�u����v���x�J�VJǽ�P����K�T��v�B�wߋ>���>���=6�=g�>r�<>�$>9>Gm+?�F�>O�>J�=�  ����=��>Z��>�:j>/G��D����#��
�&\>�=I���吸=��*>&)=���=�'�>��=�����a�ҽh/��m��X�&>S�>v��=@M�>pP쾷X�S�ž&�d�_�+�55 <S�%���B�ln�6�����ڔ�b�>��H=���<��=�ko>���=�}�>_|<=e�"��_h>	O>c�>a&�<^�ǽ��۽*�2�oJ����=9�5�m��=�h��P�N��=���=|L�=�?��M?�p3?�˝=Sq��H6����������>iD�=蹇=�?��B���z쮾�1Ծ��ξ'z��_��=��K��F>l�>�\<m�+=eP��a�2�;vܽ{sA>��k����>�=7JJ>���=��o>���=*��0r���Li��dܿۆ��Ӣ��;�l�����&��X�#=:[
�% �=g�E���j��߽ކ;>� ���[�=����̡�;e�c�*2O�����E���ǔ���� �:��+>����Q�B>�4��IE
�'�{����Y�	�>��<����F:�6X�௝>��?��/>�
�>�1�>:F�>���>��>�?%�j�?j�>��=|�����M>��->��O>N�ѽ3N'� 3�2�v:>=?��;{�����=>xr_=	B�=����9>���<Waٺ�Eн�~/��rP�oܓ���>\�K>H�=�?�iǾ��ľA���N�Ľ"�>[s>�[>�U��Q��g�Z�>,M>�W�<� ��7<�>�,>���5>&��=�	�3��	�<�K�� ���>-R�79<�I��	ԋ=�=\l��b�8�8���~;ݶ2;�ج�EU�=�^H?V�G?¿L?�$�����tҾ�?�������4�<��>ژ<uIٽR.T�3|$�3�@�z���뾨���67/�G>�>=W�=�L[>��Y>BZd=GW������e�=n^�7�!>,�a=�Y�>���=5�>�Ӊ������(S�;��Ͽh�^�($��cjԾ�i�������D��r��Hʃ>~�>�=��?�����B齰rg�D2꽓yདྷ�6>8|>�g��䧾e�E:X��|����`�A����d�'Ä�0<8<�K$�8��U};�C��r�����<ڽk�K��U=��J>9�"?s�R>�dp>�n�>e��>.�=7��2�->�$�b�>>�ҽVvr=��n>J�>��M>d��=���Pl'>Q��HI����=6]%>�0�BV
>��>P�-�A�F>)͐=���=��,�s*�3���EL��cć�:��=�m=���<$$�>������_��@���t�=�D=�_g>�������ɛ�H.R�� d����=��=t��=.��=���>N��>���>�a�=�qx�/ B;��d=z_6>H�=���=�Q!=�ͽ0�����=�)�= �=MS>���=�\�=\�=!槽B-��p&?�d?�Ia?�V\���ľ틖�8����b�]\J>B��=.�=��p�
����dԾ^�پ�A;�$��YXZ����Y>�o>��1>A�=������W��@9��=�b���P>���ez5>� �=Fʭ=��&<�	5�hɄ�0�c���ܿ��|��2��a���Q�P���>���g��18��Ҿ-ޏ=(Ge;��6>��w��E輨!�.9ݼm_�=�������!S������������4�R����o��� >�<���!��_	������zi�~��]���dxL���=6��>z��>�,4=��=n�?'�>��<+�=>{?9���~b�>���=6��=8v;��>�+>�Lm>$���v��k¨��3>[�<�ݏ=����=z-�=X�W=�J>���=n��:Ⱥ��ܽ��J��W����8>�:>ˣ4>�=?�����VξRL%�r���.�>v�%>������+>-������
�����>
@�>A7�>�4>�_>�w��T�b>�k�>��1���D�Fy�=��1>��0>oh��� "� �:=�<�<�9��m��u\��C<��=kq�>��=��<�k'?*j>?ri�>:7�=�>þ��8)
�}s�=�!V=�</>�*�=1�<�9�����ݾ؍ھ�ؾ\��;q��Ez>�IO>�,��� �<n�ؽ�0M��B�=3�>{��=࠳=*��=�>6Y>N&#>�
�<m���U���Oc����AVr��7�_���[1��ھv���紾�ҕ�ؗ�<u��!�����{!��U�I�Q�B�����ھ���;/�d���f�zAB�%0�W��.���%>�墾�R�1���}����}}B=��#���E��gd��*u��}��@l�<�?�ڔ>/�j>
�3?{��>�׻�Ia<�o�>U5{��P�>�d�>��=�Խ)�5=M=dd)>8�C>60>>�g��mc[�L�->�:>C��=}��Oֽ��Խ�w��a��= =�Ԟ;F/����o=Þ}=�9
>�-I����Ǌ?xt ����G�q���?�=`��>UB>�I��^1�j�����<���=�M�>.�h��o>�n�>�}�;d��>Yfs>���N��	=�OB>�⨽�	�񡓽H}`�f-���}=@�n>�,y=��=`�A<
�/>�->�n<�׉o>��!?j$A?��?[R*���׾U�1��߾*��=V��NS�=���=^�H:���������վ�<{�k����=�?���}�=�Z�=�l> �<ΌϽ�*l��p>�=}�M>���>����2���=M�=E�
>¦;[K��S�<!=��膿.�¾��e�J>���ā�j�B��J��j!>-��1G�7A��bX�)����z�<���"�A���=^@O�镞�S��Xï��뾾�L��~�ĭu�BK��2i�=�_��H��*Խw.s�����q���T�p��?<�55>�?ΑZ>l�X>�R�>�H�>QnG>4yC>�2�>R̢<c��>9�&����7
K���>��>���=�Q�п�S������l&�>���3�!>�h=�ؽ=�fڼX�>9����4�<
�=�4����
�=�[���Pj>��+��=�(?���X���#�eAc��z�>
��>��>Z
>�լ�׍�2Ӱ��Ά=}f>Hj*>媽޻;5	Z>�Cd>�7>��d>�u�]=Xx����=�Oy<�(�=l��=���{g�=I�H�$��=D�<�(a<�i��?�j�(Z�<:���=�0?U��>�S6?���D��aŵ�ޣ4������M�>�`
>�->��;�M,ɾ���� Q��7~��g���̮�4��>�J}>J��=mo>~���$&��h�6������%��=R�;>)�=>sN>Jy[>p��9����>���=U̿����K3�B����ξ�X�w��.˾�?����??�k�,�B�LF��1'��Z᫾�C>X^���T��V�꽫0��$㭾�ᨽ
��Ҥ�a�3�aļ���<��ۼpA>8:�)�������ü;�e�Y���w7O�ld��x=ŵ�=�>(?�%? �>s0$?FG�>�v��W�½@�2>������)>�"�=��7=�K�U�>�RG>�?�>tƗ=��ּ�"潹(T�f�i>�V�\�="��=�x:=���<&�|�>v�ruR����!�e �<7%�=�Hq>�"o:��=�s?�އ�;W���N	��Ӿ��<��G=��=��%��Jս2޴���f���=VjE>s�m���.�@�>Mn�>7`ؽ��> vM>����i���J0<���>�UȽ�=��=5�D���a���Y>)�=N�D=}�r=���>Ｆ�=��B)���>�L?+-?�D?*�8��ז�Y���ਾ�>#���<�F�=�{=�~+>q�����ؽ'��A����7�5��E��>#��>tX�=Њ�>�+=����=5�&;|��<)�>�]ܽ��=��=�*3>�Lx>��o�_�f�iO>��׿�_��HC��_u=��y��H��q�>@�� �v��>��R��8w�l줼'�����s�>s�(�,�=�`�>��!��݆�%��T������۾�V��:�O��~�&�>p��N!�u����_�F{a��p��$X��X2ӽ�S����0>~�!?��>4b>�M.?���>��k;8��>@ޑ>Ц���>��>p� �GW�?�=�����νU=M3�"�	�Q�0>��=t����4���>�z�����P��=2�8=�[��C?C�&ú��Cż�2�<�>��>D��=��?N�پ/������N߾�/�$�>�ub����؈�>��|�%m̾F�O�m��>��>�	
>�>�6��>�$�>d>�>%��<�I$�`��2 v�-�>0M$>�M>��ܽ����=��B��^�:Zu>�Vl=T�~=ܠ5>�r���Z�� >��&?(j
?�J�>�ZL�֮*����������z� C���4>S�=ϻV�͉V�軾M���r���Β��se��9����=>Sw>�Ѐ=�]4>|蜾�5߽��j='�>Z������1>>p��=��-�)��W;ӽ)Nj�m �=�\ݽ����)�|�rņ��ۇ����h�n=��ʽ�+��+)�<Y�<�پ���UT	>,[=6��<����B���Y	��OW>���<��=%��<�Z�b���ɾ
�[�Х���.�^�.>�9[��� �&T]��y*��Z��i���v��+�,�3T�'3Q��1?Um�>�h�>tC6?���>�Ս>�o�>��;?�o�l�>�c?�+)���R���=�@�=0�?��Ƚr��0]2��\��\I>�=��>�b
>.Z�?ܽl��>�->���<kb��&|������#S<ק=D�<s��=F>@�?lD~>Y33���g���=���>�]�M�-?�O����>��J�8�>�� -���ľ��;���c�hG>���>l�M>^�n<��C<p����ʽ�6>N��3��<o�7��>8R�=�n�=fM��d����ed�ʌ��y�=�X>
�>��&?ڼ"?&?��0�i^7��+�e�J�C�>��]�d_�>b�>*5U>s}���+D�	�(��Q����8��jݽ�CB>�S_>�>��/>F�T<�l����Z+H=d��=)�=u��=�`�=�l�>���>y�x>���>]R��Q���ҿ����)�U� ��Ț�����pN�g3��M�륣�w款N�����W�>�b�>���>i$�=�-M>�/&>�K�o�使��#\�b�^�����i̒�~&>�Y-۽b>>���:�f���^��r¼���Y�㽦;/��‾%��
��>O�A>5	?F?f??��>NVC?)O>�9�=g��=��?�s�N�5>sx�>��? �?
�N?�?�F'�^���^�q�ӽ=���=�E�=�y�= =�=�z�;RY�|L����s�νh����mg<7�O=^
�=�>>��>�'�>D+>�#?�U<y�'F���Z%>,:�v�-?����^D>GP+�/彯��/7,��������C����������J�>z�T>K�6>H��=!Ⱦ����j~>Cr8��q������.�>(�n��>�=�U��.���ȼ��쑾�f;��>> >;�?Ş1?_Z�>7���~c�^M�9+D���������>�*=�� ���?����2�*��o<��+�ut�=��K>��>�m>4%��n���	�=�V�>��%>��=y��>�~m>���>�X�>>�">tҥ>����O��q#�[�ſ���Z�پ�=�=��=�n�;���F�q.>:��h���%���>�͖>e!�=�GR>Y�<>%�<:GF�7�ؽ����������������)���>�f0��&D>r]	�ԈV=��j��g���i½�7^�/��j�ھGȀ�*��>M�->���>U?)�?��>�$?�Y�=NV9?&U>��>��c>��?�	?e�	?��>�k*?��?�d����&�OA�j�ݽ�q�;��$>��>���=����\7=�݈��6�����Ze���T��;s#=`��=.FI>��>5��>���>l+�Ƌ[��Fy���>;M�I�?B���_�>ȏ/�G:⼃eվG �oiC� b�Ձ�Ƽ��[�9���>�9�>������8�����n��5V.>f	���ǖ< �3���T>��5U`�Z��v��a���-����އ>�X�>q<�>���>Y
_?�t?���5.�K|پ�1�ю>�Xо�N�>���>��J�gc
����̾Cs������
$�QE�G�p=>F0>T�=��W��ͧ�=F�<!�=���=l�=*$�<Иg>k�>��?r%�>]֌>q����O���bڿ����� /�r*޾�^z>ktC;�!��a� �Hb��� p>����R���ϕ*>'��>���>�k~>}�4>�M�=��4>c򮽦qǼ��k���cPu�(���L̪�_��=��3��ѯ������c�=�Pj=�{m���A����/c�����n��>��=R�=���>���>4�>pvB?ڀ>X��>�ɴ��A�>�=��>rH,?���>��>��-?M�'?|$>%뭽+Ǆ����<7�=�gJ>�=��>ga���1�<�'�=8����<B�̽Q���g��ә<�ю�} s=�>���>X�A�[�0�1���ܼ��;�< w�=!I?8����u&���k0^���Խ�$+���2��E�|��>��=/q���=�B�>R˷�
�ͽX,�=�s�A�=7h<�D%7>��==�=h�-�L�s�ּ�=���'�=�}
>v[[>"�?�{'?nM!?�|꾵Z*��B�<�e�p�I>���P�>S��=�g=��0>�Kپ�Ͼ]����،��䔾�9����Z>җ�:C۽��z>��;��e�t�=H2���
>�:>q���A1>���>���>u��;X��>Қ�T���ǿ������Q��7�����>�){>��I����<"���o�=�8��:jw�.F|�D>�)>�a�<�|=[ˈ���ݽ���>t��=D<1�K���_�<-	��f�����=���p>����x�mx=��j�1(��X�Uқ�̭�����rK>�>�:?��?���>��Y>#�?L�S��??�'>Ot?�>�H�>M{�>}�6?�d#?lXK?�}�>އ�ѝK�|�T���g=��f��>?;>�X'>��=��3=o����:=�=>w���*���I;�]<냛<4Z�=���=D?��>�O(��S�3`k�9SX>�Vh���>�r���>"0�!jؾM$�!��/o�		�N��i�W��<`��>��=u�(>��>�jO�PQȽ+=�o���U�i҉�3F�>��=鳙�rGQ��JS���z=�zD�;�>:>�{>��+?��6?8�(?�l���B�З��`O���4�CÃ�~9?yR�>��v>�l>n���9ľ���0��4��F��Gl[>}�'>1��<��Y>�+=��<*'3�g�)>�cc�x��<�5*>�;^>�؈>��>�*>�>��=���X��3���$�"�*�ɾd���T����˽l��=G��Rپt���	�ݽ&�;>�s���C>2�>xe�>�iW>��>�L����ƼCZb�����#B������=����g=�s`�J\<�:��~�g�ʢ(� ����vL�o�=����h��Ss}���>�A�=w5�>j��>�F?]	�>qy
?�<h=-�?q�)>k��>���=^�e>�h�>�r??U�>�9 ?� ?F���J����#���\��l��3��=9Lh=x�=l4=��*=!-=�b���7Q��.�:%�<<�27���r����=�X>��>7n?�+����/�[+��˾��T>��=*�?;��4ތ>ff�o�*��cJ�O7��I���̾�k>�>�a�>�r>���3P�����Z>�����½�%x�l��==�>>�^� �a���׽�e�
��k~�=\�6TN>@�L>�v9?mG�>�%?�eι �! ?� ��|�7�����:;��v�J[�=�恾J!v=���EQ�^(��M���k��z>���<fH8�E>f�P=���^Y�=��>�o�iuͽ�+�=� �>�܍>X�> �W>\�������d�'=�ڟ��Ej�#Ա���N�*��:�=���>��;���O=�n>LAE�����^s������{�C�e�#>��;Y;�
�*�&2I�e����7��ي�������=�d��s��H�$�p�C���;8� ��W�ͽ̼,�Od�<J�4����>"�?���>���>1�?:)�=Z�P>L�پg�?��>���K��>}.�>H��>�� ?��	?a?�==wn>v��q��z>�>>kW=>[����Y.>��M�g�>�s�=&I����=:׷;7s!=�h=�=�$�<u�=��<�?󠭾+MR��C��Z5��Ӄ>�E��5jG?��6���rz=�X����3=)������XоT��V�>tG�=Ai�>0�>l!��q� ��Bu=�A3>�e>���2D���)���Q�.=.=����<����?���3��=�Z%��)>2^l>�L?m7?d?)2Z�ե��2`/��.��C�'GX�,E;>�Ɨ���R>C��w.�<�g����c�|v%�	��l>�n=�ħ=8\P>F���t�v���=��n>٦�=��N>�_>���>m��=)e]>:��>�F(<��μy�ཅ�ؿ����g��������y�%^=e>Q�2=����=͗J�=�K�=�{��-�>i+սB�<���<��P�<4E��ž�~=>崏=�Y
�1����!����=L���\+��N�clx��,�@��������;aʹ�8=��2�}�#>���>�e�>��>=X?��ս{�>����o?�N>d�6�F�?�9���>�V?&�>t��>Mʐ>�*�>"�� O��/'>��<�Y�=�#�<Ȑ�=�����<P��=��<�d�<�V��f$>r��<�Ǽ_a����B���<'�?�cվF�?�٠!�����]����>= /?�žTC��F�>>�۽إ,���9��L������� >?�>ػ�>$�L>[@�������t��^C��a���V�M>��>�����y�=K����y:��$.�{_]�q��=3�����>��f>�#$?��+?4�4?����������)��^���I���;9>���4Hf>�T�+��n�����'��Q辏�N��]b>xb=�����>(�ѽ���m��=0`9>E[��׃=�C�=�]�>{#>�R*>��>�h�=e��Z���޿�u��&�����$�NZ��]�7�;>9�O=�˾]�<+�K���t��\ǽ�f�>�>�J=ڹ��N!a>B�A����>�/�|����0>c����)��d���q�Drv�p�n��`����{�&��	��L6�x�	���\�����R����=u�?댷>�Է=Xg3?�#>�ɡ>�늾@�1?��>Bҫ����>��<>j\?s��>��>S�`>b�>�vԾ}�����>�:>�˺<g�1>��>�|=O�W�l�S�#��=$��z�����e=B�
>�3�=3�.�%�/=y�'�?�cվF�?�٠!�����]����>= /?�žTC��F�>>�۽إ,���9��L������� >?�>ػ�>$�L>[@�������t��^C��a���V�M>��>�����y�=K����y:��$.�{_]�q��=3�����>��f>�#$?��+?4�4?����������)��^���I���;9>���4Hf>�T�+��n�����'��Q辏�N��]b>xb=�����>(�ѽ���m��=0`9>E[��׃=�C�=�]�>{#>�R*>��>�h�=e��Z���޿�u��&�����$�NZ��]�7�;>9�O=�˾]�<+�K���t��\ǽ�f�>�>�J=ڹ��N!a>B�A����>�/�|����0>c����)��d���q�Drv�p�n��`����{�&��	��L6�x�	���\�����R����=u�?댷>�Է=Xg3?�#>�ɡ>�늾@�1?��>Bҫ����>��<>j\?s��>��>S�`>b�>�vԾ}�����>�:>�˺<g�1>��>�|=O�W�l�S�#��=$��z�����e=B�
>�3�=3�.�%�/=y�/T?��w�R�XK7��1ž;=>��t<Q`?�̾���=�+�>߻��h=���ƾ��Ծ@��=>��~>��1���1>V�>R'��H�H�����<�q�:�޽L�2>�>�&c� ��<ov���νl�����CN>�-�<�0�>���==Z1?a?�n<?�)��t��	���|��z��O >:��킊>Q(��AX����'��n#��n��S��h�ҽ�0=>B�4>�\\>9.4���u{>~�e>�н<!͎���=�O�>)>��h>�Kf>�F�=�䜼�W#��:ۿ������y�٥��˗Z������!���>4R���b��FC�����&A���:>���=U��<�(�<�>����nQ�=}�Ѿ������=;♾�U����J�R��������g�J|���9��&p|���ۼ��[���[�g+�(�q�{�ɾ�#>���>�F?�B�>�?��)>�ѽ>�䓾��$?s|i>����Ч>�6�=�?�?Wt�>�J�>�2=E��>SjJ���4�9Q�>��>������=�_9>��;�n�8���x9=�5�GS��O7.�LÑ=�	����En���=�#?�m�u��+��z$���:>��̽N��>�
ϼ��=�Z��лB�I'h��\�h�����=D3>���>�˙>�I�=ν	>�1���ۼ:��ʽ�
>������=*񔽥8Q=C�$=��q����=�ռ����������67��t&�<�:->[�;?��?�V?3��������W�֦���y�x6��\�>M�>�N�<�/�s����߾�5���������y3���'>2�?>┆>.��>��t��姼@ߨ�b;>���w�e>��,=���z��=��~>jq�=� >E����I�Ϳ�*���ܽh��U�<_2���&��˾��/�|��<��N�	r3�!z'��YQ>W��=��=W�ڽP�ེ�<�6�>BN�N�<����r�(�i�����a\;>)J�:ŷ��#��P��=;�3�� �P4��䚩���j����k8��x:>Vi�>e`?K��>�?��y>��>d�*�d�W>�=-r�>�.>��>�d�>`v>��=��>�9<K;�V�1��h6���`>�@=�7<Vs�=�f>N��K�=~>���;xw���{к䓾=1�����=N�Y=K��=v6�=�?��-�	���]�>�X�$}�=�5��&˘>~T�=�U=x���v���ȾE~l�Rc�<ɢ>�8H>V�>9S�=D��>�V>$�������{=%�q>����h�=N !=�s�=�+�=��W=%��<(d���k+���CK<B>=�bW=��> 8?���>_	&?>`;��������˾�t���Ľ�Fڼ�ԉ>p�>�T�<�����ϾCh�e�=C̾�/m�|�;D��>�!]>�t��������7���M�w��I�`�_����'=�>�<>@ԓ>�]w>�a�=ْ<�W;���޿�����,=I�L��~�=g��������g��/�н5��<����6%����>K�P��1����߽[~=�$>��+���h���Խe^o����m��ͽ��d=٨(��3��)�-��.m��g����b��[����
]M��/��-��;-�=���>h��>�j?���>�.,>���>Gax��1>��=K&s>C�e>�	�>�~�=�$
>�8�L�>!�}=Z��=��㽴�#��H>��@���<>���=�>�(�<g=�=���=�[�ę�9��<R���#�J�=���;y�z<�J����?����5P�?s�-l����=�Tν���>�4�=��%�]
�����r�h� �a��q⽥K>�,r��/�>E�>�+�>�">�.^=��=9kz>xP�S�&>gn���!>�7=��<�G��~�Q�%=���*=��v=bл;�2>��!??�>?�#?&HC�|���v�ȾX�̾6�T�����6>/GD>��C<L���D��F����s���ƾe��� �v��C9�>��>K�E=�u���b|<V;)���<&�i���8>�怽�8>B��>�]j>�"D>��=d2�Z�[�R��}���q��M���־�Ȭ��l������
�����>���{�!��5���}>��><�B<�kI�8��	�ɽ����=����U�
>���ʤ�I��X
��Tdv�w�Խ�y1��+"�pH���)���Z�
eI�����M(��5Ð��꯽�ex=V��>~�
?H�.?�'?=>I�>��A�`�=IѾ=���>��7�ZT�>�?�=yS>� �q�>��؟��QU��㽿��=�s��m\������V�F>=�����=��O�$Lٽ�VZ<j�=�+������_=�R=��+>�l^=,(?Z�
�[R"����)Ր��Y|�S}�����>�m�=Ёf=$������o/��jp��.�G��>��>< 
?���}iy>�C>������<zD�#�2>��5<���>�|�<HUI=��*=�N��@�l��󈽓��=<�]<j�<�=��6�T�e>#�+?1��>�l<?�e�sa���@"�uZ��M����f��X�	>;��>w�=�S�av��1&�a��ۼ�����P��¸=��>�k=Π�>�4����<N왾���>L������Br>�V�>�X�>�M�=6�A;����{5����}=��ҿ[�����R��q��Kq)��o�����-ƾg|H>�6=�����ȶ��9�>���=Z���w���7�(�m>H5��Lp��xQ�D���|K��I1����OG'>�����w�<-���<������f����o�6�=��J���c�IfY>�?u�?��>pc?ߥ?�(�>�D">�p�>��o���>tp?U)?��>�{>�ʈ���!�\z��N�2�`���rn���H> �>��$>�e�<ڗT�B!i��� �y�P>/��=�{����߽������ǽQ
�<��>�*k>,�)>�?�h�����R�7�鼒�v>��#>�&�>n0��"�D������9�T&����=Bä<�>�]>	,�>�s�>���>xi6>�?��f�����n=�5\>.��=�%>Ȓ*����=�y<!�_=nK��׼[�\=5�ɽ�3����M�=�K�<t/?�h?q�G?�펽�����Ǻ�AR�������՜�)N�>k��>�5�>RP\�������6���?��S����:�U�m<�ų>�OD>:ٍ��5��dƝ�O�R��d=`�!���5=Jz��G'>-o>B�=
8>��
>��R=9pe��q߿��xSm��`�B���侵д���ߜ\��@������^�D�<�~>��E<�|�=��:���=M��<]���̆���pܽj��Џ���D���C���w��b��$���K���1���E��Aż�7�� ���G� �&�����V
>��>�.�>`�M>h�>=�4>�s�=x=	=�>��>S~>�׽<	
>��V=��>`�t>�� >˒��X�w޽���[�1>Ӣ;=[��=���=��<��<��=�$\=[� >�]��9����ؽ���c	=�g�<+=�5�=�1�>r� >20���&�̯G�w� �W�>>��)?�ž9�#�'�'� �*=>�u�L�M��^�=fp]��T����� ��1o�>{k�>yԙ=���A��E�+��1�ȳ=!:[�:9������è=}���=��ɌS�Gy�ʿi���=��>n��>ptA?=�?�V�>·��"z"�AL.�$�_�1,R���	�J�I>��-Y>�S�x�����2��e�7;)������<�63��H��n��=��e>��>W>�L=�{�=~>��B>Ѕ�<��>騹>h��>�>�>o�>F>�"9��]ʿ9����6�E��`��>S�c�/&��E�J>t{��a񾁥����v="�̾�S'�A��KU�>N�K>&��>��#=L��dW4����F�ڽ�M�|�����(���g=��Ｕ��I¾[9��2��t�Ķ��&���w�M��2	��?��5>4�?�H?g?�7??ޙ���*?�r?ܓ?+mg<_�>��>�]�>��>�?�$?��?���vV�9�=���='>ΙK>v�=e���������=ر>�F9=K���<��<ol�<:�#=�ч�0��=�V �ʣ�=����#�7�ݍ"�j����)����>�h�=��ݾv6:��i���$�J�
����~6x�w�㾦��WN��-�>f_�>�j���=�O��)�K�/��̱<�C�^ϻ�؊>�0��:��;ký�!���/�� .
��̓=�K�<̮=�C9?7�2?�o�>�#��9�6�1b��NX�ip�T���[�>�b�=��<'R�<R<������5����Iǽ�3`�}5���<7��=a>��8>���=�����^)>��>b0>oH�=�Ю>*��>�0?�g�>���>�� =�ʁ�'���5��t���
�׆���:����t�o���և$��p\�y����{h�����=����?�>�= �'��:"��>c˅�!R��`�'=�`�}\�ߔ�~���1=�=,��v��<��i�>����� ��k�R���ݼh�n�BY�yBμJ?�.�=e+>f��>�c?�|�> ?ho^=\ԣ<ڹ�>$��>J��=H?m?�f�>R�>X?�s�>>	>�6潳����=��! =l;�=��*��W����=悲<;��C<��u=�5�;�W�=�:=J�:�@κs$�=s�>�O<4�����ֽ����G>�ϟ>'&?D�ؾPm9�s���q>�8��*��T>=�]!���þ�6=��}�>Ԇ�>�>d��5���~�������=n��B�p��>@�'���ڽ�(ܼ�䉾��Ѿl����=���>xe�>|�6?�,%?�?z�
�.��f�?�-�w��P���>�p;���
��Nپ��(�Y��jᾷ+��R�;q��=&ݠ�Zc�>,W�>�A�'Y��Ef��זV>���Y>�<�Z=��=Ւ�=��>6Ch>�X>�k��]���Ϳ�*��*���M���}*>�E�@왾|+E��hҽQ��=�{)��O`��u��V�>-�>��$>l&�=��=���=U펾.������%	����w,�����~��<��w�3�?=��C�>7ډ���ֽ����s�|�=����a������>�)>9�S>�"�>U�{>�1>��>#�ʻ�w?�p~>4��>��d�[�?��j=�%�>�3?��0?�T�>�*9=s�����l��n3>���<��=!��>8M>�O^��1�=��>s�v<�F��X�e>iG�;�+=˧�>�d4>t�@>�i<>�1�>r� >20���&�̯G�w� �W�>>��)?�ž9�#�'�'� �*=>�u�L�M��^�=fp]��T����� ��1o�>{k�>yԙ=���A��E�+��1�ȳ=!:[�:9������è=}���=��ɌS�Gy�ʿi���=��>n��>ptA?=�?�V�>·��"z"�AL.�$�_�1,R���	�J�I>��-Y>�S�x�����2��e�7;)������<�63��H��n��=��e>��>W>�L=�{�=~>��B>Ѕ�<��>騹>h��>�>�>o�>F>�"9��]ʿ9����6�E��`��>S�c�/&��E�J>t{��a񾁥����v="�̾�S'�A��KU�>N�K>&��>��#=L��dW4����F�ڽ�M�|�����(���g=��Ｕ��I¾[9��2��t�Ķ��&���w�M��2	��?��5>4�?�H?g?�7??ޙ���*?�r?ܓ?+mg<_�>��>�]�>��>�?�$?��?���vV�9�=���='>ΙK>v�=e���������=ر>�F9=K���<��<ol�<:�#=�ч�0��=�V �ʣ�=����#�7�ݍ"�j����)����>�h�=��ݾv6:��i���$�J�
����~6x�w�㾦��WN��-�>f_�>�j���=�O��)�K�/��̱<�C�^ϻ�؊>�0��:��;ký�!���/�� .
��̓=�K�<̮=�C9?7�2?�o�>�#��9�6�1b��NX�ip�T���[�>�b�=��<'R�<R<������5����Iǽ�3`�}5���<7��=a>��8>���=�����^)>��>b0>oH�=�Ю>*��>�0?�g�>���>�� =�ʁ�'���5��t���
�׆���:����t�o���և$��p\�y����{h�����=����?�>�= �'��:"��>c˅�!R��`�'=�`�}\�ߔ�~���1=�=,��v��<��i�>����� ��k�R���ݼh�n�BY�yBμJ?�.�=e+>f��>�c?�|�> ?ho^=\ԣ<ڹ�>$��>J��=H?m?�f�>R�>X?�s�>>	>�6潳����=��! =l;�=��*��W����=悲<;��C<��u=�5�;�W�=�:=J�:�@κs$�=�2?B}�<�7-��b���Ҿ�Ɯ����>@�����1�?;z���Ӿ���	�W_ ��'X>���>�><��>�w>E��>��ʼt(<�G!�j�J=�� ��+6�8��<@�������=fr[������  �hD/=�	>��9>V0��Lڑ>C�5?xK?g�@?�7��J�@�E�3Y���6=����K��>�����N�/�"���ӡ��^���̾�bR�����!>��<?.>�;�=+퇽h��<onk<L�'���b���=����N�>���>���>��<L}+�^�������ܿ���Cྌ�<�(�<Ju,>��Ƽm8i=+4>寷��4�={�>[z�>9�N>h�~>r��=�ǌ�mk=��=�,/�C,��xD�vVG�u�w�:kZ�[#ü��=�Ġ��=C�-��a�nk��2�޼I������0�ν�_C�,B�4(�>�q�>�>�KM=v?��>j"�>��=+��>�bC��k>SYC>w�>�g�>��?��>�J(<�f��!˭��۽i疾Fw >X��56z>q�>�'�=�}���t>r�L>��"=��q=<'��䍽�;-�G�<�Ǯ=G�>S�W><J�>D[�p2W��ƾ�r�j�+>B��>l��\5T�L��>S$��2��0Ծ3�P7�_Ȳ>��
?u�-?��>�M�>3��>^!ǽ�O��s]A;v�Ὅ]S�������=l��Mjs����<qT�~cM����(1�=�>�:>��p<f��>V\?��H?�:�>���6��A�6�=��=h>��?�p�>g�>?���Ȑ��16\����N�^�龬���s<�ܩ=�	�=�4�<�}�<l0�<�?v=O1E>w��=�]�:��=PJ�>�Z>���>�w�>�/��a*Ͻ���":�@�ڿC��Ɠ��,/Ծ^�>�x>|�=��F��+�`%���莽��<�=X>��l>�f>.7�=ҢQ:�"���˞>9����ν�=B�ܚ�����S#V��&)�
�Ƚ(���4b�=IH;�C�Ǿ��ɽ(%%��u�ns@�Y�`���;�`A�<O,?��>�B�>�&>�?���>�R�>&��>�0?��Ͻe@�>��?��?�� ?G�<?�,>�Md��X�vƾ���Ց�)>�>�?+>�)_>M��=]�ؽ��S=�[:>�L�=;C��<�����+���'�=j�=J��=K>���>��g>�_ �I����� �{�G��w�>:�6�ZK����>c�Ⱦ��	�g�$뾸��͠>[�?��?o&`>,�U>�*>�U�q�j�@��</N�<�%��v��=>�����8=hH>���������\=0 >�p!>�]9>Y�<ȅ>D�?��M?tE'?�I��}����{D�-^þ7(
>6�=T��>�`G>�]������l9־
�.���#�;(	��N�ը��k>��=mp%>�m�m@��N��<x�=�H�={�����=P �9Z�={�>O*�>�s=�P޽�%��ܽ��Ͽ����Lj!���>��#���Ҙ��Ӹ�a_�;z�;�aϧ�E}���G�>��>��>���=��������<�<����㽮Օ�b�����W���|����;����=1�߽�Ն��k<���e��H�]U7�1��]��	�>�Ɵ>�o>K˃>)�R?q<?��>���>�
?����P�>���>6�?tE
?-?1��>)�>��K=n3��罄o��IG>�^$>Ҁ�>G
>�F=��Q��ý�X=ї����<ă^>ۿr=g�l��:��NĬ= :=�+>��G>`�=T�M��"�7��m�;��o>��>�E���h>�7�WuC�vMk�0B5�I�U�<F�>4h5?��C?���>��j>�l�>e�=���Ѕ�DZ�=���c�9<�R>yc�<$�q=�~;��P�v���˺!���F�Օ
=��3>#56=���>�C?��>$9D?\�Ӿ��[��N"���A�|�>���w�>�/�>&��>�]�= ��fv���+���J�^���̮89�>V��=���<�=<�P�9h3�����c>dvP�Lim=ӑv>l��=l�>w��>?�>7�����v���U濝�����оs�g�j/"���=��<Qw�=�kz��[z<�̠�J%־:E����;>t�h>��=駽C�ӽ��;�?X��>�"��l�(��
��2D��Y�����<�C���3G�]�#�w�꽞���p��MJ���/�0-�x���Y�q� ��>)S>��?��>-?��<?z(Z>B��=���>�tF����>�?"�?
"�>��?EY�;]����9;kR�<�����>��n�44�=%2�=àY=�>>l�=>:W��>T���J����'=/��=Eƽ���;<�>3�=�#d>"��>������O��$��8����� �E�>*��!�  ?:i��]��i��p������	x>��>��>!M�>P~>R ->��8�A�>��:<ێ><&�<$ =��q=8������
&=�h1����O�<�?�=�	Y>_ɗ>V�6>�i">c>?kN?.�?������Bm:���B�=
!��g�>���=G����E�������yT������da���<���> �����=O޲=��^�U3G��.H=��.>���^s>(1Q>�=>u��>̓>�?�[I��.K��T��Y@ӿ�ȭ��H��3>2���<K�>T_<w�޽�Ȍ=��oXb�P;b��m>E�>�>$��=�{��-§�Z�*<�����7�P�ｖ)��l���!`(���Y��X�}Y����=r7�K�����O�d�y�	F"��Z���t�������_�蜰>K��>eY>G=~>��?�)�>K�p>S��>���>�w����#>Jo	?+��>�7�>I��>ΤW>��X>�%�=�)u�k��l��K��>f\ɼ٠�=+�1>���:�Q���ڼ.�Q>�����A<�h>t�>��3��DQ���>c¾={։<�:�>j�)��A�����@�Ծ��=d&���d?r<��U������xپ4ܴ�t��=�mR>Pa ?���>=Q��c�=p5�>�	>%I��L���=*X�<+�=���>���&�����=X����k��1�=��5>�}>i��0r=��>L�w?6
?��>(�G�Td��e�)��Dm����>�0��
j?/��>U*����Zg��^<�X;�y�H�~o�>�g<��>1yǽ$7�=[�:��=�"}�䨢��4&>�������<�-T>���>,p)<ϔ�=��ּ�w��@JȽ|	��������,μ~AO�������?�>����*��]��>����#�E�Ym���T2>W�D��Z-=)9J��Zx��mj���x�ݩ����J��Y�jG���uh��)������b�B�ɻ���m�5�,�wV�c'p�Dҵ��LC���A��U����>�7>�9>�6�>�1e?�P$?�>?�A>�5�>R�)��P.>�dZ>���>IE�>���>���<{c=.��=v�w�DF���	1�҉d>�>��Q>�o�=�%>��i����=�u�>0�U>ET��;�O> ����ֽ��t<�wG>R�.=>?�0���M0�:n��V���=>F،>���>x�V�ʾL>KS�{#j<n�Խ�!�=��$>��5>uS�=�!�>���>GS>*��=��ͽ%�<V�
<q	F>��+>�W)=��<$����;�=�7�<~�!>))�a�6�И����;��+�;�`�=�I=��8?5)?��,?�5B�D���xp���оL��e����o�=��A=�13�T�Ⱦȶ羸��t���p#�/CW�|���`M>~/1>��i>	�>����m齅�[�3��=TZ��?Ռ=�W��@�=��>�i�>��a>��~=4�H:��~���ۿ8���(n�=�����ھ����9>k�B�l����Ğ>�(������ڵ<:��>m����=���Zm�������;ɽ�
�&-}���¾�R��nE�".>1Ѻ��>Q<2����E�F��䐽�FB�d�Q�k�</�!�̳��C>%�>��>C2ź�zT?u��>7n��Ufʽؤ!?y�_�B
z>iJ�=�c>k�<@�>>�>"�>ԍ~>_��~D��=�v��:W=�=������S�=�j�1E"=���=���=y��K��<����'ʽ� �լ>ҭ�=�L=�0�=V�?����� ����5b�_F�=y� >�u�>��S�Bb�=�Ge<h�>�|>�>3C�3��=k�> -�>l�>%b�>P'N=j�־�6�B��W>�6�UoԽJ�M��F>�»=��R>�1g>梮< �M6���m�����Z8�=� �=G�4?r�	?��>zU�>ϟr�p�N��{ž޸�=n��8���45=F��=�/ɾ��W�-e�ث$��c���;?X��7A�> 0�>r��>��0>}��	1���eһ�BH>t܃�x�<`g�F�6�Y=<Yx�>�E(>�_>OYp=9UX�
пZ���u>mH>�����)���>�Đ��Rʾ>�'���ݜ�n2����>����EEY>�S-�?A�$���[�=�/ֽ�H�<���;X��^����v�U�='Qc���;/�:���3?�V�U<q�4��;�@��;¸�&t��40B>��>���=�Z�=�?���>��=����+��>Q�?��I�>Ӹ<8(��%��z"�>ȏ�=��>6	�>C;�<���+�M��{/>T �^��=@ �=vp`>�=��G=G��<ȇ�gz=��ܽn:���	��
�}�̼�s�;�8%<SE�>�7Ҿۂ�x`������p��k�>m��>SE�����14��YY>�6k>�~>X�= V�=��k>�U$>p�==م>�˒>�	ݾ��=n�0<|v%��D�=dS=��>lo�=HZ�=�W=��>a�E��D7���d�����=;�=�����*	?�(?=u)?Z�=�@�$����,��;���]��N4�C�������̇�7���i��	Ӿ����dF��\	��f}<�7�=$���{�=	L<�Ƚ���o�={����ڶ��D��#�=	U>}�>��>d��<����ϼcͿ'����> ��\��gA�=����귾�f�>累�~&ڽsIʼ2g#>�u��`�Լs�6�����=����̅|�x.=-^��UǾr���CX�=S����>R=y���4Dh��2�0�+�vY��s.c� �,�<�2���w���>"��>a!�<�M���)?D��>��<Ο漘�
?L�M�˛>|y����1�-�"�r�>�>>'̬=-*�=���<��5�6�5���>�J��A �=ΏQ>p|�=�c ��۲�����}��=��=�:���=�F�H$����=ξ=�oG>cW�>�);$�ݽ��BKϾX�=�U�>��R>�Ұ�:bM>@Y=\թ�3L��E�=���=!�=q�>Qr�>6�=Wԏ>�03=堈��k�����=�L>V{>��>;�ȋ=��;�=@��=�y1>-��=��g�5��ԗ'�g���,4=��
>W�(?R��>���>W�m>덷��e�-����H�&d����=���=��=._��;K�DΦ�K�Ծ[��*�����6C�>Y7>�i;>���=�q�Y#����:�=��d�b��=��?>Rz|�fx=gΏ>�8>�:<'�ü��bz˿������+>�I>���r�����`gT����j�>��ľKP���+���ڿX�T�u=%���ȡ��Q���ܗ�����}�`(T���վ���!+���)=2#��ԑ�=eDN�UO)�]M#��O��m���K=�R�F����,�=ְ?�c�=5	=S.,?�D�>,f3>�=R�?a#v����=ZS>>���=$�e<xJ�=��8=M�a��f�<�6�>|p��Q���G{>g��=��t=g�=`�X>mR�=	�@=�n�=$��<�7�E�����sr�9A8=�XM>�F�<�,Q=2	�<R�齏�'�<�����op<��>Е���z�h��=5	��f��㽩������2����l�/�>�?��>¡R>�֐<:�=T�Ѽd�&_���|���W�=,�<m��<�'>NF��I����"C���Ž�愼�>���="9>��?�&?P�?G~��D���M����䊾O�8>ʮ�>�z�=uTͽ%k��+Y�i��0�b���泾��`��^>>}Ӽ��3>e{=�����T=�s>/��=g鈽�Ԙ>����^(?>v'�>���>��o>1NL=F�c�����Ͽ*9����þv?;�9�����e�F�+;��3�a$�ѝ��!�¾�G߾/I�)d�>E%u>��t>tB>�4�;qJ{<�+��G�F���ݽ����v�� �k�9=�8P�O���W� ^ ��|���p�a�^�D��H%\�B\оOޜ����/�?��> P�>�n?��.?]J�>�i�=]�>>l-?�����[?���>FJ�>w�>�"?��?<?�h�=!큾������p�=�'=~`>�2>lG�=$=�4r�Ї:=��=�i<J.�<�P�=V�X��]<==�R>3,9>��=s��I;�; j&�<35�#&Ծ��=���>n2>y��ǽ��o'(�񗢾 >�ؾ�B��I޾枆���>Zث>��>=`:��뼕\�[|���N�ۓ;_g/=bi*�r�L>5}�;#_t�d������f�oK,>W�1>�+�=�I?)<?u@?�X��)y�i�G��U�c�[�"�>���>�׵>������X������)���,`�UF����R�=�h��<x0�zDh=�DK=�G����=s?+>?�+>	>l?��=є�>�7?�,�>�/>���� �e�8aͿ�R���V����Ǿ�`�i��v]>���-dt=��[>U4��Z��E=�f>];X>�>�^t>��/>NLI<-�/N��/ҽ\v�K��H)���ջd�$�����54ݽ-㾀�ľ���6��}�rׯ��h��Ԍ������#?��p>�B>h��>�LD?�,?���=3H�>j�?Z	=���> �>&�>C�>��?�H?��9?%�>����μ��]�B��=(�K>�S�>��>�Y�>��1=���H��^��=o֟=cv1>�=˩�<J%#=d�A>�{>ˣ�=�g�=�O�<�꼾��)�iU���2�ةT>=�<�?ξa�a���4���K~�Ziʾڋ�uػ�E��|X�>��?�O�>�o�>���<J�w;JQ_�V�^��18�Fu[=-u>�j&>������o>�
>����G�;���ŽQ�T>�~�>^�b>�'�>/�1?E�U?�u+?�*ݾ9��!{�y���OP�>�>�ۈ=-�ӻ�LԾ�#⾀�8���� �ʾȦ�����B2>~)��[��qbl����<��=_\f>�i�o]����=�j=���=U��>˂>�-[>��<6㽕�)�sgؿ�ڣ�D��{ �M��=�n�Y�ۼ�[���H��ǋ=���>U#e�&� [.=�h�>[��>��;�;Ӿ����.8���,�3�j=�B���'1��#��� ���<]�9�-Y���\�����f�m����=��q��mȾ�έ�Kі�F�?��>�{�=)�>uE?\A5?NF?7�?�U0?'A����<��>�?ͧ#?9S?�%?.�?�Ǭ>�紽�E�-����~=��=���>�7�>p �=z�t��kݽ��=)�>�5{��ݠ�h�=���=1��=8�5=VT�<��=��˾d"���8��,XE�������r��>�B�>̕K����M>0����h�ྷC������
��\�=�O�>0 �>n�>H-M>4��=�4�<� ���Nn�(\K�E��9^��=�k>+�$>�t�>�=~���۽-攽On�=z}:>/	�<�s+>�OU?��>P[�>.��c[(��%�����܅�=��>\�= �˽7�m���1��¾#�[�*�P��s���Y�yX�<�m�>��潒�P=lDP>�Lֽ�˼1zC>Oڧ<�����>u��|r=1��>�{�>]`>�q�=x0-�4X���ǿ���U�b��i߾�(�.��?��=K��f��F��t$W�H�0\f��D<:4d=�2�=�U��������޽��M�)�Ͼ�\о��پ���æɾB/���m���v�о	�	�l��\���ey��e�OS��y|پ᜾�H���;'?c�q>i>m�?��+?�� ?>��>��;(�=���>c?�f?�o?��?ױ(?�n?�Z�>P������H=ĕ�>�>���=Q_=̓M>T6>�|�8�μ�Q<±��]���
=�!���ս��=GG�<��=<��=�g�=�O�<�꼾��)�iU���2�ةT>=�<�?ξa�a���4���K~�Ziʾڋ�uػ�E��|X�>��?�O�>�o�>���<J�w;JQ_�V�^��18�Fu[=-u>�j&>������o>�
>����G�;���ŽQ�T>�~�>^�b>�'�>/�1?E�U?�u+?�*ݾ9��!{�y���OP�>�>�ۈ=-�ӻ�LԾ�#⾀�8���� �ʾȦ�����B2>~)��[��qbl����<��=_\f>�i�o]����=�j=���=U��>˂>�-[>��<6㽕�)�sgؿ�ڣ�D��{ �M��=�n�Y�ۼ�[���H��ǋ=���>U#e�&� [.=�h�>[��>��;�;Ӿ����.8���,�3�j=�B���'1��#��� ���<]�9�-Y���\�����f�m����=��q��mȾ�έ�Kі�F�?��>�{�=)�>uE?\A5?NF?7�?�U0?'A����<��>�?ͧ#?9S?�%?.�?�Ǭ>�紽�E�-����~=��=���>�7�>p �=z�t��kݽ��=)�>�5{��ݠ�h�=���=1��=8�5=VT�<��=v�=�н^������Ņμ��X>r",?i���6>��$�ŧ������R�����=@�ҽf�*�Q⽾;a(�� �>�[�;,/�=P��>{a��/]�$v�=[3���
���~�=��>�ܪ=����@Ƚ}�Z����$䂽? ���t>ܼ�>��?i.0?.6?�������W+�j8n��Vo����>K��=����?�ž��+�6,��9���'����<����=\i>f =V㙽n��=&��=�]��ټa/�>��&����=�+�>��<�,�>�E>V�>f��=?{4>^*��e�ѿX�����D��;�:��=N:>��T=7�>>�Ą>�w���G�<SF�=m�^>9�~>��>c��>��>��[=�Y��������>���վ���x䷾ay��>��[=k�ͼ)/�ՠ¾s��\<��d�&�g½�fv�¾��n�#��>�æ>^k�>J��>�f?΃
?�>@��3�>���ۗ�>+�l>\�>�?Zl?�K?y?q��>��H��ؽ*�]��>ڼY�>��>��N>]�>
����e��=��=���k�N=79����<bmz<x�=��=�{_>���"`˾㬔��I�+>x�ȾQ���`	?�Eg���F�r�<�_�
��m꽥�\�۬�b}N�#'?�����<D�>�p�>r��>q� >">Dn�H�'�'z{<C'j�cw�;}��R�>��I�ݫ{�)N=�="L���W�F� ���<|u= Ƙ����>I_W?���>UD����j���g�B|~�,֐�^�Ż@�a=xz;����sq�F���I���� �MJ���g�_!">\>KH	�2���t>����&�����=��>�7��-:>3�>�f�=5��>�R~>���>q�>��x=��A�\4���N���������s%> /����M����۳��F�>X%;���=i:+=�Q:���d>�q>i��>�rc�{)K>/&��͎�E�ž��ھn���
ͼ�X�f7>?���=��)��z:�E7�l(���䉽�r5�bDp�����6;B���?.|w>Sa|�i�>�.�>��?=��>r>�1?�I�����>���>�ن>�* ?5��>?�>�3�>d��>�;�=`ݦ���)���=�ۖ= �;=�9>��
>K��<��g��<C�k�M����<�l� (�;�%�b�s<a��<��\=���>�@5>�3
��W$�d�$�>O+>6��=��(?�j4�e��>7�G�c2��b>�G���:���վ�9�X:~�Z�+C�>ª�=���=�]�>�@��)���c��o\!�
q����m�E����`=�4>~���C\���Ǿd͎�w�,=nFN>|��>��[?��W?�E#?P����WZ�OG���V�o��1䳾\u�>T�=�4���F��,�}�!�I=���G�6�߾󼼑q�<S�j��F�+op=7�>40`�^�����>���bA�>�j=����)F�>�2�>]A�>�e>����b���kѿov����O%E�AI�=��zS�<���=�Lg>�#�>p�֟�I���}�ȽY^H>������A>�
�=o��>j\��(��<t@�<�A>��ۺ�/���K���=Bg���=�r�vC��Yy��;^!��<דٽ�(��
4�����u	?+挽#�a=���>tj�>��?ke?g=>ٻ?��P����>��	?W$W>��1?�[�>:BA?t�@?o 1?��+>��н׊��4�E�J����>{��=d}>���= ��<���=�g��Aټ�� �fmͽw��7j<�i�=lE>�[=>Im#>����
��#�v�����2�t=��(?љh���������q�����py+������������U׎�H_ż_H�>�q>��K>��> ����(�II����Ǧ����3�IP>W�=,T�q�e��)�"ɾ^.��"�\�� 8=}�M>L�8?�#T?��?�ц�OQ���/;9���ʾf�e>�(�>�սZ�>f�=�A���&�����Q�Ѿd6���>�$�=j�Y=�H>�>��W�h=�YK>�ߦ=q�=�#o=���=jۖ>>�>+؋>
tS>�14���P�.�⿋��.��~���>x_>�� �UnK��>��%> ��4ؾ����w��>�G�>)6>���>�N;>�Ӥ>��|�������յ��Gۼ
?'�!���a�W=�^�<�f.=�J��k.�0#�=/�w�T(���v�濎��;+�}�"��?��v>�a<�P�>�?`�6?z;?�=8f�>J���'�?1@?#�޽��>0�|>�?{#�>#.?tIo>�+��ި��v�;0�<���;A��=
�9>���h�=��=�Gt=�)��j|�@`=�q��߶�=�=�$>:�>n��>���<��@���#��0Y�p=n	���?0�۹=�� �K���H'G<�VY�$���E�³���o��D�>���>��Žl�=р�>�o`�7�/��޸@�P�y��#��>:�4ڃ����=q���O�������QW��M�^�<>��t>�$E? '>?#?ԉ>k(�w=o�Fq��2�>��c��7|��b��"?@U|�E'����Ǿ�fK�Rd�4,��ћ>sk�=v,��V�<>�_o=�Ť<]"=
�m>+���W�>Qu�=��=$��>�̪>UY�>1�>d7�W�Z��Q�_������1�n��=��+�e��P>������>�!��$������>�<�>c�L>�zN>8b�>�it>ӱ�<#�+=��=��m�KY��%n��/��
<r�O�+>�뀾�O=0�\�����{�?��R�k��O��&zP��>���<�>�ަ>���>�&?O$<?�>�s�=����N8?��>p�j��T%?��?r�?��?�?,�=F��IK��9��aC�}�7=���=��t>H��=�O@�S�#�$=�汽��ҽ��_��"�=�ȼ��9= �*>@�=2	�<R�齏�'�<�����op<��>Е���z�h��=5	��f��㽩������2����l�/�>�?��>¡R>�֐<:�=T�Ѽd�&_���|���W�=,�<m��<�'>NF��I����"C���Ž�愼�>���="9>��?�&?P�?G~��D���M����䊾O�8>ʮ�>�z�=uTͽ%k��+Y�i��0�b���泾��`��^>>}Ӽ��3>e{=�����T=�s>/��=g鈽�Ԙ>����^(?>v'�>���>��o>1NL=F�c�����Ͽ*9����þv?;�9�����e�F�+;��3�a$�ѝ��!�¾�G߾/I�)d�>E%u>��t>tB>�4�;qJ{<�+��G�F���ݽ����v�� �k�9=�8P�O���W� ^ ��|���p�a�^�D��H%\�B\оOޜ����/�?��> P�>�n?��.?]J�>�i�=]�>>l-?�����[?���>FJ�>w�>�"?��?<?�h�=!큾������p�=�'=~`>�2>lG�=$=�4r�Ї:=��=�i<J.�<�P�=V�X��]<==�R>3,9>��=2	�<R�齏�'�<�����op<��>Е���z�h��=5	��f��㽩������2����l�/�>�?��>¡R>�֐<:�=T�Ѽd�&_���|���W�=,�<m��<�'>NF��I����"C���Ž�愼�>���="9>��?�&?P�?G~��D���M����䊾O�8>ʮ�>�z�=uTͽ%k��+Y�i��0�b���泾��`��^>>}Ӽ��3>e{=�����T=�s>/��=g鈽�Ԙ>����^(?>v'�>���>��o>1NL=F�c�����Ͽ*9����þv?;�9�����e�F�+;��3�a$�ѝ��!�¾�G߾/I�)d�>E%u>��t>tB>�4�;qJ{<�+��G�F���ݽ����v�� �k�9=�8P�O���W� ^ ��|���p�a�^�D��H%\�B\оOޜ����/�?��> P�>�n?��.?]J�>�i�=]�>>l-?�����[?���>FJ�>w�>�"?��?<?�h�=!큾������p�=�'=~`>�2>lG�=$=�4r�Ї:=��=�i<J.�<�P�=V�X��]<==�R>3,9>��=s��I;�; j&�<35�#&Ծ��=���>n2>y��ǽ��o'(�񗢾 >�ؾ�B��I޾枆���>Zث>��>=`:��뼕\�[|���N�ۓ;_g/=bi*�r�L>5}�;#_t�d������f�oK,>W�1>�+�=�I?)<?u@?�X��)y�i�G��U�c�[�"�>���>�׵>������X������)���,`�UF����R�=�h��<x0�zDh=�DK=�G����=s?+>?�+>	>l?��=є�>�7?�,�>�/>���� �e�8aͿ�R���V����Ǿ�`�i��v]>���-dt=��[>U4��Z��E=�f>];X>�>�^t>��/>NLI<-�/N��/ҽ\v�K��H)���ջd�$�����54ݽ-㾀�ľ���6��}�rׯ��h��Ԍ������#?��p>�B>h��>�LD?�,?���=3H�>j�?Z	=���> �>&�>C�>��?�H?��9?%�>����μ��]�B��=(�K>�S�>��>�Y�>��1=���H��^��=o֟=cv1>�=˩�<J%#=d�A>�{>ˣ�=�g�=�O�<�꼾��)�iU���2�ةT>=�<�?ξa�a���4���K~�Ziʾڋ�uػ�E��|X�>��?�O�>�o�>���<J�w;JQ_�V�^��18�Fu[=-u>�j&>������o>�
>����G�;���ŽQ�T>�~�>^�b>�'�>/�1?E�U?�u+?�*ݾ9��!{�y���OP�>�>�ۈ=-�ӻ�LԾ�#⾀�8���� �ʾȦ�����B2>~)��[��qbl����<��=_\f>�i�o]����=�j=���=U��>˂>�-[>��<6㽕�)�sgؿ�ڣ�D��{ �M��=�n�Y�ۼ�[���H��ǋ=���>U#e�&� [.=�h�>[��>��;�;Ӿ����.8���,�3�j=�B���'1��#��� ���<]�9�-Y���\�����f�m����=��q��mȾ�έ�Kі�F�?��>�{�=)�>uE?\A5?NF?7�?�U0?'A����<��>�?ͧ#?9S?�%?.�?�Ǭ>�紽�E�-����~=��=���>�7�>p �=z�t��kݽ��=)�>�5{��ݠ�h�=���=1��=8�5=VT�<��=s��I;�; j&�<35�#&Ծ��=���>n2>y��ǽ��o'(�񗢾 >�ؾ�B��I޾枆���>Zث>��>=`:��뼕\�[|���N�ۓ;_g/=bi*�r�L>5}�;#_t�d������f�oK,>W�1>�+�=�I?)<?u@?�X��)y�i�G��U�c�[�"�>���>�׵>������X������)���,`�UF����R�=�h��<x0�zDh=�DK=�G����=s?+>?�+>	>l?��=є�>�7?�,�>�/>���� �e�8aͿ�R���V����Ǿ�`�i��v]>���-dt=��[>U4��Z��E=�f>];X>�>�^t>��/>NLI<-�/N��/ҽ\v�K��H)���ջd�$�����54ݽ-㾀�ľ���6��}�rׯ��h��Ԍ������#?��p>�B>h��>�LD?�,?���=3H�>j�?Z	=���> �>&�>C�>��?�H?��9?%�>����μ��]�B��=(�K>�S�>��>�Y�>��1=���H��^��=o֟=cv1>�=˩�<J%#=d�A>�{>ˣ�=^�?���=�$T��[�D�-T$���WU(?��>�]m��kv�{��E�.��0��H�H�>���>�a�>k 
<��>��ڼ����n�&>��L=�Vf>卂>K-�=9��'�Ž'|L>^���;伷/���5<���;��k>:��>���<�m�=U@X?�Z?���>���<"�
3��T�)�De��*
<7b�>�<�R�Ʀ��>k�E(b�_/��>2�Ґ�a�ͽV>�պ�G�=��b=!N#�g;�����f>�E=4���IP�=��>m��>ڍ�>]+�=*���{�N�<�}<ο�~��^�����2�=�&�=+�������3�þB"��Ƚt�����;=">p�Z>a }����<��k��8\>~8�>�/�=98��q~^�$�Ⱦ%پ	�����%���ܶ�C����¾f�p�ܷ�����Hq�J�ξvˈ�^=(k��d�>ݓ�>��?Ȗ�>��8?�b��Q>9��>�>N&�=?��>M$?%#�>j�>�'L>��<��V>��7�z���Q�PEV������=�}=��@0�<�q�=ʍ�<�f�<�2=�����7=;ك=��=^�=��K>~� ?ͩ���C���4���辀՛=��d�\y%?>�z���������窾F���&�"8���𿾟?�p�>\p>�/>�^=��Q�����<`>Ӻ:>�m���_��r�y�F�`<h�����;�;q�gC����@��))�q�%>	3=�\>Z]i?�5?��>��˾Z�&�ׯ�� �����t�]=��>U�>�z��9P��E��/#�yh"�5�.��{���^ֽ��=b�$> {>�nl�����|F->� ���40>��C==��>4>�U�>���>A�>� p>U˯�~�_��տ���	>侙�Q��g>�����ҽb�o�>�����˾���h.<[�_>�<�=!}�><��>�>�ŧ=!n�=[�H=hL�!xv�:�a�y��v¾),=�Z>��������<?q�	���u�ԛ�G`���;3���s}�>x��=�L�>@�>��?e	?�E?�S�2�R>\��>j=�<k>�u�=��?���>���>��?�K�:괯=:�@�a,��v�=��=+��=�֘>��ͽ� ��Z��zX>Ӈ+>����kO��3⽷���] 1�$�>��>��a>a��>n���V�,�b_B�O�
���!���(�$��>JN�=Zȍ>�<��`^������Ⱦ9�}�g�0�X؍��
 ?��>�-�>��>��i���c��>?g�<�}!=>=L߼���v5>���=>.�۾�m��'�Q�p��=��>���>F�F<\A?G?S��>�V9�%�'���c)��	��'���1���>!��n�	�\۾�چ�:n�T�=�v��=u_����=��p>;�D>�;���D�X�s>�:뽣3½5�'>����潔�i=I�>=p�>�D>�)>m�V�hA�����d����f���
��l��>���>��=�ʘ�d���ܾ�9᝾�����v����>=e�=�Ԭ>z�>4�=���<���I���-�޼v���:!�-�.X�#�D�&�F�*�G�m�S�	��<�,8�Sw޼�Mڽ�A����։������/�>(��>��E>�)�=^6�>���>~��>2�W>V5?/�3>Ɇ�>W:�>���>��F>..�>���>G��>�4>�v>�[ֽb����;ӑ�=�۞>�I�=�T=E�>��6>)��=��=�'����t���=y!�=��L>%�>�x!>�B�=<�+?Һ�"��݂��覾��ǽ�U��+?8*p��_����B�9�􍾅H8�h��e�y�sf�=�?��?Ԉ>�I>6���D�:犳<�> x�=a��= C���5=��>3��=;��:��A���	��E>�^>9B�>:4>��r?�U?�?��>;�E!�Y�jJ^�}��ǩ��p�>�6<�tٽ�����2k+��_��#S���̾V?��� >y��=��L>��>�J�{��=��!�;->c�=������H�=�ך>�7�>jL�=*��R�h��0��
�����W�i{ɾ�{S��W<�7���\�K��>(��=pA����<4X>m��>��>��>V�>&Z�=u�>�G�u�A� �N=+�N�vx�r�7�����8=Pf=(���f����۽��|�|��%����佭�q��u�2��Ŷ]>��->�>�l3=�?2�C?p?��j=n�\>#ʣ>�\����z�]{q>$8?!10?H�=?&�?�>����
��JE�E�8�m���s)3�t�=�,=�<.\>ąQ=Q�v=k=U,�����<9A>���=� >�PC>oQ�=Մ?H���a�$��F��WǾ^s�Y�e���?�������ș=m�J�B����;
�ńC�5X=j�>�d?/+�>	�>Z]�=��ؽh����Y�=MP�=L����<Ԍ�@e<>���>�C
�ܐ��l��H��ba��D�=�Y>��>>�=�K?��[?��>���<9���9����!8�6����mt�!~�=�V}<c��>��=�B	�XB���K�2�طg��[��+N>�c�=t(>��+=lf���<3�O��B�޼�\4���6>>�ۢ>]͋>�T�?�^�佁����Ćȿ
���r�ɾ6��)��J� �1�� �ú��>��O����>���x���	�>d??�:�>�.4>�j���ٽS���g4��W�����v�R�7�J��o9�=�J���+��3_�0q.��~w�_�
�U�=�(��葾�������Dlk>uTj>��[>ޤ�>MB�>P� ?��2?�3��Aڇ>\W�>���=W~>�cf>$��>���>7��>�#�>�|=�������v^8�&�1>�;[>�+<(�7=�=T>
O��w1U=j����>�~f�=�ʏ=?��$�;=�>�Q,>�Ǖ=��ļ�~�>���e�۾oؾ]n��;��S�K>!݁>����:�>�'��wDT�������z����w=7X��2����)=;H*>�B>eG>�L>�Vͽ��𼺪̽&�M�����h(T>�\�=�2>ƛ:>vУ�C���|޽
4��Y�=��a>>W�?��$?x�?��^��ݛ��,��Y(��h��k��=�H�>*��>�z>b���'iݾ������T���Ù���2�
�	>M�����a%�>;#>>�;ْ>QE>Z��4>`���E���u{[��>3^q�>��=��Kѿdͦ�������k>D4�=ξT>�C>�@�>����a���v��~o�14C>�\8>vT�>���>qq�>���>�,@�
��!m��윀�Em�����DT�|�*�_������2U�N��<?�?�ȶ�=-����ȇ��)��3�r���z�?�>x|T>��=��^>l�?E��>�>�e�>�v>�u��s�D<�eg�"�����h>�=�>
�,>��O>D���[�"�c;v���t�j���=�~��X>94>(*=?�>�RB>-�B��܎��j`=�>MI=+X>��?>=HU����޽>�>TϾVp�>^��sѫ�'ԙ��ޡ>6�C�lN��F|��I�d��J���n�ǟƽD�����e�aۋ�	���>�x6>��R���y���8�V�J>��=�Ys���]=(��=6;��Ť�:/r$> M��\�⼲ݙ���޽�E�T�c>�,�>\8?��>S��:�����-��w,�A���p	?M��>L˽>4}>�{]�d�g���S��ȯ�HB������EƼ��&>X�m=���=��=���=�Ec<�WԽ�d=ɑ���>F�X<ԡ2���E>�Y>��>hA�=vJ��8���)ܿ�h��T�*��,���#>t��=	�B�B+�����>�Z��zj;�z�<�e=/?�>j�r>��>P�g=��>N_�>S�8��\n�C�' ��r���q�ȾA_¾HlŽ9I����<<传��$g��������s(�W_���P��֗�����#�>�[�>�"=�;?R�?"�?s�'?;��>=L�>DI ����:�}�%�=M@��1�=�!?b2�>bB>\*>D�ƽ�����>>��>><>�@v>��E=�m�=�o�=2t��N��gי=�>���DZ�L�=`Dt=�_�>W1�>�~�>���e�۾oؾ]n��;��S�K>!݁>����:�>�'��wDT�������z����w=7X��2����)=;H*>�B>eG>�L>�Vͽ��𼺪̽&�M�����h(T>�\�=�2>ƛ:>vУ�C���|޽
4��Y�=��a>>W�?��$?x�?��^��ݛ��,��Y(��h��k��=�H�>*��>�z>b���'iݾ������T���Ù���2�
�	>M�����a%�>;#>>�;ْ>QE>Z��4>`���E���u{[��>3^q�>��=��Kѿdͦ�������k>D4�=ξT>�C>�@�>����a���v��~o�14C>�\8>vT�>���>qq�>���>�,@�
��!m��윀�Em�����DT�|�*�_������2U�N��<?�?�ȶ�=-����ȇ��)��3�r���z�?�>x|T>��=��^>l�?E��>�>�e�>�v>�u��s�D<�eg�"�����h>�=�>
�,>��O>D���[�"�c;v���t�j���=�~��X>94>(*=?�>�RB>-�B��܎��j`=�>MI=+X>��?>=HU����~�>���e�۾oؾ]n��;��S�K>!݁>����:�>�'��wDT�������z����w=7X��2����)=;H*>�B>eG>�L>�Vͽ��𼺪̽&�M�����h(T>�\�=�2>ƛ:>vУ�C���|޽
4��Y�=��a>>W�?��$?x�?��^��ݛ��,��Y(��h��k��=�H�>*��>�z>b���'iݾ������T���Ù���2�
�	>M�����a%�>;#>>�;ْ>QE>Z��4>`���E���u{[��>3^q�>��=��Kѿdͦ�������k>D4�=ξT>�C>�@�>����a���v��~o�14C>�\8>vT�>���>qq�>���>�,@�
��!m��윀�Em�����DT�|�*�_������2U�N��<?�?�ȶ�=-����ȇ��)��3�r���z�?�>x|T>��=��^>l�?E��>�>�e�>�v>�u��s�D<�eg�"�����h>�=�>
�,>��O>D���[�"�c;v���t�j���=�~��X>94>(*=?�>�RB>-�B��܎��j`=�>MI=+X>��?>=HU����޽>�>TϾVp�>^��sѫ�'ԙ��ޡ>6�C�lN��F|��I�d��J���n�ǟƽD�����e�aۋ�	���>�x6>��R���y���8�V�J>��=�Ys���]=(��=6;��Ť�:/r$> M��\�⼲ݙ���޽�E�T�c>�,�>\8?��>S��:�����-��w,�A���p	?M��>L˽>4}>�{]�d�g���S��ȯ�HB������EƼ��&>X�m=���=��=���=�Ec<�WԽ�d=ɑ���>F�X<ԡ2���E>�Y>��>hA�=vJ��8���)ܿ�h��T�*��,���#>t��=	�B�B+�����>�Z��zj;�z�<�e=/?�>j�r>��>P�g=��>N_�>S�8��\n�C�' ��r���q�ȾA_¾HlŽ9I����<<传��$g��������s(�W_���P��֗�����#�>�[�>�"=�;?R�?"�?s�'?;��>=L�>DI ����:�}�%�=M@��1�=�!?b2�>bB>\*>D�ƽ�����>>��>><>�@v>��E=�m�=�o�=2t��N��gי=�>���DZ�L�=`Dt=�_�>W1�>��>�	>��e��,`��?���h=JU?�J��0�o��f$?��	�@�M���C��kξ	��=���>��>�B�>:��>*�V��=��7��U9�3> �@�,ҽ�e�]N�>����\Z�d�F������N�#�>Yf>Rr�>�L�>*nj?˽K?E[G?�﷾���&�B�-�[����݄>�+*?g��=�=��S.l�����$�T�\N$�'!;Ѝ�=5eȼ'�;���>Ì=(m�=\=�=�R޽�s">�7M>�%n�6%e�P�N=N�L>|��>e�?��>$�=W���<ξ��ڿG֥��Y��jH����=��ɽL�d��c��sa����پ�y��^n���O>\��>���>Eֆ=ѥ8�XZ�>�;o���"�x����J��_�������f����>�ؚ߽.���ƾC�=���I�P�.�Y��E����v���D�Ӂ�>�6��>�Z�>��R?+�a?�?��J�/?m0�<��?=�W���?N.?��;?�$?���>ȓ�=U�ξ��X��lP�7&.�?�����==��=4�>�y���F�Pa%=��<����4��mä<!�#�A<婒<yM�=3�>�>��Ƚ�jO��W���=�Mw�ƚ=/Ha?��/�w�;��?]���ͯ�=�Ǿ�a��9SU��>�#��u�>68q>&Hս�w=�9<�!�@�z	w>����t��.�<Y��=����}U��U@��N�8���Bؓ����=��>w@>m�0?l�5?�?%?�zp��ّþ���,慾�x!>� ?w�¼5�ξ��E�P��U�v�+��־��S>�˼�U >1�">��r=uĀ>'nͽ0�����=�.�ҏn�r{>���=Ψ�<3��>�H�>
�d>uN>v��pX%����|����ʾ����ԭ�~ִ=;���S_$����=�Ι��`��GE���u��
>�Uh> ��>�E�>b>=>��<,0���S߽�
ｶr¾7��,1���ܼ�[5�=(�X�tǽ�������=CAK��(A��e�Sv����ɶy����:��>.L�>��>@,?P?R�G?���>�u@���*?�:ͽ��>a夾׃?�?5�?f?�A�>{@{=�����.,�ŉ��?a�<�>>V�>)��=�+���a> 1c>"B|<˫O�g{�>Vgs��9��|��=96^=��=��9=�;>�rr>H@I���l��j��d"�.�?:���|����A���>Sg/�����o����ѾY"���Psk�	:�>½�>1�=ɔ�>��j���ͽ�h�>.W	�h�1a�=7�<Wl,���%���"���þ��̾bf>>uۭ>�9$<u�D?��?e.?X5a���>�M����)��7�~$'�d\�>A��� a�>���Z(�u�T����1����P�(y=>ls6>C�x=��?��h>8W�=�z�:HwF>;����l>�/���5�>V`s>�X�>�@�>�Ma>��׽�s~�r�������;+�"�H�H
q������C��]�=9h��p�^c���ʡ�4��g�=rm;=JT4=��ƽ�m��*7��I����! �1��������ƾ�a���=Q��N�=ɖ���=�W�{�R�u�(��aԽ���G����¾E��>� �%ʘ>ֿ�>ɨ-?��@?Њ?��?���><�>42�>�k]=��>L�>>�ڲ>�&?�$?�g�> �>MP&�����Ƚ�_�D���z=�S8=U?=_�<�P<�y~)��ǃ��� ��=
���<e�n=+(>Y�=Q��=%�}>��̽��W�AEX��>M����缧�F?}櫾�+쾗n�{�1�����=��X�M=8��=7�o��@־�� 	�>mbk>��@�I�=�n��"�z��i<	Ҕ�k���҆>��>�>�;���"�q��BwQ��uо��t|>��e>4�3?�}?]3:?RZ5�� -��J����e����x>�=�>���> �㾤���Y4���R�S�"�nѾ~�;>/�=���>�X>(-�=J̅>B��<�|�w��H�=���Ҧ>-���%>{�H>��b>�8>
�w>�J�<��3�����ϭ�-Ҳ�_���Z7�O>&��=k�*�������K��З��{���ŗ={L>t�>>y�Y>�f8>�cJ>@�	>�fb��m�����R����%޾����Ԥ���20>t�V=,^x�h�����<�j=��B�So-��d���󽵯������p-�>��+=���>V,�>"�I?w�9?��$?c�O��{�>HW>2#U>>���˿>�>XV�>Z�?��?��?I�=Fx��畾n�Y���?�H�}=�;�>І>�񶽸��=; �<c{'�iB<>��;#j5=RP<���=�_>�zY>�V>���>刎>��?���j�p�I���پ4<=��`?�����
��U���>tV�=lV׾�k�i���q)پ޾�<ۼ���>��q>��ݼ_f>��C�	�˽��>r�h;�! �W+�=%�;=s7=a���b⏽Y����S|��S��=�A�>�ky>��6?='?�4?�����=��I$��J3����n>�;�>���>bM+�}������$1��:'����l�Q>Զ��0&�=��I>�>3��>O$�=�"4��T���o>>[����>�H$����=���=�c�>�P�>�>��(��{���ѿ���F��Q��E�C=S��<Fh�=����SԾ�@=�!1���Ƶ��DȾ+�=�8�>�<\>�>�a�>��Z�$+оX$��/�!j߾�ʼ�������;㼼1�2_2�q
��U�v=W�%��l���D��9`�݉�}�q��'����>n0=k�>cZ�>v�C?H�T?�Х>|U��?�y�>~ב>m�ľ���>�h�>�x�>��?q�?-�>��'wF=�;�����h;З�=��>�"p==��<4au=��>�˞�}Fo��dS=�>���=X	�=S�2>��1>�|�=�>�0�=�Ǽ�q+8��+�XBᾔ�⽒7?�Pʾ4U>�֏�O>8�پa����ľpu�=�����>�H��Ѷ�>U7t<��>LDf=�E=���=jWj:_->׬����=W|=d�r�1<��%�;�*>�~a=��=eEd>|�!>XO�>hF?w)A?t�O?'���оn`�Ʊ��O��"D����>]���$�<�pc>��,�׿���i<5���<��=�����>�w[����=�Ւ=G$)�@�	��G=j&�>h�����>�A>�����=w��=��>b��<�aI���>2�ۿV��������R⽺��=���"&��:���>�c������x>(�w�*����8���ݾs>ܾq�$=!���S�$��R������qM�\|���5���k��\�G�<�H�'z��qƊ�ߜG��-��K���V*=1�[������~�|�>��e>^��=dտ>�%?~��>N��>����#��>'�o��aq=���=�o+>c��>-�>�=�ߙ>ʂ;'>��[%�zk�<xb�7�;�.>�k>0ý�����n>v�<�m�+,!>ѕ|<�O��!��YP�D �=ٽ�V�>4M�> ݾf;������=��)����>�d��!w�=c��A�>��7>��Ǿw��ħk=���>��?	���$�>�qf>�e��σ$<��=�v��è<�>�Ι�#�(��>=3W>_�����<r�.>���=6�=�G�=��A�tے>ӥ"?Ab1?T0C?�|��g'�G���7�Z:���[׽>�!=�O	���=�K�>p���ʽz>���缙�Q=L�J=3�˺?�9>�f=ӹ<f᜽�>b��=��r=Z?�s�K<���<?M>= ��=.O>4�W,�զ�QH���̭�Q쾴�=���X�=��>�B�<�8�=}��T���D7޾h�t�I�P��,�H>�B��?��.C��5�;�-d�ƥ��a�b�`�h�������7/�o�>t�����ve����C������BG=��z��!��A�ͽt��>� d=	A�=ھ>��>x��>*h�>)P1�o��>���{Q(>`�½��:>���>x�j>��=��Խ�v�!��>1�뽢�B�$�>�&>��޽�e'>)�k>3�$���м՜ӽ�ҳ���wg>�-�=��Խ�9��|%��=�z>��>���= �ྰ��_ ����*>�Fw<D��>�r�O �>Vz�Urm��=9\D���&����x����> �=��>cq�<��;<Qb�=p��V꽗Z����=�������<D�(=mBN��}����� X�<>�>�=-�<�e�=�=k>uz?�1Z?_iR?KY�������g��4�B��H��I��>.hJ>���	���A�q>R>ϊ�������~�����>x�T�����s�>��o�Aw����P�Y�i�������=��=e��=�6`>*��>k�I> ���*����7���%3
�hq	�3l�=Bt�=1>:M�=��!>�h>>�S����>�.�{��J
>Jb6> ��  �k���R�I�=�B=]�:�����꠽?m�������Ɉ= ʇ>p f���9�n�<z��� 2���<�9��+��=�h�>KL�>xJ3>���>���><�=�=G>�I��<v>�r�wf�=k-�����=kC�>s��>�r�=H:�>�,6���>dE�]���с%�3~�(Ľ��0>���>J=>���=wD%�l�<y9�=܌��g�G�ˣ=����q�f��pS>�&B<�>�0�=�Ǽ�q+8��+�XBᾔ�⽒7?�Pʾ4U>�֏�O>8�پa����ľpu�=�����>�H��Ѷ�>U7t<��>LDf=�E=���=jWj:_->׬����=W|=d�r�1<��%�;�*>�~a=��=eEd>|�!>XO�>hF?w)A?t�O?'���оn`�Ʊ��O��"D����>]���$�<�pc>��,�׿���i<5���<��=�����>�w[����=�Ւ=G$)�@�	��G=j&�>h�����>�A>�����=w��=��>b��<�aI���>2�ۿV��������R⽺��=���"&��:���>�c������x>(�w�*����8���ݾs>ܾq�$=!���S�$��R������qM�\|���5���k��\�G�<�H�'z��qƊ�ߜG��-��K���V*=1�[������~�|�>��e>^��=dտ>�%?~��>N��>����#��>'�o��aq=���=�o+>c��>-�>�=�ߙ>ʂ;'>��[%�zk�<xb�7�;�.>�k>0ý�����n>v�<�m�+,!>ѕ|<�O��!��YP�D �=ٽ�V�>4M�> ݾf;������=��)����>�d��!w�=c��A�>��7>��Ǿw��ħk=���>��?	���$�>�qf>�e��σ$<��=�v��è<�>�Ι�#�(��>=3W>_�����<r�.>���=6�=�G�=��A�tے>ӥ"?Ab1?T0C?�|��g'�G���7�Z:���[׽>�!=�O	���=�K�>p���ʽz>���缙�Q=L�J=3�˺?�9>�f=ӹ<f᜽�>b��=��r=Z?�s�K<���<?M>= ��=.O>4�W,�զ�QH���̭�Q쾴�=���X�=��>�B�<�8�=}��T���D7޾h�t�I�P��,�H>�B��?��.C��5�;�-d�ƥ��a�b�`�h�������7/�o�>t�����ve����C������BG=��z��!��A�ͽt��>� d=	A�=ھ>��>x��>*h�>)P1�o��>���{Q(>`�½��:>���>x�j>��=��Խ�v�!��>1�뽢�B�$�>�&>��޽�e'>)�k>3�$���м՜ӽ�ҳ���wg>�-�=��Խ�9��|%��=�z>#֮>���>sf'�'��뜾1�� ����F<?�/ι eh=b=�^@}���������� ��%��Fʾ���ž���>�D�<2HE>�j>�����}�=+OA=Ô�3݇�ӷ�<Ro>IrU�-�=W=�ɼ=N�-�sWངz�=Pu���'�>+�?��[?�_a?��Q<�{��Q���$���?���g�=�*/?6�h>-9>p�Ҿ���M)��w���׾���t���ul�=3	�:�����X�>
3�<4��m{9�޵�=|�l�=�� >�z=�c�=@fI>~ӑ=���=Z�b<T�(>�����.�x9�gqľ2%���κ�ҟD����;�-���F��.��{�>���>�Ū>�%��6>�DA>���>8Xx�v�3��B>�ϻ���C���[7����u�=h>=ļ.��=���k=�p*��V�G\����=�{Q�tp� �|�O��>.��<o$=D#�<X;�>�t?�W?!���#
�>6z[=w�0>�[ >�&E>�Vo>�>f��>H�C?��%?X�?�J8<V�ɽ��뼦�Z<�㧽Χk<�,>�ׇ=�j=�v$>��q�[���P��)<\���S��%�=ڨe=7`)>x�a>�@�� -�B$���P��ol���6=J9"?�v�oj�BB�C�Ⱦ&�I�c��`B��;�/l�Y���R)�>�[�<<v�={�7=�V�v5^>��'>oK=���
�r=��>��;��e5�����ݽ�Gh�W�����)>�ԽT�v>�0?V�Q?��D?!H��:����4��#�y����nq�*�>��>{{�>�i��Ǭ������ 侵��� =O��>'�a��K��ve>�����8����B��=L���eĭ���>���=!&`>g�>Y�>|.�=�z��E>�տ$h��-�I���0�ݣ9=�Hb��>d�=�7�I�?��@��T����yP>Ư�=Ɠ�=���=v&>�ڮ>���>�v��<��[�0�č5���K�G����д�"�=�V�׾ݽv�m�	������`[�
|=����8!���Ž i?ٳ�>#�t����=R�?�g?��>�S�s�?Z�>O@h>@�>�P�=���>�+?��>D��>eb�>+!�>�Uu�Ɍ?��Ji>UsG>�[�<�*�=Z;>�ȼ-Ȃ<���<�gt=˂��y�
L�����r;�H>C�>۲i�#֮>���>sf'�'��뜾1�� ����F<?�/ι eh=b=�^@}���������� ��%��Fʾ���ž���>�D�<2HE>�j>�����}�=+OA=Ô�3݇�ӷ�<Ro>IrU�-�=W=�ɼ=N�-�sWངz�=Pu���'�>+�?��[?�_a?��Q<�{��Q���$���?���g�=�*/?6�h>-9>p�Ҿ���M)��w���׾���t���ul�=3	�:�����X�>
3�<4��m{9�޵�=|�l�=�� >�z=�c�=@fI>~ӑ=���=Z�b<T�(>�����.�x9�gqľ2%���κ�ҟD����;�-���F��.��{�>���>�Ū>�%��6>�DA>���>8Xx�v�3��B>�ϻ���C���[7����u�=h>=ļ.��=���k=�p*��V�G\����=�{Q�tp� �|�O��>.��<o$=D#�<X;�>�t?�W?!���#
�>6z[=w�0>�[ >�&E>�Vo>�>f��>H�C?��%?X�?�J8<V�ɽ��뼦�Z<�㧽Χk<�,>�ׇ=�j=�v$>��q�[���P��)<\���S��%�=ڨe=7`)>#֮>���>sf'�'��뜾1�� ����F<?�/ι eh=b=�^@}���������� ��%��Fʾ���ž���>�D�<2HE>�j>�����}�=+OA=Ô�3݇�ӷ�<Ro>IrU�-�=W=�ɼ=N�-�sWངz�=Pu���'�>+�?��[?�_a?��Q<�{��Q���$���?���g�=�*/?6�h>-9>p�Ҿ���M)��w���׾���t���ul�=3	�:�����X�>
3�<4��m{9�޵�=|�l�=�� >�z=�c�=@fI>~ӑ=���=Z�b<T�(>�����.�x9�gqľ2%���κ�ҟD����;�-���F��.��{�>���>�Ū>�%��6>�DA>���>8Xx�v�3��B>�ϻ���C���[7����u�=h>=ļ.��=���k=�p*��V�G\����=�{Q�tp� �|�O��>.��<o$=D#�<X;�>�t?�W?!���#
�>6z[=w�0>�[ >�&E>�Vo>�>f��>H�C?��%?X�?�J8<V�ɽ��뼦�Z<�㧽Χk<�,>�ׇ=�j=�v$>��q�[���P��)<\���S��%�=ڨe=7`)>x�a>�@�� -�B$���P��ol���6=J9"?�v�oj�BB�C�Ⱦ&�I�c��`B��;�/l�Y���R)�>�[�<<v�={�7=�V�v5^>��'>oK=���
�r=��>��;��e5�����ݽ�Gh�W�����)>�ԽT�v>�0?V�Q?��D?!H��:����4��#�y����nq�*�>��>{{�>�i��Ǭ������ 侵��� =O��>'�a��K��ve>�����8����B��=L���eĭ���>���=!&`>g�>Y�>|.�=�z��E>�տ$h��-�I���0�ݣ9=�Hb��>d�=�7�I�?��@��T����yP>Ư�=Ɠ�=���=v&>�ڮ>���>�v��<��[�0�č5���K�G����д�"�=�V�׾ݽv�m�	������`[�
|=����8!���Ž i?ٳ�>#�t����=R�?�g?��>�S�s�?Z�>O@h>@�>�P�=���>�+?��>D��>eb�>+!�>�Uu�Ɍ?��Ji>UsG>�[�<�*�=Z;>�ȼ-Ȃ<���<�gt=˂��y�
L�����r;�H>C�>۲i���?�d�>7V۾��"�5%=�;����<}&?w�1���>B�!�:>4�ܾɹ>ߢ!=$"X��վ�?޾��V}>�͚>߽^>�z>]C�:��7��=�ϼ'�;��{=��=#e��Ǌ{>p����:��~v�Z,���+�s\*��%V>�}!?��b?�2?<h1>������Ҿ�͍>#�wn�>�R>c#?���<�C�,��P��nF�N����߽�7�=�g�="Q�=�n;>�r�>6q��Z��Е�>%����z�=cS>g
�>�CS>�}>b(>Xb>�/3>nRO���տ����+�E=�}Vl�_?�=�a�=\�ʽ�_5����=�.��{����������Y��<.�`>$
�<%C�<���<�8�����pE��!|���U��R즽���xM���:��]��=)�������o���z�&̊�Bsa�r������j��f߫>���=5�@>x2�>H�?=�?�m?�5h����>�J��X�>��˽I�>Q����Z=�"�>��#?�{�>ؿ
?�]��Sq�Y⌽�"Z=b�l<�=�+S>�J >�<x��]ԽBO80&������X�;��<[�=�8=������=C?�h*>{eE�ګe�v�W��q�������eZ?�Q%�8��>Ǒ���>ȾR�a>�>�(a*��Ǿ��J=Z��>	Y>@�%>��==N@��7����=Dj>3"&��}z���>�r@><��>��=��<,~�%Y���s=�)q=��>�#!?��z?��/?)�N�w�J��!ݾ��ݾ�o��>^+�v?�
:=
7�>4jž�I���2{�ʈ��$�Ҫ���2���>��<>�hZ>o?)Ԯ>�ɉ����%">b�K�K)C�0-{�d8>]H�=�?�=q��>�+�>f�}��5���̿{���p���a����o�=�*�=�f'�G��;o7A>I��=�>���m߾|��M������W�!>�u?�?u�˽��s�_�5�����u�vA;����Z�,�l߽�3d=�����'���T��!k��	��3����ڍL��R�ѭ>��>�Ȕ>p?�L?J�B?@��>Rƅ�N?~��!R��%���R�>��>��>�?ّ4?<��>:�i��WR��������c�y;��-��=�|>X��<Tn�?�;�3{!��l��U:�p�ӽ��<�.s=o��=-�==�w>��?wb弅�������3����5|?>�G?0�3�/^>�b���>�Fi��q�	埾E 4�S���(�#=��(?Ҿ_>��s���;)y�>[[>���N��=�
�e�.;�諾���<_2�:PQ=�B�@e��2����Z��U�>1>B5>���>�_R?�)?�D9��=�����Ҿk��s2>�h�<����_þj�Ӿ7��O���z�!����p����� Έ>�j�=�O���ȯ����r�ر�Ƀ�=��[�=d- �GZ�>bR�>	��>�>�zQ=�Ԉ��븾�HʿW��v�>�f�8��2��@�>��%>�Vz������,��˾�)����x�{����V=�> �=]*����=�#��H�=���?N���
���,��e��[�˽'�$��o!>�iW��i���l�RB�wO-�U�j��O��Ƈ����/�E��>@[�>�_�>׆�>��L?W�>��=����S�>���H�*?�KܼMy�>�?��.?i�&? �!?���>T�|�Pyd��5t��.��Υ=�l�=WX>�o�>��L>��)=t��W��<p�(>}� �F*]��X<}��=B>%�)>��>��
?��>f���`,�4�U����(R��H?5qq��, >jZ� і>g�>}�	>�58�v�+[例���.�=�=��>a�=Em�=|�>DH0��?'>�i����^�.飼�\Z���L�D��=�י��e��k>�V ���r>�|M>��T>�N?�m�?w�U?���9k���m��f�x���=�_�>9f�<l���ؾ��$��BC��4ǾU�%� e�@��9]T>����>� �Q�$<�8����9�<�>1��:o>7ֱ=K�n>x͒>�&�>���>o��>���=N����ο𡏿$S(��c"��{��\l&>��h���c�4̦�s`t>��ս����{�������>�KE�
����_��;�<6��>�@�=m�����|�w�j1g��Ξ����=va%�$��=����[�����|���Q�+�νg}[��M��|��([���r>կy��R=�o�>`�8?��>+��>K�g�*u�>	ח���>ԫO��<>��:>���>Q�>�?���>
cM>�g{�Sr���-=��;=�l�=M�R>:&=�^^�m�����=�%>*�1�Kf=;ܷ=�>=fV���ݳ��>�=>��>q��>IPԾ�E� 9S�� 3�� V�+�$?ӡ㾫��>_|����>�5@�=Y�X�N�оK ��]����־#��>.�>��<C��=��*C�'ӱ=?�X;S��=Ɵ��� >��x<`9ý�z(<71���Լ ����J>Y��=�#h>Su?��W?5�?3�@�$�
"���%
������>��>�=2BԾE㾠
о�=�p��Gn��T��U�@>����;���=��_<{�r��=�&U>�bA�G�=,&�̠\>��=��>���>R4�=�z/� g���������s;���&��d<'��=��"�K��%����֕��7Y�%����悔�	�>�����c=���:H˂>)�TS���=��r���þ+@"�u����*ן��T&>�ۗ��uA��Jf��Q��غ�Jb��e�D��V��;5q��[�><�(=f�?>E|?@*E?<O�>Ù?�Q��W?��p=9�>N=�D̯>�x>�ʵ=�]"?�|4?�l�>q?�m�	ă�4����ĥ<��h>��=��:>���G�L�5P =������=TWT=f  =
��v�̽�`=�>&�9>,;�>a�S�'��?����&��'A�Hﴽ&9?��z��Ȉ>۠��S���(>��R>�e`�����о�
۽ia���K>DJ���=�Z�<*1>g�&<ќ=tΒ���
��*>ĉ�<���Q�������wO�����Q�ּ-�b=^)>�Q
>��?w�>��>�#m=�y����E��5���+�>9�!m�,��>�m��:ʾ��7yݾł���D	��>��� >�3�>�0d�����2���b=1���� S>T�>�2}�^A=W>��i>��=�,O>�x�>�>��S��޽2�b%����������UW��	b=��Q=1�I�(���ZT�:�)��V���0��e�� �=k�=}́>1�>�mG>-���Lj��>4"���������ϹݾWB=�1����=��TV�^��ꙑ�ZĽA�ν$�S����Ϛ��{�>>�x>6f?ձ�>;j6?us?3�ǾSt�>�|�=��>j�+>�>�`y>e$�>�X?��? )�>F�>_��Aƈ��]C>R�c>Y��<o��=��7>z�K�����cS�==YD>6<�<¼�=k\6>��=�<�p��t
�>���=���>j�ݽＧ����ǀ+��^(=ZϢ=-�? Ͼl���W�<-Q>�车J���`�q	���˾�� ?�y ?�@>;�=�܅=�oS>X�T�Ԧ��S�=h,]=?���=�A<�y�>,Ib�5�����D�<i��Ѽ-���A>'Q>��>ۗ1?��%?��	?쾮�_�hNF��|�z|n�Vh����?u\>���F�;m�9=53��8e˾�dP��� ��z:<)�/>�Ҷ��c��S��=2P2>̴��C�Y���>9b=�
=��<�C>'r�>���>�1J>А�;��!����啿�G�����3��ꌾ�>:>��c�->�G��sw>�>Y�$��+ξ&�>YR��o�8��1?��>cl����3>��O����䤾�c���K�ϵ��>!�c�{�����RF<u		��|���wg�Q1R���_�R�&��!K�9��>N٥>#��>jZ^>IzR?v�0?�?a⎾��>$]�=3����9o���=�uR?6h�>�g�>3��>3�B���������Y�Ƕ&>h��=���=e=�őh>��<7
�O�*;\���9r޺���|Y�=r�i�/��=_"�>c��C��?�>��5=�Eľ������D�þh�>�G?kD��d=d�{�+�`,���M��w�������������}3�״>����ׂ�<Azo>AC`�O����>�q��V���x�>��>�4��;�,�=V+���G3��F>�.�=9�'>�>b�?@y,?D�>Vir��!��=�����Zs���^_>���>�/i>>\=���ྵ4����ǰ/=��;CD�=��q>\t-=z����t >N��=jj��a�=���>}�o���
���>�m�=+b�<�o�>�%>Z����Sѽ����ƿ^�����Ü���&=?҃>d�Q=�z�w�j�:�*��ݾ�z�=bJ/=���>�g=��>�2?�P�>�>��-�R컽���H���q���k�qNپ��5�
6½#׀����<
�^�E��v��c�'�oY��*����
�s�G���>�]�>0�F>t��>�d�>�"?HQ?L�?>�� ?I�8�g��#|�G׽I�>�@�>܀�>b�>�$�_Z����JA%�<\�=8�)=�,�<7�>(.�>g�@�'e�R�6>�{��x�;J�W=-?���=��=�I�=���=q[>���>�⋽j%�,Ǿ�[��T���Y���>G%����>�;=��q��<��ɱ�;�Ʒ<.D�2r���������),>�Gg��>���q�=�2�����-��6S���w�E�>1�>��<��AA��韽�B=Z������q>9��>r�L?���>��>ZB������D�����`����ؼ�W�>���>��><�K��+%��@�}e���<����'>Z}�=D�>�Ev�#��=�p2>ξ����N=^>�Bh> hq� �l�u>�+N>|N�>��>1�=vT�9j�����6�X��u{�����FE��&M�T#���]ݾw�Ƽ��=����߿��o׾�ȶ=%	�=5MM>r�>qֆ�=����7�;-�r�/�[���O�ҋ���3���=N^�q���?'�X`R�9:�T��RO���V̸�G`���^`��R�>np>�߼>�|�>�U?�\)?��6?��]\�>��P�i���ǖ�<x%c>6��>�O�>y?���>���>ժ�=��<��0�P`>[���~�<g6�>R��=��e=�3>�� ��[f�Icj��=H���3Qq�nG��c�>��>��>|	�>���h�㾢2ƾ�f��d��<e>�]?b�㾫Y���ͽ���/�P��LR�����OX׾a��=q<>U�I�֯A�?��>��e>V"Z���G�Թ�= ^������>�L>�\�f2>���9���{ܧ���
>��>���>�^�>=?��>�%?�_�����E%�!�?���8=��a>���>>9�>��\=y��ȥk�,q�&D��}z��e>�́;�LV>�`��<�2C=1+�<�P�1�D��;>��B�<�$�Y��21_> 6^>�>�G��
n��[y��Կ	ד�qd߾�$,��>���vA����=�)H>:ʓ�)��M�5��pq=`�>f �%�;>���>SN���F����>���>&n*��xӾ�8���â��q����>V�ռ��l�p�h��A=��j��{"��7�����=_Ž�i��/ s��c>h(�>��>�o>��-?�I4?�E�>bP��x�[>?ѽ�X�=�oY���f;ِ>|H�>y��>��>֬�>^#\�[���\|���>ޘ4=��F>\<>�;?>:t"<��^�
ik;je���>i\-=ɥ;�>���>y�>H��=��>x���H;G՚�`t-��=�l����d�>�1���?6>0؋�jG���?��zɾ}�$=�R>
�?z�>�Ӓ>���>����8 W��AP��^�=E>NE���k�o�Q�f!�dM�=�}������� �=0J�=�h!>�D��Z|=�-O�=�.�>�^B?kp�>�&e�sڼ���Ū��3Ҿ^;�=�>�w
�ւ>�)A��o������°�?5;b-�S�e����e`E=�MS>�<�=ƗA=�$���D>[�<-)���%>�I�;�m�>Di�>�֨=�d��R���IT�M�=t.����[�K�e���k�9>�Vƽ%���H܃�0�=�=�K��a�޽�K�=K�b�˺Z�+>�B�<TS����>��߾8������@ڽ�l��J8ɾa~��C�j�O�� ����"���n�@s��Q��9����r��FI8�#����l=��>��>�����n>�^K?&z3?Az�>Y��?T1�����>�A>��>O&?�"?a�4>�^��䞷�!D	�Q�ܽ���B<>�&>$=�=jR&<n�n=�	�K$�=1;�=F�%>|[}��n��\�c�W����ᘼ�1�=�00>���=�ל>׃���a���V����F�پ�$����>H:ļ� �>�{S���T=<eB�ss ��ߙ�g�>��>�W?�a�>�>�>���=�����L=᫾�;�"VY>���=����a(�>?�=+ �=��Z��S*�y�Ͻëg=4C>��C>��m<}Ty>Z�#?��,?�� ?�5 ���x��a ��<������ s=~{�>Dp�3q�>Bc��)ϾJbJ��)��޾]R>��I���z>'�ܽ�����>-v�>V�p��_= <Q����AH�<u���ᾜ>�Ͷ>>�\���˙��J���`���뿇���))���=��=��>�0>���n�=?٥����d�Ǽp�>�?ڂ�>�9�==+`<7�=:�� B��ڈ�*V���wk�u����׾0ٽW�ֽ��N=�����'�4
�R;���_Խ޲=;"��Aoc��TJ��	�>W��>xpQ=��,=]{=?l?�8�>��#��O>�R�{�1>R@y�|��>'U�>���>�y->�7����׾��!�Rjf�4x��Xe+>�ƥ>��=���=U9F>�z���K5>��=C�=UMq�_�~=3��=����<��=;/�=��7>~�>S�1�dI�=�m >�x[��-�<ż�t>�)�<HH?� ��P���\SZ��9-�,P
��>�2	?0]??��D>@�>��>�5��y�o�e>
>$A�K�v=��>�O>Ą>d�]>��>T��#��a�Q��=;�=��,>8��=���>?�g?@��>�
��������+r��b
�5A%��K>���=p4z>ak�5�Ծ�e���Q��򠾈��=t�6=�޲=�r�΀=����6�>�b��s ��N
��rf���$���Ƽ�.p>�m>�>��=����K��a��'׿�Q���j�WJ�Uu�= Q�=(�'>�ʌ>7e>�x����۾�����9>�"�>��?�Nr>t
��2N���P>�7������ M�gRr��9��w���'c���F@����>�̶O��f�8�<�,��H��h%Ž��½d�3��m��D?߿?o>���=$�[?ז*?j*�>�#��u�>��J�H;k>_��>v"?N�?�.?!V�>�I�>����8F�Ѧ1�����>��m>�~w=�](>!�3>pF��C�Ӽ�="ʢ��轔�E=��=�WJ���G�	}=��g<�Ѕ> n�>��>
ֽ ���L���#�h�����?��{��ы>�d��V���(�b}8�3��0��>��>i�?�U>��a>mM�>��=��л	��<�o�=h����Ŗ= �=b�¼�R���zݽ*g�������⼻�&�`����>�jW?A�7?om?	�	�&���Z¾�Y����x��þƖ�<��^>3��>*�=+��1���3���D����$���ߝ�����=�>_{>4->	��`���om<������t�5=�+>E~E>寿=`�����beX��̰<{�����]�D�0�+X>��Z=�������{���A��+>���=3�a>��=���e�X�W��oP>�>����^��<\K6�.ܾ����>��*Z��ij�g�tFN�;b����<�q[�")��W7�����Q�>�)=~>��d>�r�?�O�?%wX?ñk�㊤>���=	��>*��>���>�#2?�*?�*&>��E>�������=!bN�@�-�L�]�=����=I�>�8�=H>!L�=�/�<��L=�=UZ<Q�4�k�=6>#�O>��o>��>�Q�>�E���D4�a�j]>����+2����>��=<�>d�ȼiG�-��[�ui�4꯼&�t>L�>&��>�eY>���>���M�P�	�̬[�c7��f<?�c>t�*>��v=Vࡽ�P%�{�����^S>M��<��$>�\߼���>ԝO?�?W�?�uC��M��kb����	νw����$>\aH�d�8>��џվ?��E68�.,��<⬔��ԏ�$I�R�)=�^r>y��>���=(Ľq��2�����=�t>8ʖ>�7>L)콿���9}̾�&�O`˿Ԥ�����'�j�>0�>�z���������_�ʾM����]�>*�>���>���>���>sz> Ɉ��Ci��FA>R�l�B�
= p�l��� ���-���LA>q2:�Ym�=w��;H��=bM�͗P;�D���>׽�ɹ����<ͯ�;6R�>3/�>n�%><��>�*&?���>��?��λr��>,��xw>����X��>?�>W�>ѿ�>��=7}E�ٻžc/����y�>Ơ�<���<v`�=F�|>@���u����J<�T<ϴs���M>��G>N卽�*�x�>(��=ݹ�<W �=F���w�q�pF���[�l�j�Y�_>�?�<�O&?��p�#���m�Cm�l���=��>��X?�aH>x��>��j=�̕=�k�:��-�Ǘ?>B&�= ���+�.=!,>�+J�U�I=_��=K������9 M>��	>�,>i�=�N(>H�S?�?Ƥ�>݀2��k⾰�@�N�8�ώ�=Bk�=�y�>t�=�)�,�=����V3
�����)W>�+=D�>�y_�cѺ��>o�l��ʺ	>�!�=~��+q>_j
>�A>���>�F�>�Z=���<�@��g,��C�����m?������!��=m�=��p��q�����9�	�V��퍚�$�ؼ�,�<Ut��II��#�
�)��=�1����Z���C��*�d�_��3�.������� ִ��/��z��ъ��ו��u��0�����¾],ľĉa�ػ�J?��<��>�E�>}-;?�MB?k��>J(V>¢?��뾰�I�?��>Z�? E#?s ?忳>�HU�
���y@�1�*�g?�=�q=;m=Us�=0ی>ͣںq˯=\��=ϏѽE�I�"�K��9�<��*�<v!�=�>|��={pu>�H���4Q���3�g�!��>��l>�t>hN/�Y��>�Ƞ���Ծ=�<X�?���	�pv;���=�@?J_�>'mu>o��P~n=\t�7�p=*!k>β�=Ay�	��<Q��M��i�>�L/���Ǿ7:��A�T=9Op>��f>:m�=w@G>�R?i7?h$?ŭ������0J����ͳ�=C|e=d�>j�i�9|�~�,=w���=���Z�߾�N��\���Sü?��>�&p�G����N�=���I��3 >N,@>1܇��#=���=��=��
?2��>��<��R��G���\��̿6ڣ�o�����侒r�qr��V�(>j2��]��Ľ�}��ͯ��NQ��3�ݽСk<H�v�Z��
�<t����$������� ����=L0���̾I���;���q����j>��H�G�����*��OR�ղd�\\׾g�r�������?� �>�Fv>�ڡ>�@e?Y�?\°>�W�>�1'?�߾��>�@?�0�>Q{1?��C?M?2��>��-�o����"�%G��I>���=���=��>�V1>o0V�$w�:���="T=It
=�G<�/c�ee��	f�=6�>���=�ø=�׾�����6�.V'��g��⾍q';I΄>�
�y�?Ꞹ�	/;��d��rX������̾��=�� ?���>(�.>�B>�DT<Eǂ= ½���7%.T>�,���v�=b�>o�X=�U�=.��҆��k�^���:>�/�=���=�w=̇��V=?k&�>T�`?����U��Đ���#�9���mȪ�e�=&�&=�CC=Aߞ=×��xzݾ*�t�&��?�=�d=Gs>�P�=����o�>�x��6zj����=��=޻q�>U��>U΀>���>M�>m�(=/��=.x������Ɵ�9�����l=����=�Ƚ��=t�c��0�<!q�5�񾦱ｔ����-�&d���{=��U��h�=}b���%����Z��??=-0����u�g��m>>��־ϳ+��_̾H��xX��K�m�Va��V�ξn��������<75?���>��'>�(�=mC?!�/?O��=���>o	$?q��{��>'�?���>lA)?��<?��?���>�d����y���=3v��t���j��� ��(>A>]׹=�=j,>5[�<Y�F��6�ڳM�b
�0 �;�(�=iE>��=��׻���H���'��hG�79��[����&?�X��?�6>פ(����i��P�i��>�>��)?[��>��l>�HK=�U�<(� >�ս�,�=7E>eY�=�����B�=٠>��y=�P��po�;(`�<p�A�U��=�0>a:B>�q>Z��?E�i?�9?� ��
"$�Հ[��>����ȿ��(��>�)�=!~��	�=�*��C�YX`�6�F���]�a��<Z�>v�c���H=l݌>�;?�#�{��<ľ�<�[X�+h\;��\>W�>�"�>_S�>�p>p���!hg���ݾ��⿃x���㸽�?���9�f����t0���=��>-���Ewܾ	���>�!���ؽ�\�y����+����=��u�ʘ�=>":<���׏�������		��(_��B��)�=�����༾v��Q��uƖ��W�����랛�lJ
��:?���
g#����>kAP?WL?�8?�ϛ�↔>�ӫ���ཟ�	?h.�>�p?�6?t�:?�1�>�]=��i��v��d�:�V�;af���=K<���=�4>s�@=��q=��=]k=4����<@{���K��Kr�=��>�$>{�L>I��>�ſ�-t[���$��I�f��۬�>�PD?�����?n����U��K���@�Y^��v%?�pG?�cV?q�>��>�$T=���a<u>��˽��Ȏ�>��=��i�;�>g��=����S z�� ��F3��*�=�,�=�{&� �ټ#��>h�T?�@X?Դ5?���N"��Uؾ4n�1Ƚش[;�\?�U�>Ri�>�g=8��E+����(Cj<�Fм�o>z*>s&�;�|>�dO>)R��3����=h+W���㻷~�=C�/>ł�>O>e>��j<����*������ɿ��p�����`��>}�p>�G�=<7�>?H=}�ᶾ�����޽��D>��=d��ޟ½�ړ�'˲���P�өнQ�q�������i����� �v���T�/�4=Dj�=h�K�1�j�֨��=x��������{��se�=+�=�(�>l<���>80�>1�/?�DN?�>��=�"?�
��)>Y�?v��><H?U�?%}>#�(>o�=���<�7�5���褽�
>��,������r=X�=��<o�=<���=T�>�>s|>�=�H=\�=�V>�z�=���>"-���O�"7#���a�j�۾q!���tB?)�������x��H���vȾ�н�ļ1���J����������>h_�=�"=�J>��F+�=d�*>I5e�z���G#> vg�g)���;��s>\Q�=����G��i�靤;���=�/?kUK?"mP?�o�<���H�׾nJ�9����B>I?nA%>Z�>�0>-����]C��g�»׾#�Ͻ��N��N�>�W6>�B�ǍS>���6ܽ�W^=�x�<��E��O�=��_>`9>0�=��z>P�>�6�=f=���=��� ܐ����*f���˽Eñ�."A�V��=!��=z�پ�r��]J��䭾�#������N>�= >��>#�~=�)h>AH>�;���T���i��zx��Y�>l�4=@S�Vx�/U�=�����^�~����Ľ0�#�7g��ۮ���>k��<=G�>JE>J�4?�iA?�@?U����a>���>>��=�\�>���>&a>F�>��=@�?K>�>,��>��j��.Ͼ�ʽ�\e�q�=�;>;^�=cꮼ�]�<깳=7�#=��Ž���m5��%2��̛���>��>'��={l>y����k��3��v��6��j��rk]?<«��?�T��d���8��I��E����i޽8����u����#��ܯ>ec�>��G</rH=A�
��=R�$> �1���p�1��>�BD>�א;e�>�n�=Ѿ�<a��=v���X����˽��L>J�O?�`Q?�G?�1��^��@�$Z@�گ���z�=w?�G?r�?��`>��?;L����_,��U�����)�b�?�x>�k>(��;��>�3m�ӿ�;��C;EM�=��<Co1>��V>p.�>�ʐ>XH�>%4>�^��hPԽ�K����ӿ��O�2�A��WT����4�:>��4=w�p��R���qѽ2�վ�NE�(�>�	ڼ8��=' >�_�=a⍾w�H��:�!���৭�6�������=0č�Bh��z���W�������Γ��#z����Yx.��^?����n��>9�k>HZ�>�DK>�!?��1?(�"?��N���>f۳>��=wO�=X-s>J$1>���=�.4>fB?���>��>�v��9��σ�D�Y�i��=1[	>��=�O=U�=~���|���"��͠k�z\��Yx���\���A>�/>Y�:>��_>y�;���7������gh�("�!KA�Y'?(Ⱥ�M�Ѿ�����7���!�<Lʾ���;-t �˘���-���I�>�U>�?�L�:>(T-=z�:>CƼ�I��S�����%><������V#�=��O>YV�=�J��Z��Ԟ�p��dD>@�_?N"?)�>?DF�=��
�O�s��=T�*�@����@<?�ު>y��>Ȳ�>��&��������������^���`%�>;˛>����GN�>⢍�Fj.=g�B=�ּE���b�>=�n>w�`<l�n=���>u�E;@�!>߄�=����y1ٿ���\-��JǾ�;����y�����p>κ�w�꽅���`����X�;�o�� ��/)�<�ꊾx�>���=0�o�;9e��)��vH�����M��h�ݽ��J>6���1C�c��ߤ�I"G��l�ԧ�
wE��`�,<���r,���?Dv>�=>����,?n[>?�?�޽1��> ��>S#�]�J�". >�3>-�=�8>~�?�\>��>���B&�7����Q����q)*=�v<��W:��=��<	up��Hܼ�^X=^5��� ���=���=�k<���=f�=�w���0�"M���B���߀Q�$m)?�]5�na�@/�����C�$��[��;o�x���L+�������>X6V>%�m��7�<럱�i��=��^=�^G�4�@��J>��=M����΃>kϐ<�Ŕ�TV=������ݴ���1E<�??h�M? $??�3���?�W��&4�#���3�=u�?DJ]>X��>}9e>?zu�^z%�L+6��.�Tہ��9�h�>qEw>�3!��]�>u�˼�K<u��b����d�=��>{O\>>sMI>���>�؆>�h(>��t=�CI��I������N���V�߁V>4Ђ<I��d�����TǾh.� ��Oz�=,
�=?1��g�(=e��=v�z=�(1���߾`m�����Xxž1a侈�پG� >��a�(ʾ�_��^�������i�� 5�d�2�k[d��l^�yw:��&�>Ya�>�>!�l?\Q?˃)?἖�ި�>��>��,>_��>�6�>=�>r�>�P�=K~?*l�>_v�>�)=<i6����r >&�Y>�8>��=*�J7�=��(<�fļ�D<�9c���=\#C��o�pC�<bYP=;�>x�>�F���T6����ߔK����2-��64+?+�S�N9����Jm��Ӿp��;Y���z�{zJ<��q����D�>-EL>k�<��t>L�H�:�n�)5�=�$^�������<��=؂���e{=�>4V�a��jP�����m�*���S>l�<?��R?�J?�����,���2����;q�<JL�>��>��>8�=��ﾐٗ���,�����&�����>%>�/%����>����{�� ~��U6>�l�=��t>���>�>�'�=�V>F��>���=�U��� +�6�ο	����%Ծ�o����i>�>������=�"��o?��:�<��<������ �R>�˘>�7@�d*>�^>�ؾ�����ݬ������	����ʾ.o�>|���hX{��㞾�� �l���ॾ"��C�C�s&�M�J��B�*]�>���>q
~>�H>2�?��?�T?/G��i�>Q{�>���=�z�>� �>�b�>d1�>:YI=��>��>e�>Z���邡��Z�=�v>�\�=-�>r��>}zD���3>$ڧ=������$��ҽ��<��=�j�w�>�&�>�8�>2D8?��N�aɾc��Ϩ.��ߠ������>�cI�8��Ly�� �����r�=:��>���>O2f>�G�>�˖>|��=w��> \V�*?��]���y>^N�<�$��������սS�����=����@E� ���D�e9�=��;�Y>=�F?�'?�d�>q"��:�(�`�vF�r$�=H�5>�t	>e��=?�>�	���,�<����ֱ�B����_���%>�ų>ٜ�=N�>De=�\�=��=�(>Giq��U�>Y*�>���=_+�=�)>�d�>�>��w��S��W�������Q�t�ܾ��>%t��_ã����=�D��
�>Ǌ��g���U�ǥ=�>��W�A�߼��/����G=��.�<�/��ֳ�����ɾF�������F����=�I���0�j`��R����u���o��f���W����뻍B�>ƶ�>'��>��	?=y*?��7?���I��>-�}>�D?@j?R�>J�=��i=�>�E>.�!>�`�=5]a���PJ��?�h=����A��^�L=�ͩ<���=�(]=8�=�������<�Jj=��L��V����=�9>�D�= �-?.gξh��������h����w�apq>D�ݾh����t�����9u/��T>��>dwP>�0	?�D ?]�>��>$�>��="Ï=��)�M�b��w�=R�h�é׽�6���L�=�r���&��\����D��p����ż���=C�x=a�=��{? ?}cC?姾�&�2s��O��q�������l=K�:>�y2=��/������V�^�N���~���=�~�>�j	��6��h>^aѽz`�>�6�>�&L�F�=�ܸ��>�)�>�#�>�J=��H�2���H���ֿ2uc�ݹ�����8�>�T�[A뾈
��1"�]��>�خ����f�������N��3�Ž �C=\ k�@���Wz<#����g��_j�?}f�����Nې��w>R�n��<�=��ľ�x-<�����F��(����|��Y��+�C��;9�;>���>�G�>OY?��>�$V?}�6?��G> �?��>�=K?[��>Y��>2[|>k��>#-�=	k@�s7c��D�<1g��i��$���b��=��!>f�=�6�=}C]��Z���ּj��=O��=�2L���q�]H5����<��>p�B>Z �=!2?�BҾ����p&��F���+>�Vw���>;����c���������>hݟ>!�>���>�??S?�|�>���=F�@=�	���v���R����=5">��>�K@��]=>ό��Z	���b=�Pv<8����'����.>�m�=sOq>�;?�k?),?f��/Z����վ0[���s����>w�N>(�=�bƾ崾Z�����ʾ�*N�K|���j>'@�>cq�>�b>���=�ű��@I���o>�Tl���+�^x=�T�>S���a��=LjI>J�=�_��G�����#dR�����ힾr��>=ś��X@���&�4G��������~>�T�����<͌���>�j7������Q��I��n{������:d�p��^����ɠ<�⽃=t�w�t�׽,9���?>N�-��ۣ��X2��z�t<Nђ=L��>��	?��?��?^]"?�D?��=%?�?3_?��>� �>�W+>C�>h�M>���>Ә>�˽7~���������kEͽ�3>�Ή>�T>K�H5�=N6`=��<�
> ���=[��=T����f�<�L>x{�>\F?�Ҿ��$�`����A�l�!�㽺�?���?��0�žф	�x����a<��>���>���>��??ԙ>by�>��>B49���3��u4�Q��<�x>����q�=��;dUG>o2ܽ�F�=,֡�`\)�k5���9=��R>y�"=�)k>�N?8l�>ʬ?��	���׾�ò�P���[�=�G�����>>��=��=g��bc�U�^�9��Ծ�r<�йq��}.>���>yK=�.�>j�>sT��|����*=��F��n�=&(=�0
>�3>;�=M��r���MV�����>b�䓑�� �m��>���Y����~�������>Nq�_i���E��1�=�{R��������Z̒�=�A���8�
T ��;�-�����侩�׾C=(�۽�+�=�r��������6�O����N�<��g���/��Õ�S5����>R&?OF
?�5?��b?\?�����>0��>9�8?��?'��>ޥ2><�>��>n���
�C.B=��h��i���ރ=�',>L��<cZ>P>��(=�	���Z�:ϡ=8>���:9fY<��<d�[=�=�8!>'y>Yw>?���,\վ����I!>��Mm��G�>h~�>MV����¾�����n���G��>�*�>�J�>R
�=
��>n��>��>d�E>�9��!��	���*>�!���Ξ�T�z���=�%o=S�p���M�}�5<#C�o|�zB=g�}<(��<�w�=̩]?!I8?�  ?���P�~�=�û�.�q�^v����>D��>�<�>���y̪�x�M����Д(�J՗�Z}H�p�.>�I>O�>"M>EF>�޽��P>0<�>��Ä=-��=��>p M>8�>��>��w<B���=˾	����,C����������>P3�Ku�T��=@��>��>���:Y��N��Rd��T��OÎ=������B�m���)��b�=��6�5��D���Ҿcf��N�=�����
��ո�S7R���߽�����wɽs'߽��|�%����o>.C�>��>d�>��?��?�> �v�L��=���=�u?�*�=�\>��q>��)>N�q>�d ?���>�N�ţ̽��M��+�=��2>�?��Lz�=;�>���=xU-=8ہ�y�>܃�>����~���pW�"���q(<i�>I?�>�~?�Q۾�k��(��9���UͽD��>$	�1.>7�����b�׾����(��f��>�>#��>��>�ka>A�> 6��[�U���B�;~����;�Fx=M�{�;\�<ty<C������t̼�F>�]i;ͽ�$g�<�a>�(?I�>)T?ڏ�S����qs�����=�¾�>>k&>�t�>Wb���>;g	��)3��1ؾ�x�:P���JQ>6�>�Y9>yT�>��>��!>Km2��m��Ļ���ký#'>r�>	E>QpB���r��=��r9ʿ��B��ս��������f��]��#��S">R��=<)>�e��؈�=#���䙾X*�����c���,��}��AC��k>�q0��_�'�.<Z>15���s>�9�(�+�Lq�	_�jI#��~H�/[��(�߽o��=o
�*�?��?ͺ�>;t?v*?7%A?���v��> k��#ҼM�w>�.�>�x?�?�>	m	>�L��y����TL����~�U=�k�<{=:��=ͦ1=��t��b!>ye>iŜ=n
�=�^�=H�A=�	a<S,.<���<�>�2�>�?"��^�sV������S��I�[<Ũ>yt�=��>r�=ɕW�����¢��;�'�>�?���>��p>��>��=d�)t����Y�h{?����ID�=_J>��O�.��= ����p^<�欽��x�[�=`5�=��>��=�Ϗ>;�?�F?{�2?{�C�fr��3޾8Ɛ�H/�8�S�n>۷$>�<�>��V;�~��5��U
�S�������X&�>��O>*�=��X>�R�>\�P>�$�9����D��lTh��O
=���>Ьk>hb�>w�w�i���ϑ�B�������Z����n�Ѿ�����%ٽ�!;M�羧Z�� ���1M���W=~�c>�hN=�4޽6Sg�H���=�!>vI��U���)#�ū6�U����-�Čk�Y^Z�!p<���p=3KŽi=�o4�\T��>�4��{��8�Ž�����->Ù-?~"�=h0�=JA0?��1?e~�>>�x>��>Y8����b��<�=T�>G�>'�>�/�>VB�*5����l�۝���x>V�>���=�.>�X>	Q����<Tt>d�=��.˽�=uU=�Є;p��=���=]O>�n?MI�oN���e۾�R龎������>�H>��>?R��e���esp���������2o�>�:?��>|��>�w�>�=�Ƚ�c�;s�R�[�<s�=�]Y=@� =���=!�_>Y��=�N�=2��=�������=X��<��=e~н���>bV??ɖ�>}��>_�J𜻡�T�pO���G$���Vs�>�>(�>+�}=�� �ыھ��jǷ�FP��c2M���>�T=�c�<��9>�C'>�7<�E�˻���**��Y���>sz>���>k>Z8�<e~���G'���߿�W�V(��"��6���ه����������9��@�	�*\���<Ҿ�>5���8�>���ҝ��ʣ��^��<�~������g3C����m�%�z��o;ʲ�����������;�%V�Ćs��o���4���!�G=��@���?L�-?H}�>:�2?|I?�I(?�ì���<�\��F�>`n�<|r�=�$>w��>�8��*]ӽk�<*o޽P�	)�sÆ>���=$`=�M���U<��<>�;͒�<Q��Z���Ž�]�����~U���=�|.>CpA>Ƚ�>���r���U̾ǁ��������O~>�5�x��>7O����J��f'�+T=���<H��>��>k'�>��>Z؀>��>w� �#I��6=����dL�sW��D�&>)�L���ս;��+��[:��\��b�=�=П>��i>g�Q?�?vM?�R�d�z��H���b!���U����au�>[9K>�>[69���.����E����߾|5�ޯʾ��=�؛=v��=~�.>;B�<3�x=*Z|= 	�<�����n�dY��bm>�2$>/#>3J�:b�����Y���]�t�:b�������c�ߖ!�R����	=���Sξ��	=�0�:
A5�ي��#�=}�A��Q+���S���Ⱦ�Ų�* q>K3X�Rϲ��c]�t�ƾ�!�������=����=�����y��Z���W�%G:�B3���9��>�#��=�P�>A�>q�
>$5���7?ɐ/? �>I��A?�ӏ<�O�=O�*>�A?k��=��>gz>6t�>�t�=g����ڽ��!�s!>�4M>� ݻل=CZ->t�k��\�G�`>6��>Uh>��`��ܽlgԼy��=�=�W>��>��)?����q�?_¾cJ������T$�/0	?sk=�W?��m�{ꑾࢳ�U
ϽF�R>i
?e��>���>&�>q�=_!%>�:���{������9�	��cs� ~f�/��<F*���N���;m?��cƽ,q���b>��=���=�F�;�<t>��W?�v_>]k�>���<��s޾J�����R�n��k>��D>˼�=\��L�*k"�[G��������
����*>�)>3���'�>E�>xJ>{��d��=��:��k��:�X>���>eB>V��;4*���X�� �`ڿJ<���0�[�ϾK�F�`8��觾@���wҾM����=r����px>�`�J���|������2T�Q�?���7����T�����b���$A�{�N>�TD���=l��ܻ��0����gc5�rp��e:�`*:��P6��@���?��W?�>��l?g�n?y�K?��,��>;���(l<mD�>\�=��>v��=U'��}I���=1�>�<��tʾ�3�k�T=��c=�=y��<��#��X��{�!>���=��F=�3�5�O�����Ǽ�d�=T/>C&C>���>�4�=�ES�rjN��uؾ
A��dq��+c?�yL�Ȧ,�i~���B��}Q�]l�t�r���E�[  ��l">�o?hʏ>;1T>�&D>�>��,�x�s:��:�{�J��},��F�<ɫ�=Z4=d��=�-��x��6j�̚�*��=c\�; �>�'A?�3-?�M?�"4�+�Z�aTd�=^�:������{V?�Yy>~
>׽뼄����{����(�3!6�j-��%���
P>}�<V���w�=�8 >h�_=
�?��>����E��<"$<���=�>�:�>�>ɾ�:��a��mw����xĿ�^�h�)1�:��������B���?��w�< �@��O"�ϾS�-B�>C�U>�^�>�I�>��/>c�4>���@�L���g��+6������윾�`F��R�=�}��'���/}���2N��ӽ}́�
~�b7P������������>#�t>���>rj�>;�.?pM?&�0?h+!=[�C?�X�>���=7z6�X��>2��>�&?ͳ?��>�[X>7�yɤ�����a��A9<�N=�n~='<�=��~���=I�K=���W;�ϭ�i.�;CA��.=�˦=:��=�>>*��>t�>gF?��JѾ����}t�p?+�?����+;籾�&��_�%���܎/����g�����->�K�>L�n>wͩ>�Oo<�)_=��<T������ۈ>��B>뤳����5��=��<>����3�|½䥄<�5�=���=���>�'?@�?��b?Tо���X�lp5�&A��Mm>�O�>
<�=����}.��Q�������􃾺&��������>�콮�=�>���<��=��L���=�J�=5��H���z�;���=�ܜ>\��>X�>����ʾ�տ�Ϸ�^��yl^���ý�\=��=��e�P�Ͻ松,��������=�͜>>ђK>D�^>�Г> ��>��<�Bžv9����(���[���p���흑<������)��)��e�����猛�뒆�qV�ҁ"�9���ߞL��0�>��>??Y;�>�z8?�S�>[]�kW\��Q?�>2�O>��p>x?q��>�N3?�x?��O>��D<�6@����w�@���=$��v��s>v�"�����{.$��K�=2>]X>u��<��4;�(�;��?�/ռ{=>��4>Z?��<<�Y�`-�֖)��������>͇&?�d)����4��=�iz>�Ľ��]�e�W��/�� >�a?��"?>[>lxT=C�>2'>�����C>���ю����;�@�� ,���8>-?M�0M �k�M���Xܽې;>m�>6��>�-*?z�?��L?�������CBj��`j�����]�ɾ��=�~=[�ǾD=���7XѾmj!���)�7'C�x�P�?�{>�+�X���8�~>?�ֽ$�&>�##>�9f> A���HϽ���U�.>��4>t�?+�->�n�=����a���ֿ�w���ٱ�H--���J�C�`Z�X�!��K�"�������u�W����>�>�"�=��ݼ�G�=[�>d�� @����p��������t�.#��Ŕ<��H���`��}�Y��0ꇾ����9h��̓���򽽈ѽ���.��>Ļ�>�]?�~u>��=?Ӟ+?<?��>,�S?�@?��ڽ`<W�(�D?>,?XUL?�;?	��>HZ��1��5���L4���F=����K[=�Q�=E{=`5��$F�*>>���=!L=�.�=�3<Ȥ����= Zt=��>N>�4�>���=T:���9$��iH�$� �+�`?�R���2Q>��b�:�ƽ��_�m�W�C[U�v�$���>�I+?��?���>h����<��-N>�14��L>i�R=j���P����=���<���;w�&;Fy�vu�O��=�2*�+�=�Z>��S>�z�>kI"? �r?�ۡ�w����pe8�T���0C���s?�8v>�n�=��J>������E��� R�V.'��K=ނK>|t���<7�l>���;R�|>U�F=���=輺��90�=�=��R=�܀<�5�>��M=hU>�z���-������ $�D
���->����վ����5v�x�������0p�k���`�>ic.<m��<�!b��� =o�J���\����ʫ*��m����T�0U��m��E�D�s��l&��_2�����¾�轭��Ɛx��`����R�p��>oѠ>��>щ=_�,?�I1?P�4?�,=4K?�"w>�)f�5�`<¨?�ݼ>�ME?ͻ+?~�>�s�=�Y> �.��:�=�B�6�0=���<{׿�Lo�<Q��=���=�R�=�<*j:>��=d���1=Jr�<D�>���=����ގ�`�:����t#�C5����(>�M>�a'��	��E�������`�I�U�A�ǖ���o�T�=3z�>�=�>��>~Q8=O}f>�� <�-��[l���սL
�<��)>M�=Č�=�Dp=��+��m$��Z<= "����ռ�A%>��>�N?A-?xk?�����v�K{��\r���¾��=|�>�>��z�"�ٽx���������x�_���U)���{K>����\+=�u>�@>�l�=��=5k^>�2��,�=k���Z�=j��>��=z�=�	+���6��9=¿��wC���	��e%=5�>
���:V�B��=��z��� >\.�=��6<��i��f>D۹�����;���;�'G���Ҿ蝷�����jO�����^۔���3s��
����������1Մ�"g��;u� ��4�>��>��> �4=�^E?��5?�J�>�.�>��K?]l># �@Cn>*�+?s6�>7VI?�E?��?S��>� >v�����$����b�|����<��=%[=�=��
�O�[=,p=�N�=y�=.(�!��<"��=W�">A�>	6�>��>�T9�	'�Cb
��>�C>���>�c��A��dྯ�%>��Ⱦ\%=)�)�]�����1�1�L�>��z>�L�=�_x��2F>�馽#�:���=��>YV<�&����_>�m��=W!>Xu��^�?�I�%�<f�>��=��= F?�8?J�?��O��Ӷ�S�L�+E�y��~�����>�;>
��>>	�=�e����������i
��¾%W/�A�r>��Ͻ��=�~c��^��=��	����>�0�E<>4�<T�>�%=��{>���>��>��s�s�)���ʿ�秿�nj�Z���>��=�
4�M��ޫ���h>�;M�=�����y���>)�#>�y>{�ͽ/��=�����S��в��ו��T������Kվ�X|�ä��C=8�@�ྉs>�c�� �<��a%�#Y��s��2�f�~�ѽ�9�>��=�?�>��?��0>9��>���>$
�=��?(u7=���>@����>r5A��(?��?�+�> ?��_�nE���ֽ��=�T4<q��=ю%>" >2G>�|�=N!=|��%�h����.3=�ۻI|I=��=�0>]�w=���>b��>d:��z~�S�2�ú�����;�>w6�+��>Z'��XI>e�h���E>5'�r��ߎ-��A���(>� �>8u>�:�=���>�轶�H��x|<��=ý����6�>�H��=�7�r����*��E�g�H�h�BM�=W`r>�x3?�	L?�&�>�����U�R�T�A�60���Ҿ��r>z'�>Z�>ʅ[����02��������������=��7=K�=>�}!>uC�=
��<z閼VY>��=��d�F��=���>��C>}�>B��>�е=�|:���B�ϿnZ���I�ǜ���=j�O��]���T�Dڨ������tԾS�����[�i�n=��>jMN=�>e�׽�q�<�/��\M�2M���rƾ?#ƽE���G�x�"Ȥ�l=��j�=�پ_�<���T�Q��=*ۀ���(���½p^�FU��M��>Y�>��>B�?B!?rZ+?e�?�g�>�}?Ō>Q'? ����w?uR��'? "(?T8&?Tf!?�~�=Pö��2����伂s�[�;�zq=@"�=����T=_0=q=W8*�.�˽(Ž�4غr���>�q>Q�=��>x.�>.,��h_�L�.�����+2�=p�?���AF־�B0�����zO�5�=�Ll�o5:�\4��x۾�"�>�S�>���>�
�~�?>�G����:6V;�r�>�^��YE��rQ�>�����th>�_��j����X׹�.�=��=�&>�,2?�?�O�>�tv���0k�6c��iꊾ�����R>Նk>���>�EW>8��We��B�6-�tܾ�ǽ���=�j�=g4=o�ך�=�z�����=�>��=��=�5�=k�]>��=�C?�6�>C��=ã<��H���ֿ6WnN�H�"��f?[Wӽ���;��;s���Q�k>Hپ���������M:>8V=�p>Fs#�D>��м*����7g�Ôľ� ��á�q8G�kw��1����=H�վ߄�=H8���>��$��hϽABx�o�h�4�Yj ?r�;�?�$?ax>�?��>�7>�P�+?p��>,u?M$�=%��>}	��eR?�?��(?9�?�|&=�G��4K�-�<>��=x��=���=h�=	�<q�>��>�=��+=9J8�k*&�����
��,5=��o=˪h=@��=���c�2=��@��0���񾲾==�;>"�Ծ����_�*@�Ϧ���>>'��nC���ʾT��.×�EC�>!�1=��<��=�Q��`l=���=�E>�2��w�(���=ȭ��Y|��J�ٕ=]VP=�䋻i��=��=�m�����>�rL?�^�>�G�<qt
�9�s���]���¾�za��@�>z��>��L>b��=f`x��B��_���������F�<�k<>ŏ��L�>.�=ȣ�=�Cf=O<�%!>����8�>�>c0n>F�%>�X:>L�����>w�<�6���\��"1���n�.��:D彛��m����=����5>U�ξ_�=p@���
�>���=��=�H ��$���Q�rT�N.Ҿ�h���_����*dǾ-};�����3�9�Q�Z4˾����þ[�D��m���<�#�=��@X��.?�		>znƼ�	�>���>�$?��>Jы>��?2�{>�8�>O�7���>�陾B��><	?��?l��>Q��>�qm�@>="*�=ݍ��e�p=�}�<�u=32���sf=^{>'v�<��=n=�1���"��ܙ��y4=~xۻ��l����=}�R>B ��}0����8�<�j�>Q?������վU,��P<`>!9��f���y��k�¾`$����=f�>�"�>�A>:�J�f~=>���:�Z�=��P=��k>J�ｔ�3��\l>PhG=W�=�`����;E �
��H>����9<�>A^?4�c?�y,?껾ح���y�j�.��Bν�.�ձ�=6M�>SPV>%4��.)��7���ܾ���!K���]��{T>��A;z�}>1h+>��G=�>���˵>���E�@>��;7��>*Ά>tW�>NS�>�w�<MdQ����f��B���7澧�Y޼<�z	=|M��x�׽,ߊ� o�>�&�c���)S�z��>��,=�u�=J�b>�o�>{�>�ـ��}�摇=�j��}!��)O��̜Ѿ�tn���:50>n�ɾ��=�����<��վ�-w���h���sT��e?oo�>p1/>F8�>�'?Qv?��+?*��<��>u;>�g?�V�=�9?���=^�?W�'?ϥ?���>9&P�0���0���(ɼ�ýH:�=sY�=2\>uʈ=���=�q=�F�~�������:I�U�>�=�/>ʾ=N��=
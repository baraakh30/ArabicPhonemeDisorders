`  �   9!�>)B�B���b��b�X���i>ۡ���?��F�>�l�sš>]%�>R.�_�I�i���I0
��PX?|��?�}7?*)?���M�� y���Ӵ>���nd>��==f�����(?��>e�y�fs��7�V��>3e�?���?��e?�����`Ͽ�������������>XC�=GX/>X}ѽ1��=�d=�B<�ِ���5>"I�>U�>�*�>�>>�I)>�->����%��R���̏���6����A����zK��M����
�I���'Ͼ����4��0�r7@��n"��'����;�a>�&?/ú>�m�>=x��j>aFf��f���D�0�>��7�nʍ��@�eC���9��������^���Q<����|�>7�*>�7�=��?�%�9�eѼ>?����d>p3�>H�>�>r�>��=Uv$�k���"\=�4>S�><�V������ԙ@����,0>��E?n>W��i�����Ǒ�<���G�>?��#>�<��ᒿ[�e�� ?�ǃ<�X��5N���x.�R֏>�8�>��=��=K8���b��5ӽ��=���>�<�=��g���Ln7�c�%>`?���ME��>�+)?�|?�V8?k�=�R�>S�=Y��>��>��^>k�= ��>ԕ�>��@?��<?t��>D�y=��V��9�==c���5����������m-��ﳽ����K=�=P�<���<�û����vh���(=�^?��/?��>��>�[�SiD��>M�ف=��u>U��=6xc>uԦ>��>aH�>��>�C>�4�=,�þ��f�>z6�>

��䇿�J�M_�>�.>�y�?��I?�ƽ��8>�e>TMu��>,j?-?�z?���>w�+����H�ݿ�A��x�%0�<;��k�>�K���C��Xx<^���%���;U�>(ɳ>�/�>ܗ@>�Ľ=�9!>��>�6'>� ��x`�<�g�6�
=�*5=UE�=�����<*Ұ��o`�f�ʽ�ٽ{����Ǵ�@=E�T�[���<�I?�;?�S�������=¢���� �o�	?��	?a�
?=M�=��>m�%���6��2�V�)���>k�^?n>?�	��F>�~��!�)�pz�>7s�>�!X>�bW��TU=�Ͼ���=&4�>��(?�̖>��W�X�xkO�L�]��
�>������?<�a?T���>W���8�f�C�?+�w�>}0��詽�����z<��b������ž��	/~>�>�ɓ?�1��@E�F��������A���A����>X>
=�߻2p���.ӾP	&��T��$�C�[>!��>55>B��>N�?t8?��b?�G?��?F��L?�E���?X��>�{F?yP.?;j?K#x>ז�=�����娾퍕���߾�S;;u��=�P�>l�`>��9>��;����<E�=K�N<+h{=�4 =R�S>E=[�A=W�׼�T}=���>�U	?��$?��<���=&{�=����&=Ü��i�>8�p��,��)�=*P�>���>^�?7��>��K<0˾z׾6���=0=x�4?v�K?1{�>�>ļ��z�m1�T+3�s�t>~]>�l��ȑd�NZ��r�������->��+>�΅=��P>��Z?PK?D�?m�B�����*"�z�#����>���BA��=Μp>�H��i�)��ui��Nd����Xﳽ�v�;���>�tI>���Z���>t�|=r9����̽Mv��[r�=t��>i0>;'?���>��N=^W�t��@L(?��e;�9���+��u辁�>^̈>�v��_?6��=��c��M��E�?V>Vk�?_��?돆?*c��PR���"?�`�>M=(*�>���#�u�E����ˈ>���=i̲�}&�SC?��w����>��̽~�� ���>.<�/dʿ��q�0Si�����_���3����+��\��~���|e�ZԈ��%���Ry�aj=Z/m;Ϳ޽hU��5��ΐ���?NӍ?i,��Ȅ��2]�i1ǾlH����p>��i�"d���ľ��ù����5��]���Y�~)�_RѾG�F>
��ߚ��� p���z���>���>�F#?(팾~��ʻ׾+-|�I�(>M.�>�*�}����q��G�P�^�p?�&+?�6վ�4����*>��t��$#?�\��aE�=b���شD�>t�/?�=*?�i�����������*�> �?�P�?�D?<��H�?�oS�ʽ[?S�?�K�>�_�vg ��0� �?x�6?�	�>�Fﾝ���g�	��?�>��Y?�gq�f�5>Q��>Sѭ>�W��9��4�� ��T�1�}F>�;�~D���T��0�`���po�>E�W>4Ok������2�>��Ѿ7,���k
��AC�Ae�FU\>���>���w��=L~T>�U>�I3��6ˍ�VU��Z�?6G�?cL>?U?��#��)�f�߽�7�>�0�>�;0>]�=�b��AX/? ��>k�辇2��8��gE?4��?]
 @�}?��w�]`�ᳰ���Ǿ�ԯ�~b><(>\O]>��7����=��!>I�m=�@��pl/>N��>��>,{|>'x/>��>Z�=y7���d����ӑ��=U�Y7��1辙�K����Ll��@��K3ξm������;.�-�ƽ1 j�K��Z�<a<�j��=q��>yv�>�2~>�䓼R�=�2��J,���ʾ����?M�Ǉ�,��I���f�����#p������ꌽze�y,�>H�>me'>���>�b��x0�_+�>C�=;5B�<��>KQr>�?>	괼��>D4 >o�>dn">�G�=!�=g�y���~��A>�u�w�}ٻ=��@?P��x0�����+��IǾ0?I>�o?��>>�q%����6i���2�>�:�W�|�\�h��6�}т>ȶ�>j��=�)"=�������T��X��=�J>|� =�,˽񺓾m$���u=>�>�&׾c�=:@x>��(?�Fw?n6?��=�y�>��c>�n�>���=GO>6�T>`r�>��?�w9?�"1?#�>�j�=�^�l�=$�;=m�>���^�>)�� �伀-����<��,�x(E=-Am=��<V4b=B�B=�u�����;��<A�
?��<?vh�>ܟ�>� F�R�C�U[�,��<a�>�':��p>̿�>���>{>��h>�3�=�z�A���8��fX�>�6�>�������?�fZ>e+�j�?�Oj?�R9=08v=�JZ>ږ>b��=�� ?�!?��>t�>&�ý����lӿ�$��!��킽RS�0�;z�<�*�M�e$J��-����_��<�\>O�>�p>8E> �>�13>�S�>}=G>��=)�=R��;h;�2F�W}M= �8nG<�Q�i���LƼ���R����I��>��*��ټ��?d>?�������8�=����J�M$?�jj>nv�>�2=�i�>�ﾘo�55B��z.���>iA�?���>@A���-a=��0�V��}�P>�?8Z�>e`�����`�nɊ=;D	?3c!?���>?z�<��X��`O�9&��=?F��;[�ƶ�?�n?B��߾5�5��F�8��Ž-���N�{�߾i)�;�4���־D�����d��B�=n�?�D�?xU�*��@���m�������ʽ%!+�lT��1s\>��=�]T��&Ͼ�z���v�ԋ^���>�Z�>D�=-K���E?8�?EQ]?[/?��?�M���/?��>�O?h&>X?Xb[?q�?h��=�5ܽI�z�Y���f(�����ޭֽ�'y��,�=��G>|L�>�DU=!1�=W�<>cv>�+�3R�;�b>>��=��=Ͳ>>��>p��=R�?��%?����<ʬ�����*��U�S�&��=�f>+�ͽ=�Y��Y0=�k>��>��$?f��>݉�<��۾hȾ��D�=�.$?�(A?':�>��󼇺�=b�����GWڻ�^>�t�������ı��@�ǽmR>��e>�E�<��u>�OL?/3Y?��a?�=���b�=��6T�/h>�T��j?>���>�&>�wǾ��&��X���O��EC�ݓ>�R��+ƽp�>r�4>�(��& �m0�>��߼��Z㵼���<y�<��S�>�s�>z��>�Y>>�������Y��Z^0?`��%��i�;�'���M� m�> �&>2[˾�Y?�%ܾ������{0پ��`?֦�?I��?*�a?����ə��\�>��?3��v�>\�־�?S�}!����>�s������m�F�>F z>��>R���h�� u�����&lſ�Z�A.��O�Gо(X����׽�@�5נ�k?Z����󴢾�U�A�r=�z�U��,���y�վ!!���5�?!�?�}��G��+bm�?*�ϧ��CI>oh��q�Ͼ�*���{�����w��&��?���)7���"�cH����>�	�j����r��e�MZ�k��>��&?͗�-[��m��Z�2=��=K��=<���֟��:�]�1S?�?E?q=���) �*��=�*�=�ݷ>���>Ѕ�(hk����U�\>��D?W?�f��������{�	#N>�o�?>��?�i?w�>#fH�(�1����;x/_?��n>�>�>u��=�%����W�>?�B]?~I�>� ��
��$�.���>��?Q'�����=b) ?Zx�>{-x������Լӷ�av=��L�t<�`�D�������=m�h>��>�[���o�bV>�6��j����d���Tw�쫌>#�>�V��'I=�&	>7lK>J@6�N1@������ߟ��c]?H��?�D6?-]:?3���+�e�I�`=�6�=�[B����>�j�>=�ݽ ��>��?�:���D��<>����>���?1M�?xAk?�t��#Ƴ�u%��?��������@=�� >�υ>����v�=4se=t5a=ϖx��8>�7�>��{>�}>T�A>U�)>�" >���2��(�����h9f�_��龃܂���!��R���� ����������4o��B����}��&���@ �|{>�"�&w"���?���>x�o>
y<�ݿ=��p�e,󾒑8=��ʾM�'�& �\��Zo�D�����������;}��H�� ��ʛ�>+�=�10>N?w�%=FD=�Y>�pZ>|��=妳=�7m>�18>g�>h>R)>׾$=���=�>T�=H1������47�>�G��2�l�C?�,S������2��1ؾ�_��9�}>��?2�L>�(�����ˠt�4��>��;��a��_Ľ����;�>�J�>Rg�=�t���I�,|��O�����=#�>@f>���9���ۖ�Jg�=�A�> �Ӿ���=\t>p�(?��w?�L5?���=�}�>��\>n1�>7��=�P>��N>��>hq?\\8?_1?���>C�=��_�m;=�H=k�>���L������~�i4$�B��<M�2�I=��{=�%<Wg=%�?=d���-�I;or=�e?�'?�y�>�>e���-�Zu�� �<��>\H>�a�>ٹ>�(�>��?��>�H>�1�ƾ�{�>t�>�Tk��S���}�f>�->f�?5�Y?7>�M�};i�(>p �>���>�)�>AP.?��i>�>�NA�u��v�ӿ��
����Z��=���<�6y=w>��4��Ĥ0<��ƽ�֚��u�ɉ	>�*p>8�y>jpV>���=�=�?1yL=vg+=ֳZ=�W���,=��������o�<�%�=��4��V>�۽m?�;��0���"�ɺ{�=H�q=��?��3?��|�ؾB�=j��8(�: ?Y�?^3�>QC>Bk�>�����LS���CUn����=@iN?��?��~<��>�0����VS�>ؒ�>}�=4�۽>��V�(�a<�j�>e�E?~N���4��fE��ts�K��]�>D�<E�q����?�V?��þ{�o���2���2�+&��I�>��M����޾�~�	z���a��\���q���@?>�?�<�?�׶���S�zyL��A���Yw�"�r<�>�4=�Y�>��>z6�ꌧ�^�(�X�X`H��q�>d�>��6>��>2�:?E�L?30*?���>/g
?B��Z�>���:@?����tF?D>?��>?�*�>1�8>��]�����k��5��B�=*Z�;� >�6y=��f>���\q��>
�>�������H2>��~�n��=��=��3>Q�V��?%$?�����=��,��7G�,g;=Lb�=K��>
.I��㽸��;E�>e� ?"q7?���>K};9��N�従��6�<�7?83?�r�>�F���="��+L����>X��>��9�2ק�*�žŃ�-_�i�>ϙm>1K��a�l>��w?ń'?F>�>;�,�+N��AV���d>�1(����=���>|0+<���x��9B]�>�h��%����=s�0�|S�vct>�Q�>����L>H�>=:ƽӇ�����A����2�< �>.Z�>��?$��<�\>M�	�?}?1��%��@���{��N�ྦj�>D�>������?�[j�D_��̵�2�,�i�$=�8�?�'�?�܄?�3���z����|>2�>�N>o8�=C�p�'�,�>	�q�>�g>ꆄ�M9ɾ,�<|)>MՕ>4ҍ�;�ȾA�;��T���[�f��=��.A���S>�n�پ����Ԛ��X��aD�:U��0��f���p��o"�1Z@�#=���� ������?� �?�8>Ay߽"Z���\���E�Z��=���0�����p�˽XF����Ⱦ(%��s�޾� 6��� �Af�����=�������΃��k���'>2г>w��>8S�g���Q��oo����O>��K>��,�����񝝿�/��j?�>���D�1��6����=�n?�R�>���=�x��!y�����<��0?�<�>�bj=`�������;B����?���?vx?>�P����f��<��U?�f�>p��>k���� .���:5?/_?��>�D��Z�w���+�>
�>9_e?a�r�-y�=s�>�?�ʼ���$�1�=�&���2<��-<Ŭp:�	E�͊�}��^�>e~E>��C>�ϕ�E�6�/��>K���n���r^�c
'�vu�=E"�:XA?d�C��@�(Q�=q��>-[.�����!��R�9��-K?3��?�o]?]�"?�n�9� �6�+��z�>�˽>r�q>`T��Tu?^�>����囿:��1?, @G�@_�k?���ϣ�E������ŋþ��=��<��=^j�Uk�=mr�=��=�{�b�_>_��>�'�>pԢ>bq>>]��= �=@���r�)�k'��D��92�����)�,���\W$�Q�%���dy��� ���ԃ��� �5_��o�8�S��&���Ǣ��C�=�գ>��>)�>`>��@=�<ͽ�5�U]�<��˾��&�v}��������s��!y��:���\~����ս��ľ���>�9=�ǐ=�y?�~=M���Q`�>�w<6�J>���>��>�'�>v$�>Sz��?->�<�$��F>�=�����R����O�%���=N�B?�����pϾ\�3�E(��Ǿ���>Ձ?�3>��;�-�����o��.�>��=9��F��������|>D�>�Yq=]ȝ=���{W��掽^_�=2_>n��=�D��PC��ѵ$� ��=��?��D�Wy��K�<=�	,?���?,�!? ɼí>2\;>�� >zY�>�{G>��= ��>P�>�D?��A?�z?��=TU�H,*>t5u=�O�
Xּ!I�	胾b� �QJs=�'���<샸��`>�芼� =�����<!sK=��?��-?���>���>�����5��!e�Z�Ƚ�lQ>�V>���>�Y�>8��>x��>�C�>8Q�=�6�=ܝ������K��>��>l�e�B�����b�m_Z=�n>�S�?�![?:P ����j�Y>�<��>L��>�N>?�u�>���>3]J<���߿��$3!�t0���/���=ܤG���j�H-b=������"�~=�f�>W��>0�}>�3>�4�=̞�=�>�)>�U!=n�!="B����;�	�<|m�=FA���'�=�S���ٕ��-ݽ+�佹L����VV������<�<'%?��?�{ս��i�Ტ<a�� �3����>\�>�$�>dc�k9�>)���i��6%�����>3�Z?�?$? �I09>�V���S5�<�?7A�>�)�>ۿ����@�$�¾�!�����>��?�>}kg���D��)H��Ͼ鯞>&֐=�M۽�5�?��A?��¾�6�rcA���)�N���ɷ=<�e�I�)�m%ľ�p�h�$��� �tݾ-�\���A>�L�>�ә?�9:�y ����7�p����&���5��>t'}��>7�d>�Ƃ��w¾%+����<4�_6V>%W�>\��=��>�K?ת5?��4?Q�>��6?�S���==?�K>�]k?�ʊ�ftw?�e?��S?�&?�f>cK뼜����ȼ�������h���&=��>��>�9Q>�E>��>C�d=q�>*&=< ���EW=*��=���=��={Q>z?��%?Tw=�.>�8�=]��!X=i�M���n>�t>��&�^��=�
[>���>�K?��>�޺=�վ�(⾝n���5=L�C?�L?]��>؇<3L{=&����js�
�(�b5�>gf����?о
Ѿ16���s>��(>Ù;���>Q�j?+�5?�?�!�=���ӫ?��*�#y=u̽��5>��u>�='þG��P'��f�҉*�R��<I�/�lt��G��=�=�>�i���X=H1�>�"�<�w���V=�ͳ>P�����>Q8?12?���=x��f�&�8��%4?��ߡ ���۾�q�p����=���>����?aڊ�]p�鍹�9W����=7��?���?��?�L�1�����>��>�+d>:�=�J�����l�B�3g>�[>���S���ژ=��=���>!sL����ݯ�y񓽯�ſ�ׁ�ͳ|���%���˾������;��{;�ţ��Q*=��������넖����<�s����P�R���2��Wv����?��?��`��<����X������}�E�V>:L��/�����������#��e��.H��7&��[S�1QC�<���v>7	�ԥ���q��Օ�~R��Yy/>�?�ڂ�W�U����Į���q:�ۨ���"�7⮿�ܮ�����NHc?C_??�������dj>��>��K?8_�S�?>0���aߣ��@k>��R?�!R?����w���EN}��>>��?*��?��M?��s�HwA��B�X'���?{c�>/;}>�*r�����u�a��*7?��?���>�ܾ��s��@׾�?�`?htY���>z~�>�=�>6������PI6�}�¾�m<E7�=L]����(�k����߭I<�t�>ag>�PZ�����9!�>)B�B���b��b�X���i>ۡ���?��F�>�l�sš>]%�>R.�_�I�i���I0
��PX?|��?�}7?*)?���M�� y���Ӵ>���nd>��==f�����(?��>e�y�fs��7�V��>3e�?���?��e?�����`Ͽ�������������>XC�=GX/>X}ѽ1��=�d=�B<�ِ���5>"I�>U�>�*�>�>>�I)>�->����%��R���̏���6����A����zK��M����
�I���'Ͼ����4��0�r7@��n"��'����;�a>�&?/ú>�m�>=x��j>aFf��f���D�0�>��7�nʍ��@�eC���9��������^���Q<����|�>7�*>�7�=��?�%�9�eѼ>?����d>p3�>H�>�>r�>��=Uv$�k���"\=�4>S�><�V������ԙ@����,0>��E?n>W��i�����Ǒ�<���G�>?��#>�<��ᒿ[�e�� ?�ǃ<�X��5N���x.�R֏>�8�>��=��=K8���b��5ӽ��=���>�<�=��g���Ln7�c�%>`?���ME��>�+)?�|?�V8?k�=�R�>S�=Y��>��>��^>k�= ��>ԕ�>��@?��<?t��>D�y=��V��9�==c���5����������m-��ﳽ����K=�=P�<���<�û����vh���(=�^?��/?��>��>�[�SiD��>M�ف=��u>U��=6xc>uԦ>��>aH�>��>�C>�4�=,�þ��f�>z6�>

��䇿�J�M_�>�.>�y�?��I?�ƽ��8>�e>TMu��>,j?-?�z?���>w�+����H�ݿ�A��x�%0�<;��k�>�K���C��Xx<^���%���;U�>(ɳ>�/�>ܗ@>�Ľ=�9!>��>�6'>� ��x`�<�g�6�
=�*5=UE�=�����<*Ұ��o`�f�ʽ�ٽ{����Ǵ�@=E�T�[���<�I?�;?�S�������=¢���� �o�	?��	?a�
?=M�=��>m�%���6��2�V�)���>k�^?n>?�	��F>�~��!�)�pz�>7s�>�!X>�bW��TU=�Ͼ���=&4�>��(?�̖>��W�X�xkO�L�]��
�>������?<�a?T���>W���8�f�C�?+�w�>}0��詽�����z<��b������ž��	/~>�>�ɓ?�1��@E�F��������A���A����>X>
=�߻2p���.ӾP	&��T��$�C�[>!��>55>B��>N�?t8?��b?�G?��?F��L?�E���?X��>�{F?yP.?;j?K#x>ז�=�����娾퍕���߾�S;;u��=�P�>l�`>��9>��;����<E�=K�N<+h{=�4 =R�S>E=[�A=W�׼�T}=���>�U	?��$?��<���=&{�=����&=Ü��i�>8�p��,��)�=*P�>���>^�?7��>��K<0˾z׾6���=0=x�4?v�K?1{�>�>ļ��z�m1�T+3�s�t>~]>�l��ȑd�NZ��r�������->��+>�΅=��P>��Z?PK?D�?m�B�����*"�z�#����>���BA��=Μp>�H��i�)��ui��Nd����Xﳽ�v�;���>�tI>���Z���>t�|=r9����̽Mv��[r�=t��>i0>;'?���>��N=^W�t��@L(?��e;�9���+��u辁�>^̈>�v��_?6��=��c��M��E�?V>Vk�?_��?돆?*c��PR���"?�`�>M=(*�>���#�u�E����ˈ>���=i̲�}&�SC?��w����>��̽~�� ���>.<�/dʿ��q�0Si�����_���3����+��\��~���|e�ZԈ��%���Ry�aj=Z/m;Ϳ޽hU��5��ΐ���?NӍ?i,��Ȅ��2]�i1ǾlH����p>��i�"d���ľ��ù����5��]���Y�~)�_RѾG�F>
��ߚ��� p���z���>���>�F#?(팾~��ʻ׾+-|�I�(>M.�>�*�}����q��G�P�^�p?�&+?�6վ�4����*>��t��$#?�\��aE�=b���شD�>t�/?�=*?�i�����������*�> �?�P�?�D?<��H�?�oS�ʽ[?S�?�K�>�_�vg ��0� �?x�6?�	�>�Fﾝ���g�	��?�>��Y?�gq�f�5>Q��>Sѭ>�W��9��4�� ��T�1�}F>�;�~D���T��0�`���po�>E�W>4Ok�����~��>����p�jG��V����=c�=���>1���;7>�`�>���>f\�����j���4��jrF?v��?�@e? o"??���p鈾f��%<6=a	T>6-�>R�<C0��VG�>O6�>��	���z���jB?3y�?T��?lr>?����#�ȿ���7����̾Y�=��P=�� >5�ؽ���=�zj>��=��=��k>���>	�R>f�>!�,>ܢ�=�>�"{��T��������͵?��5&�����.>ҽ#�� .�y������־b��G��󻼆�t	[���<��_�%�>n��>`L�>C��>���>9o_>ճ��59�\a!��*E�ĕ7�|]�pn�>��KR>���=\D�����J+2�y���/?�9�<r�=C"?>0��ᶢ=�^�>�+�=�2m=���>��=��<>m�9=:�5>�g%>�>��N=�)X>���="���USI�뀿y�H���>�_?i�=R�u�ZLJ���(�����#�?��?�tA>��ߗ�ʇ�4�?�UӼ:Ũ�M�Z�.m���>'�?��!>��������O��B�=v'> �>��!>G?ٽ8zʾ��D��>U �>{�Ծ�>D�s>5�"?`΀?�/6?s]=YM�>#i�>_+�>'�=��$>��=>�i|>]�?�x8?f0?�{�>ԣ�=L�S�$r�=8pK=�]@�~���)
��׆��k��C4�<L���TC=E��<N�8K�==���=��U�%�u=��M=Pd?#46?�՞>a��>n�R�o-T��>��|>^��>�.|�y 0?���>}� ?�\b>��F>h���D���q��7zB�F��>v[�;����7��o�9��?v�6=2+�?��?�s��ٍ��ʪ�>��@=V�)?ny?J�?�k7>�ܓ>온����ſv�����ʭ�x�
��Q4�[������qa�����>�y��#>?�>�_�>���>n� >��=g�o>�%�>���>�g�=�>����>݇<��ؼ�LB��a>v���\��:~= 6ý�ż�Y�pB�2T<��y�=ˎü��>?O8?(�>)}�=P�<F�AN����>��>�V�>42>��ӽ����1b���L�>i����?�\?�W�> �����=ʹ���=�`�>�5B>�0�>A7N�MlS��®�t��>�V�>��?��>n�?���w�N����q ��އ>*��=�:;z��?w�h? ๾�4G��R�fN���@�Op�=�ϲ�������;�y.�T,�v������d���">�D�>���?U����#<>笙�����W���v��z�ֻH�S=�\�>ب��=�h�����}�|���
����=�|�>B�=�I�>*�;?9~?;�Y?z�>� ?�!��N�>շ>�9�>E�>Ѝ6?�N�>�q?�O>0x>��,��(3���#����x25=w|�<��=#��=.�F>h��o��7�<=�]E���A��dE=�O�<�L��|�<�H�=E��=8C>0�?ݩ?@��=E.T�����)�㽻F�=1��={Ʈ=��=�E�ͯ����@>,9�>h>m?���>��d��y(�����B/�>2�?@?�� ?Nge����<�{����i�=�0�>�Z��>ֽ��"�D[��R��m�>� =S���gNL>�(�?�0?q�p?�2>Z1[�AJ�+�8���׽`u����>��=��Y>���C��Ye�3�O�ۆ:��G�<�Y��1)D�J)��ا�>U�m;-W����>��K=�{��J/<��>t`��c(�>��N>��>y���5��؛��V6�\�7?ϧJ�(����󵾂�f�[=�^?�i�->�dl��?^��3q��
Σ�h,���>�H�?@��?i�T?i���'��yɐ>��>C�=9@�����[ҽ忀���>4s�=�'��e澸2�<j��>���>1�<��z�����޽�<���A��@��d�����^�ϾΙ����'�Tw��� �w�پ����
�M��Y�s�dMv�("��Z���L��?���?<��;�f���D�SU�2'��i>k�#��e��'#ľC�?����&��	\���	�E��7�4������>���9G��&�Z��=�u�T>g��>B�'?�/澷2����>x�p>ͥ>|L�M���ݓ���U��_?��6?���ې
��k�g�>ӂ$?v(=�t.>K���l�u�>1��>HJM?	TW�����S3��k��<ŷ?E��?n�L?<�;�[�&�	$�S����?���>�kG?�H2��8��I=��1?�W?Z��>Ð��2��3�C�޹?��(?ҡ&�D+>	��>_�]>ÿ�=8���9���Xq��W�>���=#���z�",���tM>s��>�g�>����¾�;�>ӣ���䃿����.پo�꽖�Y>��>�3�����>���>ۓ�>qc�|$���7��5~K�Y�H?>w�?,�{?}F?E8������w���>�$R?y����>���;eA�=��'?]վ�_}���\V'?C��?J��?��a?�x� �п, ��]�����0c>G >T:m;l�%��g=G��E9=5���R5>�En>�NI>�ut>Ć>�Z� $>������/��,Ά�I)��`��!�夈�A.�st��A
�3n��^ľ���G "�6�⼃��A�<F���!��D�>E,�>�>Z�?�ǩ>���=�E���UE��o��4f��,����žC��F]���S�Ah�8K�P�`����aL?�[�����>��2�c�A=?:�>�)�=t�9��>�xI=��]> �=߾>>(V>e�W>�
�=w�>��>%S|�[�d�F.������.S�>n�(?�c>�M����7��/��Й5����>6�!?���=+�'�^1��Rݥ����>�>W.��!�h=ۿ��I�=�2?g?�G.��1>�Ǿ�ȼb�>R�>TY=%쁽�zӾv�ž���<�1�>{�Ⱦ�U>ɭ=>C�#?@�{?�,?j������>@�m>�@>���=��=1O>��>�6
?�3?bK.?��>i*�=rV1�DY�=�1�=�틾���*N�k�V��}�щ��yH����}��<)�#��>y�8>��R=��=SO9=s� ?�6?�k
?��>툯��J��:��y����>k僽̼>~�>�1�>���>]=�>,>s=v���.������ν>�>�6Q�,���+＄p>��=mh?4_/?�8�����~Al>R#>i�>��	?��?�>�/s=?���z���ſ�������;�N��jz��wD�^�p=��������Mw�t��=t�>�V�>�x]>^Ei>e�F<O�L>;�>�H>�V1����=M$��^��=�S=˪=��*=|J���<}㢽!X���2��p|��=s<ܖ�= �o���?��?��k>�]>���g=��V���?�m�>���>p��>��=��] M�0Q7�gÇ�pҞ>nV?:�>;*�1`J>����G�tb�>X�>94�=�(&>��)��,Y��ua>c[�>2(?�iI>Z<ý}+V�X>}�MS���8�>�ɂ=12޽qs�?gKd?m���n3z�!���F�YU�L`�=�\���4{�;��e!$���2�X�辕��~E����=~��>�ڠ?��x����=�۸��e��)���W�����E=�vm=7}�>h�$>���<��ȳ��G���D���<�#�>qȤ=���>oZ ?q�?(I`?�8?=?5'���?ܤy=R��>/|�>�5?��?��?�&�>a�a>�*�<����Y�(����<˻��_�=��>�3>�d���s=l�q=�l�<j&I�Ӕ	��y*<#�<�0=<`�=���=@�>w0??�?��=O ��f>�C�ݾ1��ƽ��ӽ�W�	�˾��n�L��=T��>��@?o�?�>��������u����@>�&�>��:?fB�>y����A��lk��>��Gj>I9�>s�ؾ	t�N��F'
�wT�q+w>�r>r��<$�>9y?r\?)R?d<��/�LlT�����3�@0M>*��>b6)>p��=]�>�@�)�X�:�K�E��\���m_&��Y�<���=/u>>V2\>N�ļ�>{���=������=�]=�Q�>���>�]�>j&�=_|�<Mɕ�ͭ�IN?��U켾�1=�i�=���>�E���h>�z�/�>��y��{����aH��s�>�%�? ��?/�N?J2Y�Tc��ߓ>/mR>�,o>oLs���l�Ȑ����K=$��=͐��C����ȾV�X>c��>6m�>������zQ��wE�7���-=�%pf�Sپ�5��`Ⱦ�ף�-��:5��Hi�ٚ���YM�\��0	��>���`\��M�	2��r-���;�?�r�?�ذ�h�ٽ�&6�ظ�O�P�y�Z>�ڽ�O�;鹾~�U1��a~��<������>:&���(�]")�X�>dj�<������-��Ir���P�8?'�>����?�:���iI>��>�
=;"��S���ע�om;�R?-f'?0~�^V-��z={�>�B�>��>���=��쥽�S�>��3?�?���,���e��m�\�t)�?���?oP?�ڇ��*���(����"�?�?Y�?a�<�Ƚ�tI���XX?L��?��A?����Fx�(�6���>�?vl��r�>��?A	>�h��p��_xv��)������->*�.�Q���QF��L��ʶ=���>8�|>>�s����~��>����p�jG��V����=c�=���>1���;7>�`�>���>f\�����j���4��jrF?v��?�@e? o"??���p鈾f��%<6=a	T>6-�>R�<C0��VG�>O6�>��	���z���jB?3y�?T��?lr>?����#�ȿ���7����̾Y�=��P=�� >5�ؽ���=�zj>��=��=��k>���>	�R>f�>!�,>ܢ�=�>�"{��T��������͵?��5&�����.>ҽ#�� .�y������־b��G��󻼆�t	[���<��_�%�>n��>`L�>C��>���>9o_>ճ��59�\a!��*E�ĕ7�|]�pn�>��KR>���=\D�����J+2�y���/?�9�<r�=C"?>0��ᶢ=�^�>�+�=�2m=���>��=��<>m�9=:�5>�g%>�>��N=�)X>���="���USI�뀿y�H���>�_?i�=R�u�ZLJ���(�����#�?��?�tA>��ߗ�ʇ�4�?�UӼ:Ũ�M�Z�.m���>'�?��!>��������O��B�=v'> �>��!>G?ٽ8zʾ��D��>U �>{�Ծ�>D�s>5�"?`΀?�/6?s]=YM�>#i�>_+�>'�=��$>��=>�i|>]�?�x8?f0?�{�>ԣ�=L�S�$r�=8pK=�]@�~���)
��׆��k��C4�<L���TC=E��<N�8K�==���=��U�%�u=��M=Pd?#46?�՞>a��>n�R�o-T��>��|>^��>�.|�y 0?���>}� ?�\b>��F>h���D���q��7zB�F��>v[�;����7��o�9��?v�6=2+�?��?�s��ٍ��ʪ�>��@=V�)?ny?J�?�k7>�ܓ>온����ſv�����ʭ�x�
��Q4�[������qa�����>�y��#>?�>�_�>���>n� >��=g�o>�%�>���>�g�=�>����>݇<��ؼ�LB��a>v���\��:~= 6ý�ż�Y�pB�2T<��y�=ˎü��>?O8?(�>)}�=P�<F�AN����>��>�V�>42>��ӽ����1b���L�>i����?�\?�W�> �����=ʹ���=�`�>�5B>�0�>A7N�MlS��®�t��>�V�>��?��>n�?���w�N����q ��އ>*��=�:;z��?w�h? ๾�4G��R�fN���@�Op�=�ϲ�������;�y.�T,�v������d���">�D�>���?U����#<>笙�����W���v��z�ֻH�S=�\�>ب��=�h�����}�|���
����=�|�>B�=�I�>*�;?9~?;�Y?z�>� ?�!��N�>շ>�9�>E�>Ѝ6?�N�>�q?�O>0x>��,��(3���#����x25=w|�<��=#��=.�F>h��o��7�<=�]E���A��dE=�O�<�L��|�<�H�=E��=8C>0�?ݩ?@��=E.T�����)�㽻F�=1��={Ʈ=��=�E�ͯ����@>,9�>h>m?���>��d��y(�����B/�>2�?@?�� ?Nge����<�{����i�=�0�>�Z��>ֽ��"�D[��R��m�>� =S���gNL>�(�?�0?q�p?�2>Z1[�AJ�+�8���׽`u����>��=��Y>���C��Ye�3�O�ۆ:��G�<�Y��1)D�J)��ا�>U�m;-W����>��K=�{��J/<��>t`��c(�>��N>��>y���5��؛��V6�\�7?ϧJ�(����󵾂�f�[=�^?�i�->�dl��?^��3q��
Σ�h,���>�H�?@��?i�T?i���'��yɐ>��>C�=9@�����[ҽ忀���>4s�=�'��e澸2�<j��>���>1�<��z�����޽�<���A��@��d�����^�ϾΙ����'�Tw��� �w�پ����
�M��Y�s�dMv�("��Z���L��?���?<��;�f���D�SU�2'��i>k�#��e��'#ľC�?����&��	\���	�E��7�4������>���9G��&�Z��=�u�T>g��>B�'?�/澷2����>x�p>ͥ>|L�M���ݓ���U��_?��6?���ې
��k�g�>ӂ$?v(=�t.>K���l�u�>1��>HJM?	TW�����S3��k��<ŷ?E��?n�L?<�;�[�&�	$�S����?���>�kG?�H2��8��I=��1?�W?Z��>Ð��2��3�C�޹?��(?ҡ&�D+>	��>_�]>ÿ�=8���9���Xq��W�>���=#���z�",���tM>s��>�g�>����¾�_?����Z�w��I�H� �P`�>��&>Δ�>oݕ�~�鹊~�>���>�)��򄿛���f�}���p?ā�?��v?A(1?�+�N0ʾ	���>��?�0/����<�uA�v?�>�?/����U����j�?�E�?��?��[?�`��M�ԿÜ����������>�g�=b�(>I��lHh=\��=/�7<���<��=}�>��T>Y�>�)k>��8=ʥS>>��w;!��W�����)�5�ud�.�!st�S��5s�1\�Q�������A�Y����e�P<��(����-uw<UI5��ɗ>Ea�>�x�>�P�>0Yd>R0�>0ө��@���g�������
��O̾z��ѹ����½�I;@ݏ�Y��</6���_?Z�Ѽ�/I=���>|�ܽ¯)=e�>�d>z>i�>5�<=�`�>$1�<Kj�=�tI>mt>���=���>���<t����Ny���F�0�.>|�+?WAǽ
馾J]6�{!���_�>�?�S>� ��ו���`��Y�>w�� V�J,	���X���V>(�?q�>��	���)����z=��>+F�>?�&>�**�M�׾)���;>P�>3(��'g�=�W>�p"?�{?��4?��W��?C>���>��>
�<��>�u>(g�>�?�:?p�/?��
?.��=T�j5V>k&="E���X��S��T���s��{Aƽ�H�������<�5�L��=�>��$>�O=���>��2?���>7��>�c���A��'a�a.�� a�g�q�78>�J>�?�[�>L?� �>}�=�3k�Ѩƾʜ�>�d&>�[���q�f��=�ߙ=��=x�Q?�!?�8$��e罀�=3�Q>�sx>�	?Br?�Ly>$��P����H��z����	�8�*�����]���h�&�YY������ � ?7��H�|��Ϩ�@�=N�=$�W>��">���>e=V�0�>kB>�_f�1��<-�c�P��r�J���=�=:�½��e�!�)��qὒ|�����������1=����d*?I�>Y�=��M�q	f�e:�'����/?��?�\?W�A?Br/>�����&���g�؀¾��E>��Z?�b!?������U=-��eqȾM?)]�>zB�>h�>�����D�|�=Z?^�!?j3�>D��P4C�1}��;Ž�M�>	�=��<��?�;�?�����ʳ�1W(�*A5��qᾐպ< 7��Dk��e׾޲D���8�j���ñ��h�����;��>���?#lL��>%<��ؾu]��VEV�'(.�>�V>da?�iq>r�ݽ�I:��<*�������e��{=<W�>�E���#?�)N?�B?&]?<��>���>Q�T;,�<?�D�<��$?�E�>y��>c�>��>�s<:�>Y�$>����=�4�z��!�ٽ�»�GS�=�!�=m�>[! =ϡ�=֬<�<5�۽L��=�Y=G�ν�j�=��=���=�e>� ?�?�Q�ʅ��G>��ֽ���s�7�Z/���%i�G�zW˽>�ͫ>�<e?`,?��">��ؾFU�D��ҫ�>�>7�C?���>��`=:Z;P!�4�3�Q D>�6�>%o������w-�_�ľ&��;<�>�g�=��j=|nk>��x?rh?wHZ?ISU�]�/��K<��0��S=�0��>��>|�==���o����m�{�b���U�Q������X>,' >1�>�~>�$i>	�,>�Z[��p���I�����=&�����>C�c>�&�>ўt=�'5>��]�g־��D?�a}�;]� c��v���l�>�y��<<-���Z�>[	@��k��-4���.���?m��?�ϼ?4oF?��
�m����p�>�T&>>�>��ì���u��A�X>}�G��ƾ�}�I�Q>�]�>bk?PFj������ ��ѽ���h@���i��C��9i��É��l���]#�i�=�V���Ҿ�p�;Fܾ�6��C�v�
�%[e��ľB$��[��?҆?ʚ���^��:L�O��iד�,G>6�ؽ�.L�����L��=�i��q�I�b3���&��),���&�D!�u�>[G/�����-s��4{�6�=c�?c�!?��P����/�.�E��>�B<=��*>z���]��_'��Ϳ��i�s?��R?�e��f⾒�k��P+=�|?���>��o>�龅1���|�>ѳ?[�S?����!���﵏�J��= ��?���?�U?�C�����$��Q�|&�>�v?��;?�l̽:/��0��B\?tj?]�6?˾�Zw�k�_����>��+?�X��p��>��?#��>�5G�V>�nF���M L��?>��o�G�=X��Lk*���>�E�>B�e>����N9��C�>���ϕp�>�_�P�پ��>�}�=34?�����u<�ʴ>��>ߙ�B|�E3������8�O?���?�u?��??m�/��Ͼ�d��r�>��>G4�=���=������>�c?'%&��@o�7o�q�?���?�� @kU2?��h�"Gӿ�
��Y�����֟�=U%�=��>>* ߽ȭ=n�K=3ؘ��b=��>[��>>o>�;x>¼T>�<>��.>e���n�#��ʤ�ْ��[B�� ����vg��{	��y����ɴ���e���l����Г���G�s���S>�,�U����>w��>���>��>��@>��<�w��s$��2���B��M�,��|ݾ�������`���U=W)F��ʱ������8L?����L�<��>��y�j>G|�>>�g�T��>,�`>�}J>M)l>�MG>h�>�#>�'�="])�����8Z>������oiz�]�C�#��>��?Bq�=4�m���c��:]��'
��~�>.�?�����T�����謹]��>�Y��d����>t�e��=���>G|�=ҥ���=f�������p�>^f�>Y�>�N��㬜�ܳ����=�k�>�{��K>��=�?I~?E�?c�Q<rj>�>�6v>�!f=��x>�5�>�k�>�J?�d&?9�%?V��>���=R�?��l_>�=O}��:N��
>�o���Z#�f[��w޽�32=�}>ov=>�Y>/3�=N�ܽ]�i�#DJ����>c�
?�>?j�?�>�<Ă�kpp��MǾ1rǽ���5�>�b�>V�1?CB&?��+?N�>L�$<�95��||���>���&�:�2�"�7{��Q>,��>pZ?�'a?��=n��4�Ҽ��Ľk�M>��>��?�Q�>�x�=ؔV=���Tvٿ�A ���/ǹ��6�qf�����������=��4�f�����oNd>�{�>�#�>8�>u9�<��m>��?��Z>k�m</�>���
��3�S;�j��EɽG��z���K��.�ˁ@��׽�����V%��M̽$,$�L�7?5ާ>'#=z�n�.��o2ھSt���?�/?t�?N�6?��뼒`�*�n�r���)k~�B��>5�V?�E�>vã�R�>������ �n��>�!�>��ۍ����������?���>q�>����A)��a]������:q>c�E=:����?�J]?���R|v���"�2cH�|�����<�c⽝\[�l/��*���\4��+��Lu��q�s|�=c�>��?N���?��=�[���ؚ��	������eK=:�=U�>�e=>�X,������B�3wϾtL�N��<�(�>Ӽ4�hSD?82.?�?h}?5��>Α�>�Z�=(=!?V>�b3?S+>�a�>}o��fam<��?>?��>_T�=(>�C��\��n`=W�:���d;�8�=��M>EfF�6�����g�y�=���xnk��Җ=Go�<B�C=ۃ�=�o�<xN�>.�>1X�>�[�=%�<R8=Q���[����[��:ƾĀ����3���G��>�t&?
@?}��>�r�<������ł(��$�>�
>��?�?���&Ջ�$S��_ة�%ٶ>��=���8ež�[5�LW���6�����>��=I>U@o>��v?� J?�?)(�=�O�D�X�yI��=���=��>7R�>�=g!�Rz>�q ��`Y�n��̉�"��;�=>4�2>��>�N5>{W>�wp>����=�z���E�	����z>&��>A?%U�>n�=����C��a?��
�C���5�l�>}���I�=N��>ڿ?��>��H?&��>�ϐ�4u���\D�~4v>���?��?�2?�D�=�v��u�7<��=L�<�3�=w�J��!�5#>��>N3c=O���e絾#[&>z��>�ۖ=�q��#L�w����)�K�ȿ�O��i���[��۾c9ɾ6�-�
O�<�"��M����>�}����l8�l�ս9'��hľ���'Ⱦ���?7_�?��/���5�lxM�*���n���N>�}轏�9�J�Ѿv&�4Խ��ݷ�춖���PS��=�k�<��L�>�*��ʐ���_���S��M|<�$ ?��,?Mޯ��=��(E'�@l�>��>Ȇ8> w��ۙ��7���7C��lO?p+M?���4�*��A+�>�hZ?��=�>Y6���-y��H�>�Ze?N2?��Ľ@#��lg��C�k<�=�?.��?�sL?����IF��L��h5�$~?z��>u��>����1�
�BD���"?�Cu?H?���*y�<��/n�>��I?�e��N��>���>�w>�k��&� �#�)=~!����cQ>�ල��Q=��G�FS�nB����>�m^>|}
��ؾ&��>0M�'�N���H���������<>�?���@C>�i>�N>��(�S���̉�S*�D�L?H��?��S?�l8?f����ϟ�����=���>Ӭ>ጯ=/����>���>�^�vr�}�Ț?}H�?���?,[Z?��m�������?������毸=b��=Ӌ�>�u��E�,>g�"��r�	�=v}>�ڥ>:��>
��>s)S>�vv>'3>����o��E������^Ph�J�7�_G־������־l����J� `��Bf��i6�� ��'�bݾ�j�¾+n���,�;�A�>�b�>�`7>U��<��=O��O$1�&麽5�ɾ�5�������쾞sV��а�>a��H��>%C����{����5?Iu!>�Y�>�?�ͺ�ߌ�<�|�>�]->xcl>�	>ևj>\�Q>�|>4��>���>�s9>��1>��н��>�웿�T���t}�P<�r¡>�<?%�&�� �mDy���˾(ޔ��E�=��?@��=oW�W����k��W�>򑃽1���������;�w]>2�>f9>C[���S=$V0�k4���[:B�=/_;�f��~#��R��7�\>F""?����Wk彃X>*�!?���? �2?_!:>u�>䭵=uQ?� �>��4>m^�>ї�>�9?Ha?T�_?~�3?,�E>�2��=Sܼ=�	�5G=l�y=L���3�3�:�]ǔ=m>ḟ;{k�e��;*��=/�⻄�>N��=lc?׵%?'�?'�?�u�5��$�3<�0�<	0�>W��>|n�>��E?��>Bü>d�>�I>�/ٽE�����>�yk>�[/���v�C��G�=��K>�i_?!�_?�B�<����bK}>����iF�>��?51?��?���>3�K>&��g�Ͽ����Z��9��S=~�l�_��_�=�s�<��Ͻ�$���w�=�h>�I�>�>>v�4>�J>�n>��>&�(<e��=h�=*E�^��=Q���k���A�<���=���
~p>��=���=+�p#Ѽ��=ʐ���=z?uo?w�&��4��?�f�;��E����>ͷ�>�C�>���>O��=�n�y�U��mA��G����>h?қ�>&�8�}ʾ=G�/��S:��>CC�>� >�a����^���2A�<��>��?Rc�>�;�DX[�t|o���
��/�>������v�?$	z?`�־��q���0���[��JǼq���y�:�-���M�y��Ȼ��!�(  �5��>|��>�?�fN��o,<>G��4���Fw���ƾ�px=��\����>�٤�\(�.a���&l�Lh!��y��"t*��h>u��=��>l?��?-Yb?B?��?Lm�bf?�W�=�"�><��>/c	?q<?�@�>�֏>���>蹥=�/ͻ4��]����J�<!�ݻ���=#E>y�8>�:0<���<p��<
�*=��0�%>��FF���E<��G=]J�=�[�=6g>."?�?�);nJ0>|H�<18<���?3->�==�(�=�W�$�>��?�?��>���=J��ϗ.�QXž��]=W?�}A?2Ӹ>�#�;P�f>'V��<��M�N>���>�/=m�[�¾Ӿ]��YT�7ݗ>���>-@�=4�>/2�?l�=?��}>+��>�s��u���?e��,����[�0>�(U����?g�t2��u�~��?4�h�2�:Խ��d��%<�1��&��=y�/>"Y>W��>DQJ>�2������#�*CY��3?;�?���>`��>��=p���ي1��I?���d�`�vо)����>��<>���~�?���q�}�����?=�W��>���?p��?�Cd?��C��0���\>04V>�>=�0<&�>����0�3>r��=�vy�B�����;h
]>_Ey>A�ɽ2�ʾ~(��?H�\��
!L�[/P�⾠ ���ľrn��WK�'���q�h��N)"���H��K�����߽� ���T������9nd?Ωh?f;����E��!�{��.C=����R�S��O�*�_k���)پ[+�������@�'�G�
����]>��'�%엿yÁ��;���ѽG�>��5?FȾ�BԾR�.��y�<[U>�a��Ҿ�����7lE��cC?��6?�ݾ0�˾�	���v*>��
?��>��<>�8־��U�y��>�!?=�?�ď��ڊ�9���4���Y�?
��?��??Q�O���A������2?��?���>�����̾(;�0?��9?rƼ>���f���6��>O�[?�HN��cb>���>�@�>Z 𽔷��,&��3��x慼��9>�������Jh��+>�-��=�
�>Ћx>�]�+���33�>Wn��#-���L�'�?�j\v�ӈ�)'?�$����=�Z�>��=i0�����nP��l�̾�x+?� �?�z?�?��뾛�n�>�>��׽U��>���mв�?I�>j��>��۾��������Ho?��?��?͇i?�>��?hϿ�B��;�����>C�= x,>����=�q=g��<�7�<P!�=���>��k>e\w>9X>T�S>Je+>�m��&�1+��{��N�;��z�'�٠^�؟�;`�'�
�������˾۱���Kɽ_n�VXJ��s"�߆j��י���=b,#?�> �>M������=gL��H�����
��/��3�3�,�F��H̾N���n�������=]��j�.��y%*?�=[���>��?�
���ϐ>���>��=�1>�o�<�b>XӁ>�/?@��>���>�$>(�|=�a*=���>������@e�+2��q�>1�\?|ց���8剿&�>�,�̾�D=R�?&xi>�X~�?S��T�y�� ?�"y>a��|��vW�#�>۵�>�I����P=IJ���.�����1�=�{;?�D>�Q���	Ծ��ҽm�M>�8?��q����>O?l?��/?�# ?��u?
�>O�>-������>]��>[N?s�k?��_?���>��j=!,�$��O��������W��WO=��-=����=O����=��=��1��Z�;E8">I�='P%��Z�=��>ƐI?2c?�
?��[�VlZ���s�:�����>�e�>���>rq?g�A?�%?H$�>��>$>6eѾ�7�1F�>C�<>����U��N�����=�CB>�U_?�H$?!J���=B�q���� �<�>5�>3�?u{�>�>�8>�F��S���.G�d.��B4K�q���2�>���Cm� =��ý��`�<�1����=���>�7�>)��=�|�=�R>:[ ?
D>G�D=a�=�G;5~=+g�������D�=�/t�����ݻ�S#{<���i��bϽ�N�wu���	?��?=#D��i��唾d���x��4��>�d�>/
�>X�>���=����b�^�����#�>�k?T9?�1����t="d�<"�>��?�І>� �>��1����{��:�
'�>b�>e�?�X��:9*���l�@Z��yU>�U/=���K�?8T[?��O�����]�$�?�'��1�:�H>�-��G|��ɉ����Q�#�&�N�c���t w�͢>�>'?�?A�O�m�ӻ]m��h�����D4��c�Ҥʽ��>�Z>R���!G����B��^)�j\	��s���}�=ё^>�>M�?�DD?l�Y?p�?��>�G߾7eY>��>G'?��%?�?+;;?��?�ޫ>�S�>	W�=�\�Q��������<4c5�e?=N�}=��a>�G�K;>��= �U���n=��1 ��:�<�.��MĽ�T���5>
u?�4?݇���ݫ=��i:i��������<�a)>�b=��*=��J>���>�?��4?ZQ?�y
>�-��}��ɉ�
��?�5?���>5�F>�6*>������'�<V�>.K��`󋾁���5h��� �M�=���>��>��9>0À?�Rt?��%?�)>��F�������������9@\>X�>l��>��H��zz-�N(e�M�#��*�N�|�e�>��(�Ȟ=i7e>)��=��=�<e�᳴�?CA>�>�=D�L>Ԉ�>p?`[*?�?NX�>7��>p%�,y��e�J?0�����E���<о���5y>�$C>!{�	P?i�
�2�}�1��ҝ;��r�>�?+��?I�d?�,?��|�{[>T�R>#�>��q<�:��M�#��z�/>t��=a
u�y���g��;��[>H�v>�<̽�Ǿ���*
J�⽽���K�d�Y������a`��ꐾ�z<�|�$
C�t��� ʾw�p����@�M���C;�����Il����?t`�?fO>�ھ�a��%������L�>����vI�����Kꩾ{	����ݾwڝ�K�;~Ij�K�~���6�E�{>
7�=����瑿T<��w�>�f>��?5f��U�D��xR��;!����>�;̾�1������:���0˾���?n� ?8-�Æ���>7��m#??&��5D�>������Y?Ԝ=?
�W?VP��@�觿�"V>�?(0�?H�9?��-���6��T��T���?�ͽ>s�?s���g��U'��7?�LL?;�>�$0��ȓ�`�!�ʗ�>M��?Y�O���F>Z�?�Y�>ڧ7������di�����,&��u>�==�'!�N��:9i��T�=�|�>�n�>!s^�SJܾ Y�>���]�7����������8��=_�>AI#���4>���=*O>��k��wI�����n�.?���?
]?�Q?�پ�ǾOO*���>���>ɒ�>�������O�>(��>���mr������D?�B�?�
�?��.?����y�G���.޸�uwѾ���=�T�=���=x�=�/>".�=G9<���0�p��
�>g�b>s$�>�ܒ>�ʇ>�v >����U��_@������<O8�P��+L��������U`�<L�\�����پ�s�0b&=r.���[��6p6�*/��욾e�>���>��>�8>�M=O�>����)�Ǿ����ꭾ�8,�����q��-m�N�σ$�)�&�$t���r+�LX���>U��z�o? AK=��>���>�.�<OL�>�>V`�>�>}��>��>�
�>e�u>m)�<�R�ӗ�>�P��dH���(V��O�f�6>�&g?��\�B�?�P�������������?"]�>a�q�ȿe���?���=���F�>�k.���H>�U?�h`�YN��3����0��J|�!�L=m*>Va=9�f��¾��G��k�=8n�>[��Q��=���>t\%?�߀?��A?�z>X�?��>|��>��M> �]>���>��>d?ȷ4?��C?��>�`�=Q��cO>�%>�����>��4'� �;=A?�Agu=Nb��C��֐p=�o
��ci=�� =D�Y���m�/�W<G��>t�,?��>�� ?^�����:�O\X��$Ѿ���=��>�ǰ>Hd�>-.2?+�?���>YSo>�|=1X��Wc���> ��>��3�<�v���=l�>���4Z?U�s?���.�l��[6>P6��7�>8i(?�zJ?��>�ڀ>�;�����g0׿ُ"�#�$�q>}��G������>���X����;
�,���	���G��[>�ʍ>.uy>o@`>a)>.:>���>�f>Ҁ)=�=�E��ʰ��u�C�k=�P����S�ѽ����E��⽟�s��R���˽&�ýu72��?�i?u'����f�����J=��I��>��>F!�>��>��=�o���U��sA�vVG�h�>��h?���> 9�X�=��.�q��:�Գ>�8�>V'>5�a��朘��<��>��?�_�>�"��d[�ąo�M�
���>uv�=��_��8�?TU?dt��[tt�����_.�V+9��F�<Ƴ$�Hpݾ����<�����&�g�'Fp�р<��>J��?��}���=S���Ր��ΰ�R4߾�l=#�<\��>��<��D����:B����}��n�T�{^$>Z��>9j�=��>�#?�{?�P?���>���z�*?��$>F�5?��1?�(?P�H?��>Z?I&?ɾ�>�]���ٽ�뙾Xe3�ETp=y�=���>W)�>��K=����W�=5`s>�)���~��|	>��绉O��i��5o�=Ө>.*?�0/?_�	����⧊<���,ѽ䬍=詋>�	޻�s%���>�q>�L?	�0?F.�>>�>����l�l��c�=IQ?V(?���>2��=�:>]R˾S�>�Q���y>KU)��F��t۾8����V�����>PW�>Xw>a�}>S��?�cy?!�>�ڽ��,�䳢���N���b�8�=���<��y�k�*��g��K�!�o�>���[6���L��/=���Ň�=%�t>�%=.T@>�μb$>j�9��+��b>z�?�@?�J�>���>�4�>q�{����Z�I?-���d�f꠾9yоTB���>�<>��8�?���W�}�����I=����>��?���?q<d?�C�����\>Q[V>=
>��0<��>��9�G�����3>f�=#�y�h����;��\>?y>��ɽ��ʾ�3侌�H��ҿ yl��#V�f& �&���p%��P%��d:>��s��?k����J���$��Ȱw��p�<!潲0���W̾�b��ﲚ?��?�It�����+C���"�&�о?�>����c���*��	��r�qp%�m���u¾⊋��݈��_1�yNH>��H�f%��!\G��~p�XP.����>>�{�mN-��g�j'��ݭF=����D�`���vŮ�׫��S�n?�P$?�����w��3�b>B/J���>}]$>ՂP>�ϾyI>6�?p-I?\P?�J4�������K3>�γ?GP�?')?�%W�}d1�>����2ؾ��>ɧ?,�?�%��վ�ѽ��? �F?���=&gp��ä�2�$�9��>��?�jV��>f@?]�>�O�C+�"3=ml��%P3�L�>���o�ʼ������>���>�8�>U�,�Ӵ����>@���&O���H�<���H�<�?J����>h>��>�(�ZɌ�����q&�`dL?�?�?�:S?�(8?�����}��{���~�=Fk�>�u�>���=���$�>�}�>� 羽r�2g�G?G�?���?h2Z?R�m�럿�A|�Z���*���nt�='d�=8܌>S�;]\3>p�G=x=����<� >Q2�>�}�>�L�>$%9>��r>D�%>Z��$���ߪ�P���Сo�?UF��9�P��뾖6��~6K��%��u���������	����.Ͼf ����E��)v�y��A��>"�><[^>JY>V�>�М�ӓ���ʽrB��`����ݾ�ž܎����w�9��p(9�My������ʾ@?*�/=>&п>�Z�=E��=�\u>�'�=�G�=�]>�_>.U�=Z�>k]�>g�^> �>n�=j�[�R;>z-��ј�����q��dP>��C?�=3���+��3{��9��{a�"�>a�
?��^>P m������q���U?����R��'i���>�
5 ?�/�>�@�=L-��T��Gꕽ[Q��Z��<V��=`˽�Nb��{���@�Cu>���>�Dվ�>��{>��3?E�?*W1?�I<�k�>1O�>v��>��E>Je>*��>>�>�7-?�W?��K?���>���=05��]��=�>����mO=C@�=���;Ӎ�<ǹ	����<���
�=�Ͼ�yv�<���=���Β��~�p=�Y?�jI?�?f�?܏��K%���;�8y�pE�=A�'>~ڠ>��?<-?�?�-
?ˉ�> ��=�ȇ�ד'��R�>�Z�>��&�XP��F�=!�:>]n>ч?��?�|��M�;���z>x>�>�.-?�b?�)#?��>�A�>�ca���%�ӿ��"�K=����9[��/�=d���| ׽/�=�
� i���=y�U>�'_>D�0>�>v�>�:�>/��>Ee�= >>F/>�U
>��l���=��N=��(��L�=���<2i����=����9�<�_=\P=`e��u= ??f?���ḏ�!Vb��)��˵����>F�>W��>y��>��='��
kV�]�A�� M�A��>y{g?��>�5�ތ�=�8��I@;F�>~��>BC>+�[�j������c�@<�1�>��?�1�>s���X���l���
�oܢ>����H�X�3ȍ?�P?����ʾ�����S��_��ni��a�=!�Ѿ�ɾ�pH���`��z#���)@��ؼ�>k��>�?�z"�����ξ��������q��z�=+����>�!<>���d����:�]�4�y ؾ�@�=(L�>c�o>�Q�>�?��?��`?�R?��?�<y�Y?Qe�<g?/��>�J�>W�9?�;?�x�>D��>6�m>�̽�圽�噾GL�%�9��7�,�I>�O�>�AQ=b�j=#>�T�=]5��/R"�<�M���L<�,�<5]=���=�X�=�8?�d%?߬Ļ�Z=��	:��o�%��&>��;>(^�=���ǉ<ʉ�>��>f�3?���>7�>�ߖ��k��}��I,�=�a?�?���>�8�=�{.>���1lh��zC=��o>�\��Fv���¾D�����ǽڵ�>��>��>98>Q�S?_�@?�n�>���=���M'��;�b�,�|>d�:.�V>B/A>�0����0���m�����.�(�ઢ���>5�����<'ᑽs��>#(�=a7�=ּ�=��S>��=i��=�t���ޕ;w�?��>�� ?ן�>>�q�������I?u���X��Š�^qоP���>�<>�#�<�?�����}�Z��bE=����>��?���?�4d?�D����\>KV>��>�0<�>�f�������3>'��=�y�/�Т;F.]>�Oy>\)ɽ	�ʾD5��I����3TH��>������৾��	t �EW�hy@�z�ٽV�%�a�=������ �ﾽ���f:־/¾��J?�x?>$e�q�&��:J�8����׾#�=�[������g��ƌ�P#��'R
�	�ž. ��_��R��4!��[>uT�$W���0��lGZ����o�>��Y?%p�6�߾ɝ0����=jJӼ�����m����z��	�E??�;?�#��^3�^C�=��1>��S>$�$>��w>���6Κ=ͮ�>CR?M�	?��=7���ẻ�$O>��?�ݦ?�7?���\�I�[�	�itw�Ff�>���>�W�>�����^��J\����?uH'?菺>��
��D���|��6�>RF?�B�s�=f��>J�>	�=�{�x\ܽ��پ��H<��J>�ʁ=KG����[���ϽCĉ=��>�u�>�78���ɾZ�>e���C�j�@�ւ�/�K���=���>����I>�l_>��,>�&�=���e����C��z@?W#�?�Z?ۨ(?(��exľ��:��]>�ܔ>u��>B��;�	��h<�>���>�F���r����e?���?���?�w\?�
{��	���Ǜ�hپ�𓾸s�=��>�jS>�B���<�L>ُ�=��-=�>yD?��}>f��>b��>A%�>�%=�-��v+�����Y��Pe�>#���?���"� �!����&�XTξ �������灾u�!�P(���ν��9�Pˬ���ڽ+�?%fg>���> �����>g�Ⱦ�v(����Jҽ�������ӾX>��ԾU��j�3��a�Aq�>��qc�>N���nK�=x�?mLԻr�=�W�>����q>��=(h���޹>���>���>�RT>��k>I�B�^F'�\Y�=�X���7���0d���߼H��=
 �?;bj=JtE�����m��M��l
>�\>?��>��.���������	?w��=��Ⱦ
�����=���>�Q?Z�;�����_ٞ���罝�r���=tQ�=�y�=���<P���I���>��?(��2~"=F�>�a?h�?��_?�A=��?=+$�>�>@�<�?U��>%�=?;o?�nv?���>��>��gA�5|5=l��G��=��<��=�<
�=�R���8�>�����g=O��</�=��9L�,�=72?e?K�?'U?��U?��B�8蛾~�2>%�=� 	?�� ?�C?��?�k?}�>S�>���B����>�d>{2/���g��QO=��t>�!>- ?Z�D?����Mn= ��>�k=�Z�>�>=�.?�9+?|�v>H��=�h�I>ҿ�(����������MvW�S������;�B�=k`�5���+,i�+T�>�> �:>�Џ>�n|>���=���>���>y=I�=�ɽC�=����[ �>C��=����<��u!<&�=��C(��#%�����v���U2=m�?֡?uS��+��7)d�r����ά�
�>���>)��>�,�>���=�/�:V���A���I��m�>K6h?L��>�8��̿=��6�/I���d�>��>9�>�d�ul��E��%ģ<�H�>�o?�e�>�l�Z�~�n�-�
��Ԥ>p5=�'�s�?�[?����F侩i�Ν<�|���!�����Dq���v�M���B�ZS�g��1���>���>
�?������=�n⽦�ne�����bo>u�+��0->��>�������6��!��(�4V.>6�v>�C>7��>z�?$Q?Yi_?I� ?�u?�|�w�?��+=�Y?��> O?��0?DF?���>��>{�
>t�V�Q��hb����d�HP��k�=%�>��t>k=�8}=d�t�6l8��ܓ����s��<\���n�<Nq>U��=�D:>�H?�F*?+s���L�=<e��qU�S_ <���=j>"=��.��V3�u �>A��>�$?+e�>��Q='�Ҿ��xK侲��=|�?�a&?���>�PZ<n��=��:�y��'>=M5>^�O��[^�E��B݅����/�>f'�>a/=�d�>9#�?,�??��?=�1=~1�Hv����G��V5>�2'>Q��>t7�`;9��-"��i?���J��%�$�� W��T1z����<|1���zv>I�B�>o?�>>HZ>]�� =Ϣ�=f�Y�N ?J�?��?���>,r�=��ߌ	�k�I?嚡��j���rо�L���>�<>�"�?6����}�s���G=����><��?f��?�?d?�C�5)�=�\>�LV>�>�/<g�>���r�����3>)�=�|y����&I�;^]>�Gy>f�ɽp�ʾ�2�ۇH�i۹�M�a���a���ɾ�Ӿ&,��.����5�=���"�+�n�ݾ��_��|���g����O��|B��򦾥Ꮎ,��?�@�?��>�.7;]� ��Q&�)��f�>��h�Bk����.����'>��B]�]���e��R	G��i�6�j��>ބ�Qƙ��I���)�#>M��>��??���E��gE�U|��Ѝ>~�Ͻ�X���\������`���+E?�?o�������Ѫ=2J	=��D>u}$>]<�<p_��=�e�>t�Y?�[;?�Z�����9����&�+�?�,�?�,?��C�/�0�\���E��\'�>Ԍ?p��>��^����(�8B?�;?0�>�<�٩���I+��׾> A�?�q���>�A.?,
�>�%F<�H�S����jھZ�9�3��>�F>�Ƀ������-��B>��^>8j�>	�)�wm���.�>��ܾa���kp��!�F�>^uj��,�>è���+>�g>aC�>���̊�a^����c���??ץ�?�gv?�c?��C��#K�O��=�<�ȼ>��N>�H>�g�^�>j�>)-��Ѓ�Pоv�8?7��?�@�L/?H�����T{���4�����!V�=�E�=�rN=
I�y8(=�3>�7>��*=��>`d>B61>�Hg>`˥>�=�>��>jx����&�������2$?�5	��B�Չ�h��qu�� ��>.������/������X{�����^&�1��������>
?%�+?9�>��?������d�S��ȾE�hjX����[�G�����\�=��w>4�{ƽp����z�>
���U+�=#��>d��=�nA=��0>d>�D>{�=>I�=���=F��=(�H>�ٴ=��%>�&��c�>u��.h��x���F�����Q�=٩E?��y��Z���9�Sʵ�ʻ����>�}#?@�>_A0�Lˎ�	[���>(���ݨ��	Խ��I����>u��>��=j��;�?������䟽R�?>��>0�>�v�����%_\��!>6i�>g�g>�M>�)?ܙ�?"�M?��=��>�>��C>)�1>w�>�،>V��>�?��?�"?^�>�=9g}�T���s�¼��D�:.����!��Hʽ*̽�ߎ��r��h�o;�m�=��@=��{=j��<k5��n�=�/=��>�?��&?���>�/\�#p=��;��a��O&@<�V�=,��>�jB>t+�>�ϳ>�J�>���>���>W����=�k��>�Y��8KX��ʕ�A[��MH>���>�yg?I]?G�>�-�=(�:�i=Gl�>��C?S�H?�\�>]��s�`����4uͿ�����)�	)����=)c!=��o��W��1d�<?��zY�֨�<F�,>��a>��>,Ê>�l>_�w>Y��>BŌ>&ߍ:�\?=u$M=Xv>�/�=%��=��M�%白���6��<�ib�ǡ���D�C��}S����Wv���???q=HD�<F'�g���j���^�>���>ȓ�>c�>�Cf��6���M����������>��;?ȴ>U�����+>�4�9��>�~?��>��=i�-�KBC�۾�jv�%��>��?�5�>��$���i�?r��f���>K�R=q���:�?A�`?پ(6��Z@ ���^�I�(�ܘ���N��-w�3�վ.o���>�7|�P�־��=;�=��>�d�?�w���->H��Ws�����~Ͼ%�|��.]�6S�>`6\�����}��}�+�U�<l��c��=�n�>��u���D?�>_<�>_�q?!A��5P�>��?VI�>��>�3k?��3>��=My>��>��>�<��������u�<�`].=|��<��R;?F�=xmX=`����Jz=��w<K�8=}#�=)Ԁ<���<�$�:�3�=�Qg=��=��>X�?���>P�N��]u�,�@�|����J1��4=ϴr>��.�Gɻ��>��u>�3�>g$?�G�>;�=©���}�Ձ>~��>�/?��?�]m���N ��1q����<Z�/>wR��+��T\%�L`��V��L>�$h>L�=��7>��q??�;?ӭ??�cw=�M.�������F�3����@+C>�^��7Q�O#�]�5��+D����2������^��0=U�">�X"=Z��=)@f>&i>n^>��p�N�뽤��;(M=lغ>���>�(�><��=��=jbξk��L�]?{��"��6J�s W��?6��r�>�W<>ID7>f|�?�^>{1V����������!?$x�?Y��?[�>�¾
aj�AQ>��>!�_>�G>�`�=�a=b��=��6>[e�=B.������
�<��>��>'Ⱥ����n���=֒ۿOL1��9��v���6��À=�>�}�������[.��I�徜
'�О�$����,�58����Z��N�����?L��?8����#q�QS����4MžM�>�R�Ҕl������Xq��M׾�bо����/�4�7�0��g�>P�Ͼ����r<��u+�1?�>Q�>CZ?S�>
�پ�Q��>�>
+�>�7�>�\���h��⨿��W�?�7?�8ᾗ�D�5��=��L>1�>�$�>�����������"�>n�Z?���?�JD>J����Ŗ�j�<���?�ı?ޛC?�~H�٠#��Vɾ�"�r��>{�?�lJ>��:G��tԾ��H?���?�TT?�i�ޠh������;?�{ ?5#�bW�>b��>i��=c췾����Es��
��'�i�rW>?�=���ýϾ�H��JW���><˳>K�f�v�پ��?c=3��m�G.��D��3">���<��>����=�g�>w>�=�4�[ŋ��m��s۽�*c?[&�?|�?��"?���g|ȾS@���}۽�c�>�>�}>b>�OV?";%?�z!�Sp��-��9?Ԛ�?y�?	�9?�避�ֿ!���v����򳾇��=%ӏ=�w2>���� z=�I�=��<���<��i>NҮ>Ԯ}>�z_>�/*>:�*>}�C>����$�.=��e���AA�o5����Ku�ݾ�na�'-�Ｆ�]��v�P�0 X�4=ٽ��N��E��e���X���>]O�>�=�>l��> �j��q�>���HW�	��#1�(2�S��T��X���Nض�򠙾�Ï�`�Y>�3�#ዾ��>�?@�J>t"�>���x��=�z�>�M�=��>g�I>6��=R=�<#x>]��=Z@8>ř>��=�dD<�Ʃ��(���"����"��,�<5?�w=�������}砾���=��>B?Ź�>v�(���x������?��e�#C��0���r�[�
H>"�?�C>�,?>`Z���Ҿ�+�=��>k��>P��;������j�t�l���	�&8�>�,޾Rv�=k�{>N�?��v?��*?I�=�u�>��>�8�><� >�&>�*>�w>6�??J?i??���>��=>�R��=d;=�/����h���7>��`�gzy<�E���=�q�=txǻ86 <�g!������@<8�<���>k�8?.��>y��>,7�F�>���L�d4�d�>�[��z�>�:�>Xo?zG�>ͽ�>��4>_�k�¾�&�L��>	$@>�:_���w�a����u>+s>��O?��1?�2b�x-b����<���=<'�>n�?)?�k�>9+>+馽�%�L�οg8,��},�����QG�����
3�i�3�@���KA%�QZ�?=�-d>0�>lZt>c(1>, >X�D>j�>�J>>T�T=-��=d��<�?���>��a+=�ٔ�t �<�/���>�cļ����jӖ��Q�Ev�C ϼ]kG���G?�\�>@p=���<놔�� ���*�~
?I@�>fb�>�a?Dߜ>>z��[Xb���r��2����?��?�H�>�����|�>I�+>"���-[>�ۇ����<�=�̬�B�ľ��<H>J��>��>2��������l<�<�`>�>r=�}�'�?��l?E�㾥O���|�8Xo��=�j�:��+��=��80��q7&���=�m�޾p����Q����=C�>؃?�D<��.�����zř�tm�� ��B ��(]y>���>�9
�
@��� ��4�����%��=�W>�%�>�����R?�F�>�{?l4|?��=+#�>qG�>[�?�e�>T ?�M!?�??���>u�=>& ����
>+`E>���;G��T�G�=�Է���n�=:��=!�?�;0�<G:<���=�;C�YIk=@�=�ܭ=m0�=�������< >K�>�ֺ>P��N��@�w�3�_����>|p���T����o��󅤽�7>��)?�i)?G��>�ѽ�r��e¾������>���>t�(?�$?e�f������"���vĺ���>�(1��%����0�S(�e0��q;>��L>�=dY>��u?(~A?(b?�u�<!+*�dc����>͆��_�����= �9;�Xվ�	���C��(~�CE����ȉ��ψ���=rN>;�>��I>@�>�G�>ٙ��R����w�Y��p��=3]�=� �>�e�>��!>�;�u�ʾ@�����?�gT����(�X-*����>'dO��=�\�>-v?�{>�k�ơ����:���>���?��?~�=?����Ł�=�h&>4���w'�>���>�2˽��?�ڦ�=�t>� >���������=7�	?�p?��=;���[����=��׿��7�:���vJ)�c����%������۟$=����)ƾ-f��S6�&�������@t�=i"��V�ݾ�hؾ�ه��V�?�(�?c-��㾍p��S[ƾC���8�V>�>��B˾[$Ӿ��3�K����䎍����S�����O�ھ�w�>��Ծ�Z��i���=��N>�5�>�:)?!�7G�6��T�=o�>�ϟ>!g��?n�UE��J��a?�B?k��ڃ��(1!>p!��?�I�>v��<�׾o�}��ۏ>�k#?MVH?^b"�#1��Z���ӈ=���?1��?w1F?� ��}�:��� �����&�?�q/?T�>"�`������ ��]?BQ?:�?xD;Y�}��A�VV�>g�n?G{a�	;P>���>ɠT>X����$ox�U�Ӿ՛�6'>?�=\݈<�Be��E����׽]=o>��>y�H�ͩپ�.�>��ܾa���kp��!�F�>^uj��,�>è���+>�g>aC�>���̊�a^����c���??ץ�?�gv?�c?��C��#K�O��=�<�ȼ>��N>�H>�g�^�>j�>)-��Ѓ�Pоv�8?7��?�@�L/?H�����T{���4�����!V�=�E�=�rN=
I�y8(=�3>�7>��*=��>`d>B61>�Hg>`˥>�=�>��>jx����&�������2$?�5	��B�Չ�h��qu�� ��>.������/������X{�����^&�1��������>
?%�+?9�>��?������d�S��ȾE�hjX����[�G�����\�=��w>4�{ƽp����z�>
���U+�=#��>d��=�nA=��0>d>�D>{�=>I�=���=F��=(�H>�ٴ=��%>�&��c�>u��.h��x���F�����Q�=٩E?��y��Z���9�Sʵ�ʻ����>�}#?@�>_A0�Lˎ�	[���>(���ݨ��	Խ��I����>u��>��=j��;�?������䟽R�?>��>0�>�v�����%_\��!>6i�>g�g>�M>�)?ܙ�?"�M?��=��>�>��C>)�1>w�>�،>V��>�?��?�"?^�>�=9g}�T���s�¼��D�:.����!��Hʽ*̽�ߎ��r��h�o;�m�=��@=��{=j��<k5��n�=�/=��>�?��&?���>�/\�#p=��;��a��O&@<�V�=,��>�jB>t+�>�ϳ>�J�>���>���>W����=�k��>�Y��8KX��ʕ�A[��MH>���>�yg?I]?G�>�-�=(�:�i=Gl�>��C?S�H?�\�>]��s�`����4uͿ�����)�	)����=)c!=��o��W��1d�<?��zY�֨�<F�,>��a>��>,Ê>�l>_�w>Y��>BŌ>&ߍ:�\?=u$M=Xv>�/�=%��=��M�%白���6��<�ib�ǡ���D�C��}S����Wv���???q=HD�<F'�g���j���^�>���>ȓ�>c�>�Cf��6���M����������>��;?ȴ>U�����+>�4�9��>�~?��>��=i�-�KBC�۾�jv�%��>��?�5�>��$���i�?r��f���>K�R=q���:�?A�`?پ(6��Z@ ���^�I�(�ܘ���N��-w�3�վ.o���>�7|�P�־��=;�=��>�d�?�w���->H��Ws�����~Ͼ%�|��.]�6S�>`6\�����}��}�+�U�<l��c��=�n�>��u���D?�>_<�>_�q?!A��5P�>��?VI�>��>�3k?��3>��=My>��>��>�<��������u�<�`].=|��<��R;?F�=xmX=`����Jz=��w<K�8=}#�=)Ԁ<���<�$�:�3�=�Qg=��=��>X�?���>P�N��]u�,�@�|����J1��4=ϴr>��.�Gɻ��>��u>�3�>g$?�G�>;�=©���}�Ձ>~��>�/?��?�]m���N ��1q����<Z�/>wR��+��T\%�L`��V��L>�$h>L�=��7>��q??�;?ӭ??�cw=�M.�������F�3����@+C>�^��7Q�O#�]�5��+D����2������^��0=U�">�X"=Z��=)@f>&i>n^>��p�N�뽤��;(M=lغ>���>�(�><��=��=jbξk��L�]?{��"��6J�s W��?6��r�>�W<>ID7>f|�?�^>{1V����������!?$x�?Y��?[�>�¾
aj�AQ>��>!�_>�G>�`�=�a=b��=��6>[e�=B.������
�<��>��>'Ⱥ����n���=֒ۿOL1��9��v���6��À=�>�}�������[.��I�徜
'�О�$����,�58����Z��N�����?L��?8����#q�QS����4MžM�>�R�Ҕl������Xq��M׾�bо����/�4�7�0��g�>P�Ͼ����r<��u+�1?�>Q�>CZ?S�>
�پ�Q��>�>
+�>�7�>�\���h��⨿��W�?�7?�8ᾗ�D�5��=��L>1�>�$�>�����������"�>n�Z?���?�JD>J����Ŗ�j�<���?�ı?ޛC?�~H�٠#��Vɾ�"�r��>{�?�lJ>��:G��tԾ��H?���?�TT?�i�ޠh������;?�{ ?5#�bW�>b��>i��=c췾����Es��
��'�i�rW>?�=���ýϾ�H��JW���><˳>K�f�v�پ�`�>���.f��Iot�wy�a[>�"=���>!+ ��H�=���>�K?%=6�fЍ��g���Jx���?}�?�m?4jj?�V��|սqul��Vt>�)\?{=¼����:%�>�;.?d�ξwe�����3!?��?[q�?��N?qj����Կ�E��(��<]��f[�=Q��= >2����=(� >�h=r�+=n�w>t�>�3>q]>���>)�>cS�=�����J#�v]ȿ%ی�1*=����A��F�1Cξ{�p߾D�����/W�Zy��v Ͻ���X�D���~�����>�1?��?Z��>u���ͧ=�������$��s����V�-�H��PϾ�v����8�\�>�S��}O��ƣ�� ?@���a=�;>��%��>��}>7��;CB>�=���=�٢=�B�X�>��>	'o=7��;9��>�pؽ,-\���z��X/���<���]>\�)?^;˼�;�� aN�F����p����>b�8?���>&MJ�r�n�o�7��O�>��+�֨��Ql,��4���&>Bǟ>,Oh>�e>�����_�z�|>�ܻ=��{>�O>��Z�CR�����=��9>t��>�s龽��=}�M>���>��d?�>?M��=��>�J+>zW�=��=X>�hc>.�>��4?�)?�&?�-?�;�=	� ���7=�*�=���nD�hJ½��8��
N�}�=�~�N�(=ac�<n��<+_'=�T=0v$;{���z��<�Y?�7?�G?u0�>m�����|�G��퓾6�9=;Ǆ<雽>�n=P�>
�>qT�>w��>���=�[����ն?_j��w��a��A��>.>S�>�z?jǖ?PP&>إR�ī�<y �=X'�>�m/?ǼZ?��>�Ҕ=I�B=���c�Z�������ݽ��]�2�2�R]�����=��>J��>n<M>��w>f|
>&�ٽZ����>z�b> �Z<��|>y�:>��>������=G�v�^=1t��a��ۦ1�W���&I��C`��Y�I�C�\C;����n�Fq�=3�?�#?q3�>������U�.�V�7��%�=��>�?�i?�$������b8�qt�ІQ��_�>�wo?Ӹ>3��2}�>�'�v=�>C�>*;��݃�����]r־0ʽ��!>�)�>a�u>ƪ{��KZ�����6���Fp>�!�=t���zi�?jr^?Y(ھ�Q/�գ�Wg���(���=,^�1���!L�Q��n�&���ھ��߾�]ɽ�2�<[o?��?��6��<>�,��������|���že:�<~��=���>�g�,����?3�����{C��b���<J�0��>{�y��mG?�`�>�&?�BK?�jB>a1�>�$�>�A�>O�m>ޠ?��\>X7�>xz�=�9>y9>��y>���Z�=�K�n���;9=h��}��BA�=W�>�E��=8�=6g�=�7���aZ=�M�=�üX��<9ͥ=Ž=�Û=��?�i[>`�������l�UQ��܄|=��@��\�=Cۧ�ЩҾ�_/>��F>��?��G?^�?u�z�����+�i�P�ξnE�>��>��A?�.?�k=����|����U���=ߤ>�E��D�!���*��D˾��ؽ��>z�>Zݮ<��q>��g?��???��^>*u
�J䆿��yL�H�S^�=���#-�n1��4�n�P��a_����4nA�wȠ��vG<�㴽�ٟ>W[>��B>~1>z�>�%p�� ����2W�>�QR>�>/�?�z�>�= ���o��g"h?������v?Ͼ��k?�V�=m>[>H>�K1?��=�SS��t����g/�>��?�~�?�Ӿ>����*޼r��=�xi>���>g�^=�Ǿ���<�~=�&>s��>�Ɲ������>���>�I�>�K�������M���a	>7�ſ�N��K�����ػ�1Yo�<G׾��9>�[�_�d=��Ž�'�="R=��y�v�:�A�Ͼ{+���M����,՗?��o?�u}�׽�83�����N_����f>0���J�x�! ��!qC��_��p󙾈`1�����H��s������>_�����t���(�cVh�h��>EDF?ƾ�뼾l�J���<���>�y�>BSԽ<щ�������*��\v?�0?E+�#\�l���Mc��u�>8�;?1q�=�B��EԾ�]X=��P?|�Z?#�^>���\��y�9�9��?�1�?WeH?��꾄��r4�F��wf�>JX?�i�>dp�����=Ծ��?�^�?�_?F���Հ��#���?�� ?N�g�e��>۰�>�z�<`�u��~˾����F���(��b$>��->�t>� ��wԾg�H�� ?���>�L��� �*��>-�辷|����w�� �� =[���w
?�)��db>S�>>ٛ'��&��v������|q?� �?]}?�i�?7lC�V;���^���>><�	?�P>K!��Z��'�y>���>1e.�֘��g���	G"?���?���?p|{?���GGӿ����������=�%�= �>>��޽_ɭ=�K=-˘� Y=�s�>s��>o>&;x>h�T>��<>��.>f����#��ʤ�:ْ��[B�� �ڤ��vg��{	��y�����ȴ���{���[���jГ���G�}���T>��Oҽş�>ii�>�J�>��>�;!a�=���L�:�s�
����<{�{�����]þ[����g#���R����MZ�E�žs��>�c���>)f�>B=��$>՚�>?�L>.@�>�|>6!`=��=��=�Υ>��>�z�=P�3�'�>�����M�9�[�EG��;���x>�0G?�>x��C�e��W��.��:p>��J?�	?gS�����j׾���>�����9Ѿ���E>[ʶ>��1<�@	�c���^����<9��W>"��>���=A轿O��L����=D��>�!ھ���=�mn>�$?��t?<�2?��=��>�
S>z��>#��=?L>��Z>o�>��?O5?$J/?�)�>u=�=�~V���(=�KZ=U�5��6?����,���#��]<�"�94=1�5=T�;��Q=��6=���/�)<��$=�>	?�"?l0?�2�>��R��f �%-0��U��¶�=5K<��>E�>��>q�>���>���>�=>��� �y[�>�FH=�j��K���~\���
>/��>��h?
�`? �^>�������D�[����>�~$?�|H?<9�>�W�=��߽���'ӿ=�$�2�"��/���1�V׏;x�;��Z�&:�e+������<�([>���>Ao>?�C>� >��2>�>�>�H>ⅅ=t�=W��;~��bXX�z�O=����HI<��R��-ϻW�μhm�������H���;�)���2��?�?��=^d$�����H��t��Vj�9�ar>�=�>�?�b���[+���[��df�)e�L��>��k?��y>t��� b�>zd�=Y�>�I�>���=�~�
���;��q�����XE>��>{}>2þxk�s����þ��s>��=W�ίS�?�a?[Ӿ�pm�b[	���V�z� ���@��)J���x�
פ� ��%a'�����AþM���$J�=�{�>/4�?�PR��>lA�O���ddn��Dξ��<��=��>���=l[�RU��nr �j��;^�T�_<��>,���P6?Gs�>c�?�g?���>E<�>�`�>NO�>��>��/?�3�>�:>BH>��>疲>��>׺������Q�z�`Ul�K�üv�ü�W����=!Ŕ=�\��۽<��E=���=�P�=�=C�d=R|;��>��_&="��=�6�=�^?}�>0����?��*�[���>*@=uƽ��j=� ��J���0���U�>�?��&?��>�2�=����|a�P����>���>�?u�?VjM���N���!x��=w�=H�R>9:��p���:"��lϾSof��B�>dy>�@'��6>ms^?��U?|�>?3�=��4�����a5�2Ž���l>��佰���2�(�`]��a�?8j�|��gf	��u��g9<�;�>��>�^>���>�bO>k�>�r��g�e�>�����<���>,h>jM?�*(>ju=�q޾;!Ⱦ]x?���@�����2�a��=`�=/
~=���>?]H?*��bb�	�����\�/?Ս�?y�?�u�>��5�΅���.���^=�W�<��׾�*��L�>>7�>J��>T���+����T>���>�'�>����E�F�C�x>�L�L+2����8+l�Iӥ��|)�ci�1d�=�?���c�=uR�<ُ>�>�n�����w����������X�z�ި?��u?L{���?g��4�9�'��R�ޖ>�=*�ʊýɭ���L��jJ+�������Ҿ;��\���J��7��>4��2�������d�@�M<.o�=��H?>���"��~�?���=�o�>��>�rH�,����������o�?T�<?q9���}� E��(��;�$?@1?��>�Ǒ�����o�>�]T?fi?Z�">�}��$5���k��T��?�}�?r�B?A*���G��-���7(�>�H?���>D\�b
.��ɾQ �>��?,�a?BU�Ň���,+�+k2?��9?=�;�B�?t� ?iV>�@ ����L��; ���H��>�0=�"��.�m<վ	r=B�>���>n򪾬�ʾR?���㦀����yӾ�э>��=�>(r����=�u'>��>#!��|��w��Yq�^1N?�1�?�l[?$�?/竾u�Q��5�d��=�Ñ>8W��c�<+���f �>���>�C$����G/[�?7��?�V�?ݽV?Vat�sۿj|��\W��Ry��L> V�.�>}6�}f�=^��~��� �}jc>)��>C:�>�+w>@2>U��=Q��=�*��B����{����jA����^�jd��^�������-۾^R޾l�k��ߏ�qt�-|(��|�0a�<!Cn����;{D ?i��>��>�>�->Iz���I��9�R���G���
��D��bӾf+��i0�=)<��M�\���o���|���?oR<�"�=��>j���?%>�>:Ӌ<{�]>��T>A_�> �F>�>��>���=�!>��=HV���5�=A6[�������V���%ݿ>�=?)ؾ���n�ྂ�$�~�=gP=�?��>cq�V:I�6莿(j?Sn�<��q�ǣ�=��s�̠>"��>�B��Xp2>�D=����d����<"��=���=:F`�,��0�Z���=�0�>�k�cg>��a>�??Bg?rB?$3�=?�>TP3>l)�>�*!=j3>�`<>�C}>�C?��=?1T!?:L�>���=�5���I>[H�=';���	=�/��D�����Q���Ž�vB<K�(>3��]Zs=�J�S����<*��<˦
?a�F?IW�>��?��U��s�\�[�ZZ�=��>���=��>@V�>y�J?!r�>�?�Jd>���:�w��@��k�>��>1�}������V���>N��>�*V?��?�"�>gy�� �E>�pc>
�?���>��D?#?�w�>.�T=}a�I_ο�?�z����}�r�A�M�2����2��/���/���_��ɼ=-+�>X�>��>d>w >'�V>i[�>�u>�.=?�'�����N =
�<ñ��
{��!<C�<|�*<���l���_���j��(��ô�d����N?��
?�^ ��~b���X������>���g�>�9�>z�>t��>�
D=��k�M�W�9�v�%�֋�>��d?�Z�>��Z�/>�=Q\+����;�k�>ͩ�>�
>��g�5NĽІ���T�=GJ�>R�?D]�>��>�g�d���m�G��s�>��B=�j1��f�?�ia?4�u��yL���'�q�T�����i��c��ʐH����t�=�c�L����~k�K��7�=9��>7A�?�m��k7��p��f����`��v�c�dH{>u	0>^wn>=2��"}c��B���
�%��'����>��=<5�>I<?�?�]X?T��>5�>�dr;X|?��=��3?S�>%�>�f?��>H��>�f�>Wǅ=c��\	U�����	�9>|��=��[>�'$>ͮ�<;?�7��:�9�<Q�i>�ٽQ�<�wa=�_�<�;�=$Df=���<�0�=��?�M?�\=�x��W��n,��=y��>��/?�̈́>x��=c��>�O�>m=!?8%?�i	?��>�|���_����������?1�4?�B�>k�����>��о�\˾ǿ����>�td; ��>������״<��$&>��X>7a!>��Q>��?`�8?3��>��?*�ݾ���|�W��{:�1�!��g0� �Y=V��C��: y��y����y�Q�2i�>�#�� Wμ.�W=�q�>��0=��׼tV�{��>�Z�H|��=Q#��f�?��$>���>�pN>z9=��������V?LN;5��i�.�~ 뾂x�=��:>��=m�Ѿ�?�G��X৿�赿�Ҁ��:�>E�?{w�?<L�?qЪ��|�J�G>���>�z
>�;��i� �!�����1��_H>T=����}���8ެ�&r�>�!�>'��>�����m^�ľ���K�6��S��<���.�ž��2��D�<2P���������\M��ѽ��=��=�m�Dƒ��Y���>���?���?cZ_���%���F��Z�L�8���>����eý��a�,�����������f7��؈�/���1���`%�>����;���5,�`$�ˉ>��?X�'?���Q��C��uy>�J|>��O>Ү�מ���O�����ؠT?(X?��)��;������~�>UE'?i>�э=�Ǿ=�Ž�>r�&?�?`��=���[����o<FE�?Q�?��B?�xi���L�d ����<?��?V��>�͌�b�ʾ9���%?k7?���>�	��'���e��>�Ra?:X@�tH>��>�r�>F�ͽy�����eS��|w+���M>���<l���#~�drU�,=���>��>�{��m���E?����q�x��g)�\�;��.>iX�=�T�>w5�fZ�=~�|>>s�P���@��ƺ��\[?(��?]k?�6?�鱾�}c�d�м�Oy=b�>�\!=s�{=~sB��{�>�$?��)�RN���4�[?��?[�?Ӣe?Կ���uÿ�枿�P���1����=�3�=;�>9���-r=����ϽςU��/>~��>�x�>�t|>�-#>�%>��I>Q}�[����~����P�9��9���L�3,��}���-�8�ʾO����a=G�n�K��Ù;���C��l���@�=�6�>���>�?N�a>�5>p��;ep����⾳}�=��<�����%�hhɾ�Z6�����fZ��K��t�8� �<��?.�<�G��;?�O�GS>2��>�P>hU�>䜻>�(b>�٬>�U�>0�>B�A>ٳ=A�=H��=��">���-����4��M���1�
?�!_?WV���Dν�\B��舾Y�ɾϿ�>�R?\�F>~{���������`?聻=���ad���=��=>�B�>�4 >>H�>�]#�ܩ����=��c=���>:U>3o ��U�H8���I>lp�>�V�.b>�!Y>ߔ?<�?��?�
>���>�T>>�)�>P��= EC>j$.>��>�3?Vc8?�1(?��>gK>��j��Gu>;�=�Cc���{��f���&��|���%=��!��ؕ=��=�-Q��)�=�p	�r�����='OY=�.?_�I?���>��>�?�F�X�<u������>AZ'>F��>`�&?!�?w�>I�>J\>@�d��]���_�h�>�p>�&F��G��h��?��>@�?��K?�*?#�k�\>�N�>�k�>|Y�>�G?�)?���>����uo�.�ݿi����ľ����L��*��%�n�%����w:�Q�������=�??�>x�o>w(Z>v\D>�eg>[�>
}m>Q���\=p5�=!��-퓽�����½SOE=f�>�p��i���)�[x½���F���bx��B�>��?X9?tˍ�����<d�<�Ͼ9�����>���>e��>���>�ꕽ��Y�Q��>������c?Y�c?J��>���Uƽ=��ڽ��=��>�ҙ>�O>:U����m������F>���>�?�	>�}m��i��0j�?����Z>�u==��kJ�?�uG?�N;�z�>�D'R����53���k���ܾ�;��8�B�K7��]�%Y�=��>�F�?�f=���҄@�嬣��&����u��:�v�<��w>�7>k��i����J�����t׾@y8����>u6�=�<�>�jR?g@=?��V?��>2��>��k�C�)?�t�>��?&�?�N?��?c?��>,g�>�V>z������L��ܶ�=c�>��>�P�=˅�>%"�=���=0�k�A��<`�����H���T���6j<,*=s}=ς>�M?z�7?�GC=�͡�HS��y��<��	��(Q>�(?"�>�$��IT>�?o�?/s ?P�?h��>v�8�5�վ��0`r���?�6N?�}�>�����՚>:;�f۾CT���>�Æ�,5=���A���XIn��>���>�7>s>�jl?&�G?�?~��>�;4���s��wn�!�5�bȘ�l��i��MWڼO`$����d���󍿈�C�fyT>3�ǽ�,���=0w�>�?>F��f1�<��>Ք�=�Z�ٺr�\�<��5�>sԒ>���>�'<>ao�=m��J��.�T?eꑾ[��/�����c	>��?>uHt>�{�����>����tӗ��t����0�(�?��?���?�?�L�&�����>\�>��=��<��Ѿ@�;<M��1x>꩷<�����
��|ѽ���>"/>�}�?P�r[��%���淿q[��13�����0��F ���:D�h����l����7:�������z�7T��<s�;[��[��%l��jP�����?%��?�m�����*R�y�7�1�t>�Lྛ��Kٸ�^@�1<ɾ���1���@!����4���F��A6���>�K�u-��#!_��4�卣=�'�>'M?-N��0-�n�#�3p�>���=�<.> Ò�-!���������e�^?h�B?<�"������A4�>�]7?�0�>z��<���
~K����>�*?�5?�͜��.��e���֥r��i�?=/�?��C?$�k�� M�UJ�|���?�~?�P�>?��X�ξA����	?
�9?lѻ>�6��膿���@�?�k?�9��DU>@��>1ו>W8����z�[���S/��db���f>�r�<�����Z�؊�lJ=��><��>�hԽ`ﭾ[]?*���m��NE��v&�}m�>~��=���>5:�.G�A��>�39>]u�����,���V��@�K?J~�?�{�?=#?���ʫ�ϝ��F}����=X�ܽ�M>vU��wF>��?g�I#���\��Q<?Mi @���?�O?ޙ��<OۿX���Y�������b$>J2�=��>�>ٽ~�={j�='+�x����*>ub�>
�>~�>y�=>��D>��5>�҃�I4�����k��B?�E�従,����(3���N�~��	Z׾5�ؾ-:	�:�<���������>�4�I����>��e>�^3>8n�>���K�>MU��޾�p�~���'��`/�f��,���-��Bz>�zl��N��f)ܽ��.��(?����3�t� ?n��n２e�>ݴY=�M>���>�2�>=3
>/ �>�(>a�>�J>�c�=v$>q�>`w�K����h�m��E�>$N�?DžtC�6-M��G �j����]~>��1?e�1>��@��4�����)��>>��=n>�n�.�
\�A�g>.=?	 =/ .���>���%��q\<��4��J>dy���1��d6�:/>f��>��ٹ�=��->�?&�?O�?�"�=d��>:�=�*�>,�=Q�>أ�=��>�-?�xH?�4,?���>A>���[S>���=���EU���� ���<�J�����<T�8��<��>�y��Χ����¼��E�#���q�1=���>ki:?i�?5��>p}a�,�>�� d���U��>�>�!�>��>�3?a�>"v�>��\>��A�wJ����!��%�>岑>ݴf�y����Q�]٢>L`>[Lj?�!?\&1>3������=�> A�>슧>��?�8 ?�'�>�1<i7�mPѿy�۾����Q>��3=�8�< ���>)�N_����G����>=���>u��>?R�>0Y�>�DN>y��>��>=�>=��=�?�������5�Aء=�����0�\u�<wl8��U9=h%%�<#�9Q,��tѽ����Ďb�Y�?<x ?^��}-�G�=�e������=6�>��>��>~.�>'������>�9�w�;���ڽ-�?�_\?��>�劾���=���_���6?u��>B�>;c���=��S�)��=��?�i?¶>�/b���^�A�d�������>a*�=A�����?�!F?����&���<�h<%�'d������\��3������:�XDW�������>��'b(�ξ>���?����,=�(�h4��<,r�v�޾}�8��)�=☦>��=n�`�pǶ��CB����'I�=��'>K'N>�8^��?!�G?Ա~?ս?�m�>�J�� A?�E?X/?GZ/?z�?#1;?c��>J��>�w�>N�=�v#=Hhj������<@��=}��=k�>��8>븆=� ��1�S���f=dּ7~�l">��=��<n@<�[��W>�'?y#?^��<����b�=N�̽���Ȏ�>fwu>���<J���q�=X>�>k#?��"?���>IS�=\'�����h	���q�<�?�G?v=?��2��Y�=Ye��B��$�=`��>$㏻�����%��)�J��Q��P/L>�"�>}f >*�>��?1P?淢>/��W�b���z��c���H퍽���>Ͻ�=	�'�@=�z�V�G+��}������.��H/콁�i�>Ksl>��p=n	o=8L�=}�N�&9>Y�N<%����2>���>���>0/�>CR�>][>�ŽU<���DY?`x��9�H��K����,�:�8=y�>�=����>v���)����ξ�xM����>k�?��?�[z?�K������ᛛ>���>J�=� J> ޾&�@=��J<zN�=!a7>G� ��ӽ�zj=?�>��;>Pb8���+�&����c<���"Z�m��?Ѿ��˾������u�s$�=�D��"���8V��;���`<ƽ|{��d���2ӽ����������9!�?��?x����8�@T����Ǒ�����>����� =�c����C�=���aݾ챾& ��`�� d���F����>Xy��D��fBa���k��H�7�;?/�&? ��F�}��^i�Ӄ�>)��=l�Ƚ��־��/똿6�{�?��B?h��\h��t>̜>q�>�B�>q�M� 8��3ؾ���>��_?�?��Y>�F��#x���^�=�L�?c��?h�A?Ry>��VQ�����of6���?�)?�K�>y���;/Ҿq?�Ɍ? L8?�j�>Ϡ���������?��v?��5���[>)	�>���>�⽵i'��;o��/�(=sG>32�=~�7�'�H���Z���9=���>��>�{˽����R�?�$ʾ�ņ���%��O�A��>.K����>F����=�>>>�>ޜ��x��^Ţ��Yӽf�-?���?|�c?Ĵ
?d��F�˽����`�p�t>������=s�~�Z�>(T�>y�>���|�Q�[����>h��?)\@� X?�4���.ֿ8㟿hy��I�����>�y�@@�=�s�p�=P��<��ѽ>R0�o�^��5�><
�>�V�>b�`>��D>9b.>�U���[�*g��-$���-�n���?�:����?���t���� ����p����������;���M5�2q���L�=K�h���>ܤ>#�>�?ؙ>�ǃ=����:���M�ρ���61̾L�����^m���[=Ef��e���ᗽ�R+�!cN?�f��r�I�>��:��<�>u�>�HL>8<U>sF�>�$�>�%o>���>嵧>~3>��c>`J�=H:>��D>+p��P��ȝ��:��&�>%�G?���g�&=�~���@P����C�=(;�>�n;!�����nڐ�la?׫E<�׾�1=�B�<Y�7>��?�	R>��|>U��-��j�wJ>�2 ?�r<��h�z����UA��H>���>(��vq>��Z>\�?��{?�$?��'>�>]�>��>6[>��>���=�<�>;?#")?}�3? ��>�6>�=���P}>@&=>{㈾�T�<i���H
����N��-��\���!>�}r=&�>/E"�,풾S� =M�ͨ?9R8?�*�>�\?�z��`
q���1>���>5�2=S?z��>v$?v�?@ټ>p	g>"=�Z���6�ǝ�>��J>�.g����Y[v��:�>'pJ>�pM?�+?���>3,����=���>���>���>��4?1
?�
�>�!o=q����Ͽ�p��q2��Ä=f����۽�ɾFJ�?��-`��� �p�F����>ZN�>I��>�li>ۙ>��>|q�>ܱ6>gv���ۆ=���8�0=���=�"�=jU�=r�=b�>�-��kܒ�-�|�^�����j�v�Lt?�?�����l��d�5��=�|���K�>ݵE>�m?���>���'&뾲$^�?cT�Q���u�>�=T?�N�>�s���X�=-]F�����'(?2�>t+�>ws^�BWH�t����=��?k�?w��>�S��3�u�`�q����_�>��=-��
�?faM?�LȾ��H��:��<�y�=�7���������X� D��-�4�&�1�0��
���r5>@��>���?Q���˟ɽǤ=����V)u��&��?�=����k�>2i~=�h��i��j�w���Ӿ��ǽ�i�>8xJ>�W>j.?	bA?WjY?�2?l�,?5�1�#,"?��="�!?�k?�?P6'?O5%?�$ ?j��>J���兽��9�C$��\kན�@;R��=aB$=�d[��<�<E�=�����q��:έ���\�S�=6���~z�<yg�=uz?{�??�i=|Ž.���HV���l>�f�>� �>��H����p�=��?ȋ2?>?���>�,�>����/�ھ���)�6���?b�V?Tp?;�p=u�6>	�n��p=' �>�[��$���z̅�����.�>S>��/>�4�>�[�?�O?y��>C|9>p��e'x��4T�r��>���6�>��=�Y��P��2HK��������_dY�5B�=�/�s��s{;�0�>�>e:���>T��>�,�=�eW�H�<��!��Z�=���>��?ߒ�>��I>jվ�N3���O?$�m���(���m�Ѯ���=�>ڽ�S>�C¾��?�3�4���E����}�#�`=|)�?g�?4h�?��u����"F>�J�>KK>�=����;��J���>�X>a���u��=m�o!>�}�> 1�7Ծb}=���0�h^��%F�#�i�@�������L��� H���������<��=���ʽ�L��%���@;_�x�e7��EU���I㾡%�?|�?�T�=3�����q�&����]��Z��>b7b�ϛ���&�1�rJ���1"���mm�5���F���:�&^�>�
�@�����_�!{2���_>�J?Q[?3.Ⱦ6	���[�-ӌ>6�6>&->BQ��_�������:�
�S?�P:?$��!,�J�,=f��>6qA?>���&_;�֐ݾ�L]��?	X/?]o?�j��秿;T���Ur�� �?"�?�RC?w/�,�G�x��;(��s?�?���>�掾�Ӿ����7?�MC?D��>�U	��x�� �H�?�9a?��C���J>j��>~�>i���j�����D���G��7>/HY���ν $c�f1p��֊=�q�>�*�>��2������5?�Iľ��mI"�Ӧ�F/@>�(>=��>�)꾸W����>��>�����=������r�T?���?Y�o?��!?s1��Ⱦ��׼��>b�K>�Y����=��m��Z�>��?i��"����l��?�N�?s�@ΰo?cT����ֿ�z��.-z�c���=�����=Q�M��r�;-�=��=d&�=��(>��>?��>c&�>�<�>À]>wB�>xă�/!����>�����D�vh�0���,��@��:�����`����*���Z:��i�ܝ��(�*���=��P�Xr�=$�>B�>�x�>��P>5ͭ=���;'
��%�O��۞6�%���v���վ#拽���=�=;����&��(c.��"E?p"�=&�ٽ�r�>�Q�YUh>�`�>�K��ǰ>�T>�6b>X2>�~�>��>Ca!>gs�>v�X;�>N>o�>��h��׃����� ���>�s�?L3�\g`�d�۩澃;���;>}�!?a>�x.��&��G`��!D�>���=HX\���w=�"T��E=�'?K(����=Ƒ�=��	��aT>�Q�=���>��F;n����!��]b� &�>b��>Q�����>?�n>VQ?U؂?N�*?�^=��>/�Q>&5[>ո(>��>mI�>�g�>�?ū)?s�0?��>���=v���#>���>�<O����*#��b<�궽wcc=��t=��='U�;��=ݳV>\�=�[��@�O��j�=�O?p3I?�8�>=:�>6"T<27z���z�?����L?�J>�J�>�H�>�C?.Z�>`��>m�p>x��z��=�(����>2BQ>2m������&����>#�>_�??�%m?��>*�оWy�=�8�>њ�>�Л>,�7?`	?Mb>�C�<!h��n>ʿ�٦�+_,�֐��ݑ����F*��ϑ���>7q<�_޼\A��~'�>��?�\r>��H>{��=3e>|�>�	>�c<���d�����>���;�W>��~���>s���ҧ�W,���"�M�=�<ݽE��"�d����?o?á��@���S�'����B3�>)}�>��>qq�>μ��s�X�/YH�pe�k?�W?��>�ɏ���#>K;6�ܼ�y?Hc�> �?>|L��j�ν�ݾ�9=���>Q�,?�H�>��z��Uh�˘u�]'��օ>�}�=)����?G�c?������R����-8�Y[�!�d���<<�	��FL¾`&V��7M��y�s��}���=ؤ>��?�d8���;�`:9����,~�&U������=+Y�>!�>�K�.��*g=�G,���\T���>�>Pc�>y�?)�Y?:BC?��?PT?�j��J�?�q�>���>�b%?��]?W�^?r�?hG�>~�>�'�=��<���m�����=�%> Y>#m����==F�;ܒ��ߖ��/>�=u�*�������<�{5=�=I�<=*�=Ƭ?d;?w��$�ʾ.���#�>�-=��6>�I?���><���a��=�H�>��
?�'�>�+�>/RD>��վ�'쾁-��J�<v��>�E,?���>�i�>���>p��N�����QD�=b�:�M����m�̾#����H>�ܖ>�QI>�cX>R�?��d?���>���>)z9��Iz�4�S�2x"=?���-ߒ>$�>gս�~�ѝX���������o��J>���{w<;�(<x.>��=�� �����#>�TV>)�]����=�j=��Q>���>�G?�>�:(>O��}	�.U?
k��69@��	�Ji"�� ��\�=Vp�>!ݳ��I�>��&"��,����{e��ʨ>@��?��?��?�T�]���Ӯ�>"�?�w>[�9�,�����=>��"���E��>#X������k���>
|/>M�y��*	��eB��+�����3�\��5D�:����;���ȉ����w=�B���V��*��^����V�?*���=�p6�N���)l~�"G޾૟?�$�?��
�#5%� �L�)��������>k�_�4��ǒ�������o��Y�������#ҾLD>��x$���9�u!�>W��Q����K�yM�a�� �7?+rK?�饾�-ʾܶn�\?�>Խ>ت�=�V������M����.�0x?��F?��վ��P��^/���w>��?E�?>�	�;$���|&���g?��C?KN?�;����Ml����<c�?AH�?��??DaM� A���_�z?��?#��>iT��@�˾؇���n?C�:?�Խ>R��������`��>�[?D�M���_>���>���>g#�F��8Q%��������7>%_�՛�O�g��;���=`̠>�
w>�HZ���EL? z&�������L��=O辶�|=�+�>�n���+�>5 ���yW>]?5��Õ��Y���2Z��`<?�N�?�l�?(X9?F�������R�>�,�g.N>0��>�����������>��>K~L��}�=+�٣
?k��?�H	@��V?�����^ο����ાs����]�=�	>�,>����@�=�#�<&�ݼ���?>Uّ> d{>+z>�y3>_�;>5}+>���<�#�|���pg��B�9�����>�������
�05_����$H��2���˽6c����Q�*�K������5W����0>�{�=Q!�>���>��t>�3>��w�t�[��(�����$�C�ʻ"�)�����8��j��<ђ��n���^⽁s-���D?BB��ű����>����]\>�%?�J<>�}B> Ƙ>�W>��n>+1�<�?>� >r.?>Ф=��>r-=wR������Gu��A*�|�p=^8g?�˽�񾠠S�|���h����=>l��>U6�>�M4�����=@}���?�X�=gɾ	���S�=�j�=���>g�>��Y<b����󑾮������=z�>�:k>����_���K =J��>�����A>6D�>O�>o�?!�Q?���>]��>X��=?��>�>H�>��>E=�>�?�'?�?���>�c�=�X8��&*�U�ּ�5K�p�׽l�x<�
=̘��nE���4���>�.�=ʦ��w=�x�=��S�(:��=R��>��e?'��>��>	&���f��nw��0v��0�>��6>�!�>���>�=?��*?�	?�"6>��@���.���F�!j�>'#_>�5i�%��{x½d�ƽ, 
>o�}?^Uz?�b�=�ž�o=xg=�$�>~b�>ٺ?�$�>Y��>���;bM�jAͿӐ�Ju.��'�_>�j =v�>�pJe���W��w��#*H�\�Ľ;�L>��>�B7>���=�g�[�=��?��%>��½[sý���o=W���K>b[<��!�� ���Z������ِ��B���<����uͽy6��Y?�?�Y�F.��z���CΦ��Ғ>(�=E��>�>7�9��_&��\�V�4�Ƕ� D�>��^?o�>Ҹ����S>!*8�o�=�?q?���=� ����3"����>[�>wW"?&^�>ㄉ��a�Jl�z}*�[�5>��=�ؽѓ�?��2?��ξ���V�M��4S����R��=���Xʓ���߾'A�&�y�B���
��F����r<�r�>6�?�(j�=�Ll��髿Rw��)$��u{��LS��v�>'�5>Д�C��=	`��1'���ھz�t���>��y>,�>�(*?�6A?��	?*O?T�(?���=��>FD<l2?v>�>1|?#C?|?��=|7u>m3C>�RH>y���4����ɽ����R��=�ω>���=�iV<YZT<f�=T�<�ꬽsŗ���k=��Ҽ�'ؼ��X���:ި=��?>�J?��=�����%�Q��w��Lݝ>��>v :>ug�f*D>	��>�?�D?�>$��>�~��^���k���V�n"?�ZY?#{�>�D>�7�>_�����zE�}q�>쐵<9$R�n�?�����޽a�e>G%�>�p�>"p=J�?Q?#*(?�,N�bJ0�� ����l�N�<�����>֋�>���=���Z[�X����\��3|��o��v��˭�<���=��>��<TfM>GP>я�����m�����;v��Ƽ�>�?�N?�O�>u��=�h��J���Cf?�����>���;���;yþ�>�ua�)��b�x?�?��7���3���腿d��>a�?q7�?��?��^����� ?��>�M>?a|�Q��˥��rhZ�>�����[=7=��Ӂ��X�ý� �>!s�>.�����=�����4���jT��A`��L���꾜P�� ��=�p�C���`�A�ӾBJ�"҄���:�1<]�d]�I(��Y�������Ț?��?e�>�z��v>���cx¾�z$>�-G��c�Q޾X���Ѵx����	��ԩ¾�)��5%��w��Φ>5��H��^O����̾k���!n>�=a?���Ī���XU�U��>d�;>U<P(��搿��]VZ�R+_?��;?d� �v2��C<U? > T>~���<5��;>��I>�=C?�(?����F���{�����<
B�?�U�?i�??|�P�o�A�XL��3���?��? �>&E���̾W����h?�9?8U�>�-�Du���k��Q�>9\?�M��Da>�\�>&��>��n���e(������+��:>l���+�aai���?�S;�=H�>%�y>��Z�
#����?�?��bn�$�Y��Q�<8M����y=V]�>�Lw���=w*�=��ʻ�b4�����pt�j�p�V("?�?�w�?��&?G����Y��>��;�?�P=d�?�&�l?��y%�>��>tq����EJ���?I��?�@�F]?�+���Ƽ��蒿�ƒ�X����>�b8��.=>j��W|�Nv��x���J̽Gv�=W{�>��o>u0> a\>�=>t,�=��~��
"��R���Bv��H8��^0����<�u�^������*���I���?��=�'f�17��q�� ���Q��5̾�P�>�B�>�j>Q�@>, �>�Ɖ>�C��T;�u���]�����>� |(����r��J���pd>�Y=�b�L�B��H�u�@?���=�)�;�?�,��5�u>ܿ�>k\}<���>n��>0�>���=�9�=��>���=O�>#d�<I�>�ܽ������:p���c-��>�;t?�|���8�)<�]���Fw ��?�>��	?��>��-��-��� ��s�>��]>e��pꔾ����*�>rP?��A>Br>N�Pm׾�pؽ$��=#r�=�J�>^Z��3�L{���  >s�>�Pо�.$>���>��#?��~?��5?��=�î>?�l>;�>B��=��\>��}>(�>��?��3?&�)?(
�>���=��~��=�C�=���Q"��׽B��Њ�<�C�yDi��:�=ZY�=b!�<Ć�<}�=j���p<�?�<��>�6`?�2?1�>5��p�Y���}��}�J��>1э>+z?yĆ>��?�Y?&�?�N?���=a;վ�(�5��>�tl>��U�C��ʬ*�1B@>�^R=rwo?��m?�
>��n�����CU��g�=�s�>�f0?᡾>Jí>��z=k}���̿���*����K�9#���P��o�e����w������w����Y<���>2�>�n>	5�=k�=����<�U?��q>$g=�P��i����=ƒѼL-6>��=���=��>X϶;�1<>�ѽ罗5�=��2����eS�"#
?�p(?b��|��Wae����8LȾ%"w>��>V?�3>�� �P%�CD��(�\�����>�S?� �>������>1ɽ��->���>�Z�>��=>�A�=vQ���$��>^c�>��?�k�>R�P�$Tg�x�y�+� ��>��#7���6�?��K?G���{+���9��WF����jE<�I�i�/��;g�mN��"d�)z�q����_���=3��>$F�?�߄�`S�>�Rν@���f��yҾ��@=�p;�ܪ>&+�>-=\ ׾��N����2�Ҿ�_C��s�>�[�>S���<?��n?E�6?orr?�?��==��>��8>��?���>VQ�>u�P?+?�lE>2S{>�=��<6\�g�z�&c>���-�B��=��>�l�=�s�<0B<Nj
��R=3y.�C��;[�'=��m=�&=��=h<�; D�=��?w�E?d�=�1n��í��%C������>
X�>r�=$�2�
m�=]K>���>}�9?̢$?6��=�JԾ־ȾӤ���X<�6?�Q?Q��>��=k�>�;S����p3��n>7-�=�.-��e���喾�IZ��w+>�=_l?>10�=g*�?��T?] ?b6��u%8��l����b�o�B�r���>���>�J>����y��C��	�a���E���������=G�0>�>�ϗ�K��<��>�罅<��G=�1�=��<�^��>�3?�>?d>��=�o��N��Y?�W���F�hd���溾O��@7�>| ��H�S�??��׾���������ip�8؄>;޽?sW�?X�?���˔��=�>z��>=�=�>?���U�c���t��;V�kx>ũ��.�+�>$�z>�mu��Ѿ�$�U�g�鷿y>Z��{7�/�ɾ�)þ-X׾�#�����l���v���R��A�b�N�0�IzH��I��=����p�x#ɾβ���~�?��v?��X=.5ƽ��9��@�x�Ҿz�k>�i���U�'i���+��\Ԙ��:��1����Ӿn����/�1�� �>68	�����e���&�G�}�>��^?,�2��f��<��6�>���>X��<��ľs���j���b"��xF?��'?��߾5΋�h9D�M�(?4�>�?i>h?�2�t��ć>1��>1[?�-?Nfٽ�奔l��
H�=��?�J�?Su??K�l�ڡX��=�>�@>���>��?�Й>6��������9��j`?�H?�M�>Ԗ#�ׄ���L�pJ?�ܐ?��̽ߣ�=F��>r>d�=�D���!^�Y�̾���=�AD>����gʾ�ʾ~ܠ����=
t�>�I�>5�=�e"��>��_����M`k��xU>>���=3��>�-m�+E�>3�þ��>�~N����|���3*���2?ξ�?HF�?��-?�d�lL彃��=�`�=��=g��>��I��%��M8?�	U>BbK���> #�T�>���?�@�	i?U�����ݿ,��>����_.�}�w>�=���=�z� �<a0(��P���"�=�j>��w>�Qo>�ņ>��=t�(>�Kh>�Ѓ���x���(���y5�{��)��g��*<�p�}�l�#��:��U���`;�Gls�E���$��7���	˽�c׾r��=;>Pt>|g	?�>]>�(����L����߼=ӿU���c���=����4�����=����A���cܽ~^)�e�G?�Z������w�>��w�	��=��>��4=��.>f4g>{��>�R?�P>�&�>��>��>�5�>�Ӱ>��1>���/���@<f��ݘ�y7���v?9�3=Ɍ7��l/�8���־��>;��>8��>9|2�����oP����	?�{ݼӏ��;�D�R��<H��>�^?e.�=��=�
`�29���mý�h)���>��>"c����5�)��W�{��>�T�p�>��l>�_ ?^�?C�.?T\�=��>%�V>C�>��>Ik�>���>{ҏ>�ޔ>4D	?��>�c	?+]�=���,������y5���=�Mi=��ܽ���<�!�ٽ8%ؽ�3Ž�ث=?��=�)��g�񼝁<z�=ߓ�>��8?-��>���>p.پJ���'C��g��9�B�>��K>�j?���>�k9?�?l7?���>Y	;�����t<����>Ȫ�>�N�Y��ZsI�G ��ž�=,��?Sˁ?Zo�=S���"�j$�=׻�;w��>�G?�Q?�� ?�$�5��8kӿ�$�S�!��悽a����;��<�N�*�=8��-�����V��<�\>��>��p>��D>§>�F3>�U�>�BG>��=�ϥ=��;�(;5F��?M=,�7VH<��P�����
-Ƽ����{���6�I�X?�1����ؼ>U�>�{?����:ሽ1Y���񾃫����>叡>�l?p��>��U�5���u��>7��1��	?�Se?I!�> 釾�(%>�a���[<�>'A?ͪ>d�6�1X���⺾�+>���>�Q?�m�>{=�BE`�k�~��0�/�>o���@B�	��?��??���;գ���9�Q�?�$�[�׻��Y�g~/�����v(��/p���&�
5	�oȟ�2i�=R��>���?R�q�UD�=&ξe���6D���s��>>M��=�-�>�j�>"�)>ʉ۾Ûc���4���ƾM;�ϱw>y��>9?�??��D?$?�/?��>��h<H�u���{�>��=���>�k?~"?Z>�%�=qE��~�A>�_��n�[�=�aT=��0>$-=�O=+W�=OB�<cg���\-=]�I=��=�đ<N�><Q�=τj=u�e<�^㼔Y?�5?&��=�?=i���o�V�6�"��l�>���>�:O=i�����Y��>���>s-?dK�><E>��}��_~�9�پ| �<0?X�I?���>Q�C>�>��&�f�ݾ��<ת�>ܧ�=�7"��'��h���3�9*v=>O>r��>�|��:"C?{�H?Ć�>eƬ�e2�����タP;�𞌽q�?���>u��>�H&�|�o�����j��Us�Z𙾩U����0�[�=��k>R�&>\�6>�>�[c:�p��ܮr���3>�ۼq&�>\H?��N?��>�Ѯ=};��j���?{����6�ھ�����;y��>?3��B�>���?�� �����H���暿3+�=���?��?f}�?ֶ���}���?��>n��>c�	�=l�Ľsk"�>j�=�x�&U{��n��@��[ڼl�i>9É�D
����Df;��>��x�K��z��!������*)�+1���f���T
��a�4�پmI�4����DH��ї=�����뻾�T`���?U��?�/ʾ�)���_���վ�ý���>�̊�U�Iϻ�4����i���;�Z��]�����R�:��
�cB�=�T������Ƙ���|E�Q�����>��X?�z<B�.����!��>��">��w=,�:���fߴ���!�B?!�;?�@���ξd��=�n?��4>T�>;�=�Ƣ�߻�>I�>��??�@?�0���֞�g��jŲ=l�?���?~�C?םP�w?4��W ����x�
?#�?�5�>����oھ�l��8?l�.?�A�>������������S�>�1W?�S�W�v>�o�>Q�>��˓�
�R�����	?�.p'>4(����2��Z���.l��\=��>?4O>&�^�&楾)?M���8���$SH���T�j7�����<gr>۸g����>���Y>Ǚ'�렞�\Wx��*5���(?���?0��?K(?�D��r���C�>xþ�'�=�t�>��4��R
���>F�?Po�����������>Po�?@b@� �?�xz���ҿ���=R���$��>�΁=2�>��=���=��)��R�74��s�
>y/�>�>��8>I�4>c�=��>F��D�!��ؗ�%z���T�O�羮�	�`��V>ܾE뚽��3V���b��2IU�����,��A�	�彵U���Rd>g�>�;�>Z�>�>�>U�=�Ҿ���&脽gI:��)A�y�"��=�m��; ���铻W�=��u+�P�#��� ?f{�=I�=r��>nܽD�=Gٸ>l��V�>�.�> �>��?��>,��>��=2=֕>�O?>`�=�(���U���!��I�)�<h2?�H��#㾴@F��W��4���:>7�?j#T>��I��s��;���C?i%�=�{��tN��1�`>�t�>nx�>-c�=�S��N���_L��E��;D�@>1K#>�ɽ�G���/���$M>�%�>ȻҾ��;>fd�>�?��?u�8?��=1�>@2�>�>�>S�"�m�(>,+�>q��>�T
?E�8?0?�8�>ۖ>X����!>U�Ƚ��R���м�������=��<
*Q=~''����u=��=N�=^�=�S=��ٽu>�_�?�G?r��>:�>�뾌b�z�q��<�[�>L�f��?��?�=?-?�!?S�>F�c��K�֖:�
��>qx�>�<a�N���_)����;��=��r?M^?�3��԰�a��<�;:�>��>ǚ*?��>�ح>�+����	� ڿ�۾�1վ� �=T^�>äd>wLX>,��<׃=+���?s��u��<0��>��p>A9�>ar>6�'�=u<��K�>�Z�=�&H��;��&�`�����)>����F��鹦=9A�={�=����Ш�[�=��vY��л��J%?��#?u� �P�Խ���`�#�g�JFX>��>V^2?n3/=�ښ�ܗ?�P[m���T�w،��
?��u?
��>�ί�խR>O=#��m��?�� ?4�{=-��="tW�H)�Xp>r�>�+?�w�>�<���\��a�����>�lE=���G�?��=?�۾���}P7�d��R6����	罪�S��^����/WT�[�=��:�k��m�=;D�>w�?�jF��u>Es��3.��c���qT�e.X�c[�>D��>���=�N�܀Y���/�sӾߴ(��3�=�>��$>��9?�K=?�{!?�+G?�@D?�]$>+��=���x #?�S�>f�%?mZA?o05?�4�>���>}��<oM >�#�@����k����;ȕ�=.�L>�>��=a��=D}�=��'=9�<�!#��S�=�7���%���<�T�<rӁ=�� ? �_?���=����t��1p��ٽ���>��)?��=q���<>�z>�� ?;�5?r4?�P�>�ŀ��N��+2ھ��F�?6?'�C?We?�:d>��>�#�����ۄ��i>cޜ��Pp��d������Lu�NWM>p^>Wj>��]>�ف?�,S?"L.?�rZ��F�5���g;O�IE`�0D���I>�>�>��>�����*U��p��G	g��Ab��R���$�U��<��>J5�>ƌA=��=�D�>�!>��=�v=�0>�au�Hmq>�H�>R-I?��>b��=���p�޾\RS?�Q��U(#���t���,��"��>qN>3B���G��Z]?�奄�'��uƿ�N��j�>O��?m�?R{�?�#�������y�>�f�>V�>���? �x�x�V~����=I��>���{F��[A�jCD>�V�=ꊅ�/����
q������O^��i����Ѿ�@��	+þ����=y��G��)���ܾ�j��Cr��'��M�D��.��|댾np��K(��P�?��?�<��ק��9U�	g�� �&$0=����m����/q��7���轾&�t�մ���3��#�X�����>��f?��ء�k�۽�b����O>��?�6���P��(4B�=�P>?5��4A۽�K�~����^��GxS��Jd?��3?����(	����=���>�'�>�T�=.퟽��-���=�2>�L?�c.?-���[ޡ�b	��0ox=x�?Ȕ�?Z @?wR�)5G����ս�^?5M?�u�>�����!ž\��*�?��7?�ˮ>���8��|����>�Md?��A�7@U>���>o4�>M��_���0;��=��p�:�fI>1|���O��6a�=eS��Ѹ=�)�>��>�2��=��)?M���8���$SH���T�j7�����<gr>۸g����>���Y>Ǚ'�렞�\Wx��*5���(?���?0��?K(?�D��r���C�>xþ�'�=�t�>��4��R
���>F�?Po�����������>Po�?@b@� �?�xz���ҿ���=R���$��>�΁=2�>��=���=��)��R�74��s�
>y/�>�>��8>I�4>c�=��>F��D�!��ؗ�%z���T�O�羮�	�`��V>ܾE뚽��3V���b��2IU�����,��A�	�彵U���Rd>g�>�;�>Z�>�>�>U�=�Ҿ���&脽gI:��)A�y�"��=�m��; ���铻W�=��u+�P�#��� ?f{�=I�=r��>nܽD�=Gٸ>l��V�>�.�> �>��?��>,��>��=2=֕>�O?>`�=�(���U���!��I�)�<h2?�H��#㾴@F��W��4���:>7�?j#T>��I��s��;���C?i%�=�{��tN��1�`>�t�>nx�>-c�=�S��N���_L��E��;D�@>1K#>�ɽ�G���/���$M>�%�>ȻҾ��;>fd�>�?��?u�8?��=1�>@2�>�>�>S�"�m�(>,+�>q��>�T
?E�8?0?�8�>ۖ>X����!>U�Ƚ��R���м�������=��<
*Q=~''����u=��=N�=^�=�S=��ٽu>�_�?�G?r��>:�>�뾌b�z�q��<�[�>L�f��?��?�=?-?�!?S�>F�c��K�֖:�
��>qx�>�<a�N���_)����;��=��r?M^?�3��԰�a��<�;:�>��>ǚ*?��>�ح>�+����	� ڿ�۾�1վ� �=T^�>äd>wLX>,��<׃=+���?s��u��<0��>��p>A9�>ar>6�'�=u<��K�>�Z�=�&H��;��&�`�����)>����F��鹦=9A�={�=����Ш�[�=��vY��л��J%?��#?u� �P�Խ���`�#�g�JFX>��>V^2?n3/=�ښ�ܗ?�P[m���T�w،��
?��u?
��>�ί�խR>O=#��m��?�� ?4�{=-��="tW�H)�Xp>r�>�+?�w�>�<���\��a�����>�lE=���G�?��=?�۾���}P7�d��R6����	罪�S��^����/WT�[�=��:�k��m�=;D�>w�?�jF��u>Es��3.��c���qT�e.X�c[�>D��>���=�N�܀Y���/�sӾߴ(��3�=�>��$>��9?�K=?�{!?�+G?�@D?�]$>+��=���x #?�S�>f�%?mZA?o05?�4�>���>}��<oM >�#�@����k����;ȕ�=.�L>�>��=a��=D}�=��'=9�<�!#��S�=�7���%���<�T�<rӁ=�� ? �_?���=����t��1p��ٽ���>��)?��=q���<>�z>�� ?;�5?r4?�P�>�ŀ��N��+2ھ��F�?6?'�C?We?�:d>��>�#�����ۄ��i>cޜ��Pp��d������Lu�NWM>p^>Wj>��]>�ف?�,S?"L.?�rZ��F�5���g;O�IE`�0D���I>�>�>��>�����*U��p��G	g��Ab��R���$�U��<��>J5�>ƌA=��=�D�>�!>��=�v=�0>�au�Hmq>�H�>R-I?��>b��=���p�޾\RS?�Q��U(#���t���,��"��>qN>3B���G��Z]?�奄�'��uƿ�N��j�>O��?m�?R{�?�#�������y�>�f�>V�>���? �x�x�V~����=I��>���{F��[A�jCD>�V�=ꊅ�/����
q������O^��i����Ѿ�@��	+þ����=y��G��)���ܾ�j��Cr��'��M�D��.��|댾np��K(��P�?��?�<��ק��9U�	g�� �&$0=����m����/q��7���轾&�t�մ���3��#�X�����>��f?��ء�k�۽�b����O>��?�6���P��(4B�=�P>?5��4A۽�K�~����^��GxS��Jd?��3?����(	����=���>�'�>�T�=.퟽��-���=�2>�L?�c.?-���[ޡ�b	��0ox=x�?Ȕ�?Z @?wR�)5G����ս�^?5M?�u�>�����!ž\��*�?��7?�ˮ>���8��|����>�Md?��A�7@U>���>o4�>M��_���0;��=��p�:�fI>1|���O��6a�=eS��Ѹ=�)�>��>�2��=��)�=?�W#����/���G�Խ�>���>�0�Ʃ>;k�;E�>���k��X���S�����>��?��?^��>������;�ݒ�R)�hU-��x>#�o���T�冂>改>[ �_|����e�><�?J�@�/?�l{�p�׿�&��\S���p���>ɇ�=�_O>*��s3=)s<��=sb�:Gw�=K�>!�W>$Ҁ>��>��H>�(>$ǉ��#�����{���##�B�����	�?ࣾ���|q��M��M���Q������	?���.�R�h�Tc��1C< �p��]>m��>��d>�?>��>V�>i���#�~��������6��龧g�>��$$�=�$��47������@��mk?1;=�D)>$��>�����{�>r�>7��>^��=�	?uɜ>!�3>��	?2�> B�=���=�@>��>��S>����Clv������־9^X�R�u?�Ͼ"�ľ8=}�"椾��ݾ�����>0mF=�A1���������K�>ॊ=y���lY>7^Ҿ"w9>�<�>Ke ��B(>m�ҽ�)�(�W�n�m��S>ݮ�=�N�,���`�R�T�>>U�>�(��U>�׉>B�8?��l?� 9?!y>I��>�x->�n�>}�o>1^�=�#�>{�>?f?��8??�S�>K�9>���(	߼�i@>]쥾��t���0��+�z���Q<�=S5���pü(1��lwm��@>{;>~���I/�eݹ=��>2tB?�ܻ>'|�>C|��J�4r���3�Y��>�e>��;>�>> �s?&v�>� ?B�>�'���P0��j3�yv�>ԝ�>�iC�y��j}��Y��>�s�;h ?}�z?p��:�޾��ټ��=4�?�C?=�?�T�>���<I�輢���y�ÿ���];�n^���}���l�Yi�_�><D���,�K0��u���3>L��>YG�>�V>A�T>Ы�>X��>[n>��}=x�=��#�󽍽�2�
>:�\<�u�/�0�啴=�l"��%�@�1=y����4��Jǽh�l<M`?z�?k���=2ӽ#�H��6!���h����>�&d=R��>mF~>����^O>�Jπ��!��s��C�"?��Y?�E�>Y���k>E��Q�)=��U?:�G?�@�>�S����>�,�x�>��=�z!?w�?��_��F�pp����ˍ>I9�=-�@����?�ac?� �?w��'��9�����=Z�k�6��G�[)F���M��H�_2�o����'A>�j�>�h�?��̾ �>g4����������u)�Ghq>���W�*>I�{>���ؾ�<b��;*��"ؾO ��Xxe>Ǿ=OLC>�?$�C?�:}?)�L?;�`?�^�Q'0?<���YM?�_>��>J\?�?c�?�t?$�r>��������Ō��6�q <���=�h�=��=>��=� ��Q�f��o��;����d;�5Q�E����Ѕ=4�= �x=��?Du?9<3<���'�	����>�er�j�M��??y�?=D���ᾒ��>��?��e?�?�=����)�U��ք<p3
?'`#?,x�>�z>?s�>���ɮȾ��=
�?m� >�Տ�᾽�ؾ=x �>I�?6l >U+�>q�p?,�c?�&[?E���	>A��ͦ��s�v�uc߽��>��>��>�7����L�w�R�{�#�r�N�+��3<�LA����'>>[g*>���p�>Q�Q>v�n�b]S���>�a���H�>��?�?/?i��>�Ų<@N�����W?������莢�v���^�DA->'%>]ϊ��?'w��i�����U�T��CQ>bɳ?��?��|?��%�Qq��}>��>��=i��<Z�������Qx�6��=W�>�b�X�Ҿ�M�=>>�]>�o1���������G�}��DRR�rך�{�-�� ��[�ݾS���k[>�]��6Wu����ٍ��~������k;�������U��&V�����?o2�?c&��4���(�ׇ ��P;���>O�پF��=�߾6��N�p�2\�G!��r#����g�&�{M�>g�.�z���B��<Q���Z���K>�y?&�9��i��|�B�?~�>�Q�X6��������Ŀ�D�I�?��R?q��+-�ݎҽhKr>*�?�>�"Q>/C�o`>��h>��Z?%�s?���=�ß����=�y��p�?���?��B?��T�4=E�Xs������?�X?�y�>����u�þ+$�J?:�;?X�>���4�����*�>O*_?'0H��[>���>6ߓ>���@��٦�'⛾'�C�F.7>��껣��5p��	N���=Cr�>�]�>�K��尾�*?p��nZ��DM����������;�|?RI���>&�T>�?%>���᡿��{�<儾#�]?��?`7|?�1?���IWؾ�BJ���>w]�>є#>*a�=���U	�>	�>�龖����S�=��>��?-N�?��?d͍�tt��R��A'���l��ȿ>��|>�Y1>(�%�"��=2b�����a�"�`�=��>�R>�9>@�E>�f>�|>�]���#�~}���!��ȡ1� ��{�� ��r��h��Cf��ھ�B��2��L���3ɽرz�Ǣ8�q��� 3��v���[;�>�;�>ě2?�;>�T�>M^,>�^!� }ᾶ�����5��v��t�� :��!Ľi� >�ks�B��oQٽI�$�Z?ڛҼ�rG>��>������>X:N>��>?�=l��>ŝ�>]��	f=+ �<�=T=>�Q�=��F>.ҕ=�ב�?fd��4_��馾��">��2?R,]�C��
�9�U���ހ���R>�J?�X�=V%�4���ҹ}�|��>X�����6�<X�R���0>�m�>�B�=�s����*=,'���E��Dn�=8�C>.�/>X9�����#p�m�s>���>Vhܾ���=��l>ڐ+?��v?�\5?�9�=�v�>�\>g�>l��=�O>`?>���>�?�g9?��.?�j�>�ջ=�[��;c=�#=�|J�)B�o����O���!��{L<O��bR=T�={�
<��0=}!%=Q`@��!���@=&��>�3? �>���>��c���;��j^��½�V0>s,w��?c�?�}D?
B3?�8 ?$�=��z���������>ۛE>kZ������=d��>S��=MB?;\?��X��ݓ��A_>�~=�?�n?�r"?&��>)kN���������ѿ] "��V-��_�S��=}�=߭,�ꂽ�M��W�H�Qjɽ��<�8Y>E�j>�\o>��H>��%>]jd>�>���>N·��Q3=�ʻU�A,�Z��=��R��x�<�Ղ��;'<^/����BH��Q
����&���hż�a?i�?g*.������c��T��<������>_��>�k�>Ê�>�T�=Gc�'jT��@�ID��c�>� g?���>U�=�p�=�75�3<�'�>�$�>��>M�f�:W�����"��<&3�>#'?ɝ�>��Z[��ao��U�_�>Tû�k��	�?;>W?�q���F���	�rb�����=��<��R�s`��8�1�t![�P]�Bk�A��^�>��>cԯ?J\Ⱦ�ވ>�d�`Z������}� � U�>u^~>��?��a>,�ɾ��?�Ώ0��⾬m۾3����}�>�3c=�?)y?"w?]Wf?�cV?n\�>�У�DB>?���L�?�?w�A?I.?��?9,�>��m>�*>����U�㟩�����ɞ�=��=��_>`̋>�W���� ��ۘ<|��=9�:=(�+��{��������=�1�=�U�>`�N>+#
?�<?#7���*��͗=��A=D�oי>g�>]���d᛾�)=��>'?�b>?�L�>w�<���kʾS�뾞P&>y��>�?�Y�>�#>�q>����f)��	>���=�c���V�>���Rپd�	��F�>��>�,�=�2�= �[?�'S?x1c?�����&�S郿�OV�LE�=e>,H�>"֊>�q�=�ž��Y�mU��dz��'��ox=�ݽuln<F=��>��=�3� �;>36}>@�U���?��T�<�k���!?�b�>��>(�>�m�<
�j�f���9Qr?���O[2�L\	��~�G�����>���>�<���?C>����cU����,�?���?р�?���?�X�._���6�>p��>ъ�=h�a=^S���h>@����]>i�X��_��1�����?�Y[>������־2>�\�������@�6�W�ξ��"��6��/xl����K�<�F��Uф�K�ؾ��4��|s��=���p�a��V���eZ�����D��?옂?B+j�P|>�"U��jW���c�GFd=��g�\��ܦ���;����վHK��1�0�����t!��k*����v$�>�Vk��䔿��b���b�	�8�c�>k�-?3�ž��q�dG�D��=?\�=��ؽ���]p�������\<���?�o@?���s��f����ck>�?�>��x>k%��N�=�:�>c�?��8?�t^�^8��&}���D>�w�?Zn�?0�??�O�
�A������3?o�?
�>�����̾I��m?H�9?y�>���]���9�*��>>�[?�GN�@xb>2��>2�>��ｔ���+�%��#��y���:>���
�qPh��r>�k��=P��>p�x>��\��鮾�5?hE�IJu��7����ȵ������>t���C�>��>�9�>J�1����W��;���-{?�s�?�g?~J?ĐI�����u�@��>��>�@�>��ͼ:��*)H>B+f>�;Ծ����0�f��>��?i�@�?�ꄿvǿpԕ�^^��n��Y�<!H<��>f����p�=efr=^ͽ�;�=:2>�>V�o>�m>�W>s0�>�\�=�'���!��������Y��U�&���֎��=�@[�������l���	�~�ͽ_{���
`�r�����#���L� ��=7ҷ>�q>wf
?&��=�>�>:��<���p��z�5�K�tl��Rח�~; a����Dľ�{۾�ᮽ L"�Ӊ@?����m�>~��>�6<;0%>:�>ZF�;�:k>���>�ʑ>�Q>�o{>:4=��Y>Ϝ]>'�>�^>Ty�=�	����l�W`���}��@<��S?^�k�"���D��]�����j�>�?�4+>�R"�����wi��3��>��=�G���"=����=w��>���=�m	>�uT������U�X�J=�>́">��)��_���eD�{pq>v��>U�{_>��>dl1?C�i?:$B?��>��+>bߟ=9Λ>��L=ֶA>?�D><O�>��?�$F?Ɲ?�'�>���=��Z���>�g�=�n^�%D��t���$���f���(=v@�<��=�R�=y������<I�=�?��,T����=�?�aK?� ?g�=����"��i�{!��L��=N�>�	�>AɃ>��h?�?r~�>�=�@X��bվS���s�>~
 >)%o�\̎�2��F^�>.��>��-?!D?��<�_���ڽ�0�=�8&?��?ϵ�>G��>MI>��-�{���$v��eh���6�	��ڡ!����>rL�>�;�� >O�� �;>b#<�u�=�<>�+S>�m�	T>;Gv>d�>z�>����)���=nCz>��R��L=��==�o�/,�<��=�
�����-ռ��ȼ�	<�!�����O?��!?�71>�x���Y��%\!�#v���@�=��*?�>?Ԓ>?�����,��-�_�K�#����՘>#�x?D�.?������=�����ɽm��>3��>v�=�F��}����ڹ<�>>D6�>��$?�d:>� ��RW��^�����p�>�� >�Ὦ��?R�`?Tgᾆ����)">�M��*2���׏�����M���n��
N���侊Ӿq����ȴ>p��>k�?#�S�y�m>2�����++���i�kY�>�7/>���=���=�*ݾ㤾��%��̙�bd��R >.�?8��=*�?�5?�s@?9f�?$>?�++?m(��k?�"����!?��?�U)?Ԝ\?��>��v>\��>)�_�1慾/�.�tM��=�V>�@p>��=������>��!>1����ʽ�2>r�=�Cƽm�=�PԼۼAOD=�-�=K^�=<�?�yO?	��������*�>.�=ki/���>��/>o�ܽ'�'���>@�=?�"F?�<�>WΖ��&���!����ˠ�=;�>�U?ee�>��.��>%������U��'P�>�>�>�㾖˾	�ؾ�$�<V�>��6>�>
f�>1=v?�@?^�l?�X2>��Lh����u-�> I��p�-?+FZ>�O>�x+�ج<�Bb�")v����	O:>b�鼿��=J��=V�$=_�{=N�]> ,�<3k�=W%q�4����=��=ƚ!?e�]>1��>(6/>m@=��������i?c��S�M�F��)x�Њ1��6�>��>�l�����>>1�r���u���&Ҿ�wV?��?�)�?��M?�;�#��\Z�>��>��㻳W˼8����>mG�=I�>�	��W����s�U��=>�>CF`>wHA�t`��p"�{7Z�8}���@�}����S�����`�}����<?���<$����� n�<��|�	���7���V���b�����Y��Թ�?t5�?��H���/���T�9�)���鲇>w�˾A�U�q�
�J�t�W�}�ھ����Z׾�)�C@7�@n%��Q�>k<Ž=�����P�&0R��KX�E>f4?�b��Z��YO���\>�m�=�����Ծ�	��M2�������*V?v�9?����cξ����c$>�M�>u1�>\�@<�rY�a�=���>�&?,L
?[Yu�n����U���S&=���?Z��?�X??'b.�=��� 	�&M?g�?���>ŕ��5����� ?�zA?J�>�|�V���=���>h�N?��N��]j>	�>���>L��𴙾(=-<Q%����<M9>�x�X��S񁾭�.�L�=���>;k|>h=M�e\���?�U �Z'X���:�꾏��dt���?��6�U��>�a���6>��'������w��Je3��!??-�?�a?t�$?�i�rb��?���N�>��>?�d>�#������ԛ<S8�>�r���i���k�>���?!�@gFy?�e���ῨE���å�&���
=��C<��V>������=��>O� �5/��>��>&U>w�@>4�Z>&S>�-">�!��n%�6��FЍ��SN�̸�t���W��?��6b��9	��C��+�˾����c�;R1I��cN�����������(P*>�ϵ>"Ţ>mb�>D�=�>����|7����x��:�'4�A�.�)�� ���9��-b=6�Ͻ�
�������.��N?(wr��>��)?~^_��C=�>�>C�>?�q>�e�>B��>b��=p�>�[�=��=��=׬}>���>u�=���D����{`�xc�m�=��M?%�$�����r�X���-�����ky>�??$p>�lC��\���Uq�`y? "=�K���^=�y��D:�1"?<@�=��?�"w2>�z��
��G�")&>H%�>�YL�o��;�,� ��=�M�>xر��@)>7��>I�@?�8~?r�<?=f�=�	�>*�=��>3�2>,�P>��>Լ>��?\�#?=�?�]�>�B>4�"�+����?�p������"���J=�,�Y�<���s��;�m�=r4�:=�5=�=]q|=F��<�?�p+?#��>k�=��伸���@R���a���>�u> ��>Ja�>g6?���>ˋ?>.���U�����"�����>�,>�6����L(�(̛>��>�p?!"?
6�e�+�>�>���<�6?\�c?<X'?�L�>6>=��h��4����e)��.#������=���=z��=[^?=���dO��3��=B�?;Y��=Y>�#�>qA.>|6>$^�=5�>�N(>�<-�2�<���<�62�v(��?��(*<e����6�TI�=�e5=c#��������`<e{��l�v�#z���L?R�9?e�2>��q�OK���;8� �ɺ��7$6?O	'?fn�=���p<�� 4�5Xp�닝��>��?v:?F�)�� >��½�g<���=�C�>m�ϻ�&�>�o��!T��ϖ�>m?ImJ?BN�>�c��`>s�tt���DB��!�>�4�=�	��,�?�iV?-C��I݉��#�D�J�K1ľ�><n� �ھ��پ'f(��U� �Ͼ`R��?�\�|��>1��>�|�? �-��01>�>��t!�����q�5� T>*-�=a�;�t��(��7ː�QI�p#k�tď�B${>� �>9��=�Q�>�&0?ғs?�Mw?T�W?�?X?_璾�~�>s�Ҿ�rK?}:?X&�>��]?¬??��>�]�=P�R��J�8�� ���1���2������f>�)�>:�I>�ɠ=p��=�~9=��=M3N�VkH���t�/�'��L���9�=��!>���>��?�\7?>�
><�4���H���ѽ7I����$X>:���7(�%2]=��&?��9?��I?ȓ>����,�E��3v�aG��,��=%-�>�5X?xeX>FM��6M�>1! �.d�,V���,>sy=]�X��^�@b8��P=^>*&Q>�!�=;x>e�q?�^(?'S'?-�>���5��Z�.��h��&=�o�>\��fk�>�s%����̬���Rl�,U-���>�3)����y=Z8:>B�L>{�@=�"<�t->S�����7.=ӱ���?p} >�e�>%
C>D=�=`a��+OW�YP?1ƃ�Xv�6���3���S�Ǿ�:K>D����پ��?2��1�����lF�/u>�r�?"��?UI�?\g齲㪾�? �>��<$jQ�����Ҩ�<�8��8>/�C���D�z���½���>5��>��/��Wľ(��������K��$���k���鵾\���瞧��#�<�0N���|��$վ�윽�@��
�Vp���½5ꮾ9b���k���ӡ?���?g�h�]Z
��+\����Ԑe�N�Q>nZ�:T��c�����Ͽ��� ��w呾�V����<�ӪS�5�#��>�D��
��CjB��]���ؾ�=�>yxA?$����`*=[Fb�Cr`>ǒ2=1�D���<��+$���-<�d,M?�(?� ��Y���ļ6n>,k�>�k<��>�b���6�>�&�>�F�>�L?����N������=�'�?`��?�p@?]J�>�?�g�	�H3��?*�	?��>;Z��Z˾"��.c
?a�:?��>(;��������Y|�>=�W?��N���b>^��>�F�>,��M&��|�����/���;5>)�N�ݮ�I�g��B<�lv�=)��>Z�v>p*\��0��#?����vK��RK��g�U��#�=�?�`,�в�>dA�<K��> �@��֘�]��� �:m?޷�?i�?f�0?�%"�]�¾��.7�>���>���>���P
��Na>�M?S��Ȣ������?�`�?�@�Lx?�ҏ��wԿC���o�;t�ž��=:S=r�>���jn>2���>=f�սK/�=C��>�ݍ>��r>��>?7L>�V->&у�M&����
����Z+��i2�9�;�R�r����$i���c�����־'� �w�ɽdȾ���\�<��q����SI��V8=���>ҋ>f��>)s�>�tb>7��;�-L��!��j����Q�G:�9z�\����S���˽HU����}��e1�P0G?���OiͽIB?<�����>���>�d>��	=�C�>���>A�>�r�>�<YB=�	6��t�=|��>�/�=�ԁ��Α�%�W���>,2h�i8z?JTj�J<��D������t�ƹ>�L?��F>��3�cҗ�8�v�Li�>�0��;�i=Y���A=�6?
�">rt<><�n;��+Ǚ�n��	�3>V?�=~������2L�hi�=޵�>C�־.��=bvw>��(?�*w?�A6?UU�=���>�Ja>�֏>�=�=%rL>��P>ˈ>��?�9?�1?���>:�=��`��,=�;=�>��CY�쳽_��X�&�ʽ�<
0/���H=�'q=�<�\=*�C=�ɼ�p�;��=*|?�84?�(?�Q�=E����r׾�셿�Wo;	�>���>jY�>�/�>#�7?\M?U�>0v��"C��G���<'����>�;>��2����DF�T�?��>A�s?�? �=}�ﾝ��(��>װF?�N? �'?t�J>�	==D0A�(y���ǿh�0���
�!�!�]�VNv������3>l��!RĽ!"m;iν�u>�En>t�[>�!�=�gv>)4>>L�>ɘJ>���;��<\G��IƵ=���=�7�=0}��x/{�ۆ��7�<8=
n�LQV�(�D=h"<�b�9����?.*?(1>�(m�P�:�'U���4�E��:#?�R-?��>�o��8�N�;�E�i����%پ���>��?��B?U�����=[��)����>k}>Ŋ��uh=>������՘>�)?�{,?��m>��F�ͤO�s>w�N�����J>��>�ͽ���?ciH?�/��������|8�[�B˓<4��ǱȾ�����J�uC���Ѿ"&۾=���I��>���>OD�?���)�C>�Y���y���-��{k0�Fz!?*��=��M><=�q��V<��ʣ(� 5��o�q�^�>��?Au��#?d&S?��b?1�q?V�;?M�i?�g�O�?���:�?��?�1?��I?��>�a�=&Y~>��}=�M�����掾]�==���}� >�K>��>�ø=�e��������=����C;����fQD�o���Ꮳ=��5>��>�\?�=?�Q�B��sΏ�%���`���s> /�>�#p>	:��N$�,�?3W?�G5?�%�>'N��!�
�V���uI6>a�>!�}?)�?:�G�` �>�I��4������J,�>��*>4Q��߾,Aݾ�8����>^y�=a�>�9�>�Ku?`�?�nX?��=�PT�UI��B-��(�<�3��ߢ>��>Y�=['�G�W��	������!���O=V����9�\>��;>���=p0>[>l�G�{��O���5<��,>?Q��>N�?#�9>�^�=�"���Y�
 i?z�	�fD3��(۾�ｾ�-f��+�>=�>��?�-��>�8��⇿����+ ��{2?�&�?F��?k�H?��I����0?�З>aEd>h陻��s�s�n���νl�)>�K;����bO���<v��>��2>��;�����3���O��`���0C�Y�Ѿe�|yU�}�+�]۞����=qp��!N��	�T佦��`�`��Pb�?+Q��R��;�ȉ�N��?��v?���SW.����o���Y7�T��>��澤�;��h��j��=��߽���_n���ľQT��YF�W������>�#���۩���S��|v���սD��>�b?�˽�#���CFN�1�>���=�ᑽ���Re���*����;��:\?ר4?f2��ﻢ�g�ýzH�=&>�8�>��=��R�Sj6>_� >��?6��>����9��M���h��<ц�?�.�?% @?��N��|A�����v0?7?t�>�G���eʾ�C����
?s:? [�>�x�[��Bv��D�>?[?B�M�^b>��>Q�>S9ｆ����"��f��еx��:>�<������j���@����=t�>`�y>lzZ��v��ĸ�>v�龘NO��G� "��� �#á<��?���~�>�i>�6>�)����҅��%��&L?s�?�ZR?d�8?b��5��iP��R�=�*�>�ݭ>���=l|
���>��>@5�(r�^J��s?\x�?�x�?�Z?��m�������R#ƾ7���=_��=�k{>(�Ž���=%Cu��H���G�����=���>$�W>�m0>V�>�:>'�>� ��IT'��
�������b9��I�7��Wh��#�BɈ����:����¾��
�ߤ=��m=eDK��~U��m%����g�1��u?<*�>o��:P��>9�<>؎�;п����<g�:�[� �8����ھ垎�&W��� 뾐N���>ʾH�S�F��}�*?"��T=��?M�>�9<�=V+]>mps>rxs>?�>�L�>�%�>K#O>�e�>gJm=ρ�>ެI=�I?�-=ᛄ��|k�D>>�!.�E�> �T?>�|��݃�2%�\I�����[<&���X>�g9<a��*앿�p���>�D_��@#>=�]��5����$>��X>6��J>�)5>�@��No7��,�=��>��%>Z&<#����������K�> ߂�?<>>~��H�%?�gy?�-�>P��=�6�>;J>s;h>? />�и>��!>[R>��?��?i��>��?V�=��i��<���7#��k6��qڽ�K���q
��!=-
��"��<�*>�V�<�
�=w�R>"	�<���<�E�=��>a�D?�>�j�>\x��[Q�˿X�55�	�߽�[�<�	?k�>��>)�?">�>?�`>X�$>%n[�'���?�>EǓ>$s]�l�r��k>���=���=$�m?Gz>?
���<�3��|��*�Z>���>�?~r?���>!
>h�L~ֿ�� ���.��6�X3��Y�=к;�u�d��[#=��9��^��t�=�%�>��>��k>�rY>�1> :L>֔�>�Z>wc=��!>�L�;�xC�:��M��;ٌg��yf=&�b�|���P�o��m���
��2�!�޽�w�<�,<}#�>��E?�S=yR��c����#]�'�=��?��>_p�>��=?��BhA��I��>����3?P�?"�%?M)�u+���=\#D>�+�>$��>.��>Jg�u���= {�{D�yK?H6?k>�Y%� ;|���U��c��s>-}��J�k���?�_?���.���<$�l�|���2���L>�{��}`<p�z=x�Ҿ^0�p��/� �پe���rR�>�y�?e˫���b>�b��ɣ�j4^��ܪ��
O�v����?#V>���7�J8�O����=��Q�8��>Z�K��A�>��)?Z�>��|?�x*?H7�>��-�\�?�rU�W��>b?�y?��>B�>"���(z>�<A�>�R��8Q��V}��ͽ���<}+>�7�=b�g<�C��3���k	>�ؽ}���?�=���Q�=y�۵�<?>z�?j�?^#�!�꽓�H�Sؠ��/A���=�;k>��8��?��<��EJ>���>=u.?9�?���<��־IƾT����@�=*G?sJ-?�H�>?�<^Z�=>���Mm�o��=Ģ>?i�������1ƾ��|������v>bŝ>�E>kEQ>vu{?�B?c�"?i3����$�q�l��v0����<U肻C��>c�>)�=��վ>4 ���Q�%�(�P���M���»��>D�
>!�b>��=��>�˭=qϽ�����ӻHw�)�>W@�>��>lP*>��P<�����,�>?��\�bB�����5d��y�ǽ1�M=�GM>�"ս�?�uQ��{������3�4��>�!�?���?�mr?y�����g�Y>(�I>/Z>o��<��=�T�@�ƍ�綂>���=cO���T��G�?� >��}>��߽	����x��O��<�����O�L����>�y	�������߽$(�����8!>eר��x���|��Qb�z3(�y��������2�ې���?C��?���q�>��|�!�Z�+�����=�x����v���ϡ�h�پ1\�s�o�X`�t������*_�TP�>Fd��Θ�s�'��"6�M"k��S�>9
?��׾�b��_��,�O>���=s2>\���u�m���}��?=GB?YW������Ͻ'�c>�^ ?�>C�>��ӽɾ�>O:?�&?ӫ!>�㙿7M{��>,�ܮ�?]\�?�Z?�À�1�x�s?����:��(�>��?VfE?K	���O�I`S>��>�͗>t��>+}X���Z�P"�:�>��>/p��mJ>���>���q�-���ec#�ZC)�HD=�d>�2 =���t���f��Q>=��>Wľ=������ɽ��>ᾌ�O��B��f���I�7p�<??D8��i`>��t>�Z>��+�mύ��d�������aG?d��?O?�9?rf��]���KU�`=��>L{�>\��=����>�6�>;ھ�Cl�X���`?\�?��?��]?��q�&��8a��_jѾW�ؾ^C>�eI>��n>����X�=׷j���
�{(=.2Z>n�>�e>CE�<ļ�=޴\>�wc>)͂���&��A�������B�����S'��|����<�GϾׯ��[����<�M�yR �Zx\�S5�=Y�8��ul<�W?�$?�{���>�Xt����f;[���V=������L�<t���j��̏��*AӾ����ž��(��$�_c.?�@
�k����1�>M2
=���=���>�X.>C�1>4�C>��O=��ໆf�>���>���>��`>������^>���=h��Cd^��$=��z�����=p�8?{����_r����Rݾ��fž5p;>��?ҪB>)d�⟂���v�y�>s�6����	�`�9���6ݓ>Z�>6g�=�Ϭ<d���4���s���=a�>Ѵ;>1��0�c�솢��� �%�> �ҼP7�>H�W�*X?(m?H�C?J��=d��>S� >��νbU=���>m��=*n�=;6�>̴T?�d?mO?v4�=6n�R���Q5�X�X�{^�<Y�0<m��<�S ={�R<u潷��<ܥ=0��A��=@�J>���S"�k�?���>�U9?�= >��?�1"��T�"&J���ڽ�n��$��6�3?��%?;��=��>�=?�cu=eY���P���{
�nD�>��o>�MR��S�W�Ƚ)L{>Ә%>9p-?��4?�oE�A�D�!�|��O�>���>��>�D%?��?�y>#���޿��$�DE������<=�[�=:�?�OIϼry����Ͻq� =�T >�2>�>��=3 �=k�=R��=YQ�>��E>i�R=�zv=h�2<GA��	+��C6I=&�����=�۩���]�Mg�O̽F
�?n缦���}����-0���?X�0?/��<��|����U���:���B�>�?h��>��>�4�<���o�A�df��6�<C&?�0�?D+?�G��6<!#>�o=:P�>o�>��>��#�> >��$��p�c����>�>D?�R�>�0(�XgR���a��R�.]>���=��9�z�?��c?R��܌�c�G�O��T���M>��O� $���<��[��=�=�q���]����M�½A�>��?뇉����>���<~����ā��屾y}��9�w�Р	?~?c���"�<�޾c��\�Ҿ�2ؽ�:%>���=>�>��8?l��>j��?�(,?9<?FB��]\�>�޷�r��=���>��1?���>�ӻ>ϴ>w-�>���=O{@>BM�M�������t2.<�t>}�B>�>�=������.�=U�=�fo��� �#2�=��1�'>��>�!x>��?H�?F�k��� ��Sֽ��?<G��=6�V>���s)}�-M}���0>��>�W$?}��>e9=�žZξ�G��f=4 ?h�#?�1�>��=��>O��u<���=��=�!����c�������������>V�T>3��=��i>��|?��A?>g$?�����-���w�n�+�#���10Y�1��>�>�u�=�Zվ�e5��>q�Ob�a�3�a�D�ͩ=���=�>*QD>\n�=��	>�=ܪ��#��Z~�<�-л�C�>*��>[	?�uP>�=�=wQ����M�)?Op���,���7���|��p=��t=��=��f>�;3?�$�&a�>R���OP���?]��?;�?�(?��}�;ٽ�3>#�p>z�1>��=�L4��F�=�DM�2Ak>�>�ٜ�G��I��=D�=f���D3=냾��}:>�Ҹ��@���j��������<���P��]� )��ݺ�=Wf� 뜾ܚ��M���QK\�#�����}̾�0L��6�?���?H�;�;{>M�@�Kwf����=��˾d��<��L��r>�9;� ����HC��zξ��۱վ�\
��$�>��1����h���*��>��mhE>o$?���Cw����vr>�>��m>��Ԙ���V���?����"?d�3?�쾎1Ͼ�<X����>D�%?("> ��>J����؈���>��?��S?n��=o-���p���u��?�??��?#4C?��e�ڇk�Kz�J��ư�>fKA>�[?����t����<���>ZT?p�?T^,�mg��Z�,��l�>��>�?��EU�=7?r<�>�t��p:�C)��j������^��>P���N־P(���Ŵ��=y$�>k�M����o��A�>/�����O��u����������;���>8�;�>-W>�	�=�I<������v�b���J?S�?@�'?L?(�������?<�,���4>�Ϣ>Bi�=<o�Ğ�>%�>̂;�m������?ya�?[c�?~�P?�q�jԿ�,��X�޾,p羉th=�f�<��B=,
��皿<��<NF�<t�<��=E�>�3�>���>�>���>��A>ۡ����+����������G��
�����SVѾ�� ��|m� ��iְ���ﾊ	D��g��������l�b���rr�*���c�<{L)?�?w�Y��>_���z����ܾJ��������uj;%'8�-�0���=����������MI,�ء]?�<��?>�f?��� �,=�_>��)>�;=�K�>��>�UM>��>�'>��=Ʈ�>��B>���>�>d����N��R��r��8����I<?�J��)�{���D�P�8�z�𾃏%='�>��1>��<��������F��>a�i�<�=�t�~#����>���>8����=Rk�=�ľ�bp�g�!=Х=)�8��=$>KT�=�I���&�>������=e!l=ϡ?�R?�G?�TF<�t�>�B/>�>I�Ž��>���>4{k>�«=�?�3?_?�;�=��#��zE<�a"=��8{6�a⼈�<(�r��խ=3�	��G�=�܏=�����@=:�h>I���Ad=cN�=lL?�.^?�\�>,w�>�9�;���������ȑ��FT��L�>�g?��>A��>�`	?.?�߃���@��Q?��h>�K ?�Y{��u��iPk>�X�=�T��~A?���?#L�G܎�t��=#�����<�?�J?+V?̴�>��>"bѿ�©��S�c�P��3��=>t�&>޺���6��^Q���Z����.�D��TR><a�>5s�>���=���c�>���>6Ak>
��="��=+�=��<�!�<�O->�Vf<��+�z\Q��ޞ<�q=�N��X���c	�=� �}��X��l�$?�j?�'Ǽ��=�i�=�#�V���ږ?�a?�f�>gm?�i$?4�-���V��l4�W���1?�=?���>����_��c�;j?��'�>Jy"?(n�>ko>��������M`>�Ơ>u-?���>A ��~�m�s�jI��Ps?>rE>[����?�Wm?�!%�Z�@��l:���b��l��}�>�x��4���q��)����n����V�洚�\��#	?��?J�����>��������F�y�hԋ� �����?�>�}�dv������J��xN��۴����9>���>=�?�l�>��M?� ?� A?[R˽�>�>��C�`R#>�=֨?�4?�}>ex���[>��>�Y>��������7�����=V�ý�}=-)>m�.�)�&�R�)=�n=7���4Ͻ{�x=ƅ\=��V��"ٺ^	�=�	�=tr?ˡ6?o�J<�?�����=k�&�ւ����=-��>>#7���Q�n=��>1m�>C?��?a:>��Ѿ���#y꾮�!=k?��.?5|�>�F=�#>���RȘ��gU=�$>$ɽGe��K��������a��g�>�>�>�*�=~��>�Ut?X�C?k� ?�~��`����c� � �,� >�� >?L�>Լ>#J&>q���Z�x�s�D%P�O\B�Oa���/V�׻���>F�컚re>%H'>G+�=P����N�����_㽷箽�U�>��>��.?���>���=.w��t���O?V6��n-.���,�*t,�w���Ј=9�>|��="1?����H�QT��|CG��h�>c��?��?1wQ?����=�7>'?#��d�=��Ͻ���<�6�<�N>�� >:m�e�B��9�D�7���>�4�="a�<��ʾ�풾҂�=�����<�X��ؤ��j��A,۾�e�y$�ǆi���ϼ��Ӿ�v�q��)��U����D��B���"苾�5O�R#�?�Q�?��<�^�=�"A��PB�wj	�*�����<���=;'��'�Y�4����s���/K�y� �\k��A�Ď;�b��>�iN�����Fy�n)�.Ӽ�7>��2?V�ξ"��J��B�|=�8'>��=�w�����d隿8;�R�P?��7?�꾌Y�J��v]*>C?f�>�&>:���������>L 5?��2?ޟ��U���1��u�����?U��?�-X?J�A=�uj���z��	�!�>| E>^qL?�_���)� |L���?��I?�h�>Q1 �����xE���>���>�����=C�>4�t>�Y������T����G�=E��>pР�����B�Ͼ��<�{�>�de>$�Ǿ�w&���>]��IN�1�B�x�	�"�4����<Jv ?*$��>Bud>E�
>�o-��c���s����DJ?%;�?+UN?�7<?b�쾑����{��;4=9�>�N�>��=���!��>j��>Xݾ7nt��H����?� �?���?�g[?��p�>�ӿ젿�?̾�DǾp?8=��>n�X>�z;��󫽡A�������=r�=�)>��-<�b�>apV>�|!>�@H>�1���j-�Va�����`$�� �i���K��"��CӾB1�r{��My�����X�����(>�g�I���c��p�����<�E_?��!?/�B�.ŏ>��p�!ើp�¾Z��=����+�b������b���T������ݾΰ2�H�������M?�܂;�'�>�d?�����`=wx�>f�񼞟�>��>�:]>��>R)]>s��>�=,>�YH<"��>�˚=�~��]�T�L�o��b�G=lkO?}.��lax��l2�!)�}b�����=�B�>�<6���Ҕ�<|��m�>.WܻRSüq�a2;�z�>���>.�A��N�<�>g�����;���Z=�">��>~��=]����0.�z�9='D�>������=UW��X�?>N�?�\?�F�=���>�>���=L��6,?��>I�B>��>�i1?H?�S"?�t>�����Ý=��>T���ln�p$4��x�ҳ=�H��rj�oMm<B�/�2�]��te���d��[?�*y�<O:=���>\�=?��f>il'?uԇ��]{�IsL���g�=P	>ʫ��i�	?>�>I]{=� �>�?�#?.�7���&���R�>�@�>_�i�A����=�q�=�Xo���_?�?�-��^�N=C~�>ҋR=��f>�C�>/4?��?G�>�
o>����AĿ��;�:2� >��=��Ľ�ӾX�ʽ��3�6��yǾ�h�����޼^�h>�>e����0<>�.�>���>�=�=���=s��=Y��=}�7۩=�i=>���=R߮�/����x6��`V>��;�s��;HY=��>=��?�aR?�*��h�����˽r��!P��<�;?#�%?j((?P#[?3??@2��au�m�f�cf���
�>d�v?�x?�ɽ�	�<�ܬ�ԧd����>q,�>H�=-��>a��=�H��Aں�"?�8?�
��ȉ���d��}�އ4�T��>��=�Y�1�?��?T�/�T�Y�!����Y�$P�!��=�=���倾�����׾W��]�Ⱦ�H�I�о�q>�?���?����BI�>Kgþ<)��J���վ0�?��=b�?�ǅ>��u�\���<��yl�3�e��<>S<>`�+>Hْ>�z?1ӱ>�F�?0f?dt_?�˝�[��>�A�<���>|�G>��/?BB5?���>=(�=]��>�X&�=�F���!��=Q �Kṽ�?'=}f�=溁>L�=��I�>><�7%��v���9�=�y}��zн0�����=���<R�	?��,?T�'� <	�!�(:�����˃�=��<_��⪢<��=*
R>��?s�Q?��>4=�>���Hl��.��Fw���^?sp(?{��>+>pl�>����� 9X>��`>ٹH���/�6���v��sS����>_[:=�'=�#}>�?-:<?�O?�䬽=�$��De�{���o�=�t�<^�>���>x}E=]���S�A��#z��O_�f�'�:��<O�?!;��>Ĺ$>99>"�=�T>'��G��}G��=[��t�w�>U��>�?gIs>/��=΍�����s�F?�/j�Ň
�n��̠��I9����(>bh<>Q����?W@ϼ�v�tx���T*����>B�?���?�t?z?�������|>Þ=>v߅=�0���;�I�����<�g�>p[>�Ec�Y�I��ܻr�r=�S$>Ƚ��������$��Z@����K���9��𠾷�|�H�ӾM�)��Z9��Ɇ����=\;վ�&��b8����<�2�=����q��� ����^��j�?�3�?��=��E>��]��$h�?ƴ���=R����Y�<}y������C��ݱ�����h��0��y�'��IO�$q�>��L�����x�v��.�U�M�l
5>�[4?;�콾q���zr=�[�=�Rn=���|̓������䏽g�H?}�:?��5��������7>��?�	�>>�N>����i� ��u�>.5*?�??�=�T��T����
�}ŷ?O��?�@?埼�O3�|;ྊ6ʽOt>���>|*=?;���оR�=Z?�2?�f�=�پD+��ϴܾ�`>#v?k��1>ٓ?��V>�U������ܭ;<��D����+>��۾dѾW�!`��7}�=�8�>{W�>9<�������>���:�G��tN����I��<���>�����5>��t>��$>|�%�T����ņ���
�%O?�ڬ?��U?�/?�/���޾p���^=K>nv�>I׹=g9�ؿ>�܈>�$g���þ�� ?�!�?+��?�`?�yf��ٿD椿a�վ��׾��;���=8��>�S�h��=�0��H1=�ػ�_x=�I�>���=�"�=�>f>�}>����
*��穿x㌿S�*�ݚ��9�?R�Z�U��t辣{���`��>��_'"���Y�ޟ�����-0�<�D����<1�B?��>�����X�>��x��j���"ξ3^����̾���M�'�I��F���kپ��K��T�&������?����m>h�?�ǟ��[g>�B?q�5>y,�=rDJ��ۘ>5��>�{�>U̮>zD�=oX�>d�9>�X�>]K�<zY���j��K���s�iv�=��|?�H���9�������@�OhԾ>�����>W>H� �!���4�����>��=��q=U���9���<Ѝ�>X�$�O�>tՒ��w��d���0(;�}r>e۾;�n>������PO8�v�>�J�R�}>������,?8��?�XD?�n۽�x>����Ag��0Ͻ�?��>��>TA?CO_?0�J?X�'?c8<]ԇ�8��=�
>	%½=�=�H=?k����ҽ/�M������=bN=þ��d�?<��6>_�4=Ԉw����/��>"6??�Q�> A?�-�[|R�ɷP�W�B���=�F��m��>%J�>��R>.��>xt�>g�>��X�n�p���e��>˚�>�a��BZ�2�� 5�;^��=�|&? d?c�>w�D��2>���4���u��>��2?�6?I_�>��>���e߿���ז<��v�pk�=�>Q�,�YP/�WA�=]L�Eh�H���z�=	��=�1�i��=��>���> f�>��>��=��>�j ���I��_����ʼf�D=�x=�ϰ���@=w����~��=���<%���	v��4�
�?=�g?��̽5�����X���	 �*³>��m?�^�?/<?���>Φ���@s�\�r�Q�f�Z�?)~Z?U
J?�߽ �;ĵ���,����>���>��n>�	>�o���y��T�=I�^>��?d�=GA��ؕL��z>�P���-�>٨�=R���?�Rq?�����|:�\z��K���;J>v���c�ξE���DX��	;1���辉rM�?c����/ �>��?�2Ͼ�ԏ>�k�;av��R����bž�Sj�{K]<<��>{�<�tT�6����+�r1 ��M����={�>���=���>O%?��?�g?1�,?q�@?��&��x>�<)�yd>�d�>�j7?�[?�b�>Z��=��>�ͽ<cX=��ཕwO���a��8�=�>���=���;���=�E���;�3$�}}�9Ң>[�}=\���=�N�>�?G>c�?t�?����Z)�=�����@����P>�X�<`���6�^���>I/?>dk�>���>��>2�r� |����ݾ�J�jB۽�)?o�@?�g]>���=Tb�=�1��3Ծ�# >r��<�	)>�(�=�V��3�Ͼ�_���[>�>'RA>�~�>�m?I�0?c(?���Xq,������
�����j�U�>�V�>�����������`�[���t���:����ʣ`�]�<�*>#��=�,�>t*�=�1>k®=kb=�`�����=:�@>���>��>H��>2�x>T*?>�Jh����_�8?9�4��a��=<Y� �͙;�k�>�"k>t�.��?�T>��#�ʿ��>X?�
�?��?��e?�ѫ�Ӣu=lh=�;W�=�S�>��>N����`�>ۗŽ��~��?�=i�����F>�\�>�d={�b��ܾ���$��
"���1A��r������P�׾ݏ��{n������pS�OY��TK���\�7����$���;&=<�����K�f�}���H�?X�?a Y�Ŵ>�#Y���z�b:۾���=�w��Q7�=)�D�`M=(�̾����s�ý�"�p")���8���!�G,�>v�X�<��{�R�)�"j��r�=>�y.?�)Ǿ����l���Hs=$�">���<��ﾟ\��摚�����U?Q�8?nV쾯���ɠ޽¶>8�?}�>��$>ڔ�vH����>�3?��-?�ߎ��P��FS����?ñ�?D�G?xx�7�[�2��A
���w�>�G�>��C?#�������">}?�>2�4?E�>i�ݾ
Wt�h*�?*�>���>̴�})>���>O�=N&��ݽ��<�������">QX��^�d�i;��[ξ���<��J>z�>��־YF��@�>�M־�Q�>�K��D��S=�Bg��f?�ھ�G >��0>+�=JO�4���l�����	�7]Q?|�?�C?ܻ3?n��1���B��Fu#=���>��> ��=TE��]�>�D�>��Ѿ~�{������?���?�m�?(X?`>_�`�ܿ�æ�e
Ͼ�Ҿ��=ܠ8>�	p>�9ǽ�g=C��=��3=?�:�S;=}��>K �>���>�!0>Ό�=�B�=B���( ��������KVC���o��F����G��Z�������ʾ��(�=�;�o0�gN���u=�H7C�%�>�G?Wc�>Lێ>�]�=�y�>������׾l(=c1���	��0��پ��E�������V���ٞ���_������?�.���bp>�"D?��Y=���=�g>��^>!��>�8>�� ����=ƻ�>�y�>Z�<�����ּ��~>���=㔅�I����Y9��[��B���1C?-��T��s�7��-������o>U�>a�N>�r�p����x�lX�>#hE�Ddn� ���V�����>���>ؘ�=^���|Z�	���z��Y١=yq>��>#VZ�J
���I��E=�=�*�>�L���6>wwX>��?�!n?@}(?�R�=5֟>Մ�>p�>�J>�r�< ��=���>�"?h�?��?
�>%��=3����$�=%>��^��d�;�m׼C�|��	�t0�=�挼��>���=9sͽ��={!�=N&,�h6������(�>�5=?N��>s��>���ǋ���z��*���KR>6�뾟�>|�L>_? �?ʙ/>UT�>q�U>W�+�����+?�y�>�I������ǭ����Q>/�=q�?�VG?�E�=D�ZɊ��P>������>�$�>�G?��=>�>�h���쿗�>�{�K���%=���>���>G���9�I�o�>��>�s����&��o�=��>�=>����4��>eĳ>��->�>�=^�5<�l��xs����=!��=�Y��"ɽ;t˽��=����#�8P�3�T��m߽�5���?�b?_0��i���|��)���
?�D�>�j�>XL�=�=r���~2D�*����*�?/Jj?r��>�_�4��02>>�=*�>c
E>���>�oa;3���T:�����=	
?}�>i�?�Lt��c��~�d�#R;S��>�hu=�t��P�?�eb? �
�C� �=����6��9�Ţ=>�͏���&S������ʾPę��3#��ˬ���V<@��>^Ϣ?�9˽�ڻ>L��޸��~���bV��7>���O�u��>Y>�j�=t:%=ؾs�ᾫD��C<����>��>-�D>�}�>�$9?̒?��<?�F?�;���,1>d�#��*+?�B�>�_>Ai$?�?G�Z=�|#���К��I�)�������\��p���!>�(�=���=�">�騽��Z��WD>����s�A�<����ܼ��v��?���aS>F�>��?d?���<v��=�&��o�F�R:߻�b�;{*X>jb.��(O�1���0�R>@�>�>0?�H>W�ƾl��P*���W����>��?5��>/����>ڭ��Rὐ$>ږZ>��ʼ����=ܾ�D���Sc�$*�>�ݝ>Y
�p�y>:x?2�>?��#?Ԍ��'���V���&�B����& �9;�>U��>��=�[Ծَ%��s��b�G0�>����^q��b[�H�=]W�=���>�.>�:>jü5ｹ����J=��^;�ө>3<�>o?�;>(ܹL����E?�螾������-�Ͼ�'�.>�M>DV ���?�f��}�;t���<��s�>]X�?���?&d?H�F��&	�,M@>vj>4>�z�:�"
���伪����(>t��=��b�𒌾����R>�ޅ>�И���Ӿ'7��O�i㴿�SI�ќs�}��T�%8�����@g9�Ռ�����<��̾*w־},a�$��e龐D����%�ݾ��w�?Pl�?�M�=�V�<���7A���0���= )���<����� �ƾ�6K=qe��Br龎��3�Ծ����ն.�B�> ��#��������<�����$T>l�A?�|���l����:�W�+=��f>��	�Ap ������:�����;�y;?g�5?����K��]屽7R=�Q�>Y`�>�uy>ĸ��q�s��>Q^M?��?�8/=L���*�����JV�? 6�?�=?�潐�B����A�˾*>SE�>�?__��S����ˍ��?�M?���>�6!��:�����4?v�%?�ě�u*�=a�?�� ?	0�=_i����������#�>;z>�d�S�(�Y�9�3N>y	�>z<����˾5 �>��美�N�2I�AT�2� ��b<]?�Y� &>�jd>�>�)�>m����������!�L?-��?8R?ɀ7?L����y�۲�����=��>>�>5�=���b�>݆�>��6�r�|� !?���?J��?��Y?d�k��zο*���Y�ʾ�(ҾC->ֳ!>�Ga>
�ӽM��=[}=��%=�\q���>�Q�>�
8>DH>�>;>�p.>�F>�����&�V���e���g/<��!�c�
�n�Y��7|~��X�R����þ�'�􊙽B���h�#�p���*�pÏ�?�=��?��>�6�>[FD>P3>�;\�T�쾅=�8r���.������������Hut��f	���A�v3���$��R^	���	?��=귆=~?Z�"��Թ=U.�>�$�=/$>��j>s�*>��=>%|k>��,>��=k�>_�=�r�>�=�.��*�}��:8�[�F�6�<ܠA?�FP�QJ���84��ʾi���W>7?�RS>��&�G䔿$Nh���>��o��*w��A�����ǔ>n
�>k��=��u�͗���(��=�f^>l��=�f̼?E������)�=�[�>\��L>��>Ha#?40r?��*?5>m��>[`�>>�f>�\~=�`�=���=���>{�?��.?�/?�n�>�� >�9����>Ö�=Ù�>s�����M踽�=nT׽`u&>�0 >���;�e1>;o=�#c�Z5��M�<���>l�;?�h�>E7�>�����4��`W�Y�Ͼ���o\Ž~�>���=o�>`X�>���>c��>�z8>��Ǿ���?�>�']>��x�I
\����X;�k�>^�J?��,?뾉��>ˌ>�Ӆ=g�)�_�}>�G�>�>s:�><�l>����}�:�_��4����>��9>�9w>5v;-��@����=C�������>�,q�;�=�H]=��=Cc�>b�>wK�=�rF=�l�=w-^=i=�c�3�L=�+<L��=��^��(�ݶ=U2a=7�=�)�=ѡy�/�<���O�r�?3?P �9������u�j̾^W#?��9?n#�>���=
e,>�h	��1�2KQ�)����?�i�?��>x���s�ƽ�^=�U�=�I�>2?�>]j�=L *>��f�#���&>�R?�U>�&�>��C� �OYy��о3�>�U�=O���Yg�?�y?��,��R�=��$���5����:�>8rJ�sȽ��+��,���|��깠�
j8����:��˶�>b7�?R<����*>&�������rG�����PD�/'޽-�?O%�=�t=@`>�H�[�t�\��FXA�lh�>�>A�>�6?n�-?�s?�>p��>�����T=�˺�>+(?t�>�z�>�$?��?��6=��=��W�6�ν�'�
{y��ܼ����U�=�k5>���=��@=�7D=d�$>�/%=����M<>�3�=#����^N<>#p���Z�?�|�e?6�?9�i��p9}kνq����=hpA>�VJ>��u;�F����=��V���>M� ?|b�>sԱ�g�e������G<I�-?E�?��!?��O=�	.>���yԾL��>Z��>ǳ������[�����?<4�!���>T�B>�o����{> �u?a.>?W�$?`��A��Y���.�q�мG�3:B��>�B�>�=���[�&��v�6�Y�U3��~���Q��� =��>���=sG\>�G�=Kz�=K�;�����'={�ۼ6�>�8�>ɳ?`�)>,aP=�¢����V+?�߄�����Z2���_�������=��>�{�;�]?���������,B8��E�>ם�?�`�?�[w?��W�>�\��h�=4�> Ł>>�=�U�����=䯃��M>��>��?�:���l�=�=;ן>?��SO}��bݾ����z��N�P�L�w��U�Iu��]��됾��I�D���F*=�e�S�¾aaz�͕`�E����K�$;P��T��j�����?�ƚ?>�\>Y�$��S/��Z?�H�,�Tq=-l:��#2=��]��g����6Ҿ�⎾�Mܾ[M�{�m���D�>U�=��#��s�y�~(��v���$N>PN.?7>��ԡ�������=.P>�����Ҹ�����ZA#��Z?=|6?%�m��Wt��J
>%y?�c�>��7>SX��i�ֽ�*�>Y�/?�(?*96�& ����ϒ���7�?s��?=�R?005�ċ.��[ɾd����? =?Pt�>����v��wԾ��&?*�e?���b���x���EC�>�GO?{�G����=O�>���>ơ���UL���>*r���G�=K�>f�=�N-������⾺�F��>-O>o�;������>����L��TM�z���.R����c��>1���P�F>�)�>��սb�&�7N��(�z�R5N��t?�2�?q�O?8=L?C�[��ž,��=�]���=0p|>E��>�f���>^<�>���Z_;����k�$?��?R��?�WP?.�p�V�ҿ#����A�ˏC>ZH>���>����ͽEG�=%�!<�"���1>��B>�]�>ǫ�>��>$�>��=����jn&�̽���.��J�S����Qѿ��Ar������ ��<��i�i�v�K�����(0�<ѿ����5s3��]¾��1=���>EX>v�>�(> �!>�n�C�������y����&����ϓ������2�f�aC�Rľ���>ۮ��?G�=��>�gu��u�=k��>ֱ�<���=�>�>��O>��p>��S>0�=>��8> �=��8�׆��_��������-�pt1�����?ʒ�֤�����BXϾ�i���rU>U��>��=^:T�����g0B����>�B=j�"��e��?����o>���>Xm������=I��%�!��.�<a�'>�p�=�4��$���Fy=���>D��FB��s9Ҽ��a?]�?�iQ?��>�)?�B�>�(�>�Ԭ=����ΑH��,��s>��:?hP?�(?�<�=��Z�#8)��f��[�n�4
>8	8�G8'>!m���=�Me=.����*����C~=��Ƚ
>�a>]�@>���>��\?ڐ(?*7+?�@��N-|��-���M�����D�dK�>`�>�4"?�??��>3�>�)�=��}�����
j�>��n>�L7��G:����5>©>�F?���>x.$��־Eَ>���=���\ɋ>��>Cr�>s׾>��+>U���<ο�50��m.������P�����3�2��<0'�=��ܽ$N$��!���i>��>:�>Q�=9'=ڥN>A��>/\>`�=t�='6=ÃK<�@��[��9����|<�'��D]�pC	�w_k��۽=�'��Kb��G̼�|?@�?O̼{�{�F��X��C���6�>Pô>UH�>p�>H��=�=�w�;�iv5���F���>�b?�0�>��.�Fv�=t����@<YN�>9��>IGn>���KCT��^��a�;�N�>��?ߦ>���6>^��j�U�	��>��=,��5��?��h?���R�\�-���=������=�F�(����o��C������������K"��;��%P�>���?�#�s)�>�7��г�����������Eڼ��Z�� ?X��=�=@-b�Ֆ𾑟Z�RX����B�������g>lհ>"j?: '?l?�m ?)?֕Ծ\�>�ْ=
ȃ>��>d��>��>��#?�i>c�h>㛖�:��i�E����_}۽�?�����>�g>b�D��">.�=������=�(��7!��pX�=�T��
�M>c�>+8�Vk>��?��%?��=���=ֽoN9��n=-�~<;��Z� <����W�-�#�=B'?F�?/ً>}���LR��No��_�+�O=I	$?Tv?=D? �3=�c�>Ml��+����2�=k�>��=6.�bD���2s�.����0]>�]>��=Wfw>�cw?��F?GB?`^���cA��h�+�!���ͽ/W|�A6�>s�R>�8>6�����
�c�0W@���#�Z�����"�Q�j=���=�R9>i>�%�<;ܑ=9��c�s<�☽X�`����=�D�>��>bO�>�`>�M��v8��@�ΥV?�p?����=�޾�_�#���4[ʽۆ1?]��>;"?�5��cC�����R�]�O>��?⋳?ܜx?t���{��L=� �>���=-f�=�{*��D��t^����=n >��&�L�q�֒���j"?�#<)C���pӾ���`����ÿsm��Q��$�bQ ��'�����Y���y����F8>�I���(۾y�T��E��i���J��_ �4s ��V�9�d?��@?��J>�9=� ��o־����;�tP��@L<�h��\�tu�[�E�����{��/-��>ľJt@�(�Ҿ.$��{����;���vg>u�?􍦾CV�W����$�.��;���A�f��x����&ؽ~�a?�/?匾����׽�=>�{�>�JD>��)>���P;@���> 9?�>�ҹ~�ݲ��yϽ���?��?x�J?L'�=a8��m�����F?2?>$!?Պ�=é���B'�BSƾS�K?�o?ó�>����������ݾ��?;<?rU7����=��>���>������}3>��Ѿ򖲻/��>���:������^�:<!�*�[>��>��=��R�dyо�J>�.��Š=��/F���ľk ��0�]<U?d_��N��h{�=�#q<AbG�X���o���vؾD-*?缲?�7N?NA?�I��ѭ���b�R��=���>Uw�>)��o���t��>a�>�澟�N���Ǿ��D?���?�K�?^�?so�b:ۿ����S|þؼɾ��=+4�=`X1>�νDk�;��<�>=n�����=��>>�m@>��j>��Z>ȑz>D�>Pք��9!�<䝿����"<�S"���Q&r�q����L�NS�:(ɾڿʾ��	�B�/��Ƨ�l���߽���D��{��m�>,V�> ��>���>�>��B�$�پ�c�5�<��f������Y�������"�$��5ή���оf������2�>_5s<��=/{?9�-�%��=��>4{G;`��=��>��>i� �>�Br>=?%���=PF#>���>�\�=�,��"Y����3�'K�Zz�<B!=?�5��@��x�5�e���{(���{>��?��8>Z�������s��-�>�tm�����e���K�<ė>^��>5�=��B�sf��.;��(�Ƚ��=G�e>i�>v4���ӊ�����w�=��>zs$���ia>
a?_��?��S?E(�>s�Z>UԨ>z??�彔C�����=wHs>��?�3�>�Q�>�@�>�!W=ʘ����ѽVHL���C��\��8O <9L�>�R���ۊ=���,�Ľ۽ =�u</��������=�c>(�>�(�>i�K?c?�>�@>��]�Į@�?�����s�>�1��>���>y��>�V�>�5�>Z�>��=�,ľX���#\? ^�>��a��狿�����H>���>�~=?Gm(?��a9a� �{�i>1�c>�a�_>�>)��>9� ?܏?_�����`�ӿ��(���*X��/~����<��\,��T����<O�������ٽ�C�a=��>=��'>�E�>S8�>��>>,��=�A�=��R�U�ս�{¼�>�����녽�&�I���|м��g;T���.��:)<� z<G���?.$!?��ԗ��wѾxu�}.ھQ�?�%?�=�>A�q>��>Ӑ��[����8�"�?p?�ky?���>����D���Q.=�>v�><�b>���=��R=0+l��1߾Y�>8��>���>�z�>�=���L�N�\�s�N�>�Ѽ=qV��5�?=.u?`����>�qd9��]8�����߁>g����>��@���i�94����սEϾC�����=o��>��?�,��|>(���;��z	��Q(�Ϯ�;li���w?�Y7>�X9=VY,�C�����ᕫ��9�ǯ�>l>�3 ?P�D?�p-?��J? (�>��>ƻ;u"�>�X�-��>Z�>��?>X?���>؝�>�G�>c�;���=��|�4�|���c���y.>�e�=�o>{�����[�<���絼T��%Z�S�=��=�~=�S>dv->��?C.?"B'>��>�� =>i�L�=��(�����8%��ݽ%�>�ƿ>�0=?΄?V��>�v�˧�$��� �������>�q!?#��>���=��>��h�9>H�{�4>-U�>����U7�P}��Cא�z�o=����nR<Q.��Ƕ>�Sq?�??<S/?s�������w�@�//��&���pK>9�?��>C�(<^O ��5w�^�w�]7�c�۾Ǡ��А	�Q>Lv�=?��>m=>�w<FJ���̱�\��΄>�޽6��>�q?�&�>�t>a� �ʾ�����F+?�����|���4������=�?�r�>w�3?l(��A[������7���	?�:�?�R�?�wv?]ם������o��}]�>?3�>�@�>���=�6W=�n�9�꼯QE>^��志�Us,���>"�_>P��R�_�t��|<�;򑷿Jz:��[����{�I�W���dƾ j��%0G�`�k�ʏ��[���־h���4w��O����x�8�r�����?�̄?�h�=���[�|�&�I��S�ɼ�^J>���=j8!���=�j�=���9=��~m|���&�Q�&�m��_���@���G��/�i�ؽ��tʽ/�)>��-?�zϾ��侈�����P��	����*�Q������+$>~�g?�P0?e�Ǿ�M�,&{>�!�>U�>�nG>��ƾf|���>��&?>Y?�k��b��
���ǉ<��?�?�WD?�̽��C��RǾ-Ü<ܑ?o/L?��>5w�@������?fwL?v�>?�پ�E|���\̔> 
?�?��U�=F�	?��>���ԅV�Z~>[?о Ă�~'�=��,<i��V�kݙ����K��=Ec���v��оd��>^��G�M��D��� �/d����<c?	��D>y�m>A>s�+�<���$����� ���M?=�?�T?s�5?&���{�̽�j=D��>۱�>�f�=����7�>x��>����Uk����^?��?m��?#mZ?o>e�I�ֿ]/���/ʾ��پ�� >+��;�p>np��71>�a>^{w�b�1���=���>�r�>�`>��=���=�)>R���[�#��D��䃎��7�]����	�PV[�L������͘�J;ž�!;����k��
���_��ś��ѽ��'���.>B�?7o�>h��>�4>���>�Yy���޾hGнv�0�^��xL9�����۬�󣜾k
y��T��{��^tB�����>?Q/��@>� ?�P�=Ѭj>���>;|�=}�0>.4?>�lB�x&a�bִ>�CR>i">N��>��>�K�>k�\>!w��/�����x�\�ɾx�c�e�j?�E==�����J�>�?
�(J>�=�>��>���
8���XW�E�>`1�����ߡ�s#I��ة>):�>��!>��<$�>������=<,l��F�>���=����f^T��$�̬����>�{ ����u����M?C_~?��q?S��>��=R�?>n�>L�.��z��|�,1�<�a�>q�m?�\v?&,m?���=��C�_���,��Q����<��M�bX�=݌x:+V>����=�"�>�*=��=pN<�L����<��$>@�>4fP?�5?+b�>����{Z�c�y�����5d�%ž7?0[-?fI?�?q�%?��>W���# ��{������>�%�>�!k�)�l���;�5b>ŵE>�7?J�)?l���<܀��]H=�Vm>Aj>�D�=|r>7U�>�Q�>j�=����޿ENP�?�2�Pi�=��>�>��~�ԽW8�=�P�=8J���>�m��=�C7>J�b�;����M<f!n>#�>P�;>��<Ӄ�=KE==u.>��z=�W�<9�͸�x�
�z<>�=VX�<��:�!�X��@��(�2��=��ź$?v?;3>�������Q�l3�.ʗ���>�@�>�>1r�>
��=c� ��eP���=��SQ����>�f?r��>�H&�☜=�	���<&�>�2�>:��= ���������r��P�>��?�s�>�� �yrV�M�r�������>�ͼ�y&��@�?n?�(�9Ab�,)���6����3^�>�3�G�i�?��/,7���о �;���t
�8����?�ʣ?r�����>\�򾗻��H͙�qm�c�z<f��=�Z�>��n=2h�=�}B��lϾ�Xӻ���V����_m=���=W1�>�+?��?rS? ��>t��>*�~�}q�>�,=���>
�>>i?y:?+�?>H�>8�4<ώ������ۉ���P;�����ܚ=��>kG*>�:��h̺�1=~��<U~b������p=�p[<=�Q=�E�=R�5>��&>Mv?�U!?�/r=�=�=D<��cj�ưż��#=$�>��?=�˶�ҹ���Y<s 2?4�>���>�P�=2��%�K��Y5A��"?_*?��,?��A=4:�>7��2cǾ�q6=w"x>��͂���N��@D,�%pK�b�>�s]>�d<���>l�t?4 2?��A?�=�c����4�4@���=]A%�CQi�3��>��S�4˙��"龓f~�ğs��mJ�)��wc�����Q2>���>��>�^��q�=�
8=�P��E5�WI1=(_!>�Y�>���>|/�>�5>���=�)�����=?y�f�O����N��w�+��0r=k��>��$���"?�䬾�_�����97徵J&>-��?���?��B?*2��~^�7��=d�>��>��>ڄ��!�<��l�Y�E���%>�A���h��$��#G�>�>�<�Iv��A�����K��5¿	a�Nu�.%���d��	��w.��W�p��;^�׉V�=꡾�^�oQ��>�0c�K���z���׾Gƒ�b�?�3�?�Q�>���=�F��D��T9��w�=y=����~�q���E�����ؾ�m������^,&��lZ�L�E�>�W��2���}��v(��Ռ��M>>[�.?�/ľ����F���m=A�'>�̴<�j�󈋿nm����	��W?��9?l=쾙)��!�߽�J>#-?���>`k&>崓��3콮}�>��3?[A-?�w���������f���n>�?��?SyI?��ļ�QD�����3aU=��0?�e�>1�>B1g<'2�轠���>�X?-<8����}��q�,���?�pU?�������=D��>��>P=_��?���v�="�Ǿ��V�X=XeԺCҾ���zy��b@>BD�=k�ƽ�b���}��Z��>��C�N���H���� ���h<Ո?{��K&>��g>]">�l(����[���m �G�L?��?[lR?/�8?om���� �����=�/�>���>)��=4 �G�>h�>� �Bhq���U?��?�c�?�xZ?�Am�;0Ϳ����{��������=2 �={�p>����q�="c�<��Y���ּ���=�Z�>2)l>Eh�>cE>��C>��;>�n��J�$�ґ��/���N?@��C�
�	��]���剄��������u˾��H���8_�9�g���.�劽� ���
�3�X?{��=6ȱ;N� >ʓ=��A���I�p>��"�v��������J�މϾ�\����M���F�"c��j������?�`㽝J�>�H�>�N�=
?۟�>V�Y>�0Z>�=�= 2�>�P�=��=h��>�a�=g�>�;�>��I>a6>�����aY�q�c�$�����+�HC�>�s׾u�Խe0�2�G���b�}>�͘>��bZ*�\a��v���@.�>����ś���$��i=^q�>v�Mƕ<{�=��<)������<Y6���>�p=����&ߓ��a�����>�l�����=7)\>��*??C|?cE?�y�>N?$�>5&�>E�9M==!��=�<�>= ?�v"?J6?C�6?���<�	u�
�@�t13��j����=����.���A��B^��G���)�]G�<{��=�V��_u,;��V=���=���=���>�Tj?z��>� >]��<$�e�}Y���k=~���\9�?�I�>��>!?��+?-{�=zKd��w��V�þ-��>�P`>_�x��l^�/O�����;��=<L�!?�r`?|����?<�GOQ=,���t��+�i>	R0?88 ?�>ޟ�!]��+ۿ	.�h�G��s����9�B��=��m����<�6 �ܼὦ��D�n=���᎒>T�>$�>0�V>��>���>	�V>y�=�ɞ=�=�9�ݽ��ڽ6tԼ�'���`=�XǼm:��.5>�0�D��s( ���\�-vv���=�&?}�/?��/���9����;����Yr���>���>��'>��s>�L�>�b���5� (�o��9�9?%��?:2�>������X������>Ϭ�>��?��>i��1�����ɛ�
?3?(�(?���>�X{���q���k�~�6�ǫk=�����e���?�t?X����M�����ž�(��!�>�Gn����F������0�����s"2��7��i�C>���>\e�?��߾W�>Py\�(ġ��w�-���*�}?����?$��>ɦ���I���+_ھ(���jн�F�<�g6>�f^>G��>x�{?�{a?)+f?{{V?��,��Hx?Yt�=uB?��>�ms>�G�>�?�?�h>�2 >���>1����������"��O�	>�9�=gt|>F!�>�3>�:>o���h����g=o<e��	�<�ż(� ���i=�3t>r�	?V?.?�q��]j=�=<������������=U�޽,�ȼ@7<5��U?M9 ?���>F�Q>筝�����x[�\D=�)"?(�??y\�>27ɽ���=�۾�j⼽x)>��>-�	������^�����K��=C��>�>���=Ⱦd>��t?�e<?a?�i�<Z(�T�w�OF0��2��T���cr>�Ϝ>;�'<�[��/��,{�@�Y�
�<�� ���@�Ȍ�<4lD>��+>�� >�2�=7��=��6������ǈ�k��;�~�=���>�>�y	?'h?>�y�;�X�����F?�E�����������Ia���D�=�q;>�����{�>Vo� 
z��b���8�#)�>�#�?���?eTi?R%%�����D>�^^>+j*>#�q<ˍ-������Y�#�(>���=�f���Ր�+ɼ�N>�6j>.��"X¾C�־�?%�~?��K@�)��Hiо �1��+��z\=G�b�Ϻ��Ϻ��Z��~���� �y������(ξ+�=�'���pQ�)Ԓ?s�?_+t���.>�5�\/�.|������e�������E����ɿ��U⃾%�������&8!�61G�R��>mOU� �����z��h&��N�N�:>��-?��þ]�������='�.> f�<�E���ڊ�є���V�g$R?�%8?�+��Q����˽~X$>��?c��>_r>p���0����>�`5?t.?m��������j �x>�?�c�?��r?|��A�W���I�?->�$?���>��<W$ھU�9�A�\Jr?MZ�?A�	?H�d��K~��rF�7C >Mt�>Rd��f�>�\?Q4?"��=.�+2�=���� ���>CPm>����q�����<��>Y��>��/> ��Nګ�Z��>R꾸�N�j�H�������ɬ�<T�?{�OK>��h>@>��(�k���ˉ�w�m�L?���?Z�S?/i8?�J�����a���?��=��>8ì>��=�����>��>�l�.tr���Ȗ?IL�?���?�TZ?)�m���ֿ�O��P�Ⱦ
"�Ɐ��?�<B�A>���֐�=Q�m��!=Z$��\��=g_�>�J�>�-�>
#>��>M\>����*,���	7��΅W�pu8����^��k ����6L��j����I��2=[D=f ;������=����'᫽��'��r5?�|e>�:\=X��>��|�G;$���w�>L#U��������2�ES_��1�g������#��]�֎�1GK?QH�=� �<�v?ާ>�	�>zp?|/>38�����=s��>������>O�m>�ڷ=�D>=��>��>�d�=����.K��`�?����߾.�i?�f����^�þf�4�S��>���=���M�<�����ٛ��˷><�4�z�	=\��L��9�>L��>xݫ���۽uA<d�r��ڱ=SQ3=ޫ�=�`��>>���߃=�̳�@��>b����ѝ>��?�2�>��E?|}?O?x>�R?��%���>��<܃�=���<b�����?�A?�K?��G?�I�D���.����ƺ<d#k�
&0��ii�9¼�c<#"�����2�b�@����=>��<	�<xvϻ�E?��Y?6�F>�ͦ>5O�=3�_�W�M�m���e�:#>�b?.?>�?��?FR�>�e��6	!��˾i���6�>�Ù>��Q��@��;]>��3�(��� P?U�.?(����P��t|�X��.�>u��=���>Z��>���>38=�S�{�ѿg�4�6|h�۩޾�������ea���=0� ��{
�U��b���`�=\-?�?$��>�9�>.�>Yq�>�/�>�۸=��$>��=��Q=�~(��`=�4�}�ڽ�Y�bS�>&�Χ������@�߉�=��<��X=rb?CtG?������z�VW>�B�K:ؾ�>]&�>���>]��>�R�>]�����n�#�W����H�>�aT?_��>A|ٽ�k�=����(�	>�L�>���>�#�>�l��ׇ�.ା�zƽ,�#?�b?1.\>�B��"bg�{���J�3�3�R>�C=�Լ$n?��P?z�'��hr=f��k$���7��>�䷼8����c9�Vt��*�w���O�D��M��b�?�R�?t8��g�>����������E���/�H)�=��C?V�.>���> ��}��Eb˾ݛa�b�{�a�*>�1 >;U,>ޥ'?O�+?��,?6�?J;:?"�����B?�^:<���> F>��>��>�_�>^�>RN�>�K�=�%�>�X��R���h����]��RF>=,�>�&>��=��;��>3�>�^_���˽��ܼ7��<i�3=����<=���=!�?+�.?8�*>��d>$������i�<>}b<��l	>��	�׌�x>�~?W*F?��>��>,[:>�����a��'����;�~5?Ι6?�W �L`��(�>萋��Q=�.��g�>г<=H;�� ��BS����v=�b?5��>�{�>�p>��?�<?k\?��M���6�	�d��zD��.��e=��>���>E�4>�b�����Vg��L���D�)Q��&��*	=n��=#�>�>��w=��>iW"=������g�޼�݇=-��>�B�>e��>��=�'��e�Ӿ���-�I?`��V<���e;о#�r>�R<>(�М?�{���}�����6=�!��>�?��?kJd?x�B�8���\>�.V>�>��8<��>�lL��I���t3>Ǫ�=�_y��ʕ��*�;t�\>Ly>�ʽ��ʾ��Q�G�N;���q?�g�>����m�ľ!v������h�O^��8u��R"Ⱦhkž�.��"�������.�+i��м������!�?�w�?q�=�e>ǫ0�������¾
�ۼ3���qO�=������6�2ぼ|�����3)��Zi�G�9�=UW���>�gI��>����|��"��tb���.>�,.?b�Ǿ=���re�T�=��">��<����$��ֆ���c�HQ?
�6?��뾛F��Ͻ&\>M\?��>�'><��Z�ݽ���>ȷ3?ب*?��伇D��]���f����?�K�?\iW?� *>!�I����`c�>$�#?���>I|I>�3;��꾔f��^9?y -?��?>���ʳ����O��U�=�v,?�zX��)��?s�?.(���MQ�M��>�7ž��T�  �>j���ĝ����V�I��xq>��)>�g>Ş��uqy��>��a{P�ՕB�Eb�AA���`=@?�{־:a�=j�>I�=��"��������;��9S?��?�V?{�3?5�������ؔ��=��>�ǟ>��i=6	��ѱ>$��>�%ݾ��c��}��~?���?���?@P?@'p����c�����ؾݩ��E��Ԁ�;�t>*2���E����=厧�ڎ�� ��=D.�>Zy�>�!�>�y�>��n>�a����$���������|E�E"�T���Ы��%<�V��{���'�g��
�@�!D���=: ��Ǘ���<�������)2?vS>���=�=�c�=�>��_���E�»D(� ��� �2��Ⱦ��ᑾ"���3uʾȦ��-��]G�DJ?�Y�=��>N��>G۲�Z�X>q~�>��0>FK>����+��>̓[>q��<V>HFw=�l�>��>ϴ�>�}�=w�{��~1�Wn��V��=��5����>�;)�eҖ��?9�x�<����i��>�s�>]~Y=j�e�#X��ҽ���5�>��ýoP޽����*%=ӌ�>v�>��b>�n�e�3>�h��ul6>�^�=kuw>-C
>
M�=�0���\�=������>~3��V��D�=���>Or ?���?"4?��/?�R�>ɇ�>f�ʥ�>��?=O�G>jg?T�y?o�T?�?��=� ����A ���$�GO�=���Pt��s7�=�A�=I��3Q>�=��3�I�=�~A>Ø=	<;=��;����>��^?��>2�P>
Q'=��`�ė~� �=r4�	�����%?�?�=?̿>���>xg��R���� e�����c�>�)�>S�}�s��l��=��>�6���_M?�lJ?:�־����r��q���r�>5?̛.?[�m>�B�>��4����mӿ;$���!�E���/c���;]�<�e�M��4O9��-����K�<X�\>��>�p>��D>2�>~:3>P�>�PG>���=l�=C��;��;�!F�O_M=���x�H<߼P�hE��	�ż��W��EI�$?��=��ټ[�?�,?��۽VlY����y+оI���Z�>:d�>y
�>�!�>��f>R�Ծ�c-�+=������>Ye?���>v8���S����� >�V�>[�>S�>��d��i�ڜ����<� ?�C�>�
�>\6��F�g��z�����	�>�S��`���Ý?A�G?L}I��;�U�(�X>���>�_�� �<_NV=+J���1�yM߾u�%���=��>)�?��&�q>,@߾Z ���'���+Ѿ�����T��-? U�>�S^>�����������<LܽS�&<�i�=��?�??��P?�?/D1?(v,?>yξ,H<?w-��.��>�g�>:�>1�?`��>Ww1>\��>n����j>&G*�Q�3��� =mYk�wJ=7zA>���>��G>wk=򾅽M�&�1=	b>x��<S�=��=�=��>���>7�>1.?&=�<1F���>�A'<�����=,�׻�7Q�Kd.�".">�=UV�>�m4?D=W>��c��x������c���;"??4�$?k�>e9սl>6��2'��j7>��c��l2=h�P�JV2��OO��Ll���?�h��;*D>��3>7?q?�E?Y�A?��h��
'�� l��,��˽j��=&KT>��>&=a>�>�����p�SE�zA�8d7��#����<|>�=T>��>B��;6络BA=�L��-E�"g�
0Q��	�>�K�>(��>�3>�e>�������}I?�ע�z�����1tϾ:����>��?>t �	�?��	��}�4�����<�k��>n��?Q��?�Md?W�A�/����\>��U>��>L3<�E=�&��a����d4>[�=8oy�ut����;�]>Vz>\�ǽ��ʾ���"RR�v�ɿQ�M���ܽ$8������d���'դ�?�I�b!s���þ{�˾�z���'���N��4+�?���z抾2h��
�?z~�?3 \<2r3>}�E�?�뾇�;���<��O��m9=+Ic����fv��ms¾N�)���%��>p�(�q�s};��ӹ>a�
�}�����y�*��z��=��=��?ɛ;�ǿ�ʱ�:�&>�,>�=������\���
�7�F?��.?�-��ē�٤���_?>:�?���>yQ3=]��1��^�>6;?�)
?o/�<ZQ��+����c����?���?t�_?���8�A�R<���px>�!?�Ȇ>QTC=^�	������3�a+C?o!M>��?:M��8���3"�~(�>;tB?��X�w �=�!?u-?!eҾ�Bʾ��>�s���'X� ��=ݟ.>�!��	~�[�����>��[>Q�.>�	��\�-���>��YkL�\xG��'�����<|�?�G��>��{>G, >b�*�f���m��|=��t�N?��?�aX?&6?�������Na�=b��>T�>�7�=��*��>��>���f�p�!��S?��?s��?�WW?�i�Gӿ�
������m��=�$�=��>>+�޽ȭ=$�K=忘��P=��>U��>�o>�:x>K�T>��<>�.>R���u�#��ʤ�+ْ��[B�� �ɤ��ug��{	��y�����ȴ��f�������<ѓ���G�)���V>�Gפ��{E�ܳ(?���=�/r>O�%>w�>^E�rѝ��Y�=�E@��3ݾb8��E<޾�� �މ���[O���_��쩾^Ȏ�\��v�?�p}<���>���>I�=D�<>I�<>`M=с>�'d>|�F>�C�=�� >�Tl>+�>���>,G>���>A񘾟Ԃ�➋���q��=%�FIھԴn?Z>=�>�=��t��,����>-y�>ˁ7>@d`�=�����_�/C>+<e��>A)Ⱦ�	:�W>r�>M4-�k��s�P>���?'s<P�	�@`�9�=�	�=�#��ӻ*�� �=?�U>EG��p>���>S�?#gE?��(?�<��F	?KnM<��>���=X�-<5'����<�C/?7�X?�U7?�=+?4 �<�u���0<O#>H��4i<�伒��=�n�;;�<V�<"e�=�G�%ν~�(��?����ֻ�ޘ�������>z�,?k;�=�>�>Ê��Q�A�~�5�:�/=�v�<2�(���>-��>��?���>@� ?}w콛(�
�z�����?��1<E_D��i�o��<� �>�s#�6?{?*`?�^��6�/�w>"��=�g�>��>x��>�?�h�=�%�=��֕ӿ.�"�*!"���������;%C;�4�Q��҈;��.��S��o:�<�Z>�)�>��p>��B>J=!>�(2>�,�>[�H>暑=���=:�;LH;gpO�0zG=�5�
S<�<E�����魼r٘������F��@�����+޼;?�D?����I�5�_�����Sm���v|>'"�>Ԧ>]f�>�#�>�*���c�MhI��v�B�?ne:?+	 ?��8�U�0=	�v�;V=���>L��>��>�۽���*�����:�q�>�`?�7�>�K��5R�܁Y��Y�!н>�L���� ;�?�5?zJ�g*B����t�6�Z�!��3>���14�by
�y�Y-�_I����	���Ί:<x��>�?ħҾ�m`>
��痿i��o-�����Mq��	?=^�> �=	;����G��:�
���;4Ib>�e<��?i�?s�>g�G?�8�>=ٚ>#[n�p��>��н��>~x�>Ry%?�?��?�O�>��>�3�>~�W=��A��xm������ϼO�
>��=��3>8=���=Q?:=G�#�߈f� |�a3���l�=E͋=ֺ�=PWp=8�f>s��>[�*?�sS:���=���=ɲ�=�o�=��m�S>�%���0�L"�<�Ё>$?�>�=?�$�>O!6>�E{��<����->c+?.?ځe>��%�j�p>�f�����=�=U߃>���yݾ+~����M�i>�>�>DT�>��>zAc>�k~?��A?��!?K(�*�-��v�,^+��{ۼْg����>��>���=��׾��3���p�$�_��/�_<3�|�@�� =)�=0�>�@>GU�=�'>��;=;������`�o<��P��گ>C�>�f?��Q>�8�=?n��¤�HHI?����-�����>�Ͼ$x�5�>��;>���24?�m��}������=����>q~�?���?�c?�,A����k\> ;W>�*>*<C0?�%f�w[���'5>T�=^�v�����FB;��X>D�u>�ƽ_zɾxX�2I�:Vÿ�<������D�����#��,=+�ܽ�E��F=�j������z�ľ�~z�"��',�l����q������d�?�L�?������
>�Q�"~H�@�뾆�/;8'��u=0�������ýҶ>�p��ѽ R��/M�"�%�֡Z���>�?X�2f��6�z��,*���׼��:>�K/?aþN��R����N=�$>D�<�y�)���C��e���S?��9?������	���>�C?���>
�->G&�����Gݏ>f4?��-?�˶�1����[���Y�>�?�n�?�M?��'64�M鍾SW@>�$?ט�>ʝM>}����]�؈���<?�� ?r�>��߾�݉��ӻ��w>rY?�1���4>� �>A�>|�s�gM����=�~]�Db��a>%�=����y�7�=,��>�u>3��=�/B�� z����>��)�L�G�A����)��YlH>,�!?�h��6��=%8m> ��=���x��j=~���b<��H?]��?��o?�.?W�ᾏ[վ���N�Q���>�*e>�	>����O>�Y�>�4���a�/����?@��?��?��Z?��T�?&ٿb���שԾ6����cH=�Y+>�m�>��k�!?=�.��\/	=�����<���>=� >܃�>t�,>���>&!�>������)�p�������eh5��w�:��g3�b��P�;����%/���@��.Z8�ό���4��"�۽��U^�� f���FF<hgH?�{7>��[>�U>�Jc���Z�O,�>���Z���'�~�ݾ	Y���/��G�};��¾#�S��N��� ?��0>%�>a��>�)�ߍ{>p?:)v=�ߋ>�!_>{�R>~�+>�=�>��>��>�>6��>{R>q�q�i����� %~�'[P�B��>�!���Y�B�R�W."�m����}>&�>�͞�y3v���\�g�����>\±���{<�x,�-�r�NO>��>�;?�"��<Ҡ>���j�5>�[�=5�>u�#>��8=K6p�2��4o�׹�>��]��9�>{�>xQ�>0R?��|?R�>T[?���>�l;?l�l�D�)�4�-�F$�>��H?�o?��]?_C?G<=7�����D� 3Y�4U=��:�4�f=�l>�@��ǰ��%��t�j=�{@>EO۽p���I>N=�"��n��=?�X>�u�>��M?�_�>`�>�ؤ<	Q����z��T��J'Z< ��-��>��>.Z ?z�>w�?��?>
a~�kW���u�lC�>�Q�>��������?e0>
,�>&:>ڎ6?�rL?�籾�־�K*>���`�>�??>�>=��>Wd�>v��gc�۠�%=5���R�"r��4$�='�R>KK�<�M����j�	nU����='����S=�И>�"�>4!�>��>U�d>��>��=>��=ҵ�=@�=���B ���<�W2�T,D��F=��<��?��Ml��"+�ڊ���޼�"���i	?ea?;�=���9�I����P�o��V�>���>i�?��?���<�@���J���2��:��?b(n?��?N7A�+mU=�-h�� �<v��>GP�>}!c>��'< �۽�!_��hU=+��>�~�>I�t>H(>�h�`�0i��~�	T�>���<C����(�?�gT?��ݾ+�Ⱦ)�8�$�^ �]��>�\�N6��B����K�����p~��K]��29�=�C�>��?�yܾ�d^>����Y��5�q������� ��m?L�I>��S=�s�Jپ�X��l�d�|a���
�>~W�=��>��)?�3>?2C?8?�?�>�����1?�<=��>~w>ڛ�>�?zb?0��>�4�>�5�=��v�u:�Gf�a�='�H>�+J>��^>?���f�=+�>��c=E9
���T�4ơ���D=�h;>,I�=w�=��[>�% ?%?ץ:��V>ɕ=r"�m��B�<���B>4����E�f�;���>�N?�?@e>vJ8>��۾�Ѿ!���"H=�SC?�/V?�CT>�(�=�w�>�N۾.�>���=K��>'`�T[n��ѥ�J�������n�>�4>��q>l�D>�Yw?�P?��B? qr=A�M�Vny���F��\���{/�'V�>��>B�>�)���f���Y�wne�s�P�'��<�tнC2�<���=��=�MA>M��<�c佲;�=�~W��Y����=�Y$>�)p>ňm>(��>�C>]����&��v
̾d�G?%᝾z�����n�Ҿc�%�$>�RK>!ս��?���K{�������<�'��>�j�?JX�?��e?�)����߶R>�"Q>fm>,fw<|H=�J ��U;�,�7>�z�=�.{�:=��^�<چX>/�k>ٶҽ�����ܾd�8������M�X!9�����`�ξNb��i�*������L�scw�2�q��J�� ��H���'ͷ�`��>����f)�%D����?A�?*�=:y=�zB�]���:�ѾE�'�����V�	������5�w��~ܾwܕ�]���*�%�H�l\j�m�>���;���z�]��E=��=�%?�R���ѾO�#� �	>�I>	�=���B��Y����R��U@?�6?�Z��K�Yۢ�T�>I�?6B�>�
<	��uX!��N>�(C?1l/?�=q=v.��?���o=�Y�?���?�m?�0)=��n��߹�>�@?l��>	9��������4I��?�ZD?Ir^?=pE�mً����w��=
w�>�1�U��=�N�>� �>��������!=Ф��H0)�>fz�=��!���v���j���=��B=��Y>�:I�*��)�?�}9���F�z�5�zuZ�G0]��R�=B�?�@��mjP>`e�>�!>�@�S`���n�8ZH�ŊN?�E�?y?���>@Q��W�D5�$�M�e^�>���>-;>ЇH�B9�>��+?�'��o����,���?���?�z�?Z^v?���S!ӿ�蛿}{�������=c�=��?>�޽��=�M=�����6���>���>��o>lx>�6U>��<>��.>������#��줿�В�*B�������\g�@	�Vx���K���Rս�8=��^y��>���G����/?�!gh��u>qͣ>��?�$�>��>Q;�=�絾������������0پ�u��(��Oe�E?�(���	��Y�뽖��� ��>2$�=~$>E�?
{ �'F���Ȫ>�	�a�>W��=�4>���>X�/>��i=y��=x*�=aO=�PA>�E�=����؊���P�E�)��X2��)d?9I7�qsž�>�[�5�&y��B��>V�?r>���e���rqZ�ؓ?7���Z}��>��b���>e��>�h)�K��=��[=�%���������=�4p>�D>����!d�Ń!�c3�=Nߣ>gʧ�dx�=���>ʬ4?w�L?��R?��9=�O�>�C�>��h>��&>��u>Z��>���>��?�9?Ƙ#?&'�>r�i>�g��du���M˽������=O�����!�U*l=�l�=�7:��Mi=��u=A>���<X�4�_��W&�R����;�>aK?�F�>?�ǩ_��X�{�5����>���>��?�4�>/j$?��"?E�?3��>�=E� �A�ER�>O��=�BE�ǜw�CKp��B.>~����#?Tm?:I�=̇�@�>&�<dX�>*J%?�wH?T-�>��>��=�����ѿ�#����0�G��#���M�R=���SL�c��<�3��K'���N6>a�>�%�>$��>k�I>��>jV>R|�>Z�J>;]=?��<�7�<� ��H���-��=��;2�;��
���bڽ��;�̽��f���g��=�H�<;?�<?jȣ�_�Ǎ��'"�󒩾��>���>�2�>�y>n�=	��a�7�>��j�~�d��>��D?.�>D&����">�B�pz[?�{�>{�V=�"��
�׾��.���ؽ���>�_O?�d�>Q�����n���C2/�,E�>>Nf=�����Ґ?��U?>�Ǿ�����$�7�W���.���Z��	ýa4Ҿ^��T�,��]��M�����짰���D=�}�>to�?�b���#�_������\��������Q=W҃>.�������'8�p���쎌��ؼo�>��T�>/o�>H*?A�[?�<!?�X?�BȾ��?4o>�0q>�>��?ͳ7?e�?�><�>��Q<t�<>s��<٦�MX�=1�N��f=]q�=�I�>93'�􀏽d�a�R"=i.�A��w
����B�fyS=.�>��.=ո�>0�-?-�3�C�q=_�N�ǜٽ��ؽ��>H��>��Y=ry�=v>�>��>�?4 _?�,�>�,4>Yy�����7��+��B,?00??��>�l��ͩ>�L�ߗ�����uW>��p���7�t�ľ�G���w+���>)�L>�{�=fˇ=8+~?�xx?���>m�t����򞌿Z�)��Q�U�����>���&o㽝��٤p�6ǃ�7�{���\�b:&>����$u=,)�=��A>�#>y���Gb>�!>��-=Oi>��<�NX=fc�>��?��<?s��>�y�=Bμ�h���]Q?$�޾[��@�޾,��<-��6�>!��>S����?�>qR���~ƿr�o��b>>{��?��?�b�?NV���ȶ�2��>���>s�]>�M,�࿾����	(�li�=#k�7��9���?P�=i��>�D=��-��v�V>�S�ѽh���c�B��&+������ܾJ���sA=������/�2�҄*<�{��	�>Y�LC��H&���O�ڒ����?��?� ��ؐ9���5��9���:־��>�����.g��@��)� >������i��$������������?�>�x޾+�.`b��XH��8>�ak>��R?��n�[ "�gD��u>��
>ݓнˈؾ�ᖿޡ���%ƽ�k)?
�`?�EZ���o׈��[�>�h+?�|`>R`C>���'=d�>�Q?�	$?�������l�m�V[�0܋?�"�?9CQ?e��}d����)��@?JN?"��>�Ȃ�懮�r^�C�$?��$?��v>��������$����>h~�?i�'��I>�?�H�>#�f=�u�87ȼr6ľ};9>�L�>%�*=��A�Kdv�����Ƽ=f��><�>��=j�:���?��&�8k���)��-��r��Y�=�6	?*�(���=&,?�h= ��f��A�����*^?�(�?��?V{�>�˽C*��3U�ƾ����&>c�K>9>�������>1�-?nJ����3<d�j�?���?HH@�fS?�K����ٿj���kf���H��^˼�a�qo>�'����<=��=�Z���4�ٌ)>��>粔>�>>^!>xJ�=b�>�Y��%��#:��������=��"�� �=Ur�,�rjr��־O9��ɛ߾��v��!>��=pI�3C�<6�k�	Y>c��>(h?���>a�>��>�ʼ��1�nԾi�o�r�j�����Ҿ$���Y�f�ý�G$���U�Ʊ�V����!?��;�}]>��)?�Mļ��ֽ ½>�"X�4�>��8>.�K>�w>�0�>sr�=�R7>5G>��[=�H>��U>-�����^�{K���վɦ��~?��=�� �+�=��l=������'>su�>U�=Q*?�sRO��2���p
?Q������n>7򐾋DW>>�>�H>,��)�I��g�"��{5=`j2>�כ>@/4�����baJ���D�j�>yǾsH>���>��3?��o?c�@?���8<�>j:�>��>֢�<@�>��S>E�q>�?V6? -?��>0�	>�倾�Q=$��=̆���ܽ�ꁻ"���g�2�*��=k��֊�W�&>��f<V#����<ꂾ��Ϊ��@�<�p
?,8N?���>�2�>wꢾ��{��Sa�`��=��#>�b^>C�"?00�>:�?�,?*c?Z"x> ����ľu�K����>`�0>4fa��I���i���>����(2B?L(R?�9v>��/��3_>ev�>?U�>k��>�b?�,�>���>�a<�����οpl�f�L���x�)zT�#��=ĺU�'y5=jp>F�V�{:S���d<G�>%}�>W4�>��n>&�=
\�=q`�>P;p>�%
<��t�>/7�=D0��K�=���=�W�<:�N�&+]=� ��ĵ5�4�K������˼c�Ǩ뽒??1�?FI�������Q������ ���4��>��u>��>?�>�M�o����W��?�a��u2?m�Y?L��>�	����j>|j佂��={�?�I�>�`�>�~�;|ಾ� ���j���>��T?�^�>�􆾨�z��w����A�%ѩ>��=�lν��?m�H?A☾�i_<�U���L�<�L�o���0�=�����;=b���N�8���k��t��_��;'��>?s�?�tb�K�=��ɾ����n
��I����<=<�;Y=֡=�շ>��(�~=�]�#�>�侓巾3J�<�j�>�6=^�d>?B??>�?��?]�"?(8���>?Qڥ>�M�>L�>sx?k� ?�?I��>Ux�>�(=�k=7" ��Da��'�4�*���<��=�PD>��?=�9�=&�<�8�=Bv��){�߆1�m>н*����:M7�<X�=�8?��?Q�p<*�`=��F<��(�'1<S�]>��>)x�>����x�>��?��6?7�9?�9?0��>�갾W�S�L��q��?F�f?���>ȇ��4�>�����ҾV�><(�=K����
I��NF=�}b�g��6>�^>/'4>�Po>:��?�!\?L��>�Zp�OW	�Pˌ��A�n:G���>�߶�L���~�̽d�@��a�N4������c�6��>>D>���=g�P=�4V>��Ѽ&4���>|\>L ��/l\��a=�;���U>���>�e1?FG>��<�h�����Q�O?�(��5��@��q�%�"%��|>	��>[?Q���?�A/>����yʿq�m���)>��?��?h�?˽������>
�>2�U>4�Q���i�!����L�>��3>E��Lބ�G��mp<>�2>����Gվ�4���A�+$���E*�_̐�*�2��8G���ӾKȼ��<k�_��ԽD�7�k��ةy��B�V��*ڽ����%ɭ��2ɾ�5�?/�?����lN+��_�Z�
����W>}S&��c���L����>�oU��ٜ�F���a����*��Ͼ�����?$����	��Z7���:��>�>��>���?����6���E0��P>b��=��=�Fu�d����]������?RrL?_�G���Ҿc� �q;??M?���>4�=���Q$~<�!�>	?�[�>&��=�뗿DGs���,�o�?���?5�Q?AӾ|a���ݾݬ}��?�l?A��>�;J�ܾ�>%�[�?��,?���>����b���'��?֘�?�Q1���Z>*+�>�c�>H*��~ɾv"�����Y��<X`>���=��6���~�������>���>;��x���^g&?�Z�=h��r�,�<�m�p����"?
˩� �>~��>��>�"����4�q�!�ν7M?�7�?���?�?�¾@���n���);���><(�>yA>c����1>w� ?�=�FR��,��i�?2:�?i�?EQW?7W����޿n��®��O�;U[>�=��2>d��u��=1��<Z�;��=@�V>:�>ke>n\z>�<I>ӡ7>YBN>4>���\!�����&���P6��#�&���C�{g�+L��!��z����a��|�ڽ��S����ZR�Q��.�͹�Ե�GsM>�1�>�{�>��?{�?U�=S�þ�/!�)���"����;�ܺ���e��%�<��ޙ��y�u�;h�Y�0���x"?1(T>�(%�l�
?�d�s�}>�?�:C>=�;>?�>�%>��>��>)8">uͺ=�>&�= �>a�������R�'e`����t�=/aN?�%J>�����A�j��Q�l����>}�?�'�>`12��a������Z�> ��J���A>ܿ!�M��>���>	[�7A�=�,=�e}=�b��>�N�>�S5=�<5=��)3��.>���>�����*>ܦ�>�5?��?�&?���=�8�> >N>�ہ>c{�=.�>|�">]ג>V�?\:5?�� ?��>XY�=}����M>�	ټd}�L숽�}��&"���%���;��˽<*�=��<]&A<V=�hG;սԱ����R���?��2?m��>��>_}��Sf�y.5�=Ȇ>�r>ɶ�;���>�5?�?+��>��?���;�����3��о��?�Ӯ��a|�w������	}>n�g>YR$?�p?��=�!��x7�>v�>��A?xM�>�ri?^�>�f>�U����ҿ�u�2)2�N#߼Ɔ�|�<=hM��`C�T�$���t�����t!�=Sk>�3~>kI�>�]=>�>r�+>���>X�p>^�<�X/<0�ӻ��C���V�|��=\�ͼzg�� �[�<����;�ͽj	M�(N༎������r�u�;�?��?PZ����2<�`��'���Ԛ>��~>�@�>8f�>ƙ<��X�:X=���G���>5�Y?�A�>�|w��G.>��q�Kx2<^��>��>TH!>��޽KiJ�d6��O��=#�>7*&? !m>Z���+Ih��ځ����w�>�ѓ<)�{�?u&n?���������3�Z���@����̻�����R�%�CT�(��L���v�%iF��&�>Ӊ�?���G=�N��>_����������}����L�`(�>e�u=�S�󜖾��J�ʓ��'z��[�q���?�/���?%�C?�w?)S�?���>S�r?��#�4�?�F�>��;0h�>j�:?��[?A�?��>�x�>���=�W��Q��Ũ�Bw}<J1��Ƃ�=>7�=���=Y�=�=C�=�:�]}<�<s�RЏ��ꩻC��7t�U'�<�0?��,?����ԙD�V;�<�y����=���>>P1>J��>�{M>o
�> 7?
�Q?��I??�wd>�Cc��־~����>R(?C�"?��?`_`���<ؿ"�@깾4�R��X[>�7��[���t�������T���>l2�>�?w>���=is?L�b?���>(褾!=���6���1����c�f=�>ϵ����ۻ��ɾ{���^��A"W�ا�.��>��ս��<,x�<d?2>��=𭽊v�>�l�>�G����->(��<Ed�i�>�F>��)?���=\��<����(�ѾJ)M?�b ��8�^���.�<e�=��T>���g=�>�K�C���{��eoE��)�>��?{��?'��?|L��a������>T��>�I>6�����ӽ���,g�=������ާ̾\ >���>�F>{�|��c���
5��B�7���&QH���U���1���m���꾌����d̼h�Ͻ3؍�#�.�u�.��`���.��N�tɖ�9��:���?Ѿ�?�K�?�н7�ܽ�P/�]�3����:iU>	lf�4�k�?���lڽ�U�A]�+���ZZ����B�T����%��u�>�Pw��䡿�`'�;!B���ۼ�=��!?�<����8�z��T�<��=pb̽�F�c���oؠ���@���a?ƴI?\H�X���-/��<�>XM?{�R>�%�<���0�S>s�d>5�?7w)?�<��J����{��QW=��?�-�?څH?�	���J�����}�,��>RZ?s�>��f��q��Q�����?��3?\8�>& ��W��z����?,�m?w8��D>� �>�M�>���M���#���~�(�m(H>�;����CKq�
1���
>.�>Hb�>��+��г�~�?ߴ%���t��dM�m䟻�-R���-=V5�>J2�����>e�q>�D	>�J� )���S���Y�7�K?��?Ċ?��?�O�,9l����6S=�>�+R>;s>�Q��
{_>���>�n����'����"?�}�?MR�?�dR?D���Aӿ�������u��l��=%_�=��>>�߽��=P�K=�f��w�<�c�>��>zo>_>x>��T>ǜ<>��.>F���-�#��Ϥ��֒�kTB�������dg��x	��y��������i콾}q�����֓�6�G�|�P~>��Q����3>&�?���>|��>�W�>�;>�G��!�Q[��a���8'�8�����W��]�R�z��9����U�=��+��&�> �=�iA<B,�>�9�=uC*; �>wa�<+�<ag>.�H>h�">�t%>�oY<>�D<�\3>��=��W>�L�=�r��")~�vT��^���e���I?��׽����K�7�.ܗ��N��H��>a?��&>�0&��뇿mi����>���g���:�;ӽ�>���>|��<A!»0�=���B�u�=�<>lq�=�lP��m0���x��=3?�� ��\���>�&?�c�?�B?K�<\��>�>��?�!�>Fѝ>ɒ�>��J>>�?\\-?�/?��|>���=AܽQ��R��ՄK�$y�3�����!|��<ϥ�,��t�=a�սB˼��Z=��=H"����<i��=�s?!.?-l�>Se�>�ө��ŀ����0�2>ւ�>P���ɑ>�K�>�5?�^?���>YQ�=�ࡾ��!�c���
�>{v�=�q�/s�����u��>��=���>�_?8`�>�N���KW>@ >v<6?�� ?Jy@?3d�>/�[>��r�\��*�ۿ p�^6��r뼾G���,>	����l0��V=���e����=V6\>iی>�Y�>js`>�L�>֘r>�+�>�:%><�<��%>V�½b;���`�=���<���9�~[>9X���~�>4��2H>��C���M�f�2�rf~=~@���9?}�?�JK������f��=��:���>���>.[�>��>�2�=���&QN�~�;���A����>��h?��>��F����=����֩�<��>%��>
�>�;)�;�&����:��<U�>��?�ښ>��
���[�	Fm�~����>eI�<�����?
:`?Sþ�M������F���� t�w�x�U�L_�*�H�'�=��c����1Gվ���<�>)��?A�p���;s/(�қ���&��}����Չ<�9*���>�Q>P-<>��bb*�@O��3���->�Ұ>0��=��>@F�>�H>?	>D?��>?��0?}`o���'?�H>]?���>�o'?e�'?��?!A�>���>�V{>Y|��bŰ�O�w�"N�=�߽6r�=���=`�=��;,-�=�r<vŴ�����^�=T�*�M�н��帇�S����o[>՛	?�QM?�-�CO\����l�e�������>:$�>��c>^|;�>~�?N�?? �2?<4�>��>6r�=�3����-��g$>f0?��B?�?�%��XjO>����j���:g�ɷ�>̙�ce���!ɾ�����U̽&�>]�>7�%>Y=�<��s?��g?P��>Ǟμ�����l�3�,��,Ծ�Ӿkχ>�ơ�Z����]�q��$����sJ�giw<$=�M����ا=�GS>���=��^���=W��>�޽=�J�h=>��5�7��>CQ�>���>��*>үO��'ξ0���uO?�@�P����)�/��/=Qg�>�HE>���+c?��ۅ���\��$Z��N?H�?�\�?7�?�����Ҿ���>
a�>�XN>�/���Ľ�>Ži���� ��RP������m����*�9�w>|g�=E~z��,FQ���c�0����i�8���y$��R��q.�"��z�I>e
��C��"5����<���� )ýU��m����9��rn��}�?9=�?����������0�C��h�����W>_���l��֠�׊�<wù�i"��
���4H��X��a!�<V󾥮�>j��"���C�U}6���Z� J>��?~�6��þ8�ڎO>h0�=��v<[���^��G���7"��X�?�e?\�+���%��n��H�>$)F?���>�$>�����!>���>xR?"-P?yl���ό�&�}�:��;�?y��?0@?��Y���H����b���>��	?���>s5���E���m�F�?O7?E��>�/������g����>z,h?W�8�v02>���>�C�> n��򕾾`t�C������N�J>���Ó�V�v���V�|<�=�Z�>�x�>`�1�Bu��^g&?�Z�=h��r�,�<�m�p����"?
˩� �>~��>��>�"����4�q�!�ν7M?�7�?���?�?�¾@���n���);���><(�>yA>c����1>w� ?�=�FR��,��i�?2:�?i�?EQW?7W����޿n��®��O�;U[>�=��2>d��u��=1��<Z�;��=@�V>:�>ke>n\z>�<I>ӡ7>YBN>4>���\!�����&���P6��#�&���C�{g�+L��!��z����a��|�ڽ��S����ZR�Q��.�͹�Ե�GsM>�1�>�{�>��?{�?U�=S�þ�/!�)���"����;�ܺ���e��%�<��ޙ��y�u�;h�Y�0���x"?1(T>�(%�l�
?�d�s�}>�?�:C>=�;>?�>�%>��>��>)8">uͺ=�>&�= �>a�������R�'e`����t�=/aN?�%J>�����A�j��Q�l����>}�?�'�>`12��a������Z�> ��J���A>ܿ!�M��>���>	[�7A�=�,=�e}=�b��>�N�>�S5=�<5=��)3��.>���>�����*>ܦ�>�5?��?�&?���=�8�> >N>�ہ>c{�=.�>|�">]ג>V�?\:5?�� ?��>XY�=}����M>�	ټd}�L숽�}��&"���%���;��˽<*�=��<]&A<V=�hG;սԱ����R���?��2?m��>��>_}��Sf�y.5�=Ȇ>�r>ɶ�;���>�5?�?+��>��?���;�����3��о��?�Ӯ��a|�w������	}>n�g>YR$?�p?��=�!��x7�>v�>��A?xM�>�ri?^�>�f>�U����ҿ�u�2)2�N#߼Ɔ�|�<=hM��`C�T�$���t�����t!�=Sk>�3~>kI�>�]=>�>r�+>���>X�p>^�<�X/<0�ӻ��C���V�|��=\�ͼzg�� �[�<����;�ͽj	M�(N༎������r�u�;�?��?PZ����2<�`��'���Ԛ>��~>�@�>8f�>ƙ<��X�:X=���G���>5�Y?�A�>�|w��G.>��q�Kx2<^��>��>TH!>��޽KiJ�d6��O��=#�>7*&? !m>Z���+Ih��ځ����w�>�ѓ<)�{�?u&n?���������3�Z���@����̻�����R�%�CT�(��L���v�%iF��&�>Ӊ�?���G=�N��>_����������}����L�`(�>e�u=�S�󜖾��J�ʓ��'z��[�q���?�/���?%�C?�w?)S�?���>S�r?��#�4�?�F�>��;0h�>j�:?��[?A�?��>�x�>���=�W��Q��Ũ�Bw}<J1��Ƃ�=>7�=���=Y�=�=C�=�:�]}<�<s�RЏ��ꩻC��7t�U'�<�0?��,?����ԙD�V;�<�y����=���>>P1>J��>�{M>o
�> 7?
�Q?��I??�wd>�Cc��־~����>R(?C�"?��?`_`���<ؿ"�@깾4�R��X[>�7��[���t�������T���>l2�>�?w>���=is?L�b?���>(褾!=���6���1����c�f=�>ϵ����ۻ��ɾ{���^��A"W�ا�.��>��ս��<,x�<d?2>��=𭽊v�>�l�>�G����->(��<Ed�i�>�F>��)?���=\��<����(�ѾJ)M?�b ��8�^���.�<e�=��T>���g=�>�K�C���{��eoE��)�>��?{��?'��?|L��a������>T��>�I>6�����ӽ���,g�=������ާ̾\ >���>�F>{�|��c���
5��B�7���&QH���U���1���m���꾌����d̼h�Ͻ3؍�#�.�u�.��`���.��N�tɖ�9��:���?Ѿ�?�K�?�н7�ܽ�P/�]�3����:iU>	lf�4�k�?���lڽ�U�A]�+���ZZ����B�T����%��u�>�Pw��䡿�`'�;!B���ۼ�=��!?�<����8�z��T�<��=pb̽�F�c���oؠ���@���a?ƴI?\H�X���-/��<�>XM?{�R>�%�<���0�S>s�d>5�?7w)?�<��J����{��QW=��?�-�?څH?�	���J�����}�,��>RZ?s�>��f��q��Q�����?��3?\8�>& ��W��z����?,�m?w8��D>� �>�M�>���M���#���~�(�m(H>�;����CKq�
1���
>.�>Hb�>��+��г�tʷ>m����O�A?I�7@��l�=AX<:
�>�󾴅
>a�f>�>M�'�I��zI���h��&H?:��?�>T?�w4?R���'뾃'�����=/�>�b�>>�=����Q�>�4�>�O����p��Q��2
?1-�?���?�Y?�j��6Կ���Oھtzʾ�|<�1;���=4�B�L�x>?��=N��=���>r��=���=̅F����=��c��m4>lq�>�g��#�CJ���5��It,�V'�ö'�����!�C!*��.��ak����žnGf���n�wq��u�v��Ъ�8�=��E���=��6?���>��<>�BC>e�<��)����a3�p]Խ�t���Ⱦ�v��lY��?R�{���SAu�u(Ѿ;h!�� 
�!��>N�?=�Q>���>w��=.Cy=�>z�'��E>v�=#��=�D>\�=�	A>�u>�>�!0>Ą:=�Eo�j��R����>����G�Ό�<<�A?mN����ݓ��
����%��Ae> �L?z3E=�B�L�J�v�*���>� �n�½�%L��>� �>v��>j��=2TA�M|�>���;5�$�A>����>�Ç;�x�� ������ܽa�>�X�����=���>�/:?�p?��4?�Z��9��k�=ق>c�=�j�>��=�+8=,��>�C�>9��>�C�>�cx<�䏾|�0�vI���Ž(Q�=��Q�y޳����; �=-Q��o	>.�8������ �/�:�y�=OT-�p��Z�>I\H?9|�>%��>�6���K�q�S�t���}?5���%.���`>�k?���>7b4>$x >Où>_%k��t�����>���>�+M�e���\}��M��=Y��<�cT?�;?
>�%��|�V��==��><i�>-A�>n4>:��>1��>ee�ːʿ�2H��U�5�.=rF>�Ő�=��Ͻ���[i���M��%��q�D=��	����>ˍ>Y���ǒ�����>�j�>�O>J�����=�n�=�"�<�B=�b�=�>h���U���m=������a��=��>Ph��W�����=��Y=�?{Q$?Ԅ;{kv��M�����eT��wT?���>Y��>m��>��]>t`;n�L�4��'Q��,?(C?�9�>H�������\������>'v�>1�>�i!�'/���p���=.��>��>��>��Y�Z�L�sWX��Oپ�d^>���XK����?��'?'��e��2�)���"��U��|�ҽ��6>�䰾2� �?�辎`徉����ܾ�������$?j��?b����?ں�i$�F���א��=�qL�>`%��?+�)ո>�"9=������羟C�����>7�>��u>6s'>,�.>B?,GZ?��r?f?�F ?PNK���>�cT�y�f>P��>��,?9c�>�x�=�M�=?��r=e�o�uH����}ٽ}h<��>D��=�0�=�p:=̿��uᇽ1��=����@���=��
=�ǘ=E�T�W�л��½�U%?PG7?w Z>[ ��ƜǾ+_�
�m|!>Y@�1_�>�gg��l&���O�P>���>ɉ?��=�k��T���ľ.mF�l�>?�NW?�=�>9�n=D�>��پ�8x��@B�w��>�~d=�R�q����콪�l>��r=��X;�f=;o>'�|?0�A?[�?���0.���z���"���Mr<Q��>`e�>T8�=�aо�4�Nn���_�=+�����ۊR�F(<��$>g�@>%�9>dq�=�>>��A<e������ })=��`����>�>!�?�@i>�Ί=��� ���I?y�����̂��5�о� ���>�,=>���0b?��
���}�;ԥ�=�6-�>Dh�?Ó�?��c?y�C�N��b]>r�U>QZ>G�:<�P>�CG��e���3>�1�=)7y�-������;|8\>ثy>�qɽɲʾ����)C���ɿR>o�Pľ4d�=!�|j��7�a����T���l��/�l�6�`�9S>�'*O�jV1�����8���-Ͼ{����?��x?�E	>v�4�����8��s羙�w=�%�T���e�]�׃[�`���������^d����Ծ�-4�M�3�1a�>RNc��tyz��"�
U�;#�N>@�*?
.¾K>������T=FE>z�=<�P��Gy���r�*�S?s�7?��$�˽�'>_ ?U��>�{%>"]����w�>��-?w�,?]�-���!���ǝ��;�?�{�?��)?�D���3��8Ⱦ�ή=O�8?{�/?��;>,н��3U���!�>m��>&�
?�����Ì����=�>��!?��28>��>���>l�0�z�̾�3����C�,�=i����n���e����=:P�=�m���Q>LK�>�,�==X�y]�>S�JDO�TrH����S���<�P ?�I���>�Kj>l
>П(�Z����`��V_�nJ?�3�?W�S?�U8?`��؅��i��D-�=���>�Ь>�V�=a$�J͛>ʤ�>�0��s�r����?�/�?���?��X?9�m�&�ܿW��k�Ծ�;ɾ��=�l�=6�`>�k��|4�=�S�:�W+;XD��q�=�+�>�H�>�jJ>��=Oe7>��M>炄�p��=��I���>�p������#[�F~��M�X�;��g̾;�侼��Q>�>ͽGK����s��2{�t$�=J+?�t�>��
>��>�ȹ=,'>4�ξ?������z�*��s�����&1�O�A<kI�%I��"��¦��;��J?8��=�x>Y1?
�>+2�>�� ?�@��!�Z�R=�+�=kr�<�k>F`A>�q�<�s�>�f>���>p�>�?��w𪿎�T�A����.���?�����������۳y��)��
��� ?���枿�ė� Y�>���Z A�����%��t�>M�z>�N�=7V�����=WH3�G1���O;=�Ї>Q��=��>������q�>�u�>�C����">st�>
�p? Z�?�uS?�%")>0�'>�V>��<|�C>G>qS�>9D?>��?�oL?72?5��o���h#��V�=⯥�;7�+�=o>p\�=lK�S�����g�g>���=u����֡�J�<XG�=��?:K?�Ie>3�z>�o����P�o3?��=M��!(>r^��i�3>I�+?uoI?��?.��=~s���e>l࿾����>{�>:��A��w�����>���E�?�F#>�*�=��Q��
��#�>ze*>�Ɉ>q�K?�8?��>KRϼ�8���ÿ��D�S��1�U���̾tb�=SXؽ��m��2�>_�����i�c<���2>�>�亽L�c�K�`>��>��>��>���=k_= 6[=�U=�&&�m�����b<>�L>��=��Ľ���Kh��½����֯�u�J=��S=5�?y�?X䐼JA<���7�r�F���{�>�y�>��>�m�>X�*=c|�D��U.���,�|� ?m?��?��@��#�=�&�N;=�y�>���>zm>T04�:W׽q	���g?<�	�>Lo?
ϝ>�� �|�T��k�$��VM�>
4/=^7<�΁�?�B?q��+���/�"��������?�<���-���q��:����s�7�sl��0_��L	?Ԁ�?���4�->�Ҿ@���Z��7u
�mU���1�'�4?���>R6�<�'�>�־�`�i�o���=+p>4Q>�R�>�/*?!YU?:��?^� ?��?��\��c�>��2>Ih�> +>�{>)�>4s7?��>'Q�>Z��>��>�t������]�F=1q�<�#L>��g>��k>5,J=$��1=Di�ҕH=j�~��~��k�&<����uZ��!E=O�=�"?�??? K�"�����Y:�hd���ꔼ���1%�=�Z>'�-��i>|�>l'?��=?-�'>�+e�w#}�l����l��1,?
C?���>)o�=��>zS;����!�<�T�>�������a�����*���;>҇�>�N=Шg>S�}?��B?�#?��Y/�q�u��&,�L`��C�r��?�>h8�>t]�=i.Ҿ�<3��s��6`�X�/��B%�YG��m=��= g>M�;>�[�=�>B�=%��5˽�!<o/ڻi�>,�>�d?�IT>o�=�+��Zw�xII?�7��b4�ν����Ͼ��߼F>ÓB>g����� ?����|�Ţ�"Z<��5�>�?Y �?��a?�^@�i���[U>b\>�>D����6�h��w���0>׀�=Gf�M����%�M�J>Aa�>������Ҿrm߾�*�?:ſ��s��qɾ���Ӊ�B���+��Ĩ��ͽ<�8M=����e���|���!���A=�ξ8|��1�>��΄����?��?��>��=;[��3)��'�F���:��?������5�>� y���Ǿ������e���Q�n�\�dS�>��c�󗐿��w���$��m��`M>�-?��žyE��+G�l�p=I>,>.��<�I��ڋ�連�7U�)�U?��5?F:�m+��Z���>��	?20�>��1>T�����̏>�3?�l,?�A�l���=����ڢ�a,�?U#�?j�.?C�����6�}Ͼ�h=�?afA?�E�>����ؒ�eA��?��V?�H�>�T�̽���9�`��>5e[?�\��/Ǽ=��/>u�=�灾�E׾�8'�"�����=3=�>�-�=;��=���2��=?>̅>� �>�����F�Xf�>R�C^�i�J��`�����76=��?�ʾXչ;�>">f�e>������;����M���O?��?��O?6?#�޾�O�ǽ�l�=К�>�~>�<�=����>��>���PT��X����?���?O��?�IO?�}U�C�׿�t����Ծ�L��S��<���=��>�a����=���=����+�xSY>(��>͉8>S��<AJ>sIr>��T>�Ć�#��{��>���&�W��J�����P.��m��v�����|¥�RO�����;\�=�`�v�%�GQ�����_UE����<~�8?A1�>��z>v2�>���=@E��D�	�n＾� f��F�-����پ�l׾��=�-��P�� �¾#('���'��??��Q=�/�>S�?�(l;��>C?�Y<>��=�A�a�>a��>�e�>Fj=WZ2>�T�>��>>�X�>���>pf���!��^���$˾�ӾD�V?�_*�Ac��8�����B�����=t"�=�|�>��<��䲿4Ʃ���>X�4�E��Q�����O�>�_>��R>��0���[>Rq�뒀����=�?ĳ>�>�f�����=�o�>��� z>!� ?��?�?c?�?�μɑ�>��>O��=�#��D�{>��{>�K �s�'>�V+?��]?
E?�8󼎕��[�C�����C�=0J>ھo>��<fA�W�/����<�r�>�缧�w=KY�=цA�l�?��!��N� >|?�HO?���>�un>�6��/�O���P���Mw;NQ �Tt?�C?��?P?G?'?���?�W��Ѡ��!�Z�>��>�`<��셿�SP=��>f��=k��>
*�>\��>j0���@��(�=��>��6?m�1?�/>6�>y�7>*���ѿ�2i�� ���ƽ���=�\>L]�;��M>��D��V��u/�=��=��P���:���=K��>3�>I��>��>.Oc> ���U#<y�h>��:��F�a�=��n��h9����U@>
$\�c����S[����=��U��ʽY몽M��>e�
?�87>�֙>��u��3����7�>��C?3Q�>F�> �=�4A�w2;���0�����+?�:?�4�>G��->9����[�4PQ>7�=U���"m=��m����=+��>�:?WDq>G��<G7������ŉ�>>��=VE0���?"U?����\؆�NQ*����ɾ�!�=�ޗ�3(����~��"��$��p��������9x�>�M�?Xþ$Ƀ>�Q��Q��m�����9���-Z�;��?iP�>�;Y=���=GT��G���!>�_��$2>�OO>	H�>�+?�?�B?�?�>�8T�<^�>�v?>���>�Eh>+�+?M��>���>�:�=���>�%>M������ᑾ��<q��=}@�=h#0>��>�5�M<��n��r�:�!0���ν�MG��1����<0>b�<��4>b�?s�9?�6&>|r��v�{��"��^�iM�j����l�>+Ie>2-����S<���>@;?fy?	��uؓ������޾��^� /?rck?Z�>����S�>A�����,>������7>� ��p��K��[�	�=�<^�>`> � �Dtj>О}?��B?�!?����/�85w�ď+��^���D�>�/�>Y��=��;�63� v�X�]��41��"`���@�}�A=�f�= �>�@>9��=Q�>n̙<���d�Žo˅<RS��	��>}Y�>�0?I�X>qM�=����,���4D?�葾��0�����Ⱦ�h��W�>�>���>-?��1�w�h��W�7��n�>���?���?�_?l�0���~G8>XFG>a�E>��=�S��[7�}�<##�>��=�eu�"b���[.��>)>��׽�g��e1�}Ld��ԯ�n;��8�����!��Xݾ�Ͼ��ǽ�{r�۲߾����5�=�@��U&��3��c����ݾP۾S��?B��?∪>���*|�܈B��D4��L<w���6�&�Ծ�0m����wѽ�t�r���]��c����_�<��>έY�h?��,�|�E�(�ӎ��6�?>5/?�Jƾ+ാU��d�g=h{%>0��<[@��������~�
�T`W?��9?�E�5.���:�ݶ>��?�|�>��%>t&���P�.�>�54?V�-?I��m���.��8ג��f�?��?��-?��bI2�|�;(S�<�&?�j1?�D�>(;��5����+p��v�>�%9?�X�>*E���퇿���f_
?�0V?6�"">8 �>�>�9���b�
>�Y3� >X����=GѼ;	+�����$�_��[�=�C�>�u�>H�9�+�����>L�꾻O���H���L��Ǌ�<!;?
��9>�i>:�>�(�*�������<���L?�r�?#�S?�d8?/��-������9�=��>޲�>�6�=����l�>���>0x辅kr�����?�E�?ΰ�?�Z?Im�l ܿ�H���־SR��BH�=�@�=|�P>�'>z=��*>��c=H��|��=G#*>+=A>.<u>��)>��4>;�4>ń�C������&��'*��������������S����฾؍���'*�\/���O̼�n�b�r�����\��t*_�֗B?k��>b>��\>X|>�|>E��M��\����5���������=�׾�퉽���sz�{{��:���n;�C�W?�u>ݰ�>��?1��^�=��9?�ѝ�D7V>ݫ���3>0��>��>��>l�$>�ee>�S�>�I�>�A�>얋��n����t��奾���%.~?cg����������=��t0>E�?wG�=v�W���������#�>9��m��4�����a5>^�?��>Z-���V�=��7�-�&=�X����>.>�rd>w��h15>05\�[P�>G����}>��?e�?�Ս?�I�?;6=��>��?6��=�� ��?��T'�=�k=C��>T�u?�HK?��?@`f�=˧�3䲾f��ֽ.��<�Q�=<�¼L�s=����=rWT���r�?��!mZ��=!>�1��� �3��>�F?�k>d��>��h��fL��0X�Ϝn�`T�>°$��<1>.�8?b�c?
ʶ>L�.>M�ݽl�������	�z�?�ߒ>�]E�a���;����
�>�n/=�@?N]>�6>\*a�Z�'�>t�<��?B�?돘>�f�>��T>�	�l�Կj�f����=2@>Y�>�%>܅
�8���q�>��Z>�=ɾc
���n���?�B2?"�5=�0�<���>�s�>��4>�r�=^�=�25�[��i�c�>c�=�Ž�
��Q7�^><z;�;�(�=o���{�%����jͱ�z]��z?�?i���X�=Σz�~))�%���:��> j$?� �>m�>�u3>��!�z�)��p�KG��	?|�e?�Y�>%cq�+��#�z��X~>�m�>�h�ʓK>sk��|�»َ�#W�>�?��s>��>s��,�״x���#��>G���S�`�L��?�?L?����Q�U�.�_�!�5���?�4q>B�Ҿ_ؗ�Q����i^������+���׾�'Ҽ�:?���?�l�,>��*��O5��hE�;A��>��?���>0�>���<�e,���Z5����,�=F8>LZ�=9C�>��;?&z8?�A? �	?+�?�z���?<���i ?jN>�; ?�?�l�>�
�>�ׄ>�&�>�R>�I{�f]�����NA/=߸>iF>qSa>V#�X_	=�H>�=h� .��ܓ��j����_>��7>��=��p>�XM>v�?-?4�Z�BA�榨��c����Խ>5�=-:��.v�"�����>���=�??z?'ip>�;�>%`:�ތ���5���Q��D*?ܢC?e��>��s�d>@Mx��` ��=�+!=_���M^�(���Ѫ�B���JL�>��z>�>��j>,�z?�U@?��"?_n�J(��Jz�xH0�	������Ҽ>��>�>&���nE�T�t�"�[�3\3�[LO��T4�0�=��=\ɥ=�Z>�l�=��>hP�<�qϽ�l�����pl=��>Y,�>�?��R>8��=���4(�u�I?�頾���៾��Ͼ�$���>>�;>�M��;?����+}�Q���1�<�Ϟ�>=E�?��?`d?��A�3��q&[>L�U>�\>�9B<DoA�������`�6>@r�=��x�R\����;i][>�Bw>��ǽ��˾���J��.���F�`Y{�c¾ˍ���jf�iy���j��ʰ�.©�)����������@վx�Ⱦ����"��~���_վ�ߣ?]��?ɒO>A����	����ܜ;������/�{�E�s7���!���vϽ׺`�<_žQD���8��^5�o6�r��>��X�p7��#�|���(����G�>>�/?2Iƾ)δ�����h=ň%>�a�<M�`���ױ��,��W?1:?�쾏G�����>��?#�>�+&>������@�><4?6�-?�������x˒�"E�?���?ޝG?�{���;�ܖ���(����>��>�]�>���A�������>��F?.��>~�޾��w�b*�R?�_J?��V��r?>7��>�c�>�� ��tx� �)=���pL��M>,��=�x`����D
�O��<���>�a>��#���b��>j[�s�N���H�����	���<�|?r�Ŗ>#i>�)>�(�~���ȉ�Ձ���L?���?��S?%e8?c=���������l�=�>B��>fʯ=�@���>:��>�%�gr������?y<�?���?mXZ?<�m��~ӿ�`��"m־�}���=Iy4=��{>9r��>�J��AjĽL.��:N>r<�=P��=��b>[}!>�l>(Ņ�g*!��D���'z�9��*���$5���&��c̾]�8�����©��"�� u���½ V�����ܦ�)����a]��j�>8�>�\�=��=���=Rj�����^��댾K,��<�-	ؾ�ཾ,��g{��f1���(�!( �h�_+?���=�/�>ǩ�>��=؋�>�w�>g�߻C;�������Vh>���=�u�>���>���=�+>M��;^�>mњ>����Bg��ǩv��J��Nþֻc?�W����־|��Aӽ垏=��a>r5?�,�>SZb��}���L��w��>����C��k�D����c�>�=M>�<x>�J;�~>|Ҵ��n�� >�u>O�Z>=Rc>�7��2�(�`>2��>�c�ŗB>[��>c@�?EŤ?��d?����Q�>lJ>Q��>��)=�#����;�D=���>��n?S>o?%��>)���O�����]�&��<��ͽ�#=ϲ>��=���=�����	��1��=�aP>v����Vy�ɼu�w��<��>C>0��>��Q?,��>y�Z>W�G����� �k�S i="��ٷ�>^b�>�2#? �?�3?1�_<���=�胾V�x����>��>��D�
���������> g;T"%?��?�'>HU��������<�{�>���>7t�>ǃ�>�
�>/�=��X�Ͽ�N�8�����"����1>dO/�S���o��k����;�k�ی���ǻ���K>s;>~ʨ=RJ>m��>�o=>(���^���Dڻ�=���<����z/�=M��=�F>J_�=k���A����*g>]�O�Ü���䠽u�?�?F#.�.��S���9��}��>���>���>���>��=r��?K��X9�tI�t�>|�j?�?�`3�z2�=U�>�W�ĺ�p�>��>�n$>��8����'c�����<���>-p?@ܜ>���XU�)�s���S�>*��=BEO��k�?��c?Z����q�\�D�Ͼ��U���!�:�>�����hO�����#4��-���11�^�ȾS��=V��>��? �ɾ)��=�8��ô��ೌ�S��7_�<�c����9?���>��;��;>O� i>� ���:٢=*.z>l�5>0w�>�v#?@?J�P?���>]@�>h�q�1?Z5�>�]�>I=��>^�?��?��>qF�>̬>n:׼������A���ս�����2�=C>5P�>�=��׽Й�<�(>�<>�h��6���<��Z=<s�����;x�<|�?{ ?8>�� ��OT�dM�Ɖ����>��X>�`>4M��*�Bs���)?�!=?θ�>�%���ˀ�.�����޾�4����;?�r~?SK?�5�=fo�=t����lO�1V>���>Z֞�[���xʾ�6���=u��>6#>|� E�>�y?T�O?�o?/�>���,��ge��)>�����{C��ϗ-?�w?�1�>�8=Y#���o��Z��8$��l�'DU���U>n>#����Z�>x��>n��>�"�Y�Lhν3�[f5>��?s��><&?�IV>֌�=�?
��G����I?������Ҟ���̾�	�]m>��7>�M ���?@��S�}��P��[<����>@i�?LF�?��c?ȔC�w�$Z>��U>��>�&}<�9��"�F\��9�/>�Q�=POv�|����$H;�>Z>�"u>��Ľ��Ⱦ�P�kyK�cƯ�טK�U@ξ��Ⱦ�N߾-����$�����Ø$��>ðj��-">󗀾IM�R����8��Qv���;�����b�?�љ?�#�=��F�sH�������!�<�Ŏ�%dh���J��f����LY�����M�����P]��=���7>����ф���r�:(�u{�ͩ^>}9?�&ξHF��y �{Ė=Җ>�PB�����A����0��ta?��4?�̾
�پ#���0�=�q�>���>U>upw��?�d�>3�#?�q ?z�=Q�s��_����ֽ�4�?D��?E�"?Й��9Y-��ɾ�v�=��"?*`W?�?���B��� ��E?��?�o�>b{�Gя���׾�+?&Ą?�%���>�J�>�>��o���ʾ�sԽb%��݌=�lt>{=&!��i���w����!>���>ƾu=�����,�Gɮ>lȾu�y�}�F�X�,�Қ �,��NFP?hk���p?�3�>���>�Ah�Y�����ԼW{?�Ǧ?˰O?�z ?�g��4�
�`>3������=�A>>#�=���}V�>�`G>��ƾ��o��%�%8�>&��?^��?�*A?Kqm��οp�����<߮�H�%>=�='RE>[x#��=�t�=��<D�e;��=֮�>V�>Ƶy>4N>��#>�c1>��'�*�pB��z�����.���h��) ��}r��W��	��r��T�ӾoBo��T��OD�z�%��G��9�G��K��`\?��?��>H��>1b�����) �w<���d��hSC��^����	�Ⱦ�}��`Ƚɪ���8|��r߽�F��U�>}�=�6+>r�?k�W��s�=�@>�n�����=����>0�>&�E>AIR>��=��F>��:=KE�>xa�>+�|�����?�b��֋1<��!?G8n��8ξ��J���VB���>�!?��d>@B�P���ē��(�>�$=����G�t�_�\>�O�> ��>���P��=��=.�������b�=C�>��>sj>��ս�=���9�\��>�?��w�L����=�"9?�φ?ˑm?*嗽Pկ>��t>���>��>��>��>�T?�`,?�4?�K!?.??C%�=������<|����~a�A���[9/��;4=��!�2�y=Ѵ;t:�mx�_=��b=BC�=#==V�)=�=�D?�:?Z��>�(�>�Ƀ���+�� B�eȽ��|;�8�����>1b�>�� ?�.�>��>�9�� Ǚ����N��=�>�ɺ>J�m�Ύ�a*5>0�>0g�>��?S2%?��̽׍���oM��o-=�>��.?�Sq?�ޤ>�K���	�[q��y��=�<��Z>��=ϫ!����5�P���<nk>�W��=�=`i�>ۮ�>��>tLk>���=jL8>�1�>Ja>?��=?T�=д=��Q�<a1���=��=t'�=�S�9��FP>s;;�>�
T���ܽ�Q��49��f�>���>i�뽅dE�sd��C�p��/D?���>�2'?���>���>(�,��܄�r�c�@R����>��b??:?��1�QY�=W����m�%(�>F��>�Q><m/>a4^>/���/l>���>	[?e
�>n$���Q�]Ĉ�ؖ���>�m�<��1[�?�U?��K�k8�L�1������Ϡ<=�F<�{�������RK�������Ǡ�=�=��?���?z����
��������>-����2@�>j�E>��.?�|�>5Ʈ��d���V��ߌ���yD�)U�>'->e�>�1?O�.?�o{?��K?�p?�Z�\��=��ż|�5>�>6q?r�4?��?*=�>�,�=��`�i����G�����0�w�W�����=1~$>�B>
��=�.&�N���\0>�ڌ=��=&���b��1=�W>V�>Ղn>�?��V?�SR�m""��Δ>����x�J>�x��ap>�]o��w(��c����#>�$?	�Q?�
?�.N� yC�����X�ܾ������ ?��q?�ϔ>�Cü��Y>�$뾻�$��"�=���=t�'�����������S8�;��>�c�>�֒>/��>!�x?B?d�?�߃����r�����Eq�>j������>��>"&?��Ѿ��]��x��W���A��xA9>��p�^�����>��(>��5=v�>�u�>\��~M��ͽ��w
�%pr>d�>��2?�	N=�p=_���1¾��9?sҘ��%��v������I���v=�K>Κ��r�)?+l���c�ⷱ�x�`�2N�>�H�?�C�?FMv?��J��L�^h)>I/�>H�R>/o"<9�=�ļ,w��Tw�=/6�&ھ�2��5VX=�Lk>X��>,�͜ݾ�ce��������iqK�V}��0������Lƾ%}��)�<�����s��,�1����G��#��6��5��g���c�	�7���?��?���<���<!�M�p J�C@
�@h>oȒ��Cf�HQ�����)���v�0�#y�����O�5����>׾5��>�XY��=����|���(�����?>NM/?(Bƾp�����%*i=��$>�K�<DC�1���i�����
��gW?<:?_&쾡F�����b>��?x}�>F�&>�ӓ�I뽲\�>/i4?m�-?�(�'��8��V���c�?��?�R<?2K=��M8�	5��+�y�?�?��>>H��o�;�0ܽ�@?(J<?e߸>�>��� ��>k�Y?DlH��]d>���>�n�>9~���D���0�e����a\���>X,»��+�>����CC�S�=BӘ>j�M>��s��D��+�>��ɭ��2��ô,�"Q����=M=?h��=#��>?j�>+�>B���3,��|���B��g�a?�.�?1:?sP8?�;����%���yp��o�>X�?�t�>@3>��-�=��?+�
�}�7��վ{��>��?/��?�}?��1����g���\����Ӿ
�=�3�=p�>�d0��I=�KD=�>-��:bXH=Pv�>롎>p�>qAs>�`�=�k�=����%�ߡ�d~����8����$�TS�_��~]�P���:Bľa�о#V��sV��\y;޸L�t�@��G���(þQ��ň,?*�>���>Eu1>���߳��|�M����<���5� �۾������@}��!��~����B��u��=!�MT?��>��=v~�>V���A%�>4n�>{�żj�=u�=oo�>���gI�>���=J�J>���><��N�|>tܦ=�����(���a7���O�r�X<�A?̬W�I#���I2�پG���(��>6	?\J>��)�6k���}w�X�>��;�I�^�<˽�X���g�>t	�>��=��c�Y�׼��}�������=���>�	>2�Իh���#��;X=��>v�վ�;>�n>�B+?�G�?�#?P�u=���>�s>Xdm>	�>v@�>؄g>j�>�D?�p/?<#?��>x{�=aDV��@�k�.=�da�:�нB��'kϼ�	�<��K=aWM<J�=0��=/�j=�A�=.�=�<��|=�"=�?��6?�p�>��>#������ 2
>n����پ(��>�-?�*-?��?��>7��B���柯������>IQ^>��z��	z�۳�=��N�ә�>�i?�zK?��=�k���>̟$>��?��6?p�7?�z�>��=��7�!����޿�!���4����<)!�=�~n�Qw��"�Y=����K��G8�< u�>�۷>t�e>;8\>ᓰ=�>���> /O>1H[=OZ�=շ�����<7��I�><����l�8�Ͻ9�?!���o�*����b�Q���<�ؓ��z?��?v�0=:;p��L��5�����4?2D<?i:?��A?��̽+��t�h��*3��5w��iY>TPH?��>��2�2��>�87<���I+�>���>/G=\�ɻ���`���^ϼM��>�?�1=�;s�ra^�p�8�=-�>\#�=J˚�Ӧ?hބ?�8+�o~#��/)���L��2�@>.�y�龡ִ����@ξ�zO�������==}�<:9?Bx�?���3�>R8���ӷ�+e*��h����=|wJ>�+=?h�=�Ȥ���a��M?�ɏȾ۸ؽ��=��,>�u�>R��>��>���>͇?k�N?�zI>�߼� S=C���`>i�<?��P?�x?d�?s�>(Gg=y����VC����X����[��>�3>��=�<3>���=�>.B)�0�w���(=���=�֣=� S<�=>H��>�/>�W?&KR?���ͤ^�R��>]cI>�>���*ۋ��B�d�����=�-�>b�8?��=?�l�>�;R�L�O��䒿Zr߾h���?b=5?1H�>9%>�}�w~"�x�˾P��:��><.w�W������ᾬ?J< ��>jC�=�#<=�Z�>�q?P+??��?z�������qq�@�=~Q��ž�Ҹ�>@�=+�T>TV�~�>��L����k�m����]>��/���I��Ġ=�>H�j>aV�=���>��=�h����Ҿr��Դ���W�>`��>���>.ʽu�g�'W���ͬ�n�$?�+���ھA3�����	�N=?z��=��!�r�?ñh�(:p�����mR��^�=F:�?�a�?��?�	��ޅ����='�!?s��>L>l%��I�����q���4�>�%������F�S�>tT�>ͩB�:��������r=�ſ�1��R ��#'ھ&�ܾjNϾ(~���:���齄�������˪�E�;:�B>;�NU�3
~�`���۞?�ߝ?魨=�=m��-w���5���Fkd>⇴=8�R�'������	��9���g:����h$5�g��	དྷ&^>@�$�"ϋ��D{��<��U��V�>t�?V���|Y���A�f]O=�U�=Ƃ+<^������b����(
��`?��4?
����\x8���>���>c��>9�>��� �ٽZ;G>��'?*?lz½���RY��U7_�˰?��?s�@?]��<�wE���.��ۼ�N�>ڍ"?f�>��]龵��/"?}�O?j�?Č�>r�"BB�D��>I.? �d�)��>-V�>�g=�=ˆؽ��h��+��T =/��>6�����c�5�=�������>l�
?Äu>���d�$�<��>�6Ӿ�%?�O-���-������o=�3?��־��>&��>&�=by:��	s��k�����"6?q�?�/K?2?O���� ��u�=�ɽ���>�Z�>�a�eE�=ğ
?�>����(j����<#N?q��?���?�Gz?�]g���̿x���ˮ���䵾�� >a��=��<>q���4�=�[�=X,�� A�sS�=��>�Ns>�
�>�P>�z=>��A>e���g",��I���-��u�F�C9����q���Sm��w@�������xPȾP���s���CJV�W0A����*�u�n�\����N�L?���>�c�>�Š> �S:�Q[��9��]��i���(�� ����ܢ����o�a�e�Q���U���a����B��>���m�=�e?�<��{�=;�I>�Ϭ��f>���7�U">>r7>�F >5�>��^>�=j�.�>q�>eW��e ��o�>c��լ�FxB?�D}��/̾�=<��ɾ�$���>�$?N= >�U������K#�>�8h=&�D�eh���&>[��>ߦ>�l��=>d�=_Ǿ~�:� �<��>K�>�>] ʽ������)��b�>>wҾ��=Ce>�5?��?03?��q<�T�> d>,jv>��=gU�>>V�>q�>�/?�fF?u?��>@@�=Um�o���6$���M[�*�������;��
��<c<��޼���=��=7��<�}=�S>S�=ͺ=�<��?H?j�s>��>�B��,0��+P��'>J$������q�>�>�N?u5 ?�»>V���6޾��ƾGѶ����>B�>t���7)���'�>:a���~�>0<0?�(?�N=�Ó�s�G>G�>�?V0C?�6??ݨ=�fļ���*��yGտ�4��%�q����=y�>Ff־;ճ����<%���|�w> �_>���;�v�>F�Y=��"=��#=O�S=��>��d>3��=�[+>����@g�a�3���5<O��׷�;����� ռ2�;����܊<�]�]���f�L��U�=l??1%K��j^�x��(b!��T1�~�?t:c?F?��??\=YL�Ķv���%�e���6F>/}?�i?S����.=�w>[�ݼ� +<��?���>aք��tu���t���G=���>��R?*�>����k�����f�$�B�:�>-�=�᫽�/�?�W?S�K+��2����:"��fV�W۽P뾴m�� ��{#���ƾt�����V�=&p ?��?_�ݾǉ�=p������J_��&n�C1�=��<B��>�>S
����V�ֳ���\������=X�>��>X�v>�u�>��7?�9�?��U?6DO?�����-�>F�x=���B�>]�?�� ?G�?5�>i�>C�����0�F,	�쳬�y)���>��T!=TN>�|�=��:>�>����m��<������K�q��OJ��sr�=s>�Pc>c>;e?�/d?o{�Y��w�>J[��EO�=u�N�/'߼�
�V{Ǿ��m>���>r@m?�%!?!��>9g0���[�x�����7���8?=Ww?ĵ>�bk=���>!�)�R莾~�>�Aj>'=AC�`|m�礠��D��g�>�Z�>��K>�I�>%�w?("T?T)? A����g�s���������@��b�>�i�=	Q>���-mD�q����
Q��)�2�>�RI�!�m��=tp�=l�>�T0>�/Q<A�)>�H��@姾��M=_�m�>�?�>}��>35,=��3��V�����p-?�������<� ��`��{I�%xC��iO>\%�Z��>xl�����������il�J-�>>ٰ?���?�r�?a����޳>ʉ>��>��:>��c��y����4(>����jL������	��p<wi�>��=!?���_^��,J=M����@@��Mw�����j`Ӿh�ھ|�a��0���3���w�*В��
X�h�z���߽�� �归M��E��Yg���@�?�ա?����Ѭ�,�^�ִ:���!����>�g6�3A�n\νRzn��|��V��������k�>��� \�$�>Ps��5��~�l��?������=��@?�ޥ������������<���F$��b5�����R��Z��;N�w?#�J?S࿾������#>D �>NA�>�|�>B����X	�H�>B�-?�L!?F���#����t��!+T���?>�?�-:?�3�A�Q�L��߀��+y>-�>4/?2ι��F�3��=7.?�;?c"c>��J�OE����,���>@�i?�Pӽ��=���>$�w>�4���k���>�����м��>��<t�Zn�(콿[�=�,�>���>�s`��Ⱦ��t>�����lV��gǾ������"��	���>�踾���>����4�ٳs�����;�I�ru=4Hh?���?vI?eVW?''边I��6��=	���[�j>a
?��>���?%�>Q�^;��|���i����>�d�?��?�Ԃ?$"D��jԿ�$��!�M�ξ�π>j�>�Q>+5��X>�,n�����K�=e`<>�/�>�2�>���>IV>!�>���=z<���'��J��Z���q�������#�I������M���2������e;�����<>`F=������"�'`@�ʧ�Ų�=��C?i ?Z��>��?�׋>���Ϙ�>���n���d;?�½O�������p����Ϫ~����Oh�N����E����>׸O������f?�H���V>5]�>�B�<�j�>��c>O[>!�=�5�>�c�=��5>��>X�Ř�>�22>+�|�x�����]f5�=¼�^8?'�����t+�8Ժ���n�2�>D�?�D>\@�6���JR���ʩ>�׋<H�E�2�-�#)=��>���>�d�<�Z�=��ۼ�v����V�oA>�ה>��=�4{=��H�BKY�[Y����>�����(>��>��%?��?�=?�z��#�>��N>���>��#=��;>0�f>&%�>��>�X'?��$?A�>3�=��i��}
���=)3��sϼ�q��u½��k<+y�<�Uؼ�^=��'=�/�=�>��>���=g�>�T=
?��6?J�>xG�>֠R�2���7��ز<Zx����>�;'?�y�>���>s��>[~�>	R��A��u�C�����>�Ԩ>j���I*��h�">��=�<��?�3?��ʽ�����T>��=�k�>g=?�a?n� =�&Q=���t6���ӿl	��|�n���>���=y�I���F�	�>�P��PU־�9>2�>�V�>'q?h8�>���>�|"=!�>���>iY>�>��=�J��"p�<��f�
�ʽ	��=�<1G��}mx<d|3=����0����ԏt����=%�? ?/0>?�<VZ��/�X8�L?�A?�6?ɤ3?t��=��ʾ߽:��L_�����Kl>�}'?�� ?��ӽҹ	>��>h�Ͻw_�>�A�>���=��8>9j�Ә������@�>��:?L��=E7s�"*h�{I��ܔ$���>�A�=b���0�?�T?{P!�Nw�<���|b�F_���@�=���.�����i��:ʾ�'�~�ɾ���d-����$��M�>�&�?���)��� �����z�I�����>�J>kf"?W�[>;�xA(���<��{ؾ�fӽ G�<��$>	�V>�o�>4�>aX�>�S?
?UGr?�ӆ����>��=o^?�|?d�?�d?�W�>:��=��U>�.=�/L��b��c��hS����B2Ի��=reG>��=m��;�FN=S&L=y<WR�1]�s%�=?�C>΁b>� �=Ƙ>H_?�#L?��
�,��k��>�L�;��3>5��,�(>m޾�_���Q�=�E�>�=?U�W?83�>���'�R�oJ������B��r?�5W?�b	?ck�=fm>
4�������%=w�=7�4�W���∾����U�=�c�>�s>�0�>�`�>N�?_Y?�b?�¾���}�"�*�EF���>[ش>6Y>���>Ⱦ��{�����Nj��*����>��"�������=kp1>�#u>�g+>��E>__Q�W2���~��w��.��sz>���>y�>���<�r<}ܾك����4?���$ؾ]@���V=�	qE�>_Z�>`*�>x-?	�=j!�cĿ�:��df"�@,�?'��?&�?˝%�֥��5�=k'?���>O{��L��ζ�y����=�*>ԋ��qCܾDV>�x�>�1�=)�;0�ľ�>$���<���rG�'��=���Q�����tH�Y�W��恾��f���龬���ʠp�>�m���.������6�� �������?��?�� >;H�:}�D��:7�ɷ�Z��1,��k�N����z*ɾ>8�����@��u����o̾<���V�ƾ�̛>c�X�W��?�|�w�(�[I����@>�.?�xƾS﴾���f=B�%>�ٴ<���R��������Z�<-W?��9?@�P����tὼ�>|?�d�>��&>_���T뽎��>�F4?R-?h�����3���Do�?���?�W??�D��N>��.�w1���?�?���>��S�Ⱦ��ֽ8
?d�7?�ռ>����)�������>U�V?�^M��R>���>b�>�,ͽ����g]U�r���藼]�5>,9�"2���c�ۛ)�n �=7|�>p��>1VF������>���V�Z���>������<�銦��j5?}X���>ޭ�>�C�>d�B�����ꂘ��l���9'?���?�1V?�?���w���hS�=mY�z�a>��>��"���.<��>H�?ʀ�&�V�5G㾝�?]T�?{��?�,�?�Ml���Ϳ񆚿q���ԸӾog�=^�<���k	���>X0=͐��6	�=��@>�o�>j��>�K>b!>4;�=�*�=����ZR,��ĝ�!Ď�+�l��DE.��@q�r�쾄������n���L��*��vjĽ�?��~B���Å���b�]���J?�L�>I��>��>��6�����0Y���پ9>M�����Ǳ�� �����NV!>v��bH���>��{ �y��>��˽$��=��?�.���">*w�>��F���u>=qV>��>h�w>+�="<x�>���ڒ�>�r>�����M�3�L��C><�A?R�j��گ�}�9�淪���j��Ů>2�?�6>U�.�
��N�y���>i���R��b߽�j�<a��>�޸>�zM=��4=�H�LV����=)�=��>�51>�J3=�ck�Kw�;aɼJ�>cp�x��>%	�>��?�?��?�	�=�_�>�n>��h>�,{���0>O;>R:�>�?�H?�=?U�> �=�6���<Wr�=G��������<����XP=|~����G�q=D�%�S��=m�0>��=�g���=��=!?2�C?��>�3�>�|���-�ƨ.��b�=�䅼Z������>S;�>� ?���>"8�>�AϽ�i���T���Kþ�@�>ق[>\Q�������di>��=(�o>�%?��?��K����|�>�FD>��?uM5?� ?`�9>�aƻ��o�p���W�ÿ��8���(�-IT=�`Q>�@=P���K��0��=�d�=+�;���>8ը>1����]y�'(��gT>Ŀ�>ς>�,\<��K=��=�@�<�:�=�F�<��Q���==j�=e�D�uu��y*��sн�6����f=�H=�>�&?�55?��>�=y}��~�"���|:?�/�?ݑU?�4Y?��c�RK�����8��	A���>Z@`?0��>������>�=/X��2<�>��>+���\�=��R��G�E��<��>��.?�!>�Pg��O� �?��b�t��>�6,=g�˽�\�?��Z?� �|�m�6!��v5��j �{B�Ho������:˭���(�do/�+�|��;Y�<��=���>W(�?��Q�=�@Ⱦ����klY�M����>�k�=�ο>U�Y>�b;������͍��5����!;;\d�>���=�>/|!?A�?+�\?�,?�+?����4�?���=��>�Ϳ>�i??��>_�]>Kuz>�O=:_�=��Eg���hF<�S��ʝ={[#>�� >�̟<�M�<���=�<[�&���$��o�<�44<��<��q=#��=�~>H�?�b?doH�x4߽��2?��;����>�ٌ�"�"=g���#���=$>q+?��P?�9Z?��>"��A�e�a^��P#���Xm�2U+?�CP?�>]
<1B>�&�I������=��x>C|}��{g���ݾح��Զ�s܅>֘�=��=Yї>G�t?ۍ]?R+?&',��{�%a��7ɾ��]������
�> �F>ɉ>��оo�3��$}��H�D��Ͳ�=�6-��� <`�N=��r=ld>���=��=/Ψ=��r��o��|/��G#=�H�>���>�2�>��=�4�:��¾9����g0?����f�<���>3�Hx>��?}�۽!��*��>����}����:�$��P�>���?L��?��|?�ˁ��4�l>��>+0`>K��������	?�����|�`>k!;><���̂쾊��=X��=hq">�N������K���3��E��pN4���R��vþ8���5��?���<��f���>�������d�de��l���tc�%(_���^������$L�^E�?��?3�=w�=(��q�6���=�B>]�5�����i`����e,��50���v����"���~�Ѿ8Vp>𜽢'��AaV�"�㻾D��=GV*?k?���B���v'�c?	>6�@=:����j;�Yo������F�Q����?�8a?�Ѿ�W��v��A �q(?T`�>�<�>�þ��$����<��T?f�>+�>)�g�������9λ?��?e�A?q@n�=<J�^�)�s�.�>���>��>YT�����t����.?@??ˠ�>�Gž�ʂ�O!+�Վ�>��9?���_v>��>6D>�B<Q/�Ã�o���[=V�;>�J�RN�|�a��[���,>���>�t�>%ޞ�&�����>��@5N�1�E���l��[� =�/?�8���>bAX>)>E(�{9��������htO?���?��V?�5?*9���	��½�,�=^��>��>@��=�l�eۛ>���>�<��lo���??
��?���?�5Y?H�j�t\ӿO ��#Ľ�y�;!�R>��8>�i\>>vj�4�">�w=��:�ڑx�� �=�z�>���>]�{>���>���>j�~>{��@�&��w��9Ϛ�.�F�]��ԇ���e�����n�����'ų�n5־K��������D�)�� ���ǔ�8�z��x�R��>�Q�>B�\>�>�=X�>�m��A�K����J�����n�bD#�B��`�'�M�ǽo�������>Y�;�*�5#c?��;>���=�4�>�u]��G�>��>���>���>�F>�m�>�>4iW>��>�x�>�~�>&��>�i>��N>'����Z��J;\�]e�z⋾��R?iY=�,U��||��FD�{�,�_�>HH?�u����j���|�gRW�k��>̐�<����̿<�?�<�y�>��>���='-l��q�Ӏ��akK����R�>���>��{��l9�˳�xk�6�>	E�$D�>���>�J?rR=?�D1?�G�=w��>ͦ�>	إ>o�=�K	>ȅ=y!>��?-9?D�2?g	?��)=�eM���0=�L=�(���/��N߽}�a��9>��>ؑ�p�۽�uN>o��(n};0+>rüF޼�U%>;��>��1?M�>�|�>�=�<k� ��wS� }��A��=3�.���>m{?��*?yG?�m�>�]>���Db߾e��\�>�P�>�T��~�6�(�:�>6�=�i?��?4����$��ߵ=׆e>vm�>f�>D�?W>>��-׌��z���߿6
(���4� �I�zj\=��[=�L!����=?U<ˡ���S�4&1<%�R>�*F>x�> B�>�>�g>���>���>1g�=��r=p�f�7����߼Z�%��[�'VI� ��= �=������<�򧽹K�yo0��������<ap?)�>io=�m�>��R���E	T>3�?��?g�?��m>$:'<�޾'�|�뷇�񭛽G�*?ᐋ?VT?�%J�����������
��?p�b>`Q�=S`|>�
��S���`���>�>��>��H�q��q�6aD�{7�>��H<~�6���?"�a?�������� ���A��F���&�=b�ɽ^[G�A���N!�X9�((׾�6��[���
��=�~�>�"�?����� ���4�����Ծ�y�<�!r<���>�<�>'�k��pa�}��ŋ˾B��9�>�0@>|�A>G�?1 	?-_*>��^?w�N?�g=M���>�s��?�#?݁=?/�;?��>o >�ث=$\x�e6���#v��n3�A����4�x�=w�=�ĺ=�~�=b�=�&�<���=���=g%��Gc<{�S<�>��4>���!��<k�#?�� ?VxʼK�>9��=r9����?�MS=>J|3>
}3�ջ����>9Wm>w��>�e ?��>���=^Ӿ)�׾`T��R�l��)$?O?p��>O��h�>ޅ��S�o��T�=�)f>R4�=�v�����l�����H>��?<�Y>�N\>	z?��??V?���3��r�um7��>G��jU�}�>/޼>�6>�᩾Uv$��e���Y��Q/��۞��m$��~�=>�=�Ƣ<i$?>��_>BV�=�Iȼ]L��[<��=V{��9�>Mk�>qa�>��B>eb:=cϯ���b�I?Z͝�G�hړ�=�Ҿ�9&��,>2�3>HJؽ��?�� �.]x�ԣ�H�?��W�>~��?���?kJe?`�(���M2O>�bO>͟>��C���D�V$���H��f�5>���=�~�⪛�iy�<F^E>֪W>�ऽ=z��11ݾ�lּN<��F�[��Fw�����
�A����i���A�
�V�~�������轐��(�Scs���=����B��L!��̙?���?�T����L����8�w�����=(J��	[n���˾v�н+ǫ�:�����P�w�{���U��}#�	�>(�(�ᥙ��x�X5�S'S��o>I�5?��¾�[���y'�}��[�N=:&�9���$��  ��Ϩ��lA?�-?���t<��3&���>�� ?���>M��=�;־\(2��1�>;A?�1?��'��-����y��_;=2��?Q��?�8?6A��P�0/��������>��?>��>�'����\���>J?6L>�%��3���
�9Y�>;/B?Y
`�u/>�_�>JP�>�R��&IR�����궾b����}�=��<W�=#_�fr���3���һ>DӞ>�"t��ھ���>:?�7�N���H�������'/�<p�?���4>�i>:>��(����ω�}$���L?��?��S?�k8?�\��T��h������=]��>5Ѭ>���=f����>?��>a�Pvr�B�&�?�I�?~��?lYZ?��m� cֿ["���ꢾ������E>l�>�>w�a�\�����;��<�û��J=���>M�->�k>IN5>A<i>>Ua>����Ǻ$�qh���h��.�B����P���R��������آ��,���>�����<�D����	�����M,��������=9h�>���>��P>��=W8�=���=���G�D	��Y8#��>;�Y�]P
��.]��8�d���Q$��ZQ��	�m�U?z�v=un�=�>E�>� >�>��>�)?vY�>w��>�?l��>��>|�	>�O ?���>��>g��>�����~����)Ǩ<=
|�fy?���>�0ƾ4�\��?%�B�/��b���n>�=o쎾m�����r�G>�>lav�q�1���=��=��)>�x@>�Q>�N��x�������<�>û�Ҽ�A�쭽>wz�S����bF�6%.>f ��i>ZS��'�n?  �?ghS?�b�>.\�>8�>���>���>s�d>���>@�>,9w?��?�X?#�Z?�绒���~_"���D�+��J�>�����i�=��=�9�V��V�#���v����=�J=�+���<�>A��>AAK?��>��?�N���#]��G�*�ܾC񷽨G�>��?k?.�P?9?��>���� > q[����н>��N>0r1�h^�h7a=_��=0���}�	?d$?�s��ZAl����>v%<rU�>i/?:(�>�Q5>,�s��!+=�F��~⿿S	���C���;1�ʻ
"�=�὎��<�uü�Q��{����Ǽ(�>s�>g�f>(��<=r�>���>|g�>�NW>���;c_=�/Ҽ��\���;�d^>t�=h�0=ὃ�X�\��<��I�'N��K��=!�>���=�� >�C?�?{/��7v���h�v���ȧ�c�>";�>y5�>hW�>:ٴ=�����S�W�@��9K�8��>˘e?��>O 9��_�=dC�ڏ�;i�>���>�/>.�������i��)��<S�>��?k4�>����Y�iMn�	��v�>g�h=E���Ԑ?�`?h���M�'���w�H�p���W��$�	>y+�+x���
���g��T�D4�#Z��&y�=ŋ�>�¯?��v
>�2��隿}���M�4|���r�=�<��
>��Ҿ���V,��F9��e��)��/�>>>$�>�%?�D!?�(5?ˏ�>υ?	o����>	��>��?"��>��?<�.?g�>�>y-�>��j>����$h>��ɒ���S=.�[�]�x>.la>|>�gI=��=`e�=d����=�B�<w����=N�N>"N��w�O>T�>�?�V'?g�����>1�ּs�o�t�=A��=
E��F��T���>N�>�'i>��?�|R= �4>�Y��5���;���uQ¼v?3Q?�^W>m�l����>��z��ɾ�d�-�=ɷ}��͚�����O���潭��>���>%Z!���v>��i?x(?�?%���d ��x����"���F�þ��ȼ���=���<b,���1�+o�0����aS��ʮ<Qi=��~K==�<>p�>(�:>�S>s �>ZO¹֚`��l�>�{=���:{?��>`M?'y�>R>\~C�9cȾ�J?1��B��3���־���L�>`~>>O���\ ?���!�}�"��|�>����>��?��?�R^?��L��Y��V>k�^>F� >���<82F�c@�����>/�=� w�eE��!�u;�cM>fhi>�
̽��̾�澴yc�����v9�I��q�#��	¾
��������={�����(���� ��u����J��!�<]ż;�2}���A���*����?���?**~��L"�t3n��þ�`���,�U։��(���;�����e���7O���ʾ���v���}:�]�N�$�>�1Y��8����|��(�������>>�//?�]ƾ7紾5��"d=ܧ$>:��<��ﾠ������������V?ȯ9?6l��8���L཯`>��?�b�>�&&>�9���N�/}�>84?"�-?D�������b��6\�?`��?GA?��5��H�kY�A.���?���>N�>����� ׾�e���?Z�$?��>��m`��N�����>	�F?�HS�d�I>P��>�ʫ>�Ņ�����3{��p���F���%B>�ʼ���fb��m[��3=�]�>��N>�cx�W���c��>�&�c�N�d�H�P��l8���<p?����=>�Mi>i>|�(����_؉�#J���L?ߍ�?!�S?)]8?�X����1���b�=p�>��>��=���e͞>.��>k)辢lr������?y:�? ��?�LZ?��m������k?¾E��=�
��>�J�>V�1=pˌ>Rm:<�:�wQ�=|,h>S>�>�o�>	�>�6�>�I>)��>xt���S"�A�����R�H�Bu�=���2I��d���yc��,پ	�*�jپ[�*�b���<ā�ooV����� �JI3=e%?���>y�>q.!=�c>�5��`�+���z���h�kDȾg�-����x���,��:�����[����������@1?�P�9>��?�>:�f>Ch�>��%=���<��>��#>�.?�$�>猳>�>N@�=TBh=��>�+T>׸���v�������žM���'�A?�o�羍P���:�����+�x�JR�>���=h.4��?��G���|G�>$���2J��T5X=�r?=�+>!US>�������K���q󌾀a,��$�����k����꾴����T~���>����-�>i��>g�F?�f?D�Q?�~c>��>!$�>B>����>�b�>�=�>��$?ĕ6?4+?�Q�>�+=�󖾁1��YG<�D�r���B�\��>����g�E��a����-�������Լ��%>'![��'�=�+>���>��8?G��>�Q�>L�����sG�WH�aI>C⼭�>J��>�+?���>j��>�k%>"j޽�����ξq��>�+>�S��r]������O>ns�>%dO?~*?�>���	}��W�=ȭ�=�W�>�T?01*?lu�>Pf> ����鿉U'���Z�ޮ��D�����=�=弡B>�'>=B&�G>�=ۨ=��G>��> ��><�>E�>���>��>�5>s��<�q�=%x�:�=�VѼ(M�W{�����=�N�;���<�ý�⇽fY�O���:���iO=��<'?�M?{W	�����N�� ��EǾn2�>��>\��>�?��="����xV�.�P���N�z��>R%a?Ot?������= *����+�au�>�8�>SS>Ӥ���K��&x�Ĥz�*�>{�?�>���D\Q��RN�F,��`�>f �=�]|��?Y?��k���վT��J�Y��v�>=<i=�q��������Ծ	�=�2�ھ���
ɜ�b��=u��>��?I�ž�h��?�g7�����t���w�[�6=Ɇ�>���>��p�q�׾� W���O�!=�,G>Ȗ?�Z�=ܒ�>�y*?nP(?<�'?Y�??i.?BA�Ƥ�>�0�=k��>�w>��>
�#?~�?%=R>�Խ>��=6�	�ei��<m�d�=�Q���= �=��:>C9�=�>V4T>��K=�����>�I>�x2=r�P>}�]>,�4>Z�?>})?�;"?ᄽpE�=�Z ���K�*>6�2>[1�=O�������="P�=�X�>2"?���>m1>ꥑ��i�Ҿ���<��?�B?��h>�R�<H�>Еb�*�����뽂k?>�w��GԾ�*\�-��R�u>"Ԅ>���<�n>��n?W9?�y�>�/H>b����~�=��pp��ǜ>>4�>��C>���>�
/�(&A� H����C���Ǿ	A�>�Lս��=<$�<���]>V�>���>Xz���LH=�,��!��ӥ�.Y�>o?�U(?ʑ>k�< �,���3�I?���_k����о����>��<>���k�?�����}�P���@=����>A��?��?�2d?D���V�\>�8V>Q�>�.<�>��;�3m����3>�4�=�y�\����;�]>Ky>��ɽ]�ʾPE�-�H������0��c�����ܗӾ#���$��%s=l7½*k��RFX��'���L���	�Q����u>�z���G�<S�'��a�?vġ?�v*�T��=��[�X'A�7�7�-�=��D��'����Q����M���D�þ����}̾�4��R>���P��U�>(a.��r���c��i0���"� >�=�w?*�׾nP��ns�,߼��=T��*�CQ��Zb��[^�oR/?i�?V��p�n��
=�@V>�Q�>%��>��<���"P=	d�>��)?�p$?S��&	���承�;�=���?��?;S@?�r��<�.Z�ʊ��� ?m{?�I�>�N��\Ⱦ��ɽ`�?�N2?�Ȩ>e$�ު���v���>w�O?&G��)Z>=��>�b�>������M+=��{�-I���K�=*�b��/����2�	�>/��>j_�>i��¾���>��龈MN��H�A��M��j�<t�?�n�z>ig>l�>"�(�)댿q���=��QM?�{�?ҍS?G�7?�j����S���s�=攦> :�>��=�<��j�>�>��jr����<?f�?	��?Z?�l�=Gӿ��������	��=%�=��>>��޽�ɭ=��K=�Ș��Y=�r�>���>o>E;x>x�T>˛<>��.>q�����#��ʤ�3ْ��[B�� ���wg��{	��y�����ȴ���F�������=Г�t�G�[���T>�>6񽑖�<*�
?�g�><�=�5�TD$>tQ�E�������4=��n���钾cO���{�p5޽ʇپT�ž��ɾ �b�B?��E>sE7>�L�>��Q>弉=,d?��?>���>��=$E�>�� ?�T>�>Nߘ>�ӗ>�d�>��>��>����ޯ|�R����-�D���+?���>��澖MG�ǐ)��z��
f�O�?�>0U"�7�T���F���>�����I����)�Ù��h�>���>X�	>���F=Vg��땾Bl���	>�\��nf�N�^���� �}.=t�G���>ٌ�=!�$?7=�?���?�?���>���>Mc�>_�>�,>2�z>�>�B?�~?A)i?V�g?�����.ʾ��Ri���X��S�=%�W���	>1�F� �Ѽ�ʘ��Y=�����Ժ�1>� �<���;��=���=��>��B?m�>��>�)�=K|5��.A��v�X�T=�_�H8?~�?�U?��?4�>فH>������澴w�>�z>!�T��ɉ�ω��+�>F�=��*?ɔ?���<�z���=��=�7[>�>��> �>��&>�����2mӿ&�#���!�	������_�;��<�*�M��A�8ta-��e�����<)�\>+�>p>�(E>ͣ>=3>6D�>=GG>,ʄ=3�=�^�;X�;F�ATM=��5H<�4Q�������ȼB̗�Yl����I��w>�s�zvۼq "?:�?M�����?���ξy����hK>,��>yl"?�\�>=��=���j(K��4���۾m��> uk?1y�>;�#�i���;�_�=�/>�<p>?2>���=�&�ر�R#!�F�>���>!_E>$�n��]�I�<����:�>6�p�	c
���?�
w?�N���g����G����A0=_�M�Z������8�ؾ�H���4d��Ad��C�9�8�>�4�?�xؾx!D<�c�"x���X}������=�-�;�̎>d0�=/�����Ӿ���ʥ��~��� �l\�>��?<�Ă>��$?pT9?�=9?kH�>$�,?W����>�/>+��>���>��?7�?@��>��r>?��>�>|���\�l�:��<%�e<x��˾<�6>��I��s
�A�S>o" =�'=�Z:�Tü�>S��=�1Q=\a5>;@>B�?A�!?7V����T<�h���UZ�)�=�%�=nH��r����� `O>f?a>N2	?���>c��<�R���& ����Q+���?~�?*#�>�e&�l�V>���w�Ծ���=~Oi>�T�H&��XM������&V�Fp�>��>\�=�f�=Ngm?�=/?$�?ъ>,��jl���n�6�M���<��+>h��>'�\>K.\�XwL��h�6|n���<�΃s=�t�׵�=�/>|�ڽ�P >_�y>qS�=i�=ů�<-=�Z��=];�=>d+?A5�>��>��?gOS>�+��Gs��J?�M�����]顾_zѾ�w
��=>��?>#� ���?�g�./~�~���>�!.�>?��?���?��b?�E������X>6DZ>^�>Gc�<�';�$��>��9*>�=��u�lՐ�4Z�;�XT>��q>Biɽ?ɾ<��A~P��ſ�MU�]���޿�$����A¾ �v��4����J�u�#�����$�%��Qu�0!)��e�<�"�w�;�����?�?' �?��ƽ�.=�$3��6��j8��Sڽ�G��us��O\��@��}������̻����@�~��Ѫ����>+7�����}}�����w�9,>	�#?'�¾����4��P=9� >��<��篋��u��E�ܽ�R?S�4?��ﾧ4��Q�ɽI�>�?�q�>�<>�p��u�Ľn��>x�.?�f?Y�H��ߎ��ڐ�����ʻ?���?�iQ?��̽p�6��������>V��>��>`��Y�������?:W�>��^=�A��O����p�>-&?�Mw�۬�=�+?���>A�c��Ӿ��=�2�������<0v��Ľ'�c�:�C�7:=��V�>k�x>쌶�!�Ǿ���>�@���N�ڪH�������J�<��?���4>qi>�?>��(����`ω��)��L?T��?Y�S?$l8?]����(������=��>uѬ>���=���v�>��>�d辶wr�����?3J�?)��?�[Z?1�m���ӿ�e���Zپ?����m>�_�>0��>�,_<��7>Fԋ=I6>aT�<F�
>�Ϙ>]�&>T�>�>��>�`z>����U=#�7ࢿ�o��<+�Z)�b�徐�2���;#X1��0�{��V~��~"Ƚ�z���b�(�I��7�����2��2>q3�>3�?�R�<���=���=�=��u�R��]�������_�ƾ�d�܎p��bս��������hh`��)&��fo?���;���>�k>�����>"S> ��>B�>�v�>�r>֋�><��>�=�=�X�>Ut>���>v~�>�4�><	��~s��8��!u�:��ݍ>��>h�=�������>!��j�kl�>�^�<q+�����ࠃ�E*�>�l�<�ƾ=;L>8u��X|�>�?}=2=�l���xھt���<�s�x�<�{>��_�����݆��ۻ��ۘ=)h�>�L�L>>��W�_d?hnz?�5�?�?�!t>4�?w!�>�`z=
�>���>0�?��D?��Y?Ifu?.zf?��<c)L�h��"5���3j�w��=Eħ<uX�<� ���uC���=���޽�B4��Q���<0>����=�>@>Ct�>3g??�j�>k��>���d�5���:�\w����>�� ��>�>�>�5?�&?Q��>rZ=�o��B�����Cy�>߀>J29�z�L��R���t>/��>JL??�/?K<e=����=L�=�O:>�t�>�"?���>��>C*1�^����4οA�+�~gj����=�>�C�=�)>��>)K>d���J�����=���=�ۈ>e��> {�>���>���>���>�>2��=;�6>�n='+�<�䷽�ټ��]�����!ɖ��Q�؂�ReȽ.{,�3%>��&���(�W���?�N?;z-������j�I���X	�����>�F�>Ґ�>a&�> c�=�F�V�U�z�?�R�F�ю�>o�f?M��>�3�*��= w?���1;���>hՠ>�>��q�G�����*Z<W��>�?Rp�>*c�R[�uo�g
���>_�L>*s^=�=�?S,r?Kb��n��٨2�?��[J���b�-��=�P��4����=.�5U4�L� �X�@�*ھ�]ɽ.N�>�s�??PȾɠJ��<o�����誟�)���̹�&�,����>O��>~5@�e>��t.V��!(�F���Nұ���>4>"Q�>�H?,?oY)?u�>�)?Y8���>L��>ו?�>�?�8?�"�>��c>�;�>�Z>�`�=c�X����Ioμ"Sp��[6>�ΐ>��9>��m>w��;���=n����μ����\k��� >�e�=���=���>�?�>�?N�.?T����#�>Ctp����:��<e��<泛<_����hIG=�c�>�?yG�>�2r>��>��ؾ�;'�Efᾪb<?-?��J?�l�>�<5:e>|���G汾āv=��>!����q����l��ϾC�=ú!>�Ч>���b]�>Âu?Ed?��>+�>p3�V掿S�4�6���j����L�>�V�>P�
>ƍ澰�F��⎿C���#6J�^�̽��c�=�=q�=�SX=��W>&�>�Lݽ�4>K�=6��FJ�� �>�5)?�n?�?>�"�>	NҽAw��=I?�������_O����Ѿ��:�<9>��8>�s���&?*����|�s��i�=����>��?���?�lc?iH����΋_>��N>��>ǹ�;�{<����*���xo4>Ƀ�=�u}���R�<&9\>�uu>8�ѽ�Vɾ��⾡�W��ū�Lp1���3�/��N15�����F���/���<�/Ͻ@�f����ξ�/���G;�Ko=9௾B)��ܼ@���?Ë�?��|=E�_��J�{�^��p9����3Ϸ���<�L��T>���,����'�7����,��u*�Q?���>'�R����;{�%�+��x��pw>>p-?K�þ���j��[]K=X�>�Շ<�B�%��i���K���T?�8?Cc����m�̽��>�?��>�:$>��`����C�>+4?�-?�S�wY���抿}����M�?�l�?F�@?9B�JQ?��@����4�?Q�? 1�>�܌��UҾ�1����?�6?~͵>b����ܹ�> �>J�V?�WM��]>6p�>>�����"��:"���!��D�A>Y���� ��Y�,�yl�=�ȟ>�n�>_����q�>Jq���T�pmV�@e�d|"��/7=�Z�>�7��D?>��0>��=\� ��v��`���}6�,�9?�{�?�PU?�@+?��׾�t��Kt���T�<��t>C�n>��=�$��u*�>Ӈ�>��ݾn |��.��x?Ҥ�?W��?*nO?�Rt�F?�$|���Ҿ�����N>SAP>�Dt>.f�U8�=�ʻ�[0���>=�A1>$�e>��9>��y>%�&>I�s>׺e>�7����&�����튿��2�����%��^��� ��Zξ��$�pV��'h��ԛC�-����$��x���yl���Gz>���>:q>��>�TU>���=͵{�f����̽Ǎ��H/�|7��kE	�������i�a���+=�=
C��7Y���?�^Z<�=��>ۊ�=��<�?\��=&�> $�>��*>�P>�$>��>H)�>����=��)>O=5H���Vr�	zo��F���	��L�Z?��H�uz�-�ɾ��z��6�=��?�R>|0�c��+��ñ?=J�'���KSɽK������>.�>|�	>Ӣཐ�����?/�����T>�9>L�M�����nH�),>��>������>ޱ>�C0?4݆?}Z?f�>$�?���>W�V>��`=���>ܭ�>o�>�?�A?�7?b\�>J��=�b(���$>�>�n���=��=gL,��h�;���;!����ۢ<�,>���=4�=�V>�Ϧ=��<>3�?�L@?��.>��>gyܾQۄ�����l��=p�>����l�X?�A?ʶ1?��>��?^�>�9>d7���b����>χ >S�y�O�����6A~>�>�=q�'?�j:?�I����y� s�>�f�>�R�>�y$?LtL?�b
?�i�=��J����l�' *���(�\���Cv=��>C���!�<�-Z�;����L��$���L>5��>��>
ؔ>�փ>ܓR>�u�>WH>8)u=RŻ	��o�	=��T��)=o�H�
r�<��=�i�ݐJ�̪n=#U�=l����l��@��K�����>>�?돉�c:-��������Y���d�>�g�>��?v>F��*�L�\���W�������O>#�?Mg ?���<�>>fH0=�� >R/?Q��>s��=�27=>�����A�5H>���>B0�>�DL��DD��rZ�����u>og=�f�:�?ก?��Ҿ]��n;���Z�tZ߾V���P���l��h\ؾ�� �SAO��c��w� �����<�>�q�>;�?xV�ݵ)>(y˾\
��X���]�1F��ɱ>���>��>>�I�ʕr����"o���W��>��)>�>	#>��?v�?$�x?9.�>�6?(6=��>�n?��>RM?X�;?a^?��*?N<&?�I/?�q=�)`�Ny���H�O�h�ݽR�=��2>]OM>���=�/=�8&�\ o��Q�q�U=�&��5������=���=��>)/?i�#?�3����P��#�޾�"/�~�|>��>�Cs����=�I?0�>��!?��N?*�3?a�>!Y���7�jž����D5?DAK?_�?���=z:y>@`������>`��=-�W�� ݾ��D�������_%"=���>7�>�>�A�?��u?�7?�%]=�����ˁ���g��I���@��<>����5�S�2�F��ZB���G�N}W��`�9>�v��ƀ	�xB���/>���=������6>,��>8�=�}�����=m��=$t>���=��>��5>?���k¾��'�I?[����j�C���%xо]����>k�<>���?���C�}�f
���J=�,��>���? ��?�Bd?��C�<2���\>�bV>)>x�.<��>��O�������3>��=Byy�������;��\>�Uy>��ɽ:�ʾ�4�٢H�6�ÿf��s�Q��|���Ͼ�w��6����߸L�������`4g���,�O<��޽����㧾l����΢??m�?�>c�~|q=�I��f<�8�
����>�3���ڇ�{��v�������2��m�m�z/i�=���>� ��6Z���C����w�gH�>��:>�RB?GT[��V߾��&�Ɇ�f�=�K��ھ��'���^����I��f?�.K?_��������ž_�
?ҋ?�1"?��?��፾�W>��=�b�>�q?7~�>U�ÿ������փ�?
��?&�E?�l���Bg�x�W�������>�<?�>���v�,r��U�>tK?��s>�lT�n��n�6���V?�Av?hLm�2��>P�+?ԭ�>Q�N� 	��1��ꟾ��>>��>�# �zc�ʛ�����"@=/�?3�>
ߍ��0�Җ�>`��5k���i�q��ZNл����S�>��i�V��=4F=	�+>C,�E���>���_ށ�J"�>�Q�?ᬋ?��?I醾�w�=�����"�B�[;�C�=�'ؽ�G=�#�> k�>���.��,<2�&?-��?���?��3?�f���ۿ�ɣ�� ����ؾ�� >�L�=2�E>�wr���]>�>�=FI��.�ý�h�=z?�>)�r>mb>��=0D>��&>|�����#�b���@O���,Q�~Q1�����U~��W�����s[&�*I׾Ц|��lǽ�t���H��V`��I����d$=��=�=��>nX�>�?�>׍�>{��=U�{��!�A�������鼾�2�V�6�@�-�t���꫾.���ýM����L�QN��Z?��A=�?�=���>m	��Q7>���>��>��>�)�>��m>؀�>[(�>���;�y�=��>:"����x>�.�=���EÀ���;��T�.�;\@E?��T��ߝ��2��ܾ�M���(�>Zg?\S>��(�L����mw�/��>I�)���l�%&Խ�>?�,��>���>��=����6,� �r��(｀��=�S|>�>�e��	���2��t��=P9�>q)�XW�=�K>J:?�΂?,MN?x-|=wJ�>w8�>B>��]��:�>it�>��>�
?L�G?,?7��>�\�=y�g�*�7��J?�
2��{?�"����	�?�=�Ң=� ߽{��<���=@��=^
C>��>m=6�=��<�%?��0?��%>-�?�d���{�Ub�A�>׺	�e�s���v?�@?@�?Ѕ?�	,?K��>��`=���7=����>F��>\bY�!�����Z��ۼE�����5?C%H?���=�@����>�� >{t�>B*?'�1?C��>Y!�>]yL=Ј�
۹�r�ƾ��:��n�ol@���.�.����o�>�5>��ɾ2�����f>j)G>w"v>"?}>Z>9�/�LH�=%W�>��>m=�d�=���8^ּ-��<�Y >�C�=
[r<�t=�3�=U��; p�����n��*�ǼT2ý={L����>�?!K��<��-�o�B��^j��\�>��?鴾>�d��&�#��g�'[���U�އ��#�L>��|?{.?gz�����=�=�=�_>���>�w�>Y�c>U�0>Ⱥ;�������>k�>�?���>w�.��x@�R��c��2h�<G��=v�&h�?Í�?�o��m�{J���}��vF����� ���W����1j�!M��|��þ��l�w>�T�> �?��߽b��>.KR�DN��aV�����G|��<��#m>�G=k���w�5��0(�aX�<9��~���Pu�>�&Y>���"�/?��>7�?�$'?�8?F���j>�'?.�>J&>�} ?e�T?�?��>7�?RK)�SŻ��n����M�t м�n�@2p<V@�>���=��n=ĩ�=���=�M��e^0�U��3>��:h��T�Ј*�GYD=5߃>��,?o�I?V�>�&�=��'>y:0� VE>i��>�ʰ>7꼽�^5���8?E�>��>�.a?��Y?Dԗ>F�=8�.�Vk�&+�
�.?#7=?�q�>u��=ܐ_>?,�\݋�2-=+a�=�&�'��i]��*a��*t���U>5�<�)���>��?X�J?ϠA?~Wս{���F��a{���Tݽ���>(2���K��{�]������D���O���<h��7A�����x>�&E��L�=�>?R�>ʁ���E��d�>����>�Y�>N? >�2ɽ��Ѿ�+��?J?��b���|��ȀݾU�H�� �=��#>x̽�5?!%�Yy�C���0'C�B%�>7��?6f�?&�l?�� �Ip�>�w>��w>6%>�֔<`�Wy��@��>�(>��=:���������y�b>�q�>y���ʾK9�+ο�ܯ���<�JVx�*�߾�aɾ�_����� ��=p�'=�R)��j���GS��3�����ؽ��\�����J���Z���R�?��{?�ꋾ]+m�D	[�7˾�tȾ���=�Y��`wݾ�ž���IË��n	�uSV��@��'��� ZE�x-��/M�>�1��[���I��'�w�7��>�
V>I�2?����\�2;¾�=H >c�����ݦ��Կ枽1�?��^?ߛ��Ծ��9�|�>�-?�I�>����vվ��V��)>��5? ?�� >B���5���hܽ���?�"�?R�G?|ݍ�z�o��-�:G�k�?_,�>�J�>�Z����߾��x�6?7a6?���>�}:�<ߕ���I��h7?Α?wI��!>Y��>5��>���qB;�)�������m=a�|>��I�NN[�vr�������=;��>��>���฾q�>Jq���T�pmV�@e�d|"��/7=�Z�>�7��D?>��0>��=\� ��v��`���}6�,�9?�{�?�PU?�@+?��׾�t��Kt���T�<��t>C�n>��=�$��u*�>Ӈ�>��ݾn |��.��x?Ҥ�?W��?*nO?�Rt�F?�$|���Ҿ�����N>SAP>�Dt>.f�U8�=�ʻ�[0���>=�A1>$�e>��9>��y>%�&>I�s>׺e>�7����&�����튿��2�����%��^��� ��Zξ��$�pV��'h��ԛC�-����$��x���yl���Gz>���>:q>��>�TU>���=͵{�f����̽Ǎ��H/�|7��kE	�������i�a���+=�=
C��7Y���?�^Z<�=��>ۊ�=��<�?\��=&�> $�>��*>�P>�$>��>H)�>����=��)>O=5H���Vr�	zo��F���	��L�Z?��H�uz�-�ɾ��z��6�=��?�R>|0�c��+��ñ?=J�'���KSɽK������>.�>|�	>Ӣཐ�����?/�����T>�9>L�M�����nH�),>��>������>ޱ>�C0?4݆?}Z?f�>$�?���>W�V>��`=���>ܭ�>o�>�?�A?�7?b\�>J��=�b(���$>�>�n���=��=gL,��h�;���;!����ۢ<�,>���=4�=�V>�Ϧ=��<>3�?�L@?��.>��>gyܾQۄ�����l��=p�>����l�X?�A?ʶ1?��>��?^�>�9>d7���b����>χ >S�y�O�����6A~>�>�=q�'?�j:?�I����y� s�>�f�>�R�>�y$?LtL?�b
?�i�=��J����l�' *���(�\���Cv=��>C���!�<�-Z�;����L��$���L>5��>��>
ؔ>�փ>ܓR>�u�>WH>8)u=RŻ	��o�	=��T��)=o�H�
r�<��=�i�ݐJ�̪n=#U�=l����l��@��K�����>>�?돉�c:-��������Y���d�>�g�>��?v>F��*�L�\���W�������O>#�?Mg ?���<�>>fH0=�� >R/?Q��>s��=�27=>�����A�5H>���>B0�>�DL��DD��rZ�����u>og=�f�:�?ก?��Ҿ]��n;���Z�tZ߾V���P���l��h\ؾ�� �SAO��c��w� �����<�>�q�>;�?xV�ݵ)>(y˾\
��X���]�1F��ɱ>���>��>>�I�ʕr����"o���W��>��)>�>	#>��?v�?$�x?9.�>�6?(6=��>�n?��>RM?X�;?a^?��*?N<&?�I/?�q=�)`�Ny���H�O�h�ݽR�=��2>]OM>���=�/=�8&�\ o��Q�q�U=�&��5������=���=��>)/?i�#?�3����P��#�޾�"/�~�|>��>�Cs����=�I?0�>��!?��N?*�3?a�>!Y���7�jž����D5?DAK?_�?���=z:y>@`������>`��=-�W�� ݾ��D�������_%"=���>7�>�>�A�?��u?�7?�%]=�����ˁ���g��I���@��<>����5�S�2�F��ZB���G�N}W��`�9>�v��ƀ	�xB���/>���=������6>,��>8�=�}�����=m��=$t>���=��>��5>?���k¾��'�I?[����j�C���%xо]����>k�<>���?���C�}�f
���J=�,��>���? ��?�Bd?��C�<2���\>�bV>)>x�.<��>��O�������3>��=Byy�������;��\>�Uy>��ɽ:�ʾ�4�٢H�6�ÿf��s�Q��|���Ͼ�w��6����߸L�������`4g���,�O<��޽����㧾l����΢??m�?�>c�~|q=�I��f<�8�
����>�3���ڇ�{��v�������2��m�m�z/i�=���>� ��6Z���C����w�gH�>��:>�RB?GT[��V߾��&�Ɇ�f�=�K��ھ��'���^����I��f?�.K?_��������ž_�
?ҋ?�1"?��?��፾�W>��=�b�>�q?7~�>U�ÿ������փ�?
��?&�E?�l���Bg�x�W�������>�<?�>���v�,r��U�>tK?��s>�lT�n��n�6���V?�Av?hLm�2��>P�+?ԭ�>Q�N� 	��1��ꟾ��>>��>�# �zc�ʛ�����"@=/�?3�>
ߍ��0�Җ�>`��5k���i�q��ZNл����S�>��i�V��=4F=	�+>C,�E���>���_ށ�J"�>�Q�?ᬋ?��?I醾�w�=�����"�B�[;�C�=�'ؽ�G=�#�> k�>���.��,<2�&?-��?���?��3?�f���ۿ�ɣ�� ����ؾ�� >�L�=2�E>�wr���]>�>�=FI��.�ý�h�=z?�>)�r>mb>��=0D>��&>|�����#�b���@O���,Q�~Q1�����U~��W�����s[&�*I׾Ц|��lǽ�t���H��V`��I����d$=��=�=��>nX�>�?�>׍�>{��=U�{��!�A�������鼾�2�V�6�@�-�t���꫾.���ýM����L�QN��Z?��A=�?�=���>m	��Q7>���>��>��>�)�>��m>؀�>[(�>���;�y�=��>:"����x>�.�=���EÀ���;��T�.�;\@E?��T��ߝ��2��ܾ�M���(�>Zg?\S>��(�L����mw�/��>I�)���l�%&Խ�>?�,��>���>��=����6,� �r��(｀��=�S|>�>�e��	���2��t��=P9�>q)�XW�=�K>J:?�΂?,MN?x-|=wJ�>w8�>B>��]��:�>it�>��>�
?L�G?,?7��>�\�=y�g�*�7��J?�
2��{?�"����	�?�=�Ң=� ߽{��<���=@��=^
C>��>m=6�=��<�%?��0?��%>-�?�d���{�Ub�A�>׺	�e�s���v?�@?@�?Ѕ?�	,?K��>��`=���7=����>F��>\bY�!�����Z��ۼE�����5?C%H?���=�@����>�� >{t�>B*?'�1?C��>Y!�>]yL=Ј�
۹�r�ƾ��:��n�ol@���.�.����o�>�5>��ɾ2�����f>j)G>w"v>"?}>Z>9�/�LH�=%W�>��>m=�d�=���8^ּ-��<�Y >�C�=
[r<�t=�3�=U��; p�����n��*�ǼT2ý={L����>�?!K��<��-�o�B��^j��\�>��?鴾>�d��&�#��g�'[���U�އ��#�L>��|?{.?gz�����=�=�=�_>���>�w�>Y�c>U�0>Ⱥ;�������>k�>�?���>w�.��x@�R��c��2h�<G��=v�&h�?Í�?�o��m�{J���}��vF����� ���W����1j�!M��|��þ��l�w>�T�> �?��߽b��>.KR�DN��aV�����G|��<��#m>�G=k���w�5��0(�aX�<9��~���Pu�>�&Y>���"�/?��>7�?�$'?�8?F���j>�'?.�>J&>�} ?e�T?�?��>7�?RK)�SŻ��n����M�t м�n�@2p<V@�>���=��n=ĩ�=���=�M��e^0�U��3>��:h��T�Ј*�GYD=5߃>��,?o�I?V�>�&�=��'>y:0� VE>i��>�ʰ>7꼽�^5���8?E�>��>�.a?��Y?Dԗ>F�=8�.�Vk�&+�
�.?#7=?�q�>u��=ܐ_>?,�\݋�2-=+a�=�&�'��i]��*a��*t���U>5�<�)���>��?X�J?ϠA?~Wս{���F��a{���Tݽ���>(2���K��{�]������D���O���<h��7A�����x>�&E��L�=�>?R�>ʁ���E��d�>����>�Y�>N? >�2ɽ��Ѿ�+��?J?��b���|��ȀݾU�H�� �=��#>x̽�5?!%�Yy�C���0'C�B%�>7��?6f�?&�l?�� �Ip�>�w>��w>6%>�֔<`�Wy��@��>�(>��=:���������y�b>�q�>y���ʾK9�+ο�ܯ���<�JVx�*�߾�aɾ�_����� ��=p�'=�R)��j���GS��3�����ؽ��\�����J���Z���R�?��{?�ꋾ]+m�D	[�7˾�tȾ���=�Y��`wݾ�ž���IË��n	�uSV��@��'��� ZE�x-��/M�>�1��[���I��'�w�7��>�
V>I�2?����\�2;¾�=H >c�����ݦ��Կ枽1�?��^?ߛ��Ծ��9�|�>�-?�I�>����vվ��V��)>��5? ?�� >B���5���hܽ���?�"�?R�G?|ݍ�z�o��-�:G�k�?_,�>�J�>�Z����߾��x�6?7a6?���>�}:�<ߕ���I��h7?Α?wI��!>Y��>5��>���qB;�)�������m=a�|>��I�NN[�vr�������=;��>��>���฾"A�>�4�f	N�vgN�r�|�;�ee<Z��>ƹ澂�
>7�U>xO�=�s,��Q���F��Ka�S>?!o�?��X?��-?��۾�GȾ�Ғ�4�=�>��>�F6=�윽�{�>Ͷ�>j�~��Q�?��?���?��G?�Si�L)ȿ�������վň��N@>H�z>{M-���ۼ�"�>;"Ľ����vr�>rܦ>ǕJ>���>O�r>�ql>%�W>zՀ�pf-��W��O㘿�e������{ℾt���R���?�<����!����W:�д=h~X�ZP���{�<r�7C�=�̹>�*?lC�>�ޖ>��=������	�n�E:�}�#����!�5��w���+�D������������"Ծ��>$�1�U�<�o�>�=�L>��r>ä>H��>i��>��{>�.�>�K�>q�>��>K�	>oP��C�A>��\=a���rs�r�l�0eQ��	��i?�[����xe�z3վɘ���Z[>e�?p �=�c7������'��6?���9�S׾`����q�@Q�>� �>vp�>?��������L�P��A�=�f>#�">]F�l����H�%/>T��>�̾Wr=u�h>P�!?��o?�u*?���=�T�>���>�+�>;��=��*>� '>�H%>h��>��0?��?��>0�=��G��$>���<�Г����꽜�$�Η=���=m���у=�=����K�<c}��]ݼ]��<L�@��?�Z,?#��>���>��о7�:���0�ܳ	>�n�>��q��M?t&?�?}�;?c�?YM>�M>��徉�I�\��>�d>�Ql��{�e�G{˼�+7>��e?A i?�z¾��>�5?C�w>f��>8/?�>Z?�=:?ش~>@������%�~4��s_��搾��<Q��>*o�����H�>�5��ʫ�nN>��>C��>��>�}�>�D�>�K�>���>��>������=:�0>���<�>[;g��=@$p�Z�̽Y_� Ŷ��,¹�,=��$���+*6�<�	?��>2=��ً���3�!L�E���Mk>!��>D��>�}>�?��� ���l���Y�*����g�>˦Q?��?� ��g�=oý�u�>i^�>��?v��=Ѧ뽰c���þ�)���8>!�
?�6a>�j�[�/��S%�=�;���">���=��ٽ�x�?�*z?��˾O⼽���[g�QG��N;��<��ట�L�C���O�r����羾����>7B�>r�?������)>A9��D����r�4�ܾ��X�.�὆�>�>���U�� ��e ��i���%��Rj��i�>���=)��>��??^$�>M��?_�>��E?��J�?�ޖ>% �>}?��F?��R?k�?�>*?$;?:�=/R�v%����ER,:�x�>B:=�>�>�F�=��k=g���=j��=y1���ܽ�| =W/%��s[���<��6=g�L>��(?fC?��[��H���_�=����>���>�[,?
,�e�=��%?i��>^Q�>��`?m	6?:y�>j��=r��2\վ�`�=}/?�&I?�?Q�E=u�)>u���3��Nі>@#��\ɽ��F������ƍ��
!�i~;�H>�a�=�"�>}�f?Q�t?"�??5�=���퉿x�<���;9�O�
{O>2l������G�)�O��c���P��+��n==��{-��>�9=6|>��!=V#�=G�>�=�LF�=��=��=]�>��`>d��>-�>,Н�B�s�`@���I?ޏ���i�9򠾆oо>��	�>��<>��-�?.����}�[���F=�%��>Ǆ�?Q��?�@d?�C��+��\>CYV>
>�80<��>�rE�ǭ����3>�"�=�y�5�����;[�\>gJy>O�ɽ3�ʾ�.��H����)Q�eGQ��^侄k��G��M��Y/���H���<���^�)�h�s�i�f���k�U���$��0�ҾR諾�G�?�r�?��=I�;=o�o��a�����2�>YU��-U��ڼj��=J"��C Ҿy݇�"JB�Y�g���D���S����>Ռv�,ް�:m�;_���?�xM>��?W�4�!	���t�W�?�}s�<�	�<���hl��J2��ȣ��g_Y?��D?>4��Vw��{+�=w�>�-?;�>�b��&�g�j�=�8D>VF?�?�;>�ꭿ\ꇿ�-����?~�?KfF?+~���Y���(���0��R�>�?c��>�m��Z������;�>��?���>̪D��q��W�?�zDZ?�_�?�}M��>��1?��a>��
�g�*��s���� ���>2ʟ>t
���1��L���Ծ�X��:�>��>���[j���g�>R���"��ݤm�q=�� ᾳ����?g��(������>��|;�rQ�K���VW{�2�i���o?֥�?k�Y?S�0?�YݾB�پ�;>qM>�r�>��Q>Ro�=��[�K�=G�s>��'���R����"?;��?ۚ@`��?����ֿ�����Sƾ�\����>xM�=ei>����O�{>-��=���<A��<m�j=Q�>��>V[q>U�>C
�=O�=G���3"�4죿y���.�>��v
��B�rq�s1�l<a����Z��ʾ��C��긽�9"�pa��*8�v�=G��2�>��
??&�>�MV>1�_>'�>�����K����+���L�W9�k��۾=�%��4�3={¾V��+ :�\�?�����j=�2�>p�=���=dہ>�:>H[	>J�0>��0��e>Cex>Ds�=:>�>y�~>�?�>؊>�i���d���I��D��\�>L�?��ݾs
�R�����Օ>�NA?�?h:��s�ct��E�b��ϩ>6]@��P�{G���N����>,��>Q�V>�������=�y���"׽*M�s�X>7�>J诼��-�-^�N�i�K��>�K���-k>a�c>Q�?�J�?��4?�Y�<��>�cd>�'�>�CT>�D�=��=�P�>%e?S�+?��'?�]�>M�=(WV���o=�r=Dl���[=ؙ �S����!=9A+<�ռ �>V�>��a���9=\42��������eH<[�?b#?�æ>�4�>�7澋t� �ӾΖ/<��>�W�<\B?�f:>=?+�
?�\u=�F���E��nܾ�
]���?�g�>�듿����{|�>��_>��T>
�?���>-�ž�Ӄ�������?H�(?�?���>c�> U��_m������x�4�HF��D�*>	�>��Ľd��/���X<QാI���->6�>���>���>y��=�O�ޘ�='�>�?>�v�<��&>=�<�y��2ǁ�F�=On��ֲX������Ҋ�=e�'��!;�c�=�Cx�
�6�/�8�/?�p�>����c4�%U�Bܧ�~���h�>��|>�$?���>/�>7�"�`#H�B9���9��?�V?��?q*e�$3�<���=k�!>���=�a�>�G?��� ��帪�V�M>��?��?�b�>b�ϣ'��)b������=��=;����?�5F??6�0uȽ�U����G�����k�t>!<�=�������*��T�5�՜	�I	��'���>�?���?��i�&=r۾������s�v�M��[�>�Yo>��?½�=�Q >��ֽ��0�<� ��)��#�G���>i�=��>>�u?��w?kO(?�?�k�>�s�x��>�V>!y�>4��>!m?��?�hL?��?��=���jɾ�B8���:�� �<��B�<�?>��>LU�=q/�=.N���=�H>��?�i��=���=3^�=��2>���=�s�=5�)<(�
?	�%?r�>���=qվ��E��ǔ>�1�=�٠�e�to�z�S�3G�>0?~�D?D?>R����W)�<˲�=����Q=_G!?fB8?��>^g��ǒ�4�L��@>����sc�=Ի����8:5��ξ*o"=���l�?��Q>�8�>,NZ?�}M?�U?%^�V�޾J@"���N�v�f>�Y׽�3>��>=e=�\����2� �>��}V�p�#��D�= v�n��=�>j�!>ZJ>�k�=:��=��\��P��'�d׽��@�H�>(�>X?V"g>��=�"ľW��yY4?|(���=�9���:]	��S�;�r�V*�>���!<蕖�r�{�s�����l��#8>�I�?���?�Ē?.�߾�8��Y��=s�>΁>�����j���{���3�=��>$�7�x�]��+ >�F�=���=�}ν:%�������x:���bL�|e"�m��/i��I��[)־TJ^�P���Vؽ�� ��캾\=0�<���U轥�[��Ҵ�f���)���??�?B_�=��n+)�J�2�l�����=6B`�B8���B(���̽(�������0��P��2@������ᾤaE>�J��ۊ��������M��N�!�f�/?�������q�ྵΌ�B6>��:��,�}Ɣ�߮���	ƽ�yK?�|X?�#��f/6���Ⱦ�İ>G�>�5�>y[y>_Ҿ�I����>�QE?���>L�߽������l>3�?���?��^?�<ں� ��0�K�>	?3B�>1��>�-˽�]�=�ý�V?�?Z̉>p���:v�į����>���?�8�.->nI?�>�ǽ}��92��r��S�=l˪>�Ԏ�������	��i�A>4��>��@>FVl�+����g�>R���"��ݤm�q=�� ᾳ����?g��(������>��|;�rQ�K���VW{�2�i���o?֥�?k�Y?S�0?�YݾB�پ�;>qM>�r�>��Q>Ro�=��[�K�=G�s>��'���R����"?;��?ۚ@`��?����ֿ�����Sƾ�\����>xM�=ei>����O�{>-��=���<A��<m�j=Q�>��>V[q>U�>C
�=O�=G���3"�4죿y���.�>��v
��B�rq�s1�l<a����Z��ʾ��C��긽�9"�pa��*8�v�=G��2�>��
??&�>�MV>1�_>'�>�����K����+���L�W9�k��۾=�%��4�3={¾V��+ :�\�?�����j=�2�>p�=���=dہ>�:>H[	>J�0>��0��e>Cex>Ds�=:>�>y�~>�?�>؊>�i���d���I��D��\�>L�?��ݾs
�R�����Օ>�NA?�?h:��s�ct��E�b��ϩ>6]@��P�{G���N����>,��>Q�V>�������=�y���"׽*M�s�X>7�>J诼��-�-^�N�i�K��>�K���-k>a�c>Q�?�J�?��4?�Y�<��>�cd>�'�>�CT>�D�=��=�P�>%e?S�+?��'?�]�>M�=(WV���o=�r=Dl���[=ؙ �S����!=9A+<�ռ �>V�>��a���9=\42��������eH<[�?b#?�æ>�4�>�7澋t� �ӾΖ/<��>�W�<\B?�f:>=?+�
?�\u=�F���E��nܾ�
]���?�g�>�듿����{|�>��_>��T>
�?���>-�ž�Ӄ�������?H�(?�?���>c�> U��_m������x�4�HF��D�*>	�>��Ľd��/���X<QാI���->6�>���>���>y��=�O�ޘ�='�>�?>�v�<��&>=�<�y��2ǁ�F�=On��ֲX������Ҋ�=e�'��!;�c�=�Cx�
�6�/�8�/?�p�>����c4�%U�Bܧ�~���h�>��|>�$?���>/�>7�"�`#H�B9���9��?�V?��?q*e�$3�<���=k�!>���=�a�>�G?��� ��帪�V�M>��?��?�b�>b�ϣ'��)b������=��=;����?�5F??6�0uȽ�U����G�����k�t>!<�=�������*��T�5�՜	�I	��'���>�?���?��i�&=r۾������s�v�M��[�>�Yo>��?½�=�Q >��ֽ��0�<� ��)��#�G���>i�=��>>�u?��w?kO(?�?�k�>�s�x��>�V>!y�>4��>!m?��?�hL?��?��=���jɾ�B8���:�� �<��B�<�?>��>LU�=q/�=.N���=�H>��?�i��=���=3^�=��2>���=�s�=5�)<(�
?	�%?r�>���=qվ��E��ǔ>�1�=�٠�e�to�z�S�3G�>0?~�D?D?>R����W)�<˲�=����Q=_G!?fB8?��>^g��ǒ�4�L��@>����sc�=Ի����8:5��ξ*o"=���l�?��Q>�8�>,NZ?�}M?�U?%^�V�޾J@"���N�v�f>�Y׽�3>��>=e=�\����2� �>��}V�p�#��D�= v�n��=�>j�!>ZJ>�k�=:��=��\��P��'�d׽��@�H�>(�>X?V"g>��=�"ľW��yY4?|(���=�9���:]	��S�;�r�V*�>���!<蕖�r�{�s�����l��#8>�I�?���?�Ē?.�߾�8��Y��=s�>΁>�����j���{���3�=��>$�7�x�]��+ >�F�=���=�}ν:%�������x:���bL�|e"�m��/i��I��[)־TJ^�P���Vؽ�� ��캾\=0�<���U轥�[��Ҵ�f���)���??�?B_�=��n+)�J�2�l�����=6B`�B8���B(���̽(�������0��P��2@������ᾤaE>�J��ۊ��������M��N�!�f�/?�������q�ྵΌ�B6>��:��,�}Ɣ�߮���	ƽ�yK?�|X?�#��f/6���Ⱦ�İ>G�>�5�>y[y>_Ҿ�I����>�QE?���>L�߽������l>3�?���?��^?�<ں� ��0�K�>	?3B�>1��>�-˽�]�=�ý�V?�?Z̉>p���:v�į����>���?�8�.->nI?�>�ǽ}��92��r��S�=l˪>�Ԏ�������	��i�A>4��>��@>FVl�+���xt�=% ��T���Y�"'���~�������"2?�^
��Ӈ�Zd>J��=H6�P���s��)�ދa?�7�?7T?��E?ēվ��־�5���<�>�OD>�U>��\=��l�fl�>��>���������q�Q? r�?~�@�n\?�E~�P ��O���r�VZ��ۄ�=8��5z;:��=B��=��3�覤=#�2�=��>�H>cb�>�R>%Re>�>���6C���񝅿=�M��,��0��ސ�m���:������˾_q���=�x}Ľ4���'��~����zs�F�뾿 3>���>'��>"v�=٬>95,>>\�����%��܊�Q�������ι����b��1!��j־�V����Ѽ�(��b?�^¼2%�=��>�4��psx>�>ڤ6�i��>8p�>�o>�~�>%`�=	��;\>[M�>�T>�g>���=>��-]���B*���v�j��<S�4?����X����P8��#������>�+?>�>M�꾠���+`�;��>g�<y��� \y��K�<���>�c�>Ag\=f�Ͻ����G��>7�>>�� >g�@��Ǿ����%��=��>�����O�=�[>��0?��v?��&?F�G�U�>�ע>8�>|A�=�G>��f> `>��?��2?��8?�(�>㱸=�nL��
�<V�=sg4�8	t�N�A��_�ąؼ�2p<���U=:8~=��<��S=�<B=A����@�;��;N��>��8?qJ�>%-�>��:�MM�1$J�ö�Gg�={�M;�	�>��>de�>���>��>�'�=�rT��M�� N���?�`z>t�r�$��2�>?&e>�_E=��M?��S?^!>�[�����=���=,I�=;�??'?���>֗�>��������hӿ^�#���!���Ra��SJ;9;��DN�y�`��E-��a�����<�[>��>�Np>��D>��>��2>�B�>�zG>(Á=(��=x��;I�;
D�7cN=O����8<0wT��~���f������s���IM��C����ܼ�E?��y?�*��o����@>�Rr�M[#�r*	�B��?Ib?��>!��>Iɾ�7@��9L��s�J>lґ?Ku?C��-�=T5�&��\G�>fR�>�(�>�U�;�CP<�k ���o�t�M?Im+?���>�E�T�h���^�Ҙ�����>Uk�<�c�֨�?ͥ6?�@�#���5y	�D	F��}��e>$�/�Х����ƾ�:�8�0�>��7���Z-;��$=���>���?�$ݾ  b>��&���y�������-xf>/�?>X?/�퍼�B�Ѿ�81��3��[�&ժ=�#?��y>����'M?_L?ʘd?�p?���>yX�1Ho��>�SV?0)>�C?�5)?`��>:��>���=[;�;��;�@ �䬓<a��P5->"W=���=��>5ե<�B���Sq< �μf�R<�Mp�^�9=���=��==�=���=zz?�@?���|1�=�H2�4A/�:�='k弢L>�@Ƽ��%����=XS\>�?�!?�.�>P����ƾ]���^�4�=��#?� 8?C�>b5t<uü=����~��%>�K�=Uyh�җ��������(��;Ƶ�>�2>�I9=�t>{�g?�YH?�)U?w���
��X��zY���߼�±=��m>�?�>e>D=c���X`=��zM���C�6�$��<z�U`D�}�i��iJ>�Z8>Bn�>ģ/>�
����=1=����>m<M����>���>�3�>.H>o�	>Q�¾�NؾkV�>{����m���4��s�����Y��K|�>�5��gP>�������ZZ���=t�?��?݇�?P�>E�O����l�>"�>��p>l'��$X���l7>�熾�k�>&j>�7�� W���`!����=ې8>
�༭��a
�W� �җοy톿�
>�c�Y��F{�
yȾ�=��߽r���Xzؾ��B���M����k9U�[V�)̯�|��|Pݾ���?�oP?��ܽs�����/�Bs��>J����P=��tg����̾򐨽�Y��꽬��ƚ!��H>�H��]���ڨ=u�O�=���N������co���<��I?����J^	�;�1�>Ғa>�AC=��
�M��������߽�EY?�*U?nA;H�$��tH�N��>��?i �>�.>	����D��iTH>�;?��?��>�C���Ý��wi�<÷�?�P�?)�6?�a�=�.�l����?Ub?ю�>��E>����d��0y?ĪP?�?�����#U�U��>1#? 9��q���B?�?���ƙ��l�>�o��NQ����q>��>�`��.
�C� >�>�F�>�b>j�N���
�?��$㾄uv�X�q���L<���&龩k�>��
��D���Ь�����,�Oɞ�"�Q�� ���o?g��?V�9?��?_U���K�Z�=ο�=a�]>��T>�!>�z�����>@>k�����W�Ia�U�"?1X�? ��?�^?|�r�����q�Z�����J��=�Q�=��%>�d�8z6>0����sS��᷼�3q>��>�5>-�>&�6>2�>��߻D��������c#��@�<'�S�8�pֽ�����b�V�x�ľ�vӾ���i�7�0������н?�ֽ�^ݾ�w����?�_?��>6S�>��>�e�&���@��n��H�����@��j㓾��#<�#�-����|������?x���	?ډ��t��=�5?5�6��2�=�>�bY>�V=�{&�K1�>@r>�Z#>���>0�;>*"ݽ���=�o>���=���������0��L�B�!=�FJ?@U9�MX���2/�Uξ~��� �>�l?�K>��'�b���h�u���>�LP��,X��J��fc���f>S�>�$�=_����Z���r��]�oK�=?��>���=������AK�K��=���> N�� ��=�'�>��)?'�z?��C? �>i��>��R>�v�>��>�:�>�,�>K7�>�x?� -?�s?2i�>^!�=�+R�$jK=`p";�8������t���:S�X�ӐU�Y0��i+=�8�=��=?�="�<_�r�����7�H�>��7?>�>Tҹ>{;�.q-����l��=���>�N=��9?�q�><�?��?�z�>�$�=k�>��3ݾ�q��� 	?w�>%�t��P3�w�>��?I�	?]�~?$"?����K�?�6�>Ӥ�>[?��F?oP6?A��>f��=0Y˻���kjӿ,�#���!��������X�;H=�9Y�s��'.��_����<Iq[>칅>]�q>��E>�_>��1>�g�>�D>�f�="8�=-�;7rH;��G�H
N=���p�U<\�L�0c�������M�������:E���9��X�׼�1?���>^]��DW�
�������о���>q��>���>.�?\?s=u����kC�ߋB�I^[���>�&d?���>��ս�]�=Z���#��?�>�=���h����I�6)��^	?��6?W�>��"�I�l���]�c���~��>�e<�����a�?CC6?�"Q�뜾�	���O2�A�'~�>g!>lN���A��"�)�˾Y��$�e��Z���U?;t�?<���Ľ}ԛ�f���,s����;܁�>&��=��H?���=�:ӽ��?<��@����\r����B;��>�.N>*/#?m�@?T.W?�#2?�>?)�+?\ǒ��{�>e�?>��O>�8?!$?c��>%r)?�w?�=����24���a��z��g��88����=��<��>K��=Ӟ�b6�<��<3T�=� c�g���\>�"I>��S>�5@>����n�?��2?*w�=�C&=(��ީ���>*��>�ݐ���	=`Ǉ;��T>��?^�;?+�_?��>�.��Ug"�LQ��=o
�a\�i8?�.?��K>0�J�&^���B��������= ��<��i�e��,)�bA�^ut�{��<�Vl>��D>7�>��s?�WA?��/?�Q�0X�Hcc��P7���;���<���>�b�>��\=ŕ����.��n���X��E2�	 ��Ca��O
=Q�3>�"0>JH>�n�=��&>���8�����(sܼ������>S�>-?��>*v�=����7�
�^��>c�Ǿ�V��j��P�ƾ�a���鞽��>�kH��\S>}A+��7���X��Dyu�a�>tc�?̗�?�ז?;eݾ��ٽ{E>{|�>Js�>�1e���v��6>�C�@�}>���>�Ǽ���ˁY�?��>hժ=�;%��w��w�ܧ���츿z0��Xh>��*�ݾ���( �����R)X�˦�u�ھ	���Y�s�ͶP���ս{#T�M�!�,qj�t>���cr?��[?Ma������r 0�A�����5�=����`���(����l�����9k��d�ھ��%�g:�����P�G6q=o�S��3���-��b����.��@�tP+?n�K��C�?���H�>KR^<I�+������(��O�K?��:?o�ܾ�	��f�i�>'�?VY>�Ĝ=+����6�>��>e>?J?�W��҂�=]��G�=���?L��?^�{?nv�<T?O�� ��JZ>���>�?P>��k>��=.*�=�F>�` _?�~�>0s?�,1�ƨ��b�x��>b�?4��]�=�q�>O�
?42��������J>ov��{��Oa�7���+�������𻒻i=��>- >6�:�̾�g�>R���"��ݤm�q=�� ᾳ����?g��(������>��|;�rQ�K���VW{�2�i���o?֥�?k�Y?S�0?�YݾB�پ�;>qM>�r�>��Q>Ro�=��[�K�=G�s>��'���R����"?;��?ۚ@`��?����ֿ�����Sƾ�\����>xM�=ei>����O�{>-��=���<A��<m�j=Q�>��>V[q>U�>C
�=O�=G���3"�4죿y���.�>��v
��B�rq�s1�l<a����Z��ʾ��C��긽�9"�pa��*8�v�=G��2�>��
??&�>�MV>1�_>'�>�����K����+���L�W9�k��۾=�%��4�3={¾V��+ :�\�?�����j=�2�>p�=���=dہ>�:>H[	>J�0>��0��e>Cex>Ds�=:>�>y�~>�?�>؊>�i���d���I��D��\�>L�?��ݾs
�R�����Օ>�NA?�?h:��s�ct��E�b��ϩ>6]@��P�{G���N����>,��>Q�V>�������=�y���"׽*M�s�X>7�>J诼��-�-^�N�i�K��>�K���-k>a�c>Q�?�J�?��4?�Y�<��>�cd>�'�>�CT>�D�=��=�P�>%e?S�+?��'?�]�>M�=(WV���o=�r=Dl���[=ؙ �S����!=9A+<�ռ �>V�>��a���9=\42��������eH<[�?b#?�æ>�4�>�7澋t� �ӾΖ/<��>�W�<\B?�f:>=?+�
?�\u=�F���E��nܾ�
]���?�g�>�듿����{|�>��_>��T>
�?���>-�ž�Ӄ�������?H�(?�?���>c�> U��_m������x�4�HF��D�*>	�>��Ľd��/���X<QാI���->6�>���>���>y��=�O�ޘ�='�>�?>�v�<��&>=�<�y��2ǁ�F�=On��ֲX������Ҋ�=e�'��!;�c�=�Cx�
�6�/�8�/?�p�>����c4�%U�Bܧ�~���h�>��|>�$?���>/�>7�"�`#H�B9���9��?�V?��?q*e�$3�<���=k�!>���=�a�>�G?��� ��帪�V�M>��?��?�b�>b�ϣ'��)b������=��=;����?�5F??6�0uȽ�U����G�����k�t>!<�=�������*��T�5�՜	�I	��'���>�?���?��i�&=r۾������s�v�M��[�>�Yo>��?½�=�Q >��ֽ��0�<� ��)��#�G���>i�=��>>�u?��w?kO(?�?�k�>�s�x��>�V>!y�>4��>!m?��?�hL?��?��=���jɾ�B8���:�� �<��B�<�?>��>LU�=q/�=.N���=�H>��?�i��=���=3^�=��2>���=�s�=5�)<(�
?	�%?r�>���=qվ��E��ǔ>�1�=�٠�e�to�z�S�3G�>0?~�D?D?>R����W)�<˲�=����Q=_G!?fB8?��>^g��ǒ�4�L��@>����sc�=Ի����8:5��ξ*o"=���l�?��Q>�8�>,NZ?�}M?�U?%^�V�޾J@"���N�v�f>�Y׽�3>��>=e=�\����2� �>��}V�p�#��D�= v�n��=�>j�!>ZJ>�k�=:��=��\��P��'�d׽��@�H�>(�>X?V"g>��=�"ľW��yY4?|(���=�9���:]	��S�;�r�V*�>���!<蕖�r�{�s�����l��#8>�I�?���?�Ē?.�߾�8��Y��=s�>΁>�����j���{���3�=��>$�7�x�]��+ >�F�=���=�}ν:%�������x:���bL�|e"�m��/i��I��[)־TJ^�P���Vؽ�� ��캾\=0�<���U轥�[��Ҵ�f���)���??�?B_�=��n+)�J�2�l�����=6B`�B8���B(���̽(�������0��P��2@������ᾤaE>�J��ۊ��������M��N�!�f�/?�������q�ྵΌ�B6>��:��,�}Ɣ�߮���	ƽ�yK?�|X?�#��f/6���Ⱦ�İ>G�>�5�>y[y>_Ҿ�I����>�QE?���>L�߽������l>3�?���?��^?�<ں� ��0�K�>	?3B�>1��>�-˽�]�=�ý�V?�?Z̉>p���:v�į����>���?�8�.->nI?�>�ǽ}��92��r��S�=l˪>�Ԏ�������	��i�A>4��>��@>FVl�+���-2�>x�h��4N�=�:������> ?� �W�x��>$,>3h.��	��ǭ��g
0�3�@?cŮ?P?H�?K����ɽ��� >JX��� 2>�_+>e��>�j�=�Ԇ>肹>nu�6x���4T0?<1�?���?%�l?��u�5ֿ�t�����T���9y=J��=j0>`�N�I��� ,<�"�;�=] �=�	�>��[>%G>�b5>ݮ�>4�E>�����[�j{���Z��6'�#����D���¾%)�P�Q���B���w8��-8���t�-ְ�a�.�l�k��i�PІ�qs`=ͺ?Ů?�G�>�i�='��>rbJ>�n�)��%C�����߈׾da���H�;\@�Χt����:�	{K��W���6?d����p�=N�?�y��4�c>l}�>Հݽ��>��>i�
>¬�=S�=�Z)>A>�l>�6�;أ�>��Ľ\��A؈���G���S<���>t.?��Y�J ��b3���c�o�5���
>�`?t��>}�/��h:��?M<��ɾ�Z/����[׫>���>���<�]�� 0]������/x�g8M=�
�>0=)��������"�=���>����*>�J�>/?�~?U"8?x�>���>��>V�m>��1=i�G>�S�>��>�g	?�}?r ?c?o'�=9�h���->�R=T~7�K�T�[A�
�W�e*k���㼵�۽J�0�Bu�=yF�<�:�ꬼ�0A;���=O��<6?ԁ>?x��>��?JLZ>�K�Ɔ��⹽�0[~>(%����T>�ă>��?��c=�>�V�>��Z>.@���B%��>g�}>%)?�]3��b���O
? \�>�*?@m`?��=����(E�Eѭ>%�>�H~>#!?�� ?sТ>֨�#����������B������}��^��(@����>��~=�*��mL����=YM�=՟�=,�7>�Ӈ>��2=���>Y!)>�4�=�ı=K_�:��?�(O�=�Hg>E�e;���4�!�*Oy=M"�<�g&�]M��j���R��2Z==�	?��<?[��<���5�=	پD�(�H�?��3?�C!?4_?$u�=����i��os��\5�[#N?�_�?��>5���r>ȅ�<��>�>ǌ�;]�=�Z0=��˾I�ھ�� ?O�?$�>��>9}p�P���f����"���/?;��==�-��/�?�Jd?�e�����$��U��|�Z
���#���LV�����K[��)��Ր�V�y���F�S�2y�>�7�?�2Ѿ�Vs>4���T��	����+�9Z��	�{O>�(;�b�������.¾�=��=Q4< )=N�=��=c��>�o1?�7�>�x?ܹ6?�1+?f#��;��=iC�>�_.?�!?���>�f�>���>�s�н]�~��2��t<�@���zf⼄�`>��=�΅=T_>t�o>�|>�6_���=b�$>��=���C�<ٴ=>�ҟ=�|+>�(�>m5 ?�v.?I��=_O������!�<C��=U/��E�=�c6>�X��&��<)�=>u�?�?�Sj>�ļ�r��w��4�����=A?�c:?��?�J��y�8>w���$Y��u�>VΞ>��-�U3�������T�[��� >%�}>�K<���=��?~y5?�g?7F�>�)a�����f����3=���=R?r9?4���1�P�j�v���õO�(3C�U@4<����,<��=O���q�>�`>��=4k����p:�so=�Nڽ���<�L�>3��>���>���=��'=\�����EH?	���z���9���{E�<뱃=*�>���>�aQ>ֳ���p��&��m�/�Z��>!�?BE�?.�L?��o���=�x���7>><m=�T
>�H8=2�����=Pr�>N۪>|
��7��GDr���>���>(��<n���<�[��=���>���'�>�ξ���T:������ü[/��h����̾T�ѽ�ؽL6�F����2�×���Y��4M��3�?��o?�笽�{��(������A����젤�<�F;H���{W��&�����3:����־ũ�U~(����D��>
'Ⱦ^2��D
{��6��*>���>j"?���������e,�ᐌ����=X�>�r��K!d��a������k i?��-?���h�̾[��<4�>cT�>�Ҳ>�_�<���B�j��>)>�>o�?Z�6>�J���ĕ��w��S��?���?�i?��&����/2��Bݾ�I ?�q>?���>E���L�����!��-���?�q?p��=#y@��S?��?Z2�?Oc��ɒ�>%	�>o	>+����8Ͼg��� o�b#̽�������	�w>0��I�e����a>��>��ǽ	����?6e�:傿��!���Ͼ�b">�`>�u�>]��0/�>�Ľ�"�>|p�������n�c��Pa?�u�?�S?GT2?�R"�����"9����>?��>G �=��m=�G�n�>��>z��wC��P�!t?y��?S�@L�_?m=��1"ӿF���荭�b��&gQ�V�e=P8>�½<��=Z�<�5�>2k�=��/>P�>�Q>2A->��6>�A>#��=8���'��]֫�]���o�k�����I�hO�"�߾ޜg����")���՚�M�;H�н&IS��7W���&�Z�*�$����>h��>顷>#b�>XQ�>'�>�%�c���p\�ġ�y@L�s�1�����M��խa=1�I�d��������6���?5�/�w�g>~"�>���:�]�=�f\>D�3�>� �>���=E�>�C�=A)�=S��=�I>r=�z;>]r�=��{���v��'_������&�=ĺP?IQ���񏾥�$��MӾ#���J|�>�l�>7�1>�� �`I���Nk�,>�>�:Pf��:8�)A��q3>�;�>LQ >���]�e��w5����%>M�>�]a=w�ؽD����N@���>��>����>0�a>5(?_�w?C�6?���=J��>BT>I�>S?�=-�5>��`>���>�,?p�9?Y�.?,)�>���=5p��Ԣ=��<=d�I��P7���~��X����;�.y�8�{=��c=��<Q"D=�a�<d����e</z�<���>#[?ŭ�>���>�u ��X�2TH����=&�>ȱ����	?E�?}�H?.d?g��>;dm=xo~���4��s�>���>˟t�鷏����=ٲE>�C>̾?z�r?|X�>�)����>|��>iq�>�>�W*?u?>%�>�k��F=�zb��B
)����<K��I��=��;=�߾,����2I>)4V>W�Լ��>*�>Ej�>ؿ�>3��=�=���>sG�>�E�=�ɺ=��5>���=,�=A�<Rt��Л��>_.���Eq�"�9�P()��s �op=7�;������=q`
?@94?�:�=���y>�F�m�B�ˇ�>�O?m�P���<>Bl�=8f�L�g���y���ؾ�?
���?'�E?���� >Q�h�cI�e�?_=�[E�p��>�s>�5n�^:Ƚ071?SI?�J�<����E� �!����>1�=M�,�L�?��V?���%����m'��d�`�Ⱦ0O�����|$���`�eV�?�����C�����=[�_=v��>j��?�����=��_�?#��&�������H�=:��p��>=��:�]��W�J���Ǿl�Q�H>���>'�I>
�&?���>˕�>�6|?i.�>��>=]-��1D?�Q�>� ?;�?&.?.�f?��>
.�=�+�>�E)>��n��<��Iľ$�E>σ�>���<^�J>h��>�Ϝ<]]�}�:�6Ev>O��~ȯ�^�<v��=�٤<ad���G>k}�>��	?{�?
C��-廁;���J���u=��=DS[>��������Խ5��=�,�>bx1?�:�>s�=�c;u
�q��i(4>�?��?��?�6�<��=���Q'��[�"=�>0�m�s;�0Q�hQ׾��R��H>>=;e>���=:ߌ>ӓY?��E?�\U?S�|>��5��v��g�>�?v>_��L>���>���>���V��	�Y��,$g����L�ki� @>q�>���w>���>|�u���U��h����<>ҭ�.1�>AX�>c-	?ޜN>]>+茶�H?���y?�I���_ݙ����T��>���>|~|<��k���[?�����f󬿬
�� O?`�?޻?�$?oo⽖P���H�>��>�i >�.�����/o��?!��%�>Ѣֽ/���W�O	X�dq>���>��O�m������Ov�[ݛ�]:L�ɧ��w��/������5�8�o�ʾ6H�=M���㼽�+o��sW���z�Ӝ���.j��ϥ���`��L�?e�t?��=+W��4�^��,����~)�>͍%��;߾���{%��ّ��q��P���8�!_�i 
�m���>��5�����	nh�vNF�������>�)?r��rW��:����=j�>R1�= ��M��K�#�L�#�i?��b?���u�%�0����$�>a�>?`��>G^位݉���=�`���qA?��+?�Y�����0�|��$�;b�?X�?c�??��I�\U@�����]���?��?\\�>����:�Ͼc���?ۈ9?J��>�H�8����;� ��>L�\?�^M���_>���>JǗ>����ߎ��L�.����e�T��:>:#�j���^���>�q7�=��>'�y>�rb�׮�ȣ?�������3+��Γ=�3>t�E?L�Q_�>:�>K��>E�2�T��l�����P|?@��?T�I?W�??r6�{EؾN޽=��>�[?0<Y�R��. ���l>x�>���͌���+D�>���?���?��Z?�`��w�߿�����}�����*��؂��|*>B��e=�_<Mg�=��[`	>0+�>˖�>� W>H�>ϋb>L�2>6����P���������*b�i.<��=���M��{�:��R��蟾�:޾�)D������<	��BW�n����t��/��m�>2��>ّ�>�l�>�G�>v?�� =2�O���q���=��K��CG�*�`�F���н�ʪ��Z�&KѾ﻽�����?�,l=��>"�&?��T�C#���>W���_�>���>�-s>���>Q!Q>���=J�>��w>&O�=�Nh>�O�=e6�����OC��׌�B_>�a?i�����>�]�V���ӾB���!h>*��>��9>��#��잿�{����>���<����K!���6i�^�^>��>负>��߼q�*�#>���O<G+7���`>7��=m�½�'��.���y��=��>�����,>a�Q>�?��t?k1?5�v=���>��>�@�>?/�=�p>��>�H�>"?s+?��1?(U�>)��=G惾��=a>��5�캽�-ֽȖ����:��8/�9��L�=L��=��S�s}=�9=������2�H�T=��>�8E?��?wʽ>9�B�BYY�d�X�`Э���?J,��|��>K?��C?��?-��>/>2�Ͻ}����@4����>���>B�7��=��_(н4��>@�>��Y?��I?�$�>'=E������>��>��>nu?t(+?��>�$	�[��O�ԿC�	��$�T�C�	b��	=�Y����O�x�<�T�I���-N=;��>�6�>�b>U�U>��&>��@>=��>�=>��}�G	�=5�>�7=�����.�'2 =Vs>r��%�=��̼��Խm����p|����oν��=I��>�)?m��=����l�z�$���L��U�W>�E�>���>Mͱ>�/����]h>���I�����`�>F;q?ײ#?��B�D�)>��X���Y�DB�>�?�>c��=������ihw���>���>�?��>��a���X���u��
��a�>��c=:�г�?r?�޾T�II ��iJ����i�����=M�޼۾W���;*�U	�aFԾZ��!�=k��>���?ۧ���O�=h��Cؒ������Ǿ�� ���R���/>���=RR��WM߾d`/�αؾ���(7J>��?N_�=��>�aQ?I��>�d?�N-?��?L���y�?��o>��G?Zơ>��,?Sv}?^�?��q=/�.>5֧>��<j[ �)��t̓>U�>�=<S�=[�$>��=S���DA�E(>�l=��
�u�/��7�=!A=��<�t=%*>F��>ؗ3?��<����W����T��f�=�l[>n#�>��=>&S4���=�Ѭ�>�L$?tE?"l�>�,>#�X�`)�:���/=�C�>A�?�:�>��*>�R>������V=�o�>�޽�2�������+�e����=�$�>��+>(q!>�-h?�?�?��?�'�����$�*����>�N ��1$>Z�?� �>8���[�����O�����P�U�>�m���Ž߻�=@�>���<`-$��HU> Z>=[1:����b4����=&��>��>\�>v��>P4<�پHh�k�y?�j6�ÆK���������=6�>|��>����>F�⒖��y��fK���@?��?º?�,?�G3<�Ɣ�2D�>;e�>�V=g��ǯǾ���=g0h��֪<�A�=�����F���0�<Z4>L��>ē��:��'��q�zS���	U���Y��G¾��9������t/�:����	��`o�=���֗&��v�a�˽�8�����l�a�������u3�?2o�?���+!��[9��t
�tX���G^��tE�}p׽��zK'������۾b���0�>.�RlD��:+��՝>�y��'��lu��IZ��-��97�>4bO?'��ح"�V�D�#\V>�>.�:����Մ�����'�3��/J?~s;?ղܾ���a�H�R�!>]M#?X�>jY�>���?������>��R?��>Uy�����������>�F�?~��?��??�RO�k�A����r6?�?���>�x����̾���^?L�9?)�>��f���9���>��[?/@N��-b>.��>�B�>!#�~����%��N������9>�s�u����g��$>��ڧ=��>7x>Uk]�pخ�ښ�>h���l�}�����6�Q�� ߾��	>��@?`�k�N"�>�	>���=�1�����b���;ͽ?�h?O��?U�h?��%?������f�=���=�K�>]_>� \�� ����?�j>�7���jn(�a��>r�?�k@��f?˱s�N�׿9>��7���u*����8<�8>��>o��U�)Q���a&>�$N�Fz >2�m>2E>͊h>��C>� E>��,>^X���"�A��MS��-��q	�����Tؽc�ྫ�A��Y�O����h��N ��՟��.ް�L�H�Ab0��v��@���=��=~_�>�{�>��>>H5�>;�>q�H=���v�Rd>�P?���7��e�<Ζ�/���4�����5��V�����%���?,����~�>��
?����=�n�>��>���>���>��>�y�>���=JO,>7;>g>�b>膇>JA�m��EvS%��}4���/>�{>m!ھ|K"=h"R�!��*4�A5=(�>�8>��%������}H��/?��^�����(o��Uy5�q�n>j!?�z<͐ӻ�M�G w��nX�Nl3=JG>���<���������peB<�3�>!�ᾟ! >{�>Bx-?.i?K�1?�=�>l�2>.�>0��=~�>�1t>�֎>�k?A�2?*-%?�y�>���=�HO�HV>G�=������$��nB��rX��h���7���"�=S�=m\�;>�;�䈻����9�;�=i�>T�J?\�?Y��>u��;��>�'`ؽo�c>�Ͻ�i#�>�?�O1?�$?�.�>��<�6�ci��3v!��P�>�J>&[���͒��ü@o�>�/�=_8?�W?xs>�?R���<��N=A{a>v}�>C�#?P\?f�>\a=���s���.�ھ�����w_�	uؽO)>(>�0T�s+�TG��(%��pF���9>:��=��=�N!>�ؤ>�yS=�w�>��>����;�#�.=&M�<|���<�~ƽp��=���YD����?B�.�����;8�p�"żX�X@	?nG$?��7=d���>Ԡ�B��O�����>�A�>(�z>&y�>��>���o`�+�S��͏�{z>��U?�?�J��rS>�a����+�Ӯ�>x�>CY>@{c=��&��P�9-�;�H?�b?���>4���LP�� w�=����>�&�=m;��G�?50N?��q�6�BP3��=��h�x+��H�=�?�X���1��"A��S����HX]�d��=���>a1�?�N��Q7��m��1��n������ikl>9W(��G&>3k�>)O�b�&���g�����JӾǣ7>]�?>� ?�40?( ?rJ`?��?_�>0S��sL[?����R1?Bv�>5�;?w�?7��>X�?;"�>�=?���w�������>���>d� >f<�=?�>�*P�v�!��νP> 63�x9Ž)Ǣ�f�=��=s+��{H�=�)3>/,?��?�U���h��5܈�� ����<3H7>��=ŀ߼�)��G�w��V>���>Ղ+?�L�>|jw=L=ӾB�����{>S�?}�(?� ?���<���=�;۾�풾V�;*��>⢔��[���}��ͩȾ�ZC���G>��P>�k=��k>9ː?C9U?¯�>�F�>� B�n8���z��5�>P��6>(�5?+X?W�W��Y�L���Li�e<J�ޕ��&>�o���@(K>���>���Г=���>Uh��F��Zf��h�==3�K��>���>E?��>��>&����&��v}?���N�/�W*#�����E�>է�>�O�� -� rD?,�Ӝ�������v[�rG?�p�?⺳?�g?+1=}O�c.>D�?���<I�<�N2��#����=��Խ!�v��3S�^Yྱ҄���r>~��>uA%��R��iʾ( #�I���{�G��	��Q��V�q�������E�
�H��fǾ��=>�꾠����`] �x]��M
� ����i��02��E�?٫p?����鈾����������&qŽ��#����=��ܾi�<i�� |����u�����U���7�����.w�>6z�LB���Q��<�D��jh���>B?��־@쀾~@�.>)�N>�˓�2<���́�zS���!����`?��?Ç��p���6�d=���UH�>��>`��>�L�ؿ=����>��!?&�	?C F;����琿D�=�(�?Zb�?1 @?s�A�Q$J���t�k�N��>V�?(��>d>����þ̰�ܿ?g?5?)��>���΄�\��;��>�j?}k�q?�>��>F�>W�
�w���$߽7A�>:Y=[�&>~}�=Y�A�����}�F�V=��>�F�>7=��◾c.�>�몾��h�߃A�ćs�l,i���B>�%?ɾ	e�>���Hew>�� �ߗ��!ᅿ�����m?]N�?��B?�Q:?*����9��F�c>��>��>bf>�d�����>��>&B'�p����N+���?~��?�@)3�?�9g�ֿ0I��������ύ=Y<�=�U>Z���o��=���	.�~�^<��="�>�Hq>��J>mvP>�	X>$�6>	��Te���ꑿ��C�(0�����T[�Dp ��w��(h�{2��4�;��!��Iս�ڇ�ã�4
�=c�xʳ��t+>
�>_�>�*�>7�D>�h�=�@�4�1���L�{���n.�V�)���x�B�U�C��=q��9������6�k�@?V{�=Ӡ%>s8�>��a�c��KZ>\�߽M�(>��>�=0��>��*>��=��<���=.ѹ=W͖>���J���?����/���R��=$�8?D�f��]����:����K����n>��?tpq>F�������$o��x�>�`:=�c����6����5*�>��>�fu>�Q����d��5 �=8��=��X> =!����W�^�ͽk->�`�>ϯ���b=>�>�>?}�|?�}:?V��=!��>�Z>ǫ>�B�=�0H>��>{�>��?��3?�m,?B��>5��=#�{���@�_@3>�J>�r�(���=�U%<����݅=���<s>�=p<6�<�Ε;��f�������=�d>�Y�>i?0X	?��>;id��X:��y��R��?�]��g?D;?�9?Ev&?���=�C��ξ3S����嘔>tbd>_OB��8{�$�ڽ�K�>�� >1�x?�=?�yK���ͻ��=�j>���>��?�"?,L�>Z
"=�?�¶��ȿ�O��W�N��<ڑǽ�{>�V2��)y��=�dM�����w�=*7>�=>��a> �i>��=�>��
?6��=�U��o�	>�`0>n��<�	t=�1������_ �>_�Y���G��=����s!��1�<�����ͽ������ ?,"?,O�=��9�$ i����쩾���=Re�>>�݄>�m=#����0��FS��˧����>װ|?&�>ё��ĊW>���t�ӽ�~�>u�>��:�����$��Y��߽�p>�>t��>5`'�c�g�C+�����zȀ>@�<�u���ħ?i�Q?wA��P������p���%�L���,=�9ͼm^��n�����=���?���Cڽ�E�=C��>�&�?��\���D�-�v��ҏ��B\��}� �=�i@����>�A>(mݹ_*���Z��p(���ʾJ��>x}�>�i=�W�>�#?�i ?��J?H\�>�*?^�����>Àd=��8?��.?�?�Z?��>�1l=1�K>�K�>��d=l�7�9�Ǿ�cb>��>��'>��=[">#��<@}���=���=_W�;к <���������=0��=g�=��c>�A?��5?�,���I�}䛽���T�d:���=T�>1sܽ�R0��e�=�И>6�?@>#?�L�>��=	7Ⱦ5=��r����=��??oB�><�Y>��n>PѾ띱�,��=�}4>{���[ԾĲؾ��������=�>�2�>s�!>�+�=R�j?P>?8q:?V3���}P�V�H����px�jf�9��`��>0��>����WYj�A��T���?��Ic>���9��^a��E<�>�=p$�.�>Wmv=�K<��¼='���^�9v��>�~=�U?5�n>L�=e�˾sp�}y�?�c9�q�Y��P����>u?��&x?ջ�={#�>-Kn������ڠ�T26���X?���?h2�?GL�>9���g���¯= ��>���=���=z=��8ӽ���o��=+���/��YR�7�T�)>$'R>��&���SB��#	��-���X�L�w������f��־u@ �A�.��C���H=���@Ɩ�7����S.�$i��2��]哾v>��̤�{ϧ?4��?�Z
����ZL��O%�YLɾ��+>���S�����侮���n��\#���H��O�x�G���A�P��%a�>� �['���
���$Y�Ӎڽ<C�>y�6?�����J���>�p��=J>n�=�O�Yu��YS����o��|I?�C'?�ľoɾ�[#���>���>U(�>?�F>MEo��#�:�>9C?�O?�a��ے�Ma�>XF�?'w�?�d<?S�=���C�%
���Z����>(?���>)�����f ��S?�7?8[�>�3�����>J��/�>�\?|�I���]>E�>č�>/�_����/���4���}�n�Q>L|x<�"��򏋾Um�pK=_�>WW�>�/������>l���e��(�I�I�����W�E�:?-��r"q>�L>ڂ>�kJ�\���>���Ø�o�U?2��?�w`?��O?n?�]�ξp����2>'ֽ>�t\>�>W�߽t�>���=$�l�l�bU�f�R?���?���?0�l?��F�[տ\b��,��Q����=��;>��->K�)����<��=�t�;�� =O�>"q�>�d>��t>��F>L�W>�JK>�����%�����Mޚ�s�@�������鸌�4	�~WU��z��ͻ��x������)�m��`2+�S�u�d��;��(��˾=���>�?"�>��=Or;�܏��H������e�JO=� %
�8���bc��Hp��8V��jw���ɾP=��/A �֠#?@>gd���%!?������=(0�>���}��>҉>�{>D��=��=$�[>q,y>y�7>Y��>j��>r�C��`���ZV��>�F�0>�wS?m:��욀�qS^����	�ؾ��>]�Y?x��>Qz�O���) ��E�>;8�2hݾ���0B>���>�%�>d潬雼�,&��5��H�
����=@,?�=>C.�<KnԾ�����ԇ>���>�ԾJL�=ѡx>B�&?��u?c4?�_�=&��>�Y>c��>�t�=��G>�uQ>���>�[?]�9?�{2?Z��>�=��Z�S3�<��=��:�:�i��û���ݼ d$��<�o+��==_Ep=��)<�|\=�E\=[�����;�)�<=��>�G:?�+�>je�>yu��)��YQ���J��z�==�z���z>g�>룴>d��>'�>�;�>�f`=j�����lɴ>Z>�^�ą�p�=x�=0ۍ=&CD?r�?Y�9=X�,��ɕ���=<�{>��>�9?5`�>��:v;�����)ٿgK{���.�p(�<��><��Ӿ�,>�T>p��=��6>�Y�=��>��z>��a>V�>
�$>�:�>ь�>9�<>���<N.+>���U�_����<wC���ʽN��o��<����0�<�0����ǽ�=����=�M ?� ?���=[�`>+JϾ&q�U
�I�>�>�?9�?��R�q�沀��_J�b$��i�>a8J?�y�>(�_� >�g4��g���ی>���=�">�e��.¾��c����>FW?��>�\>R���o�N섿v����>[�7=f`��J��?�x\?%�-`�X>�y�2�a�
��C�� )����N;��� �=�)��r�1����ᵽd�w>��>��?��m��U��n۾P���}�m��:����=���> i�>u*>�fY�$����d�ҙf����=c. >=}�>�y|�zN�>ITh?�%b?yTo?@�?q�d?f"�n��>#��>�j?K�?�&�>W}>�2�<��p>���=���ν&�4��ڳ�*E=��=n�=�T>��>&���3�{Y����<��� �p�p=�BG<t=���G�=�˘=��>?$�P?$�<���7�D>�$��ؚ*�'h�>Vb�>���=����'�={>�>���>�[?���>����"&���J���Zo�<���>�3R?-��>���rZS��3��#G� �=|�C>'Ge�o��U���tľ�x:(R�>7��>��j>�)�>&��?��?��O>/{h<��>~R��{������k>�`?W��>���>��侎L=�Nn�M�s�}�1�(dt�c[�7.�=�R>�]��i�>�>�?">̑>Tߓ;c*�`������d�>:��>y5�>�ډ>Yb� [��]6��M2?�D���о(�ྣ��[�~���7�t9�>N"(>7�>��ɾ����H���p B�`l�>03�?^o�?'@g?�݋�4��=J�_�Ӈ0=�R�=��ͽ,[.>K:�>������!?�ȓ>�����§�g"�=��0>a��>�%>B����N��q�K��ξ�e2;�vY%���ξ����񾚚Ǿ��?�S�K����»��#�z֒��<���%7�J�s���4�|�Ͼ�?d��͚?�ݤ?#�>#�Ͻr�m��^]�����f��>-g��n�%��ݝ�"H9�59���?��x���f�-2�=�2��^���?Ӽ��]y��n�|��S��2B>��>�iP?kƾ�X	�N�\�jM����I>�L?�>�vp�fS���M�����?��?�����8��{�E����>��?�t�>���>,aپ!�����>{,e?��u?y�_>�0��ub���䍽l��?��k?�CO?�,����?����h�輇�?�!F?w��>=���"F�k*¾9�*?��?LF8??�`��{��i$��d7?�?{d���q?z��>���>�����ol�S�̆<���>=�<0�������(D����>���<֢m��[����:>Fm���7�YjD�8|��<0��Cc�e?�oӾ (�=��c=s����0�����*yq��㑽�$O?���?�H?2�E?�� �W��:ip��b=,�>�.�>�>,\<�Ej>C�>�c	��]��K߾�?���?�*�?��5?#ke�戹��U}�ޅd�=���d�<n�	=��=A��_�<䡧=,�@��<�)�=��<>^�?>[~K>v�<>^ >��3>J������W������,�f���?��S��;R�^ල0��AL����_g��������彷���ܞ���e<����!):�y/>��>��>&^>�O^��u��i��?����"ž�L��u���R�����Ƴ���ľ���lD澳��<J*�� ?ET�=`�7�bv�>rf��j��'?gR���*>��F>pFL>:#P>�T='b�>�[�><��>q�{>^h9>>�o� ��s��5�I�P�B�j��JU?�R��d��rva��'���"�2>��L?�S�>�d��s���2#�k�#?kۗ�(� �^]D��3>W��>P�?34ؼ�=�]2��H�<���
d�=x?U��>��u=�P�!���m�>q�>����=�֤>T�:?�y�?�0? Z����>�XF>�ɉ>�f�=�b�>)�^>�e>��?m�,?�n?_M�>=}<>�Y#�6`�N� =����b����eƼ�[�s����+�=ӓ>.�g=�B�= �=�5���1=H��=��>(�-?:k�>S�>.Yi�Y82�s�M�i� ���i>��ǽ� �>�>�/�>�!�>�о>�!}>`<%����Ѿ�L�>��t>%vS������ �n >0�>�hn?�D=?��;�/�g�����<܀�>*��>6:?��>��>-}J�W<��ҿ1#�5��U勽p6ۼF� �ɞC�:�T�]iU��{/������<GKd>_�>^ni>ζ:>�d'>m�0>�l�>u�G>:D�=�=����; F���L=k�)�<�X��P������>��+�M����ۍ���uV��0??���>ӷz=c�B�З�ۍj��&��o�>�v�>�_f?2HY?��-���4�l{�x�����;�??6�7?r�>�7�<%m>�N��'D��,�>��Q>(h��>�9����h��I��=�3?�M?�r�>{{:���\�iP�l`ԾEҮ>������ �.,�? YU?c�
�K���'��N��k��5�V�%���|�q�����5�/�L�ﾢ/ �%#뽩�">��>@��?v=F�"ok�����i���Jr�I��|�.>N-�=Ʊ>���=�1q�����<�3��z%�L�=�w�>�IF��<?
l^?�4e?l�?KF]?c?����{?. >
��>��?e?Q��>,c�>���>iSP=����4ͼ�tڽ�^��,~��D?����x="��=�NZ<f<��<��=�q�@��.�*�jv(��ȁ��2ڻm�=�vI=ʙ�=�M?�kI?���=N�=��z=#(��4�=[%�>�s>��s
�1��>/7i>��>��;?1Z�>�]��h.�2�I�\����=��H?�_?*H?���>��S>x��r~ƽ?�>꣯>��ʻ�P���O��Cо�U�<��>���>&k�=-j�>d��?�	?�	�=��<�'��6�X��� �V��R.�wƓ>g�?S�=�ž {�]Y�� n���j�@i�=SQ2�t1>��D>���>]��=:�=��a>�?�6�=�ң�G{����i=|!8>u�>�K1?9��>�?�<'���@�[�3?s�*�X;��~����'�������>a$�>�*>��"?���=�_�������'S��QJ=6��?�A�?++i?T��g��'>Es1>���=�d[�,�����=�U>�=B>�q�>�;���	����"��t��M�A>m���Є�}H����<H俿	�=��聾�lӾ������^I(�;�T�\��������` ���U���d�9۴��"O��� ��zMn�Ƨ:?q�B?`"���껼�!��[����Q�D�>3��s�<c#����=|���㾪	�t��O��ئ��ؾr��>Ӎ��ۤ�7ۆ�;��0>E��=E�X?��ؾ(�߾�VO�������O>�>K�= <{����`�S�?�$?­��ҼR��@'>��>��?tJ?�զ>��ƾA�D�n�>�:q?�"�?;T�>ȓ��>����i����?V:�?�;6?���M5\��<��Z���?/?�{ ?X��zs6�]����4?�/�?G,@?-���'�����z)*?��,?A���y��>�0�>3<8>H���@�̾`Wx�v��G���╝�
�a=���!�C��$��2�����>��1>{
J���ƾ
�>�u����O�/�u�m��=[˾��&?�n���Q8>T�>[�>O�)�s\��S����b�&�I?PR�?��?Z�I?o}#�{軾�5>0ҡ=U�>&>1>�d}>Uy�R-|>d�>��F�s����G�PZ?%2�?w�?��y?ۜ���lο�'���~��S�����=j��=�$%>jN$��G= �<����!�<��>�]�>�V>&7z>p^4>�@+>h>�����^"�c������cR�o�!��<�7˖�W��ߝ����ľ�|�J�.�k��n[��^K�����&L�7�r�Oء=�^�>oS�>��>�P�>Om�>R�P�ņ޾q��ӾK�-���Ⱦ#�˾�����J�sU��q���j��-���	�"^�>Ն�=����2��>��o�-"c<���>t޺(�><�=�w�=v�,>�٥=6��=s >�V>A�)=�Ą>��IQ��	ꉿ0�5���
�% ¼~=?�U_�坸��[M�ƾ��낾���>�;?�E>,��닗�֏=�,��>?����d=�y�2��ŽR�>�0�>���<
l��<��{����~bz>��>�#>�\0�@����_&��V><��>��־S��=��x>�(?��w?�5?�=d��>��^>�+�>ǿ=�8L>5AQ>F�>H?[D8?�00?^@�>�L�=��d�U� =|C=%B��FZ��$�����	�9�w<:$�XCA=�c=�9�;�^=��D=.@��%��;%g=�?Q�E?��>C{�>�\Y��O��J;����h>��"�>Z�?۳?*h�>�Mg>����SS�c�Ҿ�����>w��>cZO�Uy��n˽O׷>�v�>iP?��&?�f�&���B�a=��>���>.5?�g?Ie>��p=�E���	�Φ���WH�������<\�=�_�<4+@�
�$��`�����PB=�½�^>���>��>�_�<���=�1%�X��>��>z�򽰒�<�H�<�f⽐5��=yG =�1{=��=���=���;��y�k��2Z9����;:��<�o,���?��>��>�>=���2g�X���{��>�e�>:7F?��8?�c����!���z��7c�̬��	?��k?�\>3`�+�>�|ܽ��=��>A�>:�>�^M��5վ+n���N,����>5�?��>����d�j�Z�U��L&�>��1=�,_�ȥ�?�'b?�F���5��)�
9�v����N��1��g0���)侗r�d�����J�ھY�ۄ>w��>d��?��_�=�T�Sg��c���k �8�N>Z��=��> ��=����е�������:���=ϝp>XC�>w��k�>e�X?�B?��?W4?m�G?�!�Ҋ?Tt�>bk�>u��>O��>W��>�`�> D�=���<pڽ��3��UA��eľSփ=��>��=Į�>��>�Hͽg2s�9��=�x$=U_��訜<�~�=EO=�;=�O�<�;<��=s�?�S?Py|<?�:��m<�Ҽkw#>��;>���>6d'�7_���>��?�n?��9?8�>EP#�P=��,��Y'�V�4>��>0g7?�)?K�%��Z��':�/*�`yw>��>��<�/���'���Oλs��>���>2�>���>��?��4?�0?| �0�8��P���j~ֽ��潓پ>y��>��>�Υ���*��=z�.{K�&� �Q̽$JP���=:��=0i��">�_>��=�;"=P�!���ؽ&�s��׽՝�>���>'�?E�i>#S6�������-+I?EN������X�5����(�+�]c=�?��>C3/?P�=N���\b��q]O��P�>��?���?�?�{�����=�ة;�0�=�_]����%����P�>�P��|��;�>|�&�%
9�<9z=���>�<�>&�=zVľ���!\.����YL0�"[W��L� ��,�߾�3ʾBY��5���Or�% ݾ�㽤z	��R�����U~�ym��۠��7���i�?�V�?�Z=>žf{1��J������s�>;�5<|�*��	���j�]�A�&���W�� $���*�`�C��о5"e>I�Q����y�������p?>�ws=�a(?cE���ZϾ��;�A�:>J%�>�\>�^��Eߏ��W�������?�??�N�%��N8O= IL>�?��p>�>hN��F�|C�>t}R?Ut?B��	�g���z�(���;�?Qz�?E�K?�p����-�^�9����o?�N1??�>2����	�g���� �>p^?v?+?�;*�gMe���"����>�<?,y�����>?xԱ>\����s�o+�=ܣ��3�<C��=3)C�<�/�ɽ�.���ݭ<"�>	DF>��(�����>40ξ�
=��p������/r�Jվ�O?���δ�>Xn�=�#�3�?�ԅ��=}Y�����5K?�'�?\?��|?���Bz���V�ӏT>Q� ?���>���>q���m>�!�>ڟ�.1���佾�%?d �?Dy@�~�?lm�~�ῳ+���CҾ���<�>��=7p^>�E�Z�y=�',�U��.I��A3>ڏ�>c��>�(�>�>>�@>��5>{����'�^ײ�{䇿��4��.
�8���Ha�A�[:��L��b��Il����m�Jj8��P~�_X�e�"�G�ս��p�e_(>n�j>7E�>=L�>���>��h>-Խ��4�1ɾ�U�/���޾,����'b�����ɰ��	��=:U��ֽe8���?3V�=�ݽ�;�>w�6����;y��>v�[��c>3h�<M�5;ZCT=5�/>�>�PN>P@A>Jo�=�܀>3�&=rދ��]��q��ծ��QQS= �2?:������T5J�g�
�ۥ���|�>h;?�,�>
�)�Su����K��}�>S���tG�N��<�
�G��>���>8ƙ=�/�<&�8�N�)��"����J>�0�>�8>� ����w�ν�n�=^N�>v�վ*?�=��w>�e(?�v?6?C֗=�8�>O�_>��>��=xK>�P>-ш>v�?#�8?��0?�G�>Yp�=OHb���=�E=��A���Y�����Tp���q#���<cf-�7C=|l=K��;�c=�iH=Z8��џ�;#�=c�>�?	}�>iM�>G�価V�I
D�܀>�mΎ>cO��{�=xB�=���>�+�>��?[7?p'O�ҵ��IC��U��>��X>�:��-��xߚ<�>;yj>K�?D@�?�s�<t�g���3����=7��>��>k�)?�\�>}�u>w�K�o7��G�_rN��D�T�[���m=��>ހ��OC?�&>����;�Ic�=k�>|��>���>�5>��$>Ze�=���>��>K�>�{��R�����н}�ݽG�=11d���=X��=���=#���I߽������Ѵ���x�:l�g��t?�^?� �=�d�>C#��de�"A����>9	>�{?�Y@?��P>�"��=z��2[����g
?��s?�?]m���~1>�m��m���p�>�O�>�v��Q=v� =�����䊽��@?�d&?��y>���Z9��8Z���ξ���>�J=���gݏ?d�`?Nv�v[b����}K�q���"�O�꽢N���1ľB�"�\{&�|Ӿ����-j��Y�=��>
S�?}�/��	�=EH澬+��|�����9�=��<���>`1/>��a������Ü�	Y-��K=涜>��<$w�>m�Y?]�V?^�s?�=?#�?��7���?�Ù>^!�>�y&?�:�>�P�>���<E��/�=/ז�����()�(���2$o�q��^L�=�)>r�2>��=��:y��=���;ɔ׽*�>�I��<��+=a2E;�Ba=>�>��#>��>)�*?���벗=l����d�=��*;���\W���¾�9<�	;>���>��!?��l>ڢ���@�����0�<+>7?c�G?<�?�=�����K�l�7��$�=�q >��ǽ��=�6��=�W9`>�e�>BQ>l�>�4�>�o�?6�)?�	�>�}޼�;�Z�o���ﾃG��{���>���>�G>��{�O-$�Y���Yf�X�_�����ƈ���N='��>KE�>�3�=�}���\r>f-��K��������Vh����m=Ƀ�>V�?�t�>u�?>\|׾h���MC?'F����US�����A뽑�J�*�%?���=�'?_ ��M
��Zҫ���0�9%�>�l�?<�?�K?����S��=+C*�d��=���>��G�
@��b8�>dR>�K��?ʵ>�K>8������; 	�>K1�<���^��(���Q>�����'���'��������$�bM�c�6�v㋾��(������>*�-�,�ި������Fݓ�m���% ��N�ľ_�?��?#�>���/��:$���.�k!�>�_���j&�����	j���Ծ���Z���j9-��Q��6��>S<ľ�뎿�҃�%�=�4=�ZG��g1?����`7����6�>ꏪ>�>����b��P��Hۈ�*#�?ұ#?n������G��<펓=�?��?Y8�=�݂�|k���a>��8?u�V?�u�=�/y�����vun�}�?C�?��N?Tf�<�9�� ��"
���?f>*�?��%�x{!�G���:!?K�?r��>��龉����6k�V�>v�s?-Ч�� �>���>嫞>�0��;х��D�=������\��� >J�E��qv�U��O�	���	>d��=>9>0���]R<�
�>�u����O�/�u�m��=[˾��&?�n���Q8>T�>[�>O�)�s\��S����b�&�I?PR�?��?Z�I?o}#�{軾�5>0ҡ=U�>&>1>�d}>Uy�R-|>d�>��F�s����G�PZ?%2�?w�?��y?ۜ���lο�'���~��S�����=j��=�$%>jN$��G= �<����!�<��>�]�>�V>&7z>p^4>�@+>h>�����^"�c������cR�o�!��<�7˖�W��ߝ����ľ�|�J�.�k��n[��^K�����&L�7�r�Oء=�^�>oS�>��>�P�>Om�>R�P�ņ޾q��ӾK�-���Ⱦ#�˾�����J�sU��q���j��-���	�"^�>Ն�=����2��>��o�-"c<���>t޺(�><�=�w�=v�,>�٥=6��=s >�V>A�)=�Ą>��IQ��	ꉿ0�5���
�% ¼~=?�U_�坸��[M�ƾ��낾���>�;?�E>,��닗�֏=�,��>?����d=�y�2��ŽR�>�0�>���<
l��<��{����~bz>��>�#>�\0�@����_&��V><��>��־S��=��x>�(?��w?�5?�=d��>��^>�+�>ǿ=�8L>5AQ>F�>H?[D8?�00?^@�>�L�=��d�U� =|C=%B��FZ��$�����	�9�w<:$�XCA=�c=�9�;�^=��D=.@��%��;%g=�?Q�E?��>C{�>�\Y��O��J;����h>��"�>Z�?۳?*h�>�Mg>����SS�c�Ҿ�����>w��>cZO�Uy��n˽O׷>�v�>iP?��&?�f�&���B�a=��>���>.5?�g?Ie>��p=�E���	�Φ���WH�������<\�=�_�<4+@�
�$��`�����PB=�½�^>���>��>�_�<���=�1%�X��>��>z�򽰒�<�H�<�f⽐5��=yG =�1{=��=���=���;��y�k��2Z9����;:��<�o,���?��>��>�>=���2g�X���{��>�e�>:7F?��8?�c����!���z��7c�̬��	?��k?�\>3`�+�>�|ܽ��=��>A�>:�>�^M��5վ+n���N,����>5�?��>����d�j�Z�U��L&�>��1=�,_�ȥ�?�'b?�F���5��)�
9�v����N��1��g0���)侗r�d�����J�ھY�ۄ>w��>d��?��_�=�T�Sg��c���k �8�N>Z��=��> ��=����е�������:���=ϝp>XC�>w��k�>e�X?�B?��?W4?m�G?�!�Ҋ?Tt�>bk�>u��>O��>W��>�`�> D�=���<pڽ��3��UA��eľSփ=��>��=Į�>��>�Hͽg2s�9��=�x$=U_��訜<�~�=EO=�;=�O�<�;<��=s�?�S?Py|<?�:��m<�Ҽkw#>��;>���>6d'�7_���>��?�n?��9?8�>EP#�P=��,��Y'�V�4>��>0g7?�)?K�%��Z��':�/*�`yw>��>��<�/���'���Oλs��>���>2�>���>��?��4?�0?| �0�8��P���j~ֽ��潓پ>y��>��>�Υ���*��=z�.{K�&� �Q̽$JP���=:��=0i��">�_>��=�;"=P�!���ؽ&�s��׽՝�>���>'�?E�i>#S6�������-+I?EN������X�5����(�+�]c=�?��>C3/?P�=N���\b��q]O��P�>��?���?�?�{�����=�ة;�0�=�_]����%����P�>�P��|��;�>|�&�%
9�<9z=���>�<�>&�=zVľ���!\.����YL0�"[W��L� ��,�߾�3ʾBY��5���Or�% ݾ�㽤z	��R�����U~�ym��۠��7���i�?�V�?�Z=>žf{1��J������s�>;�5<|�*��	���j�]�A�&���W�� $���*�`�C��о5"e>I�Q����y�������p?>�ws=�a(?cE���ZϾ��;�A�:>J%�>�\>�^��Eߏ��W�������?�??�N�%��N8O= IL>�?��p>�>hN��F�|C�>t}R?Ut?B��	�g���z�(���;�?Qz�?E�K?�p����-�^�9����o?�N1??�>2����	�g���� �>p^?v?+?�;*�gMe���"����>�<?,y�����>?xԱ>\����s�o+�=ܣ��3�<C��=3)C�<�/�ɽ�.���ݭ<"�>	DF>��(���5p�>C�꾱�p��}B�N+��u�w�W�j?���o�=��>�
�=��<�j��'Zm�@��� #a?���?��h?��P?�$8���B�)���+��>�LD?��= ����Z���y>��>�䋾^���U�;z�?���?�8�?R�o?�*u���ܿ9���Ҙ��#����G�=P >WK>T�"�-�=V��=%�=��<�>"=�>'�>i�>�v{>nE>�>���2%������皿�03��@��p��a�Y���Nq��K���ﭾ���n�:��g}�~�y����:�սbΘ���|��$�=@�B>�}>��>Q��>]t`>�̾^�!�`���꾫$��M�s���CǴ� �v�P���ØѾ� �I?�@�I��>U8>�O3=w� ?��}<L�e>\��>g=�>ٯP>�W:>�~>�q�>�Ȱ>LJ>u�>�Ĵ<۠>�Z�����bW��p;7�C����!��H<?T����D��TL�+7��p��I�>��0?���>_-��!���N���>y�X=��὾4���q����>M��>*�l=���~AG�z����e��]`>W�>�TL>UL:�q<��[h��}y�>;��>;G����>��7>4r?`�l?�K?�Q�Ɗt=lʽ>��1>���>�sC>j��>4k>�+�>3B.?��<?�|�>�0�=;{D�LI�=��b�������[=n�:�1�_�ٯx�%E?>�c��$>�(i=V�&<D��<�Pn���:ܼv�>��?eP?О�> џ>�jy�cm"���N�yJ�<�Ճ>�;0_s>:�?;?UA�>��>V�>�c3n�����N���>�;J>��?��L��@�R�T��>q�+>�4i?��?	�Y��r޾��X�)l>��? �N?��5?�>�>����e��FҿR�o��_���Yi�G8�O��1ӽ���<c����U߽�k�<�[>Sz�>>܄>>cf>	�z>��_>�@�>ڰT>��<�H�=�[�<x>�a���=$
�=���=�2̽�o�<3m８5k�E���[$�W����B���_�>M>?���=��&>?:��%Y)�&F�� �=�J?/�>�Q�>EVe����Tw���e��E�4�?���?P�?��H��+==��xi>�I�>x�|>j÷>t��=ÑA���	��)i>��=?��7?�[�>�"��P1��L�cE ����>��^=P�<O(i?��3?@��/'0�$K#��h��\�?L��;�¥��)� 8D�n�;�:K���� ��">��>o��?��A��=�(���_��<ח���p>`,R>�>��F��Tl�����kD<�����n�=��>�v�>g��m�5=of?��E?z�l?���>�|l?[��#�>� �>>�0?��0?�s ?�ƌ>�,n>�E=>2�`>��=L�m�ݽ����%�=��Z���>�Q0>(�j>R�/<N��iW���b��`r�_<v��"�<< <a��;��U=%I>^��=$:
?PFN?]5�������ؓ�(��о����=��?}ą>v�;�U8��O�>/s�>�@,?��>��i���ӾY��k�	9>���>��9?�&?�]����<��a�H��:C>���>��v�b���0�w�(��ݼ�n��>9�G>��^==4>s?��?D}h?�����F���L�����{[>���>�u?e�	?�es>��$��j�%$r�|))��m ��Yb>����0�P=��<�ά=�r=f�=�>�U�=��ڽ����Me;wu	>���>�ְ>�>%�<�f�9��徇;��Jj?C��PB���	��N�O9�=�� =2}�>�����>�{S�i�w�Ow��E���,?���?�S�?��J?��0X�4�=]O>}��<��ֽ E��!t�;DZ��J�>B�S�H������M�>Z?��?eoh=��$���M�P��=0�Ϳ�.K�-U������ ��?Ҿ����5/=�����9�&���aZ=���g��z�����;��@�yZ!�{;z�ξ�S�?�D�?����wD�M��W�0����>j?�7q��>ɾ�о�싾�͕�ܹ��oΙ�׳��>7�P�W�s\��{�>�pJ��u��fMj�V�:���y�4x�> Kq?����������#�3A>4�'>i���I��Lן��į��h?� ?����+x~�V�#<)���^�>�	�>S��=������=�V�>��?��*?���Cz��Et����m��i�?+��?�/N?�>�� �<�].��=̾�`+?��?�Ȩ>p����������]��>%9?ݴ*?�d:���V��Y$����>ۥn?kf|����>���>@t�>O�X�;���	�=�մ�ο�=��>w��=�C�=R����lվ:S5�EjY>��y>G�
�������>R,��M��|s��fs�D�=�|�5�3?�z�v�U>��>�l=����0q��p��-4���^w?S�?�+�?m#7?*Y� P���l�&{�>���>�>Z������c�>$n>���;h��FϾ�j+?D"�?	��?_�X?�U��ѿ.���)ǭ�<ު�|�>L�=�<>A�
�Ǜ=�'=|2��A�0=@><G�>�j>=g�>ӬX>��;>�m2>�p��H�%�0s���b���[6�j��_�	��4Z���3ㆾ���K��Q��m����?��t,-�P�0��9���u��g����R>_΢><�>�n�>i�>r-�=͓�`'$�;��=�-�$���f��L��@w�������Œ��o־�ڽ�i﾿?1?�=��$�߽�(?������=�:�>�xq�I	
>MkH>�=��;�[->4�=r�>܀%>��"=�+b>{E��$͎�V{}��.�z8i�Y'�= KA?&���׷�
�@����,�����>!�?�0>�!��Ԟ�7X��>�K�<5���]Ƚx�n�s�y>��>{|<'�J<{����7���/�ඟ>�Ϧ>M��=0!�c���' �b
b> O�>CҾ��q>Jԩ>�5?ܯt?u�2?ϰU�0?�_y>�۝>全>�_�>i<{>Nw�=�	?�k?�_%?���>��Y>�靾�f���ښ�q�/� �<�z��ѝ�d��#B3<�CT��3>z�%>*�=�Ս�Y��N	�=p�=�p���G�>��7?���>E��>)���s�9�� T�۽�;
�.>�J�"��>5��>�	?n�>?S�>�z_>Mʽ&r����a�>K�>�=���>�[���<(=[��>�u?��C?a��=��x�~��j�!>,��>��??=5?ذ�>곧=�@ ��E���׿��.��"0�:�h< �+=�/J=�xb�ԴE��Խ@F����ͽ1[�<.À>�/�>5�>A4T>&.>�8�=���>�a~>�.���8�= M���	�����;��=��a���*��i�1H�id���/�c	�~H��^�ȩ7��i�@?+P�>�e>���>B�ξ����u�_c�>T�.>,uU?�E�>�8�<�^ ���n��fJ�Q�˾V,*?�g?�m�>��e��8>��Ȍ�GV_>[k�>�m�<n a��-v���i��=3��>��?���>�(�g�`��)f��\��> �a=~T ���?��O?'���F1�
�.��S���
�)C�0��~�T�ʾ�+���!���9����8��F=Q��>���?>�L���=+���z���]r�nl���z�<��<��>Ӛ�=F������ؓ�6揾,~�� ��=~ڕ>�N���?�eI?CR'?�U�?�	?am?��7�(?�6{<K��>��p?�'?@4?4C*>�4�>�ƽH��j{����>��|}�H�H�*rڼ��>5/>��T=C�m���p��&;�e���E����Ƚ��w�f��=B�<��A�̼�t�=
��>��7?ʵƼ������� TQ�# �= H>���=�*j��ݽWp��K�>�=�>�4?���>M�ʽ/���U#�/).�hN�>Ѵ�>ЛU?��4?T��d>���?b��w�>9k�>ǽA�h��0�+O�Mzμ�I�>W§>% �=�<�>(>l?u-?^�>C�����Yej��������4�ӽ�q?�Â>��>�$;��)���EW��y�M�G!s=����I>	��=�i��oK>�"o=u�G>hb�>=�-�&mþZF��Lc��Z?���>�?��>O��C��5�D�ՕQ?��=qܾ]ȿ�����2A��f�= ��>VH>]_?BnS�����7����+�>��>��?��?��A?;��<5�R=z��<�^@>-�Q>h�4��sX�as>�$e�"��>��>0��<x8�V�=/��>3�>���<!ᆾ}��->��ӿ��G�5ɾ㿾��l����c_��_���.��\����3��
��d��=�w��
�d\�����F�ľ�}��S�?
z�?�i{�g�>��C��gZ�Hw:�Zt�>�'�������х�7���ԕ��ƣ��{ܾu���9��BV�
�t�>��b������N�l:�8{��Ve>�N?/�E���a���_<�Ns=�~O;c��Tj����������M?f@?���F�����V�'>�
>?+0�<%�4>�gz���<���>��4?�?�!�S���}�T�mI>��?���?ZF?�Z��ю@�;�*��-��@?�?�v�>��|����<o���0�>N�T?H�'?�C?�4]��.��T�>��n?$y���^�>k�?=6�>°b��䨾��g=��Ѿ�Z<2�>ST��K��B�W↾�yJ��T>#p>c+����ƾ5�?��6^�(WO�%��0��=Dʽ��:?Ҵ�Ҳ�>7%�>�c>D��}$��*��x���!�{?4ؽ?��y?�1?<U9�?���MZ�;=t�>O�p>Y��>��E�-C�c�>��v>�嬾�s�����Q?M7�?���?gn?kI�xտ�=��w����~����L>m_E>�U>�Ht���=���= ��bJ3=�j)>�G�>ۧ�>��~>v6�>/S>�,>Qp���)�~���旿?�&�Y��vd��!^��a��GȽ�#��ʾ�w�l��=�>�R����wԽIR����@�v�0>��>�v>'?��>��>�2�&�	�:q��bI���>�S����}���)��������s��|��:��Ae?�J�>t����?�)��.�F��>H*<�Ϟ>7M�>~v�<]��==�=�v�=��>���>�o>E��>`9�=�+���R�rNK���m���<�J?�E����9dH���⾑���
?�x(?Zs�=i.�Ӷ��BNy����>y]>H4����ѽ���C>{?�d>{Ί�0�V������ڽ��>�(�>��=She�J\о���;='�>��о=a�=B�|>�O&?ݫ|?ge2?��9=D�>[�J>��>��=@(,>�X=>��>��?56?#�,?�z�>���=oS�ٲp=�f=3YK���`���ǽ:�ȼ_tU�>�;f�:����</Q=�38�G<=W`_=�Z�[}c<�7�=G�?��I?���><2>C���d�v�b��c>C]0>'��=�?!�%?f�5?���>uA�=�;��Q뾽پ�>���E�>��y>N�Z��錿$�=���>a�>AEK?�PD?�R�8��pk7<S��>ǡ?�(?$H?�K>�&&=m����`�lտDz.��S�V��>N�>K|�:v[ʾt�>�P>[F�>l���O>���>\��>o�D>�G>ڍ�>gG�>ۻ�>
�d>�
�a{>`���3+��cº/N.>���#�ыH=������ֽ3 ���1
�.�;Weֽ]���BP�;��>-�!?�ذ>F�#=�ɾ��߾�T�D��>U�+>Q��>!�> ��?�B��G��׺��� ���?��?wL�>�$
�t�̼*�<�}T>�R�>l�Z>�e�=�k"���������]5>0��>�%?�YE>��X���|�0�x����\S>Cn�=8r�<���?Hׁ?���G������F^@���2�2��3t=g#[�5g��%#J�i�P��
� �����a�>ۗ�>�8�?�-�:��н���r���H��j�/=w��>��=���>��m��=��0����	`�S�;+�(>���>��<�&�>�&n?�~'?�.?kȕ>/\_?.� ��M\?>��>[�>EH?�D?Ғ�>��=yg0>>��=bQ0���4����9�=��<��\=窦>_>6)�� ���=��
;T���U������<��T=�=�R*�#�=�!>"?��:?٫��`cݾZ�0�O��{�>M��=�}�>aUѽ�H����=ɇ�>�;?��0?��>�M��T������I]4>��?7� ?U)?��O��9�>4�� �W���>%�>P\�=���NA�����ѽ���>�o>�!f;��r>TNn?��L?]R?���XE;��5W�wa��ĥ���	�>�k�>�`>!0�i ;��_��M�a�^{����������;��1��f>�U>�R�>��>��x=�� �9�F�y��<+#6>/x?<��>�i�>��=CR��࠱����!4P?����L̾������པA>����/"�>���{�>�@�%À�p����*����>S�?	�?H?T?�ӼrA��8a�>�_>~x���I����R�i�'ѫ<ѽ\>���ٓ���	���u=�
?��:?���<���p'�Y�5=����Y\<��7�� ���Zrؾ�徂���s5;�7��å�|(��v��jЇ�1u�<�ʽ>7g���Q����>>��)#�?�?�?]r��+=�6hL���������><n[�%����Ɣ��J�\!о�-��U�����)��r���b?��,�\L�>���:ߜ��au�C'^� ���S>Q�m?,���f�n���*=�=o:�<��	��'����������>??�8?�[	�9�.�t���=��>�Q?��%>K�t>�mþ��b>��?��9?��1?��%��ř�`][��3>k1�?���?5ZC?&O��o?�@���	?�ٔ?��?4=�>���Kܾ�*F��"�>/�;?�G�>d
׾�`x�#|����>��]?�2e�{��>�b�>�T�>Ӽ�'����ޙ�C���|�����->>)���ֽj�G���Y�(ru=-�>��h>��;�@��5�?��6^�(WO�%��0��=Dʽ��:?Ҵ�Ҳ�>7%�>�c>D��}$��*��x���!�{?4ؽ?��y?�1?<U9�?���MZ�;=t�>O�p>Y��>��E�-C�c�>��v>�嬾�s�����Q?M7�?���?gn?kI�xտ�=��w����~����L>m_E>�U>�Ht���=���= ��bJ3=�j)>�G�>ۧ�>��~>v6�>/S>�,>Qp���)�~���旿?�&�Y��vd��!^��a��GȽ�#��ʾ�w�l��=�>�R����wԽIR����@�v�0>��>�v>'?��>��>�2�&�	�:q��bI���>�S����}���)��������s��|��:��Ae?�J�>t����?�)��.�F��>H*<�Ϟ>7M�>~v�<]��==�=�v�=��>���>�o>E��>`9�=�+���R�rNK���m���<�J?�E����9dH���⾑���
?�x(?Zs�=i.�Ӷ��BNy����>y]>H4����ѽ���C>{?�d>{Ί�0�V������ڽ��>�(�>��=She�J\о���;='�>��о=a�=B�|>�O&?ݫ|?ge2?��9=D�>[�J>��>��=@(,>�X=>��>��?56?#�,?�z�>���=oS�ٲp=�f=3YK���`���ǽ:�ȼ_tU�>�;f�:����</Q=�38�G<=W`_=�Z�[}c<�7�=G�?��I?���><2>C���d�v�b��c>C]0>'��=�?!�%?f�5?���>uA�=�;��Q뾽پ�>���E�>��y>N�Z��錿$�=���>a�>AEK?�PD?�R�8��pk7<S��>ǡ?�(?$H?�K>�&&=m����`�lտDz.��S�V��>N�>K|�:v[ʾt�>�P>[F�>l���O>���>\��>o�D>�G>ڍ�>gG�>ۻ�>
�d>�
�a{>`���3+��cº/N.>���#�ыH=������ֽ3 ���1
�.�;Weֽ]���BP�;��>-�!?�ذ>F�#=�ɾ��߾�T�D��>U�+>Q��>!�> ��?�B��G��׺��� ���?��?wL�>�$
�t�̼*�<�}T>�R�>l�Z>�e�=�k"���������]5>0��>�%?�YE>��X���|�0�x����\S>Cn�=8r�<���?Hׁ?���G������F^@���2�2��3t=g#[�5g��%#J�i�P��
� �����a�>ۗ�>�8�?�-�:��н���r���H��j�/=w��>��=���>��m��=��0����	`�S�;+�(>���>��<�&�>�&n?�~'?�.?kȕ>/\_?.� ��M\?>��>[�>EH?�D?Ғ�>��=yg0>>��=bQ0���4����9�=��<��\=窦>_>6)�� ���=��
;T���U������<��T=�=�R*�#�=�!>"?��:?٫��`cݾZ�0�O��{�>M��=�}�>aUѽ�H����=ɇ�>�;?��0?��>�M��T������I]4>��?7� ?U)?��O��9�>4�� �W���>%�>P\�=���NA�����ѽ���>�o>�!f;��r>TNn?��L?]R?���XE;��5W�wa��ĥ���	�>�k�>�`>!0�i ;��_��M�a�^{����������;��1��f>�U>�R�>��>��x=�� �9�F�y��<+#6>/x?<��>�i�>��=CR��࠱����!4P?����L̾������པA>����/"�>���{�>�@�%À�p����*����>S�?	�?H?T?�ӼrA��8a�>�_>~x���I����R�i�'ѫ<ѽ\>���ٓ���	���u=�
?��:?���<���p'�Y�5=����Y\<��7�� ���Zrؾ�徂���s5;�7��å�|(��v��jЇ�1u�<�ʽ>7g���Q����>>��)#�?�?�?]r��+=�6hL���������><n[�%����Ɣ��J�\!о�-��U�����)��r���b?��,�\L�>���:ߜ��au�C'^� ���S>Q�m?,���f�n���*=�=o:�<��	��'����������>??�8?�[	�9�.�t���=��>�Q?��%>K�t>�mþ��b>��?��9?��1?��%��ř�`][��3>k1�?���?5ZC?&O��o?�@���	?�ٔ?��?4=�>���Kܾ�*F��"�>/�;?�G�>d
׾�`x�#|����>��]?�2e�{��>�b�>�T�>Ӽ�'����ޙ�C���|�����->>)���ֽj�G���Y�(ru=-�>��h>��;�@��5�?��6^�(WO�%��0��=Dʽ��:?Ҵ�Ҳ�>7%�>�c>D��}$��*��x���!�{?4ؽ?��y?�1?<U9�?���MZ�;=t�>O�p>Y��>��E�-C�c�>��v>�嬾�s�����Q?M7�?���?gn?kI�xտ�=��w����~����L>m_E>�U>�Ht���=���= ��bJ3=�j)>�G�>ۧ�>��~>v6�>/S>�,>Qp���)�~���旿?�&�Y��vd��!^��a��GȽ�#��ʾ�w�l��=�>�R����wԽIR����@�v�0>��>�v>'?��>��>�2�&�	�:q��bI���>�S����}���)��������s��|��:��Ae?�J�>t����?�)��.�F��>H*<�Ϟ>7M�>~v�<]��==�=�v�=��>���>�o>E��>`9�=�+���R�rNK���m���<�J?�E����9dH���⾑���
?�x(?Zs�=i.�Ӷ��BNy����>y]>H4����ѽ���C>{?�d>{Ί�0�V������ڽ��>�(�>��=She�J\о���;='�>��о=a�=B�|>�O&?ݫ|?ge2?��9=D�>[�J>��>��=@(,>�X=>��>��?56?#�,?�z�>���=oS�ٲp=�f=3YK���`���ǽ:�ȼ_tU�>�;f�:����</Q=�38�G<=W`_=�Z�[}c<�7�=G�?��I?���><2>C���d�v�b��c>C]0>'��=�?!�%?f�5?���>uA�=�;��Q뾽پ�>���E�>��y>N�Z��錿$�=���>a�>AEK?�PD?�R�8��pk7<S��>ǡ?�(?$H?�K>�&&=m����`�lտDz.��S�V��>N�>K|�:v[ʾt�>�P>[F�>l���O>���>\��>o�D>�G>ڍ�>gG�>ۻ�>
�d>�
�a{>`���3+��cº/N.>���#�ыH=������ֽ3 ���1
�.�;Weֽ]���BP�;��>-�!?�ذ>F�#=�ɾ��߾�T�D��>U�+>Q��>!�> ��?�B��G��׺��� ���?��?wL�>�$
�t�̼*�<�}T>�R�>l�Z>�e�=�k"���������]5>0��>�%?�YE>��X���|�0�x����\S>Cn�=8r�<���?Hׁ?���G������F^@���2�2��3t=g#[�5g��%#J�i�P��
� �����a�>ۗ�>�8�?�-�:��н���r���H��j�/=w��>��=���>��m��=��0����	`�S�;+�(>���>��<�&�>�&n?�~'?�.?kȕ>/\_?.� ��M\?>��>[�>EH?�D?Ғ�>��=yg0>>��=bQ0���4����9�=��<��\=窦>_>6)�� ���=��
;T���U������<��T=�=�R*�#�=�!>"?��:?٫��`cݾZ�0�O��{�>M��=�}�>aUѽ�H����=ɇ�>�;?��0?��>�M��T������I]4>��?7� ?U)?��O��9�>4�� �W���>%�>P\�=���NA�����ѽ���>�o>�!f;��r>TNn?��L?]R?���XE;��5W�wa��ĥ���	�>�k�>�`>!0�i ;��_��M�a�^{����������;��1��f>�U>�R�>��>��x=�� �9�F�y��<+#6>/x?<��>�i�>��=CR��࠱����!4P?����L̾������པA>����/"�>���{�>�@�%À�p����*����>S�?	�?H?T?�ӼrA��8a�>�_>~x���I����R�i�'ѫ<ѽ\>���ٓ���	���u=�
?��:?���<���p'�Y�5=����Y\<��7�� ���Zrؾ�徂���s5;�7��å�|(��v��jЇ�1u�<�ʽ>7g���Q����>>��)#�?�?�?]r��+=�6hL���������><n[�%����Ɣ��J�\!о�-��U�����)��r���b?��,�\L�>���:ߜ��au�C'^� ���S>Q�m?,���f�n���*=�=o:�<��	��'����������>??�8?�[	�9�.�t���=��>�Q?��%>K�t>�mþ��b>��?��9?��1?��%��ř�`][��3>k1�?���?5ZC?&O��o?�@���	?�ٔ?��?4=�>���Kܾ�*F��"�>/�;?�G�>d
׾�`x�#|����>��]?�2e�{��>�b�>�T�>Ӽ�'����ޙ�C���|�����->>)���ֽj�G���Y�(ru=-�>��h>��;�@���f�>�u�%����R��\
�L��??�'?R$��'>�&>Q��>���BV���h�� j��8Z?���?�E�?h3+?��־�ﾾʁ��t5>>`�>u_S�8��=R�F��ߞ>#?��Ͼ�����9���S?"�?�	@`�?Pԅ�6ֿ�+��w��۾}8�=��>~�=�&�����=��ݽ�m=V�<L>>��>u�>=Ʌ>4�M>O�<>(�=%d��xR%�]���v���4�i��A#�	kƾ�����t�(�ھ��.�_:��Ǻ��Ͻ�n�/�%�	=��b�E��E>�9�>U|> >�v>H$!>/U�=�f�˫���;X�I�?P;���@�|��>{�?��)N5������3�r*��G?�C���u?!?�d��e�>T��>�=>C�>[�>�+>6��>fK;>���=SJQ>F`>���=�k�>�.>�K��J��hQ4��]��6�;�N?���� ���'�3���Ѿ+Є����>�y?b>~$��Ζ�����D#�>��!x�#K$�K2,=���>N*�>��>c%3=��A��%M� �ؽ���=l�>-�>�`<��G��ec��F�=���>`�վ�;�=BO}>�z)?��x?O�3?`��=`�>�\>�f�>���=�lP>�RT>���>X�?zP8?͟.?ͤ�>��=��_���$=�0^=$;�k�[�$��J�8@�<�'!��AY=Nm=�1�;��W=�7=�Ԥ��!�;�}�<)�?��Z?�v�>O!�>%�ɾ�G��#g%�X�ɽ��G>��L>d~>���>��?{-?P��>�c�=�$��b�2��&*�LC�>�m�>I)���ְ����=�>���=��a?��j?zN�g�V�)u>��<=�=?��<?3GA?v��>;��=�Sվ��A�ؿ���� ��t=����z�B��8"���"�W��(A�0=��=2��>0�>Tm�>�\>>��>!�=�;�>Wi>����D>	���7���EE>��=��;���=O@�9���X��@��"�A�m�<�b��<�SX<-?m�?Q��;������m���	�J�˾��>1�>�R�>g��>��/=��FT\�r;J��=����>%__?�P�>�M�7)
>+k���E��X�>C��>���=���;���� ��k�<�m�>>6?;4�>0�;��qZ���p���э> >�����?�S?2���s�K?A�N�ҍ"���;�����䏾.��{4���?����ݛ��5�gi���ʪ>g��?ܢD��=5[�3˻�����_���>��"����>���=�?��p���#��	����Q��>�>p4_>}Qռf?:�V?!ˊ?�3E?D�>�8�=��c?7�Z��<0?��/?��9?
�@?�?�m�>
E>o���y���F���5�=���=$im=|w�<�)v=�͌�i��� ==�<���4�d���z�!���?:K\J=^�=�k�=��?¶D?>�+��\��~�
>��>��={'�>�h�>�^��;ړ���>���>%�1?��E?C�>sU=-��������s����?�D?��?�*O>�A=�����d�����>�%>�!���D��}���6ܽ�z�>���>J:�>0�>�r�?o�|?�?F����Ie��m��^�F� ���(]3���ݽ���'���K/���������U���6���^=�J�����<�N=�*�>��U�+�����>h�`=����<*.��ݼӞ?)��>]��>�k�<�"�.�����'X?\���^O�T��MD��)�=��>'�>{9��s�?Cn���A��ߓ��S�_���?�A�?���?\Ji?�^>D����7>v��>��i>���<�������y�����>*>k�dK������y�7�=�޽�NG�9�,j^�l+j�l䲿��I�J}��:����ľmW�1|Q��Oc����ܽ��Ҿ�n���ls���7�: \��{$�����5��r����V�?'��?�s�>��#��r"�	�#�c@�n��>W�þaR��	��xn��F���m��:!��1�1 A�טL�Q���IYs>!㥽0���dt��A�m��X��>`�Z?����N���Z�=�^Ŗ����=�$����!�4Ϥ�L+��7y���+�?u|?��l���v��I����%<�Y?}XX?h��>�Y�����>f�[?'%G?�Gs�.'Z�l�����x<��?�5�?o�??�O���A��2�T��`>?r�?���>���̾���L?C:?Լ>����W���)�y��>?�[?�N���a>9��>Q��>�n�x4��E'�c���ц�n�9>�Z
�����g���>��=D�>�y>^z\�F���bu�>&�`��O_��E�{�;T�i����?L|�'3�>)��=u>�?�L�����������^?���?#�i?kB?=M��;.&����W5>�%?�@�>�G�]�Q���7>�?k�վ�#}��f���?���?��@@`?�+j��Mٿ.8���x���u���!�=�s�=wA
>�f޼�ސ=)�<��m9���M>Q�>�Y>)R@>�4Z>�~D>�}Q>���%������Ð��.�����v���@��K��$gt����1d���c���ވ�{��5y�"r��u!�� �>�}�X>'Dx>u�>�?7M�>cs?>���j� ��kϽ)����e�- S�.5��~̾��*=盀��\辫/�m{�<���>�I��dzG>�Ӽ>[UI=�2�>,��>��^>��>�K?	ּ>��>���>�C>��r>"�>��=6��>���>p̀�y����<�vQ=���>p�\?,CU�=���FM�������bE�>��?-Ʊ=��N�g�����p�4�>_8�=�������z����>\h�>�I�<�y=m>V7��M���1�=w��> 5>a>q�ٽ�����Ҁ��D�>������>�;�>�?�oe?��8?F��=7؛>���>�=N>C �=��>>g3�=�!�>2�?l5?o�?{��>��/>3(��
yI>��>�3��0o(��7��׬=��ֽ���3$%���=nm*>kѸ=#�=��R�3���m�?��h�=��?>bG?k��>m�1>����X�H�\�1���>!�=իD���$?�o?���>��>qx>�����j��-��/o�>��>Qٕ����i�����>�
�>��R?��Y?k����TB�ב[>s��>��-?��!?c�1?�c>:�4=s�6��2���1տP�?���پ���<����/�!����Ѐ�~����>۵�=��5>��>q�3>�q=F)>!J>�;>2��>x8>��뽍$ =�v<��<���DS=T�=�һn�2�"�S<��=���/.}��9<��p��g��:/���?c+?���>I{>����t=�J�U�'��>�D�>
$�>��
������b�]����R��� ?)<�?2�*?�\��<�����6=\��=�Ӫ��_d>��>*��f�<�7��=�F�篼>�wQ?�Vk>����cH������6��C�>��/>'��Yr�?���?���7� �g!�����:/�B+˽=�K���n�h�ɾO�)�/�)�v��奛��N6�|g)>�>|[�?gѽO9����|��e��g����@��fW>ؐ���4?���<�S�T��,�۾�>��o�*�6�>�3�>���=�b�=�w4?K�?�z|?���>%W>����@}?���KF�>7r?�5?��2?��>A�c��<sE���;߾���rO����=���=p���+�>��[>���� v�1�=9�>=rD���l�����^I�q��<��=�z>�">�@?�SN?�W��T��Y��>ʐ1�dK(�T��>�y�>��C��c,���>{?Ek5?�(?�->qg[����FS�s���zӽ�{"?�oH?s�?�	�%_��w��'����� k>K�g=&�!�� ������_�<h>�'�>>�>p݊>W�W?��m?|�K?ޢ6�7�7�!^���8�S晾i[Z�ϐ˽���>h�4>���+Ji��!y��mc�<�tw$>9/[�b�ڻ��'>�*=-,�>�P<�\�=ܾ�>��]�1�T���տ�=��>�8�>�h�>%B���L���������$[??�Ͻ�+:�����)�K��>滺>*�j�;#þ��w?�覽T����B����H�g�5?.X�?oy�?�^3?�s>�u=����=A߿>h��> =�w���y����-���=*��;Z;̾�;�(B\=�>�)�=X=?��:"�b���19������}A�R������i�ƾC�Ծ����er�mk���]F�1f��_Q���O�M��g<��L�꓾.�����7��A�?��?�6�:���L�ߍ�4��m�>�ѵ��A�yѾ��������!̾�d}��[�*�;�x�"�O,���@�>�q��j���������H��ｲ�>f�6?����>$�*>'��N�<�2U=L ��25Ծ�������P\�B�i?Y>?�=��=�f�=�0>�N�>�Q7�1�(>o3��]0�=�Y>�5?)��>�h��U��������=��?���?�C?�%�yZ=�yc���ρ?��?}��>��w��;f7���?6�<?���>h����T��}j$�Ej�>��R?Ӝ?�k�c>��>:��>?ﺽ� �J9��s����d(<FH?>=���S{5���P����6�=
o�>僈>�����Tվ�X�>�������;o���X�>|��>�k�>[��ڳ<���>�]�>�b���������Ľ��K? ��?#S}?�/?[�)A��O_�<]\Y>���=�8P=��>�t��ы>��>����B��3<H�T�B?{�?vz�?�r?��߿����?���SЄ�R�>D�=J>�A�=)�4>}��=��ƽ�ݍ�v.$>��>-��>�_>~->�[3>+�Y>�����@�����8n���]?��Y�����������͆�H��Ѿ[S��@���q~���P��$��������!p�A�-<
_�>E�>L��>���=x1=��ڽ_����ɾN;O=�T� �q���	�����L=��U=6�����P��P��?��J#[<���>+��vR>��g>t.L>�x?>��>� >��}>��=S��=Z��=Z��=9��<�f5>Ct;>ھ��I����O�Q8�+nD>2}A?	�ѽiIj�v�H�"�ƾ�-㽂��>l�%?��r>@�%�Z����Պ����>x�=߳O�8g�����br�>[�>��=@��=6>�90��P4�\NT>��>>{�>_.�=�LQ��	���>��>X����	�=��>nz?�1o?��/?�o>�T�>V��>��u>"�=O{!>{�
>AZ>�
?ft/?_�'?'r�>m�=ܣ���t�=g�=�e��B���S�ս��n��rԽ,F<==ʜ���]=�Ě=��=?=��<��I�᤽��=��?	�R?�8�>�%�>J7}�A�@���;��0s>�<>>"��?���>\�?�4�>}�>i����־���`�/���>�E�>]��9R�� ��<o"?O�>%�D?��G?�0��/S����.<s�>�2?��W?I�??���>�-�<�ꦾ�M�\�����7�4<���gw����e�X<s =�.L�����W=��Z>�%�>.y>^KC>��=k�V>�>�>��>gxҼ���i��j�|�#��=��}�~���O��ŕ��N?=����༽eS����O���]�����ai�����>}$ ?��h>�Q>duc�Kr�$w!��c>V1�>[�>.x�>d2*����?��|>��B���
?��V?��>�5�0��=~<^=$��=�)>�T>H��>�d�=7@����u��V>��>�y?�nj>�U��Yc��K�ˡ����>Ma=~�{��U�?�5r?����h��<���F7�)�'��_N��t��
ʲ��HܾUz��A�=�;��ƾ�<9���{=���>T̫?	�e)A=��G�5����=��>�ھj�>��0����>en�=5|��@��]վP���<�}>[>?>^`c>�̎>Y�?Um?~~�?8^-?.!�>�6ľ��:?>��>�-?.w=?I�S?�ga?�;L?�u>���<�N�|����Q�v����>F>�>�M�=���<|o��a�=�g�=��p=�b�<ŭ6=@���gS���Yʁ=��.=+a>,�5>��'?�7@?�&�vT��ɬ�=�{*>�6>׳�=`��>&]6>�c����<tx�>��??�V?�d�>Jâ;�+���!�
��Nj���(�>n??#?ꄺ�%j�<0
N��Ծ���=6۽>�Y�=Y:������д˾�m�R�>�>��+>u�X>�[?b�_?]!E?�gԽ��D�?5� ~!��6�����79�>Om>�J>�˾ML��ى��Nd�k4)��>>�8�K
7=�#=��>
�^>:�=]>H�>^p'���t�#{S�����`/�>h�?}E�><�H=ׂ��оN���&�)?�΂�����!
�C���
����p�-�_о�y>�O�<v�j��Rb�m�e>���?��?��?Xm��d����G>��>���><&������/���"7:���>=�@>�*���.��*L>��~>`�=��3��¾����	%���ſA�`��>����!����aԾm,?��箽�L����1�&�뾯 n�Q�|�#b����F1W����2ž&û�2��?X�?B�V��D���S��%�y<}�c�� ԾU�<��j���1�����%��:���&��U�'�G�<���0�t+>(Qd�G������{�T��Ǽ�?��?V�;�����f�x-\>/(j>�j�!��#Ғ�����é=���t?C4?\/�����!���2>.FS?�?��b;��X�$�i�>�5C?�?�z��뤿x����=��?�-�?��>?G>L�rCC��L	������?�?c��>d%��u�̾��Ѐ?��9?���>m�����ٰ�kj�>%a^?xBI�3 ^>��>��>���%1��9G�\���`#O���8>����k7�l���A�;Q�=>��>�P�ꋭ�O��>��<��'���TN�Y)��`L>/�3=��!?!B����>�=q>��>O�8٬����u�@�$%z?���?+r{?U(?�l�������<�}�>R��>�
>��>&|��%{P>�?�*j�؏����U�(?���?x��?PLw?M�[��ۿvɢ�<ۣ��֤��b[>�^�=�� >�(��;y=b~4=������r3>.L�>�h>��>�c>َ1>M>뵅���#�Y ��z$���^9������/��;T��8/����� ��?y�e,���$.�y5ѽy(�^���Ǽ����R�>`!�>���>w�(?��>ߏ�<�z��ܾ�q��ጾ;�)� ��M(�'��H�~�7�����:�r����^=���a?���=�zD��Z ?��I�;�R�>�W!>�
�>w�>3�s>;��>xc
=!e>�v�=k�#��{ >/�>�B|>��}�����m��V����>x=G?Taq� ^����s�B㼾���D��>
�?�R�<�O>�J��b���c��>)=&n���
�=�}0=��=���>-H>���=���"��f��g�<E͂>/�/>�N+��a=��"D������ �>�,���.>_��>�b?�\?z�)?�*�=�A�>P��>��>5��>��>@D�>v3�>Ay ?-G?J�?�uy>/�p>�Bɾ����>j��lT=%]�9L���ꕾ!�>4�2=��u> �=�Gs�P��=�~�=��=��<d��<*�>#�1?�?�˿>9 ���%x�7$6�~��<�ܡ>�� �U�?���>���>�>�v�=0j�AW��D�]�p�>���>�O>rSs���9��<��>� �>�-K?F�?��<0���)�=P)2>�>\?��?��>ѝK>j����8�Lܿ� ����]�>�}�=�=�<����%Na=�_�;&�����ex`=a��>'�>�D�>q�w>�<>]��>ג�>�=�>�W0���H��9Ž8)N<&v�=e��=�@	��
>�����p|�:'�=��뽘�8�\j��ߘ��k��\G���V ?��$?B�>�$=X�=�XN��w=�b�<���>�SX>���>����|�aWQ��cj�Ү�~w�>�>M?82�>շb��8�=L\9�(��>{��>`�<>�R"?3�>�؄����Q��1@<�m�>wl_?}q/>r$�7�������`�[�S�>@�>fF��<<�?1Er?�����[�do7�̪W��,&�l{��#�:<������j��Mg��۾�iξ��$��=��>�[�?e_V��*�=����Ī�e�����ZE�>�\ѽ-{?j-������0�2ǒ� H��]��-�>#�o>0_&>bx�j�???�k?��>�(�>��$��'4?
m�>=�?��;?��2?�m%?��$?��=7�H��}���B�j5�,b���Y;jP����=�%,>���=8���-��=���++����¼R��D��&Vѻ,Ś=��;L)^>���=��?��)?p�׽v��=E�������	�>��> L�>a�M��x����ڼL�>��2?�RH?ä�>����GH;��U��!�`=ϟ>?X�B?�6?�w���y�ۃ0���x� %>�O ?Jj7�ހ�=B ���
����c��>p{>�(?>�ci>�_t?Z�@?�qK?���U�N�:�+�N�N�V��:7�;�KJ>�B>�s'>���I)S�nyc�ˮd��-����=N�B�_�=�yB>]Fv=�>p�>�?�>%�=�8�-a��휽0>I$�>'"?��>d����<��������\v4?�����Z�����
�s���V>O�-%>���n�>+�ͽײ��,)Ŀ��^�Y��>���?I�?xT�?�[��-^�X�>���>��ļ��=lZ�A���c?��*�>Q>����$��~>1Of>�� �f���1��i��t��a��y99�{�������2ྮ뤾��8����uEC�7��=;���ǡ�ܛ���`��fIټ7B������ež�����?u��?�F�����r|�'7 �.	���8=�t��C8��bϾC�о�F��\�þ[mþ��Q�&��C��06�i��>Bp6<럝�k���cF[�����⭾>@9�>�L��d����I�r�=-�'>6�g��v�'0�����o8f�Y?� +?uv��5�Ѿ2�~=��=�c�>?K�>�'>�%����'�/��>��U?��?������%呿T��=,��?.��?0�P?9��=2���G@�rg��#�2?��6?�43?h�@�E���\'��B?�,C?�?}d��:�����^�1%�=ʃm?����^�;>s�H>*�j>d#���e�3��=�r�i	=�
=�$��X����D���&����>ڨ�>$~�>@X��
�����>����ƅ���e��̾�s�>��q>�ޜ>����Ю=�v#?�z>\��w���cP���x��ƚJ?�_�? �?�3?�W��DϾn� >��0>�!>��>���<ߩI�'Β>��?!��<㨿U4��9O?���?���?�M?��}�\������橾?骾6)+>ӧ�=J�=�,� >����l�6���|:>hѭ>�Wy>�|>��O>��9>��>	�����"�u����0���-��P𾑞��1Dr�ޥ��)���g����/E��6�$<��#�p� �<���2�vۀ��3���䇽^�>0�k>�?2��>�w=y���@=�v���`��o�#���&�,7������+���j�0I��QG�!�湶�8���o?��c�81�=E��>W:��/�>J~�<M�=m�8>e
^>A D>o��>��B>c >#�>��=�0�<�bw>�*�>L�G����^v����9���>�N?4�꼙��9��� l���ĽQ��>��?.�=��<�}K��:�_��>��=$B��@c�敼Tȕ>�9�>B�s�S
�>LV�=��X�J<�>�BX>�?a>�oM>p�s���¾�!#�a^�>*4۾�T�=gTp>�(?j�w?r�3?g��=@w�>�e>T$�>���=SEG>�,J>�;�>hI?Z�8?.x0?\o�>˝�=K�b�{�*=�>R=H�fZ�p;������)��O&<�'5�r�3=i2p=b��;K�[=x�.=F��;��;���<ש	?�L?��>;��>���Q�b��$�K#�>G��=����Q?i��>(
 ?��>g+9>�\����V~���Ș����>���>���%��#�5?�M&?	q_??�>fv2�S�ƾXZ>���>�#?&�!?�>*?V�>��н��X���w]�I��Q=�9=ԧ<�S ��y����|�x�� �<=�=N��>`z�>ﰀ>��h><�>-w>���>��>>����T��3���"�<�кI">ω�=��ϼ��>�h�=J.y�����M^��YҊ�)Cؽ�� ��`*=x�?zZ=?S�+>!�!��a��H���r>�U�>��>5h?/��>�=4��ږy��#F�'���?�ڃ?E}�> A8���>F[��{n(=
��=��>�_D>�M�j��>V]��>���>�hH?�>��ʾ臿�˂�]�:�}��>�c�=)y��y�?��U?���C[(���a�+@��]>�A���*���$$��1���@������	"��64Ž�X�>�Q�?m�����>�R �����"�����"��=��ؽ��>j��雵��J9�hྤ�_����=�9>���>���=��N<{��>L*?�;�?��Y>a�>~�>��=H?�S�=�E=>`8?�ZU?��H?�#/?K>��ͽ%����_R����ۖ���=��]=m>%�=�>�=��W=��2=��<�==tG�X�׽bQƽ�	<? M<���<�1I>���=�#?ӲK?Rl^�		k�?@Q<%��=u�r>/�<�_ο>�Q�E^�,N4>Js�>_6?��-?�+�>�ry�T9�*_1�Ǌ	���i�g�?�_9?���>�}q���}����ѓ��_�>~��>"�1=J�޽�žQaܾ���>nW�>��=J�V>�i?�RK?��d?�M^��h����x��mK����=qI��UǠ>�E=�{���ƾ��X�#���`.O��L���<�;���,�1�>���>d��>���#>K�D>Er�l긾���=@��p>w1�>v�>��<��)�WN����־�%6?�z��N�����=���:3���+=�J�E�/� ]7?�Ӭ������y,Y���>q�?u��?XD�?\�=D�F��_�>2Sa>`��=��u=��ɾ��G��%;�Fp>�P">lz��j� �7�h��h�=Ӷ��g5��H��W� ���ÿ+CK�+E���y��շ��T����U�FY����Y�;񕾦�����kX�z?��;,���B�G���$���G[�=�?�Ş?&找�0� m���U�rg�;��ؾ8dD�B������Q˾�cq������wb���/�����]>`(��,����a��X8a�r�>���>v�?�3˾�ZԾ�M����<ӵe>�i���1��Ȍ��N���e-�5f�?��&?V&ƾ� �3���F�>��<?���>��(=�y��4N=��>��6?6>?�$�:⟿���ƕ=��??��?��C?L��8b>�Z���0��7?�3?i��>�T��2�ݾ��
�?J?=?�W�>Mr���MN(��@�>�RW?��4�)_>Z �>�#�>�ଽ0y`��C$�I:���
=�3G>��O�����[���&�>>�!�>��>��x��i̾#�?���������7x��쾶E���O>	�?���.Q ?-2�>���<�ƾb���b=���߾��;?�S�?c��?4�?�Aپv�뾀Um=%Fv�<I�Y��>[�>R��GQY>�:&?�e���ܐ�;��5&�>��?2%�?�g&?�����ڿ)5��F\����ޙ=��4�$�>/T����>�;�
<����Iě=3��>�_�>_�>)c>��=�ڙ= Ņ��u!�@Թ��N���9�d��$��T�|�}j.�	]����!��������\c97�	����<�9�Ҟ���<*,+�
�>Bc?���>�R�>Gl`>��;>�8y��P���-��㡾��߾96	��G��-H`�cK���!���w�U���%^������?�G=�J�>މ�>�-���W>+�>�N=>FA�=���= �.>���>t��>�y>�:V>�tt>	��=�Y�>�>>`v��}L��]��L�����=gw?*Qr�*K���E���l������>=�>(~�=�G�q����w����>���bI[�����u9���g>�
?��=>ƀ8:2M#�3qž%��8�=p��>��=�_����'��Ej"����>%�����>�};�X4?"|�?��?��=c?g�>�ٔ>9��>ܐ�=��>
�?�o>?��b?�3?�'�>��={y3����=*W�p}3�"t��%��<!gݻ]{6>$��<!����0�=M�=���=u��<�ć=�8j<�U?��??�i�>Yj?�s���oA�wE�� ��٧�=��G��>���>���>R��>��>2��=��X�&���߾ R�>���=2o���Q����=ޒ?��?�q?7�e?�]k�H�����������>��?/?��>�^����6��E����O�^��,@��������l��$P�lSm��p�[����n�>������>�>�Y�>�2>�g�=;TJ>z��>�U>�/]>��S>w�½˞�=(�<���6�,����2=�,��a<����"�!�ս�L�m$���?y�W��< 5?S�"?�锾F��ї����*����9��W?�G> ?,e0?�,*>�����~y��n��
?�u�?<$?pѾ��R>��>��=�;�>�r�>`�>���r$=_���.d�˒(? ��>NR=C>�9��Zz���8�v'B>�r$>��@�Ȉ�?>�h?�Ի��Ͼ�Y��J0��}8��]�>�w*><�,���e����߽A�G����ݾy3�X�=�x��>���?K���G> �֯�:�r�(9)������=}?-�m>������ξ;�.�P�"���~p,�yrv>rM>�=>�?%G�>X�?�Oe?Z!�>y��=@n?�<	=.5�=�!?� ?î,?"D?h>
?�?�x����B���k������)a�)�=XQ�=�E�=�T�Ⱦ�0WZ<ŵ�=���=�N�=v߮=���5�=�_>:�> �	>�L?V�?����F�$>�w`�h\	�7)M=�>= W7>�	��e2�5A.�eӧ�=�?	+?ޝ�>@P}��P�	�.�M���䑵<M�?�A?tL??쾼ъ���7���h����=>��>Un�=ՅN�?�ݾ�3��[|<��>��>B��=��>2΁?��j?��?��4�S�V5���Py�VlѾ����?�
?�؛>�2:��)Q�n�1��u|��{���<sK2���<�oQ<o�:>܊�=/>��O>ي���$=�u�����k?����>�ƛ>O�?rs�>�z\=�Z���kʾxPJ?�t�����x����ѾBX�H>�FT>�6��x?�����|�Uޤ��\?�HN�>O��?g;�?�Yg?8&:����d�`>�d\>�>;d;��J�Ϫ��7C�!w:>Ia�=�3s����3����`>��r>����}/ɾz��7=�^���W��=f�AZ��'���⫾En����x�杚���<c#���e��u�޾��ۦ���&�vE��X��u��u��?�'l?Z��=Q�o>dtl��\��O��2U9=`�ܾO�0�i%���t���;3�r���Ҿ}q*���h�3�3�������>�	> 䀿�1X�8懿!�U�]K�>:V?~1���ʾ�@H�����Z�>��=���?����������?[?��*?�>z���о���Wt? �?�7>�((>Ԝ��+�>qhU>��?y�r?�nc�͕���x����=R�?d��?��8?����?��p�N�n?��?$��>�򖾀#ž�^߽��?m�;?l�z>���n��[���?)g?"J��`G>7Z�>��>q���Fp�����S���7м��">�M�<ܮ� Pc����Ǽ
>��>�U�>P�0�L���x�o>�ξ�6�͐B�bF�������">�� ?h�ݾ�K���3>	��>%#�`����D��Ű���7$?�B�?��V?�2?��b���Z���Lc>�s�>e�>��>��й�0�=+N�>��¾��Z�#���'�"?�"�?�C�?��?���B����g��ʾ�2���T�>��c>2��:"j�o�>k��=�h�=͞S���>��>K�>�s�>��>�$l>��>@G�t���U���#��|;K��\ �[
O��X���1�.����Z�	�5���d�k�����M�DɄ��ľP��gױ����>���>J=�>ë?�T�>,e�>T���Qr�~2#�z�sǾ����<��΁�tc�����؇����R�݌ͽ
_�# ?ݨ�=��z>�q�>⽽V1�=
��>��%>�'T>
�>�>��S>���>%��>��G>�e>��<�*>
4>{�~��	���JP�SU��j�ͽ�,.?[�(�\⓾?Z��Q �\������=�F�>��->�b6�#J���q����>%��=��Ͼ�kн�>��A��>{�>*M�>c�����ý��ƾxk�~�K>}��s�½v��#Y��h��d>$��>h��T�>%��>��'?�oW?:h?�|�=<�>��&>-��>��~>���<� >��>6�?NX-?�(!?�Ŝ>7�I>�#����T>�1>R�y�B_ֽi�h�s-�p^e�o�>㠂=i�<��q>���LI�]��>��<������='�?��>?oi�>���>[۾��\��2�R��7��:]>�_?	��>��^>�!?=G�>��>qm���徍hϾ���>�;>7�Y���f�bM��d��>L��>�,?)�
?D7�Y>о+�=� O�=y�f>K�>P��>���>��<"����|Vο��>�<�+����Gl<]9����QO>�2�=
�K�s�3�6��<K�>J��>�5�>uN�>���<:�=l!�>%�0>�Z8>AK6:I�ʽ�=ye�=A����N���<*�`��Ԁ<Z�P=R�׽�P	��'R�q�E��R(�m��΃?��?���>)���ၾ	*��c頾�>��>DC�>#t�>�7�=�@�LwP�.a?��P��S�>�Wa?j� ?�.�TW�=΀�,����>Cͩ>2�*>:@������>���Կ���>��??V�>�D��aX���g��{
�F��>�->h������?��n?��辪	;���E�N�)�*�L_>�l>)Y̼<�~�WF�/�'�,�(�8o�6<��O=T�>��?�Ԕ�_��=�@��Rv_�*��;`���Y�=W�>�p�>��� �b����]�|�<_��>�3V;q�h>w�?0�#?�8f?��?,��>}�N�f�?�Z	���>#��>7i�>�%?_?e�g>�$�>�J�<�Q�^Ǩ�ጾ�x�=@��;��_=�J">,dºKP<�==};>��9>
%���C���� 㺱��=g�>z�=+��=�_?�o?RN�<m=>cO�<z�ս��=��2=�F><"��ט�2�Ļ���=U$?P�-?K��>5$c>Y�;����A���I��:/?7�E?ƌ-?�ޗ>T��=�Ŷ�v�Z����ޝN>W ��J�
ڍ���f�X< �4��>7�x>��$=��b>��q?R�I?R�*?��1�7*T��cz�.E�Zr���R5=H�>A�>�π=�����,�5�S�:�S��^ ��.� �*����=Rm=���=�$>>�;=+q<y3ͺZ�M=��j��V�=�����7�>�E?��)?���>mfI=L���t
��)I?���p�J���h;����->��9>P^�7�?Pb��|��ۥ�U�:�1^�>6&�?'��?�na?��G�����_>��Q>��>�i:�K�{��@딽k�+>e�=�uv�5�����;sZ>��s>ДýNξs.��3�V�¿&AV�3���0��+�����C��R���;�C�P��o�|/��3-�����8<�<6O������19̾ 6ᾨ��?�?`�=�Hz���7�c�Z�ھ?�.>�ǝ�QU�����,��^�v�\���V���=뾼�@��q)�3���^>F�н�̣�^����A���>?��>E�=?�-�D����� ���i�>4��G5��c��A�����*��jh?	2?a�Ѿ�����=DU�>�ϛ>�c�>�*�	)��!��=:?�5?a`�>j���n��=A���E1�)�?u��?��(?�ei��;E�&v�b���C�>@<?p��>~'����7���W�Sͯ>D�/?5�>�<2�KN���6� �B?�.�?�M����|>d?S��>I[�=����-�<�K�\�	=���<>��p>!���o����G=�)8>�a�>-+�����'խ>�=ξ��a���T��0�i���*�4�k�?{�پ�>��>��j=t��jā�8
����w�`�2?dR�?L�y?�&?��a��	�̑Q��_=S�H>���=��t���>���>eS���b�;���_%�>��?�?Π2?��t�C࿺~���`ܾ�_����>�8�=y��=?�����=�=�v:�����r�=[c�>w�>i�\>oVc>��z>�>�ȅ�� ��~��3$���F%��9 �����߾F�+��S���J���ؾq�Ǿ|=����K��k�*�1���<�N��T��<�#�>��>�R>ؗ>(� >iգ�Z�;�,�X��Hܾ�S��������2��u�^�I���&���х�6�վ�(�>���=-��>� ?�q>e�>ed�>��x=)�=�,�>e[>��c>穡>��>3�=W~>A�7>��">a�P=����36q�I�F�!�o�7��\)?Ί�����;2�y���M,־�'_>z��>��)>��1��L���Dz���>��H��:��u����9w>:�>pp�==N$=0P��������:W=ܔ�>k�>O) =JX���'���T=�"�>9����A=7j���L?82w?�e?Zھ>��?��>�ʹ>)d�>A��>S��>�I?��?�+Z?v�	?���>O��=�p������/��xӽ��޽	ɽB�����q�"��=��=:�=Mz>�.>��]M'=���=��s=�@S=�?r�3?9�>`�?�B����=���G���A�e�>	[��nk�>�l�>�\�>�?�*{>0`M>��Y�R=��E���.�>m� >�>T�-�d�Gt�=��>���>�i]?\�T?O����u���˽2>�b�>0�?|��>ɐ>��+>>W`�C<���޿��0���!��q<�R�<���\����Y��4�=�\R��D"��Q=a~g>đ>�.3>D�G>��>!�P=��>^�^>���=�P*>�;;~*�;ϐ���N<ҪȽt�= R�=7�G<�G��ƈ��.j��2�׽:g��l?ݽcᦽ�:�>LP?3�0�+��Ծ|��f1���L�>{��>
��>P��>K!�����$n�!o_��vܾ�z�>Łr?i�?ӝ��B�W��>��>5��>"�>{be>ֺ�=��#�UO�Z�8��}?+��> ;>U��<�R?��W�83��>!��=������?��?�d �~l���!���6��(�bA�>�#�����P��V���I��+��VZ�sޣ���R�>��?��=��>
P(�X���;��5���H=��<=1{H?���>
����Op�^<��������� �Lî>���>���>��>o��={�r?�PP?�H?Y9�=��?���= o$?��?&�1?|�D?"eC?ȕ�>��!?^��='�z����ܲ;�ԧ==�׽��=+tx>i^�=�Z;a{ >o>(�� j<z�n�$�A=��u=?Q�=�h�=j�>�s=>[}!?&J;?`� <0]m>\�=c=�[��=�fU>���>�$��9ϾŤƼǖ�=�I�>�$?؞?���g��
�۾�$羸ȑ=Í�>���>"�?`G�=�>=4���c��l�>>�>��*=K��j��h,F;v`�Ğ�>�-X>��#��}�>žb?�Ax?f�5?'
~��l������
��*�¾Wc%>YF�>�p?k���9�־� -��-��#a�.h4�� :�/�
�G���ܳV�=>��>�O>"$>Y�=b[=�$�i��e�	�/��>U�i>7�/?t��>��=�ݳ��(��!I?�`���)��⠾�VϾ��!���>��A>j��J�?�:��b|��{����<�$��>Q�?@4�?a�d?3i@��a��U>\G[>�>6U�;�F��(��-��w�/>[��=��z��왾���:d�]>c�u>{;½�E;Y���`�+����`��Y������Ú��eо�eʾ��[�By򾓝d<A����Ԗ��P޾��w�?�+���C����xǹ��ɾ���?��p?�8>6>n�W C�pھ[���y±�'�MF������}��m�ݾը��Ѳ�,r�9�Z�(c �m�=C26�J"���x���=��w�;1�:?s���敾=]��6J�����=h ��=8.�:���ݮ���K<�H�?YJL?��K���J���þ��=h#?���>�'�>�b��u8���=���>6{b?9�m>
R��>���Eg!>Io�?��?h%(?�v&��aw���2�$���W��>���>�>��S���g���Dgo>�C?��>�,��ǒ�l3��K�D?��?��)�o C>"�>,��> :0���վ�/�a ���==T�Q>��>
�'��y��c���N=	��>��>XR6��F�Y*�>ݰ�.���܆u��CP��C��<�j@?ǅ4�L"��i��>0�<>��!p}�9���5�e�b?���?C��?�p?�)
�d����>�M��ژ=e)�>��'>"s����>W>D?A'��n��؇�>��>���?gh�?�#?�&��_�߿@���K��7���������<��>Z+�?s�ϰ�;��=뇓���>��j>��6>2�>��>�ʐ>QUh>=ʆ�E*#�i���ҟ��v?X���
�8L�L����>���!Ⱦ��6d׾��*��B����)�7�\<�*�x,p�$;d�X�s>�>ͮ�>D:�>�L>&?��f���̾2
��"� g����)��J��T'��~ާ�����]����<nT$���<?YS��iM>#�?�!����=��#?�G�>a6>)bL>ca�>�?�`>wî>�j#>���>�/:>�d�>t >W'q�T�C��4��ч�v3�:�B?F�i�*龮Mg�}��O����=��?��>bX3����t�sC�>M��O&������+��f�>��%?�4�=�ٴ��`���(Ⱦ3�r����=U��>&�%>E�B� h�/H���[=n?E���8!1> >��@?2�p?�7?6Q>� ?���>a$�=�E�s�o>��>b�>r�"?��>�Z*?���>Z��<ʨ=��^��i7�*eR�h����>Ξ
>\�=+]0>ڿ�>��,>܄�=�;�>�*>@�����jQ���>|�.?��>�R!?[-?�ZOb�lZ������g�:�*�	|�>;��>��>>'�>���>�.&>��]��'����>P�><O(�d�9�"�>&��>e�>��Z?��*?|żR8�f�����=���>~�?"��>=<(>}�1=�J�;�\1��8��|!��è�4���X{�=!�����k�ν��ȼv>��[>���>�`�>9O>_(>C�>N->�ג=�M>�L=Uр=���;��=,:7�����B���	9=A⟽�A������}���?0�]N���1����>w4?4���e2w�;�gQD����� #?R,`��̢>��C?�ږ=V��l�h�߂�W/
��*A?1�B?| ?C��Q�>γ�>��<�<S?�+O>jL>��m��e->4�z���W/?��?�1��N�K|"��ɜ���$�>2�̇��v�?��h?&�!������n*�$h��&���>��=�Z�9k����gX6���̾7����zc&����>n��?���<8?󦂾~{��6)h�R`�����ZAB�=��>�����Y�������̾�k
�����N�H*=���>��>���> ִ<��]?&>;?�9�>I��=^?�?U�=<�>��&?�1?0�=?q=2?�J>�G�>�)�=����}������䟽����G=|����z��{
�j����=�@��B�8��dB�[��R`==��=��=Y��=�t?x�?6u��L�=���iAS���ݼ��n=Ζ$>�"��II�@d�<�=;��>�&?��>0[R��N�#�	�y�پsƊ=�.�>^
+?���>,�m=,}�=j�۾C��{W=�F >t;������9 �v~̾A�!�Kq>� �>���=�GQ>fU?Ț4?S�j?���%�j�u��2�I��]Z�ʖI�cI�>Ȃ+>��"�p씾�����J���Y��45�`���2ͽ}0>L�ؼՑ��7Y�>Zh�=z�>1Պ>��<8�U��3ƽ��>R=�>d3�>�T?Q/�>.W0>�7�|�����I?~���z�����\�оxl ���>�\=>]��V�?3L��}����%>=�:>�>Em�?���?�9d?W�C��J��]>��V>y>�1<�?�)8�\���l�3>o>�=�Sy�G����;0�\>:y>R�ɽ8�ʾ�E��KI��Ŀ-X���ϖ�����/;¾h����{¾3U����ξt龂ܨ��x�= n�\%�7̘�*0o�gY�>⾆jȾl�?��T?��=�x�>����� �������Ѿ���Z�����ﯾ��������)��9K�o��m(��O>�w��r5���Kp�1�@��0��*
��G-?E�y��hm�z 4��8N>x����&-������v��BrM��8�?	Cf?�t����J����RN+��9/?���>&e�>��Ծ�q�<�Rp>]�8?�8?�?=�掿;���c3�:�C�?1��?�8??ǩL�zB���zf��?��?���>H����;}��9�
?fA9?RA�>'0�����������>I�\?D�M��!a>�&�>á�>�>���GW�V����/��n�8>���,I���h��:�s��=1��>�M{>|8Z�4�����>%�Ҿ�q��?j�?�B�gA�O�O=r@!?@�"�H(>��>@5�=�H'�N�d��ɐ������lz? C�?�o?��?���g�,��t����1�=F�e>� ">���<�>Ɠ�>�kپ}p{�y6��)?�H�?��?��?���Uݿii��Vx󾧀־ҔJ>�ۥ=�M>���<�=1�L=*�C�����G�'>��>ra�>jÚ>���>��e>�6]>�&���"��l���,��X�!��ﾅ*�@8���U��-�����Q�Ծ���k���7/���u� 渽���һͽ�vȾ��&>�g?��>x�>:�>Z5>�#��坾���ξ�[0�k���2�nͮ�����o�����.1�����r�ɾ��?��2<FN>\�:?���=�v�>���>ö�>�A�=6�J��>��>��p>_�j>��v>:\>�;~;Fǿ>U�>��~�x�U��F�������8�s�?�W㽹$��I��]��.Ӿ\��>���>�]>i/����ǀ�Dd�>xM�j���`â��>�臒>M�?g�>����f$�:�~�Y�+�=��>Ǐ>�QN���Z�f��\>�=�U�>n���O.>�����9?��?�sr?"��>�U?��>0�=�c�>V�8?3��>Us?��X?��%?�6?JJ>;�>��뾋��;b�=����CJ����_�=m����ݼ�C�<�Y>��=�z��١*��m>ؗ=�t����EF ?�c8?Iz�>��>W�g�{F���u�DJg���N>^셽�
?�>Bn�>$~�>�k>�x@>���2޾������>(�T>��z���u� �=u�P>���<��?��E?'J��
Nؾp�=���=T�>_��>�(&??�;>��=�l̽����ۿ��1��`*���Ѽ��;R�ջ$a2�A!���%����0��~���=���>7��>�/m>[��>O�?>b�,>���>�qs>jL=b��=�d��=�<ق��+������c��˗R�89=P�R�����D�'��+	�Y�̽���XJǽ�0�>v?�yK�'۾�4q6��`�����>g^T=�p�>�y�>sV����%�G֊��d�������?5r?_� ?-����m>VHO>��>)�>*NA>��->P^����,>���Gg���>�q�>[������'<L���#;��\�>���=�H���?�2�?�	�`⾖:��L�=C�{L�=���=v�¾υϾ�ʾ�"���������a< ��}?<�?����q>R׷��板;u���\���>~���w?�>�(���겾�-�����O��$�=,��>�J>:2�>��#?��>�r?�7?p)?m� �A�?\n>�=?��?\&'?��?0�=?i��> ˋ>��������EV��,*��0��|>G�p>��>é�=HТ;-<�=0Š�O��=�'K���N>�Q�=��>��W>)��=�(�=�?��??�Z��ٻ��=�+��
>���>�@�>�t��a`���lJ=Ͳ�>?��L?��?���������jf�m�A>]0?���>�?k�]>��>�-�����g�>�C�>�~�����=pMǾMy��HB��)?w>��>[�x>�5�>�(r?L�+?� U?��_<�UX��ߐ���b����=nkk��t>bk?K��ѥ�����p@���_��� ��&Ƚ�N,����Q=���=�:F>�;>�,^>�b�=9�<�0V�&�&�p��<�)>o׳>`�?]�>���<�������4�H?����J�;�����վ·3���>7�C>���E?��'�|�K䥿�Z>�d��>���?2]�?��d?G�;�����'`>��X>�`>��"<��G��� ��戽A03>���=<�~� ��-�;�Q>>iv>e˽��̾�侙-K��о�|~�^-��uv���9��
������ndӾ�rѾ�9��1¾l�\�ib��xi��:Y��\o�}k���l���پZO�?d?y�|>ֳ�>��D���)����]�J�{\��$�������u�ղ ���!��-׾P�)��O��F��`��[.>�gR��2��}�r�A>Q����=k��=���>a�˾#�����=��+��@|<��ս���{��O���Jqr����?�PS?&����H�H쾡3��-
?M��>�U�>�{����=��>	B?{;?���>����ɛ��4>ip�?4��?Z3;?#�C��gM�|��KI�ڷ?~�?m�>1.��Ѐž���G�?5?�>E���;������\?5Yq?�]2��U>��>Y��>�н�����z�8&h��'���*>L�]== ���f�q���*�=mˣ>a�>bC�@�����>�=��kL�<:J�x��q���9�<-I�>�|���9>��[>'��=�j��Q���=���+�{<>?]��?��Z?��.?@7꾈���lg�ɳ�;�X�>(�>��N=�J��O�>8��>�微dq��-	��9?���?�i�?�O?��g�1��I���#Ͼf�վ%�>���=�\1>+�Ľ�r�=�>G��=��i̲=�x>���>27�>�	>rW>��c>*���"�@��"����)�TU��g���<��kH��H���ce��ξ�й��bK��c�m1���I%���=�|��q�S>i��>���=%�>>�ܴ>:��>AD��0w"��p��}��\*��h��}�ξ'@��q�9[G�;�
��C߽�L���ξӶ�>����&�>e�?�Ͻ���>D�>O�=��>��>�~>C�>�4�>"�m=#+K>�8b>��>'�>�y�ݨ��D�3�/��6��E>��c?Y9����X���_�o�@��|���e�>���>�4G>Du�=���w���>)ؕ�p]ƽT=��v�K;:_>$��>�߻��`>�ξ�vپ�Ԝ=�Tj��:q>�o�2"�hѶ�j�&�2Q�>P�Ǿ��>��=>�"?�҃?W.?�2>�;�>x>S�>x�=���>�ͪ>�Ez>)y�>G-?J3?���>���=#���2>>���������`2|<uJw�"�z���%� �=w��in˼��=$�=�"Q�#	��)=ٕ�>�_G?�y�>ّ/?j�7��g���N���&<[խ>~^'���?b�>��>�Ѡ>�?���>�vȼd �J�E�8�>\$�=�"\�}�x��|�=�> }��� E?��?Al�>	I���u\=���>[�>5LO?��?ɿ�>��u=���̿��3�9��x�6�������9E��=���]�D�,�{�,>�Ha��I�>$��>ݰc>s�$>@u>@�,>hh?xNv>~�8i�>"i���!���.�p�r=L�:���E�&��>���a�R=�3�,���~�ԼC���Xƿ���?��>�L��L��2�徴K�/U�8��=�I>��?vq�>p������r���^�d�}���>��_?�|?�1��oQ\>ߚ��H��=Y��>�S�>��>,�����6���Ǿ��=�h�>Rg? �>�e+�-�C��b����a)>"Ǽ�1�����?�I?H������3�7�p�9�Ѡ�6�s�R$H���n�z�������>�bx�HP���!��y�>!n�>!�?�d�;U>�V��<��k���U�w�;wS���op>���< q���1!���D�r��d���O@�>�'>�>�>.|?
d?CG~?��G?��#?]�0�?}J?v$=�e?�b]=۳B? �S?6h$?�??�+?�Rm>������{�hD?=7��<tĥ���=F�>%�#��u��e�]�=삛=�ӟ��@S<RP��9�;��=Ib�=|�?-U9?ぉ��.�l2�>��;�n��e>V�?�j<����X��`�?/�
?�+L?�3?x��>����d)��bھ���=�T?~(?���>C5?>�̬>J�c��^�P<&��>�	Ƚ���C���:�u�C�+���>t͙>�T*>���=p#�?�Ո?��? ��%*��~���v�V�b�ؽA�������hI>6�pe&��\d���{��U�h+a��2�=E����h
������,�>�5W=ۜ���x>�y>m">3�=��H>���<��?�m�>82?K�>:ns�ī�c�)�xJ?�����������Ѿ�
��a>�9>*�� ?�t���}��ƥ�(�=����>���?�P�?3pd?1A� C��U^> �V>�L>�4<�@@�ί��:��y2>���=��y��㕾c��;��[>�v>��ǽͱʾ^�w�I��޸�̫f�]ѿ��˱�����mT�B|t�~��>"����zD�׾�N^>i/���6O<"Yy�B���s��-x�Ћg�N��?�.�?S�ls�=��F���:��G���3>U]þŊ��D��,˽L-����� /���3��/�9��ow	����>�־i���Cޓ�������5
�>4��>^a�k2��S:��S��@m:���N�tW̾��DU��U�P�,�8?.�+?�Y�����Ȗ����>�`6?#=Z4[<����5����>o�?=�?�����s��j����@=U�?p&�? U?:�۾o�4�9Q�֭��+ ?���>�x�>��վE��U7�����>Ë?Ea%<�� ��	��Q*�v�A?:0{?�R��|>��%?���>�]þ�I�����&�Ⱦ;�=�zn>��>=QzA��]���3�����<@$�>d �>"=A�9���<� ?e���Q�p�[�G����]��*���>?���A��>B�=A>� ����䤍����??
�?�x?��	?}����a��w����R���:>x�>o�/����<U�>���>�2���Tn�g�9�3O?��?z�?w�I?�e��Oֿ[���c���I'�!e�=z >p�i>\�｠	�=���#C߽�%%�l�=��>6Af>J{�>��9>�VR>�w+>kN����#�+�������Ń5��u �<�� C��b������
�m`�N�����������n�o� �&��B����r>���>�t�>���>��>Y[X>c40�����S�������u��?�ξ���P�̾:�pVٽb��Xz>��I�n[(��=?�n>`�=���>"�$�1G>[�>��9�|��=@e.>b��='��=���>�Q>��>h�(>��>?j�>ID
>aI��0-@������k���80<jOx?�6���>���ݾ�LE���>�w�>`W#=�1�����v���^s?���=��Ž׊����h�M��>$z�>�RK>	}S��!t=���{߽�>|�>M��=C�;�e��[V��J&=��>�����p>G �>`?D��?�C?���<��?�d�;��>8y�=,�>{��>c��>�&?��F?R;1?���>�>B"��� �G��=*�n�y���"m �@-,>�����a���y.��\>��<z������=ՎV��Q��-��c.�<�*�>�M?3�!?Kw.?^+?�LM��>��]G��0�>�<@?�\N?�7?��>�S2?���>�]�>r:ؾ� L����>t�=@B �E�a�0�>��>1wm�bBb?kya?�g>��o/=[9"�	{>��?�E`?�q??�	>k��=r� ��տ.��G���	�<���M���X�l���P<>Nl���W/��=���>	>�?>��>�^�=j��>4��> �
>_��=?>@�.<T��(���@�U>G��*�>���<t�i`�~�������.��c>Ƚb?��oQ����?�P3?3=d�,�pH��f���Z��cE>_�f>�/�>#�>|^}��"��c~��~C�}i����>�^?���>2EоbW>������q?"q?E%�>��a���6=X�u��P�>2c�>��F?|�??�/Q�!�I�4�3�1/��ؘc>x�=���9�Ɛ?�PO?�q���߈�2�C;����7׾ۧ����w���K�f�_�V~$��+�Qd�2��=Tb�>gƴ?�ڽ�g�=T���<��Ax�DT;�K
<��G�㦈>gj��t@�9'���t������lڿ��>g��a�lX6>�:>?��>�!?�
??1�M?8�p?>B��f5?ݬd��U+?���>��>?d�5?C�?�U?���>�W==Or뽀$�N�8���v��ʐ����=1P>��=�&��fV��ޖ���F�KA5�zs�=���<m�$�<<�=��>d>�=L�?h�0?c��=��=��>D������:���>T>�$y��Z=>�U�>�>�`5??	?M��>򧚾����9F���="�?�T)?'��>��>���>s@�aD���}����>�%�P;������ޥ� �"���>o��>9>�=Ccu>s��?�s??�1?�����O�!���l���Q=��ܾ�4L>�o^�c>����{��#c��_�|�?��ǋ�X�(�Ŀ�<�?�=��>Y�>�{ݻ��>Y��=�,I>�*�=�t�>#��>=��>B�?�G?S��>��+>�@k��b�.�I?V��zV�����S�;_.(�UL>+-C>~`���8?uA	��{�����>=�?��>4t�?ʠ�?�oc?��C��0��V\>��S>\l>=r<"�8�?���ތ�w^5>{��=��~�:<��[M<hw[>B�q>"ν,G˾�x㾰1�����pQ��ʠ�����ݓl�u���ɩ���">�9��f�=�G����+�
����v]��2�:����z��P���c�?�T�?�����I�=*-�X���׾�՞=�1ľm��t����K��mǾ����e
	���'���H�$H6�Y�?>z���,��\�����Qȉ=��V=��a?\-J�X��=G�S�R�*>�����l���QǾא��F¿�{��MB?E�?	��WO����n�I�?�?K&>Co��sa�|#_>�-�>@$&?�"?"L�k�������X��h�?���?R�B?wr
�`�2�cT%��%��g�>=��>]?$)̾�v,��dG���>1�?�ں�����䋿^'�p�H?G<�?�-U��>�v?ZB�>lA���Rž���Ɣ���>ƽ.����枩�#����^=-�>/��>��齨a��fr�>Jz۾�VK�M�Z�����Hr����>3����=��=f�=$������e
��N�o�??,�?9�k?ߒ?N�ξ�-f�5B���G�d>�ގ>�<��G<�@ >
�>��Ӿ7d����G�?�?��?w&V?N�Y��Tܿꌢ�G�ʾ��Ծ���<*�0=f�\>�ҽc`A=BN�=�l�;~#���>��>@s> sD>%�T>4�V>Z�>A��sT#�8��������#M���%�^��S�����z¾�m�>╾�ܟ���&R��կ�!P��c3���#�\��>/� ?�h�>xK�>�d�>c=>��#�.�`V��[&q����?_׾X �j۾:ә����d%,����üT�!��M?X~�=���=��>��q�9>�֋>fj<&�=�I�>�y_=7\�=$
�>+]>�JK>2�>/7?=�L�>�3)>�����6��悿��� �>-?���Ęo� �t�Ü��R�g��=��>A�=]�����v���|��>��@=����G�o�T���=�}>�g�;��"��&`��u���gG��*�=`j >�w�=k�c���澝�龡���Q�>�骾�Ȟ>�^�>LG$?� v?��3?�\�f��>r��=^��>��=���>j�>@��>��?Z0<?Ϧ-?u��>v�=��ɾ1�:��{s������,	����(��ϋ�[��<��{��E;>��<<�>�/F=L	�0�U�-Y<=��,=1B	?�2<?У�>��H?��>%#~��铿wg�>�[[>��->b�?Y��>]�>M?h�8?���>֞&=�����K�V\�>C�8>�l��n���Ă>��s>���?͒�?���>�#f����>��6�
D�>!?�W?;�b?�˵>̵">N��$���6@�08���q��K�=�=�I��ܪ��H����=���=լX>K2�>=yM>��6>E3�<0H>?q?�;(>�	�;.��=����s�<$.��Y�)>	T=J�u=ɖ\�Y4�2n;�T� =$ҷ�M;�	0���o��`�#�6A?ă#?����GM�����ɾ,�޾�>h��>��?\��>�u�=FZھ�hV��0;��{���Q�>�]?Gi0?���%>2)�9�<=^3�>^�?��&?F�n=�}\��X�_nS>+��>6�c?�s?�T����Q�f�(�e��(�>��=����ip�?�:5?�ZʾI��"���G�9`������K�������7о��Q�$e���(�x8�� ��Mt;>?��>���?:�=p5>�i/��l��k�o��:�<vm��L��>)�?�'4ƾ��TO�c� ��⾹xL�T+>H4>�w�<���>�>�>�gA?�R?۔o?���8�?Y��>�T?]X>6�L?�+S?ط?�~?}��>�̉>tFe�_��64:��+
=F�2�U|���d�=���=C�=�����=�=.����Ce<�?���w�y���;=v�G=V4L=h�?��7?�с�K�^>|�>5]#�����Wԣ=�3?�y��}.���v> <�>���>±G?��4?�P�>��V��������"�;z6?�/?2��>_>���>�R���:�ݛ���>�w�����D���$מּ}�.=g`G>->7>���=$�l>Z��?b��?�?�C��ȍǾO�L�a�h�v�ǾXb�M�/>a �5����j��MZ�]����}��s�Vz?�D��n���0p뼽��>���< �ƿ�=-��>��D�# �<O�n>��>���>{c�>4 )?.�?�v=ש����3��J?�>���W����{���݈l�� �=��W>����|:?��a5v�����g7�xD�>ا�?�E�?�%c?~�Q��c �o�d>]�G>�
>��}<��3���X��77>�-�=>���T���A�<ՁI>N]>�<��{]ľLoҾ�m�� ��ӗ&�g���s��� ��( �V�d�hC>U�{��>�۾�=5����D <��ҽ8f��b,�S|��Hv���&�?�_�?��0���l=��1�)	-��e��l=�;��\���?���<�ܭ��w��z���[ž&Y��/
�3��j�?;F��$��E���"� ϭ��!���
?�-*�`�=w�y���<KN<?���n�Yڔ�3p��
7߾_�.?s�%?2��q���7��"U?y�G?+N��4 >4��S�{=�%�>un�>b?�ł��쉿�7���TF����?��?E�6?U&I�~�.���/�Y������>�c�>.��>��D����n�3�>eE?D���=(�����g�"���7?%�?2�K���a>��?���>�F������2��5->^��L� =i=�a־�q���=I~�>�Z�>���[}����>��)
G��K�/$���½#9m<7o?6�J�/>��>{B>1�%�+Ί�;����1�B~>?�,�?��V? �7?���ܾ�e���=[g�>���>U��=4��ކ�>
��>Zۚ���k��p�G�?�#�?I��?�MK?�^\��kܿؤ��'�ʾ�x־G��=�le= �`>3���d>��=V�.=�{j=�g�=,��>�0>>7ji>̉d>��>k=>�E��Dr ������ʭC�o:!�`�G�����S���t��p���O���Ԃ��\u���^�6I��t	���%�V|��o>U<�>�ڇ>YР>8
�>��~>:$�F��5�	�YnνgT'�-�ʾ+⺾�������� �(lӽ���j���$�WW�>E��:�
?>�϶>ٗ*�)/�>ټ�>�k�=y��=j��>D0>�^C>s]�>pl1>C-0>�4i>T�=s4�>�{�=�i��9�'�
쌿Ģ ��Q:>J�(?/����K�Ȕ���'����m�����>���=�l7�mqʿ\���E��>z���0=Qs�O�=��>�vQ>��l=0�	�'C��bU��s~�(.*>�O>&��i�D�#�0ш�( -���>���ҵ�=�-�=��? �z?�%?�Ra>3M�>'��>�r�>��>�j4>�0b>G�Q>n<�>��0?�.?��?K�=��پ�q�=���=�]�KJ�r�U�8*�<ٓ��3o==�&I�kM>'Ҡ��O	���<>�a/=��h�7�� =�?��6?���>�VL?���=�j������>�'r���?��?�?��?R��>�-?�p�>wC���I�8�%�c��>�v>>���$/��k��>���.ш�v~t?�~?���U�}>��9"U���x?�~? f?c<2>��i>�L��ӿ�P���A��<)���<��d=���rƐ=�C�=s�=�A ;�!->MVf>3�+>2��=�]�>�:�>pȁ>;?�>��6>CCu=���=�>��WZ��uZ����<U��)��X$�>��<-9��,"�NOL=��;��Z�PPl�]S��xN?O�2?��3��	6��e!��ξ����>���>�
�>^�>�X1>]⥾�{��'�@�,=��>!�J?�		?�\ž��6>R��=/��ۖ?;7?���>Mw������@��ý�=}">)�x?�Q?�_�Cia���-��V���s>[��=���Б?:k>?����l3���)�U*���n��(V-��հʾ=�%�G���׉$���]���/>���>;��?r��<T��=j���,���Jz�b��\Ҽ�^m��}>Y��� �e��.�-�Z����+���z<��ؙ<ݧ�=��>>]R$?D�>�??�l?��Z?&4����/?����P�?��=
? m?G�? \?u�?@�>Dv�=�bB�}���Hi���^�����2��=��7>q�+�����=H�=2���D;��~ܧ<@��U��o��"=A.��?h�3?�Mڽ��#>��>��Խ�c��I�>�M�>�t�#�1�Ԛ)>�?���>E?�*?�1�>ӇT��2��\� �X��<�,?;�?��s>��>���>����^���D��p>b�����!۽�l���1�{�>k@H>��>xp�>�ވ?ȕ�??U[9�`�'�uQb���W�Wж����L�\Ѿ��:�����0=��l����`���J��0��2{:�X+�cP�=���>��=�BC���>�e=�/��W>S"�>�R{=p�>4]�>a�E?O�>P�>;EU�Ә�x�I?�������}��x;��.��>��C>�T�� [?�	��X|�`\��!�=��E�>���?P��?y�c?�nC�nT�'`]>9�V>��>@d><��;��l�����y�7>��=��z��镾
� <@sY>��v>W�̽n�ʾ���B�6&��7n6�v�� 	.���@��^�G�h��<�����-=�C�/��=�O�������04��F�فԾcw����?��?�{v�E�_>ٞL�lN�!tz�dK>)�ξ�߽=L �t���g.�8z��7ľ�����l��?-��@���?�f�������q��+��k�7=��*=���>$���r=eCC�Ǡg��X�Jy������S��d��?n���m?��?����!�hy��a�>��?�\a>�"��c<������>o��>�{�>�(�SO�����.��3�?��?S�J?��'�ŷC��4�	c¾���>RB�>_ >P��Ր�j�G���>S>����U@�<"���A!�]p?f��?l5��Hn�>
�?(��>�۽��q���]��`7�͵>M�����I=�`��!�оㆋ��b7�2ۙ>%��>6����5���>�=��kL�<:J�x��q���9�<-I�>�|���9>��[>'��=�j��Q���=���+�{<>?]��?��Z?��.?@7꾈���lg�ɳ�;�X�>(�>��N=�J��O�>8��>�微dq��-	��9?���?�i�?�O?��g�1��I���#Ͼf�վ%�>���=�\1>+�Ľ�r�=�>G��=��i̲=�x>���>27�>�	>rW>��c>*���"�@��"����)�TU��g���<��kH��H���ce��ξ�й��bK��c�m1���I%���=�|��q�S>i��>���=%�>>�ܴ>:��>AD��0w"��p��}��\*��h��}�ξ'@��q�9[G�;�
��C߽�L���ξӶ�>����&�>e�?�Ͻ���>D�>O�=��>��>�~>C�>�4�>"�m=#+K>�8b>��>'�>�y�ݨ��D�3�/��6��E>��c?Y9����X���_�o�@��|���e�>���>�4G>Du�=���w���>)ؕ�p]ƽT=��v�K;:_>$��>�߻��`>�ξ�vپ�Ԝ=�Tj��:q>�o�2"�hѶ�j�&�2Q�>P�Ǿ��>��=>�"?�҃?W.?�2>�;�>x>S�>x�=���>�ͪ>�Ez>)y�>G-?J3?���>���=#���2>>���������`2|<uJw�"�z���%� �=w��in˼��=$�=�"Q�#	��)=ٕ�>�_G?�y�>ّ/?j�7��g���N���&<[խ>~^'���?b�>��>�Ѡ>�?���>�vȼd �J�E�8�>\$�=�"\�}�x��|�=�> }��� E?��?Al�>	I���u\=���>[�>5LO?��?ɿ�>��u=���̿��3�9��x�6�������9E��=���]�D�,�{�,>�Ha��I�>$��>ݰc>s�$>@u>@�,>hh?xNv>~�8i�>"i���!���.�p�r=L�:���E�&��>���a�R=�3�,���~�ԼC���Xƿ���?��>�L��L��2�徴K�/U�8��=�I>��?vq�>p������r���^�d�}���>��_?�|?�1��oQ\>ߚ��H��=Y��>�S�>��>,�����6���Ǿ��=�h�>Rg? �>�e+�-�C��b����a)>"Ǽ�1�����?�I?H������3�7�p�9�Ѡ�6�s�R$H���n�z�������>�bx�HP���!��y�>!n�>!�?�d�;U>�V��<��k���U�w�;wS���op>���< q���1!���D�r��d���O@�>�'>�>�>.|?
d?CG~?��G?��#?]�0�?}J?v$=�e?�b]=۳B? �S?6h$?�??�+?�Rm>������{�hD?=7��<tĥ���=F�>%�#��u��e�]�=삛=�ӟ��@S<RP��9�;��=Ib�=|�?-U9?ぉ��.�l2�>��;�n��e>V�?�j<����X��`�?/�
?�+L?�3?x��>����d)��bھ���=�T?~(?���>C5?>�̬>J�c��^�P<&��>�	Ƚ���C���:�u�C�+���>t͙>�T*>���=p#�?�Ո?��? ��%*��~���v�V�b�ؽA�������hI>6�pe&��\d���{��U�h+a��2�=E����h
������,�>�5W=ۜ���x>�y>m">3�=��H>���<��?�m�>82?K�>:ns�ī�c�)�xJ?�����������Ѿ�
��a>�9>*�� ?�t���}��ƥ�(�=����>���?�P�?3pd?1A� C��U^> �V>�L>�4<�@@�ί��:��y2>���=��y��㕾c��;��[>�v>��ǽͱʾ^�w�I��޸�̫f�]ѿ��˱�����mT�B|t�~��>"����zD�׾�N^>i/���6O<"Yy�B���s��-x�Ћg�N��?�.�?S�ls�=��F���:��G���3>U]þŊ��D��,˽L-����� /���3��/�9��ow	����>�־i���Cޓ�������5
�>4��>^a�k2��S:��S��@m:���N�tW̾��DU��U�P�,�8?.�+?�Y�����Ȗ����>�`6?#=Z4[<����5����>o�?=�?�����s��j����@=U�?p&�? U?:�۾o�4�9Q�֭��+ ?���>�x�>��վE��U7�����>Ë?Ea%<�� ��	��Q*�v�A?:0{?�R��|>��%?���>�]þ�I�����&�Ⱦ;�=�zn>��>=QzA��]���3�����<@$�>d �>"=A�9���֥
?d̾�����k2�d�e�-�>
h~>�<?fB�Զ�=t�!>�׻>q<��l������i�?�͟�?9²?��?,�2?�-�Z?s�����SP�>{�?��>#r=?���>6h7?�>��#����Ɏ��'?���?г�?}�?�M���_ؿ9ᨿ8^��=�Ͼ�r>�-7>Obe>����.�=���L�<��H<�B>�f�>&��>m�~>��f>0U>ez>>U����.,��2��*���1��"���Iw9�������4��9��%Ҿ1���#
�,�M<ㄞ�g^������5=o��a54>/M�>��'>��>�8�><>X���I@7�w����9���Y���<<��w$�R�j��s �7C��M�����k_��et?o�=�#.>�>)�y�>��q��>,?�����=��=f�>�h>A�>;�=j�a> l�>{>�D~>��=���?뀿�9�G�O���7;$�C?�*^������2�$/ݾ�=��kp�>�?lR>H'��7���x�m��>d�C���a�o�Ľ`��t�>]��>��=v	� 2)���u�v���=��>�>B�{�/<��)���q�=\��>�T־=�=}�w>B�(?4�v?[6?Fě=�~�>ٽa>؏>���=RL>zQ>:��>B�?U�9?Z�1?q��>�@�=",`��=��7=��>��tW��벽~pݼ��#�Gm�<R!2�\�F=6Ps=��<:`=�B=�ż:�;� =��?��H?���>�4W>c��q6]��N��{3��5�H>�D�w^	?8*�>?�?4p�>��>!��;v����k��2���@�>`�{>z���V�q�u��=��>?e�>��c?Ƕ?g�֖ŽӒ�>N��>���>f�"?�RI?���>V�>�K�v^�R2޿ŏ�`kW�S!�1+�ݼ;Bj�һ�:�����.ɾ�׽���<�>�]�>![�>\>*P�=�@�>.��>�ݡ>[�~�I8c����������I�q=C�zսZ1ļ8"D<���,��L�� C��Kk<�nϼk	���?�a ?��2=�/��`oM�b�ƾ@��Se�=6xY>8��=�2�=�o��� ��c�s\Z��b��p�>j�b?�ÿ>d��D�=(�����<±�=��>ћ���n>'8�=f���/�=���>�O4?/x_>�U[�]6O�����fV5��+�>�˖=O޽S��?��I?zg�<�a�&'� �I����т�l�d��k��VAȾ�9-��,;� ����⾑72��ZK�J�>TU�?�xK��!�=���᠘�����z��Q�&>`70<�R�>��|>Ee��J��@ �']���ۼ�I!>�z�>1�=1	�>�=?ks?j�v?���>�?�]̾/j?r��>��<?�W?q�;?��F?�I
?��A>���&z�~Ǵ�ԟ߽��u���H��O��2�<�n�=Gm>)w8=�<�x�=,Z����ǽ]H��w�<|ʚ�A�:���=�U]=�<�=�J?�ED?c0��f���ͺ9<� ��52�&J�>/��>RnD��Z��Iԍ>���> �?�V?���>ך��9}۾��ҾK��z�ȼS�?�c?��?g�=-p>�����`<eN>���>rhu��N4����Dl��KǼ�ի>_�>��=R�>�q?m�F?� "?I��_h�G���I�ƾQtý���x"��,�R�=���<7��C���Ʉ��}U�iT<�k���=knl>��*>��`=���f��<sս�ǽd��<��=�3�=��v>P�>~?ș&=��ɽ;���Vc?�����@����n4�6�=�ԥ>'�>�����?���z卿�����oD��qQ>b��?���?+ډ?i�L=�;��n��>>�?�]>ֆs>�\��Th���>�S^%>Ɨc>�k��� ���j�>p��=���=B�P��5��J2���7������wM�Ұ��:S���bɾ:��zx���U��	������J�LC,���T��獽+�=C4�)�{�N������[1�?AV�?�I��2ҟ=���S�H�<5뽾"�>bϾ����A������i���Z.���ྙ�)���D� ��U���b�>�g��	"��P?K��/u����ğ�>�tQ?���᡾\&*�ڧ2>�M�=c9�������KZ��y���|�?�%`?jΘ���&��6���u��o2?���>�F>����=�=�0>_�??Ix?�#Ծ�S��R v��W)>k6�?���?��??��N�.kA�I�M��f.?�w?��>�H���̾o��F�
?�p9?(��>'N�9�����]�>9�Z?�bN���a>��>ɂ�>��\����$�xY������t�7>j
��>�~g��=�>S�=�Z�>�tw>��\�Xݮ�\�>��d}�Z,3��?�Xg#���>��?���:B�=�-�>�S�>�-�،�ֶ��� �h�w?	�?j�?��B?��@�޾�I���t�>n�)?(m�;���=�,H�\"?���>Z�3��|��cl���??%��?K\ @	�.?�.8��e޿C���{����¾�>>ߩ5>��m��>��`=�]�=��-�_�>���>�r�>��h>�>u��>�>(e��#�{����嚿@�;�٘�`/��NN��V�s�}���
��Է��������M=�8J�s���]���Q�����R��=c_r>���>�U�>p��>��f=�ԇ��)�����H���U��'6� ,��@۾��q�f>����	� ҉�ԙ���??8���R55>��>ni׽=��>�E&>1���m+>4`=�"�=�Q>�>>m�H> c>� �>���=��|>5�=�����Sz9�FN�)��;��A?��_��H��I}3���޾�ک�ʂ>	�?�NS>�E'�������x��0�>��5�:�c�S ǽޯ	���>�>&_�=��z�B�0�ͯt�����'�=�ׄ> �>D^��e����d�π�=.��>j�о��=Y�m>)�(?�mu?�2?��=��>TS>̍�>�خ=��>>�I>m��>�?�}:?.�5?
F�> �=�C]���=�'=�8�8Z��u���&������<1<�QD�͛i=�og=%I(;��A=ЁB=�q���<�7=�?i�M?���>_�>z�f��p'���h��K�=���=s�=�7�>�`?`�?��>�6�>���=�&����$��e�>b�>	�y�p�����<���>G�>�5*?�g3?�ؑ���T���j>���>e�?~/?�!$?�C?E�x>k|��`���ڿ�^#�=S0��q`�Ԑ�.�<h�>�ת�/�����D/��+N=�Ls>F0�>�w>�wL>��@>u�^>Ec�>j�J>��<S�;e��M�ʼ��=��l>-�.�d�@�ѽ���<0���곸�?1L��g\���
�^]i����y�
?�?�]=
��L����&���R �.?�^*>�i!>(��>S;�=T���ct��l�r�%�]��>�Ӊ?ζ?
#���=W� ��cx>���=�H�>�O�����_)+�	.�����=���>�;?�ׂ=oq$�1�{�sWu�(�N�Q��>�?�==r�h)�?�K?���VB�CR!��<��g�FCn<mս�ď�cþ]%���4��ؾYS ��l��4=�)�>�7�?�!A�{�s<N>�� s������H����҈��lx����>GE>6z:�ۜ��+��˺��%���(>OP�>���J��>�"=?��6?��l?�?��Q>4���t?|IF��Z*?�o'?t(M?I?�m�>ޕ;���>�>9�������)���j=�"�=c�+>�ٍ=��
>��6���>yG�=�=��\�`�ڽ�f;=��Q��l�<�ۇ<w��=T-v=G?�$?]g��1!��Wݼ�B&��"!���=}��=�*,�_����)Z=��i>���>�M?�W�>�y$=td޾�Ӿ�0�Q�Y>�:�>j�,?y�?ɴ�=���=`��s�F�w�7���(>d�T�2q_�i�ھ��ľJ/��kp>��{>
-�=�ԁ>�p?ǮC?:?�M� �>�����ͽ��援���<}���6>JpD��j&���y����x-�T�<�7/��hw5>��>S��=x	=�;��mH>��>���=
�=މ>���=�>?v��>,�Q>#�1�[]�y����a?�g�{�.�*'�a�UB��$y>�8�>T����S?%��Q��c������lJ8?���?�q�?��E?��F���)�1:p>-��>L��=�<*=�OU�T����A�_�>wn�=�9ݾۅ �`(>�hD=���=LfS�3��h�쾅�r���ȿb^��x��Ӹ��^�|E�R :�->�h�� ~���[��G8��j8����<��=��+�����it�W��3��?���?_�'�]>dr��Z�H��#��= Z���01�h⳾�➽L=���3�H�Ѿ��r-�=d���&�W_R>G�8������V0��j����Ѵ�>�j?t����Q۾���;>ܺ>K@潱���y��UZ��8��4<?*�Y?���j���ͼ�M�<ފ?P?x3>���^��[ߔ>j�H?L�?��@�Ab���;��B�=�B�?� �?��??
dK�A��\�R&��`?��
?���>Z��mP̾���u?A?:?��>@o�^ ��:���0�>b[?�gO�Ahc>��>�>�;�Ջ����/����zx�c�4>��?!���e�q8=�<�=��>�*x>�v\�����\�>��d}�Z,3��?�Xg#���>��?���:B�=�-�>�S�>�-�،�ֶ��� �h�w?	�?j�?��B?��@�޾�I���t�>n�)?(m�;���=�,H�\"?���>Z�3��|��cl���??%��?K\ @	�.?�.8��e޿C���{����¾�>>ߩ5>��m��>��`=�]�=��-�_�>���>�r�>��h>�>u��>�>(e��#�{����嚿@�;�٘�`/��NN��V�s�}���
��Է��������M=�8J�s���]���Q�����R��=c_r>���>�U�>p��>��f=�ԇ��)�����H���U��'6� ,��@۾��q�f>����	� ҉�ԙ���??8���R55>��>ni׽=��>�E&>1���m+>4`=�"�=�Q>�>>m�H> c>� �>���=��|>5�=�����Sz9�FN�)��;��A?��_��H��I}3���޾�ک�ʂ>	�?�NS>�E'�������x��0�>��5�:�c�S ǽޯ	���>�>&_�=��z�B�0�ͯt�����'�=�ׄ> �>D^��e����d�π�=.��>j�о��=Y�m>)�(?�mu?�2?��=��>TS>̍�>�خ=��>>�I>m��>�?�}:?.�5?
F�> �=�C]���=�'=�8�8Z��u���&������<1<�QD�͛i=�og=%I(;��A=ЁB=�q���<�7=�?i�M?���>_�>z�f��p'���h��K�=���=s�=�7�>�`?`�?��>�6�>���=�&����$��e�>b�>	�y�p�����<���>G�>�5*?�g3?�ؑ���T���j>���>e�?~/?�!$?�C?E�x>k|��`���ڿ�^#�=S0��q`�Ԑ�.�<h�>�ת�/�����D/��+N=�Ls>F0�>�w>�wL>��@>u�^>Ec�>j�J>��<S�;e��M�ʼ��=��l>-�.�d�@�ѽ���<0���곸�?1L��g\���
�^]i����y�
?�?�]=
��L����&���R �.?�^*>�i!>(��>S;�=T���ct��l�r�%�]��>�Ӊ?ζ?
#���=W� ��cx>���=�H�>�O�����_)+�	.�����=���>�;?�ׂ=oq$�1�{�sWu�(�N�Q��>�?�==r�h)�?�K?���VB�CR!��<��g�FCn<mս�ď�cþ]%���4��ؾYS ��l��4=�)�>�7�?�!A�{�s<N>�� s������H����҈��lx����>GE>6z:�ۜ��+��˺��%���(>OP�>���J��>�"=?��6?��l?�?��Q>4���t?|IF��Z*?�o'?t(M?I?�m�>ޕ;���>�>9�������)���j=�"�=c�+>�ٍ=��
>��6���>yG�=�=��\�`�ڽ�f;=��Q��l�<�ۇ<w��=T-v=G?�$?]g��1!��Wݼ�B&��"!���=}��=�*,�_����)Z=��i>���>�M?�W�>�y$=td޾�Ӿ�0�Q�Y>�:�>j�,?y�?ɴ�=���=`��s�F�w�7���(>d�T�2q_�i�ھ��ľJ/��kp>��{>
-�=�ԁ>�p?ǮC?:?�M� �>�����ͽ��援���<}���6>JpD��j&���y����x-�T�<�7/��hw5>��>S��=x	=�;��mH>��>���=
�=މ>���=�>?v��>,�Q>#�1�[]�y����a?�g�{�.�*'�a�UB��$y>�8�>T����S?%��Q��c������lJ8?���?�q�?��E?��F���)�1:p>-��>L��=�<*=�OU�T����A�_�>wn�=�9ݾۅ �`(>�hD=���=LfS�3��h�쾅�r���ȿb^��x��Ӹ��^�|E�R :�->�h�� ~���[��G8��j8����<��=��+�����it�W��3��?���?_�'�]>dr��Z�H��#��= Z���01�h⳾�➽L=���3�H�Ѿ��r-�=d���&�W_R>G�8������V0��j����Ѵ�>�j?t����Q۾���;>ܺ>K@潱���y��UZ��8��4<?*�Y?���j���ͼ�M�<ފ?P?x3>���^��[ߔ>j�H?L�?��@�Ab���;��B�=�B�?� �?��??
dK�A��\�R&��`?��
?���>Z��mP̾���u?A?:?��>@o�^ ��:���0�>b[?�gO�Ahc>��>�>�;�Ջ����/����zx�c�4>��?!���e�q8=�<�=��>�*x>�v\�����X?ij�����W�� �E��=���>�D
?�t��`�5>�l�>���>fR��u����������ށ?�b�?�M?G1H?��1�a�ƾ$���6?�[&?��<'>���Ju�>�}?/�����wɾ��>���?;R@s�\?�&�T�п�������&�þo>�2*>!�\>����K׋=Vu?�.�<�R=��3>��> �R>gǆ>M>ܧ>�,>yR��ϔ&�cФ��x��3�>��!�|��ǝW���%��7ɾc�\쳾�Ӿ�H��
A��!��D�`���-�(������؞>��n>o�>��>�.>>)N$>�m���{A�>�E��?�N�� ��r.��V�.X�����|��Q�Q�3�콐�s���>K��Pj�>��>qc��� >ECb>y@���vC>�A*>�Ү=�O3>��>Y�:>��>6��>�Nn>;ђ>l��=ZɃ��I}�E�4�^4T�GI��ʒI?|�N���ה.�]˷�m?i�a;�>��?7:>��&�P�����x��z�>z��Ʌ�>��q%�<	��>n?�>��=�H<�WM�b��� w���>%�>�e>a��;B�q�x����YL>ػ�>-�Ѿ
��=p�s><�&?>�u?9�5?�!�=Ve�>��g>�ݓ>�4�=i?>>�aD>��>��?%�9?W�0?���>
 �=�tj�	�J=bQ=r&6��xi���Ž�ː�-�'���<yC���E=���=���;�Dx=d.0=d켼�^7<*6=��?J�E?��>���>�}��7�@�%P~���=x��=�Z���G�>0��>�%?D�>��>k��YX���'�u,�4�>��=I񑿆U��L]T�6�;>�T�<P~O?��9?R8M����
W>ߠ�>��?��%?�F?~�>��>��ӽ��
�.�����6 �C���?ݥ��7�<�q>+���?X������[=�V�Ŏ~>p	�>Z�>�LC>�%�>���>� �>Y�1>S�K=t�>���8�9�潤���sg\=G�a>�c��>���Q�<�e���˻��1;~�=�[�=�(G>:�?�x?�Y#=�����cn��靾�G��[�>rM�k�>m�`�V������x�c�f�m����;��>_[O?DnB?�@ѽ�} =�fo>[U>p��=�Ys> �ӽ��>v�<�Eپ��(��F�>��?	��>����!d�Nt��i���> >[=T�����?�v^?)��[��Z��P�A��B���A=E/�L�t��в��!%��7�"s�������tt��a�=��>���?�u~��_?=���|œ�Qڂ��0���|<��<̘�>�#H>��4��&��	�.�Ⱦ�CG�[ �<�~�>?8�<̈�>��=?�A?/�`?�V�>�Ը>v����'v?�of���H?���>&�?�FZ?�l?�R�=>����D5�6���xҽ^j�`'�(b��!�<�.=-yG>;D�=�Ն=��=������Ov���I��c���Q=�p-=n�0=ƀ�=�!?��??B�ǽ�0�!�)=�>(�"��W%��m>����B(��u>��?�* ?Q�Q?��>�L�Җݾٝ�����^�=�.4?Z:?V+?I�=Ӛ�>`�=� �,E��HԢ>���B����m�"����߇���>J��>i� >xӀ>Fy?T�e?'UJ?��J����j�x��À��܆��K�Xʼ��<��>�I
��|+�����^��M�d���=\V=���=��/>��>!c=��YKf>oDe��Wż�j���p=��F=s�y>�1�>��'?���;`��<���4�m���[?G����[�d��p���h��hk�>8��=�־�r�?��u����m��E.i��!��f�?%��?(H?��Z����2�>�Z�>���>θӽ����+,���v�[x5��=��ξ9��(��>�Y�<�#��W����D8�E�8��2�Ǒ��6�]�1�4�������޾�/,�b*p�P�X�0����=%������K�S� ���y�L<��B���X��b����2�?�?����%�ҽW�l�r"��=�w^=�<��2tV<L�Ӿ� ��ܾ�����Z&�Q�4��!����>�+������l�[ l�=���з>��"?бþ�Q���/�$n�=4O�=�hr��5��G���\��
�f�e�F?�t?�Қ���*�hc��Uy���?>�?$�k>����A��(�>��e?ϒ?}鵾5A���߅���@=T·?p&�?�Y??|[>�h�<��g�H?��?|G?���>�닾D�Ͼ� ��6	?�s:?�0�>I�%ل�1u���>�_?Q��\>���>��>"�õ����������k�����->�����t�$0Y��c7����=d��>�rl>�:l�![��P��>�-��z}�kk��6�-2ν���>�V'?���> >��>��(��ҍ� ��nܽN�M?��?��o?�;O?3f ��վ�	B�f�>Kr�>���=J��=���%T�>X�>����k����ɾp?���?���?�oH?��V���!P��!z���9���n�=Dn�=��_>�J��/>,��=j>e�='->>��>��>͵�>��>��>#֟=���_U��Z�����j�`�a�4�m���.���PG�j��
/������4ka���%$��#t�%B�܍��\���<�9�>�9q>���>�=�;�=^����Pm쾀�վ�UF�C*�N>�]/��n���0=R�����Sd=�E�����>�9�L@>ܢ�>��׾�`>�U�>�}K�_E|=�A(�̜t=w,&>e!> .>�>��>�B>�G�>��/>�o}�����sG0��8�F3ɽM�I?�_�Py���#�ՙ���N�Vĝ>�+?��F>����ї���y��ؼ>�I�3��k+!�s�[=�6�>��>��>=~�<#,A�Z����4��h>���>�se=鄨�	Q���J��k>_?�>N�Ӿ=$�=�v>G�(?_v?53?��=��>W>`r�>[�=X#G>�RL>)��>��?�:?'2?�u�>޸�=bU[�D=�H=-�>���N��ư�rܼ��$���<jG*���>=�Ly=�<q�f=0�3=iJ߼���;���<�?�JO?w�>XG�>sm��24��dk�`e�#R>��!���?2v�>X��>Ρ�>�r?g
=	���(���;� �>{l>��g�Ǿ��ٔ�����>���=:�S?�?4?�=8�A��&>�|�>��?A�>��1?`�?S�=����`���lӿ7$���!�7���E�j�;v�<�R�M����6�-������Z�<ʅ\>��>L�p>E>m�>�/3>7T�>�KG>��=�=a��;";�F���M=2���F<�P�b���ż����J����I��>���g�ؼ�e�>_�?tY=��������5�������>���>�>e]�>�딽A��H�H�r�=��0�s@	?�n?�v5?�'�L�>�=&=,hh>;)�=�*�>�V]>M�=>����6�Q2>�D�>Ԇ?>/�>���:��e���u�͠-��5�>��S<��� ,�?�b?�N��V1��U��Z26�r��8~ͼr���+��M,���!��)������S����=���>ql�?�Ղ��S�<�������+ ����ʾ�-=��r<k~�>D�h>�)4�5����<��Gા����U.=���>�kE���>4�L?�@?��{?4�>\ך>����Zs?��=k�N?��?X�@?�\?�i�>��>FX=�=8���P��9u���F�=P��=/܇=�%��ih>ոL<v.>S�
><�c>��k�[#�jz� ������=�i<�1=��R��<?�B:?>�������ϑ�=Lψ>�Y�Gm�=N�>��7[��0oL>Q�?��;?\Q.?k�>�j�=,Q�頾���澀=�.?��??O?^�i��\T>-��߿+��WǼ@�[>�����1��
J�I��~)�:#>p=�>h�8>��(>W=o?-�C?�_?1�������q`����?ɺ�m&�eΗ>:A1=2"�=a��� �pW��ŕs�У%��i�=�ӽX->��=<E>��=��ս5�.>ү�:��<ʨX=���<-!
=V��>�q[>��?��>�:�C
��l��n?'?'�nu@�5
ξ�[�F؏��6�>�~�>�8B�Y�j?-��Rt��ٞ�/�� ?���?�?�?��H?r���Z倾.s�>#�>�> >�ˆ�*"�<W(N����<dW�>�켾�F����s>�Q�>�ڈ>�5�h ����L
Y��s��7@�\�P��ԕ��蜾�������Ľ�¾�0=�ݾ�����v��AO�0=��#�����~���B�ݾ!`I?|�m?�~��~��m6�#�+���
¼�ھ��ݾ#������¾
	��e	���&���1��j����R��=�n��
ٚ��,V��Bb�%
���!�>eFE?����A��);&���|>mA3>~'��$�⾎\������l⼗9P?(�`?�#��h%�(v��H�}~?\&#?�U�>:}���_����=Mi.?j��>=.K�e��������=�A�?0��?}^@?�:��?���һ
�$?�>?F��>̃�/�ʾ���2�?ty>?�c�>�� ��3�����|�>��Y?�TS�T]>h
�>ȏ�>.QֽiD��{��Θ�t�w��2>f��� ����\�5�+�т�=�f�>*Ip>i�I�fd�����>�꾣�N��H�����E��<s?�y��K>�i>�[>��(�n��,Չ�02�X�L?ލ�?�S?>8?O����ۦ����=ܦ>HȬ>\��=��4��>���>�B�;dr�����?39�?���?�<Z?�m���ƿ����!��<��L�=BM`�Iն>\�����_�Oa�>��Ӽ*��<��q=ۓ�>$'>��4>>�?��>Y [>Gww�Q�#���ԩw��J�n%�����03R��[	���𼛥Ӿh��S��l>o�3jE�ɬ_�x[�H���+-'�Lb�E9�>1�?��?�?�>���>���>H'�����q���`���8���U�u׽��f���tR���v�{L��V��{Ǿ#�?�D����>��>Rw_=�}>��>��a<>�T>���=T�
>�'�>��5=�t�>�>G>E�=@�>�8;͏��j��J�G���V��?	>6p?=wF��S��0:�3�龉�����>��C?�0>5'�xh�� ��^�>�i��`y���M�;7>��� ?�?8a{>��>�Uv����J`��mE�=ӡ�=*7�>WM�����
��;iD>:��>j������=�>v�A?Da�? f,?��
=���>�3;>Y�b>κ=��A>�^u>��d>��?�U(?m?�j�>�~�=��_������G=�'�G�;�hbz�I�����-R�<kb��L7�X���G�D�(M.=N@=�|ʻ�� �/=��?@9	?��G>:��>�X��@Bm���g�yM������-�	>��E?@m?���>�z?:��>���>Ŵ���p���⾵�?��T��C�!�p��P>�r>Eaz>�b?��1?8���������>���>�.?_�>T�S?2ڕ>:g��ež�	�:��C�2�6���� =�ki���>�r�q�e����>6�M�x8���=�;�=���>_��=�j%?��?V��>��>�S>��=X�1=����**<�����b>���Hm��»�(��8��9mH���=�=���<��=��o�r3?o?>І<B����G�~ �
*Ⱦ���>�	�>���>���>�>&=3��q�ZF��`þN�>K�{?�?0�;���P>���! �oۍ>\D:>6�=�%=
(�LO����=��>R��>���>k~ <��@��oZ���{>�\�=����ۤ?��S?.���T9���� �:��ʾU��!�l�iQi��xҾC�@��>�� ���׾�����>�?���?а��K�f�/\���5~�ϋ����_�b�>�M>�6?Yr�>p&�����d������l(����>���>0f+>5?�b�>Ҹ�>���?�H?9��>M��A�C?4�輎d>P��>4 7?�v$?��>�ɚ>��7>�=T鹼05���@��q>#@��~��=���>��W>�������=[U�=�p=�ܾ��ܼR)=�](���=E�@>��=��>�m?)�?�ڰ��Z=7G>~"���k���h�����=x��=����<�U>�`W>~
?f5�>R�J?��=�m���C���!�=�a?&�?��=�G�<�Z>-L����ڧ�=4���p�Ѿ�����1.�Ǻu�m���T�>���=0����|b>}-p?A/I?��1?Z�[�ڇ$��[j�^(�AA�:,:���>���>Jl=�5�;�'��Y��wW��s&�wE�<�T�9�=0C>���=%iN�Uy=�S>��=}�����y��(�;�\��F��>��>�h�>|�Q>�H=�=�
�#�I?(���Uj���>qо'L�m�>-�<>��?�����}�@���G=�4��>Ј�?���?�=d?�C��*��\>gKV>��>%/<��>���#����3>w�='}y����m�;�]>�Hy>��ɽw�ʾ�2侀�H�$ ���O-�m�֦|��������־���=�K�p;
� �����Hd�҇����=6�����Uȵ�A`�?���?w��;��5>��.��?�z���2> M�+/�FPK��~ ����p�X���b�ྒྷd\��+>�]\�����>mǎ�T�����`^6�a>���>!^?��"������E��;�;D>G�)��S�v����:����2���-?ܷ%?����������n_>0��>t��=ֹ'��б��g����?H�"?�X�>�v�: �����=4���?kV�?7�E?��N��@�f&�������>N�>W�>{ǃ��ע�?h�:Q �>���>��m>OzN�����)�[�cn
?1��?c����>�S ?V�>Ԝ�������	���������=~>y��5搽U8�V�+�;�w�6��>�:�>Pc��������>�^�1J��SB��b��hL�q �<\j?E'�;$>��b>e$�=��,�ߏ�Bg���h;�8�B?�=�?S�[?��#?�ܾ̾/jT��u=X��>�4�>%�<�n��>��>���k�n���
��?���?��?�>?[�u�2�ҿ�����������>�>�ba>�ǽk`N=p��<���Ĭ<@>��>݆>D.�>X>�j>8X1>������'�����t5��ZE�\q���	�lIj�i��Qr����S����E�����nȽQ����QU�g"��=U�w�{����>b(?�e ?��=;�>/��>��%�M:������!"�Z�.�♾�+��3���l$h��>�Ϝ�)^��|['�����>�;~'*>���>x�>=��>[�>C;b=��>��G>��>G'���=��>_.>`Bp>���=uˍ>���=�ړ��99���J��	��\y�I�[?����M^�勚�����~�L� q�>�w9?+�><�D�vɉ�uׇ�G�$?��r��ܾk֯��nֽ&�>���>�>�<m��s)n�gލ���"<�dk>���=� �M���D�?t$=Ar�>�����M*>��=K?���?{zH?a��=O@�>Z,�>H�=�=�1>YC>�H�>���>�D?�Y?^��>��<���ΰ���u=�I�f���sBG�}r���콜)�= �E=�p'�l��<�	�a��=��k=6b{�pY=���=H�?�?w^�>��> K��I���{�:u$� �?7�8>6E>?�J?g��>aP?@R�>�5�>�䝼����s�¾��>`�<>��j�FO�Kq�>]!<�o����G?(I'?ӫ�<	�2���>��>z{?�]?b`(?���>Y>�ꑾn��:g��H)�s	=��=�	=���I��?V�=�*������	 >����f>��,>�ѵ>A��>b�>�<�>���>��	=i)F=.5D�f�	�6&��:�=.��;��<���<c����;��>���Խ��t=���my��y����C	?��?��9������N��e����C���c�>�Ζ>Z�>ٌ�>��%���&��`�%:R�//��GH�>�`i?g?�����sy>�µ:���=���>���>��9>?$ս�~4�����5���b�>l��>ȝ�>�A���T��^A�2����2>��=%�[�S�?��Y?���,N����F�Q�i-�^`�=𳓽w�L��a/�"9N���J�~N��w��e�4�0>��>m��?�K��_���0ڑ�ͣ~��ؕ�м'��T>R��>�G9?���>N�����1��Lō�c�뾆�.��b�>����hO�>���>�#�>��?KQH?1I'?�|(�$�?�X>Su�<�ܠ>�<?�G?�B? ��>4$_>�o�=���<;�C��k[�ѥ=+aA���$><9>�E�=ЁK�Ĵ�<���='m�=-K:��<�|=썹�3S/�P8�=�~>�?a>:�
?�5?�]�����=
YY�UT��㽟�=�F�:>#C�=@' ���g����>.E'?�Z?�?C��=����������I@="^?��[?�����ԼH�>�m����.iҽ�J�����qW����a�3��">#t	�B����c>�{?*LC?�(%?A��d�-��u���/���̻�5<���>��>t�=��־1\.�o>i���]�� 3��D���K���=�
�=�>�i%>p��=�!>)�3=g8Q�� 罿5�<Z�����>���>�F?j�j>P�=:ꪾ� ���I?-���([�Kנ�b�о�� �r�>'�<>`�3�?p�l�}�}���d=��"�>�d�?#��?�6d?fpC����`C]>ˑV>�,>��0<�=�����ᆽ%O3>��=4z�i<�����;��\>�y>�@ɽ��ʾ�Z侩2K��`��l=�s A���� ��SJ�7'߾Q�5��ƾ�J��U��j/h��Nd�/���z�����g�%-4�B̾߬���%�?m	�?:%&=9U&>@�(��:F�f����>�	��Pe �'�E�y�>z��x������Ʈ���J��XH���ҍ�>5����8��_����7�d𸽉�)>C2R?�y� ����뾮�&=
=�^㼵	
��m���ï�X��Y?X'"?ƙ��򃎾b
�R�>l+?���>��P>j�b�oa��h>IT?�c?M� 5��ͥ�������?b��?�>S?=���!H�C���Z�>�>�h?��-?�d�e��ӱ;��>���>�G>^jZ��k��P@/�Z�K?rє?�mz�l�p>��>���>�L5��KϾ�4�a�þ��=j��>���w0.����
[�� ��=�4�>���>|�	�n$о�8�>���K�M��g>�)�(SF�<2��>�k�1<>���>Y�+>g-��*���I���>���@?%�?�na?lu?̨ؾx�¾�c�	�=�,�>5��>���=�K��df>���>y� �g��
��?��?Pk�?cTU?��n�>Gӿ��!��������=%�=��>>��޽�ɭ=��K=�ɘ�-Z=�n�>���>o>C;x>x�T>ћ<>��.>r�����#��ʤ�4ْ��[B�� ���wg��{	��y�����ȴ���K�������:Г�y�G�]���T>�Q_��O�>A�1?��?Ā>��>A<?,�Ͼ�;�(�پ7�&��w1��5q�xv ��ii�9�־r�9=VR��Մ��o]����4�>E�k�>[��>�HC=��r=-�w>n�D>|��;Lē=P>N�=#Y>3�">�w�<U�>4�<ї�>\R;>�����f,��,7����ƅ���'9?�P�� DE�Ӑ���u���	�<��>'�?��>�ME��H��}�%�#?�gy��"������C�>���>Z�>��=��K��l��D�����=��H>��->r>�:2���5Rͽ-� >l��>�zv���>Q*��1h?��?@3?Y�?>��>ȃ�>��=[>�W�>T��>D]c>S�$?`n?�U?ڂ�>��=�E���$�=a��m���G�=��&����=�f���|= z��`�y=��<���=CTr>j��=�,4>��=��=B1?'u?�`=>��>�:@�C�8�H�L���9=xJ>�9��Q�>��>���>t?wJZ>��>�����F��3�㾱��>��;>
;�������R>d4e>��'>؊8?�CM?�s�V�r����>~�i>i�?���>�g?T�>l�P=̭����5P��_�`$�dG�ʈ>]>��Q�ls�=��=�2u�lK$�RKY�ĺI>�L�>AŸ>��>E��>��>�f�>�G�>k���(-=��\�\��-%D��0>�.z�<s<��C=�JA�Ҏս�������h�ͽ�c�=������ ?���>[��<fh�=f���L"����`��>�$�>9��>�??(�a>ղ���=�B�Z�����dG�>��P?#1?��Ҿ�>Ei>A,>Q�/>���>���>)��(���F�(�V��������?A�8>u:��:.�_�>�o;�]eƽ�4�=��n�֠?wQ?L����L��V�r��ݾm�<�{j���㾀��I�\��J]���5���e�޼�>H/	?��x?#�ᾨ%g��eg�T����y��=�m�hf�>��>o�<?^��>W�����M����	d��@�=��>S.ؽc�>��?}�?���?�� ?o�&?�/a���>�f�>~h�=ZΔ>f�>�'�>�?�Q�="g�>V�H;՚���L��U��zQ��R�m��P>���=��=�N^=��p=��U>�s�=��r�`���_�$D���nλ٪6>�3�=��%>�?q�(?r���Cb�y)>��=�{>�\=Z޾>����q����<N�>C�2?��?_�?�Cd>�]����&�-����=�C
?�1(?s�)>�jl�`9>���ͥ�t��>�ҼX���=0��CӾ�>Q��d����<>gjh>1:���	�>![_?�H ?��?��Y�ۛ2��N��h�-��I�<(�Y>��?�h�>I�:��B���K���x�<�B����:P�>��q�ߘ{���=PCr>C��=����=�J">�i�[;�U=w�=��?��>�?tS�>^[>�ǾI;侃�I?�7���T��r����Ͼ���P>�z=>B��0�?�$��}}�����C�<�+��>Er�?K��?Юc?�|C��r��?\>;uV>�>><��>�8�������1>�n�=B�y��A��TY^;�\>p�{>/Aʽ�J˾�!侽K�\���h7�X-L�z��_��y��%�>����t��ս�!w�S�%�����A�H�F�G���v���
����Lp�?rG�?|[K=/>�A�i#F�����=:����E�;T%�Q����/��Nu�����\����D�=8p�Q����>R�v�ƙ���#���p$�ua�<��H>hm?ڙ�č˾���.>�">�n=�לs�O��VX˽��M?;Q'?�h��۾p�$�7\>%�?��>m�->�I�W�?��ӑ>?�
?��<����������3�?�d�?�"N?r͙�O^����u���>0 ?5w�>:������?ǳ=�F?~?���> v��qyq�,`U�	�?-�~?�r���C�=ޘ�>7��>�`��4߾-�ܽ� ��x�u|�>A>�[���뢾��������'[>���>6�Y�Sϵ���>����t�C�[�>��(��^E�t�D=Gt
?�aԾF�>�y�>��=S�)�8ڈ�����&���C?r��?��Y?%o&?`Ҿ)�о>��[��;�@�>�S�>�e�<y3���>)�>�#�-�x��5��?M�?M��?ؾC?2�r���ݿ�ڪ�����tԾ>7�>lP�>#^=��A>�%=\��.{���l==Î>��>[��>��>uw�>��J>�����'�����jU��TDc���)�~��w���5�,d����@�ʾ�ھ!�^�q�߼th�)=a��雽in�j!D�zi>�'?Q�?��>�Mv>-^�>�Z��)r��A0�z�� $\� �ľ^V������ĕ�;R`���,�/�ƾ��
�����?�l-=,�>��>����g>\>�	>f�=�->�t>4)�=��!>�l>��.>�>	>>q�<�J>?z>>̟���b��l]�մ��6־���>�R �6�1��澵�"�&eW=���=5�?Ny?>P;1�c����q��?N.�桾ȗ{��-����>O��>�B��ۚ>8g��IF��l��ԛ(><��=�*0����0��'�q�^�,>�]v>v4��%ƍ>��<�A[?���?��<?1)>��>n��>�.�=�&>Dܞ>A=���>�G?4�j?Q0?R��>��=�䄾!	=y��m���X��<ڽ���<(���xY�{����=��=����=�`�=��=⟖<���<��?��?�.�>�	�>��(�h@4�vL�ė�<{4�>�4�>�/Q?}�!?�nm=�p?��>{ �>A+��x��M��O��>��>[���V[�F(<Ǣ�7K+>��$?�k3?OC�>10��ra�>�@�>��
?��?��:?�>�h>t�1>oq��B"��5'�o��z*u���=�X=񴻦�<�p,�&[�����p�> )�>"�>~O>"�d>�><�>�uS>����==�=jO�U5g���=�����R8=�/�<Fa���RM���<�j=����k����½���Κ?��>/�w</V།�����;e����>���>إ�>F?hB!>��#�J���^4�m@z��،>�!s?�?���N>��r;�g=$�>  �>"�>?c��������h��U�=�?�{>cK��w:X��$�H8"���=߇>@�p��6�?`�L?~-
�	�轒,��B��2�׮����?<����x@�o�G�zR+��8 ��	��k���=��?US�?�>�������[�<
p�1����u���w>�/|>��.?��>��z�n�킜��-`�V�侅�}<yd�>�1�����>��T?��>mi�?b�V?`pX?mw��N˷>�>�D$�t��>
�*?@�>��?$�>e�Z?�?�<�k5� �&��k��n2����)���q>���=�=�i>��7>�,>u3�=��ּz����8u<�.�;�\=?2>�1t>I�e>��?�>-?�Z]��]�2˼�;ƽRk�V����>�6�:!Rc�W�>޽->�[?k�>ˆ?�=�0����K�k>�)?��0??+�>ӥ+>�o�>�����*�������ڽ�����]�`_� �6��˒�G<�>�V�<�"��fl>'�y?�@?�u"?�l���+�g�u��+�V�o��<�(�>-�>F=v=�پ6|1�<xk��[�u-��=M��G�8:<�U>�/>f�->�f�=P�0>�������J���b뼯�����> ��>�g�>=�D>��=S���`	��I?O���c���៾��о]L �]�>�,;>���?o
�b~}����gE=�6��> �?�T�?B�c?�TC����[>[�X>��>�<�%:���쉎��#0>�K�=r�}�?S��w��;��Y>rw>(�˽ͫȾ�T�u�W����$%S��H��y͢�*����H�\H��(�>견�iw��ކ���h�L���'���K>��ýVֶ�hd���d�j��? �?���6�T>5�J����\~(��ښ����q���xn:��嗽z�Ҿ�˲�Z^�=�-�Q'2�3�����>� ��6F��q��b�C���=��=��&?VC��¿���m�������>�̑�N1 ��w����������j?�#?� ��N��;�����>�?�(?�$v>��������nY>S��>���>x��=�f��ۧ���a��۾?��?�eT?�ξE�/��?�me���>��
?K'
?�`����Ⱦ.=���>&/?��>�pg��r��ج��8?��?"Y�~<|>�E?j�?�I���~澠��L���	���>f�<�3��p
�����<P��>��?��Ƚ��վ$p�>��ɕH���B������5�IP<�Q�>����">�>�>�>]-�����؛���_���D?�)�?��Z?�B*?�j��ؾTL��f�=���>��>FO�=m��œ>f��>��޾c
j�����r�?�A�?�f�?�V?�	k�>Gӿ��!������
��=%�=��>>��޽�ɭ=��K=�ɘ�%Z=�n�>���>o>E;x>x�T>ϛ<>��.>r�����#��ʤ�4ْ��[B�� ���wg��{	��y�����ȴ���J�������:Г�z�G�]���T>���<\_>�//?���>T�>�>���>�Y5�N"	����������$�O�߾���h��+��!/;-Kz�k��{q�j4&���?��3�y�=�
?N;��.�=+>_�0>	D�=U'9><;=�t�=/j>N[\>�%>��=
\p>�c>��=�����o'�S�o���Й&�?O�׾w�j���;ĭ���ٺ�Q=�9?��>]�R�����V�Y�w��>l�h�q�{�����=�>���>�ib=*U�=�������a� �@\f=��= ����,<�Qྫ�X���>N��>8
e����\#���hC?V��?�/2?��$�
�?�!�>1<>� >�a�>��>��w>Ό?�G?�Q?�V�>�i\<�jR�*p!��.<f���7�8��;�~?����V>1��g��=���={\�=Y��>C%�=��=H�;<��<;?��?�I�>#��>Ib���9�>\�	�۽.��>
pL>ta<?x.?�c�>��?�>,l�>tG� {��Y��-��>��j>�z���f���2>�=��o=dq"?�)?��b=�o���>zΡ>�_0?�d
?�\?���>>�ټ����w��$�"��t�!��1=+�
=x&>�qݼ�dg���L=�x	���(�@cټqv�>��>ƾ�>}�>�>G�K>ּ?|��>xjP<9�q=�g��Ҍ������U#>�����;΋���$�=6�7<;_s�=�w�=(���Er>be���>��>꿘=��=߈&�
� ��^���L�>��>5�?}x?��;>_ �����L��؊��J�>[�n?�`&?�X۾��@>�r+>��F>e�>��>���>�fU=z������C�ľb�»���>T >������_�V�-��K ����p��=o���O�?Ki[?���Gqv�6!���F��<���=*塽�Ӿ���}�u��T���:�����t���Jߊ>��>�c?��]�8��<�Q�mԀ��"��,>��/�4>��=5f ?�j>d%���������DW+�雾��Q> ;O>�7�U
�>�?�?�C�?%+?�%.?dG�	Q�>�c�=�W>���>c8�>.�>#	 ?�>�=�-�>mI�ӥ���lv�����F��5@<���=s
>��a>��X���ͻ�O
>z�=����h��#�<B@� ��=��=�q�=7�f>��?�C?�T�M�ؽ��>>`0><>�2���g�>s��qU��tB>��	?�<�>0�4?	#�>U��>J��x�5�R�Vy�=:�?@�?6`�>�G�A�=y����.���묽�~�� B����s<q?��������/>5�e>��;3g>-�{?�[B?��"?�l��y&0�6y�Vw*��Y��D<���>Q$�>wi�=�>Ӿ��5��o�n]��)�Z����K�R�<���=��>�6>��=n>(�=�/��۽�V�;��ݼ���>��>��?3de>!t�=�%�������I?酡�`_��堾]о���>��<>�����?����}������2=�o�>�~�?I��?�,d?��C�G�R�\>�9V>k�>��+<FX>�����ޅ�K�3>n��=��y�=����;ط\>�;y>��ɽZ�ʾ1E�Y�I�v���H^T���!�qݼ�GQ����	��:��=�6��!1������╾+wp���2�e=:��B����s+�}K�� ű?���?N��g�=�|�k8�}�%��W=>�ؽ�G������}���G�����H��S���*��7x���:�ک�>����ҧ���F��O-*�;�A=�	i>�8?gc���ھ�
�C�4=��3>�;<�eҾz�v���������X?�)?g>򾬬��U�ƽ���=|	�>`��>W2<{:k��Y��Z]�>�o?�)"?vx��	��'#�����<��?�f�?�uI?�(��� [� �(�&�p�S�>���>�>gS���V����=�S�>���>��>�|*�y=m��,F����>s�u?2����H>5?M��>��A�v������оA�ҽ6ν>���=����s��1ML��Zr�1?O='9?�i@�iV��;��>�����Yd�w�W��]���s��1��I��>��?���7>���<V~=m⾌��P��[�ý˕c?��?u��>2�[?9!��:�*����m�ǘ�>FIP>��>��Kg>���>�
�,'�<�پ�� ?��?AA�?�W?�}�g�ѿ�`��=���޺�ĉ>���=��f>�+���@ >��w=�"�;�4�<��>�>ZRa>s�n>f�\>6T>y�u> ]��AV%��樂�|����?������/zg��J��r��6��T��eUľl����_���Ӱ�^�:�E��a���s�}�!>�6?J�>Zɭ>�W>��>�Z��y;羡�n�k�:�2־#�$��X�����ا��(�&�:9s="���V�q?����>��*��=Q^�>�kO��W��?�>G��>�;q>��Y>T�T> �'>h��=i:�>�%�>6�>��=Rz�>��=NF����l�=����τ����?X>��h���2���4#��ԾK�<���=>�?�Z��Y^V�A�h�0��>���J:>y>�AL�q���>�.)>��m��o�:�~��	���3ؽ��>Y��=�}>��`�����;nSq>���	�!>z�=K��>�"?,�3?�|=s��>Zh�>�K�>)��>[L�=�mv>��?#!�>�)?UX?���>��=�Ǽ�����e`�=�����@����߽�@:<��(�	�_�M�=�\�=�ڴ=�c�>PX�>�K�:_�f�p�=�0>��?��T?aF�>�x>��`��M:���B�T�F����=����_U?�\?@�?�J�>�A��l�N>��g>����@��ܢ>�U9>��8��E�� ,���	?�+!>�?�^?(>h��|�k��=3^�==��>��>w/6?@�>{�=��>|X�Qp��t@�'�:�|�����=���=!\���R�=ـ��6�J:�7o�~);��H>F$�>�~�=~;�>?��>;��>��s>w�M��?��g���y�=�`��;C�R�bA�=�⭽n&��[�z<�&�is�2�h�4���Q�7�3�\�-[?\?(tӽ	���������̾�ш�N:�>ZM�>@�>���>Y@1=�����l@��A���2��Q�>g?a��>��������d���ܼ׭�>��>�߈= ��<�+������7��z�>H��>��>z�B<ٚW�A������� ?M��=?\߽s�?�J}?��m��Gξ�� �U��Ŀ1��ǽ����2�l�����Ͼ@����`6�"Х����=�%�>���?'�R�M���������5������7`>���OX>�j�>-g�ǾҏJ��e�������B���{>P:=E\>��?�Y�>�=?z��>i,?��!�q#�>3��>��	?�f!?g�%?�o�>���>Oݣ>�|�>F�>�Z��xͽ����%�=O`��t>�|>��J>x^�=<�k=��6=*s��/='�=�s<i�;�[�+J=��*��.>�v?}�?h�<<6�=� �����>�?f>��<�ό��b;$CJ�6��<N';><��>�o�>�+��,���þ���U�W<@?��F?�}9?��΂>��{�m�$�����>�]�=ܽ{�ޕ�k�ž/Ǿ�v�>��>��n��*y>i�i?��;?k�6?D ?w��X�����]�ߍA�"�h>�J>쥽r�>�=�>o=$����`.��!�t�A=Ľ��"���<.�$���n>46>�+�Y�Q>=��<(��%�f��|�=�x����W>UK�>2��>�tT>%�<��P�kU���N?��#����E���M���S�>Gub>Q��>��9��>�S���;x������?���|>���?3��?��/?K������>�=1�	>+�|>��=v�Q����=���=&��=ٍ&�r���*��\H�i�&��Ɋ>�sS���|ξ����JĿF^U��W����ξ���ⒾF�Q�F$5�[�Ž5��<�x�N��G���uS�����'�W�Nw��S>�L񹾺	�?��?1��=H�[��O%���ܦ��?�=�%��弿�׾`e������㾯&羲�	��ԾT���22��؛>�Y�DP��=�|���(��6���?>�P/?�!ƾR*���x��zf=!G%>�(�<� ﾔ����{��?�
��6W?��9?��������߽g>�?�/�>��%>�������Z�>�$4?q6-?�����+��{ל��=�? ��?�J@?�>��K@�v"
��� ��W?�?��>򃉾� ׾�E ��� ?F-?�ϧ>� ��ڀ��D��k�>�X?��K�e�Q>Cp�>0.�>e�Ľ�����z��>��>�_m����v��AM�3S�=ع�>|Z>w[p�dV����>��վSE��63���<�ؽ��=6t�>��Ҿ�O#>��	>���=�*�E���\����*SW?"q�?#(U?�$)?�����D��^@ݽ��=��>rw�>�12=����>M��>n.Ǿ��c���
���?���?:��?�"e?��L�L=ۿ�.��+ ����Ⱦg!>��">10>��y�{]<��(��\i�nf�<[+C�3�>ۅ�=u/=,P>g��>��>���!�����!m���M��c�Ti	��a��Y�cX���6���žh���gqm��+W�9IĽ����F��ZyU=���7r>$M ?7�)?��>;��=�!�>�,��ξ��ɽ����7��n���!����A�����9/��t|�q���v����>�o��BS>[��>z(><>��>�fk>��=�]c>��+=��>���=$��>h��>�B6>:Z�=��>��>�똿�(���8o����>�[T���?�{;D{U�����\��ec��'>��U>y'�>ؽ��MW���u,�i)�>�t�H�&�w �=�GM�+P�<���>�0>\��b��=���j9�����ӗ>8:�>-�_�ڇҾ2��M4�=5�>I�Ⱦ�k->d�>�"#?��T?��^?�R:>���>�{�>P�H>�f&>h
ۼ��ӻ�>␸>��?RJ?��7?��d=��ƾ@�=�:�$�����<�Q�\�7<�sͽk+���#�ݑ'>�W!>� x>~?>��>R�G�.��<�p�>Zc?$�H?K� ?;� ?�9Y�fu��1p�``j�\!彺݃�Qq?%�0?�0E?Ѹ?T�=� �=�U�=O�#���4�2ܦ>�/�=�RP�V�N������>�Q�>�B9?:a�>{> �R�n��������>�=U�<?�l�>uX�.���L,��)���"�)�[<���=F��=�K����Ƚ<+���ө�O.��� (����L�=�$�>�m?��>ʅ�>�p�>,b>�������<�~R<��e=��*�/�z>P�=l�<�A=^�ѽjZ�=�q�����;���=�|'��n��ɫ��=?�?��+4���X~�)<��ox��F�>T��> X�>)�>���;'����K�7�4�?�;�Kn�>p�Z?
��>��-��?=�����<N��>*�>�r�=���xH�����JҞ�mԾ>~?2��>���m�i��Xl�c���>��=�)�F1�?$$n?� r�\���m!�j�}�D�@dh>��T���B�k�GǾ��g��.���z���H<�i�>tū?e�.�<x��Ӿ���6��"D��>o��>�>��?ц>�qh�����5߾!�~�o����}̽)��=��&>�E?��>��L?x@?$?5?E�����>y�:>�S�>b��>N�>VL+>K4�>z�ŽW�&>6�^>ڋ�=�5i�п[���n�:��<ľ>�H>Ճ�=�m�;z�M=�c:>��ܻ4Hd�/��<@�=^r{�	��=$.�>z�^>=?�?�'�z��<�J��y����& > g#>��4>�ʼ	:;ݟR�;�>���>��L?>"r>�ԩ�Gݳ����B1 �� ����5?�}?x:+?��ƻ�э>�`޾��Ž�|���Z4��[�,^��E.��L�Q+Ǿ��*>�v�>e�=�|>��?e�f?4"?lE�=��\��}���N�m��������$>��?�l!?>!>xO��$;��s0���a�UV������S�=��=�I>�1;>H=-�>[(�=����'+���U<��c�}��>(��>M�>!��=#�a>n$��U����+?�$��t?����.�&�O>��=��l=�J>���>S��=KÅ��Y��t3��>�E�?�l�?��Q?�f9�6A=�?
>�lD�ð7>�
��3�<'�H�[�=�.>12<��E�=���=<t�>���=4>�!2��vǾ��ƽu췿��L��x��]�#�����?��|����=d�;��}���$��*�3�e+���a%���==~Ň��?�	�;�g�?$W�?=7��FH��7��Ӿ=��ذ��.>�:�w���¾Bb��Ex���u߾� ��f.�u
 �?4�>R�S�pr��|*{�̒-�א;�C2>�M1?��ľiL��3���&=!>��<��a���|�����yfT?�r8?�O�y�꾸�ս�=>"/?���>�;>Yɟ�A�罾?�>�o/?F�'?��k�w��Ѣ��M�&�j��?��?��>?o�K��aU�/�o8Ⱦ5z�>��>Vr&?���Ӵ��2O�<�r�>	��>�a�>����=r��F<�H��>$�B?�}X�&�*>��,?�t�>޹#���󾅘�;[b�����P:�>D�Ӵ���!��,����=��>�I,=�%,�S���֌�>u���\nM�`2W�w�	�]��m����^�>C-���>ߙ>��e���9����������O��@??p�?&ID?�9:?�c��3p�g&�=�=$�;>�k�>�񨼴dw���>���>u�Ǿ������a5?���?j�?C�=?��w�G�ݿ#?���6Ѿ�8۾u��=��=���>vs���=��E=�<�=w��=�"=�M>�I>��>�ڸ>&��>���>����]%#�����c����gB��}	�D���jF� ����V�=eɾ0`��`��܈2��{b��2_��t����^�޽:O>�?��?G?��>�k�>޶M��9�����=񷾔Jþ���,�Ȝ龿������t���\7�Ӕ�������>y���;4>[8?@�=�<�=�ec>��;>4�i>p}�>��e=�<>��=�>��>���>z�5>���>	ծ=�Ñ�
d��[��c<>�����k?�Ծ�F��s#��J�+}ǽ��g>|m=Z��>�ξ����u@�[ �>��ֽ�2|���>����P����>�e�>H*~��04����a�7��J��ý=�}�>{�c=��m�׻=�>��پakC>/?>P�N?�uj?�f?�F=}؉>��I>~��=��>걚<k�#>X�#>�@5>�h%?l�.?�&?)J�=�Ŕ��9>��=��%����@�н/�<�/׽�wS=��=��$>y�9>�Ø��!>Ɍ���=>�]���O?>�d?t�A?mN$?���>6���*��I2��A1�m纽��V�� 9?�>>_��>�?U?p���f��'P澘/�����>]�Y>�KM�	H��Ӈ���k�>�q>�-�>��?6��=/=����J�=͡�>��1>7�?N%�>L�Y���=u��%��Ud;��7*�ۄ=�5->4G>8^R��EW��n���=_�I>h�=�,ؼ�^�<w��>���>9�
?��>O�>rEZ>Q?����u=�	>�Q�=�M���=�~=���=�b�����^<��߽r >��#>�������&�=�Z�?9��>���;=f�T����0`5��r>c��>���>́�>�^�=����>��88��f�� ?�Z?�)�>�,�2���(|2=��=�2�> {L>�>04>�r�R���x����D<��>n]�>w~��Лa�����S	��?�s�=7p,�p#�?rh?_C��c������'��[��.���`"�=V�i1�Z����D����eQ��7$>;}�>M�?�𒾲C~�tɾB��Q(�����8>e��E�>�+>I����,�7&��kp���e��QY�.o⼈R�=�ō>Mj?>#?��i?�1 ?��?R�F�LN�>�=���>�h?I�>D_?!
�>�B=~u�>���=7g=8I���-�����=��#��=0�,>��A>w�0=vƁ��&I=vf= V<)��<r�ټ��r��{۽�)=�.P>l�V>�r?I�?[���'=g�E�ɯE�}I�=v�>=�s<�o��w�����;J�%>ۣ>��?��?�(���� ƾ���z��=XR1?��[?�L?��b�6��>i3�p�,�>x���>z�S><��4���:�c0j���>�ʷ>��A;�́>�q?�mm?#�8?{{�=��h�%�����<�%��N���>���>��>S�>)I��pq�F,p�G;�{���*(��k=�G?>���>��Q>޸�;�n�=�_�=01���|�)q>����ͅ=�Ӂ>@u�>4Ǖ�e�6�F�׽��Ѿ�?�4ȼG��F�=�����z~m=:����>h�?o���e䌿����R4�W��>��?���?2-]?��(o�=^	=0�9�c��=�n��|�*TL�g<�=)��<]�.���Ǿ;5W��>∹>�>�֛�#��$���\G��g��x�L��,��`���m��LG����� d���2Q= *�=��ݾm����)�̟�Ce��v��v;<��6��v���?1e�?Ѯ
>w�"��lN�1�������x�<^��=�a�^鿣��� �� ������9�+��U�Ҿ!q�>�IW�a����y���'��!����8>ލ/?3J¾�P�����oJ=V,>j*�<:&��ۉ�󠘿ʰ���Q?�Z9?c����2ҽ_y>��?��>d�0>�˟�ȋ�b[�>�>3?Ħ/?$�������ˌ�ܜ�tZ�?���?�H:?N䀾�3�T�#���)?`��>]�?���������?�??_��>���`>����
�,>�>e�^?�,�`c>>X��>�\�>��9Ѽ�R��8� �����=��Z���	��Je�H+X���=$��>W�D>�գ����� ��>�?�N�T{H�����N��%�<v?�,󾞄>��h>S�>^�(�����ȉ��a�L?��?F]S?DN8?#��ԁ�Jȧ��$�=e��>��>萯=�h�t�>k �>�T�U<r����?�4�?k��?bZ?(om��ؿ�z��1oľ=n˾��{<.w=�ʔ>Z�}<���=��<f��=U%/=(��䃲>��>�(�>��>�v�>�l�>|�����$�Dy��`��("K�U���~�[�Ὗ���s|:���	�#��'���;���.�~�{�	7ͽZN�3Q��'	.>V;	?z�$?IԻ>�B�>�H�>�����.��
꾲��el-�-�(�>��8����|�e������s�����3�"?���=X�7>��>K�/<���=U��>	�>�>}��=��>���=ay> �<Z��>*\�>Z.q>k�>�b�>��t��H��^L��>M�h�C"O?�Ң=|����|J��:�g�W��X>~徽4�>��$����8+�B��>"����<��~>�oŽsE��R� ?��\>T�n�k��wQ�k�w������Y>�=�[�����o�q���p�@F�>������>�;>&+?�L?��S?������>���>�f�>Dm>���<}Ϸ���<�r>�+/?/�B?s�6?E֬��
���}O������,����b==����� 轨)��dh����>��=����n�<���>����
w���=\� ?�@L?��?�'�>�P�<�]^�:t��sܾj~��q^��V)?@U?��U?��?��(?�H>U�s��.ʾ�߾s��>�aE>�lc��G���ٽ�d�>�5L>��?L.?��;~K��?�R�����>�ۤ>�>2!s>��h>}�Q[���a����
̼?���>��.>�U!���>Yʉ��(=����f�=���>���>�?�X;?��>>��>��s>Ƶ8����=(�2=q��=>�Ӽ|ؗ������։=��½�{�<��1=)�����W��=����!�~�߼q\�o?�,?)_���_��@]��3o�f�Ѿ͏�>m�?�^�>{j�>S�̽Vk�]T^�JA<�h_��?�yC??��>Bx彏6�;�|>��<u�>?9�>�P/��5�=�iL��^���5�=͹>i�
?_�>V�M\!�ER�������>�Y>����?��m?�پ����Ӣ"���V"�ȍ�PT��9�9&z����be�0վ��޶뾒��=�>�ˡ?"��<��|=SdO��u��៍�V��e�`4]�<��>$u�>% v�(�{�@J^��J㾻G�wx���*>���<�]�>�?�G	?I��?�:?��(?�s�BN?;�@>޶�>b��>���>�n?��>0Sb>��T>�6=,ӕ=�*������,�=��7�cl>sIR>�:�=,Xl=�x>��$=e��=(��=U9=��<�n�=+]�=i`=7�=L?>�?6?�����L>4pF��c��Җ=(�N>��.:�����=�K*O�m�=^��>{�>�p>�t����`���|�~��<7#?1�W?���>���Ku�>&��a�o�%�=�.�>4�<𤤾�P�d2-��;����>�r�>�,[>��t>�gu?(`?,'?t�P<�kA�s���A��ڽם���E�>�b�>�V�>����`���]��)B�PB�Zr��%0��>Y��=�%�<F�*>�~�=�W=&��77�� z]���=r�=�?��?ۋ?->ǵP=�U������C?Ő�R������߾5*�j1�=�.>+=��	W?JZ彅~�{���A>�b�>���?��?�B_?�d���ͽ� g>�0[> �>�M�U'$��߸����p�5>fC~=��c�E ��Yd=K> "M>����v��v�澒F^�[y���m4�[���.�۾Vp���4��|���B3�p]=8->�K���RE�ɞ������=	];B�k��C�)^p��J�?x��?��>�Y�C�I����9���<�l4��i���+$������2��C#�r��� 7X���gX9�=Z%�A��>��V��⑿�|�)��"{�\�>>�X.?	�ž�ɴ�٩��c=��">8�<G��Ь���j����l0W?�K9?��뾝}��vp⽚X>$ ?��>%>
J����>_�2?1�,?��޼[2L��{錼W�?�Y�?W@O?�� �ߊ<���$�r��-(?�%�>�o>�mD�<�W��|��Q�>�t?�b�>��M~�9������>�%>?)r7���	>���>3�>!5ܽ���6f�<�zj�ٕ�}�=o��G�
�#����i���=@q>y".>/�Ͻ�,��I=�>_}ž@0E�\�B�m� �C�
�2g~<^�>!�¾{>�s>_	>z�+���_䈿�I����J?��? �<?��@?�I��p��܏��g�����>/��>�ל=h5=_��>]q�>��ؾP#I�Fv�_.?@��?�>�?��W?�u��"ӿ ������c��~�=U��=��>�6���� =�έ�%c�,�>�=;V�>�Y�=C�,>�a?>.^�>@��>�ڄ�N>&�2���:Ѕ���B�"�������?�R���t?��'�+��U���x��g��<�	�� �7�(�ɽaK㽁���%ٽ�>��?b*!?<	
?�6>�A�>Zk+�iG
��[e������	�x�
�{���:�����������h��_�·Ӿ`��>�^3�_w>I��>�<>WOJ=O��>Ny�>�3�=��4>�s�<?��=���=dۈ>��>�e�>�0F>���>�>`>�ә�O~r��jn�߫=,v0�v��?��=rﺾ-/�\��"��/�>�9�>��9=f(��X����@��ǡ>�9.�K]�=�>->����i�F�>�g�>����1�I�_���J������h�>.[�=yO=���m蟾���>!���P�Q>���>eA?�X?��S?Y�w=���>�C�>M5�>.y>��=G��'M>e�?R?�:8?��?o��=ŗ��@_x<ybY������g���KD��3->C�8�d�ϽӚ��~ٽ6�U>�Iy�kA>`̸=D�B�x{�<��>�v�>�C?+�1?t|�>v��=!wF��an���D��9�<�}3?`�?0.I?�%?��)?�B|>�Z���߾Y;��O�>� >�O)��K`���v�>��;>�"�>�>ˇ<)�?����PI�$<�>cӘ>p��>⛗>�>�%!>�y�k���&�e��F���^��r�=��=P)>,���t_��=_(e���t>�$=PǶ>���>�=�>��>��>3#E>Ŷi�=w�;��<�d���=C&=��|=B��К�����.������u��y!�إ�;Xl��?��?�Q��_*�%�Ӿ[虾%��M��>�L?4ƹ>ė�>^x��K"۾�b�{ A�痿��?��T?�X�>���x�A<��X;=o��>��>���<
S=����������=�2">���>�˻>����;]�4eX�s�3����>Y*�=6��C2�?��x?|����ɾ�b����J��~À�ʏV�)*��ν\����0��S׾�[3��Ջ���#>K+�>�a�?��N����=�*a�R#���+��\I��1���Ԅ=r3�>��>b�+= ���
�q�ܾ�d��x|�1��=*��=�}�>�&!?O`?z�e?��?�T0?p���"?��>�.�>[��>��>�O�>l��>���>ݑ>8�=��h�&�f+����J�t���">@o>l�Ž��;b��=�m����>V#I�r�|=��=��=���=
��XH�=�Տ>r?-�?R��<̠@>'���pT����=�f>�7���<�΄�����d�->$#�>!?nCt>Kc�����i��H������:?��[?� 9?E��<�v�>�꾫Ѽ�q3	>h�>od>>�;�<��׾i����>��>YH�>�{>�}o?OYK?�:-?�4=:yJ��3��l]G�j!,�!�l=|H�>���>���>P�c�ߜ��<�w�u�29��}c�J�D�!�B>2>�=�O>�>���=(.6�7���v�=��>�E=X��>%P�>L�?��>�2,>����#�]�<?��t��%�hẾ��񾋁���=Te>�6|=��?D"�mgs�������@��d�>%��?2Q�?L�m?�����X��<a>��=�q>�y������<����9����\>���= m������=o�Q>��w>@������(>���E���N��tuJ�\
Q���辺�y��e��֘��P���Kɽ7@ڽ�h��R{���w���ܧ���r�3\�nR[�փ<ަ*��y�?Pө?��?>z�޽m8+��������
=������i<��ٽ�#�g���A������/Y��_���+����ϧ>:x1��}��Zz����-�.��<�R(>k�?-Ⱦ�ꔾ4���x7=�g>���=���;���
�����p�a?�4?�����7���=��?;B�>L��=H֚�
�ν�>~�#?�m!?.����x��'���B��ļ?�y�?d~T?Z�>��!���Y��/����]?��?܆>zu�撺���n�H3]>Q4�>�p>d죾
=���e��؂�>c�	?8n���=�^^>1��>;t=6*�!�Y>]mu��O
�����tb� ?���U�l����I=��>߫�>��� �	����>u辛tN���J�����*���<?!���>�Z>�>�M&�����*G����Խ�J?�ϱ?v�U?R�5?�5���&����=\�>��>��=>L�X �>f��>��,�s�xW��P?[��?��?|"Z?o�c���n��z��9�����=CU�=��^>�h2���@=v��=o���lgR�T��>��>�,�>��>aW>F�>��=b���O�#�蛿�N����L���!��t�.y���P��v���M����e��м8=t�;˭k���:�qu���9t��	�=�?r�3?��$?�l=n��>��Ҿ9�ľ��@���6�5��a�]&Ѿ�킾m,�󐞽�ɽl����.��w��2{>�+������>R�>����ih%=��Y>p8���">��=DΤ=@2B>��>�.>�&0>��^=�����De>��U>����ra�������c>yU�����>O�ڽ�
��Ѩ�E���>���>�5?�7�=|�' ���8���e1?��ʾ� y�sR��E�>l��>���>f'?��ͽ�Cc��Ͻ�ڽD�X>O`>�����9�<6>վ>���T�>�?����D��(���� ?��e?1G?�>�`?�Y�>��x؁>o>m<�=��>&0R? �?nP?8g.?��=��2�[�ڼ���<�4�~D	�H�Ľ�ӽ��V�h��f��/2U�o0I���C�bw>B�=B�l=��>)�1����>̵ ?�Q�>u�?ܶ���O��e{���<%�>����I?�}?��X<!?�'�>�#>g���㍾��{�{��>�G>�W-�X�t�|?�����;ƃ>��)?��b?�ŝ>����{u>G�>�>>h�>v#?:?�!,>�|�w���jӿ�	$���!��C�����A��;.=�/N�E�=�b�-�8 ���|�<��\>G�>��p>OE>�>3>:u�>��G>t��=^�=EҠ;��;`�F��-M=���3J<�P�҅����żߎ���,����J�E ?�]0��ڼ3�#?���>	 <=���]�g�q�"�(�kU?4j?�!?���=�u>淾R�~���6��y=���>k�=?<�?Pjk��W>�@F>�+">Ģ?z��>�;#=��t���f�K��'�=5E�>dU�>8
7��qX�e�H��J
�yԜ>�R�=�\����?�n\?���{�T�����dF����~�>���=�����:���G���Q��������2̽r�=�j�>�@�?��!D>����������&b���h>3�=�2I?��>��O��}���R����x�PG�<�=�>�����?��?���>�im?��>�)?X������>�%B>X�X=p�x>C
?0�=�.?���>Q�.?�f��ǫ�8?o�&1^�����>���!7>2�;>6�@>1����B�HVB�*9>=�0�=>�:�=��B>�d>�P�=`P�=�
?��?�MA�z�S-��"B�����:�=^1>��v�U�;��=gr�=<��>��'?<E�>�m><ՋȾd ξa%���R=O�
?��6?���>�f�=1�>��Ѿ���z�u�=�=>�_��ŝ� /�Qߪ�eQX��p>��?>��=��Y>,�^?D�L?W�=?�B*�tz^��"�������<�X���'?3+?��Y�������~;�k�K�W���@<3���ۼ/�,=fh>2��>>r>D^>n���s4��p����I>�+�->��>�x?+L�=��<_﻾�N?�t�����d��0HӾu�Ͻ��Z>h�_>�� �x`?�s"�v�]��p�� �U�&څ>j��?'8�?z�v?��b��h��>濥>�}>����e@��ҡ���ݽ�?~>��4> 5{��N���R���;��>k�˽��Ӿ�Y�����ɿX&�f�C���	������ˋ���������l8b��1��M¾�y���!%�֒���lX>#��h,���۾�D�����?���?V΋�3}���L���־.��T����)�ؗW�4#��X�]��L�]����6+)�n<I�L�0��W:���>�|��T����2���Z���X�>'`>�$i?0R�Nh��2��q��{K�>��D>����^}�[X��B���`fU?�Y?��2骾��0=-�>>��>�w�>B:=>l�ľ����|�>.T7?0�>��<�۰�B��Ӥh�p��?K��?@�S?}����V��3���u��>)Q?�G6?��)���8%=%��>b�E?��>�V�Z�*���}H?r�V?x�9���U>һ+?t�>�r��5���N>%G¾[,½�-�>��c<�R/��tx��s ����=��?�8�>u@ ��&����>D���C�j3�;��πj���<u{	?u����w(>r��>��=�/����t����᩻ӱW?�6�?%LK?e 7?�����#
�x		�i��<��o>�z�>h�=Q+ܽIn�>~�>�pԾ�Ex�����	?���?���?��O?q�h�wؿ�����Z���|��#>�4�=�ah>��/�Q�R=:դ<فѼ��<��=[�>m̞>���>�.�>j�0>�/ >����(�A���u���$;�R����	�u�w������]��l,���Cþ:ݽ�-��H�6b+���	��Wy��8⾼:�>�\?�A�>��?�GD>~g�>��f�{��H��[��l	�����ߝ�y���`&�s�о�cP�^���}˾Z��>�BR�-;��Pż>]���c�t�>�� �y#>��>��>P��>���>V+�>Aֆ>�D=��=>/�>��Q�댚��ҟ��U��[t=y�5�p"2?,.��M
��i�;��?
���
�S�?�7?�CO>�U+�7D��|�����.?
��������S��2>��>�t�>o,�>*��<�����������W�>��!>솓=/ٽ�[���'@�u`Q>?r��{�j1T<�@�>�o?�G?*_�73�>u�*?��a>R�>� >�:�=d��>��(?3kL?�P�?�ʻ>�*#=[�B��a켬���G�r� mO��)�;E5���8��ߩ�AE��WW�=�s�=�x��JG�=~����������L�����>��!?���>�k?�ꮾ_7]��z_�0�T�?�>�G��v?��>ќ�>��>�7> �K>�y��Bص�kPh��<�>��>l�\�K�������.=��>sN?�[7?��z=���X:>��>�{�>�?��I?��>��g>��������lӿ\$�"�!��邽+I���;��<�`�M���7�-�����c��<z�\>��>-�p>�E>[�>	?3>�R�>�GG>�τ=��=��;��;��E���M=� �)?G<��P��}��[Ƽ͗�������I��>��3��5ټMR"?���>:V��S��-n�N���h��>�ȶ>S�>Ԉ>���=�7���q�� ��'U�60�>a@Y?cG�>�{���wj>>r�>��>J&�>�3��=����O�G[
����>�h�>�;�>�%�\�Q��y���9����>G�=��m��?1~U?I�<��A���q�Ab&�y�����>G�����=��Z��,��>)p��F��&�A�m��vj>�I�>Г?�>���C>Mr��D4��oS����D��x�=��?><�8?�բ>��O�bo�����}��}f���<�Qf>x��S�>vm?)��>?�?�t?��?���Td,?���=h~S>Y�a>lZ�>�?��0?%ė>���>.�ҽ��>5���n��}پ=w'�=C�$>fo*>�x�>:��_�_��=5m��܊���=���=�5T=<q�Y�l=	W�=4ɝ<�Y?h�,?�+�~=+B+���սvt,���M>�.�>��=��\�>�'=>�V�>��?� �>jEq=�Ֆ���u��b�l�7>W�R?�('?��?m�u<�l�:����ᨾM�	>h�A>[4��q>��?_�/��g7����,>�<R>�(��>S�m?G<1?9�;?��*��pT��2���Q���r@�����|�#?m??��Ω�_����I��}�U�UMʾҙ�=M>��I��V�<�$�>�E�>u�|>�x=��'�$�G��������׾�2��'҂�cР>�S=5rs>P����!��d?�WžI�4�С}���O����.�>�.:>���=��E?�#�=��T�_ِ�@ E���=eǿ?��?�Jn?��˽���*�>�ӻ���a�O>���=e�0�~}����*=�:>���e�_�a�=��S<�'�>��3��*�����>���6�Ϳ�L���S�*���ʾ;���G���Ui>�T���Y�=�	�Ⱦ�>f��E���d=�3=hk��S`p�X4žǧ�[��?��?��8�LCľ��a��о|���T>c�����ؽ�b���JA�3����@���F��z���4E��4�Qg���?���Dp��<֑��+�Ⱥ>
\w>Xh?a���>�j=�����(?��>R����偿�S����3��?�:?M��������Ib=��Q>;��>L�?P�>W��ᖾu��>��F?�=?w�_5��"{�^).�t�?i�?�X?N,���C�X�	�;�E��>϶-?�1?.	�.`���>�=(��>9�]?l�>1�7�_(t������&?��J?RX^��/R>�$??��>����]WJ���뾤-����>$�N>����e]��t��Z�#����>���>6�'�(�����>�ؾ��E��Z'�����|�sT�'�?*�����=MÚ>1��=�RI�������ؓ~:V�O?���?��L?�5?�����V�m�N�t�[�J>U��>?��=s����>6�?7��d�p��b�P��>�2�?z�?UDG? wq�0w�&���ʌ������Y�=�,�=�IP>�E���=���8^/�O�w<��n>�^
?[r�>!��>D1>�H��/�=�����Q'�����Z���F��v�����O��������e]���B��{������tY\<�ZR��N'�Tv߽����偾yW>� �>Ž�>�G?�D�=���=�9K�,����G���p/�J�����ݻ�*Ƭ���?�xS��<��]���z�.v�>��-��y=��?k9��Z�9��>�VB��`�</�>x�;�ȏ>=Ѥ>M�?��4>m�>��>��c>�f@>A������;`�\j�=ֈ��q�?ph%��G��XGs�4�N
>L�>)�4?�	�=�aL�,	������f6?��þ�վ�&ʽ�8=²>Ϲ>x�&?\
>��ľ����9�Ͻ��#>��<zw>��ͼb���C.�w��=֫?4&��7Aڼ4��=��?��?��1?����1?an?�r>=��9>8=�و>A?6f?,oe?v۽>��=�0�#<��=~Ӽ��� ��qA���>���׼�������=G�=b�۷<C�=��|�^��yW�32�;�>�?H�>B."?r	��B�G��c��мB�>(^����>�%�>X�>Ԛ�>a��>���=mp������ �R�3��>�]:>��z�ZȊ�@hj��qq=Ww>:*1?��!?KO��Ľ���=��ݽgJ�>Kͽ>%�N?V�?��=(��'9�#��(�2�����[��=sU�Ŭ��~�<�3�%"����=n2�>q�>,�>!D>�E�=^��=
��>�2>�un=eq8=�<�Y�~XA�o=32��6�E=Ź3�鐞<���(q�����閮��;�K��<�S��>#?�߸>v8��[���S F�&1
�ƏQ�&��>��>��?�_�>��G>�	�4��, ��+�%�>�	Z?`?lk���>�>PG->�a?^`Y=��?����=L��}S�}��U�>{'?}?�>*��L�r����	�;��6�>���=�.��f��?��T?�<T�4/]���$��\���ɾ`oG=e�4���g�W�ջq����ro#��2S���>���>��?��]���x>)��$���2:���B����>�Ø>٣A?l�M>�{޾@AU�.��F\o���+�aM��8p�>$:ž��?P�?8 �>���?��?h�!?wL�^�>e~����b>�-�>���>� !?��)?��>&�?��<�T�=���s��6�<&�=�����7>�me>k��<{$2>upa�Cr=;�;-�>��>��	��,����>��`��A�<�x?sN#?+�)��>��=�h��S����=�>��>Otv�@�ͽ��*>�k�>�?��
>Fq�=���������=%�$?j_m?��>3�轁�u=�&5�7�ʾx�:�Db�wXžK��N���Ⱦ�h��ܼ�>x,>0�\��T�>CR?�uA?6�R?3�n�$lJ�����(������&?y?[�6=����\��E�v�.#n� =澪nE>&6��(���R��C�>,��>#��>�8�=C%��yԽ��a��_���=��uŎ>>���	
?2��=A>�{�.:ž$e?�-�� �,��!�������2�lˤ>Q��<��>�.\?>	>y�`�B<����o���5>�m�?���?^�?��O��g��+e0>��= �W�>DT]>�T>�����c>�>zɝ�\�Dʸ>�k^>�?�>���C�u��'>(��\�ƿ�6*��B9�J6�o"��`?�����h���䙾�� �ԙ�;���m>��5�=���ZK��O���DY��&Ͼf�?Y'�?yΝ�������[����,p��1`���m�N�
��D������Ձ��	Ǿ.6�3R#�·.��5�>�Mݾ�ũ��X��|+���7>��H>�x?�����B�>�?� �}=���>G�~=�W�����	ӟ���w�#?v]?9��:�%��j�=��_=�>�c\?��M>�q⾵�ݽ��>��a?h�+?f����W���8�����=���?�B�?�LG?m��@0�G)�����A�> �E?:�4?-�2�}���j�<C�?��P?���=��L��m������?vG_?,Y<��Bw>�G<?b��>��,����6߇���V���
t"?�h>'��f��ju��������>��>.�����̾>��>�u��>�>�ߍ�`��?9*��U��6	?/�ƾ�ũ=ؽ>�=# &�d�����`�,>=��@?s5�?��B?�M$?h�I�ƾ�H$�� z��=E?F�t=�(;�ϲ?��>�0ľ%���0о�>�#�?t� @ʕ-?uV~�>Gӿ����������=%�=��>>��޽�ɭ=��K=�ɘ�RZ=�l�>���>o>D;x>v�T>Λ<>��.>q�����#��ʤ�3ْ��[B�� ���wg��{	��y�����ȴ���I�������@Г�z�G�_���T>�jq̾�ж>XҰ>l�>��4?�
?>��\�;���t�9"��$��u2��L���K�����ު�H�]�����\�������罾�l>���A7Y=���>��C��@��
T�>���Ϋ=�H^>��>�D>�}>C>zX�=��>'�=���=�CB>����%����O��N8�%��  ?�{���A̾�>�$�S>V>f��>��3?�d<�B�?������c�X?5�~㾎پ�]����6�>Gl�>�<
?U�<�6��V���C��7
0���=��+>�ᵽ�¾}*�O�=+�?����4��>b�'?~G? |1?�|�u��>X�>��q=�!>��M>��.=H�>��=?�[^?�lG?�F�>�y�=�bF��L�;�!��	'��ڢ������	���۽ݏ�������;l�=ƨ</.�=@�ϼ�l����`<h��=,k�>q�?��>?=@���O��.R���=k��>��\��	?%��>"
?�~�>�O�>���;a��ɪ`�O�;���>�>QvO�X O��^I<<eS>|�r>�/?i?'��`a9�-Z,=<��=v�P>��>s&?�i�>��>� ��mӿ�$�;�!�E
P�{�;�<�-�M��Ο7&�-�q���g��<J�\>Z�>��p>�E>��>�<3>�R�>�HG>�ф=�=�9�;P�;��E�<�M=�
�KCG<��P����%Ƽ韗�v����I��>�5:��8ټ�?���>�ٛ=6�T>`����B���O��?���>�Q?Ҟ? ]�>(຾�h羋�&�!
����>�??��?�E����F>e�h=�7�=�� ?w|�>Y��=9�=%\A�E�Ⱦy뙽�Q�>��1?���>�<k�s�-�s�������1>o��<����Ӥ?kph??�3�1���3��U$�l��)]���߽Oo$�ҁ��c����j��m㾋����߽�?�>߽?]��?H��W>�6��#ᚿʝ~�2�f����>B%>�?q�:>gf���l����;6��[�F�R��=�>5��Ї ?ل?Y;l>�y?�?/��>y'��S�>w`.�5^[>�MQ>D.�>O!?@�E?��%>��=������=&�=��Z���k=�*�i��ќr=�S�>�n��^讼o����<�U"��t=��E>N�8>Ӗ(������m ��Q>�?��?Et`<�>(>�&M���=^h>���==m0=j�D;5�:>���=A�>�o?\7�>���=�3ľ�����"�e�>,�?v�>�'?��
>ǜU��4�=���@k���-��pX� ���#����
p�k�>Rn�=+m^�f"�>=@E?#�Q?a�.?�Ǿ��\�ǔy��br�	�>s�=e�?i?�>�ù��0��X���9�>/�u�>$$�6���p��+.�>ѧ>�`�=���l�	���V���=z�q�>��j>~?$�=	Q!>|ꊾ�ܾ{�x?I���s��K���>>F�?n�U��J>��x?������2z����i�^�q>�:�?��?��?�Vྟ�2�(>^�>�p>b�>��ʼD\,�/����2>�)>�=u��+�]Xe=tS�>=��>
���]��ia���(=��ڿ�-��9K�D
 ����\�Ǿ�7��-�Ǿ���������h��P���V���:>z��<�l��^������TԾ�&�?l��?�$7��c��;�w�۾�r#�.~w�Eƾ�e��?��s!z�����jl��k8����w#�$�;��E����>QV���vq��ƪ7��si>��>E�W?:�,�D���-o,<%�O>՝�>8�V�~䋿q��� ���?��? ���+�č"=|>��>�2?2��>Mi����-�2^�>�A?R	?V���F���H��Ʋ�=���?�e�?�B?��η4��q�c���o�>a~2?�V1?�>��$���ox�=��?�Q?��>
�1�Qz���q?
V?����]>P" ?�t�>��[���_6+�Wʾ�#νC?Qi�=g���F[���ྛR��
�?�<�>�諒#J��:?P)�g q��ZY�?\��$ݽhk>�j-?0b�c�ҽEi>ɬ�>�u��~�������� 5��o,?7�?�Y?�p?ř����Q�Ώ�k�A���C���>7�=3.����?�i5?c����^྾�h�>Ѕ�?�M�?��?,p����ӿc䚿�Υ�%%��b�>�>%l>r��ݗf=[�+�~XR�漄��>\c�>�?�>	؇>�<>Ħ>jo >v����'�Q뚿L��+w:���������^�6X�Jʄ�1��3�-�˾�3�"ٹ��X��A
L��W,����1��5��>���>
P�>kpT?�5�>(Ȕ>{��Q�+�
W��I9�;DR�{v-�5V��k���t߽F����k׽$�|�&Vc��5����>4�r�%H�J�>BHE�`{M=�|>1�ϻC�>swX>�C��A>�<>���=oe�=m5�=�@�=f�=���>�f��pɡ��M�E@>Ӧ�d?��̾O爾]��Ó��ak>˜�>��0?h��=ɋ-�%㧿�R��y&?^�Za��=�龻�J>I��>Qrw�yy�>�9"�~x��������4��'>��<U-��5��6Kz�����SP�=�L�>��;�!^�׉�>�&�>|[?B�M?.׺<�{?�f�>���>.�*<g��=�^6>�b�>Z�?�c?�`?^��>�=�]��O=f�=�K�gy˻hG���)y����/=!ܽ�=x�ͼq��q]�=B�9�y�<9�y<�=�?�V?	
�>���>�J���>�q�E��_V>De�>�"�=�t?�I�>1;�>Ϧ�>��v>�:�(�i��j�T6�.&�>�*3>��~���?�Sqj<�/!>���> �5?Y?����������;o@>��>6k�>��J?9?LF�=	��������T�����<;=��=�FW�I����.;�E	�:ƽ�޽=c�b>�T�>0�l>�3>�=>�>��>X�1>�T=s�=:Ȋ��Y������;�=��=��<���s`<��=e��!�w�D�5�.��,��M=�Z?�;�>2(=��h>�&����2�N�E�'�?��	?��?Up?�͇>������+�I��!���>�>?'��>m��L�>��T��g��(?�y
?�E�����7��;�m����f�>Y#?r�>�j�Ko�>Ր���3��ل>�E�=^P��A�?��T?n�7�>�b�Wn�O�+�%3�A3�=�������J(��2i��꼾���cw���>5��>E	�?9�)s鼼��k��g�|Z�<�?�>>�p>�;?���>j���6������ľ��S��H$>:�L>�پ���>>?r�>�5n?�?;?_Q�>�/��&�>yE��ܼ�>Z�>��>� G?;De>J��>��='�<�f��ľ�(G�-n�=d��=CA�=8nt>�ͼ�<�<���=��/=u8S=��>��>�=�g�<��:M����>R\?�/,?���<�r=NL/=�3������>��)>�����G��=�c	>��>�)?�YU>����E����7	�'�=�4*?Y�?���>��=">����t���=�1o��r����۾���i\�h|/�_��>C@Q> �?W�> �W?Nv,?��>�M���0�I��oľR�=��^��6�> �> st>�O���c/�������d�
�-�4�>V� ���<�լ=1G�<l�H>�`�>��<us�=Ċҽ��S�����l���\{>��>�0�>�=�1$>�i������`X?iG�������=,@�I ��N ?fK�>Mo>�F}?��>�vn�e��>;���D= ��?o��?>+�?1�����Q�X>k>�	�>DQ�>\%[=0+	��.�=o5��H��>W4q>q%��US_��S�=���=�Y�>�Ȼ�'���ાS����ʿK~&�g��?���౾'վI�������_�k�ܽ��˾�C8�y8���<��f=���̾����'*�W��?h��?	o[���Z��b`�����C�4B���\��y���䀾aa��-��섽�)#�A$ؾ���(��#*��e�>�����.���K��r��M��=��� ?j����6��M���>�I?�ѽ���Θ��Ś��b�IH?	�1?��$���
��=k>~���@��>�K?���=�)���L��/J�=2 s?Q�?֌���5����}��j�Z��?>��?><C?Y�%��)��K�G6�P�U>N��=� ?QJ��9U�^�3>/gN?C�H?��1?������O�U�/>bz?%�'��*�=��?�0�>�!���p��(آ�9(�����@�~>"�a>�.~��R;��h�>��>�m><�=�����?�+��JM�*���� b�>��>>(�>����n����gp>���>8��2��/"����-�~.!?�!�?_O?�F?�����]&���=b�>7 >�>��S>�
���v>�:?�'������v���]K?�?W�?U�K?�o�\ڿ�P��Y�Z��j��0S��o�ս��5�S��>1�\>����
����=L��>��>+Ô>�	:>ӹ�=��N>T�����%��靿�ы��p����O]*��ؾ�T�l��x�/�����Vʾ?����LU=?m/��Ľ
���c�b�=��?|��>�q ?��]>���>"׽�Y���uF�����yq������I^1���ﾵ!��Ft�Y>���l�l6��T�1?������e>��>�V_<��=�`�>%��=fq�<�z4>��<>�ϟ>(]>D�W>�I>��>.�>PRJ>���>�ܜ��0���pK��������� ?��=�0��9��8�辢v-�猍>Q��>Z.>A+��֜������?�u,�L̐���^=�)��Y��>Ǎ}>�5�=R0�V��Z�/��C�<��=1\D>�>8�ޥ�V�5�(�;�n�>��׾;��=�w>n)?D\u?��4?�=���>c�[>���>��=�A>SR<>:��>�??o9?LB2?��>���=փ^���<>��=+�L�U�^���>Ua��� �ċ<���M]�<��`=�6�<Q�=dVu=�����D@<<�<%��>��)?I��>/�>���)1�1{L��'���>a9��b�>к>�:�>u�>[��>eyk>-�w�}����vؾ��>T�I>z�g�|vf��ݽm�\>�#?>sKE?K3?#����'��j�8�Ǽ)[�>��?o�5?���>��*>�"�.�
����S��ac<�����%���4̾R �$ׁ���ֽĊ����ѽ}	>�,?�?�Y�>�IQ>��6>ʰ�>�S�>�}�>a=l�I9+}�>̥��iӑ=A�=�xŽ]������<�H�<*S�=Fx�=�q����<�����;q� �0?7��>����T�k�sLF�r������?�Z>M�=��>Fx�=Q�'�>���E�}���bx?�5�>�u�>�$)�Ԩ'>�?�=
H���W>���=�2f>��=�ğ���̽�1$>kO�>{"?�>(��=+a��a���-�$I�>�l�=4���m�?�Z?�N���e���&��0E�p��ޭ<,�A���d�%Z��'V%��W1�ݾ&��n�N��&�=���>9��?�\��Tk@=��پ�Q�����mm��)��=��=���>�>%2V���t�@��'����2��l�>W׻�-�?_�3?��%?��?��'?�'	?qѼ�$?4j;}A�>�HL>�?"k1?V��>aD���CսbȾ�����������V�`�=��#�g��=9�>��>@��;��b>��=tR=����.����N=�9g=�]>���=i�>�F>;J	?n ?J9���)�uZ�:���Z��<�>��>)ǚ��ki����<q^S>'��>�>?Q^�>�(F=� ۾li������m�=�2?��4?x��>;�<I�h=�&���ۛ�̘~=�#>>�y}��*u�+7供˴�5���`>k@n>)��=��7>Kv�?��P?-_*?	̽t!�m�	����@��b)h=`��>�?�@?v��)�^f{��8��_[E��y��;�>�9=��>Z�g>P4�=�q=��E=�Z��8���ܼ�{>�r>e>�3?�y�>'=�¾|�%�N M?���������=�д�#�j>s�/>�֝> �=���=��=�G������F�N�7?�h�?��?8�?����� ��/#B>Vq���>֙��q��������Y�1>�V�=֑����Xs�<��G׼��3�d�d�.�O����β����9�����eϾ�@7���������R����[�=�	�D�Ӿ.O���0�������Խ{G���L׾�C���2�?�t�?sLݾXȽ��K��]>�m9w�R�����Uz�>����w>2��ν������#���x8���V���F��>鷩�d$��)�_�s�v�!⸾�[�<s��>z��<�KN=Ռ��p�>̦>j�C��&��꓿Ѣ���d?��R?��^�R�Ƚ�u��Ip�=�
~?<?V��>���e\�5 W>\�I?���>�^ὦ
���h� 	��5�?|��?�D?�#��_&��I�j����>�L�>�>�,������z�X=�H?d�?h6�>��#�����7!�ؚ�>��a?)$U��b>�V�>W�>�����fm�E,@=-뵾hA\<�	�>�Hظ@�~���G����d&=��V>-8#=6�������?���9"���b���	H�7O �ۄb=���>g����
;>�0D>֤4�؍��������*��D2?R��?� _?��?� �\�ݾ��?�ػg>��?�M�>L���і��C>��?���1q�����'&?��?���?ںv?� g�Ůɿ�����ꃾO���ŀ>& <>�!>�꽠�>m��=z䂽�=�=�^>�d�>�R]>:y:>*�>�3>t n>a��AD(�!b��������T�|��M�a8��.�������$��"��򍡾t�~�񵧽B�Å7���ý������=�m�= e+?�Kz> ��>m�Z>�&>3m�3u,�J>��F���:��&��bԣ��ĵ�t�L��b�� ����پ�M*;�$��E?��>LT:>1�>	�߼8.N��$+>��=���=�:>�zm>D;�>	�u>Oĩ>��>� �>G��>��>�>��p�Ł�Q��d�g�2�����Y?8 ��)3��{�8�x�о�ק�7�>>�%�>T�'>�/�����ꉿ��>I�3���5�)9��q�-�h�u>��>��=1��;��$=(��Wx��r= P�>ɽ�=F�`��d��UH�/k����>{*ᾃ{>(Y>�#?v�b?�*,?<4=�z>��> pO>�-���t>.$�>1��>h�&?"�6?�
?���>DJ�=�a�W�����&=�rV�0�[���ؽ�3����<��<��}���<x��<�-ϼʧ=�0q=m�<b�=ɽn=�	?}��>L�>ъ�>�i��-*�2�@��Nξq�۽^/�3ǉ=�Ƈ=Jh�>άD?��?��>G�>�?���읾(�>z�_=�C��Ni�;Q��T=cE?�4M?4}>?&`C>�~�^g��I
p=�t�=l?�>�!?x�z>q�e>?��<�'�`��J��P��(���̴�=����_���:>��x�i�<C�>s��>���>	�L>i`
=1;�;��>Y��>�@ >�c�=���>�;)�SX��7��:���d�&>�>�Eҽ��=aG�t���?X� e��a󢼳�%��.��c?��?�M齞�<7�5�d5Ͼ/b��V��>HN?-LQ>,�b?`�>J���n�x��t�����d�?��?U�>��2�@�s>3��=fқ=�W�>NV�>�A�;������=ꈜ���>��h?���>JX�j���r�<�D��>�>'\|=���.,�?��X?�U�+c��e!��P�hR���D=VR�3+M�ϙ��WU���/����Ӿ ��t�4��=���>a�?ߒ���k�=���T����솿�þ��=G:=��>�>Ep�bĂ�r������W2�i�(=1��>Ug��*�N?!*?�n ?�?6`%?��'?'�N=��>�%νx?���>{5:?/�>WYc=Cl���,�=�@�=Js�g�>��Ԍ��=n���-4�=׷�=¾@>F̻G!=><�Z=��J�+^��ℽv 2=jq=���=��=�@�<ֈ�=��?��>?H>�>1�LI�<=�b� ��=LՉ>D��v�=������H�'.?tie? n(?�[M>T$˾̋׾Ă�oU>'�?�.(?F�?����A'a�l6�'���K��[=JW�>��F���I��Z3��n�%<F�$>�З�;1>gˈ?�=9?� 8?s�%��ܾ�6P��]׾|�����C>@�?�g?�v�>�#���B�����z�lJ�֨�=�����7>2�x=��B>%	�>�=i�=�=��|��6��@�,�ڜ	>�!�>��>��?i��>�F>x���lg"�JQN?����!!�W���$��R�=鏼>?��>��<��?a��T^���6���A���%?ya�?v�?16?xl0=�	���/�>iC�>��>��>������=�z>�;�=S=>�a=�]�� p��3X>_N�>�����r��}���2ѽEe���l)�$y��(>�6ѫ�'�������q4��f��6u6�����#��&.�_H��6x�e5��>��������?Y&�?��z��:@����z�q��n.�=R>-k��~�63 �򫻽ӽ;�!�Ѿ�������WC��/C�K|.����>O������W.��b��� ��zľGf�>;��=�)K��K�x`l>[��>qzѽ��a�ߩ���¾]jR?Vw?"P(�!�оa���e�C?���>�j�>Pľ#�l��s
?#�!?���>��k��Ւ��}p�r��=̂�?"#�?��??.#O�A����uW�Ι?5�?Yb�>�����˾�.��
?��8?�W�>��� ���%����>\:[?KrN�8Kc> ��>}�>�.�5��t�)�戒�8%����7>*���zt�`�g�<@@���=�:�>7#v>z[�u����)�>q~�.�;�_�U���E�Q�1����N�>19����>93>oڽ�=E��l��k��Q���z?Ǌ�?�:Q?h
r?)��f"M���>$�>do1��^?[$}>�k�W?�>{�>?���]��칾��K?���?��?G�d?�#S�9Gӿ����������=�$�=��>>��޽�ɭ=��K=�ʘ��Z=�n�>��>%o>L;x>v�T>ś<>��.>p�����#��ʤ�3ْ��[B�� ���wg��{	��y�����ȴ���S�������8Г�t�G�c��U>���}��)�>�E�>Z��>�?��&���>�r=�ā*�����G��[���B�T�ǃ׾=-��X����B�?�A�����hN���-��>"�9="��=S�>�萼�w$<���>b�t=R7B>n�:>GeU:�i>�ݰ>���>��>nc�>��K>�G�>�J���玿�W���Z.�D�v��%>Δ+?�7��}�4�)�g�p��ۓ�Z<�>��?�ր>��)�Zڂ���!�v�>��ž6����o%���>��>�
�>>rf;>��D� ����pT="9Z>� �>6
�>�&j���̾ﳔ�?�B>�b�>�վ�>w�>�0%?��h?��+? �=�X�>Y>�@}>N�=�CP>�3X>�C�>5:?C�5?�W*?'�>`��=�hh�a6<8US=�^G�lv����3%B����T5�<�wC�P�� 	=Q�<(F�=ϙ�=z�=E%�֗=�n?x�?���>�#2?n�μѩ �q=�4���!�K:� �=Ic�>�L>N�|>^�>Q�?���>-�/>�F��_;��վ>�>J1R�l�|��ʕ���=\� ?T��?y�K?攊>Ė��5"���<��U=g��>�D�>{Y�>0߭>e�K>\�J׿���D� ��ɽ��=�ǜ���K�;a%=���$��:tj��.=�_a>?�r>�DR>3@>x�=�W9>�?kc>	,>Bn>�ǽ��M>��� �<��=�(�˼Sn�=�v�=$v�<��;8�h�]�Q�~��<g/�I��,?p�?t���Q�=�*v�����5�%�?~�>+�=ZS'?��?w���.��It���h���3?5r�?tx�>�ӄ���N>>9�C���U>L�I>�
>'�ۼ.[��#^�������?�EN?>A�Ϩ|�����=�"5�>�R�<7�
��{�?�vC?x����E��1�]�O�p �&�=m��*'e��B���U�?6������P�뒾d�=���>M��?�#�����<lv��ٯ���'���"��N�<�`�<Ä�>P>>�lR�V���r�"��F��x�Z׮<�}�>2p�?7L?�	�>	[s?���>Z?|�;=D�>Y��s�
?�H?[��>;H
>"�����M��=T�a=����pl�#7���>>"���l�1�=3> �=A�^�e�;>Tg>q[�=�J�!Xv��|=I��I��=�*��2+U=�d�=b�?���>�`=/>�"X�	ۿ�����9��6�<<){>�{��飞���1D�>JKC?c9-?�pY>\�����X��7�>Y!?��^?��"?O�>Σ�eTE��b��G�7����>0�N>;��o�`��X����)>�C�>���F1@>Lu�?�k5?�o�>�@s=�+F���!�ʜ��<�վiQ̽r
?�?��>� ��=O����L7s�732�'����{��>Ӿ>yF!>�_�>ay�=U=���?�)�yԨ��H�,g0�ǅe>ʸ�>��?��>�~�=�U~�k�$�K?�����(��S����@��'X>�ii>��<1�<?����F芿pĤ�@���)?���?�,�?>�=?�EýІC���1�9�����Ɇ��-#�AB>�����>Vi;Yh׾�ӂ�:��Y�>N>ʷ�t���Z���m���ֽ�uo��Q>�闾U!A�q�>P�<�p��ά�=�{�=]Ԙ�B���n��P6���)��MR�D=����������v�?��?;DW>�Q����Z�����]#�jË��
������bľ;.���+Ѿ@�NU ������>�P:�/:��m�>m�Ѿ�������`�4��-�>=W����?B�<�U��
=�/���̛=T�a>m&���iz�5��B
����y?!�1?5������1%�݌>ԗ>Nzw>���><7���l�Y�>4|�>�.&?E�J=ȭb����ʽ|�?Iִ?q�I?-l�m2_���!�P{ �&~�>�1?��%?���Ղ���$�
��>6܀?�*G?�̽LHU��0$��>�I�?������>4N? ��=¥ƾ���	Ӧ=3|ľTX���>�㼋b��Sk�=�ö�_��*t�>)�n>���t�Ծ�ԭ>T����h�Of@���"���پ/�V�GU�>����o+>[>����v�E��:x�x\��h��h�$?Һ�?��2?��r?d57�%6R�Z%��=�f�>��>��=�6�q��>*�=B��q��u��'�>?�)�?��?��U?�i#� Kҿ�7���^��nKȾ�n=��=�\(>��𽊬�=�mP=�<�^���B
>뎕>(Xc>�\>wA>�x;>#�!>#��o�"�����o㕿��G�6e!�K)�h?j�M��,6|����,�þ�.Ҿ�ݽ ���Zh����=�
���M{�������iF>��>���>k�>�(>��=3@��n��O������� ��Pھv]ξ�T���/��/�}�\mg�8숾+ŵ�|�	��?U��<���=�>�`���KR=۬�>��=��D>�n+>`�=��b>�g`>ϋ�>� d>�2�>=c>$p�>�򕾋���x�����O�6ұ����=��D?@��=��py��v1����>�C?���>��-����/�	����>�k��:)��\#=1tS>(?�5�>�J>��">�M���6���i����>���>m	�>�N���ľw;x���>�?���=�ww>}�?��k?-�D?��z>:�N>�3�>�r�>�o>�(�K'���\U;�4?�?���?��>m=?��C�<V��=� �� ���u�nSؼ�|˽��-��pq=��#>y�->�l�<g�I���ؽ����;,=�==�>���>��>2�+?'N�۩Ҿ��c����)�O������>r9ѽ��=dT?��>ϼ�>�c>_���N[��>�>��$�@�u����F��=�6?���?�=L?�9�>_g��+V��G��kJ�x)�>9,?�1�>.�|>�;�=���Tҿ!�)�gO��׽A�v<�º<j���Y�c�o�%��WU���=m�>��S>W[z>|*4>��O>��9>���>%�H>���=��>��1(� w���!#=b8 =*"�=-�$�|��gF<��ܽ�]���P��A���9ݽ��$�z?�?KN!�V�)=�\��U��?Ž���>t�>=O�>P-'?�u�>�=پ��T���v���� P?�f�?��>v���6�^>�;�����`>�YB>���< �ŽѾ���ݼ��=+�>��?�>��r���o�j���c�� 9@>r8A=�"
���?G*_?D����)"��G����98"=��ؽ��Z�?ò��� �_�7�qm��C"�4s��3�=N��>���? S����=����P����/���(��5�]=Nc=���>>R?>�:��휾e�/�Ҿ�+P�&�<���>��ž��*?N�%?��>��?�6?�?�/���-�e֝���>sU
?���>��[=r� >x�B��>��,=��S��g�����繽�n��wp=h@x>�.>�jQ�qq=��m;��9ǽ&����*=x}�=:Nt>_�>�V->:�->pL?�>��
��Ϳ==�V=�Ɇ�m`����C�&��=�=`�a蜼�
>̳?VR'?�~�>;���Ή��0�����˾�F>|��>�Z?8E?o�>�(���N'����D�����>�������!���}��=��fhj>nG>#2-��b�=�z�?q�"?���>��=ݷ�0�!�Jkо���b^�=`�>�@&?�g>3L:H��I��F�a��;"��g&�˰���7�=�y+>4#�=_|>.LG=U�=��,=�h �Hd�����i5����>ٲ>{?��4>�n�	���?���s�1?��ԾQ�Ҿ� �Lc'���$�>���>s�_> j?�?�$ ��J}�����48�>��?�A�?W�?Eq5�;�Ͻ1
���d==y�=��=@�*:�����V�y�(�j�ý��/��A><�E�g����>�u=�2�6*R���۽"Pӿx$�֞N>d��6�<��|;i�����+<Gm���xƾ�)�)���@��Y�&�Y����\����)ĝ?��?�3�>�O���'�����*��%�,>W΃�|6�眊�H῾��B��̫�:#��^:�7-����Z�>T���ِ�;�o���"�6�=K��=�|.?!S�d�Ծշ'���j���6> =>D��W����g����q���X?H)O?<Oݾ���.�<�k�>�t�>���>��%>ş��\D7=;��>�?��?���<�9��8�����k=N��?kr�?�H?)���8S����w��G?z	?�|,?��W�K���
��1�>;
�?��O?�~�=�M��%.�~C>���?- V����>��"?���=���"�+ܩ=�K��X�T���>Jzû�P�=+��r������b��>CR�>4�MzϾ���>����}q�Mj��:�B)=iY�=ȴ�>!Ǝ�3_>�6�>��>��(�rݒ���������D?h}�?u�c?>?�N(�h���e`��)>)*?�J�>�^Y�Gpf�^t#>�?�H��%���Ͼ�`?1��?�0�?'�V?�cd���ۿX���9���Qrɾ�Z�=���<�i>�E0��f	>�9�=>�w=�z�=m93>ᖔ>t_>�9K>�>?�>f�">����r ��:��b���Y@��� ������I�m�߾����Z���ܠ�|���������������Z��2$��՘��v��-%�>U#?��>��>��>�z�=�JN���Gk�����?ƾ,ժ�O�㾿�ɾ�벾�⢾^Д�J ��)��P��d)�>D��<�$!>��>���;��A�>�t�E<8�>Q-E>� �>��c>C�>��>-Y�>��>�b�>Y�:���>��b�L�T[=���>�wI?$V������9�]�����j�>|�?��s>0f�z��<�]�S��>�b:��V{��%8��CƽY|g>RT�>�&>��=b�[��K��Ľ�� �nV>�>&���03��̰���v�<w��>eW׾�m�� J�=�`!?]�n?%�9?�L>���>�=��=,)����>i�>���>��?YH?�<1?�?�-=�Z�E�.�F�H�
z���f�v�3���=;@�<�9�=}�}�BЙ;�r�<�|�����<��@=�-�<�]�� ���?���>�Ϛ>t��>5��,�4=R���g�$�cr��4�>�a>�t5?ڽC?��?�Ѭ>�����X����K<�<�>�O�=@2j���{���%�益>\A�>��g?	�X?󢭽������Q�ϴA>��>�C?l?��U>7�>���=jB��^Ͽ�U0�����9�f=���9�� :�>@cO������?> ��=�D>�V>��,=mE)=j*�=�S+>���>��<>��4��k�=
�z=����(?���=)��=�X*��8T�V*��Խ2[���F���o��q�e:�,
�)[h=^�?W<?-��=z�E=�'��zղ�ۈ����>D�u>��>��2?`�m>�|
�Kr���`��(����?P�?�.�>J�����>]-;��=K/L>u->8n�}b��֘����ߠQ��^�>j~(?��>"�ؾ_�{=���j?�Ҟ�>�Ð=N���~�?��P?�d�Y�y��$���W�%?��[=�Y��3����&o�mc+��7�)�9BZ��=�=QM�>�l�?���Fx�=뉝�>��")��ٙҾ��B<�V0��i�>s�.>r���>��		��E������aY=�!�>�h�=��>70?uP?ܼ�?Uv
?�`?a �bQn>����J��>x�>���>l?���>�|�>/�>�&7����!+��|��9�w�h���p�<��1>e�J>�w/��%��<>�V9�i��r�jv���w�죽=��=j�=�f
>�?d��>ҁL�I�3=���y���AF>m�>��=x��=���0�վ� [>w�?��M?�?�>�㛾@�F�-����ł>�uH?#Z?�"?��󟃾EH'�*���z�o	�>컆>��I�Ͼf���l��>�2g>���s
>��?�nA?��D?��>��S�KT7��K(�N.Ⱦ
dG>��>��>�lb>8��{�_��l��c^���9�c��T�־�<�=>�:>04�>&u�<{�'>0��=�l��",��.ܻ�P�=�ʫ>�J�>�Y�>��9>�*ͻb ��4���;?Y�M%�z����i�>��?
�>}�'����>3׺=3�w������R���?���?�?�8?�+(�����Q>XI1>�a>yq*=�i����6=o�[>*O�<G�R>M�馆�r1�=L">���>�Q����ZC�$?R=��ɿ��Ӿ>.>������|�O��%��鶾E5�>8���M���]������X�;������������?���?um�>5�]��./�R�ƾ��=^��`������ �L��('��[�k��y¾�!�$��/���@>5���S�Y�r!X��
K��\�QO�<��)?z׽�᧾H�����=�>>>� ��J���������`Qn�-D?1�?y4�JD��xc�%m���3?��>��Y>�>���� >	��>�bX?;�? Á��M�M�n6>-��? .�?̸<?�ゾ<XZ��������N?��	?�&�>�F^��������*��>g�G?|�>׾��&S��\���>0]g?d�L��4>�n�>�e�>��>������ �kK�Aۄ<��f>e��<�E��*��a����i�=f��>\��> �^��"��a��>q�8VR��mN�x
�
�ԩ==�??�����Ӫ=F?T>��>0#(�Ɗ��ɉ�$��d-L?U�?��S?>�2?�⾥�ھ�g��̓#=�+�>�|�>���=�����>�N�>l��u���0�
?��?��?ۅS?M�q�7�߿/���ܼ�-���sN>)�]>z�>f�_���=�U=����X<�GG>�8�>p=�>3C�>V�u>Y	�=�?>�F���|"�Nꦿt鍿�
a��c�t����y���ȾIq��	�P���P����k$�8́;E�<OȬ���A�XIj�2z��=�=~�"?}6?���=R@�=K�>����Զ��>`v�����������ܡ�FX������%&�>U�0��g�
�M?-&�;�u>�1�>9�
>�֙>�F0>𝞽#1=��Y>��0>�X��R]�>]��>lH>���=Q!��d�<_��=�d��>,y�W�&��K�&��q�>�C�l�����a�*v4�<���@��>�]?��>�7����Zw���>�ր=�<���1��ͭ��b.>p�>���=�,��Sq��Ȍ����NR�<��C>�=x���I�������=B�>�����>3�>̓�>6�]?�X?��=�����>)@�=���=�/�>��>>�0>t��>"aG?�@?�û>뵃=J��k�d��=>���ĩ������<#ܢ�7+�r�>"y>��x>���=�]ν�y�m`k�ǡ�<��>-�?(�K?� ?Ȱ�>u���@:��:a���J=�h�>�3>��Y?p�?���>�?*��>��>�a�:��.þ�Ž>�P>��B��_��U�&=���>�-���J�>mvJ?#�=Ǧ1��f?>��>�+?���>�A?? Ű>��>�����h�U���W2�4���+&��wa����xy��;><6=G����G��/�=��>ե�>| �>�A�>���A�����>wWL>��=G�>��r=���=���ӌ"��<��=������ὄ�=���:mS�����UxX=�d�-5����?�]?�V���<��7Pƾ��LP���>)�>]k?w��>
8����g�:���c��Kc��'�>�?f?k�
?ArH��[�='t=��>�O6>p�K>uy�=����Sr�\�=�k�S=�>!�?4�>�Y��;h�'�j�����]�>޿�=�1��4�?dm�?���A곾�t��D����X�Z������@7�8�=� �)��k�>]#���ξ����S�i>vQ�>��?�g����<���
��E�����G��>�8=�??��$>�$�����؎���Ծ��Q��b=ׇ�>?<)=Y�>p-?l��>��?���>^J�>�aI����>�KռE�>9r?_>�ߖ>�?_J�>к
?��!=�n��zY;�\Ѩ���m�����|=S�>5i>���!��<����d޽��w%=�©=�.��g���CpȽq!=x��=Ό>4�
?�rM?�a#>�F�����>P�����r�U�>�~�>��!��
>�R>t��>��?�k5?�1Z?��3����,���ﾬ�I�pƻ>6\O?ݤ?�O6�՜�>Pڻ���H�'�*���k����*���:����[�mb�>�%�=�ʗ=�p>hp?��4?��B?$��=��S�N�w��׾��c�F� =��?P��>����j ��]H���!�C� �S��<K���I�=c;�=r<�=�н=�C�=_�=��ջ�, >Cjp<��>P� ��>�@�>|�*?�F�>��
��~��T�޾#{L?2����I%��������K>/*�>9���G�>c<&�K������X;�[C�>9�?kZ�?��o?��-�^���Bp>e�>��d>�E�ܖ�����T���`>Y�e>K[P��̺��ͪ<p�Y>�'>�?�� �ؾ #� ����ƿ�L�qc�����e�����,t��e;��l1=�����6LþF��\ҽ8">��Y���FH�6xΆ��?���?m"��ٕ��k�j�澛T7>�7��OW�����Ш��2\����r�	���P����'��[%�բ��O��>��꽀Ӫ�����侬N�>J�=&�S?�ʝ�"5� �+��)�vP�>�fo����;���������=�k?�Ld?P[/�Ĝ,��4A�Z��>�xl?��?��>��Ͼ{y���?PWq?�>5?y��� ��FF�=6��?i�?#�W?���Q`���3�I��	V?1�??�u�>��aQ�J�n��e�>�	?��>�4E�����]��91_?`ȇ?��:��#g>_b5?�/�>U���)T�3�=�����Fҽ!�>�+��{���s���a�̼�J">p��>V��>������~�!?�H�%6��QM���K�WM	?v��1??k�W��p1�=�?e��s�����x�!��Q?�:�?�/�??�!��cdN��e<�}\=�N>��	?����R�-I�>n�#?R�þ+�ʓu�CF?���?f��?�,b?�By�]k޿D��t��.��Wڳ=�C�=��`>�wG���}<q��j��?�˽L��=ɍ>��X>
8d>Z�N>��>9�>,��%�"�0��������<���[Y	��j�������� &	�!������|�"��V�\q�\8� q���Jg�C�̽��%?N<?%����#�=dj�>^򂾓�"�2��)��Ͼr������Ҿ�Ɩ�'���Q�i��/����`�zQ�r?,?�;;�R�>���>*�.��a�=��U>d[�=H�>.�B>*Y�=���>'S>	o>�>f*>Z�ǽ G<�1s>�7���E�B�$����9f��0:�>ݠ�������H|������C�/9>�?��>_�q����t��*��>�	�=2�h=�@�<�H��*��>���>� ʾ�J3��w>S'	�A�����S�l���_Q�����c}�zG@��7�=a��>�E޾��\>N�>@�9? r?R?jߞ=ƚ�>Un>tUi>��[<�ګ>���>n��>�S0?m^G?pN)?��>G؂=�0���`����=''	�)g�<ht����ݽ�������\�g���=�m�;v��;���=[��<w���d��1?#sP?�:�>㩯>����B�0'D��i����>�=j��>��>�B�>�f�>��> a>�����վ~���&?[�8>)�;�vV����U�N�_>[;=��h?�!w?��">߀�Da7>lz�>�Ĝ>��>�f3?���>�G'>�>����V������=�b@}��}�=b����@$�ݓ��EҾ#���7O>�o�>@NO>�#>D��>��X>qP6<���>��1>��������1�<����$寽 B> ��=��a;\�	�����R� �g����<-�'=&�<��N:�ߣ�Kb-?��?g#��ѷ��k#�EjľW�����>\ ?63?���>��<�޾Ds�uv7�|Ϊ����>�D?GP"?�&����=�4�?�<��;>ެ8>��S>��^�T������B���8?���><.�=;�k���C���P��K �ؿ�>66�=��o�Q��?h�s?/���O��u྅�X��Q���=v��=9��$����,���o��+��p¾�`����6=�;h>���?!�����=�ڽb����Wy�ܴ��U�!>)E�(��>Q;->m�:�����Z��������8��K�>.�佟�=�[J??��>���?9�?�D? I%>�G#?���>&�>ͨ�>M;O?.�[?|Dn?�$?*�?0>b�M�w�)�Q��I�L�ސ��X�q1�>�܈>����/л��M=N���iPJ���=�>;�a=�9=���=$��=���=�o?hSF?�1t�K��{�>a���^��H�>#��>�nѽ��<W�=�">���>у!?z�>�<�PľːԾ��6�9� ��5?�D_?���>B�t��3u>	�����Ӿ����e<hB�x�S���¾�}d<f+�=���>pw=>4O��s�>�*v?�63?�
`?@9��L/�Ӄ��t3��<�F�=2�?��{>��#������!��V��z��<-�Ro�=k}_��p>��=��=E�[>#HJ<�c=c*��d�= '��7�ýʬ�zy>41�>mo�>�5w>C!*���o�Ĭ��jT?�P��\�/��_ھ������1>�Y�>u�u>\�ξ�r�>`u>�t��fU���>�DF>���?W�?,?��������&�>݆?N��>����	�� =������)+>���>�3��Q(�!��=��=�bk����=D�����1�z��oϿ�.o�q�Ǿ##�"��i��Q��Z~�=�D�w�Ծ9P��п���3<C��=�"�=��!=R��_P����⾋��?��?Ħ��s�[= �>�C�� ����>��V�DU�����)�=K{���t�h�z�vʾH=�ln=���e[�>es��#ѡ��Z��{� �x�;<�һX��>�Ծ��Ǿܴ!�Ԛ�=���>����
�����$.����M��o?ޛ~?��$��.0��(̾\d>�f?�:�>�?�⪾����n>��6?�S3?����⓿	v���=�I�?� �?AG@?�8C�:y>������(��?m�
?���>����.�ƾM�役�?��5?�)�>������N`�w��>�6\?��U��R>���>꫗>�$�����I�E�3���)�
`$>g����X��]��):��I�=?�>L�q>�0l�+��U~�>���3_O��)I�F�S��^��<��?�H��w��= �k>8>�T'�eӌ������]���K?^��?�`T?�7?Y��@;��[��mg�=M��>`Z�>섲=>�
�pt�>��>��쾷 t���1�?��?ѻ�?�Y?�m��sֿ�l����ηs�o�>k�;��c>56=�T�=��Y>,p�=FT�gGS>bk�>QE�>cf�>��>��=鷼G����v!�L���X���{3���4���(��!���۾�:��%}	�F��峾�=������+O�g�H�čս���{�5=u�J?��?�G��2T>��>pFھ�����e�@���־�z;������������=��mϼk�%�����S�?I�̼��>A�>��
=�9�=��A>C/2=�Ѹ=�>ς*>q�D=�-�=�	p>� =��<..��X��=oB�>�`���j�$%�P�Ծ�_ξs�>�=�1�ӽ�R��}��;<�<L��>e?D3n>V�O�᩿2h��R��>��,>�vb�/벽�_���m�>\��>�R����=	�7=(�i�qŞ<�A>��=r�O���?��{�L��L�=m��>埫�;�(>��x>�C?=Fa?�(? R�=�j�>o U>�+�>���=7� >-�*>;�~>�n?G+?��8?��>�=��o��j�=�o-���gy,���������m�K�# �=�G�����UK=U<{���=b}=m R<�Q����л�k�>.E?Fӭ>��>~K�=}O4�PD���
���>�)E�R^>�ٸ>��I>l_�>���>��>�4޽�~���¾
� ?6�e>iQ��9�߽'X�>5�>؊g?�uk?uF$=.֌���6>J[�>��>ǭ%>�)T?� �>�v�>�>��v�ۿ\�R�y��a��b(��IR=������=T�>���<�3��gc>�e>?���>�=�>��&?6Q	>��Q���>|N->|4->���;�9��s >&�j=,�9=���oD�0[���j�=zؔ=%Wʼ�J��r��F�V5�ꓽ�?�;?:a����r��_>���,?��?ӫ?��>�z�>^�6<hH��u����^6>�y�>��?�?��M�
����޽A�>��>н�=�u2>#$=���������ܼ�0u�>v�?O`*>=���4.�f�;����'�j>7�,>_엾~j�?���?�'����x���T�!�|�^W�������=ˎ���c-�LKe���0�g��#�����=Lm�>ʍ?J����E�w�F�u��4���+�P4d>�Y�<��>4*�>�����A������l�F�C7���G>��g=��>�2!?���>�_X?@�>��?�\=��{?�9U>4��>�c�>g��>t?RR5?̓�>p(�>[A=52$���D���
��=��<ɤ�=ի3>�
>���VN�g"T>��={�S�m!�>C�=_��=�Y:>�v�=��=�i�>a6?T<�Q�/�$��=�����ݽ=|N�>��>T'���3��˒=H�>���>�\F?�i�>s� >��R��;޾ ��J�%���%?|	�>��I>���=��{>����Iq�s�{>�  >$/�� ���<b��Ż�b��>IN�=�����x>�a?�D?�k)?�+>[���~o�8)\��v	>�D>y-�>���>:����:�RI���(�w�_���=�V#�<$`-��#>�b�=��u>��>p3�=%��=�5;�zýߋ^�j>|=�3�߱2>�v�>�+?O�>�L��ͪ�5�����I?D�����=9����ƾ����C>n&@>�ͽr6?z�����|��~���:�VN�>���?�Y�?&g?U
;��t	��F[>��M>��>?� =T1A�lW$�*�����&>��=��x�1���>�4M\>r�~>ڽ�)¾�
�EJ�ɷ�r2L���o�J��Z���c�Q�����=����mM��	�藾���c��v��<^�J=�To�QFӾ�dؾWC�?�?F��=�h��4c4���-���=����=KA���'(���;*:���֬�?[�	z���̭�N�b�a���Z�>�?���>������r�u5�>c�=7�?V]��j����߾���>�m ?����gh�]|���7���¾.�Z?AAR?��5�\�׾Ƌ�Z+>�zg?Q%?��?�F���%�Kۇ>��@?�?�;�S;�򚋿�7'�Բ�?LZ�?(ZT?��N���<����C�B�X?Ur6?��?��X�L@L>��?�-??J8>�.�G|��F�þ��?f��?��b��>�>�n?l!?h�-M�H��2�¾7gĺ<��>j7�=�	��;xھ�%o�mU���?�>$��>-������~��>��˾ĪG�UG������%��1����?�#ؾ��>��v>'9�=v�'��ٍ�Nd��tս��L?F�?�!N?�T5? ��k�K.���g�=p3�>���>�A�=A2ؽ��>�	�> �۾6Uu��? ��?���?���?c0P?f�i���ݿ)r��49��έ�5n�=Μw>���>����w4�N8=g�?�>��]�->i�k>��>=�>2Î>w?^=�c�=M���=�!�*�������C�gz���	�qr�����ŖX�D�h��d�����p��0�����?�vƽCc��F欽�\����(?�?�����Rg<��>�Ϡ�Y�)+�䅨����Svɾ{��m��.������Ž���:�P������6?~��;ٗ>~��>h*�<Ҷ�=!�>z������<�c�>?�}>�
�>��s>��D>��=��=��A��1�=tp'>������k���h6��ki:����>iL��Mܼ$#Y��g#����	)�>gn?�ja>FG�N����򎿦�?6�>ċ��{�Y��%����X>bJ>�uo>��)>}P���6ݾ�a�ti,>f��>3��=�z������}R��\>���>l�����)>�E>j�?�\?2)/?X�=���>Ni>�|>�j�=��3>M3>�s>"v?��+?��%?{'�>ޗ=;c{��p�<!�?=���R)��ɽ_8�7�����A<�TN��)�=u�-=2z�<b�=A�=�k5=�t��e�F��>�nK?�=�>/�>�����O��O>�w׉>�N��u0�>�J�:���>w7i>du>�	?>3q��
f��ߢ�z@�>+��>7�X�<��=���tN>�H�>�>V?�8?�q�>��A����=�n<>�>�>��	?�
?��W>k�Z=P�޲῏���( ���1�d,f=5̒=�𣾌���a���N�U9��n2>��=�>�>�ŷ>i�h>A�>���<_9�>3�v>%��=�,=xZ�=n�S����6�>�z>����MV����=:I:<X�h<�̽���5��-=7����4?�X?7�ν�2F��h���[���'�Mn,? �N?��+?��?�(�=��(�=� � ���R=�B?Ǝ]?Bo�>ݡM����=M�Ž8�m>��?CQ�=H(>5)�=�B�P-���,���-�>�?��>��=����_�?����z>��=�[��m��?���?h�n�Ӿ˧�#�H�s<J���<���W�ٽ`�����{e�	.$�&�;���Fg>P��>v��?��˾� >�-/��������p0���R>P��;�>5��=̬��]��S ᾵���i�����$Ʉ>�玽C8>��)?�B�>n,d?Z?7�?����p�>u��=y''>�??0��>��>fC_?��?��?M�7=�䤾Jn������Y�= �l��<(��>1T_>=�h��
��}�=/�=��<�j�=
f[=��=�\K=�U->�Ǔ��\1���?�h1?�_ʽ��A�/�>&A>�G�U��>nۇ>�΅�/h���͑���>��>,;4?�|�>.��=�@��Sݾ��?�=!�?��?���> ݵ=Z2>���y����8 =��N>�����]���]��3#��WI>[�q>h"�/a>��h?}�*?+_c?D��=bBg������˾�c �e�<��C?�T>�:���6�C羫]���m�����c�=���R�>E=L�=!��>��#>�>��<eA�(� ����R1�=�Lt�YY<>�z2>dh�>^��>@�T�����ݾ��P?Ǻ�U7���߾�u��m�ߋټ̙�>@i�=b�?\u�D�t�%���Y*�.�>"-�?a��?lr?Ǉ��ܽ.>�>�=���=�F{=W���Z%��wdu>�CV>FD�܇P��콽��>�n�>�.����{������sJ�;O��,,;��u��5����p�辎���T'�� ����mb�G����S�#=��=B�=6|=�k��rO*�e�"���?ֈ?^�����>C�.���
�$�����Y�,�^�f�">*���2���rn�X?�'%<�w�߾!�=��2%�N="����>�X��.��
�����:��>�醽��1?�HV�2��xq��@�=YP%?�<�>:�Kk�����0˾�(&?��O?V$1�P|��Ί�M�}?g�B?e�>f��"a�T�?i+a?��>��=����┿B=�?C �?�K?�f����G����w1�.w8?ԍO?`��>�n�e �ZjG=Y��>�>?���>xbQ�����Z) �/9Q?e�?�RG�"�>.8?��!?����J���׽�Ⱦ1�c<.?^I�<$��`���g���2�j)?uW>�u���4��>i�ݾJJ�S#B��� 4#��8<�<?�3ھ��>.�y>7T>��*�)ъ�f������� P?�?�(R?l�6?�����������U��=��>��>���=�Wۤ>�>����x�r�� ���~?��?T�?q_Y?��k��ٿD��S����f���{">1,�>py�>N��F��;bd�=�sǽ8�<�>T>���>/��>À�>Rm�>��E=-��=D�.V$��,��B避m�-������wm����(s�1������Fh5��$n��0��#�J�N��%�Jp��T�X(>���>	�>��>͹/>H�>����{�UY����V��/0���P�C�Ǿs,����q�&�2ڽb"�zN��E3?L$�� �<`��>�q�=n�=j�x>M9����&>�V�>%jK>�X�>��>�F\>��>x��="��l���s>r?��xxD�q�ľ���e྄W���3��W=�b]�e�H����;�t<?r_?6�>KK+����৿�e
?n�>���u��=!ḾDg�=-^�>>��=��
�EM������Z����M�>(!�>�풾(����=����=��>���� �=i>C�?c$a?gf?0>��>�l�>qk�>u�5=���=�-*>�`�>��?I?j�B?���>c�=e�_�FI�<��=�F�����(�لz����	�P=u�J<���=�8�=��I=��=�s>N��=o+�:'��ְ�>�=?�`�>���>Z$ͽe  �u�'��K�H�_>̺=!��>+�>��I>��`>'|�>q�>�����K�i7^�ک�>
�>�#`�z�u������O>���=�"�?M�?0���2���5Q�=�*�>���>�a�>��?6�&?=��>l
�����V�R1���ľXbM=x=�;B�>'�Ծz)�y?�3ñ��sW��r�>IΘ>��>^[�>5�>�e`=�C��J��>w��>P�=�̱=��G=�ǽ`�����=l<==ϖ��������&���ؽ�׽ �<�'���:�<�k0��?.�*?q�Y�W!ݽ�s*>�u�:���ɛ8?30?<��>t�?�F�:����9�dl�Y"�=	B?��m?�
?�pb�Nߗ=�:d����=`A�>�,{>1�=�qĽ��������O�{>�H�>H>c��ϣX�ֲV�����#>�]�=M�:/�?�3�?����ʾ�䟾�7�N<]�gK�=�b�Ϝ�����W��J���Z���O>��>!�?m9t���G=�E~���i��ʄ�āཱིמ>�ѯ=j�>f�A>����H*ξ8͕���ҽ�z=j>��t����>�2?�B�>�nd?Q�>)�?^>�=Yl?���Y��>�@?1Ҷ>O��=��??6? 7?�EL>�`P���L�F(о�B>��	>���=��>>�>y�<���=:|�=�K�<m�g�,jнf��e�=���=���=SZ���L>-�?;,?Bq��t����=KR��O�<-*>4�i>�ڡ�7\C�.���JN">"Y�>��(?���>���=F���xG��	��x��=��?�z?:��>[Kh=�[�=<���֒�'f9=�4>[��G~��Z��6ٙ�+X�.��>Fo>�m˻��>x|h?�`?��?? v��&����������<k�>�B?Da�>|*о2�&�K�J~���>��w$�g�[>L��\u�=���=��~=�~�>���=�Au>Y�h�-uսֵ򼂻;=����uD>���>T
?_^r>�7��W{�����A�V?�lL�@a��C�����n=y��� �>Gɟ>YP[?'� =,V��qs���n�|+�>5=�?���?ͧ�?�f��J&�� c>� c�c�S�Z8�>�mٽZ{J�]a8��y=��1>��2�ɔ����= ?�>���>Ԗ)>]p��3Vd�[�Լ����AZU��%���߾����$����ʾ)��u:��>������q-,��a={��,D=9B������>Ҿp?�ҙ?1N�?Ʒ���n���"��l �";�k�=�đ����w���J�>�N���-M0��2���U���4�Q�D�7�=��|�>��_��Q��݌��0US���?�KU>cHI?p�g��z?�r4C��6>�t�>�
?�eƾv�.���6Fܾ�%?y�D?�A�6|��齾�S6�=ya?2*-?���>e�ܾ�{þ���>��q?��>��J��V����k��K>HG�?N��?�?E?�U���!���8�"���?>`?c�>n��W��>v=��,1?�y,?���=��h�����o��~?4]�?ka`��ڞ>JA?j�?�詽�Y ��1���}p�`]?>`�¾){9�H�����<=���>�PN>��
��榾���>��A�G��J�)Y������<Z�?3��U��=�
d>ț>��!��s���㉿�=���G?X4�?rJR?�8?|��;�Epʽ��=O��>&7�>�o=�	���>��>���ip�^���)�?o�?J�?�9[?��n�HGӿ!��!���������=�$�=�>>��޽Eɭ=��K=�����\=���>���>Ko>�;x>߼T>�<>��.>c���}�#��ʤ�ْ��[B�� ���tvg��{	�ey����	ɴ���֖��@����ϓ�T�G�=��!U>�,!�� ?%�D?>�>�6?�.?'#?񼁾��?��๾,-0��'�Ђ�|ۅ�Z:j��5�=���=a	���J��8�������{?����t�<�L�>T��=��=c'�>ġ�=�&>�2e>#��>�$>��H>�#=wx�>���>^�'>m�>�+�=pK���u��_>L��&Y�9���c�9?������o�a�1�eW����,&>j��>*�>@5+��!��"tq����>;Cu�Ny��׭�[*�[��>�b?�\y=�Q����� u�p�ѼT�=J�>�j�=22���ҾfZ!����=�T�>~��h�>
a޼�t6?��e?��$? +k=>��>֓r>-��> n�>�w�>�qI>�Wp>�J?2 ?��]?]��>��>�n��#z?<���=�"���[�=�Cv�Sq<�٩��~�>^3=��>�G�=�ǈ��Т>+"X>�����=$���qD?U ?�A> �??Cyž��d�Z,t�ZR����>�Vh>*�*?(?�8�>T$?($1?MJe>A�=�þ�%9� Lo>�<>�S_�<�(�����v����<�/?�B3?a�p�A��4�(=x�$=��?~h	?��>�E�>7aս<� ��B�7�տ������7f����`��>�	Ž�r,�}9�>��-�+|���>��?�V�>^!)?��?���>;u�=��>r�=G�<
E>�J����=����4>��9l�J�����C��'v=������L��_b�2�ϻ��
>���3
?ּ?�4����=D3½�پ�;��f��>���>�\�>ǡ�>���=qe�YnP�ihF�"|�#�>�	>?ƌ�>��|��A�=���<=���C=�>��>�ȡ>����˭�����K��=�?>Ծ?�ؗ>!GB�:�s�]��^��~�>���=� ���?��G?�9 ��k�؟�+�G��_��i�>�>���ѽN�$��(�*	��ؤ�{`��?��?��*��>��?[!�u��>�������Ԅ�M@���C>�wL>��?�Q�=��ξ�^��t������@Y�5�O�==!"�d��>~`.?�K�>(hr?��?�3?Z,/��X?&x|>d58?�L�>5?�T? p?$�>э�>�F2>A6�<R)�����w�����=�>�|:>�p�=|�ܼu�&=2�<>QI<Y��<��$=���=��S==��=�V<r:�=kf�=~c�>9+3?KK��1��>־=m��y]پ����>݊>�м��O:<�<Ȝ0?�y<?$��>:�>@i-���U�(>��BM>���>�-�>:�?�S�>�nR>��b����#�<I����%��8y�B��F�iV�<�>>�%>� >��~>{�p?��-?4l"?�捽�"��,b��K$�fl＞ػ�ܮ>��>^�ؼ��dZ2�[a��\R���#��j��܆���=�.>h)>�e�>��>p�U>:b�;�w:�
�񽷅=cR��i�>�
�>�^?{��>��=�)�����n�I?�@��`��K��$Ͼ����>��9>@��EG?��
�F�}���32=���>=�?�G�?|hc?�C��g���]>��V>�>%�:<=�;�ł
�ᔅ�E0>%��=H�y�4��A�;(�]>m1y>m�Ž%�ʾ��{vI�'n���N���8��a���n����5��%�>r����k�m����^��L���&��
��w�l=��ڻ+*���	�����?rc�?��k�jﳽ�_���
����+>���޹���Z��0�־W��<'��k7���k���Z�����I��>�/�kƓ��/��v�n��G$<T>�!.?�\��~�h��_8��jK>4_[>0I���ٔ�>C����6�:�%?vy??��4��S����;�>m��>p�?r��>� X>�ݾn��=)c?dJ?q,�=���ឈ����;zx�?�W�?�TJ?�.��'>F��#��f��f^�>�K�>�`�>���=JG���̾f�
?]eq>�6��>c_�4���#[V����>�ۋ?�q����I>b��>�ŝ>�Q�<ﯛ��<�5U��rf����?>���=� 9���+1��b7>�7�>=y�=ߍ+�-����C�>u �VL�R�H��.���N�<�?ȼ�\9>�h>�1>i�%�|>��2����� ��J?D�?)`S?��8?9�����q�����=L#�>��>�&�=W��
!�>bB�>��㾟)p�[G�<�?�U�?E��?NcZ?�5m�>Gӿ�� ��������=%�=��>>��޽�ɭ=��K=�ɘ�Z=�o�>���>o>C;x>w�T>ϛ<>��.>r�����#��ʤ�4ْ��[B�� ���wg��{	��y�����ȴ���K�������:Г�x�G�]���T>�:?�)��>���>���>v�G?t��>��?V�_��,2�����-ؾ�{2��n���M�Tw��B��<��4��T��#�=5t������>�����=n�>��=O*�=P>r>�}'>��j>(5>�TS>K�>g��>X�a>r��=�+R>��==�:\>P>����]w���12�8�7��@{���9?A/������J�1�l ׾���i�_>BB?x�G>�;,��,��C�t�s��>�bR�f6���yO�����+��>���>��>��;~����������ū=���>�t=�`�='̾��S��A�=�E�>�`��8�>��=Q6?�i?��2?1>D<�>�-]>AՁ>"v�>W��>�t>|�f>?h?d�?'5K?K��>��!>䪇�^��>���=f�p���p�����ڽ��ѽ�HL>㖟�ǵ=��v�����->��_>Z5�=Y1�=�t��u?Ա?J�n>+=?̗ؾ_��e�b�y�]����>��s>��*?�7??�,?��H?�5?���=�<>�7��t��O~�>B�a>l/�v���{s��Ȅ=vj4>��(?�/3?NḼ9����h��^K>k�?�>R?��!?���>�$�k岾�@�j�ѿr3��eN��k�����2�<����ג�tSm>ȣ������bP�=y��>���>^��>}2�>� ��MW>8{�>B�>MV(>8P>f��=���=�(��|�=�pH�
/=���H6���H<Ig9���6���;�.		=�*�q��B?�^^>��ɽ��
=�ھA
(��>��x��>;�>�0�>Y�>V|>R��DT���@��'�|t>�VM?�?���9�J>�\�=�D�<��?w��>F�@>�za��~y�z�\@��T��>�$?&��=�0��9�˰<�,/��L��>�Y�=Xj�l3�?��8? ��78O�-~�&�K�����̃>n	m��4��oَ���#�#3�H�����@ڼRn��>p�?p4��8R>&:��띿�a��1����=�ġ= �?�A&<�i��s4��]�	�D?*�U�y��V����>����>��P?H��>=o`?=s�>��>��=YS9?j�o=^�/?�}�>t>?#V�>c� ?��?�?Sb1>�~K>�н̈́���"����L=��Y=�ed>]>6L<\暽��i���=��Iͼ�?>�=-���:��=+�>Q>�=�sl>�r ?>�@?������>��ǽ_�C���j������Hm>�<�>%��k��8+=�%?�{n?�a?��U>��G�
r���r��=.��>�ʮ>ܓ�>X%�=�����{G��2�=��r=.�s��v˾:W��s��Jl�K��=M�=|�=��f>_b~?��A?f"?���4I.���u���*��*��Ŋ[��A�>$�>���=�v۾J�6�V�r��{`��0���6�X�I��5=��=fX>��B>zt�=��>�w=�Z��%f۽/�*<�������>��>ؚ?	\>ԣ�=�Z��)���I?#:��Y��Jt��VξnJ���>��8>����?v4��~�����{�<��f�>f��?�*�?�~c? WA�M���@]>B�T>�>b%5<�<��2���ny0>'��=8z��镾�[�;�-\>�Fy>�tŽ��ʾ�$��*U���ſ��>�G �����㙾?�K4�����CҾ른���־�ߜ�w�o��{��h����=L� >n2d�lꤾ��?7��?I~]�m��$�B��v ����n��<��%��#��KJ����޽[��������澅L�-\�ޗ��p�>� ��M�����YP���2>'�>q�?��g�3�Ǿ����AG>��A>�½�!
������	��j(�&?vR?P�i`������IЖ=b�>|)�>�O�>�^��!㻾(W�>i�?kx�>d�=����<��7s���?c��?OQO?pH	�f�F���h�Ͼ��>�W�>�� ?�,��꾹�8?!��>̼����0�����l��;o,?�=�?�t`�=�q>I�>��>tLT�/d�4������D׍� �>��!=�ǌ��%}�h`e���=V�>[��>�4�Iש��w�>D��w�G�F�I����S���<�?�����=�@V>p�(>��!�J@���"���5�,G?��?��R?=37?�;��"پin�����=# �>�I�>���=?���>���>;��Z�o�-� �h�?��?���?��U?Іk���ݿ�Ý�W���e��{ے=fV=�-�<\�W���,>�ȗ=��b�;���Z=Rه>h�\>&��>=z�>_>?��=S����1��cэ��Z6��N�s���~H��c� ��כھ����W�ľl�7�h��Z�.~��[3����;^᪽�$�>X=�>dȷ>Y�-?���>�C?P潔�i��0�U��B�,�KT辘���S��i����n�7H�k���\�����о��?.����>���>�V~=+.��2��>)ӽ<> h�>���>â�>�n�>���>�M->��>��=�KP>�1> p��t���
�6�����������X?ad��쟍�1t8��k�G���V)>��?2�
>�G��	����t� �!?U'���־�Y��A$��Z�>�?�d'=N�g=S�dR���I�= ��<:<�>�@$>�����ξ��g�9�l=���>������d>�vN>��?d�E?o+.?{?> =�>�>W��=1�p>��~=G��<F�>QU�>�#?�=8?rU?��=Ǭp�mr>w�	>m,����D��hE��C������9�=^4ν�"���Ͻ�/D=?c�=ʎ�>ں�=!�N��:�;�?�x(?8��=6!]?<���4�t��䅿5����>���>)!�>��_>�T�>�q?ԋX?��>�Y߽$�$�7�P�wO�>�s+>	KR��|,�/R
� �<�8�=Z*?1$?X���<�ؽƵ=��>Ԭ>\L$?y?���>�%4��$��,��ſ/X��k@��P������W����E#��tf�>��~>(6���Q�=�[/>�w�>���>m��>N*<�礼�*�>Z=>���=!�>�'�=�m�=���<Q͞>5� �lf�y1鼾�w;2�;�Yl��Lֽ5�<m�R��$	���<�j?$;�>�ħ;���=��p��&�{����5�>���>�j>��>�=��H��q?���:�PŨ��B�>4f?��?<j���`>���=��O�8%?9�>aք=�bm���D����hX��y ]>�)?f��=nD���+�Z�g������ٞ>I�>��5��ݘ?�C?X��νM��!na��k&�)l>�����g�-�����6$�Mķ�+j
��x�*���2�?��?���/�>�F�����6Ͼ�}X>G=�> �/?���=KC���
��J���w���\I��H��=��ξO�?ԛx?X>Y��?Do�>�
?��R>~!?B�<�?Bd�>��(?O�>�9�>�*-?�"6?��?�S7>T�p��N���V2=��a;�����=a�>& �=Q㼍3�=&���޼g*=��A>�q�:)O�=,��=�=!p��(?Iu.?;c@�`��>�ɻ✗� *��?�}%�>��>,m*��[��@b=�0?y\?���>Ff1>jLQ��8G�ݐ۾7?	>�O�>��=>���>��.>-+>Bݯ�p��J�>���=ʥ��}��q��j�����J>�7>(�=ӧl>�|?�f??�"?>��~.��u���*�� p�:|�e��>XS�>�)�=ھ�4��8r���]��1��-�u�I��U=���=�D>�^E>�P�=3�>3�<�⬽%�ӽV3<���h��>�R�>�-?W>�P�=b���7A�0�??<:a�L���h�r챾���;�].>��>�'����>��T�O��{����%�j�>���?݅�?iFM?�vR�|�K�9�a>Cj>���=ؒI<S%s�i���kk�;��c>i��=�K���s��(=J�=>~o�>
j�����ߗо��������C��$��ےܾ�/��)�Ѿ1p��*a.=y��4�߽�>��G��{��D���ʽ-��Lh�wR���ҩ�\��?Z�?4�W�&����-�w@��v辷>�~;z��w־�u��T�ӾM����f��?%�Zib�D�e�x�?�>�1��=p���	����L�?�R>�Z�>dW?��Y�`}��3-�j�
>��V>��#�rn�l���2���u���>?;P?��]���s"�<��¼�%?)��>�	�>�Ě<�<澻��>jIP?WW&?Q�z��c��I���$��\�?Ym�?%�Y?mM	�ݮ;�H^�3����?��-?4H?|��'�ιW�V?h��>�:����L��N���1@��E?F��?�zE����>��>��>
��I@���$�z���2����>&Ӄ='�V��֥�L�|���=V��>���>�|���׾� ?x���%C��OJ��塾�a��V~=@n.?A�o1���\N>�t#>D&�S����t�w�;��NR?-��?�L?��?��	�/�|��
�����-�ף�>^�X>���=�>�>�:?��������������>a`�?�y�?Ya?'1���eտ����Q��jf�xמ�O\C�k�>z&Ƚ��Y�H��>�,�=  ��>�s�>UN�>B�>#a.>$1�=]*0=�q���}"�v{����w���F������վ�eI���R¼/��ke;���IC��%����������v�}F��EQ<��>6��>�ٰ>&?e��>:>�������$;-��*��Q�Jp�����9%���},�5>jt����И���=#?��!=�ɀ�j�p>�o�=���<���>���>�UG>B�=���=t�O>���>`��>�L�>���>�@ɽ�|>P�=0{�����~�:��Q��Zf���B?�Y������3���ݾ�����g�>�	?$�Q>��'������Dx����>�Q��f�Z�̽,��'��>� �>�;�=�Ȼ��%��x�S콳϶=���>�>ì��>������6�=�v>����>�>|��<�s%?)�Y?%}M?� =>�>��>���>H(!>,�>5�[>}��>�N!?r�@?G4+?���>=�}��Dx���D/��5�u�8�w	���2>`
�=�㾽g���NH>��B<"��~$�=Ds
>��%��n�G#�={��>\��>�l�>:3?.�������r�{��.?=�><�'?��+?��?|�K?��<?R���{���" �c�1�t*Q>!��=����$�ׯ�<�>��x>�a?}�?vV�<�E���3>�>\��>{#??2��>�܅=U�3����Ӻ����~־>���qu!��+�>� ���╾��?���=j������>�Y�>=��>�"?ec�=���=R�����>�<�>$���YV���U=GȨ=%N��=���;�����y�;��>Z�=>�S<Mż��ڽD��<��i�gh~���?��>OD�<��������ؾ����z��>��>�e�>�v�>G\㼞Eh�Q���G�wi���?�?ȏ
?Z�d�(g�>����\�=��>�<?�~9>𯘾�ؾa����Ծ$�>q),?O>Øͽ��D���w��C ����>Xr>�!нP��?g
4?�d
������ ���_���۾�Ī=T[���$����~�8�:�F��@�J4��2U���h����>���?�����^�>%%Ӿ�;��%��~����>�L�>��?z?�=��Ž��#�]ӑ�h-#��7h�\RG��ϵ>�F���R ?h�8?%��>��?��>�;?�|�<�<�>���y�>���>ݎ?���>�?���>QA�> �=��=�����z���D==���=[×=q =�#>��i=��F=e|:�����M^������ļh�L��}5=8���
��<�q�=+�?d�?�s�8�l>8�z��SL�"O&�qz½0�>�~�=��?�U,m��v2>+9�>�2?)D�>�8��꾦�������>lA�>!�>���>Zv>�oL>��2鿾`��='����;�����3��#�ԯ�=�U>�>�@�>-g`?~.?�h.?Ο%�+81�sz��%��z�=��Ż_�>n�y>
�W<�派	�!�T�z�}Z��I%��ػ�\6��R)<��=�f>�T>˫���>���=��0��7����=�r�<=�>K�	?�5?U>s>o�{�.���I?=������㳾XK	���1��)>��>����>X�=>�bS��ê�#JP�>��?�?���?�`)��g�ehN>��p>��;>�������#�8������>�Z>�fd��p���&�vԋ>bPT:<x�ֆ��W���㹽�����Z/��쁾ܖ ��¾���?���gb=�JC���(ɾI�2���<�`�@ƃ=�{ֽ#�Y�ƈݾ־uX�?,d�?uϾ4eO�HbF����C���|�<~8�N����վ��z��JǾ�j��/���}�D���,���ZC�>�R���j�� Ō�L�!���<>���1?�A�	�����;>��>�ȇ=�������n<b���&?9�U?c!�����(y/9"��>�(8?�B
?ܝ~>*¿�=o��>�3;?�d?� ~=�肿{����c���?[�?%;?:�.�Q�<�Rw��B�>0�;?�%?�y�>��z,�Nl��qa�>�4:?��>b��P�����&�T�?�:�?�X1�A9>���>��=�����5��(ν���eG����=��e��{��JW���<��e����?:X�>��3��x�n��>�n�.�`��^��4���*WC>ū�> �׾}Ö=��b>�F,>=Y��v���L��:��6DB?ʲ�?��+?��?$����g��Q��z
;���3�QbE>B #>��<�a?"?%��bT����R�>#��?ț�?��j?������Կ����#���7���>�'�='�n>T�ս�^�=���=�+X<ˮ���>�h�>�%�>���>�O>�]
>XS�=������$��飿{��k�7����4�&Ax���q\R�r�*��i���?����D���Q���c�L%-��o��6��sV�>7� ?��e>i)�>��>F��>�݁�E;�Qd	���	�>�9�Ļ��V[�@�I�R
b������;���~5����m�&?-�D�:>[�>�v���=��>�q�=�pb=�(z>Nz>����N�>���>��
>��=%:�=݄�>��4�����4^�R�C�����A(�a/?(���GT����$ܘ������F�>��?g^P=����x��>�����>��ɼ6}�o6��ͳ]�Xi�>���>p�[=�쳼"�;�������BH�=F)*>�+>,n<8�����޽؏!=��?|��G�=?��>�0? ?C?p��>Q=�6?�'�>��"=꣈<��;K�WK�>l�D?�?:J?��)?{�X=vҽV�<t��>hѽ����ò=��5��93�ny�<q��;7"��_H	>��>��=o��=��.=�?m>�;�~??�~�>��>��?;�þ0�{���U���û��r>�^	>ՀF?��?��>j�@?#�>d%�sDd�˕��k���$Y>�N>Ҷ:���:����x�T>�o�=Y��>֗�>|��8F��Yk<�>�F�=�C�>0�?k��>Sl_�Lp{�Q���	ԿG�\� �腞��L������2,��K&�x :�������ު=�%�>�e�>9��>r*>j�=�X�=jN�>�[>O�=B7�=a��H�<O���Jl=�-0<m�I=�J����x�}��;C�'���1�#�'�3����	�l�?F�>>F߽)�>կB�J��z�v��D>�Џ>LU�>��s>��U��H,�����f9�%�#���>v�\?��>�㑾��>$[;�=��"?���>X��=�/ɽ��s���&�x�X��>O��>�[�>�i=2w`��}�..��a�>$`>� ���?��K?�Vվ��ֽ��	���g�r��m�>v����x�̩��C*�]��̼��T�?�����E>���>(>�?-�z$�>j�����$�l�%"'�$>>�fi>�?8e>� _<�1T�W����3׾G��ǡ�x/�>j:#��~?�N?��->Cj?���>2��>�?�="��>�Ľ���>:e�>��>��>(v?[?sy?lv+�9����M���=I�ܼ���=��l=+�1>�O����=�|�=��a=�-Ͻ���<��>MrҼN}�<v��;S>��=J�?���>w���tV>��g��T�����C;Y7Y>�^O=Iә��)�;���=�; ?cG?���>W��=�)˾f��}���]><��>��?�;�>ԅz=���=�tȾ��s�#=[��=s5'��L�;���Uv¾h�ӽAOF>�|�>��=21]>a!�?e�3?��?K������_���>�]%��慽�֋>�?>4�=h;��"91�O�z��od��*�Z]���Q��*6=��>��=�(>�F�=e��=#ו=ͥ&�E��r�i=<4=�ә>>ء>?�?��>�C�=~�ξ6����J?�M��hb	���v�z�����1�j�&>�Q�>)���?�L<��g�`�����>�c�!>x��?��?�~?�<�8z&�A��>�.�>Uπ>��=��/��8��ʊ��Y>�H�=�TB������ϳ�
��>�#�=ş�#���=��v�ӎ��͛>��c�s��Kn������07�t�������84=22��3������<h�����=�:���-|��c�Fy����?5�?����E4b��恿�J�Jy��4>�F[�|�M��ͮ����ɱ��<"�_����";���)�g<�����>���+Y��	d���ao�A�>ŋL>?�"?y,C�
Ơ��2���>()?Ca�<M(�/����ֽ�o!��|Q7?�D?Ԣ(����i[��q>`�@?�|O?�w>GX��ݦ��%f�=}�?��Y?���;���3�{��z��|=�?�6�?p%5?Ó��A�<7��?kJ�U?y?�[�>ȷ־�T���H�U$�>¢N?�>T3�<���-x5�<�>���?�:��Xm=>�>�Z���bm��D��B,�hI��w=�:i�<G�=�̽gv�����=��<t_�>&��>&`۽�W徴��>�p���t^�6C��D���� =�/?�ža>~�=��O�-��s���Xt�+ W��??�?QIJ?^vM?��Ҿ�
�y��𡘻���>��=]T>I��
�>b
�>�H�
�m�0̾����>�h�?�m�?%�{?Q�L���տ~⢿�������;�^>��>i�~>s �2|�=�ȴ=ʄ>=]r�<�OH>�
�>?6o>j�>��->}��=�,�=B���"��{���P����4������ �GF~�W���*�X�d�ܾ ���~����������߽;� ���.���%��bR��A>.wF?v�o>�2t>
c>�˅=x��=����~Ľ�%�ɝ1�@'<�2�$������);�/7�w�羃��<GS#��?�>y�%>�(T>V��>�/=��<�3>ѕT��@�=1��>��>F^>�� >��<>���<�e~>t��=�t�>���=�B��Vuy��;��2���뽃 ;?G�s����� ��Ƥ�Mtz��@�>%�?@G>Ō7�����^p���=�>M�:�2>���&��Q���+�>j��>���=]���G���ſ�����)Z!>�} >�"y>�RK=���ðF�]d𼜔�>\�Ծ�>R���-�3?�OT?��F?~�6>}J�>
0�>��>x
L>��~>w�>�/�>vZ ?��%?=�>e�?G�=�N��j��?�ϽO�<qh�Y�=���W��=����B5o=:�I=��<}!�=�V=�B=s2_=��Q�'?�,?��">���>�8o�Gh�c]Y�NO;<��>`���z�?�G?��
?��? �p>2EB<�������˓���>ҫK>��J��nd��^�>��O=��:?G�&?Qh=Nnu�gm�=� �>Q~�>�(?��7?���>zE��b.��Dd�>�ٿτ�K;�n�\>�k#>�;>N���AQ�<�>���w+��� >Γ_>3�?R�f>���=cs�=�ۂ�-��>	H)>��0=q Z>(��)h�<R�=�$c=����=uT�̇��ۀ�=� W�ߙ����'�ڽ���sP�;M?�c?�ֻ��M>޴���Pf���¾h�m>g���>�=���=�#�����]��y@��C��a�>c0{?���>O����T>���<?�#>�̭>��>p��>���W�����E�=@��> {,?Ϯ?
d���ܒ�[�����v��>��7>~����Z?�Ub?��վw�	��'�L9��-1��ߢ�BjB�J؋��C޾�A�}�9�2i=�
��m���"*`>u?wX�?o����t<=C�׾#��NV��8���y��>��S=�o4?���>�='�D.�Y�%���ٽ��k��="��>ևƽy��>M�a?a��>��z?J�?�S?9�_�.'?W>���>�Z??+?�21?�Q>9"=!s�=	l� V}>6㽝=���!��0۔��uU>Pv�=�]�=̏�<�ݐ��U
>�������o�����G=ԢE=_vk=���=�[�=6�M>��?[�D?t"�M�i>* m�
V��hv��<e׸>=�%p=�}�>o
?*��>dVM? �>r����F:�t;�k,��B>�Z?�`N?���>��>�+�>h߾�e�/}=;Xj>o�R��ɦ�������Sk��d��>��>:ĉ>��g>��~?ےA?Gw!?�H����-�WQv��0)��<M�I�6���>�X�>���=e ؾ�5���q�g`��92���Y�:�J�i!=��=D�>&�B>DE�=��>�g=�ힽ\�?��:�ʘ����>�*�>P?�?Z>���=����B��*Z?����	�Ԃ�����͹�ܤ��d>k	۾���=o���C}�����5�f����=S��?E��?xŌ?����BX)��l�>h��>�_�=�3>�D���s��ȠZ���<Ն=�q���e��#2��z�<6��=j<�Ro�x���;�轲���z�_���q�K���*"ؾ�����1��$����u��>�����*��_��ʟ���o�=�`k�DEʾ��Ǿ��U��-�?a��?|��=��=<�_��9�v<���;����F�N��>���O�Ժξ)����������/��`ľ⤝>�TV����a�z��j(����i�=>7�/?�ľȹ��^B�;(x=�f%>�t�<"#���^���D
�P�X?��9?C�G����齧�>ΰ?�F�>.>����""ܽvY�>�47?3/?�᷼VV���2���R����?���?GO?N� �L�����0���o>�F�>n��>�`ǽ��־ģJ>��1?�/?��	?��)�>��(
8��پ>0J}?�,7�1�t>��>Qm>���Ii��h.h������Ћ=�V>9~�<7m�B�۽u�=
~>�ا>�x
>T0��ü����>������}農w�P+�����>6��3>�l�=bӽ�'/��
��^~[�d弼�D?X&�?�V'?o]J?E���������.{>u.�>�)x>D�f=�U��Im>/_�>�+Ǿ��ɏ��G�>��?f��?�-q?��W��˿)מ����������>�n!>Ʉ�>��+�[ >�π=�{/=ⷰ=?W#>j�>�&�>39\>��>>%��=�v>�|��="�t��j���o�K������������&�?�6����?!;bC羄+������ꔽ�B�!��ey��ى���1>�Y1?3ޒ>�!>�[�>]}>�����`$�e����$�����վ�� ��s����3���?�F�m�9[�CT��&��2�>�'>7��=��>=��<}�e>�D>�[�>h�	?�}>yj>p�=���=��P>��>�VF>�D�>��r=�&������9�;���X�|$$;�&A?��d�U��Tm4�w"澜���}�>t�?��k>$�������t�E�>��F�h�T�©��C�}��>�>�_�=?�@��3������꽘"�=e��>�5>5�|����I���3�=�r�>��Ѿ,J�=��n>� *?R�w?�1?��i=8*�>^PJ>�`�>�y�=��>>p�=>x��>w�?�n=?�4?l��>��=o�U��	�<c�=9�@���w�Y;�������$	�Qz;��5�7b=B�H=����o>=a�.=��¼�(<��<�$�>��8?JA�>��>��9�>h>���M�ݑ�@>������>��> �?���>�#�>G70>A�q��cþ<����>��C>Ä^��v��p���w>�ji>��M?��0?�b�� e�i��<��=ꋰ>*P?YH)?�M�>�_>�̺���p�ӿa+�FT����W�<w��=�q[���i� >N���"۽�D�=�$�>��>q�)>�i�=�Љ=->gU?��>�n�,a1>-�b�֌+>Ά��Έ�=9����V>q'��N�=�i��=���6�$��U�=m�<J&�<P�Ӽ��.?D��>��2��	��4������M|��J�>�{c>��>��?�t$>Oq��SZe��8�����1S�>*�s?��>`+~�.<S�S����;�m��=	�0uN>�>:bp>��Z<�t�>�7�>��A?h�>��k�$�e��Ƌ��B9�n�>j�,=WF*�J=�?B�_?1��p����6I�����n=��ؽ����I����"�<E*��*	�� �uG�3��=�%?"��?�+i�N�	>�1�����a؃�ܧ��˘=�Ӂ<���>�g=;#��������n�w[���X*>&��>�z���O?��L?y?.?��?;�/?#⼘;?%M>w?k3?\�,?0Q4?��>�-�<���<���7��>m�
����
�>=yѾbY�=uM >t|?>`�=<	ڼY>>��h�?�=Z쇽�[��𪓼��[=y�>׿;>��>6�>J@?pI'���g>�z�<>�G���i�!>��{>ĒP��n���W=�h�>�$?��.?A>b��[���2���p`X>V?+�N??<?W�>�ƴ>��Ծ�&X�p�=��r>��i�MⒾ&&�q�¾����i>Z�M>�=�h�>Y�~?D/�>�?��޽�-��������
.>��=��>B�>���>�?�ِ�r�q���v�x�G���Q�%���'>0��=�:�>�
q>>8'�����$�,�m��>{E�Ǆ���h`>�4�>�y$?JQe>9�=�~��S��'�R?䤾c��Q�(��ý�hʨ���$��w�7�ھ���m����r�oʧ�{j	�F?��?#_�?*�V?j�0�MƽM��>*q>v��:&,>��H��@�μ�2�=�k�#@���3N�i%�<0Fp>|9L>������Ⱦ�'ﾃ�������]�r#g�������ܾM�k���_�����.��-ύ=� ɾ8-����8�h�>��\<�<!��u��ƹ��D��PW�?t5�?��y=?+>8XJ������޾a����E��߂�ޕ��I����� ����/n�Z$�Q��#�߾���>��Y��*��(�|���(��Ƒ��?>�@/?�8ƾ�������F,h=�o%>���<�<�㪋�Ҫ��c�+UW?��9?yf��	�����h�>��?)�>1h%>O!��wM�w0�>%M4?��-?\�켲���.�� ����h�?���?!�M?�e�ޞL� ��G�:�{>��>�~?*ȼ�ń�W��=?�S?7/�>��$�;��� �A�)�>d<^?��K���>ΰ�>$v�>�=7庽.��.�5,[���>v&<� 1���t�<�@�<�F�>�W�>�V.>�����e�=x�> }��I�:�'5��5�
q��T8=>�?����bxZ>���=�诽 v'�TQu�?������giH?ף?�J?�7?.��I����'B��t!>�ƭ>�O�>j{=ļ��y>\n�>y���T�FQ��m?}��?�I�?bu?c�\��2Ͽ����y���߾�(>������>��;�]>W� =:��Ct�=F�>�(�>>_h>�R�=�L�=2-�<��&>�_}���!�#l������<?�4�4�=)�B�R��z��k,���O3��t��D������=+=� ��)K�g����y=p+����>�p?�?�T�>��h>���>���#� Ͼ�0
����ۤ�T8��Z��2\����+��r���%��g�>;!�}�?[�="��>�(?\b彖�
>Rei>+->~9m>�>��\>��>;�u>�\>^�l>K[>��">=҃>٘x=����ꣂ�ye;��\�U><KC?ƁX����k�.�����7��H�>3W?�p>!������lv�b;�>�<5��o`�by�ϕ��݇>��>lW�=	���0<V��o�h]۽l$�=o�>7b>e��G���i�pcu=��><举Y�=���>��4?C�?�0?N�ܻ�ш>�|>.�>Su�=u��="�=�z>��?'??IR??���>��=#AW�.�<Ғ�:��4��Wн�B���<y���1�<�ţ�>�O="�4=�xG��� =���=�����=<%�=Q`?�\#?$ �>�*�>FX�;��;K�{�h`��2�˼�e���S�>�V�>�h�>�4?i7?D�>���=0�ʾu'�ik�>�H�>����Pj�N�<�%
>InT=�o�>*%?1}��q�m��j��£�=0/?�?�K?��>wW��ȑ�mA����ҿ_�&�7�'�C��;[l����=t��:K�r>g��;Zv���}>�8�>V=?�>68���5+�c�N>o��>�b�>Of>�߃=�}>x<��>LD<�ޅ�W%����;Q��=ԓ�f�=��=f�e��f������R1=��M�տ(?�_#?(d���C����!�K��>�_� �?�g?�<?�c?"�>x����\{��Og�?-��C'�>��p?�=?�{ɽ�2<=��B�z(\���l#;t�=b�>���>R�?>!&|=g�>%&]?�_�>�B�H\b�9�t����h�?���=��f�~)�?�C[?��Ir�3"�Ȑ0�
��@J�=��$�pKQ�0���d��NoA�A�������<l�=Pw?2��?_�m��b>�վ:j��������\����=�@W=X/�>b�=Ɖ���{�u��O^��3ى��@j=�$�>Cs�=�t�>ľ?]}?s�c?!�?c�?��-�#B?W��=��>���>��?�v?��?QO�>8D�>R��<H�k�Y+�����T4;#S뼥	�=6d>�>*>�M`<��)=r#=C�<3�P����QC1<�m�͟=z�=��=c�>4?,(?RH���V���W>vu>$���줾�Z/����i���=Ϲ�����a�>3�.?�%?�r�>��ž�L*��~
���>R<?0X?Y�?�>�D�>����Ӿm�>�c�=�>T#���8J�V%�'���=e=�>���֚k>u�}?��0?/(?�UQ��c3�mj{�1���m4���=Hp�>	�>�b=��Ͼ	IB�P�x�`2e��}5��lw<e��q)=�
>z�I>PE.>+�p=��>��_=B6�M�i<���Pم>�n�>s�>S�l>L�>�v�����;{L?oǈ��w�J��Ś
��^W��,R>q?�>n11�"��>L��v됿з��W���٬>��?)�?b�[?�!E���Z�A>+C�=���ݺ(>Z�9���Ye����������%�Y6ٽm9@��N>#��>�Z�<6��U�yu�E���,sA��� ����������~�\��9��Bpf�
��<�
�������\.>�ɼQ��N��p����?ZܽC��?���?\	����<��a�-���Ӿ��>@ݤ���D=�0TžF$پQIҾ	l��ھ��m�$����\w�>�X�y(��
i|��!)�t��>i>>@#/?�;ƾ�������'�e=�9%>|Q�<%�ﾸ�������|��hPW?�:?qe�Ƣ���Vݽ*�>d?���>�|&>8ȓ�B�W�>�3?E�,?N��7�����+��eN�?@��?\A?i$(��=��	����f@ ?� ?���>��N��ʫ�*���F�?|IA?�$�>��2���"�T�>$�i?�N���h>�?�>Xȍ>�Lؽ�R�����9���y���c>�r&����>�]���"�* �=:O�>)O>s�~�2O�����>�m� �g�Pn�MC���ľ'X0���
?t��|��=51>¡ԽW�8��G��!0��W�5��,3?"�?�#;?D"@?ӡ!�@Ͼ���k�=ƍ�>�u�>�t�����G>Qk�>���r���Ҿ=�?�&�?&}�?�k?+�Y��Fӿ
��g�����4��=�(�=i�>>��޽Э=ӞK=)���J=���>A��>Wo>/9x>`�T>g�<>��.>꤄�C�#�[ʤ�(ْ��[B����g���wg�|	�Q
y�`��mǴ��ｾҙ��ɣ���͓��G�g��K>�ZS��`�->�0,?Ԡ�>H��>08�>�%>�ߥ�.��Jd��J�s�C����nR�V����3K�aܱ�2�Ӿ �ɾ:�<��� ���>�u$>T)>�]?gĝ�+�=�p>��`=��>*Ȣ>��>O�~>q܉>��=�偼L*�>܆>3�>@�w=bτ�. v���<��[�G��*�??�i�Wh��j�2�9T�S���}K�>P?��A>��$������6q��?�>W���T�N�ٽ'G��{>�^�>3o�=�ն;9Ah���g�����u
=��V>���=�û�=~�
����m&=��>c���#>bo6>+?��?�:?�x =t��>�bq>,�>Z�,>�fd>DG:>D��>f
?��.?#�-?:{�>���=ɧ���<����2I<����L�5�?3$�	V���f�<?������=���=W�;zr�=Q�A=��꼝��<� 4=��?�k�>��>˸?��=�~侐v��-k)�	�6���8�]��>��=.?{��?CO?<
�>�J)���޾}���=��>�Q>wQU�);`�5�0����=e�^=m�2?%?����=�5t=g澽(�>�>�4?u�>�!��4���P�ٟпp��\�,��{��б��-��N���i��h���^�����<I:>�ja>�_�>�Z%>{_�=]o�=v�>��>u�->��<,,0>����+����}��=�����=ޥ����H�t�0=K��^�O��Z��ʗ��qb���l�f48?��>ꢁ�-��p��
x!�)�h��i?qh'?S{	?��*?�ƣ>����	@����[�ɾݬ�>�;?�?��6��Ƥ>:罼J&�=���>��> Yb��w���):c]�	L�&O)?ޗ"?q�>���F}���ĘN�n�>�;�=sOg�}�?b�\?]���쮽��!�ߙI������X����
rt��������� �xLɾ�0�^���6�=��>|�?; �N�>3	������K�����9���6��=��
?[L�=�RT<����;���+����(�7�<�>���Ł?nf?)�>ٸ??�g�>iBB?�A��O�)?�	?��>~y?�+O?*��>(�H>�j�=��|�.`��+�>"rH���꾪�]���
�;��8>��3>f!_<m��;��<��d=cQ|=+a�<b<`��=I�=��+>�5>S��=��?J��>���ʽ3p�=k�`<��w�7ض��9������-��}j߽�`¼y�>��5?A�?4�W>ܠ��};��	��I>�r
?2�"?���>��=>N��>ŝ�����]Hɽ�y>H�k=L~���$���6����>���>��ia0>a2�?)?�a:?1��=��#���c�l�̾<JT>/�>�M�>��>�nG>��Ҿ3�;��������-P���<w�(�q>v��>�4�>1��>޸�=�\6>�el�?�`��=1L��l_B��%�>��>P�>ci�>!�C>&(��.��)Y?�۾��+���辊TѾ~q���n�>T˂=Q��c<�FO���M��Ԣ�o�*��#�>TO�?Eh�?�^�?W=�/�.��i>1�>>�jV�W�ؽ�s�Z��=l�>���>ߎ>\Tk�ͭ3���=�>�'H��罁$���ľ��y=1���j+T��o��,߰�"n���'��V������=�;���]�<����􌁾�y�v���p�׽����բ����jܙ���?��?$��f�@>�>X��L�uWо)�L>�뫾�F½T}�<�ľR~	��JϾ̰�� ��7��g�?͡�&��>8�V�/o��G�y��+��sϼn�8>�0?i�ƾq�b�*�Z=�!>���<���8��`"������(W?f�:?,6뾗����?ܽ�C>��?uu�>�#>d/�������>q2?U*?=_��|�������}b����?�	�?e�E?l��J?����� �(��>)J�>o��>Y��¸˾����8*?�d+?��w>"��Z���?k7�ni�>v�d?'_�����>V��>m�>a_'�FȄ�\����a����ٽ�6>y��s15�o��Me4�t<>��z>j݃=8�K��YǾ���>>ک�l�>��"�G��������x?��¾W�=���>Z���/D�����Gڎ�Զ�2�W?�f�?3>E?��C?/��N0�\dӾ��%ԣ>,��>@���lՅ�imT>���>jR�ڂI��/ݾ�	?}��?���?"�I?�L�u�ǿ������񯪾�@>k�->�X�>߱�<]��=��1=����O�=\(>:��>P'>��>�ρ=��=D�>�z�\_�u��򇿦,������zR[�&}پW��p�&��V��mX��ޘ�B����H��޵O�#d�X�̽jk<���i>_Q?k��>���>��>�є>��~�"/)���uq+��1�M��j�߾$��ޜ�Ǽ����[�楷�yj	<�o/�]�?��=��>y? +1����<�>R$����>6�>�:b=�
>BnV>�J=Y��=���><��<�)�>�Њ<FY���؉��EZ�r�}����=��9?�I+�鎠�T.������ʾ��v>�6?�;�>_��D���a�c���>�J��?�VF½ثC;͜�>%��>�n�=�Ѳ��a��z�)�Ǽ�o(>�K�>T�W>/�=s��BU(����=`�>�Ⱦ�>�h>< (?�r?X&4?���=���>S�[>(Ɏ>���=��W>�I>�(�>'N?�7?T4?�V�>���=83|�% �<��<r�;�����m_ѽ�����H����<ВC�u"=��f=?�d<��C=�qC=+�������j
=e�	?�k�>Ok>�;?+@�>V]2����?1����V��0g�>#Պ<H:�>�_?��?�]�>&��<�;ݴY�K��>q*0>#�J���d��R�+T(�}��>EWb?'%O?��Q="k�����=�=B>e�I>+D>��?R_�>!�>�N>��п�(��)����9��	�ZUK>߂?<+�<%Lq>)��� ��;���=�h�=窨>e�>Ɠ�dC>
�۽���>P��=\ͫ<$��=���5���Rt��4c<����>�#==���&m�<�h��=Z2�;�o2�A�޽Ej���j,?��>Y�t��]�j�龔��y"*<f�?QK9?eB;?��4?ϡ�>��־�i���������&?��?~�?����>��W;�=���>Ԯ�>��(�-S�����z��)�=-$9?�D?@��>��5�̯y�:ƕ��u?�Yt>L�Q=�Խ}?ϻt?��ھc�r�mOD���!� "��D=�ш��p���ƾ��#��N�ԝ
��@�Iզ��:=�?מ?��Ҿ��>�q��������B��ԓ%>�)��L�+?����쌾{3������k���̼H��='�>��ܽ7�5?�˂?�E?�i`?��?���>i� ��8?��>�u>>��?�M:??��>՞�>��i<�:>>/>ڿ�5��Xf��y��<2N��?��=mtd>[*'>|0<c��=�;m��=*�L���e�{�J=a>
�7>_�>u>���=��?���>5U%�Qm}����=I�=�*^��ۗ���l���˾�J���=���=��?f�>?��?���=G��8þ}���^�>`�'?��B?�h"?ef�>���=H�߾�����I�c(p>�9=������0���f��D��>!2�=�՜�u>�;�?��/?x�?���Q�5��J��B����j>��t<��>57?���>-ѾCWM�����5c���J��m��UӾA�d>c�>��c>vI�>b5B>~Y`>%=ν�f��H^��a��3н//�>5��>_�>�gT>C$�=�z�Szܾ�!U?�ۙ�Z2�0%���E�镾B��>��>���=GC�>=��������9�|�>}��?�? [?N���X�2���a���==��νNѭ��!.��ֈ>��>p��>��>�o��r:���9>Z��=fYY>�d�=�|��9u�#�>~W����V��<�i�7���)!q���j��x	����,>��þS���<���M�%<�3^��$���~�����P/�?[́?�D�=��>�2-��"�ج��c&>n
Ⱦ6"
<Ja������ξ��ݾ�{����� �ZA��A���>�Y��@����|�M�(����5~?>U4/?aƾϴ�D����g=e%>��<r9ﾺ���گ�����cW?u�9?Q��*��t���>F�?Os�>��%>h(��L4��&�>94?p�-?8?켳��:������l�?6�?7@?soF�z�@��'�����?��?��>7���˾A{۽��?��8?�̻>3d��$����
��>��[?�O��Rh><��>m�>�� ��3�5����k�ռ�c)>�/������c���=�VP�=�m�>��i>[`h�
����>0=��N�X�H��������!�<��?���+>i>�I>�(�Q���Ή��"���L?��?��S?�i8?�\�����������=G��>�Ϭ>>��=	����>S��>�d��vr���՘?�I�?{��?p[Z?�m��n�߽��(���b25�j�>$g<m�>������<�Ͷ=-�(��>ma�>̱1>-��>r�P>գ�>��>�~���*�֕����DVc��6�.Q���a9�{���O"��x��ع�㧭���g1��s_��U�_����oR���p��>>F��>{�>���>k>�=��>��=�׾�D���	� ���������'��e�ھW-]�K���S�l���	��?;���1?�<�>?=��=[��>Q���NȆ>*�=r��>���>�.�>q�0>��>>�>>*�<[��>~c�=2Z��3����m���7=jd��%!�>��k��S�4&���!XǽV��>��@=5��=E<�Z�hz��_<?T\8�g'Ͼi�7=���;5�;��?T�>#Og>p�(�����aBm>{�����>���=T�_��j���,�=��<qj��G�>ܧ���!�?��?P[9?�!	�R ?�>�����=a�L�)im=J?�?�>]�s?��Z?�MH?|M<y����=����@S�<ۙ�G<F5�RO-�l�E>S]�=};=�c�=���=��&��"��䏾߄ʼv���_�>��-?�0�>�1�>��Q�Q�I� �D���~��4i���8�� T?1???<?���>�=�D�>���='��������>3��=z*Q��a�G�����>X<J>�EL?ݢb>���<^�i�.f�=\�`>�>v�Z?%�?7>N(��s��`���L.�ya����ϩ=�|D����=�[��?�%� �<z�p>�RF>���>��Q>Ͻ�>` z>��>��>t�>�����,�X>�����	=���=ԙ����<~<�=*�7	��h۽����ڎ=#�<&7�
?˻?����]U>
ܽ4L��Ӿ���>\�>r�>�!�>q�>>�k��Q`�,��W&�<7mQ>@�]?N��>�*����s>IM��W�F>��?g��>7�A>֬v��_L�H� �Iq��^��>8֮<z8>9<!�E���P�yW.��
8>7 =<wȽn��?+{R?#��C��z��C�Q�<Y��'�";�!=�@+]��I��z־WS2�o����gQ��:{<#H?礣?�˿��M�=^����Պ���������Ej�I�f>�?�U�>3�c{a�y[�����X+��?v���>'��<u>�>��?m��>1)h?K3&?��?��D�<��>ʄ�=1�>��>�P�>��>�S?K�H>h=�>��=�UV�� �(A��1,m��_���D>~qF>�8U>E`}��$�<��;;�2�cͻ�r4׽U�T�vv�����8��)��-p=��=9?u��>ެ�;uT�.1Y�2�<<6�=���>��/>#�	���AJ>�Y>�J(>�u�>h�?�>�����(���.>�L?�@?�:?U�W��1������=�E:�Ag@��żP�[��D�+�"�׼��<>���>;��>��)>_~?p�H?�UT??�)��:��!��� �R��?��Y��>t1�>��e<�Ӿ�t�h�_�-V�%M���)7�T�,��x�=�s>�ݻ��'��>�=��K>��{=�+=��#��rF>����i�>��>���>�u�<Ւ
>�ֿ����2H?��)�[���	ʾhἒ�>@�C>�=�=� ?WX���y�`椿vY>�0g�>�'�?�D�?��a?�%0�5|�W\>ne>��>���<I�C�?>������:>���=��������P�;��a>y!�>~˽����ؾ��i���wT�ܲ��#���¦�����kپ����+���1��=���������%lc��,p�������L��N��4��?J��?�vu��9J��ڂ�L�þo���¦=;0߾�[����������8���)�Li¾�l���M�L�:��0�}�>��u��0��3�w�"�1��s$�)%~>c�;?zP��,���k�2���e>�$�<[��5��������j�4H?c�/?��ݾ�^˾?2���>E0�>�S�>�D�=����sG<
�>�)4?��2?C�V�Ϡ���U���_�Wi�?)��?�[K?�\~���G�f���섾���>�?�?T<b�;����^t�~2�>��O?��>􇴾Zy�}(����>�F?_�X��$n>O3?n��>L��TFо�����ľ���V��>p�v=��K�����z$�&�����>��7>|���\�!��O�>L����*���9����QB��XE=�H�>�۾�47=�`�=�A�=��7��������<=���X?��?�3^?8!? e��oR�5]�i�c=lm�>c��>_!�=m���|��>���>z���O��j	 �F��>n�?�S�?y�j?�R�_~ӿRU���˾TǾU��=?P>ļb>�7-��0>�:>�C!�������/>��>�>}>aRU>�
�>)��>�΂�p-!�*=���8����I��!������������q�
m�ʜ��B�f�lğ<G~�o����B�b8���Q���[,�BZQ>W�>7��>̿�>��4>���>����!���Gހ�-����1�i��'X��L���e����P��͐�RLP���ʽ����)?L���f=a�>â�=l��=���>�ս��=R>W�>��>,�>��>��=��>l�==\�>�)w�[���냿�O��������jx?�T=W2�h(Ⱦ2Y�n]a�4?��?��:?�P`���������E�?�q����̾ W=�v ��w�<Ps,?�M>������<�gƾ�Jp���":@+>7��>�Kk�	 a���ž6ꇽd�>|�<���>^�8<�1w?2�?�?N��.?ω}>��Oʄ��Aþ}��>����|>�^`?3cB?�a+?���<��k�{�=-�o="e˽�	q�Ƈ`��$<���,<�ˢ=�°=���=�h�=V�>m����=�HX����H���>��K?���>Zk�>y���z$��X9���M������(>�;?�/?\a>?@@/>��>�3>�z<1�O7��9³>b\�>�U{��!a�^}��2�>xQ\>��8?��?I��' ���.��v���>Ӕ�>�!?T��>�>h�	�25���ֿI��y�&�[R�=w�R=����c�>�_R�m�G�i���=b�?�{ù���>f��>�S�>���>���>=v,>7��=
>9>�_=#@T�qz��M��=J]�Q����>��ی=��j��������y��ȫ�6�������?��-?ߨ$���1=�%������l���>�Ġ=<��>��
?#��>�lľAp7��&#��[����?p�S?�:�>!�v�w^�=t�>^�>�o ?�L�>�n��֎��n��4⢾.�=Sͣ>yh?���>�߽<�O�K}�ST�����>�<O>)����?�7f?'�+�[��d����o�P��Rf>��߽q޽�:��37�u��J���?��[���6[�	\�>�;�?�����>/4#�����Dy�����lI=���>��?N ?a��锂���B�������c�D>p�>���=���>�Z3?%\?�f?X3?���>���M �>��=;��>]��>�d�>��?g��>\ؖ='`�>S:�=>(�=��3�{a��`U=�QI�ɓ>�C>j�">��<|�=�@μW������4�}K?������;�� >2�>/�8>�?�2%?� R<��=����E��}>�>��f<����b����=��>��k>��4?.�>R��<���۟ؾ���l`�=�(??�f�>,ov=��q<�������#��_>X����rU��g`�[�`��5��
�=��>��
>H��>��\?� ?�O?8�0��d7��U�1��+�����<K��>"n�>,�<�/3�(��;�v�B�j�*n#��KU�����q�;>���=�r)>>��>���>z�> K�>̀?�"�x�ĭ�=�G'���o>��>���>��i>�0>�鳾�Qƾ�F?嘾>��������ľ�a��"^">?>F��G�?��&��,�킧���>�"�>��?�H�?7�f?�-���#�P>M�O>��	>n<�;D8��B��Cz��O>H9�=�su��_���̑��b>��s>�S��_ʾ�⾚LJ�*r��P{Q�:���n���Ҿ8��"־�{2�����'X��}Ǿo�ν|���>]��-I�}�&Q��5l��?�$�?c~�?<�m>7����Ǆ�����R�-��=b���;�=8F��z���S�}���u~��)��o���>#��t$����>����h&����v���U�2�6�x��>��!?>R���G�4�ͩ1�`m�>��K���L��
���"o��OC?v�?$���.~���=7%����=T��=_��Y	E��>%�>�6Y?��I?�;��w��],�[��6�?���?�-@?��G�$A� Z�z���?��?��>z���žRe��
?��6?X��>a���Ʉ�Ǫ��>�>�Y?o~N�
�d>m��>��>.{�����%9"�}�����ǻ��6>�O��1�~1s���?��!�=�>�D|>L�Y�򫭾2z�>�&Ҿ�M��P7����
�e>�=�h?��N6>�>Vi���2�A,��!���@�
�lG=?�Y�?��H?�|&?��پ�f������Y5>@��>��>�N->@�����>���>ՙؾ6�x����?��?=��?��^?CFc�J�ֿi[��8d̾.���W>�,�=�27>���Z>y->����$S<��.>_��>/a>ah�<�6�>���>���>C���. ��k���y����(��Y ��0�/������`�C)�%����z�Vc۽�_��i���P<�Ÿ@�BW�H�6��L4>:6�>���>���>P��>���>1&=Uľ�Jݽ%����������
��ʕ�q̼�G�L����Bv�ܵ�o�?.g6=vA���>�ҽ݀H=�˘>r"=��>���>3�B>"��>:��>.d>B�_>I*�=r�=a=�>	w�>8����!���G����=q�X}?l1��6��龃��ۢ�� ½��/>��D?NV=�r;���G��>�?��l�ꙿ��,>��$:�=�I�>�yD=�%��0<������*7�/o>KD�>.��=zX<�4��׽��6����>o���>�v>Y�,?�%W?�t6?I�=
+�>L&*>g�J>]�<<��߼`O(>i>�B�>�8?),?9��>�O�=:��"t>���=�[��幪�!Tͽ�Q�я=-�=�����;{|�<��8>U�>"���:��?Vm�<'/=�x#?�75?K��>��>��|�K�v� 2��v����(��>ZP&?!@?�H;?m�>�f�>�R�gIʾ��ǌ*����>�Z�=S�Z�����˧<����>�Ԏ>L?��	>�VK��3>pU�=��o=�e�>-�T?ʋM?�o�>���>�7��]z���@ڿe�5��Q�g��=%�ȼ��=��۾��=d�>3��<Uǆ���=�S>�]�>�*�>�$�>�?�/�>�3�>�=���<`>�x��H�=�}�=A��=^#����U<媐�+��<tq|;����\���>�m;2�<�	�=�G�>�t?��=Ю��ؙ��5����U�@�x>�M>4��=s`�>���=i�=�l���@�b<�+<&?_b?R�?m�L�4�<��*��>�2��>��>t7>b	�g��t�ڽ��=F��>��?�1�>�Z�QOI��H����|2K=�(6>��c�?c&�?~��'!	� ҾXL�Lz�{+�>U�Ӿ�������;�����9�%�E�����B����>C�?������?>�B���¿�Ӥ��3�|�<�8�>B�>�Y>�{1>澗��=����& 	���Һ�	q>l��83!>r�$?8��>KR?r�?^��>x���_?	0&�j4�C�i>U�D�-6? m?��:9>*��>�V?�F����q��d<��>�:>��%>�t>?N�<x�>���<��<eƼ�;��Gq=n�1��Օ���N�i��=�.+>�{/?C,?ٌ��6��J��v��Tl���O=�Q����#�W>��>� �=��>(�>��>+>�оk��u��e��=��?�_-?h�#?��=�Z@>�:\��Q=/Kֽ|�d��y��?�羧�ξֲ�H���)�>���>O?��>x~?�=f?+?�R���B�Cq�:����Ⱦ��V���>��>��>c������cU�F�e�|�%�V�������ͦ=������q=Q�X>�)>%G>=�����!�=9�	�u�.�:¿=�/�>�'>�{>�1�>L�=��������R�G?�H����MY��{�Ǿ�ּ�+6>�zR>���t�?���%���we���=B���>�s�?gv�?��`?{l@�3
���Y>zM>�>��=ӈ2��m*��?��R�4>��=tU�5�4\<�d> ��>�R�������F޾�G�^���+3>�හ��}�4
����Y�Z�F���=h��%=F�ݾ��s�V4$��cg��E��KZ=?�����k+��$�?� �?y�ν�}ھ�<�f��	�.�f�<>�/����
�����յ������H~;D;b���ôR���Z���@���>E�"��싿��I���*��ہ�Ҡ>�*?����|�24�b�Y���=�?½י�ϭ}�����Ig]�Ř:?�}?�<����!�����>�!?
Y	?�*�>\�����׽�c>�R?�r�>�1%�諊�s���>vB�?�$�?�??�(H�>A�߹�|���d?r`?Q1�>����˾�&�?�6?�$�>�c�5������>��X?��P��fa>���> і>�s�:-��%��������o�8>��)�q���oh��>7�}T�=���>�J�>@_[��Ы����>�����J��D��B�Q�:y�<@�>c~�r��=�V>x>$f+��U��(ˉ�VK���EP?�а?��V?S'4?|:��%�揕�uM�=G�>��>6Ҙ=F�%�<Ɠ>���>�xﾪ�r�����?\��?��?�]Z?)�f�UGӿ5��.�����V��=�$�=�>>2�޽Rɭ=��K=�����X=�Ӊ>F��>�o>�:x>��T>A�<>�.>h�����#��ʤ�(ْ��[B�� ���1wg��{	�{y�����ȴ���ԗ��r����ϓ��G�����U>�;<��4$�=%�? ��>��?��>"��>�8u��긾a|�ܯվ�� �w�$�?��^�|D��{��	=�!��P9_�;�	�>�x��.�=�s�>��>-�H>r^X>�t>�R0>i�̼�,�>tO�>��=�X[>��)>��`>$����>0?A>�;��1e��)�n��j���XY�5I;?[2�<���:� !�ݴؾ�T�O�>�1�>0ش>eL����c�׏Y��?3���l�̾6�%>�=k�h>>]��>��*>B�b:�r�各��g%�Q��=��>���3wE>�;�����ey��~�>�ʾ/HB>�AW>��*?G?�V?�=]��>$�c>N�o=������>��3>��>�)? e2?{�?ݢ�>i��=5n����=i�a�N�d�:�=��佽�q��@�=�P�=���}�>��>�4�G\�=	�=���iڭ��z3��� ?E�?���>��>�� ��:6�C�q��C��Ĝ����=S�4?�!?.�:?&!?f��>�!�=�Ӈ�?���l����>�$=dof�莇�c~9��U�>l.->]�g?%�?Ff���8g��d�>O�=�d�>d�9?�O?cQ�=��V>�n->�L�C��'���0�<�6=�⌼e��=�u�����=Ђ���ٽ��K���>��I>
z�=��^>-��>�U�>���>$�_>0'U=<҉=�����&;�4�����<��+�0��;�9º���");��5�e�N���ܼxH~�z�<��;`�?|�?�j�X{���P��o澩���y�>�!�>Q`�>�z�>o޸=<g�\KY���A�x"<�֎?U�g?�?@�?<�=��@��j<�r�>ʩ�>z'>Iߒ��@���_C=|��>��?Xr�>~"2�H�U�i�#���U�>�T�=D�K�wٛ?%Qx?������x �����9%��*�>�^J���J���<�@�-u&�AD�M�vh���$r�a?�>�Ɩ?�QW�\KD>��Ⱦ�륿P����Ф��t��>�7L?I�^>������+!����ũR� %��ن>6���7�><�?@��>9v?Z+?��?�Ǵ���?Y]';m@�>�3>���>ﲒ>�>?�d�>Z�>��I>�D�=VF(�*P��̻ϽlC�L�_>Ɠ=>�w�<գ½;�=	��=��<<�A+>�A�<�����6���=���=T�<�=�'?g �>`V��O=���������"�{��).>dn�=�,�����M}�>�\�=���>��/?K��>3�a�;��jG=���=,:?�15?D!?��L>l�2>�U��H��;y���[��ʽB���H�&�z�~_ �{F>|��>���>}_E>�bn?KL?��F?-^Z=���f�4b��	v��I��-�?���>�(�=I������7Q\�k}Q���:���p��g�=1�=[?>��O>��>ص=���=W�q==�m�js��u 	�x�>�G~> �>��> ,><�ھpD"�� V?�����'_�����Z)����:۰D>f��>'�C�GN�>xI�<)@e�袚�'T�߮=`9�?�ֽ?�4?�D��Q�Y�V-�2
�>��>��5���о��>O-��s����>�J'<�l���©=�u>��o>��+����}'��4���HIN��p����� Yо�⦾/߾�sT��v�=�"u<L��[����2�9���k�Ԇ���o����`=�'��4�?aX�?�x�=�j�Y"p��Jо�����Z<�?���+��2�ľ�" ��,x��Ä�q���Zо�(���&����ޛ>I-Y��-����|���(�����t0>>��.?U�ž7S�����~of=o�$>r�<��#������ۖ�C�V?Ӈ9?[%�6a��e�޽C7>�(?�k�>�a&>Z��Y��跑>84?��,?�������*��"���Z�?[��?��@?��S��~B�� �+@"��n?��?X��>�c��x�ɾ��⽝4?0v8?K�>�9��ƃ�����>�W?�~O��[>���>g�>���c��A�8�:
��Y�v�d<>��.�#��.	[�~i7��&�=��>��i>oe�ᘫ�~V�>w����N�:�G�H=��P�Pm�<g�?���>;�h>�>�)����o��������L?a�?�1S?R�7?�P��9�cb���Q�=��>�\�>#��=/�
�[�>f9�>S�羉~r�'��o?�$�?��?��Z?BBm��K�@c��D�þ�I��l�><�=��A>����I>�e�=�s�������4>��>�j>�)Y>��_>���>$��>�j��F3$�S|��5T����7��T �I���w?��y־-_��K$�J�� ��@WʽW������e��C�����Lz�fg)>��>��? ��>̲�=E�>������������yB����F2����U׾х�#�a�ʗӽ�1����;��E����>�"�j��>A�?�X>ǁ�>�9�>:!�=-�=7I�=��J�*I��
�>���>���>K�>'�D=���>?��>�������{�u��K彶B��s�V?�x̻���~g�%"���A�b�0=�XH>���>�3�eC}�^�x�_�>ɾ���设��i>�g׻���^�?�n@=�X��������8���s����>�^��>����N˾��A�m���AiK�?�>��<{=?�6>?��D?1`��N�?�A���-������(l����>r#.?��?�[?/tv?�Yb?���;����dW>����V[���4���<��ܼ:���N��=�$���4=)%:>�	�=:>�6<�GR�0����E��>Q'"?���>��>��h���?�5�a�rp�rÄ�G�=��F?�f?�@?��?�n>�a:D=���ܪ���߷�>�5=>A�e�&�w�崪;0��>o�> �\?�T?L{ͽ�Ŝ�#��=����>S$?��?Gʀ>�h[>xX|����qlӿ$�j�!�ソ�<��[�;�<�r�M�t�7�-�����D��<<�\>��>*�p>]E>?�>m@3>�Q�>�FG>y΄=F�=��;�R;r�E��M=*�G<3�P����UƼ������G�I���>��M��jټ�
?h�?����{�^�ǡ�Jz��򒭾 �>�2�>�H�>��>h�=A	�BQ�mL8�KWy�hS?��\?a.?��a�c�=��p���<���>���>q�>"�a�{2<�Ai������#N>���>Y��>}#��=H�oe��b㾬��>�k�=�x��[m�?�$y?�%�eu��N��g/��v/��Ƴ>�ƽ����B�=7x���e ���پ(�=��R��ۙ�p��>^ؠ?�����>G�ξ龥��;���S��W����=��'?�ܷ>U�=����!�,*ľ�c�J�%�E�>ni<���>��$?n�?�vl?�#&?�?�w���>| 1��t�>㪧>n��>���>�S�>��2>1��>���=�-�=1w����q�nU�<$O;�>��a>�h%>W�ʼ\TH;��<S=Z��<���<DO5�|%%��[n=TT>J�=��=�|8?�!?�[z�B������_�V<%a����+>t��=_�M7���>�m�=�`�>�K�>� �>Ѕm>��*��޾����e�=O9?�"?J7�>�U�=�N�=����D�Q��}6�	 %>1�e��V���澤����9ݾ_��>�	�>��>D.c>�s?ȋC?�%?kO���b���f��:!���A��!޽N �>���>�0>��Ծ̇D�\�\���E�Ъ+�[b��g ��f�=Ww&=m8=��!>���=���="�=��<G	�x\=<�=2m�>땓>���>{�p>���=+����� ��rH?Fס��N��O��Ͼ^���>
J=>���$�?�>��_}������;�|;�>*K�?X��?sd?i�=��V�LZ>I�X>%>�&<��>�=��
k����5>�{�=e�v�k��6�;�8b>z>SH׽�Oξ��㾹�D�i����N���J1�wˠ�������+�d���2��@�R	*=Y|��g���ƴ��¾��i@Ͼ��Ѿ�5��B����ġ?K��?��[>�{�y�q��+�TPR��R���.N����>��Ҿ�Փ�<<�<#9׾ǉF�\4ǾwdN�����;�~��>��Z��6��>�{�pf)�iյ���@>ve.?�ƾ�l��I����\=��$>���<���r��ŝ���,���U?9?e������f�׽�%>D:?�7�>/�">�?����;{�>[�3?�x-?����ܳ���!��"x���λ?v��?n�E?�Pv�E�D�E;�֥e��R�>iq?׿�>��{¾B\���>�>6?��>������Fۿ>��B?SZ�{W>2X ?&ۺ>𰸽!�����a�����+f�d�N>N����e����-�3�Z�s[�=:2q>�5y>��r�L�|��x�>��JP��E<�a����r�ʦȼ~M?��F��=�EI>�/>r�;�������������9J?4ί??�_?��?�þd��34��6>�j�>0g>��>�8���g�;^�>�?���h��������?E�?���?{�d?U����$Կ򑚿3ܠ�+h�����=�'�=xO>q�G�=dY�=�
=܋�V�+>��>�=�>Rۈ>��>F�G>i�%>�ۅ�!�#�P����}���X�� �5�!�'��'����J�_X�i��������á�6�ɽe�½&Y�G"�&Iϼ��?��>kO?3��>��>jw�>:�D>�S�=R�1�
���4�B�1��־R� ��������|U���t�&�нvࡼ:ؾ|�?K;�=��	�Dߥ>Z�>�9�<[��>��>¦j>7$>��r>#}�>�f�>�>:�%>	9�=jb�a\�>[��=Yv����s�JR��p��v���>���� �ý�Rݾ=���j����>�d�>c�'>w�!���9}���?Vz~�H���<�O���>��?�Iz>��=��=?�t�ȃ˽�<>X|>���=А��݈˾�Q!���k>���>^�ʾ�i�=��p>�!?�'f?�x0?��>7;�>|:l>�l�>j�
>�>�G>4F�>Z��>Z�@?`*?N?���=q:��?�=�p�=ތ4��d\��9��+�;	�-���$ӆ��!�<�=��;;M=�
�=������;H�=L�?2�>TMF>��>�_���M��!���xp��H��>1�=66T>Gz/?��'?��K?�&9?̑�>@��e���8��>����}U��1�����o&�>'=>K*�>"F=?
Rs>_'���>m�?�� ?�BB?��B?�>���>a̐������Կ�1*��g��~��R7��K�d=�z��)��<��F>͈��v"�/�>-�>h%�>y�>{Š>t �>x'>�o�>�>��˽wn�����=NO>Iw �Ә�<�㫨=NϢ��%I�����X�x��}��J�;���<�9�=gŝ<h?���>���<���� �A�M��� ���j?��>���=�,�>�X>N����+�5f5�Ϥ��c?��l?�X?����k��>b(�=�	>
ޫ>?��>+*��G3�.������JX%�8��<���>L^>=���D���4}�]�!�Z�k>���=J��B�?��M?^����.��60�o�������޻X9K�#���˖��k�s�#�g��������g^>�v�>���?�����������kh��0i��`����'>n4�;s4?���>Bf1��X �P������H���7�=��J��8+?�Ai?��V?�g�?��=?�oO?o�=��>g�j��>'�>�* ?���>���>���>(��>��#>�W"=rCr��3�������c���ޮ=B@>r�A>A";L1�=E�A��G��O�=i����m���C=Q=6Ly��&>�Xa>�^?�?����-�>jZ'>�����vS���?p�>ô�=�d���*�>��?ҖC?� a?T�@?�&�ɾ8�8����#�>e��>i�?��?�ul>���>]���p��l#h�_(H>]B�����	3���/��[�����>���=�s>p�Y>%;|?M�@?P�?\	̽ur���l�!��Fc��뤽�>{��>�Fe=�꾟�<���q��=[��J.�8����S��=���=-:>]�;>���=�*>��6=),����ѽ���I����>.;�>�� ?�UB>�w=FM��!����H?[Ͼ�Q��>ͨ���ľ����l�>��>�����>����c�Fԧ��3T�Aw>��?��?H��?sp�o#c�	��>K�>�\�=c��=�-ϼo̎�jx߽����6�p�ѾR)¾Ɯ=IV�>K�/>����߾�ѾG��qƴ������ݾL�C�to���VO��ܾe���K��D�<f�S��2���{�ۆȻ(o
�(���c	��◾+ؾ�Y�?d�?*$�2v>bV���,���侾�W� �羥b#�'_��l&>iY��xC¾dz��ױ�'���\�`�+��@�>\���ܗ���h���K���m����>���>�z���K=X����f=	�1>C<)���0���I��H�w��+>?�40?����݃�2��=d��>�d�>��>@�<����/_=� ?̷&?��W� 狿9ǎ�˹0<^P�?��?��K?��Ͼ��P�{��*�Ǿ��S>I�?�:�>,�s=�����">��?�Q�>�%>����(Q�������?8�p?����s>���>=�l>3�=�Fj�����F)<�6>L��<�x�k��v��X�L�Y��=���>�-�>7��������>����H��]B������`�
P=:;?��ξ?�>���><�'>(f1�{닿 2��N�%�XGE?�*�?��Y?��(?���	�̾$��9 �=���>D#�>9:�=�$���>bc�>��ܾ"~s�O� ��?��?�b�?8W?�c���п<��{�뾼|��7vH>H��=v�>�AQ�U��='�s�#���h/ɼ��>2*�>��>7_�>`׻>�^2>3R:>���d�}㹿�8�������� x[�!����|ܾ����U�lžK����O����R}[<�ܕ�7*��D���e���>_]1?h?�u�>���>�$�>�p��:B�X��֧��������oJ��Io��)8��Ԩ��r�����[*�X8?�p�>�~0���>����w��8�>Y��>t��>�)�U�X>Z��>��>l��>�g�>� 2��':���>�C>e���j~��fh���M�|5����>SV��+�P�P��NQ羚)|�zϓ>O�>��=�[D�pݗ��璿��?����0����m"���}���M>���>{!�>�(9>P�潏����]��<0,>��;%�s8��o�����=Re�>ȔӾ�'�=�3x>�K'?D�u?�7?��=}��>+'b>>��>�O�=	YF>8�M>���>�?�9?��1?T��>���=Z�\��L=�[A=K;��kP��������l
�P��<y�9�=�9=�Fq=!�	<�B^=��Q=������;��=�?�?ϣ�>Α?-г��(^�%]z���_�Fb?�E�<̘�>�O?��8?�?f�?��>�rz����C�/��Ѩ>?�½�K�a�-���=�1��vH�>́?�:?�7I> �5=�?�?��>�H?��9?�T>���>���݈����ſ6\/�+G���>6	2>��U<�(��dS����FBz��x��e�K>��0?�3?�.'?��?|Y�>l�!>��>���=��>ze����^�s %=`�F>�-�=����>�N�;�F3����vڽ�쒼�U����<%����ȏ��X?z�>�ң=�[�<s}�����mn�=0�=?h^?>'>-�B>��=K�<�Z�Z���:���Ӿ;��>�.w?�F?EB˾&H�>D��=���=��<?�~?o�=�$9=Y�����p ���=�?9I�=aY~���P�L�	���I>��>�V���ǟ?|R�?yB�Ì	<��@���������=��&��~�[־!,��f3�Bݾ`/Ҿ��ԾJ���@��>��?�VT��o=	6پ�]������ܾ���=vi۽���>Gؑ=��ھ.f���H���/��
b�ܙ�+P�>>No=��
?��2?�.+?�]o?�1?�p,?�5S� d�>Ug�=��>�r>��
?��?���>0�n>:��>�F�=��:���,���Q��=DZ�:�%>}�0>�<
>�F��>�TS>~&�=�Ľ��<�t��=U]�=�Q>�s=ax>4;D>FB?��?{B�=/j�>��;:���R���3�6��L?�(>��ڽ�'�>8S	?�??Fe{?&?ƅ⽡վvi0���m7.>\�*?�)"?�N�>�M�>r�=��{��G��\�J>��о�x��_�	R-�M"��c�[>N�>�~>��>�y?.�S?S�4?:0ٽ` ��d�g�f��bн̑Q�؎>��T>�Խz/��Y2���u�^
T�[k*����h�'��= ��<P�S��R�=`�A��>>��A�,��=� ӽ�����=G�>��>V��>��[>Ő�=ЁξX����I?�ࡾ�������i�оY|1�Ah>��@>�����?-�M�|��+��0�=�ޫ�>���?(��?�c?��?�-u���^>9X>HW>}Q�<�M;��#�k�����->4��=C�~�jC��ぃ;R[[>�z>�jǽ�Hʾ4l㾡�G�����@��}�i4�j�2�%�����`�¾*���"�>��Ѿ��6�d���08<N䀽]fI������ǋ� ٰ?N��?k��'�Z<g���1������E���)��B����7��������U����?�Q�N��� �D�*�b��>�Î�I$��lw~�)L[��}z�|,q>�?��j��!ӽ�.⾫\���w>�HN��K	�Le�����"�����:?F�'?OD��Z����U�ey�>l�>=��>`;?8q��
����=�/3?��?�<�6���)Z�>e0=e�?��?�-;?��x����ue�2�>�?
�;?2����I��:���>�_c>����>�(�B9����u�>i�q?-�N��M�=�8�>f��>� ����(
"�_�o��z�+cu<]K�=Ss���Ҿ+%�ty�<2��>�W�>�̈́�?9����>���I��
E�7�	��EH��1<c�?z�쾛�=?ao>�T>�,�����䊿b�+���B?7�?w�V?�,?ݟ⾉�Ѿ�˽;Լ=(�>3ԟ>l�=M9�X�>B�>�@��v�u�����kE?K��?m\�?�PU?5�j���ֿ����߭��派��>��=sOV>#�Ľ&�=z�<��Ĺq����8>��>m_z>�~�>P2>�^>z�=>k>���I%��Ӫ�)���=C�v��<�"�{kr��u�J􉾈�������Q¾�zj�f���O��i0�s��ZWۼ�:���D�>�n?�@�>D�?H�>,�R>l=<��6���"�����E*�f�"��
�~3㾧��O�=�0p�ϒ��B���x����>�>A��V\�>E�>�9=Ɂ>�ɢ�v����>�{�>��>"IU>Fܷ>U�>���;�� �O̊>�Ɨ<O���z�#�O�D���@e��P>��i<ĵ
>�B�vy��Y�k<k  ?8��>���>�x�i�z�����?
�ƾ_M���F�ϣ5�j>0��>��>'��>��s�̾@^�ڗ�>�o>S�#��qq������Ĕ�,>_��>����y&$>�-1>��<?:h?߽,?��>�<�>���>0��>8��=��4>Q��<�WP>π�>�!?Q�>?.�?8=���U7>�z>ᡞ�y+=�3��Ҟ�<;������<{)��A�=��=�j"=N{&>��:=__T=s�&C�<���>x�>�2�>�/�>�����j}��ߊ�碞��V?г.���>d�P? "?ʚ3?��?KR�>Fožl�ٗ��X�>��p:e�t���Y���弛{�(D>�M�>�B?xb��\������>�x�=dE�>^(?�|?j��</
>�M1���''ѿ��,��=�h��<t�]=Mc=+-��\��)7�=�~+��H%�9q�=p�>r�>���>�ܾ>Ӎ>{�v>?�?��>;黳=�ց�{��<D|h��5&�s���'�>�(x�����c&�3�Q��!��}��m��<T>U�D�C��W?-L�>��m<��<�`�ݾ6/�Z��>`�>���>�i	?�ۼ4�#��0]��5.�R@����>��v?��?�����|>���=����q??k4����NȾ����O9��=#�<'�>��=�Vj���!� �G�j�#�4?>ɇ�=oW8���?��i?\��n��A�(� J�A�(��<=���S�\�d2�Z�C�2�S�վ��ѾH.�����=�p�>��?�{޽�/�;��d{��ď�/����n>?��=���>�b�>&�3��"%�����Ά�a��ȣ�!�>�*��3?NM?�s??9^|?ƈ1?��J?�Ĩ�~��>���=���>͌#>��>E��>GZ?�w�>��	?�zL=�.����^��j?�w��=<����^>Ş�=��>�w>8G=M>��>c�;�<��
=ەV>R�>9��=��T>\�->.V
?��>�P���\->�ʴ�%���9b��?��_��>jS���-�E��>q�s>���>̳P?�t?".�N�辦����܊�>F�?[�?��?h��>*�T>}1��Z����=z��=��꾥E�Ň��y��n\�NY�>�;~>�B>��_>G�}?��A?�7$?{���#��nt�@,�Y����;�`��>饕>��
="�;w1��Tp�ȴ\���,��N��KK���=���=1N�=�Y4>���=$>�(=� ��oV�l�#<�-�(I�>��>aj�>%8>V;�=����ڴ��u�I?B����j�����rое�J�>��<>�0�$�?����}�H��o==�]�>nn�?ƴ�?�;d?�C����\>(V>�>4<(*>�3��@����k3>�5�=A�y�F����;�]>�)y>��ɽn�ʾuA���I��oɿ�k�����^%��.1���G���l���޾曾k>�(v��C�����l�� "-<��>]C���p.�T(��j)�?��?�t���j\��4��i������.�=�+�2=�	����֛j�Z'r��¤�4k��|~E���&�S�)����>~��x��r��>6���%;�k�>u�?�vV���b��i��N8�=5��>�͒��f���n�/����a��>T?d?�����K�޽R%=x+$>?��>R�?򪒾��c�4!�>�>>?���>D������ف����SR�?���?�C?e�_�"�
z�D7���r�=Xf�>�6%?:)�.��c?>�?[w�>`=�20�����f��,?��{?�e�y�	>{�>�FA>�듻֧�j[����<�>�J�=D�}������b
X=7J>I,�>�g�=;���2��>�^��Q1M��y>�3��W)X�3��<�@	?�;޾`h�=F��>#>�.�煋�,m��#[��fC? �?�V?��,?r�㾌�Ӿ���=�W�>�{�>lov=��>�Xx�>P+�>����y�������	?�Z�?N��?t�Q?��j�ܥֿ+��䎾��ů��>�=�7�=��M>�s��=Y")=c1Q=��ؼv2>�؟>��>s4�> ��>o�t>�6>���I$�Y�������@��3�����O�e ���h�&����=���o���>u��kѼqS]�\����c������t�>G��>}��>� ?��	?pK�=��<�;��P/�\X��Y��6��<���&؞���@�!~��PE�J���Mʾ���>�f> ��a�>��'><���~>�\N����XJ>�{�>w��>�|�=\B�>N>t�>o߽OĖ>��<㶗��J��O�U�~��7K<��8�>�]�.B;��G�Wm�����=�?��?���=h��'x��YG���g?l*��n]׾�	ȼk���=�'>Y�?Lp{>��4>���$ꎾv���'H�>��E>�hq�~槽�DC�$~��P �=�� ?jѾ`�=��>Y�?ZZ?�e3?Bu>J�?'�>dκ>!��>>W=u��<��x>��>{�?��*?��'?Na:=A&.�,I=$��A����D��� �Ek?=�|Ž �
�A�:�9MU<�=�����Ӵ<���<�X��錌;i�_=�>�>z�0?���>��k>U=���W�ic�������>��F>���>'�>��)?X�?�	�>��>z�Ѿ��ƾ��%��@�>i=Oy�D�F�@(���ܽ3et>��?��a?�g��C�9�J��>�>�>��S?�9?/^)>�7���=���0ٿo�{e,��߃�V��:�G�=��)���J��,�<1�N�מ?��ˣ=�Ȍ>Ӛ�>���>N�>�>@/>dG�>�x�>,=1"X��n�<��C=��	���;[��~!�<�g���p'��"��[�:�����5����=M}	�yoT�Ѫ?u�h>�!�;�J����I����Ѽư�>(V�>�8�>�?��K>�]/��E��#��~϶�#�>a�c?z!?�R��;�0>��=p�A���?���>���F�ߔ���孾[	U�t�M>n �>m��=�� ��(��/��d
��Le>�?=ZK� ܋?�Re?���c���E���$�Q��%Q!���o�Cf��iž#�H����i3���F��X�=�"�>�H�?�C<H���[Z������P��k��8P�=�U1>^d
?껬>��UK �d���p�.x���U�>0�_>�����0?�CI?`�A?[�z?V0?�bS?J��ry>5�A=���>I�>��?iA?�*?��?�?)�h�LZ����g��L$���=W@j���Y>�h�=O6>^h=�sr=m�V>"T>}�����<��=��=��k>&L>fR>f�>��>G-?��G���>++(=�ɾ�M�oV���>�v�=$�O�'�=Y�>�?�Z?��?�`�Tj�����|>�*(?)I]?{"	?Z��>���>:�����߾�ۓ<f�=�|�����R����L��q]a�A�>7H>�/*>P�'>�Gs?��e?:k?�w���ر�����R��N���K9s>�MA>5:=�cƾo:@��`���h�������.�}z%��j�=�5Ϲo�u<��=��Q=�>����2nټA{�=G� ���3L�>H��>�?�:Y>��&>��~���,��2J?F����"�RT����Ҿ�i?���>�U@>mJ�s?6�꽑�z�p�����;�*�>���?l��?jPe?�<��H���\>��T>�9>%�<Xr3�"#��^��
�7>H��=�(��Α���<%;զV>j�o>�=ǽ�ľ���ճH�@�ȿ¾ ���P��((���K�FV"��Sվ�g���̞�ô�}�޾�{ܾ0L��^Nu��=�B�G{&=�[���ɾ��?�?
�X!��7�
�ھ��:�hO�
M��@�=h0��A)�����`ͽӇ`����Lw�����"�:�>
B����cl���K[�B#B<�8u>y?A�,�������x��;?�'�=�� �������{�����6.?;?�f��X���]�=+�C>*z�>�^�>�/?-���Ȱ��@:J>Ur?�?�g��B�����N;�$�?'W�?��J?����13��+��kc˾�uX�$0?�*3?�N=#2G�(�>k�F?���>�������􌄿,����0?��?@Q�3�>.��>Dyi>Z����¾B��0�)��v��/�>Ǡ�>�"��ޮ���,�c�B>X"{>_k�>�=ޝ��̢�><'��1?��]3��(��8���߈:?�)ؾE�hq�>�z>�oF��0��e���
壽S+I?)F�?�O?{�?$K������uE�:�>oa�>$�>�+�=�;�`S>b'�>�2~��1�?���?Pu�?U?Vqz�?Gӿ��!��������=%�=��>>��޽�ɭ=��K=�ɘ�Z=�p�>���>o>M;x>��T>ӛ<>��.>q�����#��ʤ�4ْ��[B�� ���wg��{	��y�����ȴ���X�������QГ��G�]���T>�'�o�»>��?�f)?�r?	��>1�>o�;�>:�������=�pot���שž�oB���r=Y ��M�8�K��C���DA?�P>�V�=ԡ> kr=����3aN>�v�>!�s=Ea2��uY>2n>���=�?D4�>Å��[}ս5͇>�!>�U���኿t�^���{��Ƚ�5�=��T�.Tz>	�����A >��8?�y/?��z>�ϗ��9���.����M?mE������B>�U<�gQf>��>$�>�q�>6�;䫇��V:)�B>�3>�F���Ӄ=���9k�~����=�q�>)�Ծ�V�=�Ѓ>��#?a�u?�4?Hh�=���>��b>m�>Q��=9�I>�{N>R�>(?�p8?Ѵ-?���>k#�=Nn]�I,U=owP=�aC�$[A���ǽ�����C�f�"=������)=�6=���< H=0�L=O���0A�!�?=r��>h?�²>��>q�����J��d�.@ν��>}!��3?�O?nL�>�>�Ʈ>�4üиq�?j�ZR��e�>�J��JG�C���;�K�Q`?��4?�9?���=���=��>24@>���>A?�1?Ű>�b�>4+�o�$�׿�����t�D�=>Ґ�<>�=����)=X�=_��v��k��=��>���>%�5?��	?2�>��s���>R�/>�h=Ad1�2H�=*�Y=�A���`=q����=���%�V=gJp�O�J ˼�_=�  ��P��=J=�o?�ϩ>x%�d C�p�
�����Ͽ��?�K<>BH�>�M�>��D>��8�!FC��=0���(�>^f?=?����ߤ�>�����:���] ?)"?��%>ih˽�����n}����KG�=�0?I[�=�M��u}~��0{�9�}�>G�=��l/�?>W?{/���--���8�D^�>��K��=3;�殙��ʾ�A���T�M;{��Iк�Q�/>X��>�Ɩ?�̝���0��O������_���Ȣ߾�F0>��@=���>=��>�44�����|�
�v��9qǾ�x��A>/m�"�?�PS?v"9?��?{'?�<?��۽���>�> ��>}�=�H3?F�>r?]��>o��>F��=��Ž�;�.̂���C=�t+�\S>�}�=.B�=�=�UC>�_V>�b=�/�=΢j;�U���5<��=�P�<��=i^k>�S?׹?��:�2=�&����H6�yT����>֟��<b�f>�#>���>�]:?�h>�{I�b޵�2-���͵�=i�?[A?0�?�a�>�R����@���x�MH_>V�3�t �%=ھf���q���O�u>W�>`Q�>���>b�b?��=?ؘ�>��潴<���#��n�uS�;*ʇ>ԭ>�+1�i�����8`N���w��46��}*�x����+=�{�Z1M�j�=n��q�>)P��=�XF�|��a�>�1�>�ت>�z?���=e�=�!R�����G?�4�������~�N�=�*�>f�>I�����>����_T�a�����:���>Ln�?,�?�i?��ǰ9��=�>O�>e�X<��C>y�3���J�����&|*=&u�=������þ`�o��N>�9q>���������㾕6{�5ÿ����d���0� �ͽ��f���Ⱦwi���ق��D->�f����о�e�#��)��<���I�G���Ӓ�(R�?�ڥ?�������GN�u � ����󱲾f�)�ڢh�28�bli�"�u��׃�����P�14����夿>� �����:bo��7,����t�=xR/?����!�����x�=��q>���P��%h�[��q��j�\?:!?)2�4����E��,
>*��>���>P��>T���@$��U>�IM?�;�>l�z�(��%ဿ�8�O�?B��?&�>?���6@�G����[����>�?�	?�Gw���p�c4K��_.?�9?�l��~���x�l�jn�>i��?2����3>a��>d�>�B���Ƽo��<Y��fw��_l>�;���ΐ�m�A�X�>��R>:d�>l.>�g��Z�>��!aU��\P�����* =1�!>�k?����=3 �>�&~>�f2�A����喿q�>�ّ/?m˼?��\?�T?�پ�S��j��������Q>e�>f &����q��>^?�>�=����q�@�8�4?3��?u��?EL?��e��]ۿ&���&���CL����>&��=�\(>�M����=&4������󼂼�	.>�o�>�Na>/��>��g>�i@>�W>�˂�PZ#�䠣������?�S���ћ�#������?j!����W߾)Qҽw�0��	��d�N��j��t�a��>�>�u���?�o�>XxL>������pg>���>�G�SA�5h�'�!����
� �yb��Ju�Q'��*��?8ɽ��4= |�>V����>���>g��>j��=���>�>*��>]��>�r=_@>Hj�=H����>J7G�x2����>�J鏿�u;��W�>�zQ?a1>�����M�����̾}��=�>�>M8'=4e(��9�E����G�>熳����mk��ꀞ<�7(>�X?4��=+��=ιؽ�ͽ"���=@��>9//>R �=���������+p�>Ԋ�)��=]�h>�f4?Mh?�2?b�A>���>mO>��=���!:>��K>�ۋ>�?�(D?E-?<?��^=�v���Ƈ;i��=ހӽ
����.����	9�E��<1aQ���<=y>s=a�4�"i�=��[=mR
��w���D=ə�>�S?!?��'?7�'�bfc��LM�����@P>���>2Jq>1H�>}0?�<?��?rR�>1k�<\-��DF��?!P>[7>L�.���}�.����J�>�� ?Gd?�?T�w�:���ѽ��0=ѕR>솞>��?]��>vۘ>kb��B��׿B����7���ݺ�4+�@�Q��"��%��~�Ѿ���������Z=�&>ʜ�>��?�`�>��&>��>���>��j>}��<Z(��F��L��mD��)>�̓�4і�&@ӽL髽 ��� xF=�T=�U=���=��/���j���?�� ?,� <�l<��Ռ������3� ��>�+�=Hb?o�>��>�|�9놿�h�Ə��oJ�>#�a?�k?yپ���>�����+>�>um4>�q��⪽�̽頾�Ia>S塚xb�>�T�>B���կe�YO��.��
4>�D�=Q ��	�? �5?r�ܾ�m@�}���K��2�+e�>Wk;�\��CӾ(%�+���	�����������7�>ۿ�?Ԋ��	��>�L���x���ԁ��2���B����8�>��>>��>-�������ֽ�~�����ʼ���P'>��>�?#�D?��|?�j?��>-�=�<?����*���>��?v�?��?�s�>Cu?�=�c>��P�f
��kX����=u�H>��=��=�f��� >1��=��=��h�:}�L�����`=���<�)�=��=�kc>�?�,?�<�J�=���<�Q㽃ݏ<9JH>㪉>�������<?�>(�	?jJ3?�2�>�l@>�	��<*Ծ�, ��奺��>�!?�:�>��=�m6>7�Ҿ���7���j�x=�.��`����ݾ
x���+!��"�>� �>�C>և>l�|?�l?p;?���<Al�X�Ƽ;�35r�L >Ǻk>_?��>H�=��в(���u�a*m����d�Z�<R����n>e�B>5f�<�����=Z��=�䖾�h�=}2=�p�>���>��>8[�>�=:of����\�I?He���<�Ff��ºо~v��b>;=>?'���?t���}�$���^�=�Y�>�M�?��?�}d?o�B����a\>
�W>�>�'.<�_@�`�����P3>*�=�z��a��h��;!�Z>��x>(�ʽ��ʾ�価�J��2���O�Վw��w����{˪�`o��-�;�0+�.���&�ž+8����]X5�e����F��VD��B��'����*�?�#�?jgJ�YV�<�[�2P¾�ͽ�s�>�;ǽO\/�(�0�	ý��ϾiTʾϏ׾�tK��^U�+���.o���>u�����`���3�2�v>�|�>U�S?'���6�����Nx�=o?�<��>Kt�[;��Em���e̽ .?#�3?��׾W����P4�=�I>6�%?�L�>�7
=U��r�t�u�>��a?��?��e����Bb��f��CV�?}I�?N?�f���Q�|�!��0��h�*?�L7?��>��Ӿg䦾���;�3?�>�z�=��K�2mv�A����=?��c?��p�62>�1#?Z�F>o y�����Oz����ᾕ����>��ƽ`cؽv݅�?���o����>��>N"Y���ľ��>�Jؾ�5��\]�]���{.b��Ƭ=�j�>���2>m�d>�'�=�=�= ��W�������[S%?�=�?۟F?�	?Hp�����j�=�>���>�j�>�U>��F��f%>''�>!C�ALx� XԾ��?��?6�?�,?��c���ҿ�]���K��e&��kcZ>��=m >����ZQ<ݕ�ۄ/=u����pH>"��>R�[>J^�>Do>�rR>͝4>:����&�o���󲙿�P<�)
��:��uo��1�J�}�����d����;�w�<nr��u^=�����ս3�ΐþL�g>/j�>cM>�^?�ӳ>t׺>�����!/���/�s��=�B�C.��=#�\�r��89��y��A飽�!���	?g=W��=��?��9�.��=ՍG>��2>���=e��>e|�>c_�>.�>�>�u>_��=W>�Զ>6�E�������X�S}���,�<�c">��Y?�G��%0�3�B�۲	�I��̏>�P�>T㰽�������ȓ����> �B�M^G�Ý������F�=ܲ�>͘x=A]ǽ���㖾W���ëP=��>��q��Q�=�����ъ��3L�>�/��Ψ0>!M�>ؚ ?��j?_�?'E�=� �>�>�>���=��!>�h>>��>��?��G?RT?j~�>�l�=�v���4X<���=y�U�k�n�-ʽ����Vʽ�6<�qܽ!��=�>=�=��,��=���<�RG��Ż"7�>�VW?S?���>�9���n�_��j
�
�=(�>��?�4?��2?��>�w�>���>�IZ=� �h�(�>xJ>�Y9���F��Ĕ��3�=�$L=yy?�KV?�6G��ry�e�J��x��U��>*J�>�?��?75�>n-	>�m���ؿ��&��w�cLR�?.u<M��<� w��zT<r����*Ӿ����ܶ	>��>�Y�>ڏ�>�H`>&>*�P>:��>,Ke>��P=�	F>C]����޺7�k�}�=��-��ڼ/��m|A���8��袽&H|�E�?�?�n�:{��i��u	?_�	?*1�.4*�}�l�����F��au�>�B�>��?���>{��=֙��En�LN��������>*h?Ě�>ҩ���<W>z�T�PǪ=���>J�>��9>�W�;������c�=[d�>	�>o�>�����CB���V�����؆>�!�<% ����?��d?�B �(�d����t��$���p>�y�}�<�7;�z��z��x�:E�E��b���hV�>�Y�?����>��ھKF���0��T���t�)��m>�{�>�F�=� �==�&����O���MԾ��A�LV@=�^�=�?��?�N<?b�k?��?�5>:��q_9?_�@�<�?
��=+��>���>�L??��?��j=j�>��3�2@������M�=�Cs>�&�>���>v���٦?>�o�=���=��Fz!>�{�<$x���Rֽ9�����<]仨T?א1?_'%�W?�<K�H<�Za�~�ؽ�JG>�l>�𭽣i#�%ݼnjD>&?788?�?9U)>#A��6���rq���o0=?�`*?���>bK�=37�=(��x�{�%R]��a>>xĽ%c�����ۯ�����W/�>�>�'m>vX>�6?��J?��%?8����9�,"w�Մ>�&l�C�c=m��>�M�>Cr$>�2����1��Le���g��2A��N��8��[�=���=�<�=a}y>_X��	(=?��=�*��|��='�<�<�>�+�>Z,?��>��k=iҿ������I?������� ���о�{E>`�>>�9 ��?'��Ɲ}��ߥ�U�<����>%}�?��?��c?��B�eJ��\>*�U>�E>A�;<\$=�� �@}���Y3>>7�=�pz�Bd���6�;F]>��y>Q�ǽ�aʾ��"J�����^Ia�	z��Hg��sh���_a�7N���f=kn��j�&�b~!���S��J�!�=�,u`<�Ū��@��-�"�cz�u��?u�j?>��n��=��X�0��'X��*�@>�ܱ���J=ʻ��7^�=�|�F	�Ϥ��=H�O�
��|�c��Q�>����g��k(��7;;�`�=���>�o??�:��(���4�D�Ɓ1=��=�
�<��'������8��J� >?e�?�о�1 ��c��#c{>���>��>�:H�!�r�;��:b`>{�g?"�&?7к������␿����?W��?��M?�&����,��@R��c��*�>*}&?.�r>����!���ҕ���~?�+?fҙ��kS�����W�2��QH?�H]?y[{���Z>Q�7?�MS>������S������2T��M�>��*>=�������	}澉,B=Fz>5�>N<f��Ⱦ��u�>
��7M���N�
��T�W��ˬ=�?]
 ���B>�A�>�>�9$�^���V	����.�}�;?�h�?�Z_?�I ?���d��&,����<DW>j��>L��6@�FO�>[5�>�a��>o��5�0�?c��?0w�?6�M?�Mg��s߿!m��G?���3˾s>=Կ=�>S5�C��=�X ���'�|{���-�=y�>І>�6�>���>�Wd>G�1>����`"�bd���=��&49�W��Э�T/����H�����;sЫ�15���P
��f{ǽ���?�e�-��Ct>L��>��<=��>�� >md�>�s�Ɂ�N0@�
��=�L���6�"!%��*/����x���lQ�Y�<w������ ?0 �d>��?I�0�`��=��>��^>H�->,��>�'�>��>�_�>E5>��o>���=E��<d?�>AnK�*�����>�B ��ys�;�k�];�?���=����ľE�׼����=z?_��<���W{�f5��G��>NI�i�1��0���:�6M>}�>0O>K�J�߽�Ó��\����Z>4!�>=�O>�WZ=o4�n����C =2O�>mž��>�]5>5�3?źt?�P7?hsu=��>�3�>P:Q>�Rs=K*> \>F�n>�*?e2?`)?���>4}�=��x����=���=J�(�@~t�]��� (�����w��a�S��=�<�<�.<Γ�=`�= ��ދ�<�>���>�QK?9�?�?����c�9d�P��ћ.>�k�=ո8>�t&?�G>?��?�o	?1��>��n=ݾ8H��ע�>O�(;B�H���Z��8�_��>�8o>�# ?�F?5%N�.x��ʑ8�9�����>p��>0G1?�o?y��>�5=e���ٿ��˻*��c==���;�9��鯫�w?�4Ձ�>�љ�5�D;L�>V��>��>M�>j>��i>���>�l>��(�3 >B;��#"��w��m�=���<1=st�<��3����=�Cx�VK�lK�=�-�uC��#�S;�n?{�>ZP�`8e�Z�v��H��/��z~>�;>::�>WR�>���<A������'~h�5�����>`�m?�	?����>��I���_=9��>S@�=f0y=���C,)�� �2v=j�>T�>���>�u�OK`��q^���2��i>�4=d��@I�?�Q?08꾲�_�Oz"�])J����K�_=�B��t̽2����������	��芾 :��_�>�*�?�O?����>�JϾ�睿��V\����
�I�t=���>d��=1�7�LK���J�Q����R��Z�Y.>EV�=��	?�\4?�)/?�li?���>?�?�^v��|?7�>�n�P�!>a?s�>Q[	?�"?+�?��=y�:>�wI�Zǔ���_�r;�,r>?�>lƲ>��=�Q%>cC>N~�z�� �5��==ж��=nx�=K��=Yw#>��>v*?FL�<D��=�<T�?�8��>=
h>����ݴ�%�;���>���>P�4?G[?h�Q>�f���ƾ���%W=Y��>�B?l?���=��>EؾS���NE=.F�>RPF�)�����������$�>��f>*4~>L�$>co�?��R?"O?huh���^� ���'�1�vW��:>Z�?��>�>���,վ�=���P�b�{����C�K�R	>��R>f��=�=U>ښ/�j�;�	�=��:�6��,y����=F�>�
�>��>}!!>\?�=����E��	�I?}��5���-Ѿ{����>U�;>=��E�?���K}��٥�K'>��,�>��?B�?q�d?[HA�j����\>o�Y>%�>��;<�C�g��Ғ����1>8)�=_�y�����|��;	�X>��x>�ɽ�˾�{侰VM�����o�����0޾�����j/�D��wIҼ� ��o��Ϡ���[�D~ž����3��2ׇ�='G��	�ͤ����?�_?����-�F>�_����̾滾���>�ʺ���J�R���=��;�!޾t��f(�$?�u��{�%�݌�>����љ���}��)���t>Jā>��j?�t��������\w>m��=&�Q> v˾����������k??|�? Uݾ�e־D������>�-?��>
d�=0�B闼���>&tR?��?<��;*W��f���χ��1��?k�?��P?g����I�3%�����z�"?��?3/�>�g����x�˙={?G�>��>�nB��{���"��W9?�n?{@��;>pQ*?��>� �t	 �S��;,)��x�A��>���n��*�>�����2�_��>F˹>�*ֽ�՚�Z�>��!aU��\P�����* =1�!>�k?����=3 �>�&~>�f2�A����喿q�>�ّ/?m˼?��\?�T?�پ�S��j��������Q>e�>f &����q��>^?�>�=����q�@�8�4?3��?u��?EL?��e��]ۿ&���&���CL����>&��=�\(>�M����=&4������󼂼�	.>�o�>�Na>/��>��g>�i@>�W>�˂�PZ#�䠣������?�S���ћ�#������?j!����W߾)Qҽw�0��	��d�N��j��t�a��>�>�u���?�o�>XxL>������pg>���>�G�SA�5h�'�!����
� �yb��Ju�Q'��*��?8ɽ��4= |�>V����>���>g��>j��=���>�>*��>]��>�r=_@>Hj�=H����>J7G�x2����>�J鏿�u;��W�>�zQ?a1>�����M�����̾}��=�>�>M8'=4e(��9�E����G�>熳����mk��ꀞ<�7(>�X?4��=+��=ιؽ�ͽ"���=@��>9//>R �=���������+p�>Ԋ�)��=]�h>�f4?Mh?�2?b�A>���>mO>��=���!:>��K>�ۋ>�?�(D?E-?<?��^=�v���Ƈ;i��=ހӽ
����.����	9�E��<1aQ���<=y>s=a�4�"i�=��[=mR
��w���D=ə�>�S?!?��'?7�'�bfc��LM�����@P>���>2Jq>1H�>}0?�<?��?rR�>1k�<\-��DF��?!P>[7>L�.���}�.����J�>�� ?Gd?�?T�w�:���ѽ��0=ѕR>솞>��?]��>vۘ>kb��B��׿B����7���ݺ�4+�@�Q��"��%��~�Ѿ���������Z=�&>ʜ�>��?�`�>��&>��>���>��j>}��<Z(��F��L��mD��)>�̓�4і�&@ӽL髽 ��� xF=�T=�U=���=��/���j���?�� ?,� <�l<��Ռ������3� ��>�+�=Hb?o�>��>�|�9놿�h�Ə��oJ�>#�a?�k?yپ���>�����+>�>um4>�q��⪽�̽頾�Ia>S塚xb�>�T�>B���կe�YO��.��
4>�D�=Q ��	�? �5?r�ܾ�m@�}���K��2�+e�>Wk;�\��CӾ(%�+���	�����������7�>ۿ�?Ԋ��	��>�L���x���ԁ��2���B����8�>��>>��>-�������ֽ�~�����ʼ���P'>��>�?#�D?��|?�j?��>-�=�<?����*���>��?v�?��?�s�>Cu?�=�c>��P�f
��kX����=u�H>��=��=�f��� >1��=��=��h�:}�L�����`=���<�)�=��=�kc>�?�,?�<�J�=���<�Q㽃ݏ<9JH>㪉>�������<?�>(�	?jJ3?�2�>�l@>�	��<*Ծ�, ��奺��>�!?�:�>��=�m6>7�Ҿ���7���j�x=�.��`����ݾ
x���+!��"�>� �>�C>և>l�|?�l?p;?���<Al�X�Ƽ;�35r�L >Ǻk>_?��>H�=��в(���u�a*m����d�Z�<R����n>e�B>5f�<�����=Z��=�䖾�h�=}2=�p�>���>��>8[�>�=:of����\�I?He���<�Ff��ºо~v��b>;=>?'���?t���}�$���^�=�Y�>�M�?��?�}d?o�B����a\>
�W>�>�'.<�_@�`�����P3>*�=�z��a��h��;!�Z>��x>(�ʽ��ʾ�価�J��2���O�Վw��w����{˪�`o��-�;�0+�.���&�ž+8����]X5�e����F��VD��B��'����*�?�#�?jgJ�YV�<�[�2P¾�ͽ�s�>�;ǽO\/�(�0�	ý��ϾiTʾϏ׾�tK��^U�+���.o���>u�����`���3�2�v>�|�>U�S?'���6�����Nx�=o?�<��>Kt�[;��Em���e̽ .?#�3?��׾W����P4�=�I>6�%?�L�>�7
=U��r�t�u�>��a?��?��e����Bb��f��CV�?}I�?N?�f���Q�|�!��0��h�*?�L7?��>��Ӿg䦾���;�3?�>�z�=��K�2mv�A����=?��c?��p�62>�1#?Z�F>o y�����Oz����ᾕ����>��ƽ`cؽv݅�?���o����>��>N"Y���ľ��>�Jؾ�5��\]�]���{.b��Ƭ=�j�>���2>m�d>�'�=�=�= ��W�������[S%?�=�?۟F?�	?Hp�����j�=�>���>�j�>�U>��F��f%>''�>!C�ALx� XԾ��?��?6�?�,?��c���ҿ�]���K��e&��kcZ>��=m >����ZQ<ݕ�ۄ/=u����pH>"��>R�[>J^�>Do>�rR>͝4>:����&�o���󲙿�P<�)
��:��uo��1�J�}�����d����;�w�<nr��u^=�����ս3�ΐþL�g>/j�>cM>�^?�ӳ>t׺>�����!/���/�s��=�B�C.��=#�\�r��89��y��A飽�!���	?g=W��=��?��9�.��=ՍG>��2>���=e��>e|�>c_�>.�>�>�u>_��=W>�Զ>6�E�������X�S}���,�<�c">��Y?�G��%0�3�B�۲	�I��̏>�P�>T㰽�������ȓ����> �B�M^G�Ý������F�=ܲ�>͘x=A]ǽ���㖾W���ëP=��>��q��Q�=�����ъ��3L�>�/��Ψ0>!M�>ؚ ?��j?_�?'E�=� �>�>�>���=��!>�h>>��>��?��G?RT?j~�>�l�=�v���4X<���=y�U�k�n�-ʽ����Vʽ�6<�qܽ!��=�>=�=��,��=���<�RG��Ż"7�>�VW?S?���>�9���n�_��j
�
�=(�>��?�4?��2?��>�w�>���>�IZ=� �h�(�>xJ>�Y9���F��Ĕ��3�=�$L=yy?�KV?�6G��ry�e�J��x��U��>*J�>�?��?75�>n-	>�m���ؿ��&��w�cLR�?.u<M��<� w��zT<r����*Ӿ����ܶ	>��>�Y�>ڏ�>�H`>&>*�P>:��>,Ke>��P=�	F>C]����޺7�k�}�=��-��ڼ/��m|A���8��袽&H|�E�?�?�n�:{��i��u	?_�	?*1�.4*�}�l�����F��au�>�B�>��?���>{��=֙��En�LN��������>*h?Ě�>ҩ���<W>z�T�PǪ=���>J�>��9>�W�;������c�=[d�>	�>o�>�����CB���V�����؆>�!�<% ����?��d?�B �(�d����t��$���p>�y�}�<�7;�z��z��x�:E�E��b���hV�>�Y�?����>��ھKF���0��T���t�)��m>�{�>�F�=� �==�&����O���MԾ��A�LV@=�^�=�?��?�N<?b�k?��?�5>:��q_9?_�@�<�?
��=+��>���>�L??��?��j=j�>��3�2@������M�=�Cs>�&�>���>v���٦?>�o�=���=��Fz!>�{�<$x���Rֽ9�����<]仨T?א1?_'%�W?�<K�H<�Za�~�ؽ�JG>�l>�𭽣i#�%ݼnjD>&?788?�?9U)>#A��6���rq���o0=?�`*?���>bK�=37�=(��x�{�%R]��a>>xĽ%c�����ۯ�����W/�>�>�'m>vX>�6?��J?��%?8����9�,"w�Մ>�&l�C�c=m��>�M�>Cr$>�2����1��Le���g��2A��N��8��[�=���=�<�=a}y>_X��	(=?��=�*��|��='�<�<�>�+�>Z,?��>��k=iҿ������I?������� ���о�{E>`�>>�9 ��?'��Ɲ}��ߥ�U�<����>%}�?��?��c?��B�eJ��\>*�U>�E>A�;<\$=�� �@}���Y3>>7�=�pz�Bd���6�;F]>��y>Q�ǽ�aʾ��"J�����^Ia�	z��Hg��sh���_a�7N���f=kn��j�&�b~!���S��J�!�=�,u`<�Ū��@��-�"�cz�u��?u�j?>��n��=��X�0��'X��*�@>�ܱ���J=ʻ��7^�=�|�F	�Ϥ��=H�O�
��|�c��Q�>����g��k(��7;;�`�=���>�o??�:��(���4�D�Ɓ1=��=�
�<��'������8��J� >?e�?�о�1 ��c��#c{>���>��>�:H�!�r�;��:b`>{�g?"�&?7к������␿����?W��?��M?�&����,��@R��c��*�>*}&?.�r>����!���ҕ���~?�+?fҙ��kS�����W�2��QH?�H]?y[{���Z>Q�7?�MS>������S������2T��M�>��*>=�������	}澉,B=Fz>5�>N<f��Ⱦ�z�?9���?�3�I�!t�50�'t�=�2?�����|��S�>��>L����9[����ٽ�6?�p�?Dz-?�?��ǘ���
�qXF>b|@?d�?�̄�b͜�	�5�;ǡ=3ɩ��>����	���>c<�?�> @1OS?�6�+6ٿw���̆��sƾET�=�o�=_�D>�C��C�=�==`d��e ���9>���>��f>
t>h�Z>�=>��0>���������������7�9�
�t��:#������&#������1�������-�:iy�o�9�F�,��*;��5�,~x=jt%?��>�?���>��-<������4�$�ǾA�ҵ�����Ԥ���ڽ���T��諾'�a����-=?�~H�^ٽVo�>��꼈��<�r)>��>S�W>�)>{&>��Z>ʈ�>��-=��K=�i>Q����y>,��=Z����.�k�8�7�[�A�
�7 @?�\�����:4��K�EĤ�䝇>��?��O>a�'�׳��4x�/��>JD���^�?ǻ���A�<t�>/�>`�=��;h ���s��Mݽ.ι=J>}>�>��v�ڙ��$�A��=�h�>[<۾Lb>��q>�'?�x?�<1?�h�=>N�>�i>V�>/�=��J>5:>΁�>%�?��6?g)?ڻ�>Ώ�=]S�X�[=qQ%=�L�i;���椽&1�M�a\�<L�	��T=7�9=�<��)=l�<�w���D�;Ō=���>k9?o?�>�Z�>`��
�P�t~i��-�V>w]�:�?��>i�?)�?��>O�d� �ɇ۾�+Ծh��>��=۔ �x%��eI���]>���=�@?�H6?ь�<U^��v >ڞ>Cg�>h� ?��)?{��>�]
>7�a��N �Ϻ���Z���*$`=��>�X�>�.�x�=,�>NYH���.U>+�>T�>��z>65L>���=^��=��>I>�֟���=:��=����.+������6=y�=�'<�b�<��.=�g�v��`k�"��� n=_��<x?1?ZJ�<�6��,�9޾ò�����>���>b�k>@�>���=2�E�a��xL��V���>�6?̴?�x����=`��F����>Ҽ>`��<�/����r�����ٽu��>P6+?���>�x���9f��+��]"�x��>���=��D�f��?�9?�䪾�Mi���#*�O�&��<�s%��y��q���5�=�0�V��cM�*f���p=���>�?�������<�O�����P�$'���>�������>�q�>�J��S���=R��h.��W���=>�82?�̒=���>xQ:?.x-?�mT?U?��?Y`�(�>�25>���>�=�>A�?�I?�?~9�>��m>�x����5�ݢ��<�O>=�H�=��>��=OK=�,>��=ݜܻ�2��Q<��v<|��܈<[�=��=k�1>tJ�>`�I?��>a�;j�e��7�����>���;	B;��l�=�Ⱦ\�>���>��c?��w?�$�>�0��F)/�]�B��Ñ�� �? �2?�u�>^��=�Շ>��Ծ=x���^4>!>1��;u�e��Ѿ�u��#�<���>C�x>� 2>�>��?*��>��H?a
�>�!��
A�gA��K��u��>��>zF�>��r>��c{=�؄�Jr�� ����>f5��T�!����=�>���=���R�=�R�s	ֽ��(=�|�=�s����=���>��?��>>�7=�?r��("���\?��tS�؆%�*a��	e�>V�>���>|�2>�r;���)�]��)#��0/��?չ�?��?�zz?L�C��-���0X>�fi>�l�>jgB>����X��3>.
�={�>q�%��VȾ.�x>�
>Z8>b Ｉ���/P����T5��]���Ҿ&����W���u���������)O>������8J���=�=����A��F�������{��պ?�?�:����=�#�|bK������=w�qE=�˾�cy���p��c�4�������Q<���>��,���;�>2V�{΋�9)��;�⭂��0-�?�[ּ� ��RǾ�)>��a>�{�j��H��"u���j���8?7�S?V�1�: ���D������?]ܻ>8�?����0��,[?�{<?�F�>�w��B������7<P��?�U�?�>=?;�� 6�m���/����>��?�T�>WBf��V�3�!��P?`8?�k�>������/�"�!&�>t1m?.�V�i_>�[�>�ג>�t���x���C������n9<�D>8I<T$��.N�|]��2J�=#��>�?J>�SC�����" ?�Q!�{�K���L��a]�˶������)?����Ӌ=�J�>}��=� /�nY���$�����?<Q�?�#?f1?�?ݾ"�	��P߾�}�=[rI?:t?�֡���]��&>�,Ϲ�!�BI����K�C��>���?;k�?��I?2�V�AGӿ��>�����d��=^%�=�>>�޽9ɭ=�K=0Ϙ��W=���>���>o>8;x>l�T>֛<>��.>g����#��ʤ�2ْ��[B�� ���wg��{	�_y�����ȴ���Y���Ǣ���Г���G�C��T>�DGp�Ϩ�E��>�?�>e�'?��>|�лy"=�@�y%��7���h#�;�e$�9	��J�/��R��:���j����]� D?�#0���罟"�>���<��5>&q�=&!>*~>�=>�O>�=$L>���=sWt>(^O>߿{>���=�񄿦܀���9�F�O��$�;�B?��[�������3�.��z?�����>��?0V>��&����Ŕx���>lvK���_��Ƚ�$�څ�>���>Y��=_������vu���ŷ�=C��>sD
>��|�x��	?���=���>ň־�
�=�t>�_(?�w?-e5?[�=���>�!^>t�>鰾=��G>�O>�D�>�=?�:?�1?���>�U�=UQ_�*z=��:=��?��2_�4:���޼%F'�o�<3�0��vK=0sr=��< )[=�|;=hɼ�#�;7`=���>Y+7?	ϸ>���>3�E���A�J�B����j �=������>�w�>2�?�P�>�.�>�^�=�n��qþ�j���p�>��/>f�c��P��l �øX>XR>e�X?1C?'�P�����=��>o��>�g ?ع?*z�>1�>*!���]��'տ�w0���+�� =�0%��5�=�5���q��p<=Ӯx�f�=D#�>P˙>�'�>Kl>�K�=�="Ge>%�?zxr>��2���/�=�/1=wk�����;��3<*��=�����ռ��=EC��u������k����8	hD���?�n/?
�:��l	�E�h=Z@B����H;{>ю?8-{>�%�>�v!>��B1�AQb������P??m�?(�`��f�=�#�V.=��=1�:j6>7�=#�-�0��?�>F��>e!?PN�>����{�����"�I��>M��=M����?�9?dھt N���&��7� � ���W��rk�n��쇺������&�1���!�ɾ�Z��s=��?d)�? n�����=敷��2����t�S����=��0�
�>i"�>U�v�����G���䰾2��=�p�>S7�>�~���?,�?#kz?d�8?��?9�?���7R>�&�>p�>h�>�~N?�yY?ؾ?P�+>Y&F>�K	�[xžp'���s���<o�Q=�k>���>.H8>��=0��=��V�$�<���=��=��,�E$����<�52>�"�>��>�Y�>�-?�K�=�\=��ռ�U?���>�؇=l$�=�:;a����.=�Z�>��?�3?dS�>�a��W���$��7+����=Q�?�;?W8�>�G�<��}>@ؾ�ƣ���=�6>�H�yǻ���h�����$��g>4�=�>��>��T?2�>�!?ٳd=u<���B���߾դ�+�>N��>���>L0�>p��%�
��Vm�®{�� !��	�>ä���<��>�C�={�=�#;h+�=��ֽݶ�����K@�����'��>M
�>��>u�>o�_<#��|�	��1S?;�I�����M�ݾ�p�>��9>��#>�<�>TDZ���Ⱦv��t����}�==4?���?��?��?!?��;s��.�t>@g�<^D�>�c�>b��;rO��	F>�)=1%;L�.��Z(���E�'�_>c��>��F�����J�ɾH'a���h��ܮ�|1��ـ�I����������S���/:>a�Ⱦ��o���߽i�����ܽ��[�B6�����"�����?�ۚ?��I>o]�=�G��T��!7�τ�9��������?���8��h��Z ��)҇�\��̭�~�,�'�����>@h�E����\Q��?�`q��_?潀7/?N&뽝�������dp>�f3>,=�=��������]Ž��A?GEY?�G��o�i�����x��)�>�,�>��?�y��:�����>��7?��>�!��u���5��%HP��ݽ?N׼?�:?���T�:��ݾr���H��>���>k�
?�q��a��G��=��%?��<?��>P�
��ώ���5�Vٺ>�m?�s`��>�8�>��V>v ��3cb��)��h������>2�>_�o�Sa�*���G��>C�>'�#>
D]�!�̾P��>I@Ծ�h	��7�^�T�q�վsOb=I)?)T�ص_��qn>����R.������q���@��\h#?�h�?y$"?�5?�#�гE���>��$?!�?��B�-�ݻS�>>ЀJ>d\�J��A�)�	C?*��?�&@���?gWg��	ٿ�ᘿ�Pξg���>[�\>��g>����9�=��=q 2=�!>��8<�%�>�A�>]��>���=�k>I��>=���ʮ����~l��H�7�e�-��+�wҊ��h� E;�C����1M̾���y�<�|�\��ӌ&�LwW<���ɑr> �?��?���>6�=2�O>zM����$�����v-྽�1�g۾x�����;����Q^�j&����&���׾ه	?�E`�I����>D��=�> >B
�>���=N8>�k�>�Ѧ=h�1>���<�Y�<�T >�VI>1��=9�~>Ɗ=$-���`�_:�du�A���7:?��L�h���)4�	�����5�>%??�&d>�#��R��W�s����>ط��ϨM��`�S�"��S�>,Z�>='
>�h���@��B��񘽟�> Q�>5�=���eǠ����H�=�>����
9�=�Ӈ>�R0?)kh?a'?ױ�=Ϥ�>�A>���>���=���=���=,�>>�?��C?h;?�h�>��=.Kg�Z~U<G����c�b���c|����9��H��{�=!b_�`�=z<=Ms�<��<�M�<xz;q-�;��<}u�>ی:?��>I7�>}�R�N1J��uS��� �>4����>��>
Y?���>t�>�!>Ú����ξ�Y�N�>(�%>֝S�ʽu��]��'�{>̋S>�fP?;�1?1m��$��̍=㔬=�&�>��>"^?���>�4>�&��X���v��D_����G��=�N4=^�>7��>�9��~"=��=�i�>t����9%>a=�>L�>�kn�Mr��@�[=���>��$>�d����=���=�yJ�TU���#>v=G��
��h�B=�O	���ʽÂ,�W�?=`���4���
�?�?6�<����G�=��������u>d�@?��B?qH(?"�R>�?%��k@��e�m���?4?g�c?*�g> ��D��<Y�b����<}9�>)�?>�
~�� 	�B@>6�V=1�>�ո>�6�> w>3$��N�(�6S��r�a��>ig_=����m�?��a?�j�������!�D�(����<���l���}J��K��>7�ӆ���6�[�n����=V��>~�?0H��=�j��~ӕ�%�~��=��Z#P=�=IH�>W�S>��.�e����g �Q�r��!'����>���P�?T�o?T?Wug?ѯ�>��?跴��U�>S�5>:��>�2�>�.(?�~�>���>Em^>�]z=6f�L࠾����)����X>F�=�>�>0�/=��Q>�y=J>�:е?>������C��]ļ��a=b�">]�>/+5>j�8>�?�m�>>�1��>>ֽ ��˨�=9&>�7���I[���þ�����\>�?8i+?��	?cԟ=G������&�
���u>��?H�:?��
?����'�#�����tW�>�%>C!�6t�?�I� r�����F><�>�ur���>>7�?��h?�W
? ��=�Ԓ�z�*�+���X�=6�_>û�>��	?��>6�D�q���i��꓄�Ωo��!n�X�оVBb>�8�>�[6>J��<?�����>Yʽ�ظ�S�����x�MԽ���>��>�?���>X�o=�㾖�=��TJ?\���a)
������,	��>��F>��9>T&n�\YV>c������B7��JK=�d��> �?���?yY?.%����{�*>��۽TM��x�>�yW>(2�������] >HBŽz�޾��ﾧtC><� ?�?�k�=,������5 �=௬�6;�߱���c'���K�j�>�:��h��ۚN�	{���оP����'׽�Q4��ZؽFy���`�a�	J�����??��?>��=�So<s�K��C���갔�@��нI��� S�m���L���Cƾl���L�����C��>򁘾�����'��PP*�r<������<?2俾*eھ���BA۽�ĩ><�>��P�S�9a��	7�84]?!\1?�$����N���*!w=��>��>"�?Ң���N��5�>ӄ1?��4?5o*>����9H�����Y��?Cļ?J�I?ȸ�)P�?�'���x��v:?cu'?�-A?S*���S�+�Vn>�C�?}	n?�	=!�`�NZ
��?��f?˺C��v>�{�>�?����^�����F>�Ք��һ�c�=�8@=)�罉~��qw�,�<��>�s>�)��H����/�>��ЋC�E6W�I��G��;�n?v�c a�t��>���>��:�硝�k㌿�o���>?��?�Fa?8 ?K7��H���㛾�n>|9)?>m�>Z:|�S�*�p��>��W>z%-��=��+��S�0?�
�?���?+�f?hBm���ֿ~�����⾆_�u�r>�T>Bp>�����6��<�=��T=a>8��>ۘ�>v�R>m->-Q>��>y���Y �S���C��{j/�
]����^��9��?��	�C7���˾�j����T�mE)�?�I���.�(�p4��H�\>���>�x?�>�kY>��%>/��qi`��4�Z���(�b}��<ϾV�[�Y$>�">U����������m�>煠����=���>�A2�ZE=�o>��[��t�>�8�>|�f<Ѧ�=�n.>5� >�N>-��>ׇ=��>��W�{������#�P��>��
�=��O?�[�=1���D@\�!����  �>�9??���>�N"��&��9�J����>�
���]�;FW�=��2��%>nO�>~��>Fk}���V����dH>�>�}�>2��=�~8�]���K���]>(��>��Ͼ١�=[��>��(?=|u?�Z3?;gz=�>y�E>~��>��=Ch6>��<>�"�>l�?ۘ;?>4?��>�J�=l�[�-�<0=�&@��U8�5�ýT
�lN�͖<7@��P_=��a=���;Q�n=�$<=�਼�B<D�<���>`�2?�b�>N��>�ؽ���L��2�y"Q=�b����>aԡ>��>0ۼ>Ko�>�#e>��=�z�1����~�>�E>+�b���w�ASŽJ�Z>�7�=:�6?e\C?�PE=\�~��=�ͤ=���>���>��?��>g>�Q����p�˿�^���*��+	>)M�>,k׽�l��"��<��=>��=��I>xu�=3�[>�o�>f�>ڌ̽)e�<���>��>*|R>�����G>5x��;]�6g����=�p��(>]�r�N�����Z=�袽�.�1�=��7=�Co=z�s;�,$?�`?yTC��ϙ��]������_۾_z�M� ?L�>���>B��=ԡ��U�Mo�uܾr2�>?(�?�E�>-߽�hj���������=�v�k�	>�O�=���M>V^`=^m>3��>���>Ġ*�ضe��|l�j�bd?[=������?q^?� �!�n��>��%G�h���<\Fɽz�X��Ϸ���"��7�ZN�����2�Y�]w�=��>�¢?Pڃ�9S=b]���ؘ��xԦ����=���=:��>Q:N>|k,�����h���о8TC��Í<��>)���'?�ʌ?�>�?T>?K�>�J�?��#m�>KB?}.?�E-?t�r?��,?�	�>s�=kC��I~�aF���D(��ܪ��K+=�(Z���?��>��=��=��B=����=��M=�������\g����=���=꿸=�{A>S�?�E�>���9�=�����^���+���q>1���&ʾ������.<g
�>d$?�?_�:>Re��@|�t:Ǿ�~>�Y�>oD?���>�v�G�9*-���XT�=c_s>�����Ͼ�F4�WN'���|o�>���>Ǣ}���\>A�?��G?�;�>&k�J@:���n���%��P�>9_�>N��>���>�S̽������>��2x���Ȣ�!p;/y>��>�>>�>���<�f�>��ʼLA����Q�V�ȽV��;��>���>��?��?��c>RɆ��n>��%K?ŭ������۾���
�>�������Ό���ځ=1����������X*����>���?��?��1?�Q^�~��+��=��ٽ٥���c=F���bBY�h?���˖>Ʃ���驾�ा٨蹚�>��&?�$��ր������lM����0�I���$�׾�b���x"�����P6u��ʽUn>+վ	D���ڽ�a��-<����.Ⱦ�.��Qֲ?p5�?�E�����y�wqO��* �@�=o���2�	��Pw���6�],}��N��qI�3�&�lV�6V*�	g�>���Ov���a��p��y�\-�<dfF?M�˽!��3V��zF>=̑>��=��dw�~햿Gv���(H?E�>?%�@��<̽A���p�81�>#�>�̶>��=Ⱦ1�>=�G?)��>�s|�?B��~(��~^<�H�?`"�?�A?��v��Z9�\3���>�ŭ�>̋?z1�>)����Ծ�.Y�S��>6>?E�>8";��w���!��"�>��j?�H���z>�Կ>���>�M�M|þf 6��I����%�,��=�^�<��W���D�� �ؙ�;0��>z�>�De��G���/�>��ЋC�E6W�I��G��;�n?v�c a�t��>���>��:�硝�k㌿�o���>?��?�Fa?8 ?K7��H���㛾�n>|9)?>m�>Z:|�S�*�p��>��W>z%-��=��+��S�0?�
�?���?+�f?hBm���ֿ~�����⾆_�u�r>�T>Bp>�����6��<�=��T=a>8��>ۘ�>v�R>m->-Q>��>y���Y �S���C��{j/�
]����^��9��?��	�C7���˾�j����T�mE)�?�I���.�(�p4��H�\>���>�x?�>�kY>��%>/��qi`��4�Z���(�b}��<ϾV�[�Y$>�">U����������m�>煠����=���>�A2�ZE=�o>��[��t�>�8�>|�f<Ѧ�=�n.>5� >�N>-��>ׇ=��>��W�{������#�P��>��
�=��O?�[�=1���D@\�!����  �>�9??���>�N"��&��9�J����>�
���]�;FW�=��2��%>nO�>~��>Fk}���V����dH>�>�}�>2��=�~8�]���K���]>(��>��Ͼ١�=[��>��(?=|u?�Z3?;gz=�>y�E>~��>��=Ch6>��<>�"�>l�?ۘ;?>4?��>�J�=l�[�-�<0=�&@��U8�5�ýT
�lN�͖<7@��P_=��a=���;Q�n=�$<=�਼�B<D�<���>`�2?�b�>N��>�ؽ���L��2�y"Q=�b����>aԡ>��>0ۼ>Ko�>�#e>��=�z�1����~�>�E>+�b���w�ASŽJ�Z>�7�=:�6?e\C?�PE=\�~��=�ͤ=���>���>��?��>g>�Q����p�˿�^���*��+	>)M�>,k׽�l��"��<��=>��=��I>xu�=3�[>�o�>f�>ڌ̽)e�<���>��>*|R>�����G>5x��;]�6g����=�p��(>]�r�N�����Z=�袽�.�1�=��7=�Co=z�s;�,$?�`?yTC��ϙ��]������_۾_z�M� ?L�>���>B��=ԡ��U�Mo�uܾr2�>?(�?�E�>-߽�hj���������=�v�k�	>�O�=���M>V^`=^m>3��>���>Ġ*�ضe��|l�j�bd?[=������?q^?� �!�n��>��%G�h���<\Fɽz�X��Ϸ���"��7�ZN�����2�Y�]w�=��>�¢?Pڃ�9S=b]���ؘ��xԦ����=���=:��>Q:N>|k,�����h���о8TC��Í<��>)���'?�ʌ?�>�?T>?K�>�J�?��#m�>KB?}.?�E-?t�r?��,?�	�>s�=kC��I~�aF���D(��ܪ��K+=�(Z���?��>��=��=��B=����=��M=�������\g����=���=꿸=�{A>S�?�E�>���9�=�����^���+���q>1���&ʾ������.<g
�>d$?�?_�:>Re��@|�t:Ǿ�~>�Y�>oD?���>�v�G�9*-���XT�=c_s>�����Ͼ�F4�WN'���|o�>���>Ǣ}���\>A�?��G?�;�>&k�J@:���n���%��P�>9_�>N��>���>�S̽������>��2x���Ȣ�!p;/y>��>�>>�>���<�f�>��ʼLA����Q�V�ȽV��;��>���>��?��?��c>RɆ��n>��%K?ŭ������۾���
�>�������Ό���ځ=1����������X*����>���?��?��1?�Q^�~��+��=��ٽ٥���c=F���bBY�h?���˖>Ʃ���驾�ा٨蹚�>��&?�$��ր������lM����0�I���$�׾�b���x"�����P6u��ʽUn>+վ	D���ڽ�a��-<����.Ⱦ�.��Qֲ?p5�?�E�����y�wqO��* �@�=o���2�	��Pw���6�],}��N��qI�3�&�lV�6V*�	g�>���Ov���a��p��y�\-�<dfF?M�˽!��3V��zF>=̑>��=��dw�~햿Gv���(H?E�>?%�@��<̽A���p�81�>#�>�̶>��=Ⱦ1�>=�G?)��>�s|�?B��~(��~^<�H�?`"�?�A?��v��Z9�\3���>�ŭ�>̋?z1�>)����Ծ�.Y�S��>6>?E�>8";��w���!��"�>��j?�H���z>�Կ>���>�M�M|þf 6��I����%�,��=�^�<��W���D�� �ؙ�;0��>z�>�De��G�����>:H�=$N�GH����=�F�{</?�\�>r6k>�r>Q�(�-�����3�@eL?�^�?6S?d�7?G?����P7�����=���>�>��=O4�Ĭ�>D]�>U�龬�r�O��J??��?���?ުY?|m���ֿp���5ݾ�WY��)>��<��>F����<�I>'��=\�n=�l>�I >>Ȟ=e[n>�7�>�kI>�Տ>-ׁ�D,#�`��e�m��D%����AK��HC�3�߾�ܲ����0s����Z�ʽ�%��~T�����/�᥯�7��mxi<��M?L?�9��>-�	=-V�ΰ�����<��;:���  ��� ����{��@/� ���2ɏ�����(ǈ�o��>롤=���>?#��<���>/#>Ϸ��-�P>��7��_=�">/=��O>�ߕ>|��=�=�>�>�ҽ�낿Q~�IS�_P�+)�>8=?W� �%���&ԾhZR�~�=�c�>>�?�%�>��e���L����>����;�9�����=�B ?7�?�O��O�(�n�>gcǾ3�����>W�2=L5<�=X*���V�P�4>�*�>������<�w�%(p?V6�?w�>?��V>�?��X>Y��jV�<�\h>�H�>���>,I5?�:j?�'X?]nA?3�E<	�Z�ʓ8>wʉ<�;�d7�%����v<}T�2�@>��=��W>o?>�|Μ�y
`<�-̼M=�=S�i���>�?+�?���>Zן>�i��8?���E��^Z>+��=l˝��� ?�d?�b�>s"�>^Z�>RY>5ԫ�L>��.�(H?z�>jW��[6���(�=6�>��>IG'?��E?-N�}۾ip�=Stn>H�?s�C?M�V?�8���=������4tܿP�:�ߌ�F�d=O�D����=�#��s�=X0*=���;ҁ%=�-���Es>��=<��>��p>8q�=R]�>�>�`>��>�=��]��{��1�����:=��b=j|�@���f�=�g|�����뽌�
�Y��;Cok�ǥ?А?�<w��x��C��j�f������>Ϧ>��>n�>Z�>Z���-<I��5%�SSv���?i?���>g�r����=Z=|��=�y>���>!>G���($���j��n�=�׻>�?!��>0@�4�d��Ah�a����r;>��>Q�W���?i:N?����`���/��N��%����>�[���w��K�_��n��*�p�$�W�^��p�=���>υ?��
��k�>�����Ӛ�{���
��N�<K�1=�;?���>�Nʾ��<��n+��_Ҿ�:׭=���>��코�?��4?���>�b�?5"?�^ ?���T
?:	?=�,>,��>I�?�{*?9��>N�b>��?d��>S��>�]��=����^������ҽ�N�=X@?>6.��A�=e�L�[\�<ו�=�&�=�Y����D����=<=U=��[��=N�?�A"?�ڊ�8F��e�.>Y��=wO�=�4z>�hP>�Ƥ��*����`>:9�>
?vVX?���>�5�>Ś��$F����J�J>�@	?V�.?�i�>��s<�Ӕ��X��z͈��L>4IU>{߽������M��¾H+�wͭ>�p?�ؙ=ؗ>ۅ�?"�0?���>rB<�����h����{�l1>�1C>39?�=�>���=��2�LeK�7�c�DQ\���վo�XŽ��=��ټ����=��0>�h>��U>��r<�Ԡ�(�~;i����>���>=�?�J�=�o>3�,������bJ?�ڟ��]�3��*5˾��<�>��B>��b<?�5��|����{�;�M�>�D�?0i�?�=c?o�9��i���^>��W>B>1ǹ;��H�k1� ����+>r��=�kr�����״�8)T>Ԃw>\�ֽB�ȾP!�d*Z�Os��:V���I��%\�4&�����#�辅Vf�`<��_��9����3���o�+�M��sg;W{���Y���ƺ�%�Ǿw�?��?���=��u=L�R�������0w\>t��� �V����W��8����s����h��?�E�)�HB1�}	�>\����Ԉ���x��r:��.�E�>ձ?�/Ѿ5�\���8�ϒ�)��>�7��پO�~�������n���7?4&?(Ⱦ'\�� L�;���=���>�#>[5�=:f�VU���zO>�CT?s?�06�����f����=k��?�Y�?c�>?[*�h?��Y��@[
�E� ?��?gb�>�ԙ�7�޾� ���r?w�<?��>v�۾k
��.����>��I?��m�1�q>���>g��>���ƪ����,��k������!>�,<:>
�9iL�w�JZ�=C��>��5>ݿg���ľ(��>�C󾸻A�t�>�!D��4�>��<�8�> ��!>s�G>;[ >��#�mˍ�Ĉ��E�=?�޲?�
X?ߊ'?[�g�ھ��j���={0�>y�>�=���ɚ>)��>
sܾ.Yx��\ ���?�w�?�a�?�#M?�hk�>Gӿ��$��������=�$�=��>>��޽�ɭ=�K=(Ș�Z=�f�>|��>o>8;x>��T>֛<>��.>o�����#��ʤ�1ْ��[B�� ���wg��{	��y�����ȴ���i�������IГ���G�O���T>�%���S��=7�H?��0?(>�Ӯ>���>ް����ܾX�<4��h�P�'�~d:��N��p���b����=*���پ99�����>�s<��a>a��>�Ѝ�<>HŇ>Hv��c
>�.��%�M��>آ=UU>�c�>�簺p1�=%��>M�|��!c�Pd�f�W��j#>���>\�b?D-R��˾[4�[�"�~Ĳ��J�>~�?��?����'���m{����>�x���_���먾�	>��?_
$?�m�4�>Y���E��)��>��=_�>o'�<��>�_¾����b{>;M�>^�ھ�9�Ļ�=j|"?_�?��A?�'>i�?�m7=X/>��=�S�>ݰ�>#&�>! 6?��!?�?���>�5�=�|M�ۼ�0=�A��V���:󽡬��u�����=�ǻ�l=N�<6��<�>=�9ҁ*<�E���<�?�e?'�|>��S>��=u87��?��
�%#>�?��U?�B�>���>�?���>ׇ�=�VC>�']�O���}m�>%$��避��t�2誾�}�>z�>Z�?�T?�⨾P��~�=ʭ�>A�F?�>a?c-�?s� =�M½љ��u��C����<@�ʱ.��<i�|�#��9�a_���=�	�>?>慾��K��^�>HH0=�uc;��?Yʔ>ҌZ>���>X� >���=�A>�s��t�=e%��k�<K�*�*�=���=S�J=�td�=:���Ͽ��,ս��w�u�>e
�=�?�m?|�_T=��vX�3����������>hF�>c�>cq�>�=�J	�p�S�:�A��\���>Hwf?װ�>9�C�-��=�0��i�;�?�>~�>Hk>+c�����4��t�d<}(�>UF?��>~v�WB]���g��{
��<�>�c~=�0�深?�X{?��־�V�cV3���r���žD��=!sj�4G��:�
�En��t�%@�������=���>\�?E˟?�3���t�=Ơ��S��X��}O���(>��=A�h?nY�>%�=ƬǾ~V.��)��(D�[��=�*�>���=*<�>M�?�I?z$b?�?B�?B�y�?��=g�>9��>'?�3
?��>N�z>�U�>A:=��2�NA�����kP<��Ǽ\�=�>�Y%>,<?�=�6=<�<��7����8��<^�<N��<�Ӆ=��=�.>Ƿ?��>?Ѡ��<�ؼN��>���<�IۼA�b>:	3>Pz��{��z��>O��=�?RgU?#��>/E�>��ھ2-׾��/���t>v,7?�F?�H>��b�Bn��Ծ�/�M��>��S>U���j������,����4'?5F5>AGM=,;�>��?,I?��>���>'>X�A�����`��c�=/�܋)?���>~�A=c%%��pP��`�5�J�����C>K����)>����
B����>��=29>�>5v���ϽQ�W'<3��>N��>p ?�)>e�B>t����p	���I?����Sk���-qоo7�B�>s�<>@�1�?����}�a	��;C=����>��?���?�:d?��C��*���\>�GV>��>��/<��>�5��ބ��R�3>��=V�y�����֟;� ]>Jy>��ɽu�ʾ%2�rfH��T���m@�ס�̻0��Ӿ����̾.�>
������=ug��S������M����Ѫ�~��nח�^�o���kܩ?��n?���= O(>��P�{��	꾾��>2��p��u�澂E����!��r�Ee*�����4�u�i�	�4��}�>9���wy�`9h���7�7�=6)�>��	?���TPN��+�C��a�>�W�����n��'��w���BG?��?.�(Lz�X�<,�p���>�?>p���$�/�G8~�i�>�\?� ?`f��I��v7����)����?���?1�??���k&�N��Cx�� ?x�?��>p����)���;��?:�D?�%}>��ű����5��x?$�b?��=m3>�?���>�̽j����ڽ2m��L�5�ݚE>6FǼ�1
<C[���^e��T�=t)z> �>^j۽c닾UD�>r*龒[O�D�G�r������}<?���6�>Uj>j>��(������J�������L??D�?�R?	19?*����������+�=%�>�:�>D*�=8X��D�>���>�b��,q�<��?��?�X�?�QZ?�`m���ۿ�U����¾��ھ$��=�s�=��/>�����<�<��G���<`�=>Y	s>^8>r>�&i>
ZQ>Ho5>'���� �+9��'���#D��E�$-
�8�p�������d����!�þԃ��Q����ݽ��e�1w��y��R���	��R�"?:>0?���<�[�>��=����K��=�D���D��¡�f���+���ж���������o�澙־������
?��->�=�+?V�(�V9�>�_>� �<Wu�=[^H���!>u^��J�=�>=h�>\>�>�=�
?����z��WK��=�/��G�<qP�>���?Ep>�������:��h�:>j�>��?�Q+?N1Ӿ�����ya��U�>jǾme����m�������??7�0�1��=g~=>S���5����#�>'5�>�܌=��=���=@�����;X>&��zab>�X)>��J?�?>75?��*��e�>a�=UDP>�+�=*�#=�>15�>+��>xya?��a?�;?��8��U����=?�_<�Ӽ�n���;�:�������@e�;�x<IE�=��=8���wB���=���B����>(%?��?� �>��>{u\�u�=��
.���	>!Zp=~XȽ� ?)B�>�>4�>,�>���=��ɽ�u�����2?FAN>�3��yn��_o=8�B>�Z�>�o?��Z?�GJ�������>�m >�{'?�cS?�h�?��>X���ġ	��	ѿ�B�)/=����;��_<UwP�7�=��6>h�Q��ؤ�Z�=�7�<�a:=���>-�e>���<b�=D��>zUI>��<=��>�t���� �#���o�=��=���<�+ҽ�l�9��;j̄����4k�tUӽ=v��I�<�G?�,?�7�<��p��r�ƾrS��AV�>L�>���>��>�M�=A2�;�L���)�Q�Y��X?l�z?k?�h�c(>EI+<+8����>?Ã>'�0>����������OO/�馵>��+?�ŕ>Q�'���F���b�)���l�>��)>�|��-Q�?�܄?0�/�T�k��x2�׹P��	��4ܴ>��\>q8޽P��}'��jK�O�+��-0��@�;�)�>!�>���?��K�C,�=4q���4��ݥz�7����=Qd
=��M?١�>"�Z�x���������J[��_��=\�?��Q��?�1?� �>-�?�'.?�BE?�&���h�>�e
=K<�>y�>���>���>=U�>[�=>\�?sԻ>UDC>�3}��5
�3�Խ��P�����lL�>=�ڼm�Ǽ1t3>Y��<�bE��u��]6�;Z��U���ܘ<��=�����?�0?�*������&L�H��>�U�= H�>qç>�0��G���Tk�=7R�=J�a?o�s?«�>)_>�i��Uu��&����>��?Zv*?��>�=؋��L��G��t���f˪>���=�����5������-��>���>P>	>��>@�L?�=?B^?�{�>����+ՠ���b�\��>����� #?B�?<�n>�I�h(w�����U�K�揾e>=>􋽛�$��e���=��=+�>���=��.>��y�[�.�N������X�>w�>���>M��>���=���?�<��H?v���������;��$>{A>�E�;�?q�kf{����Ã;����>'��?��?$d?S�A�u����Y>XW>��>&I�<�.1��U�������=7>��=�[s�7���%��;�U>�f><Զ�� ƾ@���'�����c&��|���Œ�(撾]Q�*Ѿ��z�+�v����Z�����2�������m�̴����v�z�5�!S��吣��'�?���?W�e�&�=��5��V�x	����>��ؾ�"���ǣ��#��泾�3��l���OM�������x����Ȩ>Z��W����v��(7�Tb����u>�?-?�ʾK����� ����;�H>�d�<G�ܾ�g������/I��eG?*&/?W��Ph;�6��<�=���>U��>h1�=	J��o�G��6�>�F?ۀ&?{��$u���#��L<� ɼ?3��?*3@?��R��(A�����^��?�O?6��>8u���Ⱦ"����c?o=:?R(�>� �����m�> �Y?�O��ib>��>M��>�x�R ���YN����{���<>6��q���1j���>��g�=�ޜ>��u>�{T��R�����>>�N�N�6�H��������g�<*|?���D>Ti>ZS>��(���'Ή��@� �L?F��?��S?�b8?�P����������=5��>
Ь>X��=X����>7��>j`��rr�[���?�H�?��?<NZ?��m��ۿ:⨿�JҾ6�����>4��=�2>�ѿ��|�?{̻��F.> �T>�d}>"ZB>3��>��>>�;>x=P>����K�*�����QD}����m�m!�Ò��*
��^�������P�v��zG�.|���L��%gd���X�x��T��9Z(>�h8?�a?�w�>r�>��=qJ'�J���5�Ӿ �����A|�����lX��f��}І����<�5��p��x�����>�(;>�=(��>�M���>�T>(\��L>�=��
>tī;��1>��?=Ӣ1>4@>3a���a�>g�b���W�7�Q� pw�{qh��<kx�?����\��ʾ#2+���;Ԩ�>Y?}=ax��ɣ���P����>�'*�9v��0پl��=���>��0?y�2�D,>*LL�m��o�4��	=��>K2��"M�Z.�F�y��ɸ>;G�>����*]�=��f>�:(?�G{?��3?��A={��>sDu>?��>���=j�=>b�m>�@�>F�?\�8?�0?	P�>�	�=�`�΀Y=l�M=)�3�B�)���轄U�������<.�,����=i�?=�K.<��j=��$=�7�� �p<��=gZ?2?�+�>�>��<=އ5�8�C���D��t�>�?0�k?X^�>-2>���>\O�>E��>���"Tc�؋��ܖ�>/\=�pr��L���c5�3ȃ=
�>z3*?�?�^��վ<�>���> ?��"?��o?�X>GBk��tɾ67���R�R��b��;�>}�2<F��=�'��[�i����=Pď�l1�>֒B>4<)�Y�A�>?^?�S]=�>Ć�>|~�>T{�µ��{���=�t�=�3�T�!���Y��ZB=.�O=��	�U��P��Ka=��=�j��?��?�`K;yl���������nξ�>���>��>�?vR>���\D��{,�x�z�u��>0�x?�"?<��=�=�)ֽ!:q�й�>y K>��=���������2]��>�>N4)?s��>_l۽0B@�$A�\� |b>k)�=�� �
�?ȁh?�S��
���_�o���Ҿ�CU=9�b��E�?��!����:����5�'��<x^>���>�?��c��=J�<��Q��\w�Z���>�N>��w>�yU?u �=�A���t����6�|!W��z�=vG�>W�=hE�>A��>W>�>�[?��(?"�?�J���
?��=>��>�w�>���>r�?��?Cc�>ŀ>&% >V��������:��=�M[<��>HMB>�!/=�)=��<�=���=�;=��Q��.$<��<x��؃�=*�>Qc>��?�^;?=a���������=c�=;��=��*���>���>��e�q꾽fc�=�x^?�X?ß0?�Ӑ>9��H�6�;�得�>4?�9?O��>RL�>#��=?پ=���b=�h>����ʤ���ƾ��ӾDlþ���>��>y��=�0�>Wc?4@?�&?�(��b~C��GY�gS0�U)>��a=��?Ͱ�>]��$;�����]�a�[�ɕ���*>&j�.>kE��^Ӎ=��>j&��|��=��6>BY�=��:�����2�<��>���>(L?��>ͼI>�⮾����I?�{��?g��栾V]о1��%�>�<>����?E��E�}�����4=�'��>��?	��?3d?�	D��)�Q�\>TV>��>c�/<�~>����m���3>���=�|y����}g�;��\>p7y>ƙɽ�ʾ2%�7^H�i󴿮\�lh$�l�S�@i�����N~޾r�P=�����K��z�����<���&g�הN�J6
�/����p������?�g?���>x�N>%�X�%���Be�>̾%s�H����2Ӿ���D�
��F=Wξ-�[�|�+���J��>/탾D���Y!��+�*�'~=��>�<#?��оv�Ѿ�����K��;f>��;K��������t�L�o�i?`Y$?�cؾ3!��}_"��Տ=�8�>]b�>�o�=�6g�i2ӽi�>�@9?$?�F��w��͊B��.�?1��?��@?�P���	
��	��D����>d�C?� I>y苾����O��e�>��;?�J=�96�G���t�?��>;�?�:��OEV>L�$?E��>0B��z��*�=�)��,�=�ܞ>V� �e�*>"����\���	�=�Wp>���6�>̶>�_�>�c龧�M�/�G����~�K�~<=s?>��.>jh>�}>��(����������jL?g?�?�S?�8?Qc��u��v�����= ��>:�>Kӱ=_		�Yѝ>���>�0羬r����?�:�?Ic�?=�Y?��m���ۿ�d����ɾ�۾��=]U=v<�=�)j��M��Z�>�i7=������=춝>@͚>�q>u�=��=>!&g>B���k�&� ѥ������w?������n2����_��uT��|��$���";H����2ͽ3b���u�Y��L3Z���Y=͙-?��*?LF=mt>M}>��-��
�#Q��^Q��E��Q)�q[$��������]l�t�[����������>����?��>w�>��?��.��æ>	Ʈ=I$'=�RR���=��j=���=�Y0>i�=���>�z>��p��?�������n�F6���S�zep>���?�A�����h(Ҿ�^������?"?��$?���>��&�`է�!R��*��>U03��U�{��o�>S�>�4?~�L��X�={ D��Oֽ�_p�*)�r��> �|�A���_���t��>�k&=14R��,G>��=�Rx?�A?юd?�-�����>n�>()�>Ɇ�>��w>l��a5>H�U?G�`?�/g?�n_?T�<!7����ҼrO�:����阽Hҽ+C<ς`�n��rJ�T@=Q>B�>��4�d�<����!=����"\?�%?��>��>�<��X���L��A�>�!f<����X��>��7>,��>��>>�>��*�!
t�++�%A	�O)?�rc>����E%��]�G=6��>�m�>��R?G i?�ľ"���>�>�3�>ۤ,?��Q?��?�@�=�4��#w����c׿'�<�-�9�5%z��.⽏x��Mվ�b
��E=��@��m�=�^!�cs>i�>.Q'=yS8=�`�>`�>3@�>M�y>I��=���=[�=��%>6�����V��Y=���=<�Ƚ��=�詽�D@�J5ؽ�����:=?�����>&-?��=N=#�aٹ�����))�>�\�>偻>Y�>��=���:YQ�v5����*??-n?"��>�3����=��3<h=t��>�I�>��>*��I�>�(v��Xt��>6�-?�l>C_����L��J�����ǎ>�}>I%L�u�?��?�G�&�סF�+�9�����>�M��ι��x�ckL�����z�e�Z��犛���W��u?�{�?{K��0E�<v%������q���h�->�<>��W?��>q<.�H��5S��@��\ح�2�={��>� ����>D�>��4>���?�#?��J?�Ts�1	�>���=�
�>�\?��>i,>׿?8*?��>D��>R��>x�Ľ�����@}����97,������=Jټ�s��L�M>�"	=�i��c�����%�=j%�ZDm����>�c�>M�*?a�O?�$�b ��e�=�3�>CoX�~R�=�>+���dd��>e�{>T]?_�.?8�>C��>�Bx��"'�3�.��=�)?@�?��R>��>C$=�����跾ߖD=���>��d'�yV��x���X������>�(�>�QC>���>�r?�AH?F��>�N[<�Ѓ�+Ǔ�0��{>o譾5�??�
?@|y��~,�����M8��5~�o���1�<o�2��bg=6L>��=�3>��>;�S>�S>;T��_�U�h��sYQ����>��>ż? �>YH�=�4������b;?�B��� �*�v�ٽ��5z=��>{W(>o�t���>����o�J���-5�)_�>�e�?a~�?N�r?��!�Y�@���>K�z>1�>��=�MX����=w�?�L�Z>3#�=sN�����7�w=O��=f!�=(ڴ�і���4��MF=��x�S�(���Z�9���N��̶����~��ǟ�=�g�w�X�}�4J=u���E���Ⱦ@7��܀����?�o{?fE>Nˢ>w�q�>�F�����x
?���X�SD!���@��{���0� ��X����
�g߀���)�4�>ͱ�����E����,�Mi��l��>(�)?�s
�o�r���־Tsr���=��{�=s���������˾��Z?e�	?���_~��k�����ݧ>��>xl��)8�$�O=��l=�E6?UqI?�'���������;�?���?��O?w4���M����!���$�>�)?7�r>�ӭ��p�����>� g?@�>��;�xA���� ���n>��$?\���`�=�N�>���>R�ｫj�[ħ�bl���2&=�u>lXE�����I����j��=��>>�S�>P�K���6y�>�P���N��HH�LJ�q��ի�<��?���>�Ok>,�>��(����"ꉿc~���K?���?."T?��7?�O�����*��� d�=/�>���>x�=�j	���>�{�>n�羍�r��R�v�?��?:��?��Z?��l��˿Ɲ��R��!|�����>�c�=ݪ&>��3��>K=���>q��� �;)����>7��=��l>�Z>oВ>I�>��z���$�?Q��;��I�@V�iY���'�eܼO*�$㟾�R���l=��[�.U�;�����>���i�k��[<>}� ?��>r�>m@�>�<>𣨾ܥ��P��R2����1�_�þNo־
3Ͼ���Y&���½�:Z��*��<徥Y�>�g�=�(>Tp�>s䚽m��=C|�>sfo����=O0>$�>���>�#>��>Gב>)�,>ޅ����>=U_�(��xxh���h�(�ܾzU����@?�c���΢�Q����|�p�<>��Y>�v�>y>�v3�ϵ��*�g��?f�D������zľ*9��Da�>�,I?�?=q�>V�>䦘�lP��y�3>N��=KD�;W>3�%���>���>B&�>��IA!>Թb>��0?�f�?�??TG��>���>M��>{{�=w42>�4	>Vߑ>e?��<?Y�"?��?Y��=<X~�}�#;mx:�m>n�hR½{�˽9�!���l��i����<��9�=W�`=�7�<E�<=�/=j�����1=��w=��?��?� �>3?�>�]��d�O�&�A�\_�kӊ>$�I��>�$b?"��>�"?/.)?��=|�Q? �8����>hS<66Q���m�}�r�ǽ�>���>3�?�q?���z���`ˁ>�>w�?ky2?���>r��=d۾�[
���߿l�[���@�j�>��X�-���AK����:�=�|��dHt�uw���?p�=�om>���>�H�>_z)>e&�>V��>�_>�>.d!�A���9���7�=�E�=��N�*Y�=JX����/=�����K��K��g�x<�z
?>?1�=]Q=H㘾�,���c�i��>!p�>���>;�>�Vt�ذ3��hz�A�I�Q��YG�><Gv?�&?�$���Lp>m�>�8��\?�� ?�/��XQȾ1�վJ����S�،>�V?�3R>9���bP�tWj�7��MC�<<�=����ے?Op?���wWj�*8$�$�N�<�-��==���}Г�����۾�4Z������ ۽�pw=�]�>I|�?�O����t>Dͽ*"��bԃ��w�� �9>�6�>�8:?a �>�:˾ ���t���i��0����<,��>��:�W�%?��H?�E?��?��?w0A?�m��m�>K�s>��>��;>���>/W����>���>}@�>���=��K>�C;��޾�X��r۽�w�=I,>�d*>����\ݽt1B>8�=��=�j�<��=���(:���=��=�>>�?��?��A��k��N2>mr佱G���:�>���>c���!۳��Y>"��>�?Pk?���>�c4;�T��86�+����>���>�?C�>Ns=w<�<��M�$pU����4>D�B��q�/�C8��а='>S�H=�B3>���>�5c?(??�d"?�g����2�Q�o��++�8�u�=��>qk�>&��
m��"�I�Ё��\��*��,>0*�x�<���=�x�=�tQ>c��=��=�C':���=~O����=t�z>���>a
?��R?�ȱ>��=7� �����P?�U�����c=X��"��5:�)T?B�/?�s�>w6?�
��I��jl���[���>�k�?	�?a��?��%=�e]���?�&?��>���>�4�#zx�ZR�َ'=6b�=�9V�}�x������=�Τ>r�Ͼ:�G����3�=<a����5�5=4��C���#���+�C���R�뀑�
����<b���׾ut�������1�;��"���.���?���?_c�<̧�<�X@�D�5�u��l>��"��, �
A�������c��C��1H�����p��(:��.��(�>q*���l��gȒ� ?B�����J�>ڋ�>�5��t~��v��3Q� ��>�ٽ���r���I���ޏ>���Y?|g?G2ʾˤ��g�>���=Eֹ>�S�>�K>v����hм%L�>�c)?�U�>�+R�a���p���w!=	�?1��?��B?�q���4�m���c���-�>c�?�@�>�R��1Q���Z =��?� ?��(>)������+�9\?�|?�~|�H�|>Һ?���>K���Y����߽�'�±�=��0>X������g�ƾ6ؗ�љ+��}:>�>9���ǉ����>���n=?�D�G���VH���"> 
?P �XϜ>d��>u.=e�)���i����`e4��=e?���?�=?Ժ?�s��U�y�kP>M�=P�=x(6>��2>%\5���?�l	?�!�+����"��g?+�?} �?��P?٪����տ����O��P꥾�$�>�?>��>�U���=��
>P�A���?�>���>�T�>���>��>"��>�>����<I�?���/��1�)�5���F��٪�ER�~�-�����ӫ������d˽����CO�<"������$�K>�+�>?�'?k��>
�>��>lt�=���D�jd��R�վ��)�E
¾���c	�{'���a��3U�Y����ս�4��$t�>V0�=��S>��>x�6=T�T>{��>^�m��#(>�>Ў>L�G>�,:>��v>_�>�D>�t >�#^>#B>�Cs���H�[Y�A���y��r�?�6k�B�X��"��;��� j�>
�?�WU>Ĳ!���������?��o���ξK맾�1��9>���>j�=ʩ�=|"�г �h�=Z�>���>�������Z��f�ӽP*h>!	�>9,����c=H�>��,?��a?��+?2E>���>u>��G>��3>-�>`X�<e�C>�>?�0,?�T?&�?As�=� ����G��D8��׈��>3��V=Á#�4�غ�
>$�[=�5�=�~�=F��=q��;�6>,	��&>>!�0~�>��,?B��>��?D彭�=�/W�h{�v�\>ԕ�<���>a�>��?g3�>a��>���5�b��A0���w�> �`>��@��K��`�=I��>�!�>\�?U��>�>��U���ذ���l>..=|6�>$��>�g�>
�=#������ɿ�Y�E��G�>��>ĺ+>��
�t�dT�=����Y~�/��ph�=�C?�.&?\�Q>���=�����"�>��>���=�Z�=��ĽS��4�E��=����U�=���ڇ�=�)ԼE����y=� ����p�z] ��5|���?�z?(Nx>��S>�w���4�)��/?h�>d-�>�o?2>�4�|� �'c������>X9?�?�N�c��:J�=�=�K�>��`>��=	۸=�]>��,���=���>>�?q��>���9g���.�*��˻>�_�=�E�=$>�?�h?����M�9Q����B'���&��e�7ƌ�_+I�[[.�m:U�ܾJ���8�FqN>���>'Ț?n2�ݶ�~���E���^�������>�捽���>f�>`��@�˾���z�Y�&@�������,�>��=��>�?�?qDQ?T�?`0?�"ɽ� ?�|G>|R�>�¡>�?<��>m��>�a>)KN>a��=ソ�� �����(�3��住���M6�=�v]>�y�;���=�#�=&�=�9�z��DC=��;ҫ�<VI5=F
>��#>._?��7?g����x���=�!��c/=��:�/>l�A�A^�����>H4�>Pl?�t�>(�������lگ�v���5�>��%?�#>?s# ?���=#�+=������U�L����=k�R��邾M�������������>esy>�yF<�9�>+�3?�U1?Ζ"?���e�������)�D�>uv?u�?ʔ�=W��r׾wI��tP���*����=�J�g���P�;Z+���3�=H�=��X�c�X��V�I_���U=��μE��=Z=z>�r"?���>��<���Ӿ��Ǿ�@?�	]��܋��2��2˾����;��=�O�>q��e"?@=+�����t�¿��Q�*�>)��?���?�?<f���?X��j�>��>D;q>ѕ�=7��
{�:ƽj��Y�佊Ӿyþ2���F�仧*>�$��_�۾Վ�o�Խw����������^��}#�����>�����Q�����k=7���ظ��9N̽@k�?�4>���<j#������8
���?<E�?��A>�<�9m��w�_���/>�7 �]:��:ܙ��k�]
2�����M��3�þ���7<���?����>0~ľ�{��-I���Ba��
>;�>�=�>հ�Ks'�}?+��NO>v��>&�>Ρ��ŝ��Ή��#F��.???]����������>XLM?[�G?)�!>�s��$펾QA�=A (?"~�>��X�nv�������R����?��?� >?�d��=���:�`.Ƚ5t?1�-?���>\c�<�M������?�G?l*G>2�	�6���i	����>�Dr?
�0�2��>��>���>��R=[����ɽK�U���V��
�>�>�=Fh��% !�E ,�UX�Ņ�>W��>IQ�=�$��^7?��.�z�����,��N(���>�P�>����)�>E�O>��>k��h����{��^���,?ɥ�?�Q6?Gz?n<��,�ӽ���=�<�<�F�<#�$>Ow!= ?���g�>?�?'��刿�Kɾ���>��?���?�,?����ۿ�b���<ؾ�ξf�=���=s8>�bG����SK9>�~�=Ϩ߼7�m>T��>lD�>���>2X�>��g=��>Ӓ��~�'�������̽�>G#�N�$�}k6�hV�D�x�:}���V�Qk��]�[�T���Q_=�T���`�{�(���V��?r�T?��0?�%?b��>v��=�����\���^��s.�p�o���ƾ�� ����b����(�ý� 0�~ޣ��k���ζ>}�=O�<O��>��=%q>{�?�~�=R7t>(��>0D�>��`>�=v>��k>�\�=~1> )л��=��.>�{k�Ff^�V�K�+�l�Sq���?_�W�����M�'�C���(ҽ�F>�?;Gk>��Q�R���X��R?a36<x�q���	>�b1�%��=�=�>�� �߽�����,��==�j=�W>>%�M����?�m��=`�?�֚�e��;��=�?PPn?��6? ��>��?���B��>H�v>���>h���>g�7?�d*?q�>C2?y%�=A߸��J��i3���$��;��
~=8*=a��i1�=��a�/Ns=ub?>�o";�o�-Í=`�/m>����p?�>1v�>8�>���������h�,�>'k?+<���p*?�YY?=i<>�d?;�>�þ�
w>}j��a��jf>VZ�>LP�`���(>D7�>�}�=؃|>��Z>Y�=�ڼ� <&��=��w>l:?�h?�g�<@��<I_N�N���w俅>V�Շ(�L(�=AӼ���ZBg�3v<5�%�l� �[Md=+O�=��$=���>S�?2�>dv=e��=�V�>媉>�L�=s��=ڡ��q格�4۽��=	�.>��������=��,��0_��y����D?����=�R��#?�>��>��<BY�B���pL��#?ɨ�>$4�>|�?��=BU����Rur�9A�4��>��-?5??0)��1E��={ϣ�.��>7[�>x&��'G\�	$�=����<m\?�M"?�%�>����27�olT�Ă�% ?�	>�Rw�Ƿ�?R�c?�����ý���ߙ�#K���D=S��o���j�.����<���¾�q��E9�P��>BG�>SU�?J����v�=`@���m���P�ۚR�Jg>Qi��R�>Bx>Y�ľbǝ�(��!��0��==��z>���$?��?�P?&��?�)\?��R?<���k�>݁>�^��� ��iJ&?��>E�p?�?5i�>��Q>t���M������0r�<ER_�����#=��=1Z=};Z8>d�=-l=s|�=8;>��>��>�wT>�5?��X/=?1?W~?��ས(�=G��v��^��E�9��>V��=w"*����=�=^�4?]9?(a=3��=�{�V�Ѿ��Ӿê	>�c?;�7?_��>�U�<�~�=�,{� �/�@��o���K���^��?}��X��8��+�>��6>�?t=��k>||?��@?�*#?q���ʢ/��ev�1�'������h����>��>S^�=p�ϾC3�Ĥq��J^�.?0�lD0��E��=�S�=n{>�3G>�3�=�>��=ͭ�|�˽/d<�FǼk��>�.�>��?�Rd>Oy=�g���)�c�J?o ����㾎Jþ۷�o�ҽ�z*>I">P���3z?��6�Ft������L��"S>�X�?��?v�w?B�i�0H��x�>�>>��>�fc=�7���RG����< I���mپB*���.u�f�=�V>�8=������꾽`$<y�����-��|��~�Ą���@Ⱦ4���gԼ,:~�[qK�j���D��w-r��k*����y�_�>U�
���1�;�^�?��?�&&>�C�7KB�� ��;B���>��H�,�U��J��������8����&辤����<���R��8�%+�>�xm��g��B$F���[�����YQ=�*.?6�����O��bo�	B>=U�;�F7+�lԏ�'�����>�h�J?D�9?�������C��p�>�?�#G?��|>F�Z睽��>#?!\?~!���|�YA����=�b�? `�?�I?�yq�}�h��B4����l�	? &?y[�>~�J�v�ƾ6 ����>B4=?q9>YY�v3n��5���"?E�\?8f}����> q�>TM�>�!��Ϡ�����$*"��+��kL�>l�������r���g�(�=F=%�>�)�=[a��2 ?��#�b�{���k�d���I�0�iv7>.��>��پF�>��_>���=|���^t����H&���Q?2��?h�J?�@!?~���*�܈=��=舽(3>e 0>gj��6? ?��"�|
��mH龸��>k��?�e@4&?�N����׿
s��������¾&�>ܽ�=�,>���T)=���=SȺF-�g
>2k�>�%�>f�>omh>�Y;>c3>dw���%��j��<F��OWC�m�e�"�D!��/��*<N����Q���R���ͩ���)�q��_�@���Nw���lf�j�>Q%?��>/��>��>�'>ӈ��$�}��H��t;P�K����
N0�g6���.T�w7�X��k��&���r��>�s>���Sݬ>��b��ȟ>R��>N��=��>�>�a>,�`>�͜=XW�=�ӕ=N<�>
P�=��z<�&Z>ft�+��!_7�E@�������-?^9������n�T�þ/�V�]�m>Օ	?e�>���3������I�?��(����7�O>I��=��b>�0�<�FN���<�w�F���=/2�=&!�<���=Ľ��9��~� �tN>b?>�������=�
 ?ݿa?��-?d]>D�?�^s>,��>��>��>W�ZN>h�h?�4*?�(?�g?bWT=���[
�4�-=kĆ����=2�m���=�,���`<��Q=˗>��>�>�|F>7��=y*�B>~Y�<>6�>� �>)��>G?�s��0`�� ��y�>���>�>0�X?~�?
:�=��X?��>`К=����&�.s��k&�>M��=2R�K�_�)��M�@>�8�=+�>�?C�=kmU����=ku}=N��>��>ذ�>U�>j���b���mӿz$�+�!�=AO��݈;|�<���M��1�7w�-��������< �\>��>�p>qE>��>�<3>�R�>�HG>kф={�=D(�;��;c�E�˗M=5
��?G<#�P�Ċ��$ƼE���)��ƐI�h�>�<�T8ټ;��>K�?�z�����=�����1���޽J?�>
-�>�%
?`��>�n���'1�FJT�T7�˺�>��-?w{?r� ����tl�x�<��l>Y 0>��=	�>��M=�%���o>��>�n?޸�>�����2�(-7��>�����>Fb2=4�%���?`?���`��W�"�.��s�%_����k���þ��ܾ�%�#�K�y����-�V�\���P=��>XI�?�f ��<�=-o�tƟ���4�%�ٽw+6>^~<&�>F~�>��[��5پ��!�I�y�j�� ���I�>�����0?�|?�&?ي�?��\?S�?�{����?�`J���=M`u>�?�
�>P?=�?_�?f�?���@���M�����!={����V��ы=�>�G�=PDi=��^>4o+�5~6=���Y>��p;s�S>iQ >�[�	��=�?�B?�$��ޑm=X�=��H�	�h�?��S�=t��Tɘ��4�.�R>�y?�m'? �m>�*2�g���Ǿg��(%�>;?Z!.?]=(?Ϣb=����
5��}A��̀������"��gо w��6�/q��;��ſ>�J"��o>��o?TE,?�?"?��*�2�|h�Qx��)�<�[��X�>O}�>�!n=�K��D� �7�m�*K��/�*���S�υ�<�)�=b�=	H>��o=�=�	�Ϭ��^1��ȧ��-���>���>�C?ŚM>��<d�������yN?c�ݾ؅��Z��U˾̖���>��=�r�R�E?V���we��j����o��=�i�?B#�?rx[?J�M���1�/y�>��>�ܜ>B7�=�T��vɀ=R}���߼҈����ݾcq���-.I=��>��=�}ƾK�;��g��ϿՅ'��-�X������`v��֋��.��X�����=��;kr����^�zL	�(�<-���� X�(����¾�K�?���?�2�=�uG�[^��������J�a>ż���佒Ӥ�;qF�v3K����)~>�Ǭ��$\#�[Q�/D�p'�>i���h��*�Y��<C���:��L⽦9?�4��>�j�2򫾏�>�^�>ggI��E����ɯ��_���??��;?��-�����j��6&<��?W�W?��K��F(�r&�q	�m�?��2?&���,���m��H�f���?�
�?6#C?���o�Z���9�揾�J-?P�:?4�>,ٴ����.Es�yC?�3z?��>�9
��~��G�R��k0?(F�?��E�=���>�"J>�|=� O��AU���p��I���=A��=֪"��˾:ku���=L��>���>�?�=w1ݾ"2�>E~�&G���3�5��~r1�^Q/>�?���*��Q>4>�<����ek���&��9?D��?cG?A�?�%�U�����i�=�y��=��P=�����>Ka?���Ċ��R��<
?f��?f��? �L?�����ܿ�%���N���ö�&ή=��=�O>��9�'t6<�.=p|6;1��<%�>2�>���>)_>��D>R�>)>����� �s럿+����?���û�����@��qe�O��OA��������~f��熽�GC�$�	�u�/��[Z����>�?L?I� ?{O?�\�>��������D� �� �2��G���m7��%�������˽G2��19Ծ�`R�UǾ���U�>��K;P��=���>E�=b=>���>�'=�7>��R>k�?>˰�>g` >��]>�&>��\>W��=�X>5P,>�倿`�t��e-��P��
^���0?)*#������1�h`O� �(�b>��?�=o>2%5�eD���9����?2�=����w�o/�=u��=��>*>aD���v��\3x��4~<6��V�>v��S
�� ���v��%�=7�?�ؔ�mWT���1����>�ρ?�}a?�2s��X-?�� ?@�>��=�et>��?D(>��5?f�&?��u?�?x��=�j������m�F9����,>������<IB0�&*��:n�{3>kv�>`����L>�ƿ�m}m��͟=w}�=_?�L?���>���>۵%���G�),�@L4>�h�>�o�=W�?h��>r�s>Se ?��J>@�c>:��=h�žT�׾	��>�Y�=sC���\��	���ҋ>8��>�"
? 4?P#�<P��A�=�<�=,id>6��>��$?<�>S��=��޽�!��VԿ����yξ%��Vo��Q�t=�����D��'�k�kK7��r��T�<��p>-'�> ��=O�a=H�b>h�=�?��%>b=B>��q>�wؽm{�<og�D�=qY=��<a$^��'����w<�v�]�s������ɽ�x.�QX@�qa?��>�}"��3�<(�Ͼ*y �t����?�¬>�`?�?1��A/�D=2�T�9���D��^?A"?�>��A��q�wT�=�� >��>6��>�t�=�@��TW>�	>3�ϼ#s�>N^>?U� ?*��<Pn���Z�=~��p ?W'�=2��:�? �a?�.
��7g��=�g=�J���;H2�F%_��u��g�"�ٜ:�v��b��8n�c*�=��>�d�?}��sS�=m���\J��浾�e�=k�<��>3$+>�0s�ퟕ��3��:��o��{��<f�>,ۯ�cA6?]c?��>y,�?�F?�h�>�ei�x��>3��=��>���b?��,?n�\?���>GϞ>!�p=�=��󔾫�������O�[�#��7�؜*>ZkB��Z!=���=4��=7�����u"�=Mz�<�E=��=��>����?+�?��l�b�=0��=
.'��[½�>�m�=x�G�e:��o� =�=(�>B�?KΤ>�(=ݾo���W���>v&?��@?}A?%���w�Լ4�謾#�7��'��ʾLs��ܾ�j˽��G���H>	���'�='�Q>��?ʃL?�g8?s_=4����{�&:���	�RWU��R3>E�M>Gھ=�-�#��v�b��*`�)�G�Pǣ�����<b�=�8Q>�$d>�.�=|��=
%�=�k�M;����=�J�=�Q�>�Y�>fh�>�c>&��=2����M�E?�`�����>������3ʡ����=	v�>������>z[k=
c��ŵ���X�#��=;�?��?.�Q?�)���z"��rS>�m>�a
>���<�.�T�i��N�vc�G�=���7��ı��(>ּ#�=�����e����H`������Q��3����2��O�/Y��u�M٠�^+E�_
����.�W���v˜9"�?��#=�7�����T�׾�1����?���?�߼��J��-��T�)l��D�=E��������L7�����[h��l��猾��6qY�P�%����>�s��Ņ����x��G�%�{�l�p�>����'�����g�>�J>�����C��p��Tv���cԾ;'F?I�V?�J_���پ���t ֽ��9?��G?���=��5�C͆�vƨ���?�&?��������c�m����NŠ?3�?��=?�־.{K��� ��"�>=�?s5?��
���z���<��.?;,?�I�>93�$��-�1�h��>�x?�B�SF>
k�>F��>�0=����G�
��=�j��@%1��r�>��b����Q��$@<��>n�>Cw���+��*�>��پy�P�Z�0� e��=�
�:a>��`�<Ԝ�>t�>f-�퇚�S���/����y-?9�?��?[?@=��m��.f���>r'?��	?���S�ƾ�g�=�*<?Ry#�up������?|�?v��?Uv?�T=�1ٿa�� ����Z>Mn:GLY>] <��>9O�=�ɡ<	-F�ۛ>�&�>.�&>#��=��u>��o>w(>ڭ��<3#���������1�t0��5ؾ�.�gY
�q�[��'̾�_��~���O�½��$������)˽�2���߽;+˽"[�=�m
?��>�'�>ڕ�><C >�{ԾL�7�妫�S��e-�I��}��Q(��������<�C�^������I"?C���I�B>��?�^#=�?=*؆=�ۈ=#':>Pfa>3x;>m>��=��=��=�Z�=�Ǝ=V��>��^}Q�~�_�%�@�?��F��>�t?ߎ->a!��FD�{\�8����?68V?���>�w'�IZ����f��>uI��=W��m�����>ʿ><��>1W[���н�����~=�5�>���>��7>%9��;���B���>��>j,��9s�=&5J>�N?��A? [/?N1>&a?���=�V�=�����<.�=uf>�,?�
]?^gD?���>� �=�j)�c��`�c��B@�z���w�<���;�떽?
I��.�OĽ_�=K�=��=���=�Cz�K��;>�?�H%?���>��>�\��#(���K��5}�=��	n�>��>d�>e�>�<�>�k>�a�=E������?�>�[=�[r�/W��,a�����=���>���?�A�?�}|>������s�qB>�s�>�A�>b�?��>��i����=��W�����L��@����=��ȽC��=	?V��h�;�D�!�1:n��>�A�>~
�>�����ż=��>���=1m����>�{>�xX��;�=���;/�=Vc/���׽\?���̻�A�I�=K:��wP[=�-�<�lǹ��B����������?�S?�	�<��F�s���ȶ!��Y���܄>��)>���=��[>�x�=��L�"�}�h���=),E?6E�?���>)!׽m\ǽ&̉<��;H9>��>ۡ*=� ������.v�6B�=?��> �>�̗>7��<�2�q���5b`>ɕ�=��%����?cPh?����T�������N���'�^��i	��@��,_��u��u7��)ﾃV����c��>�E�>�q�?�	ľ�`�>����z���WWb�����Q��=bGj����>�XR>�������u1�Q��� =�u�>:+�>��ͽY�;?�l?��B?DU?�/�>9��>���cO?o��=��>�=X?�@l?��?g?�&k<�Qʽ����Z���o�*��课�M�<���GR>��>�~�>g�	>��=����P�v���Р=�D�uv�<e�>Rc>��=���>m�?nM�>z�=0w>b�8��*�����>Sw�>��=dݴ=�s��V��p�>�PZ?7iJ?A��>�&�;.��9+W������>��?m�R?��>�u�=�6���lB�h���eUO�|�=�X�=H���!�$��
�ze$��9a>[��>&[j����=0�?Mo}?��f?(���z�龅�����:�)�=�R>R�?e�>9��>X+�k5	�*��쒿HxJ��}�����*��=�$>6�s'�=�3�<d.]>�I�<�g�=��ʻp˖>���>�v�>q��>���>�l>���B���xO��5B?��侘�ؾaA��� �<]��>���>��2>;0���?7)p>�^�ib������?�	�?�?c ?�B���ļ�,9>Ε>�O�=�{������w�=��H>���>q�>,p	���A�Y
=��!?��>��>A'žU�@�(������4K�b�羲"���E@�M��7sо���E���ý���?S����:����������������ǜ��x�]ޱ?z��?�A��:��	�4�Sq���:�>�����g<�<Fƾ�������B�ཱྀ�0�@�:���7�V��>�k&��n��#wy���4�����>�;�^�J?�$���X���2�=�&h>6t����Լ��e�'m��sp?CTc?ӻ���ʿ���U�n�ռ� �>�e>�Oc>�m���9�8�0>��+?z	I?�O�a���E���ֽ8�?5�?�G.?G��YV�5��x��yp�>Y%c>���>bjQ���R��Sh?;H?s�9>��Z���d'�:��>
�{?aͽ�>�?���>'�Ƚ	A�	�(=x��,[X�K&�>�UY<�h�ӎ����D�L��=Yg�>�}�>ZM�b�־U��>�1�lW�Ve�_��HB >�&>Q�>Z��[�Mi�>��>�0�+���m?���7�4?A��?��x?3�?��'�T���D2��W-�>�o0?��?����N�GQ>��>���v�4�E���$:?n��?n��?3�H?FM��ܿ{�������0��xP�=����(�=����><��>	�>k5>�\�>�<�>ĩQ>+�=���=��>X�&>�����$����Hi��i6G�;%C�� �g����g/���վ� '��ݕ�����i����>�D�O��-5��
�,g��d>p|e?K=?9��>|E�>���=���.���1�����o�������·�_k�������<��Ҡ��C�@����0?��=�"�=���>�<�=E�}>��>@�4>�>o�>�z�>��=��ռ?�;;K� >u�&>a��>}��Jg��_~�!�����Ǽp_�=��B?K�~�=R^���,�H;�wn����>�E6?���>������f��J�>�����l�_��e~k������> H4>/�%=A�ʤ�Ԩ��w�>�Ǒ>��=�#н!ǾUY�U�D>~��>%���2/>�>Ɋ?�[?0lB?al>�S?\ϸ>r�>~�:=��=��>�n>t�!?��C?(�*?0��>zE�=�NC��|<��W�_��҈=�����[��F|�謁��=�˽3�u=\	�=�_>��@>�ݶ;����;n�d��>�	D?���>+	?}5V=�!��'�QOy�A+>ѽ���>j��>wMd>U��>�M�>�b>
>E�\�[ˮ��Ȱ>��
>�d��Vx�̛D�{��=�V�>i�3?�;?��->j]j=�==�	y����>�~�>W)?n?��D>�艾u�^̿K5��b�����;WZľ�!_�w#�=!���>��M>�>R�?<�>g�/>�4��a��m��J��ʭ�>b�->+�=ꌳ=H3u<Ww>-��<���={s=N��&�d��8����1���̽���
CM=������)["=DI	?���>]��<�_��='�<G�ͫ���?"��>�>�>��?t�m>~ �^����y�0�þ@&�>��{?�0�>�d�ɇ�;��p>JA�=��>>F>:�,>��z=��:e	t�,Xp<
�>�-?��>���ر8���x����q�>u��=���=���?!��?���?���@a𾼊R���&�:߼vO���˅�s����+*����Q�!�����<�*�>'�?���.}�=�O����fm�3	ݾ�[�=ً���)�>�C�='���A��j��R\<
O>J�>���=�{�>w�!?��?Ц`?ek?� ?��8��>�:�=�>�>��>�)?t�?�u�>T��>� c>w��<e�X����6O��\:�<%@:�TȢ=�6>�h>!�<��=�:R=�L�<�Z�����;��6��_+<�dG=!�=8R>ݑ?`�?��K�*<�N�=_
 <h�>Ŀ�����<e@��� �N���>+>�N?	�l?�T(?�-<��������7��G�>6?��l?��>��_���'��X
�Uȼ��>��f��S�����C�̾2=žW�U>���>�l����n>2�v?ϵX?�5?>��=�] �ؿy�7\�93�=�U��`>�}�>���=Y���G�t��j����P`>���+XS�m���'�=�1>���=�@3=�k�=�j�=Tz��.�%=O�f=�^�>���>1�>t�.>�o=L��{q�2?�ၾ+���'���8��9Ü>��q>�+J�����^�>�-��zS��4������)�>h��?L�?��;?�w����>�|i�=`��=�Xʽ���i������(8V>S�>]>���x��X���>{��>�3�<��ؾg�3������:3�V`r�@l����־<����� �P�T�M��������5�0ͯ��p뽿A?�̬���H�!Ө�j����?�a�?�Zr<
���4�cC�tX6���8<��m���9�9�ݾ�<S�Lٟ�͈����	J����!�Z���J�>�#�Yv����s���7��O��=
;��?����Oz��(���m�=���=Sӽ�T�m������;f�/�`?��E?b�L���S�f�H�>%�?�V�>�>�>��gx�/�>�6?��? \������T�l�X#]=��?낶?�??hpB�r 9��3�f��GO�>T�?���>*�]�5�������`?ci3?nd�>V=	��ǀ�K\��=�>*\?ïF���T>�.�>��>#���S��O��;����"4N�Z�k>vn�<�#�X�_�)� ����=��>/`�> �0��/Ǿ�c�>ݶ��{�r�"���9��X;��i��/$?�Ѿ�3:>re�>��>��jɗ�G�����Y��#?`��?�Q;?�r~?}`Z��+(����HӦ>
wE?/��>kÖ;|�j�k�3>�G?�����l�k(ľ�?db�?���?��T?�T�/Gӿ��,������}��=D%�=�>>��޽ɭ=�K=�Ș��_=�A�>z��>o>C;x>`�T>z�<>^�.>k�����#��ʤ�.ْ��[B�� ����vg��{	��y�����ȴ���k�������xГ���G����?V>��3��-�=���>��?��>:�h>��<*8�qN��V�(R��@���������y���UP�
\��TнY���$�׽��v�>d��r����E>��p�&��:(��>���;�⼣�
�P�=��<b� ���<Μ�=�d>��ȼ��>f>�s�g�z��@����g��>.E?j4>�k"����R������>&�D?���>-;%��؆�i���G�`>�1�fbz�Y�7�e������=H �>��m>��'=-s&�Pƾ�M>��>3{`>�> <½H��eO��ҟ>.��>��Ӿ�iT��E�� �>NJ?��D?��>�'?T2�>c>H����<TOW>&�U>��!?N�S?��?��>u�#=��S��?����PT�g�K��1&�k����B���3��H������K��=S�D>hܞ=r��+ؽft�$�>�P?�0�>KR�>􉤽x����8�E�˾�y�<��l��tn=�;\>��>��>-ޕ>�u�>H!/>�
	�1�޾j��>"v>�}g���i���F���>@�?�?l }?li�>8�����ǻ�ċ>4w>&�>�',?��?�ٙ>���]���iп�{����in�[����c����飯����<����������=)�T>$�p>~�W>�yL>��=dc=�+�>�5>�܆=pن=z�<m[�;֤ ���=aN���;����l��W8;���!	��{�)�n��¥)��a�<�?��>�(>�$��|˾猴�@����>��>ž�>[�y>�Dc>���1Xi��z�l�ǽ�n4?h˂?¸?a�,���_>��=r	�>b�>��->�<>R+��Xu�ǯ>,O�>�Ż>�k�>�X��XG�ZnE�#羓[�>���<�E��xl�?0Y?�����+�?'��G� 
��y2�I���v�.�ž�]��-���	�Q���O�6��=�w�>��?��9�\s�=����L������X_;1Y>�:�=Wp�>%�i>  ͽ���ӓ�O޾�le�m�м��>�
���l;?�q?��	?:�c?4+�>X�>fjR���>�&~>�O-?�/6?ưZ?�0?B�>�����~�<1�<�94D���O�}Ƕ�B�=�t���T >>2?>�/q>��=���Y�>'�T�����n�
�Ӣ��p�,[�=a�>�!�>��>�+?�^�>U۽Ҷ�=��7>d����G>��=�~;��Q�Ňž�޽���>�N>?��S?M}�>m�;��c��O�=$�hm?
M�>,�T?���>֍�=8lV�D�������ǽD�>J8��>�徃����羷꙾B��>��x>����h��%��?�r�?R�f?Ѷe�>�v��F.�9�,�:<`=�5?�=?�>D�*�"�*�������+F��惾��;�&�=�4	>c�>)d>�ͼ�I�=�@�.��^�뼾�">�d>?�?
?!��>
�=�)���0�#F?�r���J�-y1�X�X=b?=�>Z��=�'��-?�2K=��]�Yȗ������$�>,h�?��?�	?�EѾ��@��=5��>2+�=�^$����0A>����&2>0�>�Id�J�"���5�>�Ü>��=�&ϾP��&����:޿��&���T���D�gп��A�����"�=�+<����+��� c�����=�E���M����𾙷ʾ����PGk����?���?��z�>�h-�Z,��R
�0�=b!����d���Z��K7�)�
�I���Y �;�-��.¾������b>Z�K�B7��ՆQ�m�2���� >�3?�೾�3��P��%#�=phW>@M^�Y� ����O��t�����N?��Z?�m��� �1���ȗ=�n?F��>�Z>�vy��jI�˧>4�1?z?q8W������~�
)�<�ʵ?f��?��=?�he�`r@�����˽B��>��?��?��5��˾J-��?9NB?~��>�)˾��q��)���>jfe?��>����>���>~֞>n�Ѽf脾}sڽG����.�i(>\�H���޽>p;�uN�{V�=�܇>sك>k�A������>�h!�k>����<n��t>Q�Y>%R?z�S���X��$�>��>�򾅕���P����-�f�9?j��?(�^?��?Jy$��LھH��a`�>��0?��>���(�_��u=)��>��m�/��.���?)��??��?��L?�H���ܿ)w���௾�8��TN	>O�=�:>�`�K��=��[=���:�s:=L�>>�à>�[>%eH>� 9>��*>�+>�Y����&�if��Q?���7�����A�%�V��k��}^��B���Ә��K����ؽ�枽N���F���!��@��2�Y��Ŭ=�r?iV?{�6>��M>��=����~_�BE.� /̾Y�1�1t�1��!��nQ�{d����k���Ǧ��	�>2�>�5=�J=�f�>#�>������1>}�M�Gr=�dK>��*=č
>YQ7>%�Q>D�>�R>�H�=̀�>�|��Kt�����>��m=�ǆ>�?k�">T!��)�)�>��nѾ�?��X?���>���v����4�֝>�o�����jm�;�>=-y�>W��>]�>�����T~�C��=g��>C�>�{>$N�����c���>p\�>�Ҿ�M�<	v+>Z %?��v?�~D?���=� �>5�0>yM>�l�<��V>�x�>�F�>��?�?�x
?��>f�=�O�ח��v="u�`-3��	ؽ{�u=�C����;@������=8>����܊=,h1<c�ҽlӼ�m=��>���>��>r��>Y�<����^���Ⱦ�RսP���֟=���>�U7>�_�>K�><�>s,>�h"�<y�eT�>��>�=�������޽s�>n�>��1?�tl?��>�7<���_��#�=��;>,��>:�/?��?��>_�"�]#�=ο+4 �OR����=���V����UԽc4�<�4R<����z�=	P>��$>�_>��->
	>VO�=���>�-�>U!>�q�z
�=�"�=YԼz�:��ζ=b,�,�+=�̈́��<����o�ݽR�7�;?�,���%���)=?�?�zv>�|���Խ&�.�U��ӑ<�`?�Q�>�b?D�?Y�>����n�>c��#����>4�u?�?�v���<�M >��>0��>,6��u޺�x>L8�R����[|>���>`
?G{�>��v�$�D�4�S���o!�>��<��=���?�Oj? T��ޗ��&��gL����������%˅��zǾ�F
��`#������nԽ� >I�>+��?A�������3�ؾ�mv�\�u�4�ƾ-`�>��v<LU?�6�>�Nh������+�*0!�%�Ǿ]��) >��ľT�F?��?�>�e�?/?�>���@��>��l>)g?�	?m�^?��?M�>]�˗\�d^��3#v��s8�����L
>���R�g>�C`>5��>�O�=��z��2=~�j��������j���;ŕ�=��>�+(>�n�>�x�>Y �>�u��0�>�$�>��3�=�t�>e<%��ܗ����*����vY>��E?$�W? �?��a�2]�����}<�K#%?kC)?{)J?�ב>�6<=uw(�P-(��g�=כ4=�.�g#���k���m�����>8��>m+&�����?�N?�>?nK���Ⱦ[�z�T=�!/>w!���l2?��?{�>�"���������]�.�-���ܜ��V�=?yR>a
z<z�p>��,��=BQ"�QWｌ��<��=0�=��>"��>̎?I=z>W�p=@�۾�/���;?v��f���%��H����=�3~>]�\>��>�P�>5�X�����:���b
��zI>�g�?��?F*F?t޾�6e�:�[>��q>�T>��*�վܞ?>�=�J>��>oh��uz�U#.���>�x�>(�=��ھ�����O�Ŀ��3��龽��L�d�^�ؾ�����ޕ{���g�
L۾�dl��"I��~R�Rb�U��d�������P��L�?9��?Z�Ľcp�3�[�+���
��;k>cS���qȾ>�޽�K��E���󆽾+����2�5`��+�� �>�Z�L&��'�g�)r\�ж���j�WC2?�ڎ��1q�g��:>�C>���b.��z��Ms��n��\u?�9�?�Z
��7����ʄн`�>��>�C>�8�-}Ͻԕ�>Ն@??������5�x�&.=|ӱ?���?�7>??S_�JC�ؑ�&�νU�?M�?�7�>RF�H)վ����?z�A?��>��Ͼ��s�KX#�� �>_w]?��L��H>$��>�>���5q�������n�nИ�~�(>�}8��Xʽ�!g�>cI��Q�=%�>
d>��\��V��?-u��U�� ���q�&�6C�>#��=�]?�
��봸����>{��>^v�L���=��T4��B?�Э?�s?��?����m����A��.�>[1?а>�E��<F��$^�>s_?df��م�"!���{1?:��?�q�?3�e?w����G׿ǹ���jǾ��ξ���<{m(=�>���4[>_�>�,��
�=�4�>G��>� >��>�8>>�8>uY�=�x��5�'�&a���툿P�L�V�	��K�f�c��\�3uo��g���n���N��v��l��a�*�:�ƪ���ڽ�ʽD�=b1?��?M`�>�b>;�H=�{��n;i�;��������C��.�B1Ⱦ.@��b�>}�
%�K3�������?S�=������>��S=i�>�[>�>�=u'>ez�=��=��C>�"�,��:��=t[p>���f�>�R<(mu�(�b�^o�sc��f��=b^C?��=p����Ig*��dr��u ?��I?�*�>w{�\��2,��[�>p	���J�h��=�t>�̻>O��>���=����(��<�)�;=D�P��>=_�>E��>��s��_����A>���>�ɾg��=)Z>��1?�v�?� 9?\t>�B�>MAQ>��>?�[<%��>7��>�l�>�?�A?�?���>7��=l�d��U�<|�(=�=�^Y�����q�"���ϼGQ��[n�Um�=X��=:�=xp�=�K���aO�2
�;썗=9�?�@?X�>��>���U�l�Y��+�&jU�ytz��=�k�<H\�=j�}>n#�>6��>F�=9��'G �>��>���=i�\��B���8�����=�~�>��f?m�w?:�>�>i���罵�v>.�T>�`>y�>?���>���Y~o>U�ĝſT�4���V��k��(����K<\3B�ve/=�QF>,\����e>7'�>>�`>�%Ѽ8=��ј�v�>x�=���>�@>q��=�A=B�=q8<�L�����<������e�U�=Զ��u|��*�˽W̽�5=m���]#��g;��?��> ��=ez�����Yzƾ9�2��x�>wQ�>��>���>�Q>L&��n��N;��㦼ig6?�L�?��P>s�.���=&�>2y>��>���={�<�_9���Ѿ����� >?��>��>Q�>�r=o�U��b�I8�.:[>��=��G=�d�?��w?�t��&�V��ey:�!�*�:���H���4��?��~?��h,���ߌҾHr̽ �=>5 �?i�;R!}=� ��U�)������)�>�\�<�?��,>aND�kT��`����s�u��yԼ�M>*ʾ���D?�ml?Dx�>� �?�>g?�DϽ���>�� ?8?��?�YF?�&?w�>	�>�~����fK���=k��r��k�	�P�Z��=�?.=L��>IR>!m"�|�=A�x�5��s��3�0��Cϼ�=-t^>şO>q b>2�?�)�>���-��>�b.>�ྲ�@=e�(>����"�!E4�����L>|z(?��c?ƺ?c����^��QI��o#�@�"?�6?΁&?���>��a>ص.�4�-�9��f��q�r(=4㩾�_?�N���Ҿ��C>2�> I����=���?��m??�t?5۝�s꾷ؔ�i2�0�<>E�=��<?���>|��>ͬ)�[�6�嵚�����4��x¾�����H>�6A>��|<�p�>{(�=>dj۽�W�=��<ma�>\͓>}�>G?K�
?�ٽ>�5W=�پ�x�K?�ƾj@�����9馾�Z�=㴤>�;7>�/=d�>]ӽ:T�{^���$��DT>|��?��?��4?^ ��rB�<\`>��8>j">u1E��+��������>���>�<>�l��z^Ǿ�75>��>��>MH�=����[ξٛ׽�ി=�7������o:� ,̾V�P�Ӿ���}�]b � �����v�<�s�����L�j�<���N���;K��o��D��?7Z�?� ���n�>=�P�����"�7�>��c���	��2�/5d��=�Y�پ(1h�D(��U;�ڐ�-ܛ����>�tI�|R����Z���z��e���^>�x�L?�_����ھ���@i�>_!�>��,�e;#�惙��╿;�(�ѓ�?��t?����}4�˯��b�=~]?���>O\>@�t�����,��>\Ug?�?�Ὧq����q�u/l�\ب?+��?��A?X7p� dH�����T"=�e�?��?y�?`\����Lw��\��>T�N?1�?Y� �tT���7���i>��o?;HC�g��=0�>`��>�*j�����,������t� ��=s=4�$8�=Te��81���u<hP�>��J>n��aY����>�Ͼ��H�v�=���c�P��<�	?kf��,p�=
+;> ��=`a5�c���ݞ�����AZH?, �?s�F?�vO? �[��D4��<��>�.�>Y�="�!�@C�>�{�>����7l���ʾs&?β�?��?�H?��W��T޿iv���ﺾ=�����W>�<H>jh>O}2�l:�=�>�| >g\�=��=`g>�@>�Wf>�S>�>�B&�	}�6������6탿��>���� ��O��s��+;r����ɖ�ӧ�2	x������Լ��㽈e������{�mm>L��>	�0>�;�>HG'>]O>L������}s�������'�8�ɾ���"������������0�j�轨4}�՗��,?���=
�MX�>=�����=��>N#�>�=�>&�>��;>K>�y/>Q$p>3�
>�e>�`�Z�>�%}��+��@Y���H��H�R/)>�y??x7w�걄�F�>�l!7�ž�I�>�L!?��>y�ܾb�����?����>��C��I��#�h��8V�]&�>D�>j]L���߻�A���ݾ�?S�|*�>��?�s>Lq|���˾5� md>
�>y�־rz�=�w> �(?��v?�6?*Z�=j�>_-b>�ُ>�'�=�M>�9Q>�Ȉ>��?l�9?O�1?�>�ѿ=c�`��:==�<=f?��2X�����l��M''�T��<�(0��SI=cDv=&�<�+`=�D=55Ǽ�t�;���<��>ܔ�>ɺG>N�"?��A�U�S��C��񅽃� ��$���9�>���>é&?���>L��>G]�>[������jž`�>���>�}���p�v�y��>%�>�c�?-�e?hXI�N��ó��8�N��=���>�~�>���>٭i>�н=��b�ſ�������">dx�<��=���=5�ּxO>D��=~�=fo<F~>��?>��*>�Y>2;>O旽�;�>��n>\��;ɂ>n% ���U�˪!��>�?�<�Z���������qA���?�/<���;X)����ϼ�9?��B?�6��|��ڸ�Xi��t	�;�1>#
?ڞ?�s�>�^>�A��nz�^?w���\���?��l?�p>b�[��>�+&>RQ�=n]">��r<XM!>�I�<�?Z�M��lG>G��>@Q?ԃ�>S��J���hK)����>���=��p��Ȟ?��X?
��˸p�t�2��OL�15 �.4>��(���v�@��� ��k�n0־or�<X"���<���>av?��z��	�>n޾�����G~���o�,=02u=\�?D^�>`D�=A2��O�y{�G�2�&�=�=���=岸>�?�~?��b?�d?��?Y����?|/�=L��>�c�>i?a�
?�S�> �~>�>w� =�y0����Ҋ�Q�<v7���{�=�>\z'>NMa<��"=�5=륿<p�>��������<!�4<2(=(É=��=�>b�?��	?��f��=m�>s�����=�6}=�́�0�\�Dt��Y޼�^a>A?�M/?w�>+0=1����P�{���>�>x�?�Y&?v�C���M�	�������g=��>>�R����N2�}�Ⱦ���=ȳ�>�W=��� 6)>z��?f\�?UO=?��qt�.`��O/�`�T>���>1�?{>���
1�<{�����U�Ggf���<YW�(��]�>R r>t>[y�=�wp>j=��f�-��=�[>�X5�u7�>3��>�?��=��
W̾a��YPA?	Ծ�_!!�}m�L�R�L�>�?��ef>�,b>y?�����q�����
~;��7�>��?���? e7?S���Te	>m1>�;@�ŰK=F^>�ti�	칾|�>>]6�=沘��@��&M=�x>!)5���O��,Խ.����ѽ���ɺ+�o��3����ւ�8=�����
�<=�U�",�wƫ�W,������uP���"��H��~f�P�������a�?�3�?��X=�_���,���ߦ�� �=�䴾u^�8�����g�}ƾ��žk����X׾
���?���ľ_��>4���E�����:���f=Jv�>`�? vӾ�W���B�����|>*[I>�*���)|�糔�ӡ�_�h?��&?�6޾�,߾��\�T��=r�?�F�>�T�=玙�ki7�iH%>\�Q?r�G?�F��`��X��7��=��?���?-??r缾��.���Ⱦ�@���@�>1�^?�c�>�6���)-�c�ҾI�>pX?v0$?�ֳ��b�@�0�X?RS�?a�����>�>ϩ>s��>�Ⱦ�D]=RN�F^����=��|��-8�1�ƾ����$
�=���>�V�>L��^C�R�i>h��q=��f	�����VӾ�v��P?�4��3��y >��<A�����0���jF�&pE?���?%�K?��P?�gξ1����i���=Ec�>o��>�>XG.��#�>π5>�n �>Ga�_W��b�;?�d�?Ъ�? MR?�h�Gӿ��ɶ�������=
%�=`�>>��޽`ȭ=�K=aΘ�0W=���>���>eo>';x>�T>5�<>|�.>Y�����#��ʤ�ْ�2\B�� ����wg��{	��y�{��fȴ��\���-���iϓ���G�4��sT>�~ޭ�7�,>��>PΞ>:��>�~[��}�����,��y�������@%���x�� b�������e��m�w�e0 ���)�)>�<d(/�ڲ�>)$=��:��-�>U����h��c!�>��>��>~�B>��>�F>�y>>�h>�@�=P8(>G	�=fv�>�-�<x���Ί�W��tma�4�>��q?��;�V��r3�O��ƽ���y>��<?;��>:k�����ٞW��=�>�'
��8�����pv��~?I��>��=I@�>��o<�8P���ɽk�=bK�=��+>~ �<�^��#Z��T��=]�?i�����=S(�>G��>�nB?&1?�d�׮�>*ݕ>�\�>��/=�#�>���>�y>'?�?ŽB?D�?�֪=�ý�ʽ�d	>��\��ѩ<�)�=q�>ȹa<pĨ��=�:�G������ݚ�<���=Xą=�U5={*ļ&�b>O��>Yt?p��>6�?�=z5�d�����J�/�н#�>T,>�Y�>^$?��?���>�,>Pn � �辢2�>f~<>Nk��
���`����>�W�>M%�?��v?�/�=rq��#�Z��G��>�{?��?yU,>��A�z�����Blӿ�$���!�%т������;��<���M���E�J�-�.������<M�\>��>��p>��D>��>�@3>�c�>gG>D�=���=�D�;t	;�	F��M=C�ƙE<&VQ�ð�:�Ƽ�̗�f&����I��>�`���4ټ�A?q�)?��������3lC�,	m��y�>�U�>c?�
?5Ӏ>�����q���^��J��Ó?;zh?��>���F�=�/>�p>�0=| �K%(=.5o<QE��㖽~=���>Po?��>��Y��N��胆���M��?Z�=�a��?dO?�a�Ք��4#�	N]��R���>Z�����ҽ�]׽P����Ymɾu��4��ӥ�=�?$�}?���q�)>^Q� p��*�Z��i��L��=��=S?W5> q[=Sh����呾�UL�b�0=�l�>�O��1?�=?��>��h?D�>	��>�剾���>��>2�"?t��>��	?8*�>���>��.>ݷ�=��<��:��KP߽6m����=j�P��%�>6��>3;�>�N>�#!��b=�� =lQ�=b��<$�޼;\=�
5=H��=x�=z�=�v?�p�>�	ǽ���=D�>R�ڽ�4>̾�=�
;�Vܬ������(�A�>x�!?D�#?���>�a>>��l��Rc�\�9���>�� ?��$?��"?d.��KSP����������Ľfc�<����$�J��E�������>�je=�~���_�w?��?��?_����v]��x��D���>-��>�r�>�|�>�tc�X��[�Q�A�j��:h�$P�,��.�оLY�<C�=jN->��
>����?����* �&�)�WP��い=�䃼�9v>&Ƿ>p�>��>o��9L�|��߾-oB?q�$��:;�q�(�*�N��>��0> ��>?�~>���>�A���M���2�)@�>A�?bk�?�{N?��;.�����(>9����8<l�=lc"=R)L>&ゾ���<�e<��E��� �vh5>�h>��ֽ^���l�3�=�c�<��ֿ�4�a���{�������>�62��C�'��߆���v��܋�]���o�S��ّQ�e����m���F���@�LT�?F �?�G>?N>�7S�ӧ3���w��=#���"M��B�⾠`��Ծ���:��ˬ#�s=&��ľ8(����>`̾L���N����_A�(��;\� ?v:N?5�;Y�q�Z�_�Ҵ\>��>�� ���]�a��X#ʼ�sy?��-?��*�җ���'����j=Q�?�
?�K�>�l�����B��=��s?�7`?��3>���/����I��u�?��?]`V?�� �7�g��>����@�>T?H ?��ܾw��r����1?�\�?;c(?�w�:FS�ܰ��!�?�D)?յv�2��>c�>�g�>&�>H���%�o��tʾ���%�W=<>��b��r0�/Ny�
�н�q�>�><ge��d���>b��r�Z�}.I�- �$����M�=B�	?w��c>�=�=��S=r(:�|쌿������ѽy?[�?��&?=\x?z��*���>��GT�a�>�y�>�y��*S�98
>7��>���B b�;e����>�H�?��?��U?ڷ\�;Gӿ��������T��=4%�=�>>��޽�ɭ=��K=�Ř�YY=�n�>v��>	o>3;x>��T>ћ<>��.>m�����#��ʤ�7ْ� \B�� ����vg��{	��y�����ȴ���(�������FГ�h�G�Y���T>�U	���3>&��>��U>3>翕;]�X=l���������%�L6%����'q��Q���bb�𶐾���7\U�ֽ֥ܘ.��:?i��<��}����>�ƾ�.>�a�>D�>ڜ�>��>�z�>��?>{�>>�[6>��"=�q>�O	>ɸ�>�
�J!�������;�`0��j�=��\?ٓ�Rݾ�vE���澈N���f�>�?�or>i#��>��]kL����>�܊���R�u~���_�G��>�� ?"�=� >��U=�Á���G�;�=��n>�U>c>����������l����>�=ľ9�=�E>�,?}�v? 7?��=���>}	p>�¤>I��=�{`>�YH>��w>��?"d7?{Y3?lR�>5��=��3�0h�<F"=��'��H4��P�#�,�������<��R���<=�Xo=~�;6E==���=.�-:]�9;�ZG=��?{�>e><1?����ˋt��������y���x, ���>�?�>v�?e*<?]��>Uù>=��<H�����3=��>+Q>��}�N*����X��1�>7a�>3�?Ob?��ؾ��x>��=�z>�5�>���>���= �]>��<>cp�>տ�RE�fi�mY�=sL�=É�=�E���-=D�E>��:�����:M&->)�>]3�=P��=�d�>'=~ �>�O>�����(>?��=��m=;������=��>�e����;8�����6=�ۃ=T�5�^'�w�=�&H>��?p(?@�%=[��S������r������>��>p�>ɕ�>j;�������q�g�C����{�	?��<?N��>k����6>�0%>p�T>��O>T�>�`7������*�ģ��C/N�k�>ʗ ?y�=�����X{��'��eH�([�>�6>�ž#L�?��N?_� �������^��H]�P��S�#>���"���D=<��xj��楾9���佱z7>T4
?iRC?�߾�W�>��Ѿ,���z�]�U��g90��ᐽ�H�>���>�>mR<M�┾�bk�skG>�X�>��ѾP�>_�&?��>{��?�.A?�9?4է=��$?VI�>�)?��2?���>8>�[�=������=S>-�־�s�:_��]�F�� �N�=� >;�%>b�>7�=�7�<��<�K��2e�<��"�YE�Cc2=�O=>O��>8>e�?�H�>(H��0>�=`��ZI˾m�/��7���\��7��p5ݾ�*���5>�L'?׸6?a
?	3>y>��"�R���&���>d`/?s(1?��F?�O����yǾ��ѾqB���=�>���#ܾ�L���ݾSSͽ6)�>@��$��_�=���?��?��G?��¾�\��5�Kt���+�=Ʊ�>�U?�?�J'��d?�n+��D5���a��k����۽�Ǿ4E��y�=>��=+>zV(=���=N\�����;�=r�>>��m>!�>�\�>���>>E6>jUʽ}(X�t�)��Oj?����
C�D�2�_�˾|e�>YL~>K��>�ȗ=1[>�kH�JT����������RT*?�D�?'�?'K/?�w��F�!�3rv>E��>8Uw>]�M�%z��.�3��ㄾZ,�6�;�PӾۀ���f=�=��9> Zt��(�����A=�#��S�F�KV��ǾQiG���ھ
ߗ�ƭ�yG�pBN=x���aSQ�V������R���֗�\/x�G��fC���?]#�?��>�<н��F��R�܀پ��>@�O/(��g���d��vȾR����
��UȾAS�����@����Ư>���?�����r��<(��5j���>q5?�@¾K�����˴�=c@f>;��=�oʾÀ��^��c�׽��c?K6?�i�Q���"��W�=�\?�G?�^>S�#��k"��`>��(?�g+?���~����J��kd@��)�?ߒ�?�sP?�پXS��ԾH����>.�?y<�>|t��0�>'�����>��X?%V%?ܬ�+4%��F�K?�+j?��Y��ѫ>��@>"
>���=�$<b�=��ߗI=���>�>�=�=��Y�I�[�&�6>���>���>�����1�g��>P�㾲2N�5�C��q���(�d�3<�?�F�6>ě_>E&>^�(��ӌ�����Jj��QL?@�?ıT?�:?Ȭ����m��b$�=�o�>��>��=e1�J�>�w�>y�澼�p�f��B�?7?�?C��?ЦY?�l���ѿ�3���aݾ��ھ�/^>���=m,<>�cb�)��=��o>��+>,� =I� >ϓ}>��a>*7E>e�>f$T>���=BY�����@��Z/���D����"r��é��!پt��8^�c���ξ�0����/g��V�����Oﯽc�>��R�>Z�$?�15>@�'>u�=H��q��	�Y���x��(�&��L�w|���ǻ���b��g-�����8>�y����v�!?c�/9=����U�>��b�Ȑ.=�w�>��>���>뚤>LX>9"">J.�>8�?>�߅=Lu>o�����>]�=��g	dH�[f6=�d�>�'�??�k>x��I\�zl��[����Ð>w�T?EL�>�Q.�����_!��Ұ>�p���s�����P[���F�>��>�>C�>��8�Z�/���I��� >�F>��$>��X=60ܾ�e½�F=L��>��Ծ޳�=F�t>u�(?�x?�6?\ �=b^�>��c>tk�>�v�=X�G>��M>\z�>5�?�:?^D1?=��>���=��^��=�>=\�<��P��q�����8�6��N�<~&�eV=�Zt=�H�;�gH=�0,=�B��y�<�q�<8H?�~�>�y�>,QA?[�(�J�P���4��g�<jF$��+�� ��>�Ϩ>�?J�?!N�>��#>�>��j��� ��P�>>�!>�d��Ԅ~��O;ϐ�>�/?iф?k�(?Ⱦ�YžX\���	�<�4�>��G?��?��>��>C�>Ԥ�������X�!g龆��>!+>==���w�=��>]�j>F�[>����h��u��=C�=&�����F>0��V��>cg2>���c��=��3=����o���$>�S�n�;���Խ�-�<�Ϣ<��f����t�!��<��C=���<@?a�9?���=��{��*@���L�������>i۬>`��>ġ?�[>��%�{���a��B����?1�i?FM�>�<4A>�d?>�$>��>�7;��ӽr�ĩ�n|d�X���>��?��e>�_���惿K����1��r�>T�=��!�]7�?��N?v�:���3R��L�Vn��L>
}N�����/�D �{)��?���[	�<~!�ø?��]?<�%�Y�>�MҾ[핿�s�M+پm�>��>x2?mD�>��8>\������u�6|=z�;(OH= в>Ե?,x?$�d?�(?�]?LM���?4+�=�,�>�{�><?T	?�F�>y9|>o�|>�) =`�7�PY����Q7:<Gث��[�=j�>)%>���<�)=�;,=�W�<O�4�ʩ輗5�<�V�;�=�}�=��=�>�"?A�?��j4u��7��!���
+> "i>�Z�>�;����#I��h�/�\�>��1?7.0?3K�=ע׾u^� ��<��>��?ԩ?��?N�[>r�����|��X8�>�T�>7����m���a۾#I�����=�T?�%>=倽L{f>͘?��{?�H?~K���U‿T*��;�<~�z>���>�>�����=�_ہ�4����8��%`��0��KID����;�\�>��B>�Z�=�`�;Rl>]޹<w#�z+�=�G=����;Y�>c��>�;�>G��=s��쥿��ȗ��RH?ha��L�]�ʾ�Y����>�k�>G�=>�Ì=�O�>Q�;$�m�O���4�9��>�i�?���?D�B?��}�>ٽX�#>ALp>�E�=T�=ߺL��=jj�:E�
����;*">��T�<�}�=��8=����;��"�Khֽ��]�韵��]:���U�X蘾&U�P�׾𐻾����Z�;�7vȾ��0��Es��Z��[�/�Z�����>Z��#�u��\�?6^�?&�=^�
>@`G�h�B�Xm���-<�)�����tbپhm������N�J�����Z&��L(��Y¾��>隈�Q����{��A�����>�YB?(qӾ6��"6���N=�i�>�@ >�夾F��㒐�D&�W`?��+?2���g�ܮ� +1>)�>w�>Z�=q���z@�Μ�>f8N?��H?�U�<����nȕ����Ը?���?�rA?F����!��)���1S����=��?�v�>��u�+�/
���?��o?B�%?����	}��g��P?�i?Oԑ��p�>;��>���>�8�>Ԅ�գL�e�ξ_�a���=�������ص�L�I�+dt�5)�>88�>����(�w{�>�7��j���<�3��Y���Z�8�?8B�:�>+�>&�=��5�kZ��+ҕ��鞾��f?���?�e7?$�^?) ��(��뗾"%V���??���<��Q��}�>���>��?�X����� ?.��?7a@d�_?�lU���ѿ;���,ǎ�h���>���<" >��I�м�=em�=zu�=��9=��=-Q>�H>��e>�ug>!>>@d��Ļ!�n���ȁ��8�\���
���j��{G�5����vh��='����Qq��oy ��X��!`�� a��.�>ַ+?U%�>LV�>zӆ= �=qM���'��b�����Pi.�j���㾷]��(�Z�;��C�-���x���"��.??���=�9�y�?yn���B���4�>L>�_^>���>���>W��>1)>��>���=�	>�/�;���>?=�u�������?E�`Q�x�=��D?(���)㗾mlK�+���(���nj�>w!?�>x� ����g3N����>�EJ���?��[[���b��>o�>�y1>�u=�q�<s�F�o˜�pL=ח=�(�=��=�Ў���	���<���>f]Ӿ��=tJm>��&?1v?�6?��=���> �X>��>��=��J>G�Z>�̏>l�?�5?�50?ܷ�>tƸ=t_��f =L#>=>�?�^�������S��c��羘<�"��
b=��A=):�/b=� \=�6ɼ '<1/�</? �F>8P�>�#'?�l�@B�Y;c��߾����H ���+?��f?S�j?��+?)�r>�S��z��ƥ�<rT<���>2;>��g��j�E鐽,=�>3>?��p?�?�.������:>.1�==�>���>z@�>���>ɱ�>帚���I��e���L$Ǿ_��>c��������W���p<$��=8�\>R�=�[һpV����t��˼�">�ؽ.ս=>�>cr>>?�<Ǹ=�{�=Y�W<�Pn>^h��Mҽ_����<Ѯ$�-7μ�λ%黵������(&�<�?n7?�C=t����j�D�߾�ދ���?���>|�?(}?!�T��T�[�p�+�=�V[����>	>I?��>�����>�>�=E�=�>���>�.1�����||�zX�|� ���>z?�Ma>\���L�l����S%���x>DO�=.hw���?M�d?�'�{뇾*?�!ds����[�>8�⽄��E���V�־����F��Q��z*Q�6S���	?6?35ɾ �>�3ξQ݌��ȋ��vﾠ�>")3>�Y5?A�?M�>�Ҽ�
��p�վ�L	�*�J>�҈�>n�=�U�>G?	a?%$f?e?L�?�y�L�?�^�=��>GG�>7?��?��>I�r>h�u>2�[=�Ǽ��	��������;azƼLB�=P�>�->��=��=��<}=���H$�}<=k�<
Vv<��V=G�=��>��?P�>�U��5&)�1�]��<���dS>h">@�G>es%=e0��rq���:=T�>�VJ?ۃ9?��<b�S�5ѽ�rg����>. 6?NV?��9?��*�"���9�N���g�=�J�>������|�$�����7>J��>\�>��`>.��?Cj?.AU?\��=Լ�֓{�·��>ƣ�;a�Z>g6>K�$�L�6��g���D��5���y���'���l��p=���>�7>�@>}y�=�C�=�jV�~�V�^��N�:�>�=�>Ҥ>SH�>F=�����(ھD+���mG?ܗE���B��Ծj��eƔ�Jl�>�C�>�<	��9%?:}�Lƀ��Þ��u*��	?�i�?���?�u+?��#����O�=�9|>���=>�s�i����_N�~��eDC=���=�&��	����L>���>jH�>�����Ծ�'�������D$�N_;�I�t�a2��Ȕ����⾪Žno��=z6�5V����!���aˆ�I�J�zr��������X�V�?���?�V(��a=�:��ZA�{m���>U����<YS��Hjc�Q�����Q�̾��$�W���߾�gn�>z�"�����3b������!�>#�,?�ξj����
��Ƙ=�G�=�ົ����ϣ���O������P?�"N?Сݾ�>��J��5m<�?�>��v>������*�>�E'?�0#?�p��4Ȏ��q���i?=���?(߲?��=?1:��aA�3�C��*'��̆?��X? `?�?�=��a�eξČ�>��H?<�E?�^ ��]s���)�6�?iS?G �s�>n3->���'�S�J�Z�z�<ߩ��LD�>�؁>�����W���<�bYl>V�?�t>ܲ�������>�����>��,G�E ��=�9��<y��>6� ���6>y�I>�6�=d-�����'�)4�L�:?ረ?1WV?I#?j������*ս�0t=�o�>��>(5�=\y�|�>�b�>����]a���'�?Me�?���?,�J?E�u�>Gӿ��!������
��=%�=��>>��޽�ɭ=��K=�ɘ�0Z=�n�>���>o>D;x>w�T>ϛ<>��.>r�����#��ʤ�4ْ��[B�� ���wg��{	��y�����ȴ���K�������<Г�y�G�^���T>�з��u��M�
?)O�=Ș?u�1>��p=��վ;�����=�����_��6���"�!���Ã��ٌ��v��V���3���1�ܪ?f�����R>�1?)���ћ1>��>��;>�t>�ڜ��5�=���>�?�;?��>�eI>^�e�;%>�'>�(��߻e��͇��\ɾו>� }?f��=�F��L��-�ھ{����>	0�>A���J�F��e^Y��O?�A=c$���h=�4��c�=:��>�@<=�h>����W�(>�Pq<8��>�˞<�=5��@��g������<�G�>�C����=Q�}>7�0?�Bz?V�$?�7+=�'�>m�><�>��<���>��B>�7�>)�#?A�P?f~;?5��>=#�"�x�{$��|H=.�ɽm=Fτ�z"���Plq��_����>�<>�<d<�"�) >���<��1�=%?�>�3?���> @�>��H��&�޺8���нUQT>rUd=A� ?һ?�?�a	?\�?_��>X>$>m6����
���>��!><�_���k� �;llA>k�z>��a?o�7?�CS��vv�\��/��щ>�I�>�?���>���>!��<����G࿚��.�%����;�͢=��x�z�Y���p><��=׽(p��0�[<�ϐ>�>;�>X��>�mp>Kpp>�x�>o�1>�E�=~��=J�<]���t-����=V����;�\%����=�)>�i���,��_��Q���d���K��~?�H?�!&�sz���uf�=���۪�Ok�>��>(=�>�R�>��=�q���U�7�A��G���>�hh?��>/�:�f!�=��)���:��>��>��>e���������<x��>k�?��>�����Z��Co�	�
����>��=�]L�c�?�&?�7�X"=01P�\�a�G	���L>���=���uό=��K��� ��H��8��R� ̈�e��>��? 磾�?6�ʾ�����������d�w�ט;�b=�>Q�>�|����IM���5�����R���>?p�>�́>�d�>)�?�8?��;?>�>�*�-�?�&�>n�?��E>4�?��>TO?Q�	?�&?N�l>��k=p{F�S���Q������I<��+>��|>�H��*�~=JXp�硠�z�`=9?<�	h�&��t�<���;��=t��>h� ?�#$?�=�"x>��=�H_�G���>=:w�=��<P҉�F�c=C�>A�?�NF?��>�a>�{���5�w�
�7B�� ?F�+?�8�>�<w>�a>�Qܾ\͈��|>�0`>�3b���!�R@~������z�>�g>�!^>��>��?ߺ1?�eB?pv���d�������?�Q�P��˺�e��>c��>
f�=�վh$�`�?���E�V>:�����ڋ��[Z��y�=tWT>hװ>u.��ɋ�=f�@>Ǚ= ޼�Et���>�NG>���>+<H?���>�1�>H�ξ7k@��C?;ܽ�;������������'����=g3>���A`?A����}�����_>���>f��?�B�?.�_?�Q��P��EYR>��u>�>h����!��V���+��(�5>	�=@�3��p�#��=�A>��>����@�Ⱦk�ľ5 ����ſ��V��&�?0�4�i�	1���͜�k}�=x�x����c���ִg���5��I���D)�ѳ��2����Ů?��?`�b���/��`�ox+����U�>A���E���$�y��L�Ӿ$S[�K2ƾ��8�o���g�8����6�>�[޽"w���惿��&�	g����
?>�v?҂о<� �+�h��ڶ>a��̂c>����by���p��]���eR?��"?�����C��plH����>���>1�>��=+���#+=��?�/?���>�W��A����j��x�t��?���?ӲD?��C�ΡJ����Ty���w>��.?*��>�&Ӿ1��_�U�a�O?1��>0&P=F�Y��"����>�<�?c�?7H��w�=>�DQ?��> �߽���㐽����־s�]b?��=�ɣ����AG�t��Z�>�7>�����!����>^3��N���H���l�����<�Q?'��\>d9h>�	>�`(�f ��Bى�˵�~�L?���?}S?�7?�F���k񦽷��=�w�>tm�>��=���	��>�9�>g��Vkr����0�?�'�?���?�Z?�~m�9Eӿ.	��%���������=UN�=��>>I�޽"��=��K=J����>���>A��>=�n>�+x>��T>�<> />c���
�#�fȤ��֒�dUB����М�5dg�}v	��y�e���ȴ��Wx�����}����vG�Ñ�wG>�KھB��uӨ>���=/��>%��>��d>��-��.�G�^�;�������v��?���[=�%���e�`)��{@'�w�?���%5m>�F?�V<v�> �~>�RǼ {�>�@��FJػ� f>���>��>.�>T��=�V�<�N>: N>�䛿�����3��辌�r>�b\?�m�p�9��s��0�ف����>7�>���h0���\N��0�(?��Ƚ׌�pAk�*w<mWZ>��?#=nN���9�Rķ�:>	�=���>[?N����=�ʾ�=��>�͠>���2>��7>Ƶa?43�?C�3?7�:J��>��>]W�>���H2�>V*�>2Ȭ>�1?�K?��8?�?�k�=�v�'+�=���<�����;�F������L�W�Zfz�ۓX����� =>���+=�֌�:�J�l=�<���;:��>��??���>	�?]�_�;+�msT��E8��Ȣ>ML���?���>��>�f�>k��>V��>/xB>A����|���>�|>=^g��,|���4��A@=EN>em?�7^?r���H�=Fi���e���`>|��>�WL?�U?���>�-�ָ��0ӿ'�#��!�zc~�K� ��
�;*;��/R��c:�^.��)����<�f]>�'�>�xp>a�D>�?>�A4>�r�>D�B>
��=��=�3�;�`;�D�.sN=�m�K�f<e6Q�o���)���j�����6>���;�@V�	ݼ>�?~�?��<ïŻ��_��M���8#�Q�>9{?��>�V?�#}=��$���Y�z!����7?.i�?�=�>��m�q��9)<���=�Z�>I�>;V�>m�%�7�������*5�Ti�>(?��>']=�hWp�	q�1E�����>�Ȝ=�������?z�b?�u���Ƚ_���l����>j4S�ݞO�R� ��k�"�A�rɾ\q�������>���>���?T�t�l#	?.Jھ�r���*�����b=~u�>�A?�+m>9: =϶辸�]�t ޾�D���{���>wg�=x`�>�%?e�?*�?)L2?Q�>�赾��>M>5>�?2�x>��)?Z�>
@�>�G�>*�><e�<���X�>�;p�z�Ļq��<�#�=<f@>9��<��;o���F=�#���L>���=�R��2�`;jC>���=�Q5>Q�?]j?���<�~�=�x�=�VC��(��������=�
ռҭ<���>U<>���>k�I?s�>n�=��߾x�"�)��l:��%'?�"?KQ�>�K�>Q��>�N��؎�k|?>�0�<>P��c�%қ�X]t�z9��G�>-<�>�>���>�x�?��;?[�R?���NZW�G���-���彸�k=D��>?�?���=����/��<�K�H��L�����1P�!�=�?��A�-�>
��<ݷ�;�W/>va=�ž~>#�L>ē	> n?��8?��>��F><վ�08���A?k�H��h��Ɛ����g�Ʌ�=6�>���=��?:u;�{�#Ȩ���<�Y	�>���?~��?e,q?W�&�^����=>b�4>c�d=4$=1�	�S�=ϴ�;?�/>y��=�a��������Z����=:C@>�ɽjџ��^�����9ѧۿ��_���e��¾a��`��������=(��n���Kؾ�⽾��s�BZ>���]=�\���<��m��92��A��?���?�O�⢼��_�I>��&�mZ>b�H�����&��*���+�_���.���C�UcD� /\�
DW���>�?��Ԗ��K���.�j{C�/�>�U8?f��y�־I�+��Ǜ=Ӓ=�l�= ���{��C���z��Q�R?�*?���A۾��_ϭ=ֻ?�e�>�>���']��	�>8:?B+?�}R�����������꼖B�?V�?#BR?=�%���Q��)��Ѿv>�.?���>�7��:���Y־��0?f�&?6��>�>��ކ���K�
�>M}^?8*Ⱦ�٘=[�*?%Ů>���Q�;�>�Ⱦf�����T??�#4>�*Q<W��=�p��c��<�>+�>�߽􂀾���>����l�1�Y����`��_�>|��>�9��M����>���>�O<�U���렿	@��m�M?���?N�7?��+?;����Ez�r)�n�>|��>'�y=�㻽����
��>���>����|]������>���?
�?��H?��F��jܿA�������8 ؾ�>#��=e�>�y�\C�=v&�=|�q��;����N>��>;pv>+w>2�>�|>} >����;p%�����	���#w+���	���-�R4��s��e�ڏ\�����2�Y�K}^���?�T���y���^�:�f��J>�(�>���>#�>8W�>�>Y�����g�fT��F������@��OD¾�/��=��s�8�(o��̴�Q���x�>F��=�V>�	?�~���">i��>9�:e�>q��>�8�>c~>�ܑ>�?�>��)>y�=��=�>RDh>Z�����=e�$�¾��k>> �?�m���1�G@�����Ԡ�rw.>!�>�<�BÇ�%I���]�h$�>w��=ge�D4�=�@�0�=k��>;���=�VT=��ݽ�&�TԺR^,>��E>r1@�Uo�d:�<Ŋ���>������="�D<��*?ҡ�?��?��N=,V>,�">�x>U>'��>_��>=r>��?�??o+?b?ũ >{e���>	r��B���G����a�2s�<�m^>��>����C;��@=�z>�~�=u�(=j��<� )>S����?�u7?�x?Gt�>K,i�����7����^?�
s�8 �>��ؽj؝>]�?�O'?F�r>QZ����<��Mw�< �>i�>�cE�X�t�D������:V{>�rq?3&`?�O��D�9��ﯽ�1�<.Tk>��>�O?7��>�#�>��p=�-���ݿ)�d�0�о?,����F�)aȽ�,����ü�:>J����o��g,�>�l�>�{_>��?AYI>��w>���>���>��>�8�<���=��^<�����ϔ=	c>����(���ֽ�8ǻ����S5��6��
Z;� ��u
�*f�=?�?-?���=�߁��o������}{2>BV��w��>�Da>��>rN;�Ap���w��j��1?��?�P�>E����:b�@>ʄ��O��>)�$?7�<~ͅ�����LT�����mǎ>�oL?z�!?!hn=2>���\�~���C�>u>ho���?�%6?5�2�
��H�MG[���p�pP�>+������]�����S�A�R��+������m=/��>��>��?�0����>H��Ф�>�~�C��w��=�ֹ>z4*?)��=B���[
�t�>�����"��|y���Ӵ>cq>�_>��>�?u��?��z?�
?�T�j?\�5>�>�����A?�h.?�T?�?h��>6i<�$����`����C�JR��"�:�;�y>Y��=H�=�m2�O��[����`+�,䗻���<���;.ߗ<B!>m�I>4?v;?��	���F�*;���'��=�8�>�� ?�L�=��ߋC���=�3?x�??���>��]>OO��(ݾ7V��^ҽ��>rJV?�?eP|>���=�O+��Ӿ��>Vn>��&>�%��Š��Z������F>�>�S>�1�>��?�p?wg?5�����B�O���|:�D�佘��>Z�z?Ǔ?6�b�h7��Z��=���|}���E����=�t�%G��7F��6�n=`!�>�`7>4s>}}>אݽ�(����8�X$��g�>��!?F�E?�>p�->�?�1�>��FK?m*���d��ѡ��MѾ\��i)>�:>_�'��+�>ʙ�$^s��;��APF�$��>���?���?og?��>���	�v�Z>�ņ>t>l��;O�I�������M&>9�>jv��͇����,|F>Y(o>�����ƾ�OྮTL�2J����N�7|���Y �>�n� 0���~��a�>鏾�Α�O��@'��S��T�A���p�	�nq���4��mi��?xN�?l-_=�֠�G�e���#�����>y�ϾMc޾���+-�6 ���gھ���M���v�-�?�*���>N�ý�G���P��#G�)\����>��:?���q�#����?s>DT}�Q��g�M(��-���{3��t;?�@?�kӾD��g�5����>�r�>86?v�4>E~���Q��r	?��T?5"#?��Y�|���kt��+�>7�?}O�?{D?����F�|��b���^�>��?��>:X����쾴;��?�?��?W�8>�W �_�}���?�
K?$�;�Z[Z>U?�)�>Փ!�Y���O��(�Q�;��>��K�ߵ#��$��c�k�ja�=؃�>���>l�S�B䪾��>:Dܾ�B�0�7����I�c�7��=_B�>�	���>>b�Q>�H>p�#�Bc���w��j�!�w=?쿬?�qW?��(?o�뾾?��� _��Y�=S��>�b>�_=b���Ԣ�>O��>�#��"�p����4�?f��?һ�?!�I?`�j��o���𔿅��Zu�.T�<C�M>��e>82ӽ\��=�[�=������<��>1y�>��m>��>���>Ї`>Ҟ�=u��Q�m��ꏒ� �V�L�	��Ծbi��d龲�.�Hk��;ﾱ���=.�A�O�/��(��^��O�;�Ds����=�� ?�f�>�+�>Ũ�>F*)>MF����*�&�t��%��C'��1ܾ����^�o��L���Ms7������"Y���8�4��>�Y�G/(�b/<?�#=�]�>�̪>�O��=�ɽ���>9?��>�<_>�l>�P>��>�Zb���h>sk>�ӈ�4�~���]�/Ԛ��Ӹ=�6N?�=���˾��G��ӽ�z���~�8>��>,��=!,;��3��7Hl���>�4�;��b�L=�V��h4�=� �>N�U=��$=y�<9�^��� =���=X�>^�o<&��ANq�{/=�E�>9���l>�Q0>��"?SZ�?�_?'Xc>h:�>uf�=��>�%a=��>��">�\�>��?,?-ZH?��>���=%,��\�>E�<>$���9�i9�N���:�}Ao<�[a=��~����=�À=�\����1>���=�諽hC>���<�k??�H?||�>���>���<&�JEL�{ ��p�>T	G=��?�#�>�ע>*�?Z?Q�>���=��c}*����>��'>\\�І}�U����E�=�v�=�w?��P?�������t��;���X,Q>,R?�m>?��$?6��>Cj��*��9���%�-�j�O� ��<͇>o��=�I�=�=�[�>
il����&#��f�%?Jv�>/��>�?���>��>ws�>�2>RO�=���<�>o�ȣ��Ͷ<Z�=�bm��b��8ģ=�]��G���KƦ�a�ܽQ,���={�=��?�?��=�p\�v��(���Da��>�s>f�>қ&?	^�>��r<.���l�g?���W����>��V?}?)2�����=m�W���K���?7?r��<J*��i���2���E>�)�=9��>��>��4<m�:�8�b��r ����>�M>i�^�6��?+�?6�}�4�ԡ���l��q��ͦ�=$���r`ɽ,�@�Y�9�+*.��"��J_���Q��6>�G�>�λ?G�߽�^�>Z=����u��Q����=�`�>1�%?{W>c���w��cOX�S2Ǿ�^�b/оhAM>ۜ>���>V�%?j?]�k?H�?���>�����?�>'�?�{�>-�
?��?.r?a�>^��>�S	=#&�X��	��Ub<1=���=C>�OP>���F�}=5�N=�k�:��O�Y�6�e��=PI�<��<�pA=(�E>UPC>��?1�8?~}�)��=+�>>�)�~.:��k$>�>�>��`� P�<�r����>-��>��K?j?��$>]��w$E�Ɖپ�$���?9�?�i�>}
#>���>�JǾ�����N>�a�>6 	��½"u���]�ĭ��̡>�$�>h�6>3�>F݇?,(G?�:8?�KI��1��C��3=�F�>a��=�
?�P�>p���[$���4��&�-�B��pl��=�o���3��=?<��������>�g�=��; S>�kD��[��3����<�Z��>�?s~C?�>Vΰ<�_̾�K7���I?�z��À�[⠾�j˾�E���>G>�=��?g��0}�>V��Ǹ;�~�>���?�*�?�|c?��J�~����[>s�U>{�>��J<vR<�8�ּe���,>���=_u�����m�<
�S>��x>z�ͽ�ƾi6߾Rq��੿�'7��Ԃ�h��B�x�����t�|��O�=:����n�e�Z��ѭ��t����Ϥ7�U�f���J��H��w�?-��?ֽѽ(o�/Qa��
-�9sQ���l>�뤾}���^� ��@��M��Z0#�3&־~�=�]|��_F�A�S&�>"����ꍿ��e��&�1F�����>?�j?͓þ�
���R����>r��=a�,��˓��|����G�<��:?=C?�������u�M�e��>.�?�?�	.>�`��� ~���b<�C?)?z��=kd��gR������9Z�?�z�?I�S?�~�� [���U���m�=� ]?��>�\��| �$ƾ��G?@R	?J*�;rE[�����2L�c;?�ă?�(�|l>݈:?so�>F���o���v��`b�{��<��>�qc>�S��%��ʾq�+�?-Y�>BZi��������>�=��N���H�����\u�<6~?}��C>�h>�Q>��(����щ��H�^�L?{��?��S?�d8?Zc��T��敧�eƐ=y��>��>���=������>���>�d��mr�G�@�?vI�?*��?TRZ?b�m��7߿Ju���߾����i)>�&>��>�LM�T[>��<I�t���x,�=Q.�>��>��>�Mt>�'�>�L>�A��ͨ!�#���� ��t� �iG�m0��S��w!���������˾ȣ �( �9�$B(�Q�a-;<�^���zн_zt?��@=��>�F@>7rD> c����U�u�=)-ɾ������������F>\�Pc���[ֽ�t��O|6�KV�>��=�O�>u%H?�,��Aej>?%�>S�>N�>*��=��>-�>�p�>��>���>�ͽ�t�=�$�>	�w�����׋l�qn)��'����?�/(��Q�x�R����c.�F��>\�P>�~��|������E�&a�>��G=+E������X����->�L�>{*/>�{�iv-�*BҾ�.R�Jh�=��>ī=�w >���2G�0琾Q-�>Q����A<[F�>��@?m�x?'�:?[��:���>��X>~)�>&����>��>!;�>b�+?��8?��/?Y?��=~>:����=��=>gT�-e,<=@u��.��.f��n������vV�&>��=��=0�<\cl�T�Z<[�l=��?5�f?u%>��>�%��2���^�
*|�N���S�=.�(?��3?+��>�3�=��>b�N>��=�8߾:�4����>�*�>��s�
@{�W�=x	��T�=	�d?<�I?�����շ��ϼõ>�C�>�h-?B0?d�?LQ��< A�*��&vտ��6�=�'�^�+���H=�(7��)1�v>�Ng=$-�b(ξK�f>��>}��>Q��>�i�>�5�>���>���>`\2>_��<c�=
<�뻥bJ=܆�=QeR<��I�QO�2%9��{W�H��y�=8��<�.���/u=�J�=��?�3?�����K<̦[����`����!?n��>`�?��?ܟ�=u񾕊A���˾����I/?Y�{?H?�i(��Ň:�5伓��=��>�Ү>�B�>e��(:��n�Q��;��>v3)?�?�>yi��GS�(���g:�`�	?�_o>&�\w�?GeQ??�A��iO��iM��'M�b������>
�����<�=2�'���@r}���sY�N#�D��>?K�>>E�?S޾�;F>A���R���]s�f��lY0�)�7=�%?މ;>��J�����'�*�Ǿ�ʮ�9��HM�>��Q>D�=C5�>��d?pن?��r?f�9?-3�2��>{p
>Š?�/�{�G?2�2?�? �?��>��j>\w�=񛡽��q�SF������y�=!}>�9>[�=�J>�����;�V�=�C�8����W#��C�=I
�=,m�=��'��?��;?E�[�e[>�h�<�����F�ڻ�$彄K�<h/�=g�>
��>�/�>̲/?Il�>'�+>6�$��V��w�I'���)? BO?{�>T��>q��>����z߾�c�>P��>xUy�	2��K�S@�\����>��?�^�==y>��d?MXV?د�>��a�GH�%�X���9� ���{Φ=w�=Hn�>b0=<q�U?X��-x��Dc��B�hB=U6v�����>_S�=�i�>tuo>F�>D�6�1�-�,�=���=&<�_�>	[�>�<?���>�ϸ=�\ھT���I?JK���>�����7о�Qk��1�=f�m>z�ѽ��?�����v�r��f�>�Tg�>���?�?�l?"�]����S>��G>� >�'���=���P��<��i>���=H�������(�^uC>�}s>���R0����Ǿ��=�G��~!J�D����ؾ�,���i˾H���4�Q=A�����h�����|���LQ���.��mɾx�¾���yHʽ�1�?�R�?�.>~b�N�Z�=�J�-
�A��>P7�P�������e�>��\��er�5R{�Z���B�-��a��g�>~�|��|��뉿�VE���=����>��N?ƥd�a� �{�U�O\>Mҕ���=]V�Yܘ��,����e��,)?�h'?�\龎������u >A��>v��>��H���Ծ��,>��>h\?�>�)����V⊿�=�?��?�;?�-��k/��?��=O��_�>��?a�>0O��A�ྩ�[��.?u ? �>G�?a��C�%�	��>t!Z?w�N�͔8>?�>�ƽ�˭�+�/���;I��R[�>����C꽻4!�PϢ����;7�> n�>?���P�>���F�%o?�� 
�Z�0���<j&?��a�=�׀>� >}#%�Gt��*���
�̽D�Q?Ծ�?.�G?�5?^�󾉃��چ��%u>~A�>*9�>�`=�� ����>c��>t|���fk���NZ�>	��?�U�?-�[?�Fk�˒��<[���Z����/�~=���=�8>��W#b>Pf�=��b>����$�=�4�>O�B>+8s>��~>�>�׀>�E��T��C�ÿn政��C�3�5�P/��!D���پ�1ྥ]������1��}u{=�y�����Ꮎ����0�X��9�`(��m�>r��>p&�>2\�>��!?�%��T�*�|ݤ<������qE�ɡC�@(����R�˾�S�����=�½>�/�-��>��n>?��=��?�ߪ���R�"��>E�>x�>�.>�77>N��=ͱ >k��>̛T>K�5��n�=��<��==Xܑ��)���\����\��S�I?_C���"���꾷���hA���S�����>e�>Hd��w���Î�;�>̿�=��{�3̲�y�`>4��>4<>��>���
����sRY��A�=�Y~>�6�>�Q\���
�G�x�Yc>�3?ֈ�Q��>q��>Qz;?�m_?=��>��ƽI�?�s�>��=�[�4�n>�`�>?��={�?Ar=?F^=?�G?I��=�<����>^�">	<}����m㑼j�=�Իw��=��_�e���V<��=��@>��y�����5/>G->&K?u)?V��>���>����(^���	��)X<3�>��<�3g>i:�=o)?Z��>�]�>>p>�<F���e�ɾS�?�9<>0+���Rz��=��/>OW>�i?S?��Ͼd=��q>��H���>D��>z�$?�9?w�>���R����ҿ�$�5�"�p������X�;��9���G�dҺ�0�G�ｐ�<�V>u>�>�8t>l�I>N�>�+>rS�>�I>��=�v�=��;�R�;��W�E�U=H���)<ڍX�E����ԯ��ࡽ嗊��K�*B�V�������J?�?���<��=�g�;��X���ƾ�^>���>5�>^��>v��>Hf��c�:��D�=z�R?X0b?�+�>,�4�D� >TN(�Ŵ�=(?�z�>�c��s?���P>p|��v|U�H�3>
?
?r��>'���J+1��0K����]�>`jͺ �����?��c?���E�o��"Q��f���qg>�����O�z����4{!��`��Ԧ徳���Ⱦ>M?�?Q�9�el������`��R�n�]G�=�����"�>�..>]_�'H��i�ݾn�Ⱦ�~o��/�=��=�>M~�>}4'?�g2?_b?��?���>_S^��?K�K>J̪>DA�>��?(�*?�w	?�v>.^>�/�=:�<�l�%x�����=傸<5 �<���=�'>��y=@,�=�З=;=[;<�����
p���U=�Q�<�5>I�5>�[:>:i
?(-?���(�=�y�<�wb��� =pi�=w3�>U�U��Á�Y�|��>/?��)?�)�>0�=�m�����b�	��\K=L�&?�)?���>��>?�>���Y��B(>�W>T�ȼ��Ͼ C��;���j0��\�>�6�>��=�;�=s^�?�Z`?@V�>%�!�DR�S���Y$V�2����G>�.>�$?y��>hH�������.���\��!2�$���먽���=J6>��r>k8>,b�=�8>��н�t���>Q6b>�al�	��=���>�>+�=�|��қw�D���kN?�_�����ϕ��Ѿ� G��>��G>���S��>W���`s��-����:� �>ی�?���? 0g?{M�]f��*?S>=>�>�0L=x���8�OP��j�8>	t�=�f�Bv�D��;V�J>�#P>���*V����վ��\��}��y}����
c���پS籾�*)����!t��������{�WN������ܺ�<_�;��=HxU�|ZԾMľ��a?n��?6�=*yԾ�J���ט���C�=-L��9e�Ñ���=�I���Q��������ٽ��A�57�D��><�@�����(��*�Ⱦvx�=��=��_?|�vL׾E�^�]�u�7���5�=uO�撿j�� �D��WI?m�-?���SҾS诼��=%��>���>LA!>JS��U�_=(_�>0�?_B?"f�<�?��2����=nE�?�D�?&�"?>cb��P��y(�r�����>:x"?��,?�[��bϾ�G�=���>��>?��>D7�Y棿������>]�z?��T�:6g>�8?���>fl������^d�>�� T>��^=�B���c��)�<T�����?�>z�>x�
J�����>E�r�N��H����\[�\�<�}?T���z>�Ei>�>�(���D׉�����L?���?��S?�J8?}1���t�YM���ڏ=X�>�>V��=���,Ǟ>���>�a��ir�J
���?�7�?���?�JZ?+�m�cGӿ8��0���������=�$�=T�>>��޽ʭ=:�K=u���8P=�̉>`��>Oo>�;x>W�T>r�<>��.>T���g�#��ʤ�#ْ��[B�� ����tvg��{	��y�����ȴ��񽾉�������ѓ���G�r���U>�6�� U�=�8�>*S+?��?��>��>�g�k�;�vy<��L�!tF�@����N-�����#�������߆��$G�,��~ظ>�]=��->d��>c��<�@1>�x�>)�&�$)���&>MR�9i�ֻr'�>M7�>%A=�4#�,�`�K/M>�m�=��t�l���]2J�@!վ�K>-]6?�˼�{�Xd:�*��%�˾�~>W�?�ܭ>Nh��2��b�����>itu;�����2�P�>!~�>�>�	d=��:����aY=�D�=��>���>�A�� 5ؾ,ڄ����=�t?S��,>��>�Q�>FM�?r?��=.?&ݷ>�����q>�ȭ>Q�>���>�?\�K?�%?T��>�L�=ϒ��_V�����=�+��Ih���Ľ��a/���<x��gQ	�}|㽚v=k}d;�a$�:Dd=�y4=W͘��*�>�}u?ϴ?��d>�ڦ���Y�5�J���B���>�|�=8V[>��?�F?���>��>:�1>�=��־����>�=(�*�춃��ξ��7>^��>��\?�)?]e���U��e:�>v�;>=.�>�|5?+�Q?o�>3��sj9�\`��lƿ�.L��ﾬ½��~���B��/<���0{���>b`ľ�Ծ=�ܽڼJ>Tt�>)�~>+L�>c�=8�?z!_>�2���;>����>���<=0�<�_<�E�i�'���=5��5iX=ޙ���J�=<N�<ܫʽL#��W?�?n}K��2��.m��M;�`��X�>p��>N ?���>ޛ%�kR���<���N�ց���n�>�w?�?}��g��=�6�<��=��>�,}>͂>���� �Y�^%��������>���>d��>.�
�_��y[�>�L4>+*Y< �'�?Qk^?e⳾L�8�W�,��L_��� ����=��)�w������&���1�Vv�rU%��j3���I>E)�>�T�?G;�C�=�;���~��f����.�=�='��>�[�>ƭ�e�?����{����þ��=�܈>�Q��d�>�T?$�>?X`4?B�+?Vq?�ě�ZF$?ߗ#>/��>�{�>m�>�?'\�>�?�?Cս&���'?������(��
n����=� e>�d*>��=gb>�al=��ؽ1D=��F=�Q�_+H�y��=�F�>OT>��p>(�>/D?6!�>u�<�[-�B)��J4��u�=���>�@Y�|1��»�D�7>Ar�>��:?�k?����`%�\�پ��O��ڽf1.?c�6?\ ?>b;>@��=�	���6���=���>��˟��4�M�W^R���H>2�>��7>g[P>C�?P@E?y6?�?��шL������B��"�=T�E>���>;�>=}p>}�W�B���\��e����v�F<�(�*A>��#>k��=�>�Bf��1t=/s�<�5�=M��k"=���=Wr?�v�>�8�>�w>MG�>"N��x}�<n?�������ͫn�^���|�=њ�>��[>]�=
�?�$Ѿ+�R�	�������	�?�}�?wg�?^�0?���F\��NA�>���=��¼a�>9�˾��Ͼ��U�Vo{>��(��Y�=_�����H��Ǹ�q>#!�=���n$����=�y̿�l|���Ǿ��̾�E�]:��;�о�ͺ�
@v�כ�#�
��H���ƾ��G���Z������/�Y�͉����?�'�?:;��U���2��'�7s���f#>�鮾uQ*��1e������3����Ѿ��j��k�e�8�YD6�E����>��ý����vR�����
x���q�>�?��þ�S�}�*��+�>#�&>�<��ŹAm�����ˈ���? �.?R)�i/���<>��>��O?�Ѱ>�E��c��v��>:I�>*��>��?�4
>b�������*@>��?�2�?��<?|@��|�b��h�-�=�Y=?qv>'�>E������&>���>� A?���3"V�񎊿������V?�?q��ە >.?D�>�Ϻ��h��=������ns>}�Ѽ*���������=�|�>��>��<U'+�P�>���F�%o?�� 
�Z�0���<j&?��a�=�׀>� >}#%�Gt��*���
�̽D�Q?Ծ�?.�G?�5?^�󾉃��چ��%u>~A�>*9�>�`=�� ����>c��>t|���fk���NZ�>	��?�U�?-�[?�Fk�˒��<[���Z����/�~=���=�8>��W#b>Pf�=��b>����$�=�4�>O�B>+8s>��~>�>�׀>�E��T��C�ÿn政��C�3�5�P/��!D���پ�1ྥ]������1��}u{=�y�����Ꮎ����0�X��9�`(��m�>r��>p&�>2\�>��!?�%��T�*�|ݤ<������qE�ɡC�@(����R�˾�S�����=�½>�/�-��>��n>?��=��?�ߪ���R�"��>E�>x�>�.>�77>N��=ͱ >k��>̛T>K�5��n�=��<��==Xܑ��)���\����\��S�I?_C���"���꾷���hA���S�����>e�>Hd��w���Î�;�>̿�=��{�3̲�y�`>4��>4<>��>���
����sRY��A�=�Y~>�6�>�Q\���
�G�x�Yc>�3?ֈ�Q��>q��>Qz;?�m_?=��>��ƽI�?�s�>��=�[�4�n>�`�>?��={�?Ar=?F^=?�G?I��=�<����>^�">	<}����m㑼j�=�Իw��=��_�e���V<��=��@>��y�����5/>G->&K?u)?V��>���>����(^���	��)X<3�>��<�3g>i:�=o)?Z��>�]�>>p>�<F���e�ɾS�?�9<>0+���Rz��=��/>OW>�i?S?��Ͼd=��q>��H���>D��>z�$?�9?w�>���R����ҿ�$�5�"�p������X�;��9���G�dҺ�0�G�ｐ�<�V>u>�>�8t>l�I>N�>�+>rS�>�I>��=�v�=��;�R�;��W�E�U=H���)<ڍX�E����ԯ��ࡽ嗊��K�*B�V�������J?�?���<��=�g�;��X���ƾ�^>���>5�>^��>v��>Hf��c�:��D�=z�R?X0b?�+�>,�4�D� >TN(�Ŵ�=(?�z�>�c��s?���P>p|��v|U�H�3>
?
?r��>'���J+1��0K����]�>`jͺ �����?��c?���E�o��"Q��f���qg>�����O�z����4{!��`��Ԧ徳���Ⱦ>M?�?Q�9�el������`��R�n�]G�=�����"�>�..>]_�'H��i�ݾn�Ⱦ�~o��/�=��=�>M~�>}4'?�g2?_b?��?���>_S^��?K�K>J̪>DA�>��?(�*?�w	?�v>.^>�/�=:�<�l�%x�����=傸<5 �<���=�'>��y=@,�=�З=;=[;<�����
p���U=�Q�<�5>I�5>�[:>:i
?(-?���(�=�y�<�wb��� =pi�=w3�>U�U��Á�Y�|��>/?��)?�)�>0�=�m�����b�	��\K=L�&?�)?���>��>?�>���Y��B(>�W>T�ȼ��Ͼ C��;���j0��\�>�6�>��=�;�=s^�?�Z`?@V�>%�!�DR�S���Y$V�2����G>�.>�$?y��>hH�������.���\��!2�$���먽���=J6>��r>k8>,b�=�8>��н�t���>Q6b>�al�	��=���>�>+�=�|��қw�D���kN?�_�����ϕ��Ѿ� G��>��G>���S��>W���`s��-����:� �>ی�?���? 0g?{M�]f��*?S>=>�>�0L=x���8�OP��j�8>	t�=�f�Bv�D��;V�J>�#P>���*V����վ��\��}��y}����
c���پS籾�*)����!t��������{�WN������ܺ�<_�;��=HxU�|ZԾMľ��a?n��?6�=*yԾ�J���ט���C�=-L��9e�Ñ���=�I���Q��������ٽ��A�57�D��><�@�����(��*�Ⱦvx�=��=��_?|�vL׾E�^�]�u�7���5�=uO�撿j�� �D��WI?m�-?���SҾS诼��=%��>���>LA!>JS��U�_=(_�>0�?_B?"f�<�?��2����=nE�?�D�?&�"?>cb��P��y(�r�����>:x"?��,?�[��bϾ�G�=���>��>?��>D7�Y棿������>]�z?��T�:6g>�8?���>fl������^d�>�� T>��^=�B���c��)�<T�����?�>z�>x�
J�����>E�r�N��H����\[�\�<�}?T���z>�Ei>�>�(���D׉�����L?���?��S?�J8?}1���t�YM���ڏ=X�>�>V��=���,Ǟ>���>�a��ir�J
���?�7�?���?�JZ?+�m�cGӿ8��0���������=�$�=T�>>��޽ʭ=:�K=u���8P=�̉>`��>Oo>�;x>W�T>r�<>��.>T���g�#��ʤ�#ْ��[B�� ����tvg��{	��y�����ȴ��񽾉�������ѓ���G�r���U>�6�� U�=�8�>*S+?��?��>��>�g�k�;�vy<��L�!tF�@����N-�����#�������߆��$G�,��~ظ>�]=��->d��>c��<�@1>�x�>)�&�$)���&>MR�9i�ֻr'�>M7�>%A=�4#�,�`�K/M>�m�=��t�l���]2J�@!վ�K>-]6?�˼�{�Xd:�*��%�˾�~>W�?�ܭ>Nh��2��b�����>itu;�����2�P�>!~�>�>�	d=��:����aY=�D�=��>���>�A�� 5ؾ,ڄ����=�t?S��,>��>�Q�>FM�?r?��=.?&ݷ>�����q>�ȭ>Q�>���>�?\�K?�%?T��>�L�=ϒ��_V�����=�+��Ih���Ľ��a/���<x��gQ	�}|㽚v=k}d;�a$�:Dd=�y4=W͘��*�>�}u?ϴ?��d>�ڦ���Y�5�J���B���>�|�=8V[>��?�F?���>��>:�1>�=��־����>�=(�*�춃��ξ��7>^��>��\?�)?]e���U��e:�>v�;>=.�>�|5?+�Q?o�>3��sj9�\`��lƿ�.L��ﾬ½��~���B��/<���0{���>b`ľ�Ծ=�ܽڼJ>Tt�>)�~>+L�>c�=8�?z!_>�2���;>����>���<=0�<�_<�E�i�'���=5��5iX=ޙ���J�=<N�<ܫʽL#��W?�?n}K��2��.m��M;�`��X�>p��>N ?���>ޛ%�kR���<���N�ց���n�>�w?�?}��g��=�6�<��=��>�,}>͂>���� �Y�^%��������>���>d��>.�
�_��y[�>�L4>+*Y< �'�?Qk^?e⳾L�8�W�,��L_��� ����=��)�w������&���1�Vv�rU%��j3���I>E)�>�T�?G;�C�=�;���~��f����.�=�='��>�[�>ƭ�e�?����{����þ��=�܈>�Q��d�>�T?$�>?X`4?B�+?Vq?�ě�ZF$?ߗ#>/��>�{�>m�>�?'\�>�?�?Cս&���'?������(��
n����=� e>�d*>��=gb>�al=��ؽ1D=��F=�Q�_+H�y��=�F�>OT>��p>(�>/D?6!�>u�<�[-�B)��J4��u�=���>�@Y�|1��»�D�7>Ar�>��:?�k?����`%�\�پ��O��ڽf1.?c�6?\ ?>b;>@��=�	���6���=���>��˟��4�M�W^R���H>2�>��7>g[P>C�?P@E?y6?�?��шL������B��"�=T�E>���>;�>=}p>}�W�B���\��e����v�F<�(�*A>��#>k��=�>�Bf��1t=/s�<�5�=M��k"=���=Wr?�v�>�8�>�w>MG�>"N��x}�<n?�������ͫn�^���|�=њ�>��[>]�=
�?�$Ѿ+�R�	�������	�?�}�?wg�?^�0?���F\��NA�>���=��¼a�>9�˾��Ͼ��U�Vo{>��(��Y�=_�����H��Ǹ�q>#!�=���n$����=�y̿�l|���Ǿ��̾�E�]:��;�о�ͺ�
@v�כ�#�
��H���ƾ��G���Z������/�Y�͉����?�'�?:;��U���2��'�7s���f#>�鮾uQ*��1e������3����Ѿ��j��k�e�8�YD6�E����>��ý����vR�����
x���q�>�?��þ�S�}�*��+�>#�&>�<��ŹAm�����ˈ���? �.?R)�i/���<>��>��O?�Ѱ>�E��c��v��>:I�>*��>��?�4
>b�������*@>��?�2�?��<?|@��|�b��h�-�=�Y=?qv>'�>E������&>���>� A?���3"V�񎊿������V?�?q��ە >.?D�>�Ϻ��h��=������ns>}�Ѽ*���������=�|�>��>��<U'+�P�>���F�%o?�� 
�Z�0���<j&?��a�=�׀>� >}#%�Gt��*���
�̽D�Q?Ծ�?.�G?�5?^�󾉃��چ��%u>~A�>*9�>�`=�� ����>c��>t|���fk���NZ�>	��?�U�?-�[?�Fk�˒��<[���Z����/�~=���=�8>��W#b>Pf�=��b>����$�=�4�>O�B>+8s>��~>�>�׀>�E��T��C�ÿn政��C�3�5�P/��!D���پ�1ྥ]������1��}u{=�y�����Ꮎ����0�X��9�`(��m�>r��>p&�>2\�>��!?�%��T�*�|ݤ<������qE�ɡC�@(����R�˾�S�����=�½>�/�-��>��n>?��=��?�ߪ���R�"��>E�>x�>�.>�77>N��=ͱ >k��>̛T>K�5��n�=��<��==Xܑ��)���\����\��S�I?_C���"���꾷���hA���S�����>e�>Hd��w���Î�;�>̿�=��{�3̲�y�`>4��>4<>��>���
����sRY��A�=�Y~>�6�>�Q\���
�G�x�Yc>�3?ֈ�Q��>q��>Qz;?�m_?=��>��ƽI�?�s�>��=�[�4�n>�`�>?��={�?Ar=?F^=?�G?I��=�<����>^�">	<}����m㑼j�=�Իw��=��_�e���V<��=��@>��y�����5/>G->&K?u)?V��>���>����(^���	��)X<3�>��<�3g>i:�=o)?Z��>�]�>>p>�<F���e�ɾS�?�9<>0+���Rz��=��/>OW>�i?S?��Ͼd=��q>��H���>D��>z�$?�9?w�>���R����ҿ�$�5�"�p������X�;��9���G�dҺ�0�G�ｐ�<�V>u>�>�8t>l�I>N�>�+>rS�>�I>��=�v�=��;�R�;��W�E�U=H���)<ڍX�E����ԯ��ࡽ嗊��K�*B�V�������J?�?���<��=�g�;��X���ƾ�^>���>5�>^��>v��>Hf��c�:��D�=z�R?X0b?�+�>,�4�D� >TN(�Ŵ�=(?�z�>�c��s?���P>p|��v|U�H�3>
?
?r��>'���J+1��0K����]�>`jͺ �����?��c?���E�o��"Q��f���qg>�����O�z����4{!��`��Ԧ徳���Ⱦ>M?�?Q�9�el������`��R�n�]G�=�����"�>�..>]_�'H��i�ݾn�Ⱦ�~o��/�=��=�>M~�>}4'?�g2?_b?��?���>_S^��?K�K>J̪>DA�>��?(�*?�w	?�v>.^>�/�=:�<�l�%x�����=傸<5 �<���=�'>��y=@,�=�З=;=[;<�����
p���U=�Q�<�5>I�5>�[:>:i
?(-?���(�=�y�<�wb��� =pi�=w3�>U�U��Á�Y�|��>/?��)?�)�>0�=�m�����b�	��\K=L�&?�)?���>��>?�>���Y��B(>�W>T�ȼ��Ͼ C��;���j0��\�>�6�>��=�;�=s^�?�Z`?@V�>%�!�DR�S���Y$V�2����G>�.>�$?y��>hH�������.���\��!2�$���먽���=J6>��r>k8>,b�=�8>��н�t���>Q6b>�al�	��=���>�>+�=�|��қw�D���kN?�_�����ϕ��Ѿ� G��>��G>���S��>W���`s��-����:� �>ی�?���? 0g?{M�]f��*?S>=>�>�0L=x���8�OP��j�8>	t�=�f�Bv�D��;V�J>�#P>���*V����վ��\��}��y}����
c���پS籾�*)����!t��������{�WN������ܺ�<_�;��=HxU�|ZԾMľ��a?n��?6�=*yԾ�J���ט���C�=-L��9e�Ñ���=�I���Q��������ٽ��A�57�D��><�@�����(��*�Ⱦvx�=��=��_?|�vL׾E�^�]�u�7���5�=uO�撿j�� �D��WI?m�-?���SҾS诼��=%��>���>LA!>JS��U�_=(_�>0�?_B?"f�<�?��2����=nE�?�D�?&�"?>cb��P��y(�r�����>:x"?��,?�[��bϾ�G�=���>��>?��>D7�Y棿������>]�z?��T�:6g>�8?���>fl������^d�>�� T>��^=�B���c��)�<T�����?�>z�>x�
J����>��便�L���E��/���.���< ? s��x�
>v@j>$!>*A$��<���f������I?�m�?+�T?&�/?ѫ�q7�����JV�=���>e��>�.�= ���S�>���><�dTr����;?��?f{�?�P?��s��	ٿd9��x��m^��y>f�U=�>�3T<N�<;޼�j=?�=��>>y�>zщ>�>:̀>o%�<�k<�"������v��¼��A�>>�eJ�7)����;n�d��m�����Ҿֲ���콧Ѩ�d�/���ǽ`ὔ�ƾ	�=��>�y?q9�>�<���>�4>1^1���?�<�e\������n����E�3�rQ���9��`�������<?�T�<�.v��3�>2i�^Z.����> �k>��=ȩ�=�O�GJ�=n8�>�)�>zټM�>r��=�jG>�=�=>���m��Q�jwþ�5��9�??��{�����Z���ƾ��J>W�?�>�2*��і���o�U��>x�$���o餽��ݽ�Cq>�>��=U���D��cɾ�S=Z��=Y��>�g�=r�7����e�b��=�<�>dY�j>�k>�vF?8?~?��K?�7e��a�>�
�>
7>�b$=�4�>߉�>�O�>=�-?O�a?�A?5��>�-�<�~�����=�9�>������5�����T��^�x����dd���'>X��>*"P>��=�I�v�0��<r{�=W?6h5?�?IH�>ߠ]�S��57F�聾 �>��>�z�>4_w>5<�>je?v�?-�>�&
>�� �483��-�>��~>D�V��"��Գt����>��>>��s?�U?��s>�嘾�:�=��+�u2?���>Ծr?C?w��>�_�<!��ҹ���$�ݠ꾭� ��=μ��>p��r�=��@=Y>
��ҽ���$�M> �>+�N>e�x>-� >Qm�=^s�>אp>k�˽�*<��X���A�<�"�=���=YHX��`�=���=����ٽ���%ؽ�p���b�u��<���=�?��?�#�\!��;L�������6#�>ŀ�>��>���>�`�=�9�i�V�E[?�$�F����>')f?N��>j�S�Cy�=+*L�Qq�<�Z�>�[�>*\4>+(��R9����V��<�}�>�L?���>�(��yR���g�}��X �>Q�=J�x���?��G?#���%.K��^����A=-`=ƒ�U�.�=D���6�sϾ�j>��X�\>�]�>��?���!	罳=X�� m������}��45>Kɽ}��>Y�>h6�<L�,e��Z⾖Ǿ�����>�2�=��>?�?�7/?��v?��?�V ?�:y�_ �>��<�Ĭ>�$�>�3?��6?�?�{�>��>r�	>�����u�7Z��IQ�=!��=��=�'=��=J�Ѽ��*���w�v�<�c\��偺y��=�s&=�*'=@��=���=���=g�?̒*?<.����
�=ǆ�����=�:<6{�>�	'=�˒��A �r{>,k?9�A?�m?}ik>�Ι��h��	��2�Y�
�?��8?+��>����*(>��谈����=�qY>��9��&��p��4r�9#��خ>Q��>�"�=�6m>�u?��<?,�r>�wK>Wn�\���G��}�=b��?�[�>�W�>�־��9�$�)�8uA��6_�4�D=[ U����4�=���>z02>�x<j��>����7H��m��dvU=$B(�u�>�R�>�7? �+>���>�{�E�B�C�V?�X�-Y���J%�&����*�>���=(�=��>|}c?�dj���{��߬��ʾ��>*��?���?`bQ?4Ȣ����F>"�^Z�=</v>|���>(�ֽN�%<�:�=��$�	�K�L�=|�`�t��=|�B��c���S���k=�(��W�8�fa��!E��E�a5�!0��{1_>�;Z��j<�mǾ�ݽ�W�Ǿ�\j���=v�r�S��񨙾����|�?�b�?���=<V��+�A>0�������=��>�Z�ҽЧ$�s�����LK��v[��A8 ��/6��4�^\�����>S�y��,��pkP�E�j� �a��bj>#�K?0N�����gav�
�?��>-� <�a뾵g��I����w���Q?�C?��b� ��f�>G7t?�>�>�R>č�s?��ߕ8?��?D�%?�B>5ԑ��S��W�:�
��?:��?�_L?z;��-@W��f往qT�/u�>,[?�5?7��$l��7�=ʏ3?p_G?��>\=�b#��Lm&�IV?޺�?7����ۻ>K�?�a�>�T=���v��;�:%�
�9����>��=G�R�9�d� ޾�!�=���>��>�<M��B�����>�����oP��?7���	�D�p��b�<�H?u����v->��>S�;>�w,�����T�G�=�@?,è?�gZ?��	?�P���B��ui���>Z�r>�^�>��=\�g�{��>���>#��#|��9 ���?L��?M��?0?�����տ�E���+ľj�Ҿ�|�<�4=`��>�V���\�^�V�S�μ�/C;��Y>���>���>�h�>��o>�o>+�>�+��Ǧ�s䳿�墿�C���X���8������KB�iӾ�Y���>�o�={������Ἐ���Ѿ#�=o�{>���>FO�>�
�=�>��e�$�J�Sо>����ٶ&���!�Y
�O�;��5�l"?�4�T�:�Ž\K	��7?Ė[=�na��?b篽q��=�)�>UֽK��i��=�K�=qWa>��'>��>8'۽��>U)�=�}>��;8��cn��a��:�c{��RB?�_��I��}�V�u୾T㩾���>�?!�v>G-=�PJ�����V?T�	鳾:�j����<8��>��l>Vw�>N�`�⓬�7`���#�B��=(GW>��=�Z;<�*���8�w��<�#�>�rվ�x�=�Jx>��(?��v?(�5?�/�=�Y�>;�c>vu�>A��=�0N>�eQ>�n�>=U?�y:?&%1?�D�>�=	�`�c=��A=�>�hY�G`�����Z=0�Q��<l�,�j�G=`�r==�<!la=R�@=������;lv�<�_?�qU?'6�>j^�>>�c��W���R�s�<���>������>N��>�:?�P�>�� ?x�>��J���1������>�4'>�G�oҋ�z������>��%>r�K?<'j?�۽�s�*��Lp�>I�?�)�>��X?��F>���<�M���	�{U���d0�h^D�O�O����j�>���i*�֍���dܾO[q��qv>^�?n��>F6>�n�=}�>I�->��>;�_>���=���=��׼�H��"A���*�<��a=ŕ!>G����}���A��
Ͻ�����޽��b�����<�;?|A9?1��=5!��5���wP�Ӈ�V���V�>��C?Q��>ΨӾ��5�S3��d�|����=�=:^�?�cT?��˽&�A>��N��x�4�=$�[>��>�I)��S�=�B�&9O>��>q??��>��_�R�b�kJ�^Ѿ>��=��T��?�UE?-����>9��\A� ���ͧ=���`(��g�%�r{6� j���"�������>�I�>?��?}6��2n��������/��y󝾁��=fpR=Ϙ>��>����t�����t���G��Be>{��>P�7�5�>��?�?C�b?f?��d?,�Ҿ���>Q��>�M�>��Z>�:<?���>b9?r?[I?���=T衾��x� �>) >C��=[26>�x5>�4�r�`<�߽e�.=+y�:�h�=-<�<&�ټ�o=���=��a>
�3?�-0?��<��\�S�%>�>��)����>Ҧ�>I��>	0���ۼv=�>�M�>��%?��N?���>oξ�u3��5侹�t����>�H)?�w�>g��)�>��	���񾎌E>s��>kw<�d*��7׾Xf�P���f?�a�>��F="2�>��s?y�?�/?mo�=�v�F��2��(E�=!i���'?��?F��=(=;����6\�DZ/��-�$޽��x���x=�����>`�>I���uЍ=cÆ>�������K�>S�T=�O>��|>�}P?��>��=}r�e��>�I?�����a�k�Zо����>��<>�����?{����}����9A=��|�>Ԃ�?���?H2d?~�C��G�y�\>�>V>��>!�0<�>�NK�tڅ��3>#�=ESy�����V�;��\>RBy>U�ɽ��ʾ�供 I��]����I�8����^ ��D�hc��Aɽ®�;5 O�XZ^���h���rp�/S=��=�s��G��7��� `��%�?�eI?s��xz=�b4��ؾ�^�U�>�L����\=�)��/�<y������y)��3�%�F	F������>�s�mL����w��6�`�>;R/>C?����ѾQ���m>�r,>�p��������њ����??B�0?�͇��أ�d�>4�	?�m�> �/>��@񅽵��>�C?�`5?@gG�.8���鯿���={��?u��?3�K?��ھ[�5��Á�H�?о�>*5�>�{��fٴ��ZD=G�4?l�*?ֈ�=#'�B6��^g��
?|ƈ?�J���c�>�
?Wۻ>]�����|���d͎����4��>�R>_�q��;þ*'d��K���>Vy�>v�߽w�����>�����oP��?7���	�D�p��b�<�H?u����v->��>S�;>�w,�����T�G�=�@?,è?�gZ?��	?�P���B��ui���>Z�r>�^�>��=\�g�{��>���>#��#|��9 ���?L��?M��?0?�����տ�E���+ľj�Ҿ�|�<�4=`��>�V���\�^�V�S�μ�/C;��Y>���>���>�h�>��o>�o>+�>�+��Ǧ�s䳿�墿�C���X���8������KB�iӾ�Y���>�o�={������Ἐ���Ѿ#�=o�{>���>FO�>�
�=�>��e�$�J�Sо>����ٶ&���!�Y
�O�;��5�l"?�4�T�:�Ž\K	��7?Ė[=�na��?b篽q��=�)�>UֽK��i��=�K�=qWa>��'>��>8'۽��>U)�=�}>��;8��cn��a��:�c{��RB?�_��I��}�V�u୾T㩾���>�?!�v>G-=�PJ�����V?T�	鳾:�j����<8��>��l>Vw�>N�`�⓬�7`���#�B��=(GW>��=�Z;<�*���8�w��<�#�>�rվ�x�=�Jx>��(?��v?(�5?�/�=�Y�>;�c>vu�>A��=�0N>�eQ>�n�>=U?�y:?&%1?�D�>�=	�`�c=��A=�>�hY�G`�����Z=0�Q��<l�,�j�G=`�r==�<!la=R�@=������;lv�<�_?�qU?'6�>j^�>>�c��W���R�s�<���>������>N��>�:?�P�>�� ?x�>��J���1������>�4'>�G�oҋ�z������>��%>r�K?<'j?�۽�s�*��Lp�>I�?�)�>��X?��F>���<�M���	�{U���d0�h^D�O�O����j�>���i*�֍���dܾO[q��qv>^�?n��>F6>�n�=}�>I�->��>;�_>���=���=��׼�H��"A���*�<��a=ŕ!>G����}���A��
Ͻ�����޽��b�����<�;?|A9?1��=5!��5���wP�Ӈ�V���V�>��C?Q��>ΨӾ��5�S3��d�|����=�=:^�?�cT?��˽&�A>��N��x�4�=$�[>��>�I)��S�=�B�&9O>��>q??��>��_�R�b�kJ�^Ѿ>��=��T��?�UE?-����>9��\A� ���ͧ=���`(��g�%�r{6� j���"�������>�I�>?��?}6��2n��������/��y󝾁��=fpR=Ϙ>��>����t�����t���G��Be>{��>P�7�5�>��?�?C�b?f?��d?,�Ҿ���>Q��>�M�>��Z>�:<?���>b9?r?[I?���=T衾��x� �>) >C��=[26>�x5>�4�r�`<�߽e�.=+y�:�h�=-<�<&�ټ�o=���=��a>
�3?�-0?��<��\�S�%>�>��)����>Ҧ�>I��>	0���ۼv=�>�M�>��%?��N?���>oξ�u3��5侹�t����>�H)?�w�>g��)�>��	���񾎌E>s��>kw<�d*��7׾Xf�P���f?�a�>��F="2�>��s?y�?�/?mo�=�v�F��2��(E�=!i���'?��?F��=(=;����6\�DZ/��-�$޽��x���x=�����>`�>I���uЍ=cÆ>�������K�>S�T=�O>��|>�}P?��>��=}r�e��>�I?�����a�k�Zо����>��<>�����?{����}����9A=��|�>Ԃ�?���?H2d?~�C��G�y�\>�>V>��>!�0<�>�NK�tڅ��3>#�=ESy�����V�;��\>RBy>U�ɽ��ʾ�供 I��]����I�8����^ ��D�hc��Aɽ®�;5 O�XZ^���h���rp�/S=��=�s��G��7��� `��%�?�eI?s��xz=�b4��ؾ�^�U�>�L����\=�)��/�<y������y)��3�%�F	F������>�s�mL����w��6�`�>;R/>C?����ѾQ���m>�r,>�p��������њ����??B�0?�͇��أ�d�>4�	?�m�> �/>��@񅽵��>�C?�`5?@gG�.8���鯿���={��?u��?3�K?��ھ[�5��Á�H�?о�>*5�>�{��fٴ��ZD=G�4?l�*?ֈ�=#'�B6��^g��
?|ƈ?�J���c�>�
?Wۻ>]�����|���d͎����4��>�R>_�q��;þ*'d��K���>Vy�>v�߽w��p�?ډ&�U�E�W�'�� �����b����Z�>����I>u>5>���=L�Q�g��j
��-?޽:�I?�\�?1Xw?6�?�8����������<P\�4��=a�='R�ۉ�>���>���`���!P%��R�>1z�?���?�{p?Q����οj)������4��-Y>>:S>'uսѾP=�q= X�<��\<6>ؽ�>-k>_!g>*E>5>D#>� ��8�"�1`��|唿S%>���������}�Z�!�����f��d;þ������a�x�?�m�L��~,��^j�a�Nwv=d��>I��>��>,W��@V�>N*y�3������d���2!�8�9�F�%�{��	���
-��x����뼌;m�Z��7I?_'F�h@�=W$?��������>z2;�S	>��>���>-�>;�=�!>4�=�d�����=o��>�w=�j}�(#c�����p��*�=3&c?$Th=IkھMD��C�a�23a=+��>Ҍ2?9>�EQ�ͤ��������>��i��恾+}����)����>���>jc�Vצ<�{�=(��'>���w�Ns�>��#>t;��x��3��U����>3�վ�)�=J#{>��(?��v?��6?�K�=��>�`>�;�>��=N>`ST>Nj�>��?��9?��0?g��>鞿=Xd��6=�M@=��>��^�&Q��|��8&(�V�<�1���5=2Eh=��<qh=�!J=<-ü���;�k=<y?��S?�a�>ۀ�>#�3X���4��=�>��7�y $?'x?J,?dP�>K�>yʕ��ԓ�p� ��M��[��>�/>��J� ���-/����>�'�>fCi?p]?Q �pؾ�t>0Y�>]/A?�$S?��=?�;�>ۢ�=4��&���ο(��_+�8ޖ��G8�)q��]�5�������� (������=��[>gޕ>,��>">Ʒ�=S}>*��>�>�U=x��:٨�C᡽�66�&A>p�=��û����^z����<c���
Eӽ��ܼ�8�\#�<�^B��k?F�?-�������tx�Ё۾��	�DO��w�#?��G?��?|߾<+�
�W�)�T�w_��*��>ÿ�?�N�>4F��9�>�sE�#�o=��3>{Y>��O>@�=�n�@E�����=�7�>/�(?�Vw>Z��;�{u��{���,��
?|�H=�����:�?4Q?} ����tG�;=��p���=�P=������ۨ����]E�=�۾�Q�![��f�>��?>ș?�뒾��)>��Ծ],�������.��򌵻�-(<G��>l��;%Љ��ci��|;���#�~��.�>豛>O���A=��W?��z?��z?�-?��e?k���>JF�f�>��?�?��E?�tC?$��>Y(�>�l�8���d3���Ѿ(�,=[�=��n=%ر=�.>�h�=�R�d��2*�=�\�<'ǿ��,�� .h<��˼<�C����=��,>%)?g/l?_�	����B�=MC�>��	>�|���I?���>.��[�>���>�5?P+9?ݬ?�~>�_!�>6����qc>[�?kH?x�$?�˼������T�ž2l�=ļ>�t>=+co��	;lپ'�νڟ�>"'�>��>>�Q>�d?s�?�i>?sV���I��*e�
^��V%o�0'�:�?�+>7�R=a�2T@�]򋿖�l���5� �M>2�p�] ���i=o��>%hg>�%���>��=uI�����c���mM�<���>C�>�?�A>��<�����T>?f1�������h���Ѿza���'�]�5>�B�?6�>^�[�c����1��Q�X����<Ҷ�?}B�?ng�?�BY��)q���>8V=�:��x�
>Y�����so|�+��>�i+>��B�.��KI�=���`G�>+i��SȾ�!���7�طͿ��=���۾)��@�?~��|쾏rm>�F�項�^܅��)�iL��0���;�U���8�]��b�?ե?rK`?>B:�h3<b�4���2,�H�>!��%�B�;����4�~��_z��ai���[��(���|�����>ӅѾ�$��qz���E���m=Ⲝ=�:[?Q�\��w7,����=��>�8���4ھ�.��_��%��&C@?hI?� �� ���ɽ�֏>��3?�ܺ>tSs����/�<+Ӛ>0�4?	��>����Sި�����S`�=�;�?e�?��B?(�|��*M��r
�A��-M?(��>7�>􎖾ڊо��Lp?��0?���>U�m"���:"�W��>�j?�q;��td>& �>��>�H~������ا�� ��1�<���o>�w�<o��S���F�s�i}�<D�>!�> <��J��|�?�1�LHc���8�#]�� �<��R��C
?Τ����<4�>�g>!0�����Lډ�R�:�R#0?*��?�ۀ?
?ֆ�Uvh��ϼ�勨=ju�]>p@�>���p��>|]	?	���ލ�uT�	{�>Z�?�r�?"z?�'������I��(8�����B>'<>�ME>8�|^����t���Ӕ�H^Z<�?�>
V�>��">FF�=���=E�>�H��m��"=���֊�,<�Mg
�t�K�#����e���!%����fu���$�{,�����Q@�2�Y�J	��0󾊟�=`P?~!e>�Z�>s��=�>�����#���x������>�&E ���U���!��"�����T�=҃�-o�6'%��"9?m�_<_i->�e(?��}���ǽ{
>_'��!I>�Ti>�N">Q��>�=D>��E=oӣ<N_�=��<~�>Z�="�z�o�p�� \����ϻ=y�g?�C�<����K`��X���K>��>�d<?�p�=fR��������-x�>�[�Mnd�r�>h5��>'�?�T$�!�
>P_�=�[�<���>�ݴ>6l�>�|���<h����9�'�ڊ�>P.Ծ�f�=k�v>�c+?��y? �8?,lY=��>��`>Ж>$2>�G>P�D>��>H�?qB=?D.?#�>B��=	�]���D=�1=دE�Khp�[����߾�J�@�c<��)�U�/=�>O=��9*L~=,%8=�V켘�<�G=zd?��G?�`�>�Dq>ڧo��R�2N?�\�G�,�.>����(�>Л ?��?�?=�>Żq�������c<��D��>�Q�=,I��͐�>:���?ix�>��n?�	Q?B½�vվ��>C>�>Ѹ-?��/?�C?-_p>���=�N�����Iտ'�#��g$��ZA��뉽ѻ������̦�Ri�v��:�g>:�>��a>~>�b�=rq;>���>�sy>���<�H�<߃N�� �rf��M�&>}0��Å���@��):�����0r����*�=����F�2�缀;��h?m��>����G���12�D�
��]��0?�v?�l?��R���(���W�(oR�29뽃�?u�?+��>����N>�l�=)d�=F>n�H>w�=�bS�D�Q�p����B�=4v>� ?Ш�>>@��B&l����3�e��-�>�}=7�־Q��?N�W?;���n���(��9��7�8��=�h�'i�y9��>)M����=�׾��Ox�>|�?��?כ���>�ؾ�/���R�������N>Y��<]b�>�I������|�5��3(�u�q�58<�p~>�=�>Ѱ�3ܦ> o?�{:?l�?M�=?9j?I
�{�>f�>��	?+oC?�Z�>��?���>v_�>��$?��f�Y�����%��ϝ߼���-����!>�8>�M�=��<�瞼�c=�x��.��y��ؽq;�83>�(><Ț<<�$?�O?���o�X�y<>�=E�!�T�>�T!?9��>�ף�[}̼�T�>��G?H|?Ϗ%?-�g��e ��(����(bx>�S?�Q�>~!9?����������j���>{�>2خ=Y擾�6���Ͼ���K%�>���>��h>��>Llu?f#?�_?��R=��`���x�i�G�U�	�9���N�>�Y>�?�<�̾���s����v���G����=��#�f��=3K4=2�6>��>#d���>�o>�WM�Z�x�n1�ù�=`[�>���>��?y�==��{�þ�����A?�r���y�-�X���ܾ총��>���e>���J��>����6�����Y�a�A]�?#�?��?���	2O�X_�>�=Dm=�=>�2�!>�$�����>�v�>o��
�W��[�=m̈�N�>���񅑾D�����v�����C������*�D꾖὾״�����> � ���5�N���d���ܢǽ5�߽�~�=8V�Bn�����1��?��?�ք�����
5N�������׾�á>w���;��MϜ�K<�-=G����n�7��e
�A���6�>ve��`��l�{�^(Q�(�>�M>�J?�ľI� �Ju^�c>jӫ>���V�;�穿򾗿Wfn�.�]?1mH?VW�h��v2��*0a>I{@? ��>@��P���Pږ����>�e?LC�>���i�����b`�=(��?��?8.A?W��D��>�'�ra?��	?�)�>�)��Vξ��� ?"::?�>ao��酿#��֍�>�#_?��H���_>F��>�]�>[i߽A"��AUM�Bݓ�%i��C>��y;.W��zz��)E�U��=ņ�>�͂>��H�'��"��>z��L�"UG�X�A�(���<���>ْ��=B�=VDP>�(>y�#�����������D�R?�h�?�M?�X.?4��F�⾫3��]��=���>�Ǜ>���=PD���5�>~��>�2��u�F�	��
?:�?�*�?A�_?1i��N��~�������y����G���l=�B>>�rg�{�>hF�=Q�=?���_�=���>P/�>%_�>�>dv>��(>B�u��%�򡸿o����^�L��=�����(��({�M��	6�r�۾�#���Oi=�O>�	>��P���B�Q|n=��B��>�QO?ǉ?^A�>,��=�T̽�x��q&��f�<�D��WUξ4���=�IY��e"��� ��.=������ý/M�����>�;=Y�/>��W>�R����>1�>�	�<�X�<�U����=�`=N�=�{\=8}>h�v>�\{=u=N>]
F������%����:�E��}�@=˜1?n�=u���"/�2��#���Hӭ>��?.p�> ���Ë��t<����>�V���؋�ɂF���=`��>� �>J)> ���	�}:̊t���t�Y�=ݖ�>�V>ZQ�����_�.����=�@�>Uھ ��=�Il>�+?�
s?Y�2?�l�=�R�>��X>0��>�x�=Gdd>�,P>X`�>k�?L�<?�t*?z�>���= \��	=�`=�\��2M���˝߼�4M�~��:��!i�=��A=���^$p=I"�=�g���$�K�<�A�>�Z+?�8�>�1q>g��k�,��ώ��)����=���T{>��μ���>L�U?Y5J?Hy�>�By�9�-���f>Ix?�8y>KCK���F�J?�=e%�>�b�>�&B?��7?���=zӓ��d���.�=1��>�T	?F|�> 3Q>Yw
����=-���.ӿ$�#���!��҂��+��J;�=�ZP��?�Ҹ-��X��7/�<{�Z>N�>��o>w�D>7S!>V2>��>��F>��=P��=N��;��;�PF�\LJ=�d��	@<��P��1���Ƽ%��𹌽igM���A�#$���ټ�Z@?8�?������$��B�"�����U?Z��>&�E?^be?]�K>�Y˾��g���T��9ʾY�>�e?�?���=�F�3����)K�R�>�>��>��=QH>??�@�A>�?�B?��>��P�eLw��7���8��V�>�A�=Ff�N�?�BV?��	�����[$�QII�%{����=m(Z����E�޾��)��W��N������i�f��=�)$?Sz�?��ݾ��;;:ξ�J���Qe�'��I>>�x�=r�)?�]�=�c;�覽pǾ����Z|�l��=��>c��=C�>3?��?�b?��?,�?	��W?�F�=?-�>/��>)?js
?P��>E�~>�3~>��=�2�p8��(���)<+�Ǽ��=�>3K'>��f<1=ۧ;=(�<�=��V�7��<� 5<�=���=)��=��>vl?2A?�YK�=oj
��Ĵ���>��@>��v>��K=U��ͮ�A��*,�>as(?��*?1=h�1�Noc����&g>��>?r�k?��[>^ua�����Ͼxc��ƨ�>/{�;�k<����%�r�龏�o=�#�>
��>6/=[�>wφ?�B?|B?���� �/Z�>|:���@���)=���>��>���<��Ѿf�2���g��p��`:��ƥ�3y���R�=1��=�h.>c�@>�8�=�e�=��)�'o��`#���&=�J��I�>(�>M?��)>x�(=Gv�����ҘF?�u�����	�����о7�@�փ>��5>P\�iH?on��#|�[���V<����>�s�?n��?��d?��C�w
��(a>��Z>$�>G��<�W@�q�A�=�R���6>��=�Vw��图©��6K>�o>�Bƽ�Jɾ�پ��N��t��֏A�>o޽�Ҿ������پ` Ͼi���ē��Q�w�޾�ju���r�&5e�w2'� �%��g��o6�怴�^)�?`v?6��=�
a�5 ���a㾶G=S{o�!\��ݕ�v�~������Ϗ��fK�-:���#��v �@Q>���9ᢿ�{k�Mت�.�6>	��=A�>?r����}��4�*��\]�cMy>]��>p0.���u�����A?<k�W?�0?UAfi�_�9=�m?��>��>�`g>�.��>B=��@>�$@?kU?��=9喿����) �<
��?���?`1E?ӱ�~�.��)���=C�4?��-?F@�>�Kj��D��D/<:[?��{?��>��γu�����/>l�< (��{�>��>�Zv��{ɾ�Gʽ������e�&�u��:>E1��%c<^x�������=���>��>�v���=>��Xm(��U�K��� ���Z�Oe?��!��a��gq=���<G��[u�X݇����>3?G�?F�v?A�X?=���P���Th=�}���k)>-?a'�=C�W<�I�>�j>1?	��8U�� x���)?g�?��?<�u?��Z���������?���g���<M>��Ǽ8@>���=�ץ�ߏr�c�=J}a>HOd>�^>�z>۷;>��
>޴���i��~#���wO���!����,�]k׾��d�j�eS��۲ʾL�Y���٩�Ħ����*�;���b��5w�>�6?�==?	�>�>	�=�I��n�=J���1־P�uV&��տ�~�S���[�l���j����ɽA7��;�>��{��Y>���>e=���'=>0�>�~�=���>Ds�=�]=ɗT>M5�=�>���= "�>��>W�o>��^����K�{��8�\f�4Q<\F?n	����r;=������ͫ�#*�>)w?C�>#��[�����M�>��>nW%�͐���u��`�<�M�>���>�ѭ="�d��z���Y�T��|�_>�
�>�u>���ɚȾbj�gE�=�7�>� پo]�=-�\>X�*?��[?��$?�H=��>I;>�p>�n>��8>I>���>	6?�4?�u&?�5�>PM�=�t����=m�g��暾�&������䣅��N=�����Q��;�?$=I�=��>?��=����l���eT�=�>w�?�C�>�ӵ>���nA���Y��ᾱ�Ž��۾kY�>L�>�?��D?�pB?��>�Q��묽x�]��s�>�;T>2�f�UU9�\(;qv>�J�=/)a?��?���|�*�*�f��6
>\�><T?�[�>�)�=�c=���=��G�˿�3���3��q������Ƽ�ֽ~��<ܰ�<?�D���
�UDE�3�,>٣�>�ma>Yk>�>��>�p�>�}U>XU!=�`=���<�����ʽ<�=U�J����������<E� �_����PE˽�&m�<�����--?U?������y᫾,O���%>&��>M��>G�B?��G?�=>��z�a���A��{����?�ʈ?,�>ৼ��Ѽ�̔�U��h��>F�? f>�f>���O�����>��?��F?��>���F�d�e��}�#�>9C�=�⽅��?�^?�3�@�����
���]�s����=����bN�Iؾ�$�c7#�8�����ƾ�꽵v�=�>3��?]����K�<�ھ�Y����l��J��+�>v6=�J ?���=S�&��*@�����s�Ѿ��_�u��<�o�>$	a<M�>wQ?�{!?x�a?�1+?RB�>`"�^A�>qc�=�*�>��G>�h�>9�>�0�>��f>Y�>�SY�y�*��K��u��G."��^��>��>��><{/>��	>҈�<;3�4 *��H���Ӽ��qǤ=c�>A��=�SL=�?�m�>O�T�5�ѽW�������3>q��=p�&>�ܼ��i� v��!����>X�2?n�;?ԅ�=��ɾ´���I�6��>�#?w�#?L�=	����=��P�־;e�>�B�'9���	���)�|����4�-��>��>"0��uY=�r�?��\?�l?,�t�~�"�-�6������i�5>c��>�֗>��z=�Z����0��|_���i��g�Xc}�u���ȿ>��>i�u>>@>CBP=���C����4��Ħ���ܼ�_>�
>D2�>�.�=���=�3��1?|����
�����9�߾���9�=zN!>l:׽�e�>A%����r�S ��n,�xL�>x��?���?�_?ѓ�e
B��>r��=[�>Bt
��v��i�=r���t��=���=������"Ð=�>͉�># ߽V?پ�����w�UEԿ�7�W;&��U$�ϳξ-����u�|�->F�����n�i��<���͕U��$�,����[��5��i2x�C�?�Zk?��a=����%��Gݾ�+��"=�)��Q����&�����⊆�����1����A��@!��{?j>Y��	���)���A$�����=�ڐ=�4?��c��ݾ�1��ѽIv>*J�>|�H���y�ژ��;���b?ʧ3?��4���ɾθ� X?~�?��=�`]=z�����=�6>��&?�h?�>�=���G1���7�Mʰ?�z�?�7;?!��,-��߾5��>m�H?���>�f�>�}o�H����� =gk?��?R�>/���2\�Ђ��{Hy>l�>��½�Z�>��>�L�=r��P���b=�}B��m��c=Mƺ=�o�=��y���X��X�=���>wh�>a�
�_����=>��Xm(��U�K��� ���Z�Oe?��!��a��gq=���<G��[u�X݇����>3?G�?F�v?A�X?=���P���Th=�}���k)>-?a'�=C�W<�I�>�j>1?	��8U�� x���)?g�?��?<�u?��Z���������?���g���<M>��Ǽ8@>���=�ץ�ߏr�c�=J}a>HOd>�^>�z>۷;>��
>޴���i��~#���wO���!����,�]k׾��d�j�eS��۲ʾL�Y���٩�Ħ����*�;���b��5w�>�6?�==?	�>�>	�=�I��n�=J���1־P�uV&��տ�~�S���[�l���j����ɽA7��;�>��{��Y>���>e=���'=>0�>�~�=���>Ds�=�]=ɗT>M5�=�>���= "�>��>W�o>��^����K�{��8�\f�4Q<\F?n	����r;=������ͫ�#*�>)w?C�>#��[�����M�>��>nW%�͐���u��`�<�M�>���>�ѭ="�d��z���Y�T��|�_>�
�>�u>���ɚȾbj�gE�=�7�>� پo]�=-�\>X�*?��[?��$?�H=��>I;>�p>�n>��8>I>���>	6?�4?�u&?�5�>PM�=�t����=m�g��暾�&������䣅��N=�����Q��;�?$=I�=��>?��=����l���eT�=�>w�?�C�>�ӵ>���nA���Y��ᾱ�Ž��۾kY�>L�>�?��D?�pB?��>�Q��묽x�]��s�>�;T>2�f�UU9�\(;qv>�J�=/)a?��?���|�*�*�f��6
>\�><T?�[�>�)�=�c=���=��G�˿�3���3��q������Ƽ�ֽ~��<ܰ�<?�D���
�UDE�3�,>٣�>�ma>Yk>�>��>�p�>�}U>XU!=�`=���<�����ʽ<�=U�J����������<E� �_����PE˽�&m�<�����--?U?������y᫾,O���%>&��>M��>G�B?��G?�=>��z�a���A��{����?�ʈ?,�>ৼ��Ѽ�̔�U��h��>F�? f>�f>���O�����>��?��F?��>���F�d�e��}�#�>9C�=�⽅��?�^?�3�@�����
���]�s����=����bN�Iؾ�$�c7#�8�����ƾ�꽵v�=�>3��?]����K�<�ھ�Y����l��J��+�>v6=�J ?���=S�&��*@�����s�Ѿ��_�u��<�o�>$	a<M�>wQ?�{!?x�a?�1+?RB�>`"�^A�>qc�=�*�>��G>�h�>9�>�0�>��f>Y�>�SY�y�*��K��u��G."��^��>��>��><{/>��	>҈�<;3�4 *��H���Ӽ��qǤ=c�>A��=�SL=�?�m�>O�T�5�ѽW�������3>q��=p�&>�ܼ��i� v��!����>X�2?n�;?ԅ�=��ɾ´���I�6��>�#?w�#?L�=	����=��P�־;e�>�B�'9���	���)�|����4�-��>��>"0��uY=�r�?��\?�l?,�t�~�"�-�6������i�5>c��>�֗>��z=�Z����0��|_���i��g�Xc}�u���ȿ>��>i�u>>@>CBP=���C����4��Ħ���ܼ�_>�
>D2�>�.�=���=�3��1?|����
�����9�߾���9�=zN!>l:׽�e�>A%����r�S ��n,�xL�>x��?���?�_?ѓ�e
B��>r��=[�>Bt
��v��i�=r���t��=���=������"Ð=�>͉�># ߽V?پ�����w�UEԿ�7�W;&��U$�ϳξ-����u�|�->F�����n�i��<���͕U��$�,����[��5��i2x�C�?�Zk?��a=����%��Gݾ�+��"=�)��Q����&�����⊆�����1����A��@!��{?j>Y��	���)���A$�����=�ڐ=�4?��c��ݾ�1��ѽIv>*J�>|�H���y�ژ��;���b?ʧ3?��4���ɾθ� X?~�?��=�`]=z�����=�6>��&?�h?�>�=���G1���7�Mʰ?�z�?�7;?!��,-��߾5��>m�H?���>�f�>�}o�H����� =gk?��?R�>/���2\�Ђ��{Hy>l�>��½�Z�>��>�L�=r��P���b=�}B��m��c=Mƺ=�o�=��y���X��X�=���>wh�>a�
�_�Fu�>����H�L�ǅK��g����侉�1��#?���64�>�o>>��g>�T����$M���<5�Ϋ-?宲?گ@?�]?��G��,���ɽ�g��?z�?��ɽݯ�;��]>}��>�>�G>_�2d���&?Q�?���?v�p??�|���տ%���0��݉���>�c�=-%>�?��Z�=�F=I��<ɿ:R�>L�~>�9D>;9M>��[>��>��>�݅���$�����Vo��s=����n�4[�����E�b�������f���A��A�ܽ��}���<�����+ݼ�����k>��?�?7;d>]D>�fw�����w��$�I	��������Ԩ'�Z�込�t���<�/~=�@����v��N��?�k=��=.`�>v�8���-=Y��=Y�=��!>���=�l>a|Y>��,>��>BH>� >�!k>�9Y>�q�=����׆�N2��8d�í�<��I?4�N�8����>&���̾;$�����>3�?^�P>/�'�s!��$r�`y�>ڼ[�$��l�&���2>�C�>@	>jt=�u���q�Jg�J=8Bz>�=�V��� ���!��=���>5�ɾ�Ƀ=�D>̙5?�l?E�+?6ZR=<��>�^/>s>R�h=�2d>��v>c]�>�?��3?@�"?�m�>'p�=��m�by�< $'=�\��=w����v��֫/�7~2<�&ؼ�Ai=Hz�<@Y�Ů`=쏻=��?<� P��V=-g�>Z�,?���>�>�0=�S<����՗�����QR�>�꼆�?�`W?@B?�0C>2IQ�"ͽ�I{=«�>�L>y�R�0�e�uB�>\��=2�@>� W?�:?���2�K���7O>��?�1?Ĩ�>��[=�M�<d��=բ��oпW������s��9>��>0�:�xν=c��=/
�J(��Nݵ<NI�=�EB>��>��>���>��=z��>ڎ$>��(�?XZ��ۤ�׏�<��<ꍯ<�R��J3>4�=���:�,�bFڽ3 ��7'�<{���lO*�o�����?ʑ?*҉<Yný�Pξ����O��޶>6�>f?K��>R��=f��TC��[+U��Ĳ�� ?�j?R�>��<;��H�ڈ�I>I?��>f,Z���>�/	�5�
?��%?b�?���>�}��Kㄿ;w���Ǿ��>d�_=�	���s�?��`?��P���w����?��h��E�=����h�������#�]�2�Lؾ��۾f�P���=Z��>ʼ�?'�z��q3=���gڗ�ť{�?���c�=2ہ=���> �>��7��獾�������?�A�p=���>U����N?S�R?�a2? �A?$N�>^m ?U���o?�/Ľ�%?��>���>�_�>��>e��=21��2_��������*���f|<�����[>�$R>-;8>΄y=��^�4�=7]<����ɑ��vn;���6<�='{�=���=��G>[<�>c�?p��>%���b���[��U�����N�m>�ᱽ�c��˱��鲺<�� ?:C8?%R+?���=�8����:�	�JɁ>�0?K1?��ú�x�����p}�ɸ߾�>�$�����������#�B����:B��>^�>� 
>�.X=��?%}j?�Kc?E��r�����U�p�s%S>�$&��_�>9��>�t������##���P�`�q���i�1̾U8���O	>��=>��%>R[_>,a�=�wS=���<�XO�/[��#0>�V7=�:y>� u>���>���=`�n<�h4�yC�� .?5�߾JҾB�D���n�ȷq<̊��֖>�킾93?q�U�	����B����@�&q�>���?���?]V?֛ýz��<S�s��c�=>K�=Dg}>_��=��<�����B��~>6�X�s�ל�>i��>#��>��J�k�㾇����0</�����,�� 꾭9F��,����ȾS�7��=��;��>���{	������½q�ӽ�)��;�$3����7�?�?�m#�Se����iT9�u������>�%Ⱦ
3��%���܉J��难[G�����8`�C.�/��TӾ�C>%��$K���)|�W4��\	��G���S?eƉ�t�R��8 ���:��m=
?>�����o�3+���@��2??��?L1��hR��ƉU>�]�>$��>G�>u7>PI �7���A;�q<?<|J?�a�� ��>�������C�?z��?��X?��
���7����v1=�b?(�;?��>�H�:���^�}�V?D�?]7�>��Q-��x����:>G�>VpݽѺ�> �>�Tw>��ľy�F�0H�=�sv��#�=y;�ݽ�{>�K)��5s����=��>,k>���#��~W>'���aV��6T�����HƾU���F�?sƋ�(}�>b�>I�Z>��@�����iE������B<)?���?��n?{�4?���@��`GK=����>�
�>,�-< ��:Ю>�Գ> ����q�ݵ��p*?��?��?$�,?*�o�)|��6�w�=j��/�оe��=��#X�>_-p=w��=��I=���=m2o<j�>�/�>�<>�n>4W)>̽+>��j<V������T�����((_�*06�|;�����<�� �!�\�M�
�����R������<���0�м?�~��x�k@�����`x>��	?U��>n��>_4=�6��'��Ɨ���q�+ɾ��_�þ�)��ɾ�g�����=��=-ɽP�1�ž�?���r��=�z�>)s�<�9�=Q��<0���ET>�9>I�=�&>��=Ew/>	B�=���=XS>?>�{�L����އ�e�Y���0�]v�>Z?�i�=O������X��	nQ�Yw�>�?F>s�C�g5��������>�������լڽh�����>>(>���<��(>��<�����U��8�n=��>�=���;K.n�RH�p��=�>Aa̾���=��e>Yq'?��n?N\0?e�L=�>�>�I>��>��h=7b#>�+>>u{�>NB?u�=?��+?��>��=ޫ]��f�<U�5=�*�����<���%j����u.8<�=���:G=r�@=e�t�B�'=�x3=�`<��<蜐<�J�>�Y6?�^�>��V>#�=�A}>�|�l��豾_+�����v>�S!>�|�>f_�>�Z-?ff�>�&m=����*ܻ��>�_�>1�n�{�h���$=��>�$=J�3?$M?��p���E��"�8� �Z�>b{=?�/C?���=�F��:K!���jӿY$�o�!��ւ�E�7�;+�<��N�u88ۢ-�����ʊ�<�z\>[�>Ewp>�E>��>OC3>VT�>�AG>_�=�ԥ==C�;��;:�E��M=#9�*�F<}�P�Ru���Ƽ^������[ZI���>��D���ؼ�?Ӑ?�a�=j= =�^������K�ɍ�>4?>�&$?�?+%�<b����^��G�Cƍ�ɇ�>m�K?��?j#���5������7˽���=�3�>P��>�"�mի������fu�TX�>�?Ξ>����e�>y��Q��o�>��=�y�Y��?ZFx?w����wѾU*Ѿ_9�7XO��q?)����<w��_���f���Q��e߾_�ξQw���x>ZK?���?�	��[��`Ƿ�l9��g�Q�6��;�'r>y0��?*|g>ߌ4<�
��X#�&�߾fH��H�D��[�>���!�?�1u?�m?EVn?�?�I�=�bz�.?4O����0?�H�>���>��t>F��=~骽V*���墾T~�����Rʾ���;�Iҽ��0>Y�V>�L�=ѹ�:����� >��t=S�ݽIΔ<�-=����&�<�H1>y��>^]f>�M?P�? y�����m�;��yf��3^�Q�=	�>7|�<��*�|M�+����>c�?Q� ?ǌk> ��� �L����t�>.?c�#?���>�����=$�:��{���h�>"�<t����#ྃJ���>����>���>�>s��=��?�)N?`dR?��W�2�΄9����_�=$Gp����>o��>ѕb=Sо!��+O��R�Vm�m������[>�&p>���>\�=��&>��=rE��h�q�Nvž��=�q�;Vة>(�j>'A�>�t!>�����Mྟ��hn'?���0�]��p�@�(�]���н�>�q�<H��>���6������20��p?���?�?;�?��p�a	D=C�Ͻ�*>���>z�E>��=(��1�ͼv�Ž��w>�ё������>b��>�1>z1Z��Ӿr�ؾS�+��¾��N�?%"��Ӿ�q��{_Ҿ�������Ӏ���ݽ�ܾ�V��s� ���ؽ��:��[��=��NS���H�?���?�Q�=�~��½1�����ྍ'�=������Rd���Q-�n��%����e���G���/*�#*��
��TJ>���Ɖ���R���>��>$aF>�P+?�ύ����X�"��?��lW>���>���`�z�������<��C?��%?�Bþ�ޜ�gj�=���>�D�>@�`>��M>�䢾�4�*�9>�aG?��K?$�r����z���Wo��5A�?��?�b?�,8�~�6��⾦d�Q�a?��?�K>�<;�о��P�H�_?��?O�?�s޾�v~�����`�>�V>��|�f��>t��>�`H>VU��r�V���(=����k>�pN��q�=��>��L�p���?<Ǎ�>���>u���i�C��>�.�U�c�.���ّ��$U=���=7�?-��N�>!=�>���=HP��̮w��3��NY\�ڥk?�޾?�\k?v�5?W/��́�"�
=q��>"c�>�a�>b.�=M����>��>%�<�@���$?�N�?���?^?��_��Mӿe��󳶾��!��=p"�=h�>>@߽���=�K=L���=>�po>꒛>�!o>�Qx>��T>¹<>��.>ˠ����#��¤��Ւ�CaB���ڨ�{g�Vv	���x����̴��������}����ᓽ7oG�.��p>������w`>{�>���>f�?r��>�)+>���`�{Uܽ+���yB���B#�������ҽJ��'���o����D�_�ԾS��>)'L��Lؼ���>M/�"L>�>��,>�z�>;��>�oF>u�>�� >2>���=��*>�f9=�p�>Χ齷����~I��r��
��<b>$4@?+[��+��-B��j�<k����?+%? �9>�i�弖��d���S�>}�>���;���<����M�:>�F�>�$�Oo>�+�=#��Z��;�RF>��>2�g>�x���ľe���p����>�־lM�=P�v>C�'?K�w?8?6?(�=>�>�d>6�>W�=2vO>kT>�!�>�?�}8?2�/?l��>m�=��[�b�#=<=�A�e�G�k���������iR<-l=��L=0�=�9<7\b=�7=&�8��;=��?��+?��?�l�>��O��b�f)����>��>�]�����>�{$?��5?")�>ą�>K@��1Ť�_�i�K�0�T�?f�<]}���!����3��"�>$v?�i?�چ?�ھ����^�>7��>��?��?YyA?���=F��=t��:h�8_˿v��7!5��Ԥ�����y;���ɾ��	iK��?h���n�.����ԕ>;��>z �>��>�Ԃ>�֒>W��>v�.>�����OϿ�O�����c��
>����G�&<�Jʼ@����_̤�)LԽ�kٽ��B�����W<(�>�S?��>�菉�~=�,�]#D�87�=�	?`�f>�cz>��E���ھ������b�:O�3��>2Ԏ?���>���옼F��<\���6�>:�q>��= �H>��'���X�$��>Ӱ<?�Q?(U>se�S�DH^��h�s�?Mv�:�3 =Tɘ?@gO?L'�f�<��7�TQ��ݾz��<vg��,��Xվ���N#��˾��� �5�2��=��>3��?#��=0Th��"���r�������zx>�m�����={�� c�����,�=���=d��>߽^>�Z =�	?�A?w�?m�2?�?��!?�
����.?uXS�[��>nF?��7?���>�+�>�ì>1 >Zi}���<����Tȗ��Ȇ=�J/="1=	�g>x�>��5��;�=�B���=3<��r���Ͻ�>S��=u�<��c�=ʝ�<'b?�[�>���� ��<�=��s�>`rC>��>�)c�F��/qq>
��>jn?�?��>5��������f:Z��\�>C�?��5?��?�3H�B(g�x�T�������>�=�>6S�3���g6��x�:@J�&��>�ƈ>.��>�4>�|?��w?,�0?��k<���QP��I�ʾ�\.�}f-��?�>4j�<D�3���2�>���4�V���Ǿ��a>T�C�zE9���=�&�>�C>��q�@�i>�5>L��5�=�{�=�Â<��%>��>Z	?�g�����=��־����h{\?u�<�������򉪾.��>i�X>�3�>�O���??<Z���~�|���+W �� ?���?��?�1L?)D����a�J>f�Y>#����D�|Wf�w��=m��7Ta>Z`)������v�< ,	?��D?���<f���o>�w������ -���P�;"���m��3ur�T{�<�Ǿ'jľ�V&�xpƽ�R��@ul;�*��=��4�1�k'���@z���?��m?`�۾�����/B��Z�����y�>���^��~3�sH�=;���f'b�h���0	�t�:�)��v�>�sh�������2���c��y���">O�!?9����B뽨��*>uN��iQϽ����͔�祇����<M?��B?-�N�K� �_do�$��>",G?��E>��x=I���)�2��>N<�>#{?�9��B����f���-=P�?���?�eI?`�m��3��_�b�U�t�? �*?���>�㶽�]���A���e�>�xT?�?�3l���_���6��$�>��G?�����>�@�>��K>��⽩Z��,s"�Y�ƾ�=T��=�w�����O�b��b�~=Fߠ>1�5>ɦ^�|ʶ��?ϊ1���~��Z�Q,���=�{��?�/3���>�ּ>y�W=ð�i�X��Ѐ���2g?ٟ�?�'V?g�:?�Y,������;�L/>;�0>@ļ>���J��;�>f�>�l*���l�.Z<��[?,��?�k@�B?� ���Gӿ1�����>��c��=�"�=&�>>߽+ĭ=J�K=����=�@�>W��>�o>�<x>��T>��<>A�.>�����#�ʤ��ؒ��ZB�> �����xg��{	��y�N��,ƴ�O𽾅������&̓���G����a>�E~Z�ԝ>���>�?��?���>�_�>C��R����=���ca0��2>�H�'�V�WB/�>���+3ľ���\w��̣�/��>D"B<[��=�>`g��<>�q>9��=!��>M�n>O�>�>��M>v,>Ϟ=���=乗="��>!��=�ڂ�&4i��A�����ԭ;�W?�V��K4���ND�A���t�����>D�?��+> |&�2U��eˇ�2��>
��񑝾4����a=�Ĵ>f��>���<O_�瞽�m���t�޾8=/�M>Ƚ�=���إ������=L��>x�Ⱦ� �=}߃>�)?��u?+�:?Q}K=� �>��_>�Z�>��=�<>�}Y>�g�>ok?�3?��'?���>_��=�2���Em=e]=��W���L�7���}�����I�?F::{��;ۄ<=�v=D'�=��b=�Zb�urE<�_0=�?V+)?Jh?׈�>Dͭ���P��m@�;'l>ǬU��D><G�>tІ>ȑ?|w?`V�>�T�<��8i%���o ?�>�ğ�(���͐���^R>g-�>��J?5r}?�ƺ��+���=��#>j,?�&J?��E?�U>���>�ž�v
�ڪ�������9��L����W<�!��g}r�>���xR��_)��gЊ<�&�>���>OU�>Vs>��<�ʼ>�?Υl>R�������Ľ('i��ב=��>�<v�ļ`� �=B�ѽ� ��l��׽���w��<����h�>��>?]0_>�Y��z�x�;�վ�������=xh�>�m-?�6?�D�K<m�P{���X���ܾ�A>`Έ?VU?p��[�H>t�̽t��?=�>$�=sp>���=p�=�M�=Y�K>��>�P?se�>�.���X��p��ྜྷq�>5F =����y�?�mQ?3p�S�ٺ�1�w[��v� 잺H7�<�װ����L�374�%3Ⱦf���	�,�ª�+��>0��?�׿=/#�<Ѯ޾uw����� m����=wֽЖ�>���=w��;f���^=����� ���3�>+�>��*�RQ?��?�oL?n��?�Z?'J?GǾ�+?�3�G�>9�6?h?�"6?8�>;mf>��">�	��D�>K��$/:����{�-<6u >����5e=Vּd�=�hm=R۽�qw����=���<���=o�����=��3>8?)�)?g۽�����V>�!�A�3>jd>�5�>�S�����xh�>E^�>�?�>s �>O�)>
��Ƿ���?�o�m>$ �>2<?�� ?GD>oJ�=�PV�Eچ��T�=4�>Bc=\�����¾�Gѽ��a>@��>�Q>��l>ew?׋?���>��t*G�%���w"����=k��=,5<??��>@m?F.$��sb�Ɍ��s�Cp#��A>$�<�$��dq�>5��>S�Y=�Ν<I�:���>���2yg�dS�������j%>-�>M��>w>�Ll>Rk"��־��k?��L����6o�Â���r�>7ڳ>.�E>�h|<�~'?�饾�A���̧��&�LG?�&�?�C�?�6$?í����־!��>�e�>�F÷�D[���&���3=�=���jB>�Ȗ�&� �������8���W>���>c�c�H�	�܁	�lm��Ʃ�Mn�����r���)�PQ����t�e>O����u�O�����vZ��=,3���CRi������ɬ�O}�?��?|D���>����zB�׻оݴ�>����_>�D��tN#��Y�������X�
ھ�p���J�%����>�b��
�����'���5�F�ǽ	�=��>?�_!�\��=��E�>,�>�=�j�t���-��֗��E?Z�j?�U����w늾��>�y�?f&�>%�=�^۾��;��x�><?��P?j^������).��}��;�?���?9??C��d�8�O�	��׽���>c?�C�>�x|�����ݬ��?SA?pn�>����,k���m�`��>��Q?TƂ���M>���>�̮>�c#��*���6%=a˯�����:>�������l�1�a)����=���>�܇>�}������Q�>u�2���Y�.t�T�� ��=@���%�?*%�I��>��>5̓=��V*{����X*p���\?8T�?}�S?�$?����$�%/<�9�=�S>aJ�>�J�=����'��>��>�@�*⇿�I���?%��? @� B?*t���F׿����-���:���#�=�D=�Q/>�
���=_�=�P�a���7Z>S��>��p>i;�>�U>E><6>�.����(����%����:�$���g���m��?�!΃�-��˩ɾ��¾ٛ`�Ί-�mm���F�����i����44>ϯ�>�?�?���>��2>O`���&�U������N/��6��pؾ�V��u립�Y���aԾ	����\@�V�?��H=c�5�j>�>k���HP>k�M>Z
�=�y�>҂F>��=�>�yQ=	��=�_�=D�>X`9=*x>1'�☿R+�gk~��8�Ba>0y?�[m�}��^�r�V��+ྗ�	?��?�=jA��y�������$I�>aܾ=���G���b>����=>�>��T=�-�=G�<P$�[���t�=iB>�Ll>�.�b���7���{��#��>��־�=C�w>�(?"w?�)6?�d�=�
�>hb>̼�>��=��K>�_Q>T��>��?{�9?VA1?���>cP�=}z`�0B=^�:=�?���T�Lȴ����>�%�^͇<n�1��G=v�q=�f<��^=*2B=��Ǽ�ܱ;�% =�?Z1?,�>���>2���\�Q�~�4�4M>�%>����?55?�C�>J��>i6O>m�*�'�=��p���[�q$?i0[�Z�w�w���eKŻ+V�>�?��p?�P?Fa����޾>���>=?��?w5?��>67>{�5����\�ƿY�ݾD�����Cq�����}������y��B�j�����=�_�>\��>�8�>��z>#��=(�?�k�>��B>�����Y��V~��8>��9=��=���F<�����<�=���sýU���Iн�X���<�6�}��>�F?�>/���2 ��1���I��>#q?��>(UY>������\w���~_�-�I�jn"?z�?�g�>� }�sܚ;y>n�� #=�zD>��L>�$G>���=�jV�}���S�]>�J>?��?L��>X4�;�O��[�)�"���>���<H�=�o�?�S`?v��������<���A��l���=�e�=ξ;�	�Sp8�� &�J����ZԾ�ȳ���=p��>
��?���=ꈽc�Ͼ�ޤ�Wx��AX�;��r>�Ҿ�$
�=`q�%U�>�C���t�uk=��> �>���<5??�l	?��H?s�k?���>��#?*�����	?R��ln�>�<?�?��
?��>b~�>�8>-X���ֽ)�f�|`Q����=#�������>=Ȏ>�7�C>~G<�I�<k��?��x�=~kE=���=3	�=9><V5>Yw?�?�m	��2�z�>S�����>E�>=�>�����k��J>�1,>��?�?\?s��>��<�f�����o�7��>���>��Z?�j?�q������fL���$���k> �>��3���/�i�$�L
6��{�>�F>��#>��=>�Ʉ?��N?�JW?7�9�@�;�!}{�+��՝B�8�h����>H�>�V�<C��C�$MN��!>����v��< J��M*ɼ܌�=%1�>D�=��d=C�F>
>��I�|-��_
>{�A=��&>}�>'��>���<Zԯ��q��@ݾG�H?+}��A����]V��Q�$>�B�=�9N>SX罿�<?�:���*�����1����>���?^��?Y�b?g���}�(��R�>��A>�|��D��/Ž���=�F"����>q���a��qTܾ�:�=�9�>�	(?-�g����
/��<r��C���i1�@�־��Ѿ�V�����M����@��Q���9���e���������F��=���B�A�l�����G���q�?Dz?G����n�=��+�7s� �i>Q�����T��`��5|�<iN��Y��/7ϾY����w��{�~�>}�����d<�gV��is�n_+>H�F?M��������(�T>q�>�Z���r���u���I���b?k7?VN��n�/�O�r��>.�:?���>F�5>�δ��q���>0�?mfV?v�V?���m{�Ɨ����?,��?~�Q?�
��u�+�p�!�"!�b�'?�H?9�2?-~<"��V&<���+?���?M�>�7������VA`���>��I?����&>�=wm_>�oN=.qM>WƦ��~��;��>�؄>�GY=Nv���� N��]��>�?X�>�1^��$�C��>�.�U�c�.���ّ��$U=���=7�?-��N�>!=�>���=HP��̮w��3��NY\�ڥk?�޾?�\k?v�5?W/��́�"�
=q��>"c�>�a�>b.�=M����>��>%�<�@���$?�N�?���?^?��_��Mӿe��󳶾��!��=p"�=h�>>@߽���=�K=L���=>�po>꒛>�!o>�Qx>��T>¹<>��.>ˠ����#��¤��Ւ�CaB���ڨ�{g�Vv	���x����̴��������}����ᓽ7oG�.��p>������w`>{�>���>f�?r��>�)+>���`�{Uܽ+���yB���B#�������ҽJ��'���o����D�_�ԾS��>)'L��Lؼ���>M/�"L>�>��,>�z�>;��>�oF>u�>�� >2>���=��*>�f9=�p�>Χ齷����~I��r��
��<b>$4@?+[��+��-B��j�<k����?+%? �9>�i�弖��d���S�>}�>���;���<����M�:>�F�>�$�Oo>�+�=#��Z��;�RF>��>2�g>�x���ľe���p����>�־lM�=P�v>C�'?K�w?8?6?(�=>�>�d>6�>W�=2vO>kT>�!�>�?�}8?2�/?l��>m�=��[�b�#=<=�A�e�G�k���������iR<-l=��L=0�=�9<7\b=�7=&�8��;=��?��+?��?�l�>��O��b�f)����>��>�]�����>�{$?��5?")�>ą�>K@��1Ť�_�i�K�0�T�?f�<]}���!����3��"�>$v?�i?�چ?�ھ����^�>7��>��?��?YyA?���=F��=t��:h�8_˿v��7!5��Ԥ�����y;���ɾ��	iK��?h���n�.����ԕ>;��>z �>��>�Ԃ>�֒>W��>v�.>�����OϿ�O�����c��
>����G�&<�Jʼ@����_̤�)LԽ�kٽ��B�����W<(�>�S?��>�菉�~=�,�]#D�87�=�	?`�f>�cz>��E���ھ������b�:O�3��>2Ԏ?���>���옼F��<\���6�>:�q>��= �H>��'���X�$��>Ӱ<?�Q?(U>se�S�DH^��h�s�?Mv�:�3 =Tɘ?@gO?L'�f�<��7�TQ��ݾz��<vg��,��Xվ���N#��˾��� �5�2��=��>3��?#��=0Th��"���r�������zx>�m�����={�� c�����,�=���=d��>߽^>�Z =�	?�A?w�?m�2?�?��!?�
����.?uXS�[��>nF?��7?���>�+�>�ì>1 >Zi}���<����Tȗ��Ȇ=�J/="1=	�g>x�>��5��;�=�B���=3<��r���Ͻ�>S��=u�<��c�=ʝ�<'b?�[�>���� ��<�=��s�>`rC>��>�)c�F��/qq>
��>jn?�?��>5��������f:Z��\�>C�?��5?��?�3H�B(g�x�T�������>�=�>6S�3���g6��x�:@J�&��>�ƈ>.��>�4>�|?��w?,�0?��k<���QP��I�ʾ�\.�}f-��?�>4j�<D�3���2�>���4�V���Ǿ��a>T�C�zE9���=�&�>�C>��q�@�i>�5>L��5�=�{�=�Â<��%>��>Z	?�g�����=��־����h{\?u�<�������򉪾.��>i�X>�3�>�O���??<Z���~�|���+W �� ?���?��?�1L?)D����a�J>f�Y>#����D�|Wf�w��=m��7Ta>Z`)������v�< ,	?��D?���<f���o>�w������ -���P�;"���m��3ur�T{�<�Ǿ'jľ�V&�xpƽ�R��@ul;�*��=��4�1�k'���@z���?��m?`�۾�����/B��Z�����y�>���^��~3�sH�=;���f'b�h���0	�t�:�)��v�>�sh�������2���c��y���">O�!?9����B뽨��*>uN��iQϽ����͔�祇����<M?��B?-�N�K� �_do�$��>",G?��E>��x=I���)�2��>N<�>#{?�9��B����f���-=P�?���?�eI?`�m��3��_�b�U�t�? �*?���>�㶽�]���A���e�>�xT?�?�3l���_���6��$�>��G?�����>�@�>��K>��⽩Z��,s"�Y�ƾ�=T��=�w�����O�b��b�~=Fߠ>1�5>ɦ^�|ʶ��?ϊ1���~��Z�Q,���=�{��?�/3���>�ּ>y�W=ð�i�X��Ѐ���2g?ٟ�?�'V?g�:?�Y,������;�L/>;�0>@ļ>���J��;�>f�>�l*���l�.Z<��[?,��?�k@�B?� ���Gӿ1�����>��c��=�"�=&�>>߽+ĭ=J�K=����=�@�>W��>�o>�<x>��T>��<>A�.>�����#�ʤ��ؒ��ZB�> �����xg��{	��y�N��,ƴ�O𽾅������&̓���G����a>�E~Z�ԝ>���>�?��?���>�_�>C��R����=���ca0��2>�H�'�V�WB/�>���+3ľ���\w��̣�/��>D"B<[��=�>`g��<>�q>9��=!��>M�n>O�>�>��M>v,>Ϟ=���=乗="��>!��=�ڂ�&4i��A�����ԭ;�W?�V��K4���ND�A���t�����>D�?��+> |&�2U��eˇ�2��>
��񑝾4����a=�Ĵ>f��>���<O_�瞽�m���t�޾8=/�M>Ƚ�=���إ������=L��>x�Ⱦ� �=}߃>�)?��u?+�:?Q}K=� �>��_>�Z�>��=�<>�}Y>�g�>ok?�3?��'?���>_��=�2���Em=e]=��W���L�7���}�����I�?F::{��;ۄ<=�v=D'�=��b=�Zb�urE<�_0=�?V+)?Jh?׈�>Dͭ���P��m@�;'l>ǬU��D><G�>tІ>ȑ?|w?`V�>�T�<��8i%���o ?�>�ğ�(���͐���^R>g-�>��J?5r}?�ƺ��+���=��#>j,?�&J?��E?�U>���>�ž�v
�ڪ�������9��L����W<�!��g}r�>���xR��_)��gЊ<�&�>���>OU�>Vs>��<�ʼ>�?Υl>R�������Ľ('i��ב=��>�<v�ļ`� �=B�ѽ� ��l��׽���w��<����h�>��>?]0_>�Y��z�x�;�վ�������=xh�>�m-?�6?�D�K<m�P{���X���ܾ�A>`Έ?VU?p��[�H>t�̽t��?=�>$�=sp>���=p�=�M�=Y�K>��>�P?se�>�.���X��p��ྜྷq�>5F =����y�?�mQ?3p�S�ٺ�1�w[��v� 잺H7�<�װ����L�374�%3Ⱦf���	�,�ª�+��>0��?�׿=/#�<Ѯ޾uw����� m����=wֽЖ�>���=w��;f���^=����� ���3�>+�>��*�RQ?��?�oL?n��?�Z?'J?GǾ�+?�3�G�>9�6?h?�"6?8�>;mf>��">�	��D�>K��$/:����{�-<6u >����5e=Vּd�=�hm=R۽�qw����=���<���=o�����=��3>8?)�)?g۽�����V>�!�A�3>jd>�5�>�S�����xh�>E^�>�?�>s �>O�)>
��Ƿ���?�o�m>$ �>2<?�� ?GD>oJ�=�PV�Eچ��T�=4�>Bc=\�����¾�Gѽ��a>@��>�Q>��l>ew?׋?���>��t*G�%���w"����=k��=,5<??��>@m?F.$��sb�Ɍ��s�Cp#��A>$�<�$��dq�>5��>S�Y=�Ν<I�:���>���2yg�dS�������j%>-�>M��>w>�Ll>Rk"��־��k?��L����6o�Â���r�>7ڳ>.�E>�h|<�~'?�饾�A���̧��&�LG?�&�?�C�?�6$?í����־!��>�e�>�F÷�D[���&���3=�=���jB>�Ȗ�&� �������8���W>���>c�c�H�	�܁	�lm��Ʃ�Mn�����r���)�PQ����t�e>O����u�O�����vZ��=,3���CRi������ɬ�O}�?��?|D���>����zB�׻оݴ�>����_>�D��tN#��Y�������X�
ھ�p���J�%����>�b��
�����'���5�F�ǽ	�=��>?�_!�\��=��E�>,�>�=�j�t���-��֗��E?Z�j?�U����w늾��>�y�?f&�>%�=�^۾��;��x�><?��P?j^������).��}��;�?���?9??C��d�8�O�	��׽���>c?�C�>�x|�����ݬ��?SA?pn�>����,k���m�`��>��Q?TƂ���M>���>�̮>�c#��*���6%=a˯�����:>�������l�1�a)����=���>�܇>�}������.0�>G:��?���ve~��#�٨�=�{�=��(?<'��j'>1�U��=�>�<0�1����>���%��^E?�=�?��X?��?�r����i�)ͼ�;<|e>�Ѫ>��ǻ��?��{�>��>֝(��H���Q!�p -?s}�?>� @jk?׎��eN޿߮��9h־�Τ���8>�jM>���>X?a=8�>i��*
�Fu��+R'>���>Ϥ�>x�>Ht>�:>er">����Y7�M?���长��9��g�L�N4���ݞ��⦾��7�������ܾ*���f���"�JEp���9�����F;An?<���>��>�2*>c^Z>²�>�H�H�,�Hc޾�x����у��\����^'����;�|$��nȾ���B����(?8֙�d�H�G	?j��i�7>���>�� =�
�>+�F>���>��>M��=�_>�? >�eh>$^�=T�{>�N�=
��@���f?:��WQ��k�;��C?��]��I����3��e߾O�����>��?=�S>~'�G���p�x����>�*F���b��˽}�c��>���>ޕ�="�л���"Hw��C���=�g�>(�
>��v��$��M��^�=���>����,h>�>Pa�>K"�?9�9?{��=�N�>�b>��>/V'>�e>M��=��3>g?��0?��'?/�>>^>V�`��E�=�,>+w
�����[���(�6�B�F�=+�[���=��->�}r��Dt�n΅=����$�M=��?X$E?��>��?�b�o\@��@A���վwm�>u,�;�G>���>s�)?�4?��?��D>KyZ�*��a����>�>>�?x�����J�>��s>�jm��m_?�\?���=�Ğ��<1����=�?�#?��?�M�>�X>@kݽL���mӿ9$�u�!��Ղ�"(�U%�;͐<�ZL��&�\�-�y������<r�\>T2�>�gp>�D>��>�53>y_�>��G>�\�=��=7�;O� ;�G�*M=/��*9D<�DP�����U�Ƽ`ޗ�����K��%@�*����׼��>�;?�ʚ<	悽~m�z����⾵�>zE�>�$?�?so����E�� 9����+,�>�QO?cO�>�	F�<->�$E����i��>���>��k>��/��<�L]�؏H=Շ>�~!?�{�>�e��y�y\j��a�-t�>
(o=��i�,�?^2]?�3/�� ��P���8�1�
��H�����=ġD��mk�:q<��[�f��  ˾c�_���=��>�?�D��_��>V�(�n���OV���ņ�[�>!�<��>�y�����d�B�,%
��ϾX�Y��%<<���>E�=>���>��"?:?��a?m3?���>����	?[��=�C�>F�>��#?F?��?�m>pZ>�_3�N�}b ��Y��C��=��=���<e�=�
>V�"�4P��N=�T�==��=��=L��<c���Jm]=�k�=ι>�r)>H� ?��/?6q������>�F�Wq��X;��>X��=�
���@� ��>Gt'?=\?u��>��5<�3�Ň�x�p=�%?�v'?y!
?gR>��%>�׾!`��?��;���>�<�:q�q�[���G�w�ཻ��>�>�n�=�a�>�}?��??�6??򹻽�'���i���:���=��o>��>j½�R�=V���ؐ��k�]�D�$ ��ԍ=�sؽ��Ӽ��=\�>�U�=���=�Y�>��G;;G�.�����b�>��>փ�>k�?
�>�4��b�[���D}8?��վv��c��7�о�r��ת>��>�_���?���i`�x㻿&�D��#�>Q��?��?舍?�J���@G�DW>��>��>%�|�5/���7�<$T��+k>�{�=�,��:��_(�=dz2>�vM>{,�����b�#�Zc/���п̙^�H��nҾ�Ց�#=�������`�샾�D.C���֦4��w]�%�����t�V뎾b��ne����?�l�?�Y���$߽k:����c$��=��D�Y�-�R���|���'sľ����61�q�@�0��k���N!=�>������J�� )�z�Z=n>{zY?f����W��n��%j�>Ђ>;Ɗ>e9%��i��C����7��?7�Y?�����L ��z��+�>��?�0�>�e�>���gG0����>'%W?�-?�7�����h�;s���ĸ?�x�?Jg6?[V��@P�����ő�nM?>?'C?���	aվ�H���'?�>?[_�>.��8c��N#�s ?��x?V��]U?>T2�>C�g>�'��t�������M��@+Ľ:�z>1�����D���H�����=A�>'b�>WD���Ե�2}�>6w׾�����k�$���q>�"�<�L@?t� ��P�ms�>��?�v9�6B���|���+��rJ?jS�?k�m?��+?���{��怾�d�>t�)>���>ֵ@>s�ɾ	@u>���>o�۾-8�����nn?dP�?��@�G�?	��CGӿ��$��������=%�=��>>��޽�ɭ=z�K=�˘�zZ=�y�>���>$o>G;x>p�T>ț<>��.>o�����#��ʤ�1ْ��[B�� ���wg��{	��y�����ȴ���O�������GГ���G�a���T>�]���">���>��>�S>�\><��>Ä�� R���ܾ�p<�Z@�i����&���"�-�4�#>�v�D���9x���-�m�#?v�6>�����(?��=u�7=�ԭ>R�x<3j|>S�>M?G��>�qi>���>���=r7&>w��>�=2>���=�N����z���N�)��f��DB@?�`��;Ǿ?�O�����爨�өl>A?�>�3��*��܌��!� ?Vg=�lz�q[��S�.�j>dڦ>��>�Ӄ�FN;�7����fP�=>�>�q=a	�����=�d�=}��>�+� �d>C<�>�ʼ>�?+�1?d��=Hu>�9�=��>�;>7�y>�e^>4Q>�6?M8?�*?�\	?v^�=�����+>d G>rdP��$F��w��0�.�];-|�=�Oؼ�5�<!m3=�-/=i�=�/�=C���j�����=N�?�G\?���>�ڴ>)_�9~9-��|u�/��{r�>Fw�=�@�>uGe=F�&?q+?Y��> N><M��mS���K����>�0>�-[����4�Ӽ�l�>��=�+?t�B??I�=��,�0�!�{ά=��?�G?�6?(��>�\]=Q��<�l��%߿u�&�����7�<����V�JIg�
����a������@���=Ҟ�>��>���>ʍ>�$�=��I>4��>��">��=�߼�@�<�E��j�=��=�^佱�Y���=�տ�㳽�B�OL��Vz����N�,=��>9b?�x�:�}�һ����_��}aP>ѳO>��?%��>�+��D���a�K��=���`?r:G?���>�Wܾ��P>\�{=�W>�E�>��>��="亾h2N���Խ���<�1����?�'�>�d���y~��u�����B>eV<=:А�r��?ȞQ?�/�;������L�M����ѽd։=�/Ž�n��}� ���W�`�l�r����gG�zJF>/̔>�a�?��:Qƽ�U�d䩿ˍ��B����R�>���<%�<>�<�=�f���s龶�!��Q�:�M�� 1���B>Dx�>IΪ=��$?w�??��H?8$?t_Q?�1����>|�>��>kb'>{=?\N?p�W?�Ի>j�%=����HH�Z�Y�{Ѥ��m����$>rY>�!�=z�<���=��=?���ܓ=�`�=��Y��I�;3��bz�<���=��C>zz�=<>?+�%?�ʏ<��{=�s�=��<Y=Ƚ7����*�>���=�.;�R�h���>�t?�K?��	?�!Q��7���;��E�:Խ{\	?��*?%A�>-�=���>�˯�5������<���=9)\>H�_���un���ͽ��>��>X��=�5�>��m?Q�A?�!:?�턾n�X�v-C���'��zM=�>@ܑ<�ޝ���>����d*��m�t�2W����]�P=7��5�<R0 �d>>w�f>��̼yI2>�i;]�`�ecC��9���S�<�?\&�>�?�'=Fa�z������T�H?]����M(���(�|�'�2I�W�E>r��>|�ƾ�3�>�؏��j�Aǵ�eJ���>���?&��?��?R���dT���_�>t�?J�?>��������^̽/i����>�~�>�`��`���=i�=w�>q��+�ʾJg-���(��ݿN�x��$ʾ�n��K���Ҿ�M��P��;�o=V���al���]ze�����r�=�V��S�Iͭ�q��n��?o��?AYC�bp��\��4��Ծ��d>�kн�璾�u侑(;=��ܾz��g��
���<�Y:.���(���+>y5���o��o4z�//��SF�	%8=�TI?Up1�j��B�s��>g7y=38M=���_���[���aO�MW?�]V?�2۾����ɾq�>"�Q?���>(��>�C���!|=q�?
�C?�?��W^���?���f�=h�?%��?��??E�O��A���X���1?	�?a��>��l�̾�L�n?x�9?���>_!��h��:���>U�[?@PN��jb>���>�=�>�/𽋸��F"&��7���ۅ���9>�j�����Sh��*>���=m�>!�x>�"]����)(�>�����⋿��f�����SD>ב��&X?s����=#�~>`Z+?��;�����q�����<��=?/߾?�m?X�-?�:�\x� XL���>�?.��>�%;��澉'>: ?��ҾÂ��)J��@-?(��?��@|�?vM���n�#4��Ѷ������V>;�=X��>R{�ҽR.�/r���iֽ�@>���>��Q>d0O>�>��=�+�>����F�!�Yɦ��Y��K86��Q���"��^�,���Q7����*�+V羸�Ӿ\-����E��'���u����^��(󂾅�c>���>J�/>��<?VQ>���>���0"������t������D+'�)��ߝ���\$>���[�ܾBf����7�OGe?Z�O>��q��	?�ǽၺ�;�?21�=Y�=�S8>`��>h��>��=�խ>�~�=��=s�a>$�{>�̊=����~^:�
S�&�;Q-C?3�[��ߘ���3��h߾������>�?�R>-�'�t����x����>�iE��c��Y̽: ��U�>R��>p�=��Ļ;��0v�G��B��=c��>��
>}@q�&���q*���=j��>�����A>�x�>�>E��?}78?�#�=f��>5xP>z�>{�=;�i>�&h>.6o>lk?p4?�!&?[��>��=������=���=��]�7�A�����3�r�[=���=V[<~t�=���=�X�=�����=�RW��P��=!�
?� ]?n��>��>�I�B7L�wҀ��D��!�>���Ii�=s��>��0?ɼ�> �>��=?¥�1������>L̈>�vf����ؽ��rm>�o�=a��>q21?���>�,�<��f��@l>vZ'? �+?z�!?��W>t(->]��7��@�[�#�R(���=t�>�
>�Ϟ��I=x�o���쾅r��U��=j��>�?�>�57>��>J%�=Ag�>�]�>6?@>����5=�j��T�=G��P9(>�;>�YɽM�dݼ܈���0��n=����a=�҂=`�X���>��?��=j��΃w��Y���۾�yg>|֬<�X�>ͳ0?�j>��(���s��I���H<���> �)?���>n�d�D�)>	���0�	>Qܷ>VR�>��m>�9��'����콎$D>p��>~>��T=bȂ��h�[c �JH�>��=�jL���?��i?�E�'M<���֟E�N�������">�X�&2���8���q���:z������wU�=��>!�?f(�GV���z�=�=��Nlz��Z����$�%ڇ:mͧ>h��>�fԾ=��7������;�%��)Ƽ� >#�>{�x=��2?_rG?�*?m�?�i?��C�|�?\�>��>C�>sI?�Q/?�3'?�r�=է�=Osڽߡ#� 'ӽ���|V�<�6��D��v�=��>!&|>��/=8!>��1>��;bO��0��<��o����=	l>�V>�t>��
?�q,?c_-=�
�O���Y8 �Ú�����;,?��?8�¾����?�h?���?=��>*�D�1��v���0Ծ�*'��f?E0?\ˬ>4Ch=���>e�5�!}¾����=���=���ʄ��Ҿ�A;��|>ǐ9>v<>��>U�c?��K?K�Y?�ʺ=��C�	�&�Kw��N`�8�I�a>���>	�>z�ʾ�پ	<z���b���*���=H<�β�<"�=!Lm>�,;>M�ֻ!�>�r=��|=_��g����/�=�>X�>�?�<�ԁ�����B��R?E셾TM��}I��=�	Q>�2m<a�
?�����>xK�=�S�~C��o~J�&+�=���?T��?%~�?QC�2 �i�>\��>q�=>]���Ҹ�e�M�$�=��>#�������>k�D>e$=]�����U�*�����{���D]����ߙžbN��#Pо�Q��a��%�Z�3���k�'����4����*��y�������u�������I��,�?H�?nP����U��Y0�J\c���!���A�n��e������s^>P	�U��&� ��q=�b�N�_m"�z����V>��ýŤ���g� +�����ԽJzD?X��l�־�5�͸>�2<0�=���ڦ�eF������k?�F?.~���� ���U��B�>�(?��>��?g(����!=���>N?{'?Ye��G���?:�X�G<>��?
%�?.�??��O���A�E����)? �?���>�ފ�2�̾
�?/�9?q��>�#��d��*��	�>��[?�^N�qb>\��>�)�>j�ｆ���=�$��L��������9>���>���Jh� R>�O�=[�>G�x>�]���)(�>�����⋿��f�����SD>ב��&X?s����=#�~>`Z+?��;�����q�����<��=?/߾?�m?X�-?�:�\x� XL���>�?.��>�%;��澉'>: ?��ҾÂ��)J��@-?(��?��@|�?vM���n�#4��Ѷ������V>;�=X��>R{�ҽR.�/r���iֽ�@>���>��Q>d0O>�>��=�+�>����F�!�Yɦ��Y��K86��Q���"��^�,���Q7����*�+V羸�Ӿ\-����E��'���u����^��(󂾅�c>���>J�/>��<?VQ>���>���0"������t������D+'�)��ߝ���\$>���[�ܾBf����7�OGe?Z�O>��q��	?�ǽၺ�;�?21�=Y�=�S8>`��>h��>��=�խ>�~�=��=s�a>$�{>�̊=����~^:�
S�&�;Q-C?3�[��ߘ���3��h߾������>�?�R>-�'�t����x����>�iE��c��Y̽: ��U�>R��>p�=��Ļ;��0v�G��B��=c��>��
>}@q�&���q*���=j��>�����A>�x�>�>E��?}78?�#�=f��>5xP>z�>{�=;�i>�&h>.6o>lk?p4?�!&?[��>��=������=���=��]�7�A�����3�r�[=���=V[<~t�=���=�X�=�����=�RW��P��=!�
?� ]?n��>��>�I�B7L�wҀ��D��!�>���Ii�=s��>��0?ɼ�> �>��=?¥�1������>L̈>�vf����ؽ��rm>�o�=a��>q21?���>�,�<��f��@l>vZ'? �+?z�!?��W>t(->]��7��@�[�#�R(���=t�>�
>�Ϟ��I=x�o���쾅r��U��=j��>�?�>�57>��>J%�=Ag�>�]�>6?@>����5=�j��T�=G��P9(>�;>�YɽM�dݼ܈���0��n=����a=�҂=`�X���>��?��=j��΃w��Y���۾�yg>|֬<�X�>ͳ0?�j>��(���s��I���H<���> �)?���>n�d�D�)>	���0�	>Qܷ>VR�>��m>�9��'����콎$D>p��>~>��T=bȂ��h�[c �JH�>��=�jL���?��i?�E�'M<���֟E�N�������">�X�&2���8���q���:z������wU�=��>!�?f(�GV���z�=�=��Nlz��Z����$�%ڇ:mͧ>h��>�fԾ=��7������;�%��)Ƽ� >#�>{�x=��2?_rG?�*?m�?�i?��C�|�?\�>��>C�>sI?�Q/?�3'?�r�=է�=Osڽߡ#� 'ӽ���|V�<�6��D��v�=��>!&|>��/=8!>��1>��;bO��0��<��o����=	l>�V>�t>��
?�q,?c_-=�
�O���Y8 �Ú�����;,?��?8�¾����?�h?���?=��>*�D�1��v���0Ծ�*'��f?E0?\ˬ>4Ch=���>e�5�!}¾����=���=���ʄ��Ҿ�A;��|>ǐ9>v<>��>U�c?��K?K�Y?�ʺ=��C�	�&�Kw��N`�8�I�a>���>	�>z�ʾ�پ	<z���b���*���=H<�β�<"�=!Lm>�,;>M�ֻ!�>�r=��|=_��g����/�=�>X�>�?�<�ԁ�����B��R?E셾TM��}I��=�	Q>�2m<a�
?�����>xK�=�S�~C��o~J�&+�=���?T��?%~�?QC�2 �i�>\��>q�=>]���Ҹ�e�M�$�=��>#�������>k�D>e$=]�����U�*�����{���D]����ߙžbN��#Pо�Q��a��%�Z�3���k�'����4����*��y�������u�������I��,�?H�?nP����U��Y0�J\c���!���A�n��e������s^>P	�U��&� ��q=�b�N�_m"�z����V>��ýŤ���g� +�����ԽJzD?X��l�־�5�͸>�2<0�=���ڦ�eF������k?�F?.~���� ���U��B�>�(?��>��?g(����!=���>N?{'?Ye��G���?:�X�G<>��?
%�?.�??��O���A�E����)? �?���>�ފ�2�̾
�?/�9?q��>�#��d��*��	�>��[?�^N�qb>\��>�)�>j�ｆ���=�$��L��������9>���>���Jh� R>�O�=[�>G�x>�]���2}�>6w׾�����k�$���q>�"�<�L@?t� ��P�ms�>��?�v9�6B���|���+��rJ?jS�?k�m?��+?���{��怾�d�>t�)>���>ֵ@>s�ɾ	@u>���>o�۾-8�����nn?dP�?��@�G�?	��CGӿ��$��������=%�=��>>��޽�ɭ=z�K=�˘�zZ=�y�>���>$o>G;x>p�T>ț<>��.>o�����#��ʤ�1ْ��[B�� ���wg��{	��y�����ȴ���O�������GГ���G�a���T>�]���">���>��>�S>�\><��>Ä�� R���ܾ�p<�Z@�i����&���"�-�4�#>�v�D���9x���-�m�#?v�6>�����(?��=u�7=�ԭ>R�x<3j|>S�>M?G��>�qi>���>���=r7&>w��>�=2>���=�N����z���N�)��f��DB@?�`��;Ǿ?�O�����爨�өl>A?�>�3��*��܌��!� ?Vg=�lz�q[��S�.�j>dڦ>��>�Ӄ�FN;�7����fP�=>�>�q=a	�����=�d�=}��>�+� �d>C<�>�ʼ>�?+�1?d��=Hu>�9�=��>�;>7�y>�e^>4Q>�6?M8?�*?�\	?v^�=�����+>d G>rdP��$F��w��0�.�];-|�=�Oؼ�5�<!m3=�-/=i�=�/�=C���j�����=N�?�G\?���>�ڴ>)_�9~9-��|u�/��{r�>Fw�=�@�>uGe=F�&?q+?Y��> N><M��mS���K����>�0>�-[����4�Ӽ�l�>��=�+?t�B??I�=��,�0�!�{ά=��?�G?�6?(��>�\]=Q��<�l��%߿u�&�����7�<����V�JIg�
����a������@���=Ҟ�>��>���>ʍ>�$�=��I>4��>��">��=�߼�@�<�E��j�=��=�^佱�Y���=�տ�㳽�B�OL��Vz����N�,=��>9b?�x�:�}�һ����_��}aP>ѳO>��?%��>�+��D���a�K��=���`?r:G?���>�Wܾ��P>\�{=�W>�E�>��>��="亾h2N���Խ���<�1����?�'�>�d���y~��u�����B>eV<=:А�r��?ȞQ?�/�;������L�M����ѽd։=�/Ž�n��}� ���W�`�l�r����gG�zJF>/̔>�a�?��:Qƽ�U�d䩿ˍ��B����R�>���<%�<>�<�=�f���s龶�!��Q�:�M�� 1���B>Dx�>IΪ=��$?w�??��H?8$?t_Q?�1����>|�>��>kb'>{=?\N?p�W?�Ի>j�%=����HH�Z�Y�{Ѥ��m����$>rY>�!�=z�<���=��=?���ܓ=�`�=��Y��I�;3��bz�<���=��C>zz�=<>?+�%?�ʏ<��{=�s�=��<Y=Ƚ7����*�>���=�.;�R�h���>�t?�K?��	?�!Q��7���;��E�:Խ{\	?��*?%A�>-�=���>�˯�5������<���=9)\>H�_���un���ͽ��>��>X��=�5�>��m?Q�A?�!:?�턾n�X�v-C���'��zM=�>@ܑ<�ޝ���>����d*��m�t�2W����]�P=7��5�<R0 �d>>w�f>��̼yI2>�i;]�`�ecC��9���S�<�?\&�>�?�'=Fa�z������T�H?]����M(���(�|�'�2I�W�E>r��>|�ƾ�3�>�؏��j�Aǵ�eJ���>���?&��?��?R���dT���_�>t�?J�?>��������^̽/i����>�~�>�`��`���=i�=w�>q��+�ʾJg-���(��ݿN�x��$ʾ�n��K���Ҿ�M��P��;�o=V���al���]ze�����r�=�V��S�Iͭ�q��n��?o��?AYC�bp��\��4��Ծ��d>�kн�璾�u侑(;=��ܾz��g��
���<�Y:.���(���+>y5���o��o4z�//��SF�	%8=�TI?Up1�j��B�s��>g7y=38M=���_���[���aO�MW?�]V?�2۾����ɾq�>"�Q?���>(��>�C���!|=q�?
�C?�?��W^���?���f�=h�?%��?��??E�O��A���X���1?	�?a��>��l�̾�L�n?x�9?���>_!��h��:���>U�[?@PN��jb>���>�=�>�/𽋸��F"&��7���ۅ���9>�j�����Sh��*>���=m�>!�x>�"]����